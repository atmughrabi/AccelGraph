// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WxZYFqbwTqPNZpNaS6dzMEbR7apyORIQXqnaknkBcAwohbvVEZpquvh6blUa+mUO
oTR3w6sfwme755I+KNwUl4SRNaF5JrpH8EtxjEPnsc1ZGVld5ogkh7PZ+wZF8gup
wVxxYufT9zCKSOsIlgp0l8lJ1hVWo3AH5wbN1/8iINg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6992)
wLEa6srcl/zY7R+kr2cC45/5sIXWr+44DDmDiLW1wPLumgnBH5rc/iK5jOgzFwpF
NA6tP6ypcqKxTYDOQ0KVKheelV8nokJ7CeqIzuqwZCxU4eduBBi9YGSqlkL6tDvo
cD/gYZYGI/FYp5hyryLAJzqDUUSSbSDOMDtQmO4+2cJtC/P2WTZ1j8jkuSa8BBx7
2A2FndScrKn342a02MlDiI4sZMYT+8soYeBTM1B2IJF1Q5wW45o4Iv11LkHOOjnA
VvfwyPOejIzUMK0Z2EsWZ3cUcFNk7KzXQjt0aNqivxitpnJDJaX7Bat/QgV6gNgl
qcvMoe3664FejAwHzf9xSxUel7a1Xp/6E74wnc/DzMe+U+sRGREVsMqk/Gobljqv
WSadF6JTf9YaHVw+WmUP3NNaUJtWw3zpMtCTBz6FcAlhgejcNA00P7COQtSZylRq
PPeJ0BcqfGzOmG800FakGYdg362Ky3ijNfUClYdSPMIRLhuBLoy9/bRzZo34WOAJ
vKXzlbTeb/Wl9UQio+i7SGVPFTtAHWg55e5jo3FPuAn4PIl5jtw5m2AVPZFvYJJt
0VNprvtj6/MGMTnEZ0RWolJbynA5hIQNPmXOlaVJSnlRR6sL7U5LJD7Z3b0d5RdO
Nu5OrJC2LbocHPBvb5EfYyXMe1fvG0qp5ychtNYw7g/ezgHIPQk+BZqnOhLVZgG8
d4cLgJt1ik3UatBMBGyxbWkccrbBXEKWc99JRL9xoncubdnaOTQ9CCP8ie647VGc
86bK7OW8BeK3ibNAYtxDbomoKqqMtfwELZIT8OGNp7MpEWVR84vA+JHKKGuXefev
eQCcv00BUa5jtpsjz3z+CdIGlNCOqUz8GGpNAtc5lRoDFCaFfQ9THmchPNzSkpK5
Fke0P5jied1WgJBJAkkKRuM/vBjZMkz01pcAgvw905QLaGyTIXzXwbQ8mNYwhXzM
/1zjXdFB6rdbQT2Ds5awlUExIP+yLRGm+iWS733FmwQEmdpNpHo8YZzpg7zO3Mqw
+THapAQtQxU2qXw2O2gv+Kzq7KERNjndtB9b+GLcDgeY/K+PFNtJK/EYBbgZMZiO
Dl2aAdh7K+FkidwX6cnuT8uQIXqXNLB75tWx75FF5k3Gj9YacmslECi19TdOEcc5
9u4r2GmGEtWM9BdKJIKWg5y0wA80JNbN4e10vvhloqYklsLX2XjmOF0gQZc/IP2c
Ohf5f2dXR0FESil060vB+dykm9YU9OB1oArPJD3aLPFHEbVpcAiwFuBok4qmm+Kz
kbZrg3hHW772yxm/hl43RrzYoEFprk3tOO/S+ctRbI1DY24BHdYLFJfHvw7h/Y96
oCLSCBDsEowap4/D3Lucfxmv8CVFMZV4jbPK7mZ1r1Qu81f31++j3DFa6lhn1+tL
u906U+q+kPFdkNIh+yJuBv/zQL/9BN++LI97ocyS3vb6/jtr9tinMhIJWYLxB+08
2QqvOlKDYXgUBHaaJuOUbCOPAVZjt0uOqRyIL7k/+aCGHiLP1XZpWmipixHDVHgh
5Fk1Q9yUuAXj35WEAROzFjHnQ8j36vbVypvzt+3JN4wFJN/FwMvKKf7X9Y4eBq/e
uykv1dqGQ7FSo+bVbrYzvNwrmbCPz5RR5/xw9/0wLOFFSJclcFmIzu1KkawCuZTq
Vb9k4vBxsq1FdMo68cnGqw+LKsasCSkHHWwTeI2u3FJ+yBvtsaA4Pt9ShfrA4/Zb
ootXbU9+df/FZjx43PCcmqvMxXxIJehooVr52jZjGwHI/j7X7AEZE25Vme4JIq52
jlGvv9UUpGRxtZbEATyCfacUMGUQKEFL2bt/CpCHxoXAjv8wHL+EMIcVluzVYn5H
3sN/GLomArBtvy2oL5QxiP8ZxuWwiv+2Uzx/lb3Us9qwDrwjEGvacVWa2OC3l/cQ
dZp21FyoP+M2sGnHl7u3sqVlfwjXLpNpm8BeObRGbuS6fg+FQmbun0wO4LNvPvx2
2x2tOw2WwiyMMKoKTvnrAUXjffnbGGV+9ud0ZeYlyauyZz63tAgjfE1mu0imwOk1
jpmTMtXMITnyYtZwhYnOrc0D+G8nWKfe3N0v5QFaT1bQkptsYi9eFz69tJhaWRJi
ENmXSM0iDoQj877ahe3UOPkT3SGufZtXryETzEco6TUR0i0Gd2k1jQtUmo9esiEI
8GD9ZNNvYUwkTPSQM4mD7dlihDI7R8kKFJYxFG2CBTrelqEPy9XMounvpaEknl97
103KbcY2Uj6x/PdA7L+bgF0u1mghrLq2GQnDaFAr+ZqZr2hadwOrV0R+NgT9h2eT
jrhfivROoCeZT9GwxkKxotQ2qJrVmn8sG/LgqOKWa06TBu/eTnQNRFVurIlfmR0G
Jf/tfmUEE9QrCuLJvOOOHv10qSOoOr9s0h3F4gTZ9hizSPlt1gE1lvi2hIdXOuO8
2l9dHKiNFqq8RiJNPYKZUmA+B9qGf4tfymUdQdD/YaLJViFseILKxelPn5+PPiq8
HT4lQBc5MroG5hd87FXSAiNTbFexCi5JA0W6jsdUeld8on359GKsHUJ6cm8kSMZq
0yN5/eCuWcQx8ezHQrYIkY1PIgyj00khqAGagYtpyp35xLFBwiY3kRbYPMhCfFh4
McERq2UteCzCKwMKhQ/kGiK57CB+hywJODWEXkhtUfE3XM65I1zn++8W1S/2peAd
R/32SfRpRS0cXdK6rXwuZ7Yb72dbGyxr7amDUvUy8jxsOepjzC45XY6UUl61FDLQ
3KTlq2GH9HqML9Jii8tQst6NElRrjCFCTm0DisnhFmrTyeFcw7HfWDi1XWHE+HYQ
QfH/9deZTOLa6kVQ7JPu7fMV6O6FXv2uT4aqoH4OS63bPkdGNt6gy9c7KU1axW+p
nv/ovsLMdjO+Ia80QAc2p9eEZ8oWunSh8O2MFP84SciNeMMraEQzSMCpUwM85GM2
kDXdhFMkQ43sKkKP0HLLN/o2p1bJDA9rPSm1WnWkpXblkAw7BD2XOui7xNLKymG1
cQXOIstV1GjBGbS8WbJSKsZStFkv/xVVwRXvcLGqqMwcKNvFOJhuH3/MWiGqQd2o
7mFfKCHok0SHi30K7YnryrVuHP/MnV4KE2KkRDyABPpJQOWxwEHpxkXcD8rhwjuG
DOI1GUDBRItRghp3LRJOvVNFOK1sdv9EttSL4G+Z0zh96K8wHeqF5Wparq6uzYhO
d1aE9fv77cun3nR1R0uEf0LxRjy4kYaSwnYQU/YtFdjLUQi0NXge5mzYTMMoc/sM
fR5xndUz1CfzPKd3tKFrsLjdctRbSzioh86dnh18kFnusHDs67UG0H4BQ72EFhvS
PdGe+uOzmdha4Cs9xA3Utz7xjImZuUJOYYOoHA5aScswh4K8dv5B6gZGkJT/8CHg
PqNn5WowcEe0j77kJCiA2DsIkEihZ36tySDdqsqoabQzEWaUDI72HGNQVbhNwAQC
cGmVlA1mZG5wAaDkfQhCXXrcOXkStdg/oRgy2o9+jWKcr/zuLVshZQci2krf5Gzv
bcMyDrEAolLZLGsTbKdVeNXc8P+9qnyLV85yCOifH9sNjyEzr0bdcYbD85nq4e8p
YZLVWASOG1oDc+8KwZR0387Hfcsg5QBH+/GTywhzY75jGWUkTCTn9PZTHuHTIrv/
d2IhSFUvc2q7E3ohc9PRx3+iP2haqmJ2fIWpAi+PTwf9kdUfCVRkLz4U7JsdUW2x
qPvXK3SpI41Ieuvz0D+C0bmtXWuR9p648AnYd4Huc6KnV+ScT0YxibsM8OBQ/70u
yFAznVtsW/tgJm4xH4KeiLYgvkrOgHwx75IIFyfVRN0lPSbP7dXfOI+uTkx1ggBw
2HD7ksUmRugSggw+Eb9zg/IDUlYpyEvp7PAPjiXDyFt4bi9rwJ5EcCeRlqYQofEW
c+z+/hffZoJVx81jic1VBb7HDj1fVfjX0LaVAZUgiPLPDwWXC6ebS1vkklKq/05P
Z5+55kzNErgAFzcELjVr4zvXhfMem7Wve3MjSTOPuIMGrnN3VlL8gE228S1hc1EJ
yufkOP4miD+PdOmndikyV712UyRjzerxexDYGyZqGx2INAeENdAalXhlVSuZWq3b
qjKtnc+QMj3lisWz5QxFq6n6liA8dGuHDj4nK/2qGrz7fg0Lw98fabmTyfHy0EYO
Rh+oMPpLRywftWn1glVjuVSVB4gOWMVSEhLSy9vW91VNltE2ps4vi6qN52m9MkLL
cW13GvQBetm0qzX03Tv0FQ1Hp1TyuGv1TsGqfrlPWl6kwCKhy7LXPmjc+oPg4k91
BxrseZ4IFUHwbGXLIM3LW6qwpetWlLd/i8wFcsSAI1t34jq3mn9MUJH0/Ik2Hlbz
aV1sUPCX+gT4m2OjXMyGS/ahpML/IKcu4YAYFcVCPQEkI+n/qjQv3V3i+W00OR+5
we99JzPVsOZ1qOaPJUXMyZ9RuAugoF7IuVk28NhRsWxJ1t0l0R4dEtiHgcplHuw6
YjnTAeHZyfRTPK+uLp5fhs39TnEvnxCWv4gla+jVGqu5sTZTItMcL2x5PjyClDLR
XZ5a/IoBswLcAM3gtO8fBTk2ql9ZrrR4nNs5HMGnICCMdFYPtEhT8ylkTvlX8QKM
zTWjSTujVVC2fMNJ/IRRqtdapwe4YCidwnq0Qbk0d1JntHhpQ0x5EN3fmruqw4Dl
p9ieAIo2U8Pdotd7mUAkxafcGd/+LSSdNNwj7A8Fiif2FO/EpWkpNTu6yzqb30Kx
1SYD7NHs1EOiF2BjYJzZe8rAHSqRPIBPo2+YLB7jiRPz8ApG7j5VO1WANDovsW9B
e7AuXzfQh146vhI5yuG1AjanfWh8IBkubCbmc1/p21pfcu0Ro5RDnKyv9lZwq9sQ
GVql/Cd/uXKX9rxL0S7Ow1tHQXBQYDsFwtaMcGD5ZyNLRTdfMhhJSOwT8Ut56Upu
rdEi1Fc5o/zYM/FZ0FirZK+pKhHUyrg0lbWFLVBDzEvyoQ98sl+yMN54cjkJhI8y
ChuZyaVkxKh3K6Lh3tRpa+OirDe5BCawzcP4D/0dEH9PuGasHVoziZtHvhJGe5W4
H6ThT/7boOHUVPXE+xlpLHblobwTCN6+5lQNXi3CofATEq+6htoNIlUomHpWr1Qq
vrMRXu/y0t659MoI8IX/Smk7BFlN2l9DrpzFMHwqztkZ6t+LHnBGQch6FCwsl9u1
t7cGJXVq2UP7Bd8dUCa8bGEhj1489viZjrC9DXGMw/PkV+sAKxavTlH2agJMP31y
nPynwaP6HuXZBkOaJmOHe8gRbLW72IGDYbFsMspb3uh2xOawNgchauwSoThrznie
FmbpTEXUh30HxDI55MrSVgYGXrHo5rfQj+m+WJt6mumILsD5jNscsDyRFlCCkNkp
Q5rkYC8O2WLT2+m5QgqHGbTAIf2b5Zardy9e6Aczan9+TOdIFPql9HJG7GsBBO76
CQCD+VNoX15YxcO4hgljbFfAIO6vuX7u7XP5ckqKvx+Zb0KzTu38u4ML75lCk284
KnUFV8ER+bsferlef1+l9iNU/24dsufRvANwkjKun3kVyZqlewKepdkP4y2Nx0zV
T1yU8IOFrQ/Nl226muaxs0ENSoMqHOUYMGGf+mtJ6m4/SeIuZZRZRctZPJuCYLze
XxA0/7dK54VB0PvmlsKA0sI0iXc25HWSHuqxgTiW9DCoB/HFWaPufdm+kNBYL/3q
o3ovlAsDJMTfA1Zq646Qo9/gFlZU6pgnaIvGbhTfWGodAWlVZJ4TadipXN8eQu1e
5xWO94IEtOYsHDA6e7qtj6A71Wt3jjDIXlRG7dVBu1U3yszDE3ewLv6oHe3Y076X
lbPKOrBhIOcbnhtlcqDXw8jl8mCT+4NZKgfiphAxf56fr7BGZ8VGGqIPxoyC0hMw
wH8+RgM/nDxbhOGUjlIwUAXAprmp+e3tLTJ2Iqv+LpNHK78CuMccWTaB6jCrOQbS
YiWkIjLdXWkEx87bw9mxtf1HyR8kZR0iUsx9v7Z98+rZf+jYE9EatWrdcPUyUM+S
ry0sdQ7EPQ0gXVjpSQqARzFUUIhV4zLjcf4zIkuZy9WnZ4IsqeP5cwGi4sl2JjBb
ic0gYNcOhrtWx5MMoN9yCbMg4iT4rAiSGCOE1Os6mc3jU1XSSrnmpGe2TjvzNZ8m
nZg2//9oH+Ht0PiSKVpBYkh2/d3Mj8IOgPbSc7lAyTd9Ko2QsSnlgWvAENYBNVyT
+7CFtawlnfgnMQ67Ys6G/2is/08Ld1MuKHulXi3P4WggSBuE1psK2u4LPPA+W9yu
KuCjyNtOgFGopHo7P6GddY5jHTjhe6xWiJW9NixkaPgMClr53STEYHcLOtliY3BG
quhtsDmzjexXZSlGDthD46n3Ca4iEdipFVUEz+/N6yA9/cUU2mglHNy+IwLL+p0a
LDl+udjOq3BscXMOnU+7xhah+MYFlgkyyrItRD2rlk2mw6cidrG98rZ5dX4GtLGP
FXxrsa0EAAA5zL5r146tns1T2mCgOMK4icqAnKp0XAtxCIJRMezqaWXsG7k2ScUH
vlvB7LmCyKblW8SOzR392nOBNBxw6e65BubLCgegTJAfnl+Zr1KM7nLLtejMwOXc
Rj/2o/kMAMZKcNHtaXfptbEDzRprNGLPGOgF/taDlAdov2xS5Mc1DePtSwAUvWI3
h0l2byxeS8xDmlafEbkNzHuF3dg3Ed3xL1yKlO8nUikQf8hG6sOVFno15yRVEOTZ
djGAD/CtdxATnIllGqL6IMUJmKgNIyagNwKR7im76jE4dxlVHhXUnv4sdH5m9VVY
Qu8atN4B+jvDsaQxB3Rl66e6qOA7SNPVwHigcGVyMNFG6NUr6ZVGRlouXL8pYaMy
KlzT29ucFbS6GgGUNxCH3Atc9RrtuAGMpKdlgeIqsay6Kbn7gkQU9pQxStfAj9TO
HIN2DRYBBEQxbF1m9kdY6LstrKM1SIlTvYUy2gU5eLVSQVCcYlMVIFU6gcY//21t
gyL0Twe3u/fs/Qw47jCks0iWIDobtpszAy7/ENdtQB3C27j3DfFa3YYYvKCd/yhs
i2BvXP63ztit8eb91dD576PXGOvyIpBnrdD5XGFMtz8jQNZ5oe7jWTDjrC/DzFOx
7P42AvLMxupymwCQ4uM6nJPHj/Z7FTXMYWDuew2s9zUbjEPgk39+nB9IUNEQjjN5
rzcMlaDSSFMr5S7/orCfekhFTGPBFabcrZPbT1NhKP7bDaJ9BEIWStZyunGaWG3a
yxZbrbNGEniO79720w0lljeQv+c7R0CseVmeDrCvW/Mkz022FajVqsuDEhYzrvWR
S6OM28VkAZmGV2FHjvtr8wdj680S17MKzjgTdtq/HYImOabETrJYxpxWDfzLsI5P
miwSdwxg/4IYxK+gEoSK0bUtBqG5URXxK4fzbhWljkuFWMVYACt+X+WvIjTAtd5c
E8DB26xdvMTHa3dZ59Xtc1HMStsyd/LA0jn+3hwCUFP2RbiaTWojT54YvWoJaFsG
FQudjmGbJTcPXH/a5IyjBAIasf4m6GBRnNwfAjWXwSmhIiqMzGi0OTp0gfH9+CWm
J6FuWYYaEB2NVs7mgTeh+jfnuc6RpkxrggL9xyyf1ANKyFdSB0kvedogciOaLSko
KvIL1cZoW+4DT/s2ZL/K/E/T3fMyAvA4r5EuplRI7xUGwEkxmxTjyEF4wUYAyIBg
3bCVAPTrAKhLIHcylK4Kt24wGFSK4YNj4+suG8nlnBukB4Nq2Uq96CyJjRBVAds1
0D+9xChrDgEUav019scA0kuAOA5SkIvQeewo8858/UrUjJZJl5c8hfwS44CfYKL3
EaEvzzv2zjs4sf/jaTAkhgkvUbNlX6e/blLcFNxfNACgsTqBLYTZN+CRiidc5Bg5
w3lQu7poOudy6uxHQTqlRdQLP9lm6C6bHvQfk+iFhoOmU5nZtC4PyGP5hCEf8qP6
ZMVVjtVWLm4uyTZ4e/97Zht/+fxYtQv075p4DUarPyyrmg0x/pFzNLLUp4TJVOhS
go5cDkMRB8ntgaPf7nlMn3yynXDM1Md1nPDT4lVheCygaFBQCNr60IANreY0a+f4
Pdyisf95ebYnbfeJ17LQiiRFI7rToYp5CG4otUN151FlZu1z5E17FAPoOiKgYtSL
nh+GaCpFbM5N1yDMXDDKQ6v+xRy2bhAOKc1lETHBCEeIIb/mKIZDcPIhNw6ZMbhC
rAjT71q5zRQCdAnoVbENPp6//z8v/FH6CRIui+nXUOoU0NxNWSLPH5XKYCZA/F2u
PviA28rlNC6BanzFTDzw7aKDOaOR/RXvyK1Lv9apMJGFPESE8V6NbB/uievssJ0O
iY9bFa8w6bkseXXTYF1mpQpBH6+oXga30yg8OFEe1yk+VNA88IzqVtuc7fxHWh0/
Mss/E5wXc7qSl6OKzKPh6iDPEFxe1jccraVYwPZdtTnTDKexJ1mu4kH23iqjuFSW
lZydW/y+jEjZ4bUe8rSbGyLx5+wzup5qhnjkPGCy/9f6XN0kr1Bx8iRmjTVwbJye
8i8qvIVshDpzU7wh1FVZdISLnRhU3mT4ufoykzMBHTWoo463QTdbd538whPewA07
VXODJYAiVlhH8mVLbw34JzKMzskA2dein0mV8BEUHjlExAoliS1R06nbtCQlF/qb
5Z/nWXX1Eu+91XWXVRuIsuKhicOO7AH3aJ4+RvLnUbeFXA1gB3OIGPGIK6UGmSC9
3CC0M6NddA/QbkDFMvKUCvRfDmHv3Ql/HkqOaYQPH9A45uzVhv1j1edl+tzQGrAI
BpiD1Gmzk8SfY7lKgXs9TkVo8jk4C8p3wZFUqaI8EzfBiqBxNYCbwmU4zsue7VXL
fAG36Bki2nUTlDPfp9M3G8NBASDYfyQ9IJW2/02HmiivM9IahZ30ebfNIc93aHzB
4asadtAxW/0Jzq8S/ffVIcVeSh8h6zsaWYWPzQM3jKMNJxu8xSTCpAfIH4XS/wyM
BBH2j27dt1Iw6oUMhid7FlqlHcIwNzTK2CxXKpjkCe2a413zMXIyl0SG8C5q8Rkz
XCjzTO3UwrlJtRjCIY1dES67qF2F26izs1NqlisiGDYBpsuHxnZBBFB8TBjfYuPX
rNrKQy88h1UyNzdZr2ZP79mMV37bum4tZ1va43I0E55Xytlaxyd+mEcB+G6wca/0
LCTiyPhlxveFyghysKVkRqSH2HzaH6uwTtM/oFw9m58JGXyDV3VDGFbS61PMoFkP
y+9hM02aq6o0TVfsET/kofIq+v6N5BOO5yD2bBVdLNMNGKkwPsRpLmgduoqDZTl8
LjpuljBwLHaKGngST+PI/728Dd/OU7C87GaCjN9J+L8=
`pragma protect end_protected
