// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
+qfY0cuCP3Xr1Tete3jo+QPXTZldxJOt+6Y3QkbwRvJYVWisAIUQTXtM3qAw4U3x
GouZEpa3nGPdqMZDBH0Rlil+yyJ0QUJm1t5xU+MdRW1Uvy7IfOmWRfICwg4ICZXi
q+3BgK8ixZI5bN0cnNnfsakX03gN5bFTeLi+P+DaiMS2CJagM5J8kQ==
//pragma protect end_key_block
//pragma protect digest_block
W9iHV8lzm3IpUPYVITHuDc/vs6o=
//pragma protect end_digest_block
//pragma protect data_block
PjahsW7mfqZ3E08FgMU4rI84z1oNIOxRb0M/LSZJ3ffHTkLSPMkI6WiQTkUl5tz+
/Vix99BKX9uKXoiLWc9/NaZeXAvyBubDcGxezj7RzGWCJj5onT9NS0hwj/UMpxVo
9n3JNEDsMqy6HYgG3AvAs1ScCvS52CiByc9Y4oE0VZeTJhXSkCm0wWV9WGJPBOZc
yTVTKs1xq+Y4iGR9MJeDIL3Xhn6iZWVwjbhrg/q0AKYPsN8GDN2bnxM5y7jTr2sh
LUX1nQC9LDu2pDp5finUDj/d19lQvlQ4UYeBYBr8YZGsbDvJPPw5I4uoxpRS1JMo
SOrvMi4kl2J+geDXIKfCieitrZx81eSFzBk/r56KJ+Q7EXp+9YSVtqWeherS+GoY
DSSDecr26yrwOhIBhc2Q6PG0sfS/ENdZSFg/ycIU20TuPdQb7rUavZ2DINWWcwn+
hk+/GEnZyayUBirdLDYlMudBSwfqBisrTyRxgxDC0Mr9fOFXMHmQS2a3jFf2vts7
Nng327mh1Qh7ADEMwSqHcIxwoIdyVo82l9bjeD1fMO12o+nHcyKLhMGzK/x7RvmZ
6G9eD++aw1dhz2EA5e8lA+QzisahLwzyrIkQPu4+eUW6GNUTfJZipL7cK374XUld
6kmohBSFJfPg4UaX7ZPmKEe3h+DJHnO9YARxDl8rwO+dT2vG6c476l7TPx5iyaXQ
jfuH8rarnUWG29+KPGix5ha+3Oe/WsOUIU6Ct7ylY/NbD4wCSf9dLC+Fke6gzctf
niIlTH5f9gHqlzmOOKbzijtjtjbaMe5b01ogXhHtt7D5XKeA8yhMx7V/+YmCUBVc
RS081mMlTJmGJ/E4u4jJJSaKRC2t0D2kO8iv9AQ7il/K4O7GP48uBtZCzWibmSEH
0RsTBe1AflM6SMxxRfETtkopZJR2mkJnBukEQfZdbUKOjp5xB/lS0o6MmSSS+gMn
ReDQYmMN51XVDLDYOksUO8AJJ2ph/eqMKyTB4s2ne3VLPL2EVL93ksSWlQn+/PXM
Ka8DEN6Ycuzj9AOMhPV+3YLcOHQdogh+nTu0iHP8le9UekFuEIMM61snt6rjVydg
4qdXbAtwD+8i1FqBgRKvLWXrEsiGoANUGHvxyl968cl7wYCDXLa7L1EqtRCgiG7/
RRzV2Oq8kcta5AohoYoc5tO7pL2P0wvjuJqLSGRhNTTgOzXt8bAmAAKDsenG0tkl
DaTL1MFw5gQkT1UxeWrwdbxS02YbdflGHimq80GSfaizcFKZuZ4t6ysmlwCCTdn5
0i+HWrZyL7Byx0Sxz9i0k1D9ExqnWkQC3brdcM9TLRMjSQ1Aq0A+5gztxsA0G5z/
SGQd2CLUx8KCE+Woy1JvYx7NMcVnp44D8sf7fzrpq4dvEJ06l0GkCkIrEPsySn7H
EyADPsvSva/O+PP2rYM7Sj6ObZhNRtW7Cbvk1bQYnbNfxtfM2Q8+KH84oe8g6ctn
d2ezRyWr9pqztIyGuFp8x4gHHt2nCp8Lf7g9VfoCSS7dmOnR4ZKgtGhgMzdMr3Pj
IicHN7Zco8ReZcg0izSz5pgNZQU8hIihTURhCU+6/AvsXnQKzrfS1XKMscDrQGQy
KC2IlX3EFFWiUdbr2SRHwM0qihG5vV3Amcqw3TuoJVxseBmsD/1WDGtzNdo6ea8w
caTZ475VDKury2fiUnjoTfyEDbqQ1j1Ml5/mNH32YSEMxadOqc8jVxbyvmQK4ZFn
TSEaUpBQo283Uy//iuCG+9pCYNioy8uP5qVp9UiZlwn/ZElyEf8Ox15y2ZH1J4zP
g03s2Nv973mZhG4kpGtQKHIwc3ewUQfOb/iopqn3wXDwC3uvzHLLsk1ZHfG0aTW9
82MMmqIE5LwaVXXY7QZunGDrjqgDLEHLarKaXVeVb1/ozFPkPx72tpzmmUp8EuQ+
QFRl1t10LdvsAlS++tStmMetYnpc428rFqUlvsSxcHYfaeI8Us/lbQa+/xbH4ATl
Du7sUwDaIDB2TrGNIA5sRyrvc5kbgnvV6zaCFW8db7nJzON+IZ8zLxhL1WbwklBB
LbZyWE3MDQjSVKoMrQo59RHQSHBwiAK38Ue5knfJtWnljC+E5OpwfMKXBqYMKYGd
jJXiYSE2OIY+qYg6LM3WQrCi4aPfswUrt6LaR3XgtXIgUyEexKUljQN8sS440DNA
N3Nh87U8M/Q1F8jf49qF/9G1OFgUxelHtiuHMsPhl6FWiMQi1InXGb0XdH7ghnK2
KHuwXIFFsizP+/Ae0JV0hIIODuKWXVfSKkTLvRfDk4rYRlHUkOEYi7IdDPn75+3m
jBZvCOwH/IkB9dXjrZBgBbX0xWrs66HHoeL+39TAQwqm66GfbzbxgF4x4gDTOn6/
jxk38jmSBODj0HxDW2S76T6bobrpYtFUla3lMqOVp1fpPH2sJBSXDYRpFwI3Thzc
CAsmVeMILDXMndqOEMhPHgAayWpvpnelxtiE/gG2ZAyPeDl7PdH2sCYNlyK8EMDv
leHVevbe6rAlsNKuRVC+wxtRpyIO/rY/zZEO2PG9QCCvyhkSAkb6Fp0by13qdSHq
FCuNJLizYPyCdu8TSEVXMVffKkTrwJEhfJJLTH8AHKryiy182DYO1ATg/AIR/Ft5
gkiUWmbRRTGLunibP4DHNXHSkrNqD470wsdphMn1DtjxyTLMTGZukef5Q7w2dsmJ
jV3Msaf2HitD8z9T/RkVXuYSXZmBxjEseQtXpI6ogDI0y4uB+xDcRXx5sl3iMqkK
ERI6hHEljXu+4YCkBN/rBCxMb6d1IhsX+BwwsPs9awJbpYOFxkce7FvJIi0ulEPM
/wfdJivp3+Fm0jqnvFDTu1kp6qIiUAABS29Z9Dogv5wtxUgthm/whRYHtoTN3vd8
2vWWfii+2MMFsYgMdihEm56JdnuBYHNiHxStmfSM2zkIPhhE/Bjbiw0ruywv8nrM
SX9JaaB5IKxiQcsQbb1Re2OEo310+QiAHtJLMroe0WXPDcMEnzX0xTp1/qTJGA5A
BHd5Zhwjl1X66yF1+5/wT706d2qwoclLeJwR9KhnZBGV8gMAAkXBwB1iWqbk8qEo
aMbROcH5YZKGSfNL9YaK/LBQOQf2fUN8nCiIbopCeMvs7jwi1YTIEG+fMSuC1Y7e
ut24j9BSHbJD68IRkJ1aUDSPqnY2cQ+f95Wp0xC2Aobo3Lq/u+Bn7sHXp76oG3va
WtgooZXW/5MXN74A9XtwaZO0Uz7Ws2pL7Boqypa+lMJZPlWioZ7gdPNODhUNqekN
Zb7i4VAOMPd3MiPZEqfIrMtCPT3eEgMI/SrJQGgfcObqW9P5fuZDxC8IczML5ADb
3B/vKoM5WJM3wzqUK/HpofSaY1uvEx9fUeymxMzes6zqXxJ11Wcoy7ZOwiFVGztq
JG8op0I41Oi3zKmtDKgkVd5+9QRF5lRkVWcTTGXoYv7CGszcKnp4DlsSIf4eBfFO
lwkaSnSRXKtm+CMDJd/q1xMvY/8oQcuJ24BjWAO0/znSR4IdNOzIfHak4HXBknz8
oQd+m1S3JxXj4oO0jbsi4PUGrlawXKZghyijY745ijfxfFgMw/nawc2RdHbd7B5v
51mTGVJCFxabL5shsBbxfirMByCg4lMh9vzbhZ9eXl7+txaf6CUicucYgMwoGIsH
UPFNTQDotXm2a5caeUkbwARUM6HP0rcIL8cmWgBxmxi6aqj8/UHVwa7hvArpZ//1
fogc/dXRYPVTznntmdyi/eLjwRUaEXxQbGiu8+gcmX34JqEEVp5guNarfdYH4mQS
nDmCd92kh8MoYF2qoiXjyToaY1Kzd2yQBWrIaezlvDsNTpuVurExFqTliCYbhH5P
PyeqJAlDCueTlCQlQC1UPynUOS9R2dUQLXcXKqPt8h/xGeY/yfAyrtPPhObhJhtJ
r00G9ilgzoiQ36wRxlot/zImKDzyz9TSnNqT/xgqX7b6IQslz0NjGhfuCHdhL/5W
eiNhGp3UHEL17XJpzTN8k+7lO7BsutYU3OPkflihKr+VaresMF3LCB2T4/JSmHdM
B0wCIGrhe9LyV4gNeQJtHIahxK9SgdM1Qgjq6SSqp/cMOAP122fA/MfwY8wfaCiU
dhlq9Oih+pWrj8aaGizY2QdtpvCRtIO76XEIhO6Po9X04KysKfW2VKi0QwEUDNCQ
5MU7pb9cW8baeV6g5N/NZt/NsRcDU7Y2g5dOFxNlrgbFl7R7cMf5hM9RNIIMtDYp
4n/zo5fb2MaHOb297RRkjxVIsgFDHFbRG/4KRk1bRJM2LwQBgb/b5PUlhtJEz7Ee
uFGobzVNSd/KPgKPVADmgfEs5qYEt3GX29R7a2uw11MbmFfingkZ897DAl7uDyQn
kTfIwWCV+V4s6JTByVm04wjoNfVh6drRk8LFY8dWW/iz6i7B9eW9AHtVpYXtrlXc
q8jsRozGMrDZ+3Y5NbUJVnEZyyDKhsoB6A+kZx4iaAPL8P7/n4Ncw1gEDcDKtsG/
qymsnX2DV38W5T8kevigzMWI1uMAtGLRoLlzhVm9rLBV0u+49fsYjtlHN48wEm1L
bv0MXYLCNnn6Xz+4MXgSHCFFOPPu+DNYUHYyULJoDqLTsT46mt6ZsuK3V0WVXvnf
135+8wCgcmxNmgmGiTq6XHthlb1x0FGTprf+1OAy4tJlFvmNACzFQrOOPTTYGKID
ofAbvIcoMb6ybUhD0MP+/PkSE0rOuOMm7qO00pjnY5joFdrXLqsQh+UO11vOAJt9
UDQgITDZFvTWd49h3SIizy5CCSlhKtQQG5NHiMUxs4fKAdKP/d3sfQac+NuXpXbJ
NbK0ylru45QNgMFQIqm1DtNczlTH+wFvH+PdcfVjPNZd4toGNTzNHPBu6zkhFhEi
pfobgdacAUsWV2mPq0WLPbM1VXHt2E5DRPjY5XguA05GJvk1DaO2En+6Wq9rZoci
8+J2kwkUgreN9pFIUNThlo+lCXxj+N5OKJQq3Hu2QgM9eu1QNHfqCb+gwFIJQjqx
UjfGxrxTz3GwQiPxESvIIPXn49hLHoWeJRE0eW3GeAWArAXmi7phrjkZ+9drPTtY
2y7u/Sk1MlOFwM4e92ivpqTD967P6EBHUcIEgsSzeSCLHuIfAc/rXFIfHtrBBqh0
dQg04iImLYT6DORezSOi4Oz23uqGkPcfG5zOZWLcGn0rxF5We17VSDreaLB+rhOy
edsZpMzLeRrfB35ou9K48ybbDLxvPBlm+SNpB6QUp8Mkzyt0nNDRYH8gvgnkHfs2
0zfyBeBLwtLB7ewU2NYvnOGfUfNImBAuB2EinQ2HgG1W/mbkRPn5f1Atot95FVc1
ZP1gjV3sXsmS7tgoYvR1AJS/ikMOs40mWWXp1R4HnU6wqeifAe1KGrxi/QHI0Wy6
Jp3VilZhZzEwMI7sjUw4JV95X0BtTVHhdKDtq6B9i35UKRJTS51jxQsDWJprj6oz
pyCPyloE/Z6b/1a/RS7Sbgq6LjTSaT7vYLDJmTaNWc2oxAqYKEatfQs7wbB2GkJw
IU7G+hovOd+M9efnDcNqgbj3Po/JlLmJvr36SzVppUWeaxzLDJ8zaDysFelxk2XM
xYR+nUO4hKnqSpKB2H2XeXWe5+gX/t1HsxsebLZILScA1cTi5NTobNPLCavVn4iq
D4Y8vLmJAOo6HX4KA7/chJkqUp+vFMaMFX3GTTxiRWme2FxUofD7/Vrd0mEPQ1Oa
zxc8WLSd9L4I+KLXaE81breFP24B9UnKgntaA1uU0NS40B/d8KWW3/dQUARCyrWA
XUezmJGbfGEWdfFKgR/DzJkPR9G23GhsWNfvSrrDLLM5QLNmDL7Set1lAB74gRgx
kBR2Bn5hcHsQQIHf7gSgc0fr8bCuCbFleDcxbdcp3EidejRsinpCwHoD8FC8IjIY
zAh2q/MglmVQnpWj08cj349wSKXN8IamjmReIGgKoDE6uURXjRPBPUJkVfwOolHi
lpnhvIKKNH1M0d/QUvfCF+Zn/npN4C0gb3SWPf9EE9x+QIITuF9xw/NNvtIQOc0R
Q46K0stQCA0wrrBBCpoSXsOUE9q41TCPmRNvt0crmPHR16it4+J2Trwf0OR3tewh
KCCCvAmrCR2U6bd1FnK08bj3Py5r6+eFYYO5KC+j1NAzeQZg7h7ayLCyfCNzBydY
iCoCzo0x/8i1blOcUymHs1S/6i3UUPNr5lxauNGan9hwBTrc7tmsZO5eyZA3iWiC
b7njC7OPDEVgOI5+KmHHBcFJNim6+5CNzqNF+H0driuifpONWUYdqGILzfTdSEdH
omJXrCBAGyu8ALLXXb9nuJD7X7dhM1mTBSmT/Bzg+AEaMqBDY+3uAzfDC9AS13/P
r0jhPOt41XZxLpIF1qz+i7Cls/y8MAXPTwgsFjNxPRX9RD8Uvzckij8TNuytlNuP
TaHCPo6tgpdw5Lxt0Ts6ehzPD554741FSGpew33aXyIUiA0b4RRfd/2ooTCZkgmP
v4uUHgcquGWIPt6PCNk+KkrA4yaEJxp0F6hv7gghaDNL8WfFpG38+aPuLHrw42qf
p2SX+DVAv4cRzURYqFQmu7g6fFq30f4glOTP9mzhSArPKIcPbsfN5hMNJSnaXM5w
Uxr1snI2fG3tE3x6Q33jJDVyiwCEK8O6qHUq/sRGphUwbTymHbFJ88ZYwM9U8N3W
uQxioTFsF/jOjp31AfoMpzyk9D69oxlgjZvaJle8p0VIftG+cZ0B38lWR5lSD2G0
usOix9hPmaCpF+oT7LmjmUJzs7JMnVrJh80acX44BPYbo4Me1Mi8rRnrmcSrgdQ/
6qEqrwm8utGU/ukVVQgySk4wu23zdRb4HWrEPtxhQUUvGABjZxhOA/7xOSpJhKKc
4IT6ntPKGNkUb89pCIa86Fn1H0py0uV/89r2H+/pJp2kR4waEkRbnmKPUMCFZL1G
gzVNI1FysEbNdaexeGdkWqM9upAHz0W+Q45iU+yt743/hy3HG7gZjh5d9dlkolhd
L2Ov/FPr+RtgiZbkphHkA9Ti7Y96uWPODt705zotJFRa3f7VUlB8Q8JDNYyRTpWY
JSgFiKHrRMtRHqCnTQ5nMIrQpEibiIktFwsiqSEc0/u6R5HFw2+x89t6EiUcNZ1W
KLQarBbiGNO1IKIDuLXvseHlvoQG4yL1svvjsVfvrgKGAdHwGZv8pJ7REcQuD3lI
zbnKT54/nMJ9QhOVK4DLgwOBd3apkBP9mQiEPZ7+XPrNVsDWNX1qCu4Tvaea8y4k
G89AqnyGa71BIgnw/Y3IsyhCvbLfxPAvhzl5J6LkCTnC25v/Ax6SMD569SJms9qp
wqjaxtUWQWkQopRYwvseYRW03mgztb+WzZ0gc+gznIItHJ+AJIjavGwhP2+TYL4S
XeyHcuTr7QKWt8mlBkmWHHyyJZZsYQJbnjJd15+OVw5fxThB35RT60uuNsWaB8l5
nOCGwOF5dA+viL00yCS4dlm2RY/+Ix1c8BRzzA7ELjyCn520wQU0CscI0yTO8uuj
2ZTxX0v/hlc0TpErMwACJUlrGgkRfYYfqMFuANrLuFZr7iJGQy9fZcpitLExlROh
TGpER8iVWPSpWMp2eeqpkSc3A4YKNPoGD4mUwisAllsTfBZymOkFDHZiKsfWxiJE
M4J3e/2HKI74+/a6B2PP4gKxEXQzg89p4sXAX3oEP9X+4sNFqlAeV0odyxWmJOxx
1wsk4DbgyZr3IErRgUCgn6bDdfpPkuEuND7xqGljou7/A5m8LNZULGGwA1a1kwxB
l8JYd+OpAu5IoB4M0tLMrfd37V8nxALktcJ52XoMtHI8o886oZNjQFJWP9BpQrrR
q29Kh3MVUG+v7oiRaKfDdfJRfnC+AdhaMZvGhdh0Xx6k5j55S0vkk50ykYLQV90w
aW+7ja9//t+Nmzgfkb7cgNwJpArfVuhe9fXTTv1svk3yJmOMOlpzwWb8SdhRVySu
rpw5TsCrmtj8XwpE4whFeGS1sts5KEUbrdlRNJeirXplbmIYzUqbbPUOx482wueW
0QM8e++ab2FGud6wFqEaMLqz/nzgaR8GiAwBOpHw8ROoZXZK0QNE7G2VsVJZYGZW
SXM7MU0Bxs3r0WCRkhv8bmaXFntdGPoh079JxJqIDiwmQrdJGzOCgvO9oc8ihJ5b
hvjNlgl57mi17FC094/b5f0Gi1mS2R+okPEqUFNbSF57DJtfOLebOM0ZuE5H3/mo
eAXIos/AgNq50lolEWKoSHcwwOKFmV2kV0qZhs9XCIMqaJNlVjFZCuE2odyPhCPo
cjU6NWlvubZN1d4DepaxwIG83ROD3b6LFDoIhjidFcAqzuDT6IpTh/yW44bB0VuA
FMyg+3jLzR83wLk5kwZnD04zYTt7G20xbx1vORKcQPybq5VrhNBLnoAknFzSwHNy
0ExXPFiqBI9mArP1PeCHVMG35H6uSosQgAjvbM3F7c/tzKRnTeWO8bTyw46Ll+Vr
BsblUNMJXMDHuMNN9r7UHczwjGXjcInCFUYaKMXFRQ3GYmxLeW4XkCfrn/WJuswi
Zcfjb3HepHnG3ECrqdsYovSydxrDd7E4amuBEJh2aoX/wIFtY6aMpCjUt5QzYbXe
Vws6a7pkzh8igv91vnijgNt1AkPQfMykB5dZqg5FHvSsEfWpVKJJdSJ+RhEYAssq
SPTA7E8aZFaGCUap3L3z2GJTkvPglBSrBmtRHFz78V+TGiu/d0M4/aNx72RHKhsU
HdpaI6W4MXXCQmgRzIlyMHHTCQL6JEhT548s6JpyE8JAW5tIxNTeZO7iYQDYICF6
9iNzJtDZMTxwTNVQyjDda6kF66IU/Yn8bsGCIVwFTKgdUm5NUc398WGEeg3ElXiv
PPkIs9HrzoPHq5h3lF3lErXx7UV+2TOt7g4doWi1t2Q5F62EMQ2j5IrjGX2mOOVq
b6OQTEBjlStZ5/Av+BKr4UKiDndcKddDG9nUQP1TEQzurCxLpghxZkEmmBE7YL5f
JuLsELEhrhjBAzEtWFBc0dU9j0nrH5MtqP4CF+m3+LacOdLdegbIhT5tb2afewpF
WYGILdvK8gDog4s4t3gNJKD4/WWF6PpmFSEsnVO4JYAIN7aIYcBGEZLr5U6bArCH
+GD2YLbSrBdlMzzNC0sefzoMDMD/WPmllV0F+eVWMecM3VJXKrvnTyHK9gZYExt3
9xzio7sxHxTtEQzenQRQ83P1eA/iKzW/878Ba4aYmHVvPS5vGdJt6gofYJjkvpo4
VqUumKBgXnhL/4MILURePWX7rhNBE2jfDqLC5mMwxxgfdY4x+5WgoyvdP7fsI5Sg
0GW2BQTr722EokvaumKxE6fX3iSY4KxYdRokp7UptVIuH9i4nzl520f1Q4LtPYXT
PhddH8x6VU0esFCUI1fRkLxdVszNqJQdL8hLt4OrvtbB+CjutQC0yNYIGqLcdPJS
m8xY6aoJJjJ+ZD2+gZt15eSjAMo7bOWGf6Wp/bj8cXDP5of6yzH5BrSekMA73vkU
ijUdfr6VAz3aILK7bzz93Yz76rqryQrxLV3a0lt+J9iBrAW0X785lQJtZBEMrl4V
I24FaZj+FYBCknrxwICWhWquccOgRyt4caP42VAMZgDN29TYtnzrk2+Hlskrir7f
lknzZfui1NyzpRI1E4i/SuTCHvOFACupuJ1nydNNp+eurXWlkickr47rt6cZNsK7
8GqT7jSdZCa0woC1UR+DT5V8klrJN0srrJBax1mYws7XW6BE3mrk+aNfTSB6OFut
ZOr9arrVNLn/cdi6Pn+4D6OQ+nzNxMYaazR3REmx0a2dSFqwPYZ4UScfnFGsxXo9
LbM0wkCasyPcgFhbFuw/XynX5hYgiCpC/3cO7fwiOZ9kiXu5Xzl/vaA4JGvu7sup
8esBYaQmyZclrUdVGEdI1R5aw06hVaf/1AYM5PPyd+h4iWZWmsjLQCl+IfP+dCA+
hbPKiUxC7w5zPzapdQ7GAn0oqov0n4Xyh2EGByViY2rZXR4hVcBK26ahRoBog45H
bxD6zmArUx8uaNc3XXeCYrbsoJ//usq4sIWqdQqDMQ3O/gRS/iVsmtc4dMeKMRmq
CWYoQK5pSg+32vJeu+YQookuS8JSnL9cy2c/78lFV48Ayjuef2nalRZpU+xZG1P9
QzN73WrF8oNic/HwLKPX9pVumJ1JLI9c3MBjtiN8IxqPOD2+n2sikzuOTNng0CuW
+FkxHMazsCZwmdPwBPVoVffm8tF5aHfUsmSGs4Z5J/OaTF6T1tjSTTqd8kI0dK0Q
8UqbetX+ZRKxjV2Be9jebNiN5H8gTF4FfkN/f7Z/cDTzUY6DBwsFoLr4p/AQRDUo
Ed2boGEjJ8Aw6ZZXnv22B9fI6gUqCdQ768sH6+Jcdzujx3VXaxnxmSvK4y/d5kRi
Wn3yu43GaVwNpSsDX+CDApz55wfp8cOv/bXY+R8tFNLctbP6rr3A/0ESiHPW+W7A
LH4q4KNb6yjj55G/rDOah44UeDbfJvuh2o7wo0kfsNCpmjGmlrSOqHuoKbSSC3Z3
jeN1+qSHCT7DKcsCLfqhk25Vn+RJXsteCNC5GqlYSXwCmOSN1LBTmHigW5SGpNbM
9ud7qtvPpIwZabD/HqG83d+3jPE8ZMcdlhGrxcZFg6xeux8L+RBmAmXcxA+YxnS+
xcRXAPG4fWqUsDlr8VI/Xpuf0CHrSEny94rijNpDT+dL5Y3J9ywUn7XDBlUpZ1Ms
XehrYHEU9J4mrW66gimwUag4Aj1HJ4uK/jdRY9cuBWyJgfliSg4OSQtND97OFVkB
7qFnTIk9H9aT8BnlnkhpP3d2c+tsc2cXFVKjf5s8YZWC6UpykaeFrvEnTwM2b6ne
hpc5s3esjBKHOEc+m3SSqsal7fz/Idx9Zo8tzMlnT2TAKFcEY2SIFD9T2EvO8uN9
drAgDfpBMIt04F/3DOAEaE+w78LzaCaNqnPkk0/pa/Xeq1Nr8h5bJKao9m7yhD/a
wEuvEEafxmyb/9y2xkRFdENetXCEmRtz/hQEqBj6rAfcIfE+XUFMQPnP0V5okLXH
RXK4Ehn4lenLE9k8RHe/Cdu8lNIX1aVaE1BUhMIS9e75fEpu+bwJPYd7R1QZnw6X
6z4LLk7HyFds8cl4mj634bWPbPQFParBFDcDEPnAq6QstmNN7e03S2UAx59RdPU+
fcHzuFgWuSae2QgIL8upnQSwDkz3kpFx+qu+PHuFwJdq5zzhguKKCj2NcJYanjeG
HQvBsKwaArEuz5Z8NsVqV5xCrKDFf40VXnfn6kTe2Jne66q3+cq25ogaeSpv6C/z
FC5LtA73WpRLpxkNTpZEEwvTRdcDCLcWybxX4dKznpYLsWBoBqQKNHsbTl7R9hDe
iECvVSHyY7IShXHZws4wSo6IXEUZJZEPnHL+kxNjTZQl031zQYDHd8w0JH9uxcVu
aNPSNxDY2GCvxVSBGhG9Lfb7B5yt0Fe4d+Awa3TNSSk6l7GZHHgJVPdvmyQrdij4
M3R/dFotmfCeQU3oPC+A9lfXBBOfe6YAwnTY3U/28zIc3iJV51hDbaQKCSEKm80A
bcuO6MlD9j2khU/bBvkQ1P1esuaVrWopXVqSOKY2qWAEJh8ef4Q4FtJwGgccSq7S
JCe39EO3HqoCOLoJ9JYly4MVPzUeY+6WZ1tJA4Nue6aQUYQzgGrkA1V98B9Z+2Tw
Ni2FTbK3J7KkTNkf8dZ956R9x0IDEkYJTGMwhptIoKa4PIiE3Ajy9pm1l2+zD37S
Ihrp88snAc0Sz06gBuHTDbeLuGj/+UP0RLSc8CM7tCDmjQznvTvWUnZlqS3Wg3oe
W3Dp+jChQEimK5hzh1hFNGmYua254Eurz9a6GS/q2C9cV1H5zWclBHY5MYXlDNq1
Nj6K1qZUtbWXwczCwsEppK4TC74DtkgQZzJyAEi1FQlQxkxaLHRG4RpVBUsyt2pT
NCcULdu8M2AyQgDJbWBJXeHUmwcZMHm85aWhnQa7aa4sYF0UCZKwBxuBApC6kpYk
mAxP/e+bwSg/UZr4pinbpX42T1HEqYGXEuAggWUlcTECBL8sC1Lk4lN7SSq0Ayea
JcG2KotwZEgRulli5SxC7WsWBeNch8ZRpBeTkil+Xp2RIla8NyqQlOiKNgxgYd0Z
xiTgrm2ds9ou6jXdxm+RdPaaoSO3MS0PBQi/0PFnoxfw005HDhnqhu8A2nU6If8T
ve0PT1V9Uxpb6wKSbXKHQB7jf4yMh06QSf+4uI5fgc+TH484/LJ/TkIEzll6sAMt
Q2y3zZeDld5ovzIsfbdDhNvQJ1VhrX5bIkHp1GHH+ZzLeU8+PQp+nASKfkxd47+S
Hf9kOjJa9CUUGcbJVjDxKusZFLapX89EV/KubKYW/tPAPRmFAjno4DMytYT3kftn
Z7tXHon61molSuGAfdCowiozkGQ5K+tqwnTpEEzQMeslq6I4GEU/Oxq7s20KN88L
eCDm7kTYZp0mpMC0RaLnFWr9s4VmKJkYDo+Y5Jw6Co3S/lIEq/xS6u8Vdv8juwIR
Xr1YUjPxbXdOtAWGvpzHVMGlhy2WRADKeiMW9uahpyQIqklqpBTJN0FaVvRz9Pts
3DNgWf+JTp+Dsr3wzXonr6esgVbhodzZc/qBZ8ne81IjWjAoj9YfBRX4+yT2pSBf
UwzsjuZe5qsWxULR4H7fc4TqK/SotrUqDWRgM1KFxJZ4e43zXCXWJ0AePTVM+qst
rDKzoP15omn6uSy9JM8vzyXCPCsJaUPEi+YvaJL0lWVLlAm/mnxkjnFHka8ctrab
7yUy0a7H7c4AdJAqZJPAPganm+e2FH+y0//CieFRyQqqDfDo1K6Bh0demJsASZBN
2SDOSlj6dmJ2J3CqBvkonDevfuCwyey8oHcfg0ShLkdVTGyjKK4PB9Nl+zZGcSJB
2JMGui6yzqyt2+e8A8qRrbf1Sm8Zv7zZd91QnzYlbYBoD61YZc3FkkXI/OmflhmO
vSVhtZ+L1NDstA2k4i5/LMD4YSkkRdZ1MnSJBbhvWK/yOot4h3lYth4CZoexm5LH
CVzudbh9MNw+jXQN0cmhldoA85eJY9J+UhcTXKWfpY+uQJumsAHOeprQDkJXSqoH
mguWg0tD9+tQyrEwvVG8qIXPxANnKZTujOFZl62yvE37VdiMvLZFEPyfkgVBXGDv
67JPvg5CtGNuHFkXy4xQLyliayZpYYzjKGoOHw+s0iHAQ7PF2siqcmwr5klj0IR/
v5reUUql8LmaICYuDbVz5e8bubucHWZtwna0n1L2unJij4mZ2fyiYm8oF9e7W7c1
gQ7QCCalZvsBZIU0tm1XT2Bc4MW/Qxh6XnnbLGmsV7arK+cofLRX6mH0GIhNrfD5
RSYJcbUSC7htxxzl52T/Uy5SluADf5zOeEK1Dt/X+k8mqYyK21YsOAuAAoV/K8dO
JCcwvwodY8MRMzNYYRAU/lmcyforNEQYZLptukADz77ZWnW8OKBnqemNNX5G3VA7
zpQ1ThlvqKRlQuzHzjg2daUu3cTP5FCfd2IjNbzsZc0+Og3g8WgD0v4GwleSOuNm
Ekm48qlSA99Fvp34ZC5SClj9R+VzxIobG0PB/0NG7pPr+KHpRVSZhIBf6agM/Qi1
WA5vDXX2NYI+Dfwk9M2KskH/tdDSpkGLdMYguBF4SvdHycLqC7g2j27u8iWrg8C/
jMy049G8v96fyrpBWcpjlt42najc1rqdCQAsPzNo+dXYJcB4b0qJBWYJugUJ2HjP
wglwkqnwBWozqzzKZFvy2Ldgu/CgvshTvh99Km7ROchyB01f0giBr+OvU2qgc9pI
+MhE5gKlCIJhIp2FHF56xc+2E7Y4rp1ruCS4xvyseAeIJrlwynkmeWL3bisLXrzV
pz0yVcp3/UHhRbogwtb4VY116KhqSmq4gBGCEHbrpIhOpIVryVUvLHOMF/fQ1FJT
VaD6GGsCktSmHzDhiaWmabt2FQXB+ca+RT0uNo+07GOyFMPYtxu4dXdKlkmskroI
jMUqW63pydgfAATeE+Bu8zxEnTJImGiQJrKTQ939B948t+QMeHqDYvoVRicuMozr
YLp5RtYgc0b/m69Wo6OGJ9wjvd15wauDCw8LF/odWrfdLKBQ9g5A5bxNv8gob00a
QT+2xL0Hli9aBfJhBggi7Kocj/cIO1bIEENI20oAf+fEYfMU+pDd2WFYldK+Ewgv
15tlkOxXQDqxr1QnRibKfQkWRI3oQnD4Al8T9uxhY3GiRxEJnrTCNwFwcaI0LEaR
2G4C4VVVed/+QwOUKKvVeSJQtwh3uiKbpNW8ZV/lpueQw6OrzINMfUJqLNKX9vSN
t8v5l9oGosYiNMwE6BqoizJxiRvm9zRkxCMDyINzedQJAmp1MQjgpTdk9lv+9+Wb
EzmSjkvajGGQqFZi22T2Rt8ztESkxUVrU6O8gUCWoM2Yqr6HKlPRW/gEysL1M4PY
z20vna2IkFaDYGibYW6+suF0ewCrtDhEC43EBhUQ7BrlRETP6RD6A4NuhVvhrY95
R4rQWlWq2GiPfRkh+LbUlaY+OWLWkIa43lA6hcAM9gn7X/5MH7EtpQUUV59SM1f2
Dn+cXsxjO3ONjO7yqmXrDKobxv/vl/Nw5MrWBe5U/ncmdKdS4Ts+Ni9y0fOtoIaD
wfJTWUSDCKHOPUT3HMBW7Ax3WHIqifB/KlxvT4JUczypZdatWOYsNTz6NbTXjEyI
fBu1xyRsUm6+jR3UjeLW2x0lUibClGC/gtDprejnpVjw4bP7QcFXURoGJXSpvQsK
PK0vk/pP5xtHJicqbw/lkViXe1ypMiujyrt6YmEnJAmRszunKoffOfoVu7M6LZBv
yHLr6ZQ0z6jSbnXHWnPi339QoOFIwEldxAAkN6iEuF6zlTMlu9mJc8cbI9peUROj
0IArv4JvZFX4nu4ddad4gTMyA0NLv4yedfD9NM6AtK7i4OEKhBK21yNslC9w+3n7
VdW7xk+Z1A6nxRBEoB1cCdDAS723bQvLfUThS388M/YgZVYMQKl4Wj1afEqLJXtE
VDu7PTWzvOJird6Eoklpx/aS5fznU1qeKVYnFkoalfp53XTciA9nUBNHR21t4GUv
XLb2s/r3AFsyE/a0wIhJmoqghEB+yNRmNku42O2bqAAy8G3UfwPAxGvqdBIH1mEq
V5TnxEuL+ZUi1nj03y0ixDNLTd8QHOOvWZ56nciuaziwtG99hydbLbrqsu0EV+k2
L2yj/QoYa0w0Z0xaQ3aAXg3mnbXr+QVXlYO+EmPvv9ypFOqAdnnk+xSSvhtXy8+G
iqJh5CDB0BCeDj6lwtYGHPRXCaY+oAIVkItUs1hToiGvnHPzBSEuDQzFyfqob/uq
vJb7jrXq8/u1KHNR8Xbx/gvfKDOT39BvOPKNksNkT+IOxqH0e+x6lM069FOVxe9Q
rIAvKLOZCXg03HGwZgAug0ZepLzpxrsP99VSlT5Cd7jHDDtu9zxCyOQlx7Dn9Qfy
2ceOdoGC04gBlkK7UVVag9075JmGvAfjFs7Wy6qugB0AuvN2OPRZm+o5aRrcVWM0
lMNIrCA4ctamXguM1xR17l/xpIXdpUvBCswiewaP33cSfEbBJSet+kUw1azIGEju
k/DbjRl+PQK8fRZF/rFqjPmqRz2KPTSSLZhX8eq5W8LNBJh/P0Cv79AOFl1tdoYE
RxqoiXc4rKTZhg6OWBNxM7Ba6DxT8pIFA/DY+ue+Ut5cjRoC0VfaXWj8Nl8c862m
JnqWZAYj5ex67biKyVepWtjEkcLi5j6/5KS7ep+iXclADjOyBgzHEDU55kA2oJ+o
UYOb1Y9L7p6gyAsWFrwhe4CQ4TXIxNpAE/GsHl+PQTcxf6sLaHziKFEtw1TSE4LH
iKIueMpSAt8E0DH/11VnVgUBEypOP+Vc/s4F+2OPenryzXK4cwUsolS/y3nQVOFS
qUxHsUD8oj9EwpOGuK/7cLdK31R/A9elMWZAqfDY1dnPDPZT/6QV2IDAcoZm1DiT
8FwA6/ESRiVjCDHiIW9Pqq5osO5e1koQX1Sg+p2JAc209IYMkigan2E1gIHwITKL
v/rDUyuQAsrMHPcVtQ/5zEMfbbHD1kJ6m6w4H3Dwp17/9fG4B1md5JogM/tDK+//
r4fYwiZwoGuubGLLX5Y3gE2ClsJ/AjUzSJpaMJrbO6W/ymLENG+7xti7uLB2quZ1
Hao4I0Tv8GgwOiNYENChb6lUQ/fHpeINCfoJ0c/s3TYiDoCvoFH+0pog1RtfWmoW
YDrFg+gO1CSatCq7d1MRPSewiGrND5BpTvG45tYqKa7spcFUcsOVpbzO+zhCbvr+
OF0p09PmBs2YguZSmejEV97RD7xV5QQ3kN+rKhsu0UlPprGWqTOFf+pV9y60cesN
eyC2+uJbSmkVt5ZJbbRoTwwgBgG7+VVt4hwraucOQZmfSC7F10V69CNXJJlZ0zX8
tSnl9a+w+wVaUscndZadsr46EUhmhWyLyfTrKAK+htWxBV48y9OCWA50rznpi7t6
PACLbjB/H0vXxLyPQ1SJBLIytKoAU4T66LbHILGmqa+d5L8obO0J1ub7wcvAG/oo
wPsXKdU3n9SQLlVPyZHBf5/IVq2Umf5nxOPq3Lv8zqJVVJ16x32bVRAmM84tWe9H
iAwphFrhZs0vsliIco/R7fiJQ8ZCVAzBZ4LoXBZlYoOOQ8e0RdWXJg0Sk6JA9Wmb
AAPBjrPas6+vI+aMAkHnaDm7EKkBhqjuRupWrqNwMqRkOyg7M+UYIdav9TlC+seD
S28p5ayTFczzGP+ZcV9DqVjI+1tgO5xn6p0v8KKaKGQIdHjL8NVnbzFs2aLPF2D1
nBFl1sK1MEHcb7FNpgwDIuTk1MoAm51l8zh4Xa8hEK5M5CBN9gmdmAlAf0Lnjf1D
i9b3UsWI1vBat5La3WJNv/g1S1le/wnJlUsroW2rjxpEvc6ad+dluj3wzEqxmPa4
DUOxPgWi5Q3UCvRFxoWiYJnVo7VA7MoBxQWd9td/YP4lLByCM3tOJygcfmmJLIjM
a6ErsMG5OcIspAG/N3tOAavu4sODd9ZPehdVQehLNK1njSHiWBkABCbdd32kPuXZ
SZZeaTzf8b7DrUJjUrg+iHv2qg8D56gMd95QDjOsB+HJq0pOLD/kjrBGcnweFFDs
RLNnFJBC6d5Jx30C0oynJIMMk40BN9CyHjtZx7c4InSHdI+Z9YJCZa86kJMir542
SVOBCe4QgyioliG3KIDU7eSlPdu+SKelYnqiT1eZcsMHMxHE3hHo0Tmx7uGbyySG
ZsQ+n0eObzZZdXsuzlHpfCt0XbsKDLyeJ8r10g0eOBUvE6Ohq4BiBX2L2dvjRV50
BiNRWRtlKfvG4/Dtl36sxwpkOrlZjs4uPy8gIxNA0TdXoWAEkaqZpIsr+5UO1HjJ
VOft/fnFPRuRhilvhF54kB3gjFGBzNjkYOLNINb/+eYiqIgiiMtohigSYJlkgNqx
0Z0uqBS0CLkVIltg6BvWX+35EM1FXChXSpCDljeD6susMh4/P+wxwNqq+f6FNT9q
z6Q6gwxmlMwz0GbLpvOkjiux4zzfGAAgYKRA5vQMma6tbAJRrVzKbXe3IQyho4wW
ZMUFqgJhfiZVKmcyhemrtoqL//YSXKCz4324h74WN+WvJVA/VFe3PvAAZE55BflU
TIELEUOF7ntoNTxDSGrdJxiStLjNIOIVS/YoaCv/AdjlcOXLlAo3MSn4cBAOefle
lgjA96hiLadhSF0eY5CoOUxgkQIWVVsA1J6MA2Osk+aJHY4zpowLMWmF7xPn8o8C
A+l2BwktHi5csnJbmhBBnXu16pBEY77VGX2ZcmZpWIJNrnsk3Q3OYz2UyufxWwZ4
abXikJns2J8O1bKVKjeccU5AE+JR6jtZqYbZlWfdd9UW4qM3no8HxO3xE9dhCrUW
be7U4jNIRClva1bc1nbp4Q0j9YXSjOyNKY5z0XYuXAVxWoTcHSVjDKcr+o0Mv98U
apM0vV6nD4/JnfqUjhNW2GS1P9N7hOXw4uW8QEvZ0oB3X2nb+FzO6bgd1Fsef/1O
cYFEyzcP7MWGqO492wt7d/3O91rtPEpKPxFXEqbZ38LNusvI2RZexsRPZbv2KrQc
lMm6ugTxoDbCZLyDBLkryT8CXcCg1RFmGvHE+E19Ihe6fqtcW3xv4c1Zg8uvZ/n3
GRqYN8buFWncQSjyRA29EDq6ClMyzrf1t7YbYSeLGeRcPZzQ7zgnLxuWE6r9jmqc
dqcwNqqOXvjY22t6mEu/CZ9jYKCodngytHUYKkQyINA8o1+qS5HNlXVIqjb3UlAU
NZLbp5o60X+4c91RxTl+HDrOcOKFNZEtc5viTqoUkMfoofT0U5GNSP6AjxrXJOEc
b7IoRZjDg1I7NbEdlX1KunscwpeZaIXt0IQztCCYy/Pd1C5cdaQGu2ljinMGr9+2
br+LHCEa/bsuSI98GjxVEIDrNihlwG7lYE4mh92Cdb1qwsl12X7uwmBnh9HxPO30
gGh0hibsap3h0mXKyHsn7E86t6eWNHi3O6cnNDyO8uCrwtWeFOGPTFz+4laojKcY
F/MjGtPTclvCqI4tQK362zIejT9aW6NkPk/3nUNVcoZqLLs5YvK1UMGIYeOqsTuO
Yp8Ekhx5+KbAAdOYMmP02DBxEWXA/KC3jdwM7EVQ3+MrTQdcW5wFTzHtv8HSahq5
3JYz2GiNY8eRj8nJLiS3oQhJWDPGGxp5kj2gM+2CsGwD704iAUAWWQc/26/VBKEE
6KNWeJ11NzTXBESvuwwc6GYtijWx7XlEI1a5Auyj4gY5VZ7s3xMhkOCqdr+c6PUN
vNPyGFLvPfZTqN+Y3spa+FeihJN7b6f6tFNH6zN+7n/q0+obTwtPcC5otoyOhNWt
BoxRkUPY1GLLLUPpXbRk33f5KZFQpSLhZKxGD3g0Fn3XZ40Doc4AymSZjqnNhkoV
PjJgZNKpwqjCimht5+aZO1092Rs5Z8e9Hr75Btv+oNFCk8DXPlVeaAT7f1FCdrkg
ALpvLL+D71ITwLtnJFkg4gK0WUWbuMyqhf/Jg+4jjLK0Hf1cuKOOPwWvcIs5UWxd
meL7TjwkVonqxPtch02WWd90SsFlbxqxbMAT36ShvVbZo84E+9G4JKMb+p+CWfnR
A3GSV6KZvN95rNM2N7oPYmtZO2KSVPbGlECa9ep19nwCd+6n3nCxTpJYFtGQIgyR
RkfmQdkkatT7xjsXPXYvNR8SAwnJQuW7azF947nszCfrgpQoivSZ9NSXP2dm697e
R5OD9MA72A8sMW92TeNWjV853tPbqBk9XvY1OC50J/rp3mZ25YJWGLkMyVwX1rSi
Ht6frWrTiWjR0qyHT5AEhqyoAyt/TDRi5mgunYOebiLlCqo3tQN4tDchM+/rA2Cw
b6cCoj5vBm6PaH3Ah058cEdvK5uOvtY9DOOmES2c8+kjTQ9Dby48XrzW29Ue9EQK
b72PE5aft3yCjMmP841e5+bpmKNwVsalN3VI6eFqxQl1nD+oPqnjK/dpMPr0D4p2
YAM/tvOc20kzTD7puITUlKNSUtlslyWshdXgZ7ZsYJiqr8vf8N0sx8nZ37bP/8ZB
4LggVFQZUdqrgCdhbL9AAUV5l99asfTQKxEGBn5h5nrDwxjRm/tSR3lU6WsPIQSY
s1C/ibmy231EzbFdrtIXZ+dBkvDuPl2w/O4sqIt+MFshyTOz1eSYI7XPWkUPGAUN
dwcVnB2Fv6PtwB5dYPXGfQVSmvb6nywAMVNiQTU+Nbs/45X0qPzqbdqRUTe+H1ga
bqcTq/EMH7jr2s4CuGY887OyZsingW4yql4/IQhs2HnBGdUY8y7uHmr8iDGUZ8hN
U4gnFxDEXS+IizNxfniQbMGH7uBce290ofTs+UMyesy/mxCGmVJNmVbGdAbUwYRf
MQ/1xPDD6pdZxz84bZKRpTRmBgqAUqxJMGOUykz7e35I7BhlFOu5s+ywSt6YwlwR
L9/zTW/gT7jSYArMMomryRM8k3q6ojhhn2Ow7cS/UsMm2UVxBHjbQ2L7dQ1jBg6M
eMw6wCsMavzg4QXPh9asoP4wMcvyccELZypLTbDCnnNwVecRwlT/AwWB6PtRGR0s
e8lsehXCPtW36iz3ZEQnj1Uqi5SCc1DJtpuiX/6nYKQqNXrvFzgEdIh9okwCycTB
3X/sUr64EXzLbH28gVUi/U8P6YygKEmgHbtBu2DlKX147VGnKmFExD1Mt7uGhoy2
MxsbiurQc5ggVi8U7bhlFmAJkyAecyETat2PpfqT0g2VijpyLlQ6bmue1QvjshU/
mRiO/ah77Z2jLZEAA6f4ozSc5Gf+oOssQiMrAG8Tu7TKbQdMbrJvQjikmkWDY8kM
VsvbWFPNVnyAtVDE6Z+z8T6a008tAryGCnAfMytmbL+c304LRJYtlapwDu2ed++5
vFT06g7kEWwlL1St6XvZB/oJriWNNt1GBE7VYmQfIlnX5/kO5d7h+FaJOy5lwdFQ
aHpdXox0UR7zwmZO9/WmiPtr3KjPpTPDuywpQteFEIPRmEtz7QRhyp1KfuatQo0r
XkxF95SCBkTVj4hZfWCt2p5mub8vsmMKedoVJ6a7N/IOV5aOxiPdAgLCWBNdXNq+
NUUA4J88Ecea+4fIAWy1ffe90dyvf2YftP0spN7PL1jhz6YDN9xo3KcXgIq8V45z
XlMb+/KpV8zSlW1HUUByxhDnQ+XXAAxcY7j0NDvmrnwoepYLhSeYtxVvV/dzSkqK
54MBRN5lQ2TQV5V/9lLWCQMmXYmhpo1e05qN8MFuqGfhNu8Qwo31Zl0PtJ6Rz/m6
TWUT8RuhveWHqR3mgCx2lnCA6RgO/sLEX2v2+VOkSXgT4cqkrsxGA+XKboavfLft
jZi9SIJARX2w9Qcmdf4l6YEbGMAd1RLztSqXhTL1aHpfqmzYsEVVVNMQX1AiWSA0
U+xUGORKCzj5g+PLw2nMe51XC6bbVWJ2R3Yc0obyE2FSl01fHLEPm2LrXCQoprOf
XwNQzGaVAkRkQtGkQ4UyvyxoAVNhSF+GcyM94IQpOHEglN+AIR6r4uUnLubJD0Bq
lRWThKLgPrEkWgBRPGtYI/E3qE3+khfGjbSCt2mA+FKsL70dQytVCMlzecXpqKfi
pYG0r2q6iJrxTGpKTYp3TYuUgeQrB93uE8QTSZqNbHEOw0ylY+T7aMkPbKdVVlYd
MD3VSF5EMxbRM2d1q4Ml1vUK7guv7wsAJMNcWAzs3+VgjVuAf9AyhF/dCjd3THbh
Eq5QqoHExetctNbXQASgiPCxsgKRL6a6nw8j80bCyGBfDNU4HjNN9BXwMqeHEtpd
MsQDAWA9abfU4Z2D9RfMyvk071YjzOwpCLeOiq91dx2GNWMVwn+oQOt3jXcZgatM
nlbtg2fAfG9f63jaT9wyfV8yOjVvyk7lqWzpwqpS2brJwk9anJYluQWiJD6oEKwg
BGObfzzzZFBnVXT3DuN3ZF/cWghlwuD5TFkSmALJft4zYZZCjmkYgGRhDs/o+F5A
yGZrIzAVTt7zq35x/NVFUwe6wiZEtB97YnZsSCzsEwuD4p9eBfJmDG/yP/+42reF
+K0rXAj6iFHpaJXn5LmVUjP2Z/ol1dDRsSAiLAVPg8BpWnRiM5LkAnyiR/8h9fEl
WJ7B88dFyHUpFOmgKkV/T72pTTMW2YlAqD4lB2GkXKSa7oMW58VIk8RWDJLWiX56
BvXFOZqgCD1DcIXWGNRaNC7MkqPoJB1iE6ASlpST241XsFMD+sP8wSO4b46/IXiR
6TBRm0ltqRJYAuY3tj6UnUJCI0/xO4h9Hi4yDvzsRC+5RGAqEwIYZJb0yyzML1IZ
+ABcjvndylsdjWGulH0DbWJTXrgwPiFJo0e9943X6m9wMXTQ1gLYwKi9iQVj+uli
pMA65LaqbnJZ6uMNhYYdhgnGlRMuRo/ySnzaMHlMdZlB6L5O+Pb/s0Er3XLoqqPI
nOmZUlwEYBcUW/xoC+ncfMN6Mz/D5SZnqn3pfUQiv5Zit4znWri4ipGPUERTcjiK
CbpmFjjteYL1xSM38ICaGb2Bvrg+5sH25/A6FOS4wPGDf/THhkAiFREvdmCFcjeR
kK2V8xuGqmT7x8rHRJSCp2SPuIiw8DEEYa8nL7TSecEMQHgvCUdevOctOnlIq+1F
fWFRyyPP/KZdZJs35WHEW7FKEdCyx3BEDCf/PJrCp3WKIo6ffGbOQgD5MjchptSR
wwBB3KX3l2RgMXcZO0KP8rFcEarCrpLKx2uzfDUeshjEnAcFjefDI4uhlLYzVg1w
XMjv8hVNOD50q+fy6siVUvEc6pnM3lvLp8xC20aBDVca6OqrbrXIU+FhR2qr/v75
urk6LY78x3df5mDxQcB8sImmUMi0n4NhaO0XNrbAvf4PwVhYEHJLCjl47JrFJgyZ
kuG8UhtTZJNkh9mtyEb+anOkr63slVla303JJcptqig62REO8LLT4Qsyh/nhJaTa
SJUTXAd9zTau/+SuE+qnmZ76Yp38FqRqGbRplmDnFkraFipAJlPiej38PAPfYfYa
b+iIMq0QTvfkAPl73h357oWJvjuHKG4V0PiFByQjYkrtKu25kOk0U48eydGXtDx2
ME6HTvz1htRZ8/v1SG6hEnHNXJKuogNuhFI0XFYFBy8JQani+Lykjj6kd0B2SYvk
pTmPt59fD2gtrjodahzSqHjAwrWsVsxLBzhSdgXlydlJVceSFWQP/U8bapw/Tq4B
xm1Ua16VKqs+wCRMyIFz8EEnQ0WydXh+eP35gJwc7CLrFDyLWesnpNcJB5fEfNyz
Nxul8ZZdHLHM/hIghe6HWa9iQtNtCX7WgyTe/2BcZlWJTVfYNwfyCMFJw9+CRkXU
tOx4t2gnE+lAMPlJvjpRj0uo16HMmQKePpg384NzQrrwYP78WIkAd5Mr2J5z9nFG
LHcTW821fn9ggBWKyPCAUdp+KtlCQvNvbn21NMElQHytdzHRZc8dxKtNHbQvfk04
p7PNyYZ2NAljBVScEaWLL0o1VyLWndLXSSf3KXcxwBOaEL/im4mE0kiWM/soDMD7
y2Hc70W5giGTZ4FymfNgCosXFHNOEF3fWfvgGb6/Y6XOjA6+57xaocoVbabYBynk
wcbj3zXyaWGu9PuaJ1fbcPUI06N4tlB9lT04hc+7qSH6B+1QJ3Q3efR9K4nEBaoT
HS9cTYSWj7fZUytkFadYQG67UlUY+1Y/yanhRLaqQeA9sCEO+klaWCwmada5T+KY
1Y7KRzeWvehxp7fPrcWnnYzGbVCl6XjY9chSTEF7jog1ZafIeifSBxaOQ68WPlZI
ESJPzLRiBnx8HH5TSRK2LF46woJHUTPxw+tKeW50ZlbabFDvSYGBG4IF5w53t7Dx
wY+3Wieqy6QhCVBX+/RAObzHNAy4XwUo4Uf0rYo6wVFODHUPCyh+De436X8aOLk9
8OZQBGSwoBH6ZLqoW4i5Z6IzGJCt5nfFDrOMIFNlnIUGecV8UiTRxQCpexuKMzd8
+V9hpU5WFGTesH8xWG7MeIFbFp/msfeU8i7VLFG/rl5S59jcL06q2LEGFPoIZtiF
6o1M+GzO38ghM1oZbH/upMQHIyt94mkhDyFwRRThxW7cO45lkSKLhUghXMN83dr1
OqJ+zJ1WF1aIhS5WyhGnXV7DMeLH+mARMYz69LwbdzOIoWICUEFOFe0nyY5jkgDO
qj6LSxCmQ0JKyoYxQMqzx2/oLET5Px8fXpjDcmxscTFyj06SLhHdoH/eepDyzscl
x6EOUH3Qp+o1gyvATxLRYyHtcrSmKh1RXpNtdb4OKzBXT/DRIVyV6BPl0mkhSbkQ
t0e8jerS+fvKnL2p/onWDS5XE9CM8BjOe8f9oVhBiVUE884F9rz98VOJpbEDT33C
/WXHZY1xJ6SHhoiyILZ2ZVMiYGmOviwdb8glU7tetI540i7FXdr/HJZn6+OVpGjO
JfWy0q8HlDt0Kd/CW2jvAXa473/l3kgs8PNGAtj4HTQnzWYkVIgmOEDx4Myki/bG
zRA3MN2SLYFh5lt9mteQ+EEA3/qt1zqlrSOQt4NinY8MTduOnHtZPTg5cQpXHK+2
Zza7NSZ/su68ee47VPW4KWp4vEc1bH8YdFzT92MX0WW6d4HdqlpBMQHbDF3pasIb
8dWjPX4IlNUO9B0PAJeciuNFrJpYHkcEPd3Kcp/F0sEYVmgBuVpTjcl9ca/isRw4
SYAfTkPWUm0tXRfzjOwSVMq6QhoFstyswitkGqm4gjqN5UfCirzV4SRW+O4YouSL
0qXfwI7mxk8BR720jxmA7TVAVBxXTJ+J7RP7+6BhScSd+aERdZFjJ3kxbrgMxdKc
dl6GXgqqJ5jh1agwaA1PxEnXAS/MYSgiCwSReStBmwAsCFxL0EqDEAfq1jvFb4E8
HXFunzad54NeBDiDcZVYUA0tGQOR2VuzednwaXnCeuI2BJ9EK9xcITrXdIylzKZf
YF/9bu0lDf6v5Sm0tW5Ud2kBpfu6ARBzY784xROn2AnTa6p8e4dNeqlhikKUeQ0S
4aXyarxeKYddKPIxZ5aZVvBHlHeOANKB4mCIWQiLb2qjemxrTrhHNrMHaPC3tOL7
hmz+Ec8FOny8vAMp6wymRMC7SCdRa1am2jKTjktmHU4Q7J/ea9bODhSLZ4hR0Ndy
C7DVpvFHddeHXqiuWVlt0t0Cbk2sbnvZKXW9UvEozPoY2Njcg5NeFeE4KH3bWpXo
Xyb+J1s/g8ZsnVqeiQEu0iouHpbnlEQUupdbz32cP6DPGJNcEsnQCqzXkbboOvEE
wvrsaTJBVvkEOrQVrxjj3cq/dKLRfOD9tWZLCXbkNltai0Q7ayEJIFO49egiAmFD
Oak23KoDxO0xxoyG3EHbeggI9QPtIDffpqNTqfyH1Ww0DBnQhB//P6P+eSn5uFZv
4maYcJETYJaAld+1GodMPCMZ5im5B8Tpx9zHF5lVXtnXQJOLEBK8RzkZzMcL/RNE
DAFAHGS0f6pdDfeSVuny49iEIjBg4ZFXcFi2RMVHHlByRE6DF7eGaEj+WahNLbJd
IdY/wc4cA2J+Dn+IOzfvwARNXiijXqLhynr3ebZl0qFy/oVDtz45jtr7FLf6z6uI
cIPYhr2Nxwr4Y1nxCj6zCeUNkXPIBXbJeItE5IQ+22nlUuOGtswjN6hhM8flxWjE
BxaLsMrJ5DVMRE9zcW+Kf963G+6RGbXZhXwdey/WSpxgyPW/+olfvRNp40Kmgjf7
+GnjDxHoX1iEHEe4QgwDtDTdJhzRWI+7tLoa3635VoikOWr4vR9sbUQQk1HWRUZQ
2NLNQArkpleKzAx5H0eyfzT5LfdUH9rxWmGtrSi0DUvUZuaZbNMRemntkHJMrQ7a
QKd3QkipxXJgoJBqj+3VhV4L0anw8YTJPDRE+dP0ehX/vUXP/niypEF/1Lb5UJGc
59zRXsLU0lqwTcjmm4THbSQRShp63/7q967EMl+tYvgQ+Fo1Ab+bY6P21QQNetng
f3UJmxbasha3urKhHW7ehYO2bzsiaFYLYm5/thTX8NQnAt+XFJYRrq0Q46pkr+yn
67vkut6TcTBuM//pOdS3eEQ/Wswb6GWAlyP4cuAR7VEpEBtlvQM79AXxpsp8CKxd
47jdixz4grViN0Cse41xwqiNR4g21ktsWUS4aVQu3TvDMYtt0Y4CRGT185V8LI09
BCwcT5FqNRhBqdL1cSmuabE5gxvZmBWiF9OOyIMBASJYlsDTCTJZ16tNn612Qqly
EYVMQKbge/bUDGvihVxHDM8XIHV5+CnYa3eNdvKO6oitd/txwaeKZSzbsCc9xPDy
RYK6Ip0h63PsxhvkNPlvrF/QUFBEvXC3TlgWUM22Z+6jL58t28UI3GQkrbtsJ0Xs
z+EkIQZ1/vXb3qXghzuQCVzqQIBbuHULvluBN4/kcgsT159BCJd1cyusKhOPW0ez
3owXyY6DO8Ioz3j0Ri3AS+DFhbfxsp6ZbRiTdpEsovIoZBoeDYhERKkSQn6gVuJ9
YWD/r1S+6lb2aiMTSaTXaLPZg/CaBwvN7R2HJ328g7BFdqbK39vY+FHvURXBSsXe
7jjkMATszomC2ch8LhKsbFFtV45orWEwHnAaQsKVgDnnQ0sKilpDxTJgSxcA0v6h
wHd5zNnYSojUq4ZyK0sD2b2Pv2RRWAi7a2lX+NCuMqKnqOTCCtioXaV905FUiK7U
JwZF4xzmNKxJYqzUpUcvtgg9nk7q9kliDF32rx1WeKDoUqDViR/UUpYs3di+OdVT
0HikJf7+SQc1FdkwSxxKx6JKQ+OmEzOmzO6W0lWNw37obaNOLBlJBMUIVyqrJqUc
9ijJ6FXkXulDuFPFVJvEA2brEHDG0bUVnLpO9va1M3iwPxh5S/JszuuL/8MSCZpb
bbDyB5jvdz8hiAet78Xc5DDOQjYai7OD4OmxALbZO8+uXW8KMXioNoEKfR9WCclI
CXlVUJRe6XUgm5krr8EW8pEkMP6qTN/r4SCBZ95o30W1n9UhaZ9QehkKPyno+TBy
nh1PrNeUdu8uUWXvwIxmypjmfVu+YziuvawnMM26ZihftR3sWJoYhKdsBKjy1Z+I
iZywloL08sVmsYUChbB4YF2iBYJ20kq/HBslDkK7wrfK2DllafuFjII4nCjGmXHH
dEuRm+HFKXitJyxKiHPu2A0xjBxJjBa334XRVWcUYE11z6cir1tTco8HHaxQ+0Ci
hlrUxIj/9A10roQwgj/shJsEdF/KeCSnX9TW7IsgzGWKA6UHXOGwg54qsKBfkySV
2zGmDPltzrN7UXW/DswxdKT6ftAsPdn5QyJuM/sLaFE/AVuWK3QLgRjRMSKYQb8E
rSWD5ThQbVbbY9UD8kbvn6ltggiqXjZmXUxSpmcHsMs+eWWZ9XsztVSgUFhDA4Re
BK1M+r4cyHgdpDcO7ZsdbPKbLKaMiXc2w9YtWHBozMVTkMQ3z3T7a5rlRVUtS2J1
Ad4y9o6yUV2GikoyxRM8cl2zIKcHPfEFZcPBhR7MXTE/efK0AhIn8jQJHsEv8XVU
nG28zFApARZ+ooXP35ilI96rBYLS7ZjtaVmg/S/2sKTq6npwDmL7zOBbGxoYlVHg
nrsQnzwlYBk92XlMKF6sCbAmZ1jPtFoH1Be3hj9Iw4ag8t8uOPvxHASP5nnshJJI
oEeH+/yxN2S3fI4Gkc6t7g/VnTwM+y8X2UN8ulljCwl3JwYlozfIzCXT7NKaYMA3
Oek417kQ7FS2L+zANW770J4d4DqvtTu6wczLcCpZv79nse6R+WCZvcq/FnKUOpE4
/5Cuus1jdImr8Dpczs6ve/2nDwdXGxdm9dDMbGf3iuY79cY8O6AXuPSMFFOJfrTN
dkWCVUaUOmO4/f1LQnJF2fvAytP3nA8CStUuYm6YLK18Wvd6iNywiQAPRzQwzIs6
cPXAQq8ZHLzuQNJ28m17g4SIMJXGZLfr7Tuw1r7WHlaA9xs+82dDEL3+oNK87+hn
GcbTiqBgH7f76uyjoHJpqmjOisEiV2Dr8EPDbsFT2sw31Y8EUhbfzlJji9U34XeC
qQIRXJvNg9hy4sgXqF88CzEID29Y2aYr/nbV5HBUZMuEMurv5/62R9StImYIBGlA
IYhvGnSqVVAh+mMihzI0oHOZpB6rY7gn99mwR+r0HjegD59GZDUJ9ko0/Tezs3ho
SBddvEE4BkJiucxTqeGBqsiaLCWKbrB0pAqLFT88+k2v9Ajv/XcOE6aZwjARC+SN
U+StCeoSwzPkFOtmr5nOTDGrSy9+R/tFCFqDliawWR2sK9aBN4PVaS7GMd2/UyIo
xHw4IVm14XZb7JRMoI5FK9sbgjSocdY439jDt5CCJDOsfCFgfGwEjsP2BPRoM+3s
xEqo12CJNQdKV2QW6/Py+6f5RkpRVPu7CLxfEu9n+rAwcqSiV/Y0BsnN4fOe1EA8
HV/XxfgsqF7rm+EiqcqwqQ5bgBaZrnfl5nwtKJukncFDkMNI0Lv38t/FaE+bSVAT
T+E87+23L4mkKNPp+mNVEEvzODHWkH7vkP53q7mvKLu1/LftV6Dr1ev6KZFQHQSa
Hcbf9TRskUdRVYA5x0XKhnrBuVk47Zc7wJivrX7VXUOt8OHWoYNZdA3kN4VaHX1N
nWUJNMnfe+jWKcKpaxKfik22BN9zhiazOiGyjcmmMlCc/0fmRq+eguI1yPeB6SRA
MGaBjwc6+inEiAHnZQSPj2peIwUOJzlLRrSNx8JfK44/H7hAtLfKuMkzCDGz7QT8
d7NTfpJZ7UVEScVBz1oI7/64wNlIgrjWnXbufyB26odV7tdOWGMc0TsATsUT/ALS
xFrHJgW0QHEMtos/Ok9+tG7kkDhdqYhfwsVX4qFXcm8cT/SuCm9+4HhyyPeak+oI
L9OPYYG6EtOTKzkFXqbn7OVeiUZTaFowXKoxVyGcx4H69RlpHH2z4cQOVaU8d8BL
RFRfx8rcl+qjJzJRwq4eOvXNAoh/ptgRjMp5GL3U5G8XoJT5vC1l8zH5I/NoxV0h
Jpuo8KoX8hnKLpb3Vb2C8Euf/KbPG+7P9P/dEBQMVvCu7MVAFOS9RpqP9bXx92y/
eCTJcHUK+y1cZ61CTDFQd3msZNwXrH/3rNRRyS0Vp4PlkvwE0cLW4LwzKl0E22LO
0KAU4vh4Ksf634DayKJsYK0PKlpFWCvsNWJSq9EJTINilM0H1E8s/2H7qjKmEfu2
jB6ihWWPsn8XlP2d2nOH8xCxI4Gzk1WO/D5Vb0b8ISUy/JM155Xd3ZH9SRS8OinH
kG0g18dooinUIumzhB450j5r3dv7gd/95MS1+1QTsLvZjedSDdXHNme+qWfCZ0jD
5Zq2IOTt6KJMAn0deFSIOt/ILjnTtjDzky0ZuKiNJ6Zq3EpyCT9kTn0IEI7BYe/A
6WurqoFfmCdFBas2fEW+NRrwes8fqTNIgAAwifvalL4AEnapQZIqxd907cirtvJS
rlSLYFp/5bsoAwpPOZqiEKk3p+ofX4HMNWsLWZrld6/eaaTSQim68uvMZAXZe7rz
edIuZynFjPY5qNthebJ34i3oU5gPzB8Ri8inyw3KAENPgNWLetfSNKvplkyQLnvq
UoQ/hepwJo9wnlfFYo9GRax+Jx+FUsURJsEjZQOIBO6MDwV6gmuu9VkCLAVBWj9D
uY6SqPCnbXcGBiOUNYyL9nOK1KMIQEgKC5wrgxJGxyzHmwdSWPagrfU3BfMR5Hum
PCetyqHkIfuz5X1IKvp44IZUQh2a+M3m2WlpBTdIYhxKG0xCOml154EFo9zVFmLZ
z0ykxeH34aR7sB9rOtw4PzxDzmu+jqldQ35MaKO8psTA9KIOa7nAzBISDPYmcd3h
Lnb6sMqp6GX0hMQbuLA2fJ4dMpLf7uhgdBFq9RYPzBfuN+ucVeoQkYmaMXYvlTLj
oqg8zdF68ZrGkWZWbhktTopEaB7poxYEL5VyJkj4ZYaM+IUgPR88Oav/DUoqzrd7
HNACVG6feTmcR1FYm7OxFABjbTBgsKhrrnM47N2LlC5U0a9GyZkCvllHHZOrfhuY
4zCKBwegIG8nZj2iVDy+k0WF9ctvLqD64p3gU36o/oxEJmsVLD4G5dJ8EhaHVnQE
WH6DMK1xYfXwWs3Z6ERkebHkysCxi7hzLUpoDdBcQpFNx6lFHT/hOso4mvG++lnh
VBVw+Kg3aNQIDBFoqDxCYFPmvF1PL7eNhk/QLhI7r0J4zKg0SF2YYb5DeG+A4b5m
xhEg3D/GChZmF+QS1T2/7U2Ob2EohFm+8jm6yJ0bw+0trGYqVOqmzx1IJo5iMEdM
nQP0d7GU2ihfM8+6gNMXodFqUfrOL3lFyXvwJUGpsWxT04uVCTcG6itPBr7NmO0E
aKXXKUiWMsR0HgAq416k/B9Zsiw7QW9jcyJMZAeu+gg5s4z209+2hxBjOsmn60mH
dj8Vl+K2pnDqZTZeJ34EH9/+ah5Pcn8ers0yNNWsxPDGaPRD39HQwrCiBCq7zveF
RMQ4Gb6D+VKt3MrN+oUtbLLi8LbspM1toffc4/6KNbhIeGxPZnboDZ2lBExRTKTh
kFWAN/+SjXypXNwVMB1l6+eLVyDgkNQ7w6gDze2zX+vrVKR5ByNHMeMzWk3HC1ZB
LbaE+PkqeQ5D7GMxlThe3gIKfkHB4OywiAlvkvkLJnxm82N8qwnXXZ7M9t908mYZ
+ZeokqeHDhuhD97kIxhVHYkrX3ym4A0ZO5NPlRx5PIOtktXkZh58T22nZX58g3R3
g/IlApVycG4YDoxTJNnNxx0jBYjzRSSg6eT9BDe9G0stckNApXEPMLEGwgM0rl41
xbgf0va/7nOLY/9KrmryMYrLJsH8bZuvdWj91E0C06RJYkJbwWgH2xt/BJaMqEel
MuskywI8AmJOgoAYklE0LImU9yjyOOBGQ1+NHVfPUycRaIm2q3uXgcvx3J5TnB9B
v5WmMVTYfk6Nlcu+54vm8dngBqnzAVVDIHubdrsgISrjK7whI9zHM7aBUF79uO8O
lO2Cy4XU5nGFF1+WrLvAWpVfglTp7R4QfDuTJvHvCRekseL2ju5bMUmjBQEFmFnl
MZj96gRhiFZMOlg1xRPuPzU2d24Ye1QXPwTqlJ/fC52tQsI9HFUZjsVzBzQu8wwt
imX6hZ0+Pkbrpy0PpbfK2nAmP5OWmOd+QEHJBGL8y6R9PT8cw6v4vbIJJyLZZOII
LET+SHGj5pAFIL5G3m97uhloOnQ0612IRTd0guU7nnmBCEvs7xa49Dxhr3ayfGiD
o2igSkMAzvzl/UXZPuNSuW16UgV3LoSJzFsUFbMw9+cpTV2CvSSIv0g8uQ65eVWR
gCFNLoE3AXrwc+mb7/73deJE+rTDipoEo7nF6ug/NErxlMQd8qk/nEhd3/V4c7kU
/jNYQLYvN1sXJd/O4l4jyGF5WgUYo4StMBuiNu5RXzsV6w8V27PoOKr/Tx+aKGZ5
QdZiuEWvgAD3Mg0N8u2NdB0INUYGkCSJ54SADKsw6gK2alZEI7kGhRkz+stjx0/h
kYDJ/JVIT9/CJ6fM9NBcuRLINue2bxUn1itWBF+VHsUgnN+ZnTiTia8CsQ8NHn+X
vjpfNFPULX9qZQHhEuO+WjiBzqkSPiC8850wpOfb0aLRTTYuQPrSX+mUdyFICFZ7
x8+v52j93fkaC74XOlzUPysiG59YQXDqZ1t57SqEXw/GbMDNDH4tpy9cGzTZKZs1
SPkBlWuQzcpFrFMTB9U2/6UsFt60JViv7SbptZVsAUo1Dsp+FVIEqigEQ9Ux+t1Z
xtzSsxHZLZxyu+S1J1cjEv7Xg/pGWluz7z/D90BqUoJryScZ75sfMliYZPtDJxhn
VRfw3BL49GwhtuGO+HoTVhrUi26AprLnS/jHuwL9kynB+HNpzN2tKyCtvE21RBsN
SfzRvXufEvsBdJ2d+D6/fJbIyScHjQxgWW/r/glR6bkF7/84/zkMz3b6ZKmUqoOW
8hKcNKQFvlq8n7tIYeOvDZVvMNnAxR/BlPJg9raBUBY3QBSFDjrUfuGGzd1WyxhE
ChvA7g5wiofaSZEe+TVEAvv097tV/4eBL4ub40UCtF5kf+2kGgleINu1YYcBgHi6
X0oULSNJqpQyzkUqTAM7kKZz9Dxy4PVEeVTb7L2tae2R4Xg3JfoT8aR5F612MWUA
OrxQiSJGXbkM5FB8XgJPfyA9IIiBYr59AZqFBi8NE4C3LEm2/I24sZOZ0KMLP3Sj
tEunxoemMn2FkkDQVnMvx9TaAV4YXpiiET2Du2QNsqYOGYpqU4d7jc6jkjyRn9KO
7Xty82WUlCZswBmy/yGXH73PCHHD5JltrqwmUcgsrT6oggIN61ZTsfXf4RM7w1JC
2HOHwG+vOtQ0LSKoQMJWCAzYSIOMuOkU3X/XXxu8lVt+4HsjEBlAJT0iI2ohnBb5
nB9HF20vZAFMRxD4PEgWZAzq7gcM/Bx+55tYsQMpLfMa5UoC0MJ0YgJleEyDexCC
++qQcrOJGcrYvWnkQ5r0b0X6za6z1ad/op88H22Sn+Jfa6YZZmKuk5gVgX5ueIuB
885BJB3fIk/qjVLai9+CgduKHm1zZ69wAND9Qd7oq4zQrHYT4zdMKs3parv9cTeK
PDXmeIvClLhPpmkazZQ4/8TH0Izpr5vuNFsR9rPB08XJRcgQr2p1Pr8iP7pYL8tZ
rRrW01qDCAf0ULFZ2+XcP2VxJywZFvLRJUT1EJ1fA0bWPPvVuA9iPGaiCW10f/cb
2aKiEOMB5nkpobFm81Nf3PzPwQhlKo5pPV//rwuyI0m1Y67jWJ2KolKKJoqBlRlv
fYMLKvwAvggX/yF3/7ewQkpt71TTOnyV7Xk1Z+sHRR1u9+l2T6IIowuFhKPqNJGj
Ku3BReY/o142yD/UkQDo2iSYWqEcPbbwx2LXbWiIaPnAeUPiZXaOEbhL4SC4xfWj
hfO6iIhjMuoZgffw6/0bfA==
//pragma protect end_data_block
//pragma protect digest_block
WmMgXox2jptO7d3nRJlx4uF/uK0=
//pragma protect end_digest_block
//pragma protect end_protected
