// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
YryLXz3SRjFnuFgU9NaY6dNSiwVd3Xw/MQLfW8LKv0RN94C/pnPrlNUScOtXuEx+
nqZnaSNAKLC8ePHQmk3MCyFEBuAEK8FbpGUnMYpjt+29D6GMs6RS2aFw5nEgKtj5
1pZ4vu63DCZuX9HfijJvpdwkezUwmG98RDHR5UDLRzXH4BMXVogH8Q==
//pragma protect end_key_block
//pragma protect digest_block
1F9PRHmQCbDo50YDj+yNQWDL4Yk=
//pragma protect end_digest_block
//pragma protect data_block
WV8f89l83Qj3kx2YKhQGpHz+y0YMsG2Ni2rpUliO8Guc0dyc4FtfO7ap+G0FK0pU
zbCaTX7mMdF0itfDlWCMW2ZFVqdn7JbxugdaHUrGBSS68EX5iwwKUynHrv2CIN+c
v2bJLUlGxXbF6qODYsXh76xfgog+FobBsmU9950Nv9tDWIE238wUlZRAW4XTqQvp
wpUO2MF/1JWD92mh1mMuSsrGoTcYODZXU+67xGckPJPT/JexANp7FYZBg85Mph5j
wE4m9l1NXK3JiyPjkjDrcId+i7yANv3/xusXyaM6oodIbqTw3Z7I1RfFDau6R4i4
jpa4C0BrO4skf5dS3BCEw8uRQKRl4jMaigwJ3QFBs09sUdEFUTsvyYSad0TscqwB
/D2+CSB3x9S1eCGqusAbLBVhWoCR6Oc/MtvG0ltHQt3ltchk+k0tP2HHXPGIzZKZ
xrnvleuWOx2a0K1kA96gdZXsa6EXZpQScw5DA1fYITXfOW6UtAwqseYvVnHXtKuw
OTemXIeVB+WiF7m/MuDr4k2LU9zdzYVC2uNhj6Dkl7Gl8ybdaLjY6fyL6xNHUqz0
L8ZPpwSHL+e2sT4jC66kd1zEjGXCS5UNEIGjwSvyJn8T7MvcDRyjf9mySreK3IRt
3lto5BAlb/tvUfsi82za+eHobhRLldprJjN7sTYrZfN2rjuSpfgpT302xJ3ONQWl
axfQ4x2nDU/oYNg+aGW6Cwewr696R51KlBa4xzY0900PZ/kddmL9VzKHb/CrKG8x
Kqp1OFZbfjd5fZkzMv+A8fMqcPIAADAc9KJ8q4UiA2fLNmVzhgh6QTwERzGJ3ENz
dIT5sz1iPCymAuyquWc+qIOu/BAt9bSuGJ1VqpbFxpa9w+HYC4BHA8luiiRDJ4U+
NF7QTzo2qRhvzGlpZMMSdN0E4OLYgpXx70MukdNgl+tLdysjw+4SvNRAHPvH2Wia
jmlcqB+HimEPvE5ghPWZRj5X+yPDVAbjnFxfJmivT1YUlRrczm54dNA3eJKHznq5
LtSLZVwYE7KUwaltY17QHkV13XjatNfoB0c0i2GyHydQhl+j42rdg0KJfPgXS4WG
sIZyLfzG1r83PnQW/NfQ2tGHIumnKvFTDisJeWluWLK9yoM2Vbe7bWzYn4lNG04P
tsjwkDx9b8hv+9GsFEPsVkL4MQJ35bw8W7DGcBradleX4Bkgakf08hr3NWQv//CW
rz3oElRCv0sLXWnfPq/ZYQjE3YntyOOF/JNtLFTAaENsaqU2a4GQjuXcHO9gtqPF
WcILBC5xejLw3jcfevu1XGYEfnrHmuUsodCp819HpprrBXZSKTQqLgq6cgAj+D7l
X/pDQbc0i0WtuHPMVEMkeds8sLogFYxqrm876SJ+Yq0V1rc/1za5VjwJm9o93T8/
iTVTlWJPpITbRMZS1tBInHlBy4PMOoUQ812k9GqD2xENszXPc3oztlGyMX+kN9Fq
mH28KjeDH7iUb+Hv9uhmp/icK5JsQ/TdTEmPS9THF0eloeGRxewyq8DTtwq0YHfp
ddWdbawZucBw4e4lZAJOlabX195zIhw5lmGRZYFeQK8ndj85LwwSoJh8DEKs78k3
4FJ9CaFP+t6PQdlmAXbHNywqBzcELTSLmepHrDFlm9Jfgx18FPsmSS2BrjWeBt+j
R9jgqagHav1GDe6TcIYqXS4vgLyKl6h6xO1X/b2/cTH2ZE2jeF3danUasVTiE/Lv
/jk8kv4m45HTyA8Tzugtmkexfbw7B66709lYHsakP9PEwdATbah2naHUPu3TazL6
TGB9v+S0BArj+nO17bjmNT/Mk3qn/RJcsAq9hrkpenWyZe4TC6ZdfEujWNdkal+B
wnvGapSrOevebYgYhknNjC0sBT3CmItWuo5It1gblMOEkR8xPDvzUcJVMdBJ+UVX
Pv/2x5ni7iUi6Iwk9/z5Uxgtoh9OXOltVw0YxcweAz2v3c63EMbOj+YhHWoSb8Vw
QZ2s0BmpQNNZcDk/FE+JWR+njp+PMzoNbZnIg2w5OuJhFwW73lphpX9eE+rwK2XI
TlH6fTCebtvPdbvhLtxTIQObL69E31fLI3NOpzeZtB5HHEd+MG78bCEInautaDys
qzsYWBAn+nzEyMOh6pAAW7KD5xM5Rkrx44o2iz/JoRes3ZJhuG0jrf1sNNSzs98k
LqxzZQYB1KmoHtyHAJQvRj8Or9Giq8nPHj2bCM2CB/thJ7ntj+iWl4/yq6XG14Mm
4w7pqX6/zi3ZGd8nDhGgHwUu3XhekvDsYGLp+P7LmIs38GeucrudirwhwUpiGe55
/O4fV6Vd/OePbTEqRVgEV61Zm2y7GlFa4KL1n3zhJL7xLtmbq6VO2ZVEoBPDX1sx
Cte7qCzlaFL9/kJ5Atq8Q//6r1KBJho0AZGQxBebIcUE/yFNucGW1fRmmE9ri2x0
i38zEyDcZe/w6hZMFxh9I02/dHIt36YhTnsrlXb3cy/x7b3CK0WJ5Gvf8Y+jA6yI
E6JNvLzYArKVivSXnjd9snptc9Z17AGkTLyOObw6s1dNqxVmUono3JGLDMWjrCP1
CLRMz2I1Ox3zyPf7todmfkTsIG49/rNXrsiFkEM+0j1cA0p4d9tOAevsrqu9QXf+
VqHjXj83bCMlKzbMskA+vzeCgPdchNTIqsgpfI5hlKhgMSNUvCwrt1LJucUE8pHt
KWZF6OR5rRh2k9SjWSYCFW1Sw2j2UIK5b7RVDxTj2bI+GhMXRdqlOBELNxyqRV6/
QFsNm9XJ6MLO4JUNKeP6VTcYok6gq2t8CZI2KhkCwVjISX8VtMMisPv97Fcg0WTQ
Q1M8pss985bPXlc9NCxqyIZUVuSa9xEertSTBx76jl/ASEUPXoCwZe0OE0uwqG+s
5OiI7tU49czlC3NWwL84B6xU047XJbQp9l1B+ihP1G1I4an6/1QW+HLm5iqyxFlz
gBa96+aDbwBs5ljU3w45PmEcwh5qTNS6xzW+sj4Wp6vJMD/ntoFpAd9xRsOhP0oD
X1ErkERqeElKj1kMdjfiBjO9SzKKupNIQ8vL7oM746avwlFHhXEni7Xi1lH79Kf2
GaWmoHsgBE5e1PCmCr/CBz/9wRsfIcmKn1nyrdp2uTrDldZkt687V9kgocKnfj/q
iaPIZDk4winTgJfiBveKy5sJKRCRt+s0W+xtP6BX5xwKuofLeTMXJavL0hnEq/gT
9s57jS274rTa5eFFTVzAVbytg6vyiO8PsWkYUNeqjxGxjHSsCtl5KcQIVCcRSWx4
39i3Ks5/sZlHj3tgbsKcnSMqh7BgjnF5FLr+6ihf31d2ZcvTSVAFL3PvwK7v18z2
M2G23ZlwxuQWb5UuXIhB8NqaVayRL22v6X8PGy3OgkmrCLLvG67xWA8NDZpwHYk9
F7+6gWE4tzhI0Y60WsqMlBcooz8hCPpvJYrKNmqX53sZRXx2slSiFYsfSz8mywOr
FhZkDhotGpIhAJ8tRQqKSP7ZIGbEEcNbek9v+lj/lE8aLLpRCWSgtK38HrEV04QJ
cnhgnPIuZ1hBGKmBBSieRdrf1Wpkg3BBckS35zMr86SUWE3KrEoiiMmu/2IgaRNB
FVosCNUZIzZXQDO7xXuTohSMOHgh4Rk2/Mimmep9jBurUiTTke1qxaUFHfw2E4+B
1Y6wbBtrQa7HWDws1SHN6VmGqKXVnLuXWcJGwRwGews2edd4qeqY2ggdehD5PA1Y
TmVPiVM2kBeQtzO2ujGXacgL1sski1A01UAwfqmcSmXLtDc6nPfflJbN5vp+bzoM
aXCvZBp7KGJPdGgMy3hyBh2a+oim3yox8s0R2UWZ3U2rkjT+Upog4F6JavEtoeps
kDn3RsYh41DFkHLulvuw3BSHvN1lpOqqIX+WKG5Jr10VW941n2auF5Hh9vCzIV6j
uMgXYLn1QE+otIh2Gcs3Jtjd2ErhTcb4DbOfCtHZjnZkKHkLhsYEdIjwM35tnPsP
2r68Nww5EUl66F2lFtgqkJ0hHibAYIXytsG5LwYhUjCac0NhZpa6rhG3PRLc3kgX
k2WObxBkHjjnfdNddKFsgbW5y9rebuHBdnNIHVxLclKSrPX5nkLT8qWzTI0yTJzC
fOnZyZgNQOSJ600KCtBoRY3cmHX0/mq/+kQHYVXu2/C+pFny6jM4iePZZkVkucpb
07D5I913xnobadOb3WU7tquF+H2HAiCxoaPnXVF5tpGb8rbxl4qHbpCr8EhE8Cds
v9KA3a+3Rh4jijtXrYD9SNEKb9E9IhIO8tztGRNEP6VMYfclD2VumxoZWWzpVkNU
4a1b+llyi2DB83QLcsTH2WENGnQrnyuXYK+zuQmPJMeWqzPANCeuChd6jrrpfZiE
rr90rQs5hB/f47ijOGGNww7Ky9cqaDNrBjCLjTQsYINRi1Owq5nEGxLEBEmjiqC/
oxBOmPg/AaMmLvXBJIhXg4DdaQXzufaufXTh2Fba1l4bpY1u4MoUKt/oSLa10L6e
anlC6sP0kuxHd34S0JAUOnkPMVgLMqF+Opc+NnN3fDR/MCqsRXwsMkQQvTd10c7A
y4w1eFGnXu/HcaFV/B6hozaE4kVcpEABmtGq/uTxwrO2JtBYJqZBXmeKMGONPs0r
OX+pI7pvdSKuGbtNIyRvL7xHgKaDXG2A6Qy48pAc/OtQXDIYnkuy2zEJn+rRb0pb
mYyuDCnE5kAuUivvPwmoW3vqHEoiq4vST4/ky+C0xEHc4W1Au5+d37GURuO5Qekl
xzsyHV2ywSdvBS7ABORxXKiLDV/S0kxp2AqodzpKZe2eogm3C5FI3tS9unhm5Q28
NxYSD2Yz0689HMwPGBHxNBlUShKR0v6TzULFxMrpHEW9lYYrFGyk5yrIc85WAetQ
O8a8h5RK4m03ew+GABBtoN8ucsc4kAACTlR2OlKp925E0Bctk85gMe6v/584mArk
OTcoX0iMYkuIVLvgvOSqrdhBHdrjoRo+XukaNPYOOyXtxCPgGKw8fK6ONKx/oJr7
BZTFBqtPnX+wsxvyouPETbzijbVGTFsPDMh0fOvsuweHc4toCMB0QWSjVkJrgGNe
PH5V4yvFVre8VRia6H9EK2t4spdSXQj0Dm3oeT2+Qmz2SZAKEkn5mNue0mOIeOvs
iQ9dDzOPOkDc6mx27Vws/DSMb4YFFF5cVpUkOSvoCGzgz2H3o7gU1zjE+TRN6wb3
nwvIoYe6uPTFXhej+NNi9lzCWdM2gLOh+yqYtcONj3M3UkM/9zoY3TGtUNgjlOl7
Vx5uSJo+x2r/ngmeiu2ZOLaA4w2XdtHbMJ2ZIK334TN2krWD/g8KN3ANlx2q2odN
3j7Oafoir5BAaTK5YtAyxP8ouvP8V3AHIPk+InHAe0qDphbsFrtXy4MawlGIgI9L
9+vqF0HxzDWdDzmeL4yIij6yRz50m452Wp1xRTdAl3ozr9scplE8LFF7ItmfQxrR
wRPfzuVx4jNck4ghGp3FGisO4pG9+9tv/dOfQPEMvVHDI3dgK7v/GBTo085YsJbe
AUFq1dc2bZtiaOPLZH1ffTp1EWvd/xd+7JOppbw8N1OmGbKRw6bONAb0e4YLUIWy
rKUsEzAMbK90O4/srJgAD7uwOGYWcM+5YnHrLz5VmX5kStVgI0sABx33MJTnTUTF
94Al5dqsXM1qDaJTuKlY6AHRUaevgidyxLSjNT6WvIV2JaeH3Ttt4GdwsoqvudsS
VoQHhxNcwrTfXeqe4xUnAKz+7u682K9T4F5r23//YWlhofFQn/fE6cuqN3Vzloxw
4U4SyT33f0OyZFCLzb9jb9XN0en8fMXaMrPWkT07BQiIBtO9SDY5890eobWl9vMh
FDxelPsr1lPRXnuvE+JydqxMZWddjR0b94hycG4LprC/pdejy7EYHMx/NZYzj0NI
KCl1qdsclaz4a8iK2pFCz5DMo1SuMAgRPLNTiZGydSDomC67Oop8xOeMtbO93aAi
+vXegRKhP6evbGGYMX4uY/Q12CHCnIXLiF+Jjw46VlSrAldQL/ovQ11lZqUI0y93
Or34gjBbql7pTCQwMML8Y4E6P8xUxxX5vtRpuNxCv7Dj+c4SReFyX6fyUM8sYhfq
boUbAZiNw5gJUIvxYWADDzeW93KSnPPubiiJ6Bk94sBni/5gz73iita1D4Tks990
IaZ/yxveHA12U7B7ULBKjv7O3rEuwLGcmouzE8/CuGk3PmEweUXAYz8moMums9Pz
oidK71RxjnDPbzxBrBM5UPsG78VkvgKZvEgiwj9KH1q/OZ2wiItyYhu+VDUXd9RP
DHMUhsD+mts1lvlrVquDdWGR5KPMwyjA1XMGl0I6R5vqb1ac+Lj9lPuYpOMPIJoQ
EZrl/ilPMMB/0Rmh4t9ypKsweKWriCeGBigPE5enwKLCXXww9TPXDt8CJfLol7CE
jeb4O8h8HABj+c9G9nD6kycd41Vum2CCEX2uHiEQOyhzbF7W/yrCSkntyPQwxLn2
UWgBp0IGNiIyYqeEb4/3YEjcAHAxgmwQ3Mr3Q2H5kioHS00we9nMBY3qSJx++KyZ
IGqjjUxjrOrJnSpjODfdp6O//Ck4jZdfPUiN19xbSGpMKYIbERGQomaAwUWmWbDy
PcqP0sUQNP2DIILjLtAgKsj4xKaYTwF0NH7yDBy8/3sDm7ZLevgu7323VSkIhMiK
Ix86kMl5SbrdVJyEjquZRC3R9Lm9OY5MsX+urjHHWW1MxQ2JOxnZ0T06nGTgfexw
s+B8DOX8LOCW0ksTgp6RiJ9TflSEgm8/hGOKHyZqjmUHuLeC7Al/hylwwqgaFJRC
7E0lZGB8vOihd71OzMb/y84fQLBv4YUhRC4luSRemVTWVMIvqlZhcknfJtAFGpLA
t496bXllWVUgckF+/QD1XRca6365PTRKNelRk6wPD4cAyuLLYoqA5ukVooW2MBhg
sZp/d5w7Nh9SMx0ykwUXRD271D85WKIWc49yTX68F1pokOH4pLKhaoNTT1DZ1Hge
NpeZBkp2hZgAVRYVqay3wnuGjNmJvayveGSjCrCD5HUoUQjTXHW7gZr5MucZ1lMB
2IBZEScYBuquw/aWSnKS8PhjFGQZKuCKLEFGntfGMrFK1Lo5Qvlzdwn/2OHM0f5T
kkuBgP0CB/Pw4wo9zKOgMuKG7Yj9axTBsDBVFIFN5NA7stUx/IL/Etcl/WwdTBwa
jt75kPhxg4JjNI2NPmCijElqaom6fa/lcuJZmkZJvMyTOp8F2WFU3vY0uXuwuJd8
38DDvxK7p2D47pcdd9KnMvBwRnEmKdGJ2MCiMGD98IC89E8daLAkztKpp3gNO4OV
EWhuJL/H4+SoUst/8hTqg9brfb2aOXvkO2xvhFBp0UTW3dXHMw9ewPrAyI0z1S7v
ZzZOEJMh+59Y6Vc5Iq4InYnNqbVx3U5yw7F3XpZc8teYYRTF1ycNifxO+BshOVrJ
32k/HE7zmXQagTgaQS7woU8P0MbuGRniRTjknFKHEDnQQwUwNu1XPrVuUXphF5Jc
sOUaNXiv0CyMeF0vJAot4E+qKgEdKfJvgh2gg6ZLfvYiWd1llhZZoDJ9j4fdxceJ
Bd48dQwXFug6PGqac8YsIyDeLg0Ffoq1iXEyAJvPDSSTN+PtIFGRlGqYJ/m5SBCg
0nhMu5u8KbLY6/7A7jPSoMNHo/F6OOKoG/eqBKCj5CeAvOUN/9mTp0GWBTdcgVeX
c0Da89HFvAjy5lZxDfAIK3QDlTFoA1bDWyYqSkAZ3yCGcDoyhwor0WYxB1XkVjU1
atoM7L1wPNsVjyiDCpDvIImfsvy/jL0ASWw1Mx8zA4OkxjTvMIM3SnHr6hvyd/Gt
xLyGSQMsFC8jkOlE0sUpNpEIl15Eb+KW41VBHLkDL2b1vG2WJNCmKr37Vu+FvXfk
1yNbCRP7CTr9UnvD34Im6kMzeqWvCEqd1kbW4YVrHs71ifh9qRum7faxfmBTcEyD
VEY5CJrga/r58JtIVjfqOL5FxtKjJVCzKODdbsLal27llG2D3X2WJIMyTszBRwUV
fw2SaR9aQldHkEwhFOz/MKbRcak8rlaJbawLZMUC1JOL2CfTpnYiVjdPRt6JYlJa
FVaBV4PSoq93lMdT7j0gIT2vB6O1qBZwJnXl1GgpZ61zbxYJVt4ZGdrV/JlEBT46
Y5oom1D/w1Lw7ZnD9+4uOfKG8Kh8LUb1J/VeAjPz8NLSmPbfYRXnHggRFgZtuL/x
F0ODgvCKatn0nuPVDBI0ok+Q4kGkEzfbh27ipSw32kcnMCFnD6ssDVl93gr59QDR
gw/Ca0QrPYRpvsemt4FNUzuxIdnKMODW8DKb4weI9LsgS0V7GT32i5sGsBVGtoL/
1td66ENeuVrmlUgK1xJqvlIhGK2P4BiYhPTpLm3yLcqiCPqbGRYbQSqKDh5khZ4K
1s+xDjLTRpYUzy0QpOr1/xkpUg25yp4RLFpofc1nqmk/2XCWY5Q97gnS2gk5DwfJ
Xmn/WyBFcgRtgHQHBGE0udYm/ZSKTxMPRJ7SZfvwGk6MNPT1o8mGeyFWDqx3hQs1
+QTFxA5vmHij23aFoxwsKm7XXTGRHT8fn3B+YLGzoeLtqOWnLq5sM6noKiRjCush
Ica7Y2lmuKrH+z/IApXD3adXjA3k1PIyOshfAc6r3C6SRgxL8AGmlgp4fzIIkE70
jcVpHpPMfYhYwcEN12gOkZLTGZsOza4ru3o5xsjbanbJWwkeRgFtHQWrEMPLAm+m
yP95TwW9IqAEKcRYG1RD61Nqh4RmrFx/TMfswvjhrp5BiJfbPMbyKEvYVCDV6y0s
QV75mxEqdrUYETnOSbMEF8XnYPsfrF5smjOjStnd1NNz2FefZY32gRpErS+78poQ
fYeZorWrGV0KnpMaVKUP7+PB81vU9FgDGOF72Q2Le/gnTyfyvBrww++YfvdnZ8un
9bikupw+m3lXl2+PHjLVzwPx6KlYjnERzL/UVDz2haQaJk/2t3n+YUFtKBj899xX
Rb3rw9DWSzi8glftkBxYhSEwqzl5fj7j+XITSrLVg/OEG+5t6HtJqTYMYzKo6SOU
TE93A4YhrF7PeXY6qmlxtO8gnjVt8+YL3Moq5qpS8Wys+iCzVcckOlfdNhY34fDp
Ey+XblvbVbKDiKneZHsBDFg6s1ceNqQEEt2h9RGd3oK8fAMZGL8IwYoGXAlEbidr
9GbK+a3GdHjKUXeuPDVcA+3JOQN+oANdkvnfbrhBnKk1qQ3HHELzxdpgP2TZo8oJ
HXCr82ynULZwN4CcOi03+aBC/snMgBWAmmWSEW2Oajfb7h1vxCvOjs6/pG3EW91C
+y+B52YLQCg3sfU8AYs1B46GTU+p0yJh/+t4ZlQ7VCq+IddZWzni+MM1fGAoHUAM
NyfJY4wmOVlKfWqDz6V651oGnAb/TXj//4LoM8W5hZpQrD1VAsvysOXAzLmhfEXJ
1rE+8XJ3Eb9gRKeS6E9HCl3tNBXLnPmVXEonpAg8PQ1HvSfER0RRVbUPd+D16t99
c1ybefAQgcPGOTinliyI3X6HNvBPTXgZQzfD0YAT3tEKh0GM6k4V5ZJY35Pgd38A
8Sdrej4iXAMuJjDk5ocaDGjxLTNd4XkOcMttPqdenZre9wSwjSVMpiPtQYv9bWCF
6I841DX9cYcO/NkzxX2uBOAzLYcXXmTSpiHBhwxlEvoUtFKVyDcekAuf4BPk62HJ
byxy2OLPqbS6oQyxDdSt+t5TVpfDe5K4ThLthmGq7UcS2AIeVvBXkjEalXi4aa29
kMl9+dEWD1GOUjWEs3jCJnihdPpmBRcYorlsC4+MqUhMdomn8TZc9g+pTYWpxi3v
xqxLCjGNEbA1tKx58aQEdCa7am9Fq3agEMOoD4Ua4KyquAzhlV3RTDGD9dQXBO7e
d7wTfx4XN9ZvwfGD6dd8nlc58wcJtLFz6Yuvtw6/U29eIgam81c6Ub8yAn70RFW7
o7j9AIKS8OmnHxlWdNu7yOV0Czy0NMiARaQyBs/OZrYqK8OGSrz/RALX0VuYylJj
hB7uzyZ/JsAJHT2hpbz8w2tbHjxlCn06l6cn5kKfy7+T3R8PYLSgJtN3TrQi3oj0
dg0FGZ0tTUSZkDZGSC8cYMBmSl/3JCqu0aSxzX0yUhrlaDCX3nYvnOw8M9FGBOBq
RhRj0I0tTYYoq+NnzgFKpeYaI/gmHe2Bkl/s2eRfjW2skw7DHy7vzNH53s09EO5X
FbNALGfdifXcX70m/0LUBjCrbZ0ONCjWUJI1jGPo8yXiJOdanW4TcH65j3jyXs5d
meVSm4Utmf0azUubv0Mq6JdXqlin/EQ2+lBTQU4oTHLsG8dLbTavCdA4sokQn7QP
Q76ervhkjDDjms2voY3L4KBHXFRZ2jhg+uYOq4wTHp31nlNLciN/rz+8d7KwSVC0
lhe2wct6WaxLiTy0p89nBBwP5qRBKjc8sAMww5Q3vTH+EGMLFcAodxzZ3Sg868R2
k8U3kVt0Sg3DJBrbPkU72/RqXWJidF7Xbvd60DskrvzScFPnIDUU/jddNJzmIHUE
vhxC1V/t/8JKtmnP1JZlZm8ldt69sBiKVP+I7J52Qp0hrRmvqGDecLQa+ZgcJK8G
q12RjuEeq9VX4jY0U6UmY9P7KDsfQwJD0fTsAEzqc7MXxgwEq52IW7RDDvlzItMw
TQvTlki0p91NY8AFXH+XitGCOTOPojFsQL2o7bMpv3zDJcctP3LAqlhW/fCy1Xqb
/eUeAue1NZNUm+ZDeVrCSB+jp2wxbNImxofiBvbWKJeY0KUGKJr9yJAc7MpbTlNl
lCKU1AzkQmMBHL/uS/etH7t+GENzRZwm+R32vSRxya5ynnqXn46eMPWX75d9u42u
FrFrhgVoyNodysuP7lZ1mAi2eGfq7Z4CEfwNXA3U7/tT6jUshN/V5rJJLKC/EKgJ
PEO7qikVpeM+02XrLJHbH6H7Bezzla8sULc3MBeEv+H6Xa9OCMoh9a3cbaBmrP99
UvkTii5UbG23AQsAJLiHCZ9nZwYIe96krYpq4eEWe3IBkoJPLLxwB3Zqoa6yh41u
w+T1rrg1veTkX9H0IWjXNf91vkr175Fje4tLqh0cj1mQEo8fJYLcG9yH1qb0/bKn
2joEkym6j6+XmXy3QKvGjRNMLqRk5mBKgxs3TL8PxrooyLXs1MYQDY6bI76QZUc5
l5Xe9TlZT2Ymeuh/QUYNeGQ0fPSAXBcrjmM4zInVMieMwz+xmFCfoVHAynUJCDxT
+A7cJ+0DDOafes/Rk8JboTk/Un5oTJXuSvv2iAAqSHh31X2HVytalUjSKPf9PFK7
zp+eSx2t1EpNngxw1AlcBDg234wYHmhANL/rkRqmj80FL9JxsKfshYyRDmIFVU3x
g20BMBLB+Reh07HgNiS4mfLslRAJ/yc9zhxQpJCMvXb9UHy6PGe2+M5zImP6Xn7W
doWTlCRmeQFChWLJO+5opkkprC9dZ1f+vPcOn19qeQkPEcI47LTpKwzVkPydxk5l
Cm8GeHO2Lrv1a20q0mJtx0PMVmRlyjEObOjQpipgUfJNpX9Hd8hnnNCncOG+gj70
06KbGrhrPWPcrTWV+pB5amc9301icMhCAsuMVPUhE6OCJejII2UXsmbEBLxnEdYu
FrKVF8/7ljnWPRRl53wqYxb0Xzyp8Cx6D0cRDWCEua5VXwBxRgI1+F/GJMwNSZlE
80QtiUoyGd8k7KpAY0cmR6okxYvomv494nudajfE4oXKoKA98nbxmlVAgRr5GUdp
KO3ElDzRegyqpdojWi0th6LrRlCpB3RyL0N508nOYtLjHcxWJbujidX3A24Zq8mK
PAQbS5yrIQl/LZLd/BjZ8xQa3VFe5GAChCY0BuBJjKG+0fl5+CQDSMZdjZkC/E1k
sDpQZnNaIkUaZ8PM902MbJQFz4uRjHhL+X/r1hQ9PZRk249mVSdmqaZHma7BeQWw
g6kEHhMxrlAa9UVnF+qsGcYLkXfEw7WDNhGXt5chtUWPont8RyqmS0Yq2M9oJS/v
sqsPWtd7pwAjZ67ukeN348rJGhuDqiWMJqGPtoldym38Va3QmAmorpSGlTvWclM9
f2oS8dEy5bUDWF3MhMG/bhybm0TATwc9ezHMGH/sJz+6lubn8QZfBMGWwL1Blrq+
DiA2R9vSsb7pfo2FCHyw6gBg2QxEyeoQwl+wA7jNisIfma9W5tPaqbud9kvLxVNt
BuKzMxpJ8dI7KyaUJXP8Q2hiJzbAtTExFXnPHoYZWTSdi7dOaMD8HG/bEnbTyUKx
YaHFywW+pogXbtYtBFNlMo+KoeAxJ71Hq3KiOVZj5l6Ni26Yp0zlqGTpSD4GpOfJ
uyqJWquDyI8Z5nSsM3HFoZSwH0ElIrxBDtyT6XRWvqIZjebZaV4wfuDqoqZOFSt7
r5SXl4jph6M1aBdKFjByfIWflVvJRoD3pmgj9qkQjtqd/UMpJgbc9ajgoIwx1sa8
YGEk8MAZQdvU8aGKwVTRIjfUQiyN0k0NTRXLWIbzp1I1YT1aZtsUFLLUUW7gSmFK
4qOWdXfECeNeGWap9WMK5rgPnDzW+ryYWT169kAgAdI+jKuB+GKVQKZIihwz7CXA
2sNDd8L30wlsoQJkHfa7rCE9FCTah0K4ebaP4bj52pzw2NaCYO1Y2uJlHvCsJImW
25122SK8sNBSmKnSu2EgdDqD4QogQbKxxvOUCbS//agMoRErel+6SYMrxvvvZjow
GHg8OKI6vOYeVyv4KWGy1vnCs0vsTTePwRdyE5SGBBq2T7o0lt2p02IhPQdfPPJP
hzRmRz6m7fTdSIv1PwQXVcmQVjHiMe53uF997dcG2f4wpxRy66eK1LPBFQ2QKSU4
3CtTHqXAN9utpc6GOodgszFmkjjh801DkBCv5U1dodtKX5+Vx9Kmsm+LFZDJfQ/B
xj585LyboK8h3o+glCzWcQvYHz6BjjIdhEgwAlWdh/RVULZD5MphU+KC5p+5SSls
hQF1PAtsWlLVmCb8uHTgDUEDcx1F62xxhTgpFScbDRVXlTIfVg+s3LVDgQwhe/5h
sf0cHLG41aAzulJSzzbD414tb1hiDUmzoofwz1FFhX+YYGgFFvCBMfc662TmpM3h
WMkYTX4gIybgDHUR7q89GudpyJK91lcGsUtqDHdnOQHyl5BdJdB7nde+jbYeObaM
TUZ3M/A2jpBxSCjFaN/l0l/t8EUiFxEOhXnoeoL/1YriIuTHXzhNv+m2pZhVrYeU
p0s3wc2THkmMImIgbdwnH4JD4HHjf+EWmIF3xp5RS18lPOc/u3DKdRrvykvRU00o
mMkwkUwntOYl752VQiGlDdlA2eeWzygyAgVimy6XHF7wDPDkqEF2izonZqM+Cr4I
hccWzJcP1Hshn1nwCNDv/94IMHx68PqpSDpT9jCSpiwWzgDrKRv45dfzBz8G6ZjC
rvpX5WWyaboVehpZK5IWyAch2HBqUJhwX+3o0ZtQFqH2JsAk1N7tdcyeQ9q833X4
ZYm6kl1lrwWuLRbm9ZYx6Y+SytGJ5abqft9OF/fR2/dulJkObY2jxsPxBaiWvkeX
VCumy1zhDtErH982OUXVa2jxHKOcr0bv1klLofvy2OQoZBZrViVuuzJBqoz9HBSO
3NKEOgSsIvqyRArG3OLXCo7l5p1SCbPYK6EARiJbp8bT1/UYgVsAMrd8WJDPa7JT
BrRfcE32Gyu/vLjNbg8Ma4qvFaSJADjyubNNRd+qW5yaXFZuAPfjPmB4Ft9e/FK2
QOHn4wT6qqidPsDJPnkBK6tXzRIFwDXJdtgveguUXHxSCZO4VNfE9LBHjKsJJ9FX
UnjitkCmPmt7e27DlWdIYCZQ3w08IehbfDHgLN23SRxF3LIGQV8+Kp2zkDroSMBu
K/m9J9pftnL4TW12X6SYh9y5/xLqWl9oD5DnvSm553j6x23J2K3j/ExvL2Rxc4jH
uETPUC7cc1GgVtQeh/Xhe2uKu1Ntxd509tLv/0y3BbDThrUr4PG8D0P+RSzLO2On
+Fgbl6XW5BDhcBjUqWiOExpFBzV9GxXSwY5A/dWFrARrfo7Z3D6fpDy48e8TEUxh
c65pOfBSW09Gnp/X3e7CoTIcJEc9gs4E+MzBTN2sU/ukjv18HDM7o6ZVEtyCXSBw
+Vn4isMTj2bl+jaA5XLI3vL0HdJr902Dyc3bJV8xXjk4zXFNXnstJ0eCWKYLYqXu
1Ks3JfsL4EsVNLW6VEVjKjwzz5uon5LmC2UcHVWOCkzvihCyEqqU4wcf/gXXKmV0
EZcYkisG557lpTmqEAdODzP9wJNP6n3ututrABcDpQMp+IRqgaFX1ecDsuy5lcuY
7UnYe/LoGRYegJ++My9YOB3TaaGRU9O8jis+2iBkLN1Nrzt0rJgvHLWFo7JeMSYy
1dyFxs6gjMm/PnkivICcEPjbBy708J/FW/JTJ871N8p9f1idMoqVOF4GqjRgqiMI
KHnIw6XTadoLtGWkxmH8TFjkGQzconVJ1G6CcpKzH89nS2R7pXslChJY2GyWXrGj
MIEKY8x3wwOApjUkwYKUkxgS6VZGjm8H7wBk3tJZKlJVW8hO3nBsdb8YKucHPxQ6
5fwU9JCcB7c/PSxEiApMeschKMsQ3Y1Detdpk20p/tM6BSg42lk+OUEPH78LVW6A
WmKj+MW10aYPwWKm1fQQ7WrtQu/0/ZdRvhfgwsfoFDNDK+fFftbcs9GD0Ifo18Pb
hQ66mxl9bsaIh/PV0PjTHeQANnyRtlX1l7evnETQPy5ZHbLXQexxTyxNX7eyaX8r
L1ZuCl8uUnZOLyoGYkEys99CM9vPJMIrj0G2eWajHtbwhDDU+OXa9ojOJTT3McWE
SHhQKg25dHq9GmLWy0SKYwv3an7g0iilskwQfofHbiph7i725lzzzTVO+2Fanq17
wlXH5g/h3akT5389o5ZgR7fPLy3SZ0phWYvj5MbAM+qM83WBmTDfr8NSaHFxMztQ
QxClteLWrMuTnlfD0kbuv7kZLvHtBwwDtgLYt0hKMVnzHlaYHeevGniEqCDq6d4o
PS6B32lSq+AQWQKBw8oB0+5EtWR4Je0agJmBHPwR/d7NtqjZr6gNmbFaOF7AEpNh
ZjGPELdm/hwZ7D5a7TDFE/CA6fNVenx3xyQ4DMWLXrGMkC5UvDcuFUbQighuq/ZW
kFSLXLjB71+43m/UVKM2LMoYJg6rr7K8v7jhlLWQ6p0xfNyWXir87l319aHPl0Fo
3hhEAtTix/YFJiUC1a8XNlIiijxlji967FQSZe4zW5S0aT85rCk8fIO7E8wKe94I
Ju/DpB7v0HmebYZ5nrgS719enOYtSKp1buuegN3yO5HZbmIykOt9sorBSM3EV50e
ANneX4hg+fQZyFQNIOmT+FfE29/vn4OKLy9mNvLKQFmPNA1Wh3uOI1hm8xfFC4vl
xyEU51GCgKVU6spb0at9uTuknH9su8CGnwtVLucFJQvWmXi0cTzfoFLB9sf39ndo
+WspPbfcMOT0ZADx4x+xlX6mPvvHXkmMlPgZqdDDn/vgPMgUNUpBUZgeRRTxodZ+
fEPcx9tBQvrNZ9n9oVhzXBq2xfRXoPclRgcGEA10DRHLPc8iFQ8/Iv04pbHeTCMI
/7qucL1+noWeOYAAlD3uzjNKRFm4IX8NHtIqeKd3vMmWxjETCbOHlgvVzQFqeA73
vB3C2XIEB1KnToxD9uWkDZvEmvjkqHHa5jN9RVYKcVdzmejjotpYv39HJQWe6U0e
cBQL/r01PjSBfPayAutS5EOe0rF9W1BhctR3IsW1E+jwbsn5SAOi4UAoOjxKvp/b
fTTieKPOyoEGRR3sM/9T9so2UGLHrx1WKFtyHGUOUT1NhpkotpuwZ2rxOi1C5IkV
/ZBr+WBU9eZrIWihVyUqVxds5EU+iCBokIZQ069XNdCoaChhuJ9+ZyNIhkTBzGWA
vgaJ98wD4Z1EKuUI72XZp03XKHYv1i55FUMcieyqzDvEourBSCDBABwJ8vmT/KsL
FuK1oWyc8myt/3PWVgTQQ3g0EJHBRat5Fhx5eRkbqVTYuhcthvypHjaLsjqOT3MR
ER50dvWichlXbhDb33PipmJugnKD/Cps7bcPQB69LvAf3XmX/Z31obD/D3S2mIpW
IMGy9GZjh5RClB0EMfXq5iBCeTfazWZ9uJxihnyZUoPmGWJWuqn6whb5xIdb4x7Z
mKnsvtikcT+494f9+03ogkwy0q3Kt/UA25YjA50ToSv0HFf6pHA+OL/xfrEb9kOx
FusMoF4+DKNhp0ArmtbpzA3UpSYX4HCFzxxUVnYr1f1eu7O5O1pXa5OPrrG4UMr9
fAwkVvOLacEYrpbL2VrUIxljX+/1w12ngYs3nWqqTD2bPUo9VoUblarHWJ2lbHB7
d/ZJCI3VDG0P11xzjWkBVeyRJfLXc/x1VfhGGgT/AiH7xaT3XIHeKjldJrdZ7QYF
1uapgAWcnk39txZPF1H41plgsoVrnzYUHeMRdFFqgzkJsamZbO6dqZrXWEML0Gjq
WsFPDHylQi0hzCVtbfB6/V3eZADoPLj5n4DQzpG9bUWOks6aAI/QNyahiiI+Bu9F
QVrTPQHVQtRqNYEMdKpecb4fiDbJ7Cvttt7pJgZHiVMgEj3OhWMn/S841DA0gMrI
eOcTPiC9hFgsyQNDHG8g65LHiJOVqxaANAsWi200uS0J2E+F5jttfiprpfdI/PnH
0TVrjJ2uhnEA64XxBlK2av6ncdl2dYTbWGGX9FqYAYGX7WbPRANn/JQ5eCbywlOF
zO2wG/XPewOheb983nkhbsGgGXGCBLOLX6e42t82tpybDh5iTbjvTNh7a0ZfnTUP
2YfQQwjtiVnsuvktozDTgzAafK1Wfznyt2tXwZ1waAtj8KLag0vvqUNsIomSzgh2
RK+Fic1xfYTbeDkpHatoLdJy6rzasV3C16+tGFZY50jypyD6X6f28UCJ/JlgMMjo
C0t4utIalGa1ZkpyNUyWKz7lOWqo9M+11Vhg+vTzXRvSqVvXsJIPzpmWXfcCpUOu
H3fx+Hs9vN7jNyDvdglHnd/nFDnB0k2GKOtjpeN5lFRpr7jsSd8Pdfl9ntV+3i+P
SAjXwPHxZV1E0zyGKQuu8oZjkKjmh55mKnnFx+iXDIuyAA0DnFBLzJ3JpCsPVjsV
wVZSBxRbX9TlhYqAdaFIr9f0CLLvX6gK5MTtG86lMMO3FGHdkjJIkspwP/WXOCD+
MR+gHvxMmkHWCQLQssf6Na+A4By+8NmUqibcVWjWohsNpEkjz6Povcj3U0w6XGtL
ABqHB9SjhFS6mfa9WG7Hd0+0l+WkGDYC2Ke5dUXI1+NEkYiPbgGC45e4TaKzRWDS
z258erwwfcdSKbMXhquJAX83rcK+UT7XqUGSWtDY+Bgq16Qc1UrPWTG510y27WWy
/LONiLjvG4paEhee40shqWujicYgwFvpGwVGmFUWWXVMaLVEqMsMiE9B5wV6JAlb
l9b7z//g6fijppCC/9tzoPapNlJ27HpOt+vfXI0Kmi+2q4aviM3eR/5gRFgKrW/M
Td6ln+iCxqvpy2pycyxf1xF2iA1/j2hRg65flYt7AGJsqWnUNwVco6dZgBgHymS+
7YslMArtsf/TLqC8zvTIGNQQnqkkmphaQFJg3InDL7RjPlfexzGplAlo/hC5vP5o
QcX+SKp3yPrEa2SYsc1P+BlAl2Z4gjZXfX4Qy+RnXjnR2kByxQFGoIcG6UXXQ20w
wFJSB1ToVi2aZZ6ZUKbT5D3k8iiCR6PbvhqVHPMFkSScQX9IBXvjnhpjXq6dEyM3
LlbyqdsXvRBXPg5XTAJvnSSr1yZ3+nao8DdsJ4eI1vsnzVR6WCvhmijgzckoSV8O
W+tNzcuW8JSCMvpUwDwn+luOlqcyJFbgpMVo2MRhp+nZF8qw6E/VUxMEbZndhuZU
4qlC77x/gBI9CyFMSVL6SjMFjTe0YWmJa0xVREBheAhLcHSuq/8qxtSDlzcuAcaO
zsUrlCjnPKLp7jPbsQ85uMJIJLZkZCUwv+tFXpw97bY4JbQvXA/5XXcWDS34ZgoR
2C09kz6+v2UGRp+r7iZV2GHYvFQPnDCdDYN/Rn+bGlAMvzJRovBPY/TFFzrMcqK0
87yGj3HDi5VK7U8EI76RKuT6hO4ijplx8f3G0PQ1vmozBKVAe95m0RY/ktXZPyS7
K/jOrzC1TJ+fYVhe+94YJMT/uFYT9oNl91BgJPn3biLvRB0NXtT2Yutrnwhaxmnr
KOpuhmJKvQDqpQvPw1g24gp3546qlLhfpbXMkfys2XKOtT/LtPBqu0eaJWRrmRNE
jA3vCnnkfXEp2fdvGrT9OtBz6pwSc1cFLHfq3j67e7Kgh7B14Rx53riP81kkhABt
OYDTRa8UTns2x3mbF+tP/nt6p5NXiK1a622r8V+3WuvUyz83CwyfotRVXDqTnHlS
g1ykz4RikOU12jQ2Q7uAFi7V80mn/fjFYU/Ae86phuFp8shD3Az8DmN8e0IeVmQm
K5UrGMQWvRD6r4bW2KpxGx9Tt1zWWw+5VlZDNVF3qbzY9Am0X8XCDrZZSR4pMSot
SkXJHKvMEOXL/GjtcJb+2T61fYW5ib597fD24y6XExTGu+5G3tZiNf6onhuJu5jv
CZTIRU8Io07e5WWu49HX3RavFsKQe10xuR+8hV3msD7+nayxyalXAvbGnhwZerFV
yzzfujXRZtPk35POqn4Jiu2+GX9aV8s9M7KjEpzOE1dmRkEmF77JSR/QMTnC1CPH
tJ1tHUdA/JVwtRbOaDavQpDRi+8mc6c11vtbunMqDhkMi1DSS1UXAWcCsT1YV+eF
JhY7OBW84KvklZAk7MAzqOuBtPoZjO4PtnIMcr6NpXlss+S7IG2bVctdMGCmXcgv
1mJdszYbumWbZ6zUyeUWzlQnDD6HhvKJ0wuYsIdsh/RODq9f7yUN3rnCF13G9Q1/
SFcsL8XGPKa2Bit65ztrwvWo6UkxV6lCYCCwB1zvXfyjh341TQQX9aB3DQor+/SK
9c6iFbDtj/itsGQ4X8K9bu0LpFvcJbQIOUcRJBlv2HTKaOslHtPTiY5b/USCbYOA
yLuXFTsS8EZ9gtxE5+FkE1vhLJdeLQLsfUN1oKApGBY/9hOsh/ytZdaJ6eIWS7Yd
Ion1ggjo/eyMYtd/sU9EmD6iJCpu7TXvWGXe4DddAIXUPtVSroOvU71BNVZWtsPP
S6Qm2xCDiZObyWYJqVSegzqLsGRhu2Q/mE2L0FDULLzQoWZEDeKDjWRPp4R6To2r
q23nzUqPNCuPScRtQb9Td+0e9Bu+my+4/G1yAz3hzgHRTkP61nhXuFVaJAUzHiX2
d1viOS4qPG8ttMVQB2Tey38SiBrcPvNC6I5mUVoiKnc+HcuOJfooIQvNJM1fmBU+
OOwLlR3sruqBjfpsVv5lRMHi/d/Sd6wcnZJkg0/VBUtjbetPCOutLJnazTvY/1Tn
wruRPtUhxHddUcwisDsJJ9vPzvhopsGizi+AZSCAmNvJ+dhuGEhzHo5MqSivool/
v1+x3KuDsQxvGIFgNyluQkDZz29GrSY2mUZXbQ6/4aLmI8PIxbqAecxiibqiUVND
KNn4FOb+CXsC4RAM/OBB35LJrff5gWM1US5mM05Pw0QDU1KChm3D/RKkCWqwSU/l
9VtUtDdPuddxsjByqwXCyHiyFmzAEF6bXuGtxsR9aSizGevzdX2wb9ESXtFqik5W
6JJhsg/P6DVVy7x0/oCjpoctILaHDOQbKoziF9uJ67wmQosgrRv75a9hdWk9Ag5l
LHG1+0uDUMCCpCy8jK51JifBob/brgsGzCtBejR4OGVGha5OTp3NDM+3TQLfZZ4e
3mdbCKuS/TdIYKHD34feBI79xloMRCCZhf49/Sd/+VnoadouROLHxqh9W8hbBSea
qR7E7izFgjX3ba0xeaF88iLlZ/6EfMdslI6H+M1EgAZixKemPeytLiK6n/PVvqh5
M1DkJKnilgoIkR6dGKZ2H9D8VWnAPkRmD18oIMPv0WsDU8TbxH+ucnoGep82AX9I
FpznpSDFGmiPB1lypeO1KdRX0TQm8ZWE+ynaiDrggILKai0pMGSP2bsZBG0UPEEB
JqfC6uYhw3ZTxMoDQPY/SbPPCVdwZYvUb1Asi/emJpyLOtyvhO9DaXVS1hgWyme9
jU23ay+2sBG3VarMrUbNQaM8W8mjipg6M/H0mw4PVUgeQZJKIoY7pv6BEYQNmbRV
S0QcWarXQi26pbWfb9wztQ6HWUWAbEWxy92r7I/hjMv1L/B8qHMoH/4a2ispQTRr
OwkHOcvBF4cXO7HDPcFgEPcLcSYeXozsT9FqWjBFG46b2OSV9WY6YJFWQAk2qonC
U9KofRMDqp1XUvi0BvS0shxbwqQnrMGNDwhoAJiFkuFbY/P7vUo2qsf+T0fSpAxr
mmNQqU6pBPE/E+Vhodm6CPAUL02Qa/0oXHrD49TsIOXHhPu2Nbl5vG+SGwM2KJ0D
hRVacJ73VZBLJIjIVoXfOR5PDFrrxubp6EkcySy+6X7qJ2lMSzT3WMUKMw6BAoqO
VKgt9NC/Lb9vQ6MP0vFRc1sZ87YiARRtNRJAkuGcn8aWHFi2p4owTWIOrF/spNqy
qw6FjHw24QPLEZboKfhSCDshZsUnIYWGiZm2w9cK8jndSvpyRF2mz4zPRt7/X6lI
9OqgcsRG5y/OsqLf9FT6n9xHPN+mKiwQ/HuSIRgZSMukvz05gq0yiPV1vJNUWOvQ
4GwM9wnzptDku54+iRUucTXyDt+VNXZSXHLwlFN4uLQ8Xkh1cgdhzEMGtjwcyTy1
JfanbMjwPQIPeucBrGbuzpK2bS3CNhYKa7Jbd8741SVBiuWulS85kl2qzq9paz3I
aq/wsukBHmFW2oLtipQ/WuSgZBMUtdcow5ZfhK7XczjHs+nVFqaSm36DQhb/Ahap
Lame7RTWRP+ARL3qpua7RXGu3Ljc4BGCdLIjPvDD4i3BG6BxndbG3LyNOhxVmN9h
a18oD6KPbdKKlWKNuXGZzCL6b7MaHKaXd6NLVIZtmIrVVw+38GsOF/HNi6UwabGv
t1nOcUpeMB9dZy0GhxRAF4zRpNqzSrZ1Nl2c8vLu0qEVmNqF45nFnKkyg9MSJR/R
MrunW9n3JWrsx2Ki01AYxILvi0He/n6vMwHAgaUzPnGxIpcBSiqsF3oJq2AKveH2
wiq10ROQrWSjzzdlH9VJiAZBnsW6vj9hzJpqDEfVCy2fJCWBMUvNDMA9wAfxJB1e
DxX5r7InmPyGghXtbEcDl6REHLkPNv/a5hITXSmTKnNK026lU90wWemdnkCpY7Hk
DSJe8gSXJ6x5XI+EB5++eEY/Mlv/Cf1WCPsz6wUcpQCzTUIFahwRauQJwafwqgvX
Z1u50KOx7S3CaVwq9nCVWRQrTRjc8hrDa6+q3Z7MTXrRjeT1BpQTW9+GXYKIujW4
SaZel46dNZrXJKh91MFIQXpInynmA+9iW4JOsnm/k2dq/K+wA0bJlOECAQP4ZTKE
eeVD1J+Pw/A1RK9c3sSefKcDe4QRH+DtoSGoxmJHoNfvFNvd0lmCHkQTgc9T1WUo
t2ziLhjp7jLcRVJL8Mmt1+g4wIc6/OqH2Z3OKGZYi5x5FPTceWUnuWPNa6tGQsPp
DTtDFB4fWrJ+pAw0XUC9VLxp5etzFRCKC/ioxMmH5eDJXHjFuaKzm70H2KT7zmsR
YNXwYcZcyxtFnbzSTDzXka7GkIN2CoceRmzmAB9k5RimiAL+nlF5khe0llZ2MDv8
AHBB/0QseGEggt3QzyePkuZQVaFLMp0RQG43QVPgahNzzdwB1/1qhxfkN0BGQw0u
FVSV8GGHGKI4sl/MogxEeFzavGnq1AT/Qy6/a+WfZIUG32AmBIYnYMyhYKx25Tbp
4vrbrPRmPysumgMYfWQM0EPbOXlgFWcV4pTk8OSQIRvZ3Yvf25Yzl/NBGV4Z8ac5
qmJ0THo0YcU8PZ20DgN1tjz2h0eDifgeYr4sOWBv3IOotB1AJOM+apZ2jz78Ttki
Tn/tPLaOOt4i1vMMLxUMsgJGa3HUXFaFZX10xtmrWT6xeMPLhgYDEk4pFumttBs4
2ZWJBkM0BNdSxEnlO+8JpwEai8kI5OIaaIyZzT9sbLMsWhRBjyRE/fhB4b87+DNe
UfmLwiyHoj4jP5LtHs2F4gxXbjHIvpRKVpM99Mgf5hM1kGbCENAXn+2rmtYuCXWO
O7f0mncT71eMJarqhka0+xey/OuPVPlfFiPUpXcT1H5T8kGblmL2qYjIxDIZoVac
FwsQHaGOUVNf5EmDVhJQeXZpwXUE9b40cZ4Ybl6C9G6hY2fudcueju54gEzO8SzD
VLtuC5mOnorT7X37ZbCshDXJuMBznHpG3VSL5/br3+BupATFL7ZOwHL9HVjtS+AJ
dmuHu/Shz0s7ETkJUGh4foDTgA+UtS5RIUTfRbNw4RNGtElPEQkkshNYKy30RsQC
YCZmDXirJ4wpwYqbEfmd7hLbpfROi7p/INfq5IUQ+GzRlyXSZs6xa1biF3acBTX2
yKSiV7om6TbTuoRmCB1GyxughxHQmzym+SkIjaAzo5jxI0+hHUp6lMziYxTBNdR+
1v4atk/nnjUKaacGgGhmQnMe8ma2YhvPB/1PVNp9iixw99MEz6JvKdA9GJygsBt6
mqM/6VGBFdqIHyvYAdxEG54jszOoe+rt52dyvFLCIRi4pRr9gLBY+3juM/D9wgLx
Op91eVJNBud/qNUjlgKKjCxSbJH7M3CsIiA98WmCf6mMSFmiJ3IQ1wvUSmHK5VLy
7N9fc3e2UvQpd1PwvaAPu3Ddp1M/Ww496H/IN/lDP5RBHa2KCAcF1NqQB4FrPDtM
0rb34lFWcwAe8yi2GD1BLpDwf9HpUPK1cNgpL6DphViyU+MqBdYWl4lFjJbv6pRt
2so5ocoirLXzDqAefFdQPVIUybfRo6yGgjMhFS57a595yKaTco+q6dI4epxEr7NY
MQzqmyT2XdCt+TDLetc8zvTsZf5uQO4Vnhk+1edYLQKvkFESQcsUJU0etHRu0srj
Ig5DLDYrxQl8GEApfNtXq+fQLS/CVrkzdQz5DNqzaTjOGg2LM9vYNEWKtk/dgm2z
9F38JVZWgxJ7E9zKVUMxfW2xz7DPc+xyUwZJC5PHhyUH3VWZmOPSYB73Ge0ZruKE
JQeWSf6dCpV1zZ9YapFOckROm+IufLZTiQAcZADpwQFVOxAGwMoXqxm6JCAZcQ9U
YxZNDjiseGYz/vXkXtnEKOdnbXmtML5zeTgllTIXMR+Gvkpds65hcT5XHso14ygk
kNL+KEomBr9pF2E8F7lMt8JCA6+aAa/TnPCY9vVxqP7NThk1cKJzRzOpTVaYliQp
oOHGMWd2kychZsPiMyJyVXq+jyVxXP7Myd5Q8YuG9wwIisDePJSyud6vlys8YNmw
DaLcZRil1ZzLdRmHDRvC/kgUUx4Rx+fBxaBQrFmMjLAhoMDE6e8ZdLFFa5VlkQTl
zCsE7dAG7RVuLA7517eJ+AtQe0FP8Lou/TkxmKzL4qt3Un+Brb80dWzr/MQx6HfK
SNHwSO7Yls/efkCcQcBdZlZAPO0G18LH9CO+Ih7gFKakzedZ22aMQ776b01NthOt
YD6XZ+TQJJFMc+1Xg8vflU2MKQmLRrhT06t5SW9EkKQJzP24PRsUfhc3Y02MsY3P
9URkhgiYzzgymwU/G800/ySCsBxTwXc2+J/yyG4iHAm8f60+17yHFBnIIEtZGBjE
RJuasmTNy+aDcpTglpIH4b/JjPboCwIKyUDpV6G6nOrgwZ50hbOpbpN82n4sOfX3
BUjMnk9FrCdnLqqGuvyoaUVj9UzcGLXPoh33TJIh7cM9ermzg8WeKN+fx9oC/1tx
1lQLvc/WEZmGujpPZB9U3zyKxYym7WQYyPievYuYjwcy5xcQZ2+gLlCmu4tx6VsI
1NAORTZX+77QgiqnxBdWrNHFxstsPiAS/mil7sWav+2yudzFZhHBXAsJeiSLCpL4
OAm1SBeGXc8wHWICWDK7BbmrcNeL6t1TtPQlaRX/cNCeUgqF3lcq8186qQiswHLj
ir7poiEpa3S/VvNRhLZ2876srHnKRv5hwggTqVFBgH7EYIJBIJ3ROSbsZIYs8eP5
YuL7LYm4iFA98WWPby88UwsYlxDFOMDTnckKd4RbST+Lztd+1JGbb9xYTVNL8a2s
fL28xE04vGDAPjTnt9uCyEOkmj6wtZy4GLWvfXd/ChCrF0umHn2bVGHgQvtDBVKp
KxYo9ilTtYAKVOp+ToYpXeELo+0HX76XDfl2Sf4h2m8uS0qCU027Wjo72Zcy6BDr
rz4DBU/QxBE3l1mgvbPjrtpspWh4K7lXElbucIPPQFJygGpvaTbHRpgGaOV6oz9H
LXHSRQkDIo0V1Za6hup/GoJKMUgdqFSOi5G/8D/5+FBNlxFEU2m2F/IzG5ySXcXp
/qHq7pllWmouKqij91sX6cjCA+TMKReYw4RNhzR7y2H8npY+hpWjlKvZtDJE83Y9
Y+/hTFGQXBXCi1h6IjUV7+rupHK/N4ow97cbNnCgW5PkXBCtt1iKiHr38Ocg9B4G
d0E/LljG3l/egzn4A41NbwpdbI11cP6r2VqaY65nLaJhpG2gZrNCNwzmohqPZWS5
+4yRTkVv7Twc0LAjpjnrFYFzAZyKDjs9VgdUSbeeEhEOdyfPFQsVYdwuuvMtyDL5
qpOclCY96keM3SeW/3tMwQR/ipm1yRIeaWpDzQFK7i2TmW/W51I3OF4FTlcJd6kf
iDiPuu8HaBrrz6chcVdsYp84bQPx90ADoljgalyM5pdynR69icsN3PoZK9FzCuyT
UcvaAAX5qQFMYE0L0iDDQuEpcDsLLh/pWgx59gNQtNK1yqhwuecHVFDshmxvjHfD
noC7p4raT9PD0WeWd24SKhmJmVoo3DYO7enwBv4ItuxZUwlYetT9yA4WmG+zBmpz
kqy7ql6CWcKG0sMw8I0mWcSib2lOVVAT8Fbosy6SW2oPt23WOGovDCpTgWuFkKEv
lG4y0NrraB6oZGEmTH+IVyaQdW+36n696IWkGZi1De0E9H6SnxNqQkIrm5LnhdT5
FYhenR4hkGEF6U7eRXV+utbQEO+n2ktb4P9Yq3lCxqdWR7bh/aPr2BZXpLpMTeos
/M4Kdqe6fMGh5XW/UUZyvJQWzwSTdZ5F09aWdluey9956Zbs9yEwuc5tvDMPEEQF
WG0LBL4K/tlGALnPmfMmK6jlYXkNBnOqJSb1APeU2yxDmgM9hvh7mkkHNLesHwhS
SVRtKBX2Kgna4sE5MtBdozRUpa5Hy0VcqcyV9fdcEVlduH2HDR5CL8D3sovgeHlX
db71Y+L8PUFPKf6eWQgcopbR5sena/V7Ly/U16uhhDaqGVVf0V5CwMgOuSExy6M6
b1eln5xlUKUxnXFwWKJxirSDEwu3DOGHgu7i1GkBb3TrRwlVJE2O+kOwI/A8CM+f
hgsaRgfVrSobdx6YXz7eDw8EfLyWQ0yy1LIyOzrVNyl3Pgdxl/oKXfcbkD8Kkn0T
gxWeX8R1orJgn5mfA2ITrIMl/H2pSNPGvutxh0Gj9zsbUQi1dpfd2MBk9uMNivYf
Rc++qxT/f14OnpN7o+x5hx4Uk1b3zE/6VboPE+AD40JcrIOZqoefO24zoDbNNs6K
v2TugOwxRJf3PpximIkpGarXKskN806U8HPfQaD8KORb50VYk39cxD3kRHuj2rIh
F/HC1cUsLEH027uE78VVaqsbmmVTC5JXHprKFTxCyZ+9vegtuHKJI2VlHqBLzeSR
90UZmAmBgkWQbBiLVR/hA3I8gKtRWuaOb3+lQqYt2DyVCfS7lDaKsy39rSLB8fqf
l9UpejU1IMrFCD4OK9JOxxOUOnETZrYR+eO8lTf6DXo3BpOdZFGZW6YYHgO0LRyx
6dILJtm7DKeAR28u/Yz866u9X9ANcFzZwQaiIvReqmyUzsBVTUOHmkKHE6sipKJG
7dxBKKn5wzYyPL6p7aMb8vBP/XD8IBGEkhrLkg+AoMzgqZOmf5HciFzdGRpAiagH
ItHOdt8qa82SA0fH3tddpQ+xv/tKHvWALgrhf2dB8WmfLBeRLxQ7hrZznjjnwHqQ
Ud1MSvocrIO/9ltJ+1etGT7FrwF4J6v3zVAbuVqdv/GDiqG05EEPdk+bBexGLxHN
zUGktqnYgqkTZ3Pw10KdDmhpg99DvdVanOixViZ3HemMoM4ohep1iBMFcl/qht4g
E1N85Nt9YlJSOLlc6WOto+FDGnhxfTuMqZD6nfcR2CgXDxK0WGSM17AKdF9z+fLb
dp1yKYf9Yq7p+3EIlqcDkO+fYCTkBOkVcHd46X+oycrb3H4e6qp3xs3b6IBw5blB
M6JFwae8a8XRCmaKNrE4ZLC+qgF95s+PXV1BbD/ANcOn9XdCWvAjPn/PGXse0QPg
eZHuPjh3tvaKdmiFLHZYJbHztplskiyVlmWGPnh+kBZi7y8PfqZJw6K0LSPfEb5B
q1mxqRuXB5r0WNXSBDvMi1A4zIJdkm+Ag25JMHMARJqPYI1Xq1Llcr6K5PR2Smn2
w5xiQXGMkE/v9EKRNyAQq53FrKYCCDqELG5QwbDrmXN5OouENfe3GkGL6RYuyfut
HUWqILUzgesc+Byw1gljK+aa8wnF4LYcpnkmpkrzUOciS9kwofjdUFpSxgxNMvle
8bMbAHca99W61HH/aGsgKMRwwLADhYbc5eTrYk1q3CHFTS65x5zy5JlpxVklR3J4
d4CktM2FJWYfAdv/TYSRT0gnSdYWFlHfFfHSfAXSyhyfaTI+BoY13eHVvMr/OMpz
wRpXcm4H5b96gKtU0py1/64h9W54WaMLuOV1YlHbiQErKGtSlpaoo3ADQ7Z/m62H
xMIeBQhNXoXwMkY60YeEvDiMp8dnRJb8H9zJvvGKF/fKqyr+1L3tMtM95U2x4gtm
jRjj4EUE4lvjSM+LeTosB5mHQAC0HIrJ1rjuuy09XdV343JizjvYaPvspRDVTBGt
jmBAzhBAnXKu48M5pDQQ86nBulfhDltnXG/UwIvW9ujcEnP3DscbCR8ek4h8MeXw
preaM5k3y+mKizZcvLRz0QdJpLqr4v6COce9Ca8/4s9zqKJjEjRooRtnELTxMHBT
PcLn+V4erF0cV6sidjDaUoI/RnWGENjn4NWnP6rqE6uR5+xgA7eAxmXI9+pe82Ox
7yxGbaSuMRY7JSI0oaYwXvBXSH3s81vgn1qy295jKoYcM4EnLrauoheYbiekXdGG
VAzme4ezNFCTEa39TcS2z98qvWeMcpkCBEpZvZktA6LaJNHVYWD+5fCaD0wcYAsL
cY0gAJef8/2N+OqW0OjJ2Uq1Qib39i+ILAmchXjuklboxrMB239+Dzfcw1snh30b
Qku6hJuwPGLS2WHIOIZxc8PRhlMaDWV2nEl7bAe/mn1e7cTfesnUlbZG6+Kn+gvT
VqZ3rB7Sr487rrBIwQgASP3hF+MdyZExS42Omz2pRosHWeB7s5sjUNWvYl8oATGd
qlhdLIZlcQnK1RzpK0aK6Q+TBf9mGbvW0aBsl39SUjKXcoSKkaimzroJ77KmvceX
7VXgyR3nu7J0rF9ULl7ahfBPJIGSP0dk+RPG2WlPoOF0FCTdICXZJojGEzkTK9G0
PhMg3j75HyL911vDFGtldVq1pVSv6L3YGRljvfg/0ydcxtHYqrxusSjBddSc9jGM
6faZfQMXE1e7ugG5+B1tyzN+y8INMwyoXGCreqydSOqpFTexrLIkPSwfR0cVT023
2MBIDrOCuqP+vBj9uUTyfetRAlFnPU1eyhoEaMCBm4oj+u+PnqG/FgFLE87e9c6R
bFYFtAlT5ZRGERgNSXGUrHVOBlc/eVn689IQthTyTqxknwCKd0ZQFrWbWWiLd8dp
cJCGvt5e4QWWNOCIQLbGQvhcsr1GiNATcs77ArsfRBLfc77zsL7YuU1kig0JUYMn
xlJbv66YPJuGzYnGgF3pcl5vG8+WFSxVxtV0c34ZmeK1SSDWTM/4IU0g/KeJihW/
Cz9MRRBbGhFuhfAQZVep4Sf4XpG53N19QxwGhm8ExdoaBnnX/+oPhSoKrSGya6g9
tqpLp1fo0K5zCtZHDgF5ooSCuy/rJCEI6lXLHzqLkZmc/ogx07ZFpLUyUV2ki1pC
EM3ayK/Vd0qIhHKUBURF0ec/aaOr80iSwSXGnrrop633iSrDnqXxJvWvTa9ZoZb9
BUFy3BAciECijwvF4O0yj2MR/NSQgV4fP2JoQhhd0qJOFmtKTKz7DZypo/9qMjzr
3hJsUQmaqsv1/YUOIwovx27fN++ZWj0v4WHYB+VlEoFkoTafjEmoWZkReTUs6Bjg
XBXWP2yDDjR73vv5dsxAbxKVjOsBDbb/5bGoyB4tvXlfuubsmWzTc4vkNnTAAscY
DTgxpfF9EZqhwQ28ogRilC0Ptm753O3oedif+zLtOz2lKomTehJ8ahKpqzj5eTCR
E4PyxiuAStZpQU4lUFtUkleA+x5/F9n61FvjTwd99hJnwGS19P5E00XscnZMb1yJ
6S8w9ok1Ij5tc17U3ffm6BvKxxkNGtUUPdL+XrLVDYnWI0HsgJ4flVb2aHbk1wL9
9sSxFP3FbcpcfJIAvHJzp2X/e39+roc0cWodYO6XSreh+NqfoIhjcs6rgKH8F26Q
xen0KgXVuwhiUVOK5JJEidqdJ8QusuvUkEaJ8SXeqrftxuL1LMLG5N2EZq+IjFQo
YzFtrpg9vXIcfbRy4oy6pP2z4tg68UAV+V91GxEWftueUzHtJAWtNMtt6mRdYbxD
jptL6gBa3H/p7FXTRYoPrH3TwAqsQnKo6s/Eq8TkBlSFsXIn36+kkia8LwgVBvUo
S7r7Nfl2av/XkwJ7XDXrdKNtNwOgy9XM8y4OXYX3uHQMCrB/OAtSzj66NmNXGVR0
Kiwsn3dnSdWYovjebvyFJmqPEx2hJ4mGADDZDy1KIXE0FXzb2K0z+GMmbfjlaxDN
RY9wO/zyii/HOzPrSK7/82asvDkEDFbNjM8zn870gB06lJ03lrGd5i67Td/61B1I
t+TGAOBVW83imQBeQq7lDTyME5P0Ok/h1s5/0CNX0MH3M/RWsj5ZcwJn9ETFpESS
Nz4CgG9t+aFCN3+hL+QimMm50du05Xc7fpABbMOzSUas7iF8OsIpEbic07zs7MjI
KG5SE/Rptwq4DMTuiIJEdcf4p1Goe44tZqrha4ikGC9coSfeofOpBLiTHOhdiTo9
T+pyRvQYjgXAJN/ykC7p07fZbraWgdesCaqs4kyO+gxMveSDILCZzDgvcydXpfTw
b+as3lfC8lb5ZaDAxh3fButwcqUOG0jc10if8mNGZZ7hNVI3G5SiJMpM4iXr+EOv
TsD6116If2wOm630CcH3Te7T8qsnc21w/wYLqlAGzyxgaHb6Q5n6oej0l4REmONR
gE2QuUohy7NfiDqT+lYlwZO2rMWG0kY+DrLzeaeKQhnlGwOaBPc+6kohWkT3tBPL
6dsGCYp1a9yzCSTJkYsqhi7/GTzVZsGZrafBePcAchwJzU+cmuana17dTAtTKyrz
t6nmFkxFUGusVtnGEarCwLoa0D2zeUZ2/Pp4+IIwzHVETtVqczzaUqOEIpUHYu4G
EWxdgP+fAxF97jK13d/USCU9TCA4UhOCa4OmY3uOL+ieKW0ePICzUOqs0ZlwLnH3
vlJEW6kD8j4OCUYjA0pZdqto0Z+iLripAw7bbciTlzCVMZWoKaN4uWnotnQp6oOs
MdcTC7ADM5a+bWl++DJYDUGjiuTFGzv9nMFQRpTneJKZC2+rDGW54N46AFYU3+Vy
iMcWFQCs/4lRqaXukAIFMXuYmVMQrU3WAFjS2/XRcvedJ9Gxj5Nhg+DuyOfECCZE
CKgwWNMnbl3tN2UgdPILsp2dhfNkvNtLorHIxOPePei2UxhZHk5D9XIsS0yDUqux
RV4OEnboJhUyddPbw6QaaTxcCmc5ioTFNUynY5jqNixMhcaU4eEFYLPQYnUASOeC
k19rJy/OpGK6ZEYFVJX+j4uk3uTJvzHrRVdiLpNJNic13sWMOehxqS2c16xXD2eh
6Y7J1I1ctKR88E8ky9v3ckWfk+lRD1Zp7vizDyRbhm4z5/eGmd3Yo+Mb/7eVEtG1
jcFwK96gxRBY3Luibg8tJn8fGrXR/D3kSK/+j4GGjQyTlUhjRoEe+1XMqPmJmJUe
zPnqtlJCJ3bh2LR14PlmdsuRY9oOFs6WZ4ikkXud8DeBmLPD7SIrOdtXym+IkTyk
Yrz7H4uRS/PvG6cwwd89Fm6RrrTISLm9U/v8mgZmPLFJ+2eY3jyAtxVQ1ba3VleK
JpS3+P7ZIYDwDvmd8U/b6dIavBdlnrU3PcdCqEkNz+8UxtkrE9zU9Ipoew7AMfw7
/29QABgcP618F6rmh+enZnJI5Yp0Bk6u+vpzmVFS9DbJcDxXxHD3X2Tq11Wn6WGE
ft88y2USJsJMcbcfnf/gw2aVEIn1ce/Y7pKxJI5iEznRy6l7MHFPkmIA5MGcClsQ
OZvkTWwgil47vlAHnPlFldq51tA5wt8f3JXSkqZ7E/31GMm+M6yaUers33PYcuYe
hBUN3Z55A5QZjqRXduS4PmTDwrLwVTc5/uiSI1yfr8gvDYexn28SszpNpHznhHJe
T2qZehLt8r6fLQuaCfBetluJPoCbhVwylokTUniXQgAWNTHi45J84uGmk0rXeNtJ
rb5zhNFCacWThE4YlzjbiUsNCUggnWKswC6w+3hfl02ZV8jCUI6QDp7UJ4YSimzf
vM9dxUrkDh4NvJ24PciWPTxsDfrUFrow24yasvQ8XNyRNYvCGootAirgVWYxe27t
fmrvTDB/G2pSQ8Nvi8RseLVvppDJXAL5sUFR0ZxsDtMoe6nbQWZOzpTF+9M6DYxH
WHxZNm0/hsPz6nOmtI2kUj3Qjn3fl8uOBj0mIeDwRMjuWvIxWVNWv6yKvFr9+9WO
KkUdETm2PEaz8PEZhJJ/ltxUlw7JKjgAjq+IXzAlBeyieSmUQqxD+bMm5ALOanHB
9B4NY7Xb9bHX7Wsq5yoD6VXHTD3w3fzcyL0/0TAneczMsGXwXihiCo4GUSiZRI+Z
vlm3Bk45KXWeo+7e57Wf1CFxcWe2sAaGk0z7RWdf26fI7lUyrNCqHGlY3aamkntV
f5DVBk7Rhr4900A/rfoxoWd31J563/fv+sdOzbltiOPz013d9+Gg7oOSZpm+uRIV
3Dfqzx9mwJBIFAJqjN7O66LZ2MFF/nF+asx5zfi+0ij6NTEdaYmCrfReK7fO1p6r
W9r4tNeDtANFpjM7waQpxzxYFFfJAsLLy0qC/DivkfNiLw5aLIxUgOTBzcDHjAPW
13dQtpwgXVxj7L/i3ri1Lm6zXs/qslmwbpdQ7HqPO2MZnenDtjzkFbMIexlNGCnG
fip8ClVQdpzP9xXshg3rRbwas40VfRqFKDTM1ebWqRZA+7/Q1WYMJFzX2qYG2vkS
z9SjGjfVynBIOKODmpHqZaZFuDpvMsMuLhICvz8tSnKWgth/DgsQDtNwkwrxNq4F
pmK2bF2n6Kx79BBazR2tkVK/JYa1WJu8zSNt+VEC6rw1jXZYnOYKgN+G7Lg75UcF
R7t5wkDgj0DaYxwV7NplPYdn8dqkA1bIQpbal8MbrbCu3MkIJcVGiIFoT1gNFo+d
BRlgK/afWqy0VC1Q+U9s3TfEcEDRsUuKL36E6mUXtm9QKQShr3ir60wj610WamXQ
cT0MTOrQrWc7+CrxYlqRgKYHhxBQhqgYoB+Ki942z96SFRuMf8Cczd9ZwpyLERsM
yiYKQkaI63iL174wJysJqJ78wiRHxIOoHhnPjUhxmWOMXt8XJaCF5pX/BmVUHOXE
DjoGyTIh3MSNzjJdctEJPVudDo1/chrVSxBKoMcGkgzjL6fJhDUfR54EIzOfEtDK
BBB2P+XpCYtEklXp/ocyp2B8hGeC5BOduO1bSQ26s9Y/GTMSflq5QzydT05VVIsB
wjQjdoF7lMJkZGYTmD/ELqZ4/+VhrjyGfM1gLOjmAH2lk7Pxjnh5L9yovhI8fPhV
/2BxzJTFrYoV75QJ+PiwKTVr2FW/0jrVaxKw7RKrjfi8S1NjFdYH6JjYuxYvcPpE
pQ9VmOS4T/hPEhXQjp8nKRMGM+cFngmxjm2pHCT/qxfDnEaAwYYjLSUyCCfWz3Ag
pE8fTW1HfIAyuNi7/4IicFdKKAecW2rrNBucWK/mWJv2F5xK1++nAAHUW1GTMcM/
D5wNGOqhet7IlsaD0tMlosZZ6nXPPOKaqEjLQw+HrmEC+sigJhepqbxQP+IULMu3
T/sIwFk0jBvX5JqD5UHUru9Z6m9ODW7LdUTQ5Mr4bTIDdGgxe6jHJQ1H2aQZybTx
k0a4tBhxycWSf93pA/tyQCtW0K4RVXAHp/GEGdErdDj7w7hcQTvrGkpY5wdi2G0V
nz1nlqg6KORRHALcw7XXQ3ljV15WH4KBkoZjrrG6kQpKzpmL8xL3WID96SFDZyfU
cEWIRFlkQ2FR8k9OeT38Vtk57rNGO7X2DK/ywvdVSwMKj1E5jeqpWhoQb/5XKXJL
nSea2yRc4F5zuMQKbA4Ss5FUv0IFy/fzPX4895QwJeCBSa40cs5Bz2Drc9nROBqH
ECs6SdLt9nu1yNIfYTgbM6Mbm58ZzAjMpX1exWQDXVOmVdYkleUYTm2ZpqNnjWLb
NsSeLRWVIlKf/HiHCWgx6UbKIpjz2YDG1xa61/bC+pXesqCOaVot/LyKu5HyCDX+
VA7PNld+z4giNKEvVrz9zIv9wJ0WRZ+Sm0p7o1sOInjjkxZXSTuzyytA6FYfzc0c
MG0pYv+UT7bziFcEwdB1inrXaNAAwR81qbqXWwpiy6on/v8pwpYAjYuRofGk0IxU
3IyuwnEP5IcXlALFvRaN+8y2Vw5TNzpNLngcyG1BNgeZBr3gJxansDIaoutSiXRt
VtJOtmhQyToYTCzzwAHcXKwL9otsHA2lxDdSH4JtrybwgoNm+6URhgt+fxLsGigz
qWWo26ItVPgO+eCA+eKAjsENzUS+jhhOvpwCkGSyeh5GAxqxULTXNnbSFbxXjje/
bWiyWOiGxYqiXPGYeKwNccA28mxQPtQ/e4cG/ETpftoYHWYqSNvc2ozeW5gCtzJX
Hz0sy9xHmGzLDyw3f9TfhXWuDn3M26kLnsBluNuYS2aXIuo/lg793F+A+7nPDaPG
avGeLnTT9z+T4Pdax88XSXV9bT82piPUml0LkFcdMweW6fHhpDc8iLMambcmFDsj
yC/d9JQkYCdCA2ruMluPgdmaf013U8HB4BdRSpk75jCROUhHEcFYe7cJdxK6EAod
Pr9xhIRSnrI887pWv6EmqhV68uY8xGV4ZR2okUYr6IHoQaFs9er8WVggKQFcoCMo
YrRKVqAh0rf2PcsG0Gp/Zok7dmkrTjJ91nYVwCAQUTISHaQDSA0QTVP/RD8+ighS
+79ElXU7WDUaPIgDc2LphkXzfC+8P752WCy+t4CjP8zpkBwnHMqiPIY+B3prUsVM
zy+edR191/tfs32SfwPRCPjxNZH/9T5lKLLb/VuIdGBwBwet/OG7SIwSwoiMBwfU
UJxBwjf0WTcp96sBXbHAhLJUBZ/Nx47Pj4NUhAiwGYijoHQxXFOZucKXwxzHk8lc
7HPJo6Lo0uSSUDg7o8RiOLszPkQ3cpGNk7xtaM3OFQJcURedErqnCB/vPG7vEEgT
S3MqrtCuQ3JdFABTeAdtHze+n6a2F3dYh+xe2W5dCVHRR2agqwTxRsA0jVhfsiqr
eJFfEzFtI2+box1uajK0zmqieFmRqNO1JrtWggcsC01vJRxvRjg9Mk5QSN6EVFlj
pr0UsVCwqVIgQFcFqphP/ZcbUdEJ0FKmEjRH13iSF8XasfSpBouelKeprNQiyTPW
kwHWX4UkQx+d2uzvVuAFNeqDblA2aaU+MH+tEnrMxaDf8tI5TiDLgKl+hW2R/Ce4
qj7esLMAFm4pVDTTlgzodUtJmCAg9CjP/p2Mn315YBjEguWZh5VMpVgpPDc61wsN
Z8nb8RmIq/B/k3ZHrZruPTe85iHDtnZ6mRc3gwFOR1+anzi5QCd/j2E/9rSc84Bd
zILGkGIElH69AGu2cauH34pkeWMvdOfPV5fQrQopP/eFwrzLtYm4R7QU2zodPQCm
ghrMbkRz/z+MW2cp/JuyioAVouRlqQy5Lp3s+Wi7EoBmVhzNyNAMpTKQxhMbk9Ps
ODKgMQtATWEKcofEvItprrcv9yMd6oBc+bWcLWX8E+sL2BDMbiVIfi0aJ5BPdKSm
JAyjHT4HWgm/i0GcmKMLhuiSfVp7bZSuL5/m/O5hbFrawSs3YD+GB8A437ACPWqa
UwoUd1zCtAYR15VPdNstwNdercl0COXBDF9tUCkAM9HbqLiynIaV8ocXCRPDbw+A
ZX4lXZj6AjpRq2ZwSuSXyu0IbN3vf8kRwhWJxv8Q5jOB526mOBFPrSJKI2T2TPag
3FF8m9LkHabfo7np2KCreAdAzia/cIxB0M5QUqd7IwAoqSWLIKt+QLfNO2oX+f7s
jzb0qfkAhpOV36cAantcfpxW5wYw4YEUuBWFZYNv7b3lZTpS8dSaiNlpWZNK0PBa
ao/K9HVwcVOHnH6h7euuL5O1HQZmM3ess8QdJqqDyThrAxghVsKiXQBMBZUVcrW7
C7SHAMV+uTsNnrm+tTcpxaFEPya4bUVScI1CQl0f6G9JdyAQjTHmE1P3dPEKFv+x
X+li0s1aGzOdN7JUqGGY9SloTo4mEbQq7tfTR3sdHn8/CVdg6M/qYn2hOU0obBXG
2ji6DDoeSgo6iapvnDFh/NKKOpc9p2VLk5JzUXGEZvRhcGxGH3v8Ag+xQ0mLTkAT
S+PuG71rve3o9ByuH9gw4FTTdJ4HtNi1bj1fc2wPInF240Lef3qysDtCjJE5lW/b
7TMo/YS6MwBzfKiIF6fUm7aWluthN9j/C6odF0VxzRRl5AEsPXpvaCAH4WCzvjgr
uWUi/3XZinoB+WWCTVdFzDgt3VtfY1I1LETXRSbpmD++eYd/pIgIL8LvXvDuMIg5
htw2cNmeLYn3KfkFbSo8fEHnmelUzmvA5ilqC08Wz0JjoGUmYWkCK7RD+Tqw7EfX
6WIiAApdHzcXMrjR5SFjA2SOhihnY2Z0lI2W3U0CgrSd3LkpsNKTfx+KZUSgQ8PE
ZAiX7EbxAabLC8SLDQZl0VG+RBL+BgrylTeZh+HgDQWCp11+P1tJ1Ha6BMH8UKr/
r+ioEu52hIUmSC7v3e6T3hFxWmotiXZ9EBunya1Cev2oHDF6X0QSTQHmMlRJAZVP
+PqYis1WJH5qafifoBaUK4vqcPFq8FUlLqnCgbXYOAcFYCo6IuOtrmO9M4ENBgUo
Ytnldfl6WOS+VSRF3Z3bzyEKxCU1rKzUq0Inbpp9uKfGXl14kFA0e1B1jlfGEiRF
jLHVzvBj/AfALQskFQHmk0I2zhp8zAE5KAxiz5Rhx3mZ8/XVjFPgdigbRFki2ExO
9XrQSeP4uZYA+/UvyxpOJ+AdA1SOtri+DJnkXIAPHw9URhDfZ2k1xo86v3+QfJLQ
ae199Klk15nDKSHQ70YeX+2/kw/yS05qtAalJniJbgyv9cYiSjpEBi8NQSnFJ0rk
S0PRgMxXJ0zIVFLRlPqrFajsNzTK1yk4uWONv+xNaw6H0MdLPTWMDJ3oHmgHdQuA
dZSZipVou3NYurwrzeBiODBGICX2QSS9oqw4Go3I/HtVAUXUCntF+VsITtBmKaad
UdDvmrUczxyY2D01tVgkjf28zF1N3uNM/1u/aAVnNAbt6b25qPpz+P7LpukmP6Uj
YeklqApa/UfaqLTBrZC3cs3ABqT3Ycog6GYRXP2i82Kjaog2U8lRmtG23jGXZJBu
BEyZX1AhAOS19kBqz62/kuZy6LEF+U9ORlRW/kjX5aO95kCmbwGFtrbnVmawfxy5
1EnYzDXn+SsOiUWhVR1EInLZg1otikfGyiVt574jRNeKsz01asTUdDpe12iyVBHm
tj7xTXe/OI/hFBLVfCTfxgIXdcQXLe4ChnD2e2pgRfOz7WqC4nrJ9W1XDn8nj+Te
Ar+IeWvD7jqsS6usIwMpd7RbwViOmQZlYA9ZMUp+T3+9szUgtBjSjRmsR2IPFBsT
CRyNrstAs3I8oeH7UVmMjslzRztV/AV78pq3FubKJGhfVabUXheyULwAy4vY7L4n
S1PkZ351OsdNPU5tfPhxE8uNoEZCMw9JjDJlof7QfxhHgQzYSRtowIWDHX0wouhs
FnMrzH7OC11DlDcvrjzFbYsJiJNtRLWQ7/Lmm2I/RKXxxQGtpVtWSBLeeq8jmHNC
RkBchSbjaRHuZaZZ0iDCpCNegVcFrwnoPCc965Kvfbypo3Mmpopu9riym7wOyuQi
Lbxu8J5YpR19Tmr++5894iQrapl1+nqmPgo9nrrNt8Nb1WJDAlRsn6Zw5qf1zTbq
OiqpPv0wcWPl1XiXdW1AmV/vsd0hAHwNWdgj2fpIz9QlcqM+q5EucrhzSOz5ZedX
6Pbx4aYl1Rt4sAeA5IKEcGEqHnxxQI1F7EVi9fpI35w0NKillQi5T0EAi/WtOi/3
zh5MgkYRTUlKUlCZN/Vp1EW+TzGBRFC6Bu+0JX4w3vTRcnPlOCjg9oPVhaXWLOh7
g/gDRnrPRVXI5PbXUa9ioQ3zJPg5d5ymTJvI9654RvhAHLTcQXO0Mvd5QQag9gOI
QN1D/WYgRHyiTPAM5PGO9RQTRqq9YnU1eVLlv1D+8tPkopwfQI98RyZV1hhXE/ko
NnOO/hTjoOogxETHekdiYW/KOVYdlhcRaBEj9R6Hj/5vpi/cY8O7iKZNVCJV6Ii7
yTEP3mbUq1PVTkA1SIImLWOZrJiQhRdwIjlLicJDtZDMs96QNjKdk7epiMcbmz0v
G4dqAcP9qauCoZny6l748qI/8wQ0h4iu7/5Ec5bLnLSXeNL939dOru5efms5WLcH
RfoWdex/B9Diehw8hR/XDNpULgAXV/v39V0z8s5k9PlToq/3ivUAO4TrVMDj3Eoy
RQwiVoSRNv1LVR51fZP3jropPFucNf5P1uThovfwV1eu+3z0nR44P2Su9tDj58bZ
YnJi/9zhPNHPnto6YfRtWifJ6NeDH88O7SBVxltX8qjmFHwveD/4p7aV7U56vICn
RzRWVrB+uQsUnmKj2pk9j/X7R3tSUNupG2GPapTa07SAhwyMIo2M0u65dhOwrAMo
mLTqA8KeUjcm11wbJ3jRyTUdbRnpRyWKFEQzI0HdOIRgZ8+No88KxC6v6sEn3ZlU
8ZDowOZRLKUjtC1pLgOC+VjuFjolxR20bZntTaO5l8New4mNqnz6T3zL13qAqRCA
U/DqY1OiPnBXoAusW6N86+JzQy/aNeeMcxi0azEq7wguDhIrQUSR8eU/pALj4E9J
sx3hPPFc8I8lWaPzMjY3CHki0UdCDV1hu3n7GtTzC0rVEpibfmqKmvVoRfiSVnrw
2Q1OeKKhj2AGOHLasQs5JvBN+i3tItq0fg5oIC9ev5LV+1CvVo84Ahm1AqjjlvN+
G3w2iEV89PxUrJ5euICIsonnQ3wgMjhIZK064DqXdUWiT4jhZBImvFzMixN8SbKz
bcu8tMDL/lc/2pSDSzcZOdEWB9HUFapjo0LZYISCJELj+D33qa2ojuabbLeulRoc
WI0EKoTr5IlYtNVC1BgS+RkNrRPK8t2dX11YNMDQza6X7MafV6XiB14PTezjwJ6x
9NsfT7OLsblc89sYvJse5vsdGW57zQAVBTFUCOjnV6v/Y+Fwv5ZAqJTZySVZqwiW
eTwVjGYDrHTC1fjC1nKG7DygsKKJ/dgS9Ehws2uEy2dYstk0iykgh0x0QqB8JM5T
PFJ8EZsjvnkgakK7B/p3WDm7BJcye98XjysL+LE5OVuzKaTZfASyjrbySiR+b7Nx
jJbTPiVqJPLUwPlnV5PdYqyblP1J88GVdizyFy7iVBPSuQ4YPzy66O7xEaujHqnl
A0WsFF4g2g6UtOaSr+u4uupevY2W/b5bDMMrgxV0oiCAuHRON6jDDUUfFYCjvfVP
f8VoWKnfIu4jjXgp3eDOEQh+2ruWnanW9S7OfL7T6MKKnbXyvF7N4crfp9jfe1wJ
NDVC8FbdHXWZdkjTaJjzWM+Y/unV8clNfRTxOrGU9WlMDA+ITVKxx2cVZMsY06dx
Veq9WkSqtKYW56ApbbW2FKkFIG4E5Rd0DaqbMuSVIBIea3tVQVKF53GH8KLKRboz
88IMddbcYPCLqIuDNJw0hjIhAiEgpvf1/00XL5MabpBwFs2cut9hlsm+ZNkZsoyl
trCMvuCau/G7nE1puFjUybcTqD+AipJBARa08H4HG2wvrmH8ONM+pTAU+eA5UmR5
DVNjsAdf/7rj7owtM7tLM5RUgocfTC9HVwilXb3x12gBdnraXE45aHqUd6PmHThY
qp/iMweBbiBhCjhN1GgUh/RXqcuoIa4c5j4seIwWh3XJzs6sS0CGaUdV1rEmPvGT
i3O7VIfzW8yR269Su3dGG1bAGcEuLXABw70TZI2/owzKq9M0hfErVwnzUm+LbZnV
jekiXxJxkywWT1acph1nunU/ApTApPN74cirgUwSqtZpJkdp/jZ5s8j6LNm6W+UE
Ai0MaymuUGAnJSAMWADcwJPAlTBGBkXXnhDRbJW23tAlhdg7HiSbO/w2jQ7kuJrR
abwp+cBynlEVcr/tawqEAppzNtHL0MvoV7gSpfbTtqD5a26Xd6KUTypKtUMbJ3uK
KoJ43MOrOKl3CYfzwtrVKo4keQj5J7LiuPFKEtwAiENU65wCD/9rfmsscLoke7e6
NvU2GmFwGPJXiLnteq67fGX+puT+NBIW/b+jMrQkLcpRzGREAwsglWzKczDTh5wP
7jxQvQ1hcR8rXDSpFZq6yDtUMHdPo+IIxdPsIWXah31dymBh9cfrMLjfaoK/FoPD
D1FkVQS/lW5nv+fOqHyyWbgCIi0HnHW1FrFsR/8mR7D4Nl12gArcbWN3ZAQZcItu
YHYwl/2qjE+/zV+lx8IrZKPz0auwInVOomhBSATXfxwBOCA1hdBRWg7JLLH7U5k5
HlMTqacmuaggztFJ2XVEFLtQNffmovwT1xK4z4WRIGpJJDRWABZWumIowjJowFUR
c4lmNmxpEzpTY3qxZkz2yJs2zdEjkx63bB4zG6TcJB3PF22EKndEeWqLKiGpwaPt
nRkpwcFUREdBCrwW7u7YfhmjfS1aMJxScG0njcbzvbCxd/osmnx0TRQ5bxftCKvl
YPRjiJfIprzezbRzyqxsaYuWh1kVSKyi37nXp07/fyeImUqTV4TowQ5BuwuG9Q2d
g1U1Z9RvvYMT2oPW8hxKZWrutZNYjtYkTT91Xow1A1jFmkNIBT3x1TQcNk5pPLdh
kJaCei7VE458XDwg8UcfreDLw35kVaUPjtxvKPNBuFoncnrbfxG+y98faOCWemBO
Q3PVrfiu1Mo9Fgu4r7g4kUmPvbiWmut7UZX5ewk3mRcayPMQYfYaZXIzkS5P3iQ5
PIRpm1CkjKCATqH2LE+QQHA2WVVURRzuf+NBwc7nmJUhaBLI08dI5EZFPZL7qqPS
5d5ymJoGowpf61fikNs6yjTs0CDDjSHR5+cw43oKFaL4quUfEZVgxnfd1LGQMsak
dXhFJd3QURNa8+SHkJyiSil6aLIQnfZPcQ5VXMxsTmUfqw1yQuJGM7FhnT9coikF
eBDXdaonnskXrNKBTy0htI8QIBLQxokcJCkBSYs6I93oUe9J6YKQii92pt+D6i7k
KXXVLn3p/EXy+l3iJzp19+5Q1g7E3IWY1GBocFJWOqqyYgWN2Aay4IP/jQLPVF9+
AYm8gUgjkzYvatP+Q+bavzu+G0DOVypPJC+D19tCsfArazKkWdJyDunrXsAOxxtt
oXP0jrNibTMgGwxd5p1S4e7DNy0tTiyE/oRXdioeH2DOvoRZluUrfsn+LXU08wMo
IJSK+s8IWFynm+Q4aiKYR+K8VFfjPHm7uH39eNpyKWtj0spaUlz+d4J/ENV4u2Mf
7swtjHVgzyxpl136lk0dq62K5Rrne0uvyMJFbH28dDKMfMpVkgE7b5eg8zqp7m2w
Ldecb5qrAChQUymYwNLUzBDrzwZUdpZ5aE2k01qQyDZ5v3/qLsaC2VuyE02lonEu
mrsffpjhySLPR/IgqHUG8z0h1Z0yMupLwNlKe+BvMz7h//D+7z766oxY+VcfukyR
ZrRQi4MRE9qy/6kRJVhM8qtIiI91VlSNiziuWgsMH4GFb6AO1CGj0uDEkwKJkcDd
CmFY5QlWSqQFVVOOh7ND+Lw9bWmmLNaJ6OLO8huighOO5B6E+k069xaQweTVYTPw
nNdb65wkvEWogHpRo2LAx0x33GGep6sNbeFl69AygxI8BwFGauJnBDicutJi5ly6
x8oF38FvJa9bOERMhDI8CwfKbM+1Qn8afhxP0TuhMQpjzESjtbDy1Ag2nMl9btY8
b19u2jAzkmzCUfe0ARglk/6AWPYshZD6msCPalfUUjYmoXwUIds7RQpUS/6h+uFm
WJqBflia4sdu+5EK56NjetzdkYTghEphOySzHjSP++4rjO9sq4Z5cLRP6n0LZDEp
Mk993031vBJwyyPIOojz+w3CSWxgIRPE87NcYUYk99kWen/EN4Ypc5dZwclqVWdw
Y2jR6gmrY0KDcW8Y6ap3InIzumtr+ZdwYPMpHS4H4GLTEjLnhVgKS3/7S88wDZ9D
mwYQ+iyURbRpN8pzyXXMB5g3SBIAtexWgVrj/mcnSNHHm4anw3PCJiKKdNqQQuoK
djhx38jmMsA4ZLqAn+ak7ppe17CeGCNB34vAE1O39u5jZ5lTZVF9wnrbG/9cDzvt
K5UGbESuxIcSU6uG9yJOnezSz/2b+50dNguBxGLCourtj+HhI2s7gswLpNCkATLY
m42QIx8HmF84i/7mmSZZHNME2kvZmqDBVGE8UqThZ2NrERJWiTpizoQL/dWaZSqv
B5lFElYFqpE1ZAXN6JOaALGkEnx5tob2iS8awXY513NKnh5hDjRkipo4xoNyVzrT
CH9VEd2/cLEuIG87nra6NJyCljhGhENkW7hEkOq09f8PPccwY3duaWi1KWWVtWFI
xJbpumobENXWm/uRC2BJ8tOZE60vR5AQKEgaFo4SEfRsifNSrSykXT/CT/9myPCO
OQ/MbSMLTq1RNn2bmRmdzCXsqloM1RqrASu5Vczzczc90t6yGw1vc1FoJlKXxQ86
XK+s6sdQp0cwCewcGM5oOkFvUWTNvK//0ZME9lzJye65+QjhUis8BaXL4etMeu0R
CXG0r5oe0jT9waZd1q3lHcGpx8smP86rwrNnGh/kZByw8XWpH0qkeCMtHSsitmGZ
DQsFJFFOMAPriI51Vck9l0NOlMjV7QeTvv0JHtSjJMqNTu2wluu3QlulHxzvlrbU
HrpKFPAymSInHAIpAG2uOOvSpTZViukl6SuVmYZWQn18pf9VJEZgnMpZah3Cg9PX
hAojOkT1wi728ISMysuyvw52et0ZTd1N7J3jXTDfyoQaVjIgZwhGnrRwRv3EPKou
suGHRItEv8EL6+Cm5hLAup0rRQlvm95cMOkziihI4u4lNVv5LcC9dkQ6eXYNEwcN
xNFOS+lM9xwC+s8BiryH9+YaQAbBU+cEUeLQPDaNaW5BfWvsoMnByjldxXQwtHPG
2dTjskouDMek8YakWvGT5rkfi/GsnEnZU1pKJL3XUBonbu9xAjz3I2jGwu2/Jqv9
5/tGTbBGNyVhtWou6DFd73AnTF3hK2LStwz6tHLoBi31hvwAeI7CSTHZW+k8YMC0
xqAT2Lu0VfclmCTh1R8Ta8YfTnbn5o+qA2Hz+aCl76DNHglsNSpX0erzQwO0yV/3
jdadOlVN+7cBM6BB+NaIS4Efy1vR1+elNtwUSyFmvqfQAgxXcKbE+hQiqfsI4chn
4gW7gn2vU/6kiq3eZ6mgezOuMAmCCpvLv9ZL9TQN/qgpOG1NMB4hr3qX9+MtnIn7
BhgmJ38ooDyyw4Dd26zM5jCX1D5TPOwkLtY5oMo2MdkGNHizGkhnYf5lx2fyWM0x
4P7woxMfri3dHz+t1v9jyeOglJf4XQcssZ23cDXxaTdYrxFfpWZUViQleyCocg+1
Sf0e3oj0RkBSjVVzfzpt5FIwDFXsOE43n1r0ey52tLdTc1Jk7dFWZMVisAbwCeeF
C2A7IhbXp74JAXd3mj2BpTarLAdJPy3aen4zMvy3/x7HZr0gIwYQuP3pGxvxrWEw
pzirqLBIHpil1rek99MZ3+vfKfiLHuatLzXYwmfcp4ygis/XIZCeCofw18FCFQJO
8c6gL1bXx8zFDkucjqjYcD3q2mOrlOpC7s0XxT3cn9ErBfeqi5nH2Rin+WPYeLHC
fxbJG2yC9VwV2X4zr1wWhmOxTny4SRH8GeuqbGLycDIiyiaLVcozJ9rJpnLO5mnN
azX+6euIE67r6LLAoTBHq/sXr02jlAu73qHdsO25oumAhRmalVFJJoCWLI7rIzQx
RNgefjCRJ9mLPV2Bpu9CfLIVA5LG6L/orFY0wQk411NuRDAyCUq5rBpjolRM8QcZ
vqVyKOFAwfj0WfjAXzCpHFVBQWqns0+eQt4xSyOmu1AGlrtUu+rI9q7auMN5A3nX
tvKflgBYEZfstD3f8ZGBOxxLEkJvtvLrhd399Zd+dhV6Ik/qWbH+PZUcBdnQBYz+
NSH/pqOS5DHVTd9xJWsStl2yZt/6bgBd3G+aWq3VnCPRopIfJbIxjAKzfQy/igB7
d2edz/Zsx/4ynq3IFtrddRl3TAiUeD+AwDT0VlrGBEwTALRAhIQ+5XJfNHHdDr3t
9PsiWxcuAZvIJ6AOOb/I5wKpjJnVf6FPCDvsAYX90RBvFLIkdhq/1w01J4RPBR/8
zRmdN3tzolnB0EoSufCatQx2eSYZZH8VIAm0i0TuPE0jZsyVsxwSClCq8WUrJ99f
g0IkTBYH5JZkw4aAG47TdoFrhDjSc8QLy3NyMBm97CQBFBLln2u4WV9pB6enPcHo
kMHVawaJ/OJn11I8hAH6caCbA9zkOu1kPwNrALLWqpHJ+rcy5LUyPko65S4gGgfs
Lig6fxU8clpzcRNrrkK+vsDtu+5t5WBbeTcFX8aZTtm0AyrKYqfBE+ptWrWGZDXN
YjTO6x9IQkENeZDgoZR4eJnpbZAKD8UWZfj0s7l3LJvmOkoR1vhajCGeHDA8qxoW
c4Xgp9BBfiS3ah2QFeMzf0JLh7WXbg4r9Jczm2TVlt0P1xztQmEPGqxakk3BCA9b
dSzsOc3BTeVRsNXKEHSznUB3/jlhqVzA+ILJ9psQcxDmKUh0E78qhGAmVXmb4Z24
qPLsB5o4ZBFPFJqIzzF+ww3fTMPWa3vy/Eo4zvYz7Y0+j2l/W/2+Qf19ZF8OMscB
EmyIjDB9TEIL0B10eHrHDRNUjxBW9qHV0sT4hnkkVaGbCbDEfcvqUN/zbzZy1aBe
S2RHF/bBoIwIXRvW2YDiL/di1pz4qilHlRvVM3jtsPYbEu7F2nJVC1f1/flTE5VD
Lie2NBTDgy4wu1wvtOYPkWchIDIX3+Ta5q+M6YGpD84YZC1ist2V9/tPevx02P4s
WzG+s3eFzD/iMrExvcUxxrrxF8EaC1Lu8x9nnRS1qMPljUx4drkFNdM37hq5SKer
9N7DrL17WY4MEKmCG/JWItfJ30ZoB33RkDeiNCkOp6C2rjOQM4fkKVk9+7Milwr1
yLL2jGn48QIqGUwFHSFJrAk5pLuMYFGIDEa1FhuqKKGYhJKiHH1giZ4l3bt2fshd
E1tFFtS33MOmB3QttpFQat/bH2WJZr6XiFEvBV25YMnzT1B+C1RxX1BlUw/TPQK9
5p5LpsIB0/svBuIBrTMM+ZlB1YrWlSj6iGVD44NeMqfGvV5QwCFQ4Ep47iTXY6bg
hsjTMLZbsa8butDEU6oznTxKLrnFvjXtEtL0M30hA2EgphCm2prLRk8bRK3tNqv4
x9bqVEYL8VkceRxY+bUCra/qXcmP+DrQ2oobfwrTXO6I3zw2pZ1owcjtVh1RfDsQ
QMd9PuXFYvx3Gce1z3qwiAehjnovPat1oZco4SP2nQHT9P8Fs6jCrl33ZBhXVJ7r
fdaSmTlykqcmBEE5SSJnwRjPwQNF8LbTI+eNBxdHrfPqzhtwRIGOPX6kTeNWhwKp
TySg5g08rw7YD9X4Hx3SFSikiijLskrv/MEAhGrwN4Y5RvXK690V/CfYguzS1b36
TXVCLoA5DKB9/87kMERJ/d+7e4XVNzPHigj0/dRJ8889XpaifwJwN5g83k2XB5ON
NYnu+hGlJjx0dYXlhmL45cFVUu3BD21WAEM0Z81qP10Ffuv56T9t4o29IBHS6e5b
tFOLV8RfQdRshm+ouacQeOe5xxh9SnGHCMVO0GJF8uoM+3XzMsNNdN/SappU7e/q
x8/hJkc7SQb0iEhha+Oudqi0wN3WPwiDYscAqsVWKmMNgd67YUxm7BPSbU2S5wIe
XlxYvei83FBlPw/FXb5ogNGMCeBbqpb2MNIQb8/gMFhqb6wIc/+9aGOpulZZbeuY
kp0apntI5kz/lWEX9fSAfaU5uPxUSOOiZvo/Zc1Zu0EJxnONeRhIz6VRfuGTR+9Z
KaeojPi621dA8ijWI99VdwJDJiejQheNCxSUYrJ8eM+u5t6K89/1/+l/H9YRIF0s
ih/e/t0XcjzByczs/NZI99Yeg1hRF1uKN/Jz3tMYCdqgeoPb/OAaT+2v+2Apl/W+
T649Tbxm4JoUOYYZf1TJpZbw8XYVFg7nWWZxHQvMS7JAj4VazOv8BiR5f/CzOgZx
hGMqRQQF81gHFXuSFfcl5DcsbYtVXckB79bHhLN0Rwi7jVIlSm6xyNrzw7hoD0Ux
dViSvIiupltmzoZKu+Af/rt3w0sE1J58Fec4h/FVWrOI95q0uJnJXBsJslwGd2JI
T1qhFFtjs4245AS/e8G5o7OsxtOnVJuPOAZxnDLxdUabNVyhWNLv14zh5j6bVM+B
0viqmHxcObKVIcZnsCuFojio8MgpKRNol3R1z8XJTM9M+Jhb9y8rAJh6yJf1ipPg
JeHauI637VRRsH2MBhILEOOoWEhJQY8dVwlb9Hfh/OXpMag86g2fm2+uefFxfywX
NdKGzJc7+ExZMBZnVfR6/pRThaX116fViVZcrUaFKpL44wZIXKzJysFlp00wXJUQ
sm64t7cmD0wTSaiXpRY3Y7pQ/reQo7YeGQv8xmYYkO5qU9KQEPETh9/d2MtgnYjt
GTOOM4RNYlFlVcvQlPaGtfaPdrE9jSRT7C9+c0CI01kNy7toFmgHbqr6xLHfQbqK
c+fbgbfgehANZrd0yhVLEwytKO40skV2PLbEGo0jBulLobn9ZdYm+prLlWnjpZQ4
V6Cep6lN0DuKcX1TwQM8KgeO/+UUIpWelYm+dOV3iqngkoJu79H/M6cGcJsLEX1o
gvwNmgRMDhH4XkWBD8J3XI6gf30063VZkVsmRoxxm51qDtRfjGqBCp7qrVjD3vhd
yoqk4D1BeaLq50dckLA7ZLDIw94n2tCgFvWXm4LcsCuR0aSqQBvVc97KAkcQsFwm
cq+bWPvi0Q9fKOCMVkccrMjzd3kSP9l++7NItMTt0Ss/kv13Pgl+ISCVPQZA5neZ
/pidawlbVxzueZcSI5DUAOWFppdT/8wHv6yKlP55jLxrWA0dk1fWeyZ7QFCG0zAt
IDN2gF5jfK4/dpqsBGx/EqVp3Al3juBrbrAYEmQcfr08G9pKwCTwwr3l7EbTPqGe
+Zq1B3MaeCZSuLX4U3HwmwZb3zXTuXrC/zKl9RYLJh2VX8nCj5VH3tOjL4YW1Q0u
CdEtCo26Hi2aSidiNwGumQ9qBr2sXxS+MP44NQKURUR9Db9NliWndHMUvU/sq+/7
xvUNwY+5Q8nuRrhVbA54i2xOFBXNvy1n8Rh5X3VBIpD5WSbOVK1IPQbDJ/PhAdRx
zGQf+rjHXksi/nKPzmOG7v8WyityNfsoWjIAPChdahjYdRw6cyIQYRC7ce4twmzW
hFOgGUVsLIKjI2GqVnF6mPgxsT24KLjc8IdGSLElM75/WuRpbV6JgBncYasSAdSS
RlxrJIw4S6yB3Ujbe2OCKjToV1M7hAWWajcbecPtyR6cemeFLgEsZVftuheVRUr9
EUUQkhWZgQDVhQ5ukizIaNJF39o18S/tGDSrVCCnuBkpGtHvvUIqM0+Sit8fj4Dt
YpGLe3LFrG5BFzRH/JYAYMMWhdUutAXn5jApRCOkAkPxCRdN2Jf2p2g3UmwVLiHl
dRpDJ5quIO4xNYo0mTFnmoPnC+0k1yJENkCicQiBc58VLhxoBwc1mafMZCShutNp
3lDN0NymAj9Q3rMhV1ykduFABX8uW0yJ8DcDZzWVWAgLeCVrmZccmkyFPjxB6Spk
Q8HXYPWobu4yn6G6w9E8Ev2vRx0uwDNkh4YzbNbFRIyLTStKoE3rkwZ7tzd+yVdv
tlIk5sQsP3QiaR10JCr8wtbCOsbQz586pUjCR6KBMT5PQ+RoBXRUcNE5Ash6TYq/
OuDW99t+Mb4ByBbYEnm7YUlReXIVcTGRTLEaB+DZ4YI4Ph3rf0YUif76T3mr8W0Q
2SNR+UpB4rGpa99h6NII399np+di3yT34g4SAes3slpQ+mHqHPODhkz+ae46ZjcT
1NCIVGdeCCUBrFzS+M7zqJ/la8pRsPmDH2V3TcHx55LEeaRZ6IJBFgAZ/9Htrpam
Dt2+ZpaYwRFtzaxGV6TfUjef6xFzRo8e+QvSKJnPOXrKEqomXVPFWMJwj+IvMpIK
U/ayIp+wCaK1W6QyWAxknYZHqCLA33YgsEb9XkyiTcvjZMrWRhIqxybcgJ0+YC8+
7qXqNdTproVetSL6MZNw9XyL1fzu9cFc4r1g9uDzLpw/0yg0rbTEKpCxsYwCH9ru
2/+L2LL5GuoLpn4VjsR9PGDtyagUGa52sY38MFYN5AV/3VW4wu71dTDdTGVPyNba
/Z8wYMya5B3Bnn1Rvc86LHxPrhmpQXMRq51aKMOgZokkSWA2qMNfALZHwwOVd4nX
N9TVX6pbcO1kwfx7D3/fdfTQLKeM0n/mVsVxYVvkOHHqLJHIXT9aa5G7eLZrys0k
5TfXz/Pt9KsDF9hm52vSOl4I/p9epOYAusT6lKh9KM9xUGx962PbCSzB4Hn8cis1
QkdXVCCp6OmcXF7+wmTLFaE2WpLQJ9m1h0k+Hqi+TvTFkMYP6psHHU4Uu7JBsaBq
BVQjknuc2YmT9wyKwWK1DPeBAoEBLpI72NBmhpGH+jl9jg9plzcvYa92gquzKT66
ZxEuQmCrdg6ZikXZZ436UF+0Ovt+LZdj6hr67UIhyZed7Jwac8M/ZC+53ZIu8czg
3Eal4fZsL57DRAu4CzcK0WczE3VRHCu89g3uxRKnfKSMiGqjvobNsUTYDQOucQYY
eiNQ6SBIIa2I3lSZGVazJTzmVg3JvVdeFr52v63X3ns4ZqgCLP09qXvGo4ACiyFK
byTV156xorBkB0BDCv0L0lCCQkoLeF5DdBdW4leWnDdH6/edFy80v2iqbs9R9rvr
3+xw9CBgnkgDnlnoIqtqvcQUtQ2lbFO+rxHQWs1unchmyA9yDaqUCk8R/kmT58WV
WX68w6Z+Ev9wtSXAGBUAXq47TnjJpqLBzBls7EHNSSV7e4ktulQje9fITDW8/Ws0
IJsPYzNZN3BhRu13W5q8WK/OiRhwQDB7oOKe+X15/eob6gsdvgy+YUrWYsRZz88F
jBkQ4NEx6kgK+K13Mo62xdeZz8bkIWhi6Iul5qj7unupBjfEBaGSQtoPxp4HpCVI
iU3Pe0TsFPjLJSEO+uAM+IggYTCbVVNJ6u2CyiSAzAXL6FfoPOUvU0KhIM8MMtjZ
D0EdZsoCPlOPHJEX0RPAv/ab/iTpDdvTFaY3/t4jN1pxS+0J0q2mTGJoaHzuNjvp
1b/aXhF+3L+2FXGZILHPpEZn3LRMNnd2toAFZJ2MnESJrAYZG68+BQalaZiZr0AF
FCFkJz0Llfco/4NnIjb/iv7b68frIXFRL5weSHwJi84A8lBPYQosfROOt16pgkqy
0hRkSCxc9Jhjy2fvgdSxWdzw1Jej3EQi2uinjl/N8j0qqtTxwDGlTQChkUT7XSjj
Eu1yGjTCiEqTppuELzVSC8PIXg2G/5Rp3LdAHUI4uAEdc/nFJpu8UnPHd44xlTBI
WK1LfBpxwy+t2CUfLUOFZEtR2mYeqRyd+h1JiKM6P9MWeR2pDItVtrL+PPWpa3CC
CrfWFbrJTvSTJWWkPXQ5LYFRl7YuuK2wVZbY+YyXzgAhL9BN5Sq6p/IH4z7ObRfz
ZPjgNHeXrJcb1bzlwAKLDPt/0Fl+LfRYs8mnG5SmX+pA5y2xJE9/vDNGZMr6l6me
vna1TLVotwyA92ydRZzXavJCM0yrgsgy+0F+FUE25n9wQjam7wFq2EVRbF6b21An
CitprKG4R9sYv250eq5Bn2tXVa9aAsU+dCPVCc+74sVwvVpNODu4VLXuGqnETHim
SsoClOasG9nsN5sfeieZ+mJwHfLNdFsC0B5Y4KdUJzP6AgGkRAw1QWgrImat40nH
bhVkquuxAEmi0WQ3p7FX5LEhhdi7bhUjAaEDJ2ofS0RebF/jUkXpTVoyODm9yEHU
qkrHXzMyU6XtbvG5jZd1kPQsTk6VJjgJRbLR77M0LRvj9yt7lPBQC9X1qQAmmCTD
/UmofoDazq0iWZSSfOgk6uhU6bPRBm5slXZSoW0uChxitu2ZVZCJwmIwDHQ+N3PZ
YCfwHZUt8+qBrU15oyyEyJnhehlJ4mJ8s1D7/xAt68700OrSl2ZTgZUdmriW3dVe
BzlX82ulqZ9ovC6IJP+j2CbBCw914A9LRQaK3s9s+L5DniLxiSlmRCEJ2bGbF+PK
sZ8RQ8KLCtURZVmxeZP73LQmOVpPyA9QiOlmu86lIRx2IRrPfX/D1zo8GooiDQ8h
lCj1WGmaicE95hynoSmz9Op6XfcJ3acIvrAIKG61/dnrHbuoHaw/N6Im2e5Kv9XT
/YCAe/YFedtlWc/f5EMgRDnCCakvlBPlNJD7T4l5vjbdnfHOamVdGOuSsi52eDk/
IgUVmaspXb/GlCGq/NOXpFh0rG9dI5fpoQkI6yBoP3+jTqUJlqtBzq4i/RokxxXB
87xwzx3ljR2DGEvnc2rVl35i6Y/BAdUVYdpFCA6qsnpOdzTqFDfJ8TAwuexeUBtw
cF1RzQbsEipehlWu1NApkk29441O3O7M73fLqlHpvI2KdLY49cvn+IWdELqssV/b
kwUehTLOn04Qn1mNRUumkuqtkbUFCFzpmChGo8CVQLNAmMQ/AdvvsdXL8EqhfBmX
xs+31+Y2zfdAr3I/WSgia2bJ54YWpQbnQfgkvS5CZ2Un6EH/+2O29Nb9p+2XFlKa
LAOCW0/iMm73A8VHfHNvebLm39EE1vpwoDTHM/En7yv0ywJ+BRNKItZYYmxODSXZ
jhg+1Ezpaehvam6srMG+glXpuhOyNW3Gf/hkBtR2D6Tx/Xye7TYxhT9qceEE+u7u
928FrQMJnea04OM+kRihw1DR8azu0aQsiW+JcXUac+ratdrgcQqKBg7+8UNQMW/3
68DYXx91Hr4tuhfOdUH3LjxuNGAwiKz+OPpovq9jabKzMVfbokPlv2TzSMxgbjaQ
kTC3aQH3uRXxpLdBnojH6z/BdBVDbfW5VDVq/pNKKAlI9emcPC4U5xNlahWyxjwf
lll9GNqWfW7ukpFD8bvEpQO9fC247sFgvrH167r5w1d7f9EnDGsTAmtYeSTGMAAi
1gByeKu+thNg5m2sHywYUIR1VfBee+eLdsnVle4Pvv/PxakDYBsoSkGk8GjBzY6/
J5kP2jAVk6ZhMPKjWb1AFdZFELhxj38WGMrJ1OddSlVVWsE9CZCXh5JnifF2Vsrl
oOTUkDavdFrzYzipfFIX8yx7x470ocymjIMqw4BPwkub0BwKubHZ8TyMwutGlSJ9
uqfS+sRfNrWe5cvBQ0hjxSIZQPC/Rc3iGve9YXC8GHMdboCbXDQZZonWIW1KFj8l
3o+cXEpAA78i4X5ZAaHpeQipF4z9LDNO7pbNCSlJAJNzP1CSWabHcJeq9VolDbf1
qvqo4FLNJ8SSDchNgFgKMpGGEw3X6KmVISqJvJZpo9UekDMl39iszY1N0G7rfeBh
MjZGq+EVS0tY54qfcftztBYeTNSjV9mKeJ5u0n5PmsYzl9Vz6XpNRVe0vMh+/kQ4
ZmuAjygy19WiT54b8nArIR7QRasOx0E6fxDe5LFVAUvS1YkVy43tifTqjgL77h/D
7X5tMMfMEP1U05TmtCYS0YNQQPyQaAnwkC448CD8h/0NINR17iUEiEIFWBhxCkKZ
KHRkxSkEo2Mud6Bpxphk6BbVJETfJMapS5gLqfzrmQ6t31axOhU66yQFyi2Qwy1t
T3EDL7qdx6Um1BQS6Hz7TRUMf2fTiSmbpLnDqRrKbXAfkETpKs/nLbGB6YiKBLfY
7jg1NZLWeDJfI7Olli9YqsHMsXImttcXa9pgRnDZdzAxnlsntO+FLJlmxfBPL6lh
9Ey7fsSoJFeUFuMzN854yX8rb5UHsrNiuzSGxe29rK8siH7KigtmmjSHLSKvQuah
V6/iSFaKfa9gilq1vJzNUn1x2KsNY7aMGwlGA8HrU5t8End+RC40qhbGBKDKNwwY
ZdJhCldg5LjDBiy+kdVLnex8Xzj0NVfQceQ4RdAGWpN0P29p2r8cGTcaodeIgdCO
jRbluyTkbK4zCD6NyQt0Iz8bQ1cW82T+TF6R+r2YMeBOxN+WAJOvrRU2z9Ab5h45
ERMnsmHACFnJ1nj+Y47qUQzu/G5LxMHyT+1hFYXS80/rk5b0vjbxoI3vUTWI6wbm
hAgTN3ZW4U31crfU6sfo/6HUWKdod+NLg54PHBuj9EvARrZSWlZhVzia1cFChVmm
KCgVMPjBLIPwL/KcQABxp3Gb0YyNI8ANjVPKSAAiWVtWSJ1ndVMuRSkeSJjzmSYy
qhfKpKNgZ7d97M3PpAeGbbcv9Sm82p/CDnafprCrwHi0tv4UffMJSCm7Kr9/4os6
Wq7O/xVuBkG+nCbgXkFJuxqpctU4sonSfH8W2pXjvnC9hyDtjz6yLtIWHzcSg3/7
3GBegTypbCwoOERD9Hv4rWaqLq/uShoVmyndxVle043pHKP3y2TEavIQBzBjrc5T
ijMngqA6rzorHu6/4FFw7UHlR9dwfz9UGJdy180+N7HRQVc8hnzq/X6gbIVtQtfi
QtaRZuf299N11mPRDFWF72h0dGBR3sCybulVq+WoF2Xf4DREA8OUImBUwaa20mv4
n+mvKeSVoPNQt/HbOxb/7ugbjA7VyUkt60xeipVUZULX0DI2E0+W7lRnzTcgy9aA
fZyV18HqI7bYq88yB/aKJiHCdZbV6LxbgkTn5cEkgV5kokG3pD/G63fsp8k0v14B
omjjnWKdkM8iNsJ/Up4/2ade2vkxi1jZ0TANu+Qz28lOwFIL+LHYwDQwxlobmQ2r
qZd41spKnNgqy1c5+rv+MgIUs1wo5nd2hIzShI7CQ/Z8weELgxbwo51y45soMyuI
PEKtCKENEpZfuYwh5lGHIfHRjoUkN8Qtvyze933lXg0rmR6Czn86NVWz80lPB3ub
xBd+kCS/xWwKxdXLBcK/YxUSA71NhBFsWSWcxoQkZJSQOf4EC8IZtzStmxoQJyzV
t3tH50SkxXBU3dihbVEi+inCCPNjc85IRYwy4lw/sTpYHjPISoxERPZjJUDKXA/M
ZwfAp0falkce4ZWEqdmatR67HMxn13KMTOlff077GCvR/8nCUuFr6mFPpdhD+jBA
eJfuPwQsbqJ18ppTwzwdRmFItwYPnQbN8iI0lumi2+1BwksWTAr8LIaIR8QwKkmI
VPexxQtz1VoZYARdt82mG9Pje8wTgeOUk6noPLStoiWz1Mg0dJfQFLzsfe29AKrm
A4jl20bOxBtOWeZjEKjs8/b2ur+bPN8zzPR5ElRbzWllxrWmDTHCtkCFdxymguQO
2UIxc5v24dIKGW0HMjV4nUPE79qxYct6mc0HPkCP95l1LB0LiRkkzmA1RN4O0OoZ
JSTzoYAbk/KlqBQg+qXoyd9LYLZC5DTuWUBDVNrjmoCmtlhOZRbnwTZmQ6lO98Gc
4BxtaLE4G15YzRF+/Mz2wLiLiE31uqXw1rPn/I1YUfe+VhLqEZgiL0YXLrHuLNA0
IwRnrLA0Jlvy311EHGshn3ly9bdjbzUOqv4LWfDFa1MISrqpVt8OUv92AFruxh6I
sXOgtQHKrh4n8VkM5FbX1a/qHh0anXv9nm88Yf2XD2GDuDnCvXNlQxHRBorkh+IF
mzj1aRn//GJRwaH0L6ki/VNQFYctsddoxUKKH+8V38kahGXevyIjkb+NfAniLxDb
RbknoZqrmaKSwFlhYHIF3ftgklUBj+yqNv2A7V8byt3bQh1dYbosI2xg8mpNnue3
7F+vbpgaQW2OTDJ6qMICkHUHZC8JTlxO2TDTI1PD4LVa5YxPXHNywNyjF8jwmJgh
03nWXqPAExY4VxOmvbU4NOFuoKc+b7kds//zMiMHmT56LO0rLHPq8NLf9Jobzm3b
VysBd6I671W6V/OyBqhUFcwM8T42ITOqRoL73BMnbipbPYhuxSmqlMsc3aygYU0A
GEDXDvuL118ggze8PdzNSoopcUiuTmx7MHe3gYEPwuOROkRMLfKjV0OvLA9NPJyO
u7KIJpnAlcy7+JoZggPOg0028fDD+T1pYCnqPsgfZKT/Hwe8GpXRTNmHfZlusQiX
nife4mS3axsuGC6aXb7shHOkuGYESs9EzRLAJs1X75BFsmJXRnLmQyeYPvlkzHs3
HeDTDoxoTHff2ySxp+YGVZi/inOrwXXq8dZuW0vZLprFis2rH96tm+QNUcWhvJKv
ObN8kyzLf6kJ+GTNl31OBpt8TtFDS8n4av8UZ//p65arrfmEyAh7fAWQQ/2JzRss
wmtgko+2CnoMabsEq8LFdJl+rvTM0+TOAoeVCKxYv9/yLuj7WKDG2G3WSDjoe3SD
9MHZ4XmgUvlX4AsZXVT94i/fA0sCTL9yQidy1qZDBs/tfUATJDERdFl4NxIcApsT
bSV/e1S2smoQ1ap1bKOp9zgRVy1yEJkV2i0CsROSeU+CFETy1nlEwZ1KS9D3HkdY
EWM7NEVILinKsPxUKo2pIXm4CXcxa+n+egOAkuJG8v7sTh9/zKZ0NjT+4bA4kNwW
PPuKjOpCrW06plPYv7eoAESZjAY9TgvvgC9XTO7MywV5JFRomJ73pCIcDv9TWxas
LsnqkXSzT4jaGYDvzd6SI8NB79IMH/yPsz2qnO/uC/W64ASrZC12iBPZKL32rJmr
52VYmEQeC0Utm3XRptx86ugeI8t1XGQhHaKPa+5trWd1tUAL8S3DEb7q8X+DrjvP
Tsyl8jPw0KeCLsl2hIi0B0ElYeFGupedzUdXKGPJR0a0+cWq94daO/II6tDymHJ6
Yoq/6viAyRlJ3kgl7UJioUJUMY3Waei2/mrSbB/aGNhwoYAVud1EC24kxDQ4j9bh
an0JMhooQuYwtaSeeeCslDiiT7J0nshlt9y5ApR50b/nByL3kAiKSwjRv9IhTh4Q
ID+P2QFnD3P7OZ4q3fvGxRFjfDHkr7eSEwWkchyw3N8sskCYfingtd2qGYWJaaCN
3V2psIkKMI3UNQ2lAFS2X1joHJGSqZXIKH11TIF5GT7sC4vxyZZSv6RmHS+hFWMJ
s/f0DwgRwSZOGAbb5hgsPBZK++t0B63RB/CeWWS/FyzbtHmGGtF0gzs62oy0tjxz
8LJVBZtB82L0yCh+CD9uPVXJsyFbxeBzYnzxULlpfJT33D0L1Plp6TNE1ImZ3ENr
FyUayJBqqauWbuJND97utyHhCdwjnDwsLMk/K92cBnSMkaMyhDwhGGypVgdZNb9e
x+wmwt+/ywGnqxapAdyYRuwIavkUweK8WfJ2zXUSPRgPLAsbPV1TXpYV2LikoIW4
p9ZD25IQcS/yitHgb7ydEaNLwnI75X/p+77fnGgTdxfIw1tkyZHZ1ouP48cyU/zo
Xn1pcF9ZQ+5CQoL54e/ixtmjSyrOvH/j9jwcspzrmOwsNk+tHVws8F6KJHEv7+TJ
iQZf1a3ST5oOJ9zsQTrXxsH2aSf8X1E+I6HYQ7wdrQPhBF6iJzV1kQbwSg9DQJUl
MMD2RpT3DZ57pB1GQl+sosB4jvnjPlA/bYYif2pP0tl7JeYelnxT3j6ALxD7X1cP
ECh9pZTFnj2x0cGDYLP3BNnm09RA3ZicpFxu1ehYxhpgoj4PO8d2Y4Q8A5M1rcA6
MvSakzmC679FXn9UwIdYbg1z22FGtM2TxDb0SbkNgfbMBVUHVX34iRACGsaNNKQM
Y4nVoBHN6cW1OCXeaEGiNlAEV6+/DwLPk2X2L2/UcKSFJ/9DK8dACBJzK1njWxmt
jDPK+dhSGs2TwXLiCdlQPCQ1/95rt/F/P/JmvTnXz0atUiPUOzWJuzuDlbwcuHvD
xWz/pRMsBKICZQfPaLB0o1dni2+vW+VYNfTMOiQ2PkRJY4SqkkJAnIgFihHiNGjh
mxiuk9QG9sn/LpsWyaPLkS1rEjpP72Ctxdgud5/nYTUuKtF9IgkrC9XH/iU00e+W
9TEFTc7yf4QV73/xG0v15vxOVTKOIWIguTbqotaU8g0z2IuXX4rMFvio6QcE/5VW
Vnv0MC8XE3Y+5LxL/nKzhDZA2NkF6sYI03/KPtHR8giEI44KheBAtXZNpvefx+3y
qMls0n4wUKZLL5h5aDm0nnLrRqjHDCeyz7/4T7svAJbeSbbnzDQX/Gl1Mv77HzBg
RmQoROn+sGgpkMK7ZTRPshAX3Tfa/Ll2GDi0edWC+krSgN7BKacP6uyZRYyNd4Pm
pQbUI3zQdeBWWwNZzbDFNJhladbAu8F/hI3vQdr6oWHbclpKhymwrEFtr1w48qcK
LQYz6+JHR60eS+Pjw1Yr5qyquTqebUi7T2hGeBSqxqBku09Ks9fGdpZZO4gNH8p2
DQTkaiH9UA0rZJFrPiPbtcdUlUthak1ZiQkZHc3s4Y3nNmaWwuckxS8Q1wZDCZFT
EdL/0yeqqIlEPUvdusQlHFgk9ScjmYlrdHGNkutob2tZ0RxWMXm8ye8POcNt3ClM
UyFZ9bxjdoCkZAupdqeh6lFtI7SV/pYEatJRBZ3p+W7l4Y2tV1YcdjE4VbgPUz2L
LobWJKl3C6d5vFPDO+SYuSiXvp6uWEUm7P435o+nvxJOPdj9EXBV85ZZkJc8F3w+
At6Wa8m0Lho7uSe/wufDZcrCGQjICLvhg0yRVkdsF/AdBx6RnRn0HXFWqatYmF4R
E2PvUH66N1CgYARUkk1yiwYYNEjvPc5HWUuv6jeBIDJMf7GNHhcp8+7YqhneABVd
N2kWlQzLiI2RWTMHeCtEIGF5S22ibqk7iPyqZU4sy47jWA5Iig4ZoEdHWzAjXeP3
jj9d/hkD1zgowsgtLJSgTKj8IPB6Zi7r+S5wgFdK71rum/FIipMXXiBtM+LrwNgH
JSFsjB6gCaWcVoijb4VjKjrkcrzGTqqhRZpixcN/C4BKJ4291yT5LxkWvOg6GGKY
y4+5hwJcsjBC/v0ZwgkvUlsy6CkOmLTcDkphbRIio9HpBDb4y4Q/9qhtD4V7+KLS
tutJ/emacC80NsOE7O+sQb8mRLLj/f5hLoLmWX5qyPeLhiRZZDBCD9a8S35kq6wl
ILz8ywMtKKDRNKkzrMQlpKkBhEAlP5pN1VNKWeJdu/saHmPiUwwv2dwfK86ZbZ7h
3Bq5suwsUs6kik4ZSlTQ+EJEM37RWFPl+AcevAKARQyMBrtKoLutO8vj1YHtTmFf
pdWKIa5yClQZrwv74I9lwv6jCnhMZRNZF5nuy8JoWs6NXfD96bJQx7UT8tXmt1bP
aadcS9P4o/UC9RC42n8+RXn0wA4QeIsr69h5xffLkvkVDcsgHhuirNPqGQROAdRS
bNMAGphsQFpCsFeCWl1O5+KdY3ku30XF8SBR++uXIBAEacg+TPNPp1qYbS63wKab
buNzOx8bnmyN7Hu81WN99TK/I5wMC4tXkMImaR6kx9aWRqq0ba5bNeuc1RVj1PW1
05v7LoMFVCutco3xDiEeNuNu/E7pJMBqz6HGftTywo2L/DHgIXJeHaeCPlPC581o
4IFVTQQKhDGxvpt4On0Y6uWASXcZZF4e8ovnR2DbN9s8oxoAIIMy2wmeOIp9zo7k
tarbMheH5kruLpvlqXV4JAhxVZAXUxSaD/tLHnkb3CmZ7bc4OWk+dh0JzB0eYSdD
i2R1JvNzD2zrLPZNBU7wwaw1PEYNXQlDZfkvhVZQVeRU7WUmz4gZ8P5Uaw/Uf79B
qQ2wVhhbRmbgeRNSlHMl/pZVFsYniTajVgufj6PQBgeRPn0uiHA0FmBvMNIdRUmJ
JpyGukpcyOqmLCid30WqtGZaJ/bmpSwV1j2OEGjaCWwacIACPEPVgCKBEXlJwyUV
GvCD102d+p1fEIKKyxdu07/MhkR2nWMDJa5ZM7AjuNWOky6AYsW3DyKpsVL6wriG
u3L2f9VM5PqBOaoIlSjQFIcFDS/XsIzXbNmL80fxGC8Q19Vef5FSLiS6b3AUURW8
nzbN2eKDz96cF+imqaS+mUi/UrcejiE5SmuHUXv80p5BB0YDMLEf1bfnO2BhxVSy
o6NZYYaOJENN30NkCFjrIaZixNJwiPtsnG9Z/yeOTQ801PG1P4m6rTSmKOBlCqrH
BemSac6PV5p/GE/ljA3S07uSLJ00IGwbn9e5fg24MJvB6SfyMigYww6SR4XGnuth
JsKAH2tM3wIXqkggW+o2WOtkBMvQUR/QkbG/WBAxQp5JCs3yP1tvDFecrFXwMRfT
VnUXj2dYlzk4A3oFndrdxH8zjjsLlPPCZk+Mxhbw9so+eRyuirZCgmqKyqMu/Vx2
vS4SsYZOwmO47eFfBCyvQSowsd5AIxi1/nVzzvEwR+SOEAU0XHUULub3cN6QCh6M
RP7kEblEUevD0ONWcI7vUs/o5IjYFmthDm7eb6OIwhvdqf/hSvLS7TGtA/OViyxh
knH9/CH8z5ZLzkBof41/guvMCi3NfpVAtg71DWHlQkYvGkgGLpMQD5Ah1QVhOHl0
HJUMFVcsSioHi0/co4jr04dD90Ut9bznP5aDYhu/EdYyuuNRBzwJ9hFrVFzP5dLb
S5WR+4i9574jwV8BSaOzovW/jY9VkJ2n/Kx1UY6qDQTzEJvhXRg39DG7Z03I3IoG
7L78Vp3wgeNXekfIF3Aa/1iWTrc2jrspwNNBiFv/29ld1jlDCN7J8lflTnCKyltT
NXVeFJHfo8Ax96GF7KCP6JTLC/Ctk8iW65UBGadSJyu2SxEEO8EmLA3u6YwNBamp
vlj3BiC0eLync/NPYQd1XRWVqMDuz5A7lBp3WpBY9D3w0CGZPKnq0QvW3lu1RqI4
Kegb/+k5HJbIMK0cHsqgd/7KiHWrT03WIzxLcxjLhp8lsUA/jpI55Zl2o88dtdt9
FueA8jxCQK8CvqMtnUM5worWKxH+FJurx9asdnhmSz4gMbBa8nOOsbvRDOcyaY6j
fEQYVslXn0fVlrcaJ5UsydwiJ6ccOodZziVH2PcSjy1Ll6GFRrgb2IuieXlwJsLD
tFPptgBKp5v4HdtyDHWTZPZXkTKCFl0Qn3FVpKTuq96b4pQjbSAl3SecV1sj3v9d
8N1lFeI1yS9Gw2GUGJcEK+wTjxlMZqFyLQxSNLdfC823hV2dp6odVwypwSO2xApF
A+8XRkpLv3VYO+8YEyl6LeQhse1CebJASjCcF0uTRGSZk8w6aX9c0IPeY0nX/hVN
R7yit2zKP9Kj6M/+1JRaq7NskuIq4k+I/PQdN2sBlY+NQ3LQ9x2WlZt05Z/Qe4S1
x10Sszxu3mGcb6RrUaM1D5W5oXF6EKjIyzaIjzzjGb4V2c/C4ZKf3tCO1s80rcr6
ZNPRGAb+qgYOPgFhYvxz31TdO5oWonXupSQhWJIx0FvrQcfzwKHMn9/J93L773ve
7RKdwrEnbgwOXS8xzkN3hy/Ne78v8BAFZ9OCoXhNiguBYODDuOZF1g9lH7yGCWnR
f5YYhFdF9cfHXw+KwwpZQGyDM2HRdrYuLtAnNoMb/G/dGLd+cMcgWRlDV7aBSlnC
+HbL4Z0uTGH0Ut8KP4+DyaFk9W9fiNa4Z+GcTBOmgyD/fQbipYezoZG9yY1ieByv
vRV0vx68J1KG1rUzIbrq+nql0wVf600hm4DKFgyC1dXII/Ns3/nDdEaXgFLrSX7v
HowWhh5pvX78B7zPV59A9BIuNEsGlBeo+JY79hgcn9n/s0dSAhXeidfyd/J/AK4l
My4QYueSzz+hOFWc0YP1nm+i/yjU+qh+ysMnhHgQOo30U/ht2RPCPIU6rmq1kPtq
eYWbrkfe3HqKDVXbqatcqKcy9ZDzYdoWpBoonlv7fMSfaya7U1MmUuc9XVA3eW+x
Ar/XmXjbq3Po7v/QWsbsGQM9IWCpX7XBGROWZGgPN73rAnNAdmCypFDV6TdtGGtK
nKIaNFMEcjA4T8P7BeL0R9DcvppxGtrmZZDgxjTO/cDFCAuzUOTMI///dn4uw15R
2/Eb6wDPQszkr1JFg9MNAff3SZqDklLzxqZENS9+gKq+7pTNhw5rEsE53wQJ7wM/
7sYfcgw2qbL4B7HYDXYpvNb8iutOb6JGXR7cZ21mqwCfEo3mD+O31X/bOYP/hKPj
k5cCR6eegFXYxpe5pco5pjLAZVEOazk6h3S0Rmik9Kg0KQZh7e/Z967zNmXWxe31
0nTh8uAzEc9Tol+ZL55umZF2dcqOyCh+Zhm3yTjUhakHOGbYXPmFwkllwyEbUOgx
ado8A1lHAfVaFSLtln7FzEsuXmz9S5MddGjpvR1uqi17NzFi5CdMBOiFwn1IYtIS
KHzJUxiBaWpl7ILoB4NwkYiHfzM5T0lfTTUcxYEOVq6q/QdzSVX4n8jqCoYR3yK1
8Yl1s0x9a//jf4NKGtEz5SSUPwLfFzgCDY88EOUhQYA1cOkUHFmOJ5yJZtX7Rc9p
S0lezdo2ODykjT28nw1kTTLqgSlUIdxRYsXYRkA9KGHNBU4heZ8iThdzIqhhicxs
Hfe0l55cNiwh/8sdoMbRUgcBAkV2T0Qaj3FJncXRO+4DINjFBcSG6ooD9mpkB5jY
jrY5S7KbjzqzLm+KxbEQxsOT+iX/qSnaBx449E4/Z+UyIaRPKukMvgepY3tnazAf
wICALHygDrFpneh8sD9YOm2e7SZ3V5N2USKgHzlgXwoBYIdD7l2ID7icy2bKXK3Z
lpWYm9YjrzCVFHC+6+cTTuyduKx19s5srTtJw0MYkpYsx1t2EauexLoFJ1gC5Yxu
StwCXzxL5MKzJr+LqGhs5yngnICw4SdyezxwK4PgGLknTHqRw9e3B53DjLJvz4NB
pyOEnfHGZKiNDQSv/Aa3V4M511O/+3/mCjW3YY4OJkkg0vci9ph8ckflgBlZAHhL
dqET5UjWW7+u9TYvCu60fBJwXadApkUp+Z0DnewhHwOfjpXP0NUrQCtfJjS43dEW
XvS0XxG7fBicQiFBRoyrO18Mkfyb2gUU67Wx8XRUyyFQoCAxPxQuAKOrAswdBojs
FPKbmZkm3ypGTg5QY4NxgczEF7xK7LUBXDJb4oo5z4sjECRj1EMIkdIvA6eEVD1M
VlWuqe4hUmk8Mg1ZuLWzKyhr3IqoUQs3+3rpc9qDLYmAYxXVHoPzLn/4kX/yJdaA
be5YPgHCc7qTou6eiWdHQgd+1Z5yt3RYUAt+uW1tK1SyrXX2z5neiT9QzxHfS9U6
cQg5AtAAQOOesfevKsynvlcadbmwv7hVNWgycBIhzM3K5lY3f+Fh4fQpZKnodvw2
hFP7OtpQshDjxE3XHLo2lLuFtiUSrU/6aC84B74HA/BzR5/W/auN0hFsnn4lvn6j
62Pybi+5Zt2JAFh57jQ+Fa9Dv56z23ZBpdWH9n+PlKEVWjl0c0SaJSKxTLlfQBoK
gBc2RDDElbRbkM0VDuNa2PDD5Oc86nmnNC6npOXhTAVvNkXSVqPboXMLXFES+gMm
wRB+Xd6hK08TyC0F0EYKUO78M9475S6HC7ECvlR6i2HRpubAOJZbDczcc7PpuqZc
6mx0K0a1USHh6+W/10X42A3Xp9A67hM5sYtbVap51aaKQakgvqGidbYykqpMRynd
jYodPPVzQ0PB2aC9l1GSICNQNlTqacm4+GiJYFGhMNadiuMs/mB3IX0OdPVTw9hF
lkwXBr8RwZt5ouUX+bw53KMzTB/4KfLegiA8OrSMTYYf1HQUDX2XyqeC1HI02RzN
ie6cbreiW8ZsGaConyytsNeIDfE8Hwp14z/4/gwcM6Mrp4HLAAqBzfkbbNUBj/XT
tT8uiUXYd3ok9Cq1Dr3RsOo3LqLX6UvjBCAzKeWBu6ZpYjpvVOuCbjAM8Pwzbu8f
wZniptpe/5d41KchDRSBfgMbWhCjflCw+t/OFthXqUD/FA0tRkg/9Dw7evw6ACf2
rOj0x7usUvUNiAfe74/8amUZJPYJBMOIcC7jnEIKsFpXsDcBns3NbREv+BplSUcu
OaESpW8uGoBWenqaum94vKmD+bjEcXzlqpPye3oMj5o7p23Bz2y6RIr8wInsPZLa
nC7b8uaRW6LuOjI/VnlwS3z+NCS8LINl4qo4MhpQhr3GqIjMkGdhAQQybd+EHxOR
bmRTjTNmwiiyBK2KOjr9v9gRCE9YVVIL7/hkYYo9QCSatONGjMUxnZBUZwyF6iNr
O80wOIgWRguWkUTdx34kuYrfy497TKrmD5glQYbNVRdt97hMurQ+cEQfOY++CcAn
nlA8MlNSrMllkARRQgtkYszXf1/JkoFG7ROyYlEHeAO3hczYzsaoXpRK7f0tUQKE
/i7+ZlRFlGM7WNcdOYy8lWfpfGdhUnCNlfoe+wbTnS/wpYIAASmiEUvRqj4bVZZr
esjkk6YrnKMsEmMQqt7yRk4FNTNN60yaOa7OvLGHxVDEIKW5wu73s5z8raScN2gR
yuScs+c+TF7cTaBG3Yd4nAL9wNrJCQwI92AFuoeaS8Z0YSAmRzAZ9PM8JhWOOs/8
kVp/WN/pha1mEbN+o6HH+9jWVE9RoBH+6mjUyU29sZHGuLXpj3KMHUTOHkkDD0YG
ThH8UycIgna7IdFLnME1Oh4yqTuX6MdTuAio9COKzQwkrMlE5RtJNP9XR467JAa/
F4hoAMYw7T8NcLSvbxQBmHE4hPsSb8YakxhrDRG4WYSD9lTeRdh6X6xhQq7I1T51
Ri7X+KhLiVUa/w6rB+qUpV/FHtdaLlzV25bzLJ8k+9mf0nSSUJOzzOwFIcsiE4Cy
tcTvt4WI5rAkvG1sdcnZLYd9D5qI+P9ZPRdhA04/82JdyMo/oTrmVhzgMFy1/0yp
N3HWTskowobaFhS2i4dVan8Gy+LmZUWJEe25dBl8J4lrEfu0d8ZH9HYGqr9gA4c8
1lQyzwBeKHR4tKWohymtu6dU2CloIlVGajiOfsZk2Warl/RP1isJL49kYqtFAG/C
8p8mZ/4KRdhYbqUK7FbmCfNu9dtxF/Japj457JQStjh2Xl3h+UnxO9XgwLDEqmRI
poGXLXXItFKrHfVXHcNz/UgE7ZZf+FHwWK46IZ3wZGfSVkXx7SqoHnMlfEmbRU3F
2X9U+rBrWpvVPOQLUCUvD92xLYKi7s01gpbSgJ/fpPH4yyz+vPdLvV+eNxAe0lIH

//pragma protect end_data_block
//pragma protect digest_block
WA9AVCOXoB2osQmhMAkRYRwSQcE=
//pragma protect end_digest_block
//pragma protect end_protected
