// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:30 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hASk6xlfMKQqj2TKIGmwgDZ91PtOG7CI4y1qF3EhZUgIoIlWA0WcTC565toM+CIg
sf9byYgwhxV6ZkA+4aFWa75F0mnMvpvCkdCqWX1koQxSUIwCxR/iE3ILb99hcjwR
zJZYh/3bAPRsLzDpY+Z06ePM61VDenFeXEypBi506Vw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24112)
3eo3ksYCNd+xdVDnwoWWY1vyaA7kYWZDJXrLLZrpZIGRw6C8dFhKP97otYsrGK1u
y6Oh6RJzJRRNI8KmmVQL1VbS6+DoL4cE84MasCVMwzye4YEXLSVKNkRmql45FOWy
zlubcEFoCgPfXp+waOiKvsEQq71Z0hftcrElNOrVTOwW+XQ5hybaMmVBWe53IKjh
6fNCEFflqGQlArf1iJbT/P22OSHvwrY3hZCi0nbEQ9pAGHD+6CGA9Ydjdn74q8gW
IizMiThSxe10KF+MR8Z7nzEAOt5WUc0jDzs03lv9qWLKXswjXGbhgPyPasXUR5DN
N2/694PeIziOOBTxRRSzBMRQrOF7ERuZUD5POm/usXvn6z9GnzaP2EZ8ZZ+7AXnF
kz/Gi60KrAZMU+uR1+uXsebyCrOlA18YpqZBkGYjTpmTbWVhMkHmiBr8s6/A/f3n
kZoO8Q82peOSwtt1sG338mgxfkldd0JBNIsT0C3FqmQxKHiUMjQ8Lkdbt/35Vtqo
PpAx2IFbuK5mIDfwNdLkz7xj8pyQ2zJNYqQX4X+3uEfqqXyC1IWyPhD2gQxfRoGA
8tPuTc7avn7gwaYGr9Fpzocw+7KMyd943SXi5A5vCDOhKluj9MSoZANh3GCzCX+W
Ek8M4bhUqcWQ52caFeZ/+Y+Fxky11bekbqdznTosH3ckTQ0D5mSoHrXK1hJ27oEr
0zxaSpodPJTzgbQCEuQmmVJoHtCENZO1LUtpwQthhxDDjHhVt7mpoJUsvuGit0E+
6jEnKqtCq1xPnTe4fCPjlvSmV7TH8bM/vY6+MOE6eKh36RjEWgHg08Xy6JWRiQyD
N42fnscEVcHt0kY6USYsH6Wxcppw191cd6qIN1fL9UziEqYo13Opc3aPGKG//Yl5
BtkZJy2fGbPlH3hk1yoBseIqz7EQc6GWLbEqP/fFvvw42tbat39+mgrTJcHzjNVK
dBCXRQAZrBFKWPoRVkiljVH12cZM32LbWstsOzyDQ2e7a0DVftRdMZ+Wzp+qeSmH
wtLIy8GIUa0scDn+eP8TY4lswYldnYCCm8czKaG9MzS3SP1AHtNd1FBmIwOgsUfQ
NjzXp+YukdhHvNxtyz2tzHJRYwyRLXO6DuP6QmsiWEUF+w9sONU9IrDI6kTKx/9e
UQdwwtM8RhLH3Pcn2n8hbfanwF6nT2LGggjUD9PLCrW2wYfJS9dfBUsvwVu9Q56V
sGkJaOXgPOY1RZU41x4NURoPa33FahiXC1c+tGS2bGrQ2wnf0sGg52h0XDmQR47a
Nffe8vdqd6PozFcKnw13gv71Ex5raFePZIVUEN1VUIdfiPPDYyAGpP8OCnOXwtlz
ghU0nkhwt2PKOoKSEJaRFtQK8q3H+ryiQ3LofZUamuNoaSts053feJC54wC959mR
BAZ+QszGIFdmEtUJbWgd/yJZqCOsqEo6jzsmJbltHv2TxoJqxGvaal2QuQIDqJBE
VE0XLGgeGMMoyQpQ88VxyghJ0Jt3hF04Rh9lPQlDOfMMV6XdejxQkmOOpWRXKZTQ
63eQC+QVtxyIAwUTdQECRbJSs/h1Jk19Gq3fy+F9srDAv1SDgL+DPeOC2ylajipz
RV25RA3+CnyQ+mXqdQ67jY9Z5p23jDFeALnq6MZgFNdO23ga3jd3wULOOCgqJihD
ibA1ilsK9ycZFHJPCU4UWhMVnE4rduQqsJZp7wI5M1K2umjBqPNeLUFs1XAEo8+C
5r/byweHjEBqJUW71FaNxEeR9TNbRrAUrHIrv/Y7Z5Q0aQebiolwMr7iGbmhRoYu
n1oxAyUYFPt9S+wFQCv5MxYpDqMqVUtkihFZYtAEwn+zyErDWWxDTnpmY5kPlFbM
GsymtswGLvWy/9gQRIGF9uviu7YjyeUzY8nAC+XiOqYY3YVj0212fXMjuq3LoN5G
j8teoogdXDo1RaYRfIrxsK1OShQNYtsPdsHMqcMRcEYVa7xBzxGpXe+9V0W7ZHgd
BEaAcu0n6xaSCyI68V8XmXJ4Tcqe4uF3ldr2qVif2v6WBCBmNf4wQEU4ISdInpBk
aA6CybZ4yUeAh7xJqCQMX1BsCezgwc57jXDDL6FqJQGmOemmx/xHPY838yFAoZjh
nVXVk3sfycfhpotWfOr62WBEON8vIk+/2qjOPxujwLUfdONl2UFOT3+YMkBNdK+v
LIuKawynkdLnn3u5OSVU0wO0Toesco3CHA0ITEb5RoCmHUvXfrBpIDxtxPCHcE33
ef+rw2m0PT5YpQNiel5QZ+/jstgB7WEnvIXmUfoYb5jhCphHjTmHzCozkG2XL6RS
kCcju8fmZoYFfAt7xhONS4h8GV3g4mbI1cxpMr16zrwWZB46r5aF7fXufH/Z5H59
MeGDXhXeYZTLvIaOV5FJ3S4oZOLkn+MhGMJ7OyoewXyHHvxLBOGdGX8ThK4b6TuF
L38zjGfmGlShl9ULVcbYu838yAycsvouPqPFpt8UV0aKrGj4r0gC6oQX28lMEVh2
zP/9ih60J+ZF1W0mCVzl8pPyjokNwSYrHN2Qji0kfgcnc4MQF+w1yvmU9UpnpOjf
ILIlCgh/BTCYXCxPjkKkz6lfDki1QH8zqOzyDExGy7oxTevpKJyEvvegP3xhMxNj
rOHPR97yDtcogBlQn/hjRzdpgfIZAl+h1pgMAxSIy8TBM+jyoLzG50tj/Dqz/nb1
7j9gAo+i3xZFCLl0kyQWUyjn6ugAW63NvYsgenpTSRi5jXvVRT6Hd5fK6Mfrt0YK
C89rVuuxDktoNOhQHJRGdwlZNViWfQB/EuGXfYUV0u4PVjN65deFELr5ZPEH6kGn
cfJm9RbG5U+lwY/4K25oL5BI2ggHSXLuuPRHmMOD1IB/TYVh/p/e0IlQSQxlDJ+6
6e0hiMcBxuCqqUX9t0Fs5cGf7t3/2L+DLM7OzCaDRxv7hMiKYypO5ZdsrTqPNel1
XopS3pHYzWRHfNd+mhVqDl7Af0+J0ygo+BWSMhri6l5CgibQdutm861ItnXxg08E
zmIJbYjlFp56JXNpNGju4KSvx5TICh6CNXrLv/lQKR9/By5OO77WBv0qADmlDCsD
sGT4GCd9lDG/sxZAtKp1V9CP9jQJBe/2cUR6FxgQaobc4f5aPuyttaPH3bZJMXUW
RT1scHAri6FkTE6Rv2zEXjJ9hvTMy+p8LsuHPk6cCUPi9dgWztJoVLwshz83HnFy
YEWmnKn1hKiDJVfeSW7jQDdoNaeu27MWjkv/wm07PJiTypzuQ0CaMFiyuSMlEWJF
Nn7jopUu0C61k60FP7t6ulw8nvwKQmECLPpEU0Nt9p2w4CC3yC5mpXwp37BHmBma
O9FPfsAU8UQtvvw/6Zu7kJdE6eoTGvegRtNk74dzFCZ3T+QqMtria77lKHvFapcB
VTiyQXZ+bK7Gx36ngl7iFe47ha3hvhp3qJBhBdmVcvvyPmEyQqjhBzr2Qp/s1z7G
F9P2ZQlx2ognmpB2vNm6D7RdIUgfaPraEydruJs6b2fRYd7OkeBjKVi5ETL4Od0D
J+jDKKQJUUfYMCjBpFbjWrjMDZd0W+UcrReKnoBixY80uQcT7wGeUH3GV6mC9Rgh
3auWmvke6XGh6yaZDmwNWnm25O4zbM+9mxkOyYOPlV24ohqXGRIvuwQa6Z/N5xsG
/dGLN7QoiG4sh4wmmKi5ww6qzZ/h+W9tmIJoPH+ND/W9+S37pmjp9HmBOoqC0+yL
pJjP0xuIebSo+813S3qeXptqNWImCLjOHIjd/GWZPkZWzo+vG9Rd6akYDJMTnR6Y
mIT3bZzuzJ44Em61C7pqqcLI4olgIq5Vmphm+R77a2nu4BN6sbhB1GSB0P8WKoEu
qVUYo1YjFVQ/fI/0d1ox44/OX29b4lc/Gvk58xwh8b3bLOQzIMdKEnN+/JzbDgNu
njxZh2ucjGuFtm21dOFfKfpbeQChtBoLJXGTBUNuRhMeO6NK0smY4/Fn/NYb5izF
AiCuE7/lNAoIvg3sbBDfNsG3gX/JD+zwoGey5ZY9+ybvwniw6dHNZcEsByYFotSD
LYRpJF53a3eSDHKufUIhTuGhLSpzt8LO9Ma6eNRIqkBU2q5CoUjwQAlwBv6VJTOu
2C1lEcqkF+hcjB5QagcJSivv6K5xjH+hX1jUbPa1Yc2VxbVod2v9g2cRsMQCfaTm
jiH8Kwoq2KKUuYtkgOZ0YVI3p1bAHY5dFysIzdy4NbUDCtQLC+YOogNiiEHpgme6
ZCgpH0CSm++zLWcMD5Mb/oVJJmODi+QaRaYjifv85FnRCj8KuU7DnIhjOafAEVd1
0MM1yZLUGhJvwxGBXi5hhWskretMrZaTvPL/l4nBx8I8g7MH7qqnUyUxdpgLAZgt
mjmqJ9glyW0+Jr0c+n/eUQQRL2Mo5uEefm47KVrj+NHTOdS5POAtepNTyCBi9/s4
h2tXyx+DfAKYRxu3EhoCZv1ZOTJFPLxbShX4EHU3ba3tgJMLNs174DqAimWDZiR6
THBiC1xQ/eFnNZfV6dwAQtLROjMwjFNy8NvS1h03egjnh7fFWguon+VE1Fx5FzUz
sDAjCC6SLXi7n9o6+zeyqxduppz4paf5UTgQoucv4kNaujTSsUh/C+W/Y3DC+u0i
l25SQP6OEhseH+lCDodkm+7DahO47W7A8AXpd+CcN19K+JCMiPrdp66J/210hJiT
Dngj28Cosm+dK8/urUONoBYw/HNzorqIkO/NElbrdIG+SJpB0YzWuhL8fqOdoqVF
KNvDg7iHSj7KM73G1wVSnG2P+3nptk1WNpuP9B5P7xhXemwtyk80dHdpUclb5eyx
5qWCQZOOD4lKLR64LVAKwguG5fy5rup68u0FNPZrvKwwF69U4QanztoTkR3dJeg+
M3x3/SglbY79nd6kKe4FUFSb+G49orV87zHFuk3MAG4nCCOktm8B6ER4Y/ZVv9Uk
8ZsQ9kzzxaZSSJgFkHVsH+ZEm5gEZnbVGekjUJY90AIuWzak/vtFQuxck7lQAG1X
LQ200vK4EvTf7cfy/M59DQSSZaErsKI9YuPS1Jp1vtIzZZD8tJcIh3zGmpNeqLBS
pf81kfok2I4y3qHrs5jSDJGzxO67h0gDsK2NKsQgUzFHmELmkrh5DEeV7H0LOaIQ
MQn4rwZYgZcWoSjZTsgMnKVM34yMBUra0ntSkQRpYR9F/weyGQYiIJLcS35ZCdsx
vwIt19yy41PsEi6TacR2AX/WS9dwRh8fZUwSImbTrcAvarkLBSVwVxf7OYt5nZQO
5wEQNfLP46sO8vWiaBh/drnr9RJ5Z3I4UsJmwUSzzHZEfA9LL/936FTaAFiI/xBX
IgfC4cg2uhwoVewSTuxGIJe01m+hQmu6C7k2LF8y8Dj4PWHBjNhthatq9yB+ZHtA
WqcrUyCC6uH6atnBf12YTdFNKeQtUFabXSLQhGGJB2fphu1QO8qAQSAxabmuVBYI
KPXmBXmzjSZpC35kMjPgu9M/wmAvDPB1jTgFPxbu3q1OJRQYdsuP5tLFw1qRKmi/
6x19Jptb3momEOb82+DL7pPNBRcaXflI25Lj7c4GSlqFnUPr6KRhlRTDDWzv1xKC
FXjgKLy9vmJcJ/XBTuGSHeO98CtI8mdbR39Ns7B4B4nR7SWNzOiUbBlMphjOnUwh
HE+0nfxd78LP7iM8CCAGSFzD9v9LTQ8H6QwojeYp7DV9jQrAf/r7QaAeBBtPLz2w
cz2cv5u6IZNyC7Vk3rE44RF5x11nrlCAZq83WBphx8UwfVcdLj9zHIJlV2Z8/gIS
X+bYPLxDpm3Uj/kMTPLeNroohiADmiTE/dzwGHfcrekeWpWSYkRKyCyqc208d2hK
Y73dUPfN2T4GZUV2wQXMxtmjjA6L5Pd8LlUUSAtsm/3/XBvoChlmFrbgx3fdPMBE
I+22qLqRC1Oqn6ys4ZXkxDTt57EeKIlRR0OCF9vgNlAwTMY/BOepYk5KrwexTWN6
bwPsF1G1gXPVtVxzHIhWWApyReOyVlf3ZfZjYusbIZ95lpmAoYfH4NFu+AblQ8pD
E1CJFxPvAD7uDiYOQcV0Hv9Zj9lN5eLb8WPiesKhU0Eu7WMoDoQV1yFHj++10Zt2
XFkCWvAHK8kPT75yPzw6z0GAaeAgNKxmooEI1321WxAS0BT8v5v4XuxdQ4z6/RcE
OnqKABSaoENHihNN8tm1gWKKryVrDe6h5cKSaXpNmDCWUM7T7MqUkpZK7GVneX9R
oom+44QeBZHz7LIT5BHhqrh190aYQduB8jLXIeeJCvoPzqXgCef3WX/KKS3dCv2p
YKz6dCd1qXbITPVPS/46l31/msQyuLSDYwGeXG1uT8brWfKDPHLd9eZcNAhBP9jw
dObbYAmpnPRvPrqgybSstDOJhVnma23etQM+3L5lJwaNGAMFpGIv1P4SV6ovlNeP
9smp5JVjNq35w40hBNNLe2jBtqRUV2/X5XACz4J0X3tLLEmZSVBxz/YnJ7/4RzAQ
xKnSzJ9TfsjkolrXcY21EavH154CPazVGDdO1FerYe1Q3Obi2rniKhlY55HcahD1
BNS37gn5zx016PejnsCZrT1nSB1i0oZu8j6j6F+dLAwE+XQTkb9ze0zYwf9kynf6
n13jADmV2cqtRvgOPLwu5S47hJYOXK7c8vOA31w0q6A+ubRjmMTm3WNkJv2kLEVg
t59VnQr6N9DSeEej+vqVr3R/KrSyoQMjd221TK0v4akUorwpl576oyev8NYd5iMy
I8zol7S7qx8EM/cFtB79qIr616kX3i/Y2gaPDZfGUpQKvFHwazoXus9IsrulBJSb
i6gFdt4z14TyzR789JVlPVQNxgnqKdWGYFxxMwWcmHj1fFeCS9zCaAkiB8WdC0oE
eOZr4+awxS58e8VbKpXm6DyxKd/7M/nKJafgEHuCyGaIcVGsnx63cee8ZbKT7z/f
UwQkgXRJRc6fwRjKEim9zg0JSnO+I98xG6CmrQyj01/le7KiXuqabyAhTkKH+MQa
rJDIGD3SpjlCDMDCOhPcyoWKRVUSjtZS9EfXx/2xBNyxJPubMRuM4ZYMbTtMSsAz
zkMsMaskpNd9c1eJaMY6jkVSt9mtwBisXPiz2I463OgEvQnan6KX1MHEuaOVxooT
W2wrrCLY+maE2odqdz4dEGDupeyaJvIfHvAxgqchdqqMjFJ09tlj2EMxGW8nqJYy
68lHcUAQbtGChIZSq0RJyuHTzcEJHUnDPDe3uQpW1nD1GxnY1juKiR4wRoZsy542
JSRMUv6e4pUi9SsnOUeoUXBkW4gEhI9K/qxmWmjVGu/2ZV/1WGa+SfJTYogL/CNE
WmkNG/M6x6fOdl6swPcYaAp+pRqxZ9I9tBtemSnw7M3v7WxIyGT2IKvHbzltZRyz
I+lIbBRvkKEgKzL1u2bBl0/hHOIVamn5X5OhgXJ1pIjasGgKwfZrzdlfSj+IC0Uh
seVtegJUtPIlEHJQnadGo2vxcCO9N3DTI+pe9vBfDwP+MWWEyqKKHpP2SU06p+oh
AuYBlyOnDociZHzGSFqYgcyqpk/r2Hi1nS5oSUIu5ERPuaBbkcP4tFjn+DzIAEaI
gZZV3f1HCKzJX1cxatEltA0vklW03MEvBFaa0rccdO3xTrcRfIBR/ShyosQ2pk3j
SKZa+7eGcrgDJN1P2fbgO6Ee8bkkwn3wvcCJPyQxnzvcNBhzMNEaAqxF19Z/R1E2
WF+XjERHuyG3Dtl+Hi4J4ll+Q/kIdyF65A8nt/0aZB5t1YZtgUGZpEiHlVMYUgp+
S0BxaCVi6vwTfF/ztd4n/wLn6jWuoRt7ES9PmGZ6WuYqE9GOtvMeZby19WFbCaAy
744Qf1bGW/r2B7BpaVTq6eTyNJg/JrdAyD+n/u5b68cGxtszuHczUekH+kOlt3LA
lry6teyYbfxOALAAgOHoxmPx3dKwQyINXVQyyRukJ6h0b4beSYQlmagV151VdScc
P8VaFFZMncwSizixgdww89LATbJsCPB2Glue60D91dw2V2+8bzWD9r3a8upqF/VQ
NAWHIRYE/xSjBZLB6ArimS46iA8fRl2Ec8+T4bxMkOOzzgJqXi+MMfvrVQKCCtWj
nUQmNfdwUQW9qidRcJGXkyeR13pqr3ikkCjH5EtLOh8WtJRHWUFFa41ZsDTgOdAt
XYEZ5CUjbTOwSXfcGPBILzUhhZcSWZfUrApknIGwpWlbRmwyE//Ng/8qTsxG0e6U
5X/qw719+1XQB78Z1miAUznfFV9/0/lJkp6jcM6YcspBD4xORoCGeFEXbVMszxaq
NtR/ifs4rF4/KWNg8dkcra3bD1G5X3/lQAodJXSFu7gtWtaFPJ0JqXeFD2WC99Eh
UTqoz+UOW4JumT0YCpymdfwyLLM173X3oGHUd5zhgNhMXSs0U8eODYROo/hFI0+z
ys/UOjAS+UYpFSzIA2CjX7v+Nb+JSCDvgKRB7W4PpLhl2uQJTrXuGhOzDp55kBk+
cjyjAIUULYjSJ2UW8plk+1hQWMB/wEX55PTvklxREk5/5EWD/3RoD21Tx9WmxnSc
Ukw7xPVNoUKD0/m9ocmrmQQUTmsmhKIHYCrSIq2xiJ8E74h7LixJjXUW3Mp1CekV
24cDG/30sXx9UXRS6cKEmV2AZbv30qoswrjgUjWkfLKnTLl3h1c4Y6A5hlc+5Jcs
xIaA++oJQHlBgo0r6rin8bf3o3lMclT9/myIUBajSMwMTEsTE2gj6igWUv2xX4uu
07kYELRQCm5hsbAfYqKd7EZlWN+fe2MBURZLAGDc/4cXOJIBh8L4A1vqqVg/M4sB
msFe+qSIPGbqVJn0QlnHoRemO5O4i/VWR7E4RqgEgblLWYr+jETNJ685oWmS7FHW
xQjo+bJ9AlpLKKJwK3hO/jFv0du9UDdrrkkJCmBxl2TsoGVwyJSTTbdVinvGY3KM
8N5K/DAnP6JltiOEYAJPb1fK3hSB+7hFmzW1VnIDslphPcGJMV1EbH/g/FgfKBZT
C67PcGD1zM0r4Mfu2UuG9YTyGaTUsPIIRsvVISX5grYwsdDu0RfFBx9RAxTdzmGG
MpiMAFY1UXrSnL6wc753wQttpkukCabxkMOJTqaRd8sbT4XCNQShMH5Tyhk3afJc
R9lk5u0vJiWRAS3ZAb9G4xE0Sod6Up76ZsIXvHa+3pzCaxYEvOMutTAcIpj96Y6w
voEXZNQUZ5yJaXJeaTdevTs2o7OEKWvl/xW1w4jNP+kwGKn0IA0capsMxC8y8Zed
QnbL4hTLnuHLF0sHZz0yjTY630mTQpHwsr7ApEOLT4S4SCOlcBZlf9H/RC6Hu52Q
eS0WE/3T6H3O5vHt+MpY9jAIV2rnGgqiYzdNxkMnILv8np5Zn/1+aXl0t55/z+On
pOcLjVwqxc0ZpP/c6YK8JybhCOS8W3FpebJH7lrBgjM9VAyByjc8NffYcNLH7l15
q6wQFS7yKEF4e7hr+UFdXiaiajgn7hKyT+gjpa1yA0j50BAhiiT4s3VTIgiSionR
DcYFHayoYhEr7ztYXs+GVVrfyhxyuPIJGx+6BNSDRW0iNWQ92BV7D/YMMZYlWwkF
n2Bs5daK30VxhNzhQhDm/Ga/0VqjjbAry5ib4ewHpw9RjV3wTcwFQfWQ9Jc/YqIW
j5PQuJxb9rrMfhwE1sNCGlFmGPrlk/aSP+RbxqQ2WyzzOT9/ETNEStpdNRO7z8rN
qEx9ZPAvbmmtc48Azcem5XTnr1Kcpu7Borz7fY1+3ITN3FGDpbFnc6O+hnCcBndS
9PJgnxk5cyGx+Cz1p3RLegC5WwEs2FL2lyjPXT0Ev8s2Shqi3oAXlpR2yPg7cJal
1xura5qj2+oE4w3CKLBlOyf2AdehZGrVFeMna4lqoIhY3mak0hijtQbzhU60PxO0
mDprA4J2Swb28b7rSj2SvWNBnstped5Q6RKHpM2sUqnwgqsOiJtd5to3eciT9BN4
08HQ3L2xDI7Q8C3wiotbV7AWnOWBAnuau+nrjUBC18xQFJmkoUa+bz97evgGtoEm
N169KMWo/mwRnXlR1zA56KWLyrviugsctaVbQmwH1+IFEdn2LkB4fOzcZsX7NxL/
oz3SrLcOMulcf3H6jqlJXsksDkGlUyCSZo4pUtWWfCdbfqjeVcQLkkZnp1lgqVsG
B0C8VxiM2aBK7fv70aKOIgei1cf78u3kpCJgu4siKhVNgGqORmQ66g5paNEdxfhT
y0/IMqTNYC2o2LM/gN0EHo2dGAhwABlFfrmPJaoJBe2LZV1pRSRvkrz5gahZA797
1K+ZeMRsQ+9KuAL9ogTkMp+C8BtDsNxKGJNwUp0wW2iysjxFxF5ajYJys0F/+Xu/
/mdA5krrsbAR9CtrW70n4bpk7Tkuc+1b7azQ88LrZuWnXoDGsh8FgMw28veVoowp
vCzIxnqeRdVyIrNcGrfuIXGqZBdteKSg8t4VEopBJYLb7PzMoNYUoMGbWfQkahpS
oVicvyTVoJScVnAPiMj4YLlu/jhUMuPAQ3zXREj3TuBiH5m03BEoJZvYW5P+GmNb
C2xbIRDsP+6HO4yd7SS8Es07Ohkc1zLz0z0mMImKESq+kLydiRiO9Rcp0kNEyFIr
m/8b6aE7wXq4oCyE5OPHGW5ivA1kUgMWp8hXVCp2LIOcQqAcxBXNfmii2QH6gH3B
jqX72K2WYK16d/Amj8kfd6a3zLp+k6nhZkszPYPhxbQmN54ieJ3PHdUIC2JXYrG1
38Pv3l3hcZw/J7HwmxIXdZ/c45LUmP5zgA4tzM+JCRI9VOwiC6vTHvmALzagv5q4
BHW7jrS63lPqL296te0IFo1QiaD8guASOWTbTYtJLUVjeUNzX9R1wmV4GDaJ64KR
cTBy+s7IzUSZWpmhbyK0llREkZMn7c/EQrdWT3q/esiFhsIFzzKx9TffDFiqEwfc
BB/sBzoK6gycbC0rlQ1OttVWenfnFBvCqnkTNebe45EptUjsVz5CYegoMYwXjIQw
O6oOQ9YmI0n/p3OQ+V7Dz2oXMICAXpEpPGUOq2Vmnvo/FJvPo3BSAFioSR50piCS
WMeQArz7VJkaMBcdA34F15iiTfAqfwakdo4kzmpJeNVlwHYHwjKF2+6ulIkT+clM
jFr5RhLOSIYVk00MKrYQNme+6UbgjM8mUwZjQ9c/NwTiMPFUpHSZPK4QHaqtX+Sx
wkW6MHLoqk3pKvsCwaZtu09gZCaTzeUWQk+tcYFbbsOssHa7R0N9+ngNZTx9A6vF
o/8fb/pTgGPEqgNq521z6Ki0qak7u0WXAPzc9LuqTaqBkjlHZ7/YMT5JFw7nfaul
a9cTKzjo9y5VTxbS0tkcW2vyj9fAyeKmIRYKOB5Yjep2FSdDs3Sr/C9qpw/sww+E
+PqnXgm1Pw/MAphVYjGpaRwkURclEBDCmFdN2cN8xPXfrYT54hFSmFVY2rGb58OP
kcusAIL1AXZMsj5dz1WcPmgZ02mCy4QgfdlkuSEWTRyGal21RE0dZZ5RN54cPdDT
pEFWsFizNtlPyjI44i1ofCf2OWRoTYmQh8aYAD1MHLrfhEKGoVhKPnDzyB99B8Xs
mN7gzhBgzgGV9XKWsHGL7bqIPqraxuFDgH/wUB+I653xTE0v4KG1cQ6DEBmVLahA
6tCgZaOy7OsT9l4B//QOMRVb88aDYkezCepaLSQXR0QCZWA9ao+uhCbUMledXKwg
SnEwB1WWOLQ373pSSGvXEVLJnmR+CF4vei6V5hS+FZB/4jjIYGq57p+QTOqdygLB
8bnTl6hTlujR5fvUSq7HN7ZbDPZfzuB1SlaHKtT1RgA3WQnC0TbXbL0zH+/emkaO
Y5e/zFpqT88YAy3V/ObP5HDpy2GdbkfiDrvMYYhVnjXgLxCciMMp35KpmzfEt8a6
u63RSRGoJA5zggDXKw9TJoLhzIE/k02UaZrypVNAEuVpQAp/N3EDy9ptWTlGmSVb
o2EfRRCqrKZ/zVj4YpeGUQCxA0kMBIUckAZLlBFgV1CupGrue/P5+ti2w9hizbFx
tOgUrAAb2LxAcYHYaqEm5LSXhPgjS1vbbIgNR4rzfcwl/rO+xmjq7aBqJnHkFm9p
K9SleRmfxHw6hR1BjDJadDdTM1fdhHjpziLic3GvIerq2tOQtBzdWkPHoPGE3u3Z
/YIBqOMqQldYFyTut8nmbUOVSMA3wVvdPX3URdFzdXc8+dvDQ6i4iAcUDzySSVee
p8fBAg9zIJ1AlZ0d4f7VzBkrqHYLFBHEcVoR9yfI6wwguoXkHsnKqXM8XvsX13Rx
KYltH9kNTK3ehgatTgp1EHZD58zg0fetQDYOdGgrySMTMAXKUFE8/BVfzg7+HrZ8
sSfCQ939rhAJkc3NJepECRsvLy2JOF7oD7BnH+I19avbHYGiRNrhdzwJRfVPY5FX
K2kDSO81fKJPBkIZgw5CqO9O8w4XpIuM/BqDFWCOWcWpxh1blKRQt7YsqluANy0g
/F01SJVlgNAEDmMkQ3pG+5bP+S8K0pTl1HDfxIRYXSLWOQEp3MrgqaKLQm5NmN0l
DsawW4g6FaiP1A5fopzleQKSd3tsVC1VbPFrHYJ+2gNwFqd9xdHO9SjiIlVdAAuf
By5Zrr2LK9T0Ci4hCp3wY+WW8XcLfmv1eB9toorzHRayxBLN4ZZo+K0a94VF1L/k
JmngSsJyymkooygV7R1rjQAuKqH88HjU36EZqrh/gHKKD219ajHmv3U1MHIGdwIc
6ioZgo5j1yQqvZPG0VOX9mqrfvE86s6nMniWP6FbZpr5HR/de2UVgZq6l0gcACds
8Lu73JIOjDef0X7oZUQu+7fhZAqatnJEm7rUtK9UeMCmTatF48rYDTOuPmmczkai
Oz4AaB9a0GzlaCyr8LypiScNpaDGs+NZmXz56NmS9ouZWcLbUzqTo6xreiL41Ks4
3uPviyxjEuktihPHO6MmnKwCuQ9bvipSR/HEbhXR2dsH6tWYScTeEdMygZxNazSP
sCO2vQnsKVLld68Jbu2gLIX66CyJ0sWD0Wdszn/uO5k7AoNNIbAsKA2zGpSgyOPz
HFy6GZlBdNaNGzc3cZtAyom7vLydM+p0cIVoh7GIdYLuXAFb9GeCTS0EernVTMLi
N+lSGWOSbJc2ZQQTT6VUaDkv4XdMD0RzCkH7wFZ+SRjOAyxlUeTN6DsfglP3K78M
71C1iN8KdQ7d+TWGZSwGQbj+zh4j4imFk9K0v4x8h6MvhD85OYAyywUFHAJcf1IJ
5pdADsuI8L5q85lXiYdNyM//bLj9c1tuW8kPJ7Zb/3qRpXKuuHdZqBjZd25ieuRs
BEE8kQ/UVdLSgbDMnDt9lYIUdoelA9ftXltdi04iaIE++W6cbXHFZ4GQZsT+RqZr
P2LNiVui/AW/+Hr0PFEuiGjZxirQuLj7dFlBPCBH0LN8GbI0PXo6THxYEYjZJRQh
PElD6tmPM2fWRSSL7UuC+gUMnvZjTAFu8iu2qb+D+AwQElBV7/rvAJA30lJXB8Ws
bI/S90GEBnAXvzpBR7D4BffB2UU2cF3ATQVn+3qkH0MkX3QVbd5jbL29I4wWY6SX
mntjPJzovVYfGD+aS0b8CDnMuduE+WxN3TaCM+zKPf1S60BIzTT/3zmP7p1t3OV/
EwB3GtJyXQ2CuwpIgeRXPKjdAN3cJ8z51o7XhfczumO/qc5IgYatf+nb+EoRXrjX
QtDH71cBSdqVG6M6orS5LwU/nvDV/uLaQrldV+Rgugqgk3+moxopd0xfL7YXbtOa
zkJ77xmOyBmUK05Vmf6vEOrYcusDO3BPq3nlIr2mLdk8xf/jEQkIX3E1++paG+mQ
QpCoTezNJbBbVCX509f71/DiIpgXjCUs4d5E6xKNyEQn3CC0ykDKzcaCBI4O4UiI
IGQOfm6QEVkFozytnWGP70ToMtFdnJrFKCBDsCwZVzI9z3BB6LtGjrPoOflwQ+ja
WCyDUay/11kHH6fUlcMAJH00UdtHMoGkaCbb9fFKx77MmVWaRwHTOoBx9ITlD7c4
JVfUKnY+2pclrgEMHVKluOq8l3sO7graXr9S/gXIv5Yu8cpAAc5UUFRjWWG8eJPY
UQiFKAkqDegvG/ZZhW0JjbfrQaJdPcif0WzcR8a/h+OiQ8gsRarBhPMciqItY0js
JaEkWJOMJJ7PAhuvU+ERwHmHG3NZE/rUo0hGdEsjuXMxcsvNkuO63J2JyJ84SUq+
DKZErL98w3Z83M/clE7WzNCdBR2VQHrQB5GeoUqQTCVV2c+mLgESyxM1z4umwsFv
JqF8bc+xx6nt/HLMB6XR+L2uP5Zt9oBmBYefKSt6pJz6MSSCAtux0q+ShfWyld4K
IQ+WHuty9ea4KMgU5kELqjnk86QQaG8fqFrySWQY3H2FHLr4zdFWFHU1PxJTq6kf
DfE4W7NoG0Js/c5AmMtGaGuaJHJnS7EdqbM7O1eN+E8ggaWrdbZzdi4R2nC0FSjL
MxisOWXGrpjp5KAvCzzXwrqKKoqM8jcABNJ7G0/TrA/dednVw8ryOIyQyIKlPRtB
53bw8jYDkoaqNQGe+7B6Km1dVnKQN/eGEGenCcuZuaKUIsB56uMowkQIc23EylAT
qZLEG+pB7P6boNlFiUz7i45GzCeqXPwGVIXxIfu3JX7Vc3QBk3+yFboZ2MoJh9jE
pmbuY6WB5L8cgkLjznb+F/20rzvuIXbEmgblrT3FmQjlDtUAgIcHJhrFRWatVYHr
5QkLl9yNay/UE46BVFqWkq9hyZRIbNxtPBcccuWghANx1ClkBXaMpvdYkJdmmSzR
qBsm6YEaDE/tUWMCF4OU/08nGIZ1vnFuC21Eqg6hAn1D4HQb+48ye4Ddfwoc1XUm
iaqvB/QRCBXqoyzvCM0V90SI3Eocr/csTgZDvq2mnEiyjlMj4FUxPgPQRZlQrDKY
C0Bm8EL104otysQJlY2mRtO4HtR1nq3n0UtOT8IWZ14IkD9HtLFsvgOAmG1ansJI
zsejiGn4rcCN5rT/310ECIEKuYZvDjL8h+TYwzn7ZoQS+jv6JGu6hTyovwhIoxus
EH0hpK/jrygcepTI2hvMMKs8pVmm4bJIYkcp3Zahem7dAqzVbWPnciHFhVgrcVZG
2ycMDkNbQfhQ9d1JmdtmRcVFxkBA57w6D4PZO9GqA5xSBLJNCjbbpG0C3anRllj2
voold2Kf5Ojx2EKM7Ffy8Src8eHveN+Y8Yw988HDzreM0d7Yi2xAl+3w7czNMgXC
uogZqPenedJo5UbvMFYZBYA8u1qaKX5y+Y/2Bk4aWwu9UsFXBnJaHZiXfnTIKLz2
WylWuoqh+iAKOd1kjjrMn3cGSeY3cnglZ6NEZuT/SRjQSiPQEpjm6FL5oDxkganD
1fiVtDkJEt1ev0oZW6Ez2D5OhO8doMSUiIA91WhQllvCIt3xV/tRV+W40Q26oDq2
pQz2JiPeB5weMagvz+mAc7OBqIrDGdUm1mTO8fAJ5JL4JRixHDey+xeTCWBF9gK7
2Dz/y2q/3GEmuCYgy2DNm99GMegR1utuKIOqEKbpNMRTxMhA+Al6I5hJPUlQrvYs
GFgJr1uVxkJgZRuiT0tmiLIdCtLSBgLQZ2hz7wdHJUY6r1r/g1AskQeGDfX5dx+1
M9uMAFIlpok+wDc+8eI5YULkwasRcqtoYZ49l2ywQQGgGilgjwcDZnKK4e0If5P0
NjGeALWVkZkNnMj9WDmZUByEL2jPuZM58mbEvwyTmXgaPMQPIB/ERjSWuQnxHFAR
02EWOptQGGuPQPhm8wnrFMbehfqqIX3+5SdqOGFNrM+aQe/ap9Et6On/Zs2h8SX0
YYdW6elSNHcTHVD6IOgWgF+9+ti6i8APzRVHhsubrkvJq8VB7XRIbhc+Yipj+t7e
bxBkXcmr9G7OVnfM3NEGShs4ia+OQsjly/BxSqu6zS6mHreXw2qm6rWuVz6gIAe+
a14+zf6Sj9GgLfpqRDHuMG8m1rB1zR5mngw7gffqvX+NRq/Im91TOzEae8CkYrpz
smY3uuEwT1WKugfw8FPVvO6G/EkTofv50JbAtcEVpdR6voi/SzLMNdlHDMwlpFF5
D65+2S6WpI5jGbj+/fQ7NJlOE6MOGMpe8TCPLF7L1uwm3N6A0rwjnJmNUN7n4VwW
7rFSmwV4V3VRIh4IPwfNRFp6kOEC/Qwpxihv6OWrbby3opJIlZg8CtyszTeN6qPW
5Kpyg3weSaAmoPXZBSTqks0LD8zf6zXWOy/BVaJjQlYn6nFr/zssTIt8bcnpV43c
5Hc7tqu4iSgFMGkHP+83lpiO8Iy30cncmv1A/OrouYx00HnNmKy8xipHwumi6Iak
M1nUugq6KUqu9fRuogE4Ta81uLdzZmKBCDeKx9CkkYdw7dm1PhlQXN8H88xnRn1R
ls3YBl9GUHbQlba3zLIREnYnBh6+pAGGoKBAEy/HgUBEUcCGcHcj7Au5Jh8KQsEG
04+vx/qTzPqou0tZ/r2dOoNQYdB9xOdkpoIsZVKMsf+kBzENcraoMYkMpZFTsXzV
CIVvqriJ67DSUdXeip08Q/4MAVXu4FhT2PXz1YOSJNMHO8LuaeJgjYUbYFPviyy5
/o/llE8RpuogfTftJBQFq4FAY3eJQejPH0GWLG7Tj2R84LMuUFBUT9CUsuLsdv1o
9YQRQk3887FpPB5jfPPVvm1R0i3/fabPDhctw0dynpv6so68kqxv5BVHfq3mhUT1
D88XGrzHvNCnqtBk+26ZjE4MYr3aafCqIDLVWpFm6l9MP19+LmI9uyHK7kS/zApa
ZMkBevVvD3y5osCWfhVLjejv5IwLTSsSs2Ny0HB9+4slMytkKJGAjA6C+EZ2cIM3
7Z+hZNYN3fu+bzmcgwPBLGBzmTDBqbf2SZpPzzcTsx65Z8qrq+0I9RIO5jL6O8zC
ujdJt7bpwP1JANot+efBXKUJdbVbjQMRhNY02EGxXoY1JjrVNpBmo0yIrNNOiMr/
jWOVA9x39mwNOV/TZAi5YLmuGrwEzdcn826jvUAGCAc2EJbpLEJz/RS7lbDLtA/k
IwJ4aYfVGXSDZFExBqonOKV5tIQFkVh18vV0BhxHdnsfJm9DDyrq0kjyTdHsC6vp
/bwYUIurkcwteTYJ3MvHhB9xLXG+JE6lggirhlZe7AdM1+GeenBjuSV88pIo50fL
kYGbdhB0x/Qnr7KGCJdUWnuCGMxMHFtwOhYFstaD7eSmaMykvE1B0KbhLtl+cHI8
lisxBRNSXgGTQPTPFsBJXBbCNQpoFq2amLseTACdMgyvZDxRe2Uu73l5KLDCevlg
DCnjyGmgZZ1hkShtWAVKs0SBG+dHuwYS+w884e0UjiORdXhxv2tkw4BWcp0htXhj
EEAqfsTPjo58f9c3ltZwTJARYzK5U2Yg8XQ9q8fD8dlPNybb7jX0ebnvaL4qjotc
9QVI91Qj7cfwbscXw9Lcb2aAJgPN1ernRjdQwXI+eIzf1qAi6+VZ7xptLZPizi5z
VWNhAuXSJjOLi0FGHb8MyALaqj6kWphitueNgdusPZuQ+9Zbwx4aMmRLjiT4ibPx
TxeDbbRNv0A2b+kvnfeIjqLH3Ib3tap+kzA2Mp53Zo9tG1H04hayvCpdtBfxPyuK
+hxVVIbKu8MGJHGz4vOrqYW9n5z7gjoxWZJTXtA5zOfx0otDcUsVv6P1I8fTX+oV
VyiL+5mCAhJ02ON0iNsyIrDWaCcXeDPv3JuBpDyh66UpIE3gt/ZNvU5rBSsZC76E
pLC9csH3NtSyOse6g0Ti421gqP6yZdcYLekH5erg0hHurM78WJDxMmvfGizFLrwW
eCoYMMQPhqhpVRUIn0mBVq3ZVFV7NgLVgg4ABXt4U0wmXG1UsKyo+/xd3imiaKrI
Dnd8/O/pCmmytbr0IL8egeFrY4rKSt/0dKMgarMFJ1SDZPNZl6msqVFJy8A8yhOH
LCie3T8cpS3HlORAXyqt8RDo9k/ejPNW8vp+UYqwCF4RMv5jPPD6y0BrWmhfgS8o
JUTgKpyrKTpRN/iuk+NZL7QgSXx00bUMpf3sAS/dpB7j/lkjaEHWW53nOCXzmo+y
FjpdCT7yStXGwROKcqcA+RdZmyOyWP1cd/03eSFz9oOCMzE605KGBuyyUIL6oiPL
MndX6kncld5HN22plutEe8BU71y14dk34mjK1SnnfKwGGjDB0yWJdEiwoEwu79aU
i4XNgL1ZXVRSKckRYZy0zgwfBVkzxv1JYVpZwxNTJsczcmCI/lUnjF8GG/Cm0veN
CVdmcli2NPQnMP0aHdACQoIZyfjqE3hyUwWliXzlFag+T83H9l1N+CezqkPhpW32
MltAeecoumr7vpKMreeovaui1vekyZP3J8jkN0RreSkurWlbgVpd42zT/NBmsS1w
4EqgkwtM+23ouFkyBNSvs78zYdxs97ORzdB8V48biCNfSBhK7sC3gNUMjkArZ6C7
9b4sGykWjAtWddFtQou6xYs7trQd3RGOC7Mgf2EtBcrc9VzL/tLbQHaDcSSERbze
Qiz7ixmwvTHOr+8i/s8juc2ihQ6Mjj7TfsRn6h28uCtRRX/FatEZbwXz2V5Rhles
PlYY9y8v8wmo7ThX5+tewSgPNiLVhdW14jZd8mrvwbglNNOKbv51EfyPwLN9DkVy
qYgO2fzg2i9UkanyEBEeEeb0vEd0ql0kPD3oJMAIl6U0/tIcmG8mesbaKeVTWefG
Uggm62CbSpbhBKQw1rnZ/EQlc7mQQ4XwrsunPDgXcJLlHJR55HJ+NlhiO0Fs2LDz
ZPPq8+szdwZH6Y6zlhBbkxa/WMXJOEDLsdZtFia5/lc4XCs4Eka/vk5g3nti88cb
/zA18s/BEEOqyTeq8LtYBnlneYz00cZHTN07myg4rbB4MiO7xUlMx5o4KuVCVefJ
QxdpJVjQAFAmmBRcRU7WuMAWw6BZfEwfePYjClrqM2Y2XNDCZhkxC7soZkxH+XpN
PLcNSLsKwuk+mXJ+zynYxVCNBUpUWZElVlRfGOg9Z1MzxrARDQQ46A3ek0nGPJNo
IS68ZYMxh+2YUanK1K52iGVpDZt4tZLd85KsTQjbRAxMfIWqTzkGlHbeE0me41L9
H6nFWIaaMOO3oNOcSqIUH77vw8FNIvH2nttLvznHmJeTwXkY/F8M7acSWBnCk5mL
K00fStEY/62fHWG+5jfFHvn+oL/nMFZmSyzwBEhjt4aClOHVgk+UDP9P3Qes9KcT
5uECa8wiUmXCcj9aJp083pIh5cgSO4EQzAyuDntV34i5kITczwJWTlxZwRwO5z/G
4CWg/NvSOYYje9tCOF2rQgBn1g6GwndEz3wCD4xgpArtSVYKxIlLjGCJ+VrY4iVK
4P2E1OvFvOXP97ECHFSzCb3H58FIGJYHtnxK4dfsYdH6fFvi+J6Zmrzj0i0tz5TV
uDHp5Q2s0K4eLl+oMwwdKwSxaeBDOXzwUebuin/6j+dmMJLtyMb6eGsBT+5bhjm9
qZMUAVH2glEDJG/ox/wor/TD2DEbjP+OMkdY4DaZvvTY7ynCC0YItBFn1DYQzsZM
1bf1L/SOltNoCrTBSolv9rOtn8VIOhBGkZdbDxsX97EtjB+fty/vsLjbsZHXrcAN
PMkefJcuXo005LF1G94/Ya/+4KDpb4FEkoynjPiSxzIIkzHZz3CZD+Y8W8RjcYqM
C8u7A1hpSQTdz614+Rg9PdKvMXA6xJinJ8xwysaT9spkBMrcdBL8/ml+0f1SsjUM
oMilMOYC4PjRAi8iCqGVPi2xv0ScLVhdmNYWKZS1uBlggpR0+I4GcodteUI4lKjq
cYfcf67+EFcY74JK09ygQMRWNi2tXvlPxadsx6Y36zSapms8yzzJTPmLXLZPyGFc
ECY4xVYG5iFL6vX+iB6dFV656JNrVbSrY38O78DCsaXl3F8pee4Zxc8Wx4ZJ1uHD
hpmRPOFtBa2Fdd39kD/N/FM8gHjVSdCobXg8STLo8tZmWULYxSTShSCBviYPS4st
dNvaZJA6MaOrU2NTNhptzBV0/5AvJbIdz9a8h+lPHAnqBdj7ZpFxrwJSIVTjkAki
QR9N65b+MnVmQqSIPR66bADbXWIeff+eeW0hedXc989N7MAQTLAOpmO7s4/z5PzI
eTzA5Er0UoU9jqAycfIWrLaP3mOZO4ueqG2iwWfAxngaCflPO7rv6azCbGG3Z7Pd
Z797Va01A4y/bNgKUmLMnduWqTU00liug5yDj6uUKURRfOam3WPr9zWx4ohkjmNM
J1AETt5m9gkG5cbRNAIzYuHUELImTeQsqYuMs5s0ni00bkunns8LTjQ0Vq20ROfn
VIzFC9OONp4s5iJd2uglbWNuI0SCpi+Edh6l5VKDG3DA3txkuaPr4KAGnZ7wd3Zg
IDaoV+qq4QEEdKYh+BdCOLOCIe5AWqtHtie18fkfGbGhRJwER7/YEpFC/LZeeK21
o8nbdsZpCghVsIzhldJe7aH1McQQFjkALD7j64qFUPyOPF+pz1Mnbr5PJyzq0Wnx
WWAY8UUAOzO+Sqh/yXByIfpm/T4Y5KfA4jrFrIFhrKmTgMQEztCQhlmW1Yvi6Ycr
sZ2+0dpjgt0h91g4fVRyD4lzKhN2BlnuMlXrI1h+Olk1FWj2zz/PFwyj+a1Ku5cB
+zR6uriDtoY4bqFT7SK0LCLVVbQSRZZCqo1/5+WJPQkpQ6H65yeNf4zWT86EMOAf
BBgG2sOm7GkspXcqxSdDs6LVZuUxBOJzHpOBq4BwB+/RRLLZRUE57hsPcnVrP3hE
EJa8ayPOLObM0ePwTLa9zgoadsSaH/afvIKDiV+riOmG3eHEGUiLA2kTY0Do/eT1
673s+sgPRVDbKGAzbOx4/JQaXE9GQHVxlmkKFU0scvjJm4UyDr1uLdRRsg9F3jYI
EncG3nWUBrMec4/JJfrb+xUAYzAu4qFcv6lPZ6fEYgYSxAGYMUE5SdrpVvBa6p7J
elclQ0050P18cihtLss5qT1ENjguCjgp0kr9FIBpqLuYN9k9Eu7zdGRy6rIwxGdm
j9vDAzCwI4hI4MW4tkPu0MrVtvAtBWrnCwO49wBtIY1oZ6cVoY30zfdj9r9NTKZV
csiWv/dO/lI+9vLyf27+0WDmTR5D+XLtJcbHKxU3cI2ANi7GjuEsoZ7Uik0jbrL2
hB/ZsJKQUSyKSWU2amHB1gI5Z1Qyi+uxp2yuqAnSJrfZ18TKgffPmKVqx462ts3I
5f5b7sCN2EERFQ9fdzqj2nuwi7vKxJwv2NNP4XQY828UEDqbRvBwaWJZmMAzUQsH
tqQXmDWKAaeNPv7GAsE5gl94gwffXWsRvRmE8m6sLppA+ZKrIAUFeYc7CPG9h69i
qNzbFmCwDVQLF5+McFFpM7ECNcvBX+hiOmg+91jJ0UEOVIqMxP23rmDHWFsdRb8a
7KfEdogLuXgghLtPkl/cVwmaPDxQEam0P086rM3fq7xmYKOjcfI2Tx7XQZoyG4go
bZZcGY1CwfTpbtOkskayMIhehoJAQQU5sIA0k/Op5xfZiH3boocKqJzSXFwN0Xs1
H4eevEUc48qym4x+hX0DbEvD0s2xhigWEXk4BVmYKJMKGgKn8nzBPSGu1hnTUjyS
mC9dxz31sGXqAhR6Qpcm5zW4BpFKhoCFo4cbHVaI4Mg+iQm+a0CCdRhIVfCcPHRc
QFUx17mOfsfxCigqG2mFUAITh6PAJpDW4+mS4sBvVv/Lgj+h7WFA4iTLxponqonI
q9MHrxFgZtTXeUHonRwGv88m7QcwDMJHvBZKeEEsQkixLTjrriBU3Levrs7S843r
v+MZhRoj6kojMOU9o+/zr/LP+52gRwYppHyXqqQ6gVyPOBbOLQQ1i6rYkSNEhKXd
gMT/VcSHaSu6zFM6bzgB+e8eq+cvSGwRs0/0CMTKiJZZ1nnJU9PwEVm8yB6QhS4T
/ou6TObElymY+7ageHM+YxijiIysZ92kTobmCiS6VC96PQ3iIP8sF/ozGAQ+DyhS
XthlJUWEkgVBwqcL0nXF4P2UAyxUo9qre3fU7MU/lvuCRPwrLU8TUykhvGRsXsti
xOlnmD5yAxQHikHj6GRbIsHH0CyZZR+5K3pBOirogElFV6bH/F5zWy7UftkYY1QD
xmQ1vLoxy0a77z4ufBaHACFDDbgF+XiexUp+bKwbRWEJBA6ghVslJc8l6/46jbqt
dR1hWvvwut4uvfzYaWAGW5brgUeTNrAFA/k0ADfv7Sb2h5lNyp1B3zWxceCOBnzb
HK63MhayQUEeF6WHp9IiZkn5Yqiob56OxsOP1YVWR2XFPboMltV39my/4dyA6/xN
E/22ecbWsMCCnzsDK9EGA5Q18JEfsF8QhxwKedrU3aIpd9z8Ih+X6E0LmvWYHxxI
PBJ0aZ8RhqUAssOtZR9H4oExEc2IcGY6UOC+Fhz893xDMp4MuJUf/C6mpUG8KkYZ
SIczDtJqsHHJFc5HKbznQj1650x7cLiphrKPsJJFD0ZJ+cz9NylQBBtA0NR5+Q3D
lEQBDoOzsWbrCNxEorHeS0EJ2fp69HeLc3FBd/TY0Bhj6upTeZAXU2BfKaQ63+Hs
V3Qat4Gn5B+7zlKY3RuTtC1yfG12ApAq3RrYfe+kB0LxJtuRaR65RXooH6OliC2L
WjGWQFcADJQEhsqaPF3Q39zU4YX3En3qZsVi2wJv8zHgQxdkM51qKm2f8V264aJK
+VcWdRKIBHI9O3o/CuPTC5d5gWzv4blchq26QHOqH90Ekf0nKlwHAiuHGl7zvgqw
GAD1nUnWs7cENhjjQV9ItB0LfJXnyDF4Q3h15MKYi93Sr3mmcaTIxGpsalDHz8tp
W6EIvIYgC8HfRHeOezEDZ3cJy3nTrfcjdX60pM6Yxa+JGxz17SjrCrY2mYONNRqO
UM5yWbYYqUFULXZcMbch1yqeS8ZWd8RAmxlCGP6e3zh54pcIbSXUjPyCWfg57HLB
IqtwEoKG3eW9E4FjRmQJlRWRrymnCotCd6jqqbT+3Qq1jVd/CpZc5uzTayYhqt/s
Zz9PqiCj+OzK3SWUeW2QVi9J2SmC8IlgwkEsrqKTDiVyPxj2nEmSvRrGyIH6AVWQ
ohDcPsU6AwxIkq8JuCA4DvyuVMn/GHNeOiuvo2jFawdw9vBWNiFPzwwsh/wKmhO2
oLUkB3ZEF1axwMUX1olWXu/Mno2+Pq1WobZk3cPAVPvJNHmZXHiKPIWe6c0Q3sgG
tRa6Sn7gFhaVjFcJ6Yvpjs378D5yufSTs4lDcgTu7ZiCeHIquEXASYGb103shG31
+88YkGlLPb5Ql/75q4ukiLOm/EyS3v2+pSPcx1elVQYdDELuXZkCkiMniB4+NXCg
1oY4pTGvckBSg0gDZ1lj3axwWkyH8PMN7nSbfMWvGa1H27ri62uwkdYDtfApKBUV
T9UyKmaIzJSxxR/UxJCeFVCeTsBxl+PBOU4B7z0Ag8/8pjxZDdeeUi5081t1Nitf
jXqDmsY1wph1OmCfXGrh9K06e6AP+5DowFirxejb2zB2SGWY8DhftjdNGmCrmREU
wWBFsI7P6mRpquda8iH5BJTuPQYClH404/kG8oQHnJ2rDpcI9rAR/7cCpV9oc3Zb
oKPldtrhvpMsdiJ0ANTPHyXFPURDQanlVKgcAGMdVEEPa5zVWmaNFFsf77+w2/4v
s1K6sQOI3ehRmAU1yFUcOwvK8uxvi7Fv8NWF5PuxPT2nVNo6cjFBjItgNEm32ilh
CG3Z4j3ybcv4DJorPFyuO7aI1/XjLarOlyYdEGWk7z/hr/K9cPPY0ACJ1L3L+DeS
qC0I7rwyXYiKZdn2J2HZCE8ca/KOPtMj6VxOLqC97qQuXV7+KhENyKBgat7q2eQe
cTE0A8NYSdPIeV1KQJIggXlVY1N1Mh6fwO3kiHiNLODU0yUeUXJrwOtJ9JrsyNIQ
txoa9vCzwfVDnSDpF96F2mM9k9BuSLUIL6G+asuhlLqm5XrW7gLMxgMNlLHA/6C1
f8j27acSvqILs3cNu6D1DUagaTXgeUz/UiM7TK6wNNovyAq3b4PMMcS6+nUJOWN9
4uhB9fNOQPAHkXba6pdPRaw6o0uXmOaYXAR2+AW7sPlF18vRQCcT8M4cpYzCSrmM
QNsoDYd5oCZkOkBODu9BH2P3mxKaM/VEvO3uh6657Mfw9P6Z9ZcjnQbGKRPoRk8r
6qOlTASgw7hngCYn0mAU1Y3DyJfsV5VN03oX9DzahkJ9q1XzdTbnHjIzulRNQD16
AFy+cedf6kdgyPlQgGgVmRjGM/oIFrXtzTt0mrw7WlwxrYC2jxgpyDM14Au++G49
jI3an1K0ZUvJLYO2EkuAH9Tch+G3wZp6ShiW6gC1gR4eOBAjIUxIChSeX0Y5IIVS
t6z6gyTxtAu5O0xQivVOytAjahAD4wxzQbFpg1gjzXBd+YEJe7YlVVHrSDg0gp4d
6n+5C0ATVSBI0ZDNwPiNKUg0PGz1tREobwGqJxG+tGzZ5gHZrlXZ0OEB988KTw0U
g1gbKaWNkHUp7IvDZIHPB7Lhb8/pUJnBbEzJnRueFtAJU4jyjxUx6HyFGIircm6R
w663Dsij8tCHIVYkZzmtrsPJXB458P+1nr3cVgN/mC6dR8kSu1xPsFepgeHkleM7
63MY3do8Y8YTZzoQst5nqHipyqh7dve2vm6n/7u/NRlhobUv/U45+YQpKHh0JqTf
cPtAWx08X7h5mr0hxZzuyFHth8fzYQS2esmnt7W2ZOcmJWwNKREJPcPLCw/Lx5Py
7K3PHysd5nnLr9rh5z7C9yxY0KSe7u6HUVBgLFTeZN/HuzptxUCiLRBn3WWnHC8y
2YUExuJ+cum7VDBHFpahrPQ9xKKJj07z1xnxI2v7m44cYGM+TWGpvYlGyVP672vV
eUf/60Efnt3jSjjVahrZSQ6KPyPlE5k5MCGFfSV5Vi0GlKb2Sx0MWvuj0hxrzXhi
usuXc1iozuAqniJWAcmJ9A6ud8LIgVQxddfhlJv2J9IDiPuBOYMicGj/nAL5mx9s
nZE+fY4mKohjhdXtyss8C4NMSMK5F8t0BOCtU0l4Fo0XZHjVsUSGkiXV1snWDGYZ
N4zP//mGN9+/HFCK2mwzshceMBCfHqcKz3LkRQLpCn79L6ei3Y2YSPPqUZufAA/1
xCFsn1O7vmGdEzOahYxGJpOOqonukDKGAJ29v1Up9owzZWK35Ho1SjQg/wa6Eiso
XA45+bX8LKuL/uVHkUObif0YasUYamr/wkiV4urpWb5lEdN9TlW7veZb02/5LBqa
HDlT68wN1y3LVM0H90pVT56AeHeImVTiElZfFAXDpyAGAeXedIm6Ff7Q5/h5rphi
zkfe9ItjYHb/o6yKAxF3vD9SKGVDEDd1Mjt3cYIzeooag07C6tPWqZ6qM+K6AlKX
zaBiY5H0viP/66otljQo0wQinCEGllKcJQ32F4oI35ZDFOZ7niDKbgST1qm0kOCP
2HCMNG1kmANFmyVjkLcJAF6PqWY5twchbF593ljxYl+B78+GSePwz5So3Ofrgm+7
hlhlQzxhfo/Cc47QRyJ/ievfaf3n+pl1Z9biRc/2I5S9Hl1tbEqSJ3ZrJAFIYdbr
zI7q+c2TThy2IsmntnqBmZmsmrWTViWt2S+74iKvRhkAqH1koevlD1LZTxx1Yg/i
9TpZTZUWnEkbC6O2WYW88/hF1bBnx0e0hxy3WmOmuxetv1ryhfm7Vim9rmG26tBi
Fm+9rlZgGHqKAUw/GVG6KUuUSXYWybs5uD0yUOriq7C4vwiLAYikJ8nRn5KCBMqU
R2SNBp7sgfE7Y36nLamGC0dJbChVYmzvO7eYJhOqyNHKCcUkyQhbMJ251VhLs3xX
KDRvzUdFQpQvK+vWBMWVgT4vilCtfFZXeERFOhOSFJFmJlG1t+v4bruhKq4fR9xv
HRoCUvcVGW+DdzWoWZRHJBbScGn3BJ64ISjmTrSnLJiA9DxLH8mq7508I38F7rUb
nEsGl/TXet+dPNyll6VfidU2r8sP/uPsaDhyfec3/oY3YryjMFg1RMfUll6UuGjh
bOXYSewmSgXSZ0KMzSxY4WsHDaMwz6UT/nzaw7vIq6LARApxsUiPrOsYwRfw18xl
7aMziIED1Zg5Qw9YUqK7WPaQUlXgU6S+vop7tCQ9mwTY1bYZuA/uf9lmBDvDbkSd
YnEsD/3onUOnJ/tJsgpnWZ0rhkgGnGKHRYOnN5iJuoILIgFP3hgfYhZjQ9MJNucO
R+Qfu1F9QRoT0bQ/jNy6B5sYY0SswCvSChxRHJxwPU+z8l4Iu8jdBalf0cVzUyxh
3kphdoDoHgWpqNrvZzpRIdE0syjuuMAJpFTEN5h97bPm3Wr9/C/RkQru+KqgjIBS
02ZrDqaFE3H1Pm2e04IyTMsu5A4roO8jbonf3PC/UO9Jj2RzmkDLCdIrlZ3pyysH
XoOLgYLvO00sdKhYT+FSDy/C9KEHBw9E20A5EAEFIoFdWPHiYd/DM0oC2VKRCqZ1
HnaMZzBl6/KsXCg6Vppva47f5CKkB2E9rOPuOq5clchhhra1tk5/ytTsOPMwk3Ed
Z3Kyv5OPpHGBs0TYQod1dn9YTx54U9FJqQ47/naEG+RB5cPp9pC+x+WkLOGxeKo6
+fz6GAlChnjBiyArWF58K0GpRQi7aLApl+qQAJAKk9mjIQBbuNaUSr/ISmDBXVgy
CWvjUoKtuLFsIuQOclzJCi6itvCSPQhXGDCGIkYfc44gPU8lrnqnhqpg2/3Fr7d0
NdMCjI25tWFpmF6AhhU1jpyeOP/dMDq4Tg1O8lkOAuBHHQ3vOCbRZCjvcPYBsdX6
HotNJfQebzKVr5DnKtV5kKsDMImhFOcUnxj9F919jpgj+Lcc5N2oTD11XCLtkdPo
ayJXAIlfq2dfGzimd8DsEVLSoxmtuZPIR11bYWx4nmRa9bWtuH3Js8+wTYHztqHx
8XbNdvm9+1IeTdGsBDj3TKAF4mj2idOAXGZcMUppcHdVtMsyizA+GB5WeO4iLP9N
ZQ0FoaT1p4qsJxQqmurfr9cA4X9iJeaJiBCTV10HKV9ok6uGm7Iofi1VnuxUteMp
B5eiSvheKgVdQ43UN9+XSEWN3lUpu8ZqUoxJg62qWWA9QerKncf7/ONI1l7eHYLZ
mIXnOS83bZsomicb0D312BrimZBcQhlDZpoUAsRnMqQRQJCj+8lWXQ9P0DofYW3S
HtJJCwpAzrWejneW3e5ekFFPE9m1JyLgRGqtkjmSBoYIUhnPr7LeIrfff+bwtrsY
eguUfVA7Tw+OtDj2ylWTut15JnC/w01AfAnOc3WXOs0eCqhq9IkpoS0D5vi52EqW
sj6Kqbty338jknXk04h27oSY6+09hBf3aPL6U0Ndhq9i3ZvqbF570/BEorc9pX+S
tGromB0lEExnNrNxulibHtSjN3is0iYegcAyQ4AGq2B4DgBULFVnUlmkK9EWt4RX
bcpPUJM5fFRA7Jdw38nH26SlSdL8HUNAkxBWvUc3SU+h6l1ozpzJXxB7g21lwrdQ
horS0hhiV/lpqEGZ0KhK54ZH4ycvsPxFKM2Cbm1E4st1VaP30EnwQKbtxNl6Ka1x
9+2Hh1Wezt6FcqioVv7JJAoDTFtK+baeU+olc6lhL8Xf0CAN7EHKhIsgw6kwJBe4
g0UMA8J2rxtWLafBo9H6hzmUyR8EuQvMn+N9apgdc19Lg44tTpxU0wlvLEyt3MlV
TbTQwJ395uCLPZYyQR0kwDdYr2bpJXUnvS8vXnvhO3T69Utc9mDjO5/0l6wb7WFS
u5/zWZDzCynK3sZNlvNcXRd7eVIS2J1tC8TAAHeWiEuI77isumUeBBrYpacm7OCM
FAoTaxOR6cuYC7k5YkjVjY35++ekeQYkRumc9I5hmY9v77qA+63ZlIl6EYjRZukf
eEc9HiI4H6qyzRXA64/ISwuuAEFS9CF54ULClyOtkzydt9vnIIPnzHhstoBDeslV
n7syKS+FvScbCWgbQs/c7aMbfvITXhOBaEA+VptpYQY+18OOzn/CQOpERVKIyyvd
lAU0dLAa99nK+1qoUlmdIyPpkcWl808pBrgQ0VGfAHn2tW5atlEgPKlxMNnyk1I7
5jzKTYkSGNntfS0JLwgheIKjlbAL1FRkem4oF+My0eA27MmoitYFmVQuy1ng1leX
zWVsP9WQtLBsoKzwFYoak6pj3VZIAJ2qi4+ZtiK/5Da+Xh2mOpqF5iKGnK9s7jsG
ssE4plJ1V227wk0GKVAcvGSwUY98gRhlgcUaJlttDH/GdO+jYxq3IgCaE7Hx2vGX
sdlV56/WVAUDS803HExerRHIACFZdH20L9MRCh9caloTYEc0NCm+0yu+VckLj1Pq
ABWspKLok9rkgqSTsMPnxeQU8ghodHrgrTzMZuyPCStHYTcfmiFIyKlDdVPlXkKf
WmV3GKLOZbtPutXBV898ViukcErQaFld+gAKUVqXjMNbGvyyQlasdHvibLxdJy5+
oq/RgYBlFPJdb5B3XorS+hseww1WlrX+LlHgW4H9q2pKERzLznzOSlO3LpbIpBrC
16MKF9bqGevDtLmSk3lgt1MmBTZirD1OUECJR9xULDmb2I6oacoN8F9Ix9JnUUGk
Hzfm7By2f2ZcXgZFFew1mAoFE72yrg82lKGnASIqd1YtSQlmO27KEmtEXuuU9d6O
qtJQsiBf7vDKqm8i7axAOghM5zrLE+fZRHJAnykKACfm/+X4UmsgQI86xXBo7UTJ
T/oI4TJ/g7OCg/5UwADVEB6/zTvVYuxK//h/Th3r3NCkcdO8d4zvVQ+XAm6H8FuX
k/+RvCcAN8+erMoPHL5Uun8N4GChuMna0zX/yRFtBEYWLUUYPymiJgK8qZwQvxzM
JF2CisLBBaoKY4zjio209BvjiJVXrnoh+vT5s4nSdKxMDXwXR09GD0nbqir6gYtw
O9i9bQghBCbriHJwUALZ2E4wKu7/cG6aJt2SUezVXlgWNPQbV1Ny6B/AGsv6rRNK
/a/43i0Z9/BkS8wlTvgWIbDgyH1PoJYy0aMQX0zorqujLEcbLTp02C5p7fEARhdK
EWpcOAaTGlV3Uy8YCl4NxOHDpy94qE9tfVRcw48MygpwKCT38nSSBBVTmZTzylAr
qpKt/5YEwySz0fJ3vShU6qR3/3q//YcBecIpytgAuR70+OZ4c9Mnw+N+gxBS48nt
UkJ+A/mZ/nHxwNe5sFSna/tye67QfPU4JfLAbKw4BeHoa2Hlm4//tLMHRVDVO5HI
d1xCvpi2bM6RfiW7dTqXEAnG+1Fk7aYLRk9JEgi5ysfUbzNNHgSMSU8uHUSA/c8Q
3dgi/fJOc3OlyteYT3I8xs/F9zSO3lYQIKj/eBwjbLjsjgTra/He2i3u23tGlRXQ
06o/eoWzaCCFHkodYFHQuZztLUjJuLEFo2C3yS/IOW88feTaAOqbHexNJLw+e4Dk
VCT5l0dAMc3mUAO4+ex3c1l+ETtRXmLCCGZBIGSjE0nZAIH3CuaozbYcxM3G2yry
32xs12qscxOYvN3P6c3dAhCUmVtWqbB8V602b6ZIyt60yiHx3SFL5rkOPeRZP9ms
sQhVJILc0hdIUATSjKo8iDPeK0uXi/APGi82nForL3RD9Qd1im49DFbx2ytozA48
a0x6QT5aCAHneDw3uVduhhN966Q3nSnS8uxqf6zDSHKDmL5F1LbzODmmLHcl9C6k
7hGrMRzmIzr7cqULpE4O/7/XN/l/Ajg958MA7GLnqgVTBYkT5CgV69R9+WJTSYGn
SkPlVrH4klQTlimGC9mUGXiK5aJLER9c+OWTpcwBH5ms+vYbtfagkf6iNs1y3nkv
7L03wzx8mSpSlLcsrjSecUwYs1HfMGIqiSXvSC26zz1pKnMgMJHKRMmz3pBNCVto
ml3MSdsPXoICd2xhcGqH1rRJLJbmZkRLsGEISbJr/o/C/PJYUXgRysskY2H4S6lF
avRfd/s1vhJnJgJXbjwf+Eo8sWltaVNpHt1FCJI1qtjVMYR6kFmMTNpCsGTM3aC1
rSh17AcvhFJfNmmxRJ0PLAB87C8i1SLd/TpowVDD4fK8bpBYZ3AEM7CTL4O+KqP3
xBmaZZQxhLHqVyxDw9NVAo7gZbrJ1U6TwRElgSx3RbfFE22Nbg4lTYcjMrmXGDu7
LjU/jhnS1tjCAQC4lKKpei563BatnYZiB6jp4fn8zMUB1yxsf0UQeW1+SzOHJcOt
lj8w0Ki7zjZKTOHDDTUvGnPg3F80nxbUvL1sQs3IiTcXrQDNdVxwdaGioMjwMLdZ
+5NBFc8grDru7wUAiyF0GeaSOR+VUZQBShxnwVeV0m7wnFNZGRYPnvgF9UK6rTQw
NhHMVRwo8VVn5/utBBSKb5M8nPejBEtO5spVTK4DvYiI5rZtuDreLWFVShl94bf5
ulsupa8LecXv0Us24sooFZli02tG2CRvTyJ38EInrh3F+u5bg2cbg/ZptzbjCH+c
S6/Cu6kCtD7Ds0N1yrgNr2kDx62gQaytTnagi0lVG5XXwrDash9BofDhYcbEAUoE
IWVpLxYbPOeS3PUq5n0kxdROo+2vPlMpRQp89/XX6z1Ozr3FqqrWnDQGvg84T3A6
AljCVKHul/C5ct5oazv5WD6FysDRqkxL/3nje95hWtMp0dBh7APQa+X2Ym30bMgz
nXSYrCyAccLlaXxDzwlScMX9fqo36XXLgB5fmdrF0FkIxLfFgf8F3UQkp8uNAjoZ
51CCr7xLbt23xriQXR+XhWxEjkhfJzHQDDiLF++9BOZLAlagegB3Go3W9qUhRh8j
zVGnI56+AO0ufr1ZSpRNirPttE3z37eKQcsW7IoekpK1J4pHGydtVj9kNBbuSDGA
W3AMGaEvmWj1OUB+G3vfgavmn4nUgMTz06/kVkjjkUQG84lojTAfn/IAv+RvQ1F2
EcafVBTgEqFqeyu8FtwiX2kpMaH/or+klTJUSyD9WD81A6CQKvIaBNxN37UpArbB
ldioIo48EufmHx+EaP+YrRyHjJUQLjQ2v0RTkXpp7/7Ru2Z/3+vLgjGDpv2Lz/rj
o4JbWzmvr8VyEKhpuzZGSTR6X4HETXX35+SX6+YgMSRVMiYzubTdd6gsaZRiDIeP
4lwbjLPY01yasuInpGMO1hzM/OEhBdpB2zHEk2jYHhRJ2BuPLx4bVI9+rTXpqDI6
33FzFcMEi2dov/l46Lo5nYXskZBggDuy+GHdnDNXDYniYyIn2D/QO8oF+YlQIOZA
W7XGHTJoN/vDOk6mierewpkiPgSsHM+c5c5NJUYxvClXwuR6FWB1SB1X9G2U8sx+
hCaVPCTcezn3+DdMa3mx+k5qgfJJg48a+wPbq3ZBvV3tNtObBYejynKo5WR2oHXL
z7AwHg4Wg1mXwSDhUpcfQaRis2ZQUXoE0z+JTSXTUH9EuPELuGjCfpfKh6Wd3lX+
L8+UqiXmWRtR+/36us2on3dC+WWyYD7HzBitC1pP96Tb1ZHhk88Y3DqLk5/zOBkL
qnZwI7EuPrfFy+wFcVIx7EhX2XgRPukeKwlsfqhGmm9HJ1IWICnBMQljvU4/bi5k
tyhmB6GhXTRJoQEv0Qjuq2W7+lXiddsB//dNl6NDE2YokiW6WZDxf3wMoL/vXgah
wun4NrP9IgolGQrUnPPsrfpxR4mrJgV6depqCZNhTB2MB1dcI9KKAb9KTMDceOD6
onxkcFvPKq5iDqi3qSBJiKB7wXSxpgR9pwWgSSOljemv8TsX9g3q1hkasM7dnDVV
4nJPpcrFolr7Cx48Kp9ej/hQD6BdcrrhpF1nCVUT+Dfru+yGVkWrexH3b3IBRi8H
WeQPbwwzJbWg8IzsCYX7bqNxHljVh7X8XbYr2FedLSayssszxf/VYY+sxfDmiNZD
Swv2n8lXIINW8w1DJsD9AsXmXkj3klN77zJOuEXkk2Ke5GgGEX0XMMCGQA4xIKNp
vfPTAwam4Gu8qoeh+utmgEKbBSNCtR3WTaunrjEx2WCK1GJ6Ye9EIShoxe2LTcu8
BmF9LsqKE3Rwwd+5+3wV5K9LYjwAZl+eRjbHxpz6DWKFY1c9nJrYwfx8gIYHF06q
cT+WE5celQvv8CBGY7gO4kErAyicQc13bclsT3C4Ntjry/Po2454KMx8C6NDCWhs
HRf5tIgtUF5n27k9jHbibeRYjDrQZ8rQ1fGIE/8uE/yy1qvpcKHK5tedHr/4FASv
4oDKEzSkeXjDG8xHQyDU7CNFueW9DylN6A8/4j0pMVXOiCVSgbzl97ObXL9Zx3VY
OzAh543mKeTVZ3KH0Hgbow==
`pragma protect end_protected
