// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aP/K+guTbXPEBquFRCmNr8nYGNj1JG3g9O57o31uvPlwMYSyunH1dj+wIVJq+CoU
iGB4MkHTBMHBnugrV9rBhRpXVvqfyvPr+louPQIww10fsdEd4AWntZ0UBhE1+a+v
gZC0O6Cmt7gA1d5KHzycE5NJaOT7ll5gV8/fLs+54vQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 45200)
I/LW9he5yFGik/5dzZryBKUURHbStZBu/Wii+hOqDrHK8fCqw6XFqAGQv8N8KP4d
WEJOMYWX5FrnZC3MeTij727ktx6MI1MQzXe1OOcKbFOasPqW0FuQSNDJxWIsyxuJ
4SWTowdlJK6enxaujuhSZMnQMDqZ5Y4OUUZU5omH6W80UgWjepmKUtl8Bt6wmCLw
TN/IuEtB9d+0lmbMRAAML48vHsw84ZULJeGmwjMzAKq0JZoKRFZ4lPC5W2Z0Wc+h
PJEu1K4NoQAuJyiSEMnmB45Z5zYNTTYg6OfXoY35ItH5d05trvk+ZddkTV88wx54
BcJVcs8sB2kolw3orEqLXa3eVDsGrWAPuZSy8DnFUTJ5RVSDLrtHaUkAkEI771YP
5u0CEXCsqkLwIMO7QRyfvKVTrBg7wPuRmU4GGYQ+9huYxXhyTg1ynz8DTUlkzmS9
uf4MfF65PNJ7PILuu6qKl/pEsEHNhKX1n60Ej7+pGVMZ98VYKjYmVpA1o6atdGoW
n2xQzMF+4jVBE80z8HI1juPJdA90wpSQ5j8zJhXoD8vwU+o1BBbAlS9lMDMqIErS
cS0sGvKMcGndPM9Zij+5GcOy1rnId06coGhIvoxONBPq9NdJxUhII9oR6chxNFZS
O2PIo5rDtxAH9DxKFKix4lMQOAFpwi3RcTgCyD8ZsU2uCeg0JIUYN29h+psIdQfF
y/fce1htubtaqi/lvPMl5ovMBkpKwECSVCEce4jDZ7tNQf4zpghf/nrvLSJrZ/1k
0xI5emRsM/OqWHabtlwQZb6aaKF9UNqN3h9Ead2YBwChT3n1Igy8r3A844qr77ai
fKwohOonbeaixdMkQYVxIDNolTzYkj4AAYlR5xIdiVd7j/HvfcHgVIr8RkytiP3/
xIVJvX/Di5igSDNccFv/pMhHngJNBcLnJqGMSJ2z+LT+8zgxRrBVik6yr5CzUoC9
XTGNRnYGYJMLNLvdmydViuLKVlF7cs/A5pemJVzeXJzZ5RlLnXUfOhPZqTHdFbM8
xRRHOKn/e3YokjYKv20RTphRiW2hdHXVVwNOy0L10MVNVgwSfLWp9eH3u5E9a5CO
H+t8Rr0y4Fxvd9pRONCGyB5F2ETqTVfYvQGVQvKc+y626SN9sQXn/SXb3DDU0pll
6dYwJ8Vs2naHfu/kWIE/DaRahIPU0hi9TE008k8CWKH9qIN1QVoQrlr+jCEeAyzz
aeOCw49Dc45OD2OpW248vrY+z4jp2CM4ExU7FGnYTLHTXlwwB405+t1fwj8QBu28
E350zKeumbmjEXNltUe4VnZ1xHXGQ/qeaRqzN7szH/mUJ/vg2xzi8CaslcZ4a9H3
h4gG5sAXSlt/Ynrf+qpJcRsifSBOCMtcbkkcuMwMXaZcZSldRYVVp5IHyBufD9yQ
+0tyOkRUi2o2CbwpM1ph4TyO6OpM67jT9xh/76q7jL2OLyU2GrJRwTcyBXFV8fBK
athWr+8m9depfE5iyHjDWqjCEtG3/GDCL9A4kyI1rNeyFZhA22hfeTOQtA/X+lbr
QN2ijSdUgw32/s+mv3SnyIBAuJ4/m675IK4p3Mfb4Yyaf/TkSGpol1rDwIT2s6k+
DRaVRZOz56juumRcPrBJ2yczZLtAA8F6mytczXHFeyIBU++T2H3LBRUwmhpLX2Eu
Cftw8X3w+xP9RcnwXUCYCZDPUT82tyGq4ytJmqI5vvkQfVZaddP/B8gm8LfeS5+m
ERqzDFjiGNWx74SsPrz8YHIBjjiw8iZA/TgjgSOQAaoMQOwP0idR6COIPFTt/xFk
N9pWwKg7vz4l7dBPaZTtCSB8fPYNxBfTQvSHKqvIfYGoIerstdo1e19ZgnenVcP7
f/4UZVZqeC2VHeFPYASKktvelQcEm9IRGMexy2+0ZfoDF3QsArs+LoMvYxeGe1f5
54a4VLESXpdS9B7GKPL4vImMmARp19sqFkhjlCyyLBPo+zBBFb+jsqcfYEbSBBkC
QFOOBdw8vmKvQP+6cxA2DaXRaQVZQOUeV4wEiKy6HBBGgh4nW9/Dfz4bofh3vDpU
4Fuo57OzzbXuY8Can+CPv8jxw3oShkEYowwQMHO8pnh8ceg6DHx/qoqkW6NxnmCV
+TnaxJlII0YZmU99vFd9EQCBTtK9u6s661Z0Im79nPSC+K67Xt4aWIza17liIntS
t+ssX6hK+dk/TKLwvCo61KdRV/Tjev27pZyvx+g9O9LB0Jb31My9kKl0yWdIP/Yw
fLVa3ZXAzC7tVZG01q/9N4F/qRMbgrzZ1+i/x0K7fpfrTz2brFVLovx8OktLW9x1
WeXmdLUhNTXW6I+M+pKIup2PtgeUDhcsmPpgV+stxIcpxfqy6XgWssHB9PeEleiZ
rTdZaoJvNTuqMvT9cnqUIEFG4YkM9X59xFoee/zWh3DNITytQnAF4cazdBtUG/cc
xD9i+4LbCU5uQJ1syqp8FYQngshSCdoeGeHh8kVJOB1s799DY+8wnN8iUhht7SNI
lqfs3S+WUbqxEhBcgEcPoDZz5xGwOZPx1pidAGuJtE559DbGcv0KoYES5KiM3rwk
0i8OU1MhrzFGTK/j5gPwDskYSa3hPoEGIDzc8FPxUq2YWNSLPNeBsExGAVBA7qI0
hQeY7pUZOtw64cY8GY0X3NQ5XgJIwHmuW+v0UyDOIzPO3FZunNQhrJ/QSb92IX4p
nth/WGTmnreBqLB3otLfb7rSRw4aHBrYUTjrXDvskwAaPbHVgC6Q4sE6S7/hoGMf
FDtWNnjJZmURfYyfTK5lud0qOc1+4ysiHAz+z1OyMmuh40knAehIu0t5dz8GyNrq
FUA2Htz7fvsxnQTjFdxU1PaGWdBfzxOHbGuHOrONgWBo0qWlNfSLmjutvfFhy8aL
U28+yzG8KYrEheY2Z7g/rZlBQoswnad0ygLhhJcXnwGq+b/dq2NEAWfoGiAGiZ+O
NeRLM0kVZzGusP2hosgygwnihvpAcL9TvyY+KXq22dyBXCHOchEXc5EFe3lFIKFA
bCxfRuX2sCu+ye7kyeSjnMyf9vjuN9CJlj0dhbwyawAAY92BYDxYi3QLOPeKHdCu
bmx07fq5RHdo4pf3EHnem7RjSk4v0Afhl8YBvi4VTQ7LTT6IjlBD2wAiOhmaOgc+
rU4eETwrzqcx4e8Bmad5lxJJYAkEwvDXTdVBOIs/gF4uImJgbPkCItIsjF+kSpmh
9Fx7y0BsPxPuRPTySfpuvyeL7aMcppqh2Z/J/N2qid8rfQswYBHXZTNxsCKR5NpE
6Pmt50EEmqtAdnMsAphnBxNi/9vQ/eMEhuYLuS9QMn8unWpCWFP+09WPLuVc1ZT6
0zKzMi8mvaB3PVWL9xmdcJjHeRBY4FMtpxLCFrUqrpiLmnbK5eFiGnnu+tdOHAOk
WStIix++ZfH4Q5l1JN/2f5KlMApGygwWJSeKZiaeThgtBjnrsTdcLcipZ8rAfEG9
GQPwEaQmWdDu0Ytx3jbYmfBqFxOMbc47R43cCrtK6qa+SLWWpORMBPNvizJHcoI9
wKkgnGfFtCe77r019N+YKf+8jNwrh4bH6YGwAK6+oCkxbiz+fs6F2TVazDXb7h4b
t5KeZgshsMAtv+rq/S2xwK/F4QKuuHPDxRzj0k0AM1S7PAkzXqf9aTm3hQGklH6G
TlY6+wl2Fc/ODUJvi9LdHFySf0tc+ATJrVbJs/TNu9d5BZZvL1pG7GFdHvx1med4
Fbo/H9hncjMqHgeFHRllatHzsgWKlXuA4Cnbtxt4SEFMhHYt0xQmEnlFw9H8JIWx
dRktozslQZowGOuDHW5QZx+Gtr1dWKOF55iahR+rDNnAHGJ4w8uCe2jm1T0DKCr1
6NuQK5YyQySco3gS3OqG9WpotlENfSCs++Fo2ekc3/VWIqoZeJ18pt7O2PAKVuMs
ztf5qmybI6lBwi/G8nnAi6mxIC/A/MUVFa06Kwyex7BhQJH+e5rjLD3giil1cvqd
4RfU0jyBZSh5XJ4QT6Oae1Hl+IIo/lcBfQKnnp1oTi9M0SVuGqbGDh3SFFrOYNIo
RHEFFKcG0EhDbgs00uWgeu1npcCjFbsSjwsavQ5vhcMaeNgwFpULu0EpdzCoD0DT
9vX5VHiSgdh+rGKiaz+w08xA97NogBLh05p2Pp6+7haSCyJJygOq2BZuJTRzw2tn
7KpfZaI+duLwvJSEbrWjfgKfgLCIhWuyv2Y5c077MxCY964vMROixusLR3iSFl+5
13Z6XP/b4IMx0hOH6SP/WdeqR+p4dWC6YTwZSpKQhzONAzpSDCGY/q7kp6iY63xe
WvJ6S3klEuoCSGOjyvYomPq8V+iZcLYMHSAJOhv/myLu7x6s7v395u1vzYNVZ6V1
BhhLjRXdtNXwF+qh9Lzrsiu8YuZuyJoqa+K+kcTpFbIgYKj4s3S2jcHb7vhoLLuX
AtH0SLU63Z0nBO34N8DtWvpJUL9lpADMME9ND8HlCARj1oT/RVUHkTE0cxLybhg7
N7OTupjnxqdqIk8QRXOFgxAghm81bh5ASUf7mF8ygHfQ6ws/mn+doXGOvnXjQbOL
Fehr4HiTQjtz+AqZx+5HgN6RlXB/mXGBTanBYmd+uY3yZEn72QP9G99fd8iP3CsO
Tg3424Lc45pQdq71QvvQzWsn7gsEDbXQQSkG2cNbbPUssPps/P+WIMNMbnEqItqg
JxIw+jzcA7uvvpyBfqEHmXhVi5XjAgvulLLOwlf37FJ3yZzT2za12SfAxeexmIGO
OKuGBIynXDBTgLphxLa35pOYeqh5PGCHboauHIlyvwBfurw8jm+aSIOXKU4xAaAD
Z1Gk9xQizedCynqYvUkycGCD0mc3Qy1wO8Vf8VGPxcO36ZdPgT9AOi1HTv39Hz5L
44K4whFoBIEIeuQF/rfD6x+tphihEeDuHrTNghvnws8QwDNH8+mnUoNjeBzVWjsd
5z53qJ9y+8oO4d5+QqCzZpCnoncUyj3ws8azIX5CMttRAHR0aaQv60R/Lnc/Z+6p
6SdJzq0w961uiYogGKdRNssYfhhpdeImJfE/tqfO486SMYD5vVMXguBa1QCfhtln
BoeN2yg90DzHeP4C42Gs2dVeJ0YFaZwlrLSnTF9XAqKzBp+xKEk7UDrcHIjld5QJ
LMr1+dAhc+OC5J7xcI7hVZrWq9Al0VrIOtOh613xCsePWEVdzCnJkeFXcej0bspu
gvoPEILQO631lErPD3ncNp+DUH3UGmttJbGU/C+VJp4Eq/0YdfFTBW+nXsowFSJU
3/XKlXrCrrngrI6UpOvs4IDysiYtXuWYuCbFt8R9h8XRVkjiS7ekP8rv5lOrhLqY
g2ibdSwZtU7Jr51sBPDVd97EygFX24xNXkJJLGyrfRR5cfrWwUb38DC1fxUukvbL
PJUfN0u/IQvA4K3F/oQj6F5nbObnfnQCWYV0Os+Pk3MtVWPUXYNOf8mAV61OBCoO
Ibf/myllB61jsH5qMEehvavdY/4kLANc0oshFyDptQxbcWJ4SCY/5PsYVECm3SwT
kHp1HBcXOrGCLCPwH0+94iYj2tR3e3zObkXIxNocmZtw4xdq2I5qR0f0HtGQ2D2E
XtqPxzUsnX/SybHrJC6AnfiaIS/S/8koPvohmvqBXzoV+1Wbw/lLmDou4cjqbFX+
zwVUqZq1VtOTUUwAm89sjoGGyz5Jy8jCzW4f3Eq0U+kGJptSOlDkUHsUfKDQLgPS
ihejhCeE3CZZaNZEeaAn2X7Q3wf47reXdGd8wRq1PaydY7TkWa0rkbHWYlbmGDcp
+IgqZus6jqg30u0ZMsYQVIyCZv5QjrXsSOkXXWXhL5zVBhc34wn2t929PCh8V4d4
llE23gI3onu0ggmE6uYvoWLmYp0vQGHxiNariEABcrN8zfeusmtA7XFehmazZXnV
u9x19iwwo+fmS7lQefLMoQhxib5ZTCwm1mjC15z3plSJNXdOGtxav/ZT54TEPhTK
PZOezk37UzLsmlTNJeEASZD1HQjpo/phSAl098b7QW9F5sWU0ty5Y67cs2paTsDI
HTzYKeDNyMuzpbsEbxfsMMlwcFLvD/aDEavi2hbAzXWX1zRiNKKNxd/29/6IfRTy
RcytNbaTUYGBquYB5DSkNC5h0XwjfSo5wQu2Rsm6GDdflzTf4jfwYKnevUjZo3Sm
+zwWe+a3MZg0m0a0ekE9r44jjlFxpVScvlO+VL+Yt15SRc/uJjh9HDNQEpGzTnhz
K9whPezNxmHbJGgLK7/E+TCwZZ7r2JeAdv25M0gg7OucRS8QuGk3oJ4S/ZdjqrZW
ldi3trdTZzOdA+NctyGSJ4UIiDDb5npcPC1cpBKdh9o6r6765WMSqvVvZElaQfJO
kK1xFyEBAfDU+U6rjblojZgVnNJIuM7rKdDoSMWRdwHLsjBtbZ4yl9I9AORC7SJ2
1hfQOBb8XTqgcMGLZp8n+ymNv2fTZ5vzSiQLb2HSVyZkqCyCqkKchM7xMBx2O/tv
EG70BnjrjiUDhT+HggIF4TBe79QldSZZvXhluSVTb0BF9kXrYp8w+d5/HdRhorF2
kRgIUlxiyAMBFOKqmWSEGnZVPAXbd0D6cE1DtIalRZbHzmWdvbfbW/w8MjYn+lqP
OtFeBUU2Gs7tGj8XyX/QkzXYWFUtzGMd/JVWCRQAlWZ5VafqNEBIq9b8R/5h/rDz
KZGTyxLqsfgE+yRNWYzTpRXqm6I/AZkOYPrG2wEkThTU4IEdJVAfMK6e7iytJh69
D3Gz6FHXcRgvv6hN6VpqLfcoAcidNgogV0UqI6vWBTMn0vLkFSxbUmctHHaucHL1
KhedT72Wk7o+2YmOCh1bRY8bGDhhtpE6voVrFf1xIF0K48YYoa38o8gagReerUYi
wv4A/MB8xPqiBZjzoMnLgEL3JBvuRgkhpejFDufl1dPcSSTnh6bgR+iU9PisyYNg
87dAO/LAtOEqpYS2jgbHVOlyTJfCCMHbQA6hA3SZJf+7dTKcz1LtydsLM2851rSj
eFAbAvrGb5cpfG6qoCeub9LSxp5dzuIN7IRn4JDMxw2rp3O63L9wG1fWl2YHUVTt
Vr060zYTTsoiGvREZaxk5eY9bFdXyo3YMlNkwl8r4Nfxjhk6w/Ch+2AW6J9PjACx
fX5s5b8JOwzGqZF4aQOz+KL7O7vGb5QMh/ugWYM11eMEqBC/H4zEqNN31NgwU8Ur
NkRaN0NEwIa3KIgcpSnkOYIrxV6QFp7JqvIgePUrMpjxDyyIaFO62+We0TWkvL15
nYL6UIxc8dAU9PVPIKz849z6OvZxc5P741kgwb2cml0IDuAzJx2uuJhFuNCE2GHK
Hyyu76mhcZo2hZb15LfAtgSO1bbj7JEgy9sEDtqCzP4SUrDCfWltpoKD+DSBKhwF
rCw6qZavVQRpZr95hLFIRxT1z1U72M9F4R7dhf18FBFqguIsk0vUKbI2NuCC9Elb
pUwQoZt/8JwzaOLWr0LzpHXYhAaKGyuw0kO3wV0sfY6WwvKRNmt7I/8Q9G2T6j6p
gv/WLJl+IDZRXzaaT2g1mPNqIaLsJggg2MQcVYbrGPxJ6H2280qpO9CGPg3s8Ush
CAXWEFtuG1hfDZKa9ROrvXwPJBIEV5UzI1v1sk5lSABdQPzxqRLrmg8SpxNmSsWP
uDzcqKOqEsBtCBgJeK9vdpUi+4BS+SGju980B9Njgq6uSWIqwxkLEBPzdfnWVhX4
bvOPtQBx0EUpoooqsEdkonIbxJ58AO/SDFzl+8NBwnD1TCmv+z/4Oab4cUlwpwG4
tSpNyzg0uRfiE7NsQFoRKu4WQvoPwveGNip62LlKskRO6XlAPDmTgPW0TLy4QBJW
/SzZkBwwdBmE/VYlWsziySQ6QyDor5fmkdzZd0Hfs/7zaz8rYWMbtUcfcWtLx1xA
g1pPX8Y0frG1c5CmZ18B5kXPZzCGqAB426hLAzLG/bFkkMyh42nmTiiraMsVXZXm
Nmm4DEVAyqwPI7BJxPyHRkBL3+R7Yh5E+RdcV2ntY9xU16zQW/d+MtaE+UCrfY1C
z3vXAz5Kb3jmW3ocaJXj1boe6c1X7KhWui/T1EcTgznqyu/+v11B3D3WeE9dEJzo
RNvXaAnirZTuuNYJnVzlE7DGX8zdFcok/97Dc48quu96q3PsYrMxTUplqqZU71BP
d3XjgwTVbJFqOCXiw6nGUewgZa9U/kJTMv/uCTLnOTSxdYUDNRYktzGW/WEOZhDE
YtusAERkiHwgW2fkl0nCGzokB4zWrXXgi4X5LDLAvF/zBFGdtuV1+VNbTRlJf6Kb
JvH+I6NPrQO7Ktg45L1vrsji6BtjPBVx0ONvOzpImNOkEJWHAfMRZW1EMU27q/ml
pN/0R5oH4+x4SU3Djrpi12x20MDFnluBy10a6MMKXGJO/5dFixvwgqbAhh5w1t9Z
pu2AXNic6wH+uoumflMwkK3vNp4bWcMMmfliYf3j7g/rAgd7Cjp0M3p+2ZgeHQ75
IqwcvcGc+xB6RqEpGhVeI/i9lnGeg9yLd04P1/EdR9TCcQFLSLDfRPVC/QQGPoej
69JHqyHcXK78gLej2qSKlbrrgDGa7fi2nEpwcxq+3AON6KRGiPgWxwNnZAdWdp+X
AVZa0lSdf0VHENyRb3u7eOzTzyUcF+q8lWLClgowS/ATUZ9WpUXbCWkXFCyYf+qc
g+l/2BNf0HJ4NUp+q95/Y4u0+IS0I2al5LKRgQgxx3J4HXxFlMuRjjiqVL3VR6Tl
pKp9OyUbb1gizq+082etNvSNiGeVJDqMVihXzsigASl3UvN/vRPB6w3IUiuXjSqO
ChRCiSrJKi8YTUGOugx+xW9KvbwuF22/OkDZ4ebIgPBL/apoPowrfs069A4/ISHq
uGA22/XY5O6DESGNFNxzqHl4se8wqwxAfCK0htV/OzTcxKL2zsj0i8T7biddHWhq
DYZPvzEXzukUncop/fKeQI3Ox9Dc3xunYvPMwEraqTCE3sIr09kb/UUwKEwgrvTI
dbloGMgW5632d6aJ2SFGEXPepN70x89C+6o4wvAaR3heyA+WGzA5dNb0nRxZzir8
gxFM5ZaUU5wbYT4x9onG+MLyp5o0E+yWVt/MpEvlQU2Dqf9czcXn++AjZ3Z2IrfQ
XvRWgB2ngDpWo19m54SvQ3fKExUFhw5MNuVfUXVU9d1MtVvruE2fAciIXGU8Ffck
qs1C19dXcreuZ5oP63LCOPj+mnvup0lwWmgk3kCvf6liJGMZd9zDaLzkTzrvA9Jh
x0aFHYbi//9yZ9oqlsqYuP1H3NABpiqaiJvXktnX3GJV08wypilVNPsvM/c4StNl
m5xOzMQHel5FXFdnjUvy2hjwJaP/yrQAUuKKdYnTIIQGLllXvFGl41P/pyjpdypc
ok4t8ylB93uNY5psvlnHEuCBqpafitmuq8Iv/s6C/5OsW841cEN9T92mf5tlyDDg
+KjYzPkZ9mZSu+UmS/CMNPxK58ydTSFuRxscv5z0VwedpsQb4qnar4uWlb/SQrc0
HbZAcouHBnRQ8GtogPEiS0C/oYMaBJ925IKyEOu6J+qnOIqTmvnrnVSPi9TCTsDi
O4SX1x94g+zRisdQaWV0V1Y9J/Cb0H8RSQ9KF6fJ3YjOYI8GCclUD6mIfraePRZz
bmiU1kbG8jhCBAd6nvMSfyry+BNk7qjxari+iE5ocT/bcFT5B2RHgp/qdQjvpus/
BsCNxXvPztN3w3JvJ3yeOLRZSW/29FlmVZ/kaxmMG7dd6cc+n0BxZoCTdbhOdTqB
V1WxUrRtWeQY9AApSdW1jK5jnDBMsG9gxiHdSA9OxvHGC7kZ6FYo3P1bsWHEMIco
8UrxAeX/WTQzIJl07Tce2erAZfDND3OpG+edcFW3ko1psSxvffoEVP+765ZnnoBQ
2mPAPECTZltxNupluLxmiZKVmpA92JKiPbK1IBokUzXm8WTobNVVVCRjglpizvKc
5D+EyAwOOWfXsJopZQ0rxbziirRA6tkrcwFanBZPrTFEzY3wDDGjz2iMCOKDND9s
iZqrBn0m1fIStuIW2pcLWisILf9qzkAvNvG5Ypcr7qys4V1fx0hHhw6/aCQ+ckJV
0dOG7+uJwl2QxAj0rJvUMFQAdCbKSHxBybxjEefhafcZYro/MW7g2Jus3TUr4OfX
lyi8tfpf4HZmkUU+ey12IjwAJfJKBlp9bE5r1yoEilmmFFJ975Q9tamFB/ELGOBR
rlWjjAOEyLSgoPK147bmDmzELM52nxnNdrVqnP9lZisYaXbSqAL2yYzfzfS3bGcJ
2FpLxPVU9FbBjAzgHEURGKiPfj0C14YPLz3y2Dbhw1ZDaAbZjSzplVjewU/xqSZK
VMCeo2HjLCGKLrxIsv8TdsiaY3BBn5bHV3WOAWhkp58/zGT9u0UNtQ8nBcevk3oy
zZzJwcsElIgm7d5cPqaK/x8JUP+P87xbBgTM48csvU1uDfEsaNOv6hFd80JBQ0SF
jFF/skg3R8uk89lk/FrnhFoewCcUea8bTDbA+HuIGiVSIbA3e1fezl5k5+TttmjI
eunTHKCmz1ZrgedEB9qEqRaFN5evssHmtmiJIsXHsN26y4OURapr8OEwQ9ZFUqpq
hjhAZI3POAS3dalpR28nyse1ivXGOJT/fzX0NsMCNlbO4Nmme6W4ppPY/nwsROKa
sazYzackabMdMvnkoa7LQt440L6QyWxtlPQhucdgpSzVO3HfNTmN6RONF0q5dLWh
NbNqcGp3ZUyTaBwsXVnlNYshbT3yYq+Lz3KhP4xf+8fjgTCdEJOR31dYuMthk5Cv
uOXjMbCn4g0Hc8g6dXHU5qRmdEDC5D5Bu+7mWQIoyoSVe/PNh1ygTJg4Wu1PyXHs
nRqihhBV4kErHpzLbziVUIcpMf8My/K6EktXS6S0KwNCZTEMEkHgAKTgO+3h8yfK
lLB3btPDuSwHYBTfyQtqsp2tV3FdcKrOwqRVjxJGbvXC7BBO+b5BEm4MdoAicBed
joTojhdf7dxLZB+ZEL+OhKRVTK2th6Pr7C2WW/qBHXNtjiu1om0olQmV0/qmtPoA
WioAI90wsvLOjXNhShPY+5BUBpnC5JaM8s+MWtt14HFYBUnn+PbXp7j4cD4gjFGu
4AK9fNcUhaEoMmStVN6JiXeGjRgUQCxwXTdQoWmFOUx6FLLQ6XI14w8vLpLJsLIR
kLxKMxO9VkO3gt/wGVMC+JkstSpLQ+zi2paSU3dx+4AJHqxw5KPqTZ1daiV9fc7d
Z1bMXSKktJq9V1R8YMlsFCnG4hjtckXK6kqg3aMnho0Eva18yCYE3Z/dsfcdjsI+
RoakFQcWGHGKRm71ndfVW9YVRRdMCuWWdg4kZFtVZIT8QB3ZuwgUWY8xk8MtFAq4
2RYFSGWFWLT8bw+K1yvQ2IhAHa9Tw2ak7/dOtxUzL9pEMFKbwcS8013vhwFR2xkU
M2fNJvatDSQCFFKlb+0zTuCLoqo3Rb0xm0CUaCWVFnsQeDkjaGfBgGzz/qDVygCl
RqeK70hY02pT87eEhqAB2H7YA3sx3YtElXy/j157+2COYNOAX6iEcFG0wZOKvcpe
iY7qPr4oIf1ZO9F9RWvY6BbEq2Zx6Rlf+qVHsbOxRimaqO0VtBar27zRltHvHXUV
Rfu0n4BrmxSjK4XFAtoMMApxi5dABplkN/4KaX3MYxdmgZYqqefxPCRdGnpzh5Fx
ah7CBZUHYx01NLn8Ej6Zb/Wze0ZMBBBzhwdiH6rjbin8HSeZbj6AK0qOuM2+BPRa
TTyY/aPOkwRSJaqNu8TCo5vV5QsZlBE7X6ySlW3v4K+gMkMJIFnKaOYVjD8FUHrJ
BvaEm0hOgBFlsbKvGFImzw/2cn8oPWAxA3Ghn9JwGSND6ylvPVic9ffai3U3pnBp
KTYy+Nwq52zcK/gSosL5eFYSowWgDgTp8iurQFhsqtUlYBczcs3wLa5KWakLFUB6
devIoWLKjzxTI9VNELS96SeNNYLYON1JGO/qlP5hPVW0qiXQkGpqgCMONazJ1ib3
Pt5Ax8J9SskyGLy5VfhSMQZBT80jSSy64RZq8ZtqS9m7p9f1dho4GnBBSW6Mz9V0
oZMLQr+1wevunB3rapgydOJzqgUDW3H0YPGrbFB+u/aREsDwMw4t/JblEx7t/0Bk
wwd+Afw/xx/mTnVZ+q2ok5mCu58y75z3yO3X984dFGR97J1V32OrP3c7XH2zdvV3
BMwo7shkoAvmHk8gvOZYAs6NGzaPwwfq2/8CAvxbIww8RhXbebgtCnQR6J5SRzxR
ip0dDWccUj/sKFipOD6n0Eu5oNw9vn+PahcPHpYwwe9nmUmcEslYikOyDcA8/JV6
Q7YvCY4rIACp7stM0O8pbegKeDsThH/c9qyqGq/6dZhR9ElO/I8N+6FdcAqw/NYe
tnnNEPERf6EFjFnqqKDz3cDpJmhfobknUzP8qpPSQ2xXtpILGjaDDDq5jRPsAXOp
sDmfdwVwCQIW/3BGchybxvc/voyKflUpalX3rQYhttdB0HOxvZQOpYtsHLdUykQQ
YTTJw3mvpt4I/t95xqcRq9/96JnRJY9JrxhBdbG7RJUn7YH8lr3cWneuHa8EXZS0
HM8dbfEqN3/GU1sggOnf6rrr8zFQ86ARn76uxYLEQJtJXkOraHNptp74eUnmTRU8
PNx4WLoQespi0VLIZrTCwhkoEtvW7Rg6H3/dOgPdiCJtLwCYp7PDm80c1ertKUS6
TUNaVzULDZJy39+AkOKCpWpTaedbdwC0m6bpnpzq2EXLV/2/kwJvcB6VacLEo8rX
YBj5A3aflULq09VPVMqTHmmeH2SaNGFoT0MBLX3Ea8LQvYrpJPNiZiN8y85m1dYL
DoH51/qQfU0uxhOETlGtOO0OKGyNxtxzlBMLWWl4tPDypPu13NFzs54rcJLGOx3J
+xo60FBHHSWkPCCc791zNkvXX37Ehvbu1trBDODqoyqepHY6YeuoJFfAbx6AwZDC
rH2USMOjEcLeH1/NofZiaqc/W488VDNGDzsH3iwA1yAjIfq97DJPiLV8+s0UoYyN
JxNq9tDNIc5Xwl9ntMZNVhOItaHpYvwhq5MyvTeks9Eolak6+WLG/LEnUQ2zBTui
g+NLzkTI620KoLBQvVIGVMMg5UvJg0HNhIg7KyueoB2V4yr+mZVgfvJ1HPQ9QUrW
eyzMymaRdkBsskWRNyCtBxFZ1DSJvjQmSXhCPhvdLC0eBnI4v33kyidq1GwFr7sw
EmFlZzffB/yQ5rIzZKY83mDDDm+3Nif7hepxlxkCYHn/sFq0BcJnTyC0hRHtLCme
ls+vdRMYl0f/JXrnYjDP40p7CcljWb+4lg6YpxLEc5z+9D+qGqr+0IJFIWOfZeYi
ZxaNktB3Tx1mRKaCPBesjDRUadb9YgT9qz9FfJbkPizDLhUtJgyPtsf9vjOOJVWR
PE/AKWqA1Z9L3ad6sTZRXs8mls26jZzpsDgL7uDJI32+6ny481r28+dXO3rkjLQf
JNLPk0KwiC2gCGEW2JE+AAhsJ5CVA1stzOiGsKH8jnawFulThac/rvArAIG9xBcP
5CnRE7RThqeSYg3T7zCkj0AVM3JKmpOEyR3G8efEyQKdk5FFQ9VewW4V1AOPszIH
wM+K+esEtgabM/Uj/xEX01xHy/mbJz1eXC0TquLPAl9T0vZLgJdv/KlF6RpDuNUy
y9wUOHbgEZVYx9HkRwGD6uGhQuImuSkJftioAbYEQfewDG5u8uPLSUZwbkQFNkbN
jtNtRkPoJGW6AK6y5iizSyQchPEFzZz9EioiuYv3Ng7L1hGqTFWbsSe6cnUH/hci
PAkSuTlc4CSjSSlRDEKi3ZqqNgW9fjGCOJnx+7x+efXfkLy6TRIRPTEU+laR3nW8
AJiZA1/eQ3QHMcLXYq8eLAWy7rInGFpKR5HvI+T5F1kUXF07yhN5uvxHLGr2SLZ4
6AhDxKVjIs0uqFZGr7VdlLxEusInZQQgaRVidlYBNiShUL/+HEkxjK5g6ZMGHL2I
Jh3ioRqox45eChUH6Vm4ONOM4MHPER0USBsRUp5dzEGvHT0pWYZaU1gRazafYlNX
FoiXJlNvlqKbBqZK4WTT1bw8zMsVATy6U/XRhwDkd6UU/2JACs6/aV3GtpspuTt+
HOW3grVAWEkfLhWkG15VTf0Df76mJ3A0ho/xLLrQVjrCWRFcILLo7/PfgwAwktoo
BT0esgivGBT8p+nwgDqR+MZgdOFDVe7iK8N44Oh6kIZFRqmlDkjVABQSZNbXNuCv
lajlVyt0Sv/VGxi0Kt0nFUtS7rNOKVDvKHKS60gVFw27z0Yylt0qeNL2Y2pJ3ILY
2F7GQD/U91kjs5OgFjgONKQ7t/CaTpFXo2VoL8K6JT4h7vGSscjtea//4oxgdKg2
nQu7Klr8MLg9ewk3BHIaRpnKhpwvdzkwOfYkEPG+a7IsCHBS1Urwt2ZWqLcIkw7N
illMZP4kYScExs/wxp06L98riWc1g7iIHX3XEpMP6QhY0w/R9wwXUgC6SWFXFK6F
TszGFdMq5w5z29sV+jgrx2k/OAbywmVu1IsdR9d9pnc49+vFbNG31jFq4m08vA3/
uC4FtRc9HZpOPCSSsJZqaQUy3yg2HP9y17EQrPmUs773Z8+Ok7HZ6ImpSgwKaisV
bPB/y7pc+RO+XSdREwPU0PML2WY4jX5UwcyZKxomvfzNHlHEuF5l7R/fBkuHPlU4
DYMxI3DqsIIoggL5eV7Hohz9rhOwZhh8dKxS33nA4sHL7/+kLphaK2SjAHJeCkzb
Cz2WVbrEuvDjYAyxJXrqp3o/6RsoVS2WXM5Jmu93jai+tDSw2lJKUzAyBYmAaj6G
EoOp6KtPPQPTmBgHmKx2LPDaCitNYhFgSqCh4foCOh5e7vjLhSZANxiGEgnz/4Bf
2XNfp5E6OEnSSd5Rc4vuLWOPuo036yKDOO1nZ1d3EsSE/LSv7ReG4B9j13Egoo+K
z5LjjEVIiITagKwvf+ipn7wIAquECrlmfATdf+9Np951YIw6v+lQ9od+WhYHD3hB
ZVnJFWT8mmpZFzvrxzU1GwRUx5zco8xCR1ILTn53iaNhIsDRlULd9wJPXTJbK9uH
CMRcgbCan0aWDtkRb6oaFxSglh2uv84x+FsXzSWhaWIh8a720VMmP0cePKgI4TA0
YSiUZzresogpbZxH+tl0nxIVAHmeL0GBviMY9fVdIIzJaVcqGCYwcZjVx/YVPn+R
XmdYHU48YiH2msVnoW2xyTQl0RifD4CVu7upAMTZRS/ImhKA0fOdY74eEMqP3a6g
n+dZDSIAJJ8G0WtqCRzo5qs9qYpLjM3CFlFwJrIFNzOoG/YfOG1bD62WdDx0WpDz
aViuL6EINCUGpvTxTaoChwfRLORr7O4tGLTBzfBqTe+BwmnrHhDnrdrKBMMlRyAo
j/YkEK0CirbU8W5YcYXqN2tEZQ4+fmM40GBTAfuHgfAZFPfpVj17FikvPiCoR+yo
Wm0xNamkF+wBbm6/RTglvPH9Tx5jPaRbxOIwL+kcTZY3z8H1HF17PSYRQpRuDD2W
X3pI3C/deX6fJqHhQ08IxNBNsyJ5PQEG7875G5qZKr8cnUVo+wn3M6FZrOoqUnT8
Ks6FmW09b0WbrOpcM+l0PZRzuhF7TkMHI7cCcpw6EVb5GgjCtvS9SSZpW1ijAeUJ
B5gKIKnjmdycXclxx0UuGgiHZYag26hYIXwqxthnBeC9fySK6C6L1t9aoJNZQduO
gYJk5kahzjpOnX227OTgHoR0VLQAHRwqJchpKC8qXZOCgLiepE7BvMsj24jzunq9
iyMaXfR3sXMNdkHhmbN0gvhbs12caVs1BjyBCA02JUPbF3zvrsmTvQF7FhhiSpat
fzTWnPWuGySSF0gZ1ixcjaQwHgYI//nwlwfmSe/gisAbwACxWpEshl9RvjtDGFjO
2swL/hl7dd7MoPqo0ciuvqRJnTAWQLOSrFZ+XCPXqy2lPQb+VlurDlfQIV9nwVXx
IYHt+8Qs+OkDtuMLgAUIj8Jtk1ngDaMN2IHzqbttTczJZ5Ql/lss4UvZiX6/rdJI
rZfWBvT+hrqKeh56I9+4a55xB//7dw9rUd3a6hYbPb0OuBKoZN6fBc0LlP+Rzua9
4uNUcvyzC1wOLeqVSa77prZDGylytLsFXHAc6qRizACc6EiDOMVUzQ/s4EJirqn2
vQMB6t2aOBQsavi4W4WJ9HnbI6faTju2y283+FvYT7AeyJudGBRgwEFBEnWuirL/
lIzfd2GgT3FWKn2Yb2+vaWcui2X+DCm8LeHwathLa+dQo4Pu5IFUViFgzeSa3qO2
Ym7eWwsHnwg0hTEd+UQaQD5v4VU4DzBKs+FuKifXW7Qj9D4IMr/3LdggumQGFW3k
4FY9cCn/TnvTdwt/zxXrahmGkDeu6LN13QL5mccqvbz+G+KkGPjW2Eoxhavjk8Kc
jQtAmLkx36zRu7KLNmFjC9MB727kmD2iN1pyVAusdSKZdyYlIoyZzP3XObOYxrtZ
H8zot/zzoKw2phB7Qo5QDpKAb5K+rUYy9DF4blpionSsU/7G0LsS6V2H1frOp/Rm
Iv0/69hYpAFu98xzVqf5xIkQLAz4kzDY2yXJSXVc1MFExkoqArowXfZtAhTN8opT
oC3+sMZ1Y7SULQHw3LiAC7SOC68medCKjf2K65PbJOirabD1/9i5fyR+tcJbW5om
XuALYk7DZg13iZ65ntZ3pEOrWn/kFCxPpvfnANcFW7fFenuFNpkDUE7UiDPx7Noi
q1VHRsN11WNRtQNKaYmzMnkHxwlyb75WNRWrx2UIn18HRnngF32HKinoaDdn5dwo
Q6VbjzXqqt/kqByK9yBVxd6e/uDAQ1y8jQb7/MMZ4il5LZ5GGioEeifUAKsSMA5r
qTz+L1F6JRxvXldDSK4ylHDJ65JCWnOwFj17pDGd2Ynbw504sW00TYT/6IeHO/dr
BVXocXKV6pfRVl7+J+f2QlIbfOA0tOwMgXno9y8YUeO8CgKWH60pPaV1o+gqwiRK
2Vgskpul/J7ZJTRDauXQrdHPZXqlvCGSaszOil2/j3HEG7M77KDoA1g8ffZUUBsp
+LdjhmGG/HtnEZSkWrnIDg1M8l8vbY494rQvDY8+7SE+4SYpmK2OS2MmbIQs0ki+
gJU+qSZiIGnnDa/sNrZN8+AnKJq+WEFZUSmdy6I4pwZ/YIB1r/xEg2KHgk94Vyli
jKq1yVZx/H8XRR+2r3Ln3QtQbtun8aZzh1C6D1HWt9HbFNQbOATXuon1KxwdAmOG
Rjn5hpY19KtdNXRJJ3eEzNWwhj4Hxuwcz+7+iQ2Bk76uP2hVe+3/oTNPhhIdJlkl
pc24wP5smthyoy71QUZi+IkYpK3iBVbV3OjHYzL9RuH+WGHvk0Gj75UrsI5pKN+/
XGL8UOo15k9jjzvKHdcvvTNjC9yusVxubZQfeSAPOEmNorkdxqVII2+zBEhaCohs
2iGdbQEtWq3zdBSZ3nc82yQw3gUT48+Xet/YUx7FxMlNY9FbSAf3qDwPd9GJBDjF
1ySOI0bNZEh6CpaVO1sK5nNGAI6U/h1xq+IzDdxs9D8c3dPhJ9ZY9OKtJnLmgAKv
44IO5QtLphK1ypAUBDgq41C5S5PHh6APEb6IqgrZW4gwodh9OUI+3kEpGdMXgTQc
/I3H/Az03s0xaVZZ05GZeVUC9QJ6Ae0snwFMbUrJ8zK4WR6/7d0TISvL6MivTMfK
pCfBCQ1iO7EJMFnfnjYF13Y3MmNjIzD+GwGY3CiSknMkJiIHl6umfo1hGgjginIw
J4BTT7QxypYgH5Thvasy1sADXYBBHz3GCXglSvsmUC4+BeIWkb+N1p1XbX9YvyYb
jvIUlJSCqRauwPjAQgTQfc/+mtIphvqmS0qlJsE863Q65ICmMjDM6DyzIfjl/0sV
JkxbJw8jNwZWOPydmpv9rvTF+RqSTZ6eBE4o0DnQseElJ86mtAXpQLeN1Ng4nUWa
5PCUz/pGJhvid2Fia7cioW3mzrT2FAExbDur+eEZcB2INuxz8FX8JxoFUMAYTJ9i
BKu3Zb41tFtFj+hhmk8Ldd6FGSLl5PQ1ZospNPIxb67y80a8/K/7/yqHJJI58dap
D0aQrRIuTCX7QwTx6nYY4Wqm1UCA9YFMZl5aTiVRNlXL7Vu0j33myr+FNeyAqkeP
cr2GTKIeAHdDhKoQBmPSyP5IZm+qQa7aPVHmBFY1xD6o+0meNhRgiCBMRKR54p/D
XB1P9vhsEkesaB2PNLPrGOMPI4CA0jwsNSgeU+sVfOg7o8ezeoOHI7YHI+/dsE2I
MiDBAKESkKp6dP5/iklCSlDHj+80krIWjJ0ZP6dSMCZ7170wnpI7gypMGeZmUEqy
9bnKSYbLbJdfWJ/U67Z4+5Ai6fOobByZYTvga8WH657ySWQyVZnkMJKivtNNF8Sq
SjQ/cf563XdpkPU/wmsT9z1FjZ6dqywWI3Ff9OMfR0S/tuCsOfjEyqkcrapm5Bx3
KIuo6HTbKGPH+1eYwLNLx9uUEII6zLCegFts7uKN3ZFtksOGhhg+azbVU7CKU+Is
plWDMgD4VuQw4nUdlQSQdlUsHdRYI1Mdm6eiigXJazDgkoRiYUt9jtqPbo5vp9eo
5GgajyqJ+r3T23jiYnmoi3d7CpL+fgu8sClybYXQyK4P6Yz22zWlMbBHTgf/ujj0
uBkRwWaLDBKjbza+XVpbHDUCzfJ9f0/fCMuWwplwRIO353Gpg/rLkt8I21/iy1bs
U8uNSb5A24qzFB3pPxUEvmHPCybnhPdAbAkcX1SDg6tI6BKZS4DdiHEyn4oNEU96
dNpuLb5PyiE6PlAf6Igm8QixMUKcOdM7If21XnOR5xSTHhC30UmfNUwEIhoUasmo
MuRz0LF6sPk2NKhEJXna9dnXK+PCLb8Pqvk40U3uWejue2nehvLwkWSqi4ZOSD9t
BjWjtOyZInGVLaUNI17kdNBS5QWssspGkTxejIUjo9STLdHT5KFbaZLQhsU3M57/
CHeIX/J6dBcAiC0vNtsKsgCLBDoAPFBiFX+PU4sVkFJNCbJjGicoIYOqUrmigM40
/qo2ye162yF7OKPloFmvPOy3vZmkPPcfqVg1JgxiPGPup5n34N68WK6uSd1DAha0
kR+45KzekuqyW05eEwnJFJNDW/GlhXNFruTt0a5i9Y8aZMdpjLZ/Z5iMroDHgBxj
xJGe+yB227cxfZeCzcxt2Ei0thU2QLI5u/Lzep6lxosguVo0Z3X6WKCtFO/uIbkD
tolYcmWxp39A/n2jVIXczBWnw/Io1aCUEsOUOUmqhVZ5MkgltZjav071KB2gMr/m
ZXF644pAkV9j8utuPgKZfRhz7EuPZ6L79dWfSJjDoRW92JamEp7g57+/+0fReerL
9oBazu3rbSwYETYhv5QPJItDgV6OW9ac30+Qy/mKc0To0eHydWO7oHk8Ag1eyJp6
NH6Mf8yKNY3GPc0/BcFJMC5a90tJjWhVtRGhEiIe1s8AHJpT/0Nmnc4VQgjI6SQK
p4JthoJ1KY9Zv4FZM3ih/dblopmEHmJ6L6CpT8xHVB1YrULDX1K0NIGPKqaGDG7V
tBJPpyCJit5qBSY78jWzfUAOLrtsYhGsQmaIa0EeQbtKHoONdRGK16Uk8elobzmT
PbMp4P02e4kxZT9PRupsP6kkGL9oJPN47w6J064WIuWsYVw7wTBcNdFFeoodZzoW
+si9pxQ8TCwOqysM/orlhDsM3qsnZ2uC5g3a6jv0REejyAQGEddB0xeZGxX0SVOp
FgZyrdwDV1z54/njozrJY/hmfsVDZxOA2WZYMNoP/soFsF6tX8Y5IQSBHtYD01Na
h5KPKKsEIes42JXJxu0zyr9Mp0Lf0Y876a8a40sSxWC3+dOGY+0AAhSGj+HtMbu0
p7p0wNN77VjNyklNCI6uZQAgmUgJeghllbPW1+LGvysfpEqBwdxYdoVi0SSzNCLR
AAd3gJZzWDho9T4lw6lu+wtjHafKaja6wfj3MUztpNye9iZq/L7zrwxmznAVKPn4
q2u4+3csOrwKxkEn8yok2WhsQ3cFOEde9pyZ2vWH9OlZGqexiz26rojLoKUpDbmz
4Je9gD6CuKYG5dQjJ/meG0pZdpptNtVo7Z06bJ+XeY26tch+0E7WzhpIbOTrftsm
+8MEGlYMSFPjUn9NZySj4TbkzLrOI42r1Ny8Mos3umUiouqC0n5TqHZm2igRe5vM
qv3JKZnq6n4mkM/jwKEqWEGKcqDtUgPUEX5up/r4RTkXMnDPpW9oYG34SWKH7qL7
DlfSukFZFf2+U2UBWk+bkCDnrBjX5/dHE6OgnuxhPzzAWe6FSMRbzsoW9beBwt4b
FTnUCEaGuOa4o42GdMo/zy6Zs94LynNpAtBzmMRwa+9HHmMD9NP4GtkZHxnUX6zf
CImQxsIwsBWidJTAbZqAqTdvP5ht+UhQbHfhCOIAyJiEZUqwDwwV7AXA3/K/9ilx
2rk5GALfkOv4hFSJZ1BBTDr+Q7BeEaBiUC7G9pSR+gI9iLj9TQIdAO4m6j7agVV4
XhcHLod50oPxPkYWJYEwGLTgvpRyvpaK0SP83WGQL/Skm0O0jmKNpEOtmTHUwlPZ
lVre9PdAIaFkbM4qWDhU3o/zY4tWtg9igmQy8rV+IIWPQQy0CyDybg/emOwhopNW
WvvczMLlYP8x8rG0w5ULobJOVLMAYUvCd8Jq2qC7mt+i+uDJrUMkYuxyw1O0Bp9n
oSOKWkZDAyXeyOqYoEcIJVd12LQNG6HoTseojwjwyoW/kKKHKw0GoLK3h+EvLzVc
ojZB+BV3kK8Etbx0arAQI7w0B94JwGxbEVuHxOPDGsczSyCyfP5UMnGDdRK46jmc
hLyveV9KZBAlyFT6cl+P0+V7B/XcMd2D6llAGSJVlYLS2Hb2Ltad2VZQ0QnuDN0P
H7zZm77j9c7aQhygzG/JrTK/+rkFtcezdgcKFRH6U6J4kuXQyoGnP33sOHwj/MHC
vSfYC58MlUaPJ5maS9uiVGWmUXL73n3fUfNnI2ZcwojCwcUHNaBbM/QMDxIYVBVg
16MDPnhGaZKtMBrxprC6o7IA+GqgHg/lfJ67rykihH4I8sPa3rLOka5ABIibeyhj
cRDUDC5SmGSBcPqR3ZXiBp4Wi3iwIZ/RG/oS6vSDQq1p1Oyo2huAdU4+bdS7/O4d
cSQYGBU0HUF4gaYClCdoL+yFLzCCArFJLO5ASKtgbEHxNx3+40dBOcvSE8mOuRnf
y0u2e4kQEZ9IMJdusuQ8L2EWOg7HNUBv7uNMhXFGPDe18lCHj8AroPMH4+0zK/dM
0JMZNhRn+yrjwbhQuXwjXkGEnWIatFTZR8ZfFf/uIQquuLbTf8oSUCMtWeCgQRZf
Pl+fRiYeKF4652vEv2pj0cy1XWxamAowLuzokgkIH/sRSDPb5EAW1W87TEVUG4X5
0oectgcP002JrFQvowhBsvtN1BRU34tI0oP4tutPP5eH+Xg0RrAwKTgm6tKaQ+W9
C/7OhkkMzxKeWHdJCk7mfvcCVbgl7zC6kigXCVw8LV1e/TWorOHi4leign2lAEvL
xsZ3mwR0cOCE7/aJ8p96Y9letrytEnrrRhLT4u2DBYpEyWO07I/caaL2Z18U6+bT
fetYg10tj4WIqJO7a4IoY6bdYj+gfTfdBeCRIHBm7eEpQDn6P9FRiEMiQzr0Jz6U
KpkJkpElEET8A4us5R60qZ3dZbV8yfrSYcLga34pAeg0TSZayZPqMlNrl3FC7tuX
RDRt0f4YLB6K6ZQKJdIxEoi/Q5DztkcV2q+EAyc3mjs+o0fp6Q7Ii3+Vwtxk2Bo0
WWXvZkZBusPtHjLWLmUleRYPr7HaYV4Mn/E7jLHbht2OBwtMFxN4uOdFAbPIyUQg
zZjNRBnDYICp3AKHM6CGqcznqYwEBAMu8MBvvabH4t1MrfwHhKf3pPbtk/ZNvfdw
0xM/EQJecocHmH5rft+1y4fh8q8NdtN2McaUNl71FmY2iiFet+5F5jvBCVVyRUqy
I0Fg6o14sLviP0LyT3qEeDof8adHFnZ0F1zVwMMCBJ/tdf0QYUKaxsFR3J8L5QhK
1QryUJQf6RiiWXUkWqXACUbvBPOViu4FsvU7Bx/6ItWHbORHQ88EhyX4JSK/7ovl
q1St8q5SZZoNS57v2jr+bwxuL4Li8Rfqq6Rt8MqLSQFmzIZ8skL9GcuLQs8Q82JC
aU3OEppA7035uEkBitLS5e38pPMNF0GthrP2Au8ZVI2kyGqohNXfdvVxNL+mHpY9
uIu212NMld2wxMRlDoHr12eUP465QuTWnFL80NX5T/SZ7s+L6unzjvXJOCeubHZ/
48UBt+89jHvgO/GgWWPEQ63kT0ImT9XSpg4/lN3wQFrwwS6B+BzzBOEnwibBd2QY
wwZExRDQUZTkiUonnJu9OL/d9uvjcT7bvZsHIjUVNOPHhvWrXINgixYnwDBX9V+H
BRd5jkPWDnlZLa/+VujYM3ZOgBid8e/muurqQkNtX4Nt6IkFivhXftyOtXw1VDvi
Tw8KBxKRy5u89n7vcJLuKY2dHGD7Wy0FcbdmpBy8/Pgmfw7AS+rxDI3iEHFKOiog
slegvwV5TXg96O+HyV18RbVoa4UP/YEuYHphU1ud9wvzWdzEWXH3TOipRylxkJ+2
v4ZOZ2XVKneoDDElPIsGRHxbFys2eYCXcvhmul/vh9Su2opUQ7bTbRr3CynU08PO
a9CbrJqe7ev9pNtlED/LNictMBPXVA0BRikkckh7TMXvyX4AGut1Ba/ElMAMf14a
fEsr3MIyIOu+a5IU2/oagWKXIoNlW0We/oKmAcKiVwyKiNWhGxmBA4ufFHEL8kFv
Xur4rd7KpHQJOkKtViERtH5JUi4b8UwJ0kkQrCcDIMd8HF47Lap/+CPtl7wnL+4z
tjT2/pkBbJ7DgqSK6C2Hjx6LNmhET1ZIMc/ZU8TNF4BGnjR5M5w0+SSWjUrSL1tu
DXwvBEeYAvHkgfIQemNztVaLZy4PN+hazs4kYtoyhCg4mkjqiLpQgE80MhaXNRy3
eapVqsOLJKyMy6Kdrfz5tY7tOVDm28R7fzfFTzW/Wf01JJvl/xnzBaDc6ETOP4mM
3vumUNQe/qghICDiP08wSi0i1n4vxRuLLVriBgjN/phaeHp8bjEm/YAAWAMNl+D2
XuxnBRnx0bb4SrliHWWFcbMDeohuX32r8512sEsBxpoKAO8cYi4Ru/dR4kQXBEtx
iJ+cA8vk9qL/HkSeaoWIM9U5PMLdbJmK3g/fy8m9c1ALbYrnIUjwLt8EDk8WJYzZ
7k7QaldyV78lmWARBT3j/V1xpkdOjzTExVefWUfpwKXOPGJ5RSfNDb9maWw2KAes
S2pHfD4jXivFWYucVUrjrhGdh8kdd11nTmISYhL5skp3xhjPtM4MfYYZPBFVpHIJ
7GIuM8HSBw+WiTwc5i49D2eYWQhgPl/BHlsR0jyweVf/gui+2cDje4ZTjMX48FyM
5BSL7kEqG6SOeJqzEplIh9zb1gMq0OO2TgXLULVEIsrzTmqOqu5+qcWf880Ht4t2
rwsX9pBqmsVzSYBOqDMw4TV51EPfau57o2mg4za89f6aGDOhxSXsf21v+4akI06k
w3eBwPJ2CjDQSFolu3IhBJ1sNu14/0vsM28lmBSUqb5Vp/I2KJSOY0dHNzINb8dL
oh/k+czpEz6womeYEUfpElbBGldYOxBEBcrGSW+K0aPIxP0I2a03p73JqqtnlyB9
KTwbyuK0ef8ZydJvwQymPA5+91lWI4wRNyAFXZ9K/z8z3KR+/A2r6NnQje9eLHvY
vt7lB4ZFFjYs9XdmB3UmAKud/Gy79o2bJ4AuzY2wsdGxNatOxvNOYWxYLr+kQZ9D
8iVsp4P8Ws2eR9sZhiFTbfG+8t4vkL+gmDJRCsz5la9K29wmt3dIbuAngVUEAf+u
6mtj52pvabl8MV6PAb1EXuAcIJsJhdfDu7l3IpvfpDedNaKOTC2JsdgqWEcJfv0T
C8QIAvQV3Q/Ffhi9LSKPW7sMgDG/1k/slYUOmrSebBPXebSeF04QSb3e3U5WoIC9
ewVqce1Z9ZrIa6jLVg9QIPzqUsjr4Mv1gmHYjMlumGREO6ejzVanqscrEf4/duHH
znl8uNXvOlBNf2IBb0mdzPispzSm4lWsC2jNfWucJH2SboZTXxDiN80pgRM/nzC0
YKxCpQFg4prN52ghcaUYlkIQvbwCh5BAs8tndQUwDm9FOOImyVyN9JH8OXASeVFD
5UNmm7ifbCyJkI9kN35dL17imdjTv2MplFCg0/5BRFWS6taDPOxCb0YC7OibT9cz
2+52izfEkWKQQqnEY69l6n3zr5BDYBmcKx8I0YDcUJmgX7MFsqVv5LYHewsQwfA7
f09Th2OKFr9fZZO+/NgOhQlitHLvb+RoyzKVg691QzboVvcbr4VvckOUXhdlDXSf
px+NxsDeZyFH0fqZQL5EaYwpx1mSKrU9pwdSwZogchx5I15t8DisxYRAVAtxw8pW
qwrG1C5XGA2DJaGOPtcsFzZ9kk4r1HknogSQ0iSozDJZU2WJeYlB3CT1c43NMGhk
Mo/piLVq0Y+9YnAi8rofvqCGKRolHJ0+UuBnKG7Tga3uWKMgKk/NkxWkUQXGmziT
vh0nZLdhwRDZAxKT1KNsYap0ZGF6K8g//CUcgfXKAVcZG1ZT4isa/aMn5wgVUeDg
15bYLaOOaaPGxl3ogXKVul0oq5J8NozOpJVqNa7K6ueqJhn7eX1Uw6GgpmR8M0Ff
cUTbQ875dcO61/kDgdbsfU5ZbikahhxWygoOk2mNuF0RNT76Xb/tyP/kcmR3kOty
rQ+4HiUx1sRSCGnPE0gzAWaOjw6A2rnQNLFPnJGtXxWNuXZC4axa97YYjLHTLz3V
TtTTqBXSEgDleKoTl4vBzGfz/Ix5q5ajBk9MAFc/V5hAFRhEdzL/zXzA3vzbyf6h
p7BoZEkR2hMF1wbVJKJiaSY1Ft/1XabLyAF9S/9D444Nd9V4E4eTHv25yz+WJSSL
N0b21IE3U8ZHhMVncRau8WQ0kMbIGw8c8t9MI6mpsmsgynHOJ6yCXUXoc9bz6Siu
cq4aas6b0pc+cOoW/F1mxdBU+wIHqtjVfj9PfH2cUN+E2BrFzxxJ7ydWVNJNwY+6
ShsQgFvwsBhcGpcuajRtoXNGypR8xQiLu2VZ7PA/QmsLB5lXh+WaUNOkDauETGWi
QdJ+ZveXnOTolY8PmjbnLmwzPHiRW5dCSU1gqF7RS5DtdDBSDp6VY9n8mBjWaCM/
8/pQcGZcLOhsvpK3qQHP9Aqh6c/+R49VH3u8iYrOBq29MiaGskpRWMmi2vp9hqKw
gwgIKMlyzO6vtC7N48csG/BK040lfHSAGKbrpjWUyyuvGDsf+bEEHX9wO/m/2fLo
w3/3w0amzT/ycl131bJ5NFxrP6KLjFAAK8X+vNT71qIRYf69kz1GoXvIP/tAOhAf
9CaFa6Izw9/577RNZXRfOzSbWOwcu50mh5HFZj229yGWwjA/EWzRcsELphDa02zB
VXqg4xRa4BCCn3O8fK8ClBBk9STafbyYXJ28ObiehQYyR4fh3DmXCJN2QJlGyuNs
N554pd038i0F42PCFOcYyvKSvdeSO8glV1r29oAdB4R1/czSUSnIdhydFPeYmsMm
DCqyPivOETUiDuo8m5cIwOJxLT96642Y749EpqjIOcwj1ZzVyKXbQqfA983AuC/y
tVkp39n9cZMer4aXo553OAUfD07lHCzXlGVGsECwysJFFKLldhbDoT1tGjLLpw/g
XuMZeCQ4e7KYfVfmkVtJY55wg/rWerOQFfBi1JZNz+VDsiK5+IndAgsdEqWVGIU+
17A+JHDJw6PbnX7LUln8l7C2sjJmSCtVWZuAEDLNlp3qIe/GMmjsx8BFfcNWZqVy
62E/d9HfF+K9+C/etaLsN7UcPghgSKQITcWhi4Ck9Z6+e/UTBy9QaBrTWHE2UVA2
oEp13vu/dTEb6UJX/hhyxu0d3hkWYywFdMODCaA5Z+pfdTjZJeoVkxpGur/n67rk
zEE4L3cqYI6T2ZhA2MsG/pYNrrxwbNn+/n+rsjpfjtoBwKswd/5VwY/PWiMTZtjx
eOU/t4ZnoW1mcn+RE7pXDEWyGOvZjMrJGBTPwQGDU0Opwe6cU7aI53HSlqb5kAUe
JXqkrbCDLtKWql1gTrM7gXNYKSZZHwwVRtjULc5z9wGo/Yq3ZCrsHienoEnAAwmP
nRBpiv2w0H01YDdilgli76gd2zlooXV/ltQVSx3dLCQW8VUUk2iNUeyGLCneKhLc
nQrHbrkdyrRFgbsyNWeTHiIB3Cf7ytlwTCF/Hew64RsSG51+2MYq9d4VmZP8jC74
ad3oq8jTqHBndWL3F0B4L1Qi9WvsLnL3R0J+y6NMG22y0oh6TYZUovK7rgYvjHe7
PsnkF7Jtpx/W73N3kqsIML0AkOM9pbxa15hozy5GU8ecAa0cQNKyXBKxWKiqQ4AF
1X+Wq3Mm3Qo2yM/WUtF9Pw27YqWJvkCioKJEFtSiH/YxSMUpyEaaIxVl0LtTwGa0
WBxU6mzvGw87FjNLiHIR/eTcDXwLmhbSrD7wbwURB2331m5ntjKFsce+0Nzc00MY
gskjMQrHzJPvr6DLxVCfqIor9m1HnLVZDCd82iDQsqNKYMholdTX1XgW6/MPKzQY
3mpuMFo0LG775AGOuesJv7Ao10XTSIG/XiORB46EishOYLhXi1hXnk3MdHOFeSYh
tO+abGZVF8GNUjZcL3uzH9vSr+jwffn+3vpUsuAU7h4mKOzSAkhdCaq68DpseyJP
VdEZbNUZcPVYC25YtqWiv84csrrSXhxQk+peeIIjn0/AJ/0FCIX1vdlQIJyLc4gg
tkXk96HZloENgzPolojowmqcbBiOfdGxbM18xvdNWJETCmIXe+edUXenYPxfoGRf
65S51lfEYRuz47ZVQ2nLr8Jqcpl2lkqppxxM0837vuDsgqi63rD5TjnmjuW66RRk
ZgxJ9devZJ6R156z9NM1mbk7TH/nAw9AlBmAU19T3PNTvGMYzrqrOcS+c1sC8mki
YPWTCkPbSkxY31X9kGyoHSgj5QhUT5/onYg5zUq49Vg4S+/x9NQXQ25vPgojaIpE
SMGLQf3qHwa3ctSrio+feAL5Zc6xeMZ1geVeFlpQvNeniBe+2c6UosZkqfAEp+8y
PWiB0pS6NqY1wlY3WiCFlpzanqlTxIPwQ0Roxj2qhq96Vita5CIDLpyj6OaQ9FCL
bJPqJWFaXlKovTBASVERr+SEauE0kVUPQ1TqcF9NKZJOAKaEG51j0YLibP0E5YZO
xtrnsanrMbFscPGjHTNWsfXjeRyDL6vrtii6SzSVb99PCfvOElccPL0PkQXGgRHl
nO9JQQYXQYozNIgtTUTxk3L723XjUbQwi4of5GWZpfW17PYnXxYVjICw85m4xyzz
P5vqQVQncnN7w69HXjASBVMI+ZyzzeKfG+jHZDv+C49mglDN9eSqi0r+/DJR9bK0
F35qfPRE8pjYRd2Sx5995EX+fSzNfcD4D0M3tqOxP8jdj8aafo1YDwbl+YHj2FH5
Ybf9xZJtujM/4mEtTpWlRFw+z8kq73nlG870kjrHSsRhck0UtstX3J1a5rtHfHUt
FSez7ADEto6Z1M0LHQ3P4ObcoM+8wNweiEvSkFz5KaJNBJNmhakrf0aQYSjhNP7C
63avWyWUU8OoXZ+xgo4ECqnXBav93OaoEpIKuehemV56EuwF6wdvDE06YtUCEGfb
vQIHSAESmGnB7v5S7RvDHoBWlm++ymEY1fzSnmj6zZ0ZWVjiY+i+oeTzWxxiLK6b
tvOxT97MOF2y+Ia3k5RFSV7tL9Vb7bTaQaJRE9oC9djZS1NzG2Y2BqTN1uPjnJDD
2F2kRpXaQvGM++OlUWc8LYAR44qA2uBMQ7SQQr/59pItz8UHYPhXW7Pzwbvytb3I
7hfwKRYoQbW7tQSz/MweGBDxD2E33ShGFDzhGo+zNoUxOgPbPq5FQVD42aviWOqU
uhzB6dOHamWLKeHSmyp9Vd17bZaeRQpI5NEyL/40cQwipaej3aFP3fhhgsP8boGq
WkBDzXQ9hIiD0Y3ebLItuNCoVAzev4QlHGJF0yW9UqjN8xnw4Vl3RxBhNR7VV7Js
gY86gpp7NCIFoGWXe81ZkWVMejqe03xP7596wNGVx/qvQv/zP2AXLsmlCGAFPUw3
GrHCPut8EksiWw75N4nOqKkd87euqp0S8tzyNjgesPMqbWqFNHr7aBdNf8FZ/oaQ
MlZTz81D3Lfhi8rUSyrfpqGfOvPRG46KjiX/9rs87TXpTd5xojgh+oi9bECxg+N1
wRYCGUNtpNdjMI4rrQg+tONAzwEfDg7yBvDb3U0rTnwlGctTKq5Dd7RbQxN8BZls
vsYcMGwiOD6BXTcLg6Jw3nyFCYXhTAqj9jShFbzksZAPvrc0H9NpuQAVXu6AVMZw
YLqchiLL739V+XF9jlFlj5kDbHGKmJRJwhGqgn0I4sURrCGGq4O3glAc42Nij6oO
Po5hvHrO2Ieqh531TjHdPVX5lPHCCOcU9kPjZYliE/OSHwScEOtU4b5IPvv+Ez2h
SMzVfG4QK/oqpH5cfYXAji9wNZXeoFJPcNH2FEDMa5y+wCLuKSz77++fIDyMJdXd
Gf5fU4c7bQnRO2w9kWMIwF50V9jOispOW73Zgmhl+6a41uGUSFedugbR8lDeM9mW
6mfgXAAVV6N9us+B34uaHymLn1KHaOlE7Gv0fN3P2aO18+59X7jxKwfHLMECwKR5
g1d3yqOGskpZF5kcKLorm3sGJMyZK/fG0gVRQTbSCTApn0j1OuekpBv9d4/LxlVX
JbdMcAtQ4Zsv3XdEwaITwdcK5hS+bey5nfHmvnrkTal8wiod+RlZleMjmJS87Lt3
u/fMTsDpBkf8EQQKm0+zudAiUtZ1nS3RVlcNXT52zA4p7zELsr0SazvWl1lfsJTz
dPZI7zzJr35QlbTZ6BIPPDkl7ad1J+g9nrRD2NjC+jyJ4pJeTF4r427c65dJXWAW
+kPZFhMyoCGMBZQPvDJvzZ5OVlW7mYuS2rD+HQH7N/GeohkLhx489wZ1t38bPdB1
XXLNfS8KyLwLaICpR91G2ioZ6C4jKRd2BoMQP+h2pxlun6lMhDxHChPqyj/iw79n
5EsIeDZ7SiU09eUr5kubsOOxVsC5rVbDRkSei1wEwEdRYAIIlL6xRENo+yYlrRFM
o7Q0U+hAbyTJHx8smsnj9gA/7xV+7rotQ6n3mpzMxTcGwizbffrj1UUHmegiIAdQ
BgjHQ+oazrey0bRgoGgCnAF+3dc0aKpXcnQb0FyBr1Rdn1a1kpWzbvEyyOi1ATiX
MYgv7QDbGrAhTgFt5wpewmJ3aLqZzFaEaQUnsP2aZx5tq5QesJUDFMkD0YsPHlSe
j0SQZgZRVyzh5xo371IqrB4V88X2RMsbjL7uOIuMXCO2uyvgJ88B3ZivbbIe7SmA
Q+vXorfb3U4ASscpzT/0KDmsV9+ewv56mfpqyHBNjQbENcs4VOXR/jXuGbykp1fi
iGwyU8a/OtXyVigtfC/F6TZtmMZYfwkXo1GYzrRrQ923EGybjmwV1E5ZlyfWmY47
GzA48za+x+T+Sn6ozMs0cnDQwMSNrlQdtly67YsNIra84Pc1tECIUN/KHXmSNeCE
mT5zKUrSlLjiqkzt1FgihobfoiFr91Gn3m8x7gRDDf1krqUrzKRI+XpI+/IIu1jM
FduXdNCPuX+VmTMpcaywVOy/Uyrw1tmtO8ZTTwzban75pfwnc+XPiydXo40vyK/K
Xxk0VMeJoozp82M3qDJvA+Q9e89YwytU7YzA0EhSnzww+V7bHaWB7AgvGW6NmQ0d
HLmbHS0M8YEbncuaVXG82qnMF9FY0EpYq5eDy0lnKG4UATW+r90XpU6WRnqAEjs/
nCO+qtVuiynnQfuKXF4f9zbnJd3hmsya04PSzHQqFWnYHNh5tHp4D2ZvXlxWmOHc
MCHBjar4JrunnxrdEkl9s3kkL+XILAcCdLwQBl4mS24PbT0Zrv7O9KYkvvY7KEai
fVfw4kB4hkPAsCQ/PlciF3dK/bpGZnN/8KhlDZdqzbytJv8p83Mmn6UaA6tX69Ti
+yJDcSkjMz0AG48ThDGGzHxwXYPJhXmuoSRaJ/YUgDDSbpI3UeBFu6Vxi4EyDGnM
ZCS23miESYXu/a9Jf+sYoDZooKLJTSiDDWR7UW33N93Lj5JJDWHgE440sesHbb+H
yT9Ni8f4BY1BoWXFjNx5sRz3qhaadLmwSE1u0cQIRn5S3Mm82hzkuZAoxoN5iFWV
OUmOvU4EdO5hIoWPAoH0ay7oyoY1d6QQbKr2Gte8nvbg6LKPxaTHuRkhQsYOc61K
ypjY/UIQqv8XRo5zmgKB5iH/TsfXqo9ISKTiPvaO4cbJIIfsbH08JnGyMSMpQruK
51koyHdLc5oo2C88n88eAsz3QvT0uekJ9MajkqxGVrg8vldfRj0pc8jaXysA5Uw5
PRUY3FNhp7/2HqEZ2OI6KqMKA0wQ003ixefY5hAjz5RR9ARQDza/DYh21pjqVaXJ
jqCY9q0YA5AgsH1X9AB2ezB2CggOpYCUEjr66CVWMDRVj7DqRvb3yJjaB+NYd8CT
FQKDwr5OFB+SoArGiyCUr1bVmggpzY+VBsnzTeiIcd+QhKDKbJPg0Hdsc0PT2Hnf
BA4qEeT8k1rPXfSzNGZIRr3Nt9McCg4rAGRLukA1w2jj/+7ClOjqFk1YqhE/FVFW
dhiFwBO1wjQH7LG/TNZp72f1SDh0lhSUh36nlHb2fHNzfo+LolXDsEBv0BFJyaqk
R/hLEPYGXBxZ5NVQaj/irGJ6Y32Of6dXg3OzJkXNalPMZGUxjdB6IeqIcfoQiQE+
TVwm/6HTE3I7eCWkXuKZLq9g+uy+KGbD4sgTvm3THfDv76FrsGeqK212e5RQZOR3
rzFhxOlT9v7/WMAP1IrpfB8sCAXCSYg3yGnxuAeEXtBAn2b0eQKJt/TFzC93K7hp
Kq6z3HdLkeTLUstTNyBhCkADUMh8wm54vxXQW/cU3+yDzxJS6o2xBGh40o25uMvs
anH79BHtt7wtsWS9fLfj0cq36DpUN0ia7973WAZ1aFtK+6wHJdv/4iUaiTw63CfR
8jGyLNbb0v+7MSCB3Zfe01ZfPegjA0xZw8GuFA+nGLueLDClsO0bWiGKd5bPuehA
hZKcgbP0pWJDl3vM9tvAc6S/03MsxXf/x4ZCfdDlBFt8YBgFYn/YTZoVGqvdbaA2
CL8nSAQ2Hp4iTdo05Zc0wfFve/+ZV9Qn5Iiq34AEW3LQw20ui6BAmuRy+J3Kkpeh
tStbiZotdA9O6RttGwT+QFavqxyIDEopKydOZUcyuqOF2GzOj55SiOIq3IBMOnal
obKjnww5eoYSehNbF56cr99Qcfe4RUBxXvfS7q07RuKfOWc/euJjNgGd+dYhfT0B
scBn6U2xugODzSDkOnt8rfzN6GCe2ZP2UC6gaA9uEQniefvkSsLesSfMieWDWr20
xA3CzW92LuWYaMu6qSnKfH8MkKC8Vj5ur6zvLT93vkVGhvnVfgZY9kgpb/IgLr1e
RVIx3lwi5Sbe4ELULmWGX7Sw+iBgXcA0A/gVMsND7XhaSOVJATUtXdhK6ukvaNSA
Blu9GR0o9gUheaUoLHtyaIdXowp4YC94SLpq/CUixus9nrQsBSF5EsoOb+Gaf5/g
dnqVbLU4Dm3KzoxOZdO0iGzGo0hR/dqOrMWgOczJaujGYey242Na2t0lrGPHJ45Q
hv4JqiR5Z9ypJDswWAG2De7jxyqY0EzcuLNEGcK1gIIml6TGowpPsEDIL8UJpmxX
P+tl2JOnyq6cEVj4WM2ksS2pNeByjB1Dt/EZePEza/gAJ7M15FS6L2mUX5UQB+SD
LkfBWalnRwQ96HC9oi7M8AabDY+qzePlf8cwyts897s2Bbp0+zrg2DbRiLbPGs2s
d/FsgecpVmVyDsru0pIbbIXHWoR/yDg4dBSGiqQirv4nnHuIOYh1vL5UcjEcC8Qh
5IBUyaFrNnISaIBYCsw0qE5hcXQ3HN1Qoc3QVamsqObGuvp8kd+6LvFWSNRJ3wEf
NWRyZws1CtMV4zOUWngDm+H0M2ap6evadUY5kBUgiUAvFGERZbcZsRFR9DpCPCw7
cr3qC/N5bn2/j9ckBVMf7DM8E/nqjmPXiSsbD+Zbm/zNGeUjPBbXYDK+fRk4dfV9
McYdj/sbZyKKbJbNCXQQp1Uybdfptmql6YWobvmDl+6PZ4eiZDtGsA/3pm3wI2rQ
xVqdAPWru4Vqsiuzb+LOwIIrzjI9ooiGu1Wwjd9S0S0G1wIr4RgR4k/T+iVCJ9rY
vnanFzZ/hrhH5qJfqZPuqaWBEfSuCnav0EY/v6U37AOZk5TJqQrBHV6M+X7s4cc5
BbmZGAm7PbuyA62R8P6f0u/4epg4tKRqY6+/ge4X9z9qh5XwFaSSA48Ol45BcNKM
vrIS5dqURni+grvqU0uIPnurajJz7+/puM8glwdo3E0JHFanZhDQCRUrjbUId34F
dIbVnv172Z92nkQFFdHnYy5ng455UTJiPjtp9TZFJv13FWd94fDoG/v1DsTVyCUG
aFVqm4F/JHHgBvyOZ7PbiguFQkNPuIZx/KrTKP/DTe0+aUW/lgZmUOaDI2VU0Vv0
1YeQCsooPPFJW/9IvugD9VXPnMIBP7lqeeGDd/nAYnboiofGqBy4BSJ7c/eWJT5C
KzBmK4zrfYqr9gdqHalY/ZawMF8WoO/jprjZtaFKR2BizEPtj9bOXcoIVA8fMZnf
vV/p5J1u+i0fKJBKU9wjCoUKxIAtRdsOS7Pro2NYiZBZs8Ki36tFaj5AJyo2aaWw
VemBgI6FWU4WXwfX8BOZIuZvZkTm8moJ9wQCGnQ27SKTHCVjNIIDMYMXfXOdwmiE
vwiJaPjLgTn9GdPP4YbePshz+wBrnSGren/R+KDc7UEHL2oe5L0AC0ioY6spvecy
ovm9rGrkgJAyrBgYWUMif7+QOX8c345GIERswyGNaLPkoUSa6ks+KAnG/LqYR5uj
kelJdErqXXp0GY5OMvtUSz79NCsSZh7/WQdTo4cBUH3clsltprlsIKh0FLeszEvr
7d+YSaH6FGm4RBVMypXShZwsoaa0I+GTBPlEqDXHcq83lLSOuWHtArXEzHsZ9vZu
U7yRjyU0Ksl/vYCdSqyBeyADqasDATxghZ+UYV6XqFSTL2SBac6Bq6JDuFFXzGbg
gEmYH9jqbuIfdeJNQR5c6MDCY3ckLXl2R3Z7nqSn+KpcwfIKnRq+lI2qsmMTiy1f
bI0x/wNgsQTnX7ZtJhGA+ZKElILIhKrPDvy4DjTViWQcv96aB1KyduH7hUG7UpvI
3dKKHaR4KLiiFj/cC7Kt4Ri3ol7EvoUMw1SfxqD20+23DALIbPzc5AIYQTUJE5CG
1o7zBFsYfNVBDfJ26RdAB9DL16K0m52pGe+ytYZlTSP1k73wtgLKgUIpG/tn7kwr
BQzsEclEOyaFbZbYxMilnIS2bees9MMWteZQ+Cf/GPiaGCWf4Ppo4ZZMvlUcrvOm
zjRaUiJZzwE+/mw9QXcPcbHgeVadyMt6Y22L8qRMXCcDvrl45t2mIb/Um87S+0c6
YzGMh8ddFrRhNqlu1bBvT8Jqwoj0qW68d62ktw0LVH3xH8bMbpmacUjd6QeUSrUy
speiUlNcrDTby9rw3eZWaM3gS6M9P3T2xosXmxmlhl5c4jN4t6hgc7Tyu/aI1I4L
QxuD4eKvVQQ/58z3tqVUo4dzuNstyqWDyKQ6qphBJfTwuATtygSLdAYUOWDZ3qHN
Pt4n8PNj6WWNDjURZxYVs849IVOLKD3boX+N8abwXVrgrv5JYH1ANIOdEwXdzeX9
tTaqR1E7edTtYFGvKdN83dlOAAGxZUglv7oeKX+I2ogW6wHDH1OQclxQpg+AnS4c
1ZTqiTlCD/v/LRb3mFo0krtRQyblAFITBh0V2HFxeWSoYjCbUy8EbpqC/h8ll49t
48Ip7OH6EI1dxF6Bu0IKPzz0DvdJJlfwqucrBItWVMK8EHLWB74ggNBT1nKpYdqr
+7Io4/A9QdbV6U0RZY3STA4g6600RpS2ZYzdDt9upISOUV9hI9SL/Cdj6P1ez0Ar
4qZRZQ8a4I7d1cdY9FdDnO1mHsq0dzz2sUFJNivak55oNntwoOKKmKysFTqFZTZk
vHD4DXlIu2fam0c1OO0nWL69nGGvpRN1RNNfWRHkl6FhL0QMay9lpVsgwJVa1CA0
yjDY5V56keDzGGGuq9eCwgJaBu8n10kvA7rApYFJt1iTC2/9GAz086O6FmYoZO3o
tahL80KAwzqyiYaO6WjPtEVtqE30MzdYSQNRb3P+lbOH2jofQhFlWbbC1Bp5wKI3
3fvOJ+LLxwVrqtVUC8SQF4xq1Ds4/rw88PA4jrxLfg3KBPPANJFSA553Ecblb3UN
EO5KLpJkG/NigQNpXFB9SAnMQfaMjQymSHZy7DDk+UDPBBvsgSfRFAbWpk7gh5uD
NuLqJwr3Lwh1gfrvNUND9Gw6E1ESHlFHNgoWmci3oIOhW+WD5ndZ6l8PGsTUzP90
w46Qa2ZuOeJTcsfl5/UnJqDmc3UvMmj0XFWoKl2JIcLmAL2bd9JJq5iZgW7/AKdR
vtPk1WKBWKcvRRTJfVsZJih9MAO6AAN930uulOPHNhOE8yLE4M1Tq9mgbBfaMeVm
GeFmfb02lpJPrh16s8VGN4fCQFsjmRVBOo3iOTlEkZZ2gvkgAYQ4YAlr+aZVldP+
qzYLWS0iho7fDKtfolqygffOzthhiOlaxDv4j/bKbP5dEk5/z8h7OeMwvcJBe/Kd
ax2BTq5vMQxBpxI2sAglo1VBG2QhB/2vxT7A0Eo2XEuDFj4l9NAcCAWsE5MsPt1O
xKxdPlkCFP/G1VPNF7L9lRxsjqr8TodmsYZqRKYs09qe8F1kDov72O19Pv7yHnOc
N8OR5e3qSWRVAa+mkfDQ1iP+dymWMbx1xhR81wLDtffyrNUUYE4LP4FTQAcu04RP
x1u/2p9LrYw7pWQI+rOaqK4yu2YqK0gwbQD+T09a/ngU1d/9IJG6Haav8ZraxCV1
ituo+0NRN9+gA6xWKtObrySojhLG1Ob9p83R5a/z6L5dUGrlhKfh+QD8loP8cZyb
HzzQYqIdb9diGBV7/PObZZncrxoJoO8h627x+1VX3AUa51RQQOC2WnLmX5RZgVHL
dwPlzswGoxCM4z7dpKEs7vLS/Gj9tdOdgJDzr7AyNoK3wXfCd9rHljSplOuYYBTe
ns+r/cb17Fqg4+1XDwkKMmhu9tXiUY/hH4JHM+LFNyIMPdFSrAYLRMiJh2ZXYNZI
mCFPhKBbmmMNfD6p5P1uGmZMdrsJXszk4jgPX1bszRjD3il/l6Z46XUfoCc7gQQQ
XbOgnKuXkDgcWRY+lsOTL6XvvlwUrDxHSbK8hdcph8XlCms4Os/5X3S9SiFUDciL
fs6pw0G0TsiJG6kSl16Ye3QjvAeYqHfk9xdRVqCIF7v00DM2Gk4NUgl8kHJ7hGdF
h2F22KAMtBPUOPmKQqrPnt31rflsNsXum2C1hVa1lSTKSMjKGctep9h9UR3BUi3y
XA93/mJoHoeVG5yayBplnjKTH0bF47NfPYFZR2vHx3DrSyOoz34KNDbS7KwLPUdK
/OzemtS+Qxa8obnQOJgiOG4Ngsi2zHokevtohHyYE+ARM2gunrk0p6pD0LHFOrrQ
TLAPbMJN2Dru9HDHF6V4IeLru/saSjtqpfT42djuFDpPX+kqo3oC4v5LddvDnAKl
ymUhYvZFG1q6obJG/WTW6UpoYT7fGIX2FWXv16sbBPbhjdN58Ay65jqRSNxt5+YS
IlrMu/TUO2hukxEP0x9cYcXjHNwoOXWciiee0tKtQBK+16FsUtsaIbYXY+NQeQbl
ezwNGAXyzWy/R0ctICXk/xVetQEkhLwYqVFCyNxs8hiH9nKWe6TKScBi4ogW7w4s
QZrL12d4BfhFcqR6iCpAHrYJaL7bW6qg68D+AOSNF5DNLYbUdvpMvKU+3BxGznBy
YSbYnmqIiAuQS1P0aQITA+3qjNd4zy+96yZwp/Y4We5coPCAfzFe1TQK7WkxVKot
1Yc8H4vNnmN5gaeEM17Uttd+BGH2u/0Ua7R5j4wdUh+NBUCG1/vPY+8x/b9VNkbu
uo6xMTURgztFY79vDC+yGsjrFJBgQ7ROgwUrYlIo5FANhNOs3MSaRfpOxj3JWAvn
1dSVP1vHUeZAnQBDJk609mAiExacSjIZ4AoYvX3NsRkbeqpcgWI0+LgG9mNtT+mZ
4LsC4p9lPH+yX4DrV9VWlqxqyw3aT0+25mpOCHzRP7EHKeXcUq1RHQTmpxxrkHgJ
LfgCXsVgv2WYYbnJD0b3gXicbjhp+9CQFnEfO42m9BiG7J3d45Ee38iCQmdainE5
yTHl/u37CYrdyOIf02mPiXythJg4/Z+uYoKMDo+YTsQZGFycKQn+/kduocqr9dEy
JBemx7OwiaaOtnDpZw8I7Hzoga0/trWnzXcCfyMH4kfXuXoOJchJQvxKdHDVePlb
Dy7s+mgyKFCeQbJP63NpGkACKJMrNsWNste2u8TEBiFvxfOGzcTx4/xXILBll4VT
3CaTmmigBhCkRWsBN6Sa2K6p/+1Dyap/bd2fZSwhIwPAqLYkuHRauy7XAcHwQZS0
3RaMDxd67bfIyfgWIjzRjgW8hJYul8wZLM7NLwHIfD/aBBk/Cohhke/KwsX6sVFE
e5mjk+vEiW2EEPGJoO40z/Qwd4O+j67BHcGKRdMaa9TqnBqo/7I0eqSVfdWD3wbF
aTELR7oFEfjuXNR8bW0vFALixjIk9aEAt8Nkb1RAA6O9T1GaqayS9J4IzW4cGRuj
RRGRZj8MXGEU4N57lBEYHv5GUH+XjTh61sYF3qOwklmvDDl6A9bZN8/NstT7XxQ/
Zs1Yx6F054Rh4maI4BcsxhgW0bOph1fzVXI7bHRpJY1L7/mEWJEF+JugSDREwFLs
02lsFSdCg1oDfTdl4IH6dWdTar3Ic2kPedGG47CMgsAnByTc30v1MZZil0JvIj7u
Oh5W3FmnW2bt5vBiYuNt+T/1BGUkchQsjZpmUZCdQmOqPfuAgkozcVUxZxbXS/1I
Cn63LPZGsiyy3CDk+dKkU+CRmOQsa0K6Uz4vKKc5NbqUflIB2PdDRku7yd3DG3aF
SYXR8rzd/ET5zZi3K+wz1jOmBoviZ89ni5D99pk4ibLlrlBNQU9zE97W8v62hW0X
4vPgSjPHisqBksyKaJ4KkZlQXJd5H4weChOpSw3UoSGQ1PH7a/Hv/AszRdDEOTof
M7L6t9yvpWQz860BCqsUJaPR2lOct87efx4gjSTmuphddh/8x+SUd8jFRanMhpSy
0piHY8A90pP8WzgK8m9XIQCeQuJmpa3ySQgzx1f2jJHfc1YDH+LOUblH3dnvvx42
pCggtXTf5FPOfPqKXlsFbmCgsSfywfKNrY5OzizBbLo+6oIMJUkBx6EQkCJuGW9S
bQfoiF/LZ+jiupmy4ds8iKSBSTRR+ROGCyeZMm2PczTKDX4ywpLeme+ErWWWLpfo
I80BOw3R5C5tc0wpx7rzXEBtbiPWIypse4MXfjAADXyBwCJcdvLrloYzjPoj0Tp8
8TAHOMfMrINxHeVNCn5iyrSNzaFL8kLr2t41B0Hyoepc96ISnzyD59LpcQn8m80I
AN4If9AlcL+v8amw6C7j+07nvvpTj+ORsUPouIF50mEZzyPmH4Fqz2bmpxLSl8JW
oJqrTK+M5NscYWTZ6C4356glf7agNfHNjdNo3lAtcZKSnNPOfyot1ZwdDaBDtai5
Vi9hldVxelvki4VJNB7DN5MIN8/yU09+rKk0dwcfYBE2WO+xGqIlnIdiXvMzjwk2
2CWWGh5SK7WNUDcC4heMcPM7Y3WTKuvRfFu3QNQP7Ct2uHluHWQQeZ65R+kFmD1f
lsKSAfJC1/oHuTBMUYnOuStJ7s/LP/qvjfV6GU1PSNrGmSCVSfyCTdzWpG/uklTp
Plm4TrHEytoK9w0KQ+vo8MRCvb+WnmVDRhzsF8/WeMoD459n3aVeOmxT5zjBrlAl
U8NeLPZIIwQ9T0ojrbe0JgjHG5V8Rut19lkiLK0NmosOvzJzdEvM4g/dCG/HkjqM
bRkPAqrKfzg7yc2HAeSRyHvUE9Rv7z65XQx3Q5HK8YUz2zEPpRz80cDSAQ+s8UpG
fT3K5jIVHrJPXjOyzUqsWgqa3ri1pZihy19y+PXFq7coEf7pvimnHOugi9y7LAyF
BLwapgBLG8IZHnOwaJ6qwrDVc/vff09za3pOqAFLUNCdZXn67Q5MPmn+zcdm7A6h
gLGSKIZuPKlpMXpQ9ICtvTB7GNB4SJDq7MZurIZfxiTW8YsD4fjUo7ggD7TSwOCT
a+f3+XXZmeHjF53ZTm+JnUmspuiQ+p4+tVZgFvs1b0D9/21aaCrZHXoRwWg2XU1L
MokfSX+l+TjAD3y0upnLPe6E4pY/2vbRDCbp25nLUcE3ty1stIAX+XwXJfP2GRAt
eVwlFebxuZi5iwP/a+9+OxJ4QfnD9ydecmOPMn2CHE69UALiZyNaw7MwDbnzT80z
8yzXxv7u+rx6mvli0KD0JCnPfMm+6qVJyYpZasPrp0Wuyd9Klk0gVw6d5vo4tX18
4hoM3HsMjTDe0D0Xz0w+jhOkwwjJLhQURqREWNp6TOXxOyn8M3eqprnIXzbbYxM8
IZLpeuzgqp7c3GpRGLqnIyk14RPTMq/kl3NbJf9Z/20xlbUOpTiCMC8YBZnWR7ag
OwAhVIQWgffw0XGm1OgK5DypbUHL+H4ZKdlLHRud00J/kz9xHVnv++oOXDJXf/Jk
goCwDYHWdIHSe7ydSpMzeNB5P8a3RBw2DX0LY3tSGL8mQMNZY7n4n55f30KMgYCM
owNyYKKWc5OAP+9QH6pwWuXPuU8p6rhDRVij1GKoCsZpBHqdYq9lDZPcbAY4zCTL
h2nSSFuQTUdeJ3K+LBgNYvxNSdxzcJGIw3yALNKy2fR6SdzE8mbVLs9oST8nLK0s
uPi261JR79kHHgv1SY03CCRqtyg4uAMjzh8aicM2r+ghd1GduIWvzocD4sNA6IV+
7LMBDKKsHfn+qXK/FRt7lIfnB44as/k1zP4wOT7Sq0HbSgPrsphUPwiHiqrrkc9Z
/ABBT31yPWaJwJG/k/h2UWY/ZrRIU37JUX6TyKQ6EkUb0BvJ2cQr+9cjaMyCo/gI
2JpAD+Idmiqs1J81lbCygwaUB3VnzeXtXxqzelY5jUKvRtKHPjbsJSpoZamA/7ul
Vu6dXEvklt7fOeIyNq9zVVVkjET3VllQnH2UA2sZDkUkvPRf4jsT28vrDLCoijej
SlHVkUOYE45f6fRHnZh9wJsA6IdB7vhzIZRLU1dn63ahy31V7BS7FZnOrC4aoBdB
rS1nur3/NUzQq9TSu8CfBX/sXIHzvthm8krlu4s2ByUsTI5+Vviq4LwBqDlj2/Ch
P7ZY8fVjX9qsX7dTjelrSEwZDK3Q2z6MDSqmY5Xm2LlzJVq48Hvuv7LfG/i/6tZv
sJvrSL2BpZQ6gMisP5RKoAog15e8gc/B8Iq4gyLEYKs1izfGG8foXAE/kOvFB6So
KVtBgewVM9fmjDNl7n9f2BeCitXKQoob6FxhzNrUXC9KfYgLnNTGw6Q0iFkEiFh1
H1VZdCEDzwBukp9fZshWDd54VfUgUZg0CrRY0ehKbgnjVs22w2ufDLYehH9bvgYQ
0UjBN4DxNq85Xi4GQHpUyrj4ZMJlNIc2REpvE1XvuTUKPDOLWvVRbEXHu8BDP8IM
bqc6/5MUWsFNSxCsU850/Kscw+4yxEGH3nnNNUZCCiW+xaBBoZeOZntnQCkPc2ox
HYFijIbK4KvAYP65xKM2jijSUB12amiIPhwylyUuqu0bDOpetOvGwpNOGHs6fvDT
oE/NVVL0qEdJp1j1Gz243+a/4hyQ24AYFtpXzVwTh1VKG6moCLWIkElyJ4EdxPWj
dbLLA0TKPIk1947mdHVwNnPjI8KjvaEabCQB1jw90l0yj08FRNg1Q9LPnRPnDr04
mS9WVm/tuteCLLeRykriIBPtq5NOAslejsvUUk2WSiYzeQwrT6i9YKdDkSJ5YjmW
OX9RMKDmOPwryc64E7Y6job22tTPYTf2P6oRsj/xh9p7x9p9QAZfssODIBrWdtFf
mI1xdFYMM2pE/l6HQz6Z2HjA/AXKVZpKHKXONjP4ANvqCxIwqDEDduDepdRFmE0e
4tQJbitaGSEByk6B76kr3vp0uDLKD4gB3sdSg2oVOq39FdQX/mzvUPcedrVIYKo4
elMH53Dhyn/jQkJpnEFH9j9E0qHCkQgy1Z1B4iqnAoWcHhN1XHWf2CYOh3iZwCOd
EYm0Rh7/E3YTKL/3xXkST9d3exrBF2MLzc1yGc3tZDrB4hIQq5Kgg2lLixbgz638
tg2GXHfj34JF3V5XzMySBrzdPfSP9RxGvY1ecfKiZXsZ0Vef8zyI+wbZ2gav/BFy
4vZOnC7ZvrDaQhNz8gm2Yg98rfJ603Ml9CupgUn+Go8FfXyDa9i1bbys8Sc2OM9r
e49E3XSdi+OYC6kerAExmpT+9Yo2dxMK7CGO/pjV4Uj9YstW+8q0trAxyWTLvCFN
+g/+9knBVKeTHDoRKraRABeA54d/Qa/BZlpr1c04FUArpF6EOycxPZl466qFu37n
urSD5URnz+WW5Q/CUICqxnC9eXps5A/edIIuYPPZjCPGtb5yAmZ+cktuZ5sCAro6
9pu6c7B5JinxLtLrN6heqP8Tks8T1TpVyHQw/tB5uSabszwTDAhQyyjOYWLnDrXH
jr58eMsyJg0p2c9hEJRoUTji86OCYW1sWXcJAZh/ROrVTcWHoQLyY69VKnvmO39u
Jyrwjvgk8zQa/Xv/chRzmP+TElu+TNQafPtZ09IFc+shWnf/HzWSBe6b8wUfFhzh
UP184lFnj8MGi+azs3OHzXv3LQTSnME6awagFF5Wswl+tIKMO7ageEdNvVFFZc1U
KNNaFKRTjjDaVNxyzyjaDczszcq4CEEteL+gqtJL/1Y3wGGj+oPT9RXO1+0etcz2
cyUo4HTBfpD8cU6aKrNVRfVv/n4TjLJROkIFnEumuyYUeAJJAfiLU2lh5wzM0+gX
gN6RvDTDV4t0/5rmFA9N/tmkE73tUZjxetLyf4cCQX0lXDZpUcKtgoZhiK8cZ6Pw
9rEBQFRCYzV1tZrfSgVaETu8nbmDMo17fILEOJJznXpMHBDjirQbqNTcKhw7zGas
937gtNhN70XKxYIBFTsFkSn674GJkN5s6dxIrKJ9GBzkbiO1oUTe4Tk/VPUyPkBx
jjPdlcpj6BF7wDkzxMyn5lan8+ww/1EecDF1XK7/8mTSZKqThglgBZ8LE3gfFvli
V4/P7uH/OTy4iHarUl+wKzkwTFS0nQHeWAn6mBWAm11swn721j3Q4K/vOlpG9CnS
MTmXV9JBTAHdA3klk1iANsPZgGXgEHphGCo24cvNhL2gAnqf4qc2b9ErVNTMszhD
jlIcEtp/EPtexghM1tHfkxKaUF9DUNPWVWHdtRYohpHF070qMVuTbLhpqrxC6AJ6
kWXyi67DKsNpnbOu0PD4xSzP+bpSlnBfciyAPwNer3e8NJ3b9q30xZcb4/YNqDeo
5be7sWbG1xUugGNkZn8m5Gi4U3jwmxiv1TWqZFgyZBUSm62AAX/NNmsPaejJEjLc
TzoO/jPmWQyiyJ0x2EjwUP0f+4IdxEBPUKhgVGIhyH1iAt/3/Hjz4DBx/sxI/DA3
2yZD+AZ8PR3Xi0a08wuwaD7lFWC1uO6yq7UnvWo5IO4LCB1TGTWI7cL6gFEIuGQK
EUrjfCgJ3mqpshooN4V98UEVCOFdaiygDrol+c1+4XIi15lKx6UHRou3wxahsGX+
i9KUjKG4bv9zr272ir0EYmu2Eq3KEfHrkkv7pjQa+HnhHuiktMb1TA8kT0oZ1pHn
K5NUe/DE1O0HHDAlIH935IeV6lTEsS836zVI0cROwL+ECV94F1edJk1bxC7jRlxr
QGc8bfTGIfY6cA1eHfE3//LVtSBQ1J716niYxGTXwQSM1LdK6Yhy1tX6map2TDwl
int8F+GjPM9qfkPe5HriqdxK5ZzvnIw0dtZdK50MnLlT4hbHUwJDGLucwxrpcixK
hEUnHsBd11OXPKAEIOeIJBf9lLUKCnVphu6kOYKi3TClXDM0ltg+9JHVbDSPzp1k
9rbXB3MKRq9elzaNLMbVXhrmpQ1ZQqiEw+VdDhcA8NSDw2v3t5tKAn5BAlWoBDCQ
c0HkWNkE+fsTz5oTCN5maqs16l5jNyPAXEBazRq+Sq1PoK6PUNTgX9mmkdSdf/aS
JY6eFPRroNyCwyd8+OnuNxBu2ophSzHT6ISI5riY0UjXXrg47QwmwrU+ZDBNEsTE
GAfDKWPfRSpCyv1NGKw/WQfkgyR06WprFCeUXLYzb0JUXhprIZo0tWGgulfIA+G5
sx/82Tcmx5V2T8WEN2yDLzDqYjgDyJFQNXRRnQ5lhniDmQU1d4kIv58+gG+IXxeO
BEVpgz5KkoDBAV6ihHXdGbSTmqnd2wiBxkqoUVQZGIZEXYrPXjOHFJHsColbNWCb
yqaEaXjC+LbvUBiuIjIDjDQY03mrdrbwvPRGbinc0tn+b4Yl+Ea9ejHcxt8AHYIs
kGfOk+J1z8G4sENpUoC18gmXow+FJUAbiOnaoEOMf2vxhQvP8jddasAN4iLbITC4
V+S5OemOKbI2b9nc3tnEAefSTxTPV1XWlREa6Q6EZkUrGUqFJujlDoQI5kOQhBaP
WoiArmnt3pJqgVHOEJWl+Ch37lS1egDSBrtsklrQVtX7ddA/jr8X5kEFLLSqUxaT
6sh1LrPGyKpTdXW2lnHuFulx49iOqYPGShs8FbWM0sOcqeDjgydYED6liv0M0aNw
MAPJLEgWz9pMlvJ7v/Muwp2q9H25FPkXkfRIGh2TFAMJMkvTHxjbNTxT8Ouu2RjX
ozC/gtDuba3ekreMZ8VmYcpApkiTMtIWkxhDSG9OVuOqrhQ9Rs2gsJbPA5AIjeuq
QTfT9Yay+0Mf5EOwPyOSjA6k5R74GgA13us42rTH3wYxS0snbKLb1YblE93n/AzZ
IPTvoup4TqCGBj2CaAtC8EKk18SNy+txMXjS6qk9Jtj/dYNSHlzKYjoKef3Yldf7
cJomIifSO6p8Z4by9EKukbFGLtMM/wvPwpkPhWQymaKh2r98tm7Vo2ksZndw4uO9
bp+D0/REn08h3h+8+SWUayPHee+p6yhsrmhDy2ZhScGSv/k8Ir6iOeiDzXr25Z1L
QV4DjfGFQkc06DmQ8tS8k1OS08xcQNDkSWRiVQ6AlemT8hPlNc8IBPp3DuhxAZ9i
Fa1IMi7qFdeti1WiiNuUrdE88MVvhSK0LONpQH4YEhEqKZH+8bixuOvvcysI5W10
ZnSjNF/klXE2CoFa+ucMU/8SYYQe4VKMs4UvJEoW0tC4z3J4zKYXh1Hjm1u0EBZS
pZJTaF87A4VkobNGj1HfivoJp8QvtMnGpdzVwUaYQKK84D7MUF6GmAQQSCs4pZ4X
7Cjo0/iKRzuvhyRUV+dZng9vzgpl9Jg6PaTMFHClXUnNHv2XjOKqUkW3OPxmqID+
NPaRz/jt88SvZRqNdw/JpFHz9d3J5GwHw6w38oM+ieFW4JKrBSGxCiB8wDW3nNLj
u1WrL/7JYDlg/Bwjxs86OfNOIp8L95VKF5J59e72/SMtCYWPyJcOqRUY/YfPiWbM
zNOwPBEypXjhH/hBioP4VkUY6wZ9gChOB6ADRpwS2BT/v9OEOLOsD5Xtb8TxncmU
WTaRFCf0V2sbf6+kHzdUdRbt86sEPbWlK9I2SGG8hbRtwBxA8MeHjfvRL3NQPzGR
xHWcVpD0mMGLWJN6Ys60IpyklUElJ+HWBmlbqdX4OmoIgV81nFb7koTKUiPqNpXw
w/jXONxidEcNQjidGwV+d6dYjxGTISGEaqSxS9QrD/NH2GYt2+x3N7ScSOSCvgHK
FnY+iv++tr9cuZ0pAXLMhWaODItsquJdC2g8+MhsQCRbW45Yo10jZvWC+Iay6QAW
QC3/3/oRcBqyFHAXw3KGDGReOdUu3Uej/GpMYMjcG6Lxk5pBap6Q/OIVoZJMiZTz
D43VoJ9lvQylodloWD/ep92LgzrN/JLMMKyEOJcbrLsPhmaPvBYgah0rD861kvp3
6un5nxKvMu57PEdAD5GleoxuSKEbr0S/gbzgYDoXZsYeeHzMbvursJccivxViiy+
I64pVWk1ajRl1g1w27+THQtneHiXhr59w1EVMMefKpVefGfxrbFdJTctA8qeB9UU
QVPcHhnYALxFC8GQEAKnZZn0IvAFNXNvk+phuuCJt68/0AJ2D07HnUTbCDhoNPqP
7STfHviP9uZ/puDjhy2GysfEN0KlpA2ityN4/EW6TQwv45sbhqYkrs5bpNBIJE0Q
0crB9jpkb2cEn82S3lYDpn12I1tWCz9le07pA1AtlDf4S/0E8wyvD3sAJGJKmPbO
a+yPkGGEBuO9MWxKQdPTldOleKZD20nRXs5uSc+wWYNkR8w3/lyUfFvisLKLuZPg
f9hVX2Ygr3Do0hL8d5FempZ2EcQbR4NgoCJxVqGR7obbSeWuPkJloVYtUN7+etdw
+ptzw6GMcq3Eys4IBH4FrLKRa08kg1YGPc0nuXUyfWLXiSgr4SFlEJqRzGbcy19R
fNusu1spGQFgHCaizOhgl3b4vqukN4cWp4x3770FGzlpmXrMvJHGKzus8nfQuGzF
IlDAl1K4eUUCKGe+lNRy1t4COFNDyM2DtJM9kFHZbd4VKl9swdaHlLs1XgRnq/U9
SQ2ePnfrfVXYUwM8wquyS3d12bi/RBzR/Wa/KQFfiwebq9ifVGvL3GTxps5GYIVg
h4Wz38kMNWoTEHA0cUP7JgV5c5lUPTpbTTw2fl3BMojWIoYIBCGtPXHLHNeycNu0
CvaPnvDKIjv1v36tiZ7hQoBg9m61xmmnkQkiQrFeLCVsQoY27bSGAuhB/AlDEsX0
R6ypzQjz8i/wgg17THHaBSfrWh0V/iaO4lnIUXLAnBdCjcFVEsO+MAYcjRKWObhD
EuzRb3O/ziXP+cppDudCRDs0bfGTnkEuT4N4rOh0LgpWCTjvsbDVaCvVXd8q7BDq
iUDKjqzNcvncjyojqBuS+99VnQQrgx1SRwo+xoaZ2e7T27FZ1fmzJD38Wm5DXwVS
hyXPThqzViJ7ZTkzFx2syLjTIo0N8wmTZ+mSLe9nrev7WgBm+8YBV57x3WXI6kxY
WzUEuPIDegwt0j9xlc801ICGedvkuC729xVlk3IVgrGt7zsb7HxiYxKS7HqyncxL
b6GiCK2t28z61h/P0TkNewYW9q1AvvB51IJRKy3TrrH4/1rDUzmXykcQGiYt7uno
3SNT6LhuEvhHM098KhZSbYO9TuX6VV2FH9OEjExddDNncjghjAeR4TYyzP0BxN2T
Xu2mpKbrQScsUS2r3a2nqWFZA3p6DasTkiGE0hBLgBJhBmzCl7x3xIIBrcux3ARw
F1w9/cd25ZIpFsGguTzdUJ5DQUunC6TLbj6Yxxox0TvOZoynz/z0PFF68/mtYxMB
JGklQFBtyu5E8eJhOAMFga97C7lauhNfOvuhB9T+zHakVgxvOe/NI05v/s3bw6yR
uwmFkpPQO5UOFO74ZS5vi6fuvDkDSXIvIbjW6/fMDKAlTJfDSzTVloU+0lw3kION
Z7/WmgkiSm84Fkt3sbrmfd2nCPYqiBJ6vRFXJkFoDTS2IR8Pl5K2d2cZV8Pk1e1E
23YUyeCWc7CW9AI6/ot5Nu1r4REozQE+Nat7xT47sn31aA8POpnv4uOZyfhH4yEc
zewQLVYOn/EdynsPA/AqjA+FRAPWkMvuXMneMp7zlH0f8QtewvCURWAJ21zFfGYJ
pkhbk2YbfvgX7bBfSbfxdxdKJBhgdOtxYHu4QqlKkeb3b8eiSdWSXUkI+5FKfr51
B1aaC+ztazwClwQvMdJWBSw0TQ/zLTyCoV6Ap3ZtpBx+wZGpY8h4qH8Bt6hc8uCB
PP8xUaXvsG4/QTv/haKHxUNc53GrSE3Nu2dk8XkdPyQq2dHvaWdgfUPIKQ98qORV
EZ5xLBLic+0CiOo3bqA1wbeEY5YC+HdoYzRUofVJ5SRiEWo7s9nk0KskPThxZTpV
SaawzSkaPZEUtWfnYBVwr6coUeSr48LYDELS6SAWsV1cxjHcl2CEYlC9R0kl7Yyv
xgxTTNlwyEhxC2HnSWwRjDCn7j582VfaTdygoHd/r2zxpHDtDXXB/ii0AaytfpEj
y8aD1vEokG//DMMqQZ4HIzkfuwEH/DAQ1RC8OizeUp8PjwC6aiHvcCw1otkU1Ugy
2/CMWXdmaupmzeX+3Fxi8Kkb/+xbFldQG9HpI9G11US1TubWsjalCyUFH7z75grh
hvXIuSVF1RTzwUe4bxMF+MqjbWg4NgBGTzvRBdmxbACuQR2Q8o5moZ7H5h1fdaYE
3sRobm6xIIgh1a+q9WyLcdxqhltdvCf9zAMQ3hPov86/mP68dUXufsmX4iFJlnnn
jniU0agval5G4MXrhDkIQ8CUhQKN4iSDyrtUFyT/ErmKRYLcd7LzhGnKfU1/Dy6F
AMyHCwwMK/O6c3lOCykfk3A94ZTyhLCTqkR3x/Npuz7anFZPWFqwPTW10LzM18RR
XuTvIwWKWlQSv0ZH6bJvcrZqCMDuAPL8OWOVpUhRx3OnYeboBtw4h3Ce0y4OgPNB
VkvRj4q9elvvbL8VmJn9FH6hZZA9aPoHM1vDH74w9ehvRwBNRSS8TFlpcS5RwyOh
LXAYz4CvJcbPAhtXc+hG+WS80vlZoJ7LrNblFrXoC+NAoji4J25Pfa4o61P7oCuu
ZN0bsOmQqGbcjD4YIFIRQuxX+Skg5Vk9Nwy4F16x3MHEuCxVEGJPnlN+wqjyaFFq
Z86IJU8j6rOA6xqRPfH5ArPHUH9d3grTHyLhttxqjHwWgLMF3mZ9VkHPdk+USnCr
fFBRQcRbRTi6QxSE1o1W3dBBXZqMTfC5Xy/q76sfv02BxFvH6ahBGJHfTyXqtnjC
ben41U+8rurXwUbRr+IniXS2+sfyTyEIC8jVaIKMkTatpR6ykTvKgY/uAP7drD53
+86LFP3tfoQXdLk+sla6R932BrRYyPPPUYEh6oSL/RibxU4QblpWvaCWjVlRu/Q0
5O3vDXutfe+xQdHHpQkLwHPaoe/NRCUH8vHik1U2Cqc8gvO6ulLf/AnKvM7dv4V3
WpCnc8bxemSjh1yBalINY07I7Ii+Dyt2fOrYCpOhlRkoCGvB03+2I4ddI3MRV5j4
ysNfJkUGrdBwxHbRXxkraP10c3q3y0UN20/ssdKNssvHCOdDa9PASsGfMkUVSxMV
0sCMC2vZRrCFBJgo+pTd+7woPAvcLykrlkVoEaaO9acowgV9JIPUbZXimnGLaiq5
+tWgDC97Gy2PE3GcitxqEUSyLIRvs8A36sv+F5YxWtsyNYAimM4f1vzJfPzYLSPB
sukTuvnb+RjQr6wg9iCyRhIsGAr5dSEc5MpK96G/T/M5K90irRpiZPkqaNvvfgIK
uEBB/n9cSfRVNMehTSKEt5GM8uucYMtn7pYZnSC9aeFiriddonDdIQrlgAjtNLZX
go2IkkDSHsBRJirC31SdcHFOEnvpmfvF1WSywcU+JA10m9LyziEgz2jyb0mLBEis
W/aD53FSklGBadTFuhK/k9x9OqN2E9Mb1ZxnaowG+mXwKce9rlMAgLVe/KwYVqzI
4k5dVIy2DeUUMis28I/Y5zsjPy4s593/hSDNbUOuS3ZYQ5TLENLeNj+1cWym5K7c
dIxGUiRqhbMI7LxfETunsoXWLWyUTT/vJ/cbkrpzZG5W2h77vON3Hu8/wrJyaKxs
cxLiJDQ4wK/JHdJJxGYTx3nSC8Hs+muXLkb+o8bI8m+b/Yp2o/JyPHuv1GlJJvG4
ndQc6tWkRQVxEES3QWwJaEe60txlPyw4xF6LRNpHgRlbVTgk1vWE8TVCbEJqSmYC
FI/1FlVLZwjLz1Tf2l8z/31NbHjknCC2v58/oorsP3qbxNKrgNQEu/GlhHo4O70a
7Sy+aJ35/rsdXzC41Ji1/RT8iSqR1JrTWxmdYWAH83ZSwxh8g8VpyDwTD01kVyud
1YBks/222nowfTEOy2thBludPhIiJN041SyQ+mI4uCW7SU8BhRzKrWR0eT5/bG5d
7XrwoGlaqnQrqCmG3vu3wR9IJDYV3bRvtPENr5d0og7sqsfIJikLrfZ79nbQisF8
SLLlGkArO2+SgCH3aCDb0a9+Kuu/f+D8Nnr5JrHToiBCfs/DI2aTnya1M1xJvsxf
q2+X4iCnskwYY17zkxJ+/6JrOODHuFuajGlr1nTbfhp8A4+EexxsU7pv81cGv6O3
RlRQE3+cxzW0xtfn73jBYcU5xyZuW9aCMf+N8zzmYl6o7tnluv+hLdhWdNz/uqnx
4nrd938Fwut0lcMpniWVR/ltZSm09qQGHZsAhRnNWmQjRbmrdNbMoylOF1yCEnuM
NUXhdP0ujMfs0PuVFHimzL2gIKZpUzfYduYPneA+seaGzTYS+6mb3HNb984/uouJ
D83Cb4KsDKkXH5j6wsGYEP9IKJ7INlVfOvEkQxRrC8asKHnoDeSLLnV+HfaH4l4+
yT09a5+g/KSJYkdgWzV9OSvUfJWzC/URjufAKrcc5sqkEq3utb+W87Mqh6ctNcHB
HRz96Yd9LBJezoV7pQxRPgPdkl2Wc6lcT1JK5ZFQKxdeydg/HAsJ4Nn4LQpe5EOS
FNinZrbs1DGTzSRfZqwmk7WnNYIbLFCzqeIHiGABMjpqmzOG+lc/hD9S2rEcG605
yLGmkAYps2vqcef49qrY1sYY7p1CRHXru6KQrd1yPOEv7yM9jKmO38D3ogVHwp/D
pnHMm2pZGudiQ4OZPAVoMyJbG3qbTUNtOvB7z2FErYipZY4z3IEVd2A+aNy1fs1u
T+Xs54Cz3okGSGM4hOS4wGKdHzH/wXBD/EwfIMt+dwgVJdYcnHHkIlNY0gS0jV3w
3BNvc5n2EuopBTniaRlMimoYJf8N111AyyKWjmHPq3F4Kv9q43ChyHob2rIF/qM4
b2YbXd6mD9PaNzgvupg3uAB805XmBFGPevjSXUVT9tK/bYDpNN0OmlMfONaKIX+5
0MxYUnS/Km4xx7MYGgT1jP9k/Du0rtJLxa1J3lZxPmHEhl01B+yjVuUtUVdTB5dC
RVYb1sX/cpCOi7TOlGzCsNWU7Xb7pY8mnoPNPFqO1To6V0IlIhEdMRI38ZJZ6DDU
juT+TF2TXt0zKOCx08Ls2SD1WqpCGc25nV/utaSOKg+eIn/Xlr5QKUmM+jLbnEAJ
MPQdCObODWJocxoDqS7qYQ9PfOBCQwHtPCyUBqJZ/ZDO99ZJ6H/SJLhSau6PifCP
XRCd7qLC8FoYAri0mwtOPKjXaT0iVjEteT5yvFwR7fylaXIRM+XlpWVXp7f3+u1k
YGU37uJWtAT5zRlM3QVbMk1Hxg0h4o+Jsf5eX9K7O7j8Ldk8xzk9INOqro99zBt3
eVdZx/SbLZwwKsI7aotTfmujKEgkI1l5SQAJgDH2q+9idqeAFYhAoQLyVoPHK8pZ
Emwl2CKaTt03dJKMIJcNzVoJii8fX8pUpLXQV8d4AlmkEfORmWC91oQK6KUiUMOf
S6nZaFIlw/JCFIhSUwVGresWHCS+EThy273QiOHirnGX/6C4Wy8dXjZPT6KFF1JF
IV+/COKLP40qFnuvWE7qFzZPqPSsNXN+b6fGncueLfZavMuWVGFeuTewT3lhTOzY
bqqRIZs+GRBHfq6DiD5ole0bhZojMndtE3csg/DMQKoD6HLyKBseQCptXDyquL4H
TFQvcMQe6mBifCc6D33eXst16wp3a6UuMaFFQmhJN5+c2QAG2xG/ERcvo2hi5XYS
jOAjPG9rSmnssZR7Wj2+YbLm24wtoPWJl4r2etgRnwarMkTkT/dDprn81HhYkrtM
yvsQkW5ZczFFKztHoz2jkWC60rTY/yq9/VpnzvAVCzhua/vzM6ExKyeo5bsGaOjL
x8ieK64GelkAIPdQdOt/cSAtQpVBlECckLhi9Rro4daJBjGsjrGVS/Sx72IozT2p
ZUM6TDoZ3/MCqHGu8XHzZ+DueRMbgpNgA28EM4n/UVYb0qOgXinaY+9PrTIGrgaj
hrF257SbIIIc7WYvNZZGhlxDha2fMs5Y90303J6LKX2+KNX9XXceRZmPz9B+MjEF
OXb/2RiS03amNjB0Ahh3aEiF8Ewv2NME+z07R8CbTF+CQp7DmzvSe2IY8nash0fP
B92jZhhq08lpusvQ/uJqxxag7mYUiWpAnYr6Wm5RWmyh0DMPdqPxmrE/ZuG7auG6
Y/ZxXUaWwOEzzAcmyc8D6l/xGK8iLmV5D3JdaYImZcVOIYAIkWUz6bMdCddgVYap
LHHjEaNxtwvbgQ39z/wvqW6bAxBJKy0bsS1Mur9GvnYUJOZZfX1MG+2w8MGKxmUd
SL6sdYAcBYjfaqIQwLDxMEb+dWFo1cT31+BLyJNewCs5JqHIKb1k9n6kvdQUZZOE
4YFp2FV6FgeR2tud2Tr6I6Z/rWgiemYHz0mpMbJ+OabNW6jjqiLIQTTeY1lbGSPW
M0WgBCUObxkvLq0BNAGfKjdanYJ4hO69ESS/aMBKMwalOEFSndEdweKywB903+Ma
hvEK53osx8PbFhYiya28b4npsp/1SXbbZa6JJ2eiqbNL/T7886ZaK+dtUsj0XHrE
XIK1UvDwlBnyl/h2cJaB4+Zrk6GAjYLAAFQjGshXjHirrLJt7uoDXmjRfF30IOZP
v9z9oxsQ5VP2SRlZ9XTHQm/Rk04ho3Q4i9aLxykT6hiodVUlPCEWWg5WOzrz4+n2
BlnXX1K+aqOodmQkBKSbcqtneuf3Nau+NqxQggyxiJa2TwxubBC8GOs/ZnBt7m6U
bxCD7kq8BliSWcTGTl3vq2y9O4DWWpU9w2DfzV6QftNCMNfpMz9lQrlzffWC6Z7y
TfV0CD0pfdRgBQ1Gr/DpoidunOK6NvJLQ9ot34VEH9Tvur1JsiKOdLK1e0qjeQx5
aGoAskobLW+TcQXq+ZgzMb0ABakvmsC1Wwa0TqwVBmVCvzS91WvPLaw462CiONFp
AUQX3Xu2ZaPcqT+Jzre/90NpW/AEVH1cAG1/oxb2KJ9vAdzMSx0lUCsAxDAk55Gj
XE2y8qVlbvvUuI7YOhMwyE/AN1epfVqcvyZpIxag+bB0hE51ytcEoXlxYpzOvV8o
U9t4FSqHGV8AxzjKkCs1jKXVL6UkcmJ+fYMPwzMyYarVBEpoVc8qJG4dQZPbBEAO
BVvOPOFboJSxG4VTJdTFMtaIXZJpC9CXZqpCosXPATwr2mSY3YUGXmYaBHEOmvll
/DlaZ9crHB/KNaWjvse2ZZmEBt9cWobyjbVsHs5qxnAb/nCIHTsk+6sjfwchliKJ
UmJ8T4gYqCOCmQyRhmMptN1sbT3yDSHlV+psyBdWikjfnqToO+5SiEaeLd/GgWtz
EbDx1szE24DH5e4SdaTxkAd+T7lwOtcTsovw+awveXMcekUxZNPOb5bQFmgi/4Oa
1MXuJGEtOscUUuFSAezlJyTaiCEkjjPNOr6l42qROn+Pf/2icdWIkKKCpYla86Bd
g5J4Xjk25ka6MaFHff/8YBS6/9vdiRlLZvJl7dauhm5UNuW/a3/xQmnncrop/v9K
4x+NaI7UMyzRhP5/kfZYI2tlxVKnKDwiD/hu8KHfsaUh2e2A8n7Z0BxhSI4l75w5
0M9EoJcmYbg//QSdyLbV1giv3fYTkV/uECd2tHwgyU4tYFxQ9+6v/IP3bzdCxELk
X67IDa9/sqAdaMLDqxMadcZU49EG9r0obponx36nJrT250i4aKeoyRCBboyOhv7m
ZGen93T0PWF8mbvgcKqJB4rZTJBBlgqRsU4cj080Xd1JKUeCLAaUflVNe4lokJNJ
Gn3MheNGKBUqLRbwVp6LEjmnwvaGkP8LAbVc7cEVUYqH6FFNgkLepuVsyLVK/0Jm
DTQ8Xq2TAcKMX0HegrQAOLWZqLK/FAm8wntPvlQtmmkGxyLCfmbhmarOmfvReeMQ
V8hPSf6cmTifko07egjVooz6EMtLpTUdkxhcw64RAy7wEVCnB+tEQjjsqXnSmS+2
VZ2EcDfJDd9t46xDnMDDuk2l4Lw1roAIuNiMxFQRKFafOQb93wQOlHLDTBCDcWeL
MaxMArhIodofZjLyMabN2DCGUam6tOCLSBFvfuOKRrxKJX0hK+szO62elN3fJgDv
RHqw95a5jDmSZdq1wNhDGACECuEf1JUw9a/9LwsH17WKPzRwSWvdf5fr6Z7Y9GSY
j9rtFpUVf4EdVaGu5/fXi4UptjQ2PPx8pxahTQjVrWL7lm82qoF0zBHM/wKqOBjQ
T1wXp0b6PpTKsPcYs8fMPMuHVEZHLUJzk1bkZj/yBmgU/nZEw07Ga5R86PS2YJnW
M94Br+2HqYZMjFSn6CsyMLz/J8Wxdkbn3dNQKHBJIJ4407SCeOxfHNQk/jeZUwDK
pqHkJ6vsofnSBBdET69UfkukuIFhOSmw5r9PpjWn5DzX6oPTYPE7fjsDkSdkwM7/
EIHdYpoRCr94D2UIZJCvyGRIzSDWDzcoaXAwfBYjMXc87zSReGeAcnTzI3sOLWdO
SEjopWcnQheHyOvrPHJFTrKh+UmOpLO0dy3xZSXcq5jfew8fVUhbdDWy3DTR9b+n
b41danyZAgIaX2QnRZNWykJu9EDTc6WmhLE1EBhknJ8Vu4YTpRrc4/V93oW9yq7W
9cEsHKdopfVCmPRcq4HbVOlikAIPx5DibN+qf+X2Q7llICoRGLGcEmPQzU23Bgq2
k0Igp+0Cj5g1Latq4AUhZ0Er/4f0kTq90lj4YGA9/Rr36YRB6vEaAYhc8ODCQpmb
O4k1RAEHK/HPttBkztUiVEL3d9MmaLhGm9ZXCIddfQCJGJflef8AdPLO3ccOIMrp
8YbVDpVvZKzDbxzdp8Zrg8dEeVj2jay9Wq9ooyvqDH5n2VZcEw7qHRbBhMnQIpBy
CAepTa8xL/DLjCe5sS5vb73PwfuH82mzpzy1PiOcjij/mL0bdr4WeCVgK34YaK+s
ONWKylljel4BbzajE6SS3vzIvdBELHxReO2Lyq/fFY4kfc06K8W1umhIDBk8/Hbg
QYG45AQ6RhvgLGTpqdPpTv6OfcxL70Nrt3UEVxxOqfqv1wjLCZXFVv1UK8NklDxC
aZmsqf26hsa15ocppjmEpnQgu6onma5bCXZ0WLFm+ZO3hW4I4TkbQbGSdiMOPIF4
WbhaPMkarL5dtwPlpeg2VUQzgY2g2DhS8IEy9NQj5yePlSThuDltckAFQh16Rbb0
MfdrCuLf72ULqiOkviKHiWY/3T+pwgY2hrRoYS5JYcjrfX8EMAdKdy3BVNj6ulS/
MmqFTls6mS1n7Xn9fxrEZBPxHoR6MPa7TjrTB37wR4BQkScwgonRVosTrM+309Sn
RXh0UCOeQVzV1J901H81LBhG8cH/g6B5Fv+Wf2gZwqvLI/KQBpOJGZn7PyMFJbJI
OzmsLhu+8EWGAC9U3YWS901cKW4R+hWEfOyruQbG++zRQbSvtYybxknqpDWbhd0H
wApHDQJRuHcdllTs+pxZLHkpyI9YXTRVQ4G8zOcL8E8939KHJi9T1ojcrukQZopm
dn/WhT/PirRKplpq+lcfYcSKpRhajxtb0ZNo99uhlDCpC0owSfHxcetLW20SGWF7
vUPjI8xdeZBBhXTHk+V+KYJVboCjBexzD12TF4a0iCl/RUsGmKtzSufR3KDCTglz
HqSVbPKYFdb9GDmGn0ViVsSc9zrcUCzQ54YzNgR4xoGhEd+RE0USB0nstVd4P5X8
0Y1TWRmGP4ytisrcpR4NOA2KJ23tolIpXiuf9L6qvAo9GJs3ZeZdC/fuUyEaLGaU
VzXxFLCb5EsA64JMnrXZHeH+nGUXFNPWBkZvLdw04o9Vz9kzx0nKqLp0S1rYpwv7
YdsugIS+4b9yJ0tilfGHqej6fWMme9zrJgD5HjSy+gokmHpFYQ4HzS3niWEbCVBc
exaEnJoeZTc0yOO0vpTe4yCq5eX1iUhaTM2QydLhimNfRrjWT6sIz6wkF2GUmMPb
nntk7T6P7aUxXDVAJuF3CGsl1har2CML7zbGrpZsoEPSZTJdNm8Nbyn1M7m+v6jH
5rMcj603ZTvPLH9WfmVI3g6pagsNcBFUMh2Zx2oFdzB6P7WZf0hdvQEaqjOzsgmg
wrNIknCjeFom84JeGP5M8enGaolyOkIivyD7RjNQ7VLZbz4241fZiNHHS/bfYgCQ
jxXoEk9tsVQvBYr3R5HL9stj6+SzhNiSg+VQGAnxdQ6jtnyzg2POVttd6XgWmerQ
EVHXuTL/uIfkeHYrvFR8ElwFFvsxHMdvDgO0NbM6oYKMr0P8xjEb6LUlb3eGIpZB
DEAjO24VaPlLF+VmHPbbRAgphx2YbSukLsbtdUmwsKs4owc+bAJ9XtpC9Owjv/FQ
Pj1R6CcOU27n+1tnmwIOFBiKosvC+OOhi/qbr8FT+vxc6eNXyKNbUtsCu5200sum
5b9THu1K3AYOxHdNehYwPa20gPAD2s2IRXmUTPoiqYnHTyXo/jn+A22tw/KyPwo4
kDlQSnCm6I/eW2VbvQJCfmIAUo4UGO7uSI5L1/Xb1mwF4zTEY9NNbr9GZ/nPO6ek
vSYj63okekOcrwGzBhVIF4zKxkcxCi66F++OGav8R1BC5x1WQFRrAGZqdxXasF9Q
d8prHe9w7MYyvmTiEQvmtgjmNSrBCk8PBiEySGjQxMvsWIJZfvGJ0WCY327MaKqK
p9D7EshTTGlXCblPFhXFmfMBK59snMPelTWQExKIz6W3qjL38MOcUlwch0O0UgJi
kS1jNenI0shu7Jz9mxd+5RKfCDpqhlu29nYxPzVXzcL9TWftqTGYsA2FsWRiyh6/
YuFvrAsd+8Uo3oqAZg6WXl7KuDs9k6NL1bFiHy9LrcbegVj5KmSlWvi9Z+RKdvP7
jJALlr7WCohS3t0GVberrkJw8GUt/KQENVDItvp6k4X1CsfDjjgpXwosjAOPI5se
Fo4IcsF9LXrsQN+vxhWPDa7kwhQMvTCFq58r723qiEIiNVgfQ+C9zmuLfEYAzTZ9
yKiF4kZUo5ty4LZhUtFhwBArPUbXX4XYQHWv3mmVce1/X37VghJ99jJQCZgxu5f6
fMKnzAF3Bn1dllfWxf8l0+5rSV+i5dXvEXEj382eMvV4g5ByAsVre32P3hIb8pfF
Vl5aYoQysj4fthorCEHYFXYDH96Pjx2V/sppUpcg8vCXa9jGucb8TUAKVprjgrE8
1pvhCGRKySrxV5+VQM9/D/LErnf0FEi2rOn7L4xhWNytYu+67o10N2FOOSX2phas
zFCsfwMnD6pAP55O0Y0yYXnK2bKNMc9ive02jQOJa0i3wxVS0dWmo51ViDcnUC9+
hKXf5apa8EQ8z7rqWrH05pMyMI62ACS6/BmSmpc8w9/kZs++0K+6PiQ66vzpEdYq
3LLP0eEKfL3Mk3CIJ+bKSkgPPRw6MZezddRH3nTr9mnu36kZWVtrWvvEnhSJLnUp
Od8WNr6kEf/QYNEslUUoH0Kjlrl2BXnsSc/qXm2d7zYG0mUUFFNctUUQ/qtWhOBM
yq/2OUqApjnTppFh37t1sMBzW+R3WA/yuvs1tljr3jemam3ZAD2Obu1xcHKrpRU1
31uLfBMmhvbuAtM9DVdNKgzo+/GM6lhBziLgKREun8DcQX5voT0sQuTeaFqrzMQz
8kWZF9jNbTLBy6cQ8EolrBjIcnKXeBEBG+1hdHBQahkkYQo93vYXdZw74ueuSP+w
iuRU68+bouT1mkFv0+wZKvrrvucHNAwrgt7gCYYEh0PF5Q8AfCf7qMeEuIxsqEwp
cV2f/0hgo/5jFJq9WSRH72f+u+YWW/WogcqBXoynpDplosb6CZe5ln5H4E+Qhr87
/Rs7ROxFYuS91F1hVAcVkPwCfgZUclDrSLOhUrZqz1sz+AXj8f1NSV07oONaOj5+
q+ZKBXbpb7z8x17wE2jf2ToFrGLEZTmYgw9ThbhUlXkR0T+WGYkirBiZJq13Wcq4
epB9jlKR3grxKqvCPsbOt2Go0fGUA91aGE4+ATAQ8yxwnEkydyl9kXsMl+WOmhRH
DTkQTMi0UVOJI/B6gS7rBWwEziU3Vi4wjxP6SPRXuh9fFc7ua/Fa5GV73H9zTlSA
YwuTl6oulPpYI+Tz4ZXvioofepNORV4FTURwkVDgNwnWN8dFWLQNG0CSGw6t2/J4
eOcYidxiyHR6WjaUNzuc/2Oc1OZ8jwS9hwgvSWnNxdRXd9UL1q3EybJsDM7WnJpb
gomAUUfcoBGuKdY1TEqdiHZHfi5sgPmVt0Ymo4usg1Ufi4Qr9CC6a7ISFN6AgXAn
UiMkQBUgZZpARXeJiEG20SSq7299w5J1Jg8TMJw8LhMVHIyqzxuCZjRaXAQ/knyF
74/kUe/cacBa7k8x9xiqcCc6Ib6djoRYpgTcgmyTnHSCki+VZEe3hgTC7nlMIdv/
JfTISIUsNyQViDBQQgE5VMdCdGkCF8cqp226jkSOgE+4WkAzxniCKEqfI4rxnqmP
4FsskaMNaN1tGdQCvpBPHM389BOiyc3jOHPUh/M/e7eaCdo4eK8bgGDhYTLi0Xnn
b2u0oA0JJHPegLT0yiXN0evVJAJm6rl9KrmQy3dHUo+gZd/UiuRL3btWZ1WyQmKp
JxVptc+AnXfFPPe4vkABjUb9hXdSK+o/9+oN4Uu9i1CnEPjoQa9gpmM/srPmAmvO
PuEoF9k0Z44ZC7TQJNi+oVxd9AnA/3fnviUo5BaK2r0gsW+u4104k7IXVCg4Q4Tr
GRYfltpfOpLZcnxzToZ7WbUlDg/U4NsndoayMgNmPPCmSf1grW/zGA1TePsdMqS6
XzrahXawBoCSRARC/6NWa9kI+2WZUGtITCKjqlj9UDrcV9Lt2nrz4aThes+FcCIA
AqiqY2CSekht8NXCVgjvy5HpYe+YGbsbJg3MQh0a1H+Pxk7sxMahVroCV2zc4EgS
h1MnzScpgKnvcWyKfmfblwoepRJhhiNFFjGyQwJUZjmbbt1HAo8++s2ZwitkTo/9
uBMIuA0AUwA3/ZDv7OD2fzXT0flXACeYaBXddCkZVjh6t/YzktlLBab4kJjwwjKi
NFTq56zJR10pdcVdt75FUGy4HUZJOB0blCr0teOIR/RzqnW+iMcuarUeIant05G+
d0YguDNVB+ISYisN7MnWxTOd3L8Aawoh6mW+v7CYWGWI2/4IkFJPAohf+CX3Ex4N
HDm40ohvpXLz8VVwawdgdVCpMfYiiU0hfKHAUQkOdx6kt+gJYtbiJRe08cJgX1NS
xaeEwzZR5qaYSkMEXZnF0S8XVRP4l5Eet7bGf5JV0vIlYXzMpBk1l/ydfnBv1U9v
uuSO4aLPFlG+g1osFxll+iUyn9KY4uqRKpudkSskb/FIRrEu++VATi7vcv2AU+U7
XB42k0Y2XyHWKDUrIYxjnbwy0ndSDkuF9T0ijUhphKPcGpw2X4dXXJGnBFW9PHib
7k3Ir333gwrEkg2PB9ZKeLlC/mfE+MwIGcnBo8zyNjAX+i+jo+bq/iqQCVjHOqKB
z9+J/k8UiePazVJ4tr/X2yyrMJ8GiDAo9PdoU4/7v24KyIGTmYZVD3nbPU/r6ORF
jo/KLa0eB1jKsO6k4H5bvzmf1+Md3sPQTPDZKigDM62lLkAzc9yzaUJKz/fyVia2
T/QIxgAgMFxqXtLc5tedvXMl84Y0uHBwOq96+T7eIwkSYdD+MMBbb2QMOzG0wKBm
bkhGuVYVIyk35g1RNrrAFf3YqI+v+aD8ZlAmJ4+hWv5eFGFsqzgS69o/h26nhbcs
/pVnuKO8fq1S6uEYCQOK5TIXMSPMoq9J2mfC+mDDZdAp/bYYMKUTCrlhvTT6KBCb
9TU1sSt0QhvsimNceTTXOo2kgjyU8uxN9fZHR8R3bMomKFkcKSsO3Bz4XZUJv2xZ
oSKc6SlMamVPvWkyxBSoixTJlvJFNr3Bc3mxi8UYt4fOHbWyoekS28vmG7GPM7q7
QSGFCbVnEoYLz30ZtCLRCOf9cK/iPKh46HKsc/4u8Ioupezv6ZK+MMnAz40Dmg2g
djhBkAG2z1MacvjZ1MP2s4QHKSFrwZbDnsg0NJINOsyGFkDSSibzTOgWSA8mLMN6
uVuB2+KztLDbqZXhZCvOSKdnYsARhSY5pNkOl3uhEPEgX96sPiY26ox1vkyZMNmj
sLpPOtn2h2MoxsA+wi7yPuoESvSxF/zSHc+yyGrU6IY+rscJo+Vezn7qOCr6P7YS
MkCna1FjvjNE5fAW19NhawevOdOpv+XwEsZ/t3Q72o8I6uVY2ZM7aogjeSwVu0kD
rAo34y5xBOkyQGU/fwuMZJu6lChqVb7w+dnGUWdRArn67cx/ygOp9yQJmEsLyWT1
+RPKj3WQGTJTUN+HI5GieeWPurg55bljD/T1NBNzwS42xaG5bF3wAlEUJay+VSHU
pp8imkeZTZXllOzehbouyq4FJ0HTm64WuzX4LaaahEaF8pBcooZEBnvAcMVSQGPQ
fm5i0+4Guv6j9MDyZd1si80DwVWruqdXy4+HkcnWVLIbpIrzPzdMubwcLuyl//J4
SNiaXjARxnq5r/VWWTYv5YQY6HpxkbqHmNtJ30+o6+ztigJ236kI5w7LrjPW3Wfq
69haRLTIUDIDA6jFGaUn2e6wlYRoBS9p+OCgcP8I7NJk7Wic7OSx/4JLdHUaU6dy
9bXCI5cXo3uhEtklDe/rdbkrqteLCSsjGmuL8Rvv8bdDrShMJcwO7dBh8XaSxWng
xd+PB6LKz9kr09vC/p65XMZsg6NwuiPKZyB+efsCfHFIzBaWFWF36njQj6KEADmO
dZeUzrB2vgoQbXh4nKHTaf1PgrTlrsVnCCpZObHUHzuiEg+H5VtPlW9fodvwUN9v
bqvUN2Kk1BJFgcKWpmsw1Xw8q6D50Ym73A+AphsB1Lf5ugTJ19R27gRgoaLoAZA5
9z13FcYf/PW6rnOpVukLaxlevFn92yXeK146BinvHzZP7u5OK+C3aza+n8ThUxdX
vLjCiwVgNqB7ZCdYm5h3/9OHjXbRxNHbnWGAjWjaj5kopBFZqIN99yq2UKh+ViTl
poltPwJLVFjAdqeHX0gmSMpn6UD+Zve/MCgFlOGk0/arXFfo0H0cKQ77K6c7QUQm
9kMipa0lbxnRVom0DxSbWM+LUhGvrYAu/kBmHlQC01YwMgL0k8xg3SfSXsZN6Xey
36nRBRVm95PHPyZRcBM/uCImuHI6fkmcsu8cA34i9L0UN6MVOZYpI19IJ/E9grm8
TTK7tweKZ/6+bjvVtNd1qFme3KkB0hJ9XcXe2YU+P+6XFzIKzWt7hswf5cNboGSU
LloUmNnnEupXIYVTM1kvysicZHsd2sfYWMeUoaEq3A6XML3Bwc24HJ9Omwf5dzOA
Urhyh7oYGFgPO79bvS+EVAyUHwEiNx5LrbbJe6okEVAUFzEaUQ2ZiI4MCxtCOTQc
4YJ5F5FWoQ/MvQnWB8AegTySz3TIMnSPRKnLTsEdU/S/sikGVVbPyKvFe16w/WDz
XQviNrp1lAyas8hJScuoJGtxXKHckZsA775PoyP3XOqHUgIAKj2LqW7iT8zwjuH4
17/a9g81L8KNaGYyYmjTOmVI44/mTnuvO1Jv/5RGv9+lU6y0GMDoZ9qqniPCTp/Y
AB9pDLV5tCYeZvT//lT7vOwv7k83T27MJyi4O9VC6aYfqKVnwld46qH30sMSi62l
BKbWH0uvomkAvF4q3vm1HMEAy2xzLBRFHzhEOn8RE88FD/dh7IVwsNOtiREA/iA6
r9WKisZGSLq+2H3RsDwHWGyNBhze89tJ1KlC0g5dUlhlxPccqdTKbcDAKpFJ37/i
mPb05JuMkP0lmWkw2M6/V4+Voy37ed+HJO3hNhmjShjmfPKAdBZIlj5EI+g9OZYp
zvUj7d5L7B3iYA3sEmTBA5hPI2ezD1hchGFuofGMc1yX40+4lDJXgH/AMjdG3tlr
ywmrqHg4bgIKQyNVOQsNGp49F1d4jdC2zDGy81UfXcQLkjrJ4EmzdmixLA9w4asr
VFdxe9eLld73Gs2NsePs5UNXUzK4Iwh6Mn9daW+xxFE=
`pragma protect end_protected
