// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IUAKGigE0NdUW8rX2WwEHeBeWRdA7zQQW+JKZ7z1TtJJyB4HOoidzotdevbUAZaJ
gCwSO4Mx4CkJGSnsrNhKlTh4fXBnzWCZDUVyDR39u74gAoztlybHEPJ95kyWlFXD
eIJQdbBSOOF+LNNKo/eo5P1FDMy0i1/Q9lH+yYgJY0g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19040)
vJ+yKyRE/RqfRVO4ts+0niYdWUohKPd9FNEJRqz2QhtLQJYdlWzAyuTcqGNNJnZm
uzYEfxVejsIqx9rR8NNb5QoWLnGcqmu7Jj6yMwMmOiaRei4sxYow88aqV5anHrHg
Up1ZRofZMEA/DwVXdo45D44L0+0sQLX5XDBvFV+HT5X+npxz7Gbd9IHP3l2qgHuv
detAvNMfbH5Tjcf4tqjO7udlyc4PdBODv0HE7Y2jFHPbS+68E2Dqgcvl8zZkjcHd
2aW0+Npoej6iTqWaQepcGFCFZkMPoLvqxcWHqW6sUhv19iEXK3ENlVgLXMQkqmCO
5SJSMrCt2rK1Ik+GZpj8hn7R0YWE1uDRHXwYoKNPmxj5RYvS6+hwaPMLN5oVX6Fx
GdADyCjHf/q2hs0ztkN21byj/TCmIc2quO6OP7kPV959S/NzZtl8d+BaB0Vy5s2n
uoYYPcG7WoE6b2R0Mor55IDDQmgTtL4Q+olCTSYwoncAbIFL/ilOpbjL7bF+lpkV
da8TdOiZDnD84GcSTsGrlJanBE+ULfTGGfKZM6LNoIa+3XHqdlCnXpAA/O88T5zN
Rp8iVDPoOLkMTWzVmBA4C4sjkoM/aMlCrpzEMyRMOYHroaUhAk8tBNCPaqkLAlWk
3kskocOYQ/77ZWdbp8JhJrR8cO7qKNAf4+k54kmvCHkjDQyr45OKQNCB9B5b53uT
7956YN6taW89kq1bbUbYsttlf44KTZBQ7pIt+5RY/h7BD7cnseLJVgz5DX7AW0gn
8QoWwfJL0rlIjikuBlaEqqyPfbjm2qWoKUsWyo3h1zXELq9NHY3Alkoffzbasf8F
I71m8//YViU+IqeEqOPy3rMbhvv2A20Rn8tJ8DpYgYbDzj2euzyyvP7APUweaZPU
vNcUJ1/Fm7DYpOKBONzvN51gLzEZ505BP5cTXoEkNUg15gJK2q0QGmb5fPBGJ6uL
atIewWqp8+JJ9DNfCwkP8k11ksUwz3Nz8ks58uCwHL2St4W9kj8DwcDz7c48Fq1N
9JkX63uP8ZIS8n17L++BzCwabMKfp6DYWZ5tsIjRSH0ZbdMeTJ650V3lPh4JdU/j
+pd8u9tiLybEMs/FN0YIFKCmVB3PV+NPQFUdgVGswAbF4tPDj3ELron4Oqr1FTdy
TM2FGJJZ5ZNljwB+pV+xmM/mFVOYk6AIL6qSga4eD2cfC4TYYRret23+OvZ77MWZ
XmxmSZO9zLhcNM6feEpoPlECJxji9wgDmh31obz1A7WsZ2IUdlHM7v2sq5F8oehX
JQcm7LrLHnFfpWpzvo+YWvs1FgROMWJdeiJ242wnU9AeoofOiSMZ2YYDHRtrBIkI
XuyrJXe15NGgJQAZeeeDet0oUPCXN/FqcpzuQ2ZrfQkktq19ZKfHKtSfE2g3Qqh2
4sVbrtMsEeJmoLhkOwsCQJhiXygxspXb5PMdhp+/J9KkfurLHx8G3sivo84nms7v
9p6mz4zdToIrmwAABKTAorqfNhPPA4etYEXKb9pEbgqglAOs2b/X6VttnlorV6Rv
9qkcKernznYtQqm7fQkeEPPvztEQPAS24VGZOj8156bxejhxkWcLPT3+Df6BVWlM
Hvzgk074TL+RuloP7kcPzJUGgsADRPMFxD/0WKRu2na094rTkG+2+FJIa68BUJd4
OvrbOiAFRLZAXluaBsLN1cCbuyxOsFkeBFCj0A+gf/0kYPdOmUTM2AX+cMHH+WS9
CBYcji90wt8OcdlIurXqnNybVSrciRU1bRI2VsIuJiwFdS+YXVvYYQUllUnwwZMH
qme4co3s82G/urEga7isXbTB63ccm9JrKHsa8anarHx2uBOz5J19po5Dam8QPfb4
PcXqjd/dQgiCWtlP5AKJ24lay+vFOkulgv46s7OIXvIM8QHqLgNfcJRPz8Y8gTGJ
fqfVtrDiWBqwraC8gJZL2C3tF20HSGYv0sIYbZn1D9hiim6MryWQMGrCjCVr9ttS
bYrOp2BEVQ4S1X7BAnMfG77d/zPiDJEozmMLZS0pQ+tckhqO1n6iDjiH3tBnHrV6
V0LsZk+LnGQ6Muw7/VWoVatXKcPNOMpbERGWFThI+Moag/njqpx0KL2Mx2JHOMgC
hEtYW95B6XqwVTs/Q4c+XaBX9lOfJaEEAxzSWui5/+7cqIOOUbSagYpbRJYUUpHl
HyYaVQnboCCSF4DS9q14Zdvt8zEqYXQqDLdZlOehEQy2F8BlUl7L6jQJFIwgj1Dg
bCbZmeobEMgeDrbvLrutypGoSs2hFBbqQxK1mttkAZY3spnpfNyf34WzVypy8JDU
1k44sO6l0SHnt3FCE3b5/+R0MsrurYRtmSyBnfKHDzO+PbxgR0G/1khhkbwcqDPt
zv6BSJDOJOyaCBt9Ews9so2FLXAXJNljwa9Gr44hfA/3lJclhgizT7S0q3009e8z
hugd2JTEGusKIKdQhFDm1dqqHLUYSS7lRSgCSz7RBY98UzDldi3IkKeg28JHGmjX
UAyl4E8sAhToS17kM76HfmJxso6Jpbe7wThgJfSqscy/LEQr9bdoIdcn7DFLU3JR
kpA+jKn+lBZS4PCTdUEkyb6/hKr45X/T4w56MqZ2HihjOWPAYjGZ/6HMgAedX6r9
hbe+w4gg8aNqjubZtMT3KJNtw8MLMZEKqY5pRifiW2xEmNnuUAfvhKkSHrMzJvmc
US/wYPbztSbcKDAmMGZ8inFQW0lqO+bVcy0P+yrsHudzRsn1Ele2z0BvxjZ23glt
AnVekca0RePCX1iN8P+Rz1+4Fl0aENzTg4zLXHQlklcaWy1qmvfndvqNxCo8RjVZ
Kr8yCGmuxHZt+NWU7/1GsJdqsKDhrIcadPNmbBvUzNFTv3Z6CNnYHYUWzg7zoJkh
J/Vx+rc7Cp/h4o5LuRx+eiRQePi2hw3frcAV4xCdwen9eI1epcuBJ4/5ssXEOs3a
cYIap6BdobUkCMmEnbP0j2GeGEM42QeMl7rR0Go8YTvWQoZuFfkbcpV7R5g0a1M7
nf0iZEGNejg+Xy8UwH4mj3/7x4gIBwqPSHDu6u1bbF8tSEYq6xwT05PHFZUk3RZL
p5OHtX+GvpdzgGe24ROSUL3t1RonGg1sjswrLe9qwrjx25OfWbD+0F6ZitYbpptp
1IjvJl4A9M43fgAPmL3SX8f6BHORg6hnSiGXnPWkX3ei3MWlA3+y7O8UvYnoahHC
BFI9aty8g2GveSX3dS8D/tLtrilbaXWDTYxGG5IbijXXwTxsgpqjfRZm5Z4CyoYX
yYtj7rifH3EeaB9r1vZHrY3HFVkAk4z049caOl1cH+0r/756E9CiPXalnNk5Athv
dYoN0V6goGzdtafyL3eWrFDJo7w5xspqP0TZeXqg8y+aCgtNQhoPPNuA6FdIsAGi
FMK//P32Xl+olvfIXwA2J8zvD4dAEbnzrPZdqItVPhpfTITaSJOwvK3DvXnWvAcr
xvGyOCe8B9ecE5SHf7H7sD2E5gQV7vWMVH3VsMd/FLpA9JKJsDMwJggX4AwDwYrw
erjfgXyXBZcmGmEi5fPFC5j7ZBxkyxBPqsJEWjMjkU7akukCgkuayYgsWmEQrl6W
N1zrl7MMHmq834oStmMVAbRuw2dX4dKI6hRVOQmLjBV1cXQfxqitt7ymoXtNvE0b
VPK5MuaCFEIrA0Z5MKdtfZCQ1qXBISmuv5eQCRYXPhoKgUsq76aZMnokJ+lTNucV
l+oUX6qdOI6Da3abQmT6JqgeNn4S+XE2xCK2RFVv5CO7nHqSk1Ooyrvntno4vMBb
fu2MeQX5F2Tu9zyOzWAcgYSn69k96rin/5sp2s8WD0cePQQ1VF0V0Z1ZrzTh50uY
8NE+wPEKpQfZyklmN32T84H/BRB184s32gRVtLh9OXewz7oGKsVIeiHZoS4/7ilA
HZFnigLE+hvWqmlTtQoy8fqLQBE2KyY49eL++xUr67jhSoI9MbypDMyU7UN47GTn
BmCzHig0oycxshYKMSXDZczQbTNBbsLr9H9bHfqnbuhzDHQ5MjgcfGspRVbmGfeA
OrDOJ3VB8tTsNbN97c7DK/5eZRQmTxU3L6mz4AanLggnmAdgsaTP+l/N4YUBO7+K
FSkXHWWv5eyTjA4LCmi5DiiEzdQkNtq+pGSy/BT9+08MXEHXoWbX9oxzDJJOs09B
1EFzvGbOxXKSVqo7RV4DUSfNzI7V15O6Rny5An0OF+y27WwqZg5vazOz/p0hSp2d
tdCqRkabJTlwTSJR92/R8DrXBoM7wrcqd4PBt8nvHCr++E2VxA/ACuTA0yUcYzf8
W7QgsjDoSFwL94UakH0HV5A7fpkgx8higupKsSh995jJ2j7YkI3Rb9Jn0sVzJT1P
2mZIn+jr0jRrIK614rzJrOjwoIRd4jycxDfPg2eDJvLzJ5k+sCGfyMkIQhhwf8Xv
EsVymRv3nlhxN+FL+xr8AsXxhM9IA6fqfp0PMgW9YoWoipioAclFy3TnNhg0Nmsq
WPb5UGd9jiFKnV6ZL2pcbcFyfT2G4/cuh/lM9R4lc/M8zCcHry/HPDDQFnSzDbh+
31ze9gahIzC6igA2TAwQgef8KZ/+TT5aPPmVjDCg335Mqu/w5hjb9NXJe+IlLuLx
IjlRh0jbXtC0LGHAdBHk7l4wxJJ+uRVYgMhVV+G8mhpNKb4mZabC13EdvTSunGYj
dtY+SrufsQIIJMEmICdKLtGQNolhY8LC2vGjiEtALxo3xxSEdrEswwTG+8Nwmrii
83tOFrTa2KMhZ0wPXn0xyk0A2zrKfJ8GTHRbYMOnTyowdjcnDNc65isC6gLcawBF
ZHuFZFYRJa3A9Eqa1dkWpVMpu6a77Xr58j1BnOK9peNrfFJPsol2ZrA22oCZTpV7
wmgSGMuB5Q/cuKgFgz+qtBzSkUX0vle1rUuvYQO30BTnH1GK8K+eJlBcMyfCNQYX
mXpWWwt4Ng+RaPxfGTzuwGXikuV5qP8Rsl1yVlIXc3OvxkWIZ3c66RTrQROwZkMB
m1QxgKx1VZmrQjvAU/n6SP8n/v7pRLX7lcPwMFE16lWAjdeg0sv/6iGs84pSJgMw
wsBH6rMJ2BLl/TRPA7JL47hBsdB787sTWg6Z0lU2/e4fV6oUap/z7F/Rf/pxaho5
SRFqLnOpOisZqS9hjsUjFJqaXmI80vQPATFJsMLUFLGUITf6wPtRSxtdIrPFTMFb
pf/HGQLigAlmOKTOCU0bnmFfw1O4JCTDV4wD6KtHIDhOD/vQ8qrDP8PsCLBLpq2g
n3qFvsvpUw8DauZkHdc9lhUNxSL9IvKLaIizeG5TrD9MHtGcuKGuf6Ze/HoAJhh5
D6YhGNl6BsGa3RY7kBi3aHvXT6GeTPB7rJDgzWZc5Lrg6Ta1liszyHu5KShKX7iB
ZruLKBq2T7ehmLoN/CkA0w3xY3KTQ77L3RZYOXzlNu5oUxLT9wlVvgW10Hojh7Sk
sa4zMEG8UKYYNQCLqmFde75Ts1qFw3oeXi+kUTh8SYg+paeLWuD78EneJAgtP9uC
KqSoa00fpBeJ9Ebfk70ahB8Cg/ZbiOAjKEu7nW+v3zYlU/0WM61WQr22PkYCZQ5G
Rmtdo/TnUXVtwbE+AwmlNwP8Rn0QPuSCqg2y6O6g4gxgw6sKmmen9qfzyvBPwE+X
buGWCqNo8pFkr2a/8c9Xh/nStX2G2PKeP7ZvzKaiBFeLzpgeYSCXgSBfT37JAxWX
rskr7erZiSxtEAZfMKS0oHvHq+DaH1t2NTe2WJ7JE4ske3cp6TqaefOcV85rkq3u
9oX6TyMWBooSQvY8c9jqGipdA1eu1LS2MqyhVC3jF2qXkgfTGpxQc1EwOwn9MCZ0
H5chkX61mcp85XXktNONydwoGLln0n98migBu59bZG6YdPu+EUix5W76Xf7AGvJh
Hw3ykjyWvozmfPXja4DEL7p9ZZi4KIEcqsjmbjILajQyFbe+n4PLfvVgDxAm3fON
C9qF3xY1+EOUls6IXGCV4bSQYPJ+Bn1P427XuUxOqxtWdpZbWcgQrX1XVkL7NFBY
sdd0x5SSU1pW9Lw4id0LHl4EW/YG1CcS6KGVcFLNjxQ231Wf/5v9njWR/hBKYV2o
DknWx7yTNTaL2KW2w98wIjqHz9m92AmVpWjlpb7rjTUSvOd3dISiI6IZYkrgg/0j
zjK1nCSJmfifMtke+aQ2GHMQBg8m3jlISHuwEr0d8xUaAsOSNCZWKWeE+kcfmnXq
Rqm6XBunjJGD44R1jaUZQmasMr+noGxM8LoeYuPBw00BNd69hAx5eUiYAM+bIbTH
dsnRZgop17hacnzLRRU4YcWT2BBpTMSfJx1wHx/V5aF4JsgmyeZVLfvzl/IdcKpz
qU+4NtOVG7pKg6Unt0HSOMMd77O8sw9BxbDYB6a7J/WwKDANHWe8epRvKR7+AKVq
HxXPs48YrJEU4uQVPd58mqnTmkOV+MdUbAYiDN/flQrvSKfgTyCxxjKgnAo3+Im1
yLorksvmu/7B8Cee9POeMGK9DC0zqDbKEux+BHIqTMkdFW6pbYUjOPdAWwGNiRxo
nfzAZBU08CX348DQfwTmJqquFeUyr7C+if0jZorrp+cdMP0nUUDssTy4Xv2jA/KC
V9ixvdaDCc+HLXng6OqnyOA9lKwGRi5UFhzWZW2mSfcAjUQcUyfTxRRaTi8YjOJK
U38emBn4T0iiGAAyoqax720MGEz7FSel7n97yuz6TT9ZIJ0Cu15q5T/iTB8+Ul9x
tP/VrGoIyOKsBf6q4wJEC7AZUfleBzq6BbD43nsnW4ntK6O8KcCJRdf1VqpoouGP
JwIVq4Wbh7WGspDXG2TQQFpCDX/sJs1DFw/ur393NX/nFVTiAE+jk2h/v1ovJB5w
5lNxjWgOhrLsuTq//fsjMvQGcEaQu5YinQi6XvnI++w2EHD3yA5KYFuCfiOcwEfO
zBOLXFH3P8RQwCnyPIuDTufhcXhHgGbjh4Gk/kHTEu/4loOjJVKp6xve6oZYjWCG
mWWCuBbwZfy3fDH9CHnu/8cfqDKc1nSpP+Vo02zWEJD1+/U4lYstXMl1I4XaWhFV
ljgbF8S78dS0WMnES+XRn2BPpi7SQUtR0uGSmuIgrUt0MUJG1aHRxciWRXMv8O5z
7PdLCKBYJoV9ee+5UQANgyYTVt5EFONNM9Gk+XeJpo8yL02IQg3hKOYxYTgnA0vV
3oDkR2w593lAYCQY+zcdJX91IpgASijDgLe9V1OIiJ7uQbRed2Bz6vyJT33saWqO
XgfXcjDLEu2Q3XqSHTweR4dQhCfjXfi3pV1n45VoLm1BojqZ5gtyXYjqVuCvy+qh
aDrriGUC9S9FMCXL7D8NhQ30GgTm44vbb7Qf1X4I4/X7lChWKKCmsKCdIteprDkw
ZAEh3kp93lcLCW/ndqYMiAUArw2IrAM8kvajGlm7aI6zM+5r7KmyxaqoMHwiiTnj
xOUJOEvFHInEQ4NRVvuCLxVLuNZ4ZMjXZX9ZpQKFQJhaUFAgKmwMaAGyQ5TUN3Hs
9sf2D0+8TpoLTaIztwvXhyBRtGI/vdbw32j0eF3c+8+Vj5o7XxRBHw7PFxhYgGXf
nsoaxRCW5MBhG2krblDTOcidHOhnrVFeBZ4Z5blGIc9mslc3TWw0/J/QInBGCwAy
jC0Tc709YvIpTTmfWDJpiRMHPEBhlJ557nTf65/dNRUQTWbTnRtRgrHetJd+zyl+
SV4fn2oH805jWFyLYSU96OLbyldMZHD4qNsNNRKxPnpKife4UFdivTls0aeTStDH
l1iCi4IJCn09MmdfNBCd+uAfFGTYLT3X9IiZ2IMnYQhMeaj1CAsqcs467HTkcIJB
cPG5+rZKfdl4fTMvA68EsJ1LW/tNhKUB7LLjWm0wjD7IhXF7BuMflGR2jXG2PhG7
0+TRXMrq8Tm5DOpxHb8PN2PijcqcbyRdS7PZxipO8qQ34BWDSs3wVgY/nrk4Zh1L
Qkb9J7HuiM3EuiVqNS/bQZgpPRli/EQrfUlqM3i9ZfMT/J/aw9jXt5e0aDlSm8ep
BmyP/2wnQ7yzFnGQbJT4FaW8O/gvhlznh2lWlR2ZRJF/joKHdUIp8pzseVHRjlwK
ltsHw2KmUUp9YLtUUz9Jt2ScNhIAN7JhptT/R+e3F4mHDGm2z2aR7Cr/+sIpdzWJ
MypbJqg9TWDHEbpZ9jxHCIJXIFX3HUU7Dz/mbRb0hlzKYFVnANyN9QUN1faO4NPG
zsiVEom5ieUrVYG4ISDH0BRNAb0TTx3iy6yzF0jRfAcQveRpiTdrQZia9XE+4dMQ
CnUMNCZ/A2iIBFwOoxcfTS/7dSbh1uoy6+2sPHsmaPfphv5n00EcpFXgpxYP2g1V
HWA3p2+aCbcyFvJYynhgZf1Ec9Gkz/nuFlXv6+F5nVVtvNydgi2LSZOTV0WJoS7m
fb59adSMALuYplLkscxHYuKlBmPrKANvfjgoI55ClKMGxguYhol2M3k3+TxbwHCz
vWIOovaUSxCEnfG9/IweKf+gChQdpuiymGqTdYafm6gnTrGpz028W6HFF7c9Mixz
Jy6JAnra7SjiGCKE5YdxemLriM7aiAgdh3u7CbAp9lbeStdpU4PkJd0OCRly6vTK
607UVpY+t/+VL37u9ndrexsvDmE0jQgxdD9Gn3ab1A4ALQsmepP8M4QKz5Xaip/H
iFSKTS26qAEhrOwzNnZ1MGCTUmhOKq/my8V7DA0yV+bSSiJ/o/rIfPiAey/MpTa3
HC5Lb6/oOsCievM7HUJmWdn7h0BeSGxEcDNlR1EMGqjIiOGdfdxWm12dwUwX2Jvz
i7/EUI6nlCWnt7x5VlyDX0H8RvQ9HwHwGJNPDKb9EMmSnFEfOdnocE2Rn5ZlDs3c
rUX4rPBJjxIujKWa7xkcIJxl5gIQszX8toR4ZlyhKFnpYq4P65fao74+d+WEhA5/
606Y0y2VQV8hw8egiLoM1ujzijsiGLEpJKDf7QkWMPE1Djl2VVxTMuT5f1xbLF8k
9lMP1x/qNCEcSKli8OKCsMS5b9f0DHg3WyYzjGCJ8vz979aBaV2UVWi2VSzUZaJ0
bsnrj8VkuHsS8UD4fyCMwG5/40MPyu1Z1jc+Qsy1a3IaJNm+tKvGXapyR3fvxVyk
fdhoiMT4HTpptsCgcsIvldUwsdSoDnIhWPbw+ZvL0qFFe51wHspVCQgXShPTzSt5
mb+0mpydn13ZvYrbxKl34+Y42I8C+WXCNFKa83HEZUEk+B95yc2GM1gNGaS23ROt
vTKr1cUycdMuMP1CKzgCO6RcN6gqVWnfZTQ2EWvS+srd2IRad/WsUbLheVfQy5LM
4T6AT3AIPMEhp2YjhrQ37zeYas8kayX5EytZgdl+u2cYOMF8PXgnTYFK4GBPHGgn
X66cH6EnTa3I9v1r5jtlvbkuNGVZ21+1j6Lu3mAk/5Iah6Pz5sPB3rVfHnUCd1j8
UwMitMQKtTBR5ipDxA2KBCv8hz3ThDlxZhTlUTe9amFDB5sjuBKifrsJGWj1WkVb
/hubhC4oxi2HnvRHO5LesHL5VCVSnWsB2eOhK33wVRbTyoqxvyMaQna607xOJdcY
Hha9Adr6GkLQyRckQs1UGvtBAiW6ptGeHRSI48wqg7pJYW7JgQbPdVsd0W7jWWEb
+BS1Nyr/ViHEA9tZRCkZQmDgHh4s7HMInlaE/Nwrp1ELuiiwmSHC6OTRM1jVklw+
IAUv8bYwozVS1YBo+khGq13g4T1FDnboYhGDyWyFU3mEbv5fx9UmA/u79rEJg4bV
LmFomfGZlt6DlF/fFl3zEZ9FjB6VckxL+Z6aBeQYUdSBVJOCNKP5bfbtklb3clZM
1ISrv3iM7WSQJBWlfQYR9Betv7LuOGfEZxo+2tY8yr69sLB1JKnOC0//b2b+vJa8
rFP6PMGcjbitXQCGCRVsUIOirveGo0WZyl2UstokF/szvqpAp5cRVqjztzwqbsKZ
Sbjx37DvCzFYpKxKM0XUl+yIDR7nlfVu8UaBa/H75dIMzuaHicNC9bhr+TnfRST6
PkUrV4TcxwqFhdP6nwKVxTBZnbOAwMF+BClA6xRk6Fp0Q0nHfEHlUKRGp+a754ez
+YgJ7g8YDcqpIOhlD6+ib1D4F7tOmI60ZXNv69woFR7l/K+oSI6kBjMe7K7Qg0lt
cew+2PUtF6I5dpULOyr+L879f6vnAB+M1VJKvC/hdnCUEfGFOKPnpi52w/5ZI7Q5
rLVlQ1sE9J9frwgmKU6hWsWd5ThcRGp9Jiw9VSZucwwVlMjVAvU59B38ngE9CRrI
zuyv5bZxVXTnX7GlemEePmTHnpG4qPMg5ImU4AzDP5AcJazuq4oCNq3GSSMgWwRb
yOA1MDuVca/c5HokYTKksFhyRotVFARcotpofgXma7BP0KIxIS6+2Vfjf4bCQMy8
NxByDMKhicw++sYY4vwp9Y6Ir7kKPxHsCxsizkEYWrbCTaEYa4ZKdF7f3V7+YV4L
dYovOY3yXL0PIedEF8G1c3qo7L/N/mOzouwNFDKeJ5F4VxM5FxxR/5d8PO7dFePm
foZLCRy3L/oM5SPDBwM+xuR88jvdC18/Td1/Qj+qpaCGUE2PkgsZMXre+kNYlb9q
E/S/6+br4dG61nV1LM3LOH9OimheDsCaYwa5ubMqeEGjJBZzWuQ7ENUZikGCPU0N
y6g6nC7c2MuK+1SHvWXnoO9wVZa+uSd+zOhO1pF/Y0IPEnG65lBz+QudBNGLuSIZ
ERjK1fU8gnRgSOs4t1dFPgr1cfXO1eyPsmdVSrhiWlj/bjhKL9pwbsQeSmoMOlxN
+4WbSNAZytsmwsn+lq8glZhwPYv8IVV5771t9HhfzD7QvrscQvbSNLm0MAjfJ9pA
3plynIMuI4myQqza4vroFeTZyY2D9NXaf7w5SitMu7TKkcuLUyvLmeI5222Nm1kW
IMEFd6vF9RZNruDO7HrX18372T3mVvdVLVR7UuzjAQnnkjS03uhTek0BkbuqNDkn
3GK9qLO73UMwzB6u3ZBhc33FhpOiOobTf0fQZwTlMI9CD5gsm0+JBEC+6fzxADGN
oxNGgLJfHdgaENHfz1jbHt7nin2sN8CcXZnQ8JBD86W05LnQH45f3tZc/bJUFama
d9Bd0XPAJIi0MiTiCvUmrGi1vT7spX6QfLQFKKHzmy8fOJdNrvyvrdWzZWFL7M7Y
JDO9HCI8OAuimVlVGqQiJ4eoMgd9prLuf5JU+eyCXIJGpkO0uZOdv5Nd3+gYHqER
FACtyAhfRY3yQqPAfkZNRC8yNwaVJx1sCKQ9VF4RdIWEzTy0yDQjkR0ECeEv9Adr
QEaa9y780AOi9tygg0oNiF/DQnvf3JMI3PwvZJ8SOQiwagYBiOboKr1SmZpde7nh
tDFBBXGDP1YKJcmMppfZELe8Id98qR+NuXRhqLVeTq/TbArQYGgvr7uRDlfV0Ken
6vTnx5SukffeRLUFQ9gySy6SERUzZK9bPl6jdjcTvyeTEja9SH88gNyfrTcJrgsp
Sj/TzgiDPQ9AtDu84v4KDmhqK8gQxHcm7T2cJdUd+/+hWf+1L9gQmJ9xWygUgiuP
lipBPljGsfxGhwW1lI6S5uXsENWaxNWiwVpYQA71JZUt7WopEauekt4Xe0VslNqA
omeHsGUqJYVw00lnxtxQCZV48Og1VLcqYuTIm/DyJcT2eu9S3IH29TNUrrlGKxzW
mnIzjx8yDG6pSLVGuCvXm05QFWK58FVDeEwkauorkErimMbg5ZfqIohpaS3ZcGxl
wvK0YC5/1Z/OZogPp2L7m6kUdIBoBip7qxJ8Ybq7SrBf6xJXOtA9yuAyjoBMvwu1
+8HuvT3w8B6qos93wqAEBHp4ZXcQzwb6ZIsx5hoNzAvICKEjh+s7E2XqTdWBd+A8
ugxF5VAfrW2mig5AVllBWdS2Bt6EECv4lOL/W4e9j7WfgJ1yqkVy0asJkwymKIo0
xtooZmByYW0hp+2JAfGK5DF0lO9/el/u2P/r2X056WuFacjP7WpjzRxYw3RlVtp9
dXtD2mpvbm0vNzLio3R9sLOlpDtc9c5ZkeXjt+zDccAPqLLoBrgT504rw8zR3VoP
lEonegcK1S5344XzGyu+7C5PzVdELLhgWopWJUOqTNdykJnMgfXndcjpg+gogIrY
J8XwuBT2+VC6ARrFvjfibTlCJ1c871VrPgoQn4bduiDo8rpFEO5hNzqdJJzjKZrt
8acjJPuFdgm1wcpXB6rw0lA2ktXwkBHyaDHt/dpWCTpsHvjwJqvMVi/orhVVVpkA
rEcoiDwoqkDjoIrloC3oyuNlg9Wzfrvn2WCh0i/jJn06+haxGwsPeJv1Rb+e+crE
/i1S6sWcus5AOunbpta52RicK6ZotvX1CWvcSBeO4Ju64zEFNdxjk6lnwrXiRGMN
J5UGf8b7NPambyFVcdowuGEMwTwIMuhEYpNAZHqCXxPpixbY2NBbyR/F/Bc5TvcA
mNOH0bh/BezTBjwINoPJnYgQJ9CFxXdEko+7AOnGo7YpwjgXPL8OPkmuR16UjjNY
Suh1YYGCZ1Ierb6ltXowWMqEQ+Kb20dodTxAkL3t4tDAwLqCAOfZ4jvpvCJTj4Dh
e2lVAOWb/7Gf/oI11ijywz+pEP58Jle2q2LyfvONsLoUy6bM8WQyBRpWZAkxyC/X
ktaukE1c8yBdSLpwmLb+REIQxBUZvGZDNjin7AVTohUNLI0Ao652fwDhZVu9d/Uj
UFo8xX4oROKeMq8WXc1QTxkkZ9KU7FRbYaoWIEVdUl4sbBDETw5xmm0qnoHMTU4P
sJL5hLgRsyqnRHOOLTv08TMVOMsPrFxQtCv4PHRrkMrELupsGuEZWuI4bPxnoKLF
lCzjyB4VQA8Tcdj2UBQP88NbGXNkg3FYh+XnKejT21kquLIU2Dk4wEp6yfjWzQx7
4XaQF1vnHdIgzJh3rFcm0OTjyxa5mxhH6MP2HHofqZImd5lfRaLGhK7cOX00FObx
netli3tpIxrx2jwgui751G5nLlsb2SSTmQe5SSHr0/XGHQEm5/Teun6uicr2j1LB
T9Uplvzosax2sn+I6qu0jDVTHo/su8gNgytFk04T/Ed+qgcGqpY1C07ZbSJdiyA6
Th32IMKAb5Fmr+C4467rqhVSw2oKTmlP6ksxgpTkAl3devmQMZ8UVGUHT0tLwqZO
ZaLJCnkQZEtL4YjevtH7RvDFCpMcnb2Vit6+d+jATtLkNTZER2gQ97ID8uN8ixBL
FVcweeyhnj1Et3av/OMD6Np9jpi45wBRaOUivwvwhZxP/lFhzcIrqSmKemJgFL3n
oxZd9oTdXcSwv26sHTjvHoLu0IEPjbvTZ/7nYxxpTL+4y7bQxGMdh5COtoUYMXvK
RhzNB/Xj+FAfwBY1AWtB+l/6vXvFxdsxjJ5K8dv1uQ3QAsiOPTEIm8sjc5tkKQ30
dvmsJRr6U8v1csj62/mCX4UFANKWmI7iFfmeZSZzOh0LZeCRSqbQeeYZgYsirQ/Y
0ByG9H5R+RgiDLP8JuMcUhb6YeuT4M+ih1znhiUsRnC+Yd5xPuL7u4C1uR54pn16
B/Hg5v8T2EDQsmoPhzBNbFb27H/I5HYo47t7vXOzgppxcgV+jMefUoBH/sQ0WwsC
eoj7eW+nOl72q98kVCf6S43L24OFAruDgQ+H8p2/AfCAIlsqU2n2SbYM4qWumcjY
1sWqXuGJVsA4eDZcP4xAU1H9orQeTCREdScht/mpXARBx0D40WPwO6mYZyR1MXHE
y6/8CUer+U9yYBcvig+wRGsYjiRbs7RVS8PpwyjMEKcEtLTxDqdw/RT9SJ70bHU7
aeWWIykgeaziA3mbjf9F96ci2xWzIFPuBPWKOMAR0NEf8LrsDgPqpIHfDoecWKff
xwG5DaUkgsI1/Ez4yte+jBi8kv9pwjG9ZNuzpEp4MkVQ9+LAW4n33la0fUzx+eep
WiXN04BwMXM+Z/abxjP0Pfy3cBAH27HN/tVdLiK678ZEAmay8Hhlg/NbTStOFmwK
bGHaQPeKjH8lxpVriLzw1uBwf0r9RHAxY+17q2ptF7PudHSkdY1gjjPudTNkAiy+
sTiacfv5nqKFqpyjBkC/wVzSR8hUrjyKbyC75qeHNm/vQ9swo6J6ERKKcNB0uUDs
dfSgxXrDKi8u7CDmQ4XLWo38TxRp39YiS6bDjXv2YQbrByZGgkzBGF3l7yJwpKZM
9Zpd05qrKpuco8PQu+viUDIhvX7aGjV8i76x8tTtSXn90gUAJy8e1bDfEbgI1/yp
T5TBD2xRfWzCs1SJX+iXIGu9htJXa7UJ3Pzewk7frT4wmDXJD/sKkr3liK5ymAGC
r0mLD89jjlYF9x5kcYx1IyJSftYZKkpHjaUAcoeToe7yEnFnaNl8w+DJkrBCKXzE
R7BCkjehDxqM/Fwvmvdw5UjQPtk9Lnc7cgWWyePqQ2AHh1kfQ61fl9TrtyPRbr8V
PfkLM6Szqz8j+DsQw50BVE9ufkLN2lHtoIrxdRAHsbzm8qxtZH+WOTaWfammSZlY
UHyB6KZZHlrO79+VTxtZcKdhYF0nXSIUAEqth5eO9pcJAadlHUZgsLNq4kyE4F5C
V26FPK+pC6/KarQG5Cs09QoOC684ZUiRzv754Lw3d7VwGYwg52VP8xnDhBJhINvY
/x7i743VhQw9d7nxgaF14EXECPRFtDU06wyTViuAsUMdCaAO4S06X/RuC2FoEhoI
wGyn6uEy6R/d7B05DSyn60SbuSjlxRBl66adpeLynK7IF4XE2YPaTrPwbJiLTKBW
srZ0UvkApOGfcYG/JpGydauuCfOHLYgNS8CcqmHuhA75B9mCDscZexKE4PNLqZsa
Am2WGnZzeHwdbJ+tY+srPgBkgbSy8iF/Rrzz4EmFsXosPzwB222XZpqSkjFdtBdC
pTUgMLK4POU6TS57vBKivG/7st6Q3j8StBTvR0QiQpghFEw0jLaqMcfFGLEm+4sM
Z4dTnDnO7pnzb1iKq+R7jECoMnlbg47NYlc3C2C6pFRIERwlvp8NYZ4a/4zt8rnO
MPQLkf078/T6OGJv5iJ5aRFRE4d4Yg193Bnu/NRoGwjS6/DD/KdX+iavxtT7XiJV
uiOjedNffiWJncVO03D7KHIsxl6nN+Wo1dsjhupSYVAbXS6CD/6rrcwW83tI/dON
Y1zFcLKjNQAdkNkYWGTnDZ1K2JGaWoOzufqEAV8W6Zk59yb4kx9TPXskLpG1Def7
5k1LWXbEXOeKVCLxvQLykLtFHMe1WbC5Y3vmyjOHfRUaX2gNL2K0Q1RVdiZ2pjpx
QUw90R26nKcC+ZYGyww3VDd8uyc2cSHNaga4Gnohwos0QxUBFRYdwx4g7uLi/Njl
XcSUEgI10MHcDrUxHr9kjCisqBYx69rCYZ7cYPbZi1oNs5sah5Z4LscJWge6vOHv
RbSWtbqWilLf6pzVzHTDskjTzlhHoLi7ahpMafzIRAoJTFJx6zYXjcoc6ddZ/Q4a
g+BvGhDUql88YotsrDQtzQkB33Jd/WxrPM9+d2CZmui5oS53KKQF0VDyBDXP8bu+
NUni8Qiwr+cVzkpeWI2WGwV2R35sOp7+KGjDwqshBRYxJpGT4LcIGZwbEPdm0bL0
VYVqeuyC6aBNdOTrG9JfPWM7pjgx340JbstXHGkK41NpzAYpRcu5rsI1k0dPwLTK
CW6P8eD/bwpe3tIUkTtRX5/ae3zPa44LhJoEsXdCTyDl6tpSbAWMivIk6nFj7Iqq
jHbvSHFhK75LVfjuWOGBwqhyYJvgzW8VEzoDnyE9hXQpoBRst2u80N49HWOXTRq5
uCeQGdMwHsi2eKzzRl6KsmcQL4pRV3RsdzXHg1INeDkoxhr0YXTFQzBPqB+sWxQi
bwX8m8MJuTucsuFLMPTfe1i84orRFHmjE7cKUJBag3bQo9vKLRohsYYseGd6D+3I
yVmQeXIg1iLUxD8kmdHnQoe38pT8Q8odrypbvcPzPwYm/pPSQKjVjkVlYlPpKFHD
aE8IxKx193dXy13BqBkKu/Rcluy3LDvFlxmDySi5OFaLsdVe9RZbgswnhgLzc3N/
6Qg+lirfVPngWidzdBMeNIbIu11A//vWrarsrNWT8dwYnaial1+jYDPV+2e26ffB
oJLCDA54MpY5z33vHtCZk49qQ2M+SCk+gLDpZaiy3r9pK9rjf/YlrfObp3q3LHQX
42m+7/PkACjPr0LsK3H1MJeto46OR0O63lyXwxIhyD9jjyWoKKnV81JCk7TnZs2i
QFokjOpFuQXXIpIUfwQYtbwDdzgbQPfvb4LxylXvIUegDQwi1yyyJwLta/zhmRsl
HdsS9Gtor0ZavnUU0TPF+Qxe4bKxUlglfCjQIG8cU5CIgHsJG8fbzmkAuQcFtOBD
+0wHkVM8yF3lRQ4/5yXA+jQNWSInXav+bdmG3mmEgmdr6UGiVUwh9ZUexwb3Gvc2
b90eBb++4CH6XquIVoj9bbwA2EkUA6EMiXT7gN4fs58K5C77pFVotYTZhG8QOS6i
CA+UjgpUUxQaZrrbLF1R2vvmm3dqlTKijT3CCa2IKxByNGw4Qnwe3V6+/jpeAfvn
tGoYdh+mKzmfoQze/NOsOtXSHI0jX7JRcizCO1hf6Fxng+4DHf7HJhKNZI5Q1Vh2
asU744GpLdw5W9aDUOmdhA/WVGd9rNPfjV6aM6JQkSS+4AHsmtvWbK+G9SvQyrbV
vVd7+9bdmkleoynOOrz7TpllEPVYPW6bITaKOnQvFYF5kr6aC7WXwTzZtOu/o3KH
VxgW4if7CjfJuqPuyea+Aehi3XoZXSnx9zs8GASjK5MW2C3KdlC29zm+bu3zvB64
Zb/JayQQbx0MowgkGG3KdJfnehxdQ+q0m7jTZt6IKxpFIBVGRLum9Fo51GSa58hd
7OgMjPe0KE9ksorhW8GxKC9nT3VvzgppW6AOC23eCp2P9oEBs5mNj4HptKr817tk
DYeLCW4oI9p+1iTanRKwe5TycRldlnjxsIpdNm+tBMUTQd6nEMQ1j9WCF2X5KbvH
dFrivOz5+w4Wz4qcTpqgjZwiK3TKEKDu5dm7kp40JBKuGweph0LoW9u+mbQMiY4n
4SbBZugRYSmHUwlrILVtsCg+e+wm4nmQeBXwaAQe8Gq6LDXnYFclYzI5jKVtuynY
wgzfY5S60JbPJvfZ34pOh/bwvJm9iw9/LgvqU7ZKIXGcYw5l7zGsGqu/dNW31O4I
46W2jkD9XqFSvk5thJN0C/EbRHa094r/lvjvF/4dUB86oFlTgYOEkUmpwPmeS+ZX
p3TTZx/p1FQrY4vF0/mDGMx4fTsorU9L0NgmEA0pEwJyOKjLV6eN0pRRjLRjdFJ+
ea8GuI3S5f1nPcFH1JLvMp4Z8z5PRcDVUJe/505+ZhyJZCJeQxc+jMW2jyalgU/2
aQjkD8I3IAJyEbycDBjZBE/LSMwMTJKYKmzfLAvrAVAP4FbnxJxXOy/emK+6Gpd5
Ifk6K1EWdIgIb0XDuY0o3mDFDv9+GU5/fB1Etqqq6f49ppjJkVhTKiBN3MSxcP38
HmwqzK6NIdFLiYn7NSP2T38ftZAgy9k2GszM+ohx7rMzhSKI97sFsMtOnN4GX63X
7tkefPKIDC2TBX8afS0TbsGMxfgkCI34ueYY31f2FWm5uPnmHTRijrxG6+TxG0pc
4DjCr0uDsaKFvYdJi+dyg0EXnvsdBJYTpNtSNHkjK88mULQ9jro2SNMicHBQN9dX
fbPVnpoPgYQC26KcNiJ4nZvZTo9n4nPAc6TrwyTe7myiW9IbT8rQ3IUi/A9wUHZO
DY/0RDK4n/wUaGSHCNYNm6qYNMP94bLaIrL6kMVt4kOiP1Jw+mnOccawhSq1yMgX
jypn1nIjoUObv8HUo/xrdZ5qMmRkj7rWkbDt8CgiX1pDTrYfnRgp/1PP2NuNV4OL
MIb/q3Ia8lmdagWVChZSqgfj4UPEMA6AgAGoib0JKTy8yk1WZLfmUCLHNfTgu4hQ
Nqks18ewYBCC9XptbS3AMvgsTROTKMytw6Skk50ari0+KR8clwmzXf4Hh5UZx36j
K1JFZ+MQZyfgZBS3W/U+As2mc2F2UOIEo+1v7yrCkD/MGOQn6VIy5ZRtOzkMdGQV
uc3cMUwgTisuzm8ZP9YCAboXdzhk3ANncz+p4EdQIfqqPOfL38c6Mm/IzWJM4+fj
uV39mSo9yyoWTNbICU4ncEvMq6vVMlTOKTL+GRuHx+5ibkA4PO41GrToCNljpRnz
QInMKMCFiwk87+06YbFxQhe+RE1msYBCEi7eA6u4Rtxi2oBiwdkA4ioxslQIZkx7
2LHitH7CIvcJvvSR0V6f2IJL5m1J6z01/gN5bwqTlDTZ0iXjFser2dot8utdat5w
1hQnICry6ZLtP8swuUN1JPg8eD5J1N+6KI46NQlGS2yWieSvk/6Zrg3D71Fg5YXA
vsKF84ygieFp75lsvbk/f9C5zqWF5Hye505CQUagh5L9SI17MN9xxEMoQFhy+ozz
3mTofH6MwQr8k080V3m3jJv3/zClnzFL6gl7bZifpsTGWVdls5RG7kXwTKU52Nuy
+bQGaKCKs7mmNVBxpwfgAVrcQl+4P2Se5Vsq6ch9wSirrYJBgdFa9Apk4F+pPTrq
UqbW91FUySVXY0E4Bxi5QuzPtMLI/3edA2U5f2l7AfVeoPS2ifQz+G9p8D/XEHEx
9SfaIT5yFvj+cXzB5DLtAtfLWNtRau0fUQu3lEkCIyKz7zXMwWtGbKo5gIjgzAIk
HFYQrY1Jz7law5KYvIlBC0PAZZu28EVd0YE11PT7zTEhhAfc+ybP/54pMUHQcomC
mwAKUxkyaXeaSzeMB/5yR3BzuISNJoat/zDWBUqdzrxfAFeAWatAmUiUKaIymCoA
cKt8r+pte7iL1xVV7ZkpJDXLPqP4jAW6F9/oDIqfdXPf8dq8JdaKGSSBk0hhvlLv
9UXrdiP6VjSr4EIWiDQxEU0BzbHgeZtBIym+xQnuSd+G9pkWlEcYnA70TnfdPhb7
W1Es9QohsVE5YddfMfG5+1419R1cvWNIeO6v6dAJSd4yW67fTLkvmjmTbWqBIBie
Rf4irvjDpYg2kwj9ij/ldvdWNR/n4oTMkt7I/iKzqT7ExCwm7Be5Oho5Z2o/S2qO
srCdhnluoQrJ5tWbB6RMo9AgBfMEjm6gRqa4IbYI+wXON2Ww7HdMIneTErK52M3r
WVb6fCpMbLNVfed7wo+pvWEXRsK7DD3wWAyGKuP13CDYABGske+OOulCN1+MOC3L
wSBDT4mphYBklcBiw/cjzSmp/LHVyBDnhX9tCMoi6VmE+G9CV1esrH8xyqMxerPD
I5wwKYpMICGxMeFehGr2ZkMFKNK5aN9qKSyABHuiglfoXmwzxLoa+h5rBCZVUFzf
Zn/CKpn+yXwYYh312Dt9tJQ603ZrO2AIdFPUiC4wCmIIVBEwjoFqNxSDLIy63jpg
zBX7JficYX6K62HYjl4oQeGUZ/h//Kn9UtVKeXRMAIU+cD5Bspu+suLtgJFfRBJg
l2HRWT74NJAalg8MDFi8hGWRictA8fUTKASNWkdRIZIXvehf/ur5ZIS8xQVtBDP8
LwR/scD/OE+faAPMRz24wGdCAgzhcxq98ztb6rnNRbajLm9N1jgurJmjowZRHfOV
1nGEYPXo+6eQVjpP2NrpWByKuTZAElfwSIjt99cUDny4T+qPwbwpYY1huqrjmyLe
2OfxQU1/lOlEQ1jnMY5Pfc12E0rZ/niFpDSNAxsQD9mSTwBqRKJ5wuKtz3F+Ix+E
cp3cOd5fIwWIg1lFr9HYPeY2BX10nun5l6lSveLA8ruJ/oo0cbH07bCIccJzRnA8
wtuftVxxFG6qwgTsn5BYmQ78wS1u/qx8m2QL2VRdSfu9ozFmxxBVLaeiwTasDk5H
dyvTphTppxzEKINGYzRpfcRL8gVdWh3WwlxBv306f7ugKcJDzOue/IZf+OVSM95d
TSOpq2f03NZfbAoSNjQzgovKhYs4K1b+W5RRiYOxKBPa1sRfSachywfzIR9PYYZu
4koh/xPU17XcxYIAPBmL8VkpoUAVLCYpD8pIe2pue03upO+jwYZnxyl30khoZA25
pGD8kebNT8lUU2FNVSAmjJhC4Tt2bkI3+tpXC06307WZKuDwCiYGeHyA/iB654uu
88nPnMk4j5Y2ZidK+BcPWC5V0oJeZsON0qCWC8JlW8ujzV8cKkMVsjCeac1rhoaK
HHS+TWsh2cEMOJdPdm3SOc8MRtM9iQRMwQEw0VEHQuB8z9AdraIQoAsbI0ibaRyW
BS53ZcM4E2C3FICFmY0x1ws7/gytkJUy1VcJRM5zQp91A6UKvHMX8rpO38Sd3pCr
Dj2RTduQr+otCS3b60arpIVjOlml1DZcvVNbNcBUS8r+X0k6yjGMi+6Y4hJMuLLN
sj0EaixqKoz5PjppV5NrZmg6QH35jVWd/XBtG44KnCg4sXcilno+0m+Efu6TjLYk
xk5YEQvLVNzAWu6+8aspn4Z8V2IDLcDCQEvlPV+0QSMh3OCfCBjATKkUImk079y5
qDncOu0B+dGwOHDiJ5BpASY9J3mUZ65FWp2uUs+9CNsO75VokkE6buNcN7Ofi9kL
9ILY9FL3jffhBn7cd3mKOlGFNBqdUqJRxrW/mhSU/UvzLaFFTackC7MiDFa5FOa7
PCzpe6+3b43csuGE7+39w/CedZ43QW/6ryP2D30ijY2HZdI1Q4LD64mCAWfEijeY
BCpeW1U+gbn6rgOXGAluiaoQ98ni6mU7wA9MuZUSbs+p1cU6L1bmn0amLF6I+XNe
ifjU6EcW1P+OlbESS8sacQemVtgnjcYlish5/nbtVmuWk5WXmuW9/I0lg4gXQZEg
vXfhkVMvMZ7XYTvDbvbzhAglmb8Klaote5D3Zn01pFY6qXMH4FOrSUAFPDc+bbqj
dQhg8oWmvUuRG5CD9cV3loV+YBAni7b3caDAr9IqkVPEFSKwIYSDPePfgAsoK+RV
Z48oZm/LxZPtTlTaj3BkPK+5Wwe1Eb1Sn8ERxY27e0tVtU7t29aKuaRjQkrCbC5G
mu6WS0z7PA/J33WMGWI1VFxGWx8qeEJtWJ7cVDabut82hqJLRyztohgsIKMJUbwG
pxi/lowFe14BguolJSWs0IIRbD5BswqL35H62B5J6V1aaxLFmi6krOxmfr9lDOik
E3bIVgR/spGAabqG7yIy4YM3nkqDK7erY5GdInFZdv5c3Zw2GaFihsanV5XM9Lf1
wX/OWEBIykOm32hXCdDgBV6N2/iCTVbFpDFIXHSYH3iSzIwLwVEBkXuZOnCAggnA
jYJR6+mJjuoj/+khZV4urC9WTL3kBq+X5K55YQgZwaSGQw5cyRNIPVZAMyqCF3uH
9Zmm55kyCFAq63cuikcxU1YIBg4rDYu4NuqRM6DVSMzVT++4cR11Qks5rIpXUl4F
mRydZMDsvQxzscaB3cf0SPWscXKkypymATC/FWhK4VNEQM/WsO80UuBDNUhQXLxu
FCUP4wKGpxsgLruX6A697E9RZCSDICd8ms27DWKfGSJ5ebqqNoFu1sareFA6E9u9
KlsXKUs4TXjoa5rx791cj6wNSuZACQMtmpiYce78tdxv8n3qLg7gX4MuoSOZp8yv
clxkrBKXUGICzF0E75prRh3t/JFsLimFXAo3RyniN0+RGvi5lGlnKopGQRuJZpOy
jOCPyvGm9N0CEDV1Ul0vZVfqiW4znFz7xaFHtM33h3C8NncRCHc3weOCCnnfcT93
oWBPVJbGw4qWZrKs76k8aLKqN1O24JrLfggcCiOoEwDKyY6PmENGCewofieC7fkp
twxd+AHk46EZq4HuO/wkTVSK1DQ789kT/203tf5o6l7jWfyTZXaw8ZMpuJmqCtN0
0r5gn5KMvh9hOYOa2f2QxZIH3884yoxtAX3MDndI2HKWp4hVYeXxps9E4bOjzkzY
Q5FCVXkg7c3umEWMA9KMwkjXMkJ0CK3opMU1BodYhjFuggsD6XcQvH7yX/wXXOsy
ZcQBfU3sNc99tO84qjUAwTxhCreHFwnlFVsIZSmo6dMRHVbseC1H3/1vaBE2PuSe
Dt0smYHevlho5lIxfRV39rF8FnThVvom3kdRYHXSadDzcn0DQNmJrZMjRKpVWdj1
/Zr4WThB+UtaGZgGIYuYCMIVtOy/2/0A2PTQ7H8n4/5QqxZIwnrZO6BI7FusiP9m
GloZCGt/Rz8mz9pC5n2W+pMDpk8Z94qpavQmnKdMIIdVcTUF3sfTbQTGmxZ3VN6I
ANNVn+PNTFrJiko/FoFqVe9bR95v/5FkNj67E7y4Tsvnp/yCjvoHszEYeYY20wYz
EzbGbioUFsN9dle+uT2iIHtebQwGw470nnBEWITi4blQuMlKpAMaSkSpGwaZH+g6
JTobPgppP6W1cdJw0e8ElsRljIBRNm93SkxmY8ZhsMHQNyvRFXdB99Agqwe/zObf
2ZyeFkucerm1WNK1aQjc6r4TifyTBroepx38zGxNqRQRWFrreKjE5fgPIKLy4O0q
nqyXEerm4d2ueZhZH6dTinXrDrfTszC053KM2UapVwMUp4mt+olPTA6vVuCFf8NA
ScGdGwjRWc9i6lLvejzYw7SS14mGbiBnxU4xLQN/1jJjpj5gTRVhDxnoNcTD505E
IfDVFT1sbymGWrNI+mxg6a+uaZn4XQ5Y3fBOxIpVgMFd/DiDlGFdAalGWieHiedg
QF9tlUnhgSvlxnACnusqQDadmG51ISHk4+3hJo9KZesdcuRK8tMG+psMDRb/ESda
XPJm84kZVqDHmo/05QvZZozPrXgFfhlAe02OjR91NhKOWMYeOvQySpxOS+/Ku57J
g31qtTi3LGSXz0YaT0THn8AlSW+CNbTgMNU6L8rhNYj7RycjxMiLe/h13nf+BsNl
kd+MardSXA7ftmYoIiCnr0v35w9jUQwA+vCGVrYtzyEs2q5ZryZgdfuUYR7T3VYS
SmyCf0RxQuS6JPvxH+WO4GZsgHXsrcixVIvjoduzwGxszXJSSExH6+Y5PIT0On6U
wcsWz9zkmunpF493olZuONqIHkq49BGlC8lreTQsWdatEuu0clb/XUeMWzpyRrng
vZOXfSl69Oc/0MTEkS7fOxHUYrntlsBL+rcS4etqwZqRSgGviiqeLrwWYpXfu/Gn
+edIdFOABxW0RglihkbgCN45PAfsuzds6altxeI78VZ7vK8ksjoY/m3zzD5ZpjoR
lgU4CHy7adR/bED8Q6U3+RMY6wSNRQ4DD4oYGDIElLmcj0oGnhlPS2kasQY4hTHv
TTicgE8r29RNam33QXUhUBmutwf5NceAERd/3KEVJP8cqZiBvbytqCwev5/MrANS
6N86hHvRfSuKR1tFhF0U5a2kxNqFjkRUfPw9GY/ArFJp+ln8mVtFC5le8bml7eOf
SXocWrG28ScV5dujyCQJkFhpjm0nrRUGHW4/urGZVTwAFEdngs6fPaojqudhgXOh
sWWLG6tbFE+OD9doxGZrxTss4ozvWYJMWPNUnAQGOuJCD63VJtaZkHS+PPlylW6d
5C6FSLlHwPk1ZWRAXP+SjPgR2WGQxnJexWhy5xalejToBD5EWctFD8R5Jx8KmVuO
ETO2v2BWpio6sdMsDFC2oiySJe1QDZbRrcNyuhzG8ntkbUBK51IFYb2Mrgu8tf0K
Gty8kLtWG11wLGglMX9Vq9KMvBzLVwp3xxPaJBUcH/RW0M2XbpCMg77Nh1x33OQQ
PhwKrVKjudvIpk08BqkH3jpSDFg6cp3agXltynSV+Jz7NhnTo3+6HMbKUM9JlaSQ
zCN+aqx0HaE7tRCRJ261pXf44+RSenrBIT2dMzbgdm187sNgr3tTkGwmTekjclik
f8Ou2eegTviFIvXA2oMcW+pnVpzovkNX9imQ+ror7q/myB6A53DHjjQiEtF8gQws
A4sSNVp8YFCe2YHu75XxujJaL/Ssc50/BcBpmhbTmHfOk1tT5ixY0NWfTp1DfIX7
EYsjQUqagsefFpZicvK4G758n4AjHnaf/33Xrrkr251uTArwCC5FDBCPHeAoavnZ
V1yMl5p6n4mkdk/AtBYQr3FNv6zKAKJsk3OFuq4nDQqyaHjTom2iUAsE5xNwW4az
2UAp2thGqiOJPL25mUL9ZXAopb/zVOqLPUmYwXxxi6vXYMu+V9+fFlqSN2lvL3Ke
/xaRrdvDeMoGntHLk2c6a4eT5xL72qpPYy35BkJwdySJgyDnwKHb5wGBPnEX1gUk
qvZ34X1wALBqstSpyKhTnQZs/aDrHRqdZD3J44lKyLRjoKmKjlDdFfbkYsY9IatM
YCJNacLkCDEcpmdRhapf/w4mFupovqyXWfiV9JKrRKVUI0NeMgOKouEjSEwmbUft
tNXVWAp6pXnejBMPEj0pCZrwRU7yw8wy9MDtfu49eioJoFkxaE8ACL2K8q8/cZVE
tAur/8BNpZtKjlX1T7prq2A36KGIGjaRt6Y6/OnYiPttbJCOePi+IO47CWw9t884
bFAwZXeKsuItyGQXeE9Up6FrdPL+pbAcc56yCb1PQl5tr5u+/Wnmd3YMMbQjXs6Y
B6omM9a7ZBE7qDDifYBlD4vyJD8QUT6jFDTOtEbWaIZRMQ6pAUTdW85TXfo4/KSh
21fB8XXptYuHCO5fcorNTZ3I0R504zkT0+TsfGIkqDUQpWJYl/n7Lt3Wur97yFgW
XaUOG26CB026noMqgU49i9JAWVENp9BKeJO1FRUXrFxiU6tKjcDh6HDaNG0sMnqW
/YqCpZdPe5wa/CtDQptQVR+3VHX//tz9pRUNULlfK7xn+K2OuFniYkxtcfy3OUcy
0+Dl85O2/qIN4UTIkr8hpUDyvGeMyW5zgDGkGLCLC7qrqo1eNn+odz8Pf5UcwHGD
4yJIPQWwiJfqHUEHpfQshJIF24lKPt9kFUq4M5LwTlsaDW6VPTf7wx70q/MT8v9/
DuQdvlqNdqVz7TVno6MpBSiF7byRk/ijtk0yZgG+sa7SxFp0yG6Rxg9YFkng8fTD
QqlwUGSl9kK02sMVUkkgc3PRzQH5ULZgic9XOm6wRAfFISjUX/PVsleF8kd81SW3
1W0QCbbQpWyRlHcujCR/vMuim/jrGZMcSII9vcJAHnKeNL7Sp6T5Rw07vu4tHWbt
lIj5TR22OfgQ94LiBfxwiRC8JZwUa/XEeonEvXZUVaewYn/yV7UXhciyrX2jhszc
mPNd6FUHFZwTq47O8WNwIOwT8gAT0qOxza8BKW74LgHrpmxA+VZS/sAir9wLCKoQ
mpjPlWjr1Eb97+QqNI6X40C8/rAtU/x+zaSjgWd0W0xyKClNHEFxN7Xk3bPkvlPs
/XZMaGESLWT4AxkGq1JBp6FERsVsIo4CYKgvYTIQP3jyNbCSx5uzlJnLO6wCwevk
DU7gVZkJm87k8V0RRVX14HtyiTnXw9tT3dtQsWFdEhw=
`pragma protect end_protected
