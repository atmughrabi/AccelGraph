// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mIEBgxBsKADaoOZaDp1JuwZZ+BJhXZEKyGIWl2we1e3Q/ZOL+CI7CDbuBs2zPOac
F98+QgcENXpAMnS6acV9IVq5tP3Tl3cBgSsd1SVn7RGZ2RqcSmGwqyVm+3Mh1lok
ASIMrMABQXre3HF4L/AKzROKSQuK9TDYRawGGQqMkiw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 49968)
JPVPVrlZ+SRUDoWBQsn607nm0ECI8JkupAQRNXrAj/2Bg5jes0/Q+Sa1fTQReJ3/
YA/ox0BlXxl3Cl2mKfvZ3/RmPrqhnyU5OhOgsF/1vM3ZPm9/OGuZSJVxmlFckMbN
j7Qxa2RSxX6txKPBEDcsjNoOhKmj2YnVDyYIITtcwoH3Y+Lne5wKmQyHU+bwsrUw
nsjlrjckURXTtcWnEZr6jt0F9ulV1bvLT1RP2jSSj9pxeEf1q3xkNLeASntKdEKc
ZsJqbjuthWrPX9TAh+b9xbt0rOiwmNnH6l1Di45rZW0361Ign+Q+D8VfpKTBC2mP
U+2xisHTR5FdJf0G1cPEQGan5KcAc9c2LcbYRcW7Weip7ifnDtknhYtFJTa8P5cS
KGsmqmG3Qr1L6wMgWYO/r7cRtwLW7Bc9JAIyN5Eitt4f46mZfo743zGhMk4E2IPN
EP9lPbZMlTJJUNJhMQHYmCq9FpD4QbI7jhZn/veIB2KqkMMCNDbOCYTWgLWyBUAv
eBIyZyV72x7UXX4uCZcpm5Gxe6OLOQolW710TfqHL1UuwVR5OXIXZirxieBow1Kg
kFoyHAGPXVPzO3TvPufRnZJqi8i7N1eH6XEs6rwYFiSv3MCQAE9rELo9M9KT74VI
vRN32vXXT6UpK3sOcFZ/kt+py8IGDQIyG1CsoPQAauypYMojcreX+cZW7+ensNUW
TtM3WvpDe9NuqbOex1ZdE+Js9XS5jwDT433Y7675rjyDhfbJSSjLqA8HqVEMiV29
D+2zMzmmIpjli1nE8iYWT4Yz0mrdTAVXqP1GHumqiPvGLsyG9K4Gw1akXuAxcoGq
Snq3XxtNCL4Z00R88MwrRdDo3npZQkjWKnRdE8zZ2rVmi9oWMglCQAlWG0W3W+jS
DTGzF9/EQX6nhV34D+4BGTJj9Qo5pBw6bTsV8qVpoMLeoVuRYWMPNUBT5N/ddMVv
HgBfJAEqBVYle8pk/qGaInI9ybY4LU+UEtUa1i0ZXGVIgjkoSF0IbRTxge/rW/TZ
DYuPmh1nyII0Hyg72+AO97/PPIvdmGp3s1J9RZA5JdHDEqP0wKaZrBVX/OGhKKR0
hwe0YSo+uQ9EgOLwkv/cxqwW9cp4DV8lLnuZCu40S3nTMaLsOWAL+rjOkFWSmK4R
uiFE57bb63qUfzihdD6AVYl0PYCJbfevf4bBL0eOna6nayaW4rRJA4PcS/BZOJ1F
ImQ1Xh5Tb8ynQtMRHhWi1R2gOcnSCELE8x3jhvA73bFbowRr1kjkOzDLaoThTZEj
KGHMGMaFSpRCoHyNI/pIJyqw8gdsng1iShLlVMQRbRIcZSANLCLFmEorgDDFpZYq
apH70mpZHIJ1l0SymHAserM5VEc9EGjErgT/xIv6xg5aIy7JpMnuk3lQiiySH2g2
AXjlZuGWyXl5OHKtuLBUeFZiBAxywdUy+ZXBko1GZ5/FLf/oa3k3I8Ro8tBOazue
cfQGu88RfVmZbbB4NxJZa76LgHzhhcD0n41S55IpQcUcB3zemCtMRHqspj72VYq+
HGqAGqhFSy56lpB1ZA/cE4uC4cWyZwE1Tjxo5IQeGAJ27Zt73V7hmpONR63kH6Kx
YELASHXI4Jw17zKiuXyXdf1SQM3oJvDPYPgEnFVns+Vi5mgjX2z1bK/5JBtBGz+G
K+3TKPmpYw1ZoKh/cDkUoD3eVu4VUutVTI5d8Bsu9XceroQJlzEhl8+Ub/uQxgI7
8P9UDEPV6FzgBOb+JXJjqT6WjBX3Bb34O/Io6Bz8koG6fKT1GkN2g1Te0dUdjnx+
nhZ6NcbPm8k0qDgTxGAeycsuKWzyMKSzM01h+XNs4OvuK72Lk5E5Zx2pkOxI3E9s
yNB+o92h7yaNvPFeOFF6Off0sIj1ahhv0SJhZntBDQtOT3tFv6QkR9Ru/rx7G1vN
Bt+1TxsRBOLoUwkZfVNrUwz/U2FZWPBCW3U001mW2z6mx3RiB+MpjUWWDsWsOPiJ
O0zlr3hm38x94hpOSa0gL/+1DkYE7GXz8phtfQPEKn2iRUlCcAhr/isjCji3lTYU
/gt0jUY4YWyQ6UnO+8An4uTcrM3lgAbkYxD1LOA83Kh51uapUojMZnlpUs5Qft5q
iiyQK8QPdNaU2f5TYrlo0SEoqlyk9QfiCvYKb4AWl9uwbPWUfbFnAiQn5BydD40j
8pBeQHMMgv4UmtIKZ9oLnHC4FPquVSRMyRAqY7C7fTglTyFc7fJVVJJCZmzeQ7QM
IvrfWPriMm2osQqhBf3zLhGTB9gyj2QInnrgP2nywpcIUUYRNPTqE8QyesFGhEQt
cP8MACd4HwMAe2I24uLPpjJ+5IQXqlKLslDEyPXu6IYKQd4ePID66OPDAAeoWSfw
Kk5amJ9rcyt2cnqA3aLqi9EqgGafBxoxNYh3MGFAJ5tr6TU4AyNnBVZBzv4NrA6z
5vI39I1dUhEvJ6KkMD8Ds3qSNSzLMRoohebj/G7uNAZCmer79IrY/Bi7qE1UHkzH
AKqjcx1pfIGqP9N4XFj1fNHlesq+ax14tMfCyxU63fNZ/57B0n0nmPP0Ovu58D8Y
errT+qJvoYHR1j4s7onV2A+zDPip3M4G0Q4nn9E1MbeUpQ4uDhgQ+aXX+Pkn1wxX
Qi+NfShyNp4D3Lm31/pt1DS7fg3La68HR5fbalqkyEZJH3u4ojB4DeTs5S2n0tQ+
NtTEAUctFQR3T9m2yNle7QnUE2ia26RKYspxiik776tNW5BN6k0LUuAaFDLUBYE/
MIHIARlTAFdpNKr8HdMVd2VBZvVWe/KaMNT5Lp578PRhbewbAXwYMLfFv83LkutQ
zPHj6r+re9T7f0sviZ1mDzBgm41qIO4GlIt7VxgziXFd2FtSgP17eS7P9xVexKOG
g4A4ocuTDnYn6r5e4c14WfmGGiJEZ198quqtNQxnYYVAvRA4NfQw56vHSGLK3Vw8
R8yprfwNEPXmyKCR1DyTav7NOHscQULgt2R6hoaQAdyc0yJsjznuhzDetBn0YiQy
JRf7J6NqllCs8Rvjd+QpECemKL13d1sRhwfqWigEvd2SEeu875UdOwB1paZIHlcZ
rin/j6GmDZHb+IxhlWftIrOyoSabhsPqpix1sG21ieyOSJhSWU7XONOISN2uyRt0
yt4hFJNKUU9FrDoVv60fUnQ466Eb259d5kem/0/Iw80Ofw89hGFfWTNovPrLnZ1M
24Cn3Cj4q8QugyESDm2/cVJmy64rMMapAc09HmuzoklmrO91J6ZcUnFeziV+rG+3
vNzfsCj4Z0AmzTWhwt5AqsVtgFw9GAcCNacQn/LvJZxYZnw5WUXhOoqVZp8pAt8U
oSOzUSZGOi4cdk0kxdi0le4+Yw0i2e0E/VB4NHLoxDc4RMeXT+IZ7X2ta2LCcUPl
EqacH57h24pWxZB2gG9D4IotI+3SmUoGWXHmhlX4haRnTcGQIUAUh2+XXIt8eF6Q
/2g3/mw7r8wLk8fdkxQ4L2LabA6ZfVgHIjDZl8XKjl8Q4vR7HqRPPmD5Pn8+bu6h
dcdVW28vgd6OIU6ohC5QFpHbkeJ2LynZdcmS3wGGFgCf6440kiNlABfbSa1JDzYK
I0b1BN9q7KzqbDr6gLPPsVJGH4xKAan/PJ9hyjntp/MIWJWP39WzbKIP0piHxbSH
SVLVXAIX18imVwH9KUJ3QzTUM8eSFiebIfueEFsB2PQozUp3FdL4m1zpNkZ8Gzeq
kDU/ON0RdNZFxWEx6Gq4WSzD95Ts/spLLU8VZIZfHpOJnNXFZEtWTZIQ7+67p5PL
3CTkRetAkCS1CecRyhId0i2UJSb+0a2EDtF3x5lthpUHVaxAbERMkQQD8KWSJdk8
luG7eBqu3zPn107QQHg9ZPDKxuiUgI7WVR+lQEFay6YIij9jt2JSAcZM3YnPdgcb
BqZ2X5tmZWC5r3qbS4GQJwDSd34ABb7I62wWwOhC2eijr2+4gDHmTFwoDj4ekVoq
k/d/PhA7RdB3JNHspBrmu6g60MwJjagdBebdWDgBJGgHMmJ8UcSznQny4j2vfTgn
tO833QK3EkFfawG92AIStOs8gCc8G/9UZRBNv6mpKRTrU6E7XwcLwwUVx+YrPY5h
pWC3vz85I73O69e3+Lh16eQO5mex5QJS5+X9Pwfexh4XDSTRekBqI0Mr0fSyRnPH
9ZyjKgX2uX/S96OblV+mD+EIvUL6MwYGoT0r/DUb6sLAlfIY4xesdrZ6eT1/I3Yo
+SbjQ6vyR653d4SM/SAfw5psIAQg632tnkzmaVlsoYnN+qVZHfZ4dQO4mSODrBMw
M1rJeWgi2Sx2myTGtOoU9kc0eNDz/B32HICuZ8zfda8cpEVRUdtVb+1bGvplJtTj
rLiZcRgwfq2KwHNmlN4Z/N6SBSwShi0xAwhfggY29ck+PKw5Cmqt5GTe2foubk5b
Fp1r/IlrVS3z152MBSEkCkAUFupG3P828IBXwl7G4ESk4mOgYvPWsoquK+Zalj7R
XMmXvzuHHPkLvOgnlFWps/vpKDznYkRNeJt5kx1/BgSc8YYk8F+md9atrgQZ0QFi
2XiKcSUQxr9hDiMrfTInq3wEbVSu/d5FMWGyQ+rBZMY0rmAip2xuhQ1oj2juBSMO
t5Di/OAjkZURjN96iHQg31zLXbVYBrTr4KlY32e4Oy2HfJEhph3klGOQ0Gh4aZBM
3ewrEHlmW2/gu2Rykw/6z/0obfh6jBYNKg91LWCh2PTgsNfHiGljZOAk2j4wvX6G
gy4KLkoW137AmN9NG2PcrzTdWiV4khklhb8T+hYrcazAnlCYRnASrP8h3x5Dzsc1
9IsCaZAoRPkkBq59NBHV6Y9t+DyHNjjcENpCdk0Hk3lVGRr2XMCeZC26G4A87We7
lJ40CfSeJW1CgTYRxhhG//bYTBx5tNaNvW39NfhnDfKoemIrJFGjuDj3ePUShl4X
9yoJgxngf+H0BStcUb0fm4PLj+JuP5kDVT+fwkZdO87daC+UHKsFmwO06+qgU6zg
YAqYrW++BzZxjoIIeulQ56H0+7J1OadKOuNHlN6LB9X7BNCjhESweSU2+49qGMJM
Fss6TRjlxmRlmZDVLgKxkFqZYT9DNA4Be3u6EC41fbtzSieEBwaXIdrpmBIIPDqT
oLDAbMNo908ekinVawvw6iB38m39S17O5uQhMKb2DinDoslzOK8ldEaLkMe3Y5YY
AbIrIfhnX3LdLKSLG71ZsnK8s0btBFblMvTPEIKyBAn7N95dFGwdJU2BPYfrO1WD
e43MlWenhrnfi2IPg1TIHgDfiAc7jYpOTAeXNx6NGW8aRuE9Tnb+53CUrtuighz+
WeJijkvmT1V0Bsh/vZSi2DSA4DVexyrLIca6HYDsrubx6J/BMUtUmDnq5RSLwdxR
yv776uXMdJojPOwjhFNTjdAiUmMrmveKkSW38PhmogKuRKLzuJ1R7xVDZI0CAHJR
BSKMCTUx4XtbwuzjIQzJPdilHl645hvq11OaJmhYnWycSX39IEScKBSqWpbtB2OK
SQbruIZQGhNDXKkZYc3Y+F+2XTxU/1tY5nQS+RfFri7pI1gBRLzjNzcMgEQVfPSw
eQ5Ko1PLTlqa7kMkJ8pAcndRXKMfQx0HtDwvw9tUChktgxFal0yHEAO/9sJ91fAO
ZWtdU4SUVNj/S89Jcspyp6fMWxUDxN1mBQhT9JiP5ZuQFmk4JViwObFQ5vMZslXN
5c9bH0k+lt0HEJ7MsVP7uS3pHiCMLcSJK56cDH7us01ZZit2hBGeFRuwRWfq+wYI
QxWZi9s0H11YwtGpma2ZTTRBa/mIhP/6kw7N1gBnfm2ToIuoywb+3Ov4mFYS7yDx
xQQ53wDFE3wpzEnxkaCC+1O06tlVkDtVZlA6GFfBMdBDvPizk94q7HklNwaslmx3
dmnsi7WMn2NUD41EGayj4Dn2ufOc+Tdud4AtT3s5aJKxgQ0cGgBDIiPF3QcAQXxk
KC72VArDSqwCMVcLwkjxkHvc6gJc5vGkTsZIugt4PQMjSvLuu1tqnjHCD4g/GQNJ
YYMpym9RTRaAJ87BaFHz8s1cqZGXBM1+12xrMGqsxPvfAHHx3KNs4dBtECTkL8Sa
1KZSDvMn+Do8vjZcpw3SfY6/XvSdr7X47N4oDSno374tbmo0t1xgfoZt8jv1OA7m
9T+YI1omETWTSe8HLjDxuQ/oAMe8n68xQ8YwWd0iCqahE3tZVdFhK84cDIUEqxrr
pXsWAnL4kduNE4k8eRKHIlnOPyYuhipJ0/eS8Pj7kiGMn1eH1FLZ+gMqEToXlQiU
KKDnb5okVsw3gv6Am6wtUvB1dCubeMwc01YTEuodvorHARAfIv9h6KMUmTbOuGwp
cbjh1dI20bw/iej5cK4EyMVH6skbzmT8bWHI024b/Gct4QwyPTvbTscl8qGh/oLW
ZvoF/MwdUC6Rpjati36Fdaig27l1uk4esGTcb2vpUCpy7VnfI+tnkZEkBIG501A8
7PTdxbz1x2uQlyeskl1C4TuuPk3fpmL4IHDVehHL8vKdQ63avTt1dEXkG1LEqnLZ
iiU5TLvChzUplttW/mP+a/gzEPUp5ROHiU/25dNH8aE9pDfisy70ThyEkLaaQ7Ag
Ngr1Lk/YjBqCa+vnhupiujpzZQk0Q6hXw+PO7d9d1T6W0tQe/zMHlEQGGqvzqeyB
uW1u3IdVHrX50lirGvpUxx2mXIeamrE4adGKUCXyRvJ7QBtQwObiw6u9hirIsLIV
fmUL0f8H9ew7iv7PaP5nIf56gvPa5K5YUlnqmFh2Uxym0yAt0clhKEeRR6VlFJSJ
k8SS2oF4TmqsSsIs44wyAOKF0+AJ2NVu8nXB1fbQjusMZ44F3PqyvlR8i+ojVZj7
x/bg/BmKzjt3SK984GlEcvp/41LKmTdsTnVmcXEJJenLe5C4qxt0PNAs5PZgfM+A
O9bR9MjNpTU1P82dbWnZ3gHHB5APkMuy/SQOcTXVSLHfpUmhHHb6uhi7JiCaNN9G
WEzRalXw2/WMFEQAUyIFYAJsKhRidhiekAj6vCKHgoLENwce2VbFrnT9P12+wQPz
SAB12O0dkbWmrV2bMI5LilQtEfoPQ5HVm3X11/cE3ulFZtNoNTG/DcgDz1BXa2Ol
FC++2yfWrJkZSMlXeMOPmwBuQHdNvmasDELU5U6BQpaoamaLlNviEkKYasOB8jf5
4bxUgJFYkGWEfofx87t7o6+Fz3hpJrraqy5IRXf8loeUV4ZjheDy4qCL7xZUj/IZ
yAaNAEW1DCp4eCPU8xvSvXS32dGkZBqdozaFBYLdlpt6cWDsxxnkXI77d5CHSYdB
N7jvxCi6CyjYNaXMH+Ed4Sd0skcdlxZb0DTCJTnH3DZZ0RLl1gRHnjMtGTYVu4rP
lp+8fYqsDZZLnVfrs5mfNXthPCse+gFrDgPEwoG0LsA5kI6UObMbLmmF6B2NFsF9
Rn2bblAMlTok/TE9dBVf1lWSg6abtoD/T8TaGuHyU1W6t+vf9EYvT+gKa3+fn/fD
utbom0EwXJ7SWRzls69aMSQjbK8IyzXOD2LF/pyIsmCSAbYy1CEBJCbz4yvXli5v
VIzwB90+0t1BlbOlg+rvoBdZeuPo/DcLe5c0gfcJCH+XisbN1yJT/j5LpFjaRgm0
fWGAKZGWtsfqLfiEkFwzxThenKdS9Z60Wq9PNWX70gmqQu/IrkKB0VgZCG+QmSi4
hapmdC7NOThb7d8x1tTlONNNgfVxhtrCsAPqGK/4bHjv8QF5pC3pwpPr8pctAfKe
M8oXt1ZPc4QhZh22laV6vru1AsEXV8LfYolcJMZhpJ+ai3dYP8nh5U4vFJXtzHFs
rLh45wFZWlFUAK9zAAQtUPNx2/BvrLThl8kx697l0j6hG1tY+mcOvP2W9xmUDKxD
hgwUOEdHmCsp9Q0A6o62qgt/5lOVM9l7VcaDAB9SUfYbdlFDIaCPzSfeE/c1z8Gx
NC5szVXxR1scCamN3ZsX1wIUIEetu8KD7i4mMD5VYNEAV4aQhPOctCQnkX76SJYW
IJhmri+0RtDcXnfLVviwOJLMrOe9ze5ln9o7kG9zszH2C7UcrTTe8nwN1WRO5JqK
wL3QHeqP7ljEoTGAi+tDGg440mVJVbeTLkiGx10XxGEj+gPzDGbxA8TlAwNDds6t
/2J7jzn6megiZ2ODEVnmNQcgqqobd67A8VviOj/9wY0tL4aNyEEpmwHF1In7LOIm
qf0DnFGQ4pfTD1vBqeIc1/F/0JRbLZxT/NS8OazDwcmrH1zekZYq+ycq82l2sLCG
M2NDiI+WkXALwxNCE2YQwNCLg0uzkymdEA9qrwzi6h8RS05CC8MrHpT6OOTvvrgP
M4wAPW2C6Q5LSEZKwUei0jSosdPgoCTChJp11dMdEAWbsfa1ZFnfZ0hGJzLyHJXC
h0A/2aw2ADdsdp+i7ndS7I5ad69BDrU9hUWqDltYQ7vxHYKqq9s8aIAxOi6X9d2k
s90pGsS/Y0Sf9QIOoYwlEHj6GLZsPvFVgKJV0MW2OOUUFOw7Z7ozpCoW5po3DywH
s6+kwyofbF1VhtDYiuht0BJLZ7WsfPgFPRcDlHBFMQvQ/sR8BumMxtvGvqrau+5z
DPpQX/MwsvLc2Yd8gW2mFpFWsJ6N9oStZrMRutmg1qkLfmAMOGJa8V4A6Lcz3nHA
qDE5wFvF6vqh6Cg/SorLwsP5feDYHTlUDnyKNRVRHNtlaA6ghku8GCp5XrB6ag4r
G5avl9ZrVGQyjIqGkSokrQMHhSv0VFjW3NpyibuYSHFXjz2PFX9b1qGyUQYYDZrE
1Ij00jkhBeW/cHOe1yAU+4dSCo95aEymkGOJSngDQodnJcrzw8gaeJ7MJ+SAZBbW
k+1xY6z3Da2axJMbSF8JtY6uu81+///r+DKvVSSo1wA6gJUFr/uW5NUrLx0Ucn8V
F5M4q605bAsuS7LiMmyOBUkplIu1DT0ZWDwdwfL4UMmvG4hfVBmAKkg9oSalfwzl
TWFcnp1cJgTFOq3z3BpHOmMT1JVujFGnoKQCI9ahaJcG3/wbyLgId0FNV0I6tgg/
B+9Ke2sKdF5vBlvakyFOVdBegXfYFdO7vlPVPwies/mBg3+IBzilSOQ5Z4Am0EFR
myJxNsyxUULN5JE6t4WFSBvS9iDfpjg1ye1i4tefHYI29M66FEcqnW+fpyPgKxiP
MkmJilQwBepHtq3uaBytfyOZBr9Mrv45INW7nVsecXXG8rcxrlyUgnVeqKI9B30q
0edjwuvfd8gfND7WX9M2dt+Cp52K2iL0KT4JBi/rY4CmflJ0cgXGh+2mk2X2lK6r
4AbszeN0uQc6Ljhz85dcetv7fOQzVbXq0mhn9I94Jhng2euIvUgxZidFdxNB8Rnx
lvmtYhGe8ZM0ANFyK6lM1tgePYqe5UELdfeBUURp/xvS7GKn9oG8+Tbmy6BiDeCD
bwtdUEGXJCekxNPi+Kqsr7hNrB6n4ca5j9E0Ga69J8unQsdnNHqoprZc/kMFgMWh
SOZzUteYvhUyEg99qlaqE2psn8K8GQD68FFNbC1S+Oqs7EsJflC4OBWLYGD1V3WD
QxxhezeWf8AhmYR0fqAIyc2gnTo1gaIbReRJXrdx3B2C2FAAX+e31/cOPguDQiwd
TcgOs0ELAzce67nWYlIdj0hT1mwz+fXlR12/qDE/mKez5eahlKGDLhC/b73lsI0A
/X5YUPEoTfHLuYgC7QKIet8k3wtqyd/+5Q/4gz5LP8ZHZoMdgvOhZbx0hu432Nlp
3Tq5wp/BGj+8hr3wbe8GT2cUgvw5kwceo9ZEC1uOWRYdvEbnlwtTiGCRbf2IIYPU
JksLj9/wPItSIWGHBBWrdZxyKXbQkjiNcdNtx8iy6Mk5rLFWLI9rjG2aOYfy/FpM
LC/SIwClelamrmQiDiaaqov5cCo9TqlNJtKoxlXacx7fZNuMJivDoXpsLtQ2Eldv
NIRoje/wIrVEu0M1Ll4K+lamnU9bhZCxJWkeiWUhSyGageauoD+foq1kLAxE3MUb
JfJZEcx3sFHbCEAxtIh53ayoUlxSK7tIRSxz1mAJp7EDj3I2xbintjQto8pZxvwo
mT612sK+8kfh51Zj07xbf89ADHDxLSBP9fIW9QrkQXDWiz1JFOMOPQKWX2I3KG79
VlMJtdOyzRU1P3oMw0/DgriSbtr2hkG/4DUL8H8jis6xQjaBqgvcZ5pCPA6hwA3s
rOyLPs8IQNoRuwU+czd6USPapkhaM/4wNWPctMJqmnlxHv6RdkYEdbac5bwKHXUq
r9CpQ1uybzeGgdTCDBGYQb2DtMHgqP2ZxRiy1hEc0jDCiDsB3mpAeh9IoocuXxdf
DRbPok0d2Sa5ar8R8MKDg0OUbJpTwvYYb0tM4FCXq87rAzInJLrRUNyLaPioosHn
dTg6IgNPpY3BULaMjoKdFyVnMS2e0wG+zGm0iq7L8wN3jLZr4n/zGBKYcrum3fh5
evj04AkwM7feOFRA/k5VJw0rgOlKULzRP5I1QvGXj7ZAOfOelQJD5lUjgRxwYGv+
/aHNxlGqW+1YZsFAEx3fy/ED7hUX5gh07plgyeyI3UjPkgijL7v4iDbeRTFIk1q5
ZMpgDEiv3kEELqGDvAvE85vo9QrcnIns1o71uagUdjQ5gvdotf0MCRmmtVtwvf7/
eOj3gpYjZ6byjDTpGSSXOPMb3ou2T+MeOWrOTlIi1mgyjh8O1SVGxCXO8DmUHQ9T
HA6e/9xpP7zLql8Xe0eLrrXGbM0uLWenj6dMPHnOsC907M4pt78GAwiI5N+ERN6M
Mo9JLOpBkSUT7IrAwGmI0BKIGb1jbnXMq8cjMNLwccpMTMG4fpHKfOKX2NI5z9dG
9qS3hYpbM6q4c4SA9VVLJICvTpUT0mEWbqNgEgmHlPNOSuuKsTn1A5LCJ9tN099h
CyXpdvCBqnubkDV/2ZObESGZ8HlbZ/qAjDCbfQqK3Y4hIKzLTJIwlmq2Ostvv7bb
OWguGqTl9oR3Pk7IgE8zpd87ggmQGlW5AinGGXvgchd4NYNnRacq36GO2gETvbOC
2MCMmZiwq9lCHqUea5mlDjCOELHFupC1diVZeHtAxH89Cw3c5Vbas33/lThCn8Ky
wdLCdDQpxGV6vec+mcw6+Tg4VJkoO7IkWqABYVm6KE7050c9zk26Kwb7rdIfyN8M
LhKAQrDcdDJJw3r07FbmfcJxfYHlTywnrxuJHjsPufbLMw2u1vAPFvdJQ6qQnyVv
j+iQPYCwoE9lVnM64aBGZ5fsQRNPsy8EtXtWuYP4WPOwoGrDVSAP6GoBjb0kP7t+
Jx18Ho/Dt9OOrhQJQsRFi3NJSMRzraP2MZK7NZvH8LEsOafOKutVjJXzt+/QKz1c
7AjX/nm4BcAmwpyE1jEgtS1wzEQLaZuIqfOqrKSm+QhoTymORJWY0UoiqrI5O+I6
xbvIh6qXq4RVDNpALTDBqR1mqt+k0CzmUNGcq0mYu4RK6y3H9NUfbHB2O0yr6Uao
7/MBSyZ/fKtuXciSMyulRlX8wyrLm9TRUVpxwy2cx10I/H2Bgcw9qbhFsTPPqZt1
vYjkFQt6IPexR7k+8tktGLJuugijhXiAFfxAWESOZqjwVdA56teX9fK0dJLdVmhk
vTPe0Bf/lJeRXF2WrGv4cNrabSL8kT2N1fsX7pjEYZ/mbeuNwXPLq73ecm2BTGSD
xnVPhRCq8LzJMTrcuSxLjR+isbhDdfFSa2JX/yWauKsng6ivxUY/FZr9cVR+q7i0
NYebQinpluiH53srAP5EH5rl3yw29xGvFqAzm7pdhbS1IjA3OdnujoiV8TXD6G1c
E3cPLNVWMVOTDBPoVK9dlsFeIWUPf42+gH358KMecg7rKTHRugBk4L3J0Ru6QE72
9C5SQNRxbQ65CLaBWEQgP4yMl65oeY0/xgqIAoVImwVJ2vqdYsSVwWwQxxW7ofjp
tBYEgnuetvNBlKd7w8nebjj90bp7zW+TqfICKyuH4qWn4amf7qtMOEeQaayLlDr8
4Rn0wZeaoIn4JJ7JzpI8X5CyvR3AvscYTMGghqaCTwSiQYHJJGd8WH3VzP47g/eH
V9/8MvXZMtB+kgBOb4Q2NZdq9tQuXAnzJ+m58SLCXlFoYhYwsG5rVyRhJp0zdVBT
5h2EYd7qXokUtr7Xi87G4kgIt1sYd+XzhqsX3kpfK79nRv0Dgt2mr85PKcegCNz3
3cknjdL3HtAAlGTYaBKDfOyn+Ayhcp2FN3sPUBBCnfUZ3HwcmEDHhO0Ogc7I1h+K
34KNHjXkgWotAQ7MoskamodF5efuzTqXi/uPGiXFexVcvfRk/ylZmVJqBWqvKg5o
F0qcRzhgW9pOcv18oqEot8SQLRJNaEYa3eQ8fFiI/AqotxJf4HWHehfh2ihhqdd5
j4TYpxTKtLs/hndUcRMVvVe9iFCPxxVVza9j/llMzHELFom6603TOywX4AGEIVNH
+uczBUqoibNWU0JYxBtwNmyy15Oq2DPuiLIaV10P+3COtDPUzHYmBOukfZMNl84S
yXgdrG5T8LJIw1v20fu61wgdKVge9wivGVwuRBpoY4s2YQmEMK2YSJ0C+gwI8qim
N/KnS/nMREH1iD3VBsrfdEus3JmlsdfcNtdHxJMshYKZIOyNn2gN1GkNEwqAccgJ
IPloj6P0ecT/4HiaMFYQ3gwh9LzkuqIlPPedBG6YdPP6UWTHUJ58l5hVLwITBVHY
n2Qq81Jwa6W3gsRpTAqbFyGl82HDG6DRsmEGngCJHXz0V6977D5/zF8JBgWS2NBp
XzFUHZFapj7NUagaLR7I5IFcjPp4gPebwGBtZyyHy4GlJg6kgI0YVePNbDuGsV/0
b3NzLdz8nBpo45QVG/WGS8c0S6kLdm9zs8rFEc2+SobenPjotICgWUZuzg9jlSuB
CdlCNcCEEG52guL4kgqZeFsJPf6rZIa9og15mkH/9j29RILS2nFrvraNwM7uRLeB
jP719wyu1597Kv1fqMgKx2r6FjOCHkLOjPF9hZqCYzQQ5kmGvdxkfR7xfLd0n+kB
pMYbCtsMDhKA1VgdHnRhqQw/9pNBPH9p0jbMbiynah9sfKiG5Yve49n+7fZmST1q
rfub112onzsXJ/d1RoiF6sCpI3t5vkb/i5dnjsfo0h4Ynh9HY7xAE54XaEI8pO0h
HTEksVmpCvzmxi12j9q9XYtJhRVAj33hZMqArXrxdtVa4yqTcjIVcjr7FkfnywOF
e7t++IlEdZDZ/Ix/wykVKijzRtzxuxIG5NFH5Q0KkhGqDevpz7mpG1QYYoori0NQ
KJ0AZx6Y4oPECO4BUgnNijCu/Y4Uf95mofEIAAguhMIQxE0jiZn8uO2rhfC0daVN
jZxrD66BJKLdkDl4bFx25hEsLlnuyaK5TNDk9FiHtvFLQQy2vdM8V9gnQkIgcW7e
PQOOQpAP/Fr90NqBkW27YY0lVp/l+gZMazxs4gsnIPE7y1vdvLYu3nQ3Blche/Wj
1QrkokWZWahBwO8MeQHHdi92RTt0MDyQFGbIUcaFFfJww886SD3RsNuWM48MkgaI
MJUatJZid8K55K+UrnICaQXaGd9OjqxZ+K1KiEnWN44m71veQPEjreoej9vw/LDb
5mxG627CPNzeR6+BFRh3OyjUW4zO0vvutN4MbEQgcoLKver4tfLj56M/x7KyoSkT
f+86/JZv8l2S0VVvZ5J3yKS6AOB3eAT4GmouS3POt2gBvNZXMTaLc+5p4OUN+Cj0
nbHu0KYoZcpQ2hmUS7zzclcmK5xbVfM79z4bBMzRAFbV1S+/8xvCyxkl/5AjMkWb
rsPTkAYHsRiCKBli1EudErg+DfMJQBwPmSQrrQytyZjCx94v6xwgORoBDWbyFTEH
W9xmjwKKW9Xvd6RBxpWq6gwxaJkv67FilK2GbM1h+xpleajEiHp9KsuYF1pV5tDO
iJK667lvOU6xO6NKZkpbnHhd6hDVBBfqlEp8qHgfo2v3aqdd8DShIHjyZ2aYACbO
I79Nuog6utNWX9neq7px8HlcnFZ5uwaze2OgTa4LsMwMFXHdYS1+1xsWF6r6Xl18
Y2IutO+A3AgIn8KmVeGVNE9FdjC7rAi+q2tBsZbtbaGAs4q90JgDqjcK0KkFOstM
VlYjfYAZWedZTd0i9wJBrWqIAyWCxaKjrrLTzBEvoC8MnmNKJDPPIxfSsHyPGD/P
PtWf049jqKRKVPjCzzy/VkM+cuTtOGta+u/nO/Mnoboec7wGdKE0mY2HNBilo2NX
w8RIADIXqfXyEGgKb0M+TuhbpuuXOvUx6hcR0V6Sm35sMlhGVihHWwg1gSxomKnm
jOH5BBra+xF0aHHEaKWrmNy2aSDCtIn/SIdh/YwWbUtEOP5iAGDGthf7Nyh/0/I5
s1JRoAYSY7atmiu9yiURgxiztVWd1jncKS3PLhZhnNKgeHDMsNE+nLmx6uehU87q
jyDQgOSr5S55fq9P9KkpIDSk7w+ZMZf1LWQplxsOjCpZ79kYD3+uW7Smp2ifESd7
+5F49F1ENsNVcWw6hK9ESJP1Ezj5ylrg+wfFRkzqkQ6pDnIHXtPFWtHOJxfBF8GJ
akUJigefsyuSraDXjhG4W66U79Q22nq7XDTOm/Fp9zVvCtE9UUnS9tbbdgDFqEbu
N3f4fFH2/E00qWk7lGAEAnXYJAoixu1PjkdUv/IgLgsnznicIe3i1ZpSdUvGPi21
ftFi/+2UD8JlVL7C7Q3yhn4Hxgifynp4wzWSY6EWjp2OrpsBdfPA/LPZ7abBTN2w
Z6ZA+hZgouHBEXKEL9EeZpbVX1WlEb3rmFhlSJscX9zYWxrDYhl+vmSYN9sp4JRA
HQDEV6AnsA8gOiipwewZk4JNduaj2vjcsUXbgsoBs+wirdxgiEpSiOCZk3SgEhfp
ZYRAXDWyIqY1rtiz2Gvhb8mjwrZGFPLBXNG47s4YsAii3wwkuVbzXJ+4MKjDitXk
LfBQsWmeQ/mfo7uKVwbVcgNcRtuAaA9aPgj4VSld/858Y4KcHLeA/BCv26xGMLrx
a8D8NX3tdtRc08TZoz8y/ZECsDNqH7f7bVcaNWi0Z7NqCaOxkeDsfJs3jqwvjOeg
r4zXvpiHbdSj7gCvJb4zL/vTDp+LQ0sSptw/k3Kjhk3lVSgwqv4uHnFEFonZjLvS
RDWuFqVd875Syurhh+/AMo0B2pIL66O+R9xBXa/uVaEE0kMI2/Hg79T9PPqj1hoG
WpBDe6HmRoMbYZyy0vOotq+FU/ORovSPF/CsbtvYZweMzXFVsqI2BpXDxeupJmFs
QjhTEuEWdQRlr2pmNJX5y04qaC32BP9XU8H5Twkk+4nerCb6uoME0Jny5Jj/BgDA
XdYWQIF3F2iE4N7QHjdiwiZCmZa0HQhaiA7UAckvs6+zDWWfrKhuCrWsht22h2kR
td8H/L6XmUV+WwKmBYwMklxyWsxdSDMAg++/Ggq4JboGoV67WZ2eXFtF+n/itCN9
hQsomwplKCTB/YuFNWvRIVZyrSGAm79HTrubs7InjXOH8fJjYe+5zro6u7nsoVP1
UNtyjgcU0visc9SHUMpV6mJLb7AThoXbVpg5BSOHmvLAgq00tvqWKPK6HPbG1pfj
kLs8aYKzX0KbzvuzVwHHOovDt46tAoU/+pSyLfvzMtlyIcGnBRh00zaXixywZC9b
tqoxvCpN0Y8TLaYAyL5uYCdzgtnk9Cmg5DdyTtX1wWLH3hGhCozB8Kt+prrA9lnq
Tn1FekYx1l1l/AKDcYxBRGd/geZ00h0pRpF1gRC1eDiK/q504evMztvVdzYS8WRN
glf1eDx8uIZFpSplo9Uzcw1RxiIgdlBwB8ywjOlZ/ytdUwGqVtM5DsF3IxBSJYjG
BUx9s5Et/A4U0ysjTKjcx6vW8PQule1NJ/vsacofTrW9xboq2itkrHSz+gaLPBc9
zUMfBry+MNk+k6eaawpw9BbJ1ahA7bFpi1xPBf3ayNDGfS+6dmqZ52XF64q7JhXh
exRRJlybQOLDTBfB9FG7kbUJYNOOkwr6IYBBaFt3OG39ivGq8KuiNIOodGuep1cG
+7oG/FS/5qL246Z4vXgj9yj3kY+5QfRaV8b6UN3eDAhoX+RcqpUm0esSri/ReCW1
A8blzgV5RP5XiA4yG4vfs8/ROtgVywJ0Ula9ga6bZx+qghSm9wVf/5oQOOdZhPER
Hj5CEjht62umOUux+Iw8kD6sqXhVwos3umwj1j3CyxRYu5NMwbFLjqMLkRYe5jkX
DLT37aPI6DQlHEarQcivBNvoqJWnlYfyDmBGIhfPSprahfKBLGcHPeu6zGdY5Fwr
JlZzVu3lJMIdQMrsBNmJJevuKIkmNVPW7XuX1iR01CnjpMZKUmhxfyjfjOkurIuV
EBC8I0hYHswrfij5DAOpjEcsJoej730gM8GA5wqdw7+re3Z9qGK5gF3dQGfMZQM2
sYBJYlXGRlNj+IDvPJ5N8AEpgldS4CaMsX+iy6EOLcarvgCuhqHzLGGWY+Tn9+8g
aMN1Ekjd4r+vVOC4s0xR92K54sNhUpETb8VY7lLB25PPABNE4mx1M/hlU64HniKJ
aEpV55SV8dRQk4AySTeBPaf3uHmub4JP1rs1SqJX2nIqlg759w7HIvVfIrz6hfBf
lo8lJgkozxDCYbchRr+4yytIDGYe5ZOi23japmBYlrj7foADO/1qUCRKwZTJgtLU
d4iuprNiCSGARU2AhGVTS6+k2IvdyEOXQQkBPAZmmLfDKtlSV22rwiUXDuH6AgGk
3j2MnucZM5gbTLsbWICjuBlonKtLQuzdayXpTsvKVFgfrXEp6IfUh9lWB/brSMhy
P7jqSi4WKwRSSN5XxxENaP0ONIp0Knw9629dm2Qhc+vs8tUnAOYmZydMgzIQHEhP
2q7/sZdmOtTAHjDvxiSoS0W5W7/0lOSkSAtp0pwbsyO/gdEzhH36/ftKvjGXlFo2
GvACu01GustdUiRDwm4GdEvJbipTYp5o670hD5caMjluEk/WM22P3CbZNuEV0zjj
ZKgSB8c+07EP7oF9qRpOwVxEdqBU3H7LvRcpTdyfg5dKvksEvlC6PZFWYOE1JaCq
kpbbq3U0qjjmNSdUd0kHKusa4HeUwVFJ5oQc3p1owobpCzhppD5i68CrPCc5JpmG
Ac33eVP5ho5YO8A7OeeYDcoEsVzqiODEc/Se7jk96bu+O5YKATNWI7NhC6jAPYzA
O3qPWiWqQNW+qeUVesq6zVu/z87l9NVrcOUXzW6zsaXrTTAkFQa23SDB4xOVN/8G
6xpT9ENWl11DeZVSrvNiUHDL0dIC+pVnqXc17np+UhORUhbSv4ExqwtQHS/wM2sX
/PHUFMwbLelASlndxy5P3zgBZzk1PQORpsE6HDymdk+96zerIjmBGRvO/AGDjsNG
qM22boqLoIgkCJ63h+OYRcwrMcsW/Msc7FTKMOEFJx6ZYjtJSL9BKb3yJ35tyncW
EAbxflUsF2zHSGwLjegaTH3flo3EI/QXUDlt8rIasK0HWqhYVi7VCNLTrGmkt2+U
2s/z/vU4dePANCMrr3Ghb8QmnFPOrk49iQliP6+RwP6U9ZGxnErhaGitS9EezAuc
6POADSgnKq3P9yCiE8GGTO7feLF+O8y4TAqEg3tKak2GFOPQgtQYb3h0+pZl3AXJ
fBsTf3yF3C34L3qkkQvfUDp3LVmjIEvIN8SrF8hiZ+3OrjaOmXC5dBs6F0g20eNf
tXyKsdGjjoC5W3Ze+ahRuOrTBTDBpMEHh6Zs8sMPv6KvfbkxON9QhrpUYuHKBxS3
+/UX1Q+VjIH+MOJE0owNhXC69AYCUFGee7ew4NA2XaTtZCR4iJ69UP4W1FI7PSDK
4uxHJ30edGlbiOgV8/I0EE4e1h7RMsD8sSZXBIvYpPoH4Wbc6UCNpgzlu1Dni3VA
pFTluSK9i1iICbr2Ax0J2tJVOa0qq8QNbWCNAbhkdehKLMfWuXvec7sOIoBnU8tw
bFb2n0Dh/SM+y9d5k5hL0NAkUvPTl9/ja4orrl8LuXKf6brqoVFZTfhSHWjyI4oD
6GDvvyeG7CVEhTbTER9jKjiggXrBSk9lBGd9/HIQVAwwLkD2SVfkt4hb+JrHkJF+
/BckIWYNVpOAtJG7T47wInQ6ys7NDA6Pcq8eS+3SFbExr+6WhDJo8Fh9S7y65TKr
bUSd2uxS2npXAppoetb8tkisMgRjbxtTWjT9bUVMobKnLnEQ1xmxoHeyl0aF8R+4
UWtdwKecJp+G5WczHGyn6MZ2co7khjQPmpRoKHW5FFyAoz150/Gf8bEiI10to5h3
hOlWQaKk0lpyssDj7ktJOl0B84OgyXwv0G1ZFhd4q/SaYCS+tI+Wjypy4m9LA9/q
k73w2Zlluf50HiPfps1DMy+ob0IuKqVYtdU78274jLWSDk+5IALPV2QJDiWg5Rjc
E4EM32OkWV58vUzag9HkNP+5tQJ3f6y65Hz09hLmWLi3DWrFZZSLfEywNsWLRLji
pxdUAeeGGcFoT0QnxfPQ05mFN405WrLkIIfTCgZhlcknLG4OAH87xVAOMUSgyMBL
16R6KRdifCciAqS4xQZFTJ4C+YoJtdHcNf+TagepytDi6Kg023i4ILNaM530JHs7
9rlmZ4wIGBA3h2G/PCJl9WWxLiFZPffZEs5YLaMjsbQ35jweCNebtWAmV9ydcZTt
azEl6tDDI09GGwDOWKA1ekYbymrdIFfSsbMxNb/4/iRYQkCRTPBodBCEevFO3Trb
TxI7VEQkMokBvh0p5VLgrLEGoCXeXc3jg1UiJBS0TDfgakUp20cxgHVOODkjMEvJ
Hb25E/bPwJeRc8InQbN9cpNboDhdOqHO44WXxrxg57b82eUPfPpdOWoLSqYFhCY8
FRYMFABXJaqMjXPsXb1sp5Hht/4wwwxTkHlbtR8cRJ3uDXZfyj7Jr/txnLKqVXoW
0SZJd7+82TihQyhX0ZqbhC8t/OCp0iSsUpftJOM6JsFD2/mbVCWHjlZN+mFnjrlq
YunkgLqlQSZlLKwWRF9jIJO2KIVBVFFIXIsEPbR6J5xUj0X2ltWlxLLm1MM44MXw
DnwX0Znj07J5+23x+ub8018mHth77WdqkAWIS1tqCTr9epQKzS0vUykXD4R4KriD
hJLiskiw6Xw4ha8+8ye7WGk4eGbIH3bdtoqIrJPqRhAk2AVi7FO0pz48wqxKitY0
Cj5qvqVleejtLKfXFJ0KGCkvOQifTssVjghxmma/GJSC2wb6PGQgSIygAYft8vSy
78pivU2dBulvVOYUhZvRGio+cZqN0XlB5P/aztwoOQ2vQoKgnK5IA+At4JGKJqd3
T8Q8SPmzX/a/bobCpsJkHGQBVPCR7nvSyhqLRqn4TXO2g+7TpaFQtDpWNR/axoJt
wJZMuS9pq/KYxf7+H5kvPzzan7cjmOOb86yWM1J/BMqfNK23VRwRcBdeuG+UWk1r
KhBknEBdFNPXENhFHqX0rHonl74ApejckDrg33jmmirP+b7aWqAHdtfjkunTGDLG
wr2lZd1IP+gjvN1FIG1J0tcAVcFRKXHXtqUDn5tizGHPEplFC7/jW2LvMnXzT6P5
LXIUR7AzzQVEeBfyaVx9MNmcYP21Opx+HiOrx9QWPmxvFyBAQngZvB5YWCTTatMM
age0CgGUIe1vxRYHQZkk45BrHW2WmQNAXWSs3W1QVmMjvrRL5qHz2K8A+2duOsYi
eOmMJ+8N23rH01gPTIL5DlND+f1Z3UftYL60p2Kn4iQrpfNew0deECZGrvyR6aBk
jq+I47EvD2YhmajJllX5mWWrjo9uiouxwIGhZ3tzNKwwyBKXOhTglfL7+0UuwkCM
FbGB7V1HbrebmK56MVu9/VlnPtHTg+3iG2EyL7cTRHAuT7jZZJtYyjOb+nh34M0F
OCdllG6QQlVV02xQUXznqP/xgwnqjIG45VlNXjSYLOuRGoEXlNCT3He7729uCxrR
xapf7SRCpGZEmh76uuCDJf1HK2ia0yUXjqdt0ZoxPR3SX1ilYsTV4SPW5SGSin1Z
SFc18O14gI9jmf4+WdDCindl9ikX1p3oxggzbhDz8GbX4AgfQGxEs5OOq7IbDM4S
sE6ktbJ87VuAJsw3fvIkG58FpKLMtbvM1OExApyuY9kT6tes2z3FF2hPRMvqmg0D
HbUHQbVUgZChpmXaZv4UGWEXYyzgMXs5PRe7sZhntj3MbXDE7CFyAH0WvHdo+DNB
q3Fh2jwdYAyPbgFqJAxwEAjtqcjMxcUx+EJbv072x4eRI0ieSxMD9vWVd1iwuawM
j3h510sz0tvm9vq3n+5iTqQn+M92AddMk8Z7azcy9R3OMHMgFDNJZgldp6+RxQKz
YzkYmPXhQoXZ+VpStwVzkjzGXTg9jJfUWEu4PMCA6AQRfgEuH3GzONhXasiZ07Gq
4IIbE6b5q4S+IAFJ+G6JLzsBJZO2eSHp8qOIWpCZldTc77BN9M8oVfHU3ZMVNZtn
vDAYW2oGltvRyO4HD6cqP+vl9e1RjnIWDppWemKHibdibfYe90sOpmc4G55KWV5S
n1FR3RGPA9cfuy0A9txmG/dQ08mIUdP9lotoerfQv1MMncWD1w9poGKHXg5Nutn4
aeTECjrK4JmhyONv2RuDRTS6wWpUFLp5hOYJNRZCwYoSw+V3JT20z4MHzv73OkLM
6/NOfZXBym3UeY6ntStC16IoDteMZZ2QgKm4KaBEuB36sYvuR7bhasND3d3pGZJ1
vReKChuldQS3Ua3L9FKEAQTZ/kKH5ZajshoOhout+ZO9Y6kVT+h84A7q1mwz9rn/
MMI5hoR0a5ZVu4CwuWz3UQT1Ae+npPRCj2PrA8var8t/3v9VZSGPMR3hxQH1dzVF
ZIj6fkr6WPX7SXJXmso0h2KcUmN2pcSvEbybZR63KRFDKA5Daia0D67GZB2OZrQ5
5Vkt+nIPF8aoBFE26FRCxa2Ohtnr9hgOkvde+O8U2SV17USMXMosFC9B5l+i12tL
NvZ4BfWj46IoMp6wTWqBoWUMqV6fbfReDKCaFZTT7q5MUqPDJj+D+k2U6F7bargY
5wsYs0f7FGBdqJH6R1QnKiARSXeU7UtEKEwm+lhjWd16XXlJla3BzvWPJf2fHg7Z
Fy6GxnaKJbU5oSiPHIJAY1vAT/veFvFdvkcyFlSGsh81RxoDTjwoM6MIO3PWF+1a
JnN/H2Oe4rgahO1dF7OezUI+9N6EgIU17p/OXjyaU9bspr5kcmDSzjHj/wZh+PWx
x9j1SrFBRaNEEzM0azrFy13ynM8GcQN7fwP3WDfxCS9HsEIiMa/wmR3wiFHGEkm+
xiC6YFImkgkz/rZOUH5f8pfB/aFECNRbP02Leahob6Tyj1jl/e5DD8bBQzbRiick
Ww0EVFwdPe2dcMY9WEIUCm/ccCqX+PtFNA61BVvHZLYqhi9exTzkjAOOyK7Y0/R7
opfXvr+b+YEKe2ynl7bYx+S478wKb1jalAxwesbTNpfMIFUJxwkr3OjvnjM+1WI0
PRiqbKTp9e77nfyp5dGIn6UNj+iNJpsFTbnYV3dM5ZDl8WZiZRKCJHNoSE+mObE1
Emny/mPVKM5BNYngxT9j+tg2rOf046H21l3V2e6uW5hfbC8bxPCCkI6LsC3pnnIh
DfcP9/z+PMBERBYW4YAu6CFqWP9aD5be7gBLPyrAi0PzvwRB+aUpP8E2DcT6QECy
l42yHUvPtQkgTWwlmCjvM3/P04Efuu0CZR9RZh1FEPNLjclz/rE7/bV3r93wUaTr
oTXY2x7ldlJLwnUcBJH+t1DDbZayvz4IplkJPZNP4dpJinSzvX5/F7HMdUWYwueA
L5EaDJh2/R7fV3OhL9mBXAFvrYLjA8JHuYFvFKdUHXieRl4oOvv+XpLl5e5My8UZ
0SRG2oul0M+F7jg+mxkbvTVWoNoDvIrCBgnDAign43iqHgaFSch8MSaBRJXmJ2sn
/Q6XatyCns2oI6iYL5EJTUUwwisVQZFHeXABbOg31kz3FQisAJRNuf8icwSG156R
AkeuQkOcd2erqc1hdOmiK5HXELMinUQU5JMUYsMWyxEhQ9R2TOddOinkcM/VKP7s
cQ/hVFgNbztu14X8wvyWA2uVFN0MzqawGC8FJhw7TDEwC00YlUKj0gVRystCFwJO
wjyaL956nwJE8rPpolgRJ6bZry1RuLpeBkEl0LwDdGtNQ3DIE2c/zIv1cFqqXw2z
XOmmkUx8LkWUQIb1CsyAhZ/5K4PDG4WwPEmsMqajRwsjUmCp9qIRuTWG/M7mYkKs
odPbPP2NsWyJMBJKWIijEYkPx7yg0tus91K9UfPEAjFtcRB4ncEpu7iO4djq4K8G
yF7VPNcN5FQoAGY0rBV+VghgXK/wEEyXlssF/M9dZT1eVOnBaZIrfKXCSAkt6O44
kInXEYFIvZzD5CrLu9u9tlJuFw/u3B2zvpYFQWN4D172VJiFds6t9aCYzlzzpkjB
omadPsK90uHUt1Ay3rDYErBw28+9HGPk0b09U9uozzUsmgTE+/rf60BVnH9bUJOH
tXONG5Ndr5UjaP/milkGfoAXdTqwzLoqACaE448L9OWWrPEe1K/HX29eDHGH3ogF
n5O7IHq62jJzJS3yshX9Tqek1y3aTEovqWjtykm1vFE18a920ESIP6bBq/vkkJ2t
Fe2bapOPQxe4Dmo/hLkjgx98k8TOcjvo2owIByLaOB1SeWApNPHxBT4vCg13oiA5
Z2oVy7FZ50sk6JvZI559e5poddALDccsg9grO7ZR1jI3h6g+Ozr/UZvkhqXbHAqK
2tNtFzRxA90qW+CmksPNuGHcbVElf6VCe/aXY3o27JDjVa3ZuzTOeifL5qL5Ucmh
yL/jR4acuMk+VlEFkJ1PnhG1oIa5quqso5X65+4lowj9Ec38pgl0RJsW3saHikjC
AzeKk6Dv3vxMhkYhZSHDobEUmn03nXVXv4mdmfIuD0flbUAiOFKosOVVgDpSFEuk
MQexRycsYot0cOVl2sygSZx6BrBu8KY3Fvpor+B8bCJ0WlnmYbUsRQdPFAzKkvLt
fQYjJEf+nn7WonzkeRSvJbtyiyabN776Agus0AmwKtkacuqAyiqbQXXk3Q1Ga/7m
hHRfnYlWFCCr5OQ9LCFmZ7Q90WOsOlyNxHabdY4WXxg5X+VoQFOk0/PAwO8VBqRl
AjU0J2+4KA3Z/BdH5qE3j6uNpEPJ3fLUV1jSUl70p83APTuh7wQWZlvqvlfLpI1l
YExsF6rGrQemXV6lADiuGmE2Y0yyxggAbjdKYV/U8ZbUM0kfuAVlD5T20294mAVu
bbS4HYUS2Al5yWciizGAVRu5G8WsiftRT7ugxnaYa5WYln8JIxj9XbphIYboPYif
VRLjqkJboPxuNsrkp05fErVDMSKYUn9bD2Nwc5GrZlywr/PcxNGMDHVPm12eOOkD
FNBD7n4JoqFCIjrxZz7TB9F0jaWRqvkh5e4xwVdUrFipbf6BwOP1gTWa6GavFSdQ
PjyRwBD4kyvyRVadXzvWdMH8JHO9cAttc13epPGNMIIP5WNvAHDuH4JlKjKIRPKa
UF0hzvaKpmIMqQybBAnQIDSOyeWBwaorMyk77FFL/SNaa+AtMEl/3mAUmq6idkiN
Nzd/yiHpczyAg6H1iYBHTlCYoGOdh53drUZYpawRcey7sAuH2jq0rkvYgRRVJ6sl
ju+G5+lyygIHtL4SadbnJIscF5eAt7lGFRR6yhul0IGoLYMfIyNunUB8tlYlyYoe
lZtEFfeK+FSECeqt14uJo2IfCCo/a6k3TlzwOOVK3LEBtlts1BeCgNiS3B0K58L9
yUlpkG3ful9Sf4FETwBn3SkMW1sxy2Jn9NO0BO7z81R4O2PrnNP3lGKONAP9TGAT
akRnB5GWwU0mvP9vXEmZdduz7Tm1yT02SnL8MrnLYThgxFfRgE2nJzQyiezdOkbd
z3laWFiJd2z0L5953oFkompyJL8St6uzb6JIOgQxsAsAoQ/taYL0oYL+3j7xmBYo
ZMOYtwhmLWvXvCKMX2wMQdpjSKCtgoSu6vLcMWC2Es45sYNuLWA+EjWMXmdsyc7l
xhNUiFddstWvDijlT8SKG0OR4mOpF+ubLwWAaejguSYc9Dekt8CB/hlxfVb/3X/e
Dpe1q76tZUBQJzW4cy2fpyNXa67a6Mf8U1md3vD19ziOAvqDh/3CNu6srblcyIg+
T9aC3dzBdWLF6en1N469n7/+MltD8oRt/tQYxGzAoPsCNxD7w5h2l3ns6QDmqqtA
mgFJsU6+bcqx8LQ+cGaYzMEG2pQRbNdtH0VV/I7aKsz0r3nvpf+Ynht6ck/ETyUa
zB1KRl9jT52tYEoXaErHX0eSRJgusL+BKj/jUTtTm9VmELE3nWsXQL36Wf/qxDxF
JK4S6ntTRyG6ImfV3RJL+f7Y/itxgqTBMOS53dOLm7iJJGSP57cFOZIrpQw9O8p9
l9XxLioioTQsaHx5sWMpKkK04qViHTmiBf6HJ78W4wSruIyUAzrh1dEoDOXqqzbC
/0NsOBoJiY5Fy8puRM6jNk/t1h4g6ylirgnnU2540xMuUFesPeT2lKy/0FU11V+B
3C0j4oqrRKa4Ko0y2pkZCS90/UvS0WiqfIHrCq2XC0CMH+wrdhc0GuJMPInyYtD6
4rU3E0T57LCU0t8fBFjG28Qb4o7gjUN6z85+AuhPeUmqqu8GdUEMODC9RXcxOL9Y
Fveev5d2b+EFPssxDZYhhrAWAMyeXHLBZJuqjM8nmxVWPU3lc5ooKgjQWIwHmXUy
DsxZg72jKa4Cg2ZUfyYlN/feUUd4+xCvvfxaXb8rgGAt6EoOJKJGspO7sTE6axDG
WdFLC1gUHFYS/pCnLXddLop50jA/B2uT7iMJyyUHgKEq+nT1JI00AP5QVatvghBH
6wuVHXiJUgvNkdv0XpjcewpVV0tvQ/VPvNggFTREFFF64Upj9HD7UuXq4/FSNUNG
E6N6fNnABCeDKCOPUOeGpRNUUnAooABzYPV44gFq1tKH0lTOxH2NfHzV0IpYYUN9
RjwpqHL1rAZJNPlOwkJnTmoTOI/g0e4BJdsS+ZVP6izwx2mzXHktVRTehFNNM2xr
VUrP33er2nYpANbc0hKyC8v95jofWQhodBrchL7zkIggm8FJtqoAbQMkvHjQR2La
ewctk8AYESkK7HpQvrXZ82PFHntX/oirM6IjOKS+DmOskhwPwwNqqdd8OJHwrrev
DTrjK1UujjHQZEvliVtYOVI3avKH0GBiMER/doqkqg96jknZP9DxZgrpC9ITWqqt
MGOXxCfIkg7H678iYlRZOCeoRfYWGAUZPOEFZcKIXRYIt6LqQQwhFQWldXtf/daT
dc2EIk6D/QfA6MVmEABpicadlSc+2Ad1eQdFnQBejVsduT4GtMyohBStMHJXhNCX
vWhxIcqb/QZ0ySFpPl+fDJTet+51qtdqmv1K1/J52jpUoCS/MKE5L+EAzopzVGWv
3GcfxXPgbpZmohQucnHsDojyna2z54We4a54vZibyO8vEt9b8ZQZoUqFnekcsN82
Ihwggq2vaVLqB52h9ajpwex+bPBjkhaWS2jYNodnq0tXJeDHtZ0eq0Q4m24k1CB7
fJD6O3cmefoK2kCzhCAwkrRMDg+xdkksLJdyK1YfP/ERO49eEYRzGgALVN8Xjuc2
jN/+sYzkvx/82VpXYSNlJHnExz1v4UPouYjCtHkwu8orW3wYqNiyYqgrml/d8cKE
iTVM1wyrO46Nxu5TGAloz0/SZ4KhsGNPXcQS+o8BkcYB1Iu/AH+dxzgCWuxhrMC7
S69lu0NUBlKmcHZuVdNk27oDbfB5HJlxyvpaHcO9V9O90goPk40pGPqHiDydOfdd
Z38tWrsk/f6ZzDLnlqLWmURJdOQVqGqPTo5/2C5xTRbmlNIkS6ocfI/ECCJcqMXH
qyY0yP9sUxSeG6u6IoGkbaFOhYzvxhBaQ1AFpazTOD1n4kYNtcX1h1+frLE4GePq
liWC5uB4rQ/FvGa7GlbrMSs+J5QswR5SOdtKQ6Ay3sj8tfZrBhNw4cWk09orkuvr
TsszXtBd4rksqhHPf+bvfoFaJZR5DkgLO3bKyPHorqbJyk4bP0TcGqid/PnODs1K
x6cHE9KtaNgnwOPO5OI+Ovb0rdypPXBQwgh+LM26H6t3oqpADDmIwMgDH3VbMTFj
gceLSBAG3mvf4waan3z/QhnvAWgEm0FyesA6dF6FZCygN94FaH08xKAecxGPILbK
Xq0E62r2H7ns0DWKe68bOs716lnEmmy0VGJUFu42SPvO8Q6Z+sQTQEGMRBAK5OoS
Q4JNG8LLOo2OL6l4ZUIidxIuc6zrdFk8tfYrpYkSpBAbDI6oU0kH/wsR7S6jKpSj
H3yKt5tXMmftmlbHWvsWrdgqsibZm6SNw6dyVNiQam9EER/Q16qLIhG+meehnR56
smGFQUGZbrEzb2gWrXXY0OMhMQpG3LgzULb8YggNZ6o+1Ps1vrVpTlBqMbBsZ96x
RSWL8kUFFq1Ab7h8g55IIhjjQ3FDijefRKGpkiXdCYw0ZBpkOokBcXWhBgmlXzmr
0DrVqErxVqYC9cMyinEHwRLvAtlPSKvgWL+/4xxgCs3dpTJuZ8E9pjdpJBYttw/i
N9pQ+LoRsOrM1pHJheEEZLhuD7tBAmRo1HyZuG10Aqx5M2qLS6C/c45LDoTIF3k1
lDwLlK1a6NTQzTqTbyTPv/Lng7tC+S+JtXxjZE6oPBOxL82F06FD2Pwel1QncML5
KtqQSg2E3sQ0ux8x2wWxqbaeLq+TqAcm6PLQWkCOTHMgJKF/vRipvMGrQ+n4x7H3
4YYA6DSXxPWbd2fehwLDV0VX100zMUr/MrjMyzJCiB4utCfLK4r/UOTajXHgG/UT
AcU7U+wpV6QWODA4ZgeoaUxZdUspvbiZylNVTEo9sUxa458Vl+8G3eWxlHRywiyy
K+ePKHrWXFPV0dXpBCg20CHYNnIKTfZSweoJik6L/9cNiQapoCovtDsQpZTlGq4Y
zZQc4QCoQcIV13AOaHQmEPyqGkHJ3ZqWe3ocwDBXf7Q511UTEIaG3+hSuUnwC/lW
FASgjsCTy7YGfh7mQK6WQ3YCgDAzhs23dKe76wozM0UABXCcEpwdDr/DbJpXuZwB
27BVANKP09pzqeUYOA3QV2Qu2zDrV98+NKlnNtKzS8cnWlPORs3CUdEGAnwMJRbQ
z53/7Zi8cTlgMYPSU0MK6LlqmhranZJSZBBAgyQNpGFhVTEMhfJTlROUzSXW3+6X
08Hg7E21X4wxLVv/xTweUGYdJfFa4KeFn8Ebd0jQ/78c5RP29ZEP/dtIx4qb4a4z
Cs0HY0d2O11MwG8hfj0E18BItM2px72BBGH1sByyUm8beHjLbPDBnQyoXLaaj6UI
Z6R1Fnpn99kurV+I+DR/t0czo+gfM6Sa6WHR4fkSQ+vAUTu8TxRHFVsTQvcPWHmy
AYiG9sdY3lm853i/bV0LPCbRDyrc8Z21vCca62IuG/0kFN1PRmQUft5pj+a6j1NL
mZgC1iUPJWmlerdCxEQPBKsoPIQFN+lHJn7D6sVAAb/OexUnwu1jsotxx51WK/8X
uC7xWSEtG0Ziqry9NV8m6SJDsEqDH3t3/O4O/RTX8LpgdhzLU99Yqo74qLpKLjyH
ihPR6QOaoMj0eDcbtbhI5y1W0FMT52/qPCgbge+vslZk9QMeLpyDKBF6TVlRKHgw
fK2Rfaske2xrWlYtRHJs/N01Zb0z8JLyjUDxfofsfAYtZVP30nrC6dw9p07Q5yi0
KfPcBynlVun4js0132HEt8PG03wmZG6zdwb7xYQfrbvVQV80QePQ9kLENbkUhlW1
APcPUGbtr35d+Mo3sLdtt7Sep729eSN2XoNPpD8bTyfnBF2XqvEWXkTFshwrEpz5
vcoSBpIBHYCC5o3/lwMsd8mLH4abG7CqtvoVtz9YbG8Aa/3QuucoM+z72UtuTqec
o4NOPUUc43zsj3IlHrXP53t9nm7t7dVqzq9s62sVJh+FCo7Q7PQGDvLV8kLn6lu6
aBJln/+y26uO3UeTgaQVaUg4D+eE5f/nRwt4Gue4mMHKthw04ADHi990tHokF3Gq
XZKoIrst/oTcDrxbt7KR8ptYfJhDK7u7IMV+pJCWBPdzxO7SHeTrISYnCY1pHfVF
1Gshme5+dg0fD6DIWEx6dVuXRv6SgfVc2ZjnX2NtIIfpGKDCsG537MJUoGp6Fbcj
B8Oh0TNHmLhP0+1kD4PJ11sOTRn8BNHR+HDHmsIbgUjkgD+16QSdmiS1A0T/xDRf
JWqQThSmRANYtOER2zk7Oa07p/tNcoJ4rDDjqOS1K1wjuv1/EJln5TTvtd5+UbH+
qu+ii2q3WsUeecmu28RMllIt4P9a5AADLj5O7pZNL6rk1ju9p4ikNZQkGhUjiPAz
rz5/zWxhjm4Q0quB4x5TEoBrnoQudrdomVeuA2Ql+1W8C1x7HQxfu3ttMexBuXrw
/I8enkawHXNuiqczlnEIKlPWD63veOAttWalEsGgxeHj/0/zZQqdlXo0/ROc+AiR
+M6r7rzyoYYa7b5tY7rvk4UI7simNNGQgwgwhI/LABYzWs0C/VtbtHPPyp25cEBF
X7brmT7W9oFvZmCpZu1SQoo/8BFPeuFcqVvtwQsd/XLVxlXu1TjR6Kv1DrctNbAB
VfEoF2Y9dppf9cy/kkXS2pMaY0xMleRuS9oHydiXgcxnZ9iZn6krq6sTJuoKd+TD
OehIuyz5xYcgRELCnKFoMVN2wbVq1aiNmJAzzyREdH14D08Qy8//npKLX5CUl2Z+
ctiyWtiHuDBrvgINJyq/GAykLI48ALrDZ1gWJNGn/8ldXDbctnEq3RHdaXCJo/N/
jae14St7MlAamLS3J40ZRBtvcZFirEPThiTlcK2XDE5Au1NzWGaePKYVPU+jLM1G
JN7sX6FXkPJgiJq2/iARI39gDihGJ58fYOaOmxByhzeCUlyDkLKmzBfajiODYO7r
uF5wAJgqVYHtAYSQ92mrAxiwMHoF9FSM6i+NnZ9gW18nHxazPrRdNs8aCQy1457n
NOzwCFJd0IB8HSimm47ww5D4kpm24NyQVJHarfOCB1roTqQ2sdM97bOjbtvU2WbR
F+3cXrl8DEuHueC3xxUJnilaoINhbw4Am8cd6jcC9hZNaqUKvMkyu8I66XWYXH+4
t4RK9QoqjqOhXh9ji46ZbhDtKAPKUS8jbMuH0bx0UeBJZN7QNbikXm4K1L4ZLH/e
NaRzENM02j3dDgxoIR/FJ6za5/C/JgoDFC9FcHnZRYOUo2LfU9esjDS7H6lWPpUC
QyevvqzIifxUbcOi/aiJw7sYodoSomsJ86RWraJsDZqwLgitjGT3gzla/my1FoCm
apfsWYZxd9Az9o9UzqrFO97YsQHzIX91EY/CaIpe6JfvSPb+sevYNuGlkyLdJ0Yf
IYOQEYRkryecP5ZVQuZHfh/AyZ3jINvhS/8jyQ2wqDG/woDJIGH6nVJ7lBTMhY/i
lD9DSylsXK1Bc3GQHfezvmGO82mnd1RaIEY2MqHiZEWrAp1pzOi9msZy6fRDQvty
QkhZsDl9Cs4HT7ifPW+6fpPAfhw4HtmEULsP9umwMjZoop35az1joP+bE03o2858
VInV6ArohMkbX3leKW2uDdVCKt8CyIdHVbG1jx2n4eKI/NuJf7TZBM514+4YM1W6
Ni+ZiZjUGht81IPxIpbHFvJoFlSak1AABzUmgkk6KSd0H/CH7Rivi48aRtX1sIct
GwOzenRIzo7XorlKX7h6U4+I64dnzQPAb5qGCb+TPmIShPgoJaLtea5LipPAi9y+
Asu19OJOo+8XSt/5wvN1smZn+I7Lz9fr/LDyI4aOfyEpfgpriLrluQDVrvI3qwGh
X3BN76ZVHYygsw8Gb4Is3JrmVQNb3CwTa286Bnd+gSgA3dMlkF6oNBgGNteSG2er
hN9aOg2BQFBKizttFwiVvnTxX7tmYHoih2gOJL8yH/sF8wFTr7WIroHYl+xcCJGm
kTbSZngfDruHMrCDL4K/xzSIjX/C8b1aRV3P6rzICQsYlrtCbphcx6qeEGj3sZUT
9R6I2fEojCQJdpYYaGobUS9gE66Ri8olEM5zCer6xgtQnt4NNDIji51GClmJi1cu
4DZnlxg1cWw4fMMVYkahhAOg+iiQboulcvM3j5cIPpt89r2WRuzBPVaa9wALjl6r
7xMhsYzsZT+FywJ3tqZILL23deD/Gv4XW+jvn3+G7+DIRf8CPteOUYFX96sMEd7W
tkzy6rCv39fAmGj6A2lKMwErTH1hpCxOS1fzHRdxKTqESJofquT6Mgj+YuvdfB4u
Loz3TAPGU73SaUB9MQGIuxgvuXJS+DzHw0/O8/g34Gau6nnYDtDmFH8AEWTRCAdM
4SGTt8uUgt136YNALvjevpSbQyjUBJUuWd5izLfROSEmQoID8dF+YKj0iIVd7wEO
6VezjPBgbPD/oLphC1sfd1cTxT8Vw5cFuKr6rxby7pGiyB9AZHuMVStl1YG6bJFv
dpHouS6RJOH0jj7c+a5qdCQU2M2btOHggZpk5bTUc8Vsj5TlvRGZby3iOiyM/nHR
Ptm1B932bQpgWebY8bcoq7GWZsiUeJePwOTRIwPMTD0bCiEZI9unY9xjYkmFDNnG
ymCaRzJQCO2fgWwkZ3vuggcGbn45EZkXj8QzudkpwhFzc7ymdw1nZ2XTZyqPQk64
P0DemrFmUCpNdm10OnUO3r6ddI7PhM8e8fbvkVtQFjzDz7jV73VCs0cv3XipGzxo
Yplj/QaEwxmqaD/SjrIHR8uPTvwSyet+O234k4NH2HGiwgPVSidbkA7XBWkLvAEs
aZyypRdeP9Spf1JeM/4OhL5/sx2yOhdQLnspBO7NFVMhTkwSHrQHujmM400ebbDE
UtEeKTrEL0FNCxdw1e+bkx8yQgxMOxhN8N9pWNj9+aC2egxGKRWF58kZGRCxT1U/
8GWl/jD6GWvvY/uuJYXJdlM0eDVp6YtrrM7LJ1iFdbeuCQvwQ7ngM3WvBZnFjuP1
ccbWudNw+EVZDmXQUqIs0cGBoXKJMXbXVj/dAGs2miBsKxInWfm4J8ys7W8zZx3P
IcvTpObeVHXuBZolOH+VX1DvL8HSiQZM37nFR9V6HquO33Krb2JdX7DplxfhP7xk
Yhk9E21DSXQ8pgbStU783IyAYNKAQeZJrXkb09ITSQ5Q968hrUlU+Th46yffgfRU
fl7xRnJwXidNrhzWiaiLCqxKdfBnuU3qOhy0XBklTA8cFKYFtQQRxIxDECllZA1G
+ZMzsAUhQxjccxRZba1durIA6UPq59RuijempAhzQ+rJT7Yvexb3UdP5VgjUrvf3
r522s5U0W5XTne9POhPDNaaUXtUVg5jrbzFYDwP+gdraj9Cr6J24xzwMxrkEXnlX
U9kDDsb78Hvp00otQaQy9+DVAiNv1dlrc/vPVKs3ZX2oMEsslkXmRVoDCbjs+Rnz
dA5E6VVxdFu8lVsrsWLy1cHDt4jTLVs4SWutkKam5u0O72ollxqjcr6b570nJcEi
TSggAjeqSFxrdhOJmaHqkb9kfxjCkm8PxJX1Ph6mjBvcYcHeOYwyN+++bw+/1rzP
an/ipCH0Vzhw9NhOaqZf+mn8JzJjKRraloFSVcC61I0Sb8SeAyPPbe3uGeIkAD18
0M7a4i5T5wc77p538fdw7hfY43jGWFBU6N7zPHajmTKLA1gcK3c4cXy1bIEUidaD
9l6C6lmsT+vRuZ+PgVlN+fZCOJS6s1h956IXBCoPnm8VJjeOQ2JmevofgdUeZZaa
bc4uiwNs+fXr+bEOTTqc0p7oO5omNB+1WW5mnDjHvFNpwfWR3q25VrXLYzIdlmrM
op0O2xkF2LoP9ExGXvk5asjfROVWw05GGxKiki++8sDX3EaZF5twWE22jPdEYXMk
UKO1BbdP7kHkQ4uPS/gzkwZnBmz3I/AhZX4P+h6CbGa0UwueNbI6tK4bf/Gap9Ie
C/JtWibrZx2nXf9UAJ6KjGfaldhc6WaLzMuQBSr81wgl3d7D66oia1JD35WG05D4
9tbNcf/Iu6ALtMs9UlDq2CnR9GdCzHuUp5/pFjTfbONZYRJBvyvuYAImAJGvLdgJ
kLz9LyGefMxO2AacPmzmlbpAEg4D4saUueTLHRvZ2NA74nsf0gY72XEUJQtQUzKr
Ulg9ajwHgSS/WgI6ROnmzTP4bCVVcCR25brIedlh446CkMop2dDbj9SODzMTaRPX
tMmJsx4cNhhU6y6Zl3NIZAKmTWvooMeXYGYrYvd+m68QAyW2MIgV4SdQbO698a0a
a37/hVfcc2DmiYwMlFMhRJnhQvZyPjwF5WYCNX9oq7Ybhy4DYXf7X0+huzAmRVSY
Mj2HC3gsQP7z6U3CWnYKxVmbgRjZhyn+FtA4OHJkxsaAw9SOLFZ7w5Ej22r8GV9J
KLhUesbrg7nsecYSfXoQbpxb2yBSISEb+KR9AMFGDMZjpybt2+ZOLa7i+vuNxYRh
dG2CQdsqMpjr8r+Er7CeRReQf7qh7EsA7wgnExbOViKAKFV9ERV8FlGFrsU/5W8e
WQL5HeJMCkvNrp6GUQ01JB9pqmjHhLCPNqxk77H9h84IDl1EnW2EHTRKEiiS3tFc
0816Ib9wjrViseZdhlHy3Kd+9AprAzeWs8NL42TamjtH9MCLggYQ7h2aqZWLyXv0
K19NOLJJpBPGHB3j4kBz16ounxpo4/WaIGX2s+QzZYONmGeePP7gTY0DdQSOGvgj
uC585/ZpaZjS2qAow4g9FJ/EieMNtqI9UII47vOVn5oD4qEqEggygBZ86BDSf2+Z
KFyTJz9v1ENo9vPu6IKjJHvzSyWaFqagpB2kBQEvy4AE5x9ijhvYL1JJINW0Pz/Y
2key/NkIPdxM9ltp2C/Z9nJ7wZCu6/LSTIG77YV7CumGvqRrC4W2UcM/4h4kmOu3
kvQcjS4OM0QNPuSnvlZpQt1o9DqyCUFvWCimvrG8G3+nE0Sb4/tcVfdqXLBwP40M
m5N8kX0AZZ7wl1/uaVVEOmNCYqs3T+GX2/wVMUN6acUh6OUtKvY69txcy0DrNCAi
gEquas/Wpvw8576hwTruVupnvfWw861hh52oMxU4+U+7NHASrfg3jRnmqiJEW7s4
A8uytw8NEEGdxDiVFNULSG/4cImuvIUxgYmI7wxdpn3Y+g9iAqFp0YIrNzBSgFrn
dH/JXGwsE1rBI/VmQOjHnHSzLIX9DLPbyytQmtpjQ4aJb5sWM8nn4UUUq4Tf7llN
QVjenH0I84+3VRMuN4PxitEJH9FPqXbSTK92d/E1WPL4U8f/5+VVRAc9eu7tLfSU
9/rYb75h1KGkU6Vj/uyQaljmxS17eVGQDjP1NaVk+dWM549vam2jCydWLypAsyeB
BGuf8E4EpGiz9YyMIX5qzfzQ61t3zyuhtOmjI7QOB9R3M5wowUgY740uSLLoy4U0
yBLe30byGgLd7AemFSvWFiTwgApGA18AkcvharnTuQg7pYq5Vr6j5ctyA5nIQcgR
aHPM2fRV8rt9xiK+ucYREpuJQNLFbMD5fx1ttip+IJpwKF/S8O6otPT1oTj3YBcH
MuRlarOsMXC6v40VjPocXPu1W1Z38wMzS1pErUGrtSkmsHN8d1UVjZH6T+ndRrv+
ZdpJmfaBOk0zvmOY7I8sEFz9hKrM4IrCjQ8sSRBbJtssecX/n+zsHWgTc6sBqzWb
/rWNSKzHo2NzQraEwECoGkXNQt3yVy3V1nSLoNfDX5qI1Ti7no2bculz6Lfm96BF
CdFkVLeIDClLiVInbqdEKI1cYZ5g+aeHdIfFv+0fQVBDUBUbE2Zt4PQmFL5JrgNl
xvavypfBSGhgt5K3HAC7VBxQ5P7pgM93t6a0fxv78rX7bOUrwfct23n3WDfz+q34
U0yhEeoDIL5I2RhossN2j+geDGPu4mqU+dnmgiv2422TywU7UnH8Iivj1RWiZbvX
9DR7jJQHcfs90KnDO+ngAks6SI1h0IEGaNxpnh4y9HkC+a9M/X0YlvggykP4SucI
T7BjvrI0NdOvP8YxX89yuAVLBfvzULYEmt2I+O51eF4cK89wL0YqPj3jPOu6eV8K
RrQp1l5kKY5qG8ej+2zO31jMkwR+yrffX+b6LaRmRyLKFllEl/71opCr5bIzlHc2
5Pz3H96shmNp4N0fvTU8IktWgvwxIbuol2ulL/e3iS/2jkmyfyvC6AVTEuOqz+aw
E610r9+9otezyoyMuWo8bBBTn/PGcbekzwKF0mDu1zwv7wNdDebL5RwCKCuJLGbA
9WggfrYsvbwU+/7RKVU6WFsS+9SsCMy/pesIE3JLFZuBlrHC8iiMnkFQCwDxoXT4
vRgC4u+rBiHBubqipgrkUp7iDRQyROXaHsUUE3N55w+g+x4E2wylepl2QqT5oBDe
GiD/5OM/vtBz3Z9jXxaA+1xgktfRxS9vHldzNeN+XglgLctV30nnxd3ZhLoABodt
vPhtwdh9tYp59miqxE2hr8Y+nplho86P4ZNxNy+YPXTCd9Va02FLa6+tbDEq8FZK
Ow7ouTeEnHbkm9WIcYB1HHmbvOTmK0kWWx14R2KWMkIq2LGrjHTNSWY17Nxq3fXw
/Jpmz3ENf9EJowTHvmsawvAkCgD7Jcg1naH5BbpsmW8QQqJJXGmkUcj/kYrzx2ek
IGYOZHDuXzoYDplgVWvvvBoVAv6IuRw3z7LdQmWIoXeboZWDVPWIlpSnKXuBA1sp
y3fkZg3HWaioUgZVPjBsFEVpu+4JRHgBIelHCilBWjaljO25gq+YnNTNbmlepLe+
g3UXVcH7Ts4YWExCHf2t9fV3kYmdATuQkidfcuHZWa4hX19suOpTHb5J27bQJYMQ
GPUrD+LrPlY1wO55XqpxGLj4Zw4SxokZm9ArWmcGE2rKE2oXOumuDSdqhVnqD5eW
A5vDAnp/nwHFblCS8HaqslWaYioDNV57IzaqmhM79r7worWFzHQMdEqS9mtYucRm
Wfki+SVbZeGLp9i+phUzLmNVo6HNSebtj7XiOPPmuESsW6sS45YeeUeGL7/7lvP5
tFD+3YwQyNbM1v10nmpePFB8x0DM1C2kZPxF5aAlsAJc+PwGvClQIyC7aAttbraY
0+eOuY1Vt3z8GHhE2KrGk10ILLTD+7VWlIue1+O+PC7o6j/GQmaVYUTeT2sKyKMB
Cy1rTAXowVk4vlHygvZF0xlklApqBcIpHhaeiLl2hpsksOWFgkwqBgUepPJbi3al
sGck9QKTYAbroz0ZRmItT2xXrsumHou29to7Pt6mjwcPOwUlI6fMLUYz06EDRHhz
/lEYizSjnOUFjQN/Q3pdBgI2Kt9uxEayN1MyXfqJFAhhoQMr/SLWVo41kjHDYmiu
zfG697PFLzQMk+0PsrSVIxMtSP2LGtfcgpOnBKnUidwQQ17QpnURxnLNJ3gD+z/0
F0hzJ77+TYD5jy6dqq18VOBN//nX2zNsEVLLyW5xJ09y++HRqMUiw2sGBxqpjXY/
zqygGppiGRQGy5bVg9f+xSCDUQDH3M+8thU05kpAXhDmJFnQ3rtieUCeMHOGzrj7
qdAwj4jhRRVuI+zxbU0XYe03C0EqyQjuI+njRaVDCdRvqhiX0sMXuLIfV5pY7SjU
Bm83H1EP8HBJnZ4IE0sZIQko33d7zwL4mR4aGRX556qOMtQCwAspvcfpmMfzrjpA
X+uDclESQXeFjAv8pyYfRHQRrFjFUbCRmF9DngDULZmzpZYwXfqCZsdZ/YhnGWlh
eE/Xaj+71UUco5S95sgFrgJnpLJnlhrpbwelX2ETY9On1rvTf3fEI8Aq0L+WQTyY
2z93gjCCsETVh3Ug0X+vV+UaZYKqqh3AKcVAbNVcex3NbOBcbJ2OO9CrwO5sgoTz
800wLYmAkcQJL/E2lsZG3LuYWh4NwodN3yiWNsOXwb3CCbqs4uB76VlEgNdDo4hO
DpTyQO0IFZvNeVpGrpo0xOFsPHTsmUGMj2tzHf+Vk1zObTZsK39cysSrfPxLndVR
fWMZaGi4uFxUDzyjh6fy1+CBM/C0j/b51FrUCoiD93XQef0DC3Jn8kV9T5M24iz8
AVnOcNP3ZSwxyMnVhmWLayL1pVYIwuVNprlUDdfIMPO7tGWgyPkOrOoOVVHBxLWN
naWuu9UT/NNA5PrWIxwvZfmqgCT9K/DsIyx40hpXrX+Vx5dI1X53edWNc0ZPM/NJ
8hSBT32ct5RVEW6KXP1hKAV0CXu8u94xURI1rn6hq1P1Coe3C04+Lk5eQpX0468K
vYZ2j6xbarkXD+3NYictOu7kTAC53iY9qy03GmgGO3OxiUzR7NTLU8t+AKNRHRA0
znBddUsnNDZeZkQQ/qbpeOgyGsEIFcbZtGgCV/++4EYadx4gNyXrYDUy83Ww6rv+
p792xiZIu+z6U5JIE6OLEEYY15tTBCNJ1q5E43PgnHnhQBzqSYbcSi1Z6cTMEua2
qmkGmFdKn6iveGY39kR7Z1uAyOhKTSasG8GBPEBxFXAQkQyXeZ4D3CxdQnm0E/Et
2VOIYeLK32GAZ/IDTHG1D/cyV08Sa2U6uxaXpxHc4vguoWvup6yzGirlCTxNq7ob
rTsoymFZnKvV2quCbELHpck/eo+b7yxMRNWhBo2dPrNaueNeBooO4UChcja3i56X
u/i2UlcJ/665QVMPJql98Edr0ijji5ZEpPTQefEa9MKULfn0PGMA0oA2j5zQQbpW
/usDeYRqHbcgzx6G64d6DvxxgmxRLQWFrL1yb8xxk3SbXkfq+fZat02huvl+J0Ur
aEgUYBFybDdTeGbEXwWT509Y5AZyDVUYASUVW4sRtLBzBlU/+hle8DJHMGeIib0t
VimVqnZB0ova0eztDwM8x7wqEQRveq7GjbtWsnnkOpdMpX8nC0++FcZjzKoLe0Pp
VNEvvXG8SWR9pqWioFptPyhhskK7Aq3uPJqizXJctIJ7vQ29Ghh81NjcaPje8S26
/oDZyTvsK4OBM52bf/BcVef7ZbCZGWQUAY/l74ZSGfnlNYnp6R3dMXqEPOEdserJ
hSRkBty9PLfOLiiairJvoV7XbhnOQa0RJ/X5Zp2Ovhifr5PdoS90XUHSTc4+rPDa
GH1a4UuUHUsmNewrCrLI48NNBUqVKjTVO+8uTUPy1tfmnoVw47EAljBzmihM13mm
dzZOXFBBKppUPd84RvwOSLMYYxmD37XhNyfIjsyDQoZ6Mrey9aTVseUYuEMEt/xW
RNx94ixiP2WbdsvQo2hqtvCaYjnS88MJ1DZcnef0RGEt1o+UAS6jG8lq+za3Nq75
T9U0oDJ2kZY0j2wYB9499liorXDR5DxitLLXGQZd+m1yXQ8fGS8vkYU4ryNSPvhL
sseRWPcgdx31a0CGshQ4KLFn3BtCMArzWapIYbmxiVWMcMVUNTMU6vuwU0WQX5CF
BeSGJWGpdKNAtXpIdoTtqawb/QMRAOIjLjX7X9m/s8b7k8tl+ZoVFfWBupiJb7SP
qFZTjKEhqjQ/Nu6YIv7akRqrbXthYznE03r+jFu+euQFdqdtj1jI6n8E+j/mvqR+
HtWmD7XaytfZFks+p2jZu3+ziUXzwzn7NsG/0juytHjt/VrTchQcX66+4e9I+MFc
+6GG9g2OdLeeemP7hYvp2RjdXC75kQYkh7j6mAVgSmJqeK4QHW+Qgz3acjEkrgYr
6lxT1nhlW1kzdTVxhuQh1moXhjLhI/1DjlbfWdMWdRfrGZ4mhYZqAApL5MMuAQfG
/xVDc+SH6iFIKjyLBLh10auGam27mMONQ1ijQpuzwOl8UD5lqRE5/yLYEeUWfPDw
BnrQ8gb3AKvtSxhNonfH5jCJPadSU/dpL2xRzqFnMSZmz87lT0ajvYhMhK74YFqY
bmGqdaxeHuwVPzodj5oWz4e0GTqGbhsOwSSTarjfiLlMh4TUUuIYil6UcmGZpaYz
gtEsgz1G1DYT9ZjeQysZhUPeck01YGObx4NtHd4+RTkz1nARS1wD6VHP1IZRoqkO
ys9qAuPztPKjSDgdWvQ9p6MqtnuOewrKBPb3PiVg7mP5dqbLVjyYlnkiT7jlWzSJ
sAnemaK1hGDL3jCe3DQqUsAdzlLuFTQjqRsFEEHG1CdZF5CielTbR9BfkgdkWEcC
r/HOrCMBDPdubmq/p5UXfi8Hl7b4QNUlPtY34+q/dlrZjPAXUEM08Ip4m3eM9wXS
Rnq447FwpuUJqU4A1FNSHOAriCg4aP4Hb4uM5LDH7oy55BudPS/GwNjpcNW54Uvc
mLZg2c8aVeG4ApZe6dgtJ/UsgoieKMXND+4BPy77ymMo7MR8Ll8MGSAhY6UThrlw
v5tKxJQDyj6zmKENgWSrty4khSji7aDZQLIe1mUGQWyL4nuEqI/wmE69bJKLC9Dt
XPeLV4xSuBx97ZDqZ/aC0cQqRBFmzrfETBuvpIfTeEajqFG7rhstlwc2zw3Cy+ht
H4t2M6kJx5okuaazDCvAWWGvAaKFCaYij6tOGB7+hdspEr/p/lw4Q1SZsb4I+hfi
J1X5PJMZUJblj1Sc3JsueD7w2pZzMe4ehrFPp6o8lHRk5sYjy5dLlEyxfJqm3TjO
BAP7n0t4I/Noqdt/BfiYvJn/CwULhMdj6cwEyVtoJQgXaL8Ce3TTEhbOejIVBRZU
1pRgT+aueF5Uh4JmftnMulEo1d8hJacFYrL5C9GW3Mph+fd8cnUPERz6yjfHRqCr
opaFfQ7wNOqvCTsObZufHwVHuUbDHjDlXhr+UhP/3YQRRu1A+NpL7NH3cTO01P2C
GZfdL+q+Ipq/BrEQhTwGa/0LCRKhHZlntxyxXNVEoauLKSFJNBzxX0UrmwdYTTgW
aQc+m3fWDR0zkQFFtRWVmwdVnPZdgFgzeiFhfYTKryYHWR/WMCgRWUQtkBwjx8VP
6jJoIKwc6YztuzUmzPACsYpPlaFC2KDnNAPtQHNuQ/HT16q+1QjTEBIFPLMid0uY
4EngRE1s6FxwIbZtc8VAIlPXB586HmBqNFKh1w7trc8kTyNT+raBhIClKSHpRr97
FiNo4UIsRsd0AAWVmwCcyd7iOfusx7UIVkCK7lacnhGidbIbovpa7jeuVTuMOyFh
MTs9OX6zqb1wfKXMhU/5DVwap5yBUvGSy0H8cm8M3VLQLJHh4L0v4f4bq1dxs1+X
Vf6fx/C5KiLTSH9a/DSTwtFKHQrv+HQjzezK/GlT0jOtFvZz8E2zg3xi+WH15TM2
YQvNoUQCWF5hWFg/JBI6bmyxBw8XCyAK+ciwJUz1gsYPrIDBCd0huyjeS9rujqZt
8XokhUpYimzGMgoc6gWMY46KF2qjgPpYnXa1X+zex5TrYbj/GREDH/8EVmsiqvDS
gGchn/7EDPXlxEfMl16P2eIpZQWd0oDmFtiRU20shmTHZSlb34BXMd9diP9vMD+p
958DfyVqvM5f7bI3MvihgPhYWPLnknlHg2eXgNzSx2f5pTNNlCylho1rSyaZLOv1
iMJb6QKoClmQBdQZvejeuOm225Z7wVnjHo9BwEZXaYqe9PIJ22dYJ6zlhWSKJ34m
nJCuJVSkO33t2ac7apOkaMIJYqCgO6NQMM5cskBsaFMJ6eGP6dlVVIsNEED41fph
mkiQ9Z9BhV/0BT1+qLuBJgMQu32QAyNBzXL4XuXpSbAIwQZ/Hgn0/yalx83ofdfd
FjTQPe9hXo0yaL4RdPqrimJ3thsguFHSIhKufsA/pMBGD4eDmQmY/xBNsmqm37ug
3pqY3dZ+8zXiFpNQQVjNALMngrThoWqFQvBHktAeh3RBqr7TG34K1o04+f7PiYTe
oplTFnuY5Ligw/f3xrZ1IsG3aUkzH+7Ckldqtt1KgM3ITEpbbOrhUXbbKqqVLQ6h
47P+y+nRzyfjmtRtP7U7iD/fqMQdkb2Wdmk8p8zcS8r37DiVAZujyaHqQBRyWjdE
gs/iuT6D5R/WTGqwNv06jGuzDMkgDaH+9M22GMXjNlSFsfkQicJ7YjYZ9ynxA47e
bKwBoV7IADz0asKxRtCPew6K9W/281s1bxSQQkhhEr/bQcMT7huuDl93ipUJxbIN
ZwYdzC4Y0uTe5/9pKbR3YgqE0M2g/wEAijquhEatOHHx98ROVMi+EIMZWKiDK0kG
5v4YPkydE4HU/wyp/B78ZiK2gf+dOjTOk1YSgz7275XJJ/orh6bXc+7TEGfb9ReT
oLWX78KHrh9Q0JPe8/WBUzx/X7WdoWzoP16CP4fxNihfpUIRh6+cjDObRIiLtiUj
N6N5TGi5WdAhGCUXjrfPxywo61wWPhtzzwmL5h1MTkxv5axq1a7hkmlZJrqmpsgJ
UukRweLKE/3JGPRS7SR8mXp+OnzmsDupPelER919gQoH8LH6amIgYnFOxR4yQoS7
H9XKKHpSJ79OFaa9Dsrb4Uj1KZbH+NdKkUD3sv1YCcih5GbC7YH+GbFCHwGARNCk
gPoFUxVpJA6UTttiQBoj4ZNfKssQ6+BRF4/avma8H5D20Ex04wEfjkiiD0JLmxJ8
RGuP9v6cy3Yr6K8QKEnIgF1MYy//WW/gaA1OlNSNFkOxU++hq4PtDezld43wNf/s
Qq0irUq6+POpEorO3Qtf370g6etPrCNiOgObL/Kc568hzYEd5pjUTUKcGDa0jytX
uJ5VA//7yzhjZNLKS6CEWyGi7axwY2nt4cnwmeb9T9xZ1OmuLGiB7zgurQqyjwAX
ErtAsT8O/sVExRKsgo548+psWMQ5lcmOScXPZFiZrc1jv6FAU5fRMO31ldWjjFF/
rl6wVTEwrq6cNZgTKtpP9wBtj1KYOBc/PKfAb5AzZN3tpuVaAwaZ+/3RFBWm8try
smuqKzm4doMBKos867y35aRLO2IlcPnpQAhDetw2ybJMcnMHs/0UlhhOFskBSENa
tyRwOshWQfNaWa1xu0QT3R+etyPoGFiiaYc2QETnjj7QkLqhmfiSI2PbUf5Ml1gT
eYNW6Qklo1P06IStRIu4ASC7XD1ZPnFTk/7yHVmwwitUnJlYKu0Jymf9T6OQM+6V
X/IWqth9GlYkacVVbA6PBdSBBeF5EP21bvO+dhZXGPVaKKrBfg7xLVb4KREtHZLZ
G6qtgkOr8uzr1FWMU9685IpBTMr62K7H+jN2lHXav+txEcMGIGgmjgjeln8g4mZR
FW2Y3p3bVjEOrx0WrvMwdm0LgDdd8K3Ek5rZwrUTZVyhYRwivT9ijsmRbhIUTmJL
gBVfmKOlExvJUuTlb7L+Gt5wJw3M0jiGFPgMAIeQ3LLvfKBoIiES+0fDscyBieQx
DFzjliGt1ZfZyKGudOW3jDA0VOyNxbHqRdJiRRMNXmHDsBVGmVK+yfq/PUfQ3DMa
XxzWUAzlU2EiV6EBrfera6qaQm47qdwUxL/CO0Rjc4OScU3hdwvNky9Tw2qwHsUA
ITi73cisW8/3QCGLPCQ2299x4rF9r4pr0ltGaFE4ZWMjamuAQmxpc1pdAR/67iwb
l4+x0zCjyTYOJyHjlsWEBMQwSSUqq59YFd/wTIGQDovnojSSWUDMrc1tpdX/ZdND
9uYmzcgsFdlI4RhjAmIvzyRNxY9FAapIAnmyOZhaqAO/DpjJbp34nlgvShZNnC9F
Ts2ulhY3HZz9GNSoD3NAodB7AC2M+fg/sbisBABR6qPRIyT/k3Bp8gCr+b6AKvRF
jejABQsvFrYeoOpwwB/XkmUHE2s8XU3GYznkKN3CKt2JwU1AYoZxZw/jrG7YAL5M
7RFAMmK22J6XC7CSyAw3qI5pvd2o12URdn9fonl9qOkXkFU9t/arZZm7UfyiVp5P
61RFKV5NWq6qSQkEknce1hjBF2P7vuBv1n3kp5AoZ5MMSkOyOq/1nmDHYpuvKITb
fMC650ICw9wCNx1/eaqH4B/PWXGHSAedanhhO+Zvxn+en2WAQWqNPp2GbIcYYj9z
zmz+MfdpTD6EUdEbCvRA1qkcJkeULEdAXyd847Y6S1cNLY64f20Je5ypZW81bUHJ
gDwkyAng6MAAnypDmuHM+Om6sV16CM0rnOVvV/8FBJGAAbcojRxhkqe7mmvOsyM2
xC61kbjPNXLsjre6u5v5T0F88QMsmUEZNiKlqLOWS/wZjhSpGBnFC7RIXL8Nn6/X
1wwSawJr5OYTbTIyuGhKLnQUF+doY1cfvhoCIoXe7yUO2TDkWow80Rb0SexY9jSl
68wVbhFobYl7r3spfuRF4FHZETL3tgg0OF8GYbBUXbCBKbOK0+irapAN68tDlZ7j
BU0cexKp43Bm1ezXzKsJnvsO9mO+Gwc0Mv0MZu5c/wSjAN6OKmmaqotlVw954sFE
4sNelHL4cN8ochV7GnPLF6lzMCDoz4QdEW8HPal9KKaARIha910tnvJjA3a6Kt6Y
GXUViPX7oGeFCx5hzCiGUHv508ZVAFRtmpaY17tstyM2v0OejHaCHmjutFltDBvs
hqS3LXXQuPSirnGzUdh3PgAFgnvqHibN4XwrGQIQe5pFBnoOsvO0E8qxEMrW1r1U
lp6nJ6reb4l244yQQLDLlIYS3fg2/LqFsz60WJltehK1jPlGa0GuO6x17EDqJA8A
/EyKH1qW/GkG5mV9eXNFLD45G/qglsCnXe65ZU+LW3JY8dDwEdXh9zt5xZ61tjmB
7MnptYsK2ybweqzfjIPbD1PGHOnEi7H0oaDPDJY6iuckYHPl41dV2irE3rRuMx3m
VQU1AyP9MT1Q19PZf/0CUBfS0629H6Od/T4YMHoxna/4DVszWbN3slTDX5ABIzWm
t61fAsELZzV7Fi3jTtfyjY5XiKZNEqQjOKb5FV5RBh8+cSEEKubtKhY1tu3XKZct
qfswN2gwC2j7o3g2QWDneoYb12lhGZkK+vulr84oENVnb6INyaI1b/MTokcOlZrr
Dcdfk/IkxymmHQQKuUvhuGzP776sp4YzZJXW8ft6kMXoZNLqrqjJt4x/3pw0fEII
h3w81T1dZ+uIkv7ezuEd3T1ocIoE3SnJZ/9kp9Y0NBuIv92zwKMZnOIwlkDTE0Up
2xAo4uAlhmmRGl3Hrow332LHw3D+4cZP0M1MteIhMf93PUbBs5kXwXy9XJLKrIB2
XH4URULg1L+sjblyjDn2rtuwUmnZbPLeGeBc/eg7n47jKb6pIWMhPOuHjLXRILLJ
yZYJshRzW9uDm9951Fu6EWflAIUVJ82yNAToSarxyJkuPQ5BTKfmb3T2I0B/d2Ck
VwXlLGksl9Njb/x5CodkDAxVVOGpXL9STUBhGTbQFvirY8+vklmLVdqX39GW9srw
AhjbEmuSMCexlw7Uju67TOSi5pjmq+QtcdvtR3iosWzgRsKark6sGZDvZtXLbjt4
uf3JNkJNzyahU0PAIhiweCPI/yI83q6cO4arEwrf1++WNkwlq69ZYB/XRYpdoadz
Gyv56pslkzn0+ZdMyh4foiQ6C89FoJXMOgQnouPggMx2/hf9VymP60qfOf6QhpAD
3izF/dTn4UAw7STg7sgUghJQNNanVMGDl0Nu0o5g47TGmiBY5erRwoiuZ7pQLeez
Z3z1Bv4RhOq63n1M745WBh0hK/7xRBSyzEqmY9mfbaeC+hk/sXz37n51YI20p3Ww
CO9oFukfPCA0KvvcaIcP0BPc/SuoXynfnPnnnJAOANtwB0KmuscADvZevuHiRvJQ
hYpZEYihcHcgve+Rjgb1IOuKM6w32uon/tS23dWDKinp57hmtTsVm9FLNTJYgAnT
NxnOpPP1Hubjvv3KxpoN5JXMatztoaGFlg1NXiZPwYJ+PnOpZI6RUE+4K0L77P/0
oWN7DAQEOKGFA/7BZwl2PRx01SoP0ajYyXYmyBgjQgmYRMCqd5RReCXasDRATfLZ
s9b87ngNycGcZ/Xr+9cKLR2zsFCNT9oAAw9b27No1Qa9rzRO8UPAbvKsd4drJZFY
OwOs1M/ZsVPuQUKGTJpxZO3s3TVhHE3hsm4yuWEEa5Xs9K4Q0X/Z/UT8KngTWwRo
V97YejzDbWn7EYOYz8X+LPgxQaZTnqtcSbCsr7ExwPzy0cLETLHecZhxO69nkGG8
pxnQ8vlDCQe91bm40D1KelJ3cjAjStpbMfa4NSpj8pvxExXgFqUhQ+cahsXISsNA
6R4eRgRXemp0xwUjUGpvkw0tbQ8BDV7fbj0GmzFxUcwsk5kdNRkJQMvb3AhEWE4y
wXHXZf4UxyL1XbV3YuKv+dIw19E3h+XEWQvPzxjnxc8IpM1LzgwfikzwaT8KaP6O
9eAz2y77sUX2NG87Oz+orbaorwuIJROx1NRbdK+LnYbVJfn5ufwLnhbQygLLkF5o
K+qJsL/kadobUj0yEedrHmFZcP0Ji1Cr768I4lmXhxvANYOLgk/is2UtM2czyfhj
+SRnmvCNhFu9V/ePinmcKatSI8D5Jw2L4CNHGMosGOC1kJXLK7npVQ6YjQRCAl90
PY0vhoVM7VLcnZgYQYqRpNHHRNdIhcFkdO03bqsw6y13/xNBJDV4BLr79pp5Fw0T
xQcW58dZOyJfk4sa1wwd5btwBwVaunf5sVan/T8Ntd9L4wOKnMcKEd9R7CwxD4BX
Sie6M1P3SxBySgNb+AF2Rmcak3pxZxVQxTeUnzIX9JJ7J+NdIf2undCcmtgddn9D
uQe9IztX71q5r7/4X/zVbwtovmEjEjpAizjZkqkrfGlz82rb52kXPbq3DWbHqcbf
gmDwjaUQmTksh56w/Awdt4uU2sUwUiDYPI7wqwyYb/gnCijRojKjCIjw1XqT6obP
kCqdHM12DoGcgoPqtky+exsp8aIR3/dgvqrJA/grKuKFasQtiWBXD5iREXYYeF16
5GX0ghedKIf+qBCxyMp2Ttq3dN8V9LsCFHdpd1Xvp3Exz859+nvyRSUK3wTy2C5I
dst2v/Ce3sjn2XSRm7uK9g9B3M7w96wGqZ05ZwlzuNQrJKTyAuxfiFpoWETWQKpV
Db4BtqBjvfA3Ux2UPIm44pp7/xsjusr9QN/yohulqD/R2dIGrHs4E8k0zC08JREK
InielYUXA7zYHI6oZLNeYsD7uf8Bkjgzw4vr7YgoINga2kEDkAb/Mzw8iLLaHZkG
xwbEScAjO0vW4in9WzfJjw71BY1kvzLotUTBK6OLTIxYE2k3WPnCXsb4EoN6nxZm
AHIgGNtBHqWird0tFuYCrEcJmRkM+P7UzLzrTCnWTaHriWMRiBy6VDdshL/zHD9t
0cPm5RtxYV0MLUa82BGYx8eiTjnJWXJFgKobUc/qfUTUY9Y/07gKep1nGY7WoMGC
v5z9Bp9Vrv3tK/yaKrJtCqJ3vf7foCILCmlhFKX0n06il5vnOo0iPO4l+ozkeKp8
+I7HRH8MjPArpcStK/7EGjFOagYHrMLkF6T1RWuc7F2R9Qwqzmnn4KZuMmKRVcbn
Gk5bj6gZkVjhDM3bLFEG27OlKxVWimRVmysePaIA2egVdIcck5v/xALeDj6VQFYb
ayQe8JLRTbru81IEWX7x6mpHc3mrWG9Wu+7AS4RpMrI1ubFrw4JM5zat/BVzhJHL
oPq50kKTu/41ax8ZI70EwNyRMol8olL2GbAFVWx8HpzQNMUYb+pwadSgWGy+WYWO
JC6a8RnXHEiR4wl+JewP9/8H1Dr9PkFgMnGN1/dRY8CMTrXt5amOJhMaZrWRxoCx
/rBZkBwnMop9Gkaaq21wEiLFjeagyW/iOtxWi3yT79UvXD69wts5GBm+sl99mVX7
lDFSbnZ5AIduAWu/zFRqegX8522lHiBrgg5CGwy6H9Uv4mm2xLsWBzJaj2LjRw2h
ufw/+HvUpL+Dp0xvJOc7TBOJQzuzZNnVpnRKwlvEGPQM+cMCAkz68TNiSgAWqLum
nEbo21dBCLP+mUytLg2l9ZHTZcAS3hGmCihOGdGJNLbP1FC7HW2Y5uYfw7oEPFYY
BtLtWHJ0YDXAuGp6ZGO+YKzOQWz7wgQkTWGlR/onZVKL6eFPWPQj+QIDQeCYp6wK
TDdg9ZG0qUARVtP3Stn7YBHlxSYpohGTePndkuvg4d2objgHJhhuGH6uADURdbAe
2qsNzTEMaexjXQgtHJG5dFEoHb25v2VdFOfVEmSPnwBacVAma6IxDfxhhbLvKCM3
5Txcz3HJZzECXgz9cnYz+NR5yo3gwnjCI7lE1aH12CuHCqpO9iEAo5wburpPb6aE
r5iUB3+QhYF94h0Ht+79mKi8XQwgY5WfjN+k2zcSc6lM2MFW2FC06iKpk8rwUUbT
XXOs5UUHJaa9K0kAyZOGIBB2YhdhwivxTdNxJmRpK7XWgzcMScnF3wyQwUDT+SWh
mApI0Z0NDCHSrEkEpZgCVgCRsZWYSZlcg7tYM0wc4NWxZVsRdrhLssNLf8g58WjU
qOOTcndMAW7hYddE6pVx6jyiXls/axEDlKZ7FuFW35D5S1kaOR4UjyoDRzh/Yvnw
8wBqiU5UZccObK8WrOFzu8qoWYncsJ0/DbhA65tVhXK14WaJdchQbI1jkVSxeYIg
PuRQTLOf+J2uPUHSazntg1WTggqSNj1wEzncSDdG5sbUI0M+SA26R+4UTRiAVccr
XTKD3HMRQKUNeuSQkfQ8dA5UIQbLc/3gNu3yj5iKMXwuFUe0nfoojUmobTXYTH63
Wp+wKpkTfaKVcXHN6YGWdE2/qhjw/C3fLDJcGEqVduqtci0qeE8fHJmFOkh8huy5
RKWfZbv5/xkNg6iaVUBEI1hOHxCIL4GvfmZDw94OWJel8khIR/zllwByGaeyxU1j
YCVrlbsF/EI67GJ3aBjxkvE5esohhSV7JQBNjJT/p2FBSqQh6vFePlXTm1H4jks2
U0Vcw9EE/YSB/Sa92eAXEis9g7ochhZ5IhV6PvsG024F8VJZAKBxIC2YGDBD16Gv
we1QGq33hS30YYh+lUINfBbuQPxA8YiwiXU35ASxoEWhWHClrfmQE6//NKQgWNcj
KNTD65D0MbutaxbAVgiWiuhIixChNxwlZ74uea/ANuOPtK9vR8rKCrhvB+YQugh1
ksO0UY7X9UYi3AIb2N65e7z3nYtTZdt3gkwJ/wwdB3UB//HFq9vh1SBTWserv7GJ
SrGdnTGOsu4/NUBArmNMpowtgkyLjgQYtf2QMudywaPRvRcC/LmOCb/yHspoCM0/
8o6eesOESu+MMUEl0wIUvDAunT9ysZ5EkxGFXAKPcIjLppSYy0J2EQ6kfz1U6/YM
3nOWuRFvoyvXSgz8jsjHGB1LX2SaCgltEBVRyvkDhXtzx8s/BzIbwujU1w4ht6QX
VSF6sHMHvn2yi7SCkR73ZKRxfZ3EPr4/WyI1f6m40o6JXZCf9/XIxqVl92Ra9hRS
rtA6hCBpF76r+rtz2plHn4IFNgiUgRV/TSiBS+AIZHuowB9E04fiRHkZE14DYoET
OnKqICCfWfN2R4RvxYEr7kJvZIbuTmnN+EceuqsasRRKY/iWXhnC5++HMnHpn0kc
E3hveYNVVdCPeqBhuvk/VXDuN12ijL6Q1m/yCsk0I5WVmX6agb5XrHA2WVtPYjt1
mEtIkU22SCwexdg9KR7i4YL2IpjLoPDqEPBmWgX9plKcFskWtKP5SNs3rWTGLhQv
dIAzPSmy+YwygAgC+kzGh7BRtvGkxxO3CLl0jCJlOzE2ILNwrGwyDUdd+E68iin3
bRzx9KTLp4r6Ih1ZRLa/Ule3DQ3qrRpBOVvbf2IzdkJD7wUikaYFINHPOjcCitqp
vaubNy2wTfxvu4brxNLasE/EZpnSI9RkezUnmlHkRCL9zKFjpFRKEfI0nCWxs5ZO
V9O28vFb41W+w0E7NFBsB8SAUeDJeQRITHHkjLIlW8MCYj4yJkKBpL4ZD7zEcdqp
WU2yS1xoid7k7ksqaUzk/f7Luloovumo/PVJy2RUv+1ZHRRrK+h8WWnAFf1NLPwX
EktF0h1BSRlmyuMfx8Ho8TJMbMXRkn+n8Tbyjcnu035CwLzYoULIAKO1Fsyd57us
U1voH1IJmo4YSNnejoIrMU93eI6kCMmUNhWDCtYfuSrBk6bmYIwrJS9ZOglf39/X
HAZa+u0DSG3Dxzp8KexC9bXlWVst8S/+tMii2HqdW9mH04MYTO+RrVn7NntgiSMx
4YcU4fh97y28GXX4oNoRYWY2CDHS4J2ls5xfv56Qm/Q9ycYXhuMah65z+QVCxmsq
KmXVBMtuUrK5UOKt+7Ey7ayUFHdGsnBFbBYBxs/0JtEyNurwxJuAQT8IKhTmu/86
PvsMePa3SXw/aoAKESDkhbJ1m2osqpyf4VnNqvWib8PWQal6HOHcKvdo+YTCKT2Q
zikdTqet8LgTsbIybKf5Gs0KDdb5XnW0SKnxjvOtMx3Ip3BAonLuYcMDygqPOEHB
osDy2eAjBsPBb2/Eztvmgd0SNJWdzbI6eqwjiM8QcEcHsJA+Vi/R0M6YjAWYsPex
yCW4JEEP+J5XcoAdEurw2DjBAJU7X8Y/yTBCiRUI73AYo5Ub47CV5+wXfzYaSfND
hao88rkoeJwJJZbavQxrXG811zm4p6zVRGdnjY6HFO82K1+b6Jvm9k3zZYnw8ZYz
v2f9NgxQfvNaaKty7eTZZ2YULBTp7Pb6KrmNWK8d74uXxuKhocW7wkqr80c/uXgo
BuNVa7pwJUJlXTgXsv0olNFCHiX2lxNor5IHlLXRQJRYQXvP/gvjzStrI1Wkeg3x
prAqDLoES0F/Qb/kDPNUTLARolNNqxP58wUhcpFIdehis1IG91FPHNCer9XP/giD
1gSoVVr1KrG+wC+VJ9ushFsC0+a9ba3shlfHPNrY58LCjsSOLlzp/M/XVPZN60he
ZpmpIZVdauP7sDpYRyPHrRgpXjytQJKXtP6y/ovHpYaFIXhJVK6w+VOrT5vORrEF
VNIz1DwjhbMyPYkTm3wLnxwfzwiwsEKuv8TU4dhS4ksGohNWHxDROd8QGPf4sERn
YklfGNIaoICKh9iWCY3bcwKNG+REZAArHoRstTM4Y7uhTTDSjdQ5G0kPUyJvHmeB
XGqIMahp4sbLhbPiEJvdPC8O8i2FZ8T/lzjyqwPfEXh5fgWWcK+PP0yI+IsTHRUB
zfd6+sAfYT1BOMzh84qp5yxGq0AUvE3Mehslo7q+yUud4ueE5acUBTc9FNFb3nH0
pAsB/24a4Po3qckJNQELEYJgRkuoXsfrEX2c0N/xJHf2Qn9ZE0EAeRVLt5vrcr/c
scrBJWu+79Q0mErn5QXWWfz211r6kvUIJy2x6VAQAKzJ5/F4tTea/PWyevUlRDPX
tmlgfUtYaV5E9G3Lg41zrW6/Q8y2e+m9IJIuSZw8PGYLkf5jwlSmGA25mUDLBcBb
6U4rZVsRvhHA81M7qJ/8WiUXM4DsLqWfkFK+8lzdOF8qoXNp1hjKSPyTd8xNb3h+
86XFWM3VirU9YappZUWPzWKlc9/sGSpm7MqHg936cF2uAvL0LD2yMNVXFm1K6otR
bFKdEsVVxjlbyfsLAwCfOhe4ZXQ2TbKcNtwrUKUy/vnmD0dza+HpoyMrEtxbpGfJ
hB66+NK1jxDttzlClp4UHW5h0ZbNgF0GKc3AdrcHWm0pvq7gmZfcUpi4+neiuUSo
LCtmIhYfZ6TMjG128HuYclVCmB6qHNcTTBpGk5eStT7UuCTvZ8ur3elnhk1d3PwP
IALkyHQbMHCK9dAhuuQ2EPj2wSaW0ajkkf3TsnR0VOPtgzjmZYIppRmmEef//IHd
LGS5TitiffTBOL/xgh2cXN2hdy3+TUh1jLIXOwnANCIwTs5+/5UpCT+f2MxDOuJI
xNvYkTQbbu4FyT2du+fXVORem4WadItIlUjv5310PUzjzTuJ8AXj5NzL+xkbK7rz
1+6RLIWOk47zNIGIPzYwFvCDKzUah13CQA/GeW2QB7or9SQujzXhmO/sPcTCemi2
QFq7/33tye98mdKmTDkK0ujI53cSrwHPBoqXpHIzbNOHj1jVcVoCOz62IpqAX1/G
cRnoSBuMWO7eOYwwE6MUrU8GnC2G2fYbxyPKMGKnKu+ptkAzrWzzT7vhTLs/zoT2
3yL8gVgjfQ1hY+fJX/V4p82HXJHbWyzUVAL+7JbukSdCDKl69XKEIUnEPsQ8OvsH
2sWrDEu49oysN8NpjAgYsV3IIA2raeiUvx6D9AhkQjoeAmjHZXXnIOeSps0LSiIW
zP1EVAuy6YNiUnVtXtfOg82Q34OSPxHfZGh4609eDpBO81ZAr2uYstMyJHAArrKr
vr1OAqIWRjyFQYVNDrzqrx/WaSu7/9GNlPCSBiscr6j+g+kGuEXjzP3CgwtqcrbR
6E9W2EFF/gwk5/c6j17/uu3V7VTT50O8tw/FRwtPn58lpL0xrrXebpUpZOdYAUft
P7Qg2+m3fnQ9FiR3TNIRse9DP7r9R7+ph98r0FAkf+PuTEhrTZarXEoLcXVBmy8S
s5ImR/FwXEMvzuVYtKphFsbkkYLgA7H0Am5UKul+G3Ln1/GtVyRdKFmimUN11Z7j
+3mcP/Jh+V4GHdb6//vNjHtt81Hll81HD4DrIxg2/bYnbyG0aYs6DsSqrvP4lS9x
2jgetH1Veg6fththuzT5qmCZ8Hf0NT1R8ZLyhkMiUDVBnXHNdUc4cyLM1bXQNg/e
HAXdRdZiU85cz7Gcb/v2wLt8gPoISPOnW4OtT5Oo6a7XgaLWULasfuuMxeHLaKZQ
aVO+2pNd6+cXFISjJqMWUrYS+pGfntghY5/PVd2SQR49hbkFuVTQPaehWDkvJ8+s
wJaFzxmzoYcCV5DQxAIDpHn7BdG6lx5M/WrvugKdUO/LmL3BZN+H5OAgndZy3TIR
F3UYCDyKmsJeUH+YDPTIZDFuE4uMTFl/KLEMhJDrLQs66CJVpD8BTJGm23uc+lo6
OLVds/83H9ZI2PfJIlyEmperT/JwqwIEesMCnGilGOuIr2T/p2LbgF5Ped37QFVi
bmyoJNLRtnTCIxjWpRm2f/8d4Gj3WCMrB5Rwijd/HKUoSIRIkuQrUsPqhtUwsAl7
wFFYeNNYd1PanJYv+rDs3hPyxsEzkeuCuJtRX8e3fAy9MOybCxgP68OsFKRV/1Q3
6BuGgMOd+ovfAek3uGNsdkrQZrYi8QGszHamxWnLCA7UTMn0piHkS6GtoVsW/pkb
xPqHUChr6YjuD+eTPjqD0CeLHBcgM51S7R3+DzjNaH9GMvQBOkeBJ4L+zsMjLQ1C
Biu4zwH1+19IgueUmRDVSCDCgS+xOsZHjCF/ftEig/4PKIHIjk/QYcS81e7B0eut
kmHUZt38wAvCokJj8BGI32cFcTskGNYbVsITiSlnw1uWxY5MB2LY8zHuRWjBjefm
T9igtYH4XNgechtUdkkNLOxyHPrL45FS5wpy61Ekrh3wXh1NuUSZ6NFmC3eEX0Fd
fAnYvIEfKjT2PEC0282c1STWV4nEmwfCJZQBTntobMIELLLxWYhMOZgCTggbMz1N
goWerxdBMAyi4J2h8iWJkctYfUVIVHoGKDKU2ZmNuM7eClfe5S79VxEPuVq/cs0R
jAPMHAbcGY0WTXKEkRU+wYpHUuZvfqUlvDtYKPCpA5pHqAFkBlFIf0u5dUV2qrOi
CfYlAiXvKC8QwB2HgtCJWZ845W6+vDcGigCjESRHsgfQlpncJsWjuV+h2kiGe3uD
p7Y8n/kPHvIV+rf5ilH5+rpUGKTXjPboWa9Ed4dckeI+xaknX2MScvwfzE1Gk3p4
e0KR1+wHhTheTLlDWwaYzGOO9l7dhLFB6NVk9xPXSq++Wc4bYWNHnGXMvfeGpSjC
FKwCjmR/1tVP1S7cqFCUCaPJU0ECkNWN2muUKHp8z25ogvnYcstG9mn3Wh8AcXpi
FdRX/uYEtWD4KxM9zsX8NIpg5UycaImPDHoIsBWeeSVTvtEzxQB4xfueMYN5BYmP
o0JIwlAgMHUggkkEHBkussM7/zR89vLPAqCvNvRR7qCIHUK+ehwUjOPOPEFNGrJ3
F0l8YU/Y2m6rPGaStbIZX9iti8UK9/5zMvkvc5VNKpb5EebxoyDq7DeaVQbX9WVp
6jPIUOnyVfIYC1VIMtUL+FND/EKfDjlt1CR7vt+4Wg1ZP/04EvatN9M4vzvcSmfy
vIbFSSbtYHDswU0dmREOxDewdtpTrjI3JJ9jEpsWPcd8rAJDmndQVZpjQh5R7G6X
KWIF+QdwbP6ITSp4IGY05pgQLmI8KkytOc4Ad0rrXv5zB1wBIwRd5iW8LjD3cWNP
uW/djsumh3Pow5rWSr9VuJnKliin0V2NNkS3q8lTy8FPOjVwwXbwkIL6KaQkG4hH
8zRIsSZBmOTjEdz/ND9NBNiZpaONgkadrI6Z7oy5UZ/z6YbcMn4efrdjG0dED9FM
F1mgPwUMSa7R0nQY2go9WsyRRJNCx3tG+pJkDT2eoJGvR7UpR3nc14p9tiroU7Bd
4ltGTSUPrIOGIAHQoD2eDjutRo0PYcvzFuMRASDKH+vbp1ciG/GgGO4CEVH9zhcI
C8idNHFQxbxkTQkVM/nOk3HTtHbd/kZ4ebx0uelJMG7UE2PP7jjxHCkiKkLXG1nk
iKujHywtIcskhrq2yeBpk5AYsLHKVTaU++wJIpCofL+pOXlczkQL0ug9Qsadvc7p
uOND5IKObWvQvqR9BUGKhgpQNVgvQuPM7FnRs/IIs02ah9dW6p76IFTUH0ZX4k++
2gcu2F/28eoxc8WIggqv5aQeJ2doDiFzeKKf2gJQ98iqSCuv31/SXRyFXRoKTBoJ
N9IFwzDZVdkIKc/9pYCN8Qcg1Y3Yc3h9T+E84sw5S4KWSzfwC90GDrorS4dtRQKe
0l+Omm5hz3ZOgGsImm0Lug8evSxDJuyVw2NGAiF/X9O4Ss6m1WNTa889rbU9eH6n
ly9wFD7L4rwv4EwqgZr/39E7g1hhcKn5Kx5mr+cnWnS+MhkmenFZAXZ7cog/pKw4
c4ZRT+OoUDIJ7UGu5s14fOFHct3ZOgg5wu7P738BC3cXms3OgbgKAjuEdN/JFoO0
LNQDi6sV1Fbh4JMp7S33IKFIGQmkoenNHW8jmaaSnizBe3pSBXFbVCak0+1RoyvI
HSWX5IGkzTLuiTMV4lTMB+2bX4wuWz1dOG7W167NPVc6I4/HybryySDmu/6OlMKo
INwlkDrXtzJtVHj+NGaV5C9ro0sHn93lrnLgLwzw15SRBMcstAlypWV+A5WPC7uQ
daGtr3TWb/bqVPiA3YlPvpwaJzJwezC/aPkb2gQVzvbrQvomQC8keYeHa+yRXsyW
kT7YXxsgANmbLs/EGxuzwQ5QlhSIws7ZDSV0vBUsyyljYgrN/iHXlknOSIutH0Gi
A/hxQPWLf1/8j4qKwU+vYR2sqZoo4O5HLjWFXr5770MxkKyNMnki0oeogcELcJm0
2tdcEKOtgGFeHDzBBrN7aLrwcIf1vsv0QQG/hV+QNqEaiQ38r39TL4llLSy3tF1t
IHRxVTM2VZ/gLeYDuWEZ1dHZsJTMcKP2LvdgmYDxKARuUezsZHFy2qlIeBgH69qx
gilcnpKnbInLjcHtE/pyddb5U32GcXeZCDu6BgE9yso01dmsqjR3qKbAnTerO3KL
+2/OZVVq7rs8b31CygXIYUNGImxmPG6ZDAOw708+COVzrWNYdFkAXZBp0+iKCr1Z
nYRMhk3m46u7AUhqozQCTR+NellAT3TqDoVqMx0Hl0cL8TgBhHPCngN2kkyEcX1f
by5aJm4ENP3T97iA8yHQtpF824QYU2lnDljC/ncTpu5HyaF0HHfSz0uiqVgOcFEE
B2RfD5VxdzixcbSz/QEd+2Cn4+kvXahjnbPixMkE/ixf1YhdNxqPdhDPzPQBN42U
emetW+LuHVf0Lj/djUCVbqQAgfr2DVNbgnTmNz1YFQbQbWJCy2eKJEun51oyGWq7
xUrcSBKsvdfXDO0ISggNG+e0FzTPQxx18rhy1Y8PNLzZwEFJSfsYruPBatpoWffG
Z0z6xMEFkCXKjTqs/MPBh0TK9kCvDtokbW/pxYq/+aGVDO28GQOxgtZA1mOnpgdW
ebaaXHyjiIz0mMWHDs3DEyT3zY46YswU41iKsrsO5s+pbAi2aSLe9xBD3H2NSiqx
hGUkaVPU5G8otz3xiyWMr9PqfIVcWX6toe6DroxyskcwIigEhHdsgd90HabHvBbj
e+L5x5hTC5jFkY1yij9HXq7dU6JIqStK/ve51QJ0vVOJ48Sz2dolEC8xvG1FVTjK
KoXjLnPH1jlhHlYhOlzB5i81FkwCzpEtRA+Z0iqJP2u2qlR9KsxAAcfHKuFc9Wys
MsSBPbmZTDYAd6WdTQpwhgne08e4Y1Yv1f80NdGSJSniQXDepW7wlpI+feCR/sjR
cHhqDk61QXEL9g/Jg+j4FVRrRtFDqGwQUjskJ/aZMdRrfODjJsEsgDcL+0b4D4U7
shXY0f8wt4NQjvF/mjPJmDm1QpMY0utaLWaLQTyuQKHkRyRjuITNYvo1/+hKw+gW
XKyWZClKk3tD7O3w/kUTHEumPUE19KRkf67CeOmEOggjd3nIdBwEZ7TjYNBLMvlG
Rlc6RtvdN8ZFahd/yjwD5jXHXlufk3ddn466M62bNazaJefiuB+g8r3ivYcccoHC
5jJ3jvafwWsa2W8UhpNFvpUP+3lJKXfH6lbkj/FU+y+WXXu3iUvsacWoYj59d/nR
i4ifIsCkivUBRzNvHJHSYqFHEBerK2FQbr+P9nXI/EiBkwlfp0OHZAiImhj40CCC
1L6WvyiYJUEz1vCrQDGbo9i9kMXrPGJJZZWFcJnCjnXG3Yrxq0APxewBHKLWp4GE
byNLL2qth6RhCe38qLuspNPO3Uk/cB4BD//Q93ZZGzFGz3Eap5D3Mn6csbZyxwMC
zfm7zs8Y7Udl0t3GUx+w/QBo8Mns1lqWZJ1cfzROYaBSVdgc5L9D5OGlUvv0aHTy
GFGXaPvKC3xtHeT8yTWPzZBxL6+HCTMUumDO713A1aRuhOoc00w8pp4lOSc71KJS
3WdRkfyo91v9uvA+Gm0ThwcsfFBTcd//DbjEvaaxCfpaBgBoPePQKux58UDoEP5I
CWvA/pzokAmw8xyxn/UlX436Pn4xD+5bH9/mS+DO+NHt2MqrvihMX8rBoQAKkEvD
ZcK3L0cn7RhSGQOlAAX9tzdBuo/R0KE/Vk7OcFlGTT/LwO6CQ7tITP61jgs7hTKE
gZdG/8aYFFi6YbtpTZJVdoqTADIwH0HtEmlgWmVrkjmWk5kWLcF6KaBqZlSGryab
9ZQktDmrtD9Z/D7jGGPsxhfnQPF5dxrLeWAYcfFieFkUcRow1nOMf8TCKw99i0H5
PsOhAuK48Y/ddWjujPxBa0O2W6bKasle9tdDDJkB3tRPz3l7F9numFuBSq5FFEWv
32N4nMud67NuVIhQlUxxBUi87Zj2ZabDCxE+14sBP44Ho2lW2EPv2cbnwWg1yrzd
b2Hed2ePZO3hYnCxcwrqtLqk3oQ0OTor8M8G2r/WDvttHWuwiBvMZqx8fdVdrR+f
SxWDJaJIYp9wvoAtGrgjdErXgOaaK+NVf86oFf7fGWVTl7dOF2YoDiYh09oBMzTA
Nu7Ybj4xQV1KfIzzNPb5tw5QB/9+gIexDj1npiJhZgqaz90BhoDSaQ2hgN7MSDor
rkwswwon7cvLoBuGgyVUxw1fogPcsghibK3l3CCQ+EBxEt25/BPRyPZQAzL14V2H
OtDZJZWgUm4OasZQ47TcLpLFEe0jFoAqNsrlGPbR8yYORz49xGWOIWMQcfm+18SJ
OjI0yCup+5xw+TVEKvAOqi2hjHXII4JaUy+UKagrO7JoMEwj6j8KsoIWOS6w6nkG
wPHBwoJsZN4EGUGVSV05K2RHGET5IanZai0tcifQwnRb5CDrwEFUcNuc8R6Sybmi
Xbd+PAnVhA29ds3jlB+LIF9ZZ1u66GnWJ+Cv5CCNYygd4yJ0TBPU3dGpBzKoAkhW
PLaBZWsiC3lF+AudHV7HZwFffM8owFtRdPWsuor4bY1ILMj+le47JqEVVRhsWsqO
hbkaOxHxLXzSpxqBQZ42e9Mx7EQzb3eN0IcfDUXwFHxBHZIQ3QYKt0ARqOJkopN/
L0+pfQZ4KfSC1Quhm8CRY5hhxKCDkHPe6YpV9oXa4wT5hBoeDejIz+PA8kk8QZAx
x6AfIxp6y5Jd+QXHY1XtdAlKoWX9BYOsVwLA/cqjGmJ0QkSdIs0peDfl0y/YwVeI
ZDA0VI6JFN+8E5wvGZtRSYrSwqBVOLRRKSjKpF0TLLOCfO9/LpmLi5nHXPtduMMd
T7Va9nmoQJsI+tleOwvA188nzwiHY8Mk192GC6T0QXi9vnR4yt7KQXmQQm3RVb9o
MbNVgGBHD1vOSH9J5x5XpuhuWVUhSvPaaLZBRnqPb2gYkEanhwDYhvhAbRAXl1NR
hyjMs4jWDLtWVfJ0tW/euCzLV+UglnnEXWmvzHkZiu2pHPULhTV866f67nt/RJ6v
MFAcZkB8W83hQdbpR0j8/kkQuW2UR6HiWAmykXLqpdWKxwE273VqqQS1usvywMH4
E5RGhkQY3Y/QjtIn/3wHBPzd890aozYJfmiQpKi6YPBNzWYCIieV4PJm1khLRvfG
3BdvStDorHjoccr816KsOIw2SK0g09cAbZQMoF8NVD+cVwER+RJgsH7L8Yoeh/Yn
bb9lGaQUM8pPtIV6ZQZgwxF927ZCRceqNGNty2kLaSo5wAM+ekdgDfpNLTuIw1Cu
YjksJ07kPT2dCc+TeC6RK6iF9ktGb2YkEySU/Ovah2TRYt3X9Lz95BtViP7OKCDS
DJFv6HpWgjCpyaxYaKdaqf48LOh8Hu1XoRa8OZHTF8rbK6pFt71oKBumGCaD8lLa
zkw1T07x+XFZA/Qw17zAvgoSX2+rcbTqvT36mICGEsA200qd1Bl6mDwtmeNvgsFd
MEDBUA9qmytzDWi7G2ZOO47i3kfxIET5DRzjMwGej4sot/ZWO4aZQoeYDHVkrl5e
CdacO6uO7aaRMJWnmZHYzPYXl2Gu8nUnfKYk82qym+WkGoPncmgYuXDCqUSYQoqj
FHbMH7NurTv7hqTXoB2v8L8XwIZwJDM+XmcQl8CnMircRsdhuNvO8Ll9mlAw/RSB
hRrSOREehgLUhLq+tzJbi7MIwk7RXYsSkTOrH97GKUdaIp6Lc3sgAOoeTGcBoZPj
ldkFcjvdpuu6Ij4TURGJ1dNPGkkSw83FZval9T+U5EmPbcvn3bWEXewL19F1CAtu
8ELYjihPEMV4yLVEelcWsgGce/tp6F/rtTU218OWUlc6KUlVU3PM6BLO9crh2pE4
XCAjVc/Cq+0TWyKF0nkj492BYJ1xF8X5pYl+uUaADWFpwZztRf58/ZBClaEw8uN+
qUb4Ayik36GPe/63DyzGaI1zMmsLHbJUab9Ru3VQN+ugepdJX4lZuKTaCbqjeoam
NhH4YpYe1zGJ2O85lgBmdsrRwd0g+ddfJYStlZ6Ry5r60BOG+PqMILENbMmJwY5I
zKfC5reisKfj0Cyes8VzIzX4aGmUK+0adA4kqjQMTq6OSH4OxC+QDQykw/K1icbk
Oe39/uX3nhEdMI5S3nbD5ae8FN+Lh/7mBHHkpNjs/u/v4BeYmEJq8XkNIxNubmzP
KBPhklJkpZswVF1rtaq/ZwX+yfGPKfG6ZLm1n7TxWyLa+0sO3aZy/QXflgnSegtQ
ylid7ypuZV8SBJZuBotWfH1+DA5F4RRZGlt8U18mUcpPTBedE7HlyyF+LLhXCL9l
ogbsDj2Q+gDvOgdnn+7f0mT0339030uCN5FJ1O0DH1JJ6QTXqRe+6xW3Hb5AmkDm
fPHBWnYmjjHpYH7+2qYkLdcUGgQ8Ty6GIw6skiUjsSLDo0je4ZfVixtVzuetwrYP
k95aMnALoWmNc5ldqP69mU7hUNTTjGm8Jduf0cf7q2w3p7pCSSMIXxhX9u+7EJQP
+bEkoeuLYnaISIh4anl9D09XlN5tfiKjq8jWxYls0UNGPAWsjqFMFub5R0Ki1/BG
G3dqu68Y0ZPojSVWCXbDoQYNIe/VEXMkOMKIh/tzsIlnMcK81eOK0kd8bBtj0x2Z
n/eq3+qp0j4/+s7iZ0D0Y3/e+w43TeFqplEb6njV929+7hfRvUi7M2ODbyy96z8u
we3ifQNUrmr/bdNtLMMZRQvIRfIoMYmRvNF+UpwiQkhZbVYPdG66HcSsKrFkm7OW
QPH06Y3GJ9JHwrDhpgWKqRnmIKvulNdcxmaH0V3Z0sL84nwOT48eUlIQbbKipwE1
hXjHJWhz93YEM7GQFTckyUvXn0ttck9QNLaZPDNML04Lzyh2JFnypui0s8sTXNSw
kRH2Ar0c0a3vHlBLCvOqw1/1oVLdDon7kgx0ZoyL9vQJhVynDJjEJvsHLmdYX8ep
87F4nGW4UKE+rPskqfvIRLqWhhnNTscTC5W9Gj9UQ6K/uxZYD/fE9/wWUub/somY
IcYOcSOStHYHE6uvh4CJOH+OtUA2wDc+pZmKdUBeOEfzjSbX+CEyMJlYndI3nNoI
0RxFGt3AoUEVP+loE6XcM315o2Ft7HVyaPJ5fwCRUVVQ5uqAssE77iMTXo5D/Qoz
3Dbc5Y9XgC1a7GH4y4KIRELZYVXSRyVxPem33azGds8q5nJmLF6+0D30ff951Z5A
4ZgCikzdB+hmrEw33IesvIZnOXWsmojoT73hKqw7/qAE71fwjMBnvl1oz/0JMEbn
9IWZi2l0ldtcivDT5zYM4pJoxoOxohr7jOh9Q+UrfvfB82NQCc/lC9LilGYiAP5f
tXnAlmaZpdaj+2vq3dbwdWer815Zkrmjuq54x5V/tFkLJ0J4WRcoJRoEQwfZr5F3
p4YiS3jWhkzAk4baOsAQtMe0lyfJgIMKCUQ0N1PtYX9LnDWnzNUHwGcOaiB5Ka+9
pDltv0r5m/Dt8ziMLim1Y/aRafeunqw6cYk/xtOzCSmc7YXX+nPD+EOiGIuB4JPm
oGCwC6smF8AZFB7Y3CEnxBaZwg52p8ZWyKgEefiDx+lMVfUr8qTOO0aZkE0dlNWC
SP266d5/1KApGXGaoC74VedbC4JAz/wpsFPszvfOyyHLhzHP3K+G3yiPc7V1f4pq
PY82rABoZLtu4UntTR9VNSZ5qhwADflZt9RVAk4iqQzjgYVLCccDC3ytsZho/2Bm
+2CY8dr7o6Fphgscw5C4fo3+qKFkjh0oFweBWXS24E14VbsuBytDTpe6M9SG5k8A
Fy03FxtgLqXcxUBnzjS7OhEPVlVFeX59WmpGDGUpOOoXUf+fk81YYJf8PciYZ1fM
jTW0MVom+X9tRe1H8MMmWuOkcwlEHBw/zCjKcEPT8fpklWFT+Z1zbPplephhm5yy
zpa9/cGejeKFUT1HVze26+K9KcZgEyKBRssmx6DvpqDYTdxleprN2v2LKkEmfFB1
h4PjEVL475CgupjOfgk95b3cq3kTmt5w6SoO//cYUYqb1W1O3HNSob7p+fEZ2k+E
1jt2zLI1l+M7mTVy6y/vyipQiWwVNNEBNF92iMSYvzXOjjFyOYc+AIBkREFBsrSh
Sg+du09ngox75HMhIRs5e59zbJd1MNFO5EXg5rermj/vGTiXsK9mOTFxBgPCihpu
lm+Jyzt1K0DFsLvrR+HUUFV1uo58xf8ZPP8x2JCc9TCdtlnQ645nsQ9hXXMur6v6
WFxulOmfTRiP5QKsPYdSwj3oQybL30plTpJdB15oiG2ivSp9yHnV5g8ZASoJzZbz
9C6CFLCygu2q+TPUgB1uWU5QwTBD5RBcSi4Dth7Nw7qYzfZ1sTmG+MuffTbeeXOk
pJ6YCxBNbN1o6iKIQmo/6iP3qWn5rslejmMtctqG1KsYYPAuIx5rNRz+nkoypIsz
ZbEJSDu9Yr2fTFbE6zRM48cnfE9YNDnslT2FFxO3mcvftxPgmzHNrC5yuiDkfmEX
Z12/KFlkUak3xsifE6ElyppjqklKpv+gDm9gKLtYQZOkwWHsVCy9DN/k0pBV/wcN
lVppKCqSbvzuAIbN2+NCIwKvxrSZl2/vZeqNVDgc5WlghBCsotJv3AptihuFftcm
cy79Mr16o/05d42W9Ow6bJJJ6l2Vxew3bxIzgEholT3In+cr+ZNLyy9vRs9VwRGh
lh6ZxRDKSrf7LhoHH7eBkInc8qJ6kho6sEJL+aFoscZaV+/AiUxPSYsWnvzPYpSb
OTUH3Ts37HuGpVP6Y9Ss7vSEXMGh3xWdViek83H0VQxTtwqHP7QaHrAiAInxHiEi
b4cEF96ypo8+CFS3i4HP+pk8nbwSrT9cfRJYvw/SrV2wOJTVD2dCGSgldvPct+jj
HZtoAxTHo/c7EtzgWcnTFRt/VX1DISysSjDEJWZShozUc7VO5mw66MNrKh684xxK
ohWdAElu0mElC7t8qCSoc4IpKMKD4LPr9RZTMCyOH77PLd4hw8JCWZ/R6QDEtQch
GLHQp9tbRfuobrDZqdekVsN0GGm0shK0+HEuB1HihCfVo7RCjys1qmDSwC7DYXeh
UT5kJfiOxBAD4rSWfL9Rf8Arap6PhFTAfkp5/EgVtNBwCn9kQ6J57xcibVOgYIpn
9P7Uh/ZLL4MZLzALa8kQiJ2oY/9PeT9ZuIL21spbuc27pdCpmXmmApr7eOaDbS2i
gSenBcVU53nayJTED2TfxLEu5NtGfiHZBlEocw28ZF4jnMTCFQPsdbxydBnlrYnC
5ykPJSXnpRxRBhtFsvvfIMZFXX+0ZAFIBjStQe+5npYCrFA5Wws2w0T98/7qHXlM
lmaHDA1IEeufHiVUQxHEyF1AbOBnf/X7dKsRm9tyNV/2ESkB8WIHu7Wke2+SK7fQ
eZpa5CxWNHNYLBrLJVrXhtkazsO+jj82ArsnnSyhF42AFrQIeo0pKD+pMIzqv74E
DWCFQYT+xLWCPsIi7uIiubl4NXPyLU6f3Jma/VGouv4M5FKR0zdbrIXxtsZos9YP
795NDxxghQ7iNMr4LLQtBqwbgsYVxe2GGA14Bh7BTUMhWEB7kWhi9esbwUEWXmVw
l1i7VOHm6D3JZ4zaTv8vQImPEzL+Qm2M5MTS3EVm1+uYt8IDsw+PPMlxyF5xVcny
SBlp+hYeXWWlOxz9PopfaQD4ILZ5QSwDTLQiROW1kXIqo/yyiepmK4geVwAUII4F
k25gLDxcbyUJ8jeyN92RCFFLhp/tBeZ1G3B1hkX/RlhcUvvP6oRsEXTdwzu8eHmM
iOaqCX1gZ0btG1H08Xlj5HHJLXHj8xGVFXXggM0OWZk8WQE0JhL8uQaxd9tB+8BH
89/LF8fwfT3VcIYJdJeeHpymtfsQdEencK4eVEDsuNkYZZOiEAxLEeB86/curSuC
7Yt53Soa7pV6fko/cSCgfHNA5zujIKywFbrA0n6LCJlzp/zcWB+/zlBUK6E+MDjF
X1DCK6F8/xIRGz6ef1Hf6xPcx6Kft31wCAclSDy+Y/OFPGQ3yjR3hvXWlqx80NSc
o5+C3m3QyPazghWlPqbMzlR/X88OY4+AwLadvd7Mt7kLxiEDuAdegLFPlB2REXuN
sJm4k1Iy1Mw87T7TgWrcuhNG+MhXFEIKVmVAiXiLrUkeYsjdT1u283zfpwFH3cap
VgtMlLTXEdz4RCeKrIdWiGVwqry2DWW+ocEpTp/QIfj30kiQIWnC/4Tx+NvZGy0L
djhEl2hnzzsWmfRXgEsZUoJqjOojWnwKyQxiWaKMqPk+41nP947NvLV8uf3Mw0tU
XBXGQGDgKMmnIaAC5wlaNxiI6SiOenJ49aJIbR+2mk6fsKXtXcOBFhGjjVbGa84j
shTy5wjmCjLF81ZH2PG9RKaSx8M0l+EpOZSOAt9xy9fLFaszQlMU3eh67frRg7hU
54w7jzhOe/nY00N/QDKYgH1asYMb6l7BNg6KNZg0p1USdKVpOy1vAUbJPjSKT0/B
hXqeLe3NDlJfTqa3Ey3f0ZB15Wc7EBud0gWDVDFi2EVihQ4CedeFcq7Tn24O994G
ivcTeBTqEO1lIh5Aj1968JvgOAk2r+jwfrnOkbV6dvLuQozsXnVzJ5WSI8NyfcpF
Q1P2r0jo4cpwGwso7HIQzNWPelSc12Ppcg6SZ2E50BFWa3l6BDzcy2QuUXeujfrv
PAim0lQvmYfRvF3qO03c1ZuTzru84It/0deEyjDl6DK7kMFG/JoeVWIdgzHdDMiO
mC0zZPsEtun1VJO88UzWSPj2k4ln3Jtj0nFI41uhCA0IOUUUILj2myY8797wlYgA
HBQyn37JdOKjLPAFbMbI+uK78UJImuHAz7fSbL0JzheC2/A7kRq3QQkPcNcjqy4D
Ahl9fgV4kmk3pjFINS3oAJCjACyUYRC/KLMCd9Tv2irH6+Boo4WrlkNoCbrtY3/Z
u1fubXyj+8xXohsIDQWePPpxh+YsuSnMJUOvKl2QQyhMm3enfs8pNYjiaV3Cotc7
/eRfic5aq7jWLG7Ltbet3Q3A8xy99QzckAyXe9sSaNAYrzoj0MAiGOGwg/jd1lVk
aBB/K3q5gAlQKZjTWeITS0a+hctAO8yZYpsvGvKchBZgd6NSLYPeaCqJUwMqM0so
8hbpj7BgwVZYgnU1wrERAX5QFVDzkUqjZEMqSAtxArJJ44wTcopjNcWmgtlDRe1M
zh0boFrFP6uYZFLy0SCQjjTSpr0xNtgj2Z6Hm7ZWpqOzFaR7id9/kB9qD869D37g
p/zj3kB2y5i9lcbNlCgTnUBZDcbjDhTMbgdJ9VSablx1JVu/a0E9YptyLPL2MqII
8X06P3Wuaj1bZbtUHMQezpgziTdHI7gxBg6XxzZDsG/OpjGfxLurnFLxR7YO6rWr
/xNi/G9R+Q9F50vmox6g5CBWcyxHJLd/VGLTsNlbw7aHzpmB5SXJRLcR0c9yy/AV
JbMSPPvQisInIqTxgpTjabyyIeiQ/JGBwlEuaM3dcAuiJ8i9R41IgfYDx6lYJYxT
BfwxjbHJDy/GhCJaphPLGzyaHOLzfX/NKH8n3SMv+iuLtcxWcQW4zVuhNzvdjdOq
gZz6sx7j5actX0OAx7ydr5mr1yIr7Cmsmpbz/OKVZteRlfwGtEV1r6IYTOnoCYcX
IZd/XSQDhOZy+HOD6Ioqndbxx7WB0bU3rV2ko043r86UeqOA5C4ZEFOrvmhWCpAo
TmpqGn/uh5pi/bCrwi1gCFxERwa9AI3EHRS74DagZC9NUQ41wKATTp+pQofBgsjk
EQzQN8EVbEQXAWpvN/gstrJCRWeT1EAwk5VyCDLrTFwxoue6NahUN432OUYHsI5M
jUb87l3QWU1ja35Ov1334+YXkz2305i5CR78BL9tJgKVMwtcxyFE7gmM3FLUg0Se
EZrCr8tpVm7XAiL6Isu81rV4eTYYA2YpVA0v6oi6CbylWqU0ZCL+w9RMTPXETFps
xJ3Odo5KiBnymERI5MJ0TIMp6Jm5VCM/r9yx8Opvm4o/xXRxHyI3uHrk0r0gJAh0
Mw5XHmk2wu/MUZRwK17RvlFghhG7jG/3MiVwNuWjXWIYmXnJRUVqnujH1avOpXss
2pW8oYYHAwL9NZCyWCmFY7M8me4qMVuqn+j6lOO2NrsnCxXMIgYMVrys84EKyHdF
KkIksVi8nwejaNvXSbnZmFpWVgA2L1S5iy3edYusKEYLjwzdXRkOG8EoTiR9DGFi
abCfCd/xyptEehfNZG79ZIYr3hzEG+hwZwRIMJbH/vMjGhldWSUIT1NJIV+T38dH
Cx2YIyeTy0RKd6iZ8ChH1w6RzJNVGCyfttoSmbSNSno07EKLewg5+yMVq5M5XzOz
OLNb7MxxJMuWsl5MCqKzGtBhLaVKlsvHZDbL4XvL5zbZKjOoMUL0Tb0awk6sSEyU
TwwNRnGyTkr4nYNz9D1nGHS5TQ/ViGQRGuXzYvA+YtnGbgCyNkiO1PHiwphPRwVM
atzOFk5MXXzoiYs2gxKSe6UrrmN9Y0m6lJQDPfiQ6SUDMoLBTSxgd4X3Y2k0LNQ0
4ZStPgWuOZ5x1S/ywi2RH9phhXhIcnHr5K3/fEgHWYOWUA2cTUg6Qo/E3GxmtiuR
seG6MClPkvoi0p6Du9kD9i9q7sCf1TFB+7+DyMLit0nH0/16ED/dOEj0bSLO+jt+
uljoa+jVlbwD/9joqwdirz+vu8quKVD/1rhm4958nHi9W5xilC3pm0sLRzv4Lrdu
vC2iJ/WZRSRkKxjpgNcmfl27jjPrKWcAY0DGyJmMg9U5o6Nj3g9qn/l0cAYcX/1P
HXre5D5MKKOgT9Z/tPuMg636nhdfpR+c/zS/iUF6g2pivlxUIj4UIDvsUoT1Hf78
sXDdInL+wpbUcubn7RApP77uLL685Qgs0jX1BHvspfTBz9QGrYbyKCv2BCKllJMH
SCAcH/AtRFglzEF3NegMvsxINC9f/KvFAqfWK5+JVe7/gIZe+zJqBRe9FIp8WglI
CMgjCPrCefSIl+ZLACLztingQyP8kY5f6vW1ot2WcZGcdsbsH2MIKOMqpybG8YhA
6K6BT790cYbk6AV6kQpIugYROWEsMhnNlGA/cGvo7Z4/4RxtWL4WnZUNAGkyjDPD
6qmJiHaIj1787OQxHyI50tXejQgjcJUxdW1AKrvtRf0keZ9G8di/JBq1BzCWAuKu
d9DHjlIU8S/K3b+W5g2f+gaHObIQ+qd4lJr1hj8Hayr2AhSyTLGZEoNZ6vU9uVMJ
p5Q+nqifDfltUwAdambj7OmjFUDQS9A1HYoMmUGlF2OTXbOF/lVFdMnm96C779Fr
bSsy1+0224sFxMtzTOlHkBBRh5RvlHQ4tTDDW9RRhZS5RqVKGbzD/WUhpyDwAOyW
lZ6lgRouYHjobndEdcs7Ah5v8Wiq5fIQl+h2uQ7DhgowGd7o/EsCecF1i2BK5wwz
5i6co4dzbHOCuwC0SMSOyGq9f6qPYDeVxnsARGIPSgwk4OZnCG8KjFGYeDxMvxg4
W4+854a7uPAC+N1I23lLfKYPFTDE8vD/iVahgEPV6x5aL2Nc/qAD8oMTDvlS04pK
vTrHlXBIePwehJeutdEiUrQE4P2S2PRYwUDgMU+sWibnrJY5owSW+VQZak2RwKrT
dCd9MF2UyA+gTY20K6U8cpp7hyZHbXbrNcQMUyLcDT1rDZPy9efJk/Iz17vP0AzK
5DIPWrpn5mr2czkbgXLQA6IuejyyJkQgXZlpSgXgWvnf527jVeGBsNGbihnoJrcY
7jRPrTPK/ChakUNMozlMig7j9n+cEy5NycuPFCmGaihphNf2M3SXF2fhxatgOR93
qBRcJQ2pQSafCRXdGcyBjd5DTkD3Q6JMUJp/3eHVRcrawujOA33DqM5yKRCQ7Uwo
3lEXt1jd+bWG+9VqCksszgm4YCBPxuAdgNa+Qeu0d07FafM2edzjum/I9E1Z87Y8
SrRVBv7mLTzByRgYjWNNjyuwbx+q5EEG8pjmtjnpMcAI1lHa5XvQQWag2/EE0v1q
S7firsvkJGkkfDwBxlaSwDP5GECikxCGyoXVIsrLU/DCP8PHGcF8X/I1cXjiJ7ln
6kGDD5nHwMERmoCZGcAZevK2V/LYYzigVbt2SpfDYSImwuoy5gK2Nz43fXfEjn1D
RSjbAaLvyyHpy97NCx3vJElYlB3RWpqxsalq6pn2aPjbTFCWPM1km1bvBBLh0RI0
e+0upNn/IhSJ0xD6GZ3nGR9SAcrXxkVu9gjF7w7ztcvCTRI4zU55W6jaYecmyKJG
Gn4JIEka1aamMxG7f6+46X0xa3hy3NZC0Ykq0pXubCRTcR6XqOWD72+bzk6k5Unp
mEQjUgtBSIiW221vrH2Yoe/BqaXhlPbeW7xkOJGbylarBmNcDOVt/2EtHtj2ZNko
po+DREE9uaQDiuRJkHi2359bOHr8tTah6SyvrMvvrRZ4qDJtP24WUueWkiUJNd7w
5kxOZWM840uovnp3xNmxroPPeIGPT/6/HPTEPcQKd46UNhww+POURyvMTZXFIzlG
aX9qlMGf5PHuMiY97UqFC1fIvyPPCnH3XQNCCgwFedF7xCeOZmeMGU1GljXEpz5c
GMI25U6ularWZ59PlU8k2hzTCSS7GREJVipBYdM3I/+5cxs35k4jjn3tJVoXH/RV
0BI9r+mUPWJPLMriFZ73qTKfJ6Z+v6H02XLuvD29mFuQkvHXIxEQ6n/WY0AyX3Rv
PbVkjq88bntFkJZRH8OFX34zcXY/pVZRUthAYt7yR5HCxAqTUmgp6OIBwa/2AnPM
4jIaWzwYAbWK3TYFgx7cE9uEfED1XHPpMSdvrdg7zM5DlqwBqccHXLof1vnJ33g+
Hy9mUF1lcR1NfNywkW9wg5jYdIYZj0VLv3ggIRuF5DuZnpIqgfmJKehp/fuS26Ok
qUACfJBUdcfgHInJmNtz176xIq51u6OlY2HRTyty776/l9rRU3gk88DNsWDW2VoM
/OYTmEY+r5tjB4Lykj7qScQPo/hV/7CdRb8hKWjRCme9vUd7ptJg/rucHvpciydH
Bny5b6oXZwkykKBrdy8V2ydO3lpErz6Ce1YZGj7nQzZph+gxwMLQmo0Rq9eIQ1/0
aJnSmSwnJXHc0wfh56UuLfbWIJ+nbsAIQ95pRs6GTYtN5RL0xU6d7LUJUrym6Ll3
WKkLPwiIWTz5yya/PkKT9yiK+kHGNdaBpjMjHCqGGiO40YsagoxkF2F8KPAp75tC
3niEtAK8awD1RmshKrWeXukCz1+Bn9Q2ESsoovARQpIHENXCLhJTry7/f5BrIfzK
vOsQ17B78KmuK+Ik5NV3zSPwE1mc6cU6IF3L3CrYQ4/64mxhhqCAM0yI+acymE5a
`pragma protect end_protected
