��/  x��(L�5��i~d��jx�a�����Ȳ/�t���l?i7��6w4�o�ȑ��r��g�+Sg����	�ߗ�-|t-�,w��+�F���#T���wl��凕@���>�H��Õ)�BC6f��r�������q�1�[A������:[����Ь������Ԋ����H����#{@��)	�<�:3eE<�᭮��yJ�Z��X^dݭ5W�!L�cSa�&,�q��zN8�[�cӭ!��K��,#�U�������k�#!�ܼ�jH�i!r��$�ۃ7�g�ۇ�P��J���F��dN�[y��Ov�4�eC"�Sd>S�}���/�;rȅ�d�a�e_�Qx�¹����xc�u��S�@�����w��n��M�֮a�G�����U+�e*���'V�!�}W�j�LRQ�=CpY����<��9UK�V�"��	RL� ���a6�]x�_iX�m��rʙ�'g.E3e�v[��fS�@�	$�%���U=l�\�|���-���h�YL7~)4����x�E��1���L�W�L�>F6�_݈�7�2!�Γ�j#dC���s)!U��tY$t�lE��?7�n(L$�3�iB��6��s���˶-7SOg�ș��,�Q5��Ɲ���#���w�����g8o7���8N�$K~SfdI�k2���dR�p�^=r��T� ���P�)�q�e/*=�^E9����Z(��V]�:[.��7��d �N�<�湵�_k4C�oBG��x ���34����|�����6p�8��ܩT��yW�=	�b� V#�����(�Bk�w6���?�\v!��q�� 0+��y�ØVi��s�}�r�yf�;�������+d�Fu����q�s{���I�O�4w�*�����a��n)B+LQlu�(K�J�
�e�o�ʬƯ�� ��2����v�G��n�fnW�� i�Pw���%�W�
�u��Z�-�m1�x]
��1�.te\�JW�e�i=��%RR���մv� o!�<�C~�R�K*j)�$�a)�V�%��E��������]y�}�T��>(r8�4ma��vJqᯘ��𔏫����1D�Ԑ�$��'�c��_AUvo�����N�g�4�39H�偽'�odC��e1�z}���u�l�J�W/`��|z!���k����`
7���x�z�>���c)c�i�Ԭ\b���q&��<�9���:�.Nvf�@��eSʹ@��o�H�Z��A5x��u)�=�g}��aC��&.#^�1�Iׁْ:�z����!�L�՜嘺.*q��M�^�����d���q&;�"��BX$L�G�Bٌ��+,��M�[WO�6�B�'��7�6Xܯ�,H;{��RV`U[&��V��	Tx�^�^��TR|Q�V~}6�躆�[�U��c��uB�����k��~p
Ŷ'���j�,-e��?�u���L���/F�́PSͭ��K1�:y��1�`�m�u��d|����%����M��/�2xL�q��