// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Eq9N5CcuoXTDNEiAi0hTaYghG7yrOITENTN26zJfCS9z/bU7z62mdl08H7yWwqI7
F3hJLiF8nlwgo32OwAzNmCwTKjdwIkiFvxr6ugIDYGjbHq3uD8rh0+mtEXY7FSuS
445jy14xaH5oXU2FH7sovw3BdBwPXwDTRJZ7gLqOiOg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5776)
FHukAjY3E+fwkBsAZuu/70nLhHaRpNMZaJoaec9g3qqvhP3XdnYFM9TGCMyt3jCk
p0+6k+a8HrIlJCYNrxboC1TLDPuZrDcYu40xu1K7XX3XKK4JN4Idt8n0Ad2TgT+T
fRQLC4Riqgdtx6Xbwm9Wc7z1wGUF6bt9EWZdr6mVDmo22qTXDaXff1j47TJQwtIn
9FjuELVI1BV915JprzZmbySl59C62+r9fKg2a2yjA0D0BRYk6jNLZHwcgSPO+sQw
1x05vsG7mLbpZRFzIsmgEGnN5bTnZOBUXCOnqOGjAqw+DODAgbaUSNGgRq/aHwI0
ja4nar7p78iFJ1Rl+E2tL3CerZJIqq30avkDaWV4Ah6OF36QL/6q9PppHDgApecY
jwvK1b6nz7+6vCK+rgw1TMA9vVjoQ86eVh9FfpbU/wec89slT9n+8M7Smj7QnCkH
itRlwJyIySMOguj4RviSe/rJtoZ4grX6OGLJ3ort/wNof0gO+xxHPIXsVJt6fSs9
1FNDO8rL/FOzSZG3CfKSOACm5HpNVt62lyd4rh28NsxJer/rg2fDFALHcTeKEgdG
K5YtvkI0Uf91NtwpG+/MfViY1cLYUN400dUT8pf+5HCZlq/H0aH1ACHH107z+BMO
GEABj92469zOtj3P9WRD9LiSDoZxK4LmYppB98OWceY8XdDoLj9vB1ibFNYI/9tu
ASeirUR66KtMipogVJ/WgZ3TECXyxbsSL7ngHVZDTZKHZPFVeUn3WidGY5i7pq/2
yPzBPq89ASzZyqbJlRVEuk7u4pAWmneVWn9cD+st9OFPDXu4LMq8GT7MNbkqH0wY
ArelEKAWQi/EgZzJB4abuY6hLIqTBWbO25Nx6YbPA4waVnjvQQKhitv1iakEnZzJ
U/OYVtcvOJgiFz4cKxFavj0FkfhkMoRCzfk91POXHLmPzA3Y2WfQktq54uMMbg/p
umX64rVvwz1Ko5VkL1ClRuZUSNZkXsnwKCpA53tm3VnhDYTiRTbPQV8fMy+3uus+
0l/+QCD2V4Dk/7ZwwMyIguF4FG53UPkxsLfg+tf+RGVq94GlozZW9riC/dv6SDlv
qLWbwjr7Sj56c2eH8JZ9ipb2blU/a8BvqVoxWiTTMxNc2Sx+1aUWz+QhPk0VkMjg
d2oTzGFZ/RYVlLsP26J0oo4HUKMHBKxPR4+9ZEGPzBP0amdsCrkmmHrbejd9xXW0
wZRQX60vBB1jZiSn70urazL/l3C1p5v83esPavNOdx9drg8LMXjSFmGcNMrqlUP1
DPj5Zv07pRfGzgRWtR3IWYVzySf8PclGbHbjrfRn3vIyMFhQQMBauc9WPrNDmPPl
tqY407l04Ow6bkn5kDwDBpeb7Ak3SH7gvRh318GOsNVWJmxKGQVj5xAYeew5RMGq
DTAms3A3pG6hbHQ3tCgOYhgMav5dEiCVziUiusMQ3o/GW692thSn0EC1v93nfD58
RpimwGXK/xtFfcDvfIuNI8/zkwm3y3xW3rhlTx3+X9CDcX7/qoBnRXg+Mo71uAnP
VtoO0vMRSRzvM4JnKeJA5P0Cpi/6U2caeX1U5qZ0OBUne1OhtH53vwW2v2LPykLv
NFtV1/WTgH8zvCyC7fE5UESDeZXszZgtwrEe0KjHAAlURmp3a7Kd+Xeu0dTN7uk6
e+qODI29R+p+xGQddSXNWx7PsexdS3mZmeVjna9rAZ76fCma85/YQOHDhMlMJFqd
X6HgH5ONi6WA5tf/oLjkoDJ1U4IyaBjLbWjznGkeMPhxM1ycMBlEJXmOmzixU6TS
PQ5hIcW3/ZQT7fVj5z/6+x6zvifKyVJON93IRUiAj/fg0mFajW+0ipKeuNPHpnsY
HcpSAGMNbi7h5ruSJX6Fuu1m23SSOfEhkphzoO4FHk0GBchst/VVG5Tjrj4s3JMP
FN6U2g2qrqY/rTc3h6Kza5GjeLfSbU3XNLirh0EEKY3AJm3EiC29VUGKgxSc9gU2
2FyPcFOeZtEuaXNUb30DoJ4+Nd/7XDXgVn4jq65eOMJsRV3gn/evkFPvEXVPW4Lb
yvv2Lq8oqLU3WpZ7vfKXfdginwnCW6E/+Fnj/JaicMglyRbfL+QNpBCwawbp/TT0
bfT3bkgbIfihnd9iUIZQV4y4W2u7E0eB6wiM2j+FmpYlC8BEy8xu4nOuHGjWJROk
H3lbG5FHAUrYJZAPAn45OFBqNFnPRvzmE1HqvWkWH1+BGq+JlMxvQDQYofdqu0Cs
WSRVzJy8h+ngapuLx8QHIoX/QLTj+FJmWtKSHmpZtCFjoLojZyr84vda/TE1Oz5r
klT28nRMnar2kRfbRcZdgTdjXU9bYWiTRP7/GhtdPGoip20wfC+pLQRZ9JnVwpvi
PZ+KBZkryEicBnsHbZHwDpv94VrCYB0LUGCtQAnV6mczP9JHqbje5gQb2iujJxi0
wB9ae5WXoe//aDbis6zhoTFs3mnTp3WtEJ4wKGG1jQ2bRBcED4Jq9YOnLTkh8qHb
Z0CT63Hmw/WR4+Y1zBj0SmcoTiNhYZoQ/S97AFsqe/CI+e/ddkR3Zm5JKqLOhe4F
PpDCYzL1OXDkEEHnJpzAXH87GwdolT7onRnmMJf6HhnGHkYAIYq9xzMjKVg339ho
ISg1k8XafQqbh3TMQYpiTDtwRliV6PnH7wk8x0Ms59tWoOiPRFNx3gGDdOrzhTUl
apavrC4BCpZIIOK1cxQmvJ+GEhrm/gupphpYmQENBx5wKD+t5xeOyM+iAEBt1O1t
CyCVwFbxpyAEBPJyi5Q3HBJSSzxXGTdGZn7NZxxG0CZRAnWmQX0EXUt2Dj6SG6H0
6x44041UKVjX+lIjs9WaZGeLgB1FWwhxqOWywcREwynSe9jgCGjKIC54gIso9ZnB
qWhePLChQEdiRsD+O5QOAMpT3VoSpJ/9AZUgqGdIN6fRfmXAyqjh7Rv5A68kVwIx
sBc9Lw5SVxTZ7ZTD1nSmRaZxrhFAmDdytnVv6z25c7XfrRqT0MBvAokeluP5Cbzk
6xz0m3RqiRcK44SoBPNmx7c00+lxg4LOGPTZStYa+T+M82X+Oawir6LYznSHm4XK
+LCjSEzv8vQrwBLAn7H6wZrnwPdIhP3nWP5yDvkgDQwISrSDnp+XYLGOuR4fcVhh
WWzeCXU4CgCS6U1F2p/kVkSABLPLh1MXD1Z1KHeCG9gsUA3AVWhAuOyehUegYeH4
LVj+pRkA5sHdcbOoS6dUV8KpTcAhG/hxAZlZij70tr91qcORtIWilcnuaqVZC4ha
yIyVfcicEkpULVf8d9mnLjSCxAj1BzxrpscWpMYgtGy+WSxmmVVNxHk93o3+qFj0
eVrig2xZ9KBFpSPeRh5ycN5gjByHot8oe0uRa2XnfmernH6kYLE8vVrdM2qS2GGF
YwHVQcyBaH3btZJLo1DUGwKx+7h/HvGyH/vRydgLAoyZQtXrXewOsdi4Yb95Ws++
2BR2jVBVkOZ9q3zvga+q5Cf8Y5lt6VVfz7vlGyePq32MG2g8/OM+eaZucUYoemW9
rLtNT3IyOYT2RaXH0RK25kPBzOC3L8Dkdh7lRFXyqXLc0FYl1Pum2Gc3TqlhN+Kv
3gHOdF9b5jU59KexwVcMv7bFK7PaXUOqIQj+IUQZb+nLegipdC+6uE6OM2mdYF6Q
bMt4RbGzAoceXTOkYdKRmEfdh+Crwf4ueFubHSO56Zsa2MFCLEvlZg6t8dDyl6gD
v7Tvnh/hKtOwWVpH4GT0uz74T30Co3tDfh9zsz3FEWbSw15OSV2gW25sLhWaWflx
M007s41gtG9NTsJXW6TGyxPrIVaixaMYM1gbeoJ3uvW4GaGc58fBwl4JsKYyKPBG
SAH/VD46P3yoNtgIu7KCYTef8lJNvGRgEne/+44Tw31tw9jFt79ABt3bAxGE7RH4
g44UVa5AbD+4zobV+j+9xbuyr5lbUKAS6LxuRAVim78logNx3DcDT6Ul5gEvhV/r
nXMOBYZzCfrsEVewnV3PnvxTa+k3W0jQD70CR4SWEp6JLrpuf5Vz/GhyRwxb1NzG
Svw3bquwv5rQvgM1PAwB/wyGLSCt//DTBGO25VDlH3Y37MmcCTk9AMZtvH8VBLkV
CU+vvESAGT8Usypqk4M8uJkqdMJmvK1u5DnhIVog3nzNdMsqpaqZIhk4sNdwjtuN
HhYfgy08c3bqnqLxpl5hT4zspAtv54PjhvXFQekFjAlRNgP99dtZsDpFpuJPa79t
94YSXDjCMDQUwneDC/kGpcdSIFmK2+Gk+A/oCtrM3wkDFTS7HSWcfxvhEj9YNnsD
LlhIjFFID8jnuNYYopn31xmomlreJYawTzEnQsjGPj1AKcuRBaT1ZEldyaD3gX3k
bsM4bQNG7T8HOd1a1mRYQQZ6rn9w4BbmMikrNBh+DMXcc6eOpmZ9G4qCd58CcspT
BobGIm5T8RH6E236f/Qn1wH71D2GNgRAgUb8R0ZuOtU1Z2+4NK2KsPVncPTIDxAM
T9/5Rq1+b2PLj/2m4T5Kj7fOmULTpcYG+y38R1ChBBP8fRCyM7q4Xvd+Bv693QRx
f0dakeXMuAjDP/WSm/lGKfGuiQqnA0VemAxMviO+0aIh7KiFB1jicwKBqsF5y6wQ
XvqzUnELiNpBrjxJD5AZUu0chjwLr94TmrNYuQvkKUNlRKTkMF8sK4axL1aR9TSx
IQI6U2vZPlY/lB4TSrZTt61wc1dKbYkJEPQ62y+GTPbfR4FYaDaO1hI10K5NT8s5
ieK4ZUpOMHd4zrQo3M0/NmpQI9SBUCeNS8PBCBe0x3LypFEgQesyzcfODIbn3RbQ
BQcyo3WRJSC7t/CfsXGYblbyvSSS1ZswWUhZG/rUPbnKyoxlad+dx1Eou59C2uA6
/PxM+H54c4GVJyuASkzXbe/pcnynwJCTZMPd8rW1uOkZZjqI/f14YXTVjAQ8MWye
U/6PsSGfyCQaDO3aGykxcJfEEgdltNxQW72mYnSKwx1kM5os6pTtw0WusozpKif6
SM0YEqYDqzn1g7mUhEeB0MtRZ/N7+vhKbPTeePbseu3wZaqtjRotyZFxh3Tor8pc
cLmZcG2HaDff9rYAeyXfb7qu/xUJzX/USbs082XkGGLC6ym2mjT6kEHLluJDcEQf
yluKdjtcROb8MN7FQwLRUqTBSgdDMMblu9v48kJL567miy4u/QtCC7WrBNREPR4O
v/W5bmvX7oczR3L6mV+fOEskmdqButJAhnDuDODyMh/FW8AX5b4m6O0DpI9aKRWb
Qzeho7kGi/e4h5kYCtOF7bmX9fPq3G8IbyZOpRBDFY3cZecS1/BP77bRMJvYDMRI
rcOaT8Qr4ZhP3/dWWPpqy7MzOWGQFUVFkCK4XKEO8U8+qRRPV5QpaIM1yBLAFGJR
KFl9w1gaULl7q7x9ENvGFmPMK2MeyGAzhGRKb1+mpQpNiuNCx2SKWLZAWGM0P7Ei
QVRp+YQpb579JwW9qtou56Bt0lY3s+2gxFEL4v4iUk2Q2vJH8XliHWWXJiSGXdIV
XaC7Eb+MOfOxw8pgzpenuYhhsK1MoyKWKZG3ECgreZhVrDi6+gSxHNSW3hUzMbWd
pfarbUL2XVsdq8u31eDzZh8TfBT5hBo8EugL5MNzVrbwe/zTUZw8ftukvWPYWt1N
q4/zIVB4+zc82sdVH1wrRNxmpsiFv51e+STKfOezqIo7Gj1biQzzOLLkTvaq9A4z
D5BnEbL8FwBQHSB/TZWiryUP+WXII+Rr0HJAzUe325ZXRW8U5AuFaYFT26UyIGl+
rLnjahxO+VLzHxdM4wCPrWw2n6H3C0uwUXnglGacO4L6WWETxG+diJc4M0YovHH8
FxX5Zp1RExdhkLgZgF8NwEpl1dvGaulGqKPfDrSyWp2d6wAOwft5Z03G/8IOHtkm
3Tq48/MssrMYtyRPUP7LEqoZaQk6XmJn5Cu0xyrLaXLSVPm5HeRxj3xlzTK4cj4Z
Gfv7aABJZ2ICp3DmOje1/eGcTDJCw3Ipdmtyrn6HUr5WVuHLZ0WgAr6rxW8sxaP4
TDs1Gw33VC6xl+aPK2qLACOLZq0hgYA7oeKcDIFS7taJ6kegniKbPHFOnCH23kS/
/MhY7FuwkQmyQNa6qiwDbuDmebiauYO/mpyPWqRvKJrtSH5l/yBqtbDdKEWylIVE
GWGt+Fl/E2Qtkc951AdNLrNE72WA2vL4F29B/WViqewctfrhbYRtGGWCeH9wuw/y
MGVnHbsJ7LwlTSUEmaxhzkJEuXrwU8HgK9caCckexx+V8z1Q2LIfVTRF/TRcja3G
T5xLogdMjdzet/JsE/UHLOQv2KSeGnX7UCHRBGg7hnDpPYoYnSoyujCIQJtAfhFF
pQ171FzGkwLyIMnde+Fm/OBESWqTwMc6vb8+hDbfp1aPc+/wR6ETCfoJBcaXzSzo
MlN3nvYcYM1Rym0Oc35otQ3xwI6CHvvyTFDCLDq5BVzmSpQmkNmCEtGTXzbbNkaX
sx37Kl6GVruz61mFULcFUSXL6cHo7zmoA1OsJsHubinh4wSZdo8ku3AyORQPaLCG
kIp7EI1i8XS9p+cJMDBAmCZOAdvJAg8pNpAGLDWstuN9Jfw1oXTBxWYxKixTxmi3
royKMA1RIEiFGK01pYTV5VQmA8bemjRn8RseKFE7d/brCNNjhTfG7T1t2dbdUs6y
FdrClLowNx56GpvmvvKpqyLKgkO8R7q/rSBQ5b4oScVeqylcE2KSkKWWlk/pdRV8
SatylcQhkJMueVDhkdo3Ct81yw9yjYeJsXjNfDWAO1JYwCWS9FP1rHb6b/68FSUw
EP86OeVk8IWjjpNizoYZVWZzA9rdI53zDAUPEi1Jab1xZPhkuodtyE+l4sEHvqBM
ruJ7h41EAmPQVwZi+0E60G1bjC4Ec05N6eARaeQS+Tellb7xgshUA7mky2sPz26u
mt8s7+7GNDEzsTt3CqBbARY0YYr5HBAkTUU8Le2WbWmlE8YJIyTRWDzzz1xH+q6U
kpBZWpMwwMmoCyE0wVj3Nlc95/GXzVVWtbF1hkx8itVI4ZFslshthNBEzZlTaN7H
1ln80jmAwJEmsfvprYa7DRwILOrETtDQYnheyCvX36Qs7qEzq2NigvJ78YkWsDbt
e+bHv3Tknaefti4gYlATSN8ge1ysO68asFuwEPSPsdaIVtBbR6Veiuvm6BIfiLNw
fEWvR7XHzs+v00baa4acvDSRjTLdMxspkMKXOkVkMmfdO6vT+aYeuHqhiAJOsFzM
z00CMnNVwB0KXY5kCBJmGWaTJ5mNuGWLu00Xl35kLvjilTlCzX9vduesYFJK00bW
Oc767HHVII1QXJXxSeGhBFIx9tc2D5XC6Qo4r28/JG3ECtpv6C8Ymt26PWH8wuzo
WmRX9eaVzMunhsP/0zObtStQzblxBy9bYz7fRiIqrFcDKK0yW2Fbc6qU6MTA4GVI
1DDluWYVdn3T5AO9KaX51S5M51qzH3sA45QovcjxFMA7ny5XOgE6mla9gHzshPTO
D7wpcxjzqh3i88wNVR9EmdlzwKY/QBqYpxtg9bmei4Ml3f03AVPr09+EHbiDG0/E
i3WLhjRoAYBd4+FmLmlzCkea5AspdmZFCH+1xbuQgkstWe/zv1FhbdULgy0672Iw
lSIrUuA1hLFsx/1YCc3e5XPKdf+4DDxjA66dXvw0S+iWSZzjtMq7ML7KO3Jrnhiq
C/n5/tlWm63LjYS9qcS12g==
`pragma protect end_protected
