// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
h37izpGuYNHTX1mL7wiZMZzsC7mEMebK7fTh1eNo1HrAGwhPWwCS8slCN4BaVWln
jMVWcVZJ5OtZCeoy4S8w08c9dugwAgpCMYktoXioufpyF4n9i6FX7yAWFxN/6t05
+/7x3Je94kCZMBDeNITl3NCYV390OBhXuXObqxbqpa4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16208)
CYL9wiOGTDX7LBF9idIPTKxZ/yw/rU3mF9j15hYbUWAPgPPteGWYU+wA4v/Ug2Ce
oV17CV84z17wk1VpNEdUleFIo6AjsRgBNBEygXWYhT6/kRRbSHw1pJL9w+0GwPQB
OXdBw6Yd+5O0liMbyPeEsVYaaTDX9pu1vO5psBGM5AP+cnwn1gFfNu+7vcQmpDLf
fDYGUuZG9utD93bErDnuwMocr/r5f8oOiiianVZTF+Tp2RDD5ttqXEdVB5jzkJow
MLKi2vSk5TKFjEjJLQsYZjvSXXu5AlvYLSjckDdrBsTfXXFORPxhV1D9bNqfX2K0
rj0iyq1QAyJli706Gp63qmC1mAOdRUA1sS9rkz3IrLe6O3rlngyk5FEWC8wsRnR8
GCILjkRZTvoNODeJFJSt8/XvTzgUNETZemahzktujfcTa9WGbB8SD2N+gzaq3/7v
mHB8a0DVRqkDHp4FzsPZAzURy7DLVnMre93ejHk/autiVfDqVousprNZx13C9vPV
QW2K9GGGc1oxgyCUJr0Ro2HbeOHPfkW80uPRup6KPiMXcHYfYLh7CbPDO9hbDJ2r
GmQi/GyS1qWlLwJW+IHuMJB/LBA1OdBHLQOYuwXItDEBvhbN5bfsHZ9PXuevMVTh
gJsNzqZ1ey70gYrTU1cXT99HbSYQB6q0Hh0F2wrdS+z6OGbuCMs2L/Weq/d2A78q
Kj8jQ9F2Z17HhXUTx1ZQkLUDG0icmKAy0gqOPJbAH/tSqULF/8QGU8nEnE69hELH
nb1YIbHJ6zvGgOcfKO3o9F8pxpbvDbYLAUKQd9Vcs+MPFJEAU0QTPF6SLiWybhHS
y6o86JrOagaKBVrrV9v+DfpoI+gNpAYVmuwzsayIIistiATWi1aODa8flBZexXlW
JMK29NA2rO0EZob6XF17aKW+He4vky54VIz6CBDPH2Tj8pl/31nX+9IxVtGifFs0
0U4P3z26ml9X39uUcXWiysiV4nYN+33JHQGfPYajEo82H7eb4iqZ+Dqf4ehM40RY
m3dzm/GWF4Lqt9TmIbtxKODAyiPd6cnkMUsmaK0PaFSxqzfgvuhu8xFV7W2FLnkC
OwD2+cokBpaiYPy2Sm4hMiHQctTHZg6PdimIgyCmqBXD6B/rifLyKlJxCmfiT0No
vS4ofUQI5XcL33INvqMjtSN3+t2U9nm87GrM0b2ova6jIn2ZUKdZcMVV1bs0RNo/
XThoVjZBJDFvD6ZiNnJ0XmprY3bAHdWTLdO9KssnaZOpJK0ZSaG82cleIc8kwdAj
xfCB6BNPtv0okL4dwds+2wkciUiPJesdCDRog/hddJalrf/hv9NU9zF5u2qk97ef
bfDu8vD94kRDL235AlZFiTb7di9z99hqLR93gzIbmqDr3lcuRDbABuh3XpfTiOW3
YESLMQEdWbNDGi7b1grCOMOIIfoeJitsnhkZzgegbeXOzv962Psm7p5f6uT/gGPV
2ZA+zxyXxIPbklxF+uFXQO5rx8bj1Hhw0r1yudjT/DsAp4DlVxyBXnMfty+YN7nK
8vCTAKTJ05YZWtcbCyZjE9U5/+zzuhfVQzB0okemBCBW++4o6SSMo1uFLs5Rj/aW
23ClF+gEx+3jKha8JGEbfSxLauYdTPDpEvxCXVU58igq/VIpVwry2j8KmxmM5Xjf
uD2A+gsSZs0GZTMYyHsdzeqMf0Zz2kmAiqemGcAgLEJ6c7QVfn988maJ8+83mLv+
F4BhB3Zk0Cd3msWt28OqrEIA8n2KTxn4YJmYrpI+pHDfrCsLD/Fzi70G0ALKrSNg
wjxxsjLS9CBmPR1qSWcp0n3GYyMEVyz7hqs9iK4rGG+pbJllJx/ZTip4v1x0ymYt
FV87RmUPey/FeSvd/TWg20Cojghjz7CDPrMIe2VW8jO04yP5meWCk45vy+x2BaKz
dhak+DNFx96QOF8w+nIbpR0erhfsyAbKSHUgFmmoUuSd0PTo0ZI+B/cPLuVWx7NG
L3Q+IHR94rjy/+68zA39Pdumwf0g7fU2eImKW5JxwEdnR34es1rrLWlcg/vUOV1P
lk1Ar4Ulm9BUnTUUdAq9DXLfTsjb1A/C1A/nsc1OtoPoLRP/XL5uFsN7Q2ZUKie8
QZ7MH9hDBilHwd80KSd1ZbLn2m4dS8zzbR0D4tGFAN5kj7IXBD+lSx7Lg6e+EptD
eiyF4Iw2jMaxAQ+/8ajSmmyjH3tLrh7oRw1Qy4/e9Q0BFboJAW5V+gurcHilSMhC
6Am6+ncjsjXBX+LHMWfV7tsjvrJOubdfo45xay69M1P6+NnssbVnZ6aniuEDIZlx
u7/mKfUk1v4ZGTIkrfrEm5xFyTvx9QSHHWT+YD9XqCEUdRrRWw1BNp9wjgBuLpQ0
zuqSJTf/knAY++WHuOZTlhJY66jcF76JzY8PICjVhac3X/YUF6vbsnw70hcx5FSW
+L9haZdR+ky2FCjKcDegGIRo5iyNfUYaZe0nNo1MMCL3GhDWm10nG3xHPxrQyt4w
GwtJVshMAMsEZUHZQ6TMD6YNRkyXsdl1Gq18S0ApC4Ms0jpW/gbdC0t+qhVpvw4O
7L55g20sQQGWfoS/0a1BADci5nxYnqv1Z6c4MjvU44hnIjWIn1mguToYSpeTI6rF
MkyNKngfGE8CMb2RuuHx1r2/ZO9QnOvexRTyMW+P0+ui1aRCbeOW9FJ/DsJgChfs
MOcMzXljWRzFMjH0hxn5ONAYhSqJ4q/84iB6ZLmZOoyr1xSRUgDxV1+b4kkp1wFz
juKx1IyELngQTyPD+UXVowfaCd6VLkDx3RqpzrYFojU+Uo7iz80lbY6+2WxVex6c
rtB+oNYnlwDk6vZ/U4lLPpT+evCpN8nHpEMYbMJDRh3EKU26rpbIHuJGkFiKkz93
3Uf/zP8c8cQOctRdz/6ruOGTHSSfewWy517+wg4RJr9u8xHUj/+lIb/XSkWdDm0h
CIJUavnI1/CnF1tDlACSYPWA6GYB9mziqKuSicA5plUYb2MF5GBcPDK9pQ12rm43
Ltnka5yN9WufBWpBoaQdw68pOvU4SAhtoMq7TMLHdePzXab1i0zh5+k7c1R+9Ldx
qh84c5hCPLAl9tNuJDXeobjt2+0WanhwaNZMmbeSyn4/l6rUIo6kavwtvguaQ1xz
BJe7FfnHv2KiMlyvtZiwZjEHVlb1LEnrEQOR80BG8ReqMW/hiyKQ7gmppw2iMLjC
iHPmI5R2IQT34Opky7NCamC227IRFrs2L2K3TZBeTUaekKvU+/bcbb85OHaL6t49
Xwzh14ekoBt5n5jS2/l8QKHrGDSCEgJgtWISQKfNxeeY2c4dwMTw426MLWVOMIKF
jXdzQ+Z0gyNTs3J+bUfb1mM4J1YdRci6jPF8E+oCHdxSy+uCbiv1aE7hYzDPdbW6
lZxLQfrbSDqv20sLI/VJfx87NJvqDiEJynMsjbnuehTJWYGOkzXlfrd6nPa/oYvR
a8Hsv0kASZg+Oe0lKUPjSzXoCLetUoKFWY5M6fEWb977utu2OZOEAsrzIbKlg1a3
jbFAXqrjj6YJFQpjZv2rgK46gbHtMyOBp138ri1GQCCtYBRcKBo3OdrEUgFzKqCK
KVytVKOVPx+LxjDXyTyzp8sD05fN4CQhHSPtirWnae/L2DFt/YS8mHUq1FUqTIko
LimFAJ/ZVrSrntXMICBLfKY2u/GUhspEDYoQMfXjjjE8YirksxmedbXYaxgYc3FW
CTrRaS3DUdqTjksVOonMfNwjUu+mourkD+LpACv1J+7eOIWzX7SUkCa585t1koRr
KLESeUwcJmlP2k55zI4nULqLV0iSi9vsfK+Ey8cFyTi77jHgGGRO/Tvsvxkyl7sJ
k+Y411R9F8tpbJf5IDOKmxjQS/S/M6rMkHbiIQfdijnh9f5D6P8XZb58VKp6aSRV
QNCJs7l+m+g9bR/bm/dvKUDh2fS3pG8blNFSJlUtjyon7MlD0iq/QGbIpcKrFI48
a8665QvE8bxtKtob/wr2B7IaAeUW1ylCR71oBvywS0b/pSnF3DDvzCgW+22enJaV
uUmUH3B3ei05wOb2x1vHwLAOSPfGuQfyhPQ+nW35GkV1PR0bRxjD4eup3LMuwe6+
Z0JXNyoVofKbAWX9Ze6nDKKJl+t+/pi6piPjT5j7FwoJmrAojOirlepcZ5JKEYJY
nqATMLZF3mIJ/MoD3vcn1sFuUwzD3/aOJnYsBluyTAMVvZcBbj21U0frt8WPG4Vg
doR1Mpnb1HsoN9h/2bTJt9mAa5mzDTnPLSne5KM4LlPtpzQnTexwW7L3HEjtR5XN
Fv4ZrHmflp7Wzs/4Pb/VCYLOE8e65rGpoPMxOQWm0j/wV4dJJDxOU6IwgiZOx++S
QDdGUEZYsr5k/iGf0IigTKErtlO5hLfxa7o3uqyGyD+A7Xw1L+wfhJG85wsPVe2D
3HPODJ9FRylYC27Yc8htGxELKclI3jWiDQsR7CVR+4ph0x0hrHIBJwcxsrOYetN6
7d0c6s/zvzWH4wNZrSabjh/94DgPXKvcxzJ6EIGLX3KmE7nITv7GIpYsx1vcx6S+
ihf6HzMQjM/L4JluSXAIU+FehGIBPgUOnK3CxIs/274MrJI90zAH8oXtCwEvL67A
pKHe/tw8K407ubQSa/tzrlVYlQr3k2epapIZaiaKpSjYmrkqAW7hTndTFliFnvpx
H5IFl2fr76sNbZWIssHBDW1zJsexDfp8wcLL8v4QcsBPkFgtiSww/ffwgIHpskxb
kkcEfkLBNV3i+O/7qtLcf8LGCfaAGMj7YRTXgOUhjXMOwC5ygF3nm/DuEsU7f6W6
ApoHymRDviBWVcBOSB/yrA6ugjwifMxU4UbDVEpp3mE7w2Mk6LHn8/e7dt+E8EAC
Udyqsk8fi6lVPiBS1muheOljS5QLZ+Q+8zbU9raMaId0aenWdPzFSETM91SeCZJt
u8mLpJTAaRqInZj4T58hAqzyTPGLb59IdcSxBCUlLCryOFTz7+ghNyxqj7OmEhrH
Y0jHcznew8Xqs4xNuId0fav4g03htpnRalv0Vh6zPNXDtTkmrWsmvrHZxiy2S7ke
Zzz9Y0lL5+hY7pkvhRLTDSNsIDpAjmfjV+9CWsVPYyH2xyNyIsGOnhS/NstS9/R9
EMGGe8H3zP/fYuwqAUoYk9Sq5eqvrVqQUYJgWDJ0TRtpvsbLz8buHNGiKxZqu667
E3bvysQV4MxUjbpmpXC+ia8wIA2VFizNETFENz4HPzYI3kwSE0uKSjYeoq47039z
FchnRoSLQ1bKzjNIdBMHygK1QxREHLdymH6SvSklUZVaO8cSC2EomXIeP9+JQ1B8
UrWkgbv51yOHdbWvQFrmUzd1Kmhq1+3Dc23mov8VlDab3LLaF1J62Xz+B0Mzdg6S
e6D+WPXsezPTYdz3VV3otM0Es8Jbn9GU7F+IH6IP5fYQB0lwnclD0c1lHtqBoQAi
9jF1z2odaBJdLOPL0jnq9mztruZhtB0RIpydusLw6hqMN0TR05Tm0RhLui/Bisfv
UuE4MFKG9Q1xxQXj5RfmtFgJeR7bZkstrDvuFNlxgsbX6D+cVGDPtnndSWA1iw7y
lTYkBPQVFehb895skL9NYSAwgjNQ0fAvHiEkORzoXcp93ZTcCLeC0GnixwMYPbN3
+CrwYWqLK53oq/YED5zT/uSYgYaNqr8OxtmW9sQblC5iloCioir6cL+I6OAZyWUX
uVVLdyyyzGdipg0QCs7GWV16wr5jV2O/WQqH/8M/D92+IkD8yXhI+lq0l6oScFpA
b/Kp886Y26itL/JcTgBXPeXwwrGjZGpUNrFhgKwrHmzu29HmfxMtGTQGtIuNqxiB
fxtzDsUbyZjEfy1lM22jWx3v7yn09DgYwF+Jbrmyp2+5948MDegFEdKTm0V6zt03
pnHN6tH6btVgY3K3tc7Y2VxjEpNKtwbmD656HuzDw2jWOXBmmF1/Oe/XCJc3SMBS
4kSIYwlROdU7Pwg4NBGlMfvAP81QW2+Oe1QLg5R6Q7XQ+Aff1tyd3xshl8kX2Rld
PUX1JrCZvXTBYpZqCv8SU2CukPGPlC61oEGJL/qjc9ceBfhZ7Zcd53L8XfrlTIcd
WstvaA7+jODzDmPpIDQocfSRgDn0EG6z7KOFoTrwWdIHDSwOOOXGjqvudNW3zEjc
2R3UdgwLVqMwNrsY3TID358YVIWWadtpBUa6DKKKrNGGZUrsAzsXQJfUUPonweuc
KvHJA6X1i+FcrBni8ZI4i6AhtZ3/3sIwKaXRxhIdpGoCEbAZLPGb5cxOhZqfnzny
mvwEehLa34ehg1CSl/zj4gLHRRC0lL25qxhEAOqKze6T3fjq0bet1wghR30kpBfr
bpmGawMyDiGzjPaTeYKzPbS8zswv+ojLeskqFnaGn1t3PQvy4+Z4Uzm+xccUjFYN
fjoEc23KlIo2fe+LqCANiA8JAnJdkGUMhiUp7qoqT/0+NQkgHxqv6GnH/O8KflhB
+zbACHBQwm7yLS/nFtRMUL1efE6b9wQIKOImzOX6CnxhXYsdGHp/J3Ss/tc1P+LY
aFJ38a9yIdf7DAbvhrsXtJzJ1NctDUkRg0KjiBh/4EAJ9x8EDxleYXzcRBtnFB9f
mDkKZVsmhA17H664lIaWobtytX+w/fJA5BdmyZq5bbK4iRZQo3glqw2uwkhiJBlT
N2nQrj4Yal0wz/YwzjxkFUEZkRZ9gQNLPTvlSVYZgtBHzuF7F0/z8FFprGVmn9ya
fLlg8x5rObywRB8dh78jn1PGmA9kFwmCU7N/1NdZq2Fe5UwDwnOBPPdtrcpRjcn8
iLkFGbHgvW8AL/CC4+JDQTapurRUpZnSEjdOh6Ptq7xoJPC1ntT5lMqiup9KptJx
svDKBjsJcu/+nSgKI2pAvSw194wI6Xu92Pq1tvVRHTArUxFNuTISijIMKMf3t43g
k0E0jS0ehYRIGeYgLT/fQ3xAlGOrZRXJEG2J1AX4N4G4vz/opoyFUR0EJ7PQm/7m
RZwRMu0glHlUdaf1jJw4AOnZzdSmTPA5h7HJEvCt+QWAd//qQB9MiqOdbmkv+vzI
IAk7YxbrRLY6ASij2MgFUhT7RBDZUBlFGHVCey5C69sodHSiqZvfPqYchDiH7xtR
qzAZdQKbMnP2u2Htd5OBHTJa0/tekbYSKh1F5N4kvypZHywqpqBX90lvgQo/QrNZ
VsBAbQ79cINxtZZyK91v20pDYNXn4f7p+jULaQEY3KOlSN5vVXu5ypUSVpjM0RQm
NWe8iGRLvY9S1xRmL42Z4Cd+e6kIY4D83JDD5qqeK7yEeJ9BSHdchEoTPdkPiAww
V9fPCyaxY9VTfVM+CTdDi42awM5QRvI0b5sH3rkmfUB1NTTtsOxJOayYLIXfgq1j
NkxoeYtIk/6bGImbWrj0RAaA0hT7Uz+TXJi0HiZSjd5rTsUWCuxEUFvEGCL7TKYC
bcfklJax5+a3VBC3m0v0LjiH6Ix7OVqyALBSoHuk6zxl8P0uBo5ynLMFX2A3YOic
Uky5AEOh8bDNcdt/reWESOXcouoEzZqMy5W5ydepYeOivVyx3YylNjyiBepX1JbE
9nk4fMWInFpfv++uiAfnJ0acAeoIoDoKkow0vdj2nytaM45xhZTvr6LDKdxpvx8H
e4lNJOHmZQj17jVgdgTRXlVO+jOrwGaxvs/P691zYBtUD0R/3z3gQEL/b0D7VqT1
CNa34Cvq2shuWgvDQ78mYwAWb+Cwlf+8UoqqBelhaOOi3+WqbkS3f0OFb0XMoyX6
VMNgNhokOgABfH4QsAqLOdo+ceW6jl8RpZzTteknP6xl5MB71q2hNBsouUvIaDtw
oHEJhhENglzu2Sh12jrsE/aeyAg+MJld7kvX7qj9ARYKSvo4OW/Suzin8mgm1bbm
dURLLnNPTuRCTx3O9uqhXGmwEZ95qxHEQCG9Uby0kIoEa2aYyfepMgvHIiACHya3
Xhi+ay92HRoOZZ8HcclRM+NtwPjoddmH3tMdI5pL/kbFA3BGBxSTHtVYg+3fKW2P
RNMVvc6l+PQNiKx67AxdOKQaQz63xedhoe0Lv2kTRTQIAk+yFwdx0W71h39r8ZjM
V6ve6MkeSCP89mY2pxx4bcn+nGNUK/i64FS5VMP/QFu6byjc3FW+aQBsXfnIC5Sw
Jw/9ByE+KKlUzkcYGoo4B6fp1dKXW5NKOGG4mE0jU8EE5XXG5ikLu/ut6B5nvFQV
phWyDqjCNT2qdnlupOVH5PrYieFgI0tr+oN/trQiTHrIMvY1rBWNhObMYKEinp8A
1NJrJmcSq8sqoE2scUjfTliiMbgeSymnTj0xEZeEWCew046VyXqWFktSuOrq4qZc
MGsxuKZ94vUktDsYAkVabLL2uTMXWc+SPVyUowBAYISKEHfo7IcGNvLkIO+ImOxB
0ZmGVBSqYsfg0+8EU17ctO5ApZla3Xn+ck1fRTqZ9id6ZYRFTgapN58j+sVurAka
7szhDt+utSLfs6S4Y3wHfshqSJX46XNrb7cpbSkSHNXgrimvwKsN8cCaiJ7AvnC3
pFSQWX5sLHFLAkXJTu1OBDe4m7L6t9EAtdh1se+ql9dkovew1O9lVkxw8riIfUfN
CsDrO0cteO6RSBoOH/6oXCYtJXrLhRT9hp4UMz49OckRRZpiXqQpDNtRSKbzXKn8
KOffBFnJptYZkcDNE5swQ7BouNwlrIrFUHI0P5hoqL+pP/nkiiLxFowVK6ei5r54
sKP4sgfeq5dDx9UM1G0SxypfJT+cwi8ScyisoNScN+JO+r82G+zjkCtme8A41cRv
eyoFDgi/P2ZNeaLFEIACyTKRTR2fsYNmJrRIhIbjTR3HfIjStH/TZz94LDaDDkrh
qCu1dfcmvnW5YUadxZWqwyofdSmm1xw2Xq9v4jb51V1dM+vMZwZug6jl+wCzJH+O
XUxN9BSVA9K8kU0EROqt0RhLGAf5VP/140ofddBKiqW9zbCNIpsXEo5ELUSEyNM4
R7AiDBt/90MmagnQJiIXnmE+vvrLYjFOLHQqndNKsui5++AcjxJcwezP0dfTH7e3
amfCdl7vU7ATP31JPzfVbwnEs8vugXwdwINvvjix1hK2jbY3mIMCk73QGJb+/W8n
xknxKPqKAq8jxZAG7B1ccklXeVYv7kN+uhAufgxR+8C/Hah+qbWTJnJcENZq+2vd
u0z3VJy8f0ZzI9Cy5qROS9IDlHfdZr4SiPcWmNURmqxXrFggS5yrgz4sbsWRrM2Z
e3ct+YGoLDf9jAthh+fwICB3xRIXg7/9SyocK3agr1L1dNaR1vWCNLZDhfGG+MBI
2RRY28gDnKLaSxz6dDAAl6FQjG/L/ffn0mobPVs+Kb5SQDooTs6NN4rIRvOx+Ta/
CgdjbHa7YVZ2Y1zDpEhJYe8rLFr7z63C5JlrNZvtaJJbkcFTryeBkMXmDmdaIks4
hNuujTwTil9ty3n0yISayqvgQ9kYVWv9M4TfozzjPMndfpfUcHi9k20obRXiZMp3
H7WvF/Thv1EaJwUkPVeo2ZI/KgScGjvE48dod3Zd8sWmFEaFgrJCGJVYjotDpPVS
OAjnEHj4tU+wfsGhoV8CZylpT795v9H5XClJuSEFyVk3ubUXqNBK7Fm7c+11xLYI
Nbx35+31aRR2bTvamASE9lsAUZRXIk+TIvYTLBIE6hHqRi9tjbyYKjpx9uzXISZP
jgxcJq1AiCxJt9NItmQTg/WZ4p4k9oHc061cqnT8+mtU8cIPZJKo/sfQBWzeuvy6
FEcXr4yUgeD2CmGmqqym5E2kavyw+hLprpHPT2qoR8diQDu7sA5PwRe9cFxpPI/2
+nO/qAS9kQqYyQPPcRTMT3ZEnlFfH/o/ks4zQu8fHngDg6btV35EfBMXq8v4Y9hz
U0dxgRqE/4hIUYgHfw8HcRbCszHyKRDVoxyr5SOrLTGbRFbb+VDobbS6Wjb0nj3g
OYWNJ+tbTlnt+ojcc2yrk1oOsWmiq5uwzgYi3/DqYOQpnYrAfWp/d8sh3KuWENeW
kPW2tvG/3QLhKVqcjn3Tc8ebuDwg1Jkmu1k8gKoQpUYM4tphVgU+cQ953IXB44IG
BrZJrBnmtFjHQnV32Bek+Kiq3hyIE6MyilC6i2EzxSkmQ0qoY9rTeZjqdGSaroZh
GHNCpbH1KTrYmWgRZWjNF2m3oujcNmaBdXEhVMKffhz+Lai84nWml559+lOr2iNi
tVzhZa/lUmkJBT4wwS7spfANTcBPPwAiskEj/xogYmxcRzYUAgzEwIhMd5ILhGok
ApJ2lEvAtBSWbRj2e59HywTmjOVYxkO78cBq+leyJDswaJJ8FMleyoM6hyLK0T3n
NmK+O9eFlVQ5QwHibq2ufJDJQiX20QuMB96ikGGqwyHFC/XY4cv0RrWAhSTut5aO
2ahSbLXQ6SfSPrCeZeli3xJzXXm7XC6Q+7/pMK9spsmxz+VCXjE9E75Wfe2ROr8+
MY8qwQxQ3c6QtLz5yatdhXA/YvQPUIvXAl2QWxuhuz8Dsgmcn+HMtNf1BDsljvdS
mSM7um1vQYTYmSmBrIEBoqJMo5GcoNR5dTHL7Wmk45Dj0RfjUbHy7XPu11rOGtTQ
VdK/GfrzC9ncyx7n9TeiOPU1VSOJJL1LP8bHIWXJJOglWrK/cIBoyc1xeZv/WrbE
NlaYg30lF4Fe3uP0C1sPqqTIvLT+UYFRmMqoRhzLdt7My6mV1fsWqOHXbNFS/7WI
mmhzyAtZYWYJjqQMRlgP8aLTy9kjSmCIpnrw1xMl/cwchf8Xu6M3YfchDAf9tbqp
sL63sBL9R9Tj5JCMHUtE7A4lhl9SN12Tktaxmcfby6nbV0U15aAB8jzsIMosWuYK
4dn0m10JkDUmleN/EhoKS/yn0OSvXpBzraCYoGwWMKcrAc4Puasup+uyaPgY405y
22fcJlNDh9W5ydxdkJZyRNRtpvndPp/Pz3cAIWU9qjel0ZOvoEc1jMIKmMZjUdBq
J2iB6h3t4PL1w8Upr2FkEz3Afr7PkBc4wxJvUc4/yJXlyNYhp5l1YNHNN3jTiQHE
nUgRImLA+TKlq9M/63vez1nenCjxSsja9jL//DFilQ8zumbKb9hmTK9Jp45Egfjy
JnIw1Qt7uAdDLSunR4Fql19u7moK5H8vF99pRYR8P+L36zDBf2/OCNmYeufqFhZ1
hh3uYMoGVR6MMV9K5mIdW3ZULMnk/g6Og6CODTsqV6N+Pll3/KX2VQX5igW+FqQx
ANwtGcIKZfsZ4+PYr9Fyg3pblwrX8Utelhy+Q2uijlxrAX1tZWegRB/HsBFU6Uto
KGSS8Bk0Ed8iDQe5HQJlyVk2XoLj6bSLHqxa1Pbud24N2WJzgkLuWERc2I2nMH4b
pmhoYKAWzywu6yXbxc4VkqS36XvN4RXct66BYbb8gO0dg6bwpjXz5nfAP0y55S13
yUQ62P/CNZ217pzY0x++Gh70CkkZdPpGNricnYKq2YbkCOdJE7YOzHqzR8kgs5tV
dLXCs+eCtmrRIoS7oRiZGa5wSuVhp7+dmqbgqP0kft/frv3Mq4iZSq2kb+iXFsuk
MNS3ZMmo/7nkyJ3hgnODW0rXsYrOVq9pbhiHaXvpwR9QMTpzDHNRYF8zc0FEf0m3
/bvKyG0SwvLKFPjKnx1jy9KLcbhHnebn3qD7e1C3TRcupg9UqiCpV/3mvaMXdMtV
pikHbYBFADzUiE44xIX8u6SUqng3Uw6RWUTOegG7cs2G61wpOk79DlZrHO7dHi6a
n2V7JeMNt0R7zHGcI1ozgpGQ7p2zEj4IvPPveIgRYTpM/kR8IAOytycRV/WTnJQo
BKbAWTderWOZ/SgRsTIjal1p+nOonvWHVe4cfDSz2P2InN1I1pGoJQeU6pnPyhJU
lrL6wkQWbo3i2m6G5SjV79sNDFlmdsWmNV1MwOG6crhw72Pjt9CTW+W1hoge2+e3
HXqbbU4PB+0M/8Kh2B7ZT0FkxMp4Zp+KM/qKuiuers+DwNozUUtd1OcAcOk094G+
fV3CB1HFowGovsj0/3xurwZnqpv6LVX7BGyY9+F9r33Hw7dNJ8EdEN351mINP5gx
5ILv2R+gcht7SQ+mHf2iX1dR1MGWIHpXlxXhtIo+nYTxx/Maby5YdRjuLwjMXuc7
8QzLDIpgUPCH1yZFOF/SExpmwtNd9uOVMM3HJ2z0ZrSk1J145G7Hobr5zJaRDsbk
DQ6w8jTErY/ZeZFPaX3nyVempWuNwVFYef88q8XpzuppNnfjiBWwvcp0LZZ5l8ui
k0AXCSdgvjAkEC2JhlSbYHhnbqnN6+j0Ij7jtzuLh+YWX89O6ptwNuf15nL8LSFP
aXoyEAxaQLdtIXrjNTRyrIrTiItE/1WFimPdHDab9p4EvbtB51JHVn5fYniBwxmG
hxVcvkyQ0vt1SMwgjk5DWFHEdjAbJoRAVmNK+mQoJpd/u3YaIrfElrdJHod8zYhq
uaaZ6/+YdX3vY4diaHdLxzVgWFD+umWvSmnxSik/rJ5DrWIsBJ6hWxYjhnzbpvIW
5qVD628aKjbb74Wd3oZL4EJ/HueR9XXoFnBhYK7PRiWhqRrAvqFU8dNw3VBCTQZc
0g4M4vNpied0IUsMaWoKxrtW4gM9N16EYKNUnvqmamgKtnc9z+9sWbonATPR9H9l
aOlaap/6Pfh18DQOv5XY5TDvidbT5Db67gVOAP3PxzwX78Oi2huG+qT7ih/SVyHH
dUrql0lKan1F47IQZAGToEYQtZ3oSpIGOHkLYlAeciAaEdo1cAbARVkUAONC4of+
kC25wa32Te659g0WWYBoHFGNwDOrxgPm7cjRjoo6jDjowGl51IGAiclJZpcZ8beN
D/cpUo1bpzFPwMsA2+8j9GQYpcUfJs5kszwJLPxygQQYWw3IxAzRSSTpP7XPljJ1
YHi5MhHx0Pf8mnKk1mGRdgkmIjkowqtgqTAYFaXeEk1mvBM2g8yW3VYvkyHFxk3r
fXIYaCg4ojUPaWTz0ilIs4D3Ur8n6mLeJ7fmKiV0Ivu72L15+hn6rIs1KkEOZE9K
WbmksQUsCVG46DKVd58HoYi/ulArU8jIwSi7++55fYdRsM4bNjSms5CjvtSgE9n5
KUe0FQoT3wsIAxrQzJ5hHc1yfYEllfrgjb2WtBm/WC7hwQtTEdTZCwD3Kx1GlG0h
IrSmfCXm85+zsjnQhg7nmW+6/M6Urv6FJB1MUuahAu46Ro7QXPnxU244gaf5/jBX
FZo19SfKj0oqGmiGX1OOvKBVw/X6VFXKXkoqboRhZzsKU4OYWc/ZIaYZMmBzeJI/
6/tUwB0uJMEebsd+ths8WNeavdbnM5+DflAdT4y5gcy/ECKps3+mIvjryiXXeA7G
80C7d1THJ7BDT/GUGkH/uTTuq3j2RGh9IZtFoBwuX8G/D6LCuwK68D7XJhka55PO
V0vlKWu5nBVd+NPJte0rimr5jhEHjwuY3BNCVGrv+++G1iUjCJU572EQcHnYYS4O
VsLPhHeJEj9J4nreDP0QDHQmGREs/TYp26DF/8q7jwqStuBJaf4LpZmNKSlzb62/
EjBY93Y/P1iMRNBUU70dfYmPNC+gjGzYZXVPa5KakDNrTU4D03v6zjIW6dV5KC9+
LKL9f5Wi59+p90QexDrsw0RGADr63l+ibyBzmhry3sfjQSDJeJ9hE7HKc+YxfRw0
cUTK91zw3iR+KpuhTr66p5qIXET1yyHTcC6E7YL3IhzaF8kojS5wKObq6V9JL8HZ
DZXr2fRE7IZqufNtlLGnlR2X5Y+ssunElMnMjqkAosjU4SOKfaRri0N83Ty6YC4X
U2DO+7+2wzsUVoca5SlGCznVVeuVbW8YIeej7OAQabqnitsYROVS3cr5efNXVprA
RnU23LAv4Xru4HsDCnqUZBQojs/uySuV9n40+KQg7UBmsq8A9F8JHMNrfmh2mQoK
YTLTc5BSXN0XyZg/rnNDqugBMkTzIJQ9lnP+qfeBOoYARRfJqwoFdzG0VI4IwDWr
DzZPubcWehBrxCb2ZLuf+S8snhRRB/f9+zR9VNr8oSrSsIyEJVxQSIY81Q9CMqVC
sX9wsWBONbXHcRyfJ7hgbjydxhVzt7GrtuJOPmUh+oUeqqh7MjdGW5MgsscbBMJQ
gHmj9f/SEZUR5rfpeuZYi5jMpU2xWGBnP+w2BkQ3tWYMfxGz13Pbi7yzTc6iSYbF
oPcLZknHHR6vdzkZzknvIehtGdJtbz/lWPANI4oT5ga346gSZm2EICFm1oyL5ceu
laDdfJ+fDT0EZSsMELwvgInq3POzNvAhVnSZsyfoxQzG3bq7E0etc+EEgC67GPgb
COHn4k4EdcDDrG75T68jt5sofeyt31gsmk2jgCoCF0h3pCON/7Sks2dI9aPWaoEp
9PFUZ17Hy1l48CdgU0BzWgIrZVcSDU9XE/phq5NNd6rDQO8E+ffqsm/rkLBjRlG0
Iy4uMINimBKsXhVLIwThxuObkDinq6R2HUq77ul2dl1mYQMuBumXjmaxu31kSDSu
VC35ut3mg9HSVbOJdMzU0OksNCL8ZIbWVVlidVc26W7skZIUAckFeCxuHO2M0cQ4
5aEXQpBexF207cE0L8UQ+i4fKqL0e/diSkKs/M5kdnEa3D/W4jLH4AWyiTQtavpm
7PLWXcWFMVv9Yks0kGJim5N7oUg+L65Ff3WDdP4cwNe2lsPkQ9gsv5N37m1TLPlp
Lx0E5tUqIbuzofYawVGxZD7j3Z8Ba4TxP8rE85j9DAALQR1owmWTNYCzQ9VF4vWE
xhLMFwat29MEs8dUk4cu1XM2wO1p9I6cqd9y6yWz72uyG2RqUh2qbLNgYPXfH/m4
SeTvP6JjDuSryYW5EepWg3oP9zEJO7e8ilj/N5r1l3ukDHd2ddPyd1GHdiojqvid
9QQiE0GlO4vmMsgOlCHd+n/yMuFhOfTZS0nWUo02UK0X09IDemQsxDeQerpODnZq
oRxCYQ+5AHgCaq3+er8XbTs16hvXHVmUt8zGrMN3xyvdpQIrgjHGHDuLWgfyDp6e
XTEfqXgJq41kg2L0oiYCjeS/Lg66ELDg0GY1Qw1cPWboQ9+ujEvKtzfE6lMCKrvF
wMLDTQVvnZXHfVqlbb1dxTX/DsV05uYh7mc6zSwiin9OeXRxuqyHqCNlF7IHiKVH
d2oDbvyNxUgQZcHhPYfnWduvWFooL7stlC7PybLpdgqI+4vW+LiZkwQ2vdq38Ix4
Zkhe35FaplcaWuiWvi9g6ARzRKD4CBNN8YYo19RODwVVJfAu9+wRG+p1L/cuBcip
Qhku8C3XWFCPc/j/70nsGOM8Le3hZxFzBQW+FeHaPGIrLzbzuhgq1pntMCECPgOT
Jr3GbVpmkBek+9rlRJRS2siiUzh0GokUr8pZoIA2dL4ea7tXqYCBjK2hPx57b5sj
UiajznEY9FR9sBKpeIko73Eao+LjqOG4h7qpTbBdzs3k/NBGzh8n1/+9ZfZyy6UK
iMh9Pt+NOLa0KyQjGYu1hAsSq3drS4OYdICULruT/1OeL4C1a35z/d56Zr5fRBnn
gwbg5/feuzAtlsCbGFWYlyeJalE+YwA3JjVxnPRp2yzKkxprbC3yLZqPtK5/Oow+
1dfn9tveq8He17KyjCpZZ2KgiKANYcXg3UAtvsq1QtbVAJ65QiVx/uSP7bZtXdRy
lkD2pCcGUGJ1MPPz5AZZScCYoUUqNW9GwpqR1zIN/PXyqJ5MiLp7qkowr5cfh7+1
18tLOZE2A7/gwh3xycH/M5qwIWLVS+1XfL3khNrEB5E5U3U4VddWqKJ71/V1GzgO
ctwTBxDhHrlYa8TRQyI8oWg0vFXRCgCR0qkO674xgq8nNGoCGMnpDil3DEsYdFtr
S1NmdHcsN+aGDZCKDzqW7fVvneRxWa+DNl7ouBfSomt3HmVqAFQDtbVnXLxDWVlu
HnAPlS9OJ0fjGL0KSCty1j1W8sxNbt++ZrWTExu8lvXGIFsJnybaPX4GGjGDp3ru
4Yd8hi2EHL/POSGrgljZPfH5ovO5kQYdNiwebHkmUIuRnlKgYuaSRfUIVgd0Tszj
ypWwUWyXa+3zZWHIbSzfdJzy+DGwTg0idxWFqg4v4lo5LkzydRwwVEGGSOcRk5sw
nei5xPGxWuyPcuCRM+Y6YCoIqRjSSowPIkJmN6t5+h0vxN1cTFqdyV3/x0bTu6bC
Zuf8AItoxqPNt3rPPrm/kBJfSnT2lKFlF+0cXaUvwLuV8J/e3jM01JF7ZNusLZws
CYm3+S1mp8W1rntCX6nDqJtvIJJwMQ7DoGLbeK2Wn6nPfVQ412PObEH2Zi5EsZyj
JRzX2EpMnslYtjLU0ggO/pzJQ3Pg1i6B5QHexBdMR9NcEq4tZO/7WM7WzIZ9u/pn
fnxUNlzcZ85RxY4VX+zMHqw66Mu3JImzGhaxcffYNuRt3d1JwwrL4wbl/G1FO8fJ
JBEEL9fh+U///1jyeH8oZ7tF7IgV21hsAB2BlsCLHiM39qa+BtLZGLd7TiUK0nHi
wp+RwV4a1eiEE+R6DXZL4z8R88tlZa/NbXxaXdIH3cIDidsBsVpmg6J8YoIw4z9G
ebmjwDeW2O51A9ToQ+ititVg1I9/3yIGJQ760uriqGn6907H9X1c17EzzXpmEqr9
igxzEFsLh95CD+OI3cVUAKPkR+dHPmh65gmYUSBKjZkOd8VrW86Pfjrg70hI/XSD
PD0yxzFfKNwci7JSnH+Y0oUi5rmuqCfXabLOpW+eAEf+nV2xmoV2p9qzMjwj8Km8
hDUyShhT56/pDEfc2s+Lz1lxwKz3/hGgupWlciyfoxNBKTyt8m4lDyDCwm3RzxrE
7rkCRAglBubc/79zkT2JdgTgaZmdoeS93CknD7Dz+gQSFddz+TBj4lU5dgl8lXCM
KEd7bw2Jnf8dLW0Wyz8y08DKioCweYDNJvYzl0/kyobh80aPU5sGJbZ/Anf7EyCu
7vThCG17Ej5UkDOmoId1LHqGB+z4y0YJk/jyI6uLM6EALYRP1juIUxYac4uN1hU0
Jlo++aI52A487eBZ0GMeSbuKrDAUbouFKOpEKtPEqBVaRksdYrwI6UsZeqm3vW5F
kZYncnk0qW6GndSD+BELLAITwLz8d6rOD3+mwEbPuUkmbU6ss+Tni5y6Ax7BejPJ
hotWZtVMbjxPX2Enu9FcfptVNlvh0uaMgfTLlFUaitboVDkVqXI4W1zMp+4KBcah
2MKLssdyaPHnwHSbH1AjB8tFDBJSdR0bkKba6wTg+Rt+prdLfvU/UIdHc04WxbAc
1cCcbo2uoL3a/nKqkdZ2l1biscLavHV3fIR46ETAVvytUknOciLMb+JZSpbPlOvt
qOufQ6CVDKm19B4iBaBpNRLcOMzPhIL8VBeKzmCXrTQ31whJm1yPCLfe8RJaekCc
QRVVS4h5RdNsJTcIe7cSQJ30yvF77qnN1ErHKo9tGqJV1caSxVTV4jzdMN+ONDuF
qGuOSzxDkPc1AWRf+jZqFJq0bS7sm2M0s2Ct8xM/va5xxdv2TIss8M2sI9WHsx+H
lJQMugLooFw7OA5bl0xTro/RyJ/LLYUiWyVL+F8gWPl5KGT2Ii1qr2cI1oS4jph2
I7pxzfh2wCGWj6Sg3WY/W0BCNZcSh0TplcWGPtsFIbRVgLm7jo1QElGGD8sXA+CE
5cGDHHNUjQpo07Cd3xtAo8J5TbEU6oWR0vdrqQV3fiRpoiHF0TAb2Eqa7QS24okq
M9e7h4EN+D19OTC5sC/cXtuVakluD5+8IVdjMo+wDQNeHlxFdc9qqz+LFi9zNiph
ZAgbPFRFARth+pyCNJE2CUHJckAWeRfucHomdxbpDGqBzsSfOCu387TOvIU/0mas
NtbsYN8a1HFpeh/9E0xrdtazDgrsrn9u2QpCGdFYDrLIwtwH2jV7rv4bA8ITj9DF
2u3gXqsIIvmDJkJomJPBYLl+V91pQ4PcYD00EDwQG5MbMGKPZN3hKp4RLmUeXCrg
MZ/qu8fY3vCslcjQ+KHs4/jrL7Kx/b63A8nEaTCfQkUPCKDMjQP4tgoCB4OmngaL
JyiFlDia6g23/bbzJAsuoOE2CxVktrgI8/RLWr2pMhCQCItMIFTN5/Fzv5sPSSgp
PG8uXvwQxRSHRt0GZ3ilzT1yGJ37GZmBlJhElqYhhRxx6R8ymyAS131BHdX/OXKw
QYNBwMWA7UAB4MwGWkLXnhgZzS+OOSsPG/OHLRyOfd6mY48BNE6UFlgUUYhEJnzI
qPA2V39g2openIwhsjiR0JmvbPfOX3CGGH3bLGlZVQtKyXr3JsBpP+aceczjYMf6
dZbekbKcE6lecQ/lBWxL6bR/YxCWdi5pnLMzgKONrxwxYObp3FdFqtbPhvtmRg8+
vdSN6Q3Xt2RXmcvvC9Bi6pKR1mX+H8FStC/3EC3g2ALjogiqp+VFxH4IW4KOrcy5
wAKTFd0f/ypt3SQzArRXjuCiRwpbZXtyzsrz8NsKEvLu+0SkFRUxO8aOlnVAsMWX
UwuyGK0MmA/4fL5KO65KNn7CwlIKsiObJ5V7MQL0Yy1Ox3KUAOZtXL4Q7c2GNPr/
/aRG9ARGTvmF1hQVAAzwCf3EcXTOiNMT1tYlZfgui61DmB0B7K+ZfnHcHJAoBYMH
kyKY5X0/J49tNGJrxRgqnrgAfHoT0xoKjC8n34DUxrjXgAnpWHr4IKGlGfbbLXNP
lHAi24cm8g9vcprHhwak/2OIUYv78v2R9pNSRJOb3qB1VvsblhvA9O+K7+yM6nGC
V54islLe95Dg5jinuP4vldl7GpymzzTiZ72JDHYKDig9xQc4AXoXoDFfJFbpS3xr
VCpm1Pe00DFEHZaRsP5L1zQPE0BQXI8JxmNss4FlEb3zHMVXCpvJnvooOhM5e/py
nWSgBxoSam4GhCN3PK5ac3YPtIREhhaSZPOyqafriF7IfoPj+kn3LcX3vwr52MR/
ooz1z20cCVauR7csJsuDUAIDEhs24tmOUd2YFVu9dDbZ03cyDXZG295OlVEhcnBJ
GqYUm/r58TBHcAFe/HPeBiVMtBovTunska9mwkbqX5W/r0ZENZM5DcbL6qtMWpuJ
vV/7zy9zTf2iXM+sJvduhK7N+5g2p1tchlJUWneM3R3TIyl/eX3vlOckUvGHbupX
fobtOEgIOFXckRw+YSeS2GLU/sq61BErrmRQ6VKuLcnMCYES5zrsvQubcFRhOQT9
0e5aHvBW8rmjdju/wZ90sHBCCGvqFl2Li+ZzEeWooKgdx2KitcbI2Suhs78A1d4P
jt326M8HpxAoEKSbufwkY9pCpB+Gvl56hA9s+eC0dUYnQg3nmPj8fDkDW6cSXxaB
X+KFR49GM8RYYw8sHGCXET4Trb7xCK7+4ctfTIhGhXmBfKwEPRX6OmOzqEy6oaK7
yIy6i+4N7Ptu8PeGrPLY1tgJ+x6Mqx94dKAwESeDYOnpsDgs+Gt8gKHrWmuYv2VZ
xsF+geoC3nS6Vkxu/uKbX7UXI6GzZlrYqJ8ATxTCkNlJIRMEur1/xz1eKmvtNLCJ
giFEmspV0BiJit2uAf6fzb8JKF46p8kCe7e1CWOa19VC420M12gJtorTg3fGqjrV
cVb24sg38bOsbZuLyjHsrbL/kFZ2cVPcvRgI7CVdP69azyFFE8DsVFzv1DE5/mE6
da/8/j1S+unt7mK4Py2mxsVqiWWcdBpjuPTrT9i/85uzSU/64mDUgL5wKgKHuH6M
Sym4TDxciIKyHroOQ3mbpcgphBvJz/zwgqUXnCRD6TQhsfosHu2tXNPbtdO4+anQ
TYj55E/880r2nlUbEGgUGotqr0FdjZ+V5bZtgVgUzv089PjdDPEaSwMFDQGnzz2U
UcmLac230XLyCI+9onGyEAwa6XD4U/Jv8GQtrFOcOo2Y2y4DOpOcTWFL+JyAWYhv
xX6S5MCh4On9CQuBHibGmDv5lm5pdDbA1UVXMUoUEGM3aT6Gjjq5EysV7GhZ4W3V
VBxaIoAh1ldx4Gj/zg2TD0kbaKx1oIXByTpCxccpdW5BbBERg/pCnOfNHqztLtCy
b2LSvvo/E96Pn1ZJgwlJuJfTx8Z4QbQN7ga8tksNb7Hmud2cvGmpTgdmPZrOX43g
Acj5Zfkn00stUHI5yOwqqByfmgYnLeCU8Eroxo1nXBPKyikkABdlY+JjCgKxaR3V
5AkjLgBnzM8btIN1U7w2GuWstNN24TgbMQAlykI4PlGMHMmzjhRq6SuOyoclpl7s
howP2jWJ3OX7ECyP16+wbsHI8ORKI6fQCSebxlQ13iVnydnUkkkG3DVon+x8EIta
7e4y3kTp4Y2fwPUAZWqWGh5F3Ng9FIXVrrAnNUzH7C+PB0XcQ7xpCrHdW8/3Hj8b
ZAJB18QYeWf4vaySMZDrsv1fo+FdiYf5DwHd7dZ1V6a9L1xZa+y4tMnA+YzmuJvw
Io8N2h1DQFwX93XaFBVKmK6jnpE3lIia84XRTouSQXtD+ry2u0epAFX1asxzzKuh
ydDwkKBYOQehX+fITJgW792ivg9HIxU3M0dirPlUYeL55rHRL/BalrWcNjxaSLVq
NouB7GBUUFfXr71ZXFTFInahyUQfkEB9U6HfgDpCqxU6FS8GnhyowygPnEEAPCoW
mzM6YwbGEmP97/eGpTEgYkYz2hGQ5U5L7s+SRAemaJ3nHJbzf9XkWpu3PKtS20AQ
3q4h3i8UAlwaldtAVQ2qWSLyz1/kXqV7+39q0/xUhCjqBbpp01+G731l/6m1U2ST
8XhRBc8U9si5Ndk1VA142xL0mP2Ac+jMzVuptB5o/JEH7T4SPI4oaxXjdIJPVpQE
TAHn6gVX1yutEr1PNU5zND0GU6Tz1qxsnjJKzxyvblN7antUcTmX5ygifSmWmodf
2a4m0IjShweDoFDvHc2tF3rPt2bzxiJ/WBS4bkfBKUbC7XtCXiszUzbYqMwevKGL
pa6KvHWZjHZt1NJnEkPbdjsP81RS81vBHIdoMXAzr61hYLRLqKwKfOrq/Us5K5tN
T3TnpbBf6Ws4W+Kr+MSHQ/7vkVBK6MyRFZSnOkhZretl8GOKc19QgKDILl+9XVxw
LKBYo6inZcJwzJ5A7/IuIF9pJBf5Dwn3suN87Y90pKYpNjaRvdFbjyaXrliy3AnV
wb5/XGgJ8tx7mvvRe22Z9rOB0H8a8jmgNeLwsXdhid6LOKQNO+MCeU1QQMub7QT8
SILio7t8wB0eajyiMFdXtd+cG5hVO4+xB9s2NERszFR66zz5pHe66NRa6a32djft
RyGd6F13rdO32ecW9v+MOaaaFxYjpsL3RejnjS/T2kab24Sgu21AJRByvq/iavWU
gpK2HzkqYYG7fEGq275k0bYlFxy+mjOCBNd/w4QuNYJkAM6uIEO90MCGKHgkuufn
mOQ9aiJR2eNcwgvXWvotid3y9FXtdFcXd0mUsM06HADOEhckhPiTSWDIRgBVeO8q
sGeQRtm9nlSXB2hsmXtueWJUdJMSo5ydgZFViDyE3iQVd0jmnRg0YQmX0zqMB78h
o4sjxFQxzUF0L6y29Z1YpGJAaI1XknNLjfFbPKg88UswXQs7NxJPJO5IJoOoyPvQ
rgrp130NDX5mtEfBlUeBAdQD1SJiYy8aYKBBGkuK8KG3XDb+iQrQoe1ty+78PMPB
RuUAdRktnSdVB1664R9uTbp/IFX/WERnY/9S8zL47Oc=
`pragma protect end_protected
