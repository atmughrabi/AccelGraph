// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dA4ggx/+hVm9Px0NGeS1QOZFSDxcQRpiOe/k6o5Wgd4xY11sY1IogwmKBLgwTHNH
XMYNGyM3WYZ+ruwqkPUGZ5TEfJOt0Avym3NrcZLasjxfv65PYDZlrz+PKLn2VLFy
Krq2ePmsa6C9t2ofTgt+DlJ7b1rqeC79Y2PliH5a7/o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5584)
61EgiFP+ys5cUQi9znAjkjzBtJgP0U53lYGCwoXuRXDHXqQ2QmVpt3a+tRwgyjZ3
+VgRcmwG2HRrEuEvpir3v76t3aKZiQJBwUCqu4gY4O0pbD6/OjiRS3LsrirU9MSX
jt4GFJNN5qSZNio4ZYj0cFBp5aFaC/TKAJDN0hHLM/+UXNJ6NSYjf4awtGM3GW5I
zgRkNdfqjEMA65g7mInVUqPpcXhlGau60OXQDjArI2ONwa6l4oCcaJDT2NZ2axC0
BYXev8FOVoa9lwvybVbPa0/+6YCs8hBdwMfgdGDFnbKcH6SUxBnhoDcz/x5sUqo3
a5TTONkpfiT4xatt7ed0Q3vwUA3pGzmnAH6K67an+5aChwm98fk3B3BJBFUFbiBH
5tKPjyYdhcapBRxtK87rtOA5Wee8L9pAEGZPAjA44U70jCXv8UhDDktsAna9gl5/
2edrMeRcCU3AQ0JAoycdfTkshpSClinNce46or7Pky5DIXmZK+iKQFj28l7OK6Xe
SlRv9piAnI0XWGkv0X1nvhV06UcWrgQrUE+Fp4VMKQfkX4tY5S7ShfNDgVK7PUEs
wAbFHVvyYxBZ8/my8/PgELyigGIRAwNux+aearw3Xy+zEM7geQhpiZJHI4xOeAW9
jbAfirV7TXGmDV121/AmBH/3Oic/GZTXGLLGbEFqOPCf6N80RnH5ujpia/mKnyyj
T1tPq9coQqwXeds2aziW3kL+tZLM3yuz8LI2qYZ+QsHuHonJZOoKlXKYkm2H4XXh
LfzNgruCor0YFoWYCR1ue0dsgwoJztludV18iSd4NFLViZIDr09SOGHoeO8sHiDH
x1PjVLO3dyMjLG/AZACaPbBzjDh6cUep5Jnh+Ge9t4GNXKbGA6irYDEyGh/eV1qb
w0xSkKzv/V01R7jU20dE01sbJ9jWNwID0qI1tdfehpmW2N21TVE9T9L4VQTxO9JQ
/ezjvQDAwwW3aCcnqZ6pEJHHLgxf4XCm0O1fuyZ7gqUuOt6yZCNwS6QYD2Co35Ix
rfx0WcneKZVj/YIg9tM2HfYyuuQVPIi5vUrHNHnKLcQybunTnl4CmzCOgWRzebeV
uAV4NwbEFOd4QrH8s1Um0Rb+IhU6bTsoLnCZEPBhu28O9dvirkOh9GjiMTaBDYNm
gRpuf+32hQMpB/fA3879K8Rr3AZIaeka0dnXyvZ/EQAtLJSzgRLoNMkftg8xgNu4
a98OZOUz9s0SVaZ5x0zytRIrqvIRxgtDTe3IuurIwk0dcdKpdcO55JK7/eUpC+IJ
ZH5txIn7tL49k0EjoTKX6W/ii34gGB8NzCEBTMldFpEUQIMZczSoakc5jDjnls4X
hMDxRkA/VTNVGxi6CORnQtQjHVyvXBLM9NRqkGbKvQxy2bCq8oo4MtL24Jadfd7i
gjxbg9mv/Z4hw0KxVAtuUdSV2re1e1YxCSFPJzAU1EI6J/KIQam23LVumD4UUxxI
RczP5ckMPOGYhn4gCroJQfNCXILUuTmhYFlovWs3y/dNPCoIMFYuQfcx0QfJaDUU
g8zMZwb1B2IuKOGxNergJDCwLxgECvBQzid7IUnlIgWQRYNRY429X47ByFiii/5o
KdSyS6bsUNMuoPrPmFa0Zql+NJWazvcOi/uf2ubz+1fl+O808heTXn3Q155CSc7F
HucgOt3CPMpIuVeCU7rgflx4lz+I8TiaTw77HUV+1QWPLxIK6ZJ6zj2V7FvJobZn
3KseSnlWmwEVPDu5eMpvQrTscF2WEkv1VNVGGWklxiU1nu0fqQtqFegdWx+/CMaZ
rsCdF98oFMKFkWmeO7lDu/qtpv5KBLUkxGp3u4R7DLTLXB116oJR6r6JHQ/fShFQ
MUoTu6zGgdQ9c59g9DVfSWeOYXVlDSPs3LWa1S/JUtH/gd9OSd5mfIgrcNtSUIzI
XBgDqe0EjSuXZa5NJuAyUAZBliwnH/kXP4IKju0afiMNV3u9oZQtazIZM81VCFNr
UY8WFAz160oncvtPc9UiqKychP/w9zXOgoAMRg4ZgaEYAoDmgPm9nyrwN6Nf6K6g
gYsdhQaGW5qBk+exAy/oIILjKUwMKehGoB/9OwCqIyx4K6f9bAe7S5JEkAYUQlp0
qN4Ao9HEPAYJAb8QyOr5zeelMF41nteGb8j6MHH8JPqLf9MOGWRhcPpJpz+viJdz
Mr/JQjG3c0pAjfl7OryxxWSbcvwHJKOCDL505GBv5m+J7KkTuDfkOFUT2LWefsVE
4t1VowRUr4Qm4jk6SjBCYIduT/WevXzMzckpXfvFMDw6/6LYfzU3ld4chipGtDzR
XJ8jfxsreQKzqvkJcDNdWa+460Syq/1cMzD/iHTVsVmPYX8ajokMnxX4e9JV5OyK
+x9nHmxCU8bDc51Gm8Pv9ImWksipjVvw4ni/4FzE5MxRgCErahrWul8mwxD6H8sI
oWmRNczZcdJkold4H62XD512eEf3/WO3h271B/0VAEvHsy14y/2/qe1azhnjxFVY
05mQNOPusrmNExtKoHibv14PwWk9t3vWnW+zpSYgazN+XLpkhhRHI6pg1IcJMa9C
5IrocDBpu3897NarLvjwTv6jJidOWwbqnE1/MOlhHvv69HHFrNyDfjTQNo4WhFjn
j8IP3Yyw3kiHlWrQpUCCi9rAgUsea3C7grJFvfPNcs/hlP9qdgifgcETjPiDaKDR
7DG2GQfkbu9nSHtSAB9Y/YN2Kyu4doYKtBSvycCcwQRL0DnrtzENwMw/OSZWyRl0
ERfrCnfrzmxX0gG3ANp3pxRuwZMFaL2OQ0MPEPBCADc5SFrlBorXac8OQsqd0WW8
dO4CQRqYeSkZfNYBApWgI4EnSsrkSKhWa840LWSGxkOTW+6Ncc+zYnQBcTzoKkWL
iYNApTzmhELN7P0Q+UtvzelLZIq9iRylGBqvZ671mMc7DKoLPEFNngACj6NVncUb
x6y4F6+2q3bL0052b3Y3rXChkqnRME3LV+9BUpGnJBbDRwxHKSwP+hrg4NxUVNWr
y8ag3/FYKBMEfLqYPC81hf/ynpGyOpwT2h3COyKoTtzz50o+tbLrMbvTGvWv2sqP
HxDe/Z41IogRXVseU7inMx2fRxo92LjiGY/u1XlWhIin6Unucd5RNI31DgKsxbu2
vEDNXylCklEksAi5iIaRVJ539xXvBrYovw9ggmIehBp3kLQxIs91Dn2dznyhuoFI
pUycwqI/CX3jnPHQ6OAzk5r0QzIQTa/dWhvM2lAhlvq9EYkDBcYDKyCzzAT7QeWe
Vta0yAxBI51fsZXoqVZRwCh0OqM0xFw976Gpzp73q1rqCRLcEAvLrrslDs2Mqisc
Q5iqzuClLbhnLcwmztq1uUUh7AHIWgryWP32aXSbdMiviKj/DsWqKU2BzQEFSl6S
MHVxBdLWFs+CHCb4Tgsa/RdH/YKwzVFX0hrGiuYSOCCdgPawyvGcx0++3aGfoI5D
rPhYwop3A8PNHVCA4TsVKEZ1muVU6v5kulRUOCUO91C5PnfUcR85EBDq9Ztv55b5
KpV7z4LLZtYjm/lR6ecyKX85t7g95o5XVi6Cire4jKn4Do0jM/LuygXl0turQYs7
2T7PXL2WB7yyLJQA3BrI4C6tLPDesZG1l1yg8PRanmm3ZUelE7J/hMyTrJlbWTdw
P9Bo8z5BP/ZX69ydPmunync3nk6uUo4pDPbjjWnJDDAJ/nEfovJKOTRPLzbDpuhJ
XZGV66WooHxwARM4h5sMK9Gtm0i+OxjETAhXGzp2ChjdXEKae2GZyU5SwE9e36CX
AAaeMvCBESGmH1SCSxoEw4Bc3e+44Y86ccNISeHrC15di+foEEjXlrc66ICwGf6v
swjuOCS0kUJ/+P4IESCD/4fAOiU5TYub/WOFvZCIE8J8JcRpzBNc467NSHdvWhar
ROkSIcwyg2ds8y2z3BHxep62i9jIcF20s3Ks+PUMW9bQwbK8cilzubuij3TrZx7W
5xo0u/D221kaYGWa1OhsO6S77mscoLpzFcjv9Y/PPT3tSkr1ZchmlJlGHWrklLPT
fBbs8UEJgjG6JUmli8+Jkl9z8hkWyxhoOMfBC9Y3Cp+bmPLChWiQsTbRXL0ZH+gK
l12mYg9lvGRNSR9U99NiqanzOAQuA+n2qAYdctObIIi1gpZAYVt4jCojKg8Yj+y0
shpX2pgQtbS0ZOinG+Jir+1uZ07tqyllNhmWtb6eZ3mi1itjV6TnmrCc9orHjaLm
QyyemJ1MiX2ho6Sr1nhISdpacb938sLaDHinE9jYaytWQjBmx784cfqh06QhacBx
RHZ+Orbbrr/55fq1oyXfKeMBL8kUIMcdjzxJu0fG9f727ZyzAfASpcvj6g5Ifcef
RFRer0bDVfb8IK5VMRg+glR80vfoMdmMzLEPOYW5u80QGQpacaoZJOxTLjUVr0aw
2IdztRWlt3ba4JXcWOKzijrtNdRAj9TrCuXDfTFOE4X6G6bwbxa8bKgitt+JnnSw
GS2mOqs2NLkexhrT99TFLq3ppxJTFPzN1ENFNmgdVBJW3IR2TX7snvrGtKeOrfoA
mkOh8y4itKy8uu0keteMwZUsb8xEyoXz140B0JyRVt3G7DT6Ya9zbx45QhZe9rPN
jYI0ZAE1iN8HT6qu0R+PmhSkMcL1FIia75r3BLhGNwqeCEA0GiXHxJ2yiooNFpUN
QOIH4Hib0l+aEJS0ft3sRiMrtRsVR63dtuC8pd9IHz8XUzfe6zNshAIW7VrbxeWb
IQY5xEHIUDius1bzqEz3peIjd+jNq0LDTekP2v9X63p4EaOdZL2HyTV9HyGD3SOf
rpmp9QjuwB8h+rQxSl06xY4vQcD+cjU4S903nMlgTHcphjfMwltZ45kZfiVsxh1n
pqxKXHAg4DT7A9cVzdGaff+mdEXyjQy2jOe0EE6cdzMXtfDDb5aPJJ3l1JoaxI5e
r/sXHRnvHWA28HtmwdAIazV4VSjXAyrd0ybNhV8DvHuxRL2ECZ0Djd1LeFM6aBJT
43YP92wghETERmO4ozN4vuGAEq3sz7Y0AnB9xpCixfHJQtt/AQK+9Mo5ZI5GY3sf
85R60mwNyzMOXjyX7FCG1KQdkHgJZQN2+fZtJ4nlFZpSeJllEarlXbZzTGASrJnY
T2HAv5IKuKNkQWmpikk3uGNl9SYXA2BkPJIMqzHyGYkHbdPyuLyvvvapsQJ8cZtd
NZnnbvTkT6FkbJf1eXehLvSD1LAzMyFS2JVGtGx8oIITbN4HPByjSzxba9Jd5CXX
vKj9KQV4iIICYtNGCXwnwPf1wzMtPl4E9fD5jH6ySr1+DQ38LMncGEV//Ptps9Aw
fFEuEgmlDTZtcM3AUg8Sxlg25VQAAKIIB7LZ/HaJSMH6CwnAJuSqezm70nSaO+D7
ch4dFhJg/TuixCYe0Sc23GWGx/VW9m6yIuQN5XH6FDTbmM+zVwT4P8DBFFLScb3o
6rg1+cduxAtbJpPVZ8VkT1aKiN6f2st4Q0ClhFh2/MS5hijxfFjjMOAdWngVWNb5
NqdnbZa9IGR9foa4tcEOot2R2nSEzzKeRH71JAQavdz7lv+iBZ5wLYAGTNHuLmcU
sU7Cyg7S9ukjKakfD8TfWTJfyezTfHwLUpgXlUUQc0P1EAb+OZdxhbYXLPBNRPmt
hDAg9HbtJq0Un+RsjgrfdP61XXraecdb7un040OjT12IXAktagvY7EE/k8g3+xPp
SPfkwQFBNMjJPfo7yPCA0+AaafaH3kaj8tKsp7PPkn++AlJeoKcWiEt8KH7e9IlT
OzC/UAoFgt/h7rvha436nwWfVKKmWPLKtYUMo1vM8RtvyRBHZZKTdlwVseyK0ANR
KikfNupYXkqVmJyeFV8UUeIvioPwZ9//Uoppl5biLFhqQqrGNRnytDR7ssEJpQJA
MUOfSzKkr1rKbeaoG1JZX3eSegdeXS3nxdAjKz8NBFH3NF5+Z/ZwIfB7V95a/cd/
OiIzKkX32avxW7wIwgr5qoqWmfRIjEG+oOn1TjkxRIR+PLVPBeLKov4PFubi/6FH
7AhwKna5rXWbQf1fwMda7/Zi9E0jBsfiwRaqywlMeHuyssb8Vv2s8b+uDWNtyxgz
0pIg56K1dRFllfg7skkmCQMmnuyEPXd2UEXaMFe7BsekIvBLOtu3UGAHgvgRq+9Q
rsJBouT8KhNJrF52C63Zy5AF6aH73YGz+wtZR1rOWmYtHqymI8Q4svcNQDhnNkQi
iiNkdbaO+0NupttXr4+3AsEqp5wiSplcKBJLRi+qXnNqmkbIiz0ipL56JctlCzcO
k9y6UZpfPDggYEgvErnlft3XWtXOwkJ40SvllWy34BYo8qgE6pWLN6R8KWUmr2as
W9Iurkj+gb6DO0+eVM3uBHLT8tBHipF0tHPhnvoCbrBkEqtIkTyoIABGhzcCKZyD
caohUZjJeSXCpDCiWKOQe39EMgJtWLjYyFjFaPF8nn3OCfpORCJIuFQVPZeh/Pv7
YAYeCPVqkK5OjrXggACw5aJV9fNhz42NlgxHbJIcDZFADnH873i4iercrwGgbmzB
omFZ+qh7iNqvMtPaZuGL2sTQRNVqPcRtT8aNZnm3MDgSOWgHVWS79lXIlIfjOqQi
ChxGNzJcZ7vHL5SbfeQ8HTfRd5qThGzszsyyNtUFcIke4FpWobSbloN0A/adn/lb
qQLgzbZkzwfmvRZCFQitCrk4TUsxvu3kBu1/Owgehvw+KU3J687ZUZdunIb+9/D0
bruqE8seD3NvuTtwjTrfLbGzQtvN62c0/qC4BG4tpr+4819SM2cTazyG6b9SqyIm
yXQt6B9psSdibmmc/zdIepnFMyJVzwhT+nS1av2lekFLsOSZwPwmKyWr5YXBGLbn
BfwI7DJSnvHBGbcgrvJmoWEjVgNbdIa8G3FleAqMv7YLE4WDAgMg79Leta/yVvcF
pz6a372cUAfbe90dxiS3fMzXiZTMO/h+K+40bmNHA2HGny7JPYu+grd+/azG5xW/
iPqN3DyN7mlFBzwVQZypt6HFfRyOLkMpUQFtsGKZL0N9C3O9NYZyKJiVBgdp3hOD
P3ey/53P+6LOP+h8f4DWp54mBb9UAaE8w18vKeCVIgDo9ykh79jJJMMamMoFckRw
dfQx8n5XZLmL77F/FtV7f8XtqjrBOtdDuYfGBlDXgMcvqy9RJEdpwY2QxptvRT1y
uScLz4iDYZ9HRrl1qp283sj0sa3T/cadmhqcTcpSPJ7h3+0figBWMoPrTlXeMDiO
WRQMqp2+UnGrFooTK/AxHCT97wcEs9obsjQ9dFEFlDKf2C6aW8hfSEPTW1ZFm0GY
7xXnMC2u1nfRxeBZlH+zuTkVhz4J+6l7H+j/gXr3A+8Lr0vJrhUXWAMSRGFvuoFy
MKWJx2KFy91p+y2msJKUckaomSU02r+OJXbQM+g2/2scGTN84g6ku204LS6rI4ry
vkYkzCZrJvpYzep8M6ItoQ==
`pragma protect end_protected
