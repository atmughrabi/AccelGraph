// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YAdwq2ebUa4ZvTqxUgYnuNt5qhQ2Y1fEQK4IYi/UBhzK6o8MN+GE0CF9IbxLQJzh
imUikdu8JruB4rCGGyrotSTmNV7jDJ4Q5fdqjZIj/UkR5hLQONQPRwiHYfbVEJy3
2CsYC0NJj6ZKUOQxGQjI++uLXVOGiKqE9joDCZNmn3M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30976)
lXdqjdSnPguSXQIW4qDVOH8/sy9dnsY/rSxF17K6oABHgesrosb7nqS9H82BjhDA
UqP1lxxfF3zlFFsSruwlmfZ+OWcKoe6AGP9aLq7JllpZ0haIg15bvlRKmovsz1k1
QmD4s++8UJ1ZzRMswQwtExkk5k4o2eeB8XnsalKEkcXBTvLHfcVzT9FwZ1OnZFzt
yLm2TXhx0VOt1RiGJW84ocVkTIEU/iD36p0gdpncnr+QlOyAnJ4KBvT8gXZJSs2E
IkCwiiGzZTMVS2ocuuCVCmkrPgAPY5iORSl463vwdzLAFshL4HRSDDfJ3gO96qpn
0ri1HQy39thTKpeEzdrD/+gfv6e7bW81jhQjlh1HlcL1jAiCWAvuCYHozx1K2zma
W2zWCE11utnSR48+n8KDVbSo5xroiKSUortTzAuv5hBCROpT5bssBbvGIpE51KwA
VbJozYwIgQ0zacNPss+CgiKlfxiA5o3qoLml4fw9qV00NvKWOSmdCjXhqjjLB83O
M+fmip2foUoCtKHLcJm5BOMkBiqYL89kv5vCYKnx42ikdkdsWS1StbPRkbqFDFom
P2XhCi1Q2dWp0B1EZ1tkmwK/XMV+PYVDMo0y4rdGdfV6pLPLfIDEI1REYnfM+kd9
Vcgr7JSp2dKQfgyr39pHL0HUissUAX4Vag6fpPzF/gwOk+0LKZll1xnzlA9TXAmI
nbeCSgKYmrC3ALKUPm6ytNRaaoOprcSKKxygbC55xe8KZ47QoKCG6ARj3C0MzK7L
r/4v6EWB2frS/uLS7VJuFgVKEObZioiw6utye5kB2OnFBjOEQFUN+W3suKhjUmWR
XamGS0hAUR0CHPdGzJxVG64XmeKPL9PU/vWCGodINCvkwGcmfqW2wncRJEXvvSKe
V19koYxoTM0wXxGp2fqGgWUuAqQPQXuEB2crxZSGxHPrUS4HJFPE1ApFujBMyNzi
187nibwTRsIyeO5Q0i2FsR21I0/M1dZZceygFdfwz8rgizQmxO9NQ9COxBKfJ8Ut
j+3ltKwUcq7WHZSjbSS/gRpzNdh8uRqbhpqyilN2l77FIp4sD/9vNJFH5FyeIFsL
kFT/peZ6s5IGYqaVoPZehvkHjy7I4Rejjr+XyLp2riVg71hwdWXf6yE7+D9glLbY
OP9OKJ1Z7cmjLFrgeTopYAv850jP3PCKO2uVfQA3UT8aT7Gj10LM7zLLY/YwEz/E
H5y1YeMaSpbgMzTl8lf++8Zr/1AIj5oKO8j04TTV2vLIc4bKSZl9cLBadjzlqJXQ
8lIXxBJounPh81LJEjF92KX+K0cqaqks95IGiQb7iyn0Z/Uty4V863yQi9bQGuNm
J5/hiKy5I8sCEdt+7QN/cg5EZgl0YO2wiJE3lKCjoTVorPOkztRTqUJiQgiSXcTa
sCWM67M9/MKaUKZxJpnzPnRMsGkDKZGLdacPSNHx6mds6XWat35BbcGRJlcPei6p
TkOMNehrO/xTd5ZV1yFE4+fJeLx7KD2gv4JxPazsbFExh506Pm2jZ8MWvGZRc1LP
HtW3KPUPQRGk2ghKXvE4nFwyCn2wTnHvfWsdtP0TdhTdoqEtqym2ySfb2rYWks9M
11aNGHdl4NaiD7nQZxsS8cfB2Zilp4CtkUWVltvAKYTV0afSf1fzVGYkHXQSuk4/
UWd9to1ryhM9O96vdhvhHvyClzBb5zywd2G5umF1ftjpRkSUygARW8hY+Et5BIFu
73hvZNhSRqw8fo5ZLGseeAbBN8cWAbQ3KU+2gQ6SsjTJ+pXpbSusII4tZ8zmgNZP
wbXia/a0Nszv/hkLqWit3FpBDU4iXi9+oFPrUFuBYeXwvqVsmzTU6kjeRV7XG4sb
NvOjUoE/590hu1J6KVmes13+leJEiOVowvLAqWskaKMMN+yuIA4MndKpFO6IC5NR
uKqKQ/xHVKePOli3qk4SurJrOFZFT/5o+uFtRFuwIQIv4L6AYyk1jiI2dLxp84cV
OYZBYDap4GRjdyNu8x7SHmkskio+Dh8sicTy9SCJXeIud8ltCz2jT1XxTX2RDPCt
vTnPiFc5hHDpyGxzskceJrpqnVbEfz5liiOKT2e/0aJBc0Xt3qtMtpnBC/TvH4LB
vMjk95VN890Vg02hmK+tRYb/iAnOU5zojFVgnoSno3XaMUMLuUXj+fuCsnX99VoA
9heUVuM5QLeZ2G0vlb6g4xHWJ3kvjWtMw6Y1PFIXWHKioRu+ZEMMsfLtTzWmlsVc
+yi/dJ4x2OTADu14Wm2sAFt51JFQqgiqbrrPeLznrUm37P55WFGR1u0mq2AWNl1V
ILCv5NfHXbfSSkIMUrdBLln1CLNuGomJQKbdd2kH7Y4VP5/VooxygD3tqebtiwUs
pU5T15AMKxN0DBCE5q6Tk7hkIKi4nhMfZCt3D+EjrWxU/Jm1krMyPMyeCRdOAHiK
KdMdZ1qfhZpss+TsGRbua2IX7qRwgVqcVvlxA7StC07gvgG/4GEJcIDeOymp90tD
XnPUosDsX2HWHb6nKLcKMqo5ni/TnBVddo9t1SiLH/TWdcTzJ/S+e1iF/yltLZIb
PIZqfsicD7+QFCm2uJOVEuGFlVRN5uoVTK1lDRgit6OYV2xur5X3wpUgkt2xXvoF
V6qC1gwjO4/rie+JvcrTI+fjMj9muB7C+AnO2bY3FoyJH7Y1A8WeM+wRWWaA/JOp
aqm1LR2H59bTiCrfpFnzwr+Zp6+ceqemcqTXrjjYIPmfZiH82lP2fg31JtxsfdVi
G0PuUAlMKVCELibxE3QR5qi0/ZBsLtplhwq0NQ3NkfdJVJBa3CAK0MPR0L/iiKHH
RngVxLJF1bUkq1mpjiPoqAtuLWfKdeXs35XR08wQ8odkqNlzJWoF32AXlhomg/OM
0bY5/TKGyAq8fLa/tUod7RbF5f0tA7Jj3Y7Jxq56b4Q0QOPzuA87MhyCcipVLgEP
NugMKPC048dp+1apwKGN4vEKUcF89c36qtEPtDu/alBal6PprRXP7D+kmjhAlw8Z
jlK9/vGRHPoFwLLsMe5+MQKYhUur6aIzE/H/DT3sPfZsDGGH3eeWOTSboEAHFH5A
6mSr5w91lrVvrY48rtNq7PgrmhwiugItK3ThzPDU4S1KrKUrbAUacCA3xGgZxkpr
q0hj5DOeSLK3jml83ivTznXix5saB80zVeCf344PCRoMfroITkAHiVie/+xY6f5c
/9iMhRrBckSNnQRdqlvBm456Km2dV3NU6AwPD3z4uC/BnWH4+Xq8uYGDjERiWdvc
tKt7MHHYIr0yS//HkBz/N3afmZEvKQRfVHYM+BUos5MYJUjMiGuIYP8GLGSMIKqu
UZR1QCYwIhwXOpcnGvxIcsdWUvO9q5ONJdPtZ0ziIceKuMvefSqHcL+oGnbIkU+m
o6dmcse79YjC3N6TflwmL2TzIichBapFD0e68JbDhjBG4tWbTLrqZ1JnxMe1WpCH
m+enmAmJ0DeIM6lc5etwz4a6k8aN15RXLcR+uahiHHmSFWpNdQqXyLU86o6Wu46U
axNQRTE0W6aB95fgqW04Uuc0lD68jG5HDlJEd9ui1VvIqUXNBp3ZvqZWyFiZsUXF
gPL0qR0WFjKcyHLgkdx33XQKayq+CrbQpwRBm5aQB+QMQD7shyHCOPTpUQdp/TSP
LbSQn0FZ3gvKc3Jp/9RlK9Ps32tUBAv9t7K35u/Iqi6hNtiG2Wnr24KFdmc+IwHt
BJ7ugjco8vypSTfqk3OUU4X5KggF3mtDGAskuyAApEyYcCbOewYDTaBjHOQdx2RA
gM7KfL136KqHSlP6qYPK2Z+T9ZnYEGDXucZ/7YCganF+zGk1VV3h4lhTSBOSDknj
loBsdXl+D4aOZilJh3YtXH4fGoE4Ici6VByGkWRGVlBwqeuR0bP6FGFePgjn8THj
hmcqQec5wJgo+xdLqBjEiHm0vDD2hIDUEuCzvRgACe0JbSH2KxXjMQRTQiJjp16x
1uMcPx/JT9wGKOKXu3dWB8shgbP9UDaA7C/HthwjDgqIQmvo11ZDlT7uVXcHVyll
ospK0rdScwY5EHQBP1AbhlViIal49+qY2fpmSy07Qj9efvBfA4AjNAGop0aLRqVf
Ke0fnexACYQ/VzxqRcSzLMuBRXajHQFovqARf3sBZr0Ei/IRmJcXBh4mN4EO/ZLP
rgpFnvJXF0Nk3B9+uS9/DGxzd+A2ePFU/t6JAZ9Zf3TMxKCKhNODnx0cibQIr3vd
i1aW03k/3aaOriU9m79hKTcl2qGtaJ3MmrcJTRfhUdY6PAGJ0JB6oyXM4POoD0qF
ZBiaYVnxd0GtWtybyK1P0bu1axT1wN/8zQRpd8fPH6HSEcx2apM83JdVUoqCcRJh
jZn69hPdb+NrVvRSmNeuODYR2graRljDjwRzp9zA4FIu/SyFc7Eon5thvDWW8uwG
kVwmex1C6CZVOqcwEBTJUr4z9Jg0gYNaMMiP4qUzwlkia0mRhGfXSkoGc9DTV/QZ
y03aPG6+G2hLsoe5ycbQqPaIhTmRd5xh38NKyybTUg6GlkNOXH86TOSI1axONvGD
Erv1CRecwl+2ILfztPUDtG4wgCMSIfZNJ60LYjGrVw9fLDAiOtOgstcM8nChj/w2
HY6d8n59g43bTiuK5D3e+lILwMgsSR38KI6F3jYbFzB4RvRTTAl9QfPzO17UQMGX
qIkfCkkjGl8G6WVueS6Ik7Uo+S9M3RnNuPAo3kpZjxwpZF0L/0rQWVY4FK2s4MCY
XC5QO/zD8/VwzjcGtLyT/YXk87SzOufo5ApKNAXbk3w9GfUdbhnUjmELQT1NRaHQ
jAcQwg3oOlA5QbHe95H5Y8GA97onbc/B9cGRiN2l+qr9x1g517mkxc0nQG2mRhev
e0JnpBzDISRJQYZQ6nQ5/FtE37RpxRtP36sz1/vLDg2M8LtJTVpXNbSzGJ8asOUT
vR99sMvSCDL5MSCUftP/q5uImioYTFpdYSU9QnqAc3YsVY8LVHu7MHXAxSyZpNoH
575FOZHMXNktoRwDUlmotEwTPLHsp1rY5mTbyPs48wW7QGFvruo9SQenHSj2HrTq
0Ft5Zke693fKt7JQj2O/a6JCq3VOhdDcdsM05Hfm55JHwdJyKu/BKjEszEO2I+0m
ispoplULJdWMt4vc2WoBhNRVmciaRH4H74VNcgcPCOqHOyVmtKTm72UDrrDV1IvR
g2sVL7opYusdFQyI94xs6+h9p7pSJRgin76sM+v/RRhQdLOjd5XxOEqHPq5qvI+J
ohIxt8iBKblyJvv+Y0C5WQMszXb+e73Y5hBBftcPgg5C9YI9b6MQuLIQseQMyd+v
YADAOLN8gSi4oj0SPWLtYiY4T0BmO6TL+5A3RONDPFb0XiMlC+jIch/Kb7Fkn8y6
tymeOKPM8iz4TvBw80Or3n+vH9/qAiOSojnbx+pj0Rsit+h9f5D37K7DwIzwBU6M
b9rX+XPbReoynvdv/grLwf1cXULp1UhfgvZjkX/12Inx5KJNrKPReZulf1bZrHvQ
mLBvGUpWwEmrHpHyeBEtDdSSmLaN4cefGNRxCpf2XC7KpHnlSemnyKlIHCs1LbUN
9r218l0dGREs6OPNbVzrgzbN9PXyDu3ak7p9ApEiV4jpWWKb8cQJ8aMuGKccDGxB
h+bycDgnEUVQMOSPY5AvtagvkSOHRh8ejINwGPlIZFrdErmuYmjhTdoacjlTQNQJ
d65llnlE4iX3C8seTOaubWaMJtDN5txo2upi2srGcL8jdIrs3Ya3kFkocQvhRvEm
t93naPGCyi0NhzJa9+EypTgPF0EuOkVufgeEBGeznDXq9BXUeXDCO2o1jMKBegD8
Vq19jdJj5/UXPxfkEtdpZvaLhABog2xMuP9Wf0uf8lQfDoiIA3yPLkJsE7ndQLwF
kZjR8hsltWiWGQFCthaeOXk3FN3UhKAJvhhDYaKN96MrOjUzTDCFXy+FXHwQ9Zuk
j/RUloUGqnFRVZ/Cvbuyvvic5j/neHKNKUvV1lSjLlAcjjqTb5DJtHnliDdJwkFx
v2on0T3ktFgFuRn0kh79UV4P8bTEi5S5Vs4J+F5YgtW0DU4gQcBKrsbBgjBD3sv/
CUfKokFkiQjqml3I96TSsKIgQIOid1fdDRkKlbX4/PEZlMOSQtYPpVzL1HGlb/te
IaVZtlGBPEiU5Bvenddpjv7IuQPLd3oTGz5PUJfYMuD4eytSCtE8LmnSn11PR+1F
0JyohYm8Q4CoeYux1V3AbeVffSFOrIZsOCZZGGNsa4GqYFOC50Imp+UG+u1Yk8XX
rs0Bg/qhJ9gJQjWrBALJsLcP98kvKzDbOxy3PjClaZraoKlcuCAJiPVgqhqdRGWA
t9B1pdhcFDPlOC4wTyk5ms8kQbEeeWOSuv13P+3CdrWSHK/e+6tY6YeMZhy8wPvZ
1cMScUhbmJIbbDyescK/rYDtDPva/ph2o/DPHTR2BZC2YgKF5exXX17dQWcEjVfg
Xq3a6t9RDDvOUJrjqQMUUSVPpjxhANrJRlcUpOHzHgbyHYOaJ4pep75AxOga0JZb
10sdm8SSLlCuAeBUe/65QFuxUBg0eT8ZMiqflL67avZPRnm94Z5fkawG7tdMG7yK
iERW2/QmhB9dQdinbRmWB/ufXebA7XMTNA6ULTYLhXT6Qt+ySHJ55KtrZLJcUzz7
fvJ3IXqgT6J6vIufSzMP13QhqgMgVLYCQHZkcPDQhu+TLnwE2baKzWNzvYh8/ZVs
tcmNZIquinXQtdThoYFvFvhI4mAWen5weUvJRXj4pokxBRgMzTiTeLJZZ9iSPyED
HVH/y/uJtrUBGvOHKzU83el7ueqwU8rJSz9mYGTJbpDmhvYZPEcv5dYyoNMOn7El
NpFv7x+H8XObBfsg6tMflzMoVjkfYoUKZUX7YHxIxzhM8W72mQTzYCCJyoTfFU3h
OzJArVFHCKPQ6cFpwHYRxCYJSEAe+PUMktX6dUqo8X1Vp6A0KSAgcDlWZYoW0JK7
b/uAgLueYE3faTXUiroERI8qjfs2Y71mAII3gNN0jRFkC7bRgeZz/a1W6cEQXoxi
BtaslkmknYw9AHZXwJfAOsAYEa0WdNXcWARmAoGD77+z78bhRK4ou35Skcz0kTOq
uG1HlzmuCNIP5YBndPDXkerXhbmNNZ6XataUjhDWcFLlkRqTwr8TbT7x9wyZZvV9
8COBvJMi4lXGSs2/Os0uAmPTccgz/O+BYsCciazO77r66lgBE21V5NK/QpH4urRE
iuGpDT3WT3h/jU5pKJ5ozTX+PT2KrNHAKRtd1eVLyy3Oqy01bVs6NyOTJZksv12H
L37tH34SCQWfyR4uwKA21DVF3XY6Dqok0XNruv2Fgf4MQccboUabpJyb1dsHEsh0
gfgmcTsgGwsM9ra2oRPxxAbI+SLRkg5RTvwYfCPr4KG5+pJaxkVe3FyfrDwqmsKW
ntGbJ8JFFFZc//cdMw+wWCizf1okGOuKFVwHC7DHxAfxvqdh/ptCqfDgXi8vLz0p
d/JkxGtWelOBSh9o7PZOp6ePN6hX2YJ2fxzJCCLg9u20CP4evOP+r7CbchVXa8JN
PtaJjlwbry3wzq15Hhwb5b87gWPDs+v7J2uR4wcO4O2ngNvbmN4TEJcS3cWgV/n0
CzBX21khRb8BPv92Z8YCdatCnQA3AT14tkpwLJJ12cthndbStNtUJq77UcCwEtGu
5PVXqAJXVT3mzJBV17zQcA/tCh+NeS7NEGjgnDVk36lpxRk548Cw8X7Fww64nIQM
L/Qmfq11LkmmxIF82PpLA8h7uVhht4X4oePOG6SIDniEDIAYypfmUr2P74TA+fPx
zzvHzL5G71NLw675xmJtRCq0MQTXh4YxispLXonEFpJg1kxZ1u9g2KEIWVxcTZ3C
0DjFfExVUKWWw0YVemwE+WCsMJ/P3wicuJokKqNky8HgMH5VFpSC6DWqd7++MyP8
zygEFvVLU1xhSQ3ZXbiuFmGgiC3MjOZQaEUa7ad+fKSYkDmu4udenvvc5hd52TeN
Atd8OdV/1Cbg+TY/paXmvaWQofwkNfL6f/6v6odJGmdb4Jh0v9h4K9T5jiIWMPwB
VYWIRtdt6zmr32oT7ipotawjFcRDnjizj6YdofreYJTXU1L0HC7U9WDt+C1szwrc
UGivquPe/BsPX7D0kzKo6Lt3cN3M4v4UJLAlygOdb6NdDh0ijugcEC92pWmU5dN2
00BnSNWzNeQVW3y2QenLnTg0IGQfUoW37+L3rOZTVWQZJ2h8EDPplJPNLz/4rxuk
UnNbtWNYQOZPbYwi6133T/v2Gcd6lK5GiYo49OzaY7FkPugczpvu3Hpx/e7DD4uL
0kJsp0hQmYSb6R/JuXCV4r/QGR8gu453B6lG4IclVRZrgHT5OWFBZGYlIwCbQCNj
0BJtDCJsOhsepKl/RnuAZ8txPbLd/n3nXZ+s0wIf/OVWY4ue9Y7fJZeK4uXcIBjn
U/CLEA6sl2hnPuEuy7hesCACzGoGMzB9k7/vBMwHrJzNeZGbe0IP9+IeY8/JWzsd
vriovesmBCsJJw3to0mf2Glqe7GX+70Eas+rPlK8Cqd1hIwACUaWnyFndPY/tuzV
xxS07F88vEFr7OU/j8NooAsVayrCAmMF2KKxOU1nmLTBkGM/3fBR6rhwWDCyHO/y
qax3XtLdqyFNA3jeYcR/A+g9enremft8gYOF/eaUNs0kyLh7g2aeFO952COLouKM
azhkUibiPW5gwr6Jqfeq0NKN/ayGtVpyOU06eDtEA9QjFYuqHx38zZmzLGH90IZO
7dycCoMoJm1tBGtnI1/Z44P/XBsYt2gFXxaEhhNMNi8uvOTHrptlagvEaGTTj5gL
kTbwYIdVSrCd6r3/1MAHURj/9irMN4LliC6VwCPCvOF2MFa8Gym65SGy/2UxTcLK
qBhZnk9tRPo6Q5ZJX22a3OofXJcl9gMJhW1jUR0oXUavYebMEesgrYjjTnO76hCF
9/J/qBKcVnhuYckpWyG69f69TljoHryCX3jSNvGiFFPpUfmeGf0HDAStpGu799BB
iQGEx6i6K0ltb+K2FnFspMUUcQ1d80Lvp9/bUjYPzGx5dBlDejXVYA7zjoYtV+9j
ElVbBR9uGRPmXYlVrCU+FzfjJp7HGIlo67rZr5MHgb+CKh0gGRACRQlqYy//3KE8
dmSY97NFfCM0OieewIQ9IuPJGXhFB7dg2fK1Cd/nrixdtMw2XEdsqlON0DgfVOyF
kM1J8CLfMI2ze98BLTCYsVYo+WT6uC6L6Mi085bXwmnpDwK5vaZCsHnBoN2NGNgl
pJyIrPcv/qBZrkw+tf7DQciI3geiIk/leT+L6Jaa8N7kukIHXb7XVSKRoVzsMWmE
iR9YEdXwjZtcaxaS3Bsqa0ywOjOgBfNddcUpr6h2PYhOtXxMDkNYiNU7fwm2Rvob
stkwAEtBV/z5LtLUdUvfZBRp0qsc5F6232z/dk5cmf0dY1uZrPzLA2i7yfzTb9+j
S0U2M7IG/AZaW54IMagiCP2fECfFS66gMYtDN2BMLB9aPqx3xfG4vvr6KWtGcU8l
fa8DiLeyQ9ZwHZO/gid9TqJ/+yjoUI3bNafY8GPdIDarHHlxrjVF8Tbk+Rwb6Xlb
E6JZzQYF8uuAhi4WqlX/WJPg5ZPXLXDnMTXf64U53MM7yiD2F7g7vLmACVv+ZF4S
6jE+KcgcqhxIoc4WMkvq0kcfYWNGWo0rJ8t5MLLbd+ZvMBg0hjH+VmNwrIeuvaUX
RjxNk9O0eivmrtbVZtyTwwMuluD1QsDPJxXq6ZZcv6ErrZckI/CXsi1fWeB2qFZI
KGkWRYFXwlvZvsAZXCt1ff+mpIzI6k/k4OwGh/4MIhnZhVChs45gNBKwGOjkICxc
gpOgvMuqXiiZOlGEixhcP8AkbXY20zj00SZrMDJQDC8lqDrqEJ4UCAnSS2Puw6tN
jAe8mMKh/XvhdwusjoSLob3WYozMVDt+2Eo/e/t9fPiXn8iu3Be6POScOqiYcsfZ
Csj2LXGB1tULe/IcPrFDiSmYV71vMxMAS4yw1v0YWuUH5uitrVElkTT6EBtKbzPi
UIygNiMklhGvLtXbb10h4dpgb9a3/HBkTp09JXRuHAuBv+Vl0AQc0FJizIoK9vNW
NLhZhEbTikhW6aMljT5HFBkS6tx9IkQ4tEz1dVrt41LFQJz1WQ8URV1Fi9tPx5aU
zHQac37S3VuVLIh3dr1T/qPaomCUYjQZ+G0kLzEK2JMR/OFJcm+ExUzq4oiMx1dt
BDcKdGQY7CuYJ22ZP1n3zoe5DoqEhzAzpj8YQqPkzqN1xWuIC54DizA9wdyPrAj7
YZaMSa+4AicUDPJUW8NspdnfhmqWTSIVHB5jMpcp+6mhVF/2lC3werK5X9R+uruR
z//bEMoLRjvZjWqA2zBRu6C7v8UeiqblO712XXNFUCOwUOtmltT6n5FZCpd74zzl
fZgukCVb6rAru7LHuaeKZUioptoOXbz4rWUMJqLCgrtirB0tf44mGyOO5d1tdKSB
wbMWfhYgyejfZhyAnpQFbegr5cNzr2+DaDa+nkU61two/lQnKw0sThSbx+Kr4YHq
WTPqZ9VVaJecbod3ZCaia3mQcdgq5FJN9STZ8Z8503W6jsGVAxZdwcR3xo0powjC
cYWKFDNWhXuqi+SJQ1zEn/MJhmRWNHE4iVqxe4Tv2HG8dWleXNGHU+8h7oC1CBxw
jvN1Z577d48KXnBQtkoyW+AbQrdhnYXWFCA0omChHqPdpOEB1uqBuAvXd0nGmjw6
fLRfSCk3YT/e8E+I3DDJ9lNPnzi7pstqrkH6o/ciTyoJSR4escMGJNXA6VC8jUNs
2md8SVFkhyaQ6TytUovFR7jldPmb9Gy40LBmTq7vcqESWbmxExZEW50oaw7MUKPu
kRdT2h0bWJ99kHbXMn6UHW0mMlMNK8e9KUcmZnmqRM/omJ/cmTEj/wWYae/YLZa2
EUqK7n5GBl2DuS5cYj4m6TszB7zFcijA5sazAiZdsnR984RGxm1x/lhWLKrgS2Tl
AeZx4hKwQLi4yL+cC+Q27Xd2ZlrI9cwOgiYjYEdwfy155bVYg999HnbaS3u0756b
sCnZDQA03iwSZCTrCeBrm3yFGOlOPiO0MikMtIq6Stw+yjuz0SZj/XU/ZvLSWoPc
fGtsslDoXIb1e/dYhNT/oumSelDLI8mVInNl8w7irfCN9u+EZhTnRALlty7T7XpE
yyXTzINl3ncUj0yWykAzOE9dIowbpH4tvAXy2+smXYL1GCOhGf8HDSg+VsWfsoXL
Np7umHeNtJ3UvYcLfxBBloRnppDfK9k1DIoWESAmFCBIOgVLLM5p2IQG3wGptOth
t5YaAP527NLSFpP78vyA4CWW3ctHs7qit3uh69KVmBhzwc2t2G4c7aDNmY8yMQ5c
+OyVjvpdoU0azPctpCoNVaK8GMFOdX/1mw/WJiVKbFqET1e8L5ZFdNtQg/Ujo6VO
cBX0oLtWeZvvlTRKlXObJe4xIDg4jsGDxtgEeuL8lp9hXzqDVR1rmRghIHKqA/Uu
Ymr9/vJyAjmAs/47BQMR7RSDQs3pCsqXesC9IaUx2kZDI2JfQGwQkvokg6MzE5CN
PCfWNcULwYY4iRXfSmRI/LCDXwq17qYELb2CMg78jVSwpXzRMNnAInZHtGZyVRhj
/AiScPbOY2loegICTJrw33ro+e2XUQyMOAsN5zCzlwOpDbiAP4V4d5Wnu4kq2l6f
SiRN3rWfUosVirJ4WND/bGa0RADDm+93NwJWTF5Q2H8YLs7b68Sejmu+fOLYRT2G
Dm4CdnjCjBOwCu9ajX5g0lwx8hpE95ttVLQokk//aRZRMQpulEzRMglDcpcDXI/E
flf1I7kYfuMf28GVKsMaJal0Eljk/Ja8oXutdI1bRjiS4JZAYT20NSRKhbnQSh6F
rO/02e1SfVWiiGl6lEHI88criE13HBFH7igWXvOFNogMm5SVbxKYpqVSJwAw+b3j
RC88yKMuVrMiu3Hn/mfXnKD9LjAO/OTDknvJsLItkaZYdMQaSYyqC5mvRFoHgRR4
5mxZSBDD8U7vSLjWaQ8Upmhhz2sE3pWGS0QL4u+M//f3h7DWpmHIxemXY/isQ3pc
aoaCyWa9h5xd+oQ8hI0JzquILn7Upa/hNpeYQg66tTBye9FU/PNu7/yrN1a3eTEA
ofQvXJrz0158cnqJOyVAn4giUjxP/tYxvZXtb2ouWdYMvFmI6MRyaHVvPdXDWH1U
nVmwDqXpQ9Cp9Qmu3F6T5+ZzDsoGW3LPfGUfnbxYjfweZl1OtHyGLpePxFg0qsoz
TEuhYitQfZ1eUETdcMW05Pi2o9LRh/EkNIV+Hzh9KhgXWmJnwuvO6VMMKleFeM+1
kImPgO8QALDOOkis+eFI1Hk2Rdm7NJChZCZmZrK0m8540e9ctqZHd436fUUsYtC9
n/o+y7jibPv1eKhFF0+aHz41MuqBvfSPrIgUlpm2CibVyLACkHOboZBNqlOpHPDX
MmdOfOXHd16nMH+Yr8Q1TiGlM0v3Tkc3E+iWRWzTl5B4uoXSNRQbeCoI9wdlOdLh
gErXQXq0s4KZIkae8V6o8YmI5PU1ShIuYdtAYLyMO3edpuKrAvrwQuJ/Gkvnjt/t
VXbgZHwsmZ6dVxkpU1XZSOfKqOnE4UgJFPAwpwfp3ACugUaEspvaHxYKOlNyq1Xm
fcPst0ZtLx0es6zrSB2TxOY9Th/a2FYmQ9F967pfhQJQhKXzgQx7f12e9NAiXGS7
mOwI3A24nSFEt2B+OmG/adROZVszUmJGxruvwe8uobfwshS3PAhme1slwllCb52/
+pHusXAkL3PqlvqPgQOcWazajFP4rzdqaQrbP+8vh43hjAOK1sW81KISEZr+hegC
BZgO1tKqVff+RXYXYbkRIsprlHrT5pu1XnvTVdWfCLVli5wy+m6m2QEKAw5LPvEb
YMPSytC7djaZWGW/F8IzDEqvH6+5TuXoDnzcT9XRhWCrTUk+uILCMwDeXGL5vP84
EZ9wRnN2NmU8KOTcGV6NaIkvzVOR8O7qPC1DM8NOvb9fkaYSr1Zujbb+NaHK8HfR
LmxE/ETDRZNbhOyEksCt+dDaFAvbnhziFVVjixLOTM2vdg60Zgc8AV/Yu1Whckkf
x8K6p+UcZcHKBys/5AUOZ/j0vlTSOlAw5LOtiWntsU6hCPms8SEFitVQbWPLNZG/
7GAMExZGNainN8e3HAI6jHdAtX6jvquE1QUZk/o1YKa6/g7qHqNai5Cb9Q876HJv
CE7qasUaxLgUZ3IPmKutwoJAwyA1+s+ZjWKRhWzkklRgK0Jd+YH38jkvA5HVXTp5
dlq7f7URMRO1ZFsFW17+vQYczcxZqn8WOeIu5B9njG7cofmXYz6Z4hwwg90+/4f1
jLeD++d/zhvPjjq7lkVUfzTncjQgVfikL/Wp9qvYWug6bdNGEHafOoS6ILNiQ0i5
isNjWWPh1mgAj1ux8LEPWmc6I/5kDiu9eX2MDygBKPkY805L35GR828upJqDeCqn
k84KaOlD5/avOizYvL9qws4S0rsX5nVcWunELNdzwLIgGE8Sg5mrzeQIeZfwkDdS
TAzfr/2IJ22rj6Z84n1fRWpFSCdp4SBwqTZQVreNuHEbq1Jmri9WNjDfq+LVrLyN
JKFW8CMdp2VZYnuAm3ut+oX4d2sgnfuErUefZr+b6dIrU1YBqRMy4krHt+38ftw+
Zlrp0gNhd7MWJF5HVhISTomndr8cme91VT7dHHLylAjSvSM6ZSPgEy30AFjPYZ/L
kJsRFTnTOP6SJ6ZO4boIen5ediI0Rftfhkr8ApHvrIZBvBZx49iqjvgmsBheLgdK
XNIYpBR8i9dTtNdf9K0jstx1B9R5toLE1oqLFWSgj23WB4nLfppJWFmR+Dl+qrVq
YdzJtHH5qrnLFCGI15PKWalpFpB4I3rZDs1yba3ujlYgRNtsY8rTmenz6myilDWS
jfyslKnXZV+lg+XNlAFHp+Ybc6avqMRe/FB8gEG1hqtdtghtoaoaomvWMXj3+tk9
bumLAWIp0HX9rPBySsO2g5dZanIRtx6aYlXXv2GJYXUhgdBjaHaJju80i78EHEiS
GvAoIAqAfTPqCYhBqzGEIdL38XNokLUauwhNZURp/5Cu2VUfguR71O3VOp4dIK3L
UxXwvGpoDc/L+JIrcePItSVsFChTBzHTUuDIx9Nr5ut2znSiZvhJjajunedaZmH8
LSnf2uaFoQuLHld90hYKqNGv0mv5LmS4oowpzjFxZiCcK1N0endEW8sik+esBJwf
EO/xWBU19hHKLgkRsLeiKD8antykG2KUDpNVtxeL6I6gFKMERjH/5QsZQa44LKin
UedFnnHBJN25HdN/pxQCLOhKUvUScgeU8tV2pZqRXiCw0SMUA+mtEYXHh+dstmY1
FNjq7zbxu2mMRK+FWkc4cirN32CgmtRFjKRzxq/LlRRvr2mxEMKEINoiVbkrdf4z
e2DZlNKkymmNmGb8R5xP56VQ2hGzpj/gyrnKz6JYOCxgFURjtTmB+S27n/Tr/h3o
yEhG3fgSFllODXtySRZKpxUQFet4ZlVHlCgjRGKNPNlTW02+ebXe3GmMBtXq0k5d
jRKCzAxrWT9hGWeshIWTEkZ7o4YYuhwaTRr9WsYuvzIcO7BN6q97jdwsePJYdr+K
TJk6acN2tWPlhOzPzqRYIOwnuhh3V+CjlzPNR+UBqQinUvdx6wGFDz/3Z/eTtxe5
Nplg0Q3xvTAlCKaM6umZmTm3lrXixpK5yWOeNuGbQeVHjc6yWzn1jbE3eJuStlWR
Jxm42K4Xy/fhbtu2rHjvG8xsn0A3WJCCJtGxzgq/XUngEKqTeMw9oD3WbesJVdht
WupC5cGnOBpr5UpXzkyDJ2xKHGzz2vzlpptnzRgsFRB5Us9ftEIJx8HViBPoh1gp
DKbyq+ha5/u8h3UnvnMVDYE7yEP0iiecWe1DuN2sxqL40ZlGQCWjDwgmTX+tD6j4
3/vXPu/jDEdBrPQgBKcT/Ih0omUb/FvzXfgSKAPEVUnxbsdKQAJrsEmwwPyvvI5B
V0wkxPFWxeSw3bnlE2V3Bp44A9dhd3XvIh+4hUb5olsfy3IM+w65194zAL3fepYv
fNPbyBWC4Fqk5Fvi8FvWZezJvomwMb4zekomzcxoKyFyYiBbBRRVLmXBQ8yxvWk3
Wx7rBNu8Ec/MjHOlUkmY0dXGJtaJZf1XHmlaPlGv9b7hZbdrTD6zlewIGSyahPhA
W7Gf5KNkvPLntGkocqr0opdvLJNKVFsQWIbyDGxrcITd+ChpNCYCK6+zAaKpd/YW
Uz7nR3PaylGhizEeyf/qPXaeSdt4/A3o+nu4u4KcR1wcP1+NEbwo9bKryhrdVySm
aOTuzvMaJwArO6dUWh2D6JdOY9ljO/KlpOzPs2dako2NczGHOzJCABeBvGIGBuDI
LnA2P9xoiKqkebXMw6opWZwrMIqrgilhWAnGG+gVPRx3WkwWoVVzxelylfKOIhQA
tkWhqMutkr8J53QvlQTzQLu7CTqYH1A/4VJT8wAOFfqAtkOWv80pU56K5oB3n7RW
E8FtgXnu7yQNmqJrHxYeCQgEFkdASCDWjIqiYJEfbYvT1Mf4We7vv0M0TKSxyS27
DujCaUZVA1s4wItrZDes2+dNbJe0Xf+n3wSks2W+xY/SWW9qcoijyfO2AD9aKDUD
0j4eF9iToNVwSOARx52ztw9Q+7xo8q4gHxqypqXVVs4JOuHXMyX1HbVI//UBNbMh
cpqUPmNSIIW9ggJ9BPBlufcc3Ekv46oJ3+LdookWutMKKN/A6NFQRyiVZSsYsWxk
7W9kCt5s8xjPB+OssRANMhuTXmWjg7xdrVYpt+62UXAeG7pIM70XMfP7R9rYkWjv
NLQ+7fZNbpYuFLvAEjdnpKYc0sJvcflOa52FOd2jibMjArctJrwvm2fVVOQza2uS
SpEGZzwj8IqwqtbQazEuyHtD0t6kNbHSeapH4ieDcNp/koYWjMs2J7VMuSxgzqbA
hlERrTlnwW9zN89HMT0AoPnCQGIl/41QqnSf9x+s169SXyB6rSGvhP6rvgLkzN3t
PtqYzawq8qPe8GO0Re9+v0rfSBCRPW1HS/eSUxK2l5X4uDfTx0PA6yQF+j+t30ry
x3qA9jTThdPWzv1LHYqQnaLwUgxOy76FJuqGNZqcHEGtTmaFEZKM0rFmsdLqiTZ4
PdCDx7KhDfITR5wnPM87M2EE5WxikyqvANx7yj0lUwZzZYACEnfSjlfCbZAM6KxU
g1gHhVeagSmCYdWdLwF+8Ek/JzBS8RLZtcuL3sWd5+KovTZUngLG6Eigp8wHzxfx
MPz3xERWRXRjbjBPCuqmW6NNYPuogHFHmIU2qyRYJFkTyAjbC8HynPQPnYKIep0O
Q8/d/cFrhgsbWi1MxsQnhbO7optqB93mYOhMyvHFdlOPbmYtJZu+hynuL3ohBRFt
d1qfM2l4hQygEucDc+GsamQFPpvMKEFlYjuRZ/HTnLO593wGdB5X3U+cax/WVcnW
Nao5NOihxU0hiIenLKQFWJDBudypfYZbWTtBOOl98t4AxJJ0LxM1bNZoPBbRV/Aa
y6UQMsz0ydHGa6QO7klfKQ46qfh62O9eztHjocc0UdLLsegeJPxW35MiwXHoDkqA
j9imxJyN4uJXyleyFfA5FpYHNMYQqsJ0vYXZrAter+qw0PaCI8gglsvG3P8z28db
MrPTCBFyu1u7qSg/El5l5GTVIl6U1iqFhzeMaqVXqYs/j2kiQAG8H9DXOTMZE31k
pTHtXPYzfEdXeo504S+wGqS90F7AFyA4GbJB2E0BzWxmfoo7bCpCWypKpNEdHlK2
qyOPJzujTaI95lMFBhVy6kl8OtqZ4KWrx3YcLwKZuLeabKoS9gb8eHdJMhwxLcdn
I0aZkbDPMJaZFPIQIDKJxo4b3o6xPS4u402YoGc0aWflnFbDZQa5nXU/ngKaL5Nx
hLuFoJxIcRuMQmsIaiPA+oQLecikNWqY5zzRDZ8R0G+gug1U1JPE79J4GAvEL44M
CGQk4B7gB5oNkVXhBbh9fi8f+8c2YnDLbiQIQl2N2mW6jMRrTutaABkaD7kIwgSK
XHVZpDOyWZAfaaH7kMIjlIFDeujN7i02npDUeRs3W3Z8TEkW0yn2QVDqi9eLYv7W
hI9hAttuGUVf+nTI67ZTMkrXGPnARsNG+JFqu9y1EI03bf/ylTpwk2CWLozBeSm7
P7euN5Qml2NbQ6pErsF5L30nNB4nhaGKL/whZ12UaSlvcTJLE6sZOUgqecrz3/eL
GfZe5KjhZH4dGOmjfvdxdLqrnifQzkFONl1tQSoj8fzSA5nQtg79DmINal0c27E8
nnZpFmrMe45RprOh5tDHehP4779dNqmuBCKFMYtj5Gj2I+WVQRXUhXiUgSnCM9Zj
Z/nqVUeMZBYhkA3K3KAx92MY3PbdnA2e+iDJRywMWmRNxUhOxyMFtogl0Dfn9EGf
VOfDq3glmGWY/M8/Be0/astZ5uMpwjdpU4VkjnN9uIUD8Osf29GsmN31zNU7bo30
bjaKm8pwwY9orH1WPODMYH825ZZSAU+oZwrsm8cRRJUROQDf68jk7nwuOBYq8JFe
5ks/uH5DQYn/UnLYDz5hKvGJ6GH7naj+3eEFJofXCAWMJypZP0iTrDyLXBwuWEUj
WAjqIQvDelz0MCPBBOlZ3X8MChGG4pCP2EXVy1x8FcooKUfPJ4a3A9zxLDduN7jQ
/YSeBsKjMeWQcJtXoeQsYO73k8WTB94A/JD0SGKB+1AMkXV43vRf59AocpREvL1J
CMuaakaHiDWdmrtNbkl7yHdGmmhSuXxBKaf6ABQ05cP3i+I3AV8esD9T7/TlIt+T
iMy2wAWx06JEm3LBDwc2KEQ3b/CPumGRg+Klay4Wpr9+HIxTLnB6+yEhYZ7WHkrT
x4jy4oT65Q02D5+YUcmVfrt/9NzdOcBfudejTYcul0a7RVLyX7Cu8bd3G1dft8sY
5fjcGWq6A/xtfHoY4DDLnQArVs2L3AJ4qwGwEl+wcNXbr+8nDSYVzowjsP+0I+/n
gFy1B1sHoRsr1P+B/qf3Gte9ekQTEVzb7q8AZ1smNRKfgWlZBhb9gjjymPq7sWuk
fXe+k9xTHOd6lwprMH2eWkX1QhyIB63JkmDtdKedZg7hAfhSUzeN+u2z7r5cW9LJ
1CS2wnFPeRRUOosxNvYLjaME+G+2Ea3uqEGjJNI96N58cJjcav17TENniu7+80aS
apNDOfPF6qjP6/y5V3MFt71YbjOZUERlMlYXsh569bZdyfoVUJtmPef9GcQEWNKr
/AaFO+ObPaqYN1lwkhMT/7yJkmHhrq3W0OnPW97AioxAIkDVW6XDlfV34S4HbZib
l7AiHHkiVfdn1NIAM0uZHQdhzwujBwnN0wsXR4Z7jm9NzTf3t+n8N/IE9g3zG2BJ
R54YN38uMkfBtun8HQqQqnKjhE9+kkE8heougNgD26so9JYHQnLWUhLMqNQLrC26
hth+3xSY5iZfEBRhJf9X1Ntq1fjlNwfnBP9VDLYyd/3d+lH+PaNUFkwszKWsIT8k
WsllhWkhA3LmKRQlvl5b7RGQ7yROQHNHdwT8wiiofSVAgx4gVgeuaDqcLPglA2d+
qzgsxjwyb2NtTDTmYjroOl4gjPGFVAJs5uzlfBZOtOQUXLQwM9NExbpkJNGTIZPD
+DVD12t7YSADtm4mEmsn5dQis6pWxlXPiWF0fXgRiQ1X8E5X4uaRkh71xenc++Rz
hM6PzBT1K1+KcVa5ZnCZ1EZGQQypGaG+Y/zoffxP3i2Y7P3y2fWXvcDTN/IsAcWx
mSSmQRKUEdMmbBZnDBnIl0XZhPTlgmYjXx8Ma4v4dVBvMOWpIeM2d3mKPazDLfUf
0BFmTyE7bUrzmvIuLVghKJevzanyzCFZHDQqjaE16G3lWz6h6yavPwa7I75IDW7n
O5lQYCCnmKso5W9UIXqJd1TPLO1rCvXR/Hgm4ZEcXuKUbF3NAplcDMBv93IpYzhA
LvP40+MyxroJBmhhrVZGz7IIZADL8HqbqbNHwfiJ6EHqlEDCiKPMu6w3R7LAv3Aa
UVKJSoYTK0xPNDFYipbB1Wpy9indR/W3R0Cuoa+rHjcImnE7Azw+uL6me8+pp+Eo
O5cxh6s2lgAqEk3leKjH9FoeGi2iZczc3ALgwvQVl5jDBasH5r5k9u8sz6pbgkOX
EgIAZNOnuqBYBSjsdGr0A+rypdQHGeYtjIdcDgFvKReQPCPg9sl4I4lIDBb5txgZ
jN5JbK5u1vOzMovX7fgP94eUnEGTFZTwypTsNL69IxeucfA0GyrZieF0CsDGxc+/
DtcT2fcsiPptYYQaMD09VvwY6+YoTcBUssH8Zp3L8uHRKutQfU4lkfaOdIcRt3Up
g696KOI+ZkaX3xyWLE0fpzk7yd/Nt5enOoRbTlcdHpMZaJGdsZreEkvGrm/e/RTa
v/Uc87w1L9UaFdcyZxyu6tDnMwg4Mr390pimKR/9aiC7uHXwy1bQOOwp1lNjseWx
vetSGEUkVCN92A71zZqAGV85VvUY5Fwh0cR9/8cG0ESapPeCMeluNdSuD2bytP+Y
eSLcNaypOntpYMHh6Bvzgt9Wz+AbVGCn80uYbbSJ7Vy03NMYpIvJyjOjo1Es2Oub
C+buuPgwtu5pyG8z49Ya3LMqzn0Ys299yQeb/mcPw/HM0YDAXbi7XhoBd1SHvTDi
ldnUeP1VFR6gtYtLLPMPbieP/br8mbOJzZhG50TnBjR3hycx4JFdHXoOyC36J1iZ
QeYRBih/JxQnCuh9ByCctIs0TyPc1D2UaoXzrd2vHdmuEHsQHSreWZ/wgFp0on1d
Kvwkf+qbOrXrGurhnAwlxomn86ymGucXMzuuXe0JKq1vQ6HyehNkWszUs0XECg6C
R7TAFMpNgumuKeH2aZSP5WuTgLx2ow8N6mJ7qNbLVK5CmPQTrD9Lr9fUPK/KtvHJ
S9agwi7Pw4Ydivx8Cmn0ornsPlQ4alP4QzTYU5c4FgJB5SDtlmoIMdDLCL4GNWZg
kY/XbNZmr1kQKdCTp5OnqSrVVjG7r5Kt070FpNyfhn2WkE/Ia+etNuduP9Jczfec
uX+w1XoLM0b9S+IK9f0GYPEhX3QbgudJhUAprErh+2lMS+QHfXZNhkcZ4um6F6So
nQ86BaEM5jCcuFuYriJ8L4nkfHfGuPmlwAF0DJXNG0MG1KerGZ5wTmOU+SH4yVQ+
PFjhu5zr82hEW0u2e9h9mVVDgWvHR//uStH1R+Gh5S4rQFrNOo/C0gK1d/IPTf3S
Ho7wtLmCnhOZgXCBQ893ZWPdUup2s9m4d9XUkoLMiSxnMYzxPXl8Y9AXqHgCv3ka
2XWOb0JMStZKj0c2608fcAP+9jdOH02z3XhLNbd0zJ5r+ffKrXF4BcmS7ek+X/Zw
olWAkF6dK7BLU/T514deYwr9JTthtCoupEKW14HPnHSKsHgh7Vxc032jVoN6Mraw
VDNHj9LrvtGaqKfIO/DV4NTNLuFaKcx0pHqmOllTqW37y4BaFhi6ZusTf3jxXM93
sfbjU21Vf73phZS2nJEPyzHkE35W5x9lq+lNW0Za/+nn+yy/B2dRxc/L2X/CXMIE
Biq03TcqCTvC/2zxvvtKT5M/yzclZaaT5vYz8VAbYliDl9ynLOV+xwrAUzcokwI6
8IsqxvauQpRle7SrD0gxmSsVDQx9iLzauTRZf2W+B9iO6ROa1TryXi25XObC2DeB
Dn5DBgadxYd1OWKP62yLe3GlC9Ua/FPLHFCWIVHlqpGrn2vNEVGPbMk4LN8XZYCO
YGbZG0I91P/keYDE80t6nuLMuhe+rL2+l6xJnyu7//7HNl+GPx7VdFcljAjNHiDk
5v8qAbOg7RxPLTUJ1anDvwqaNRvvsLkD+HYUkHHi0+C9iyoG8aWRy926vnm0Z6XW
KdKIvl2FLHpk2t9Dx8kdtWxvwsLqBQNxA2UD7hYn+g2DM0eUjW4sGr0RYudsZLod
2gjBr5Qgjgm9JlGmmM4cfh3Kz7ZIGg/udwHj4s7/81nts9pl/NpjZrEh7vQgSLip
LP46eMIbEAK2c7gvu1yCbA6PT6xVPha2Eza7EsAk7GyA0sqkC66rYrfZ1T5hBfV9
GOCHxpmDQKRkuE/VHSd9CkkytHr0KTpJ/a6wCVt2LkDu71HotmkipYPNcYdzE8oL
RlRarGBzNUtMxp+vTn70oPs/hJ4TgYNvzdZzDjFEmkmF9Si0m5qeYEPeGe3gmDoI
86ufEgI9roL04sbWMokIgdJjbDLtAvedNDzUba2soXrNPvASZ6x+IbmcI51wWPky
oduDeeMKh8cofqW+quMllUsr446hlpkBax6DJm8c3SYSPHsC+h4AjDtslmi5Yalp
24NQIM4WytRe+pXWZDn1aHLFSvg5IlXzDyn0F+8MsLVeQIa1BAiJarDPY7THGIF5
f6YeE/14JVTPvs9OhcZMmsttVv5phE6phbcZYSbWxc4vnWmUE8Pf+727cLn63T+Y
kv1ZUhDOcuAeoCn84TVAMK8Uf5BJ0FPDTJ8GTFo+Rzii7oEggsuDNE3Pp1vD+E9o
vTxu5cL8OvhgB+AFbIDPeXVqxnPV5xUHBfjs9lb7dwLi4fHUmlH2vpmBsNPHV4P0
RmqkXVpk0pO0Yfk/riuNZlnVIGvBErgWCuVjXc9IH3IzswNEPmnsfEA3QYZvB0q+
Vr6Xx+kW8Wki2t5pKezfO4oH/YpI189f/jdtQ8CQsiORfLZn9fm0qYBMnT+wZomu
tSNqiUcEXUm+8U+WgAK/5hokEG4OlEIUgHbxnMEsfxmuprS/J54b0wD6qg+yQZZj
EGrc2PdcfnJLPbD6ivrtBe4QS44+yZ24MObVzHgpj/FahLXCyn3AKbYO0ki+kGn2
UbbAwcPLPqb+CwPK3J00lB+ZDbqeAM2VLFUF6e/rWZmMCnXsxytd8wCKOzy+9GbT
02qytM7swX5Pe+IMnZCqQcevJjtKaWjxRBbEBJx1aV+fJ2T52HxA3Jbd1T4dfBmN
V2ENJGKLUrNLz/rx2WQ9rvI5Nz6CKzfBVMFYFmnO5baSLzDk+XLJJc/HPvYNvPNm
4ErmoY8FtTmiZrIYGv9lrFqLnMkFmTKEke2ju+ZAITLRHl5pvWjkQcaCW77LUatM
YvZk/+LBOWSOQUJKKEMMmyr5TfySetBGI/+3KPNSYfNjD2OKaQ8SwsKNXFNcYdeK
nIW/jeUQi0A9bgtpNvS3dNanlcrhriZMdVt660esGEKomw/7T7oAVa0nz6A+hCCX
VutPzq7+VwdxYyhJj6g7TlvG1xGB9kV07dpeZQQcTufbusm/Pap1xP1dwSrZyd0p
lCd558EK5AK/iEdsq1WWZtBqr3z0YImwEXPDHe//LY0u3im7M+hSWP32e6mwPxHj
VkQDDErYQsjbelcTUJNHzHeMRkHymdV/G7QUpWGUUYNVZPtNlgjaSBNC3tNHL/5V
SLGkSRcTgWE4BCtIFbF3WdmhJ1GkxpSqcA8itfvjrnIyts7n97Ts7HT+ZeUAJWGp
pKwKyjie9lH+XxUeZCma3zZ4LkXOqlFQXSyHoJ7QSnnf8hxsyAEOk9zgzMD5jPVr
DTlF+hhLWYKNJI3iAb5IL3vQwFB1VsvYxY4u798F03zUqh3ePmFDnik3z/NTw1cX
bBkQHaz648dUKRC7nzGyM04nEiJP5+E4266AwkE/c87nHMcraJNz5tH0aQ+CulqR
GkqpC/cIQA4GaYXpJCRSnMQqQBROk0z5Imnwu++RyFEHVvStL5T60BdbnUgFzQiA
ULy6DLSxuynQ8IIR1V/d/yue272KIQmLxpaKa7zHbRk8qVdtP5odbr6syizFdGfZ
JxjS4f8g/A5V/AEojy8E6Qg1b8QdXVJ9+EEb4HlHSzTyodoZXWr3gHG21Jm8KG3+
nqktCdi/Di7ztE9D7P078BUgK4TrGsmUNBia8sFPRLSIyji6Co6woAqBdDQnWDWs
NTklbwrr7Z+05b/igaeaVd+mw1dqs7La+KklzC25EUbj1pYeBKWyVYvhnTuMlph7
XhspcxbzGl+YtD0+PB8qZiFzj7nDrBK+NJcS1Fg1joHCphySAe6GZ8EWyXFvM+3B
BDfQl0AgqkCAOV9jmJcZuhlBgfIdDG0buDPzipLx/bmOi9PZT/Zq2kbbtGwyDrd/
IGvyVCWRJERS4gkivO1czSym3DnyueKEltukvm559nP8y8XNbD0nFynSmOwHK5qF
RI5W4J7/L8m10B4CQYeiX8lIwOXx+zdClnpjveYnvKLS9T7EXBa0YQ0qbvgZMftA
8pKRkcYhFRSt7iCijkbGE8ZjxzJKqqEnG/cfHterjitulIU5kEKzWTYpuXjwoAse
PQDlNmHNIQiVWxAwHzibAAKbLAb3rXvsOi4XLARFXSWSST3fuF3qKqZzob5LiV2j
76Ybq76o+yKQMWXiykeMGBknfPT5Po5gw8OpwXc6iKfDQ9wu+9PUGkmoTbRfXlPU
PDko2enPn/qtnpOYGh2cMaK1vKz998q3ZmOzHh57FS0+zztdmugLTwj++0Yueow7
25kqP6rb2fMrf+fyXFLWjSAk/SBstCqi7xlDUZAOBSYWcA4ju17WMOWMdi+FtllO
bcH2zBp0R1Bxoq8nRvNyeGCbcL0/EN0PXfqQpdPt+UN26slrBTp3P5hKV3aCftIQ
NzBKl2+aelT0CE7dOlyghQYcnDJzlHajjiSdOFuhBDigQQOF+rMXQkgmzGROCOWh
h66paCIH/TsSmHr2+ItYvqSWD9CgzY96GNC9Hd78+Z5br86hSP1tcNR185UCxyen
o6kO9imDMhL0ooydoBpywqb4YJ9GCKl8WIUfjrEETAo17MPoBm0Y53aFgijbp/Yh
ugkTJmxgQAVnlQyjuC811tS2gVhgjQwj/JrKoPVLBkwzyBy/DhzMBfiR1FabQLcW
Xvb/wL6UfIl7vUWg0fcWYiBmzM8u8vQMD0X0L4+GqyBDpy4/T0a0AJOUNJXICPr8
GbKchKGkNc5AF6K26Q/EEde5+3s18Utk8BJtKLGdb4N1rE6EwKXt4onc+nfEwC0E
pSj6lYEFIwjMCj2i2h0D1qUfTHPGqMcnRzXxqfrCVuN+rSXtGaayLkkllxDh+NeD
SjmZp4WSfibY/Ps4pcQQtq9/Y8NBl2WPYZwO+Qhj9EMZdoOcOBXu4RvpChEjETqy
Fn6IxQGKObyJ/QmgGPpF9aEtPHBPT1M4+BOhkG+ERRCgGjcWYRXgBNaI5JW3/+/f
IWmejZE4FeyAIBWsXhXxup2mJ0MV0qoCK7rG1i9yb+j5WTrPutdsGcSnsQZIgzhM
URIFewyjlvpvdfVeo92KaxBdhTho0pEK4y7rI+YSluxeffMrX34Wqkg/fjTJUaXS
bEMSmMCHQobNzcc/pUxFBeYHSgPJTBRj8JCnenJHbWff4y8YKniMmCqEZp55kJz+
cEWUfh/+WSuBP3B6Q5d37Xi4RU+2fqTxmBmxzGfqf+8su6t5TQwOLGsie9g+XP+4
Md4yFON27QrhyhR8ooxXxe7rO/KTCQau9crCMEWQN9nE5bHZHq3KvMqyQVHFVmC8
g6Dp04IzvLwFP/0k3LksTc4oRtgh25oKCooBs/xC+MkZndBWcjLaSi3GOiUrVxVe
GSQptZO2sGR9EbRcRybpWALUGgXGl2iI8MMKmQ2UsnOGFPwcrrd8i98IimDHp8CQ
b4k+mYtq0lcUy2zptCQwKGpKA/8VUtEVfFUIJOnNHBZIyf/yKNYJiC/mq88HK4DF
eTnz5GtIKXvmzqGT8xmni7wK9g4FE0e5dc3vF9eMJ6rxT+CxHJ5t41T8kxWS8AhE
XxKGGfdgFX7cD2iIuUeZunGlP2ENNE/X9GrJWbt1jCVlHuuanuHIkwlbcJbnRuDn
ZhHBfm/ZrrT0e2Lgxt2r71ctUa5DdeB1OZlduS0GWm6buC+Ap150clv4WwO4IFSq
PLuQD33dmhXZpGfdI2psGt2Gt27fsNLKOrIzg6Ij/mlcwNkLGB0QMbzFtMs2X1y4
uRSlGNtqIyVX/YYr9IKa1e/0nO99MbaHdRTKw9aKiy0uWvzRh9zdKEl/jTTxzLbU
CuWkMfrLPqRrBzicOHFp9WiZ/M+R+1wJuLCZlxl0hoPS06+BtLJ9yuRZJmHK6+c0
FqnZQU+oJYq9h6MzUUeM2JIUiP3g3qS9ZPJzm8X0Ub3flhgp2g1x7CeGKFZo46Pa
LVkNEaIv3XJZ1gShieAV4y5hy+hwJGdnQb8UujD7AG98sSHX2lBszpUcpQrTQJdc
GnE1bLuWtrrJ90iGstwsMgcfPB1+AmtT3kA7ISI8+b2X8A7nJf3QH8v1Mka09raR
QV5OI9OPOqRe/IVxNa72g1UmYUCsv1GhbOJlv3MXx4yVXWiVOp8W7Te8YgcOTYyf
FShAr4DvOQZEMXuS+ZeK4HxqBzW8BHkz1oEgE+p+C/T3dAY13boDilnUH0KnFpDh
hUwJoohcNuCBPjs5ZZbPUczDLeJhttquFT07Ca727yjxeVAt86C7S8zXMfT7+fAo
JD6RT+Z+PvIUBAv0NRFed++wA8ONgt650F7wwgF14dH9+Gib66I5CIEUP+mTMvVz
HFinnaBgKpSlqO8+SBp1YXqLpPaY6DO1txjBbdGq0AtpPjK17zcRKfZJoO4Kj2cl
KK75RhY2CctMkPKbX8ydrG7ZfTxRYVWZr25XiexiSLR+VegOJBs5AmVj1s7o5+N+
+91FquC/bc02iJI32oWDAsaY8P4S6jRWju9HyWOCNl/SZ0G6jTZYjp/ibJrAB1ZN
kSaHcTGEin5kSMzLoVPnhcmrqi0JP76TH6GVa1DSqmOT513hQpp+kmfTnedqxj0W
Oa3QlM5ttVDW+2QTxxnTtMJY71FQHl8kdRnHZVY4w8j64WjmuqVbiRtj1Za2IBpe
tsZas3Av9VEx52CS0I8ErBabdsf/BsXP1cQ3Ts/kjDAoPna/gQa/zl70P2zaJpW/
8mXpd3hkodnYquwA+qiPja48OqeN/xo/igp9eBIHOJzmccikrtfRFxIjUBJyoHZe
1ykux2fgJdnoq536uSgrv8EjQVrn0v4AgrgZ3iE7gFcIH4EyzTgU8LzFSH39G8VM
ROqqrqgtEhDhQgETJ/xVYEQ8i/nqhQZO5BPHpzH4zOqckNfDIBcecmKmww5B6ioH
5XYC9ZnymVYOmFOiF99ktvZaF+89rfBe+bmk+sLAcrKdGpRgDhmQ9fMCie3zBZSm
kBCOXCjAaRAlktgz1U5Ciu9Qb8mfXM8vlpOuL7/Dr2I5+wEG53PS00wzRrzUGYse
Cl23SAp28XFiZ5nalOBwXjxwQ2u740pHI9ryTgN6B8FslxUGNFv85/oJhNNiNxmO
eC5jR8Fn5wLFC6fqEY+/hsEuIp6hLcaocmLuKmp2SiZbAPAAyQx0GGDh8YMVWWvq
z+rejUK3RZAlR7Rw0U/AyiL7CCdp/Q8JL/JDkBC9QWtAjBMG4wCeY4/v4TrWCmDJ
OixL+UfUYoEqw0GTb3W6k2ZZbYyq5fUC6/xjVl/a/EagXpi/Alvh3Eme/15IK5qk
izcrcOrTyZOvAXc5liFpGBAbLSl9ZyW3fQD6QhP03N3Rrn6HnG8yJTpRIGnz3cce
bjPUL6DtM/rcF6w2iPvCq9H7EEQl43Z2GiY0Qvtc8H3JFh/E49RGinId3mg+aayg
wt12zE1w52xbBrmk0ALUdfZ5N82vK6jE+5bz2RDmgIZ1qwqPqlUaE3c2959d1i3/
v5muAwmE9a/vRFD/Wc6ES73Hbzz5raLtmKqHkExVKlS8pSMIwj6xwTiUET9dhfwh
1CN4nc3UICP/bGm0P906eqa9hSqXuRQXh7J3levRCESLpNRPxxk0Dkty8PzaTXeV
Q5ctYSAYDjVw9ntCgtDpySXyyNAbczSJCewlusIv5jE8C+ImW96NXBh3KJ/Qg1vP
OgcONytN/K9jCsXNT4NnwKgqHtxab9DFl/bWZ2Jjn9hBnWRtCZFKLizGS+lzVTi6
zBQeR+sR3xYPXpemPqXEB73Hx6ivUezZJ2CXT226cTpt4Xip5oU7EXhP16S18/wj
2h75eKwBA44s3tqjCmyqLR5/tagNJAKacAnNMkxd4PrbpLLlIxwsoGgBcETMjr2E
YR3n0PdKap+iux+PHkB4bWSP+TnawgYWYYVB7Y+WKTiAGGZvPxa2WrEl+PIxxcuJ
n3V5zDeeYl5cPXdEz9+cD1rN78+1zntkSkBbQAYX9+egCy9SkQJHKKMh4sg8NWVd
J8JC4smhLgLe1trRW/l3iBckUG7RewyxHOt/8EwjSXHQS+97C3H1ZHactlmWU3zL
542OmrtjgUIApwS28sA7kVUoJiy+RykDGBS8FDqlNVS7mZCBbb9Jqmbz2LkRpRES
pCEA8ThMIZTXQhf8Of1DpoB3M4PoWC7FPIBX2F/GJQBh96sLeXXUKKKcOdUU1u36
f/a9bAxfJ4AsEAids8+0ZMRgmEcgxN3UNsO2T3P9dk56j1Z7BmL2iAiKvVvSKQzt
TVUlGhvT4QlIM+sAQGiy6Uw9GTZI6JKt6uYZ/PiuL6aFzE7+kAjRIsJJyErzRzF0
U8N+6LhyLiWCm/b9pi3U5HNNfYb38yBxxaCY/Aas6Xz4hNmWA646v9twShhs6A8h
8x9quw3UIM6u0s5lQDkJVwkFiNJXem+kf09i1qAnhIsd8USlq5Q+K8XjPkozZgNh
EMUsI0jMCTNEEbQwzQ59FburIs94uEvUpyo4lITwfM7krOh3xfN2e9d9rn+UxWeq
wTqraH9YeeqIts3dHnVRAvaw8M40EJsxzyL+xYHAxEpG3mULRTRlm6XXnoKRBEW7
KLhxKw3hbW3k+tuuvxzZpxHPcgxsDpnaHg5GQYv4Z9u2TOXjUOIxOt8s9rdHKled
i9jhCavR94momkklJ0UR6+8bhVvztLTG538wWAHh5evhhaFSxCv/LVROSXBmPjIZ
B/ttXt8yvG3Tp2uvuQBTqiBDm8Z4KcCChx9iMlSkW4s0KLPQOgO3y8/YNAK8LhzO
B97D4v3WMJSl817ywF73K9WlMso3vAeXPnyd/lhc9DT4Qm1QZ0TfJ0AfZXbI7Cpi
aj65nwVrJpptZ9yP9bjVCWqUCFr4oSTu0vqzK+JFHUyceRHdONkckeHtNCeX96Vr
LDunt7APo7kwyA0Z94OHde4V+ikTrhbvhe2xM12ol5nndQfBMjfTg5P707YAwScC
FsBkEc8h3ayvIMNfY3LDMTEtF2+YOKEOV9nu/vd3HVjNz99U/6JObA30VUc5RQV9
oYUJvydP+dWI6Yj51QrV2jgJNOh+CGhiggLcGjW3V5RmfKcb96QtlyHXgoUVvrqg
1uW6TVvEQYoBOBFBhmEuFVDtwaB3WAettruZMf4guKtvSyMkbEp3JofqsY6ejBiy
8Eh3KAbYllzM9iICn9TPMIF7tjGpXlNTIlIHekGzaImbA4GuCe6cA9lCCMqiNwok
3KWpLHZl/CM0gDoGlIS/EKdiRA8rqwGCyC3lGXEQ1mQMIc4GZN51kw3WdD6GqiF8
G/yRHf+6k1IqVN1rNNC7o/nCIXyPyB6HIRXXPoDJTdnZaRagpWtwLe0UK0IwFqZN
oyODZf9YeyCdnIhaL98lmlzyfoQXt2iDrH+zqX9JhYF8e1WqmHVk8F4ulUuPX48l
PDZaLFoPahcbuutH3DaEyLsWV6Z6OBHA7Y1lrMqF4DxF9RTb+D0e9IKa9LRTVUKF
CL60TI5juribzW2+fGMm961WBVnYz4pCXxhZcHIN32x8aO0nJz6F36UXOxi1MJDc
Cm5kkxjctgQpiglByFKJ0SQDm6tblqvE9pPLhdYwO5ABdLx8+7ZbIr8di0d+yOdY
eueDAI/O77ityaE5i2tAn48JsNXC0HoiZQjLHp8nOPVwyB8ofruS0nLDaRXUx8m2
LFfuj61PVeSDQBXnQRiNcjuJ9QPCFv9paF9tdQimNWvlsRYH+55WcdC5gtZfoHKO
o1tBnbBGBqnO0la8kS5J88WtiLSVbt5e/7pGXE4fAx72D3rHnfmRiD7LOIZWAkHO
kknTAMyEV9OEedh0RLr0ZJn8uzJj3NoiFDeZGL7ucgjJwyziIpXoljhCSQMH34oo
8zJshAdWaksQAxByv1bpsuKj00MlUAQLlEA0r9Rd2c/Ni8VtJv/xSjijRws3Tr6w
lvanfbhSZzz8EFe9sWTy4zr1y0pcVfpK1mJx7nsSyu9yif0XYPH8mhu68J+yhHoa
V2/cO7W2TRMo0Jq/XXEdj6DihTifsTUfJMjUwPdbM5T9tEJCAIx60a2QdTR/Nj3X
IX6hdNHBMlrPPFHbUppGQXU7bW5ydAZ53XUXlXcrUG+5epy/qhyltXRyWlDo4AMq
GXHzcq/NYL7ubP7kxC34FQ97jscOctlx3sn+P10NjdHhwByIjvnaY+V8Hbm1AQwY
jnCLkHc0WUA+bAteZnXZuVBrQFFU7E3Zoris5YiTEjRjOjB4d8hAuWyFuyUO5yn/
8MzvVeKWmMguTRRJZ9UkZ69R+1SvXbyUCwABM/07YXq8O85exNXdrJ53oFxADS7n
P6TegwRVylf67mJeI5BvaIecJS2CD4s2ztiNmjZgiqHN/X1gZoHXOi7Zl0eqv7wA
au17OnodLZzdeYU7uMDKU2eznL+naKzhfhGZtCxu2O8IG3gb4Aj0Hh7iNhOLZtdI
lOSzQv4R3IekwknWJzIRgWZEpOjUbrHASNseigNNjjlUXgAfpMeHNUlVeCeXdSIj
ZoR7zn5do41N9EFgac+pNL4q/Cz6EyEdk1ePPhizyRFxtMqsvc+r/B8qpv9PVjXG
WlJ7+lkmB9bSyk4rxlQ8ye57y2gvzPzZoCmKDXKgx0AgjO7B7bNJxkCXoJ49sKjQ
HlAafS6HhJB/b8cUb76HwFNccUMCS7oL66/+0DSbb6GfuNW6MG28oMQBf5X2PQe8
CYFLwbwUfBGxahUYrxZUTDtHEroaIVS0M+Eu/378KDmS8uvvavkJaYIU9nrhmZxP
OHOP03GiF+Np/rg4nkfQIfzVlVUR7AJwe88Rx73I4Wi7D/KhUw4xp7/eBWREwgOX
nqBzg3BNLtBIoDrCbTdqssTgn2HUjxRlNcLnERwRYhybtMp6p+JHan4ZGaONLyg8
vm4iaDnH0gKSL54iPFLpwUYbpzTuInbwwfjngtxjI6igqhu5Fp2VVSXIyLo7AN3g
1VL3Ba7BxMHqRVTQVRkDX78wLPgSwwpnETLcnCLnBSDPcrVWKDfV/53sdPJfRcGd
ZJhfwtMTheFrXj65eEJYPS3sCop4F2n4X4R8V42ehO0yiII8+/Cn01wnunwM9Bya
BhTw5yUotaRcaTSfF0uuli3GEkHf9aFfTdSuw8dp9UU76hKnhhhgNHkxF8PE0jbG
AZNQHq7UsV9bDNyMDmTY1fzF84Dr3gALcQxG5E3k+aEAy3ZhGvj/Q4lxRV//n2HR
Q/1uIWbVk+lVzwE8aWO43RgXNaVvuXG4BcVj9Gpfr2s4NYSVrH1A6hAFvS+O1jAL
qq7cy4anz2pQl61mKxh4qe96BrZ3ccqv37mD/pMBbU+usr+/Ck7mHLGp59pynaKO
M87KlrEqbrsQiZEoBbwX4alR9x8soomC037UaTVcOyLSgSYxy83p6OWKA1Er5Ued
s6qQVARHTkfVBeQBrTowXOl57bm/MQD5eFoohfNOgFvPA/N0lBFg2Z3ki/c3yyQu
WbejSnhD3i7ChB/pA6OI6y5Whke7brF3aifCDeGZSuygVP21c+cKabbtu2JOVnU7
hfSxuAD7CA52ZaVDtVAvfx+rRC5tFUq+3ny0sM1e/0RTWPq342ia77/aVEog6cxA
uqxA7l1GhHQEIUtVpQBUtoAGh59s0H1t5SO6S+fniqE+ziV9P7m4VrIZurFY8cB/
TbBrA0ijg9CqT3VyXaObB2IO9++vPmewBRQjbnqZSV15uy8XXc4vJbWZScXefwt3
Z+9LdsVzMEnDj8+HHHWUtc54ud5WVRevv014kcps5EbQHeogutFMbn7EAvhKCAdY
ALCGEncbfAqBt5Nu9zEVqegcRjSZpD9QOC19QlIBO3w5lZItudHzJdxRLk6aXWPP
JDgTjzy+BrudwwvJTUmbi9gPpI4zQUL1aQl3ZiOtdHcnMckhC7fZPDgZsYaNZ/0d
iaY4tGfulXpOFc/h/lS3mxK6sjvCiwqvdc26aCJAtdIJg08USWNzV5EWrzjahlWg
EAT31Vc9kl3yj/KfS3OnpEB65AEIGmi0kwMJbchvG71K6ZM+ja6ZQTGoe7YFXbWA
f0JfFMiBWi5q3SJIQxhU94LwFEcxARf52++G82nwR0tqciZba0NxCejgNUBWVyM+
hsLQVADXM2gH/3Ygqz7a1KZEQZDmyKdZVgJVoKHMCQb0jykpx0dxcgQZW9XDQM4k
Xd9gyuTSKkC0ZNxj1KzGKMM/MUrFtSsN6Wo99gG5ykBa2mSukqUoLwAD9+WpzdhL
2KzFR9VS+r/2hgIwdNEnbdo06hxVRcMuZHmu9DxMhNCF6J9cqPrMf2Hnv6+HzC4N
3e1rG0L5tNLxH0cPIzRembzzRM/z1yL+8Ri/qzsFkRASLqBn7VMSgWuY2n6lVRpu
uYd2Rhs4tRd5zlR4TYioR3K7viyCSPOKDW+jpKbC2YF3dDn4+EkyiEQzGyczOWCO
DIqOIlARxEKyd/V5/YO4AG7dCgvr7mI4AzI5WBm/aHR47d38GkWE5hVZXPpp4/BY
cWCfZZFMVUXVlZyMc2vbsoTQPa8cMy4VNloESjhu1htJyrkxOj/vc420NW+daCuz
hAWaVBaWbkalVlG86dc77zDTPL3SQmMzdV4tExHD6pl0rVemFDyXH/3YiDvRqKiR
DLn5lFlKrH8lOQd5UOCCwyzNsLOkdqYqTXSpDQ4X1LB5GK+jVMbx0PsTNblo3LzA
SVs8BzOlhc7t6sDQiTojwXRQXdtBYomU1kpaFIh4gb6rFo7Gv1XwmpL6f+FLMuuo
V0+3ZNyDXUldgWEYhkgcnRgPiFrwrsCvze96ahdhzWZHCnk5NzDeSStxadxhAZjE
cDU0eEatog7OGeU0r98A3GNFQGh+ywmM2GojUysIKGSZgkiAUC18yu+K11Zl9UZr
GZozzkGR13i1Y/CGewQszfAlRe0cplGG/sYl5u9p5Y4kqwMwyDPsEXv1vdYu6HXP
EnmDRQ2PJilBAgQ6JgauE7zEsOMFVLhIwVAtBKCcnKNRJ9+5SCzsqiokms9tBLuF
Iu36FsvqtV5eaJxiB/EMJBvj+VWR6EuBKCmlOUizQJVX6OGZZV9ZwR6p3C5HW2dQ
2FpSSYstmp7mS0CElBlgpFRniOo7Dw1WjIq83He7ydkgqgDwsIrTuZPPldNyE2Oj
lTn6ad8d5bxe5Fy1iQr2w7jctqePNn/yE7i5TQJ3bZdAwmte22l3pj6JwWa7MsiN
atRmqkwcMzs6IGsOv+nGRE8FyXuvUME67MqJnz8chgibTsU4P2ehHX4LVUuP6kPM
SR8n7UVueHy0k5GkPc1KugdPXw6alvhGXmfisHBfi3t6j9YOwCyyKPTjwdmGCy6l
IGli8XjmiWJmZiKQj70t75p+Yw9kksXO8xN/qXvkzjE2NbyI+kPbkx6Sh7gd9OUw
7tRmGk1oOJQQjb2bRaz5UgGYRtbdkfiZvaT50/nd3f6zLrH0bw/ZVQn+qB+6IkV3
28WbSzSgD6G7WvkbZhfdpBhtaYiEH7ISQ2ki5PPSI/c3NzuVcLxnhLNlQfhNEEhr
+KbBg0stEGn4ArNT1+cQqtTyKMA+eFEOTE9ua5ZBQRBIZfPFX+Zm1G/JW1bhNv+U
o7zKozzLROheaVkfttlhe2nmLmfOvByiPFQHjRap51xCR/gwRdI4GFg41AnIxSA/
Y3IU0Knno+clI5oHmjjmD43FcdJACxTzARNWmiN5wicrdbiTG8UeC+ue+ZPLzD+e
iUVOeuFcjIGdQbx25NmFslksTiWSsl0cGWTDoY+ucBzeKh3lvosJBVUw6C+0p4Hc
nSOWYcDDlDsHuH2EPUgxPKNybyXom5iBW4KDldhKyAxZqQ2kyBu9WIZFDw5FUnLE
nwuG11wVpzIsHCdsWSfcUFnIRUAxVTuGc7p/2Dw1C7un7lbzK8qcHxxV5ooNcYRb
MvktpC8i/fkzPZal3futVKrGTrVaFtibFiYLuUaQXnlnB6oEngwPaFIMKx7JlaEZ
NaeVgtpTAJh05gNGEsIhFsdeczEXgXXPnk6QH+kNGbNsDJ9rMWBwtuOAFfeFr4mf
xBGBU4s0WuVRnMk3sMwb/EFj3vuqR2ct8c3GbIwO2S+ss/Jy+itASuaDZwVFyEn2
vYMZs/puBeQJCSaYcj4bJhmQ4y0K0pJlMYtPB8OiB9QwgFDRbcDJZOwVxR1AVIPD
MHsD9FhYjHa4jaC9Hv6XS2VZbjtORpp6Qv53Iq2JS9ST02jdb5Tc1QRMSpYfsDwV
ZD2j0St9i8rVZymeTz12AYOEvsKSYw/VHQ/y2TlgFyuguEAtGiA40DFo1PtQO/l8
xk4GhoGpjtKpaxMtJtTkelXnCLzruumiJ2KmW6l105ssmezej81n0X8Fkga32jyT
CwNQUUNJDefeTAn+o3ppmu5q77CXvpSp7l63BW9xy2J5mWF4HwYwFqPgHRmkEBln
GT68DuLPwngr7c0ED25mDZYGe/au7IMRG+IPXUBZdYrX/0cC8GKDfbc5HpaZjTxV
WPn+WrrMhmFN4vE8iOT8ajSeKUUh2OuER+vCQPpgfqk+5kSGBs7GAPI5+y5FqG0L
rEK9OLz1S1StsFh5ts0pCTiBIxXQA7FvPwV6/Fs855rwrmyerK+ePHH5GsiMBUI0
mViCJ/2Suy1UGHexCY06vGO2wd7MqxcuQfZV7o7VTELOiAUHVWodiL62FDwqE3/l
x5ErAyG6YZLSyN12/9jCkO7E8WCrAVhia7dJD6vUjqYl6qOh4x0LMY+svhGG7NvN
sSWI6+J1X0JwQFk+KQFV/GjsFlNWFSwphXCocP72Gq5c8LXVbxzAj49BWofrsWXb
9xCWCP+W6HAWJKgtlVtXJJh4TJ9UKgBPppuLVb7w3BgKeYKT39uxrfhBhflwntFD
+ELNn+nUz6Bnrvw5exXF6DoPQFn5KJD8fARg3ho7uMaY3nhltKaDgzmAGDBJ4A9/
txNxqh2Fn2ubeil+cklHt/V6hdoySocGCR5Zuq2GrBF1izBXJaR+c1p1lwFmMq8Y
DbS1NAYfDknO5pm9YvOplbqfVEGO50B/yhovplzaGXLiXzghmMznasloovklpzUs
C48i3lGCTKB+L8gkVODDhJelhzePIBusPPaRO9pVYqQ3Do52OfzfWQ8DjwPLiLPB
K+0kPcklcar0bsP9f4OXxbEE1ejnvp9lk7NzRqMuY6zevxAOK6t/3LhJT2OjcBbP
hOVXBdNbFntHwZVsC8vJBRiMqszQ443paE25kwsS/O32deSYTrqCRLZ9k8iNSeR8
MdLPxSx9iCeiEdLeZIB0SRRkqHNFkQfrkvkXlV2JHsd4suhlyLsYI3JoL+wEAevn
j8q+2ejRisdFpAPHtTmDe3EKeYLbqOGtLdkLV3j3rAlsod+KS2J0E+cVINhre47E
Y49IiV4AChuUkwKs79lp9rfLOBSf7Dq7XZC9foj/pcbvBzLD59WKhtwZ8aTgkwQt
0yBeuUkiRKWwHyL+eQLhaFJYZ3VvJWyVCyQVe50sQO4HPTgCwqpWQgy5AU/5Nizr
kHukZCmN0lOXXvndtGpdgfgbbG41QLQYf1ZPIPbrpmd/mgRVY91cGLSBc/lV1TQs
dUufLTVdZmzFGw1/9eN9lYQEPRgXoFbHEmPRVuR1bR0jlLH2iDD3/9JSJfFqcUC5
GHMkO0TdAha8RiXC1yCPX+AfHV5oxvWN/DR79Lo/b25k1ccdDx1rFvD4dbhWtSrL
3LGObVJ4uqyBZig15fNzafk/EX4BK+F9FpmpIF4ti6F/avPKBjp0czbdOJnoWInz
ChJ/Atyylv7bUp00ajz4ZlOxboZJIOJHga2gCUhxfEvrV4JTpsjCcZJI2Bve8wHm
EGT1uXe6uugd0DJEX5yZo/lW6QJzPunhiqFRIbfaCBMYMeJoZ6e03aitYPsj7pMH
pAchNHOAWp9Tg+N9xapjY8WbwZxY2GMwFulzz+mBrrk2aSdOJspusTg4TR+iWPyQ
xevP4tLP8f7fNZwZtzR6S18lD40Y8mGPJZhJ+YY90BnLoNbpivOqwC6PYYZeesGY
3nf51erwaGFceKfZPxkqJkn/sdf7mKYN72rTOgCUvCKSyUt37NZ5JXtDDt4RXMPD
vtjrQeALJsnAwggnHEL32TwFWOgJU2bZfWx91GrnvN7WNhbANartWz7fXkWOtBJQ
o1WdYjSSZJERuiEr4UQe4EIWiunyzo2Wo1H3J59JQ7kJg89FFXeCe7dWFuOpEsL9
mJ5qfBG681D8viKKi8E42+Oqwh0P6NS3jrAc//Sl51jez5zXLybD73oep16RKBKI
4Q58gMEpprhupUJ99YIVwcSSkBbYcAXuJKnTv1pEh2Inp5DjVw4uYMqWP6BXbbHK
0HL+18NJy0yJxaOK5TmfdqxrcxFQlh7FV86UYoktDEKpCNXJFgmynn+4AMcg39Kv
SvjP7PdVgteMQp/WRkovS5jRVFJXrplwCO4vi7Y/TXqC47sdT64//MQ1BjFfT5qS
MPIAZx5KzZ/fy2A5AZiTKdRIXyIjk9aQ+yfzc8bqgq1FJpTo4twrvs1BesCA0/ra
B2esmjIJyogN35mg1JnLUGlo/Id430sXp9pu3vyLq9I1jSyB2fI88pfNZtVFMwpl
cCdfD6/3PzUBgG1U3HpoW8Exwa+d/eGBHYTd1/gGvd1l9Kv7ZSCGPy6sgiWMoHeL
cDww0VZcJiKaM2xWlrcgapvarcDHxsjDd045+QEBMYGiPtc29h9aHg/s44M5XM3H
eh4jZv9u15C2RfxSv8Mp5NkZaq0YjUoowsDZXxWf3rmfbdw6OVAyQrc5BiuOMgRd
1Gogwj1XzjuXjYffUkA2E7IlRNxpWjj4kqeNSD4aGS7/HPu1s13TKyuajt6Vj+Yi
hFBjknpWeTGh7Hz7cLQqnetZkNdtaGiufRAHcRweRjRTlYoD8iQpTqJLLFWHON6N
zKhgKiKV4e8RgZ4dyWX65VjUoCI3WUBOltEq3rju5hhZtp9EYDFydc74Ob7j7ENO
+9XEH5zm41R8G9sTiR7r7+FrLgfDJYLXvV31cJt4K2DEM61+3pjDa7qKFKSF4YJA
3uPauqyBwR9ODhChvVDJvtv80Il+is6S0qPFHDQwseXBTmOUtQLHV3T50vpcpUAP
wDQu4aKteRqeJHawMZ1rieGy/xVFCfTYmsDgxoyG8jiqNeOeSRqfROUPMtxXTGUg
Vcz/F9PFH5US7L2YBb3aT5HLYwnxZR6ylCYW2rlYn3Q1J2CQ/VUoewsAHQLfGoZF
VRY2pyjCnliYBbHSWKhvQnCUESNJ52GnEFlbT7aVdMrdl/NeWBflsjyx1/LaU1HJ
LnriGExyaDhiaY+MpMDmq0NkVSUxpoM2Xyi2JZwvyO5pkRfTPVtIS2U6KM54g+k3
PyoF5xyuL+RZhppEuC08LRVYCOIXryik70jj/B3h6UJZiPO8nh8xY2X7WrFrFNS/
JciSiMls/tIRipSOt7SBYJ/8ne2/elyDsjupMXkc/2xvdbmMfGdff7fTPaNisq0d
c/z8o7szmMkGRBgaeDwIbajQLIHq9urc+Sx9NrlwmR11PlDpyaVZW7Fy5KhPgZ8Z
/nRs7jp4j0ggW0PhVQ8ZqzcXSpQKdQST+0PmzkG20y6fqSyglrb72Szle1V50S1/
ChkKrK7diJcj515HbFAReR2ZwnfJwVWEcVqYgNQKICwjwKgidLgRkMHUkBC7Eenf
uXaSWpPc32QMrctm5U1oIb1HwWz2yZNiFuq5JLJRbl7apcVArejL8o0eN3H92A+M
JrlqgXd/90cZGlkSIRjm4u2dVnfMHytWMp2EXrTW9ekkXpgejhfeO7Uw+MDs/Vw9
DPxnwsQVnMjj1telUmbCQ0lazYiMWkdtotVLQHq4pKcVK3nUOFJvdWMrgMaUblVn
q33y6/oHqtOtLbRvzahNdzvt4aD9oUjv6gu5MmyGE/Q2VMKnKXjTxw9bU9aw4BzZ
8AoQIFZI7jbNfdDKJWtsda6WJu5v3JV5k3atAut9nPju8AeJTShc7CuZCD6ZwIQ1
yjlIWhJWsB0j2ftmrzp4aNGUWX8FCOJHLWCwUqGfKQiNHX8EpRT1yxK0ESOL8gHc
wiEkVw6PN87QNM+Lwm73m3C8R7nA3dAJuyJouCJ/LNmVB5mk8iB/x6PN8dEBSzBE
FFSqEQjGSc74hTz40IFEpYKc1RjooLYPv0CpGcLi5Qaf7xZPV7Hs19B0664enCDK
1syUjSc3Wr7IE/CHo/MWQwrOmwnvDljLBfzNWdeb925LGb1DkGgep2sgp0ggx/WM
6gHAy3PoFoDiNcAP5k1jYm7PC8RpIGJ6pmKi1E4NUl8YLVpr/EAaZoEg+L+kVX+B
n/TXnWL0rvHG7fjgG36VJrUKozEzoyHKZOP1ZC9577K/rPzUhYFngwYbfrB61FV2
IADBLW5s1G7AkLM0UwFCyy6EueHbZAKQPS0/VgP52Hz+oVQKn+rGTQzZzgCA01dh
+sQ9jMt7IJH8uiOGbB6mu8bMqbETmPZ2VSbbYZlUC1a73xOPUQBoLaSz+AKkcAvJ
7lquTNCKvSCYUtiV81i2fw1PsF/XyL9rf9lKpLgHjQNPr/wshvnX5TDjnUntcseD
lI2yqqidAIQdFfN2KpeT7t9xgA9LU5C/C6fFnKB35ToyZonNSeOCs5xOhfTH17pv
6Cbnq/jo3sr5ThEncqykLVuLDGE2Cs2Q5S0kHZN7lS8ckgwCbf7jSZgQjiwC2UCI
wUhwK1oucpHgiO//RrjXoLMLCZDei03Ve/Y7SoTcLcNi36ArUbD01xK5SpuN8L3I
QIqd7LDU4khkEOyg+rClaBKmKz/MRWzbCOsxT0ESDpfN16KMRQ1/eVadZ4T0ER/p
aDiIugjbxB6LgFwiNStNMt84ORo/ynVilibVqdVerF082VxTjNcC7j+p2qsrJRwh
vyjVfk52B9YF2rhbQQiOE7N2sByJ2oVLapgiubsbWGPqfQMMjGcA1sFUtduob5fH
WnXdTTb6CpbB41eadosQ4WZAWXA65leoAcm+qcsLWPcYICWAyXppJYIvnxuLHYu2
S0RQhE0TfONQGOvPWRuBC/55FXZZ1Nvhc9LugofV6dbaxQ6JdYNKwSHsfx9MXGE/
wZ3/65aHKyd4tOrg15U41a9zM6FrROA7xl+cJjrnrtpevyKits7HeWISv4U78YwM
KtEONFi0d/ZX7hryn8SAxjMjUElESPMgnn7YAE5s0WihGjdmljjLsArl3oYfjgXt
Oisk4zs9sWFp6RzXP8r2rWhNvJV/9TX1htoWzZlyputjovDfmus7RJbb8Jvs54mH
LKhoXGCzmHFhUyZchz0HjdrUpAQoPlJeWZ5fqa6a1uF89Lw091XykM4xcIFZa20C
XXIXmWkvuaPsWkW/AEJ9jNtyhDlLKlwzkNbdCoui7gy0JYntYX+PObOqDl8ugbyA
TQFrI2nmIRZt/pHetYl4G+DDs8DdRGb8zaeYm4mAaL6rZ50keeFj8mW6KsiC7c4Q
v8sqIU8+PT/yLpSWn/UQYUH06Adfwic8USE1401tK/LuhfASwP2Xn3krRtaTYraJ
YS3mj/17eXwtg+DczpoQUR43/zmgEgu6hKgAvfrF8Tvruvsjj8eyOtER6Tuv45nO
8bMYmN0mVWgYH238e9+B5xLOt1MWjzLOaaXwUmz9X+B9IbsFEd5o6e/DtNghrgVX
yePeqKMSWo+WNvGCJ23GEUOtzFtNFByaaJwb6An6YwVjQ4R13xOsNOWlxcV6VUnG
oecuDfezbWPxbGiyzYQ22UwOmct86WnqEzzRsMgJk4kyxUeqz0v0CgKxnrBAPa34
9jkICgWOoztHmwu+e56UfJczYGCWNBEPIj1Fp+Ynmp3DgsSrE3lQ5ZWSfIrevxqf
SkYhE0hm+/Rla+4gs4frC2RSHfSw8JNDrmGIOpiLKSKFsTMJzJ1D9SbqR+PzTOv6
Ghzuufuaem0YJiuDM47Imk+IzX5g7vpalx8f5J3FcgruEWb0KW2tEm6HcuM3pKgx
1kxRGYgp/GSowYZd/Qon2JO7KyGBF7RbvjUDObcQRAwVGcX8nLvpcQp8NapTz/Jl
kedDZ/ZHUxJRwQZ507vF46P0JQic/8eD0jqJ/Rbl/J9Zfte2wEUWg/IOHf//rIQT
TIsygAOR0P9MvUyfMga4WYSzJLgSUFvI/Ao9a2fna8eTgw+q7+1KwOeYBRf0XYaj
/qanUe0DCrkVI/Dxrdzwh3HpbpCCLVSh+yV+oxV+3pdx/NMieUZYq7Qlni4KJT3K
r8jQ6DJGaN0rzHmH0kSqPCJaGcgRgMJiJr3kO6JweTVGHX39dRmjfq2UuOf9m8NT
ZTs66IPeZmI0VXuccAaSp145PbNBRh3eH/lMIAWTAPJEu76EfgciCrUhsXmmSJhc
zQIwkcmbPc5kb9wHbSC/Xr2CrdQ4IZdKw/Hoi47ABOoZrFO7UsJVd/d6G5w5jWRu
FDJ7ys49gt5VSALgESKudrPwQvNtLqcDgLBkWmRdVfZHmpr2h8N7DYHT5A7123nJ
PnbiJX1YGyMlMMHFs2UdpJ6l7nuVKNEUp0d9TRfo0lnOG9+zzxAKvNUejTQITf4X
l/Mh/nFAlqz2f91wI0DC8VbDXVLcxdCHK51bdY1hPnHeFUe2hBHyoY5b0aV5uAs6
T0sQXgrpaa7YH44XIYhKzQ59Z/H3WjoAKJ7SD2c8F01PQnJr70Ko5FbGA+1i0+Vy
ltEGjHoBqTFLhNnbHbhgmUrp6Qb2IXFEDaymVnbQCx2+7gHxUdzS4+JVpm4cCIYA
nDxhU7AgaZeJeyzjx3Vz9YqDv2h4DSQfuUB2+QOKSwpVzpYV8e/DqARvO5cl2JQP
Pij2F4bMP5YGpken3NfcXkPLFQ8fQDO+bSJlscQaiISuf07C4o7OqY6Z6h1bl6mC
/VnxFSpDPTleXx94aMY+EIybMEDn9BNgQq2XRVWdb0/X4ZTqYn+JUge+m/I+RVxV
mVeaK7ex0T2MU4eeyPb2pUxrvRatoPyYaBFitMDsHHnhhYjqfnCQCRgaTb09p6e9
B0KDyU8FgbjZi7kamRp6qL1GaQPP5ZVFikiw5t4xhjzNfk5LhisGlMY3OTav+eo/
424d0iw+ygioAqsYHKAfw/te83gNb5pFRqL8GW21BBNfdAnZH43UGY8FkTyO+iIC
Su8lsUCiumMhZtKhWh0UQO8HgQR0b0jRQEHjcaTHnkHeDBqTcz0SwL3LWDgYAAaF
xPJyF2IMBxKnMx7rMenH01gw85uEAMxHDzWQgSPJb5x6ibPoVoBpX9UjTsVsgOvz
hJaojc8wNieyaFSF3xA+L6eypfDy+tgHauTufIsgTPhNfBfOwa5UrxVDj/CTR+9p
qFiLaBsvmaYFyjc/XmW4QuCz86IakbGHHwQYGOak4xWaYs6p9Rf9HK2t58qu+0c6
bokP3lluiEpzC6/9MTJ1UZ8qCeu0Sh5BJCOJwW2S/glVRZLm+KCeWT5BlW+fLsbd
zaH23EbjqjTgnZ5u32UhmDwaj3X27ixQj7TVN+FJLmABw3uVA6vFQD5lOscO10PK
LqQybiXIQPx8yeUb5LdQhv6JZmB4OEqXwRJdzy1/U7Zh0+l/9ytW8vaglYLUvfgK
FCpS77S33vZZP+o6Y38+9QlArqV++YbFf+2MK+RmR9mUT+3r1q2OemcDxoiGHQ1P
fu4vgE49bfuZ2knOC+siSKT0bvuPHhM7eFWaUkC+Qd2DEQ98ppTWotEAgPeKNiaF
xZ2YqJGq3gkXjHV7HgIfUb0ngt9y+5VAgToQk9LAtd62unPkaO85wEYpU1gRqH+g
7gwpHR75s0jXWRdw0q0c/hKq43t41SRw2NAVJck1NzSzi5MtIWYRsWhkbBqtDLmY
IiQaViXCrXRj0jvCgBQ8g/v2hszLiYtgr6GW4kfofevyNTETmtBr1RQNWBu5u8RB
kIEHMAaAH/eh1c+jgThB7TReWnbiv6IUeNecMWS5ztIURUAWrr8zm/ebt/M9o12B
UuP2+CqTdSRCFPsIMrfwbQ5RBj2/ecvtjDJrMMWfG7/v7nW47kBFzmkNNrLl6QY4
Qs0JivGWONdxqTAt+RLqaQ==
`pragma protect end_protected
