��/  y��:�0�	]�F�#߰��eoC��{b��r*��q�)��}�␷E����]�,u(�[�/��.��#'fhz����m$�"QnȂ �gl���j
����ɿ/,E=lV�0ogQ������԰���E��u��|�ɿ���w&S���Ԋ����H����#{@��)	�<�:3eE<�᭮��yJ�Z��X^dݭ5W�!L�cSa�&,�q��zN8�[�cӭ!��K��,#�U�������k�#!�ܼ�jH�i!r��$�ۃ7�g�ۇ�P��J���F��dN�[y��Ov�4�eC"�Sd>S�}���/�;rȅ�d�a�e_�Qx�¹����xc�u��S�@�����w��n��M�֮a�G�����U+�e*���'V�!�}W�j�LRQ�=CpY����<��9UK�V�"��	RL� ���a6�]x�_iX�m��rʙ�'g.E3e�v[��fS�@�	$�%���U=l�\�|���-���h�YL7~)4����x�E��1���L�W�L�>F6�_݈�7�2!�Γ�j#dC���s)!U��tY$t�lE��?7�n(L$�3�iB��6��s���˶-7SOg�ș��,�Q5��Ɲ���#���w�����g8o7���8N�$K~SfdI�k2���dR�p�^=r��T� ���P�)�q�e/*=�^E9����Z(��V]�:[.��7��d �N�<�湵�_k4C�oBG��x ���34����|�����6p�8��ܩT��yW�=	�b� V#�����(�Bk�w6���?�\v!��q�� 0+��y�ØVi��s�}�r�yf�;�������+d�Fu����q�s{���I�O�4w�*�����a��n)B+LQlu�(K�J�
�e�o�ʬƯ�� ��2����v�G��n�fnW�� i�Pw���%�W�
�u��Z�-�m1�x]
��1�.te\�JW�e�i=��%RR���մv� o!�<�C��.��`b2��j�̦��)�@��ިY�	�y�.�C�֦2��EZ�g���Z��>aګ�(9�T �!jL�<���x��B�PKĝq���\��iNsr$PaW���;̀$������@���_�r^�|̀i������ыGk�Y��}/Sx��<��ė�av����w�*M&�����Q��q���߉�� O%ͪ:ri���ԏ���ډ�}Ȥ�>QvGn-��"H��_���x�A!}�}��&/q ��őZ�qH�]��x�	�઻���fC�C���K��I5�W��`�jl��{���:5z�`ZK%�g�=<�$��/��iG��\��};4-�4 _�
18��X
�;��u]�1���霮\�^�M;��|I� �Z��.	��2�� ��G�0���bc���]F�6�&ɑ� >%����k�dOgDn��E��yR���y�[O�N���Xk���P��[��ȩ_�w�Ti�N���89V�Մ������P�x��ی�2c�p��tzF��b�!I�-���|��K3��i`�>1���GYw�)q@�4�
_>n'�ӱ ����N�+�!e.��X��7E�����0�; �1����V5/J�R^� dj��@��L���i��ӄ�&M�׭�ZZ�o�ZVnu~\�äw�������0EY�pN��'ϭ�[2.�l>� ��C',\�M�zQc�*�6u�e�p�}>����3l����U{�'�a���@9����- ��
Z��U���E�M"t�ߔ���n�|��(�_F��M?ɑ�X�e�#�'SΩ��E�y�\Nh��j�*K��. /`��ᐤ���yſ����%-q�#�\�s~�V�	����{�_�fTj�-z��������8?�!J���bMu~�<�BY�����Yp��[��[�i���3"�y�_�V�bJ�e�e5q5�����"U#vO�i��3
��X^��L��'�'�� \��/�#O��6xs^9~<[.���� �W
9�[�R7�����汇5���\�|:��\�鸟�c���K'-���K�>��EnF4f@�L������u�w/����0�<��Xe�ع��Q�L�>���Yt"�?h��nZ�V;]�������7�_U�T�+y$2��T��o7��-/��wՉ�|;s��Yh7�劝!
h��EφZ
�ު��HR	�K�tKA �Y����*�.�é�G~&i�Q�4�_���ʕXc�S�oõYx�st�
?N��:��Å��`Uk�Z�K+��q�B�:*@6�L4�
��A:��'��.ӕ�J��ŏ3��6�f�7�Z����������V��7^c�pb-=�%RpϽ����m$*�X��ol|$ �'2:!�4�'�7kl��%#��jGџ�dK׸�ICF����{�����b)R��b���'��k��C�!���A��l� }#F}��8�7ҩ_�*���K�<֠�vn�)���ǣV$�.����Z~[�������k�O��������s��g7�+I�D^1x�T����
�h�b��+fD�nڜN.��?(�"��'C�e�b���!)U��_\4Ѧ�a��M���J�sE5IUhW��������鱋T'�_y���c�v�N���������k���X�����h�|T5�(3l*��B2�Ϩx�CPR�u�s�x�!��Ъ̦6�pc~�s�,a,ퟺ_ԍ��Ɇ�c�'v̯w���1�1I(%{�ɪ'�]څ���K�Xɐ�8�b�^i ���}����-IqB�4I��u����Μj�	���P}ʱ��ILk�{��j���]�1A�����
�~SBެ��G"��&Aьw�"9&��6� ������IZS6`oFȋm�?G:(�ģ/%�F���.��	7��[vA���w¤�@��@��R��X�c�M��g���F�����/e�4H�zf�
������
��d��o��>8�fԮ>OB��w�'@yP�)�b9f1��ޞ����;[�a0�	I7x�|��_:&ȑ'�đ��ɶ٥/���ba�0���f�p����(�8�vu�S����iܚ��/ʳ�����(���`z���A�ޣ�/�!����ĥ[�C�(�ݙ@B �hŚC����+���q0����N\U�Ǭ<"$�*I3�y ��d�۬4t��1;�X��ֆ��R�	÷��q6ԝ��d��*
�!��R�CN�g���:��;{�k9g�(��5.���;�
�����S��gj����z�����Ђ��bm���������>�ۓ���Y7�VC�!J�8�LC%>�7ˎJ�F��������&�� w�L0����%��N�G�n��oU�D�������v�M#�ɵb^��<(�9�"G����+�0N�Dyڃ5_�Q�+��K�]��,�%����¬�E�ki˳�~Q^2�>�ʹ�[����_҆�����NԾǠ��&�5s��ó3,T.�8HxÂ,��2��_�f�\��+&��	"�q���]i} E�SB�V@�*+�=�צk(Ӳx��ض���?�.�Rl�Kt�����E� T��T��ZJ��w���=���OO���C�f�]�|1S{>_A�`7�-���Y�]fOj�j�S��3��߿���᧏�]�~���+ɋ����ͫ�i�����E��D�_~8�pE��ک_��G�?
1|D|(i'���qF!����[�Ҩ_f�*?fڧM6��ubŌ\dc;��V�GF�՛{��-�J�2��Yp�����]*�ؒ3"�$�_�=k�5�*6��U(ݏ i�o��)�:J��vl�{���H;���CZ��]��.�[���D �2��Hiy)����C=9c"��U ݠ<�D�F�y��������|�9Ίcd���Y��ř��"�1@<����Z�j�?-���g�V�
Ea��?<�!���U)�*��}z�'kxk��%��W����o�(�M�߮o�v�s�����v3`�����d�1��]*Q�T�Y�1���s���z��PM�Wڡ���orH��RV�&�fE����)F����ʦ�5Q�( ��\t��'kJa�ϨJ.��:�����Н*�8s�B�~��.F��J��������K�tFŴ�Jg?N���۩uR�<�b�����X�Y%	��4=0ƒE;���I	s�nn�]�S��{j�ٜv��W��XHƅ�+Z1���l���w��+�o��zp$�{'`��|U���Z#	��߄ٚ?���E�\-�o1k��o���ij_�q�.!Jc4�Q�xgԟ�~_oͻ+C�싒B�
����]��(��O�/̦�BRR��Z�='��@Hw�$���
�
��GSl~�p)����ɝr��	Ʋ��a҇Tb>d\쟚��X�fnߡiU�H��Jl.v��L���?*���m�3F�C�y�p��f\�}7s�`�'�6vE�պ�W��$�Îy΍]�韣^�pf�}J���Hf>��H��3��,À)�>��x"Z2��Om�uI�i���O3Ȗ���IBd8��'S��hXH<�N��zU!lgs76�ʈ��Ċu~�����Dr ^�����߃ r_���/�%���!q3T�[�K ?UKi��%��=@���I��R����������>�t���(Rh3��.�@�q�N�?WP<iHӼ�p	�DL��d۸1�>��_ԿDl����ճ��L˿��}۪�i����%��w)X׃�	}�"ܮ+�Ea�2mj9�����b�~N�rzl�k%:Y�\B�;�k����7M�8�s��%W:@\��[HO�9�z�a��3�'�0�>�u���ć� ��-�-R
~N�6����^��G��:R�vO�1��;ˍ�oq����ʊQ�k|���> &:�*lC��֩'ȍ�sN:�ӡP*�b�GU�GF�ռ�E����&��j�X�a4���g�?3�$C��|�Ni$�A�{�H�6a]��.,&]��+0g�W�
����~	"��\�lo���9{�{�v#N�aoF��^Y:���+������S���B4���p���U���
_Z��NP�%:AF��=r��-��fٵh�!'@]�Qaj�zD�ʛL`˗��/O�4������k]֝|�������c�(����*�m������?Q3:Hg��㲝�ʚ�e����WI���}���>�w���b�����x-��۞L@�=A���ז�$�:�d��ҕ̺�d��J��:��F�I�ۍ�f����5��Pŉ*�} �eTn��ptz/;Ϊ���Q�މ֢��3���	�����m0��n���%��H�h�p�9��=u��r��H�����b�C�J��:��A���UݫY�h��=��5r��ߛN?�&�R�&�c���܉��h#/\A���S���]����|�7��mC��O�
��� _ҒO3py���xPk�솄�qW��~
�xN�XRҗ��������!��찚�l��+�>�x��[�$��1Q�0\@�j�+ �ù�f����W.�zQg(��V{奃{�9��f�\	�o�N1�t��v*w&*樾宄d�*��*���}	G��>"M3N��Zҗy���5��7�$�v]V$���7+V���m ^��T����;�͹�S�����B��z�!�L�@��^�Xq������1�c6�2� �t_�p���`1c�"��I�5��ǍL$i�Gb����b���*��KRJ�lق?�P�Lca<�s�.�jSB�fZݷkҴ�te��G]�c՟5FMSq_����X���f@�IwS�������#�l�5�cP �Qg8�;�n��ɗ����+H��B����lq����a��s���� E�����1�%��R෨ȏA�悙�s}�*�jU��B����/��[-�sE0�r?�!���,|���i���0�pԓ��4�3#�)�g�
^w��,0�����HY��fPC΍����T�@��{1����:PFXsݎgSG2�U��S����9����{fT=K\��ɠ\t�*ykҰ򺐸ۅ�CS �C5��?�q�_��\�-܎c�]W����Ѣ٠��u^׍�;�%��!Rf���#}5t�YX>�5��AY�N�s��۫P�o���#0�/��یF��W�m{>ovX%#=؍Cg|��\�h��@.���g�?��БV�C�E����\��h���f�v�Ψ�*�vmby�M-P&�[:MBx	)��g�E�d���ϐ���b��wK.��φ��Ī��?�z��Ʊa_g5��OS�����B���_���I�7^jwu�-�L�<�B!�����J�qX�%����Q�z�if���;J;{�-#�j�����ة�\=��Se��NQ��o"6}al��|��@G��-r��yd�߉��+��+l\�}�^��A]0{��h=`�s��q	r�ݡ����c'��T̃}܂�$���Lр�^;����Q2LJj�?��ٌ�
 ���9�e8�-� 2�� p��0X}�(v=�P��@k��ƣ�8f[���|��Q��K{��>X�����0`-�g��
��ƝTV�'[͒S(-RC 5e3ǕYz���FKշn����2�0��uCt�۸/fF����z��F�|�h��#�bN3�($��_��E^P�@��;=/%��{�E�J.��m-�p�sרTa�>%?���r��nq&���V�y�]<��Yu3����d��2�[���P�~�� @�0�n"kLD��| �A%:�EU��e��𝹽&JUdx����y��dL���a�/�ʣ_���-:�d�m!�{vG-��?LD����8Y���vh���Sd
%�x������� IR ��/�͡�Ʊ]��0���贶�5�cǿ����*~�{x�Gw����cv��}��z���Z�r�O�D�R�=�/�����<�!駚�*��ɣ�} �|S&}7�������K�N8�����M�mŢ��
�k��à��M�!�Rtٗ�{c�e�M�}[&=������rO��͚?w^Ի�B�O��*��ۊ�̊���M�N� 3�XȌ��V�bjt6�����bt��X��5�Y�u}���K'��[�&\�W>����fr�R���4,�>�X��k7�Rx,�@����a�+ͦ�:n�ЧɁ�OLf��e��k��	���<U$��h�iϮ���������f D�iāP�$��+E��B	<��O��2�	�ՠ����U-�5��}��W��وoK��W�/Hp���%j\��[���A�X�[����4C�s�wY}z��ȇ��g�1�u�HK��f���s�I��υ�w���I�b���⠎kk��ia�'�2���p����g�J�����h;%��L��/��g����ՔM�6��e25G�A� 6���8nL�Ή�/"�����A0�gY����1U8��<�N?L�v���~M�D~汆��:���d����g�k��.h 1yS}��+��/���� ؈���B(*�2���yz��BK���a����=O��&��g,�8��~dF[r? ����+�;��L�<!83o�Ɋ��:��2���� �������Ѵ��6�!�֡9R���#��)y��7-��,��o�o�+�p6���*TAjz�jV���B Pl��c"֗Tq+Xl�xrfL��me�y&�������w(�F�ޭ������	�k�>1�Y���]���pp�0�@��.�|�ڜ*���pAK+M�|$��̏ȭ�^��sZG�Va���v�!�!ɘV/�05������̗['���>oy83vБ�iS��L��h�_�9�]�$�`�nnDc��||5�R'LCgXlu�h��f!R�h������4#p���9��HE��9j6&%R∴�r�nVoBȓ-6nu��K�5�<�:΂k��d��S'��D������g���k|瘧m۔���8WU�3���b�%������xv�tb��[��(o �s�p�^逋�L��I�f�f]]$�|8�h ׮�$Q�L��Ѡ�&b'�֍<T�tw��J+;B��\I�;�3�1,��=�9̑x�=p�+"F�q���%Fƶ�H�^8��t1��œ�ϾV[�`��^���ܛw�ty���J(�[_�O�.0F�I�D
��itjR�w��.���̇���1!�Du�t2��~�#-����X�PW�Ȣ�OI��J=^����h�N�5�+B�c�3f`�iTy_���ď�<�N�W��,��*t�po����-�ai]#sz�����i-���ޤ�3r̀,_��e_bx<zq�K1Y7?��/a����Yɍ�ԱjW�/�w�f�eW)��l�pX�A�c�vA���5�m��|O�c@�Y��I����<�~0�5jh��_�*�ʸG��/�.(L{gJ�콇|IY�O�j�a�.�&y=x��Y�����C�� �!�2��b�OVbR�(<�hj��2c�_��M<��G��=���0d~K^�6�5ka/`a���5l�>�d�ң��Uf(�ư�J�0t�5?���|��۞�Ճ�B�&I��_��O[��*CR�̠$.%�4Y4-�g j�D�hG�S��L�Ks٤�Œ4����o�%%�Vb�"pc�1+�����q@�:JW���hD���;P	��L���X��]b��	�'��t�v����e�-�||B�'�J�A?r[���#�Ԫiu'���l���y\{c�$C`ò�;k�N���AĕNv�bb��3�W�E�B
��3�̣q���	вJ�'.1���$����� �O�}ϰ���"EL�\����J.�K
^HOX&��f]=X���WXN�j^Rv���$��yg-S?�����ȅR	r���Ր���Q#mJ��ǰ1v����� ���z� O��"(U#��؟���VM��&���yz��'�d���si� {_:����>�
�@�T*\m�ZYq 2ly����z8yf�7�{��4}1���(c�7*d:� =��A���a�eJ�����B�������y*b1'76~���Qt^�xVs���$�v��������3L�R�lRY��C��+j[t��	���s贷��߬�W"�SZ�E*�CE�^�[�`/مϓ�s5W�\T�{�!#=��*D�<��DWW3-y�h�Էu���#h4�3UJN����f{7@�<ShsY�6ϊ�Q6�|���Ć�dm�A��}zDd��MڡTt�n�y)�O�i2�Pͫ(�j�K��	"F���-�<�Ef������w� C+�4I�(��f���7�3��mbh�W��;4>�e��ۼ�2zP��"��%�X@1
A�fl�G���T����0�	�I�Ө�W�ꤳ�*�����
t�������wMΦMQӭ�>-�O|��1�O�z��l:�aV���r,�=fƵ��#��a�������4�!I4!��*%�-����"���v4��_2�&~���t���d�tj�i���0[ �Fʠ�� �s?�f�w�v!��z��Ͱ�)u�KCJ��f��2~��줞��ʛ�?� R+�V�A���ݬ����[���R��+6b�s����r�J�7���Q=��	��,mX>�Ǻ=�ϿIi�o���ݽ�rC��K����<dY'���e���#݋F^HV������l�*85�cw��q��ƥ�S���P^=�c�ݧ�O�&'"��h]�$ Ҩ�2e�HZ�r�n�{8�@f�7�b�p�&��o����7i� �ŋ�?*��f�^!�V�7���g�{��<ҕ��	�%���Z���}ծM_?b8U�:\T�v�V�g��լ+96*d�&!��l���!Q�th�[��f��Qק}ڹ��P������Ӽ5&�(��f�O���a��:�]������yL����@Z>
d�n��X����be�R:���A^��(~i��ږb�7 j��q/-RA�����.��_!:� ��p�����ܢH�{y0�~�Ҹ�6E�I��خK�Ǫ5����MY-�\a_��;�3����YO�'.��9�=��D��lQB��P��v ��s�	�J(b�2n*Z���� ��z�f��ʰ�f�����T���h�������x�	�mZ;�zU6:HH�q���F���$[���E's��� �1�]�aT���zk��r5�������'������u]S��QH�ʴ��n�w�� ݢ�d*����%�8��"V	�m��Sv;�&⺮��Pu��F�_VF:Q�<�ȵXy�"��(����:�yaǱ���!$&��g��K���}�X0�
Q3�9<z�dMn{�R�wo�J�LVltɭg߇0r����	K[��ig5:���C�����q?�U�,�d2����ԶĀ�na��h��e��-�����fT�m�;��X�6~����*>R<�=�?�v�Zȸ�͡�4��P���i��^µ�<[����]��!����n�T9�X�qvJ1���v(#[N���nS�&C���cq1��������5��f���~jv��܏�t][]�Ԃ��(W�HHߟ�zM��e�u葉�DCt<���'�(�)wOǘP5Fe��j��1\_O��-�d|Z,��R�q|�ݬ�2��^DۄҸ��EX�����eMQ��"UL��C���.��}B6��-��S9?�66dcaU���HD�� �T !���L��Y\���3�wλ@��Z�-=�z�o�4���H���t)1�ϖ+�^�=�_š��ز20������V�_Q�t`ǵ�-� ��E��=(`4 �B�m���᳛0�#0�hd�-�Hi/���f(�8�r$�zr�������o��x�K�����*,W	�z��;� V<�#�%�������!�X�� �=L}V�����rz�0�Uv7ËLJ��cŉ�Y��Ւ�k�(��Om��Fn�i@��%V�����IC��P�wQ��̯-e^Ȅ���o߻]�c}lTQ���j� ��Z���I}VSN\_!�#g;���w�C�3�ĵ����w�Ȧ���'�l�9��A�)�yT׌rԤg2H���}�vB�-6�̭�y�y�`��r����y�˪�'L�6�������8($�p����"]@[��>���,6��l�o{��5���pIW�t�bԊ�5�!.���=�V"F���$+�r�!��5jݛϩ�m?ޞ�+�/^��dIҊ�p<l��L��b�E���8���Jǳ�Y�<�׼>��lB2��r��S�����*�S|�0ej-�*v��K�g=�i}!NJ��/��|�-�Ǩ	lQ=��u�X8Z)��͵_#�ф�t~��rn����$ a��J��iF�P<g-�y�`�&]�2�L�벳(ꃢ־���5�����~6��Y"G9%w�O��Ihai�U�/�O�T\*e�'x���	��x����Ȣ:��Gi{T��?�Xv�X)=ã�0���ʹu�m���&���E��/m*��c�Ѳ&|�׀�Ҏ�Q	W9��-�Z��k���lD�������*?^9���09|�T���{ ��$��.8�W�x��{��C��5���喍 �d���k�?C��ٲ�!�����s���+��(��Oӝd�;��@"������'<gC�����(� g��g��Fz��ŝ�\ڨ���z�^��W�;a@���D:��j�0�ʖ�O>�z7"&J2u;�|. ���br�$��0�OgyݭCאkdn�lAZAJɥ̽��u��6�ӠS�t3{�x5E�_X*���c�_���8�A�zi�9����M��ff�T��치��Q����{a�FMuPU��4(#.Hk���
Vd�4����
IG&����F�>����x��ph�բ�hi2-��tN�Et�X�p�m�9����!	���I�'T��o��ň���9�?�=�T#�+䎎1��"���0��&7P���Ml����=9�����0j�盐t`V|
��$N��l^��%N�O䨋R���$��%��~Fi�N|ٸ��s�h�}���L�f�+�I�]k���@�$��C�d�dMW<J�
���l��G�i�B���'=H� �N����8-���AmO�v�?w�ާ�7?��˺��H<%3?:��_�]b����G�����2�pD�� ȁ)l�ϔ�b�?Y�U�����Nχ�@ﺒ��0�����%�R4�T&��h:V�>s���
@��|`שU�,�Zf�Ѿ�$ЖHgJ�N#~e�V����+��t��+�TK�r��H�"���w��C����>�[mMB^!9Eֽ��8���^�Ʀ'~3��噶5�\<���Œ�Rk��±�sy����D�F􀖴����Q�YOx<�+�A$���H͇N��p���-ǈ�*z�Op�Oj�� ����|��'O��yx����j�T���̎q��~���Z��6�<3%��p�����J��_:�~���ͣ7��_��S���⸠�;��q<���S�!z��O'y^4�e�Uj�H��%���-a�G�6�=:?$�L�`��G��Yv� ���A�ZSٚ��h���4���ژBbG�ѷe��|k4(�|D��r���x��4R���ۍԬ��<�{�Y,+���O�f����5
v:��e�N�9����"~����[&&��t�လ���vQ����g���QL,O X��Z.�#�1[i*��X��<�c�� H��s�6�Jhwc���+kkes=�g�2�tHE��F����u~˯I-ݞ+��!�W؎g���GO���ށ*�%@8Ǘ؋�d��Ej��W2�Ж�.)1�@]G���\m@���K~�e;I�R&���^`�����
�j�c���Ǻ.g����v,S|�W��k�^%|�`5�@�U�9��E�#�q�+%Mo�ت�S)�y����ޝ�ta����Ld���>�h�h�77��gt�l�2dт�D��I�������F���������Dz�c6�f��]�~��GiY��kaiYF'���C	�C&7%a�_"q�Ê��zu��m��4�K��vN�4��E a�3�^͑/z�&P�ca���ēȝ��=�k��_$k�Ͳ��73EV��[c-���-�#�J�4��I��9~?��&:@cr�/����[ R�m�x÷X�n�ZĄ8���/q�?�"��H���x�
k+�Q#���\�� ��a#���i|(t�M�?0��տ%]>��a���]s���`��)�T�������ka��O���rߣ#^�uF��_w|IG��(���.(��8�Mf՝��o�2f��{�^x�.O�6�&0H��e#��~k\)GE�C�j\��7m��wbE���Mv镖^�nV�ÅJ��3kF��v_�3x�A�@��jpP�}c<����@·��x�t�ͩ���9OK-���������[O����^ВNd9D#�r`�l�s.-��|i�����l}�����.���6�����R>��"��&7*vX�x�N�\O�{++������"�_U��$z�����@�u8�aqy5��IO�W0����b
����n�Y�Z�CXꗖ�
�]g.L[T�Y�(�|z��Y�7��f0b�(��(�;�6���W�{��&ڨ�����h���"/���J�C�\�y+ȴ>���_�Z<�N�\�v�?��K
R��8��bcš�q�AǄE@8���l�}�\�=��1�����N����R��aٴ�ȹ�yJXq�{�C���x�Zge��{�`ʷ�"S=HMrY��v<x'C��`�!"�$�]_�_hݫ��Y����q�3���1���p���J��YW����u���j�$�Q�N�h4��� 7�^٢,�.���t�ge�q�п�A�mS߃����1�V0U��%vo���:3��MP���^�M���l�D������?5�1<QxF��z����A@���,���\i2H e�ۺ�h5�g�ȇ�R%��D� �wt�.jfo m���1��5��Ǭ��"҆�1afm�^q��1�:m/1��Ԫz��˥)�V�JI1ݻ����}R/�X2R�hEcg.e� �7��/53rP.->C-��5O�5�]�et�V+9��b~�
�`���Cs=�[C�FW?ѽc��r�|@��C�to=�Y�{m+eB8PRa���H.����#u!�c���x,�����R�]vǃ�8y��N��\�u��c�b}����G?���:�V��u#�1_2+)����$��v���sO�Q
�`W�
�Ģc[,LR�xuU�g�ҩ5��T/si����\jvnQ��%���� �,�H!��������u&�['�� u4��/��#o����L�G&���0S�~3�l�6#��}��^U���3q[!(ޏ���P����9��k��$��TG3E��y���01����);�=աN�$5Вh�IY�H����]�>֬�)ϣ��Gy�������\��h��ῑ_ӭY$�����ja)���T&oI��=W�?=���h��,D�dl�"��F��K�	��Ӂ[b�=��p�:XY���o�*ng�Wnl�&"�3#j�>pEVh{E��C����8��Ӎ�0'1��}�u�&�M֩C"��?�Z�+�n���[��%��	����箄���,M�E��d�dnJ�?��5I�n���J��
=A�>?��dE��y����'�;P���k�[k�&�-p�`q=��̾�|;��G[Z?��}��w�մJ=lf��$tЊ!����Pټ�ź+�d�V����'��-��	�K%�k�b���Y��d��]r��|�M.4��-=C����Q�RyU�R��I�A ����S�n��]��cGD�@����6����^��w??��Ʈ���M�3����7��FJ��:�a��w��E�8�J����=92�G%��r��S�,�>�yԴFy �C���ب"��r׳L��o {5F-~�����8����$�k?|<�w��8^>Q���-L5�R�M�e�̵�<k8��k��ҽ4h��a�g/�!ܵ�9}l��K㷳G!����Ӓ�a��[i$Y��JZ�����m�ΣTNf��H�5�;���k8};L�ة�iFqG.
s��/�'l����C�����6"�C
s�ב�2�������`c������RK��,3YEDN/�Z� ���=�Ȓ?�{�&��M;�:�A�%��NϏ�_��-���RB��~v^�P[������z�Ǩ���w���G:.ހ��@��~�������ͿYj����{��������.��n���ʾ��G6"+��p�2};����!���·R��3���f�2[��0��F4$X�z С�����Dg����=��.�L�Uʶ)���X��r�ْ��~�:bN�; ��zٞ�)JO�=�ƫ�a�X����,מ������m䖉xou�c%>����Õiݒib������X���~��i�M�]Xq�f� LE�vg�.�bw�?�V
L�t�����Pk~�q�zjE!Ot��3tQ��������( tF��u�72�{\)�>(5i��U��t5�@q�Wi|k��m�:�|�a}�׶Cv�����<�,���r�QB���!�&#� ��&h
�5Txq������2k�&Q/�W��4®D�VG�����č�'�@���3�CF���ul8Gi�;���i�,H���/�ǘ���U��u�5�>��+!Z���Uډ4��fyg�W�v�>%��b?�ҕ�(�J�^&��+ي�r7b�/-���a�h����	�b���#���;s�Ѥt�#+O+�DTD�^�&����%z�mS�*���Z�A=�Q�cn�W�izs@F�.f&���b@Մ���D��-��1Ep ��Ȏ�Oa1W���U�ʐ'��s!���yB QM�"����M��+�a�Qp \���F�	��_B�L~ox奆:u���m�qt�9�#m��,��x+��Y蠔L�������\ឰ���J����.Zģ]�������~z�sJ񇞲�Ź�U�:����=����cOD
��I4]7����I�ޗ�f��*��?Y��e���o�Syl���b��(>���ϊ��Ex# ��Uw�"��y�H0�k����q^EZv��ٽ�W`\��}ͼ��
��49�|��kjw���LbtU�
9+����*�4�
����,E��hl���y3�|4�S
m�Vj���=��?zA݈_7>�ҍ���{ha���Exg�s�*��N�l!#�(���ٺڳ78C�ia��n�]��� B0ҷ�1Z�@	����	��Ҡ�qݘ�o�Z	�g~8(�=0��q�O?�WuD����?�x��r�3��f�0OQ�^�c��L�����O哴�7��?&�	c��TA�b�GBF����w�W͋kI��y�HD9pO�rv�wG��.+��7.����z�����{��ň��SH�"�o}�#`Ja��J!����׻V��41��dg���*�"<�O�"�|m�1�G�$�{Eߑӡ�[�ޅ"��*�CY+�' ��k�Q���k�%����;�e�6�d���N�Ι�s���,9�=6R(%m;.�R��􃅖�i�U)�T^������}�$"=�U����0���ǟQ��+���5#�t�<^�#]ǔ�Ѷ���Cs�����U����f��Z����kj��,��6��<�]�4�<�d��-�G�g�50нp9)�TE0i�J�)�W���(��Df���\��]���^�c���R	1Tb%��+�L��AH=�M���O��V|��X���t��ˠ�!����,���ĺ?P��� m���jN}�=_��pw�;G��8Ձ�n���Py�ub�����KHZj0�|+�iPY�
�k ���6����Ќ���]�}�~O@Gخ+:KTL+f����B���m�=�ˈo#x�W��ۻ������N�����Y Qp�t�(y��ָ}���Z�=�o:����
TI�ht����=e�է����*]���U��^u��Y�27@��S;|`�\���J��J@eѢ�ʠ�E��������2��鴑�}t�ˑP��6z�+�-��*?kZ�2�&K�y����<ͼ���֟�tH���20�΃2�Co\lw��&&�=����U jrWE}���:l�c�����������>�e������͛B��tD��"U	��WƬ�i������\1���'y<붿�\���6�C�@�7���Z��E	��y]k��{YH�-�mz��c�W�G�3��S0�=%O�?p��"��60خ�Yq$0���Kt ˽���l�7�p �'���J,�䐬���k���.�Ή!Y�l�^�Aw�C�!e�'-�_5hlz��m���toȱ�m�邿�K�e���j�f��i �A쯯�'o�S����Z�8��rR��}:Nf�Ҵ6�|T��ٖ]p��;I�� �����|9��vhcrN��j�F'9mY�c
(�q�eųh�'�@�l������c�t)�?�!2�=o���Cɋ�kfK�c����a^苀����O����Uh���bdx���/e��2�/�=X�Ca;��U��g~���
��VK<��V�,���pP��UѸG�&�����"H���J�S �űs�%H���N)W즳������6{~2%j�W�Mڊ����(;q|�^��,ў4Ho-�P���#T��=p'E�4�u��m��k�TWM�[�$Ö�Z1�#G:R�!��G��\���GJT�\h�a��x�PD��g��(�{{AԦ�z��|��g�j�j|[�NDn\��P3�D��*7S�y�}o�����1ȝKK��8��h���n�����.��M�\^�UK9S�!}��^��D�y7'�#(7��T�.(Gm/��{^ԯ���Y��[]R��P#�e]���|�V¯���#a#���������
�r�o�Z�T8����FmRn�s>��<��UX���6=]��a��^�AV�Y�b���^𽟃z��-`���`(0W�5_rR8膉&Ѣ^�H ���S?�A}�`Ye߷}?i�QD�V�k,q����\�nR q���s\ީ��v�n���	ύ�$�]��G�C��%�B�1�M�WF�Z��Yϭ�=A�_,�*
���1:���/������^���)�o�_�l(���0N������4��!H��F�ET!f���;���C���ξ��u�P�~�>FMȖ���hp�i���L���B`be�^)-�K��Z��dm��T|�����{�}����N���JGp���5+����p�Q���1u�/cj� ����V�26o(ְ:@����҅��i����8o�8��8gY��+�?���%�n�"G�<2E$�z
D�O��q^��y;�yӨpC�������
n�/�[�v�r�'?�������W�y�k�Y�����C�+�+�	%�֤� ���k��V3vy�ܲ���+:�� Q/!��~is>+����z��HB����o��a��<y�h~H0���ʓ�]�z^��P�Yr���ʁ����0�r-Ha!�G1������T��
:�:�'ȡ�{uW��>�����3�<I�(��{�����t�ɟ6o�e�U ^�Ҡ,���tOL���� �mk*�R;����]��Z���u�ϕ� ���;S���Hx����bՋi�D���7�a�ް]�e��OS]U�7~J���Ƨ�b9W�h��-��'IMa���p��Dm�����ƘЊj��Q,�����G����T����*�Au�,�wB���o���hx��d�hB���T�7��[���@�\e,���1��OM�#���5�gE���=By,|fX�^�'�V���~�Df�Tj�y�Q�crl%��A��k)�h�_�����IF4��󿵎�&}�O��cۺ�)DN�\�I͂����6����E�!����z5�d�Bq��br�ۀ~��3��3��GX�?7�d���89��!^��!	2�k�K�#� _wJ����G��M$����_���6���q�D��A�o�K(G5���V=(�P�(jȉi�9��jƅ
��C�`�P֐�����'u7��t�|ݧe�/���W�a�&�����#�]8��?����Op�;G�Q�fs1�u2�*�ͭ1�����R�G>���W���뀯J��n�-E~��3�� a�%#�������6cu���9�@�]Ӿa�Z�"�@��..�+b��B&�ވ���@�7t?y_��ˮ'J;�Ĝ�xG��t�����_$Ui��@��i��Wښ�Y�E�r�%٬~w0��)|g�/Aѥck��<{lG��zt�_�9�!���i����I錌��M�;;�^�C��Ư���N� ��L1�A=RM���Fw�gS��Y3,(p-倶4B���Ie���J�[�ǜ�`[3��i���R#�巏�GԐpX�D+[kdH�d�{y'g�V#5?��ڹ����"�Ru6L�
*	�Ck��w�� o�ϵ�db�5�g@�O�I�8���̥s28n��%}�S���WmO��*���`�/��6u4�0D�K3��_��z�ŝ���Qr����O��a�r��������؏0���=��T�FvU�����r8-�:[����l���>��Hz�lZ�1I��b�bn�4�G@&����.w5�/��i>._W8��O��+���>�df��r��X���L��ޙ]���f!���H��[MO�(��e��s�^K�e��Ս쫌6-���@G�eD����@�#A��"�u�n=L���*ŋJ	sP�m8O�u�p.��(S=W��V��v����3ūg�՜�!��J��K���ԣ������#���y®��|��'ibJ����WP��Fe�H8PP`e�zT�҄�����f'�����~[pa���Gp�gs���Ҝ�n^��Q�-֟����t�j2Q���?'$Ã ���.�>��<�K��ť|nd�	D���s�w
���k$� W�f����hʠp4��l�)>v�����<wd���IF�� .���������P��GS9z���]~���q��a|l<������4�+aO1#1#�r�h���.n�q`AIc�8��yR:��|�ńb#�*����L<��^X����m��I;�����n"r����8��r��N)g�J�>��	�m�X!']�Nge�G�*��-��u�u��Okq��2-��膻_k?|ݷ�%l,<4\Q���o�榘���J���U�^oDQ���9[�����Oۗ��^E*\�\/O|)�_�X�m9�W��e�gJ\�}@�J
il~�H�kK�m�w!���������:�Ǎc���B��輮��|m3Ḛ�����>���X��nY�m������jjɺ��i��Ru�{�n%�߲������Ԅ�n� �0R����.�ɶ�~�Z�s��e�)Ź#��i�&!S�|�s����g�4U���g�+�bԊ�u��r(ǥ�z��o�-^���>���RB���Oh�~t�ϣ����,{��馽8���4i���L��t���9��ofϥ� /P��z\����fKp�ġ���`+V�-�=	=��.[�,:��9I�M^SRǹ��R��%j^c%3|k&o���0u
*t�Ք�+�2a�㰦����Q(��f�9ԝ��B����*�	�ͭ��$��wc	��n:DBYX<�h	��'��<�U����C����Ԭ4� l&;�Š��8*�|����J����Ǳ��a�)�X�[P2��+�� ���@򵽛|�#�0<qO���O���_ɾD��#���E��*�h�3��>��{�:��qB\�|m��+�Ӏ�\ULD��۝����*�4��.�<���&V�q�2�)�I��XW}��̱���p�t~��0ݪĎ���:����͎ꉜ�f-!k��h���:������G������=�}�n����H�B���;Z!��`�.����x/�������y�H�W�~+���fp��2��zN��Axr<�\����nh�;9��Z��'ۙ$�
�%����4
b�������-Ӟ�pMG���ڎ\H����r�M�!��i/��=6�kg�
5��{A:Y�:�~�k��]�Q�Yd�F�E�pc[cX����E�8Z��wp��OJ8�=���'�-F����SD.��ܩ��%ȣ���^-Cl��t�<5Wfr��Wrt�r��G��4VYo�p����5_�E��/��L0���R}�	%��ך��|^H��o:ՅşݠT��F"�T��!`���ڗ�*V-��:� c{|�3��Vɼ�H4��\�����u��Bly~g+�Qo��Nh>!�;�Ϙۜp}#j���0�5��(]� �ʜ�Ƶ#��}�(	�(W�m��W�T�n�#I��̂�z��?��ӷ.殑{n~O�g�#��k9�y n>�n镘������8���ISהrbX�3V���KP��E���Q�Ym�$ݳ�~�F�Մ�'���LB[�UB(����G{՟�f H��W��2n��rqW��P�U����m���ǟ;�����G�:���wPf��oa�yN'����{�@]Z5�er�}p��G{DCy�N���@Li�`��he�$��E�IB��=YQ�.ג���\r��g��鰞���eF:B����lJ���뇩�:��qL���~���1�ٵS�<X�),����>v��ٶ͖���{��߷��SZʘ'ʎ���V5&(�����+�Nk��MCJ7���9����Cp4ؔ[��*xUIny�9rh�#%����ê���E_ >�éUǌ`;��\�@�Ϭ��랪�e��Z�c3��'����W �����Z�h%��߆W��jW|�:w����r��������A|~m�a����[d�����Q��f+�1�=M��S��j�{�Ƶs�ګ�(RU���2��e����)(��#�(lQ�h�+�#1�{Ey-1�b���f��,~Ø����%� db�9�@ìXp���@ӷ�B�Y���
Qc���B�X۔fCٯ	�/�!K���q-�%�ѓ��Z�R|!��l.�ܹ���0�0�ׇk�����?�#B��܏�B�(�
��P��~ֽ6�,�h�!j�*��ѢU�I�9L:���vaq��@����a�b�z��� ׻��N�K�L�_(���a�f'��)�W䎎<]pC�e	�#���惿a��"QɊ��*Dqt��W}�7��^�8�$#�{�X�R)��꛿�ǅ�2i�&zv2����i�-
�}�ӊ�+:9i�����9��#��D�u���$�k)�8>'����<����V�[�e���J�y��R8R3%B�O���Ygn�-+hKcoB��J��=�$���M���G/�����5�����%n�j?Ш�����/��@��T#\߆��T���fo�d4s�zF�_)�M6���$���g#�{ߊ���B숚R�sQ�ć'����j�/�}���y�lΰ��s�����d�`t���!�BI�c\��@�����7����!�2�s��L�]��6p"�u�wo�_DƤ��q D�*�I�*��sa�}�n��e�"�5��+$�� ���MJ���(�Mz�����0-[���̒�E(Օ�cur�&|��-b2ur�H����2�?2� �4�A����p�Ю�r��Z�Ĺ��l�����o+<i'l�ɛ0�[~:,�^UᙵEJn4CX��ެQc��Qg�z�5 zТ���v���vq)�pP�/ao,i�ʟ�]���X�ȿ�|�qZ��9T�N�*{��^�����y���LM���Z�Qq�4�_�(Ħ�� M���H���OzR �.E���^J1��^F�׫� �5$$��������Jd���̊9��<���G��� �}Vߺ��L�/q�U�@+�j�����[�۱�5ͩD�FϽ�������(K?W�@UaJd��ۙ?��U�o�n�h7���)漮P�|4��e||5C妹�w��N�\���P���c%@����[^y���B�A�6��+��;�`�r�4�`�@;���ߪ�]����	� Wy{�hbF�]Oj�}��JZ�h�s��A��*�J�1�0��28*���W�"wkus;"�SgVD�k��H]�hH+\�[�c�wMjo똋�Q���Z�?�t�pyYzg�%��9�>s�|{��i<�R�u� ����j�K��Sՠ>F}\OVN�@��[*K\��2��zd��#�4��ݮS$���x�)1D��f�z����i��Y��i_=�]�6��\!�*8��m��f��c�D�>ȤP�_��Y�.3oKw7��5�S?��F�J��T8�������H�5�u�5>�g"����
�GO��J~㙸V��<`��ϊj�^r��(��'����lYA���hmxZ��ĭb`����*���i�"�uX>�h[$$��=94������i����ԣWE!J]����x0O�n��V�/�ʃ����w���}[f�|���ݠG�{8�e.h��)et��w�y��,��\��g�iSA�	:�a��t&���9L(�W�8ly&��,R�n9�,�" �E]�ǈ=�t���_K	�jë����+��T���}q~Q ާH���n~*5��A�����ރU�#���JJn�"��!�3'��x	��i���) u}R�\a��U1�=��Y�|G�rA�a��i8�J,�#�D%�!�����&[d��?U�V����]�~_>t�l�^�Wq���Sy�	�9��2R1�/��J��`��'E8�KE7f"d,�W����w�.(A��y��O��[c*�ċ����і~�%��AK���t�ɤSs�I.��v�(d���� ˜M�i1�+	o\[�Fb4��`H��]o�#D��6k�C�\��ɑ�A(C��m�Fcnx��+b��_�`����kj����PE}�w�x�����~ܴ����������j&�"ak7�m���59���o�V�������
rʲ�`�����k�}����q*����H�(�Q鶐�[��DH���ҫ�2n�&��[J�+�p��}#�0>�i�����m��n��z�Z� �_V$�W՚JJ��O�ew��ʞ��g>��'=���5L�ԝSs�+���Ї�C��|�T&���|`�X�Џ����T���}�rw���`�sc��Nml���YԿ��ƘFWm�b_E�f
�֓� K�(�N�J�
�}��E�*��t�3�:=��~��O�+t�Rt.���*�~�*����
cZ@����=������K����j4�9��qx�ý�k��Ŏ��`Y�K}��3�k�Gm��"^&�6IU��}d�A3؀�
=*|w�$ӊ����2�%7m��d^��w�*`��9 =���/�r��0���o{/�2�J���_DW�ǽJn�C�����{��<_<�_�S�.�{�}-CZ��6���}[X�l�kŋN�R� (:+������p��4!	Q�"�9��;�ܩ@�Vy�����\;���	J̩9.��
���s((Y�ju.˯���	����;4K�H!����Eh�h��b����\�cEН<ܢ[RT�q��,?~��G.���D������3Õ�SH���,?5��8���TKV�9�/1M<��y-��f�Z��Qsw��Z��.Z������'K*OvPB��C���C� �s��S� #|�v�x�̆Z���#��X,Tf��(�L��m�j�6����9B{�}����v�HM�f��vx�%k�~��W�k; ^e����8���ũ�3���Cb&��[��"�)-$�^$�vU�Q��ݷ�`�9W�:�T������*���v�detN��C���A*)4�T���] �3�t9�מO��s�|8����
wZ�����ʓ�W+U�$���H��n�ˊ�$@�\�Hh"A��me��
F�����X&K~R�g�s��:Y�/��_�|������#k,&w��gr"��v:��e�0>4�}س�+K֌�u[�䨾=��v�z�8"c"s�:�G
�aZ�:?ȃY&׀ᖫQ>�}���'ؗ�:�Q�p��R!��#)+��@�#�t�Z#���[2ӥ:��}Р���w־2b�R�o hm�f:�>��$���Q��C�JįA��������O�l��DRSmQsȆcrf4gm��}˩X-Hr�S&?����Nl��[[�"�Y��Ѽ/ ^ԉ��w�O����-\�_��sС�W��|[]���>�^���i���F� �I�(�&��)Dl�Q� ~���}n����3�s���`%�z���&�ŗoCm�O���PU����s�4�R#��ʓZ��� �d�<�C��7��v�G�Ğ�A+?����p8"��Q�tk�^������vBa kv.+	�}4#p.Ρ�,��x�ڞ�dez��(��N��/��W������є�m�+���pL,?�=�8�I��n�������O��(>�ޛ(�_���,���6�l��?�9���JF\f9�
Z�\̖ �����*�9g"h)��R�P��LB����ٶ-��qN�}���<��[衰+�(�G���.��g5��d���lt~s�׷��^:�[�K�v��0a�g��G�3IU��﹯,�b��π��A ���̣g�>p:�$GTg�9����G������bL���\]زv93�=��5�Q�E�t�7�V���K�������N�����[��
R,	$=y;���P�vd_�� ر�$_߭e����@D��f�94wr`M���f�b5(���]2��X�����&�D�"�sn�'�d��r����/�N��B9����(uށ*;t�9x�8��v���^כ���5.�51oB�r�, �n�'���	d=�|��z㳸��&�U����Rl��{�_U�:��� �WrD�Ѭ���nŻ��"��1�P_YS��p�dUP�QE�>ĝ����Հ�Qb���(M:ؓ�Ӕ�Q~�)�����(v��gcoY,L����E�;�'ޝt�BB���Bƾ �x_���S;ߛ������+]���%��35$��`��+|%�Թ8ԕ1��6$܏�+�Cz /��<��jS�� �Pu�0-�d|u�qJ�o����c�N���D�M�����:L�B�x	��5�l=O���)GЎ����|護�e��^/�b�	�tL�cI9���?:�K�[�o�cӂN��l�rkj=�0�UY_�^��}��:�$_{�Y����P�>F{�.����A�&���c�����I^�W����T<cX���c�9O���^��,A�����ڟ�Ν	�guxK��h�5����u{t����V�1��ֈ�]�׍li����J�$*�upt%";_�l����KU=��ǃ�F���IR�< ��n�oj��ߍ:]L�y�	?��=�
�*ıWRL�g*�Q^��jv$�?�
x�����N{I�^K̉x{�$;��,�����$���S������*����b*,��9[գ��o�>Z�@�(�Ϛ��U�c����po]j߿c!rn�o��8��7����֙����ƣ�I��p4t �%U��Ģ���Oޮ�A�۵d��������Z �Υ���Ph�f��m�Q��X�\��k��A�6� ����R��$5�g����S���k�'_@�&@�̤%v�8W�1��QY�d�1+�P�-�o��,Pp��c#Ts9��'t��"v��s���#�bؚw��1*E����0�#}{�bߙqh�^�u1uե%:<��f'��jak���*����9�z�<Qo3�ev��!St��}�]f�.��rbk�~���jW�Y}�=�tw;�x�!�z�%K�]���w^~�L`�Y8�^�V��
�GL=���L=,_,���\�V�6;I�Ǣ]���U*�fXG��$o�sL59�����5樕�?Vc萸�~i�BÌ"	 ��.>�@x�J�X2�aƖ4B�^ ���
5�D3,��#"��py��,��v�@J�<47N�R�vs�_j�qo���@ì`$�lx�l�l���+ ���V���n�k�q+L}u�XrI��W]*�L	P�[	�Q��L����z����&g��>��|�HC<aJpΝH1����5$
�_�g`'X�۠�yW����\�|�g+�z�#4��ߋ�y��R?檏�R�9�*��D+��]T	ն�̬����8^j0w9��ݕw;i��;�؞���l����k��T��6q�/t�+5-�P��=�]�x�ȐR�c'�*�#_�0t�(M�mm��]�/��$���^.��1��M�����Qpc�ѱ.(��Bd��\a��޹�ݍ���R�y<�2zIi��ü׿�j��	9K��	�����.]�Qh��nK�j���V�	ؤ�#gۍq��ɍ�	6υQ��$E�ֺR{��ZD�n��:�=ך���-ř���W2\[t;�}g#k%h�2V���S��\�E+ ��FԮ�2�����"���itUT���:A�{�k��ja���t�a���f7��IJ��?rm�4Y[ߠ��4c��ǘdQ�ZK�RYx��t�H���7b�
��=���(Z&��'����ߎvt�@�J	ص�x�n	ȰwG��33�l<I��S���?z㮐�j��_�,8����L�^F���G{����$2���[�e���]����pӄ�Yb e�Q;_MCu"~<[��?SjW�>�Cdrp1���|�,GsI0q�����Cw��Y�BT�����'��G�SfcS:�W�̸�૬���|r�Ci��W�]�s��bIb?�&.��?�Wc.�"��ޒ~�j���kɢ�''Ҷ�a'���/3�c��eR�TG�7�,�����rB�l�w�ݷ`�1[)���{��~(��0(�n �"�� ��ō?�=�����,q��u�v�4�	!É�x}8z=T�"U�.�W���ݫ��/��:F���@�5�D CJA���
P�zZOW�vz@�J���O��YD����a��MrEP��}�i<��y&��Q���&�_'?��#�^Ѫ��8@�IA �5��J�|P�L��%���]�`�_����I�%���}YX�qD�o���&��A���n ����g/��+�{���6�Ʈ�m�/ ������^�~��W|��R�%icG�k�N ��U�}{6(�M���޻���.�u���:|'PC�R����I35(�E��s�Bn݇m��#�+�H�����a�R���O=��ްN�r#[��\?M��|b��Y�㼩��QO�d_~e�5ɬ rƁ�tE<�bm*� �p��f��u2j�}��