// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o8fy/nHdHIq1avEYA0x2w95UGGVev8iW9RQyuVfRH5JOoGLGvQMjRAP3MOnSL83v
KAa+ytQtY0jpOZFbsCRZYiszSK/YUdb1N15Uj9D96zv+yJLieG9e6/63w4kfMbBQ
k0ZHXwGsX8EAQxwSrVyHOgA72cjUS5HYjb1HKe2JJ8A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6336)
fOUKgPoYkXuWOpCPabxBLy8EBi0cNNXu7tyaNKYwXWgzm9BpCUciUvrKShe59LYZ
JjVltNsQiNRiijpbO44VMkgWW84HKwgGlXmS836Vn4ny9kNPZkoevFN13Q+QrZjN
kHDlM91D2QF0R0TYweT7KBC9LVuecMT2E0GimCSOyFfFjLQ76BgTM/XIg3eOntyl
DCn62Xndf3ESnVerSB1DK3ScVcEHMkdBeXLeoPqHeVtg90OgYmjKlkmnjScCU9Mw
dAbKLCPqRQfR3YJalIH8HMnWLZCyW5qCnU+LelG9h2Ky1cY1qoebfXPkidWcvuq2
by6HOUjfIViMgVJCxmtPgFCnIt0zJW8Ly7qkFuDh/JIdOcs3hVvep5BmnwJQGAow
QYha9RVLV96n4emhFw0TF6buWEjZjLSxpiHTDXVOrh5Zdseflx2mMb2WHsVKnPKm
FBicgHONdYfYvt3h2OCT2bMxlpJnCNWnnKAfrE9RghhB5efNa66uqhF0K77tpBm5
tBGlwnttxMOxWjSgchwDQAYM8NAlgBFAWWuwKx+oDDdglz1tUGJwoqPpzGQqJoTX
l/UqyXLMDMZUQzLIatxcgtxgPtbTSvFfaL7Zok2Nt7hIE3RP2XG0wgl8iMaW5gLe
B+Hq8dl1fqo2cyzR4QrjcdzA/GujSNm3P57haZpQaHH57ZFrqU/jmDAe3th1mlrQ
RfmHb56pmt9mW88pc9bW3FSXe8CT/TbtYZRJD931E9O5f1YZiMQgGneSUOtM6iDw
mfmM+3wfkc+eZoOxi740I25Gyndwd3Ujm42qtJ/Ovm+XQr4fPv4QIKknjgkGuFPR
yLFGnvxaGUy81b/Q5ZC5gw/CbzqyeAymiAsdmVaho55ocg9+SXcpxqd4I5Aaa+Pp
tMq2QZg9/PiRYt+LqG7n6G4Pb/GE3b7OOCIFdxL9ybSTI8q86nMT/8VL1cWs5THS
gNcQ6K10BKxvp1S8g8D6u9XFWW8i5FKXEHHJxhXI68GtGnadl49z83ztr8g3pbPg
vofsp96/egxARdWR89ppUL2YvgdbFELRC1lmZIImcKP6uR+sHtzF+MrlMsFaaHVc
b+8MP5yvDy7PLGRl0rd8syAQUmVvdc0wUh/kKO5g8WiXdiCgrcODWkwyQTHZcRcv
kyLkxs9Arr7dt+zOW8l3bmsIoXD2367REI9ytgQrPHFdH9csDDBYNwKW9m6pJYM1
x17lyyPIzLfhmp98McgJ4YJ54vSCzJQHzgE/aW5GxD5xxYPlLnKfWg5sjOasYv8g
k+cZDOJzhbtdSKAQZK/JnduTCVuUr5/0QyQ8Zc+NhI0yn9syq3HrdCgaJHfTCngY
XFyGBUsjFWNno/V1I9TRTH+2kHzBPA7FP0YD9YlBt59o8jXMQv78IDuoQy1SCitq
7Amnvux0OeeyK2/GH9cZl9qAxxqfs6uAuOBapS/hqbaCyVQoR+c7/1MzXvE8Qqsr
g1f8Ia3oK0ZjhfJxo8l6WDOxVbYk7Hd9ivVpJ7iix8bdXJD/g7Mwg+e/xYJ/0sHR
W5DWlfL0GhP6gnd3hXFHQ8BJSkTiM3sq7vwSIYnHNt597r6KseJvT1yKa82ZHG+V
lJh0Jyh0KH9EQyXu0hq4JCJ3avngEMai9jPPTTRpcTDTb+ujGCioJohhosfTkHty
X07uldAV4edz0hmyGmhPTcCtKZxLIO3ecQv7DpjwyCLkZeRJ5HiZ/3AwqHt/XUB6
btCPSJT4Sc8ti/WvCelV6bX8IVYoSDMHIcm90Wzr1O9mlj0T/uIEnW5hIoTzCMbi
T9vpSEteqsIvG7gIMbBUnYkpcif8j4SQNvm3eqAetHzAc6m6T7Gax8GWjnQniyb0
RXm0V5JbAh/YCIX5JXVQ5n96SVGTdHjECB3I2PhktzLUqSrnSXInobqw5oZhanN0
3jY9By5bp+fAv5PYQMjARFeoz3/+35LPB2u9TnWoLVGw/sWuqZY92GaI6ZQWy4MV
qvGtDYlu06E2NzLSH8K2n/vr7Oidu/dv2BR2bl3HloXX36+ifW0hpioBaERdfibp
KG7E/EIB66NKNjgsVhCDnXuRAJoVccrnnWgtZAR0hUpO0g/uxKdflItKR9UPGgJO
Sp92N+RfXXrd+/+3tJiNIK5Y0oD+TzsHsv8xgqTV9GFr9FP0QwliegVbe+wPunYx
WP0f+2qEmoPsTX/ZmZPCshe9GzJdqxMVSQuxiaVa2s0zZWqC8armRVyGm7UokMwB
21g+NBSk+DM0nBDgQgUJM4t9NVCgpJnxlUeEPawrWlNqtZd4Tc49X2mT33IZ4nBu
wQLCH8Li+TueWd5bPHfKrQw5oh9zpdfl3yGGnSvbt/xAxvJh3b7m6j2aE+ry5oct
hvmfFnDcmd+tAqqg5k8sun4cEFrKfsw8uBAYPW0FhsDeEfg4gR1u7/GZT+Tk0emP
TXZVYzcHW9uivNMAc5Hgh3NxPQ04Q/xk62M2yxzEVtdKQIDDI/S3FP191Pal16Tg
WDibKZ+++ViM1OmMc3pgAOuqTvebVmXfFfeILE7hkFM/cZyFRc+eNecHTRAJ+AEy
VXO9Ak7X1nZ9i7KEadFYpBZ5Wgcr1vH3rJqcyScM+vJjmgkv8KgJqWRdqqjxGKOW
qwwowcWvzFdReaFtBvrDj+f9S1i3e8l2m8uixoZIwqb+tADVcUTTVNMy73D8BUPe
npYJgGPAXEDDoXbMPf2tkJ+mEFwzngp+ToNzdsLBXK20vdEjwpGmEU9QWDN2G0lE
iT1DQ3y/v+avVbxNgu8L6l9vBDUxQ4Oh0LajgB+DzUmkKA80LYBv2t2AZimfh7O3
CHHsYQwPpBmNwvTCKMgeHXbG9jUD1Q31M/2AgGrdBqhN+/7fDKNNvsON/0ngixWM
IB3Jv9wZpEdIUf+XFPhFGIS7nWpe/lFeWenvBepW12KCcuVYDvfvK8fq1TMuLCpp
MuE0lE19gOqh+ivlehq8y1Rd7iVDiRG1Wl9bR0wNt+pR/mjF0iHuNgZhkmX9ll9r
gCjDXiJZlKmCrqE+OP1zvw1aEKgiMAYEdOgk67LaOI2HDX5c0AOaT53LtWGz3aed
DQOS20QFz6bNj9jqIuDFrqK9PAU3MHBqJmSL2G7Pjm/7n+5+dHYcKG2ULu6jSS29
F43/uAS8UFxOthbmTja7TMo9DrjNSsg9h0buein0HdhkjwkreVs1AYv+tlj33Ovq
m0WS5j1WBPkZV+9Ov0bYxHJt4Ie0S5+QJZgyIWKB7hNiME9sGmSarscgQ43cAVuM
gSIzex7xMCR+YW2168YsGKlOf+IdU4x90to37idM12MimzwnXBxihRvbccmh+gzq
kt57iYSoWmWQuo6D124GmL52FFgUWr+M1TQ9stUodRAZswmxrvJtTgtIbXCEO8n0
+ANBDAyA+1peaHww0reORBZKjtUkHjtrT8r9+1D2cpllij57spQ9ELr6ub75kXnZ
EjOlXQsqsRISLrgZf6ctMaykokCMSLNJPwHRtamkKMhxwPcY+5GrzhAfryHOTbp0
rKGJaIFZXRNfVb/nY2FStgtIp9K0j0Hq0T5u0hLwX7v/ZQ324vSGGlvrNjypiNwT
CtemBazaj7ax9BSnjLOLogXU2d39JOr5517kDAKnCZr8mFp5tDQqzDnGsklfsj4O
lR/6yF+siU/p88ir9MjybnH+7gUqogTULjOXycKl3ewQK0brkjz5D1dC1m0+jKTc
qQxGXnVL+5sB4y6M6NLWBJZk1tr3dRnrD4AaYuqXD0hrsyAme+wDuRTjFrGXZXql
cwELaK31kRSPdzlFJEaEOhDbIDKxhNtiFSXWx+4MRsXd1WWJJsUsiBwxTTHHfGqe
zEC2Bu8X1GOvkGPDZW2E4A+GzrCJ69DXPiArp7jD/kw85o/QLf3ZaAjPT35FZtS4
QHRDWVRPMwVm7hRQkuwuZWjeeQtSFjV7GDTYfoEGAXhRIZUf6ab228OFMChmY4Bc
by3W2epylQI3ouZdjztU2p8/+Fy4jCTTX6dpfpDz1BkV8AloLtkC7yeey4Gs/fwT
903SSORlvrbgiID9yWx20ga/9V8fnvmmnBj8NbhWnyNxQ5/AzI6oA1IwmOeOkg8r
KCuGAGTto5W6MkTLpGVJfx6W9pcOXDxqoKYbhE6CVIyTRYwTDo+ZQlcfhjYZbnqK
JLOMd69CSrOheK+8m7ZdcnO7swQdnz9MyWezTFlAET2QShmtN5+Ss01+5y8P+B+T
N7L4LtmOGy5TO5oU8cuT7MYF1/yOiPZByetiy2SUIlgTVWvX2ZqAkEOaVDdSUVeU
+DjE5qX/EGctM5xN3MfvAIAG640noVbwm2ERI7mYGEpinvBkmqf3A0BT95Uaz877
gJa2UBS2LrXxh1g9OrIqttjXZQTD43cN/atn4i+k8+Mf3C2QUwKybBSgjMPkqUS+
brs/oStTiheLbcY6eA5SLGqhUQw6bTbF/74AciaZpTnWw/zxQHJxwMfk9Aybivy4
SJADoOZHWCWAp6fyLheVLX1KLoVNgQWe3lBRt2DxMNB0SJywSV15rosMabjFJBxL
3ARZIvm5hmlaFhR+AcNGyYChkNz3qCqxVJ8sRWigLZtBCDW0kqG3POX7B+oOUMaP
q88iL19DJf3NBwoHyvqnPPY2tRdgbLyZXjJe3S1gZC9mRDrjpsIzfeMwPOBSSbei
x/xaO+Ebq3HTSsZzHwjtwgEL2qBjiedziHHgo6AcumM4nBqpt5HYf/VU2IVszO32
qNUVG24X8NkwF9uOZoGSaeW2Aghi+YMJwMIPJsplf+NveK0rrEkcWnxkCkW9Ov5K
rv9L5+/gtqxvJEGUAWrfh2gYa5bJ9d1Vsvj/XcFUd9J3Rt8fheTd1/II6q9unkOm
ixm/NvQGo719AAj5RLz8bfmmwzfCf9UJOQnZD3ICRzjSzYq69rqC9W0W8LAdPHXM
MNEktI1w2FrBcZBZA0k/mSX4egdTKBTPU54MX+7XeLmc4Ropu3cm6V1ACywQzLqw
8Y3Q4kklaWgTCKOvGwc8g2/f7kfE2sLZZq4+MhVotDwz1Z9sy2dGgTbnieKVTFo/
rlD7aMj6Zpu6dR9MAoS/kn7lmVVCDO09joEYzYaAlUqkjlacBCIuF4acJbR7Urzk
AOF4GBuC/ID1ny+lAyCm43y26bFeld2S1HKkyeKwsM921bTT6FkCMgyI68JDbxOD
WDIktmugVqQpu2ewbszpsk6kEME0WIwayYaU1zTOaqkPv2k+SyJWl2YfSJ1Sa6Cd
x8gph8nEK51432CH7XvoMg0NB7lQ5GBUkBZ0qtI+AuP3t6ehg67NVIbIAn4XpZme
/DGxgiWmiJy5UGe0XHP1xhZXIgUCQjFUbhJo5I4OZ0jICF+9D0DTMHCFEMjndy4s
7pDEZTJTprWeJRxaYgGRcY+1v3H3B2eSCoynrveakiAuhsnVsT14D3wpqb9UZNzY
iI6vTMP8QjUYm8el9HSGGbzL8zVrm4QiceVMh4t2KqM7YCx6pETsKKVEy3w73jOV
csbkO9mbDZOA2+sRo04IEmgMhm1b5aFseUUEl5T2B+1HwNyejXeNInQ5LnXMLo8B
oUq3IF+UntqmTLbHJg+5GWiF02EVp0/GYXqja3g2kI/iEZiQkdSlmeVD6dk0bh9p
hxWnLM+lmTO9NNrOSjNfYH7iKhppiZdSNhAWI39fkuOJqvrs1TB81hVinIKFdmtj
5kmb3Nr4v2O2wpAD59YhTsO3H8Fg/A0WeEA7cafKocukpiExb23FS4pIfP2vkaz4
fLC4X/BDSIMTJRpR2gScuctBs3tgYBOg1kRb1tFXysOeOM6gAo3I64oidev2tcJo
AOlsd6stpddiwr57r6jxwpletybEdRJa+oyXqHcr56bcxGw2w2RJJPZlnUSOjxqs
9YFGeN6GWfGR5O/ljr+2ALZr85tuSgMpwrH40lSuEc4RaHibxxhEpJQ+oJCyDesF
TKWOKFudgnrMTzb5MBj3SoFLcuy9zsVHzweTakyAFcaxx2FO2Gq0ZAnDTVsoloct
OyN5H8vwkjHOiVfUTR+xsp4DSHgF+ai1r6lTwRtFawrjNAJXmzb0XEh2D0sqz1Fm
ZIghHu1bhk3Ag+umPRdeZppGYaWIwH8xnOIwt103X1Boy48+Yr8fPHbuYZPRHqKI
URnr1dC9B1pWK362s6kc5kkWXBsgWCdo7QmL3IfpvwOtm0l8/CuK4MUt6OXYtTUf
pvX2ZQSyr3hxMDRCZ4kBU6YKRcAdpS1oqEtEkFKYxOp87v87AYk3H1O/MwkO+CKB
nrs3X1bs0/FKG6daSEP28ZKeZ6MY4JgrBH/1nQtb3uJZqAKPrf2f1gq80IVIxfEg
aDb1nCLcp7ZnayJMs3LDJG50WEMCX8mfFO0huzZ6PIp1LzQPa23hlRzmwkSH5lyX
Zwecp9CHXOeseOKieHR6EJuP9c9zn9fcsYMR7wcmKgl1n+KiuIlzhS+G9QsqsLOz
sXKbgbng0VBlESIz8Xa0ALX8bp2RRgPM1PO9Pen9jHxVug1nIHIQZCtqeNpSNk5G
qyLKfbahxotxTHHKdsv24MKuDQMt19lCtluN+CP/uZmOO2y4YkVuWLP4C7vemmfx
5REJJYhkMvB/cIfFtMxK+OxUfF/ZlOevdzo3zFHTgfqoK0hkVtu7vVfKZjbVV4U3
jqTxbcBaPe/NPYKUtNIjP7oUm+pMbEQ2bMTKQAl+RxoSFpH2NAffBNZWTx3JFeaA
ZlayG+OPZ90p+qyJOv9U5HFF/vvsexdLC9L4MUMHGy4aC/8Jbz2f0E8lN+z9Rh/4
DxmHyBi/to6uI50qYGk3LiyXc3ZrHJLJCqxi87wCcA427707RJp5viW3xGb1Hd3z
5pUggTDCRXgAsaOJyso1+XVskLJ03+HHGcAyiaV9dBxY4v4IsTskmgfZ0GfvRHEV
gyPv5zonZ0ZQODcjR6Q+9M1IHRg4/ul3oYj/DEvqwZjc1t5rGbeo9VgTS7t0Xjys
l6iL/szB1+QnsB3QUauKr3plfxe5yrDN4JjZf2B3hA6KI1jkRB34pSj6bnUmCMbx
d/tfe+w6DiXLJZaPL7hqXHw0uTa0Sl/5lIi+Xc5kH93T2UaXzsXYe1ev5LibaBlK
F+VPvBr//IZaKrQiV2Hfi8oTK7e6CnmSpCWrND0D+AvZ1p2fRZAdEWKcPkDmvrlx
KgWd2H1f4Iy8kMf8T1lLEb8e7BOD1WVXTqlhFnnMRjMswqKAXqBq5+bjEl6q+VI7
NGDRjx9LnYkAkMLLl+V8hEox6is8MSOswvwCfmYwHDgIcMJzDIFact3SPv+39tph
XX49WKZumS3EfR/FvB5nGU6Xeec3tl/GRhRbz2oc+BNyj1Accwx6hrvhM8KeRmzM
V8lnDXST3qOyMY5+rCoKrTOCi8+m1y1e0AX4EyLR1K9JhnzR/6uR9czsGk5DKHcW
AFSGmUn6tVux6am8kFrdBBZIwjC9L75SNzJvEdMFspCQFJ41eftwY8mWoywxH5s/
7G+PyvwLYsLp2zO9BbXOwAGBH5eBaNC7KIBlIb9rVSAGgpgGLjI4i/q2VGM+8+ar
1jpkpvtn7fy/tr1kaM6QQNkgm4LoejM7xMYEeIF7+VRDFu7p8XhB7kWZMQZyZnx3
WO5VHJnVPNCXhu1XO2o2X+agcmDe4AdacIbL9XF7gmdN45RK8u7DR32kXdo0y2g3
VkaFemv442uctwpJmODQHOpkB9c+KamA0FKdS4nk3AqTHzDqH8IrrkDf5s7qmvU8
aduChvzS/m4cdX94q2F5ddm5mom31loAazSH/6FjKP714SXutOq/jleWHmHbvvdc
yyJqeL/FUsy7DKNq+MjtdwUS+ZkqlNhV9VHZSVaORsSa0AlPcR31Mm0vZ17/dAPm
ORdLBsACNaGJdF2gXnQRWO7sh0nEQq79Y1Q6JlX/ZmlgKyXcJtynFbUGyw4OgcGh
NbmNCi2T7JyTmFrKQ7oE1+xldVs5BQijNQAUqS0W+C7fPEyQS2TaRcaB3suLkL2n
LYwCDJChwp4FcJLxr3d/R0u+6Aaz8V1x9Yxo1PGtlp+XRggif5nQRzMgvBl2SrNH
jiG6ko/MIWi9OsI+XlilcVJSVassgpx0UPT7TkRFXIxNlwbk0Xk9wjESjPObbL7M
bBxjY1w+vN0xjqMvZxaBzaJ3hbkXkFl0tFqP8JYXHz+CvliRDNnl5bA9Ris5C7Ma
AYkMQq+dRW49Z6GIWRkqRHRxL5OPQsNxMk8gCfWTOePlsLE+gd/vAcUUndMEjrvM
uNbMdCkCqhk0vQPw0O1cApURFscTKbWjGAvQXvxNRZXAzvbWVrf6Ah90oyisc0Ez
hiay+SFmWRmJMYvr7IJHkCjCZuGI+xE6flHEQsX7QBwshZMYECxkoc+3eLpsAuEB
Q9fHPTLY9Out4Rc0XpAa9iRIckFIn9ZETgBQs57W5SrPBb77N9QHCK+y3k2UoHft
`pragma protect end_protected
