// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aX7VS+qIy4YnzKoUUmESciNKaDiLiK3PWuWUkqM6d3tbvGyvXGafKcPFFE1YD2JI
mnDoIrU/OTt1P2T3/FYA17h7r5Om9U/gZqdxUYuazT+nYHa4HQP+CqqgLBZDsV7S
TEKe2oQOoR14p1It+UyVMUeaVinkWfBfse+3T50Zwec=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5296)
D2u6fpGrf9/D9/wlx87wfQuDJ9U337WA8jtzkmecNSDxoNw/xlS7atTV9ACiMxme
i7TROpt3HVYvaYIGvgYeTa7QVkl4DuwqqKgIC4NWT5Sh+MUDrBSy60Y2qQ6x0gz+
Lx4vp+2FGd7UXimICsYUtUULaeEFGdU0faZBC+EXyuamGddIYAC2izdmygZq+/ZQ
PtQMy7kUPQMRZ4XwO2fC/92bZVV6t22F5ZvWpQ51nf1yb2R/M22SyKPLfcIoYLsm
oyQJVHmSovSgbewBsxV6lk6rWbCYV6EjVG/7BqGzARnQh/nnvJD2bQjRF5aTyiTI
2f9wZ3TvoNdRv/QNpfiBiX++5p9eNoJ4AFFZFFeGIKPfMPLCs0YISGJ0R6IkSk1l
6LwEkKk9G36EgbfVOpFbPmFkHoRPkT9KNS+d8UlCTElf8Q25ToPMQZrlS5sAToJd
MwQVh4IfkYyMYBUfgwrNq2yPeqVJVZaQOSs7XB95zrd6d2SHF0qdjK2OGDEkEpZ8
6gQg1UZ8UoxKcv8tgUsdfZmiHie1lwKi4hDprj2OP6ppQTFo2gAGp/b7bo1IhVwt
j7Xj0NQLQ2UGNedcXmqeHlqQ9YBgAm5/O/CE1L0h7BrwvJtOGrocc4pzxNbjHdGe
utboQHDlIK+n8958A4y6TnixT9vIf2RFy2L3Vfeq8iuBG+lAOJdtuTwygr1CJXv0
gLphsIz11khOcJ2CPfV9APVq43zsBtbGKy0KES8gQGQ8RFzgnxcQvXM5xxOcg0AL
KgVvc1zeM7XYsL0E/Y6unyrykWmyCPSqtI0JZ1l9fSOiWNJEgpv/EUmb5YTEFWVf
baQMlqLTrpDa+KXuUiKwYhAvdLirVsaF2+aGaNVqm2O5tyMpdVHPEZqe5zdI4KF1
i/7h6YlxIr6KP1oZpl9vSxxMFmuyGUsAjPZJZJf/xgh9ZCVxk8HCKG9WostzBKj4
dZmwgCehe5fIfx5kGv53pWTJmEHIpJoP9tNEiCoC2fQH5F7zYRvButtrtiAfvIEx
ae9WnMYSoVEBzKKd7yzHb5ALknQK9Tgl+gUKFjzua15EMQZ/wXL1ETvjJ2iv9xJN
uU7v84clpy0K+ENXVpcdi0ushp0uWxVQ/bnxIEfa+xTI+jeYGLyiRGXVGT3dAL55
gQ2kkOjnvD7mY1jeu4pou1ggWk+CrtNosEbi81gGw9AwODVNUxeu8H//o5N7Pgp+
AXtxTQbkSMiM42DnkNX31NUYp8U7VNQ9egb8PsaO1cMSZw8QOpCXM3dnHsNDtPrL
Q4tDPAY1eU8bo0Xsp3TqAICZXywI68pnn8qv7QAey2DXTwhWCYHd/oeDooCTkvbo
UDcOTYlmr1RaTqKLU81wbLO4FjByRtTuTy8TWm1bTa1hvCdEbnuJ089RGEzfo6DI
lDKpzZc1soznzrn4VmK3rvMYF9XCD8MK3b0y1FoIlj5oMJzRef0M6jRJ7oXXT3Vr
/qW395U3Amp/LsbcMtYzB3hBT3kjXLHLnei5DPEYOGFYz4BB3IRaW6PvqxImRJCh
WnVkvXOa0FLWY+mFpqSIz2b1YoVOXuiaiVv3jPVRw+fGeQISEtjGpwIbpSgvYb+8
1v39c+HNu2vNO+EKGpE6ibzMTBwnqw7HswMtymxx1n3WpoQ/XPehDWosc3UX3pK1
sr960n9SX35IF/Xpn2YOs9gZgAsK5QZlRayuH1C3+Bz7iqUHbWmIt5PdO4IKAtkA
pI30zfrYBUjENwsGixDjg9KZj0tUhkf1U7FjPDMBk8anSBQyMAY0WNqin1Ze7ouL
xPHQhGV4dJhhCilVKIiOa2zs9RVH1iV9ahutFGAi8mjliRPbiyACNynN5ggccaIn
EqxcjtAYYvLu5c83gifzBNbqe7Ay3ZldHKpASM+IIN5GmhWdzel8i3KJrZux7VDN
apBUb2Cmb6PsvY9aDUquD7L8r59qYmJ066ncj7TJNVJirCKfSYyaQpLhmYkkGN6D
EFuvyYcBc70f0eLOlU0OQWS0wijDvR7GQAAcFw/cwC4NmcSXdppdSFyhZlybQnN4
eUFN5SLeUSG7QBczypYw0S5wTpJEP0b3GWSsFCe1vqiDzOrTu9AWumZGAPasre2/
xiQcA2F13ssxZv9HxRf5XB6w5N0fEueuc2y17CzanuRb76hcO3/AoRn7dSM9KsfL
0kzc9Z7lR+y2dNgp0UcHhsvyv6PbK+3fLIcY22KvyY5iCDB6L+tEhxZoZAHyS9Q4
2u1x2P1eDUTK47w/WtSzPyEn3EHtTzwYS0Jx5MXdmYDc1Jsli+Lsj4sZIfAxInuW
gEVCpR9eQGkrNMYiA34a0ei6f7dGpF1KmGAA3z/2DUOWE88bIPJcmPCzI5auZDv4
5E/uf71dalBvt/CRgW/BD4srWaNXmgwsX9vSRfN4u7oyh08t8giJlrG+IcEqh3pO
0XC5V2Lg9OATNgWiov5KVS1r/1rRlOZh+jxxu7v8j3l5lJn4k3964P1tJotIg1/s
Hu37USs/++FDVCA4B2CgBUjx4w5AxaypqKqQodtpcLRQDQBMfvkdp/kl2KNlX4Dc
shnw0Zv1J7Oz92XXGQuF8Dp6mX4/Xw3KkunIAjOt6rIum2hQDBI2xXhX1RRT6ciN
m2A68VTks7rTj77kKfAtrfrB3XPFUTzdhajDwM7k3nHROZdtMMZbGPIl9XItaANS
owii4538AAH/Y4+Ao3tIU4W+vG+3kuFFjqOjCDF/X7ZE8MhwaYmZdzCN6dY8Rsms
kIdX+Es7XNErJrnEyDvuAfIP0VEenAjKtW4B0aGM38QysRqJYIMqAgWgo5HXoUB2
8106T8zX4kaCJE8G4Z17MTzWm95rR2RPt058K1ciplcVKuLvLj1NDwsAed/A7E7U
Gsm30sAgMXB0+z/SM4qiWqiLI0nhv0KFXYn6K5ARNpRi453e5szAY0Y0WiBXJFdK
yMQZCkGl1yxARvKrWmPoJiGTfaONCp5681e5tJHRvWR2Tf74tetazowHfPItIYS5
glHCtsv9uwGhO15pEdtLvUG+PL0QR1v+I+zM28jzdp3zLSkI7tKbxkqLmRfN9u8L
wTL63pmLSsJ47jilTZqiU4t55WUGQeJtTkXGGAeURoZtd1OyiRxlXYdLlRO/pjyz
pw0OMp/Ki1796vbFMeEY/39whgOhM/4iaDcd5XmgMdbTqTsZKZVs7HOTLAzNjn3p
p3cPDpYT2h0eLRvyA86Tp9O+kiyHKoTkYskdqusbl+bLoaegAZm+e+Z+igkL8aNZ
Iqbjh6nj5ur4cqvyk4QFj5ZiTsAm3QvwMF07a8zRYkU0kfNqojZMa+AI5tf8Ersk
b6ChTk/xYYkO3DaeHEqYkSfWUwQpu2+Na6qP4jijLAwWT+aA8Wz4nIvO6RPKodJa
9lr0YfXnpOC1LfBLmzs6u2ks3Fz4dk0tqQdqVF8/puTRw0P6+BiEvK5x1szBC9IO
hmCAoZFsxKnGKyXbt/j1m+kzd58zvBHlVGjeW1y9XBNDptXOsw0XvFTcx7gbAD9w
uoifqgr9Q5aUNc02E/VyBcKjh2UWMGlFNJ5EbfrOicar4boJ6AWMrrmcwYeTbN3g
49M5D9xsi9iqS3uarbeod4uTcIlkuO+JibIp6UudV6bl7vrWAqTgQBkWFnE8sLU3
ynOwuyQMiZcUm/Fy/f9CALf0xp2V0YjrZ12sZIRqbONuPx26q598lb2Wz8en5vZ7
Ty6SJC87A15r7/lYJ2X8OR71ESVNYaDyT4IO7DaIwWhz+WwumvYBhNZ+fL66EzJ8
PsEZNyMreyBtWMti1cqWtnmOmgwFPv11ahIQpAgWzGm5AXqTC3WxB0ccVBIN3x4p
9pIpY42FZn9pmx+nQurYvGiVbfrxpGSqua5i7XIY3Pkb+lhetMTEwisEGsBgp6/t
1p9ZCRI1wwGPWkJcOcY1Y853vOLoThKuGirttLUEztF9k7MqR6CBwH1JIHTBmoK/
9CKY46d6OlvLmev7pRrJBSmwjdyZatUVdEGCp0BzfMofKTtHMiySwdCPd3uFJW5m
vjgwMraPVzZsJUPrsQAvo0tcOOz1gcxRf/XRYZG2KR2/O58SzWxwV+EabAXEHOVH
97Nc4ph6B6G5/7lSYOl5S5CxJqy3lGV/Dpt3k4kwBbGoKimFDUSCHsDvxt5kvJAW
dnSQnRa7jTiMFCLrYAHYvI9eVNus75lMo0y6HoKbaAfbHOGmPBHER8uGBYwMbi7k
qC6gGLb77zbmGG/mU9UfGoNIMsr7yANr/6eTQxLtAXaNXfajiOagiebifIkm2r8E
fM0EY9bjeZq4TFLvwmNC6iVM/etso6CVvlDigcvW542hupnnu9fnjHVX4jU6OkZC
HnNhUovwM1G7dW6r7btpAoWLJC3NKOvUOtyJPPgrES44yphVmj0rXypOj0ISflsV
DwrOMZIbsAIVmJMtNgrddV70ePLKC1LhFPMdxNrmZahPskAm5XDcO1WeTOCnTWbO
yRdfWWSDwZOOKZYptLxQ3aDDYGLmAarlvWGDRzs2gxT3+rKUNObfhK/Z66MiCNaD
ATjyql76gBG8XZbKW3tbZVZic0tObhGlbckH7uc+cQmiH2D44dMREQgpBTZ0O6+n
rtxmzzoM+vB/wv0bp2Zxc3s4a5FrjLQCokIFCdZbHgW+/6QLh5jL5nraj2FtgNEP
o0/lJAZcVxMEzz2+3O35l/7CUhkeggeJqZ1g5LTpHFSgbUZJp0LTUneMoNKrDBtq
7dUtHSzHowd4ZzhLhBwxsSgDwQX48H8lxf/4QVoRynOcDHG/W6tGXSBWgVBEhn8k
77t/jIzAQeH/qdk9V/Xr3NPETLG6vaIenzF+8AoCPJp15vjW/LiF588tWT/gv8hx
Ad6ZCk61/uzx+E2yoX0dYQ2uOoiIsZSvcWnPvgxI6VWbketpeYttL0y9A5xbS9tJ
+2wPy9MNw8bmCsrfY1qmv/5cf7h+R4DDY1TJ8y3BSIU27U6TYZx1U7xeiDt7Rie/
WxD6PaIl7A+B/6dRarmLu3O4GR5l3oZ6ubO/P3EPBlegWDLYbjx0H7soIurh/TJe
QmFynsKsCMsCu2nbecCDJJULeiXKeRZzwGUTGObDziWKUMkbFumNJtrpMcVdU8ED
HiRc0TbgmRO9cdVHE0O7CEf0UzeKUnUoSgHrSBiNHxroqTO16BdpltWVNj6MTgFi
ykCVTQKIKKvenkAs+E0uzsJmWLzf0kvwuuSgp7xrPQooFA0GSooEouNyQeI2g23o
+4kIqi2QeVuP2b06KTD63CsA/5c8Y1qqHXtocQfcVpleAaGCzwGKwnIBQMUOU9r1
vnB9KfTL8miljgH0l4CCs1wSqiPaYoxCSDKJ942b4vNOunjwg9EX+lwSsnTpntG3
U8o3WLMW0T4QrreQekNDxTgFHhX9oMmTYIqM2gIIwSGL4aJqbS92JXEe1mD5iEIL
7q+jpgGmhJqs4EFP2eGnYJCCTuVlmlp9ZpkMTweJ7hBbLxVqA8zEyQ+oeVVfsKRM
4yNgaXCzWbLokGiNEGXsQ4BgszRpD7ZGFrC+usvohROHyWQQSKtXTdlzVaxIErhT
/Sfrp82qJzY3QncfDSd+AXB5XKsmacTGnP0m0uSKz9LX6n6/PL6k87WN81mXOIdy
hgNNqtisZAylD8mq9xF3FCItk/wgW4DMObPr0TX34Zinwp21VrdcpQwn4cRAMC2E
V8sPX/fPyyLd/dFoiB4n4yu5xYfuLTyFk2cx4nopZNthCaCQ8Iso+rWG6BTWm8di
GG8qeSLxblgXKN/jPDpTu5wZPIBUVWuusIp9LshbJHzDLrqmsVzIykp5LRChFyvL
lEfqYmtuSnv67VU3H2OU5gbVoUar0g+lT686NoZfKG3QfIl4Y29Ug6MddWEuy9oU
7gBVkcy/m+h0Sg8/yVXly601v2qJxM/PRpuy8xwE10IiWnqkr3nbsOmwZRhWXD7B
nBUShF2mx4QnbGYM3yflqQ9POdmY5Yp+FpC8ii3j4+1I1nZB1/g+sbPUVwmWvoR/
KnTf0RABe87jUeTTKUCROhS+ayk2eN3BsmsSCzFWVpXnD+SUvRF/xFJD4LIjbo0t
T1nFGe5j7SDeuYQSs1vhiGFDOaa3fnzNc3LEeHuIXiO8P0dtTi96TaCL+YIw4rNm
k75KVo3DA8lHixnS+WWhv4gwQL8KsS5ah7d8xg3C6UxCSzz+WSatNZduYy1dpg9M
HGlEdqf6E4nNB9Jui9OYhQXg+/tR2es32AtfyJHRIDFbjii1FQ9p5Ms9XC+xxh9G
kCAYhQQsmb6NfR1OuS4bDrPAXen0VbWg4IU6LUCb6MQfPK4pFRcB/7IcdHidY7sr
GLiUG9TfVq5sG1ii1OM2/AEJcCsnzNoUKuG+tvlt+n6/3tv9U6drKD14wGqMSMIr
UQseRLiil+ULUj91+PJzTUCrXUFEd0tRWNTOs9ETwTxQmhznbIp09tnISORRISNE
HFxK34p0NIwmrpmbs+HorY2GPcnI3LGh6QRS5riDUK9BsmC3stXznjsmUiRlZaA+
uxmUjhpvMFqly1rK89jUn4SQgCxOdJEnHZ17vkeRAjfNf/Kph6LUhHffu9WjNCS9
OTT3WQ0MHZ3qSWVaq1y2ajjjWcOWeVu2O5xR72JF3eVfjaZpZD+pmHfD13G0ieWL
ovzBuHRU2bGsYx1B8qPxvuFj01GebHxXPzqOsW7yTiOGfMjujzDv86F/U7Q4af6c
+0+ekzXc/aDfWEHUy7lCKKsXWxptVRW9N73SbuRnb0DdgvIyY5WBlrRAKUNkCfS4
4rsy/0Y9qhP+s2lAkFiliPFyjYPUiXXfGGsvie+MSRMRDA/535C3oD+QE44fqWRV
1u7VQjojKCmX5nwDnOEkRy3EE138pZT4vY1lHGCU8fb3pJoDIerCusnUuWClcoyJ
RYW/afYsOHd0eJtG+oRKNToIRgPrINBT+aIEe93LRv8eVc+XQ63ciw+KTz5VlRTA
23+ndne3dQUNS6rO872DloexrrJpwdOTCrleJcVTrSXEiKH7sqs4IFnlkKIGrBh0
LtNJnrFKguPKmsIgI7LYFw==
`pragma protect end_protected
