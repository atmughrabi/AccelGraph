// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:36 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MJqqaXPuKPGCde1KVlvi2mi3kP3wJLafaw0642nPPs3q6WC/HU8SRjbxsezskGGB
rOL5tBar6YEG5l89L/nxIlA5y1VkUlrl0cLpkL59UO9/Xyhw3fQYxuV6gmNXGlau
uB1y0sSBeChnJ+mBvmr7OaKJ6gWb83dXTLX5mwakrRI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 54048)
6YwbYmOOSXf+/gxW88t6SsCx/5KPoGOAX01A+Jo00x7aVCx/fCzjfgGBOfQNcjnX
ek3+9ZiKwlXGdM5HOiQG74Buc0hQpqSPU1SCeG6RUAUncIWs1TdK+ahtBekMvA5/
Hm7gvpD0eytRE3U/HOQshaOeOmCQJVRYq2BVzluD8/RJUFcoO8RviyQ0yZe1plnc
OzezVG+d7reTzNvYcEL7C0uY83gCbd4kk/PJD3uetm+x4YB1GU3qJGF9XzXsmYV1
a5rPutls8i5a0jt4dijkGLq3Rg61eyhGpU6PWi/KzBtg4QZJT7Jj0jmPbtLtfFxQ
m7JmQgNJWCGa6gLaPlY/9A/NU7E6Vwyw1ZDoaPLCv743jmOxtS/mSAwNDBkhc0l1
Kut7LKB9sf6seQkcv8GQ8SZPJBwfwup2og7uaH7Eu37Yah9ymEqOz6z0drlzy3u9
gJcCnmdfjprZaFM+FXPI/pz2T3AU8mftRKZtNn3ajzbtuDdwdvJSXngDcPJ+QNp0
wqXe5HJ9Ln87YlzKk8j4gLgXXTJ39B9V+qN14yOnVeUXqDSOuTKdbpc9whijmsl7
aNeNYj1OnzOflicB7ttzsgjdBAmCF4W7v9X/GPYZYIgFsPIQoXwR4TBYA6qZbW05
+XHL16H99UGivWsMwtC+1MlGAjvLHbgG30l79ZzD5nrYiccsg1RAe6KIX/gPt0LG
Fs7m5hvQTFgcQ9mWf0bNxpfyLnQRRCoM89+Dl+LU+rJNLfOmMvfOwdwGBmIPM/2k
usETFyX1sziX4Q44d12xKGc+cy2vtBKu/E3t4BDiUMIXICmO65yMBE/Tx/jvg4tw
hm4ZcCWqwJx6XX9HBarwbr0IIkRrbzO0AvdDvgB3SY2M4SRkULI7hRtz1zTwxx3O
0ADgTodzJgi1VrITdhr6JtLUBQotHZ/H718u1hzyISzLt+z0ToR6Qhz4bczUtWZx
XKyow/qKMl0pXwtVCRZlqMRimxvvympO1bm1KTtZdK4H6NFp5tQKuN5Q5Bv0pkEV
Hf5PbdgCtYlTPO3It9JwyHf0YsE0MauuzDwCks2ZMW+7SZhtrPA7XCaNJWZnMiQ3
DBK/fligL8CWPTTDBidUCxNdpSPn/IBTRrcUqQi642KmcI+DOGcU5gEitN+LxSRQ
4ZrVi0B/hJRKnCBeqyYJkaM+xau9dOuUb4URGuWghKt8a6HmF49fjG8ipXI17Q1y
BswfFi+Jgv/RHAziGgLne2H02Yxbp1oLYfo0EX6PmZpaHilMK9+y6HfxXcrDDQWN
BcECmLSUyGA9i1rCuOXcQy5UvETSRKm8wnWwbg8MGi0gyTbhAlPGagFqUPnTI1lZ
44EEfN4e1ZYTTvYWxQAFlMr11bkVaOe57o83I8OYBMOeXjU/iJaUj5fKieHpc0yq
u57qBWs3o6yoBiOzxqogu6pVMtdOaqQMWL3Zm0wi7/r0QwC1d4jBhikncGyfPhuh
i4MQyEE9/yGuTtvMqn7+RsjdjfttpWuGnJPK+Uze82dWhIxZ3Clp3qK6QOV+L8zV
AdYIZqJshMAE3F3iFmsai7s8UHD2CN2Pl6bHYPUBDKaytPXcp7KTBEQpMEAff/gU
i0sCj0PPgSOvlEIES6eFKT9/lzg619OJyb8jKvaxSj7C+tGs2V9oGY5Kz7ct9r27
DNNhtpn65yyBfNbY6IAJjqL8g8Iau7pY2AWPYxcjK2rdcO6nKo2/DLBMauKD6oPs
g5dwBAaRNdPRnS290I75zE3NqV5irMdAOmXLBP4wPah18X5G1pN6afyhrV9YpStP
wcjJGWEF+31xbjyg/SXcItCJKbzX6SFe1Aoa38HVDCoHDyczjYCPVOgJ5p9+SQ2f
t94j98X4JZ4lkvtqxQrSB3c5NZcLy6lRo2TKrmyJquH4looqA0J4OS+1AnurFxkx
Q+1Fr/GwxN5+c+LSd5xVXzn6KsvSA7+6FcL2Wul44yH2OrVfWMeaauLWJC72XGjT
E3KWPkVAOKVa4MwlVRXDhKqNT6SxtkIOjtGcrC94GeF6U3Fa0ZIQJ6EFtqqZJYHj
aromBv7+pdkN6DVGRD5zuL+jY7BsjWq88pZIgOUZZ/tq46FDDMV41ip6uZ7i6mGh
OY/17J3rSk5nO8HA1EyFidLbt5thqrl4sKwWc4bNH4jouazwx7r7EJ9cusNolJdd
XyPfuCGntqa3228D7ahuqsr8p2IXRaxuMAOEB/b7V+NTtCdFhsLX0+QYPVT/lvYP
7CiE0GVfYJ1xOgn7vRTsPPO+DLhjycATMhS5yBqp248qr4Vv68ArQCzZhBi/0fMO
zm8uRmupFt7jwaBA06zno8KDlBPZFVWU4qhffl/mKsk0ZDyYQLXIzakDIIZAqgFK
Lat//1KuzAU1C0mrTIdRMJglybaRj86OT2rCTwTehO2JPKogLj7b/kdSHs4cYFXd
6Mr80FUypAY6Xq48wRP31u6dIOKSYp6+jYxAWJlg1Vu8qyu0MZct1EBGKjS0BA91
c1+ZQIO+FbvmPsOvJWpkABvNGWesCLxy6qHf7fCqu51wzDR47K1873zxJYlGNN2D
KFVZggzfCoFiOJ16ycf3Vn+k0d/9zNawRkfInMoLakFEZ7V12D8fvR4Z50OfnBQK
iuDgim32U/pNUFSbjWPF/1MjJ7v6ZsR7IR15vgD2+FixlaodlhlNg1BoJUkUley4
hEuLF6m7+HlP0ke8jZ/ldpyFcIWPSokKsP0pA0TlAph9ioSkIwTVTaMaXh82r6f5
P2jarzoM27goaLg6sPbrED5XePnN8tvpw5sIlMNxJWwJtXwOpUlskrt/SkrelX8D
GPj9uUXQzPq0VCM1NMzRvzYhw3P6Ef1AOCwQjsoRuQ2FrxQvCbMELN/PoVBJ2z/7
ZYRcPbG73ngHE8K14FR7dsFv9HCPDO/VA+JtWuNMRuQRzzzaj3QzDv65DJKCL1VC
l9oN9pSY9aujufADEW02XU3FaMK41UVj3/Tq2BJZU3jeMCLbTxKvCCZ1kpYorJap
OCDTREEdhcLG4gTri9TwWEDUR3lBJVZd1xNb1sYCUri6KTwxZWVkrNsxKEtF5eOJ
w5j9sG/bkOFe0nPIuTIcvdNlViJ+W4Mvs+K3cxnus4466f78Z9QHLVfkCYnSIknU
osYCSg2SIBM33UIm4RzZhIpcl5gb7zR769x5CrJJohyup+16KsfOKLxS5nw0qMly
xUXNNJpV5aXUFwVdN7nKeOV7eWkvKqjd2G99BmYvYkoSVxvjsDjNAjCCFi309hMX
P5KoTkjA2U0yC4osuqbhE03WWemQ4zOn+7sjrO2KfP6uVUNsaEOBWXZ5U4NwW2BE
dSbqZQsZskjCEJFmK9ty+YIo9B7hJaPFT4Du5y6Q8kZHQSA8BXaCdqQgAU/uZQiY
s2o0vI8fUPK/TDdd/v3Kvrj7Riz8JPsJyqbfTh4jPm0WmtVeDUqiLpwg7GWaYaas
c0zofPYdFa+7nP7dsoP4abjMblbJ06PiI+SJVXYNjI3qDMRxH/iKDUJfbiPE2tDM
YK9zftKVafk0fIAtRvfJU//aj/5hmvsCxkBkTksM//9zxIGKP+j0lWsxzF75Kthp
/bN9NTsqSjgXznICjYvV1dgTTrxUThg9rYeNtIwnr+Fuh1ukmiwGosg08R4KKEGe
vLQ7ORTFOzB3dSm08vq096/s8Letd4w6HDb8AD1R9kSNe12/nQ2Ks3QSHKLu25H+
PDKJ8p2PMiaY/rkem1Ew7Xg37MlXElSIS+BugKLVAJDGUdj45/ykQ+9CGjgB0YZN
x01nisVhBUfBzix/CynxFf9uPZIWR0RkXsJz0szQca1gyw+E/y5r1Gj1oeRWlNI+
mbWulMUpL+sMsDE6Vz8DA7KxcIi8HuLlH91kVfOSbWQvWlXMjvJsV2Sp4L2tewDe
G0/uPENMavZk5GIzJcvl8U5GXLeztPJ76inHDH6rcPC+CigiykguSC0OA7VhOGaB
cjp+V4yXlsEW58H8EQVAowpmXaS6dzhvr0qBXlYdXoeNxwOwybdGqVS2pLHXsid2
GXif9ZRsdtoyOE05S21REApFMocqmQMmGZ0c/T/yIRDY0ciwXymy3WhQjZ/0Zj/K
vUumopzBlUXMZvJn6odGCqr7hF10Nf0aY99eZt7tKIn4/vBT9oLJ3cZmMQQdzRI1
/sGD7EiVe7+x46CoHop9qYnbE7SgkBIqGNOcHgIMdBaaCYyKxCXNuA1ccr20iLuF
sbtM6hfzE0qLhUAsMXQWd1MsXNUrltys/ytRC4TP4PqwgY5hf3mg+/+cgzMEMOM8
bxB8zfrUSrtA/d1sSeE1MiBIkpDyVueva0mLqR3ophQp9JKYm5fmeplxpm9KOPLP
1Fg+ltMwqBdxJ1MWHDOupkaoYGgElILxPxTMnLT8r1Kyk+LvvoGAtfrvDHVPcq1/
IHuwTFvT+b0+dwVn+CAGj9KMOQ/jR94fEwBUcIET+MRkGqNNHOB+gdtd3w6hbZIs
RVjL8iSCwBTh2gTcnru4SAZR0pR3wH5hUoBiAwItFiLVGSE/A8ncwo4exgRsbyJd
k4lH5bBxQ3YGMjxS6eE++3yo2FQ44PZO4s+493+5EtjZsjGJwrGOq87JyJdOywqt
aUesPxEgycPYgg6xD4Fe/Pge+9WjCBdHKG3C3k121kcMrYU9y7qKW1lQLnZ6W0X+
fFSLpCb4uTbTuWCZ7AqOIBf9Mu/lqew41sPoKQmUJVQJa0aMHdtPXJ9ti8NQEMBn
Gi/DEjP7jU/qiCeikE4rcpIgu6LS5vWGOQq3LPhjWiMkhqQmmujT56YBuDhzxr14
r+6H6LglIBMAqrl+zjicroEQ+PBrXfCbUqG+V8EK+7tNW6Aal5RdA8EAJIOeLuSL
pekT+2S2kY58pxsTV6VBVqKe9LGYxMN8EhtZJUidh/1HRDI6q/SvFOy2IaN78lAL
3utVIqlxt3ipjRDov1zD05V30SimVgSkuSetq0u2Yl9ET4f4O44KFVN8dbG6uIbl
8LRSx6HEppPMHd/r8NXjgozKcjDEx2pXbBjYx5S/ajyV25emL0ahW5mTBApvkPhv
aqRqBSRe/ESDMciSGQtxZAAGL2Rs2CHfO3ljJF8f5EqYBRbeuc1jMcudX7UHVPxs
8bBPN9n5erqdXB+DoPlCm9T7zagznXdr0fkjdbS31JIBy3FXr/G6e2nrn6E3o3TH
+EMGCCkAmkSz6IwvyXDCVVnm+ep9MChQ0G0U67ESWNqdzVpw9qRkUTu5Lm3fxKAj
f5n56IsoZ48+Tyk8MMNP0CUth/GlGvkAf3OANF+UgNaQ38Jc2yM4PcPNsgKKMyl1
vJ4dYbuiUICb7gBlbSG3ptT5I+Knt7zBCHJfbfiWJdmnUYmEuJW0Uh6q4s3UEx5y
Mdk2+VvfaoWl5MtP5mg+PKOV6lEnImRXcApgZSLBEBOKVr0Hs6qUTvGuB9I6Yyiz
vx+lvzcYn3V7/nkfC3MhuHC4Q8t9UGFUC7gTBnF1gE87mQa59MGm0nqL/7/Kd+IV
zFtlqZXKM9K5pAtYeXy/izKaiC8zp45Rj3NWuTVsYOAYexMwBIWjyRXlLjP+0Lxj
Sx5jbvyVN9rLnMGRQEEpZVlwK6MU8BngKKQgikILi0Ss+Detv3vit2U5c738SeDc
BbD7XpgU5Cm1rIfGugPnQioNDWarm+k3pdfGDX+cG8CMaaUbTgOMBPCzbtMQsB/X
aaunHFB+xryjFjyH/r+mihHKIr6o6ieVgYiM486uYcuIdGX2WOq+o/P/5Or8kBM3
1OTum4qcXT1pAH424rBGaW0Wf123NtzIzRKTOPLTPo+gIMUwv5r3nUzi8RuT+FKO
j0J0MiRXAj85nx2eKOD2tHc+IHt4JcmI5g321u+fw0QbkQcd6j5kyhusGwnBvLen
g+18aOLYJFg/Rd2Upf6ygfc5tMxOySD5Znz65qZR70Hs5b/nZoMKSpXwWgenImUr
185c1IjVlpvHszANmkAjFcVt4MNEpry0YUm7SAPqqdF5OngdyWHtc0ezshmC0wXK
WXt2bAhVUa/ze3Vf2FaSRN86CLiE3pb0BQDATqATkIZuYqHo71VmdlBdmqeQED3p
ibAmE9n1p1+NcOfzEOAfYx+CZMfXjfaW05Ji+sf06eze9QRBtfcOk2xxgdo8bvUb
czGsrE6qSWtKXBWGWqAFCJ9J/npAVViLZXy8pvmij3ldojxKKiRd54YJTrtTV6dR
t1cIQDsS515lN7U+5Bj6hVIphe184oY+AOfwy7fOw0oFB7y6q7r8j08tunmZlMt5
YCCyszAxbdar2lCG90Q9yXkrdRjiWI8C+KgOJFia+AL4STQiePI44m5HjLYEOIli
/hliF/GTJdz8ALGOr+IEy563ND0ZOLeT9vAlQ+fV/leWzs2LAOA3MElw1eu244qP
eRqNxlB6THYX2fcBySSsDcz4BHTgYqZRFGhgXZ5g1l6mZ4ajQG/A1ohuPVGUGE3a
Z130Ekl0rfoSxl25HElJHOfpTGu+EHTpq61VrX686jIMqgO17g5kny8YVszRnAU6
8Y5uyAsDsLI9CQplOHIMWbXLBkJby1s8+N3jmqKyEPwIEl7LgND/UQihRE0gWZO9
WU5/J3SgPtqogCZJJgz8MvxMgpK7q71W8t96qq7xsEPn14lGUEOlJjBMjGPE01A0
wwq4d4wBQwM18X5ZYmKHnO1f3HGmC5TW5NxZ0KuQIG8m4PoTHre1NY0hzj6hHwyV
9VK+iM3v0lswiqN/zeqPQlKxHXz8RYeVJ5DlDHS7rYGZMVTWDjryhfOzncIEkTNU
NfX5cj+4oy+NGga0hoLw9Mm5nG82gJFbdi1rJFDfftCXhhJ0HFYODr8S00rFKvrT
JfgbNnXX42kJTSA9eEfZGU8JEn4BxckYkYJVG3zfUK1MDPUsOqfnX/TjIoc82RFC
gGqE/uHHxwNFZA+g2dBpJUq6/aYeoQZJCfV+Y+VrvjFygMzPjVu8iP0PWggYH4Fq
nWHwpSB8+/sMm5zIJLu3znpbdJvMwwVh9t8l7grjChFFX/gYk3OsmSeZrgK8mEty
K6+Y2tB7Pcps757rKxcmV0mGEhn8mN1AB58oO9SH9wokRaVpKK+oks++GpJzemr4
gv50T2RP5QSDaR1SmIjYQvPEwPjaTSRltg60+4CJGbgmW0eqS1ueYPIpxorDg16p
gYhTVS3R++Gi2VeBSWV++DD6y0J2vbcAz3YvRoZQDA6iGHNztKEZLI69KIc4wFZm
ZIKcENgOvtzy2Ajk6cQ8VEnxnPxMzKtSN0zXyDXbdyCZfcfy6GtoJgUunxlEQml4
BxDG16Iqp52OXtsMZrdRKNnTlAJRFKt/eVG1GvFO9DeYNly4Scesx4aIbQRabHE4
kDS+x72nh5b6U/orl5BnPnNc0CP7NYFPOlYgWEIb0cpeL93MhKQN4QgGgHUNXhEv
RnDsFEx3dthq17rHx5b7NYdTmjFLyBbAwu9en4tSR2JfnyQvWpWGEKhyWQJ5QHGb
XiUkYjjB4YfrxlmFcW1mXcwxEdUAfZRfsjfoNs87/8d2XQNo9t1FBZseOHCkePax
lKugnlaMO7xCisyNxcPuX5mswgd/I7sZyE2ixUcjRPJ7l3apbf1X2LoGo1duo/SY
zl9M4u88hxfdykrt+8LHk3+OKB/OVO330T+zbicDPR8JUloJlbWsirgFmFum+Xss
5XDeTirgRq5n4FpOypAzR+xl59F13snqX9Qw7MLTVgbDAGvLs6raRr4Mxygzq1Cb
9pMnnmaKveUavsYYkG4Vl9XMlY0JXmjkBNXwig6NFhA4SuAXvEqJuvM2RUcqEpW6
mgFkixjCCuk1J88l3nDEuSVZLsiaQvkt291UjnvKF71TWZZmKS5GBHykZaNn6kXk
IAJhWm8zIPbg2cxC88lTOnx0rHqI1XHp9OZq//7Aje5Klt4HEUzUK18ESdsvxmth
btEEH8neIA+2Otu3hS8/3Tps4uOaE4zHp40YmvjWGvmjnNlSH1oi15+pguF+hg1P
+vNNs33ZMDMaedEZo0o9ZY4NgH9iGuUEMT17s8OPt0Djr1L8dvre6cA01UsOL8/J
hkfmQIfjQ1nSHwajFcdkkZlWO+KkqzGVnoRGRmpU9OriOiEiOX2/eryywHT1IYCV
zaCrEleMp2LxuBfc+WCyx8S9GgXhmNiTWC1zB9zDsLb2mnHZN71uK9mnlhIBUb0p
3peQx5NaNZu6A2SW+D2ojCNR5ogmrH8H/8oNG8QA/WgD2OIG+zsUoJEJ2bnWu2JC
kQ5fcQnCQ6++58xRM/MnQhz8zBGFYZOaMEaBecNQawa/Q5Az/3ieWzIqkD+S6d95
vq6oBiVlJo6tH4sfnELC5A0zGZsvMBaolGerox4s59ALRtjB4G6sUHULWCOZgCDw
6kp/tl9x3+IGL8vcLiI5198hY6hseRUYwk74TCSimAlzqnWUhH2bODJRF9FYmwng
Y/BhX5J1qpSlw29R67uweaKvJLoykzVh1oo71SxlnA1bgtI5dkqsnX2Q1+BU2zbb
kkxhd7aV+L/p7d6iGdzLjrc/CdxZ3ZS+GAyJ4yjoyTiM5fVK5lRiX4ksqnxxU5v6
98u/MzoC7fOptx/O/Lq7XFrmgLVZER8qOQG00w5NGUKakoL9/h34SbHUK50a9rcs
0V+8/x7c/VfwEgk/hkE8FcziGhw8vYzOtDsFwTmZsPB8F+gMBIml6GIiHZfrKDJq
PJ7W2ydPI7YDtF42rZ9Ygzxp92+Sey8Q0VVkYdoI81tTA/s+pwTzmjG3s/s996y+
SHqsYeRtrUDVyx8Fde4cm6PBQYXMwXmC5wMynFZQyPtC/Uc+l+qiHhyjGsfphE02
h9q7EMV0Eqwk0muNpIEqrP6/mto1bK3V4FNJfKA9q6cYiwVDv1GfcdsOXqaV3lAJ
H7XRa3NbZ07P8+D4D0zSKO1efyIhitSlqrxo4f0wyQF7ARgkb13SliDuf/1pSKPZ
+/lFsJ1FoM5VT3iIsZudah8zjKm3uQNvgAgvejrcOEjt3f1xHeZN1R3WePubn9XE
B0SL2JaiEJj1xq8KsE/B/XALJvivdHinUNyc5mf9JSi3TwTk3d9dhIUO5iFMFRd/
28cfeYXy/OX0RJ0an4vqxJ4KPoaC6qHcA9DB60yY30OJAYQtRaUJU6M/VLJrypvk
ojIlm8tjq/9He4Mmq29zvH5bD+XtAnYTKP0tk3Hd9jQsky7OhEjE1NAQa2aQTZta
TlMy6t1NT+Mgb/PCU3KsK5U55IY3A3Wrge4BOXMeBcsYSMWKSJlnSPMd6PfPaXOZ
WC5Kxd/Wibj7GufW2yAbFr0DijVR0k8tnakHoOvcdVZXZfJzbTCTpo7u6nEOxQcw
QeIu3vy0FEHJY1+/gjh6nP2wjT5U5VC4E8aa8FNVLLZTP0GLdX8rI+qXBECuF+Mq
h7zZMZkONYUET8VdYaydkVgbKImpb5mNNyid0Gw1584phlMxbXYlGHI7oOYOcDXj
0+miiL/ikjdaNBlY1uVqAYwzC8PCNpEvaNKMjxlNZpq9/YxbEmRBHAX0cmzjKZXG
0VxaY4dHhr66e5KiRVIimkPIGYmpgpSiVluvWqGe54B+wstjyH5fezLNPaXomwc0
a+4yWkjvrQKfRf/+AU12FrbFxAXEUZQ4GkGc4dO+m2rKZia8ljv3FpPqSD7/dMvV
Pxv/Y+L2SQ4BtVdrfjQ8Kbs9Ti8iztiLLrrpw3cVhg1yDCV+oOpmAJxbgXUkYGPO
y/zFjW8EpPkS8Kou4Q8roijHzGCgL4Mj09J+baHLoBgSKuAIJ5yf8DT9uioJJD/O
OthEThidHETAqBcoTSO522f3kOf5DKrunetNFyn23CkqwZVJOnE3DNfgrhGqiShC
AVQrj1tvbInWP/GkwnUdFTn+SX4zl6S+O3cY2lvGX8LKn6vfbCv1Thzew6eVpThL
v4fm+Ow/v2GRxHKoAmeESvbEK/g7CedKPwezx3FkN7X3AMS+XvhN1ub3rWorowa4
FYtL9v9+ORa3vulEIj6NhLTxbWAaZVj1V7iuHGWH8Tyodvzc66rIcYiGzai8YXNC
zWpQ3P6d9m9rnwMYQdWq8X44MbVjDqHLMuWZsZaEOirrIjVL/J/plzvaIgMQ4X3Q
Su+4sRhjdSCnq7jCnxMb+LzAZNSpP+nUkAf9yUYsSFKaUyNLL+FODdq91WbiuJ9p
Uma/r0Bz3bE1jla3bSfnEgnCisOkB/Q6GyUpffsBUO+xoufvbTd1W0es1kW+bxS1
XwTkP9mkQc/47xeQRWIjEmCSygCMplWybme2RBaC9JL/Y9GJHBuEhMEvQS1BjMqo
lgIFFipoRgPYZflkG0D/mN7e1DV63Thdy1BGqasDc61wLbpCJxtdCf/RcPUbbiAI
Iuieih8LGxHPtizwVvGFQhBeGefkHOrSwGhKb1ILYOaSS7T8hx00cuBATUUHgq7Y
Se9Jmx3sYwr08UXS/fPjd2iSSMC2ImunTyX4qzxNzthKfIEFtqQIzm7PTYW/PCeb
4s7VW7er7uNF17Wdxf5VA1Y98iL9tSWlLwqHtkUfaKDSB+onIu1XQ6xvu4X31cHe
RtfcqaitrQ4Txkr0hg70tXhqHp65+s6t9N2ZijSXz+lNJJcaP+m4KFj6On/JxNoD
WPmxlFtY8+6uZXQw9Hi08EX6Bg2AY4aCxSCMO667TcM98zGXs1sXXC32dkpLGyir
AhiM7g7xvNn3QkRkBR18hKCABfT3np3WYnnNFQUnU9l+yZM3eluyhesS4mEtREeX
trdF73Qhe76tXogn5MwvF+zYm4qVvPqbpicIA48mCy+EeZb/WDOkSlojFD00OVzM
fOpSmTecG5GGtkuP0u/kwiaZHiu6UcU9pRJoD4Oj8OJHEw7qdyMIH4Ugc9JEbyJY
xUgaW57ngqrzKmvMIg5ISkh31w2Tal1LDDF6UNK/KRv2nyjS0kHfM1VX30Q2Se2d
4NPf5NpjXU3zOP8Q6ofeOuQO1GZDMBAzonsaHshklME0Dmqi6497rZjME69jfa8G
x74j0zlJWkH7s7qgrzn9C4xeQEX1yGsGo3sidE3JiGQ12khQ7P74o8gLJCqAvnUw
7vVVgKD/Fg2ogXEdJP984aBwcFSTWSHBQn0IwOCKhlGqix8RSURch2P+6VIT0jhT
Q/Y9ZaWceTWLDIFBW6k3ic45bEYGiPPg7Kwzn2tqIxl5rVOckAwkMU9ZIwFhlkgJ
iVc6Vl0s0brUmPpuiPdqWoLRwCMychs4w/INUCN13/lgteUO3ulID1FAg7Q4rq50
kCcCtu/sKCTQKXgYv0+RO7jyf2AoHcCr1ZTu3J9KJqWdEcdTu/fg3vZcxk6I0xZf
taeMMkdi4TEfmCrkFyx8XZrRkyX5kG72TnScrtjz1NDBU7BsUxl1H3G7NPLmsGL7
oMA2ChtyGGNSVwUQzxlUHnhcpx718QG5qe0Gvu9PCLvrdyleGPykI6Oe0uWgfujz
4lgu4bVZixJjuYhV4seMLXwSVwwoXyH64GhaKAbKv52jCfVObyFLjqanvbqZDVFz
Evx9b9Zz8zKYdCZMP6D7DsoPxQ5owm1hb4YD0oONulUkW4gEgI1xi3vv+67IoCeq
yukz1fjobwfQbyt91W40s+x3iRI3reTGsk3YcQVysJNtNn310B7U/uqtant7QnA7
w4JvUe23DTEYTrf1OWdxaJEOB0TcuFAMUwju/BBdQWI8qwgE1iToUhV8NwGmrdzk
MK5/9wqXZN2o1AIbyUmujKVczFauki8d/GvUExoJzvnXeps/O0a6JW6c+kk1sxjo
Rv8jVSa17VLQi5g6ud7wukdor9aLpOwP2lB+PpuhBepbE9aHatPZP2z7kIMysK6q
vzX87ivPVJRrm/FWkTc6QRBDOMLUUgwLFYfg/5LB85h1tuBCtoXGjdB6qgxnKIPp
u+X01TgrUQrhs+B4iz9ZxaancM6fvIXPACFI8lHtjIul9lkhq9ScwEUDGhGYKR66
0dbf9msa4nbTND6mwFwZPahKdvBAEO70BgzT5uauUWgDqIoaq6UAfuHikQJUYlZt
QqYCwaF1VtB9LU27MtiFTH8JtPJ++pcbxfxjdrgEuxN6sbJ+B36FiBRL/B3sGBY1
v93BwOqPq3+O4QCd6OUb3qm0OBy+qNJnoGuNoBhcRAOpdxjjxhJ6NoI17F+hsmnZ
Feeh3gRVYjudz7e4ut0d83/q9XvZKIodsAaDAmM9Iafa96Hm/pvzoTmZ3B3cDEL6
GuKwiUJU0qTOUYIEdU3p76O/BSDQcUol7lQdMYpE4krLVgEKTc0/hufYA5h/S+DC
ClrxlH0Hc0h3UQMuW6b0hHf7t6HD5wJ5KiLVFpkGaGu39J3iqEo9UwHUaJYk3uLX
XYLg3xZ1Bt+fVALtE4NxGETe2GDskt+p9diVznRXuUTUac8UFFdONfUW5yeErxs3
RfNRw/pK5k3R3/iKZn/AC2Ljc+y4MFNne6HWouBcN4vad7CTEkkPAqNZGrXmSL6O
/5cQReDU4GhX5kxRTiwCHmFRMzwHd73gseNxzmhrEnx9mbtzUhU6vSwhv7Hq750W
/DZ4P9LQE8XS4M/RG+FcK7rLrTL/YIWG42phJpdk9Vvr7AOhD6ifKROxsfe6K6/r
8crXQAZYXMSkazotYTohVvYGWeg81+20dbZpoTcvRxL+tRfJFOhKWHxF/yCtlBig
UQA9J53ojRLy0FGCmuedcBrb+7KmuoOoxNfIfjlCSDpkwSOU7uqVnyYiNHAhNfYV
d0pkq8MKhZuGMMH4+FmjFzQboc9qcYLLKZDAyMxyZy/TDRQkkD63tVhu3vZX4Uf3
hz8+MQziqzOg5PrbExiNCBrZJjH47Smro6EL2vITfBj22IkFWZ1J0eL0XM4Upxg/
fyC2ooTK5h4fV9oViXL0rxNU/GgZzm3da/pCwKCIfDs2cJd1o5QYkoZtuHoCDOlH
BMkbj5iXVyoVavtUgwYudDyfwIqehHI6achnHQpeBMtE0W24FRRiSejSBfZhdYl5
gKE8SNz5aJuP66cH8SX+A9N22Yc2i2I880KE2/TFmLvKPhWCMlvoae9QLVVhjhEi
ftE0unaiSoW2IsGpoDXT6G3hRbae6MlijR4IRNYxCb+Tz3zrc+EUciIUCZANPiVz
s9UAdLkwG+0rLQz/wgxk4pbPshOiDP8a3CtiWkei337buoqw89KR0pnNnrkNIr6Q
b0yPhDKcdkKlEB4EEWwyNxxf2yuLNVTy0xlH4ZBxcHDtH1V8aqn31+huvxklQQ4C
5j91DKEvbOyWhAKnlMCevHixti9+WTVKQhNKm+Spjq7u08LmBXFXoK5YHehtv8fG
OmHzYoX4gBmTuGoQW0DaPf2Cbg0y5ARymC43GbM5RIOmXqEhHCa4/eShtvxEpjq9
ncWzxEmNRe/stL4OSe+UX9LSJZRxLhYcr3JA1FVZAnbY0ZktdrqNbnH5OwuljjHp
gJe49c3n5C8QqGD2dI/RMAXdn8Prt6pBlI0VgE8QoNEpuEiwzmCJoj/N2wme1Eq0
0AGfvsc2lH95dXpyQVKpJDf3sTuMwNaFu7j4QmSOK4QRgvfSXm+DBxLbhu6hpGeM
HhWtpOaYWr75oRBmMP6BDg1JXl2WxbaTS/XDhktGGaAGHRl/yJg0Ti0hUJbZvvjk
NFFV2RsXmte846fRcZPeCf/3K3XaZ/F9tXGZcQp4qD6yHOQXNlhaeGXRViplmcxv
au6mOnrz6ujYzp6tHz1LaY+Ys4tUR0q08NvFDV4/6pRrdCwOJ1B0MKnkXsdWvK1w
XPcqSV2QI6KtLuhb2Q4NCLxZznewpb4IFX19onozYA/KZnRNFUpDzcClwGBfvwzI
vSyI+NUJjyItmPuCysqSXas3doIuMJHw+3iZkXCMlqq+lTY9rhnEhtbmO/1kn3vW
NAbb7aE7g+BIj7Goi8yYrAc+GWUPJghYTW95ycjcGcdKmi7na9ndWnIFucNkC35o
cybZrDKz6cH883koaBwJA3AprwL5PRX4l4K0sz9Ev6tvAQanP0SSViPPAVBwJMfa
laIipCWL39EsziQy9c8G0dlQSHwwuEmjsyZifGh2RRhbxMd9CgMtSvfiEk58cK16
rNwuNxnLCl5ss9uTICUe3d2sw0sRzGo+gkoJ/UtKWaGkZc4653qSWnkUWebvn7p5
ea+ACHjHaji9UxudheaCkfxmLcBylgu/cPneM30xS8B8HtSZt0yukSt016E9R+z9
STKqeAbRKCdM1/oogLNlK2Lx0FsaAXttNgtuJp993K4scKtTxumxMQ3/aVFkSsfi
OVaGwuWxAuoKL1mlCj7ps/mlmq/vvj25v41eM63kHYf9KuqjCSrOHfkMfr+tpT0T
n3Oj0T9e06oWCPsCRmvZE8NTUkETR3ULNIG3rItqIWqaJS9efDMMvtUdBGH1bVnF
ZFiFMup8U9EhyADQQXZlPMHexFfd2icEthy8WeWokUWuUoeVJu6gLmTg47cwtLIU
EPVPT0prZioGC62YdHNoO9xvkNsBWYv+5iwHH9MrcpPa0O1go7nLeSe370yLVZWG
AYzzvHtKMXgKc7njqqe1sx9ncJA1eQQL29K4Wx74pr1S9oJbCuV9WQXHSJaOAgyy
kOkcJrWsLGUrVW1IVDPJnhixw/R2JyiKIntmsEzWBtO6GqLmPBQKnYylczLvYcky
+8tW6s+tDCgzUwH7aYgIZNGZnym6DyZkCaffh5om0nYp1h6I+gvOOBLH5smdmZsJ
YqB/xteV/izRnr0DmM0uTX3O+Teu4ly3XiJsW3G9Notp+G1ycEK5Ahlywcx7oqwi
Cm4vqQ6eIedONuqgD82cFJsP3Y1NhuVCH0MgdnafiQ1FY1VJOh/mt60qeVE96j3P
pMDmRApFOf9qT5ley/5faEwZwdXmlpo6Q30hAAy+QuJE864E4+xS1ZHgSBcpOFBA
8nKAcEyyVjY8wIGcXoW2Ug8IJaG7y3tkIishIwkKkfmx6LYSDCK2TYtrr59vaPMU
2MdyP+62FonEepD8IYfTmICa7SdPylwuZPot5WLMFkIWE7SjdLoMl60iv9Li3NM5
OnW/lP+ZTSqBXrV8KshAXXIT8vrWnHsL2rnWz15vBv5onCwlcDyC32EkQym84hdM
dJORJ4A+zTBonyhmucEdjrvrix55O0cq/der5i77E4yxlGGwE5nXH1IF75XXw2kt
fr2p7FRR/7R0d1iIUjcFkQs89L/jVqH6NYkC5lZgkbcCZc4xCeV6lFbfFeBsNfDq
tt2KxMI2NEt3wCsuC0Nvl91tQs+fY94dh+rG6FzotB/RFnIqJwYi02AiPhI8fJhp
3Hzwj7ResEV0d81rcOoUMoTUFxPso6DuObhx/cPAYgrBYNYDlJXb8t6e1uIaY8de
B9Vz6K6X58fHn0NGPJtKf0JijTd2QsXneQ1qWxthzY7UMxPvsswwpFw2AtygkGm5
d5TLgc5vzz59QKYiryYmRKhRoK9Mach2LnTbS+Gpqt+X0dMgrSY2/hzm4fYXxniX
t3dZVsPvszBzLaWWDl90E3Vm2O0Zuhl3RzEasDU/ve6FHHx7VEOn9KuwaFejJJwF
GsfOb2MH9bidZaOQ4opyuMab4xLHfRIujYyGCnE+7seiNIsXgYi82xFapMPCKUgn
jvLAbGBbXCae/tAD8S+sRRKLPMzLVRdi7cByDt1gPFoWjHUnPd9B5scr/wistJBK
XvKz46WZLHz54CVbgFY1hgJRm5u0YcYZzPjneufEgCoCBxqQax8a4z7982PZZyk7
WJRb6gdJDHgWTpNuackABztGTMPDNW7PI3Br90iuD6KEK/GjDQNpwpMBrkkx8UKL
zGEaDN0nF4F9EtsRlu5LYHN8CMAsW4IvUeLoeFCi9E5Bzi8oMI0uIBlJNQ0pMzDO
JeshzoR1yvTeocIgIEYQ4jK7e27WgID3rbHxpo5XUzLm9D4xk0edwqhuXv5V/XRt
dnsC6B43r2YeZM4RvkTdtgi1tzidJXudkAjv3ARBlObMMGIIgweVPXOF/HY2bKTw
23gSe3+UAxv6OdxD463Iewf6CMn21LS4vSfpEf2galYc0cnJgqvSzPFF45TrgX9F
9cODnKn8GWM55uyVQbFfRfhokiDnZncq/Q42lEiMAfdtRoFa3RHpRldtYo39xPt9
HlkUdI+Br2Qu7EPwX5Zd5iOPTI1xKPA3Ymed7yWpf1S/c+hzmJ7v6/7EDCFqrBuh
fy/ZjOeQht2iqd2DMZ6nvNbqVSGJXF6XFtNY8YN5XrBxwQfyQs6WMIVTuiyeN9UA
LdJZay8xWQLKhSGuyMGU+xFV+vTgAoZT5H5iq6pAKxCmIhoDrrBFW1t7DP+2Dsjz
9yW6uuKUNYtrQ5NdI2iqFPzeZktVValbjpQjvWUKfWrqdOHlof2CyUs9Sgr0Mrl4
nGKy58XTQ2e4/fgMCUJr50Mmzb+TGp7N5PA5PzmZhbcEQGNM87oZiPUoILRKMRkN
aTJCUuU0JupXkINwp0cUUMJceM/3uSoxl6YNsa89wZ2UZXP49Bz5Cc+P9Olz7OBL
nlJPqdnDD2oeEuO0XlVo29oDB50hjkSa7HRSVjb4Q0uL9iN1xt7j5hD9jm0KPLLZ
a3dvR90D5d/cDUbxPLl0BHM7RvzRRMRJvIj0A6SjKWJI7nwhoPZhebCsC9rxK0pL
UkBI6S9nii3Mixf587jCQYm49f/40krC8YdQFFkS+ft81nC/7w4ZTxFE2/Te3Xoo
I8/sLqnqOZrX+e9JNQ7OIdTgFkrbZRvOQiVHMHeKfRQIEUzY2Iu8m10OZGnR6Sm1
ZI9gdZaPZ5pwX53gi+p0EGnJ+m9+Xz1jkFs3ngIJVOvXDlBmxftR7gpQ/b6QjiKA
xKwZ0uMlB9NWhya2HVx97EuIeRBrPQXzJ75T4a3uDjdnjvVZ+5c+XAxVaVdn5eMp
dW0TmEcRNG00bA43qlRSzJkgtWDrgQNuD0vHNZ+YlKm3++6elEUnnqLHvCNMIRXl
WY6+lCigxauBxtL6sqCa1yzfpDwQH+Xmbyk8gFFArsbONKUUZjXLW1anywPBxDLg
wXS2T/2RG0Ni64iUy0kfdYn8ejN/dJWUdVIaYuTOy4F90yzvgh7BiNxkIOtgIucl
E0ayI4wI+EAD32RHrw5WVbU/6/y3gCkdGqkPI26tnMQnvvgBxWz64vln6xhEg+d6
3E9o3Fd++G+fMQvOT1ds5ippaFDGLtI8jUBVJEjpaOfOEO/ZStbmKrgpgxAjRh/A
aVFN9UNBn8GuqrB6dbWWnI7+UyWx9i9VA7F8PlzAR+Dn7llKsZXDWoLQ1H/cXt5+
UYuKaXHYT2OlrOqHiBRgdOU/zI39igK2BqWqlAhNRFj6Mm6eIPH/32ErCI54LmQs
G+pr8DGlIDHqZV36wdGZsVu9CsFPR3MtmP4HZluHmrS9EZY1LDlL1zLG+28U2vK6
5oaX30ThaLFVuD4Y9Z/HFS7XJp0vQIhbkZZbccSFpPR8QLZaQhvgLyUJRLxDWzOE
GXFTSfMeicELmpycn1v2nQTY2vH3+fNC8uqYWbNduqwzM2QwetDcY1C0gTepcVm6
FxoI7p5b4Lbj1tAzxbN59734vw75T0pIjWGCqoWD9KMn3uoIywl+neFnmH1l0WaD
N4i9CCKY+aiLArIMUgjMMqgoZj4Bo2xn9vgb1Z//9Qcd/DV29uH0CS/p7vSvae/y
ALpUCOq75fcaAiSCQh8oCEGesNnHpTEwe6+1BkSHhiHI+AK0HBSTUVK3Wx8tx9yM
pI7tNNjcqF/t+dQY1xKTy3GCD0GnKsr1CrRkxsnZeHSAvP2opVCULKAGwb0dfQeD
faYJZtMqRLDr3/TI3uTHMGy/BA7BgOB9+t/xiTkobFhYkF5jqjhS9DjLMmfVp56S
Pn+ZhYpTorETl4yVCZkFeUIMSpdPwA05GWNYIwGIMivRKt5HwV9OftOwwsw5VwSf
r8QeR/iL6H4+7BGVwo0zGh/BaELCvdfxyx0/J+SOkDaqm2tn9MMBsIMfl5DzEDoq
sC6iiWRQTUOqvT22BaPUEnPit86JMcFAzYLpG6vNB1xAojaWHQYIhx2Mv0NvETtr
wb5vxaIX0uqw943IZb0pPWKWrEySZq6LJlYRaaV4etilISY1UuSIZ9bGpshpb/yg
iCdeJ83m3yhoOYDDDT1rM8aShLOprX23giLtQ1bklC8BjqsO9SdBsrB492j1pY25
9kjbh6teHQwUQXRp3SnYoYEHvBaki6mNPKrh5BzgDWzh0XjVS+sokw6xebZqqf/d
NGL4SK/elazKwgwHNUvTpQZXOy8jZ594FnBgeTmNaQkpgi/YjlV3KOFCGAsUbDVc
9a2aPensfrWaC18dMqTb234+OOtXOzPsK8P7GfAQ2Vky/0KKEm2yxIKrE4pMJyWh
mf0iVzxR7rKm89hA79j9oYADHeL8PD4127CH6MJawzKkecV/Mipe69FX83fTIZvk
jsjLnn6PkzW/up/fVAU/HjSBjinvVGb2Hz332U8/zrxck5vb6d63zKe5INNSKGZW
gAA4U9t8SyR7Cxg0CwIwbcTNmUWsvnT1spGQP/vQ3UHwXPKkGfqAtsrJNziPa6hh
Cd2LUMw+E+BWsnXu2488uZsL/x8AEoG8CFENEN68YecTHzlQaqZLQ4bgMdOKUhtZ
aVneEotZUkgvaNhDx0/5UoeTwv/nfQvwZVaBoRkbvSSb//R6ASz4qWnSyvYlSY5C
nsG5pyQfyTWUiGtCTeDAOsbEW66q6t9T74eF5aSm4VveAIct3gsrANk5RNfF/Eg2
jBsCDz18Cs1oaeZi6kLkFfTaXA0RBeO1ykTev5z04C1D/ba9xFTa+TV0Obxmsw+q
zCzqshjvdquy7k3sBxuTw9XwjylWuO4ZCI3KlYs+eskUnpQuqNTowYdalCoTGLRN
g101Qge2V1F/ksvWvT/9BIiFgvMwQq7SGWlHj8/E8cWVFMO3pNMB9PkN3r9gQGMb
04cM/yjO5t6npF4248DHD8TuM6Kop+ltDwJIwpz7S6o9xp9GgallNT8LpyEtjv3C
XERTPj6koTt7ZIVhII/0x+jokrtLbWq4VZ6iYW1W7OG+PPIojvUmh4YNKvl8rbOo
+oAx/ZTvMdMeiDuWF3PC0vYJndWf2KUKki6AstlrueIAAbJBR/0tfOVbBR4wKVTy
8CMXooPk94g46ST7O1mlxkJ371DYdJ29c+eat5joW4tdWBJT/8LyqLY3f/4X0uFQ
mQxVmi6ck68cty/H+nrOs01C3RdXspUOAiF2psTq+mpDsyYSkP5bP9UBnMl0CDHu
49aN8czneO6WVE/HKPNubWnB4ofxx1nsAhXLdzFSxLzX2rJZagzdqrmdN8x0Q06P
6B5SFzQMulwFyyGNEoRYCR+sUHiAQ3rIwzI5F+fqrdZatoFXhORoFMjO6HpypnDG
cYa9snb6MdtxWLzQuYHuNrqV/kneStSuwPZ4Qp35k7sMqafmYUjP2FYabbl0W5ep
LRYg2PtYPr9Qw1rFgnPyTJ/odYd3qCcdlOWQcD0foqcvQDAlAcJVeXM1fSgymEg8
b1pIZhyyKoKTwSUAnI9avvJMjz9U/wQ9euMx1VJuCCKTu+G2nmHKNQTjz3jJnN7H
hsvagn7BjVkS8ikWPMiLC2/+jmZuoh9lq9RtWQugBquANLVMikiuq4l1o5Y78YTZ
rAb8RF5ya4eunmh2NgDwB7pTHJ+gj7vQDJt8trV+/cVZe9BzsIGHi7yFDlsEu6Rq
x28RJQ0KpToCg+KPdRJPgnqMrEn5+9c28ivtZ5Kwz/KsEp1+7xC4M7VUvRAgGT/9
oQA0zn9mIkzIm+kEchppao8j/P6kh0/Fe+RLRLA5MN5WnglT2fX+mJUkXNv6WTT8
MJrlGvni1tata/1hKuYv9/zQ+wSHerv2fEzYn5QfbScHe2LtuC3vVXlwZgXx8E4K
+W/vT7ovEQNHEpJhPMvXcn54OteykAP4sKHCsPUVE18VhaJYt1dZZQim+uTfTWjC
rolVWxe0QcgGi3vDhW330MkJyq4B/jfz4U8F8W9XuT1QU2mY3YDwtZXHY1sOuan0
m4qi5bocVLt/s1o9K3q8e2x6hd8aXnH2tFX48sKE1dlDgXpGnaHVA0zfpGGq6Ns2
TCoAOxgIm+SfaI79Ypgowt0WxYsMQ1X9rNB7lvJMZsgjSiap1oZJjQWLGiWKGYvz
o6oDHQ3CgXJAl7U3nSmKlVefKry1C33sOr7D/K9mKz+hzukOyNjItIJTrZAcXTUW
Mxy/5Ue96lLKRVegppk69/mSBgmdCRggrSIyDLV9+3WxAV9Hn+2BOtcxN0Aj+EYK
tZ/cygw+mPl0eDdYL/ISEKQvqWrE1Cp7SrqEKlRvEa1Cu7iQbVSmLci54srJggZA
/AJoKLQi3aeFFOqyZxwi6hrQQazqC+Az2rTU9CFrex9dJPkzVpVXBMOWwCi0j+MG
7RI52es8xhJ0ipgNB/U7NKwZFE10sMLHEalG5IQNPRwesLdKpLYphGNsAC7tiOd8
2futMvYRBYnRR8raZdc6HEK0HsdwJoP3IM6YSBXVgWMg/8kx6+b2om8OOfZLz1NU
btbzaiuHYh08uv/ZtIN/9B5uFMJ0mDCurOFoz1KelWeMevoEIaVxTqkN6KfK9QHF
mj/QMOQI4c21X8EEHReo6OSQ8SsUpU0Q1QBmL63qSF/irvGE8533JDL+tqD0PYnH
ParFAopz67du6v/YSoSe5ekGV/BQmEm6QwOko6EXCsS2fqB3IDtt6lgcXP9RkxXq
NiMgPpNyAWny5UmzkavYJfPWRGKv6dC5NhDbQ0uoxU6RBn8698OvsX2TRTDIe2bw
ejbCjLgt4nq0WTv6uW8h10nu6Thjx8Rd/4l+nhpFe+NFDeVwcKsD2v6D3bUoHm3C
o6oHwi3/MUXW+wJpS3SFN2Uz2FHHDxvrvt1n0x3lDUZFc9vo96fir/HUAtu8qCQT
2TXsvaZLnwCw6o+LmgFi+J1PF71ngDivlG8W0FrG8so+WnOjDBLAEh4K11e+QBB9
YaNtgEHxCLiVv0AsAjsQFGBfsDLDyDhJA5ykLSI79UhjelySNl505wYK4LLCHkUd
ZfPqmYbD/6dk8zKhmNhXd7SW8sPr/ON9atXdxldV5Edm+2hNTwdsEzh39an/atN1
XidEEndjI2J6ts9IPbp/41yqpuLPqe7uVzhniMhsaX22KbzvUQkbeY8LuKYknFe3
EJF688+4depVQHtVGV0Zo3E9RQzWB77qhBynh5H6adMPFXXznpEkthW1m0dn4TTd
92pQUqURTq+sZI8e2Rdk+YE+bqIQCbhcaLjLseWmmfzylv2IBJr4Rf2TMBmlOHfu
csM73MBBL98XRLowKwQkNik3jSNgilwaA+uDwUU/QEcLcto31uy6osg10mudn5hB
sBzWXTkMTW35F36BTSxSW2jmf3tW/9vrufMYwX/Y25/eYy8xLSTlYsQI1l4DaII6
LLLek68nWkI5r9jTTfv4kLp/vcwJ48oozEcWLipG8Yagj6oFxai/9PGN8dh1rACF
cire1p3oEV3H1FLQQkSVQWdTSNa8hkHom5b9Q6sXmWlRTLTboVJ9vKWvElOagHGX
LeKIGLtQBgyRoZm1Ir+bo4lsVJxhwEzF/KngbKnxRt0cdb15HWlIDCRlryMQWCkc
f4FhvSEMvPlbKvRYA/KeX1o+8eeZGwrVDEj/m4Y4cQhcnKHylScx5DDu6ctQbN0k
v+fm/QmpTf2kNFAFgcVJTbmiMBb1wO8JUt1HUiaIXBdwSDo7f20XP0PQrgsCjPrV
CbISvCUYir9uIO1Gt4N25sZlLM/dgGMmzHunN9pwHiFUeGeLobUh5aDqxks85tnN
gUQzg0FUk6prBCIIMlIbd4YCgui7OWeIeLT+9qXey2rj7l15io25up/6DSUGVke7
9SnXoIU0otiIKpoIhjFzXUw+s4c7V5UtXD5O/kJOPbP5KKBkRhvOSNsap9mvnoIM
qLbK96s+lsTrKEABHwm0Yo5Q8ThrwKKsIxZiWvgquLBfajmdFdjlb1UDllEjNrfq
Fsy/J8eJrTKnqlJkLDOu8NXHF50CMbMHqoslVZ4XM2uFfrynx0VZi0JdKqy6oQV3
PyxNuRXWY/L9hsKHElDHM7MFI7wUbHWdYOM+3+j5ovNyD9hTdboko3iiEY6qOFrx
oMuksmXJP1rpDdX2DIR7xoR7L7JDns45SD7uNjxL0+zcgelSCnGImqeRtelnIQ0j
58mDVpNXbuXjqsCMYPeRBGvycuXKsBhakL2MRsC0VMvqdOMxmYfyIqZoFJk41goa
dW8bFdOIJ/9+5UHJtelgKp5d8KGq7VT/XUqW3JY9yzNdPr6sF09aYY+6qqZnzjhM
iEat0lHYHHqk9bNhTOY9PjI1GvNeO2Ioh9Sj73m6VV72v28eaptiTUIqggBuR4RN
Xvo8Gq4aX/vQ5gflcRN9PZlwD3wvfQQ5CjdOAK1/PXfqQv/fTTvy3xuRf6NcBD9h
aIsmPxTr8tYF8kAK1IpqLXGeYsZUMRkHADpuRqYUfMJi1nA26o+MZwGuT5h6OjSy
Tbm3RIXF36YsqkroewLtqF4efBPdQR3mcj6Y1eyH0fY5IAuHFm9gUN/3H5itS2xh
Z0Iowlud6vws03qvj7XUWxlL72Uuch123XZqv4uGBHwwX8NYWuUOjZpJpkZVNyRK
QO/J9exqAqdGlZhTJ2W6TgthZORy1TyPAk9vOB9QvxBwJ/MGSlHvGTmvST0C1EFK
dEjfs+LeO0Jim+vrc+HBIGtwcBY2daMDOLwv1AU6v+E4YolPzVCHg3gyvWJX39ae
V7ty6KGXSPwyXhVQFC1N+pKSpp1fq4Cza9hjYSUcAE8s8YyFxS4FsHIfkVGcrlVm
eUtE6/vk3abWbpJcqxXGfOL8Dcq9AxKqdarfKkqMhCh9EAYJjGPRMMhXtaksQRVS
CK/mfi4Q8+UxnexKDqdU1TZQXZLtAEf+naXU/OeF0CNBqz4HSDSUPJItYbqrZ3vU
o5R5/eta9DsO3FA/l05VCVmKlpeeLjhy9BB1zkYc392rDNMl8wm6AXFW6Mi7PMFX
KRN9bFIUqoRo7sD4scKYFELeo99Ef2AXStJzU2Lw2rXk0n85Nr/qE0S2tSG5v9sy
dov5Y/yfuzdINXL0WAhvNfo4Ur2a1rC3DY53SnPYCzbYXV5lJ2av7hZuOjP2WgqW
xS3KZxrTClmA3Lp5UU1U8uoQsyfwfkfFM5HuewgF7WI1xWXwScE0qpKZSh64dJZZ
qVtq7RUYIM3irtPl72nxjp4/3pYcYoXAIZFMyZk+eoaIpGhezNp/2Hf3NMbmULxm
AH9DbWniXOLf1UhbW8S5DVG1fcCvoccJ7+VZeY3O6+LxpxD16tEfhjHg8EXCB/dT
tYdYqQ3DRkUvynCzQ2uYukSEXuo9kF7N3CtQZMxys+TEVFt8+8JboRlVLPmX2x6A
dOdr9foEcA2mZNYnrlwfjCWoD5AGaUQZ2sziXK5KCBy5PMCm9q4c//kwssblOce1
wbja5NLAIFLJ9kGrx6+Anz/FuSL4/2zdAeLGAkEBft31PofBj/3aa2tloi2xZUut
0g2ZYjx+Bm7QwVMJPzUw107mPU0m/4WDqWZ4V33rDuvuWr6O3TN5/NaCxhFi7Zi8
O95Hbli8SyYTQDoEf/ZIWEz3mfq2K3QnCEXKteDaKQUfRvA7t5zoFnjJiAdTL12y
++gohDVCrB5GkUCfvCA3FVUA6M8XJFPgoBBpu1Eo5pA1QX0eCXEsps+g8vf0aURw
rG1FiHEKZFff4Brk34iLpizbN3R1UG0mvfsdCYkTKchyKrYOeKzSLQ/9MKmOp297
b8FlDuvzXSa1QO5s/8Y0g+wHoqXmsWd6LeNw74Fjulx52hmqea1X+7cnSs7k1odV
MmV1uRKD7IBQaRMtfdfqC5FxQw8Fm9LrrB6N/nWEcedQ8EJ+WbJl4nTEv9FJEXsl
vuhQ+t24tYEEKZ7Lob7kY4yXmGIxsgSFI+U1CsmXv3uIzUyVYJYxt/6chgxfdI19
QRMxXHJxa7jv64+KAI5iZn/CUpV7UTQnZDDKbO/UqKjysnFtmkbZR6cU3DSwI/5Y
TdP2i1zLehUBj8GFxrvmACB6YxGQeCBZboExowSv6jVrnrUvpgcJ/6vHVQBv3Ir9
XKW23VYJAR13WHqVbgkaRs312Y8exVcyeUBfSCj5856BuycT+PX/R2vigkSyfK6U
SXKqHD2+z/fsYb9Ur8VH2BM9SxxMeFFIl04q7FdrSD+jntLDDQKEHO939qpXJtip
ac4J7+mKPVIzH3s9lusVr5psCegNXakGx/orKMzCMkXsHqPeg6Toh3lbqh/Cr+wn
1KzMqkNDikCDdi/2uLxCf17CGfNRbBcTjVVGzsVH9YR0jQZyjoQyCfbzmxjlz3Vj
/a4PMyKWJqmjAbI0+ZpiO0a2ivjPCukTrxL/imu2yWlR3Ym6kAs0vAyqt5nZ2WSd
t5ozCZ4/DJ7Lrno3qxwC/GeHzQdKXtKlVIR/z0Dd2wHdwmI01n9f9YCs77bWsoV3
QpEco91ijuHNWOqBRXbpD71yc/j3rxY2+8g8IzghUfT939KJjFQFGbk/ytr+TYP0
xLAPwDZJfxuSGf4Ty/vk4RLne7M2zFPOS0WQkIqHtQFcWGqcgvuTN1CceTVFwh7x
zzDa7auPUwwE6DBUWvt5nJhSDp9OPj+jeNwWac4ysv9iYc2j1X5TjmOFEMWUdZSS
gFXJ0/MhIh39ED6BWgQRhaY76fgtpHauIUqxDZcaSL7kxtAFOaQlbAQ7mLw5MU9e
dhcSoIX71RZmDfXdqs84VVrUCwCsCXcp1FHrJ7dPtGUVjdqndjhhcMIfZmQqjd4q
juYUTIKJJ5CTeYbP7fYKhUT6IH+qwRLjIjnWthlRmRmEnKgf1ApQgQOTufANSpWL
8d++OP9qohlrRcgg4gG9TWX/cK6lNcGO6V1C5XybwrL9+yu4rfpp2jULX7ymcXFR
KZp2CtZkZxPekDm3rWy4Q21lKdhSXQ6M4fUyqbPNAYlk6Hw/nPGIebvPFzhr5h41
KCODAe0qodF0qfVjUd0crhQYyFelNCYMq46zAH0wnNSaWn9D73/hnDs5WWc0SmXz
1dmAucxhC883EEbBFxFsTKOhKA7bGZo3WuT+XUsidKMUBm6FevpHCbZ5sjJQU+Kg
hsBCJC0rtNvVmGyTGpnGkHH0q2fBIlFUerilCLhI9r7zQ2yo8aJxa1xBW/vmvMA0
/gjrqzKH6weaR1NCgFngJo2ZjhQqlGgAh49JSBviLJk+ZIdL797c2Y9aWSCFBxlJ
9CKA0piSQ8BeSlTynmiBbkcfGeUy4fcaHVdBHhALYNaBEwe8L3wUh48B8wGtBG16
2s7gMX781Imv+RuU5ItWPOA+eTA86DmLsXxmoXtAL1MMqVMSeKd6sKaVqICdr/J6
QQZMsgXCSGdaFZNmhSgfKpmIKz/teMQD8YGbloQzm7tNyWcarppFWqKFn7/7Au3f
Zmn2/sqB6ASC+PBJRXtCWiMCyXUOyeghSyUzzayHUN5369XwQJGyGzZlhyGtdKI5
MHNp6SfaIiT1dOa/vHBmV+gSiZGVmIk6iCLwqquLiJpupdGScc5DovXlAej42wlW
2biP11ptr4u1XObIPqU86e2F8P3jLefE+UDs8Oxt8WgL7tdLyP5jiHJoS26Qk9bJ
os1gZNlHUseChM5Hfe1kF6f8sE0wzyJVpJkT/ALxVh8dZdXcEqlo5W/AkMB3DFXf
7CXBD8HEHk8u6rQJ/aKmy9Td+RbD4xjkyZkM5UYvgUWqdkLKJu+n64dJxkX1RNJo
4BVgfmRFEyaqXb/WxQG2gJLHyqbBkm7V2FSIed2bsGRHScVq/7UjOrh0LmnSR2Es
AlwHG2cl+MI1b6bO6SEWWarUMEDCQ4MpAA45rNQTvCM+uzmk5tZyTRt55oYAhUsO
kRsWSPqvORj5yPNAS6uykuVudBTut4rb6i97fc3k16MZXaig5RsYDdxiPa3E5BZ0
8k8QkqyfnyzRA3hcugVFwHoy5DKd0W4CvPFAlbFtMWH+31PUU/cv2NDT3+5PfZ2Y
y4uoyzONLMOZsDQl8tlymfRPZjumCrYimrgy4OeeoGHk5cjSKl3+oiMaT/forZAk
Huf0yWpSJG5ZnCkspj0kMU+jXpLBXH1XOxfN38D993ZfPkgbNdB1wwvwmQDR4LDB
PrE9VGA0kKpnGMAu29mfJHSWO8PnqYTbMaPT60FbXHAVvd0vjfQx8yaihZJZb3V4
vflRMHFZlN9k22CPkL+j2tplYXDTqnVnxwxrH65ZCtIJAgUyb+lMjPLLdRpquzKH
mVwCslxwUOEKI6CwgII49H2DB5nnIILVXYJqQ48mVlX1OxAKAI+dWsfWe7g3UTbs
1zGt7qkWCQncTbKoqQV3sN+X8fFuJk6EjwaV05sxonsvHhEtqK9X7GIA4wWXf8hg
kMqOVi4d0eYv0FxfW3Pim28n2t0T6aQzXQOu1oqEBja+7T/+HcWQ+EacAmGrdWQ5
8tOyH0zFpLHf6WWDCewNn/FRe81s9nPL/Dc/J8den105AJRmNRAZFJcI79a9lE/E
Xm7x/jjjFcZU4kaBF/AiSvDkeUK7y51ZsRFi3H8GIxJfOTv3KELJ33GcfceBXmq7
LkfyQlUauVZ5CAwAPHAK29nd4Vm7Pfsjo6KNic2F/k3LFzhY7cWxB5eU34pFfWWL
2ResBaaXLUrWU9j4wR04CbVWoEW+mBrtThf1DW4FfiQ8pXHD4dcIGe31STlp1+0B
+xRUxC2kMVGAAYvG+6cmH8tV/Nka+cUMq3VADTVJAVgpnj4SfY2vqGgTdfwqZPNT
vIPH+Qqe4lOb4ESnJ+7MyqYp7yq7s+AEZBJDroBU6DeQ4H7AIunv3I7nWaI4t9gt
LEW9KAkPSQHbRFvqSeqA8Om3drg+P58YdUaYOhJAQRl8yTICAOGHmA/Ij6E83ypT
Pzg9+jg1nl6VenQa6kaomf+rvWF6U7JDZWjBv8aDTcJB2wE4rH0SR8/7f7Cf0kOi
sidLg2UIwwXhiu0BUsLDW6MRwYpPhSYP+Y6ckpDdRsEPXeplmGes6NQGgR9qRnbd
RYOYV6PAJ/nwebecRsc56ACZua5r8HsLH9nZmgn5PVtcpStL3EpE19kewP2ybCQC
oIEbGhE9nELUVQ2ZHH0pIn7JbV5F+Y2f4wlgc8+o7odslNBmxjM+Bk514/n3Cf+K
Y50aWBWT1SPWZS+dGuoYb4I7o3k39Q1Z8soUky4DHko+er95afBZF/xnp0b3TsFw
RXDSSVnCFxtO9b89DbV9F3uOKhTajniAgY9AyNKBUPhExAjWXgXPID/7h14C/o9o
nRSb8XVQBkeJ56lsG/k+s2uG2ukqujuqOKxZ+caopsnnnEaDwH9mkkQ1jg1BvI0A
AeS4xgQ1KySjSOzTo0OfsPIUClkYWrVa6JCI8uKkuKJPwm/HgjApsecbX8jYvf6e
9Ni5zYd8J9e9SVS3T/ubbtI/8kCpK+Kvl5iKKKRIF/AN651O2VdwAULYXpw5FppT
M3sK4X7AfWv0rB0b9OQhlOQxWtfMqAuS2GHnGX9onJY6dG54pyC/d2feAeTTlsLh
VE/soBImssyRg2r0H417UvusLrOwTZoANE0gjni5c+714Wx+KWVj6nB4lP8gueDJ
7YC4NEWFemIELP74hU17BEE+SLTJHZ+xUxxJnqFL86pSw5lHmVINAUwbe9Pypeaa
QVUHCUUEMZNDag6gpCsbx1/lPSrqSc2r11qfoX2tgfSHiRs0/BRbeHm8GS738K2b
qDGvmZv18nuDJUmvYEVjALbNF0tGV2+4Hy0pzuYXZ6lOrxW8/NWi2OBXBuG5J6N5
o1obgJZpaHM9BOG2E7UAcRZ73AoT3KhikYRmSPWQceI8yn49qO3SJPzE3B5vfCFU
9MDIZkW4wgLoCQQ01KnGzSsuARfo8DlN//r1YBTGyZ7VHmd34EeCAEzgi77kCLBh
U/GLn08VLzVCIGEYdXHjs8uKJ/49i2+SocP/7+LcBWvL/Kjf9fzWjeW+76FCi/aW
0BTXr9o5WBGhLQ8i8PdPJric3Hj/CuCKAEI4wZq2hyxPh8bHCAHGvCc4CrkGDiGv
rX7HJ9sOBJ88Z7glrEm+xZxYNY3FfEoIf4szJ+M+XI56UsEqLoLgWD0RohsdXY2x
th5orXk8Bp3rfTfq0ONgqWyBbkRaVoynfC/N4CtR3S2h9RMly38s1O4u+CC0Hel2
IZlCQbVu5e7ySAG1ayY+wEce9Bjr9knPncgbi/nW9vpRFHGSIGz7tZZgPTkdsY8G
nXguiMPbSpTl6gmKY56qiDqhTyRU7PcR0uy3X1v5DTkDeThrcVMtCiXV5DqRUt+R
gqv5GaCRj/RfRfNiTs2BsGACIqMbgMFlNj+uBNQOV8XVxUJQxI7C2/9zBV3eCcmX
TccFZ09iTFCfmKMAgADZw/0IamsQbLNEtD33xFpLYzY1Wh/bDgCsbrl2QUsaAgwn
Zyi3yW3kAGo8ORKcgeGG1TABXO/AUm/6afaAcxzHLHKZgLPRRHf5b0rZocmvNXvu
U6f+OiWW6hnYGjGmNpN5wMQgGa8MxuCvURA/oKBKAdFnOuhirzFDLCxUGbN8hYjU
DML0Sn/4ah3/rvyCE3Ub/NdZ5u3yPNn9mZRNhY1tjaCRFKk+RYgOtEHSzPMbNLdP
R37MODBlvHLDrpugI32aSfnh20ZEKjNl/RYrTLHuR4+PlmcbLB6arDHMDQQzxwbj
b5ozQuZAmoerDCwSkDqffJY/NP0EpSeovSCyHD8aWaFyMjDM/H6TzMxiq1Fhl8jL
WClB62OgKQi3H2tPDoawnoPC6vItz7TOIvughjvvDjtgSHAk+N2PWJIMCWl+8lsm
/t8Py7YjvGOHx6LBoqbEimmHQK134Di8r34Cmoa5zNM9SAtWegZl/Z2X8AIs/Tmg
5KKpTmhPUHwXMDp528u6Er510YyGbLfhZHmZkZzRbTdI1hTdhddpiUGtjMJ9DBPS
INkVYxKTjasvbLAV2p5VZf+oZ1VhEBuA05lvfZAXplyQHmAeSviXGxxUHkZaG4gn
lwk/tGaQOpUgoz1mYOGG6DQIT2COtipSqzCaea58riS1clRm32lTSk3ODVWpSxbp
erGofE+QMeStkRpWqR5XQRPPUOrNkiZgh+QCUZHniNZneJEYKKRTbXVTouTFUi53
aGOI5B6fAYTadV3au6t54iRnkfk8ljfYdTwPuPZfD+yIjcNAsWcpSs+XqoD+I1eN
oQU59NH85IwEgekwhDNwuSyG6KwKG6vvvBbo3//3LS+lZ8KztXJfpVZeuEmdRyjk
utYsD/m+w3H3MctCA8+Kuoid0U8YUtTK8xuraWyTW+1c020oFV1MvYLMIJchoPqo
70gm3dsCnPI288n1o//FIcHE3m0Dyo93xF1P6I/RbLYywwtVivBFgaD2pRBGZgey
yr5gy0bUc+bapdjJolIqK+eQtPJ2xVPliCZS8nvWSm48vQPwh/eAT98KEtD2ibC/
fY2ShI9NMuN4Pt4C+iPWD8JPUz8IhpDg9+3eyxsvo+mP71cvRuSIWOBeyoHCHo/K
tmBuo5lMhLZQHZtTheX8PTTuPefWx2Jc0pdwiBr+8ZPYYraYH9k2tuZgWu2kOBP6
2V7eAyQxqSVNxcDZ0jafsKFGWxjdjdh/QahrZraXOIC2MWmvZJDuPNDIu51ijwDu
Qv3t0u69Yv4voj3vfb1MCT8TA1aToAfCwC7GGEM9+XyYedQzFOJ72fXo5wy4kega
GOLS1szuGFsIVd8rk7TZCvwP/KT+kaHbQApMXNQqE1qX9HB7Tug4bv3FEwEyl3ra
gIL0CLjwKa1PG1mwpEI9H0+ZPHyQv7wb07n/m43n3iotLfpLlK5YS4vA60tXq+o2
EZwDemmLU43yLNzmuRkRDkOQEqFw2t6Be8ebVrvALqCCOeXSrnjvu/O2lm13vycq
XM3WTVBe8cBfYiU5Ce7yg78x4BzCr/CEtXY/LaEYWHa5icpgMRY8oGEwvoh0hjAj
jF4sPDJaUVbNzv/q5psXYhwR/XFARlHx6zZRy8e7ypk5XjtGxrTJ/KgrNKuQDCnX
ttQVOJoM3Gtai4O2PYeks1J0GeQ0cLHK4KLvh1Th0VKk8ql1Qf3Ry++9MWEqFtH/
XtOanoQXpuztikGg7cPMcyS2tSZ5pdwoqd0EucMRHHO97wIFnTt1+HvLYKUEdTjT
7J+c+iI7JqqowFBnqPy673MgTIFUksGMZpINXyCZXyvU31bmKWqcw/+tsrBqmc/4
vppZTQ5CyfXpZqwXY8RyAkO84dqRwq5jlnQA9Ga0Q2y9LBlt1f6NN9oCwl4iYVJZ
5EXgp0HrvZ15OafXkPVQra6dLnUJXqjbZ3oG6Oyr2Ecc6cWjmo+Isn6wloNeNs1i
1v0ZU67oIvMVR0J8b78Z2PHoWpSftlQn4c+y/zv3xI3Y4eST9ChEVm4yExB2lK1u
eCWfY2SzcRsLclq52kWkJDmpVu/jfpEi2ipnh5aACuMlDLC/3jDXgqxQd4q8xX+q
VGernxeYmkPqMRQExMNniq4ouvb/ual4bMzkV5hL37nf6nhw9TV1uKnihFetdzxS
BpgzF3GydmynLd6e5c4d3H5IcDBQ1esP7thY77GDM2JuCOeqqwMcWD1iJYPlqQ5A
2TqAogUydGVACuuMPu8hc5yU4yN6moyQ95JX2+06IViY10zungVm1LF332VF91gO
fqNDRkywtL2Mzdtbvfgmdoyot0+DYDSXUsmmB27aFgt3KSDDeNe5NIHTUdIliKnm
FM5iuBa8mUDYWb3CeT/qt7rdG63w4mL67cwxc7NT7Ij9Kruo6NJAuePSTyGqbTDc
AEf6IaLIobvcFPFoLygfsZjB940pAtor859u4xHcprRpZQgPnqJRdroZqWaWpVmj
UdvbcadnJd5/1snK5PuESEmGtEUv+lKeiWX7hZ6gyHmWTRWcWDiC7MNyijNJ1h02
IHAze4pCESbWJE8EvEZOG7yGhdXI3xw31Q9VyGjROMWpIstFVLdcgcKBPCHCVvcZ
V5012OMXy7WesL6p43CPT+Y26e4lfxmuAzwTgngqigTxy7GkT7ITlvdUZ30JURjC
DYg1Ue8AGNtSPKtgj4LMOS519SR8eJO2DHTHY+9r90ii0mEabDzDMbdVMEMiCNqH
TU4iMltf6aI7BLFAxI/ZbpQ8ntL0OZCpNLU6z40k1P9aHKVzH9mnHGza6FW31SAM
AO5NK/uo6Zuh0eEs/aFM1e6OA+aIuqBPRAIIiAEJfMs/J6pAdLRjhkeSyyUJ30Op
EVb5nGG6ZDGuUQeatVTd6fzv8ch3jX/TaAxHHo9pGVXH7MjVgLL99qm+EJQtCLIV
vP54MPiRwwvNEV7kKuAHX8t0ZtCuIrZErGM8TFoZlosZQ/rLGiYxLYTgANhLivH0
/yN5GoaCFsmXhzak2wpSLk06aLcWrBWgaIWW3NWX5nTsXGNoYrqxGl0mbX339sLJ
kDLgS9gbiB11f+NekBzHZr1djS6PaEey2CwwNIX8HGtYPp2r7259a+agQfEbERpY
vYZ+usEGGCy8P/BBk7zK8P6BdGHOv9tKVWtPiOHfKK/xQcanzNQPtdlILH1+BsVP
TMc7ndOg2UnE6QgHOY1aEQ4fmSrz6Jyqaabh3mVHqsi67xYJjlPie98lAZ+vlBjv
Mxd17M+Jj5bd5rOr8mX8naiugeYAHGp1unhcMbRC1p0WEpzdiH/DJ9ijlWE/gmgp
1+9m+BS0TafYKvVkWYH433/pyTs5MS0MCQKd315Wr5IURhQDWapc9ZSibgg0JFxP
hqo01qtPpTXWHbanbvGm81787CIPpDcE/twpji1OsKgc/5epB5rV5xkOx21G70Rq
7uU66dqZt0j5HqxNgRl4HcylE8FdOJQFZE+EohmtATQ1jEgKNcxTOX4CGzJ9Nlip
/y1i76X5IQL5TiWz53nWlljZtNvCUstfdmlQ9ONlbA7WPxoCTvs58frGlPHLo5dv
c7CxJ8mIUZvldD6MV44ZFghdb49QDoKoyOu6+b1K5cpxa1JFdIBwEZS7bgxF1mON
NndDKPRBDxiXQwbkHFmcaqA3R+nnvna1EHtkzxyR88L0mBJ6AW8Gx4mli3OFibR9
W2hfpblhSA73kftdHPZegjD6OLsvQp2h+HZAnaiqAWDngZHSMTOBfn3Qlu06jR8X
8uIo2drqT24KpIwyNzHreQrtXtvz1PxJj6AqFlCwdXtbf7rjB3EFECNv2rZK4qiQ
N2w3V44owX0AA/X5FjV/CF7UgvHIQ1LDg5BC0z1UuJx8Ut06oWOk3SiL+zi0077L
Z22ms0Pf4aBwLO0W9IdBCdWalEK5tJDz00zLCeXh3c6hlo8TN5QRNVEPiRZNzlsc
W/chL+8V/CDtC3RWq57bhDNhjktWsZQe9n+ieB/urwyASTE9Vk/nFHxha3siOrwn
WCRM0tFBNbcZ1fTdG1ZEIfCpv/cY9hS2TujC1auimKZeiLLKbcF3jvG7w7ixFt6F
5/28bxFWVgwLAMMJEQ/qoNRLA00mNHPmxRIchomFEqQN4HZQwSA0oKqDfuwuI6Dz
AApUIdg33IRdow6pIOn/5gP9QPgM8qIb1ytXTjDnN46Eax3ssxqDT5elKM53Fp3j
G2/UVUcN1tjJ44uCmTiPXo5sIWhZGsRgoF/bNTNDxBSTjFMCFODlEyr9kXZ8MSS6
IkvQg8sBvYXQsT2J0Pv4rlSeg0KQMY9hg5c8DIEmFYNsugeYwFbhgsBOA7Yn/r4n
FmY3X1V5OQAdKZleqnrUo9nqdi5fr6Zk5JN+XfwbEDdfIE2W7yNTtDboM/Ca3VXs
0qNErBPuZoBHunSYUO6i4VYwcd8auuXvXGCSE6IOSs3nyATdysFWaU5jwJE5Bysk
VCAXxuUF+Sp5/Db8a5wDFh+D/uedAapU30qQyw0N8tPpV7ugyGZ/GrEzqWY9J6Uj
K78gs+RA/AYf8B/MDiMArrtZjBdpGun+LtZwxaTKZWLVMITwAi/kK5VJkNjZhEwj
D4vb3ogj9sbNAks6e0M2c+PaEJxJBHDE4yyNpoBMltpIVtXv05iCUa59kheTJvbI
U4ws86e4BM7ZbWAJ27m8HmzK94mk3TnSAfRPIGl5ZuRhKworkJjgun2qwQgoEB1g
eGEn09qTGuGRnwv7AwdxpSP9nWwNB352D7Xa8by+QF/MQUdWrrkfhWYqiNtgFinJ
Ay0NVY+2jw6SIjvVp6rhH8EumRGLZ4NWP1Yg5j0QscA8BWJvAb4iKpURCifBOZFr
L+RbOGWFkv+0DZ11vcyWXjjE8/uBHnCvRiwOkr0gYfyCC0tfnu73iUZhtLeKeZYl
/J1PJIkB/pw4c1a5s6LT/4dWC6z5LHCEDZxIRQY35nh3CSxTi/3jmKzVfbQqe6gZ
fR3MsfLeFjaUCVuTvNxxsya09wSejDPO5eaCYouN30kDkncm3PIKScX8Dr7/IYgq
jL3ikR1qfQ0EETcMk1I7WZHpQP1w88UEDNEoEHyiSebxnSF3gsv73OJsDrYXPu0J
ay81+46F+fSPKA26tKCMDWa0yoZ924gs8KG2zr3o6Ot2jR2CMewhFNCcbvMepjET
6y+b2tRXTPuy+xc2a2O9GRxnvSPUwWj2k/ULrlY3Q9bhLdcnndTvCf0lLR6WC39/
2Z9MD+pLbymzRsYORc9QCIi/KbVT5Uj0chnNlhVSeTSaxVJFxKhAZXqdtrNvGkn/
B9JXTnuURHBgHxsqS0oROIQSgauCf4HSFK2DU8NSv/seRpW0m6CoGaI3B90y9pbQ
m2TFb+vjeQ+WMXkb0TMLABkZBPV70Tx05at4y78ryk+AhxmExjDfkaDeDAgd9urs
FmwrTnICU6c5bKjIf8pkQvE4o9771kCoMRzPxn9NrFsldN+i/0ETmbPtsYa0PfQn
Kw3JtO8tV1jg1tpSzLxyUJ7FwZWRlaHS4WvFBZmhUVV5Ec6GXt8c+eAyYmc12pTp
L3BrZ7qatQVzFzy+cibLgf65ZDDxDR6SvFSVyoOwFugqwcmaLHNJo/kblGQVkbTT
UFGTiJWhOJd6nQtQG7xfFMGP0PO2PhjxJCZr4GsQq4X3ZAjZ/N+XpSKiOPXkGB4R
xEqJ0dYicYwk2ScZFxyfiBEp18b8Cex6cUQ0+JIrbI4RWUNvrJCz19jgTyGECty2
//oWEsFoXc16DlZi/2Jb+07yxpfUvU1iLfarZIIl0ZXn0OFpzIG/lw7NbrCR+lq3
bHIJSB4SQj05+RmGTeAGPFpSiPaueRPD2tR86Y+xoDE4xSV1NwiKSB6j+jhFFpzq
72Ovck1v9F+N/NGPEDm439YjK4RDjAMPLKCeNYkN/+ef4UuRK5hu4uW549PNM7/u
m5POrUzzG1zCjKW325/LLt1IhqE0qAqAToydpBAwMTjATPVGCxwZr4UNXE/7DSWb
kc7Bvvxu/DE1oYdtfIwrMbKxgJu2LG9PYzg2fQl2WP2GbRH7/Yu/fVyia1IwJKb7
9lJpI1zPt9JUVk0Ei3kDddiYqTklm0Uqft9oL0BATzS0tWZkxXDDiQt6RCx/C6Ug
oJQCzlcmiLzevGvuCeNgsuYAZ7L85bp/nkvKjKoXLHsV6TA15imenCOU8PiwJO1L
lL4t83a64peY7Z5ir5EGXOiBwaTZeYJow+auntWjPL/Ad7GEhYSd3iSnewJ96wzw
zMhazCWYFraL2hWRHH2zmkdVkujNnIBHUZO4pT3bnIxn4Vp8K1VAN1QhpkcbaAme
A3AXY+VQTTUiuZAXW43RQaxMVG1LLQF/petZFiwY7s9BRsWXQtQfUpUBDawT7zqs
wpwLjdvIqwsQ3vPsVE0fMUUh+6zmZkowRF/Qs+f8eA55nf0CBVSbh50AhOKVS+IS
t8jvaaiiagMHbOjk+K+hfynGxwZ6VtqQd+BpB3y5gntpPAFynRPf/x7BX1ZtHsqZ
8yQl1t0ZYaAwKLagvtjwLyLpoz6lh7k/W9dO2q04MTzmK+69PPz69JkdssGwegQl
HpSeFJiGfA485dlwwz4S4Uhd1iG5x2W6885+zi5fhxfskCCGi7nAFZF3YqfVkhgQ
HXVdd1vWUwiul2JydY4sITy2UhpEQY2JH0XMkafkSYSHVdVNmlUXt4S6e1halOzl
i72vAsFLwGXvCUV/z0bLBZ17YC9DduOrVuL2nwTUSMX7imG3EaSTeQf5AWxsGFTS
+8mBKGlSYWy2tWeBoHjhU1FwB8CUskQIhc2sqO+kAW65K6lYXybr3VZGY0SJ+88Y
/mEevhg7RApEHolVXrCTah5HP/L7SyeVU8jssYPiliHORGZPJ5d+DgzZHmvvQyRL
R4Ssq3u5c8AtEPwgQiJ0u2UixcftXSIEaTs+iBAbSY/0KlF12RUBimYC0GRVMBzs
f5B7eNiUj+YO/n0ZjYfDIqlHEt0AJMUdtjoBkoJof9eeSMg+gSheMU2WQtSicU5O
t4+X68DEbaik8xMJnGoeT5lq/vU4/8yZPk2nRm1Jgu5I/Fqu4Key/MMMPPTkeCfx
jlL7gJbiMGP5sNhC9zJ7yQRgtXD5JaA2keREGhVLB4MoZ4wJd++NTHD6ABNnXeL5
iR7f7NNIt7guQVacDwPyGCAlAHga/slVbOA7HxL6McQRh1JPzBe615/ygouf+iuU
Ph9+aTImLnpjg7PHGMK29NRjaqq8VzuOcxHB7RSPyx24TIqyG5l3Wol3VjElh43P
PPdSzQ+swDdVUTzwQM8Fn3R/5W6/WjZv713XX9k262hn9abF6EoVg8vBscy2+vGt
+M4sgfyHqNwxbSSWxIJdYbaFL9AfB2Xg52/3RsvfWNqfRgYpgeCtPJh4qtn0Xf0j
CH+iKiCzSPUI1hf3LuQdX5ioDzwnX/OclhpCeGu4fiYhljIP4DeUVmLrSMy+3+04
MCiRdA/aj0FR6PyDp2RGFMxY1v2PtNROWlztMqfsy5P0VVxYISWG3z4qcty4TH/e
tepWgaM+klC29NzJtmCve3XNZ6ZDMVyA2VgiQgi8DE4kNr3F+CrNgG62fxcvV/9Z
rfJyM6DPvHTl3Eyc1fXlPKVzTEb8HsVubXwY1AXc/PYi0dGIPpDQDE659N9ul+Se
CSUkAxxhBWqlcdh8zTz6u8/YjB0IXkpUBTfPqIyDOv931d2SRNahTPraRm+j8SEd
nC6GiVZfAFLfeF07DOsMqIHMqd4aNs4Lq/61NSSVFvwMemF2oKIGcazb8mCGwN7d
+QBL0YA7qzDzXQLauQsYd3tva7rRTYfyC+4VE4axTslzbLOs887/ZKqs5nT1HQ5r
H05NKy+/Evk9I4lYfkM0NBmjQPuD5JAvfllmNQ7v+0ycDhLYCnRIm3ZSUkI5xtTG
oD+V333D5Y+UqxsznKncxoy8jfjQYLeP7biLBfs28pG9ZGKmpXUe3fhRpFlGY1aI
tNTtmOOZLW+7+rRkv0cjR55lN2+XXMrc/hg2RwnvHJVpDmJEjzaHdPdBQJUzuOnV
9G7Ko6uj9ZbmGQMaMGRiHAX4G+4np7/+G302bVRU3qXgBcGfYoo3hImVCRL1yxpt
7MNZn3RNKIm/bmCn7M/ued6S3UQBue97hbaiJULgefB8qimgnZgDt0gTQ4ep//5D
9fKJeWOn8/JMjh0VXSFm9PBtvCDCBvk+dY44Onc+uW2ATz+VtDpMk4GR694FXiy3
G8tVnhtwmSb2C8rKVjh8gtxy2ag90llkHi3jthmfKjzA7ptySuAYTVEbX8Mjpelf
lZps3dPMB34le9JzCoIYdsfdRNj/jjMeCWuFfaXxvZIH+WHdOCoesQby5ifxu3sB
mzZeqSgz2J1b2elri8cfCa9P9/3EzK62OIIa6iOACVySoGyqNZQSWkciDeqdDHvN
aVWuWojXENlQ6SsNKoSVysTXmqF5e3/djcfDN0BFvjexoMYt+DZIvaOYsjwWBv+K
5U1cqMQLOfreMCGIavdx6VaDLFJ78qkKu5zjZYKjhYtB8T8QbRNehIAlxroxxxEz
TNSwyZR2cOywr+8/Fh62DP4xbdzSltNousLoScdKVI7BUpXLsNhX1z32Ibo5BBhp
runlz5gl4Vsu1U7rC8s+zLx/+8HQ1u506ktS77Kx/Ia5rCJ0koqIEt/AIiUQEtZY
HMs4Xc1y8y7Ai+Kc5i6Cs1OOveJLfiHkMj4izblHOu/EbwS2qkK7HZ3qI1YvyYv4
1o45bLLBaSx3m7rRXojiaKcE5lr7/vzLbluB42dyhqrtfe9kN3A+mV6+smVPVPpP
SgwJGvVWTIpVkyfo+1XALYG0Fbur5eFhcM/8mdEpfwd78j7hpPrmwvjbIt6oVB2a
EZmiD6ohjjelf08A+fN7GxLcr7j3OeNdZxJWg0WqiXR/06sLF7G/sPjGMjygp5QS
wxJf7nY0VpYDg3kRRuDCOxINVWLxOVJnhAJoe6DgHDyvpO7HUTfNC7ykvBMXu7qT
ppyKJmVKCT0PRGQBD0ri//TjmNbKWkf/OEAIFo0XC4EDnUk0be2IDD2fpGhFq5z5
JQLTBacyVEN95zcQnjTssaXL3A3G65xx2UunoSem06FsQI4QoJCx7enwhpojM5i1
QfPOJWVe7d75FVnKxSfgv5cjyfvJX1T7ZQXYoHxgzDoH5UKyDLc/B2EP1q2ecKYi
Q0iCCxGMpoz76qHumsEapVZthvjqlDdEOq5gJ7KwWT2KcOgBFqQcnelzs1ZWppI5
rMt/XzpfYE860j7Q8Q3+yEsajyZO6u1eiV5myW/FdMj3OZwHqMEgewgk6fuWN6Xm
VNGzyeG3uMiwsw2EsGfN36j9FqpOybTDvXnphLxB76c0+PntrcM4Su22JefRgrY0
pfP8yyKv1C2wsq6O2cqW4yEGUbL4DhmCxrg1xHA2CrQCfepNrklMIIuUx+Kehxua
FnH/3tfHAbqrkc9aCluq1HfDnd7NEn19MJ07+ncwBVqsyKo+O+M9Occjq8ABtpfJ
xbaDDyjiHN0rf7R7srjAgMQ+T4/NGwpsQ+N8k/99V2Q6j5yakKamCE4WJYh3Y5Hx
LFIR4mKNUfL36RW14kjeLJxMgN1ZbotVKP+GNW82iqOuGysWvNTkZLlvkXpGEk2s
JbBYaVXrhXr2ywDg9AY8I4MWY1vVCtpQ5cZUQqONMGKk8UaP9MeRrwfqJk7+eqB9
N68/AiHWdPwawBwlvNCfwxPQb+vlclfrzVbFzK9mUosBNM/ZO1Q92OOyCPeFd9HR
wAGcOws2TPBYa+YZLerL8bHbcZdqYXsM2nQIA09yJK2/iX1LKe+Ps68s3khC6q+K
Idr9JmWWK9/dzvAIvp8HIbNiQ6mJsv4b5snL8fqP1L6LtL/g6JFgP2+CEapmbg04
qMW2HAGE/RBG1z2F2Q6luCcHmJcWs6uxyeEvv+ccVHi8H7S6G0LTOiPcnZKORtms
X/ha3PjAJkWWmujq7dKhm0JvPreUtVDfcmb+CnfDOq01NtHHMURS6mfLU0Emt0Jb
1UerxMgdYWoEPUChA0sjL5Ye4G3P9O9lMIcQeYo4B3mlgmJXphRRjeWWpoXEq/ni
LL84+JTjOqUCKF+OcH3MQFviRDlwKBjyZ/x8XyxAZXFG7o8x1GtNfU8/l8gRmHIg
d96dwykiYzVKZJ6kkoANzZblE0g3cNY0S2+kMX7ybqYfZyp0U6ihfjzCPXcmpnjt
nkGZB7Ji9mAZg7fwvAmXwSsvSuO9cn2M+9LkWXuMEgqoFbeWK+nfgUzkbLU3Qmd1
1M7LThhDfqCnXaqLKfvDu5itA+Svz/L9O20pbRwtXzALE/TuK3YHGOUK/k44ly7L
Qd9Pk7qL4SgwX5HT7lkOgyoxBRZu4KmBZ+y/miMA7jl4Cw31kdmrnPWxnYbrXhHK
3zu+PZNpxSBA/zs4P7JPTxnIaY8+GmdyJfv8z8SpNo3JUDrtOkfFJAzCGzyrup8v
9JbzN62ZSlLF17F2NGHfbM89mn6W8W3udzsQlpxo8p2cVa015RK+tOPK5EyTaiXO
p4usTtp4q7ttornejujRdvYVMp3XjKJizjWtVk5jwy9RyRnioaCEGwsXW1XMENe6
ldSjO96OQP5ZfiwMJVAx8jpmkGw5OUHw6Wgl1BAuU7FGhKBoPj9XIfkbuhwIdwEx
jEnx2Avg/a0lvMgAqEuHeegSqEMeJSVEM5CHbR9p7/6BZGuC5a3A6YsTCSLZT8YL
4MQT0NvuDqGR0jXKwU1b/2I+yqQfvwqpbGDSDuBOZI54wlRHWl0oTfQgFktXIT17
7Jql5KaC3zYNlzhm2lyNf6Xo5tqetzinDzKIaDnrMesQCpmZXwmyXpgHybPHVGkD
M5MCwliJKek0mQB6hRg/9BGa7H6tdlXX07IuVIHr8pY+9fCWPu+Xwow/2X/PMAEW
e37FC/nIu06yZ5LrOL+rWBDXuQG0z/B2nzdPq1YcANFGtJJKdX7+shqOK01rzDmh
74Mnk+rFwtPUXqOMtD0RBhEGiKxq6khXxQxQF21Qne+9zqZYrG9aw14p4mwoBFnA
9sRtaeAxWt16osAA9Rwq6PYXSktpnfSDXWzeR1atGYaa1QTBJ76sistF4tulu5Q/
dFrCEByCrAv2xwXYH8oTb08ZFGIjB0het3TP5dcYtv/iofEd4VS7DNC8xJvX0wGN
ppfcUoDlAm+5efVCZnmM/amwGRnsjQKAjXvmW3wvxMthkC4EB3A24GwEpoQRNvTS
K0oRBxINtuDorGhcOnDAJoyfeOU9GXWaU1gUVa75hWGOw/nWpRQ/yFpWXJ5a86uY
RvzoPBRGagu6lhYukgzS3SdTx9SEFTnVC9VIKyM69p7kyDxS994iDfWp56flTxxq
vqEYNtktBsO6hdJMhVgA6AvJKcPeK2BxDrXukkyp3KC4wFD+8Vd75r2IocO7W7Y5
jmCwzHuCUMw+x7TS0EWD3Wi0kE+DSsbLt9fKQu8D4H1hRfBLF301pCK+Oki5Fw9Z
RQAkmviEV/DVvljm7fX5VHfUrjSU0kDOVMbBrLLXUfbTvgBgSwb0ss9kPN3Tkqk5
9vxPPSq5abSLRWeF3x1fMVaOf3u3H4M/fHFB41CHsH7+89XF+kYtYFthPQGz+Cvj
3PDxgWWNYZ5fUWMnrWhIfJzBX1eGnqjd3Fl8C3v3Mt2UITCnOKs/Mq3EUdCwQWp8
64CVuOY0qNEjJ7pPyhRgOLa8mawNYFrjn/1DOKhL2Jw5UFPcb4raqQc0iYY0bPwO
0d6Uf7bSRwuZ0qXiIagwSp7+Iy4MIJoca8o6ZOLCeuOCVXpPitCvcGx6O1bJ2LVR
5FaYfypgj0LiDxbYZmLKneoFZTz0vmEASxAmzbWsLwwFR+VBEiutC7HPuxxRYB9j
GVggh5cVRKHcSceurd+8b6ZXnl484CkUve5f1EH1iQmdS2rH9yNS3NGK+2tNQoFz
dVoSoEYoJa5V8pL8ahx/WqO2XAHVXbl8Kp+c7EWge1UwxLHj2tIzJYyF3vms14ua
OayCUq03/HhYNmOS41VMM5gsl1QlTXEJxiMRCHja6IyNk5xlUBuspnjuVJUbErZK
1843f7EDvW2oAEuOjJc5GbwiR1nuIBlG5dxZ5+oxJaFwkiaiJF+j51Z0hCG1LAL4
qjIE/lqO0ryvJLzK4B8WQZPObUbia3t7KB8QHWrBgJ6AHiEr+1ZF1PtWnxFjhHV/
F94X4IC1CIPOFGiWOpiO4ALPEg0X+0NfK+w6ShzDEZg23eOqPHLVVwtfJMvHAZ+P
3j24OmzbDdnyVgRPKAZbEt1d0BR8bSD6QVrCQyr4V9xdgawyuYXE93CtWZBWTjtp
5C2k2lDaNqQJjdThx+V7kc2i9iA2Km30A+LDdOeejREPNy2fD5s1nGgc7VbAY2hE
3WSJpqdjHDti6uWBrzDEOCVzrKMP6J75OQRM9c4HEXealiM/2JhMp3uWZPqNhCSE
UHYJRripJASeMKZPG0gS4zDBJWcdHw6b8mhYdLVfwpOmRwnAbg93unvIq2Zgw9SE
3bzEFKAZzqZ9OL8taYJs/b8qrij8Y1SL2QVVYAQ8QVnWfxl63LAM9Bq++7dwpCSu
+QBmwVXkdgAdJ48hJXnPxogKaMyEZb828fVGJoh1ZGTjGpRr5I4tb5airMfaV/3L
V4ifEOCrUiXyQc1ONt9WEsHnhqpKRBMvRBHXMBWfCbkf+OG4shYxZGf20F1SZCn7
LgJxqU4IRiqn08tdHjhlxNUWULSUf8QfU7ZYSDxYVBnHRk6LCB97D80O7wOA3a2X
o67sQu9bYGpbq7MFlJlh7obTmdM6Cf0+Feqk1iGrXr/GOqKykJTO3qAfNiMpmwBg
th5KpEVIqsUTgVM8ObKH6XMOghO7DVHXNhfpWcNa6nvv5s0ebfj76J2hRdtfrn5N
ySN+6cNir50dibKrw7xgp0/+bdFa7M73C+L61gxAiIC+OIKcA2LcFgQyjJAAY7Sd
hjYYTx5n4q0udkSdsW52MRi+C7plLuhRYv7bcbnJAV/sueApCyrlZkIMdxAx3en+
rfI2Vo3pniJN1e2GvWGyGYAhbNLtT67/jilQppGa80FN4n4QFTZVOVpKpJDTQZjz
UqejaDotKqD733+7yZm283UAjDYi9XqchcFiZUf7/ZXoFK0t2aaAh3mr//Yyw28O
PtHGk9TT/R8uKQp739+A8A+haN7MSdMzSJQjOCp82h36+QESGJ8FiX+DH9A744mF
RPxAB71Ew6oG5jSrsCT83eQkAJQlUEzBj+0k0iVfl2PUxKH1FLHXMhxvGQr3je1V
NM7bVT4pihPxtZ7wMNjIzCicF0WyQcHDaRGSHU3tlNznZpcVcVSMAYKzIM5sxss+
RGzEEX8NduaSvC40mf9/pEHjg9LyuIHcglXwwZBaUm8yuPClZei8SCdNSVTVysGW
L0vj+un6LuM+NR57gAv+JRqTjIRyxnuYux6mQQuuzcrnJiLp4sccPQABNBzGRSla
QbV2CaWuqJUV3JHckbjnzQOE1B/UP14jHAk3miTNDT7Lxzno4YWkdzYm3vJLHpcN
XjN6f+i0JVWAcQ7a3fIYlKDGuX3jxLXHJ+eLNqYeJ12sdfKuT7DJZ5wSjgGfpykW
kvM1LtO6k2Ol125XtVj8i+TxKcyQeHN2VG2d7laACPDoOJQ7IHzy5Uu0v19icBbj
JZVVBfIyACPfl6xcxsDi6WrWa/q7nXxFxdhRDRXq+/Bjh4ecCmIj5x2Ee1OyCRnq
m83gPQTata3ps1d42UnCb6Dehomy3Jmsrt4zpGhvRjVbj11opeNNl8i2B7/Jh7QF
E9nBm1DKvdFyOalz8MZDj04OGb+zTscXR1r/qkiYdpDoayHxi8oE96sJnm5UK/hS
SD6BSNmVA/lzH2XcPB1zUg+r8dE0p2BoCKZUN/BAFDK/4l1LAuhwZXFte4NobFBl
BxgTe/CCcvBGhg9YR8GMsSmpNldWiN+VX2HeXqOpBfD0A7npaU3WBEoKkHCWnxNL
OCO3OONA86ovjNHMYCwMd1gDBnl3H8JQvuBTXMMK9msG3cjNUulYUn8HS77gOmey
j3Nx3HwmuU6+Rdw3Wx06wQE6ruamygttXXqB5Usp55oSaPi2OCWl8LJ5Z3ppioGA
Ode8+Kob7HZjCoA8ORefa5HdtM+qTr4Cn+FMECXdBPcH/jvlqLLqlIvF7+FfhymI
qrTnYT6cTLdnI6+Mdd7qzvd31+HXMrb/MbL3sGT6ezRVv6piCp2KnmL40jfRfnwn
PFDV39u+HOdf7bX+w3e9pHKPA4TQJ0UDB2krqzB3CPQxJ+SabTx6ipA2CChYnbUZ
v4mkXrWhxKe1N5OVTWIUXN5Q7KPDh/Bd0sAKGgUBcCCTgK6ZtU8ywbGR++8x95Tf
ovUXylMcCICAzJF/JUopQuBz+M85sDF1F4VMHcKjWaSf8uUNigD7tAHrj/a6gWHj
Fl9PS+bBqCrOcDESjumPsG6mgC5nYWveEyzRDws/Cep/fC5nBZFpn5q69gZg3+32
cneFv705dZ/NWvc1dxEtd4uUxwAAWvyRyJsEueMxVdMGCSXrK55bLnUim4m9tl4i
0zZZyAIq1RTeg+mBYyOyWy4wCDBZSnRLUng+hkMcUVGFC3qQXYC6XJJ2FukGD0CI
5vu7gHIY3Zjv9KoGXaIKTYAHJsaDnQ34jsFpwmCrYEjcPvUUT69tJysdVB5cnGQ1
5OY1/A/F2ibMearcz/M791AdTGKGvdaMoScAAZkiwJgNpCF6FIdQzmxEM0jpwBWQ
Xm/Yn2kZODCjrVrWHkWnPWC4VKtKJO5ImJeInRZZa9Gk8cw7LLYv8pT3LLdnFDet
Dog8Q515RGxNKYc6ufMgq1ebc88sBnB5RmrMhV2PqAAP25dDxGhwJ0ScM+FU3ewB
PTtuXl0U64eIm6W8mSUkeOtsVt8Z8vnNYkxK7J70wTrYlBBBR0eSNcqGGs2+DiB3
iDDemr1UZWO2GKnt4BMZMXYgbzdvNHdj/tPq+/glfu/ATFANIcf750Or/Vk133DQ
lZYdlhJMOuDNptY1TatxAe4SdWRHwijiPXVymTW4bM3rjMQIC9WMOGOQ5vwAILrE
KyEatUcAAx7omdk5+/nyxsB4EPnkiA/N0NgYjXF2Jcj8J2CB+zAL751jeSG3Ezp6
K9UHlukEhTS6HHv+5BgcCxh2AK3ILoTznsb0R7IEgeo5smDZspyy9NHo+FWRlLKk
ribl85PtpJX+BycitOWHsnKTksjs/TMtSq30kviDxkO/xyKDJ0ZlJcCof9M59PrC
yhrLdJY3vxFLVdQpu+LDlx3u2XDpv77tVkw/6KvAink8NOoZpyeDt+pvdXqCFzGX
Djy+afawDT8FovaeV71erDOPp3I+oDvcDC1b8E/qzWFN2Ue0laqvE7r3BlgYKgFi
AYzGYzM5pUB1AxqKJgDH1RgORhb39yRJQ5E/WRhxf6JEOm/AQ0B0C3bCkC1vGO65
prhmUPB/6t7ukXjwX1NkmJiq11u6ptPt2hFiBBcy7yJ6sds5o9GqiO4Oc33wKTGJ
8tS3Q9+g0qeyIUh5jkp+wY3AfkDoqCIaBecYvQsc2DCIESWaKrjsYU4w8l/oRTJ7
c99DXHgM3ashG5GQhAhQr7TpVgt3l09UUp8aP8mX8nHw3Xt7xN9HBy2bxJY7ShTE
wP5J0LmbwGHuy9xe+gQvy4vaGnlF5n9Ef891caHO/xxZCQlLysx0X4phHQ0PH4Wv
peNlGZGvM55tw8UUVL+wr2OUHFBvTDQOhFfjxzb0LmIW5pcD79E5QvTJ7jihq48U
2iFVse01Lfm34qT+jr6MqTQfUENrmS6cY+C5t+yokVeUk6cUXMwfISvwU37GOrLJ
d/phVoTG1CxTyDmfdkF+ux+TDNZ6HN+cThyRFe9hd8N3UGdpV2dl6/8vPpo85AZ6
todBs+YelHBDXe+1yoEX+vyv/6lviudhFOq8RnANNBt3Q0d+mWXEg2JAFCJQJzmY
kwdtUGviOzdk2QDHTHPGLsx/3B2QntHzpAaBCy+3D/XkDy/lXcJOYiDoFQphB8Os
nlC2ZKIl00yUSWc3/Elrtjru80oe+NSzwOJ3A2NRtjTpgWettUfY5TF4TjylzD3e
sp2sX61vNL0muWEZYBQsO7Tsfu4AAC3a2jeYDPaI/SIqvQZrwD9MlTqu25HyCPi1
gzr7dk/+qiGHW8va/Sf4GcyCMQxaeniu97+BI9+ha/VYlLRz3LIUgB3wDXezuF/V
p+ohj2MshIFqaWWoQMsUtkhbOGkemE/cL+/E1fapl9EnKhh1iwgGrMh4TkTUFQt2
qrPfy1/1jCf90eyXQAkQSrdGVBYHjUf1QH4IPpshM6jNw4f5t2j5XNpbTNlvWpvX
UgSZVODuPqxAczGBMDxRMzqoCL3bbi3m5cBWsJqeDJXcze5VvgbJkuhkI4cf61Tv
/Lqn2+FeLryVI+JhI25JAeY+1tkALOklQS6tTFdddY0qngnZdOiuZvq2ChJfzvKI
VTNRCaAOUikwRMrZztblczOZZ0xfXmPlxNev8IKlmyyIyDRIG5KS1wsMKsWN5AHO
RFsGVFdyzrCkmlKja8M5+Xp9qAYHA/nVOhI+2q+1PRmJkhKHu5VBkI06P7cDxJaG
S7T9VaALLVDKrRYSGMl4zXuWAVaHmvVf65X0dAz9VD2JQLX5qQ/oD5QxJbhXR1/o
bXkhfzHK0iJkLMy4931mzN37IxYbkrjhXvXv0ADEyh2UzImnjVOSaHNAQUDB1Qlp
UqpWMOSboLH96Ps4oKO0EO1ld0NpZhblr2KSunzMEDjpAyHIlCkHshI4Ks2BsY+x
jEfyfs9N7h0s6cV+6FcbdLAs8fVsMWMeXdK3y783lIDQ6qWtGQXhG+VDOsRAFisR
d7Azus92nVeReeRhQfVgeq0WHuQDejHsk0dVtE2HOuHaJW0oIy3zaCplHAIlFaeF
7KgwIxNEc6GDpdjFoYUODyLm0k0XSkgSK9nYJZHMc867Z6ugVlqc5Z6HV8Tn12Fx
7WCRrn7TeunyVDI5NNDgjQSaO3q4xHZz9aLxfZ7Z9gUaqOuEkblXVrSaz66PrnMH
yaPEaGRqotU6c76c6OouFa4v8Zr2HJNRcZdOiyMHZMrTO52iuD7aTcj0r0t7Teea
XppO9RnA/dZL2wo0T+6q+mw276hY/LA3sMuJqLrJ85/wzqXBSyZBj9J1quZiBKXz
Lu0sCpvEuLe0sRWJc4i3O7tRWt8UO26Lp1zKInHGwUtsdRp6LiJ7ou7DF9Q72U+j
ysmGB47rgfDAEj/1GMOWd5QlJUA9GYqBFYhxJbGWWXlB6XvczObnsQ6+60Ls5SXL
ByxlzZGFZ8HC1OfuOSIzL+sCwKpr+6c8wNYZEZR5LM5LvSnQoBBqnUYAkrIyF2Ev
pJ6YEDsub8rfX4jB5WQIH+te2JT7WCekwAUwNf+RPDER0fu1Sz8nJxZso94EusXa
Vf04iOD0bc8W10j20q7VDj4QZgQF5Rd/XPT7Mc/7DKaTWjg9OMgEHLvIJpAX8/yL
J65zD2OpYge3ev/ev/8d8jyToiLUDmVKDsN68XY+q1PvKHJdLCJYR2JnqX46QruA
m0s5eCAjn52hK9mtC2auJCPXWUmzD/oftuSkNyb4Dq4dkSlhrfrZuwQbTtRn4t9o
AEldFfddJ2drT1ow83V1a5UrodqI9GQDafQdDJwvKaxhSsKCVTWGNnZTPZuLGnWt
e611vjJEEjw2IDssPhZ4nT6/XWAnTeiTIcHahs+tbYGJXm/QTxbfCrV0FnYwvIaP
Zw+9kmi0S7k7yahhpLqLB+7Km1RcpVZ2aM5Q1W/9NqQNGuObSex5tzP0vugUhMEN
y0Uq9h1nxtqJe7KCYIkfalfjcQVpyscUq7luYOYsoXyIhsfvEVaZIX68sYsSr1RY
1V3hUxi9TuqatzYQmw3fC3+bdD5WyV2KLgfeaMieWQvl9Gr6LADJifLDIckMs70X
+HSnNwV/Zz6Tiuz2aseyWWtN+ZRh1+o0ohmu3mVPKcpPONAq6YUsxmsVvWe9Rem/
FkxALC1rbxx8bP/5cFgIJqsScNAwgFM0rQF2MdfvTG4I5RZp8CUdl+YKfAtFF64b
3l+qZbqRiXru0XykWuoSKfyYzjHKiqYaB1mCgRxtNQieoxzRH3M797WacQer7lfS
bRRuKlD86GNX+Ne6MQLlZ2b5Tc97lqlGlSYX1PhlOA/PJ6p9Iy6lJLbnuzdi/U1d
0Vamm5A/9g/dmgf7dhqWhc4FKTWntflGtwwuqpeSCxXYhBEjjce5s7InQGA3rrcW
f2Htu2rEfhS5X011lRdAQdiur+sgNIjlee38x2ZMcWEdgvmhF4G0UrBtDu5ZcMTs
jyf0fGoe1jPiYEFEooeQkbe5WG59voRMTgnzKK4waDo2/OSSe81naMbvt5zS1xGH
osbfF1yXipSCEkOXOGXABqLGkUYkndRdVKf7RWOM7C/Ifrg0tLpcAXCQOyuIASoP
zvbt/8ort3ApqXfqskuPxGd2pKHPfFOHrtjRZOrsN6r3ZRN8rh6eRDGEWKSBkW90
5JCO1ihxe21ZNKAyNWCGiOSKSBrS+QnHSQvw1iga4A1uu19HQhjWeCfS8HCP2epU
spMfKTe9vg1ul3F8BLYpW5/nenPwWCtK+SjyUzUEhO0cMgwbLk0XCPC/Lf3oySVy
VxAAd0uWfGqjOH4TjXHP7zBafnMcBU5K8oCONkd2uPjoab3vwx0+xXThC3yyA4mK
zKue0SnVJ0eygYRAleLwd/gFc4YWK1tpweyxguQ6A9ZnMHLN+3lJJvQfes3Kg8EN
7/w7eJZiruhTV6TzBJ18NKulc2oZ5sbt3rEEsYSBiceKpQk1tBDpdtnFDIlg4fvD
AplutEpZiMBzAzPqsoHJQbidveqhEQw4+bxLBlyadnbQQ6N88YAyCotiBig57Kvi
JoueVohNn+Mm9iXe2TU/nyFuRe7xsal28+NcTwL8VaoZ/t7sRyUaJA3bS7z3OWnc
GJ3ZB15Ub5luoUZjRmOb71YJD5NJuGJMOx1w4rzy2smho6famXBuNUSTC4Qf/DvB
S4yRNis4ebfwcVyDb7Z5t368pjbquwM8e3tFRLfDMl2xZTtdwdl4nuO0zjIpTWBS
3DCtLlv4LjE+cd0gF1o2YS4WnDDeesa5EobXWQ5g6NQTIo+j0JeIZYoNF8Kebmma
qhARWjdvAiRiYWldKJp5MtWdqAvuRLd8ACsCivDwJl16BAPzTzZkoSF+T9USW1uj
7AEKDzeIS2+etHBuyN1j0brGSesCjN6z0OBAcgVLtAMPR9X7CdggITrVaPsryYsE
SjzbOYMHS+k874AXzNeIN4R8Y329zC3BwCyazEZVOgPgdpi+PUObXPZxHb9FElLR
cdE0zjcdp88k1nDY7J0hXomTVuCgmHm9OoafzNS0QzjvnCKa/cQugVMJYPGS5vWe
9uyB5HmsYPQ0IpH5lvJo+3TkWczjtWtGcmt36KxWbM4qLss3925+CKxQlUPLmdHD
/EprOP0zGTcGVZxx6zDJ7H9KJhMd1Ye3AuKCYVTgjc8Tp4KbMQW131VlGTJCIpMz
/DIK5UhfnqKITocwLCf28Tez8bxq+l5cWKevPK1ROL952B6lWyItqdg2k7PtwB3e
uwp7FfX3KLBfmSXXIgTuiYRw7W0dILTLuViCMOAfb43Uyc+k06g+0eFaQXv4t0SW
CKJmjneao/9EAHv4uJgY/yOJrlhyNyXvyL64xu0fiqcgmnhARgYyvF0YDYZKDiKW
PI71IagmwHKlhjS5glFcDBNtLXvkECnUAHcnIxWh3wCbued4ayq8R5mQekuI/GL2
6p/pg9sSsUcB5cPj1F6gQMXFP75vNEjAcu+iEco+/WQzG7VMAa25z0Ef/+gjrNNW
NLgdsC+sg3fxpVSRAhT167nxcu3wNg9brNbOBZAJmGj6iyvJdfWfs2plJi9fFGyL
0GPYwWWfFNCBdLV7f1WMX2RVBp/C0JKHqewiKq+OOmMzrI5XVJNRbjn+Q3YRkxLs
O8HZZaGFflcmiijk/GYE7wiig4eohJJ7iAuvxpwlXbaTRidZfTMZHm/mni6io73Q
CYzeOdouY5ZvhxNWB5LU+bHw4QeV5u5QD2d3B8xpg7E5uVIbeGV+/WyO35cE6GHO
FUgFhfZFAIVbh9kAFjfpLgQoN0cRwMyOkjoDClWDdJlY+8XCO0kdQqjJHmSJGZe7
00aHX+PCuNnfqLDU0+H/eAuxts00El1bnofsbQfgZmoPs6r8nylvCcKkGWOfT7aI
sduxio1r2VAFr2n1J6gWAKfRQlDWSyXH88qcCsjFSms0dTk4fLc+V7LpuevCmzF5
6lqtHD7n6VNcVH/PrTLKv+Pi3jo29D6TH23EzpcbBmLYu7+vl//yShYYXHj4FZ+C
m/itbW1Gf5eZNCh0NqPetyxDITrwRgZkXW7RuJLXSm8p/rflFVzp3piXYG7RDpbN
U2iCNvtTvzjFn7BBE3LiRIVbogTyMG/VNB2ctE4nZo+53BERZJLbCrFqSJgkW1p0
oJKTRSSEwDIorZorBAHsKvinP04b3tT2QfdS/yXwE/imwfDhm9A88BgIQCuT4gha
oihaZmQmOoD2VIzFmypwFy3wgE9TBDWg3I4YmXpKs+mD0X341/R9qYtS4AavK/02
FTPXZ8T/2acVj5OWcznn3rl+d9rpR0B4JMwiBpLjp8wJuYQYEI9IPyKRXxOGAI4x
Y/+JcM51QIyphya7Sp3LmS3CyvhAPqaI660gOKT3NEatD2VBAIGVWiFPEOCx8hfF
0bVFEoDNRrYbp6CbIe9SU+xgQ23M1sjp4+l3d/IdsxziKF/lk5iE7sLnh2h1BFme
oMqu8ess/1rjL+bjrs3IyflNKh15G4Kx4UvjblrVANWQqKIzwT5LEGGV3T0BA8kJ
g3oLK8BghKCbLgW4HfB1gwv2sH4/L10lCgmjhUwYDG4rpVt6/AcMTv26eQfdpPiH
p+KuiBI3B6+TL6QlWdYk/fjxhwG1N2UN9xrLW10flFkUmgz7ryIxNhwBeA+rVgGF
i0wtioGIPZJ+IsNl0CtFQAL0lWwxGXmaipQBSuuP3QyVEDXI2UKU9VToT0oJbo3Y
lU+giwNVoNh98B5gSJBs0et6d3StCNvf670CNvQ9ksaBNyN+FB0K1QJfIaAmXDqr
gwGD6u+nQRCoKNhZXrnwsTMvVVs01RuJavj6QGlKY9Ih6bLHC7vLk1XvE3zG0Dop
9+hINs/UjMtXdZnL6aqKoD1pGGMmT/kjlfgvCF5wF84HchrMeZiVMptdWIkvJ4KE
91Ika7VzeGN20jIKdkIIOZ0LjxbB45/8i2HZmfp+4cgc/UVuG0dTClUes9oQcwv6
ahz5TOd145l6FDi5s2Lw5rWmoCSq77YmFozzrK+zPGxqSBaLMbZhEtMKNLA8kMYS
I4k21zo2A+H9mrKkzYTmd6B3zXn0Jx/kt31Zy3IZtA69wAHqYNhMSHadHt0qL1Hc
qKiUpR56hcR6u7oDkAQQRfY082x/DRITl1i8LoUTRwaI34YB0MI+me4f1UFgISx0
+7QW0pKmrN0AEMQ/FNVQ+iJu3H9qWLa4EjSPai1M4Bzvjdkab/Riv104fIzDXFgC
CaY8GHLQzh5D2bUEQsGF+AxZ0ep4RLbP924fod63YKOtDU2NtBCr/jw3HEwYfwoH
r5ACnmgkW0XfNQByzTPBXSLHxRepeca9RJM8I55Gu17/782HatYEgR3wyJ8UcKWo
l8r0V2sRgWeuB0pW3Lzhd8NaTo7P4cPnh6P919W5N1/v5NZ/Xa156qBNo2q21oTE
T72+h/+RTDut5DzIIXIB7EiQoIqzwRhsJfZ5B/V8ld6pg6irv0+9QqYG2fvQgRRp
//L7lPjLnMHm1bEGI7nmlNOnO96luO46+pxx7+ObcU4OIN+xQZL1IqvXmXufo+pd
U79CoofLBZuM163gj+Kyfis2pIClCV5As2LojXdTnBc+jWpS1dtoiIvGFu5bgQ+L
RQi2X2vWITCSI6yZ65v+cKzsyPPdMHKC0FQXG1Iz8USx8Dt2naswqKkxn6OeACyO
P8JmUudfNu/YnuQLx0FxoYayJP1my15liFwlCW+9aaYOW4M6478pLCsx/99w5ZgP
3jE80/lvoRdI79QAOHmoD7l+lig5lqFMFLsVIttFqL0TYgdC4Qakc39cbUgs4t4u
xE5WfmD6jx1ZFjdbM76uR5EBpIArG4PXEscaeW6KoY5nSl+9XGANhXXCie+2HFtn
E8ALNV156NV53zXzia0BI6Ao0eb9PgUQqdod+00XZWDOZeuVzdr33rhWSxVgVOQG
ucskEMA5BE/H6MJAHLBamcCPjO1cWiSOtrQIotsEt1lhmT7/9bL0y3lGbT39jYSO
AZds11q59EsyLPD0PMWALnWjj1kp900zSApZVHX0pdhupku2SXnBze6s0UkWdIp9
XgCF+3klW5HGexzH6ekaWLrN2vfDsQtqjlqLElM2cmE+S0/b3/HlYlPY0XAdUpps
eWVehPq2Z3lHdX6UeOrfDxNn6xE5stuD3ZCeuQ2bOVISD09Vd3LcApRsSNmVM3xJ
XPjM7y/29twlBupmaesKO+Kc8OzitFLuY+DiJj8olDgBlj9B9bSkX8IiyN9FOHwq
V3wfthkEV9x9zYahV6wNYlMijfM8APZefSvdiDT/GazAA2ayt7myBJNB7ZzCMRn5
GyE4MhIYYnfM+KrC3zmILAdxvpchIAox6xMJ7qB9Liz/3tZgL/utyhqpNavCilPY
uaLjzvpw6cKpszF7mTX7C2BiR8vmROUWywlScAYOtYq3NvC3TahpaqGq6e6244o0
i77IYZIdg8tk60etVwoQKpK9dqQ94kq1wcRGwc9kVUb9LZTbSAi1kxLARc4QR/Lj
QQ5g8k53Uu8+yg5KrRwpY3PO9IbU+CwxG5d8eCyA/qkKx8ttCYczy89PHXupv8uS
dGKbUWgvsuTc3YUQhfI6ocF1h2Otj/ojPp3CTiUYu6LVxn+IThc6tlOeOQ/+5/9o
rPO6eZUuVkhD6ZNPRTtqnWoYv2lmL+qsgYecQOe49Q3G2BQBJ3T8/fTRNwVg0uUG
K8LWZOD2MULxE0PeB2ghZyY1TvjBB/CR3IirNH1NAhx4cSkUTeJZjH02Tla1VMQC
Rhxcwe7ELQhdbNkYMpZe4/EnQLsGMem1Q/HFmzg1hZU55/HxNP2iics/aKl3Gfa6
TLZax0CIs/0DFaI44gToA0CkrdKfsvX5Re/z31go4HKmJddKkgdQHsO40dajkUWk
/A5HuJKbMj/OC8LIhQ8knrIhML2xX+syRG0UESc56O8n6QmElimu7/ri6+gTz26U
BN9PEyhftAgHDlSXFOKaLPX0MT56mFzDMbYQJr0UDl+cmPXHO7mcPsyF/N19EdT0
B5ov6VOq1Hq742u5adlFKqOM938p8x2aMHovoUGwE/vQEF6GsBtQeiqGNcpLu20K
W3+1B7uiuKtXgUd/1MEIpl4Zeg3mmQj+6VzkkC9S884QgsJ5GdTaHkSpietmfP6T
d6bqC8r8rshYt/zJeh9jXp0/DByiOVuaVTGEFZD4fBlE1Yc1nEanUdF6oy/MYLNF
r+9vBKihahyIOB/gxjvWTxOTKRkRnCPya3MiS46OuLPVokuxwkH0Y+wZ9mDSKWwu
QBOzMDvCXifEG5vUVATcOwXs8Ie6dRM655Mazi8eSMpbSU5uLHCGK3UrSpwoWfIy
tGrJrgF6r2ppAmKyIYrH9eahSEU8HIoUEra+LWDzy/KTRLTTCUGsUHd6rMBlWGTg
k0f5Htv+P32NoEXIYlX2w0+t0VllPhlB+It+FmIllsCutnk387tHIyB8AtantRkI
IbHKSN0frkaGSE7/REJs1EOwoWeNDJ8rBCDvNfDqNPv5iZ6MFIchxQ5t3nF1Ntaw
9upJRWYzkkGTtBaDdDLucWHMSGenZnblHQvZITY52/pN4ac7jBrQBd93m9ZBm4Dz
22lHGs+OtihjPto8v734Jy1rHt/fKzdkRv05R8Vnwr44BAneVgkmwvUTBnSXuJar
TocC1yikus36kexFaeCcliqLzFIggOlG8UlIU8qQzrcWh95mXrgV24/4e5pdIjGa
mIzPLN29V34rg/Otllwyn05Qiy+Owuwfsgwy1hGwShsoOlXFx7PZYzSbriQFOUyn
9KcNtwaJHFdht6Ec/rIBzqDU7FBzO42MxA7yTP6Hm1E8ZCJ7JDs6ShpTqw/N/ube
vZM316TI8vrga51pmHQXvlRMuaY+8jKRlPErLWDMSzexm5W+cAYZLcFjMEghbbQj
DiJIZAbt2VuhjFsaNUfRzAn3btN12gZm/emiZzQvpvlsqB44LqEwsVEyCjbRf2Fe
4vEFdcbBXmBHR4vjHZAWPT5RlojhY50A1GyMxKapHZmPBvOGz16OJlrk8YzxuiLv
111upL52AVnXrafRKmMwtl5UfLPp+ZoTnW/v8nHZjvn64pNsPOtpHNLaqcP7qHVX
ojxdMbpv7KP8bWs7mel0yYMtAlvWnO0fBMCfN6m372gLWXaQ4ZGXyDxkpdVUBYwo
1HHKF78/Nm0Fc9pDzq9wZeSIUfJ+R0W4/pFMXJ7QDW8KGl0qH7+zqYE2smwItYMF
3UR+JDLweazfDY9p3mL9DNm5jRllNF6xyHGG1N/N1q8UOEwTXtebZzRGzeT9H0aK
UpUNR8FgFwCMSKLdOopHQwmqpTY5wqaO8vsI+XnXRC7/hssSpzS6stJ2xgo8SgpS
CKaNEHcC60pwmjUUeQ/3y19d8GjGwjwXU5s8VvyaBvG3Q50OfVQEIbGhEhjmK82o
HejYS3kIIK59tl5MLD4gJhuVT+3I4J4D35qHUTmLbIbm2r0Cma2f07E5HycO2LQK
U8UERfsQMs5MHrLY7Hs6p7oFuvFgmFh6Xt72UoIxxN6Ros8AL/9pBbeMMN907p15
2ZEtU6qSpWKUCL2N8/Qo/rsBADrk1pQyDveXJovjOrZnfA4dijlrycQeVDBHFfsi
0lTDuG48HJIiFQdOU1axVWYCzveXMuOKo/MIrgZhwq4foVHkx9sK+7+Th9FXfxAq
nNwlnw1jllf+Y9vHXsXVa3aCABgfTs7tIpdhUc53elKRJKfeY/PI+T++TabJZq+B
8GF0mEOlU5etVv50YrqkSXLXkq+PThbrVXotsttxgz7Kr42gTLT49S/Gzk0qllzX
0m2KHe+fA82K5k70V6SijEwTmUOoE/v3uFbRNNWntlBfGrdSnWCXYTQ8FQdw0aOn
ku7W8KRJNlHVkYrJPPRyECd1+apRHB5cf7Zl85Od7VYgh5jWzOCZSEUhdpoKubjy
tnyxGAHXf7FwVkyZIPCgC2cacnjbsqP82+A6khq3qEh1O6Vh712p6vMis1FStMnT
3YOnwcfTNOhULHRYis93gyKUT8ABEp+OYCQqn8+SQseNTVuWNhlRDkAOtewusCWE
IRHVvwxWhTZM9w7RlcGiAakTk9CWqcP8L2TwMl1/yRC2HUNq3tAmGYpXMDW9Ca6O
dDQuFq5YP2MV5Tr2tm6o5S5McMuIjCLqZIfMrdlABd7RbywXsASA8sowPdefPnqP
x3r/PgVeBMKucg5BY6ykWp6YLELuc+dksQronzN6ovBQKdPv5i4hpL+Ue3CrGmq/
MKBBM1V76wm8jvG/jCJgpSlgolgjeYr+/6RYyTGyCdf6u5qdw4/pFZpxDck07fUw
Yz7bKv+rv5jP8WrgNJLYeHZtkp12s0nJHER57d4r3ruryw7H2SBN/lTlVRnowQL6
3bGCEkjYStxQNb8v6iJZw867N5RY4B+M8inUVlp3FKsMxAi0MMbmfX2si15lBsQx
6gjk1n1mqEGzgtke+1VtQSREy/K794gOIfs40muqegqvlT2QR10KGgfBCG+tmCL0
AjLg8Iq8lNccq0U6FfypNf6InvNFhMP+WPCKKh8ppY90ZQ8uFhzNCO43yrDBK6g3
TDkfTxcvHJc5RGO5ZWq0G/GyqchblnwybvLdopyqZN+QyDtgk+Wgyr/Tgu1E2vGP
Xvy97DtOUwmvuWlBYWiCnMq4ebHpGb2QfhMzbTms4RM0jYu/awvKqAjQg0SWAwRB
ad8vpPiBxTXIecJcsbkehcgmbyPfLnqv7PchPGOxajIjvzlpy9Ex5BQT04GXu53L
1Caja/xia/EkcGFKRAuaK/UW+GUrJ2RPVrLaxOqF9i1aVUIeF6FXfi0mlOSrJz3q
DwMJWsXdWt9rgTNaHBbvavesiFQU59ayl/6RVft7Uy/ZJUcw07C6CtrjvDF+q6P5
ifeAnyzLwAlljoD9fAoyzuIvd6RqaYApAk6nyE2fy2bBwMQSJRGbLHB/ofSlOH6O
tZo8+lthuQnUitwaAFFnpcbC2zn7Uk294P/OGn3A1QbjCD/Y6LoFmrfPJVS7cSBI
wfFZ1HnGljpBk2Frtw7ZhNunwxPprCb+Tqr4lm5RoJTtmA1szam5qsXL/Vwh3SgX
bvOvWb8csgHvseEA3bphid5NrfY4m10ZdF9bxJB1C2JH7QBloPLaUrkqBer4jfQH
zZbpCGSyyWdj/rHVbDAiM0bIi8+iQaZCg5fKFaHOWQOTuKrhtAsyA+/PfoTjkxZ8
P/bVtrdPBC8l32EpTe28OApX9J2Xj3rc75FbZx7EVBggSHhVzCK6+R9CFdPZOgjL
3OTvRolnX1G7UWxvFqwoUAPxhZ1DbrdbnN+ZDdN3O4JqfyGXo4WPe4Jis839Ahpt
MCc+pLE5rYF7a70vdtfnnoXwLPZ8ieLmxDtDiTHtRZO5BQ5dagskVK0Pve3+TD4e
8RUYrviSEBWQK2ddCqoD2XqxD/slUaSwjth0kDimSXa1uWo+KyKZt+aFTQfKjYlY
DkZOlHLs8822LwWo2taGeufnq4Xe9LbkWvxXcS5Yd2j2hxYuyTIkCGrtPdwPD0Ou
FvRBhEw2ZYQzd5ywz6Qm8lyAy5c/aTy0Zl/8hunQ5/Qv7ZkgtD8gLl7m5EHPN0rZ
q5Wtb6ToyxnVADUIn5i/fR3Ur0rPPwhWp7jnwv9xl+mdEmxDjm8osJSXltD5K+K8
6oAfMVRyJ95ul+ZlIDclidzisd8FAiBtjNWBFJVCcMGg/5n+EvkcNukPRFUgAQA1
HD4HZN+CgSmZiZAlF85ai2s/S6Kv4NT1fEExkPw3V1s2ZlsfqVejrGdijGXfp6mE
4HWojfwPcmIu/rdL9N0rUZoyg66IZ42hJ05equefqdO0rW0zv5l6YqLeqSOI9snp
gH0yfP/JmuYYePg3WcglchuLD1xiZGalrR4sK/50kCZrHZ5wb5pndmby+UKtcCpr
i9VVr3sNgA1B1bNdc2c26FV/kvM2PlkmfpfggTDKoFPba/61EG+qonxeM/iuV/XK
QV8IoPaQ5/SbwWwQKbBa5ZMZQgYcqRKgTnfyQMQyOPcQ+TNi+IIMK8sBv3kcmMoo
gGM8m4Q9uM7JrUDgKf/hcmG+zkdgPjQae1aDdnxncxSNnZM14UkGCbcaXNkOkg+q
hPsIgUqTFpcd35K4H8cvYVAzBhhs62JfFXP3u+Jeb1rtjrGSHhwUftCBt1/R1rw7
KnQpS79MW3uIzC7Ha4IREeue6oZpO85KJt5H/a8pgo3a9UJcT/EAfNxewvjQeO6W
lJZAjgiK3G/IQha+8nlPUPolpcaYZYZjT+hgxypnC6taXEkUg/J4DLP/NH8grZ2U
9uDCAkFiVxcHgjFOHIrDPk0J0BeWWJr1sYUmaUN/Kobs81G255s5VaSl7tFXvhXw
5lgsEgToXiHDbKZpFXqHlki/ylb1SzHQEjsP07AsEOgJENWaXXW0pX/k8KyPXbyo
Qo9aXngJ04Bx6qjjGzJVA4KDxDGoOtKl8T+Il2NiDRg456yI6VwWEAOuuqwH4vS0
Lc/+1rQ+F2rBeON/4/QnVhJmdnzi7e2OUSJ4xCUy8RAnDBUVEHd6IqdhCiNUhd3i
DqhC7NHEV7b4YV3qUlglqGLbKzlLAD7lBkDC6+5FtRcEH/ffLblPyYC2QLy78ul2
MUcMF8rcqngNZ6/FzVpeMUHgdObrbVNr8vfLev6ubQ+GFuzJeGjFTNol6NYpXOK7
4KugNHgsh7Y2z4p3/I5r5GH5fFVRaZ6UOlGRBnOSGVgBGhL172DpOFb388yImbDe
kQl1jZIQXPFuyXrXtJ7oNJPpPyyxytybHL+gFFmpobTX/tgne6N+gh3VM1qj1seN
PWjYLlJJcqQFkix5GUMZHXR3vnqT47rBdP8xm+PaZwP/rNQbFVexqT4Q7PdOUqju
fQRIY2Z/XakneZMl32zQ46mW+N565RJpx0DFVBUlRE8Eop2CX2s/0dQ9CVX3JxTy
QbQy3D7bu3RqaUOz24hk7pFN/V3jLTq5AFBWuNomxXjc3o3jKMGGIFwHjtYPsQJa
HH0nxEZJM84RyQE1FDztwlcA8WE7dEqnfWw2P++VrG1HYF3PlxaZtOILabTgUxfI
c3SNTMBAhP7SCX2RQXTnX9i3qfSKpq43OlRGtg4ODDje38fomjvQkYYbIqN1AnwC
IpnxXbVWgG3/7v8UFTDGbnvLirpjsLwnFyPw2Qy3I7n01oQ2MH5H+XSzclWoP6nn
XPpSeRpVNtMVFSJOZZk5Nv64B1qoSuhhfgLbtU70hhxku5Bfw5GiSBxYXZP3CWp6
QrqkCfN5BPNkm/L/PsLo4Tvo7VHV10arPVkXAY82oYT2gXIvs8+/P85Io0/zoJrL
FydPXZ17JkjfrzO34/Ck5UlxCmMgFp7Pxal7ui9RtiGBS6vcuW19Oo+dcizEpWYO
xM3SNMWSU3NhYtYkU46XD5WKJDBdbsWHgE0Ra8F3vf7fWkQGyHBy2en23jcHWut2
zhxIQhi1NpyvdeH4m9COrxQfhUwUEDN8zv/vzTuTCPkxo+x4bybq5hVRdvKqALOg
xVn6fmJMm8EDld3ck4DtlZPzlpgZoKZDSfXAyByHa0kXea7BZCPHU4e1Pv4axjDW
xq8A6vXmb2zAEBlWFnsRGGispeHJzw2K4Igd9axEmioBXlZcE9+T+V9sGuUQ3gyD
5vhwWgAm8AdYbDcUVSl8qCk8MsbpD+57BwMhzy9z0/BuRW+SuJwJKA+YGmy4n1D6
ad0i5HP8EAVyDO9KKxheJLmeo4XPLoak5q/NDEnkGoDPDAfACl1IwU0h4emDkbHJ
U/xgHNUey/vFhadbITboHk0Be2+WQCu8xB565CW/ZGRmWCESXCGTX1gW8odn5g2M
8Je8BhRUA6V/7j7cQARINq0OP36sg8VViCeZdz170dXXvad7xVxC1a+VgQIlMbj1
CmUu+WbrmTvPTFEYKRgiv0s0zQBYrYgJqxUEE1bElb+++sPF5B+g31SMZgOEuHJC
fbKdjZfY5VcO3DV/Bb3mcnGsgg1cCaNpxjw0wUJ6bxOZenNTOJGPeyOXfHyZJt9a
/hOK/7VKD0SGHmft9Il/CXlHLSvL2cBg5ZZ8hJtFU+/MpW+E+eCBKsYeHwjiDBSv
zaXi9JBQig5Fn1cToyt3MeTZtwHjCiOu8xpb9ALDxPlfQx8DuEoS2o1xZXr3BoWe
bEWFnstKrya6IJZmLTaeuSxYNq2Rrgy6Q3WMVVIo+ZENuOJJEfPxbslZBcQPc9hn
+DJfP6q/RHtjMGnN8HOA7yDb2lQ9gi3rywAbdhx2MQ9zi3kf2HI9H4l8+C6WhA3b
obPwdKaYpoehP45nQJ+gNzkCFdiVpn+YtxMm4cEKM32bJ2JO0hV3tWHLlVnX4G7O
OT8lTXEQ9elxkD+4ZWjxUb2WJaInlv8/rWSkrq32GJnlEv1auytkjVCiJBCqOYwO
ddSHCixZnGYFO+ztxgg1/z/C6wMlHwGxqH+3qUIFiDoIc0AVdwDpI146nvv+5Xtg
sYA1J+fWmrHBv6vik9WrDQS2FZE7AKfKouL9IeuJUDGcMsTCXbX6LaPDsvFxsEri
6XaG8h6rTsN3gBJCBtuWiiTEkj865tMUGgYaAMEvv6eFhvdMu/vFvaqmtX6ZZLzX
JLVl9KJtObMsdxnP8TZQlshOmasuaSLaKRTCc4oYWiOD0YUyNwY9S+8ERhkou56U
EPGxiQ8HFFwa6cpOrEuczg04Pzgiq2DiK8jjA/oXrGmLVvR0O/OFMjNq/GwtGB+T
xawVy5dxWsB2kKgOwoS+lkirSUYHcMVBMlHMMdIsQ5iSXGbqEfEdffPVE/yMOIqm
7CUqAnTNY9MyshC3E76H5HVI0M3vDBejHfSlA9hEXHbvPElmcH6EOopM+2DiTiu6
G2t8y1akU2L4OochN4KmwJH5UQSOTGMMwMLKKMtUf29Jl6jWxB1pxviPJ6TV73WZ
aEjNLq13SOTe6mblxjOrquqy/CiwOyhQfycU0b4FTPEZofKyAbHJNNpSmRlJOw2I
hnChb7TY+MOK4JAlWAPJX8VKBUt27QZVsWzehHf9SzQT9PEjNr3XLI+/5XdTRydy
zpbFa/XmVWPh7kZcNgxbSW1UQl73UPYoTi3iseWlF6TVLoyPk+YoCWcFq/C5TB0M
9E/TM5OqPxpSuRzxCzK8MdkOptPcGUgYXsFGbh+qIarBwQcjCXcHbhzwBv2CBcKW
T3lkFXOu7guafUEzHl5cFfl1dWQseAZO4SC+BGtZb8MOVVRo+CbPWl8dILezixxq
opWcxfCR2/acfOdjJ2bZ9fQ0S/x6nnzufWl+wNuHZN1QzEqV+U6jOf7ypV4gD2Gt
Jfj6L8xcf4Vs7LPAlZMwkZplDQmtw9y7qfrQg3xeNSLvXKm50uHPl1BFFqwBndKc
ialLvsphKWKDwr0utCh+9GWHZOAvJdCLOtUs1YF8TGjBM8fdcaA8AWqjFcfqxu0J
nzOytoftcwmrR+8sP91Bc+/5/x7Im7bSq5rGqF4GizQS78mYbAyzp0lCL+0q5v5f
SKbukvPLgDp284F3hpD5ycyzp8BZuEFKLdyWvXrHkJHzdL9fM34LOa/LD3nUGwXy
oUnNOlWkdh/Y39JK/xY2HMC37+MbOqhGuJOWD/snZVZhnLFPajoT6xKIlJFR2rxc
C39BUkux2+S5iZP0KkgB4rZwA31XZoMOGNMPKTD0Kw+4tS/3HDIz5GXSLtw0gXB7
VRhwDUQ6TYt/2ymkUXHg8lJKr8GCf7IeAIwyiRNkpwj7R4m8xbv/WB1jTkSiEdQM
jZTVYV0HGsLyS6904ZZGzwP5GbC7Rr/Vp0aBwSOqetJ8A1tXXQWC1D9/uRdyBCNi
eTxmrvTlXSFE7dZgD48rwKFDCYCuvOkntWgaHdNsdA6q2xoWhZspEPBFvM3GqDuf
ERfC9XambI+I4YjnSOfbmIQDtCGSEg0QbuHXpQ42Kat8aK/1tVdKo9ABiRwqIIP7
nqEdCJGx7S0I96oEem9rfOxeukOW6Itv8+d8yhQ7F/SkUCwMcqxCQtdCrYbT1lrS
KICahT8w5+NMrJ8uHgL6HhqqfVZ7Qri6fL4hDZIgNlVPYHhTDFZ4LUyLxEzmnhiZ
odbEVcLTuscOwzP+jNBkbkJG+a4TTaGejjxy6IV7+V1XWsct7yQfJcd0KegYb8l+
mfH4xTJFE0R9sgvVsZ2ENFduxuQPiow1aTbMvXNYBnCCX7VmEGPJUI6yZhR8ufyi
E4fjqdi9iMkS6hFIiZfzODwlhPG8cuLwUdiOIz3OauAErbEG3QIKEaZtqZZJbyEx
6Ry1kzc1pR2+AlrqRxR/RXGhCVsW3+b9w6VrQfio+myC/KMZkM5fFtJLLxrqC2Ob
wLQlPVzqina/RuZipcJr+Pmtbul6XWxEVicZI/urBDCDQAGapu4d1Nm5xTU6R9Qd
i0VdRbZHx8Xrz4Aq/11x9RUe/bqdMTR+Sj2Tn5wFIgekCEzk11q5HNZ8xwSWTPbW
5bVjDJM3w5Jkp8mQtfyl/RajBSRcVLr6GxoXS0KUn/tdrgqwnu9WTdxHhlFtX9bn
b1bEPUTTzcYc9grbcZegQ2DJr7cm9HyCHJxLNrHHM2b7EFhDbPy3EIWuVkDUYdqC
sRr/eI+0GDgCcB2OwCLjZY06lpem0KQ4ZZU+BLBwdju1CqXv0bY8wLHVLdX/ZCv3
j/cufR7YVhu3roE41ViHQmusKAyyI6K2/xJTYrf5WN3UIskAolRYBSKS7h/5I3q1
to83qwqg/oPidEbGXYN9JBIxS8te6umKyOInS7EmEUVt6vZ6ozxdrUHFB4mwxNpr
j/+6EdPcEMOxBwtETsab2RZ26/wB5oZTXmxVHTI0VkSF8EuFPe7QeXa1kkdS7hs/
faHKX01ueoTF8l5CiR96fHIwskqiWSHmtJpas6oGjvg1fuZ7Ha13JTws5alnVGc1
zEQ+En864zkiK60RqEvKCYxK5A+4XwkHRnKB4bACCesgR11RWXWhocDxzp8Rc7Mr
XDiOyilExe+i2BpAyLuVQ0UJfzLaVcekHLRSpwYiH1NoZrrT3wq85p/lqNOxg/Le
OkY0CgYbT4ihHpHPRJRfUK05CGR7XtvyQtquoRclCQD/DN03B5QEVyuM3j1XNm4W
4oV6fdfVdaodb4n2wUdTsSAGGWtXS9pVRkPsAorOFKgaiXliX3tFKs6zvvqRDgSs
7LWVWbYaTJlsgnBhLhF+YKzgY90/1G55tA51a3sIVTkKx+zGE7E5LGoLMj5PhB3q
7KmadaHHtqLgV9OZxqsGTsOFet6Ur0uskEbMeS8xdNgZ+89IQOacYKgyXc88s5Hc
uYki+hVUSfV17sURNUvc3E6oaJKDUdYL+bahEYnO+44s797xYAZnA07GORzxdsxo
+Mo0jn58gV3zq3V6AGWNXpFCH9AqioZbB1s5oLBBtb2knaqV6KEHBA/FCsVq8F0n
KtG7gdJRxRcPeUOThlr4kJ0ie4/OfvfewUBA8WyDVjFms93mppNRyRJrps6U/UGD
UQNairkbBRDCpxW2ApBSnfksXdppyTbLmKhrHl2e6ftmPJs5aUTvRjKlDYE1HNWP
qer9xI6aODocZMn+N7sKV4PKjlG5nnqJxeh4fRvFvNL8S/4A2UJ8FQpWezq8FE5X
v3dB3gXh7HPB0+5g9cqO6QVKhZaETkTkn1XlI1wL7Hg1muigyBtHXnhVLj4BEmNu
m+RqPo1w1bYAv6pay5p67rQdx2K1LjF8ez7mNytyF6vPAhUsXN50Jaey6jZFVCU4
zNbtgmBxLIrDahfvQd7CfDWZjugSHEcg7LclA42gCqF10AKKLe522+EJYYiD9sbp
AS9UAO2EhljO40dksM2G1ZLzdl7Cnt3ro8DrvDNPFwDUDVgjSZZbqMAneTYpaKxG
Qn5fvlkFr9ALWB55qsAuMeAKSIpKQp7SDUn8MjZH+T064fV5as1R16QSQS9kzHB/
C12FNwB7Etmr5s9uWSh6Cw6DJUT0d5FGu/93pGFkNXIhHHOO49rSIvOwBWxFusJA
1/+ryDaXh1WFO7Bd65z0fYV3Zi9sDC7e2OpOuHKfzrNOgkTeTHlPB6JVEBHvuUkZ
GUBuvDmsdNw/WCz3/6mT+aD6Ka/y9cTSV4LVOnG4Hf4baYyneShT3jk9p9QfRAAh
ju9pliAIcjU5c6pY4PK/55HXbgXXN/S1g9cuavwqanCIQZYb1Wy+q4LTKdgQJmyL
xcJXN2wz/+dPZnfU4PH79VJXyNG+1Dg20/72mMy19QV3ZKV8S+hdWJHF5wjq74ly
zitiXc1ENqY2g3H6gMAR//5RaurD90mqFj54hORSBMAD3094uEJ4u5Xilrq4HKmo
gczVwQZ5GUfQorsn9JO3RW9yfE5pu6/QLvJA8AYnTrdwdSdMaGfvueb1n/V6XiI0
I6n5F0LxKo1ST/zYu10fESfI+DNXcwfAFAwkUils1WZqVlzhmhcgQD4Rls3HTlFz
eU62E9LgWhRBwwFu3q/GSJJKDshnXmvFUWDpOZv5MNJjESqpt7ZMZtPTnBP3XXNi
2fe6jgA3rn4QLOFeRV2EQmsHNIk82yYUtFso0cDQ1quCLfdk365fbyyOr1DJaKC9
0hcq9JEuWOc+JtdtXBQLO14gbLXx3qT7CJQeFsvJrcW+yAeibm6LqItUJTLNcmpX
ikaRX7PKpP4r/cPjtbjTel1V+vXV3juZJ3M/0ONIc1aoWqyyvRW2ctjNj/wg+GhR
TEA2WmCf8GbJ1WVzSJbDgcVM3nzmCx/RzyMpwFMVIodI5ldezXBUYgZP9L007hTh
xJgg0So7Yov2fKhIHEe2Zad/oaKHMY4OpLp0l0IwD4OyoT7qcHxT1J2R+QpuXv/6
9D4vtptMMC/AYHGwRU9lrJUnZt8T+SYGTCs+JAwuAgN1zfuo2FSiQNMC9j0Tg3Wm
DAB8fPfVajeCDM4weArMaqrOEFPxiLUGtkUZgbmJAB4TIbnxbrTekS6m50GPeSQS
EwK5C85tb9cs93Bqohrmh8Y8ad3gn2IyXLREJgnq+61NIc9NGT1pYN9KDuNtfJIB
wXfJtcY8nfWqcFCvAP1xROz+/rMtB99SGqB3FPje0i6eJh4Znsu1/A1pAu8wsUgR
/VSyaeQ8BYmY23qDXcfYL8OXZdk/wRz+oTE/R1MmVIDBXTetPEaFLGDLpdiYFK1V
gccwroEg/EsAGqdwcXUO6N8eTwEu0GNx9V/IZjBv7hkNpCXFuAk3+8NtaK6ZfU0+
4Fo5qe8jCz640wl+7VqDWAXP7nSRTRMhkQZHi9+cZTsdSr9zlTZ0Vf1z0To+AUnj
ClD2tldjsGRtx0ncXYRT89y2aOaUtyl2Ey/ZSztXL0V+FHE/J6FF/4hulm3fN/5Q
cuWNYty7hMNSj7PzXsbSonuNBRx4fFCZw6KOgaMzfu+Yv74kQNgSl/xS/hZyDnfK
aSodpPq1ADIOELKznMptI4CzzkqkiKz9WL7Bc4SiljlZoQFU3F+3kk6TLseOCo+W
wjj0VkTZLcBAtcNy5ZVpTIKJ5m0gLtGncMfJQRFduEBnK0QfTKoE0sYt4VrxJTR1
2Z9+NlVyB0CjNgpCVc8fx4GPLFrvsp/ya45/Bj21A4hBMF54JFZQsvXYPPJ6EGsV
ZftpEI7yNoX2kYNo9CHc8EZCesssca9I5Xovo3ZBF4CkTuPQwebp7aQ9h1cLFhPz
GlSQ9615dpV4P10Y7ZRkMOUarirV7bPfpE56CONIzDb40ISY+MuE9l4S388TwhTz
5B6Ghy1vh9PGEL5PYIRJhJZCf92YckwR5vAT1WXXAJ3n/YRU3d67Had8nOMcrP9k
S79lviI9pSmwQ5MRe0U5Zowi2A+PoTYAG2Y4vfkxTxD53zttseP5XSo8Z+zURzuy
awCw9X0ARKz3h3/N0q8VcXM2VE2KvgbJu54KDuEOhldGrYGBxR249xO42IAJMrnL
KRhRrF1hZeFLR9/xM/2aL4GoBALZUlCAjZhXQk9TsRsiWdnA/lmhq9BJw3J4aJu0
l2txvgr8LeRbkpb5bY+ufQGjsyQ7Gdq5R+FAfOWZWO84vwCNKuDcHB8bpTTZ8NDs
A00d8CIIPY+HP9d2IUmYNJHsg+WYah4gfaKtWiM+gmjjv2HEtput6CLPtQIRESYo
J0/fhvytnqUES9ZiiB1j1xEVYSr0Og1CkEv70h6aQBSIBjoBUlyvSZ66eYzAA4sl
pC4aPExvOcAzjo/sVyPREvJX+CYSmGgrW37yqHKvmlFg54Q5uAf2eIZysWcZlosb
kz9d9wLv4ylzARnvbC0/yno0fxvsITSh9htiCzbSKnKMSkXuQKOuXxkdlwDS05wc
S8DhYQXk9T+tE/0FTb7wOXuxxftqpWR5wXrjcWq1czwZfbVwA4SiomHBxj+QdXj2
unhe0hTsYUkQkqIbx0qhg3vLH1unQ+exzGA+4+0e9USCqNR2Pt1wspiDL1DV/xgV
1h4nVe7uNENhyjFCjkPxV6P3XNhAif3N8s82T2BwSkfElvdgNgI/7RBAhlrvM00I
t7I+eaXD5O1w/yokkYz4YxQ/JBcF5AuFEGhn+r5fsOiOlNO63NHGox+t2ArgRiIT
sly7mSmysfFwC3SGg/ES3nqbw0dha+u2j37E/Lt/H3IoAOiDoTovTnwdC8ACbkbg
TtRLjyN92yUQNWWW1aiS3i8g4zJ9cKxDegISUHZ8XRXy/L7NlqBAZBnMSy1alYu9
2psOUJdFDWToWJNSEEIn98lfS6vz7c5eaAO2ychpcbg0Ajc3zyemYDtwcRtctl/D
FO80YMixjTBjOLNtBSSJvIZ5UnNWntBbyr/Tni4oXilyaOMqOOYnQ2vIT0xbkR3W
uk0a8F4MQ8QSBRjCFStJmG8bELCQm/ctffGb5tU42ksInHmhXIeNztRppEYJwuiT
JI5QZXBPiEy9Y8rn0hTp8mm47RIwGdzK2Bsefu7tuAc1wjP+jyqdE/T6FaToE7CC
oco5CLiRUd7/zmVTo7CBsVkc7SoF2D+peO0Ih4c8omP+CQQE2ZBRUcYtf6AxgjkN
zc3owatM3QJBOWSHwLq3mvRxSSBy6sKUQShp4Tg7Z+Jp/IZvU3sYu5Gex823Qtfd
pDaUJQfa7T33HUyfR6iCzOpTwnNIXk4WQeBciT3u8wU8nE8HxQqeX52FysoWw9T9
p8ADYUeHuZZHNQh7nupPPMfH31JsL2zwKPjTvI4obwCbG1dN2m/7mtkkRhL9HVED
Er18p6uX9IqZp1PU+c6aCB4HYnursmQuhP+OLeLJbBy93Of35d9oajBoem2QzAxR
JIy14LfvyGPPGYCAaQXUDB5XrM5V2CBVYk98T4RWBUHxPV3EtIy5iOalGbtYvWfA
PRKGtxx6ZXhFZghDZ2dlj8ApVp/EGV4Tr05IdKhvsM5Iq7wsh2gGZfFR6OipLh4W
9b/JHpu0FpcIzU9ZPNyYMytN9B5Q8sNjCRwBg263KFdxyP7w0/QrugM5F6Tx4bv0
JAlz/aBz2F02IR2tUxeSZ0L4hSfu/vJkST73hC7VYq2pQTjZLiVkBGRP+M5phMcL
jOl91FZ28TnVfF3mjNWPnH4ULhdfmdGY4kNguPdr+U74LYhiyGvGsrplNs47lDU+
nr2tK7WuCNx1yH/kEKbfQAmQfVpCon0tOhDIjDbRvOKZq3w1yRYUw9AM4C7jg74K
tQi412WoN6X1g2nW+jdqyePBZmeWad9WcYuzDkiSJJNHyEoHNjmTu+ZelOK2R3gW
A0Rs3L48Jo3/lrvicZqNgTfQ1HMvJmjLTkmMzyW4I8aUt1cleKvpTplJRDfaVcGG
/N/CXYe2rSSniyfWEjdPxuPSG841Csbhb05870S1ZfZIo3Ce4L9xlu14y4Zq7p7R
BZOvAc1OWggBbrTP9GAsKXbuamnKupyMFOA/sC1ToKtRvP96jZH7vrCUqSX80Md/
xXDsV6YVeyXa8o5pCy7f6EPNQR3vgpuObaFLR46oDKMXMLO34oa7BQ/vpBOPjscJ
HMEiDmtC8k8lwt9nZab2szbxFWlIC11rXFrqKzgDEaslT6SjYPbGisyKj5XbhRBW
Rkb7x6eQcfDJOtg/rNQRVE7WUFofc9VTUQVbDiTZvE2hp21ZCcd8m3ovr0UOPJXp
odE8ksYead2Df51Rxlowutmrp2GUSFZTUuQUUp+SPRid52Q5JlEd6o9nshfq5nkV
fEJx4UhjKKxQmaTnckbpm/DGCrTlJ9G3rAL3s30QoRS6jV0yZgBFakVAF2J3r6WC
CyFPZXn/ohy2b/xoaAvJd/NgCZw10Tyn3AZmYM1eJ/0oZkVhXYJ9nYl4Y2ezAc73
6mOtXVTkLa/TA7iCJhmDwzb1HuInSe1T0keNcjRuCHe3lq0MKs8EkTI21u7Rp2yQ
da76m9uY8dNlrBtXRUEDau5QsnUQd2+iPtYJx+m5GiISKCoOsGU11RX8aWo3BvmO
PrL43ZoIHT7+f/F4CLD9nQG0Uo5SUwrlRKCiah0Zm1QvEbbh0z78OAijR0s00PoA
DI7fun0n0t/YRVurb7j/17P0WucAJqmj5hR9BGRwFo6BhMJ/Fb0NwXJLQks8k0rM
6rc99zJ4qftVTD8nsLUlY/ilCwqrNWRMs9Io8L89bevG/+KsULfKJ22SFk2rrK6U
jbCQtqYQG4XPQs8WDVBA9UDjHr4oKYC7Ub8+PET34G85GS5C0P+NMKLvndbYk6eI
qJtwjq+wS7+ILZ6lIZZy1eh+eSNsRBL+Z6KvyVMwRoxhP7l5q7TaxgR+vL5dovra
lx7QQbAKpIVy8hRsbv0ucrDAS+2B5PnwAJ2nhAgCByac1d6SGm/AhZwvKkvROrMY
bRVelbT7azg2CCjHEFsFZO9QNFnW/U627Jh6LL3h4lHWZctQ5tAi/ovBTBVsg69z
HmLwGupIgdMM0Mk76AdbKFqrFzCoMBF5Jz1rzdEIvLuqvhmndv+6yNmO34jb+LJt
wXqHGY8NuTHOHcrwrEqCydkz7opwlUDedDyjeo83tPEWDvyd5Yk4ZZzUR5GkoUqg
Nxx5osNQ+OoUnpUCHXJ9GhxtYWUSA28B0w4AWZ7U2P3Gohi8r6aiH0z6vxRtrSMm
8N5IespoAYfocQGZuynFx5TlDR/6NTUK9i5XqRh8SNHTjxVRxqhZ+OI8UYvcDvjt
c//EFHXGj3WVVqpzAkLazhrD/ul3XC4V5F4Eixx3ryv/5gsmJBBX1jsJJo6wnTxy
OHlxBtDwtK6dL8SYXeog5yvOdhYUaVfNWVMM7jKNqrsI8SpqcMdLnsnagMjFaolj
EFYmJeAqhEYIth3PoJNET/8aYaMwhORIUlCs5iNZi9mXS2dIOq5soyeCewhJkss0
crGPsqNyIFbxzdwXN+De2q439PVWHp9DCFdKm4/6qbcxhFCGEfFkvC3CB1oaBi9v
LR1DluMrgpcmDifybCQCjdOrhjIPzjsaLU5xJjycf4ZeUQlm9lJfbJkSyXBAG0io
Tfop4pBkFxqE4EpzgiwUtn5lYMWmBlOTn63B915U9s3LBbocfeDFkephMWGnHVnq
mpL+DalFTL0R4jqme0WQZXxbRxUkWY6bTD/OB4He2rP9OKJ1zi3/Ltio3gB61Hnr
UOvqaaLM7jWL7buq8lH+CYvI6yWn125pQDmM1inCUdFfzMRQSTw+dwKEgpbfnQc7
9jK/yngZSXTkRiwtHgldfy4MiEjvH5o8MqOEBBhFZlsXsI+5zXiGWE5t09L3IPZw
FPTS78Z2hYbr1kJjwlu8hCW90mDqDCIk9MTZzmDIf9aNCIhn2qO9zGX3MBq+OWup
mMNltRPf92XqXTsLk+nzP9kcnzjYRG1jYs9aiW+tOJ6a8GWmcPFQkqaqvMNWIuRr
suMyGEnU8x2oxeuX0GZqIiu944mNUMPk0+TH9Pdy9yc8VaATPSAbZpqbR7R0/Kxa
NUGCBzCqZ/MH/U3r4Im5B0jNTz+wy+nW+4nzS8GWMfc8CE44kA+REzGfAU32rXU8
8o9ZZpNVIONH86C2OvBXHDLs/lgOb7R6uV1uRWo88klNhWUyLEYdEkcGBhSnwJV5
yUBDAorfSxNbrZmcMECAq4Wzs1VDf/I1q99Rw4eOjl48c2DKDLw7k8w4rcq6ibt8
cqlKloNSpAywWvtewTuGFdqdnZbz52gHe7MUDOeqQxQA3dv+X4foZzfynBzkcZW6
6drwgDgSCNbIvj8dBvM0Amuv5EHxgifi3YwTozWQro4IuVEWXVXWu0xwVUBriEUs
TlzFYxiWIJ4VOj3lVFhfcqYveQgbgkdYA96M45lYZZ8r5Eye2gRQAY6SKgBLEpbV
Vb34hkMynqAIF3D5bP+MZnhmo5oS3O+MXHYdMeEdMItFumERlktyWqZAX7i3X3KO
VK2kCcis+q0i8E2dxal2sxXAx4hIj8tOimoHmqIjwqKIRZzKeht22zSIYuGzyYDW
sstbXD5f3HqLM/I+6mVgFlA0or7ITe4vcCrC5ezdvVhIpOizGM9bk3DKFzcsaJFN
40JnZOZSQFnqEXPFJ0vmFfUtoBpH7ryoybxi6KUYZwbX/VI/PKj0E4uZPq3nhsZ5
EswSrbty1titQIxELujAk7qf1HxOWxBjSSV9enuLtymtJbiDZHgdJazXMdJDoH78
0zFr53cJZGOOBdDporBSOIg0SyEeTfpNpautlNEuvY2xqlXwOc3CNAQXNslxm0r5
UdmqeeMmYO55HIKl7ZYSJIpur/QQ5BbH4zEVCh2OFFXtc2HjrXp2rCmX0ZPsv/PW
H5bTdedx3L7udwQVzB30hGvU4DtCTXvpOmERMDFx6zm4guujdoeTZFiNrdFQgyQu
VGVr++k3EJx6LHVYWznaaa1cdYIphKOg1mnmEbbDbs/o25CWhEf0PnDqj9Xz0eSI
xwXCW2x0rUCbaXHzyJK0hZGa/nkalhjuqip77wqIlubXQnytF9sBKGwIj98+pu8W
Y24YQR+sBYjkL2eWKVeCtS1eXBXKB28WZYz00EshAhqFL4f2nA9Mw32Xht9vunkZ
UmNcu1ebVAjiCNDjThKrpwJs30cY99ipjB6Pm7MNJGt94FSPd0LwS0aFzVeGg+fF
TBJZykkkE/iy9OzAeK41kZw7Bs0iobj8aifLSc2NxtG0lYWveKGKGvQCApdV32uX
eM2S5jV2CKjNKzMQGWXrGZjiZVQrHrYcnrmmSAm9yS63bbk70DpyX/hlKRJ9PjYQ
15LVb9MuSEAu7ohcZSbY+gvPDGToMIgaWgsrD2REF8OXnesoM6Z/F6NydbS77Urr
lmY+5d+Q+ayuVZ7jqbPEhWV7LFZAagpKosyEWd2R7CQgIB552tDhhWQKzlNxDauO
X7+od5xNbnyu1sEz4OZndswiivrXXM9mS270hMtSxNu57oa16137sa3b+iHaC3/K
aX4KXobJEEF5u4GFtVkLfqxIOfD3kn6Zq2+u8HHbkUWvo8Z1o1yheySmok7p4XHJ
ItuDm30gUZ7QPt0KkXES+iDDZGl38nRrySItL9peDM/mco9gg0IRqrVvajvbANSB
SfcL2ClZ15qWiWkns0bTkxj6AAcbff9JdbfHiFNZkgsru78R5aGnZvjUAPWtWFx+
1EAjmIYE/Lo87hgThXlJvyjGOKSu0mAkqm02KXcbc2t6TzjdUTQwtfDhzCcgGman
V9WwMmgFhV1rfDzcKbmQOvUMawPyuXQOpu33BXdlpxM3OCJuJgmaGVAuEvQbVdQO
NWiSrj4L5ztHdxdaHUMhXQ7yabZuEvv926dKsQ+uXNM0NoIBXWnBz1toRAcn2nwy
AEn4ENE60tekXkKrkO9iYpo8OErkK0XlC3SbT7ReRVmurbHI39OxQcP3ZEANIL9E
iAQDReFRNPZyhlcEs/KiS2Sl7AcpWqO1VcJgXalIUFa7Wb/pli3Pjkws1qh710ko
mDEGwJWbL2HspWucsueAMs+83D8KSGZ2alI+poUsBVDnvAnuSY0xr9A1I0POu+l4
MIQw0bogDh6Igg4sd4xCIl0bz2ljX2zg8AnzLNIIogHzfMNz1c4AAKEP2hXZ6dmR
8RSWR4PT50hpeoPBq2VgTJEpB5vQp3HmCJr9jL2K+LC4oW1TQpCi53CHPcW6zGpB
QAcXiK/dMnGMSVdA2SdonVS2o4V1KZR8SU3jyo3DJki7T0+xsPewi9hqonB0uuj0
ELqVN00KTiuem7R7eanVaXWaKQb8r11dEzQMT06PKXnJgDTNJ6paRpXDuhkfwbMY
ego5E55D5tdBMyb4m42ID5mnp2OTwsIlHokSemuPQlF2fWXvLjjjgr/cQ01n1REe
YLUc1RQDVARf2zMuRsQvnu2r30uaio/H6aqlPfcTbMjyoLslFnNX/X4kwP5KoID+
FrrRPqB2flOlWes7EuA4qW2CglrjRzK+H9FuNGge826BMf0B2QCXaNSyoBeEMiV8
zZrncaPwCiPPnDdbtK4F9P3VjMKTHGtSjez4W5jYCsbT8etJlcwAHFcHuwsxn9+B
sl3A7NBkGJjUHRaUMnxZdQG7qPxNXb6JWbhrPFYOfS3UlubPlZaCiayJlrkof4j/
HKbQ3U/vAl/f0xsKjt5/FmX1pLTUOospU36bkdhi/TFfD0tTtXY0LL8dsOsfmBG9
9R2muv+lsS5ZpAEA8RiqLG5Uh0kT4mX6YazHC+GSM/VGuuGkhCGOC1AEfaWxnRjW
BaKaTazpEvGcg+biPWoxMHm+Kxaq16I3+pp/4/e4htKzpJiDJv36dJ7LqP7Y7KPA
bfe30O999xpn4I8yVdT6mPagquBG0bHm8gbhJN6SctthsNN6lKmycHd7bu9kTWt8
YFRX1hSR9PBxpN7Phkm2YmDE6AkJa8qL+zbEhAiZYyRwQlb+1e/IfSiHTwWGiXGk
sc/SaO8lEaucXDNg1Q4pRfltcbuZraMjwWNYb+eiE+bxrWQmVLWSaHeFNgVbkEdV
OCtzRZynl8fmSp3alMXvSQZYBfxT+OSlDGVT+ece9w6yaPPjI5T268UTlfZAMFGz
8gvPyCGUH/mDgsOuqsK+9zpCGyA6d8HarKgcQQ3u8V2b7AwR/Oqhp+6mu3Ta+DAZ
C+7RpjZV0NDohzJzc1AT1qo6/cyeUKX3Nm4w9vC2om1KgHutebj8FuNwRqasXYPg
il7TJdSgQRTTCOa2xXa679+kEUgyDCSZKPjkB5c/drbJhIdlkzH074k2CkbZrRHJ
q1Oox3kn15IXaENE2i8ifai4EqztrxKf6e+J6VeWIrKAWNdTKIIeHqCChMYxkN3E
ZKANR7aeEDpp0f2q1b+tf0HjsUclyOxG2X1rR5bW5dBhRDk6zFn+ml/G6nye3UZG
/RpqZwHOwnXl6+rVyQHD23VC8dlunL2btAhPdvwsE3m7UATtjKKJ6vbxnVcjVvzt
/TO+1/WWwBUiZRHvS6K/z3iNCZf9dG3dqVkCaW6IHosPKuZQt9y5qRBbzAZ+cRLH
5gNM+9g/ORoxE8DReUjHC72Q+gj9On8NAQPuMDZr2SpxwdRXwk1INU7H91Vrfnu+
+K1VrH8cO+kzAzcDC3u5mVK58Skh8CR2oHjywusQYENf1MGP5od+spOQ4AsJjDQ5
/ynRg3lZ1hCwh6lF8f9vcyy2/VgJOYM22VSSncjF0ySko9+iNaJ8GCQz++ubeP41
UxIaOQTGG8woThhlwYgq9lOBzZ8UHdDjnoFohYHo2/0GjCwzgLeUaLb/sXbDa68b
cVfMBk17NNhML8rltNf0v/jNiIEhWc3qGjWLWeinf0w7Ak6eqV5rHpiYEifcq0Ff
xtOtPVdJJn+N3L2svfK5zJ/yLeryeH1JfS8pmHcSequlEyw1nRGlsXnTvl/OEVjw
xwfE2Vc6kvU8DULsHrDK8/xymzEFR6wdKbq+6rWCCPSx4St+dYLcawZnbehLcvUQ
HB3cCvlLpJdPPgB1Cg2hl4n8OzQ7UIV7OoxVl7pGxgAXKTFOnx3Zd4V1bpmygE2c
YB04md8bM4JGjLPYrneFpxEkegIpXqpdUTYSaPtoCu6Z2fdJLG7J7kaqflkW37w2
aj8Bpb+Bn6M/6Taajpbf8nTyfGpROANQ7autVb/sPHyDz5yzKDUhObz1uUpoHHsE
0zxpnaMGkoFwdhS1bHXTZgmCCF/sF+ANP72kb5kwjzYj8pkg/CQe7qt3lGy3ZTGF
9pUA5jf3ECeq3w743bLT1c3VmDthmHVawahdSqo3ANNSJWvn6UVK8rnqgrW7wjv8
ZF8jIBh1yyTrxVk6iFnCZrA1KwtruWFgC3lfy8pdl/gXxY3rTw4rCov6ZV3xn0Cn
`pragma protect end_protected
