// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kjVjd2Y8c26cO/BcbhX2fnzK8AJS12RNAEbElFJYbMQdxkqnN/eBIFN3vCLzp/8h
i4mRmFkZTL/jyX2UTw47sfVBEEj/+xYFGyEG1s+dz0AXWBFsCBnmL6aGpg0+/YKs
U0or4aL0NCWu0WhJQxfW92DpB0QfmGkoD9XrKZC4xKg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7120)
7S7a5qqJwD/Swr+zGZeYqfKZYCvgGJiTZMwvx86XA+FScTgP+GYuopFbOd+gpxi6
sMAsdsU5wv3xBqbd/RPOuDd0g0r2E5J8pqg2xX6TccmcA1TjSe/7tE5t1eGRc85g
NNZIXZfg2C9b+Y667FPeSpYOvA8FcBCUog/THQ+jWDtrT+zSWnezdK+Wx1h98a6G
QkB2TVNTYqcu/RW15VnQKJwCis8FSGibzJggNuiHnFjR+AddHccI7qbPgjLRDBgO
RZ2e+ubY359C4Rb9aAG1R+4YuPV7DkNb9IftTizqgGXVP+V45BGXDbzqMpU7kjbB
QTa3LvdeyhkH2SJ/8DOJz+bX9pZuBwDY7xUe2A2OifhLyrjgsaK+iHhcHaHdv1Ih
C6UvXN5ei61rQ+Yx2/H7eXggwdenreWYfqkWTfIEA3F7LNExV1ATb7xePjvGqM5X
nwvrD+g11iJlgvy2bpzUiZwXO+UBL5WhwsJs/Nk0kmRJk6cfKxV3Fmi1SfV/x+f8
tdKPuuQA5BOW4rIf8RRIMWOZOTj3GSVvQGBQr7nIO0pbKj1qdUJ0XrzlCaA77oYZ
E0ezoF8IA8YXsmNnENdtFuaD27nPXgTmakFpXPwk9+H4hd/Fm7wAuC4uul51UjIh
HJ5BUf5QCp1zzdslfoemnctfKXnaj+aseOv4DKtJyOWLffQGvjM3Sev8oNxtQ2X7
PqyvqX4WY6u/Ht7jO/WI2lW1IM+sTJIURKzUSTv1ZFOGuXoGxBTZs7c5rGYtDHLF
wJJyLu99lCg4Zrw+IkXkQ/2R/5V3HGGb78bwqNiIOUE35Ly9MdvvczrhO5KlxJ2h
H9+XNd6bCWfSKsozaslm2Jv5kmC2aCzpd1Y2w4Xqf9nfPMTq1SfYZLzzQP0uWiwi
T2/p2L0zhZbRX8ElbNH2gJJ0G3bGSzR3fQCBa29Hi7BpJU3LeREop8wBQC1lXC/r
6s1VvwrawY4tj7O5T/qR0uzuHtjTNEEMha6SzPSxSjCFlFcj/sKjuq2v9PlfBEsw
AAvzo+NUqQRkj347rb3aeKppY/jsV09I7HEidVPgPI28vIv7lPP2vrY5yslWEnLb
0IBiLgxxlOQv5MsFKUuOCTV0ngM0VdgQw3chFLuGQwvjlP3Xx1dc+OvPGs7JwXtE
UxvYdtoj3Iby1839eSYU3A9IdaL4NcHBYS1xCsEqmz7dY1opmqaYgT5SWY3YpfzW
Ia7CDOuEL1irqWbywleVs43NWN9GZ3A11Z68ap6uPKFPDhcAm5ABrgIuH3uuh/Wr
Ew2VyGObiSOS3NrvibKGuF7UPk60vpTpIBSy5B3M6qIppwS5Al9+qxpBg5d/uiQd
0oK1Sa8LrWiQ0OHLq/PGSuWjUpXMSaJ2d79xVctpdjz2DCiNWBOJGlCY6iZ7yxgn
3XqGq0oWrf2slZ34qaxbeUoaGJae+kTTMD7xT2rHztBmWHpKn6zS9/tPVwv7JQlA
0tRiuz1MzMDjQd72cG9Tz6FyOBYbXjXvdMtWqxpnSqPKX7uf7ueLf6sigC2kdR/j
e+kuH5TUjV6CV70ZF/CSwq163EGREYpoDow60cpmABnM6smKN09qA17HLCH4bDyO
P+a4A8v0C4rTndDIfv+duyUujfDhNZsal1tjGUReWWnS0CmeTEAI4X93S5+HP3Rs
VJmlG2icjVmNcnxSUrfF+J48y73HOeTWRpwoATGoAR+BF8M+iYD4vzOyaKNbsrx9
tlPbRtAgIwwSMcyN1Ne6SRNYbPbqJNDmKnZhCdtIGLwpJsOznKGSD8BcFAdhRxbV
wIGP3dZVWz39St+W96+eGBXXmX7lV4kY3XecxpfTqxinZXQPbwsetDy4Zt/we9fu
wa0cbsr5iAKILg5FesAGJPOfZxZ4RFj7Ui7Wb6ilCJMQVhKHrcvWGf7ibkPsIyvp
yH1KwTyCqsWA4anLu5Zk6fJ7yaYHEQVGOguzNhF/akpMdy2msmMY4GSy/gSO3bmX
PITedK3/de8AxUDUJ+F9hoPtNRpSpKEaI+n1ZoO49WKvjCKHdwDruVrphekGL8as
Io3X/4Xb+WA+PaT1dLFgTtTh4fixcqai6FyS0ufndPgVMN3Y8VMZkTYWiNxOBw/w
YgEa70v0B4ERDfmCgob9KjF7drbdk+NbjWeSG8a6/aE7EOBkgNhSIkZdaQtZKyiI
GNUPPFEFieGAKFgKLM46jLm93v6kEDVrrOxjpBaxX2qiRhiQv6THT0cttDqmKop/
oW39d8+6bDyf20nWmj8caS7YN3o2VQYG9cLkI0R6vn8XGlYnFg7noTNZkOaDpTYn
3Zw5ymuOAostSciW3IDDyvXJCy+PoTKioQGGlEyICwv1eq2L2kGrFnD0PrYVCIEV
wDAuGMsm2Ofb++SLX2iMGMGEqn2O1zbioLq6Mcrnp3QeQ+c1pFRlqvuEFf9EUXuf
ZWjfluQMsuEWqqrc2OyJPvvockUtuNxDTeCmwyS6Jh0y+SaA3qAGcD0N0/8CjMzD
0iab1g1jAIfy/q4nnTYxSacGLZNxn+VcDMqJ2qe3C6VZEd1elKQ6FLiNAuj7wIeU
cE4iUtOM17oBuV3BDsuMP2P8eCj9vZ85vHQI8kgbN+bSyVng8Wrek09qHW8WSwV7
XoRSmARpvwquhusLCYKpqfcCToCraA85a66v/LV3YSBiRqOAo8HUlBpzeSnGCwIo
5HrHFh0LH6czjSp3iovidfhX+vrgz1Hi8GpNqPGmk+Ip5w8rWLskqlXfL3Zc9uWr
IHsNvvDDLwN6p+f4P9bCJV1sNCVW5ATQgvTM1LDkSxrhf5P5YnyIqE58ELC6kgHo
buXgp/RSJVquasBtFDONqb3eMdc3chNl/z+S9fEYJTUXTXYGqggaZZWMOM78uSMh
cQCtkW6XD8eiqjyDmbUZR17H3dSU6SMWwnfHV1/gt7LbRURT5E5onQOabe1fnBVT
++Ca/APNHCzbbQSJeQIw1XEzjF3yg3W8L4vNAj88XL/th4XHzZ3u1BhY1PTXKdok
sMHkNfshiy3Mv73g37BTSa3DQcvDKwkLjE2rL88Kv067SQkD3H6oGRasZb/MrJLQ
yH7y4bTIhbzXMwJjmQ0AehygSRCPVtCkhfC9IlaXLNlZ4+NfuhWXCFEH50OYMpih
YuRBFz4ItkkczgducNoM+6oZz4Gx2brV/2TL2eaJAQp68B1K+Mx9+ugXCofURgm2
EtAD1xUt7pcz0hy05xijYHd1esVQPYCcj9yRvA8XIz46J3yZkM0sTdvAapjLVe6u
215X83w8OGMGxQ7Ux5S3N5hqZTUrOpIhiR5Z1wnZIIzfRm9GbJ5U3nHCGs7a+KB6
/49vk7QmmUmUePeOAvQyC4ImFw4XQ8PLJomrRP1SIld70/eXzJ3D9qwPbrM6IEBa
9VYptqAU2jZOTAU/0rMsqWR2fXISFv+L2TmrCaQYWcEOsdr3d4F3tJqojHqG2bUo
RXfG1vOylFZJO9lDVdoQ1BzDwNTsa3GjmGFgRw2vz+nu40XVmJRZoI2VtXdaPksB
E3HEEwVgLdJyDNTv6R/kQQLlVyJTgnvPvkmZYGPqqHA0wnOTGEOn7cMslOvBsr5O
Nn89gjuXYHUisOX/GEprcu6Az/gvA2lu6WggR9nZBW1L446FlSvTUMGxNkGs9eHc
v+rM3FFFVieVXG4xRWHPfxUqK6Ru0uvE9OkRfO8EEzXZwmBuzlW9XDG8yF8ZcpOr
POqMBy4FUMEfe9lvpr4G00TRvVUbhjxqSgTv6RPS+bLDG3E9hMSnGeqFyZ99OBbH
yOWHUVK70MzjgAnqrFMpzniLKzx52h60SZXLqV2pT73uNxPR9hd+hT4Be+43I8VK
szFnvjNWqKktID+bV5asqISQRFIvjXvRyPwSJ3DbFWqEcW7xZXN13oNkPkrvKbWJ
m+hgl8wPm8twEkXdZeM6HBzmQeRpVsTPUG5NtZsAi24UFRAlkPEDvk8eYgXty65J
JEL1/famghVei+60tEo3QPU4iQSPEU41vCr+aTlmhjhsAs7Q9gStpkpJR+FmLY+r
MVvcmcGZXTZzP6dNYTQpxCuPd3VDdpjxtcetu1ysgT2fgO9cNTmiouV1/3MWZFZQ
5TuiLhtNevGySRoJ15mCTd4Z8vHjmjWqqE0rz4WRRvMIYpUpigRwLqDWVRtSwLcm
bpBqcf6qg19gggH8kmr+kx2YzSGJxsGBqWQ48xlGBVdcAIocv63aoeD1iL4dZieq
/zHjBXR+KmyxzYCcdqN+nOt2mpIRQMFSZSl5bPx0ar4ilsmqCIHpc0dn0Iuo/pof
Dc7ZwE1FzCAhORlzsWqiauvdhDR6rqeH6i1nt2ZCEUJ2Bzykc72A6wcqcv2UE12o
rPEvHl6biay4Rv0I4bMoaMPdx5EoMIeER9lQpSmwkORZvOfmYamHIayXWYKkXrGi
tDff3Ae8dHhHo+Es9gL+jB5wEDzbJZpWMd/S7XxjF0n/mMMb9uEpiJL7peOGGSn0
7u77VZ8rtq30AD9i81ffMbHLVR3/d6/NnmTVJ226mIycQ4MObuQA2JV3IfpUJNzs
F/zcNvhGqnprWoF7qrJL6AiuKxcS/Wfwn7vVQQGnWE431NdJalvHpStiO4Ar+Ejm
XexFmVD5ZaEAvgxVLAc48ux8THoMV2CNvMxmq0aIjzLfCNqkzbJS6V7scAWEs6b+
SqzpmSXHBu9VRL7uQKE2uFmWpimLpKxsFzRmXvzrJQ3oovzWXGbHQPLwItzEwGTH
XggefRkocq/P03V/4ITDC8i+IAFHtm6nbz7mI5DxFlpVW6WS+fkDorUbJQSz/wTu
9RO3AVYdMIXZKCMjkb7BLDU9w+Xsop7W2xPlaG9/GiAbOyPOed+Jpzy2OMwoLKCR
N5GJSXDYDcgFLg0/TL2eJYcHRgSBZGOsPy4tw80ZUljDBG90dVMF91LwQfgPQV2U
oyxX4ftntHd2pUnnkgLd4LVOUVLPYgyDM9yCnCPcToVeNudrXC/7o/Rh45f3y9dJ
8Ub6SnkHg9GWT+sdKBwt4g0RMRJw5aqnBN2ciQKDlbaOcBgq5cvgn5Lucyb2thkX
1vOG2HwoZr70Z27gOIjRLwHxotCDZPQSoE/7Mstz00oggwQQuWaoLqYdpzi9vgAS
qY/uZKg54qxd6v2Y0/kavSumoijhIO7EvS/kIPu10cdzMm+qG45FimuwlseRunRX
eoP8acuxWUVgnxGYH/QKPMRh1A6MTnz6vDyXyJ+D0zVzJ+dm/40OoqNsUQcU7fOi
CB/xr1FGnOb95ndv7xz+h5alJQgsajm6nvGPTwzVpclVBNn/EvTk+Sz0jpXJ7gb7
uY9NuuWLkYqiPPG8IuC5x4QLBwYhRekl8GhsdMfWvB2fTHEpTOnn2XTIEsLojdnq
IhZiU/bf4ymA5eRVE7awhKTg8ynk5oKCB1nMoIJtTxh+wa38gjsO1Kegmjjx/GJk
FeB5cQ9hioDW8vxiu06XMyzqK4zvzQPQb0hKqQjsPjvkskkVu/uIY07iUoqeOapE
fUBE2qHvg8S2XnJisf8ayH6z6rYGgf+fCT3UTCGD65couV1iVJXP9woJZ/+0AlLM
xQePiLKJLUfepZkdrxL7BvVMI/9aTI6bSTXhWsrvB+xmR/w0U7HrlQqBOY0tK5jg
+zrhSuxWZ+o2KwJcJQ/VqmQ26Ye7ZSPtWNfjl58RdHi5SxBI3UpnpsugeNv0e47P
vg5RhUGSghffGEJFl3s1hDSUpXwAw0VezhWTByKFivmwoEdttkxeOtAebHqBIls2
sXKSQ+4aPV9pnwrsYz1nfy9jzHgkQk+r+EJuHx1rxntlyKozZGdPy8QusiK+3gPr
M0BEbgS1567Nv5uBqknoVmlIC2fX30PJq6pHvVPu1E23c3TyZlvWDkmxhT8FeAn/
J54pB58yU3RmdQ2C8vo7izOjsxZ1DPK1IaLMGgaAeq2EYrfiZQfPGQAdGyZxz379
bVzxIZYnRfch2RqvCq2b1jlx1mbVhXEuZGQDjlUbzvjpIXXPUajZUOzBBJNy6Bep
KLyiYqQML0bkQe7x/ZqDMsmlYB8cWhnOXO+CCXcSYmtC3pp3Qib6Pfm4NE86Vapr
jLNtb+fFMkS4kFTRIN6eBxg4gI9K7DQQhdwh7H310ZOeJm1jtWnDVnEoX0RyKCZv
tOKFGQM5PPEsccOG+kpkQv0c0WObGQ1ANL8NkRDUOXvgfM+L6+2EXgynmV0M0xP3
hUopsSKTJXXT9ts8c9BX/dfOkAcdMOPPWZuD2mzDiGFXYUeeQmZHJqzakCgAcaL1
KrwcQ133rKPxEc7fAlkWhjjJlNybU9uTmriGgkIW7X3jn+2F/mxKuXP2QuKc6h30
NmSU1asDJR6aSxdcxWS6fhJMY/n0L2WG/h7Hx2xTkExWnZBHJ8upJbGzWgAC/WBO
JUWyPHd/a4VTPf9/olWCgQnGbxOqBE/RhjFvcXjvpWAOUyt6RxxflJdDuDTSYNiY
+LpM6pOvSFh4GeZooe9XI1Q2SLgvwb7rxDSfkiXXrlZEoVtKzk+3PQDt/DdrKBFZ
8IS71OY7BlVVyVQrP+o8WF+eOzZ/vUF/Pkd9BuB7xRhGfNezbDwGxsfS0oJa4Rnh
PC1dT4KCMlMfX0OFCzy6lxBtxxzPbIEvSf3+nt/GKfi08Oygs9esLsNOy51dD5ra
k6cc6BGst26tr45YqncfgLFKvrtVlNKxEIbOUJlbbJ4HC8ir92cYGxB1SyNDCuEg
Pyoc9oicKnzu+1xd9SyWTfDNZEHXapZ1A3x7YB0o9SYVdzKjnRJTx1qjQEc14DJK
VSYgfY/hONC3pxP1ryEvVXEbfxvGgUIj5p2Oo34B8DnUftUaWmw2Tst67da2IrBz
jc2Uu1aZkRoxdtqCmPMLqgAXU2jyXOFeILjy/pRyIdKUyMtpOXrKyxTcB8lufGqw
gbPtI8OTh1HkFLYNlCppdtqZMG0YcDFgFV3lSUpbu9O4NlU36n2DOpcQ6BWfeyBY
UmRV9dyt0UGbg+3Nql6h8At+jUVCqkGU+2nGGEVvlKqX8cVjSckV7ujZ940Oohxh
7hewcO7csC2A66gw1cjqv3SfIQkJXHGs+5kOZ6LvChHj7uVAmWWFFsc7YzDKF6ry
NdVoi9cYHuxGTnoYc10ozzmX8gt5SSnxGXG8SWibXslXldZVDA0FG+tqdK6yy1mo
Rv2pqyt0WNr2edA9G43Yz2MIy5z5JYIS+lQfV6VAgW0xuqze9kOEr4hRuOXiO9r3
R4z7y59Wjd8x7Mmy9736X3jCtx6uwdemmSC/W4GSGgKU1tvZ20p5Oa3MYfJHb71M
jV3L6x1NQ2HEaecqo4f5XP51OGsNK8KHbaVVWxBW3JIwG8Vpt24FvHqlCcMjwOc5
4SrM1BhR8+4d0Kak/85V6V7PvQuHHhUCnfGyddF+unFh9TPLJbOCYH4uA2NowBF5
wk359+w3X7/P1V2h4+jZDzfRbOWz3+hIpzJu+dPhmppyrxZcX4+5OiongdJNk0Gu
VnYksxk6d+UGnUxvrdKrfGRNkciJphc6SByAcnzmVUU0Frxr/nYYM+mqZzU74sdv
vJ1Q1TUS28yGIUkWnErqC/qZXn/l7qSzPtGPTqaGo0T3p8ujEn0vJOFFeHrHg/Ky
G9d7qTvBhsEAvMDLmomdk16GHiGHeOv4E3GpAf4ZQj8zv4PhWQfJEr/BeDCXvZ6Z
w3OaIsuZbOOwZvCakmxPYMUNJFjaWyTnbqj5m0TtyZifXIaYeED33GAJpszi619v
EuEfPOSVTKeSidiaWdgNTvLSrvU7nwXAfNLdR8W7+vALGe4R9VTKW4L1Ric15jeb
2cFX6f6SBDrOG81Jw+gmqOGNPJRp9xI+D60o9tBEiJKcd488O1asYqVXlyl5v6hq
LM6vZWsehBq2AKv8MPQJWPpudQI7Gds3t+j6jZ4PrrmBSaqbg7IX0MYXkva9sdkG
HajKPSLLxbEurrVOxE7YscKG7Awe8kyTdW2xXwGKmD8OTSQLTCCXctG0CiDHpBaK
q3opjFosprWwZzGjSpehx9+OAslyvP0hzhaF5TmAPq08fEzYjJGWflwY/Jq4tFRL
4nuzf+Wom1k0qTssW7xc/BrE/Aob0fQM/5bFZ/aitFBp6kgQPnF2wc/0stUx8R//
aCNZtpssO2zph4ocAxklabs2jZk2JX9GSo+JVvU9EdnX6V+smqLuIRNaQKxWGDGU
C4C0vC1gyXHeAudVQgfq3Q4/iIm7jA8efg5lhpuRes9l+ri1ODw20M2brOYR/LQR
EmYwPM11WkMOrVj12ePze3USzEwdpj6IpH/2fmllca2WY2Ujtr860PHJ7XBx7LSJ
WNDe6d91anw8InxHkzGMyl7S4X3WkawxOlpaMYJIoVo5AZNpPQBi5gy0mKvB+H0M
6TeGC+bGXImY6NM5H2olzihkVPSaeeC2wjt5dMl5Yx6NwNeWkMexb4p95EQa7ijN
LYhgsIM8R1L/zJUh+pl1a66hkbysLQ3Ks9tQNY1hPrKTJ5bVKvbRZexUwu0KzXxq
PEi6sCr4ZZHTRV6xhsQ4jNInSZBhAOc//4Uev5a56AhNInpLJm9xt8Biv2DCJ9xl
xnn9cv1MvwJNLdUV6rpPp/paKFfoP2vdm4dk72d3l4jnpdc+qgvLvBJ+sWzQ1Zfx
QkSm5W784zLDEEnaWTP5YQh0IqH4W14kZmHOX2YaopAdMDQcEePaMJOizCiWpeZF
yo7ylo0kdPjOIGvRjnrky4rh23Sm7HfmvFACb1VaVHDYugsZJXvKv62Av/OOwq12
sDQJdSFndBQ8UWSYyboANE/EHyKc6qZwRt6vLxwnH+e5USGoJ76/bpNpyDPviWV0
K9VWAx4KDIlak8/+NxaTyAVNz5aD9fBtOaWs+3VFEyvtAjjx53IqU5/+OMRCuy5f
9/se6lZAaaQms3uBFHktJUar46E47pCy3URnNEfZcnZzB1qiKhzlnjy1kGdBBFFk
csXQg4dQ5OpNFL8GoqrRB+Qk2O3TKfcnRbdSrYLN6PfQA3mX2KBvPXBXiWcJmGlU
Vl5rrLsGwgi9ZscnyQ8LU598OFDjgDJslOcGmGxKZMx8JK5bGd8phO2jdPUvMtk9
mW2fjd5A9b8HRCyJF6QNcAb/qDatVgk888IaSAGiPWGUSG0KRDPKVm8Cok87Esk5
o8Q5RoHqoDTm+2fUfKnRyhLlsc53+IakcOMhhuzR+czt+SSoqu/pdJV8U1mrUE5/
ff+EPw+eza4ShwrX1tOKZmM5LyoaI+unca2gBg4FRnuzQBTlrfhEIC45cA/3Ge1L
GrFkBtY+AR3WWhEMuGpyKGYfe0ivbDfWI1Pm46vgpT6apAo87q7ym6LMbEZhYmFD
S+N14Urfy+sI9xBVVFRgytu6xET3/+UNMHb3X+9ozEYzp/zh3cEOtfdtXZ5zjXkG
nNtmfw+d/p0OHJ1MtrI2+42M2fmgiMmjh7EyMSIQuBTrPTfxHmhMC3VjmjC7McX3
Q8RPzeX9vHvMfibS7IzJig==
`pragma protect end_protected
