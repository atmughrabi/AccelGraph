// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XnuP2Eurx0ca8eIPjCP9CyrolHnk80jafZbVVxO8LXPx5gRaW2oNf5Pph0fiT11j
6WbA4HBoewJajQElOCe/Bv2/62nLrYRBhcDqkuJKbh/3jQpQnLcoy9AhlNOYD5Px
lUXw1xmImnu0cTvmgnN4Kp/w6qJiLS8pgcL5T2mjyiA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21232)
msbpVmXoRM+InG5dgLDgE7qwHDVpIAt7jhW81/eDU5pa03tr8pIwP7nJFHnBWOXa
vdVZM65cJdgiL565WYdC3MXG0oKtgGgJp/CW9v/RWr1Pj/7HtEMhm1iMW2SdQuRd
QKxmKKPPbg0Lxyw9k59wriMbj9AXBdoxpAGC6fDPOyc4jeva8F/NFvssklTqSeBG
7/TxTi0o1Gz5vnSBy8Nt79yYPCtepFh7RvKy9QlHSzl+eAsZMvbuUExkR+4jSZBS
uOC6r4J3b0CeHG/rml8wSnailAw2/f/YBLc521Q4cVAxjYB7AAxqLKreBgCc3ZHN
cZL52ZVxUPpVe9YgSpteyLfmQEk+i0UKmW7k0BqQx7CBfrhetZPm44Nc8uW3S3Ma
OevyeHwCFM12+POF2OVOf1Pn/SCuZe5hQ+izT7BvK14qdEL5Is1/mKYdMUdgpkph
NxQJgB8oVIAJWiwQBkF+bV0uZ5AlV/bhRhQDU2dj7YNrdRluAe62rQM0snZBf+4p
AN/Fui6mHuwBDAa+RVVBBXff2J+mbRT3WxYR2CYyMwFlZpJs5yThOkIwuuoF50sP
n7BtkOjdTjnCR54llmf8tZJRcrmGJ5FoU/hooMeve7xpRtID/UNHebj7x9hrHzD4
cDZLCUE3ERBOJo/+jz/uXEJYDAAAU9rDovVybbUcybUCXsEKtg92QNoT+VieLcoJ
52FQNkyW/HmdHGmIpVoCjhqpGopK5Qx/DVwoeAemfQ0RyLbglKzuV17jo1S3rSIS
aoQ8VksUkF8WuLHcfuBT0sBwDo4eMOziv9QjVQNhNFBqMV5blkgvrOdUSpYB2PVv
RJg7oViBN9O5SZ5GBsgiYYPdQlM2+L23SEJOl8Oe/MLAVRSkp6nwGczbU9OlXDDV
MsOm1nxlIw8EUtmtf3sLi+R4AsIdA0XOrT2PKL04YT9tzQBH2Am9RrOjKXiuXsQI
GFWqlvGi8Dy5mTtMQLRCuDQWy39irRhy6MGPlTyjlw5h6/oA4xkeX8XZQtayikXY
+0mbJibzuETjG4fdw568IOpSQs89Og92MXaJlmDJB4aT3qnCk5XomSOL5h+bckvd
al9rA2livOQDpcFYB9TnAvBbnvxxTUPBSdIX+iraJBX/PqHfHCT6Ft16Z8lvoQbL
b6zW1B/LuEuwkAi14B956LwVyZ95tQ1Z5tCmPywLhr9DrYOt+hHREIxhjzn5KUW5
ZrnHIVXDho4wLo7orN7jqMIX8kTiVPV4FKjUOGKU05Th5rkXHttggxX4gCAnsOQc
S9BE14PTW5wvSsR7SUBRSsiY5H3N0tGrrxodnU66XumrkHGXcTkV6qv3lcNLp5tK
3rSmpqdb7vmk1n0/H3gFSor+fPONVuG7nIEwbVjwKa4MuHQu562Y7wresj+aEnh+
BRJVT5oeLLvmubwhni2xdv18lZX9qEAyGpoxj/CBCPl0M9VIuz4fj3wJJfNY5zUY
z81mzEZ6hRfiOjv29VoFfG0QhKYp2urieYaNZwR2PFsytR8ff8FFXtECKj7hs4q3
9dOxUv9jk30pBt2AV7/E8+qYIMoSI0FI6OdeSIBWfSTQFfhOJeRNaGhl574jZWRO
+7iLuGbBwjdcfwTDxpyWdaQJYhf87/THmJJryUZnU1ndaJaQqMYXDWUwB1xyCvtQ
wmVWBHx49vbZWSdZTJv4mbM7htlLkdQejY8f2Q6FSVF0DZZgZP59xuvZvy72kw8x
pq2YHbZZBq9c90t1+E84jZDcNn8vjuQeLbcchpZtOv7VOpaXvTOfw/xXy4qGjtuI
uMJ8L/NQMcWvgiJK6Zhg+q8bIqEOcun+oPYPIqtOtBkVuP4I8GiXoHZDlx/o/v8p
hVm9Z8awVZQNF4ohN8ezYCUeZiNX2/Wt/GOBY5bGQVelztomEpFrAaeJGlNtYAY3
7+4U1gw+FHuShvadOBcNaLEwTLiYDrj3dTdZDYqpr/Ua1/aV3+t/7Gp6AmuaBvus
/F94oaC5XDMSbpKZjwSJqaDENOVuZopiwY5VzdxLKLYFnmbTmOyG2yB7RHGRoztG
r866FBQjcDYxdJescQUIRX37LqPhkd5cSZdAhhhMgdsbP6aVWyw7XnYQ0Gbo8Mnn
pX3n4IzdmccBTunbt0HDwSOTMndriR/zEqba2glupTCrUyTOBC5ZBSqGTed0HykS
K5oHR97p13lzoZc6R+QWg2QVS55nKoayZkkeWE75WdFTo5zzkoNg6frbugr/mKc5
1YWVpDO5Oxf3GbrJJyuAGnBRqc7Vr07NRyHELBdkBwRhXzmJZeK5xMSMnQnn4oMC
L9avOfIl7a/EOKbhr8lmKyU1spOaV3LHGYvivDZfjgXpDVgXsjlFXmF9skkqJrFN
7QSI9ioQJLEZgfj5f+fOEay3NZTo+8zfCIg4c2orWHiCiOd1UAr62YffLx3rl8ky
77m3oxV8RyEhDXtMdqIJGlb3FNd1NIeMSF0izu9+ELLfRXRn/ybTyOPp2f+lA/TS
RCzy01lDK4bJ0RhDcFocjWLQzKF9IVxzxQzwBrXKY/pBcxfwtxdwokeFQlk+yvfy
UbX3wGg9OnAq0PzDmiCYOvQe1a5g0i/0HD1uZLnalrch/2wus92FmoHtIiEXkNJm
h+BaqmtjKd+kdM56LhyUFGUfauUVGXdYI5+W++0dmaGdVoTSAZcMEfnZGsSrI/xA
9j41mrs4CgiL9Sf2NQlJto4XoMy8z5tKqqV1/6zV7YnyUcEe3j0jSeqBn+ryt2ai
fCjYUXSIYocn6KsvcVIrygnJb1+GzKorRz3la0i5XlaCfagijyMNU6swXYut3aUK
3fccgJA4dCePpEgaTDC/7WH8igAyjCfmiVb/VnKx9czcTMkcB+hPAkJaJwGfirHC
TPJ7mcZMlkIl2YrY7nWrfq9ZfH0Uzp/DntHZ8IsLLlh5ULbZkJ6DUJLMoUn0TcUH
jAywiBEpXqAg9M3xG2LzgTX3IG0JCecaacT4lyJjD7whjIRubtSfxDYkPagSAPYH
lrDjOMp8QSpPKrur0DUBPgJWiaV31X+WTa2iNG+v0EJTjHw7vMawwOwDreo3zSZs
VVz9ap97OP5PnZjM0YmDra1s4d/8CzTfeedaMm51q1cy/i6iP5vlTVM5/nnfXspV
j1wvq5+1LKlZQauJePL+p9Xq8kuRfQU1n1FE7qL+TjGnIdkW7Tiy9yr0TRZvxZBQ
OQ+dLe9s/7a1wQ9SCyaF4ahIy5nIawfaoKwXCpl9TvaYB42UoHLX7Lw40knJ3Sro
jATstPBg2cURl1UEo1qXzZ39xrhFPSIQoDtL0ns1Lpup3O/aW4o78XBq0Vk1YcX3
QbUCqg8mEHSftSPaYmJv5dKWZTNxrsdW+VzGyXKicARXSFpzJkRrKhngG2XSG1ae
u+gZzQ3P2ZQYEQeltNVjFI6HlMO1XSuTn0bsQ1EIIkyote3Hw9OWusg4mgHhV5v2
Ol/7R8azc4tYvn2xfx2WgW35nzylkKrdgf0hDwzV1LE1Rpsenu72Zf+MNGZgEMC0
6GAcpL9y+wHF/oCoRloCLpYdWuWIYyuomi+ePWIPzN+WhrujOFC+5xDnUAYKeHuc
J/mTFWabllq1KbdaywsO7rth5hTKZ+B/1PIm+lVRgDwX2miXq0U3nd6VXgx9rUwF
WtO2OsxNzxoBmdbxCUxcinSv8ArFMgQbJCW4GIG8Tl3uO6xMZ65cKaow4CGR2EFi
Iaxor4q6SXS7GRiATEAUpavPWH4ez8HNc7Mjgj0I54RYy3s/KUD3vHQ5ntgU5HjS
oGuY0zZ4GqzxGlEC4xOgWYMIy2zaF25Nuro3we1dUvt+buf4HJ1JH9S4sBqsj7Xu
3JAifeKnriHy+J7CvVavv6Z1v4afcdBm80+dsL1ZAP5lhnCZsolTKd1Z/xuc5b2t
4Gk9vn7oN0MJ0yq8rh4TZUvJm62dzMydVmsZz5l75d8UGNm+fraG3Huj4DR/zNmI
FTNclKr5a9n8Uf5FVxqf3mGqT1OmQTyRRwrUp9Ve6cdZBzziZ4jaNRv/vL8FSP1X
mppUYMVMFQSYpRZbZ2SnZ9lUo/loQRYM3PPNc7m+cW13rOf7g5bHOF+AiFuXzRtJ
Q4hk+tw2ZhK5ZmvvCUF2U4Dz1to/MM9F2JgkZ2YzTrSQa9V8Ck9fHYGV3WPRrJzM
KhsMHRTe2vTL8CgxDUXSVJLHk0C0PsAxbD51NkfR3oY0DFiZoULjC9yedY3WCkpi
G56i2eQj+09OAdS9iBYUP19oIFd6uPT+ZwdanM8kdXblBMyioU2sDNm/ZCdBFUU8
emhjKLYRqHPuMDOWfmsd6Z/ZD1ChFcxVzlaL+PGqu51ecx5YEUBOfIoiSOzBqd+i
RQ+VOUooeVV5txbg9aq8c0PHtlD7PIn63dqo4grkJiEzG/OeEuYJaVhnNpuA5FUt
sFWoAPFMVQTM4R+4R/UVZbIngKGYBewCGEIjqzxvyDLNKQzqioeXCS7LZXO3jCPB
aQWaMSiBu0WZIV4tejxfsPK7+HT7PxzAqWNAD2hELTVeF+uZ8ssM8K8DZXzyylju
SBYeNYfD7RfL9tD3iwgwdJPIbIgO0eeLKzWLjrpCE3qJO4SizjeIis/FS8NWahCh
57n5RBrN4DiBupctNdP1QFUp6JwGRBYJCdOkckkw/y2yK7puRHNwQjR8zTV+tYnm
H6+arbZQjX1lBl9H0KoglnfvhnLjpXzmJFm+F3wpBMoy44l4TNnNcOJTUdsIHR/d
TGKnX4PGmZtz0exjKJazVLVH0CClUNJlM0IxFxP0wgRqcfHNIXZQYd/dY1zXRvPH
p6ribBqJkZez6ZrP9f6As+RoUMYNsDRnPYoO+6zpsS3OfSzulimrCPNjOSX0cCBT
BAMrfE/TxmgDxgnfHSKeSC8tgVoOe1UDzXLQYzpV7qGq5G2wKZPSeqV1J4nN7KZb
vQXYe0KgSvxdafKAEleSqyfCp0kJAlth6hrzskJ6cuzgauac0Cy85Lj2i7EyR7XK
Gs2XdFpj04gQIOuGKcofRSfHe4TXE5LH1ZT1YOPsFCXA/F+QIaR6PBc50x8np4zE
tuuAIG+kxWidhK75Pw4qzcNGfQa8MDWP4+mjznxrPHa70Ed6yOcLRTIuCTwK0fgU
rGSguLQMEavM/OcA+xq9azZitCf4JtOPcvLwe+hUjTRoIUls9ig8GnhKVe05jjul
5L/Cc18dEe9lSpPyi1h0gy6n/0ZBFe6E5GcQzY8umw28nenkJcKO1gxnRRJEyRg3
Xk770PFMgucESLju7JVFCI5L6aItSWziGsiyBuiW3XhnvqsxMeR3SACfcSYc3Vek
a+KS09AKq2kvaJ3sGhSFhA+2vJ5wDsL6ugSKEwalLhOmgtMzC+v9oZD5xeHqI0ZK
N/c0TghI08hRaBkyO5p6VHgmHT70SGn++DhnYoKgwrl4J8Pw33TVNPZrcr0pHdRJ
sbgt0/VbPR3wBsYDmOjuA+NGegN74YVyZFkOmuFddbSkGKI9ypyqXuAZ7/N+9Qlk
zvlKdTjhzf3kEvsldzyeq6eONZcI4vxFEiHVbeC+xtbcEuZ06qZrcQnRqYjEqU5p
hbiPqp7fTZWx3v5ctVWSwlSns5FNKpzVuoHN2k0EM5hvoU7l79cnrbtYKb3SlIEs
GkRH9sWfilyQL7Jq8TKwQLX4u2EQyVHGo8W+GJRLuzYwKfn1U1JiDCI4+4nXsh3J
0o8vGkLjYvYkL+jcbHRbNWv4YRKPLku+ri8LZW3vDng6LdrUijgLnQWlRNHAnGoF
2ASC83LNyQgrhg+pP8DeduEQ0BS9OZWvaJqFcFj9taqhfIgESxXa50XqZkkDIDel
V9QYqq7hGep3mZ25MChqVFisS3J9JwLY76xYKTXFfbo8MVtYUJhb76JijtfH1jrA
wtu2MperJxjIko8BYXMV/cw6vdIUfIWtBnv6DTBbFKF0CozQv2DCotYdhYsIXjQX
psrDGfpM9BjV4eYzsVmihk5q3dL7ycasjd03JvNFOPUzET3r6scajYWrvIucJ5ec
BDa1hpR8aB0xghI8wlq4eKxT/QfHPkxrIu5GNRDLXx1Xs7IlrthjR5QFgkv7ApBc
MVlz00xkBet0VUJcW2BaURndwmIifr01DYVtX31F/M8yauqZJDsDrHrATHyXXLfR
3GKH7w53gDcqAGTryodhsWgG9j62/DWVevKhdVOyorvLX0vJW91TkP0AUuOO1pCl
cHNUJ4BITYqAlBgmKuff2+CnjNKmSocUfh1S8YG6ejIZ2soiCWbf+bL73Bb2DpiP
xhliC4CzWjMWypH9V+C6HCkDhzTiNamwr9lHmq1ckosk/TJjU7p8KQaVCghw83d4
EB2E7UrGRnuoZdQcjdqlOCnzuoLLGqBJ7hgC/YPlsGxENfdxpFzG15OJP836Me3Q
xA4e17dRcBOjoxd8bUI5JyOmGeNV6jGvPqg3It/7mdkir7yEZMkA4NxPeCmaeSvc
XDEYHTu4Yf4G4Rn7ujF2jHzmOxbT1GNt/8bnDpoJmfFP6oHTJiE/aBgLv8Une7hh
5DLA+qfyRTVVKfsaJ253iq1/Tv6lmhWhUUHZNOJ0WkHnc5F/ACPEX3ltG1qeARk2
TGThKHKkBY9BRAI/DVMn7zeEIXCW4BIZ4BLEK5WffHB2rK1kb0IhEqR2GuO8vnqo
DVI1w3zd+//DhCCMuPSHheehK9D088A9gHZA6wtGw3vakmlDkbn4Cqza4SSG81WF
gSt81MROP+5M2xDo64lRt5cJ87UFNn33g6JjZE7su8PVvlRxo5Gy7EBc3sDsZF8O
QbDjmrkSkQCfCoeTvENNW69mPzGORByvdClgEj0DfJbVrIJHImznuzEOb0UhCOCr
dF6I3CwNS5tYTD+u71i2eAZ5CGF5wy86vuZ2RlgbT9AovmbZvOjwenDLsVbyJcMI
8ZrHH34/sJHAtDBdqgAfYEGCEd/7/0US5VdEWh8/Oae2J84ws7Ix0aD/UAWR0Wt9
eqqouyVXTb+Hn8yJ23rOlV5eD5EzFES20XOC1PVMclY3dTNAtgCRFmEbbAImQaV+
Y6bCVopk8stmYardZfukm/tkfJqxSkAYQ1e9S9HfCIjA9Y1ZsIMfk8KMP2jLs3A3
NDDxsSvDuU2yzYnAMjFgMk/GLwvTNQSPBMhP9ihT+DuyZOQ2nyF2Vhjc735xs+7p
lAT0k9p4posWSbiccfYO4UnOeCn0y19lnfM9ndfwX82ug4gGx+Bwkq0GucdhgRaH
Uygp6/xjfkgHOmJR7mpfiUAbiFPvzKsCsIi5k5CLm8NDWhBUWYdgjGhTt4PfUZSI
xQktREO3I84mYZ/AfNmlo6IDtMdIZFdzNEpL01CwjCjAhIO9t/LxTntrjaqeZ5nR
NoL8kCwWrH/BPbhLkGWgquhW/8O++jeUIVeXblXV/IvlBwNAW1gzdftWspyIOb/V
MHh4xvR7daca89GDWpOTPouwBdEhwVhaakJ+8EMkV5Wfy0LpVZsFqvH9pUt488yc
ulxfh+HFg6Phsw59Mw6TLbuW4/xrBQOGvzYie7/yjuzaQz6qDiqp+gtwQ1enaXt2
uzLsyTZXYC5k1rzn06cLr+8zRLvUaIwV7jxinBQBWOyixcrlCtnd51Vkgav1BdNJ
0IBOsYrHZP4CY0GH0G1KFDnuEWR8/YPaAEJOfRH3MizcnDvR0k4CF/OEKgzeokTR
KqXw05AsZoU0v1lfmT/fDgPJIjEj73sFHewQFRdL6tkpYZEqdF7x5FYoDL3cECjo
HlAuXrr1Ri3Rf473awuWGubuDbFwo4g8xnd/mHvMfu+kEvh2CAfrU/WD8+ftCAl9
PpZmuHBlJtudNEXIEkLyZrpOEHUoqqckQhL3MfVEeoGzLp7qi+Gyv5V3gH/QOuyb
+KpNSLTZ7TJYQWCIYHbP4o1aFvYmvmtm9inNEod5cUSn9B101xO0A6uelcfCawlP
zwOx78r8nvjwTg0qx1iFWkc1hnihws4BEJ6hSiTjAagOL1526rdNnfQTeX9GabXy
1UMs5MiXWs3FAs8bT2/nb0xKWXnjLpRgogc/KNn7J+jt9GESYWcKfr2Q9CtE9XUS
dBgGGb9TgOchkrO0f7aRlpmX7IOCCiIZu6s1YYvZ76mG/MAWWYgeLy409PFf2RDO
nQXdb9dzsTLoYVEJ5JVbvwGV9c7qF3EMDrED29i13m2zeA/KZR5Ae6ZliE0occyc
PQlMnbX+BWmA0MNiB07FiNxEc4PHJaN6kZ87j0l0aXKACM3BY4XOEZ3HoU1bqydQ
rBcyhBLpvlsRvSYlGcx+nBrHMwEq9DrlBkyNgYbm4NOQKfRsyMfo2zmljqgl9jba
Vh39hoZE2ampso2/aUSjn1jGK3Y5zkxBhR3BW+DeAcRoRG3WU8rUraIUA1NkFN+N
/iG/uhzdMYpeKd43E8EEOWjRpM7QA31E8LF6wNl+8WcP0P+JvoxgjNgTpsioSr/1
aAv06/YDaeUTzJ5rEtgDQ35O/CBJWl/n4cSoWZ7dhza7ajUO/ZgXLvu73VjLBA+S
YleFoJnlzAXYyWXJwDx0sPscBQtBrvEMumGAMJszvK2HAYwCkWbTceW8nHGveKGZ
hmagdIQG9bbNtE5x5eF1wunDEf+j3hxmco9b/BgLaEAYPnJVdvM/1V1uRn0uvXJ6
gBCU7zvEyC6NUub8cDnzPNaR5xkRvynvRiXAAP06YFniaDBkwgoQYhcf6fY1Yqyl
lLQ94bbROrsPrKEwsqgHRYYaoZ05F6jGrJyGmt4HkOxMDEoakpe5OW9z6RhbHgl0
BTklA57QVyiqd5tPO4KIhu5Xdu9iXErZGMvoSTZlHipebK3rRGZhDy0/LoPWxInT
mQu6k0gefC9tG+o9t1IY0GnplP8ShcRsGZIuh3DQ/u9AhcrfrWopy1K6/S1FXYZX
cGcIJjJ7td4JvxTP1OP+zLmNIDgxH/6p5mcjQFnG3XJgNb5TJk6Jtn0Un0P3NBKN
dbvKtuBpMXob6z7AiGRK2B+o16rKghNcejOj0e6EFq981ZoKNl4LSKxe/3cxyfon
Agmqe3mOvqmm2D1Fao+78ohwLm1twvxnCyl0/qF1xN4EJPPWaBT0btbJGYEHAbwP
Gg3gYx1oEk4b+HkGpDGIZujwGMX8fI8CLTbZouPLf4DNuh/yasy6XIpP4+GluVgQ
RAdNPcosQWc66CZyKRnWA1qdqIHFELgW/yoPTYpxqyyA/HKwnOmWSrbjvy/6s69K
WusNK1de6EERvzqXaiRKO7wBgAUbsh2ksY108wf2ooldwxu2Ngr695mseALmkgSy
pq7ek30kGvSIkF9vExW7s35MnWZqJs+JE84FS58rrrJ2PQLHneEWu20qYpVHdxCb
/3MtvpYmB30zodzi5V0di2HFE8ckMOZV8YK8gIVxFtMi+pb+CFL7X1JuKEP9U2zF
8HRP+v1rPygrCC5wMziCvxuzYox+/tr8+ODFH3zytUuRThupe+qqbRCiJqxyDjSU
r/Ont27yY+0Vm75INTfWaD0HuXd/xd2VudIPheBHa1TBATyJdYZS49KbDCkPSSRr
rj8paaXAxhABj0CYp/2ovtidGM+8XXMCOswciNxYus9Vv7XH8KOLQIwOzB0uxnMZ
wZkV82LnXm6dXLhe/6MtvNv81IUCOuQNKqsqRxq/KBdEGJorq8jp7RgfiOSqwiJT
NLIrB5VsqrVQKPHiblZONAa9YRIFTgDxlDS/qUHMtERAfs3r30GR/6UXGkGVSoYB
enKQIgMkIjDmoWf0rA4DUxHAd3KZUjPqkgrfEGUEoClKwt4Pgj7xnXSDQCLY21tg
9lQLtNrcVh5xf4YggRwQc9dSw01gcy3UlIn0L8Mi1KiypMfhThHjvpJE8Gbc/Ws7
47LwzSdDPm9KMoxd6R64YH1/HxmnmZ1Z+Z1EtOF14QsnfQDP5CgPSIEFG9QtbZsI
OM/vAFAnG6ajPKB/pZZ9kBiG1tT14238fgnfetP/B8Mqfdcctx7q33cdRIvoedLM
W8+Dxo5eX1I7/40s8q7cVO98uCSpDoCRY9b/jNv7C5uO4ZSrQavzS/Vv45kACAF5
O77BL2AnUSoqp+cbY/ZSWbiBAPgwko4Smobzph1w9fG7z2UZDAkdJZK1laVvUExX
uA32utza/+YdiYWfp7OsBK/CNRz4m17nkBSIMAxC0Vuy7c6+OnSWKdd5n5ClHri7
HRi2TKKOWbVhPXc/k/F1OA/nbzKm6ZzgJBTC1CsY6H2Krz7zyR0cMkICH0vSwx5m
VI5gFdvDSx16t93MBq2cdD9ua/BdGxWne1Mua5z1XfuBA9K6/wZtPGL1ErsmXFZr
TXsweuWjH4KR+hJdjGeykJLot+zMAPOypP1mRTafbfjIYePprskW+gYhYUXdbHLf
zFqIkR0quf6bwT7cD4BcqutAEGV5T7iAADa7Eorxzz+uEV3/0dzeEE1TSUf1uKoL
+HXqFBpyz1fcN0PFGpxkzCsV5f5/bC0w/HVaq0+ouMd7iKnkQOstl2yNGrHxql5o
boD2MCzAgsDXr3TlM9x8Q+2kpUk1f0g7HbmPiisxEedfEE5Q+OoNxUZF11287CS1
FEeGnZRSPKUcMA1pduVwkktirrAlJ2Hig4e+6ZgPxWHFgVCFrjjCGbnJzwXHgn4I
jzoiLI4bvBV2WMC6+kf/ohkkhK3AYoljd6VMbtisxg9aCNmBzMBeql8wEAfugf+G
TJzwQqRFdJ4OHMdTjyDDJkhBImdRuqeKFFjDkB/9Rn9xFWtJVgTzetDAafZ5MZ40
bfGVqkOS9my1bNcaScD71nRAxcvvtUV94qX/xMDsU7TXZPYDzsJU2CmD1HYbCU3E
wrg464kT0KEXkWj7x+5X87h0ZvViJeow0l1zg6C+buHfWe+IckmCjqe5MyaTEh6H
LduiX05VGEwXKjxEBfjURi3Lxx3OTzMhJMGhlc1r59Udo1iK47Lpfqo6elrPfmJs
+f/E7IBjm8HTBNRGRK/v5HCaAsee/lvZt8CYgIcTqZ76rsIdIvfCPyPN1GGv3169
tUk0sOkb4OOVTJigYLqs8mwxiNCWdG/Hzqvw1XmhRmkqtO3dMi3pQyLnuA2Iqmfd
oW1XUHScLO8kjoP6CRr76qxoZVGU4dAYj7Vu5MG50oUvQaWWT2b8H5tkE3/YzPoN
QBpNb8r7NzhezCBy0SFmSqPoNF5r1NvJonrKHDYXCMtbdIJYkZQ3Go6gXzBic0f8
C9ZXDAImh2u0YJaq97QTGQ0W7O9fbfIG7WVm2XEMMvAc10XgQyxi9eqaInJ56FOP
+0xlxFYI3AKzBVW5H1Ri87Fgy59guGVY/+eBNqSUlfSuDKDbIAmfis12KQXnY+/k
7S78LQoWgqR1T6tfdCs/xjD38W0ihqzycTFqK5wFlSla8Uc6+brIZnMyxvMNVplO
ojyBQVnDJ9vtulSjIKDeVM2Qa+geOuq5pnz6OOQRho5/Iu0WCUvWUF2+GG0sAEpp
AGiim9jkQBzynH50h+X1bQWvEsOYnuCuCrtYBmrnTuf4XcA7CdQRjz8NeZXqFPmO
vji1lTnvfiPRISVUMXsvDPMkbs4mJQl/FNL8PY/gWQstDAP50V9z4teBtVLx012I
TecotZfLFhzh0t+vdf+qNpu754lkRbnKWgW1fC6o1WRtsLHfzP2VIdvLyExtD1uL
QisF5KahQVTA5URe1BMUv+mT90lofk9khvF3CO7kyy2BS6kwex8l9iP1V4B88L4M
5D8f2k13wMaTSp9HOH6SajRCgQuLYJvGDV8rBoPn5c+20/rE0DyuLvyBXMYmcOJQ
wNTg+6rMpBogFaK1tO5/8xLCpkF3pZb/Z+rHYPHQlypOAHlXNZd6sWplCA8Z4kTm
wIt/XfbrrYm7ItPkK2IoWWi0VL0xZzrwuyaaYWxdVvf3YjXyu2Aujvmq9wW4gfRS
2R5VyGOb2FiXQY6E/C6691mJ6pgbQikXXx13HkhvHHLoW4MMpUq9GZNq6Dp4A8Wd
gYRpmNhXdnmdtgqvT7XXqujLlb0zimOnTmx3gGqKOhtApzw0eyxCqbHy57NRfgA5
QtmdAiqUK2gxtK15rIiWB/F3D/WGFIeCZH+HrfSka4JW8w34VAsEK0T4GovhYEQi
JBzxVMduw16iUefvwDg2T9Ns6tptxzBOos7y0jcSv6y6vTbINVBdCGIT9gJWduSe
og72pLTzQ/uJpEyvha9Dke7FrwnMsZmyyxBNG4UcNnGSvECOO1eZDv5fPh+2nWLk
TY/V6wriLIL7eYPSNKtQadzeqTe433rfYenKmiIq5nNJ0Zzwf+hx/UOaLX/ILwGd
gr3Tczo2m0JZzyNtPhoHy/Tto8H0iS1mUWSwMbV1gba7BK74YCCeff4jD6e7IfBE
AULT+vxoric39Fwoaz1oqnIlIJ8VDs3oKLqrPAYUXjLA/gNrqW+SptZA+UEsbUtR
t95BFoMgFuI4Fjd85mZNkzSz5i6vFBcEBye6U+Zp8nd8HpuvXDsMQTKJC8OBb0vD
BUEnlsXMg0+WblNiFqoxULPntH1gYrUKO4jvfVXI/3w75vdPtx5xOgWYyFTVyVjq
XnDSdbGLLj5L8f3GRShpNDbjYL7mrUaKU0qj+E5HDcJ0cHDZgUOY2hqC8jLhVvzb
W3RqSI0nfMv4XCAJ+O/v6RT1fRy4duWhV4fq13LUQZjWfNniVd8D/jkMNHOV0RC5
zM3t5frK+jZdNp7sP6ToyKDHILAVp9p3qpla5wMLLDxRdL+0LnYqOyEBhTKyH4+0
cNdiO+ErAsnW2eLhoa5Dba2oCYNl1sGLKWmjg3rrR07+GaZiCYsbffu6oBOxOQaS
mlsHmaEdKIuPtQ4hfstzef5YPlkhdI3GtGma9rDPdfzuowretAg6Cn+ETXImdpjS
7gFa9j1b3ZHVpQ0R+7w1YcRlnADkrIXeOMtOo+59PHY8VHyZByBQSkURO5fbqUQ0
qJlEEN9FMmcSZ9Zf/voduFnT1Eom0ZRKXkHXfD3H2f+VSo8HBCr2PjeYok7CJyjk
2sHfvNBmR5xhBB/2tJPfm8jwSg8y7NswE65CW+h78GMptSqz2mD60KEVPCQYNXXf
IImZdUDrqP2/BrkMAlHF3DxHoD0aK8bAsgzzy3ZHf4l1fyujcbkYdsPgyK1H+eSb
sywZ3ncPmdnED7ogAnADmlT8131OdR1n++qQB9c3cfjyherHCOI0GjHO802A24td
7gZxAySsAjl+wsd5mWWkFMT4kTYKQw3Q6nN92slilUqeg5oHhh5dGiZy3UbDXZgn
8UOfelxBVGXjdjKLSXqtPXVcJzXztu/EuEWV20Q166w5oJtgVvTzcQZ4YnqKq1R/
sEUzL+wOTtlin2qqG14wA/OWuRPKUMGNW5SgdjbgF+cLVdshPNn+q+lnqKICGXGQ
ofxplslGJONGEXpSrJ4Za/rfo6m4JwE1VpsT5p4WwKAtghHvXaKiZBgqD8JDjrUM
8PMSGhPD6N2V25WU+NFBZl/wp1TXThA351UrgGkPtZkvRXaOggGvAfAz0E4IfvP0
Xn9KSGm84hVu7C+3zsVMv62ZRfw231E49njV6gVp3zZ7k9LtMfRu2F5vbp0DxzEx
UYEHCBoeWu7vX4II9Zaqc4dpYrzXJ2qtRhQDKIUXeBOy/TveUvF922GbjpXEk3G2
rCYZumpjbV3zBTtWSFDci5acERBqnfUOOaLCmIjOmbc/YAkS6kbSz8+DfqmacemW
5La/1TU5jcrsJWD/1OqAYd/VED30uWe7HPRzff/0s7Shj26O0BANhXerB5GML+hU
Y+tQL1EKAHgvSmgrPEMIFOcrx+WnXsMkKMNfjBPc0J/pOT+FeRBWiOeGMJrHnb8D
lF1SVTcsbrwhQvRutKGcfs+0Z7//0xqHocV/IgH23Q/sDDrXFl5labNPMMkDpXF8
iMO+zvhT+BKpb/HDMNhoukt5wJvstO2Greki74o9ymyiaS3i6UwX6ZZSz+PGblrh
IIAaaz2ht1xrkmT1M8GtO1oTfgS/dN9e+6oPWnZZznX4+gtU8j38J4fWuYD3+7Ap
hMABLVioaYngJaSmMIC5JLB+OUI2y49jJXpJhUqRK+PEdd8Ev7kfaX8BYwOh6awy
tGZlFyD1vGugjXBJayIgU2foCl/XMQMvtuxPgHwlwSzq9AtaEvmaqdsd1fAnIlwx
DXJWtrpFXQPboHo2ouXfIpz+myhrhlWRuTM7oY7Iu0nkzTZg06J6RZa4xQI8e/0e
ZiIkUxFPGj/4XU8WoTn9I3qsBOjiLMWyBxS3W3WNmpNvHhak/DlbxV8intBivaqi
SGoM0Ab6fIMxedAcN4h4HKe1Xg/jigcydxTKP9GreQlvCD8B2rQcQ7kGUbpzOVIk
MsiDrbFK05zdhFyPWGBRpp2VW3L4/BPkOiodPBESOPmI3a3qYV2oDb9qIc9DUF+C
KlxqN1JLs3jjJefUpBfq+FmchAiO0KAdDiA10f8NAo9aR7fLKrHI0hc6CtSeeVB+
yFe2W0JO1Plazet1qjbXmP8UqrnnVGLJg5eKS/Aa3BD5/Z8WZVR42Iuhf3tLS0Eh
NHizwpoD22kBZBRf7Ayg8MjgZJCYxxnNVPOqNnnYFsZ5dOlpn/zZoToBAd57H73o
2UF4YE8UoJWFa1EsFmseAQUtuLmcZWQQSi9q5dT0T8Desiv4ZGYK68H8dlH0lBUo
Kw8yNdnc2FpnBzQhb60/3Eq9AM/TsZPoUkKHkwq5DzFJIgmilDz6NJyJukrw/IpL
W3XMey+6pwVvMRLOeSXKbKVYqU2HdqK09YBCiRLy3dNDbBxfOarVoFM/7+NO2pTw
hEifQYBvX9SVS9q0EWYuHzrn1Dsk1C2Gu5wUDDmcjXiUU7tvbcZ8LoN0o4/4mH0o
jdAaq7zdmWnhw0YA35X5eSsrQiZOqF28lSlvWo7iCD/tR+J4XwTNnmunYWRKcMP0
0hsQcwZ6bIUB/u4KvnkBDdOdDjoVoJjhgmWvbS4LehPsC+238MjAVCxwLE4u+5o4
Q6At1hrcQNttUnLAjUKUUNMsXm73OgtIixN51qLgtrTjY8o7fM1uLfpTgSUPUwfe
nP38TEoQxLi30hBrosNA5PaPiXwzXCp63gx09ou8LrJPCPsIxh6vqh7na6A0CclE
1KnM/LvjvggtbtSqPhxqlqjRavcykweJ0QO0fI6xxqMfcqCOQ0Hvn0e1z6thS5Rv
sZQipoEdlWy5KewHXTv+LZuFKxrARdFf3dTafezhfZuO85FqxOIsVL2co00aBfF+
dn63Qq0cnA+qD6700jNh1wzw4VytfTPmn2aVaAH1aoj/5NbdBiwJNoi6HASnC7Cr
X4AJv4zx4CSWw4Skw9JfbCzuKd1WKuIJ74y6uItbaenAHU6vXo2/BKaU1fuCo6xs
VYi5nNUucEmdeq8+Gy96rimEVNY+8v7OBgT2PFt/nL8aNSsM6NX9d5yin4UTx0g+
Lg3eq0T1Msp/BDQHwlaTdGmezcJ488Vgxwdu1KfkNeldqRI9WcXvtsRUtPOy4PQu
NjK5HA5unk1tkoJdLMQWuqSkTgX/KSvVH5JbXXhqRiwauyMJnjHjBcsHfErTRQ4R
8QRGPTW9rSRXhbVWTFOilEawQCligPxfIGMGRtELBAaQLhg6U2JzBVfEIgoxFsVu
bFeccQZPnR86VpqC62xWQpIhI5RkgZBpaGconkYL+gz5AJ5UhlhCoJ0FT/bfRO3e
DtmT2TUolaNPf6Rct3tiFoo3/67bUdoX2IT7ZrZcJG3yr3eztEdIrafzTDh8BDGz
QE27s4K7FwZo8UyXx3UukJ8oyAPH2cSQJrv9yMCWWtxmZB+tnZJNj6o8rz5zxScI
hIvO4q+7mMLj38pBB5jSzNeTyrUw+3IjMi2mvRB4jJ7Co+cSKjN7FLXLsbs62F/m
X2RCxDf8vDyrZv05NcGI9Sgw78gJxkkHB7bWkDunShBlWRDP6m9Thn9e//A+3GG5
J2jPXo6VqXHtmvsSbJBntgnsLLZsInzZlM/Ka2OYreM3n6XwBNpM0yid8TNnRoKj
dBJfe+pRjEiOV0K5aqSFZpTW11fdPikI/+8Lgmc96/eILj6vf9UBB4qk7gddGMzl
8ZxiMYutHfut6hwW7jOk+LR2pbcPk2/pc1G0KfbimDvD1nPmlaorWQeDJXOelYzw
EfmUlGQK77c2xPHpIQuENkcF8AokpxTALU9huqDwU1tnUXXz510AaNCEePDTCyMx
XbriLA3/47qQY2qEA7upJGi054+jg5doFXKvWGJYr6sZKOwr6qVQBkhhIrkuv8Cm
Kbv0gDIlJCGpta6+/HEOwMF1Vf62rbeFVOeR0y9Vb0cPRD8qsnpNOyalwAIFr19A
NibwmaJOCdwOJ14oKsxkE0TGdB5Vr9YKGDVK5A+mzOGa2QjyBIjHEvo8h16oZRW0
ngA2i0LT27X723HmyooO6DUsqVY8MKCZMzegxlbojpeSaM4udHGKD49hCLuD2M0c
h2bBWVZPqt0Qonqo1NIxeJCNXEFOBQGKdUms1Gyz2K1dnggBIfNC9bhm9jRfk4bZ
gQVqCvhzLRPfVy3TW0LK7d0RbfmmXwlaX5tBdqtx7WZy1vACJ1r0EJyDz7C7pC0F
69xO8VuS/VY1D9NyfAIujpSHqfLMP/nKwISXPo5NzA1eORpfaXwKU9XzOpgngU7A
SvCZiCf4T/LmeMJHXp+kHb7ifNIXvai7Toyz5Th7tPT8RkF15fdYqAa4tdpW7zit
XDLnEMwCVcxe5qj6xnn4Rd15g2+bYcehAlt9B/9kNfYBRuDFDen3eyMHAkT3rKbv
XTL6VkGk9jR+Z5ThQusWWR5CD2/zZ1Fyk4rZKE5ZyqeVCtAFzgCd+EDd+mBHTGFj
ik1C4cJU6J+kZCCdAH2uJAD3joZhmW7kr0ZsNsV3jHNtCfkCAMGvCZNS//rdb9FG
Sk40QT3jN6GzyZYJnSULN474JZKoLWJjJcD9cJI75RGjYmfokH6l+HX0My0ZcJPx
SA9vtDiMaQUtsoYqIktTsJWgpGkLmnmcbkrXOXk3Nw78Cx2kGbzSlZ/CiT1nK+sA
lPaRlJ+Xzkz91x+rRlxvsDh9ifE/rC2gwaKoGYTIL2pZTsZ23emHVUNr+NJ6mxKb
lu99AD6kpLMtg5+W20zQOk66wHQRfXfM/c6oUqSaE7sAb83pCT8eTaUeCxm2Onid
zsT+YMR4VI9m3yPeltee78Q5bArE6+Q8VdoqcoKyItJ6mvuAgnMxBjtaFk1Hr5jJ
Y56JMMWipbNsxKajtffQz/MdzHgAkLV816d8yRWvJJKF7aAL28iZp2Zwmgdk16ll
7MLqOTvwv4PUQP0kRlQaFsBMJzJLgII4quGgfhFW5cTPGLsvvcCP4aRu1dPnDC/H
N1FooDhD+xNHqTly5sDz0EeurbyOYhu1qmOEKn+X64GyxiLQ8KpJGPMo0YnXhQk3
R10CsLq5ErtfsjvuuHWxeGWMnqLvwYyGjN6crB2+7IsQB7HF5nrSNlbkV+z1xngP
e/OeMI81USyDpvlv5oZslmWEyAJSsKQOhpDEdBmgs25U4BFIhUeVtQr5jwx3kzpi
qmt3WiTtkxhG7mtbAVMe5IxYzngzz1VAROrndMSWcbqelbdXP96L/VesDQLD3R5+
+fpSIlmKxotRd+sUj9aDjXpII0+wz0wgNYiJqLz06HZj0VMxHo70wyuMxJH/XaDo
akR72Hsx520b2ngwCBzAmF2pCEi4t7pQdv/Djk2funPwC7rdiCPAP+Ky0AxqEviM
gyAvGvLXbEZ8WdM5wjhv52KWi3iZEF7QuqSoha2PL0yCXp/qjpirbsl7h8JUiONQ
XQ7nWlgP3SUQoKKO3RWD/lvYFX4JtE8+DgkabxQLpQh80Eh8SlAETI2241sVBzZJ
ei/Nd2bFyNdJLY+4O2qKTRrq2mJcYFHiKzCtJNIDc6ZvHsRDR7G66LeQ2jNDA0+g
1ydh39GM/wdEr2O4rKexYDP4C0SjzhlxDOuxptbVl/M93WCrtyo3lUys05VPX1U0
rJoBh7iVyRT9jLIilt8xvILwmL+++kYD2/TxkPRhzdmihafb0dM800GzZmS3SqvH
rS/dLUD93ZPJIk/LWyToHZSWrLdmvD4w8wS4JbedNtUznlYJQDYiaLQqYidGy0ay
dQPDUCyz795hXTQxjd7xZ6emr504Vvfo3Q27XRRrsCsGMfjjiRaxDvdO/JHTc1wM
dEv8LOzpo9IN0o9PAV/Aq3mOSwPXuzdurST4e6Oqx9dOpG5OJpEKa26ZZjKADRhQ
gx4CUW0Mtni/arqeW45r11NbwNWas8HZ4g6quVQ+Z4p/8OaljtzbsbUMvHSCsjZA
6ecxGdC84EXGvsHm6rH8YfwVetOktvyobNwRlAT0wCxXIDt/1zJm/Z8gPmz/tMxw
TVh0s/nlJLLT+5k6OsI7L0sfkl95HYpVJKpBKBWVll1Q6c2MRMJt6FrMEre2ZUZZ
WiE16N2LJbP/0at4u+t0zWhGWo0neP4Zc3qIA+HyYbFcxpPe7b3iR3DQBFz8XfLg
5D5bBk4RvuxX/eXTvH6vhn6Ickw/gfLOU1DnmFRS8UvsFx9tVhCSdRXm2gEky2Ch
81YWim/1//NezWpK/iq74kP9x10UpmqAjM7gcpJ2ptN2uC2QGCw3WXLDfS9mQBvL
YVeJQu/kgCCQTKk7vXkparvcwPAMAwoF/KDDJL0VSlS2WMqbFzrmy1eFH2YxDFps
NePtkF6p2+fQl8E3ZuzMMeNkpZHuHGg9QWlB+qg4bCFB3BAYy1Ej0N834KHnsXN8
3+fkLUmzYrMAuAQgBCDp4ewMm6DqQxxEK/Mm/3RC1uiU/TLVIT610Y7vdJO8MFoj
gWE8hywgRFPTTsLMo8CC/yLdFh+4f6pzevLiBQNEWv0vrcGSBmqcb8xm2pRnS73/
5XipMQ9q2gUiN6lXx9K/889g864DwMbhPTNJdn9f66jk73kaUsEeejPOJAJ8/bs2
xQpyO9WsvI0XbcyDAztl+Et/qC5kdc1PiDwQqIFE18VI7C8yJnPZlwYpbeBGYvWA
mpB3Vc75NTd0K1fu3mW5VjniF3qkQMq4uGB3MxYyJcXxMYyDk7+cBjQNLWhzjzMQ
3I06GKO2xCv/KylUvnbGqnCbG1mpGLARpIr+PuJmVvuOBLPg/fSV62xNphpeG+z/
aoatjlfkTmzgYhyNPT3kMvdjCRnoEARHCSa4AQ70EZG9YXqQdD/6yrslLvkQ3s5u
8CuhWpusCdqsMG9hNsz2aBGoqQVUho1/Dk40NQHOu7p79nsXTe61VODB9YezXKaj
r4StT37yN1LFJYzp0gV7L+cYkH3+z4fjAvpYHsQrIsYKC14AQHFRwstdzHSnuzew
LRIwCFGb1PcrlrdvdkeGoRKMxc4mDZP40Ce8S5gOu7Jra0cg5zWzTPqQNmhkisPL
A3uXqroQYkCry/5bdOUzfDnutdu4J+Povp+4SLT9cS63k6kNv9VQAQaK8TpzcwPd
s+C3xtT7MCD274Y4nRjhfrq67sBfOQKnKuqXQugSE1FQNIV9Q5gPNo0Ft+HnI8KI
R9GKE5+/+I5+NUZTy8FvkEcvD/v+EIVzfjcu2D83vjPX5IRQCHspibiMdJGxrG//
7jV3eT3WfqxHOlQwJs7GG2cLFaJyXtr2OlhxVXwDNW9VBBStBHZXIZHdSDcmFOUW
HGrCKduLUJbKjKWhz7WcJUNtx2puusTnb8vTdpr4xW3/ZS9e7uJVWM0pjyH4f3Yd
bGqlGnH6G7+yvsKDghPjHlXNJ9aqfJoKV0zhYB9qk1BjouFvr1I4X0Ja2iuWoXDE
boQR+io3SwMgrAErSLJThS3cBQ20PMuk8Af1gYhgjv7/x4wq+h1w9yakokm5heAn
b6F2Ih/E7w0oECdzNauKCzqWMFOaGGyinsAWvIRhjaWQHb7P5K8v6RlB75fEfyGq
/ayWfICAPaqF6o6THyG7bQxxH+MS5zMlbzHZwq03Zp+VU3HwxR4cNXnfk+Nk8pUu
JzpJ3xdrlzadnoQCp8z+nLvtpRFk/2OgtRNPG1sftUJ2H6cm+qXTtEUBI3DxI6ZT
lzfznme1ksrbvlJd4Ws3f077IYvB1ks3mHXLhkW/MA6/7pnPH9LTCAKSD2Vn+dWG
iJf5Kr/YgjoOVY+tOg8JZJr76LbAQ4CEWPvI0HTy5cLNI69O27i1fUqw+hHlm7T5
OLja9r6WZxgp1UVnKbfQufq96PYkp80QHhalYTA/KV4e7OWQmxtO3aG5Md56c11I
VemFN8uhXus2SD7ZTseSPpQfldhOsVjMl6U1rRv6lGVAEhv3WBWQZggnYYvaz8j3
I2CVHPdCk94LU910ztnYtFkTiRF5G0sqOM34U593kOL3ywdXZJjN+0xnXxSd2aA8
oNt1SeXGEf4sf5t01JDRVaPIED9zXzQI+9Aoid2dlj3O4wl83MwspYPj19oI2g9j
k3qfFm7l3k/E7bWoGMtH6d4gx2H1rtx4MtksLXvP7nQGycsnt2Tt4aGeXLWPDDf0
iViIDg4GQ0I4cJzfAosfmYQJWRIjqNjIruHWz1Ec6WvUrwDd09Z1cFlFw7pdcAg3
XDAGQn7/rMZDTRKEM8axh1sbl2Zod0ebLxYD+swQgXz25GDti/Yor5M0UhDkbffb
3NlgWznh7w6baG+oqT2orC2YfoxRXmMGsnl4sTUtWVJZ3Fw8lOs5Lvz/JyHmk7mJ
t8g0lwBn6013hnu4g7or2EW5ETqihC6Fo+Nhd7ZHA0YUYiAsPxecSm6Tnb6Ar0dg
DLhhHIJouM0iKxEJNP6621+C5weQ2I67vF6kwO+MY2TIqK3IalksCW+IXDL48+uw
OTU1Dtt47H4FKBfEsYX/Wi+Qijx7LtWmXbQ1su5qBW4kfoWYpWOOYDS1nNrZ6Us0
18bX8UpR7TohHPkdYF8/XPBViNB2fCjfHuOEqxwb5ukg/RN9pJOME+tfS8UC+Pkz
wLkP+raCfXDZk3QXQp1/Fzt8GloKFw1iTjYg3G76VP+xnHYs/N+t2bwPLS98taI3
R5IIKE7DQg2Ot2T0uitElzEZeVgizHsTX9SmChpAkqAnebo1JKC+CnI2pl0h8aE8
ocu8v6xFRR2tx8rIrzfAyoKsZO3Eo90D1nGr2wqtiD7rUypZmJTj/bcMUVKTWOn/
pwPQrLX/rJrxNqCr+JoKS0wofXh+avF31Apa+nZSuPenmTUpwQsy24Rz3nY4QEtV
nyxhPk9grb7TsAIN8e+h6u5mQc5QDMczzOT5D3CjWlH6dYYD5txb9cJvPYYyFVBa
eZDQW28Bpy4nOVqED7pF55yBSGvKCYYMsskxQUdDK6p6m8VHV1+uii6a1u/fVsHy
Ffd2yTKEF8cq1NEFetzRbtjAacm12o5MYb5G/8VfIyLWEbpNdOvYGNLn6Nl/srSn
q+NhNH3OurFYBCyw0m7q63iP2Bn4uJSmtkS2MqIvQk7DnN8QW2xE4TyNHw19Hs33
TC+dtcKERK6iF9qcZeJtZlwnxUGSgcjZQBZLNZyzhDF0LlF4JNy8YtaYk11hm55I
r/w/i9mGj5hcdlZRFfGeUt3RejzcbVxtU/HCLZB8z1qPt1ia2JGOl1/JKZ3i9DQs
31qs6Q0gPPz7np4B8nQNY6XLZ5cM1fmRoF280QKZKahV/7t54y/Uw1TQKZdIccXD
ZR4E66c6ziU2nJyIMDWOZRAyYSGviZidJz7TqnOpSKOYUMtKLaq5ED0kaqH4zsdB
lzz64HPlA/VR+0I0rQ9FDof0B6vVd3TyJLS1a+qBEfsTPfb1q0PbkI90oinkNfQ4
DWMmtFOpDusH8M5bBVw08guA2ZBxLuw53WXuA0Y+wqtXeXfEzDoeNxho/TkUuNKS
Cq/Qf+ksvN5kbro6QWnq6kMEyFt/cWA1M/f2M6/8MiRTNKDvb0jAA6aKcbvOihwG
9IsKKSIwe1dqhmrmS+U3UTzj4tcUU3G5VcHb8GFxl3LKFge7nkwSPmrtVICQEHTy
/ifxHsjRB539yM87AkWLWJUr+s7QllJgQKe7WpXUlyndQbhD4+FX9yxoqP7vGWs/
RA/sX9JxW4rlLPKDz+4vCv8QrtCArfoPepli+NKbJTyPMLLjuy4XHhSDqXG5Imrs
F9+o26mQs5GQQAXj6xTDbii0yIP7pX9hOUqfUm4iXJ0UyIHvpuDOawoRyYpKlyyb
imeGtR7s9N1cCmiPcSDfpm7TR1vRtKQH22HRRVwnukGJZB487zJ+DPopcfJV7tns
54EvAM+Y9VjftqgsxxZ/OuZXVZdqp3yXwNqYzMNMY7HjGALJ1d85ObGKAvuTsfnz
ZpY19M2s9upj5loGCXXUmwwFORyixlYt0cMVWp4k7sJxbyfPp1AkRCFnBk2wDpYQ
L9Lr1K2MIYc825xsOVfuVEgyXFDpKNNrnbXPSTRY1nmL1rKYxMH8kfACq93UYG8u
iyrKJZmBe73l8UjMKeO1tETw8VpDGmBhYF3lKtxGW3UbsLsv5qlEONKq0WSoslqc
GOFX5bU03ot/SFObWCEsdOdZMeIbAVVdJogqqPaT4n/IO90alXmUaxo6QN7PzbSY
MTIM7ItWGHFX9jo2HcuPK0ZCfm4cbMh6CiHFXQDg0f+bsd6WKRwnmIIhKCyYpZ/1
z+bPAzXQ2PYgXglyoCcSpWe7TGI47PK1F4VpfdBYG6whiFkV2esEJL61CWW42pv5
IapdNR7endOhRjsLwSj44xfeOm9W6RHXW0+zo+ffbX4ctZ81SMrjuJLSMHs1j3OT
5c6r8kt9jo077YsdqauwaxjqvUh3uLoKPHDtV3GHqls8tKDwI6R7+N9I8rn+D1jn
zLU3Wp+kFAPAFXrPhZ8pw/tK+E25B2LLaJRCd4JX94zyfMZ4KaWlaA7c4h9/tYus
yLfhUPHS3MArRqZ9b9g/jIneEJDHSJilWD/KEMS/4lwHz7oPArL98NiR9GsRjAfj
sfprHHeF9AGLaze1KhJvV14lZUsMqikgmezpcME/pgplP/rOjiVncW2jsYegMBiv
DqsWg38F72l70QHB/EmO+7p6fge1Wini4bRIpxTfFVOW0vljRYr/qBtipedzM1lh
r/Kmh6Pzpm3abkEXuXFZT892zVjY3Pl+TnKnA72sPZXUaLKVjazpy4mPGcupTvLR
HQYT8TW3iCNdWWxGEcVUSijmkvkxmJqw9jJueXYBljMqigZ1uu3JSxllzqAkfmYw
ZTsaRaRU/YEAX7KQ7NRUnVekXcggtnsUHqSm7SvzeQDXsEAmtfFI+fG0Y50oQcEa
pJ4U3txOlU+eioxDzxYoaMdtnkEG8RJIubGaWW1wzCXjCWwhQGW0Mzl3Y+mUNhMu
XmIt/96a+P96Y4bbWvMIDD4gzZJ7xf8lZ6YcCkBrwWCfM36O3sEe8Vb2R2hLg0y9
ypT168wPjeDrPduwJ1pF5VOrX01W0brDUF2qIzudg/8Ph+/smFBvuDEPl1PHEVgU
hyQij3AByjLr0etlabUUkys0o3x9NMvZxJw4pj+Iel2yQc6wV+seMXr9Mo0LLU3Y
62qa0Oj4A2Pb+g6wiXcxDqdOg2TyNGlyaeZBapm82H8aWlcxZ9idvUoV9JQngo52
BKQfY8Nt/F7WaO5IP9zSpnhwA0SC1WtIzJYrLxI/YZpngWz7XejaBZQ7cgrocTGu
yyjBz6hLDFSK5U+vv+PO73UTE99ljXEcEbl1pGDMvrC/Yms/EuXp8m8DiTHkjA8F
/n2z0QPbgA+021cyfvQMNzU1FSTJQH5EGONcmQplo595ZoqZ6Sbzk81Gd+lzMT00
ibHzgb8R7FJg+alfWZH4yFubsz1QPtEMNexYPWJhGkrrT537dSOfLeO3SUyBd/iX
IqrA8S4Am3b5tA2k3o9X26GsWLatqLCAd5L7z8rWYhy4Y+CQuz8dxTWiwG0SUYUy
yswYQwKlCLxwlRKMD/CHFbWciHKGXnGNNZzK0Ys2uybCDEPAjz+dAcNhhD/mu5Pb
zeEfcQcuLbh1jx5cttsBq1XuOLPBKoV3IYDB1YVJSd9FEOk7tz1MVHejbpbhyVyq
TXPqwdyUGjeui+YTNWZNosm+uz6f3huyMM0vrEnz0XU97+QifXOOSGd9p7YR1fbb
ioFY6EpbGTmdkf214vDp9T+3lU3ySHS5yLUupCr/TVRRrALhp2zXPsl6Iy93lwF9
LoG+ZkhgXUm7+GfvutsLHON2QAoSCHPYZsE9jtfHyKn02lpcSIECj57T0GlSCnHx
mBbVv5VUbbIgRpD2katCknTAvM0O5N+0PexIXHQW7f/nJixA1dkMhR9onpN8Jzpy
cYl2hfY/bOcFd/o2HkyTp5POXNC8KkaCbuAr3s4qeakoBDa+aW6lzrdaD3lwL585
KQucv1qbRQtbYZjYZkrribwhp11sHrGt50HNFcf0QOkKSN3QfCzegj216SZSs++z
6he24m700lpO1vUtikFGNfIAhXNzHAP+pDJjNGRPxgfH0OXlF8TrGSgPCk4sWUN0
MYo44DsGtybB/2G20D0qehB4gOOGWzZRGBiO56mvD1tGgc3/WdgCASX956yxjDws
RsFo2+3v0NaisKLtHGTCjR+qWJKyOLigfodtOhY0Es6C4RKDaBuAk9JN1noseaFu
91uJQAYIktiN3KlJHh2+VjOS64YESEJ7GBWuTq8LvrS/5onQhWaPIo4JiaAagQgM
uHolyME/6MzXhxENDdbJTSaYp3rgqeEYrz4rQ5/YngPM/FZ4aOeWbY0KsvT0j80H
7mEdMr7KuHNqd69Dy9EVCCiUaNKlzknjTNiM4I6Qkv1pOzFtbQBYh/IL1L3DgOTy
bD/IJ3q91A7fixefcuexHSt/KZovW0KekxKbcru2pEzK2HmRFC80KI3arYQDhyem
6OCRzvzs5EeujMvPr6e7ChIEqJ7t/fqQ2608KpKvi3jmy/kdmXM1s3gbP1zh3rB9
UBYgKqbOR2ffiMN2WvaZKFum85f7Od0cA58QJnEqZ7+9o22ZJSCpWjPMq+P3kR9l
IdROG4HtGMbOWOjqoH1fjHi2+t1jgrYEirZM+eYznblcmarz+7yBAiELAvtp7hrz
tcp3lQvR4d1KLTHGOlkqK2yxtKuwGutKkIYHCMi9m3joo9baKjsBJKZEGxcBstPv
LTEU+JtWNNf6MKDJyJWS3zwAtV3UmGIKjOg+/kXB8rZc8FY8wSaMcaLNYOU7H4Oj
MkZu/LnkToW7BocBjo4a8JqnuFzAN5jSzrpQrJ4Tj/BcWhO+NXtdihBuUnzNPNjq
ZIz3AOUQt4X6zgwbLDaYmxP5I1jtlrajo9cMWd04+O2TUmoPEnxBHZGNdc71uW17
bBoss7BsId7oZSeVHemIL6Y9pjJKomZd/Z+y1sXO5Ej51Rcui4JFT/1NOyJL6Pkd
WPQD7tsmbWMnZ33/c4rTELdJ3+2oSVJ/JmOknpQRRa0Qh3DfToF2KA4zMriGl1jG
V65lc0xnEqkRegHO4C/gfOM39l+uWEV6CY/+CuE7FShA2+P5H5P2hyGc01U0AZm/
Asf5TnvNiZZQYDf0aKCQ0J0m0skq15wV+hxLXWFX6qii7qS0Wi1EzVcd3pEztOUS
ylcz2i4myO5mBqH8UyDWtjh0qcULiAlyhe6ZeewETp34akDFdoD1s7JBOZQ/T1E7
qUALOv1ObxZ28zVHITLFWjIX+M7mj1vWuprgopqjd6dykeU6JCi2LkJC4Ijs05FR
nakYxh0Zcu6obE1mMpoLPebOyqfC/17WGQPNc45G5OU61lkQ1gkcGK8BSqlsMCKs
AKVUbDChnBqQPXOVJt1G2RKrTjV3EbiHhNpQWPPCCCDDXQoaHfg6h+qdP7Et6xn4
eU7R9SXwWmu7XZ3AKIdRGSzIWUjtFeGxnHSJhhgNwudnWkGxQ1gK2JbS8QXTgW28
kNETQHtmXpu/l4FWloj9WGORMt5ydJjarnViVzg5CV48HwRefDcw0eVnCLUhXrOT
fPGXR9iPP6wKfMwTs0c/KhRlxYEI4pqHvBZMxefi2sROfznV6he6dBNwr9vp7HS/
mVOzhfQZoAJ1IfGbjy7z9EC912E1p4pAMHMQuxw+7E9A38oh7m0RzL1RsGMIOz7l
qRjjogX4xQMUJKGbmEEu9Zf3JEfnWXUvtQYXo8I9DGrDCSpGKmcFJWG1ExfR84k3
NCKADxUWwcViIA9fOBaabecmAoQbQvSzhGEt0YtSBnNroUtfjp3gjLJiTsABYcBY
rELiu28WS+rmTbhaSiPe3z590VbSRyYrM5mFfOTDFvCYSzD6EK/crSTVjAZlbmvd
+6DWQbbkO8PsdTeft9Z5lyZWg6sFqmLW9dNMRzTK75p5NwLf3wKS/qFOhDbF1NWY
47gLZHq1VxxJD+yiDnoN5tsas3JapAkbjSSZblw3o0DYrJUZMRBidOo/cXA4GpeF
wUZPcJGtOs27KgE7pZoY7Xz3UiewdZtKsFHY1tZikUxWF+Cv1MjX8rMa8xrXjqM5
aq2s8YHbRc2FWrMiTSPV5kzI0NkMNJbHH9asIbWso8jQK+KBvXA4BMzovbppUIWL
o1Tiy/DyenIrcL2mzUeoqbz1D6vYlf0bAQ49cOR0L5GKokJZ0TWrHg+uiYXh2iRn
93TtslVjkTohMQ9Bir0G+/0BBHqQHrUEmttcNuWVBz/HnwOHIuLDKpaKR2Dr8tFy
m/oIQT+qgs+/GXky6gD1FiYTgU/tr8H7n2uQJqheL/92MxB/BsdtG/PB8dBnbUbu
3MKz8hsg4YZTV0Z2HDT7/YVFpe9ruYOLmdNLJEh74Xn5AAZsGKq/w4oiKV28KX10
kq4B2KbrUL1wRhkR/xbu6Dy9bNcu/dt/ThjtQpZw0Hk3qt34QnOyUU5QwtZuKJQB
ebvRK4hpesx/8SE7EQIz9fdA5zjlHcC4GGVQZ00VIfNMN2BC1SIefdcEBpAkvYcU
5pOagueSaJM3LhpUXV65/QaAfync6V+P9BYRSaOsbC6LjVat0l1hx+UN4W4h3k6q
vASh1qr35zBHmr8yD5J28cpkPOZjfLmgxaWUfKdqIURhWUizl06hp0ZlXwgvUj5C
lhDT4h2zDhe0ncUBB5bzzTmaPW3EUtB8dKE8+f2hFeo6QaKnWqNmPE5ldI85JSuR
aKlXioNrxzDuUdX34ylJI5RfWTV6jW96WCZWhDlxa/hM0x6zaYpTWEi4OMm7VizA
Br2QENw0xQeslnzY5eLaMtnEBg2IzNE0VrT7NqooT2mRhad9HAQBfCzXZ5wq/jb+
wzlYuEC3y+Pr6VFfOtMiAR1/iheqRocaklZR/V38QE8Zgi8i+8yr7Gry1nt5eLva
5OlWt3mdRNmC4GW/3JiVP2KBzIjyimW0nEcu+iEP9ZaJZ+X39MPz/9yZVBxwvDPG
IQwOYiOVZ747Z6B8jGS0EiC59RoUTL2xDPySS2fWvmaV42fSqjJrRSL9pfVEU6kI
/W3aSb3yBFhcZnKiiHVEm15M53EzLpsqRvqiqUJYw7gl1FodyPiLuyRej5DqU7yS
/qUZBYiHQWSjs8bXpMLin9+vUpQA/rUVZNGGN5QoZLDXG+FLth/Hcr8wSvihEcgy
zj/NiGLN7SVyrTibLyNpnj6d7orTcP0oIx4qh6vAN5m9wIzllJ5HL8iV8hiv/1fk
r2VQO93X0WjmlrUaNUxeM6wlGd1Hjyn9R0psEn7vwgeC6zgiRc2XZM8tUJ3wrruq
W0PaDfW4AGcXW/Qs/Lf9uN6oY2QGvL2nbSI95gXInTTYX9JN9uzfyhYRkdFGUU8X
AoNjPmc7YBEH/UxA1Q5alysxorUIEaTQ7gG3SZmZnA5Ka+/9pRW3aVJvExPJQdV1
L4iT6eqzvc0bIA254n7DlkUIcRQ29lsV8RBzWtOCEvgvtpnA1NaGqWgqAYI8IHLx
oKMTJILTS4sgmbME/ahs+gTDbOOo2qF3DuTueRj3pniVZN9vHLJrgEE9m69wRp5E
CcSocM9TmWR8T+ziHxSV558K5HVzHHRPNF8WByoDpAlRYcWEAEs787V8LKjjLnlf
gMb3Sbw5hKhIx5NZZLN5ONEpvfbnNPCJaYtgsISvbVvBH9AfrJX5/tlzlHemhdei
/4HiczfQhgGizlMcwWQljsPQkDrcrQeM8DwOQSKCDDucMzIuAoGatLKHPPPDBxrN
wuB4AwG+LOqJoQog4Il6+msYWsZ3KNZKlIEA1Dpph7iYsK7a7bMIkWBZAFG5ayGv
T32ON1PXuuiAq/ajFgzCnWE9uwOQIhkYv773uUKYfCOeqSyEaV+zZmt4wMGBBpnY
nztSZyaelswpMnIOy33Q8bSygDpP+VVNqpaYZGr3GTU34aRFLTjSAcD2mqDbi6qA
S8SCXwOy0DxCmmntbDeRBw==
`pragma protect end_protected
