-- megafunction wizard: %ALTIOBUF%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altiobuf_out 

-- ============================================================
-- File Name: psl_vgpo.vhd
-- Megafunction Name(s):
-- 			altiobuf_out
--
-- Simulation Library Files(s):
-- 			stratixv
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.0 Build 156 04/24/2013 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altiobuf_out CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix V" ENABLE_BUS_HOLD="FALSE" LEFT_SHIFT_SERIES_TERMINATION_CONTROL="FALSE" NUMBER_OF_CHANNELS=10 OPEN_DRAIN_OUTPUT="FALSE" PSEUDO_DIFFERENTIAL_MODE="FALSE" USE_DIFFERENTIAL_MODE="FALSE" USE_OE="TRUE" USE_TERMINATION_CONTROL="FALSE" datain dataout oe
--VERSION_BEGIN 13.0 cbx_altiobuf_out 2013:04:24:18:05:29:SJ cbx_mgl 2013:04:24:18:40:34:SJ cbx_stratixiii 2013:04:24:18:05:30:SJ cbx_stratixv 2013:04:24:18:05:30:SJ  VERSION_END

 LIBRARY stratixv;
 USE stratixv.all;

--synthesis_resources = stratixv_io_obuf 10 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  psl_vgpo_iobuf_out_h0t IS 
	 PORT 
	 ( 
		 datain	:	IN  STD_LOGIC_VECTOR (9 DOWNTO 0);
		 dataout	:	OUT  STD_LOGIC_VECTOR (9 DOWNTO 0);
		 oe	:	IN  STD_LOGIC_VECTOR (9 DOWNTO 0) := (OTHERS => '1')
	 ); 
 END psl_vgpo_iobuf_out_h0t;

 ARCHITECTURE RTL OF psl_vgpo_iobuf_out_h0t IS

	 SIGNAL  wire_obufa_i	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_obufa_o	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_obufa_oe	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  oe_w :	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 COMPONENT  stratixv_io_obuf
	 GENERIC 
	 (
		bus_hold	:	STRING := "false";
		open_drain_output	:	STRING := "false";
		shift_series_termination_control	:	STRING := "false";
		lpm_type	:	STRING := "stratixv_io_obuf"
	 );
	 PORT
	 ( 
		dynamicterminationcontrol	:	IN STD_LOGIC := '0';
		i	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC;
		obar	:	OUT STD_LOGIC;
		oe	:	IN STD_LOGIC := '1';
		parallelterminationcontrol	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
		seriesterminationcontrol	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	dataout <= wire_obufa_o;
	oe_w <= oe;
	wire_obufa_i <= datain;
	wire_obufa_oe <= oe_w;
	loop0 : FOR i IN 0 TO 9 GENERATE 
	  obufa :  stratixv_io_obuf
	  GENERIC MAP (
		bus_hold => "false",
		open_drain_output => "false"
	  )
	  PORT MAP ( 
		i => wire_obufa_i(i),
		o => wire_obufa_o(i),
		oe => wire_obufa_oe(i)
	  );
	END GENERATE loop0;

 END RTL; --psl_vgpo_iobuf_out_h0t
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY psl_vgpo IS
	PORT
	(
		datain		: IN STD_LOGIC_VECTOR (9 DOWNTO 0);
		oe		: IN STD_LOGIC_VECTOR (9 DOWNTO 0);
		dataout		: OUT STD_LOGIC_VECTOR (9 DOWNTO 0)
	);
END psl_vgpo;


ARCHITECTURE RTL OF psl_vgpo IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (9 DOWNTO 0);



	COMPONENT psl_vgpo_iobuf_out_h0t
	PORT (
			datain	: IN STD_LOGIC_VECTOR (9 DOWNTO 0);
			dataout	: OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
			oe	: IN STD_LOGIC_VECTOR (9 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	dataout    <= sub_wire0(9 DOWNTO 0);

	psl_vgpo_iobuf_out_h0t_component : psl_vgpo_iobuf_out_h0t
	PORT MAP (
		datain => datain,
		oe => oe,
		dataout => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix V"
-- Retrieval info: CONSTANT: enable_bus_hold STRING "FALSE"
-- Retrieval info: CONSTANT: left_shift_series_termination_control STRING "FALSE"
-- Retrieval info: CONSTANT: number_of_channels NUMERIC "10"
-- Retrieval info: CONSTANT: open_drain_output STRING "FALSE"
-- Retrieval info: CONSTANT: pseudo_differential_mode STRING "FALSE"
-- Retrieval info: CONSTANT: use_differential_mode STRING "FALSE"
-- Retrieval info: CONSTANT: use_oe STRING "TRUE"
-- Retrieval info: CONSTANT: use_termination_control STRING "FALSE"
-- Retrieval info: USED_PORT: datain 0 0 10 0 INPUT NODEFVAL "datain[9..0]"
-- Retrieval info: USED_PORT: dataout 0 0 10 0 OUTPUT NODEFVAL "dataout[9..0]"
-- Retrieval info: USED_PORT: oe 0 0 10 0 INPUT NODEFVAL "oe[9..0]"
-- Retrieval info: CONNECT: @datain 0 0 10 0 datain 0 0 10 0
-- Retrieval info: CONNECT: @oe 0 0 10 0 oe 0 0 10 0
-- Retrieval info: CONNECT: dataout 0 0 10 0 @dataout 0 0 10 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL psl_vgpo.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL psl_vgpo.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL psl_vgpo.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL psl_vgpo.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL psl_vgpo_inst.vhd TRUE
-- Retrieval info: LIB_FILE: stratixv
