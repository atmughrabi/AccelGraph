// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DGBfFFxxaL6pgZqr6W6kNf29Ykjtjziw9G8JSPMhfjHlA9vR9ppiqj+sRHZ0iT9o
79BGLTV6ikoiY7orCDg/YcBH+RKvql8EgUhZWkNHm5YFNuZfun6ekJ4wuy/xRyGT
Wf1L+rNouZzIZbxh3jPuK/tf/O6dBDEIpu4u1Hgb0fA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5200)
SmqUgIh9+zOHWSujWfx3LD77JTC1dPtiXWcBSrunaJO1u9rLQ5+/xO3JkfJbWaxE
PnXIgsZ7D7LMYhPYWw5A71cyQVWEkBfpPNqVdIUiROJQKVFNNa/RWUApixfr+zRU
t4lDLBqsOBNzlA6fmrF57sy045fiOAKr+TdnTSDablqOrw1IvH01OzoywTLopjER
t8ZDC7EiYWgIHlfk9QBLueB1XofebbU2WR9Wwn9U7a1sSmIj2ishvTNkZgoIhKZM
wHE9LkNhTG1xlaSyxOyUIZx0uglbKJlqtotE5wbDwDris9kO/ROfDGPSQvu+LJTb
5hvnAGXC+IszbES9hjyFR95Houk5djZnhQ1G+4z1Xqfee5t8+T1BW5LXGqV9cteS
CCfWlYHsDW4Ib8AvvnmqbVLujULgnDEE3ycqiFYMb0yaFIvMWnlrADoEr8PAYp9t
/Y6slE5NeMtVhDHcDF/rp43GCOPPlmThs+HoTu9RXKRNcr6J0RcsrlGaaVYyouSO
wBzpac3Tl6UDiDtjIwKfRwTd6ZbHwvOBIcFTKm6zq0NdYmu9FM0Ix0gT2GuI1NL2
sIWNFw0k6VroH+I4wsbWexomrWBqM86udVURALpH54cuvaAjmMJUYiy7VA+4JxYD
4HQt3aWPiUHhB7NLj1eHLs77o2DsO8cmKmvrWD3I2y152H9dZPsq8CwCakfL2O5w
DMJwKEpOr2DikaxckRPDhK3OwLEmDI7SqBpp28gjveSq+Eve7USAQvDRq4y1j8Cc
ojfpq5FhYuFJn/DnqHtWs7yn0CW/AReJ6vUQven91RNRufaGMNPQOh2BBAs0JKmB
i5IKrmmp7ssV4LegdqiJwtq+a7rhoPYxWtaqIVFIPgz3k9wY1IK4lVO6kyyBHd+p
MhutH0Vz3Q3keJD7F7fUtLeODEXpAxhTamgRtPgU/ALWPcwm2wGeze3DjYl+DEhv
pNC4QoVu00T3Sori4iwyVgz2M2OCDRlLhaVOd/FgqDl9Lr+2IGlWKwevVkqxpYix
1Sxv0ilvPQ/gf5Oc/ubr4h+HMqkaEfMaI1S8XU8gPP61d7P4hFi/b4BGiFFtHT9w
77h4Agy1n0TPqyXKqr2Q8kjF6nnJvg2P1DTpr45jS+NPQM2leHVopyWiknfj+zjg
z1KjIj1fzY9pdAo+UMMOxnc9NiT8sqPrh+VystTt+pAawRKCE3o+DSDPGfxDA5lR
8ZShuLnE6UQOtiv8nYprpiomGXvlV/DtKih/Ld676a/3mSA7pNQEMHIAfniZq0a0
N6XtgVDxehkQi7JuA5bVJVH6CPTj8ZnUHfc1qMIz3i1WcQgfjMHzBkIvdUGxgV55
v5XCVfgBCfsCwAWupEQF+ZFQy7rMr+bmCFmvDWpb0ENFHa27K7JxqfGGWx9c5Ard
80E053BW2ADt6RxatmDm0i84GgD+f+RuuO7QAs5Wzi2G3ghACTla1Z2QAUZntBiX
65j4CkA8tR9ckLnyYojizSur0jpl6S/QCj0+CwTgQUP3/5xmkyCaOJajk0e4bDZo
lY5wvumqhIOCBxQuw65MioqIdUCzW6CZEozuXD0GzvKq+XQTr1z8v5haR33l5th2
paQAerDaZT2rOGFPPo+q2puG3w2x80HJP8JKLc/elYtO7B+dC7ZBA/slk5FtChe4
VmU7rfKug5q/3wTvufiVIrDwgBBtLvYgD9STUwMzVvHZv2Yu/oHtKrVxBvjaOpt9
DWA983D/0nXTyIvaiXJj1sJko3HG+XD0cqFihZTZppSehZ0WHE9k/k2dXhqPS2hU
YWL1je/SflGCnLr4ExLuFoNU3q7PADfdpThHevEKrnic41sYumGjs6bF6pBhOIzT
1S2tEODSNHh+gHjEoObV4NMd9WjEPvWztiZhSZUxQ4YU92BwZk4Liz2BGWBPU201
1shwxHwVq+XhdnB14uGCtKGi+Cfvtm6jyBwXQ8qVkQor05crmdbXwL3gAqmhGPfV
ysLOHWn9KnZixDzQ4ppLpEl4spLoyAeHGSfCE+cXNLvZgO5dMHOY13x7JYA0QVg5
E2BaskeBvJC+mnRAU34AFpI7KV7mDzLmqnY3hzbHgrly0No1KV/5vmcnbHPlEzQn
4D9yqAq4Ur17yMlpB4ng01nCGeaZVM/REiWnxkvcNHoOhYG5K43C2Xn+wP3qxErL
NtU0gDJQL/m4I3u+Tnku4hQ0wiRGGgPeDd5JoBh0nWkCLKdAe8Pd9GS7S93SXE1T
78YqejiS4QDgBDca94BF6sakG/pKwawiToE2iiEe6hyTrJ+lZQcz2/TrM+17Itvp
CwL0xNdRdRoB5gJHYMicYv2CNpPwOvDqMGb3QM4cepk02ufv5oqRMMK37EbxG3LM
kwDOM4JDhp1RW7wdEjdIOCEeMthePTNiZT5fTQ6z2M/fgx/HuVvNkIiw9ZzgyDMz
X+Ay++aMeGMMcJTnR396YPVfE2EBFISPOsEZXI9U6CJxmPIdwrd3rLnrGNvsz0CO
R2AZ8GyZiW/repWr1lIo8cf5g54wCsypMWo5cavV+pywvYN7r58RBVbKP4ufk4ln
3Iof5hInYqI4x2V61GpZRh0L7qOtwV2ASROodQP82UgyQSyAzQ44nx2mVFTcPMz4
G8xy+nJiDpcI4Tw2RgmAyTb2m24obwFr03+4TiMUyd6V8+ouJeYPrTPaQcltCjEf
90ouRdICtqqYbW1JNuWC90ecMOHMh3xJ0anjBUVoCNV1/WicNqDeqosdG1eiejLe
wzKxRqLvF17k8EpSVEclPDhWGOv0l4FCdubwMNva+ADXUo+XswtHWbjt2baLjO9/
w6inJEtkZJoS3L3Iqa566ikqAEqKFdap1zcagdGbAlq9VqhQOBoUYr3Hfg0YKyb+
nlGLpzp0krgYikqYLRgrxYj77HYKKphKsU4sOqeHCs7aDfLyCfpgT97VUe5bxP1U
hNtXhINOT0A0MGqUvWVztAlujLYSRH11Xqc6mSOcaMiK1LRYdzPlyqfMcI4EGJnt
2PrqZnEAnRr6r4iMOhuotoHz6E/JjILxSUD/U/KWBZp/pYCNggiSEd772BBkdo9s
GrUxuydrLyew/7V6aQiEiSjK7ZzDLo5QtdkmFvxnNoEree+7U5JKX39z8ENcTLQd
VIUfJQNFRdDWLVwI07zI5Excr1ob/LyLmkcxTraFjFefPmJRfobsrO3FbqrgSv5I
4jnE5cBm2NQI4Aeri5m8o2TCo2t29nSsD3uZS7FcUT+AoWABELTz7M4raz/yrHiM
UdKOQ1FdhZXNafxu0bwUTQ72lfC+h6IT+LNlY6YmuvZPbhG91jyybLRloqsL/Nxf
OS2IfTv3nuVdHptjdiNCP9i3l872aEFszUVvJ9jHjyrl6gXclUFhtI4BoBlwZY+w
zUbc5VDubwrPATB83eL9Tctn4SmZr8vBaaIXDaVP5UogAfoPFUTEzRnz/yjBYPwF
Cy+S/SEIr7EMBAIToGffttVD/TMJQp1ReSwZuKy3FUBR/StAtOkoqJjxRWidcNLP
3XMGZQ+LBbvxFTemdhmMSJxDMHXEH8/yQ+snVfgrzIUXSu0c5nUcMC4OsdyL7nYG
j67egGnjtg7CaiTFceKeKAUu1+2WXEFbnNwVVKxtOm+5WtoJdkEh3F85JjR5GlrK
G49wKMbI0IOSLDuyzzAjtoyBpcUBaAZG3sHUr8qkukKiVs0GI/M/OEdMOUEG9OJT
kbEgAULgs6EzubnW8QCpYRaFBGbbDp3rIuVMsTpthkHPs05Lmx8gnumi2JU3JG67
lzRwamM0wLJEZTJ9qvuieJggeh3gQiqMCQ6IJXZf86plzH1HS3ZF2akDhJg3ZDPH
ooT1elT3Nxelsfeb3tQQwCnoHfb/D0y9o0yXIA0HqStk3sNf4c9kEutglKy2pz/c
f2ven8zgdHj5Y/1oe2fp7R+j1ERRQipN/IP7+nHdNTf+cZzzA6ySnP3zwIaOE01r
0RfQQTTyG9VAIkF2BhTMmBDh+XT4FlsjMXxBgK/DUS04I6AGh5P11aUTD+Y1UjRZ
yh78nLFAIVM9d6swupTlitCv3B8w0Qkz4Ir4FSd1ckIlAwW5Sfajoqt3W1NBGH4H
Fb/tqt36EsJh8ogyntfdyNrvY9QXZdJe7cronsXxk0c0haUYDWlGTXfFBVUqgqJ7
WIiXwnCDiJSNL3z5LoC6s8d9OsoGqp6I4bkx1hGFjcYmfqlwwUdZLVqAaSH56YyQ
tioiKyk2Ko+MCR2nt5VcYeV9nMziWiLJubL6Ub6JHF6DSRGNsZfKGHMTjd31osMW
hL5vLg7oMZYyk1OxXXjlHB+eNCHUnBIm25SGI5TI2VJJVlxXJ7rXjcQv+9U4jSzg
lmilsSkd8XHOkmL8okNbU1nXU0UUChYlQ2exReZ8pp7SWIk/To9NKs1k9XhRpg3d
jBYbbqElHr2GfXCibkb28UFeqp1b8mXAGS4jI2jFDgrfIE2qm+rJKG1VUwa50b5m
ZHzKl/fSwmJNy60Durz7ogjyk4993H22mGVnK3N1f3lteCNtGxz42MF/mjATdI5V
ihKbNJ6EOQcR4pMbUVggbtAdtlNz4Sd41U3faxON/oH210aopd0Gku7GLafighLC
M9+8h4RZSoBqBdmoAiWVLDBHNxWgFg/riymLlbtHskz0FNorY/7SiR1IuIro+rHg
ZvL1Pj911kQaxGSJXCm/xeKnf7F8KRMlp96neClMprORrrzuvumYHvVpr/GgrwIx
gxwloqBOHTywLjTlAGhOUfb1ULPn4dGtUcyr20bNJzcb7j7QUrSS38OKoAZ/Yiw+
Y6E7auBqNh816Rcm1Mu/qaMztRb2OXfEuoFrJTZByA1Aaj3h+ddqIZPT8p2GEIPe
+272cfmYeKMNUXoxih3THm+LvdG5pM8akeY9FLvKfUw43MvqDRZJlBt7Mxgk+iDy
Gzu8un/vVM2CXy3cIJExdXD2vrntnk059FZGNKspImNWcKS/2Sj3Zy5fP6lCiDyz
CjnaANiqWcChZLegQLyYt3wW4XjzQaUY3bDV8bJAMKJraYLtbjaIoTGPa7dPNMMd
sfKVEEiC1BhiaB3ybPow2nDv0X4xCuA0NuvqZiBSc75CO1G8nhy6szF8ys+kLgQj
vfYxXau9LIgoxl2Vc2oUSS3dCWqiw+nJ/J2/NjhQ9YW55Dk2Alf/6S+Yh1vFlMds
oeB4qfPNT5FadEGRkliqPdu7vO4W24/HJVyjvRZ7NCU88AR63fr80Kv+CnbOPt0B
WO5qAeZBrHoHXoFhBay3Uq4zSEwbr2Xs664vwh2+a7BySuwXwCPfP2Mq2y28Fq4h
O3oL/RHc3zPhV8z+M/Xy3560ou6ZoI7UvEHWCncUTddAz7rMtuYSVgau+p7wWokB
pGS/UpibudehnsFZqNew8TwBlj7sK3vSDK/hZ3Li9GfsKLRcYV6sdV/J9wBPLYNS
hq+8rIcv4778sOue+rIhd/OKXzheSIzgi9h6TAi1qlmrBnPXbTqzcTXj0e1p1vZ2
CvpUFR0vKKHq3cYH8pH5HuqkN1JUrjJfUOkySNjIkgV7zmt0xYdz48pKgT4Bt6Yw
iMIBk/LCgJ5/MzjnSjvUV1krEmTOV3K8P81f1GxBcqbDPLn7JR5MiTIiam+LnKQZ
HmhoHXW7BDjKxkHK+9Mr2F8iiMhurEr3eG/RUMU3HxUfXqAgfy3ZQICzZiLUEGpp
n58YtBlWSi2fDVKSeaGBX6N4kMTzhRe3j9lB4LhvZVvXrIJ4QLUvF6hsIcQ+doPA
zheA3fwHrxW8TG9sp5+41aV+NXaauAdEi5Pngwr4hDHZGhSapAva7NDsD+ClkVe3
z3f9o3YvrnxrzdMBThsd6Kvt/QnqUdXdVxqEypkn6getdqQHMiBxh1kRfWgkXwM6
qrGVpD3KwKIw6o3UCeTzzA5z1pW49DAhTvZoHwx2GgrRzc07g5DPbxcqaTqB6LCc
JGO7h4Wv+CZPI/RllbaHfiiSdiwK9NLQkFV4C/KY87nUbIaYJmXH27gq02HSetkX
uQrkvFJYdF5PNrT8ckNL6EJ6zF5GF3UK6TWF5ZUoVvwCOsTEvkzkoICHfukgDmyb
dOQrawjudI147o52XFgasndodj1qctu/QR84pehJU7lYxdmgd15ZtUl1V3PWtvmR
QeMtZI5O8ZjzfFajTbcRs6T7UCkDl/8jedkodh5MxbRrqSJbWxH07SDMUgaj1VoZ
iWaHBQgsEAQWnnrEk6x00Ds2LQBC6KQg1ELb/N75/0o52Y+aN7TQmeN3VFxh0ft7
EbivYI9qerBmIdSCBr/c0aAQObtZXKvHE7QMW2Pc6McCxOTnxB9f1LqRIb5WJYuN
VsVt7tZqtXQeC1n3oa5m2R3Ld7YL15dXoGHQ7CyQrgpw3Yy0xpHwp+0pt5pjRpqn
rl5GyWAJvOoFdgBUDEftkjzSqzEJvfkpRhZaaigcMrOKOFh/wHbu+H8c5JFyAifg
QlZWV0blP6WhrjQpXSwjQLGEUOjZJwqJXLYb7ZY2nkpxbAdM2nrFkHEdeKgNqYoD
Y2o6aCkdkNv1q3BxZrHXnzvIB0Jp/2A4IoCcdFDQVNT2cQeWu/lkchEaCni9+nV8
pmOY3Qd1QZm5vYgM74oT84UX0qJax6HPfZ3n6mTLe7OnFNX6XKEF5BgWd+4We/3D
VGZbWOqmZvHKztKXMHx+exkvmfGylDJ6sOmbYJpWpEzmdoTOm+mVmh04cN7nF+zS
MVm5Ih3slxaxk5Nf9CBxdWwDMbxfIwbN3SQC5u1+evL3eYFCOfgTKDnM5/dqh/4N
+LJhxjTmvGHmdAekRTVMwhfy2+o4Uo5ZRAR7ihNN+JZubsvKKyuQvQBfhO2e5Nd2
mLzqUrL48xYiOvVCczyWhN+TVAW2jWqpGlrki6ElG41Ge4F03Gqwfn5tZJrLxxGW
syiB6WXPjDx9zD74T9GA5g==
`pragma protect end_protected
