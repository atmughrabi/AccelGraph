// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:31 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
enrxuCaN+k+C/xpREqdkavN0O3dnrzGGnisgRZK2fVeGnzQ1GPVS5krtm34H64L4
nHw//38M2+Nk6DgVl8TpHzeHziBBZLrXdwwMtU9zb0o2gf3rszRDBd3IhWe2Y6++
rRA7QORbaBHhcbbGG8s8BITPHfjBoP8XEmje15md5Bk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20352)
hbAnokEW0T+iZM6cqqQ4q76+SxSOpyj1CYwNsa1kdjCyhIwEW8BLJgC1GLvgDfco
71tBsZ/T5QOQsBqxahlGb8C/otnKR798ebMhxM5kEY/Bym96f0r7rtA5skEDfQB1
ZhkQKNdiUcvNOEEiM4X0j/SVmnKhYH98aqpTp52fS7aIkxz+Q+h8Lj36kvCcmeSM
6QMrPn8KkLdDAfnBNbgtKuIhX+wG57z2XKJszNFhgzyuBK8TOcdxgRjddKIXszu2
umSBEbEHGJGm2IgQrlJH7V9Xvp0VsReIOHBjJrlr8XnTkNIMp+qeyDM/ehxhjYT6
oD7Rf9/laUbBThd6s6utIycT0kCFEfjVwbf5EIrCNazvZBS03DJmeEAQ2kofECef
SOwZhjid5I1NtFPpttOkNjjuxHdKGnVbEeS3h0q8tzKaTSXaGCx6GSOkkU51HEoO
Et6hCAF9yHqAXdFHcxeFzlsWaE86YOyE9FZHa7qkvL9vHuB8udlUxFqvKTldcs60
mejS/gNMV4UcYqmq7XkRzC8AjfgzRElPV8UNbUdXS1ib1bf+hT/S1dh6EmWsj1yD
k6MVgL7a9nV4a8H2HV3EQDUeBPomdR+DoCmCVgWlKMKUNCFnl+Ypd1Qig6gU/qPC
sBrIgLKeKa1nFAISfgDOlL+AWR7wu1aHF+tmGDih73ufZfsH27pjmTUuYiD0Ka5M
aOElcJ1KIPXDxNrvHlv0KfxCkB7jxKrCc8GqhrEprCoZZKfkFz5BvnnEsPFaLAYY
sfZ6z56hbpa+y9qYyjy8i99vsMVPrvZEsQmxHtgQcVMkw15mOLbQXTIP/WAkn10W
ao8HlvDk18QyhE2Dckq/m5GEN0QUnDrMwwXNie43MBcr/cCe98QOMlBcUveLgBMf
XsW78yy2IrsXPuEnUfrUP93VojZWmam2+7vW9UWK0452UPUr26BshBZ/rDkWP6Bc
bS5SZoWTEkzd8tkX0jHsEwKPkobUAxyNv9xkQ6hyrAXEyxoNa+V68XJd/Vyo5M0W
lNxpb7xPANLd5KNsCzbPLx4AnBAdvqb+eb93QzoW7Ttf34GrcrM/EoYDdvsYZRTK
4W1kzMxGpueo3r6KCTKi1r07imptQ9ncAvIzaOkX7+PlIrgylYfRJScAZeaW8+Nh
vKdGSENDQ1VFS0jA1a2Gb0piUbWwHJGfhBF7I0HZErjTNZua03pKwqokPDuMXzMr
X7ktZjPUg/PBKOi8C33Xz7zqNUQL1Y9uSYkvsskdSb1bW28bfaKnpzlVdRnva9bI
Ja5JhsDZ5bjd77JtyfspnDqxRZieMCUqCEbC+DpHZ45u5JoQl5GuJhVQoWMJsr5x
tXLAU/8vxbuPjMtPaPutAVODNbvbt24QQWlqXNbNhdjzcPqD5RS1D/uw7HEdKY7f
ndE7y6oJ866+AEp9FgkxM5IRBAVWP4avkwEGSGZ41Pu0r3kb71/ZWwcQ9uLs8nNT
AqNCgFKENklt9ZOlkCaLk+RtoVcpwqJkjkkzqpvC9KyKKrMbiW+esTo1pCmfWvi7
XIhqSMcaIFO8f1n4SBA8FBQTbvivpTDBDIcyjSpPudQkp0EhwuQRTEckGGNfJIwf
lPq7pvUQtKAQo2vl0X+c+9zCndrYBiyyA2Ze35d21txFOAQIR3b31w5vpTfCcMuG
S35ROgUPz/kZbbiQcFT+soGo8lB/uGNrdEtL1go7EFlqiauBlknw0Z6BytureZ38
ITYI3ExUQco6JjFmpdC4/TtiWIqSi9xIz7OKbGLhthyJOZRxcQzgieCDjlvGfRDh
BuzePZh99VcBdxP3aGHENqNJHV2lvdbSVAyyVmdBXYm/VTxbt2AEesbpSqla/MAo
9mBVnJMrLxyScTd8gkvp9vrpQiXBHP9iwJlkTLQ9ELVZYtjOYA8eamn4WtvFyux5
k+fq+of+tYj5Ulwi8XxLV+75BozvRLSb9bZ+4lH1vodQeiT0hHPHEyHZxzbrOzGY
x7WHK3i5wODG9p8jLqBGQTpp1v3sqAKcWZoUCG+3pze+sos14mrrU/ByUKULiNjv
gJGZta9sCAHdvoAJREu7+aVMSxfuHcOYqSJrpmEqZjPap3+HpP3KJ0TQgDUIOHPs
imFR6ekurDzigaGm5sZeVqrjPNlNWQB2n8a+ahRX7Ro97AVddX3pKevjB/HBiKnE
AZffyScLXnGlSgWLbM+JWNGbD0Y9yXTSgmYCkYBpWOHtUECFo56ZX2UndgYCWQEY
SM/oowXa0MWnIcHe+BhmbvcFgLdWtrCwd8utOKvmSzk86JXjluR+GyKe77Nqthio
IgnsHGPRkd3y9Q9xW6ZeBEfKFKAOUSEIo4q07IHx7XYjLEFQlFIXzvyC7VAhPfZd
ljDe4Aei+XErVZIayud4ytvjwVthKfmUp4pmxqkAnO6GVFL0qapBDUdchb0pwHrR
Jp9NcfTWSZovsLZQo/YaImtz6/Lyb3y+DZgeTGeesV/SkG5Y8ZptuYMINCJDdZCI
g1WX7XaTe1UWKn4HgP6TzzZz68UWKDFOJYPNe1U46yY70ide+IO/n7diygWAt9k2
RcKJM894iXjoWX3yV+lNTV0l5QHSSalbXApC/xH4sg8u5hi9/4ZAh0R5DYCdIw6E
in6TzI2bO5Z26gO0v33z3OrwiWc1CIq6pVcOYbja4QZVpfRLrU5uQZv7KEUOrFOf
mTXpFOuwtnpL2xhCoubc1XeiWvqp2ciFDF/7xW5JT+ZnMN+1BSyh7zPIOKOkBysE
6lucDP33164jECFqjUMy7e+RqBBIXyjnErn3XsAfWTBu84pveewdZwD2YrSka7FD
zeqFpS62N129zK9O4mLPh6IIQJOVhGeGliIXJ6baGUL9DgIRwJQHiyqwbEe4U0iN
uYb1uXFG32F1JnzoN/KA1ny1qSmSv1fPyafu/yf90f/dF4dK8u7v+ugq7nkj7DSL
vhA/uBG+7jmgbPyIClrejt8E6jiBqBQTKm0E1fKQWP6J5uekPj2rLb+VrbAYb+4w
xD2hWS1wJKZBhsHRgvQDAXNe4WPqQ9tAsc7N6gan5MmVDwVb84IMoJdKqqrOvwww
uxvWK8f7rZP9wr8fipqB6tvBBCFrOsv8DF73ijOw5CbB7Y8sfgv9vqhsK3ujk6xD
Dq/ef7CtyOELxf3Z8qYcFqNBlacZ9RpuPKPgU6kuA7H2hEtioskCuKLsqR4O79sc
lCvUfOW/WzQxWN58wUl7rTLpKSo1RrEFySiWvTKXsOGe6Q8NJhYNf20OvihjBwKm
EehdjxvO4A6svHAnjtp0V+SX1+Rz6OtPujUdu3N171hyDXmhtK64I4rQTEYMk7a7
0u6LZJd2HeChfjmIaQatenKcmq5VtVoqAV4ZpNFS7CBDwnAsZH3JwrLZpsFXWFmt
P+z4AAmoVFIBcHcNiV7LZFoeUxuqi9CccDgji5RR208ZcGhMDcufNNeP5x7nmNrC
lhWhpjz5VNeAULlj2YjX6JQ3/D3jm+nZ0wL03AzupbIWhG+YkpPL2sxbBmWFUsdT
yybVSysIaeBWz9atp+ZvPCaPNZU3xaepN3pG3ZG49q6t824L3I+SGcFTw8jHF72i
HEgZgjn6kn3z7zl/efmFYPgwkmP8bH4guq4jnHOxxU4wJfBdBYy8/CCz5jXLVTyK
yh7BR54dqTklz907P/mDqkxJFgb6bDbmr8kkIZzGPA8BKao68EVcybi9YxLUFMwh
eAb+RGEIWHhBG7g7IWx/C9tAghVfoo9saYcuMzWokRhFHxgxdXqlZprm/ORWmyFC
KnVP9bK1QbiRbQB23+8zWchnB9G/Q6AcNbEOMp/pPkThhlBIzp8jbtaEDKFrTFfT
2XYNF5iq3X/F7IgWqSqtuy8c6K//FHLv8AcVPlFVdqjkli9DzwyQlBA3KHX+yVFW
klL6De8CacFfnolXauUtP5e827GgD6dtESnQBli58brLFwyOon4uqwIWUIOxRSLs
gIrAhmMXpIB/e8IyGlcOK4OUOOddYP+O/kX8fgX6yztAfQHMJcBY5Ng/GzkbsBky
mz0daCjJCEcyoN/2tUWz1qUD0ZN/Aq8vmDqR8sr62W1Pqz5low4WsJUaLFPTyJv3
Wq67euOSaLnqbWrk6bxyM2guKqH6EFdaFPfYl0jsL8ydELMF5NlNKuqxj+vBGp8s
d/U9ei4OcH/mE/ZFtDZuBy8aOYelt/CjDQ+DSgK8OgojqQn7s5xu1+gy6cwkWLuz
lQB2rIbT70V3hPTfv4eQjhMAng2ETDiDnU8nCLILj32mpYbQAhKv0aIQvA1ELbbq
UlhLzr2dtK9fp900/6s/3Z7DTzw1SLDbMKzJEPOJaf24JHuzRKujao/3vZULEA1x
o3qYutqXoOhainNgsr8eqQ4I9gzdemKBpIldJQekq1Q8ZKUbPlPsX6BbIwtgKquC
hd2CY8i/Oxj1rYEALUtlmbfftmP9j9j/4f39OWjZclcyVImgbySc6HyWD0B/yExn
HEP2kyQ8N54h8u6q8+lF2EXUkHI9bo87quyTHM5O0uW9l2xES9SKlclD/k27lmLa
X1OMAf8bQVdVeyEDlGjlnPp/oVVVSp8Yr2a9iIBw530JPY5pJrTXoqBQ4xuptoBG
kgO4skqijo883twuiY2yOPwwQbkXhCsql2L07OcF4Jwzaz3bvYTx7TiEZIcT7mAH
QoGJVuz3grn36rW+K6CwfIv9VSyp/kzMIBmK2OaUK+PoKzLjLKjEyRcjCSPoI73B
be3KdzzzFrCT7r6aOJiX7n8fp3llevEF6F/koHsl4mSGWcRzUH76hXi7SVodIhvc
xJPH3hhzbdWAML5K/vi1xRhLDKLevnaX+u2mOd52BeGPABtbbJ+moWRvozIq966/
GoLisjP1jn/oDof/1CJFP/NkA0ZEp90BK5SsJvfpGEfUB3S60ax21h5Gylah8WR9
cZayGy5XYz00VZ5StG0VPaNZK7z/f425BtnI74N7LEaTptOLamWuKblL4oZvxbVK
O6jMvQEBD+d9pPsRRUhrcaK7bzqMNYjlksS4ldUn0HgXVt7QSVx9FqozuI3ElBuw
n2/JQzR6ST6hAxKMb645La7LD5A/nRCQLIWhCc+Lo+1q51+s7QhNa3EUieGeT8xz
fHsLHeNZ6SEB8Ow1K181NUqSk2EJ1zGr/q5FfXvBHqslhjQoD/zSaoqhYozkaBNI
bPUlzluXfT31DJ2V3hx+TKq1Cpk3aXKUF6+/x7zDiLN1SL/lSok/oP76T97gNRO6
8FrNHbLd5Au4SjwHqCmYUhnNDj8nMpjPmU4wKWnWsq/WdRdTdnr2twKXSjwIV6IM
KpOva/9UXXLLeohU7SCgUmNY4R7oNQMK+snX58IpI4r/45+vaUCU+G4I+1bLVsZp
WxgbOLYiEiaqv/M+wJ4YBDIBWKD4HVq8pefMDICVNrctOyNRmiHHaCr4qoEHlZc8
M3pl5v6FyHHjBscxHQvgRv2GYfWWNZo+wTRuRAFUUORPJ1ZVOTb622MgfyopT8F5
3YoxqFgiptckqNryiOD/kUv39d0enG7onPkcycpBH2FitSE7dDpwsF1VN9VgIWWz
6F1hmAJ90POM6e8pOQV7ZGo82PVkRnKy7SEHfkTeViX5f7XvPffcA4IPStWblsz4
qbqLygZYU+cjX5bxd8YJt9IxZrlH9HLS5KKer2R+epIxDzTsBfGkzBIvFZakTh2T
glQ23BPEUFCS5jSnJYTYqC7lbsW2ScfsfvtmoWJvCRE/2N2/cSffvPYb6J1HakmS
SalJxfc5gLsLiAdzc9eov0tG0iC2hpSMiVhSCJopAr7AVh/095tW6sfRstFRNAUt
AG2X0gRJXdwdCdLxU2P80BWOXgqsNTW4nJMvvrMn37OlMw2WXZiiQFIzURFeVrN1
O/lQw4sWqPovP76cTVpQIG966tPp436RgUoqt0snna0EOyHdu0cvOfRjJ2tfZODg
k97noDG1WtzdgOunELSh7fw05e4nt1NoO8kS1FXb32pqHTD42257qMNHPhcjf+ap
NJz+fusCdNkHUoW7FjNP/GEtgi2ckwbiK7YsvICtCX3LBsWJPtx5cDdQE9HTBh48
AWYHwQ57ybbeG6KDq5E6DI8ihprfFMeDIK7GhyLL62NIH+d2aZod72+nNzdXKZVb
OmKDcJZFkgQ/PIn/SDuj0LxxjY/lm/gg7lUPgaK8GYVSSe56T21S8YtGiYBp7I/l
B/7UlP5Z5bPRMrA6a+92T7Q75wRcu0SaNZfaprpIsyObku51sAKHZfVONJZ4yn02
+QamtcxjHswlToUAch5AOdRHpos36H8WAIC9ltnT1++hfhkYqG87oegysKosujfu
i1hEjOODHW17xVSLYNgcPPcmFPJ3RcBzT7vZ5YfifAXCfme1GBm6hgNj6lwp3moA
nUGT6EvmPz+iFvTw5iCM8he5pgrULzlEYpi/YIZI41eWFDtJNz4voTfzb6JxPhyO
DaOvNSU0So/LxwKVb+fjMJ3o0otLLj40vTxrSKXyvh481BkurxEoCuZmbMuZLxDb
RcGOMOsmbHdmxUcPu64efK8MGznB3ROPwiCGcJmxRWtwyQViaLozLbZLeNFeLVss
9OLHuDWoETqk0k1Q4cV56G1/WKOUXQ9VKi5WqS+F5wYOOlNOOUq8p1aI+KgX3DI/
UKMxtgwzWpwqhOHChR6lYqt0Wipi4zKyYd704vhI50GdP6raZ7YLKx8bqxs9bpfF
DIC/YT6QE8l+RFNrkd0VA/X6elP1klj36kMHXk0LQ1Yz7FCUxvO1o45J4X9kpm40
nE84CgF10PfdlLhm3HDx3Gh66V6ItKi4Gh3WKt+xaJq4urHvdQSb1DyTJPse7jmQ
EImAglOvH3EfcxdVkI+xKfrzdytDoKpXaCm7/QUjPhg2NVjTCyDo2TcwYUKdnnZD
If1PdxZc4Dc+G8ogt4T3vXX0Mt8OkcxHiXdqXcX5m6HAFrxysQH6V+JZVIbhxzv/
Nej2Mgs+Fxz3mXkzwoF+xTNWhG4BB3IrBwhlQUf3huGwvEcldQbtsQa+XnXJ+Q35
UqeenhpDL+K2ZxYI9W5y15/577g5uoUyDEEcly1i8fwwSIM64uBGZMIW408tN8KX
mVw6zjyE1CK2UobX0eEtx80WTMAJKlkaCW8Lk6WwC46IGeKcbrUNiYoH3MBUDpI5
7dfjyZUZCbLuu/5cs2nRWCJDoJt7azBVoIGiQ/tdoiCCWypr+c0MEXsIHHiwoxyy
7eDGBp0mi9jwwJ0ykd0tSvHnZ+M7+JvmajCpbXhkzF+LZCspcQL9u/VJuFxGP1Ut
Nc7MURzdSkrmF8vzwvjykpXs9L7/3SiNhA7IZ2lWsnKwbmfkXwp/NzvyRn1Sxp6x
cGxwdFZA8yUCerKC6ql5cEyU0V45/5BI+OEFR6704v9PFQFIjvEPajYPr5IN5/wn
2Zb4TCr6JUVWT+7V3vt0dKA5FqLrP5yLs+hnxYhRMbCjFAbqZaHQ+SgNLuR4ZB3I
pRRIIxtlE3b6ik73F6R4j1VvI/aWZS8kBpBMMvElcs70AOgZ7m1tmVK7TCFsBXwY
K29tlVqHcNRy0Ud6ZxmslM6HjsVbb/p1jpCICOVZFaRPBrTdmlmFnxJ+k5zN7Xaa
ahcMwMb+MHwT+7/dG392tiPrQP/qwy8vrbZM3Bp41K/w4eaG/FzDQ71h+UsWI8oT
Re7iKTL6+rnmw9b8pVWU5xuJGCcfRy54YniVAFB4im8Aw0OTzKm5DpOp9eTSpW2H
smgZZmTo49E2/HJF8NwOndO81kpKQ2UE1F3/LbwNC6qCCpoV4xJqm2gKqALNVuVN
htQsi8DUfWmdSozbwNbRoe2sBz4PFhizb65OI+Sk6tdRArj/61DtErZVSCxEuVT1
JpUxkTFZ3KwpXDQilDekhBQXu/5TwZgjx/xv4gnj8nU1Yt1WS9Ve9su8pEhzdZy0
TbjAdUdFQWcD0h7pqpz2v12WFvo726CBSW0gCtEWrVOILmP/nLv7T1RYXtmafZD9
nn3eAuIB97BFAbDik4S+6rD3hl+5xoqirk0kN/FNpDbZQ8kF2DH5+ioWd0Ezx0fd
rAKrUDUCY+0F2Tw1BPoAtm6UaBMVeZREm2+eWL+QWwY6kzbM3uj9BpbW3i/vOxoi
xjf230JEi4V4O6JUusFGChx/a2sXtXitK8QU0dl41NxdQ/Tb8iNmBrZp6/yQilCS
gvzoIBTGoOG3ljlVAsZ74Xbzw4DFFXKJ2rBonv7j2NWC8zxXIxBK/B9LP7t+v9IF
s7lTEBG/hBpq8S1tjZuLDM3BMNqrVQmE7yPP2iweb0s2oxE7V//XzoCYiaWRsTdT
rs5fRSHUx+h+QRQ6oEoGELMJ+3vFDxvmDI2MfQ8nrnY6zaUMkLr3FHndTIhhLH1N
yYARU2zvsorToVIG15p6gMUoXLbG8gP9t4j8SZvYS5/2o2YsZvfq7cvR25qDlD97
wH7KiHJpej8Zz8pq/Nx5ZufVbgWgXLpBj5R2Nor10KdNEojP8YEjkpliBL3TG1p6
NFqCqBXFPnd6xWFt7q/PKvb/3gH9FDCUQaiyCBvz/M60BmiBkdLYqglGhH3xqJ7z
U7/wEnhPepXucn6dibKPt1vuVkt3zwc3cSr7l4tYV+9+Cfdu5rvmc3aZWxWQ0foL
sfouE7r7p+T6pMSSUru0P3iEE8MODbIltRnZs7LV2b6Ex2bAIIgvGcQKy+EsAREJ
s4o+wlwEiJBBgckwU/FNWDFpBRs8SFQulSU94AhPHi1F612jSNn26716+9ObFr7m
aPdaeP20H1WDuiy5VpSmPuEKP9oUGacMHb/mFfbb39rsY6Lg5/2UpaRMJRhUxlxs
//VYGvXwpcnl96LAdkJnVE4CFS0ILCFNTX8knkiCiaq7pjJmEuNGSLkIwyA8EhVq
KBpTmELyewaHsXoWXOxc7go7joXP/+JH+4bPDSf79HbMCf9m/DacJeb4sJeFoPe1
CMWAWOfuj8LlbZNBgBiPUwgnr4HC0hA/OpilNIMtRrQInr7hGfyXL0Qxkd6U9Czg
VCN5xfcCksiw5GfdB82dAYTiMjz6I8GIig7WbOcMpeZ9CJAYA4UTMn7v3EsHSylh
LN3kFz/8v2A8A5sR+k2aG8m46blNpV7aIGWu1F1vtzyZGqENbH4TrRbWm7dauVxF
KdL874uLpQUmAmCAR98H79A8yxTuP8tf5g8kr7kbscwBig5IJ2ePSKGmd/0vRuIn
DgXrWR5vFCHe8pSBJznOAwSOX1P22s9C8r3xGoWP/NAGaULggNh5iG0nE7pWCBCT
JmY9bJt/94vXD4q8XJ5dKQxvaAqKQUpLpe1YaSSyJXUl9rdzzsYzUdm80lnkXLlo
YpgDccQD7sXdenioK4p6D6r8dWpFWhlKlBluPwcQk4rYh1zX1bk2grDDvcpS7WEr
jQUoxLji5ecYD0b/y9QVas4MTF9c6MePzArRZ028PQAld5IFpvi5oF2h5I2eAoTk
LZkBsc57xtjLsFOPYnOBqJC4s7ag7pe5Fkd+9mnPAfrGqq758uUZTO8vybIq7Bsa
FUYoG6F5KYIWdANFDd0hbKmCf5OTEWTRA6g1TCT02SIISUwxGoH3meMkPH8tz5o7
iJ5I1lWvLF6FlyYreJlfiixA8bL1kPhE+5bQmFjeKYLyHgU+gan4RS9EHtB071yy
mCL7e60Ky6pI4muPkoYLgksuSaYsxI0SVcEpjZuLwmVr8flluPRyaywQoRtcDloH
R629KY0ie854JHkT6498DG06ue78hRoLTBVeU4uoSDtvITqQ/Zy31vNMOs+K70Yh
+EhsGhZJVp9al7Kl+dQu9j90ck7DPhAFhaCLI9F2virf157ZnCPCP57RHeXcBjGs
C9X4xkAznjM0Z4LTIpWpEMEpZFdMMnnUtr0i8WJyrr8O+ExKCT+zf/3cFm7TqafZ
/nMc+3Hb9r8U2irrRDv3Kk5uFoR7pCxodIN+1uLVyugVZN2iFgfLq/Org6OOSszj
kYmeH8PRKGiH23q8J614nJ+rzU6joSc43Gmtul6YzptT8xrqUQnWEZ85Ua9psBvu
gnN6wQLtGivbToP+bKqvuuyKeMmyuivvVzG9UmQjau5i+6nxbAezsN7RcioIPUSZ
1ZPCVbexBlbR6A8JkcH9YDTqckSGoswb2JvhZK8ohTmBvtOcE1owZEA7msuymStW
qEmoLyJufpxQBLI5R0Iofv/whTE9tMgdFTP+qr36wxyiJerF6vFAZ5UZR0bG/uqD
BFZmrG7x+I9DYFyzsuk4IFGq/D9V92a6Q212WIJerWBxtI6xDRYy6CXI3JOvIrqR
cXmRTF94+n+k02OGl0+uCo0XlCo+af2vqUx6i8a6XtuWrExoKOssL0SC54QhqTD3
J8+doJixeF7bGRcQC3kEgf78GDOYDfZu/kEYJIemv/8a7qyWlnACe4He3B2SRerG
oXdWFsaicj+53g09a6L3ne1EIoL4ken5yhs8dQaR8u/KtyEjVIMrVx3uUHfdDiAk
bLCs1dVVC1pdzRtmtKe34EU9gXFpQIKTZtnjABQi0SPiyo3KHVhSzCMvhNhpwsut
ggsltafEpIN8oqwCqrNSSzQ4sUX3UDbnWGmIhEGPC8SD/5Hf9pBC0KEVDa02p9Th
n0IHHnfPbmJ3Pmi1VG+nGHbYwUKx5UVysog+LYenJkTMAVl0X7GKXHSzTBcZMDnf
13P3ScHxtENWW4ZCZ/3ZPcZTYuXAOo4kbZDa0JbTqFzG+dZpjumBGpHPc9VyHo1R
SQAx3LTCOSqCm6jF6d9zNT5W2CKINoOqZ/1eXz1WwIw8VNNd1b0scKeCjQPITVcV
ZNG5rmel2D7s/HurYYhc6rBUzgFgTFAn6TyqAHkC0TGFGjlxDb5csGbuNEmL++hR
q9T++Y+C/5QRu+iQzfeNHLngJuOe3q896/yqET8ALWx1jgc5mBGtI+e+aVBtJMXh
ECaCX9iMtK3BAS9OfTOHP/NRu4BsgM80fkO98cuFJa1RIJAHCxUvi+Xj3g5/dFIp
qINw7DH+xwi0DnzbXZFLWwq4Woq55105v2ycIB5ChaPftSAtqbm/k2HjonknJyzt
SrzuLWi5TMl24DpXSnaqGHiuXb4ZLmGv7LzGJ8S3lqlOU7Dg376d4uabddxmBgY/
mdhiC683q9PSznbTMgjiSJsku/gkkGZM/UgkKLqETSxsCcRiZLwe4qROdWAVXUAD
7SGrlWDL6njS0AmX0b0cWpWHa+u6wkxVmSrMKDU8rgwzxn8adWXyUqSRoQIb93Sy
651gv/r/e5wf9HRmUSOmAf/r4VQJHdfo0SB6iVnJCbrr87sz+eeq4Om+1jxnHqNK
bkdAGlAXSh6yk7JAWA1kwV1dHae5RlMs+UpWmKhE3E5u2WV/3b7xPl9yFvQyTz1E
rbZSA6nlpsWnwUebtQ3+iYdKi9tSQ+RJBACk6kxm68du4pfM+95cDMnhLlSbZL7F
GlMYIiyhmZwi+I69l0dA7fjwjTF62bSYRImoKNhouZkO2ylxAb6MRD7wcclnwxj4
2KPuA1ojsvuTvAzIg3kyjdjDahYQFfad670zQT7yc5LSgVV39gQk9RDapxmSZe9Z
3dzADgEol8S5shE5sfRXNEi4+JVoS2GLXB1C7YsvmlLEudP92hscOPLPsw6x2nHz
XXIJPl22lhVuwsamY/Focx5qbBps7u/dgZrU/kHLrNCs0DKAD8Qqp0dxzWn+JFb/
k4rKTXtmml7dA9K5ckB8cIBYeX+zQFj7uwHI9b7F0JuMoEemrNMlomfeIxiJoZ5B
TJ1PTRH5SKkutfDr0AN5HDQBK73YU10BwTGtdVs2ubh7cyjaPJlUPb0hw6ggWAQh
O9Y/vX2F2z69L4JF6FEGEmcRObj5sixMX8Nwn3W9wNaOr4A28ZJi2E52s40Hal4B
WMIFCMqNkOaYPFyvGMOG/QFL1b1sC5O68jAqdS9SrFilP1UzGldUpYAHCCJ7KMI/
ZYiAS5BSBhEo41EMaOVyFRs2vO7OQQyeOlU6hrZgW5OmURD3LRIMEqr5O5zbuVDv
X5DD49ncMN5x93i7s+HFdonwhH/VJiJqJ6qSU5McY2DdSOyWCh1E62vgAIueTB4Z
85mIPEehaYCZw8GMsOQbCQJeXyEpoH21+qJWqa71zoMjFpNBgJyEjgLJS6Q7jiy1
6unxLLdzBSdFX2hCE9vn+IB9oPsS2qY9+tgAa/qa/9xtBNN1Ho+DqWFRiCFyCvWt
5w2IkVALYmIdi8oeowU5Gba3ZHaHDzMUT3O/Gg+8bz4MI+VfWvmYI+ZkQdZMoOCZ
lmay4OEWZ8T6FFwH1wBjWOq6zxabAavN7JfVKPTnLFnEL+q//SLYlHujwAzmFCy5
26eIvhtfsThnwEHWrRXrODXCmpB/5SRFe1O61mJ2GxHfeskVMtlfsFG6b08s1n42
I34I9fErfzRA3oEMVov97mruqoh+okSvuGJ3BIdGiWlxSFAQUETfwWgHaVp3a1PL
Z8fzYet7DhN0p0MOqz7KAHlAFLFrPvg8zFBeQCuetDoKpvZDycKiP7JjvL6ONnmJ
jNGxX7jWc2c9rt/44/1BUa1TET8twEn1AalP9RhJDKm8wRE1O9iDrwaRzXdPFHzX
eXx3Znha2BBuUmRD/eSsnn6GbdPLway3labgFuyn7J3+3b+4WmL3z/EePVY9fEY4
sj+0BpoSlZrOHK8W9aV0u+t4fa4sI9Ro1V0/E1zK9x59rgZdZ5NoFHpe6hy2DyXy
5JkRbYiVOBkw/rmM6PBsPcrA2ebA3U/OXQJKnUjEfj1QQpGfdoN5VlHDqbWeB1ha
qWSosUNyLG10JHI5vnuPGB9MzAEqPubIfbTITsgFerrmKadiyt/UcuRFfbfHV/H1
4Q4D1vUSRqv9xmt+XJHGIH5ZIOSQli0eXR/VBUY73RcUldTOlfLf+Dque51ZnZ8B
+KPA7rvJ/u/ajjv7DNNa41Z8LEqxhP8wMG2o+A1V+fVR0i9RnLgslL4repSvCikv
O0EYuMhATS9U+iEXtLTrfiZUUnOFR9XJWJ3uuMj2SBwNHgjd82B9pZURaC1PsJrb
EqmntEC7CqUrlhaooReVpEg3DOsq0sUEziFHaAsorNLuuxOKS1DtTqRp7aJpuVQA
BoNhkFDMzufwCgNmYqgckPUYdMuy+fMr4G5ZXEP64qd3A6q77C8+ASRQBJbEzP8k
5sj8hcCIk+KOv8fOluDWSSmSDCvW8h++dirMtsOEBc8AMsVBIyqsZ9ZSPfjOD2cE
t/hjoh1s/2X2kYvr/5/Q/EXCJdI7HPaO2Tarf4vkK9o1FHqcGsHgyiPH1UFw6Nm0
Oa+ygrtv5cHjpXHWjy96bWEro6N4tbUYrHhyPXTady8DWzfY88C7ju0hpWtfZ5lb
zQEpTnMtWXrj52Wt6Rz3KE8qASG9WC9vs+6VNCt/hvP8zgiIRG3vLaRkhpc539FP
fedPtdeTtQciRR+jPZm7NvS2/iRrWO4pqGyAnwW/7OqlsQMr1LI0dozkfMXvj7jj
tAfLUWsRre/3uszkjP1bzGC3FQi7zGz7LR805t+Co0mblIf4+rrr08wHZzE+L9xp
iBArWi1ppqKM6g73vxwjNZTU87xk1vbwlRdUy62BzoE1svP0WJ/6+YjMqzsQbp/V
KziNbbnaHAfjnbhhsYOe/Klu3XL9Nrz3PQV7+xiVzhEXbSi3NcxLXyzbSJQpxqpB
/P3ITvsOBn35gWPH81E9YjzkqGhcrFSldOxZ5nFfrn3/Y1SacqaBPERyTBzb/pFh
CvpM7xG0nNXR0UcMdU2vCe44Bdk+HbmGiqCB6w0H2QxDOJLx1rZua5L/294DU5v+
auZ/91gasB+X9GVKAUBZO/pApxPYozz6QU3je2pEXuWq14sFdR4AawGi+BNXoJdg
GEsMxpCkkCaUJUnPcCk1eULlLhmA77APTlpZIWAeaIe0k8S+179+vpuJQ8BEu+qk
ByQQ8rNQp9elbZ66sk8u6CNbjlF90nW/KeUzsNgbJ1BuqUhAnYOsVAbsFToUjIYQ
mb/ScCIlXP51TQBy975qmjvyvZQMNG6igegoVvkU0pT9nbGbZDJZnaDjLB1lhmeW
iQBojC3vP5Ds25KoE2GL36/kln049FkPQooQTdDwSzWuo8gMWQPvkbjpjmV1ByE9
84d4A+2ON66zu19pRtwQL7TAAglbSYr5ONK6ncUx4uXpCw1ZdHHDbnaUkMztAW+M
Evi1kpnKBPwu8F/NkK+uFaA3spvByMmSlrA1TNt7+KO8yng16DScNdLCr2tHacQA
Fg4zHVtc693VVwDQzxs/aEfZGlcihCQNcOAXo9umMQmlUIKYV+SLHwSSI/LK1NjI
A4kX1VFA9hRHjsqlyLUEDogXgrQeHW6btbPQcM6rrnCL3adg2cnmMli33WcYz/Wt
BwSyLPpkTpzZy3C8hFGkLruyoYoRakmm1e2UnYEjZb4WNHHvTP6R0hmZv4dWhO0t
OfrVqVMkPruXqZNL6VoWym2swFRiypRjpXMlmg1mO6h6indZ7W+MxPJcaG/E0p07
kd9z4iJj7ajEoaxeia9N5GYPgqQVSuvzzZ+4I47PK8q+kHeFuJs+qBMTBIW1cvEH
oyjqKts8AYAU5o4TH3AZuZ6vdHz2CsrFURWLez+WSt6oaGCTIUaI2JK96QLi1jGR
epjmuKNVXPRjs+pp6hZmm7b0B6Jvr1b6YGjsbJ3/DeyTZAysDMsGrhlaBegX/j7B
rX3o4zdD46qB3UwioCvjQyYKAZ+Nm6hvO8zEIZWxVExVUd/U/PQ4/XzcfWtsgHoU
7ComkZrhtb1QMvVFQPdSZXA6FFt+7C7ddtqZPJTigtF60lB0GLCnzQdbhOc3dL57
0lGQrmVainMc/vo/X6gi33zIjwY2QnZnM/2ptk31Ykq8IfuiQ0yeGeGOp3APo1jO
bsDbHgLqyYqhpMvltnAUbqdq2MKCPl7zTF+daVSs6M6RPRS1aDccDpRQnkJKBOgV
v+Sst9R2WiWbJyQgzdAu9a3jDEqbwSmfc0t4yJ70abAvO46S5z4Fke2XZXYVQuYT
ETqDAKwgUcMpDaNbeehY3D4NyMxKvKFcLKttxdqvTk1e8OZUs4Vsh0NFA4tsBMg+
nR8BTCLS6OrzF0wPYYUU/ixYC/0s+K2PjQwsCEQVK+k0zCk3Ciw1+SEq0VeiuREa
DPwNt6TqH6XgcPhjvhKzg/8lBJwH6ARX5uMGnCfHcJ/MJ4b0bD8SXn6pZ22MMAsA
TjPSj37TSOZFtxO6pngc2je9iDvM5jEHL/jif6XXcUvhWRKYksoCGqWWjAaix56o
t7560m/hVncg+heemL94Pqy95wA+V0zUJcar7a94n1RMtJ0NR3MTBmAFqvyKWvZR
n7kC7qHZe0wgWT5c3UCxUIAi1ehujrDY2KmkrYQIc9K6lirqI2Lc6jRCRfj/cV8y
Y2wnXum71FT1UbpvdZDLVoxBLhTG1j7IrxSR4sVxnSVqQefhBZ7QeBNqAfhsan1s
AFIk7r4gzXugluyYPUMamrbFy/fD+1EdmuXjcNKZEkO545UdWiYXaJ143oyfBeXU
wHr5b8Q9QKxIwLHkB77q3YTBRyCJxAMlCFyDqSbIFVHmskPCrp8m9W4cxxqnkdtg
robhol/baZKhjb2z4WJShFBMhizts9dwdomMSQfmOr4Xtsp5k6vSEYdKPQWiEIDo
He9OvnEaiZGtARpOtUaFrG/EoL4tBZgBul1IcIp7/SkWLBLilvTh4YhsWUGLoCdJ
unpPT25t5RVLCfIHW8xD8EV2nlHxaLFWQy5HtiRoMhIBOpRtWi3irNXIC8s2JPij
U40bxOAL7Hhg6e1rcLzIP5ek7jhrs9EfxekVta0FKlSbzrHRdUbrXR7n7/EQjLtB
/xhao6VaExmU5pSzCX+RdLqir667nHvNC7izvqIf44THgEshKyF6QcPMAuzktNVb
XbIdoJtxcvyaEtIgEAHdpCHEx5cIl3UQwTc8w7hRjZ4TL4oPOpFCxaJ+7hFFxZkk
BoxvKRsi+P57ahEGh67q588oifdrw++P1jnDDGJ6SpzQ/tRzG4wwb1R3ZSqn9ZS1
wfySi/cBZ/myIqGLTvFEkjbCMzvkJZ5n4N+fA03q1lzjuaE7Y/B9jIxhmkBWhw66
OQSYwp3CWcz1JiiLTjQZbelg4ZpF50RU56Yt9ONmxMbbdmdVIxg4MwevMLQ8ozW2
bXzsaXF/em4Z1V5tfiZTpleHnisrJusP3Y1pqrhIZ7tCfLCcA+6Zg9vDkOzaxBwF
QEhcoqBG73Xb8K8y/s0kyo3/J0YV51+2f9GZ/9r4avtE6j4p+lRXqAXyRxSZmCLe
BGNURg1rP17RWxC5fgekoqy1KKuxmkrSGDQ63XA2NP14L4i0r9RDpWQ1NaVujlXh
V37I2xA6t65TDFlTf+IBX4QsnzJW4RJ7NbKP5pXVOhWbD7lRlEAtSxwupVmRcBCs
G5/slIAr6BfcGPCGxudDq9dMpGGPdY25MH1yOTIpRPHbxLRNdKaH7gFsX+StQipc
cN2smc7pgUvsQ1eRnSxNGUo6/hWwoP+7QLBTZ/MeBcNMoY1y+s0SatvBczH5q6Ij
/KpeOZKjMHyWAF72zxbr0MnbWP8ry+tlK224BhDqhLE1oBWeg8Q4Q83yhEHlD6T8
ztDgBy+1SFhjvSsIfJ8fg1L+dAHlIT7QnKB6mD12TnOfyLIco+OmKUa5Y951jZh2
WfmWyfiP56H2ZLdKFmKJUUE3rLHzyPsL8K7bPbvp+N//g3muITHto/s99kTxcsP/
v6BUxEaUfhGMmm8776ip7KyueHAzR7r11t4/hR9CtaJBkOyc5CGCQmbELUrXCKE6
neVF0Ljxorn0+03I8mwNbfE1jr/Qp0ea+OjAFGk30b2kEwwc+mxXQoWQ/NxWO7bM
j9os+KAw3f4SC9RSg5eHY9gz0zYOxndAKtvOzuAsS4l3u+aW/m1vPJqKZek755Jj
sk4YgVzY7wDd4J0CLUTDW8gvL7dVMSYsFzq+GluRmVA43NHh2DspJAGzgMHOycoM
xoPOOm5mv9RVtdnqPttn9hMpn6DMgKufMji//GSTMpsJGMK1yc/7ZDgDNVmVNZG4
C9Sm5o3nJ0hGf9SJAvrKd9ydPQC+j6eVXPohenSiIG7aUKF3kXOriir4arJ0SYVF
vj9IPrAowws+GRjsta2CK+Fp0jE8UyX4MaIAchTSol2R0UWEuiE/UW9L3xYSdqJn
54YLGsfyBkTMPw94taohB/3FW9PFeG8DRixSKdngPGyjKiKhEMKMkOB7B09kMWZP
24tbzzVqYEAw7OuyYoT+zqgM0ZXd8XQDN76vrdGw2W8k0kTl2Cwf+sBHvV5Q4cBE
j+SEobzpuPfwynmLe75+34EPRulUqCaCLW5pRbQwrUZBP7HhosXAiIKNa3FJYAQq
m7k+19Bi4kPucoRuaEAZtdJXr8X0XytnDBY268P4A0hhz/Ik0fKAmC4gFB7q7v10
9oLErRVKBRYX1yHdoLY74jpOJ8ahFIxRyNW3E7XEqPntfUMtQQ7ki+w+HkPoJ/KR
3LQ6rd1htsB4IgAbIBOSb/MZjG6U6Nta8Mi3+v5JzonmslWktPIGqr9xVmeC0Ja8
vppQt/QsYSyZ+9IP8Os3RoXeaH1QMJdzsUIvudhXyYEi/2m+a8OgZ/kHR94SxH13
Jv8QiOuWQJC/I5BoTByDZDfa5+0kJTyB2G+JwV49xtXQwm1chl3b22604GhuPp7K
K6aFBS3FWYfS3C8DJTEdEfahdQWpyZzuL2epWhURniizIbtrn+KdMPlfTHB0VufV
3oet5bDQg0Nu9m7i/zHZq1qdQ6+uKy0AaTkqxLpIfICa3smveyAPyl/pBC9ZPK1t
zlNHw/U52/068BKaznVXT24Y52vAuiKYpLKQ3F3JfQVPeOugzlw/nU+e+MffWhoK
frsP2UJa086QCUhsnMkjDU1o29d9+SqEmFXn7iWAHXTPZZX07JnLzL4/2FaGMjCE
0BtGlF8UdPIwA45lrMOxbyBKUHkZwKW8ch5M1ZLZMspWS6kT+xg4N2raLi35AHMx
uLcvnR5gUdMJb4hhO8i7CW3rj75YATpSqn3eb2jrb+DS9giQkIe9zimXm/FAKxo1
FpwXDO6Lksh1Iu3Lm7sbyFb3XYQeewy7pfyw3G2XEesGAy0m8Y06D7UiFldwGSXZ
Bpwu2jbw//wYztPJP44pqd2f3CDxmU1MYzp1WgsCRCr5TDFzsiDTAZOA+lfPbRpK
Uwll3cZSLK2EC1XEvGUkBoOYoNa2fRnBpkOn7xL2QG5+uGi9zj/Fx+IKhSpQnbWa
tXkdg/tUvqJIdKiY2ojAvvBqHlzFYtrKEziTqBwkTy3YqFIfS24+kuveSuPd7AMU
JCYPTUC+461HM2UopNaOj8PVesE6iFUCxmQQFtrIltt6W3NIdOhnRSNcQg7/97CR
DOZVRE0eqSsgqSPUdis/JgCiBxrVlQrPpGJEvj48e6rfhs9WYC024AixMwR+qJ0s
/vzbBLqMqkfBUZLVeMHEgL8+Th1H+H38m0UGBFh3A7YCPC7t/RsHQM5hpD9WwBvt
SeoeyAu7j1m32rqEvE9xwaUEXgwFIKaSnb3L+ePPtMraDlplac08n/f7cHnhHHuU
qj+bBRQxFizUE/cHXtvPLOW3hufI8rWdwqMYq74hbpJw7LFmKmPBsQqGcr9mB/lt
T6QzY323TVc4jRaOGueLCaXoWBcJVgC9wEFxXHdKdfnVufg2MIUQCo1Iq6LHCJxJ
UaPTuSJUgu5Os5WsJEaz+vNdSu8TPfV7jczDePuqb0vZOQQ1r41mDvZSztX8ZEUC
oEBmOvDLym+GqfGh5l8H7LRLf0coaemgO5ctE3Xu5tiSvUCF4Jkit0of7rsWMXGe
td+cUSF9KecZXh1pHMsLZWyXIWHQfhYJoWH2Ti54lvSy5fON9TuNaYLk87DHt3rE
4wwVwWTlBKNa6QCWJKPTyawsQfyGas490zpqh9KCcGajZ93vm9x8PeU2xiDSyKcv
IbvUeaUtAoJrfqZ7VawZbA3GUcZMpcEe/ps62NIgggO2UzjEJ0FfrX42lxeoUyKk
udh4YgFL4RedHoQHF+WWRpHh0b/8W/fOzoklXcqQkfnCtwo3P/o0JIlbKEbgcLL+
HNdWtUsmT+2rnQSMrPP7R3MkGg0Y0OBWcKciBrgybYoWx8xXus/8LHjnkSySkcMK
V/NmGNBq7i+D6B6KkGMnRc+TDWl/u0tPusw4+0WQBvOLj/1LDqbgUnECzG/CeLIm
hXorUrusH6rsulorm0stKkA9sqacxRndm4Z40OvLVL7jlKUSdJZF4MXdcpWfZS14
SIg1WYlw7DhGhGX/nA2BMmrMB4oovbx5A7qQPvTFDcjONfYJtVRP6yTqtDCevMSe
dzGELbWuDYmVdZQTl67+iCmcG2TLev3+OUfKLNLDiXhLmt0+0oycPqQCW4gkF+Ld
TYAnyLGYSUUXpnziJZ5c270/ZJm0nR9haGHYeYVf4lh0FQ+3m+XA8jWQeo0AHPJz
nwXUA4gcJJ378IgdJH/ISNt2ivAod8SpDEfur0UX1tx4On7ZoBsLHIgxMzewwXOb
RE46OXOovNVtwCjoy0iJ8Mv3BR0GGnc1PTqcckovfl+YVlH8QS09oJf8onx9FDIS
xVYQSB23I+7bQSjLjK6ynogsR9JDRbdPUXxDzQV7kaPCOzk1UWVaoHLSU5WghQR8
RhHlJlscSVpYb3QrOcYHKmYsc15YYFQlqQuiSfVSAMCtD7W0PK5h0J98HKWIT+KA
653LiVYPJM0FTCVfLydFd5xPy10mpnqjkffSjxn3GOt/IpVY8djyLI2u+2Ifec0z
8WLtGRloTD2jVEno2E2kdG4e9PSKAJnegsKxGzEhV0kWZnhGyjFJViyN3xBlf4oA
stdWwt2oMycyBs4GZ0DPzcDvzVLCVM6a6g4abmJ4T1WBxOV54yxCKhjXnV0zAC5j
PSnb00rxCkpcdNp/+5DthcHauxmphIZsx1eByIubOlvSlG1xRUe5KxRhP4FL9p23
l/EDAM6iwLRLufMY1Ol2JvywTfOvAgmT0pKRIo8FBILyFRlofxEprmknbC3NRWr8
Z6EVZOqB/IJUV8CRBOD8CiufqcRRbYY1237aR7ng1Ea5lcuW3o747C2s8XvMW6KW
PxhRrFk1Fh7PsCclKbHSUDL4Z9NdFOSTDbSdeUnR+xIkgwzXtgf8I2lZ30p1mxHq
wDhWGTDSQCjpWIy3Eur4H0Niqa6x0UL/JpKbaBuND7bVEH+lFA7eyJsp+1KUT0Fj
6lEeEQ85c2LkBqfFh3G67MiiiQYVg0YKaz7I9TdmSYjZU+W61sKgy6ekpcasKOYd
ghC4hUwQFZFKj05d5rYeXxPRMPUnWgaC5C23XiH3r95Qt4y7ml+cv1K3PHKgKhMa
aixfJeL8+jcC1bmg8q25LLL/mZzGea2icNyyHxTsiPl21XtjO93cZN/vS8oXMRSX
CfowS/zlusA17AOKm581obJZkTH5qcjz7fSIFCjQHHTPWs1xYzLul3f81N8sifcG
4fRDuQ+Xhp8ffexKMRrGL8YYEt24P3lnO3e2248trbccoSKr4NdY/2+FrjxifufQ
y/+Kh0u7TltS2e1z9J2T5fHsHrLR35Ch/qBsEKtBzzuuGTF0OzB7XILDXBmiu9l7
tYnDtTu0MQ6J5BKtz4PWcVG7J0s/GuYIK2MBU6lrBlg0HoHfLEj58PRWf/dtQd39
dJl+fsT6dEVYz37AU6Yp8ieZ0CqkR8K0JSjMK2jZTaJxT89X3Dr3D+LZy5WjddXR
0dLeYOyxa4UdbEzIDWsPOc5rHZ0VeApTN+xe5iXJsEQmgQd6MJxub9cGYiAtLRHz
+xsQ0BWxa9bFOyiStFLa26rVogF/6Vqg0zxNrL/mIOCIZ9CBMt6JeAYFNjN+a0x+
YtA0QMqwHb/aktGmbPudxHHDKTzj2tQUJyK467ZI+WAMVlaUnMLafNd/afgguSz1
CzjqFSX7jJIwnT5+h8Z/F3szTQd+ZKwrhXySMViQaqp+E5VmDxA7oBms0OH54lki
i+o6mmlGJkeHNReJfO5aKe1ysVlH7iOLnA6ckOTvDHvbE/0ZwukU86jV/6lLIAvd
53KJi1qZmHxoTle7fOJ10NX1+19gE+sM2fQ4klzGMskAPk10b7oz1LZJCecvAr05
aX/qgPqk6vbaTFUXxZUppvttU1PjCosm6F/eVr8GMgFA1qNsPp6zTdgDSE5QYxJC
yOgg3sWxpaj4NZcd27HY+V8rEJExFzPY/OjkkJan8UFRVEO8YXMReviMQ/qjaUoc
eJel2KbsfIaLatkECfp9zTDk0NLtWOHMncun0GcoFDQfr3OFqN1qvmHTajpG/+Wu
dj+kyYvylwlx9y2TBjzMBCkttz51btIn6Q5780/vIX8+h/rbzT6trT0vh6O62gEe
GrsR1d/3W3XhG4x5sPWLr9bkYC/kQB9VwBSkpJJFCUZ2+n7vA/m+gYl/zRwJz4d4
TYYr/5eW0i2xRK8oY4DqGnvV4OeC/hVBRIAQ+ln+GknGARFM41EvWRpFoxcFi9Te
VjLyg8650qAFp4iqEPcBF3CB4bd5gLKTjTxYhTt9I2FBhKoenk6CPoDrRyjDulL8
6+arFU5KlLr6lp09Z+Iqg6e5hXYEA8ZhR7moEDZWif8YAFd60BJExu6E/NqNPZ3x
JlThZA4jmf1f0mpuetItRFObxL/g4SpmMCQgm7ci4/1LsJjxX0XwdDck+sifd895
MDJmHMkqYll0UNYWpGXHhIZqTLEmMHCIDEDxOCxwZ4hbjE3rhceeG4yi4w4mAYgH
sAB3Bm8cyCdWn5DfYEi1XJ3BMvsViSJzz+IgubKeX9FNeYUodnybVy6B0K0HCumr
VqeHK2UXBreBI0rFw/mrrNHLn/drgKRJULxT/QbQMlzfqT1LP8BGggxPotbdRxla
Wn8j/svZADFt5SyvTUX9AzbTRpmX6+PDJxuE84OpAEYpwsqizkM5PzqG51kqeTG2
JIFV0rOc/2YONU1e9QQFvY1iV1EcYP3j9rOYLwslgm8KbwRYSsJCnp5GtAkuMQ7a
ywhGmwr1RN0LINfyEfx7QL2sJPE5aZwqFKCZwdTrzoFH3CgoR/l9q77L4S9Z8/6v
8ka7Be1Ad5qWjF/KcGpsbiZmrEewy7NHSDdHyeT6chK+Kq0qO1i9ZuzgdNH+kNW1
vw3MRyR+iil7fx0Kxd/NZa+ud+e2TVLAUUa6znuJEOeO77V7ldFCONyADBA0X5CF
ouV5zKEwRvJ0icsGdpdRzSLLGEZ5fBVmg1sIfU9LuPtICh8uPMiWdB5TLj2g6/AB
FcMA1IF06ONMgvUtNhI7S/VIrNQnABhi9wNL4HA4B1/gFARThnYPm0GrfYp0xQt2
rMjRcT4NqNrhQ5Yv4A9oCpzWhE21kNzc5gP03dF1wJo8lNI1T3C+dz1zJ5FIkDFO
uUaJdffeFI/ILvlZk2S+IzXWesrEexOkQgxnjz2SN4kNQzWHHi4SLdtZuiOVsBlz
2zSuapOLbV1T9jcSN785jV3kFfcpTqrQfCE0mCBoAb0ibFrgkKkl18fv9GWSxMU4
U8PksQZHUiEsrzF43j25eSy9kui0j496vP0tj+o+6h28oKnI+kMo8qODDmkoRbVu
ssOee7VrwPCxoh53ccZPAIADdRTYYI9y8AhFZFqUvtEocEvpMCtLUWP5Pd3au7Yd
vondWPXsOHS8pdFvXLk8ZcPG5sjvA1DDClJZcOW6gxLPQQeV0LSu2SawiAKlQFgk
U8wlrITVd0glkQSZ/YdHA6u/AJjxoBKAnOiUp+VbLtg+I/atMTdumdbPV6PEu51Y
+ibSlyXYgWwWDl0oajsdUeJnBMT+Ea8SQFdWn0p1LvSuLgTb50LQtc550GKgr3Yj
AIMNFtrRr0h69jea+LKzxhYzwofEpfhWZuVcZi3p2lXp31TyrIZ7tYgXJXysvIgV
GqF7OUp9DMtjqtXBfOAU8C2KegxWSTkkHj2kbaDcKTUaK/L3dzkpBPuyYbbdw/S4
5tBWY+oUxyJh5Xff0v/8w+L55qdq3uTbeVXv2E2rAxU91+zR1KKxKZ5cj52Ledw9
0PjRogjR7B+DQnEJSjRMKEQkfWbsCd50ZfWwwn4mUMLJx+u4UyIjZbBD46fN8Lc7
75TbxYldo2qzAaWs2eiWl7T+VZuURVfw4bFWwuowA7jK2E3LVJpwoArDidP4amnZ
QvSNWe+Uh3M5I5/mPGqnuTeb1bvYrOATz4xOgzSc2dxYxikn42qoeoh2fnVB4KD3
kqD0qcHNpVnOno2BmKJX1MTetAuNE1KLm+UORT9Ro6AbcvGjLa6sh+iikY2SNYCU
vYNqfYw9bx84L5Fb22543TQYBlIgx7QMprgfXomVXGBSwsN5eEtreBwx5NhKSrV2
8UmfieaNAPbrnaDgJ4Tn1h0sAWukpkx6MFUDuuQkEKgWgbLQicyB1FJhbQ3Sb8ml
IJNmSoqteotZeo9juGVKB5krFZKmc5VFo1cVhZejl6vDnbPyLErQCyu4NIfscxMd
/AdojyHIbNYhhmvuqrRanm+L2uwvP55yPNYcPaONC15kN4jN7WQAe4+FLMS+l1+L
3OFHxlnp/A9EjpeYhwSl5npmExUDRmtQHqeZ7/l2K7avK18tQ3Rnh/eYk601/KPv
MFUzWTF8NSiPa24qTn/Z332xzeWahDTUz5den3x59iOyhZYtF8XsWJlZ4wPu3L97
mOQbg9ClN+RFgC5yjRBoyfhygZQoCt3UieesGf+Vc9d9kaVyLA+ja5a3hITRT3ae
a4aImRN5YSCuQhKPg3Ra0HTf0HHXNxylDMp7rWtuWaYiLgTUJ4cKhAaWGd6UlE9X
BB6qT/WllsS2BGzLdm9l18E1IgbA9LFyHJzXpLSjVBOuHr+iczKsqIudrbZ34hWc
ODTHXbBsKJEcsD7EitY4uLypfhaF1dN1hqcFHHE+nUbzGKs9+dTLoPeOO4JPv3NZ
TnrelEM6yxmbfGJZPbbcYIF6O/F6hLSCO43hOXW1KaagxK3LWor7pH/djJQc1Vkt
n9SXfPMFmDSl/V0TgfM5/qOv6mqcmSGvd4PgtEU+3FWkeH6ZLizTlKlRbdXh6Yhe
dFo9n/sV3N+kkQllo79F543wXPpKOGxz/G4jIcKZgBLIsng3lUPlg5hBiT8rG0uN
K3jCO+sbcSTNOei7xSceUQavjTMWJboN1qzgna5gxaIgbU8fxQQJKqs+Qoh0nLcs
qANN7D9rJEQQLRUKG9Ofoa7NbaUZCZBcLDyVKNUnZRN4y7qgs4+FO3c3ocIe8hLq
P9CW9eSQ9tMNhePsKXXml6R/Srcf6ejPd7GMsUXLXuTgOI/fsa9C5lLjRrXYsxbw
dXX/l2AAd4B5moldVXO9dyz2Plsr3rqlsbh2BEwPNdDggleX4qNS6YNe3AEDzwS0
XvCcW5uEzXqxia61p9vWDKLJqrfl2UutgQ4fteYembTNLmbpWAYO9s3YdxnRGel2
JzYGNbq81SSUmVedyWz+FTDHZ6dNlfAKxP3MiupEYJ1qb3xfB4N38xpfXPwowgwI
dX9ey9Z2IJpjFvnuLRPAz41W51koYfgj9Tc8rX7YyeuE0Cm1SHuaNu2+6NRNgqWA
HsaLfG2NQH4kmyFnqm6iwtdCZU/EzFePPnC2qfIMnbm/tCHLQmwMwI7k+ZK+tUZ7
CLFyWAlaR5ipQMwcmNHliyMAWEb1oczIzGFIYp+2t0th9DIcpf2QW+rAMmeFeY2r
yriCU9ptszsaZVZxoRoemg4QC+5+yXTg5o9KEo9Pn2AepSj6XZXe+p+XW8ArGKUz
CfxGXRbTsUorgJg4g8t6AHtLJUAHhZaCyc5e/fmZnR1HEGpYA+zN3lVmLXx5+Ncv
6aZNi+JRqWRfHKwhlPVDayiisMXvKO1IEUqFeBL2MvPJzfeW+QDNtAXgur7bOy3a
/CsM2mz1vWOVnwnZwOuEzIfvfPJOwUjK0dQ+dv2QXnbjSlIE51M2s2h5SsnxUu8v
89/TIfpyD6+W06+bLAS+N8g8YsjzdqG5SABV5LNftgFFeeO91++9azu/EI4a44i6
9nKcocEdbGwPKngbjNliNYO1gC5SBfZlkPG94qzPmSKAqzEz99k+J2bBPe5Xqike
wwf8o0Ka85zW0qHaej7dNtlZK0BcpSqrKxv7FDYsNy/0Q9N5Z6WSGG0UZ4/iHD61
ohNBZCLXRMvJk9HIiwDRV43lK3+C9FyAXoBE1CBTgF+aKh6zJVACTJH9C1Oyd4ik
XCRwQROikupUeJWrc6SM9ZvDTB5DZtVhabJ5KQv8kryFND2a3d1gyhDzlDIQft7d
NC0Xtp8dgtE5p2BoewLaI8BCWA6TV9yJ4dXxgQrKp93c27e9KC9s4yaZXuus24E1
IV64YyrgD22rH+V7wp/+mVDAs1LIG8zqzQY9rJvmPQnQgs/VyRMwQuU0FypQIq1E
6GaPg2COlq73xQuqIEfibKzQGwkufdHSdHImvpiIDcoV5YoY2XhUixx6NParrJb0
ewwrzSiOzeX80nOcHMdUQEoFxu+44Jmcz/497LIu5Q02DpnObZLn27XYwpvSxAIE
NSVUUy+vPq+v8DridbRniyHSONDhc0q9ymbDrMLoPV68zqTX6OoN0itdTMjyqKp3
6W5lye/5Zj0Mixzfg20XKki2/kne9nSYDd1OS5JxVJDWIHc5inTXYG8wvY88RkJR
LMChcQ9qaGd4ebL1mbjF712pD3wtiauTbbCp1+G6bbw8c+zxvsF3y3Dph2lKMG0f
iU6xx0S2dV6SitSNzsV7cENd/p3T6eNErUbaXoQONIE7+TOOn8zPB0g8d+vcV0Cc
KnalkovqsLL7KXBka7rDaVBXzpjVJ/EBjzHygEulIh82HEFkQtkZ3GYpxuC+uMye
ZXrDcg3DN8pt0gbzVkgYyWzi2ILbvWYOZF4q4WtXtp+4BNO2WOv0ueKfENtqn+zk
ih9VEARJ9E7BNIn0ORUg1SnxSwLEFUlSFay23/5Fx9MdMhhVDUAjrHPI9+H0p9yF
xut8nLwG2jAEWpuflzVRUXsnA/21rcpTWztgiP6NDqfftLAx2i9iQQ8BHGHiudz8
0SRcFACmaZYdSFj4+bg6C13v8EYKLbjKrHEM3+SB42YFz9dZpPYyoFM7SdCSybgQ
NcBgKv+Q7cI+qeadf+HFYXbWuNqjhVMIHyG6fvkJDso1CmgcQJifDRzOwiOs3Gzb
oSz596TTBv/nUq2D1yzyxZRPt6uMuPqPwKZANWFAEeWsJv86kviOTj0wMAnyH5al
2LWELj8vZDWxqFpkEGTE8QErpKVN/oiTKpbrKTdo27hJIFGhotPCIeb32paIGF6d
DciRmUFQHJp0qXfqGSsuo1Qfm08BI2LrhG4fQt8vFd8OxxjiTNEsEDb5vMfk7X3j
o+Ia45v88oi4D+UhNlHuH9g4SuH+60pIu9o2v5gDB+Cb+0V/a7aFFRdHC0A55bhG
9ZJwD2EyptKoFR7FnHDpyOLdFMjNYmWalRVQ+szJQ5okPJ5BE+wJHWGn6E2fjU7X
d5rn2N6mid8CmxS1OIBx3Dv/6knj2FfJXnuOTE1Yg04I2DyMKpzUIDVwMgcGB9u6
oER3EKmWgS73bNZDPME7dlVQCyVdDpsgrxdpyHNz5HQQO+qJKsmkcPkw/4V/AzTF
Ixdu6K7e8d/cqYJ57N170rLFKJE1+RuhC4sj6E1a01qoR1YXAxa02t0zSZrc9o+n
FatrmGt2ELpe3O0YG+k2DDHEtD5LV4tx10GgnM5/CtBIvWAlpagD1K696hDqwMIh
9P3xuVkFNIecLEfJfuBITCTDYuSrJ4MFEokVqnhZdmwB3vFbOSw0n74bVh6Bn9fL
UiinW3BlbW8LGB+/p7LIlVtsxvNentpcalldG+Nt8vhAFs9pdNHHpKXyszIJbf3M
Ap3wEeLUyyJtBpg2RFo2qh+f8t5ZAMVlGlDPozFqPx7u2RyzznH+vdrAYvXn/UtN
9gfx38aJwIlnzvyRfaHzSq+RKfKw6ExecQNuGVUEw7umFaprtJCklapB1GyLIG2R
rhPR5nvb/c/DVj9OIsypC/TPwZHsfyt6owUE35Vw1rny0E6fgc00soXGeoXuNyr4
`pragma protect end_protected
