// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nZB3mYLTW19QoMua3nqAoJB8vxtZ60h2xC6uKXjVO8UHvSQUluFNWPAJKk/8mSMN
LSJQveFquGa5NqMm6zo17WF5Zs4iNh2s62Dpq1bVeDNv3EgVLum4VKKwtOqSPWAf
lt0CBXQyYpirAIsPARx0NJZJ4VN/Ri7kGAdAS6o9lxk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16528)
kmt+ScgUnzl7w8pqPDD9h8M2+vOrBNJhJuf1DGcyREt2ssyxRL42pGK+nc7eK8nG
UMVABEjcPXwbgs/abmSDZPcf/HM8bMYiJF1BVuAREIirSFMxLeRKgQyQn+MoTF72
qBqHG5YtnhtICiohGGGZjNkZJLMLgggsMm6raCnhZypknspoO+1r9Jw/BrPP9+VH
cRvkF6Qf/zStfiBoQfY/KKmmCSzpF7/1pAgVigKraBaAlLWggB7O1AYBdmDQf5sh
gzo+V5/vFnoGPsyjF4dgHFueq0kKQzKYUpszPiVZiyode/CC40BSKR6l/cfN2lBU
rMYj6UHWHu0U3OuqEQfc971xtKXPXCO/fl3vqSGRYXY/uMvM0VfO9VvrougbKNPV
Ok+Wj1Oce4EpUApdz4a2J04RN9Tr56IjLIOoDVaW5lCY/c2wBnzPS95BcCFjZPJy
YhyALBFCMOnjJ3g59fFBdFqX18C1by186BR3CLaeFpoqtqYuyNxLsTYSoToxjbkY
UJw6qjBx/To9d7R/b9iM1ktf7I36r0etfPlgGAirW9kMSncr7uCxpgr3ZwtKxTLw
vD/2Le8iQhKhESd9RRNd53YZbe9jLWpzHYXw82f/t1EnTVvriSV2yBh/qs3esu+Q
ABxpC5z7Ggto2SbU3LEFQSZyaPIDzQjPPiMT/jq2biQAtwFqtwk8BjV2QBgFkERi
bsKBr+2XU9PcNYbss5kgmqkcyNQG/DghKpN/X4SEE++2hRXeHnD05pB2j5NWOXlX
IzgAaSMIZ/K/96hdL/u/5S3DFqQiuTMTF4XPuBfp+NeUyDzWaFrlO/nnX++cFSPl
8wyodMEd/c1SJtcgxiQzts9r7AQWb6DeBFEZJ/jrfbLVTT+aM446ftuQxFpKfDQm
PViZEXbo1ciHPPNf4PCmzeUYktab9FtjRGuwe6b9WoMWpcG0F7nE9zP7As8qGECv
4td53azgORFWkCnYjadk3wk4MfBIIh1VIk9mY32tZcH3Na3Q3pNZg2EOqVuknlg+
x4cR4+O7tlJJUvBFfw/k9lBD/jwo8f4ytPv1Vrt35yISqNNOELEXPSBZb2/+Wk9q
36HaYgDtLyXS9hBQvKCMu3JMaorr8Fxe2Hr7XuEzKm4s3zUPuglWgCHmWL7rZGIB
UoMnI3CF8jVvpCV3gFbZyvoHVPO/W2HQQnDp14QgdbsO6vZ4eMZnUAucoFlimVml
ja0qeXaUE+Gm5rZIlkG9uq+wgIlUm0ROLFP7eFjuT616e8RrOd5+nYwMiIMOr1Y1
WYNNZH2qVuzerOtuhZg3syLUnqtaf+7yLsFqRZ1AkaVAzLQ+aykUiFq0/guIy4kw
fZFBpSpZfhBlZlSP3lTahUD1pc6qLXPSU2GVoxDQEtExKaeif2AIRuNFHpwwWfEV
chvlJiW5VXX5b6nfaO8FfWBDa7QAOr5jGTjADSGUo33+/RF59rooULx42/qAcg6M
qNgQLiWygDgx/BL93d0J3dhszafETYPhoA9mKZBWBhJJ6p1y/jJMbSfLYbjMkt91
OweNflcDltYkJX4B/WUA1JCkjPgU3ipaq+eWrTAJMV+8NX9VvSanWoerIdf+T21N
JzW5Qx7wt+EfaiJ//6Ie08G+/m1DCOLDWjm6915OturfBEe+9COUYtg2+0KFqQ+i
3pddRFmVPgMoH2EP4utbO5ow27Am/NlO5KU6ld/KCxCmTPt3AFPq3/K6vKPjjMNx
HgFq1Hl2pa6Ch9gpMVwx4JNaTbM7wvDZm8wVzy17MpDuQ6YAb7IqlvWjhvBq5V+e
FyfPQ1pqdKytJYGds2/R63DaKbAsdbcYQ844EZdLEnvQrcSHfHGs5S9PaSg2iG9I
Py6rm6XOA0sfFildh4QZZj+cvvsGW4Sumrcx4bJWn5na1GM0ZRr3KXe+IWNCpaKc
xnGodsagNTcYgX9xySu0Vrn4hK/IoDsVN5X6gD2387MLNZ/hbbsdX9dDDQeT5KgQ
v85b4shB03QgQL6SyFp7Krc3r74kpopMdMBXqfgX1SfREhevS0N9kd9ePdRMB0jL
C/HTMCBtsLpzT6QMFkne91wKiFM+ZxdU2ouPO/d7nmko736GWMYzBx10MoucAX/F
05Ht9L30SUARvayk1c0dEVMWa3NAHfeoBBiIei90PrS0R5hBkWvlKL7++Y+tiNTk
1ikQRuROg/Fq//Dez0MS1q7Nw26OZ5Fzc4eg5oEvSGyqk1YVvkM99rrMNPaiL5GV
ubv3DwpUTWrVBX0yRDSrMfs47W9WFy+F5AFEwwY/3ZK8iDS7GuMcOK8SBnQiK0nj
mclSFwpFSsYc8uFmLlbkAZGJU8E2fuUAsh+yz0QUDrhUjOzpLFnkoW5dg87pDN8G
RztN8bcrkk183WJaPOuL1si2czVp23rO3I4+GSNOf3LIBl3IVK+cPzn0yavOKmFc
f8Oe2nwe/2Ym6GIfAVviffWEaYmpdXe5MYRaDlvjtfRWyCeK/pkoSSQGINNs3KWm
UKWsZkjgmv5WIsTbsqISr5i0gNes/HDCYUunhX+cZIk9WVNiPbCK1lbEBCFY65ct
yVqInwx41AwuH+cr0of5k7Gx5oceiDlk/lChKb5vXz/lMjO154S5soVqVl106HS8
n2+jkNY1oY46qiNRPzvLi+aenS5PHP1NG4/KLLARoHOmec+15STYhaMQrId9Cz+U
cLji83w7sUHGts3uUxb/12nDvTEAuvRFp9mUa9pl9dm/Hd+o6fuA2umxzp9pWQaG
9b48KCriNS9jAKDbL6VJUD2Xj8qyBj5Vo8rl23N6c2i9tuTvMo2HLbYpp4VKmmk7
YPDIiZMZRNcfEf8qcem0sEaLMz07KMj0D2KqfPU99l1RiK0U1UY8bQZ/fuRT+8jY
cQCvCwZKSlhIEKYPGZC+hHM01Yv7AcjcDoC2lUV27MKSruW0eDsESMQ+Aekf175h
NUMwWWfLsEfhW4FhlKrcDHeqp4kwLPtBoSaItGSgU7qb7IdEeYpCXocshtfYl7Jn
sMLKcxYaJHspSWqsUv2mcKdqJexpT3IAOLaWSka0XVkXB46dfjjj6oQvj7BLgv01
D11lMNnDL1JnXRniIdWx1bcyYetA3FI22faWA+Xf48CARZRY6E2z8nXFVKM7Qw50
Oo3S1kpVgzooPs+DHnqjYgwCOKtCTy5LwHXaS9bqhYTJ+AMWGFtOBO80IY5an17V
vULVXgAVo5jV2rNKCabLpq9pv9Hs6jZ2z21gcl36UfZtK1DxwlFkaLXhtYfQt5wt
v2vIItlv3AvKxnt44wYXqjo4nit4QW7o6ATzy2YvY+MBl6Psc8Q9539F/rHYCLGE
unLX1ajWBjwlNSP+kdhOgioUm7+c715dwQ1RsHWXWE4n5PEMh+5+PJLa1W8I6OXN
bs2jHdl2eaoT/PA5Dgu68Lh8og1yzcl+yCcUEqDaJOGAoGM7NQB2jgB2fattwplQ
gDHGs6ABATQiMU6efv0Fb4m5jn7DDgMbX6wUXD/VL5gtOPJGzceILwCj2uzvmKos
yRP2s2EqpBFykY3EwHqTRxH7BpCc56nPjxTGyJd0SX5XLf0Nz+ajc4X0GeV/sg13
kzfQYGCWVXP5vqCwYF/hbSdIL8vjCH2yYiymERwWzilfctLTuoMfbj5cRATzTsmA
Mw9xwKub45zXQRL0F/5AJLEMsx0k1XsWm9QZli/vqKSJEQT6eAWD/apKeGF7FaZv
eOdTc0AJs+BGlTljQViBKLYcLqvpQoxouhR23j/N8moANAtyATnPV/06L2LZl4YR
/6un79Jvh09YvfU8DhuFXoUcNKz9ubeES90ajEfQCYGsSAXLPGDdWDqctRLarDj9
J3amCqvyX5jxfOBgv5doTAYH5lwCJB8I+KQdlbjRrjo0nHMzwKXYQIwAeWA3Gqqx
iFV7VVbPCZI+sS2Dmda80wLBDnVMaiDXONe1eNGzC/gZZLaEDzdOXvHq+4vQKHoB
0wwrqENA6/VBN8+iN2FDyJejyWm8qVZ3kL8bN7sfWxPVPRxicB9a/mJjLwlpVwwJ
rrRX2wdn31DsdlvTpf4vuALmFIZTZTfUEmmn+nagZ/mhZaW3HZmT+/Wu8Bna7gB7
y+jZ3NkjZ1MisQXTBqNp2fGyflcW+qKqgLGUwqv074AJJdW3A5Pr6hH/ZkUUZK1l
oO0Uf9WKSerDHd5R4Rl2SEtGQos/oDfpi5d0COBAByvML8K7O49+I8vC2yJNM6to
w4x2PGaii07Ue3OxV/xlxU5NjJ/KM0lXvoIbSlfCjXKwV5nSGDtSU0ztYL6JB3uT
8OFAGKyNBs9wtRWY1QOLKHqATscx3FPIVG9+8Z5z0h2etuYWXEMIkizgiKFDlwk+
efPWqjx7Su5jYveEwPJZb59109nEtPKVwBIcc3WHMSV7oO5KvQHSbsdB2IqsgYeI
016TFgs6e4xZAxAkC9mfuRObu2PAQVaBJcAV/nnPinLvR1VZ3VOkDThssRrP86OK
JsOHpR9VTCP9SyAxqFmVOdra0n7CvFXTvBIiqtDn1G+77tASCokhbVPDuVVfoYUM
cBu4pw2llbT/0OE1s9VJbnYNu6duJofbHM/fkP8FiRBIC/DJlMwel+IIlCgGqFN/
LF2q+jITHdJxzxprpYZl//bAtPVORx1aPS14DhuE3ZlzOh04IuFWy/69hJDpjYrK
ug7G1AwMm7udYFtfXc+BlWTTCgaPJyzWHdhVozC44ZycjehiMAHar1a0wAByAzBG
7O8BAs1RLxm0vdbeJGK66J9RqOp/rhmjAdIw1YGBefdpPqCZZWG5T8FQVYJtXvgs
vX7TOjqm0SQJ85X+AE1na92vB4T/bBIHuJd4aHpd7U/KoFbygivce4ZIHLVQ80nj
liI/DUFgfr9YZT3ZUnmNi0Xq1OPgndbbQLQakv59o/hcwABT9zd/6oUx9/RDEZV0
yw6UFDdly+KIpm7obASu4DRx+xsLk4/TgwLx19SW6/1LzaLe5R7eDxJSAocTsbIY
q/3gAgFSf64ea/onHabux+1ZxUOEzIq0vElbTU9gEQ1CyVfZp1UpeWczYfNKH2Be
PPQTFsY6FD7iHhdgXubksXXTrWAF6S4TILO+RP5K2GwkGUXH2MJScmrxqt2koK/x
2OChqdTMT/OZpm6ra942nnWE75SjJkHncPLlm/GbpfeqIJ7L3QOvQhgU/1K8riJ4
49n1qP6zOHs9SmuxLbE/fhZWqdSnhpIZeqw06suWXyZ930gcyvxtwHPewh15YFcF
23hmsNlkXDr82gSkznH5iZKDXMsXjObEN/c+w09g8yS00bGnGtKaPLi/IFvTEUPV
vDDgEcyqSP9lI3yo7erEo9/Otis2gW2UZb0yn4Mxh6H3+2szR9SOMy6G9KPrcpg1
jmonQtUvTZlj2y2+w6SwdG2ond4ZfwARq12NWqpnQboAwXd1RnOHlU8r+GWOyGoH
YVQbvWEodH/vxmROjoZ5hnsB4CdWioHNi8U6auTliUnLaN9ZM0x/huxJPmqyCaC+
wQXe4a1/XV+m6WB2OeExPyVh78lR6TBjQV2Vlv18dmAZ5WOCkLL4xP79bj9W4HGY
RLmRJlRsZ2rUIEhmal8R3rOKXShNp2Jm8fvS09Ij/S2/F9u+dyrLv4BJ5XW2ytcT
Gs/kBUwodqyDlK62lev4n9O+VU8zA3ZrtRmfFCH+bHeQ+f/QVG8+179+wEa46Qme
e4BzHEMTU2Y+E977C08Mzcn6cpmByAn2BmrYv0ZXF/9OJT3nVIxttJc7aVpRDB93
0jYNohSxL4C0jI7T4pzHuHXgeYDsLWLPLGu4K0DOFlp4eK7Derl1JUx0LvWfBBRB
Vzwso2RFri5wygXxaOf6lbrQ4rIB3QwpN0we4/bTzH6+A16jSpVKCgkmVNKDYPZC
81g8uXzc20Sy1MZmtJBpJ416t+GU3Lz78pAjSxsDNht55bdM0JkP6lGZ+KQpT/Zu
hQTqUF4bQ8s//yejFKe4l1f4gvNScZlNmp9ZgNHZ25V2IdW5KfZuG3+V2hqdVezb
WbMfg1Qe7gPgRfUZYPjjCxY84k/WCNGp5mDQPxiCafM9mLECZzjpRwDiDB9wuIIW
YF5JQVn1/qUXG2uV9t4YWf3RVueHXaDBHdlWm5TCXquBUBon5aiA/Sme9/VCr6El
uTuOLuc505vrqpFT3+ehIbt+/yp90c8Tvg92hST2QTSRvgmirN53PNuu/LVKGPp9
yemJVzC3SmXnm7Jwsk0ZXI0wFhind84OyaPmqWRJr0mrt5ASdaKOQZhEAO1Ad8QD
V4e7Zh+KHrW04JI++k6kpc+J8d0GUc7WciyrqKt6bodwDtSxCUapPTTI8AvIxIHk
bc5drox14euUJK9hDY4UWcMUDDmU4W0zqrJKEmS9vI40/HgRRqKSKC7QW/vakYhM
Wov9pozhYFtOiEnUPPde2iq5XLOtpF4GrIxvurtf3Mp29BgHKL7ArC4e1iUMyjTl
Q3Yf7g3rDmVqzax3s/zAHkZ+ivMx21uZp0QbCXAZeokjEYlwR53BSBbj0pzzZedL
c946UWrfMUAiUw91ZmQAxiwuYRMCYibccd0xP8DVEaUqyY9trQqHHMGCSc0cKlgM
QVfC+bCTPg9qA5FgdBvdXVOQubP46ORkyxaM184Fgu3xAO3Ts1jTeOcYHSoKnLVP
b4AkqfIZ7CpiubOkB0oiMVyQo3ubT2pXLtKOt7wf7uLsicIPwXbiPqR/b0QLBcra
2ZflaepclczlNUARyQ03AyWrmz97Xxl/cB0AYV/vGkQQYuI3edEjTVj6InpbB+WX
XwT+F8JAqBYNHRQ2DfhoGJ0Fnnk6XDSaWuRUiEoCfS/IuwPnGPZss5vxq3cGlp8d
u9Iz87+3tMzX3g/p8Izgx/z7ce36c7hWEyQC0wRSBimaZDhvew8Jc5CBmMq1iVIO
qQfOHIn96v4x0lB78t1jo7dhdidXb9YiOCqsW/cRMbrufMNykzsPPfXiGR3A+Rsw
nPdW7DCdYiGYBoYxwt9yhiPsZ8nTeOLpRYAxtcqWHh3FUKT4yMp5blp/Vkk33BAc
fdlJpC9SUVQbF1TuHTVQTZBgeFfLllFuHC2WO3TppL6dKOiPagMOLB9acjsdN/P9
NE2KQTSn61HgLrZoeOpacHotT9NU0sH9zx4Y8m4zrK2aLGxF35KUOhZWncGfpkPo
/xoB2H5V1oL+xFYNYEhQCrbn2KFDNxgttXI4DsRad3+o7qiBb607kvEnfLVOtFUF
B5FYKMwvgvS4L1awwd5USwqIJMuW4gVlkSiuy/j3FmToni+CPSED7rRgrrFO3rNX
OvcMi10Bf+fVLDUEl6lfw00ZPS15/q7ktGHChongx4N0FP9T8Kyo/7kfnL3d6d+7
igVGgK0HlZrQAi/W6CY5TU/4sT54xoEZaKlapvWD0CMy1mj3C+p59tMEKgurqeLj
FxeynnzIVM2003BFklhEc6kfG2gHRx8d97mpqszziNrgMyzTcaj0sof871WoXnPW
/3LqlwjcmQokpxA3D/2b3yj61j0CrEycKj7pM1/9iCL+3mqmIMe3d7vsR3kDk6om
toAsAqipv92KVMhLkoFqewZExtSW5bel3bNkPBOZZbAGQnS4a78291l7qGOldQKZ
/wYca9G2zYOG4F5x4sx50z/vb82S3AYxdmWIO7WrKN1qNqBNwwdHdNp82zupiLji
S9wrXzS+60ufwPSSoWlf3qSrU0Jf7xhUAUtju/LsuhrSRMSVgbo8xWQd+uJ+8Xzq
sbH61PKquEJgzK/CPPv+484tqcPkIch7P6eDHrYg/Bonkq/kH7BvZTlfS1eY/OXh
GKKFvbaHOYP+wnwVQYd6pI6Jx3VMzyCpaQbj2gr3YRmgK1PkI+RftREuaJP/Vxo0
3nB/RioineMf+ofrgjhn8/6NcTjZyM1aGckmOhBwhyLRrbgzwpkneV4IWdIRHImT
/D/OEjZ16EVLvWBrYODMgZCRiGGHUp35/6mI5CGrYpKvLcrSYRiBttJfyn+Fs5Ud
t2EKIuAOQf0vj8rozu/nTVEZukUEkpaGc3egeGpZM5e+uIwn2nAj035WZQRB5Uae
dtb/HweulYEJmSWRgyybweEElgeX1RjTDHz7qpLNQ0U2QzrX8G+2AqzG6H9Xi0fn
hghGR/GkamZK2RyGQ6G8ETXPC8Sn9vlBhRq2f9vcpEnLDgJnkd/XRCvO9d4n12ku
OLqNJVAdFV4dYU62ijdWAqcA4U0dHwJB+su8R4raCY51H9aR6a0PBN9yFI9qww8c
uAcYGBbIfdLZ3y4sVAE1u6oKS3+yhIVCt3laDkgFiOCo80YwXCnzuWGd5naEOoAY
uevuOvlu7cML7486fxKq710fWOg97023BnQp4Vh3MrMtD9wWZvtndR4j5EWWswwE
d35qzmfIqyFaa4iEQFTE2ZVvKi7nKpxxfDt4lndb3PhXt+R8XCReQbjDZhAWQ/uD
kWDidOn9zIvL44dZUIN6ZtjWBXyW4QZZfWuojmOpP9vKBlGipr9dWA24ViUKf/h7
u01RtOjDGsl+BkFx9lI0bRKsobnMH7ozCyK4kqVtMu/AFDieBC8Qdq76+wjzZmR7
a41RmtqhJXTwsQ1FomeADPer/P9LHP6WsVvdFRpuQGBVpuys0bIDJVbcwCDxD4aH
SEzeVLPEFB4126EP5jzXpS7b8XuwIEVgzBZi0IEBaVpAW/23+A9EU4+v1KM5494E
UmF9dmvJtROt7Z+sdJXQEv77LmQQmYUGoofe3xSojLwCMK1cDd1f0L0I2mUj/n4w
rjXt4oOUVXzasBUBuRDjUbFdKdNCKSptVK56dObqms7sttk/j9Y/tsMRDiTrgIph
y/fRdFUzJViPN4/KexQAVbBkvjw5+vjwQtneCaHz5R5EIMoX9F9YnrruBA6x4NQG
JBfaxB0bqRjdPugsei3ZXhUbwV9m1cPNR3Hlzh8FuW5Y26XlULWBcGtUM/whJZ8b
C/ym/82WQnRFAdBeKKIjibsj2bTvdVJfv80hjLz/G4mg10Bgh9nBZEV8VIvrK2ly
ev8Tof2w9I+CLJ6PwmcB0BZsam3dwbc5kvA9bEQ16RAiGhT+ftX74e2Nu+7zorIU
FAUeEreClfgRewD87KBALsHNBmv9Pbj2eL2AjZrqoYw4w2+hYOaqwPOIqICrfocJ
TII7GIuYOhmYZGSfZSPwBUKX+jVht+0BsATcPPhjIMPL24FjnCdi979GZV7v621L
W6ct8Q4/wjipD3NzjDi27IMtUPg0iWjvikNxk77W4MhmdAHsP5cd9pKY1c4b8Ng3
SjbFJKm6AviRpo+VF5v3eMmzsMIzzBzd0VvOACbxhyiinuv72/+ssFR6lm7fq6PT
2Yo8itOHcCid+PSP5uALi9XgD8qZFyUaq+RiwShUNCtyX11yv4Pcb1lU06VWmyzg
5jM8ObmN8VUPSEMPEuc8I13RKDMAi+A6NrU2fMo07DXPmx8xjefiEGS06rZ8z1z7
ZoHStKWHvBSu0g/kKTJZ4a3RZwq9F/hwmkcxGOysLU0C+v8syZ3VoUHeVqT9K9YJ
2oxifiz7MJn2lUXLmW+UYZ6vVemMFJjE0+jK4rMbL0oSsYgyK8AXtios4JkEWigg
MCi/MS4ELHIj4HOg9f/HQKlOLXDFIp0OEAHswNzuLNjQ/fEWV87JcSY0l3DA2X28
gQQbrwTs0q0O5Ll9KTgHHmz6btOtTatIS12vw8WWNq2wF242TnHMkV4lPRztznrO
+10N8Hznm1/kQmKTjV4kHZZL5jTSJd1vKmLiZL+kpbgsGBRpD1qpR+Mw40OKWKPy
duAjzvSA+XFEXYSkOxlYdVes2vS7KkHtudv5JzhB/n1SZZd+KJBZ73p72c81o1U3
ufCjFvJ95kdsWkV4Rs4Qi5+JhuXRGMLMggo5kX84RQb0gfKQ+xe/c2o26zRjXXb9
8fWq5vX5IaW89LydT8x0GreNwxgXQeBKoySmH23di8wsYBLmoMMiG5v4rtccebGO
b3LOhvM3umXGmpf7wiZihTKDUVz9fInxs+Q9A+vyIUkfLIPWBJ13j/WYxdS9KQho
JGWgTxma1CW8e8nde4nrJFEysoA7Dm83KTlKuZm5BL0i7BjJW2i5iSSxUxZYzj0x
yAU5rkIRrAS3O8gpe8uIlY6FwEmvXiJhx+8lo7lRxLbnbeXQdumomXtuc07h/sBc
fxP0QBWR1uPsbmB0FFGOcJJh4gDSMyLO+ByMBFEiOsVBQ92+oTlWXANZZEzejYWY
DelV5L3s34bN4nChBqQs/TyMSY+S+iuIw74bI65lP3ftYGC96QNsYnLq1tjh8Hxb
2fN65Fy1q5gjYye0TEaFT2/qv7B6tK6CcSpDnsbTprN4BjItstHKlYNc5G06R81I
uq1sSzU4UmuLVgnmmoAx1wiJZNuEBjGt9BF+2meiIPML6ZFVYIeBHBSKh7gBmnWe
MZPjKR2VCS9ROoKDUxc6YaadT1tPym2REmCybTvm5KWkYXhV+pBzumkt6YD3gBHH
hXqG5Tka2lFFDfG5qST92dJ8fSvm5a9fipVXnvmDAw09gshLnuReE53NqPRpgfuZ
52KwcAY6Nqt0z52tkPg25OM2bNYTHobVvE91FCm++LVQD6rA6Zt4rcjS2lJwh0gP
bBWcUbbyKsfgAyNp+5giLTuTLwB+d3CfmmctJOeZJ/GOhSzQ0P2OUhjnCj1Rb62c
RhrFghAodxqQKPQ3lKcWEk4GrksbmFdF457zvuz9XIQmMfDX2LdAWt9uR7HjDHMF
w5f+mtN9e+5tFyK+Vpoz1fd1zLQlVizFC6SYcob3B55QkYCMa5+vnrbaBAt8CY9n
v9elFy5uzqRHbZFg487JvgvvyywLEhmYMPSAFWulVj4rh0PwoedwD01Pg72/38C8
3MmDHEXQ2oFwpiyMGDqKljaQRIuGCI9wd/eCQE8T9Pj+FwZhXRLoBsOU3hTZ74Xw
Ugjjnb5hXGtJxNHVPL+wjoEi19PLiObP5ZFRRwjywuEoqNNANY7PuU0EnfcAKOe6
EDX62gNqB+yY5zaWm17nlnfoJb6RDwxAKWvY7PdH60fZuS58FwOrKESLvcG6z9/T
V7hQHCTZudkubX1LXSrK0ZYFO0qInME6wuKGgE2ONqECehmNPPVk4wB+GSQmdxbL
bH0WXGSiaQ0urrvqqsQNN+xV5FjKTtenZUVGWHWDRr8OoIHPiWxfYlhOArK1hwJD
qEQ2A0rm214pS/uPTgctXYRb1esuug/Kmyht4YQn5+RmdOxf4hj2/6uGtKpij7cg
LWc0Y5y1SBTxxoauPU1YX0kfClIEkhbXZvgokzooIKmE41t407pZZMyFLkIG2lQJ
fxergZNNgaXZSEFT+ssHaxb5zWcRSlCkbK9SxkR8fnWtovDIjFnGNqrIcmekg1ch
3ZYVbXyJ5V6O6SxsySAUfHxLLA+x1XHBzmNTMnqvw/SJ1XFCrJI0j0lbyxflXTG2
d7xRE9lfIWxrM1zvsPO28EgXVFzXMaigcj/Dq3SBnJOL2LhuuC0aVQ48dkEnsf0U
uSr9K/rMblSe08Oro6xC5C9h1qE6BLRnYd6sDIc3OaO1wbne4Xg4nPb9l3MgedMC
Ukssd5WLZEAGZm9IrAmDHPqOgJjUl3oZOEeQ81CPpSoH5HnUUFKb2G3G4YZuP6Pi
S+9O7wS6nLjACC7RBEgQM6yU+9+eSIr1tFKBztqZoEG1skxzWi/AYLfVwR/+vGTM
xXDEJTLZcq16NMvGr897SdYnfpGiAc5epUwAtzjzFi1hLMx1dIdpymIGBdr8kclf
9lGg78K32k9p37EyQ9McPx0goEFS+4Nf0hYr1R9SZc48U/mX7yqcKK9a2cNORan8
QAbIFM2dJ5+10F5uszPf2Gzo+ZbvVEIAfD72nR/4LNb3GnhKVxh1i7ZMdng/x+1j
aMrCi5lSNpC1U8VFhMVinUg9e5STp+a0oarsZMLcbfTERN0xvdvEUyFzhZ1cNxkH
cTlARgdZ1fn2qV/ssMaepu/aIyPmEHflqKdySPFx/xMfWWsbfpVXLxteT8jIt+i2
wVKs5GVvYhOSeVz/DaKePNEekbLAZi/N78r0ODUjb77iqPM9nDOK3wcs3RjNZr5E
Eor1MlDwyOHDRfqiaoYT7uql3u4dIXxz9VIB2b67KOp4hPer8Rkc924sQG67JvGj
xwF713NeqzmtJiVKLFCFvQHMzOmLQQCIiCe2nkBGgHyd3y4Ncc+c8xtZuukfouOm
DXIvAka4WDI/YfPZaaHC8ro1NERLOS8YU0WItKSOt0CpqhPDqric25P0B0xlUXy3
8VRk0qJaAP96o9s1MGzRVuZmIqe/49X4HiIK5/2JKbYukuVdhlvGKkXtjn0Dj88D
Jh90vzFuM4mryCWjp9z1D64oV0aN+nmbpqTnr1PrFlg/msG4pEf6HSvp3fNOdCcq
UfjNoNdqyc/0WiH8nTDDT7KWBBHteAjYWwxdODBqPkVo0gPxRuSdBZrcVl/gNllo
BIyja4dVw09yvJ9Vemy7XubnLMo3BNd3xS3Wzr/6bgd998g3dQKj9wgnIYTLgZuN
bAFFcn/1/6aXoBnQjmSrJcBkW9CYnVoS7Evuo6/sydwxhtRrxu3c2vVvjkq4UnVi
HMSyzjwImNIC/l+d291298Fc1zVW9o1HD9If27Wfyd8VhrGjWYodFQpguzalosCQ
4mqM/toesD/cz6w8RYZl4s6tJsdBMplQaBoW+oiXPe0dPkTxHhyJ+w08s0bULEZS
e1G7xqUCEp648qe3hhdckGa0ca/80nIt/oDOMiRnoRjPvPP03qS+jlbOMpAwjWNm
T0L1skQ43N95mCseo2Nw0Bw/w/xRIkWCdnhKRL7Ho06SWBXMnnxd8wFG+2+nfXWX
8ccrtOsmmpRRFTEwMY4Guk4jQjn23FZ3Ll7A1oXxpLh4DQcfMXblFbRQnUpEV/wi
U0Pe0Zp55lLYfz2D3se4/RuYmYoqn0EmnMOo3KrsriJUwlCoOAsgJXE0tsp8UJrn
1G8kieTlPtKqz5z1LKiD2LwNd085+INLDBtIs2fcy14e62LczA8hmMGemt95tXZX
vHkiORCowNCKxeRUrDoagRpb/fKupd2UZfudPH4YKYC2wtIKhF6iwd57vLeoQ8l5
2wuq8NHF6SW2vwgJLbinxjxJw+NYnycONxmZHsrY6s5M+KuHqHTJrzisjd4KywUE
paQMK7UNQtRqm+ij8PpHj6PwlS/6OXMDF+JqaOsDF5/x0G/g5bKwhfKEOtKA0A+q
lFYUnnHhDJ2sp9yO6i5+HQ/kczFeqv5AilNV4ska1KgGScb1NHKh7vIoUWuCC/X+
66v7Mq6xdqjg95cTa2gGmcVD/VRKjOYZLO9lhjl4qH+bTvQJ3NCeAsLiQvoXHAnj
dbhp6Nqlpli9lVkZKL3Yc6uDZSVu6W3URbWR+Sx44VOSPT0hQDQeGVrrNo+hctbM
GKG6B+ICHQT4bND2hFMXv07uDXN2C8WXcZL446Exe0jvQZuK47XiT7c+Fgr5wJAt
iKEbiyV85+QFKdqR/5NKifZtXs5g1ayDDs4KbauVo6hu4A38nKd59VMb5u5Gpz7H
6vELsNleKTN4VZo+1VzPJkE83VOoXlP7w9mPfRB011H2JmoNpGVZfqGs+b30I8hf
3axi9ZkXRtKyBfVif9zh0ZTQpdqwpFH9l+ZFnW1fo3f7sAE0k26PfPxktJgCyPsV
VsuLrA7FDSXbdCcM58T4qGnLf20RoubDZhq6Pz5ASyCCFTGc0sqVb0KSVBXC00Vd
DO4MnMunRMjjSI31jLbP1q6+FLGYsIbdsOB/0XZZvd4cPb7QqpKnYOqK66ca7Rbq
BmSkWFrcAdpaMgd2GszxWai4p43/ZUhdjtjspq+0CJ/Jb+gW5tGLXFoaNV+BUi+t
/mIOOy03l/OLfT+yXbT4XjDLISxInBrY4TverijfBVdNwG2p1x/9SzGhA6CWodkg
fgcuWipg0YgUwwAZSm4jEh6Ua/9Ov5/nzRd+TnvvaXWdCO6oZ7EtcWn4av8hD6Kq
qvi+hPJw0ozFgFfgGCIJgPQC/bwz3/aPAtzfpxT4Agcs1EC9N2TKK2ku123maSna
jknOG3m3Dv/Jc9lIG6p+7dlWRY6osxkKzWHIrAvGRtRvmPV4XQdYT+CJd/dpgXfG
dioAXgNRbG3t+/zgp2qwFa2vt1iqFZNjk7vNwJYZlNmfRTYq0jVqSyU1o0eerLcA
W/jff0Xmu0fMCG5SyZxwCKF3NIaalsyrURtTL46qi4yypuLMd2WqRqg37BOWWyZ+
6ER+T2cwDECH9+hQFy79xQ9F3xTqdWBwo59VP9s7Ql4Vy+ouTJeO7XmhkozLqZQr
sA5Ho7pDA3eYi1LaK8b6Kj7JbkMTokpNfmVqBGfY3gVWch6AlksVpWwA+Z/BAsmg
3QdaFQUf4jX4Wz4BphDAxopLBUELU1ccgplX8KdlC5GACY6CHXpBUQI8rm6XeaWp
B3vBiCVoMtyxAq0Rs+qHGJeAIsoSVm0PbjWieP44qC8mlMf8ZFdgb14KrjDpw+PM
mbGzCnaDofhN4B+nxdt9lEVpqIIu+9Wof9unGGRxaIZxeZU/Sqe9QMYWtpwyqdOj
szO2WW2WvWh8YFnJAptJgmS0M37iI73NYCaYO1gmV95PIan62DBzOvFFqsXONR7I
k1RfO4qZ58jQ/LqI/Pr1VzgY5OVrq0o7ARYuKuD5VRjPZz/LQkpIFxGdKys0ou7y
dB8Y0+yQ9bKATbT5WAeAvUqzpTZdsjaysPPkfTD8U1QySpyzJGAs3v0ylg4arn4x
JA7CupsMrVU4OVHd0LVCTeoadJxNN6QcXktmYHcUMix3C9IhrRck3JgMAa2hQ0Ct
s61OvVYhZJ9zl8T3re2a2b8Df9krD8B10qHUMS4X15DFDzN2DyqZqF4HW+IXsAlS
EiKA4kki5/FAbbbrjvHB+G9egiv6z0QY3USA97Dcf03bz1Wv/Ht7Z7v9kvje9LZz
IHIOnnNvXlO1hRjUbJkM7enc+irO4l3vef39tjTxnII3FWnp1QVmxbP/0tGomQjb
0yWvwJGQm4biIB9/LkTeBbhhsArGqzhlcE/NH8pqDcH/hqApZ6qm+3wAMFymuvih
qqYIaI7pTXspO2rpNRnrwXLl8g2R30zH42FRDkqjn0F0xGf2Da11/Zg0GQpDMH0m
BLZpvpPLC6v1B+NeZ8/aQ3WSK+bzfj/xsgUsGcwfze33WEJXUGc4vvMNV7/dxEAq
zryvPMGXClH9mB5L9eH+M4cKRlxLSzxOPR9wuymA29Q6nO85yg++8Nm4RTqpb66u
HW7w7DtAQFbMmvN6jLw5EYp0GQYo79ZDLIHx27kqulCBI/Nev5rSiKz0HDZGWjai
XirfsPMg0Cw5G2TUXZRqGd6V3N3oRxlRPQpQBxHbylXcHzaG8t37tLFu4o0VBk2P
QVpLW8DqZ6IpM1DJXmHYeikLMoF0Y+wi4eI9F6ettw78LHnzrQdMqs4Lt/bJHApS
+4wgaVcrg54XI1+9cPA0CgyKJnV5dQpxJZI2l+xIgPPe77Y3UHuo6yZSxF+kxah8
zDTMHJfF3euBnzMQZsmtveOXdy3WnrXtW0rBKf9nduDycHsgP6QPdhMRozCLx8DN
BFhqMZ8SqERtS478VyqHq6qOEn/ZrNqV4WKUUT/tkUiJjUc6KlvDzVVH1l6HlANZ
4Kt2icZ+akHWP2iZRw2RQpMXOD2zTrzX+0J9aQnCxiF4+4vcPZtBLfRG/NLvBXl2
J4hVS9xC3DNJbjNAS6ZCbnumMFIhYc5eYpczIEjb6iBwUKZkTF+a4hz2Y7HjEqWE
5h/Rm9uf54oe0xCdfKGFogvUl+7K6kC++ZBeKvwXJ3z0Amk0UQegucxEi2LbsgfH
wXHYaobGsAOM0D0s9dttSAh8RJcCV1wNytn1loA65/uD/0yp2X+q0VDEE0o1007g
Kz50j3h17ZPeMpBjAO2iu3fMN74lfgM9SFO7oIHGujKtoGKlcPWZFgUkgyQdmPVM
lxR0jYtMSJtUQiygv1Xl5kCbcu2SrQS8ZEQpCDAjn64T+Q/DRv5Cno9iWZOUzL8H
sPZoJ7l9SpNsB5L6TWLdhzlhPTgDK8Kh1yOGvqpwUMy3pN8hZXU+pVpNNgtZXZSr
lUlRdJjdpM+cq74NW7yJUcYyMXFmySc4ujObghrA+tI5OyZfrC6MH9Geq3Pgi84Z
tKu/jvJMyWN4KFXQbZUpQB91I4uaUrP5bGMG6WzLJ4+DXFcgVhW7S4i0R0PCYiTv
8JvBuZMhzPsYmsJGDQyo06yM6glGnzp+C+0f1QKtaIWq+O4Gpxm3vgal/LS0HqRj
c3Zu4Do9iifa3uCp+rkPn07J0Wm661rw6cBxvBclN3oeK96U6Nr0VglT1Vs1f9ph
2KMffhUnlupAWcHHsdoX6ee8l81EdRhNRtBwamw+0gJ4iu9TTIbsmWZXQB7wHuoI
fLXoqHl1o1al/SuzPqW1q9yLa0ciCcpwE+0mjp7dbfg4oyw0fpTAq7RsXsUeTHTL
qAVcgiLo8vCseSDjRxcAlL0imQMrhveKaMuKwqTb+w+a9iiH8pns+BhBDmuRhVfF
5u4YQ+y5rg5HCC8KaUpHPy02j5qAIdWTeV7KoP4+YWetraALCsQR4bRfQDx/3Sip
EoZehWw7aOmjaNQxoJDNZHZXEeh+21Unr5qy9Ry0IsQuFWj1Ylic8gDOLeKxn9a2
NZnIPHiXwCWIA7D+i3L7sZNjUHWkKw2S/2JdKVRGVl+/uwpqf0rT2n/UHg+ixRUn
bO0/OVSyDohwyvJIjkg9I3FveLz/2iSdFFBIvGHXAZHebThp2HvXmRej+3iE+Bty
xx8YLY+5PoLAsW6vONq1pchSR5boNNXr9uxEFYvBJq8wRT4GYWcqyYXUgrSSZL6+
g9sHpOVUP8JJdIG5q01buF/uoNazpTBB+UHKd4mL3UFU27sLtKzdHA1XcCHCp+f8
AV8NM12AfO0G66Gug8sMHPy13tn665tBHQaOZ1ZXz8FcMyDZ2WM7U5BZCGyFaJzJ
Tq0ppXj6F70iQtlPTjOqbECDwUuUoWJnxRuljLIJbKTIb7jYeOgHELVLFxCZbiv2
w3GFVD3Wwlel44aOJyUWb4JEusisL1l/yPksQdijl/g1tAGfR5/ew2/iAwZYIaJZ
OxultA7h+WoFDFwZDzI0UH2HslOZBxV+c4UABIDAX4tCLJYXuYec7kx35lFk4jUR
NUCeisAqLO3wHBXML7LFcq57IaR9LW6eqEtxuFTE2VFMtHX+6MKZo0Y+ZT3iyOE7
DtTol0BkoaKCocCuoH26zVlyTL3yCPtFujdzh4/kEaTDpC7fxJJRpwwug22J7d7Y
dBoILLxBLvnQgf3J0T2ClfHcMx5cFHJpH7zvOWaseEb0u/rALkVWqKvSd23/3oXw
Pod21U7jhA0iS9xGJH7DmlqWj3XzkSAT2HObhWsdPXBW+lTMTvUxiJWFRL23gp/n
sHjMU66z1syZrS8q9uHoQ6OqUFSzZ3/paE6VNmlRVlIzv/N/v1w7EDEvWywUstxs
03RA01Z94iXaggWtaGVSTev35/1kg9EqkXqnebuNOZoDiF26MOoImL7hlxe2sstO
3m3KuGOPhNX5LjEeG/Ua/25BiHjofq/xQjLSj8irreIsb/0cwyJFD0pSJeDNokCi
l24L3SwMiakvcsEhNvjeeQdeoaz3+5vr5iQlOlOOHMtBl5fDAYziyzjSpSDgG9aD
cSGIm594K0cVu0VkV5xhTvHoj3kZvAmtkD0JkUliOYLr+QMrp8ehGE3wC3ovR5YS
9EzhVU2zrmreyNTQoedGt/OdzqoIt9baTfSNt1pxclK6oa2SujxVQCjUnLT3yPXq
bug8R2oEwugeDtIf3+Ru6SIyfNHDDo7/wmQP4dgTJn91K8TY558ExRa060QzuCQJ
L3SG6Ft8VjQxwEIciqLomSmIqOzBj2HSFXXVd2MUL7J4+qLIUhUHK2vXkJvdQopi
iy44sr1UcIhWORyU/nvzNfOFr3koQSNAfuEOuoIg4GmE6hLlxdk6qLnzpFhaq5i5
Ir723IPknQn+8TciYfNGhBq8dh0YroNYapMpKOSOGouAVxZuurtynkodJbVW9pfa
ojBxwNlc+EIyYuZonc8Ddo3SVXUb8Qs9TFJDG0eDf0ifZS10PtbY699n8COBsqsF
1KRIeuxoVOK4phzEEEyKR5l1IwxTSANzM9lInGwNb2H+ywRonNW9QGEXwgtpB023
6f50o+A3bJNi4W6ge388Tc1MXAvFwhN8YjtIU14+N8fUIWEu80/VBXHtTJyPz7G3
giKLWVY88zE3MZ5ygM4Shzp9peJYxRjKzaNkgl8YPFPWxTW97gUWIXMB4kBB+OeK
HXEcnNk58Sktk6W9xrI9UZfIeN7DHQukSRUJNd8oxFp5M6PXn8UOwavL17KRArxg
V3+9B8qCAMcOrL7kxy/d5HvrU2Lh2DIlndhrDOrOP3gB5zRAZ28nEH6ixgVaFApX
74A31Me02cN6r5qXoFd+dIKr6iSE2udAwn5UiWpHTvCLxG3P0O3WLZHfbIw5BN2J
U25cWPsklttZW70UtBUIutLWPrngOeFrimw6sWg8RtF2mwFCo+DmBoqkQHrfWMxa
YSn4m/U4dMYn/XvWOJjYVHwOZwGvfSGVRiSR9RExtbRUJHX3aLEh3uTNm+3+JNPY
X6VjpXvEP3ZOaxfq+S2ik+CGCm7UZMJ+bpEdxfoHyQEyzH+eqTKWqkmqkZIlzzJz
O7pikWfaTrStcf7J4HsS7G39hx4RBkMqZyY09RqypJuKaUPuRTpZcoXOd0Xf1Vlc
h/dNwtOCWWgLJRbt20a3eiV4H4w4lWQXmo5nMCKiMIZCmt1Ce+Hg/w3Sc/H5blFC
z5YJmZKjbeO1UYd5TJSP+Xlbkb5gMwZqXszkUmjo3QKMI8OuZnz9KfxrUyuq4qMQ
c6Yu+4/QvOA0IffMJ6Tek886mnmJV2VXP79fItdCm4I6/E1Cu5wrV8PzzIrMEtiy
7q9XY/63eH/5r9Ua2hJuYUW9vdRvuz+wEa3xtZhVp159hddIkg2y+Hzwei2ajViZ
csBg0kTZaGJs8n3HY5T+P+bbSKTUP97ZGo9iqB9r36J08g4r+0Dh1789DXgMNgeC
alMWhZQywZZlfHv8CfmHhGmk58V/TGg+Y8quj7Er95BxlIHjPZrcucnQZ3byK0vM
Hg8Brxzp+fm71tJ/8Z8BT73hXpmPpKB8aG64rODasW3WIbXXnb266ysylTLIVdas
kbqH4xbFAnDdNFKLssKl/L1OViY3vSJmWYBO8lMk+pX6CXuboE8V+Cton4tCq9qL
RHyzW3elSnw9PXZNG6J9OkU6YrWZjp1s5MFMNfvVC1Pz5lYdpKZWGdXq2itOZD6Y
mpwivLl+sWAP9tBZ/b/S3Z9AcSyl/JsiCieV8s37lu7uaW9Kgrsj9ZvOOPJ9kRsI
1VYQuPpvGuO5x6tHyBEZNontMTjlqNZSoQBGbW06umr/HO7HVg2YlYlUe1yrB1q/
/wTL46unZInALgbd5XTpOGnKai0gtDBlrUGETWg2HltltU3uexy5Ou3NWvmqk3km
qO83S08nneolSlt38qFFQ6YzTfjwWg2Ymo0ZVAYPUEhrmebfCQFzVHonuuY4MTEd
vx1xgaslSVyIBC9kgbhzZV30TTb+BTHFtaUI0u/QFrlpvm2ZfxvGqn4oPTXpzMBS
IXYkst26Oeh/kJmtbU1cZWPhhD+WuC2cPJxusPRhRGe7mnzd3/UXymmmGNgKS6jZ
zBBIUHwV6oy4ttHuKVjjXvS1UFIJzz31haDy4s53zTXNH8MaAyGZQZ86ajyGWd5x
orf9cV7g8Rcs72nTdE+YzLex9DLPJIJwnXsl7p1cgglKz/gTzubXJy7A48N9gYGX
a6aSAPvSGngGI639W7JYJ5Vfa/MaUG2D5j3CefUuuLUyEekD71CqLDTa3AkyX8pB
fq21gdSYAlSw2Qd089PBNNacz014NbRPUkjv5aRgDrJmbpI46b7esBw/zJUDXL20
pup+PLAZgI37NooLeTcHWUnfjOutNhSU+js2AaLEBQIS6me4MEibA6sdDq5KW6KE
S3R/jpQhFbHm3RMltHYFJ+/EUxEQIwUUb9zmzl6hdSgsWgB+hYCI9r7pHLCgt/2Z
YCCKGIHUqWhBSrpFwif4PrkxwRPTPIjaXv5x3A85ZGCnH6agYH83oAynxVEm1iK7
dNvQy7Pi/Yugm0xhRhTNy1eXxXTx+5NLAank1fKhFshNLMr/C+kvLH2shtScg7Ay
kVDS6l3vQ581xMWBMDr7PMMaUq59cnqrjVtbs8w7CxhouLEQCFTAQXU8i+wazpOY
FXxKj2eEoziIl/I49SzgJRabHIBYnkvqb23Z+l6dkfnEhX0pD/J4R5VaBIcqloDU
1E2Hq4Y3eKL2c5Dksc9ArlBj05ycjEkzVBiEVEdWE/32FEoxe9oGYpo5mapH+Qol
raGfJSOnzoV3KWvvXAcuZreLvFtolUl7i5MU3v8pGM9tj1fRqDZ0brUr+CsUGpt/
1IEdzqXJEN+JiteF0xJe7yPUWeTt61MKSh31I5z4WkHs7+JZmGWorrpmp3Y2TWNh
dYEcrQnFsuVO6XvSKqHg3GKFpdobVmEg71zcDbGUhZHXs8n3vicM1LL46y0FeAOt
dWDxH7TM4X1uKAba6s9JqxGoM/zkJU+JHLp46I0d0KNUUovmGg4p0B3NvfYMwwBU
O+Yb/QZS7pLPPXHRSd0tXmr2gdt9Odu1bgiw/mMFJIl8Nng7GwjYrvnl5y3fCShm
tLBCnFB0K6Yp0hr+UNapZ3rSwTwAUneApuM9ebnNNFhh6Korehbq+H3xL/sDsdtg
MtkzTQKqgi3ZYR92SEh+/P/K7epQ5sYc0PZRBbRmfvgk8yY/vPy8pSQ4Q2V8WzaP
1Wkoluc05ICVxFqqgNb3IChXbytZW9a/wjTousfh0Ersvb8dd3eHIyXzNdMlQTfF
C3X0uRKFInyW1bHmPKVe+A5QgPyA8NY/LYBbmmGK5LEIeQ9kFYRDh162DjrLGwgO
WiD9OvjYeIHu9TTS20q+DWS6jRzjvyEElJhCMEQK/AE2CvUSIHZBwQhADdZw6gHI
nT/YfMnB0kdO3dNamEo7iTVorDhU6wD5UU1e/yVJJHuHd8FUkP2cVHHh+y0izaDB
gdDcspFthXHrQSO/2xCx2QXxSmniQXOhJc9noTU8LwZkNZgmSl+8TjIwLFxRNPj4
weiQRpItmDH83dQzd8zNiy7IiPd/BW6NZbyso3asBaE1PmPV4/ftVw886KtMZ1jH
trQJdER4S/tRuq6f4QP3PubZNLT3d8LT9YWdXuE5tqoNh9P3pdqpD16PVhIb5t33
rnNQQbvQ2T5PGN3BlwvDKvOw+xJs6HqAkQaecQ8NyrjC7SHqX7pJKXAL9fNwkaKg
OGWzDhbx/jeRAIlWISBu3pr6k/HXc046HoTxnNnSWPZFsvo9FkGn8jT+aihYrTU7
HqFNduLOZk5MRCxnIYbzz6yTAm5LprRRaYyejmCDckG6fEnBaaipsGyyydcp5uIl
9q8iMyT2nAHZzT7PLq+c/rTDyi9If66R2Ddy8coC4J8iFXeY/cCglnv6toLMjfs0
hTP14MDWBrUlQ52OeuzvoSnN/VHygj+OXubUe3+711QTJmsTJddWch8FmOQFMGht
5fnviXSVvqyAlBSXgXr6DHoYZbuBYglKILraQPlMPlR7VxmMJ5L8aXUGlbi1Jb/Q
p52rRqnFoxpzKJfYNrSzHaN3NPkWTxiTLVJPvacD+s8b0YML1u3uyq3ptdfFMCGK
iOFfgxSAAh/hoqhsuz4ktg3yL5HkYo3TrSd6BnogdLVoVMw623Ms6g4A3nhl1/21
15nsIFCBB/+b1rUlDDF+W/5pjqT8ZGVSDmklJYTkFwoNuF57eJlsiRplhviJ11aD
bjIbfhX81KPvxS/mGpJTg5Z+myB7hFhkPXSk7rzNQXZRT4cMrP4e/NFumAj+/5Xt
DampVe0X7BlUYVKiS3odQQ==
`pragma protect end_protected
