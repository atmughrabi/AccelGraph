// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:30 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QU2I0Jhn3jr7qBwQzVJXaWXdA/0JnLiGe7YFyclroTiEKcmKlUCrwlkRRZLTWojc
NSq8jdzE0Diwr31CVYXh7NyC7wgpRPaqGQCaA9t5isf0x8xruI0KkEzUrJ+KDF+L
4Ikhsidkx3tzqPBndkixdSbqy2QjQ3uS08BGD/jCaHE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 45088)
W27vWSt8k9+i/soKm0ovo6cyyLrIlsk4UCiiSDEl+3enUhpB6SAPepIk5Uyfi/42
0kh5br4hW74cphftDDjikcHgLhGB9Qpe/BXPL4tnlraoR+aLnoARFbXXX54nuUnf
YwwNIf2taKYfV4m+Jlspg6YE3HLZQxGhyc80rG1hxIaUBa41dSaQKw1LH7yX5NsI
NnZBY4oqK5bEZm3UDmEdysj86Q3T+/QjZI5VCdv4nWYQDohZ8pR1IKKPKXDx58dU
3CIf+MQuTXWlLuwZfcPu6Iq+bKAxXciy45QToRl75v0w0bwzXa8Osi6nYWyIr2m8
BOgC30tjlUFfGbHeubjapbtBqb37N478sOfZzAmgF+8Enb87jCuF+xhlKuoAey71
UcJJwz4B4ZuspsdfcY8QHWB7cSf5ft4UIAyN8ASMUlqKV2Z9exmM12+Tzz+1IB+/
DZP/83QZ1DGqsCuGF8ZGth1LbMJE3K45O/kO3w5BWnvC5HASBGdar9niMvHz2oBD
u5m67vIwzw3fjXdfl0jH/98kO8C43fngOBSremlTWEWKXq7fxtuvM0DMueQmB8a0
3F78fuR8a6GCegCJ82xtXCRt1dlEgEz5M2Uk6kggNC5YSat/YF3CbOeQ0NYk719Y
nrp1hcVZs7TT/U4H8npLKQvM2EeMwrVV5lTVTHwqVWCKzaPV8/cROwCeQFSZ7KJ/
IBIrhMUCYA1cE2GCMREACfEzQlLNBJNY/9aKgMG30Q68+s4yiOP9g0pN4+6b5to8
foB44zU4hY4lO/kdPw7+P0Fak4wcd2m1TTNzF1yB1ICVGB2NR1RzTPwS+zFtSht3
U/XSuSE5dG8sLgghDBude3JrOLwXsNYQenR/CXfhj3wAYeyeqe8PTUtZJuAWwd6w
mxUTHAnPy1T4P0OhsmGByizb0VJcyaUbtsrKWnsRmfAJuLYaeDUqqD51rTvJPfRq
7TiJxfhFL1bFH0vZLaih2QjvCFnDWFKHfGTWGvPaYj7Bhbk5ro1zXkG2XIoZDg32
/abkAdEldFaAojpCm+bgygk0ceGZupHqSoX3ujEGn3CX+Dc3/jo9xT8Ij12sSOM3
K9tfWALaWe9OvfrdCdrNOiowxmtFsfoz/9wmufd/ypMpfVTVa+XWylzMc3GUXIts
IUGLWAXxM229B+JA2ozffLbDcKMvoJSKieyvCU8SJfNqiobQRb4d0KrjMTVbO1Me
2n6rwiLtQN4bzOPjql2Hr3Q7D63bMZG1pkQzERXICLrH/nDrX+PvW7UDzKrMhIec
8pWPp72f4i0LW2wdFG9VHrvM+z2bJX3t+R4pQEveFVuKplBLfJkF7or9xMzd7Xfg
gjrgj5ChByNiuGjFmEz3OUdCH/RTCUf7uebgAZS/3C+9Ju0Q5t65oQXtWO8ri3+Q
pEGFh4uigeMfAOxJFR78pZXORcJb8bNtop66ghwfWRhdqd8pD90vhYq3Zg7u3UUH
lc/KIRBNSIFhB65QUCI3X6KW6A0izSIhnJCuBhrn+vYowS27h/uox52P5OnYv1Ln
gtZFNTh7zR1b9t0TH8O7jRzocHS5es9J8sAydSS53ZmPx8pprpK9rP7DpQi+B1bF
LAQ4GHPU9I0hAroxHdb41QPlA3pGo4onvFP4wxEG5on/1njd4oN7Gs+6o1TYMSCP
bSfbiXrD9IWb3bN9NWVU2A0NsSkQwOQ+c8QdBAb1iWtHUGx3mHEqSlVyLRwzUpB0
TR0x8rPb347XMLbOPkK/SEzD86Axhs1qel+GyK41ubAfL8UrqI74gciFzF+OkVtW
37CKM0SoPhzdvRUSB0omvj9zxubNoIphmMjL/q7Kn2oi4P52BeRPnaBBVISlxjZn
p6T/uJxvzfnxCYw4VPQg+6OPUbr8KtW/8kW3h2PdvQNuNYTsUgPAGobmA6hhTr44
qP/pLC6WUw4V2/3Bvignk2AEPQYdUiUn/myNI50oz+hhtKuMaxQMFObITNcVWWPT
Ozk38McptootsaUBqQlo+pkWN8dm/SB7gbGDfbsS3OvDWfYeAJ+Bd609eOz8H8FA
JMOFhNYSjnuGkXF6WN03gvZAQCtxRuRoUU9SoBl6cPIF2hxsje24g9xjASEm4owU
kglWqwqOlsoZV/YDg10CNEHnyco3p+kov5JF+q3rrJ/H6VSid78J7QtIV083cZyS
PbvmOcbD1S/r7aJKoGqyDRWxXV5lHKWDbtKeWJOp2HwP8AWuIYfnUaWrARNjWrOA
lDQKp0/gPLXVPMGuQdNQVUdXF7gpO6AOAivZI5L0rsBWlaTUXQvOTgrNeJ0ShP04
V+mNfb0Zxc2dhTHqByX2Kc9bhao3x+0rNk9iT9hGKjl1N3o4AF2acUnbhX8oNcLG
jgjp4gGFAb/JSdhKNRIQ01tVcM01Jtew133iUBm9SowC67CWIFTpm1myIzO7yMKe
1Yd0T0cofdIddDFGDzSSdloH1HcDD5RMYxn6JWdppWzovfBwKGNEm1FlPXrrRBHz
DhJnMaTysYbtO2MuCBnCVHq/hja0fr/RXZGLEijF6OaVdJ+LFuvPNP6aW9SZYIfD
PzDZc0J8SwnmqhNcKrstqrxHEtRCu+A1xhVxM0q4VNrK+FaZo875yxQA3MWMFKUf
Cjd/VtHVfLU90RxhfsI+w4nvhEb7jKUkxgtwdw7uFTTBTN2T2dfYqXLnEjaZ9wnt
ViV+jZIRh8xEiNZ1r4+m1ByPoPTeOrx1qZOxibJqTSOL+oA7Daztq7w/oRBWd2lq
H8zMC/yDE/Qn26sCEUL94fR+DwGxk4iSdpAHhzOP19JjpAhVqbuFyBglt0jcRYrV
rcIUZVYIqPQdg4pRUDhKs/oT4SeifsGz4pWqfGIbE6xfKZITd2qolJW/jwHVLhOi
nHmOAFOQfz94Kz2dFeWOC7aoHlpY2u/kvqQvLorDjveABK60+84yfMFV+pCmrM8x
HkT8yXojhda8EELMM+SEgK8hRWpUAlmWRtRowuvZVDbFWB+4S1dGp6Xy34ITjdE9
VrfLXU5w8ci8h/t2PLqmGgFSry3dMwDAt8hGsTLDd2MUxhwTG9g/p7EcprliaEge
DE/egCr81EfF/0+vaVMLs6v7U925i8ns5Y2jI50e8kXVdyEc4kwAl0lRfMnvXYPf
PEeuVNIkkThyrzUzJHVPiP3RkXecuyIBUiEvC7Npyl5HjiuuFxAMH7+04oq4ahsC
nPBzsrtfSI1/SI5bMX0bsKjaw4rR9Y7k8uKcFLi5BP06RXhVJ2nSjbMSq6nO6bA/
ntIhaxXzCrF337G3PsiEHhJLBhsswW1q9MR7wBVsu5nn9mYaJjjExKW1FI+kZx2R
lfLebb77hw/c17afnmXIl+ntZs+Ld/CfihPuu1mQwqVlipUCQmYCFBSVSC/UbkYn
vAOpwfc/ahZt4UwngYDKtohO9k5DTVyNUfXGnyWrbZyV5exUxK0kZOXwT/WbDZNR
8UkcSFMWXLWIxCEOg4DJAUn+qv9O1CWwzomC8n2xNsWkXt7dhb93/l5AemxcZE1o
D+K5uEWL9nhAGSTcr8RfKCY3PL6I1DB4FYI09HX7pilAdBMLLOKDQeDqcd2RSdfp
C7nVH3wN0Njm1b1cbqkxJyrsRUZZaIApgK5tAzauidALSmuqnl6ulg+SdifPLiDA
U02Xmf/9y1bNc1PKLvfqL+ISTIsAhN909wBIk4IYuqCeZuFFiEEkp3DFs5n4JmTN
YIR5y29hYgET+IRei7y1aHQjh60tzhPabYd4IjqHolInzG/UTSROd4Vkj68dXCok
L1vIVdWyvL4Xf/SV7M0mNwwENPxaWcSXdtNtH9TaDs7he5yVJKQ3zSUtQiGcE8VJ
1Q84F0DWpnIvvlMgvyZGtjs7jb/pC0jjTrmT5ZdqTji8GvoBkszn8rZkgWG26F1q
X8J3PJ0sN3ynX24xJfUJmpTFhXvsthLcIPpfLnigP5fC4gxUYoCU9Bm4Or4sRtNh
fi0WfpFycCMdoCMKwjwFPBNQ/II4Q18281WxF2nmIl4kfjQK23QG4+eSxBuRZ6nJ
FqDziiyIT1nadlc3dHvUZJkE4BnB7w2E2McXlmVNsMrsF3GZVWWVGsKOykBESB0W
X9B9wgI6fxLvRooqxylMQAff3Vy0KlYLRtdk1otPkTicgzUTGYG5Baw0WVEL9l4v
4Bed7AcVasOBcFO2YTiIo42LK3dVcb2E5XMkFnya9WfV47tcylR6+rT+WibQLRkD
UhHlhequHcUJxsizzBdoQEYZTB0GyfBcgNmIhJtFGWzKfN6s9eE22e0coldNmLYs
2Tla5I+QfvkO6uWb3MXGDsoZdtEDxM3wivV8fxxmsAkHlu5+vi9Dhc5fiN7vyECj
H17gaugeoZzCHs+z1eUSE58VIpsj4AudABGQdOunVQD86uD0Zv2g4uHy5ROAKXKS
fiacbMknoenjS6iwXreqS0QwvBrY/Q1+1q+Q6tnJNYu63BBoNlJ0S5x3VtJ9fZDR
BsWh6oFWf4ggsDNDK5JwtNfQfG7rpLAJaY8bH3RNyra4i+aCn4gAUCBaEGbzv2Xc
qH8yoDovyFrz4J5e9cnMY731GNaUMriFj3D3ap3uAKMPkLfT3OvVLfHZlF6TpRjW
ZP5ilbx1ZYrOLzzG3LkTpADwR3ebeypLv0gJFR4zlJpKlg50Z/MA5N+44jr4FEMG
wjCQhT64RIRbdsqwlYEgwejj2NtXcUGFcw0jz0hTTXg/y9jDljfdDunHmqo8q8+h
KSUiM18gvYnFOBH4eJYGvknJt1l62l/cfwqKK9qaEF2Ewsj8onfUHeVsqILx2GzO
fKtmSFO2xu2qWgY4530E1isDP/eUCxw/BVwUddsr+PfTnuy/RGsP0cqL2Si4shqU
nBBcFRxPgWmObU49NcZLqjSa93iQ1mhFmedOAxYPe9xDRhX2qkt71TtWzAidpDz8
WEQJDhGCYgdBQAub/zr1UuFHsfu3B6ZOM7/tiUZw1gS0lMLS8BmT9vF3wWkQIG6l
9/VXAcV1r36JMyeZ5wxG0VHyEaEiG90/+KpwSEyM63XXE48w3rWuZik6fKmq+w5t
F784vOcPfzy5ZheUHHZkH6/R7JUCb0GgbaXS85S3nCkweqRStyZYQmDrO3Ez4QMz
4GJvmY3p6eFxEaU/iej4fjJf48d5yG+Wxn4qtXpGZKhLWv4TxMX8ipSsGPV565mE
TRLfIKPwHoyLtWDjO7r1QpKSqCVRF5NZixGLN7BFqNPmsGW+8JT16oGBscpgGthQ
uQThhtSALZle0AdnyIaCGCyKQ36f0wMwSvPAocoSnhDFZ40BtxOAAHvjmb3MBOUl
igygwOGhH3P14O3j72NQmFFsNbs8HAWCAGBGt15rjD+TJJBs66ylQJwgEA3rYPMc
ZDlFt9Q7KHiW95IJ7gkWk5T3Ms22h+6BpH6d+ZZjnL6RcIllHKZ2iliV7uyvU/gf
5X1AY2wts33m3IgeIl+jKX/elGWqen5AtlReVoEVuuhD9gM4hZyPcGMA6HzPPN/R
qnR2qkbhJ+iiPAZ8ca+tsVFbR69v63zjY3ISDA+xRDHRaaL+7YTdijVxbAwkR7gx
+x9V9OSQAa1sVHDBdo6v/UsFS2KNPFneuZUZbzAj80rksu2qYqRPoUaSj9ysseb7
pfqxy0CnqugdHrRKeBiWXHIzqdy2+npInMOOwjkYdwAQhxuYwsz5E9qTCmMqMKvQ
oxvmpnHl2PiANTEz3Hl09tIWtj/L+UzA12y/L57+z9XzWOWeZS4CCfkaXB0Ve8kZ
vCYdAhaBj4dew/qJSN4os3Xxv4DH13TIJ1jzHyJ5oYLIHywyqjyIJxUGGD/6tLB5
mLjobvgjCBQsLg3k+vACU6Gm7do4kKT7S3PBbDNVVis6wt+zG2YYContjKUooU0X
ieEuhZhAmQ9i9Tx4XTY1bb/s+oJrgku06OTRwXups17+jsNjEqcSval5q7fQzm9F
CkM3aYn/u+jzL7A2MdKU+jGaFPFuW7FEe1a7l473qSB6l8TWLPuTRWsM9XKIEPFz
kjBQ4wQMWEiklBH8ZKCnwNqFCnn3XpsrrTbvLGNvs1szjINcAQuvXbHcuBRk/PiX
GEHCT4qGKWB0X5ZjpQxxHurHw4wHSKbQ5hykMz0ZhXHnAT8FfVv4kmb+PMm8G2tA
rmlLHjOHum2rZJahu3CMne9hAM0gng8HRNrT48xYitU6cpwqC+9zaOVfqszRqz3l
8hnfEdkX5snstKSh6hDhy2O3xDK7gWrFTtRAdh05hA9iP1P5BIamFeeYqRHxdARP
+k+tZDGivutuMQ5ryp74bcO1SEereejuHv4qdB5yA6mlgKUQX+CwTT5WMvuEQqKC
uLO8SfzJkIvWV+Rt/Q+8Of2JIFOeZ6r9JaxQfAHWLFRXLrCzpDEdI3+sPPnBc9R2
2ryYgkwnugHE5IrC6ts6H9akr+k/o9SPfsTBW3+Ly8obyK9/bEQg8ZnIrHOlrPpF
aXM2qAlwU+cMY7FCGGZryXBTgZ+mT836C6Y2F6KP6tKOCgGH24cKdDcuSIGn6c6g
xLjpvNlLGyC+grkCUhz5yAUjJ14EBpvMfZtSbAghvwbCgOSd0QS4SwADuOWnY/Kg
7XHpEVUEKH1kITSDBIG0g8U5p/PdP2qiesyCKH/RpfG4rN3ImSIfSyMRq7Uis4NS
MryL3t3ykQkh/03fP93kmrfIbMxP0Am0Ic0JI7JEzc8ohKVy7NpUtt32yDXIT1r7
Doq2ahvX+sv3lsS492n2xOZitC5Jl3aL+w+HlhIzWKiW8ZfH77pG+eBSXYullrXm
wxnroNvITcDz3SQruyXfEoN2feCkqYhxjmPVBA/KtzNTHjcugnqD77NvlUNHD3Tq
BIgfC6ix7us8AM7RKGDSs97Bnb7mlz5DMF6Ps2d+91FPZti3PgOSSiGOhDX9pbn+
NjkNk/K5CUoRvW07AU8C0lWc43BlzkbLCx1Ob9Lwf4hY4Ba/vZWGhMrorAYL9BEg
BBomhJZYNwUsJ4l+09yCcvORg0U/yy1iVr338+sHo5HCYdOa2WuOnYs9KSPq27xc
20P+HdSWEcMJjdiTXWmERXSyHjwL5p19AjO9T9993d3EZRELNbeuKLzpYTZDXsTE
NITkUftEJDxe7EasJ6yUnR7Bq6qAFWcU1xv/WDGyrHqHDzIw22iuMLycJ3geU/D7
FmH0kE6s+CzdM9MgzYqKBZu+wVx4rjPKvjIe7SZpkTpAvryO+ydFvQiUUrNbJU+z
mK0JBFwPWV05S5rccqY9fJ5LoOqIINmFTyEFquSvNvHQQ+HwpBRVeY103IKeXBRh
Er9BNzd4oN+1rR+/O4klnddAZlcjgcFR7Toh95H//3Y8grwxTEa0rTQIy//tt02I
+aejc+twKW2JiNxUEqTzH0WRt36uIG6pP5jIwhJrSJYfcx2tgwBqsyBOb4dgkNEc
JrXM8qTYGHx1GOnplt+n3FOigtS+ZmbOo340V592xCqWccZQhidWUBiHE/G9XwAB
XyTxANXsrTE4wDO072Ns8bf9godRjXltoZ0dF12+qtLYCljI9KTLnfMPmuX8/5LB
iqZ9d7+rh2aAF5CSwSH0FJIr81ZigjNRcCos5MceI0DpMrEVp9pTbFpKs8CEvJHF
iQVoU+J8gp4yf+aCTWn0tmFf7rBsQdadkGq+HBHc+JRrNrh+YldUCp/QEQHTck0Q
pLpHzbDX9g3D87PC/Z0OKgKdaQI54X2cCM8Qhk8BV3P6oDs9UA9MYrQpkOfTm4M+
xa8e24jTQtqnmmeknNOzq2A3re2BI9qEdzEHfnokD7reNLDb0GKS3Gm9xLC4xVFM
lXVTUaj91WUC+B4qP9wgGhI79GxmrYTO9OrgYEV4g57vnc1vb3G88BT+Vr+6Gy2R
/K4AB3rrbTNQl+hg+LWFde4r/1JpffKnGHqcJPfU7kgLP8HbCKIlFvhrAbNYqOVc
RaUUnvbbWP39LGKh/SLJlvpPXFOnuSbxcR+g6q6cv8XAwCQLg/+8gwrb/awi0z3N
PDYuXffg0Z6YlM4O7mxh4Cg2Bskc+GhtFSrPUdWEtnGY2FS9rLKvIdOtudFHbYgv
Ku71c2v/YN03Ws/0hZFTLks2171kXw5MRfnt19XBBkvaXa44H1PydoywaLh70Drq
mXCaekl7lRIf6VioxGaH713MCgQ7W5YkOP7aFrHDGH1pojpnnpS0x4M9Yow/kEuI
f+H6d3zGj6UmwAC6POpgI80RRjIwOUpwC8K4aX2fXJkG5hA+zopVE9ewZhFvcV1C
H2EblXGbi6C93yHWPPK3DeyxWIt8h0Y7gY3JBxQWiUr0Nx6z00ZGH1HkLd7N2XMR
99gaCt/JBsxnmDYOW6CBh5hODvqaOcib7owzattOFHKhwkHza8pOI83OVJZZH/P3
AGXmNW1fVuTcHU+EX6vZadwqWzm+cOLJ9koLzyHTy2U+545N+wvVpis4OXJjmXjb
7FeNJ6EkabHoRgsPMJNKiPEYZryV0X0g6y2aIcnhw/1FWcyy9jRtdLy9MNRCU/2A
OOF4ZpRavSMz1tYtOKCzG9NucUhPf9Ba9UBh6W6MZJKacAk1t+fNTWBWNzj5RRor
vFqcis1s8puLVSUghSQYWoeT7XURQUFvacwcKIOyhCDmFMkW1X4HZN4yGwLixLzT
UpMtBi3vMNvin3dcNpqb5ALTndbESMoHPpv+qS0+sAppcJ44zAUoyJhICHWZdGif
aiE1E1ggnCCyytbUYngtzAyS/+f/HTHFj3gv6zfAxhYfsvrj/3C5KDRutfFK8/sE
EcK/qwb4xPrm1za7pAIeUuJQG7QkjuRiSeSB+epob5onWy+A1u56soqpTG2oNua2
z1v1+3UKNYc/rwQ5PD2PdVTaQjJpbsyGe+eW3M14cMs1s8RvIjh+K50NH4Qdg7Ut
EV0mIAKIjECrJJFKOgAuGfgAOIapYQpP3r0KAUdajhoLJSG7McovMwp5xLDE+jaW
s6tBG8hry4Ug81IwW8vKGNtD/DJbIBTm0JTAdZz7YmxZ6Z3KucahVUn1EJkExLn2
6F1zuLKjnkucZswXSFvHmmUhjjYgwgIQh67OtmGB5IRlyM8QKOB0VZhRj5DENGSA
yIcB1N1WGhckH5Nqzj63pLBRRdok+KAx5/H3eWgia6bhh6oykJ6qqh65CL3ulYfp
k72EDDwNo26E5ZJTcsO+KmwEsHH40/2e+LMPLcE8keu0gHzAtQWFIeayndVnLFk6
WtRNlFzkcCymJXBgLZ6YY83jUZLfN0Gr5KkFiUwMoloPPLXfnL1Z1lNnq8aAQPqw
1UeSA3Qj53z9LGApf8KZ5fCmLJht969Yn8hjzP9i307mtTGaGvObq+M+1BBH9iQf
644suAQO8m6U0SIvQtub37sAomVaHRtpH6L5fbkwHFJjxI6qw8Y0wjo4f+oFhoJo
j/ZD8BGKdSgkUxqkZ544wKH5e7C9YN4IF1xKU3v5NsJhsteDTuNOVPuxby4PWgds
Sly7a5qU71DmvLyVTY8abwf/zPXvyh8f1b1YLlj6pfIrRG/opW6VC9CaymyOnJjc
dWuBFaEzfbuasWe0zkQmUSDFRLIVXPE4fpK22c0ZwkLeadiZl/owzPtHgqaJeUxz
fYOkGZ3qptGC1q534vBOhybR+3mLn47CqPRIPwzFCWNDw2ckBbatk+ASNMa2ynR1
kSs6lFtLBDddQw2IsSiGWpUpBTSP8jWo5Zzecu9gw2iAeq2aYxAKMV5suenz90DU
PQrF0ZJWWmt+61MrxyHDwjokafqzUMhsrCFKkRnIVBRKY27GaAjKt/5pmfZfqn2G
abhBB7qQEMc50AyPSV/4IjettigJFI8MKU2gi9aqHprzSP10MmTDHntYpJ0P7tEA
7x1mQeMkHjU/9c62Gu1xgfePGp4W+EeVYnzKKfBd9VATXn0E9lLk/Q+5NAzKK0I5
ugN1gEZPnWvNfvg4dXNJkcjIOJtffystHMXjFcoB1nVTs+atoUBbIcDXSyv/bZxr
Q+prGhFsDOmynxGmZ19n0A/ll3F80fkNnXbACkw/XKHrRPGlkUTjhgYxaIt23Kqk
MH58fsVhSGXLBiROEeVsMEf/0ZNRudOP+l2b0KfSS0adswRoUo4P8QjibAgZt+sS
m3YTvHdaLha9vpxHTzzcYvxxfsTYL1m8zkEJuxd5QWm2wflWT28v0qj9vH4sT65B
jWykFwbM64JzKV4c0mev9wZ8z+KlDJXQ6mlzPS4ZPePtArEHXamokOafRmT1d+3Z
NuuPA0MyO12xbduhirdePUfacMzHdfTnZnlpwCEPZTIm1mrMIdVo9sNNZojZpyzg
Fb6Qetx3PJwihunY0CVHZdI/L3dmaZklAB2T7oJdJLdHqnyfjl0ojmL4oDeYd/Uj
qsxLbifMZHkmqfLy0P/3gEwmI/bZHbg1/ZUwRm81kZ5s4PV+L/vpaEsO7fbyyOeZ
boH4gv8qvM20eiihhgead4mbbRYd6G6xNxxQ8RPQpVDpL+FKpcjaEqr95+UYfKcW
/TIDg/OaIBloMhGREOdIIYTXT3cYdpnRzyYp31Vm32fP5ahRbYCW5Nw2oc67y/2H
3iDEheG5kLGSm7/pEshzUWWqD5o6tpLvwMz29RXirzFhI0v5PzzHe3+xz4a4/A1+
rtGJXOEvk01gK8r974OyDNlTmNIsejhjI2vDaR+BLOG8of67WkZW/cJ9GguyS4wv
aLqoBuwbM0+iw2BkrCJ8x/Hl0KhfB+DrB+i8UJd2w4XbtlEc2VK9RBLl4jEzUq3i
fTiK1XHhWjWHbXb7MR7vaoWSMtKZIJ/uqcBfOVEJ9PL3U/Vcvq3WYpuk6SWYn8ar
e7H6jgCI4skJRZOQ20tt6V2w52Npi93IsHOjtOje3YPa9RMK9nQg/36xgFoMpb5C
+lT6vyFNEPQ5L0WNn5NeJAP/5P60V5ScftSQhQ1/AcAuXruBbMi/D9oQvF4jdjCm
h6nh1LdsRZTdBYl0OavTeL9n8CAVJ1vIMFLpZoWuVdupT86hdw38HGBWs9gjdQX5
zrJZKY/2uIBb+66hJOCcM314E0bSk7J48RJbFdv11HETJjWk0yI11XO6I7EFMioc
HUKm8Kx9QBdGIboz0MR2267TFaPhsmrhrDOQmczeuuz+pvCWAD+uNkoyaXGremsC
4ICic8yrJ95SixYJW1sEO3NiC1UkhZorzFStp57MO8QBfyvmLC/zjjrYWBFTGtZm
z97J3IAxTHLEAi7JusP9K0wE4XpXOmQyRAkwhrl9rKZ45H1VbctjjXVPBFZ/0FIb
WyG48wFLMxxxRINGYSr3BCumpYwbZYGEViVEk6tGz2/JWfMkZqfee11i+8IPi/gh
ZUB7bKjtXQQ7XSp3Zdf2gq3jlPnj+mIWjfZJCoocghBAMNzqSKC3Ukau+OgJs9Yf
qBiSdO8rrNXbjKdbFItmgzRSsFPtUGyNOu4MXWOCVrRcECc/jk89YLlLOyrZx4sM
GOQdAzOeU0Ultb5Og1tqOkabo+ZXYxg6ctwEsofdc35qas82nSRb2LBT7HWyR9LI
9i/6wsc+hbY6ijmBBqZzU+4X5hvpCXtuy9Ruul1agLflu1JpFMTCk+S7359pez5p
ybfysLF0GJbKTiNQtXWhAPbUroiEMtkJyxR4k8M1gmcR81I8jBba1RXEEjZy70Qg
ODBq6u42juBvB5hDAxrXMRB7AROIc5hveRDudompj6nW35NG87Dh/IbsUoJtWIey
ZWwq6lLtf+fxxl7dOQyLvY1omR9NUl7TBrn/FkVT3u1dcqQjmJknqGxVPLiOCKmY
SImARgS9TRU3rihA3x4yMXO7iURostQJVjvemGO6DCnDnvzzu9vVU4mRug0wpXQl
0JjI+xBP5eu/W8Ai18klHv7P3pJ9m1xZSP/59AFPMNQwDNt8zBi9T/5dMeBZR17m
kiiGb/hzYneSgnsjM8/zFfq6sl/whi5xlNbVom1Hh20iCt9hWX8qsy09FZQJKwgB
uuNUsARK6NmaVHdjc4YAo6JsFGh2t6A0b7IPyPxE8/a/6Gsykg/MK8TJ6dZ2DzFP
pILpfKRDv+kpVVhewutaJsdM1fx0ZvUUhA7empmP2Gwvu/rPwThTx+3nFzo0dfsc
GQRxdHfBVTSLX/G4GEpxta8qk+yI0V6kdRfaoheMh4VvkBCmIYWMY0lYi2DeIZ5l
EWF9wGrNR3uBb6vIbYh/eilrakIRIje3w/E//Hap17/jbqVN+VoZZAFspD43kFx5
ozFeOAS6r8ZxGq2pumxKRG1XJyhk7yO0lLG0+9ARKv3YLf6op8UxsgK0DysyUd9j
sKK1/KiDkR256je4BU6Sg0qA3sE7hwL15khKHqZwtSsTm2bNp98LpeeMo4jAxhjA
V/YtBO3FbmllVk806+5eT+9NGEWep/MhknUD6cd1uzc1R3/BIYAiG5bWDv78bq/K
GjXj8GU1upgxvltCRDv8Qi9dK1DdOuVzaUmSs3/ETY47mYX8/akMnWFpkXf1Jxz2
AQ6ntPkctW/CkDtqqOOeRJGh1AicPfILVzXvVqK5AOUOgEVLc9d+JAyOfmk8FMJl
5R8H6ibD8f2x8i27MEczZNLgib0mbpTOPZONqnr3l6H+EUPDEex/FPUDQWgOylEj
0KsC/WoImEU+237D3ycz8ReAPnHtyjcrZ5bzDsexCMIDuXVEg0Cg8L2nH258aFjq
Ag/6RNK5yulOiTM9EJZ8xJzlj9zPEQhiB8ogG8djd2wDEy+wWLLNUcTy4/vStDom
2ARiOlhiRvWIaVm9cC6eMMsi74k1+yFQmmxi5zzXu1MOlujsAgDN5mQArr6L4T+6
XD52axKDr0BV0m1IadcQhwqZRRgSqt7eMZhKbQ/iGcXF8z3jn3A7rwo2FbQsG2Z0
AFJKY+Hh2X5clR2Q2q5367lqXNrZL7BKciNWecgR5KxUfenXJdXsm09q4SEZwqvi
izs+dTku2saz128hgUGCn2YJXVhZDzBIdLZVIF4zk6E47NukAcocr/Xxft20oDms
dt44qG4UQGu8T9w0rpLj08+Ru8ui+f3ePbkWnfaE70Gk64W+KbQvcODvuTN4whVu
6tORwbjrzT7LC5ulkB9Wd0Ce1wkJ2TO4tN7oyHh6QDsNIYw4mw0ejZql9mS7gdla
6af/3CHW2Mm8r/Z0+ZiJFbS/K0MtkhjL6UuKLc2IkHcg9yfbF0NF9cp3nodPLD7I
NslfMwjpRiYUJWlY/EWliNWrNPE9HYq5hQZqudvoGdJW8Co57kVRpIPysvVuAf6c
PBGm4TbDWOhlbq6oV+VIJtNmDhvfvi23pVn35nCVyc5fYC5iksSleT6TVz0tBThP
DuQVHjDJ+KBD8sSGX0bWJO52uog4bVYJ0J6mqM27ORVrEXsmLU2ul/V4L8KEDl6Z
99LBamfA2IEVNXErwdac7Rf2Kb1zySN5gUfnv7rONfGDOakroTBJn23mJ/cGR0fc
cLrY57XvWAXDUcqC7EoJoZ4jKtl+Ezlsu1Tjbig4t9xTP2sly0V9P/Zzu2NqsPie
MiRWc+S+JMzPgwFk77GU9Jd2v6uq40hB+sQgVKWkTCFIO4PBTtbqmousq9FVmi2R
nS7eP5oY0y9VuDp5aGuNR8xXEaLfmVrS6zIG4fQYhQHv2CWCcKJHs0EJs7MnGb/W
SB7kOKb4sxsnIqjg2wYLjiokJgfJN80lrX0FpKhhLMKtjf3Fy/jSXbpsPle8eNg8
St05qEpVklT4Am21UemQbhsraI4+8umRm+YJKobkOp1r7uTvIkCTj5G0wvyddc8M
ZxQpDiBrUmevaDRBSTagtsVWWZaY3txZyn1IuTLKvc+X/OIJr5R+/OVSLHUJYS2b
pPkG7FF35Qxlctpk5mtVO5wT8CP+JyxIPT39r9Rr94rlXMpeZstlvezHJzV9C5+A
+KldZlxc/YcGal4gV9uJL91TKymbkXlEpw9OMYB5YpWn1AbXG7DtnMKtl6CrWMBM
Ybx9IRP8Aq8sAgVHYRcLYTJiCQVMVW2cQqBz3HivUGy16ARCwGuMpBT+Lrk17ytV
ABivNt0b0j0aDwsSpASpcVqOMjA4hN4RNQGrUCrx9diU+hVhK58hfCnt3KFWQHXO
JOhqyz4Elomfar41NvUOpd668qXmBuBKulVHoKvJ9O9E3hwahl0/hsF8KR04KZP1
aWVFdQ6uBUshw/uZ2L13ETyze2Eg5TMuTi4LFXNVg2bXagfD82Vt/FfxRdoW3IbI
68NHBhDKSGUFCTEpC9KO80unbpMaxtLHRXhXKeawdTr+D6P2/0LvTaPyAjJjh+55
YCDdrBN+7G9MtiW039VAKTvqt/Ugwyj0zz4NclNuVBORBwDvngQ7j2BJNraCORVJ
MzxQH5D4RhbP29a6Wq2YnRuyeZQjMJAo2Qz4m8d8q8C3MQgweGQYD6r9Iu58cRtq
jcFr+7ijLF+FfABxCLmuAV6BHtDnd4dIVofiZhrIu2kgnpixjSt5Wkqf+MUibKiX
UEOTcc258VSS5QT+q+pQEFM9zvBEyTSwM6AsWbsFfJc9tUGSVpb7cuaOTU6TMJCP
Fb/VsKhMzYvDXG3gVdmF6EgjqClcv36pm6sGKYOMHA7sXVnf479IS/Vzx7g5r/zK
TR8J2TLthLuR5l91hLPaNsh+s/XK1Hkg0LwvpgQK8gIzO+ygkxNpX+joMn74tG/1
kI0JZ1OPQwlUnueGRGEi35b5Zsf/pXa6VD5A5IQb+EYX96MbzaFwgjbhBnI3XS91
BI85gsOGxk+sNJpBzS+EFZojal6SOdYDexP/7yFoeW4Z3ih0n4+RkSFcDdAV/+QN
HrlYfR9M3P98jsn3FH5ai46f2d+6ZZtaq3pAEO4/AF7Ck9gNk7GI9YzAkrStHrSB
aegjhiRl/2lDbnjZQ7n0JpBp4TuuHQKVMz3z2ltry8X+9JaQY4JkQ7ahgZcSTTAN
KzWxMn5wSXO0jr8yEgUv7eRYYZYlwaqq+0H8s/lAk4MwaIh67V8v33l5mSCfD9vT
TGfUt2X1icDlTpm6TdoBt571spDf5ErDgDTMI7/UrvB55niJQ71goe4w4aqRszKS
yQvQKt3xGZmld1SEj4DDRdeEgd4njQAYxG6ZDQ367B4ZVkPfZB817uxtOHZn5cpq
0BMEZrWr+DCtORWHZLB/qahpdj/dRJdWL/FoSqmisz+xLndL4P/5mn0zRsKsJoax
CUOokmDtPF4rgjQ2tOf0sl78/pXKmWKR50mRKmvWc2tgtLMpV1xM+zsehlwrmmPT
YZx0T0+q3RTggCgYPZ8a+HDwUW3MGZ++awA37vrV8Sy678W29Fe9nFqFfHzn2Xw0
t6dhPrm9vqOj17hCD/j8UPKLyEICDNGknVapDIPm1SDMK5oOwCqTnGXsNpwaeEHh
3ylTAOwsyJa/JB0kXrfVxX7nZcwSPEGoNQigRDwH/NEgkGcu/cuuj60aUFKhkv4L
DJ5SPEdCC9NOszJqBJ5a+A1+SkgJqRQCeDBNQCrkrU8U3gPmQhoGjGXpq60IXM1A
EYbdKbK31+WrnmNiMlQwp/xhAmG98YDwTBq2VCzGeommUDfuABuFqV0m9i6LaBo8
WKdGGnq++PmTu/KGoaiJMDla4suC8Z2dyoxWFPisX+DpLT8rDf0SWNC2J8w4UZC9
Du7ZnIhT/cV8+TUExtmIDPPnNNiQBbgSATyIK7FC6fPwVSNT0FpyTfFb4zY1bnPa
a0eS32wWMgRXqNv5wZv/mbKRqkRq7e/Xm3iVpsry4w3VEEk4o+K1TTFMo27Zr385
jDb5xKecEHnHeQsLRD9USm8enPO+ZKYKFnboXwhRRuvu1rkJeLUGG8lZB87BE0pp
AbfbaJZgpcBrKxBX44fpi7klFWB+3Q7Y0AyAgJPz9hk9cZRRafejws+DuASX/gD7
bdZrflHkyf1dgIWi5bS3Mmzkjik3H7yCMCMbIod/JHMtpV1EY3vn8uQHaN8cFrMG
ziVAA4wOwKR5h2X18+wfMXH7RHz/clifm7+Fhg4H1oemxS37VhZraeKxCzxwVII8
4CMpf+tFMLGTd4pFgwO5g0KeH9ZL/rkylsk6zzh68rmsbt9YuTMz/KNUy623rigE
2LAETXSEYt3XdeoMbw5OUHaHUTmYhajCOouXYtROpo49rqSN33mx4VYcYS8ccc7L
aPPJQOu2BmOAiKmHw4WUgAM1aH+5Vq4rL1BIkzkow0yvi409vgKUd6Rg8zrhYV/G
0G2+dDzPRtliEJ0wwRR5PFU34zJgRrEAut0lNGCAfqWNG/uovRiMDkiIiTF/kRLe
bXytZINy39PWC39/xfT3HkWo2k6P5cY3HXz3Mk27r97WZiwqLEAbOtjzeCquywJu
pv/HJQ9tV8aRok2SKYFpUddCjM0Hggnm+CPcKLPV/mZF3wRkwFaHYsAdjWk3n8wo
fwVrVn0xUTP1NeCkIu3NceLL9DezI41G5xCHyVMfdSPwP7mO/jKeRq5xApTb1ZuQ
P8fkYV6su99DLmFUhS5awRLn7t+W1ccsnHP2yLuwkrBku4//bLG+8Z9bYRgWYhfj
xNwOiuy6eMdnLb4oyo9VOag3w+zdZMVRs0aQgrQsXN9it1/xwsd3xYkCbEaj4AMg
fOLZg52s+lenQDmztjmUzUJqoUO5FkBo/h8ddcm8M8UwwM5P0AcQupMOOUl356ux
Io+fihSeQf0LlNJecaX8YJMg4HrL5L6TwXWm6WNRIFmlR1HAGlOZi+V7W3E08yF6
bxlmV6nuIkQxUrjRgXvnpGch/nnjCLjHP/oe3xNZeIVQKC9aTeQXOu6H2BhRenqx
Q2eLWObNSydSIlk2ge6FeBpx89IjsjJZbekxnipo4T/ztQ6BvQLKOrDx/RMqXzlM
nHwmlN1yJuvey+Ulp4MI9sncqyCtgicFNOwIUQEew7N2bph4z0nawuVU7XjopF3J
8MmHwKjfdjN4xgTbBVNiC+L4+p2i9zTomyVZ9LxW/Hyv8DKc5EF1wSmZFVhj10w2
QS2P/HA87FtYi0+sgNdiCM0SgWL5/cehlkE7SlVPWVsaGQGamdwj/4np7IDDr3dA
nFsAjNSv7GAiil1L5tjSzuYOhNbcWPOccU8F5rsRYQRg+hWN9ry6eDlqs9ZTm3LI
bKec5SbsrnYmmPgrNSt2RS3z1qYMC+pGr5sAAuAwLl+qEKNp2oMG+k21A4DNvUz1
ysKgc4nDy/pqJg5NooLw9hHrWaexe+2D1yNM1fw3yQEL510lvIha1PJFMYyzKELv
PMYEd47cWw5Fd9RLnGq/WfspttRC/5bQiVjSa1Bw/BAuyIJJNjp3M5ZqpRXpNggs
f+8rFkI1NEl0vp04g8I2NbsjrKZhWjnR3Q5i/1Z3eyetApjc/QJTA/jsaiyByr7C
FV3bhlAS4Kth8f0c3IczkdeLknxdOP5Byyx0XMBwDV1fnJ/fequ7euGQN6Gyu5Vh
ASBTwm2KZfYwMWRtHQuRh46Xf3hYLbtLhkTAKUheAbE5jVMFTvl9cBf8EIp28rUh
rRlEKNq9D2uA/c09tfxxIX4+8S7iZ/RVbgQnGkZ3++J2XDj5X/06LwwkeTNG6Wi0
v8H6bQveBWTtLgJD8XTFVXb6ZUSXSTAPmTjl+e7BsW2kXhpXc0opgos0CbHqMrW1
JJ5ADvZkQp3V3lPjIyVxZZ2JvT7WZs9cjuRP+tzS4lyU6AMiwQgDYon+0lUeKVna
jk820lDcv8mpBubAtaPzG2hiiqI5kjIDfxuiQZdwSbcSZs5FwqXuexdT4lvx9j+P
bnqwWcPGgUC980VQ62fv5xUJLdOc2J4qY5pHhg8Ps0PC7UxjqE265hjuAV+TksJH
DkgxqosnKla0dRA3ZS/8Wm0M/etQ9h96+YpzBFb2WDlMsQH/9BYk/fMqoggUcEpr
9uLi2wA9ZcXOBfK6SsoaZMAIKffOXXt3dK1T4BOvaHxTpPfteTU23sWC5eeA4Rd8
zquK26x6RHUMpdBpOK/lsTH6ik6mchqpPKMaogH1glXuRNKf+n+3+wwPTMW8wINV
OqBkKo7qiXfP3GZfcEDtilMw5d54ePskPlSYiK5N9UFDgcl/0fOU2HCT1Hrq6dy3
V0Rm8GcfrOaTNUO4fK1mM3dYpKx9BcF9SrNfMsowg+gD79ylfqoDoNsNEKCIleRH
KWrTAkrm4NUrNc5ZKh4M02AwszYJEhQ7FSPaNv/kXZoB1mKYsqi3sW/Jxgdqy0CC
3m8JD7oa3xYapa4N9ZR8TchfNqkBK5gOxGYuJ5YWTi6gYmOtvAE2nur8OULlHg5c
1hG/C5A71873/cU/MA+r1xvQDZU1vda8z1FDGElAB+PzZ/YjLpK6rg/FMAk7bAsZ
wwzadkLQ77RtN2d49EeJOadcbHG4yGqs0mUzN6x44WtPMkSnlDLEsYl02Hq95bs3
DhOkxNZz3zaZIOXzhTmSv0dd0ckzRNfJNl4GQsa2vD9hbE2eOQD3rVniX1P/LrH/
wkJ8pXvXZwbP+M33pskCATIvLy3QJw1OhHhPhFgoNoe3QoHg4yPAyFyQ+/N/qkAo
VYPIKtwUfkwqTvxhUbShRwyDbjBr6NLXLOaQtF5/oKNjIGn4stXFKlkhJ/bv5VM+
fpdhW/1Zf2m4ibpGX1L79qcV6wvDu4miB68ZRT9UC+dqLPd1bLhdksS8EiJ6shKf
/vZZ8EjubZA9zvpWqWPd/YfUnQm8bRQ5DP9+gnJ4z44pYD8Mp+bmppWw34BaZd8a
9v0TlZJeLjERPeX4rESJX4FW1r2DUrTIBSud1PfO4u3Ni4yzjcYtfYDTEqK9zaTC
hOE3X+JDCJDeuMoNu1LBYSCMuVtUFvm/gDjjb/fG+OUPfrz78h9gl/Sp5R4UYz2w
ibNQJ65gOMQoXTxfkY8vCxK/CbtF4Dk0dxjN0VJjWmqcHt4r0b52+tyYpsxUc4E+
K9hNnhv3V9GqfV455a1st1fW0b2osmScYyDNMRxvXjrZVSUMpORlH/OeZ1lVNW0a
/iCokC2yypqr2zLSH13nZRA2AOkx4fHsKFzZDcaMi9VC5jQyKDk2W3Fd6kELiqfa
KZGSEmggV8ofmfMUjo4+7pqd8a1wmhM6ReofhTiS2ieDkAJy3GDQFkcXhZgZrIS3
/j+JL8hAwidjeb1rt50VLyOSYIftof7/ZWPXsYWvALU0OeIdifC4gM2kxGL8uzJu
IWSvw7HWkan0xCeFGPaYlRuYvjs+kVNLU72szxKb22l0BupL+9utYwIWfhhcn9y/
o9kPM7nouhv1MNp2p/D2TImn2/ekn2+UaWO/Kp9VAJRVskJxoKFbOXjxxuB2rIZh
eB0IEQQwuIey1nxeD2XHdj9+E+c8AQ5bJuAnvH2o2TY/Ekq+H0fQZ96UOX4w2Bu/
V27c6xPTEbkXNiMgGrnfyzA5PUFYUhyatJtJalIWS6OaXJDZycGQkF3UFgG43rMC
4izNFN+6HemHSW/nXmNFFEhCIVIDBr6oOz9aW+SxDSw7pK3Y4r2CJ71fw+MeyZ6e
on8AZkNAMNXw4hGIcyIhrfFxZjZNItj8l2KZn+KOySGQQefso3J7h4vV4rq38cOm
e71AIT9wakNJCNwTjUAFU7cv+65h5Q8BQF3dlmWHIJ6XxfK/uO0idx9Y776DfnA7
KUJKN0STaar5WWkXEcTk7xdlPjiBschJWD583Q+TZ8biOOIA1Sr+jxaCjBl2hyGu
jccP6MqjXkWoWIShcXUF7rJVIBG2jmPdg5vZ9FiD0lAtubEsCoYB41BDWDhZMXyp
kQcaXXnVsoDxav8BwUZZbF6RKnCcPrTU/7RhFlTfMea9nWHyodsDdq+ZtSF50iGp
S71pfGyhdgskRK5mR2Y5yqz0hFQmWxWDlaFBkqaWJILkGhp6RGv+jz1M/ceKVes8
FsyywBdySQSq7T3zBJzfSdTRNHX+UR/pFIArGyDcKhGRkfbd1KIKdM68/lZcJxzM
e9Lp64+VxwclnSAyA6bI44wHVvjuBJ8Sf483YSLxSD1GCddIrj6VHr5eQP7nIUqd
4aZp2dio5bjUumiNHBH1X3zF3ITFrm/clGtGxRKkie3P/VefZKoUHe82cyAbFYGl
OKttlVrBviGiUgLZLHfQtl/AGiF21tmu4LJbr7ITW4xeGYwX6XfmbjjQLmCqQv6c
ppmI2aCWt8Ez2MLkg6AkDt+G2lI6uXqnkINHaHmpAOi9q5PLVQZm65utPnNICr5j
467gyQs0olWksoUCDHmlLmkyAu222c1UJ7rgp9hxo8986SyPBwDo3Y+swZ+tmB6I
LJ593DXNqy2JoD31PvRp3EBk6m4TIk2GsrSxGB4aJ68DH3w5wwxCAFVzY7eIx9WS
sQZkc2WmOUpWS4/4Ic3Kh+GRqIRLnuqSTVNneVAiJBPmwunf1HT/QDSGo4QtCnaN
OpHTOwsnAEtPtWoW5t+ai+AZPBOMtG6okD3ymqoFm0T0LlmAsVxItfBsy1lG8bLs
Tay0yRfPDsMas+bOO8q8uJqg2VvY39170qya/DFsTbOmoKafWNgwPix+iXddyBoZ
KdMNwrc2LsuYdfEK/uWfnKXeYQJZWH4Er7FBCOvI6DQ289c0gKFFERUmMyvuZFwZ
prwNFbRuj4w/VaKiBMXxJs2rS4Fk/tyk23YlJ0YMSGAt8DMAEED9eRSULcCUO1V5
58s/XLI2YHl2/VQp1Y3bByxw4QAIhpyO3CyMhf/ODYhDNJ9E6fGZAb1M6M69uss1
0ZKSCOeTQL7ixJf0Ls76GOXXbQF3CU+qQst+8dj0QdjtbN30HfGSI11gzCCdH0Wi
yWOwDn/eqnjMR75rX2qKwidZfpZKQIBWZKFER7kf8LMzWNrSO+0LwXhjUqzKOfwA
VIO1iaadI2ULarpuLaeH5xLY471+qKv2CA7lcLlZV1/XDIhRAZYPvmjqh5rrd6M8
s3XUB/wPbuAotwAfMssa9ve59Xn5FgVY6lgwjXNYMN1ZdbVjDEOnbIuLLtavay1I
5MR3Z907zULKxZiWRmlA0oBizV30w3az/J5cvnyHUMg4SS96AFnE2bX/Ihf1eEsr
lnxcRShA+rrCowPFDAoUcNW4yOWhlt+ZGcAi4ifeRhIKH5g4O3bWiGR3dsf13JZr
GvbCQDvjrfJlpL7SapSXdQvUkk2c0gIxaB8JnmIylnImh5N0h6IH9KaPAz0TlyIn
37uWa8Qq+1KsqDQ/R11BgWxaSwSSlCSP4+22sztgrsY9NWp5UJPxc+uOLQFNecOF
FqZU1fTkqjbl09e8Y73hJy5Ss8EtC1MApuuB5CAgnYRlYXFWPAt2sm+li7a/Lu5Q
57cdLPRhjW5IUw805KhAFYDzZoQCq8zXuG0R4AUWHkuUMMs7+dxCoPh4X63vb73R
nFes3CnFwOsKVRGm6ody397NNrYWK1AfqcrjK5f7RragdzlYycJaisjWZNvPMupD
JzITQP5kV5/uzR1yWdDkPoVyiynQwxJrmhh35u3HkaTko/bquCYj/3vNe5XwuWbb
udTxDOYPeI1F33tNiCroXp2Bv4Q3eJZ3ZFKCrZs7lLa8x4lVk/hJBVsoEfBZpFFr
MkQsCnocogajHqlZYH+/J4HGmbdS/ij85pIle4XAfeYjFE8XEzcBUsGU0p4IToa4
Ooz+QH9N2njMRnNmxruer1zAvzdY+3bwjJm0L6IRkrzlcvpTB8PDs6D3RypAGl61
JuteiuexTL1IUTPmo36Rxy7Qax1kKoujDATvcicRWoPMWqVTSamg8iQsGKO5Iv7X
zZf/dRBX+E0lJRF/l0LIxjYeQfJPe8d006vbPamkm8u2oOKz8gIUstLJlJq9ooO/
xF8tibjq5yR9dHtgR8zrLpmYzmbxihI2x5p5/nEl0g8YTTysEBhnsAeZIAU44Ek+
OjMCsJl7jEEki4oqFwM2wW/1mQOWef1gnyhlLWy1LGgGbB59cBag129h08ZO+T6I
GYKPESqanMQ4FNTqvBM7LKbxGyEtQUHHXD/UXwq6z4z4oPMOUeTZmE3+lECguF8q
Tx7HpLD4DkOkagaYCHGwDa1aryuD6g5tdIG94PI06XmpRQY8phESsX+NdjtLwkv0
n02etbvqxnG1WvmHwewwlKOnyYHaWJqGLzECDc8gfTwTrbMuRAYLJx7Y45YGR/kK
5lW6HiPyKVQw7kW6msf9/ih96VU9oXL1Y+JeiY6S7Aq2nsNqLzJYi1rL2Xju5Nww
qmKICyepCVq6Lm7XHybPTU8BdxpAlHvu5ipCwSYe/MKiENe40fUPR9IMzs0RLO+q
KFuKtXPhH8t+Zm9lgpB9HOu2fUZ197Pkx0Y+RspiF5/uEcbLfix571y04ljHkT0M
ZkV/NrvCma8PGMVgMoOimQnh1dCKuPrWOrN62OicNyL743gv0aoQYs1PvdodbqOa
pIO8yBT4YRuU3dPkdemriSKprWUfHKHO3yNq1L1uQnugFIqEKEf/BY4Ex+/MyHov
EcvBMq3vgmsnaCoJ4TjR5oBdiB42PSeN/t/xy+Rftq8sfO4U1h6GXHwNeq9bDiXK
arkwo6nBBE5cH/xGmFCRyetBDoYT6nj3M4+wG9GHFORT7RD+Ng794LTHYOOAWKan
PbujwfVr8KVuo2ongKKW/7/WYlw5SYbAOJSJVKP9Fq0evWRe86GJ7CbhcEGSUFBb
IDKFTTuPlVlLjYsm/e98S3ELj6tI/bAS1K3qRRXghW0pMQpmBm1O58WLQvvvpiTV
o3//LTqKY1tKwe5SF3It4L5qu38O2TPa1hlHLXQcfMqJflNrYkmVR0WCkZsHiwne
MKQWaflc4Rpfi67LLfFo8CsNz+XXbGgTtA4yf7YO3Fwk/Pz2KeAV6fByryNAoKmt
sD23RQgDLzLAM+6OCV4Rw0Cx750vrR2EyvWjBXrXhjvKH5tIYt19JQNnmIXEuRva
716dcWncHiGspi89kIQeDYc41bq+8K7DdAG13iEskbHZjVcrIYIgUER+KFmmZwvn
7V6llrx44EI3APg49TO/PPvvyYpYRtrDRTBrl60lfNZXniaSeVcONDSktACvNNVA
wxQdsmp44g8SCHm+UhHCHdx8M0SDaEupDxOQv7ViH7ZRnfVaVgh9cJisHAuKnZer
qoHcF8OqP5+vOJhSC3qRoiHcMEbKCLHEvgOXb/2+7MKmF92M8n7WeoRtE8kKof28
MVuDuSUT/UMrAAevX0PKV9eZcYVv2QEWUPN7KelqTAsbobfkS7I7hX2ydqo+Ca79
RHH0Eo2lXyceYWIBM5nls3vQlO0JjDuymGlMxMtlAAGq9E2AsmuOl9ZIH4KB5rvi
Trli1cf9L1v/BwfWA8Ajw3j2uXbzKjBMKUR0V9vH/kZb1WClr7F4MOFElYThycDB
lHlH/LfOCToza6kZewXe8GGBXLxOjj1DoIfNoknTyIeSWsuJBVVQjlyRYXwq+/zI
pC/flFU1mV0iDGzIzooHjlczqar7m0Aq875OBhn7NV4n1vR5QvzYV5v3fsJQbaTt
ZI9TS6mg88ek9KDKKZ0ujRZyjw4/fKNwWp81TcvyP59zI4oARIii0YLe6GSXZgvm
mN5dUQFeqhf6nMVjYvqXPlzPeKvI48wQ9I1ZoBPaLtU/8pEJnDUGoIoz8aTTUvRJ
wYhvj28zsYrM0TrTwTmut4KvaJ6aEyQoBw017F88zakDtntgWLmb9wYw+7/B3pus
mANZUZRfn+QnULcUTXgexXs+VwzmkkfKdyRbfpfbl7OpoH6WvFg/QZJyGbiOlJvS
VJLj2iu2nYjOhr0WAq4+MLZolVRvyVLNGpmUQQb0rrH83Z0Hk77b9vll9LUucPSv
3130kzkYKZGRDPumJ+DjfJhSSuSO7D98YPT0NCbepODoh59CSxlpB+YFFgTs9rlU
d3Sor0jVHlUwTnz3MWoGtEdbFHatJrJuhi4PeSwOBKaWPwAfqgb0/NNhYe2l5WGS
T2Mk81tYpn7nKnJeLiw9C9ooGedID7rK4SZsyZpdgS+6xnZ9CwBlRFmR0UONWP3y
bT9BoAp7YVGJU4xU9xJw7Uc10WEMxQ3RbGJpfnS7OBntMRXriIP2GE4NgXzNfH/x
c9KptfHDuPybqXjDKdZeQz1vYpH1MLIVgSb1DxZD2wVU/qfN3VTXf8MVtD0ZhO/S
bpxejS59KU7jwgdEY7ogCxsAohivYxwrgKop+j6G1Op4NFE/0ifbHkUy9Ikt9iNt
oVaR0fAT9SInrQQwYDT5z2y9h4d++LaAELnql255BCM++tiOaZnRjrbLWqei7KQV
/NixxSj/go5bYGshnOIYWp/uH/KUKeH1P1wvCB63NhgsXZxac+MclkPM06ucTW+U
d/C0MtQtCiCmBIvabOQMtWPP3hLHonBXzV6+RAztoxhOSVD2MJQVn0Aa08QJ+IGi
XnWJlQtTVLD7MXKHUdsUIoksy9DrbEnTFelA7lGRXf3lh8S4rXAo4+1xO2KMHykg
8nfjtr43VJHdIS5W8g3r1wkeIKGtDQKHzEKWkJThG32f2266pIIeApcHq0n0ePXV
tecoVsZZySBp+pOHfFA2e+f3C3fXEcDg1GY+VYUeAaNZe7gaGeZ5jE/iAZBKcxl3
/3/sxpiUmAC7p0xXQOk9pPZkIKVZuIqV6JLynoIGpryu0Mlp0uliwm4IpBZ5kQS1
q8DDdHTiWFwEDHzXI2gDhMUZpkebQLSmq3ydUe+zSVcLDc9b+iirZWVEySGtVvj7
y2R+bknbO20W2bv9HYzGR23KXYf5JSP5ylbA0e45pbt3iC9zOeokls8I9TQ7Icg7
tp5xFa65Be6OAN7gqLG0dCm+OfbJt3RPaLR8cRSMo+VkUdluEXPsqVWbhdKifps6
rCd5SdwrlbJs00veNF4JFYTFIckJTps24GauQP0mA86UV/LQ62Qmz3s3ipYW5HJy
3JXRsuoYIcvWk6p7wa2Qqz9eX5gFMTJC31U3c2n5hU8bBHcrxeTgXhqqfBApVKJB
aJn09gjSvHnyineSAAnKmjsbqmkzjdQ4EvjG7pRChwRvPlnggUfvbIU0YKfjEC2V
dH7iFXxOEtoH+SWVmAVxDoubqekqIq1ISRKZHViJ9Spay6Ab+0zdDME73MtLoMNp
6JUSXjfMajieyiOsFyn0dE+WxlAfkBhGu6Byzs9WGVI6RT0hexl1F/VQzKxYPoxV
K+1B5kbvOG/Do3gQWy7yxzRvk1YnS5Lly17sdLkm1Ban6pxFdWkv3cQ7cbb8rkye
HwZUC5heXK/CgG1IJi0jJIHl47kUny/q7mTKb1w4NmhQQFyj00NnmRWhdF45DyJH
rf20Z9CzKFenyaB/fmeMF43s/Z5+c2BNiVyYPm9E1QRG1KjulGsbhE5ft8bUeg7T
2YxziHJ0wxBoYz4Us6sxu9vR7xPqVp539yJE2BYzFgeMg3950S4AvURoEtK+F+hO
TusFKLC2EKo1Ut/C7Jl5qaeioxce5vfzE1zhJXhHXozqHRIYC9UdW23XLINNhAt/
MA22i9gQTrFZwwWdkAbHdi1BhaR9WU8afb6tQyFE1+TYj21fszB1RMRb3JxnkI81
8G2VnxRtt16wuOY8nkfUy443HPivBeQ9IcPU9o+woy0TrHaIL7gb8KherWraeT8l
1WxuqFSQwkWiDp4zLFveNYhjXwTsBVmaX88zitQ2FSCz4Ohj4GjDcb/yXpeCyQYp
FUW3W+K92jBVUGCIAk3wT5+8kiUqIxf5cZwuLzEOAgWAEmim8eOy7fFE95exIEBP
6xLH8TJFyWJHDfmB/xt1sUpz8N5CE7w79HstkkdSZRLNBFR2hLLscBWfdRAmoIyH
RH7RbZQsPejJwpcxh52Qgknx5TMkR83gaz6dX6bWUNtZ+FO19z3ay2vnk+fMIq4c
PVfJy6GDOq+YmyEDcFaGw/9ViR/0CBENuW4nXp41LVq/HSnTAmP6ViSxKcisKQIU
WGSnkX3ImjhZBuUXdflIjD3pCg0ptR6RJffw/GkG96f8/veXCVOPG6fb3wsvpvRh
WB5EsrHzvM+bXSloczO3JpwoLQc2T5VmbqP5UhfnffUDpFEOM1JG6Hm1dh6/DuVl
jsnZzBYylZTkyw5sDVmBr+yfalTVx3Tx9R59B/P5mNHIagxiF6ixaUiFLGIbHX7B
2dbrZ3q4HK1+Zy5tWtVzGPBotCoAKIN6vLVZZkx0L483MnQJ/sopyE7hiXUwc8YN
0QoQ1Aq6gWnBgZnzwlcs272gAUjKO6p0+EMcu6hdU3Jhsk6ZvqQNQ9nWQCGOda70
WrBMR9mQc+K4HF5InZPCPOgjdIVtyHFKQ+SHVDEWf2URO66B0eObL/vEoFKypmOd
rKkgMFO9KlwAgC73dE/TgvcBNLsKsWSI9sk4VYb7fv3F9N+BtgxANf0/sTPlq3x7
t+6pIzjVKegWNaiaRzDziEqlzQaof9h/gZzzvnnHPSW5byRka94DsSAGovhU7Pyq
mecykW0rfon2ZycNfyp3kCQfPNncE5m+2CA/pnEPYLZMITBlAXdCsoqgQd70bAJo
uClbIwLmtO2NGX7GRfs4DO3b/VK2QiquzRondwhbxwUYV5wwWQ8JRp/fW0S2gQuF
lxyhlOe4FcebC1s4BRUTI+xgS9ba5ziKCZOug4gZ3JmaHNm1XiFMIa7BLTpdI9Hi
pOv1BybF4mpyjTat6LcBKeR6UDcKt1v7rh/6Kudk5UcJT1CRVKxCSCXCxlpxiBjj
enClAkxa92satrvauEIPULJQ0837nP0XdwgKfiYFHoVLdhac4HyEWjXXMIqfUkml
UHTS3hC+pVFUSd/bT+3OY+f55lZgyZOZ7jEYQjn/qIXuZkE09b2bCvn02teZ3zVn
BzzrZmKdsYQ4iBxwfljlrdYafEMfAXZ1shWmUsMprEd6AX0SI28R78FDn8NVS2YF
wUFUkbnZeAXitLQAj2cu2NWuPqKvWOiX74mXtxP+HVCYEdANBHiIHnv1XQUKyS2O
50c/vv29wT0WbPvYHsSwkujtmyGGCRgBXishUY6ZtvjB/p6fzXULQJA+1wpDI22/
BfmczgZNVTBLKLP6fhry6kFflyU8ZYuIYtcodLxiC/ohaHTXZoXHb9NbO6qTdNM+
ZznvnRQlZJxas+8DJB5+FzOa0umWI5yexBhQ1mlokknKESw5X0ZrLtKU9axBr/Sh
V4fY7FB4ESwIv1Dw/TY581egzyCWch4kbhjfVPtnk6pDNtLU3uJRNCJLymJLCHM8
aID4iJEG7aazEs+RiehtFReuYttJZ+IJJnDWgBnYtl8/W3s0uuxpa7I/KDQGQWcz
sinLcxwGKub5AkkfUUg4Q3IB2mCgtuvPrI8QcAJ4L9ip0lecVATdnKUnuHvZVVuV
N6bf14kOFIFKp/6zdDkZhtW11A2lv4ARTfaKhxVTMCLr1+QPjLTnU1MvGAWIOsc6
KnbC9rQx+DdwsDAuXehNK1uqOY4ygACBT5K5WoEnNCKpn/udxy1vVmgLCFL/6ZX+
4Ad0Am+ENjC+Zt8Ouz/ia+wJx8Nmukcd754qLG7lBWXU/BkzgywrgIZOftGRJ6cT
rf1GxOvc/cBUunmHQmzplfUTS+RX00Vd9zesduUDNPL4DWon8Y9oBuMkSYS7bun9
iSGrcOy6W12PRF2RaPdDwMQSH8ij5mdzeYOh+FgQwrhytsgffEsinbS56vGRhQZS
OChVqH3TdL9KXBTtyyf6whzLWMqMVji3BrjZQuXikc72zCS7uXpYr0Z1pr6iD2KH
G+bL7DNaJTl3ekKnhrYxAfQ/uuwYCn6AG3znMYLsqCV1qzIy1zPEaAaJ7iPAt2MX
tLauR+6tZpAL9UVrGD7oZQOH6xkxtFVibF3f8pGm2D0OPxaedTVrEXd2MwzLOHKi
GmLSkOiDx9ccVcqL9TMi6zdq3KSdxOormaDLp+NfRUKmHa2IrfzfIFsc4meFWt0K
twblN0jHZjBgtAeZPRSqdjMUME+Cq6NFdpnm2T5O2u0vFGz7NzWcjtdECcxkeJrI
NGdhiFdQZ1/NMlwYO4FqJVbFwl2g4xCWanZMF6gYs5Uotr/hB2bA2jR6qZ5NkYa/
/r37GxnKSeqTYuUgeqhRRZLW/WDvhAgB8vh55KHOmspQwojCmTAsfFv6MTh5R9OK
1zz5E7ZAsmCAra7CbWzrZnaBYHKafh0cINpl7y+qkU4ri+v4zlwt4XgQw+xULolR
VkfRalDQwmKYs5VzrZPMI/LuMe09f1gxGbAsdghnfvlVkz+WcjbEJkHBQD+yzKtk
oG9GH5rWdVRvU5zTzbCeVV29wZ5iD8B0MKDt5/p+S1FjkwUvMpVlbS8ow9RGl1Z9
lhZitQco5BbE6J/mepMu/EPBkDzmOPr57TFsXJ8PH223rKYBlLdwjQziEOJ4QyK0
6KImH/NZoXVlf+daPNCHS4FBqA72xdz1sZDx3VqCFQwqZWKYCdrMIS51xg8/Uv0W
U8zcr8VF4vE9DnNOG2mIs+me2CpPqfW+TT+Lj791Nb4ZFkzfACoLB9OqZeJmqbvW
URw/rexnRK0CpEEOhBhI12NjwuYBYmLQEaKEvw2+9gG4cSe5fRnm4WBKyIBQWmu/
1EMfdTbPcd2ym0Dt0oLst8pprpLpbRLJ0sdGlR2WqOta0jlYnfNCM93g0XvetrxV
JJX+xJczjCoUrDjV42fJprs7ih8qnClTERHUIvY6Sx6DhNBATnklH7VBLKcpc32p
p9hLpZwJxwv/74G452TW/aISMn9M0TPOEjrI3LFS1UjEuH+d1ysB6LkteKVqhnVk
7Zt7HWsS1m2YY2tpZ+5tJ1+B89FcLZI8UEgwPty8C7vlUjPnzlXiJkJxkfO1GDaW
QVO7A/xRPwSNs8x/v0f9KItjijelM2m8uq07ErkkUKclAcF0a3ht3RMqhfYrEHsT
JCasRFtEvtKEMxTi56EgHcB3FEmXvcvjrPJMYyhkEUaSzvJqmbmsxCSgLORup+eJ
dWe1XDLSudQwUlceJnf8a02eUq/r36ItFlw+VpBLva1cjmL1nMAGhXpFNJ+puSHk
2yYTpknnHnqGS3pTERXP6kNi6Fv5ZE6/QFwS1gW7kynhs/HGpbyaLZYT8OCvW9iv
NagYfYFOEZJO8Y4S05iTdJDxvn3DqpNxGI3AJG4YpnUwp4oii1Zw80rvM+4QgVyh
ivYcHKRDMJ+SyI74SHGtfmBZOJ5TTkto9K89SEppW5OIWlb4xsWS6olFaY2Xh563
WSWEwmbP/H4+kW2XgGb5gUafNSSEl23iJTy+15ziS5QOJwwnYI30VaunsLS/xa1f
FieE91+ytZCigyY8pM5EZybQJ32NV5DtC3uFAa1xpIsXi3IsDjkrt3WxqhiK360A
DqVHSrV3S8lpJ97Rze7ISWHKXTJgWS3HiUYmoA5VhD1nA2kxQgW173OVeONG7Mic
Qh+67hfMoltnYUb2PEjhbbffiZ+hCyj8tYQyGsEw0PfzC4kbuPTlm8zNGr8yUpws
utvrppAVrYloHamGPcH9a/Mb+dQIO0af242BZSgLC5B5Qi8kgoAo+zNxVRXSap1w
zoCk9EqT4LKdEu+PDLl82JojDvWx4h/FrTraoyA7iT6/56A0mieryGthAYYOa4bx
4kzs14MfFT62ocLzih7We397dt1dLVcXQzxrCOsqarenTjlukCIC0iquZ/VAArkG
epZbrnjx31XfFvLBWKk35UzGx+qoyFrp1d9XHiUhIH79YboFRhuGKIlK+AR1h23C
+ZDuC2LEBeLDY6sAwAfD1T4OFdhLnxh2A1jyZ4JUsNbNqY2Q72PgAxjPHJO2PWOz
uvRYMdf7eneazffHYaL5VscP+YM52oX3+ukD3WaBxf/3koRyLi3B3WzUEIDWN/K/
xBBpU7mtmCzO4zkgZnWpfCfW3nWVyC+qqso0VJ9hZ2cucibjvY3tExpFy4dky+Kz
VfRg9b2ka53jWajlPBHRFezORZdoljTJWMdbp4GHOrmks28EQWVY7Q5qEDbr8ixZ
vBMM1uildhN2ybHQ9WK69Toqyz2t4eZJEM2rHZQ+Jule9C/5SQXmfLfBCT4bfgxv
TyzRr0T3Z2pxVwCbJNLhQsf44M3uUeK127obfhnJsnxgz3hbLwCEzki6v7SQcJIv
8TO7oolmjQ+2EiDC1O+SNUiBwgQXruDELnnFMRy5uk+Nh+KQorvkx5c9gYpVwtoe
8Q+1vu/fMBWzisgVgtxpIk8hI3nwm7TjgyzjHePHFSLkpfUhe5wP2uA4dXfENcU7
Ot/bJPo/dBzDtDJezDdWxIPTUJGUVoUCHnZ1mqILbftiir+qHIcok2koc7e9ctlt
jtgYk7X36uWufPlTk67pY1OovV61pHFWCKNAWg038UjulGWoEou7auMJS03MaNGS
N+oZ2dob8OyVbQFqZ+mt7cGwb/DrrRnLCDln5a7KS38WFx6ERKy+s+x8+WHiyWbW
FbHx9M/2oYh7iEDmJj5gAuErNZgtE1amh8S/v1FzolHRo4dYMBUhTb4NVXv0pDZ1
OssDhlX9oYl6GR9MoqMYdeJbPCjmnPgpKIFwMUnyx/wAYuIQWtiCCZ2xvaVTeD8/
URMNZ5tCglxdkSyK7SIIZniNa/rjBmu3UF2DFjSJkVN8S5bSOIIqfITA6lUsc9Fz
T78rlF8IhxFD8LrUCRmsaKxzeUfp/b5oyM99/+cRTq8EhScZ5DLTYB9MCNXB43kV
ezQle/IYG/9xTyulnr83AxXcA5QXhlPT8irwj7RQ/IOtrwSaE9ZeuY6r/Y7c57Hg
LYOrA4PFjGlbDjWbtw/gPl68BSWmIHyHiUnnffNbmAgS1a2HAY5xtm+BvQiV9OWn
SWB7mQUkzfzGv5KAqtUd2NP2q5H5DudcIi6I3Uf3dzbb+1VumQ5HeWwcbOQBwMq9
R/C0GmZ6/nwF8kGcYyfvttQNdmB8P416caOYfeRQ7RlZvgyMsD/injxsSPPJY+wL
hpKAcDs7ZTcBGo8FT5rEC590z31benfKmnZHDrZVvz//ZMu5X8VDwKHz7Uy1cVQ2
kXUb9SYHamPTZe7dNoUPS5uXqSS6ZpDv1Yh7U8m8DThWbcfyd+W4oL3v2++iEYv6
RZLVFkFswqZIBwK2sAJhEKh5j4mdBLhkZqlZRxm4HDbfaRyEzqlzYJ8lZ2h1y/3g
ZiRakIHei//zRv0/tX5DaBpr+fCgm2UhAKbAxJVNHX1OTN8o08jikmUbYV0KtHxm
e9Vov4IJ2FhDvtDg9GA8841hGT/R7CZBQ/wuQRl70myBJyQJuQUnfIidoPIhFceM
Q+5WVx/jULURejo16RBVGt5BvGT4PLmImtOGWkaQCkxu9WgbZcFtoCwizkHmXLwU
rW95Ea/Z4uwgc0XnSAv0h4GUTIkNLnNLnCs88Sw7ZNMrgggoDyn0GrLbZ3/tsuYb
EY4rW2AnSKIu+bCXFaIpELyZICHON8cVxHOp8swYcvUcfjdBQvrImhoascEb3RQg
2Aht4Rh4Dp+QIdF27DU8C+C2XgqQjUYxwqGoK5HS43yzqNdJKwCkGKHgY/bZwlK7
gXAWPHKLAUmik9Hv5KNksdtGKoR5oaBbYVykWDzG9rJAjmXQfI0QrEQLntMnRcc0
BSu8GDhOLceWYBwJpGHm28gqDSKl1sXqLaVS3lKbf/xenAk0GYiQFIzW8YLUzidb
TDg6zKyj65eLBtxaapOu3qMyo1E/elp1y4l45Cg7xB4NnxTh5lo004AjpM9InB28
10GE6hUBtW8hHXo39LtsV3QnKPPEzDwaqs7wp97XdAsyWuC0hoArHbgICWXLb2Q2
RSufQh/wi833Op9vmItgaBsQa2YhY6Ph0N56UBWsoJpCHsL7Poy93yx3XdtlP/M0
cJKwjwG/o8J6YR5+62t5wvHYu557H/57nsoeloyMPm9EjrgNiFVtE36rO6COZeU/
lrUGeLbV/f8StGSfQRRRmNd7GkKUXS5rfL3cRGaBxWVJ9NyriYZkbrmyjUCgZVk5
kEbGb3psauQ6IIvWJ4opOBgDWIwoQWOj2QFCm6C+iO4DlhhaOSkFcdxPK08miM4T
fFDd32CWDc0ZkXG3vqBSlR4xuKpQLbJPnia2QK+cj8fTRSP/V1WHIhQHCsM3K33F
DO4QAWdrCIJf6t7vzCvitoXfO1Zh06ULdhc0jhuuAb1zFLJZSQeUBjTriJf7AHCw
raGtPTmitCxNadm/bK9O+93NMO+JhC4U3+hwbBJyzBYuSV0tWZW4xrM0J17kFpPG
bYa7augHNFuZr8YBnBRnftQY/FSZ3WM0DtSxW1OpENZTkVuhbTGadKhAyx2eODSE
gYCNlRzavonQbZVeBSKqw7vNZzW7T3ogckT94tzvUioUB5w6P+c/WVb9WnXia6M9
jqNUmJxPy9lXqcM3bP41CyVd0GQLaK7TwEV1IfEsw8MVvoSHsrgWS5P6JZoSY6e9
t8RilWjWweiqj/OuYJ/kpixZ8u0FqHrfLU+vLY+dxZpJlL3090Oswxc16137Riqe
52Zu8Prb8XSeAQVQM/h1MdKV7pA26jlNP/7UNK/bQjR7RWGeZAU6kLJ9/g3u6Xx5
PqTJHWknFsI8aSYLYktsuFD15VJM92cImrLojfrFTdIcieed0Ki8o4nFBRE/6omf
NuHyUT42M3Uvek2rn2Fg/MSy960gKyA0axezBfi4F6JtoRf86py2IohqU6IpYgeb
GuPllGWmLH5oLYAxOaCzsGQjetP6n6rNjnliBEJXOWusJpXjBsU1RmDcUJi18VJu
pQ+WCxHYAqCzB+ygSkSYTb9by10SzCT4HCpxqbeVVHDE/gxhRMF5nlZs4AAfbLRV
tW+MjTB7TrRf6s77xlIhcIUSvsMiEI41EaVDjomnff8GhcnttY5tyvIKH4sHnkTa
XxQLmk0rZic5m8dtDfcw3vVBEDnB3krj1JHTl6VaHLRKDRVMKFaZC5xWLI3BggWs
hHLBBXg23BzWAi/mnlIrc81bdgf10+UI99DISjjkRGAPrgsn1FHw3MK73H8UdoRQ
BxgmbZEe0cJo2G73nzKRvewEmST0knU0MNFED3j77T3wOwFu9hgBA7V/LNgcSLy1
8h+8qJ43XKqs8+XgTiRLtlxcrZRd2SCAR+7fWclntzVI1yOGwk1BryduLIMhNaqB
NkUhUlgD5Zai0G+Ix629bplKUA1G7HDUKWqJpf2QbJuBFP+hOUCGFV5sXE+wbpl2
BWjf9capXEnQTVMWAGDZS+Ncq6pjuQFgsnXAvrBkI44AsiQ0RrqRGRXG2GgetNEm
yhXFB/ihDmothXX4ApRDhZKk5oHx92aBwz6axzDeMB0vov1Dzn0CJJEh3g7/3BIi
9SM3T1nTJjkKe3jOkfJk8Z0VcBA9gA/y1KIgTc91MtAV+zLGWC+oLs78OvFtI1Gy
6rpvK3FnKIEb/IXBu7CB6tFtkwiYtdW2RbBnc1PlWBJRKBmT0/3rufBHnuLnamic
CIgqIF3pzeH36OJoDmt9oarbXHua3y0+zX02YYfdtU23gtTUjm8PZNRIKO+pvIYB
v1zoa9xDVCfTxiQyTrFNcOaqB8RlchrVuqCeFMW6IFnvgpKEIwukp4CAhd6XddfM
t2cIzeYkgyLx1cMIJILb6Jswg8p5f1UfddxKRi+gsWjrKfRkDzQHvFD+R8mRmZOp
twwdPXoKr4UoDGT5jChvsmITrX5bWQ8c4LLgwD+v4BWfn+fnrcHm3LacNImt0WIa
YVlpByTNOwMTVOgNh+iQGcq+X7CiRYb336qsZMlHC8CHHP1ehzra7yLeUrvGL65G
wBsehqJGEpIxKWuNM+O2LBxxLW/ujxFiUAWHK3/wN0R23A5ocEBB9mx75VJDvGnD
IDNJ3+j9x9P88wnIVyPs1vVU7AQ2w5fZm78JkDeYPOrlnHc8chjajTuqzH/OW8x7
NcWbqqeonV+orFeBorDa4+hE6RO3FpGjyiFPTGzbM3cbaAUysuAMLERxX9ppzIh6
Fquze5FFsuJ12VvqHd71qibEpkvJwvfukvoDTonJIqoV1wtdPkrb75cHkVoPZxde
mXTgCTCzgMRdJGuMs/bYqc796d+8l5RvbEayOeXKoVPxE4WGtu4zsUesu8Ui38AS
yRLDGSrH5Nao3q1tssWY4lGQFW7YrFc+OIR6TazCEShjUB9oo9PlU1tUJSWF7RSP
o/PuPhwdjdlWvbEu9nkUYOh4OmRgx/peX9UTKtjU3s7H+6FfSA069azxtByRC/zh
wQ3HZzX7MVGbfHktLP89FL+zSmMCmJOJX+b6mkUnYJnpiQ33juvmuU53ZxKismz+
4EUPlitB+ToNvCDW3X1RNXzkMjQgO3l6Kr2yg1uArTPeQYH+4eSPCpaph8ty410K
2ItnNo6rvgXVHdToMfG5IvTBeUPuli87VQLA1kgBCNXD3T1iaz5BBl00SvE447Lb
8r6PYHB1npIquv4L+GdjKl1bWx8HRtB/6dRNp85E8pF/EawxIaM/voKO1jacPjZZ
fdhObVyJHOwuuiM00SO1ShNsNvhaXminEpo5+oZm02PX4eUXXPU6DeJbyxwdFBUh
lP5/6c2IXZZY4/ELQZSbLEaVFJKQGbVT16vPpYep3wBiZGdq0G/yESJr86KXhy2M
lHx/ZbQLsnV2XcDXNFDy4zbFkvHQqcmUPgm/sXc5NCsw4SdTgDG+umX7hMxZkBeu
fPMikAAbX9L9oVKPnpD+srUOupQ+QUTx+oBa8oREIB9snMMrUmtJD39FifhymlK9
gKlgor+/0ZBoXHYu9DGmLr9Y5vrkBXWKIpYPGW/V9SfhISAaFjIrw609v0yapJlC
tiS6+Uvhc0rvrMnPJEFIPCPOc51P+9uNv6W2WVKY4L4YvWPliHxJqzu8TB7rtv62
2R5ycrHIH32uqR8atj9FaA6jVM7IceUNzKxZy8eWFOMYKA6Cg4eFzujfquD8bEz4
08+L5TU8j3aqg/0XpZhPfof/KNf085lmofXwHC5NdQ4fMKGyR1+ZrnrQzdyBDa9L
7uGMne/8iCZQXbExEUNVFzGZk1XKM7W1orq805vQw6TTieKsVwSLE4cMHffz3AUE
7Iwzntu/hyFwNrR6meO8Y/JbW9PTXGFpx6hZSKT4hBuvWQWkk1NzKIIYD58/RryK
otr2FBCm91aUo/Dd6vWDUe01PBlVMHOO0ZqZ5iwfXI7+fguG21rMbSxyekT6DhY0
udvrUYwzdyQCZbhOXYPz7HJqdRzgMUPctK+nkQLShmg8nS0c/MXUVekPEW+LdpW0
iozsJkfnZ8awvim39stJrX43cvqbpW2+jW+Te55ad9ElgV0Q/HTAh4LG+vRXRYPE
7RkDF2aaejUpeJnyT18q0sq3CtSkQSLcZYifdOyw7sFa7xD1OpMV+yzCJDKCVAkT
FkguFjbFA+OOCKofNf4vjbcUiaX1n//HqodTtcnIJ6GI/u9Kpx83wXHJChjQKVTz
cpn2d449ne5QHOncT/3CI7olVwkOopqdhjrNAAx+WraKJyOSdp7t+toUrL/bY3Y3
8JnHLzUdBtBYvFNTvsaMr25g+DQ3Fa5nYPCCjP1BzRlOdoHmfJ53hUVXprFhcl/D
eAVsnCr199gBQsn0cd/W2P1p0aQjixI0/9yJG7F9GrfRB6FNqIf09WMrZ1e4H5ga
XVxzOyT2qNp10Cc9vfINualiMqE3ZvbTaGY/rxhv1BJG4wva3OoCGgMTfIJ3ZBJz
i7eUqCr3DmliN8/VuTsqvpT/BzOYh61o5nnRloMwGboNfxZaX6/dbCwXIhoWt6vW
mg6jVxXC5WG6kdXcq9xlUvEd1On2jF4jlkptdCh9CebPoIDxKiQGHTJKBbJHKaSF
WPX2IQA/P5TJBXWkMrsXxJFt3KEshF/WKUCOjXTASIdvGQVFGZHMx0T8IQbVx7+6
R9f+GjGPRCST1Ib/G7pHNT0Vc9HanwIuYje5Mux9I24WGsIStjZ0vPCpnZ8pwY9h
GK6iJUCqCE4/cLPqbHaka2TiYvK1qsjOzTYPGxiRHfVm4hqwMteApow9wpoC3iAT
kb9ewlCUhUPJDhjaXnNXRtVJ+xTvW87ejnO8UdnrKhmvjbGyHpmprpA4yLt6X8Pd
6uMk7p9bXmyZyiViA4+Cd/e000ZmIJuL4wepoxsJ3AA8bZhdZRRI+uviVvr2tSjg
Q6luaVJayelivfYPbaDDQMKd1qMlPqqIRoOoVy2Nzicgat1Mkz8W43wErEW1QfsI
aSB7HZ4KFLwjVF03/p89Xfp6VpUh5n63w9qC5dK+ce2qMt5s1Ys9jWJ5RdcZmRSp
AiMi0sOXuMQyYwWxYxsDk1xjY2PN06itHi8J5KIZK79C4aTuHYGb8UelDGk0Hm5X
4WXoR++FptGpiMyyXF+mNyb3TXG9srI9Rhv2z2gJdhLx7CtaoHRZOMUhaVaBydLR
s0A+frYwqblY0H4VcHMb8XIxdud8hccly22P3zEm5hWkoUkOCgeJOAmzDsrwq3G7
USTtGhzstbAo9RnuuH0UmKPimAwMFkWOcu+5X0zRRiiMxWtpkrBTB1v2qCN4d2BQ
76taWvIjPCmD7bY0CcYUag1aR0c1LGdEXS99ruMJWHrje8DPuA1iLzTZi0MTsyYI
cUuxIpUtYbZ75pofN9cqzKGx0T6rLjh2hDcs0OW/TrPpG6mSMrNuOXpzGpgGGA51
rm7ZG3bon+ySJ6rK14MTbDYtUG6WNipDj7k4ffnuWeYe4XqqTpnQADLyPO43izLj
EfBqHfTV8UmfVdSSl2PPG/BswBnT0kvEjAEpyDQfaTOdL/NDI+Wc/e3dlIImJjRQ
TUqotk7/RA7G6ndH2Bv35vNRlHtXVkx/nyhxkHxN8aycjkFZfcQF/3WmfQtdrH/S
BP84Dd4rFDYhHbD5lP51M9ZOBTjdyCIEI7YeQS1k1AQ2DwvOU31umt3LVGPR8EX9
MqTpfAWl1pCCG6zhlWzlW8vIP2jvjJukIFW26NxvOZ5R9f8twOKKZ1FBu2Z6SrXM
/ORsBPw7RGmeycifUopKeTXfH0Eg1IBi948wcUy6GiC++TFfSyefggf49I2W+LX9
CiqTnEuEaBVysEGH9B6dk3YnEdZbDgjPGJmPitz6EbVBJZWstRic3xUJ4mZUQcJY
hBcixEmNeDQ+A71LK2yxFulmlHEDnY9K4VlIwchqIsm0SCzeTuXbsTxQmIvhKiAS
P50zPjWQOzw7yQAlOzWWTd7kLMea6vjmQuePl2ZC56dfpZSeFz3uGKv6LIeDvCgy
Pa/7LpIQFSJg46M8wovwv0vqHGr/ejJ4PG5RvvQnQxdyeWK6ulOQsPafJ2M+NYJY
S1fbPKfvjvRACinTTsIX0h0AdEJXscf7sulFCOcnE1jcSv22oJ2mKU12E2AuoWk/
pRmC8uM2Cw2b2wyqQ1oT3YgCVGcKR3HKk7+D0osEsS+cM/L3i+rxz5EE5NVRzVHQ
+R1bryy0VtLMoBGD8JjKJkI/FDYl2wWJqBwHDxbj8RQoISvIlAWt2OKE9TpSgM86
jXFfxDhsFcVdpkeVA/lVLOwEAbNTPD65zaMYSMDewk1yI5PfcwgOJWlCvQg8LAlC
m6ZAqJ+5sf9MPAbP2MPYDA/QM/eQxj+rHUxb2/qg9tBAW92wcfouqWXKPeqr7DFG
i7e8+fn/8ndkxrhzcjo+PiRmKnWyh8EK6+akfQPE9X4AAC44wqk5NvNtVlCmD5OZ
5B5XjFCVh6IltkUPjtsEVwJVxkjcr4d4av05SJ2wVskeFga6US0GfMUfGQ7+qNRs
Esrkn5UAGosN4ovbA4xRavT1hP33Shys3YrChJ/uzJfPmnTD8uP9Z6jcpq2Hbv1X
c/BjWOr5dftME/HU8S1GqQ5T5NJV/jYOs7J5Hj4Mr+L+9C1S2X/4VcQTxVms8hlL
DFi68e/uFopsU6oa9J32HKJRCkRhnLqs3ECfoIyfFwjCXAkGwe3kiUCTJaxz80a6
7eeKgrftz/M/a6aKGUEAdP8Nx+Q3lhoX9MKFgssC1AW5NjFxrXEXLdxADtGRXOkE
zYtxJpyGyiDjPL/WgLQ9Hq7icSJBxzT03zp/lLBxExcpYGtpZkG9gntzFsms9NIl
hcXE84s0zmgu4rY0021JvK2e0vwvQ9uGMlS2ja02DD0GnVlrM2RoBhnGlEK6bkzg
76AHNpgH/DboXdwpTU7ubav11TjUrhBYoJxCGK++ZlWAG7AJzlqzVXnzIFsykhIW
5JG+KM6PpcrtOmMmxJ9aei4VYssGBM2Jn0KVu15mr0q2LVcCT7aBvsElZXROK2il
eTxc5CQ0ZneTS9EA1yYPEi+RNboM7lTLNTsgHCc50eje7wx5Y5VZRN1Hw4cvZSpP
5J6zt7g9v7cywSo39U2KoFa6udql05CAZky95vqDE6Qn9Upg2pkwfjGF6eY/+pWY
K6RcmoK/EMHnX+kwhrqrDbB70HpKkdEt9iXNoZei6+uqivIA/2Xj/xwZT/9HWk/f
aSp8lmmvkRVxFsMnkTTG3iTdqJdXFVfeiaXFwLB4HWxUueZYyfereMGi55uNO8wD
nf1J6ZfURzv0879oIDLIQDBgM0wtpOi5z8mzmZxVzspo2oqvIsh5Laew3c56glgx
21f7MI6o0LTahduHPaD3mJ0iC8bDuagkRwu1XAo0SN/MU5vwOgdJiznuZCcWT2xO
VOY4wuMnlg+e8y1ScEjPTNHk+vJ+4Up5B8ZECqj+/0PNzN0zBXQflFRq9fnRwADK
BTcM50fKzgjj984CSnglOMHrPKgh2nAABidO8DE+TS7Sg14iRY27TzDXgozF9Gz6
tz/yo9Kv1s4+gmbnX07jLfn1tJ4JXUmm2P5h2t0X7Auosh48DWKVe25wISSLS96+
gt1P9Mq9sr1CNdTcnbgRm6bBbsK6AssTPZrw7D1LnZnNuc6VdtISjuGHUM6x1J8q
ydX84TLu2quXVklB1o8yR/r6iSrs4f1rBV2mfRUkfWintCgibH5w9xf81zV8kbzQ
qW6HQCQtkdsbZKdYwk/oWGygNg+9U6ambccbRhAqvoxSvkHDq5WvQ+Ig2uwqgX+M
oqmwgpc78iQOeL/+w/ndPJIsUnk++uyyp82sahACCAR8JjLwjxj3cqB2i103SREZ
8Aw88xFz2vT7nLSPlzKiJ6/G9kVU6bCSDEq4ER7//6iXivRYY3NKdLbAxGaYDBxM
pPfzjP/yiIHBV8xaD4YFRvxxq4Rofhr49NXOHO7+xl2UI/7lgqPvpXH3GUDd7Qyc
7QUxCcrkN9XgDWOGs70ht6xhfsqdwPDLRwKTgSefF3hLxXQ8U4Hz3GoMXKdGbaWD
KV8zSkfVcNmFVUI5eWPcqtSpOlTy3o2fQditaE/XLMYbTv5rtuRCYStjacinILqD
TdMai/PhorpW96UDJxgjMHVD1iFEDnMDAa8QEe8d2CG9XRxxyDAOUOlLlE5LGQo3
vXxIsau4GfQ2LvZvxO34R1B4T+aePPJe8lZ6Kl0RkqU0CKox+Hvsn6vjVv4YsIv0
o+7s7j6L9kFPS8VjoZm91+YgWjK8zMr1SreLWiiNOuI297yTBbJaSL0gu35Y15ee
NsD8fPmFvQu/y/DajEueUtTZLnyckcfA/M9Yf2vJXv7AkBb56rW+cbGzcJBqydY4
kg9Z6t88g8VkpnKKBw43xHEISjsYl4L5RATvEN3yKmv4MUBIIzjPZXw5MfpI3jLD
6eO8YOgEZwYM26VR7fZNyNsTYY08vzgOcfz0+E3yQvTDGbJub3CytNIVwRVCGIcq
1rWbRFuCOHEnRbo/EQHb7v3IxLpqJrW4tBq9opkqK3RULB2Nd+Ut2R7kcj2lRF5m
Cy2SrOAFLm62YTm14vSaEuypsiQW3FKPbbtEwkIBYezOPx5l52e+fQPwnQA3oZan
Vq4xta4wO8Z8F1r3+D5YkPGkwnCgRstVEDgl4AU2Wi94Za/8bERuDtd6bCxlnt3i
uvjdlFS9I/qMxR+jsp9sVNtehQEEILRl6j6ljGkA7q5HPBMUdYk3/InbtMBWAUr4
vvQA9pRcUXpurTBA+kbSKxbSfCVmVq1fF3NEcuhev2aELhz8teOqhaLTr3N4nLDf
looniN13V4FFRxeigzlPCLRCADI980fpI0d4NEprEFn+qa68qryr7bW5rG68aoDg
NzJE9ztHvWdQijpmCA23pGXnGay363h0nTBnTZ/a8L8h7tgdTVQRU8xc0kabC6e+
jIBRUa/hAryUZ0O38Rw+QO4S8T2KuCtKbgo5riYE5aQ5ikENB9ElmLsI9lsKCNJy
V541OVk+yYk7XefqnLVFirHGs0M9lJxodItedFvcm6hhizWugeCpRXC3h6I8xA4+
znuIdHGAXkXNM3HdPdVE1DTmb8zSM7li55bitXLOs7iEuyaPgv5a4IwZV0vTBz6U
rtzvaUi6gcJSnSaz6yFnhubvOuLEbGAh5kvX5wCC8eUMgtIk1E4r5qEXbLJnAsSn
xK7fniM7c2Bp5W1Yq65pRh08nBgVNnRMwxhzN08NrRteNPMv/uflx6exf6ucTXjz
hXIgFxoK6p4nFEQ9r42Id05Awiq7rigRTfSYR0rDp/G2PSeV4OM4iBuFRHtBtXU5
vL4TA4CzOLztCUQgKvi7+9q/HEdzbdAvUG1UW8yBrePU4cdCNGLRmjivdPj51GZh
f0+7IV6eIZIyQz2IHrjieJiuE046bKdMiXcb2DGSiXADvr9Pilb4GXHIha0n3Zcu
woNWOUMsC33NiiqFtuAlm7unxsgaK8pkRViHaHn61AFDv6Z1/lEfmBLpBIUjg4pc
xUR6WMQ3MnJ/3PwScbBoBfn2Q5iU9GmmAr5HYQIC1VmvO+aSsHYMhZZSeZHcCNf+
SJM04hW6HuNUJhbS5EPgcPNQ+tCt2ebvrDfUWikQDFcTzdk/3ivsM1jiT6xCGfOX
g0ZZq3XDzcZpt9gNLZ20Dl5DPePEOmyULhN0Xju06ZXiT3e3z58jx+I3aQQtZrXY
Pq+jS4sD4HZin38VovBzRicLYGKe0HukhbcBow0UvpO/kWwp5ahYKJc6WZTYB48C
+L7w3e1HIJBgnG91vZKAl7/3iku6TaBbgTBQxkxi+vlc5ZnWdkvFidmQ8fo0d60E
2oz01n44Ymd1Yo6gcSuetZmlqN901SHNpebRVGrd6DE0NhaoMxx95ycCEOmtXD8Q
F3vo1MRr2u9/PQin6U+mbJf2np5+XSVwShgGben/ph/xa/J1tfgZfEQKK41Szqps
9Xy1CYtPV5eZPr0IDap7i6LFXRP1rTdufWUGmCCroBa0gNxYkmaa3ghStHI8hZ5f
ldPZsbtWUaBdxdRt7vM8tJzfwsQu80dPjL4fCIqpYktXdXapm5GQ/tAeSDMahliM
+ymPnfD0gNYp5vDbHvqQTwkyqWcx/vGEu0cyCE9YsQBQZ2YpXg/579Jy8XD9luNy
+DNiT0/VO0vSex1O100hj23O0JTJl08KNiUC+114cb53F0WeVjzys5cP895qPba/
JaekD6a8BpIOFN+vmfLajYrEgfbbd3WiO5xRiGlGvWYPRxgThPwQZqNxvj5Ylydb
9PKsw3cU0UeWsentmZOZGpN/rHnGjzLjttdd1dEX2akSnrb06UDHPanfgtHVstSm
ehyZg754GekEC64/sFJPRuFinsUl3xe6Vh7CdElXrtp170NYPFMpdCUQcLp5AgPF
aUYR1NihZqAoBJ5KhwWa1w1mru8TIHbZ5RvXwJt9Ozp6+EPYmfS4Dym6lyLWzYYc
f+Pn9+1PoI5AZhG+UZMGysfJLN8pd3sTBFGRL4gZEOzTybNwmmaakO8Ysy2x3eRR
yPvk6cNp4P9J08TuCKlyA4FofPPiCRGdQ0ad6Ls4GSBITJo9CdhahWlt3mNyTbuq
X2txfgC4IAQdxSohQo0K/ihkwhJ9JLePs0uyxVKSTBdNh5JX82YvS1jO2y+V5zdC
E/VONY/QmZDLT9k/Ko7RNQ82pYVvuwrMKirWNhxgGlUF5pfFUOuN1ZQ9hi+0KVhn
4sFqL5LPQxj9PgSAkJxtcgYejyYCtXgrssRKBkHLQXh/YCnyVvSEq4A2yOk9DXP0
K33s3aK1h5toQrAWDembtV+LDaoMPPKwQTLgXq0DtKnLHvLIvIsjcpqgtag1s59U
W5tjYIr0jOZMQ9DNYRa6MyFfLjqrxhYJwJAuYh8i50gjuax9y3AL2wMtgLRAVDkf
QcSdDr6533WENPX5r+ptqp2l2YuUs1GTfGhUVUPM04YGPIXeNDXowBancPYNdquA
7A746fP3N5XIVXriQNP/jvHvmY8gzm961syaXIhfghRCVU5SBpz9og34UxSQCV4d
sjCOAoaUIXBXlG/jceSlluds9myFkR2i5uQ63kAB90+Nc5pcn09LhzfOTvafbTFC
2VOGRNI5M5MXeOrpNgHRZnc3RXez1AIgQCwM3PGBhkZGj2SKi35usJ+nNMfr4rVR
ngIy8GSdOCkBf922EWr4NaMN/OYtOzrAAOH9qBWs2zWb4AUwrGO1A2m1ykBuMGZZ
MqHzy6mvxPruQBD+Kx0xl2VXcgzp8klbwpDi/H202Ypyrtmyv5f8W0P313MgNC6E
xaubbsesd5OM3gkqKyVJ77uIXH5zkODbYWaEVP/HcvnHWZmZb4Wa6/iLRLcONM+h
/02N7YBrqQ9KjjeNOt6nWbm+ZMTR3xOTedT8Q16NQWXbLn53wIQ0SZetpQWLQSYm
lDzOolIhSMWq0Dg5dJuHzxuwnhdFEMBxSd1Jili3B5sjyiBW/w/DEZk36ygvtkTE
sY/w7IbsOX6x+QiMVHsuIEPnjeC017SRA2+uaNFYd+ZbRYFMpIx296AOGQELPQYT
CFC9F2BjpSWi5EyNKHDqUWcgg78V2w5Xd09iCkfiOWkOjoyqz+LZZoPU9ts8hGPj
G7CxX1xjQeC726qvB4LCKU9tC+Moc4AkRQ8p9I8Y6HGgD9/0htTT3JrULQaZ9tQC
9BgTDSYvpETJt+MFaFsZZ/vmmVBvHIX603m2dNV6dR2uAhNSZRwrfFW0Tg62h94S
PR/YJ5n7Z4rKR5pvZeQLloQqdGX671GJys0glu5OWe/vfSch8GvHnGVQjIv/L2pl
gShoa93HFCJkTju6xxxaKS0SLs+QrkLo5SuJj6sRMpNVKrbgr+vyLJUnEryBPwMU
ayM6IS+dcscuSHpg11qV4M5X7w0zBjHd/dplMq2Nil0Z7Xf1VqxhKBwaGMiF2C6l
FkUOoukvxr/+OY3PiOStksDS83970KwQJzoADpRED9PclIO+BGcNJsASe7FaqTKl
xWm0//edXqLoL8THpcADi3tQyhcFJcX7jAaFIdZqFOvQPGiJawZ3Nthz3hF+JJvE
8ycvOVdZVhXIXIL7p5gitSuH58K4ZVmekKl/kBhYrBneIBVsQ9GWWLq/C614McAE
PWxiS6zagFrart0duBVn8ODhKef3BWRBZHADPr3X+APDn654mtPY5OnvSJsF+O3S
0GUCX4zN6W2fmet2XWVt7EWw/PfM9OuTN+BibnbLbd4b9BiCVfrMGotM5QI327c3
P11aPFBEm2ita8YNW1nY2+khKIzQ36MdwlRIQNWoKgodoqbcFYkbbIv9/3fmXMY+
FmpKxtAtKTAOIrmbCbLGIuVjqZgKcigwk1ofahthtaHMSGR00QonxdV0Nz+uLTl1
DITrIghD0aVN3xmYI0pfP0unkxxE+79+66eHFnYn8uZeNf7Sc33GtaIv8WyDwVrR
8luOzOBo4ps+4XAkYRWdews2oGdUCfi5zPgx6v+G5kdWGUGhWmYW/h9BQuN5IrBN
e9JPLTsJ8wWWNBCnRr5V5/j0//GMRBoOXjUsId7L6tnGAfPc1Nm2FCJUnxo/Igsz
wE8wckc+ZbAcIATgNigVv98z9J35wpzSOLlMY/WIcIKWA4ufGi2lh59FSzA2BHRI
yziJCWJgLpVdGip/C0zybZwuUl+9oFXYXzaf4HFOr1bhwUAAi5OBgIMLfzIE18gA
OegS4HvI0oeMoIs/HRCwlJaf5lvdd7LSnjFqGCAfMoUp27uVqme8klzMEE1HEDMm
r+dv87H4r+XOhr6l8V3apqD6cYNDqiuuQP+dVplClA1iZyMCxicFuGgzISNZY7E2
39diBOI+5R/uNC8i6C3J+01vZKu9Xqz76uETTWQeRu3TwOR2zeorVugziIkp9BDo
NgvJebQCMjqcxzRW96pqPG3F01KW9zfjvbv6gItp1yh0Srq7gukSimm6XwoPZdEr
6TCqi+q3uTltvpgqx3dnYfMD9hSOIjFrc2jpYW+4IfwirQRn+N9IdVXcmaiDd9Q/
5w3lHRD727p6A0y1Db4Z8pl1it8cq1lTlkAYEkZOdT6fp4PuGoAv7+5LeER5QVy6
b/8/D6GxSOKXVkKqUhY7gJpDI7Ag9u1q5+Cn4GgxW/3HdiVliI5JaoeBYKv7qlk8
u7uftjA1Xk6r4Q2B14BAT3JP+5upas5Lc0X0ANnc4FpWtUBtkqOdGjLN3k4gGio6
yKCmiDrPtuhZNzB+HWDGUL4I93KKVayDjgRWPdYtIwH0mDZpeDjtP0Rw+zZHKbJO
Jy1xPjhgmvdZGqNSDZe86xnqIpGcG1J6zNMvV/YAkfrG8BJIpJ6DPWYUtKo7jLbb
jLy9ntXNbPP0zxbgTET7bL7NxUnlzUroJG5Q3yNMZBFg1nsa/XPsOv2UOqaTnlnq
n/2H/9XYA0PiFZBFbp4xHRxibAXMTuJEyeLrnrBeiZ3nKcBsYk8fPa8qelo8C+Qz
6c87XJ+9th7T570QM2SSNFN+wrtRhAdI06M54iLrQSSluf9uIR+svU/VjAdpflwe
WqEGhIJNxdncKhe4Im9F1TYRcNeeujcTXBvtBrmIL6rD1muGo3sMa+fhczQK1Pex
PhEGVljJdjE5Ye4qdUiqEfVoUlGC7DgGlCX35Y5kD45wstoJHyA4Y71wK91kq99/
nmXAQ/WLwwpwoU0RPqJ1O4Jr8ZKWxOtlN872ModkKztTYzCdsFL57I2BC0evZgTE
iqkoXppqxP0hV0Hc7R940wH4YYcyj9ShnRtZ7RrknlACJXLIDNLLZLGAbid8tz+b
8uewXJklT/NYRnQ+EQHdk9WCqmWksRzE2/qnFC+bRVtVrGxErEnFqa7kUHIzTxFi
RBiji6kW6fA7DkpbH59l+8EB2EOpbhc6sXA5grpibwbLaFEnyxQvbRLXhYKxIX0Z
BkFInkA5go/vBt2jUcUNLqtGAwLAG7uxnS/Q4kWuChA/c3rdN0gm52c7Vmz8wt32
PWKTJtkQtb7drNpAl+z6NZ3QQC758TQNXlMp+lNYOWg11XsRJB77gm0L/u+jCE54
VJcgpidgO+gpShbbCmjdU9SjW8JtpmMM9Yb7pYWw7s429BOPSmmONL3K7G3qWGAr
k55lda6Ao2ZGLMU5pqXzksHT8uw8vCSIHfP564OnNA72XAXLaIlyj9rq5d/WNDLt
DYSdcss7t1ZS2/pp8cvxI4JQZq5ktWiPmqLNHcsIx04+KlAYyF1LNdBbpEQm/Yxm
nBUtoIMO8J8FSGta4sJMq56+0qyr5N3r4wGU6efLY+UpbxUN9y7cGgk2KuQVg4JF
5UQ9p0Rj6GO/b1DUOyP/zESn0RQk879anzdRkSBx+t2SykbFbD/3Gc9DsfI7itVe
gER7g67g/XYR55XGTvnu2MRKemKhLGUjHKHzU382AUviS2FhJb925MpsqHKPX5qw
j7ivQ6Oe+tmH6qXgyalHxNeaToybazi1WJERw3rW68gvE3VqoYywB6/BIQqJXoCj
EIWilcXrxfYeir3DzytXpwBO0FDgBHlr3ftOJfKZc2uBX9PkLkS0r8KWGozxcNKP
v4P3v3UQdsX5qjVb64vwwfscIDtSlCGFSCvNnCDnMKBJXJcXKyCUCzXdbWt3Pmvt
q605nf1MUoz8PTm/MQY/dxPYKyd0eAzJQM2HUVGyVl23JgjRc5pgPWAqAJp72wCC
tHwCR7Is0DThPER58V7wGOV6sUH1DFzBJHbS1lJ4kdecGOL++QfYO3QonFAueahJ
AlOvXoO4BjVG16hOjPULCahFZOtYoyKo0O+24hApDYMIrsz9AxFcrWr5Q2HWY3wx
XfEmflTq0FVXpngclZgIhZ5Ue/L2DUtYWlcGK9NVYMlGv9F9ymsdD2yiM6Dzbsvk
dpBBlhX++HFjUguHe1l7rC5YHNqM2BPQleU+bgB479D1B9HVEFLRlPcbyHsFXrCe
I7Fac38Giz42hlSwWzxIQyBgBFDOqdjAOGd3cpkwjUbOSS2il5sm2M2++iXfZGFQ
LwILMf0pxlKKX7lbs8nyR097VL1V9VutX+gNvGuMivjCagfY8gIOXPzYhJ6oHM95
3oMGzNTCKCrV2D3kZ7aLFASyFpQ68YP/s3rzO+l1bqhvid5uqvdOIsmIZ7zGCuQl
/hquTdaW4u/AN1xIwmVQVMm7LoeOA/NMPPv8HqaADzX8x9TuJAWjEQvWH0hFYvFK
1JKjiO6Ev56Z18wpybrFLsQeNqxb4Ww3wiJLCFNj5BcaKaG/4Lo+4wVkCICnK5iH
bLU/h/gs/UAwyhv+OSmygx033GZHTSZXfL8cLaSOCJgCBk1Em5HWz9Max2boW5RN
me7xONyFNBOr7Nn8SsJQpFq2G94ArDhM7Qz2Ome9QUXv9ejHwnj1oON5T9IBsOkX
6FYYdKT+3t7Bl790KSemrvybTrsdeEXYtRPtMsTaAKawlgUU/O+pi/f2e9EzXGJh
LwPjL1PubUmOb8TiEyDKKiGK7T8DEJHrn++ThL9/JgFCb8Na4tg/IKkqbxta3gt5
WgdbGCCe4ggInWo7MLBGa/0APC2liorJD7tfuPhJhCdMy0EeeZiSh67n8xOB1Zt6
sjUJT2UvNAmCNo3ATG4pXtAWRs3lHIxJvj/SY9LUv7ajrJDTroWekSG3kXYvaRF3
ODf60g15Vdijp0GbzNcKx2bVPXQQ0Gmlqz8B0R5b/B7AZXsm1vx407ymQlTkKXvH
8bvBf6v60OM0Tm8Nk+P880DkdTZpmQyvy7Fi85SC8Gdzd6q+B/NJKlUL85iEVFxj
rh/9Wq6KhODgETbjF9l5Lc3b9bHpd1CqCn/71VYLjs4QYclu6J6fBOc7Jifa5Dj/
fssHXjaNZpFZATtXjR9G4joB/kG7m5yUtd83MZEVzDmyQCX7/2uOM8zcgZonbCk2
1oDUdoTBc06JHQilfD1CzYUT15RNO6Sr6YLL3+/XaNoGErODnHAUdiMvSjXeWj7L
QSoY8Fc3qu5hYiRr05ANBeyrhwfYDz8sHrbJ8/hoC4y42v/mPW35rjwqJP4gT4jt
cYFkzTU66lJeqKLMdfmEPvYbl310dmmRwYuKfQ/gWQZ+VgYdJy//zrd2fPLxgAtq
XNt71uSLvVYLGV3KGizPc6tTVMgM3HS8ehhdEuTKGX7nIlI7hETwAHxsarhHWHH8
js4BqxOF/KNd+mxycxwc518hkpMVprfmOkBLa5Qw+ln0y7wEjshbHJGRIc5zGBps
Ix5OoX/rNUfJM8KQnaANzSrVa3VXFc6/D7WxPpuM4Km+1N8b17wFwdXi3JvBXkEu
1FUH1HI8xyU6Pbnee0Ni/PkdH5K6gK/o5qyo29m84YX+b52K5V0HOzmcX78bC3oE
N+umgaqBUwc9oz/DXmnHSaqcdyPBG/nCHShLBeswSyeftk+SBDUZYpaAKAx1FXGF
2AYChHC5ip/wedDUEtOpIqLcwRZAunT6UiAOaJPbEl22fa2J+j3XLZUrylQPoVx2
GzVsnOa4tZoBnvHlrU73tWfA+Gzv7nPEkZ3ieoznlkhqmRHDRJuxYgy33hYI1loK
hraRwlGqnwao/pYA0icFT8/JHq6MOWZpmVWlYPnXqLn/YIxQdH1L9SbrRUmb5loO
XbnDUfWBWOQfxzaQrPOkmMEMqO9YgtjzeHJ5x72zmsSWLlASKqt2jgVVptN5kCK1
WKXZMY3KWqyO9IG57qqnZiHEVFV/iJWYhywbTksRio58FyNAKwvJtSuylk6v0APE
o24WTIZTanj7NZmQPMPQbBSLn/Fdx8HhxdE69vsFlAszlxXE4E1D08VEOQ7nEZti
8Nm8067BHzUECr7Ky3DT88X1MtIynLM6CIsDXrRyLs02pS1aPuJbudvPqx62l0QP
v3+vVhB6AlNYttOQbNur+xkeo4d9d6uF7otP0cPLoYtPtkxwHB8cm1kamORPw6vD
6mZ7xOgAGpXMFQjjbn5qgL8xF7Zf26Mz0qSy8PVb04XGE4vs9RXfotdryB45SoFf
SAkSCZ/dAYYNotA7uJ7L9/OrnAUw0h1DU9VMK0xJL5CSM2rUN1RT2HruIG5pIggZ
yD43GjkBFKSNgrwSazad+znu2W7a9zs4L20NJYO2lrvQMCWjmbvwAq4wDr+WMbE1
+QeYrd7TRGaUPtMkOwuDIHEa45k31QIfUeUB65NXCrvmIUSt8+LukkqxxYz/ZIVT
b28MaA4pXYOf/Q5UwcuzFHhAfE1+tYEIarEflgyQz47NTDebX0Js71IykSaMBUxH
Ptm7pA+CITgSDvJGqrL6316KUAsYuO/MFo0EXbiINozaSXT8cOXff3CTj0SIGaNw
XhoI6yWQW4ZjM6B+Gyk79+M/aOucNmdM8upuF83ZJfbgMTdCNkdtpJba3HR95ujP
pz1jKwMoDWgk65ygHlrUqmikErJ4F60+SYSYnCivEIP016NL7u6A5OhGpikuDekW
5c7VJ6giOdonJxq6vv+VYWnlrXrqlNP16SqUnwP3t07yGtq8f3Oop+fBueWP0X1W
v7yW5BXLjMgHJhU+ixsEkpNZk4MbGxuvX+NDeJr5FXgqBVrT1glbLDfhiNMflDOl
6pvP3JF3nIjaLJsIS1cF4PiYU44MgYIHnrC8puJbyMgNFqUVKXdcFKkm2juBCD8b
VIGJBSakayXhqXHND8xwfMEqfDeflyW2+wQ81n2QNON93Us4pB1xLPwefMlWge2j
VKtuyUJ+hqmXlGXNe0OOa/oTclo1K3wpo2B9Vhm8l63BahMDevYnYnjG1qwY9rrB
rHm0sG9gwA4j5W/eecXAHkR0RNAF7+h1GUJ2mCdbshzebB8WONqDdefmaZF2t5Ar
EhZ/sDbEvSFFjbl0g2gVrlHSxmwHp0P8Eg0Kkjv44q9nwMK9EgtV/5hmZjibb0F+
3O2ToshyJyVkk5bV9k2mq97mfYBWR7yX4Ilcx4OtmGKyVWMpcK0mfKSeREeGPLOz
/M3Gv/fdyz7djG5YrqeFk0weJnp4iy2SfQarM7GYYt4U+5Db8yAdM5+msMErH/RQ
+ZomOeJKzDi+M1hHeK7oSq4jaXY0qPPgA2VtLKF+N7zWKN+ye626lImV6zpIW8nq
3s3UBEH6vrbqTeVeaASJdhyqUaLV6yh91NrB7eB8idGWhBd57ObXgrS2QnqOX1nQ
jC7H24WHCbnFoTsJcQ71okwPndZ85eQQ/A3HVQutNIqOvsezAkCsK6j8pbkl+CXT
8tYMpMaQO6tOsnwEj9dPJP3c823/zVzJ00PH4jqqDhxixON1JvqkYsWnyvaEkGAw
iwHNHWSMe7rd1M4hfeIOGCRtW9Zc+kJMmGh3N0H8+1f06rrVKmI86PJZhYBxjLjQ
aAG5pjQcCmrIwSibEb/Z9Y8ogGDZLdKvwUR9F/ziTpY1X4lP2ugQ/BAbQ9UlWtyU
b9eufVC5JFNNUHteclGrqQ+H9Igy40Jii5njRVpwQ4qN97hp89qTczf39boHw50B
9qa5REu7PvjoRM0ast2cdgktxTF+w1hUdMl0d6DQyKi9sdrjs3TREDMbAhecBZ//
1KWyUlo58fWqoy+lL7xCreu5Lc2SXmmUfZj7Rkcuh17p4Fdutlxt+71vDNwm0RY2
2q7rXe4XYbT8pW9AxTsLfBCUqnOiFySILM7oeyvNv/Rj52Ax2+fVijXGwjHd+MnX
hFDXSGkWDonYq8JNHpJ6FwVcPilj9Kikkj/G8weMDwaSSaFWByJvEVnb02j7LeDI
kiRPQbyMfgJA0r4rOA7QyIx9gzajK6xsHJptR9a5iUvSl6KzZStm96sI65X8s9+1
2nRwfx3MrJInW+cawUAky57ioVMQEdeEGujhwC1VUPcsn+wXiezI1dWuOTiu8UJu
2ulY1W/oTgJiQ/rq1mWvg1qAmjOMRfDRsQ8KjlDZpaEjR/L2zDZ3S3aEqvAIZcCF
dpyrfIX55z1ut2lFtktz65nR9X8k4dQJyybndXq7wEBVw7gmaOL0NBYEPe8/L+vw
gTnq+F5DSrya64K0sd/m6jbXEaU+1Hk/27nzwI9Rh5ZewPfi62f3HzVT+FH5zJmK
JlWiAQlAWs2T47ykckY0nzZBJTyRvWrvNVN0L6VvruPaYPqdlTopAWZ1Pn0y2cqq
lwvuxbxYTv82oagxbQhKrZ5FUpvyWzSPqhr5aVUuaiZVaZdBLejrMoQUf/+yoR9i
IcBiIlG38JXHt34tugkP5uAtmK3dtcvli6ttg1N3aY3z7uAtz57NMeTg0AZAm6uz
oHpY4VqVWXupzJ08l27h9EQWTNbc3aocTfjSHhSpz2rPsXyGcx35CfqlzZKvbGBC
okNFWPrnVqAKLvHhK8+qKTEnouA1uaCdZefk8lu7RHwhN8Nkn9ih750IB51bTDAH
LHAWuYG8KvvEkGTsPZZBQKq85E/fytlHd+TqWd9bgg0ahdnEihp8OlhfbYoOoyVe
TkCqEs5ePsbZqQrgSpqfxQpHL95AgAp8MNe/KDmI2XDvK0EZCLlgTG6VIulzPyeF
oTTRqx8iVePL6LM7/SNCjDxaaCy+Z1UiC113JEnq45h7vnLOvkNJiiPmMRP2TiJK
tdX2aWfCcxHeg26KlHiBJzQAdXBzmH34kl8sG+5OmfnmjojBZ0fhSyxECRVA9aiM
+l7ig8ZZuIumxjwoKEJ30GZ3OdncG5S2OA8tj3NtVCgGismjmCyM62I1m2t6JDzl
zkXgWIvcsiyTxnR2PvIIrGGBOHYVOy4mWFTqbDCl21WN8UsOeR5pABoWvEWtJKaT
Ia03eJD/WrBCiejT1OGhsxZo0g0Doe7C6jRp06o96TwHHmERYx9ChKJnu/eONYxc
x8gcMvojCmYYu8PJF6yg6haO8QoW83y6M1WdZPZ5NuKTOS5ui5Ceo7MxDznTkAf9
urax1ANhp/v78zZkxQbYnjyli3jDY68d8X35w/23wzib7szD8w4GrG1ESIHdg7xa
HmSOaPbiLADbs8AfcDiS2XFKjG3EkmaNIxnk3zr79h1TMTFO+m7jHfWeYvEsmpQP
eo7/Ph8DSAp9ZLa/58I/ZpyeM/KI7kJyP4X8S9QfkEO2gjsLNugcbWdrDEm333DP
KCmNt6ST/bxxXZ9EinRwDJpsHEqwiwDeOyZOgqtsh2FekKtaRu3x3iaGnllQJ9gO
tOMMzfRXUieHw0AUccb/OpZq3auUZghL2PGg/63P+0Y7jxGVW5wfHzGnTDgN12vM
vpwMQBwmddCL5BNjx+wgvRknNiO3qDdu7cbnN6MQXSolOv520ynB00wF/4wpfTil
oPWkL5UA47S/1Im5A9CbZVr+ZARW8JQDRCClvebAQnuOUpWMAPvZhmb0YxNy42ZT
1V0SfNWbME4hUMkERzxSiOX7iautz5aVbwOr0JFGq7bHYSos0kOrXLBBlTpRpe8E
5qt2sWER8Mx6TqwXoHiBf5rRz+kQddzbaSTIGFx2WFBp8/BKCgDGVMr4Pgh6Xq8r
4J55zSUNjqDk78HSXlaLEv91EA/mWwuwhc1DfSV5N7Io4pWRnQYgnMyG93xIksaa
HvX71RH1HW009/6bQvVNDw6xM8u30Qi7GVAcjwWET4dEUmGUW5P3st4vl3R7PD0Q
VAzxeT5qe0IdxUkS3NZrmmSk9KVwyzQBaKvwAvVPXrrKgi25W4EfKFbMnexwaEWH
pTFhQBFvunOE+Cn+OfJjcj01JyY+trtIdaaEcDCROMFQUeL6wrX0wKYlHRvupoOH
duPd8fcBC5dx/5iL+cnTmA3NlzNcizxqhbz8HRANPxEuQjHmNyvqKtf2s49FtljM
GtBFdnzBSVy8vu6Tgp+kYriAt7h4wd6h3MsP3aYjtlMRyyHMfI1zmAz1G02EVaDa
qhqCFN5Xxnqsh65URAPzWBil2nc7vxO2LnwaU8kaECWfN8oX/eFetC4eM/32ShDx
zzZ9Cl5ZnFcVPNdMZlYJthXUM7H8rh42p5ls6OXsialC0ykFPFAuYGDTRqmJlz1o
ZE5WvcZd0OirvYaHttGKWNZm0MLcvMFz129J45KmKLy/qxLmW2F+/YFazQNwHqxt
A5648L/KFAvOVfFWg3tDFPBBzmDA3Y1MSz/oblzB+UMDlaxLL6MmHo9ZjY8RR4MU
a5JPy02yTqQuFiGrmqQAKbeOYXrjm7ROWmrslgQF1XZhy9qYjm76nvU3J68k6ZK2
AzP8Nn0DECbzOISSJPQMyOHGqpHLiH4pesdXcJCigdeRMziOKi453YtfSK3h9m4J
Mv50kuUX+DmQ4rzw27PJ+3ikmiKsqIGxzUJPcUlioS5ihLAdi90c+hg4ppEu2CDD
ZtgG4vywsLXO3Xacm4RgH7rEpQHmv6kKjEeEa/ozKLNSIZXhDR2kyr5e7KUDFcxP
RvLOBt45ciAyhp6/aHiyR7a2J9iarcnO+9LSsEpBWJpnV+P6F4SvhKSqIHSjdVX3
5pvnfPq7QvHfQJg8sIueM0hF+7ap1d0BfdNGisTIsxiIcGoD4TQLPbVxIZW5UwEj
9dHDfcbKm4Lroq6Hq/ybntDjsNNyQ7gbEYOsWNssJt0c1R39FWp6GixkAo3uivoB
R/yZecRcu7dvwFG5c1IPexkujzOYHZzUwvQ/phE9TJlfa1oNydvzCeBaPhs0Pa/0
kw0MdXp6qWw4GQQbRCd4vIqBw6ib+zgRrL9djx5UZzaTf6yTIUCsZFelf1e1LNVO
UpEp0OFRpLKpn9vuBN1tDtNlrZf9qhB0qbk8uIA9hW6Wq4uiCgdc1nIAd29j8S5P
vLYb+Rt1pC/yqWFcHOZlseH7emS91DPdu9nge1CyCjLUMcXt7Wzj7xH/FU8JP7UA
Fi//vuWgVqKupPhvMe4i7zP/T7OI/q5Je4V5MtatKkgTQk1Pz0A/WcuLVHRKNk6u
Bvy3nFwmAMTIFeDbV2D4Y8GMWLp2fWWABTcSAE4toVGHSle9ptSaNiDoi0cm9Utl
82TI2Nv7axudYOcFOStcHhhdsucoQu/OZiIB7ybf8bebMxEUotgsUe744OqAWUpC
rltiqWNC7E9QDRjzBlAWTfYmOR8uhHjzfmx5EuqZHH2zKCnUBaGNP7vIW5DuabsB
MV9HVb4uysrRnESPJOfnQhGQTuLqJZDOUc/YyhOSzDbqL4eSicy+GSIK0VdYu7ti
jAdMeI2299PXPOGh8kbG75fAnyPF+B9R8db3+5mHZTodbHx4k+VHlKs1XHDA6i25
ugRFWXcYcZzgt14zlExCMB9aCvDozmGC+9CQpUWHh7qIsctDwB3pYZqK+Z/geonf
HRQof1UBcd3UR8F+TMn3V8lZrRUnHcd96DznxqUfm/ny8g1Za4iR/S1LPhyNXQHd
0EB6z9z/+CVVKKwvPVMmGJv5yzDyoQoa7yi4r619nuzlhWIVzxF88tTqxxVAkV0s
EWJX9BcP+NiS3Cz8t+XLfqzA28HArQ9FlRKyp659HvVYNwrTMUFW7Za3W/MmMTFV
wXlB9ACs9iuEFWH9arFSPekRGyH6O/TtdRRvKPLoyvfcVGyIaCpO8bmeSfzPvI/b
rOiGgG42to/xy3wCJ3mZtG0gK0RnEhKgK7EmhCVPw3Zt3/nFg8xJYwju6HgGSHm/
ES/4Zdyfz8D8Sf8K6kmMTtrLUspR6LiJQt+50LILyR0HpKWvl4o5ceJDFI2GIvU4
ITRbMEFCtZnOKIRpmzjqoukI8Ndh9NjIeY/jeXJTuUSzcfqt79tKAoAWfAe6qdg6
q4cwm+UlhV8vzuPzBb9Uc0ziF2dQMs+M22NMB8bR2vb32nwx4h2Bh3uLRizTQ9sr
QDTPUQEiNrFuXmtYQXY2+rDAr0nrZQ6+ahF/Y1CgTnOSKKOdjSU8g+UjZ5CyhAcs
Ql+uZSgRXVEw4nVaFGysjJ3COOsJas+7nyK34DSr2oSwqPE4yfVZTKNzIqbsxVzb
Jcny0ZgF6goNzu/z6k8IMCw6X/jL9O9MLvQ5YUwCtxyHjGRM00O79SR1pyo2sPmK
V3vbr6TZfnQByC5vkMiG0OEdKG10sOiy+d/HqCmJV//54t9EykNxbm91lHxPX+ll
3uhtaISHTRpe+xsQsIjKwBIfCUOZNeKClaQxZgXmpsYsm+YQR7CXYqNwrxe5k+Fa
12MoBXB56vF74MiHLu1WD5NstHBBK1GnqxtrirEWkn1NLsgdaK58ExzF8GR9WJ4Y
VbzjEAsCzsU9N62ABJtZjna8mIlaf/zyo7Gkl5HX/wc2Ss0HiC9fvlTv0s/Rw7+U
fluzQ+/VMuYNDsI8co4UATHdw818lT3Wczr+d/j5K68h5tJWyCM6m62NWaUiuwTb
sN2EwkQGY61ieDf2wfaKcvqPw5clvaI6NMO1PGMiD6ORv+KGpocYW5NmqNlhBM5W
Tiwkgjy8sbIiN15IfrxuEQH2QDVkTQO0E4Jt11atZovl4BrkiqE/vMIRrsKgfUx6
wYEGiDlV5PO/X0Hmb7xTk7xyEEWNSp8/1e7IcvH6MdQ2A7sn1wCsH3S8SuPark9t
yoOOPM/jnn4+PZ+jEyQ/WVo/PjXjH2ca1DUcsN9c9PIqyp2TlCfjlDr9Hyhl1zz9
op73bqFL1cl7meWWggQ3Jr1PTT4/RYhGWFiI1epeur2ahY4gQeCI3N60d9o6bIxq
QEi5WibOM8YGvuJBGqusV0f08ZJGVZe2irveEOuhgYuueh4SOwrxp7C6SIDWd+bE
AsNnwmMRKQLdM7EFB55C0aAk0vNMb6N2spGFQumfYln4DNFTQhDQ0k+AkzAccKKw
19fZrED6g1pZy0VhchoBv1NCVssnqMegmnDx+mFW9oW/z9CpkQAP/vLMioOe81dU
0zsRuTTTHrCIlPK/JqT8vbSQ0kG/uc2i3gq9ElCPCHjfKOUmtgqdKRTDC/XUxuD6
A87UKX6sFMhQsLjVosb1TrVM2eYgrWuXOoPBnNhi16B7zP0CoGWsjvxkdJBY54NA
E9hCbPSxjC77Fa+vR3SHj9rB6z2RL7D4vmaGRuzwryK/oZqtJuVU2txU4A5kj5hW
J0WUmlJeqSwi/N+OCzS+UFbxDJS81jbymnAuHUsu8kzb2AVtCh+2bSfb6UR1COIl
uuVwJuyaDWRn9NpogRQR5WM1THtf/fh2odj/pWPl2KlULpbbi4LcY9bLj9gklhtI
woui7ocMdG9L2p3CZP27HqCxhbopRRNjthWqtYuFtGF7eHiH7EX7OKvJp1C9LzXD
xsAH8YDxAtNVXCRsCfn8j69gHmzEbV02vzlTaWVgMe7WOmqQ4JtcSLL6ARTmaEGq
bYwzDG9BVUkroSWcb4jMnoxNXYsiB3rJ5zKD9wCzz7TDaXocuQH8RSuomIch3QI1
bEhnEFGbR/7rj/AVpr0RDdcSgl9lTo916BEhMKH92FM/mWfbNSU6/990JsnZgZq8
CEzD79++8OWj1AEv/sqRUgWFqGWx5H1+c8zQ6Cf7RZne9UlwgOQRormcjuwwIZ+S
9YLLnPcDvd6axR6XB0OKGebIDQRhdXsmDu0jmST5hW8yzjnCoV0IZ3Z7RQy9CW1M
RVYFh0clD9/kxcPYc2A4xp1ZjV6wRhqd+a6i90qF/H7BTMXYduwy0s9QqqnqllgL
dftts0ymeH6I1nAMYaMh34ft4HxiiDGAhCoiAU98/zp/OMtKIB79xFpl3l/2Ohk4
CAPLX51/XFruzGOwKZCQ1mFX1CcTB+Bib1vZ+8UzxkZnnadR+6BWF4cMjanPTk27
mzlrD/jrOMRvl+iff6IqLUbauTCRkYjd1ILY7+GcGCNwg+INe16Lec4xNvCq9HC8
wT0X02ZrXRST0YoAP5D+DRw4B/fg7y2BUb2MFBhwv2jLff+r2dfISrjOyYoyUZ8x
wYIYVnduoQEGZlMh/6siz8vh5Ujmdw9MnHQ2cTjLy8G92oCmtWzReQP/ucEaEYWr
ynUMu885cKQB+jxp7IDpGmRHSF4u0NHtNrH8re+Z294F4PwJ5kmJI8DYHG52fP2O
bAdNPnOUoSxT4d9eyLv46x5k5ClGw1R1AlVjpj+Uek3OD7JfXhD1xhfU/DY+Utn9
c1MySHCzd8TXqNuSvWpGNkhXPxeYoHOO5DRq4CVUUL+DpwmLtTW50hIO3xXT5enH
oTVxKgUrE/rxBGaXPgJJfBPuX4cdvlXx4OMO+NoObHTPbvxlggreD0J1WPviCDTe
h7J9claqEUxaKBcb07U00HZvH2krShP7RCI4GhcDNyoWcByhSHV1nb8bXRjFSziD
Jx6R0al3OeqbYU86t3u7KQlGP4KdI08+Kylz11t3wW+ZXeO+m7idxONPPvWfNrVE
fR1IH8cUXqWoOdPB5LoH3/Q3LKpYhdIV/Q2+GDcgdemFiINhqqYIwY5KQWPxYLyv
ocKL9fR2Zp3zDhUX2dSzxbMp7DnzM08YKn3j3Swx8oyyh8b29OACRxguUCMK4osp
t5OkN4UTaiD0b6/7CWjW5FxHuOorzt6y37v6InWT7BTOd/6W5B+WR5zE3JQ+uDjp
a10iJj+JyNWKmlT95V0d6LNkWLSRGAkoE/bn/E90RuFt4A4QiNLmgu99Eqt4mcPO
YsUi0quLbjqsaDgJ1bRVv5fzVRZh9m68X4IqyJ80DcRuaJHXFNLUsDCh2sssGhES
00XUpEOuLXKAUGVvz09ro6dSZ/wm8TOoo2qznpTXYPY3QaTa6UkUCDJgi8Xo2DIR
qdg5B0SVKGEaEiHTWdtTVUTgNNsHYMZWbMgWMYoKqp620HvqRglWD+pzgM9BmChW
oGt936YJGUmmcVJvt39K2aDLBp1DQL9emQcicwd3GD5TVHfwPrr19skBLIU6lbS2
2ePiEr7IWHTbDXbdlBgauj8ja8XY4x9o859KhvydLWWltycx1uKOMsmRex5dKG8M
sgtd2DfNNUbmtOUIS+VM505gD2BoTP/LKOasnriJj9DC+vzu/3V7ZZ2eX7z+X3Qg
/i45UgAFAlEUSdlhvIZykr8L36Y1KObioYIY4L98tKZS7zXb/0qjhLHazql8VFJu
KOhihQrNjzuCYNztQjy0UsioIk2wcgAmoAfmm659t0d2iDTeH3hTSY/Y3YAD8TLH
hmEjOiWvylg+ufIAPc2CzgVdrNihOBkil2ONsbZl4/68T5HNEQIingTzq7k/ZiHe
hEuia8gjgLBPmJfVXBfBmAs9IieDTJ/+GVhfwUm1y1fqgLnNxoBfUgl6OCKEGR1q
dJe7sREw6Q+SlaJX8SD9njfYchsKmPq98sdBdTlaR0dmqWwsYx889VB9WA1lknhg
sXOEg+ZnODWQ/VvEM0yflJmGQa4Z191sBQwqaB05DiVC/6I3ZqimNhkDPArqh4aU
r5U1jHTsYQObeqSlm+ph0G6qnJugT3aebaf9yG/7gdoqFv668NGCr8fGKRFg9TFc
8IlLRPcaxLTIc/koaihil54SgMMDn+82tIk8kEbRq7rGAwpfEyFC97CcJfvOR6cR
NhJ92kz30H53acibl6P3yLogbR90DwiBZydUcNGXvOKD+0H4bd2FIR1xCj6zOJId
JUHV8H8EHBZMFtvpkIfFytX0/gjBzZz+4UQYU6Je57uTbyOZab4cbMh9kdaN/l+5
bzLBdYMBxh3a7Dhfitkt6FODszfZi5uSaj3FVPRwQnvQxeR7VIUH7nRMO/B762+U
J4QjFKejukWuUAwn5lO6sHm7hNiPG4hQGIia1Pig/ZvWOhsOFB7HU5J9YV0Dzz9e
BNjReT24RcISUw1RPgeKLLWYF0F+EcXc2URyudzHc5280U49ZbusoM7gVeXpzwLJ
hXHibCpNPv95E80ydkuvbKp0SWALecHaq94UwaLHbm8RD9LieNT++4BV+dEEbOLF
T9l7z7O65yCCdf5uEx+xsGAaOLL9dCdcU4mI7OI3fqOgtmBGc313/znF1ra9n22W
5N1/IU+lVxYAJW0ufHchJ1OIv1tfuP8y/dI7EDcdQdx7wd2oY9H5TSMo+tGZTfot
UG1fZPFS6ILdTqTORUXQ7AdK4LGjC4dOfNfmYI8pZQjPRPmKpAjqIU5pZWE7xvEm
7djafvivLRSo88X+tQt7T3OO1AKjdNzu7s7JvUhl1WEnQUebL+/OExrQDwlInP7O
n+dUGpBxHF3zEbzISHh8zVcJbW7BipV83ux+h3+U/YHrN2Uhy6taiMbQjR+nQVgW
M3v30uLIvHlI0qMtmYfLDgOLShcDv2MWz10i869XPJW4zKofHExIizYDUNcy6X2h
p6tME3m2FQkxuws4nFLcKjvCzSNF4Y3M+7vi11dDTkyeXX7Gck0dmOi1Hb3pY9BC
ynGjCYj2JB+J1Sn4MepdD/fG79Y3xlAkeNLY2yi3tUTtjKLXNkYH1z+gUODtsrs0
MCfN12QKfxBo8H/QAPqTAwRkTFOc/I2kF7CGrztf/vVl/ixHO9lVUVpHhrtxKwkm
zYXYs2jRw9uX2pWKypkfCFi4+OJOT0+6Qxfh42yMidsoLUwz5BcuSrJgHEqKfg8F
nRMAgEzKz59IkBf/sJmwzmV9+vo30iAaVABG2G24p6xk3+lgBoURMptK4NfVIuXG
0y4EQyvv728yPWRnQ/81MjVICo5iha9thSy3dMS9wup1j2+GjXYncTQdt1qY/mUZ
HxuIfpdinck5jLTVj3LPdYNGRIZQD8oBALnD5ev+wlbFA8DHg8n1vPn+HOx3vNDv
nK8Cf7wt/wmuFfNFW6mG8/te2eG58zeJjhZmk/WZ1iU7vhX55/cbTkCs6PhZsY/i
0XUhfCM2A1fGtWX/Htac6JuGsVOZoluKIfk6GXqA7FPfRN+uOEQWuW+63XHCUMwH
7Oe64Nt646AOhdzoQ8Q07GyGcL/KD8b3HEvSx/E2GvFcAHqpeWODgrH8gkSpf7QP
NfUGjMcWQg5sH1uzZ1JVs99SkdHJ3o1bjZaWFrCNYDdA2PU5DPm1H0kGHJP+J/uz
SBahOltTh6GMU1ALmIfPydxvGZO7C3o93W2D3Ej9ZLbd9HkuGq/49Sx2fxa9yMzp
pIyinbUvEUOpGcpznqKCBohkmLtJNdI9c4HzOoBAylz9wMNYuKNtnNmGZvE6G2X/
zBwUXsZB3a5F6cITIqji3jeIgiGWRlZUxWvGeyrGdU0HCMH0tZHRZo2fzUN99FVo
Zyu8RVbtuaRzNVry0zt1m/kWBnlHKyUkpvjochbHe2QF9sMWUqJIylslw5SER34t
DYbgNM1Oi1acX6FMnhoiRy3gZ1UW4jI6AJ97UQE77GJmvn9bTbyEp3ElO9JwM359
OYUkE9EK1FQa4eKQlrI+TXI/qwm1u33cPQ3cbbBB9aPMlvHq0KuOo5TruZ6c7xtA
Tj7hLwQBY5Lg/gAtccEbycfjSrkhXppGvqLHKsY6A+OkHz0suCxqpuBK6QYluEsr
Adk78bzJeQxatX2536fMI5p8pZnYPHOBFZU+yRc+vhh6Yo8pRqPV1gK23OZkgKL/
WuBSDyHLmbF8dgaAgust4bvgmwLD2+XIsbAVuakSMm7Jp+oLCopH4FeRL3lFKH3Z
Y/wndEUnGa6AMzOwk1/kJJwxzJqD3hiKk6ozrg36iKRTTs8us47nXFzkoJ1wyxW4
YIIIyda+T9nUnHjIfveuWek/b6Lp1fUkcJgRJCJY939Wk1v7r13WIj171MQdf8Jb
/t1VPfQpYX2BJHZ8bA7Q0XBr0tXtFaHdajoWkN/PaO35jsP5dE7AOSD0OO38KG7G
d58SpVVmI3oZ607e4dnzX+ncPZXuMz/KsMKNOKYvvgX/64gKHxssL5i8jICYh9KL
yscwxmKmLQdTNrKVXbdty1OHlQTNWn0FwLQUF5fat1Qs+dGGBL48Oc30s8bXYK6D
3ihNdeH1/AMGXpP0nysPprj/sYuYmIixyDvGL+vy++onAaPf/+t+KWlSgbq0082c
0aHeEawfLRbljuEDcRhNuSmxNMC8wOvHxfCDtl0M5qyOjAG+Mn8WJU6sNfl2czpl
MXW0zH8ZbLllS+NLl20oAf12FHharPP4YKUxrh5G/cNLS9UUGMFXPJ1YTcZVed7m
nfSBXe00Znek2eOL1E9mrQ==
`pragma protect end_protected
