// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
1zLZbFkTfMLqd8KH0yFoYfvP58cIwEy1rMwTx30eilQUDlW+j3Y9pVuOyIPzN/np3YLcSoN07bJq
AnZhYAgJZQLMS4JpY72H9NR08PtX6WOFDBCa56tgQL1HoU4Bzbfd7GvxKXiSd/sLwhuffSbpyDtB
wY5+yOCE3MVifRSKDLu15D7CWZr6fq6akS0U77mWbYxPOKKy1oTOrS4+Xl+yAsx7DgxtCiC53er0
lkRBekN0a5aHwqxVw9FF4/Eygd0WPv9zY0U1FCnWkBeS9wX3ufOsBMjsFU6TYkIV4Bh0cBpaBzyO
6DH4qG4CuzsC8IvCCgZG6o73/H0PSaSsTZeSQQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 24016)
7mkZ9cK/6Bj8kUpA1hVhkZti3dTrv+8zVlfvSlQB3DnP0LyG+TXcQ7e6MEEp7SRjpyVRZmgLmbE/
U14ujkZ1AcdBvZ3EzoHU4f6La+WUi/D6NSPmeZGVashtkzfj9cE69U0138hEnKydgrzA+noaiqxf
Ehf16ZR67tsQUv19h5j9/LxI9zXEuZX8z24ftiLbpFJDUvDmw00hvLYVaMBEcNt81gZ4oUkwpXLc
yRXCAVklq3JwTOmTSZFbZrMQKDA18SOuxW1yEpePsbHkBjM+QMO0bQsbJvFxQAAGdP4GPtSo2W4B
d2S7SFl3xyYKmM54GPirmednWFEUNbQ/jSbfj3dLlcSHykcfcO2kQILs8WqQMqaU3DBy2mq/IKjs
//nLEwnz0d/j2GDcQovie3u6gKOlEwSMOqz9PBYQfQriHPYyphINvHRfnXHWDUdEMGUBb7WqsbsQ
jPBbkbQSwfju6c1kwe+LCErpGJJ6Ij0fm5ZSmjrL3uyxZKR15GLHg8uLysyEWLFA7Sp15qaVBAFd
GWNgSVBBqiufzjLngOBKT3v26jXofsONOkElXPxlB1vyHWIYODr1fDCQKfT5xQTEgliYzdpTGMwq
dZ6K9/39nDc9+0xjUVaSywBplblUFvkQ8kgQsPLp6bd2IKar1KNmZ+8ljzlT7daVpRMmwQv5s+T7
7TRpG/Zu6VDWHeXYZZtblgdrjKS5Khsl1KCHYgF5NCFx7xOApI9QFYPlxMdd8FHWfYkzOX8C+XGo
KaMmimomZvlA+RP0P2FrBguICbmqIDV0aU7BUWyiTdWkyN4RIN5pMn6CUlifMJM7G//vnU/Bi1jn
Z7/2wMMubTPAILn9edPCIY/5Yq4feKuhmaq97bPGpp0JnaZCf3n2jUoLhQQBnXBN31cc0U1IsBez
7mH+LxvEz1y2G9QGr2ZzQi2uxDuvwgWDSEdPDSpYc2BlyI/wnVk3UEHMwG5jZ7j2TdWuXow+uaxO
dk2m7yy7awvJGmLGT/xILI7j6S5nlXg0lZlhPbhXylO2rAg5aJZQNmlonTsvV3qCYDLE7JNtC5iJ
wQXRvIrAr4s1/XCEIhQqEQ3w5gP5C2OpAKZMnVsJjgiI4Z1PiE8qNlARrdkbpvfL5Iv7A/S3LCJ0
/HtNsGX+udfNLxEc77QG8qXiY1q1WWmDSqs9hAwWdta4Eqo77dzVHj4LdyfaAPiWjdP4llaw2JTh
GQv9UMT3K7DnMPyz/vNy4ehwtT0p2ryUMRj69AzpOm0HYuXoINNDA4rQ/y1EzKbrJvWmG5O1BAIx
S1Qg6bgSz7qsrd3ZA8WeSD7HN5MqDVLbi+oAobD6dTuOxrJkXAS+BOfBxgwGa/2DVgnFVO8aiuyK
2pxi+VrzFABN0Pa+cjJlnJ7Vu+dAqld6m/ZXZFbMut9TmLopmAP8g5AjMmbSZa9Iyt7Zmcs8leFo
h9hysrG0sv1+1QR4GPSmK0x/e0Pw+V1ODbaAomBuPhztC4GyOxR064kHe6rU8ZUQklGNwTB4T50D
A35czrnH54JpkJKn4UHylSnX7Xz0KlcZkJpQKUqhWOtH0cnNh9LH6jKJNYxnfnVXp34P41+1Lwk2
tMEfLcaf5yp2Xq9QvLAJmxlmVSi1ehLJ4SE6V/3SAfFc1aSKcJjmFwtNnyucaxybI9aonatJt5E0
HAp5IRoKklAWAADWH5I+Zw+e9smgDIDBe/I8qoSR2AZ14GP8mIKxi7cV0YYKxfmfAZ2htRg7NPCb
5Gl6s5ZlAT4nZVqXQs22wL2yd6Sz9q4afKbZDgWL+RnngQTee/gy0lz/eyTZQjsrhZh2h1d97yEs
oiy0A9gADIMPDwxGFncKq6+Ldg0dbE0zPT+lWP4219MGue+rvGG0+zktuIIgKIluGHz3yPqX2Niu
z4DCwzvZL0VcEoULgJmHQvRZrSiriF8UqF3I9hEGh7pyG4PcUVDsZFySZgKwSMQ6AGRtIJbYsW6U
5kIRBeLyKSjycBe7fT/MjLHuSwtmnuHyqDcSRbYQymnWKkAx/Gj3RuqLssDRyt8r5VddubVYRz4l
ixhfnwoTBxIe3LwA7/Kk3NlOuTXtRzIHh45dZSCyGLrKZVRfZPu0YXJFsItoHP1ay0rBjdA8MAR2
gV68RoJPce9JkwD8aha2znTTfvvmP6tHNbbt/kDV19zvH9Uzh3ivgVIAo4LSEd3jrSlYHVLQBEp/
FD64epO3hq/ynjTyyUr16FBuinpt3N86f4qrxtm4yRG9AXlyls8oKnDLNPBq23SywWO9dg+NoQK+
WPCTN9r2Vvm+mJmFIvy0xpvJSBlXt3zl4Chlsot+nbtfZGQyUGqQgPMiAndZzs1VuLQTLS6hXmwe
oPK5U6tvhpmQBtNtrQbzXChWnpttWdfZmnSGcVveuWf16dxg3RQlvUKVGHQPGPIi3Od0S6X7tD51
3W0qHMcEM3+91RP9qBoaNhX9R/ZOB1FqBoEzQJ5T096To6A/rv5m5ZIIjg3B3eyxrdQ0Jz/UAgJ3
NS6JmGVneFdp7OqmneiSBcDGGyh86l/xvjsjHGWLsCkx6OdBrA65TGvmokewVMJM4EPhDl/DpJwm
zK30wQJQA5ig3zIZ0r3qPImH+VfasdbhzAmmqiGzusUHRS0yxhcOeoG2OZE6vWlPEreu7rV1Db7K
OLRImOI9MoB2drxCYD4XfGdWOH2sB1XKSrCzAcwORwO5E4Y+sEyFFR0N+TCVm4hzh6fWQJjDDn9K
KFGDjcyZnrcf3+pWVI+/TvrNlab44NRRz0bBJoSZinUMjByeFB5/yTUoBeZp4yVdXjZZPmPN7tTN
AL7Cns8qN6Utuyd46obUusVk5Zx0gJc+6QfiCWlh2QcVoZiEC8DxZSdQxzGJS+4Ot1P2P70cR7Eb
5omGxm6NQmL2NYYK5O3xeBRbhkvbDYUrztNz1oII7ESpZzNZ9BZStfkby4ZBeD/hJiXbSmQD7Aj3
fV8BYOezkCKGSaDXO11OKUgWB68sMf+W1INHjTgYqJGlOLgEHTqNbeqQGw45fZvjFKY96ACjulyh
SFBD5w/gTrqGPeAWyWOrmKSZS0YWdUibTmfFTz1YGhGTnt4MbMZbt31O01GL5L2IwQjDzIO01HK3
RuTq6g8h2AUFFyzVApye6M2kt5kkhGlGkaT6RGuLDrsufXuE03VdHibmlj/fX2UYOk6Xlu8luTPt
Gj7aqU60WiyTOMSFWBPhL5YIEA9CPG8EOXkRD3OyR2If3I7spJco6biqubtN3xF1R6S4WxiFlQ2t
Bac68qeZXdqbnFy1e19f5axI83ZOSmFsyX+2JCLuqJzkM1pje3l2GCpmuD0j3rjc+nxfsJpmckTO
Q8L9kWRIqcqXnsu2wy70IAVpnDVBAi6iACIy4zcM5TJG5e/k/H93UdBkNzoZkRVhR9VHneRgpurm
83ciXC3JSVy2wJL6rY/3WjnvWgqRP75yIoPUa8LwgW036D6BnFupyCq4gPlkdJqSRKnEOlLxfLZh
vyXCn7x/4M0vVAJXuuUZzjw0Hw4tC5vHcMxE5K8H7L77az+8QfzIOl7/tzjuwG3Hxx3uAgfv7mhz
jcm/wF0pGdrswpaNyLyA3hs99K4JTDyYWbwgMH8wEsVgKqql71Q4QOGKaCu639sMqjxVNjE0VqJi
9cBQ6hm8fBf2f01L1x10wFz4UnUJHUQ3LuDjq/1utLDmhCL0VWfcmTn4Ij6ldiw7jNbhThYVGEA+
9Ems8q08+NAn05+Qa+H9uW2Hosv5ThbYB6+CcxQlIt3yKtkVH1t1QYvNWnIwwvv3ZNoHsimSZpFj
/ArHFA7GaFHoiuVNynqZGFg8N75lhJoaqHygQGPRvmw2+1ObKmPyswZTudaH1W+Ka12bGXd/1Cmy
DFFD5V0j9wcj3F0Dx4RO27RMkdvl2RVPDyIBetTNrBjN6835bnGWYc3nk+TPHBEPy821XxA/Fbjr
WgUVPFpCAUdeBbpwmh7lBCf0X3KUL1tJJleIAPlhcsZGWGaS7CT/tU90m7r5XwqJShRC+CO/C56S
BCjOC9QtfwK+5qYZm/SIDhWZ/QWIenewe7d7RN6P/uGYvAAP7r5YqZK0UNgqKN/H1952GIoNfxcI
HpINgi0/fHLVQt6ab7JEZz6zk5hzNwTYzmhJk3ClZv+nyPGHIVRKH6wyCa79LXGwvkkQX+WM+o0G
eYvJUv2UHNFUU7nWdsY4ME+FcMKQrA9ZJ/w6erGAnXRdUNrNX6Q1/5JzRBMPVUjBHRCCtZAC+Wht
cGTaQL5nvwAmQChJL9L3n0vy0/Gpdcm3QBKOmjZxRHJVtzZVhjA0uNZY3w7bFW8RrDWV3Rn6bAaU
ZRUD1u68Y0J8u9ftYbfM+MwDV2Zj2HKVqCuGZMa4UiX2ne9L9/KbOUx9iDgPPM4tFIB+jvMxqf3m
suou1j5mlgNFox9rl3XaXnm2c2wcv+Lm+PKylMprgYAC5EzvOgc2/jZMqf2yVoEXYn4A/4owmmmn
UQQRfCfGeTZ6zUa6CobBL+C1R+sMfWOxW4smai9hb38omtc8TJ8CYSr8GHl5JbRA74+hJLm74feb
IbJDcR/65Pc003NRlJMTDIBiM6GKloshC2NTZC9ldUDkvZmjKXwGHXhMUGH1qh0l/r0KYkYPAkmb
FWD5lkKzgE5yN4Yw2XM2DGqB5hYYFsPH+yU+D1qU6YDr7h+Ltv5WYeN6qSNTGpnxocqvlDXRH39x
Nmv+SV7QW5dm8syZm90nEGWf+Ch1O2Dlex0Rcc3Jt0+QuGOjFHp4xRTqKi0oXurHxcipmah3PTIE
3xdsh1awCD2ioT2aqOA6pJfWdfRp9DW2jdTCjoAl5m/UqFuBLUPngvMu1+vHmtkf6O3oheM7wNJf
l2cTf9xv03hu+b+g8yOPieImW/1xKjyFXOzeV/x7Xty5Ud2GNNxbltvQdixPWFtBLqqKBYwynSih
UgtWSiWERhCf8G6BJB0idbHaDVSj/y08Te5DFQ0WOkeZY8AviTsQhNGvU/kFRXuN87f5FuE5BWgA
yidEfwM0HnluQaUr6DR7XoGcDc0xU1bKYMAcat+BPaYT/5i/fJDCg6zqzWFl1k5y8SiXfnT1Bt25
/B8j5j+UKQzT9CiHsCmw4KN09AO3lo9TW/dXBgZj+80SOEbwwse0ho7roX+ZGizaoFfCwm0XKOde
w9cw3beSqK4AjLBPY6WqJLPPRg4t0kczuRO6d5Mc969UkHosr0Yt3w3pVKhdqAx+k8WKd7ouwgsp
2BaP5rX3l+dO67WWAwr98i5Tl8JZnW0QP+Zm9e3zgxkevj1oQ6cE12Ue69PO4jA7A2y83VUQLXhF
ecNT0Jyi5LJDhA6wWRLp8JLHnmFt1jKs0XCITtd8letDVKqwDAesd0D4LyzP8NuiujUd4DfWjeeR
33EHPtsynO3BLcFoRDy+u50P4obkJuh7UesE7X/PrxTZfJoFg/WyzQj5U3wF3dDBsNs7LRhXZcVz
O4xCnp/xwn/7ujv7rgVG2y1+qbT+/kCu0y3DVbtxUrtLUr16Ao1S+l999dfBEH4IrRZ9J4Ofo6JM
LTDJU8RschX0uFvjtTWzgmDDB1y2GMVL4ytf91ybCobKeihmM8UfuTVj6vys8IK37JU9iRmYNljI
UMqYTsqaGCwUx1c/bR3Z/Kn1R4VXaCE8Q3H8+zyvgXQg3YfT9+ZitxWNYpmnWIT9nuhpV37LvUpF
Ds5joaPhilqxfCDCdbmOBJnTMVhyzMMSasjirWDPw407fpEQO8CLsvowhOUykNqZ21c5RLny3vA9
ZWbzA5nm3TZv5646jbi+zsyKjp0vTM6/hmbvSx25pepeeLV43sXZwEgq/2IkwALvqfIwbosFEvhK
6kFRCfankVRHeyXPDKcvbFhblHWLlfC0WbuAn+cdjWVEe6fFBD1iHF2KT/hBIVQolfSXfsUGpIdx
DwSxNoFdRw60mD+9DW7ZSxoyF/QKrN8EcwSeojMMAE1Q8Fz8ngTPXmTIyhmN68RMqDwsjLCiTKqI
l+jK07THmsg3KhWmblrHR3M4xxHtaSxMQ/16uvG2yvnoIHhyXauLLgQMnebfQaAHQjVMoRf1bjEq
ckomZG4jyIPP60iQOKZQi/aBdxQJWhipYib4dBRviloWrMpPbOwA4tX7QspQC8gEbyb0h1vYlsBO
sapzA65kTzfesR4RW+0Q0okJyCRsJMn+bRXZWT2QgoDUwna0B5l995bdnWjRZskeRJ1vzUwU+8EA
CQRuSc6ogFP0utm/mvQjBO8hD53hAyOMYxcZ/75f/93L5hri5rt0yl7nKCJWThGmwkzgwnXKpRoZ
y2bU7tn1YI7/OIVNixYIKAPfPOIPJSxie5JEKoUi+ZhCbQCdfs+jREcDy7ggPZBu1M5FMi4HCLz1
AVw+5q0BiLqEABne+/pXf48zVEVgWCjliDTCJpzFDlUhMFByQ3wqjBBmqsAPAQ1UIzT0oIG5FIsb
R1BpPdzDVrSUB7gQzpUgLFyJXcPfkBypXD2dKnZ0g00yEuuAAtcYFdBBWCNfXwIalah3sWrG/JBs
cvu2Wltc9/DlCIkRzl6xEWrNkfs8OVCKhTqWGzNw6i2Wti6QipSD8zWTNkwg2iGZNXjYxzOcQDmj
4w3LGYSSjFGpdk5i0hZEyi4AEMrVYLVCetkv13Jtdne6Nyj2kCj4YnkbxJaTik5n392Q3cDPYZzk
dK5Ajl+MR1hIs1SRwMWfcyfhaOU6+RBXSMJgzyIgJikTmmUN0Ah6CwcYNEBC2MOU2w4eQ6qex6kx
vilI58O3vROEiGQs7xRYL3rBpMC8w4WzVmqmHXRHLEyDmb2gifhq9Pse1QZooztDtvuFP6X8qvBk
h4V3URqi3ZvupKtfJEv7nGPso1HRFnZl6KOJ4jeJjmOFh9agfAbStVcT1uqZO0CFet+tRljvGj7Y
yOF5XUl9TTlCOlbwJaiuIuG4NiAgbZa1/hy7FUJssSK0cDKv+gv3fF4oYrmbLCJV5svngz8K696Y
UToM9o2J6ucwriOaEpNDmZXTOQaA245aG6hzScPReJ3NQwAzVcg/a3xiVuPYIHHkA/JKXDtzYGey
pn5b8bbZ/mp9hcWnlIcyG0f3atUHxaurtilHAPpejs4gnx5XGseQ5ZrdS3Fi4tZJX8LRF3ZLPb8K
6jrG5HPWchGFnpuARpLlyYUsYBSvwxmFpogkh4BwTUKx7gGCJY6cPvnTIp5HooeXH1z6mglljVfr
lenXnbU5Iq9Ey8tRvr30YUa0ulIw/cJtbgG5ICXRg5pK2zmgISDVaAk2Av8E44KvizVHBsVYv/z0
DIOUOBwpVfIsmEiwKegOtV90meNKAOfFIzoTv9KewtECB2ziXA5yQOk5kPKCHWx3d7Rmf/dzd9Op
PuVHcGOKS96WuwajquRO0UrLbMHNR2S2o8uc2rmwet3OErvHreJxBZ5kkW/MHe20TECKlUnuhmrp
UDpIc8DFqS+5T/WwdMt5td2gpIQim056JNB/Uq4dZYoFdIszfvhyVbFEJwYiIgOx6iE4WIe5IBaD
Ceoy2G+NXkUkf80I04rDHpcl86rwmRn3TvHw6ZVXfMtG8HAfvCaSrzEm6Hie2YW754zyo5XeWIiH
DMvrm1+BFPcCfyX0bd3gYA+7PWCR/tdlVewkCKny3dwq0dJItaFOMWnd9QdkljdSkLcEjRAbDS/O
5n5lHa18ajhecO9Yw1jwMiQrsEebs44qUoJmymd+vwxe0jF+FTj3LRFknzsGck0sPCTQ/iLUWEA/
jqzSgPoUj/DXu4TlEoD+2W/zml1tOJx4uxTr7DEl/VaS0R048KbbU0LJGIMmET6aWic9Iv4rPsZz
v5yj+zosE4n4u0PlNssTtPnoopHuA1XGOE+dos61tPap15N8+J4wnyfSWChSFWxWAbSFRFpUMo57
rxITT09fyVnHwrQ5oYADhCUx6GVAYuyogaWklnk6dCx5CHxxcL0huO9KOlg2Tn6daBP5TT35ON+A
1T6Y++g1ZbNqy6E93GCs9PdjCYNusKb+1vPalh8/S/iXsiFGM6WnGCgqyEjdR+K0+R3isIeKlYwa
UZz14OjTFfuyZPQHDtO6An1QIH/uNa/XPGFoiZpUgcON9Gh277zm0jxx6ry6RILBS3p7jY3mGHbK
i20ZvPtSEIjOaKwpr8Kj7Y6zYW7KvcTMjdWnAqDKTdeDJ+HywlwElxi5rGQsF1M01XsZ+AjJNCtn
AuLMEtAtKApVBbZBs8WFwBTG74O+TeBRK2Wef/xsYGpEAhU3H4C4WQ0wOmVn6GrsppLbk7XRDSRE
xyLIP7Uh3IEXX4PNlO2styZ9JR70cRMTCe/vNIAORsBKXhPYnMxb+40+0ALTPaEBgAepOiXo9hra
AnhoQqPKaJ7q6Or1aL1WbvJdC74prdnJ8gSuODusTJcp9NiztZ42evATSayEcgggGtvakXdSSNaQ
h+KBBrtpVe+emFzpyzcV5dnlQp2/SQG7VbILuRLZbEXwOtZwgOsuNNIJVZX3jQ1JpCXokqaCA22m
GMaUEtAioWf+/YeoQ09F+vwdRcdPE6u+aw+wuI2toVJM097hAnr7QxwdzPLf5bf2cQquizUYNZRN
J7KfYqb2hKVuvu7ajuorOUtzfCP6fwgQ4//WMHcRd3xnNvlizdiR/+CKc8ENMdTFqie+/et+wShk
5mUvrwCIHwLt2h5zz+BokZR0zZRNv1A5AaZAQR3duvYLzNK4BtAKH3n73gJgaIamgXP8Y6624s54
pq9pIFPpSz4JW+HM3HBQ8t6LHIRuchVOIJS9eQ1yNneFr+xcsFHEY5XiNLh09PrT8dhKHXUOqzdA
kZruGtUhtw9iyKRP/lleoazrf04Xb8q+GXHNUncqlsgTd+l6G2V3h2a4zUssSP8ZLZdDdkU3wkQT
mk9jEphrvBljf/nJbZHd9EhZ5UNlWoinnMOqMjDngFhulUlqDj8U0XwuHyYgMEj2RLM9inqmO66s
JgRg1DHF73lbJ1j+B5ogIaPHwssIx6iUbJOIU3kge4XGfgL0ZEc/tUZ4bJ/6TJccuq1TtoVk9aJr
tMZAualkhPJ/UABn7aYjEDxVK/eWuU+H0njzkEeNOVv12URJjZuKEvdAtj3J/o4LTV+KoarlX3wc
7UuZ5L5fNr9eWOCTfv/Fh91uFXZ0eeAQ3xsciSneW1dfhJ+9HDW6niuMpjdNVsAFnppB+ywfzH8B
rOK2zNVTpU5U/P080VBuneAczV8BOgvFdzjU8CMTw+XDmHLUx2YGtOkAoC2/zgPyPrrgZaXEyNXk
kQXO44sNhg/3bAQr2cNujKSIjQ30+ViMmq4eaKvdq3kbGxCgPazyNaZPFCIXizZxOhdZSTe8vWIZ
/PUCiQdc9LpZNbbqCum4LxChWbz9bAAsyfk0aAug/PdG3YLRAMqsYKfZkORHB8F6QdkKvvGLaGvx
0l3kmkmduPn/fyiGXljYHe3ehZzhp7OIWpp394X4ZiXcLaKxIulwZFZpOGh4bhisSSBCOCrtVF1O
Qi2rYuTyc0pYla8/HT9kWfPw668tWZV0Q5NC8E5VTWQUuwtRD66It2xIGBv87twtgP8jKbD+p9jU
EdLAz4AFQOqa0dkYOT0K1xmX0rZxvKUqVTO8AEhoYKKy19cph0yyqAZWak7AjpJ7MsqCVTLh9q7X
z4kPTr6TvxecvAs+iiCicgJf+Eo3Y1vjvPu5pjFGVs9bVBGTQzCaRQr5NkkDwbxz7tdFTrWAmYaG
cwFhdi6zQo5Y4PRsdE36GlK47nC2XBXk/0Z9OVh3FXUE1eitbHcLL/tGaLX1DyDOU+w0q6JtoWIr
TqwgMrBVaW25i6PUKp+8QrXDkz27bYbqhOiIbrSNuq6Lk9AKAn7blghGYj3+kurdKE31q4FAbedE
H1EiDXS/rVF6SkntK3/iEbJUUcEhWreREMyveR36TquoYcKTQlK6RsGGPhd5PZ1FcpB/0Ch+A6wo
57vdXTBohVnpc4Otj0zASLP685Ao2gAWglHK8tfCQ4fHjtTKodDlG98EiOFh9IMrP9mNTI8gMxI0
UJ4IECNhGwZsDnCafNCTojAdQp3RYrSAR5TP/zpSw1NyKKWtTq5WQGKJgF5IEHGC3sTdXhW0toR4
+Gg0YUyhMtSmYhaPCj3/lSZlagWoa/5LRVM4zU6bIJxgk++ILwWWq1Nit737Xnxdiwb6Nr+lCMjD
Wmzuc9whQsXYcPzUPPC3W18F3PoK4RAlMSpgFBFA1EFYiJvSJOQVxWVjbrvwiPu1HSZ73XvPEP+i
Ffbag6wlDEFJWJIP/KcPLkukZGqhXnFLT/atfP9cY8d4ftk2poHNxUuK+s5H536JBNfT8oWeyoh2
+CM5Bdly7reCIiAgAjhAFPiVm3dhtZfR4Ewj7jOVUfl+yOugMxuXbhDnauLdpc7j7ZyPZJ9NHy/l
EN9J5d+135Y6D76nT6MKodPAf01S5986n9CLwL9E3+sm9ZJCyWHJ7j/a/1XzCZe0wl339GQKsXCH
foWy8aZnv6hRuKiv564II6JvlZ7Y9+4TkAN6kI3T6lyo5eT3SAjDSjHeNgHmkAAA1fzPNKW4SzI7
Yiz47cMjkYvPGdFFSSvpnCNHFm7SK9BFBkcAExRrJbasjemB7syuUzncvvy1CN9f7JXn/Wnr4FaK
BmtH1q/wljOgOKVHASiQxPVGPvati8sJBbY3VcHzmGGJFAt7/BMIjBhmadeTuTqatFMDyRMmaSUu
AoHEHDyCVMvZhHJdPo8w+WIX2tjB7eUhtT8Wnl10/pu1Jd0260PhdyeGiu5k0BGn9UG8eFtBQT3y
5NNJWBN9IFsRrGXq0Gz/e+dUQVborK97Zlc6R2hPcjfhI3OUCGjeYXQBzQoqC+k3MnUsqj6A+8VS
0urq54EQu0R5cvHy1f5tSRBmKgmEP5KXffQr6MVriBxWBi7lkKP0btNK6GPLoXhVFGdZHYExYlQ7
aHgo5ctCu9+1KGMkevrxvtJ2OR/JGlAp3iotsg8hL9noL4iU0AzBG26s1bxNNSMWZkrX+qN5oMIX
WP8HSZdwZ7Okq02LubnXcbXYkv5wNEpcoIb/kOFgAs0usi6uDlV0j1bOpVRZqAJJmvZPAWfdo6+g
0iEWAVPks0a1TOm/j8Q2fEW0LnhQwDZl6a5bXRCUyFTURWCg/SoE4qnaojidqKdnvdr+pu6y/hrn
htLvwbK6NXxVidjsrWW9DaoDdEfANb+xevdqMawBbCBTGK4xABeI6X/w+b3CPIxX+GwE82KdcfZS
8RTcDYpFuJ5jdwbYPIFaaoyKG9jXzeRyFSwqALaKAYSpUSqP6uGoOtHGGlFJMPCU3T4G3XEndty5
jQkAz8v1x+Y5Sr7+J9jiMxOuymSx3cCKObSe/h8LcpvCD0T5IA/loNML8u0qgTe7vCdWB1tSoFXu
6xOYh2w+rbUtEngSMvWVUbb1VPkwDafz4upChLj2kRHreE1FX7WiGYD3mL0THMpO+uI7VF7WrreX
tSkI4W+R1K7R6wUKqeuu8oCapKITi4Sx7kx8n3Nkd/VUQ993lyb4W5pu5beOG569WlK2TbVSksZ4
SBQACkXCFqBWRkye2rQ0MEx5GPhcMo2k7TfFXzFnnxfASQ5759vbX9kfvBJYpCmJFlokjj9Yqxe4
39/RlLWnhmONvXG77+OPaNziSJ600FaQgj3OYPDTIcruVusQoMfGDPTauAE1HOljervQUUvjk0AR
wPhAEbudsJBjlKz1n+clNdsORAWHJmN5dg0wxij692kQT+ey1tUxFx0ecvB5jodAkhjt/XZtOepd
jyS6lc3Hazh/ErXtvGw8PUBNOt941DPJ2EDtuJuj2xKy5d9FI6HtyO7rd5FSoTi1bzYJTQLc6FSd
49fnyK5H/+jEsMu6ZqqNB8N93iiJZDWDGPfBj2lAVPz2w5cAp6xNs8dhPx71kN+yLfPP+5HfOUov
MC0S13ADgbZb2zubGfsZ89siSwnQIQOOtgjKrIcH4k66PumeLku4bbt3u+xG6FwVPxL37rK/U9Dr
d+JvTiL0qENF+QD5J8G6wGsjAvCldMOtCv3djEnsYgtuo8W3PJ3tKq9+SspzV6tQg8X7DHD4P9Mu
H2XGO+rh4AdcqtoNh1qU1MKC/OVSNSAVoAbbt/mvn/TJYQOY28JagZCekjuoMOQ7aa0atfuL8dUw
t5q8NYiHFhPSr3kLxS2U59Z5pFSGhyehyMuVQigUfwRsFaSnxFNhrcdR+Jz6UMJT0CI3HQBcLuJQ
wJr44rm/iXEHWwkOBws7XHQsspIyMmVsmsL2LLh3X9SNDe2LIjl1WVoc6dPZGwWQyZgXZsTwfMK5
rdECLlEehnG229jfW1VvpCgN6ITBjDK7yLQEqQi/X5B5ZCdjWF9AczAItJMRsVFk9MazzAqkICdB
PtCzV+AYJohOLd8nmBwH0TyUiAXl4oHRbdGLtHW4PJkLKYRUYeRC40UNmT9D5xynzi78L4ZBARAw
CAH5Sb8knwPFOzuU2F9ndIsSAyUf9htZPi5Yt/zWxMsLqSLktQnnecjYQRyaCv7cmlvGg9keZrwA
wXVOrFOIEJV0XuRJJb9BZG66WqWh3a5qNLSG7LkXQr2dhiqHIK8luxXHSWeDP4N+BVgdcIAVKY6b
0Jj5UBrfKnzsSTTBP3J4THGOZh9/48hrxCA9oXQvzLkinAiTkgm1BmVHA/bBrJbYsKTT/efoETit
Xbv6Fj1moQjTExdYzNIDeOp61Um74JwqcNTdJr4m0QZcILI9baeFgwaOjfjjrnM6XasoXS6Vd+Wr
lCTh18dDHAM3COl7YKSq+Dws+Ixf2uT6dGE4w46JIqwOur5mzsrQgsXBZef5vGTE4wEjMxjNgueT
GmURTs13935zamvuU68SRVb9VHxSRDvJcy750BqZvm43533ICkx59bJf8S1zL0JSVMk8xmUQRzBD
OIwKe6x18N5I3mJiBm+eIBxJ6K/h2z+F9V0L+wVklchQD/dm/uXDMrLLAbtxSI60pw87KOEGiqSD
UN97agh35iD5OcGnsGRTqVJRWNsObAtK1RrfqE0JduRgdjc1yrF/ukjmYJP2M7V1hYUQp21EfB9z
0RpmhqRDDlRusG4xogBYqDc0WH3oCvq0CI7HJ/RNtByzhUPA25Rz1RJ8no34OKmf5crs/Yuy9F9N
QLvhtrf/UnX21hahBEm5mx9FImmwzJYduUsgy2B4D7KaHaaKdV8OPU7d+shDZIG6KX1LCvuhUlaV
XGAecvsr3i8t2Bbw7y0GdZmXglX3hlMlfHFegO6tVVz+XA9QFXQjULYsr6jxqfj7lQJZnOrqyLjY
W9o/56433iv/r8qDckc3FSZkY4+ZAXHh/2L5rQTqVc/XAFY3xWNdUa7FiVcUjTTRgcn3YAKGDDvW
Wp1SkiQaOto/tfwzxnAN2jwNLj0mY9C2AqzxzUUOG5DGYdcUhXQjWSqH3TmTedftFNgtKf6QBUSa
DXN20X65WUXAYffQM7EutFi21ikLy4BgJKZgpkaNn/ZU0SQ6cS2F5PAVyaEIcBZVQSFT6BZ3wg6W
XL01ctFC873R3L7T0DkjpNxNIV/C8yQBGfhadCY68Vz9Km8X/DSj93lQHGR26djdXg6ixAQZV7dN
lDVLdFQeGWZY5sVQh7c6lINdO51gfp27qDeFj1rt8rQyM75j+WMSQUwzhx3xmxjga0zJuHcV8fa0
TcU3q9qBuHsxX9sIaKTIC0uGrRn9se2AYFHh8kpsFecl0z64bLOuMhYQuBykqPLZRsyxVWkq8+HS
6G71iO+HiRJVGy206C4ZpdpYOyS+d9xGket6WoZ79xLioW/71gjkmNkg187KOsp6MlYbhU6YjYOa
exOdFYyMaogP67x5hmqC0AKRI2i+go/ZKR6/2YxnLUvnpfmazeX/SKp8V/ulYY6Rj+xvAPli4igq
PfJ33FOJoOQA7yuAGOAnDUX+MFb0B7aPjWRtbLXY7pAiYdPe19fni4ZCQ+5cvb8F7GuQJJ+DwBj5
bLXOBVj7Y8QI7L06bHSJQyzEjpXS2YvatZzbib6Vai508oj2tMoAqlTDHo/CcflxVMWG3XvBQqFn
SwlPkv21fbbeUtKHLZq+oO1EyqyeUux8UKbGsRlUzXrae0fhEkBjqBqNffEFDmkmovKTtKhJdpF+
j1BZTGcG3ij0Iy3uVthzSMSv1/f9hpTYnE9dHu70np/BCkFwVEoehLffgWJpUje1k+Mp4endhj2s
Mmz0KGQUrszMDxMyjcebLPimJAZBTnJFZcBj+P3mq5Tbe9jeDVT3p7xwxaqooUs0A0RdxCzPKRE3
S0yYPnZNBZ7EnEZMidINnnduc81Jd4uX4xD6YL6AQV7GUNut9dL8vpsDHNA5K8a8z9W8TXW4M3qs
+j6BKAP/EtiFe9F0ksz9+9rCpf/1/cF5LcpuMXP8S1NLNfcWiqQDPnIogq/sscHKZrMsr73DMi1s
oyf2Kj2haHf4X2duQWQgiTQCEKOY1PkjR6XWiYhigCS6v8pecrYg9UDsZX9BOO04EsR2TEQ03afO
SZPC//yeDlWdIRVe45uxwAmmvl41g9ilfxIscj9yCjQYfIvt7L5Hsuo6b7PU8EvBv8f+IaarIZhb
C46hgFgW49JEyOvT2kQKiVW9eMNnxSEalvRlzNbGia6Ypvf9peOGK0d8GLwUvZqoN4/fQi8dedBY
QxaEcv79XcwqBFfZuCXX3ubmexShqSHC9Nl7Tc0tlf9bxB8HqQXkWhRt+per5pF6O52cHwXcqxGj
ZST8Y/s5W4vRPbA3Gjy9yeAvpq2TbqKG5ddXf3NVkXi3/qyvB3YKfaVMQQmj/rZ6fG/mwvpYLiSa
nu9wDORxEV7H8cO9YYrI0HCB0FmmNy1XK03sVALtfuhk1jlkXhJRb9WbXpAbrW4KA2EGd9dBlfki
kr5aLUF+kuB9fmQeYnu1bdcf5ZyJX2o+17joXc1eWNMxV3jlMLGfHfppXQbwFbALQptD4H1kuhRt
8qrx+DN4mi50vqNBiygnd1O/sBYPPUVW0qmBDXEe7KzNZQSZdgPTu4kOZH3l+D1b8X/YYLJCj+VQ
1ZjpITb77Nz6ljeQYeMLWDHE0f/bJXh0KCmLTZHX4+F42vkedvbiWFzRKKWYQVQpOItYoN6Z5CVr
k0TLScb2wP3ZKcekhKkUiFcF/9++n1us4oEDolzguspVAu4Pg24enLXNi81qVXV3zvVH22csxNnI
wLp/mEwm2/CqMyw1okG1ymgDCdL0iKpCplsGjuy+Tx8a95O2VhS0WMRYq3b5dBoVeaeBSWy7EdeT
1r2/qXrJNplG1XyVlBWhKpAq2BtPK10Q9ePXnxMMsNE+tJdYAPJsKYsCrcAv2K0+5zfVDcc6WkcI
a4GHRXmKCGfnTkXh09AXkDrGaj5YB4ky+C/CdKIz+vS33OTLzzC/hZr7HSeXviz9gIiKWokx1crJ
HLmQl1DSuyewraTTwwCDQC0Rv1yUPMBMSsPCnQpkoAfHW3tdZH97zwYdMODvWzP7DaVpn5gQEl30
yvuzIp6OMNgFitatbwT003Pgbs3dJpl3vGMELFwEH7W8GqwlfSH1VkFwDA8REbubWbJBrLhZRMDf
jYEnx2sd7NW8LebWoreJiHXqudYs7n80JNHeHY0YheF6zmGDaYUoVreBwBjOzpYsY8/B7FP2Biub
luzKwSrepX1AC7pDPWXerF+Z9BuJSaes+8/1Iv94dGrdU8w1HAa/A5UNr6HVjcu9vfJW2e7QWr6Z
I4YkvOIB/zEvZ+T79XBdMBxwnAMnK9Tit7nRuoPsYLqCHK2gudrcfrrFmNsS9ggLDSpCrEzFvFCs
F6mYHckLin91RiPgc6kMXXd+p7H/4FjLQHbqIfSMNi/9RjkEwIc2UyC6T0u/zlDq9moXceDiJX80
gEIvKaEdh2i3I/DfKfhfJQ9nMT4Fbn1x6BWlgUeGjrZFYCoZhesH73naFxxLUSTG4i2L3/cx3+HT
lZheqzq7bHciY5oZXHIwt9SJIqU2+uoBOziXHTTqCRKEpxHMIrCVDAD9/cRjlAn1hBTdkhyfZxha
aoKlaNKZ4GwtFmJs87skhHoGWj9EMM++0ZopyhsYwDIAuU0pjlN9+ZenYpmxeT0/JKuxyk9DpH+x
r7YwLTzBEXJxLO/BHsCWNRn5JAIepb7hzhlW1NJp6x68c4k1LFL5fgvdwVsH7S8/OlzwRsI6guvP
qV9mQkgDZ7IxyEmm7twN4l2n6/E5h5Qf2H9O0g+NG+Cgt7juPAnU+hIaEx/KvWWoZebMmvO6vFZB
1EZ2oXREMtUCJN382SOGqxDWK8jw7YmHt+QbRv8qf1yhtDXXpDC/U2SP6tySbvHdpBXE7aKMHw6G
4DGCnZu7jaV2HBkPmPF7EHECIclXJJ0bfBrbl2Q7zLIJXlz11M5OWBHLg2NmYwgd82iUI5/YBcGe
CEkNfogOjNHxFvIIXHNBh8rKwjgcBE+B9anYzaUoSaH1PPp2bb56y48WgJm69a6mHeGo6rocd/PC
/ISOX/1Ogx/5jYSdyjZT42MfRRZdUzErkeRdf9ZKu4r0aFnf4DpPNbzOZH6wwn+TVu3rWlf79WBN
FDMUSrCYr4NKOhZFuQ/xGB1VILe8mP/Ov8qj/W4lo0lsFEogAHr6v2wMXtGU82D6pYN4FzoDdCCj
D1aDUrUjbvqoBVLS3rE5hwCagphF0hR/2VFhsAnldfzt/cRUIWRA0g3b3UYpjoWlGinTs7E7+QXX
2YmZ3lxi4FIu5k1deJdP5TqluWJUTN6YTMJB3c535giXcmAH6vIWjTBT/XXw0v3YkzjdTnTQ1MdE
V4AX7RyXt5FYMrlY1J0iJ/J/j2DJVbsolQkSjQvB3/Vlh3RhufelvHZtWuurEYsnH0Fk3G6t/+HH
v7HQ6xuxZTpOkltdzF+QNBMBoVAmI3eFL3QUHMzGKucWfiTOLXJ0jV6Xzn9mH+4upuMZCdkQwb2b
nuFpyNdnvbhYdYYw3JMqEqdUgpPtW+gMw0zmRpQdf7KXNLak/Ie4ivrZKMyo8rZYbzRePm0mu5Iq
jLwvRuM8QodI6qFfz7e0kcUR55HU13vcy4Y4XdbVr4zbdhA8nZFM8IHrR+qw5CmpCDjhBuS4J9G+
fESLYQvWB5LguTuD5jRtLSORles78vi60cjY2ub/OsaChh8AQCzI5VFX30FtSWjl4aAWTZon+4Rd
LTfXHCfS2gpxXbcl1GTQYo5j/UKYBC1IeebD7PXAMHCUFpHeAQcJjEobvunYBZsoFz0iY1rcLtpy
LBIhlsosrUTsJIrj2e9IesNl3ctE41fRpDB0OGhiJZb78XdxxnFu8xx0yCxbuomh8HeplAgwZHR1
tLlv09Eq+Y3c3+m+RipxXhaCgzwtY6xW2envp3aQ6wEENOVYaBtAXg/MQEMXSbXnWOWzIOcMmYIr
17GgyDRNFoTU2EH7KcA7M6rN8DZcg6bPDupLreynOT8MldhpXz6P6hhrT0DVoQ6vubEEKQeWvNxb
I/x0tOKNpe8zwUDsK9KIpJMVH1akKZmpmSClNHGTIfTnQyoCn5BFcD0TywXnqmqHybggB9fZZR6r
zQF2LM6MTZtf+mRHHqzHmiV+MctgkVu3SLOKQXyiEiITJiVJ7ASoF5ilolKDis79MVRgGLiqIxqJ
HrzhW5zi9ba/GwnIapO3eIWp+KNmh0A9PMV+d5V7NvAh46Tjshp8aFHuGKfEzNvWqp7YFtpDpAzq
QOa+iogKMRNAHfJgmwvXQqyt67OzBJ/jP1ghSX4miwQWqt2gOG+SNEzAznaC86T7DXVmyA4Xa8/n
TbDGfr27+5Mnuo1iPyFCsL+locC3I7f8CLdFhKUE8oRjrR7eMJZhdC7/CEzmnr3KQFPzMre/f81o
23sTmeHtCQQ8tMSJV9ExYjIMFUOtBwe4E1E/0RjHtsNZ2DdYyx0PCBcScfaDzMLO1T01TfVNLvqu
Mm5AJs+elHul2uITJpJEmSKiKl/lBbMgTXLyIIyh0EqGSrOMr3I2q2XHU5uqjEqK669ZCbw159sN
iBEBaNloeJ7tjaJYxRu77zMCkA17S/9LKHK40ES0+2ycD5JK6TC5clWFswASD8mVQ/ALnwYQ1sd7
h7DljcIA+2HrnrBOXgqKdG0BZsAJfUXE0c7RYWdAGBl4VXXp4Z3oDFY75ezaRVQNg5sYgGyZfx8D
2XV6WAo3s+D29OdZDcwRf9UJzGkmWbmVa+gvgMUU1b+SewPIyOkr3y+TIOWqlwTAvL/oW7xugdzo
LpVu4Bu/l9zqzUq/L/cmAe56Hxl4jPE0j2aiZlZ+BCmAcWXy2gJEuoSCdA9/WesFX/cnpfSX6kCI
1Bz7laefm+Fx3Fy5a4s4+H/KrLcm7W0iet2aBJGnubjeRP9kULBEz3HSPBeOs/Sa0aoImL3VDWFR
aJtT30yK8ycYpZ2vcdLRQJLfjjKO/mTaLWt7ssYdCDtiA6yJEMtS9eyJilYkfWgRwhQ1M/X3zRJp
KNnvZONGj+ZKzHXFdcYKxYg7kSsHnmDODP8BemmWLvk4YVYSL0AcW6HEtVgN6IXc5Nr1FKRHj3Kd
3PwkRQvUrLGQaDGX/3WensBd8bx8K5g4YT6bwfzUpEDeookPA+ELNOg1f+aa0axQN87bIEYUToSt
9pIJoAlGNND8WRnxTHFU65qFfGfwYg4uML7XcPUPoCFnbv8VJBGqA/sm5fH7OhMm2bkS2i30PcHO
cJ0EI9ytUC0AdEhjK9KCEY8YSaz2lB+Dk20SzrwayasvJdZiZDJ+8Mn5kNMzfHS7ZDKnM4yGBh8o
nea5nH9i0gVyfXIofG7wlcwVsfhJqTBISCx7Dyvz5h3Q4/0gzOFmtVVHC/xWSWi0PzQDxe2xMhxV
U8j61QyCpJ+rEaZzGF1kLdYT4JYSenJbi+MRr3OtNGBbYyn0tCStb5S2PcNUwkm6BEGzCX6ewtEO
nSTa65Wt8cO5lUxGY8VN++wuOcoGRkMoKJbQpjwV039EpHSn/iF+xKy78WHbvcUh30NNDMGrLdBV
1Ftk7O8lkX/UeQdQZUCdSetk5/1gU3PUUSajRwsmLF/pOVH279yQwNmLVLci4hqSzdsAuxbOQqd/
otXEeLh5ifD3+MPwV7y6M7KbEZa8fh56Fu6gHsO84Oeow+6NsMQgJ2p3cQ2OwkkD4tqXaGLoA75o
jZ4loN0Pj53Gb2FluiNbrcEvRvUX5Dr6lde0Vx/uBTBZjFId8oTOsz7e/IXt1DknFbkFfSKLs812
C1y8qtjbni5kDll0TZhAyaoU8eWR/W7wp0qNcTQgQAmdpBTVUftFr26g2lgO+Qk1GGcjT+BmpxRp
Ki4WwiVxvybOCTZakx9BBOciBpxFM+phsIt2AqNYoYuDjVcXn0mlZXSAWI6j731gd6i6HyEZpgCe
yucHogg2izqkIKDijPQR6XEsF9vR9EFqhbsCXn7DAkcagIHMyUIVxcS3kLuEyf+lcQkZfhzlewm6
b5kJZPtg033H3plTd23hZR5CP14527HtVmdk/d8IvLvXEqPCf0nVSa4xjkmU5bwDEENAagzWBCK7
w7Drol+PWgcuFXFt9JDe/5/WvX7kYt6LoJCDYwHA+qotkcl6urrj88oRan8GwPRmzvVXWtjRuq97
C+aReJ6rpb6rLRsJPETACZ8IjJ2YqjKtRiA2Za3vlSeyVfeNp1euFLd25eZk/gtHs0yDWPxBhc9g
y2bt8n9eFPS3QFfwSW4+ZjYoezVWQYRPEXVjHtcd3NUQPCuK6ELTJ+z1uUaLm199c+psrlYEKa/X
RvTga3vpFOua8T3r0Iwys6xgpTBs++plP5cnTc0/MD198yesZ92/wgWx9oHrusHItGrYUbqG8nx5
pocjaCboskpbEDwSl3LfH6iuLS18p+EUMFL3PNvdgKChrvwoxmLTAljBSt1ubSrv5hl0qZsI7MgA
nIUi/9WLcRQYJ5Bdu1IZdBKok+hcPZoOM+oJu1NnCwuqXsf42f4MNTzNTgOyqMmYKOPh9FYwvgqx
EWBTFHEVzyl6FWdYIM/YfohxqyR+kaaWq5r8QhKpa0TgJmvvFFJwnrFoCqMk0aXHm9mzyE0fSq1Y
ZjElQiI66FtcJwkWFzhTM6S6Yw4Cw/QSjAW7411/Pd8/fTFW3gKjCUm4CcE84botbBSxttttA2x2
KpjjbZdsoLZe7Lkr2iF6WZP3p+WnbLJvVqxcXIqnpcGZAgF2EmmWKnI/liuKKCp6yLPRlqFtmHxL
Zyy5SCZ4H08GiB2Pku8EIYCRlw8YHp/90gz4/uErSZYTvSIr0t1woXIPjX2wqqwcyLJIjMNp0u+L
t3I6bC/sTU6O3hxKSwW2l+COCuVGiTdiAeOjyRyjjiKR1C4ydbQKj+b6IuNE6b/tI9IiwTMSKAmd
srXY5iqxl3Gb9Rdfd4h4OFPIIrWS1kU7h/LCMBrsaxbxOhz55Cdr9P0wOsAkGSoMKa0F09LrH1/a
0UeVZ4HAvcrH4LboutzMVW4ENK9PEa7FS0BrdZ/vPniuNG6CKoYlCseMQgCKLrweqBHUm9wXT9D9
Sxpx1ggePcNCjUnURkodDlCevAY8FjzCIXwt8i2Xz1mQW6BGYrKCHqi7sn9EAOhdUXy8RUoxa6Pm
R1Tqd+ArQ/68BsUSRgHkA8CjCorw+f+vfJ1h1Srplgu7DI9JcbGDjUy49/X9Z4RcN4+gecY6IAUk
mVnPqYpdgXYi1tPJLaEY00aNHgp+bvJNyolM6hrlTW8/xwWZt2DRweNts8gLS9oxjkKACrIfIhgm
thH4z4Fwz5s/2BaiffzeO71dHWgVMeVMgan9sguhp7WRQEYYqITqYvox+H6jQ8/aUyOahU/nIbjJ
Ldsb5aogBQeDmcXtvI+ZjwX8VN+B3P+GYLZ75pKDdoOKD9OGc0Tz/UhDExJ0w+/ZwOUCCK42iV1U
V+XUmMm8E7OSY0LR/nB0X8kbTljrGbwh0ShU1DhcLOTMg6nnz3vQR3bPGFlvnyn48ii2rfcG81lY
8pE3AoHr8xY/h7vwRpGYvP+i0y+oV4UeEPp1yi9JeXqvJiIvsEnBapkbSjOm3pUiNBicsX7mZRcG
cUacTf+txCr5B4SQ697suewYDf26AwiKpbaw66i/BBjL8mLpTqlymt6UjUcUSigpGnh1Bp6MYwBB
91Qn9I8EO67h9Ks43sURp6qLImpUy1qItjuub7suJleJ5RSuSuxSGvWZ6rsn3cyFaMxXWClYUrWc
LS4ZYafliazMV0ro7YaK03AbyxJvH9v1dOwLjGGN4GtN/YUuixYdAFZb6RYzvu0rvCfLFNHJ76EK
feRcOhEkPgu1ABc3lhjHJBJxhvGvK+8B42KwhNA/PufHHQ4Y98EKhyVqlSeSEeVMHsY0wLsagBlw
pDuI9hVwc2bTemyrpxqnHzTHLfHr7JRqyhfy0eBbY5HBJx3ZH6Kf5kERlOT4WxJcDnzIJLLkTS7q
aJ8WfzA9bqa6Z3/xpRpZgfOIYTuKiSVNpOuYlMu9Dc9MtjZRQDPey9CS9f2aYM77xE54dfHAo8Qi
ej1j3iWN2693ND7W9BYOQFZq9kPsdVsCOVoagzZ5O6/bxs+6SZjCneOehskXdUYVhwLAtsWSjnX3
MmweyZLTjsSj4ESy8TzrM20JyMb3U0Q0Q+Wf6XazIfdPL8bYx97/XUOR07jkAkRpIoyX6PwPlUvF
FS5kw2V1hzqzL+/NdM9KDOGjRvBX/Rdoedoy0BjUv5WuVs7oDkK+y0wI+bdt9PRnQsh2FNkUmCjb
d4GEfgZCqUBwfzdcONFoPH9va5kZaVsEQLn33BPUawEKYKSgwYPKT915UUiBjRk03nz0jy4J4VxB
PYtEQyOrvOi0EyJ772UCfRhidKzQOfB+J69+MHXvrfPAAH/G4JIGx144JLukwqIuXj+X1pMA282J
8aYJUzbIzZk5UDz6QOlusrgtxzzod1cynvhn768+PMgGGMLpGWnF6VstJRnuTfF4O9B2kBVNZWnx
yq4RtFS3JoYE3KtRH6i2o0nPKcQFii65/fqPPpDQBMOs9s4IEbbB2YNchCzbsObjHz0576Cr0Lk1
A1EnT9QJ7pnnFRbGlgy9W05DGjHfhlBvuHi+OEwaqn/WjEgBJpmesTPKbDfg9KHPsm7fqgMysleg
N/nIrzW6275cAGPIYqTLx7geB5MJB8UuAULyFy/JTGLASIWALQffFFaPxdsYk04AkeVVV6Fkn5bZ
zWVmHD6PZBJQrvd53ZPl2HoJwEUSOfjFjVvNq04bwVDmhVs6MZmLuCSRpG+xUvvgecc4F5bVN45z
aqI/bhgDjqhG8LZFMbBc/GRIPJ0CDOee3I4ki9Rt3nviiKjBQHC/7ZxeXrLNn2grE8LVaolRdkIQ
19FXQQQQXDtAroANrqE+KfHR1ij2pFNVXd8nztV6XSLxLJUT4sbjnaWHW5Mlz0GLgSEk+3te1WQ4
bBM6EGw24ux0peYzxABSeyIqO8SClqG5eANVoi1ZHxIrHzPr0x+1u1v+nLq4vBr4o5lz0czoXRyD
zQqKNh9REZAn30QrsjQJT1htCFLKNf4ZODGNxytA9VqF+CWNQHBqI0nMzmV7TnLcBiMjGPDKwQfY
XZB58I62zDK0nz5MDm/rtqWqzCYieCgKqJeoUPjrImQU7hcDQaIk+KltzaReXodsw/PBmW9BryN1
rTqob5XC1EAW/gb8eSyHxd/9y29xmFm2G3ReWL2WuWZP948jOMoQDl4TVmcolzqSn6FWL9rODb+u
IsO4udq2ouU9YcTCfkpVMtqFC857JX36kQXFq1tFh+soMY9D6E3ehgK4BIGi0fP2W+mM8ab9E+c3
YhUyxJX3y5utyl0dckrjH2orT/EpuuawRvogCd7Vrt2ZjmvYVJiIILIleEb9v5UgVI3f4lYcniKD
YeZi7BJaauZrjgSugi7n1byO1ojFJuTfJ4vIk/o7jYUSkEpVDR273xKI88H4p68F6xnsnC5246C8
pLBWhzsY5hRcrpa/YBxt5zZHOP1ZbTjxLpahvgTSMU0QO7GGIQLmIpydsTYV6NkM9FV2LKTlVQfa
ozWus0UskrDlcFE+iM4fB35EDN4LzQyD5QYURLnr3flQSkbuHW6h9zOOw2BW7UQHircNvrOoegGW
OJlq1VjRCq0z8kdLdQX+Bif1SMomQ+fETwwNu7J14GVI6VfFpYZnYmq4o7ISAy+qKLFgdaTdzdiw
i+9/4AvORfs0GSFW2lNGpNZLkHImPhiLpdYN34glQ5WsSmh+jacNGWb8na5h8r4TUk3EhABWnWrZ
sVgm6JHokvNsIy8OtULBMcPsNfw2nakS+ZqOD4gi+7KsmwT3Uc/AVHTWYCwrLZLaFQ5CEDb1GMOf
sLiID3EvyT4+oMwp95CillpQMfyBHu3nuBZCSqSQsP0x1eZ2y+64bg2UchGyj/uT4HVtc8e4Jxoy
oPjlfnhwcDuzwe8i6E68T5k4aORQId7x2Tzd2zQEaV16vNrI/lMYoZNV/bqXUAELQ3lZ3OLi0qg4
XMQnxKhn2Esn9zkK3vBubHcmFXt04aflmq+wl9CgKweaa/rfi5KtlWILqp3fOHDBWpG/ss+nxQgr
/FvU/jFMSS2cEDahVI3tnl+rKwH68fTK7egtLMdjoRxUfp1oWwN4RCNv/aTKw/nhTRIpvXjqY5vG
J2CXE0gPmmDebhSL1LFyQuI6Hofg14h82t4hfCKJgWXQQbAxS3O2fkkfG7dI0i7jj8Ir39V+Waiz
zRSWaQYuwLLcZOSJ/Kl7TboNhiEx6vc468EVV7psKY42wEsM2NHm+xly1kMiJXZfKY/xoRT4gXzN
HNww57g1OlMwL4j0xlkUUFJjz8rcEWfzhZgJ+dMGIR6vDGr+m5n4zPQNZ69g8DZoXRlxw3h0xuAu
8H/0J1vvvCk1cFYvqiMJzcBmzxDa5O6VvJyQRKXizijN7U88m6ygx/OE/V1beb8TmD3wHeDbvRxv
5pc/nQ5vHliCnVa3+wGpBNC1mCsCYMZSrXgFF9zxcsXqSz25RsPDK0SqfkoXfcU6PR6qKyAxjKyG
OG+HB1YhoZFyj6P9YRhUToihZC9yZ7Bqx8sXK4zC2ET+H0vSPkRXyylGKmOtN9NNAxyOsTDaZpmw
GlwF+R2Rr3tZ+OXzmipCBd4WqDi1F7XHlZ/bgwkdJegB5jDyVtTuY4vmGSvsnClxsHwpKxK4u70r
I+39ZvPW6gWx+8TVJP1WTNDV9EAABycvm4ywU/IRAGBlqtAZeyz12a+lhNFaefQkZmrJr0OiOJaZ
UCZCHerd91xN9fQ0S7JvHRwx7OkD+Hw0/kqGyu4FAt/kHsZZlxhOps0jizH0YvUA+oYa9gLsWE8l
ftPlAkofKdVlbCetIxeeolpPyapuPinbcMfRJL4paHhkROlRje8tvoHXHLHbLmQh3qd6y5k0gYso
V3B9vPAFamTbFFRf6qjB+DqzlcsloEhpjIJQ7CougqmViUyul6u/zDp0JQXJGucxNDUTms8xatIK
9qtDkTcOIPHnts5tBIhFcQ8+XPg0QbUkPiBqgw9WKz7VoHEH8+pHMx2CDz8vz16VrRHFNGBRdGnc
MuuCWUnVSPbxS3xwogK3FDcv8mJ4ESawStnI5GMLnZL20xql+BRwdGv3QjGeyCJetY7HdyyhKn1B
J5ELLiEWZNTwY78jmcdSjMKLC/1Nt8T2h0dmsX5dMdLNRHvWiVeMH90DoWoEXxfCweKa7V+V1aWr
4U+n/EHDNogv/MlNS5/qG9wIimzecxzr8GYzCgFDIbMetjG9LfSsTmAUsVBeaNxNXH1iwOfWFI0A
8AVrJ61tG32WkpqtSwWZ66mAWpADg2df0Pw05Wt8dPHuK8QVhE5+Hmc7t2b3kOXvqOa01To9jLNy
Ys7vg5xQjmCS+Hifpc00VNBTAdO2u8IDzyAoyhNCOUqtdRRRyVqJ87lEBpongYrYTTRvc5eHsNKB
rP1MGn73MslB4FAGRCWtf3dNuaHw3us18GxLm2paoZiNs0czRuidC5na23gBWqpTHV5t52aQf6bU
nWfpiG0+IvczL4sKg1lomLyDhlM5gIuKi/3/NjRBQJnpLW4YACef20mRCJUCDuDOGJTQaDDU0zWX
5jxUnOgW4m1oGXcbBGShNIPkm4m1aIXgNIBnt/XfxT81nb/VGMnKBE2YdYOoOdTtDyrubg/oa/DJ
m3kJL1hPXENIanmLtIDjBrKMvLBcUkY+OGBFYiMN8a0EYZFP4Fa0URvg3Sjf1jA8Qce6cSZApKFP
YeOADyERodsNEipI7d3Z1vfgyt0bhiv753KE+pkZeUJMs541NxSBMMvUbnmvYghq+9+xwJseDwXE
dcyBnrRNpFqUpscvjtT4e3NvukPyzefBYyVjtoDasBGg4yGtMp3YUu9Nw8yQNgDD8wpbbA1hYpH0
rA5cQBJecftF6PI5/m+KyfTWSVDZTB84DZ0vIwU/WsfJBQrQxmgCx0nHCmLrubdNPB7HM3+fcSIN
vZ4a2BN2bOSLQOXuDXR4MjXfbMaKTuJQrrJXHv+2mpRzjJu8m1BVYM5jk88ThLsF5pmhjwaoVqlD
jf/LD/KHqO0jTSVutZeSZyjHnrfhF/0PfuUd0MQQjJlA4uYvnbgwRSGHaltjpi7YqMjnI6weVgDJ
3pQpfCGPyqSPzZBYcTw2WrDWqMWhAeGwGH9CvfH4gT9bmPQ3HmUHGLTaC8ncHzbon06Am65QI+Co
zV7Elfv81b48HKdn/ZesZcOzFvWsnBKTurwho5vpCFQk6Cyct4NUdoJScITFuNhkOKNMA6uy1pSk
MynB+b6zY/C3OhQdPMpZaQOmg/n5NBfOiIZsa8LwNHOZtaItz0qBU3doLlytFoQ7sJms9ZTyI0KA
YNLeIsoLM6NtTYVAQv9owB7KqzlQ6kYbDPpUIIhCvuFekET504CV4f+P0XTsZj6dkMXKPNb3Ag9k
ZfLCsX6kPmWfi5HI9gK9tvN7KfasbZw4OjYZUlNTyK6JeLcj5CVdY2+3ALujH/z7V7mq2jCHqSYf
Ia/07M+q+7EmT19iIkt04QjSq+mcE/j05EOJRSJms3lfc6DyshBj0Sfri/BVAQwdKiwPrusl4VIC
YGF+VjT5D3JOflw4TXwzld3deJKT/KA/G2NJeXCZoR7xlkO3A02/wHhmcKUVb8caaPjKgtLYP8FA
8VzI76jjgFQAK81PFT4+Pj8H9zFcqP3p4zo3VVNe60NpxcFKrXcAQMOFfe9WElTpmooxzOcVKAPH
z3O+UdwA12SpYoKYBwcDVhaB7Voq0Ibi973yeGBVSBotkq9iasirEh7Nn2VTtzuT2EIifz83TmJp
7US4hzcNdWCfx0Euzp0MBadCWjXvaNv2taQDVVbu7+j64TnEFCWLwcRKSdxMsxwb/xWDXjJF6fBL
Z2aFpnzAg7r59iHxM26cKgpgoajCo8PvjirwYotBNMnlzaVWkyb1k7D31wWyqumuhLJAnG/tf/qa
MIszNOz80e67zCVJKEIO37HS9Llqy+oDrcthkiy7Yu/WZt/WWkRkSF4+bvEa3hOtAPPpOm0KCVN6
Bt/3SW7KhPiuT6hJVJ1NGA/SDRjK9OAoKtSUkMrgR18od/g7vqu6eHyCc8mecbImweB/EqP5DiKm
cNgd2/jNq1g2XOAg8LY6VRiQrkDousf7Svi2l6jsjdu4xdIuGESD9920FKWTdupR3JwbXDw0Krw9
e6yu5LgSZC7MJOWY6H+mTsaLa1Lf4eYfOyoL6HseKZd5G5c0Q5xteRDTwtrrzw0WvsaQVoQhokpH
0Vdf0SG2fv/fPb6XgK9vDfG3do/TwFTXBDm4+7qfos1vGwSReN4vsrR4uXjNAzf5zZ4/hkBILKs3
mn6mOF7ijlRGe1iL66u9BOfec+U6DCsvqL5qqaH8NpRm/gfreotGcFXrASjIUeuKyKgWz5/K/MZa
v1CreZUd9ZeFFV1LV9mo6RxvzxxMc9rRGNHMxK6xPNkGSbkVEacH2KE9DTF56OuoAW1ZJsLOoE5p
TLmgx+Mf12/hml9EBGJ6qWouSAQAuKUHBmA0ScgYE+A/M+ksjLwf0u8/p2UJQzP4y291CjwdJk4q
UQCMG2Moz72pVdIM++GvYdAMceZzYO93Nkm2YSN/o7MQ8t+JFq3G4ULlKO3yoJVYSPg6+2fMV2Dy
gQaQUohPM1gWSp6yhkYTWvXVCsyB3RrL+Bktw14xwvGAYEyHCKlsUryI3Z9U1gJ5EQxuDcNfHM6q
Gf3vhz2lzddDz6cq8UnT6JxrErqGE42pySX0jifDvRMu8zRHZrAjliAdGQuqguGLEKoHVD5m/wmE
AQZEXkcAwgD14RAswf75ohavkIO1fXrsCVyNadKfnSDTBt7ZwIo/ncF2KIwZuTYWt6hSlbQccLam
A9J8c027JDYTETadnHk53NjA9CWYNDfBgLXsp9VcNhBzbCVm65gs+SzCrq0qiy20SJq6ANxQb7kt
rBSW+rVnBYtc+LsadOhFCY9/lhcZXAaAWUhEDH8nRpTNIPbHPCk5a6/1FClJOk0sk4K6LGDwpY2M
/59ap0x4/X6qIlpG0H6T+AG8N8tPAtJTMA16wMlceGWotpG0TNdRY6JjjRW3phIhHTjsRt5KEC1z
suw5inCK4IiS2p4Xwu858tXWDg2WZZ7xAant2ohWWVfnRW5TRyDhq7IMGOI5fLl34HhntjZiC2uN
AZCnkbPVPvKCHGuyAccdG9xHs5EmULXcY9EfOPOLW+PhQuTn9lyK3FO0KAXC6lg17/P87LKPgNAK
Cf5lhMZT0KwP6OWosMV0oHWJyyhio5400V1H11lZ8yhcQ4j6gw6stOdOb1+Kcj2Cr2LYRBZvYp/g
HKWc718qeSUHcaVFaeoFKxvDDtnN4F6LADsmRcL7i9ake18Azn9H5MQ6rAKDDPwnSegkBUwahY0G
JLFQx99uPSgb8TFPDkMu27z8hP2vy0/D/qLCA0tc4DnF8JZnni+lGQrJ/kyoZDbNufblrdp8u9ky
DphhIhh5xhCoVaCUaSDvixNP1dpfAuq/o88hHKrIePS5VjXevbrqIGjeeka+ucAcuGnF5QOSTYnQ
wJrPmIL+6n8GB/VNGEjF3/9jruoLQzMGSgz+BjqG0k/1MfMmuuvhRCdfWYUZW+sjv9rFN+DFoIZr
UV8sApTNCS/egHP5RaJCVvHDF14wxEZlVi31Ge9QpeHa5gseepnRR1/Ebo6l3hQlfgdfqydiwq7p
1Q3QdyIPouyePYZtMSEIUSIGgm2tVMk8S6fIVYiDroINFz+4ZYiKOKLowDOsAMb+q8PVoDD2WMqr
/1mhzKtkH2GpMK50tAE2QxMastWTT47WXt3/GUMbsINCVaNg37BPT/pFIOTjV17DwfFHvpaQmUGi
MRC1OwOV5n4qG4rz6eZeXLIx6mlYL2We7T+9FBpiDdcUK8zZUzprJuFtSnTV2/HgEsRj8zYF2YQT
5kvTJBQslXlXv9BmHMNlEvwaYrpB7O4dpaLQfNMpyWYIP1XYO3e6EwFVj9pM0LyjU6d/+bfF/oJK
XWGVWQRukP7Rki0wj8ydbBgeh6EgPVicgc0aFTBNdf0cy+xRXHGPZCiNFfkGpruYp98/YTo1RGBq
GIXInomVnCRU9lAqxgXKgv7tcI3wPhiJ/y/S5ocXc1OCXQqxuucEPpPxfgqNiLTFqfWmDvMs4DYX
ACsCwtkhXJLgBvzC0bnCiVZHjo8sr81acqVeF1R2ZRDz3Hh47ufqCdspIC8yRapbfKjB9zSuIB7h
flLmgjpsCwG4gPfAhgM+1yupDMQv9sNvyzgMDzSWGlZnjCC6zVOuZZ1VCgq4BggRW7s/PBUKh3jG
H6zpY+/YtDuaGbAh5lWMTO4GlfkEZQ3jmsb71cfhRr8OZ/hVBt5s+3NHzCDJA31kavvrMS5/iOze
P+ttYsu7/oEfwfVew6JpOHSQeckDa7eWKWCnYx+NFJ9YnZjQTHyOo8BQEHnMxkh782DmfUTl//B3
2VvoBMj0yuJ8rUhrF4nzWG6ewmeBQNHml89bBfVGU1Apo9Kpflm5bkK61sawHRbqpIY2dToFpj4N
Fyw38dKSNoE5jBmdl5TfWdcqltzM3HJ6ORH+yacCkFkkb5lQrWq87yVlBhs7thvIJczrh5sN6t5L
GPQuFWmWQLfaFsWr0zDFB7wdE/aXY/Eoswnz1b70TPVcsD4+2/nvJ5IYN0QPiNPCDMFc/e7PPD1E
V7/SusL9RD/7B3CZieoVsCo2Qvy4DGn/43pvwv5kH4wzWYjBhvGa6ENpHn0ycAIQs/EHJVb8JBKC
kE9RTfxCSuniCL2UFa1SGI1NqknwVHLeVFh0J977G44GTIDsAfRWfWCkwaIPkWOT4/t3IC8ke/N3
sqkhKjxpAKGORHiF/U0RhL8shIAThqz3vLTAsi5EK9MMwak4BYR5M7UP+0CJfNI43AjWPNoC9mGa
CfXiByoVIGOl3YKQecXuSMg37px9yLVwDOlqpQFnnDR/e2idivJEZanOVF1qBykUAf/0v46f03pn
SHz3x/GEEdonIqtoJUer5LM++0nUtMZWedkSqns4fDpzHGtpwKDrz5eC8WRiU1Q2k/0Hj9t1g8Ch
+80rymSFfj7A65LqVgmuDjiDhCf2R52us6jhw4zXWk19yxnfKqiza/i9WLd322HdhGvHmQAbAOek
bDwM71fPMMFkOVzPzRMG/y0r0oi2dkuTSMvdqLti+jWuaVRzIBHD6p2NUMgvdY+7hZ9DQtnvoTcx
m8+QSdCFhR7AM0WrvJYIs5kVMjb3d7LvebRdDIds0TZewD4RhwaxWZYF4rZLGF+MC+vwSs5EDmeX
iyJe3J5PWw+qf91M39m7Mkffg4eFjEItyf1hSbx/nEgmZIfJVgfi5HCc1R8FnaghjHGdsc6kQDeV
LsbL9V9wJoKt7U7kN3r/ZIgvNqFDbw9KdR6GBYpbNOaB4UoGMRTLUK9dd9VKDNXmLvFqc6gzlwtR
5UhHPKNr/aZO0+X1qNwgRqAkw7WaA7aR6wgoVCc5wpPjCMqyUykZQ8ZCGBpsAgqhE1P2Pg1oDoKF
Xffw1vnXfVg9fO2O3RNSUFCvmeVtbxu+QPLK6g3Zqb6uBqNwKNQgbbz/2Nahw9xXdNJ9eoWaZKq3
ajEqRhzUlpZZiXO9GyVCTmu2EN8lGTVwJCq6qQRr9zBkKcmylXCEYwwPxTFSZxmrB5ywZbGTfvSg
IfV6rj/WxOsPhJI+MG3/UuwF3GYInLQMWyuGAjNwnyFvmzob/SeNY3XUh/z0ptcQmnzU7dCLgARx
/kxzWyqxzx/vP2174mMycJ67SFhnKPZRopaEaM3smkyICiCMPAWiccE8xK8AHyhlPQWZ5vt0x41m
Lyq5HqRvJm4DGyaIJBVjV9/OcKyLfCCVz7XjpjQhfaxkTwHpfzqBakTvIy6RcQLIYzLw/kkOOKb3
tlAzxowkF1fAgc+nw6BHQuDV6BFD7+B7X/msnmofLQz0cdu3BDgLxTe8KS1TRffJwmHUN7ZJWezx
h04HJtJ1niagfswzwrDY1rQpoWeg3yRhFnL2T3cOc9T3b7ht4Cj8iV0ufp6GlKzgvuOylS1hqK/E
SQKTmaNAkudjWlcRUmggr+le1d7K+RK8eDHcqhKwslEsWQwmuqGunDPDEGFmywO+q7uDSaI4xc/I
tTzECD/HLF6xgeC4L92OEWC6/MeaTDMAYCZkO+YICGq3cyHliKfgCDKaoBD0iinCQqQ35jrSKnZg
hSed+Jevi8ADevFh2vvD8XQ69PTyZ+N9H68uDoSdAx5PXv8/+xXIWoOInftL/NZGF+q8Yd0U/Rds
MAPWxvF4cOnl04qIAXZSlpQIoeHiSbOFIgqsiPbd8vMFPadTnPdGxUPbSfg4N2RsE0VfzptiF0pn
3qxdWEaewluzEbcfRMXHumRXP5tuhFNlXRmgjg1BWR2Age6jILydli9cw+FV2j91EvTvRfZRpV1n
pX+mDj0WjvPUETL39mmiJdXt9nkk2hyqXT9uZvb3dZY7sRRR5EjrkzdJBoLnEC5EPBydC/04qC+k
/cXuntFXJ/uRDsziem+kqphYdJqCugF0fXTJKAodJp3AWXIU76ic6xt7kfdVFlKMWYSeiAkGY2mU
1pn8AJLBZGgUSzDiQ3zPEEMgv0E3LE5QbS/bPRLkb/Bu4VDxehOz4pNENLFQmezBVPcgxnRj5n6L
xIw4La6b3v2sr/+bxdpQ/7M7vgO8cHzcO6NLNn5rKYYrck6NFjAon3KTVMXXcsYsavpz9srMF50b
mkO8YEoXqc3coYY3cYEell8eH5Y5sns9Xtp0rP27+3drEatDzjd8k6wGTXdrdQ8pRr4BtAecBLDK
QXGFcLf/wUMcEw6THa37r6kUwANpko8pG1HlWxDejEf1wFP0cCWQ+0QLzxm4DVJq9uwVjfqJVAX2
qYnZAbDRQp4SDGQMshlRNhhNBA4gVPu98Gqb1cdOC7E64cKY9W1s2xfUlwjWKSto+0UhZukmGETO
Eq4Y6Z63HeJczugq2kQVmbsE8AltOb04CGtJpS32hGkgkKcYWaVdG5eR3f0Y+GUN9hwhdBQ85xL6
YhAg+3cxvE4dwfgNNCqEnnwqDqCyp1WL3DJSvO5WSLjgK8oFDSUgtxrVSd7NmkfChC5xJmi3NHhv
AavlIf0SjtjqsKfH/GAy+CZANq5lii35C/jlNPcdaSw8E/4xfTg8xkz5KCljezFO4TfaeusgOHPO
q2QaQy27cQasLPUMnlB0XlAyDlIZw4ntczw0NJyUIsJEg/doPEXpk40EgCzWMytRsIOuDOacK65v
9WW/bEH0G8b/qMRcS/oP8v8Pr4CYvDlT3VyH9rjqhnm2ppHnW5rNXEwCuBO5HmSJVZEDNrh26oG7
OKjMcBoHTOgM5vlQyqKRyq/FB7JF6Sk4vjXoTZprxI1TTgam48PkKthRLRCTo1r4cseCtv7CL+wp
hvcUbVLog0Qpkkqr4GP9A1UGnMb+nLft42uGPH0Z51AvLCFxs0hHQQeUmgC6RDD6SA+4eu9vgehc
W0AtC6iGfi+NCXUM8eY4yAn9ng==
`pragma protect end_protected
