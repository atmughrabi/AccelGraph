// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aw9b29mL+WJlNWcJ6eeSspDFaqRCafLDS/9nH+juf/EXpVB7JSZheCguJIpA1U0V
D6J4ZxKPqz48Go9hkRzmBA8vYbtXIE64UklACx31zNOKyC1PhXKPm+peDXbLe1/g
1LPRCfg6QT6lyYFrBbxTNUr6zR2nEw7mz71fK6Hzp6Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31808)
2SGsAg+kWIFK+7YhyYVKVjdbKSENZYpIGJ1Qthm0w1MxuPpxFhUV1K8CwZhsGryG
aZUOv62woMrvfw4jAGOT+WDvI2xG9MvjpUjwovcBjScJVEOfVUmeei8K+CJ/A1Dd
RgHIubQ5cVvTC6N57Le0CfaQxm7UBs/If3oN/64AtJGVx/WE679s1N+nKs0i52SS
zSOCqwqjnqufuLCik89l+yzN/jUYdAkTEgV33wcVUhEacrD8RyEmooEIMTXNaZgx
CRsqPQzTU6c1Hmgb64shQAUKkpu+51zJLWP9+44DmseKh5U7G/z6usFW95jXeD3N
eh5o7blgkTSQKs4bNLN+6DZ0lppKZXisZEclo43YBXcF3rbQK2W8/MNcMlk5DqZj
sZ3J7ZGm0lSVPL4rmcZEUHAZ1gv2OVUnweKchkXtaWOvpuTLxw0AWTjGPCUpPA5e
ZehMbEggWlZySvqjsOwF5ORUF3khIJULyLi2nn2+mcKnDRTqolAOo3ugNv+vAf4+
iVDnhBScF8XdTRXFaW8kYfdiBm3dl748VORxf7ivmYqPHq8uRGv2sOCExoCMqukB
Y8TYTDTmy6cCRkQk6Yg+eDxb/uA4aq9BUxi5WUpshM9oEaE1zHgrS8Z1YyLFYdy8
PfzrGNX2jcnb33e4DOdxVv72OfK4Z4q+zBeHTgIGKPsQH9OvW+mm/NuPMYIrPMpF
y2BJ4TcSt9hjU0TmhjCq0OdYUtOCF0uUVzU/A0Ey1q5G6zrB8duC7ZglukTLQQtd
/+NcxeSFY2e35DdIxbDNZEZDcQwtPOOKGmshPmmRLqmmTYHQDeuu7e9fiU0e1Kjk
KKMeLH0UUL4ToxM25lSy1DnhJwph44/TKUm/sy4SUxtO841awAddJOfr3YJ8RvqN
x9q8LvV3A7kzKwGNv5xY2R+hwnwBIKMbPtd3bVSyJveLMncLfpnP/lBPfkCXhzR+
VHz4LMAVFPQnL5WcRIg7/rkWiIt+4Ngc1/sZkp+VpSLnJnFHooDFd0ltFlAUj5hP
e/pLfFqzE0QYKtt1QKylqugbvNkrJave1uBzAhF89J85VmJdvjC5XRXJomcnth/j
8Hr57O3jiNXVmldq6G2xQhLoltcC7slSW2iJq0ZVDiWn9C+mTW+rBZA8o0GnIJEE
Mww57PdeZQ6BcQeFwdfX7ohy6/5eW8wdJuTbd53t/2ocfJiS988sKZOTVfft+Nhq
T5IwXXfI3AYhH0PNMLrJWWHH9KPc5pTHS4NY5CgzT89ukA+3s33HBiE2mXLy6qx7
jOu/uMHzhFQcQwvX6JUnNInKr+BvaED87IsZmeRhL+7nwiRw4G/ULCKi7bt0xjBm
hywB5wrpWD8YvkszvVu7Ea0E8sQEy9l0r0/eeTHUjNoep899U4LC5tZ5AA7CmcVA
qhg0KeH38R4eIOUxpCEmRpge1Dgw6WNK6JMwI3i+blirHLh4N68Pr0JhtBIRBHmG
/d+TVQt+4/zWVFiGOUFsGIR7Akox+awMqQ1WohM8GuJPRKMrKq+NOOUmrrfofRqo
yPd3LEiZLp2+E24RsEo+DUk9WxLOjUJM4p/OKKgJlLE1xcK5F5/ZkWE0Q8UlBy+X
QsstEU2aakPNuP9YAxdmurScIoI3y/pu3mCQSRlCELRjOHUuYRJvvtRpBIaAkKI0
3jfM0wpVekHwoOrvcKdMuvKWc6RX7oiylcR+oyxAJrnnwXJ+E0Du3GAozG80tt8J
tbMW5k+PD9g+R1a2xBv7JRKGMaWGW4aietvQfLwbTTrMyMxYvIfF/IByisdeNcxa
F9zf/g/Pf1bzHdWPUkehOPmaweRpN3uDksr1n4NNEgcdHVSO/BgTDOaQDZ3gXe4K
1pPal/1EYM1ic4Arquu3MqFt6RyiXCC3wXgX6wLMDI1O68MgLkSKrlhCMF9IrW2S
KwX5qV1+VSAgjkZOd5wddg2OQ//Ye7lB0pJ5NGnNo58lXEsuhDZWtd9xJfkxpFx3
+ppMx5qUWSmiwhii3leV0eZLMDrflGd0B6SdOGmR1zaOj5ku70yUKIS46ZfnzOmg
yFfa009s+xNwgrcjd+vWZN0cj2qbJ00C1nBl8oaC+gBknqXckuS0rU33bcb3/3Gr
iccNHo3lBHTzVxHlnmWAzcu4DZLTkUKooq6+vpIS07aQ2GXbxQM7zYF+xafiwrUt
ZYui+Zw78uKNO/dF92gx6aa/uEW4sG+AzB7Y0BZPya2TWeLyUXrkjKGKvjofgdH/
R0rirZrXMN5maPVz6fhTxVR4MLrpMF29X+dFtgGCWCcuWt67313OSo5sxcq24Z76
rt80PUg4YyJ8zn+YLohlUMhbgQ1MBjWdjHDJrofL507cX7w8grFSoXIBwauX82Ow
4qESMw88uxARYKvfQr6VSrvmCgPzsLixFV71rDU9JCVIAnUhDLalpk2Ya+rJOkn7
YnyELgmxhz/qwgvQKa7k+B/u6Y7AdwYGBBD5KzXSR35qQ5wQlkWoBEoBBHUxN3S7
xSCh/nckCdieAzFz8KCvstTNQMUiAbBYLycQbkLAuxhnpFYG1tP+R1Vqt9ZxA0kH
+QqYeN3AcQqm9XDLBL5Bv/w16ZHZXROeV8xXBZOw+x/G+YyQMOabHbLtF1JFNeKK
tgwRujMrS72tjyjIq4E63wt5r4dW5nuTz7BTeJq7GZYAg2LCACt0NvNgk6ZGZ6gb
IMnc7i2NdDhyBLA1hO3q2SlQBlXNs7Ckt/ZUrkSlHypaq5/GdFygYO618/t/P2aL
/aOQskhtIZDdANMVoSEFlmEQ/xAro4jjp/DagOkiD/wtR28+7VK5iGXbWV/Ei5V2
xwvQouyhLkWhJVo1WKFsEVyCqIw357bw2fQI3TtiPA1Jo1LjMFcnpnKC9fKGgjCm
LFLCbYKUvJmYqyoUHP/gayO+pAW9qsjKrR1sn9LdM6XcM2dJoXY8veQ8c+qVVDcN
AMT2DR8qqroHJCbYQlsJ2TlFKQl8HRc8zK5YiEk7a5axEI+NqnKpzCgz7a9wKeQA
M8aiexMrUAwPKbi1fUE6VRUCflSPrIrTvC+1XfWu+mXklvFT2nvXNtfbU4l10rkP
mRwZ+UPqQIjQ6aHuY3tVC2I2c00SVmPkSjSegvj9M3nLXLC3VEiQPFQVoDKP/1/B
qUXf0cVpwD2RnP+08VgWh1C73SYT/AfQiuHtJIl0JAPBQoBsr7C1v7xtmvWtBKlM
xKjAkkMMXf38GDvCOBQE195rxnl2L+r2rOnvS8A0DV+p14zyXu69QrUauxpEEzNB
VI4bFKj44HphGifNFfISNaPOY1DFA4yldfyDB6XN8o6hVbrAWp2t2fNub07dWryP
ReWcI+o0IwPaBzagoLePibYSpNtBw8fey1GDW1GgmZeBz99te082s0nMUtnuOH2z
D3MQMAMdAJFz51NhKaq4Yi7mu7lGIb+IsZexQxqFvmcf5aYo1TubAaY/7KXF86uf
3d/uuBYzphn5fR0jYnBmLjFMvUyUZwxkG48vVNrd3jBZ16W4jz6mnzymgaYLR397
lBks2JdnOz9fG21zYG2dki/sCwdRcaLckol0VioWQ71dkK1mEHqqVnrpVRaVcu/d
9DDrXDP9HzJpctPUC9GyfZB8f9husTraHiMHJVK3W8cpNuHAzP2nPNQuMOEeBGl2
QPbaHafV8UgFIR7A9WexJPeUDf+o75lc2SBibO3MlZCdcGtOd4pBn9pn020cwhEJ
nAnSSRDvJutwNxKHKeKXfQtM4M9ir6exw5ITPg05V2wInVcvJBwbwmyru8OoeMl+
EjmNLFgOGaehT1tC1v8yWGMhwFWbS9PjcCzcB1O/1Npqs/TzjO6Il8EzdaTidXl3
qop9gye3I+VH0fMxlBumWpj8xWUxz5VvGtM/SmUtnr4AWcDOuD9bUUleTGHU6YSK
/Hl97MwJy7qwMMM8Et7LiuFSNR3SsGeO0jp9gETEo9XJhD6U1Nuff1LPiPOXSuyf
7OR/BDIZ8qfzI6zUn39P+kwNa+/uQI6+t9JACIzuKv9EgrTLWtnqONGW1fk5+ehn
MKv+cm/HaaLQQk31WMr+GtdSrZbAYgz3w/dnswUNKnncv/7RjvYMu2mf+lqnGhKk
xCmXHAH5OkhzuPN8n1nqqNfJ7Z3MXcKjoDj3hNO347Km2M2ZNqk0C7m/BUEqdEQ3
6MVrPDZPLq6bMDdz+RtESWdLl/neA1nqBfuYmXN/IsSu++Np9UqAbE6nqIRuEKeU
IwQz5iEWam2zaaTpjII42NsgQmzvpBC+i7+Z1QPQeJ+sRR6Ed5VnWiAnev2fvXYG
3uKOdERaEtcLzho5RFcPXSWYcik9aZ2e5exusrYRjn54MWABjcEK9TMlXM04YUnp
GEyYvsPxDcJ02qTw4fjKC5rWhEomrgwkjD4fU0+we7MsA/pGLIjyDzvNIE5m4Xif
gdp/IVyQErvfGzOlcYjAvGKWvouXoeA+f3aH+A2IbOC6DxcWYXB3iKrKpFl84LJu
HyPrEqumNnMXBh+PXHeZDZG5qG4owArUgWofgQePXpdJa1WnNMdUwoPcZHJUTmMn
NXVTT8YLXTE1CICO/2jameGSuhk4yzKu5sdCXHIkonnbjFTTXixYeDKnRmrVg57L
JGE9L7LGR7ZyQM6rHG0xlmghYznyCAc1tyI4c1I7IaVOFRI71NQbMLKjxve9vXh4
5lVKf0pr/gVjasdP5WM630WUgzXxs+DY76+3NBbOSt7p1sW9OPae5rrM+Hj7uldt
O33m3condF/NG6vYS3Z9HCB730g9sRd96PqJQfE3i1k4/IlJhUvaJhnV6puPQzEH
nzC59a9SHO4TZSF18JOt6plxcSxXjFpPxSC6sGH4cgRZuVwTtuvdcdemBX2HISsN
Rd8S15cZgSYlCx4bNvxZc1HQAHJgq2FjBEbFU+ihaHSlhMGfJpswZjFJyDXCdO4o
5qLmsylQsb8CDsdCLmzpZYi/NiuSWaeU2TolzMtYFPGSzA/gCd5O7095sONtNTxr
w+3G9NTAALm5r7KZnIUhqRG1wE339tYZQDOqynD5aol6kLkuiZCZlFEhbmoug+zF
UTOdMdj0bGD+yLbFKv3pXMTMUH3dueDew5nokTxvK69AP2Lt52aVEwQ35ns/2i3Q
YDOMTw2q/JDcTdmHRzj2ROqjNdXeCKs0BRjfOaEakJGMJSW3Yxrjqcg+7T90PcU+
pDfX1zhTfodhpb1Ygfy8z5Q8Tz8gt4X3aSiqVMFpaKd4rwgDtCwKzcHxPmxel/lm
AWBVR4Dvgk+Uyt8rQiuzGs6fiuDH5fsbRq2p7GYe2LpEB6BPvPaBagxT4AZV0jX3
/OWc3bf39ti27Kuken7pQsw8NX89XNDSOg793P/YGxryeS4pmYddpTdJet4f+OFU
Asn2b0sPfcncGmUgjN6nsTSOhGLgXbdBNi1Wur+qnJHX4dyzXUpr/w6PXAC8cal5
3715xrt9MMFxODMmje8wT279elzS840KQlFSUE4Prqev7NXIJJaE6YnPawyWZH2p
ecbRrJm96r2n2Vk4SrezbGYJi1iUbS6Lkpicik4TMbsudt3TGEFevC7ceDV/1o72
l77jIVDRnjn/Ml4DlFvFMfVhot1Ldorqh8WZLUdQ8Ial8PUSYHQKlzD6wYVoR13Z
axuBQhXI59bYM0zJ+3tfRWctJUpZp0s3WIX3bSi+J3ls+XZmF+1xrSzyKoPSCvUL
ZZo7kp21t1HytgN+3Yc32/TGz0pjjb3xFc5LOlzB3jbp+e7dnRQ+UTlo3Adr/6IV
0ReLvl503+Gb80DYOoNrLapFlFVXpmp56NDF5AxHYEBDFX2c6PrQGEeeiYMn2d6O
rWj/yU+GDBAH5LDUFxJ9iMYHyNZGjIykbSEnRYYpm752WckwH7QUmBi0z9T/XhDz
rvFwILWlpvEUuKW3JpEAYUenkVl93ayzHgxq6IeYLajnPX2hhekkdtyEzVnHQl9B
EaLqaRueC67qe4tKCVRIjMThOeFUq13aUUwronQ6DqQTEkp+HSYpArBqSoQ6wgHQ
LcMljSnoSedqeEEAh5T3cii7GvDdnWLBjEc4G8GROpoiY/k0xTAED4OwHTXaOiTI
ck4dusztmrXuDp/AMlgh3ekeTHECjfzIYpvrf2vKHRDG/xk7McNmnjtulwOyEwBT
+YMaKACT1GtOS1EQB3CVMyfcQx/Aie2EOe0hqt0M1/04+TskneIKlDJ8HmB09xAk
wNFH9rrBmWztzqrErri3Tnr4ApkeRHdWlcvVEV2GGKu9/5pBe9uumpSYRszmJsDc
C687FJPt9+5MZa/l9ZAVXW6CuDhxto2cIW88/ytAhOOl3keAAn3Imh/10r34Nzc8
pfE8xSkiOQicItFMcj7DCpY9+ztpAbyK66RQBfbyq3PxdD+W1ZM6Psk+pK80WAKh
4EJCwD1/d1ur8j4MOk5kwUjbkB2AUi05clegXd8umoA1dfjySgs3NmetFj36pbFR
5bbCgXV3ePRoBIjfCjvUBO8175T/D60WkEv5pPh+mrzqVOeTmylCSAHVTKphyVLh
1ku2FDpPK3HklbHtjnJv/bdeTbnFXPWITUxJoQBnI7/x2UN12YgZ8zy68NqYqg/M
RLYA3aCYAa+qBO5xROlM9X5yyF4HMyxUxeFzQHC/5ztDI7rhij2saLMAQ0Xr4Pws
G0L+FXmoclU1LI/UkHKByV/WDPfcft05vnIe9YcMnqSgyYhKslVLN+jDLakFGfrH
8x43QOL1gXsiqZKW/+rZW+v+YG1oNBmRcsInAPAc6loLpXHui9ePwHT+Td9ksAkt
htQJ1hytOjm1s7iWrUSXWXZdZ/1SwtybgntigXoUIeTlO0rnF12/uEXJLdN4lIWE
b/5TaJhCQFsgg9i2KRsWLBzUTs2SS5Ayq+siTfBQIdHiCmtJM6zgzOBFh/oHVHpe
AxEJb6Ys6ABTzo5/Ua+IU6gipIDmtmihGlOU67Auc+ikWfRrlCjb+2NqLznNFu16
8mhAEjksQJ04RH1cwTZ4DllGDIxuOZYMwa+LK/kzwJ4owqpw39vFm0A4/XBXS3rb
VvBvLi4q3H1jKHtDC/yIsuGbzCFB30l8VQ/HvEW5ceHDarbu0hyWry5FzK5fQXsk
UYl+Va/6mMBIZTDQ4gaD+kVLqb/TqFSeU3YFUJho59TGqZMH29+ZYAepLJjEKLXH
u7LiJevTRfwoIB0axlzljWBGYBh991FRf3bpbJ4iOxgCTdcYvCjnOQvci9oTZfjm
55aZzXiureFz/tgYO/HJUpC0wKCFf4yiZtTcWPSqlTOsk7mAuQrN9hwmF2KNXzG7
55A1JpWR0mX3MGK70Hitb3NXkaOe+ioGNKKhPeQzwaTDk80JBCcS9r3r51rg2/OO
SZcAM+AgauEA+7CHgKiXkbQ/JjlDZa9PrzjQEJtX8M8/8y0ak/dTpl6iCmfhqItX
eOT38HA05xMypirlahNXBPUpV1CsHdRgBCkE9qGu5txeS708Rl5D5wNRhcJuCR7O
cKBc3woXgEj5n2+8PafY+TQYtob5T1L14t79OBPp4+KvQQg0z900KPQsYaM3JElm
XSUra4mDU0V0l4nEZQJqG6ehxOOJTK7itLWUp0ISIOsMFjYU+zF/AI31X0qwlj0/
Eb3sQZITAro/3dX0fWMl6TX4PB/2tuQjfxjBGv3eNgPbEufhh9sd0vNhsIKtUFUB
CVsAaorMI/JWs3eJZHp4ql2V6XPv4/xzhYI5A+xN5W6Mu09g+TooJPHCYXTumK71
Jw9zPUYeV6TreJ82dT6eJo4d/+wgy/CXzNPh/unSLyfbeHWzT3J0B0q9W4WpkLb/
VIAiuD6u+32i0BpYweQuz+SxWtceNN3T8CosBcmZK61gDCtvLkDwH7OQ75+v/oya
iiWlvqm2iXQNen5zd8g/kq90AIpsEW4i2yzrz8y3Xlu+0LvLoh4I4csQY7bCB3da
qZR14RYd0M1uv8K4cEZ1+vwtLouSXYdKIlyNIvhUMYQKLvdFyHvSvXGBqQJqdvk2
Is4e0NzeHUphfvuUzIrG7pPtoFNuBZHp0M8Xh9+8GsM4SB5K3FVIwO1k+n7Zv+TL
VEPTDn6us1qH2tWFSLdE1lItp9wl//WwDD1L8oir5qq00MXAzPNdcSyfSV5U0HNk
jljb7J0GsGPYYn6Je+w6WRFQGbki8x23vxScwrEjAP1/bLkxZo1b7ANKS56ERvBT
aLX1wvFMvySWLfl8b7sMACfBb/dHbwVLOwl1QkC4vxbKtGNCUGuj+37oXL7mGQS/
9/Ch7KGWxaB9WjP3z2tQMnPdIFPUuYg1FtEbTKNt1Jh2hQjsKUgi8/U7jWD2fQQM
Ci7UAH7zueD26YlMY+0b+2OzTsUB3popHyaWtjBnxJ/WwjRDCbldhI58YfEzRqfq
Wby2SrdHuf9LGGNSFVX3vbrazsxanOfFOzVMiZuEB/Qsl3QTm9F7UMySyZqKJ0/s
5YIMpoxThbRK95mYtkF7uxZ3uIhCjfDJQUcUYzglvKt9Zou/ZZagoFEflFZ7yYOA
7U79qX2BOtcOPzDi0oqyqms8mcRvpSXphf5n2ADrIxodRtQhPZRYPa2YRSzUrG9l
KZFWXViIYXEhK+v+ObofPXYIWSCudo1Hq5bRiX6tGKgkFRpDFnBxL5B3fA91Xqoq
aoqN5Cq9KHMTTNSoYqUL4wxHMTLiXTekbtKhyV9mjeUMoUwEh2f2AbTw/ZgRpCHI
iNc3SCUkRQS3tc9obLXH8+1FCTNT1jxb2Mu3xjlNSzQWP/ep0zHToIIoeqj5JyUs
X5cdqDpqJ9ETtY/QwX0DXdqFa+Wj9V0yrSLdAxo10cjjRodvqpHEwbBO8to4HPQK
c6JmC5QCZ3moufoWLoGZOg7ouUS86FV98tzKunVFTKe2gUm2MGcLK4w6XtX0Ydjt
PaZVlx/IOgH6FIKaAqSo4nHyXEzkhrMfuiN1Jll05U5JalTt7EjjWelHEGS+RTg5
qgLsiKlUwH7mbuR1OfyYzbfM/JCWRvNyrRkNxEEVGzFn3lU0OoUNsQp+hRhbiBDS
LoZwi0IrjVHXG+coTw7RgwBa+8f6ZnO5HbJrX9kKex06qf9QTxf9IDvTmUHZdklg
1bygjyhXsYXxPu7Z3LqiB5s1lw4pWfOgUMZ7mc1qAm4BEOdfxec4XC0EExYhFqw+
50byF101VzhFNZ4IIQMwvEo3URVWTcGDF7ihHdz/xXxpW+07hkQakUFYfpA6N5x+
kzqQ8ZxzFivNrWrmB9DFjE6JqDbBmEQFViHTDhqIeoIvFdzrzMmTy1VnknBB2nVg
11F4jXxNQKM2hsb3oIDlwgrxubSAXvYypKuHYUrkeOjtfgLe0bwv41M/o+xk29LX
qIbyJvssmK63rzF2JE4X8plckSwBcmlUQEaedIBzCDGbkUBM6BbI164GbH9gXp7V
rSBFHifNUtqxFFHOmi4bfGKlYuIVf1sS48wYamB6HjM5mg8IWlZLX9raVxofXFDt
Z96ooDtz+cGNx9swcj9E8DcSNESl+EqyG4wohvIgWQolmroOVpt2bkKK/eCK47bo
2RCzTIfDX8n8xuPe6ZFqGuEmtQWNe2UiSHUdDswF0QaBrNjgbiz8PFNsgpn9ZbEE
74leQfVTibCsib7ew2iA24xSEQ9b2HMHjWq+bmu5XlrHbqLvvm3X1e23DHvdfqDd
dXr+xfHpBBGJdL2BFMf5DlEfJXZQtl1bYetZjN64Qz+RF+vd7L1skMDWgdjekWkZ
CIY214KpT9dYn805V6i25gTMOrRgxXANiWvMu+OtqAY+dU0+jWbNWpQtBLXeOIlk
a0YoWfS+vNOQpsNIPUiDkORoJBuUxNCWqH5GNmmAoqbmGW3QIhh/E2EnAOOgkzgX
xrJ9bHo0IqfkwKr+/vz/9Vs/95CpSe3mSixSNT/048k71uzzDjpmDCI7IZqh3Zbc
8z7Rl4vSle3yCYnLvY022tYmodxj2zGKJIcA6M0fl3RJXANaELfsBU+kxSjtjbbo
2qNyYXdJLvA7Uq3Nrpvw9VsRFlKIZbHjjrPRTbCTUkMZY01lYYuc+PfghNykhiUu
Z9h4ZSnq8Wv5SjjQ6+zEVy3DbnjDS+YoF4Kudtv8bvOD+GgpSTCBzaR24EusUOYL
ENcgfaRFY+HlpRNnij/pJ0kOc4ODJCR6DluTU1nBjpMVkgE4VU0d1iDVRvikYGQ9
nKiQEwgVDK3N7EH4sR23O3JZCQvlbgFoXA0YuA9nWr7ZOQWQPHLHTnWPjHNr5giL
apxLZycU7WJAtfb56s4QO9M1F7abyUqRotJ1cfizAAHJppvoTzExk7ipC6u+NC6O
Ge/1NR4m9laM6i1q4L93jhBPAvD2qG3ZIr9gTzrurd5zGznuSqbEyFtvLFGix82s
IFwFp5q9/sy40/aIGTvsTqLXgSPOIcKNdrkUwLmN0uuZxn43SaTgOzutFsFoKAqb
A+oW3s10boeVHPJPnOWcXJwhW4nRywgqZUU207eqdLaNcBhptqzdYCg7p71zxjwp
tKiPSam2K2e6SXGayiQQZKlPAji7jeGaWHQz5ko/vwbu84apOWZu6uakYlsqkMm5
7dNvwXnLDcnO5WvCnIcRg3jukuQmt5XwlE+arbdcNoACLK4EJpqLbvcZ+16II1BU
taDwndkvKXlNmrphehBXDeNhz1doVpTFe0Wb5RLU0SPqJumZQSH5L+aC6d+R3uxN
Sv0rbo/aPDu+NjtqaC8dY136AMIFJBfBos0me/LM367xcYlt23tIJcqM+J40Jt/D
GU2zyi52DCkhu6DMPNS93X0VjCruUy4X075mZ9+daJ50RNvR3ARkSgMDA00aKhYC
CHHnHb2X2Hlp5LTT3X/n1XIk7pcL8IbBrjwvEwxN6W5uGG14ZBVsB19CNvj4rWmn
iEJ2EKjud2f9iW+u5LEryXJ1FQ5UWsNL+s78ifevdCImoZNoH3AVNyN95avyuOn1
SBmGCs9BIY6nRITnKb2aRCWKeeEOJ3nqQGPjJq4fF1nqQwplkaYJWnAjQZGge8YL
55/APH31v5lQWmo7KSNNHq6GaNaTz6BktGBdak7uc0Q8RI77LBP1ODGO2asg+KT6
TyOhFXWOsRUOYA755eKtzH8QzQsv20TqxfBNipGcAHA2tiWwBM57elX5L5YXjCSf
mBikKqCoFNJc5S8SqWJcXgxoeiBv1GYLKE8cw6NjdFdQngh4+ykquJRwM+p+7r9n
le/Gsqzf/oNeQMDZZrJbHTownSqX1pzsWpUpWztYJBqe8i9vTFc6D9CpruZ3e6LM
EiZ+USys6dPoM0XxBKm/KrXTfFNBpqrrUPDkbpxnz11euDiy9CPCrYQ28nDUgrbs
+SN6sgO6GAsSKjWayfcs693SNrZVNIKawRkHbRO0W7kgXz4sDlh8s7zvVirxmar6
TuX0HucGtad28mrtpOfBtSZ/EAdZu8u6bo0DP2ZLVrpW8o3wDOunaQh2dOXxJczQ
Oli5fTqZuMkxFDwoFwZQqtssj1WHndZz/lAy1mBXCLTyZZp898zoiYs5O4JuCaCt
DGgD0LprFaqdkOIeHSOzZ5ug/e25JqFdor4cWDy/2OJ3NqQ4Bda/ck8mewUyAEPI
g9roT8lZBC2qaio+MaLB7od9VMhsF4N5bVAu2bsILv1TXLibbRxPOU8lOferBXCV
7d6fv0ZNXeEMuRlwnJrZb0dWDuaMWhag4kMFhSAY2zEV6YQpxN2NWr0xtJzp7o4Z
GaCi0x2IGeZMytsXDu4wfzIfco/JBhm3OUh7zHegFWuzRjxir0HwLBj4PVz+yJYt
CuoOBNdQIkadmhCc+bU3D5iyPbKsd9KR5jLnKkxz8pet4PM469FTy4HQeHn8GWsf
aKM3GGiworRMi2EYx4Wb6x1U0ei5WTLR3T6n0G7vKJ92IEdBjtmyKjZ6rS6WyvWZ
KWcI5NaKRDs5l9d99ApibZ2xCc56cS6iyoW85b9WrUI8i/spwk6xvoHFqSdtpHp2
r2QntZtSZRYw9FdYpVjtAtrASd7mn7sUj3bAMyyakFmeK0y92I6yhHeIjOigvM4b
mdb7L8UnfmLan/x+Q5cGTBRMw5RlqWlT2ibUnWdfUO4eS9ArFp5WRZUvEue8Y3lo
SAUZB9HSU9U02t6Tu0BdepRt9Ma2DBMRg84E/JJpzuaFcMmEksWmHrNEm1yCYi1e
GnKEBFMQso+PlRdFm0SDZ8UlU7iDHZsq14y6EzN9pQLnkS6RaKmjNKSzrG4xERSz
k2OFdlMlSnvTCnpyTPUE9JXSxir2oDGuTXJg9UNk/7g3Xyq93mqFzuvsNxUiqlgB
WBVvtXbts1X6uHfDuMiRRVvwKfACjvF9DjSjir8wYE6PXOndUMiqFxifx2QvIUb7
4kxo5Ah1AQZkIZmrfku6DX3VqtN1IfnKJs6ANRzvZtdD6XKmt98L5qcVJ/udlFxw
wY6WxPMHQ8CLb47ToWjZan0DWz8++A5KyQt5QsKqVl2caAcLX8LcPbMn/JTzmL+l
VdSqMMAAB0OXDuud2DmRnQdxlsQPqD00IgU21vPvfEalIn03T3E63/t+renwwLNf
ifKZbrLcbLNYB6XQ9DC+H/W60keR2XTF6jpX3mXi/4PB5JXJCZcqi+zVX1DpNhzj
0lkiZhqKjXE0DrKXZ31Pl/k+qgHNllgj443HSxpOyGYZOgrWlH3urEJAFTe2g6VU
4zIRAAV2vglNLGHucjqQG8nSXHKHPCXZnrcEs311dCTgFuVmAL50EIps124KPoiH
WbhQ9QdAs+6itTZaGsXtakftn4NPjJ+dICL/KSQvopPw3jxR2ZpN0SIsPcMDJjgK
eaQFvWdh/0MzEa/O6vbQ3p152gjMbhIZ5/g9xRa34BilpQxZiSKE5yl1qdDAllZ4
5GruSw5S0Yrrq/0wpXdLKv658DFM5Nsf8hm1kQ563JmNh6zmw7FGlEgniUBbwFKI
VBQ4N+QWcYTOyClJO4JGbc1r0VA6zcxwllOIEeJHwhpRYncBYxng8s9paAYgEbfQ
blxUB9PoWo/U/R6H9oW+MsYXUacRu+KuADRmu5/9KRvcSXG2t5ckxvpDtecqNj73
9gCJvSgLmQ8xsOb4LLKQoe5uImSQH75jQn/MqS+1eroVLw63xj1fZ5c8WrgsQJzI
HeLQL+682B6ZX9o8fmefwkAkxJR37fCzwD51CG9P51JoziZXDiGYlfay+IYmWBhz
2suoH6XMzwnRHo8YdeIcE0B1NIbBGpo363uRaYinKfLq4xQNcL44LzWQEJ+lffmC
eBGD36X0q4YXYHBXC03VhzG6D9RTP5YwzIIx8NT2nL6EEI65agNoz494HJYeRAOO
PigV8tsoL3MH7mNeTnMgONnIFWXGXyyZzks6bf/tUl5CyPFPDrAxO1ASVj0bUr+r
6wQi2Sc/WxFygbN22LQ005CsB3D2E1S1l4DA273vwcuy7Cl3VO9+X76JY3a5G+gr
m5RWbVRgs8HSZXzkgxgt1kIAdT+Gs3c6tkk8YFrAU53GATwFs9PKuty6H2ME1LWE
RfheOd398Mbkx4LuNzUFxmsL98wKvXgojl0U8neHATgPdNjTNRDitcMcOfaJL+/z
y7yawJd+Iwwuv0k6eqivCRbWJdsOoJEGXvHxeDA7NIOwmjXvP4/nF2YfRCkIsRfh
8rLQkr5cxCbLYkNGA5LaT1tF4Xm36jzwMr6TmIAqk2yhs1hEQCl/66Tn45M8Nf8O
jaLQwdvz3aO7z42N1mQRbWQg1A7jM7e7v7+Kq+41UiyINqFOJ59Z4HfALY8uFD4x
nQpkWMArA9U6PGKE/v78yetv4vNrWGb4/R3DQlQ/KmIxLGnwj8V3/HAYBj2B9jvS
esJDG3ig+BBfljl+i6Hxte8jnoXd9k3K1tl2RJZP7hehONfDa9BjFl8eWMLLO9NP
GTgM+grzsMqdl0NZuIl4Zw2aTQS62rhqZy8QCz9HI8ZqQymW5qVJzW3SMriI/ta/
Wkrhj4uM61FVPVbWBMupMsm9H/Q1rhgfdTT91o98COki8XdUAMN7DkcNT3ueD+f8
Ved79yBGyN4J18jKOwmjizlRGX0SxehGrLZHj93sQaGWZKJRFlGMKqIOVXqJ28N1
UxBMcSPVp/+cvF/fp0kLD9BJspnIozeYNpZlVLQJyXFfvdX7y78dKLVQTBDPRHCk
n3Sdekb4LNq6ugA+5xKsgmDvQrvh+W65Euuue8MBs6qzzKAt8XS8Xx80xJG1E2ac
TXKGYmcg1+M1wGkJP2j1tsdVJCHZ+afvkOMfgUbOWTMetAwEqWP3KjWeTNI50JQM
vSRGC2InmHA85zZwBL7vv6rw/HXVOEKh679CLbzGGku3I23XurTmiXiHhRNEY7mK
nlqozlrGLr7PjsZL68wM05aE4FrdDDsAgqUhFXmoWuDP8VajYzqUwLMiqU5v0iMG
ZlnbNUkxV0S4S35dnyeoRePn+iWV5ClaeadfzxCFVc4LUnEmhb9sxEWJEOTBL5RE
f02dtYbagUq4d1JyCJZIIKRXTiVHwsRjvgiL/OGvaB55reHW4A2KRJ0mzbLjXuyb
Gna8scK8sbFFB6fcscy8sJJJ44qnHR+i0kOLrmegHi/XIERZbFJ9jbes78zc/wHn
ND0dlfFgTSCabXeu8jK68H11aqPWtmZO0ZspjRzTuaVFO5LXMOh8Xk1MqWMMGpqs
MKsTPu4lg3bX77hS8f48JIYBaQLXQF+4dcMdfwcUz1fkfwk+ELACaX7QCtsq6UK/
wfJKKzsYn3wQ5Jj7iiABxO6sNY5QzQ4QGAALrGRVBrVSXdA96pg6VtLtTaXtQ8tf
jgIgKKwOZhV8t0Vg00NiphrZH8igQk4B4ZTMMslTW+bJVT5g7cGuWy7Se3LNRmEW
ff27Fgd+uHxJHLBwv1M4Y5sXDCcvrIihechOAOqJdOd7lw+6viN0iqJoGw6bRLcM
hJVGvRGoy9zEg6BAfTvMDptvI9cCLl14vXXsPM86142uifG/KLdzft/v+X/J7XI7
olDN54SnlwGojgt0FSaSH3AyCKEgKUTWHpLtswNBLDvSUlDkhw/TFcC7jwX/SCUE
n8x3t1sqkALwuy5NvAxVsyQKBzWCfl2Qhae7frKJBXkfYZQnDwD6poz3lvsSAszs
dkP24f8s1CK40RZLRgeu83via3f2rzGpK27riG4iS+h8WR9AAv7gvWXhnNi79w/u
VYT8ab7HrnWvRdv7HM34nFOoHl8BS0t8F+raJfd/xuuA95W4OVDI9S6R9BImHO2i
YWBfliHQHG/PYqUGv6WCU7g5zLX9JSLmdnjNHrjUK6l8bx4rru0s3HS0ubhDMCZ0
FUDdInNBcHJ0Zl+HZ74OTS6dyaQr+WgI+dfEyW4DHJ86xV1hS6PMqTeRcx0hYeQ+
21/U3eGWGEu1cfIsJhWOv5b7kwIIT6xqE9dE3N1Caneha5vJ2m7y4n7l4H10fk41
L9c0pR3KPVs+4aDNyk5i2nrm8GvoWEDN0BbUmFzVB23wL2D0kSSR/qvCBg7LANKm
3A7umgrC06ZEZJIpdGHLXCmXZdXiYGyyZhO5kqmEqu1mn+nXG+ZhVoFwGTbq7Az2
0t3Xj5oZzi2qCgm2QrZbyPOzmmV1QwpRQ/NcCwSeqUHG42Q++oJS67yieGO8aHOY
CYUlNAApsFdEkXLLC07RuLgdk4N1l/Qoo7uC3uEuYSwUqee2aeJDrGMcEC6dnZSp
dAcGogCabEUe3q3BSKYS+V6Y6CtLK8POnXNGJUy7F37Ns/QY/W+MUGv9/0Gp6S5r
5siGXXzQQ5Iluz6OAZS2vRSJwiFJYu2knh9JBNCoABrXsZ4AlFU3RpHePv3X5l6j
lItRiYd5c4JWdoJBcshOSEuYBsQij/39/zSvbLtnfFNPhrL3jrod0xTY5w2G3UOy
WxWJxr0dIIS4smM6f7rMJCtvweekB4GTHHBzQ3Ntb008cKsaFCza+h6zFbtSCNBH
a03hKfkDedibCOObJXk8UUYSOTFC7WgBJp11VWX5avdTroLD/A63SSgkZ5nndWeG
M2p3BU0eZahEl0fm4+pwz01Cgm7AHrjePrkX8qVeOYWmpJujkLJ/sq7e8DH9+aog
rgZj6Iy4zy6FmZ0ix06vfw+5L3U7EI1ssOW43zZLPsgJIrTgTC1j2tH1mWtoBTZr
yZC3k8k+AUrppvbztXfXrKJ3avxVLYWdDVCxSUIqjTjNF4n4pizMjFeUZXf0+X3v
oH3lh1M3FzLCAwNU+DdNwxpIbouwDmzHA7ek3qt93JiodtX5oj3azNVK5gkrokqb
u19rUIwfjvb7F3/jAYgybNSmplpobanT13AbF9GRmkffhAWRoP8VCa73JhOR8TFS
ogWsfm7mYyRl0hg2rowNacyZOf36WdyLwrPG8UB1Bt+8tGIaH6U+FPKZeXRYW5+/
JXrKufAD1FTL4c3Dxqnwnxk/OkWAGGyTF2Qg8LsuJnTu1CAjOLWFT2XFPpeSWWhz
l7s/EdiBb3yEfU6j77W7WhNwJevWrhsrSRLQz0hYMlm/WsyIMWE46KvGBDmPvNiE
pkj5TSmWju+3oE2TCzV967fyfqCoxS0kC3WYy954LETD+xQJPTg8aHtJ3+kTdq3A
p+gwTaFGeWw7/hc2tuVs07nwxiomlFXEITwsju6NFSn1kn8sSLuL5vjnWHap6ZQU
alAPAO02+ZIAwPPw+b0qd/O5gxdXJFhwjTq17sXfq4DHfgvH13OO6HsFvKn3Sou8
knIDDpfakZFC6Snor+Si6g3xwHWyECpVxEv5WacYbvw22Dlaqja0vgl7L+AO5yjd
VB6fnfc3zfpKzh/t1mCWhB4cG2iOrEeAL6RR7vL0J+oaekDUYb9EBrCp4G7lGExZ
ZQ3nn5ua5mWHrcq5G7UykEdSTNQjCsrQoQYb0/SJZ5+UislmKPXKYl19M+AbJqht
Z4X/XB7l0/F2BOou2/v+u/pKMPfVtGu8cWkktTJtgk9swE3q3ogGyIRyW7fJafGt
cYgq2aX7Y5bZDqOTG2zZSYuIXJvnDmqFrlrcK3nTuaSz1DEZvh6M0OIxMswmFHnS
rPn7r0JGEWDcdlGX1o4P/p6yy3yV+mNKqYv+ZTgJcu0qg7P+KGlpczMOO4ZJGvub
YZzZHuNwy5zE+keafsBd43pc59UM0NOgcz8uRtZNWU2dQGNu6KHRa/9pSNMRPsgZ
rMRcUsmnrhZhRZnQCXc5j+imc7Sg/W7Uzhxm2yrk6nKTSZ8fANXwooLHGA8F7ctw
EYxCn/wKhM8V8RbLq6zTkNjvKSV4LgoL75p6YYbvGi2snkdtQdaqzzcg4aPu0QFE
4df+KrstVPsJU0AVZ/OFsHgFTXTUlOKbJHrTf95t+0atUR/kfyYMZ1W4JxqNaOA0
EWopb+9+uZ5dr78deIMAiOZisVrdw1QMf+4b6BjLNMOtAUthYdG0cmRBgGv1EVAp
97l7ZWkSU1eROIRO7zolUtjbO2ohg9onlbmy2tP/ojwO/Ow9s9KS7tfCaGQsISe1
qXQOxMoKYX/5Rpzx+/xs+Y1QMmzNZTDEX10JvL4zmdCaVWFiwg51Z5nowhei5QYa
b1GajskncoH5cwGqAjnrCpHzA8eAKPDJ+h7p9ikwIw9miEpLORgwW1FT/ZtrJyAd
LXOcG/M+ZaeZCul1xEo/SrY143L9cCVtos/q4Q5NqyLsCxKiqiKBTdKkOb1MSM/v
HObo3HTLYdCQcErCCwpN/gQaFlL8Pe+voXS2F7uG9Rkd5nS/MdHsPMnD8B6AAdE4
4FtaISmDtwOPSifV0/SdkErcwaqc+Q6EfOospxW2h4tRMt/3zQ5cF0O4bYfGoMuP
YxPlRqIWY3Z82ZpQ2liFOGbZPuR4oUqTAimSsbPOZbwkRRquoOapPGyYC2hcR19N
cBPrTCD1bhmWTvJkT34GLlNEkFqX5Uaa5ebbQhZA1pZOamgcJVYGgT6W1D6NHqSN
8wBAk84/9CQqdbrMHicO1TYkCQdNXTuYPhSLS4ieOrniY+wTKto8zZohaJ2t8mSE
pIIeYsd5pBZycY3Iy/vJ5P68aN9+io2Uc2CzcrvMwC6Qyp1PK2HkY7UdASiqtTfo
ktKDcvAZlEJvjfA8mSEkZSZ+ltxCICsKw5yygglzx0JGXtVh/PDDs6eCm71HwRDK
EZnEs1OqeWPG5q75q4OLvUEcLJfoKPc/uOGVGUYE6Wyn8xVEcOYdoVrlz6AjC5u9
hbt08Y4hAtEoHZIu6S43BqcQrT0aYXMaDrmw8Y6ORsj3BdhW/D5UUSM31IRGgLsl
1e2zNPx1S9tgun2mLPQLee9QkQ64mCs0JAnaoG2PD1v9mEofEuVSCGrfIof/Uytp
OSZLM2w3EVN/f8o8vyqJcffXCMjUvmk7fw2VBsxm2IDilquGyBjHddVdEJ6S5817
oWbaGfYDuzCZzEHC09KKol9hgc22PMA3PBmWbNuYrnPmGhwAlXzcSSMP8EzgV+Cg
+Z/7yH3cL4xNhojjaI1poTbVdfUSTc9oWAY7tspAFzEpZSr4S8ywzl+DIGkNq8Xl
VnYYfWwKLuxNnF4OPfcpfQoSZMgk9DKAWMbcnnk+8TW7+3dVX2DwqF2+ibxWNTix
K1BynXVmJuU6Ex4R9KzlCnKXdRIN8i34IFrtMYIGFwraPW6tARsgvwnQbIVooIIe
cgDtQBE3KiXZnmuWp3Wlu2e1Cxf7Rt3PDqvxXJ//JJ2iPO9U3dsFmnAiHKkTH+Z/
0+I+lLbebbNXjIg9yXSUTebyIsEHy9BIKL57j2UazhNza6Wkiu6E2ti3OBfEoAou
U8irnqEgcftgEH4Qs9YU/prMfFe1ryQwaizRxYoDW2cKaeIHT6hDyrYNaZSxzgXG
oScl7Y3Owoj/aL7tSsmbvxFpkT5fVqDJqK2XsELHdnBh6s/sfwbLTUUtSg8nFCg4
idhwEqi8Ex3jTqQXt0Vo9w9XwCq3jf2HpgliT6qG7R1iy3kqibH/9bWpfs9MkiIA
27HTAXZvp7NOT/EjlpsDH+36tmFO57jtDB16lidWAUWXbgWQwv+EBphCQhYw/5SX
aprxh6IUDY86XSicB0LVk1vK5n9JirypftTjOl+SaZJte1R4C3U/SioHD9xhQXhV
vcoHXgGmpwndQu+vTWoZN17n8FoU5GCTZlSAb3JkBGcIpEFPL6fHqZtj4w5Ym8gi
iNbMaczKi7A2MZwurM6ozAvlyPjdykZBm7EPB9+kEfR4acYlFG2T3XFbxkO1Odlb
nK8CFxSpRm3dgvlNyx50Ui2NwAqIT00T652h2DnKMBgirxwvH4D5OeFnGq1RgNO0
EgeZQ8tMtMILT2lZWNh+d8rHl/+17Sm3rCOCj1IUe0grVdkreUImmQh9nITSJ5C5
CXgtVkT+p6lf5EH8D5nw3YNy1PLNKZfxM7jm8wIIwe2Pn+BOQhnq89eQqWKzy7ET
wm6szkgDQN50YPVbfMf6hV2MZvTEGmEHHSks/XvE4TMfLQU0GE0DLBU599IHk6Tz
Wios7LZHjCueZd4jJ+m2VKZCVmfoZN7Xz+wRotQya4TvmBCZBJY6GFnxytnYD4E/
lCKNxG6FkKkBTTCbTNW82DQa52epFCFfbt3BAGOhBz+xxNjW0Gf4+khhHvizBHzh
CtJb8bEp3Nz88yCRCmFSjd1r4TFZ/j3CNI+ca5AHmsCwI4/kg7XC8YQUmbDX9m+p
lx32z8jDEeSLHkkDEdwfUSAYlxVBWt+/dK7Rg9PsFjPMTsgjSMt3AcQvNQ3dsXAg
AlhYcu313oG2LH6/Py3X1WkIigLJJ8GYyi7Il1T1H9zoqSq6aAWj8xJrJZ2ugs8r
KUpAOwWvuYAB1lp3iVqhLVN0nQBKP47YzSqzvxvk9YddP460qtahwMLKzkTdSP3D
CaasxQYCQzxZLoa40BPjbbq3Cv3CONijIauAWsql08rhwkCoJvtxFZ6A9SVMkNiK
jtAH60GkA+THVheP1bbxhxSrlOMbbGyXT4vU5A6q6J9MVP92n/IMi9pjnxUEPtr7
JrBURKZYkenxEgOaNKuVk1kpiIXuZDMBbeSSfy2DCXBZZOPGkj/nwKgBSlk2/kMA
Kchv1DTu/l/rik0HeOFMDwHE8qb0YKSVJo6bzGAA0JlKejM6lUn2QR4gaXwuuyoQ
cQjv7kcNg7Q8GpcSisrbfdxzXEriYTX6eWBUBCD8r++LIBTYJsUP9hjqVN9jWKGg
8INV3zEu1oxlMLm5AG4IBJZ5XV1/lVOh5CNyMdPQ7joWjQlNKYhoTyGYMSt7SA1J
8UJ4u1fSH3OdGtcisNUySJZhZCKVxqmELFlvbKh1sKRyoxi+TP29lcrxajZVaju3
hl33jHaBmdiq2ftwWTmfQ0YKCan4s143pIRX/TPIpLece7sUFHtQI6AF03J2CFY3
mcaGqPCGbfNbHH/mZjZ8f6CgBPDzkE2f01yHeyM/J9ErjKud90NQ8pErJhRXHin+
iAl0e+XWarnAvKR/FlqhsIowV5efn2mHkSq/WTXi6+0b/pyWLy8hZHc/jBGShpEz
P83NH2IVGKXP5xIFl7YJ3aIxcUh18FmvQlk0UMDqxSfP1O8ZyKQ50hkKaF6SDha0
TIHbrf5zZY08h0VZ+dbZ44i+zaTNiJK6+AG3NDpopKQShTXN7tDQISxCezIXSo6n
y6zF8HMBFFkfR3lQxLuNtVX4lgNgGFgBgK63mEh3H6Ln30QCHCIds51Qtvr0J6Pu
dyTW0Ys+QCN8ipwqMRstYkW3QqR59lH62qBVRH7qW9iDxFlQhmvm8zAzW7azZ7i1
Odg7OhYBrHcrdoF90c5RvscF6Dk6ywgg98xmOzePEEGdRg6WSkbG6seOBNWLI4sF
+SPN+1wzARJBJMdjTLXMd0wNweXKIxa5Inybw7ArhPUu8IO2m2oqT92XEce/klF5
Xwr+bDPZGWYnUagatC08Yu9JDPZn+rtQMQA5nnAfaAgxIgJVv+Z/H68J/2CMa9Gi
lMESKt+6rW/Y3mC0WYw+3AdWw6yzeufmKaQCaIZUm5ECD2wvRieumh34NT+yKzRt
n9q6fChQKMm+z9ilpm/jhsJ0YZCNxzUctigp7LfPuaCYSXkUZ00oZK9PoqQ6p1J4
PoB/YmFsRdXGBO6FAGSopqnGHJVNFuI6/YBYIzZ27zbPzhpNiZea7364tHK83Biv
Il4KkOTRVWHwTrH/EKWwrwGgwbIgYmpikeOAe9xk1uUEfamKE/v3RU2Fz+hz45b5
L8IO5eEl2YIKVmze8hxbqx2Ivj17ZA5wXrOW2QbgXzbE3APR44WK5GtUSQh8op1w
j6BliHMrp2LSbqvoljZqKTz2ApEe9WD3W84SF+YocKxnHM9NA5D3uA1qYTlzycdt
h1Y1DRYhytqfqiyBV9Oow0YFXUaChKtOssWWiWC7Y3b7iSVvskV0LrmZSvJznm3d
Gq+6VKhmdcN2djSZkRBEsxHuiGFbUxJOG5/PMGfNbW2fjVwS6nlEhYm+B+cvp6uF
xnn32piOW0I47BTyS1d3HO83ad5YqjGCJ3TR1JhXO7qVgmmCbJFDVyPes2hyNWdx
kjqllG3lBH2iZtxFgk1u7aleG8XBNBipkdJ5VQIwRmaz8zOEo7u+460cXca+KoMN
7+OqkG99swamDXTTIsF0zA8WP7obL+DyDF72Pbsc/kO95teIY4cJAS2b94bsdY3E
SB02gmbE8pNpnQaPOzwluR4I3YVHE47cPev1Go+V2LKHOrztmR1zpdxI2+MAPGIj
DgZKvX1rHhoCSTAakeOB2z6BRS1FyMS0rvWELeRVIhEBxko5crbu5St/HM6Z66qR
Xs7r6+5ivosinvybD5vEETjIeYJ6libduuQG0pr3NAlgf/Aw0N2BTFUGszBZnPpA
kdGHJyLrmT/BA77pIeeIP5+eKv0GYtbCdmeNwoVjNq7WLW6xXj7VBQgtnZ0dSSF5
XwQaYLT2zXAEg4B6JeGfJNvSPUQdI78RIvO+WE2avjx2nfpdN0UpJ9xlveYXZm6X
qxqeb9kR7us0aOC4wpKTdV0AN8Zy8ihUzBOPTahidIXouILgbMRdfUjntjR3CGm6
tPzePGlUNu2/ZjP/Fjj1jrYvmuOK6oVJVsHnSJvJyjwLWb6vTZTo5TQum+8VSmGM
bZ5GvXXM/Kov3/Vv5SW5juY+mvEN1PjC6VvOqc6i1wyAT0CKWcRnn9bFXG1U04cj
RtcP/7jTCQwn4Ur4+JIOD+MpKYeE+D91N5WnApb4LiV73ISe5KdIJXPJ/Y5S+GpA
RXuhlqC/KbzAzlZ0+lRrjS0STs56EEbXKM6MP+F/+I4u9WLYr43dBI5oVuRYbr2V
tccesv7UIe8o0NG3Ao6nEEugIePxd/1IHaRK5Mma6U7G58cSy+wd1UeYmLj0C2NX
9SJ5ZwqXNECuGEMyqcGswSrUmoj0JwrV8Ngh9nYnoBAbdVD+We1HNM+uhoDoEiLo
p2lBPdkeV4rZt1U4RZuLdYsS34sqEnVkMVyBj0HvLJha7kXJLIVhQFvhxsLH/IfF
sFNVwI2O0yG/SGMjj6jWeF1i1BbnjW/4QSamq7MlW5wfL6xW6rmuUVaa28FO58mp
jjUWnNE//bsdZdvvBSXpqIqAajJASSaUNoj9Skry/wMZts6Y3+FmaHFwR4oNaaYg
lWDEXXe8COgc3/L2xQ9nRkmmN1uNFwjNoDQ1Vzh04b6Ff9l58PqhRvbciFMjBrIT
8IPwwL7jbhy+UbfsRFGMZ+DKKhg/KbUQD/216jl2995A6mG+QwtRIpQTIP5O3Cmc
oHRq4ou2RSMAstccRPLj67MQldBZq5UmKNiLqzzCkVpYj6u/Fqo1TMaWYjQc3JfG
05s9Q6U+YhfMk3zxWUc4Qi+zIKixxiJTGf1U/uAJvKL4z7vkb/Esp4iL30TpAOal
iJD1X9YjO1uDTAKGF7vBnbX7/vBS0HM7k3wWeu98b07l07ZxWE8TXQ+Q2I23JLMY
/BkMK4Otz5NGQnBJkB4k+Elg9+//3QTN+S34pt+celYv2Y4kpOLGoLHiKw6mzA8o
DiYEWT9Qm7UjNnJ5MpFx7GA06PtNTM59qWP/wRK0WdpC9Djc4G19iSuzt8bY1U17
DcmH7e7SQ3KIxhuIDJTdlntsndNiQltysbuUwfPZ3jp4AJNAwTRfkMGqox4ii+lA
2TQgTALNfAtPyhf7ATDrgRuQPhlXv3mOdlbduMjrvhLhy00UMhe+8oFNwjF4n/Ft
qabP4jl7SBuov4cC/otnA7cddgZlds4Usn9S8y9hJ0Fj2KNvoHSFFjudQu+m5chX
+c8MK79FIQzVcX6+WlPFkwkghbiZl0DrBoIdkp0/wSArxL0DdKfZmy50KjZ5H05g
IpmC1hQc7xyti1Je/k3zECunkOcW28ZhZMG3hxzI/InGlo2JKW/s+6WNm4+8Ze+I
M4kKC5jxKZf0NREAMPPI+vBbTLGJCuUlh/nIS5ngvd5OCLz8AivK5HTuqBtxe55X
KVDxzddQ7ZlFNat70+pTcD98XlV7P6tvN0miGQJ2ZyE/RDIeAs9SZsLEheFWLj+i
SMzdCJttSXUrjUXdBuTJpaGvAoc23e0eEHsg8uO3SguqRQreVukv2TOFvjJN+PJn
UntfBVosrQ9EdPrwIYGJA34fSp+0AulNvqe3+Jwj6MUbqYj+EEIWpSMswG3bSdxk
jnPjRAs1Q7CSsxER7TBbCY55fVCpaO4OLP+bVu4K7uCd9nZS+PFsxiXG9cnlyLpw
+Fj1807gfrTblAktHbuz10J38779iHzalzu+kljUJh4v5J/Box77BbLwMHObFPjI
Uc/0fmYfKcqMqAidcYyrlFBlMOLuhjYXspUfWrFjKnlaE8ZowoV+A10XMMSg4xvX
//oq8YaQRaip04Yjiyq2gpRzCktF6O7aI5Su5D6xmvFlM73EIBrSH5GM9wwBfOzt
ll4dqrhpBEu4IKWDo/gBjX7ANmt6R+kvae74jczwI/OAmV3gij0oiM/vHea9MhsX
8zZgkBo8flU+gynKZxvSkkWz1xkE1Jhgl/8CKS4V6XCCAl/8NkzqM59alA8+JT1z
jYujvRBMieeCUq5Dhb0sksQDT8+cE1ZR0rgZrnBzqd20knb8RVG0uP5VoFDbsWEs
fWPtYKkCu9A7jm7WxNzYG947F/NrysQlujpWE87QK24iD2I50yDriHbI1ZLU0EZH
lW9hs5/juKdLNxEPITqk9mcJFWmpFgx0VX5aR9RBWkiKXxDfoAcxz5qD4QzoO+wi
FCUVf7/ohuV7kE4aUvHLrmDiSMfq7fwiHoOAWDBHPMDHVse+dZBlnvA7l2JWwA+h
dztnQQaVAj5S9hZAuWKPERinY10CsebyvwVVYld0hpJhwbE+76rtN6+Ha73lNccH
w9Mtky7ov93Aow7acHAawociiZO1nxwFkp35lFquPXMLrcv4egd0qrIS4Kn3cTJH
B3BRuaj49yNnAXxSFoPZq4X6hU+YnaYd23fqSIUeXK1EkKEDXBMf4oTT0qLeulIs
P+nmNhkhged+SxYvOJoXu5oX1/visIaQD1O1jKVBCk9giBFI2TWKggmLwStgL70l
aSrLnDiu0r2QZ4nL3sWRQIkRqdCMRyc+9Qlf3bdwpqmmnEaOx5HM2CbLZ6pwsu9p
Fkcbr7V+7QYTxC17xTxHDJo5pkRbbDqLPhEMlx8hf3VKSZyHv8cxoqof9KrCmQ6c
YEH/UatfgBufkKbiUple+8+bXgsbe7HVXxfihD/JXAvdv/3/d9WtLpEqjYpVj7iZ
gJjg0wsseZgOmWPVEW35kYQJjf0ckX1g8u2CUnUthV5Hi72UmrUs/Dypv07qfanU
a9ApK4y+DxOoOaSDkK3LBYqTKjtZQsAYFUfbsfW7ALkrU0+2fV/yc/BiMMu2NA3c
5sf4dbI7IqgpJ4ACJetyI4xXWbEBSuuvBagb2VzcrAAMH0RBGs3KpL9c8lw6OXsM
5+Eqsnr60t0FtAhOnfYJHW1yMC/evtswc0EcxVHiz8F+dAYSSBbxJI/UztNsTxE+
pHgnjygJLQ694uVFzPhjMzTdkN30DPNVJk+5B0oDSQfEenxCdyRAlTuvbzPdBYW1
1u8xJXXhQywjoJdVtPOJ6hCmKOILAP7sqGuNKNTowp12LlEkB0szbC3og4SLzGZD
8Afg2iqKmgjE8RP0ZW5ZGqCeYDA8JArDBu/NahiL0jm/SsMDNlXH1eO3nTmRTema
paORSuJFotRGHFnqVIbuvFxWQT8tCDavIN6NyxanPsBOlij2kNNB57CJOnSv0S9n
MGRFHZDB4eF+2BKIgI8CwUtRkjoB6GsF+MKCCoA45Xfm6jfnQyiaUWSK3irdpGhu
TbAY1bBzTzOhKcOb5MgdQR7nVWeZoD2rzCHfLrABGscliuLFlMRsonJDylyhF0tA
sSCG7nqWBfoQIQa+wIT+Dz+nQI5Reivc1zFR4cKBrUDRLfkr1UaShTsj8eZ5WhLL
niEhiTdyaPNssITK0ASffSxeeD5BqS1Thj8hZNvlxLuaSt9BoKCZrnuxrpnCc5bN
PRcJkGOX0YOhy5E8zIea5VOoaWEacPF84fev4fLZ2Lg5YSaxMjkKjnc+9fNCwb9h
4aonV5sXHMuLtydsDbhGCO2/XVNOD+lsrFuW4yMjfGSvXkuSo/dLwZ0fllsYL9UT
7MRA9vyqnJ9Aluy/zyCKzVllZmhHvCgtB8LbVytYtHrZn5hch2x8OqMEJ5MbX2Hy
+Zp8k7dWW9RME4tHqcNNBjGpvM7CUW/RrMykrQ4YLnzrua6KozNxuCeqJi0rOFCy
DXGCENb01bpGXcgRIRIfIeEOkSOQ6yccC8e3Hwp7FcwQVgPRVuOivbF4tfFZJRZ/
dnE50H2ykzES0rrVO7sO59qG1a+BVtyTu9VRxUs+Be4IxxkEOlDiQoLG3wZZCXda
qTNiiz8LPtoWS/1bnafXeyrBsVvTuyTgfbt/M8yE8k385lekNdr2UQFKoDNLGcX0
DTCcO1jWFlp62Nr4loD9Wr+gLjjTIP9hCFeouq6+jDHLf15Tlom+8OED/rlHWfOz
Q8x8CE6OZ+G5vecXBYR+5oMPSYJn90iPMXK4ilkcCLZ//gscgRt13e5zA+8/zhYk
8FxAdE1F5c3d9H6xUUstSwfc41Ig5X1OhXuVs4vo7M0m/Y3Vuo+r9abqMwtHqNVj
dBBnGd3QMlECCVxV+pDZVwkX32aJx6yapV7CSfVWni3LrBhLn91MN6ObdMsGkl6A
ZwtE1HVSIzvCSOLUdj2xp/WA/CVY8Q8K1pyeTRKUwfHAYIBcheJmtvPBQsmQ1CV/
oIzMcOg1bcRaz6+lzGHAWOrRUa4iAAos/JP4QxMs5Gan1snBgdTTMkynnkBDeyq3
BfPelfDKLow7ACv3qXhGDY0x0A4g9FqPALN18Tw67Re0Y1go8RzhRgscHP3twj5Q
xRihrfBEfuyBFtRQwBDzdH+zYQAAMV12vtk6WRH3dSomjfSXn74ynA3TLcLtETuu
AvsxVHiQsIIezrGZb3+zZ1Z8gGf4NwGhNvYXjoygv7t+CAqyWBsTU5U81nL+6ee9
SnndJygBvSF1xCOa2y/bmYC/hlw+nfFgSETQ+QuwOr8wtkAwo8kJjtWz8Peid264
pNr4S9Ku9e4MJlucD3Taqs7clrgt1Zd7bDKbINFLdSZEiV27dTjXfdo9X3Jj7iwo
5yXwtsO4SsDTQo2FXnCzoEwQfuDidjdU3ame8+t8k+6jKa6gzdJ1Nmo2dwn+yx1R
8JQSlmQh0k9ACpK6zEcl0xhlUWTJk683AVuMFMWQOEp2LVASJ99/bUkmTmxrfn0m
ld5exBysgJuS7KLrSaf/84SyTWfq/43gw+HcWTX2w0+elNsE/MVXmLwGTBQOb8Al
LkS5bSNaQfi7aq8BmJNoD8qw/XmI4ERCQfd6N58m3KDMFftHic0/d16bBZrm0cS9
7x5W8C4owqCWGNyx6OGkC81l8Yxqe+56EtGt4owTHMPWV+yXZspW7qGwAYMKsPcE
KXG85bqSc81Tscfcm1P1jtgX+9f5aKT66D5oDGsJXVepmJHklb3iR5x6OlK5TasH
OiuOoaaZ25XGMf5afeb6ehSZyk+vBiRqoJakVH4SMZh6Si8FudqH2FeLBOT7YFlA
lZEOzW76WIlGRZmHhJjm4OsUKj4auTpTA6tYT9z5zMFXaQav7GgZo7JQQOqhoF0p
So7da+gQfSDHtmfoV2VtYlTbVwB3gQtysWLjNgYgSFy1Ay35cyGEuZ9jtwLxtH4H
qsHJetnKs2j/Xm9wZQbBYUDhDVclzUU91NDo1xqWoccjWWnRW1vP96s60HRZg+OC
yHe803gmLdwRelODZqLEMsl4cEnilDsX/wiaZCLjn9cwGqs8S4fecqAeXg0K+g/x
DFh4btc5L5PNhfHMeufgA2yU7xfH9YI8cwbF1EGQWTAGVh2/6LaaYIBapFbszdQi
Bx1QJvPXXae0b2ThXcy9pqk6po684m5yypLIlaFBl+cQP6jr2xWu2Sn+vlyR+rvg
Qn/HitrsMVdU9V+IOTq/vYcFqAPk3hOl4k1c6KhuCNZhAO4XA9UEj/H+pL87ECuO
YUTcU5YhIyiH1UjHZfB6LSNTJfkKsZ3VAuczMmV6JSmgNuIoJBbDNW2OEi0QUQRj
FeHvqzacrAXUO4Qs8Aee3GOoqBmceiivOmD1f1q8fkFtBVVfOC2TN6t+ozfL+Gal
WXvYAuxA/tj4NlyURpVw6pMpPlBDJcUSMU32cQhkW9hSWcqwcpXglafqbkGtV9f1
8PzSjBCsJoqgF7qKdyN3ODx9r7XPRSqS3LCVrsNA6gSKbT5lBwDdKEpwCAHW3z18
jVzfeoNf0KsU3AApahE5xBscVlhSEEj9qtbZBV1b1j4lnUdzubsw9m6pz+4xP9rT
W95eSRDAismgFsec70X2bRfzehz9FJDh7+1VqWiaNuEFQ6M6RvkuBAgGuEfUb+QR
47oaf/sTU8unfT7ob3W3p4/iOP3vrTtY8MhLt6GNJMdqR9del6QgCh7vpaA4Ahl0
oft5SnNRYe2IJ/F56n3JGH2c57zw5IzOhT+GSekdFFavIXBEhTWKhHeL3Whe4oqg
4Nhc+rrIx1NoB1hl/AZ9Ss1tv/ObH77yhkyUIi8bD2T+tGyWnM+740fqngaFctYy
qKhVEuQNkS/fik8zqJ07D19cy8S/W1JyteVdA/FCGQCFTLFpEziOq4VbqPM3+0Xg
A4hP4++NBHhfvQaDpLhtR8hIWlsZKBobwQgrUFPNu3U+zvMOBDoDEM38bMnSQcyN
bZuBvaLGMOccrbXFwkDMgQFPEsMY4gPs1LzUyKRuTsIU9GOptfZYHsXONkLAkelb
cYENwEuJ/kT8qWNHRlhFoizTNrDgjJDNeQM19T2O+l300t6miowC3j7PZM4/FMZ7
/t96RZHmXtERn/fm/BW0SvlfVpLOfnfPNZoXvQLrJAtDeHK6PlPIp6j8wQm6FEzI
nOlAJkGrMDKU/JO13q/0mAoxsX+zJoWiudPXciEKc30SPG3CvOvt5QCIiXojK06t
W/PCw5/s99Oxu56ZPMfFWySrgId2u46d0B4UQFNC78PjCwYz04i7ADPAPSYF0PhF
3PFqYjHEYhOe0dK1n0kD855LXP+zQGPq0xWmbdl/KAOi8k1oA/MGuysP+MRC9WHV
1lSoEWt4iQw3ljDohRDzb1JM2GdfZ4c3aejloYVZJRb5y2fntBVUF+59mntPlaCP
1N24bp1yVpIjNMw/G6SHHQAAQ7/mt1nQkt2ZJLLs4TL3xOa5InTZ8aBsWaSPcwxZ
eM+bAC9ZaJi2kPhDIozrcg7Mqyg+Ouk1eascjtn2I5Ms7EcJ+A2ub9fh9PYjazVX
RmW8bybAkhEZqADLClGAl15Q4a18g+X+RQzbI3GLSkXlIUqhObhn1sxLPRp13fTQ
F/GRbVLImkbzKHeVOrj2bHk+RR6i/toHk+6LhTSl2Qcx2GW9sONdtQY8spOPkaMK
JLjn4BjjWs7+VMXJp2w0J61YpABTQMFMEtONokJPBEHNY+vn5povKPQrFFdH6kR1
3wqcj3HD/TPNn+01rPN2/zOW/dHHbOa0pSIDm7nIps+GiP91fQyo7/GE1zsWeepm
DVnWXewegFo1Oq7nCXpaq56gte02lybyv0G+drUR3CVYtSKlAg0U/qgHYJHreScI
VeCnp4iiRn4GvFYu05BsvKNr3+RJgcMFGstrY9R5nkSNeGQqPbCSZr4+NM2MVH1k
5h9xEM95GPrJpUmtXBucYvF9viZT7dtrz74SbGcciZmK0cBQ01n8eXD7sE3OdBAt
vnuI11gPkr18x1OWRUQNNpDloNxOxyX3RmVdk9nwNAR5paSIQgAtz5KZzGt5ETtw
klOy0sw3zX4zqUdjOJp0yh07HhSoE0Y2Aq1uktPKzpBGm3kl9OhRtpvqJHH+8zlA
1j7CI9IH87uH9tSHMToZurIQ6dm++/Fc3v13H8S/QXQ3guJBYX9M4BVc+WRoyvoc
D09+xobqcjzg5FZrlx72EUo3mipOWWwwRbnEgRqdSJUfFHd/xwsqsnp5tx0R1NqV
w5IqlwAmVBoNlONMc6p5i3gu8k0WPxRl+b4g+BXBySAr0sYPWJX2x4s/t5ci2WMT
4hCNIRGHyX8EQfYJjJ9KTVqi4GhFQ2K7yofqdgzci4e3q+AI02IcjtnQJ3y06pFf
zmw2v7SrX//rUfsY2mVdU4qj3gcn4GNQXPbelRhvod6jrMiKubnJeV9BmyQm56ZZ
80FJaLo/ETFTTPLRS5S9xSqlQbQcbJMWUacvvpJ4d7WBu/sz4jyMAXZ4V/hlfVEE
TuSBZM0kigsfO7GySNrSrEnBcRS2hVc7Tp9CKYmiR2fWMEtTdw8C2l9qZep4JZaw
3sNlpkckcyz1/kCPn9OtUXFejtm96RfXnbdEAtvwzjhRe/X8DJGrc1ENpQ1WACbE
VCLxdp1NXLP/n19gses7Cdjb9Cw+1wp1SfTI99nT4VkzuT2mxZrOmocSpQ7G1/qV
tE6Ep9Okiw4wPJpA4DTH9wZkk3WuAS0seX+7R2wGearAf29SHurqFiD4y0/OkAon
36N+rpiSWKgfMeOjjFDv6McRGA9YZPT8TYxq1kkGB0+cJaPqUOnBwpE7FY8tF4xA
K/UKVQ9X/50zrrsL7EtzCGx8Grc8xJBajWRx5xs1x7/BsXZ17MalgkT7rqlv2YRP
6szGASTGvANp8sDgDZD+NCK63s1L8pUX/Qyv/QACtHow4vzC+F3cEbCU+FL3INh6
UFVm7VccErC2Sropd4YVBGOvld8BYoGNxktiQx/CcM1zXOivRSLfsqxlR1JyvX3A
Aaz5cnNnSXNDsHBMOSRLyWOnv8b5o9lNczjXsdyaY9TCQVM3+azkf589ixAh9Y2p
rwUPHQPNcvl180XDn3EEJrShQCFpY5t+vjYbi01PehoRP/h/Pbl4GCKJH0URcmCW
iI0UVPRWk7Htjm3vu/qTJY5crJlujRDHM43PIR8xwe4ll213360YkSaCKdDmXiHA
pvWhXXOXF8CIx13ieRQy80V3A7QuytUKb2jbW/kBL5Xqx2MLeQbZmIOHOB6zWUpx
56JxIyvUaBg6rBhcylx8tR6ni52FoJb8/cFgOAWG8m3QU/GUGlklpX/M9ceO2H6d
CXhTAifQmIp/HsW76xKHm71o9iHeD5VI/Ku2oda+OoaPTcwuNbhBW9MWJrxOXnn/
TNCPrm8mRDm5xoRBtd8JCDR6//pMfdUMz8FPk+4GI/tvZDVRt2GY8gU+Ib1xe+LI
OPDZAtneYNPS/ojLqmsvw0XUz8k+X4AYvn1yVLrkf9GneiWmvfda9cO4KLfsbZPm
59eD4kJYBTSFLkOiESFWTTZQ18ZmKmsVjLRYOXksF+k/3v6QvowfaopswSYn98hk
4JVjPrjdJ4RpnEi+9MgcCB7xYcEiisdn707XDxPHVPiTopLHChz8g8LOqXsYbzhu
ZGVxARErUmXe3JQ6jhldHCz5ApnwcgKZ3x0hShh1b8NSS24oySLMK3x7SAUPLZaN
3qkkbBwUeSOi+4Zz83kcMzj7C5MgGEu5fJ86rAmrKihaI1cslVGjiVgz0nzzJ13R
L8HlofU5WAivN1qc6XupnejHxDh01Pv22ikc/zqbofkKUeUyumkmF805VTbGuUX1
Kuk/peP7BShKDx/9D/Tarb/NO//dppfsroqCYHgfzUvjM+DNJeBybwRyjr0PDQG2
PRQhrJuXYbjWfhqWZ6ZlMFZJenOFyMdAIoVsF/2y+5RHXuYLYdsRXaehB1r9aiPW
KMq0T2dq982Ss002t4M+xgSr2hz2H/TepHtRY7p1T5ruRE2MM819l7PVebB8qrH3
scGNiMq/mbdcvPo7+UnPcEmfhoxHRCY44wEmF7IWOF0jU4kHP5KB8huLKnPA5Lz+
r9JeYF2zQh7Hk51O94hs1EgNkyBGo0nsSO98E3OFUFPIJGnCC5ifQLm534ClRhxb
jSpi2OiTX4g1wWoE2zTC3p/f5XbhGHOwdMRlLU9iDZw7GX6MkwuW7EoV9GV7LJ19
vExYRTFNCueDW32TxDI/zsmfWyp7gDTuwf4MJD/Q5MN1MoOLbVaC9ccBSLQeU0U4
VCo4oOc+ru2Vi/OOFr8gX+HlURzvgQBNt31Mfch5gfX9CWrkZBUP4HNqrTs/kOVP
Pet66xgV1CdDuv78IfA14/acCr8A+JG4UzjeTSMLrbCWzvFe2SBPsEm6dieaHIml
fBvHUyb6lekY9SAyZL9k4UKzBS2SUWe7Jk3vbS6QWtNZfGZ5OqZeGlLnss4a4UVM
brxZdwC7TT8I6HhfUe3L2Dig/7wJUqZ9oJRsVW2iOtpxZ6lcPCExJMdO4bgxeG3L
YsY7MxlDzAk3RzAFfzD+7ybLJhoxAnKSRWHPZzAMsyeAjY7Bewm3ppt+PKqOQzzP
n4Hc8U60JD2NQ4IycZblMZXHYWOJCiSyDiRq00xMVUm8sT9+dXZd1jpZxPy8uU6N
0R8352St79wljeseZFFZ+9CP/OItyUl0JtZ2MPIXU7J+MU5FrIezVkOD+TcowasN
vmPHnT9tfkz8Ck/1ghDLhYWpTu27FeAiJI1al5o79DIUAQpz8tY1lfFA+DA4H7xu
f4padH9NNOolqxGvgft4+JiFwhpLjbvkY/IAJE+0nCSV0gprXxZ7v+Q/9VkSo87y
67foPU9sYaYELF47MKfl61fIRNa/yZq4son7Rs8jtV6r0b1lHYozVCvGQuOd5JYv
Gj1M1owmnPjMtHFedskI42FiJpJQef1IiPf/+ojCesY/bsHScXNNEPo86KqISJIv
1eIoapCQAEqndJGhFRGZBEgOg8L2rzlj1IUTJbjGQtn9W0VqkqEFk9gIK88Bj0fx
FD2tZIZWHbNvgmCcrmjg0PHTY+/k2DLqMpMgFCJW6keZBkCTv0V3zAiIYQzbds0N
cXjY99Ya9iTk+AnI9PEzzl0FLMjba5+2xnM6lgN/NzTLpHgy7sP/HHYuOW8dnSzo
4FMkmxn+RNAJGlbU+e8oKmm3cT9nKId0jCmpBD3YteS6FaK8RppaUSju/CYGyvvc
4C3OagjG84dSniT+mPho6UZjq3QIMRWphAHny2Pz1B1WFfk984NRH2IuF/AzYW0s
+8ZSaqx6BsF8oNXSWR997hFJV4T5wvD+KZB7PLuJNuFL2t7SO+WyOz/YkcHBF02P
kW+nOWd12Xep/+coT52FhI0d7A4g3fhkMeaecNtgWB6a/V4L/3oVeuxNLLJ67q1L
91OfGEl/ivOoZy6+KuDjDRlZy4PF+tx4BZoZ/B6zOe5tHeyptHfuD7o5KZUameCM
uskxpu+vihNG+Irvy00yUPLSh8L347UHoIVh8ikKCy4gJJ+EncUhGb0TD5JQgc6D
wwC5iNolvMr9MQCOeXQjfT11Z2+MY4eWm5KEGfLdc5slAUX/MbwOYjpPHuooEdTs
ksqbJ8bvuswxwuZ+McBMw8xiPvfH5qszYLTkJxG2IBMdevkHT85s28zOsn0plbvS
/08+4ZQ5dLtjq3841HOUFZGd39+YD8O/2R6uf1pPZ0hgq2lbRZI2cdlFjoKPUcvY
xkpBPeA+N/l6WHQSDvky3MqxMCp0LICzqz8dqVIVNs52BYhH82hF+jwCaMqPUy7+
okMxRHlqyMUZ1gIzPbmw081ttRe6XEaSmd6e/S/+9KAvBGypqgddPqlNAueNP9JQ
beh3T9cb0RCZfQkX+CJ7LRZNgjoASBMsc/4/KuZMn9TBmYT8ZVjND7JCDVnLdXxZ
qiEphkIWQtFlc67df0B7CClc38gAk10Tf3l4Sm0yE6fdX/0wdXZzGpCYw1fAWHcv
7ZlFCItt+7/jb58Szf87klGoOD7mh46l2Elaw/EAN6eztojRskZQ7g++dDzqsQS5
hy7iaeRu1BRyqq7NwB25TKFq1KPD8pDcxMDYmPm0EWcY6tT09TPduXmwxOkMzreM
a6VTmmEFMGDxxZA+639gIRSadxw+xdAyeWBlDDUj79JGWlqHq44stVzub1LnJJDh
jfWwgGWvLtV3Nk6RySzS7+g0tJpmKvdnQBqGT+epIXdKTkdVed3DYt1UQYknWFZo
tgQgW74Byvt4Fj0VEon0OjnvR7jRD1PxDM8kjAv8lEca3c8uo5s2QCRWdNRuJBfT
HWzsXUt5zGP20bmxR5XgCqixvPv7Zj4pcoPUWhff5xZzRS0N5IAIujsvExtdPN9A
3Q1zoMoQo1YMmYuwhT95At2djSwt+zUnKJsOUOZJ9JOj+cfdA2KCovO26mbHQHn3
5Xn6DfRFv+UXxg2cs2ZXTUuBaJgSGUHb14gvKCZBfpaaE4zKyKjuIB5sRbdi6TdM
HAPMUMIGkt9kKaLlOU1WhDOkdOV1yF05OhTYRWdr9oJXrV/j18an/luGp91txwxj
mM5WI2oAJdkBs0UQHv8ddUwXhvsgf8UPDlqbYParimPT0k8aGmaVZefgxl40b2vw
UoPB6qCd8XWcyQu0TvEObo1446+XsRU+csFFH1+xNKQneYD/rHs4A6J4WyCkI4pA
qQ8Kj46J2b0/J5+d5DJ7Qs31QgXCqDczJhpmTNrtvUZX0kRHGfcH2nY+wwoSXfq2
e4dNAyhIuVccg2DgR2HrQlW0U7cRNQv70jZ+uQyL9TSTFKdpDjvIrlNsvDD75sD7
H0D9FEWmA2hVD8o7C1lJk+nEBXF6K3tj9sp3I+L0CcccDpyf9fyNaFdJw+Z8OeVW
c+C1Tau1b1+LphEJBai5poHwXut8JCpuQRlcaX8GsnG+EgbMkmdRvUezJvBVvC0j
q31KTW94rDqi1fBqgiBR+lseaoXIYGY6BgtcDgxebmtVBX/lJkIK24iSPOchjNX4
8tRL0PQVYBJg1c9y339WPAp/yXeVyxpCjlytKKBauRUDVK68MbIdeFSB9yAWzAQY
/vjF04J85F32hRDzH0ErQG/uQo0FPmC54LfPR+5wMghoFj4/D4DZMpFgxjuW8LWN
pcdfrtO3QgElEwSjhhMPbntlLSZfYpWEa/GPjzgpDGK5gF+ZF18SUInUXYEwPg4a
MWvxdy+6KPeGzrJdVd8mDH00CSQDC/BE7yrhz0yG1UmDm2XmUYqxGgGd199hvzkV
A+JIBzNmudRBK4hFZPrbeP0rlO4aOkgzgYRP+ABLixGOdUG6FpDloai4DgYvFNew
A016DPdrMilMho+3Ht1HvdZxWNyAK3pgnqVMUzN66WN43HuXdD2yLXPrt4l8V9kN
MmbR/pDtC7zAH2R+hvECmOa3JZYGrSBtw000dSZ5wpKPWI4+wACE5kUJieSdAUjz
mG3py88/DjxUqCMFyx85gjlAqDGrN0+ebsMkw+tX/D4zdZcpaWOzdMsHcAAglOub
P/tMXqf11MIsX+poEYwc12VOQm4LgKDolo5qDiJGr2DjEPPnty4AV7yDPuEBmF29
WhkTgDFPbp2qDtF8CFzaLyF/y7oIyJRYCpt+c4sL0j+tT3ujdCRMoFb1nlH+tnxF
35eOcDPhLcGLS5ohEr1BHCUd/2c9m2iy+DP6yXrYm5k/FjnnECdGxi9simtNFxIx
jYVQUEweSvQj6xs/jUB8D40qv5QnJgEKcWpjSzDDGd1dfGWNG0kNM5s9rr8vku4w
PWjYpbYkUCzUlcL87Na0f611ZRlo7eOKjvScp1zkIOKkdDu4olJADczALhdk8ahc
l4FM3OofV7UHfLVLyuzOTEPhiQHocxgdH6qxqErutvGhpvmCJ0pKhQPuumWcDPAn
/6+PUi9xed+WppHVx6dz4Sl9BaOav9d6iQFhakGX6dSd9IKVU01qMZ8Ct7LtE053
NLgsGhct6QXfvq/J8lwd8dQw5rMAhw7A9uj7UdgtLLIrKznjP9an4afaEMis0krb
bEr6yu+A8+vFQ8wyUWj5lPFSKNmjDDTwW5Loc3uYCxpKSfsAhq+MG+PYlMdLNQ/G
oeGwOv7L5moF6oVqv9kxUeNXKUv/JYerKa8ZImqawvJZXh2XcnkvPILg0FIaz/Zd
Ou2XdLu8NOxICDKuamwTuei6tVtdMHlWs/yJ7AhI0eX8inYAdBelqujMtUFAsuHC
EzpoB7piwiMtQb0LbV0t0VWCS8RRxHKqeAZQIGIqEWkJLd9Zjl/uNejofZTza4Ny
YTAmqEZVPa+n6KOhbpYDaqT4dKSWybn7uvzqU8QiItCRLCr8pZGlrZB6RMDM29b+
hAzCiLgqreGwhEUYED3RFko/PLaT0qo6Eo9n+3U6Top8TIBj5P94WGG8aoJ4bWgt
U5jil2VKtdBb3JXtfMBY1iTdpfT2JHn0jBdbgUzjqtcqKSF4X42IMUvCoI90t0J7
MfCfDtcEYHTozJ9tY4PkQFxgNh1LxoZgMPCB2d8p+N4f/Ygd8cZk/zvO2zcEmn9E
Pv5FHrmETlm4aUZerEwdiARzOM5dmIx/cftofzZaPEjoe9Ivq4o82feyLfiKgsX1
+iMMHSAFx0sLE7yf3+nU8seEHoK8H/3W64MAG75sg8lbSNQV9OzWIFvDNBJcl2Mi
QEqbcDergVguZGaZrFdMWL84ThI1+GAGgn8UmmnPsPt4hR4SotAtzGdpw4a2rHke
T032Q1TfIcgD9PFebCqCNmDnJTcWX+XlOv2Rvrf1CrXdCposmYagWVnR5jeJOBMB
bigJg0ijeBhiPVnH+ONngZIz7z32oPP6Uf9QdRppQbDRvCbyZz42yb4D7QA0DmbB
b2kpozpUXKaLiOiqtvOUB3muIPwKSMY6NlmSQn6QL5IugDyxBfePAA2MyCDvO93R
P8tkBVZI7iUV+159SxNAMrtHTE1oCagslbnpz8vSoSlvIfuSRZaHjvd+838vt8sc
+2QG18cMWjB+zbZi7mHeSEahaoMRPwEd9XYZqJORd8W60O0r0thm/zxYmkM0HMYI
rLwz5bBa8sUHCgKZt0ELxpLSOeaS02mpztAaQhESZl3hI3IOyHTTlcrX19Me7O8g
Pc/r5MG4jYDxpNnFqKGONjJZ7s4bInvDAnyVBy0qk0rV3IG0/eoEzMJCtcZDRQfE
Rf+tbBA8YizL4THH+kFmYj906PqzMaqEv4pE0Z3Tv8MLGx1L6trn2YQcL8E/xd58
LQL/2lQE/MP7pemuh5vkF8XYSRDphu8WMST6V3gGX3y8SvdJ9yo/d7fAyW6I2Jsf
8Me4KlN7FL7YbaYHgG2Hliro1Aob0TYwJHyUcBD+Bl3D1PCfpZl9hfUmhTGVpCRa
cPLD3Pq8ONSHINJsNpiU2hFAErqOuH4t7LCQLt9d+qhLV4B+pHC7SYRgU88K+8Ro
ifzxu3S79mSq4poFBPcMz3nZgXMJuRg9SP3Hy3HGl+UxCnyqXnMvVNPdY2k6M5Z9
sCwZsCKOpHPX49fxF+WuJcqNC5WQDV/89Xv36RtuPHYjgyCaiJlTXJCkXWzJY+tc
DKZY09V6S8FTCzgpzX1SZyqdHTmxr8lrmxBbo0f3CsTCLjxCDKvTH4ICySIZ3ED9
YuvGL+eIN8pQlvVsqQT6wO55ozTlnOZ1+gSyGOU8EPI7pqqhZKMSzJSXGel1nI12
j4x28aTB7uiFA5iNOBh5vG+ZBNFALJOuX75sswuRnFxOrqZBhWQFfq/GyQd0sk1z
RfNZ0DHW2OTQ2BFRURlRhThnf6KjkaLA6/XpwJ0cVEdaTdjgS2PYbRoZbRqOAYOS
IYXW36+IYyF5F95ugvtPXHeUunAJlN/B/osmga64u9GRmmW28LWgIN4EbYfj9Sbp
hUZkePXc3CzBO43KW4KHShMUHh0kSBw5HkK+FQlnIFnUCNvsFgpnoX5KAdvRcE1U
sdl2rm/7+e9a8ArR5CtC2gf4vFMqSXC92JNxxCSn8ZJt4MD+QQgAf1cYR8lukg8E
m5m2BFE9fynJVsg+rbtrbAnf6cELu0S4H/2C2XFgOEvxnZHF0rke+S/Emyu7mLCI
7CLL27f0lnTcVfvYJUU/SD4C8kMpskUZEUwYhCB50wfyE0oEq1AgDctOvc0QqsAL
dK0MWAXyNb7IXBza8fF5lO1sWap3JlDP+wavfpR5ulIcpu7swl+UXNrvQmDyZKjk
Lvmr9lzBwqW5QQPfxIckWTt+iNuNB/gChLRcGZPjcn14BHnqh9J2i84X3tSwKaZJ
dqEOvG8Eu2fKfUR94c0miX3MWFPXcRCEetyNjLtE5cSE8cZKYAcp0Un1S/oQEXVl
ROs3w80bMiqTIifD9QvA7OkKw0SmFiaZC+K4ZpuZ9sjYlwoRummHozUzUziFqQvR
k5DFh7IF9cdPN/l3WrY9P6ZKUwsQQyPCm5Yae9Soh/ZtYo/E84Jg9zERvdf2kiv5
e/yxnD9NukkZUwXGXEu/iDPmyLuju0RUl0LPZcKFS9KTyvSFAbwD1dUNCfuMUOJP
84B/YHeIo71R0faK6ZEHztRBOsYcpzYZWA/p/4s5nO6AwcJ7aA3w51dehBHruag3
Dy29FJNQibbd8Ey7VSwBBgbu2jweD91vVLtnAOX4ZnQKvqAKuSsyZfhymFvjZWBD
0GO6TB6x+CBVWSMM3q38ufOZRV8xMqWzHG75ritT5FHOiyqPppkR+nZdJulE9PSC
OOAKWEQ8r3ov2wr6uQNt4ZpWx5DG4dKDMFUsVnBPvdGdiHVa/YYV/2RqE3aFzt3M
kJi7iTdlVUuaEZxI0ArrDbV2SDJNDcjA5Eq1yII7b6LTnZ4loyLuv5Ma7EFisV3M
xAkPrniiQNG7pY/e076nM3Hez0KFD3ISZ++vceOebemorK/u/GHCwAzi1fnxUzaC
SNfEpo9yHs2DrILkVLfkZbxUrI7UDUuVcqqUXJnkuCYVgPdjHmWluf1v7UA1IDqM
BMnQCSmkR9X8VoDMX68PHNbaA7SxmDJ0uoGcjXU1AB6Cy+LmHMfcD7rbYFAfuJ7Z
wx9B8heTyrwK/KB7hzptb/yo8T2kIaI7HYv/sEq7VLzMTdoADQJbFbfGQnoEvZWD
+wkX0lO3hHdqug0YwjxG46R3NkD8msImyEuxG74ziaNnD0VJIcGr92Ix6wvxcV2W
KBtlLnDbXZB0u5eDchikjhqhcE4O1vvE8qfbD65wCFBD9V/bgnRWL7l0feFciJKs
7jUQZWSKXUwCHjL3JoQVJ4li3uyDB8texh02ErOePguWKJuIKPRpfRFIbcwy1NeV
Ud1h8GZRhWE+ZQYNdYqtE6fhOwCWxico7G5cqfhdDoE8f7N1xd26DzmS3Ot3H2VE
yXwpBesBMroPQSoR18cq0MTJkiRrXtK2lIX6ShRm9ZLF2+XLdVqCNnpJyehDmwdC
AjT/QsjbVWHqHRPYzb/f3q0nxuVLsllWKPhgNri/SRM1KNZOmd8OHrBfC6C3ldvb
jM7nhEnxRbGEvOVKokNoZHUzcZ56FyLQS0z4ATucGpGlmYVf+pdovodDGgy4l0Og
nLVIx/BjSy6rzzZj1e2YxO9DSu90DrDn6LrdhtTb6mkCcfVjeiebxjO05bkIJWvS
dhOpgROKtHPWjFXn6Sk79a3jDt0h3Fm5f2OJg5goUYc/M45Zooh0aDo/27ElQBRT
98hfwhpAojAyGNDCEEKKsruau3LpN+rjLrAi4NCxGgnsd6BAoXkBUo+NAIEfHW6n
AxT7ILtPkQoJgQyCbkQVtuVBJgoyvVAYHepFK+GcrkaL5g2R2uRAtjgXadRciHf4
/i45swiu27LmG5W5Q+AqbS8qtNCB4Uazi4x0JcYmHyhrgHytl/NXKQL1KUaFQ4uv
/p0WvHP40Txfnoa0bMeTNWdlrpoSrE3mUqJsihhJoAE0SlEQLeoCUgADr5T2j/OE
MPmcZpRBe+fp3xcpxM8vYWVlik3blcujKZmd+qKo3BDXtU98TE3g1aaOreXL4J49
xwsEuOZBYLuzUdzzBceTa/UHc/n0hDl9HKWGgdF3VTPoceMpZjp4hIagwJQ6GWay
z1yvfqRSNPY87ZgwI8omeOfhin/a5B4hLnOPeO0pQjMqy4tZImr15QSX9XrJAvJq
/oGf2hh40lAcJMUMXDgBizPXp3oHQEUhbu66QyEOIF4047bkfTIBBoqmdrD7azmp
9PKxqFDDto4hX3EskU2Gj/eAGTy5Jb41e6wdOm8nKh5Mm4aC1pC8PMg2lyc4mFWQ
Qy+wssm+EuJmI8F5EjRerVIjwS8/Ui9Iw/2+kXvTrrLqD7af6u2QpXW1jJm2pj4t
kvWipLV5BzU+xoyai2RVDdg1H3V49C1gkLdO5esbCWq6870G5/PTTu01bq5Q2vEG
6d/W41edi4lrhdqYcTs4YwhbFIgf7ydQogohwjEvrnWnbUsFwChWzIAygJmsjZwU
TeKDyYmhVPfMI02ENUorpwdSqT85lMcNHLX7r2S6jxTNzvGcl+ekmik3Fjl5nMAd
Opug8J32otYDfuspINrryBV0acUO1PgLUveRYAbyS2SiF+weU7P8dweNTRyJ6ZzE
Xwb8MEyRh9MguthgujQ57yCb2iG5t5uU6itZbSC0GhXYMl2CB/rOgxHonXpDPYcN
2o5srYptlF1LFrzw1cX8Azj4s+bb1F+eauu/Zv9qQFT/xpFFd6XABurWiQ4YwvvW
Yt0ZZXsuHRWV+TUPqqdzgKLr7TwQsSma1NPphkHGquLTCLUwEC3OlbQTsMUJnQL7
PRjCT6X1Zs5oNVIbk84HehHiffBCz634XtaCRRbUK68yf30ragAuYjViMNZBundo
pTh4WqmLS4/5087fuG4SFFIGreyTWUj+4ig7r4bbnSoq9ujmRP/mc15PkzQNfHW0
zSdkon1kiN8HrdwIWk63EKRAUmGwJuqry6d8DAoZ7nrnbJ1itybkt6DPqNbPpQPF
dQApzyLZpZhOJ8IeOUnSNjITBiB/VYOG7a+Qm0ULMg+1CC/8PO12HsXrwdF98fiv
V+DNNTIJhfUxI/999U2JfGEFschXygR9u8gQayhmnjQ8ouwZeaCKB6GHpDJJpgoO
x0y6eAxIBgZU93jBmU1m0j4UqMxHK9zCDFvJDW+Ee9oimbjXUJUmJaNfkqZ66tPl
hFxuBlO0zSuxRHZX/Xvm45U1KEYAqRxvPN4JevFffoabgxvn6HAfjoGj0fQyQo4U
2TbC+JsYgBo8alpu8tiLqe/hDt32wG0jC/37feJ1qfkO3ClHdV8nM7+EOOKSpNxX
i7Vn+2vVMTm5X5Si+LDSae1mF9GKhb+3j1PRFlMpFPtkb+TCa1LsMUiWlE12qcL6
YQLJ17MfYBpwMlBYnqm9KsiCrM4YVSthLILwhehsaeITvr1FRCYhrYw4aSwFwOua
FR8lrKlg8Q8XrmEEh9NlxnvrdUJUK7UTMQaKMfVk2IuGX46RBZYUWCoK+ARXsPs9
hqC10vkQfu+kw3NvXOsWoCbwvdaSaWBVW0OZqPXYG8soDUnvbZO51E85ekGebnEa
hrTelXywTb0ezHSyvt1CDKQID6VgxVi50I/wrh263Bd05qZoe4Tzfsb5WD/s8Uio
lhr1WKsrx1QZDZNw3aj95SNC5CVTMmXroQu4wVTtBiSLUrtC9smXaSXeWGp+Qi32
jbzyCuoU+bvdhpVOBtm8ibdcq0LL5neB28qQIWP/b/wcZdc7/9zS9yJ6XAIFmGR2
ktk6m/QuHdHI3GYmaLR/Y6Q915Ncbe/bPNS50gVkHmZqD9kXLGgRY1Fgshci56l5
WMZ2NakJZS7iZ9m2LBp9Iw1ViREfMG7nli2N2rXeQ9/RMerLtStLQWZIFK/6lLcb
w1tx68d1qAdAtXwEemR+ZqK45SiB9+sHCWtrUT4Cr6VxaRXiDGenmNE7X6OahqXU
5SOqakTMnfs+fUwbo57iAdFF8siGfuSsVC9bzCKLr76SBdlZ3dPpWC40Cdak1XfG
tZvnmoCot5lzs8ZZ9dy13qX34o0MMvCNdHxboYSOCD+NT6blVWA5rdy1bMB99UKb
CsdTvRAow415VFGSV3hDcb/hTAQFfo1k7JVI6HRZavf8efC/RjdUepNBVUo+PTin
/8uynFFHX/xvhbZywkqKpRUOYke28cwvFp/n5hyDhL84eRSiBhNzi/NrV0I8b7u9
/3m9kOyjYaZCFNj3BGTlMV3b11YM4WFgBQEesTByhdO91mUVtQJjgGKcsaCu3qui
az1BE0DV4za1p2KIC+IWJJrsjslFdXDgzaSMVw8WZ6PKMjnE6ndT6W+zhAyAlfBs
UKW6nrkDPCAQecx/gDTiFwGBAiFYgm69QyzdezBMzTjOaorF8spLNWAXwIhsE7NA
kM/Lm9bKxXqD/p1aiybw+KnA/hityQldGqiKEx2YdExfIi7AkzGoAkRGrICcABqu
srVgwmDVYEWfW0LZ0Od26AnOQLJXGWuSnCObdCSXm3jI4hkDGAVraVUgw6UhDv3B
9n/TMHLx75WPrLWRMWnv7CB+Z3ZLAwl3Ed7LgrB1QLOtQ96S8s+PtMNMkSOBfLv+
7R3PosZCs/F/BHH5m0UQTvbWVefEKxuGcumvo9LwbFi0M27RmEFaV25yti0poFM1
bJUygxxLXgYTmvPJvZDOsOwYENb58pZC9yZIJRVFccdlN4OkbT74z+y1AGh38hLS
h983EB0hsUQabBSjb31i3LKg9mmQHPbC3PjXWCv0ez5Z62ajRrWAjHldEGLn2Iio
sRVoU9Z5vGMQccXoZ2zYLb+ZNSDmtVxf0qi2IBcoR+/Uaac93HDTThAal6AcC1Wj
SrAfYwAYpHtLRXGSpihRgbXUBoP1rNlsOqMO+OkZMHfBiEMFcK1njFIxla2+UWLY
3d56U79B/LHHoOZ1e+tSaeYqrrLWvU4wRtQA0i6t/+XA9DZZT0DRP2wXHdG1XkLh
V4fnPEWgxL4bDTe0pQT3F9np8xhUAE4h5mhgul0LDt8vL45FKGYaQnbSg/G/4O+c
+XIiCqeqD6t2qXHhcDsaPRI6IxOImV5OQDDXm5gUedea56nYHV7T5u2EsPIuJt8h
keU7Jh2KisBTWslPN7P5GveBfoPmP8qEYpLH/ctB2KA=
`pragma protect end_protected
