��/  6����p�̱]K��	�s���yƻe�q�z�ѪwXG���0�{h��l��0��$3�֏�	�"���3$�4Tkp�UX���ٳ�J�d_\�J��-�D_���(�u��m+k�'��{�7[��g�L�Т�� �s-�v5>5���݆�V+"�@���Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9��X�q\�U�o��8��d�s��e���ڟ���]d�R��e��+h/�deonRױ"�g��9P1�VR���c̭-	�~���BN8W�Y9��$?h�G��:�33�Wַ�k� �Qj-�����OL��i�2U U�&Ѳl]��;�Y˛�4.1�_-@Y
�s��˴[Ks#�"��[���tw����S$6��Hx����ɯ�kjXC��6���X�X����ȃDl�x�n���`�^hրj��[�� �\�7WmE�/z���/��p�j���/�º-��r�8�Z\إ�8�p��E����S<C��_ O[t�BxF�y������S,s/�$n5�D��9�Cwf`�r>�s���X��t�x嵱����r!8�u�-f�T��u��xQuT�㥡���J+9��؜��0���HRπԣ�׼�62�6[�S�ͤ��+��k�G1_�ŝ���o�$�K`
�>�Z6�+Lo�5	ďmI��e�ڡ�)�v���E2qt����8P��d�[~
�Bv���,O����Rۍ��Z��et���#䨾4j��5/���O'�$��E�^.�6f}X�1]�rfhX�~J��P��?GTV��^�\bJs[.Mn���Q�M
L&�ʻx&#��==�#f
5*���N�C
R��&&�nL�j� Y|�@���U�'Yq(�c�R��>A�ӅU�LB#ϝ3�͓�oI5�rO��) nG3bZa���I"O�3�#O�̱�6g�L\�M[��MϨ[�b�uЕV����V!��.t�:��R&Q��'M��Lc��!�B�#�]A�R^eݗf�@i������M�{G��+j�?)����a����1���;]Rn�UR`v����FY��lP˽N�S�6�I|;B:�3�,�Q��u7��&���@�g��.�Ή���&���.m��������s��p�c>v?��*����+&��4�m/�f�I�J/�ȊWg�md���C��h���� �;���*;ל.�/'C>%��rX��/��'�ZTn�9��)�z�v��PZd$�����K��N�iK\G�B��hP[{�X���a�6�V�L>F�0�Ӟz�C��,+CO�b2�&�J��+��4���H����Vp��`˕���Z89��Lf�D]�g�0���s��В n&�g���@s���@��a'L���s�㦘-����!}��t����+j�͎0��l��y���6�'�2X��7�l�e�����d�n�4��i.BKX�6ƍ��a�>Y8~�l]be�$���8϶3�Ł�y	=�ɶV�>JTc^b�`�'k�DV�N���B�MH�-�U��]=HX;��Ki��ଢ଼�4M댭E�r�a�}���C�b��T�����n�G��X�{������f7ɜ2R�I]1���ܫj�)#�J<o�^��C��o��$������k�DkM��S'�g=�d�ܣ�V�A'�3����{�ȍ���V}t9 C�3�.���qi�뚋�����-� �<S�B��z3[����2��"b4��$I�����9�f��&�'-W�: �;u�s3^�����o��O�RX� �B����/z�� O�Zϴ!R���̂�$5��Y�o�s��$(	K�2o�'~dr�S�GU���Cȓ�?�H��R`������l�4,��˅?񶔦���舑������O�9�.\�J3�
E��se�zMÝ))�͚�r���]B��iݱ�X��k�����C�eA�w�M�Wh��$�L/�d�:f���z���ֺ��(Z�˗p̟,�$O�v�P�<LlYP���S{x��6��W��z�b<���]���;��4Z�Ԑt��k��ߕs̲3B�U��g�^�Ys�)q-�����g@��aG8 ��OB�N*��%�P��_2i\#�9S���7.�����/f�\D�R�L�f������A��Yp��E�G�?F�~'^Y5��W�N��3��o�S �l	*x�u�{�p�Rl/kV
c�b�ρ	F�-�J���C��V��<�c_���f�R� ���p�r{q�2�Q�E'7ɛl֣�md� x7ҡ3:�R�K��W�����"q��lP��*<~�'���c��V� C3�y{����|W����Ű$�'z�ܪת~�nnv�&�����TV�p{\a����n�v��9|&��@�f�F���Mv5�i�5	�!x��lۋ�N�ġ�5e��sNvx)�3��dU�*̦�b:�{�`�ǡ�u���&#y�%�Q�c�@OC��jM���S"E?�1��"?u;�2N��T�*hD�����7N����kx����1q�ʭ�ϰG��S��H��s
�=4��a6�u��0՛Ǝd�
P�aG�>ŀo��Ǌ�5^���_�.|�������|.�mY�Īñ�Cx���H�������FJ����T�Y_�yӼ�P�k"�����''