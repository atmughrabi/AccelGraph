// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D9j2GVXXWcPU6CNnAgcKOID8dZgkPiqLtqTOyvCgV/muV7gEF0vN29NNaTgj6uqu
Wb+bPLMBchv/AVLK2rmesfpPINfHm33bBD9Bxsa0v1c9btjnpLAXXSOoR9rIcYy8
sgLCSGz9JzEBNDBkCqbzLcX/M1JGqrE7/A+cJu8S/Kc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10720)
dw2nfz4tSqf2JWT5NP8styifqOREqKiZJNIu1PD0VHcge1q6YWVD6MAdkvNqBFOr
tvKQa+GmD4yg5UtPKtJY6Mf0qxaS4E0YizuT3iAaHKTnHysWnssIEWc5XmstsJQx
TkfnFUbjt6L/v5MH6KArSBF+HVDmxhAaxP/dJTvRVzBPUbLcsFgGsOh2Z3MdPH6m
F5qpnfa5FxX70ev0Vv4tInsFZrC4a50PR5gFf4ME3bHoR0+2HPA8S0Z2yDOzd4Ej
67CdHdtN3xwna9/nCpmk8HYkOx1w9kWAd58FK63TwU4kobpmRNFP58UZWg74bakW
rfunUFBdL8A8lQWPc1VnApct8W4bE/I81xXc1EHf0VanKce18ZTOMtwmkLgWT6LE
YYr+jPmv9jbCRarUGJXtXe5MjJol7k/8e1RIg0gLvFM8L91uLPFAIt0WWFnxMu40
8SoWHD0dNdVxhscXiXQ1X3WpJ7NuRwQy5q5NsqlafdRikNGNsKy+d5Q6IJRMYAUS
4eU3/FnZI/X6OhCG8wC8iI2jCqF11BS9nJzBbPeuqQKsyJqH31RESImyI3xyWA8X
2An+uWbnQAUNzvTf7GNovF/kS5xMJ7WaLcQUX76GkoK6s4wqRoz/WIXwgU9U9Jo1
tw+f21sf8skSukRHj2WhfUWtBOSp/UUr8I02TB8uNR2VwefVyfZ/O7p925SjwyF+
MzvPhHNkiCA2x5cQ5KfaiePLTYuEhPQC+koJk2LtnU8g93QfTnP1ftek7WUMfJvZ
CK2m9ERd2x5q24YWsBm8SR6yQbMC3qkDMlCgKUnXQFqxEvGU8PuOgQggZbNgM8td
OyrIDaOsp09JupUxgin4boGhs5rbd6X5JL2Nquc+oQHsWl26uaed6naRRYOEegQ6
9u8XP9sK3OIJtF8k3qeeLU5sJob9z0U24fSEeo0PezBiqss+onlNqMTKF8doULHU
DZxrBjRbsUEtY3yKSRSS5HeTvRCOEyb6aVnnNAfXOSj7d0fq5oFBGuj47qKUCJFz
l8tUKb07iAixEjwbseAaHWYU6B1k/5wPzkm2ykTI+JzUJ//WKcMdv3a3Ot25rz5X
Yfdp7I7T4jpj/wsgEkQ5alc8mWqJjKPDMKrDRARkB6ax1mFFGHgp/q9FeD6/Q1pB
z3mhTnTg5qZbdrpBLYH/PCLSIZTzjXkwbkGo6TP5jdQwqxZsB2Hyw4zMoTIseaj9
tKp7rFefBNdTDnQFfvDo0yIo1TAdETWvLxBWdhZo5E0odtOcWdkpYVH/ZcQfbRkz
nKlghEdNWIYo/HVP18ivCoTDXxoI8zUdBhlT/vpnESP3HTybI8J/c8P6vqiIY9hp
1VmjDIVMJeSAUChmoxAycnUIYV6tAHjwaF33dxFym6z+9UX6nNhLikR+4p4g/L2f
L5NvmJwgioFhh+RJ2S9coORV6Q/UzDC1h957TKqaHXib0grCjkhQQqDw+m096yf9
6bTgljt/D/iz14QpvZMCfmcS6WunEEuCFxEmxkHlGEosCaivQt4EDmAFfRpGyGJi
iMYRVw0H+C2hN2CbGpDBcjKjSvGtQGWQs8MHf3QGpTIoxBPquaFVPyY9UrxDFBiu
cUjxLEeSgeblFdp58MAFzTB0ANUGKvzCm2F4e4lVEZiOYtbBw6lsgHAl0Atv8cpx
IxaVUB/f64l/B0ueiHEvcXYuwWKIPLbq9HQgoigrRRXFkFoJTG+5kYSUZ1aBVBZp
FEdtEQIqgbg0JcnHSRl/y/SR6gsqeOhFCiQtVyRQhd70RFGkTr5Lij4CIFRfqe/v
hKeNhIRjiMeE/R892QUmTZWJcLHFs40aHufFwC4pGmPGO6jtsV1dHbWSV9F1gcwm
2rCLq/5ATNUJD9GrIZuJs0MXQdNy8xSLShuoa5TqLBu5Z1Vtk1/yhreIfM426FEZ
ZDTz1mK+wIiGtJOlzF0dLOI09gLs33i6ocFphaQxE2Kive2v71R6Fo0nQ/5TAwvt
W1XjpLvwCgZot9en2wbkZxnB3Fq4WhkqPCTS6DguT/0yr1cynIeUR+eVDjSntSok
ZzlVfb1r/N9H+yUoC356ChnSROUbqyLIG1Ze+AJ3jQ+fhzpSGSkRHHWPquu5KqqE
y9dr6zOg8MQ5ugj5ctMALoMNj3r9QPvGov/sf3dpx+TL67T6I9Ik+9VPWiq2vCof
sCCY6tfJPJ4UZ30nhLEKaJhMFMvT8cCMv7P7/4K4n1dF4S/5XqrgwMrtaEbQMsIv
s69Y+V9Ii0qMjvUpmcVPHfOqJSGU5g4dtSlg3MTI0ja6oS9UbjLQQtJ4eBJTXhUX
Q7g11qupL7Pt+otYzkvq2XJpD4ZMu/VrXhgHcP7ypGl6PgyhxuM6X6CgeTjFdAeT
kh+z7InerjAYkaX40a13bGzlhQYP1APj7Lk8PKHbvcnJ9vn+eQ0VwiynEQqlakRt
K5qrZO1/mt1rKCgM+j8Cra/AOlx4G5cLdtG3K13vJdVMbDeIXPyoxua9SCByztfw
cvA6kpGPE8GPwOJerMQywkfGANpxzoKzhwC7fTswXyahXDkdIonOMdZcWfPust0r
rWAMgM605y6CjPINvaUT+Q/sly3fSMxsSO/7Ae4YvMxPCZW0xo15MktlAfWxbDUb
CZP2byGETL9k9jsLueYjomH8ssZ28CZiM29Zc0cJ39Fz6CBVJqGk+HTc4F2BGfP/
FfCXVBtU06ZwMiqBkkYmvOkIa0UhcMlimap47ACm4NE9a5EqNSSQNCkHmiWZ+7Bn
vlecULMAC+jzx0uEH+YWIme79LK40fwS3KGJ9aY2x7AnS7YUP0CC3KHW7xoHn3rl
F9kZPpQxqFoASzCPBpdn58cWFfbMpIHyWQ7FO1ZnSLwuTo1lrsXbPfFFArRAs74u
2R5FaDcY3vUQj5cpk6hd5+ofF9CRd4EPPrCB013/7h1XWBPq0RpQFZKd/2EwjQQs
ZH0KSfZzctifyuYAdh3VybSJdDbonGJLQPBcMd56uhHENuds8K5QaYCB8bNIvFuu
ZsmsvfkJF1T+FtDfV1xS2gYq/nXNYhyIce4YKXJ1I0CbatWzRYrA7HzWwjHt3tCZ
ISGJ2eH6vJ6ftoSBYEPjx6luuX0vUglbPRDOE1hpix5ud/ww3YghrxEhYJP2yIuX
rsvwB3jX0HfZ1oOP6632vC5SYrR2qwoXQcdkYohsMok11W1Fo//cQx4FXZ9LzqMW
b+gOiQHkSNGEjtqQ9Q3ERDbXjfEQy7zgDglangYZZjFB+DHScRRgFh+aSzZsheyP
R62X7oMZfGd6TUUresY98dwGPhkjHokEDmmw2BzZgSOKPG8mjbnAS1M3xQFcJI4R
RvGOm3CeYDcpdQ0WgKenjxs8Jik4ZC1eBILih7KbZ84Q2a6CrAQR1rneT6kLzCaW
TJ6lmJt6WGwyILXrQe/L4kAQbba8KL/vurStYj6SjvzmGV8tgkuSkX+tgs0tQd8t
wtm8OQVLhqoUlaSFcPj6+86pVUni8lhe8JcpKgz24PXJJ4zt1WALxFfE+JiCbY88
SEuthFk1uyftinIYeleG87eaRY9WXEktcGDzTp42wBJtZQYx35rXI3TaC0mav06J
IAv4/GB3q4mvXBlwAYhqN9kRyF0GdojQBR8ULLQjZTfvXja7ix9wE3ZYHUhw/tha
cg0XTypeATmof912+KbGFlsifdEuiSDvlC8BvXrr4sdtxUTzlQDDyGOltIfcZoYp
2Tgt2+vIgdfWZ508VXigqnPQ6qbpGmlMMzfM1w1/snL/XIKpUeMnI/n0fMeWej/G
8QGxLbRPeSTUsQeW54KH32xPktlJ7CCn5N3hw631PBYV2kqKiJpp8O6oMfW6gZZl
IlZjrepXbGPNdox00tS2eg7l7t+BD5tAG+Q+i6QzGdd5uE0PEZtnxUxc5KraoneP
A1K7Po8FHWdODJlQ072f8Zz5RhFUjA7Yn5lUaJZuSVVuTnBiniMSlIXjvl/ubQAg
Sjvzt10YfNEeRC4cQ2uWk1rsFa4mF/S4dyl0j3QBQVN0Pnk37qe/B7FWcvRKhnNk
HOTjJztt8PF3vj2Di88iA3rMHZw8RpawyBlb3JXrE7w0XGABM+2ReedNM+6CrlJU
zFHPjtPvRIcUBmiRGIl2aW2Q0WJ6nu9Zwrd8PPRsR2Ay+j4pZ00cEFxhjjoMt3di
6KCZTT3aS+dxT+6JuxlCJI4QP/tCpZbRPDE9eOP90K1OAzD6z/UPbb+QHF2g0EwL
vgYdMv+UbE1Ig/NOxl47wraa1v2mMnI4OR8mmbUgz8UtsCGaJg1ldTe1sWvHQ/cQ
aA05miTbxbnxJT416yafaTALxHu9xlgfPUre4Yi85UwcyUQc4L6vGmo6qWaky81z
3OBaHi/E5XP/TdePAE5Kv0EaaB+HmcdAMW77AS9Y4F6nSyUqt2B+qyeP+qlVo2+e
u6FO+3nznO6EJKksCX/+QPoMpuQ3ESKpN6cqu7lGK+nkLJxfIRfFR7R4XgT3OT5n
cYDtZolXarIcab7w8PXYUB9+bHsCQo7AOFWent6xsDukV08uPk8HzDZbPShm3+m5
KZXmU41aKiEAY7oCP7oPLZEgDqN5aaXekdeCLoNTScft2hmfyi1/mJok+Ht8Q+wH
mi2J6lIzZPf85GZo2fOrdqH57QU5v5iOx+oQ7gEXyszmpB1Ru2gCLGbhvBVQRR8g
u/LKwOIvL/u8VK8/FIyIunIXv81tWne+uQ8FXKvFtJAxAKKpAc8ecVbYeyRID/qb
Xu2AJsxczjbgQdlNrxQgmZDBirlphIRObCIjNBoutGxnUoOstWOjKX5lltDK10dz
OHK7sgsFW1urEWvy3wj4F9xD1lB4zBl0sN96XoESlznWzUEB0kdIQKahopH3XP1Z
5DFfPU4B+sTR+KcWL4yPE++xXwt4mTVKuzf/wiHamVmSy3flVvk4Ad/0iZBpcwh6
tlP9L7yWXNYjFTZzZLfhPwShxV/Vi+J7dEdsCjTsHiZxdHRNoU1yKCkFie6QZuTM
TLaM2Gc8VZDTeLxjrZmFZEzfqEuDhhwSRikook8C9D2nOBQ7FRA6y5t4NXywYf44
qdHUcKNLaJwTk+l5lRg68b7Bcnw+3wq6MyxFQjYOqZvkiV3BgGxdU96siHPHvEq3
leOpATpX1+NIgB0TUVFEZnsiS4VRrfwuw24UM4qNe641/Q5dqO8pJ9Ymnld9JCo/
h4RBPpKkZ3md8ppDz/OfzeI4fbo1eKZ95rqr27HLpB3kvjgcf2xzOIK25ouAMNhz
eugGyVbbQwBFINl71Jc0vRVQG1rOTXWVdaoqk7PC3VLj4dkRtXF95MZM1wMfC5ID
LoUhPfepSGBhM2hEdWnC8aFnMJVnkHVtZLbAHCAp5OnGJU/2P8O3AESjz4Me9eL3
S1RfWs2xSxyOhezdOxWqw01aKIGv0UXm0MIAajeLWp5o+o4qLxlb/1X9ZiTr46Yn
ch3t5FDG7RowK6ndNrP60mOOrGtDWf9bNK1QV2/43TGl1W9tf9+fh8f7Xy++lL8d
iVBEx2YgA3+luQ6OZsTSz95ASXA1N+wh98KU9IedqE8m1oYxG+4Zuzibz8+IxzA1
0KKlI2S3p9Jd+af2yts4Tv5SD19bR0g4KtyvwfTBr/qxrN8u8K5FfKNjhUJolonr
ZOYSc5FI7QMP4wo7Gd+zo3tbeB2jnCap1pQWswXZmwAg/SfHd32mNJyCfquKKkyb
dIbLg5J8JECeCEM0Rf0QjtsD4rQPCspyJNYsTPVlbJfcWEvzGJKLBLOkIkFj3bI0
zvhA57MxsJ0EMcukpOK8CttVXYqE8HEfR8oOmdKKaNI8EWdjzKIBWY8FgU/4P3qD
qF1oPHzSEEplujUfdw1p3SqkIP0g7xAkV3+prHpSqgn82FdaUXRAp/ZtWKakA3GO
OTSJuNDvjfQyxZ8bdRxMLhDLAiYPytTZZeMQXbJAsRsbXKxThqfaoZ5EJ3ANqvNt
jD0sLt/F4Tz+ROZIqoXMb81rR/iXpL05QqfNiPhkXiSlja35+QG+uAkJi7n7YcL2
b2wA127YfiRh9vGMjD+bFD800UZijsPNxkWGCZ02ZKcwATbAkpFYD6RTcgmiIDMJ
xmdtKuzCGmDMHlTwCkQeyOaZNz+puEh5LW68J7ZfMK24lu0W/gKRFVtEzdArZERE
Zdpw9EzB1kWRXfegNWMuCvCtZ3K/3LEbpaLYHrhGG22I5ZV5YumFipxL4f+vgEUL
aVM/EtpyfRtR3t9BRJNK9uAA2QT7v+klqq25WooH9PHWbcIm42+NxgSm3X0oM46H
O0CvUAVbMktbEbaqYyXiwkeet7xLAh3WTXkgVqGKzRW2z6z7/SMglO9MaihvvK/h
Ok30pD82Gx5MAjcSc8EcV+9VzbnHJEGMtvQHNbRP4hhKcuuSVgqHXdP1uAMhrSXj
IAZo0SoSPLmPs2NEszLIJtjLs1ajWRilbWJHrJeMf/wtxySdZNwXpyV34RoAhqBF
NTmrZtWY/Drhz1UDz57QRuuA4PRHFRp6wGwdqF5ooCNTIKk1PZA0UQqXr7HLkL47
y7yS5a+z+yugimElX0uCkPYhNyt4PlsOHWHAeurYqc8pOQ6JTxc0IUPBciLLjbHj
9TbnlnGEZndjM/+BkhoNOYpEFYuqshC0CgOnfGDQxtQ0wjYR+7Yf1TVdnDHfapd1
yKjLTfvMzkfdu99ghOGN2AkWqIjAZhvILKP0NMcRaYWy0LK+62Ie+VsWdMC0Asiu
1jiNkMR3y8qFTBVptr6fR2iJAroqbyjn7wiKMTPS9RbKc1cfQvATGHtv4gZL/yuC
V+FIO7y2w+cur488YKeruc0tGBda2Un+8iiAu9HOaycRFR+Oe60calZGvX+wESCj
uIhV2sFsabunXccA/eHfGtpkY3pxQi3IlkbucblEfcvWkLXYOSRkD+0IRLjAncK4
5pTbc6l3m9Mnz9JKQMqoJQt0v7YYW9u2zaVbfwgxJ9vffFncKhzwZcc+k3PURGPI
NE4j1/6g2BuTHitME3PbO1vrKDuZIhyqrGvzY+WYOSBYYcyZDBxFDZhbVM/elosB
JJuxmK30Gb/LzrITUyzz6kL3UoWhUiPCGN9kc0jqWX9HIIrr0FP1WhCCKxE90eTc
hpLs473dlu4tyLZkjN5Fb5LTPFpg2InaeZXebxrJxhNkjJj0HPObVKwnogAJPkku
5o0cVclBvwhN1HynS9NSlVaqLdOg9PEErUJshliJhlVapQNYh3mjK1gF0UjcUXhW
jJpAIE0cfLfwtLo1SZPevOVPisKC9VNRWaAm/P8CWasvSYPo73ecnDEnO715lbvQ
PteE4cN0bAFpLcg8ovvvA7UriM4aEwct15n1QFDHier6S3O4xEqONhrGJB3CdgCd
0DKtNVKFW0Nw6sOjsd8KSkk7AA3VNIk3RmFVonwy1FrLttLwYuwQVgyZE5Wwupc6
4l3ZEqqEJhnUYUEd0jgl3h33uNfiA5NYzhh+qHNAijCCRr6ZmR8zaORrdzAcYove
qGEHmqWm5pkhv0ImrNtGvBnUaq6ivR68vYoEKykC8RIol1oDKd4gwbrCfu28ZDG5
sr/4oLnxdtEqMlTQBrRg54EXKWC3nHJWULnGL9lcwV57K/zMzf/0Y5LwwpN/+Ffu
XI9cy2gFUU7eJYPyKxiykAYnDorLs1aExsbkct6P+3dy0qOG95oquAteXephEcUD
IGcOEFCoy2bcqXsnLmq9mIZPJe/uB5LwMYz9Oig6LFaYMWD2DOTgsQcDFwDNgu4L
8uX2xTMuw7b4/KGtkPXVQdYu4FpnKoHkD4nBKE6f2TdmGKtMS6Ul+HKvN+b4KV+p
BSOX1vS6gangQ1H1F6L00SuXX+tghktP92GTShZKjuzRJyH1Q2c5pDV9NY6P8Bwb
ueFS6zKt4lkPSpySl9/iESToMTT21yk4Ngw4E0FMtGbi50Pdou/MwXhu2S3dFvJV
igJlKE5IwvMpUw54w+TH06ReinYJ4JkIUhNPBPepewDvUqjwrcgOlgTSzTlJjNGP
tet9DphPyO9Pr3ND5pXH+Jqk9NXrwuKMf5xLbOYZ8Wt8KaSsWkA60M6NiFZL75B3
Mv9AEvvdu30mqjLA4LLGkgARSvCrCJ+zme644LSY5pV4hl84PCXpSYOkNWVX4+cC
t6o69viyqoQMxFmkkEaSVXk0TfI6fQVx5/OrFp03uivqc4jblWDU/D/Us2R7izAh
d5LJKUylRmty4RJIGI7d0Q05b57TxIdXplL9n/NlWg8ctWjfi6KSsgBqXVXTWGVQ
DM+7HqPaFQFBl1e3rgEeeK+ll/M0lFRs+BR3V0sSYtAy2EbF4/Bn6yMTibdm/bOC
j5B/VvP5zBQAMwWya5X3onYVRRNQ/eTng29vlehZN6sLOa37YbAjgCyevJzRK6gh
L6dtqSCWCSHS8GRCGpLVUmbidD7I1uAYOTIxuNbDWOKgKrgzSkwlu+Mt+C1Gh2fz
5fJJn3Yw0TnAqrNxBAqpWKQj7rJ5q7ourpRmTEssE3PKWe6A3xYjjzTHBCNf+2x1
yQ+Xjzyswp1vg/NHS3QbOQCvrrdo5g7y71s15RX9iCxJzDBmSLb+Cp5G+3VUL7ml
SAfSLG0F+flIKxuNyCaKrvBF1DELYLcQB7bT5Cvhlpb6l/HMgjVHZkmZBGPC10uS
svlXW/87t41qkmkWouBSdtZam9rxfxs4Ab96i+wCmBYKBKX+8Aacvbi735jQNN5N
RVhvZ2td7xFdGnT0GcALvk3nSsNtwh2NEAWq3m8eIJSGnl/ix6ulry7zpCuFIOxd
4N+y0svS1Hu2NYVuzIfAAevOCZdRGWhoYCXyWFW/2aTUVP0upThzXVwEJounbSpC
IApP3xklQwG6NyI9WQmZfjGGJ+KvTf6YyKUEfqGOvBxOtzFkoFzlnm42yqJDIDHL
7OVAx1AAwKwJbgovG5cddI+rf5s8yc3nrqdZaJoOXTvc1lNycJ2pzcqzpMDL3tfg
uCSNFu7kket388TPf5+wucbpPUlRF2fRYh8sSCMKfM+ptfCzbxgY4az1IIavqJl2
8qy0C8F0gqPtDkVH5VK83Br9bdCQe0gtqbxc5CzDJsmaxeAZB8LJWozjfKH3s8qb
sct1MAn6K+5LObRZlJGR4Ys4gKF/nD1p6LN9e6zZuqafFpwjd8Oa8xBd5fuoZAzw
zaOztsVycxT9ElpLMCtCQh+R9I8NoUDRg4oNR+TyZJn0syRhf41KyA+aGH5vcizY
67Me9e1ut57FgGHW90dpHfQ69XHMyFkP9USbMvPk4qmCvzW9NYj39p76ZF8S7f1o
UH4RrRDfTjP4lD9mu8AHHohPHAHwWg9su0coIH4zcI/ONbYXWMSRBPM9BGUeUqny
W07c+BpKEdqUgllkCiZewk8pYpHS9lXeo7ffERmQheFMBu+8R02XMbHAoM+BxjWI
7wH2kZJsr4SFFYgd2m2RsoKNYQxxjbj6uFS38zKi3mxfx72jVsjV+uJNf1x76GGW
sMe5b4aIIa6zXeVOlNAKdCIw+ZELTXTnz25v8xwEyGes2BugOEmu2afwf/+HruNY
4JwV1aePkP5lbrZgOrPmSFuppKSoZ8zBHeLrLGxM9VyA+71elbzjS76zcql0H5ye
b6JeGUqKvFCl761t1GB1dU/CkEubKz9hF2pN4S0fXganeh+GwJ2+IC73raal8WN1
QRB80UDVPcsAP/+OCsf+xOTuByA4HmkfjmkSylEgKQMjWpclDbE/spZptvy/yEaa
bCEPbDaju3UcNWZMIoQmtXVE4PiTOdfBfsS+1Dr+x9PjQfQ5PzOxjS87qgU1Uwbv
RpTBSzSZh9aow101Wt0FRAHtl9oSebV3CaIOrnCNPR3K7s2ONUv1etWxSIaHvNM7
N5GOda5UQLJfY3NizzK8/9jgg+Xxc5T6hE+nb2sWq14qnue2UuqHF9iGWHWNdJ0k
VgOit8xY2pVvGgsxc8Cm4ZG8Iumg0q4s15RuLG+g5Uvn2tcjL/rfaO4z4XF+5O7q
rhFGkZI68gPJUgdTtLxvD0x8NPNocuA+3PjiudW6QjArvvB9eZw+aPTesTuzfRjw
fXDNJdjGoK8bfaOymKZxtK6IGhL0us+lnE1lxm3BPkNj6bo7iyWW3a5kBoOKkz79
JDUe/G/wQ0jXLm3bp7hBmdIpKFlnwtauuavInMCz0LY2mGPuNJ/Gt20ssjE/DANn
NtriN6I16A7oVKXpx5sFXalNKkLRiwMDmoGnNZbniwUTNDrMu56okY736di0x8/p
sRx/pwuFep29JzSNVQcQTFBoDdYhuyxNJnnbf/SHnfwh2AUVt1aUGN5BbQ5SGXxZ
7E1hrNiIiP+21VjpUkgjk1EZoe8qeUbJChH2z7xNL18rNqAlDVnl1LrypYAGdshr
jjY85KUaY4G9C/7ztA0LoOjlTrFAFlpvBay8IWTOzZ/GqduSYzEGtusU/4EIQo79
WnwytG7L4iMlguXDZbyrn4ZnoRJCLo36FqBDYTwRhGA90wL/deh/SY3fHio0EliW
ceFJC5ldurRHpzYGZgbBlBjXl/bksHZwJTVeZV5Ek9+1od0+st6k2Cxt1snDO89i
xSzaslBDCT7+p25Mnfu1gbuGlAwn5trYU1qbxudTVXzOS10ZFA/WnVgXeLB6BEMv
is9cBsqk1YewDPs12y4SkpgJCmgHle2JntM7gs2Hmwoik0Zt3G2G1tUz6Q//p+j3
O7XgELTFIx2XHZ7TL0KQggVSyJ49OCdr8S0IGg94BGYOnFU8JginTE+u0lInbcW6
7hu0FYJbYFRY0x5OPT7QflZjUDpdkwKxGMYjRRYD7BVObRImEDFkQeKxSMHtLuW6
puF+zkMENIW/uLZDZQ/+8aJShjhTpy2Vzwv42Ya1wRctReeqgJNABn0RJhQCJ30j
BlekGb0kN4rH9o09m07pIuH4I06MC5YWmnpBMRy4Cd4RRxjQnmT+FhRd+l+csE8y
RRPL2XgPShvSpzV/LrliknHtjXb2DNYBKkSW3xa0j22g49/2v+oNSzoWhpHq/88p
5WuYzs8lDx5DZaIHEqpJidQkhQA6RS5fvHHK1D64Pclo6GJ4Q06zxFr2Ahc1jOoH
+6dmHbbZhMQ6+L2m9yzMmOJ3p8Sz7Vu3uQTzHeF++sUJ4PenxNVW0mCAGElnrVUh
sLtQN2PaaD741H4hDmE9MBIHJ7CgWB/fbenTly62Qo8CFumv9rHgO3+Z2xSCvPZV
Uf70mtB+2nWH7w2eSYqqY9gAX+dRuQYEykbhQayDfz/KJ9svyoU2Nw7F3j1+4idl
rPqazIsnkln9uw5rQFyeVxtIQ76AowirnZFdPhyzCr21QKUyomQNEL+F+U/aS8va
jLR67oAr6FEl0aY/d1kIlHP3YWzzqyLMeRRvtbDm9sxoGhpOxkTrfjIseYMBdAga
tndXW2d3mUESzd6yxggK7kbVz/BfFPbail21ophcbn3vkCNdg1bKSZxku0ttz5Hp
vwWihVNY490MIN9gxq3YhO2f4tn3FnTyGe4VOxk7yDHdEEBkps+6O2u95QOtvZAd
4Gdiu2JxIxg+aHBz9P1DI5Tprh/8hJDxSVY25cSAoEC49pTr9Zg+hlPLGxk6MUab
omjF1hZJho7r+Dwui6CfgMRV/6FxqDbAxTk5g7l2GtSQ/pT4WtMrjyqPuU29G0+o
ZV3LGjDse1gXVyLv6SGqr6LzXIXQqvdlGZ4GZKeyT/r4T0TVvLEKhjB+DVIuXnyx
KgBlrqX2LQJ/0QVlZy8zjgbbW58KOt5ao+I98K6MZP7QB2KpCMeeKItO3UheQnaR
Zj0PvM55Lk3RnX4xvfiwZrkLJnDpgL1CE7CjtNCyxjrGMGT0ZUzcEI+2b+00KM9L
3qJXNeDJDX78sp7LdMz0zBfQebIzPM5IohzAcsHZ7/yngACvYCw4/YHxUgs8mlHn
llhfIkkyjrJNo7Gck9NWLjhDHXo6icvx0QD5HBmNghSsL9LlyL3EriZyxGUpWJuW
IFE0D9YNlDx7q2SGmgQPwIimoIdN41yba7NM7WyjlMK3FAMxYBLVWubzMPWalto8
gCycmvAUKyA1K8EaSmPG9QjOoluPDdfqts6PdMiyrchiW5SCf/H1wZVFYkdiIgDX
SO/XK9+EdUU2FDTvGEhNIt/xU+S9oONz3pBsR96vuIY4SVZK3UeDRJdCeP+qiSby
W+NWjRpCv74K5qjEJoEStqOHpJ+Q0KHisElqjVyDztb5rFXNgTYovlcymBZESo2q
QW57BXrgi+C8CycSe19ml8QwFAVXsAz4RFv+3bInQxJYhHDe+N0N8zLNgD4OIKnj
pmZDOoMz+K9LeXacdzp2t1diiKfUHVbOS+e9/pihjYyGib3PHVF2SsKmPZvoyRbj
audcRU+HkpG3zVI/MmUL7INdhGTiE88IjDwQ0QdtYNuY72CYUsjyNxMUnjWVR0CW
P7xtJ/8JeazUb28FnecKI6mqUAhd7cukqT+Vuey4SlDjH1358aXnxK1MiA67+ydD
OrvUOpOTIq+TrcpusaXYCGtsBFva4julOwSA4f/hY34IZxixfgUKNnw2rxknGA+r
p71uCXBUjyQ/3Dhf+JJc8Sp/atDNF636gF/Kb5arp9kkv9MyfclgcaILACyQdhw/
5RcoGyz09L6h64kcLN60DO5p6KnbgogOSFrELLxvWfSTlNa/9x647RWz9wmHjRXJ
XyPNljq2HQYPrW4ZqlUGnvNNK0t58GLI9uR86QSSOq8rMHDO0JororQC6/bNt3tU
DD/CYbWuOkjcnpVW2apuabHB7Vc9cZECGAacQrGv1HgNxO4ezthfXYnDrtjTaXgt
GLZUUZuM5HxCv6Et0I/qamloeUl8VI+CAv87PE+TDLMmZOAwztdyKZoD4c3jB+wp
4373+QsSxLiTV+BEUexMO1sUj4AOxjwqRnj+CS9KmtqYFw+CDem1gSovnHfu3sqW
iBhnr3P6q22RXsZOF62QpsASMfvIgLeKGrdF27iwubPObC8Q1v98pITY90Zl+uOF
tI8FoYDsI00iYQABFFNorEQ03X3B6dlXhPAMYjt7LdzOAeXn5JKPyvZHxByqnkP9
2W1hJSlACz/drfxvpzXLPSKEQwFf0J/qm1NuiBHdgDlff2KyqwL/1WDYIH0+EI2M
axSn9FhAc+0G/cY6UBoz57lEBklzoGvOaia8FwVPXreP6u2G+AHInhqjCN3/wAXQ
rDj9Kg7S9S1j1jaRMZMeHoOD7MxgxGzWYfgpGTtAyq6eXPGsrgL+JTgNHoC+qK2g
/qGMZGMr2DqzXpE8rWCnYg6s+W73HuR10egXm9wiOxqaDCe8ExajnhwcpFvOBccY
6hE2JF8UIBSO7R/jxmf0DpzAFT5IEiYzftZZ2m+5bImxtWYojIyzSzZNuQgr/QEP
ek/j4GZE+JqFhktGx6KocVtQI3PhVvBQxLcnn90sRXrYJTkrB+GsYWKzhvax9dAS
OyjiDkBglo3qiv/lWu9Kps38JBFNvZ3SIPOUSa3si85HXE5a/E7jh4Jqe9aATVju
wVSqrj5n3fKEGwdg+9qztn8YuTpkwFopXJckSQxO0BhandqZoSs0U0RufV8xbvCF
zX1ZBeczKav9mjrcfBGEeMEs1bdaWpLCauwa2eU7mbG2hKuophYwadOKPt7owiY0
qXGa49EhubTaf89XIvSYweNPcOOuqm40SQU1FmiVFCmj6O8XTQm/oVjjRQoYs1Tw
+m6d95XwdnGs34Y+62f+gZIjTVEv1LCNKmJUWS6ekJok+2NcQ0IH7hUDtIWp3MTM
2zc2z0aS4xd925MXV7vp3y4hXS1MvNua0HWvU3qecONEWT8l71hFBjtZP9UUqRrq
wWyvu3TPc9i70/qHuv09qj/NlkPHYL34YjnHtNBScjGAQ6GK1oofCKkcBH1mq+Cn
xbf72obp9IC/4p5wKtMNZ/HfPY/ky/0cyqhfD0APZ0RYPeOTBs/80MJz+Pbdub+s
G8y5hGTiLTSxWH0Nn0Km1CYTJFY33QqH3w7Krxy9pq8VcEmHK6KmWeOw0+iKznMA
/QIfG71h5VbtQzd8Pw9l0DZFIm9iE9vE3krHsOlA+E0AiBzHcvzrNUn224AomFyo
JRM/HZcz5MSPMGS4V7perO7MycFFtPT9unlCULjr36KHjeHUC5uKJzPBnnoW69+Z
HKGdqRb2p2OXKa3MuOT16YVH2wKBZa5YBOS6GZXobAID3hEQU62Dimbagve+J6cO
ww8iluZlXAeKywS9DSZuN8tlbx63f2OkV6f+cV3COkIXfx1UhKZzLq7yfOvwBIMU
oiKh3j2PYFkEp5uIFLTcng==
`pragma protect end_protected
