psl_gpo_inst : psl_gpo PORT MAP (
		datain	 => datain_sig,
		oe	 => oe_sig,
		dataout	 => dataout_sig
	);
