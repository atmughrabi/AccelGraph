// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
H6K8bk8DaN/ZKKa9k0mWAS5asH5eY/soxevkp108yf+h9nOepfVhCQTnN/TvTe4K
gMJTh6bFHzozxy18AX2ndP9jadE++qfLI9mpMI0s1zIptzBjEE0lF+JB00IrfNCl
WpWwB9qpJq37aAwF3CgZX6h52/iyLNb7wgfm7cFUxeg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8816)
iyrXjRzCK+nng8o3Sg6eW1632G7xHavog1WO5w7hWGZxIYPty8Kn4eMXfOJblmUs
7/atmnIXFGNonYlJsUVP/bhhytRVN/bBg4n6poCxpKUmwp82LAKuxvDD9G+AlEhp
IdOf2+Ex46k54g0L+eYc5hUOrMaCwAG4M7k0aNelCzlaqOod+paEOnOqjXuULHQE
IQmsItSr9898jT4mPQRjN1/v08/Q5u0CxJ52zZhLlwX9zpK3YOXO1S+A53PRH5S8
EHDSIwPK2QbEPipkGU9CPW6N6fogEGA9z7JB4qQAXvxWgyh9hzYEQNaWPgPAQugc
wLQqnnaDpMRNig9iaJs58/Rl67vCNW0xqayheMTarkU7+ghuTL/DdImNC5qFBzuJ
nBwDN+3MHSHQlh/aH0xo/BX9Lz8XSsmBUc2ry0egRAf9oH6vER+F660iO7NAB3kU
KZt9dEJZUAqovKHP5ikLTW78Wdgffg+VHKsWuJCjPq2MIYwhc2wWRrJHkKo83cYx
sWwZSNI1mhtahsFhlkaOEZiVDp8b6UnXIMHuxSuXA/vMLOliny3gMq7NmSFG9q7Q
zETGCca5jKLAIoGalvlXT4bJ+W52cx7mhep5Gnw9oFpYQhYJ3BQzoB4U4/8U3OtW
H+TgHDJAZj4qe+FC7RlxgqLfnheLrt5kqeECU8Qo5g+zhIxfnFF6XhOSkz7fdzGg
A3T5AgNUoOZqwy6mn3deUfamwu2AZKK3DihvMLZbUyLC2nuzkVhhCuPZhMV8Y3gv
cVVVLUOhTZR89fZpGGQvRq6BLHTO5LoMs9uTguR1aUvpf4w5uYhRobiLb3nlwZv/
jmdQCfHU9k3z893N+tfcef6FjKXrAGBCIRbCLW/dFCpGxkqrpT1OZMn+opF3uE0m
jil6kbZ2ZHD5AFCaE/g2c+krOrHt6t7bJNnF+GXBdJrx23uDuZqCBMLmbAb8ow7+
i4aljkF0vJpXNk4UFAAoYbe0ODFZhlvnOFOJTDkTdYwhEkIK+02l4/vbpBzI0xCm
Ja65OG/EB+PEyzgt0WtwcPOBxn31Q0UY8oCE95UR8U8F7tF4kIs/DIe4IdT8jg55
TI8iIXRm6JvMLZTBVXBio8ZXVIFU7/e18/7ML1SAIpbT2XpC1DH3qMKaH6jN/0R7
gUZyXGvFPyyNldrr8IpcMci+GCWlL+ER4cmNsFJhCxMHomjPpiqF6eBdSqUPWGFR
7/2jgVUi0Eo+UhiPF1ZRwgOWiCdSGKU98Nl0WvDZt1wWNogFE9lxVVrMic7CyQ6Z
dFepsCum1w8+BK7vmewC5o/zWXl4ojkvfY2y3rRe738mahaetQdwP1VlaqF4duUB
tHgBYs7jBHRvOHYQtpsKP20CHqv/M0y97Jav01v+q1SUdACp8IM2LDtkQ7bFlPLV
hRBLTrYS6AfaLflFQcFflMPtk0ERENF8mxoT8afQomqru7W0aL5ByeoG3qR3tGth
Uk2xPShy5ZEtxoSXQUnwDl/YFwvUTGMlY7MUuXgCeQJHWT1VAacqDT1hdgfZDea2
HbiZCDmVm/ifrv4HmfEw8vcnIsHrafrikm/NbrzkPju+XyXCdlvoteoQPaPP958u
XFsFheL1iTf8rGxK9d1pyP0T5ZxgB7PJ+xZfXl6fmi/CHKFXdWB/ue3mm+3R9gti
3SrqFxymYeSPMLwNXCU5B/liYKwM5iTBbpZ6oK4ON7kPmJyGmw49NVcQkq92wV83
t2j0mrbl3MFGSx0O3vh9/d8Byx9VpJUSdD1vKEr2TjsmJjqZHKgjNo1ndsR+/vxD
q/YOJJlrKPCuZ4MGVNhfSIQlkmds2lLxJyWEJYGF7Gm2w6wb1qU7VYf4YWrQ4gyC
JhJqMgkrKxohfVH/sb6zcd8ZcfFOsBbABwbCNe7a6zsv7gx46c2Ktfv75y90+tfY
7H9Lh2pAAsKJKUDx27engPErSk9b7D5pnmMIqbHbODetniS1Fjc/l/pTQORSYvhp
5KrTWDNAlZCOfq0X/ZZ7tDqr9StwfAomD3/HnSpCfKFk1zsQS16wWbWyYKFRR0zx
bJ+T2fqROzUfmIxPipqO3pwvVoLRoRaQ+reCBh8cbAjATScicu9DZfjo1YuUw72B
EicvGlaSdW/JgM+mivFxhzNzEZ5InjPCMwcvEi+MntWk8LUJfELBRUS5kMUaT4T2
JUbSYdxwizI7Hzsuz8yI1ZoxkMbjjbk3jjWW33UlkTvdVMDCN7B20122iWtOUUJk
LwKMFjKAsR4h5HOUNDJV8fsIMmvjvhaL6uanF7XPy/8xl33EE39Lcl6cMreVerXD
OSe7t1jOCtWjnwqBWZVPTlx0WJaNhAoMxDmBIOLgBJ57q/J7BEa8JaIzve06AFbf
K7n8WQ9SQVWyTvvqVmKQ1KMvLaQ4kIQZnHdIKrvc1rfSs211WDCbOLEjuHktzSnx
/XJZ+DmAX+Cff09LM4r1MgOFgv6VXYg3KS/1yKB7Jaimb8uL+ryUX+Se2wZHMcvP
QnwZmz7KC5lalgYkrtogZfHYab+/7ThifVRm0LQYeFUFzXWe43zyufH7RSoiFViq
8fQ5GGviJcvsproUTuXLzUU4CdhEZLVXVNyfgLmZrJxAQEnwipT+5bBhtw0NJ0S/
F58+LxX+7q/utx8O7LG1qp+bRpUk4HE1zX5oA3G0i1Es4h1wEbFrVuDof9zNt5Sx
7XsBfd1yVsYo7Lc1FyFA+m7fzGcz5Qz80eQYtjrRlXtNFkkDUWDy26wpOtpMWKGu
YmE7eE+39uI5TPZIBUbU/pLJeKpBkqm/9gb/oXIQ/fSuhJZQiv4IezIoL8OMvtMQ
aUeGKJyekymdAN8huYcGGdOZiZ+Wt2/vkUGasqmoJVgEK5JL1VaQjd64JzrhywMZ
wfr+sPM9utgfDYX7aMsXG4mPAVasGGChRKmqVtBCsjUsheaINNJVMyfTpQcZnF8V
oo6938VuRHajJ9b0qepL4qCQR+YXfmMRHpSZA/B9KoUgwkvy0NMhbflOvME3mVyO
7Er7sSszqgdHFR5KZkslYY0Mk3QF61JU2PS6od4ropfxTA6xAg6+W81MJU3gQPtz
Q9V9v2bia9Y/7Fg656D0+TqWh91lsBv6XdSSXXP6wRgYpOJSdAYiPXBmRhCGlKXO
4WvGOTsLzrbsUfIEThv+GH9ZKU0iVeoxO9Fvqi+zpASdGxiUfQybZI0ehRTlGrtx
Q+t+Hawsf8GLB8v4ENXYet3lJ5OPN9tzYoMhJX4y8FGI6o1U//sLTr+vGiV4YNl1
xZlsdYrPbol7NKBppejs4GQ2cnbmeLGofWk+3hPMtyo8nQkA9jrzgDllyv6cB21D
ABfM1CKYXDqCqqw3VskY32VyUynBDDwVGoZuGdllLu46XVaofK0227KCDXavy+oh
tAodpWChLLqsUEzozuhCf+j1IGeLIg+EUk5JbF3Z3oO/ByrfE9Oc4fAM47DV61e3
C4uFCxlV4vvbmh+nxs9VQGkfYcKtrv5aEDERFrCpn9onU94H6fZAy98DLdu53PwF
bo8NO1qcGODHIdz0EE5Ckb4y9ptm0pB1GaZgDqqjX1veA2Emc6DxCtjz8uReuBmN
hLxn7KFiy+fQmqdmWH/GjkPtDypnVDbJpcocpRaqnDMPE9VCLL8PSXJkmtqtSj0Z
0/hyJm3pyL1w4dFtwWZoCgPvWF10aGySXpVD3jY7HSSBZ8oKcNuco5z8Ina9IXyG
JmbeMOXM6h4S2XNmHkMzzLojJ7B/HSrTQ5beboh5OgAN2No3K7879FQ01ja6kk6a
AR5Nkk4kT56VSuZOOUCll/hI7pjJfoZuHElakVdxZdXVuXJXuqK5rv5xXG9HrL/w
mLnqZJIvYUP9KO0jZ/jPlEwvnF/JJRakLsXMhFwwQ0iIauv8o0sSw1XcAciN6fQP
SHhwR5ehgbiAaAMGwjzh3/9t/+0N+c+Jds0Y8j0/40DZhXVtdmE87V8EKk5wti2z
RqE8ZvNgcmbTxgvmvlhl2T7BuV94s5tRTmpK3AIgXezsLjFBe8ceAQhcoei6GRXZ
SFwtgqg1yy94BORQNTxUvrE2hjHhIZYD/SXhhUkM2MAo75VqtVJUUxbjCriOa696
nS57PrWUFA2dthnBDa0oBuPTdkD0HbJPg+XWZuJCsp/Jp/zfsOVtmRAgN6MjE72s
n6q08Wj+tPf87sfhWuOM5sqI9AJnKMy6LfhZFT2c3TfMPifAA+JwEUlsUShpfU/D
b4TEitKXrHuLxs/u4n+wZBXYGKjR0bcIgKuNujnBIILp2OtU1WKS7XKr0/lN5E5W
j8mmWWZa+/fAFgyMII+JpZ1iOTEeJIILRadc2h642mpWO7qloTKw9+N0R9D2XMkQ
rysiMEpVqL68a/CCzMROHhMWjA7thxDT8exQMMVlNi9n+lJ2pr5I62ABom4ihSk2
HG+gaul5TLswEfAbX+lq2G6cw3kkSfIufisdnYj/9PDHSxxiMh7XQZkVjF83KXmS
+0oQh1AUqdHnDH1Kz7pHAIfBzsLhKQG1FbiB9j1Dei5rVzD0k2Vwr6ueNZCRV5qp
XPYDPWOyisFuftlawL4qML1rFqNKiK29X/sBcuwMR6axMhDqByfIL0OI8REUI8zB
WoQvOVzBvh89Znvr8xuDN8fUlcA2pIVQoCMF+yFljcfrRSaNWQAoqTf4az7wi7LH
Vaus/VUf+WtJ7V/Z6R6FssCKH0u3eYku9/Owf5fItVN00eUXZCYxyT9E3k2c2CD0
2pMLqkMr+++IsDoSGzK5sSKcxwg77E2PIHLQ2vPguWURNn3cFlUz5QWd8wg4+XaR
gAGZv9U1Yb5/WOoSQkdHzqINGB6t6FKgTfSPZBthIasYtYp+r6M/Dz2kDYI+rNrN
tNcCo98QOwP/GEtQDG1ixc2Sr1EbtM2zOJTdYeddzbdfIH8zSa5mFSQxIunHqF4Q
BiXX7dSD+fEjnKXnUK6mwoiOEcCR+wdtEY7RPXluPQTTGx0hL7pcjM+5s31pgUAT
ibVgyvBy1CxHapAW5ODF0ePLXBDKSUYChEz44w0+BLufeKsHm37anoGfizBb979N
hrM0BG0yXIR0/zI8wyvHBHsJ1UdeDGzywXqjwQFMawXm71R+wDTK4CEyw5Fl3ti+
Tf5koTx7Uw99U/31lQLrrgIxTVzJrg4p2e8EvAOUsCQJwlF8GfP0nfD2rCA09Wdw
w0kEedGciPqmAQ9ThyS4fQ9rgYkDReOgjHJjlzrsyi+LIxc3249itBxSinmufqKD
0UnoMei3M1eTJ1TMbUXv8BcLVu1QGxFrYWTahTuDyy8iiUidfrj7w7WNJWFwlwdU
p6fLSgX6imzotqk6XDL5Kiu3zMjKdxOCSW/6Uz5WMxN914iXa+v5/BgpmclAwUHO
fN6W8LdGudfsbI6gkY9EEOuDJhvU4BFtKtAioajQvau0LJLmM101yZhTYQcV98YR
4rKDC6f3i2K7bGYyCQ3KD9gI0doWIlBtNv4+aXeSCCAD3I3bIpSzIVI2BbAQ14fA
nEKWgNfnOoIHljDPQVQmtlBqx19LUXhFQYByFpcGDKsfHRYBz5py3IR0xsh3T63O
ABzfau8fZpn9oIptYvFKfzDiImvY0c6NLKsiT111olsU33ruZtH+vdxjeZ5jes2k
3cw+WKt/Xl31kZ39au2dRRyQ3u6QE7vy+BQ7FA6HN+QRo9viX+jB0aN012CLhnGJ
Kf4eBWNnNxPehngz4NwVyqbcK1v5cK036EsXGsGLXk3LiSMgVaWwddBqBB1lOXf1
azxdTcMUOLVWMcGjwX7n4FprhU5T7bD8p47NoYGmOhW4t14ldMBouQFFf9rTK69N
OUHMy8BhXWxkpwoEGx8e172iSK/xqclkZGdP80DKuv5gnBPixI3TvhIQIVs7ySNw
pLVd1xTzhCg2d6plXIMPzE7d03agPQVfnyVTWqnWidt09OyVdi4nVxYUQeZhT+1R
Uu2e1XgefP0WOMMny9Vu5i715K20crTgQMX9aGuuSXnNPWGUt9khyj2St56u7x6S
6glWAyOLX2XiVMXHa9Kw7cnk9m4lp4dYVkscND1QGTcmGBcjN0oIMGm/ulQUzgxf
H5CvCkgD5IvPwLZIt34336lvxu0CprHM021v0P4cI+dYpAro+/c8SpSlgLq6JY/o
8q3ZefSELWOPE4GfO38UxfVsUYDf1gYn83zwlu4csYwkzybRWopiEeeK4Z+meeW2
PoHoVDoWsLvCHjGhsirk198dWtZg9ux5hQnEH8WcjJAjJ9Rzbgxk9Vkcsh+s7g6y
H1uYGm1sIl9ktNQzbPyCUF5BPeMwH7utYoRmKDQSemV+s8AzVYuMTUqib72O96lN
pOcp/h3y3I3ED2cmMGNK34BGpvpnewHZfBnOptt2h1Fq4moMd5YkQapfy1Uw23gt
8A9GxvSjCzfttQXQ07fS9nFrl6Ms0rvKr+k4LZwFw9sjWkFp2DzIm+s+CKs44Kt5
quLSyObkmNvFNkyf9U/bi1xAnRKurisFRefC0zvg/aOtyScrsa4tRe6J+eQohwXx
9RKY4Bh/dn4KV00RvEvf9MVBaCA16t/MDzZJi9heK/EkCLgTXj2lONBv+WPGl3xo
cEXyFLiVhTc7oBVUr/GHBvTCHWHyOBNCLt+7Y/rGEJX/LATNUTivknLWSN+VlK5z
VgWTNMVWh5lle2d1ls8uRx/ccEh+L8LpjDpo4SBmsW+KU5DbHiSuCVMMQy1ow7m6
SBnA7LlbFsPUHEJmhsYpAod70SUvAXY/N3LkNU47hPHoptRdfp3DFZmZ3ijnaOOI
rqwePRTTFHeEuuUH3xAuyDBWRfX58ZIwDx+xirbzLwBHw2cRFr6Wwqo+KnDMk4Wz
Iglsaz5sSHOtzITD0V+tR+9kWZa0yYPMKOtlpA0EAUIn32S9/WAZvPt3n9r7/ss+
+U2+fZEN20XWF+9PykPNZFrVEH5q7YaChWkddhuO8WYoSuN/YadOOb5FJVtkc6re
IFYBK9GRLQMsGokGazZwyPmxvlupz0YqCf5UGrSlIIKFCDPQjhPm6PWsP9/1aLdA
QTJ0bTT07FQKWuITxRC1Ug4OM2TD+TG1b664AXYGQjXGQ85pjgPoJqzYh4qkrKOY
cGsigHIavWU1m98LNk6JDwiyJlrXqO6NVSdDmQr+P8YXbp0tChxWSWmEtaxacSJh
61Yj17OkLaEakRaBO8b26JU8a2tbVhTSE9zQnF6UOCu3GaTRk7q0SvDYCv+IqtpQ
WVMYcufoxK7XDf0CfKh6mJETMACxRMqo3DqKmu5FfNyVp9yKdZERYAouY0GE9t/a
+dROCYHqgR/+hIrUlbrG7s+ZAzHp7g3QLJg0qaCY0JWBDeNEqGwtFEbnuJXDTbMx
KqlbVOdLS5bRD3PY+dDnzYpLSMcC/Nymn/G22dw1eFQ8xEvkkPZ328LfaqLgh+D1
5V5wLnSFrOiL16c96vtwzHvGsmGUNWRQ+Nb9FUG/crSQ53bqdiorIiHK0C09yruY
2j8PV/oT7AAbjO0syiPBmEMCAgVTPMHHZAcOjQu7nYFms4tn7hHfTt+WbOo/sG/K
HyJKMmwYDV7r2kC5JLfigBb3pov1bdNhk9/IpaZW8s+QYh1CWUez8Pq8nXBvmztS
AqAmFGrs/sa2kdZYF2q2Kw+DXP+Esq2lMq08pKupVKSLzI9Nf++YUxct1uMU6j/G
5H0ByfFYv7CN2EfXbDj0eMVIpiFB4POPChVahchxnF3VglAZKN9HybwaTDjNJe1c
73yxdEWJmdNA2qo//jivfpfd3vSnu68jQr4Ha9Sh0GTUI3OFZzhIk3+JIzXDSFVy
LqHjVl+1ikn/TzT5RgyTQixshWdZRf57CaSwxtJKOTpi+bvbiCb+Vy5nKylZC+R0
EDpcLItR225d+Vbi0bsg+1pwbmIRg6WSz9C9wZLejlShVCFa29Xo6iWjw19nRyaj
ORyLyYqi/hCujw9cl6Qbw2BN6f1alXkNtIWFSPndtB1T4aQrXfq5p2mlZ24Bpt/p
Nd9XwCuzj+AX9FBlKS5k5ZvH047skJEpsqLw5VDkwjHcz8WAoyPDToOwdqukdA6Y
ejQVfSLnr4NzcIB5jkBDNmVKIcyGnCYqlGkxMi/xCMbgBh/iBo/F8Ee/3vAgo128
38qiqF/AmlxdjyMjYCwZJR85dWg9m9Gp3GAvi7S3COcgVpTON0cS/1L0LROqL1r1
UJO7taUdlNHF7FwmHbDgmgCdwG3vesCpvM/uGFWWacuVXOco3FTaXPG8lF+4J9cW
+ad/pwJTWJKbzxIPNRtnWaSpkgRlWEemlHDX4cpP1iFY0Vm4Df1+rEbaUfoZFk6f
hbz3YS0rKrI7Ddfvrcan4fpqhpHBhHCjbok2+202rdhH6k15Ig4V2MchjJlPzIJX
ckjXC0aWmVrgcV/rBWM+6UD6QD+25n2jRiyPBjE0kume/cJI6AOcF/OTUNeoLLO+
j+uCqBQoeICTVpvsP+foaqylu2otFSG6IC90iqiez2H+ImaHhvh4nYP+tM0DDdtR
DIYFhVVmhFEAc36LS56t2q4VNGafC6CPyIIGed5tkh4pD9FXwpwsa2Bu2VLm0Edn
P7qItxYCJlBYoFM8BukSxLcRphYv78bT+HKTXCIBWGIFmc7sraXq9iK4/NFA/JZ8
qGc3z4JTuzrflq/CKq+opahlafIpGCH7Jm5zfPwypOyng6EhwrKqN/cKApj/2Cxg
Nv6ByzgR2tbxIDXEmG890V5P/dJW5KRJXOBW4tBbMLx1J4JgZmM9EaUxZUamcBbt
tWHnUKnNGPMoQFI2EaR3WJjorN89eaItkX3iEttvTRUTFpqwqZ3gxEXLBBareU29
JyTGnVJC+zxnJkjmitdv9N5klXQOdyhd2d6/wV+1PKeoW3koQOcLr16uCt6hzzMe
z4YyGMdlsNwWIuWM1cqsF2SCwM1qUcerzdzEDegcFvmXfAAX9DIgPVg+RK5Th/U9
bw31tyB/FgXXaM5aOglpGW6EEk5AFUSuhGaWR+q2uacAvaJD5RsV9x48I3gk0Sd+
NDN/EFSw8hlegc1F2/6IjqVhkEmDyzLeNMFLDe+v8MfmcakYNhe7VKcHNoMM8/qL
pWebxwPxtGFnVnUnb1ImigiQ+MyRg919MYh2Dst4HfKAWOnjoblL6T6d6M8xs0qn
eJtZjMbaghVKGXJCZ+IQGGBkPtF5Mk1DSC9DlOnx4QekUpLY+QhEAmXWk/VB6zEy
3ulXIpdQ0EhurCGs6c620Vo/5a5zkoHx6iLElvXNXDVFItBlhr560hoND70bgD51
fv3qCAXOF4voW6IuL7TW7F8hPR81gZomGAP/RuAf8ZhkLD6xPZB+o8LWvC9vOsP9
msuQiHmWSG/hbqccBusC3GkOnuFYXUm2N9ueWhiKzaSAKMmzB3/ZVpdIFgEEZB0L
rljTQgwVSwJFAcJt/uVUgeGsqu77+YwqQKMgfbOv3IjXqsxUQkGvOAn5+L8mCVUJ
Xx5Gabho/kvLytQFsCNb2QpoibrC9D6qa2+fp0g9YoY/ki9TA9ZQn+77/9ma1RGA
c2GJ5HCF4JEexTT1P3oFtPwozrNU/Quh+jKriEMOGQUFxnJ0Cr/EAOHXRdfQoOc6
Y+jZc5LdO8OduNLcyoaeGee0A++fU3Ev8a1wZf+PJ0WjTpfxpSIafBhBFROoMhXT
WpDENBds0V/XbgJoWRjWuCw38vMLQoXh9c9vuMinFSmsps9Ls0CaVkAHfe5HRjEX
tWSNF7UZFlHj14HM4vhmXENFmJBrgkRinGCUJbrsXN/EniuqBBjmdu/3bDKdJ+lW
LrSJJ3dSgkOhGTBcLMkH5Ns663wtiVtelC21PUblUGaxKQ33rVjmQqeMmZgXFQZr
sLIBhnazW/MQX4fEdalqDjBQnfKEqSTOHa5NwNxwiPLoHKwJGyk5ca9v1fIM/+ZA
z/YpPN2CKURp4FS6GryhtjW/oHeXB3HhY7pkyAf0WfGHgLKpXJrbNq9sNhuGM77V
/2SE/P1yZ3k5wtBq125r7sLC1RdbcLiQTGJ8kLMRzAAv6rP+qnUqrzLQwff6gs/s
0lm3q7BsLIhl3aWFH2D2vF/vpvJYA71boX1vmd+MDDADlwf7hkms5AcVFX8T6LKE
JJh+BFr1WiTVsYI9eRdUFJ9HB5Y9UzLJl6qoSbN0h1NPAopnR8xSR9NVenuNsQJm
7KYY9a2YOA+VvtJCLwlwreflfoCSwZ6ff8zYuJHll+l67Zj+C+FihQ0vjwZDzYN6
EuVDuCa1L5hACmopBTShEcy5CnLrjpLTmge6SjCCl8XXGdI82d9TsAGYcx5HHpQg
n1d8maCTh9Fcm4sHPmg+jDvnkSqXBkKDcDGan4SRMfkmFYFKzWfHzuJhR48URgt+
mGhEMZBTpyjxtnLzdr1cfplMVVMbYejfZpeRoLLYhf9yLBmQmYcNiruuOZGFyHaV
fTiv6CX68HCg+N1z9zOIaNIcfxlkhyDIzv3Bo+jVimsxTid1mxFcv4jWRhvICqTc
qO3kg1UoFdTwKuG1Uipk7yXiLIi9LlxCvxZzM8MZrwX2jPSjfCPcIUfyi8cNzq+9
FYBqs+xi8he/gDPBoP7RkP7yAzfwdlHkFrziHoI5ahneXTFQpTVaiJ4+Hcs4w6U6
pRBqiFCLgZrSrZzRSI3V7QHrVYBqMKqNXd4tFiLWZdIDtuO2JUUw6J2AWFA7cdTV
VHcpHedmMEIh6mDyIMz+BPULMIBSzoFlY0jZdX/p+Uo9sy/Y+glahBoseb4b+cXU
YmT3oO+S0MA5c82xzlpxGywl14yzxCLSOWE+dylRGwRrrC8Fm9y4SNZUu5pewW0u
eNWt0S++wKkV1JmHJL1omHe8q4zKr0HYF6AagUDWYfsjSpOYO9rSvqmLlqXbnBfO
PyGRitpBHK/FS7Jwh/rty3iVY4iIC6Zf4iEH7j+jilENwobdJN5dQHEsRdjsPI7+
8eubhk8/fW4RfFztVg89xJhxIYIsvniKZGIJzDrumKemM/GpzTiKmqYSXeBc65Y9
s+uU1d2G3rIC7gBb4f69oAjen4ngH3p8B6rNRaGYR+bTo7IhElwWxDWhwlnToDyD
l9mQdCwBQs0fdaJ4O9TOQ5QCymlb5p4nDQlgfIadnC/BcPHkS00iSyAsRcfPwSs0
DejpKlc1W4HlYRyTEW6KFx5GMxYOsdKl/YUAhgr3np2QOb3bSYozx8P5nzITKFd4
ESjLsF5Yfgv3K0cm0xz6YAK+gk2W/qPKBOg4ipkQD2P/wCtp78j7Oub7V3DT36iq
9XuoSKY2iKeXxAPtpZW4svLJFyzQSGzLDIt60bGzQpSFzCVWq8ZgG42VvTIbz8NI
B6DEn3Knym87TFfmgscDj6stmLZOXabLhAuK5aKTmMCUJJCnbWm4TTEoOER7cgGg
BcfSTJwi54EiES7cqlAs9ewofb4K3un2ItAt618Wlh9JA9Runh0ypWnYBYVxzitQ
BnCG3vXsbNYg5swIv7eDTP++v0D002lG01eot9L4845GdfvnrTQDDm5cVtLks0+Z
+g115cybHw9gLnpLuPwG3ueC0fatxoadSFuCpdepPmhhMAMuUjKQucHxG/LvLNES
vSX0RyOliJbm592GVqn10x2tXN9sCztaoTq5Tn5HHFr3zqa1S0sD89jDAu6v0dBI
VGl5QvxcRQOXaAbdjbro1uEYFqpGPJhw7Os68tv+J2/yHRvtFrlvNYR2wBXVWGiN
IiNLKq8Pf1ou+qynkJOOaopceEPWkTnG2QtEKCw/ztA=
`pragma protect end_protected
