// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qyijg1/H6XXtiCTDjjKNjLG3d+xlqr+LRSUHmSluqiR5KDgav9KKaDz6US4h0jfj
0nW0ENQEVy5GN3eAI+wgSWjmhosS0DjIw6+pLHr9uD9xLrvLa7OCPbcITn4pT0E9
iCoeUFcZCikg8Vee6JX/oXs96LoKYt0phnXgRKCpSMw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30512)
MjzAalfw+f+PlPuL1dtxxa86hq5gK7LfCq4vGqhNpKIKwyMVY3wSkMJvfqT0HCGG
Qbfo8q5gwx3SsnpyhrwDhNfLOKnpOZ7J5vnd/jMqoRyVWTyKKhGV58HP/HfFs0HU
pcT78bkPncf4Xum6kcM8BNH7uCIX98aZRSpAMUKYba/DKxAMXZDb5v0HTOVWs+UV
RWDVaLpq3A+xGCKjYZoApzMtrF2vrrg5lLbknHvZWgya0bYYl5EP25jpdJrHgX/t
Htqe2uCvj3M+TB96KxOXNPMR0KCK4f2ZRBSoy7rcinvvmclFmwl+27M9lhijXPwK
EbkVRDUg6b+9zaeUirsUpIHifO0auyrCNTrUZRfb2J9EBqj9YutuhlJtO7mMkX7X
uJD2NLjycVYLOBY1lCCxOErJr+akpiNFfEcr6nSTJKMRhFaKTO3WTIAmxKksuGHD
LIOMkZmNk3pBKRHjMKxe/RzagGz47blBQkBxOLeum2qOzxB+w+D4XY7uniPuUFEk
CYzztgWlUtHWuVTQ3NBilogBVtutTeeXfkemaSh5GCHHTMkt79DR7jBNs76yxvAu
G1ztLywaSWtjoVoSESlnFsTyF/de6z+7QfHv86P6yCKy6ovgfB+rANKuRGbyWtip
cl4XxJRIB3uK0XZMQ/me0yi/NbTMI/vf6h/d54lFRlLsnoEu+XOh3BcjzJjFG5pk
QIksRvysIZxu3qC5Z8FnhL6bcrdzPTRfbDwiBBampdfFYtGCuHcP25DPDmgpcwB1
mcIwpBgVOAZ3OiazwTv6Wys2wfpI+lGNqQAY4T5k/stOVk4Iw2vt5fdqcygFP69M
37LkmMgHKY2iNj+3yqH5zn5kNf1jDPgoK+gEd8YDi4x2fIxb8MitMzG95fGDPrZd
exPhwrefxmz0IZFO7AhGsDDJwA8sFdOgJuEqeqTapqAixqciYYyMftXo8T13I4qS
Tnbi4hmE8ygwUq7PILWhKIpiESCN3cY2gquPKYqGFrco+vSybxlODbsAxt3S17zr
F9pgCNJUxG8scjgOLJjOyqcei8SDKI8UOkbyJkoiS2bpe7BZxvu5IE+3dGelAA5F
2Idgc0K1VraBYHB+TyW+JwLhyGVUzzC1eAymtCnYoBlPXHTzmBeu0FCB2xQGdCWy
hgWcQlJIw/+l7NjckiHrjLsS7cc0xT8hvz+7/RapDQ40KBGrhR2NG4w63ppom1Oj
4Y+UTJFajb/naiQDiQ/FUpXTdb0/5AKCgmTa9dFr3gnk+7Uoq8ishZ0BJhh855kQ
Xo9RARkh5H5wpdn5Sr+PTmC2x0GDFNSGV08m0C4KvhSQzjSlvP0fRKvnZBs8AQR8
FIDpcBY9B8cS5kWV8v45YmAUG7ms16SCrvwuoJTEXmLx2pjZfUDasEEV23yDdvxp
83iIvJfVjHWQQo5a6cFdjyGUDEa9VFDdv5ux1qBx3lbvVa+LwjyqbyiNGKqT4evy
+XfUgv6EpJocjRoioHYa0Uesxttux0uhaNXll4AwnwUBwcL89sIsg9akS9m2/13i
1rywHawVKjgnKo6IKCc6y7WCV7iFd7TLn8bDVlzef2/MpHtq+dce6VIEHcCTnDQq
MI8K19X9h1nQXVXLchaYy4i9xPDxbcV6ddSIshUKGRvxzYlbc2aURXnNJyM+oGm2
2rU5Z4wq+bhyCCwj/wQWemh9Pld73sa0TbT1Wd1/O7S+AFOIVlWmMj3XpPc5Hmmd
HJamhDeDyOpPj9qY+Eys7ZSJ2JOnmKXFfUV6GN+Ak777/eDQMk28cm1ewn1rXqFS
QwMhK7cLCEHLAoiN5AlrMX7/xQX+C8B9ls7ZjYvMMbRZjTYp3ytrhjsPB60p9xNR
e2tQscNW0s23rgNCGDS240bb0nt1ZjYF3Vhl0ElVDlQBJokqS5z6iAJwipt63Wps
/uVBdqGo7DOxXH9w0m9Ygw3f21q3uobFUSZfWcrJRAUlxq1ElFb0zQlPGiRyDGA5
iz8IQBauRQ65y/8kuPSct5UAfiBa69sdwCiLMdAEWMxKL2TEeeKngr5lclIwwXaD
09IR7/9tp0kaDlTPNgptqeAVCZ9ahSMIrLf4VbbYTIsKkkVdvCOZbp9vT9QfPOdS
z6H06plUGa3HuD9UOh/viaPTGohdJ3ihqDy5aYU9e9FTtj0oBcFrxuLvpoKYsoBS
3ljipqixapdyDWOSm1nImOTkRiQbWZBGJdpwNtgXtmL+SH5GPyQGuIL8z7ag6/03
rqCn0WVN9oLwokMCZY3pLc7PgpJkZPUdxkg5K9hElnSZOR27n8pSruPs2oRG4iut
slVQ+/7OZJmuGH77ohHIyrNLQOLNFn5Ghj8YiKeuv8J1uUAz79JI5aoTsqSAx67m
9OV+jCSb9mWSwgUx7ur5tk8I8Rxj+JWSAYuNqbtVK4QB4A0dM51TsdX3hRTe8jBP
FdPFNwFW1DNXsbBj+YE9nsPo+0GqVEABm5WK6UkTZ3QUBpcP5mzH7Lw/sSFc/OsP
wfVjZiwXqFv78jAwbeUZeE2/C6Oz5AKVKNQKEhGlt69sMklGab8lEv4uPz0lrbfD
/Ho0cH7tlwXV8rHSedDgsxspjK9ubYoF7WObt6bsRFdqU7L4YwL755v6amTW0uKp
aH2ZYHPOweFze77wEjy0IyWVciTkfkotlyV99ivuflQgWRw2MAkeKD0Hv31kHgJk
+yRZJicXrCRint0k6t0iWk65mnq6osGemz6nRcwjXt61c0qhwz/c8ODeqG3AT9Rh
J5+ABxKTxDBy7xi0wkoUjgazJwVcfwudRK0R5VN2b2iOaApvXqNyQfa61iyZ3o6z
MvfoNilf4o69/o8sCpsY5R5KmfVl7w12Am0nWAY6apHRLaUTtcyVkkIsM/jvcmyS
r/Fdvp3sXAKlpp5fWmGzX+9k9nai7tGCW+di/45GercZsr7yXHz2mcyhgCvV6iZB
fN0sixSPaF000/5E4JWHCdsmspR8gwKdDJb8Bi4fScmfgkDgXKvguMmxdj2eOBu1
Nr587UgDwYXujguT/P2RlmEToNk9pX+vAT0sdC0pXClxtmywbwdlRKTowNLPe9TT
1JQ0Yal86T5+o3Z8BM76INsFm3J2TRSZ0k32M4BDD41cFAdycZylqQfw6D7R9QDA
UZwJ/3V0O0jssZfDLgYi7aUvAgS531QsT5w95vr7KWzTTzQ6lt7g4s6WQvf6zWIw
WNjjPJ/na7tCzr78drES+MeTa89Oyr6Jng/5o1Vpgc0a5JgDhqv3g+YLgK0HfSBN
/VSZjIOqtzCTIcNiL8MOSDv70XqKHKeqhu0JpXWyAEYg2yMXpiEKAX1+fTXfwux2
1iJZ9bPUD67Lz6U1DNKSEks7pRHYV6wr3FLdxfk7QQyZbVoovwG/Ecf++nToCktG
Aa54Pxfi1AkauNAIFsGCmBRMhi89leCWdHF+9lFJ9Fv+v5c6fWwtSNxFK6KOIPnJ
RtY2T4LGf1iQcIkTIPa2sW4gmQ+hpvlYCwlPJ+p1wm6cbBh000IGxlCvc5DVV7i0
20+GiqAxoFLbp9xO94pKJILh/hcvjTZGLwxKhwi3PtlwNvQRN8DhxihaxsaNxdNK
GMR5YfZ4lvkYXRZcm6dO/ubbrOPf4fOqE66KKSrOdLWFs9jKBOxROT+mP6W7rAlr
bqnBScAfCCnRQOI0L7nOEqz0KxPUZb9Qd0J41L0eqqP80OH75w4qlXbEYxZnk/Nt
bl/pXfBC+2fTU9mVApcjdH1qDjYryCHz4RidEiMmVdG+xJl0ONuiTWQVQoSxOkwv
21XUyk/ayhNwlQnMj5qN41PIi3wyPWVoWQqgEE06/lNr5d8S9rHBJ6tctKhTHxtr
jC4B3ZhYbNpNQN8mNdEdO9/wfCr6IZRzI5q7U1ZhUqFRB2gpUDUyKul5p9AwBMyF
Gd/5zcsTesiT0CwZkKVzEJoQbTfX5fHZPmKijwZQwjEuQmMZD2AHr8K7r2aibMpM
POVVEyhH9ma5LXMQd4HwNi8XrcVOjs93GRR7XPKI8/+7X9HsEeU/JrMDV7ZD2LaP
Eua/edIJuyttY2EFgFF4lyJAqGOSzsbqVZrzOjAG+py17xGTUKengoQjulnT7OO9
Dwdo7rcepPIqIXO4mFi3bLR7wlk+pGIXlQLY57a0Hy13oOuQx0YmXCRqD8Pfpb/P
4MbfUZp5gXzVAU8mWleFvCKErfxmterEigrAhtYfDKjSIUkz5fQ7TUTKK7+mIZXs
upyzwWAV5AE8/vCSRRVak3bTSbP/r19Yc71ZtdRLJX30Wgqyx4piXUhJX4/ckikU
sOPDEgbL+9hprcJ+Ms4yp8vAXyFCiTmFhLlMvGiCsTqwxr/lSL6klEoSpV/szRfD
CeBVA9u7uNCUwTlm2YZ9uKWmgbMdP4f36td64p03UxCzl+spnX/hwpISfsfxxa+3
qOrojpIEckljZ48YwCBlAOOWT33upHX9Yjwls5LStUkLvYA2TVhxHS5hLdczQ70a
E29BlbFLKZlwFeGUAlWbvFztX870UMy2+R+OHOdRbBBtv43dCDYsVOFe9AVSi5W2
KG4jbM89YMFn/Q5eDEJXSL0B+5fAPbTU6SIjcGpniD0AdWerQZV1Xh3QR9S2SyRx
2YM3zxJv8baWOyQlYbA5moSbAJiLmZOckP7T4fEbu5mIlikKaYplA+caFOkmK7V3
dJ/e5NcSElAABDvQ3i1CXmGlK5A1vQYFDEsxQT8oTbu+1jT7KiKdo5vx6PVoBGCt
G9Ewyu8m0hgV+aJmBy/SuqHtqXOPWwOhpwYmSa1ssjMmwTVUMl0p68LPX1CLxjk9
Ie8BWwKBfrZSIk1iWEt8tVrEb5FY5SGWNH5ktUdK1/eIACISWTozr0VNsuhte9cL
jJA8lu06tjGcmPEgqs/6e3hHE3sw5UNRD+jaL130jsmoER5qnG1Xmegj6Ge0jsFa
eA84Rxd+WinBcCe/ho/rGhlP6+WHEO1J43ISuqVXhzo9l7n9oBg74d7xa7ISehGs
ZakNolISP1fo3e+XK9wx+Pu9UF5rzU+ZZuDXCOZcNB8z2pUXE17Zd7Xq11/iNXPK
ytz9I7NSAcCBGhuPrS49PCgOpEzTg9OiOyOZCevCVEiqxHnd67OQf27tR3Pj8a1y
mSNyfVduDtBknRzLoLMh5aKz34fjZVOo3IRdmrSh5nPkqnW/UlqrQoLnN5DwyC1F
On3CC8AoEiQp8XX6xG6Pm+6HuamUGCu+pXl+EZq2b6kQFbc8iX762FVUgBZGm7Po
A7XbPEWU1K9OT5W1A3fy2SSyRAN/wStBhE7IaA8RNZrwwZgNZDcCoH9tWczAC/dq
Y+z7MufR4zXv+xTfA5vrTQek9R4LR4ri70+CSuZrpcceKZ4FrUVdpST3XV4Tz1XB
8ehJ5kS0enNiNWOg0tlrbosX3sMtbMCf74kqH9RR1Fv34yj/yeXqWY0wGg+U3Xiq
0rYp4zFjuosbDbrbL5tChkpU0vuFa5rdQk/pUXSqDSsA40W2hD+rzL1WNQARdvwr
5nKnjr41GS3+WEchGFVplNQZoAvN4Sut/bR7L5fOuKSwmKjP0329kH/DnyGYdgpU
3eDYTml/4Yd5GFnvRN6MrcNaNeeRbawhzLukPJNOsc4fjwZepDmJeiwsGjAFR8Wp
YIuARG1QjMiEz1kobwGH8T7QGdp/0fu/K6b5PZIr8tXPIGhVpxeT7ur1PFsKr2ar
hZxmiMBQojSIwKbmQTnGc1F6VxV7SQiZdF8b0Ob97dUJ1fnwA0VWG/mbG/IuVaNF
UIoGmJW72Bz+/YZy6g7iek8jsCxQtXs698RHJnhYMATPv1LdMTkXtst+mgBHAWow
aueVWNMF5NHDNUd1WfXqBOFSJ6eoUaQGrCYcWccwhm7aTS0kmRNBuLqyJG3RFinY
DR5MK+f75vPvnSZUmTFMYreT0NZuB+7FiPjfuj+t+6R2YKSo1piaBHbxAlqz3giJ
u+ujs93rP8QCNdrYgr+latYBowoXldDNEmdiaImnoFGvJqhGr/npRzgaBSkb0UvO
KnOVw2j0LJMapN9NG6bL6+BnS6/xBq/B8pBQg/9LGT41PK31iVdp+OUPvGZtv8TH
Yg0JpkjVHbbnNCD3G3ZAYbawWTEfiCGkJ51O6hNqDio1na+5gKFURA/xvX8VGfXU
WkP0p7VvwsZd38+NK2vKZqUxeKmu2MGH/6FCvC9BAAGBKJxRa3ERdYbRyA3pLigg
aoc1TjSD2+rhm1t9WOgGaDwLUmdMWCRndqa+LfrgNg8nX+deb72xywmGdKePQOEB
nQaEcHmp+teJb1NDBXh5oA4CmDrRHCPbCFSHavy16BYyyRqfVwyWMKFcypDQSkeb
WPBCgc9nKJzBzL/WbztwcdKAl425qtDk8tb1NO55eziczK0PByjZcpouhd6kbKBN
ILyLrNEuUizHMLaQpWg0Mn7BrIyq6IYr6rVByTIbOz4GCroDQAzNUFIh18Dm8wti
x5Z4G8Td+AjZpgRylejaY13WD2+yIYhk4hAVfBnw1BhPnzaxi/UV7Zgw/Hvd+7CX
tXGErLm8tXd2WoD6mZj1qiqD0vq1yeVprG+3RNZpDDXxHgrzQfHkDDLFl8EO0+IU
tWrMZ0XBxdI1FJCGieUUO9Zpdkb7XXqBuss6/E3JGipLWhop3PIfsSXN/MA5w7Vm
9s+Y6aWQS2TQMC2CmdRgg7hdmLKT85j5QOwy2AqW2siix/Ho1STATw3hmWK0IVKR
vog6n8jM6KcxN3G/sLS/HtU8QO5W/30E0vLYu41/R0RPOKnB66CGCPs1Y+GVUAjW
8IA0WB0Gmqh1wabhCCH5ze8x3e0z+6SthB9bVD2C9yRe1siHKqwIfmxES5sT5oUA
uQVYYqxIYfue1d0Snr5k4B5dBCCxqvMa/ndu2KdfsYHZL4slXVS8JmWxfQGU9wOy
uCBarxBv3a1kkcq1LEKXKToD2g395sKGcE2Ex5QDnq3pucxflRZV7ysB9pyF2ALn
fJ7FSbp44rUd+PFeSA575AlinK3C7mm199jjhJOqttnIYR/MIrm299mOgN+SDQrZ
C9xICkXhekR1wwACi4IiJ5RAoLhMicbcj90IE9s+aEmvN0yYCruppj2za9GY/dTq
gDXramKp0YcRebrJV+id9bPS+YKeRC8lVQlanJbwSsq1F8zyWOexQww+6Xlvinwb
FhNQCXLm4SsB8SmHNrc4zPk+NIeH0sWjz5zX0E+UWcNHrZaZMMEZe8ACrTL2HEQV
whnn8ErrNFeC7/XFAv9lXGYB/MciEJ2wnmvUgfWyzkHDvBcIwkuCNaNJw05HcROA
90RVZiW6kVW/Su3TlXISPguzz3vSwwGcAorjaHE5EAEt+BDpzeaQLKzajeYV9kG/
0/Mb/RRxItJlRilrA449IJO9wDB4VbUgx6kvkjUFJm7OxVz6Mlm+W9rYFYCNjrI+
8mrR55AzFsR5KA4cSGtsffiMBem1o7Rac6hWS5xHQeF1DaNZXDhlUdztIGF4DDfL
2o+ZEDT/qH4Ev22wBHZamDL/bt0JczdKksU2iA0ExbAKdbSds2y5wQl9PBwJVGc6
5jS4f8yYqx3qIHQlbU4ngPm9s9bf4qiEOHqS/K0IfcXbQMjObP4GCjJCCfEKxx9j
UuORIA26Yp1AfMN+HdqvNHtOIi5IArz6Wz3egmYy8nuoZF8dt/K7yAhpVsAeJrlc
hyJsvefIzKIrf3blQjagNzSd7hv9Y4buI0wISUBvGSogD869f9HUifQHXNnu2tLl
QzxZxrfEDFR+rixzKpBIyxJf0z1zKuGtCBCdI8s3y+DgheGQsBJpd3yq2v328FJZ
RSi9590hcxNoOzqXVQxK6Rrj56gsyFjV7WCdkv9EdI0cOO4mLFXVe1Xhuyj1zmFO
NY/w45gPemWg1w/gUg7t0iMcsFrXGsupxpEqhuF/v3zltPJXBwpFJFur9bBRUirF
bC7djb0nOfqpIoiaHkCplYoE8LpejyhahCS7/0z4lfKsZWIEcUkof9WdnFmyHwWZ
9yn7PSSnCMGgQ0nE1frQ0aCG7PDnjf+N6mQej2h74RLTXtN66lI1rnt3UUhTLTtD
hZSfNRNgQCg3UnazgWAdz8D2xaZ2Dk3GZgroT6b9OO5nA/U2CGloxfLQ7VKyKNAA
uMRxVpxsGqzBkxMo26ltJ4PZTra6XMPtuXm1aCvXorwKEjni5zJE8Tsf/0cEYaPU
GJKJhEpNrKvNm3ukrE4oeDHPO2jV+0g1d3XCk5fAlyKfVpsh2MNR+VwYIL5s3ovv
umpLB1v0iAMegxjKqZBT+rAdbam7044xTApBzckCTUV3rhTMgZjMMkxkcmem9RKW
RINbDafo9I1JmPNqRG7msPRIUID9fh/xlh/fI+fl2054BJiFVqpLPULvhdwTsEAp
3TECIXlIA/5XyHAkeWNeYekt9S14+LDhRYohNUfjBzTIDyGrLlhDSiuJGidAnFIw
sraEZDANEcwgMI3UXCLrSP4Vt8two88y9E/GwIiPjnXTahEUVo4e4IzPW1QB4+l4
aBY1YYNoQ+ADMM5i70kzJ+n/y+FhrkN31pphcw5Hng+wpWBBPMpueebMmmceCczB
DfO3Evk09uFhl2keKtKUUL3QwiyKCJJWrGXKdnI+R1Qew/VwL+LiOy8X6okxkSSa
ZQIdLd8eClRRmvvwvl8SGAIOtHwmGRvyGmLWFkC8Kk7RDgIbhfUwSFkEQ59KLZir
m/nWC7jCr00lrggq+VK9hAaWibV1U+Ar5gNrCWul0N2UcECE5mIREZvy4XWImMHb
5NijJJI20O2hVmB1HsDAbGm0/Ts5q6avxgEQoHm9YtQWb5y/QUAe0d/qRJ8wFC3o
y3706wRjrp0csZIWKsEPerlqcTj8vXngG5YiSt0/EgtAUVizewdwvMBQl7jFtISg
w+uEhEqJAFGge9DO56NV5ONtRWqfk0BMg8TXWGQbSDARGqpfghDWQiU5sqIHMukS
v3Ml7zsP+Ex/hQAI4FbEwnSYx3vKHw4IYyi+aR6axR/E8rkBv0uhmt/II9xy53OJ
wNNr8qat6CtI+pkybpjfBPJiy7YVqaj7M8Ew5080c4emJSjRuiVleDgzNzWigIr7
bw24dLtN95fV+2+QBaCUmLqnOzh/vF7U8sePfz4u+SfF/g4vUfb6PS6AwtYP7KLw
qeEGB02nkF2y8uUfQgG13VgRnvojsnaoGAmFopl5WBYaNVbAgD5/3KtcgNsKFOwQ
MDvPCpSc/2KkcRnaLer/JEgm3QD8yLSUX3imNEMeGpTVwRkmS52mq3c2CdrNP2Yt
+7ey96A/Q8eh0hr/h/gTXZ0EBVkSA7GAYoepc+LZJChYpNZUsTWD7X4TNtRUK6qb
uD2wJmNQiacjoJCfOEFTexEfKl3rb0HCD0GVexDu3oW19nbHzQyW3mYVxs3JFTEa
nb2dNdRgb/4a4wWHmi1QVvWAZwzzxGsTCdIy5NFgA8a9UA9L3OQFLGQVGHpDAWBl
CdnbOaLn9cbXl/9qTsdeh7Yva9Z0jfWfqR7i9wYluxC5bnUchojNZ/AHUST+U1K1
thzikyzlkuynhpRVjSqJkvk7h+L1PCcyp92O+s23YmPFJoRvSOO3JzLqlZXholLm
u/5+/yeWyvmrJb2A2+jDHS2189QPYtc56tmITIV/Irb7epWpioAx3ztQRsONLi+8
Eqm1HvpUK8NYOAZhvYg/F31Knx1q6JwsYGUzaGlM+m/KG0HzkbxPYIwAHBAYUFCj
JhMea6RNVHqDaP/CHitpJuVL8iR9kZ5TBpkpH4OVPdz1i258uRR44il1QWXYZbzI
MZPY0N6zf6dhffxBdVxL/bY3DpJ/oeUYeO1WXBc+yb5jgQFcag4TmP72pQrR0gKe
lz2F9Qqiv6wzKZIYAZejHvilL7NbLUXwtbbF8hxwKgGUMFf8ybpCO9AQVSdlChBB
xKpFrcEd2TUwIQ+z/qm/f+PpdAo5XIPD77oPW9j8MWxT1AFedjFSsp+7LNtVE2Kc
D00VgABE5/QUDeBdj4qVnVIhWRyP093GBMWk9l5E944mJJfAhXh85fMrEfjhxwZ1
g/GvilpkuporsOX1Bwd0VCUGTzbbnIpLLVHzFuJrO+A50oxlJH6g61LtnX+C+Vc3
/6tW5uPBrcG9zPVX7fSJ498uFABvu6+A7k9OUuVN9iHmrmK4jzzXedK2MUEwVSLw
CeBi0+NEySep+kyRLBzZypJ9rJTAva8URZu4utXmUfjFpvZWVpcgQvzLG/7iL9cS
27gsiXd20rhLWfpWcUZU5gFDp9iufSKMyU6wofc7Rt8ExmC0cSl8Qk2vsGNP+WPY
db1wG5BfG2iemJ1OlW3INx5sX2xq3VVGI4iWHzA/qvNEbHxfHLmaBMv1VYcjn3lq
ci4Dx9M0cYJO2/K5l6/JdcuHyqgnk/e1HZ9bLSK9Kagv5Ze0kZJw5RqsUCRkYDJI
08PAhm3P3C16nah2Z+BEtoQQLFWYMLFEeQwBcILsRFJZ+k3IWJ/lHATMiAThhYQD
OwO5BjSKnGT0QO4zp+szwnuHoS6SHsHiCyZY10gjrgilNyV4uip43WfJMGhSvS8+
mClb8Tw9jAsUSiwoZ9W0JofA284BYJudDVSA5aPbk601oTfTpve1ZFuZIyYZNTV6
UwfalgDXzzvkpg6raogo2oWhmLLMhFMeY0ldqqt/h80/mKk5al7Feq5lxcm0Hl6E
7ed9sE4J+4EKV0QVpPivMQFaXydQA7GKydCcK/QE63YkIJNbUsbtpz+cSsz4Zara
2vGGSDDIynBbm9T+aAHWJ2ObX2XMxwNzmEhJYG9d4chJHjvp8k91gR+ytShesOfG
rx9ale6SLGLECnuB5KRJ3e8vpAhmrAZlTLTWn4n+TNyaXgOxiQYTufHg6FX7RVg3
fCDlmNo+17HISaFH5mJsitd5CpzjjrbPMbIMmmg0KKXi60+Vc9bhW9S9QhWSkXW9
WlO7UuYlDNWKUibOph4ptw+w8X9K35qyLadU/kWH/OMLPEuRoLkbiUcM5wSQD7m1
/oJfdWcMUVFfV8R2OQ58PiqxMLEsgDNS5yG1vADbdKq4dj3+VOoQinG/f0d2nAkb
bTASQaLd7gUnGNmYSK2z2LPXbnzuWG81SDu5Zuk1eWmKYZNKj+aqY2pwliyeF/3z
KUtt8C5kxlNg5+mdPTwCh81gfRY0I+i/IvybPoD/m9L/aLH7baDn/cECtOdhVfw7
N7UMyRlXHOxYan2CS3IT6ovor7kVzb0anhcjqf+DpqYTB0aKSYoBAG2aZ7BL+vnH
KgR/xTepGHWYE7CxSE5BcJYfSflYJmTZQwHOCxOU35wbm5T0VZ+aQQXvKIIKTUb+
kn+YcOqaOMHllXbKP4MoCKFPFbrqYvfdlJaLSdZzcU2PI6v6D+v4TBCeTlmRRkXh
xjFjyCxPqXUOz+LUKg5XGYaGK/bOFwYCyfginUssuOFk4bpkhXqM3MxOvpFZCYL8
8+JEQ4plx4xjvW3bZQO2bFAsYfigsjfRhQK7w0fVif598xK/oO4OzbofiD/WKtMQ
42Swmho0i8yGrZpw3GqoHPML6ojhV7KFmYFqbxebSmdZc8h20wFLoubefFJZOxnQ
00Z+p4RFWYhvtBOhtx+/OKFdMEveF7XNXIL+1ht1HnNDSnE6oZMBW8itAIrw7EWV
LdGF1ZzY8y9WLE/s9IHnEb3RgBrbE27KhrKzKTBKWAmcJRVu5+G4q7Vxsh0l8QpW
FqxsD+pzzvKGdFicN5/D3jSBJRWDCRk4a1NKOB4vAnKpn0BFxUn5k1Ca//FjHYgp
QPsb+A2phFoOiP5Aw/B1s0RO5ZxsvItXduf5FSfKEt1bvl6QgFbzMlxZzVXVhhz/
skGteAutV6YSQfCMaFfwvdZF2CIYDq0xc0ZVrXgoBtJNItGnQW0PpWm5h/W29g71
rJ8qHnHs8WVESiVRYkIltQJDU3G0sgIeQ9cZ5SqzqwNsZ5zRyq86XpYrk8pCDw+z
Hofx9yM5eUrBT+lJZ4kVOucNBggMv+abCli6f7xYx0Y23CpC/HIEPDWYqHZAWhCw
mQpyKmNa460vkMi/R+wH+a93I+zX83yxLaunO3H68fcz32zrE5NTxM99LmCXKOhi
Y+aqX0bkUFlU/nKbJ68OhGrnvKaLdBc51I5KfNpuU5VcauSZ51TtxoVQf0ZRhhAD
N0nga+X+cRcbC5lrjXdDUYbZAQQhWgxuSSHuHaFotFPprH+0xz/o/b7QJl0GsZM3
dEqm4O+q6RKTWCyIpjFdOoieXYx17HykLgzod0go26p+iLz7AAR0YlH2sGogxSZh
9JNxhrAL7laBFFVgrs1D79AeJ4f8wt3NaUx3N/6DhuCD+36IbaRD6iMyudKizwgK
6vzjAqjXrvPpQLMcLHPQ1Y29t0Ad6g4NbzXR7O8O7BAwLoJdcOLJ5DQOv/cMaTjV
OOpRPPXne97BJGn68YyuS1tAVy//sDfG5O/B2MzuvcIzFT1HLITnVztdpPKIWwvH
LTJQcKSeu+gLJ+ydW9O2pLMwnTj0QzjOHB04hcg8U7I2OHB0ZLcPcwN72Axf8ZjA
pAHLkkm+EfgwJ4+LIu5SmKohFE0JMS/y9WklhV+RNqgQPap7i23Ka6iCBv8vvpeX
Bv4cwf3mY6nwQCE+iG14P9iCk7PzdyKI5v+q7cocJa0/T1wBWXqLxOohVr3ZVg4q
tFJ5AbeGKIOxbl0jjbIt42cEhIcybqDjSffzWg4eY4evVNS04O31Ye92pYxw4mTD
e/I1JsRastkSIbqAkm86P83unx0uZP4v6nnWbi4JXFY87Pji6CMn61vl9foeL9uk
jFAeznBpIFeTVIP5Qi9U9NtorihzTHsmulMQyNXoE/dEGZicF2wzpc+mroZHI6Tg
jN3Yc681H0igMPlsYkfkOh8mMGfDUzG9C9KAL1ZsbxVH4YAGax/TuwH56gE+XXPB
wpkGA+J2H3sSXdYI0IbsogRq7f34CPASb4F1JMe+r8+KwCxtZBjLjYiH3LBAREF9
v6RDI+lTgHGy06Oo64rUr7PJQDij9W2Fvby6GN1NRWU5QOIsGGl96pHd9OsCotDy
/WfcmsNjvog+WN8WLPitSqotaUUEIAgvM33jZSSN9rW8oYVYa4h+lyfFDaHu031W
tV77bjNH3K2m1L80q3GCQy/UltH/VDU0scR23W24ORb/t/ryEh3hxATL5bUt3HZr
+/Wqyz2so0za9pMBnrxBh17VasknpT+34RHLSE1n3YaOwxYMoAvkhi12l9WXWgji
XA+18lRfTaZerJVmMOW9mU0jROsdpGNOi4bh8XctJJwpNv1SlrsfOosV7y4I8Y8R
Rk/3zkkoOtFB/urzU/lD3PuG/JuXNejv7LEOAWXaPCdqXJd+d1lsk7va7hCEtwCT
yjlNNU7lvOzt5ClXGlTMDzo3X2lt8a6lXli8aWgpWqavXDTrw3aPJf3ZLh5i9AEQ
YWkdjHfXZRvGgTT/bizREXc0g0CCybYQmEtB2lYOrikiSyxZlXYWC+/6bvpV7vwZ
FzP3CYuatMYLI7/S6mqRiaOKcg/9xwGLYcfQjbzFDcdHpTAh0pBCRYliDlskcDcy
VXqvqIAGfuKaTJXSWzd0sbM4mxusLb8XzyMeNEu+9bqiYTiztzFOUJXeUgS4EgZX
ulpscMw4vo6nkF1CP7sbrd+NSHdGqFIkcQiYgpYQZBjzre6A7SbtPBXrIyCBKGhv
UYi3qy+AvuxrR/3FwTcXa+vi6jB7kYpgQL1gdGDsjlQA3P/yqARjC2qFHXkMWyy+
P1AnD5aVe/kpiT9Tm/wCUF+AKlHhc2RVyRzS5o4zZPQdKtIGiKiLZYxz63uXxzPQ
p2kFclSliaocCQnIz2GU6o7Q9zQnr2emekIp9FDKHfmkdtYIMto2yApiFquk17Y7
cHtKm7cB1Khlz+iP03DXFTKScqh8rMQN9k+BQdBVQXFlAGYaSehbWTLa0sMBXOml
k7Zh4P12U0f96iafrc4J/1DTGthIzKapWkNKLf3XM/lFyv3TVnlShnGVkWOYqm9t
4EbLeV+1YUlJ+LiBKOOBSi96C5u/VRX6BcdvJ5Xk2jH4lzqVXrdr+4/tkOmX1JPN
dMk6NZu97Mo+63CwJGJFgAbyEWtQVAmHgGeQyHODL6ImnmDGtXGAorcFrDTBQ3q4
8pf5wAPFiQ4TWWljI3Vvu2k7RANqauXdbB5k1rAt8x92QCeCOlwkTzCcjVwhPn2i
tuIt5bk8aJBXj+vhWiXsjTlFPo76+ROPVkF2bPCBtxQ225vdjnf278G7MbX5aMAb
R2c/5+Ptn5Q/JYVKwN79lfuQxYnzwnhQW4/jG/YUvcURmgsCVauuW2H9P5FkjmnP
nNbfIDSNFMEMwT7V5PwLwvey8dn1xJsja9jz1RXdvX0IAgXyU6ypzhynj292T7GK
yneEQw6zWLVJp5h0vocv+NIX9F3CvahEv9jJls/yiN9lxLcY8MA20LdicDL/J7A0
jKZMgA9vMpq3x9NOGHEttmTuPki9QHR37qpF32BXrGpqXfiikjNnKtuJDQvVZE9A
YjxZFffNyGP+iy1jXYwGRgO9E1POtnEkAbmtnmseJe4u/v9f7ImxPrl79mjkbYs4
CcIrBALJt49zuj97r+T+h4V7TnC/qM4ke8KEzdiXe8DTfsVUZhi7j6H6Agptw26q
fTnW6lrq5AHHawEid0ldWC9jI1mkE7eRSZCYBQjmMTkbbZY+Ti/7ZHBFXgRQohrG
eaOxv7NSipkeJFfHXoY1bUb6wc5M2GZCHoC3kJez8Ax9EWiCobjEomRKKDmhEXXO
BSN7SullFcNq4zhjs5BzWj427Uans1kNAjh+9p3scAk31jHBFmW90ptTwyOhpOPW
sFuy3zcOLhDJEmEkpLTHY3UGqn+3YACpJv/uLopV0pz9gfvCbfme3m00QlxDJkFA
RCBWFPVHxvzN7y2eG/HWwm2L6bW5BzlSXtshOP3A5B9siWwY8204SK5bKaQQwPo+
OnTOurGH2e70Vv6LGrxMN0WSWpJSuYbjpFaCU47ganlix3T+Swf5NdlUVsZ1zgYc
12VFCjMiO+3LKOAJAc5w4t/SvfpIOuexWPzct3Xhk0KlXnL/GNMr35eQ+YBMkRU8
6r0YlHD3kI0SKaHbS32bjzMWWvVwj3Ds0sDnTzpdGdNTgyQjyTPYKTLXWWkEdLA5
sNPUorpv3pdBmaG70bmmlqHHxYGdUiyV6OviI0qq6aZfb2+PcR0hmEJErVd8gPD/
F4UlpZ74cBHqe665ePb0342DvD8b7k4FD2SZCCiSYArf3KbGfuiDAbGe0pFEAEVQ
wVwLTXgYd/NN39a/Gpkoh9AeYBp2/60hsdWq4anWmhWaKY5YYjuCJtD76drEduz7
CdFWSeDWry10uIaGm+x46Qq2R7MuQO4vaT4epcDuuROPjySP6sWj4+95ajLTdLcx
GN3LrcVWAUj3DTXkbpqZE9PBGJLyQVBWVu8n66nr2L6fxhgp4TUUVu0mqLANsjns
sL7AaT6wIcdTgQ5+70e2qw05PZ0N7C0tYqtHQz4g/LqKk97paD6btpoizupfuUmS
leOqRgiWoGAeAbRfRJyoiJfZayg1hQSS3ZP9VPQwGNcVm6rzrL21/p9hJUuuRzNJ
CYKlRtJzmz9R2qDn24bTKlyjo136Xeq9KcTct0LcU/kpzvxI1kg4b+uDSrdYM466
hsQ3Qq3HSj23iRbO7bvCLBFLAdGM6leSWczj78yjWTwxaD1aUqcCwYekoTQOV9NT
69Ve18RzpguqQMh1KtmorEPE8Iq69ZKpsJGFnyx3ezP8oikKPC3Z7zTs3XSFI4+b
Nq5yo0zpLK99Yg2NduPaGoJao23JShveCncewqya+LwiUbJXlDRqSWD4MZLftN0q
lopFB8exw8UKd56MmyJIr5PBRLQqQPbxm5XABI0NMDmWPrd1tbBMPTqnBYTHsDQq
RKfFDMFyXlwmEgkPPKEiHCcPBTMugDssGNgehHR2eL+Dx9YtcQGSkGEg5xx0KMyY
A+InjvIcgsc3TzMNdd5FiCCSGBfBaDNndT1irBnFF81BBj9h6p84nKF3fBXwfb6c
imY4gnpPoFn8ooKFrVKLIXlFn9BobnzzLhxNdc7gmIb0NhvBuSrUgssYVXlDONd6
Vzih2Mw8upMHZHCSNKi/RQvYzPrQUgOvBEgi7vWkrcZwWxaTqb6zxnevCRES9Ua0
ySCOQoQkFQKV6c104Nrs/cZUzTG8B48V4uJsMkaditC4o70HN2hz/pyrKg44SLun
gG6d8O60hrTc3gAUNRD87dFczuZAw4WNpYmQVTHTX81IyXmw2HiFMtNVo5ImReG8
RaVEjWUCmOrIiLJIsz6x7b7Hrxktyjo/ibZdt7ycuoVgYRoWLUYbyVcYbscxVgrg
sJ2n2nkksCOFtvynrqBYClMxXooSPOwmnkI6pcK0QfNHBSFQy6kHepvKEvn2HY5o
iP2evlka70Oib+knJCF1TJBJhmomzXhV4ugH/1CKCc5pbghCNrBdb9k0HGtTHvTK
dePvJ4iSUn6NN3w1JgeG2VK3p2Cio612e+LWbUlZSWHGdeIpj9BlmQxU03CDgP72
2viyASDNO96SuWY2u2zeHLbqgFI+rXC6S5egRiWR26e0OCNyFnqS4ndDTBr8XS4M
svIy1uannLVWToA3+q6xJNfrEl/IKnmWIurFEIZJa9LIdZytt8kAiIdxBJXDU3lk
k9RWOOZ1wXInj9xJzaIedGA9N+IARNhw/2Ed9Hb+RZqpOgl77Urp66rPHzmhx5mH
cdjv+PCmqQO2bTUgHb5yFY5AFKeNgw8EYuJ4SEwhN+QdfDomTOzK4PZ63dnF82d1
Z8Z4pgf7rbe/vglRjcPBR6CHBaz2HnoT3HnuPQiu34jX8FSV0R0bchCuuQWgw7JI
Xm67U/JK2bXHyh1EQ6NcZiJSSw8BMkN0209f0wGzkvdbKA1GEZr69sc7taN5NMls
RsFAhziRl1B7ETDEaSWnuTeNwf9xSRfLk0A3YXnom+VzK2bgp8CqBQXwtoaXSb09
Ckr3IrJSYYMMBvF3x/byRxqmMW0qOisqnY28ZQUmdFuZqpuqhRTcuO9nXv9M7zeF
HgV5QiZwkztfcfqv1VqvA33OwhfqyFTe4gpuqImLTfET75oKn/nhs44rDqSrNZmn
bXGHThlU2CBy/0S1GgdXQdv3NYpWQ6ds26bdvwIPZc9g+AAQnmYdHpLa/OIfUfPp
Ct96XimmhXFSDi/jCrjzOYhLbx03goClvdKeQ852Yh036Jw4eMdXHe8vRZQV8/Bn
u0nyl+Ra3q9+RpLWhxCZY0CSbatX6fo26kv1UoL/Qn7wIzvofTLnhZf4z2/3dQJV
Ag7qOkWrUGsLw9s+d73MLnCFR6X+eilO0sj29HuxH98cOgvOVmA1uebw/1mTWq2h
eRrRh9OXzGR/KCmxL5XgoTfpfguFxESFHZN4Pzjc/cksm47Zqz+kdBbrNyXZFokO
adcxYG7l6vo/Nf5O41qrzdtGZmVWNkW2HxlxAd5f3eqd9os4CB628w19Ocvn+znv
t9+quIMK2hTNTUikJ6lIYIvzpQjV2thmKwtIN63C99Mv2Bj0HvN2HM9SdzZ02q+i
LSc/UHow6Ytf/9bld7k421FnemnG8QLnr8jT2oiNIqWhv+ZdTdcTKjOqAhZbBRep
HXJzUmdpg/BMDTQuXFmuCyl7UlFtfOdDegMv4CO2n06E903JEy/KeLhNqvwPhWad
jeSHmeuWdpMenao4lmULMoGR/sOD0XHGT3d1myR/g3d6PZ7I2cvqUVPFZXwxoPuV
FGxZCPyHYN+2PeBlXIzX9lqBM5hShnFokGtAp65qI28UyXeH+WXAzQTftBBCbn7/
lLcSgwFu8e7mqR8NNDCbU73Cw2QRLbv204q7hKhxvrVnUhFGy13kzIlxl4Jgj1Oj
H4GWKPSTNLam/UgugOmgfklN/vU8r9Rm8L3niSwOaiBrOoCFM9P7yI9TkNNVc8Ir
s7GveQFX1HTR5A5LMoATVulsE3RnqgNSK5bQu/9s074kOmlRoaRg25WaY1SEU5GO
DA8khc6psMAoA9ChUB6u6YoDlVcNOtqGJxpPP4xfZu5+whlCAT8yepL1WTYMnqAb
UftskbaUE1bg6/FRpPDWyF8DPed4Shp8hLsqF9eufdUqYt5Wo1gFC2nTLDritF1H
YU+d1g3ACNy0orRB+99ZUaqig2czxQl4E10oiU2c07df5DA3UzNhA++U/+33QUjW
1nupOilZ1jOtJGSQIqXyM2WKAGvGEiQp9lFRiUWU66ZOEImAIiWkW5bpR3t75t24
d2/do3WnV3y2FTRwwqMyuuHu1faV7DAvBsBMazv8vW8REFsNvfydpe8eUx55K56P
wHoC2YYoy+z/Et6YYN4Im0Gj4f5d2DYP3E/2UZTZMee89qa/RvDC0bzpsV3syJW4
6nUuINkyRyDJq0sUj703lkx2rUuX8APa9YeqAKcgaJynaP7M9xieyni+6tFA1+lP
XkJkuk+0Y3OVKHg7Rb1iXVDgPKNGFQVrPLA6pCMlMlcxTggWY7FcV6b4d6yggE+q
d0F731Qbm/ruP2JvYb6eFBq/RX5nwpa1f7PSchMWC7qafW1gdynavE4Ouq37wnxd
EB6PKPJf1Qiba6g4IIQ6EhJwdgh0UMeiVXBOdq8Z1erzbT/CACf+8yCixRBOn127
qfwhsR8SgUiumH9BZxvctxUChLBPcn/euhazHUQNGdLvOVJODLcLVYb5pSHGUNIc
uywg94Te8LYHeH6BmFaR3PNGaSRsQ8GpvgsK+cRrcWlyHjLst8CrwN38IhLekkAB
AnBUOfGJheyQl0UcmKnil4hJF+HnFNLHHJpCork26EGX+I3Zae62rdHTCpNr2m5p
8ouyjrZz147obWI/zTmcxtnx1yDL6/e7NK+DuVw39UOywCvtqi6aT4eCS3y8g9x9
ARb5Km0K8oEMlVs6wa3w8eVRRo0/b9+Ae3+MQ3eGs0ZCQIDh9ihLKzjCA/XuI7Li
rW/gTKuRDIQsofbHhuSryoNpKtHbnyYLn3t/JlN60eeOm5D1Zg9l0Sjb2fVOA6jE
4YDnfGgYVZ7/WBCwAYyhudqFriWZUOwO/95Y2UqBRHaFL9FHku01tzN8WGKd0r1d
sbmE5QUXK2DsibUjJBepw1hv6dPhsB7FfIJ6OGoDTTojkQQ+VBKjta8nA8zlX/aa
h6QhWUvS9RjrGxQ9o0KHZfEKmlDQ9MphOGubZmBHaXER7Ar4ZGixVM+q5Vq2DniU
Jze7ttJ+hcITM0v2KM6LNYZR1H5kKctfe2YWPeirdusPK5IW3iWiVIv/Q9s0CrMJ
7iqH5fuHFo0fXRaDudoPOBXi2ijboDPJeb8bnGs95PV+cibK4+YZK/6h4j9St+Qo
zIW5iAwQpyxYd7XfPZu54qP09935szZ/imz+HY9RkDzYrG4cH5QhEJEJ0T0YvD6+
k53ZE6ojdKBT5N23IAng5p3vLW8Xo3YntZRosR7by1efsOhRG5tkyu0IECpYX5h+
hkQLsCqnCfa8nHpOQcIHtZFxQs5cIX0CORrossxlhZHCp4pBOasCcIMVYmquJQcL
doJDBjPzNSjbQ1i38oWFM2Xs5qYNnEHsnV/fsr6VkeSUVzSllpnjZ7ZAph0MbdyU
QIhYLuPG2zY3E/3tSkI1cLwadcjPoagztJBaz0isZcurMukpKZcmPYkIZqZeBGom
vtYAj+AOKidDTnTk+9qg6ZG/RKShAaN3aZCMmR18UFuM5v+VK9On2v8sjPc0zAh0
aPgC0Bpw5AO8fOZ1mofuL12GqDDMiY/cAdhARoEWONo88dcVZinwOxIZBtzF4Ken
DYWSHxZgDZQ128hJdutZ/8TcHayfjXzxJzN367qqd4M7ciAQdvIYJj1rzp0gaVlM
0zhX1Bx1AK+D+9O+z0dlFNhCv+mGBY/V1JQbNfBsbdrQzyTI5WexZRFb066zdhPu
jtffEdAjrWZZE98nkMx8CasPt5AFGwUIsNg76VWRjrrqqoRcFGn7SVu0M0TnmchA
pdJkrd+AtjvfETgkS5VKgaNP96AX6bgLOgbZdp78zc1d/VDVnE01KH99ucqCwmeF
4r7YTRNUjD4FenPMuRwCU7mNEFr+4pHkhkdbcsGSHqiLpaf6wMWOPSpWWTlBjWm7
deaBvM6rYEd211YPZjSl7qgJQOFnVgLcooc2YnW+kTcB1o13KqDWsutRM+qhmyhC
H5A76Wgj/HeKY+n9/1NH7mrdDn59wWkzcLsG3dlPQt78z0YUUrVI81nwrzDrgzk9
L9UXUvMOtnvfN/qLayoHhMH5RoSne9QraHDXleQIOmNgrWyD7Z7oQuc1Q4FhEfpe
jfZ5BwrlHwBciR8nojTs3j1iZaVnkQEfHCAYD8oqzDVJJMx4hTVwp8h3ek+6GX4Q
S9RjvaieKSGku8/kWcKX7nygAqA7SSIaffWUGFpd1R1TqIg/9In7wkWIL+3bl4+m
yPxN8GpwKKgeWDYRQwmkrx78P/s8Aa2v1UH2d4Pyjg1Z6px1b211IGuE3lhvAt8f
M8ut/gKODjHIOh00kHr9JJA8lkaMX7tXtBZe3+SnTs4/3hIJVuiyWiIgundDGCiS
bKoLKFY/JaEudKMu+aktKgYhMp5XILngyh+rKSh5MslGjRcqBvhvd7IXgKhRKs+R
HLtbPFFqpdji4NE8nfioqV4E75vAQHE9C3ULwQ9H5r8w44C9qsDZZwUGk7CKfGit
sbdlbOJK+MjOI4V0N1JCiWjwqHwBBm+BtrzjrxGgC+49BpX27pHZr7uAPj7qYp5+
1U/J4xylCIKLRQyWaUpaaOoltNhRXw6htHYw/iU3PMtDSvwS2Cc4j/S/eF8FWPr2
/wMtYNrLSZ/fD1clhyi5pOef21chubMfIugGcsFMd8BPWw1NualinAKfbcgyqRTU
W/IpDYT3O+99CjM+YBxhotQuBJ4R8w06JpyB1dqtEl7ql1JGjX9Ij2rPSaLLsra3
DdgvTUNzSyKqgjCtO7vwSwDteA7D/8YQJfary/LnTHsMyXe1e+iAPngdFAR3imdP
PxfpxXfXu3ngRm8bAPzH5nkR/SuNB+2/HwzNkjFVYZvFQ9fnSj6lzxPkd/43tl3i
fqdnQtZU7ugWrQen9DbcyI9sjfq+4ytjMimBbRQH4lXWJVAH3A7IYfoCNeeOAgZ5
rxF0JkR3N1qd1E/iiGKTvl6oO/iXwJ5h18inHOVsBxKJN8pK8sdpCC4aVMGd8d4b
9HUqSQtjCJQBsDxbNMhj1Cvzp+l2nrQToyPkUSrcksOttY2KvwH2RPrxOB9shrc+
TQ2F0zd2iQU04hucf8lCp8F354FMEbzZChlVfjt+c9etchHdT6lwhoLcT6otvQtv
Sdp+8CYfzMrVL0z1r6rPNmsN7FU+XBUbnwxaysAnxBKAegSZmdZ5BqxALidu48yG
N37CpfzyAT9D8P099NjO/PZjASMAAFAjsJsQaX8doU8a5c/QSyP0OSA7WDcsCnq8
JNNYvirU0qm3Ke05b+5oVJGI4z54n3GOZa2G1otLDKYQG8qO0Uoc3zDpH5vFZeKN
2/WFLd9IVuKwjYmKaXBTnIEvjFLcGX/yvIdP12Kt2a8OkdauTz2I6cAVh2l8Hs2E
XD7TNhMlN/1YCrFdIaDm2fIcoI2r+C4VpKqYCA+lyMcmkG1IH7lQ0/1+PGpQoBYi
+T3P6eycH0dVUn8JDry7mNQdWTVnkJu1hdweBuZ6DXE7ObRCbHdap8YYLrWFHZ+4
TSnivb+kWzveyc0NZXRssuZl1K41inwYqUEnXDMYut4Ql5fHcLrNRcvmjfNJhkdS
iXzGpWWHxUUOh6bm3nfPo62Sufs4e9E+saA4knZBjufjGd+ICMpKAdkQ54G1sto7
yaoHO+X37NlEypdjwQJIo7TYUUSaWXl3jnN5SSdPv9gQfB+/CGMmBi3jPnp/y8Xa
Gyk1DkRnldLQ2wPlQ+PkmBa4NoUiwOFlRmo9SFkhUDmlqeMIir8rwL8W2HjlMAG3
Kq0gq60b2pehctAm65jZnRJ2uszNegQu5RHnJSD3Uo5jW52SBKdeTsxBbJEUJAe8
bzGM/DUQ09hf3fdGZx5y//zbs75pL0mvCtRD4OOYDX0281XpVK2QLr1zrmjnAhow
5H4+0DQHs+EQ0MinccbzptKDxhcrmvzG+TS+bLmEMnCCGeRFnhu+d6+gWdOyLGDE
gTCoO+qg9FDswaIY/aLvrK0dbehRRLlyrOjzTNWHemsQ4QGMtTKk/9iRqLskYJYN
pnLQZjPLsAGbhnKK6/Y9Bb5AnN/sTEku+AOJyuq40TmzFkMef0VEkAvf5c22NziP
G3fSGFJUSWGIe4nglEsGcUSiBZyDNM5MZG9jzNoKfMSmFyzmwM6bVVSmyCOLqgYd
b9WSkqURCC73UB3cx2v+XzGGi730v9wNfojIUlxZ+CNDqGuYNiAeex2dXkWJTuta
kkJ3NXY9y8WyXZbI1IaCTUqG88rObQFXn2b4FTF9/KDi0F4bpgC1mHKH5DV9n2a9
Zu/TA5mSfSRKfeMzFf+xNoFrOlnCyztfl1rkRbzsX5ZLB/VlbSeSq4AyXJFSpKYj
EtYb/ZUq+CShJtI2yiH0Ll9qfz20dlu1LFQqS+BvOIwrpGxmlb/thQ0oBhBamXYi
GxWZwJ1ddprleK+n8WEdZSQxkMPXDwUpp4WnOalloSeP+1k00T9y0JK2xdBS5Til
+3t1hdD3yt2VLrhiBncLxN6YSWnJw05lrD0g7V4lTXEYMSGMIUV6Fo0H/8HXgMqd
T1fwAGr4WBya7dDICEbLfnRvdbh8NAKWPONQT4bmmlUJyj9by+QlrqCPe1yK9cL6
n85FXW/Yk4YtD/9FKJEdORZNTZSMcz1pvRT++jx+z2Nc+30m43b0a16zG/dDFnlt
S8GpFvQk3V9LwylUlXgOpOQe+ZuzgF85GEGmV3WTfcmHdekj1IeeQNB3pVVOGPVS
qt9veq+9TFOspHxva7WoPvmuklcDRaqwrLysrDlucrEUDJkonZl1UM4xGK29XthQ
HfgLrttYcXMDvyE0LlwOpN2LKqRFY0jGWJPuwqV3V+jStAUK5uwK+19xuyVRk5HB
0r5/ZYwqu/MJWapfs4MRS1XdMjMf8Ibddr1CAApJilthPH9KyJFi8nIfki3JRjbB
tGXNE+pwKs9dO6zz0JVp2XZL3WI2YXQCWtHiHQXmQBFRSvOMYMD9hgoYwBT0Ubiv
/xHw6Fxc7pA3w6grI3GC9IIujofIYc4vYwc1g9pLQU4UaGmZAcjDTUYy+XKmMG2M
tvdH7tyDiJdG4lYmYuhj8H1Mtzl06Ig+6F+cfwY/l9OyCM0sQ11/Kbt2ImL071dJ
jXnHv3ap/fGcrCGUz/NVRfgbyhBEMlmNsvoUBTqhiRskh2UVe4tB7E7FYVQP4rVw
X+mf3S0vrFkgaOBZ6fqYUHCD/X6+rE91p2CePbykjZa6/mZzYKvkZ+tk3Nrq7SZe
YgL8dC+KFteu02v76QTvIsdvC0hKTaZGV/bzRQXWFI+PpZPugqYVxG4MzDzeIc1J
/+P503V0I6lS6+7v+RQ6hAXwsjcNOPRsqsFl3m/6yxdi2gV8knTUXnjQ8qUy1K/5
LVAc+xyp1rjcn2T1b1KwcNLg1sU7zDFfp1wVRehARnqZxne/SlVp5R0YomtMCdF1
FUrChbrN/owlI0UR0cKL2qmTJ9D1/Ath0CXsVyIqUxkm79Fklzj574qoMlgm1VIT
FM6BBh5a+opjgQ8sSCo2PGr7bJQ/ZW+jNESsEsiCJRRHTZs12gqZobFG78GepxK2
em2yQH/zAd0EpSofDmDz/9LRb8CbDSjq6teo4CEKPPkCgMnJJrda1o3uB25A8Fxu
XKhogi/5aCl5n7qObTZ/M/2uCgQX+I8HZtHPF+aAb3G6iAoAtUpomBlY6oKOSFvV
lqCYd/mepY16gau65sxjYkjf8NdA++mlbGVSMa0ooH5KJcx7SqOiVWppLjJU+T3b
3eP4SDKpy5Imdj5TeJGSLk/TOArauZpjzSOtOJHfoGJ6F7h12P8J9CgQdhplnEd2
v+IwdEuWMWk7U1AjG1h/hgYvY4x2+eTS9bKttSmWDPIL35ntbBqGC0MHUpX0btvm
C7oyt0Gm7UWmMBHIk4IEUKVwrnIOz2gIU/tUrp/BafthOhDj/0+0bsqMSIlFrB45
iux+QH43r+rTfPv72vh1bFhEmEyaFzsDqC3f2lpAdkhL8now467kUC38bIEmCxIx
ZeAjmM3kVPYJj9PkQdI8OXBPdZmman58JqtkR1kHCHELsj5LE34kcFBbPR4uX6VS
SHBYmmXMOkK51tTD+Py1+hO0ZNvc8N06+6AgADVPeIZMQQ0UcJY1LEFtbr97pG7O
XUlGNm/dMgdycf9NoKd8srvHNf+l+sO+FVApehA1WpTwz6008I+WQVrGZPgZeU89
llaemY8GQNPJhc1gXGpob6B/obZKiR2VZ1lXeos8SueONu38oJvg1ieE0yVAt+DP
U7ftl5Ss6mT8dg6lUfp9oWYUG5hqU6bChbMKVyZWt8TvUoZW1FM13zZCLilv3w0/
eQI/w+HQGU1dIXfVUdCA+LVezac4xYOU9fi67C3+HO9dnlK2fUgATfm9o6HnfL/8
PVQwTdg7n1XjSGYs766jx0S/KJyp3Ne1HFAgmUsAWwqTNKiH8IUKZJ+C8WV/Wkqo
nwuLPJ9+OCz9+/SkxfrIktdxaS24p/hmItYtrAcwJ3bemHpI1crQKkaM5fv8GDI9
nlkoP9bg8gs1YVK9Y2LXlA5JxywCn/NzacLBzOtEaBFndSIXshLQnl4FujQwl54k
MFt1ZQLe6vXFuEEyiEL3xe8F1vIrT0HRlbvSZKa8QYx1H7/Jhs/nc1r4jtZ00o4s
Nu2qX7N0jRWanb3puA8shhFAbT4k5cfQBfWJkEL0NXjr7nwQqvFXCCthd4oCTFeq
EiF+A/e3lM3Om4k+DPVOvDtqY282rTcCODaGxfdKBY99I23dzdEgxBwzFT1uQ1US
m2NMJZrh3fp63VIQADxJDkjX8ePzy7KfWPpLNUFtrQ3LNcEmjrgFC5FrHOvLNyNm
OVZ1QCCjZEQe2nAh6EC52X+JmhVv1DlEqybpKABvGAV8FiloOXVgeCaM8d/9RR8G
rHUkEG3ETkRKWhnOVJTML/hDrSGfL3Z8BliuFU6bKTjzyo6me5CSU8HpqHAJenBO
j5hz4IZ9uoarefqRUGqPyOS+AKu0PlyvvjglLG3Dcagw3KrEV5pIzzdHpY6N+eXT
NgKyrd5/VAN30gSNoHEjFOwplj3JaZq7G+bX2EuW9qcXnUf1d7vNcToYhDXGSxSR
jznRt23SMi3YX6T0Zk2xsDw5LGNgeD/1OgRdG8QVziQB9piKyA/0ljBHzD4X3NJc
lv7n8O62um7SGJtL+W8wp8VpNiu+Ixqw/gVu0bWTZk3tSU9WcLaEcW+qz1QqgXtQ
k0pbyo9w1HFP1wqMEKwLmhcHgYnn8tVKLBz10HocPVBBp//QvMaMOZN0DxB4m0B+
YBKV9Z3fptyyjma8B1P7nN0pa0SUFLp7uSSCw7I17fNBWMGnL5wcv9zPu0SSXnel
TAiqn5pFdXEEhi+ptkNUqcro24wP02GEkBpWfB0AtNqLpP+N26TQl++3D+9Rhf1Y
1B38Qz1ttALdS6Vzcpr9yslcGIBjuUOKVRJinPI+YUDvChXbCB/9F1v+WZ/UiNzt
nE/ahmmyicsM63QKtI/snHdzJV9J5b8vv4ZVUk5iO8hxrwZU+QNQ995EkSStYqcJ
DyFM2qlMCgCqRs7+DkeDP/sUFo4UY9wY4QDtp6CTRiMBHydlKJFBPzJWPUGtYt3g
XTz8e6XG27sVjucAIYrHhmn+TtSSTy1AOjiZFYd4CeC2A2MC0SVXDrkUqRkynhM/
pPUmJljp+Tx09q2PrXIm6mGf1eeDiLHI4ivJtF998YU4/evuAHxDhljKhVa7Iw3P
ytBPvoCh+7UheNggSKHIJ7a3SRRCsQ6OdDAzylj1YtaizJaqNLCFQXgMmICyDP54
GlMMW9cVm1dpOM/N3kUih1E+VwL7yoTfTEsnuxycillZvbcGDt7sdFHxs+HuLI2p
i8ELbi89pgGs8KJlSjEOq6ijMHPXPpVLP+1+nq6Qg1N2rf1/YSOFgf28iHHLDHuo
edSG4BMZnIWOC/tw2LmolI7vzdSBTyO7/oP8TBfztRi2DYHzcR2fEnayzxsbH547
lKfKOZnhAMRqlXJRowfetOrQGdzE+ZxrycTeeUD1fToPOiYrwUceuCGkx0d4Bepm
41NaGeYp3feih1/ReRFK2naHlgF9gsAGPx6S5dobj2qsMjkU+6KZmC4EZB/8Es1j
2RG255rdNpOy7CypLDrIpZO5PBcayuhWSEwygioUCYla1EjFE4pbhZE97iZFf/Ix
CUVLJCuO1j+adYdPtUK4fMTipU2Rsq/NqBdACms4h0YHG4r2BOtnXZPSKU1lRJYH
1JRzPBrnHu+7psA66FTG66WH19cO/jJe8O2wUhzMJIVthRAfw9uhSyUs/eeekMPP
j2dBLEFdSJpN7Zi51UWmt8KWdlD6SdkUBZjpxpahnbknFo6dwnFJmSN3sVYBITjc
UjsWHMQ2wp/gtRMdDGD66hnDqJWsQwFpmHfFd/00WWHvl7Whq27SVfXXTSi2H4u+
IFczJ5TVlnk+Sg+g/5T7yQ+9+tWU11EFlOAo084J1ijIm1AhHT375TnFc1u+TRQP
raBrLU5fKeJSl9gChyoBDKioj2bq9+vdPbUwr7WDAggrzSE8mhSt0mE8Di3uzSh7
Zu9vVVb7PmGd5pz+AIMJpm5Pw0V5b8E5wPyyLRfa37HmtWbkLRdnBkJK6V8+MZWm
V6/t1tFewPgWMHmhzDSaNvHzE7CkGlit7jj84rgQZ3wL9l94VAo7P2koPvmsfLAK
hYlgQWaAncu3m4XsdXQGXDBHA/RwNVieh2iiEIMJVntFJJU3N6Arva9NgVHNevac
jhDav0vuykXAC536hxe/EdALTyWGQFt+OrblmBomO4/xyhaWtL7lHgeRY6yJXchM
pJ3GijstYYiNMw391sIKXpYw/wy41VvKDB1zbVTnD/2fSpPc5hR1/mhcdq8smEBy
0TxXG3ueOB6hNfnVrM6U3Xe0+g+7WG8saTu2BQBpnvc9kEt0QE4ADwFMygnOgULQ
OJny8c8GFlZN2ThaZJmiaQftssg3km0RimHm9ciuwnV9EqkAByN0LAtdQiLZ5aXL
oM0v6YW0Gd0Fx6vgjiO/Vcce3VY8hbS4VMfaOtCq3KgLKo0Ui93IndKYFD6sdndK
w55Gv14lalAQnrBmfqqActVEpgvgs0hy5HWqhMW6QcI2f4nRxIyAhjpfZEzdWTYX
MAJYtMdydOUzxtX6JXbyRxx5exMwriEmllY/xQcdId1W9a9AB4nm59ZMluRe0RdA
3vjh0To6ZscdCnMAgBgx8zMl5To8hnvK07SpcMZ0Td4MLxmmG6geA9Pethl50ey8
6NVb46YWNToEE/nvTipjSPF7qocGrZjKh/SOgoirkTZpCv32cVqzAP8SgXABzhy7
WbYO5RGh7mL5oqDdVpKpYKBueYBH9rozzA6pQpuwMZnyKg0ECD947zAuISUv3XkF
9R/EqkQo6zv/2HBpji6C9cxF91ztnNNmRrzZq4K8j4mdExIbP3poX5cpaMWqYptS
D4+6L07Ofw7W98v5FCKFi2FrmPY0Ir5ugP4OFQK/bofQD8Jy2moThgPXbN4KSu7c
qmnd425Yl6bKHqS3pKqFbfEENtbIFJIjABVF0wcOv8IyUs4ti4VTSXjsNmvONe8A
HqdnTYsi72JZhEXMmFimtOcbaOEjPF4zb2/sejMTxcstB3omYHRYPS+0RgG69L+6
mQr8u+wcJZHjwF8an7NJGlmYp+RiVqAkzporxu2iiM1o9dxgy2b7pMtVMgPzJDm3
Ev4a3aU54CMWKGUXV1wmkuAqE1uKqM2Al1Ryeg9G4Y5Wcf3mVx5iT/4jhiOo36Lu
To6u73wYgtMHJfUlqc2YdC7oJ8yIKHr2ch1H7AK+ASwRDdt73ly5fWaR+N3e4kDB
5RKUxAZZWY/61jNcn1Jbom4QRFuQtlvo5M/6bCRcB8xlanMoHrurYzSIWNo8Jf3x
KchOx/ou7e9RU46jppn2lKH5l2TW1wjl7YGZilpoOyeycUsJ9FTuHAbwfZE/uF0Y
DoG+xDnMJ6EyxoasIpVz+DOlNiBejs6OGqjwrQCw8TW0Jb+5lkYiH0A08jvOw5Np
DS9x1Lbat9J2FJT015GyfsLZHteAg6cN9zPVhfUMGuYEqibqSan7wq5j+wkw1fpk
9v2Cu+al94JPjcS3TmBVbCmram9GeNka+sFb66uZ53LoTi3SSS/p4BtDnMIiOAyo
fWqnsQ7RUkhfRU36ydLNiCRoXFxA4DXYlEs/yoLyQ2m3PyKWZKKONkbM3+n8RgPB
ldWv1bBrIah91EoI/r9O62AtqbJXycQjq9RIyAN7GoxPSt95+okLnfjOC8Ct3a46
blUL+lJOKbwf2aMkgJ4NUl8KhftIinzdlvyBQX7is24qMLjgQcttgbYKUmea4U1K
GtfwATjZ+MtZ5eA6UHDwUlFQor3QiOhF5BaaD3UG9WRpZqr5hGcb547HSUDsFuUL
cl5DoBoS7CyjHzm5c/0GLskartwxUEEonIENTsv3PiDngv7bUD2Vqc8BBToWoeR0
ExdCSn0Zj0yF8OHwJI4vIf3nnBZAJ/vm4UYLXf3zM2ZtdapHwYaltSm5wNAiIEmG
kXBY+7I7Q0svbAHSrKo0yhecHkvXz5IEle0fKToSCcORxLBFWIA1B/MWMdYXymLr
jOo4Ag6Mj2QN0p+gqZ5RibY6FcEVV4r4k1QloHSWbl38U6+w9FmUb2r54SRxvVP/
jcaL2nwAxH7QRD5IsVKO9bLGjVY8KduMQe4P+YL4YvGXTIRyxTm7NejSqdKa5KgZ
oaCmkFK+/0eAFJlrPLl8mBahuTcDoxH5b4McvUkBqQUSu+kGCUTwUI1cuZcHtuLb
9zTDQfcWxKJgl/rDIgFihgXSSmoDxeiQGTn9ricP1Ka5wjn3yaNYHZYO/qb2AAdF
KHMK0NtK39qKShDJ20io2O/no8/NIDqmPv9eZ2fWCzd+x/ZQa4L30P2Ep+hkXIuv
tzK4O6bIBPvRq+NyW3YBlVgdUggyIYeeXPfhqf1dbQk8siIpa/WTyfzZS6Iy1vSq
as/IBVmFWvf1N+R2nOtx0o+uBoq+DVgQjHqz1as8BGk/59Ni9sTHZsHxNIAmokgA
mp0ZpCHcniWi6CX6BGhCS0Q4+tQQTZFQa/67180olQrHFtZ178LRnnzrqZ1dL8rX
ySDvBNGj4uscAwknA0gDvEN7cPIb7r2dtBtVRjN6JgoVlblzRIJInbLmGOKaq9JX
20KvTiC/AiEKVLeSzk8ZoMaPfGbWox+NEfPqzp+O2Em84jGza8DEaIQUNo9s6k1z
v0DlXrjLIj513iW2ny0veh93OMs5sqoThTHtwMH4FREdyljDvkYGpPlsdwAO5Wgp
55AKTMVmqQCoS4uh695+v4SwQRlTQnScZFmh/KEYn46CJW35DEFAgJjP1TcaVnBm
iRhz9DoIckoDHavVU7q8RMHjJumgpJbNvOi51hfNcsSdyZclIE+W6A6HCHahn+Sm
PMjp/tDKbO9YX6CcGvnYZ+wQSx6lN9LcyZ8z+VPliWvHhU2Z8z1VfWAhZBMnmha0
jQfy1r11HEPvDvekD4V25CX+bWQ18zDEzFjxNqpgh52hFrKQ24WQVai2Wiz4CgX4
wtWBUM4lTi+yS4H4M8JUgYdgXZKIQNGHgU4VDxlD5s6Vn8rwPcwwPFFevBxkSzH2
sa4Gh1CppxYGPyZ9iFcHh9J2d+Xq0o5GCQBpTM6d3rA1DPXxbDf+Y5hyEnJN9b/K
ucKArKp1Z32TFsAs/IHsChdUutITf1YrwMaLWckz+i4x9MfKvcFKjnrhi5+vul0k
zrsjCJyXmi0Ni+YakvoX2SxpuWCwxjnBkBdSL6HDzD2zkHQXk8wZlpThQpMqFr4+
kr6kQy2cBaa8rpptv0vti/MJg6s4OGCG74IP8CNp9+zIsw0G80h4nOyIKmHFBP7o
1W6+ByW4sxjkwo8l77nII8DHI2ExQT76eMQ+0VJows9W0nT8aCsVSc2EXCXfvxuv
xNqyZ79CWUx7opOyvBhyi93+jY0DctUIKC1ot7jkXOV7r9HuAeHLqo+qX50uFYqe
9QRIjPL11l6NDvneqBcYz5etlOzNt4VluWpbkkUTOKO51OM/xzvidCzQIjGdvZUs
5QCUrjQ0OzSLv3I0njmiS18omarDzuVmE/U9V5C04Yd9kI2MPJsQCemOmMy/oBLs
JTBwCf3rUfv7OlXDN9OcC7siSsc3DGPoYSQxYOHic6dRfppZ8gwwN7D5JbS1od9u
MCRv/z0uEBHV4iIFIkxx53asXbU7E7B9itEH7Vfo6FrCvIuV8rj2MalzpiejUgmZ
OuB+34psPAGQKW4IYP9fB4mhCHqLhRywV8GGnDYlfB/1Fv4lOD3BWAz7+3gC3R0N
Z8DTqb+wzyvrZi1uteQwqgrju2t7NRZQyaYWn/lxKpQ4a2v/U2UeLY2Mi3iMZhis
LZY6UY1t/UpTGcV0ktE5s0LNwubrs2a564YWmHSrumcODmge7IudemeB7E4mgIgO
LsAVMRlWtEzUyMIuZ8V/wq0UHhfOrkLvHqNuEnivFXQfZJfBxxzIu+X9PYmG4ZeN
8Eyrv8jep7IuNygBarnSS3lrVaSNvyriH2dgXOVIU+dXotAxpKytEmgTw9orgwk9
eq79kSJuEY9YvFuyAshN0tiFDu4qHab6ebcOC1jlYSWKv8aLz9HBpAHdbEQNZMOk
oKs2rSNm/LDBtnWMaUMsaTRVnNUPRoSgHITIeLBlP5wQc5iofAyVHVgC+yjWZqyx
dK4T+GbA3ZDQF085Sv7jZNXq57mHs/BnD0642wLeUDPBenrj+zORufMBG22ojbq7
uf3lIWq7sX1958kRNOsFbEACldV73aYlBtztzubzsFvx+MmeL8OqudOAruQzcBfZ
VFJnDhd2Y8UCsCBnYPFmV5n8VfmvyCnje/lMRoaCJGjchUPu9Tz4fyYRboQn4xDa
VLPSR3GZMO/l5yfjcJf/7ptcir5H0lru0FnFPCXu2MlR0ISjOrJDJyuvSGQ29CId
MU+wyAXKTRLK/G1gfGyQ+xh6XSbW7dwEUqlgcplyGrzcrxQVOnw5u1FvZYoqBIu1
b6+/Yjg8tb1Q4xQ2nPA4YNNfkcblviccrr/ykouaiOeNUVQptF+pXZeKAKsHbasi
1+oq7gCQk476jRAbUNrzA3pnZPwlVnKzL2FtsqLLDPo+N44XlTTtvSjaQthCfJx2
o9d5GNw2ATbYQAyFyvzaCe0vsnRvAF51eI949EFYt8J9fxLCCM6BjG4B1nRdGOws
9eWBsV7fHgNtX6Z/iRp/a5LgZt23Qe20cRuZ8spwZP2SeZpQ0uxbBb0SdwdMd1eH
ucvhT8J6O1MJ0vLd30BUuOTQBBe65ZQ0B7T3UYAOXqyBxfK++XiZPR2EHc/Xd/i4
HtpIfXTT5n8qj/RFewt50jIwz18kiJm6LVrcoujKZMTB1lNqQAXXArQm8j79stS/
6vvCj1BGb91UcMuuWoBLGSdnIY+yKtR6UJEPkIfiCFcGi/8tjBu49BRVMcOYJJCf
ukRwSSw5sZnET2x/9z1bbU+JSomBtqHiucLmpXtE3qkrfHTW/vTaqqwsNM8AwzsG
j9W9g2QYrivyoLBcOH7gXdL1NXkOo5anvFcxhqhNsQ6QEQvgX7wjcGtPvSMAmMKU
EDUbRf8OQbDmKMnfE4TqsgIHZ+wLhfQqWX6tVyE4SfeJJWagLe07uFJBasGA8eB9
yEFQa7CZ9hAbiXn99xpn7+tYpKMmevDOEsHQc/fif9o9lD4tATohIe9BkIG15tBV
ea2YGJG4BnrYmd5s0nUrLrzxscAVmwGtSWZJXdhwIINw2GT8fY6S6P2IGdF9lXLN
HQKUdMOxqKhJypeizNsF4er7gVPGtyIfnlASOaaSVEX6N9BYPulzu9vq/4jtkZcA
xtItwRb6pxyZFKGD0+qnTtCasSh/gN7apNRO2S+AgQ1pA+jF4HKeXwLwNP93+8vC
Vg0aPfSXv2rrf9yRScLmFrzdiaRZwK6CD2gQnW8TufCNGMqdakq2Q2Ybw0SCoZlo
xWo2kRGCtVO3ne9K7iVUEvtGhDm4PPUx9p2YPTy4D5fVSCQWSO5+L2wxklS3uhCz
fVyu7/JgTyEbuLveqYVgy5v5DFNKe5w1IZ2/Q69tX/zSAI6f9KaERwFkX8iY/67n
v0tar2LQbodBbzWAJ8iE0Mp9WNBBMKtWsQAhA4kiLcP6H3WSlnStlaxHIVXUx68E
rUNeQRV2eJpn0DXbWz8ihW5yqKAzhoW54e7qAQDlxqp7emtQxm6NSzZDr04uKqL7
6BmADDnDoS4R2wxzRSgxD/XeIKx0CIlqh5u55QY/PtbQslwQNkg2rkkNSJCwfpp7
ay+yGcznbiIfZgsz7r1xVtbWA3iC04hULwOyAtS5HyAckEMOy8ioxGjzXWiCckNs
wJp1VsLhXScXkxOG51HhCuwlHD7CRXkQDAgFpZkFRWZ3NbZSjvdxQdQ/WC58cnjG
2yoY0V5j+xa+Gi5dSJzzzf5bZB2vu9h+jXcdlBmqClETsYXYEnnq/iDSUAgIKUfR
oJOCvpvqEfm2xxognCoAA8PRPx3fcE9o079+M4/nXs813QkDjXWeZIt66H2T5tIq
qioHr0GS6R2T/NN+8dSj44Wijs0Xhzo3Zce2VqruZVfMljaLv8vfOFxcsU6lR08z
5HjWgTNYgSzq3xJRa+ZBJCpHw6OhURhldF9NxK8TST43M4YF2RlpeMdNhsQkoiBb
EzS3wNFm/aShfBmoonQB2J1BiZUsEiVC+LMW8raoa14iAWULHyBcet0+6wsF1nAz
bxYtKbH0oJfsWi2ifSse6M6f21nEem2TPxD7EE1YAN9vmGlx6b+ynF85XqKvoAr6
ZVKKfPmzeflS3rlsOOyM8P5ErLtoeGp5emQP4SDC1/JnAkDnXG3C+be7obXOsoSn
ocPsfRySRvOBATkY4u9zSC95iZWaazwxz+lj+aQH7YiUVSAqc6He+4+GlOHgrLIo
sF8b+TDcpmoALe50fljzRDvpRWFkhNdXTlhKUEsVAxf7qmI7QIGy9fkmQ1giYlaL
Dl7VjqG4KcxB5GVcXsy1BbUuLgAPWAwJUDwgi9fkYR0N3xhYgWYf9q9PB0DA6Mjo
dB8nLDwaO+KzlCnb+tb3N/srlCQJTwg8AJN6lmCFW24rKUNEwwMm0at/SP1KjQys
lgWpoqTrMnqVn2OKp2gdzshKLH6fMNAmSGU2PgjsjansAae/mVthG0Iera7ugXFx
bbU1kLw2YSE0MArJWgUO2BgQc3Hakqb8gpV7XDh0HqPlMy6LEewhKHSHBOFeIgyt
yy5FVcqtxrBWxT67yw8BEOefXFn9YZ8lt745KfdpXVMhDhqrLBG/S+q8JbcjCgtu
zzvIkFpnboy+raRoM9Gf39yJ8BhUvzQoecSGQ78zkfsjKeBtNfcAyY65dGsnndKZ
1URxMjW9YNcKBRb4eBAE0HKHr8rSRY3FrOa/GASNsVwLDt5TrA5cpwhyedkA1zYW
7VhlP8eF7MYCkA8SOGnY4kUr6Chwmj8B9a/shHJU7ONuXBghGVg8XfC24LrfU9EJ
/nByjE8iN/nRI2e9WzDXTg9Z61dT6MofPLvuS0S/Z8QDQAI8gE8qP5a2UxlJ0QKl
HYhdmD15pcNiIN6uF/+BXdjmMELrtKvwuARDBaAo3qT/7PmQb5v0ykratpomMJnB
02uD9tzWGd1vJ00lx9v43FbgYpAodjbfxBb/BNuY/NGiTSVjxGPcdIRXeQYGBpxi
FOJoOGO187RLfvhkiGk6KIrFgaHYW9fWNYB71n+sgfpSVAlSe41TfMr9pKK/wPHE
Gnq+niNZf5Rxj4UqSLDx1bNbEHSd8P4FWoHHriA+XKGNCsF1wgiG+NIZbSK+LHsF
1nLlZlWgFDE2x+PfwLszltJCf1PYzGmMtMA3ioZFFPCYmoMewROrZGbGARJct0wL
kp5KHnf+FxZsGMLWRLs3GgJHXV0y4fD0OqjWEEXt4K2a9b0fJ/Q+KzOzP85ZjBCF
7gY79hcKDrwCpDqaVwElVyrtC36OJyKiW2nscQ+h4o0680qNN2LBJ3en0pnCev71
hjS9dMNFh/XA/NL6u5eBlZXYrPwkqsgM6MVuskoHGCapon2Uw8IeZPrLuDijqHew
PfH92EwQf8yRw1OqNK4pmgeTe0TrH2rhN7HnKtyHKJgng/W9wj/wJE907KMEcWMf
ZALoE6ZMRlM6KBfMGwrVJUZEqrQN1lTiXn45iQF44bEmA8foQF9XjR5qcGpmR5Io
sI3EsWXMHgQjobeDpwkq5DFEbNBhpD1ar5x5mcYZ0JjulOXtA3jif2L0PWJ4dak7
+p69t5MSI4CRj9Mxpl5TwHDOBYnCXcJYMuDN+jzj+l6Fa+fbm31qGC5iltTLbvvB
bIa/EjS5IaKrr5YLv24/9Y37hhciYyc1v1inXqyTUIQ643fcFipy0Mo3dczO+EZ1
qFgmrvJffNeQJRDK6yrzltilWs4wDmOE0T4rMH3iNEWqLUgjolfzGhXvZRwKIPhW
Ak2agv2DlnbPupb1UlzNpj/vYPvXwmzLUAAHDRnSFSaaZfz2bnoyYWGBVv9wcR38
ujHx2KxvncaQjorYWHzFoCVwjLqRN6D8FNIgfxmLrwwcLbpwJu9yz6s6ejWP5K78
FtLpQe45SzBo6bhKsMOE1UtCZa2CzYXESOpDzwmm6Q9xDqnh5/swW1A1ZEBxJMaj
YUNpHu58OgSzJ0FYPcHyZJ+MIxGyW4h9L7Xip14q+1U03YQ1dqJqqk6xyBlVEJIX
UossvVSb9Zk35+gxYsixUGW2MrxX3QMwn+6AE7NsMHJ0q9uGz3JYh+qe+KhtAfYQ
dXIzb0f0Z+jYT/VI2SEcg+eYp0CGE1MGSoj0ORH9+7V14KXiTlsHNUOETxdS0Ad9
boWlBpC7vMU/ZLk97OHc41TJV6tfO8SXErKCrDTVVEXtCJKLCe5hVjsgdsubMD6I
C5+AgJutb++H8U4ukS1QIYYJp6c0X9q/aRwHPdvli6pMusSNh/b/BpM3qAM41Ib3
6xRhaS6F1qGlR4SU5ZmTssppdxnrEPmFfMLgNeNRhaKkOppic2zm0o0R8N2pgipQ
cxAxXWXbTX78cNcTAQOmDSIdOwL/Y/D6fbnZjGHxBWzsrginOgI1yausBS8eZ2mV
ildkD3ZNf8lLY+BQ/rGgMlcNcc8FzhguA91mYWqiq9CIcsIZTWoHA7dmHxuMCbL7
P/AzCzS6zYU9ctneDZbBdzPKccbHEuGkKTDx204Clmu2b/vwHeI74YC3DneEABYY
e2ykE9VyJ8y/D8OohHwV2mG/kNbRxmhYJZxw6DlWsjObMk1y4ZvxK5gxMH0y2q7K
9cQDsufJoP827fsAIog5F8snfPyr3mj2RFky4AOfU5Lf3bzZ6nYtM3ED0nB0RVly
AlLOzcWggW//FyhD0aSv+Mt7ByAoM46ueekYq7s1QuYV47Sh2zMZ+h+l4dWxLtDv
/G+oZeZRquUkJztkSq580R7vIJNHppqobtxR8gZgy2z9v8wPRL9W36Lpro0R8O72
hkBrt3wtVpf6asynsR5a1yyoBiAEZaBhsrtLTP+6uOXL33RiHtHsU0lyULr9wdsT
GR7nNrIDysy2rhW0udlLEzIsdreFkhXYbpq4s1ymJE3Sk3GSp4riMevkxLTsNsXd
CwV7Aw4ZDiFGyJc+Ld+W//iM+IKRcpoAt3ppbkUsc4jjDDXo56wJMLmgenvcsd3I
hVjwXsIbxHQ3Jd7g4CSlnUOEpKU6hweGZjnkhw9A1g/9wiGPjFW7snZVSXD6YhTm
0ablSrem/3eg5yFIQfHvCjCBMzyF59+8b7U+PjyR9Rxy4RvRE+ZdxPeYoZzySP0j
yMDywM+qK56LJEsK1SvDPpTfUafHuNkpp/dSaMFJ+fjJcsrZRBt1lkM7BdWbb5Xp
DlQQ6cvcL86rCM7vMuUAKnCcpEWpAhPlENHwc4rPCTAru2P9/akL36sXwEFiMJWA
XQK2a/Tu5atloLBsWwZdfNiX9SNatEjhnPP1A+k7jmHLxjvMNzyb0RTO6p3Uf3XM
ME0URLMSyJ8tCNrbu5tjNv4qAnqFkLY6JrSMyO3zLkBUTa8E+5pw/3yFzAaUn8wX
YNOc5v8bz/3txeX/OcSRMFqSEaIKxuFdfpK1U4arUp3e2w70WIlEU6MS4Qx/WWKm
oK2X+a2i1HO4c5T25AY5VVvy++1m/7ndtljYscA1ORMcuZdmYZs/ZQYKyEPuQBzx
3Mi4jt+zPkCGlKM9NTPjvpfHeHtlJQ9dJswF9nyVqAbtxaLNzb+8001nGRAxpNQU
WrxmMVd1uYQuTElIwOhwsj/tDcF9gNGcDu2vtOa7oNS2e6JKgp38viMPAyXRE+SS
fFNYa0gcaW7aRcDpzVrlAw3P0VUVA7hq8rFqvzrOcVsddbKTpXswYyISqh4qo72S
e2/fTtN1Q7L1VE5VGBiYoo7kTUxr+8JR1tRvfVIfewxWTszsD+ZsSD5i+nK8Pc2a
5jfmsG4hESYgRGhLGWGDYv0ffoQk2dYwB3ajGt/KHwamYvsug9D8RnYz3vXLhCue
phX7l6KNIWXZ0Cgft6fbwb3xBhhHTBqt+GMY+hQQqCLajyolfoJEcgSmKIkML12K
8iUGsnsc3zmeaLhpfDpW2hC+mNpIGU6kZbrs0Vbij5u+Bj9wjusRKJczHbbqw/K+
xlLUWub69ibfxPucZnY21PE2xSBTCHmIgu6GaJTLPzHnvC0FqnOj/1G2iehzb6mA
+2bVcSeal5kpLZWuvr15Ld/dH5BTZqFtkOPiqxciblZUW0vn5KK9O7YvOOuqoNcg
Sys5k3bOcgxIjBvCUCfM5JMk9/nsu+WYfpWtVEHuoNGwQjWn4eP81XBZ8PFGt6ZT
1NKRGmUdwIfdPK0SCkdiEtw3MFodzQnIlaTSM/Wq2Fwvh+5awXlRMQZx1yE/Mzf9
yG689wT3Fefq0ctIuVyoleS8dysUtuKvrQI0kEPkoDCzNr6egIbRVxETgTJFq00L
T1C6Fq/aCUrHKRfb87y97VrljZf908CAVIdE7kz9u8XvOK6SM9iEkKLH3X4JPk5l
sN/yJ5wwA8qqcjDv/EO0gV/0JqS1jfq7kUo05sAWZd08o5N3l2ndt3sA4V67m4Gd
Rx0iJkBxvD0cf7Y8bk4YRUY9xUAydU4t5cNN7jpxivV0P3f2HjgEGXXmF6//mk2W
vW/xorWSi9qL46gR4fc1+o1Jo3gpZqQWxLUdwVu4MCW9g7IzavfqsBP24mygihPk
T1h1soMlV//V7GgaeY0mhz5IYu7K/eR0xxTnsbi7s1RqjnTgkcgdnMCruHN+6j/H
oLNBWKz8F0+64ZLpvWX28fPsPGAlYpeWW3asZd139D6m5kKJgOCplo19Yo0Ob7CZ
hAHRADl+cNAM3TuCXpVPePEpDBh6JCkMh5MzG0yHGLouQeckuXSx6u+mmTZI0+Wr
vOxQv5gx4LqZoIQXNKQNJVxHXG6YYi9B3W2Le8cpsom0BlzCSyWF05/K8RMq3fBY
gbc7U9ykE8Nvfr58GWWZub3C+j49ONejCVUELokYNmSmT8wjaFcydbcsyd3LXxx5
Ff3b7NDB+9xHm4/U+rKBuhH4BYagIOWzWvFLx8BcE73JVAQSQ4gVkrheReOyaGw8
+54eQHYT3HHuYFRSIEGP17LBXm9zFKI23RB36hyBDXvggTRaBSgTWt6tAhEmheb7
qstqndIh4++Fewfs9+5iM98k8qKM/JsjhJ/e/74PpfEt5f0v/LKsj1RbxyVwjtea
qjyEsMWYN3SJbPKdpC/hUizahVwWlyivN9Z81fq0xf3epG3D+0JjCOUbfVGfZrIb
KBaNi/BbXi6IssjLa/c0+96tMKAdj9eVDxKzhenqjRV2ktXsStWx9oN4BgQsC4Vw
7opCcfL1lJkgJW3skjCXEW9x1pvjwpGbc+0OG3gGDlxT3pu4RqhxQvXgF4F3p+rJ
HWgS6Hl/r0HtOKwB0IYv0pwlphg7RYexIIybyZ28vbZchNryWwmth8KYMR3nV/1G
7X8J28HIWBJSy4HCDOfKmBFM8t17SB51Cy4SS/bNaulPcqWvgQXIQedqy0rMb1zY
pc1mePG2YxSF5fy3bGqyHCl2JcXD0lnViMKjn8DxY3wzBEQtPjvrRZ98OdqrmYOP
VcVxkJuk6/EkG0ZQujQ9FI6n4qcWAqe83UKd9szNYMvtnlYGXLsIDFN5/gLnA7xS
KY1aDMuW6O6w0NGwBKXOkaMNH98VtlEeDe+lBfdUpjMO9+44NGWpw2obeGktZcP+
xZ2eKM4v3ErIL6ju2X8whDSh9YGu4hRn6/7pC1WRIhB0PWBlbDJBK8TIZXCgWgSG
ohtIbIxLP/823AUSY29ZbeNmQe4szSEvqjflteuqmQ9BlMhnZnr06+nA+oT1wLZx
AXBJFsH3udODQLmcYXCazC+sl3pZGczgY9xC3dgnUaC2+xP0ufaUu+bo01kXD9on
1UGRxRgSg2gyfBOWSLs331TNGLBDSPKOx8JpAWAflmh+xlkKLx4F1kXnEUPOZtuY
rEYGFAPzcQNuFiMfnWzlfTbGGwqM0mgFAZhx+ZbMpdX/nN2vpZHBl8c7nw3PKVqu
ng1nYoVKvThkL7soJuXw7p8gm0AVoWt6aEJ1rNVz8X7Fv6FrGZkz7RpjLHJqBMA9
5Mj/kdaPTCCUsJHWqEx8R4/X5tFySqYlUr+GL0/uoLQ/br1ZaqsWZCMzyQFD0lS+
tgxRoNSaYo4fXjGRPj982UH6Un1mxZlpGebVUj+MUiPOmW7zT94SfcxuaM6kIlEl
oKJXa5RfEVP0k6fHMFucqQhyz520bLBPoJX3a8Yzr8W9MUhNxKDh1yqOvYcs4ASX
VeZY3KipOQo0b/1vycGKh9Me8X9hoOJfrVMRQ6WOm+CaqsslSPGlriOa9t12OtYC
b9U6ufQJV1bjiA0ZDFGthggCRU3iMxj68U9cj/3Yjozh5JDdqUPKpKkMIYzbhqi7
EV/NAvq2MoTX6iLB4UVRaurn/S41cjGSdkP8YNonyXlbp4VkW92tj5ynjndUUPH7
mHEzkek90ay8rc3jUyoaAAuOFGN6elxyK0OYdsCdhz+S8JpY3Oa5xbNRV5zR/cdx
DP3zdIcNEVC7vJVxyrg8GcLVDom2HM/axbu9PtdU62CptDNZF1pKaLAn7lz0FPrj
bsod1wVS3EczxQyikCBLKiCP59SDdB0XYcM/LKbcYmhJeIaCOME677gNLppdJNEc
ukD8TB+Ct2o7bsbAxCT4sV6KCF2YYjSwhvSVs+vUn7QH00nJIkNUOyBYrm5WpqMA
wfBHaF6XjZW/IF58lLG10wXa1jsdiiMxnFisKRsuxaLMKkow0USxq2ZTBX/1KCSE
9HOC804UEndPxVFAMSdm4KM6CAW2khpbq8z/bU8EZt+pQEiX4MSD4UcWmbEblmXl
q0YxyVvpqDQVNBHxIAt/tsqrZkcQWNJh+9AcM3scgshjaQXJ0ln62JGpZ+J5ra/M
PZ11q3pwivrbZmIdLuibqvjXySHMwuiu0ps/3pH8cVXqkYpVyXat9To/2M99Z+mS
+D8NZx7UEoMY6PVNweGjbw0WzO/H0ATATlOvbvlYMMGLD1lkrgvrNdSK2EjuXC/f
ycyzFdetICP3ms9Atswbnebael7GVEEvVYsdz+fBZPBpXujxOqkooF5DH9uBskkb
fQKujWPAuhfBgGE3XZaS3m3Pa3IZuXll4EnG09GJAqnmy9YnnSYlQMWe5ExOjBfm
xkFx7LwNCiVKNXuBIk6FKIEPicKMpJnKp6X2yx9s0pwtlYUU+BjOU5qBJnQ0Piu9
QrO64UmBrMuZdgRcEK83VxBY3StwUz097bVa0R5iibzpJiKMaATkQdxe3j70/p6D
DflM1PVp0cvWIyMobcevX73Xf0h7Tm2Pt5SCmpQnLZOeNKjQCJjcAB/h0z9ytx4+
y20RSDG05rYY1BJlqhCnQBReNo05TbYzW3ohvgXSLIpsJ8BXABt9OVUFVF+tvgEQ
9NloQsy4HfiDPhFD0ytkZnOX/hGRoAj7AKiGTyzPCYcyEU/DcWWNc4pCxCkw8pO7
c0NAwvMXaxOxso8+uNABAu6heWwJQDLKQwiFr3lbIImPY3YhFm0sEGu0IjuZoiLo
xGABlw5LEtM3WzcCUdetSk+18R1GwEsviSxZO4bRKhaqTEb8sJfBA7XVx0zqZqM8
0cCUzTt/v3GUcTizk9/yvrD4EwX4Fb2aOYMI7GsdZRas1IjKV3kb+qIVHOulpLtT
rCCEh6JSf+6ZkecYoLWtn38Azrq4b0UCAv+VVukldjLKvE7MYX0DmhNTvVO+zFb9
q5/4rYq0k8rQ8MO5SV9ILMWuWHi4SP8HYK6GJYnwr84mtdCxsjIvaYykOpfHKMor
nna4RvITu4UFRP+8zp/Acdp3t37eGG2EEYUDdIqLu5k=
`pragma protect end_protected
