// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
a8Xrse+TjCbT1xXqYUbiXnQmOPUpfy23iR+27bFueG41sKzZ2c7d51JyKN5mquhG
ZXX+6ooQuUXtQ3ihENmG8c/LlbapuZLs2irIAKopgjBzv62eOpFryQibFs2LI95R
cPfvrRNmGgDf4R8MiWoNvm6rNPaKGrNBTFp2n/7Yaj0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14416)
Jwez72cSeV2ALvk9KdE7To4te99BuIDixm43rOi8bh+wb2z4+tYZC68HoCW0Ilur
APLhB4AojS/m6oVvpqNj86wvgeDglSNl+AJj0ixWvDi1aIAnHik4Ao7K7Uk8yN4f
7bkZLWostRY4oxf/1vBN+UXyDmCmNOv+MtC5KQ3rC7n/DBxIbt/D0Aafb4kkeH/Z
8aSV/zFgqPIVr/+apSW4UgOhdYCcU4iuLYxWolnl6Qqs9yuDVT0WjUVzltNz91Is
9N6oSiQ34J2jW1M02yjqQG/bAbE9DFtG27dcFIJQji4XacZ/kn86ZWjCP6cjPS+h
y3CScSEqIK0HZ3GBBIj1XKV6XlEZxKHrk3Dw8gv2IxegkfbYEZT0CsJN81pWjAyC
1RkPMKoSprfiWYo7rSxrx/knQxwoOKXxyu9aFRoPBVYl1LUYSjsINB5eHGCexGfv
fPJB3Dhx3FfJl3X5g2yarCE4k2ubjVN4Ncl0xl1oANolgy67FvmYW+isw1ufJOk4
dtiA3Gi0BOXjHCnGvWFesxTeFXhozQfgh5LLYMkyQHnE8PhH14dPyJCZnogbEGwA
DrLyfO3bNm92q4S9AQ3Vnqb4oCnkWe+MBiPFG4VDX5RllSWD7OIpvEEdGlHsaR4o
NMyD6nRxZUA8OOJiFsAH0nkdeMruKVIcnr8U5ZQmWy7fCpnmmMtE3ylwdzmemHuD
5YLVMV/6evqxyEprVlR+Jj8euFVKon17I2VmhxaYJ33TD18Dq05vaXgJL0/AdStT
t+yiOWUUnziS5NVJDlh8l6pZZsaZTg4xiqreksNyNNZGrH6hZun/dkwJ4W0vd/pz
ha740HwlkB7yJWXhTqevxy9d2POtk79WVVwoGddNm91qZUielv0/ecUBgaDiLWsz
OIyiezSJddCByr2HcnI9LKwSoJcqt1lss/17tGL4aegUJREW3IgyMSSe2by3tj4s
tD3TRw8Y6Ai46npUvzGyVfSyXz6NIpVir9SzgixHLND+NyYb3ziZct/qiXaYD5ai
j5qxqw6UPfhvNZ7FwR7ZuEVZdhhtYs8WGyXr0IUGFmDDsNYfxBOZMuWPMGRchBub
qAMJpJCOZzAVD6bF3ICajA+TIs4yxsSwd0XAvm82C9fV7K6KsfrakiR0HdlRzzY4
iCfHHHXOW1aYBfrKQXdSXuRtiOz1OFqNP4N7jnbTaVqcua6EWA9XJCwm6wAOiTxZ
vhgjTp6iBnc7Pqw74Z8+93KhryHekfEw8GEsOyqnNeWuyb5zlpsBKPQJtgh6I/xA
uSDtRAZpcMEi7uCFjnyVx0k9ysdOmIHx6vIT2Q0FPZL3GDUBuOFylfif97FWHsLw
EaIhpaWCkGeyrKXu5H5Mmrt5mlVl3g+Xlc0Rev3/d7TV4cmqmE0AayMO012RSG4o
KfJyPUqQWjLCEClbLilb945TvcusXR4k3+IpNKDKqjGMcMLESTOJRqc4b52xL8Un
tATGyvfo5Fz8Xjih92m5aLwYBnuNfAH+eRII62A8hkDWgBbCebG9uM1lngS1q7lX
UbltuiRU7D4JoAP1IufxTAV5EzNPLNiFd/0AscEMUun+KSYwIexbIFXNv/1P/xEg
Z4aOckwpmc++e4xVJkq6Flw7XJT5gDaVOGBQoNpDqHVr1SnO/Mm8XH0CzZwiyIqk
sI4fnxDV+H5GDyDrsdEki3VaYvaXh6UmfA2QezO8os8zR24IwRYNEHTin3kVWqIK
TIa/QAumIPEaGnGakRJQbLfvN0jSYDGvsM5WS1BruZdnJOcct7nO9lf0ijz6FFS9
E8QwspBLPDjeOgf/IHmzJY0GRULaZtqUOq7G7sgPezUndDakoLpAHawOCqv29F+v
4SMovV5zEMsscr+iU7Em89HdWbHMSbAzdVfMuyuJRBXnZH9mMk8eat+liDnWljeJ
8e7UIk0Da/HALvrRoju87wfTTZOMi50WY2WdI8CDo+l8WM55r+qJFZAkfvV5Ily/
gc6JD2NwJVvy9WBr8KoLqR7nzbCgpaZdHe3+KzxKlKBQxd1ZFvPjxKi3Beuhjj7J
g+FDmCUYkZFKZtn6GQcfxCpUKhm+yytnK4lqwVaIC6tAFDUkCpKS7Vsy/VkYZTqP
kdIyV2Cxl4H3B/nnPk0BaC7rujI9OoeL1yy7hKgzytkG8yBJRlSSlm8kkYXFhn4K
Md7/onA44UzqdGDuI3QciC3wTkjz4XRVMysTOu8b/fdDpVM0MQXBIM4igZzeCOGH
4vQ3IorUAKS24OA0/S51Al+38d0GSjgvJDFizD7sZeUxHqiOAuaVLzJHF+kknLeM
Ghpzl/0Q/aLGevdPZBRHBU5R0TGRR9WAsC9VXkMQD+bYgW+K6ZialGvAibSAhH0K
cvN8y5rjsFln9Xt+WXt9viEHYe4L896Ot7iDhLS6wQye+c0CbulnfGV30unWWNjT
CvmY+FewgMCdIu2jvw8a6T5f2p7TCeesQjQWteyq1OzfkOjm7NSPbGDDM1t+JP9B
sM6gWtU8+WifY7caCw4BumkywkUXG1Enk0fYZ21WKJCoad1+2ASjzUL4HqcXg9MG
zPe7RaHIdNDMCePPX9QlixJUydDMZy5/jjYKejIfmtu6jNCbeU44H6vKhK2B9SzL
3cLVCuXdemruPcjv5/cWVg4zw0DjQU8Coloy6G/8s4oe2EZbPnqwrITSc4rVdvE3
iIT+8agWnKQsUtsiS5gYKdo/bT1ZOLZfVqyqsG0HHP6lAGKzq4TYDNV5uZWu5HG9
l+YX5b09oEpljlo/OgpMNTqDy+kjqvcCFTxl82kZEVRLdjzLn11iFQGOmtseatcD
4Rgq1SMFS1hh4aVhbg6+I31ogWMKq3+jMed3AGoTT3KbRKqsw2gPrHq9pIdEAfdt
+9IF8+iy4eY+3AKhf1EuICO7rABo0qTQct/Li4SRAzzL37g5WS73R+ZX1S6UhleS
94UGsmpuAMESaEV+fzusriKrEeolwgIigi+zrHEuvwZtDcs0cj8aKvOXP+GLt+RK
Nf0fkfHjEHNkJSa9ooU87L9GG3iE000vUUSIKeAvIbeee2ouYwhGQcAK+EEFGDJ6
NfH1be+Hoy9xdd4DFN9bHxWYb2sshQPT5dPtJCz1QqlCr1vSe7auSzamcwNv6Yry
P2wzGutQGwmBc1YWaa3HTdarfDBWUTs8RWcRbprwkf+VBThp7uSXFIYMV546MZms
mHnFGsE+ipSL1R/YcIy9Clx5y4KGqkmb/N6hx7HtxF5QbbFUv6Qhh5f7kQGAaO1w
TuYXgCnxu2jS930+B7TfSMDsi9V6fgwSWb2KAqUYKf9GKpAllMc0CWOjVI/vIyrZ
DYmmUxtSER8R51V4gR2Nc4IzGxKN0QE5bIjlsBVf9AAZwfFrVLegIhdBsV337jUN
B7Lni9GDxCruv8+GpswZG8u1781gbrr40tm7nKevznCcPIOuzVvPA9YJj5Tq5EJl
3H8V0FwsLnyLUuGDMKBFrDiwdHAHLcfU+5vVGDOFLxG4pK9bJo/SgCJpLd/AQlwU
WVXKb2oJ4Ot6DUwfuspM95PzQ1xpXGEwHzCls83T+eYlJ47oohLXQBHHv1va2h5O
HvWYv2MRnnfxQpjabFno4vQ++M3PvWJWcYs9GXKk9dbPg1kZFBXi/ECbY9HkDKDP
v9/abBdz2iK+eH2PIiHbj6lfAsxVdvViWwBa4ESEuzSmap1bKz+AUoxjxxKOH4zu
eqDNXVTBRn1V328QcQzBpPOaRLjREF/9yNpCIhsADBkA0jz/17wgH6lG1psOvhuv
f6gbgUoOy4mvm4+dOvnEz+ceLUL7bzANsQfHMYAO59R5r6LSpWRiFFQP+5Xp6hdc
Xm6dIRo2CDlaPWj1A8fw0pIhrlv8EDVqbJJNt1Nc1x6X1pyGShAQyna9xe5UDtIC
GD+fLynybxLlsJgwe768BNih/NTZhKhwGNubznnMPdXr4OT5BUufXj41T4x1Q8wu
r2zj+uFF2b8UvTsbfEGb1TrCPsMMIPczriiY8KeH2xaf2u6SkCP4IX2iVqY/I7JZ
ywdr0uEJ9PfXM/p88FQ4HJhiKKdK9mj07DZ+4THjdKhrG0vYHx1aklRp0a9dhw73
ZpvAdYcjFzsL1HqkKT/JHzPk1/AeUQG1Fj1Bd0noAL9A91XNHBNGcZgbZ4cs+Hed
WNcSMgWkPlBdKwru/sm2ThmaYCc1CBSK/UoRJUR26h8BLhF47M0/dTdfDmJmoDTw
tOAxXGpxfr/gETHN54aLzO+HwqqIibf6C7FjTO/GQWfsCsvameT5M0zk+j3KgAHX
k9J8jA/wZCeJRXltLIL88uNcIglmjAJHdp6FE89W9Lh10Cgxj1cJp6Crbbm22A4/
z7T7RqRJtNT+70G2VAnaHpVjroWrTHmhJlhL/VjAhx9C9P/U/gjWlBDQL5XS35jz
a96eZ65o2pslBcbLgG/nVN4XgG22lfmGz7/gbK88MLMia5bkmz5qvmRAFCmPvjGR
poS+Z1OnaTg9d7EREBP8gk3NoFHzB/58CbzW/bpIwbSJOcw82IKsHt1HWtD+75kI
ftkxBmONyJSYVfUa4gFz37OGv9u7vPL+tuO3WiVuTYSE6Lr8h47N9u0b3FM5ctAu
W2FKq/tAGjiPoVBZWc6NoAzXzB5y4lOXzlsPsfS7K9FsNz+zzx0C+G1DK5fVmyfw
enQ2FurDAx86ppQjF//oqyqe1YslIZWxcNTIe3+nk8rqJflz7+YdG7U7bn458NIU
3LG5JHQ6k7WIHe4wqZ/R0bIgEhtRUf3qyaj7VPIRQI4w6Md/6yI5PHtX/RW4JVuK
j5QM70KrEOhxt4OLd5cws0aJZZHM1GPajVzdE+G9mvqAyTMQbUvdWUWL1uZXKIYg
rm/m00AbnZmGAhumiBIdsGwpDOdROu8TMlps6ydwOuXE8Gm4fkEN7ymDorwx1qcY
5m0xQfuCVra/mx0oFkcPfiAGZ0pbsTkhGSswEHa5TVXMyCuU5k+CqpfualVz6+EA
Axa9yvdsIBlJdsiTQ2nSgmn4YOcslbt/NQwlNrXOBkO520q2WT2YNAXGzVrtNMrm
totCG/4/AJBrT4vnqXyJzO+0wYjdTt5B6rfwV3v6u8TjuaiqCtBPcntPQfbbYXQ4
OtXYlqZQN0WiqRCxWM1Uk1cyJfVVtC+GtekPQW2QKHA0V2eVCMK0sx6hPGmBgoQ1
9zZZDdbClkHVEUdzg7LhB46tLqLc2BqEVTKhDhQEE2b9UA8E1FTpI9zOJw9pUyl+
XWd2TK1t736NLHBtPj863CRtFHCfMrTMpfb86Me0YkbhZB7x25/MsdMO5r6Nly/+
NUssh0uuGz1vcCfGp99/QV93xQinGPATvpwp/qSLCafW4szPKRUojindt9rTOAtW
jiXJzXZlbzFqjglGcafQQkq7yyXvqzgVu/Q1HY9iyMnh0yH4jKYZ8ZDDCoPtmd6D
CsdgAxfK1IbIkmjQ7NR71YhtHaxL9JZdKFnskH8Eo8v8G9X3gDMqlQ2kvwq9lLE1
w8rRAEkqChmbNA1YinnVQ3J4RqK1G+H9/h/rJK4GzhT4i1h4+QmQne3Q11fVStNH
OxVP66lj2B7UtgrQplJQsRC5RZLdYXQEM2JgFz/2j/ZyA30FKFDtfZ0Q1D/uKWWQ
khO4CLfd/jYrM0IV8QVAZZxM4pwwwR5MMCUuOMRXBuIs2Wq2Wv8BRmONTeK0IdVk
+SJnfTFsQewxQrJoVxnTrQhRipFconYlzNjqIvpsspEat9WWt+ZOWTTtiLxnfu8f
p2s/w4DwMAfbbgoQX107oRDS3ilLc8BCgmS9cOZg2osjhiDaxjK7udP6jocCbq0O
kYz1LwwyBRlhTF7a4stXdhDXC3mSS3ErB3DTrImYMvR/tEG9e0n01gYyprnRts1t
uUjW0xDvJxJuIS5Z6cAeYsPefrKLqLjs+haBTlQQWZFsPUfYjzdmi0nqfMFWjdpt
NP0CmF7uj6DVSsjowITardyMMdvnmOtu6NJ5KDiKahKbg+P5cGWTgeE/M4fta6Vh
nauEJqRCljtUSZcKzPPXZeKduNmZTodzyfK6Ldprs7wgb7mOCsfhM7d1A8cnoqFl
mON/SAysihW1i/AB33gd2654U90f/e+/rxwrVDto7XKY4mYUl91n3hfbU5XcBVNt
VgYZ+LzLQWMXI9PwnB1+p/ke3MYrY2JyHlP2v0e0hHiB21H16kfgDlDRq/7HTAfy
w8bq9X0eEtExbBqd8Yy/yfRvIjvDvevUFgm0+cE4eIJYsgCND75XpNI7N2bQYGBC
oJyIDSefE2bP5Mx4qk4Co9Xp3CBTY6N8flI2pzEQzDhQEDdbycNLVSSXBWqbSQvZ
T1VSC0Z6sJEW8Jr5k5kPb5xPSz41V+6pjn8VPakzo6F+tR4GOuGnKMU7gb+KwJbf
EBi3upX82/lgl3F/822xPIcVNWVr87S5XT6i5wfQNkWm3b25N06mdoifM3qyNgGC
H1CT5adyr3BUsLsg4onF4Mq0mMvT9l/BieVf/2vkv5ba0aoLsVu29r9JAzTOx4LX
D+UQ6oi4XgYX6Kg+7GMUEvSwbDh0ICZTCbzh9ho0+vm6vTfTodg4qnsJBj4beu71
/WGSGskEVv7JM+EVYeKwuAQ1k3EOge7lOJphYaSUC0dwP82Cpx4YQxazLwp91V7K
v3hvgsHOxDoAM3NNElO1x7tQYoufjBduOMZslrSNBfcPLEU4HBsjVh56LDp9RXqD
BB/vEipPOgdwkQus3Lq6+UzcHQszVSOKaYM8I2EnDYHJzWGynlNqnLclAO3Tqnco
7TTc69kmcdLyVnosFPYvzc+F5tP9jq5ASi2+VKRDQgA9OajiL0tycc15B/VUCXz6
0kPo2u9fXFqnd3w99stdmePHv8Nz21MuVXOBAoSPGFyTvwR41m5EdQ2Xs9Ale8x/
YUD5uSDsd4/oia6z4GHUFidVODegatY8sZQlep64fTY4ROSolaO0C4MPFyQMP1nE
XP+9QwqftpcuNXW9TzV3xs9OUuyW07jnbT2oGIGvTVJVpnY1MjJP0eXj+dVRqUuO
lO7jlnbGx60zhzThyhwaHYqDjrwTwA1sQa1qT4LqJtNr8F8covr3WJJEHgO/uJMV
rgsE88Op2JIp7IQsUxh26jdiJ2dbv9rgeAHENk6hl5ysy79PWARctjcp9Ig61Uso
FYOMD5YgoZxxamzceocmJoLVCc4dbXSg3MmxVqr0UxEI1PO5TTBLmyhzVcshrdE8
eKPiRrCXIHUOb8V6uZaP4EYQGxGGoTGzIuFK9GR892CvKg2B7raWKNEEuGH/soQu
gWnB4ha13q99/4oPUPO/Et0f2UNZz2IRwFc5twSBfuMTwAuE+YeiccswfJPn4+iA
9ohwEAExmdl3oLgcdvUvDIFYWxFsqguLEf42CdD+sI4wQLkJ6l67c4xXZMYVyC4X
mXVwCsxZPMkeQ7QDavqn/Dpm/s96LOQzSRWm5cg+r6wFaxBmQvUi48XTEbEInpsT
HIxaIMU0/121mbmS+lPZDveTWKqUIaGqi3kLJCmr7u2sgDhwX4HedWbFNTmK1A+d
TKhUkb+hEwixja9sgr2texxmxgHNQeLUJHh4JcA1glRrLN9uzXdghfwcuSAdZdgu
fCdExDkBq0LxQ4Rpgc75M4F9bOP7RKmnefMJzw/oAu24jcdiQZ+0JadV3pNCsfkN
DCVUF4UNELkfpalrXGSdMObmpVLUCQ2TEEGDBJVaeZouISJKANnAP0f+8uWqzmGg
vAn6uGqgUNijIDAUzUy674HnxguxfVP87+KtKS9TRFyDRX4QecNHtY9/lQVvSfki
9JEP0Ca9Y1/zP3Pu76SjdCIWsiPR6wJFHOWHMommSWxixXlWEx38U/bqJLrwuxfd
DyPVuhNIom6qMT0i1i7obNQJKMfbupOB7r6EWSQxut3FVWAKcR83rwvLHMRKkmdQ
OtkuOCJviALREqkyPXueCCui44A4TihGRlO/j44S8OohW3Jfd6uU2foQf1xCzu6V
rHT1a6CvbM3iumg1hM2Q9wv8rxJ5hghtuyqEOUfLlZpsaqgqyX5vBgnXtcFnRx1M
OtYqgtTF2PNIP84KUJs6D3CrVcjeihiLHURkmAag9ejdUF95ZBEj2CHZPEoqjqL9
tfGaa+dQAxe6Alz2sZaLePFk4F7saxnlZMnFlq7V7org1TIz5QbnwDlxM5/OFQ4p
BJe070nZWB1z4Kb+UJdKIuCtcstczIAdtuAUrY0j2VUfJl2LutLngYsgb3FuujvO
p5TMSAXievnVhapn3IXcHCv525ZeAQ0tiX3uOAFKB2z9+I8hjYn0c+/ZjTSjCLda
oj3NP9R1yuXuFxvzkpO0Cy22OqwEredhh/XzvrX1SP8SiZTHjQf7oa+HZmdBtSUE
BefhpjXBJqAhBuNy/p6byNX1E6D8mh8qUVk64grcMuOEbkKnx+AU2jlXXzhVkszi
pgLhrpVyWuTGVxWKOBDFE2Zdv8K8HP9OVjmsb6w8BQguf0WbDaeCm83qhY9Io1zn
X84ahp1TP2E6aiYjBy+mncyGuSOXZTmgGPnpnDICFyaIEalWEvSwaFck2T8+xOU0
pJ5e6hLdWmO0ws1sfool7xXZso4BO3Hxp744Kg7HzqE7WdM9t2MkbqJ+atKQz5vK
9jUN3oz6MzXwbzcUacPeBhAkIFz8gzeJ+rPjoHKe4XbFnT+n49x5Xu6kqqpekci/
dKtAyM+Au/5kxJXA/FJhJso4Pd6kfxXtWVyjXJnz3TkOXNS2EvxUG55ycnZkzy+z
CTOfpCxQ80fDMDYeICUEondD33cKh363Uhl2lBjaetOjV1sE31EzZMT/2wor/dne
qiSPHUeShg20mK5RAKL+HiG+ecKEJ0BGXtWwakP8Ks8msIznya0Rc1EAV5fp0zjX
au6mKOtGEuM+dkMy1H4c47DLag6Lgxei8Yg5i+F1AJ2Fm3q1bYhtNS3KAZUealgZ
7Dg9uikpbLZ+lf6KOi3KV7VBNKb+8Li4I2Er8HwjrYIArgoTcP9yi+keTEc/xaFC
32bwfau2MNLKehckc6vhEObCryHiVFIvFIfZhaboLeQC/svv+tzBm6hyPZ7FoZlF
Mbnf6x2+hFchIBmaNWtt4UnDWepgkgf3DY0mGC1ZBUkzYSWrL37jTM31v4Qxsv57
CvvSpntxLtIx6THP1PS484Bqy2yQDrb0C72jwslCewRjAh9a7VwABsX58S67Aw5h
buy9hW/lRieRHABiWiBtrcCIV3Mjc39koutIrA7wwmqBJxK1qGZzsNXWTEvA39S0
tN/QNK9XRdI+so7/hLZ45tc/1TIgOB64E+2/E1jp5aPedotpCjgg/xGXcGlq0uPu
4qBqWrDYZtkS6U9BLiomgSC0k+gkO0f6LA3SAXKP9XpvVtkwotP+5VhQJ2lqHnIw
Qf5wVoXVO5vkQgrFEp17NDTJx2taBmszqk6bpclUb22Evgt7r/b/sZqXVoV6PtSv
4d0HToTfsGavVg6h7rsNClvqQoKlTx0vlVGeIJi6M4k40E+PQ74qRzr0FaRp3oh8
i3LLE3GxpDDmZE8nLlksPQWy6w5f6BjifMX126O+OJydR8SneBW5nKanBCceAzOr
unMah/NORpy9QeUfyR2mWQ/YF1KWKLztmj1yfdAOwkkxMZTcC5t77gHpcSrAqeiu
wnizQH6CHijEi96f3anfM3MwnEr5rtWiP2h2RRixR0VmmtL8fbMVdPfCKBanlAX2
Wa/3siNedyw5usLtqZCLjr9+6wdt/f2E7JbCruQesUZ3WFCbynORGcu4GbYuweF/
MKac6XhkV1mHUv/dOL7TUc84ePdJ1HfMveKO+Pt7dYF0w2bzCZohiLCzqqYl5BUk
ff9uSou9I8X+YoLubjHzBjdEfUz0fabu0wTJhav8vtaXC0utYe5AMcMtKDrGWwJD
UqgeG2M1TErzeKNyL1BnSat0VQUNPcb9u7OFGSYB+EQEg+clau3vgmb/zltUd04v
cdB2gZCu8qJtq7C7L3EWmjsZoapsgW9Va6EgqH1FovLxyfByIhb4VjHjtz/U79GU
c/v9iBqDrvkD5Of8gxeR57uZNa49e+csUoNrUAH+i0BFfvHWxvUigYGw/dmcHjT0
F9sTIvNX4JDs/I3LrXCc2Z6WSz5nkTNy7LATszv0Gkt+zOimY1I0oNyKpUJJSMMN
o2DcEmOHpWSu/kKQbctHrzaX1aTwMGVjOXARYx5ViXsIhKpEfowApEFOj7RUc7kZ
SPp3Gzuzav2HVvxN45qaiBZqdMqGkXu0J4xGzewa13IDfnw9dhPSPASEcQKSS51D
GWpiokirONKM7PWLcyVO9EA6u9t5D+kj+TmqjdHoAwq7qNJ0XL5Q+9T5RdVc9s1+
WowIedEYbRfq/K9YIo45X+x77cBvPwOcRqDXBcEYykgJCH5xUqurxaHyt/PLGJuM
c4wKGNGMKZKvjXoGgb4xYxT0vatuUqlmasJTubhwf915NywZg+TgKnYhxieCIrqY
gJSUNEQ0j9HEBc5HhkPevt5IWpun4nWcYXyDSsMIQL3ma+KKlnAFVjQ+1FU5e8oO
Ob45i0mOL4Bw1XM7AozjU4i+zt9o3wHLT95CkL4EUhH8zvUX5dR//0E1fZZxuxjF
Q8hxFkHw471hX0UDVqT1aP1LywDrEvTWgrf+4RIKXw8ERxpJKE+Dg3CfIuePR6hM
x1E74mOiapghpVDpCYcsBVxTgaFzLNREiHyDPXVsYDoea9T3KkHgLK6agmoh5Y50
VnFKKliLPAU7wiSNZ3xFPMCOcUxOuSEiGY7YIQk93s5h32vw5A7Et3wiCMoEn21O
5WKCa3CZMwEW5p3dwDNs5C9nLb/nrYW5lEOYSqz2GSgHys9In6lUqn1bR/Or9PmQ
krZjyytx9UrtYEFp7FZJwMxHH+cUFkKJtUBIVcxNrU4NdUkTWS2XXGgFUOTUhbdl
3//nbk3y7In5IgNzldmzysX1q4q/to4CuoL/Z+7hjkrnwKIo8y8iHaJu5P6M08hv
Tgx6IkNtOwXWwbw092B0K6LkuE1cKQ+LXEEvjmee3thLVS7iR/Wq3UGwAuzGig1m
TawE/aJCqbvzbtt25YoJhBbVYgGtdE6qtC231yIDbJpzzYMPIqJGYZ7wf/7USD6C
15JA3c+wttXAlqD9cXQha3CvpArfHHYcLJiM6lqmgOusmazjHAGfQcRtQxoqHeJN
+ktuAEr2wwGdEHzgdcAydL3mRYsxLafEHlvjt2qlYiU3nF8mCw0vC4vt6IHOQRyq
zpz47Y+7KGqDu8RkuVuR+n7wKb9lNAIS5T1xdzOgPA4jbQ8hD7q+FnDZelXU98me
qLdBy3VGLZGpw9uSdgmIWkUxX9EkoKWc/rKo/M9IgWzhUOvkCAOiaOYbmQvD2dIS
RqlzqiWeRZz1lRgOi2dP5071vYpWOz95WS5KVccMdyodlcLSqB7vBrKqTb80eK5V
0KMsAN3cP7f4ORjidyGqRzJ3/fsU+UnxJ8fmHAWTjdWvt404IN1rxY7+OxVlabvE
uTYbaYijonvFXSZdL+VL7vYYEBuHmedydP9xX3oTbiEpLUmOEEo0cRkQyFgiQnps
8qUFLDworFc8KDq8i8g+YFpErYclE4lDQjMBl14lWN/CFD4XsaU2lJV9Dny1Apyi
q/e8OemHMH9y/PfMNZXEYazweAZknzDAKJrx18sn/bOjWLTB2ejZKS3IGU9+1KVM
xjUVNBsb1mlUT7UUm3+fVMJAa8s1K1Op/QrtveV3RuTn+4+TlV6h7LbycJtjmAuw
mQUl26JIq1zZFkl5626O0Q69HeGhnmdwUVRidb0XG2Jn+ujqT5HSQVOEFZfTy+c8
KTjGHNaHtI2DHfaLr4kcytlMBRuCgG82P3fZFl/B6SdBw2vehWk6uqhvagUx8ik1
CnOaAftBFnApfA2bW5yrvbhlz35h0Nnd3sSnrgZxqiARnglOE5dpbxPRCPNBS1Zi
4CWB+8fH6EWOirzb/Oik0Wj03VebbyZZvDGZZqrY2Hw0Tu7KyLktdt1ieEG7oLbk
njYACnt1hyfOqwoVhkIvsG5XDAlgTA0qDcFFBuzsRG4HBm/lxeztiXWSRbh71+vd
hsb5kvjak5HYFsiOuPHhChhd6Vt49H7WGgwrvBoL9/vjTt8afH2QN1bjSUgwgL9T
gP7U/iaMGuwMltcAeh8d5x9VlwgcblZol+Mgu0/MSxB/A+EuuTlf5hNBsj5IT160
20wBruMUifz+q1YyoRH2k4DCFB6pevc9l0VE5uCr+B4qDQlTaLntTkPL1gj9DK/T
tS8nHcvZwbUltOJ0TSgDAoPDUEa/UBcQ7xkdFVDmqnAnKxughZqu3cZW81KCnO5C
y59uqEXDWtV2XtYfteX5epR4haEezxlvJmghri9rj+01og5TE30htRzu0YY7w9U2
nlCEyxqMHayQxBvKCaPBQVDhpPVp4MznPy1I4xi9sypm9NsSQZttDbEcqcBuNcC2
VBzddn1mZPtZMl+uFVO5MnJr/zLPpAb1C3TKTL9eSMY0Xz9D4nDqGoWLkk7SKxiR
uxsFz2ahkAAvu9h5VqSONzSI8YKJUHOnsRMTfyYLcrNoAx7eIobUV4D2YyU8Zua3
fj80rc+oBSjWOIaebOwfkmu8Ka5ize/JbFgXDKY6FZOH13/jbQsve4owD4TiO+fI
rfn6RD9W0ZnydQWHMZ9nhkxV1ON6gqe8m5zqJz7kr5Oz2DrY6T97B37Kjndokv8n
QYIOSy7DZSKJl2V2yIVW2cMv1afZoEqFUnxkfzKJz9CVxtg6BLukDh67cOpRrRyM
YRIrUfml8iCHNBk1Dblg4i7i2HjLRIT4a0BmyA2CemdS+383W5mR5vEfkVIWMUnL
X2NziFt1KCcglfLG/7doyET5KTtYfb69uOf8Y4e5PO49t4jM2pRSNcukFTzXydUR
IE6AmDbd3cSyH4oZec7W1WsooScKVqCWUuux6FZ1Piz65vwsGq4H90PdPCRm0w2z
qPhNDqjh91PwqAviZeyCYrMaOT5TC14fV4blE0QxaJzgGghuLhZZMIef0YPvx4K3
q8z3EUC3yyx6t+EjbFfwGFHNmomsNauaKC1Fbx+e+d9mQ/g1/AKs8xS/kWpS3jiV
8vZ/Wr1eFfHrlA129sZz5HNCublOJSG39Zc9G9eLDkjjLyfBcuGW0pA8HR36SO4F
THedPb9iM2Ta0OGxF7tkhAWtPKChqMa9BBZU1jH/vjwk+eBuSNJO2oBV6S+sKkPU
NRbjBf9kskU6AwxjLQJqltaSK1kPTl6VxKoy3GAWLdTnwp42JEO1WUwWj3FuVhBP
icyR7rEkqaeQxUYcYutwl12NAvYYifgrnLtlkb1fjbgxrqNWsOWiWGZyORd1Ds6Y
boIi6rhhszIeSlWklSNzGkLqRcpmufwsXB5vjUR2s4WTWNsH7YWjs2IJG+/zrt6N
gn3JWhu+0U1SmolUO+JVkATN6eMUFM0GKjrFuB/AcZPFdMPvvaYkHLxaZVWQAgzJ
t/GPvSwRdHpi5qG85r8gpa6px8V8KGPJx+bzwZfTcYoXinkx9+13h5nckMAEtNSO
1jPeD46JrkhOUI+MEJpt4NvBFGgmOtPEvMDLXcFplB6LQp+hzHM8szTJ5cLlqkC0
tiaB61q0VTwWgjQz49MaCSlrHL1AN1hmZleHYCd292hftmYlczKWs/X8NRZ07cDy
5ha9DdxZafz/zDwUA10Y/yr/zBwptrOnM/Yic5Vo2QGsVpF+RU8SQDgRn/R4Q1y9
fNzFN2ZO4qJXXqYyMR/NJ7+p1u5u8zaj3SetPNT74A9BCzTr+o3eoWXfEbkoONqN
2sjYQWkkhkfStJt4aLMoLdmcOmG632+8r+T4JvmBYsHLzCtyJiIohDJdwJJyXjw3
XZmOGahX7eVcaGEKrMZGKTyL7wwWRb6D4nf6QLeApuvYXWIwpAdfuI/mt8NmiAw2
X5nj0YtCdkBX9NeGPTnPrSgjSAsGtPm4Zep76CbNBf+eC2q2Hqed1bEgrZNZqV0Q
P57eksiKPXhai4iQtDKxPoo6gNqQnNxmb8qBjs8otRxH6UxjYXrMc+fmKmEwKcgk
OgI2ITz9/MSILn0nwz6c7NYLtuM/mzExAJCr7V52TNXQ7owypDkO0Jz2o3q6VjXL
88wNiGpe2Lq3EUnMlGCVKTJNg+25gNbdibLNhMwo3lUu7+LbFwdv+m5IfNZ3Nsqa
WYvil5ZSEDAG13dhwv7S7efruZB6dtmckrlC77OhXCbPwzBdPUaFLcntbxGFj3CE
R/zILasMtaYF/1RxnA89li01mmeX/7t7Vhw3FrCM6a8QCyuSzeg96ZEwrFa6GjnO
8bmogVhKJAdVIGIdSP7C1+0WdUhIzRYVM/MOMHFtKq4hn1Fhb9bioIJq30GzVBkD
MvNK4ywAdnpaGcsiNHYMNIcGX4wgjinvs/MKABBdq+ehCU07ub3S1t3F5URTmZv1
Y7/f12/HCcgzcVidW586rX6KFDsMW8KlI7eAyAE36FOydQmh1OhKxPDc6sBU4Svv
NBn/YNbVC2e0R2M48Kp/MMSOqh7Qau2gAA9EyQvI33EDIRV3K9/6YwFdo4Kwxl8v
QdjpSgtisdj+XjFO8xdGFs15W7hWpNXGlpyNktjCMt6notNkO13MWAnMLwhnQvVK
r782gqufJX9+M5ziTclrJcZvpjI72zRWpjUis1gJ/bJ3ahEez2jUbh1YXkwkkEj0
eS+n97MtYgBRttcsONwSaMsJm4SEQzNaJqQKwdGbgihyet8feZ+mLaO9qkrKh94t
3HIr5dbNIqmtpL3q7dPhRy7YLjmIHLufAefv0KQZNgcNRHj3jkd7NzJIYLiL+qxH
+z9tfOvH7TiYR+9iYp884N5T4XhunhTdZpdCdKFNpmQv6Oo0/qF7mwR4cQ0/iovD
rZ+1v/U0dUwPEXlhDsFW/5/nKZCgODDKQmsK+6nvxyGSCO8CtB7PHwEq6faxOCXp
da69tsxEC0VuiUb8LMTPt4E9Go15bmbYYCL7FlEn2qmwRw6V5hbSh6rhPdl8NVGI
Sv1LrWjI91lSdb/bfTzSh7X19xjgduzZaRhkEQmOOeDOooZmrb5lFxDLBYNy+yH9
Ev3s64ja7v/zkEH6zadLO2oXAPkcZWaZZFLWxXtnI5mz5XlV+FDzAzuWP8XXZuq4
ot52sYAbW6ylycy26h2uqE0KZtkATWONfnYeRLvc/H/mvJQOfuEbqWp9LHt+HnMu
9wDYltXXnauG+wSvI/UoID7Tg3gdZ0qgOqgwntJ1PhDYWhg9W8rumHodw7aoac9P
W4SYczs5vqjrltHpaZZQm/l6swXLA+OXXHC1zVq+SxPKMcLmkiqmgBus3GNgqbk9
pPdCvtHzcAIfAKcF7HyD7IE499RW94lQazbrJp8Ly7+NGYuKuxonUyuDpBPCuvwN
cSQSk3hPpF8KA3/gCxsHCE25heqqZfuVzSKYv/gtFeoA3jaQK0AzQQePgNqn5GWf
O70uf7CN7ulb4bmprq62BHSEPXOQTCLMj1k1r5eXfKRRe7/RW7v2qzsC3bfnMvfT
sX58r1LvMEEwNRn1ykzNKU5XFps/RX92u39tkMBFlEeIj2UMWIVsuzyp9yaswy+N
vD/5QM4i09EPiG+KrSkHiBtbnIjiLJiKvvTDmFbcdMREO3SvPB6zCw2ByYlQTUvG
8EfyM5FpTiDP118vHbw08aXSWBwMwQ2D4RphQKtNkis629LHYy03kKjjN+Szy7zG
z2bqmPAQXVpMRWrl2ddY2sMJ8EiSSiwL17GzHiWNSy1jafGoo6BAHus9CSjwkVCy
A70Mgdu/jKsyM2OfTy7j+/w+jIn6Z+Yx7fmR6SzU/pbu/7QLJWMM/oDHLh8BOKDi
rBu05DG1bqO5n2WQ27lXDcmwQsFy8nOLLaXD2ey/pdiXgsRS9ee1LUXvRbifE58w
9ux0ERO6HlGiDbWSOTntJcRJWeizn7TFf/mX9YOEOm0aJs+qoM64SAisgMwG0Dlw
5aXGlitN/9IRhytIHmPDRPul/5xwxhcnYsyaeuwIjLxcq1iPr7wr0Td3RLrOyvP5
VCGU8NrM3lwuhxAU74e1m8PqsLpVjv1erLGGJxeywIpPMplpGySS2F7PHJIvSxgo
IwFkPb99ItZuS/l5LxLOvYsFBzgTHN7G0hKHnp1/bB+7V4GbBJK99jZN7Vt7sYzt
ZOKasH20iK/Yt8YKaUbbaSMPMjwZQGRUp0LQAp4P85Z7bdhrabUQBgczZzOTvjZe
f4J+isE97OrcfmH8gol4DC3wiUGORKF+htKFxAdwtbmeQ/DWt0PH//8khxKX6GjR
ki6PwwIIYVPGOoCMB1pSYz5ZyiWQV9qf61P9fitYG/mGY/nzCfQAfwGI6vHGE5S1
Y2WQSEyK7wbriuWaxfFHF1b38uv+0SkqFnrKEQ3TDlMzro+Xl4fUri69IXHjOD4+
u/4FCrnwQwFI+JdCUVm9ZGZeMosvIVsQCWXTXpMM5aaMjje5asgIW8dE+/LvLNHB
P1bucm4pIujwodGNb5+NWJMcoIS1wRaBcibWVhPv2nQ9Tb4AYTTEdR2PEQdvDfzA
F/mk8T7oN1dpDZwoLLUNO+8JrHLw2Jjmi2D6SnoqQk6nhKtImMjwxsv6FR2HrWWc
+aXQ1F4TjWMHqlOQSmbiyGCjIrw+ZgGoXAsBdE33FZ/VgX4I8g0kweV466i9mIl7
n+BXiuT79lN2iN1BMXHmH/Y5gtwr/fhvLHfRyHtL0hlOdsH1S44q+5viK18dxGIr
B/1XVNjGee6oAufRQyKtNamzgCv9mtTtDFJfMgjTsjGQeJTolmgqYW/CnOH9wMcY
AlvTZkrJWbjiUbuPr/VcC6lN4+HeCqzXw9nInu9F49WArPmAq5IbNk3Vk9Ir4TvJ
6Z7fXumsmUZBJpbvfIpEV/OImLqJHgK9w2M1HRPr5TjXQ1sDvvKHcsLv+ORD/pwg
G5kwHHJGIlHsjqIDkfqIEW8znGKKEKN6Dve6+keX8Xp/b1ocXrinqfdVuLHHG4MG
JqGpzgBXYvC2mimQvFbcvsu28IqmiE1UgJvIUpgXUNE7UZRW4zVCEqa2mggyNkxL
jmd+KB/4TNUI9DvGQ+NTLvS8W1XFPEsxkZ5P9F7DfTdl9Va3u/Bvh6qWril/JKtU
PxEZn/Tt/hRNzlTBST4tP5KC5XSZxBmN9r+0/RURa1Wqun5lBPmDf4v/arFTUPW7
3QSNtL6pfBAOLMCKHszDeZevnrHE3Biqx8d0zsZnJ4KMg9xrE0izwjdBcB+c1FPo
B8M8cqILvC/YP8DLfvIC9uLTbZKzC3L/0RfRouk2bE7jS3UbsIHbO0z4yNPUVXBH
uucMiDj3zkVMCklP+hpBe4snXETSt3CJQiD6esYUZBipAvr+LbgiPpM/LpKdWoSC
13wBa4NLfj2K801Y5/T2Ps6fAASWemoBYNlk/hsOXSFxWRhq3ZWjXnSwjE85GRXA
ckpvwMOiMYHJHaawvZyIevCzI4+JhbHVbVsleTzPoUujrCBdwNrZm5xqTIyfxgsX
T/ywB6APATyFsCcWIFHfTD3v1e/aCq29CqKBC22dMzBxR749UXHPFwnL3ZWonhfp
8K726i2i4Reb1ccVAjZROtfUpa4jz/Ku1Wct7J1VAv4AohkD2T70X83vb0CHbgj3
LYIhg5BkRao6sXp8s/VfJUqZuhdvOYItYCBDXRiXUuxc4fRxFR/i3+MkEr7mzBGr
oWhANUeFXDAlbujhVQEZwN1vJ8Rt806izcwm1anoyKhY6AvTgO1PjEBKrUJfoRW/
CA/VazQ0Nof4Tj+vCT/Ytw/fCaiOaQ/vtcDEBLlUJXnEwtW/elSKBOt19ts2zxEJ
bmNsT+x/DR6NMiYt/tsJpsxuDophLeFdup2SEbpxKFBC3Lc2uSz277nnMcLqBFwK
JoLB+toOGlMKDVLVClwjcQjBxVLJqRkDaLTt2SsRmyizOFplglsIH0W91E1rpUoV
0Kj9e6lXdn7KDKrOseIX49tnjbDr6D3kI1HykppetS+wF/+grQeLMNqczMpyczKQ
pawUNssUocdxtUCUtjRge98k2ouexTG343yNWZmBvnrb/1vVP7nQV9gjX531zPVS
hg+S9e6Z2YyBsMGikABUL9T+Ig3K84BCHkF0A8o7yglAWxIFCff85B018TeyTmdk
68R7p6kTB9m0p2WNHyv7ebB46wixQURWVpWc1Yn4ozL+GMCojgF8Amm8GUdc0S7n
fnQwBYZYBqCJc/RxNUdkPduNFKod3ltCt7R9kPCpX2XzIcwNoQOSo44cJJwvENcf
oqwK9Xtj+1iXdPWzlEb95EJXLsll3P0+DZnjBzexIQTf3e65eOc3/5ZA8pI5uuo9
/TmrRggwkzXWIi+Nznfpr83i5rpSNtvS1whD54uetAIMoMijlqFlH+YPNQzxV0pw
gAKv2mC7N3r5i2D+OQrsGsRT6pBxYW7Hq/B1oRPmELankt7ZEBoE1NJmkbi1KOVa
Jwvdxx9EtGjAVRN2QzpmSA58TzIDR10GkWw8XL3mwf1lWYnspunRC9sWn7bGlhHs
VlF5xUfSt5xMv7b1elhIpetfg+/AfHmy9pVgfffJGa5sIx+ydGqOm2urFtR+k8Ct
b8gazkjGcLMqwx0O3m0Xs0ky/YZcejGBRylRqKx1Eh+RnMbQnR48S5qLRYrcehGm
ruboz+ORRi0h4Gs5aKLp38sMfBo34aFZDDQ+/X7GB9A+Uua5NhUhtD/jZJ9dT+Qn
WofANxAS3BCtZQ5Xqhfy2sEYu8Epy57TZio/vpunXRUFpZK8LFF0c1cu4yfH4682
zR5yxoRVaiVSL/7qjUgLSdOyueiVhqE9HdrkbPpcmqU+oyGLtfxBDYLagk/4x7oz
p14FJdqNjheoGUPrPUDbQcsjTi54vXiyQzkbQ7fgSDeFLjmJNIdRkdqRdu3D1uNk
RycNKVsPK7aQGIUeuoVOrYdKhuosEOOJnF0rrzwnjAatDgR50ZXKo2OMxnhL3Cfn
amFgbrDzGwkVV7Gy38C0VMOebBoAE8Oi5Ti/pkv/CpYDX9IsOdnfMxi1PFsjaFyJ
4OYv4GW+ipoeatdm/4u8HZp33Q55GZBvc40sBKNtVq3G7QhJUg1jtTjjFcdeHZtR
SILL+gut93LgDkkEFPcntO2LDQKuMjds3vWK+ZNxLxmH6SpTGWahotAMwivyBKCi
7XJLJonb4ZnOVolOA/sWuw==
`pragma protect end_protected
