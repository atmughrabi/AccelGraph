// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FBUs4zZNrpClE5EBIOYoWFyZphLbu3m+6nGtrsfyq6WIcxdD98Ce9/bKV44Ka2GL
Wj7Wn1HLUBYxpxcgI3eI2DaaYGY27Sfhd0xNF7qOvP6STe3WnSNliwjy94+ZNYqr
lToo7nlp/rvIZGYk10uVBtNBLGF1jN4IAbR2+CHW5fo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 319840)
NeF/Q/byu55cJC591y0TTIjVO23RZUJOax+xCVhyt16V2BOWknFpNsAfoax1237T
OW/VF9xzxJ7vQ0m1LNu/tu9UB8tukLDdYcAd8360vgmAoRd5dZXKhMVUY6T/cQW4
42hENgbaBkjv86o/TNsBBFbnX75r8OPqUQnflDRYDkI7aMO327OnrsAVap3RqRxP
VBTryqtceQF2alu2Qou8lrtgApcIHATv51HIgrg9L79dy2j+NcQIFT2wf2tEO5V5
rugHrY0YlrPTG46wEePwnAhGMnMPIw3hO8LGPVHXZmAJuV/o73LmvGTIucN4oEvD
5wRz24MQsY9FeGbPFumRlzjj2dvZztTCc+DDjJpydAsdBNcRmlkgadxbmAXvcepR
AOr9uNDDgLqmXImRP4R51/6jPRP3ItxbhLBEnjsTe2xxn2TzfqYu2P7r7nuo+Ngl
Btrnw//Au5SPeyXXXd1MW7M1bq9ACvw/mulDLoYjqmITAVEtnB8XcKKE6N5ijj4O
d7KZyzGk60g7LpuB7JpODqcKqsUicattZhP8rhD/nN4ID4RzQ60AR27PNGcgjX94
e1EFwhlFPoj0ko4BRcqx/p+28gsF0PmA1OWRtovXU35QGdXn8s4U1mNW4ymh+tkD
ZSe8oGnMN9n+Tm4CiIUXtBIvttZZGb/+PUBmVDV2YGExgYVt+z9Qz9cZDrjQPo4d
MWUdxTrHsOxBGeKtMymITFiDwl0vE/U7u+KFLkYGu29V6HQ7JZSbGn20t0EB3z9v
EWyKDX3O9T7IQYYzCrzvRzkD+hPbgGN0jSNAOMCb6TImHLX1k1OMaxsUo4uf3p/Y
+EyvLfPleIUEBUyzcZ0zJDW1Lnq6O1+oncF1cEOAXUOZTLSu6mKZx3lCmiQvj/ru
cnaJwHtHYSbmka9Kz+ANsKYHCDtMjsOI7zV7IbZdw+2O6gvHEH7Iu9OZKBElXyh3
F7F981LAvILwGmkHt2CtWkypgxx8VDIOHhJnA5QdZX/OptPQVhR9QK5kAg0RkV9x
gkaS4FO7dB9xcXbccVE9vyWESnDF3fBzME3sNYYrpIqy9JHyAmFAx8dYR2eRoVaM
oNazrQEhx41+p82Ld5aipJRaqVpA5BgKbR+DsQpnsYhADQsoYjLxO+d1kIMRj3cn
aMRKtt5mEGtXDzEMRCVaHeQIBck1nq0hVo0yNybXhrv3x2gV8FksBqitv++PmffA
x6UXMRqcXcOmNviR7xcGu8YLvzsbH+EL7eaOIyoZlmF1QvYUDwVKMeYsmCAdb8tX
ZwojFIZRxf52scTZYz/m5idwiugG8OdisoNWCgu9N34hq/xnhpYuYRfkZ9jPmLyA
LBbo7+gPngZKVqPNhI2aze7vwLyIW1C8BnHudZ6ocsn17R1EmpjdTAFOUAk1/MM/
cTfgG/mUqGanm02W+5MbL8RMimUzxISPanDrldd8GZxtvyvu82JRtPhBE5sRmQSs
zr1Zx2fKgg2hzTrLIEC2pxi8zY81RLit/Tp8D3Z1f9QWsQw4zHdmsuDtQwVeisJJ
i9lxfKT3SnXIybmUFkFFxlDe4QpgKTY50QdcHjnKyPG8YsFTLYU7PEHk2VKBz7fa
Mjrw0H3Zm1b/wt6hupE3Sv/esu7R5Mu/nEemOJP5dTR8TwnAdB7/LfEbmgCmesgN
VBxtvmj9NskmBzWtk2e2BLbtBnwrF3qUU4l6uI4QUeGb2TffZYpQshMRcNP4jSxE
KKpgXGkAbh6OLvEB3LaAhnbN4EMUX+Gxpzb2Vxr21pDCjejDZWiV6RgM/1v9bFCg
cVXWMlw3CVqj0S4w3UJfOqCpkRxS7HdwSO3SM609MPHTrPeqFMQ4JXlJsfA6SY5q
IdXzx4poKsD2fjRxuw0WqDR3nbVf9ZI0oOB1Y4ZToKPSZL+vf3iloF87nYCgttEC
sRWuQYMP6/0VJFWSsxj7QUTq237JwT06WbqmxlEHEkGo2zNq9Gu1C2P6Xf3lcgQ7
dfyzCkl9V/JKi4k3VP0gAfTEJmG05WnjYAc1OCIXF3ocwALY9JVNXyVuGAP0W407
+pCdwr6/2zSZx0WiOfRhGnValCoi59MUQKtdSuD7kq4nfns3uviAa/fKadfGB+kd
90VWEbm2Hb2gUmltO9z8Vlt9Spu67BmpMJzLageb8+x/+DCxJvDGYAcpEupeZnYD
cbMHXANHhKWoQaL8sMNyULTZ3rlwBnh9T2BFwkycLmQmOrXEZ+uE1cJQQ/oGOFmv
i8cifE+Vo40Sx0hJn+FalAqLibgZyP40F+rnf/jiDj2uNDRE0JNaCVI0pzaZr9hY
dSWiLlPL3zn/qa3CH1Nr4I4pBt+HtKtw6zRCANaFipiNBlh9J/6UPB2NqDGMERPA
kcdY40iN8hoCwHqymYAXGOGtbDF2EWrE0yfEAMuru+tr8Mt8GwjEfW/LEk+MGzNE
nX4zJX/KpJSrBHvo58tedi8djdlXJBlUYe46JZCwc3ZKsJ3m479S4AxK+60/gkZz
B6WRuWpOcpqmXAsJm3eRUMxApRBlhhIaZmp691MEX0a0RHUJaC8SAiqXpyVBTlBK
a4h3OC9y5JrM/AL9qoTYViADLeyMTtWe+4zJhJdLXD1kq+YbqJViyzx0IgZumjJt
NNbMac2Kkl2bsuRBMS7brkca09Kp0WeGQ+VAgtDQCxjzLKFbPhHH5I1T2cp+6Sjq
kRtubjdYC6HYIV6LI4xYbYC/zVLcMjbLr3bNGZOLf3+uq+UqAgJWLjvKBgNNjx+8
pmzOKvtbOZdKbcIqc3QZ8fFqSEbe3lkx1BTViV9eTOyZFz+uQth/OfQrtHOjzXX/
2IQqcXRnnU+rZbyHjfE0TrRXE9wzfEb8zU7xnS5AIuChHOo/MsIdOsqyCw3xa5Un
pp3pZpnr+CCUi1uSW0uCh2Hbd8sirse4PeWmh1EBDPzkgO7fK64c5HLSK3AVzN8T
gkggoIcW9LTrLQvMO7VlY8t1TGQP98FUwGlT5nJoBVGEPAeEhUJdi8amrQ+wMsdn
5REfbUMwPk3qZ7ImZHIZFyv8qlVvTOfjTuBe2uWG8btz9y2JH1ihHRhilul/x7by
prsptktdWGl2Lervj5ztwTMOrWJKUm2CAqi2KhwSuza7455grbmE2gw7RphRjfuf
9mwNUxOkPBmSYk2qN0a9lUnffDpLTZvKYXcBIkPEDUyyB42gfwTpp9M8iDTCMifA
j9ZDMEJOswrONHHRSGbsKZwk6+gCPWE662cKhYN93fcygq+M5S8k3Xc5sewxeXz9
aX2Vht8L38uYWZJTY0hqfIwTA3fEGlI2PafC9lYB9PCAgF6Mj2mk+ZHTYsl2Su2Z
Opn5fg6tmi4PfAc61yEzV9w6n8nS1csuGxowvRu8Vi0GJx43itxZJ64ezRLtwfB2
TYuoCcGLGczf7iQevHmqjpOtm9WyoyaMhYiud53TOidU3S+bc9mOwYSjMaVHFksJ
XjzAQtS9XoU5YHAsUCvHcjPjhWtUV3VVz7J8vqhuRTPzjAWk+HnTy9oqdcSQTmap
V4DyxagnYAm08LB02NR+Da0nSr4VcoK+3yeJmf9UPQHVdYufgbcLeSZ4CAV6MbP1
Bmt25dCJBXAaolXFwaW8rwoJJlL2aGvcEZL5V1OYyrU++oOzKXVCNfbXG96hwpiM
12xewa5jJwY5U9OHxt/jECNN+1LnfQRmjhSYK/+TOrejmtICje+vk+HXcJn0cfzw
yQ4n7hva6VPvyBzi9HTTb2FRCR22vQRPhXDqAX+GZG9KT0OFKSn5FEyqfcoEmvLK
C/NVRW0uKt0GW9cYlG8ltmqhPbzOTHDs+PG9pipPO8pYppGuU77oJpGBXiwo2Y32
QLSgOhC9m1rpUWzbiB3fbhK1/i3/ElW9Wc5S35Cp7k1cV3i2wllRaSIpKkOlh1d+
LvULQRgWfePqt3JfvqnWaJMpAtVRYSy+TjqGJKYO4cLg383DkiV+/A2ZvCEiQddE
0sGK98CzzCiQN2b+UDU3B32zCICJtNpUzYZj9F9tyPJd/gdFvMR7etcWs9diuqG5
Pr09aOXUd/aTZqp+4zbU0VRvh4VxsCWsgdcQ2qEnG4amXNwXbmWh4md/GF9F6vaq
ZvXkUZqsjnWYffu09uJM+PYNVka5Wx52NEnSQTNuh6sq2cXL9+y2LYiTO4ROFdcG
2mGUASltfiYyk32e3wdOmDkd70Hx54jGs6zM54zpYIWfjGwjaBg/PsWLU1HFZ1Fx
7izGFDsQZbhVJbSlY8voIbqyX7HQIdqFymw/JSBVFSeNosUDYl40AS9KSsR7QiLQ
WjYp9oL9FGQxnuUapoSycQcp19CPpd5KMOgi4I2JNIHtB6pRygmFN23S5sQ7pjwG
m33tG/vAixE0rdPUzBg2y2urRlaMi6n74Cu17kisvN86fXPrh6fv58znhQLkSKBR
BwsnedLlSCckd/YvmBw6C+tyXLMN+6+Vqn0BStDAFwZ2OiwYXtjlqCYaWBEjhV+S
Mj/pszJlKdu/3vJG02/tgI+M/Ju+4QCnVzC4wfZCM7ggvUOIki2uICsNzpfI0aRp
Q7mGSEuh4Wb/4Ja2JBie5P9Iwwlx7kft5rrvXAkJvwWdQ9ZGvuNTak8dgFYe5/rL
dRfEDqXU0dl2HnF/tOHdFhnv5v7ZtaDPcn/16rnJ+Vg/pFo47eOFrEHrYix7DaA/
sxloQT0f1xtswD+igq2i5LGBjaeX7tzPlYVGEYX95QzbNnemQS06lxIItH9+S4MT
ODm+bnqiqH73aZgcCFtUdyOqkK2MhkAsBgbopT5xwheM/HAoBhG/Yieb9ZXsRrMr
F3Gd3AYh0LFZXJT2dw4rnCaJoxfcKWT7allBCU5HKONiCy7E/Lp5jUef0hUUr62S
SfJqXuQJERBece+5gxgwrLcXwAHLKtBguD7OmgXdYQUru0Q0ISfoBTaLh5S4q06+
Mj6ZeK76loABoucksQzDoYODlfvYU0E/9oP8dXhT18PfwrQNdGjZS4aRDsAcldpu
3C3rQCVyNax5VIICsLtjFT7t4tOqUomC1oO4k4EBRbnpUjWgX8uYzto1/nwOLfrQ
0vh4VcY9K+nEQ0MnBj/ekoU1dPZInTeypo1zZIPI3MLlhReJC6xSXEdwsI10iKpC
ir/P72gKaERMyxOapL4aGjKcfMAeLaxMOJG24MRnaKUFjreKV+g90v+7gL5bPY2j
Wz/3PxW0jD+zEQDG9M+LwJp7k9IWBxGJSIXXUMejK8vlJh7nAKW8LLwEFHwuPLlJ
fA2sd1z5X1ryWsjETUYzUObfKPZkIDK1+jQ1kaxBg1p98rRcZxdEHwvv2Geu8WoQ
juIW28NY3TUncUwU4mDMpzgOpmsJEVGPaZWTDNJYPQt21HaSe0oBxx31dsb2qi9x
QmXe61Sr0g7+BNaLdaAdi7TCx278OhO20UiojQZV8HwO5B0+EFaJlrzJoAoJTYlf
8DfXUrDqabqufBwkfWrSpujQeIBld8znYGyWpxkf7+Lmh9179Fjk6eIG7EQiF0nu
zMbcwt+I+yrvQB0ueIRskooBCH7u8W18fkUHA4s+GApS2C5WIfUmVHr3de38T+Fx
3CyvF6zk6X9TC7rxlD3f03hHslKyfZpQvVRoE4WjQ65bKua9HbsxSKH04q4SgIjb
UXzNCQcbzaubECtmW/e47ebkXkCEOPekcmGeUY2Squ2ajaIfv01HlfHBtyWfrQmL
5JijOT0lOswJRc7MtACBXHH20oTXKMRTw2Nv3w57IRCXrQ/c9T1BctrJKhSC0O9C
Va4d2Tzx7vEpjemehveW2zB6VrKo6GlNCxuinLFuAxlR+3FY5z0zLpzfhfGVl1fh
Va0S0DoeZ+nZEVsbfTYWVc8AGUQGWeMnq/0T26kKBBHmI3uNJj+Pz9CrZAaoZfoK
qK9ZoHQLUgOVTSt+PMvANZPzqL0487MHx3u+zhfpucZ14816hMM7FOX5aikdfsG5
l9v1kYFrp/7kdjijBAYSbqvYSjz3u86SH4I+Z8GEyDtC0c1uITm/NCYOYFGARi7C
F89Q+Jf49ja46x5ldZrRThk0uMh8OTNIs7WgALYCgFkB4pDaniUp0Qi3Lg1Tbhld
0aJGj8KFs70oUS1e2+m0P4WOSeQtD8OT4guj4PLcxZACXgdAaZvwVRhgTJjFOcSw
AeXbCUFaHmq2YuDyVC957WtRlgdFTW7vxqWgPssVkurfLTUIbe+u1a1tp9m7tnwB
MMUlPL0LebcTPvwazXcVp50p2c2DOvQ3TP6c8LugZbiAwmwrhzHM7lK6D1gnzXMV
c1mJlic0/LPmo8Rp3ugTt1HCVBE8tF42WhmWXBRQq8gGmb6NJLxi9P4RECGmDZ1m
/jA5XHMB/OuxrKgzO6JjXkLaYT+cc+n+3otDDLS8tRbszHxlVfrmyChZt44eFulp
DLnBgNfY+yEaU0j7GtBYmzwGLk0SphiOaCbaBq7kHIXTDnntjt7O2TqgK7uuOfMS
vqTgN2G6MLTApSWQlAM15todQ/pERET5PB/hGpebXxfHI+6RzcIHdg5kX69Slrfr
hViMcbxbkzXUqyPhPPy5uGM5UdDn9lgg87Mq2suh2z/i5n5GaoGGx4iyjx5oieog
U4f1X8zy/3SsbY+93RinCvOOPlUWtwoYsD+El+97P87sgVf/eRQKQzTX5ymydNyq
L+eHG37O4XqLsexppZpNlbeQ/5TFqteg7BrQ0JiC4EltE4bC9fO6syvf+9YifvVw
W1TufokaHyWVZiGu+uuxRNkyT2n/JMmIHHs6CeJ61M0hupOk3txaIwnwHiXY8sU9
t+UcNEAVytv4YDRaeWy25hc4IDrxah6h1Gkx0UTabiQ9XBHbITT4HndQqfc4O8t6
Fz9kQV/9Hke1vq4xnGBoEFTn8m1BUtKVXlQY6pXxKc+VBMfTMuX5FI1KqlNCkz3/
qRRt4NGGp9V9L+u7885nZYb952aoLpo+qv/KuAN/cXUlwt++S1TaeuQgeyFWsPLc
DrAUEUt9h9Y5Q3xMtydxnbkuIUDqspWyLEZHYsckNv9KbypBlKqSGazxPCe+9F0E
B7HnP7VPQr2uPpxnbeBuG9VQowuAzFR4aHJfNLlN3nmar32+UNE9iZxvPZY4bH0i
Oln44z1wruax+IUJTrLcRNA5u5ywgsI+3tEsDzkGyeLv8fRN77+CYLNulndnT6Kg
ceV3+tKhhlFEhyCXyAshDIfD5J4VwoEd3a/7X+gPKCpE7PO3XucSFa3Kscr+y8sF
XIAbmJUT9LtDTdPNc9VXPDY/Mmit20irccPLN0rUQsOBHhdP4iE5oiy0eOpCNEKX
kLWyoyEJgdZloUfOi6Dk0q7xrivoueyu3kHEhu8miDk3jgKQ80EQbORaW/e/RcRz
ifUuIUxj70mRw5xaoXzjYHLIgCUEyyt/xb9+z3zI4QXn71mTZ9SFr5CTfhxoZyEm
pXW9IK12ExIjhid8wbkQws7jR4a+4aCFEDa+h6SoQLOKftzwNyOjlt/agL16MyNc
TRcSp8JEnxRvDWt5v/NfMhrj27Wx/tH5kv8byyXTuyXCj9m7Owga2DmOZMJDliJB
JBaGWLGk27ZdOhBonnVTIgyGZqJMLbS95C/+dWCzBJgEsboaWofV5wBO6cGN9ey+
0XNhxD5JPAECMdeMBz2Va6mcDjG5E1SZI24q8S951Yo0zmmk30bPVFAK5FbA+pC1
r3F48VC0iP6v+MJFrPpiEZkc9Xf8NNe47hK9zzi7QsjEaO64oTnfkrkiEm0Fyz/K
ytJqTqZEuN1nR1y0gdK3BvBzIKQED9Jtpf8H4XrZ0zV4E66limCDzZ3toRl7Knue
iU36OirlgHwtH8fOSoBy6xQMys+mJ/Y8SsVHy4251D9a5ADF4ImInKWLWQV6G7XP
GjIK934iE8sx+aqad7OXmO4JvdbKz/vtyhzFNxHoehX/AFWgIBYa3DkeP0OtCJKD
jKkYrQCofTJ9TBWDNN0yy2wxNredO4nej+IbQ6b8wdoT17B1XFeTRdaM56Y66Ydp
wsSgST+BmLt3PIyytEJgAJOtXkvehZ/S6y2srCkdYRZI1BLtLjKi8I1Ie6cdMe05
K7zdmxO3qee8pUDbnkTiA18SJ28PJgUU5QoNn2N2dpW4wbUy2Wlg2xkhAwH23z3+
/dc4/BruNwX25Ewg+czLnmuh0bupAu9FWMSFJ8VyIQaXEjdSLnmVWmM6D9p3/trD
Aa+KU1BaXmiiBMbB5+02pqjWlTGPsbDzgzGytzPfX6W7DwIHrPYMIdmcWEF8V8OW
9oFacnnCcj+sbeotGk/l/AUqq8HohighpJRBDqgFxMRLIF64Xs8X6h0r1SRYcWds
VUQ6CPE4YDJRNvcuLf/4fMj7a/hrklor7PH7BrhghWJsuB15uERs9i1sM9IUM2b9
uoAexkGK/k74QdLEzfoHfeK3pHzOYSr5Su3+QkOCe+0kgXd34eo+3vRP+PETrzX/
c1zyCiHZR7Jswpdtx4eDq6SGzlCAW34PVBGvegvJVKI/eMWXJNOXgoqtN7MTumkK
cmK9kqE5u6sW/pRRGo93akk63hJHqugdo/j69CrAjS+lvZ3gQ6hWK+wyPQhjMRZy
1326ELelennco+cjtp5Xm1JcI2010zNfGpsgf2qHBDBCpjHOVbIt68yMrUyK2V2H
Cf9fcaKZW0Jb4c0Gx5x5oiA/MtQ0V6ZR6JBFN/X6fL34FkBFaQvh6dtuRuzCzScd
V3jgcKX8i+Gio9vShBTHoFasOaeQefFdE9iptGX5KeiVgUut/2xOE5v2xsNpYgKZ
JCG8QBjG5JwWZ/wPDwnAQOaAjPolu6YMRvQAEJR5BPi2jh8iubpAW2NA7mRHCGaq
zQ3mItuJzvj614NTatB8ntqMmastWuwoF4nrCxP9e5FXi8WWYdmzdi20ilmH0r9I
MokTv59CLCjmhcQR52thn3VAVAX3VBSKCoLTk5br3iQ/2d6OpT1EFKrSUm0eF7ZD
9e9NoqA9sk+FN/qtHkbIicqXxYsJomgw1IUZap4RinrkIl0MlC/3o23zF5x4VRFd
n27vQ+lvOu1bvfZrh1fgMgZnsCwjpvESBh6ct4IKIL9uUyKN2a7EkVyXSfjM0stc
izHOp2rygyhGEzARIYWmFQJVUny/XbEzQgIZ6PzcNe6Lhw/1tudfuEsIpML57/Xz
pIihHu7jVZNA/4XnLgghfiwxWIHwgjdf39npmcfiwwbuSpz6f6BpDOWg8u6mmUS+
IACDoeu1hBIBhKKH+RgWA6rVzqb1HGqT6spk0krh8SOHl1g7ZddT8i7g8NeP20Kj
FKErLOpusiG8JqR+HR21gxIL1S5597n6bflo/hzSov8KtGQhEIbk0mFrLWXsM5oU
Tk9QT/w09RiPqgtCRVU7T3LlhyohskSN2Cjr5fQXgVn2sToK5jRlZO3h66kaOJVE
ztzT1TWU2IgeTg+/V5q3Ma7lrlPHdAlWeiqSukWRrEZxwWR5bRt4IDpy94ex+ihQ
4+1DP0lpCBLpt2q4jlVF11XxpqVQ79ERNJQhdIuGGme+JJjvLFI2g6P0XZvdgOmQ
3ei/f0vyX+ZMN6lqQUZvNAT7guGO53zcd7eBGWzIKGUHQNGWSG+Bm+62EC5fWaQA
q8UcUq/qvax8raFWaEO3TuOYJdMtnRlqBV6TuGsaXirUsVtz/YMcoBWyi2LUI0XR
fHuUzeRjdZP2k2jqV1j/A96CQvWDnjgJiKhD1vtjKZ7nP9xYbTf40ks+3iCWUkOX
HSCV1MuzVR3vVQYOqK/VToBPtYp+DOyNdle27oJrMCBJ6Ij+L5EIREVRVdO5YjbD
vbi7PBS0V6k0ZUb84kzDvb5ssS9FShX2/DPWi82sVHIYILHPL3/JFAEV6FUjH0Rk
mCsx//eNwM+yjD5WEuhwTyyLdbZLwEVn2LGm0xi75Ht8uk7yivJ0GWtXzHxdsNYq
gJGaHTH22L7cu6ZQjK7kfgkusaxBKeuB+An4SrV9d35W44AY8FNywgFq8U9URxdI
m6Cc+YA0yw0MYPEcepuhUGS9mT+zy0OS3a/ua/tIZvzGL2PnbvSVfmorw3xC3eOx
r5zC5gS/bttifTCyOP335ZIPVaOmrj29vRi/wn7wHnBicZDGkMPyJqzo3wbm4kPC
h2wuDp1GC1Xql2PuwRe7tR78fKqq+xudvEUMiwNS2lxty8rkr+ro10jViIfMUXhF
rXQJ2PjPPqIEWjUz+FtcYrxZrpvM6BLcgzzop7M/DlSfKJYoPCA/ZVVihkQhimRs
x/gb0Mmo+0Jg7xSNwpW9DWr7SX0Q3QikMUsUsVrXmCRnpDWaQftCW7qMCRoj4vEI
zISmU5iRKI63RbVKgWiGDoOIupDXdhK5Rz4VktjUPBh2koV0DtN4roDsld6bym7E
bO5GSKpA1I9TDrvqpyyqIjfRJ8Te4oowSXNg+8PqieFJaPeXR78AESRLgq+LdtKR
JONe0Dzy7dCayas76jCYISeuSS8qVbnnaXfHa9HT7NMF4eQThKBQK3Fh22cQqmM7
rq01V1dsS+B7H3ZanG3kdpFGmdc7bt5mKqLSmzPxPZ38dcKWxWjfduWzaZgT6yBJ
mt0OmLMaFNbkz+1w3L7HSqHHRqKhwaEwub34HefuNEERQw5PDvWk5xWYrZg0kT0s
toVqXxVpOjJLeBmso/NAL0YOTwDQ1n7eUN2Cw7WPMJUNtjgYtlR7+MWva5jv+tPB
5CipPppoE9/pgb345qrdYaIs3tOH100kI6Cq0muKv5v0qr1rKkSiDMpcP50WovIY
26INJlj5LoVQZgJEk0gU4FXSBQRnc/u4JiHp7moKB6X3OhZOe3dLpng1u97Dw8Lm
d1caV8Pml5tcPETn/QFRC6Qx2OXoXwXAF/KfKUNLKV/Mf7Sr50hadZCxFOTp+ttX
/rCaMUjv54TGk0YPc2v7Gj4CtPq8qXvI9G2NqeakX2cjublXgiPh/jrD5twm58gi
3ym+6FJ+jYBYkuB54H18ObYjZUdn+AwzypNut/qxRwyvytOiqriBGTiEq9s2pVBX
A+9j0BploFPyAOjHHK0uWtmbFaUfLQws0Uaz4Ksg/bwapTmc4s1z82d+EBh9gaif
D3WYzsGxD20EFg7LH0lubary4B6tiD+YiyqHTxIKA3HsdIFSct01ZG1mq8wOmhyp
3EmeRLkpeN3bR3km/afQvVb6FeWHZmd55tGFuOp4kmFIJF+dpQshSuRrE4OPcE3P
iREjRp5xh/sUt5gTS8CAw6XKpmKjkIOsE8jcBV1wXWJ+VvQPpk39DWuLne3BTet3
bahwN1IapzDlGabDypHsUQKmyItTVyDFbevgyQVTfwt90IdgEqtQqjNybaj7gggV
PtDn3kAzYZjRzp2iagKh0H9G5FmuGWN10W4AUfBoPYCTpzZ7nJzta9aXc+6+yN5X
xdWccHDTTyoN3/3U2KOrA1CJrtM9q60FeF7Lx3bTL7qTf51Steti/cBNGO485NO0
wZfnxXtFQ/xXjtY9KfQsiFTgHicvJL7MyeP6Tl7tucUVe5kCjYSfleV2krXpTe+f
FVDyzKBOwdtmqs1TsEllc16q4FD6yqGao/GZYnBppOz2shnOgiSuXANIHPXy+69F
H4l01+ixvI+ljDS1O2Vqrd1akv6y212jyHz79kgWrNThS0sM4DWS6pLC2YAOohNf
Ndsbf4/h7e6vLQK8aSGrgSPufQqse0xW7sslV9bYCiZArny+nfzEpzGiJWIvcVso
UNlhUDG6FYmswt9LvMOxQ/RParBizoiRaSZCHLI1YlkormfMv5hcQs3zN5o/DR8E
eyKSXSW8GlM3L7TBzlux874eCgpIPJp+XR1AVfAuVGNVk18GWw+TNiJOJ9PKIFON
9fE61VL/F0FQXwvatzC32loswqWHvtL0JE0WGjcj932unMh0Ep0yRplw2izHL2TX
ZR75tbiGzfbsAA+NgYu1u/uIMw5tr12oi95qUZ5bXRAwwApkg9s4equ6IvkeNrOp
aQTmh7MRKR8DxgzUWXx8Kiywr0figrOgVMZSxybY/hyEgN5ngPEKOn/3PxiPpBOe
EEmK+PyLeewDsrRfkdpXM/G53owi4ypyfzo3RE3fcrtnef/q+I9I/YNfinC/HcP5
/2eCm74zvbm5/kSOrQcx6/sg0hzxj967T4A+xO1bme7gZE5jEwncpXagE8Ua/PJ1
Z8hgJA3S6CUoB2+jAtg4iNZ69We6RXH60gvQ4uQ5BZDHpSHM3wtCF3TRJmEl3k6O
wzhxm1FFKeFN+6Qy2LOwIwdSrGK8UmxjO08fcC5I5pY2b9NFR9B4F0DhGPE9ts2F
KBZgBlEy9B/d/IgY+cVJvnMtV4tknQ3ZA6X7es1ImJGvmxTPbhCNS1kNfg5F/jp7
EzWzc3j2jyMurXEr+dG0es4m/9wdY2i0H86dOspl7yrlKuQ4cNAV9ORdKS6cLuj/
ar5TMXck0Ag955ZtaUklhN7NTur2uHh85V4xuCXAlu1h5V9pKR92ERtxz5e+mTGO
rX8hY16mg2JYwPA52dhUmkc+xdjvjTneguMcUVheT6Rra6ruu87vwd6+o8HYgl7m
x8EtGEtfuqrwTowiE9G6oZrlxe0RzzgTuqKqxiiz+mfNWWJRx793espNxri9iUQi
54USsXw1Xeww+8C6vOERZRt3FC/nMk4pu9lhFljR4C9OV4P+FLvdAmFzqKlxBFX1
HawMWGEZ7D1Ir9GMsYxuQut/vrupC0rRT3289yIK2dPhgkU2CpQQUE4XzTjNr0Kd
fo8Ttik5GBwHt8aqcO0M2HmhW70l6UYtjS+8n+/TYJUqwR1hURvw/fUeMerNDb/4
t+3fwsBL6S3+0lC0EK06g5dweJzOOQdSPE5rvC4pR/9pxHbDSadBNFcnKPGqOg+a
nzfusExs/K1n23o3YQZYlWL9m0i78bET4RFuGZnU3PxrGvBfMSyy21H/U6Skeqz2
mDzD/hts8y/Yd3AmVLn3eaOOFALd8ZtE4XcLLm95VgHTdEdcUnNmrwoSmnvRtGrA
7pEDlAic2nKcxi6BdJWzh1uvYpyp7TsXPczDlqv+Eihn8zXYbyL/cRM9hD38fr0m
z8UQgfO7Rf3YuVvbkNrBV6iiR+OesbR7AnFp8ntqHIYryg3mzaEwQfQC7I+fiSoj
48FXfy3SGQ1dU0FOZpD9fW+GFZyysjGmNgnwYqiGwgEFHq5SLUKSumuLG3M6Cbfi
5ib6zB+lngrG/eQFaa1enQXokCj2n/W1+2oCq6vj8sB5i9WdTswPAfYLetZ6MwJu
WQHGpj5eNt+aQK9hgy2Mrh7uLXisuJ14xlbrERS4Kd9sXGqFH+XJs+FmshE4ximV
sT0jWjAGDQjW4cAwLd0lWCAMHdUaJfTWj/1NtExODmUX0/XXvC9bTPcDOgRgLK9p
N8prfkPQ267FZhJ1G7etxSoE5J8qWRnxjV6LFIOgvL4w9JILqEBJfDOVLw/I4V+p
Yz3OZKWJ1W9lWJnXdLAMG1kvrfcrBCGJthtpS5PjddMY08zpj8+G1IxeI59K3DEG
eYmUyL1E1vrllsGsdNW9n4ao56vQ3S8lReT7dVBjJJkzEfhksH6pr6bdW3VgHuwR
/WY5HvEP+2yQFuJIuheCjwSeC6nmJkqlU8BOpRBU49Vx6KRX9rD30DltblwIbKVY
0+vtP/lY4EOAToQen2g+6QZBQZcILqX3o2kofZeGjyMsWxoIPDxMh5tcXJEWg1I4
dUKKFzRWkJXZtB6na3ocjd/0pkcpZuHiGQxFoH/cg16oxc4JvigAe8ZB49mNb+Rg
nJMc82P5N33mz/7z/jFiF+H9B8T9+FoiCn8IcdRrU9O+eAQVMVOoWWrTm+adtuTZ
vDHO/VWiXwN/nBBxmS8rILAgfgG68YpRXS/Je/bu+sOA1Xdn+mc7CSsPFrvUNpOj
Zl24kOwpziBQtVZVLCERIkN/tC3PJ41utfGc1tUs/le9qOM85W+qGqKbqvEfQrk3
gcTmowDyi6hUR+ZSrqkvP3YJRpkR47tQO+dWvWyGSY2WQwQZ2uXB1vj7xG4pz3Wf
PSkxilaUXkll0wGil/5C38a49VrgH0cx4HHrZmnZtYRlEGDq2nwXF/zfENp2OhLO
OFWKm/f2GWoAvbMQ9CFDMSshRW9w+FPVhJ4Ep2m1vyd9I1GmVH4EqqgmvFwCAYsl
mU11PJQbatVCCpU1pyG6KV0Ayq3tUZuRnfsa6erslkK/r5vui1DYfR2IlWzuWK8o
COZVPUyIkVnxyFx+50hY6YXevsTw8//w/wLz+aNUYxPelcizJQwg5nOjuuKavh8n
6dC5jtVfGzUYY0TQkx/+1gGavFkkKwZLamQaHFR9LVDiRfVbJnlxi3nw2rlRRZmY
Zr6OndgE2qqhVAO90aV9a1AbnOytQFgs5cp0yevg1i1zIaWfLdieQlp2RRVVES6H
sDqohh0q+3+IIAt+8ZBrVB45eMXEwj0SW7jD9GTgfRwifAWUzyhauTbcA+ZQRm0i
mJfDh3hjbiiKq7qPbzx7fUvWSTTUeew6tAVqtXb9/IgaEzRJdq0TQ0nyorxlln0B
Pp3sl8N5D9bI9cRXOS5l1xNE9cPgaW+PPGQ/p3xuIxto7t12iZrvw7lzzMDEiVjc
uILv5tr5GMGUOQljg2bxvdQ7sT0WIFf7SfXPbBhIf/9DSPRJIZppOX/trfrDb83R
gcJH0BtByxjTmIhjREXiF6jutn/6lq9eOD0anfrVSm0vB0J6wXnJLDg611YtTFoZ
mCQ6rLv7Z8rS+gJaQZYSdlUHD5qJWCY0Ws3Us05acY1MkhhNPsw8z2ZYxeMRqb6W
vjOdw4XfkBhe1ar4pxIcTCmxsDecaOd8HOhR57KQbWqWwFN+BHB5k5tDW3ffPWAd
z+lol3iVlN5DHyv5cKZH3LgE2TPYKTgDjjCGH86CBihnzei3LYEf4ma5kZqlkxTO
m2qMIV8cJFb/UrTQ55FoVgi29pO3qeeuJe0A+5Xe1n+v6EwhlXQYPmTIYGhCBXzJ
ZRQldLeN/On+wT8rSj/3pxBJw10b/R1ZyBg5rllPwu+7UP+GE5JrESiav+89M+F0
wsuo8+U4elKhl5htN1TIPedJGYhagd77IP/3y8W7yb4iKx7RSkSY1sNEd1foKiHc
oUbHU32RHLNFuotLET10IWzcZB5v5IASpclklcsbycvEVaMX0ioa0L5s00M5jD19
bm71AffBZbNdIPoh5iUis5EK9AbKDQ54ytFYCbWQ4imWXo0fb3mPAttoRYK1GjCm
uRkOTxf/qW3xvePh2v0DoOyg9dfo3kCeTHdvgHiTTlvCNAtd+hgj+rfaZD9ivcR+
HtgnTw/lAVliLds1kwPh3vbZywKHGa4IKs7uPsglp+xlzUZ8/AKNI3otGxKCJT1G
sLp87wVa7I0rnowp3tmkWV9og6C9Uo3bsb2mPj+uAovP78dpNX9p6FOQUeTbPJfj
jJl0/6d0AZTjFG+CPADtkK6f3n2Hop1iT+iLAjS+UZ9zl7BAlPPdff3Y2DZoJA82
2rNJyyJjcK0S3YcZFWlR1OjWWZoDRQjmIx69gp6KQAPr/+MSp0aQexWSEQHHCW3X
SrDj1ZBHGpguW7nm/xEBc64cDdlmTOn23MOLQfSUlgYaESgcbHqyhC7L5yIjqEtL
oC+jznoUdk26K0NozW+ZJZXuAkk1AxAvlTsT78eb13xi2jJ519FnYD1X6Yylgdda
47Zbf9o52KNGgPUZVlKULvIrO23L54p7iYrJdEN2vKPNrnadBJEhVCwe5K9l8qeb
MB3oEuG7v7OLLlMRN6xqrw9VnlEUmC57OeyiYdVIC/kqh5KNZmW7kWoeXIKhKEMQ
YLg0v0TDwOQLPLNMPQObZZ2keVEpEY2vwkwR2B7WiIyY7Sv4f5TDm98HAkl5Zumd
paGJXKEIhkcZr9A7Cc/F6M2VU9oJaaXprLSH+ontnY4dr5NJSQI4LzWI7p17JOM7
A+dJg0Wb0hbZXNOStRUxcKiG4UWg5qvAw415o1CKsDoGu+iuSPsHI9+jgCFVsP7N
M5KrLaMZ8yNNrtAaDE07fqs+fXyn/CIpkYWwnfUca7gO0gKHpFXlmpKDQkk/mzV/
j4QEuB1e7gZXoCYf5k5JH6rXZ+RJmt+iWmoIHYHYfc0rNw5EUaa0GIqJgNSyJzNv
jTr2TschOkkufgvPbImIPpkyfkZ2Da/HnPnklRb7lujpW67kv9Fws7oQFSlp05Dg
hQNEr7jeuiV07IafKDYv9KaieXZHikTLs6znuROva9iPEEWq9v5st9RW5vSdrQLW
bMJHzBKzfiR/bmSoJu5DJRH9msTLtcapXajsBhqE6NC57cg3J6BuSC+rZxLUzOuV
3qxKUiQzDPFWyKepQpvjJhLMiFQ7X4hKj6k999EVVlwO/dK2c5PSMdO+5lUJ/DQc
8tANWmHZh4V/GyfzIudNluXJ5lZA8kmbS+XA8gl/ut2z1sS1xYHGKpV+GQNC+W6l
Ke6b+y74SXzaMHsK2Jc8wgaFf1zDKuJVcNjhl7AxWUOVFBX1EMxfCtGNSS9WV7xl
bcn11dHeAZdFOFfSxdLFJNk+boKsPaVji7uZs1x8hm0hWP/V3X8P9DLR8UHFAJ0u
RGqeF1Yoh+kRRiGdd69HylurvEqMX+LZNolJB2pgtRDBmfErfjwB2n5PCMdODzn+
XmUik8/AGglp7187NKfpwvlzFiYSGCP7VVBllTThqe55yKqO+HUBapmoezNSvowZ
JD8WyzRXe2bc5I1Tgzs8y4H4/d2mLnwbYBvZ6CSYoJETM+1MCu3rs/BiohnbbIfc
wml86rYCAvChAwYHuHU85/n3AzTfkC6R1nO1eU857mpfRZVIdxtYO03acrGYJex5
AUmsN8v9r9+vsdHcP9YPJk9vrrXlzInbK4oXzi2Ljw4C6ROOvUZn23p921oUj6S6
30F/26MctZ3ZIEIPykiMvTqBDHeJuHkCjly7wZdiqDbpHoNvWIbqO14B6F7nnC8K
r9dUjaM1bAAxwidjDFttBEJNyPIJ9p7Ckfms1nFM4h/RAFDMIWxgwHEJ1jLX5Y7W
czqpVLdVExX5y4xdcpdky6diUqpMuUCeqJGeumuiZifBJXsOSj2LZWx+vcXhRfMw
jkG02zRyQu89IRx3gSK7gDcWkSYIitev2VpT8Z3QiiO/OsYI+8Rf4fi2wKyQwa1Y
Y8BeTI2u8K47t8/S992f55b8I/x2j8/d8vrH2d5LvYXuVUnYWxH7I0n6YdVorNhv
B7TITEf8JYlJL0Qik+wUpwCsLa1jzdBIlZqSgJjEIY8a4V8lxX3B61RpdUsEWrNe
9SQUqPPhRvhbUs7h/fPBtffvmqsS7LHu7SzvuwXwTM4zLB3mfTxa0vtwpoMgddk0
LpdqRN8ymTHsN1YWkkKNzqIgm9AO6zpieJcZdZj5LqVFgM/avYhcnO6dHSQ9tHQd
anCefdyXKon3aqLEMsLIgNVpikf8DHIPPpe4vSBct5lZ4dwRPnS0FLlibBVGOXlY
HZxYnz6aXwpIhL9WAJnSFv+f3D7hcoihg9J+3XPH774pzAqpB2NfbnLgu+tvxiNv
sO1xq2G6dzhjFJWm9GGolJ9vnRP/Pe7Ang01iGVtL+X1RnKJHwxahnjB9/hNcGYM
JO+bHqZDkDigbtephcVuNsWIMzR5QXGRFBmfS3oxi33MXwofQ9ryNicanTFrQSmC
QPTg4FXcekOC8D/6D8YzFKD0PNtwgzTaJq+xtsGO3Yb6MpfW259XrmZPAX75aZ1L
vqqbC17/d8zpUxZ4j/NzvVNHNPESkTGe030rvoorXj8VVQfTW7cMvzUPch2o4Z2Y
WS84BeQajolUSiOXAqHwdEi2r6oos4hUins2vxKwG/FmHa6w7AfQlbf7/W4kvuCy
LKO4i9mY+2ri1R875T9VrRuc6cYRUUq4BL7al2YbjJ1ILLCNQT49eM1OfbUbYfAG
8QIzpT3bI99+eL8xWPjtw4KUruwKCSHP8MfDV8zdwEp3KizvamrK2P+ooVLaFAKo
34pDwhWcipVUGqnOcmRSMsrY+1pXWyj7PZwx8rrLcuG/ya/y7BKCGoTeKRLckoVW
9s9xl03ldDiqXu8Cz67QcO9dOjNSky9xf711Q0ItRSRNlT0LvDZmzcpk/TqbRElj
g0LgB97H3rjntb/UXFpr8KWOfEm9a7jcHOD0QaEU2wuCz85wnV5e88M/vOZY8JU9
GU+ocIqBUPuhspeE/CEkjEXWqpvK/N9/kp/HIK2FywtewOsLP0cpcjG6fkdknxX2
b3QuGYWybtHl1cytWQ3d/gTN3rVl+0PMKOlG3c7yC2eu197FM59QmWq/r5BwbM5L
LR7lVQoZLW9/Dreltfy7ugQbbRjaDJcr3hZGPZIlPymHfFk5bkQNvGv7CyPQOyOi
QGJoL8MF0p/6cAYQ0KTt48Hv6tlanu5mqUx+Iz9XiRvBDe5KadBmeMoIJv9HRhPg
k7R1iZRoof7Xcd9GRyzkad0oVyUBzZIgR7kxe0KTHpsoxgg5X/rVBEY0M4RBn2us
xo8Itli76yWUySl9zA9wWA5o2Hr7ZlAU6bxvohBjY1XfUfkNPLRkNnXChP5s2/EW
AwY/vMydyRpPec1vi+1wyqefEhChaiA5W9ys2oqedKkqCf2beIxTalrtaNd0NAZq
wMdlBg0Hkbskp4jGrBJIjR7CBfbvbd3NvRvBCF0K+Xqm3LbOPgC2tfOqQxwgKQ0P
gEjti36T/Rn40z1bARwePiRgIQ/gYhhK9xP6zAHF51ufAQcHe2RV//ai4tTgVBKW
Hrv/CDoKti9lmjsZ2pj01wtch8R6WLK//S7QCoWuq4p0nBrxwC70OKqb1HVFjc1W
qrKzWx5ZNdacj2goH6g+TSeFKroHYJaQrIcsIW8Z/7qX/FjXV4lzyJwuBkzTVDwu
5npCOVwes3d5ltIsGP+J7B39lb2s8tVdOaav3uxKGfnyMqdNPKZ0KgVxCrhiW4Uj
dDO7C1CN2oCVFqNnZHM6DdIjsbu9zcw7KxggNs5BACIqTHyHXQi7CCQJxGzLLW9u
TSEtVx6RYhd3k4NSBhwvDP0DlhUN7Np1v4QrnlIudNcGusbWq68vLDBlg8B6wiI6
hiBvCn9/fJVWCWLe1jsKLMTEUZsX6fWRVz5oaOva65ojtkadghrvgoXwOyrP0V+G
IjWFz+pa6IfXc3412Aks0ncCfdeC/ZfcEA1vz32uN+n8XSAYIczOn3uJdg1++Gte
W+5uMMLFBatgAY/qOmWYVawW+7/X8Ck7WlvC+sVu8Cps0Y3u2s9o/7IB3SwSzqsy
7/w0Sk1W1X0WsQ9e3IP0YcooJy4a9ztOj8iKTkzkekEvY10FIs3jHbwHJkmwj36R
YaQASWxKhgdDwXPzb8Ry5x1y0UiQS+LCOBVyylIPheS5DjhO8AT3lo8+85S9EVTe
Pm/yFprEjOMWL3Ih/C2hAqKCfmLlkGSDEnpOMGqiJ9SYrubUWq1BhVilq2+YQpLx
tnsDpvt1ZW+YCgfwFIUrnLRFLb43roieL9iXTowCVjDARUFKW8ueE6agCfeFO7nj
yyUytElZw9eabIfuw6d1FkjsoQetX6o/j03mwJlrMdoEn6Oih31Zjl0yjPZ591mV
f/sOL8qPxOxH8AD0tcuPph17aJQoAF5hT5W6leQHvLTBCQLtZkqfm+8RlnFnxuUg
uxPenPt8ilhiqSLY0a0955Ab1PPsH4sywGCOvjZYQy5Px/rji2F3b+y0wL9TwUbv
PR/IIelFjg8i3nO01/l+VI35oZ0LG/D5nWxJo99ZzK1IY4kQDilez9vxGltWooVP
UtMGES51alZ/6gRuEkFY+imRyWGv0ESn7Nb0OGCkjoI9C1bHzm11gGfQdxnxAA3y
eeqSF5KquaqvYqSZq1oakLjVW2QrzB6IOhRHPjDw8juicdSfiU616sFZdsMMAUVq
Ky82I8JSx241nZOCKstRQtuwNW+laM4DSF/DRY6s6hG/MgOUyJUS94Kd/Kg0GcEz
xM9d0Jj3Fh4cALuMGcDBq7Rv6BFHGTjc40YV4HfKQJFhPe5LK+61fNY3jN5D1NAX
Gs5ihSvfrd8PGjPPhd6Ix6ZvGXgF8oSFLnysJWnek3h8j5ICABr5+RVioKMRX5Pt
TFi346NETOO/PqIFXAttpVr5eY9tfcQqimQTuIsdu04G2zZ8PYKjd21UHOYls8gB
fcjnQ+p5Fpl236zg+aiP+Bv2oWrKlJTK6TauoxA+4VcVtpLjku7xN2hJvncJrCfV
R37WdCg8T3ULRjEDBRE3zq/6mNjTva7edqL4bE+1zMJNNZyKDRWjRwrbHc6B34A3
bV/MOS/clTNyxPXEYlyab80fH6EM9+Kg2Sj4XLSoU3OJlofGR1TFdNUrBvc4k3JD
/LtOU5bORBTkkjJp3qmm6fZqZ1b0nfNqFe94IF4Jpl49LpoMQLw8hwOTj3dHVd4A
9ZS6V8YLhnq7fWO0A8G9/gvAyYyH4X57n8L6j19906Yq0kvU0a4MjlAoHHp9A8H+
MGQqZzlW0hFUXGdQ/g6vD8Dd2a2rDeF4FNNT4/Wss1wayiSZSvsCGQmAnU+OWW45
+e1TmrtDFWkAq0Jz7TRHC3BSC2ohdtvngU5B7OWe5uznIx2Pa9IU2e3/eealnHuq
ymrKHLkRmXMUb5kCvSZoVa76eEURwrZSduPaCBRmopn1lkq9G4NfWVTdCmFpFHjC
CnPzUXKuw/oUlJ6dfM2HOIJ7LjFOvuXkIqr57WwXWx4Scw4ECxzLiNiG6NGzV7cT
fTJBYQE5GAi1lCE9ZghGkokbINs9cJ/AjY4q9uPF5vObE6zt3L0ATMF3ZqK+CFa+
2HM9ZFlScVpyeEsZnCsaAUVV0dhq+P3A/7pjtcrbaO0e/QrJPOSMB9Mh74UOyTv+
m2Fhqt/wU0nZ69NGgGXvovtKaKmp6WdjELGVdtC0JBgt1e2e6CDcRvPe7dhLqbFb
6UAhg+cK2TlHP4td7z7inKv5F+yURMPWL7b0ftuImu6zKEF+AnwaisdFq6QThbuE
5BUjpestEb1JbuWfU/NIgHkYkgpzKuk16+84HxqHOpsQaBCxr2Dvqr+8F1TGKp+p
uqW14ngbLag45DzpTGjVJRK4l/cb/dvSk/YDE5e86stHQNLGWTtwD2GlOCNem3if
ZjwEk8Q8aUy+tCUzY8MNegVL/Ud3l8Do5AoVEUJ+0bK/XvNjMNM34eFOl+wsfCAG
j+nmXdtf6hnyE7R1LCqfZ9mvQRNUaM/Wr0sKSjF16kDAnIx/x0TrW0/uluB/7JK5
14MG6F5EtwPb1iN2IWdQxkM39K19b+v8d4bHiHMZY9WPFxoQLvUiUbeEWyCHVrYx
ujvlLhaXt5UXB75nXFlOOVRDuXXbJDAEXnHRmRMDcJPsOYLYlPwy7cQtJmFNw9+J
b+ASYbY9dBaPatYsRlFBMrEAuLURMpS7hpmVzjtHPB1k5O17sNn+teJuqedhmyGC
T5QJiPy1AQUObrmJrsLq0V0WS+HOhQfpfi5LJRhO0lDzUz2gvtvretKi74zrl5Gn
zpZPC5wqKaHAwEuAVVhR4dt9m31jHDB9VL8M2ts8Eu3spVaQPzYWKdCIk35shX16
qZZ/fUbl0LKcYEvnCVrDlv1hj2SoAOdWnI9c7L9suNaZA+mDsPoFEQeON99HCh5s
I9OsNRYTzmrd6OGInEqOy7X5aq/+i/bCHXIRj5RgVThb8DwpKABJI3URTpLYpSpT
tfkipJ+rGaOohlIQPPoGqBgUAxUuIZJkmdz5qepRN7FTmBIxEPY65TnJuAOGDWTY
YNHWaUnc+CzNwiSWp4ZAa+Rjt7huSKsxKpUbMIT9aB6zjS7ZohS2Q1ggmhhnyoHz
CpoW1XL+JJeV4GQJ+ZItVIunHhEfZW5gzuP0+78aLVK1HMnq3RfJU0RxhDxBt/wu
EagvQqAym1jhNtXQsLGzZ4OGBPKpGFdYUOou92yjMUpIouvby16njPuLMRQrX/TW
/lvpI+Iyw7Op5r47WumeBW7bIiWbyXMvVsv42GrSWqdBUSum/REnnpHb6hUP7g6Q
p9deo6szdb8o8D/zoItOgcc+kboStaMg7xwAZ8YZPCczjFb7qcN0bmA/FOFy69W9
N88w1KEOrLFQWLqt+U0Ab2+/6bE6YVWYoiRIKpYvBm0gGf4B+nOdVqmoamWor41O
jiRxEsbLMRJ5wOrNKkhXkYadQZQn7kcWbjLKpYID4qyOeZxd+n5B0nKeVvDsQ98x
i4xfMIFM7REpWokEn+HiBqjP3wCWg2s8aWWJtPf6bLsiNhQzXXkuxhOzC6c+fcEr
SBuYBVSnrnX0+t4K0bPc8XRUhikylUBqNIewLTwectzJ41vj+bDnV8EdCKa0xzF4
BEy1xdMdFVFVK2P+gIYOao7XYg2iiDgHM7nfBfYCTN1/fCcjqRF/lc9Jcy9/Ka51
+jtvQEltIMX+8wdEnKnmB+895nxQzf9SZrY18W6ZzOxnFFBz7T7FXWDIa5V7Klvf
pRuBLIRdh4SHpb/DD+OiGvEsDo6bT6lrqg0I7Px/MaeOYLsnQClowVafmeZxXriS
x8UVPl1zUAiHkQTAxdlJkBdcN4EzKwJhDGqZW4bBK1dN1icbVvsz49xLVimLvKEn
3+2lZPqjt01HyWQHhrC7Y7GJlii2lacDV8I1Wenp/VZQLZFwyhQ4CUX10UKQFSh/
gbUyl17vlhTyGj7x2QaVar5U7uqHJLChCUMvczmFeshFgOr6pClT29JL9Nx1iz8E
AnogzeMFU1324rBjBYCskkrrLcmJov54PA6Pp/pS1NbaislL5zc51+Q3KPYWdf3+
2IUURKeCN15wgXeZz7wzPAITUd2JvDlClqJTkm4+08imL17uG1Z6gEmYhOFFPCyD
OvlculPsuTh9D3v0pPd90PRW0dZBhcHEG/fKqbeyzqTtO4KTpQUvkihV5qCBZTjn
ws7XdUyojXOvQCYeG1oZfByV2Jif1iwzT7Z4Mmfw1r0Zpei3dzCEmVIWDNNajXFt
YgfhXir8AptBcoOHkoHS+siZ8vLS08sxXyQDoQwi/PB+4D/bVPK1r/pJtLlVvrQv
CBMVhu88rHs49r2cGxQLbAEKlTlwoSSRbyCbxNtPzygYeC4G8tO9q8+F9rw7SyVl
dwWcSRyiilT3PNgvrT7nOnhJ1an8cUDOc1k7N2OMnUbbcdS4A0bMW9+oqMBfNa1k
UQrFPmJnarLd7xCSpKUbaPNoQwRe7NmI/gCmaqF7x3uq3t7zSpWjVqz3AI2FAjeo
DfZNvlyBQoQ4CymNwZBOF+pjNrDgfK35Z/ts2Nz5hJ/AmzWT/J+ZrgmZGk7VDxJZ
/qWVuB6hoduP5poUkGykj3wEsgGUQs+zC+4WBzLXwv9OdaulD3dXTSyxzNPZxNRQ
lvKyr5oSrkkV1y5yXYcRPTZ3u30QmeOWXPAAcu7YLlNCSTgBC3jjg/vVYVa4s70m
YsyVD0VEnxPnT851/eoBPSqklA2+mDGXhnp7DimtaOiJrx+a9/x9jU8ahB9UZqmx
osjBfTKY01n9PSsL0KQ09v4S9dZApqdBEc3ge8C8WyKi9Cm2uNrTyqu/+QZUqw1s
3iY5E/dWbAU43hB0N3M+nLZtP9wM17WnxBATVC+SKmK9GnhLz6Q9wWtRxKt1f+UW
78JtM6sXr6s91QAgCmyd7IdamlgQKVs/lof8Yk7gnM+KN+DejI+rvf4CmYE0rOhp
QrE3wP9HuITmuAgDZDTIyr9SmfW/WlWZKr87Q+f071u4oP+QJm84sasLWWTZJqmo
TN9+mK1SvR4rTYkr6sCScxy1UwkCHjpdVmzMSgzDn5A8LqgCo2/Ca2f97OKueVM7
dxs7VzH77oKMV/ew9U1ew88I4i+OGv4ugKrQ3Og/j5nkLbht92zlL2E0dYhmlotM
9H9RRcVaz4S7FfI+zXW0e638V+Nt3zPK2To7pJ2TfsKrICRdyuEtXMeeaNRZlk9n
bKO/if/MYO6aaOyp1Sf76+3PAMaQOXqchdaHB7rCMBFN/fw2/3UktwztCxzxS3vv
WfR5IrK35BmmCzA+nmOrvBzE5WfWuY6JVuQLL1B2YGCYsE3b3AVsZ3UwRB0UMZoH
8E0ERWIwBe2XylOqvqDJI7IZQg8pXSR6CZo52TIQpMDrN4nI0ns2umGG0UStQJAp
RIXnjIK+k3p1KnJcey4aDrTeRGwSSyTh+YYEhFX1SwncGl0zjnwLo++sdsJCxNal
B3PX2sd8rvnq+mFaqn1p6ROWNjAWYuPjsXb+pNCIoKDQ4T1kp6njEM/4r+ojYQGu
xdn83m7BkiLLoTOxCk8WvorSPSjKsqTN/QmWJzR5L/ahYTkxyhlYaBsClQgkqlZi
YsG+ChHKS/9VgivsYGpXskb2EP9FRW5bpE5+I4cszMBZXBBGYSuA8ZpNsl6Q+rKI
LATcYXApYschXiBc2TFrX2OZnMf25oiOHzzhCc0XbqiSaEfs1EP47SVZx3fOwtTT
nJhKT330emKODX3q2E8Yuw79qep6FEDULBin3FjFTH6K+TaQ2jkDaXCHtWEQWjPe
4fAhiIsvX7FSsmBfFep9ZQQkTZovU7MJcUQZt+580cFa1I4edRyT6mM30XnpkstM
NGQAOPJV/0biEVppRWdRf6QJtZGbnhhSCxuQnLhijB7a7b/LCmfyLq5W+4I3qNZe
2BxaBXGfkKwLgwnh3TBg4MDg4eBOE9XbwDO3QqiE+q8zsO3UOkkz7CKKJvAnN7qL
dVm65ASuTHUHqqafdqaAIcZdLQ/ak+IPaSNnMvl6ffchuZ0rPYww9hP/N8/8780n
3YqisYs25r/gWzPeOLG5ZVa+LqS8sJXSbO6F6iTWqjF+qdXWEVZf3qHxuToZolxe
KGOIYymEekZ9ipQOdpjZLDGuCRf7fWG8sVN+xOn6AbPih5T3ifaP8DrWvKRF8bpI
c4cv2RT0Vrtkw+S2Km/0jVxAqd1MMJb5EnDNRzfcR/kyyAstPf75usns+U30qp6z
khYtqiKmHlXuYIORzbpYpC7pZuyhiZy80DjvVextS6XkT2W1TrJrbYJACZXBSDAH
MwLWKPxDXoNzOqfiQQxX5H26T8PEfRIRzMEyo4maeVzvhFHEwbuiZrqesG3OwYM4
/5BZtHE0XWBYyT5TB7hI6LHPc4AY88EjZ3dbIdq29JOfF4RbHFYEn00CrYYoD6HU
TqT/mNEj19PVrXtOQSPFkgIGaX3s6HT7J4vi/zRteY1/gkXsUuCBcA/wW1wuCm1W
ABWBypvqQfmI8DQbVmu0fL7moP522kJzQtzuG6vaj+FwazBoXit/pDNmLtd8VQ3h
rFqDpE8p58DTm7V4/r6AJVcLbbrEvddm5f3IHe4EKgMawsW6yU8XtcLQ+suAVFC9
le51zDTEj7EYQbrdWXTdSsYHbEqT6ifiul97NYPZL6R0D+CCIKp4l0z67QLqlC0j
zeVT28WcomQrjol8lkAv+e8gEGDqz9q/BBTtxdwcWsW985CG9MJGz89aWSlhX/FJ
DSdFJOtxbhf5T5l8hO3K51rABEn1UeVEePWMuuyR8f53COsgTBhhhcOdX7+DkzCI
5WWT5Wz5pjp+/8Hz60AisBtcrVrYOrEotT0Kx0FQ6YTm0cZvS94CEMLVRoodJu9F
kSS6TaHeq9JY+GjH7MP1AM78+MP9+8pMiyeS1TwmTZBvWmGzzy0I5JteHPa90SXa
f+JmqWMD1p0QCy9HZ69ysAL9OSWWiWFOgbzCtMkGZsrUNJosoyaMcT1OrUEEreU8
uTfM3VmePJmYHaDudpMjD1EeeZT5y9ssQOED7KjfkgQoY78MVw38+JlMpgXZt2uF
tnyfLSSfCRxSdzMCv8/cJqT1hGI4LIrb9ys4zwJBFbn46bBQc5KI8e20mfT85RLb
KRyKJxwZinkEVu7p38PZ/0qMZ/LgI2UlZ0TCv4W7GxIBnL7tJq8bYeOATcThblH1
JSkCxFxfwV4lwOJ9qS8AbMhSHZ3R83KQJq1UY9cDG4o+qSWOOV91tDupj73XlB1Q
BL3cVJq7Yb0li9bbI/K5jwKPRo8Sd5D3HzjceF/nYuh/Ky3KjrW7mz697SEuOcAX
HNCetMFQRbGScZ5U02elvOCnLLu0GjgcvZfUn/icjxDkTIPtVH3K8Z8Y7cTumACg
ERs2QU6RTVL+8RB/wTODyJCQMpUPo005KQFC+HJTjpoR8nXijy4+G9j3t8Xg/SwY
jqv0j61n6kLcwAjUfh0NRJlnKeGuNcDEawO2A21N3NBY1JT376VlfSDpoLBBjZvQ
ujROt2FfVmpElZfJM9P0sb4V4H7NUzEbJRUDCHlYS9Cn83Dr+589xZ7hBUkQx21O
EBNW8LaU/dcy1gNEkIgf4mgn9ngW9JPZngg5OmWdQDLbY6KfsnUFxNNvuk6KFPKl
TvsBl6n7PMdvogOLWIQw1XEFsIbleHlSx3w25pDepBOBWmrpRUV6axx9gaJt2qPN
Ek6eDy0ZXpuxHCbY1m8AAg2wDx3G5+0I/VkMnmSh+7zr55dkN267dZ+rQDDDdM0K
p1jCOuP3NGL/JhNwbmNWjwVupayn8f7jg5HKWXqeig27P1KAshgWPQyOPWRvgF6/
irz62EEM+/nqdgA6q0bRwcJOFM5BNgI8nDE9rE7FRY0+6MS9Bn6olRAjx3AIcet5
GXIftRMHJW+EwvZ4IfafuuJBqE2QAk9u4ExbS/L3eJCl3y+Bcdbg/poBP4n5mL08
4HaaaUFusLYwQWLyITp2Kcj8IBOKVaXb4yIk/rhoJJxsGXE6eHR9H+5/8oT5QMjd
pljEmhJAEa2nNztTKvunbwqaCEY8c+eOJplaXVDuEa+0CZ79A0AQSBGXk52f7UFq
i5loii+2G0uN0t7xooGw19kXSP3QwYyZOJU+VCx30o/ficM3yqVKmeXtatyNouia
pZ+++FUqPIrZl98YJjAsR/daWvSfgFfxM+zBuw8jqeiQRP2DEZXasfvTf3YV0+2m
8GBcyku83+r+g9n01bbn0Zq4Uu1PlxAVRzND0XRVGwHzg+i50JU3YhY5+FoBNjaj
kkE4Tva4RAiczXkjUt+58CNvkKnDk9S2dv0z4SoBFOZxHD4GgoDM7CK3ly7y9nn8
Tr9vNpMx2KM/uje2nQeM8WHYivGZ8TwZTFLwO91KGgTjdjWDhDnyIaw+7enK5VD+
ElAx85a7GD5B6Os6FDysRwMp4E4tfhQLmc5dC3PosYyf2KRlUKfaIujS129/379p
FItDvu3dzqA3jc2zHlGUOXpdtpoAD42vOakiZ9RNWakb26H6jClPMbrYYYgPlh8L
oNj81d5gHE1sWbrVzqPCxblNn/K96KJuhuQwEeptZYD+JlK1hb+6CbX0lStSuReN
FFOWJUyqV70snsEpRCxv9srPDd3g0JyEFZfUfslqOyfqi419UmgDviP+kqtrf750
2G6Gu1+XyfIbmmtt6cokKluLDKHg4WAosg7eeEF6pX67jCTsfnZh2Zt8j7hkVo5W
5cy7jFZOI6OXge8AYFJeihgX7vksbxwlyiYi3TezZ3hYZTeIfgIALmOblAQqNNT0
aBAOQHmjg/C93eDHXwxK+dWzVw+ehdJC08k3ia6SAN6a7O8ciuTfrGOv87+sXysj
hABt+wo9+XiXt/gSTavOc/Ki4/9NbhtSXFtV/4zzUXs633SdmCnoRFrX3Qn0nzUW
M3MUSC2i0a/QrOYRGkV5Ay6/SavZkMyo1UsVuVCNBvSPF5wY8bHZRsQmFs3KpDBk
62/TQSUlVnhZvfGcocs4T6vM4+PkIBHQgG1hlwN1UaWcUcsXjo/6p7va5RNUaeJB
fhoH8+sFi9W8fDlao5rgwds3IgQAtCdsgPcv1I456gQDxV17Inv6A8OGLv4Sxchs
bDNg++gzWkIw9hLx2aPAL+TLeqMLve+O/cuxpuoVA1tuqi7amafPMZ2cvatGDpM/
eAUgc4UyXgMfqzQY8OAUemnNyHMCVjf6NijXm4Dj5PBPvjaKm0uvroluxdIPlv6N
yHKpY8kgnUQ1krSN/HXPsAiRb0+xxwYpuX+0p75YcDbyGUk7yecc0r5Fs7+tde8a
V1BvOP8OJqt922kthuWDmr4th0cT/qupjHbqE/QWYoCMD2EwOFxuIwxyh4hNOC2M
fY1drd//dWrfRwYcorbEXkBEAmHwYcDrqTeP4ttGNF6N+4x9q+NfNy7ffIqO7T/z
O+ljFx+Wu3nzlrmzRpCHIp8RiBO5f1sWuJk3d9ESHcNxYgH13yX/JwZAJiG2btrr
sarGsbc4T6jJ0SxtgJ5S1h6IOyHOhVV+XGknVtJ+mad1IPeK1eY17Fjy78lJZepl
XjT/nM1NkuK8c5f8GyfFa5dhDMWLkwKaBCpAYam0yH6y8QjZI6QxYK6MLK3kw9uq
sgdpESjheiPFejmAepUnmjGVC94W9jspPaYo0d4xIlb1W+NVSDWH7wU4ELRk3jpB
Lu8EngcHXH/ILMa0D19kOOJK9RzLsww3aQ9KbfRgLe5S5coX+aQ/n12l8ldH2fgt
u+l4hAupi4rUc7/D5tHhiZPmhTYa4pkPRp6BUA3wGNW5jufN4Gm3gnqoD71Eq8kb
y4BQoIYoas9JxJ9VnOXlsZE/m2RseJ9RYTFoT/iJz8JnV/YReRL2LS+Aeb3QUOT1
HPBtREtDeGLIFWcfbaslh1pFmko8luVtrECSVADbBjMADb3h8h9jV7SaH5ylCOHT
mYFiF4wcgc4nGzI62gVNpsNkvGyDhhe7JcpRHPbr7nVz4i8VjW6NUEgGZstzC8gr
Q90Z6S6+Ir3Db82TXDXFBaWULfu8IcZgyWzVNrnH6QX5Uekbzwa9mtfl1/7kHHmp
rbG7L1sg/cqHnT/1WdVHmQhUitDlbUgTQNqmE5qeGOky8dNG0Amhk0gbzW/A7ubL
Tzd1Z7orYDYKN/bDcYfnEWRScpCzZIYANOxwsuoU1cmAmpR/4SxTiEYyxoXGeGRc
6JP4GJvPnzgQGK+qsgff3TeGRh9ddgGTPmyB1pZ+NxsdKysv49KoYZZW+3VfTS27
NuZLQ8KRQiiJAfvpcizeT8gRfYxbC5U3P8j+XL1qhO90bxISi8RH7ymRSiCQi0Pt
bSWY2KCE9AZBgu+tQfH0kBKSKb4fZZLxi0M1RIjHSi1fQ7Uew0jWo878ZnJiIu0G
4qgzzeCLQHW+puKEv/UCRIFqr3mo+vdr5XHHmGvCXionAF9DW7zGumr2BzUZO6In
hHT0f/QCoiCBI5OTG4/1VJcTTn+e7huHo+xhwJS2WyjipUt7oX9lVj2IaQ1wOiky
8zDEf0ft2UjXfXRmL4XPvp5oC8qD0kZwBRJqvRIyanBIYAZ4cFZPMPCyveJ15NhQ
8kXgneJ066pnh4gnZW2awUyB86UwSEG1jmuuzVBMzlG3YSYbzFFpos6wQnSeU6ke
rK7bwbZ1I2gA8V77UcGmYHEM1hdmisKD5LctBjeHX//By8GSbuMB6QJ8VCrPyoQm
nSQjTzQY6Yt6KhEsU++k8etv6Maj9gt1c+1t7yKrn+ARIYz5DzlCy3K3fHnOYXQA
V0zUuxGhoO/a93K+QjeqSzr1uJntlojI7G8pMFm8gtdQLRn7Y++jsDxglE7+DDXH
/8ktWo+z26HKJHShfs4dQ3/fynDjqGpn3/L2z6oaI0eHUSQyZ+XiePMzPAQpc/Yd
o22jwVbx/3ef+ZPlTv3JQSX3XmeTHbJ2yKdN9hJoi6vSEv6RAYOwkVffgOe7n7qD
f2S5LVrsCtGmow+vayA/vLBY1ZdKxG1SQKcfcgQNMdh+oT3gqnFyCb5uZa4Qn3KM
vBGraGLbH70cCoiKdi1Z05he2R1N8IscPzC72ckYrwoVyvHQUazHWxBARc6u6eMW
IwS6xlPhlNJAe71liKJTiTTVjAcHUvDqGDhAL2sMP7ZRJNgQUZi+sj8gHXyT68G7
YYgqpCCOnPZrrN9xnEYIKuAlIGefqrZEx2XoE3K67u7Jo/hhCXHd50kJ76fFHb9W
xnH326OAy0nxOMfndFh3xttVWhdmy03wZ/NVXhUmwgWbFhujjua8ZJxXhp65686a
DUqBxVrKqWNZ8SiMk9W/2aBCF/Al4s6UnOc3xC78OBv7ynLkEpmsDlKEVTPJJjz4
qsExY1CIDRt7Vh+KqdqtfoojPHfaLyxiFjyx3/WEQwWWsB9NS77DYBN2NT3I9hrX
bURIP8T0OlNVaLhqmJ+XpBHPfrCrxok7ECzpjAgRqEytFghHR+timyEseZpxW5q7
3WoeQlDFgR+Vd1mx4KRGY0eioTFaqpdSYtVt0surNVq9pVR4Ad92MgXdbEJ8sxCU
gvhSyCXSBE/Doxh5ujWwqNd92IjeFcOBHhsVZgoC9vodQ9a4vOcjtGQ2u8VLHw5v
eB1mchcc+SMINntD5M49mb7d0XBgtaT22h15FIiUI179w49XBvCvHZ+L2ittxJCr
zJ9VBvobmHvhokQctK1/qHKfDvZdS7+b6EocTbE8IX/Na04jj6xjHMECs3q1wWuH
HhCKZI9BFgCAIdi3TdTogF5HM0iK6wgm/u/9KSh1clgli52/zGiRt7+7T4Newyx6
NZty8TqIlHACpNtKsAeoCWid4/x8uKy0fi+uf4zHhuhVgb/agyEPDzb2FRZy0+67
ZX9A5Qfoa5rfurodDqwFQlCLbym6yaCA5co3Z+62BkdPNeDS5wtWA+oqL5/tQQtT
UIYcda4iCxHbanTvxRagtLwYLboH1IC86W10uusgFNnzIqGfVPbZtp8gDV6OJHWU
4ocouOZn50sunySrPjWKypwGSO9V+LScyNnehrZ2pEczL3HSjTkCIg8eI3Itadmn
YaYq/ZeRfFY+kcp0wbFga9RddmwX8asOaI19Pe87AMnEkSmkkJFCLGxADplOVKlb
R8TWuTJrB2JIcVIhN+1IYAJC96twfYmcO04erC2ruSZKZm6hlqoRDVbE4za4qcp1
GFAfnfAFVbGxtnpWnVsblK9JUatUWPemZAcjmrzvVNVSSN09OlR/etINiqM4Oq+6
4qCDZf3lTv8RTjFqQYvMyWxVfjhQngmZvc1uofvWfNVaFSiqd8WMVDOAXpdPrvkA
hqF3uVjFBhuTv86JCSgy4E1wKjxMK1srVMYoCJ7lIeHr5yZ3RBBtVlVvGzTjY7sW
8VML9HqCl/dXWq08+XtkFdJZ3JJ/02kbELWakp1cU9SVn3KZYdyb0sD2LxBqyMBu
vLZNH8vSNOJwmtkhOiYNYWh9NOrQ74Dfudu4tFSpuxG5M6VKPuXWW6huAxs8YIak
wGRbPqPHFfgQygHBF9te14YeeUORz3sYF19mXHITrnOI1OiONxx8pm+8E8BCTZIR
eCkecUl5dyVrQJScztCCsr2P8qGuoRdiQl2mIHvwx3qS9kXD/+Ciab6pqw7T0P+n
JwFfFdXXZWche0cba4cmvwqi+riDjwsjsuI+GnKN698V81cDV+iYelrOUgXMx4o4
ZJ4cRMRWcEo10l2BEQNstZ9TTt4B2zF7xGD7Qz+aJRTCLlbtsTb1dFVHNDHhLOS4
ZE7L5zddoHc74Hg2xrB7xVBvG01Q2mTRhAlJUS/HIgGWkQrOddF/Xmo31RHJ18mF
9RGjwVBvetGVj0vJXVdoz+quaoNXro5JL5kPzRWZM1ahOZxjW4o3Ulddni2fEYmv
4z95g0pUz5rzzZPAUqLFTF37jumR/Ha3hDB7qQNzAOrxNao31gbYqj1q31z/FnEU
9P3Fh7BrQt8KC49+pNsEVBlAcUOZksllMoSgrhsXR2vCVVycu/PrKMcRvDzic9G7
wEP1PlHwiNejqnIzPEj1bkCi07GqlKu/QjzvDcFW0kovuwyvZjvhuuHYKn9aQW38
DKYPXKFv0pRxlGaImrJVJHIW/PjIcDHZIHlJdC022f+/8GqLv1SiSpaD8dr4JQNp
9gfGUWbw4gpRd6cW4PQ7u59XXOCt15i3sCp8XbcTZ14PVM3wtV3smCZZLAmOBWSa
6lpOrhmmxgJpEq+fUIYLY6lo7lpKq7bUhqlx5+50kini5eGtAQaMfVz+QD3kx5fZ
GZQ6FJrFe+iln1MF0N/mjvYcMJVcLUv99aXQyS7OpnyF4BagDrHplqXL8YJerOpN
6kCMgpYKBAWRuYvnuog/o0BKEdJ0jdlGUIqqXKHLHUV60nRzigMK+c0z1dbE1/+P
NH38alDz3Yj9HIVtsYJOXMLwbt5b/zBgFPJuovfrabVZ2L8hPQI7c8AJI9mxickY
PZXK08lHu6Ga0djIsqOpp+7/HS3IPhByK8iG3nEM9Xtmd0zVHK9pT4bGEosnQGtn
xpHkSY76UUyEMrp20zea8POp3o1iMG32JC96tWtCOyLDvILunDOERkC/0UmxX0XZ
AX8kWx7H09KsesNQlQXz+f9nMC6rE0XP51DWqQ5EbVfT6U6PWQFzjXSMxqN2aOVx
p4ATF1sxIdkZLGziKAwNJ13OorxbC/BdNnvti3xrw6ToCi/MLIXALeE3ydvC3GzO
bGHbTOy3LNkbfJyGIKgp6JHG9bHvnDFmetpaF7QLEgOL/mQPLFOBBijF0ZPB1rL5
as6ld9lQPeG9qlCFywQTnatcDTNW0FQEWkRX6LVL8EH1PEeWiZNwCaroOEuFHd//
+NG4WNZCNpnOStQwp2jOwaVJDJoE5BJWuAYU1R+traOUvmzqn8+CVOy7yMfBbqTM
KXPcg6CkMFi+wcU62rsEcRjZoag2WMJI8Qse3ZJeDfAQHko7bujclu4A33ESlMc/
Q8zQiVBpYggCdQVvqb+MI+CGvu2r0Ees8b+4g6X0lpajdFrLEEOdXGZ3Ig0An1+W
z6DjF/Jz0ldB5R7ygl+6LsfHt3INuJCVjkREkgGr8rCVqt2QVOj8cf8O6omDQ/+E
u7CIuO1fL7bgPsgFz3ldO0nbQfQJBffoDD8IL6tPXbatB9gnIsTm6bHepg1UaR6x
t32U+yD6rvfBeYcOcbTrE4BdXoV3HttJwnq5W/xvDnO3lvkurFVdnnmKlGVUz4+z
wv+apWq/i4h/dC4GXl3Frb8CUefZfmGlCi6m1Vp5afz2wwR+97FFGKewsfDvZDpu
6ZuXS0iHh4J8xrI61jRIXQAjJ4HrRtqORomKRzou6TQ0nnWN27paigX0KWz87wRQ
a5pN4a6bA4F3VrIt/9kmR3L+xUYAyg/xbspfR1pAqOvtezXJX4RP+b4rQ64yTD1R
EpYmTG30v2Ukar3N4VrRiLhMbhvTreNUtJNmaImbjRczpBLv2I8FqVfprwN4ojjV
vpDPpyU4sxl0CqpLi21ja8q4P5YQO16ZhM1bTr4o0pGvuTzcZ2vMxPfABXgnaXiE
v5hcbaOG1+MgWJvrmbg6CaJ79zS6GwtXswfJCOO0UbTT/2mfu3rJAo8fZ5H/u71Z
G3RyuzjRuz0ddETTnvBhjPRPCViH/uyCAKSyvi7qPLXEW2ezqkZG+IUTBi9EWtsM
purAF9NUe6V1+Mp2K6qc3jDKMUmORWfTjB7s2r7nvnuEUKvFTwzh+AKCdvh2gyfL
H4OQCXyBnTbZH+VKs/W7GwGUmVy3Ndkw+GKvD/sMKT8pD9/ReEEOPkCJFXCeTi+o
JcVy+a7juIl8ObMebTIsqtVbXsxkKkFtIrPEsX7DtRZG16/TEtjhGOoyJhO0dmd0
iVxMFnixDEphr5Phs1uFSeiaTmeaZ3TaGQnC3sWFYZvRUodT1PK3oW+/lfhDHXO3
X8WzQFkPlwnlrwsRntwbXBq58NiNVR3fu+JEkkv+iFSjOo7WAdYDbLI6h6xLFhbE
6hy/rS1tet2tWg9NyY5LyTTqxK1TGIz5cZvRze6mqaYdLLJmp7RF0vKkXHIGoi1q
cCOVk44+soArMwGUR9lXJCM/Rk+WYnEwo71lqvh44xNVde1KdBhByGq70zIEDwMj
nXN/L8I/g/NjvAp9SS3FLuOaKM4o5x1LbCiUJFCT6G4IDK2+s0dUYUBSxmmmaoLX
b6DJgtvT7aTJFARVbljavy3hRnUKwcYVSnYtCCh9GUAGtYH1At14F0wfCWV1yU1I
Z+AAHkqV9oAuK8/ePhB2yY1znWe2B/HWOGXo92JkFIthdCqF3+qkaaYXBVL0bXO5
+qmxOeY9+/AEhRYCk+mlp01HjF8UVUQtgCXq8UnrXqEL84a1KIlulvdYn+UbQmZJ
0JntAcYbSYSqeFjuidnSz6N+AjXO3bcRKmYbxvs7cjYGHCLNzIauySTMWIPQ2lfJ
QF8brXn9qCM4clgQq3zh0D1MJkZQhNbXnXhiLOui+sURzFqTOyknkfuWB0xvCgHG
RG2X2HYr3gH92mh6awt6ShKvJ6ttWdSdmDk//GO0c31L2Iofs5meNpae/o1P/bUt
40ioCvv/y9TTPPMfB5BF6yRzIcB35aQNbZoi4ivEX9Bxe0opeopm3isgQQK4yMmx
nChP2oEdX313ERiZlGVP2ROfX9/xuDAd7ePtbu1KHlfXXjgmuuXDaqddCtxGUFfg
ABHmjCX4G4n4hDjZ+6Ck9aaf0l56XlodwFhADcr8jFh23Jv0ty8zVgM4LS92BTpz
0hy4RCzB1amNuD25O2J22lwZXxTZZmKkrcC5XTPp1MI+WCqeYVJ59OhL81X/87ft
CKrc5lWMHVK3EvRsW26ePY8uv/iQY/Ci53xX6D5MaQn3xavJ2zcvUPH3FnHj3NNn
1XZGMczokXGqml9aJQxjvxyRue7qHmra1WtdpzGcXbykw4xINVmrlU0wnXtVBc28
XpJ47HHioAbViRNi2mL2g9dN3lrYDi6oiWd1+IXMGmYZ3j2A2InMSqwpDa+d652R
PyEdfYpucEVZEvTpgLtqOprH+Jd5JjTfqY8Qx+RG7dn7P3DRGvd11H68xVuxxRRV
R+07g4+Vz2iTbQ82t0WducgqZroMnZ8ZIpCDgJOJLCb5KT17k+LiMmYrOCtb4F2B
X1PvGkWXOvw0OagMKZL3zIdd0S6qGJ0WZ5kDvP5KY5K7Mp9yqpx9x7mIGBj0g0hO
s/b1U31eS9BjO/L7Ikt0bcVe3BBE9Ox/w+zxCV6XDxm29paSXVoW4gI9zazkDUyn
cDivfz28RoaUZIq4OpG7UM+uHzC8qAJdslgzSzjA3dKvxnuRWKB4Wh4RY5BYDiDl
ZYOL/4s9UV7WowQ8BtVlnkt3bZdgokE7wiXuvJdQLwrsHcofgXigcdZXSuNFm1Qw
q6yXeixgysVDWqYS2eHlc9lQmh2149Jz1bBAkIxIFQwcOV+MUPb8FbQ3XI8XCybc
bEc+WH6W3KouTTMJqWrndylal4aDMzawH8YQ6NKw+nj7Cs9lzupMGxDLQes1cu4C
f0A8eja2qOqrZmlAg5g5I1xtEZi/vhUoPRvpR+q48EdPITWosfoKDRBtPfXF8Kuk
zExXaz/0NZEJe2Xfd4WV1ncOWFakqpWDzF4rj3f9eNERV+QuPHHJRVLU70KjS8Gx
yyaR4Y5YbFDTu0WxyGcWkVROoLRl+YFoP+749t3TYBDT0hVQvjg4gVNsJZDv1W2L
2QD554v0lGs0+gbSETP4XTxUi6foROboe7RajCA0Yj+5kmiQSaSyhLwv4Xf3RyHd
73EwOgNCArP5rMg2gDu11GU/Z9sz7XY2tkOAwnLveZEsQYq0PsXkhL7dp0BCv1vS
xEgTZne9ai16snxDmWHB2VUvS1vMoF5+bNYF1X5dE8cbrG23fENP7l3tJOfKYv9i
9Xue/ouByldeZRKHxnFUC/gzndJ4N1L0EDAmjwtyRM8coCjcl/9SPy9B5Nyfsxfx
reAHXYQDw4OllbRbVXmJyq4ksK3uNcQO9i3QPiujQLBFOoQfilMICyGz+9Kxwf5H
unv8qcaAXgIBER18EX8wjY62FwKOciddspnxfeit3omd++RxvQWRJYN1XgMmoR7r
16CoPSH5kGzvBobk5eHmJ17jdGlsvnmiJbfvwyXmMh2vcPwB1rIHMCEcBA2elIhu
hSO/89fVsXveeRP1vR/1+t/0o0pBY/QXEnkAFBHmiRP2bJo5lndY5M9t6knh0nHJ
g6GgShX93so12/tLZFOBInh+09nbe/dlSBCde2T6g3lHXvaGN13TdYGu0nfixOjz
5D4nR3I4mk5OUc0eOL6yJoY4qKeRzimIzH5+fbh65G49iKnf5+8vceB+58t/cbKO
aAYn6SydYadROfehz7dyqgx0u4fKzcvh2b16iBA59KPTX8drynYy4KRPyENsHXOu
BDaPMHPWo/BgTeZsBN7bDap7y4Tj/5EWymUKKfy+SjBTjnHD0LmRtFyI/23w3eaZ
N9Ey/iHaeDs3kHEC6xc0zGn0Fsgh8NBV5/mbqcqwgmyuwIASyZYdWaoXR2f3Q0DZ
NwP7uiv/7G32O4uRCfdt/FNonSf3vD+TiS8tezgMRe7qWuicvL5FHbZrfQ03xd5S
rQdteT7aUekoN+jiVJX1Vd8vg4CRcdcPZLnbF6vxrUqKX3v8W5yKQYi1/1VR1Vee
Evcwcp8TShzYyRTL3ohTRGjkxi7PqBdeGHM+1i/NCVpMIRISw6t+x9lN8GafGEgo
9OxHx/bEvT0prEn5YtZFbQteElkAz8BkQaxTx/ovo8eIPKsWkStBzU3RrvbU8n6u
HwOqjBZAuT3l1CCbfRoQ+PQh21SKPxQZg2heW9K7N6v4S3MU2x8Bsyfb40kYVGsy
i1AyZr1R34bubOahelYnLfvNED0QE/vrahvjglvD0fsDHFS5yrzV0cG2M5DE/xlK
29Y6Mauls4KwIXiRQU55NlGXiERsdyMZqnbprROUG/0tJeg1nG7kTa4p4mh82l9Z
AsTCioKzZABydrnsU1192xC7JSTtGfrJBxVxjD1kSShZed14TOtypWuUQugzhcEE
2QUm9DrxjKMUd0xEit/FOXxZoPYAYqgd+RiWrnU/QJc2JeQZbJ1kRJURS496X7hj
vB4bQBg4hp3hpPtZWTKkJA30lkCTgRm79vg+xpzGsBl5ThVO3Adm6G2BErLSH86y
yqJ1GNLGimQkksDq0H/nunZ5pChezwYjpkm7KccvMJuJUGy+KFa+Bn+vQYz1GyWR
yFPnVY68o9ZBv7RcHKe0206BnGqe0CuZYGhLl+RlezHWFhdgnGaidqZQh9VHanUo
vEoC5aTVgFX8vnsNVjYvTpyyczNcAvX9vGV1cDbWhrbbvgYrMp4XgROc8BXUuHsK
hmOVkBu/zK/GOjhVLxOkzPfYeBP4kMvnnGxE44NmhxFE7AdBYTgt/KhZzVQy9Ut9
4nUlqQxMtQXEFrWFTiLaIjIKDgQsmJgc0iDTbT+lG/tbdCQeWqI+RiHZ2CARuVl3
X5zcaFKtDal6QOUFIYgMDTKigwihZOjVjmp8W/ZoJmasG85lDdHavRS8+d6p0ax3
O6DQkPJgVPJPsjAvFNenoAp5UKrqr3U1592SJIAVTm4b73Z1Biclbkx9A3q0t+mu
qK1xiQuT1UO6edgLyyHur2h63rGHPnWjhe7Xk+c1SH9iyq46vuj0r9jHKAT9+S2q
4VrnrAL5TpO1u33iToKOCnDEr7hwDbcPGjq0X31x5SCK54UI0LgAmeEKnKT9Eohc
YSF1O1untG/9RYynZvaoDz/ithu8LtPXN0weozlnTT2ajv73NLBBh/FGnVnhV7RA
+NxKhlx1vvoELJyqriOHS4bVKWcn9iN/veJ3RspDj7fgxmchLpd1QUXsYmm5ZDJF
7+n+K6mOubWJiv/e1phGNWHFF+mnlrv/6Fs9aymgG12/hpyNw2LcFf0GL1ZCC8Lo
a+gXke+dAE74/9sB0+cUo9Yv3lMgnu3Hu6QzoiGZSrnRe/hAfujlsOBpjY7CeSFX
yZed7J9kZ9HXwErgfYt9Yof9/YTXeTaCiPtAZ5g1/fUXgM3MUYyhTOavLmkiGhy6
K0uIskqb+ixu8O57mImciof3sVfqMk47/ZMk76jRYz2CprGVRQzKhlGjC+na3vRG
RKRcFeb5umDM/9OydqL6NxNtx0rUw0jJaRVlmNoeTM/qmm3oOExTe4tDdEjVGDEX
K6I7o4kJDr/JvWTgTnrg5psCCDBUzTsEQFMzq2EUFxzVyFU6ZrRM/w2sphkH0MUy
C5Qe7qlqLDqIdn5nIFqvk0aMDB89fIA2kVxanKgoV2dpUrths7GaIdrx8oIYdERi
/1Xsh95Z8f0MrXtw+wrYl4EGol9m6p+ycHx/rqMCjlBeH6slL0SyxNwsONqbolcj
N3npEfJX1cFNxXvPWlGeUN9CTa3BtSum81iJVSZVmg4yK+H02tsUpPf1m2FBeiOT
h+P3M3ibBgjc3lqNrSP7JCacNI64LuQLm3ZlGrq4wwDGJszsaCPQ2IfQcs52DBG/
/PnoQlQAbVbXK80VIQ6mmJV8soHd3D6yAoi8+tx6IrMgE3tLwx9ZipaDCB7A3Ikz
arnw+3GPC0UvVOJYfJpDpteVpCF4HSVT4FMOzYpaqghS21VDFqosPNgpH8cV8beI
FK/Y0PO8uIjO1hCFshZNDJ5S9UZqit0z/jxoubKoYjBNtP8xUaYC/kiS/kgh+6vA
4WPr4Hxgpf6uMiP5+2VqPxI2c5cX+WEy8AX66lI8wg/kLeoIHyEUcm6/ryZKjFuW
L8UMczM0hbUfyTahhm49OLZEaSXCTH4Kg7pTuy4vcsjyvEBUR3CBP9wp/R00x2dA
BCOJYLQKepB85Im5cw+MxiEgmOptxHYJwK364jVw3nFvs4LsfEzY0lD5MFU3hkv/
lTXSkzu7kmXeMQZjW1l6jAXNnlDVomN1omGud8c8KuSbm86oinzoLO03RHJoVWBo
o4vQmgXAtLxPfrRP2HvMv+I9jjMy7K1N+aM/1rBLZ67JwyKkH0frQogA5UxFXu72
qLHDcFSR/b58bSYyKN9hk14vUGfvrA+WL9ziq+jDN+OFRvp5TAniqx7muFCYosOL
GY8GASWQu0b9h0xZp4SDN6SR2nhxDmFx9lRU5hPmso+CcpSSzJOL2I7+AOenkiMe
UTBkNYh9+1TFvHr67hrJT+MaSgCG2uovdw6LyeK01YtBOpW/15qv2o4QgI/GdxT7
c1I5MuyQ2quyus12GeEKTQHdMzXtTZ799bEV70JYyNAAV0E/Fdpir6hnP3Ppq0I5
jhmlnf4TXRYy7ULhyrVm2Sk68X3Ih+BlQPfj+Zwg7GZbbsQfPYP5FyJmyz7VkK/9
F+xlZy7F/d/RuSsfg5qVpyHPIRjWcnNawUWcSTwGNjiQu7ItYWSppGvaElX/SgEi
0aiaANW7byb1xZ5m31tbbdxcB0heDDKmicCGWqECukitR07nScYvtNyI3Szw4jBc
QjyawTlp3TUa0eRQHfuu62dOF04IVXeiF1+F7Ig/RcHPaAvY6H8N3WtT5synnCyH
U7XWPw8rbGauFWHCtvllVILJy0vQEKq5CTeNV4MBUVbUdRiXTgRD597SySKd2BTt
Gf/C1zawU300WBnXjLZYvUaodIZY2P0k+WmJudVse1/nNfOavIrQy/LH96pe0d5b
wT68RVnUZekYXhkMg517Uz9/wD5UMmWBo4WxhZJ6D+0JFZveFw+m1pRxcXI5hwaG
ynZPLUTkFTC6Z92nn6qzkFZeryrigrty/3Nq0cUf3XISeslTpjYH8xUHPEB+uNge
GGUv8Ao24GEftittE0cFpoKYGyMoQQOZ0iZx//EYOFaFhs7FynOPiZPbZnpns+ze
/aOoygwJGRiWInVJuF1udk6BgCOJizl/fmHg5O1tIV1rGB08hDtpMx157nUtD+Aa
UX5cT4jUOsIxlI56Mp+kz7vl61Hr7MGfoSwjaM0ax9fJjPJ6+P2DpcG3vq7EyYmm
Xs6VLqQ6B1Jo6FWpLHSCfanrMx6adROpH6ngC4qteS/vC9fCI3HjYKY0FglE8hdA
shSr74g+AqmnLqOkj1KyfPvYV/8lccDt3+vfL7yNB0jMJb8ZnyJFIXCSJT/xStXC
Sp+aMazT/olit7GFisoW0jzeKYxWs/jvYfV/WwUU4r5IRz1SH0t2SInqHZ0Qny6n
n/0nA9Ej0ttpKxk7+GZ7EeCRsClZCT7mJ05YfCqZeL7uW2fuXqu6KB5rGJKluPdG
j4+xYeTVb4Trz4OhyPx6x6GBJYM6I76CJvzS9GP5HvL2wNb8hvAka++X24EBdFsU
HxyiTC2i9GvrY5L9XD04b3h49I4a4L1rjl4ZQj3wTW5AcGLGSqhloS8viiwKJfrq
4o3sJ1QNidVvhTsEIJw9VmT4I3HQAZ9kjF3vZhElLh82+NyZ4KHRRfqV9CFllbfv
T9IVxoB3pL99JOkcFKRUpiOdU7RPU8O2nnm/woBlFE8flTtobREEVezVnNvRodW1
M7Y9QocMEMrzj+DJSxW8/OEAreYKDklUApKD+wGEqYO+jcnhVDxC9ZFr5Z+KA8mW
hhmEmDC6io+3AxODwzmlLx0TUddIrS2nB7Mw2luJB2wEbeQxCUNI3HQtTLqChcpi
oVspkEu+6rwP2OGeyIVKqb4AdEsM1PEYDdaxfYnCZgMzR0g82GqAAyGDfoe5YL6i
eTvCpY5/6mScN1IS647F6OK7/4xFemwyD5WkFX8urc3IaLOCkrqBx2s5Z7/VZ1jl
awSLVM2V2o9LIGL4rIzW3r2QvTS5FNqlU/vPHE4vzumP/Am8CTAByXjq6YOFpjeQ
SC95vbC6Vwu1H1YV3uew6q79Drw2Qp9LYnSTqQf1ShKLAKdZYK0O7dYw95HvWNAr
KU2abeLbhL2hQMadB0FogUKK/pienGu9WbTF434vTJah1Hi1uha/o+OJOD6d7DeJ
WwUxFs5S8akD7H0KuRBaRYr7d4Tbnm82fbORmRoKlU3Gmj2dvKMr+0fjFY854QDI
H832iHnqz/Jn3WxnzmqvF8/LLJtAwGnC7uiL2UgzQKwTuL9oCHPN+UneHtK1PRfz
WPakgU1XtXcV+12EQL04TgfMHBOteuWyhVFJKuJ76P6G6OvAg63VxJ85H5USaDmu
dBg98EPZtTlFWMtmUTuuXMskVzstndzuqHtmYcVwcDPFuveIbakUN7XJAhun4iLH
ARfKiUrAzKIwrpZCZq8o/mXB4QDa3/U8p1YnPzU+aHF7oGB3pVKqvY8AUWMz5+4h
O2uE6MqvwlKRTuZ2BAs+r0iJcwRle3gkV3PD8xY357yn2VwLdJbI8zG0wjRDuH6x
QST2FhAPQbszDNa42dKUy0y/rIGLoFZ7krkPMwOhjLZTo4nJr3di1ZLwOjnM0t0B
FZX4Z864yPIQgxGyGEfuL3biRaD5kaFNiW82/+uhLg0MR3DP0hdMyzmoENbOkxdc
F75eepuV5s7HALIlzdX2Yjf6l0i5HS+448wujl1wvezMTHEOHpRoewGEkErJyKy5
PVnWbHi7R8mJhM4RcqWnrVVoTT23m5Obr5FchjoJw3S2pILvHebV7jPNqahSwcb6
290qv4gvxwHE8cZJ6IpfkOmHtKSlgK6oqCk08pnCE82Q62qajGz1TVlGF4GRcarb
xjxP9xSE4JV2RvsEUGSg/HdTUt/LJ/4ZFeNfxuxzN6LJFODPwHHItxttxE13seZb
F8XJpS89+oSDBJHhVsDx1HvEFLxQ10l23QgLsZIeoe0sF1p+OKOeJDutDx9YFvLo
tQ2HJhT8EhtP9y5CmZXN7tMPynIudl0ukFeF2V32QrRM6I5ovKvByr4XDHt3Q8YZ
+GVapIDF4/YP7Ff9djM84czPLlwUBy/kX7WyvmzGYoH0OmzPEEwDskHGb1J7hjK+
pMczfrlhArTtw59oc6qZSNrFCaYBFO/beAqpqKVN8B1QItYZYORXWl0t/7U2HDgu
x+iag2P/SVbp4k5iiVIy4RqZoUa5bJuzt/EMQhnxEmZJGLaIV3APLr+Bg4Gr2GA+
D7FmtIQ6uXZ1bjNepqRqXunWzU533vrdA2aT5NhQqZByTrx1NFhk1EYaXH/INt5N
VQABS9swyFL2VAgxtvV3F57EGG4Zt8jaObFI1eXh+1JLRZe8ZLL+2LYCdEaOidiE
L956esz1Sh/lcj2N8mRBPEwtt9C798GAL5vk9OhQAedrxgrGR1OkZu1jOj6OCv1N
SwssFgbUyf2PLpMpcdWwrGwdrZfJ4Gx/tse1nnN6D9zsEoYa0iUxdWIIy1fPpJW/
h7r7gaW/NiZmC1+4qF0DsrQdGHlTSQZqbsPOVe1AMARRHyItrIzr2PvHD+0AwvW1
h3NW4O4KAgR/3PUT+thhco9qao6DxucB9mzmxITNHzWzpZZRHjG2HWPNkgjfzfSj
9scN1LWekrbvF7Zvrx73fWwx9pFekLiWomvTq/LZBvEhnDjKRkQYJTYq7kwqV4PG
20T88prbMWmraKu7SP/B2HwHytMS1embCDHWJcmmWyjGuy7tgdED/sbPS8eu2eEn
J2puwgnwlRJX4MVqXugS3HGFXZwmUYEx7zWJuLUplsYwOnueW0OvTCMfYqTDVcuP
kZxog8FDZPnP18LnBlsHcfUBCxzMovV+kyY32XYDky3/mp1mmjwoL+vO/qbc/9EV
Vcllwxc/IZ+56DrpsFYd8SNnVXfWZg9xVCxOpzx1DYAV5TENw33cyR/+7YsdJTGk
/ZAqkLlFndU17ncF+Dgjh8BDmdoeq2cAi8X7mMA7pXN5ZA2DMyidhGjokvLUcBzr
tMZhHbkjVa+8PvaBBGhp/tWD+tUD2BwapJq4ohyRGE3WJz2JujNgjxwwotWJhD/U
EV95ispT9YiNEa1QDXsqfPbqXR1OLSjrFSHFQXrzJcEcWg6g5cCYny1MKZaTx0vg
lbeKyeWGIXlIVSoGKnF9WbSK7tjezxfC6Cm6cRW5ebHWUePxvg4T1pAcrFWeiyvt
7v7UL0oerJx0JTZQT9mXekRBRaD+ADsirwtiFLFf+MG1Q6ZoLTHwYsxu/6agugZS
v364VfVHmA+LWK9HowJnQcd8unbmcBqFEIue30ugFzbflfSgHNbbqqy1RauwJBYJ
9PpEkPFWMG8J/DpXMAoKvzwIDJbbdpti1lVrO6TrnAnwSn22uAo3XPhAwkt6GAa2
eydjILeVPQ24/1qZsi0CexO2cyFJ1fJQpbXgyd5vLEPBL12LWnO9Vcnfj0qxN9g0
Abu3EwPUlzNiFZW+fMFCmN5oJb7P8WAJRrP3pCLstAycTQ/1WZP24G6J5LnOsw5/
NZQky2j4xbZIj8x58PhWjM/uBe+2TScZ82SUXJdSmR0hnjvzJc5yBCXyvircIxFA
O1EK4ilOSYp4mZhaxif53mfrEPPqCHLNjo3dnCWoY0nBKmyiUebTYHlWx5XXSz0q
O4IlKveg5EbMBFtZBe/MiDEU4vuoMT3UrKyK0o8WyCIDIS/7a7xNrVfaqQVvzVG1
XiDE0A+45IGN+6QW1VDiUTZD2JDoi3RzRFaAQix9dHY4eqpFoWCDI0tl5XitTqp+
KejluZHZanIJrCYaZASQQhURDpHdtNpEVdxgxPLi4FfQByAPT1opkBAmpGoIgH9v
vXqEoSeCml61JSOs0y4XB1WJrYLV3JmOmtSwWSgoSd8u3w7DZF4ESmInEFrvVkP1
w2BWLfu1c5azxyKyXCtFF6h8mo9QQEIfNiSyA4MI/k8qBJT6Vf4R2Lgf1eRaTm4n
s9APnvncih72hswhc11WsunmNS8UMbZm2kLnF0rFPMq7Z2vwSkYhpyE9FnhyMa5H
0+jdH9cGTJRc1XIsFKOhlDsulbAG+w3fwKpm3egv/6wbWpu51reVqAfF9aJEwaVq
nr2H62mq77Q6NoJOwwsfg7BmutmdtjpjET1BwQ7D23lh6Udj9qJYQ0eQ3mD+G7SL
q0CBIdRRTRDWlB/yoCqPQliYTXBc3ElRAX/Qsw9o0KK0xlm/SU+qFTwUWxJC1GBv
Jy1KFtxFxs6inFSpt3JiAIhgBDgnpui2WiFSU5uT4gx45MrzqBm+CdO+RVmI3BLd
4L4RGbXYkFFVgIG0hm4iSXJbjvpQ3aarhVLn5+hjAZton/rM6rm+yS60Zsn5Ezp+
1Iu61SeAHuIlKj7D/kTBs9kRHvHXjV8JBbUY2lb21weyDEXkGuFFpd+5kekAOG5V
u7ZoNHi6kY1dHOJrKhTX9jvt3O44sOPXEB7Dp7oEIk36dHZtacwKBeTSPEDRpGbC
XBKcLoPScWFIraJxmZqQW3+cmaCpSQtJ4G/uarCoiLhiNX0Vx7657l6dRHcioIt2
JXFiT54THKjq+qIsSS4gqBHdea4z0dOv9It1Hi8lmEl2KpCpsqWnbOngGEoWeKKg
Ds8eA91TjB3q3eiI6sWM4qJQgaG+JXecthB+djLegidQeiXItQgd5m1deA4Fe+4G
BpWs1jCM2ECOTd8tGeZw07ScYnX7eqnRWG2CWv3C0xNwIOuYOpjh6KVJC6nNPMTE
Oj0vsNdn1Cr1V2AIV2kpdOTutL3c/1mm//yeb3ZLi4num0fj9ilPNxKpIvIKwR+c
n+1yNJYZqMwrpLb+QiQh8/xHx6ne80Gq7cTKU5xK3jt6PRZPrjdcFclvI054l6vf
xLiD0+SdHHkQ9w84GQzu9GRCDDMMmVYrCtKQ5rEo84cicn2HsJR3pKumZGmOR/p8
hwwkC7YJJB9Lo31m4R0U11yx0oINj29K4mVjFqoFAggWut3pt9PpSpuV+Q5DQ2ZK
7VuEJd7zT2j3neGHCOZ/zTc2gq0zWYeCIWaGsJp2Eptq6qshQ5aQc8UbW36+3C3U
iaJKTwobHWrMjtZKPUmocN7JDy5bePze2p9eJS5DhknjzYhGOISzhDEPNp2deD7/
/j/si4j6JmirWese9dAX41GIW1IETeRSfzv+DT8tNjTZUUJXlqla9WdBhB+OA6fe
Z6XErRnPiuDwzwuZcLgMTSH8NlGgx1rHugnuiJdh+VSx9/gDSHxq8krMhRwFy+KL
v5CSz8qghNvUAJPJOYMNTK8X/67mOACyit4H0fIQxaCiIdzzFc4TLYcALgptfqQ+
2+6PPC4GP1Ugeq2HYQZT5nZrj7rFjWyKKiKp3iNU88MIg/OSTzEOdEvEEQvX+XYt
RTtinAs/agsxpG9apx5aPZX9qXDFt4GRxmFOBLTQKum/rPMnt9LMDl/Rb+xiKMSS
bFPLYrbMxr0bvG3EI/Q1R/1+Klbg9QJJjlF819/rlDx7zMu2mDNKJwLFoViqsWTQ
v4Nqg1fZLC5U/tjd4cczm0GZub3vK/aeKAqRxxYHx5HpSyLAw+Y2B1XMfbjfr4lJ
qq5LZKaJxL+r0kEn2mh2/SJ6/Q22FPriUqU5J207owI7OjjaMoR9hvv9zpSUdESH
gM8D3MIA0aHcLDx3MQkigQTgqdHZJU7F+212xhR8vvm+v07GLWYxqK4Im3QgcEop
BPsaBXc9n/eu97Se5AXQdGuHoFzThY+4QoqGEzKQN0AzW/JscRRqu6faU2KwUYFV
IEdZfg9Rjwe2SgjnIr/3BrDMRBqXV/O6ufZXu3ZXUMs3k4g+0Q/WiRLdVYAnooU6
LNQl1IbsNVn1+E5K1kIl8jSKw0CRI7oAfB8s5gTHCB3hz0iOK/Ys2uP9eUZGAc8r
z42dm1F2k1qhswDX0alQ+rsEObqOSLiwIKb8kTdugi/eezLzUn3S5O4zENcNMvh8
5Wactyw/k+rajpeOiJHJ1FMmcmo5qmkHds47dR+uJOWMnSUM5GlxYfoyDHUaeLIb
Ydo2pCFKAkib3B2B1SJbza2cAcPXY/TwzVM1CdLPPiAbgHv8+/+C18E+l8MRSRXQ
EEky5g1/7YYgf4JEDGoJJ98etZ0LMWXiH0fdfUIAAg13zOBjeZtTlxITRs9lyOgw
Xsqe/ULjCGqlxxoSJ0A+3pOnJQXxoRMMlUPEHFID2RtJ4R3qe5g40fRonTr6ff2N
lBlmDN8J5/fsQANPuA14Am3z8hx7QKsAPBbzT/vCa8OylhcU4spqF8DiCu33srWb
GXTKvxBG8cLrNMxN3sGmuofZ0tp/FbjHJl37e2VgOu02PppEF4lxVZi5A11WmbHU
Eix3Dt8cJ3hwOt8n7R/oYZFpPCPHiH9bmoFwiYQo77Fl5t7eo8cgD+/553lNCigi
HRtKrH3J1lxbBCpl/GlDYZR2JULt5xg898eeOjOTv6/GGlhFAdXGOMkcHn+4xciJ
dY21QMxHK9eUD1C/XKBnWA/5zIFBWC1fc3eDWh6A62GOxxJVpBV6nPVDlDB9sOv3
Xk6CN8gt9MC+vE4i5qb8aVmNdGVWJ+UfY8JDKXOO6XOczixScJmIF28xgM5EHvIb
OinY0DkK+LvWYABQLDIILs7zWPMQlOr0u02Tjl0NslVyTorDN7AZxgdkIXdB72iD
6EsTu6u6ghrIO66XzhWjlcKdk5RSvspaWCyuS5WKuZDIsJ8Pb0SiKBZeh2ud71ME
0lzR4td+yTcWyE4i/2GRfYP1DMutiYdrJwhJyT/vYGE9YaNlD77qEo4xU25fk+MJ
278vjD0MZ8qMtd53MNyh2+JZb38T7FosDEz55a/yCjm0nJdXq4b8zxt/QDV7YD0p
VtaJ7Su2jKvATJa8zEz41LSAHhBNNq4O2ozmAJ7z3viNOpPVvOmInpG+mZz6JNeY
BJ1W+HOhwB0hHmY7VywCZXOQBn+Wm6GBSFQ1ryLRuHF9spgGJxtpvsvGas9+JPRh
JhdAOPg2xITuZF+cHmBa/zjNDOTlMI1XSVY2FrY1r0DJXSkF0d/ybny5OIeWRKIj
vYreiq1bY/Qiex2YjW8UqQossqMa4hTbJ5/5X4QwQLtAY386Lhw4A8yOa3ymG/7l
BfeXrsFrelOnuQzuR2eHe81UIQPzUB1WyM+lEvqmlDi3c4to6TvFPWf6in1FrcOL
Y7WM0IQEBHQoGjlm3ij7ZkVP2lIxyX+syg4QkinjMC9x6219dLu3uwr742wk4KkW
UsOS00wp6Ko3Lrf9p0qBoepw5BYNZoxF0rglZ38DoDkP8dZF1mWlptu0ifjMWOAP
pcCkrncXwZv31SVxDOzjMIWFiepyv5pN2q+RuIIUTLCrRh2S05TeLBPwPm1mYSJ2
LOfw5IQLLUw+8CwMOkB3OkrANMX9Ian3wo9xFf4HCdZBIoEDE6Agdwv9d/aKsKMs
pwjGnPEQolOgliqqSR3YX7q/dfG7bo2yU//2Ao4jdB3a5HgBrsaE1y00LsnYPjIg
zRy3sqEgvJv17NkgxUjNquX7MaBPdU/wTVWusqFl74AH2lUQEXx2cQYM5w8+xBzX
hX7Pct2iGpYxTmTjerrfQdktuk3ReYkv84WjU6CVa65/vIabb4dJsaSAZUau50Pw
ywaVMw/QPYciLwQiioR2tXwoCClXqmctZRuKrcRLBUpfex7+cUb1Rk2THcl4SSoS
xmSEhwS9vHGvB9eQ3YxLdFx8HIF8xwgvaYDFx2WFS0MTvyA1mTPFhgD3GH4Iz3k9
hRAkL9VNQLCUIEtQilifHLgaeOOw+OqjNz3mL17mw5/onP1naI7jyI6gTPFVeAbq
I1MYq7z9KdkvSCWtJDvNQEPsle/PDVWToE/FCaPEEbnUE5/dpPaPhHpa9cQOhgyK
/aGp3NkpprL/dp4bzgjwVBYVpG6vPVD5KDsMRyO8NBNwuQHPiY+KOrBfvBLxBkqN
AsQC2qfSsZlFWXqF3RQefaKefzkag9UcZCEsp2/fjZkrA16r9bCSoZOAOI/fIBxF
58S0r+2bWV3/rzVdNnhFMbzHjpeWsA0tXa2uPK2yuNOjSKm4dL4mvulvVJEOsQze
DggT+JCBvSQ7DTQKR8h59PInUfBEtJUc8lvQz3HX/uEIQha2z35nNSAkIxL32BA8
b743IODjoOKfMZYJHfGx73Dbx5LUuacLn4aUAZbPtXFKHb+u38TFmvqF85Rmagga
0j5Rz43akT8G9YKiKTjHd5+cKC18rbz4ox+8UFKkfKZbwF9olWMQho+6pmVtXtJo
6xZm/QdXFeB1YdQi67ZlnHdKZX6hmT5IdZKI1/1KzZV2uttQm3VDzsvtzjT9grqF
hI6o+EjQvlDo1uYycOrTzCwa7REdGUjMfcHCVc+HlHCQtKzYxlCkqVY7/ax2Ztxd
HzwpWygZ0zqpEQl9dejx28KtwfnYQoMIw51++qSxwSfJ9xT/ioN62nt7tAjedysf
l7PgFg6U+YSZvt0HjiYq+tircKHD/5HLTQya1sWTG4+UOgPcgQiSTOTaa7uhDClT
X2pRVT+zVGH6KIGyinWI77fMB7JokEOjgEPF5Of6yROkNtlnxYd27bYOer4uyN7F
JmiC/C7wvmmj4PgVJjm6P7hYGCegNkkTwXeraNyCq3aDduKYkPVZbDXhPMOFG6hT
B8u04icMw4gETLSNE+sa/gSqBIllM4h6/Md+tQWIaEnt4MBGGazS0HIz2HScUenb
ewgkQZF9sE2luZoLaolOjJuRtCLF9dYpTiAS1lQZW7BbAmEuDLBPNjo38NN4HWtC
lmM/27ugd/yISjURDPr7Xu1HZc7IAf7kaZXcxF7uXaOZqHndMmtIto2Gglit5T5k
RkLIQdLpMAASnDCKKAV3ZMJRizaPu/RTlnVYqUtMENjgYSCap9WjQDs5Q/AVZuVs
tUrE1qAzRVkmILbHOA85Lv3bEduzWb7GwAzgBh618pu5e7BFkl1NHwScWMBCTmNR
e3aHozFswf0VxlXW1hf/1xcf77TvjU8EQ/iqJbgilT237ZWWLA1cAfrvwNdqBHyl
EA6AVz2oOrOkCwKYfIaF6ctiwe5qTBDD31YDCBXELSYMVFsT/TXSA0lvdd6xzZpI
LmsxqI4iHziWT8H2zRfSkuphdspXVqTxiK61sgAvJLDaKNvFyg3ze3KwAy99ZcI4
wIQxt1ca3saUexgEpGbQH3wEXG6s05Jl+MxI5j4OvuCqxVc/g9RefPgDva7qNo+3
tLcb1ldfLYWnCZfLem1ahKzNNaPSAgQK6aq/elNxLlM7aoEZgCyHJ6mgKoGgyyc9
n7Tnd4XYmvp7SgbxuI5ksLcO6xrtb5+FtkJQ09lj7cmbm02UljspuRoL0aymX7xT
P69ZNIQnkBgV0oacwHHwkAXeny3iR8DF/UelilOxwJirtC5FUo1Hh5U4OD5rOvcl
r3gBvTLqVqAnbwdk2WfBOeI//sZRL8FM8SXQIhY9TlOwZeOz4rwFaw2j97oRlrig
YlkVtFF4VDyBj0LfjTUKusTuBPHiKWuuC3MnO83TnmzJgDEWdW3X2tTXqN8PwbJs
HNDbXpPUCKgWd6pDSeobYao/PvoxWloWu3pw3Y5ioqAT1srExWGm2L9wPOZXtbE5
TsUao9ZmcnkxcZGSNOpV9gPytxHvG9wON05uQcVpG64uz2vqrLpqrkXs1uqUQEgq
1udiOPfP8I+TFt4z3VZ+IHzjOflN4fpRZPsuMFYHgeXasERnTuMI8PDbd5ao4rQs
qeImyD5w7k67FWATVHnFP2MVMKg2HlqS5/p/Jh0nScM84wZgYnlRwR1txULlZMk2
rMEntBAIZMvwcAq0OR5II7bcs11qVBUD+NDv7nQqvIh6Ziyg6QYF2EDt+9oXJhUC
hv5HWP7414Hk59WOXHAhNVTbPpR/uUhusLjQ/iZ0bLkfrQ3B7HwTnNobMUje2ZCv
FHoSN4mUffxSCW0xPnMds3LUCuUcIphnTeKmhfJs1kK85OW+w8sXLLrw/IIp14hJ
75BBZ02mBfhddF0uAXa1EhE3nMdjBAh1ilwc7oKt8KgRw5cThgqqa2ov/k1F0ht5
M3PeC0F1Hg+l1ILELvwE9HELt7cc7vOJdNCUwqDB+12AoIXJnvjbrXaJNLNRQOHL
D/RG4gyMhTvVF6uXO6gv/8XKnEt2JB+n+RQW7RqxiO/mWGBsd04j1UvAzoYUmUss
//XcgyqvIAJ5dC3cLu31Wckcn/ernVDH+3cmbbc0gTHf2jpunXlBtBYvEFXlDFKI
UTazQua7kCrr4bprxmKd1DnuGniLX83GbtBRibZsWQTUnHaww/uel9dw4U4Q3E3g
PH3GIkmghtdLeOte4sqKS9DEDfju9jKC3Tjjm1QvQgxTYQbYcsxOsEswCisZDdk+
DWFm0+nu8bdzq38s1hDz44A7ZCA+kpTT7Q/uqy/+Pgb33oSI2O52DzhMmkqqlfoM
LoedOCRxIkYO2q+5x/xXWSLAjVxhxHxBTClIyIaKRVfmwWpZgir8nXB5CN1B0pE3
o9lLYMCDtfjA1phRLBi8r6VNNLrpvB5aAsHVvI7xFRWHzUHP49/TWPsJ0EsOdGqf
r6seW3qvseSPKk3rpFJDTw/+0rOtOACtZOCCWjKPJ8YZN+DOcFqzux+aOC6qe/pf
zCeLr7jGUHh59+9t1Gv5ayvyVbzhom73ROxS7NXnbkpLIYIbXO5WISRUE/Rpl8Yf
lNN3VJ0TmG/11yBUmpxTteyMconIUu9JJxicYKObAJWdq2032poUNxZYOM1UuPY8
ib3JwIsf1GGQQV7Dpo5WQOL7rFP+vdoO/7yFDxCIpK8DySAhxm4hUjs9SLvKdv59
WQxG+JQhwVgOc0JBWiEtvKt3uA506+6juhNxtEvP5JSaIAsE3ZpfGAm3KYd6KdLc
UC8SXi5pGFvcLHHE9c+3sWkgM2MzWmzuQRLV6Om2ZpzeKKugdsVdq71NnCLTdBRW
fwu53vo4uHNb1BEBlGGr//1INRX1KLt4HEhHvIVNYuIt3w6aEqPX9R1yqtonOxVW
49SFKAw9jxo7KcMy0i9aprn82E2XxPWPH7XDoki4zPhgTHBEMEEx2wg8HHxBDkxk
z7v3I/pANA2l/QPbTGQOGkgASK9T/41YuZv/FR22Za/N3wgJL7EE6GB6TUWVo8rx
cIvMN+05D2Fut5BSzVipUfQLSyFiw/5B8YMIAvI0hqLUPe0DnEWh2T6Fc57o3ssy
2JKCllPDCxkxNRZf3qOB3Elj+XbrFbMQ8KMEy66fKNoVsoCs6tKPhL+k7bnuQBD9
e3ulz22ThHBSBHfnxb3aQf1d4yvyVSVEowOAMfUTO+vu/ScfdCNcLimbqXJwE7hy
oicTjeql9ZhSOrYiH8cM4ogB3vsJumuhprxU+jjBb3LpwAFfLxMKCzurBt7g/2iz
GJBFJigM0s64Rzo3gdxIS4MUgn4LM5xQr1becYvb2YXm24Mh3Fog3viefk/xZ4S7
Pdt0suatomG7JQRtW3yDI8/xNaiClVnqwJA6oySRgSao/Qc6DWUmL6YHs9luyTQM
VDHyKwGnuggx8YkXzEcL28dq00EUBdGeIOKSf2QxX+WEp2jZNzQdwwecQG5k0PYg
NJrruGNORwSNimt5K9vJId+vK9fufpkh4StHuck8Nf57hxGpPEvlnh9g7dD4KhEL
sbNraqIcnIx29kN75Ps3vMzgQyYPEXzW5Ax8tFiXebH7NHAtnvSe+W14NJ1+LneK
9w1g3JWkgABvGqi/DTJgaWv+xY83C8zykoR1c5hMRHcx0Y0QtS4N7V+IEKNQ17UD
VVsKklMjoEBbzpehkLcFJUXYhe5k9wiynoYuMkGHdbyA5oHzSJB1BTOt1djyTkqy
oNZucAzEQxKhMhYUMBG5/B0j4gk86hg61JOKI5IzXXZnmqazoY7vshzHGfAoAO/O
Rxg8rIBuobNli2pF0hrxZBxlSiMdF5LX8y8U8nse7uuF4IUetEG/JFeoW9HVloKo
RYsY29vyTKdUOHYQCl8ONz3K3a9DpIYKKGOYxdNFRvvgsROAb0AEZcC5tWhrCtKD
QcFlk5OIHMcBoOXEHiXXoO2yT5bLyHUxUwR45NXdO0vhF+XqnfqkuA/UmdXqY4eE
S9xdVoJgM6WfI310tvYLlgosACMizQJgldcbXR8pIs8VgLKENzAOgD6DmUE34ky9
j4sbkeYnYEV+C14srFyIvdpBRkbT5RQEHbDDdDoTDSrHspX1Yg5cy5fy5oYzCVfq
Ey85XescL7Wuymbn5uJzotIsZxZX1BWDeAzQcHs6LK+igHZk2NAW5/JALjSGM2MC
uVT//QGFlgPNQwtTuYEvSEGPJJ39j9uvAXKg4MbK8UhUkHnH6M5qVsBhApQYh+0r
HPOkkUJWHTaAwyEzRJSnG5sSsBa+NplzkaxzLrd/kYgAY4Vw+VK2XPWTehuIisdt
Zkbs7bjDB5LjD+5XFf3nHKfF2c+hUGbatGUs75M+st72O55mPoZPE1+MABZxSa/j
GybYvqUyLYDEvc2wOpH1m/rUUgMMqeqLbJah7tS8A+LvIDn2OSiMVi5eLhC4zfNE
Z59gU+BkwNjKNZBGsbLVXt2DR2Hn5RDyXPw7j2HRuC9Q/VCsbk4585QApPFp2KaV
OiKz4HQjMaad4lxEyECbGR8FSTgYko5bCoswQELuz2CE4JwkTQMoMT/7dB9FM+SO
Ncm9zdc4wkjq3xEH51Rq5E3qxsJ+ylyqHbbu+B3ENUF6AniedJ+hLLdzIq50Chwc
jxzHgZCeDbsDqs1AJskGaiIb/ip41lqwNgjEgnITspMd6r7t8mP1pYx17klCDFJW
Hv89vGfp6RXepCgkwgSVM+S/nl/p8ge6X7KdJYwtJ7BHY2osVvZxX/vB4/D7FvW8
qXQ4Mz/98yzFR4xnySu+yPih0gf0NHGOtj/XPqHZugMGBnb9om9wmCc+QQcb1Pjg
NOQBId2Gy/6Edz4l6cbhaxm2UVpGecrDOa3FLQ5DgGPrgA/GkMDwr009D713QZ4G
CsinYXkgFInUNy3eBHwMLOogLEdK/B5vdsnpunUqQWLgtbvhyrmUpmcZe8YuGYWI
HD61RWlsI+AldGe/W8BwPvWJO+8TidVS9MJ7IK9OW90Ege24iAvmoVeWps5oEk2M
Ep50pw5z8ZqRpKkDAFG0Hkbh2byFbxFYPBiwpDnmsNwkqXKetQyj1NFOg9cU6wls
kWxKXH7r1pwt9QrnhZ2/S1/6U8DkkOjRY9dDVPRcuVA0R7oWwSRBkO3TedVqOg+i
aj3cixedE/etLlN2jZJMf2OlyhzNz8ypxt72Cy6Y9q3Zhv8cHY0gjuIc9Ldzv7Yc
/iJtpqFiPIiDtT3nsGb1x1HPNUo0qE9MWHMWHBbjMvBYtOr3ew6vB7IMPfGHd3QV
qV1ECdGWnHuIqUZUYyUND84GswWk2nENlFu8cDIRzCKcbA4lNrLCTsmvcvL+P7jY
ldMaxxeReoQ+mIJQUL6k/KtGsak19ZtpHMZO0IO7iWkc8yNTnnpjs/jRniW/Oty+
pTPh6Y9BdJ4rxpRgVj/igGy+LIbiDH0SC52IV1/eDVmgHk3jsi9mxVAGo3JYbXhs
SdxyKZnGBq0m2Egj9quQR/JOr9CqSu9X5UryHY03vQOVWyWdxOuXiPi2fy0gTUh3
nkx/q8KcGBpZbpp3lbF//44EiGaQfwCEBDXW7Ur176/U0MFf7Cl0cYfe/zuwTyqX
G1bLkKYFRF89CmIISlx6JhEvqK0UCPhC5kiuIBtPHA89jUo+EGNwUw0VO+QfzLou
NE4lnE3vVmukhgg1DFZN9jqtv5elL6bBVGdBxbrbO20SHcSEISabBmWblC4IxaSk
0MLYC8stv7QvGYqQdszoSSjorZi5harpq6h7ggtwJbdtr+pTM57aR5LlOvF6Xkw2
oCghaD8uUMEUW7U2LwDG9Kw3bEhzi2d/wS5aljL4mXUZZD6ULNFdhfx9khpeZkaP
jstn2A28qyQZyq/3giaZ9Qz7Dh8GP5MWg94HPYK7IWAKegC/CrfG5RzeTcqn14LQ
gBHcstFWCv1z9uyrx+FHuRM4ZxAC3BDl8EBmn/JBF4oLcVPok/eUiYH1YvHSoEYD
/ov16jUwf1fCM8XbbiwVdUuP0+2F1MALyI+elLOZsJj1iPp+d0aACGW0eLq96NQC
nv6g7MRpK0layjm+1V7B6J1A3Mhl9Bu1I8LNM5meqTAnI/kxGxJMOkKscW41TJHQ
WV9q2n8Mq90gtKkdBcyHnkkLSi3e3RozIQmxUgoSJeg1s5+DbjoRhLArbFGT9h5C
6geiD46HXyPagYiQSDlwIzhMYE3zicMPdMH3o8HPlMr+3N84eKDQJOg4HBp3LG1e
K4q6gUXUj0jIxcWrHakLa++B88oK6mYsz6BLa8eZB+bSeamfmPnL9LuPzDhgl9fi
JR/dhffW/LL9AUJ2CPbguqHo6BnkWespfofiODp3MRRzimxj+panJjvDHs3i0g4G
9R0r1MVJPp0jvq6ICMD5SBoew+nTbUy8O3WPIm9Du1yE24j6cLG9297vbuUWMKTy
8AlIwEkc9tZAKGFOQ3PKG/w87ijpsf2dROnI9ADw+hXvxU57aTnIdn/Iu+13UlsT
+WsX9/V64R5uSey/7qmezZJBg9R8dlgGlqC2MB5Y6srGDJj+zFiAXDeKoTtyTDKI
jzqt4F8hektvRZYlg98pBCtZ4TUfwwenLMRAlt+A9/miR4XHXUGRjlFJJSaR78tH
I8b0eKVMn1jgva6oCaBFQlLI62OJkMIwcRY3W8zZjd0bvwo1f4Nq+w1rcllGfFwT
EbXGPWK15a7YMyWp9eDUxE+OJ5VGciEAMyJfQPg8ibKYJh5xS/wlXudweXi8u1A6
+sddUWlIkr/d51JDy1bRlvqT8aupapNh/XN0QXyKCRyFd60pFIjpqoiGnt5abVcH
GFMR9IRbiO8dEvTsKH5viVu6zLgjA/AT66O/KA9BMDcA+1FAxhdSaDuRhGik/UYa
F9rpnM7wdAjg6jTmXROyh8bzN1j1MFcXWArIbStxoVDhACFd3esTQmxtob51IwXX
qyjRz4o5qkExiDXNhLIAZLUhJJCHW+7OFZfi7/gEl1e4L/d6fAZGtiUHot9LKCXL
abP36v44gZK3zD+R4g9OTTaznrkExxGELIj+IDbeRHDnBrWsSE6NUJGw7SudgsZ1
PwOh4F8VozIMJl92QimW5nGa1IMYNq8GQNInTMv7r0UN5N7YXdxJvFhrOBjQpkWY
8iYQRLgV6J437QNWDrAMNa71gOJGlVsgwR9gWIG48P436ow9PF8P9uoNA/EI4OC/
ccFBYt5ouhwOCwuxJOshEldGt4cqxeFDYu9hsrl9+7fCO+QqtSp6sDscEjCYeHwY
DdPjK2dAe5+TVlPaPBhqc35Vwl8DSStobXtw9YGA3FDGa4KWob4CHHrYyKH+Fh8/
/n9qOi6iUe1lTb8qVDLQAAZifoXO2ghPlQtR/NZSqj4i4f+zVQelneHn7qwXkKpl
3auo6dB9tCT6XEDWoXE7CC/gE/9HSPIBAAqPTdUKuYunZL676d8ixKto2IES9SCC
H9fsF0fo8qJuF9yXxKeCQT0h6+xbKpeWGHKaXgn6OYY6jgj8im7dQLwNcwulvt0e
tQjXt1VCfceBQ3zPfVf7VhpTy0MPOBdmIT2XSPucrFbPSjkuerDsebC35E6rdkKq
GcdSmuhgxI6haQCE7Iv0WXU6A8sn55PxDn3ZP/PFMjLIeM1/6pbCqafBMZtS4It8
CHDE32H6U/h8Kcw/tzw1miZtS0kra9Y7Lwi74hxqaEJ1BAevTOIx9geqRix7acPn
O7YwMB9g4PR65K3pcXRxWAF0lIcFwOir5i/i6ITJQBUFZRYWl6jI4JIpN1S0byzv
SPosjRMk6XoK1cUVAsBr3J+34mqTH8NAQ5Rw4IWXxsGVPTqZ/L7FZfV1GI3zY7j+
j05GNVyM9YHtlYaM9S2GITfhnELNZ4xrhgz5+5b2IZW3s2V/OxMvw8zcmgh4NsU2
Uj2lXVBS06JwayPfJpKoCeXGxFXKkGM+vcPrF03RDtT3Ppqn4DZgd0FytXeC5oWe
PVnzK/4j8bXuMj5pfPbapFtmB/UGNUO8GpadbQt3GDArxA5uiZ2Q2BYQYoXdhcsz
TvUJCUwfuu+etUeksjo2/tgH11r+zb3Q9ZPWYz8NL4N92r9eqoxfJVvincKWTwxU
7iiT5wHDyuIBUPWxYHdV1QSe6hGep9ff+DzXV2mgNmefyzq5rhleNPX0FbXe+oK0
r35qGblFE2zGxZE3TczbRpT5EvlPLQXioLlCP3yDQFV4VAUAflZQmrJ5Q5iLs6jt
0pwgFCAcnqbtqdVlauH2UAFOlGZJXTJy5+pWIcUspHfjOCUj6vyEGIDMV9tmA6RR
53sMVqQ4L0RoxTQ2IuuWQuY4PIG6fTHJN1FrT4+7J7Z/XowIYgzJyDPQoOjJ8+dd
589cgsjJ1cxNMIafadLR/l0T1fMaAVzHKdjVKIyi1IqX1pVzJIqUWy8ShAuJ3l9T
WBsjJnpqY9YOxZdger7Tqk7jFj6JTRup5ZoJMfzWM7dWI65QVoySzu/SCfCpQFdp
Z01eCx4WMamfS6LA8z8iRYjjTYszvTwoIi10ELUHUMwxhp858j+695K/traAHIQb
0qRBQ9EP7xGN/79jFnDDSUb+E68Mm3JCbXP2rVNRLv20gnCn3D1LKV3iyrcamI00
IJ/UcP8sf5g5VAuFq1NrPFVYD2Zi42SchSh5RWb7YgktMTd+QH83iseuODrEYIBE
BDCHoaKHdixZeMNp7mqdoWrKddYhhOPzmUPq48qMY5fluOTLhX8vnM2lTEENp51Q
QRkOFLTvi0lbJXBA7eCxwOF2//1FWkzZKh1Xpf1RM4b0V4es39UPohRkA3M3vABp
MR9XBqcIa022oxwO8pfy+2/NbYTtmQfu2nLR8Jv8JxRXNZMpzCxy98dxtFm3WXWV
o69dfqww3X/vLEYn/59XFDlSSZmQ5ZQVb+hY0kxfXP65JhZJva0j7xeBYgYUIeM7
bO5FuBtxpb0Km/rjBE6dmy9IXyIUrsozLpR1H+k8ZTRd79w9q+fJWfZT5BGocUFn
lslrbyE+HMQIuuck/20RqjMNztyGpIqTRE0yo3WKRShImTyNVKwXRHOFdmvEVtxB
zJL5mIlbaUN/c8UntTTw89bgapAqE/bXrmjD2mDhPOREuPvsmL7cWyezHN05IER4
RPUR/sMNbP2uMMy1V2irBgocBzVsHjtdduy9tdlF2DxXFkncYEdho3qhBd6sQ+1t
eOhaEKjdePqzck6U1D0NfesJWuo4dc53hb83D5ArCmw9TpfwG4viNj5xIUxEoHjd
SpkXxhu2rgXMjxO9Eknzh6SoBWx67VSura2Ni9KmhMECjfFpMZUTsNcD+oBQEish
AeL/zU5u5+b+370naG5M+voijPF3RL35BcGO9HQPjsAox7i4syn/oz7xESJ8y5by
NFg7QsxTlwEAwW/Z/aQPtTne938WS8K1yfbm0Vby1Vi7CZwF8CKGFT16Su9LbGSV
cAnFqCwgEYhFVET+SpPLbrGpVtuWDKgIoXkhImM/gpUHGDkHyyvNbkbCZBoodjRw
4XZUWyTAlrz4gGNTrgB7k9y8DEpvIQtzXSf0SpGiDi/3nMcswUxDAPgFLEvDpPKP
sdb3Inrpxj3BRU+6r4/Jn/VmUx04WyS37HIf9ISc5+GmhsiRd5rcMRTCOydkLNFk
80Vw/rNlFgjFTlbXTf/LSevzf+QhXIJKA/XJq6oWIvjclzwsfvhbnl/nsUkROFKz
BTzz9Ye14HkScbdNZSTkkKUZb3btXrDHlaIQBlH2Eefg4E0mBcqQpXRZw7ReW5tD
DeWhFmYWaTi0EhhiTlmnCy1oaHTiOJR/zzQ6EQrNwkxTd49iA1MHgjOVEE6PosuP
XFdE0Ea8IT5OzxYaEqz84ZG2ddbG88jLmGEyMyBwXQJ20lW9zbRq79+oxKPShe4C
1G1cwXFukunGikB59Lexm2MSlPPbqMBuUPTiwO3yTNcq+SWExMyq8iUDPv8bXCw7
WXcGZyooD9biiqtN1ZluAZPy2smQJD+yALGdxzIfZCcVqQuZ7kzB7j0E4DDEjnqN
g4iSc0eql16qcpn1tv769L/wgdnvhe1ZKpdBIwMGbr5rRTRyU3cIukWDsrZ+6Vp0
Dp21vPL9JzhmV7trJnFDHyNMExpS7Gzd9w+PACUUEk9LnWI9tgkI2Pl9FO25pSBL
11FIZDjhZe5/KZwUv0WaEkUB8x8C+CvqIe4pSQQXBlZID0qrbuMmFJ+t6wCVMtWs
wqaEVGkxiKWGVLqYAMIjboKTf3xp5GJoF+DUq0oTrHO2cK3jmTWuXU3UxO1KtVdY
T/b1OXBeaP1iYyrq6szNWcdU6p+tXDATLlIav3JNpuO6C92PLS6hoVa5J54d+i37
nx4YI1EiH/1kZAZsIa9TVz8QQK8pChgb44eF1owCjoz2A0DAeq64uzZlnrKwa6Vi
c8Icf8MMB0Si/dEZfc0XbUpWmY8+o2K0fnxnQRsuYDzMtXc3u85UnfASAozdYGuS
R2CIghfRmODCknRaP/dOY9osiBCxWaWMNlKx04fGkRhPKmVPBnLWI8KlCkX+Krg1
j0sSoNQV+PlcTjlAnwIGK22AW88qQbtQ8QdEb8I4NYc1JCHhQTVW8N263rZYugE+
QEG6BiloWsndLApRRMJnFLm2M+s632Hph3B8aYF7UIx+ktPHhoq14yE0S+WrElIF
PbsuUM7ljmcmUhQ41Gfk2KNJNNQAIFZl1hpE99JKBJXuHUZDV9IRvRhRlgzRZ3rU
xj9mG8AJSuR7w0WIUCSnINVRBfb7lbtWDzoupClL1zbHJo0NbXNgy9D7lVJTcYcM
HT1u1UsPmK345KRGI/YJdPsEKHW264ni0cu4hKXUHlpAoD5ZOKdDDkUpbIXhTKzI
0J+jFC8Q0ssOFdw3U2ufSPWpsELsQ3iPSAscSF48uJea3hfQNcaa9969k09aKeRd
x9cLyuIdHvdQosQTHqFY6XO5+tdAE9PYOmwcZgdrWtqvfOEYUkI0htH/DFKMhcUK
DP12GfObRBfagjI4jxfJEgLlx4PJ8jdWrrSUpD/O1oy97Zuw2XvyBRK98Txt4iIj
xq5rO72zQsu7csnYIjxfGCWnlKyC+4G0wpGe8WgNPko7TLLfqTlgEHYatCk9DnZi
8K8UPgcbz6YyVphgXDSITkvGqNf/TE3rBu6xJ+sCw+yL2t7+i/mWz7Q/SPTVcMgA
69WCEcxESeeqedomIDGvJ2ulscILj+JDvpfcz8A55s0jVUD/+ZvZeoUml8S6LpQf
kzgRDaiq1L++NDzVqKU6Xt0Zsg+tedmsQx5BmvQaC/Ui3NzeAFX+YaGpJu58DmAz
gSFIiAGvThhbPM2dnMW5kDb1g+elDsLXYkTZJDj8xl0I+B3BIBbV00vYZDdI0XxN
B+b1S/0awEP2oB5eDfPcN6DN3pZPNRPn7K7d0jDf32YzQ83+LbV/dn1PQeIkqHCz
JFeJzBH6sZjlHSI2Ji/In/cTh8wGG3fXtDuHN3svITfNzHhoEdLeraD7WaMpkPE9
CQlctaoy+BE6kyaXFczb2SoQpj07g9Lx1+XVVw5KTVdFfm7hFP2btAmSPeDkJYh8
PT+HsVd8hKpWBl3Gc7eBFEsnZVfA1QkD5x6cMqa3XXfDoyXeSqnNfcO2ANLZH1yg
RNl2hEGXiFWRLNeAEX9Im3bxGNo/7A0siHYU5TvIMpi6mVK4CAhzfyXRZWq4pJP3
H5G51ly/F6bky6je2gMTCaWkLBGYrfiidRmFnF0XxrqUUoaZA+tKkXYVaKrjr0LZ
FlpB2xPAsxQMUHSqD3raR1DgqH+RdMA8k8XfJeX/wYAaBidBrMYYHhqtFCobv+Ar
6AFLAy+Jz324VF4EmXdVCPgJ5FMUK6VQ5eVKwcKYS8muEaCaKBP3k9wya8xDvzE+
EQ8Hhq5wMCbbsa6vEQj64+VfHREfYWmxI1rw0pHYeTz87SGVKnItDVIiKubUAM97
+Njl226xsYHvlN4020uir83ba8jRoTTsbGBLBr1m/SIDYxXINdUcS8KY3crj1yM+
ehF0J8KDwF/Cv4XcDdUsOmfLBvFMME3qZQTskD3Ff4NctP4zmSlwtF8kWhSCF29m
SC/mUdjkj9Tnng8FX5OFOB6JHeDamGDPnBWwj5j3haWI+JOp+FdyNboYrrUcJFMM
FhSQRpy6K5JhPXju6w10dmoIbreoUJ1BoU6jNBjKE7LV7BhKB41n/10Uy0YtSVlO
MR1Y972NJR936i8mu7hClSNv2ieqsev0m/8wrFyEfvKAXhULeHooh1MM0q0saZ3Z
dB/8WwA60SJIC196zBLO2XSh+Ac4ZkjQL9oJEAecXMF3kCEVREBuUcX6ouyfZRT7
XccndCLM/EDiR7nOgeufv1ewpiz1n0V98mUbqz5IRYPIgCxocLH4+T3Swf2mLPNw
UiNzYCVxOC/i41sg7R+pMFltcatsz5yQBaOw1IPoc1/HT6oUEGZ0hs8VSSEI8U03
Ff3zdud1FkrkHOS0Dhlmqey5dYNpLH9xlYg8hOeBM5KS4WdK4EbLUypAIWzXEfPd
QqIZsnKZhUpQCHh9vjkea+wsx2GzwUEb68rZEy7ZB26noVwTEv/Ew8jL8U0bgSCP
Pe74chSeo7k78ozxpdNKSdSv9hxe6weGhQSV5wNloADBAd/F5PKYp8dBkcwX6MdT
3t0m69U2pG2fPckG4m3h21g3ql4d8OP+VnwoxUH4l0a/fqAga1rgD488x5KhCPk1
DAO3RPja9UDEiKXCIX+H3C+oX/XBWaByOFPhISPeJT9FcEAhOtmM6KFcMYdF0lLi
1TqMRycb3+dZwsiMFUDaCgrgTy4qvULAQ6hOZiGjHuPWA0esNCFcCXugyc3otnLU
HOTCbSobUVIo2SRZlKtixShXVoj7+Y6KfLiP20hraIVuG6GvGaiA0yNzs1QwDNGh
59+SmdUuwduU3uaBsTtfRnKiNA1/CJmAzZUwE5ccZCRg+DX1whmPQL9owZMbvvci
bn3MBvOixRqi35mos1oYcWdEHhtk7wunhF2p6XgENSMQGaGudt20Fsr0SVoYz3Ls
0RWrS3zqgETC2vqDKSEJan3ZhaQcN8ITpqoBLwbw1aaayP58YPIExirDY5RBA0ax
q3EY7XAzdRiiQKb5/56ZO+tqzo772LyNkKkEebhpkgrYgvFERD/YmBUAHCAZqa2+
TDXystalYRHolkbXiOeaq2JVJNVOB3Vylz2yD+4aRPiHLnasHRVrCZCm8j7j36nK
SxQ1DbGc8/m0MCOnHa6Op1jQjHP7IugfpVibj8vk2dKqETN8KVfTb+nzFzmSXasr
9ADf/11W80tzUvTTG0ootamewJ3ppIzgjGFVPny0r1LspnN3FZwxuuo1sQslPAbc
QI3x/OdaxgHl6FBd1Wb9Cjm3JKoqcOnGx9bySJsoFW6dkoIFaAwOc2F2OoBEP0bt
t7G+b64eNgeQJUFcmFeOItvqbZNFkKpi+HccnjWopj/l2SZrpcDbjC6JOIu9nhLm
KD2MOPsJtV2PFSHo12Qi1SltKU2kiSmJ2JePHIUhZYe4cAOxHT0S9qep729z2OK9
rO47EBWNV1vgMmBxFpD/DLlT5Zv1JwOib1iS6DrQZScI/WyMYniiVy2YqhMadd4W
u9aKnmv045Xk202tJRjbY8SXz6lewiRwJt+7l7PySeUgJrSYf3jXcXDYQpESsDbH
d0TNORrYuJEK5yO4c0gQFVSk1qpFdJ6KNNkBJTNRUY3cwvtBC+BHBZWD3ux760Ne
+X3HAYBkXI5Bzfo+X3+1wFvyNhEiqU1v49LZchwAYhGIGLf37fFxD/KdCERCKPSN
KXECiGJeCkAGIRIHJiC+p+wmQHu12lm5Z7Z9PvelnbtDiMWh/kG8xTZqQnxL1+ce
lAUu9wJqgzZvo3gkMBJ6gNg6w7btlZvreSia+sxHYJH+HiYIcbEphPyz9M+IFoWb
Lft9E7woLU4RfIRwmeLgBR8E2o+3MamqiLTdCTJwdpu0XSDwaLx4BPHJ+OAoeZOZ
0DvE4VD0nQU0ZqbZbQEzkRBrJZqZ7HFIPUPTnS1gS2BXEKt/Aiqzz6I+YT61vcIW
TMqX0OSkaGRHtPwrppTqR/aRAKcPpCZBW5kMVNP+K6BJ1OqaJP3oTAhYZrnzXsHQ
bDmKguFzsvqX0UxZmGKM0w5sgjXmyeQ3Zr8/bo47E/hzWmu1ByaBqhCD5ErjRCAt
bpF+gksF85a35yotfu+HcHim5J+DcG9XnfTzOA4QPvsL1jk7BMrWYV2cl6JdCw3c
1Umz5m2nmJDPKPLoU6omFBMBMuJni0bhIvqa3fxPrfgEsRkFLt14TRxpp2cvK3Z/
qsaCy63IDE9VEVA8D76DBag+LYhxJzhttz6GL7vduqsN4wElxof9b7/WGRhUuRMh
IpxyClN7NSaX7hWe+BLqIIqgQBiPnOI1F8J0PsCjK+1xhk200apW8JQ3nmZPuSDP
8GoV7HVaxXl0aIonYSLnWD/GESY7Q1iDnypwTln2CVdb+CX0Zdy5gpuiaAHVMxC0
1ksq2yUbanTVI3Jgx8eiUIndzKNmK1payriARocBZ5ja+hdm4OKGX5CUtFWfs5m9
RvwIwLQdJ4JUtwNxEdVbU8lARhvly/r7mclx+zLwOAV0Yxn4/pq1WVtVbOtwJCYI
5x2W1YMy8onitj8hrib1NiuScM4PIkEyD0wrXJ0ruYiAahfABZRIxMbuGNW/e9Xa
Wj/bVQsIgKBpjYhqN8UPwexmK9fvJWKr0rZ3XqiIFGxCHIXYp2pOsQEmUz1d51Aq
YLpHfHOqzi+wbCMB9T4PguIB9ENnbhGrXATwzBvF4UqF5brL6ntVoLb6YTmM9pJP
la0eNygXjpRFxAr4R88leD0UZki6TG6Vc6XNbQIoFIPkMjXcQaT9e1Fp8ShmFNa3
rbbqSz66MW6U7Rd8BFunHfvLgUgmS2NEsWBe4E/raaa5wPXqhwF84UrjrvhAhQrH
zdQysYT5so+9tWrKdqc5XhN/cUSaPOLQMXLW0Ohv1P1iyeImUJuZe5GUYl9klZD1
BH41DE8VmbRfsb6DPmS1XiZ73qGbyFyFL3xqud35vVUnye5sFl7J7B6oNWheDPXZ
A3daXRtPG1FBiWIOAw2efdk2quxeH0c13TOZSzonAOLAUeA3Fhp30eJ4ssVVTcT/
bm4Wac3WxXdTyUFgsbGDjmeUPLuoh/HLm/18jTIYefr1wA7FSYS0LpmK2ofBga2h
gTa4+p3nkBUOAjLGfmrg6HcCPNQg2ZDU4O3S7G1ILHtIfJM/TaBO2JUyQyP2d4dW
CcHhSfDp+nG2o/lXdgCeS4rH7Rir+KIwQUoFloe+nYNb7XD6/3JxZd43JdtamP4s
9VzBV3jNYyOdoUFBP/34f0JJ36THpqlIC2/JzhBQ+JXchcU9iv04wbuqI2/FnxqZ
jdi0Jppdv+Vr242n1cMhxSkkGkc7Qb76yWTwa7IMO9Dn3wYjHst1Guj1zUE5fY/U
TDeXkgHq0xIy2UeLxm2jjfi5GffpfaY+nu7mwRpuE+LYBLxX3iqD/pV1evRlcjDT
7rcqAm9ssy/YNrjWlT4kykFBCDzlli/dhtMQYcpwfc50DstGXvpAsQSB4vY9cR9Y
4yGBT3GOIOROVCR6Alz/pdqF5g12pU9TxETx8iBvmpkGs9yIn0SUKmx5YmzuKAW6
Hd3XQlCn6/mkf2oshRINetlvxafqmazvZFPF/hc0VpCcVoJcC9DcwrIPvHO6tGR6
D4O88qDCGIsdI2mawwUCfHFlBNbSc3KoGiHzCrNwNejBKCBHs9t/kUtGWVYOP6QK
jnUhpYBmu+Aix/K5nb/vfel3O8d6REhs183z7Bdy6jqGcvF+fLC03uWCMUD+xbd7
3LulxUUcqLbYbz1SGkBC7y8yHBCsBMLuyvDgWX6f3qg0SvUP/wRu1CizxBkTlHFI
XXJPZxxUL3HlgvCDyfhzUaShXoMYIEVrXEQx5m4wNhuBore5/A1krjUODix547ju
FBUTkiv6f52azioYgnS8a+7LmU4/8H01QqwqVvuNCZWAUPh9q2vOo+JsvyUimODX
qBAFByO2f1g09L23iiRnf4n7uhQUE7BQuqh+EZ8hkW0dXOu2Qe/bhO6SsKTj0SUU
V2jOgXquqArPB1NjInMpZ2CxJbeJ4LljBJinbpvNpzdMU47OawGVl/kTB+SNyjX3
2KB1uhaWEqAviX+Ax6mieQwSs1Fi7scLnwnL4VoNMF0/lrG0MxxmKPBZehxYlIN0
HARyZVU36tfc9XbJhQW87g1JkCtipeGfU7iEJGKgWn6m79taJkAitnhBRl5S1/BA
fJUtI2ld0nyzrVcLdcqumoxfZmLHFHnkbrzXwgsk2QzR3ywV59Smy+hd7osczEMa
NJyo8Q4ZwEOo6TFMmmRSnAHRt38SH7ijdJLS3S0ms0pmUP8uxi9ayRBKU3nUQ7Z0
NU496GvUCqv38P5zFptZaVTNkI7rYJ21v4VQy3xs4y9ZHJsX3+lUzytfc2OMMZ5k
O6Q8ip2tiiQDoOgSIqZAMRQn4siog7wxgUWotpMjwg4RfNIQbSPy5M4oiVeW4Va9
6gU0sqOcM6W63YeH9n72chNjB/7+Qwa8fpl0JCAnkoRCqkQi6mnXa4OplA9h8SpN
4PaU/GbVvaO5o3HprfbQ/9bTp9cUbat4Q3X765P13L0bD29GTEtkxBAG/BZ03JNg
1z+hCP2EmJ1WcoC5Mr65ckGX3+Z5MPaVIM4QkAbCjh9U4KOZ3dBmjfNhSMU5qn2E
1V2gLzP+lR2ykGJ6tVEmoXYbRYfuhETHd0hx33Jwi3N5fKv9FZ5nhBLwlqzZK8uG
+DCj+de3bXkgmjcF93xsKE72Tfp7I2UN7CDCkwXbSu1+IbGcrGZhZyJN2wDGEoyZ
gBfTuVfAuIlR6+zXMGP7tlRHjc5mBM8awYTb+NQWLJfAiS552Z1AEVtRzoIBTICs
hHjtGlROaiD0veoBR+cJ9FF3rjQng5tlawhZNYgCrIu7MWBe1ppXJDGNq/Pxdwih
cWSG2yutULbdMrxDHAZBbIJsF0+yKFca/dM/2gHpoEOs+bmWRfQhDMA/LJZJ/gmL
sw3Jt09KlTGmIgG5elufpLnL5CFQM6Wg/IGbGsE+rrW8XKyeoyizLuMrBHxm6phQ
1qvY36L6cgr5GZEpYg3OZjaw8qOLL6USgB4kTcy7dXrNlB1N2+7ho5muX0YaGxRx
52ogXn8FDlzAIThVOw+1P2F6tv+MLTIar03SEQxh4TuycKkM342gSIvmbmG0Acit
MeX9QuI7gdt+2B+sSU/LPmF3IjrtFuPaqalJBPtNpE2JETqSlrrMEsKwo1zee570
sUIvqcRuFiA2XuYC57Gc3SUj3lHLW9bYNnPLrdGQEvlxdhhAtfWWchV67rQCeTNe
DBR9iO2M/ePjyqnX348yXVVZl6bGcP2FE1Ph6BXq30BFASce0tdTglglUM1CIyeX
hh1OUiyeyd08wXoZX/Zum+sI28/u7nma6NJdSkZmSFueCNHEY15xWaqMQW64sOcM
qzL0B2OF5ssm+GfDQqXi78cqnBawN+5TON7rlRHYIp6fizogFQKm0pSJmwus8GjS
eCpDT/476MJG65+mfLr9i5Ltwyu4GbWY2UaF6XNrdlT16wUNKEcMEITVcDpLpjCk
AOPn2N/a83ffrB0u3zFION5RyeTs1zsI/+KtEQVSUHqcDgKlbyW0ujtO98iRVwmh
wVBh6y3ZIPEyVWK9arIJSCIMU7L5EYFXeGl9o4BxCGq+pz9uFz2hqyhWLryG4Dpl
X3mNFcCgUMHcG7yU8C7QwAHMjzhAZplO5W8GUx/xWX1JjVnV//zO3huu/Z2ZezuA
L4Ke7UYsOkG74+bxDpGcaDcD6L8KPedbDH59OPmDrxRUK+0eiv440rJT7LTFBSUu
/S6b6Mlh59mZUpX6rDeSX/baqluwa8cvqcIKECBu1TFxEa0WuoYKqJmOzN9keKno
17ig+/x/+u9ReikKEPK5cn4joDsyuqhrvEKyD6n6VUyPj/HM5UDnYZzPpAMV1xMB
RtC0TUz2j4UY8WNPvkq2my/5NtXaZ7sSaYmPOrPjIhfiHNzbJ0xtpLIt71sVnzi4
ywNupzuoJEYvJF03+TxqJD1U2ljzjV/y0bf1B7epo3AsPZ8XMBQoWBYHXyWYP0LL
qfWVtdirdEuqF/xdUElC8wRb7NX4/cokLW+t2jx3UvsD/AcS4lCyhHf0SDQKhAz/
BQ0ClQRh6iB0VFNmMH6reNDHZxBFAImui94ZXoFgtZVhDJsYK36voltA6pzpOcWy
N/t7XpGup+W4GFmb1p6UT4HJJB47z1neP4l/XhKX9yAiSCMXPEKc+wJ3T60iNJhC
CMFdP9FSOM9iYZG0sWNtM0msXtZPoI+XdzAeY7P2VbaaTpiicyB6m9Pewucjaqs7
VwcDheyTjQo0Z5QkAXPC2MlHW0HeVRzZkrItwHKtIItrdhObx5DxJ3aroLArz8uA
/jKqIeYZvNLG4z2U+KSoo5Y7G3ujx4tF0OVH7Es22qPo/py3KDD4LjNzq1EWke2U
jOsH94haAzj/mvQgU511DSrHL4rq8zIEDTdm+vuSYOxSK9JQotGs4t5Xpe0MbfkH
Sx63LF6p5ua2TAiyJXafhcrz22NScBFoN1a+32wtrgMuHyE7gArpyYjjo+b9Dk11
RqLMbAjjBT+iKkJcxFGcpBFClng34+lqWCkxu2DTQ6AUcayVHHSXkBiqzObE1RUZ
OUbQht8UcVGPruzziKohY7qLTzZXKumt1oG8kYil6S2JI86lVetBhVnS0AT6Qydu
rtaC/+Tzs7q4yHR+Yt0U/8lU7MWXbwz9+96WYggH/b7iMTqMY8D0mkQQtOuXzTc2
N5bp+Xbj+76ywVvlDhk+QtU42IrS0Xt9VXNJXhgUcs6XJm1kTHSXdt7ITjiAGOrx
q/66UDIsxHnnP2KbxlopgpyvIiifh0TZJ5SuDioDSrKbwxp57VD1jJCwO7MfBkPN
drOGQ5AwYKfSZWhdJZqdb3wy+6N4GBy1VvRswz/gxvB4XWBmdFY1UFBCs1YbLiRW
u5mzC/Htox2Mhum/7nvyfP1HnpWcZGkJ0nBE0cwvB6JU5U5aBdLqGewbxvHMF8MJ
htfZX25BiNQOLUeDzIaNqsuhvdFH6zQCw2qLksyNUDCQFvWxWzu50m0P9A59SLZG
4Dkmd4WfaQkwTNgCEN1DRdt3A+tjKAyArD1WhH2PdR4Ifl17on3Bycy3tcUfwBK6
pEeGAEbjDC9fQZbqMbhmCoYbPVIlJbuqbqObMEJ8qte8Kel6qf0FKXPhrz2FHcjz
gTmyYibj2BB5SVOxATS9G535WYqcwbRZWmhz2vfEvG4ltbecWldIPkD9fBnj9VKb
D+aHpFcbs1FvRwsUpHaD5UsFKXGMYJr25CJFKIfnsdEQG2/CG6VFD2dKByUcc21Q
ee7y7TJoBV+VBiegvGFC/tORApyObgXUDKSaltXIN35Dgl7rlYq/zi9fHANNTDkO
GVxidKzkU1tnt4b6CGl/XPvEXbCZwh7v85sj0VJL2QVn++hRDScsgp4krHltoaEC
Fz2/Umt5hJzM4FqwVdnnLLyAxj3N1IicXuz2e6cWBF+2wFG7ARvTP9KNOhk834HZ
BbUxP0uo9fQ516JepQdaWpr/NsWVUiTakpcdIg/02NFEYhIaeDSWDt6AcxrxTutX
M5BJ6c0qwtUVC+0fKKT/V0u/+HIkU/zpkrHf75AiP1k+rKi0/ldKjo906gY9VIc6
MFZudeJYBJ/3OkDkCrl6yytFaGcbCzSOaxOZlAI6hMfHjckQQ0XInDOqzmIIjj85
4UNYmh/5x0ZC7e5Z9tEa2UXdYjjOVsFUij2fugNVpwiByfIS7U9iegkPLTwN4k+s
qWzs18L54E37gLuO7aVcYJs9G9DXvBhbJqg1XIQnBRoWNaL+8xmu1xKFHGW5YkFx
uynvw4xexDitdD5o36fLXVnPU4EIqBb/n36vql4Oer1MwA9V0GiUWj4fvX8yfZNF
IKWPjWjkAyN89q9i3N5wgGp+e107wusvpZoNOe883setELWowpVk5kbnwY6+XFHD
WcYIOLol0e/3VRuHM+wx8mD/+e3nLcnXNWgZCtlHPAmNDfpWUSELSLrF8WfiuPc3
APDAc8hJhSR5kNzHU8tDK8xTRiXWmwz4LjvC8EWg3a9P7jsZIq3Hbvo5zhW0nuJ1
8WQBIwZiF9IMCTkJZJITrgglmjjUlC9N4UVw30xCP8v3BoXL1e4EcDFJ6F9apGfl
33qrazAXO9ArQA5POo1+KtK4WcxI8AMrOawibtlJDTAcDtmoC7a9kUcxclfXiiKA
+/MOqqeu3XKmIG//q/Z5ZWtXWIWvI+kQPBz7OEp3KljE6GjVi7tLnXvuRrtoSQtu
Y3HCUKMJNaEvILFp6xnv1e+q+JQrFOHxAYKWNOqOy7CWZqocgeu9HVJaMbT/qz/C
aJ4rED0qAEd82YOKG/dnqWNalRNTeXZIAIh/vximQNjPHbSXczK57Kbmu8+jAeVI
u4VBVF1yWew7aUMqtNzVIUU4nXThKdgEoBWv0yW1Ka2MzfW828DAKjqeiSY9J7qF
Ll5wG71h1Uozbeyhva71DdPFMgK2wjdS/92O+i1R/q1z2hYyWJW/67fs5mCFUfwW
thYJ51syRjY/gRysUwa9/r4TyucrZEDWhQgPqOnPyU6oMb+0U7ukuhHFW5kfD91p
M2HAlFOTNVMpOOcFcz+XWem365s83Y3DcS2qXtMMEKrkZBAUDYSZScleA8FuV61P
qBeWEtqXRhG7tQI5s2+9Bt6yRVMWt7Zfy43y9Y4zP7wQ+0SyiMR2JUWP7Ae4R92I
KowV01MWQeP9ey3/AGOJuWIaTm2Y+3slvxL2vYzQ3+cNzBoQy8hZuFn2E/wUNYiJ
w18KeWKb5jjf9SOEosQ5YbdkVR9UpK+FEPfCooCmnWNKbWpauC3hFcHq6ct52xQp
ZYiDr0ifWDQPXkLgHYNpLOXGsYB68WphTKu7y4giV9CPHE6m4m+A7YZvKmRMLasW
HJkiu2uZA0qVYfEUqNs7LSOo+2/mRrp7IvdTuIakFvGAG5gUbWyIu4jya9Pvb/nQ
2Pf6WvMx1GkbcNvorAlaMTxBI5KYBeEERRqSC69UFgOoCB8LyzsX+/AXD5v5IquR
f7XSbbbeg+7CYNnmxabf8yKd1XcynOKSu+flRAi1t/YVhOAaCX+kSMY2afgS/SR0
BWq5GpPwIajYwz/X97K7IKXLErp26gvoUk44S+yo7yvdtwOU/ND6Gvdn9ir03W+e
kAgmLkCNMGVePHtaDryPSsSbf5GtQv67lRSGR3EYSw2ZrmUA4kb17GNBlF+28qrM
RtAG0MrhF2X3I5XkGTQJml+D5QRCYOT5Uk4DEf8ISJxUCfPkMWBM+/err8t5HyTM
5WCdSr2Y7cQlE21XhHUO1vM3aoVwWX0xW86YzpRpZX+GqNgAKc/LqxmR1RnijceD
4rDLmtQ5wpL3ZznfKh2WO29Zq83FhatbC/Pg4GZPjfxcnp2Kg6BPnnhoObBE47Ef
71nnUPvpz7NK1+4HnSo7gfmS6p4ki4+Du5RJrZ527ZuLfJa0nl4JCRRoYYLOZ6aW
HgnOH2Dzw64+wV3pIgTKog85Gfg3iiQ0RWH/yymbZyDkksPVJn8zo83p0YanzAWB
WgltvSVdN6aNSPTSvmMEDuUhAlymUgLyE3nMJB2F3J42sM/fSwnPrvJml9MQMQoJ
BeCFZ70Ge2xxQN+Ra3y33nrct1cvBH+ZOL6K/wmjLg9W261MpXD2zPkLIXDLINmo
/8OdrGQpPX5es+3kasRqeqeRYV9ylGomEGQ9oMMqce3LnWpC+vcxgsvZYr0QW24q
DOfokIj83CrslG1x3mJ/IYRhrC/wz2+Qk6M5qJdzaQlcxuwcy6SI5Bih5fVeQm+l
B16/54Zka/HdTMX0WcDisK3LCZYT4rwPKGiTYjN0kKEuLBvHoYrSFtq9CB7QXepJ
D52+wf5e0wiswrNfqkGA8glj+JDxudf+4WkTFaz59iW6bQAcdqckZr7gHi+hClKX
fpMxvccM1qK+4XPDv+fAyEHuKlxPO/LOkpSdk+K6hzpQK8d/UG4HTzjbvQW3xaYa
vr3yj70v8QwJfZ8CasFiTRn+UWZK/D6pWcnc+onx63Wo8IpN4jSM5sibsep5UxjB
JbAWaxuFdDoxkRJLt3g7QbB4LnGqzBooTgRNdYKUYoj4WwKWNQvpGg5Jk09GxDIM
yt7kOFi5GANy7ndEnABmBw2BmjAeeYYBjVu/yyMS8Aq2PAMmfDLIETKnBZWEuarv
qwMyUfcVAuUSxZUxs/mtd9BcSxRKa9NdeK1YKjpGnwQydML2tBZBChhZqDVY2h4O
ftm5+xVanK3Lb0D/3kImAjvgr0kjROGJ74do+FuarEYwnOHFZFXkj//3Aov7ccCV
WVOb6N4N5hFJSYLa+mGxdwUxHlFjzQ+WFPrZr7RqffdljX3YAjuWb80h/Gh49R94
SetJzektRMu84u4WoOepaC1LRtV3gefw6Kz5nJNRpLbXkP+SgLEjHw9cMu0SJzlb
HYvAMPMJzxu9YfRiNaRl1gG1cZabmBHbEKJUT7tQ+SiCEqe1RU2B88ar8OwcEDQM
NIoFobY9PyJd1TmgQAzP8yQn2ZGbbSZ7h/c0uaTQ53mlL2rjcsp3rBhaayhAvJ1T
3Qasp3IsqMRr/ZhWlJD2BEEcdVA6xO7yb1egpXD01e6wvoi+LkpXszsZTxlkw9PJ
vZppv4O20chPxypQlWO52Va4cZFMdX+ij4mSrmAh7+Xq4RSJcY7/IyYRRe1WdfvS
9NbSMWcwrhMzTiU02/OfzQ3HBMoInc3BIHYL1Ayn5CkAqNGOyOSE07OyruIaK9Uj
0bCfKLuQm0SElhvqMl0Oezsf+/dtTdslTiEZLV1Um9EfFC6KiI+FuLHU0TUwsAmL
5DyBoUMzuNWqaXnngzjRCOOHCDNBk3O4rqHKWKmoQbR6VmbL6xlnw36u8amxZQ35
gGfKO/SaHavIc22DJWcuXR/VbDFRPVq1OP8ERNfj9JT0WB4u9OermHiMWIP688mG
9BvP16nJ7ENotR+FCjfstBtiGLRU/kTUG7No6kExgFbxwlpcfZrqAgzdMJPmD1Vy
+82gOsqziLe5K+RBWc7w/n8HZpLTYHhGlI0stQI4kHwrK47X5QKK1cSFZj64uWQF
/Pe7CHMNsyebWC89bDuunhsqrvBrm3Xuvcjqhru+uAONb0JrroQwJUI6cF9MdCwe
6QGpP7jvNGv3gaEMW1aRaYHJcDsq6R2tLeXGSmarZlE36bori7OCAUsGNG+xiW+7
upoa1CsMNy7Rxu6+b7V+Pu/r2IGzNvMTeGbxkz4PrhlpMWDFVuNFpfLeo19PKBIL
LXL5tPLdZwmzokQeZgAWvkWuXa+pEtZSy+eRy1h0ViRADsKlQ9AxmSS8/D4t51GO
rJtz22t+UMuYV5w/7Sq2lvbCneVSPl5PsNeMwj+5nF3t00plGS4UJHvMdXcqHQkr
4Cky/ZAouHOKcLh7lq/Jse54JReNOPdyQecowyqbq2wDLzCFOnzxy6tRD7GgxfjO
8S4SsXJzTFq06omWSChjLHTxmbSJAecf2a+s3N4SvajYQ6RglSMyKi5aTM9TXQnn
ks5tdI1NRc4oGq64wUdjJodwzwiZjEOGJJ+Xpv2nlYJHzIWstuhEzqlnYwiTa13M
YKLaMZoEsHDq79d06q2xmZc7wilRkg/AYj9LOEe52sIZvjX69F0x6TTkDcIx3NML
jAT03/JjoeBvgJWNlZr+7Q3l8sbfk2Mlqv+Y6fmx/D2/y2pNluMVPsYKxa2wJ/xt
EYm8+dDJ43wO+GoVjzZRUOrjcsN1fzcmQZLD6xT4Zhd7BZlSb7yP72hp4cIthDig
GPDf19y02VFX+6JM6bGZ0a5OKlTFe+5B7FyMhPAwNMMIfDKUmgjzbm+nuvklj/bp
5YqhVCp9I34zltcB8FAnvGrJ50ve+Y4D1m+LwFwPuXJQdpTjkcDe/DNPkCRtIpl7
DH8f5t2xOGtjo5ilI0gAa+VQ6WuYFCj2nxQHufEk+6A6Bka3M4Y6P8NoS2OO1qsR
yRnmABRIycLleiD3lxWN2L0KomR6xlGa4+SDyZ/RWLhh+SsEVoSTdCf9vgAV57WK
09YVzq1L9CWzjV8Yqk88diU3moV99tMpeNdhOHJ5DKNQ3Sbhrchg7mUSI9To04nL
KNhvj2cFMKTJL+KoZp33f4nuGuqX0clYe+dvoGWX9P2Lx0+cgoGswrwQcw1UL49p
UNs0fWwDYF3yh1a+l8iTN6Zb+qMEvrqJfAwHoJm4r85qMy1prCXMm953ImTLFCd8
NhlFk983ANPGCDpMIg7ekeQ+S6vILOq7E8TuUvTBKqAH7RTJJLouyh0YBFpM59/X
b87+Vj0HkL/nr/bOdNx+qAJhlaWxp3aqrApJ/UHirSXQnwfCMkFlg4BCDNqPxfHh
TViDow53cks9pf/ndrbMrpPNMXcxIa9Y3shjzjxHXXQkDRLBaq0XvxRX6diECzhJ
jZ3wIu+9Wz7IbYfKyPXfZGgRWploBLeIm2ieICUneDoR8f1t2HlMWoU0XmS6yRxf
NufH1EYU5Hf1xeD3j3hNG+uzTj2aCCL9B5mUCDtTa/4cpLodIe9obmjSsrhhmSNr
BJm2Eb25EZ+Rr7pGeF/517hrthwCrBqoxZn2n75Mi0O0u97Q7UMHLFswRPmnLbeV
xzyA9LHFyk9H1/dU9QaDOccyfCprTTCew4ApxLgGSBVXm9qCTAn7ykvZ8blEwJv2
9aezdKPRmpk/xWR96hiXomSoGcSlqzBMtHr4bt7b/1qlYuzGTBKSSoST1yDPlrfE
NSVAkGMcG704RwdaAo6NzqaAhKSqvkd4y9opzwSg7pWsN6Od8GwYN0C82KsU8Ld1
po3OHtmjjorU6m7LtO37I3hjALrflL7KuObnIHfc4stHBF8wFIrIs5cPzlvOhHRB
zEYaOAHLFDfOwhH+DSSuie5jl4tvoxz7rbf9vini6J4UbxvqX//QqsKLEL5eUtyC
NdH0cTOHRHh/jAZoX2QuwL0qSuWmFDFzonFtxgGVa/FNJsGTJIltCxyw6/oaPdch
67BI4YXXKzNvJh6LlePBtZhkJJJfYnNEH3a9he+l4cL9p/vHNAbDpxkYhHrkb7nF
GjRRvI+xvwkMoLfIV0O/zUXtDjA7zZQPVZ06qRIPXCYKxhHQg+a8ovAN5FGL79Bh
P8vaF21FHgDjsKVk7osdmIWVz3+0OcOnQSRoKJZZPorJsJC9Rysz0kuPQsw/LPr2
/L5ax8u/EyhFEvioqOFqiauweHOhP8MLTqCwOdsqmfVLcxL8EBj0W63HTTLRxgAK
4d0hxP0DTqbni11SECmzr5huIN+X/x1VT3DRRPRos4CSK5QgZE7UBjhHxRtyoKgp
KxsbGRw5ijYF5QwtielHqNt3VRheMLh9m2oqZlqx5xPJ+yKSROQ4Bx4obnM4cwbK
KBeIlRm/OHbvi6X8p7uM4orUKl7JBH8VuZihLrjoo/WKZDC0/gfUQIQiRo3Bl9ny
MlBoYaivs+2k2YOev727LHV+xc5a1tDsG5sioXskq6eTWKA1nd7OnJ95AykspcWH
+VHNGOFxGARqezjEfVrZFigBlY9OeWU+lBfqjJVa47f8U5f3sevafuY6zbaRCRtP
cL6kWBXJkg337UeBl8hVPakB7Uz6xe6YFe3t3llthCpUlWfPvcxG+iXrO3E28Om6
QpcBXAkFjHW0wmdV3P/UhJv7g6VTx8zFsQlAhdeA72C4o88G4lAZi5q+pVFVED4c
O3D++fV2QsoBpAg7sJT/FrtlpqAkdCBSNzsnFTtpoaNgassi1VqSMTKQbfpAinc3
kjrv/yeAmVpaYp7kfrJaDp5FtKqFVPV8upQBjQW2UhbaMkSLURvKAr39sJXrRzoL
D9QwEYCYtHqrQoPY6qGIhVToIez7hrkbuI3EkpVRQqc9drZaRRkBsjkIkhw5x8v8
0zch542OR2UmFR/MCsvlhLDtYVNwTzcz5K1quA2ssq2wtxQvwz1GZSpll8gkDd7o
rQhSMHgMCy0mMDRUXfayhh7ppnWdxp8jS+4Hn1N1wuzAVDZNXAuQAE3kJ0dB/nRO
FIOoqCnEEH030OvrlMUslWJ1rv4376PUBLj7P7DpI6k7F6NEJ3ozqaFVjM1Mg1jA
AG9psVXUkSdk75rY4qCprS2j36KwhO8npX843Q2YZarX1JC0zilTVbud/hAn3Vuq
O895i955nT9Jv5lUdpUJRgvB3YaFxa8uy9r7esy9HnXA3/BjAAp6LHJ7V362ggEG
JymLO54G3LWhiE1pVoiWrUe3VBis+6ohMAwe3AKFfyDVGAI7+jw6A7GI8B/1k7OO
nLYcN7iHwy2qgN60fbCJVeN0zecchrvvp4KukkhCukHeoIbxMHPGydNWE160zAVG
p252QuGXDxftZYi5RbVVrTLMp8DmveC1G19SiVyv9bdbM42w7O9CekTbADKv8mCG
AiXgzPPLlPiteLW55pfitjcZ7EE6EFpTkgtf85g5ctQhTsx39fw3rjKRKjBh2xJD
llBBwP3AfIfSXvXepRKZlwZPzWvQPx/YFvWiqiGrIQnm+o+inQgti9HhdsSkrbau
XlxYvX5WtLFagLH1ZsdWVTzW5xvULkZv8dB3BTn3SLKF/UwRuz2bNjgnN6DRyLE+
ZfsUOa7cCUUczddmJmf1GOv1kZVnRzjiVpP4Ml6PFQbjcZDqjej+OLjWbxIIfgiX
9UxB2QcP+nVPxJIBabHZjsszRcoCO1jAK389BGiTW+zQODINL82Tcl325pFY5KOM
7AHx1kOHa04w2JnE2sS9e4yRPnkIEfu4s2mOHhzWKm+NYgYPWH0EdpEXz/9HuoGA
jpYvH+KhfKkR0iKZ1l7GePgzlCrj2WLkbRlcOz9rZD0LAuYeEOJoiiDF7nVg9pSn
+yJ/kOI/9T1DjNBq6lE5/H49fJWHGMq1T961r5A5BYiSr0AmmWsoJv0ughEvx9AF
SRagZB/qG3L3+GiOcrG9YSgt8CtO77t4i0mLO/Vn6YpbjiTrWIXKpzGeMaaz9zra
gMQft+1P7dj34qCIjcohOEnnjji5PboGZmVmZO56Vs8jGvip+0+IpgNxJadyehFY
b8pW2HnSdZilfeETQFeS17iQGn+NxmNRfCHs/h18Gzdv9nZgMZEMtVrgCEA/jXZh
dHoiO8pHki0Tgd2iL8r7Y3eDN4AiZQ12xGYneDr/Al1l416lzHMdgQ5FzpNZ8wez
NN0god1edL6Dk0BqL2gCu22iWkkTy8h3IVTPOWZOVzm7ORp7bDf31rgBHCkQ0fNQ
1W5aXCnwWwHIILN3vDeNg0WWa9W7+17x+YaFs084E5Wo0F7vqVlliTQ/Zr9Ln+Oj
DYlLi1tj+P1U8saLjHZFr9mMUxkzOmW/Ho7HjAkokz2liyM0y/xWp5XXkj2tp7fL
/gN/OXSXoCyz4pGKVnMmeK8njHDDlhKPjyd0oMHiCpd0wQfK+5+P+WpoG5Ygfw43
96zICE4KUvWOk+ttWON7IYdmDxtm1MUj0DXzAAvufeFGYvPVNUjifd0YMcDHeCvf
K8482lToI99YjeEk+G/EL+fXUkE6BOMu8vPIwtxXsYLWN9YWjx0Cxvbaa5iwend4
dgH9ZbLKc3lSAx6oTNH80lAjekIyuF1gNPqWeCXvIw90VIy1z20sj1fwJ1ISIcya
TsysMZzz8Mfo3L3l0BARorzIOtWWlb6Demy5G3z38nCTLHxyADOnvZdsDTqDBb4R
jBOsjZgbfhkt5GaHriYVzCJ0n/zn38r1ORcSne9XamHBuQLhjjIq9gLwpOByZf2W
m1M9YnLLMffX/pTRXun223U58wRMNYmFVkcE54+S1tCm4v0i+kY6D15SFqq1cO2Y
JtfSrRqNGvJkcq3ca3/qwBBE3ofTx/TDqSFTlq3EUY8U7Qq0RxMODeu0BlECCz25
TCUUqDZQGApUnFcsmQxHLe4FEOM925QOyRTxnFxa/4WG0srMnTKAt0MrRSMxN6Ga
Q7KgeSrLcoIozEKjEvKn2ypCLdeWUChIuvWXnUIKnRLCtjmmTtQtJWIpualhj6cc
q2GL6s/hUNPzQDxP9kmuU7+y0cACikJu/aBEIilqH2t3aGydvuVGgN1nJJy4RgP4
Ar7JHXR1bZHDOKBVrXSwERX1VolJo5/uNSudTwDzM3vbOshPQ/YhB5rl5JgmoGlC
kQdNvcYA2oQnkE0izVjA71u/DBhfRYl+BHsRHTHHb9fqn0LMlCMCjMEM2wLtDotl
Ag05ahbor7Lipo7O/c3y0rgzeNrMlaAj0fByTQhyhBzY2iqf0231usGqZ6l9GRqN
vIeRq1whjOY2lZe5e2s5NRr21gij+wfEj/JaReU1Y+iSsAzteS34LcKU5sojw0l+
2RK0UauVU5YveRWjzJaKXJk4tDWSMD+c4zeoWMKZfzyxfDAfl6nX8eEXnNOIPaWC
hfrgFqfYNm2Fmii3O3xx9AgDzb8/fcIzej6OYACY8KxUibaKhDWgSwmT4AHDIQnY
UbYgkrgGvdgTJYwSm4FPqbxQP4jzdgRbCZd2vSSNXgwLyfYpUXysP0Y62udYJ1Al
3tFBUwx5G78ht4hePaBseDlNnTp/jatTDBAU+Lf5LVKEFEXyzg125NrLhBKBpeKK
4NEy1kFhbp9grx5pLM5rP26uCPlgHFkeKpwpCeltIh19Aqh55XFcuhuEQh3mLh9c
dJOMqyq6zEyGCO+r4ZadhGwwioTARdaILmHJKxeKAEe6m2r8apl8t/P4tRAgJKS1
zH+Dz9eqr9c2hbm/dowqAw9SgMUg3o7Dv+rFv6Y6Y3K2Hr1T1pgAjVrt3zFDzZ//
mgbCtXA0I8BtHZ4zAuxX+zRtnAmLU4GvRpBHCjOxJ9acm0Gy3btO3LvuqQQaDUIW
Q2JSVcQvo07TaWPqyisivahkQrBKmotg2HxmnbuBisCrI/ddH6r5A8VW56g1/ScH
QC10ICiI/MsNqYUWUFlpKEHwPAba2BdhpRfVYrMVeIaKEX80Q4I9t6AbSVwj0w7B
SIqlMEIXomgakhH5ItniJAGB2laiirVt5PtxoKpWdcvWHcg4dUdEe1qcVkcZGVXa
SC9iFkVdEypNiBAKvqKsAZObdYsR/XyWqfhfYk0OvUCyWHQWYFKDW6CQrrZgvs+I
Qywl+itSsxzJDECKbs3Bwnve2CH0f+dkq3VHGcpQJzLUnhVjWyFqnJGErH7oNGLL
mgrgM1jMAykGk4JDsIck68rMNv9u23OsWsRlcW9b7wOeQK0W5cs4pDQtUgXLoAPW
peMzJEnCvZzNOGuJV012deiOQZMPbGVGLU4gBNY79qfHOE81LqQlgedtM2DPP84a
MUOx3G4poMXOGPq++uEY6tUkr/PCM9ZDSNrq0MPfdnoeos/sbnEFuKFR9Bbtxvry
TSRA1d7ukXQPrEnQP5wcz+BYgqs3uKN2w54oMIddlfc1dNzf9ezQrCg58tSCIU5N
I0J/YCSh93svd8p0nGyDz6ALCq+n+IVTdX/jFOrxuJ7m1RJvf5CIs0xFsyrNObx0
NyJFbnPIyLmApH8v6U0s/0ildEr6WWNfSey8CqRPKrCKHTPWPjqS8DmRajeXSQI1
+DfmPVKdGKlqryqgLbw48hYH5eT9LgcdkLyvBGjBQkKI5Pav0Zzt/5PeUi+zOq6e
gTIFWE9uTi0Yglc+auU1Z/wLki5c++U9q9GMr78HDIlg0L5tOZ3lvjene+EX/ljy
aRy2Tlw6+QvjN3F5aUXxL/Foiz1qYuUYctdZyBVaT0zoU6ApXeilgEiR2RzEm2Js
i3vXM9G/T3X5u7rbxAVSqoLo4eRBapJmBBLa05Ts1I2BNX+lfImoGCftNdbP1wbw
NNoUHXhmRY8LjSC8/MtN64+wBy0VCitV2G2drXIb5t5djnBEG9nh5MbO+fIgNsAQ
tNLOVXBmBbZgQhJAPvFfhHWLZARGXPzJbuOzjPvpDLUqT9HiRZLERlfiC5Q3ibWe
sxztkEcxo1dcRtAkIZm88zSDeEAtdszB8k6u/9RgOVp/05idxY4whFBViFyB9gjG
cTkfyxia+yLiQ0TdKq/Mdkn1QnkfWsyl+zIVN+IKC6kbV7S6oVeqOBvgluV9CJ/I
F0RnWuSh4xxK63GRJB2cAunN7fbmu9zBAigaFCn24KFUCLGzb2k1ypNjNpAjIvww
NiL9RrYIUYuvHYq8RsmN+aK376Oag6NA4OvFZFWYg0wXHXizBv+CIAXlWAofn+Xe
0FFls9KRaaaM5bX0TaEwzs9RjQyO3sAnqc+kqzSWUJIhocrv6Sq2/31y3WNyfjGm
PRA/CO6Hk0VnvtVZmibNM2lAinZdCydrf77H3gDgDExNtA9viwsz0/ssc9mpEznP
zIw5KrVlmPlU1h6FvoKAGfK/0jJL9Et0vgNBYsPDN01hY88zGlYr6wQWvyw/k70M
QTX/hGg+uF6MWv4QeVMHW1idf80/UGHYzotk2JzkuGAGKs2T4PnBW53lZH0HLrPJ
eQhK9iaEJEvDoaabSkbTKEt2G8EiLIDBPxyPeju9R+MKHc9c9fORqG2yPwnl1dFU
+M2d6fK+y1tMuP43Uc+oIBFL83QysQCDfewY4UODV+n8iLeKpIbxTC94F8txDKsp
G4295MS8+wCV9eHoNNc8ASM6qpUP2PAbXBSjrqnnwrWGqS3D0tyM7l9GxWXniibg
UEMEdF8yjkErmTPmlaG6Qq3mAgIsBeNI29LuIacFK1QqtdSiWLSLdSZdEihBGWZh
PGimDBEvRHRMDume+w1Lb698XeSPwq31mx5mC9UTcjYY9arYTHV19AKYJRWVXAeM
/eOSTkZmtaNX8igNLFz1AaHGtAPLTiSlYc0K8+Y9V3i/n9GivBPGwmgG+rxYK+k9
Gc8/IbUXC5Q52U1uSXcSC3zDvvlG1AKHm2xSZtYh0lzmlTodH2HhoY3LUZ40CAX6
DTYra5RK1HUrH/RGBWzINTp6mRSLJU2lLGeSsl5O1zBC6r1jmwARyVAnzmPnsq9G
auVFDwt4O6CeRhHXkt5oAWztWpx2nhY3OgoYH/bnYuSKFjVGtU4X7S32du0XF0vG
Th4d0MNVlMMa/nukSrgcLUpn0L5Ag+a7LXwrD+jNlsqZyChNnNGT9QMRbcrsX0Ia
sbeA6QxQivLD8R9gi7l3X5EXjngd5FL5Js9Jsy2oPGHXWNtu7a8b/qXqWMcEZIg5
jFNR06AvQq3lYgOtvdkePhPrmbCYsjtZvc9uQNsiFuawPOdvN3xCzUkQy+Tou1Vd
Q+l/PzAAitDbIH45a3YjhvN5baWSGHFcwY7AY8mIipOHjg9ALYFO6izMNOqkSyVw
WfWq8qc6Ir0SWHCrjXS7S/SQBnH5Jr5GWMvv8x0/xKUdHW1Cb0QLeRHm5PxlE9WZ
Zh/qnDz8ZNZMXfb1Rx5vgeCKCZP5EpCyTi1sa58JyMUAZBqlmgZ5Bd0o3IPS/4RN
MBqWxorIuOFhtHFhRH9U6PRCjKR+G1/6ehkNSvw0tiSu6DtzOD5N0iXLbN8VDlML
0LbgQbnzXHt+0a0PNvxe/p6zazywUZpb2/xNLuMjaEIVEoeaaL/1LFUpDHigEn1V
YyhHLDeWBj2+BRIVAgvRKCI50AESRLs1C5hVIrlqwp0rOCBZ32KK2Ft1n082kkbl
qg8pjo6jZv5tiPMsv8s/cIbgc+VWVJKa5Lq4l31KcnqEnLKesbwAvA6k1o8gf8If
V0ocDAVX5pYCdTkT/uIL170WA2yPsvEE0W4GF0XR7WcjAwB0DrV4MpvmZAZzyC00
vaEAzzsYVbObnxwwBAByXDi0IzGWRDFXDq867Gn1vIAFkT+dzLVguPyCJpGbZ8C/
rKzKhW9uj5UJSoIVZICFfrgENxDmTMfdPoFjgh+MChbFhI5ZuioNFi2YBC4FY+fQ
g1M/caO4hwvvkRbUI5vr1u32WSbq1kkagWWQVkF8m/zWE3KPQQsm4jQ9C7BDo6np
hQqChCkdkbTthkKTuRHL4xTCfNsCi8nH3OFY0C8jkjGIk9MyAZXdf7oQ9njK4cSG
yQhYok7xP9l3iodOJEGn+w9XRHPb2pEnj80O0fmICSLqitwt/8pNMgJhJEmqauAp
D3dspF972a+TLLn2XE2TWOH1G7tEFUQK+g0qasrGNx6IGXHUL+B0G0BoxTPVHm+u
saOiWa3UYW0OZpzrAhJRjk/sTRck0q0rtX0bcDOY8vnFE9OjTlBCadMXsXZbVyBF
rJwvlARj++Nvd7I8eiV70E92CpuFWrPkskftXpLTp5CAvhwLDJDZRNopgXIwd/vX
zKRh+YJO+QMnY2dd3054MPlIwlV4Iaq6WByfUuAVIMG0c4MxHayWPviF6GBUYTOj
B25gDvlQg36akCWD67wS+Vq9tO9g17hBsMDpksuwxPkezZeMSjdSeVGDzhNcOulc
VUtT3IGe1w3Cs2xWSVaCEupuixI4CuFPLivWpqblQNRUTYmyP6HEMmp7XimAatXX
FoaXh9/CEiIXgGSsXcm+OITVjAF+0zQwOyQPitIySBhEaFmYXuiBUuTKKL/+seE8
DJztAeGm3htCxQb9PAwIc3BFMZmTfMRkhKC/HkE5fy1QMa4U8svkIeo2jgKdf6oh
pAP+KmfkqfHBAL8FzQTCpvsIuTyeb0HuFHnuwRQEhF4d/UmGMNEphtnBEKAlQ6f6
miKqyOTwAHRAWlsLJLlMWV2ZkeBsVRGP7V4GIvUCm9yE4yAgHqn7jtach5TzpJyb
tNnciQlsBoDROTJpME6OvF/o429kKip5SL2RbNAiT3TaYP8HhIgMMF9cPfaTEKL6
EGeqj2FsaCP+jo6X7NDubYZCTD1bmOxfqK6+APCvg2PdCDGOK/SqJWlEQk7TDi5t
QIjQ/PcoVmR4hH48lULfplT3xkEqCct0/OWREh8NoiQuxIFROnjWTvj9/hfb/2uC
G5WTzgRGr60mq2lNkADoDwK+CFD1+q5TQV/qijyC3lhXyw55akPPnLIEV3J75BpW
BRFojRwVj9hQgJzibtOZLHKGTYp6qpCDJSHY9BNBCms1YHXgti2zafRuAcTvB+bF
rLaUJj0JOvnCsgK057tbLgIDxRsZm9CiOz1IwkQVN4qs2S94weZveSp/xVW+FKca
Tck+bzpLzHfrAFL6YgquIC/l+pa1I/SudQa2fSQOhK1TikdYCcKZgrzgpEAdvVcM
K93F5QeSuyThgzH7kGmZU2vAiQZILiyx51B85snrOt63z/YOkN7SYmyG00xXXgq6
Ll4v20X+STXgq8kRY2E1dwgLWNFJYzLxYe9o3kjq+JX6mgQEsacJWlbUfeRJDmB3
Mindu1MiBQrfGb3N7sanibRaZkcENXAH4DgHf9B+2XYFP/kP3syBEMSUBJ035mRL
k02s5wzhIv+IjW2UnC2LzmiO5wSckaot4MQMtN4mb0bMPjmag/JF4MZd8FIuvhXY
2awT4wl0YnJXfyA1w3cz1/LIaJ8dgXy64LQTeLF4iEZnsopwbClOpAysRqS2h4XK
hAWzoLvpx6NPNWWnE+Q27yhNYFujqgko2rKuXBkcIsCiF4yPUqZoxmb6YFtUV0vN
+uSfPZh/5jJDmGLv/dm07R1aeFMKflWvdH2ONtVjnDGIZ5LR0k/bXAALKRuPH6DV
vEwoDAfEz3Oh0FUybqjpG4hVYbpoxLa7zW5vxul6tPdQ+h2gdnXDD/0jrnkfYy5z
7x62ygH4OvtwzFdXo/ZA9K5zBaVu5/PZCdC5kU/rRr3yBiak9kn03KfU02uvZLHE
/7uKytYYLEX/s2iy5E6RAl9BemSGXFog1p7uKjUZtFNUocEePOQGshWWQkZStKFI
gW0YhlYRG/bz3zYWAZflJpR2ebZuZvz/aCq5voF6PgmOYQmXDeJUzR9wJch/wqWY
Pks3URscmDu1cjtW+dMdFLkXSnNdguDGPoPVoNgI3/+loxQK+xtQ5/POVDBRmhjo
F6LvPdPK1GfH7ZtWVhVy3TGZQ7bx+NhnD12eg1ozr/3tjCSKQSl7DZxTS59FCSHe
jcJOB9aEdq6P/n+AFnu5dGjerbDC9bDp4ex8nk2nf842r0qEvGW2Oe9OlbDIbVn6
tJG1iSV5qxmuVzTUKGrIYWx8nRxIVnHP4AMwVJsBCLvg2mg5F2EwQm+km2HNIj/m
5JNXF+/HioslqeMzrFlQbtRvJm++EYJUSOYS+mQdimlG4f4zuWINV6F7/wNs1JWY
wgKMKRacNR5hzdsolcSRhUlP0+LE7esCST1pGoCA1CfYL5p8IGqoQYiSui9s/ump
RL3wCP3EhvLwXw4a1OrYQdkYlZIt/icImvl2AwcwwJlTUR00gIF1FpgDm6zvsDUG
YUnHVZezvvZmya3xX+n7clLClqcHBpTDTESQ6BR9Eutp0iUMwSvPoiJ+oXPG08kT
cF+44XPkRqjlb4zYU0GM8oJ1aWfWru7aiiim10E3BnJJ395ELalcM0ci7FxGhqdv
45tcf3qTq7CqvTMbQlcRYFepWzx5x5ZcyPhpYyZIrETc2PCjm8iNBA1o0CA9d76g
HvSxn0n/ZXemIp34FwvJBKm9SrTA0zfS3JmpafWhvRkhtflMCMEtZb3qYBrSL24z
/DStGOopm6drc5zY8ga0cnC9oq5RTlxHkKqLcBYpazLXJ1PelJxxlaRUiv/TyXMg
c1Baqk2/tvPFYg+kFGcJ6xVatFflvYH89nRoHSpzHa967Mya/futLamsHcCzGiGI
LZuM5ZEzvfSNbvFbhRQSQYsnI34SluCfT4NIL+CTJ7obs4KnoYid7CtOuRbrTz/g
kZVWZrFe+P3Ko6kRMi83gR2QZ8OPbZcn53fBIAG4dtkeJayLTla9xBg3a6fLzSzQ
MFXmnOFfVwZWjbmUCqtcjxQRhy4QAWuo8Qj609iCO7jnv64Ytbcp8AqFk0Rw8W/c
4vlJN4SdVdprgIUwEbIdHt128jFWuOgBONyhkn0/QB1C3mnzCtcvG2f8u7g5RoBq
ELxjaqKlAEhjBbbVTpeNA/92SOPZ64VMuqZZfhb2RW79oJ+Eg/Pvuf9aY53vCCtf
o1OvGqIKIYGZC/BDRhX37kTnOw8sI9vLrgFxk12movmLNLGWP1qmZjK1GLTVG8SU
qnIy5gDbnQWbBd7b/twI5CI4OUCpd+g5awMp/k8iqeWRwy81k5XBy9CIhqKa+bNe
lJmzOdv67+ASwoE3rC7/RJQYh/bMmLuB8toP7pbZtORsc3wOIGIIqUPQSkaTNWSk
/1AdlSKa/ugru18zHEFn5/ilMA2iwmmtR3WeVgQCeLFdMocl0hKwAoKiLkBDh+xQ
ginTHE/A93u8ilLcYLMQKjJT4Syr3WUkxOte6OL/K5Ohc3YrtKSskHxDB5i9Hu1X
ZCVqfV3YGznyPhNdG/Ctx9LapY1tvDs6TILb1Vr3MgeS9lY/7X0e1UgWSVgcPN2m
jEFqSDMLR83jkTks7l50UvN0PJMboXOz3WE/l0BiHnRk61S+AWzukq8VSu+NmQNu
2k64vTfuod5FLpL6D8XeaGm5XE/zInMJQ7IrprdAtGZ0CjMpSchM1r+hegAWNzkV
DQdxNoLNOVq/ykd/IIEf8s2+mIyNzfu+c7XM0dvL/hoyK7MexVIJ+FlfvgOqm1au
SwE+0efNPDWNLicjc+787phGKhaf9G2u0YQ3xk4xuGC05os907gwINPIJZvBUvef
6O8hVCyGzItkrIWg9MM25u6wiWcbg8ydkLMzBWK92VG53cOuAFD1qHO/mZN+73J0
0gsvcCovQdR2/AqbRT1OQXSHF02R/WDFtvOu5EpDjxXt4eQKz1169im08avkCxp9
gquc8TeV1mCv8+V/oxB4aaIZqEVs7v908ZVxfAEHMvuRv9EZL9RLIV+30la8F46c
28sFMfjfX4AUNEWMkUlrTYZ/KZwJy5aoTHplA3czpmW90OoG5mIGw0rXy5Xpsvby
9Vj5pMcDNjhXCvhK96+DOcDRgDEFQ2AKhtA+d7PyQgzG7k0LLvvEkPAfATWiPrNK
Rk3C/XM5poihFIwX1nVdYnYt/rv7PqR0IIjeCSjciHzdmwyuCZdo918/xpSaHs2T
dc261QIgb65ulV6DMTg+S6jV/FtLDTd4UpbdMk0KOnpRgng6Ro/StUA7hZTjBwZT
Pzq6nt1Qtv/ATy1oNR+JA6JgfsaRRY44OEXBaCW8jiwKIACFuZ8VDPhya+8JhssN
5xCxrdaF7n3MIHFDqo3VaxxVyf3cOcvHG2nlyqR4faGDUFzv6yB3QZzr+KVRXDas
v14Gd24sGGBfGAz4EMolNXQKZODYq9o3K+Nr8OeH5nyLzQvskCRGyPVvs02PkGAu
N2oZfsvQHCrEMCEKATeOSFTedCZQ6Ig97P7Jsoyu/C0hmVZTCBzHpwxpfTtyOZYd
lntWqODlRM57xb6WWdnpD0/mtRUVRpjbV0dZNBDMnPDJYVmB77Q1ava4kbz78kRH
OBEkPIKNbvvPLJF6UImpA5fi9brejDrxfFVLNjCS0Gacjbsp+d3m1IA3Jte2YTiq
9VTupsJl20N5q9glSaWLCja2b7ehiEIY6vTVu0c2nPGAX4lvq14T0xx3qJSMtHiB
pxDanzT8fptVUPkooFQ/OTq18SMuc327g01MubyyBTv2HaoWOBSO2OOkG3U0sjhL
7MgJih/6TjTeVYLAdpH4PfxKjGJg8LfXgcFS4sHkEl1GBwgMv6MavoKMpxogr1L/
5ErKQkuC9Hd1QaEUBbj+qpPVvd2t34KpISkQcYwbU9H5H/TetO4W7sbw/xw7FqXj
Ss7VsvKBPfniUrjDBGuERQwxFGBhfVI17RTHxthnsu8GhEOwIbNSJrec+6QHvHI6
LXxnwI2isGuAjIKnJh9qwdOsrsSsobMTFoFptlXg3CdizyaY+Du091bsufEeUgaK
D06YKbPdypQUhfM+a1tTydBHkyAgLg2B+Km7exKAYRJibUkyViJc0jS93/grKx/S
+ePyzdrq9Zx7zOLRIiSk0wLxvEV1dJdwxaRmLHX5yZtzoVkC2Bs4fDf8w7hqOBjn
t+GCAkhK5msNRyMTQD4lW6wEkL2GHcS0CDENQXtXVaCaFroixEewQ+IuvjH8j+g6
wH+qeX46YaX5MghiRsrl0hZqNsVcZsobcPygGQnzT9VlJyWYtdXQQOMEpwNAjHid
d4h/YSX+mXpuOPzmJJTKF8C6lyArKSSEbBnRvriGwuKM0oc940v7GrtctNBeBCaR
cvLEC+U7Er2f715Konah6buKghEyx5oX/wZuup0sIPr742rOqClVIvQssMVyjI2B
uMVfE6jprsgdh8UMR3J58ZtdFOmwK05ZdT4nRLlDAJg5DHZk73g4cqczA4f6OUP9
xV1twa6YBym4qmRIPs37e59fQ7zEJPf45JquTSk1q2dgJl31nJklP9Xzk1pkAkNR
iRu2m6nb82vInAq4z40Cm/DzQ9t8/vzn4Z68DtgIOcfTUBN1ewqYVhAYrqnsBb9a
bern9Xrw03AOZzVRZTcSlvvumVs/eRkzLlUE+3TYCsa6PgmOnvkAYFLPWuGraa82
+8swiY4M/I6sFGGcZz1BmZ58tLpudt91eDiozJGvX4ict93YnrxWQtc3g76J25IP
Xp2+kzBwM51f5XZl5oGvtD8ZC1QxWpukw5lra49uv8CJFHRj0fu2aTU2bELKdS/r
mFmPplPKB5oNf+sEkI5RmsLCtLpZ803RoYEoml9wkhXSKf2Lmqb3X02TGuO2kx0V
Uk4/4NftnDqAdaNJOXIzcM/pwKO/hA9PBShmGMJ+KLWN6nouTdGzTepWoarPulQ5
OMvD0r50LkYC4hUHd95+lNIjxnxcYH7zFzUGU96bgt1lnnnRDOdStTzJrX/1OzXY
JVIhHnclrSHapY142TpN1hKtfuRfTHa0w+WHDEK6HD3s6G8jAe1HheWns1k4acKV
Iwx7XXCyv4nj9PJ13zC2shDJLcJ6JioLEa4ULhl8F1xR9mkYKLq7jNV6bCFn81K3
VPVTmBWAqid3hYfjGTBEE46l6eJRaFipZK6oRxoQiFLxK8aSHJHEw5YO4pZ9XmAM
Un4A4UZs3y1iQtdWjaYmDkJ7ILOHvLlYFAGwyfdPZDooNGlZkXiI3JXMMzFlWWJ2
WlkW4ZPz9lthu1VZ7PUsRfwwsJL8sGex+0iYvqEYCbGDgGwOkvGU6KL2QM47M8Yy
+wERbdEptqCvWDsJ/xmWeUjnv77SE+PfsWhc81mWv+ZMGfFSeKpla2AJgb9OvFH6
rYN3Hh0xLgnsS7s4mSVxQA+3MZoLuVZ+5M7dR/2Bkntb+M2f0CCxttXiATsDB4Sj
UDHmw2sMk08iYWlyG5hB3Z3FEk66ji3PD6AMgr0o95Hd3w2THxUHOeYbilED+e9m
Uq8QWnDZHY/tn9wjbT6oX7O4H9fsOfVo8cRrLzSoBdGIyVR/Xjp7M7V0Qc9i5VcE
gIaZqn4aZgAENbRfkrZN23zaZRFQ+ER8KhEk12jtNRzxsv7Hymbieigh+f5PiIHJ
9H8/Nr4w4Fvb+wbvEtaLlVZBDqVkandh4hv/pjDllz55IXIXbGiTaIk58zvWk562
q9b5KJIQqRfvVNC6OUrOuQojl67wzPWiMkolr6lcLcP+MeeyddyQkxLPBlzOR0Ch
c2kCKjci/18K0Vf1oRH4cQi2XW73cnUIZi9pDuyJsJNY6g8O29FAtEUUoGMDzSKH
3++Aof518ZyCGww0afQOWBRM1hKPbyb2UHAUTY29pO1VhMvJseIt3rsLYoS/LTtj
9Gg1NvL2DEuH334idXkFj/S4finjN4zlLMIvsTjh546yo7s2mELKIU6ZkG93lYag
/CcnHXyFuxg2yitrr0p5AmicpdOITGjRX78FQ50V9Jb4S9ftOZQMYlBY4pIwWJj9
YoCsEKz/mzDZqkjckXn4fakcVEt6f2JqiKGhFBL7TTF3H5o1PFe2n28idHuMlzrQ
/ZCDzUoNzHK8vM9+MCRkK51CoQTMyiSdp6yvA+fcaQOnPy9QS84Risznm+UoiCwU
3FbhgRdO7V0XkPcSzu3wA4V4JHnjY5WzlQIz2lHQzrBQkyIXZISjxqufBzEyr2JP
abo40YXAiiVbAP9ytWNlqVVdoqhmqglFJQtAQTxet1j2Wfpeb4l7GC4q1gKdo7/C
GDUs5YcAzMEhdrkLVbtjH590mv5V3JcxhrXDEm3iICol+d8OT5z4dtOfJOnJhk1P
5YpiTrobNeRcsI/us7A9EMnXiQNhO9SHyG5zMrFTFH9Skp6TmlBh2s0Dh7SJW0KI
J+VcNnqvAhYy2mQE8lrNh/3GmvI1UES9qH6N0h5c4lJ2SeBjjZAUV8St22lk07a5
Dxy1n/BFH57FcyFEQeujKNOgWXrTtQrFPDvgmIsObIuWdw0KppiyNs0MB7qU2XaR
kqugp7Rk2WdwGV6EYoI5vaAr/WgFiaNgzTiUTb8M6feEoXLB3i/N4vunMtIQM3Ks
43doVYRf4HztPDsDEZ8GRymPqgWw+ZDATU2vZQP3q1Fo8etXy1Ay4FCcKkgi0KgV
XIsJiyUz1tE4IAumypG0Dtf9mbMSMv79DqipXSRfJWeEtzPMr0DRjotLLLj59MPH
GCKRkeYLaknMq6/dnhuEkGW+0v4ARx8UR7RqAdgWaCb7EDc/0HfhrVLzLYNnIO1z
6ET45TA8PQe6wIoeu9T34v0wPYqrjD3d5cDiTSZHaAyEf4CV0aD6gPgbjfS1PLGe
anlKsITPX28dVmUP2d5SurfPpgpQPOPDxOpAfZyOfC/2mIYtqL5+8bsZncdYJdoI
paC6ozD6304gvS+Nke9XrqQO2X4nz7GelVpIWOrxulV5qu1ZZ4kgURb4SWdnyYuF
S35MFORrJFnj/Jcd5lWaGVzvpfPemhKoy15Wv6Qc6KcbCbPSF/annigTwn07BhnH
0wKjXEbPybUX7YMRDn3EXztynDAvlEgTnu1P+3EACJsN4WbsJF1hp7IDoYuz9yL2
dRpwQO93QF8QO/OnS6ekMAAnhD3uA/aLTIj+AYIDt7iUIQqzlLMQG6PNtlL9QR7j
+FRRtOb4ejee3eFKjkzs684KX3zekB/BJGXHvXRKRg9UjYYO1RbYfoe5erP9Uue2
NbSDMV9w6eNAzWE4UwUXwoZTzydXTvXvHpLCO8CBA+QO9TQnphs0t6yMYNJ01oOm
C6qy8Xxp5sgQUDPfU9nirS+MkTOTC6vpiemaq+ThtWsUtWzGIdhF5NPFBpzsygpY
Wf4cQBKo0x3ZBagnv7WNmIoZ9GJJAIQUALXOFwU2752n35RB4BC0xB+OydFQaU/u
MJdSA83oa+MrD4wSGPwQ8z5I3RKb2VgfrjX14XQWmEsvmP4Uhotg479EZspozS12
1FWpXS/6p3EWPN1KNaLGr9YTl0MZ0NYUM9ym70T8iVEoj3XUIqY4XXMcqumzMr8a
5HIA4PIfOLhTl3ZlV/KRuajHelR24B1Ypf9BS36Gno4Ekq+Of2YS/q35et28rbIc
bIew35JQzbAhiG3W40BUjRasS1c4o20cjZgubKq79kZquZnd49ElCI3tRDpg1km8
FEgoV1xSxiu3XzV9Dq3pfLC3esLGWCN5ifDEjuaW6ESBpiUb6v4pHDbglxFu90eh
lTiwmIHd5CP0Oox/rD29NVKkoK2vv/8R5kVnOSA52oVjQmvDD74xd7qA8aNm1K4L
KWsR7CgFhTakfoddXZFpG6nXiR/6MTVUG88UTj+MnzlN50aa0zpL9BA1JRdiSg81
KicKTFYFsyKIpYy5HriYxD7J5ySEUZxD7u8Y/fxoRZ+EP57Kn382zxnJL88wPSXZ
COZ9HZVv4kqq1BB2hPxFg7sHJvy7kUssCF0m9gup19p5Ump6zFq8Q8aFNWo+U4EP
qg9JfSFPBfMGFqLYJsTJAwQCxuFan7lycZF4n/RlgwwQJpXyKXbMvc8U9lfg5pSF
Yd6+rt9idOwYhX75MpEDh2Dy4yeA81TyqCFk5ERezgYWgUrVaGTL0mdWkurDqAWQ
iGMC8GMSpm7sHNNQcH7uIhKOpnoT5y0ZNkkm6H0Ru8LgbAKA1YVTSDdISTcmcbnk
7B3UuBRTQS4MOwQqy4NfaKwTWkmbktLn+3XGU8BjyZlo/ynYUbM8NATfZp6Tc0IF
4Crfz2D5md2Xo2kZg/nYKK/htZY1al31h7PA8lnSCwr5nKXXMzHEH/yitvALlPlA
4yTYeZezshe+9GbBZkhX6umSqzMepIIr32RThVDOPD7SftEMoGjLRdD3g/OuGL+2
J2po3vGqxu5hzEXc+MN42EZLh+Selb/L6yAtq1sjviRknXQuTOe7GhFBh6EV8+x/
HUF4/0rurzMTKxktc7YRkcSS1v8mRDZvlzyp904+neuQ7m8U5QKNpo1DpKgjXzVY
Rlmm9gro0prltKxaf6U4yox3oH3tlI5swt7onJ1WzZJOJmlkBLleaCbNQXNvEXSd
tCQG+u++C3pBNKpMlUn/GRI4BnldpLJDLDM9YKHgC9a3rI/09NKVLRtsR46iSrAD
cMvprCfZR7kZ5p8b3OCbkP6N+3BvM/4qEFCLpGwZb7X74hNCL/3clyIgR3qKYk3t
r50IyfyhdhTVV99GT927LbKqQzqFWSjoFz6O7qm/O1g+no6jaRM++E6MlZfrpavv
4WWLkToYC1mJgFX9+4D7aj4kifujbhBTV9I/httFu/i+gk0TUUJCVsT8QCb3l8Yn
94j7BXXeNkb0zhObpYl7f6Vl9BhQfphXyyVCplqdLmKYBlIMRyLPxCMIWfUDf42R
jKj3CN12CoM6Mrg5FIwHBWbQb8o8LAsabZodkvJC6S+SlREyqUBp2WjLwH09qRBl
8qc2rNYy1xo4lrolnUDPDL+Ga4WujgJsvIF08/bVTwlFoik+BtSIotYsiDP3UlMS
w+4aTdTclT1egTZFn1H8MgXCGBNvFKfj+oGIfpa90tFreKDg2gsZ5EZnkPMumly4
BS+tnOKAd0Hf5u0mBkeL6lCOXC23FbExEaR/InJ03dYGNcOQ0P4jg+kRnEBd51DJ
T4sLOnWRtrj6DMa2bBpqR/JL+X5TddnULS2C5T3Aqu71DYRNM8Ut+/R3RxSCTf+i
xfkknbzMuXz64O+jWPemV9PYBRQiCPmPNu66gLcznb87GDIUrMsUGRj+btWJKc8H
UQBmAdlS15+zwVB1bgCgPPFDqVuZ3VEzZH9rlTXYAzxs6On7pf1hSbWQGAXrC6jv
HuQD5ma46ZXs9eHvP9MMNHSndqPQh9oSPgR0H67A24QCw6bCyrYfgwamCYYnnS8V
lsWqkJRjvfb71dBaWSIGDO8NOxUgU6apJZUKLeXJrri5wOJz3uxp0CDWuaJkNRVU
JMKejimQ+cP0w3ZZ6u2imyJCHar1QvPL+VpMB5me3SuqUNzLUhSj7yLOV5la/zbT
y3pSd8CN809QRRWklUA9P0KGTQiPZR0qfMe8XP4Y3q9HSrJtij66FY6fzcCZltdn
B5BMPnN+sXkHmFyodvl1CZMwbsM+Xv64elL9M8OpQsKhfMclGYuAyb+p7uQDCqIP
KvBO/KA+Ubc45iJjI66XL1WM7CF0RahSTpZt1+U6LHWUXTxuO6LgJxJWtVBFCx4A
AtiaGlRpw3izsM1x0rGPQI5OUa31feRcHK186/A/4V2DEI8Dkrfsm+CFebhzMIeC
clUXJSa+hBR1m3xyXYpicGZc1jOHbBDu2eGJZ/+14uf6yoNzGoCCBUL4rNwDfaKJ
S2Awrrc121JjaXLzKE4PTSLajcFsnUDtphvwoXl9yTR2g89G/0i+Av8mb93byaSF
zvXoCwn8mvOaRU55MOMscRnDULccZ28+nOROAbZ+Hp0Rals19dUicRSCT8nCnxdb
1opcGDN6VCiwnes4YDyM4vUWpLDLGMXaQjvFPB+0biFGxciHyEb2zXTwcM+gtp6f
ZbPVN5PjAKjx1uc4Ld0TSnicm137SYqHAH38R/VMTBDRRW8v+gg8n3aKW9n711co
Gl1l/u7dOzgL7NlP8Ip0aVhhyAQmxw6vCMcUWD3hw9WLUXkv2Ur7O3+OFDUSWHHP
CmKxXzhokTP1vTXhWK5/QqhwC5PM4UNGgw3qykxMrTEGmIZ0lQ69Wuc3Z5eH3P6R
iZD/PzCgjW4hs2LZvI8W/JmCdFVZp3TTHfD0ys+B4sq8vNko7fJRjn4pyBROEpiL
3wqvGfVYxWtB6VfYrdxjcdzzEn0NJFMbKX3h7FeqmrZFBAhwb46Riw++/OeN9GXL
/B3scUNV+FipKjf+KYALAdgvW2lkorOLQkPktnpV846IZ3sBPrZUrbJsgbW1K+3U
Ux83+Qf5IR4fDxFxtXcU/TsvLCgxH9+ewNIe8HT+ZPrgEsA1LIL9Qc3k9iSTralS
C2USKa65MAj/7VZA7vLD7U3FivLm995+L7XUz0QHrQiMCkdiBc/0KsOeBjaP1OfK
hxwNQJ2A35rugU7GvTDcd9N2HHcszU5T/k34t//DeeJly2IxKzFGbPT+FDEC+UaJ
71TN+VjlFv/VAwz0fDrzC8P9MuEuMAHiHXp25h/2me83bVyqHWsu54d0gaGrDVWA
6ys4CJHKrtrV3INDJjPxEUUB79Ql64cwKBr8g1fPh53cnjWIBMm0hlnoK+g+0X4X
i6qJ/twHQGZlgfCLRcGrJNTV/zY0wsne7qUEE6l9XH5P/7tPo6Os9xlaAeDNGTrh
5vx5SdPznLNn32xfzGrzrPUKiR331St+ssauZWHIxstCPtxUwv5r9x2Wdsz23/3B
W9nSdum6UjAYPk+pFbEoaVkudiyJZHsi8DB56ksQVjJzfvOMdeV8IvNiggVkgLZV
fH/3da4EGc84lBBp1sQC1Xn6Cn8MNsT3ucHd6JqJjGsIx3/yP7FMj6I/QyNvHHfM
FaMayZC/ljQNLgJ7fTeXJ3jAhXV1WhDrSLi3wHJrz2ugBcj1Z5/ytTSptzBiemQR
fBpO92JDa49xAE3MPaXQIDNssQysueKoryzDiSri0xAgabf3Bvq1G4JGfouZTWnh
qgpkkPIZJfhARp9n7kUhaqXZ28W70N5qpfyXNDPJPtrzUmKv+6zmnnyWVDDB05do
H3EY/8UuKOseqNXGXTX5f8Dv9102d9xVoMV2Mvbba2mNCrasvoSYzGDsE1gH+Txp
CP/pr2kzuFuZraQKI4fzY3rFiBsUAbVYFcb08htoZ6a6PnU/gNbIEZFoY/IQyfjJ
9oeyHcVHivseH8M/sRKFPR6RntoCk8gQJcpNbaSoirXtK5/gezoH2AIOJiN5MDbc
+22JwiN/pGoPQK02FtbV3fiHpOkPTL1qIKDxdgeH4pks1kY0cyA32qbCtrk/7uZM
aC5DRIFMXYE+lQH8DIaE7flYHavordhw8Tk1F8VVu3bIRopPK1MHQrjsRs5o/qJC
p5qrPpwksGX37WPbKSsbFGZl+mvwCV3ECUyG5LoQXSlI011FZzb6QqN9OzVEAEt3
/fc0GOHGSemzkTJxaiET+8OeaIPUNF8h8aV6BtUZzjHgDa25U9d62mwAsFliX4il
bNAlo38CQ/75SJH7xhDVVn8xc+HEY/gvFmExZbmmMNo6Jbmk07sUBjy8Vn8jKZbV
htKhw2sFbPWuKVy40SsDlLLlk8uGEX77dlKVy3WtS0s2JTew1F/FNYJ9wygs0sby
GT2HDcFX2Cl8ARkFDbjjdLLEy+yc7acyNzmgwvOTQj8dmrSTCeT9+9C/r1NG9cBT
eZ4gt0PP3u2zm3nma84yJiPoV+CmldvnIWtDHyqHX/OUlJkKyjBUjLKvuQJYqVH4
Pfeek57t/pzQeQHP5zWjzBC6X3Klxg65VZ4c33rz9zS5zABOuTcWjusZ4E+8entt
NoutxgqV7Zjqce9DBV+dB8PO7iYr4MZo0vmfsGBRUJ8EFXKEVKAIhnXiZ2e1TRP4
AKNxw91UnvD6JRt0eL/fcI57biqEjCzuN9TxglPNOtcIPvCsE/FXsk0dXnEkvjUR
gA95wUZHGsjdx/k+2IzWwWlafOAYBwIHguTob7QNGyYvSlL0nSMKlBWsCqXSnppE
aJ3p2saxQ0L2DApeE4MhmoLxMUGGj9wvz7AFGI2gcF1bFtn4mhBWsQuhtiN6SndT
+I604A+Syj6greaf28NWv35zqdl5bFAsWosQnD3SSKRBC/MKojkVlgln2FddE5Pb
LxzdSNk0HV3y3CjoRTZ2Bc9G9H5uq7gy/Z3xgXsp1TK6fX+JKBx6PmZS+w0N20We
LVDr2h4Lh+VC5xbU4B+o/OQr9MsOCNHlNMuxGnrR/kZBvLZGg+/cj8aOOs9SBk3q
TfgbOMVxQsKqAJiA1SiQbDU06hRlP4+mT/KxwkbBT7znnbE++BCmJtSSrNgI8scR
SMmMn0Nwu3MVEuScDZEwYElPc1klEWnjBaISJnFcWzEQ26pY0qKdYSLKNnDy5q1Y
/pw5LjTx0vkWmCDHS3j4Y/g86QWpz2btjZnLlwT1Rmwe+hGqKp1AwNkRlkqbZWyO
j5C0kqJzbsRtHQwmgO3kYJqovwUc+wR8RFG0F/S+/oCnjWIw8UX7z958Is82lFrI
+Ney9So2a3v2zpIBtOREGeG8VSWjf04rbo4KwpTxvz9EksCB07FezjPnOtFYsmq6
quHyAf8KQAMy4Xn8kuoitvH8jYANLm+RHshmqx6xzR4v4N4Q+hYTs8FL4u9HK1fS
xioiiTZEDTeL+fyst0bn9U3mKes+7tfN1jYPU+zi4yi8hLt/70CClbq+QofGa3HK
4nS8DxYPILX7j/QrpIhv7K1I1SI2Drwn6uw6F1lQMSAvQ9vea3sCXzTbts5phS//
UWJS/QQThlOWqweidac/upPR/2Otv9zHCT8Z4mX0/HuSTE+r5Iis6170ziSa1Dg6
pQS7ruHvQt9VI5E0JMmnPk9AAIAT3ksPD5Qp9KnkicI4nCuAw9NHDDpQuwCQ57Yu
GGPwdDoboayZ44UN9YY6oV/5DvXNIXVk/r6Y5ZQqfFiThUgdQuGSeF2rXxx3AvWn
o4jG4XYBXULQIWMf1N03HjOoqrPzMrTWnIVRzRPLcQzB0je5spFNj2SFntEtnM8Y
rzSQZFPrV9il1kfPhppxAiWpCR8P8+QV5K520kz64qiR5V6e4ZkL3SHx44HEB7HC
HW1MFb95sVniaPxiHXRaG5Ti/6KZ0zXK/yi3h9ES+80T0MJ8PE7d66BWSBH5LReh
hxYUd0AdWlDYz0RvN0LVSgwXOQ89JM6iS0rZfx/ZwQB8YR2HHr3kgNow39KetkN5
agdDQIO9dYc5tYxZB9bbZnFqeJ5griWLa1o6i8QSJMaMI5oY3Z1qo70Mw59NpSGU
heTlGySKJGlpr0mN5aZ9Mm7yPX6Ye1w9+1OkiSM6NBJDpuoZkhO9Fo1C3g0fBV+j
C2TOGbF9NgwD+5vgxygV6PWNMbGkJUI3Rs/cGOcPnmgJBJ/o3oCVRMGproeJHx7C
ROJ+FkWEQm5PG/P/OVoRgh/G8k59wwSwNHx8RRzhTdrKFkhuiJiCZvCYRXrj8UE6
FxKbsYRH8Qzc7KbniNlfEH4/37DMgHJjYxHufz9jkL6ElPRrqloJHzrhYMzk16Va
w8rJ/gl0qrz3wjF+u0Aqs6Cg3IyuQ/+99sY0fr0Fiq42w0wctpnUT+ZfnAG3lk64
OuS0IOqauEA2tFBY+u2asqnTcK3xVwrPzdWihHDU9whPrik5aaWmepk68kECfKWE
XDLjhDl5QlV4wlVvcBtgBYShbNTGqQDcuAu3agtkm2cP6VWs9GwsTL3XpzyMVpuU
TGsPgQHOCepVPaWo/Vz57A30IQErRnF+IrT2pFH7UxdcEGvn5WLSLqViBg1ypDE7
blZ7RDebvBVm9XHsRk2EPWGoB1ds9vCKoTLegCew5M+A7bgDee0OcIbM6SNv3644
1SeMx0njq68w4xU2TPQGPjdfxHbw++Ifq53nkLHlAA8nFtXYizwsUehJeBgKb3ZB
uk3KNfaUU9FfDU2pAQM1aypRXMAzKLyvbsubFgjYPACaZwD5RhzyYo8unrJxllDD
MkH0vikDJJRjJcNNFPYx54SdtUGbRbGildh9yy3h7CyGMmvqjxoXbAaffDh+J4Gq
N9Opj7Zk0fGWeJS3thFaN7rWr0L5Lu363yHfVId8aDTPQ35JLRA86exFE0wZi4wv
t8vS/p020lW0UIuz270WjXKlijNmI0u6ToMQS4s6v7oiAwO92BLKlJjo4HNqDeo4
mS6bwrM04L3iBU5KQ8qiICXF5YDtOPDaJbppI2OzZKEaVU72FI1DWdek7R1q5lG2
c18uyH6Nvhvcs0NzRklzCLi/vi9Sq6bEKB9TKp7awsqMTpWELqOURrz+02YhlR89
2RGoK2qrgD/rQaB7+gsXNVSmOiFZRb0RlS9nBSn15VPKDS5lEcGIDcgzSUy5G7kr
b2j7F/NhmSpcqpo2cuxL8GaUZxGQe2SQvd1z5SRxd2ezn+HKlpjw2kuEXz8tO3yz
mZUNXPEo45sYOwqm/H//+/JiBiqSwp3TsFiJqiYODf2dOLhbrgN7iOyEP0zUwKw3
g6IS5lKgHdE5q2CxINXlgrUTUxoIrheWGHz0r88pWBS3jeav4fqeYDeRvDv7YeNX
b/38G1V+5v3Uw1nhXDZUjMbntyDLZ3stKe9vMFBFsjhXIvev7G/1m9IOxk5CQ7Fx
kT3y/TLrTpfbiEKGk1mk2UXs2ThjKviJ+GugiyDodByIkmabXtan6+bjVmDzCRSt
rk7+iXnuUXIbF5vZ6rzbO/dR5Qlr4rRsoWFlyq6Aq+2qd95E95TJptFZRM1ZwxEj
LHOmH0ZjIPFHYtEgXXrciXz/EY/ABKcy91a41OXQGFfOkmrTu5Jfgxg+4I/ccvRO
BFy6N/4h1dYEpotyhlEf27Cr9RA0gz4PQfA/kWs0hsD0kc6KORDRmQ4w9v1OIsgl
RmlWRUVADVMv/Kkg3GvGzF31cmN3bncmblio5W7f25h9Mn5+zsqAG2XfynXOoPkd
YDQu2O0Jldmj/GlC86m3JID9/+F1Vzeuvf0MHCiQhUQxYh2Tq/Y7fK/6+IT+K6zh
3TTEIfUkKgu0B08BgU1gWASf9vktmphJlLFnaoeCSuH/g1VxBaBxBG/Sm/YouFms
D3gylsAfJqn4Rn60EqLuLListjL4SKe+/L5YW1Dvn4oMsVuiIKSnYvxxCX9HZU5k
Xz0mngnfMP7zQDmJf3nSKF3L1734Fu8kbsE+CtTOgs53fIdZ+APKRPkcMr0awvmU
IpBLfSRwh9YTpxDvf0H4VlqeDzcp1D/AzX4PqkVPXZtQ74jShRWRjT0nAcv3Tr1N
sebm1W76ocIIerJo2hLNiV4c7ksEksJW3BL0EhmEzMKYffSjoYkEW0vm8douTOJc
MCAyHRfOIJU0T3GLfsbAJouO+6njjUtMw3DNOdU+Ppw4cSs7tDLt+7HW+8kbUQx9
Q/MO+8KZA+ktKYUuCfU9QoG4mh/kVZNxMC1gh+hb7ru20cT8vXyYWJ53C1mNNPob
ypKWWPEgpvjfwocUdfz6HtLr4Wvetwgc3p0V/Tekqzq8rADXk2yLfGdNZF9LgK/C
3WlV4HZ0wMbbQ8ZJ3E1RVINWB+q3ViQ8NvNJlKEWSP94ZrrqLqPVsxOlChvcv5lt
PBu6sfafc4a7OFEpTxx43Pg5idQga2BtZ9N/Lw8Zso66wLMf4CX7CMxoqTmgWMt0
lB/vpx8pkvHArXbp4kZ5iD4Y1xqO1FmaEZuJaL1pC6Gjmldd/W2y1C/1I7hwtyG+
8oRPiDg2xWs1UkCVL56OShCi79I9X7KV4r9pzns9MWqwA1MNYIz06DtyR9Ebfhxu
AHJI71Bi5vW/m0FYVoV+53lwqG5VQzx1W6sdkuw6GnxWgRBiSIos9kgsEjEyj/+b
blS+/jjqqQw3NiHy08IqG3hTfymak9+pCobMkXHq0ul2qZ+jEcitqYYSfwkkiWx2
LDiRk3ftSUDlKSQYm3LElNO1+fwlZMQZxWMjqtz5Qwdw03GNkQElPVyo0p+PX/he
PUsQ5aYKTZPR4YI9aW9jF6JQCMAPUuL9TbuQusqqMssU9b1+Otq8xNIDItA7Z3GJ
btLyw+Mzmy8RuwIB7mY2EQyrV4bkYKyCPPHD7GbZOtj966Yv2xKM+lS/LqJWSYfv
dC0iRMLw8/FfL+l9Boo+WoxBspJQTJqZnvm1qecWcs8vlk0dR6yWxbk+bS3cDQJj
fp2WhtL8GOsLrGGWXOTjVkkTw1SrdVzU4DEvwJBz1KimJfm54pvMy860+1ibzpRM
di9lvz+tzoJxd4wHtZu/yXl+Dvlow/AJT6+1aBWBXU08pWcz/+b4yFadfhgOD2d4
j8zC/gI37gwsDmFBsM0U3ggbo6cap6nILmujcYgOc20jB+RC1Yk3/wuLGEhZir+B
OxQIoCBDLLBfEeQiPQKOxxoyPUXCplzeoS6LhR3TDnbZNzDNo7toFO7mnCOEkzXZ
6BZj+/RGBVeHewmGkU4Ra/8UGYBkbDpCuYA5zmzNcGSX3klD8UCSg8M5i1+JSCt5
29eVlMauA1GHwfEz806b4N6uvdus0nXyR2UKYjzQ2KgbQjmYQ8UKJ9XDdBBDLwzv
88mCatX5iFYG5ouhioWGoTN2Vtx9Fzx13d8vN7M8RmQ1BsV00OlGsVj1TGAGbqSc
UbltTw88xz6Z1hqAUOcUOgJGmUCzPR407wtfhGiHJtBZrzWbE7a3t8/dK4nv4Y6q
sKjuFGdabQGNdL8BM4d4lQxYpuxT6ZKS/oaDMvXMLHlfTAVVMr/JH5ANF3oM8FiD
Tfqe2LzK6dLsdbrRojxkLLc/0cTMemPeQzst9RuP1LDqPjIa1x/ebGf+/pSR9dWX
hh1zk+Ligq36aYvhwa+KzbZucCZIswIbvqtrnwKg90sK8Kaue8OwzNLygVQNU5Yg
oSEOMBOc1mbBUIuCdT1aBI4G4FNgxp7FucQEckOQ6Em42ZGp+anAGftCjXlwrDSl
DWxI9sVZXErtJal/X6LfYxq2l7KjfjrC7SFCJlNrpLxRSxXgrRdRR7jQW/wwFaDn
B2zjEYrch1Ak6ePr0Nos+k6EZC9k4vqGPbM/cfETmaXbzzIDeHvQCWM7xk2QjmAv
/5mY83enm+mofweovRzzMUiGTxkhRYUfm5aCNGjiMTNvX6LHIkHR57hEzb6WUmKT
t/PY+qQFLKN7UYGxlITOmG5l0TUNmTstguj7wdcmcvqVKtnvYIvs958l7f8+8Elo
jQgmtEpFq7fWfLaMGC0Ogfvsq6n4uFN3qy0vi7Frqw/w67XyRHJ8Y9fCI8xvMwTr
23dHacZo3GINwAcfvwIDUKJZCpxU1MkbX1t9z3cZCKlvCuYq5PiXBkJ3U/teBPEC
bn8EdD40aeS1lUbuEFJrA9lrq6hobCFhm6nkCz6eB/zP6R3WM3LsNq7KoxMZUekp
hv/Uw/fYICPAnygORoqp3IOj9mO5WJgI+OaEj11GsfKRhuBpqsYHxVo3RtVzdi1b
TWJJiZ1XwOxWpBxjVwU37PLYeEXg9fBIX983yhoHvNhLDr0sKpHo12eo9KvclveN
d81nQqJLZ12uGwdTl4KauT8P2n6W8vhwJXJjE9pePOeJ1Z0Y9SIozs7wn76xdhwC
ognleUvIG3QVUCLEghFlDfDNazH40oPesAN72IhPkvKDPQ91kajRznM4G/gO8FE+
usPESkUltMOVnryY+1Yjlzr+NfzrfoL4LnXsTYYVNCSDVHFAl30lNKXa4QMYb3du
7Qxpe4qszIYUAcM5W1GXCyhaKcMDvYMHp2DfZWCYkgml3+wXr1EfpydbEooyydJd
J1p9OBI6GOkxqsZu0abvIwA9gahxr+1lVikd4cVcm1IUZpTmIhEtAPIH2Hv4TQf7
tftzV/B7xwm2t5BA91m62Lg1Xuxu8jAf1zVVijIWXtat+qNlzwqRSH/eYY+5QJ+h
myCQUlljI4NP8/j4+ffLrPb6AppeGnLQZt4I8QvlFw3d14EyvS/Tjzv4UZuegC2w
WW28At0oxCohiBYRM91TrDeABihJII2VkQUhHvQ9oUT2TbG6Kt30Wse9wSlzSuf/
QhhQsL5S8uZC7x2ETdVxHBzA6MfuOaswS7AQ7+ktbtSCkG4Nvp+oMvCsATZzPY48
sFXFZA3z+coPumadEEnXs60h87EyEIcy0U2zWhw0wpOHAexthZidqAbyAW9XRFk6
+3usvFY11sxzu/Om2pZiE7R2z1zoGsjllTgSwJ9F6Z0AFichGR5JZ2/YtQfe5KY0
JR+7zMxFFDsvooG5kEmBAka0l/H8dvyRUn0gABAMfkROKoCbDkEmMd+LPbwoHPNg
0WY6frkHU/10uv+nmfDEJJYAY4ByF8/jOsjAUStnsRZRuUTazTxpAJPcatryVhQ2
UFnMXbLoos13puSxelA5V/cQ8CgdBhjBdK0XJ+n/+Ys/kdCgjHa5CqwMmsqaDvV2
yOtghMNHjZFEC/G1RXPRWqSymGlqDFask3OEiTV2mSejZ/xbGOKH0dLBRvhsMthj
iUxUrl/PF2xRK3nwc3NK8Qp3Xzz6Tfy3Imsnzc8ESan0elOO4Y64PEHk8Abkjgy6
1NKKCfVQ2Bi55WS57N05DkKB8ywF0MQt9afkj64gCaF+pzKrFeCYBqDeDBnIrxL6
CFJTxSOGDyfs+dv9ScGciBnzDXdfAWNrNKf0bxE12rO7hhGaulArkUWb+CqVBnmi
qYla6JKGM0sOnfzj9PULm/0zThNO0Bf0jOXTThMTgKq9U7H2L12kSYjMli4cvgJy
2jG/EdK5oMIYAkzRypyr0GETt4W6h9J6xiiXGHhC7nfZycziqffNWuxoffs/eu/O
Zb1ouqZoa6P3t3guxawh9llx/z9AERcVoklMtyL0w9+JlFLNQgKZqRumbFV++M3x
maVFyGVs1yDrHbfOjNjEVtwrYIer4YAt4OkbIfj4mGlMTEGQMi6yfyMtcojeMq89
NgHn2Cy2yI96w77/iu0KJBxYSylFkloI3y8QAHqy52WT2kS8lbjA9S7g4nneCUVC
bv7QXLFyPlLjTh7v/ZrD7MNLrCRyz6DCSIQySQLnBtkr71o+/7FitN5i08uVyJnA
jCxEMAPKTRTm61FLahl1eSJfJLsNQ//g9OFxtt4ZC8nrNzgzpu7/fgadslzyoVIl
9uVZ0ZPdCUKL2EOqPuOaOS6QNKx4WJp7tf6bQ+w8QGeYIfgjOMKywLeGrdor/0Rb
UzcUd1Nr1a9uxv3ku5PEFKz109EuND9sEoT/HDFBobaAYq8F2TDrDr5eMZ9988zu
bTLoM/FL0IAfAvcXMHaRHy1wTRC2CkPjPbUa58hiTFkYwJhNB9pIDTahP/TxzDw3
9/Ew0ipVeMM6eGYMjvHhMncec6dWotBnmQ/u6RkO62LKD9uo3yIkLg8TPPY7Ge/z
d1Gtkf137G4I25sLltkM7F1JPAHZbDr7yPhD77BKxdk0JyuWX2ya74MM/Xy+9bZ/
zmVQC5bnEDjsppPU+6LLME3/3plwThAbTkrzvaSuPX0Bk3/R/Mhm1IDsopSpRZL2
jbJPdDIfh2vFOR7gisI5aZeK3v5zW/FrGOo/I+NgKNZI9rfA/qadj1fmhC+JWi2t
uQdMccNNSWB2JwwpbZvvVdrEZ05UJqep0ifdT6585ftkBw5Z50TUGmp7tD+7zds+
4Yi4qaMuL63wOHuz3gMTnPlwUl9C4hAg/2PH6uD5mtz23nBEPxlQvMhAQ9YWVlEq
/21QVpvbNzF5qgqxFV3nmyO0fGcGUKTSmuSGWJH59cshLX43Tw3f/HtP3Hoc8mdv
J3vPGgq1Nl6r8OH9IVtSkXHKdKSnxfxxDIV7PiNsQv93GpiFaGol+A8NDrhXBgG9
QHrvdmn5a+zXI3fXv4KBDRE5riOpwjmB6/GwQrtiPWLd3OBtcwM2s17+Py9FyGvB
gQ8P/o+oifQaI2VVwHgaBH43RtYG5GAT+aRAtU5rA3S4tuJqHnnE4oqbYO3+eG9W
N46vO3xK4bnu114Za0T4Kdg/upkYH4U5IkAM3oh6o7xCrEaRAbSelIiGe1yBxVWu
DANCAaNj4Sk2xRds2cV3Lov8U22YFlaybAXkEbSJd1vKmnJR2KTZU8Hg0CYxKUW8
GAFnohfyyYIJakzBmz0yEKpLXQyHljv91Z5CopUNSe/pdcd9fw3Ko+ofDz1pRpl5
yWyWbb6KV2xiKRbpq67K9cZaxsCBncJyQpt3f2SSVaZ+FH023Ge8hnejMGHxsOFX
zGm/YMGFf9zNS5steTJemdvQaveSvVRwXTSSg24Iau0pX7CGRbbIiJD7pfbvCzlN
xRFAtJimz5m/E0bwQq/cZRBz02C48RQ4VJQA5CmVk/B2a02WLi4YLUGm+XS+QMnt
4YTwX/1IPKbWbswc8k7tvaz4KKfqj77Yq203sX/RISvvpHhkSlwru4pGi4kxLvL4
/kqKUjvnu+/f1lnhc1+7OkOaQt5stnfmIufmkyDVCDVBIze/9GZAxYSYoSvft28j
kPFUmjdizUym7FJ7zZ9MrOXspvKfonMLPW+b9EuqrQ0MHaFLtHlLH0m0V1oAsd5D
+oj+vaQcHhmtuw5mbAljoPEvODHSfEmzrvI02VCbpDa0FFCYxAhw6x3LwhK34YSb
/cOidGql53qRgml9j05yo4Ij2ThE3pAOMqcxtJbceVNsb342Nbdw0OUOYXnllzaH
CihE0MuUiUcaxj3RvgGN8J1l1u6rVC6ZZL5O7KPOvzfoTFO/kdvUB7hMJzbQajJ8
MMpUN0SSeqhNSzjKe5iS3OAWS1zZ+wdo1y2pgbGY2ZtkLMEX85QDzBlWJ1P1hZiC
67akTURnhfdT6ZmRt6sHI6oONSfR1fwmwzc5uXkrf+K0aRULa4SdSem9Z+awSmRM
65IWid97+S2FVALWZ/k9EHTJT18o0gMoMdIHM0OIfeGZ22q0wV3RkD4gzpPQIAmI
kFgwdYt16BtjHd0Fw4C7EOGFs/zbYnv9rvHVH8pHSgLD1aAYPUtHf3DlJtVAgBrX
ALvREAstacyoWX88IYyK5Kakc19hz7tHmpJj3RH8MwRYb9X+CVzzIQMa7vC4pBxK
qp8LyZ8UX/s6ILvEs/UjzbOpeRp1aNHLFMhyiIaLJm5QinCOFtvgOkNosaXOXOnD
bl0245G5YEgLbNh5jOZzb6ej5CGnMTUZRtgJZ2nLh2ySpoLnghhXYT5fT/e7vL/u
uf/9BfQVNXhE8NP6862S2OPM2kr4H9VJm3scDwli07khS5L/D4Gl7G81aDHZsAQF
t3t5Anfa/Zc7bcxQNNPb0LYGnymuMFfs3pRXIiMFTEAUsZ3M1FTtzLyZmuS57biB
kfYfPju0QVlo/08rBEobdRqTH1ShT+tZteoqSObg6dttRdJX9mLcqMF0rgx+zYn+
ycxP8pdlHr/P9C2ZLd5k2/zvH0E0QYllZkPogKUYuKDqDuCQ+D/y1iB8KnfxKCBz
RLxXJbNJ2MhBCuN/wVrE3RzD7tCHrg96b9VnYHjzU4VhJQEmI3Z1Bip/q8aI7Uxr
4t0BnhOSzoHXt9DgAHpkk7Bq9+VguEIbySHewjc+kzmBG2mXaqu+bR77EjjX5Nk/
WTsDBWNOBWMzJf8GloCWFNblXzzWOhjOZwOraESMW8BGbL0dFVuJN2hjgLE4PlGo
qgsiHKmBBleXl+Worrc8RmlaEgXiS0WvduIg4eX86A5LIlRwLA56Io2vL4ax7AK3
6AwTyNfBKn+SAitO8YvBDXJwpepuXhmHmDB8PViHHk6Y90OUqVvC0B3KM6JzRmgs
jHHG93qL0nSGm1JNHsXW7UIi9QGFx8z1AUEUHKHB2hxS8WQnTbamAj+7BwWhh1X9
WFbX49ArxF/SN/5iTYsXJRd30QSbzPpflmwMbizP/u6GF9oXqzX/nBCivvKPrD3o
n/Fw/2Z9m8rTyc+WroBPUd85ADrU+AE7vDmP0Pl1Ij+1B9guJ2ccVXzLLTJaQdkC
DEJZn95dgZBhx1laAETda4pHGuLgysJuB3nrjZlrkDs8EKP0za7gv25DdryNh8wu
GhPmMGdQh6U3Ui82qCNKBjbCxJLCKh8i0HQvPEYbvXYVhuJpPmvoUPBE/WLnt1vf
OH6U7RZxWPcdUboKeKuZrvu6iE5S1J/zGQHEEWgwAPfgfnUCodFboQoAE1Brlg+x
Da36edDnzFWWrKB37YoRM7xLWABvKbR5GLffxsRpYGDMAe6nTzzLgPI/cLFVjYVq
UltN1sOCEOiW0ziZmOxSywO7hknoOopNg9voPAvBuHQLBSSao70DjggLphEVB4nH
aNdQ/c+yRpsPpbHAuU6vPiYuL3vRH0Rt+joKsstIk3xy/UDTUo4QJce+/SCSfYxS
KUOvQ+kEbg8KOo0YB3jP8YeuQrURtvDCyOPwVqZUTjAbzXCalO6JehMeoSOrCr0r
+1A4laT7sSDxcw4yxAI6S6VVD+2rHTZ/CjQ1nBOl8sbsofaA+wdSUAdNrwu8BOo1
+l0lPRBUS0AsVkdCJHdefrfVvvZySUzslUxRuMD67Ue4bYYwvVkM1ELYVQ8xk11e
scUwe7E2ogEJ7jGyw0aqONLCH1issrKhCy6/o5gb6OMZkJGwrC7Du6bw/X/ih5N2
+ZC4uplOI9c7hapWNDH3JnMhs+v9v2s3wxLum8zHo9dQKw1hXwSWV7PMhvQbHwNK
mN2tB0Nqjc0CbAUEsfU/j+Fj2XMRevZIG7JbJNRHwJJrXZtneTfnifKrConeZczO
N17RpcwGid1xDcBRiFdjKQU42hcjMZJwVNiER3ghk5rGRL6C9PnWz+cBy5wRQtLo
Lfx5b1GFDTIQ4qTagVL8qcCxOXjhDhgsL8k37NLaS6YJuKVfljc39iUplTwn/p9H
Vd7x2DB5yE9PtEwhBiZjZTWKWdK/tQzlpmqgBrKJVhM7dq2b/0hcKwy2q6/VzMpU
Q9J2l7DR2pbs08/JhN7DYeSaFaqrvPesh+H0wgzUHpXNtvQ5q2Pcpv1ciXKziSRd
v9f2oHOfCxz+7e0KKX1pYCjsgD3wJQ4HnOFaT8p65z4Rw/yuBEMmDa9Os0uGz2or
/ipFUXEhZYwj2ascdYqnv4E0IoXibkND1puIcIoriVc3Ikm10d30U8GbGMDHRuW9
3tyGHTixGlZdX/YQyPTzOYLl+xWiAD/Noqa7B+40OVjeYpMSypg4XC2MJCSV/kB3
oSMMNY9YR9jjq11cfTzrhacyNvm28qV0t767AZiAKUWQRQu3KTSjkLN8SWAJVpWf
xlJ6hwKYDaU8EBDI50VQO0Z5elsT1hh+k4I5fkolaLBWZv02ejsnwfFEiYdB3AWB
SF30dW/bIYEHjtstmS3FEbP68qQWNAEqHl1+/7eWIlRJcxaGnbJzUpfINdi5Od80
uX3QfUWkI0acCxXsx+L2UDnTTziAjYVqA0Ai5PZ62lZDLupTGbQ+c50ZYkXbK8xp
9cGmUaaM2ZcCxQGH40W8QgTGQxnEIClpl9/NpESSCkRnzMjaf60leFTis82Y2Awm
qZAgnt+uYCYI73WrIYtUAm4pcsIPr84aJt6JT1l1cWkiWjmXgsg2kqVWjx32214L
59B9NI9vU1bDH6vSgtC0sll/tj6N6AsWWNqjy5W48epJRjhIERIljCiu7eZuGqIQ
oPc++Ax0iljr/XvjJDNItji2AoZY/VHLmyMbAndwJEH+Ltu9gYk/K5jGEdZAtLQ8
V93B7XhGg3IMWgK3YFMvmL0w5UHePa0EmeSXwAKzx3Jp/azzwwynmQIv/hmPWiK/
p3nJxkN88qU60wVsd5t1vi+RDyeWHaG4mffU3qy5Hct+Y1N50HI2aq3eLQe6uCtG
MC0HfgqS+hiGsj3wbbUPGYhxiffdww6oOgdHr5pKnXGtWSO9Dvw5WPrDc6ZTWqvH
vI9mqsvQs8rpOD2Kg3sJRFzvimBq4NupEiq9iHKyddLAuxCHyBudoJBieDenckS7
E/NwttuAlJk/VLMGYovR8nsImKtzQCxKNfyZpHYFPBz0cxkA+UvTzrCMjkthlPEJ
f4nqRn68Ra3dgx5+OvwUNgl0Wx5gMk5nddRNa9I+eb9BeznZ2RfIHIFZGbqxzWR4
yY6fFKpgR2uM5jyxi6topmwSU0+y/ViUBx59qZp8c0n2+Bghwy4uKQyJLZbtUleK
QfHfgezmTlhdEEaof+SQy6mkkpj0IwR6RGxvIWtRQGE2PlffRW+ulPhzHTzeVIWS
jBjmTkVp5h1K6SfEmwyq8iiiRVdpqzE0ebsrJxABiVhBxB9PXeIdTxPmZk3h6KGc
gHq14tL5EUpWMYeY0fE41SHL40Sj+PmNWQPVbKjf1nDv8GsjTmhiFnmmJnnhW46Q
wtTfKzph6tWxMhafH2jN1FqwqHUvQ+ATjFwHctuQq7p0eO2U0+Aa2/3PL6ufvlPb
HCrMozfcKP6Y5CuEwY83eD+1f/2j6JPRHtJpuPuk0laWwJASEh2KuOktRejsnHdZ
bwFfAXPuhvtJ582i1GlgcqWs5J8MQrkoVBtuZ0xG70VfttfIMOe/iRzNwPMwZ8Mg
8lShsu6+4a2gmYUDNYX1WDteDrzwPSZ974kSf5Hlb115lMCvvpbAdi2iIoW/l7lk
myobt+0ONzLTkqLrZMVbdRlwJLmm/FFBZSG2RDeFvGGVjmFr5LZHzVjAhXTx2UQi
hEhBrGlKTTwYwqAZoOR4zFUZRtMcwjE6B/PoyB2Gs1jPsPkabgULA7T5DlHtLdDj
oh7p08Yw2jl3jYYiiYv29e+IYzldipEogH6/mFkphqEgY/bc8LzaTgi0RRDDoxIE
DNH3pVzlk9JUC2OLaG36qjpzNgMT6cJqW6y+JqpI6hQOjI1/ZtwOqGg+rkET4luf
dbf+nS0IJ6ADE1kmBEluULOg0jhz2In4GqI02+3qR0aVSFfCjPRjxM9Gk5bEXrHV
+y9bV/ZKDlkCERpX0pU3oPWKuOE2zXEPrUg2p2sSJJaQo0nYO96hAvrp1H3umAFH
LGfZpa4RjdnxuhZTxlK801I+B+uabvul3SZ+G5DmOnmdgjye1TJiDVlAV0P1WA0U
fN/TPLzvfeomZcmP2IJLZmlkl2HY5dZXynoFPYHJyrOFnx7H6iSMXJ748d+Bg1UH
U75rDWaqqrgq2bRkCf5G6HDXykXG9Eti4j3FpIco3/boO3FuUv2nCaZvBdKfrvkt
BUJA3M+Mj8TbBQZj2bfwaowgcMx0dA/lxL02c6zmhSYKxLfs4FOaEIPlWfpF/r5b
MIkxaNQ6uqD96Bqfyj2J/PrtyXS74cXOHsrU8bXonNbfBPV+bEMW/JebcxGTucsS
ruVufccoIql2OB+C0eU04D8tI03bcXkPRQsN8DRl5754DPNWYvyE2/6mEwqrjirP
gPEQWEcGYGk+YZCzBHU/HaaJxbEyItArPLKef8xhC0XkgoNiqVFTCd4GbqtsyUHD
gCuDwxvEefOVbLTs6onPCMZJhVVhvtt8uVV+3tgKxaSdWTlQn45YfqZTOyOgWpEu
f2NRqMJH+TgTNU5KI6QG2UFT9WbmFa8EQlwZ6/BWs30FfxhKStp0er1zH8lo7k+X
GncSVPUIUhCYgIT0IrcLpiD3fjm5htGjm5qcb9S+jDn7TPZZ5clSl396y0Q91bAl
PeS6n1qXI5nzJh8br42McCt0XKUZ8uwHEx2azpnnOsY4QOdTsTrAte69KV2tkKRn
B5JHnNPtFtQGGJqsCvTQrgUZoZUZ1ClaFShUp/TdRtDkAJqWGVIt2DQBsIe4jl/I
po7lCJ2HdbLCX6W91P67qS2aE6CLFjZ8gtzxjFf6N1ESsinG0bydQpBHDg/fuVgn
Ffyx6vKYjrzBxQP8gyW4nESWc+/fMW6FME9QnffIErqTuR1IkNKAo56ga2KNC9Fw
Uuh+aoEtXhGgZJvbY/BVo1J8x0IbUviyjKYg93P2XCqIbDPAlQurrTVdBgaa3kSh
fQjcujFNOKpbvzENboQgdtZIqcHJRsEjGDdrXw8IqUFApip6Feu86w5bsU8gIM58
YWmh7yBgNKGpS4XBiMtv4HNKyImvEK8srTS6/mPFT7fDDQC4cfkWu3fw0a5mxXKi
nmNFoDCmO1j7F2wisHCxtW/xsb1LnlzkuNLnX/vwB+zytKWqlfNXXZF2QInB8A9z
E0aa2gAakW3t1YuPEEGibslT2nxJX4RKUGUKQtFdIHoim/r2Zx+fVTxp4JEP4dor
5nqL+nuXd19POTm2FSCTKZq0I8aIgz+MbU2M9W7vdpfm0K6omLBk434FLhwZxQV3
7DEoDyBG069LwlYeMk9AEL/wxzm7p9nPVvcHVOZQPyzXp49OVO48at5y2260W20S
PedRGWXLbq7cXJ1EF9CwyIl7x+OtAlyB1vYTGBNfUY88A+vuLSwG4uoW3qWkALCM
TTd6Yv9vZP6s7tGEc5+VCK/Eo7Cz/OA8fXV1crzsAoeJIN+LhSU0/Kv8nFiI1DW4
SG2zdkHccAfQIxIg5ED8cIjmrVm9Js/FfcIfuLtsUSoB4HR9dJZFxXxoxZwvijfk
TvUkkoA2EgBmqyJgK2B5OfdLGpiF2V1j5VkrN9RBLKmQCwYCDtPSORz4wx82N2C8
dAmsWoVGGCsZrRIa2mI3vswgy7F12UgaeBXDrrMlI14p0ZsUS6XU1v5HPs/4gc0z
NYtHXTqfGrh58u/hWcWRH2ON3uptgwz135xfDOakDB8gDjeCddz3gFsrrggzoKhd
XE7aaIv92vj5BzL42l9tTYlG5KapKqNAHmMBr1BQ28kgSIq3vKd7VPCWub0+VZGN
AqXpqnOwHN2ZqNbljUGQWu+P7M+acbvWTWrkaBh27g5QGK+tN1QMjLduR71HFIAU
+8z7UEPjfHLOTUyJ216pT9Vj/bJiQFed/lLlxFaeFCx25s411tFdtNajDuZaTPEg
RkxgkOyU51dH5ISGF1K2vjFOUb/Qv6WpUaNJjynRhVq+mlTSmwetsl4klSr+8TwW
Y3zY3c/cySG6AIyLub4yN9/Jg/Cc8Gkt7Izr8Se8IJrdqIOw9YLBR989EURb0Bja
Sn4ROh7r7omT4+Yio3oxcw6eLoGBTBum0SF0r0JKGX+TJLIDG/MTCZgaL3c4L/0+
0GZXUHU1A4YQVBtN/lTyYrpiOManb4TE0cZzxsj4rr6pWZBkWqUiDdHGid01L+wb
DOFNeKQtUBYFPuxk3tdsL9HBTGnae/MXlgyQKDzLbNLpF16xvOyyFZnVHQCfQ3ff
3PjDt2E6QKyW0VqmTqr/vcxzA11QMttCzw7nj2qCsyE6eAFtkgNqsXTVgmYN3J8j
PHl/C5IURY4WouTVfTekQrGMC5OQNr0u2sBCdTKhhlrJADaNyJyQa9prGJ+nAZCB
ZNiacs7/mvX7/dE2En+pZDYkXipKPut1FQI3f/QiUJzRkNhVNJTDq6IckBmyINo0
3TIyZc1k+4PVrGuoz1/QH9mEEqL5ssplsS0sR85iOH5OFYrIzWlU5hbpOlI+nKwx
xmrXcBapgEfgUvBCeF6/uvE2+JnzyscgEmKJzFRn3/Mi6oGX66u8nWdnuhi1qnfO
RMd4hyPm6RCvK3Dquax5XF1dm5rH9cROTmMUARtq6eBXNHzHNza1QZIlxktM8xrH
WtsEwutF5ZPzAmadl0IMVw2snB47Nz0ObsIw8l1TZAeZ/letDYlrvUxsAhB+II9L
L9+eD05dkpK9HjVNV39pdkBI/NCWuGejuwgorF+vpw8c4dS3qMsXbbLa08ltcPmR
g9LAZFYqrsfsbKSaZGQlejMw0xCodBUf+QQSDE3vnCUqoK+w5oecERXgx0fe2bGn
QscVF07svBwjYbgExY3PX8+pGjaBz7NqBKYNc2KQZIGA/6WFJJPAlfHhvTBBK5BB
+x8bZigc7kr3wTc9yv2nfXaa36dUSk3IcUbypreCTwDow0XxoMVbAqlJPRIdKhcQ
Ls9dV53UhW5tePzDRE+Y7v19TT/8kuhdEN1SUEPKtPmiORmNzNns50BwVtWWiUOi
INta/yodfCIetyehcWJx7UKW2X23PVEmqFxS5JUsbJsfuyBL6Cdt0i1Faqc2+0Eo
5TzINqmsgrIKqgYuNTNn0rhL8+c04yHqCaArA5QWO9gfXncSemxUgv21pFnykdQY
3m93hgr3bgqvsF5XtIr1hvd6nTpHQ1n0/JMj698QwsWKY4aco5wLBmQ2XKRMv6Ds
fFzN6LV450GnSLDNosoBj6h9IrwSztO1UfrQ35dQgKYbfK/kF3tbjIcOoSyXb408
eUIjlcq9Eot0WcmD38BWDrtMEMd1lN8MOA1Ly5McpMe0IlItpKld5pZm9KBSxEyy
mVfhfKncoSHAJJfPH6kEIlY22rBVtBCbP/LQEDA+1I99YuLC77z5o9HUDJGsfqvT
m4Qa7zl2g1UdhD3w+13OfVJung27dBagyI+/Tx51gP43DCXQ2Dr8/p9EdXAjPRxj
pjteujwzfGzkAtuzaA2TAmaBvz+CSA4tMzO5kpvlEUhc2Kqs/iytv1sHpX+3dkRg
TniwwaVutgiT4l8u/w6W6oODS/ebdVhyUovtQGJSRpaaqQ9cOzwPAHqvoPoivnjJ
CnFxAaGpVVVMAx9hcT2RuGtiiwOMFl19VInUSB/llHKt0aC6kIKCp8yOIeu5SCOq
rFKzs36zZCyqXJCcTEewNpDttHIgwmqi3szvVRC8sol7oHrchzeGLjuruirOEBxS
h2iUDW/OG6wKxBZL72Q+2UQ1LUURehhWh+s4PrtLPJET1ie04IFOj8qomE2X2j/T
fz//WgOTkAr5pnasHk7PnIvX083/8WUCBnjDeTE83b55dt0wiDB5yug/qmBPc40L
ha6nzEo2tnrMa5PDroprulSvJWEFvSsAOQT46wCiNbu7byvNR5XSyJ5oF4J2YTDc
fEHy5rq4SCsYFnzezUPgzuy0Yv9jw2O+fClFd1Ble2KGaTFghPQ/8zws+lt+e/qh
fOX/Vx9X1K/96in23GzplN+l5LIvjsog5CK4eWCnwj3AkvCvhQYCrL9L0BEQcXTK
eTh+XPs5KSV4QXfmBW5rVUWLDkPaGMFcwgnSfx8dUwyAzW7It3FDrD7Mygkhugzf
phm69rgspKOciAXYpyyx73LbaVCfikDUg5reuAgqm5BcyHk48BXxQa/1++ROZSe8
9NiOqLOiihNz2MDK1dnb7oZ9zCTgyqZKaSfjKL4KsMWONKv0m1OELY36DUUutZdA
RJxYn1OsDgwI83axg8yv9EN8SmkUM94Zhdnf+WtCJHpHMXXmdm3NOR5gSr24eXEs
5vKQSOzxHP3OkaXOxzfRYQu/XCaYHvp5jhjIlWASI17+qYiFxBaWkMO7lJlklxiy
fLfb8eN4UV4E8wE9E+JT1srmpRzU3WSfQ3tUyfVmmMjcdf17j6OJMS0pr8dS3e5q
6UXaWG9iy47NqKIla4mVsigUI05g6hwbkeJqMhMVpuaY7eSjWFf0y0thGFB2Ij+s
hNKiYhS4Lrz2SpFlR4gRcz5NuCE9G2aQuDsXsKDecJ+WieKcF7kyBwCGr75srDFN
ke/KQp/OUN9eQ75rCa3BK3P8NjWLvAN5wqaIet34DtRzQpliIoT+X5yjUPM/p8Ph
tnvJNNaQYbOcJYk6bNPO8COJCRgF/RlKTJM98t7ZP7gYYgJfesm0Kv26RYBBkLWq
u/jVoKQDUdl9XobDDfFnPSlc811wZld5Yae9qd/DVwEzj4nu5Xd1AHTaDUg/vJG3
5JZoIcTGXbI8SY3QY/yvjw/qZYS63gRS7jZvvdu21ygnkPexmb2t/0Y7Mccmdneh
j59ML6iefn17oKFAWHJ3rQ6ovwNOiqDc4TYUgp/5fG31xOTZ54wigJ8+H7W+vojC
1qnp3R/30n0uBZvs5aP0/mYEFFnHN0LpFa/yKGgboxz/08xAW+sAtTlimwIP6QCl
JnZePaQlFjZyCKIOtqPBzpQRTix+KD1m/nPcE1RxCJtKoTFIxvIAtJlzjdVQXKdv
3+OoI656YhvRzf1zrDUbS52AZz7sz0rMDcg1EBGc00x/DKh0FTQUbLdzUf1ktoPp
hOsyR37zg8qXvwqfZGgcFvYOsqOEU9q1X+T/Au2b1pO1Ta0KR9iWzjxqBxgwkdh7
Fw3UqSotJdIZxAWD4cwA9cK49j2Km91z5VeAw9PoxOnz5aUdY6Bsuw/OAiEHYl79
AstrYe7QPyqyDtovsEMNhgkuD79od1LXZkIy5CkeHNRwZ5NFI2zdrghfbF8lI7nV
fKyzaMIGzk8XhGSLiTGTV6+zSV3JMAem86pijLsfiOTP/4eihTqQBmpeUIg4hycN
PIEwPHaxVgaehZb+krB9Tz1jqjwF0JYnm+PdVzvSCSH1Zxy6RZ+aCwAWsp5r4oTc
aYhbyTUMMZtPFmGNkUHNfS5twgKfieNZ1nNk4fHBEPa1t83PIpFtk619CjJUN72I
WocBHZl4O2TFnD0rh+Uv51nooo8hlZoaUcRTQVP25ZPtK34c16+Boo/nl2dCiHjg
uDvaa0iCl2nk6JOgumkf8Al1zm0VBuyE1R6+psdK1Fz6HY9lOl2+QEWfZxOQ5q31
D9b1+ob/zm7xDjZf/iHm1pww+GW2PC5YwCEaybe6vyOO+igXdMwhhxTxVkXJyyhr
uo/mpk8aCBFLvI7tmhIC4PlIJm41CJG9Yucw1RXuIQi7UTCtU6l3lNFv6mFl+E27
H+ZzlWXusC02oNDqV148NR2UruNoFJaHAZEK/ZYyzW2XugCVlbEnWcUMKa1LpQd/
dhdOrCAWwktlSKBZ07oqU0vpxmoS4qIUavKI/n1cvyKXEXBJXdzqrYlcZgkfXHHt
2WJHa8j6oUCxor4KuSqBTCdihyfsc+SvOqWwlEd11vcVuz3YvDyft6zezbefL0eE
Kzp3HDfjTblBlZ/TDHv+z+4s61swMoX1ZIlM5LISoEunRnS6FMBER13ROoQUuXoT
qlHu3bapdp6oFrvp68hWxVWmcBj4d6eviBw2UlrcEGeYakrZuQai85WqKvl4rZed
TLdHFAU84obL06saeJFFnwkFVpLRxJfDilghCex1RVHy7UpxIKdW+UCwZo8d5VQ7
Y84TaD68NRIbKzbu+L+5vP0XUvMBZeSD4b57Q6xb0B8g8lxOJm1BOZNabSXjkqk5
vPYqtr7rF21+AzFPpxty9RtVyyHR6Gq9Ocw6eyCW64+rd6gt2PjWPa2TVFMViYIn
gs/pZe8nt2RreTIT+7jUHmYqaXMuq6bIWjm2Cx54rdGAnJGnEwRuWQyCzlL8LktQ
BFYr8kqOIgr/ErpeqSDQujlq+d4YBOkd0LFmwwMk+p7KgZ3oqBzoHzBpJXZvwoMr
yBD2tch3HW8DwlRPnJMAYiiwgDuwA30YdQjfyc2QC2OcMqxMXwaRpKxzStDOJ7y1
71t98kDRmGOejx3XBGQMozx63Qh669F3JAULczzztR4lQegwal73fOpbSkJMt/Mw
ZC6fgf+YxskeIU7v2vg3fKHo/QXT8KKR0v2gfsDxkQ/gf8n5nvRgHSkTqj39Oilr
hXI/3FsElAAKwkLhka/dhd+mEmswtHpSHOtemCjpFsQeqetDEY8ONkUIy2alExQm
lPkQmEw75fPkqXjo0SRT0LQzoh8PHUTiEkE/YDCfW7ab5WDHHk1tQkqSO/dJJj7h
8m70mZn+bHbxgL8nSQ0h71wW7HIWxHFN6fAequeUjSAK1Lwc0deGo0AliajkTvNG
jiwNHdk/cUAN8z5r08LH4iMwOzEW1ClTtbbDNi2qE7iWt4Hw0oEDZ+HVX9rTl5l3
++nlA5HNioFPAuzdKJ5fXMAFogThPN4nGgx+NusqmpLZzRq9wnrNAgOsG6ZPGP8R
oGxI3d+c3Cts41XFfZY7A94ZqLuB9izNxX2xzQyTTaB7pJNe2pe76RxCjN59Ah/6
WPcnropvvSWnHGm70X0RPp80x+VOEiEmIMhz0g4srWz6j0aKoGyr7GznY+8Emwvm
G3y93Fju0JbqB5IXtrAppQ74Hb4K9QzlnU54dWQim8dAX1S8NB2fphvlTzW9Lxps
xi+SGr8QIHKkfTxBA8LT32n+S6h0Cjajapbgd0r0oVmLUDelkcVI98ef7dudeLkA
FNqRwpGpjgMzC4gp6ujbfbZHsjzhoSvxd+zw88IhyXJuC2W8Jua6uDp6d4gw/p7M
uS1HsGFfwZdNHQ4g3l6sQgeTYhAKlRl5kvb4xjFexqI9c7hSeJvQnh9kFoEfKTND
UcQ3MumZ9PvGVzgNzR15/q7vUzBxP1gjrc5D04vFi6ECsPR0S+r2khw0n5MVMkcY
m8eIFKLp1zhPInlUydUHvsNGQyt3rI10Lebi/pEq/J7xn26CircgCRxx5VqwFDTZ
5bpp1hJa9OH7xhqnI+jrt1WDaahvM0BVANPONN+yGMNRz8GWgnN/9i/vhVB3HvWQ
G7JMHa3iEu3Cvg/xG1Mn+CQ5bG8XLkbaOZMoWEEfybdFyDFaO98RlEAdbhv7djzf
LpM+7ZL7K1CSfaY/L2c7nfAgHyle6XuF6q+1ODN7nldNx5ZrosAFWzQiF4mER9pZ
emQSTUba1NhrpJkDFdks7OD+Zilm9j/B2KzVdmaEBtBu+6nUHT+lmspo5Wx+4Ql+
j9C5BL2GT7qJVCs6e7+yu6iQyMjnFIu4bULKdTYX96Dkh8oZXxu9yxjrl5Mn1CQh
EIDqxT7TCnVaKjyy2AKm2Kcs/euXVsDVWHlNSMy0k8Ty21r9RCiV1ozTCmrWZLDB
l5gIkO3PF5Jpd5S7pofA6h/KWDqo/H+W0yjJMDflfIRAkU//DMIqP0tYxG3s/2e6
2X0zhJw3XfBAUmVKGK2CP7Ip1NNnEXZTaVL7yGAnsGPhnCcqAbUYLwpAReCRou71
ZWS/fFsla3mkjeJNb5LTl1PoXO0h6fhWagqG83isCALH3oTWXmeGnEw+/BsDTUyO
2EG1PJ1jDEI0c0uTXHV+7N9O3hJfj4XVDL9JeV8QRefu7mlmZtgROKff4owB9v1I
F0ZTbwZ2X29y47ajH4f0DIcQJ2mLWomo1ZeTuieXkuOwBzzX0EB4DD4ZOcLoiwRf
4b/B/8CeT98F9ut7XCpI0dhG0+diJZLeWpq6LgzadSoa+HJldL98snUsY67OdijR
IqEPG1PEnQ0eMAA3+I1W+v5uEB22W/cXN9kRwsahNjkU1Lb34wupoihIwgOb4/NF
KMplfZZv32H9eHdCfDDRx46/GANKMwKG9vR/ayTbP/V/Kb2xqDGXwKFSyVVoZAQJ
sev6ITQh9l8ouMVCm88EfzGR2ELQzh8w2d3pOi/9YDdITv8FZ4A0optyxzym9DKB
ULDYLxsejPuvTYdL3uBRirWiIJKJJXxV4Z/Md/49/5AGcME/e8YH90V8zizoz/Xt
6YDbWQYz+Mye8Gae28uopwYuvVHevyFxl62EHXpnwAoWb3IXepqCHg04teR+S1hZ
5CSSYqlbOpvHQA8b3BzWW+UzAn/isN/Es4j5c/hu09U/rJBc7/U9Bs8unQWuVKNH
fkrPGQJ6ThKfy3tEwjBmSfB/MMPBpeGp4GShSLA8E5W59OJz0weMrmUy8dLehyh3
qms/OOOyJ5sqPcAUEHzxJ2Ma2YPHDVMU6HjoPPu5YSu7XCI1i+ZcNEdqR2zlB44R
GaBEkmRK/zwxk9QgY8UPpOqO2F/BnQ5DD9tHCdLT+lQXi5V+71FAyelVcxoGsDKB
9fTdn15MPJCc9YAUn+7fpHrRkjaAnC0kobjvqiDry/ft6GxFSeWRMiBFkAHi1bx4
Jdd8Tq8Lg0x+gTaE+4k9A661/DOMG+E1P00qByXpEaDXjQL30c2TiOuWd7ZuknR7
mlMGgxkIjtyCxQGvSrfcIlERGPdJ6fKpT7C3NPgiZDHeMpJhmQlAcUekdEmj7PpA
u7vPc3TjsQrh9zYX8QL74UOMD8j9774eaPnOJSW9jiOJh3jD9eLHWQXwt8yCC2M5
r7MUSXiOAeHpARLi/XQDk9BticuK/y1ezdaGdNbD3MyyZQ7vjlq4Xpa3vdxTbVyu
U9b1XX9AzAx4m0OK2LsKuao6F0sSFxblO6B32+wh4FWQAlQxbGDqOSb66MbOdtmD
eatrrE/1chC90p86OsRqsHYDPfbSVDcscqnLmTzCGHLLQv1suj4dUDlVDGROml0m
OkJJ+I9QbkJ0Rx/iZ5hRvZZF3yYundl4jI8ePvppQ8Xrr1WGUKkJDjwL0iAO0R7R
15i3TwyOmNYIM5aDPtVVx5exRHGtpYQyeYswkWpVP/5SOqpNlKAAyRrFU/OVhsFm
BjN6HReWzeoMvvO8CTPcr40jb6gBaxrsNVLAOC8aDan+eB01if8NcG5UOWIj+y/u
KZwIOuphdBNUPY2Z9u+oW5OfD6luJ3v4lMI/KPTNKi0wdRhCcrQpEp0ZTm9a7gdK
EnwkWgmh4cbbzaUZi0c1lcVyWEbLTbAidfL7OF9dPmYh4P/cY7brxSkeVWjXHuxy
Tuwak8mY8SEoX9xIbFEsfzvlw7HP3ddEfi69hJ0B4MZHcsrfkTsfESCEwUDCDqE0
UdZuiFJpCRZXq0ucRiYFJFzKciY4q/tHTvr3+pQj+mTYoJ6ySeLC/JlwqFVk47bk
WdqpVUu4vfEp7CDdkPJJnRWkwCn5/8BdWjEfhW0NCKplvK61RzLSSTYVSkrSPUuG
UoZi3sFn3C5QRXdVpdeYEQkd3VXIlONuiOTvbQwZTwf4Qu3LRpgzd+QBh0MtUPx/
Y+N6qIlysBjxo0vF2p83rXoG/GMf4tuJCiXvOEqRiCX/JLAjNt0MXnmoyrgmYcpg
GmklAXSWGkTIVn2oAU8nGWWoGUpSuDLCAH5CANQLsQERrrDK6/Lh3I8OwE9eY031
+wF7JdA9fnUOj5j9LhO0aUBMeHhNcfbOY2pQ0do4IIT9z15+7GNwIzur4v6jf2Y0
sFi0BeaBREHrRQ9v6iLzmKjVzDpkm0R4VaBBevsER2yUfLtfOB2MDbxHknPJNPb1
vwH99Vcrmpt4IrR9/czknavQhH6SsgZzWTawuBMXq/S6UApant2cMdgjGJI71IPE
aeJdhoU3882QtdbU6R8TTC1/TQ8eGs337/CW5ztgavlr3aLo8sqFEavVLQYQL/Yn
bGLlvlAeADZ+MS0ekTvDbnVBZcEkUvWSsUF4LBLF0WHTuN6BYet8apIJqoM9vt3Y
f+1VtRAkBr9YFPzA3EbgN4Q3eJQGtAR/dQl+y/9+cpdmiTQ1dmpySaFalLGdyLhG
XHQKJomreHcTmLYUUU6RDVnoMer+WIk1DHkEfqY1zYgy95aLNfwxi/oCfMHXryXM
SH7fSjajRr2KhxcdOuTLCD075hcbLuv7tZec52zqTcKdAEhb4W+X/bgARP4/wFYp
qfSC681XgdFlVB4kbrhfmII5wCLQ79awRk1bc6TasRIlL46qTgLtYTrTssuQfNee
nJC1qlzTg+D65nKaGwDxgDXm02Km3RTc0UnlO+0yildKI49XAIMA8d+r/GeE1UlT
/MtOmcdm8U67fxBjDJB16eMUkILk4GKzyk8MPybs538HTP/AHmKPjrtipjQtzxA4
YotyfUyePgxfBV2KZ3B14nnN8vqy270utgL5xPRsQZ9CRoPzSAZLdDN7BDqJRX8y
k1TTHh8aLATUWQGhGbBMaFU8d9mtf59Kmc7cGv1+JNLxyxddOHEG4NakS4dwIPAl
a9tZVaP7xIXxZ9camUf2EW0ER1gMHUJ/9j819JoBZEV/Z46xQnxK2RbePVqbLM/9
fBwJlazC9Qcst+GUui4plvfK0xaMF6QgkHxUAmc+wngymwoNtKP3TFgq+uuEXk/u
61Nfaxf9ISZ5EGt7ABwEEedUsLUXZ7HWDMFHp93MIFd0D7CJK14zTowadHDOSJ8Z
IT4M7fCL5wXjdClK0TS3Erg5UuIfYU1shm58nvjvQVayfCIXGyer0RXURnjrbEbd
wzmmdJpfw3W7cyNDwXxIV4wGdmYIVxbfwtXMtJqOi+cS72sSzLWNVwTmz667CRbJ
fAHN3EQO+WR3Hx12BN2fgot0ATH085S2h+oAhFOB+2d0apgx8/tfic1JJ6hXO5B4
axHmItwrs6by16M6GBHIhcQjIODyuf/UPymB3lHGiIbI97paPpYyWPbvoex61cYh
L4XLBDZ8TwJTXm1nswSpwKGQMCCehdgeFeCI8Xl+Vnd6DJiOJ4KQF0kOD0uSbSWd
gSuYN/1X5/OnizhlNyFFLqCkChvkySLlm9TvMFWYlfnZvS73YI7FxvpUZozra+M4
o1O6f7gEBQ8mjz+pl2fo5TyxHQRcNrqUOeZ9m49AAkba4kZXpZFN/92vUfeZ4CTu
xLH8Br7MLRzKBrQ4+1ScPdnEdhp30u7oxmxXtcz3GxALj79/+zuc1Vw5MCzZWoMy
wxqPP9KBiLZ8wpBcvBjEwuZ89NtsKihAi4CePl54E3p/X4kNJ2x6mYtFyTljFqPI
I5+fQ/DEDI+AP7YqdVbhCguRWVnTw4pZOYog364YWz/Hkq5isOtzIiAiwAiWWmHq
skb18XAq9RUYM/Lqg11uRpmBkv4RJqbrWw1veUVWtP4Ku84pbTW3W2brlqicuP39
Pcja9SsQHEn2tXY3JTcBW11vv+rvxT4UMovndroTBz7Zb5Wg/2HTYPv40zBdAqN5
2VBXzxOPa9Mvy8qdlOCSGVTtmnXbdxkERDs+DfbQdCLb+kp7Z0xnn7FhKQmgLi8H
3RTswRQFqoopx995AO0APmIOICwxXOgYvSvLuD58HBGvJHeBcu+Os75b8JbEE8FR
jIzdk0L4UvLYnVqhdjaznHaYvFf8OQmtMy6E5nwpxp3AvFYqUWSagQtHvT+oOYYJ
8Nk5ahsAtvSLftegyi+picNq7uBaODci2j4Gtzz6V2lR0BHQGmIWNw4Cf7dXjoGb
+VG/IgzgENIQRco6K0a4xhRgFfb3lvl22tClSEWuNYCgVlR7vacwHiZX8sn5qbUJ
ABezdDZjMEBaJZ6D2Ek/IZM4yO9LjBLCNg5k5nFRoSZmiZH9ZDVd/jomoCzaCz9G
vYBOqHLnKdAaQeU3H+UqO3JauUrJopTUEKz288g47X7Iz8IYdfZj22covFMNJ/sL
rHjRELOoSBv/Z/Qtzfb3N5pmniPf9DztWf9zY55aiaSs3fyTSD9ZW9uNalpeoiu9
If07+Dd37gbOS/5AX3hPrQTCXB+PoEwTGaxLN+0BKGwkYzuG38sJSWwLFLHlHfHA
457SXMV6kN+uML5kNZcKX0AIu2rU2GwBpxJ0aNMwOfH9O1+p4hO2NyZp+sHNkoko
WriBz/83mIO5jGOO3xfOOT8eto9VGKZspknPrM99D24uV6fjyFCBc+NuQT5V5t2M
Q/JRTjXx0BxXHNoWP15ZQwuWUUnauZUISX+gXtg5IPSGglztlnFmQlne9ofSWRVI
ScrkqZZwqmDo8fcbkH+/J2AKrRyKcI96P/SRzJ4KBNwkFvK0x+tbdH4yNJf2SCGM
aAV8FWGDsHx0KeAGHacIIyZnLxFStpBYJkVqz7MiFlMpmAUTttHPpbworDxuS27s
NziPXpi+TgkeU/diBsd7gNj0LVx4VaX4FXjo7EqdJSWLI2/nwZwEoUrPnKp7uoov
Kd2sFS7eFeeZWkle/FzYhmftAtBAA5XZZZowHMWWlrZf2cCwPIHfqk00hKzflNa1
z/9aCLlgJjYZ1b3EHCYK4+hfw9/9VvWMf792CblY1ScM+3YX0HgyX8HhZ9wlg9bx
ZWIK2Fl8xOrcW//tIKFdAWpSY/Dju4ZFZxItIlQMTrFjcDr5W5LOCCXZ4itUAB7m
mVcCIQjYc5Nn6oFGCU4WPjqnvCbkPa1Bvedg+RU6JWWZY4fQBaMrMZUZZ06/+DMC
awUnA6oes/m4anMdxqp68rGqQceI1vMQrVz46wsVT/D60PxSengGZz3SbGN29/ux
XJIvlUrGDqJ85EtwUtsoIVZsYtV1EqQflpF2cBF3cUrjoc7lX2e+dRFoNdOtzSi4
YaKMtGpkRSfd6tGS/KGSKY4BN8xzdlwyNHUQysbgiXu3JXAZhq59XF304CiGnSck
p3wI9Fllyn0yctDjFUtLsaHgAOO2jwsAYQNDadxI0vUYs9W2tRBPRuPE8BpLL+PG
FhtVlV29kKkgJpHba6UV4haaeE0ZYLJNzTPRW30bOoKPWh+0j3jVJMcBClN4793i
Nl0s+bW0/FePD18EQy2TYiR5Q8yalAmxGXkCZecLb7VOSjjwrZkft2KeHOkyKqMq
YRPHFU7a3xQuBe/IP7+HdiOPUcJ8xhHf8XO0hy13/6XqTngF/lYAn9FOZd/JTNdj
5V7Pm96EpMlQfHdBqZIL69BqvAyK+aiRoWUcoAyvRG4sLYF4989//lniDhuy/n6d
iFU2wK0Yc8Pg2ilZmn6n2yjT3MS5nrr8sjm+CwuSAS++kupnGWsrU23u6wzdSP1U
GAfcehjB6LoUu9pKK6JYjK4F5F6CKvH2R1glEhJesbWl3tAhFb83+UVLqhDCgkwW
Y66ucRv7KtS8ODXPO1DNSxpJsxd+PtQk8Km187qstcODWKNo71LOFXONTvLdRzwu
dOuKIt+kj/cWqX3tAxiG49eEOo18zHAOJQebjXIFwwK7+l/0XDXdjqvT1Tff2dPs
BTGxlXxVKBjUXcWg2sBxvUtaEE0ksiFU6bel+qHrijahCfg+f+mzx9Ct2kOPXNMl
yLL9P9kiIOSxlrgwmuNz20sXcQ+b6wF87T+ob+TPiF5m2G4o5ymbM69JcVEuHb5k
K8EX/tVwxE57JpazS0RC2pxxoQV/AR4G8w2DjCX4eA+zbp7yEuKqWF/FCUnbnDfB
ltnT0R6kRCWik1ZQ85oOb7L2Kb/7olBG++a80sduae+FWnexi9L+2wKURyzw9zc7
uu5jA5Ailcl4jSv8bYa4ZZ4V8f+zsbmxmGTpmhsKXgHMGimqWC+dWfFNVLyl9/jC
uMrfvU2XCjw+o+utbusozFwZDS2gNmyCsERI44Yx2v8Z7bVuoR8/gbdh6twAup7j
2D/5vHzDhrshY59P6ByQ4pyPWoH0ZzJuuqv8pUUzPKAWJEIspSBkHimQJbUAqbqh
VfB/UzDXtrdHxwdKrgetES9lDFdAOB9xOZQ+EqTJ3CrHzWE2RhmOdZygxM00pbei
+CrAvz/TXtWZUAu4+F0hIWkPpfG1HVQeB5bY384dnGLwh6cbfmIgYfas8O/zSfYG
b0ufe9D/H6XVdtCaHtbkIc5ARCAEwW4OXwlOpbuKD2hwyU/EsKm2ifKGhG3e+Em5
FgonUw+lmWnaIyf2E9wIw/wOMkoIlwtTpOyASXuszGiQ1HMzgjsPMVqKPmaBiuAz
JABPeP3ClhzS7kgEk+9HdLleFc7kek6Mkq2pRGh2GmHdE24ehSkMGBzn9Sa5n7Ll
/IltBlhRtSAgQCQDAZWXZYr8pPqMGAa48vf1k7bqbgrkgMPLIp3k9pSyIL17B7z2
ZaJ9QyOzJNVhDt2Xz/lSo02H+Lc0uGy80sRg2qIVqbRu7gYPukn5yPGmnLSCqeH1
Q/IZSfyDae5dXDEykXCZIWfOm/s6bcHdQj7K7Danf1c3/ehQ5ieqi7LyUT3GXcYS
J2M6PZ+pzlMaAHzpD2b+t7olOPHUl+NQYEFoxjxNm+rw470MU34mxfOqxsFEE84B
ep4AtJTWSwIBGk31+ZwcX8CtvFOrOK/5QuiYk5GmbvtknXRlgW+soiXCdGyX4yrZ
OlC+2AdbHZ78YwSjaIyt68PUI/m+xmR+eY28kOP9HWKFHPs+zpCvnMv7M7BBv/tg
fSNAFsof9xL8gPHpO5HBwUEFgS6XZVRZh7qRs1j6wfwQJ6+0wIx+PCbAVGFrNCa7
QcDy3WxiJ2rnN3gdgEszc9vq8aWLzCTpD1Bfbok+KztkMlyEZPR1Dj6diunf9MBv
wQYw6Pe3D2FdJ9lup8y+pPbKs4VCM/lRg74dxmVk53vGUcHllrNZlHCofEPzz3j3
0VTRCMHXHz4SHlIXprMFnSK59JuYT/0ggLs0r9DxHkdE5QdgWm6v2PxqfvzBzlkr
TXFeHwVXDVTi51yNEkq4Q+IOlOGdvstYuQJ5+t6ZbYd/Xe3vU0z+KT4aq0XgOXIq
EYaGGHSjxKjE+DCSlz4Qge6GMCPV+jvu+PQZqWm4eknSlcIUGR7Guk4kAl8jrFth
NFpeGKzvMafQRVV3GV5YCufmsTMSeAL08FzZ/iAc1YZBgowfBG3nbKq6iYDnCndM
gTfoukQGiOGPDsQaLF2fj9WQQV1AqvIZGI4QmDRdsd2lOAL8vPI0Vws1HfZFPqS6
IAXqpzZyC/hwEzABFmEw3XH91CRRjefZIsd1grg6N3wg13omZJYp3jY5ogi7UXmB
9i0LM3D8uJIqR+sbGwGVVcQSAm8QRSl+yo5uSZodTJEMZyVsmoNkuyTmPAzlwz1M
VC6qORP+bdJBnkl8xfOa/PcKH0fL0qywcoRlXvwJyh1RYoHGf/K1u4h32CQTD6ss
KP3L+GtjwXzxB/luyJqWZmC25SOpkI+nqFt2TCHfGu0mrgCouDATKt2NJyPAdqzK
e9za0GN02sa/tUwA5Kmh0sIELuZxLhC6cqovbHUptUXFhKTYeRy4C/Wi6DV5eAJe
SwPe/OcoPjCtH1LYL/aPxYGi7/tn3VG+qvOYWqZ3HXz5n8Ql22E7bkFNBJLQspCT
cYyAJKa9V0hglvCgtrr8MIq7dvPIGZxBX4rxddl2Cddk01oL1cp60DA1HFovgHY7
MDggW7coBcge8+rQ6T2XddBuDGR5ZKL8kBZfNECV5vpl6GyqX5Nzx+ns1GPbb7Ae
eqT+BhVey9y9gAzyuhG8O3YzvFenaULVwcL1YR5KLPZJeZ/l08bj5mmrxv9C5uJn
kfxMzNxZArYqZ9gfBcwJ5bTTmljyIp5rlBK5Bc2pZ/Fpkk5gD+05F7Bn32Ry9axd
wHN831QofA1xvfqMiGzEn6VYLtlw3u386r4g7eznrt7zCHh9byr53AhusnwvLrTZ
1wc1iRS3Dl+BII8b23ji2HIdOs3BjjaiXbwZdt7u8JmskKmTzQw6OGUFqiK4uJch
0oXfO9Blct+uwO7/1TsF9bN2rLuXBZwfoMEDl8kBHXiWmwxmUkcdQvXL4W/ySiJX
aHUpPyxxqQN0AMqV0Ems/SGP3S+Hp07Ve1riAPQxjHY9EUZb/ONIBw5UdRKOlmd2
VnaCDlPHjklTSEacnhSUYIweZJpBmGehnEzqiPSKKydBc/J8DJaI9iRyKHKB4oYH
VnIIu+WBBSFgsaQ1mqy2910BSGKSwF8veHhunR+E43ILAT9gWOw2mozEaG8cZ8/X
AQ6eAoTBwDyZjwKBK/IlovYTbO6POClVCKO0w2kmAH8g1ZU+2SMTTeXjacVNDGsb
X8tMBm3uVfDj/zmih2peJtTy+G9G4FIZvbH47FDAgAMSf5kVm65RAG1AvnC3f4jL
J9grBkuPQJV5AhEKzA6A/Nxlbw/3CkzmpVAUyng08GRrEDFDwP6mr87/gyuWxJQj
7VGlAGkTdeOHXuDAXNLpW4m0torF4yp3Zj+AL40dBLZoijcI5G3ZhER3QtJ1WqJ2
tLTVM0AGFaZvbQVVFNve4T9E2BsxBQGC99u+nSw3qzBtWD1Fy7yTSvotG+4YfpWD
Agl1o0dVuAoV/LdGkwKhuKTYCaT9x8pmheOqSXqWEL/D2L+lRvDGiVzulC4ZVXXG
6evwlq69jtwe3nUIlk6NZvcuufQUhAMaFFS49TniFMdRQFL+CHnGIeTI9FEBvq0R
i06zvXXt7qtk3sSYxC1GxIttbki5GiKqMAZ0quOl+GssKpVkyVEpTyFAzHIK4TZf
URyHG4bs7yb48tFqAqMw8idRk4UbskABukYUZetl2LRhJS/xJcV7NN3Z+q9s44gV
2NCqETvnk7Ayy8Y8/wF1Lu0stRcABIOzLsAZPawXPBaQ5QSfMY+2AorRn0UqP6Zk
HAmrIQ6PPsU0cIuO0P/XTKFcSK0d/QrGVXhaw5hNpIldyUqQJVaIW9SkRnRnhaz5
diBc1tPoZgSV6A/au2kLl8MAChQIoWlGSLxTHr+qQq/HkWY58Kv2vR+Dp62L4brj
5HNIRREH10McyKi9wt1dPQpqitFVABnTWcJ1OtjGXURyxm7oiq1X+CGl8hQ0Tjse
5w9Ktmb7DU2T1GdKCmaKtrmxEMB930N12MrFt5cmoTN85Q1vAy+dFaYZzyRcr2fv
kAwhAllFmZ9JJ1kstTiGmLKQu33e+tslOpknJPgeh1qRi2YRGsEmwmitYVesiE0P
wcU5IBxV5m9q/2zNHS6OeNSKhiNh1oaUlsHsTgWpQ12hC8UZqec5Hbw1B5fXxZzs
pVNL9qlXDmY1Jhp//3891Qc8TRxksonfcGNkceyCz+9bazdt/FE40nt5oJ+244ex
EJ4lmWzSULGYkejZMJadEd+Y6cgJl4gd9xyzgaiLj825JjyLsItCvXo9nbTZLBAb
VH6heR8hzkYHHhFiW0BPrhzuqgn3cIAjRwE6IdxuBIYcBV5/0GvrjzFvaC40lArO
KxXvh2wdf7AyofOOpESM7sH9uHbqpzdMeSE+z10JSQxiIG2yCfgfa+z4imvzgfTe
NiSB62wsBA7qkKybE/ToXqUq8Xh/fvtsGOIz84ngsr4RJem+IecHvObIqqfm0ymz
qpQMXR8GNtcsrbJLxHoQoJKZ669mzGNBBmC6z48dDeVerdsO1qTBFLOKWYF61vWh
3kUtayJbmFq+vKcqPLQePRkhXw1RGcbrYUOLUW7RjMD75KKLDhzAV63Z2rAGEg28
mZW63zQceUtEpw2UV/ofCBpKMp7gj/o2G4lVaCEgRFl0JzBG5bCpH64vwNHdDQcf
8//Vs5TdKJiq51SrBeysWoVYNIGEUJxXoBIUivIfs6gCTu0tnc8tiAorDvVJtGd5
FMquvW7tMt81dqTjwIpy+MLvek9GppPra5z6RoTKFWLkKrdemwwQqkiANgAgD5ix
tYyDAwjGY6v2JzPxCh9Hz8MYIRLbgHxLxIZ5PnVIwPptHrMcfMij+q5dyqr9GlB0
49SJ0PJ7uVC7f0ln66324tlWBzz7ASUFdh+R/OCNC0n59dS1UcktRQTnoK9TgHX1
2dvx2Bfd69qt6iAyE8//wgVb512s6ORAdQhZIMWpnydJp9y5My9n51dRvMvGxk+C
AiwzW/ovQpCDYVSenzsPF4YE4gwKPbKTZSJRAX12HJPAM5h9KfjelyDzkgDVveNI
m18RLM08qxQW+M2Z5xjvuj43rphluudygrth/O7HUsSaM3TKbBuVlomx8ttNG8In
o3X3xOGlvBbJPmy8ARNrWk83maXybeonIN7ADsylxTYucvEw2BUdaW7kXCW4KHgP
MtQ0fxqq0821+M3l5Sspxl0TvD2Xe2IbcCGsghEuai9GLlju2LWUVOx61S2QJwgm
FCb2P7nkoAn8Ob7oFy853k01n/wxuRJl+UtgUvMiV3teYpZ2i0VfAdJH9ohLTdW+
9qaF1yQgVu09z/ITozuBqtzhvxZ2nLtXJIOKFooUvIRN8eustnMzIUIhS6QQN8rI
4Yfk62luW/cwQcpuIG4ARZGVEEdekV+hWX/Z78XTu0R/tyMvQiXFBvm0PoBwfWlH
ibtanIwJ6XC6rJPUW5VJsYUDSwHLNW82MZcmqt0j/nNuhEvElX46UaY0GORzUEcs
IJEVKJv3wJQpob/mS20Sa2AZM19q96L07b9BPBb4XQ7BC4+MZEy5OgAEWI4ehMWy
gZQbF0vLWD2poi9+d8fVTijchriltW1MN3xz7mLUEz1KeY4V/Zarex27PYxRxJEc
5kaGQFTryjyzdlHvWusSbfweCnTd7CXOhCaJ2ZZrSe/OHygki/+hzh/qMgEtqxnE
vaAp/PRd9gZ7RStyDLPA8u0OVF3hgEVkh2naMB3lUMHz47rS6q1tqcUbtEvfNRJg
3pXfLhWOgMiJoEAjkiWbstIkWxmE2GA+BaH9eLW3MggFuFERw8LCVMX5T+EeBDpC
9UBUNfb7/HPYHO9vVjkgolZrFMuNtkeg+EXMvvSJhnm/Q7cBXJodRip5KI9whY1p
cI5Z6UgYMlgntYQgIS9bvwsP8ND+J2YEY7DjepAKv9AxcmeLKga3G8paIi9tKZHF
Wmyq091qVNSYqZ9cyMfif1dgZsEC/w7lJpAv0vt7Hojm8DAZhRsdXDBGFaTYSbF/
wYBuu+pGxs6dmJG1HHkgNlA2NfYdM6KZGgqvdu7klq9/cUa4NEIyPH/Kk60DqhiE
cYhDN1xocqTVCPPYrT7ata9Rjsb9vti4NZlBG7xMrAz8wsO/UljMtBM5xlfff42E
ybsJrez8HFuQb0bGZBEVyTu8SiLdTypICol8TFRcxc7m1d0CN+cqp6+7WmcM9Gob
fFEoiUZX+jAfnsWmwUDl1PlwNSaw07Zc208SCQ53ccf6n+sUs4Ve+2BUnYomw/Rc
Rct1KMG8iNMDn9Lmbp4z/+mWlwL6O0g6oomJYBhXFhyU9WWuhOt4sUkx5e/8G5Hu
+NzrIUdc96R70fwJCHJ79Y50X/KIc76y+yfvXQycuURkcxWfRfqrOfwotTonV/o0
EijC35miGfgg0WQMj6EOCDq2MLIF0u8SLfvyEGR1jCql61h3t6RN7V6LCaFBsWph
3pyD6PxByrXXdqV76B150J2I0zvx2kkI1hppg5hkjiX317nzgHfTaQFT0u9R5em0
a7c+eeauWqUeQf68UEI4efXS5ATcVozRqbL+qOSycLJQ2JA1/AM9Ms5BQnqDWv58
jgn2q13UyoDie+u2y6wX13tnHGhPnXv/tcv1mNKwv1InMZOqqUrd6MpINhFaiCRz
Eyl2RlWcTFSO4djfMnH9iLBX6PXd7/JnRg7Lby9tXIUf2oZmz0TodKYZKBDmjq8w
DxyQFaxFg4tEfQwA+v22v+IZWUj44rn4okujoPBayzXku6vbMYnRb5bpWy5pM+Uv
BzGOmK78/wkDHeQHOJWUTELCM3Z2zzvWbhKNkaxBNTqlpE/nWwhTsYjVQrt2utbB
B9CJ570DHnQDMTRbh58qB0PMXbxdVXjjPT+YOByeaMCspzCRtaLnTLjkm6rslNNP
oFr8NivEJghmaN4EG3HrCzc4csawCxEELEEWL7HCbS385x4HRfVDpdg0h5qUzSp4
A2/PtbyrL0rqFUsWrduQ+otfnAiw1O8aRjzRHXtQwwRl7Y+I0/6HFb41IFaJT9HG
CXspxOGYr7M4onH5AqgK9BB9hQH+OI1LYD4COWZzNe06tDVCt0gB+o44kczfNZf1
3piushdp21GWVFaIWX3iZV8ml1I69rR66Q08ny88MVXBtvS/0E/DIMD/lxJfZjuv
6k11ahtnnxYzX6fy01quXKM84GPHMBlgl8/BScNONl/ZwP3uqtE5fMdvCMP8gYfq
2soP+aIJgp7KLLhjfzAe4m6QGnqRUr7FbEGgjujv1961Ih9SMeX86sPgbK4H1uTN
lrvgELW7mSxe4xClFbPGEV2kfSjCC8yeFF54swJFIy9VSaqhErmp3X+fVVes9TC5
H7ALMpYv4xkJe9C/wMwFvJyZs9CaZA+p1tfrAPFJsMqX99jS+mQIYIMbvhHw8k37
Xw/HwDxFv2eb+kj1fAohw3ycxjSDfJCarFfnRbl11HgB5wQJDUkKPe34D3kQnXUm
MM7lORxG2TqknzSGif/V+8xpI5/w4wFrHMr9UuAiCfEailp7b5Oihguwmmo/1qZ8
z/rBI+wfPDZ/Dz9+GXrvCksEMgV0b9/RnP2lDSHIGSeWGGFp5ugojmhJVANM78jR
w2D4LVOE7INUeL/PlyBCVSeTS5xsvoV9tBGKGgSsbx0nG90thxg/hT5pK26r4J+k
Cl7rsLrhicHOM3CAUxas89ofsooiA6DW8wV9qftZTp0bwyc4ILv/SX4a65CRvALB
MrJ4LatD+KExS7y/CLwzckflzhux2CkU4AWPVW3wOpVkQxMi7bKfTO1F9pld7/fq
KKQA2OPyuEsgZ9YJ44BtWmzkRUm3tun+Jogo7bH0PLEJL3Hn2BfVcYhesu0bB49D
dl3Ejm0j8PM9powP5T7CxayXjUfQ5JsM6riq7V5GxSt33QOGejPF/caI3xCNM+nh
EmyiAT0RM2roskiShC0oQC5tp+3xQK54yEWut9CI98Apz4B9BvxcKVsUZXm4d1Z/
6+EEmuaYj8w3F66UK9PLwLUihtUDQG5Gx7rErlwW3P2a5b3r48v0YZkQYfkmYJqu
FUCmANNMN7lQ+rgTleRmzABvJ+oCmoamGFnshjg8HSkAwe4HgKwXVIVL8aB3XMVZ
zgF66SzA30vDZzXVM1cglqy4pg+qnWm5Rj0yd/vWCgJvPCx3AYv6hsWOEkKNB7Oo
RJ2EB1pjjx45k46xbQFEY98NkfgqfLcRkJVyBIt91E1dnCEsHENLNsmNgRpUDiu5
ovyxfQtyJ7/W+yB4Xauc3G8InN1vfIa0kbM4bsaxSgfZ5eLKb8H1fXcM3INxzUAl
e0mkXM8fVjWx1VeBBTze2xWXIBWrIXRvsZhOi3plWn61sinZ/LhnyPccl/lYngFi
5hYvH43lUjrOmSndDeTdywAT08fAWL1/oSfpHUI+MnNfSN5Ge5LIY3/lTOAttWUH
VGUNyGTheqhw2fHwD3YZaQq/ozNt5j5fwmD0wLvZDl2VEezwagVHYcyu6cyvZ/tN
ImAA6klyB+vbZkqwAEixPEsLz3GNWjMtItakzV3xzmnuriC6zeuzitD9rlHNgIjv
6SKDT5+A4q8NedwlV6aCvrsI/OzOpZM02l6qSPNBoN6Zj3AJQjd4toQ5OCFrO1ui
CRkmMvPP2D9hSgXpuI6jR86jd3Y3V1SGQBYb1P4UvViL5UCkBpXT01oxNH7Y4DNq
QkhuavtkOJqWIae4S1X6OEkyJueXkmjRAOq3S8nPAp1D3YLulAF6k3GNxDdgDaCz
pzwyPNql9Urv1RAPxRTzbPWHFU8z8PoRmphCvxFYfMNDJ7EvHm+TQx0xeLc8X6d4
odVo8UbU2fr3l/L2q/WiQ+sZopiljpfp4P2jbyLCD62AnQcJBsb0Yk6WGJsZGeAO
G3K85qN/hmUbSfpNk8GalnggjU2NqTSAt2KeOsgrZHyJhyIaXY4mRj3Tce3+vX/P
zVQPAfESgD2h4BdQsET9gWs8nf8JiYTZ/BSRH0EFwym6ebOFBeytN4NVtNBsN2hd
9ZbOkzxr1jd21otsIGe19JljJ62XXxkBxucFD5L5msAkYB/Ji+hkoyf7twn5b5hv
8tCz6XIuUQjkewFHaicOPr71I9VTViYxr3aLZdG7FMypovDX4Fpknc0gGAiVy8Eu
JKx1IrINFURnEvmb7qI7+yGn9juz3ewmP88q6+tu87qpgFeX4uXEZ6FVpXHrezWQ
orq5B4sTey3y37Tww0TLc3a7KV8dJ/DKi1y67d4ThKzpT6LC2HOuxj5S2nCF7mO0
9arnsWdELRsn/7w/OtuHuB0Rh0loSCvW5LHaoaivYkfdUhNg6+C36IeI2PdvsAW9
yAqPOPi+vb6imzRMMajD2TCzXC3kJnq0W5X4h3T3HBuqiuo5jajaIUPTzmEYcaz1
fiSSI5Ro05xde4uKL/Kk35XWFeUmUK1jvxwAnn6HQO1FgCCskf2YhYjM02I6c96O
beiXiRCAX822QYO+wYIxWAyvpa/MMdTQb8YTT/JJ8eCveYqSlDiZp72hThIc28wl
UHqPdbdp9t03D98V3bPjFDo4e9uhSOHEMDIkrykr3e27uiR9xmnHyn1/xN2eeQIQ
ci2xXO0QhlBr55DUOVjSt4d66rewzDdChzRmBNjTstKVI+tM+yq69oCpoRBY27yf
Oct9otYpb6LgsZLvVPwe0Ub0qe2swBO33sZTyS9NhZXClqtjVVYI3kRh/qr4tJbh
hrVUThyDEaUHUXP9z2+mu3jEot2tzmRt1ic7lgfH6XfzHTC0XWXFEEsjOiMX9gMZ
CiuCOElTzqwnsXJ11WKct63//VJ6euOXZU59P+esQADcIRsIxJ9UB4rPhtaKXoiH
9DkQ1ynohFcL3DyyITEpkNG9G44E6zAsWArZJHgrDKLUj/m/zzIppRV1L/TlEZSt
riTJyli3nXxn4jzMEGrSAqUX2bsdVlFkWkCjvzvsv1xmv5nV1Oc1BqheO/KKudgO
AXYKST97AmuUZOgI8E74fmJb4dI9XrECgiTkFScV0c8+H6YhEhuiaQkB3y+xgQxh
K9Agln0gYtLvLzFWtEYfh8PqYPgcVIbyNA1DuabB/lKLVavO1+jKX5d/4kkdEa3K
4IzKLDjO6oOzDYWKsMMWqJa3WezvncWDJSlSCFSQGcvGYZoaBWzEJ3U1w7B5u7cZ
/YK6HcuibCmaEQLtBzRR0lVbVWRVmrcwe0YXf44J0/Ct8uoA7SYMuIhDB3YzDedk
Ui2zZlir+VR4ZDNsCtm6VuS5mHkThM3fEOKBXjqw5GOC867Uz9uyyO4PJkxrIemt
Gnq/oa+t5CLc1NgAQac4rHZfstH3/1KuwIcxR2X/9Vdq97gQF6y+AP7Q0weJAPLJ
OrIgb0izQU4aAPE2fGzHve07Msfao4mSW3VkZuP3oF9GoJXvSvVWlNzeTddnpIOJ
g7bXPnHI+RgfqkmtCzBYBPGLWsXQsLJjheaFb+KMWF35P6oz4QYvnI1joS2TTuN/
lzNtjOwEnc24QK7klsy9na47c9TOsOF2j7QzgD0fM8qxmdQt4yn4ffAYFEgdGh2G
9JE2RiURSix7vEBmdRo+SitUREeV0npMXIb+No63Nd8AYzXCc6DNU2DpoXg+pm6i
KU/D2CMy1022l3AeAKh/poz7DtePxDIAf89i+Tjet/8lQD65vRSslXvjT7UFITKE
/iQRVSCzjPHBjEFNAWFtVmuLjR3knv5R9GVJc4uAcZX3tm46mEg+U+xHbthK4i+b
NRNZ3abL/ahmXNYZuOPu7CwWTCjnV82cfkMrpy9FmfD41ntvjz6D6+HFP4age2RJ
N3siBGx2jHo+JsvcoHo3HdcasTgi1DujDgDk7byzqvz+s616+Pd83f/6lLHFpQZQ
+LTTyK2umH3pSbLzNdNJykE1g9p1PQpv99b1ZIw6P5+/LictUF3AZwIC3jr3SeRG
9RW26zzntDFgLlKuW4yJs1oY0hovu97vw0423z6YlN4kSfYcvuTEquMVEEc343Hg
PhULkCYnDX9imxXbHJR8AhLaRALPfp+wvZcPs8R8Appzze22zwWdyUGxixKUwGR7
oaNW2TLwKjxP3PkE2ynasr2ozr0RWBCV9YY7PJ5WpMQ00ll0YhBorCSj/9c2M7r6
lNKVBRtJSu52L3FtTEqNlQP6mENK14Hicjb3IVRKjoB/aHduwDIPZyvvs4JSmJnV
sIyFNE09yrMH5Cga9ML6DMk0q8oA5l8jZER9MDlySmV5/jhM4Ad1C8rIJjLc3ZdQ
vYOKEd3IJhTIUm8j/dulvbaf0+Kp3noRc9GmyXSYI7XZ99S48SjUp8NcCcLrJfyD
4sjFWts12aU/oN/Hw5RGV+HIUxmEBiaZgh/tYk86QeNX9Waae3Hhj8NWg0thYhEE
dob6ls3SJr4GGRMzvFjEN9SQf2R4FmlB/EqPmb1/ejQRgbh/Z+jBM5HsKNbHG7U7
kZqY8gaVt232fm+pKivwj0OZmDemZKVIAD8758ys//zqgqcD/q6sUpJwKAC84/KP
/UIfONJyJDX8jeh4YeI09mJA7sZmuKf8XKG6v2oRLO7q7qGtxURexUDTLumpPGAZ
6dI6icz8cqnYrcjmJn/PCxfs9KAQBk2cY5q4UCACMek8cGrZVhEVHEeWHHJ/leT1
2Uxpwj5NKzl82pSnGA5BU2DQ1/J11NMfDBnQ7gPHTgTGXw2M+nrg7Kk1L0b4z5G2
L1zLhTR0pLNgz0mp82V08jdmUCIwIJXXpHYnqlUsxdOCuTF10v8Bko0TGa2eF+Gk
BWkE1h+OTqN1iuaBssCmU+daKdXZNuZwl3dt2n0nDumSbmY7FoOkY6qMmCiEeQx7
lHsHD0R8g2MR/i0I3L0BTqbPqQ31cUAWp+P6zr86o4BuHyzaju2j1JBB6POFkSeS
fgg6fml8N2kpCQ1Y//pMUZq9fJoQueXNwqA69ZNO7tD+cDbBEuZMalgDTMHnLaqJ
i9/hYV+eGkLS8J3PkPIUC57P4juC/tgTTyKSbhNB3jfKCTtbfr+JrRA2sWnbriAI
C3Xa567PyNWC0LsSvPwBVmWJLEbl5iL+atXd9dyILrF2Gw6fKUjt7J5+p6qq7dzc
UVTWlZUkzYUVguMjFP4b3nQF0dS7n6xaB/kZyOIw0DK3nuOmWmbJK6os8cooOz84
FPuc+lzvFSp6izaa6L5hgJOD+QfJ9XhvZKzUfynztfwiGGvmV1rf78qLA7W9rtd+
eBqJue18th/mLG+weerXSy6bu2N9ambnnU1qHLDF/NvCdygCdFyWb2ohrHBYDMAV
B7pVP+VezJNy9nFkeENk53g+YQ/u5zvNR9En44UMCzaL5j9U8uVst/1R7rMv2SPc
zVNyRqSnl0Cv0azoQY0UVDPkGj8pUSqLy90m/2SCUYbhWQb5UZRq9K3sfpcoQi9K
RF+B8S3w1Ik6eZn0cou5X6ibaXEOK3TmbBcovKAZi1nmuP/9VuqcfQ/qm9mcldYD
u08ccptk21UVqnTWp4V6UVIF26KwF0aw68RPIHQG0bk5YzhCUCxfwjRDhfB51Q6K
vtj3Jrl/oj6EYPa5ESMR6rRbMFg0Weq3EfsK1ZxPzlH8PmEV7E4mB2OHLbrDaBqg
vSTAGqXFTrqwSs4wHoy56UPabAxqgBdWFar98KOKB8pkHNFRlq7ugfw98aEMX3Y2
jvMYwRU54F9zZLAVqg0WvJn8N+5+lHgTiUPWWVdKBRKIYmoLBCdYe+VGel1NvldA
qM0UMqBvQZd/qmOB/+KcxKnRLSFC/sXVVHd31L2UXN6Sfs9fi7hUtVlhNciCf9zH
p887/f9esPI5KS0kRuZ3aSHfHTGxE3zOnCDn1MuOMyeICyhD/FpalA3fnP5IbcEH
N3yUAAvNklPFabIyGBtLy6TkZ0KaC61XRjvj2EY7tGRTESrwLGhMomoC7uksoRWE
ahw7nk/ItVcE3NYNvL0VkT3wlfiuEbkBMOhhzdtEbBrJeyaBBVfjzaUCzFMp0qrW
30BhlSdfEw6dKfwLp23scQCYpuJD+M2TbpJptX2bm6ll8wrPqDo1eR7SlcgGJ+WO
752KHe6IOWUAlVsRmwOUQdelTFNw+nkeFpO+drq8pi/bjIFDG8epYX5vmS1B10r5
JuO2afNGAmqtWdq9f1z+/sYzpQgIu0asV1ODAOL9nswDYkhlxxN+f8WF9kavf43M
v+zb+6XQzz45cQO5dgSrOlJPm54zLtAIC8NcLD9I76BuY0V+KJ8uOiZEVW6GIm5H
5lyFKgKM0OObHYq7lVk8J/6DC9R7zSCiPk4mHaZIBwI0B5eCnUyV27PGiumJ0v+n
SZwtyK7O/6b1Bc/i2yhXZ9Iaxf8bmDWK1tsJcNmIV6nnRxKS35NkLHmZWXbh1L4x
I3QxXizLaqALv+cWYkrP8d8rsfcUlTvMpXEw6CJNQo4Y5SBu41TvQEAf8FgzlFi4
w1dX/uQH3I+0hkwfZDyuQvwHqXNM3AW7P4wo/VSiwTlD9PRxTAXVw73fSbVFEzZe
tlMuG4czViFoz2a7ahD4IxuYBz9Zw/Argkg1pdj648KP/gxHnq3KEJSAE8O3p7Oh
PWmAHuMtdq1nPzFk6Z8RHMHfHmPZhCprxrpe+aml7jIoXMp7Qi8uDEMuITE0fOGB
mOHD7ZCWwL+NVypV/3OEILA0PAOJNKKmDZOFsHGmOuIx5F7VTBh8c1NTKEoXx+YX
otEtlEJyMgfcVxq+IlM61/PwUyVu6JfdSWsNqUDb8xwg/IIwZFYQJR/1Bj8o3WiU
owvVrD7T4EJCULofaJgOw06OwjJOACdU44IquPM4GduyhCi26nxtq+1gSe79NJ1z
kLWjOwJuQKsQPt9mVB3b9dzzlS4AoP6tXYi2DRZbS3qEsjR0oeC2lz4vNCbnP23Q
9GHSU76LneuoKRXcu6ETuoyZ3scfterZcpS6xn+g91CXA+5iGsotFoVXrFpnyxCW
4k6sZGh4cqAPA8zes4vCAW8wT7I73En7BXrMrX8pJgnCkcdgvNhWWDy8JuRgRe4o
tly7qQK0u4J8zql//fuEpY6ppA0Af7b8jp0z5Z1y+aRP8QL5I8tiVrSVCifP5BIe
HajPDJ5gilEtKRr/6uypPBkdRxk7mYB9eCeAat3dMmk4XVFFxw0/eP+OQ0Qo9LIY
PJ7Tu9KvwgkTcBwmk4BnsIER7W/3Lff/+5Is4P0kdgV5qDIi8MD+IkbRR2kDMlgu
+QDmJw54rZAifzgURxefubMuNRE+dAsmM3G7Q7UnK7dOPJIB6i+Y6LDdWo17HKbQ
B/8dOXeta8S8QhOsVw36c30r5aqRb/e7zqEzruwzhv1na5vd2AROpWuf49MtHN7q
DoyjqNNXlMVF1gLXJCzW3yC1ARhjOwoGcJAbL1tDHgXNFxNiQrau+5ek6Q0hogPL
dWA90E4cUotyFMboWdLC0AHeAI3lGUwy8KZnF03y0fh7jhT9PIn18znplKMxcgdI
LA/jNWPIdppPO/kx3HeAbOs79dmnfc2JZ/SZtC9ejXfoxOF8I8serHB/wowtYqZ2
+k6USzLAuZ8GsBd2nyzhWIFKXV9rRXIn8xgSuI+szusFHXTlKOTuN0miMg5UAT8M
bkGKRb9CiUfEyOmleNkvir9/ThEAEwBUsejdiNGEnzyiBiTYq/ywvXlrG29rPc2h
NX2p8d5TXfXPouyhwvfhrYav1mEJS+1XqqrLWqOnK8Ur02VLskLwG7WKn+JJsU1v
1QHGca5xzlSHGXqY19IgR8q3dkW7PoFiMmV+yGI7JR4m+zzSk2jI0l5NZEzKVFkx
TV2/iP4mjYwfvZwqKUUkQQEABEs3dxuRdiHrL1s5r06nVPGNwHE168OKubRtbvbK
knfmCEfTfb5T1O2qF7PezwpnNaMacmd1Sov6nxW5gFDy0h6+8SVnAuX3NhDxOv0N
COjHofvQwmB8s3XEGL38lnd8SXcxW0mVKnP3xOV0NpkaqZQkiTweROo+ZzFuvyyQ
zcXkW5XeTB967uRMUQqGVgXXsSI7rb9HMxzOPQ1rm/RvhTu1XT4lTAS/uM4XWUGg
vLPNTL9bzHaTEgDcbdaDlkzRex9xoCFlfO/6HhtZSo9K8dNU1na4raZGfYi0W06O
UcPmPmMSX9KeFmmv4vpwhV/dL0NJe/Fb80TYUntFgNPUjBCMfa6k+vsU+rQFQxLj
DlECW8OTGafwP1L0/gekWa8gRbrr3yi4V8X5PKS5JcL0bAb+2bS7Y94Ndt3CX45L
P1oDvh3eaCToNoxri5cGbMVBhIgB+9k/4pPhbGFlsadzfxKFIVwj9oW0UsUxWRnT
7YZ4LE0DYGzSynODHJdW2Fi7ByakkaGkaj92boyCac5uMvSndWlXg6KhjPi7B5Oi
lxtnKfIY106UrqHdU5NX5Utq068IWltUswekZk1KU1Y9/9GDUCeAfTuVgy2VecOT
q/9vv1t6oPp0E+9HXTVYRi0v4+pn+5vMs4dB0KdHyV/U0bfTN4kQqoD2aRvRl3eu
OMr3BSubCqLQFZuORYsPazTDHJUqKpakbe7MPEQegmy2ywRXMggjHCeRkSVbWgay
EUAfr5KrP9uh6+ErfWbFBpPuz4jXnJembBn+XOxl/EKHnRtGNIRJPPKJEUHMmhYc
/taVT6HH9c/FxXg80swL1MhB7++0LfVz0qqSWj46N9dwh1EjAMEYwTwD95QIaI8C
2MtswNc3RQNi7UI8cQ3RmRar6y5NGyuJooz2qtABmH6JIC2wWY57ib7iSE3pxm7A
/fWLCoL9mrmQbdLRoVRx7Tq7eHw0K0yTotats96hKEefYZ63DDDdnPcYuH1Ngxkf
0fJRwxuAADVuhdXnKh2j39hZC5x5DS51d0D8+u5jj6E+w9CFOpmM5iMHNbz3Hfxx
wKCQ4LkOOntZCZaKpJ0LGz0eOsPYPmtVUNEtqZ0ZieFNR65+zL616bMc8fR0uQRb
boeXVx06B+wwzT7cN1I9PxdOdiOjYAhSJ/7hbAbpHSHujSkpkhkoZaweo1ycqEf0
6MYU7MNY+L8ysFHBMvKPPTz3SJKBzyeyguXrTjb1iULuePtnEW8ASTOg5cRukn10
s0PYgRphMW4eZm/0Q9MuFu0JRoM8YS7kr3jpwhLw8+GtB6HDo+QM2ybYrpWWkyIZ
x1XRB5l29XNXb542zIhoVEJhQKNbhvKZ/LQXyHNGx8mZ1jLhMN+1kxlK5xCv4Y3Q
2C1iqkqJnAQR1Dr7u1+dBvEuz193JWEs0+oU+dtMIckOuhnNon7wAk7q1M+BI2Vl
zO8JI/FJkMv88xDohrG4ngYlq75NKBZSF66SwJMvJ/Qt/pVKGwUBIBKjhc+yMAO9
HqCP3aEhsFfMbtV8FdrWmY8BgqoQIJX3c8YFhO/A+Dn+I4i4GDxm+aMa6RI3oyEB
wCi5KdDBPjSpMP+LU+9LbM2l62WkumNi6Qkzs5egGZ8NV0VrF+I274J9kxD1IYfO
xN7wHVpoWxxc3Bsc/HYKzTc8b0XcGlZb4AHhaSO3jT8nV0imjG16j+ffUuvzad7u
MOSUOHF802GB2ZOOw4BKSo44TyD/yjWAgmYrwOc/m2Aq1SubOtwq21js4r8N2Slb
HMUMIhMJOy+T3bZwUkZciCDag2BsXN94hriXtDMLwp8EBY65wSU+4wIc6uDAbE+U
9fGjesKJu5ZTZs4Q+vKPo5S5ZoBqfWvx6wS5v91SJ6YJit2oOZ/aMLKzzjnI6aiM
xw3GXrp+SI39Y6csaLdTfKzK9xjGuAlfy+QYXjDtF6XjewwoY1XkGnlYxdp/1IjH
KOgYRbf1zv0tCYBm55QBZDPWdkdquAthU0pIztJvxZfiW5xMAkXy66UMcNvDKeJO
kwjWoDh/eMqaTN2ciUygoiRGxYR1vVtUSpImJcYaB7SSNlqW6jSvsBWKCouf3uhH
TVpUiEb/iemAfueMMANhYmHnX36obJn1VPuYRVRyMpfW5Ae/WlwlJhaivI372pEM
v3U4akpz7Nd45cO6dt777zud9u1Q4qZn+s3H0n7er+wrWnBnT0e9fQbUKTUCHNeO
/kK3X68uizAl/88YlOM6Ln5pjgHK9nPTlLTFqF36PfkNbkI1qi9jxeT6qDASTeda
+n6UBcxhYVlGEefGxQZv1UH4XCXfllh0/saFjhIn+B+ele9ILhYN3bpo3TqGN9Kl
sF4y4FHaHRmiNGQfsqVtkGxs/YRyo9WDquMe3E7XM8LLO0r6pCTGHBACf+e9zSie
p1G2U/daUurewq253ubILyoW1kMi6oYDbAANIho8f/YXCPI49lS63oI0C28iBJDj
tEQr51da9zRjXKnZXBQyVX98yUc08J0fIZjtzJlXgjkg+IpSQQb9yc56FQK5O6M9
+ecV0mQ+lq87iCfKY/ztkmuZufM+DuAuA3WB/HWceFnnhkg9ss4Ge4zePmBACJt2
VCyT6U9K07rbl4ceQ/gIbEaV1RrngTYvsTa8hiJjxw1p/Pbf4UaPl2E5qZXVK5jW
BWc3l+DXhrg0hCQwyr5RmOM9sgNiZhg33TSwajZqX74RwS1aD1rCQmdBiNSgfrYz
USup8DhQ8///Pq32wRJbsmxZvXu3da8H95iKvMHma2h/rEJH/o38SwsDCSgMZgeS
3dSkydMuu8sBWkIThGH6G52/Ul5fdu64ViY/YF6/fkQiqQXu0nxZ9esZdZkH54oT
wI6AFVhTQ5guHAOWvNEQ5NQzfC7XL+2CQYmfvH6J/RMZ+YT1Bgq//kjN4O4f60kq
ZkFKmtY4MsLb9jtt3yAdvbGAbLBSI5SvLnoZjCzqqZ9TBJhQn7ygip12oI0RBpkE
5pWi538yT9c01Jj7/p1KB01zV7Vr1MuKEqIXK24dqCdLRD8xIKDv1CG8498e8hKk
pyeU2l1dVzUFCD2anraxSd8Tamav47ODARsnGinTHnwnjHvwkPJyNCF/aiZ+wj3X
kgW8JnAIhaQ364xltN5ivlPGlBL5ccLqDq37fDjhlZzn0O20noDpzNZAmTgALa/d
ZH5sIuFRMyvbkQWm6RC8kyn/5TamQxEcqz/tgiYXgftCDWNXUak6B+bi4OUL+e73
RidnHpbAe1Iqwc8r9P300cF+ClyfE3+3M9s37RKNmPP6AEC2Rp8CwzxJcVBpq7It
QViEMvbY3HqX/R6rrm2Ej6O1Y55XscI8lUO9Bo3yX2pJ1yMbjPS7aVrisCki7pbN
LnZbBSXQfCsz2MnETesWoAQ6sddLkHkUCTwRZOVmBYtBUHVh8emn1KeC59/Trqnd
HuK404crrHgoplMtXoJ828Jnw43x7/qrk8hr4ZTWmZBXVwErkrAJEjq0fippSZSF
aXjIu0Y9YyBH/haHFxhRznBhI+CuK4M7LEpJOAu3AaJaQXxDdzaTsTJ8vSzzdGr9
um/O7IqPqSB2N0K67338SURHb5pj1AxiusGOp6bf6mCZpngzJ1WciAXolIaAhASP
lqoHtZGGGlXS8j3efd64GRaceKiirdw7NWezsR0I6zcqKSRo7pO21O5u1yumN1Ce
WBmHgJNIptBF4xKB/Jz0sC2f3sOptT2EXibw4ILhh2fyR8m4S8z2OVBYiCWUZlgh
gpZMDNLsLaxiwC1xpVfh2XKDJfQjIsAjx0T1bzzlUw5awl74Uy+8f5Hjbv09VVaS
aZreoOI43ub9FcX5sT8ZXI1cVoik8pwpz0oLDQ754DqvQQNdFsg0m71kIzMPHz6j
jYZbQZPmGOVUgtYX1fJxLb8z2iHj6IP+rfbjacDgjMQfzxTxWOGJ8O4f/gICZbYf
GQ9rJdGKMiIbu6ogomiwdvgiDQSTuL/318Rj6KfEcpVVBGcmZMNbQVowUkh6ozXn
nnX7YrD5iRpOPLfJQ1oUdn6nSExVScAaoL6kco+KoubkO86CMQ+3JJKStgupu4mF
D7+EDNYs1J8ROxfnIG1O52bAikHLN3nSPOqTnlyVgXc+CVp5KrmxCo8Pd+xAWQkr
g4YBB6RzvVnaUOLJrPcNjk1KEANtEZV7TMZt46PyXhs3QI6nw5t+r+JD5aRjuIA2
8bSVIczQaP9QlSRyPuTG8S/iPKMok6/at/am2LK0u5R/Xqwo+GCYFeakua3ucNB/
97VoGczWZ2djvFI+iO/uuM33p8YihZ4n5sqqbHuQDNfR56N7LbaqmNFYqAUr6xKW
HOOWDxsgvpkox2cR+w/R24Iqynk7m75eCi9HdekljNMYn/4gf/kS26sOLrBZXPb8
VethI2P0yMuhurcpCbdl3cb9Q9Conukl8985LNXF6lk4OyUzBDehS1jtrpYavVZ+
SZCJstjNXkpTviN1xwd/5kBbTHQEVnVWnMRcLxsA8LydCp47o3yjjKNrmxrqcqNO
/+XtBnrFooPeuj3c2TJ4jLSQCKTY5lWwSAjAwVbkEL5Q3yNI+zT6owsDx/g3CdmK
XEJFdssStugggP1L87+mzygcfIy4lZL3O7cscClSIB7ICdgWVxfw0YkLl1qdam8S
j47rADgSyLiHfgVifPm8On4lqkvwhf3l9sRxWJ7mzlX286V5wXiEzFR8BxsuNigO
O9juC4chudQWmIdsrRC9GJTwB2E865JenC7qEBMn+xWx1NyCYIMP4nOcbDhbhbuK
GsTnqZLbcNvgJP/A0YqtlRNk68r/5otpejX4NzKhA4So2RatROCGdwFmpLMJUM3B
sk4H1nZteC7Ma0n9kYkt6YnNBuKBvSVmeWfFRrPlRK/XovAGTRRbBlYnPManyRqv
bF6u3dfo8Kq58XBVySzWP5p+S1kGQ/YQ65BsJOh9pFWb8dqSv0Yqye+YxDXfvugf
QQwh8v/ek5MK4H1a5xIi4m0ZV/7wh+lxKqeFI/cyHrjG7d0XKgZiztDpWcgbgWEE
EDJ8sMzm5m9PrR8KIzGL6qZZOMAciwHs+nXBZDVaOzoUtRju/WQRDOm/DUfjh1xI
79sbIMhzu+ZxuzpgvRfu/eBfhrUAhEuTZ0PbBC1U+xhjEPVKOKJi6ux5u54MIBJI
CR7JvG6laFu40VwAdXtg3eAlCfzXT0NRGGVAWH/6cZSAdJtIZ381aBu4hInQi++i
43q7m4fJazrG0XIgaRQ8sqsH+SWmMGCsnZM0xaGTMrcG9MfQ1zYKFZSD91OjLfqb
XyzUGzwTgl5LcDMaINKV07IxTZp1o4CZAHfYxeETzb1bAEEUETBFyJApDJWfQs5N
7/socSs5w51b3rG7c0rhaw4LuwofV4HDIe6/WSpWF+NfaWI4xpD03O2GvWhm38Lo
jrZ4j+uM/YFc7te46TVJ8FRoS6p2wbiENpuBq0+IRaLScOQWcmA/kK51EbBrvcle
Aj4S01bVX3B+nKeOLa4wpQxe30Ye2BU74EpG74dfB7iSWT9CMjR2Eo/e9WLXew/I
TTZD3lZ95s+bswR2yY1KvPMqqjODd+9YY4Ko0gq9TceC+jYKGViKkCgOHkmXlvNx
Uj+sQU9RavPO1F0GygqQjaQh8z2kFIm260i9/y/qHnorvboMY9q8cHzvqTRW1H1U
RAW7QmCEITNB6lxDTikktLA6fZO1rHLbDzn2TS19uaI3llTrhErBmWbqMfHdZe4d
I/wNfNBtoxNByXEtfQuiqkE6iOUs3x1O5QlY05J1f07jW+PLpqRbCuf+Jr1xqMdt
4mqR9gny2VzuMyisL6GZ+HtNGw7zQ1U0hig5AQOyuaq9Otm5bLGXCxgldTzXPCMV
tZEerf6CoMIEVi1WFHBbdfIGAU20bymaq6I2YCryPSSmbpifsL4BvGgOz9v0XhSi
RtYNrKqEGtkHDqhXqhcTZE04lTt1wdotVc19fJemgiEWaOvfT78AgdyCkyqBkqp9
vIVkBQCwLN1/tLW+47XHRpFz3Qu1zdu5AdEaEAJ1ss2epAIEHaZR0Q05I0ORrl0p
Bo6NKxBbe2+5OeZ/I1OMELk/9p2pE5KMNLb8nghkGxieLzySTbjmIX5wE/0kFRHj
4manlqXLSBuRdyTtX3ns45iwKkbLmGpU83uCJ1MPpXiX3WpoH6BKJI7dYkPSL8IS
T1t3SZQVqc3jM0VcmQEOjsRV/6TqFTaF4yFa+29D6Bxc5lpLYt8AX4j20Nt+TGsW
oqSuDDgfouyXgECG6E0YeP5pW2c5aHQPcmc3+cvJ9meZ73vidFQED3GeeTGwTkEA
XxQz3lauxKm1KyjQDsUafFAMnuAK6s/WYoH9pex56QGs8UXZNR/xSX3o5ka+9bhC
0OnOHmI5o6/UHZLNokRRPK2Es5VAzP6QfodBIYChqfPlW9Z7BxI3Aeu/ZIpyseFe
KeXaUDJlU2pA/FAa+j1702n7M0LrbOB/kkgvYR/OzRhpcg6dkL+LUl4EgJYmyQr4
oWyTPflDXZrwkP7PLpn4N2G5LVngDEnOimOmQQGSz5gcYHXD2NfKX+W2Y2RWg9RG
HzNi9oFp0DoHUuG8l1LGxIgsLWDtaRD5vQSopx17KTL3soWxp1+0iGFqShYREKkC
Rx1jynl8Zm9JPFj9unHxZus+x74uvj7QrWBYNS9upb3DPDenblGlF6WP6HSgCI8L
Bq+Um05zQ4aQblF46Np6qDPDfrHznMWtgE+FwwTTU9WVIDjOOZ8YZrtQi2jXHU4m
m3LAMYx5LUjXMucKbBsahMkcvnaFL0dgDWgZCkQz4+6tZ3iGJpmVTfmIBPfReECV
0mLKZICx9P+SyK3EBTFs8DVoggz39QJZS7Z8HdaEQOmVYl2vTSCMoeqogoneLtjv
iGNhZQvUaB5e3NSMzv88egZNI+KR9EbHWlTrlZ+8pUyEOghnQyefYicSU7szzboc
ho6DHQTjJLSrtI/B9NJHaewoXvLyLd6auARitJdEqfvKqxJSzicI8pLqp5ot+C8D
jarNz+7l9A7X83NRhdnIJsR//ZWkfH2SnorvmJurq8leR8nHgNIysTqeuHqvNZWB
yVgGhZkoXARuw7lmbgHdKy0489OLYEnAkIgsGuiqzZrS7SutNROwqkVqJ54BLaxA
tn6IE4n71JAxCl6o7AuoegfEP4LsiV7iHB8dsOLRH5isgamIsja7rmBdf3OPwMLZ
xaV9lsNDBKkt9PCwX5GDMx3qw04hdI+ltCBN0tswOYzJ9xMBwrx26FGAQtg7Yzp9
oAqW5y0inmdtKWTHGxqmjN0CvY5Hhc7qkC161/Q5tT9pUENOjSwXfpT2a8qigZp2
xewfpc7faQlYPDC5YFROS3Mgn2Bawxy86F6hoiM2gQy7RxYM56uPoRoJmZ86LCDt
e53TRonMUCPTbAReb/UE73X2GloodK6Dum20p2JCgqW+jIO8PVp6A56XPZQMQoYM
T0Ye5kjr2oEXVEwnDueVHHuSXFNl3qow09Y10g+xQg090r4eFzcY4Iz6VYiMF+6E
qaBMRvJv09rLHfv1e51K94EExC9Ka8Galpg9LJ0kyCi7KWs5q2wfX6o0Z4Q7Ci+d
O1SvojmLZ5qwXwi5/c+tPyZYg2B92Yc5pa9/VOISxKlEPfNJELihAUUtHYwrtdwE
SvX9Vv+gD3WfJ1ADpVrHSqmLJybQxS6LpF698p/JCA8GolHYWv23R6u+j36x0B78
v4/tFQFxkeaib8r/v/GDDJxfHEKXeNu8jrrozVZz5Q9qO+MgfASJR6iRQv5j9/KT
EAF3vBrMFATVVDSTmAyFcmO/1nFxylSQHoyCRbvl7u3Zsa9mr+TG6ZNuNo+cja0q
VJithVIQvx2Jrihk3XamGdKfxUZq/jyCz3szhRWArlPAKlGrFtrgdqArOaHstYZf
q4acnRQqyl53f5TvKE5LYU4F01J0VZnQZYtKE0iSF7iF4c4QMgz/6MkidOsRY2d+
iz8ohEktTusf8CKSWPz78F/lPoXqa/nzuB0Gg2PeJfqGD5xP2MNiR5m48ZYccUwA
W3xtb00wM4tXQPBKHAq6ElV7MyZ8oApNmG8L4oVWuTfWA/RhjInTWaVNsNA/gNoB
HEAGXIqf8ptanLFHmJP9kgGUxzbRS6eWyZ6291UN72JmakdXWMCn0cMift+BUC9I
ocqH9ErzDH+6KFPU1CkMmwPHwlk3l7B54a0v7RdmPWcZU8zxw+18IfZ+Q/xvhIxv
ddNOtD2yxdynSEyW1ZDkEBazPjgAiqQL3k/cVCu3mhqJGYGwQnamgLDJ7V8Rt/M9
a7WiQKuAI5A2pejjs6D7AXokYz2t51R8weP0qnGYZcW4ECA8l3XICXNDB6Jfv9VO
sVXvpaGGT+7/8PALRqx6yHqoyBJKCBDf6eS3W6e6Czm9YBGbEj8sSEb/tFv+qCzE
3b4IDDCMk5cQUXQGSMGNYv1Q3wdFiSmXRD2bPsAOt+F9lIisQcsxkZTG1pno2k3D
MToyM+3FpiKNeW7Gf4C2FhQrR8B5xyBGWBmjew3kOo+yolXawqQ8mfVBb5X3St9u
Xn8ZYJjxOcB2XqOz3pnhG9Ueesq+CbJe6ZCy/B3RwMDtIgvfj2VtWpllycSV5dr8
2EIIYYT0GkPvh2hMdaUXGjk8DP773koZ+MT7uEAEoP76Zyatjr9Hb2KE1GxQu/kQ
OktDuiMAUwGN1PLaL5O6fJ8RkYdqwZBZiVmsk3tRQwVfEmh/MtsvLgookOVpfDpk
m+SbCcEU6605Q2K2kp0ssvsX5Z+vNyGYbtFwpGE0yPsSRWGhcn1AR8eyN6nKBqFh
hzhEZ3v5Of0om4P4DEeqA5mAWfvilFs+7hg9VA2LBHfo8uXd497T9FOV9fygMjiE
loRh2hwK5Cts63enkh1kaZKmzTajX0nqThr5pE6Pfw/1RmSU6diBMAZhBnVr587E
03LZDZX/0F3rlX3lE6kjk9XHflhb2etT2v0Fgq0DqlnDaC+zdtR9Hqk9Ia6nIK0O
3GXTg1ugky08xUk055Oy4VSstcpCW1LnIZioItvpCbYaItHr9W4aUkwFAeWd8rwt
htpdsbGaRf+I366fyJnGtmUhzVo7m455zIwQoaQUx+Yol/wHih15lndyuZ/R8bsi
xeVPGFGGo8L4TFPaFcjExJDXaSw10nEmV8bUdNak3+3IUOBsS2bHDYwmnFVOptSW
tnN2IxlLXT/95jWKy/efZKMkAgmVmnz+/RmiM6U+hwnficjJPJMUNg+cETmDS4ws
jqyDPTIcgvGpmnS5TsfQjQsxqoKsqb7GSRSFkikhpLRPthuyeABgp9qW+GmIFDiK
4JmNjVpAskyCJMhbHf/Q6NfhRJSKskqdn2AZUZ75QroOzr+GBKbbkhprRIUDue4V
ySa6S3eb4fOWsOaF0Zskdq+UpyzqOI8dr93eghNGh8BQCU7+NjFxMGCbmA6ZyguP
96qCEOXtRps+T2CO9iJD45JZGyQuQSj4PAM9i5OIfnOYNjB5RivhROpdsSg0pgBC
G5gPgKm0vi+758NZ3yndfKuVD+P5nUiooIuvrmvEcn8YZPWZyIHVV01qprcMDDY/
pUJ9Z7WZBeqfFTqeXfE0hEtHPfuYTS8Nu/8DPdlSMWyS1HgEOB75iz888iTtxEw7
qhlSXzPzPxIwAZRs3epM/YUVbSXgoH8udBCppJ+KXtz4mY8Dwvhuey9MX8Y6gf/K
2AxDSbgf2dEyYBnMYGy3njbIiTtNBjafiZS3J/SjedyeWTrW/pZ5WpgEhIwEgKig
Sy1EatP8Nge+8en4ygKT++d8/J5iYtDDaD7/fVOZgztXT+B/N4ppcx9bvBi9bp8Y
shIUe/frIUBlA8a4With6kM3QleptW4Dd9DKX3RjlrzFLTnlSAHLtmbkGxI0ilmf
/gZo9X+VoWr68nkL6zWYXeX84QI5dzsBqyZtOAgpj2HadVE75neKN8HZ8LsR4WSx
iT6lZFGd7oP0NVwnQB+ro/1ORhUCZ11FYd7hHzc2r8JmELQS4agV3yFyctJ6/+tu
q2D0L8l8H0D5kvWxuaY7/9tisZovvXX7NOnBhcV2xAowdDINnymD4G/D4apcV8G0
s84KY1LdI2hTfvsZz/wAXx+2bKIkjlWoWcYqzr8GOHbIa1piCzQd5jKVzvpDA5ZO
CnnyVWviTS3zWWfpRVHIca2gEU6rV1mpq6QC/rrmAU9peOLeZ4+VGIqFQlgyxJLv
d21UJdowFy5y7uY76QCn3UkNoyJ5Ne023/5zxpRtP15HGpN9Y3YiQsONJWa0PflU
VN0ykd9Dak+Cq2kkgCyW5jaBPihz2V+aIDcmf0q1QqAVqWM81YAyP+XlC+Ls/9nn
NPFHGFq/0YlpXrIF2z0uHardQ+Guqs7M2DNiMGiiuCmrxp8r7P7goyOJiUMdWGmR
7vu+EM2L5e1jrTtZFZIlqPaFTo2OrgIiHrU4Q3cB6dpSbzWwFCH8AxkPsNCk4/ZD
5KMeP5l4RCV9pGAExyJ3gcGlkjo+7rkj/DEj3xuDaF+wXhKJBMpiFU4jVaR5Phmr
HRhAhItTNWD9FB5rSzRBoezPIQQTsO9fwpCFkJGRzaBGDjMHSJvlPcPkYBPoxpHc
7BsLIsqAIvpN7zixdtVRdD+yY1H3c5ivb7bgzwAmhKkWN+YLbspmO+qCGDNn9t8O
XAA3C4FgkKrvqhsVjEpwFOsAgInHgVfSMvKfTKHQ9I4l9HTJHSupDd9pnxKYrcgl
p/GS3FKDcjRjM+KS9Ms2k/aUf03nUQ4oaWQjMlGXvWdbwNYk1h87JNYBbm4zkoi9
Y80Sv2qiPpIjimVyQe4KAlGwW8/CWgXFXIJ2LecGjKUkCdq51dV3rwbRKHFy0w1+
A55cFHrlik4GEq4xa6FHsVHaN0vF0215zMOH7d+DFws/7GHkR8hv6sC6R+h15MK8
+HzrVTAoSYpc6bEl3N31fDy6Ta1xvmQbFlt/fGCCPw+9e+cfazMDHJ2/UcG2JJp7
Pe8VmeMu6+o731O+zCHWsa8oxnyg2CQC37IFRvKiJvFFGkjD/1AZGrUosVVzPWOA
f4IZHGdwb27Y4YKigSSpirzFnK39Y1tXRCoDgF+8U1rfCGrlKuSvL4pGDoFHrpk9
nkAkzL4YDA7lVeYx9Lj2iOxzZjOw0rNdl1wrXwc9Z+ULfEqU29m0JtaQQB3nVa0E
UKBIyFZlRiKN6Dv8SxfXFkpCQLmBFC2KP9ns4/3/6Wmac3lrOKFJzj9yxJnwUiCU
60wspKhCXkca1ukkFsu/AdATNgzfjP/PWLv0CvXITd1FRQDzsrDKTPvvHj55ISJ+
v0NQfg7KS0r+38SjPpNK+RQ/7FRDekWv8yf7sf+9pWXcC4u25dapb+c6pQE3fV9j
OdZ+VAfigaH/sdPlUUgwh/8xGRvr3QltJVM9kJ7g4JJZsVfnf//cNTQE59ADNBnt
oeBGHDCEwK2NapItNh9Yjf/iFOJl6jiSWE9wLDu6dzV4acTTzqeUkeksTbEWbwzc
6fhm2eaGsx0/OXwk6WTroUXEAIYhSwdYCbaldpUmsdnziep4FcleR9eWmZG5rQmi
3fODWcuOMAiJyzRCr1yP5m5yl96dkjno9sZemn1TK0GinB7sFDg55hDlAoYGs/gp
UVdxnWpf1V9xQP1eYUmZFRKznvxX6tWLYph9ls35Yn3hOzmqqXjNh0sRv84A9RfW
AW99OBuGY93NGuAyDxGYQGopCcUtUuIxGL8OH4TCrxIHYAxZJ/PFAouWsxqaGVzr
PKTemLiWHv0Y4lBFpb5kfprAwJiIWXEE9xOXwEd+bxKXKCbzcLVbfga/O6qsG1Yi
3jX6vL5n+D9TLzNrCTH04H9CN77UQJ5EmQpK7FaWUu8oIdDzJVDA9shEy+OcUCKU
dmOExbExkw4yUT9jarmFc7oIHaZpJtgvcMl4KfOuyvLC3GJHxNNeQAKAa+igx3zA
6wTzkReF4U8b/XXLau3QXHMZ2gLK2/t6ALaqI9utsmoXYG8jS5VRgNIShXI+gJDj
BTOTWwX7UWe65ae0RRu+I4rNIlArY5xFn7S8ECh6Dw6m/SZNbjKYyvzbChUh0SXS
kdLwHOroYgKrcGVJUqYAWusryC7b4znUwaulsyERJ5+ZI5o0e/dO2t9pbwOvY2kl
Ko5DGoschCvOVyyU755BFWC0Z2zXU2CL2gcri8PUc5ISe+jdI9JD9LN4HgLn3M8m
LEsOzQ3m2H19r8mznFdwNYdYZ/yLUBFSXqyYjG33ijrMa6ni2xld0nE007CnmqzU
PnyLHADvfWzB1KkPGry8tMYMUPzGOwP5rF9BVA9N84v8dLjE3zdeq/efA1Jvg8wm
XgyxLWYxfwk5rcD7sU4TB/f8tuv0c1jNGqfvXjnfN2MKc/Zojotn8KH8DTy7rMon
IbWqRA6SeJdallMwI1c1CEtf9QhdJrrkoYrFyu5QBe2pGv1dURyX+6vNPLxNo5rh
K0lq1O+w80quK5Cpe59yb5b9QL09X7wP4qfJL/OpfN/k0BcE+uuFs8/FBwwBbz+l
xvz/lxkILHZftbFGBDF7u26ZXt+G86SEz94mXQ6pP6m4w0seZ5BWoWlFaQxDM7vA
eyISdZeI+ua7X9FTwpBrOboleVaLea87qNsj5C+UCJiLP+7bev826HogUqmJXTvF
HLVdX6A2J9y7ZZR0FyLcwSFpqsXxB+k3htWPkhNzslF6RAMYiLa7DNxBt80/nYxB
nrRljE+75W64Z/KfPxu7x5QkPMSa32s9UFYAxHnfmKl2Xrz6sK6RaIlyEptrv7cq
3Se4/4xjvNv7WzHeF9vmj5M1nOzRd/rgR4buCO79DWW+W7rHCejpOVBtBDemq/e+
dVw1r1nA0qaggBBYimH1TyXkH7Lm2mAjfPiWPqkfeOXAphIzA/s0SbuBYUc8Q9Hl
SArpQRDjMJahs53uxhqSqboG3LuaJCcuwAr+Btwv2wwFiV0aNd9lHdeh1GGV5hR/
w7rO/xV+9G8advYtM+WSRDNsnrTIM7xHv6IVP9uiyWAyR+jT+Oa/HX+lIyzJsNu2
ireHw5+8HK1O+XLq8iQ7stBNjkTMseoMb4DzngkXQmJE1gVKt9L6cC0abdwCJ5or
g92nBB9KtKPDGyX3SSmY+H+tLauUnZXKmim2Jak01aFrkjii046gz5IdbEY1ZUeq
MnjqdXlGDflGV1xd1Rv49b+tvG5w11O64rwg9nGXJdJ3JRSkdnw9EejzqNCDYf/J
7A8uljTEHLaJiYsFegbM6WzY4fktMntJVRW3P44ngdGsVS+D93K1o8fZVZNDzx7p
SVLvfvXpv5RzaxdvMzqSk5D1RGEZKw4bSwtfKcVQs45f/DxhmFG4hZVl1fl7obGE
fKL+H1hZDKsuHBU2oRi9mVki864Jff0/D9p4tgZhKaQbrWp7K3X0Dx+FSOUS7tfR
8PelvUYJpXV8Bu9n7EdyH/pbx+Rw5BOLvdgeN3CLViQYti4FnWuz3o639qsm8E69
hK2631dxE6WgNONlCBlv0sQ2MJbrKQeLUHBnCudUZT2uBJMfCzQP/URUjwYfP5iV
3NQ5YggwMyYwqGVLFpYd7slVd4Y1Qj8Jq8h8YlzYIWdENR8LNJy5k1kMYGTHHmEE
l3SyOZa8Ig+1r7BbOLjLU+Jd12yoP8zgTIMb6PwCbpA+7DRF3w+Xo8BuMHXTBBxs
HLB86V4mZ8ZB2akBD5xKy58u/QrDD2z6c04VwID/uyvMlWnttfNpKyO/ujwg06+F
px+5aDWvLPyq6dkXmBWG8faRJN3IzJHbEePoZ+2ngCM84QqKMac90DtLI8La3hld
b71+3Msn9HIu1zTLrckqhzyOsKM/vXT6lkzCEs/upWxKNIcjLFOTRvxzUuWi78zU
PPOk8EUj7N+Rb9yE2sKXuNf9Q8htSZWDZIMhAxXNHLFVaFh4Wi+jeQrzDch8Ti6A
9s1rqdRuw1ItSTQmQmPMrquSsPU55Iv8BQabdo1Kl23eLaIXOkFzLa/ze5TGrLPk
8V04wjnMsmdMhUdvR6VSZ4ysgy1YwD/NNMSSmdh1Ie5pEG6YREHhztEXy0qY5Hfi
GfQF8dNYB8nZ2okNCavLup0Uix98yYJnrxfaf6H/4xadmclyPyKoPixn4gVf7Pzv
zAvJjLCayrre6HcAf2AsbASPYKeb2lBf8iatbYvQk2oUFGjF3FFmkfTyACjALfie
jKFXEO2ga/2+kxquB9Wbw/D7G6Eanhv5rnuBevdpzFsz9Wy+T+PkMwpHkmQ/4KYv
DV2kYvvyUxnULp/rsB3FgORcT+7uHVzLJY7ZuuEecfFiIVMvJQUwHNLQZuOQ3+Nb
8C0UnvZlQIySX1jo3nD1aQVnoZz0F7dE2cEg+gsyZrazxqFDSYX6XQLsvK2oMbXR
C1nTsTulIoQC3MBEmySsdH6dZlbR+eiBv0xfDPabZcjiUE+WgdGVBRHMpcR0Tj09
4FkOuS1WfMb8q8AdyNg/i06KI52xiwsttp1u3YXABwv3WMNdg6sI6Y4Y47UFD/Io
v20zv25EfCDWvXXqr3KIyy8ptzbrYfsxGURzBU66Gu0cH002fCaNV/cRas5WJEYF
f6mEENpwLYhiyDsqtxsqMZRilspvS7I/D4Q0tjb+Pn4v3YPz496swPg2wuqBJfUr
s5wKIz61UJNm3vJdg0piNxcHFUeCU6Wxe1MMVIxIDF3ZyQ99gpIeMXH8yK7eytfW
T+7rooI6KBdharzbLLzOhmgEtthj1Z2lrwsRcsjb6VFjEiczrIIgJ2jPZiGzmN4m
z1EoOQsEPQ8xWbXv1o7OaHYq9jEiu2aqvjl9Fe5MmRHaQWr05/UzvYs7D8iG60nD
vrQMj3LHxJcNm9EUli1rqHthgjP/y9tB4z9lMX7/s25Tws6McIJjnpK9WlmAPMj4
pwfXbIHV0hJjD2Je9qwk6kcdVqgmAtnYj3KFflk+HO2934f5ui73OfRxwwq2qtIU
JsCjA2IohC7Ra7ytK2sX9NPRnQUjAPJTF7gxAqxt3IOKOXLqnuaZsL1XFnRTqE7g
LWC9Z5xx7UlL6kv4OKILftw6b+35vFOxfXnmFBvak8kDLTeGRE8gsWbNwOqOv+8n
GpL1OhuMV01DdmOBsGdsmIsVKbWDbP6BiLMTeKu877mmhCq4SpVwYkSScIqRp7Fx
s3FX0T/kSMEldJ/8oeg0PYjv17pu7nKr0zhkgFY7QdVQvoAFyRrDNzkVoQ+2wZT3
5HN69lCKWh4eTUhNiY8sEmVOgA3TGw2OIEa41x4714hsxop7/Ej+SlKmQHsfKoa2
0PUbHzdvmVgey/8WKVXa/PlFuOeAEUwLKdTC/a1P/mSCU1km2mIAI/6GHrVED++W
gvfR1xm7bzf3aqUry0qLTZRpMq1ukipq002OXd3pfg/fHDRf2y7mgaAoWR5kvV8Z
dECB2r+Yj9LGSrtJyhZ+HEDwgX7AAVgHLGAbnR1frpfMqXP8ggVkeV+VlEmS2/mc
rwRuJ+53wm6p7rfqQ/mPk0mNOn0Q2pb2bV8k3iKehhkvdighiqy7qDUDxH2QQjIg
mTGtowfSHMxuqxR2MjACKo6nXXVfP4wgxElGqHSOYAdx+8OpWZikqNnUPnnO295D
EUTFlJeIbvjxLPBP33QBSI1jN0WQ7simbrh0IjeKZbooEZecGbxj/4nUtUN4sQgu
NUaFWLLbaXrwZcuQbC6UmkjVQ11dQkHimW2l1SF98qef7fDNw3iLzK6YLwUmeTCD
k3dKx+due/7PTtGG4c3mTwFzNiQvPNxu/TslxBUEstBBGhnGtn9s6sA6FiombhQf
hPiHjgNIFMWcQk4+SbmcDepom2C8LhJVYUuqj4a8h5Z+68dNzjA7B/QWWQJW8C9z
Jce1xKz3g3bDJIy5tJALdzCnXrP/EfbfxdDahYjSCfKeUvnrZSHFXeio2Nf4okwR
UVdlCGLfwdbP8Y0iwKKUhfn23iSJHdDaKWJYuqkyq8m/Y/GUq9dgg7qOTT1Es+px
IsvrBxGH/ydtwav8z+bPrgHvi7SL99Uf/FAkoN0TOnXL/zW0mHlAP+9Ygs2e1wOP
zlEIjx8hOoMTBukvLXo7lllBmyJPPDBiri6ng3IGamP8CZKp2ZpAE3f3iC+fc11/
R/xPVOopFxTE6RnFHp9QVJZkt+tUMdxgL6H3AFp5hWtKqFjNy/TgDjrKmXWaeRSz
em8OZ7AzP7QyAvYIFEV5jQfbdCTTifFpZYCp/Pi5r8wrNmFdkpxLZH7VdFfR5ZLr
HISJ/HoG9+VM5En8uLovlSdwJHJnOCH56u3dkJyuXci++o+AzOaXFCvzwherjvxa
C/OZc60sKR3paDrdGE8L6Z40mq/8FwssJntHiTfrK7Mh+pF9e5sAOS4dwDYkUIrj
0UHfp++IgnkDJajENtWaOY1IJSGP+DMMG8YS7NTKOUQQr4BwoZ+y5hjACzZ/U/No
vkT6IgwfYeX6Xa2kvvNSyXOsNIvqtfCsER/fEp4b8vRUV0VKN1WPVOpXtz9EE3vG
Y2Zcjj6guG/8v4L+VlvRVvsmlLxX6/TPtY66hETb1K60F+8V41vmQOEc9tBKHMK2
KIYwJJxHXgm727+4ifih4uyQZZr00vQws17nskiKRRWFEdaxBsIGCzHB5umyDC/X
isOxywUibDxbThK+qx7DDhbGbno3vHzDs7PvsybQyw+cwcT0Eqp7i0FqyLt+bcXt
LkC+JtK3WUJsWkndSZKn681qlk6DyFGu7ozMwXXrD4v2pF+pdqcQDVU/cLweSywX
Aa9RQYaVM/oXqc3Eio5CS7BC0rOsfOXWO8A2RwHwcvskvzw7/e40d1qz8Q7vDQY0
Gwi51aTlSAtJz/bE5TJfY+WFNDCFqXQQLRgXJfeboHDmr3xYiqNKaEfwxst5gUbC
cq3OMT6hV25qTRmc0CWglnIDi5DKhQuJsIINEqbb+O66XNIRzcCdYbdET6TD+RN9
nNKTr5j9FQTTaBnM+HTA9I09cpMmLOU+1YpmQ+25gEFSvM3iHh1VnKyfSndPd50q
ONINn9iP7JDI1ROH/+mNypbzGbuPgF/GpSaTqfsl/m95fufi7UY5Ps0WKepDKBUz
oAtwNua48YRR2z80MSom0PkN3y5QYYSI7VrRF9rcmNDkILT0nCgKsfoKczG+mtM3
BM5oAnUORij9mMQurjDyUHbcgX3r7xHIkaK6OG7er3ksljG38ERxzLxLd6ny35JN
s/NQzOlf9qE9sskBKzfncHVFTEpajKOmUmXqlG+J5TrbH2AxikgPlKty2OF59GpT
mY9Zkfq0erweu3jnIh+qVv5AYK6kz2qlKiGvzO8XfRj5uuf6eE/Re0BAqQZck9et
FcR6fnfs1Y6r/0dArq+fcYpJNx7d60L65+tmaRSixXR/45GYPqApCW1wTLteJW48
9rpLFKWcUq9mVai//B+yRIwWN+U4ACFS8LOZtrmvJtA9S7b5qkPJhdOPim9Z+6nP
AfM+CL4rvzmcMCpMyH6J1Q69WzYo7Uht/oB7SWt0XB0tz4aRTwc6Q/GL5hEVM/76
YqVn0g3y1CWY3RkBlr6APvK9Ujv/Bq7q2Nyl3uPihZSRqgEkUVf+f6T+u6TChsJE
Ldt+ck4y2it0UzZ6FUZKP14o34g+3vRZbGe1X7rEpunz7LklF+k6gxOJNNVu8EBT
buiLROasivN6IaDC+2ZGDs87krosVTIrh1G6QAnKPpXkwGorriBukM2BZnuncn1x
97L+EmFx+9B7tOuRK9S9VOTs25JMakaXNXIXNg3ygoKZak9cVeb9u2aSvnLrWy7C
i9Coov9Yi+IV9LRxzUG8lqbpUZcAZv7TbcO/Vkv7Ae+OCEYmfIKLEK9ax/D6P5MX
1Nj1ElgUxSRJ3RQUqK1VWIO2+2QvlgmlYKCAoZDvhcxf27LolyIVkAzG0oM0O0IO
przZHD5oKDSknbrC0P40z4YPW/WfW22V7/zLElCnSsLNsxiZ90c5OVL3zb9tYlQ8
Yehlo8s8R9eKK1yHGyZNzCwt0Q+L3wVU7RYgTBTfjt/D26KPc+Aj5HEiL3F/Bq2a
DqU9TuXHunM1dCclBR/+01wsXlOd+FEVq4tjYlh1xxGXTYvVfEYWU+BAUzeQhXxD
GAXWdYrax8IvsLe92gB8ctoBaZTRZJ+7fvLjD+uX0OGWfyZ3zAF98In5MDdTG2J0
sLOjlY592qHogqC6DfYxj0par8ryG001NSXDI2CbkV4IApihddn0YmIG+LIHj1Se
HPJmJ77W9qQnywvFMGQ+VMVXNHQXFFjy6v37sRyTn2Ri71dlckuodrP0EZOEEynY
n3p8OrZtsYHP3BHEdYDyRdzvwsO2gbyVqmu7Z9dqDkzW5DLtkVrCKCpd4XuaITSR
QTg16rUnpDJihU9LyzsnyPHmolBJDsIfsIPKlk1/Li6cwCqF9zm8EZ0KM7Mmrilw
j7rQaXKpSvYSltpU39FFGzVHdE0r6WLEUH8nSDMkG8TcjSvLQpGJ3QA6Z9Y70TK6
DtWyeAtNA37Bg6JIjHlEh4u9+LPnToNJM2d8lwlJIJA85gn9HoojUDQJAQMH+Qvg
eZVnaeheo4h8GcJgLnO8y0js90pHHVnvQhKq5O2Dq+ZVRM2hZXeIrvzSD9mLJ1/O
m1LAE71Pkf+MtGaNeoNCfKHdOEPRyyT8NyBVGMIRb7V8RO1YIzwgzbF6sEolshi6
fBriDvHIZZ61jD/TlouVBX+Eff2DYM83tjJCKHDW05kB20AO0knDm/Lr3QeszZEc
G1xFax7E1ivyYaFC0+dfNwhwISS9ZA1+KrU7rQRF16GmtI8oVl1EFnSiLPwgwl5x
jznrOU1lfSXZfeaM61MERPzalaEXKPtquc6R2u9H5uqdVLvxMz3s6Lkyr6eW9KdH
tTKA4GqxTVcVcQbCiQbG4C0NTFVmSnMRZwnNCNf1WKJTCFYlZtQr2+uF2oACdQn/
ssocaMbvJG884GXMN6/500xeiDr+CsjxbxWUkzxGSvtfjNNHK7AwcHNcW2/33qFI
EHVyKbjP68zNQBBGwvZgk37tiMokt+/bJlSe/qsCezk2ypUo7AkUSmRuxvmWR4ou
m3si71gfqj6sFEGyxyD+kRVm1GqyGAYrpKv3H4re5wNva4mhIFx0/aOzcyUcyjXQ
N0Y1sbfalexjDeVW8IYXL7vgU4DC24f3LMkLesO8/aJ1frIqehRQWNOnAMbPr1j2
bWRIB9H9GIRIFk73xFgS9lI5hWLA470K7RGyl3IvMt/WE2wOUNhGq3qUN3tPS6mz
G7rehNzc+58d7Rf1FStRQhYNVQaiZf/EWwWKU/SFnPWrTY2X1i9tlQyS4aGpaPXb
2wFdwSxUQf99b4aheILdS6Gd59lNvRDHAXzsOb8He30hSg4LQFhxtZeWvbXHsMby
oORU0N14JTpxfcT0pC30Zdo6IXGoBAUC310Bb+Su3Tdh0W0poVlaXIin+L2endDd
X+FbZi3+upB66HPlPj0/XwH7TNpJ4swFLcu3nsK0+NHlKRWzKwYYROHmFGO/82Fr
Nk6e1F9gPmia7paaNNlyg/DX3E5rrGIGUxyRZmszhN2gPWhnozTeIUCRHUDm7Omq
pkQDc9T3+Nx6NYJngSv368znLI3ENVd/Y+p46tNkqlw3unBMsOsr7KYmDCT1bC40
BggPRUKF+cFBrpwOU2XeJ4wsu+I47DPm8ngS8a42tQOTm+GOv1CtKNKDJF+rIrfD
uZp69s9kJe6+uvt981CNLWAYHCw3Yvs8VHCtI0zEI8kYmWfiGnGQdTg9Xbylb7XX
GZlsM+3nNEzDTjhoxkEv/EsxE6YqZ06P30s6ndPeesIlDVwK53RNqqe3vit/cxuQ
FLq8Mj1Qjm9LJNFXHFASvWkTHK9GQgn4WJHYS0CvCwGHHyIqhQyJiBxuj9czpJ55
8Z12dx3rgJ11Vwa1S6UBIZldocs2G2P4iSBUMWeSEvU/UbCQy9nIPzi2pYxqYQBG
mKUtIdfx/D54fqxySxJhHc99BvSnFdDMHtGvRnt4pyQQPhp0TpSekr6dMzNnOAj6
LWZ3AIK7av7XmAoWoeG63P6yX0WloI0PaoV+UnfI7EJCZO1+IJBcYiv04GR1vAcp
ZElTxaffelRkNnX/Kwl+qT42Wzyo56EnIpa/nqVqvzYOHohsVZFPMP0JWcodNVq8
RNHJDffUgZtcHlPtvsUj+I7oUQisko9iNVsiaYebS9IriI33b6dOEcKip9hnpUp3
Lp1CO4PO70lSkE9vcvvk6hy8Dn1Stim6KdWPIfozqM1s5+osDfs1SjUvsmOM3oSy
gYhyl4bjrexvXYPqEFifa4+7purs4vdhq7Gnly72NquYXt5NaapEJwYM09jTOIpu
9dC5PUOa0UpmAW22y85yOZyHUAaUMDljKEO1E43A0jOviwgWgWZz3rRBFcZgSQmK
E03IHmM/TuCjl7C142KqNgy+KZ3w3Dc2qqyqs60GpwfWJEiZmFUzEkMWHaOblKd7
GoXR/nBS08zB1y8Q5BIgdRLS9RkKUM+t+1pIOTw4Y7PxYK34R039X/0dBTsK9Ufa
XyOqJFXNJHz+WP3BFpraEemLfy+knkbYT3xxboDhTz65TJH01fMxIghW9pIheHSY
Fwuqd/v74b4c4BbJipqnRW5qeCTsDXXN0PpgXjTYmfPq39aSxbKnAYU4l4/Gbja/
PUaGOGXIVcq/ZnOj4/MPF0QSxXIvUB+SRjRBDbZjoO4LkDETdPVtIfFZo6J18kV8
LZEAHkNSnpTyhia59folrNksq2u9R8ydOjjcao91++8cpjcnRnox1wyzXOhPiDV/
cUA1mbr6uz3E0z8PUPqqeXTEE7uw/41HCuv9unEn+odAG+uhd5j8tLeegtt927ar
eubxKrAQ4OyTNs3Lz+L4Ua1HbE0WFVowzy7VDidImoj5lovkLm/vzpPZQyNwVPvG
yC3VygENrWBY/CHhZVNITdNWC2Txv0yIypk/CTz3Z95MLzQrx8c8Hpnym44XV3vk
wBqo07VMMBNTspJXoBeVPqznHISkEc1p67UUqdPkDLCiea/UHxnTgcDNAWTR9A0o
sIkIypeFN3YxMlN5NXhUqyOnGneIeWwZQy3BozmwhO5ouFcahM1RCLtog18B7+NF
syxGGwLiFeL+iwlY4srZPx1LWMuah+fUASJ+ugLwkWf88Lb+Vgp+/T6GzdWwCzG1
SyTmte1FXkGzYYCsxPZNfm+g03Jx0zUF3wN6o5dFSEec06+qJcbWzQojmk85WMif
qHky8tQkzqkgwWcPMCm/vXvI+fFkgpvUwvJz3G7IE4DiFx+flR7WwhmYrncvkxsv
SDjmSeDBDIwY6zPRgbX+jSb5ZqPrmbHuIu99FMKSX9618YQMAaoDmlKaT9BYG/5U
7TAe0oK4YiQaqNsgbq4rApNi9sIG7V6KCAn5lCX/+O/0uNOhIV/3T8fvcQEFxDvF
zPhPH+Qpy5YQQjOQU/amfUFy+fl9o49Sp15W1zx+lSmTV5lsZN2EuMi63XdNev1Z
F1rSHfMxAP2jwER3v5G1FOEnVaH76BPRqeczgxI2j/4mh/Kj5ubtQZXVmI38+6vt
F+qPhGyiZJE7HprjoZhur6LKILT18eVJhNqk1y+gfdAAUc9FdxJPKbnXGuyOpFxL
bv0C6d7m4OaTvi7fbO7bnYvc8QVJba4fm0P61JF4rmE20FwXvDJA3R4PlJAlOB+B
fpAxUmfNjhYt4NUeY4KR9yyHW/xO0/v/v0tARdf0DKAiNhopZBI8Eyx+rp9K8O2W
bUV9Jt8EyQpf+GfO/f1ipkOjtoNjkoB0uPN2shVqtUMiksGKgvGKvuqEkYamJ6km
2BhwZiPEYrKhP73o82vZLazgr+lhL2XctGtbl3Ian+/brc/BDoaR9H1vjFX7gh6N
iRFmCyT+HxUV/V/bFu/59TrzA7RH1jqmE8z6zHiXP7+O3dgZS4y1twoHzo7f3GgS
70btIuSI+MP+9plP5WwwWas1QX9l2g2QhTqKPf0Q4/aWFSZRRdECUOuGT1p8ju4H
ZB8kBR0Mfr6t1DcxAy6iD5S1PDyqdooEL78A/1F3LPJ+rL9nqeCNHyd8dM8egplq
xgztrTWe2nZi2lrr9WIqyc3ZpnNFz+ENIocbSv6pSbDtT/NwAqtNbb0C4ab4zc7C
EEzpKt/l8C5gBt7JpxYaQ+DRIj0pXmmx6sjHZEu8dNriO/9PBZAEA9cxm7X3M07H
57luBm7RaEMk0Lm7OrzZaUo+EH+eQ3uehc6YufshVxxf5fb5xvXn9eVIU4NGh66y
+sMG+6cMJ/1hJUn+gOCId0O7c0F6XAJ6wLr2OVxczNkXo3g3bnbHmyw/EesQzXR4
N5lUk/b57sDBdV71cKknyrudYcVt28rlQxWvqtIpolJtzaKzCZ//qmgXA38fhPaO
hfSR/CWt3HQIVu8ZGtgJoHcjwWWG8XM+wGmZA1VFQXi7eSwLrxiwoAF5fVO1xVhW
zanG+E8yO9M+roqMg8UtHCu5fbw5KW8zE+g0Lek77/ozHKT/wDBQtJDK2VvIrMET
rTVQP8SxM0EJzHj2NssC8RjmNHooKeAyrl1lWK2Z7nPg1wExZUoq5iSPKBUB5cdl
s4kuTLCTpH8iw9O3nRpRZaNUi5OVT188YrOjUFeGuO7cTgw7tw0O6FigzW7Kbmki
k7TkKp9jfP6ZW1EPjbfLrQI30VVkHc+6b4bMNHKQk4sUFH6ZCDFBo7qJQU0G7SLd
6FZrd32wxxjlCh7R7DUgVdMh1ZxjfWixtBaZiQVQph/Xz5RMS0vptjSYbv/U9Ssb
a8KUsSpl60+jvKjyVTFNfC3c664u/487+tfeTUlJsw7Y8WPB23iWP278zq3cljhv
r3eIrtkg+qqmkArufJWx8tp+x4vqJ5PkYfDlU/6fqWLOtg/oPcJKucSU0zQ4jmGU
8naQUEaFKmiDiVLySMkMoJM72A/GVMKD8xT4xmTF+HYy4jaZr8ugvFtVWAoLJTId
H0ytQQap20ionrYmMHWwq/saHMSVYzkGV3wbCiUqHkJIdFb5aVKl/unXI63puUCs
rPBIBhIe+9PNdLg/2Okj+fCQqGWYCqIOOTg3zqCabOQVpel9NbRjDW0Z+5ULcWFn
BE+rBRDayYvZB1PEIF7t0xtNA7/L+UPaIXVEhPRCLcpP7VO7flQWoNrXmzDR9Aof
Yg67ijsg6BL6pscfMjpL8G+QvpWs2X9ocJL1LvtBmX+SQXvdywmJmo5kVqotC7xi
W+bglV7JESvPBUHSUicbn6x30k9Mb++9izM1CKFVy8Jam1cT/W7gZ4SI85n1DgJ0
TrB9IAgtKetaL+2ltf56V1s2w77+lrcxJpBUw0CLYdPJnV9B5O/1np36BIqvla3X
WuWU/7VWbFkTsLGjmpaii34/lT08yTVegVxQZLX8J8hK1BzsIY6r8Y3F5/xDiul5
C99kZ1JVvV7rgYQcrxFLn9gl81HuAGlR1bZXBdazfki5zjLgNVx684oayeDelsZv
yoJvEJgQ9oIY2enbwgthpPWG6vs0Q3BTgGPzbHBYkHMSRM/472nPK6Jzs3vbslum
HcMIlROm3JFB/EjALSZVXBtnni//Gp5yUaycEhxBRAPwL3jeJgFuACxFCmvxsFk+
f7AzEp8hOVzpjRfp4nfxSzhPre4VB5SrUBnx2uZCil4duZmcNrqbtc4bzwcPDAKH
7uK9imvEH+5qn5xiTZKNE5Mh1QCTVqoZECu0s3bFwn7Mj3HiI7ko93x3+UCshl8a
cVGVrDQVL5C5FuT8XGxCk7oDjyQ46FyYoOW0tF3OFVSrte9MCgPDkOcUBUXdqd5B
CJjr4801ey2gejNbQTAY9HVLkk8slIDJoJ+3QfqGJw6mA4gt5/KSbi3q4C15GM+4
f4buJWUWko63TPPBkMGRzgDnW8nWCKd+cGxKxnZaeJ4KpBou56GCxBKehelYN5eG
ar9cq0nRO7+dJ4e+JHz+4ycRvhzC0rXLJ8UCpTcE0IeyMvw2i/18BrVTmdremZbk
JDqZuFFKA+1ISpidTrcGUBE6DZJsAyGbsWrwXxuKCdaM5vS7o7/rpoGynaXMxNrm
47RvmtSvvzZ28mWS3IlliKTimq41FnPFEP6nYw56ABg6QX4jNQWboXqKADHBaK3+
TfHBryKNRIbbOmVyURluNPkMsl7y0mVgsDnD1k38CsrkbZ4rOvLZ+vEj/mZi2ZYp
b1Oq1in1r57NE7X8uB+IszluZ1i6y7sBxdGKU/ULLgkHg1y5wt9vNseF5fm/77t8
+YNZYDXHPYo1sZUvizL69Abk37pB5FYKdV9Y+2LkjFCs89/dMAAhTVL6CUn4C129
YXfiN0vRPuEgznD88cZ0d6Z59ly9m8g6gofhd/TKjoD/gVjdLmAkVqpCtPtUDa0d
KeL7pabr9OesAfoM//mptXF31oIXhDTp9l/L3yV2vkEyvu2IcRKHhCiC0+zDLrpM
LEjVgKBiJnO6QBJBIPqlyYePZ2GefGU6p4O/s9iovutzQplaZE1AIMrmjh4C8TJR
kiFeLWFjLuXsdJXVHvFVvsK1GsFQ4BvYsmNp8SLGtkcvSP40YcdyasECN89Uu/RY
iEpPLdn+mD02d2p78x3IrTZhI+vLLKyHSlujeNs9LWBaT3NsYNvZGxR99xCO6Qws
QGJxzx7ExDcSXzd4nxPQ8mdqk9NZOdNhIwOQ7mWYJe0O/155COx3XUEwJUK6SxHf
ZB8EeRegf7bEDQu93LuyW5aWW9C3HQMlWU2uh5ZZNvqv3/e3oFeB9SRGjMgNDeNp
3nS1tr/bB0arlj+G4bC3w0/azzPtU1W2Sok86iD1DAqaf6uFecNqc62mRms6SLAj
hAkWDBstzTFqabLGHNwE+pvFtj3v4Z/Ggb25k0OmeJCn9Jucb0DbGB6qjWHtClEV
ZsQ+lgh9I5Tf7DHMUbbD8JPHz14/sB+yfTblymO/3uUv3Wq79lxIFSDHP5u90TIR
YgO2z6xorr9Xj7Sybyjduysjpv6av59DsrrfXwH8swEX5Dou6FNWUcCySZZJnEpD
Ob+r0rXay+o2bjbWawj+pWPCz18TfTB3okWTnmEIlNK5Wc/PVlx/jsI/o/UmaeFg
dONCHRHkU4783JjJNCF0cBr0VEtQ+b4aXv9cvijeE0sAAkHJDNJAWFVlt/9qJjzb
2FecAm9uzpjffiojFvE5wsObCM/sRGCrqlSWJmxxs7tF4IZrPqwq5gbArxXF4ViX
R2xmeyHMvEqk6CxiEscPkWB1v0qYxz5G5AfwsKSc9cTLxfg8YPNcUr+QyUor38ok
i4sxYJGWqES9kbgeVk8BjP+gOuv4jqleHvBxTiB6fxkh2xjeuSIZkJxF5vkzLK3m
TFWSlc6sLyFnSiDKGK+kF62S1E9eXt4LGuyXDPtchqpMry8gYjgtfKMAmNY4O1rn
Wg2CD3P4xldeL6T4JOKB4cl49FsqJawUu0JYt+Q5gIyjaFWzHsqoVc+bzKawg29E
2lUbYpfM8H3JHur7w3xFddEYKgFIA8DoE9NQycsr2myrBkk+DdFtoWwjg/U5/3p1
3Vdg0ZvBSb8DoyPfFysdCnaeCMbA5epzHf40OaGxphtCq/gMW8yxnUVy3uz0MKkv
ZQpQtOxKG1ykcum274hglE0WXmvOjnNT1nTiW7bdaeppA/UlYYtpgwc5yWqnpMrN
RyDXBdYesX1qZw8Byshn6N/UmcATaNmoX7wO0iVYFarKoaq8Y3ptGDmGU/LyYZO+
o+ocHlRmiE1EQ0bIELdEsoSJCM212GLTHCkFowCK0ZGayomSPD2uf6pV61K44CDO
HPwM5jYFCTFmq/eoyk/DRBXBOqIANux9A1w55hgZpllmGHbmy0WHNRBq3YiUnkiJ
F8dxW+BZD9xidzKxdA3lKrIg1HPqZpkbu4xXfJQAXOFT8klHvFuqKqFBvP7f0CwU
xjod3LhUUyoBMzo4izMn2tRMhPcB0NPZfcu8gf34vEUQXUtaLRTNLxyvS+Sq552x
EDDUAJKUlzdkbMQj5ic8gbSaUxKl6X0MhyiL+tjpsyYm/TxJCj08vG6JJQ8781u+
3Ojo3h0iZqovpTwp6HjvpHY2tmHG9ebvfZIb4E09PrUJmi7TAWad0PV4R5nJHYUE
xscE7iaSKa9KwQYdn6kxOqMo4SucK/Q7DVRE9hQaGOOHZacpVuXWZ+yATuxLBTwW
/Q4nI8RV/OkhAwsSU7x74uXpNYaPR5FrPRvmcpvu/q1wXzO3FPDC0X8FJxLZ/eTL
v/vRyG6IOvWueM1S0nDiS70DaANFkNktLjHzQq5shQBnwB55WctjLniFlkY1qXYX
mOvod2GSr0VbM1bs3GwOuu9rSEcmsXFhSf2grm0TBUIP1IKqNPSrW+IOzByn2Wpt
EF3W/NgekaGz1J/1ZTM+0f3vyz4rGHfh0LtFCeXt9Z2HNtw2AA+h/iLGdPrK8tm7
KLELiMF76h2klwbvJjJyhlBEgENpIBdFWU7F2BMmCTwKXzJFOIU+0i/ZBGuamQ4E
YMZSraGPa3k4UeKMauNGnqqofEHqgPcriBV58SBV4xtJmjHfWZcSAh2XIKxHI+xL
PoJDBE1CAcl0GrKhIAi12cW7ycA5xLm+as80sCX1y3QTrSzWau1PeKoDhICn/qE2
L6yhsCQ2nneuO9f9+EulQg8BdnMDNKo+yq3en7KBHC9ss+kaZdXrxiDcq9NDEAYK
MW/N8Q3lXpBvbRwSgiG/R+FUFqP/qCF3IJRzBCOTv+YYp1XT9YgTMXf7Aq95rD5w
Zqe+YtTczpRGV8T7WE+N0R8nxKeJn+u3yhmI5IwXQbS/P7nCyjfzsRnvmDzZKhQW
padYMFGYbRVsHa7sNP1URr/jlGTKHgAw3A3hZR7S6ImzmHauvOwCyuF4FPQCqV33
6uoWTCk42tP/HdetpfOZsaJpUjf0QVdKNPOdttpHafIjQOQmI9md1D+F0HqF7OBT
RtGyYDJ7uPxwMlyEd9472zE/dsYHHMVbsj7CXREIGphojGyb4wb+L/MaMstc3uNP
X7VS9ZPsD1RcssDqkmq75r8/QkbxIyYvEKuN7uSRTrOwjLA+FEAYvI6AWjJ6pJ2l
N2bfRw7XbsYjqWcZGwzCrXP0TFxbIqicFmHESgFTeDnnrniqCHCsLutBDnTBoTTV
p5QKGGOhPwSu+L+ZYRNj1NNMKoESIrlAMD1wegPXTIqAPqOTlq4cbrpvm/NLhe91
zRuWtHK2oeTIW4BfmNUuVZB9yZoCqOfteZup4kGd4Eh4BVA8XrH3oBAbLOxsuRQ5
6frMNf1jiDOSKP+dsfa6/DCDg/Gs/NUWqpSqd+HzqJ1lrtbD0g0r2WXIzsHp7GJJ
9SH0z2c/DgIhqgY1H/lbY42n5d16lgYRXqXYsnl5ogjPQWtRWLAhcRN2bP5pk/jH
Rhm8vzEGstSi5U8C7yAJ+4QM6kOUBp9DYxBmpYORFhMBXzzteOHGgR06OK51Xe3U
pwwf7OwZ/jmHSnak2COinnIIcZUn/QPmFhWqXB+xfmkf+w1/Px8iY75OBuFLp9Dt
aAJ8UlJH72eodz2f8jpnXp7lM6uDNfGC8xPxsw166DTlal35cAGuUeT2Pfk/CBDU
a0BlibqtWgh544KJM3iFa4pES9CDwEijrzmYUD6yJLXQdQ+WZ/Vvi0Rm3D7uIHIP
4m5L0grbDbTG57DwTFEigi7n+N4jKUsKMxCeW2hS2JZ7rmZwMTt+zeWvaC8TIePG
EU5mN5VoPhDRib+cRkuOT6UunyrtDq+ZQV+on1iixNXKQ4Y0PrIHZKg0eZHIRq7+
rTy0R+POfSWknS5dVIQDhu2aqCy462TFjqyRtsyT3TGMmWOUsNHAJeRJAm0a2Mbz
9l2yJER+NdJebyzxRNs7L2BRRyMWX1G90o1WbtvAwQ5u93c1uTqrOPU9m4oDnVDN
3ZIyKhNua+pSR2UtWrQf7qY74hw7kaknf8Zmu37q9N1i4sWiiayAlf9QkHXErYrE
/fFsI+59uttLrHovzLiah/7SX2lSl2xH/AkBDPzjre3e1ar1yTmdmWqXH2co0S26
IpS8dncJAjCsv+rAwPqYCTc0UGjtglPjdgxwFI3cfd6FHeL0uvssHCbYciVlut4P
xfGgL+42HnswYXTtFZINPWzKsDh3As1IbipN32YQjmTwBMmffd5vardoOz6J7jv/
wfT3ElwLhcLJ6b5gSec/B0WKlg6kgq7I6gb28HDqYECqdLUx+0JnoGQDlUIzcJtf
yYfpuaLftcefwG3qu6LQuM3RAO9d/9yIwQ0g0JJg+8qhFmzpnCaVsARAkt/3C8qO
pqrSxzIBoh0JzkVTKyfdL6QNOleWowQIIoQwptipsAVe+q/qSo2W2CKZpMWByf6W
hWjYuIAOh0c9oVPJdWkUZUOU4Y9y220qhBi6EGlze/QU5ZIv4JaIAO7yh43xD61D
extJvKINtZoMv3piDYp3/imfzbRKKz8GbA8h6F2NXDAkeJgFF1YPgyTpbs4Hftdq
4Hs6jLUC+sNU3my6jrUP7GfWeXP67x0PpkDPiMNA8hg9z8bWsKEXeRrTSOT3rZBc
igzDn99lu3IC2gX7xJ5bx1EGi0Qv6LYXoCQOJwXLz4vBaGsRQ7dK29A+L8w8x7rF
pPqjV3FYRt/fUNbu4ehU6uhwfFajBtXo0txeBIhV+Xd3fwRKjAdaOukyKGfkjcWg
WDH3aLY3tFaMknDG+eadKZKqQKPN7ora3DWT0atq0LThO0/opMaj4oRNrt027czw
utXzhy3gvMmqWoapUWdsA8dmDchmqVx3FcmyGdZkdH9KapsBZi1PbX0XMTXES6OW
1jONq9WBWsnOGmwNjL/+qWcgzmwQwApYcAfsOgwOjtyRZy0j7Quv1n9LzCb2DrMW
wR0Q11WEIjT2EohY6hi25laaK2hJJ5RkvH8lwNs0Su71njM3Q5mNfcod5Qa1e/mY
uPcWFSqXVpi60BMO5aoSoq50gWcoq/7JVWxvyDSrcGYfZgJmTgDjh1MQHxaHo82b
CnXSnG3ENZ/OyWVnwf7s4W1tLxxtw6L1fJ8a2Cz3EyQhq3bBE9yyXvHTstRQzVL3
wOCoI8OXpTBRaNAlkAKRyBVc3DuQ5v3BMPYomQux43oYTPR7ZoXcGM9EiAjm/UT3
JyDExalK30az721WlFeU7OKHu4q3AU/g4XIeXza+VVThEjCUftEP0rHa4ZW1VIUY
24lMeKZ+CoBYeR6wBbC+bgHJx0tPkXf+UgUteEAgRHkS+cnPhEp7ZH+c6VmQ6KNA
uv8kUTALQUCJRuZdReAvhbjUvGqmTvSba7AkEG/rng2Ql0JVZy6c6m9ZQTtkJTTj
3zU0BaaBDpbrXO9UIItZ5maFqOiYJ60ohRqlU/ztDtDkM2hkFtPvpzVsVe5k9eX+
91z52VpmSPckr0CDYLimMjv/YSnhlSRcQ2rvlKGhFXj1cmRj/e7qrSCN0ELB/biR
+PmuckjjRG42VJRUTTw1ypcYhhvEh+khfF9kaK4Ze6mJiU20hNLe+qLhv5LRRQ4U
O5wdWcKsaggymJXWhE558WLpJHT1fHpEcrfR2hk41zUx9lkamdagDIkaK7l/4UvT
zx6XHEKSCfbfWIrKONlhaqB7TBgYS2BEWR+I7DV5TDAUbCs/dPOozylsUtKBswng
ksK8JqZlNY2Pg9samCSh4AtgId+OGCNUH7SigXT4KzX65kl7RStXh0m7v4AJTe06
0RRhScqUs5SBBhOQHOphu8+d1XIQ755yvLan7y91Vgo2UUCkRfnBKYBpDafMv+M3
Nfsux0e0MOyRMgpnyRQT6IpAjJy/clZKRk48Jy838xQa+9rw9BSOo49+G3W/XQA/
WWnHECuCjGopd3RpQ9iTn3LC642Q6wRHDFc/QktrjbX5ZqpDUyWhUIDz50KdGbso
vMnv/3BmuAoHJA26zMe+Sq9WZ8CgaI8n53kipo11+obN0kjHKL5SaXZNSTM5388f
CkYShXYT/uMHjsGDZl5xi8lnPo+1T1vHHCZJqSnIh0h8ZvXKtgurFlMECtMaTkQu
lZvyERcAn16sfxPr35iKJlNya+CbMmRMNrFLINRvs9blFTGkyzjbDLDEDYSS/RfU
Oh1sH4xMbiw422TDtoEHw70PWO1/Lxu8/N4K1RVjWlgntjMYB3bHjE/FZlSoTcv3
N2LbXBxphZfxRiZT6Qy8a5qiNW0fs7rf+EmK8bzZTMvhxOC42JS5raZ33LyVvijx
/DvavK2y/2cUnaHqQQFIj+e1Nlax0XyfpAYlOuzQLDHvbnXHLBd+C7ugJxWBbi4I
APAyQvdVJ1V2oU1VE/u/apVNaifZdwtDkqDKDCl7qspsZaRUDtPLzGF5UvYa/6LJ
nAZDHfwCRryu1G62fym9A3NVEcohoxUR56UEoqo+EmT1WFHACUSiEM/C9OMWYbzV
flKAdgCuNMfuMYiGboiHmFo+jjk/5FVEepJOtilhpStnWiN2fWceF1HWpCR5QboI
yjrtly614Gpqk65OhLUVphF56oTr7mF8lznLtn1Eif6ABLuP8jpERETVkL0RN1sX
VMjOlZJskc1uCcOLp+oMTJNTuhVRAqZeptbO+ZLEd2F+IOQeg36OFNaDVwJqdwqU
a0Mao+uNf/XAB08Z6DO0TWkt1oM5Px6O1uTTJ4O5x3vt93TMPK/+mtpKDivee6me
S9znoZ8kgUQsgjEtKpbu3AJXp2knLgZBEAVSpcJ/A2bp1OdFTNFjtH19IbG1xc13
fif6ev/WsY05HWsj2eXG8/gO95YPdKEd7BUgSQULBveyq2FH6oHTiOADAXipUkH1
//IuYgOtVoptqou1v6I6tmLev8LI+3260rwcD2t2O+nbtJfoHs8zp7UKjGdQXVrp
rmCRXIQfnJleNo6eu2h8+kiLkgiQtYbKDrkR9l9uStzr+u07DiHFeklZfV0XLH9q
wICydlG79lkccyTAwv/zSN0MkYqKiWSeGhblJNwz8GF8wvV4+rFFKMG9EncGxpwg
K8+JOe48K1uYfi+kqGaMtkHBTahwlr5XrtaJc6f7zv0HednHsz1el3hF128FKnWQ
V3T605YCK/rtD8nIPEjetyYvCaS5spDkZ3wqbgccdFMhldT9x8YuhfwLd85heHML
GyaaBrPXDFaBKyn0+xrMPKI0wXEZrtJOmDIO9q8fUGmqnS/mfvybr+Zd3DYCgCoP
33LGJES8YtTTX0w0qlHv8Tobr4jroT2HjWYBYuVTBwtqi+i6MR2rbyc0S4V42TVP
rKrIV1t+lbJClfN08SUghvrze30RwuClzDlbuIHUuS7XS3zFfxIhXc5nqmcMWVir
YDMzsEvgLIzBvVLF7K/z7c5bBcorqpV2HjvAs/ZekxPdVwfpVh5q/hb4OufpSO/Q
/wHJP2weRCrIUgrgFNlZQc4GskppZS6+PVZ85vAVLiAYVK/HJUiqt0djXG8IV0rD
pE05bPEoBm8WYzlfm4adypWuNwESY7pVH7pS1LSnBWCHNc0tpI9O1WM+CO2eh3zN
bNgHhqz/vDqO0ziZZ0iXP3UU8G0hQLoTUSlJm4nQfTWFpvbOmrHY6amWXJjDjDUW
y3olPgdE7yZF1HCf/mI0NEy8EKopTr9IG2iup52FHzyhhX45j2lhX0FPS673G41k
vuOQmNUY/SS6Gm3AYOqTYNq6Ttvvg8ZDbbR8Ke9y1GxDo9rPXPifEkPkL/b+wfn0
CD6AvQfbKRqAbbSwPmQsU/xcEsHZ6y7W+uihFxWVplXK2VRx4xkA1RHw4T44Kqbt
klab41wqgKLA32NOt2oII73aUc49x1omFk1iSawRhOMu/F5SmWCFiQU9YcQ2bJIL
OjMmW/yaV5p2EvHf2T9eCo4Il8PHqEuY/taQ+/h73XDIHvG0sPnJ+Z6ZTJ9XYoOz
FZ/bschS0gx54X5cQPUnAkNMkByoz35EEnKGJtLC0kdVF1pFPzQT1pWYcuzERwDD
TcGHRoYXj5XMDEejWeaJoAi1qhu/isVKXJAiaceROHMx8CemBFMvp4iiTf6GOepO
zttMFqNaUvUxlrmKrwsfSk8UotgCsEYaNE5c5eQKi5kaLeyLGohycC9ves1uqxF2
gMppwW82JDEJcvQmqDQ1miVAVPZJy9rOmdnoRnfuVgY+nSFxZsRZHmilnG6P3J7x
vTWtqU3W/qpXU6W4IhBUK5DA7+SjNZY8T3LoddfG0CMvDp3dhC0Hl4byHeQ1KUuP
L04SZdPJRCL6Bv3Ezia3Z+9Kkvfi5p9JLV7t4TywIKThYyTYS2mfpJG8LMEMeZFk
SXE0clmfS/Ag3entoBXvEV46LLDKhm+ejCd3w4brpHfWJSVG5uVniTeHpkCcEHI0
WEn96h0KgsAmJgLssU1WYVd5L4mxVNgf7xNiREuYIPO11otBuet5bFEexO5R6LkT
HAb1AKJg5EVfhuL+Yl+tt8CNita8nv1Zs3CTDHngRjlE45Am0dHkzp+x5NSMXERn
7mqU9FH9PDey9t+V1WIc+4VgXr7I+GDLnZRvtYYH+7wbz1FsyD8TTtdKg3/xqhLv
tLMCpJVVWuFjZBh+YcblrjWKIE4rWH1PnWSTK+ZIQw3Z2a40xQjwfrPlm1QGZRq6
n5k2mBZ638j0n6Wd61Vw8dmUR/XVh0Tt2nyKa5yn7UcnohjJEQP5/b8p5Xa3FndN
9YXZk4cPVJ6GB+kp6lQcOJ6yrDqH3Z8wvKhh9RfhtbjP28IyLjTAE/kiF6Wfo5pg
MXcnBLAJdH6jDW112iFP9g6GZ9PA5d8bUgsynd1tOtEVmypSD0cAF3Nb1EqULkjd
3HHnUCrVpuLuVDfXASdEu92nH02lxHLzatIHUdhNaRrMqoEC3gqW46r7os/oHOC4
HyysyO1ZlZ6AxxhulQZIHcd5jdW5pWnXxrou6WxSbtXmLMiOVVlJlDmy0iBi78+Y
dbPpWWsTiWNQN32vMB/guzI9Vd8nWq3FhmrKVnSaO+p7s94EXMpjPyVbp+4Buoo8
s7SVpjsXg9vqpJ1JjrVktdHZ8PPcQq3x/i1ItEUBIVKQ2yJbmtdY3yV1kNdUJzj4
k9hToZkhi6d+83YEysTiGugKVaxwUEULogcqM4i+b4dV2XIhPFkOgCRKjlhNYY4h
T/FVP06PHv/bz2RIK7I/ihpKBPG241Q8bOKqJlCgqTxQbTiKxk5QWU+0HrMjO5Rx
dlsIZkGBszaZyfVYakHSrOKhbOEGKW4WUkzGsoKYor9PdO2an/atX5k0EqPeo63m
3WWWv1LJcQZEX7BXM+EjP5NwQOiwF4/tSm42NdmM/Sggc6NIY4gJNRWZeqTKVv0H
oIGn8xlWcocBYSCdGYTCw+xyZoZLCbhLYC5jbvxdAqV9f+nYlFhMFlHoVChqfP58
HHjTncqkpB5xP7jbjB0GMUIBJ1/YYcAs8wRbOe2vVxO9kBctJKigG/3XmH3QY4t0
TALGW+sBzm91ggkhW5cY8BqjDyEPN/Xr6lYAEz3mtJtvhMQ8epj/6hLreYJcUHu2
9lwVR3e1hahrYJegTXbGa0kSAKRhV4MS1E2eR8ZJF3mjpl4uXbFQDpQrHZMxhb5k
Z3mIcAe8KmKtGeum3Y4Y1n40FhysGAKAbcnYiO0ny0fTcVtbak9ytuJtnGMMANsj
HcnpdwqquEmbTy62FikZMUdjuMgmmZq6aKSCH8duF4hInM07LducUB61/Mf4j50x
n1OGSETD2h04h7xB9RyqLRNFB4jM51JqDhBpGvDe9eKw8640enpeJkCcLPQJKTEm
uG6pJVDCh586FxEIYq0uTDJfuEmenTxSPRaH7QwrBNi55abXkIv6gT82CdYYNtXS
IMw7fgjg35nO1ECBM+Agrpk5ymSBHglQoaO7R88QOQ0Fvh54m2BRklB1zQBGiuPl
l/y89kclgvH1h0N3d02xvwk0rB5Vcc7cHqaXcPZNCQ+THTH/qzyK07vw1Dr2LKhn
UkaDpCWBjBiInPJufoP2USBj9ih5gPi94/pCrVoF4UH04Cp8SjgJ8QzA1/IfOnLY
W2rio9HbdUUXt0iXDYCgoZVSm2drLXPTJ14u28M+sNk0qiYwumLhW/DzekloH4yK
04OHMaGZflohhsLIOV/4vrqwm+pZYq0P6m6ea79Di/MUC8r+QQu/oB73PKg98Lh2
V4fORyCJ1dbZ+9nw1ehzt1YQk8rW19WWgNPITDXmuCLyYyWg80PL5rAY0+QD3/1u
VJZicupxrApzg6k5PiyHO6ZSh6X1aOcvSlxPDmddx17d+TC6DFS8ki54Eq8jtyif
3LJIkz4b6qq+kC8bLaE5ZKInL7WDIQrovMxAR+VoOBruuMSIDo6mErFcTy6h65wx
0ND+o9MJEgQ1PdiyO6+5PaqewVrAHP1CzQMuBXMXOWuJQ/IXCpzUzWYEousO4ZWX
azaOxDa+XcNn1vo5WL5Y4E1ydXZXnMYBox3wQd00PwjDSbMeao1Itfw1XsPCroCX
dpS0v35aAagWf98gHVG2xHD7OmSEtz7xx21Vcq5PP0UFmzuxzyJ/9F2OU7BvsTD4
QxovoQLo4RGpmlza+UigCmhCyY1otrls8mLuurcOFZAn4mv/SNiXq6W4Ni/SNtIS
7/sVRHjsDZ5CcKQGt1r4JMro6dL3Y7tnwPJNX6bm1XgOKz5DYd6WYgRMbYkAnOfI
WXZBO16tt8JpNUmIg0GhI5owH/emK/Uxnl+8pbQyls2gOeoAUbCaIi4CF3va8o4Q
2fK4gCYJDN1UPCC1u6DP9WDEmjxsbBdm1GfTRz9gOIklcwJuNwoPQXqJyCj9sD/x
LL4TRNEzZnbo267Krdha5YsQ2NvC7tklltQqxGY+uMLWbqkyTHuDuqXVcLmRuZ6i
hHF87grhPFucNYQvrByr4ORgDG+Db9UCx2ihxkRzo1eW+smRngCznIp/JXBUCjhS
8lLFPrnBbADBlp7sb19x2f7zhY9Ttn0mytuc5FShiLwZPnC/wNYA69syLqPxBIeM
55EtuJMKVPGezQQQDroWmI50rmcncsw/aqDBxl81CjNWKg32MNa4CV8mZvGcj4Mg
8G74WM9JrnCoqVSUEAeJCoFH018e9irOuC46NaPZDBeaSu2on9qpdjUdF8shfbEb
At9kT3h4NxGG/oy3wtw2WRuxHCbkuzx0/0ceDpTI4YzRfsqeQ8yhyhqGjfBcflFc
QDnI4jat4V4bxkrcDgYvBZ6+2x28WL7fi8XjMZs+BVM2POZFD9wTV5D9AQzy8hQw
BnvFr8frAgrIGb8XhFVsGmZu6X3rMJ/KqkHJIsQfbazAPRZAj9GgVHMi38HmO7z2
8AegRGYrPjRFybE+cb9vtAocsefx+mb9tXmK1AF5/uExxWw+YzI6Pg34anieW959
nw69tzaZPBcCSKgNf1W7FjPtk/SiuLe61wAWzPTvIyqLuebdLDD3wTxQSWSYdXVx
ZoM3vGIiLv/1Vw60r7izp2lmO0ylB2fXIqmcjhqSKOWaqCUZ/1JdCErTIqzc2zs/
Z7uORuvJq2tyD7TN6tehX4ThxnZ7SzfiV5sKbIbFvjEnstQ2tSy8jmOj68Nrth4s
vRtJjwUFwk0hgWOdhFhE7fR8Y96u024ujIC3nLRcJhP1WvBYTLd6SzM073Zk2+G5
QosM/LPqj0i5FqbqGpHVcl1/KXNUPud4hnKcCsCIzx29e8wK/GQrig6VAEaet9R8
fJn/8y+PlmLrJ73X2ZZ5oi1QdMFcCc+zyoyDtzOwaGhhmwTHSiFz+n0dJ+pGQGX+
L/Z/hGQ6crJoaJrhzoJ9S4EMPxbLoCTtPPhrOrPIEZM8pT1nkyhoNI7r27Cd3ZLQ
y63RKnca95R8nyCGtWXzF1uHN/X9YS8/P/LICIWUNKKcNrpcGQ06+x6MYNmkMdJe
5NurWDO2vCF5T7EhSnw653G15IJjrvlEonc3pBUCgPtzX5wzoDdXFZvLaci0zU2S
eSAaiy1tuIvRVdfN09SU0YNplh+QuwKNf6juSp8jWUVYN57lsJnXVm84Af1qW0Yl
Je8PCiB6LU6LUW9wnazk6fxOmYO+fbExANtPvud0sO1FpXUItQNWu5Oirm2HgXry
21fxNSzGrD2PYiPIGzubxhZiGBejpFP1IWoMRbai4Dv6TXvngATupLc6qqTV6wet
nmjG7YOak1nBIAqXmZ3qdRyMGOkLNlVZ80ikRd/pol9Zl/lhP1t+a1nJCxuDSGGp
Ct28iPpQJUYcBkSBef6lDtBYKjvbVH+PUtoJZsxkEFz4xUUOIUF7RCqDVOhq7eKz
cfNRy9S5DUXJFUUc5x10KEUtwthvCF7vzynU4J2vphba4LCvxDTDkybYOaNbl8mA
bsAg/r1i5q/vglEbOSDN/xGHI2XPUyw+JmOGvtcwT7RfaUEWr8qlL01o5nYZYkOm
aTqGEgnrUaG2c1v9CXfhW1X5Dyd4mt4DbRO878Tk9RBlKHtlD8WefyOO8qAelbd6
LO3p5sdWWb3/uwR9CkH3fx1Auvp7hc4sZgesdwiMLog4ql0/r6a4/C4yQHUvUz2S
5E1p4cz168j2No0H9FkV9ElYFdisnBRQpaZUM/3mD6hrVcPGNtC3taBvw5qiMpP0
dnGfvLEj05YXn9flXzxqIIk2zakvZWKhh/KIpqf7E8W1FAmApY7x4UAMGC7J33SZ
Wesn9hZDRwQ+S89NR9uF1DkjEymx6RWj1jhHOqF7bJ8Aa5pbPHKjIgocVBTCgXwu
SHQkZL0mifmERJx1r8BcRFDLjuLmk1EikGryCHzHdmlWYdGSnsawpaAGbXFiJ+eq
rui3urK3oLCc/iLtbcxZ0He7jOAzKe1QBs/6FTDGVItqbpOAPuaynixUE/xVot9i
POcW2oc5S8AKgbNA7Se7Ct9Mj8O8CAA0I4/C2JnQAuXF/s4DJ31UehkuMPkGQIez
70GS/i9UvtYagAZqQ1cdRAlU+7ySWJ48NTCMR5MWG4ETJRg//20pUka4o5+OKJ7E
h1ialp60jWz/Ph+Gj4G8A6Wnkxen1uFondPc6F4rb6HBE+9I34xFK+GmvXIm0XUJ
pyK6/9yoYq7/wi2+e5BfkyTN+jW4MMhseqHJfu9lzV9zEdlfPq6SBiPe5URMtflh
B6Q5k08SIE6uz+xzUi6tLZwRuzVJ/q+CWlQQtEacR5fW/xy2bYgieJdWqs1lNkGk
Ru7Blcg2pmTyj4Dv7ggcMILq1MT61VkBILjgFtvqholkbUCzDkfVbbJfZLfe30s1
n0zU6MMkEycLkDh8+8YGKaKS/zC5D3TNwXyUwaMW/Fcxmk5ZdeFp0Hrj9+DwLYDk
yPxI4x+5vyL+xEJae3UyoDVQWwdoTiAHXNydfTUpgUcdAIcJkC1o7L8ELiyZ/bAA
fw9418bAn+UMyqRkkf1SWdIO3hMuQA9H8GFe6FjrgM8KJNLBP9ll1aKqV+GY86yN
ulDhZaYRNip6L7Paq94Xltz4jCbJ+baOtRH9aIBqJB/LwupWOOdB/oa1ARc/fANq
m6957TEJ7rg5VPzuK5BM541nV54ol+YKF4IqbkmRK3yWXjohXvZGZBZUejl1Cqao
hjK3gSqJwBcNGMDk7336qpQC/eovDzZ3a+qfCTwlqTrW8KC1O2PJQzQofBev2chq
7JwHZvenI4HNSSbAszmOWnz60JiqiJQOm5k516s3VkNe8F8iUjhEykNheSKwKPnO
2G84IvzYkGx+SgcAthIcUDIezyo1Wh2c5UdXyP5x+fkEwszukYnqgtP12Zv12Db1
f+P5qTNHV9yH4EwPkauKarOTdO52jacYwN831qwiMjWwzn6oKdbv5geUe8TeUHLe
juACLnV4e2w6wf1dcSFJAOzh+kFBPViScy/fH+xX9KbETn7+65YOUw8+GETiP1Z/
sp4dcNCyprYZrbcSYU1/+DhjUHyljqV3QdzoIETVlc3PfWQORq/E6qa77+OH1zNh
cXvwcESjHAQliulZUgoTwZyOJdPwhN1Hbu1DJuYeWsbrfTCJv2ZO60B2WFxWLmK2
wsWWvxh84dq/subG/gG6qH33gWIFkqzVz9BjtOwpGpWMmgbym9Yf5EuEdp/lRCtV
BMxZqxojk4dgE+tuZEUBouX/iobwcs0j1+QHWfHr+4WFnyp3BfIVRjfa9DEzIgZU
EWyGhBzYNUippJELKD1cCygR3i/i5F67dEspkcTx9YHu4E1QQFLO/4jW6Z4W6fDp
6TblZtwBHe+WThXiw5TlxyCBcnnMvNXJbZGjzltKDQhClgZzV1hFkDxnztU2pdl8
vyTuc4pyfx88fXlvPncLOqIAAZveMGKp42kxSQrJbP1MoTgw+iZdQZuPxqmqoHc3
khyEjhYigIzVBT2hx5x9xwtHgDbzWDTqAM7lv6yv4T2qJBETcoZ4TshywvstHlgn
pvOFpfjLUqv9ricWGb0g5Q460egeUU8xfsCcwGmd++sfgagr+Z8Fh/QHlzPpXwie
TzA6R7ngW7p18ETwTTZNQKyXfeCvbJtIvRsBvKhj7nkEzrm5HdIv5gDEmWpUG5UV
lZKvvodZfPlOCH+sW4Eh9dKq2aSFqYBsQzicfxle+cgsJlpJGtSOshZTMWmKuwKW
6/LR0LnUM/G+1Yw6gXV25/GVqktJEO5c9Gop+h4omhbkOZY/8Qf19dzmUgX1eZx7
GTFKHLrGcUISedj4STLtUJcOCFfKExJ2owkEc2//YSO6tKbSTgofjNUA5QbbzdOk
QH1DjQ+cn1KBZY1UAOTSpmlabdHyvCGZZfO1jvFBqaTA6AWqXwJn3IrKFcEloTcR
IbrSezK3gtIJsqB0zPPk6FZOAsVgAvJcmXmWa246qty3Y5ixg9r2Ty1W/+3Dxf+X
c0wkabBgfkbzS1ckN/r7LEgQVNvBUDz/J8onsXo2LOkxh4366EBVV92BxQJSs9A8
Bkz8YIvmzNQ35ci4Duh4KATXbnbK4X0hABK7rWYwNtmsWUfU8IMRjVtGEbPZZ2X6
1kglGY86tCbL2pxBQl8gHvqWZPxRNb4iUCntRXfAd7BCUTLSRBI5JiDLdtbybWZT
bcbq7H+lS8vEl1+wBsdBaIzLCxwHpgo3qzjXYjkqAdrxvHOts6Rl4CTnROkoeXKq
ZPxKaDM7J6L2Aiu6trG461/Zq9/ulA2CKgngHv+X4uoVzwqVjTBrH9RmQmo7OiJp
WSqE1OXVTUsPAblm+Gflc1QuVCurJ38oNfeJ7il54GaiM120m4Yk1vasNUZQtV3f
flxky8AirRMiE4+vBpwqA5JU0veisGpNX1GiMPYLm3g0HUBvguktsrC78b7pd7Zf
HZ76dHxcsnhdm3GeD4DMqThrr7UYjUuNyYm6UIoyy+upGWvjR4xdQrNrciJ6XQDI
2zR2oLTg4flWmA89Mygrkk8Knfz/kn93RMfx4CNh9N+ezqbP2RJGgSnYard2kjXT
fhtL8VemI00XTfutoVTrmPRGHnAYxul9DPrrLVHCPWZoFxb4FBk1dj23aZu4FDXD
Znr7hYIfHyBs/Rq2fo4l7Xiq45/4uypDVq/9Ie9f5uLDb8DGry0fc/hA6wickQwu
2mjzN6wbyUuNu+ln7sKm3+2/RIVQBR4aYmTUTmysC/xZNqdl43xpU9TuXJ7ZVIbx
ieWChc5L3cgN3ysO8L7ik27JdbluXuMvczNIXqvc1ccqw7toGCtsDmCt0Ri/24Y7
6vdcYfQISVaSAZ7vKPXG9uhD8ODgGeMJK5TNXR104c45QXy+etIc1Wyib5PvoWUU
NXaaOh9YZHGoIOGRdlmgW/b9kK8m9VkChNC0aKblr7mDTDLr87/ezcf6IpBha8wz
0C1XoFuP/DJjeWQ9WklbNZwkbpNMiVZACNiHu9dOKAH44RvmZ9epMX5EQ0WjwJGJ
Y1QKp5uoArpT4WowoDwwbgqG9rk0ZUoO+NBGQGJlr1hFiC57C2TTFHgI8rmF34Yp
GsWnb+q5HALjW3k+TiBAKiBe2fsyAkwRN2pbdhkOo7zriTi4opZhGAvyN8hDZ9iE
TexA9v4GlH3Kv5UkOBygqP9lQfBRnjit8qiBSz+O3kuLRGZE7R5q5LwhnErYkfTi
+lBK7lag/4HBynI6qeIaWPoB7g8j2p8HwpTTLhkn9qrXWG2AGOsI4yrHsWiPWQJ/
pyHgJ34Bp5AXFqRzgUzMEz7knHyIKk5HfUDNX35+Fr6IMvc+/Bz/PW2DA4Ak0PXh
Ddz/xQDYeMXu/ivXVopIUZ5Jxq+THtEXAP7vs6rAhcCCHKH/VMEXJpavJ8o21Z90
MkSkGzOQQJfliBLgFLQLlAwc48Xoc6xmo1CvpUumiLeClPlPlb0ZSEx/yUl5x10x
xXITBXh09QWugiDQgK/ne/4N3Gy0cyYH96sOy6aXzG6kmQc9N92/65TXAsunqTFL
FNJdAn8nWmL28vIa8rQqCMy/BLz/o8wdfFnZnlIpo+TYNQHV7d5pPx2fDWJ2i0id
LOrz3YSVANr40AfRdF7YfXRUN47gYzCSWvIUIRVxU4X3AY0JVx1TnFs1W9NmdkAz
KRwXScolnBKv6PihJQh1pas98piJ21h+dA7otTLJRrDbODSJKHCuaR+sGUousf/X
mwvZDfbtuotgfwzlxKfE/mExmmBnMrw661kBk8XkaAGj4E2BXE4P7SIlXjsTUwuy
4Ao1dOxnkOa/n3xB4Ow4O7GEFwIenOJ55HwKLcHZ6qzvF7ITW+cJqT1nHgYUWNNd
E3CdeuXkPIlXlhP/fYta4wHrhypQyhLzsO5IIdHkqRqTrEW2KpAP8wP9/h9SHZCL
esB7eTy1LDk5BePYo1yxXxlEkyjkU2Sv47PTcBCThHvyv11GKwNSf+e0yW0TspSP
W3s46uB/S2H5zQ5KEp2rFN+KDc+wp4Yr43U63xSymM3N4CJBTJKZTiTOL+rnZG5j
oYG9DzwnyTqhVvW/swUY2TPiH6tNkaigATE0VynZuAv1xUOrx+fsfBdZgm1PjEMl
4BqCcyk5y4WSfYHWXiIbQQ3P5iMOqVeCjRU+kh86EZ0pimKPfa2GV2XkYJMtF0zX
r3MNjG3RUbkGZIq08+RK0g2wGg2zaiLDbbcibkv3XZDiMsLLzBxuwNBf6mt3tUiw
cc9b0co5V58571rOpu9mKn67iEtNLQNF+f6GzUL5NjoNsMTDoVYIcf/ckmkT+pzR
OCKyU5Huyfa+uQ4jvCwUAnmQrlFn+rZaDHvJAkjrpIxZg/s8+ylnWfTtBVZAvcPW
FyHMx6QHEu99nfkbcH0uCmoS7xCjXPAmazH/GoupRNJh/s8U0aufnNotlm9kr2NH
KX7MShs/DJ0TdjmnL/lxfVTqp96sUoVw9HLViRGq5hhFfE91TJNnLdYXUMAYsFPK
GGMTYViGkAllWgG9LKlOSwF7vLC1LY/UIMqbUnKvhX/FmJF205fJY3ZXpyPjKTTY
z2Mfv8C1Ey5IOOVZyxKssme2JaPAz0hOHINNJmDEk1kwtMAdUIso5Tp2zO4KrfwN
ymOl8c/aKwU5ONLMeaw5x8ms1b/inUHIWQOAWWur42jBINhJmOtPKC41C5ODG3YI
VMswqz/a1pAb23LTANDncyOhWYn2ideTY41Az3cJV0WdVMQuWFbG82Nu4UUxPFT7
Ud74v1swNEhbhSV+FYqMgA1sJlpvWFH0i5SMCPi/FbdoMfZSKx5PqDugh4ryjEVm
ZVr4kloQJ82XQckVefeFkUKYXXFqzjddPVYHPlypBoynj5EDk5uf31LepzQbmf73
pWA7p5pNzu8CBZFGkNnuyfjSszQOqd5gtjt4/XtpCh1B1txCV37RmgXc/MajbikG
q9wq34GfR/eYLHtvuvxR/BhXhNsH78zF5+UKRDQ8UsODpmXyAYSNklYp5LyO8Qwb
FLo1evUG25WwKPNLLHM83Amdj9Qk7xZQkDs4ONZ3HBb4xO2Avfxim3J1SAz2vnN0
8vDak8ySPXdZBdnyJHGD7tYw87XVZDWM6qHv7SZ/Xu+0fB3st0tDsz5uLg4h8mWs
1CT1b2dzf+aVkbKVO4Cfr4bLvsAR+9LwwVDyzaHy4gJAOzkD4Ma/XSH73LO+W54o
JcSfYm1/131tHmZ8353e3Oew8UvADaT7Fw6dUORxYe1cLk+3gGUHYtIe7WSbqD2o
9IRSeUMqPuf5dspQXz8m5iOFJaNnV/aAQqQmLwVuiVE2QEjT9NLbksx8y1+/JS6s
8rvPvH+2UrMh7swfpNm6rLmCSr9Sw2Z63whvJ/7wcBL2S4z91HG/19mam3UDfUcV
QIXcogxJ+1oVIlhNMwE6+iCuXA6DXoS/YtV/wlImXT8VfwjezqMjw8brM0bgoFAr
rbtDYMd/ki4F41vxBDhZe2iBJrkTPKZ3cJdv0VWnXODp/o+uxkg/ew4tGR0JKEv1
Qn0aUIhKgDiLxGdseId+6KXNWlnLZvr2hkoAV6ol/aD4tKe2eynloQlAOpJwVnth
fVs4goHZp3fMSkDn8dw/4aCIXc6ysmTVCHJAJxPAM7ZZhsO62HLJH23wEPAUq95X
SEJoWgSEyOyB4poYtKNdbelx1Bd1MSyskjDieKRJBOXNhUU6xd792xmRPPg6HBWZ
GrdQRY+1ARNzPoKTXMtUaR6PnamS0hLZNBBsHHh9H75BEFpSjXmwRcO2zvP2rLJU
wLBhWdU//uVq/FtZqaSRH6ku0Z0b98MPH4uOUdGe5xNhmtUBkngCwShHGQFw4NwC
qHsGFW2QG7diikhjBKpMV8hQ9Y/FS3WZlvjS8VhU/hO6LlENHgkhWLuO6gxDKKrf
An05kn/jx+ZM7XgJ2087+2dHtKkki+hglPqxSVpf2vMiMr2uNvEQI+tP3Bv74h2N
QQjPOOqrXp4z1PbnHaV4yhzKPdniytxgUH4S0oNVS4gBmlWYIrFXtK7DZhPEPWA4
MMRyFqptBJW6xmPKhMheaUoHTe73+G1j0J2y4Wl8vTBnlCsFJ1xiER21JMkuMhoL
+0n0BoUt3c0fkzrc0RFUGOfikzvtsSSL0ED8PQsIF00sETH5/ktxGUCLCtbkcsOC
xCmUqarqQf5I78t4bK23NQCipe8VkE5I5jDOHGHPOlUAoNzYiZ6bGjLKVbmrMHpj
y+/s3+uEJRS5NlpcfMBwDfTt5w2U2XG+DKmyzqofJS0fodAq8fb8a2ChigF4VLdm
vTYGIuDQjugfHYoH2LYFcQRAS+ZqQx23fcV7uNScP8/B3wNmEWE8sSNvkgywXFUW
57amci0Wa/Yx5baMuxG2SPZ/+ZV3cX54N/5t43RvkiElob2OqB85AUcT+meqlQ9S
L40NHdcwoBB9iemBieloJsFRJyyfJhoROHdS48b1i5Y4t7JGHfWZubPxquRj6bmE
lwpXpJDpBvng+zW7LzjUHXArswCSrXyLm/44S1Y/0qZLIe6q91AR+0kMkW9LlzUg
Iey99lil12fO83+5hSr6reZ+ZziFuDhF4zDdV5zijKX9Pw8HKnwxSD7UHZ+9Mioo
D/LT+MyRkZ9wJWaaMvM5EuiFNkg0EfumkuuXnVMI83z65uYoiJMHChl2GqLWj19P
bL29QIIZACLvYY2RWcjcsmoaIVrEuvtCF+8QeBy+cwRPVb/9W04Es5qhIb+ekNmd
qyZYuj1vEyPfprmdJK5G/oCtGKPGCtd1AX9TAm9jlW+g3ClpNp9eApIAtTvHgFra
Hsg4/FHpz7z6XVKoXa9mMlA002S0G+hgIl2INlITF0hp+DoG45bzb/8CSLeGyfo7
4OQUHE19/wXKdkKL8YBUPqlFpQp8B4Otoau4RisFMKD8XI4gYuWgS7bK7vmiQcxX
xWDxqURuVZAk+p0OTD+aW0hbm4SlzQ75dSgmywQaMr0kDR/Hd12P3qCqWPypzQHV
QNpMoofqLPDd8mUKVQJtWU4zMLfeqmVnl6UYc5XBYks/3J4ObYARJ6vteyvro8QO
PLBw3Pt3cKlk5o5DiTiyH168UKa6NbTYHgXYr4GaA9jPrbLZT5H3ydZe1q4DQAGD
ueEfbtIg9FT0OzEesgX2gICRopQootIpX1HwFRZVWYgmjqYxnHtoMMPKwXGWsmj6
fhBeisBCoTphHTUp7DlN25Kiz1K0/PnGIgLA7+aX+up5g1OJKXKTZObkMbNOnK/J
P7JguZNTf0u7TeI3eImMPaL6zvN5x/4nX/bOvLgy3gPCkKLhiOWzKLhEReZjNbK9
UnYaDZnmuQXqKWZPi9edwhbzm2GknnmozWAJMtRA7RdFALzg8bKyCrLOqH9RUwP0
2GGLElWg5/cbFEhlzTuxXuEVxNuatC3oXK4W2JQn1e0lNp/6UzRNp7r173ShuL+N
Z1TcRU1SLqYiA7NSO6X9BRSuLNfzxFxZ6ZMSlPMUJ85RLlGk7ZG/FeFFRGZk3OVs
CmwiPm9PqnqzcaXLrCEO2XEg8MeX7VkRFNcW9nPjz2nuf6ah4DICHbduh/iRadhc
qAoygcaDxxJMgfVSOqkwUf22/kdCJYHx0mzXj42P/GmdIo5pGchwbssTRWKGH/Pm
qQIfrlLN5epSS55xG6QcoLU1BC0yHY2+zDo/L+NRkP/JELxNb9LCAaYRXXoYTLCf
x3owHA1COcU8hmSFJBbDsPAVvqEMTQsO5fhMZktE3JRjn19UJFXvLsCwkltG7a/p
Tn0BilIZRJTku3wYBtIOwbbGSvWR7cYCm5lyKFIzP9+pKO9D/gVwnxH6FqzcBOxX
RrMSUHSGD6knZaZ08QmMNg4+IJkPQ512BS8N/ZeDL7wEAmykAl3z3puvRFRRonDl
DwlAywm020GPIEcGMmY1vG7kGcWSJRMpn7u6qClTIWiUsO403OlmVRPJaTOGc+Gq
Gsr63qvZmUgzd7zaVVVWGRL6T20uPnDmK4Q+nEIrrGU1l05US08Mk1PEH0AL2SPD
Dl0yYdabl6NvpHMrZe+bRJ2FVFLDq7FAhmCaIf3Q0SA787efqK79DJzSS5nfid7A
xofo26V/OzbCXklSPGSWcu5KJ3zwikQnHbGUoAqQKMCjEcihWtarpvmuZydBDyDj
mVgb4JK4rsTXvunZ+nO8Qh1Pegj0j7mEwdwVOGpNNSHw+q9ycCIaelnE+nXy6PpB
NXmff3VFI/BNNIvDRc7jHQ0/cXHzeQ9LPo0KPS3yzIA/HgzrZHqb+NQCZs+uzoVH
naBDyN4/N6QJpgvPFcIRSpA/xhU9cB2hwt4sxBK3HTwwxEzzk+BFE/mJ9+OKHCE2
wpMn7McBejcbmtpIuFoq6TFX/K+yU6swUoheXUfs19cAxfAb3fYoO7xazKPjwz/9
2iWgcjbqgM1CtIUgyFFsy/8K1xvFXRsrW6foHaBkKi5PLqhfWrsHnLqvhub79ASf
l+Z8Zzt0pA7SnkWmRmug7UMu/bwzriltyyv2EXEK123eBD01TtMCHfKcvh1hRbyb
+Xk3Og4eqFfTG95rxy9s/vZ8UbP/grV92noGRx7p2CIRrH6as5vjSn7nHOjUiXvY
baU9yS9ytx8SxSclgqsFzLzbiuhL0zsq7fMFX/PPIIoMsgBAu4DIA+RDjrBcYHAb
LHqK+UkRWKRakXQrydy5QIRhoKEB64tBLxVHCjFe0uUaEVuMXTYNbTj2sapAOYRz
66+5TlCwdV7SfiEgQyjwak5Q/wrx5du1XwSICziFFH8lxRxfy86zjd3cUQocnSg6
2wMZ4kyV8IDgq6d/IzbZ9K9pK4zNRC6VX+QX4xOlziDEVjKKAkLzAFy73NfnCOIz
9kJ8ppUdXS4049Cp+7EU/eA1lNPLsj6bbwJh9Hs78P5CVlpgb8HRMF+HdyzmqRWT
tQdr6eDrDV792cYE3kLoMQYHh7cL/PQtTHlTDnUABTKcm7gpkocQDidUucSyUCsR
S6Y/brh6JollQVEB/kSOf58NEYFAIIKts5cMnraX6k+yX5k68rKpj1E3/hCOxsF3
FUJ6gfApH9NxSNWx0BmEayqE60cWZpHcvZWSgUFJ5qT+W/2pYgmCijt0jDJ1jkVY
hFZgJ7oqN7qoRAg7hOPDZoeASadNetQNtIqEXyfMlY1skmJIRmkpqmZzlWWMA3Vj
8nd8UAtX27AvRaFE0cQbxUneTsq6/Jkmm/5sVmWub4ei0SEW+LZcQPwbWksTDuw3
2edpYGiTcoqloiK6ftHrRXviQzDC3h8qwcv1U7YNDoycFZXD+Wz++td2MhxP+Ywa
RmjXAB+4Xmi5kiKCqm5i7tNAa7oj7ASt1cxBRpzVFCrP6z3uqZd7bDivFoSTdeTm
bWtLifJ20gf9Ax6GK7tWnbbTJfUoJXRH9UNGtP8pINezZ13SIR7zcw2KSnKm5abn
rlGXHQMJXRniwlkSRwoz59oug9sLk84/Yux9ytSGc9O5JHwqmviXLLtWReF/dpRf
qhjGxJENOFmbvmCjcyjzREAuS2DOm5JkvGPyuXpfo2L0oxoOxBcKDpBBYvCxdPFp
jv1JxoETEWowkjz9/fQ3UV4M7RAP+XpUhThCLr45pRYgY7mJbwmsdBqmZaOpJFf4
ERfKIUwpRJOjHxut/OeAErtDkKysqvSo3Ra/cj95N+YY3ur8RUPmhd6uI6Ebc7Lc
yz3dakIfGJSE8JabAOb2LIgMeDtEhJ+xArOGpCq3T/FfHrgmkFpww7nL4WxxFns+
usHy70lI03oZ9Rp0nBWXI9qJdAjoqXNkkGo3lT1Uv2xyPM7dQAR/JQ3hJNmUtFgT
GD4eRO3jAFhT9+tonIeZMDVb8YvCF+s192Z1RQ70kEFDe2B0M3KPcTCf4nlzaODa
lgPPerKXxRdz1stdbCfwXWEguyHeaRlCEDreVzs/R08vAQHEQXstBbdY752HG+MG
u1JSVhGi+8kYakbYydqUbRLptZDnkY3Ca/6jbA5/KfYLQI/xY9JsfVC+T9f4FNzy
rv7w8g6mmu/tZyo7Rivb4ifD9NuhnKfsh3xNtkvhVrKY1+Hlkej8jm4694bP9Fpw
dSSKBTA+Qyhvw1YcKk15qjySC/gEAaf5pinlQOuGqOqxYjWK75OLSwK8lnq/HLha
6yC9qi2OluVzoNZV3uUbSsQeDMWxzvP48GZQbs0Dfi1PczKInQonQIXHlC473OoH
Lt/641Lb+yu8wWF2+kUXiIDDugusVL82nZLMJjtg25gj/Z+azz7Mi1Z64CBljHF5
LHk9ae+WlCy5jpm9a5PJXXjWJzUls3AalpZIY8ICElQVtuSwh8x7bt0Yg4mKCRLR
YQ1/Y8ANfn6xYN2NtgwIYBOWBA+ViUIL4lvK2zQwUXsTcPeirJp9ElVkL0MgKSg5
7M1QVCHsjIX8d62QkD7KLhPVcOrwhka5ZahuLkWEIC6+ieB5e8sKVLL2yNtM4dIG
g5xukgHF4QdrUsxYTuMpKB7la82IxcLTkf6Apz7FimqrVRjwlTQgddKFkqas5Ets
14hDzIifavrzeu4tv/1bgW5AJ+VdZ/o3JRCcx4nJYzRcl5uR3MbdhC6qzHxC+7sG
wd8T/csh1cXkQL3xpN3RjwcnmrxLgEp0TFEcYeyt1Fsihv4jQ2zQkllJ+AZUYAMG
Ctrq4X7MwAYotCEedhpa1uz/M0WR8bu7AFs24yFGtqxl+tAX6Sjj1DepkWAhJpwc
SCSEr66uJ12+F+isQeJsNI/U29DHtNUz2gM2H6cWrtDHRJWWtHZs3uhR/JdndrGD
fg4g8d6F5xPdDs7+zzOpSbwtOBVwCjU/LT49c8VqbEzxd/wi97zQNMrhdZDKy5EO
HliYXY8CyNC3oDOAntgG0pGLxLST3FYSDS+peVsYtHKr5s2ClycSnTXSrcb7mE6G
r3X418bhKFewNy5N9ZgjfJ6RFWDHKwUjtXpmojt2d5U/zQGaqigTJubsEUerMIip
XexktvsW87/hBrnmr9n5S5e1acxxXsmU5NFbRXmQ80eiF6tx93ngR1O6pPpT+ufu
yqN2Qf4B8/4Jx4e+iokzYaMm9EmRaQVjCh9cjzBl5gChC5vmhbQlVoSXUw6w9GQI
CrPP1965RIkV9vh2rpptWij7F1Xm/RbAzbP5JdcH81I7tJkUEqm9McKgatq+ehcM
MAmRirs9KYzszSo/MbF9PPH1IoK77Wij+11q/DhR48F+sWUgbQ0qoUSarINCPsV+
WMBTepLRiOhgZfHBVnu2TWFKz2SPIJPEA3XFyJd73uhIPxFNwoa/YDOr4GXqJ1ne
f6YLe/zlmeu70PwwSaOw2ER2SZTDqpzilAAtJbggw4+cg9ZUvbSWicdJJxDqxf2U
4Md+P+p2A6BAaNhs6AXz0ki5Ntg0+PxaegjMkJ36rIx9McYpjc64eum35gvHqBOd
bVANPdGryzkdbvYf96Bu5bZJ5aklZNB2ESDkNUR3BHOKUSgNtJ3OnwjRII7fXIvJ
P46CXyxYdlIj5qpF2xMcCKcN25Rehy8M8s+zY4FscRTlrxAVcL5r4HtJC2F1+olH
w8md/jG53KprBdX++x9BTIARJv2hE1IRBUBrVCWCBxtZAQKGa/mhjie0hwUZSvBG
rcteaL6k0fqU+Zhv3qTtkxqSH9uq7BWs30cKdxJAYZxCrhspy34fUJoUgV/EoRSZ
Dtphvj9uGHdiBegoeDaZE3o3s3+WHzZb40HJ7N017gDQIDKMuukpQ7JN81jGbyjX
XBL5UE1fEpkqX4xnSoya2l1JyrbmymoZ4uOCo3enEEb569TTD/j/4WZmuKO93UYN
dD/C+nyjC2Zrn5Qwi6Mp3Z1ZSajXk7oeoYZdEMrk8r6bUQRABuephJaADsldIiBP
D/Cr8mX5OFmtmr6Jr4WkvhxQc5QP28rEVXWV6BSkFGTtEKoSQzV8vHf8WEi/ELh5
1YOZgsDaEZZM5Ub3JFUW5CDxph5nAE5pB//ELxENka7XsEWQw5tuSKrAqOTuCvp1
TtmFpeNrCFrCL5ydGOn6JmWayJzrsbpKLcFKoIChEtS1aOb3GBR09AmcUW8zpxcL
Wwx2Dzj2f0bmevi2b2LZQW0Pcb8/Q6WzOS4Hd6vZThix2+eL7ZJBMGyCNVzlc3Tj
p+F1d1QyZCK/ezurBYYY+j7hMGxIdfUaxaK8RMO+1e3JSf0cOaifbW4Mr+JmA6QF
M7Q1Qb3EU7IbbCmC6YWRQU28gIfMaIpzlqm5DUCNHnS9KahsYfCBcSNZb6gregn2
LQYRkPuPBpdQm3WWQ5p9ro5nl7CkuPVJy7B1FuUZrCMd2fd9+IiKthIQLfKh29E5
YMAusI36/+0h/j37YtbZdpTpATYhtEAi6JdTszZRbQu8SqZY4ZB9k2XBbGUTN/V2
pz771N7mbOVBsGLvft10P2WBoTctRoMfBaIUozqWMhjKhdv/WStkb4dUO+OkHGBu
G/d/Ng3Ke2CACzEYr0TIQO9eVsxz2SUSqIF17GRZfjiJkN9DV+op/6TAAKGEvfzV
72WBEn50svuNSFXl1hzCL02hVqBytZtfx7lHlYdDnpg/JUTn5RwvoYhwoYDhZ4MA
LyqdPAmRlUMF0xJnO5kFoPrRQbqrKk7gf3a9xYS75dIIdyLSe5m46d+TaPl3vNlp
DZ3CREgVnD/z+CFKWKBBsZA6dtVx6cL5f+NTbihiZzQ2VyGAvGngYmZY+1o7cG7y
P4wIr23NuV2MsfpwE8T3MC8sBPI5ebswhaw/G/3yVJ+pO8kuWiMqZg1BAMpU2HrG
ZteUkOK4TPW4gV+UfLO/CihGRYpNd+9CES+n7FxTY0uZ3h8wyDsiecJojajTI+yR
Vj3uK6XFPCp53jQHPwessu+wo1g53p9DUllz2T6CximqcR5rZntIUPQ7zf6iOKVY
LYp2Q24GAgm3KZkYW+J8cySAMctRgBEl/O8TUAPJkDWLvxtfDlyjBaOdbctzgT25
qqaOL3A4+VCvQu1SfOshLry+2a5aYaH1G1/mwQC7FR2qiPWQiNh9JSu1kwVgujjR
oY/Gbwm/Ost+DfMdihTKJ8R59CDNKENJdXP5fNQk6q/sZUb5/H/7K8ZnRRt3UkK8
zr/QpxXmPfURXelf1EdWW1KqanzrV7IKJVRNo9esd9iEEnmeqs/Rk0NfjtPhnU+I
NwbMc7X+JQGzUmg8Jf94tcCiNS1/9FXwI0aY6M9VoWsOxcl8uVCTjS3HIIT7vg/I
K0yVADxke3bLT33mKjVuJUhynXbtoAVt8Od9ogsdB0ZOSw9XwtnZrsRUhyPrpPUL
0uIdT1x5yeG1tkWhkc7DOBIczX/jbVZa37UzHPM4YVOs2IgngBtQcWATPB0+RWRE
SnFFZSoo7NawokcsIkfIGGdvDFhOu84ogx2tztcUsd+PoPINui7tEAr4IwuxDKJi
fatTWhH0r0epFQH7gwca6W1FocoxIXj5cx8RsRszPRKTa7OS5P6xGmuSfVhELEzY
LCppOri8ks7rEueJjw+poX2qkoGuSawrNZtMRSCT0Ho62UnLkkbgmjoU1CVQn9q/
2nO9s9ZoxdM7vymHyv1Ggu+X1mwNGO+NUHfMJ9B+0iuRFJ1X5Gnm9HFiYrZIfxOt
+gYiSLb/HPZi0395h476vBo1CrM2S/58JFmN8GPeKfvyklAKECP9+Dw26yLgP94o
tgG53NvpZNWoygb1xpbZJNeMYVdZfrds6ICDHD+B+2J3/inJpn6jOwUuJq8eALSY
nJ1ZpteDRq8iq12EnLZSojsgWYj4QdmBjLQ1gcfNoit/YXXZf/j2gMecGubGwP+4
8UrfHE7VtfssEj4lOns6zD7yVV9BzBy96kjPKKHbBtYCYQQJ6IoLgIJLUAsrfsor
jjFT3VG6K8Ey6QzOimqDkat4j/dO4y5NRlkSFsuk42yigFJLXOETlN1keNWD9Pqt
4gQmb7XqK8v5NGxqlic+Oen33uNMjqXyDBlufobgctvUE4IJhCj4pAuCKUyGMjoG
wRhasgw7HDofyjtvoP3ANAb8X8iGJn8dNKjgPellQzFSTgayTlH8m7UARmg+bOC4
2ZNc0a4ERcPIvEMdqcH2fbI0ykKK8hPmx2SO2IwJRqajwdStoUrXP/lsD0M3K4nG
tY0vNqpwuT8Gve6G4TYCIjrG1tBI/SUB2YHMSfUZOTf173On8IxQgdWd+7cGeGJa
lQEGjCzr0z1VskofZOLCHhFsTNiDutIUfPFE0izcDF1CwD6HaKT9BAqLjb2oxAiv
YuKw3tuTri6aZpsReUjpQSyxPrPiQLhJazhVL2v0oQY3rcxgLCDOmSV4DjrDxI1z
mDDjY//VsVyySAKvyabBQ41SXXsxLrwEY/n2PSKsFakRmRg3fRDPQ/saFIysGrtJ
2JZGfGNuhcCWmN+qmYr+sH5KdC0i9x1vjMUhGBSiz429tsBpW1MsI8PcqobcexES
YKl8sW+ZqOJVcGDIou6iTgr235/zOdRVoW3dXmXfHzTwrWPBGWjhAAx2J/HNR7ie
NPjt1bW0bPCEovbyM7GjH3VNd23rHKm57u1PQyXNY/0s/egjpIGT6jNuc61UZOrt
A4TKF5U9/o0ujLuhmehfjDlCYEftdVlxeQCHJTHPdklsu62b947mmQnqr1QlpsOA
W6KkXJtsBZQvOTeb5Jg49+/aRAyxVeIP7eD5/RsxdliprKGDGKVwuO7u85w5w4GL
D35noUP24k/6g9WlBtzQcrUeio/MLxHOzsBfrK04hfgOfYS7By1Uw4QgW8eJWMnf
78ytSTJinfuqswnmv23JjllaTKLstyT+csxh5eoMuiPI3B1A1N+t53+m0liH8m5S
gSG3/iz+Lm4smMOTrygBlSiFJRLAONaxMjDkylzSMjJLFGOyhCmw1Tzr29VNzJrL
CNsae4ZHc+J7bSw+RUxNuKSlLuzK1nkMXA1mX4VfPWQ+zXalD2Gc2C2K88RUCcv/
bGhCVl4ZC/a5D7bUMslibcZagdOXjk7ajfoYGKEazXal4eWRpSAHCi3MlbumHc5l
/+qWukMVxvzWlGrEAmc30C7fGThSPjQcH/OMw7h4S7rST6UbkusNprOkF8l1pnKQ
0hsvsaC3i/Od7+Q3mtFC4E+1fexjxrctO5Qycd5t1KgxEzkslLkN7PFU9iUyqBXK
uVJmweEQSdoDbPYXQFhwQTf5FyQm9gT8y+2QSKU4WLyoFTAuQZIxHcf64nAp7Xk6
JTsQ8FffjbI5/DlTyKqi0g9T9cE9jeEphnOCb32HzPrRCGJOAzp5o5VrAGdvGWVu
+0xrEjh51z1y/AvmPHKEGwnOSEoR1mknWBh+foO9YhQ2RucgXBSHsodus3xGCOk0
pz3U023WVi/tmtt2hfShGI7TAD0Fz0Jap+wNEcZv+oYmuXgn1yKHDjOf5meFSfKF
fumXv475CnLyuascAquU5T23sRpIu5ZgNl+fsQXN7wfWeNVl2ZWCx+BRTnAUzbOP
UbJg+uKobpK8lmTf/IjqfVdQvXMqfNndXXZwP9clg50ie4V8AxfGda4iEQdoNgNl
2seK+th20Fslt7nn6o/7qY2pIFIOvBuJfSPpRejQD0tPzh6WfQHXjiyoWnOEc17S
fdBn0Fou5mLANALoaBoTeGcLfzI//etQrfBKgW7hkYB4vRssBmhJXiRvPTI0Aoxx
YQjj/jUt4k0lPzTigc5Cwq+bC4hRD6+/nMdkXYMchjxpPAA1/Q+Too20nprUtuiK
W16XE+ZhFJI9VK1zfM2YKP0qpTiM+3an1KUbY0lr67qxnlyq8y9Nj+tqTN4wLfM2
R2deuMdFI4BZJhawAkEdae7P/tbIrII/vxhlVcc7/XZLWXuYoInChBMKTI8jMid3
OHep8H7e/JzH5Y3rMaZ+s07jdnTympKUfdoyNh96JprI767FTopO/pL3obgtbnJi
7mEcCD2ahF3lVJIe0AgNTGLDfMpwFq7+r5WKFni4+FPWA8IM709QXiZv90UDqQgz
1rOZpwW2ko/+i5RrsYRJWtkPfLpZOXFQGsFYs6CbNMst4soPQqIz6UcSZ6hqKjlw
pIpNQNWzsEdNLOlrS7g/U7h6dPvOboEudsmwqlTjH+MhF7lmz/ynKeAUiaFFoQsS
z5eO7GGjUsp4IMPF/v0W54P1MGH5T7N3ppDoj8pD5AThVMokiqcJnJFYuv3ci7fp
/BcH16ebd/qLf4co8ZRV3fz7Z6ZzkZbZRrgDNVitMdUchPOJ5I94c8DS5n/yTWAH
LI3lXuTd1LYtNgUFyiLEvLmmH7pCIizteJPqfHUvJAb8UJSSITEUU4iWVh7o5Brx
2gM1VGao3sc2k34gCExpTqfnYUlB1Og8CrUya4gGogv3OSv+dUlLEp8tBnuEbtUO
KuahYIxZd1gnH9zQanFkgmy7r7EhqFnP/Dtg8LM5Q+BZ3q1IKBJmD5AJpI6vssvT
Vv5jMkjwKGghtB4/98ntpwgpJHHGQrwxoHLvGUjSM7H323V38UPhqlZhNbuoBL6t
SvB95NLGs/9RNJmIaqc2FMtL2z1LOW5l/B/RxJDwFiDDntc5DZnBSWNraNgd9Evd
9ChDuGZXVMFc7lTJQb7jVAhFgiOHPw2c2m15L3wGi9eO/+1hEAn3g1ni2IC4m6Mn
B2EGmGNuHkGbrfnQrV5G7sYflzhelucPXExGX1i9cZOmK4PylK+qPcTPfi6ujTjY
/JXyuYHPzIGZJOAHAsAT4j7P4TAf3g4pBEZYbi/14S1Rto7Fb0p9AQ9cPcmSa7n7
K8jgMQhaO3sn+zGiUFDGeVHY7r0iN5slFB9lODbwCc845KfgjAqx2+GIDPETzjG2
uklH8O6JYOLpMtPYUgZF8mxPczqvCVLZtNNhxexVuPQNsZSncth21K9YRROGxmY7
90I02zsQoaRjgMyrMN9r8YGTHXSabp8lSYADmwvDUa+1SMfzcyRbomj/AYWw95Ab
bg8JEXvj5Qyg2lZF2EQ360iV3/Ko695FQnBkSxAq3hBntIHdHr9paDQ+zqvWA88w
FEYuj8g2y+jUaan0+YHyHlkMUuz51hiNEQJWc1MYwh+c79WKYUI5bvHzos0o91j3
2XVSJqdra/a/u6iE6No0bglPzyWfrQnl9mhwyJ+gSqlAEIHJ8aI1OcOdeFLMfYD6
eL/oxIXFREoSD36V1FQwiCs2Ae2gAQaeEIgbYzyQf+yC7BxhGuV6ZbyJ8rLUCn5U
MKexU5R1ACt3A8s4DDdk29q/npMflWtsoEjuwnm+R9EUtRpCWlJeWLemkNX/+PjK
/31DE+cJBqI6HWS/f4adrMGuR22NaaCDjOROIyT0XVki1/dgBCUKWuo/oc6bRWHd
t/dnyJOgIiQGG8XDUZuj5ellAx63RX97wxjbEC8Sya+h1G3hmvfl4NHivGISRRQ8
i+E8oEFrXOBRQIHeljE57vIdPem7fOLtjedCupqMikyKpVHiKggPgL7oCbShx8cp
HgR1MTGoDyRXg79k64KJtvws0n50cpHqId0eXBLFOH2n3wYO18Nm3TaHUyJ26su1
nua7Fw81l31B3u5+qqz2We2sSD3VmubmsIug/8KUSkzsezpT6PjyAPQMiPZUqbc3
UxQsJcB6v81Iafd4G3FXSx8E4gLMVCQBOm7cclZ7N+fFLmDDRcupWxaGvBwRpzCh
9p5TkMvvscwXEV5yL4WS0wkw66bEE2irgVqkRaoxRkKrC6NP6QlRBHbGBc+pERY4
sYgXTCLf9APRVv3XMaUFYp7UI5aV79fmBMypTz6aamYl9Ev+wCk4CURJgYkWdK/k
eQJkIHNlH4+bNixHrwlwyimx0hv5vRmFATbyntDQVB0Y51FvF9rOWRha648x/g5S
Sr6X6fMrRmwUuRNZKpsSt3t2uKK3zICZ5IqvxG+EwXrqI9dIihMyu46KUpC5s6Ed
qc5E+7gGR0NsMakMWIidz9pZHYO/gXAj1t34i8LxYhMhJj0ZwGeGoTOhZBKNh/Sb
oleIhhBTuP5Mdh549XCReN8ruu0KRfvsJlxJmSB4JSouIY0Q81b+ge4xroVFoZas
9lC+V44NGFeFI5sKuF90s3HlqV2Id69VgvbY2IEVyaF+QG5bVm5pB/WbREqlXVxh
nkrw6SCqYHxtyEe+82lVMePiEgkhsnRUZPsKgXQE3fTvffXMZBOF7VZ6+l7dQJck
2Sav26R5lDMD2skDGS8CfkSUyoPR2iLNSboLNaLKJgB6XgF/z26NUiI9kCJfkPLa
rCBMvk7BjinOs3wQpp8ikh1A5xJm5Kt3ymoMtOkEyW2fFD5YkzeYwgd8wVzp5C7T
hVFRHviIaUhRtQw8tt+le1VPmj5LmR7TaI8K8ihwR6MxYAA23X0Wva6JliA6Pq0J
gVzqckw2cOWIaziKVMymvNFVG+bj1bgQ5cdhZ8spUav635trxz4byrYrANTeTxWE
I8JqXDHZq1CzB84rqv0atWGIdWc9asfsoz0CvRntZNmdoCY6bNhvzmsqLiGrAVi7
6tGKw5ZyGnF7hAwJQVw4bne9DElbln5Z3YNKxsyaq5Fwn3uOixlo8oLm/Gw48h6O
etRr69JdGdbiNmBH8ydRNw9u5hHybhUVHkOsJNUjhDemq3qG9UkhFF7Q95LhrRI1
5hAXszaW5VMfSuzHdQ+NvVusAgAnPyRF3i8UOSdsQO1n4B2mrDtlQ7FJc9ZpgyrV
y73s4WvvWxi3P1NmsJ+1FHvJUKFaQ4389t718ioATpkmCnh6LpjQRCTOAI4drRlq
zH1VHWBFYHDIG78xnQjHg6+3Hn3ypaL5FK7tV1+iN2IoLuW9suBO6PUllwLqsAsz
n022TLTVTDQU/D1bAs9TeD3hSCSxAnaez1VJ07hvHqk9E1RfA1k2wa4wBvDWwb3v
RoQgIxulRT7CIYx9QqkX5R+itBo6fBoHcn2kjzFUVboR3TgHwYNkCZ/CfH5u3edN
/niUVNPFVcZ1q+uC5gMrAwzMUP7wAExl3Y+vG7UjjUufqhjRWcACWnHbb9loWq7+
Y5LeyQaFns2mOSixbjvrt+9rFJVolFIjbo9iaWR4vgHR7whypkWZdnjp0aeUzFwO
AaTkTxy5C8mbr0Qfg8Zzncv9XRv8DBxZdDhyLu0f/2bY458s5wgINocjCJLurYet
MN+uW9gSK9WSPCfoEW2JkbOd5YWI9oljFd/M9yi6FveXD+uKUPH/NSIhhEt67Q29
PNAlRzxYLJJw6uW7n1/0l9ceCXiBXUew8ihWPPrdiapoXihFcwgYlREAIDkpxpOO
cdI9MVkLFm6CJdcjWIUzoBVzgh97bIcER+BzQ79M68a3U16P+pV491e6xWFdZj0d
AP1626N5izPz0ZmszP/NM0KiiZV6BZwlKeIUiM1gVJGnU6FRlulWNOyFbTe435A1
kPEHhwSnrWqyGtkdkSpS0YQIfgoECtGfQcj1M9tkFO/d5PpcjIIweY0mXFtk3Uxg
w2vXfWvMMcpEYM9d08XKcRpnrU9I2qTGb2CpnRfeSdF8u11cxD0RTXbszsp/hR+B
ag15bqB94TgOLNceyAEzCAXn2YgOjMbHkIiaIKM8DKCbgEz5WRj9/UsUult68cgS
bMRh0FfGIYtCYx2gxKIV2MfzHmOyIQlKP+7bmlgIKhW3w2XzSCn899tB/H2yTO3E
Vc4OrPbYwIjgmXORKETNyw7ayfpUj1HDqkEjrML8oAYvSHA7YaHhDhIHC1GvLwrG
HV9m/B1zoVt/6QT3S89J3b1o1xpXqFbJgW4Xn6sGpd1G8jW+0VUT2hPv8PUr5Qxy
6rsdelTPvsMs7OaL+ock5SzZt8G6qmihba1pc6yeoWlyVcoMF3PEmeo7sdx+ErTZ
zHYAtXTsBmnLXi4Fa2aKG0pFBgcll53Q8sbHYuqE8jsYqveKF7B2yWawIeS9n8ez
WxJf79lhS2AFZH9RsH3B3noDXkxXYrQ5I4n6X1V6QdocE4K5XGTBXo8mdM7BBHkX
Ke971h0nC6jM7hxMn29hJufsIsNu7GoZP2eB7+bYRJC4mMuNfQf1aYnCXrkG5yQX
Z6boIT+d/K+M8JqkMck7hnbAKCnAQmRkJRS0YFWrJ2DQxcGWZcknW4gCJdyJqc/z
YrzLyQuQ9HkiC0seILweny1mIvDt1qlEazDxvq6p5Q4yLZmkBSC3P4SRVF30GR9Z
qGhU3zZTlF3vWF+zN+VSb7tUxd1ZT9rHOVD+RHWd8LOIh7WQWGrz9EkDzrAHHria
WOGuz4RGrP/prHIHHhUpcWRcDt+r5xQ/SyfrwlTpmPX4958BWB1sIqe0qHPZi/zd
WwB6Cka5IcM5Al+NVeK3rQ9RdGoYDMIwgxJSCAYk4cb5lufRpsV5AS6k5s/8Jo0o
mGS0R7LnN+OH5Yi7xUCpkbnzxOllwBKjm1e7NtotHhsZ439du9T1sOsPl4uYuzIx
2XHCXpo4dG33Q2VoQUbZpYu0o10Qr+QcYm/FXSq7UyIYuTNCqg2Odfg1rHedlAi+
QOSorhuqY8ftXp5+9LJVtD838yo9QgKgvqM1sasBmZ3jZmcz5T3kQWM5Nzp4nvns
vAAUfHFwSCFeRUW3wqc1ONG6mQpnuQtK+SaMm9QZRIZUCa7/SGgwk4I6ITAO/yby
HpipoyZ9ZfbpmfGgE6miXQAFAJ2VkAscQh+3OJkPAbkVP3qk6ju02LinVQtNi6L7
bFP8o1hmpReEAQdb+lpPxTkRA5p4mpDbYO6LQs9fEEjMvRXRcrpgSCRO62vlUpeX
0lK/6MtO2YHFNwe+2ZI0M3Y6g5z5MEZvA2QuAhdOJGbklYl5EjgtrgyiHAjivrP7
INGaobNazkHn1oOX90EGAkzvb1sQy9cvbZWLDQvcrh16G7htHhDlvp/yDTQCBF2y
LQzGlcixp8ItOSXQ6pG9ZVOY+o/oU0YmxpGrtKrGLHxOODRD0nQig8OOstJSUg+S
IvgYNa+0S8/rNtt9t33A1MXf+4fjQIGB6ykIO0MJHRFaKuvVJSr2K1kLeZc1MEAC
LO0LLuBD4mi0NxeU5h+0/pKG/qtUA2su9KquTnWYppvn53TF5aJcfLFV6v0BfFyw
pqb0w9qO06U0qyaBpwqhzyY+d8e0t5PGvzwcfjmSubQvK4Hoc8+hfA1RvmM6nNj7
BfTnT6RzBAJL8iw5AscSim2+pdNsVGiiO/ZxtoeApDa81uDXqXbQhvbVIh5ABm12
OAVi9uypG6l06TB1x8A4wvvvKHUtCTtNDWtYHrtkwYJYoub7DHhLP4z65/wYCQb+
wyw/f05+dqw1Vgn0Pvca+M/8pF/uWiJ1d3UqKUOFCGnkwb5eyy6vn7EPKjss3mMJ
ToKSM2m5D7QLZuTbXqXjvdzqJFrDvingfZ6xaFD6sRwHPtpssoIpRWPL/o3B6uGX
dWrkyTgQ9MTQrphHdVXfqtlzLYI9B5+YsLoT8FpjxYsq6KpumIx8yps4pNoAwhbG
ogOfLwYH3onVHD3CFJFZaeIQuaOPHx9oIYmtuH9zVNc9vsix3eFvrIs6MMD7w7vr
J9MmDya5RytaHkNX6zOlwC5/PAsIqU4GffSKIhWuQUuPcHgpPXRc2Nbr1X4XJH5O
M++uMHng7B1k3yI6wdlFuK4+TKaCzW/M2fxi0HcBF3djRR6e/KnZUEQCGduYQXOK
VMGVHlPJlwCOBMvwzl5v+qmUxy9TDFRVdbrxaQHHHWENxPD0zXzv65D/X2ZeyaMI
2iGrvpyiqTGIPXYlpyCdo+3u94C/pnddbC/E3LFydQ9G8gswbtd5jXVoOm1XEWpp
j8ulCHF/Nsp6YNGw+J3iDBkOVvc0dPmBB6fZpfuPiUzOr76ZGWP1fS0aky0l4oGi
1Rp9PwAW3qVmfkTNmQI9MnI5TGq9EJE7vdEk7g42CxVWj3bLRJr56aWGEV1ZBgHY
6yNu9hCWRPHlaEo4jIvX01mEgrrmhAMxDp0zPlGRohlqqdbNFpnQlCpWmyB7lwIF
7XhNaBwX9kIS21oTalp6dnCm3Sqv3ArsgJDIlUJATMM2x3kOYGaJ+jrQMvuLQzDH
weoW0FZxjt2Lv/onoOI9cM5woGD5Xo30N0enuSc0RMLNvIlSHl7O+PXN6IAprlR+
pUsMqz+NBaf1/POP/xWL/q2cBZsih+OG67JAIpi1xdbEacVoHnVX/yM0l+KolaB4
TNDjrcT+8QdDEr6ZXwcXaIlbH197qldoW+e9WGLKiEOl3GdEzxkqAr1HtrRf87rt
2hWHpjvAf2Pvj4V455gRw5RQMYK1YwCGCmKOH0OrnjAvL3nAumjfR9bS+zztOd0+
LcBOJaU7EWmPDiUuwpo8QC/gAXGMImGyd7NavpXE5QAsJ5QcV4fr1wNt/GGhVMmD
cZB++MS0Mgml/mLDi6IcFe7f1cYR8en9ASi5c4aVkTp13EowT8HBHqaFkpfBMrmP
E3g9dDrTMVHquyKWvgxvuNCc/G/Flja1vErIP5ch60pQalbce3GVe9foVzCfE9Uc
GpAjqQC8a0NxV8YdYEg/94Op/f3u8vyNuG0PWvsbDfk3u7FEZoZKCGTp1QwvecjG
PmsG2HEhOb313JQ5kd47IBuQLxISgR/TL4FbcecTuqGL43iJSJC9PQSkj/lS8sBP
bsSb0wOJ1JCSZJqDDz7tj7Ijl+v27mjJMP9Q4B9A/PlNpt9gREExgSiUeCgBLkd6
lIHJmvnFF+24TALATlQwh2749RCBsfw1FvtSK080cXBXjJEi7bNzeh3S6n/QRb7l
00h+LQ0GLd6Q4ZJfg1dpqJQ66j2fPo36xDVozkCwjQzafD9Ye75WovPHpMpEQoLc
SnR+GfgeWxTUbOZXAFW4vozjfQSH6h+r9vFcACW46dRfZIcb1QTc3W4PT45CL/UI
s4QZ0zXqLh0rJtKigm4nJSLf/pZtU21mloJCfE6AsOP2go2wiAjPTgm6+e9zPHNw
xcG7OsX+k9RowP8dlohtY2MKzfrORfb6/ELQAPBSwSd9MdvWzUfsqvAYvSS7X/4v
Ac8Kha4ydAV+GbW+wXhjpCK2XZgQRibq3qAJ/Rkv8x92+s/Qw9pRTEOhzsCAm3Tz
V99qheMIAs+dh3mGY0tqDTs9G2OJe4lWdNly+K6ku0KMe1UVYSXqLGXc34+q80+X
QmZ11fLiaCFgNfdHQlt4TRR2N9BbEoA6aWlUrZRlIfCbVRd+Q3PprwDqfx+LdOWd
AwoPMI2VyGnyyvY4Q4VO4AASh5SHVTe6zThcdg9AghI+AQFNjcMqVILI99nM1NGS
0UYlPn6o+HRQwHlnjM9wBiwcbD/k9rqThQn7yMlUnB1rZv5tJJNqvOpoZdfL9Lut
k3eos29cQXaZ80474H05bmaGsqdjG4De3QCOa6GfBPd9pcQeIwi3g489Gc1avOLy
Yx1o4RVAMmyhYfZ4aQpMY9NAc+HrbWcuQ20V8vSAi7iwAP0DFcH7MFzVV0/TmoTC
lLuLTWtTs4l4FTemZhpwnlmIi4BkRMMxzOoVwz++eFd46w2rFWF3bOZI0n9vLIXZ
N3Ie4M/plzPtumXVjJe7gWDX0YqKKVclJ/vm9GQuvKkSM+Qlysck2BCdJUK/G4G3
cSsj5hY0OC4ic2FwNE0CHAHqVQ04m1Bnf86yLtQgr/LLtLY6LmwBnSwKDodhnAV0
fiG4+G4CV+MVOoauYxxWqefYhBeQP5Pn6CfFFP2ciBbrqkpjeg/3yTRrthtzydx9
3tPNJW/DFtigMHPwBx6lG8Hb0IGVc+S7zGcncdn112z6VEx2H+KMCnLPKiaMQE/R
N3ECw8/eQsTF13WRN1I6js9srkDBm+Em2NuGWgqvRkiLucuEhWTJIKDPErSgpcXi
NYo501weMjGkaKZKuv0JpgjAUDqKJmcQCndnnCQqhlmMLMFCr78uO+ZaBqGoe1Gw
5CSI18kldtVpmJLACLhh6oT0ogCYWtvevFiPa5pg1zTkwOm94Qe2AGTZ05blKK++
aun6/R5bHqbNTXEyvcc+MG9PlxMj5J891B8Sz4aEvoGm3MNXwnCOEKvZ+sgvQi7X
aR/wKCOkyjCESJIa+LO8P4bQay4UCMkkpIiXmPF/uxLoFzMTimRBRI6Tbeg5EPJg
0IDtmP79hIazeDURh2HsqXaX6RlIs9BQfDo1kDMUQB5VMKcEvc/eeAYuvKafhxk3
vEY7BjWoxgOBaFP3laRDexj+dRgE2gOi+QAFE0dEkjx2gJ2NF2vTJq6j8Mw+RtB9
TYH+7TFpZuDiFOX3DsD7DZTZbyVeijR4C+uQh/jYOCdmhc1EsL4tYmyyWn51glSP
zKfbFYf0R2PwZyIWf4v/hz276auNCTNBzB8zwZFrhkzni8SWWMgebDoibf/ETtMw
blzMcxZ9q004Q2tuGJd6fjDA0PA5Q2QVwL0dTfMvmj2whz646mMpCpX4kzpAYViH
cZI+os0bvd+sD4mLZRVH8Zf4dVp9J/4e3/BpB7kKs9mMSCj0RnddjR0+wXzFU6TD
TXIdvc/L4mAi3eh/FmYERE54MRI57+3CPZCn+BDh/8zXv5oGKlPfKGkGEscl4qLe
z5jiYt0Cd7g5VGxSMVX/Dxz1h1sVE165Xee3B62kAQGNbGUuXBiKDNQFIK0eggLZ
H6X+CyvCt7Q4ow83kh2pKocHuhYEFk75dV5/lERyDFrfJdD6F/fMZY6d9ZPlvzU0
pvYXqRyvGz20ae4vpTZ89221zI4RBwbcWrhZ6Srj7bcviukxTsEr+keabQoGknxk
Eaqlsd9RuQpraN7MIj9inBEJ4FrBjeraCgekC768ZiXKBXzUDmHu43EMpr0+l4AC
4cfAt/fcsL5Dz9IDKy4VKQjPByHlWCLIU3SktoU17WUUOLlGKhEo4OI+8Ha6Zv25
Cj47MLjsrC+crJkie7+j4oyAll/08Y7LTKUFOvX5Gc43MtNHn5cFEshgloZkepQR
VQGPqMK7YMsntotO8vRqruBoDI1xxwFrS+vJCWCPBnXaFEJZX/tpoOuPiBHT6RHj
gO7/OU3S8csq0HPmXaWfmWtnCXkSo3F5SNdd4j2eizBpiYYvxgwkSkA6X6hDs868
68+dMRJBIcUJtsypHxmWdFic+vFW5WHUj+l6HSoB2A0OD8Df9Tr3jDmQ+J00lCXd
JwDfYW8YyQhsmY1jsp6OjHuyPNzXw2v6zTC4dleM3vpPSUbOqpEZNtPbuW8p2kqN
2BrA8n6eqL2SclDn3XLuBp58DlmndOJkfQHLQsYc6UBmNQMssN2mEWPhVgbwW9Af
txB4pK7jSZllb2Dsam9UMpRLKIm2jco41Q0nSJF4Sldiwwmy9b8Hy+9SFTh86IS2
13EOtVx39NLzJ2Cc8hkgxLPQCrrpANWk6HKYjG9bG8UHO1/dKswjNK94qeXqp8By
01DmdkVEhyXUvzOAeVZxboVE+kY50AxnqeSiFTzNNt0v6LNetFxip9w/GN3l/HOz
iR/DcScRCLDuckMGs1JDGJeR0GUDKt6Xvc8X7n23zdhexF67/Ee9u888hNM8mnrm
txYAqugkKHsx8lFPysdUbiqrjD8fd1b23o6GtHIG5NCF1qYa5jwva6G5XWIKknom
8/YNhk6HpJxbxSI2G22YOp1/eS5Ilc1Q9+nEY8yLEtIoibI0gr6muOqPbHplDqPy
FrzaivoDWfSTJRE6degVrbnQ/T9W6GBWCkN+PkMk2MsLILmHVTxQce7WN5rWMQL9
BFi34H7/RGQ2QOqcrQlCYA4bxvtdtKhJs+7BHrYGyxQR9ulvq66r3f1XVV5+jO9x
2iM6BTD3HEzY4XOx4KMUT816c1GxJdDLr4Zz5sgtAbPB9Ymw01rEsccuweKvGO9Z
G20I4c7gJzeJMb306qs2/C61RNeJUa/oNSh2ogQojO5iNuyPO2TOGNMWWGtwC6fa
sBKJrfjxQRwVKBifeqCTZfk9KYq06uzbz7bBKODhW060f0Fb3da1qB8jG/d4zMTX
8q+lVF6C426Gu6xHTXkMIY9aDTxWZgTQMKpSerPHrR41C227e0w7btMU+bsWwCZq
IsKJ/YHNEaMmtD+jALEz7+8FmbOKKmkZafA2/BdZAHxnTIdCecjOZhAmXBP/PBBY
eVsRsmCaaLvnjJj/Qdo5K0Yur3p5G1X6PlDG/dFKr2vldu8ga15ZeDZpKKX2iGBB
o5RGClZMtD/4oN2/phcJSu8sT4cXnrYKXdl3uu/XRhDbzTD74AHjF4u4n2BeF3x9
iHg7SGKKHm+hsZJTVvw14yv/FchmRrXxHdpdy/N2ubH5J/GrQtDd7RHi9fKgyE1T
SWEw78yuDCcU7Jig5P7672d6TMwA0VetuSW2qsIrWybmIZcw83jMNB45YEXQf48d
xRjjBL+zpAtJ1fKeGtjkFwZLEcBNjX/4tN5pcW6W467X0topIAcANzoM4BscHGgC
nFHaDueEQgns/eLnLrXZW7fkWgMhUGHUm1zTob+xKcS6RneX1HgmwpmsuBgl6phZ
poIBhdaGOD5UiuP/PAwxCVU0skpev+OValK2eeXb/QaxGvLF6gXPWN68HXdAMvgo
e+r45+96rqnMSAlQguo6GbLmZbFVvfz1GnBJFmLBBo9DElepXy8PcWKLSRox2RX9
putSTfFSf1tJrslEdQFUrJGoG8R2Psr9zx9AvBK3zhihOKnNhu0fe4VeZ6tkaEiP
SvLVc9tTMzMVi+yOPa4GBUYniYkjaOKmNyzggOsUCqDlnxixAE91kFnSwxmG9x0a
EH1/8uPxgQ8r8FCe3q4A39U8uFRzX0hd5uBDDbOMqGPC6sJabKvjI8l2OfQrSI4A
sg6LU4T0Dc1slW//aSD/vrnFUsdBg9n56VHI0IA1K5O2UdR9MmbE/JkfC06zcA4H
t7dBcFhCEwIhWMkvcvclevlXRmhqj5RcKghx7CpPAnsCwp4Of00HRzraKydu5tvs
tVKbXPAOdLX+S/cvMjzz1qpHfV1Ygs0iZaTp0q/y5Jb3BSS9l4w/RM3Wsc2fDktB
7a5UAiRvrVa1yUiVr7pnAz1wtEDjIlHpg5vdrTnfyB7K+kvVOF9G+tRV8wPbqZ5m
Ef+Yg5dFzhhOx0NvtnAk6+9AEAbEBKrgUezmm0GCZ0RaLuRtn9dQ6X4gWpBTxWJX
i9dUsHyHZxvdjbcigvjk5NnER9o/NXX/O6i+rZTCP2QHL0O+lbfMnXLde5Ns6uVk
LgmAoftQddtM2l4zplYJcAqaYUkPbO/If1oedZoNxGeOc5OzNL/vBp02FVIep/wA
8oiA1dKFLy5clgYPgAnANxc+b7U4dR3bpw6aekMNDis6Ma+gmKfWR6N4Et6G7FRs
I3CbD7j4uAIQ/UouMGKp00qYJWESUSyPU5iXP4BMQZj3hKm9tQ3SzRFDmziheKsM
tbvIlx9NTQmHmun3FoXUJmkoxodsXBBsSomzf9KtVZvrugzCrMnn0fIVXFszUHne
feku2a3jr+GHbTGaQetorGSiPc0AtN7OQr/Aahxc5c8XIW8YBSzcsZGEdPGkFIxD
hqjW9/bjBCb3sR23FT1eG4dbcKMIZyoltChb6VcGX5ft9wJ4RsEUrNCp5OyNujj0
hGbnJSMUeE0aeOVL5F601zSo8753Rz8YO6x0t9crrox/lsj/FCxLkwxvWqyu3liB
7zzEUWxBTDE560AU0kk6PhRvSxFrg9GQjbOqbbxMzM7W0BoR3C5wFXFFOhkGhLrN
wDX6Y2RMlLM1hK4xnR4e6NmfvwyarkN8tgnAgir6IM9ngVTmlHj6+E/q0DOsTnWx
RblzXT4ItjQ7rBJIY9+dIuCsU34ztBBC7epSRf3sG9HHDo1vqYkPJiHUvYuMvbwo
Q6WNEzjlPBJLlxTSbxN0YBo0er1FdEGfkTEeztxnT8XMc+VbxEqbLf25NYaiYg3W
LB/2bhFQj0tXtW/5GkFTFi/o/zlC9sxhiQ0gP7l8Rb1SUrWUjVlCQ4YHIugr9Znu
LGqmtNcMz0YwHO2DXwtP/TwUDoy1fxG7D4mrDlQmxfz7kWwqkvfMXVQ5e/BF6+y1
KmFw77s1+/cZBm2qDsMdSuBebe90Be3KPM60zyXzRgY+6N1Pnpk3zkyYu1U8tWeq
SKlno5JvaUWLaIqMEtyw3NExOcq5s0SsgULw26DwBu+2L49cYBhyO+BMBx4uNWeE
v3hfJ+DdcbyxmwNnEm+soCsiSVXOGizAosf54pjOUiq7qpxupC5ImoXgQhleKsjG
1SnKDoVt2N4sUqjKTcbn/2jOIFigRbteblFczbhnF0SfTZuddKyAOBZ96XIZwQ9G
22Y3BN2z5pZ/mIq0HcnyPcdt31/VYXp1YwKtXV5iAjJ0V7uIqz8nkbrpnc4SLbLv
H2LwPV2S9V1Gr1Ha3fbtrcqM5PE76SlXdqQLp9fLkwGUQjLeyxgKUl2NJeoj2JEX
2ur6eF799i5VutiviHTtleLU2sZLNqTGAF08hKdHo3QYzbPbQETZ+cKRg4sYqiR9
b/wjn1MjPWveAlSpSmarrOe6Fl6gkoLjaYF/OU1i6VFLrmBkFfIOg7VGdfeE/Cej
yknTSYEfuLkQ8fjqBjHbB51cwxUkyrlgGKWSo1BfpktyBxOumthLl/6QNSohQPcF
um5dRQI/9GgQKJDfsySo0jRBfvReDhVxcOk0V0iEGuzJuIRuHXHiMJPWruR/XnWs
YdqUhD8K2Sd1av3eK4e1SfH3jXoCXPljT9iLhnuV2FIJGCAMRVOWk+4weqJjQkwg
S8e8EANgu41J+30F9jTlFYlY+OHczvhNkGoY8BNwZYD2mWm/5Nhth6zB62lmNcva
GFcqFjK7Yx2A2DqAr/9XzHHfPgkB+KJNIW21gUjTAQyAyxpvBXwYWBcG3O6XhM5L
S5ibCqX6uiOGJBtEKBTBBnswOb8nag3tL2/Ao3pGyqxtOLOO3MWQxAciU4/G9GyN
vaCUraM1/i+EXJ6Ky3Yhsdm9jrSzq0lRQqGRo6jb+8UlRkqdFUTpWAbQKgVeIsWm
BbCtnRlSFXwlw5qh+m7gIezCT+KvbSv1w1YIe4IqdtRWrQc3NIxqOPg8FE1t7c7q
BkcVz71lKmM9tmWLsDbdTT3rHnu+MTuVJ+7/bIX6h0L8NALf8373hgVWtNNwF74/
ISb/jBgxK57VyxOCqb/hry/vAYpRVPPP6uPLGf3ZhsgxklSPZBlMjERB6Wd6Yabj
3RqwegkxRzU7LR9htrbiIYTSujCw0C/nvFj0zIPlryOw37Z5f2qpY3RL4XVHTWFM
7gJuLYV0/VTGWpbgqCutMTR8ryjNJK+hU4w6G+QXOBj5REbwjGUBCm9jilnlcFDI
SF7R8vSGX2rdPk4fpOX5SutQtXV2JW/qZfTS2b/j+pQZjLBJg/cm230B9dYLtG6Y
AiljQ0Ow0HGCoUYfzWfI9MwyGPTcpmtyc4YnSGvUd0eneqpmBsOkT1zFS+iVcWVt
O1rYN4bZ+eWuQKEQ6H1epjbDyqoZXBQUWkxjPYljG4mF08N0J+CGTKkLvxL4CqxG
0kHP5G+3mtXcO1LmXZQuVVEoLVZZrJL+ai1xv16JrXh1DGfZd4T+UEFbXgI9vd3c
fqnDtH63IhUNDWwnyFv5WPERplwgHFaAx37r1PaREdGKiAVBIBPb14DfXiQsfXNw
d+EWM8gsxqBQ1XfXdBWejQ57BopQtney6VPGanGruQ+27ldl+RY/ctbyY4drXIQu
Dq1x1tD45VZb8wKhlWXazAxYF55F90XaFc+5pQevXgLbi5WbmMtW6MG8W5hSoabO
TfXd1M7M4a8f5LZWPZn0Zi3A48FbFowFZIaMOC1qJv42ZZxuk0ml023T/qCrbdLh
95CWkoejIiPv9elkwWOYEnEGsmGkUw0LgPpCihy4AJ0itHTxisRVE/R+2vyDhcy8
7n6g76zUH8YlGbPmlWjodlox/BaYFZ2cECRXnWnwD3iJPfQn5heo46blDbkqVnh/
A6PaFI1PZNaijOH5EUtZQTF5c2ss4mdiltRemdX3PZM/vXHHGXNCWfu82uhZIF0s
EjNJC8033BTKpJApplCX3BbLpib6T69gd0G8NFxUV064Qwb9J9+g48lyTAeG+mUm
Axn4XPyH9/ZFVbSRtl6oPqQFXCqK+lGM0cI1i9msBDa1YXJaXhaQGyIiLxzjfDAF
h48HpOKn8QgsIBz26f7q9p+LS5npJ8xeQSvudcvrR6H5+pJjLID6cjQ4j4FyriIs
G9OtATVMccNZfjuixzwnSyH2gcwecv/XGoD39RxpfgTZwI8ZR5fM2k3T3BdbKeiy
NZL4omCfEy3iQgRJcqq7OVH8IGHCWbTf7whG2TMTp/BCs+1jRlKqVtE+XfJQsOzw
ID0m1bcJXLgIe+l1O9BzEvJfedB/nsVN0T8sfPboq03bfpOVbzydnDx/bqhLQ3Jb
lxuwvNAMC/0rAny6AUq5nsYvTMHER0C5oAUK4MieRzNQtc8q1GlyaLuPHDlag2UX
JPKMzUmHmIEX0BIZGR1OV/u/m1Hk5QdJ0TOVAbh8KWfnubvAHnU8+oqkv/qIJdLx
87gxzC4JmxobiI5LjIokDpE/jSETsFjxYYNWT4LE5wDVeIgsLFejpG51cL08pTu4
BZyES037ktJ4nTo/1j9tGY260nzKm1di4NLcsbqxp0M9adshFZagmkEHkDno2zn2
g6IbQFXyQRNsWUIWUv0E2tiXnOF0uesdWwaOwW2P+lvnLlk7CQMAlOGg3HTUhx6D
EZ03JNZTMvQyZP8WiVPm27ajAhuMyqQ7NdDeJjPadw+QdbCVEn80KEyd+pzSR2kJ
/ToIR5F4yK6rQNLfAvWqFoQdwetDvC6RqCl1a4B/K/VaedQUFkfwqAegYYl2KRGo
2AXa8rJUg025WDwMF95Isaacr4/v0WGs4FqAUNmwDSJgDvnSXscTff4+3EbZ9c7c
kAchxp67JsBoiMm/azaALfD/8AvBiqqekvy0hu2A/F7Hnbbs20nMO6mvWagXzW7k
b5J8ExFifwu1dSaShqmngBImUrA+LblXptTq2/jgQWy9IrDSzNDywmfBSeSAXd4B
PW5qf/Sya9vx6j71kcQKxm2Mqp+0scd2vdTgrJNgo8rVscK5GYo4dfJ8sG4W56JU
IVGWIonWzRfosYlGgeFaSMg5HNY1TPgoYi9qBaNdmEFaC4/ree0tKPN0L+6UYJx0
pIOND1TDaepZLXdqNLdoqWcB/SiAHpyjycLRiXVUKJXlE78v2RitQjFOSKoutL7H
1oToicv+m/Ju+++anmfwklUyXQweFBk6jlIXSA1EhUPrjGwwMcE/UJQ/bfOoIs3k
vBMwn1Kc+PFBg9rGu4AisRFFtBJtlM8LGV2E2CvJzNOBKqyY7LQOigw0g50Y+xR1
iPCR8y1QYWFZGrafbrsJ95BkNc+m8IaatuZb6y2oBR7x5h3MejgCIpaFEVk9OlOp
P/UasjmDklox4z5vV5mMMONFvgFnkxSTPffXTx4OzWSTEbKdkzC3PGF/uSC/ETQF
3XbOtp9sXfulbbSGErSfIPGPAVtdfW/+f6S3zf1yN1M+2yr+TTPI1ErglBuny0Ax
mBGcFRwCMC/ohSBRUa6YFaqe8woKyDvfnyPM5WbGXecKKbOw+fmR2HvIpu68KoeF
9S5hX09qClxmkz3fCit8E9mp+wiM9k0k7AVK/AHPnOHnMUM1YsdviEjl5t2jJIez
7Zddy+J3gKsRjB7vohsTkDwFMoETJimPjB5j9BVrH/LYiqVA89wvD4UewBY6PQxs
BSebtIj84iX/LSFkI127jWDnULNjT0YIAHQcn2pcxLd7vfjtTnrhoCFVIrFbMWmq
ZUDEOaOjT0IPmB8gTbqqgcmDXRjRXSDAi1BZ+OKyOgoq02BxkAz7Z/MoFDzUrpy0
YwsOnjl8UCaMjnR6DlnfO0E34hgmmGKw6WztqmHroHoEzDHFdm2qz+BiuTgECljz
rqC7uB7/g/is14G4obu0ivZVawjoWKrRRf2xR+avyRk4Af4N6zgcYUPbb2yIYAz6
465HqbLxEx1VfauaFo16Jt91nPdwUVIhagyNEXiUNT4AdMKMYjN76f7QD9sxB+Xe
0Uyckf+fuaiWtdelgPhAxbniJyl9piAWn5YsZdvnnrHptOpv5DDwV16Vm7ITRLKv
fGhtqnGse/f1XzkC7rUIDIdf/7/N7dO7Vr/w2lLbbajBZzK3CIOFFrqeOnK9pSZv
URWzuTOxPu8kF/mwqSocBg3omeCC0h+rl2btCibZUY3GncbB3EInhYGjZ50ufJRT
7LgWxoXevcR/GkcjVArB6dthB5SI84XcE+7u91t1ZvKnS35f28borlVyUeRJI3T2
BqQqJYU4qF4hrAKsOA0P9DV80OmX7eJ2sQWxcAUxOmYxtdLkRBo1JF5MhkG4xPXZ
jCgItdsEmNwqrjtkTxYKOjoCTcGwQb8BBinNSr437i7yQxO3gvCdMfb0UsddzoJU
VH9NkTuHC4jVsH99q7BDzsrnnJx8ynTyocGOZVHps/YnQei2577NpnmwZESDv0J9
uf1p4qPR1++vadWFPuWHApuPjvUyFhgPN4oBryBUD8xlNaadV70ZUx2UgTrEQb48
CpqL8RXsBZ4YVtrjOlYsVRSpxH4h6/CXBPlb69sUcNYeqf8lAuXmdIDs1Mb094Pg
LjR5/MzK7KFu8fT+EuzJ/nwmOlnwtRWIHqN++Wnes52Z4m0Fk5feog0Mn3rNtmYy
k9gQJIwWT12ko2RHYS1UX1RnOWUROkwIdIIYpupEPb0nTZyvWy+4MPIhgF3SeAC9
QCiBa7maGntztuxfXevBSmXLW9hNcQVtQpqv3oCLbBpamkyX4B9ppFiniw166SIp
WfMPDTII24GT9THx+3cnf0yR0u5a0Yi+dBA9CjAKih1QVAbP8PM2BCDk9dYDCH1Q
yhu6QA64bmyP3EzyJGIDgrKke7tYTCvY5oNZyTJp/AoJxtfbsWlkQBKS+FCxP4D7
THngxWm41pGwJs2q59gZDtEf/ZHgaPmmTRG5mk/CLW4wRomMWZMNL8xj1EGs+tle
KQY7NwsXPdlBfgAv1ohQ5JJ4dMifBa4XrGyJi3CJJVbnPLjsWymAp8r4YDMYgWLk
swuhC5TISZZaIKk76dxs7Z1RqfNKDWzlTyar89EEH8g9JPIryaDu5IwJdctLgxkC
cnX5dHZttQZjke+2pG23qJHmggXKA9CFYcvPftPKr9cI0JIwJgNgZGzBJVVI3Jno
2y/mSmnf0zvzzqtpgcBdq89ucLCIKL8HVTD6Mp4vCzOj8RnKtkxkPsHfwFvkM9iL
LbgmEa6D9LW3H0+Tj2Hh2KxPNZ0Qgpq3kKDSCU6hSxn+bWOhOt1t+8bYrQXlnfJO
V3zEFhW418wdiWEbeBVQtphXcNybCVjVWxoR4s7UqGwmnYV7HRManiIzcxo0PB0Z
eC9gK1N2L4EWWIz0Na1DumhOxDZqoihgfEJyMHaWqDEY09FlRbv8ZJ/0VxvYo4s0
z5QU0dNMtyME+R4Ku/dVHF9PiK4lOYPVopxTNrGX1G/fKAKWgpiCX0Hwm+NZPJ88
TRgRwnLdbMgI9bX+Qz0BH9SWZBS5GZNmL9pXT8c4bcKlSmcdNBnR6YxatluD0wNm
GQI0wFD6tyQxqsikakkRQ3YYMOUfgnRwlC140WK/4D+94hemr8EwmSdan6+g4q0A
Jn7URdBuUevBlgXbPuON1pbbucD9e7ERcq2bfeXsjgjEBjSc3nc5EbBG1oo9p6Yo
JemMaUUdIcl6efReq2EtYxBGvNk4F0LJChny1FjtydfFL8/CyaXULn4RaNUtsvX2
RZVQlXNzU6PFx8pi3/uXnr3wjsP6rBblyd0evgoaa7GpGh0t2niiD/3N3ubaQn6B
ZWBv1V1HgeDz+1Kgxs24+PUW/01JG3bShigs9TQ/DJPfKgCOo5CCILoQ3JcfatFP
Lll4VKB7fjQVqV+b6k1Es3pTWTu2gu5PllvMAHV3+V/DKqUm3jvCNuCrZQH9qIuO
5uvjnGEV/YZCZg1810fXsDX3K0+TBa6t0E/8lLKeL7lAIHzPVmXHlP+07CNsGRXJ
ICKNz5Ugzs5gEIbe8a6VFd9Su4Sq+f/iXt9KHDD+FPVNf9v3+xU1rYALS+CtjfG/
yt80+d1gxWmEyRB7oGcTPDPL172HQR8D7RDiMa1QQq1831Zln6OuVcC4esR0VrJG
7e9DvGgt6jWDjKYYLjFxevUeV+uWbNAyuPONcEr63tHlQI7uXaYZ7OkdbvDJaCZT
2+L14rYVA3Zz1HvtGFiku9SW6+CV3kFIZKFRYF2HY/TkmCrv7ZrNOxPlU4v6heOG
eL5xQUCz8vnRzWvnNjSAO3RItLBTGJPUC7brR82xsfSf7G7Sjf1vtR8xO3x3tnOS
OUJxwdL2qVirH7f0RvokSmhPoL3xTZN89aRcFo5uKsQmOf1GtJXlLxxRCKS7E3hV
+hlXqI/cjAwFE31A2tezN+YD0ggXoS6XWUNyqkhgCwTHSVtDitD7HUFCBhtCaJ2S
CCRVCyVAFewjFGrkIMKGIzSnTZaCPMt0s1s6Jm+K9HgpHBW3BPr4XFcx/4wgxzJ2
dx2UHic0o3TQ16s+o4Ese6ZfwK/pv6So1hqN2dV4uXPPe/DWQSwR+0Q9L272nAJK
OTAwCPylHGXY6YaALVkVrb0XqlRyvqyLSVMrRMsgENT7LdLbOEfMf0nv9WbuZQfr
+hkU5jgdXipdjwZV/Z671VGxslRgvfnIwmuE6WsbJw306q57LJL9W5eo44iZbGVS
eRsSQlVYk+qawkBQ77X2N4V/aw73hIXRm97yXaKPsLuHSB00+F5vfAAQs29/GMnP
+uJcG+9Re2U5dKqgb/DsxtH7yo2wljtHH/Y0tw3ElNK/5EMu6MTGmJzCqcBLgcIW
1VE6AucdGkblIHzPKfepXn+TQwfwc5mlo5/lHHuK39DGHz9Uk+ieJ9WqENJiLAg4
9FZ/s3C6CTJKy7lpik0AaVejLif49dymwxj2Nsl8bUPU0VVTMQgjGxt5c7HOlzsl
x3oHt4j0Y0p6w00HYFXoTdB6QZ668tkjfkWnC5FWuArtdcMf0P2lUV++vs9y7oZ4
L8m65dVXm8U5ASMfp0OMDJki/hDwfVxjXBo29Ce68/2V0aWQYPCv9Uyath9OvQG+
FtabhyeeEO7LByWhttnoj6I5Enu9LDNlKb8yhkyw8a5MstptylGghli4ZZvXa77O
1UgCNJG9FeXAbKA5jqlBZxPW/7cDt6nTlaN2D4BGNVf32j8Pdn6Pu005fkGFCleo
fA6gl1sfsPqVKaAXfH5If70QgtwVPxjDHme6LWjINpvhMSG37B2gq1P8L4Q0fF/Y
WTbt5OqiiX4DmzAeQlM8Qh28OnQJPFdyN0alj2m4wDD5VGcwtL50mnF+GK8TfQ3t
t9+I1eHBnwZcU8zjjYeNRmy4aa7rI+ou0QoGiOsytMZBcft44GaGgKaAyK5BQqTu
SPLiCWUWO8rwjiFMWTbXZOjdaQUR3KhkXe6f3MSbv8nN1FzuuWeQNtEWePbKEMNO
FSSBKmbvbqFpAxZat+VbvNnavIacsth2cCcuvS58fRRnU0c/9T9eOx0wHeKHoKs6
loEWJZM+BEa1p9VO4MRZ4mEB7KBw2YuPw/PCxu8GfTumQeLx97dnL6p6UM0NDKxm
wVyXr2yM8mciMctMUFIdGjmS3RZmhyYAYFfJRX3MNX2vczAcXvhKM3P9OMjDXBYB
Xerh4lpF34fg6/rItX/mruv/hclSTKHx/3F5YvZkYmNT2OE0vWEozGhkBICslQ/J
UrEmtmd83QRHgC9OZmcHJlvOjLyHn2urXbRu24aZhk5r73jGhXCq4zbGsrLoHui6
jDiEQQmeg/Z/peUZnHD5V3rCUnF0i59b3xVfTAECxi76PN7USQVDzupIQq7ho4B+
mp1FvZ4HGKLbHGa9kM/08RH6WwO5PTRenI/5aKnrmmQVKC1SmcojyetT0Z1A/ziO
hZj1SpchGeFqaY42b8ojdQguZmI6N0VYcRImvJTPVBMuNf7GHGWZy71yiUIkYB2Q
7qQns1f4/cBw6bWcKNCdvxC2QQ02Uv1AVp8GdXVQweudfLuSKT8E5lilapnqbwt2
+eeG/Znfsp5GiOUvDBdihWaV+YuH0y3rHld0KyeDc0gVnfU2amsviFGHSKnszxXp
pT9OeeWcIuNLWN4ThHxJSkoALsh3a7xqXIov1vtEU79HZpfSeEshLwxAUoflDaS4
3c/RU/RaSq8U7AGc6Kz7vFMbVAnN4Jx0SnSBeGzxh2DueQ83N+DahatECHXn1Wax
NNTuSNo40VkhkJEeLWGwXssEhcg2z+myysKF9sg3+KY9R7STQP5D3kDakDm+bfLY
BBevOPNAeSA2o7W3NZ2/JlaCoqd3me0sE9PP5usxt1e5LcyE+cgryslJmRA7aHv/
/6yFSfmNlonFUL8i7ZQxZ58p1SB082ua8JNf9Hi3rhC7uzs6mxELFuYatIbrjhJu
/kL5WkuhuiWTZ+78TviYsQsAf09nHINQ+Ti/OSJQNHED9qxEXWNQ49ySCMFRjkYL
g1hJ0mNmTEoE8tydaFg+qoZpw1WvbEZkqrKa1AEo5NHv0zF1WsWOmZuw7M/Mwgf1
svGXEEvpzF0ZpMP8TEdPwESEAXiPc4h1Qxyla5EcUV//1Os64a9K4ZTMIMFB08u8
WN/OqthFQg7qtv9L4FenFnTYa54iN2A+qc3PYbJ3lVmFB8I9doPMZrFsKh/5sGT4
6WSQiF4KOJSucyrykkUCIzeSUb/BNxmnFOZHf3wRzoFwX7UNbANI+6zwvjV+P0i8
tchpCreiT64jt+YCrW4FM0zs+TzbqJdt84iCTZB717NAToGe4ukcVEEWlbNZZA1Q
5MRujPNBSdVL3xg+twIzgSFlUmXt3PoIo71YWLDgsrA/1bjZIlJKt9R0fsDlxTcf
uERzT7T55G1+gUHc7c6kmvoPDcNWqn/7ZjsFv6JN007ebuNSzFZUOvuNitFcCAGd
9Vj3f/rVc53l57XR1SumYUq5lz83BiHEI4ks14c4JNOLk1yN8W7AGE+4TxJoYBhi
pegOCdLiVIAIMNIfpIesWh/xImWFnOZM8+m3PHJstdd53Qhs4cGF3Myox6Xb1CCP
g8a9fgPseg3NP4PO9Fct6W3gp+ZANzyygoWwsCQ7XfAswC4/zznJizYx99FGhdgt
mFSGHI7aATrsm8FBe6Z7y/lpHnxF54YIhwwJPlMMvwux6+MOHZXtSEmJLeofVVQd
VuK0Eyj60tFnGaVo3yvQbDZLM5FefMBBgW0oOWe3jT/pt2T6MA1qVQeH5jREhri5
y3DHNb2HOQYv+VDgDu1IBLdLTwv1cECrArao/521ZWaZjpsqcyhYMsKxy9uig0mE
RerxqRDUmSUGuHHAy0yC9TT9ccC006BXwdSm4l34TG9zEvqBEgvIYzc0vajVF2Ta
3/pUi1WCgf5QODQlz1cmMh4sgNIvI72wnx3OihDldBBhVN3VT+3mOHx4wrXPN3jD
3wPPk+sMmsk0JlOAwulT7Ly1Ewpm0nvp5TO2o+Va7cAXzrHVPp+84wXhSuDi8RN7
Vk4qly/fdqbalorRM9OPsM89O0EYllE97XdR4Mc6SpBiZmxiAlQlBO73C4tZzD0+
4JEgPI6/HiqWZmL6tixhZCGM42uqV5uEf7AR0+W2YA3xs3eiAH7KzXaCaAGY8MVD
h0aV4Bmua1JdjnPsb4zSdMsjlLlNkQGa9EwUE4sSs0KbMKh25iBPQPHAavhhNKaF
KMen+O5Oxe49q8/XP1SKTycGYaQnp34LDvaXpxbRh3rnqZWmPMVKrAFrm145rCpf
L4zxXw61tGo72NVU5zOinGHGfZZBsaoLjuqmkc6ctV7yjuBT8Gbuzpi2zZSwG8Gb
EwTdfarm4nKBKsiqlypQPOR/L3L1o+HIC5CrODMrWHtPwrdgdiq6lgFcexZWegnT
fTPC9bD98XQZtPhykoyaBJ4xWNPcDYHL1ZaBUh3fNduiJeKJhQcR2Xhje6s8YfFv
7STs/Kuq1xrzmripgYtJS5mQyp31b2oK9E5XU7ysRZQd/jcVF8K39jQH9ZTXLO8T
WGPKLWBWoYv1pcIDPr/dGyX/I4GaT2HNZf575GAuVw0dcVffyhdMUDwlItTegffA
j7MDj9+T1oKXWL4sUl1wxGQOE0XiQI777ZJ4KbZ8dpmlTmRhVZkvc7dL4jLYgEKG
bV0iiN8pPMgwMz9UcsenYbdWKSwJgwb+kAN9lmdesSFARlbEgVs8I0MjttgC6mDt
nT53RfENIUL3EhzHWjyLn09sPJfb5g21oZt5dM7EjmSXM65Ta0+IA3481y2Z4vJV
HOOnqzY9fMA1hG2y6U7F+Za8Ktki45APsi9umHMl9Vi8TUhI+EAHfA6smraevfWC
cUMeU2AP0LRYqyf9B6gAUAlQc6wnepulQd5R9s6OigJR/kfiXZeNZHhxhQJMUeAf
gXQD4BtLKenP0LGkohJXjp7Eo7B+LR5kG2xoWawC9Xx/Oq/AhuoYYAX+08nbtxpa
tYTs5kJ/gNrkja/7ddxynHC2XckRQhDEklKUs/cWjBqkm8FUL116rc+wq8AryFRn
cdqJW4/qtCC4kAbyj87zavdbh82uAON5Rc9Xd9uxhH4SFYC90M+2/40MNKLE+oAx
gokIdUDAaombJCANC5ihxekFjcO+U+QjRqpb0Q2ZpFU+TpSEffiH4W4JtjPkbXrx
gVMBqM8UAELQQpDAYK/Xhjg3Gxta780o0RvHUUluDh8/b7PplvclbAS4PI8bo89m
AR8WLM/EUg81qQuRfovEx/LnhGBYaeTrpEaQlMnY4mPrKghb2ayznJyT7vUvy5Pd
N2GZEQBujoAH/FYnJJRpqYoHtEIOsy01njCOfiJqGrRNOLYP0wJb7Mu4eGwzarYY
qmnlAMNxUKRSDMzmorvdovKO2YBYlAIhv2K3LCccmjeETXZ74f2kaAS7UY2MtT+e
72HbVQGMV0fXmPKlCusKzvlUGJ17+gvc5gRCZGWc80cppblX2Gi4NUKpWcx4FER5
VJBXPwZl4owMLuvlDRNT/lGWwZPcP8YwbmgJYmd05vkAoKIPga/ZQ0nfHski9U7o
eoANLIs33mhFBCeuvCyHjc3sgeB3QU4VHMQ0BbaV8WWPepjeU64XRME58Emp/HxJ
9pt0+aYoHwW9+XnCD1vGWAekCDXvI27fgDFwlRZtQMEPRbJOyAH9TdG0l7BAB24f
2NE1p9/hrFp1eusUcXg6ViVT9CUZLCQEHkgzr/z2EtZJoXHk/B3tmrezxUQxPrbv
FFjECULFenQCGCSqxqkj8+rFXAZ+Ga0jmEoiBwFXypDFFg+LkCU3hWjl/wNk0vd7
U6R0BR1myTKxhrlzXBl37AeNO6kNg7b8EmIsYQFSeLksIDJNoUEWO04DNRpaZtpd
SnrNYPcvL9iVVnPadVQdXVf/xfRwaN96rpKHKJ/cX3K8Fl76fwKoeYmWvx0GVPcw
rr4cmqZe4zvGe52gfaQwsju7ZQxBxOga5BO7PUtDe/mxfIJov/7WL+t+55lDMGAw
1diJUXtKCx36U75m4DNA47OtSaXcxXV6DLNveU5HM9ctfg71MXQpeTAb1FyhzoMh
y7JThR9h2q2W73QZ16R+Go7Lui/6l7SOLZmdhb18Togl8BIh8PXRIkoOr3l7pF7F
FoWjjcS2wJGnZPJRUkbkChahsBRqKQptNYiw/P82TVeEaIUOI8utikM5uylYFVft
BmN0bIKquwQlIcwLNrUd66qsc2L3jyJAa4crNdOkYYvpDbMrcAswfSPp2TzHnrkV
yhcCl9hciYs0XH6BgOFHmNXWuSirMl4k18lFNghREcuaeUvmHNKVaP6sQBCMcivc
cPkkgC53+CHh9Otxto+HgFqj8dp9W2H7d7STm4X3YCJfqkw8C5ykx/2XnvqUsymc
anZ0ObkcCk+t2lP+qBFAnomyA2GZ/qfJLnFhq4z4dTowxdtWdSbaZjB095pjPKP8
Zs1FOgq5yhAoJGJDOJ1Y/9IPnUVblmFKlwKciCEHoG1ZUrcjRYPnlR8VmUvUvLee
pnvwGW22f5cBi+ZSLEB42/GW83xkAcRdyM19weWdIpBhc0LiWl2547tpDfqCGoRB
Fs3rm1CGr0q3IWXwV1vRkASrEXRzXQW+NT9yz+rpxE9lPbXGbbmR7KPEHxSjB4fH
w02avBHoWBJMLKdWRDhcOECAkkWeDJfoyGV5MlxmnOMT7bLUMQLSZDjUq53Y7TWU
n3VFshrG9wVLxh7Nf3Zxg08bibrih3rQYPC/eynWZgrbArwpnqdt1AdApp9B5vdA
SGg1AF3oOGfPOy3vjtBXJBCTGq3b/WZF1rGfGdG22xHBC3LUKDYFPSXW1+VME16y
2pSW64RfD52829BQepa0/T4qtYiDQWZ5P5PG5UCA2ZQUdDT7tGryrfpheSiYTQeB
7aFWGtEawmnndsRSsrH+ZACB7PGJ7jVrSq9vq2Wf2c8V1vlZF5HUvxe1T01tWxGs
nCq1Zjou5xFyyhBbqwgZZb38bITt1CF3bRhLFn5NSH4Q6dudxmOd7pXycd+x1JJj
iJikTtMeQ4MX8sN+9pyS0OjzpS77NWVKgvNOcsOSQZhBzKaEMHksKSROkFs2RLPQ
l80KdsMVRGaEnU2VWOGFakT5kusw/O3oWflUkC8TDkyMBGDr6CtC3cJGFOy5oe86
3XqAFwYB3S5ksKSwnCYCnIdxEhzl4M8/kd0Tf2nnvIgeqGSTBCeJhDC95jzrecHg
Xy2HvcK2ceYrJvOHmc1LikaWQrI20DyhHBKN5f+gH6elW7OFZ5UC8j6bJoTcu3j8
QAiji9hPZ8z/7iOjRec0nz/XGFOBjIMp5akkJglxVuALhGS1RuY/nlAAUlkOj2R0
C/2XAR5THSz1POTrf0fJds8umpo4AcZUD4X95NcFlKpJ8SANFBTVcKcQ3Agq1Gtt
3A21uGYYLw/ZKfjDH19AVCCVOZA5MDplwrjF51ahw2W8KHm+841SjIBWMZUKa4mx
Zk5ZM7QTwoGvjhXHBcoa7GSCC8Xcg1+h2Q+XpHdDXn25MAprJIyTOU0Kc3IDYgWk
Ze9wkOIzq9tDaTe3vRSK2FyXnHiOreUynmXvIH3Jv9rCUtHKsAHoyYnw7IVQflpJ
x/sQDtHaPbvmrNDty+/VAwlJSL3Rk6bTH+7HJ0CtLgbOOJ2O/5iEvsqfMaB76o4f
lttFtGHFahQ0LNq7Nj0TTlLhxXP5ZH2ubZLP+5BSTNF/VEvWim1LIszbOt+i6U2b
TkgdZbbflKB4tl2cl4qbTWmaC7e/CiB5AnOd6GNz5LQQD4NX3g34oI/wyRYadvIJ
x2B2Y5RiwPiq7GBbM2L4W/WGkPMiMUW5SxJw78wvagAz17DWCP+IcPSBUzFjzlK4
ohAI80ar1O7wYBzCU82h5BW44FGywF8t4zYRRkQQQkig4LkoGH3M6LTK3/f0iLoo
i7RyPSaqQxTFnFvA6zR6iuLoiw2zZYorJUUqwbTIGchnNCFC/TSEUEa5fooXJjJ3
8b15fDGGnZ7YAf0S1HjmlFdV8GBRMIr7nbxy60pYUGVQfJ2f+MlviPYUqMehJcD/
mLMsMLYHKGMxRrXs9jogkoBCaBOt3GZFyIp9tUi/97YppuuMGMnRo8YIA8ylWV1s
tYWI/c7aw8WBal+e0etH/avsS/Y/Jrfqk3+Q8+PH+LbboiwXXnYxh41kkzivehqC
VawgTFvbP4kzc+/Mv2ez4a8xqZ1HYSbktJIuqIF0pc5DuwhiJDLgfyR/pIdP5Ig3
PdtdZOPQfBVPwqR3h3IbD2Q+DdVWLRD34bYqjjzsF/AqrNiuL7Jg4sou+f/oVruW
NgSkx9D19zvAChoCrWqk+vO4VE80EbkG4MMFztPVRQjk8ZOYGt1OAltXSYMtMADG
8rgzcKJJIElnVp8zCrAshR/hy5RRXp+VZk2e9kh3oOFJdvBcVWQLBKG64pdpuSFL
PV1P3ltxmyzpqhIcFkWpWy/X5qxpNKvid71m764fyKgY/lEXAY0tzbYSBoTfjuSw
GFqCZVkkZAkileM8tzTFpaECwGtQ5pQMJvcpzO95ZGd0/cwN83A3VCkxcWLxF+5t
0g7awT3z+XWADwkF4iGNDxZFM9VO3I5ALcErmjSmFHin8/xowSYSzqnHSAlKpnlz
LyNxNswaVRoOhs6BR2vw3ap4Xu13PiI9S+LYWiIHmmDyjxToqmTqPhcF4PYjw2Vz
8zcQM178aS7XF9mrC2lcFDCw23FiUpC2AYuAprXVHzBX3XHeI+1MwUJhqntnKnde
v57xBmTKrLVN5Bkm/6OEH/Hl2Vt6KCIcmJxuZOTWspHCYQOHnCVdn6BZlX3qNadA
rJzmrhoZzNA8WyMQpcGKmJhA6Lo71hcP2CZ1QRkMc8iaXS8tVlRwRuM6NduGkaCE
1LLbzgfZXcfl12C5FczzqayWaBh+Kt6Fu74z92R410oywLCsG77pADr+gZiazbuz
a+EnwaHckF0RPm3dgiOXzhtezFhHEoIqpCoNB/rKON9IDAf3IpfQoisbLyXTO25S
5dCilLfsPUKtK8vthr2jPk3sHv6kAs6QIxATvd1j1A2yYb7bcmTWnmRr6R3Pw2H/
h+dqEx5ReUJQ/LcA4CXviZBiAtNGA50o/LTgc6NYILqCH6s2QcvpWYRUzMupbSJ/
IfUIWvxE8LYnxo5cn4j6jJ96YOdw1yd8rHbUbtrk1w/zTHAan/YeQKmBluDBSg9X
/FpEKKrshbz8KpfDG22U0wAp/j2rkV4wxHhx36XN3rWJAF3BkvcpJVcEDnCLNkir
t83oWg2BWJBAVWotR5IVcbGOBR2eTr7bO9J21rUBLUMBZDpc2/uMJULi7DHZKU/u
1ZweFoeuwcJPCZuWUvGtbIvoOk0CeUWtESzNQoj8sanWeClhsgDXRyw/HLnyGdhC
DObAzB0W3VgZ9kSyj0+ohG0yzcWLFbwOFKDy/hQg1FL4Y9Z+yhIeNWSLr4pq7Xl8
FzERaGHjTadxhe1Y3fXCnw/JhV1hmPGjEGb9ZpZExNfedhOC7SgkywsneJZ+hAqX
jSwas04iSgkloSe/ZLGDwuGjl0Cp+lUQvwh1q4oga0TEemn3JUAqqqKS/Jyrcj9v
vVsDhTQFGoeY4/6dWS5W08XgMU5yk8kfIAujX5dJCrFu+fU1LNKCHA9abHiptxOY
WiEUuoEeDwDPNIOudVztyBFbXdEg2wkFNWhe63ooxwL9Q1785vvyWTwRdlOFhnrw
M6iTr0Zqsmg+vartVEkLXhysuPi6iJdxxz9Dd2GXhgMvI2R5c72EQgReJcvnY8vp
voYGn5KrJ8AYcWl2XAjD3FObe7Jb+mOzHC42qcS2QF7acgTUQQgDB1JWiXaWVrRM
FQeWs4ceFUXMADNIw8IqUNhMIqVEukDrm/1VG+1SBV/6JyxfP0/Ru/Jtn8btoZFP
AzIJ35PNkLf7v1pjzzMFugDaXmoEWlDeqWXCDsZwfhAfGo5nHGmOWv2AVwfTDX5I
I0cqRfPYyXFRhzjh9DQfIhnAhmS0qFcqayBscx71+x6vfWAs6NksKesaGfhz08Qb
bY9ZCM7tVpWTj4LgGM2zOMmy1R6+s8O7OmUn+a3tAAkwLsrbbWZeEaoY+pVDVyy8
cs+eR53UtuHuiFCcbBPibB7V3Zn9OiNk80KZNavHoxIK6dp41g6xEHkbH0dBDnGz
JvTqM9l8/PTRjNcwljILt/9vlCX50xHF+YQd91ztpOzC7g+xzBDn+h+1I2zbio2S
+ZjD0eanzWtDGwMgQWqCKUjUHd8iOjrGokm5fjJ9kd+JhUtsFeTHXtCz4me7BK7y
DDxUmwesm9K8+nXFcZkvkMGqB4M54Z53YxWCNNdcAm8R74rMlEAlGUkmRLkmz1+z
7P5G40XJGZTBJaUygGXeYN/s69prcx7tFpWn3Z0FFtc3V1lRzN7BLNLiOeAsOpC/
nWQ6xszMdmdIe+H7UN6tmzcpAe63C9rbYyb6MeKaTxEbhTOpBosLo+Z56YRDbqeK
sc86MgU5OC1HFRYucTr+rDAfc4G06aeU2DgGzAbtzMOV/OTyhAx4RbY7F2uZcCYT
fE/2ixfJ++3Dq1btS9jw43bawVPcHjelexwJH4AUCqQwymTXVflOTR+FiAZdLpHa
hmMtsOOsauOYqFMGrZBIPDOV8xBtIYHCQBM/egcFjfqzYstWeoO7Y49dBhpY2esg
z67peGHyYzRs045HAGV/Dgi+FD54lad7dPWuW8mFhEFpCDkzIi4ncxR+PX9f4eFo
2ExPJsVBYxpI5r9qNxB5BUk810o3zvn+NrN9GfxpPnbGg8CZ4ulohG1XAuitYcMb
l2jhVrmByTTLCbilusrgH9od5K3GUctv7XlJu8Kge3iBrRy91SLOw+hp2yYVM8Cq
+vCeNCQQsn2Z/ZTyWzNcLM5VJf0fU8C4aLiPI1X8RVeRd0MlFbmmwcSUnlvnJ2Y1
v20uuR9dv8rwzwrUzV39Gx8bBQlVS3lL9yma+PMsq4/7SpgUEeIBa5MS2C2MxdPM
q5hWqAeouJBKEALVcoQbLLBm8sk8J4HGJ+DgFBCSON3W7CCXzfsEc4moGAuJjcKX
N5SYtFws8FCVA7u1E6Dxv6sBrVFyyKSqh4NE1jjv67AgfinW0swx0Kc3bj8QeDNG
oyB0Ol9ZQmUxmSUcGVH9FIMtznwhb9Rpur5cHaiRatLQzhQXP2UNDG0zeFfII7Za
WBkF4931yQ3LiZS2MFBeKHYv6u6ZODOmRupdHx+KIWPaH86m04oVT4YcMvBmkuBS
LTY0ldKEiCzeUWANzrUpLYkhXTa7LJcXm1CNvr1zCjfUNt/JGnCuFER9JxYYonyd
3fCPETP4XVu72oXVHYAVmXUNQRKYO5/7LubK4YtdcX2L96QJ7W98/btbN3JgRUxN
47NSAufgvYQWNYfSpGiJ1OLe8PWWwiKphp0Djwh2CAolF0H+Hf/EHse/66Tq7VQS
9vuGM4OfHzF3+0hPJg3em9/elVvgZ/qyrHM00XCPoG6l1fYuQ0UHHcW6AlL3Ec9e
m1WZokaKtvwo8E818gsSo2V7Ho+uny98lHzVAVuAjA/XgEVeYjXqnAujkbhtT58r
OyZTFh3XXsyeFVQ3FkL+tCUjEkiTYOEb8GnIfdSgeeMjehgmoEajQNGvPDwLgqtP
Br039cRRdg5sA+7Iu0JV2wDk9ojoA5Yd7hCY6V+tCy2eyt6sXeiLICWLT1TRZ7Ly
NGOYtcCN+kjNYa10RJuVF94mXEN/LKTa+jcKDKshCsYp0euxk7Tss64EDXlR4oRb
sAUpov/QX/0JOfVHZyJw1i7cUg7A0Dk2jN+dgifn1YJ7Gm6f0FAsqyC/e1xU+5EJ
To6wVpegzrQ5hsWUK9g4+FcXvIpkUhgUt2mNn4oUmFpY2ci68pmZoVtqO+lxAht+
HSHQUr0fxrdGeoHUls2E7dnGvilYoYnbl062yAMXULzG8svwVO8aD+0Ar/s6ko2i
ybvpHRCQHdQPwjIl2im0ylBSVdWz+HR1MNIywV4xXVyMl7qh2VuXuqAwCK+oRb3U
9ensCQw4L3Jf+P3y/xLHnd/cAPFor07q/eKcXjDOAQ1akosJw4COqyiOzyLGvIdx
fZ4JkKUiPm2E0kvDzX98z7vJi2AOpGQlgnSDEgsUPHYX+EKh2LtX+Ovx4Rv+L3nn
y4DbP2J+c0g+dm76HAFcs6LdpnmoHqripzPr7Sml2DCwYtGXumiG36t3WGSCOQ01
/zkU4TjsTHO3OkepdTChwv5tf6fyzRdvxlJzq2wPUkWVdNWYSqkUWkobFaQRkEDU
b0WdvwAsrmFyd68w76EOMPs1WmXb4W7LpJZfoEa8etDbO05Ncx2TzTmYirLdERdl
9EZ7cHH2MP8QEzFHQ62bwJLMilxb6DPwhjwyI/fDYXkop2jcv/tlk5ddWCY0GCeE
HUOrJYEgo1+i+QZz72/PFjrEFMpbSQ75qizV9KlNttX9FyUpbQOM7B9FabcMbQzi
ysnJ9O6Yrbws8fv2GI8MmdM3HcPDmkRFFeeMAAy2PSXV5/UaRTXqAAS3We3vaz+H
r+kSJfaCjnQI3EfSPa+AJ4AWn1Zly6w9BWv8HOtobMT3r3FAWo2hYQfDAdOpDj12
ldUJl6W6hcLtjGbdRyHjvqTlVoMIoOh9G+fLwBTuKS5sV/rS3LwhjvWTAluwfYZr
LEHKEinU26ojzlxhib9LciYqccgfVBMOu4in1Pj0j7dv3C+pdSr6NDc1/rkHtHU8
yhDQ+n/HP2svgKDhjMySXjV2JClQR2eItLDlmiLZhG7n4gBrD8mrDJqXV7jg6Rza
R8vDwg2AH8xtmCYHHjS1rt93Ii5lwljNLtpdCpgy4e2lI/B6azaeWaY9c4+djyFk
4fl4kBR/GC671nCysHdrmy09kU4IPY/k3GXC24fvjK0zfDLfci4GmZQ8xWF+Z4mH
OG0oj5LWJSYl8q97x58nase6FstID8gadMHfA879SIl5tC4zBrl0d8KVbO+0CGV5
OP6zvtn3oYClTB2YmUFiOCvvptfJ0E2rH+fYkPP6d8H5Xx0LaibQZ1NNsDc7zWFe
QdMY0cgVvN77TZXoQrsxagbuuJhrXW0oPxTcZ/bx8kVcc2iFyQmM3BfyWMtNQkhq
nIJ2uLcN0AT4R+drTTSw7CpPcky1FE8/q9JNkP5AbcaE6Xvu8XmqMcPRIZhw4s+e
OnwHdRcs6XOGUc9rcQcJdfV9yjnjeAjVSObdWLwtoxuXCA4ZLHLaNjCjNJBlO2wb
iz7agkfHB3AKR/+xOCAspq39azK2JBrqZud+fQbaTXGqeFHOtep9zdBVSPnszBiq
eWrGedUZ1nSVDfzOXit9roZ5cyJ8Q1sLrYUjfs7UV5Rt/3BJLAbScsDtYiHvjrJm
KUFRUls5VC0cdzqFu3w1kaJ5dcIyp6qJxGnDgot4vMMMLsdfyGDhv7bwHn7BwaE7
KcuFd8B0cinmi/B43HGdDxKijvgSxxUSJEpowxtTH7I//PZO3IYE3kEaVZZ2TFDT
zoFBvNIcjbAbK/GKjVU/5wgEOVHK8sf3AackTagy+jB2/IcZ3UeeHRA9Ef3WEbsv
rmZoo34R1/PDrTtg2YQc+o0UsQ0gfZUu97okhIwyLF4K6ArttljRY9fuvHIJl03S
Mr8ywU81v7kPOMF7wJGTs1J13IrEUnfKQ55DuCWSHdV9Bu++F/wWnPuSBhYtY90B
+DjUICTy1GHOL1ntou3Ju0pP5/Gg3uSPCXbYWPeNXSsPz2JDQyiD3O1TkngG7acj
f1ZvOqCakErq2TXs4LhsnGAnBkmGZ30gqDHYRV++Dt2Txc5speWeAe2KkHmmPn8f
iYMPRUZnG9wJmOjr8LuC84tK4OTP+fSXefQEOPWNcxUfwWZAx2s7eZBLjY1nkNJS
UKKCbHaqkyXbLLAqn8+QF5PZrOIXDyO2BhXiaETWeE1wIFj6fkDRufF4lgTj9ZhJ
fAE+A9V7TjDqHNuW7jGDn4V/oQlwI7PN+SYzcSgudVn+ZFbzk04TvpNcBxQc78g0
ADyOwnDNvkltyjSr/HdcTIwTM5v4Vaw1xkEqSszcVyoovXI85WldTN1lgPJnqgmr
6UYMMvJrJgukvMTJPqkgriz1J1foR3yjHpxmtTGJ9fQD90HXQkrBRNcpdZZoZbOe
IK/FgNBAXdmP8+2Uh8BKF98K4ThGGMCjXUYgvLLgT+6wgPeTgASnBjOWRTStFlor
wrVXF0+jKp89WjpjarZwAG8pzD3nGyuv4ipaZJnkMsnVH7SYmWjmvQP9QyBwHFTM
Qpul7m3TYVK43xmcBlcCKVp0bDNfd10jeVZyf2U+kIBFVyMZAPp5bwkcsDazgMQS
br1NW0Ejfw2O5HMTmzFGpehqGbEamHOlNswI18nivfvfeV61kbDUsXpAkOVBDeGq
4740OBBGpCFIHEEh3sucFUVOqQR2pFz59YMr0KopoRxPlNwKy/OnAQXdUmR9PjT6
XDYEf+k/wvv19AtKwSS4kcdeZ+k9+Q3W2SvIYDLWXRXdfK9K4fr8d5aWmoAoHIGc
aLqqOrkytkn37h5+0spdauwIgf2Z/w1qixrjE1mB+kLgWJrBiTnKtCa5CYkVTyc8
d4kUZdDxxiMGsd4RM9haoG3/DpUsFFUIhp2U+bY9oaPYDq+KCh9nSyJrkb40sSct
E9DZF78y7xlA+j/9411+xgXYIUx13q+5VAmUH+gLcKm4QEuivTc9p7+vl3R6cwGm
z2WSv9GeuI+f+/8De7p/qqb0aNUoJDQPbFaBQSWOyB1o6wC7tUh7pt4FKYCiQUlK
OzrJ/OhTQsN7ad6CcQqbh9qzZPQtJwBSTtBkJEx39YHe+xj7tJVP9x5srZtnq62l
cqccAwgAo8T07mZaKM5A0M3kOOkp1WCMwdpRMJJMS+nC2fuUvZDY9dwfAUbJrZtA
qxLiTEry7wZ66CSLapn2UO0YSPfriL6AZjrXp2NuON8piGijq/syK0Lh8bjd/+KP
VbJHQDw9BqCZUO9GkbbLDXFXa2vB3irprEF8GXw/hGRCFlRWMvrVfAowCk0i8Y49
PwoUDTryJuSFFljZ2sRhWQYanJ3ocG0fvO+Lkow6qAH3ZFjyxfsPvoKg8Q6NM3ez
UgaYmKwd32tx0SqooN0UyiVr0Wv7zFtagRNMOmuR1OqLzlWRp0YLlT9xkNS6FUEo
hrDdTqYNpYjTNNerf3l29Yw0wLyLw8lLtX5DigJ0+cu/kTq265HPo+Q9ZgLbPI+K
nVgyQoZ2cW2Y30groGr/fgz5oFkYJNzv1PHE+LIXgAxtICLIhZcFq8dz3XYFwsV+
rdMgzTqYxMsOO+Ao4m5vPAeNjUHYfWNet2u4CBXdsb4MzM/dutEXRl1GfuK5WMYu
AtOQb/se8Sd/tRgkT47+HBrvrSFqJJl0cY6pLyKMZ6PCWCStCNmTJ2+e2BaWEIJx
nPMSQT2P0TfGJ6WMWu4OggOIV7dLWTxqpxjvFG27CsAgfS46TZCMk2NpEP6j18sj
gBLM6JuttdgVtUfhg4aLwzSqwIKA77IKORGmfkeSj6cA4owpbZzM4TXsohD6JEqe
G96ggO3UM7PaLPgwQJS4UQCJwHHGlxsxmSvnLfY36V+OFnKocxIsGfD+e/oeE4+w
9uRyMosqkp3QRu5SPhmSAXayi9T5vY68086NU171t2RoQsY/3QzfafDAfzOqFaeN
fiyVOcQS2thvq5tWwHSZa2eQLojoCFF4jC0i5PEsPg0AiMk3oQ+YMVEAND3dgdbK
v9nlb+knACGMrd16LlXHlJyNt5fKaMuCBZwkEKZXhUEohaU1lD2z31i1GX7V600O
qovCSWFYRM0RjLZ158e6vm+E6FkCvs4jdMDRQ3h8ipeha7aqtyOJxNQQUwrt4Xlg
zOTkxGzlauV6y+5OOviGFXDrmSH5gpAvw04uc8h66uYG1Pg8mDJniVHatQWjTVOP
/1r/8Q+aJ5JEeULw638Joy+UaVqzkZvktKsCXRdidLyvkyFJCCdVjMIEfM9FpFoo
V0K0qJ7PvC6ijQgMZ71XbRyAdishr9wD/wXxZ+jlSK+AWttHDZ17v52HwnGxuwEz
Zn9SueayMatqg6ig2+IZ+us1KtQBR7DyZMXlgFJiD+/qVioD22FajMKgX8WCOAJ3
VlMaVk9v3GpfrQKNscZFDdVwOPlWw5qf44XwsVHg4eqbxLt+A3rGLi4dagkyV5cr
K8NJ0tckVU7ECHped+7McFgXXSGpvAfpyoQCmWJ0wQRpkSxt1TdleHOlZi+sc/az
Hx5bADLA8quvAsTaH/YOPRtKT8bbw+PnpC7Bdw+ZyUM90PKqNmGEECjzMTSl0J73
DfNCxizX62CQlB6EQ7bdccfDtR0RUMZxo8suDrlBlBaprqb68hdG5ywNZJRIf34u
R9H8imd3A6DuCU/Zi59M0IY8hXZjppHcMb59d259QHK5FvA+LTGJfgcHf0cuJv0K
gC/RxYy9xtLVOI/A3ZGn3t22bPcYrh5jqheNda+hTPO+AbTrSE4zispia5HWOqSb
T/VfxZEsc9N3ztk9qNP5SZGM2c1KV/7TjaVURPQK1GCKZy6ArWCxI1p3OeKrYY8G
ZPzTy2BstkPnfuY+i7IAXyiF0PjBObVLNc4Xyy4aG8lz59lD+/b+jbMgp1XXaaQp
7ikO43kE9XJylwCPCsitAd23LUK4Op3lUePQ5R7XL8bgBL8NnXIIZRUppbJe2aL/
4Z7ApaYPMQGWo5/z8dRuk58iFQv/QxRLV3Y+o8r2xsj4/IeYcHtoIvMNCfsTwxWn
DgeqCI4oVPChObQXGktU+skmplY1gG0hsAR/sHKBd8jfvcxw0crE7C86IuZ0SN+e
mO5LQbl1WkgLXWr1xrYTmt9BPM15jrH/EAF74nkRPn9mPr+e7O4NPQ/Ap6cbZ6BG
lWF8XIFyh233gigHKNUOtO+nyk000WR/xWqWk8Y+Tf/gCHFbNcaBxuC1VJG+sGhm
NiSvppTgX0FD7T8K/mg0L5MXuoxa6F9YJxqBdzGyVgYdFW6Inr8RUcZtLekp/04H
KWpOkyeSvgkupU1T2XQc1fGz+fAnw0Qq/yh0yIL8PPRWhiFd3NItajFVaRTzgiap
c1gtQlyEM/PLorlITllKcLAukHRB/xvC5BAovLKuK7Xv2cUBR+Jddr79GuNQseoA
G8x4QT1HNAoEgLbLMxtDxySc6J2cUVKWog700qLSrprIUtLZrOmHuVjvZ291rv+S
BPEiYHUars/H4WVy2TjEPo7RJZaWmxybZT8vh7zeam6Q47Y4jXd4WPYdI3uP/OC6
0yzm6+JKNP+emUdXW5igI7cesfx4SNMwvd9EfnAGpFgVP38hxcZLXdptEyAWup87
KIoTlIfNSUb+miGYDewq2mNd1M1B9m8QoRkxrgimZ93GMWBCL1FicFJHb9kdN+s6
ADWPmgcmMUZQ/NeiUxOlp3fAnXuEGbdrWjqrUBtkzeGpJLpxTxKG6IPLirTTjK0C
h2mSym2OWszdnhE0eqaLFPz3xySWnOvL1ASOGHqFh2tqFn8IDE/Wwa9MBZ7fhSe4
iIOpOG7pYJg7HHk7jAsZPukZ9jgjHezoAmoDVQk0LzQd3nAfQN45t3u5CH1Tuhbr
QNct3ywc2f8cwET03qXuoPQQkUd2BB//IzHozJJUiogmfMd245GSLUOlqhk0xYrE
sWQ6hfLnV+hyoYA+WqcQscVuAxc6PP4UuGLqDj+9GhgNbR6kVOFSUswW77sY9Sz/
YJE8ZMGbw6x0NQv1GiaV+EH7YVc8BjAmh0sgTRTUXLz29fAcfzJkARLgKE/8vbwJ
Fp4qsg4e1cU2GtHuiiVrb01MFAGuYOZKBjT7CdGqO3GxddtPMmXAhYbYJtNQnJMv
h+RFDCQHN91w2301nbadmLU3tZozim1Q0TG/A6Brr2fAVYl3InsuUzR13mvrK4CD
6xbtiUQsivl31rvjnHcWjXkypLVcljjBo+0nekHM9+WeEfRLBXQxYUyhvIm4woUG
ALXD2tsQG445bB91HrvFvRqwifBkTbjyRQ2LPApSm7kAZMwHf2Bj91mJ+4XZ1/vI
/+MrbbHMh1tj1WOPGUC5jmmXSQfu8z8XZ77myUQ8kttqOvXayEQ1kos0rJaVJPRv
HLnv+911Ck8ZvGhNZgJ1+ALU7um7uuEFR9Fe8EO0HcAD35GooOahCiR3LzwEoh4Y
mgJBwXfoicmKuwT6YPlK3yYD9O4gwSOFhM5K1jG5w+OtmgbbvhrHS3RI6hXO7oPA
/fjObZENqnVogT+O3RO2comkjXjg7GSrLccUJHQLXm5L8sa7ZE5UVPdzeXn738h8
/SogdUZ6CrqTMsDhxbf6PGakDiTyFwqtxS3nJvjvmEv1/9Oe0ZR5N8xOI+IQrp8Z
ZHe28xIE7HFjgX+LWKGC2HNNC+VRFkaHp5RyiW7Px4mf84THdqrzPn6vYPQrpgYR
7fMkQcV/K/Nq53m36rzMPaN3NX+8EXYoJ86tD+DntAi1En2sn+GTM0ypKroeJuEs
8uwu3TqZHPMFSzGNTDSQD4X2v9kgfqxjvYRys4KJVFF/T4Q9/kj7HbQC0JUr3I9/
uK8eO+9dEyMMmGczJ6+T14UqBpRf+YF2K7GfcGEb8GaPtfW34/sG8DOc2bRYGBie
rDs6AQMw4bHv2mJGMxroC+MNDLoY3sMxmevlyPBJuXmbRHhsn6MC12XAB7Wvb0Gd
wRnO7hC+86z7wvBUjBqgzkwAWyhk2BpUTLF+ba3CWpINIMm7quDID7rG5r/fm/bv
MHnfQhcv+ksqG1DS5lNo5s3n/Cn8fDLVX1lXMi9y/rndc440wiO1t+duCNpaiUgf
LTiR3lR+PPneVZpLW7HcewXhOewlfcH20nYSwe1TKngHDRqtJ9/UUTpHrp3v2XGq
y1sPpkV/e/ZwBV55WqbvXssRiNSHkoElhBYebroevSRjxGpBDVbxu4GvJ+gcsTT9
vQV9ltmyd/nj0/mh5s86rbFlfYvamRy1W1KjXzpkRsYwpj8XeEmjT1y6W7JP3Fe2
1aM/5ptgk0NvP652vLGLNWIzDEQNg5P/YYzAndIJApvwYw0oYY3AhjYwpiqw0lfF
xCuq7Axi6C1E2DaVjEQ1P5dX7mLqUt63UoaMr1bqMV+HlYQ+/DKm2AaX0KOtN1Hh
QfwSjsJaR3fa6cJ1cvqQY2loh6R6/8JGfpNTsJHuXkdk4WrC5qZND5Hags69ZN5t
URM2VMImwDFViLraLJTjRAgTZePZFenTesqWGh353Dc/cMo6DDzHWuzP41lkfCcU
X9kqcW1/Giwp5x7vRY2h0uG+LCJpVlwmYxj2ZfXT/TU8skwiPWZ5wVOrXGx8Gtqj
eh1r7Ms1q15dLVfjw3cV6Y815rRtrBlTlQAII5Vfgski8T/B8xCWdRssyQleJIIQ
1Mv4jUsPcBTSXvjS3fIVppiINJ12dTiqlXLvk25eJspM3bEzJoPdDeM6V7xBZ+gb
lfNcihgp/AkyYEQT7Ui6tkAbCV1UdhVUrxf4dAACeo6od5PaRKQ/ENONlUNM3xvu
C+DAwzZwkkpoRIU2oyC8Y2Dfyro6cP1pddwanzYZehSqgnwJPHfc3CCkeVtatoIQ
qU9SxS6LUOAqlulqMZTPv17+Hta/NcIS4ikdrcCR3lUZ6ENUx6dbhUDpOpHqJ4X1
cnxlBFIoNDZAI9zzFi9cqwU/HZt5z/BoxaXBTdUZEtFl+JckFGSHJPglOD/giwvs
GmhFADjsr2MMCe1fklhxwYOWhm7suNGjRlMIQISvN3BwqqVINhJmeUVT67HP9AhM
vgB1c+nPCHctZuSY1WxPFsxI6FYmL2gBeb05IZcXuo7d+TMOrC0eCfs/MVZNs7sH
ixF2nxFw8tGtmOebia18mZW7qg+dbWcd/ioC7tlJf/jD01A9suC0ohVwmu1alRyw
gE9GNwCPNDnz+ja7yIhN3RB+kNZ8HsM3tofh0U/2O6aC51lkHV2se50dVAQmJkeM
9ZFGbS8QzXd0HpvVzOBsxfAiuG8XUNYmSVkqJDgMsWVoykGDbiyMjuM9GfUpqBoG
s6BrHoUq4vkrr/BSriyW1Ck6UDBLU8fOX9w9KCGUZETgHzG2pWl2fFv0dQc/r30P
RV6cHNTtpTIJ6pLPf1qLhCv+k94r3U0MOhtXKR075NeCyNButV8LHj+TlMf2d7Ls
k+Pfmp9dAImd9pmZeZYyQmTHwHQrI7fhktV0EgcNCYd+T3H5/ML+8vJbZvvYoNV0
nxcVA24qv4qeozVCUbGieNpOpqVg3kVJIQV+G7XV+4dki90D9mKyqG/Ft7gtxdVW
wJoJAbMOPxQ1xwl8he2jPe6VLHB7YrAKVuc/egeL3Cq1ePzJDa6V2edyQu26b7v+
iGTUmsPuF4ZqvLJLudeMB1GD9ZHr1Z53LnTmluqnYx6gdg5w0xvA0cSUPnmHu9Wq
mY1H6Ee4MwwGCXl6I4zFfvgF9xW8MwPjzk+Fh11AItjo2KTO7329mWDh82v78Php
UKK+aF6Aig2rAcqunUPMq+QB0VbtK/1pPjoL72Qjyel4nqardET2wjg41OUz3aZ/
FPxh6aJxzos0yQUqhjPtoP5okbBZ1t66yDT3b6o9AAEU1lq97evSXw1JxOm7VZ7g
EunpW9kalyYVx/zjkujcVfYXVlIAekZ82M5TCNSqji7sx19zWi2a4B/xRrhThpF7
RrdA/bAOTRP7dUPD4692arQoilLUUF4wfxEoG7mxnaOEQvatPVhc5ez57t8Mi6N5
OzYTxNJ62A8saFthCsYCGUldp858HZSge04SaOBFhL43IhUNBMlz2CIBhzR+kY2p
1AQuia6aGQPCg5TzrEQtb/PGnQJHiMyaPZBJPChYtKu36N2j2+//HBE7Kjxm3GEt
fODr5+Eab3DznToRmZcwv/Kt7pF8K+nxonCzJUJAHC1lzAg90bxZ8TQ8Xcm6bBIX
6lw7uMwvufbuV+EVexclAHUqrVYaj6ZoMmJAcRdTJKKIaD3Dhb2zpNiP1c0F5RcU
+WM3SDFR4y+7wbGAnqRM91SCcJfkxWuMlGHyD/pNhfZypPcrH+a6XqjXuvrAZF/c
5B4kqZ7gHdLFg69feVOInL9Pfh1xA+ONfujDa399lSAX0LPmUZgxXg0KCNRZ+A/z
vPcMe3UpqNU7uAyusRQNYJ357F52zzSMSOJLokCA3n2YK71ODqdVotGy894igWPO
0adhjGfbWXq9L6/j/RyJ96uZEARqKiNt2cJT8/QvwQdTarawE/LIawzSkI4tHTYN
F+FyCTzezL3hFcb8OXLZ20iP2aYWIFyJzIHch0uBgI/QML22FJepK5EtZqmPb7qk
QL+drTB0y7yuC+8JN8j5Yi1YRyTYA1+BfoDrhbE8elnJOOGhJzur96wVTO6eRGFV
64pfESVTz5zZ2CQKMaGZzYbyyPrWo4blQvqNBjd9VkSFrMwyebL0t1sxxuUSZiBn
gCMiPKY5Zg71pq7fMazIKUXKNN805D2qdy+vR9CIurSNQ+F+D+KlWZYej67lY2Z7
VVDDJ3orWV1tuxuEnInKP/G/SYi9dZjjrtXr93z4/cm0IaICGedmp5o5x2oLjJ7f
LIZC1AZHS4H752jUlhDbeKV7wrzrExEwLzqHKjrFmI8BpFyDjUmvx8X6392ID4O5
uVaHaaPJdbRn4PHeKAOprOMDejl8h1ZeObkJpW8uQfL7w9OCNxoiFOkrFkekw16Z
C9KisqLDZA2noYIRnNnLCMPWgh/mXWRLkn2LjmYU+WvOgyGlImjOrTo1LFKjCuKn
GwhiGYuC0BU7ATBAXSpjXIaBPsT5/Eaoi4kBhwF3S9/fn8GhEgD0HBp5CyMV00fS
+GNqsjlM469c+oD9UPTrftIvUonxJawGzCEMW2keQC9blFTNZFIOggo4/+24Vunm
wrMHt38m0VDoYHNellRm4kRF24AK8KqdR8oBnNOWoNdudwsfZl1mqsuKP7Dk/J9f
9GWccR9bABCnP5Mu7sD2Bp9HBBZkGJEBWzaPR0EhMXob1BB7AthEbWexN9Gcoolv
HIYn5xtGkCo5LdZDPcLJ2MZmomp5DUjlY7ZIAnYOsKhc+niaJxDs8mez/eW5xa22
0OSaS5MxgKKiaT5CK8h9qF2Cc/A1LanPKi1yirBjkKmlcY5AI++maiuuG/TsMqSd
p7qGgVi6O1hLZwPHiX0NGQuavwYdJ4jEvB3M/bqTeY/BiFfC6JA2vkGFJi9/XrlU
qEWjTCO0hiqpDX89b4idoBdvZUs/hyyj2gwrtsrGsUfguMlJVA98MzJzkN0YO0kA
9icyzH0MqaNCQujWDr+aadE6JcwQhXUuG6ZezJcVaKi0UX8ySWy6dirIYFZGS7Q8
5xezl09o19EpjKSzCf7Fab+eNnxBatPpG29aQqVWaUnEj+IhA7loS3OugtrTL9Di
4wrD43Tqdsxdlakus5PLejj19IVptyUCDNIJkf0GX8/3c1VKsl6N/H5oF7QEa+et
kP6qyzCxR1YABCRsVEXydFRUcWNXtQ/0M2kojgdbjzB6H2Wpo8mxaejW8C3UUZ3m
ztsOSe8qZJOfs+mw1D3BHz6hSJfEmTJnGzsO1dA1ZOIk2buFkwpinRjLR9zUa169
BA19Dzxt8BojcTcXLt2+ty44ESOOPkPCvVS5NIhylYFAaKh3aIDQSwzhWoE4/pjn
kCG/QhZBdrhta+MlA6WvU/oO0OpoIDfT9Mzbg6+OHHdahZZGQXks9XTcUwFz+Szj
ZnLpcaeqQ1ZTgt7n3oBErg/bGnGJ9EOX0IPmxoFMqqpR4NFZRtxd9Px6qZe+Phrj
9noJD/LImQgl6/2nkLgyjq66P1Wz3vTQ8dv5mpZ2jrMm7DML6O6KY8GAa6azFcnQ
1OiKyf0KYztBCmMnT/Fk543IBzCNV0l2fFMRGlptb42LvmjXE8CuzvljhxdZhBBI
YvQNpOswsTuKMtuEKfCHOThXeWBXKvz79BZKn4CBbvo2em5ob30sIT9OJ6I5c/N2
tLsVwKvfhmsQ389qSwvzvuNip/XFhgtq7e7uH7MiwKFFFXxS4J+XWdNQqsEDh4hj
80Z43sVGL4D3M65yJOhHUanGF9h8dU9nhP1MWSodA/AiTmOKz+Z6nk7Cem7DUTiR
BB7DEnMItIVKwnk/0pPncP9FHsZlabBoy13/YffikZyRKVbRS55PRmOMDL9ru9hN
uTy0Jfz5BcoykNEUNfULqD6lvlAnqo6eUe7mFmCf2z1IYPhku/g5l8KyAt9gmHHL
0F3nUFPnyCVRn0PvFfaqJ0GBkOolzAsZrpCPIxr/zfZxpmqkOHN/1fyJrSygHxgU
NcckJBxvk1M9hEWAlpXPt9Q2pAIp8RYgmVoyP63WnmM7PN5R80X6FdP82aCiLxyT
mHGEH3tnmcjjfp+z+HhXYPl1iLOAJnvzdbZilth7Byr4UVKwXMsZZy2Nw2mDSuA5
9pdT6LRm/Vk0m2ne/wubcwu/ZXO7pIHZPQf+KK5GVscc2VDnjJ4jqm6Tv0YEWRPU
NfgxM7fbDupDtgCNI/7PxEy6oUiJxAB26TAqUSWdgMhpdXio/fUJa+C3u1tuZT0N
bbsPTgjOPY4ZkiG9pAr3zAI9tI+kPO3p41D2fvuxKHM+6ZNZy7/FowtNdMx/XyTk
ZIr4bwvI2GDY0DK/05+5zOsFNb9cjEIC863LLvgvLscOHmiDldC9smg+mBDnu1e5
3h93y6dEgrrKLEs+wUhsNpNVFtcXgZEC2bk6LrBxxmMnPF/nTZwm/YgO9hIwSbhe
KlhX29dldC3YX4cFPbwM6jGsrKLTZEc5QHNjzkC3nVjnNjAtkfN9YPWQq47FsfiW
dBDa/vfnsE53YKPIMQN1hOTko+qSMY39qDjbBoiHoQfJ7HRfBrcFq7DBtVRpmH0P
MiaSu7IEqQqmCuN5xrKeDswn8k+0OfAejF8Jnm4A/OQJyVILgO5/OKR3O7zU0epZ
3xKLJFeBPbVYtPpJjCp/foA/qRnNLYp9aqEQ3eabO6hGtzl31cf8GhSlNSnMtQ/w
YPjs4PEPSisk3HXWsmVaBJW7O6a4Kr1ZCJyxZehyzAbXN/ps0l5NSNrW/rCdQE5S
tSDBlsJ8LqEu7lM1Y0AAIc4lxLzDZ+YSSPdERo5XlQpKPFCAdN3Z+J5CK34EG2mk
PnavWoLPe9pr96srZ65t0NSRALJUVZhZqTQMJMQ5VjrvXmMyd0Nzn0sLAlLLMfAy
FmPgAsv0CLSD1cHHTjmeJvFVvUyM05GGIpMAeW2bFwdz7G2U3Cm42aiwJ/JjI5P9
AK2ZCDpBPKE9QaiB+GSaO10utsOHRuMdt+C4/3veOGg5hAmyPLlauNIYasBAMIpe
LIYBAytmZ/DOJEJy2MoygbDMP57DacbR/stSmEM14lA0DVg5Cs9QMMGXCVGO94Jw
dezC9ZtBJicIZK2d7kcJERJEM/zcnuFn7YO2yk1W7fWnjgK22ru/k9BJ+9eYWVsa
yrNOPbrJ5Tew5tK5SKR/VC0ltMSYeYLh5paPFSvLdOCFUroZvqIOy5ZOphAnGHP8
xN+AT76/0EunFoRTP98ZMFAH4N2JomiFrIidIOXFb5deyYoc2GpxsHwAZSnrDPwQ
RvCUMmBL3RU7j3Stj5ZX2xIe/NrXjhvN/GUIyrsWUlmrrnZhCwMwJUsR8iNfaq1w
Lc1XG7UiP9hj0qngoxiSfWc4+X1C2UpovZJ5qi4ZFFFLcukCDKK4L6yxqsCkiTHW
KM+7sEZavIKHKyIpkAyTR681gRuffd5o0UG4fRBisuF83304gDm4QP20NkCctzYk
vflwysse7nac2PQC5E9Ok2t2kg23PedwliwjWL5MBXKd4PFhXkxIE/++ce0/icK8
rR1CwS5h3GC67LTUf2f0EZtqdVgSiBt8Eyex3qfKVnCCAlDcvA9IXGYCLQyB4y88
vhGOmbHQtu/lqjIlKMgxZtAwFNJzkyV49PXTIIp6HKZCpSty0sddTj+yNjaC+2ri
qRFZ3STMhq5NiWnnrKpt9XiSM5gStwDfyzN960NalEHReAkYThLfLUW/alOYAadm
iV1xx6Z6+DSVdKJFdfio/Yk4sqmJhY3FMwmzRFGrdeUqOOmu0cXEe4cc1Awy8uGP
pbFqxZmjrwhytw/OCPRvoM+IgqJE3E/QgIEVInYtlB4UGJSqXajJY6MTzxaRfIyP
NwZbMJ/nd+ZJnZLmUh3TfYoYZ8Je5mIKTSzbq3On+x4xUoV/dHlyfWpPL3t14S9c
8CRR8N0zqm1fnUxc23is3DA4KVGNBMlKHFFrQBKQpk4LZHaQm7TrLr8hTLMKH8dF
vO2DZuCZySipEk7agOprp7z66KIPGgAGfBUB7WrrKYgEJqZT6bxuh0nyW7F1jUXR
ov7HyFMPtesHVfVd+4NBwagKIaoQ7Nsx3nt6WYDOBzJVB6rGuT9rqCqlTqzvPlRg
glt1ab6KMnqnN1REHzTlJ4of7ymcxP6WqBskxbDPLTqzU2N2f5x1niebuLKBd5Xf
UG+iocCjn9DRoSNoI7r5Q35K5HiGgPJoNdRqyQ0Hcf/3IAnvqcKnoIOFHawduEXH
SJoy3ritD+YX5Sghv34SglaIy63IYk8Ge55/QSguiAjy/3N3ukKUFXCybFvZiGFw
dU6aRpAOmhhZYD2OXBl8AA1397JRagy2HJwiTo0JhzhTSJHsAkK+2FI7270YWqPn
h0EfHwYnK9zJCNMldltIfa0dUD4bw2njw2lrDVgrnKvOh+Bta9Fgk82aStqXdPiV
xi+Om2Z0PNAqbiCfo2Pq7FHf1G5XCYL5n4uXOvTeE4JJvcgxxkdGdM98buNuiqAx
Ly8D+qXq4qwKvy2WzVnIgos77U/mNbXRLJrmfoX1xWiTLj1RlPGE2P6eeFRIpsKq
Lrmbq7QWuLUeg3zHW8+1LsghYRNpuBVQjRYCcie5wE64nHShTaPnBu2ZkYf3a4BW
K+l8gaMEGFqQCD9JYLuR/7EbtXNRfc49+6EUQgkYgDJcMtwMh+Oex4LPWCbO1ai8
hMCul5ddjQE+rP1ORnzj7u6zC1mK71L++ibvVHJ3XvJdLLvGChDxzpqHJATZxOlY
hxojSlv6XPm67y9QBEmTQvSUCenFCyVxumk4+mjon7rztzwJf/wi8v+LObz/e6w+
65PUzaODJp4P2JVAZpxGL/iBw+kMKMB22OkhlTF4YfLe9oBHZFPfeRGlnEbTJOKa
Ol1r1pwkmZ8050zc3BYkSvnQGr492m0n+P6WWAkVkhOhAX9cUOqlwL1gFGUxQynG
d10dApbskRM/s5T7hS83KvZDucKWt5WqtI83Ae5/zlRP8PvGGZuxSFDtTDOM+N35
HVMbfChLPPJlVbc8W7t7XMwkjDT9WYAmMz0RhQ7mNWKZwuWVv1FDZvZujEKXPuJi
ChAacE6mh5laZp+6OrWpdbD6l49Ndok9009s/pM2NKsNE0VjK+D+sUySiW1RwY2/
beikg4urYiIlBMPTLPZ0BMBirP5Y0vkbtP3hUSUqvN4lI/2YCktMSIIX1Bq+FgvB
CBL7GVE0ZaaL/lCRgFZSq40Y78FUks4dLh7RcpPYr1GSMCEO31e7Rn6AZEdwNkw6
Mj/L8PgKaIgYAq4n8RE7J0j7UB8BRFm052niIhbtfDMcBqyUojYnJjCCCU3s6ysG
l23hPsC1OdFjBIXEo/sfQ+m+wf0XbyF1/rk87ShBa5bm3iC/9yWMtpIqiCqiAunV
yIMzYwx7pH1ZYd4RcaFnnMPBQbHLPUwVZL/PK1W46RQJZDbqMx+oBCfIf69pm1te
dZv5PkNQY/pDQ4YkGNpLYKjPpy6+dd+LkdsgBwuJgNAHivnYAE73mxF4dj+wTOOb
ODd2Da2fgk5gr2qVPf53wwwcOB1keJDCAKp9ZPIIgI76LQN4rjJSaR5F+8QwY298
s/e2Xh59uop0r+BukcZnfQqisYqYbKPmPoI9539atT4QkkrR9A58cwJRKk4R/KgM
rPYPh4zoNvj0b1jB6vY+tSmWfljDe9aBt53IK9J5qqYcO79r4bwaVxL9s3hP+gLp
vJAVOn4t5KuTYh0AxkrxMErmPCDL6GsXRfcyHNUMRip9wir3O4qHFAfLEeNHAjx7
dxv6zABOWQgguw+uDnWaxuXlUbJfHCKMSXP84jaSYFuSvpiQzFyWOty2gNbrGffE
0BLX4B9q6vJSIo5SrvohebqOl0tRwaqVhOh+tgUK8n4F5gfVvejrC3t+v0yksMxV
PXNbySYLpi2STbjEs77DIka9KoqrszQtjyhMYRo8+3ViDw2s+6iTThiJdesaLXqj
QxVd1FnkuWa8WKzkm75lzVppAvv+RyeuIfdFiESrkbRXsewvFAS1eWG8ts2zQOJL
JiEGqU+cxa+Ctk+clpv3nQ+qyfLdzvRlpZAFc7h0MNhMNGqtHkSoAy6/YquqHHX4
8xVvOUciFWU/VpFjO/RlrVt1mWY3ep6Djk0TsxqM2HdRJZwJ+PsaSvIsWqk0R+Ed
1gSD3RKOVXNjMwDlzXD7FnAvyawa1t9LDjwbOlaIk3zeJVm7jbESuANxtv3N+Z3f
eyA2Q6AkGC21XodkRatWr8Qk0o9qU/AKKNu0ZyVVB/V+S3/Fi/mtMqsHp+bAGGAy
O/3vA22ZGw39Zld2CidbACdazxo5NU2UOffiU+ucLjtLO7D5tBZ/YpuHhExEAdJs
OP/bym+h6R/jAM+m6gVVBtyLWVrjEMLNKo9o0MTETyAK3cmKuGgKhUvEmYP1G7vJ
kKTIN9wyUq03gcgH5Rld/EJErcyJaZJdOE2iDpAP/JFZhTNdmbrxHLvrah6VcQtl
Myq2jfeHmdMUhQVyT46V5gPbuwR/369YzGNHVLJ9n7/O0LjryNl8GHDVZB3JSjNT
iBY6mPrmJsMPmr0i1lpZ7dpUW7KJd6czAIVs0UF/naHceTBrRhIbcSQ4MDDwE5yk
eVUT/8PfUbocb5g6PHuEpwx+EXpls0cyHcccVGxEQ+D7/EOhjvp+86bnft+LpHXN
48/7FDvBABUPCfqJH7XxxNGCjgBn5Lc83n8+dYeyUtgAgsDdAA0fIusht/DXRv1z
O5qAzj/V/6+noXpnXK1r7YUW04HT1QPTS0RADNhmB+6pORhtpe85BlHJKWqWK3Ze
QBrB0bY7mvQdgH0aAXdImzWbKlWXCix5malHYBQ31ApuUQxbtnq83cXHU/TrEGIn
lQ9V+x+d66Eubxv6/1gGQkyzd5h21ImkeQa8AsKaWSIwPDQHmacgFN7YJv4LBUF6
IEO9gQIuiD1giV23rIOPO5MhX6Jd7PF5pjxrhFYUJYKdAjSxo7/ifGw+x8/HNXlQ
zymlOp0/wAIA1b5iGFleuy0rAlGk+0NfN5PVyrQDyD2KH54hUt4QjhB8H9HazTGk
x8WtED3hUIryHly3pyWp9ay/ZpffOHTfXOxeujuRVJj9RP2OWQ0ByIqaAlOOP5in
GtiA77TTWk8I+0sglkkU6tJyWyGXuFkzcJlprlcErGRD1Q2CS8TnCvPj896nQ+iX
QqCTvA/4idJkWBbCX5ktnnZYVB7O/AOYZvlxC2CEEwWkzS13RmQ/F/8hGC/Sq269
q1h1eId/0Lo0fHCICGdZM/bLS4EE6DkbLjDAoi0Ab0zDVcJoN5phzqvfs6WswKAm
9EER29UXVqlHyUW0b+u1/dSAyXTwB23h8larpERIP1e1i4guuF8QP/LoWOdeBzFH
uZEiqbQl3mHiR7YUKAJMl3kO1dV5xY2hyaFxzB9DHAwo86CLD0/SdPOFdDQaxWZK
dSLC6tJLpVV0SFNbRLzbEzsx84lERXGayrCVPAfaHF7braxrDh8Rhy0XMfT012l/
ZSHwjw1tyTRYStBeVaFSoH0XdrIPu+DJTemL4JmoIS2UyNEi47cFfCaJc3Yb/+BV
1D5W1qt8et++D9p9TYPMV3yBDbQV56wspRnOu25ztQS3vWfL8wnJPNsb4wCZ3tTn
jfHR+/gLVLgDQQsIIYe6SK8QrxoEy7hXqm53p9SHPDMtXmgO5pHyDg5lb7m+npYt
GBhrbg200TQ/8ic45zyBr2uoiPgefN3hY68xCCj7j2KfjQ7Qr+c4XQSqAkfkIay/
CAswgXWtqp/MLkLtlQLFL5hUqa8ga8bT+jvIzIJPeTvqPZmJ/wr8gVgNXAzvfo+q
MAhiukKqt5E9n+SfB8YpIQbp2/6V8+FGmhJiloGO6tkwyY1M9rQon/y8rFf6Lhbs
JMqOcd3lRZXp5PFfAtZXTGbfwF4if526rY6w93CIhYWcUtEgCepPAiprZuthjE06
egV4ENF8bX+PE7B0UEmMZU4Bv1Vw6n6eN0vzCja1s0gD66kLRR+oxwrPnukWf8EM
bpqqrOq5IeORPPAJLG+wN1zeoGLzHa+hXNO3dod5sqaJwXGAeURq//p6R4Lv2e2W
oxpQXEU85By2gmmJld/GFx0S/Zd68HIfYr0vLFm2FMmbkUI9MUDwqVjugM1b5ndv
hVwnswJ3UlJcx0WIc1+eIo4vE7umyGHO672a/P/NAzmU+zHohCBXEAWyXYZz3W47
Inqqfy1pYxKPDg2D/39gCzivIarfXgAmi8H1xFFlzwH2Z9lR5FOVZvOcYcHXKyXh
4WVuQF4ya1lWFUNg+/zqzJi611fAR8hSM+ZarRuTSidAuKKMhioIPqnQZkSLzeBH
dkmSMzDwT74hU+cHKsasDDhWacMbHmvqtnkv9ah/k0+Kk9IMv6qpQM9zseCCRYZO
H+4mCVFDyDw0XVDvbpTHzEkQPWcqf6SCVG1OrvSdADS4Cv/cdbP+UnPJkiUcH5Dx
hIMAMhjxdFmhNaVnrDrS6gB2OYywypqoZy9TTBUQbJ709WoaQr5HG/fGoOV+jK2F
gzS3So5RjXFwnlp4hV8RDhkN/gFvHZwknRr8s9LSg/gKPvlN91T2UnHmAJlZb+jk
da8bRPhGxruVOQQtmkeWJiFXqYqxxBUcusENiUX4B0P4tC6D2SfUl/zWQKnVOGX5
CtDmSATG80c98PZnteBnVXpU2FyX59V1QSuyfdeHZ3OOw6H9hPBxV6mVYRBzVUUJ
nNNoogLltfJEjJ51LqqNvLkHORc2N64j1qNPc7Vc0JJi5mv09Q9Whu39DS9lrhK0
LKNQ6P4bnJp6usvVn8rVjDInvQ0WTFSJ4y114WLR+axCeaUL81i+9V9QuCW4pyCK
k3Bop6VGBNL3YBdH2I2t4yMHeayqS6lYmvwCIWGdCOoE4w0GBUy6l7Adk5oYdBFP
RoZHTW1zks9hAAt4fknF6oZQ0QmbLgMmgEXGndNHXwKYr/+V2LcTbAAnjOcAOWED
eGf3gB/mmUV+FDXT8YyPn/dsaRs64dhvFfs/+KoNxT7YIphqIQGgkg3nCdF5nCw6
3DS+iSkjmDvh1U98pzhONg0T47QF8S7i2w/EkIuevulSFvd02kiGYTa79FE8MXoG
u1RWokw+BYjjwU85WttVPGUitbPPoCsM+h6vVJ/FsK40HIi6V9heHFzaIQSmamuT
vHwagGrEdGHYOse6i45Nw00hdOgeeDHOqV+p8qXapAXn2GB7P4uDnnZOklQls+zL
LMKzMboWLWJS3IxBXCUyZjA35sDNddcSh8hMolZQ28MZ4WicfD0VcM8Hq3MCoQZY
fRD6zwSs7XSocffeKgftpOc52IBTIFEtZkxA2z+nzVc6+9A99pitjEi0qqNxDdp8
ejJS/RVaYPy5fqvyqD/7+QZdDckiUYwwQ68uRGwiR4Y5LlVdnWYl1f7n+DJyYzlr
Mp6rSbqmsRma72sEywyRoxK8B3Uj/+7xagI52Dp8/soiuo57sjML4jUg5DvXpk95
bMheYVDs75nHm7IZ3VuFg44VrCY9WxtwQD/3vLktvhYaOxJO9tJih0DgOtVKFhfm
lfuLdgywZP2WSF8ZsiM07wYJEP/K9IryYaeF0yXiJ224thbH5InSL4akwgf50WkX
HLqEmB/+dvKjf4NzOvtkN10jNlYJzfvhwf+4DrrJ4QMG9aJdP8h3nXyp69jzaiJe
fuH8EEZoxoRSVNwhg0DoAiBPesj/tTGgU9A1/PbUtru6IryCSQfaylxzYJAjpsjs
pAE7S+tWZDUPiBd4XC2d3/LFCOrxxPq+Fz3Ateekph/cMAKR+HPj8ndXo2xd9j7u
SorhmQiiHo47e1w5SzebR9jbvr4leud5JB4y+S58n/7k4ysYPgKH9XiJ/H8RA52h
xhFeZz0t3fmwMDEkoe5Mq+ad+ZSU39G7l02rqMgOvbXHgDA7vz2wlxqGBvUAVWyx
JigMytbVHKUUXAM28PrPVPe0uk7ly0nuGR/cPfNLHvyZmvdFjy3oLmOvUoskwnHl
VFCAg8rCeIR+FJbkzBUOEa/fc5h47kIPt9rmR16i7Xcfwb3zlVEVwosdceB4//eZ
WbU9Rkf+UcWvTvoi5YULbjeEPs/i3b3r8fe+AFHBZQhTF19tKAwo9EYeBpx8cNsW
c145HmQRWhCQ346JGqrjKqf9dWVSZp+oBMArL0XWehHtF6Y5Rfb2unhGv3FUBoM+
ot2iH/uP7V7sNp6AakWGvVeDXpID1+5wbAU2yWpu2sNQp91Nd9/J1fdusTdAzyv+
+N3+wr8uN/dIzUnBwV8iDZvE6dRlnoAYTvvSgY75/dei9wxMwyU6Sl/NXIZkXIqu
bqTR2YcA6gl8jl9T9gL0sXQoaA94a2ESIt6R0WdphMt93qLoVIAymvEaaoKP1tzj
IDWLEKUk0KJeT9w+fehI9lp+d7rPNw1cQ/0hD6R/G5EMaMveM9axDkwsXbtL1Jxp
497OjSd1bwIJkBa/HexLeyuSJnMVt/tUdk4fCemIrD/ld7LEPuYuHxkcN25vKFWS
TxUhG/o3os6GZX7vwGGhmlruPqFTwJhRsFKm+WMpUk2s89jQcmP5uUqbo6JmUj6N
sAJK0dsEamAkqcz3VxZD1vPNiK44lqmJKq9a3cVrRX3J5vwcIU40tEK5mwXYttNm
LIVp/OVfJq73cLLtnJLHW83SIdGFdqUZs6yxg386h23vAhO4D0Vo5i4e3owTBN5l
0kzCK2qAdblVd/V/Okx+yqsmafYoeUqkz/4HTmPKVtCsOx+IF2TDlBgrZADpwm7Z
S6MUGsMoQ3nfIrdwnbttU/apxb6ZfdhXAhBRJZDWica6c8LnKX9G7LaFB3vPfRPz
V8uM1CvXiQAbDQxoRnhLkcJXrNdYx3s9z2CcnMvp0qJKHgGHGItDCzf4/jHJ7XFq
Nxs0nX+FcNxbBhY133WXjFZ6EiWW6cuSlCagZaYQ2QdH6AK8PrdxaFag+MpWw50Z
ZhISolMgeZwDNa5HgNhxSdnukmfXwu4v1t1/xj9leGybJeTc/6qvl+HEteblA7SA
HVo7hkpfFTPFUwtYsJw3vyVFyDeC1uycpROVMIbj6ZZUuNnt0UsnPctRORoiS61f
q+SLSQNa2WkIoSxnQmdnjnlwE6fzariFoNGmzYLXGF+nhsPUToAl4qb1+8NsJPFQ
2GfY9rnC6Nm7oN2TWDX6b3hD8cBqMRj9m504WB7RIICq+artVd6TI9twfcKmYXWV
R4oJ2g4p3F7alFSZsvshQwoZFO2Mc18K5b61EYKpy6WhwXBaWURVO0iB/HFjmVej
fT/5kG6JtoG4cBSOpcxQo7o5BCPK3+kiakTfv6v7d4o8Z7QaftIy6yiLO/XrdOOU
MCKII577Ot6SouyBvmCcxAucmptV7dOWq9hRQFoL0YvlgPKi6dnFEEzTUDOXLek/
TzAn+EbIavN6vOjGgBO1kldn/+JOoE8/XnBaCJP3gKyW9+WHP0GzSjfV7+/INFgP
bvrH8ZtUFTWwmpjYjJRusxIW942wFXUOJUfrs56p4BOUAYNiXG5/3a9LObZ8UNMv
2DO4dwavhPM2M34P4LiNSbWVbjytyUsxqbVmRzRIVI8/qgKXfycajgq6d7JkUW98
8pR0gpWteMi3ooNT7OVD/dZkmHmkfBAWneRUN+u+TqzrBR7pVNjnwxErUMGLUZ4t
RQJ5X7QGmUTzqzvudB65rLOsbxrH/xKClVrjKNiSReLlr9UvqrTrCgpMHZr7Wk/f
KrL1MQDVhXf3opmFHlKAja2zq3l/chpBJO7ovtgKc1UVFt6qTng+o/3rb1d3Qp3P
nRrtZRkJJ7i1/Ebg4YUMJ1ImoQJ24KJja7tDVZMOSphZpBj6OCtpqg9Loew+rBiQ
h4gAMgKL7DACnAb58ikukh6fHcsR4Yue2UsVAPtKWsUdEnGG6wEcISvZlyU1QnB7
mH30++UO/aIhbSZNV4zXvzV0bFA7UzgOw9M7uEHvgxlsHMQnSYbjkKiLxZS8tdeA
/nzGQ1MdvBcSkNQUjlRtza+tYifM+n65LJ/g+32nz0QSnfLBmO1X3e/BqzfBAN2N
qhG5YCcAk/NX0yGKdAHnmUzpLwUbNrTH7UvToyQf2UB5ddSLLcKnfF2Erz1NAvzW
NDIUkaojy5jbdPDBVYgIcDD7WQKki3Rqmu+iRykrdewllx1RUg16fGNl2LDQmDXO
BS1GFXqDOAsWJFDXk1V1jGEd28ssq3gr22oXv0D3UxjR8kzC3DZn1wHh0FQ4YU5Y
sMTI/8/xR+w1k76Pdr2hqmLziW9FT322zH7F0X9Kxy3O+8qfrGc1VXO44BEXH6yR
mo5MBz9tUM7ziBZ92ZvedfybbtzVelfXHOEjlJD81fkWF+ZLY3ZUurPJkpF7Pp8x
SZ/zMp4IheukrBJx13jjvC6jLwBijIt2C5DSF+goSrJK8BqTSvbsJynzjO7NFE8p
O86SUC392M1AXtu7GIrMAcmFc61xAUNhaeYQwLhgf7uZyCorwi0gpQ7adnPTFo7G
rL9aXF72slhqClSusCitlhZEOYbIHnlxjphI4l3MUiSgr0nVKYAKspHXKQEDMqIx
S+/q9bdEqqOnf577K83Cc/ISujScXLqpM5sOn1HejPvp3RgHUgw8nhqGMzJxZ9VW
TdApBGrDtp0u6BPShq4Npax+F8xaF7ZKWgDkI4nBjM/1x0wPbPRCD7rgMyj1HBHZ
ni/oaCxxyTheP7VzSiEY5xFBWebZSm5nJ8ifGFdPgJiWlP1ynunEQ0fy5YdjrSTF
zAvToakceAzSjzyWevHDUIDO94phHqYqeJnzEVzG4aqUZNfu5qeZIczpFJfzzRtq
Zq9f3aLorDfEsXNCclVWpLxDc6L4xXlhlKgmHG091L5b6VVA2TGT0BGH9+jWVokE
8XJPcFLU1UYkoxa1Wb+0mdvSn1FquCR6N3JAYEEhtEmS6sS9h6ts4x7C1Qb1Gl0K
Ruj7vN211eMs6krQ9bMCPQKpml0WrKUFreczB22Y/VxJfL8EMf6s87OR3bPyVOvt
vp7XuVGCadCb1CEbS2sbUVr4Deip83z8za4cFeK141v7ZSsGxQVJqFHJ3DUaPA20
vTg2qsajJ5RjgKYMliehaRa2ptGuU2LClVw6Mx1kNNxQeTKHY3AmdlQ9orm//FpU
0o4oNdNteUCWq9CXt45KckHTXue3uf6+SqUKfwVBd7mcO6OsXy0GWNa4+HbpSTjW
gKKsKy9/DEXU0gPRANXwVl8xoFoxfXomSaLy/bMAjBJXLEtl++hvpkJ28AOIM2bi
5F5RzF9j3GBWl/eFRW4zIfkIvd2HP/JYyqTO/hbnetmtzzl52MplH+GL0xCv1m2x
7XGWiqtBxPDsaGGIH0pr9czDUi2fagy/dkOeyIR0i0Kzu0QQQAKWR65sKNETj6/E
TxRhDThClrsKkkMgynBtqntH3lo47OFLV7RNwuJ1OkLwkGUySGaxNyuEeu28jYtk
AxTxazPUPWsg5u4Gh4HxGBmd2/0hHOrbpaN2IMomFQXRnepe3sNLu4AuT0Al5VUd
aTWcmM6elaNiZrjk+gIUOTV6WKQbDJTS/B1PWzxH7MNl6xr4tzfeBLiB3dWeRsLp
q35DP38tTnq8kUdj0bc5NkHfOFht5fFTqZSNItg6XdvYkXJF/q0gs6C0/EqZbxV1
xBmYioClcfU+U2nG33flvxA1tGxwNwnjHtWQ18My6o6H5OxLNyZ7T7ua5wXLaprf
sIKkGIRSsklrGIt5yZbBwhjfcl24d1iCZMiUsEz9+tid3CPgBlZymOYcOkU0dQcs
RK2FeuO74tGQ6sbLNj6l/mCXb0aQE+sZ0jEKAqb4kXlis7RwR7QuSbvFJFR5k+5y
wFGQFMKAFQ6yS/OfNkluft2dHUOwoVQew/9KxsoJDe9y/l931btg8yJgDW3WdR05
uswVvOriHrtbQibz24+Rwzo7KwX+s0WlR/nZaIaNQ/5oRzCp0vP4W+V0OGTe4jW1
mlnQDJzxx+pLXS4mm9CkBslOcBC0dNIO70SG/KwN9LtDeYbF8wqC5faN8WNmRPdb
ejseg6Ig3qO5QW1fDvgV3pf1voGIW1IrHByTmAWeMnF3fYBnX5ewXRGb5GoJ194R
768f4B5HCOf79IcgzkUBXh0QhYGJTOFxSnonUG+Efj9gvjXP5JFXB15e0Elp4cRl
AC/i+4PNWs07vEn0g7hgBc4se6UqeJA5+yYLww62AtxaQ62Skaq0RQsn9sJMFyYE
6Bg6uDHJnf/wnkiUF31rFIq+Vpn/h6y/jY2Jy1acHfbervqK8y8LekAFEdcKLOh+
LBJ1p5c8jKz3eWg6nBeFrRfAaGYqVVOKyXbvsRV5kIpb/8zHU4cdyq6lUKyaPoXO
3wgGYOgsXH75PjWqgELr16KqFTCHb2vTlBcaUaZcYwLdtJjZGzuhOMu8c4B+axrH
H96Isj05FY2vRlbIJEQiIWWRBTda6Px/APLICUCVJPRH5pm+fOfbylOs59NkSyLf
mhES+mWrVEvGxCzz+C+/HTOmZwiR6SShoeCXTJM/DJbCIGnD0N0iAF2GkJmxfVra
Rb7vgdIurHj3rPpaM+I7BPTMDK2mEa/WQjp2ChSXuErdAcLl3n4lKjxA0iPcrmeZ
BqKNiLcd+ExK7jLes4LHMEcJB5zj8pP7QGsY5GMTvBFtdTEzB+FL8RX0xMK4T6Wb
rHxcSWJVPaF2NaBeFF5OXTWa1addGEBXxD8JS6ic1phvHVAB4wMF1gYIBQDNvCYX
l/pph7hvREpHTqr96ko57hYV5DzDE6JDLmKW1doxbazv8UEQH4q6MT9KQXdMz6GI
ynoVwJzUEJCbxDKBLDkWIb3yONUQlvJMyvXhnj2O+z4oHBqj9oQyxGCPmKv47Mjt
pT9GxjcR6LiHkZbTrsMEd4WLE28k23U1t9QAd2bsybDQE7HF8GhoVZs2ltOTab4s
Q/qrc2PyDc7wTXvPWqmmYxMDikHrgmyypLvmQb+3//ce+mtBoNml35m7a0k+ld3E
Wy31ct5uvaqWFbnte1mVx8HHOpW2itiixt9vOhjDqFSxj8iYl/oc9B5gKrZnIU38
Pnf6yDfWsQnJPYu//ttIkILm67XiBg+PJ+HDsRPEbMDwqC985KY4hHAJ/JtvJDVe
gtxX0KgjYhsvk+pGUoM4JC72s+JJDC9KKMmjH/jn6q13AwJKCzuopCGugWi5rLNR
/kKfa3/PjJpboTfNIS8EmitwAh2MdOuA4uwteVlkgQHiQzfTXWyWYsTYt6DUVzTO
YbzvbEq1T50ykl9PhRqV9hmd6BrqpO6/vjUkDV2cWNbZA9dKE1StsHTcy+UgBHzO
b8VHB9M+ah79cfCPAc3JfkvcbAkt5t9Hd/RFL7yky5bRCpMtJvIoz7b5r7qUoQzd
Zddt1J91OfXHDhejSdnjU/pPNgoUXgTgn1YQCMhK2bO9eCUq84EP83MT7P3etNlq
oAT2pGqOUw9YGc18EBWGaJabRdMZ0Y6CrmI3IOghgq3K7wqq9HyIJlI5Nikt0Z9W
nioz+wmzmPgGgi9OCIzqZGF5ZQJfw4vhbqWH2m1ycDpl8kGL1Gd38ZEWwExuES8Y
YJ26Cp2jGXw5u4MmSsruZVL1R0CVP36H/hYCcnQLTtTxmMEctAiDCv7IfEEC5hT8
q4JFDDKlZb7IdqxuWJm9hlTkMSozK6+MxYgIrIlucsu6it1iZuerduUAhLLaJy42
fg01YOMDu5M1bajf6O3z8VryYOiZQXEnbynp+Z++6amdkkROm0hjvTkaAlPWavor
/AS9jCSWjQcopLK2/Ux3lEmtydBY+oVcKQ9T+1qWd9+fyHYVbqsSJzb+cdud4j0+
viwoPb6CXUSl/TfLtOeg2jel+Bg2mbw29ALB92+8XT3iTbEwhB8YkiqGIFNegd//
V9EhkPx92tgSPvnB5ZJmmEowBVqPUm1NRuU0mh7zLgoOVlPiFwJH9EUSdwWFkl9d
iC4pCd55lqgIWYa6buD7Lh62K+wnfOcsWiZd3KBa8DitsSsEFlh0NpuMslQvnaTJ
X8j248o98bBgWUWIgTL5N35LbYg0MQDqSWBmWhkoEQkcWyfvoXwER4+BBFO2RRPE
bfKpoTlr3Pd4U1VO4pS38Y2iDpdThE58rnERXisAL40hx9J2LW4twLV1EWhNysfC
4Y8kgieVEDAaNAXupvZrMRdXF9+7zslu3YnnoHYNlNUV9d/N5eGqYbWLJqEsZpi6
5rnKESZtif+CF1on2bQPSaHo1yvakrv8EWLgXDce/gLTXzuM+6NnSbT/EGA7QnTO
zRPPxO8HLb6PWQU5OocPT/3BjXOANIFf/lwvMZ6oclWlUNbGe11Iv3AMA0WtY81l
Kswswd1uGxJ4w0vuyfJgyaT9g0+dW34pbp2EtoYryFAWT3PogQ07vYZxnpWe3mtG
+AG78AnTwJOQbs8DF3DQW4lBvbTCQObI3nd/e0WTIS7S4XVERaomXDPtvfLvWSJg
ZvPPlZpS9TAxXnO5h2RmKjIXTmLz0XbCUHyaaRX3+N99GkV4wEyro0Imn4UF8ZBR
j753fP4JGltxXg7eDLHOov3KJpxNmQzIaqKKcMHPlqqXQhpqB5iv6t801s3PebE/
AeoourFb7jyl8rCS/N1ubjGiWI9bDM30DowO9Tceip57rTkXzqyyrLQZG5knM6pV
AGVyx5ccuTjGymdKjXczLHwv9G1ApUp6lnpCmD/nIxmNezGOU8nQdT+j9aJOiRD+
Y4+oRAhPdX+lbE3u9ixzaAqXu8y/vVCsJQr2NPCExR46Q87xB5kSzUJxTOAOJPHR
VzmhNJP+76i9s3cTJJNUQ9sot7GhjWrm0qyrk/iHeaJQWusID31dFcfH7Tb4CXXZ
UkVbr+WJxO6tQ+QWw/6g464z/9GohRXGCGRaQK3MTQHON9gC9fk7owiM2pUtaV9U
KB0a9r5cctuV3uQY6RgSYXpywO9ZAyovH/NtDuJexzQ45HJVsVr/7A+2YLmwWozP
oM3wu2l7COOLAGOYi4qnYAKXzdTeBLZoNou/M/gj7CFZc2687P/F2pWxSUhBTuEv
gPHDiF+8u4WSgEC0y0uUNFH63wu2gxCxiSTqJlV/+zXEfI/+NW3cdKSJQdGSpYeN
WOj4I8zjhvs5rqEz+gyxxpdT9o1/nIrCVLnXKrHbxpYnujoI0fPgvYnTx7nb0wur
7sMzsX8VbRFKC696DRBCckKiQzL0X8PCRhGpnNJmKT/L15lrZpUN22VM2+4SBzbm
7gyXVdvsS+XDQ7GMmxwqNCr0O0dBmavSqpEVExE5/lj8ebZY2MJpQ9fFdRwlVnY8
x3TwrnZ2HJRqss0h2h8IuTaEprRYPxtXV5MSBAXzskGSSCu25jQEdh+/lwj9wWh9
516vaey4Utao/hn6HCI3X2i9/prhDcIAEnDSmi8KlZnsQ6tc1MFqiXee3Xh9oXFo
MQz9o8NQCzglz5+nz5WXWOXLfWIIDt9q9z0Fq/fFdLFOIFpAgIMarF1q2pltMqXj
9EFGNqFNDDEoUOC0mxvyNppIVkL8VKZ54CSndmSWAD4U23mVWyI6UAIgJ8bcuCeo
1y2QGTyS7ksp5BvdKs0C2eG+BVofYyAigC/Vzxma/kxTveRForahoqulcuKoDSJp
p6YaSMCHQ1wrWvR6GycEEFqEOH8n1d9LzvUqG6H71t23NR9s5m6aSU1aycirh4xO
NeLuyjZ2v2H5D8/ot2gy8ct5KJ36X8KoOMVm2Ja4qTTjPDwGJ5eOL70YmxoJrJRg
/c4etC/mIYKM+QMw335dBRhzRlBlgexbdQP8HliVDPax5EYS8kz2Z78Qe0ZXAxu2
RLZyRw2ley5V0OrNyKbmttEZuZgjSPRUJm5UzEpxHZv7yD82TCwm89mx8Y4DiZ5b
JkeRdxbJGRmKLYp5afPeiuMmmf3mERvZm0kumdI6nm8FQk3mVqF7jvxLL7WIglBR
xLYtyNugvexbcnLMtMWK48CE2KiLXAYwn063BngUHfuUiMhtrwkYijWubfo62hgm
yJkjOBhL3J8TSQUzVaZXJIYKutXkNixIKeLwqo3kls4HtkjJLGYnV4qVKdRCDg0t
R+eaQCyRlhPna2ztvNhGlOA7d1uTp3Q06mvjXDZr79HfiAP0g0sCqdxLhXmwYWjZ
eClGKa4CeI82YPVRSRh6MJLVDZD/lrAPnf/4Zb060LcMKOe65GaaJYCfgTTDdPnN
SMXnNM2SsYh+Kni/eHcc3xiJa90XV9n1scpGTAe6euKz6yuOuAPfXbRwzorpRJ1T
Sh+ygBqO/+0673Apk6NutQP5gqDbQfNQW5Y8KI8ELvxmc8+SXVXC+VRzsA4JOam2
xolY/7ocE76SHZxB2lldTyW/uuZOAbVaV1UU58t2967mFLQzmqLZYpUYs2FhYxyk
eVSZW2CTKse22OOEeqUGeVSN3MsrTZ9CuLiEHvN/VOU2Z1fSG5e5Th4jIZchJKqw
IBNyo9wqSPhSR4FZH/XwYKev7hRccrytfQBgMYDJv1FF5684/RZ2Zn45+ui3QWKQ
jYYZsHlf14MzL62TuRvD163Oj+5TKgqna1eeELEkAd6DFiFer1Mwy6I97kuphivV
TH/5tdjxyAnIFjdnXNCH+9bLmu8ZzXx7sPUtX4up23EEGqfbA7eVQjfBRQrpFh1P
UvD3ABKY23ypgMLf5A5yRINnm4YfseRbd2fTwIcB+PPV0RpTsciThr1A4q8TcOzJ
EdwSj45QLefDl6RflHyWNNbbCJc+pUwhL0Autvxtk9sW88FwguSmC//HakDgYQsH
TKkvYydccQpOsq0udvRKu3qjEAiI2WEMXdpY0rw3kgXDgTOIvZcFUgxDbP5JrxnY
y/EmZvRXN+f8vGmv0t42dQeSbaJLymxnT7Kq86ChMWynQrh/JQgV3Rwm/5uhqHJo
1w+od22Q0ix1/lIc3UnLOztZJbVrYzxXkKBibq/3lZ4hGY7rd9Pn6GxKjFrfZL2I
IS4astMLnJczMN3GgcmoO7Rp2O1CzQhuyn4H6Li6fCczo3B5RT7j3+5JqEkF+vml
IXyzKgr7bVKXEvsRqBGveKTAbP8Ek9cAVeqZyAjx3N/Dr2B+8aliE+hD/x+a06FE
ntDLTDhUTHDnNoo/mNshBxS3i3j/8CzQYgNEwpwtj8BzmOS4I/mgeCCb4jLMiHZj
LG+MgfYFEHLBBgV5ml+uYkoTr20RIIDemAWcV6/FYZhKIL/wFKJ1PZbFbTIkABGG
zTyBfJbSXdgieOaK9OK1D1iuGK8eX41VE4ZVT7bSlrNW6tO35TQlvOgAgspz4fpf
+rWB3333sZ32Y34S5xR4qjPgNqORNla0tcDdqCflgu/jOQXjRUKnBko2SwEyucr4
VYDyaeobc7YHC6nLWgOzyjSoF/qzTHG/f8dYB6lu1YQqAT2VvfK2kuvGUeVcytYY
YwfHAEFGS5GNTHtqI6cwgLdWOSDWq/UuZXdUXKQiOyQ2syvfCksRiVif7Z/CtKcI
krz/VIgCU8XHFL58U6cFY5r+cePZ1eZadXaGT/OkLKn7x7NI0/7pPi7jkR+9lNG4
nAHBHjzYMVpZCHbfn989ZWXFzFQILRNzlEelooed2zzACy/4uFBxDp4BLY0tXQmO
KOiGDp7n6bMCaiw3mPLtDw0zRZ6g/ohBk5xhnbCjdFBB6eDGX7RBscRg618SA3PH
bao/ojVCmsmI/A/88EQuq1jYk1gACw9JCN8n3SWLAdNEk+JwIgZWupdq1KuVq9c1
6oDcdarOQqAAAiGxjVCxndgt1xRUT4eBIr6XCajYcFOIXYBtm6OG+nQafwSRvZ+e
+kHK9IDtzScfU0Y1wUth6stBhYcsdpkAze025MAzMlykHnji6Bvpgn9/J5Crz9Ln
UeiJd0j0lr6A8m+PrIX0VNUaLQGr5PORV+R2xUlJFQ4adqaJVmnpBupFkgAu2SYN
uQL/6EyVkMeiEMx/bfUhpJruCiU3o6yHAFeUZk8lMqxJxh+60dqsN1j0Aal/oUgB
AvG2GcohsCgarutkza3PcCloqnl06WCswhmSw7QxpT8C84D6FV7UdadlJpg3qSRT
Tjd13MkIDSvjKqEpk6Hf8baSStf5YV+Oc9ln9cuuOKSMxVRoVIP0IncuCcJAFMLL
Dcbd4v8fQKgo+fUmpsE7sf/bzAxhAcH+qNln70L57LAtMzvHEBmjI8Dy6eZtdVZM
gXDQpoiAEymJaQPVa0kevi4w1hRld0ddAusVJojtzp4d6xtCoN2DNPanJTDxLBkz
cE4jjLODMA6i1b8XhlKlCf7C8mCaMxYw7beq8ZM/ShIRZJxz1J2Jq7ceYQFlUq3O
+p5+z+RVFHwPRJRKJQ4Z70wVHSvvHGjNqSTNy8mkTO4m+qhdwkVsXQGc3S2gZrfG
6vhNCTaYnwg0I8/yYQfKd84WQ271ZuRns9JqtB14XUPMjhtET6A6J3H+jAnBLt3a
QCGA6sRWSKGl/ymlwvcmDAK/wjD9lx4m39hPq5hz3daaGLx8i+7IFea2pMTSejlt
1AKqZM/FdN6z/ozVGsWn7FqLMefwjleii/zhxgou579z2jSLvIA6Gm9wSH3U4pjh
m13yN7Th2C51KzK2Pj+ASWkB/xfKi/w0BjFMl1015IM+MPx08dIdwpiFBFUgIxxk
mO67zqBKJjxg7RB1Ww0FoMNX3Tmdc5q7BPwUYVgvbXv1gGoaF3IiEnD7pDHvfjnY
RFzh688hGuccLVsg2xV4fpH/oDSeMpvPeZZpoZ2gtITLQSYEBbkbZ5vOEqllvtJu
EYlltgClKCL9OjUdUSlDw0tWXCJCInpYCt7I85hFuXnylkI3p8T/vUNmMRJKbneI
Yn4k3Mam6lL85MzoBEzN5GDqOPwBwWlOM8WmY67U/6IftHkeXAdG3YXlDXTeqrJ3
IhkzRBbCfqnIs7VoHfJY8Su9pXoDAGzLM76chOsLRINJN2+146WQLjVEOE/vMCqq
Wc8vb7Tb3eTzcKqYCt3rWyCYYlRSn2oV9+GJVzpv820bxaBMXrj3Qtykof+HwTtO
THkwXgA5HkgQHiGf2XycfVnsW6BZ8NcO/sSO1ORagYPAwK+1i7838KPmipErCko3
yFli4cMwpMO4a1bo3f3sNcpYqfc62Md7MsrrHRKpnZonGr7umOCfLz18pbysYjK/
boo4OErPr00J94Q2FdXssIRRVfONV1JSqwhhnySwtdtHBjEVlmXPepbn/rTBVVxY
5MbbKhT0sUdcOEw089dMODCEiGGAQWAVqgqQkvMDhhV9bJM0IunuDrG1VpkAiITT
8VgnSFrP4JbD6k6R6Pll2BhGnnkFnZoVm/WPf4gFQV+fJ0BofiFWaxMYFPyQw4LW
vs0ZMzNROc88g5W3PDB7lhZ7qPH3/vLn1riGY5/14jKl1YD//nafHo316ZLF9KrX
8WhqwgERBdBJTdHTtkeJEr1JNMWSSGow53wU03euo0r9Q70465HuMATWF/7mJWyg
rnH6Lrop3KG83ykF/qzVBu1No2BU/mgm7sKd8m3Hzb+E/SD9NX9UbPTMDl5nFi/D
hjTgR5TA1pA51lJ096oD2uVdCpco1/TRFdJAf1W84zLHLRdsaZn/3jZPWuPAkKMF
w9g1HPkGEyTBf4tjiBcUIPluObzQ/yhf5Iar3wnaWq/nUt93HWVeCz2NCwUXa6Dv
xlfvFDTeBCpVc1dJZ6bfjLbeXs2FrxrwFX+YexZu+JRd+7lzqlubAUyBULEcra4I
fJgJ6VjCM8pSdF7NhGcGAga6vzAOhoeL0q6vpu6NJEP+Czlwpy2uFESCQg6ASM+G
VLpXWHLa7ti1nfEulJ70LYgkEaZ6DKjXDieI/FvQlns+t/VYxGQsNwRizZwQyYEO
lT+kspt62GnPd7VaQyqJ+Aql+PpP8rzXn9LQCQih1TfmCEZmNDZ3Xk0EjJMVl3yW
CdyoiDZDEkbhv3YkR4sjoylxq/9rMX9qH+8qYyQZxQGn+wR+KN6v0ZzxkUmTsave
21FDQPeArkY3GgMZiH3aVcNAmC+jOf8WGou6lipXTlCFjzMHBIJf1vlrVkKoFAMU
zcYPXqoD/0JGKlp64sF7QihZ7scksAgvHr2N2LzLNpUIpBkD7tx4UH08P+WloKo8
HkUkuoB9Sm/SsliTtERSG+yLUrcA8GE4tpq/qZBdfPjbTHwTElFNZyS32jMEHEcZ
F4YX1gi3cKveiRqvO0F1Ug6225m9A/b93WmKivkLrgYDdaDuYX7kZVNLmxsPRP47
xyx/y2eexnD+KiRv7auPmriE7BqNXWOJnuQlW3inMsklJODl3T3NS63vbliu7axq
dZOQdBVSMotV3QPTq0HnohOAeVIPt44/KLBG7UEznrb1gsIMewRWIDzZqzAViMng
nbzZWLbrbUO+6+gv8mtc9bgb+zXAKpFs3fnh1shEW0/TALCJbh+CDz6jnwF30PVb
uzZIB6eiIEVal5gdyakmkZvf5bixGLx+xOWumeJWau2yWqIGcIw+StaN2B4RXw5Q
y9LLL9S17MNLRWX7T/Y1bubtJEBrE1EWRZe8ydi2mS8JZxuCoaXinj5bJfn+Pa3l
P/0H+ZEtf7ZDdfDNRjHOCVqBFqKRCpeb4mbgej22mvKETBNDQLirHJwdf+R6CD2b
o35X79uhw7G5zBKy+lI1O4j0zQBR6W5WF7ctZtXqlEGOomVavkd51LtgWwArqgIW
V9X0mV0ZxWL51muNDKvI2PvULNQR6Gil74hjrfTCYXfISHfNaDmHe0OJFS6OL3jR
mV0EWgjYa48wm5OLOmbExtH3MBe1DbTJB/4uBQAzDT9gRrszoiFFn782hUF+BtbQ
JBIXp1ypTTN3H8x90Icyz3mIJli0Z3cpoc8mOPNz8z92CqhGMwbztbrgS3kBmvoH
m7FHFn2wH3vr0cYrsoERb5Vi6j03dNdOkwuhRiGSAzbQnskchN+VN7U0QEcbZklD
3aWPic1TA7lp5Mae99lGiAN/CsRpnkza600Oo6p4ZRs3s4n57x/dIfBiiW+Dtt5C
IkZ+dHADePxp8aQ8UnJnbXy8QNH6IBCZksUJhBX5LydDhg0u91XESw4UI8vTW3rP
+juIVXY9VuyMptQFWCOzFEZr26oaCsor7OTwkAEQXQf/2Jamhvu4B4K3B3b6XGwG
iuhclhy+OMPfPihIYkI5JiwKFTdut1BUU1sqRb38x/PM2jAYmZbtsPcCk3+CoWkk
+dlJYSwl5pOQeLFwUocuZEURgoXd45gAUhxwHlAP6kujwwiYWvfXvm6Hp+/+zJKQ
wPt6z9/OEs1cHVdQVf/6Jg9k0S+4j2CU2wAh7NUiQQ1aw+rAGX3YuKZep8MGu4Eo
0ZDHOojxjX6To681xf4hXQ8xofEerjIKsWJfGD4OZME9eVdcJk24wv2LwDlp3Sf2
mRyEzwz+OQoiBinhjTuoL+XMeW0xAk56L6XBsMn3EUWqtGF/blMuGkTR1E9LA/zb
YrS3KnZXMVxIuI6NfktATlKBZdYQVQzqVAtMwW0FbDrkFC/iEwlvJuwUzBy8quGl
/PQPl4rhKe8y/Eznob9mJ4rpa/4rbRT/2YWz/cdcIiEgHCrVei0FIRGCqlRpc9yR
kvLW3J9RT1CXx6NLjtosicHI55OJD3xas2o1wrr4Asy+AkN2Bn1Xhnt2xuE5Xq12
PXP8QlGjIoO+pA/50z1aYa+QCbRuHl5jsSnvhUuFBTxsJly/oMqMwI2xq02ViOsi
xkCh3ldELTGXEqPIgVfXYPymBAo+l5i4K/s92YoLgiy0JYMCDJR8DPqrD7LLsAV9
GydhN8DAiEd8YfmqTlR1FbfW5KEi4CZLCdvf6gH7kMO9oXraMo67TCoalnmETwX7
gN8sdCeeEIvhM/llOvZv/kRmBREleX8Acd0aeAJgmaS7Xf3dRIfL+a4Zy6k3GKl5
rCImhht6c52XkWeZsjyPocslLdLlz3J+qeE1WmZYhCXpr2/MlQ0OyX7rSm673qtX
SVtCkwSexbV0uSiUS/FdnIlQWzPPwyPC0HA6zT0P26GAOM2krxnecHOefn2ybZnj
nh5WSX8xlAMVpll80NpVZK4yQ/RRY1JN5V5IOSKO3/L3ZVZdIWj1YSFW7hC3HNnn
s6WOi12+5TWpnG9khlh/Vcd/QeNbAESftKTtT+60SXMjKFrtO06vDqpFsxh2E5TP
T1/b6Dzx1cSzUL2/NgtkEyoZhEYm4Ii6zdGq5lQekYZ8pum6MrfXbv6CCHKFDuoH
H7TjHI7mqrf8hOrQJSPxFX5FXF6F202c9DxdbAaTR/5gBMxeNqVz7B0SCfPo/dRw
b2Aa6unlKBBYiXjdGRJ5zux30GcZXKyfwRnCOjYjOjDjxz1abf6E0hWJRo7s1YMF
xbnuaDLmU8LhnY2JL9f4itZJK8G4TaGAYhakFFXMFDrh0LPqIIoU0ksdTtxdQV0Y
mT+bUbDnlHWE8t7kRo8KWrHdPrLtsOHGAaIa5Avx7UawYICnxskmdG0jr7gAMuJN
fnm5mLnaA39QIyGS8lRkgGddOcgW8hYAqrwkLvsOLteSaB1u+ovgUodReSfEn3h+
CaM3YoxJ2ZiSKdr0qK6Wn7eWfsG6+OcvuE8Dp4THpnwW33rtm9+eadeztTZvaqIA
i0TCTJpQsV5TzcZdYArC9GAeQW/9+gy0Fbib2D1t9IKOjBwz2/0JgO585HSSrQmy
PXbLghBNMLnkoTR71jTAEC78zAwFMeZ45ZK8QV6xfgofGEpodizjgCUw7bZV5ESh
tC78brHlOtkiXqc7zg6kd9kFI8vl6VAK62dpy/fhYMA0O6Pc5trGgYhT+97fteql
fTdxc6EyY0DUKpr/uPUNAQb6ajKdqxKn5XH0MpFKRXEJe4N4PMg1MGlEpflhGDub
10xWtRNihmPGAl/kw4DKW/tP3rECbVD8bv87T8W6GD+LAmrZ/5YQM3huOAtnNlFK
ZxT1wnMn/W7sfulFp7FLXhBRb2yAHTm3iRV75r2AJrXOUCQlx/Me7YuZpZ799zzf
O5PbI++do/V/t9WXdQJCxjob0IbzuoE53HFb9mGCIYIs2JYLVutLvvjKHfcRj/GO
VTVNiHOJR7p2TyHRD+esX4Uo8hd7KW4ppgeaC7K3pOmJt90PBLZlSsVtKOnkFZAU
ohpWpZSJgVmWeI3eWedPf6A5F62XlIuh/0/gHZMDI7q2QKdswjWTNODZ+6ZpE+nz
RlwJxpB1pxUx65CG+Ye2uAH9PlNB0ANYfXCFVQjpgTQBhjnMKGLx1BD/FWfdgQwA
N5DjHZ05bPF1gJ/WXpehx60OYuzwkNkZSKYXec4M+4ZZZu2ug52/R392zQJQkUQz
ip4ei4CvnyRUrQyXOhjNytUE7UyMWSEtcGXV4yS79nITYszwnrQorKKBpASS10YA
ngYLPBEDzre33rDE1D6Q7RysP831svMPiAN0BWHCVvYW0wx4gZDapRnnyaxRT7Z6
1imYAG1/pdxg/u08BGFWoFWsb9gLD1ItDO3oaVsRIpYqUn1EiSzCzWHrpMGHzbNN
OilfMgw4xbATemSpmTxivgoaE6umj6x9L6xJQ54t87/NJ9Lw1rehiVO5/BJ/aeDo
v4Ov2TKbgwTZdbaOHrJDfB6xZBa/qN3OhBwIKlrZ5fBekZe/tkGaiTjDl0GhVo69
i9X+NuCAtMvM8qMslWDd9QyLGDwEUHoGsEhoQANHh63qbiF0tTVsKRdWovgmGusc
8fVSs556dAjelSSSshlwNhquSfKTKbqTkRY8kPCG5GFuEE37GaguIdEFxc+JnYMB
IAt+TI23r33/TtbCLY9g5kifJxu6Fb8QgZIhE5UmbdFpUrCiP1Phjz3J0+iB322q
iSQoizYHjL2N6BDcTHk03mfGEoAssdO1+vkPOmvo77GiJhb/p1HlZPrq1erVB/t9
ySF3IOXinr3JMjKEW8KBjiXY8dgiyejStcFRO30KHFWRKxL/T4XJUWa/7JRWNDb3
gRiU2VVaTIt8Lje0fmvCvpPisOuiADhv3rADcjJ2DvicTb6a7Ds366lW/B8dtfB0
600ibHHBkaSI/h6+5nvM7oE+B8512rKKRanr94GsSQL0TOU32DwDtMsu+Y4+Gegl
7TI0BdyrIE9Nl6cDIrF251RQjk4osQqEMGHOWfTJSf1u9whS0GjNwIVDmDrxHzNL
JgzUJWSNaCn6w1aWqe11VTmioMA9lJghBDsOivzXf7SI5SUlfIG+qfASjGhAFTUW
jq0mkOuBDTzpqyAVy4EyCWRuratsJkOTTVdgZOEDr6RHCvvTSYbeCaAlzaleNckA
WfiVu6VjXCqEMBpEJXlgiAAvC/MkzhQvG5O8X7LzLst1dHkERk+7EQqh8ZKTzhVU
2UcRxHvRJWjm+sKsYO8Z7xHl5rs2xBlCPq0s0Lz1lAmG2/44t2ZQpYBJxL0TvoJQ
kkVjsyuWKPwJsLPG63Pde8vKIQSx7MP5JMyPceetS8xr/20U8NxFrCoi410hPH7s
ENy2YIEEUrDCvtWEEyFl2K98tM3+TopGIGnpGqe8uciQAaAsvyNF28oYVJX/4ATG
CdKwHBWZvBOZvwx0gojiu8mzRFCS/m+SssWrU1/Wx5C4kiz7IPkBNdatceS38YzA
A4sqs2KT9Rk/R/J5phjXfhUduGV9F9B6rEeaJ67Qz1rFz3t9/AgeWsTFR21y0NlZ
7oRfx8KpvgZAvcG7KozymnDoExeBPpsrf6rT8ugpYI+cxL/ckH873O/cRdUiwALn
7edZZz5tLf6r8lQUof9pCJDDFHZ7edujXwzKGJ4jsS0u2okG5AYKESzvkuaVn/QL
B7EqnwmetVoZmLds1LSs3adbCgdVwtbszK/k7eSk5GdNUqOG0AiurdjzCZiAFK8v
oZFcrlxjNTxi3LiwrJm1AjaERrq39TNYlrrpw58FEgJsIlonKqG2/NO/Gc8rICiZ
Hp0rDhBS/XYp8YQAowxZnHulddYcLrSbzd6gjrkInrlcoYvlRgf0HiaCi4VpRzsH
yi8Yzzi/iBCw4PkptX66KAulysRF5fibK5eLmQvsPuoy+dvwe7sK1AD/8as78FFk
3nJtXmUyS2dIvhnOqTqjL4afqdTnPDC5jU/W6GCwe1sWjcZ9CZNB220SU8+AmBjx
qv5GEi9KWtzrA72/rcKRAFm9Qnj49eRonYqkrT10pw3Z36yzxJpoLiLW7sHB/qlU
JxXG2W+CwsRAGFjIQtwyiiYP2w6IhFGZS/mOipFpmNKuSqxmiojXBrzCy7wcikLU
KY2od5pDhGw25vlEOwlQAtcX7gRnhgQdtnvj8GCXFFr31M7jMFMpoR4l4NO9cHZW
N+x3j98Tsj8d6BBcAufwSKnxj6l2nUJiFKLtbmvfAvqdVtilIoZfQ3ku7lWwzfi2
6Sd3QHW+cxZmcOZYrDKZdVxBvtK7OEuWDTocXL8THdsgbGxi4N86VIfxyZqJh605
vdHxISELe+ucEDnParhOh5kHaWk+4CZdp+1Hhcoh1V8RgOsJmPA9T5R9uQESsslW
3M0AEh50bLTE1fu+9E2TgoIkuLXFqn4rZth3vvyWFq6au1Ufjh5X0ev6b+S7vrr0
kztHbP7rwtCndXkWUgysYbwA+tW3k9g2WWSrBZgazrnj0LrV+8ZM56f0andPGQd4
RrPRrpIdRX+HpLuTueAJdjJVcF14bNod4p0rKFIZ1xErS8QP32vULNq9QwNs1ZSB
pgXgjJ5ysIcpgFLtz8NwSwkoUjmZhAddebggAcTcoPeR/eIgvNIMtdI+YC4rHkxo
2NPuXdzQ2m0msY+QByGly3+5Y7CTS/Ixx8XBM63RLL3EsdBzuzQUddsSLgNJplCM
pLkcQyVYi6xD91h3aWUjHcXrMvoT473FF0+eLTYEj+MS9G92iILojUN/OkkIeOFM
dJobfNyHMM97FzMAGB1SiXcDjnC1wIzwcmcCrN08LdmpKoBBuLpu47uBNgK+Pw6S
8AisjpzYP5mgunkvCW2VNDLst6dQK70xJxilwNccQOdX9JdUqLOAAnUR91hZ9Suc
+OHjt/1eZar0NRqjQLtKS03JD+gOaSpv8QZcb0DfY0IE2L7cb303enwEGHGmnauU
Xk7yqaUKQij9ZO06beNkMQDu0Tm19cQa+1bKr/8ZSrljF3UwENL70yQAYIHk/sOt
/gXLJU+ou4k4LGml0IBA3g7YRYiHYwRS1md1SxHyaajRu31Dj6tuWYRD9QmXvDoL
wIW78B+4imCmtl+eIxUNAF13hy9LW/X87ZAbdIOC5yu3MXUH3kP/skg0KLyS5uqM
TCJFtcY92lMDbita3Hj+E9YmXnbXP7enDz1CsHCJBASTio7e86t0SisxwK4idti1
Y1xp+JmoYhCVmWNHbkniisrXlEeY5XeXmvREL+sIH+jodESQA7ql/oRJR4ksiK20
PWINLX4duPikIsAhMiT4zGBiyER+B05NHmkKIl4TBZLF5+G0flyyMGxA4De3DNKI
Q7vo6vktrFHhB5DTDceanNPHiNsA4OFHWraUpUrEOAtx8O8PQFWBGbzR4ekNToK5
LjlX2NSt4GEqFRlMF3Wo/Py79ApEx5roeOuIH/yv2/EsvhpGQd2AwAvL20TdmnpU
NAj2Vl5QWnzbGu7w7ZyYjle9xrCSqlXOHhgry+500zcylwD8if0ZEO4qQ2PATxxD
N4Ku8d3IkbARAtYEDeGe4CBDiFf7HGoqeKhmysNZCzBGinUwGhz2oPP/lQyH9INI
n5uCuwLVAPBz9i0e+hBj3U08RLR7aeE292aDFY5MpU7fi5Oelfud4eU/L0I7LzeF
vFrhLefjysQWfbqj8XUSq0GVz9U3UeUpkRt8ew/yTXwrj7fiYqGf5QNj6Mkqf6ly
GsA4BHaRpcRhP+X5QJMs8FOwVvODidnhl1fKvKjxRB2006c8qHn7F1gK1VsBQ/jA
Q0CD4hQMu+e8bn4EzFfdjTK2P/aSj4Mpe3UXgztqsvuh6DYyAmZAU76gaocnXs2Q
WcrboXFnKffODcVnzt+/4aZPjkpIuBAbvb4zgxakmBroJUcg16XEUVdfdAtL61hU
aVH9tY7w3L8CooZoUL4A3JBS8h2fVEqzh/p20yKEDeALoyI6+GsJ+O6H7k+KYS9n
hDLQ/4iNsbPByax+VqMDEyfovBDXBBqMIx6JoFZl0rQKEvEhOOpKepVMeKT+2B0N
EtzhWEABOIxhu7wFajRoGZ2pmaIP8FtBWHs0UHB+WwtGokEAFnPFR/uhVV2MoELM
KVWq7Vn8QOeHBByhnMZSPSguQ68sJ5vzwgy4/uFbCilJ4WUIu7cYb/h5oGfIUARU
0+4hdgb3180BaOHfRe7nXGiM3fQuHyPSNzZr6F1Rxyyo3ABGnXwfQMfM4u4fPZXx
0UohTv8OJ52oX+vvZfGse9TLNT6WV3pg74DI10qzq6EgRn6eh6WInS4VAm0xgTtF
DfaTKQf6g2Zp4DbrHphZZaZVB97pxd2k/f+gmpjvtZCLuvoeKn+kRZj+tZbQ0yul
AQlItSnm+23Akzc90bR8j55WTMpSlL+NCVu7el73wRPmb5eQTw7fvOSyNs9GiQL9
RnHGo2tXKn9DZefl2nuoMrym3u3hUMApN8zdqpqyKT+2iFj8/E1+amSBPXyKA00I
7tlMmJdqcfqatJEC//TanURQa9PWaXHNrvI/4ZpJfIv7ReCy/CEeI2xowc8tvXeu
PpyggjZar2suKzFkRhB8pYrBdhOqn5d0avCb7lm8rxPjDHKEx3Ic6tjRWpswkkdf
LIMP3Qe+8Qr3+XJ5rzAh2wBirqk/3bZ+AZagd+QKikfd0yAwmk4yT2mM/e9ZdwpK
q57XJDCu/auqsGs7ZqT7R5TcBP/RAgGyCaxvsjAPeO7MOv4oKbagqWq4vkDX97dM
S+6SWs/aOeVwy53WVQ2/BU15Rzpunjg4hk1/GVfpepa7T5IBdhthrFqVpQScK1Tt
ycqLqoaBP2ZjalIMDaHClcZyUr662c0Ysi4VEwqW76mHi+AhsW28RF+kYhkc/IXt
hJ2HiYma1rozQRNXeItH52oEY6Jb9GbmOd+ZLi2DC8n8ShpZkYiGErxKd0M0mziK
Ll87Y/KEBMrf571Toq3Bude2R4N8Ee0OF/c6kM+MWlyn9RVFGT3EuXDtcHFOnPHS
4J+pdIt1IIo/FGvfzlTe1u1ehcoPKRitWZ35yGgIyUiZOTWChmDM8o3kqbi2tVAm
VHR6shQfv6B4zeYhFXRV2tu8zfbdCZG6xooN/piXizLPpayD0I50+bawSpzFeq/W
YMpOdEwJHmFBhKHAtQ3OTbAqGi13mMif6FLuuEgJah9P83Ry0J0caDqAFq49cGAw
ooxkaNs4N66mDC+MGK5EW3mNNCAgnz/7WHrnPxpPhAQao0WrHBrtnU1tcrS58/j/
z4IkKHBrs9rCcoMeiEmXXXEFfjj6UMn7QJRLcxpK7nNna0Idzhw18j4gFaIN28iL
sMmg3yAWcXFHfpB7WgQOlXILpKX6ehd9HTD3l9kaKPqGUkn3CusCGA3ai5PIhE39
grBDQYmcFG6fwC1CmYo38zLtUOY2p2wsw/edrP8ewkMm7V2TLZAGvbnFdqAN24fX
tqY0JP8Rdmnj9Lq556FwmCkcr1pNUFwU+DUwqV1qRaf4EJy/1NlgWkQx9YCkjOnq
KBhLfb/aowjlqPFFzdEZ7hlWN4Fv+kVIhRwluq00P3zUTPQoP1e5W7KLb3Da8SHI
ir0t9fKiMJU+xouTaBAoE/12Eaoav0p+tveUl6qv+9KG65a2pq78EZT8iKetlqwE
PKcEQr7PGrunJn15VJjHy9P2Ns+2b8z2TMadbLNYUBL8qZfS/Oji788UYYS1MYh7
QPhCxvBDbV/zivfpSfHh3dy26DrW98Y4nCGKvYb4v1wKR6ku9eZFd+zOJY08wd3T
dYK/bOQ8sd/J7bPMjH1IpZDrmWeYT0JAaq2jlmL/ud3okvZEulRCgGVcvH0yCSrE
S3Dtl1V/vXJbc8bKspBZovJk2PoZdybwwG51uGvp+cDFhSwN/7mPyR9knAXh8a4V
0arhokgGtkM2FNBEfSBojiOMc8Jmqlqahhbousas4lVeY1JKA09CwOVvQjgAiPal
tt3S5xW1BkA76+BlR9WUPRq5GGLptHJcRTbr0g5L4qZvOtje/3JHSjb+FYQQivHT
uOnhDNXt+fVWiEa+cu9jER28FGANLkYVbAt5FrGJIHWr+At5S8SQNqn+8E8yG+Dr
ZXwjv/lyZeGbtjOWjflhkZ8Yebrsa7GCE4qyVvO+KF2MmhFIlRymwUBJSSz0Cv1k
UHsCkPl7raeRtRjbaUMjzHL4dC0qa27FomN4nM6jUTm/M2BT0G9OhKCKhdcOiqEk
OHX0drtQffDHNUqrVBnOaWaaz33WyJrrZy+w1IuN/VDsv5kvnoTCEP4lJNNPbjun
h7OxopK69m3R053mTCy6RSR2VtP5dDxI5UYNwIU8mKsFgq/PJuEPczg5Ss+9W2k0
DBaTMZVyRqW68hf0c6xTQjTUWb95OhQ3AVP4Yd5+dXJ2OzmAXCV+FHVRa9VeDd4l
Tc92Za2/jDvRzQj9btRfrc7RgohlatO5DdPCyvYWlpATGQakPFL5ROTlGVjRP615
NDPvKqy5+vXE3SKhda9RrEeVrhDOrE7pLzpeljb43s8lzZ/SAikGSv83Ux8iumJN
e0RmlSZpAzisamcweUnErZPeC1sg8lRaoyw7zPI9fertJhovOHArmJU0ve4qMim2
SBbLCFmveWUh0nlmTMS+uneXhUUlAJiyikSHwJ/aTzlozAxFlWXOUO1ZwMvuAPTX
nsDEMHd+fiBgHVzwGipScAqcWwVESuKYWdceelJULfsgsK5NDeY0kPzbbidW1uyW
g7NCqqo6Q51HPr4U1I7/GcwWWWifkrAQZ2cgcEy1diz3S3TqWkh4+tundPTXE4BR
0GjS+SXMeRqbZIyl/5PZOVEsFuZ4JDGSs00lbDtDSlgGCWKj8dIC5acoMoXk+SFv
BOywUeWgM0zdUrnKe1PnxV9/rGCi04oiQjXIXgVy8ImwWRA3nPI/d6dFvL4Zl4nd
Pgr3JU2/ckAUdVcH23hjNFwiSmdjns8o4uNYse6LgsUC4zO39Y7vsRNieTRBA3lR
dgCAooxfTtR0MV/dw+7pHFzEcClTCwMmf3j/nMx06rO3BzEN9x6PaBTFDomA7s6u
lamKM4BiDa8V14XyCNdUuznk1qCp5KLspPgBps6azD/zQ54J18FzFerjU3tQ955t
0s9gLAoqznmpxpDnBYKN//tHMJjsxQCMAetBdJwrdJnrPdM5PMDnimyv4P8xDhQc
SQ3uu9c4Ub8iiRjIDCN6AJlhcefH6624sXlkmXKzKyqEhDK4rli0JWV70+3EI9pP
ceYAr62OQi9S6Za0Zx9eZpw4g+B1ba8dxxgfGx/4R9q2DDMoeNSr+abir8MNpXv2
TvIwFrH7brtmvUxUC+QyMv7tX+MQ9cj4PxLiBwS+S3RSk0Mw+8a/ovyV7uQV3AWk
ZuZl4N4AdvlThoKHjLVJpRYzAuCAsPoEXTu/1lfNEqFjijJlA6O6/8FKy/LjahV0
zp4QBA34nZmCp0oLTv29GqR4YEfv4H7BXBI2lYguL4Hah6UX3f3Oi0Wid56LPR1Z
wFJJ48zC4Vk1kDoZOQPz29TIVlqDd1jIUO7eCHmIvJ1KVouVKdNNFJkZ970G+0D5
hC0+Yfy9jWu1p+F6GpA0iR73seenCIo1UxdjxrNYGgMMCT5Cmmtjj0ITRgwye0bU
T6X3NHR5A63YwM/IFbOVYbWB4Qfx6BT+gaS610n9WN/oVaf/NmAj65Tk+FDamJoA
cB6bkb11mZhhEezamUHl+gegoEGXbRT07rFmzZjI2SaE6FzJJPeJEkIzq5FpiNg8
cdBVFNRcx3zDKbAeZu0XDByS+mIQp0g19uSIdeWYYA/9sFeAJlBRgIHJ3OmLMG8A
S8zbc60fJDmaDaHEwfD/AbNpVXm3lF47TZOxJddg+npboxUSLCWqXcQt/CuluRu1
vfqdlWST1LMSjP0sDoIUjqPSaOJi69MNNwT+aUkJ1kyUlO1Lt3IPYBv5bcqeBpgt
nALRy+39xtAa2kzv2BXcfuhgzAS6hfrza84+RaojKKa2r47DKidF2lx55/t/JntA
q4SBpaaj4R/KXhxIYIzEw2aWD6eszGHDBD8m1PR+a06LC3mJrNce2MyTmwfD3M6b
ZnbJXHX67E05Z2BzN3wvnGJeU6g9sy4PpH5J4gs7ryV+d0/xUdfJK2sMJa7D7JgJ
E8G8vk0V32z9ruBVEy6l68iVUUdLY9IgJOTwQLUoUMl6Cdn/S/q0/VNIpivI0OLL
m72482o8p/wh9+wKmuVptNhXcsbD0YqX0OYNrw++YWOlnbDqxzj9/ZKfgCUAm4fK
78RQg3d2QwFDr2kYoVFDNu/B04rIZH7VoIzrvSCM1JFc4SnyUogb6VePOjUYvj1c
m4w3ZjRC9heEZedAim68VF6S4MP0bV3Y8VkYAYTvC+tig4j/sh1KSUqDAXWuFnf1
B/i85X+tW9M6PopG+igHFVUCZwkQ1P0NT2KbUp9EyENbSgHg19orWT8RWu7M+aO7
evjUajAKptN8NOloMU5eUtKrdfkG/uZADzAia7TXZ165V39E7kXKHB6qdAr5/VUT
dFUvXRIcQUPoW5z2C0wVJOV9GZFXNL39StjQol0KgVKl+Q8VRyXKizmwC1sW9nYz
eT3D+BZhX7VxqFjB+AzOqcWpIaioC0dSqG96oFYqja6UGUvf9e5VO7WSRDFO//Xg
211pQcQFOUfY9nOeTV3RsBEFl9PfbfclS1fFms1MwEKbPBU5qnmtzbR3Xd+vC1zX
7kECs4APObieVXnMIm1x52F05tZLgGpS5Y7SsMFtpSirG0/Nh9oOY49LH4j3koVZ
CJCw4tUTjUO+LBpzWTYlq843nVnnJZvw9ZdyPlxj4Vjo9vVCmM5iQvtj/0Lc6BZO
AM0vkvzQ1r1TqX5C+g+cF5RYnEra5jioNB+a/ONYC3fZuElDmKXHO5kxHKYTmjRT
PYS5cDMbyVTY6D5hclLKLKo/N444rkpFhAnyOw92mn1gI4ihOOXO9NOjhsri0n2h
8mfVLu5NvsXA1A9646GzT0crUCGQl8Tyw8wmeopwz1qnBaQ+tqB82o4ZpGCUxwmB
aiKSc5OGVkGKAqhDH4XAb86Rddtk57/M4jBFS1UYglwzlXiNsgFIXOBvXJwIvSjb
5eaER83eRO7gcNRzWvfT+VzGo/wl61sF3UQa9G0zyzHql9QyKteFxAJ9HtuZ6fdA
OxVaeXP2exojEXKPvImPGDxWyzOP2M8bL9xe/YPHRj1frWFqvJUPUDG15cjIwE5e
ZpM8jLk7NZM6GmlWD7wVzbrY7T/T/DTTPWcJ3UF52SHXpWLwNCuBq9bbPIQlcwDu
X9y1QixZ/0qdUeNpOzesA73Gc3P3rurQJGse/au4gp6cUbotEgbmHsUmcybcBCvi
KKMN4SjSZUH4PnvCdC6bTZJXqSVNUs6AMz2HEzLFXWiqKsSDOyGkhLa+jfa52Y0d
eiPSzG/38YSqOoUs2Ofo+DM0rQMEbIwf0pPcr1kNY+UA4g3eI6rmeO7iaQBGqEoE
IEC//pA5CR2JbGnB24ZowjllPyvw3RKspdhMArCP6J/Qd/hj3AsnyCNii7NUmjRM
1s6nOsAMYwF/O7BBCLLKAk3nXQAmWLPMH/9hHA7dmHIUfIFF4/v9Smjxvk3gjZYI
Bw6tyQ5yTk4OFcfjHJVWLcoUxIgOiHevA2SYWgpg4TOwck3d0Vc9y8PMFU5Zz/RQ
3voWpfcLOY+J8AIgpo8leJfNrt/brhuuCY99HTzCc7EblyTnB+RnqGd/Dm3jyK2m
0FwGlfrDS8DpZeFITLWxjMClCkdHxrCvcgafV+XBqmXmHduGsLaIAEJ3fFXmsdRD
AkUn4lokcE4t9ULT6mygBBLH6+O5FCpENij03OezoFlYLQGTKIAIuEcanZntZtTD
yxiISCaViL0sesWpDKm8HiP65FhgOlbuRxRRKxVYjlDoOGh2Ashpn/D5xJetMu0n
AOnBU4iYI/Wh/uZ05tnY9iAs0xhuN0Pl8CWegZS79mvHbLsEZswj9MR5sTyoET8l
Hocark/OZV9C6XbXVKJOL2++6nNNSJZX7xsihtgSz4j5FJpgCd2UtdH5dneSit1w
jSlawDYInsPGKKYdORyNZvoGfnvA2CxszGiCCyrB+++4r4dgawE5ceLBBfxsieKa
t+oEqJEJkX0gqyor89NN9ZDbljsy4dgRuSRHlMGqmf6QtL0Ja4lVSs4bdb9uVPYF
79c68f1wTjjAuSJpVLJhbjJ37mGFDEjvzSDVWKKIAyk+AfDgy0yy79QVt24Oj896
dbIbhkMJCeE+bq1SVd2Ad3kK/Q5VKByTvgpdw5B+eyGM8pwfwfdzywWmYD7DvxIg
EtpzEJ72/wk3wLSw4UzIHqdRvclfCd53/mwMlbta3EBImSmRwt6/lT0VxhDE4ASo
fE/cStyzR13qufh6ZctmMfD/Fv6s4EA0oZY7Dd0EerDT06iQ1e3Ovd8Ef2z+7hId
ExXg8AYzugc/HRqLtJg+e6cnxUq8RTM4MswFrjDW4RvdGlRsN6kzbff5DJl+v4V+
eBSIS6YmQss/phULXuOg2LfvDbMG3xzqcjH/LjnE8+8rGXQRNqhFqA0t2amSPpAY
exXdxPbOeK9T2HS3dlnKMAhF9kOpTkt5ullhQ6YMG7NwxN6XFgGueJiKeHvx8+00
GbBFe9I6RhkC+4Jkc1UyqmVW85OghEwlg0MyeITy9g99Gz4Fo2rzt2dNDsEj1EJG
Si8dwXJmT38ZU/5Xa1QiOVaXRGY8pf6dEuSGapfhyQRm9GWia+XUiEav+Vrmryos
KLsIRrbojcW1k/tqT0n+9VMsfSL3FpoJ6dvBpREyKHsiIbEQqChZxP5YoUbygobO
yId4e60+Agp5gHYpAvyst3Ou+hY1ubbMHYvkkAFy5qDgNm2eKXvl8nhYH8at8CKH
u/3kH4oLRDyGzz6+yI4d48ui5gEI4jPe3A1LwMdAwqZsedPr0BcZgWdDe7OkGYXB
LLZjvZeQ3jujAiXSoBwLpMKq7GKbcS3m3WGrK/phS9n2FBEAt10OniSlkqrFQBbB
E85a6jREseLQtktWcZFv1NIz+kkY/KVRc8iWVTEcQn29Ixx9a+91n51lNgO8t7Fm
EFYiFiUQ0Qd+bNSLxN+LUZ8Be744tQXGQrP/131JlGolRxH9rjIb+bejmaKoWbyj
wGgKj1t6HGbvvKNrHOldNPSKaX5G3/hTtWSqHEEnEd1FcZ5EQ0XKJj0IAnN560H2
5aZjmsH0D5oBAhCPpvJI8WZadf1L4/kJYI0dHtEmIZG3bvj/z7uzslyIR5IcoEG4
mRKVmpD4aMrODYsnfa5KTt1CIUaTJgmIWt7arUguSlfXNSkJpf3JXXHD/3V5BmEL
X66YdHnOQkgpcFP7wrJVdLKkhLyx9QSgKcCWkG2HGs9Qos9UWD4MgIzQeNk/lLxS
hRlmQo0F5YqrkjBD34fADxaHwoGMy/BL8SSTQqXGqlg6fbOzJ9Ll2eoqIp5o4TVa
kwOMitSWR8O4s5Z1OuwEJT+jOkO0QX5A2c7wbOI4IQUmNJGNHy/nPjFOeR9i1gCk
DtSrMn+0YdAJxa9vMzTexUzIH4RKp+B5+t1dZ1AwZj+Lk27GAbDdUbsd7V60Qoyz
UmBbXiooMLpc6gUFn46MtrxNUjkvoWZUhqsJvvT55BxbcI6vjng+KQktysomdKGQ
6Ow53XPOaverGo3LeHdFkNg3iEbo73fdRtru+AQ+tcZ5o3Etc9HjCxMRfFLv0oWz
4iKYRcRpnJzWl1E/DJh0UjHbgFvFv9SSxqmw2JMSoy0ml9dtuqS2nKKp5i+ftS/j
+iPhJciYYCqo/nW6WZ+Ws5mG4ESZSnSZbxL/crK19jVDOPsks/DpKeVZX75nFnrX
6KhmiGsyzz1rZefvJseSlIbNizCuA4RVD91EFfSsJZHGtO4oTOog2VVt8Eti3YnG
TXpmcKIaOLyFV2tlr+wdmBiKoKvDd1FejJd9IVoFZ2kht5wNhmk9Q32f9aacpFHT
9Qxw86YhCCdqV/QLMxGp7v8bqI0zKTiUrUmTPL1Ni5ZoxaIk69NyCg8pnMEHCjZa
A+JtoO12yOIrNtaqg5AhreSOHa5LKeVbI4oo7RmIrLvAg4hse4Yp55MfzN7tBu55
iwwtc82ZYGFsI9aS+dUIvIlmD2DjFp8QPQkS2i3XlV/MdXpRpEgUH6i/9v7skfs3
YEanT8XuPXbmA4mc1Hx3BC3289q0C9mp9L8849GIi5xSY3IObXQWfyBSZfliwpzN
cAJP8yGZjvxfHkpqlL4GwnofuUpX7Fdqs8+JD6dRsRE3VwISYRp4vn+wrWg8DFny
QZD8YgkmEFhqMHKznVOJUGcRGIoj/4jdbxi0CGw2awptubmKRlISouwW88PCfdvl
PZXsgTxffF7wImH/6bXj/EGdbPdPSt35apVmESKKHGMCdLMEDtsv0wZCJz1hweOX
gPYIoYGXqwlcgxRDiQ96VHophEpysdrQqid99Kz3n9pNpNxUHH+2IAVmGNHpYkRv
C+b1p2OqHOzGkAXaYRiov3s2RU5RYAQctTVoopmaq2A6uLec/e+YZPWZxPECRMGz
ARKlzMA4s2eRxxKnIl/j3EsxS7HCZ5MiwKRfWT9zuo77D0AckkArrJd384sKxDon
EEHLQjqSKHPfBX4SFATM7+GdgeX50itW2lyREdW/8IES6Nf3SjYa/0S1oX3VXPkk
B6VMGboCwQQOA87KjX2LabfHKC125fJEQCfaV3F6QZrjV7DCN7+aRJXjjqIWfw6w
SX5ibExRC074cPF1odSudfgmNP4GiD7/eQZME20jp2wKSysDU5Vb5xhQCm/j3SX+
Ic4dx3BxP5RuxVDWjRKDCx5Kh/fS53keCB8l11/Q6ojvDxaPKEfQzWDm91YhdbpN
LWEGFR8g3ozpPNHy1e01S7ilV3W0mOnrw8plO58rHSc72gI9TJgiIMZbU46s8+wV
Zt7/MvqmX09dMeSrcFhHh7DdxWgThkbolSeJKF4Hupotwd72PjGrSe/9FMlx/9vW
aL3YDDdWVdf9L3ZnyVbBwJRlygXiSJCZ/4/ktmeGpmpEMjzOUjGnFAvkgLol9hN2
7t7YRYuAytOyOMxz8VNwOkn2RGl7+V2kbzKD4wfV/YiZoqrgtGi2KBTwyGont7CI
Cyz/3CALAShi4JRHE9H/eYmmEoH2Y/jQItqFDArZR00VWAxXANrB8HdCwCgW87Sy
MYaPl/lKhvY7Rc84G5lA2U3N7pZVi/20GGyfpt+ksvjYoYLtFz08PeSDAXPMW5HS
vweSbeCB/ssTA1HfjZbOLOEjcBa3BW0e0vJZXfCM4ehtBDL2LJSkz38CQBHF+MXa
jPRjKzRCxd4KLFPpeNf6wTrCQ/ZyrMZRF5I9pwCe0KQ46Nw5f/mGDGOYORFEMOha
UPohIbNt7Qe0H7LB+0+v1zDHkXXpfDa0majw5xmh9cu9Q5TN4hnE/n0lnByPkWnO
p97FJGN9rdcZTT8gRTfSv57T0bFRDKjRueZft2hGhkFFJECtZGxhQqdngL0YKlRx
ELdtN0XjNGEJMOwbpMufxxXJtEawsJCbWAOvyN4BnPiyGHxAt2ZLdzp/+/cFRKST
ccKyn7hFuL/UPSlXNYSuEjCiE/zNXqLQmsD5h6aPMW94Hq1XVqGVhrV2NREprYQq
RHMPAPMRcN9S3+qlrj0CDPEmhhmbK58yi67O46slofvd80c/kBTwIMh5b5lERf7O
NCBgt0Ab+S0ql8Z8ELP4ubNaypb/FIgsRcUJPwo4jnjim8fKGsvtjdRk86UWao6R
wlQwvAzLRMawPkuJ/E9FZWBjUf/ENKPkWuX1ytPISo6HTWNo2fsw3wwUqG7UJFYf
5FVbaL3ZZ4VsBEzKJ5fjDBLj3rpnMwm31vD29hQyExY35G3HBgQXlGZ6cLQLNihK
Ui3H0EpKiG0+Wb6gWpY4x7X/Z2dH8zTVV0ZQfQzBfI5skCY+2tmeeYlrHMmB+Isp
VQZIF4OIwcSnpw/JWlF4Pv1Cd4WWxe8gaFXhigdj7tkLQLx/xqUB7N4qB5iPpxCp
xiNAEwA08jDNMLkHxJLaBjeZq3Yb5GGRy77hjZ26ynwuPsbbA+FgRGiZ5H6UigvT
3SmsCU7DjBsrka8EZZ71qitTx3/T3Nsjql3sC32MvdXE7DtbqwSNrRyURgywPbxs
/sJBTfpKN4y6WaJ8AJ3qZeMOjimTQZ9lg0mgnFydrmKZmRIhIMKKgoAiUaL1XHQY
r6BlCYmG8SA59HqX+j/fwOqUGzA+jyM5WM6FVF4s1U9NpXhpr8UF3FvNOjmTuyJ3
wP7EG+OUtQiv5/E1Z3VOhTXQXeVV8ZKYeudHBIBmbOyGjpf1IXMhhaQ6uwU357RH
oLTD0TTPC6fPXj5vDC8oxvKr6U1x24b47wuYwd4ACmBaw+rPKPRbEMwV4RhZd2xT
8LdUmU/RUxhMsTz7Q6fiV+ML1OenydrCV5WkcDaaTScEY/OhbBSL4NjDMvvWvVzI
yg/KrwWO26jdRUigX7zSrK/Jba+XjiOKYHr4EdOPF7eot7KNzWjHc+VM+zdbjMxX
AMbMqlFcap+UcrBveP3QGKq4lZQbW6KL7Kmn7RdYZhfk8Prm8YAwX6uDyI5Sxr65
EAObRlgH0tcD9vbpG/ZXXtr4g0MaGP9PxQmrdttQ89KlukCWotpUkG4rKBqWVNd0
Zoffq6Wnxvdsg5+BrR1Hnkgt0mvoMGRJDN2dMLjwJaOa8FXOq9EZwIdIAcYJO3Dx
2mrg7zNBgI0EQVLbSiJvOKMsxqXHts86LSYppekI4RUMkRPZC/ZadsiWV6pEYwgK
TLPFwvgqoqqHVNyRTPq1e7xPzBxaQyvKHd+2GiTEAoohfbVCOVD7/vJUkB9helay
/7JJ1RGY9U7al/UAvqQ83bdURcPMKcxcdyuVuheiGMcQlEDPLRMyWDUiO6Kotg4m
VNT8VJTH+Nx2KNBC/GM1lseCdyqP7nKMazExfXdBtTOg4lND7ywd1IXcTmYBUdXB
K2Z52alAi5BhEtbYLrmDtzrRuVrXrxtvjA/T+uNqS1s5+KHcUdT/gwpnMzl68U+i
aAlYZ9OO5VLC8ZEO7mQ/f4wn5tTrcZSr78Qsy2RA8AFOZoDutd41ojx8padEfMF8
i+3ad48bqhmg5+kDpj0QgsqGoXMDGZZKuhLUgD6KTqe2vdybRyRHCgz2f2iUSuPt
LeNnn5Yj9l3fVmLlwhFWbhAv0janrc4RPRFT13Ze+mpazsi7rUDESq0ar4BYd6UY
eFH/uPXM77wBMHwDgIk1Rhx/Pw3LhUbqpLsPm+kmXICY51qlDyMDTLa3aROw3rfE
9vINd1Tay1vGD5/gianqeUbgEF/7f7zTOwC8y4t3bT0wWs2nuuj9QFludQ2d3Y95
WwWlJfcUSDwyL4N/trmZxaGyFJX2qVu/C/Tcjh0nlF8TZ/5oWsfdaQ2FjkMeHacN
HlbiLDxyLH1UT+KvIeH3bdMboODR5BnsScXN7Q3fAesIk+CJq3bN0IvKvUGHwGJn
L6bXHQaVGLTsto8CQyfZPJY9JUwrVNiZlh5BqQ4nPSrhs9N6KEY4kLfvcn8vEHV2
mYII4OvYC4ymYgQVlzOlWTJw+7Ip5ecD2fYkA0sLGFlXVfK87Oc9etqMqSgrSxjt
G2+uwRqO5oIHAP6T/8HEIuYUPpYk2zKF4ZOAX3/Sq9c3QoU1SPiB/zAtWsRyfRHS
tdPO+ohzfyaj3wV2eLjwW+ZaaQ5HwBiuAwln6b9V0YCYSN7T/ZkKWLyK3PILyi0L
JXiPJ2tlBkfodxgtaGuYye7IAAnUlSLK7rPegOfzVERzxtyJB1kwgmnItr3vbCTy
5PjVWcmhu1MWuls1p94qcVChlExdFOzcXOF4AqSBbjKK5xFwZociJppZJtcGb2V7
7Yjr+x9IuQeWniFJYMqXv6fFgAu0TylvxgZDhGObXTJowd1GuDRqi2x6mgS9WVIS
iK+8fWACLKx5kYfHoFZFTb/j4TIFAISdPzjNzMvQuwIDaNyK4vB7GUJXzQXhgvqQ
n//Vt4dAPDpYz5X/Ne+fY5MnLACGf6Et/WqOHrZKySTkkaQhsNsUuBoStZpT3M8b
NPtEh1o1pcEhsCYC/ZCUUctGUyNcylDW3SLdL8NFX6FUwBsfBZsbxEzkNUgNx2Y+
ZgBLCLaUlqnkpRorTXSVaejthxnRaw3EJHho8vPNIbMjxFcFGi2N75czWFoL/Brv
jEpGmVFI5xdyfJC7jDlN1qqt0bF7s89pqEhHSLs+qCtD6blGimVlOW5oBohTOfwU
QtN2R699phQmQ/MXpSQFu2HimHPlblN4eZVsC1OtxuihrnpX4cyph2YnxaHzaxrp
HBCB3CybChHKO3123KdyzxiEU0hv/AU+0XfWQicf6cvkKv14fIzFWb1BUAolQX+e
VBbd+zew8qVH8UwA2i2lrzGecSzu8S8eRMRJ2uoxhi2p+31NFdAivTGMZzhK5b6Y
JgvLS70qGhnV1lyWkanRGY8yjCe/ulmbKz3Og8fwgbnfEPynGB/TC8LFjOMAtOqE
yS+M5EK1BGmhk/jrKmzUtNyfTY8XLwxHcBgwgPEdz1qhTx1Ehj9+1TKLUQAylCxP
qbHzaz3TsuHI4bqXhmcMkdDmd8AaV2yKCY81+0GKb9cXl0K9Bzd18JE7auglSyWK
ms7zxawj/Mo1I+D4KfvS/MF6egtJPTbqCMMzTGQgR797xEIY5MjwhlRxnVoXYiLj
16d3kwgFgGOiiLzzFXuzeXiDrDaeETKpKRBUrd9VqawC5G219TZ3mGU9X/7rtxt8
CpDWTUiDPFhbKKHuakAe9ddhczhDw7TkQrvn4GsukW3ckzUV5o0JRzGOjG0U5hgj
A7RWBWFeG1WKgTjQsv7TOQrwFpZb4Is8gZ3Pvk8Dt+2aBP7WQz07jb6FMuLjLafi
xZhyra9GlBb/18r3AnmO7gu9bHCRdYpjmzzR3a8hVzHR3mL2BacrtGBpRx+hw42a
dT7WGunWb/3bL/Wz0bXJNlzfIbOdBEcdnVDYL0aP0A1X4CVKRyHWlZsCglB2S+SR
9v2bCv5BjPxmkgrAo/C+en9k448OivackgSl8cKbP29IRDZifpZbNDEnx51aNg+Z
pDqbW7rOk6ZZQKv22FCrfpJyUVk76+WqK1P6n1Jik3jFboji/6mF9BGJZs8phSYS
q7qLFQ+8ui04EDOJR04N8kdgzyYBoM0ihyIByA06uXZ3ukXA7T3WJEjej5yDOp3h
hyt7SLEYuV37gqD9SPhMCARhd73/JNNA6ta8AHPQhDVIBRmQkUZ271pLUa8m/ykU
z2YymULhniyyLR+ItaXBEoLJX2x8HVH+7los10qBJw/a6Y/e8KrxfOv/OtsQZ9dQ
sDwrOBSqvdAcK9dLbWXlMNsjyu3tRAK1AEjd4RQfIHp+gt/eQa+GS2IjZ16ka82z
yTytYQPRj1pAJ0TEMWsn7CCcVavrMwbfUZUM9uULBEYOj5B9yxOJP3sGj8MupwFU
7IGnFScVYYdSUGRyQDO+lPbCH/Yp7aq+BlcU6qTfLBsa0FmXodNOtw4DBxQq01Ui
xFDCpGsmsiWgaZK5DQHgun/O8Gg59yjudqudr8EN7PH8lumlmgIf5pRbkx1VLvvm
WEkpygWqBR3GeYrAcrZZftK9ikdBQL4NvIz3fN6trmulJvx+HA6jFCJqsIqBDp9w
/DW7L6DdL78BE8pKlt+CFSOeQHzlRN2m350NkKr6SQe8biRET6/1SYwYrrN4m9be
lRecnpYHq5lHlRgWct68Hw95hHCm4qf4Zr4sr2kwOPQwIKhCt9OFUSbBzDrGH9eV
+1SEJ7c+DPvAME0qHgHO4waafECg8F3yKAiXQoeP/1y1/Npk7h8JB457Me3h0eJC
Nt1GJp5yNwG7OD8knYng8jvID4+I9Frsae9noDorFJAdl97e26dEnRmDCC3NSfF7
1yqMcbQbIt1LAYsao3oqvQL8VBJ4j6vnNabmwEoMLPVs+3S6KrEiCqU7L+d120Hp
CiM0lAPdzZ+KwhmU6QklCx0+o9334WNiJdjFFsYQA4zvG8EhkJZjNxSJYezp2z+Q
BJAay7xeD5mDLTqgjWCTJig3wPaPaotb4aeYvmSM5Z8P0zmrDRG9eOM592jLgG7Q
XZVO1v9zqUIYFXEM5RiINg76cPTTI5YQcVk0tQkvBDqaBUmXUpdwPDLxkfZ2srpL
jsOEPXLducZofzW+mhN3lSJDHdR/DZU3I7HHuwcRVL5uvmihGnn1uTvgwzc8gmJt
lXPigk9TWv+a58KEsgyUyEYOqrKiHgw+/PH6rRz+3ke/Jd8J3sPTu4YegLSwSZhO
8LTfVyBpKP4Mlb3q/u4F/b6u3mH6mxfxNiG7pYLHCgr1pufP8lHWR65jH9hHxcXN
Pt1gcCnHTP9ztWtxNXvGIWBB9PDZwPI2LFSGti2JgDzRrmiLmJQ7FaPAPeqTswo1
+hO9BX6laTKkQrIoAHiQ1JjeJ8ka9/npQg66I6hX/ANg5YjNKFWR9WlFtDhDEMNz
hGRRQqpeJHYZyt+7GYZzY9FVHkx0UmoFjMhVdDCMZW9Qxpnhy+Kls1vexEvm9KAi
TKafeIM6+t4Hm9rWv9bxjVmVV6xej+hjH30QvYQSQv92zmaF9iVxM+NtsMW1t+X/
ZHX+3jbB6KShZ3918ph0y1LCOct/2+kCcK6yoDKloC7xsyCOz0KfMzrBeO4Eb6rY
YAB9/Mo280+u8BdA8tIcgDNZg9AQpPK+ovPGmGrH5KvleIzMxRvK1pfESNcBFEkj
fN6/HS5oNNLXtjWNXeVoTYaxyF0JbSzk6/wI/n2s4BvlixoVCW8URcAQrzft4O6Q
sYizyCXmwC2fBwVS6oXxOv74FTWSND5saFb/fhb+KgxoBL55Iq3l0Dl7xKphUAaj
cEgEsC9Za5Zz/1wcR4Gk1zAamnQUpyrl+OJWSmRYgTWvg3jZerKut43fXRTLl9xQ
Bj/QDHjfEC+lHPkmTOPc2gIrmZdz2H5KITp/crEJiXU40G5zvN3JoAD5f/JcpYl4
rdeY/OhGuAfnuJpcvhtBztwaQ+CD3Ztd4/LHAmPn2CWHKNhKaoNncs+3+2g1OUlT
tAqLRj87BEVlMHr9a5QPbF+n0GbGBzRrvhBboI+nhVVPpTf1bEM7B0MfEtnTHQ8o
iRLAYY37rbP83MoR980+/e+iU4iCFDr6g9kvH8oRgIADc7Y+xQOVMr1mIujIgyHQ
vUcRZyFXTdsVGG1EAUZX4j6XPtqHAHciGDyB6qg05lkkmwHM2ffgsLdqk7hwnvGm
dhFUFp4gwpcp1l14YMVwEjuU+XfvY/Nfh9NDF2nUeeiuzOv2FzG354EtdY97aZEi
N0oWtIU84SIHy29TAee32bEXu15Yqsw1KwdeVBzEyzWODwwJFdu+/HD96Ul9RavI
sGf7MoPsp7IjBBrwhDAOGRyZFAsZa2LEsNaD9RPMhn3Etlac3jG3n5jzA/ey2ZQU
IqKxP0or7JsCd2QAWnjMkI8A4VU9ICLXkisaEuAp/kB/UUQm5f+QinHnqeXf0e+J
tU6qPX9DUXL1aeW1D7piE7Z6/ZjRkz0BUrZvlkjqUIJwzKv+WHvOILxmnDvQWUyD
VSJwzak+zSGgz0lU5W3VwLCPpEAa7M2Gq4FUXpiOvh7u6wlZjoc/FkWtTDKA1k7Y
45qWvLWZ0kUVnscM32f4EpItlaUzjegW/HtOmSsvYKu/ZEU2Es6llUJJM2oyPlo/
512dl6Nag5PlTzzKwIj/xdbWo5tsCfbUB/8JFzdG3ZzZuptsgdxco6Yi1tOD0ZgC
0W0t3L+qj/x/H+ORhWQBIqo1x6j4MC7n+sPQIphj0xbxwNendEROgJuik0fFTtZy
HWC+iQH5Y8UDP43909l2MQMZmozxn6Fv11Ckmuex52XUoNHypk4XF5N56nGqJXBq
tlsI/tQYSFs24fnePQr6+F7rVZD0ZxkyVsnWm+UZvWCQYAgShHGgCgJqoTtvqzvh
HnKfAMP2s2Tpzivu8FKPlosuwZiE0JEB0FVTHBt8F6MYaI+1ZxTcfKXIg+/8iN/7
Y4M2hUBZXCUKY3+m6DsaY9oNAmNXrxJEOHdMyzaUCk3w5GEtWMElSf/k5AZo0MAR
ym7zTRypgC5QrjtMreI3IYoC8WOpLVZgb3l7nVGQZj6CE13aUtD1x1jvszUEr0Vm
gGH+XCMSDgSgryN20nudRoAU1UkuoP94Hf0kY46Ik7qrrwhiIuKJuJZah79qekhv
EPYYA6xoh9Tpw4X5P7gRMddmv6F/Eqn+VRxELusLshOUHKZVNlZ9mCG7VlY2OC4c
7ZahNlySujMBqzDwC0es6G+4+UMCEaP1BiONhczspJ5N3datfGPstntO9C1/T1Vs
pa07w5ssvy290WndhLHVYQEY87Ir8v5IIKU6l54ooGw1oAsLhzoyE8PJCCGbtiNt
LzPoqKPNwQxQsuTyXBiCl5dW8XuRER/U7V3Lxa+346/QYwb0y/2ZDyU+ik/B/Y8C
zWz/Lff0ELDQH4X0ZAjfW6ww8pZTDbAYXkdoFdXPiqWVpvxOcmUOEApxPzG2Nhdi
DVIEeB5nCkAYJNRsJ39PJxvZcKxDCZqcm8IeIOXHYEu0ppR9zOk6ExHOy1nJsl2g
JjjBbHohZPdJEdk2Nq4OOCmv3OueY/CQrAU6RsS9c0Hqt3MfAlDX0spS90kx/GR4
AL47eUEiMoF7go2RMS1e5i7tg4lnKImsCX9xBK1HP4I899nl350j3+n0C88kbyPL
adoOUSkzKxc2Q0vhSg+pWDL1fcmmuV6iHxo+lxyGpxf5uJ+lkac67kdPInuvwNTT
n5llPoTgxu+voA5Zidke2q0hO6KKU+kJoISZueoaKxNzcWMGTO+Yx6h3IoM5fLGi
/QWtYB3u0GfmURlovmEarYDUz0YMI7baMDJslb28qMwCFu/86xQdaKTWWzPnMIIs
8DF7noBKXIJwEByBvphDS/4GkSHPNRjjgVyIIqf0+9yD8csGQ8S+yrDvUFT/1vwg
gfDFkO1QxMHhQg1tsIIeDogzDSJ6arEuQae1ZvViCVWxieS+Mwh/f1CJbu+fqpJ2
UKp9LSyLpjZ9oK6qKCc3h/7bKbTtv1KV25KYWA++KBmg4zDcKZj2dVoJm7oWMRhl
D4BvtDokwnAQH5hvu5u/fsOdPbwZ5WXczns4eAU+/ig/ITC8jaMWCC6z7HS1D+yQ
zXdGDXc9plSUSNE+l+PGslbu8TmKmuov6M+IJRnl8qICA77HzeMz43ckHjEbJu2M
HXqCire93teFcoQ8HuOHFX1gSDx8zC2PamdgCM9cTEdqORDFgw6SRqPWAhP/4307
A0CSeWNNTvByoN8dxsczYhpDgxu631QSJQO9Fw6q/65kzO5meaqwPx6TZ/QJ/eL4
BE7x8ws2LCVUKDQgSaUB1QV2Bao79KR3qZ0p63MHRnqieB2LQ7UzRKUKupNePHfQ
fyOYgG/1cwj+qNN3nV3/VWu7zBn2bs3X11Nnedu+7PuwwfENcNpcNd4t6lduPbQE
xsUSm+16cOYLAJ3hx4LZUpJeBPANekTCyg9xSCdLcJrnutXXe8To0r6PfwPIqzWB
DgYfZ+b+WMT1G55g3E6QDrORgdsUwXeikzTVH9CgT3lZzLT53cEVzM1SvnmrTx3p
VZRdcn5gZyiVNZ/awfdnd8Hw3nD86M+1mg7lKRnff+WR+F6h/o2hgMqBTy2/Ub0o
7qEi0Up1VV7zVYZ/MjtNJ8MuxheLl3Kol++/hyLiPGKHxnYKnBj2ZJWXF3t3ALlv
ICmRzmhRK/Ddo46/pt7czPFuYwNUdthPMI35ax0IR9QOy9D1l9Jh6IQx+dxFO5Gs
gmU3NHh361ZeITzyZ/1XPy0aLTno7ktQ6tJ6d4QCjoz4V6gxps99XWYVuFR6llcl
T4KYo0/MtletBow88FoTdbRbJEKE3yTXRhhU7nLabkGOQMXXuiYjNOhIJTERxzmk
QCpmO7AHRZTa3Bs2XKURVbRUlxO4kVY0Fo59kWn5r6jOuaVCm9l9TwUuyLcBDyN6
XcRJjy+6xJz/pcqLhue7eayx27COdNACzsEtReJEdhfuCfmEXeyPUlFgJr/p8B9O
G70wWE5eMWi/LvpbWvx/7BPqnFUYd7ClIfbKHUGaIHRoCCSYZTBXH+jYmMOBKF/O
bp2WJeN7Ty2jc/CDTlvGzooLsOMdO+glLpJ367Fu7ckOPvAZw/oUOX3QZFgWiFF9
Q/C+uoKHIk931BtXU/yRDY1eNqqMNQ0ER0KS2feyrTIOkz5DVqTNJe2zCr1lAJjh
iR1ftkLZNuFnTlFI6OwoxA+yuouwrfpTGiHGn0115t9e8cHfEdPTHNX3sYmsNdFy
BtiNQAYMLVokbOzyTU1/rdh+ENvo/kQKbWU933UUQAjyddTXX97fSjGL9WKUyXwz
JHtRXWOL8BnVqxUJ/zhqvX8ELE1U7foi/isdCtQNoHqTidpGzzW8y3EDF5Ro3T65
rOSvOvjR5rWkkG6DAP/uioWqGUy6+gaSE5O+pggDMe7DGle+5vowTCoW4qDp9sDv
H2rTOrRVzjPF/ZYpnm4wiz9BTi1/mR0fET4UHOl9dOSQiF0tMGSqsI9F4ng/jaAp
zloFSOeWI3J8MIAYaAcC8DiwY8dbqXTqicQvurlcGyK2HO54rTAhffBdAq4/hhi9
Jvn/J1sLrrSB7ykEuZWhPnOLsGP6YldfFhNncXv/QngHCdxmIfpwDbnW49mIXMOj
y6xsxulAzujAf8u8ksW4l/wx4XmuZQc1br89GDmVo2YUsSkGXKAdlFuQgbh9MFbb
4sF1NVkMyCiWxpFZEFGgExqYl+rng10/1zCX8Jz/+dGpBFtU+oyX6W3WFy24tmH9
1/hajDx3f9ISYy5DA6LoI4sOPZ5BCuwu/pwO/ymY2ECJsZJTsC/o02Tthgxytnrm
9d5iNrxl8h2JivsuFA+5XXXpAaWA26mDcwhEe9JTtQhL2ipifGq9X0oKPR1L42F/
vYZXNePaoQS+JBm7W+F9DtNbdTHf5QMbutjcrn6/w4VvgFkPxTIDYMGni2J/aKcb
0aP7lKJYNAbXfznJYdGYuIZtSnc3y/yHrosGkQG2x/aQWvulaXUf79GhPBvvy49o
JCXqqenkD59YA8X961dectyW8P/rRG0B9s/xfB3SWF3M5co9nZG+EKr/K3EvCCgr
5SUnAFGZB/YgXlHDjxM6GF6RSa+jt4Zcn99l57ql8Nryel9Yg7nl3iwck8RiJh80
K5KrNdBGP4ri67Lu81HtzmIGuA7zOuD5K0eLmX8P2cHZ3e5mAoC15omdU+dwZ4fm
Gu1Dd2vOmfKUm3XlbkSEj6HKzLKoUPcP2qoid3cDzvNGOllW6VEG5mimr6hfxzfc
6OP8dWGoYJD6fBfR4jLfuHKG4Qq4p8Pi9HNGF48A31gAzSYPzIrRHdAJX8pN8oXg
mq6MgWHYUr0CoBf/z8MqRbPGWZPdzr9dZzYdWPrquhQUMlnhGQlblGRQ9NR7PtKL
O/BVsCr0T3kiaUpHV/GTQZ27l5oEmcDb25QNE+Toz7BCUpWl3ClYpcRwYgRoDMb1
LUrSxaqkDIErP36kf1C3CSLmN42ki7qpUXQ7XKOY29hTsTSevQB+EyayNPoEUiN4
j4TmgGoWbue965txrPqS2Rfx0anLtORVJpqynmrIibuTuu05LxJ6asExkWRd0SUF
CXgMrvl+4O5wZpgwMM3l3cAG2vYnM06hajbg8PEcxRzSHsqmfrM71LCycsOgVoIV
/r5di44yMgtxTlVO/7/ur0/vYHlJtLLiudhB1DGE95DIDwWQTQYyT9otW4umCxsM
FOAdyIeqyAyMOxPFM8Hn2oAz8ytKuwTmhSDJmFNx6FOYitGUMqy4LnnHRnTgY1Sf
gmZjpGNRAZZK5z7YbkXsoc45m9vLB90DOJ0pH08ob6ULBp8fG2QPE+WUkOy9wifw
0jyhBVw3TY7e3PTqx26u6GOa5Rrp+mlXkc+wvMqIAy+nJZCnYvUIAGKxworcamUO
ouGZbeViE94oG4Bsq9mcKkoLMKyVqMtDqcQ5cDHkI1aJI0RuY+AToTvZj06cJ6Kr
iMrNaAq6rVnnf/iShNXaoCjNuDqThxuJdTMD6g0ujWRYYqSLs6Xv+93lSdgpNjr4
OvmXJiFt6+61JiAEOleJEt2rbO1+UxEvG7Z/zwRLU+WMeRUXoXbGaAFgUTxy/lmz
EYmMrIJsvOJOuZ046T0GuPuEDiHSpH0sCcX+P4AJFtMlGUSqF4aaeQy0IBrrJP1Q
XIIngBbhVXC22NfSH6O+ZB5A9GcxotXSigySgPi+bq76mZIN8qtitPFBejHPnrQy
chVn3+2zI+2vCk7s35dZAKOz9r34BI4kjVveE0bZMGG6/HBQ8No4xssuJyzH0MZP
SdLoTb/H591FOZUt1qvhlHKKrMtI+QFrGg7N4J6gkAXZy0rP4xy6ikD2TwE7lehG
dRTqMe4QguqmuhuUgDzlBzSjbZVP9hBZpjAAQWHbG4Bdn9VE3cELk/WGBemKGL1i
AtBJQwOkcUiiOVvbACvca7W8O3ioObGw+PDVinu25WFYGMRQZ49nS8xUZrF6+g73
N4sNra7ole4HHwgjiY2U+3SrCKjTKOZ/CIMD8V1Bd2afJoSYUpduv8rk58YVeUud
oa6B/E8b3GWLe8GkT9esiWTpdf226G5BVQNbB0VOGVyXjpYwnPWTDzqUy0EFIAzZ
1ksF15TpIibLmI+CWjRz/2X25P9Bgje17glMvnWMn83usIzTOJ1dzBwwCLQYxPrX
16+lWPOc4UrfsGc8mkh/bjUQiUe/kWdzzHW6cK5/KGz0KvagZmhJnTze2re2Xhbu
CGEizxM83pVQRve4uvSTT7BFQ5OP5VrfiFj1B3PkWSc3pFY+Ub4dtZGsQ1qzrXBw
2HyUtKaZW9yJM5kQC8X9hRpOHw+9uCWpuAIgf60zQg8+obzz2NIaze9zJsF3Sei1
PNjPelq1q3mjI7pAKLsuB0olDbSI62lc7zrvNFlG7Arilb/Qd1vnsM6cq0MJvVWd
aEWKwLf7EHFaPagzHIi8PINuiNcQSKsnjJoj0+Vj2znROCovCNA7nDnOmVDXSIf2
0Sqagzu8NaHCjjg2UMEhBi3ptDAZOsQaS+Fetp+w9Z7nSapwyWzzF5dgSCHLVfaB
OdTbwnhD3XzoXr0bWiSWZWtnKcpxTijIzkQIpjUrc04voTX4Xa0mMVD/EKghq1IX
Zjaomkj7OTx5TyYTKOCDR638TWeb7wJh9dtpQux5hPCPbzP+3UgVw0pWmSLGiJK7
qxWjjw/k5SftoCuti3x//ZYsjP5c/gLZ7tnTxW90sETiatJsaQtLe2f1l4FZhAJ9
UdDqPnVwrYeyVVAPZM56Ap4p7Pihhs7+iBjCHbrFokCP56J7V/KGVGbA6oBAFOMO
JUbr3aaAopiJ8MctQ4Tg2hVyhVw+iX2vhTXdJNT+mNJC9fwChG0Q+h0EJrPRhcHE
Xf725YkK6c/QKexoARggVaI2dgXSeQsKLfjx/7i/252lV2MAmt3DU1x3B0pSvher
QxxPb5RCgLWrmCc/0SaFpYxXt8vb76YHBK/7pF+4Z9/OCZVIFGSJ11UrwEPtnYHV
LCjDfdhSpY2wT/vmH7IOCx0uDjurSHJs7Gd7UMHYdqkhcW66OejULmAv3E96vG7r
ObQG9tYE+1LFPCyXiDMUfurO16a4peDcq+3lHWBXlS+ZTsjGI7IRhT/EFvto+be8
BumxT5LvYeqnz16JLUnAxJ1Nw/myXmYDBgAOxbKFaDC1KnQZpuSlY14h1LZgsHwo
/+d17lUYy8LB2plb+Od8/DyFxFEzuFZXoo/QBANNyJVotBOrgX7bsdxdWxaDqkH5
N6XsdKO48ji67GLeCEzgo1r95DLmcnTkYg1/ke/JfV/npQmb+0HDjSHBYUEtMUbr
wmciFljPOBYhpQHdp1VZpdhkuJwyjcIC8lASPSIgeXdKJsIekSR14V3imEf9TNCI
hXaWjUDbtWzCgcXIo25TzV1sJSFajtk+STaDSqJIyf8AatP4nyFAQR/xy4uYLS3m
8lgYgDb4Q6fylWtkWDa8SzJpMTcnl2tu6uMYenFa33FvtBwvx6XE2m1ySGXJ9S7d
wVaf5PEgkwrHeKNQilfZ8Ycs/K5Z4Nbt/nyVQ+dh5C53zV0+qTGIxYb1sZ5cQYz0
a748esD8n335ykaMU6pHTPoK1/zeEHE0pLsEZGCIvgPhoDizsC6HcubTcOj0wAhR
GTi0MgzqnW4L/i2Bbvp2CcwVwCIwB8RboiUAkSDbf86YjR+fs3KbsIWV8L88wiCH
12ULiq5kd8tjlVx8OyMWYdsLuAwe7Wo409JTsqkIZ3yzb3hj/k6ZFqD6+mlANa3S
bA7+OPePdcivKRKi3LGrxxdOe4ELAKm2Q1gc24Kvsi7jPcMyvHZ0z36oTYZeW3pz
THoKOeESzAXsvHCghSeNFc1YuqQ6TyE7qbF7m6VoYmX2ISJs+K5xKO4H1aLXEvWr
WtbfP+woOduVH3BSS8IqACknnd8kIaeNXc2OEZNsmxh+o/3aYM0VgyqKt+Ntamhi
Fzyj/vYMjmxaIzp3fKG9Z9yXidHtek6BmvYVJoJjBAlubwglN5PlkfRvwA2GTyN/
sm8EoMbIDGfa95uyS/EftILBphMQx7J80hN0EkzEOwDmed7MFqcyus+Dwjoe/vC7
Chs5hegQ2J0Iw51qu1qmZfDwF6XELaJUFr8rerB6t6jueMSnyDliZqafY8z5vuGK
8qXa8dX8rVOdy/h43bjGh2xvfRaayOCohIj/3QdR3GE8U98d7a/5j/HTbFf4DYSU
NE1jCyZa8nYELmNB9FSMTP+/x4X/vQbZ1mO8R34hxHI39XdAxT58LL3Q17LNnmfY
v/m64KuwlVXZMVF1dbIsezE3UAOvhrGOgiuUUqkEvy1xIWheR9SRIrVgddwTXaw7
TKC9XqZLoJHhjKQggV4Hgny3ytBm403fMjBTljmJC3Rrl16AycOKTagmYJX+oJdR
q6lSbKzQYEtBEa10MjKaW+E4li4s5M0emNQcreeBMcHNUP9jiQmtzL+9vjO0gZ5w
IJ4jpQNvkJNMSFTYmNgP+4uYrqONuTLWJ8Vwiy1rNixc/5KhvFUmQVaLCS3CUzGi
G9n6a34AFIk7kwAk6/h661Wb2bCR/nD6M4Dwz7h/XxnOVHHM50eyoZUU4KIHl7Cu
E0pMENg7qW7Ij6Qtf435DwlhMxat2UZlfB+p35NasJi67aBCJgWu3tYkdbb6p+PK
YoYJqqJG43enDq+erigcnCb4HCBpk2cgdg4i2GPzAAQZFqXrO4dLC3XDnBJ89EoZ
bRj39+ppGFOdhvJVirPAkshepEnIIeIUL/VF3PH4Cioxb93VNt3cdHYeBY81w3Za
iBY7cmRYXrsINm1a/FLz0TiLvF0LEfY9rnw8VGbf17O0/SbpCARmLAa359PLfyrg
Afw/cvr4+kMGPlPtxRCf5BVCW1hFOrVw3c8RHD5Fz/MUMjaLGGBMIBczDQ0cg3ch
VdfpDCSj21SEnoy1GB4U9Y3PvxCduydr9c0iKoVstCtKnVsMRukfhu4hu12gDZJN
Ld3GPc4qifISZbwZHZldqLz5GkwWkd8npedI58hFLWVD73aftMGD+F/zeUUWJLp4
hqG7YmzMJORvj+yqAOg+Hfk04G9u5lmKcQNIbrFyLfFPhftlTifrs0UDH7OOft72
5YDWbM8enL5ZUws8WZplN/5zL9mUSxTmsB3TE3GolpLyVViLlgFUSeXNksAxKCCJ
IQGLqeAwmYvvvF+QULEZwonjAYnF68kz1BnVQBYJ12pczQdGf+gC0lTyVp99pZqk
0q6DkW63MhmOZwvgmzUINMQ/HPshl3+tRIaM5+3DP0BLk4fugc+Sgi2RREqtDOfM
aAbVD3FHyW/d88+ltNaQvIHzy1cZah7VlYtpYhfLNnuXW8FuuiL1Hxyx7113t2TX
Po/zA57OLPjNK62rwzdofnITi1RZ2D/Y7S9cer7ZvzU091dqLiPwcqV39jzcU9Ep
nmEA1knwwoSdvW8dKqrUUjfjsqy/nmWyfZRL7RFX8/G/RDdc9VnrBPJ24dWS91p7
YhWXTd38iJTuupU7i6Fwb4MaKtrXIMUzbcjEQJulSzyyg0a34jBJm3LO+y4bR9ou
Sa4tNyFD2tV42s4nK3h8VZEkgfs+5UV9VYCQkUDecfbXA5nySc3lAjdyWE/970mM
YFwyQs9tBfidjmxJmGNLrRYmDk8ImCBK0dQNY+Itx3lSBMM5m268LJ60pTgDf0px
An75KfRaNNPx6mSuSt9Zduq9GybX9EKpAVsEWSTCfXVBBF/GH8bJtKhOU/Gv2FS1
2UgUH3WKE04hSSWqyEIP4Xsi5pIvNI2LpFbh8RRZPtRVrOyVrwmgQqJfIkFubosL
jWiVE7AxdDyAtEdQEbDngfASVL2VhG8S8Z8VEnuLOAv98sJO2Kxyots9c+iCq7Uh
Kf5abB5YyFBxQ4PfHY/a5J65cx2ji4L57nyWQs3iq3jOpd3AtQG99DiDABDJJKOn
ICKhT9qJxGCR4KPoWueW6aqqoLaMZyTTfGYdS1/3TovjosVG5MyCz5v1mMefo5L+
/tE+qFIF6MA6znq8vDNzXMB/r0rS1S7SnNwACxJOIotxbBurrPXIh2sgKQhvPSYc
aQDCIFWE0X15GsElw2zsUJjYLvF98kBd9H2MtqD//HnmgNSio69IVhHKBB7IoL1m
44BxL/Q8/kPC04xou0+O/M/8rZXs2IAKmplinWBXrLOnwsU3k3n4begdyJ7fb9FH
vicR/gVGvpKS9BX0Ewac4Qfi8yY/U6VFrSa95agLgIexoDZVEJMjMu9x7gR3MOUh
uDuKsMDH3jToI1F+Ymxz27rlrxGpzdYe7KtxAXtNwNyAiLbAs5ZnyIxQl8J+3WD1
pA3MXs2CJfl/qjI4GXQgZmy2X8MDxnxm1IoDbhYiLuPNyTVpWTun0+8bp1Pa6DSu
tOJQ8aTothHp2TDHAGq+n2riJVAb5NHCELJI3gK0GTrPyp9umcT+hCF6dHF2qXS0
Fi3b0Xx+9N30PM+nG+wl2p5/3omeHHckUHz1nn2uKYvk63nrvbK4mVBKRb+pG2xh
2603U722ZYQJ7cR1DTBsZUdu3/hsOR0+kTWHBiy3sZIP63Io2JRDXPB2d8lAxp06
kTjF4FApMQSuGX9pCLQ7P7S1qCtrVOC4VxoPQGqb1Ca2o2sSWrkk9LbWQRn0TAOU
FyFFFkjlIeee3EZWFeW4J3qTXmNUdXaCIrMtdc1BvZnQhqDsgp3sEVnHFn6EsakV
zIRGQzxs/KtkkSTpPwKbliS05obMLSYqTP/j40Wg1tT/5BSdWPL2fzeQfpcRHRBG
oVTseRGUJqdr89YXGpnRLvHYKEJoJU4ryq0J9TAGhbBSuk0ve/K8nrn+9VyRKU/U
8PvGsRH+y+G0pwAxpmPvZplO5Uqg+54anM9SLWr/zNZWe9furJwST2i22PezXcrr
bOPDgIRh+xSOD4It6hvCuW9U0ZtVpXDPKafs5zqi0Nl9ZW7vmTpJiYMMibVbtpcf
q13OJ39DwgBKQwbAOLvv2NWKatgEGCbR+IugEjlkzfK2YuaUBMRXanU2C0BeruTH
k1PYuLP8HFuv78gxQlH/QtbOOoE+qUfpBJFS+53qptOjLw/6N+YXim/WO1fsmse7
JN+xbdyJ25jLYGRwrXVqpR+ZUlE6CV85Lh1VfsvB04CdJbI4K9aE5UUCn/z1ArPF
VGggAT1iEQel5FwocXEKTXOJioqlvtX7lO4L8W15ysQhjo7xQxsRxCXxbn6B0m/v
k9PJZ9qaYf+xaHD1iRzsrNLb2rtB8nYNYoG66PclTf9+pUkfLVLO1cZK6VV4mB5b
l5nQ9iPMYMSkFbc2SUI/zWJ/IEMeMB7w9gD4QBorukVOMpRTb8UiJNszlVSuFMVu
fk0FeM5yfiO/iVUAwwsunyW//SIKA9a6Y9hxflyU4642nn4hkHDN4DSMm2mBmkeN
VCnbVgp1h0v/Ft6IHYCofujrxpuLSL0Bb8r/VzB6vm9cxIOuJwIJei5kqdT1rodO
GGO9L8lGWQOJhFwfLt0amldVzgZkw3aEznvMztSLkBVM02NCzeTPduxfLV6P9LKx
Cvqvr/dOuGfCYm1qX0kZtY5WoFOoiCKQ3vvqVW6ntMmTJQhuflqI+fadY/2bBKbr
OYTFWKYb0E4XywkJl+pijz8XXUSMv+BGHSVAnA/abL337OCIeKNHhqN8qvyF4r86
zz+32HS0+at3S5Sri908oyVxKJoAr8LAXxck3x2wP1IrvljyVAO2RFZPCbUTWqWR
/4r2Pbn+VRM1XPr5XeiR+2U5BzjaMta0Ss2VHwbblyDeRQ3KhJS65v1mGkrryefb
xQxwWhKOdS62MQEKqncLIOf8b6+zCWMUdPcCKe1JVxaUwFSrLV8tz2gM7Sa5ERH6
1szzeaflYBHfbMDTu5OBHgMnxJ8iCgbkYtV5gEASmdGtn+XiYNqnKQb2T6zloHLY
JwqnQJUFJewQagXZOKyZB1Ho1OonZo6DBegJmuMh9Pd3SCzhXoIsHIKmDY5jRNJh
k9M/M3L/y3MT0CVR5GAYF0hE3fk7CxZidsWtQLAFH/C7SB4Io11/vu4I0AnvNkta
9cFC4xmf/GyAiL9cFirq/NqML6c8GFa8dMYASQMOgQenZHcmtW02JxlUEwNtHoi3
c835BC+UZZGS1oxVCp1bXeFikNjRAfSHeTP6rOcPbbPj768piP1WOB2dcnIDSq+y
/PteMt/POkGfMkaU4y4G278SpSOIekZ8PXTvRHnD8NPhsqCUbhrUmu81PX3qMbty
ydpToLF1T67wAVOVyOg+r2N57a761Wfy8jpRjXbbQ0KVvEdpN+rDE7BSL4+CDDWq
zzxE4vlIg4CZWhjOzWP26R8KRj2wuruCkpmbpkVF9ATouK7G1UxSi3FNWNEo7zVk
BYwMOqKOPjWqQLjW4ORnH0rkxEYz1CW6PdsEJFHFxkjihs6SA4X4OW3D8KyW6HSa
QLmLOtPJwz6AxFrsR3mAxiJI6Nx6vD5UgqJC7Ltkx8/YLtrJuWkO/OtgRoKXPThT
fVgd4oWiIkQXRx1VQCzrSDVSzcURZD2HM1Gis9lDOfUzBrLO6vVcDNe3w3pVFRDH
9XBbjAMsClG4eJdppFnGi44KxG2ivx3/pEuhsQRGk2g/bw+zD5EwuTQ8I1l1PYs+
/Z7/jquHiNm/DOpWptTnW54BzUX3u/tVMeQFUQIRQQ+7w6f7gYLBjQVcyzIuozWo
qdOtUvnZOCmUUZUAOwMxwK52RESloQDuhhsGQI/BwxZBEOt/GazX5nzT391rrJFN
KZ9aNn8BNOwIffjwOTaog8rDFMWEh5bwmc26HaHKm759iOeHl6yLNSTh/Iu3tD5o
WeqTFRl2eSl6P2mm192iwFi1Ac825/k3fMv97eQk5rXMUFmcKjkumxeaimotLIM2
6O84fs51XkO5w2KoP4+6MEsqP5850jaTOzcOgVj3R0ucTGNMCWFBS6DjyU8BjWKu
l4oHnPGiDhI3vp1ZxJkJTGwsfYa8UKBKlGNKb3qSBiP6LTllwkJY1Sd+rmFm0gee
1Tt+VEr/VGyWkBIDBauA9JgDznkjjl9h+mlbEiNvBDYB9pGxstDrEOR0yRiwkFlW
ntmTMb7fv+N3jFOeio9lsESk76ad2m9oj5ytg3gaLvUutkeZf1VP6BRWWksBohL3
8ADjBztr3jQu2uOnQB+EdWEWwGtdh8q/Cvw+QVBwG7MuNtEI1oJqFV10GEdUR6ik
CfVRCO2WT8J7SSiYW8aadEX1HPt0XuqHQYZk5tdOT5inONrR83HBgMCLJ8kcRPTy
sMDFQqxptINBen8VE/dcrgtVC0yhJWG5CyAei0JhCwgu8bJ71dmA4i31kJ2cua2A
UdlnTMNBJMqel0XEQwanZUo5qekNbI7fy8kWZ0JCNjLzcNmb/AFkdHLstbS0hc72
ONexZou+cBddAi5ixmxS1xtasmyCyPm0y41VAKar9GgjEnwtc4S/jWkjSqGbeobh
Eqko7L9cDXS9LxxfNYPmIzKvEKBcWFVaSfsD+Ed2zYf7jCHkDokbGznalsS3piVP
YW7plhcVsiipjBu8xC2A+bEh7tMOu2fLHOrBLrIwtT0r7m7HiTLEy3axj13o4kO3
h8G7mbi+WURTiWP2b3KYJLSha3Q0dWfXJVncc8hgZUd/3tX9nd396+vosk/ZOecP
4x0+hD3D4gipkWIfBQs2de6mvybCU1P+Tc4UEh29GiX8YZzvD1IxUpZWCbiW+nnC
nuDMCaQUf3TSxpVmORhIYn+g22k7Jmifmp+CCQxSnFoEnnexXUqh1aclg4Rn55Ph
nj86GV9tOlGCZIioGlMEWgtg7Ja1L3v9aIj7zYjtiF1pSy6WT4YH1Eh2Owl5M+CY
dtZObSgS9P3hxkRT3a/+oubln3GeseTfrmNjZJ9bSK1PV3p/dvyQ/R/8QFQcq7/D
rQoMXmeYV5Xt2t+PavzCmVTO0DN3hm07vhiO+p6jGbTLL1FPGz9TampiAQd7SRAh
omA0so/xuXJHM5XbzwV+KbdmMEKHMjwDT27nO0HTpNg+iVtT+RH8DQxfp6fWtXId
jmuRFvOX23XUSiCxhqM5z6DpacKI2t41NJjAb6cAdU/1rvgGz41fioNo7i//nCbS
0d9FPtEvalux9l8tRA0iFQzz6qQGsFeq8P76yQd6xgzx6CCgCEOs7Pbwdg0ReOCW
gi4229rXe8TRd1meNJr4S5nnM65u8YVI3R+UC1IoCJPVLjQCg0HU3LO9/v/nXlFv
NK/CxtiT8pxRuoxgYZ8wfFvW3tJ/ztwLcO2MpxlbvfpK+6C6PzzQj6JBX7/M8bLC
JFmi+/BSmRztU7bclNHkZavo4pMPuNBwZfS96WHjBUheA7v5mEe4fmFhsSwG4rU5
oaitNVBVenG1vdkmDMRDTaG8FSmDbjTewOxvpzqi+ulDfxauGtW8xKfl0dBc/nUD
ga3Cqb3+0m/L/Cl+mJ27hKLvW6rsJRHHjo2qpS5QacrWLY8eers8jdSy2tBBfi/W
NoTvwgf2xkrTNchEvtsC9zFeDnfU6JohHmTF/8O4syu/3Qx+TwBuiLsTp/TEtsRx
1IamKeoVbu6pClRZln4K2YFujXs58k4iC+XQMOEHEigu4W6eePQufaHxnyoXvcop
8Ez/+MHSFZyAT2xWw1HBT9vF/63C2Yhvp60Yf0pZzec/TvZkKsXSQlb5T0u8IjhL
jJIvIhVzOaPoScnOQlMUu/1nfxXedF3wsceySrhYodvTtWVw3Iac6knVS9JuQjeR
SQCUGI+rYNAcVpVOCJr9TmUuSvpMcBrE9wMRt2xKmlKoWmZ+rhe6U84I13GV2A/z
GqdUflvybmK7RnQBEH1E3oqWe9LB4+OUqvd4HQJa+IXf9ozzVaLciolgj/AB/5rS
pcjUd0RgMe8p5EBlF8pAcUGmXWM6J5RHLvkKJgGKzy94dXxTrIW6l6Li4le6TMwy
28jyUQR2t3SHNz7Apz7nAFMNw1cvegSRnSfWCsD3311YID0W/Jvup+VVIU11s9QE
ztofz92eyF851u/7sU0DcEUG2YTGBL3W3+/PX79cdN0ykH8VhFh+TSg7qio5NXTj
uNDPxJNplPjRqLRPi8JskU6poSIiF3DyQ0+xI7g89foDnickUrJ+y2R9sy6w7RyM
R9lFzf2mQXUTkG37iDCA0G54/w3q/jkEE1G4gz7O6/ZtJ5oC/jX3nq2TWabHCb41
v6Ed+QQ3EXVQw+n4v2TUK4dL8BimuW5xLSB5lHFihRhGzEYfcJONlntMaEBudjb8
i6umcxU/ScMGT/RrMLGxdg1it9nr0sp1q98PwYYkOl0oeJ3Kj+c81uGgl5a7YeOU
fnKBeLTrW4POShn9W8ryBYWwc/o4uLasbhm3OOvlDHuEgCRJSfvzeqt50x1SMZ3p
KGQZdZOVrkd919u8OAxvl/2WZTFJ9uo2QV4Yum2zSRLCWEOMm2BSQObHHdtaMVI/
K1ZCXT5GZh9G2de9zt8NQnCj15QdAl41x0rvYvDMXL8OO2Q1oZWcmAG4fWHi0sl3
aNXiO0PrUZb2xBon3KDGJ1OBTeb8QnhdbYpmN/rsKCkyWcKdZgIItCJ0dZTYb+ZJ
toWEGVAesgOGDJuY25bFAR4kVjLjCr20STCZVROhecPHUVwSijrh5fJvwYEzUdIf
IJO9aC0nydc43po2jMQnTCfshys+1sZ6qZHlMxGgkpO1gEZaiofWvqQv31B6IxCW
BLlpzpbot0fZyWQQBDieTDGCdQKSJe7oK4N+BjuAAZ9g8aFQmxij71rDuSPtvBwW
XEL3uaq3lY5L8gAr0y6726js3peR/ZFyni6ZOWAWuX+Y2V1LuhFiVoscOIFDIN/c
XC/KZj7CYkmzBM98V4ZuWsT9ZA51f4mqAo62pBikEujZ5SZwxs1fe0p7Re4fgZ4t
iogzUTg+S2hlLRw1mjB17B6ixYROKpyLT0u9G4/jMsKU985yx8YsTVFTAwCAfJrd
h15r8jmxbR1uWNgBbk29N2fnaZXliENDwC7rHchi31QBmO/77yz2RMK5QMu3aqxa
0420oDVZ/tF7EWHorToLZ7Y3PRfLYr6FTHsjzk1ANn0xzWZq0zLPqJBIbv2SW/uC
dOraJOdmGpTOoXSIaj6xXVElXwQDYm22BvfrBHgmun4QMliB/oRXq+0I3eysgf6V
HJJbcJhoEWyivWx5TuX7q7WnS5nLrZixWey+HGT8QgPYSeLGO1wD2zykWifePH1B
0c21fs1X0GnsFZ63B+E0KWCXiOTl4AilZgHoBEXqEVH8UBevdIBO08lKMbzikQxB
DurSHwOIIzJ2J6K3MfzTOAhb1xQ8P6OVB/BrUt3ohQGTRwObCtI9948qkqxNf8mz
JDuA9Pt7HUhbRp2v1LxetrZYgdsI56nc0fZm7eb2fGNvsCKGmTPNo8sYVHo7o5ei
/uC4g+LSA5zAdzAnF1JC3GR2BdKmlEFIwYbokRDLtvJDBfEFlnN6pmYIL0gkJv5P
Nv5O+rVjg9IzGOh6OTVbf7GLaYmTob8wSD7UTvQGIYFO9Ru2ZOFt2DPhRJ8bSCvC
xBiOSRuLXV8vLWc36t6r8vkim4HKncgcOJ6EmQNu0ayodsIXj8PRIpoaxH8a8HJK
WZQs1osE1e64tgDUpYUwO5hqiX3R5PZTB9nIrX1vqOto2DFAVUkXJ0E+jjSCiwqN
36Lhb2c8ioYBWzFb6NT4jzJToT5JIjtECkx3B4l8I2Oepd9d/7ZkBBwDiSiguw57
g2K+JwmqyfBPWFbaR/fUTuQ9XXTAmI3vmCFxsfWSkF3cC8dW0QhhvJ/iiZO25Uwo
pnthBVveObPFUsqRIDd3fJu8gwJc6xksBmUXdyk/P9wO/Sp+BJJ23B86uiGPrI4J
1S59Ac2xOtv5jD+kooUxitjpz53/mhAkVcau0Dr0npJ4VVVeT1ioe6S19hJzPj4I
IAESVVYsmAmgJyV0y64JssUFZkWJ/U/NGy9w9K7k9tGPEc0dQgDYDJJ3y3uMS5ty
VfltAFTywA4Rj63w7YC9RH5zZGCL6WlXxXgwfPqU3WEyV8QNRT/81353WHc6kfxR
ML5VsxiRwYXS9qHhdNOzTi67GWG4NKl/TZLHt3h6SfjxWtZ73QRdB/bKatuNQBYw
0M+sUDGNzTMYyRgUj9T/rCwLVnKKVrHbmIfvrfwvrY0BxqxcNuCY1YOx8SPi8/jY
BMEjCZ9KTJ2Esel0OMBXnvirJNOS990t7PPcS8B5SGWfqAP3nxyzk38iaIZQ9mnB
uF4tyFi9nF1jTKE57f1sq7lElY6HNyUW8O9N076vOmceCWBo5vCawMTiVlZl7yhY
x8dMf5Gb10a2jgDURvI0+uCFIwc7q+1MEqA48FsqX7pNcron87HD99eiEianidwM
RhD/ietuE31dVlnrePdSe5cW0bffM3OMFe7L1FbNB9GKrBCDYmtvmFlHYhO2cRGw
cYTGmHRg7PkY3TMIZTi+kdzl7uJ4B/i7em3UpgFaKNlCAL6hpfmII/tSyp59au32
VskagvwZmik1vYIrA1MX7D5yAnQzVbhB3RdzUPtdLT4fosZ0KrNORWqhlvlbzTvB
+4YNHhc87AMBLp1y6t19jStkT9gwsZlv0FgO1j6MdKNX/0jwJ3+pgVIrWB6RCckh
IE7FDHK4qB9RLjJurvOpXw5z5L78HjppVYZWm0wN8GJRXG5n0otZ8a3PkFF2v7Gd
wpzZtPcf2qzqxKOOWHv0lsDtx16aND0/5ll20t2Ji37gtCI9+2B1epNpMXiFQSYH
OdHC8aAgJtY/B/DzAFM+K39XCcZzD8WRuSqQ2sPZz5QXjYGjKRm16IHvRLvq9VHw
qn+W2lEO9P8DkvKDOsiA68wcdsp3BkCUXAH+nUqq1PdzuRNSfhN4fk7Kx7D5vP6v
D8DeFf4JmJh5OAyqzyPvRtuPqxnHJAIu3HSGpXJkTfMxvHTd4dPH3LeW6NzGfVN+
veteOtsz6xYgxrtDpC0WSx1QuPfkLJ9JdjFr3K46xEOcG5ImNI/sjiMgNYvwe5Xc
e2RLWwIoTY6nAOjVilWqXFZJFm9jq9Rix5lhpvuK1I9qjRGChXCpw2W12GN5vE2a
gR2TflngMtss5jLBYcqzkEMCWF95DEB2xIFXPel8TiAdhZ0GfrP/XeD5PEK53t8O
lXW3cEf9M54h3XvtA5XYiqb7HEIS4T9zSt8g7WwNqFO5bS2DoDEzv1huum4ieDNI
QP+WGCVFU5Q7wZ5X3UjPkaXtmnJDfg3uoZMr5lFBljfwLezgKxATcBLZMjDf0X8+
5gb5V4oHMeHQpz4rQT54oW1VlAO2XUZ4/+pZI6Ez2uamaSdl0Q5Me6JOLSh3YqcM
blLIE/9mRB7/HZCBN6FIR+K3jqduV1GasSR/RGRhlCiaazXwLsXpKykr4kxfktSh
BncqcmYkhcnrXYfKpvqfcMvQ2K9/v9rbG4ztXapPnoC7kPKufCC32z1mJ/CWF3VY
txlULrudPKWvzGXAVoB0M+ztJP2Mik4VV95KU7aE6aEqRBe35nwev91vPcOQDDgG
0Ibyf5ykoa6qw02g30TuvmJjHrocS6U6198jxsK3O6MF/jDNxi/ZCV/owNqo6r3e
NW4uI2WqC7tOd6Y334gSvVSQhXncCeguOVSKU4/4E+3PEa56czZ8JxSPYqqQS+S9
39G7yRouTdhLFEAIkChlOIi+I8tFPPkBmGqdLmENXPZC/5x1k7mOTaSrT1qLuZJB
GjCzwEIaFiVx3K963lELp2qBTdnuSen1wldz4aWRb8zfd1Mp7AjJf9yhOiV8p9ab
tAqA0zYur/2oCFMuemi3f2Q7FJwny0r6PfAEWqeFzUZ3C5Kf7wqO34BSOlkvvgDT
fQnpjMkhkxH1c339anae/i7+emng3aELY0g+Xtoy0b+AOZY9mO1W2h32llTUEDXV
EaZb2pOom5KghNiZiJi+EUIyOYK+BhsnO4Yi9k62EGSjp3LhKpzg8Q/kCxBBta9H
EXHO6+rKEg+3PsHmr8jHzACCS4vxVL0nCfw8rxvwrLzIRpdYuEFCl76LOHMGDjSt
noA2IlCxlvuDw9ZE8xRWbFFOR2SXL6BYwzZNSUhkH/14w5G+9yhkstjKTZurLim0
DSVvBLR8cR6rMf657LTB+oaPp2MmjME27l9liz9ZjChk8LoQ7AeIU7PQoCjQir7A
te6Pel8nNhs2hUYaxMkX9DfJ1m4Z4Nu8+CXV3A/HuLpY0bs9TGuqaJrDvexYn6t+
h9odeqodJE7CgtThyJno6F5AYKnYILuagSYLZhVB+jAM9MkckxhSXs6FVL6xghxt
ydm1YfvacnoULeXYB3xyNvGZAaqdoc+lOTqWIXaCprvoP0Ol5YC/pAX7Tf3lcnuc
xad4afUj3KixgE3wl0SKT8n2Q8MvlFQidNxiPLaOR0+/N2aFoV3fHNWYoGtKcO4g
28R50kBS//OD9vVLkFdiKcB1beIC5Ck6lXcUv3DRzQuJQukPHcELA4pdeMMnZMRM
aOf2a7E41n9t64tTyn5f7BlpvMelsnhe/SuFcijDdCRrRy/C38jRPWswUmp/1WPe
KvewqCTxZCk149SkOCqwD58KDpBkcPQS5m9E7Y7782Y7LdFMldJUZvPly0uwfQyl
dX3MlvBv8vVqB3A58C49TCkBtKWa/noAccjYvMOibSosbPAFi97HZHi4xjvLOiWd
1T4V4g/bmsFmgeTq6V/ErfG5chhb/zgbDhpS6Ls0LbPmfuAEaIF0rEswVkuzIeLz
+5Kv2uqkiJVt7N1dgjIgwzK+05xPAjd0eVYM0ZcLAP1xmRNY3QdsGXJlaCSR/8xm
LczKvu8GrY6vi8tHHN6LUzYq8zrQQwOjQa4V7/bP4r3G3ZvS/kj1nMKu5+c+rjT9
yFDVDFCbTGKzkcc9xVeJB5VSyJrI5Uwis2DX3aKNsehTTd5lzwyMz2ySodTvl/ti
xQ2tKNcbtz3GdWLdipJ18kqCKiGSCMrSiNyBq7Pummuf9BZcXtzIcc0tFe/0metz
FPqnJMX6YVOwnvSiR1mgkWhfdTpzaYr3RchEH1IQhsKpKSwWTjz9hLIRWaBPQZLM
6cnQAyTW3MXAalmAJ1EUQhQwtwLMuU6h9IHbLpEw4v25eKU02w8ns9snmtDN3A7I
M1BuXaFhbSudii3tcFCje+HEiDyuZAtIWlJXBC29kmisQpOvYgHZC4Lj35D5tBqR
G6JX3uFVcJKJbjSZwZdGiZPVgsyaTSxW5fEYXZZdYdyEB2qVZBy9U50SNFBMVo0F
re+SqRFpzY2ZIy/OKpfpjJKdeGFK1oTtZtbtYwzpIP+h+Rz+AOHzsOfdqygjO0Af
R2df03QUyELeSj/DKcorgRS9/OiGM5d62IRL3wBLAvkeoATVsylcrF9zWE1jteqw
Ni6ebvcoHRNH30fcVPW+BSLEo/tOy5v1ZikHkTFlfLuHV9z52CQG9ir16T2J/NKI
CYt4TS2GDAVztdmxiKAPRq+5Op3bCpHREaxscqOJVslNeTnVrApR7ViL1jj5kuKR
/7hYDUSsaV7TEJ0R2sDUCxbjpL2rVMk9/v9rjXq/hSFdvgXMG7HtsXX06g78/5yo
weilpZnv/iHLdtZWlSQj0GOOeLjZkoYjl4+wDjPeL/oJERLAt+93f5QciFvZQhUc
185+X19McM6u23fHDtU7soidswofonU1de4gnpWprkM+avxL9rv2H6omAu12+9JN
0EDl/9vskCJWgOyGXwjD5Oovl3N68Q7ATGiDZoJBqWmYpeXepdqkpJbYuzzZtlOj
KevKpn3QwSHOfBHinfDIAZJuHF7SmcL27GIK1docSCx4fJdL//ZSehfORdezqfBP
pSZ2jvwKPeJr1rXvZtMrufrB0YYTcykvHaUEb9qt9XpaPv+8SKlmttKwfsZIAPmH
nMYfhzni0oQOOJ+w+cNMAPClI+VGmTsxVfry8wSOxKMwXP51exWf/o32acs4hIgB
gkYybICh410Z9c51SLbsaPNWXRBSn/KG8GZJefq227k65fyuINDDfp86WrQX6y8Q
gEQFbkzSAFzbqgfn+zRXDeUzpF4QgYHlAp3tCyaoxw57HYGwaDxN9ybyIJx6UFZ9
8PXWOBP5p4nF2DpcvvrkuUC3nb7NpiGf3K7zm1eml+KKSCuWuOqH0gjyaWNgUH8A
HMJzO3fwW3eH2+lXa/JG/0vdgYRLRaFUsBoLZPAgloByOVg0GLntaCCC+HcY179d
bvgOiFc2krlgOtoyZ5EIdwcWTzGQgRqTcUBNtiWRb2rBU7l/6ORTfPHzIcBJcjyY
Q4QFB5fh5dZqySnixf8pUClnxUxDX0IFQSmCaQPKypyWW23XfpHbQLwR/trmWqbf
459kTAVMM8JdTiluHDaTSsWWlW1nvvGVQUBE4mM2Zl8qOuCWN6NgMj4Nxxm8ma7O
nPYTR/w1YYu6lgiSzLe1FJvMDNipX6+oLpXAAvehg/FHp3Re9KGh+WcUE3neon8+
Dk4TWDQaAvhjUY0xUtko+D2Q/a0mZTh4d3/UzUnfe9airA5ZFTv6lxtmbn8rIICn
ybZqeKTX+AI5j/2ZCI2U/C+dtNg5RULN1jx1xC7JiFx50n0/XMbKwKbf8WwIM4Mn
+OG+OJYmy04R1MBAdWx15jLRic4wX5qP8jBufoBxTrkSE20cb8Q7ChNJe1hLIijL
SFzNs+pZalrFh8scDOTwbXpOOEAexNSw5vm9OF/Taw7NzctG6v8p7IQ/E2UCJ5M+
qPBbrhLEEOBYFqKi+kavfq1i6ASmimB6dzUBuWax1YK0bmT6i+bgmQNTt85pgpN7
Ja3F3gmY2d6887TcO9sOU/d24ZVT8x3mnAJvV+Uqk+MFJt6y0l9hozA+gAQqc4z3
1dtjoqBZ6dG9pcFD78yTC/kLbQ0SScAwOQRo4nuFrWGpRSBd1dka3d/p8nMgJLnZ
F+K81kdCtnuSIPNF0yINugap57Su8qb+s1L8HiV9VdkG28FZp+JYlmm+PfjTHiSO
5K3+8D2FP0xoNq1FHgSCd9qv61f1Lv/JcSjiBWgsYY9Wp/fJf+t5vXSST/SnKOD/
fuJ1tKoTLjNXUBBp4PQOI8u5AvZI4p66w0VfbiUafXIeLO5yayp+Udb895lStx6I
zIs5sgupdPL+QkwYX6eoN2X3IAg+vMw3Lkf1UWyeXxG2qJjSPUDk/fK+jZC65ZZe
5dWjCwpyk2HGBmC+dGmwcqHaDMGp3gxwXtmNZoEL7+0bmtkUCRH9Xz5bH+AaH+kj
e0703gVg411Oyn3qDSmpt7sTSuj6FPCcECNx1mCUcfzyNuuNKwoSkQBRdB0l1AIN
e8XDO7lNA+W01AQVVbRrx8xcO7ctvbIeOqSwBPik8+e/LfRxBBhe2k+F2XC6swBs
6MU8qRqJvd6gTaWVUSKQ04mOCgWUqeR/ERvPuymeFzWM0NT89FJOYip2IvuugkjK
3Z7vBsNP+6JpdpDcSMF/++Cj9OkK+AkrND5e3UQ00EZiNO8XYALHGvty1ZBFCACt
A53h1ahtT3UFh8Z/emYi1asObCCn4fJmXcSlZzL9bAbBs0bWM4ISdYDE+5iQPrOy
QHC60Bk9Hyfl1d5LYMJ2ep4FsYrpCRx8qf4hOU+e8Fc3oe1xblG5NbtuUM+PfppF
2cQg8dSeaI2FGsA5M7UJNbUv24mIMpBPp3PzV6AhuWaF0NyiRsdFxf9YVQyi9TBE
eCA5LE8p+RCKjj2zChy6JD4lHmP+qhO4VzYvE3qNLkWHYZL9zQiPbs3daAf4KFZe
C8vOIcg2dVGefq9pJuIKp1FVPWutlcAutwSI1SmQl1pg4esR7ma6bEDA7TW+m+ed
y3ePB0JbAbfo8QAB23hLaSCk+3TEACLY0y9BBqxnwTQpAGgIdj8DdN9KJouFugi8
8CLzEpDIXGm8iF/lLoKC7VaY8X0LSvsVlXryZ1bq6RYJ18N3pfAlGMWjAsET6yxr
Tqf6emPlbf5d8W4bVGr+2VXxNu5tFe/nKX3UvExKwPVESUPScLKIB1DFaBwVfubT
k0n8b7it7IsuaFmIwrmD8KdMakOlCueXIbv34jebk4aFD/btFiBsTIFznboZ4w4w
tdwYo/W2c8bVztzp4Ypm1s86rrZB6FcJQku3nM9EQwyZU9boqnY0Cxm8BLa9ByNE
sNlGbvEopa5xN64H11M/QeFSjTYcTKZZiIanLTBC6xdAfdU02Qk0sWKLGCOQPoa1
4W8sXnSqStlyfqhnhWNQZ90gz3PfdNSJQc8Ur+GhWWIhVzE4JGwhCFu4CWKHCk9w
2joKThkuLbIL7UnJ0gllOpnwz/IHzMkyIU+xgSYnrVKseg/Q/Y3W4honZpzt8rh6
/DUB3x3ODSuZCWzKM7TX1ZwK9gY72ExaaJsZQIiPqrCms4ScuZdfrJz/F1zQRxNJ
MxJyRCaHxz7hPo3UwybfOtjVhmEV4yRZGWdHr9IUvBH88B7rrBIHduJUxStklY+A
0WvyeJdQjcQF7mIsVIBjYkTrzYBBTSyRGe8k/n11kTO7tweWPVptXqEzIrFC0fMG
F66Y93bxs7Pg9Wc2+YizcXTuo6QSVdhWSlE4ttPedIZNFW09YSMseXe5sl2ilBmN
6J8ZzE0ZLCTZ9+fUMJrOVUXL3bXe0qi3yPQ4kFzga6TwliUaLJqqIs/XG8j2WlE6
GozgxvUSpTbyNe4wGGiDt9CdEoGZW7fE6CKAeQ+lIhngMOBrFI5wHpzrDrrBOHto
vQgy1LodedyOPIYMBncb2qLGNozQlCg3GgsbThVeOI9lfYMxWlIzXcFHqkE9Gmxp
PRZ9SJdgIEi+q1abLiSrLUfPp3J68Zj4+WZ45oz+MXFbPfs9QdVfWThDeWnU+8tN
VfmUl6A0ZWyacNfelKGI3v3nifbX1sg2qZedqQx58RDtxvUlcwhQCnJCAERApRAg
jyGVPctC38s9yYJwlFlm6l6G+ONHgQK80V0Nr0fEojM+hOLFN/pbs4zSzibhlCQi
9rEgsXkhmlkfA/+Jeuu2hXdFNkHib7RcljyI09T/7nzENA8VXF/Q77nLzcgUonPu
ourLVfwU8Sv0KPuoYJa26kgEj3XJfxzmZ8Un7uE6YYPxMu0SImnGgAPVXKhj+YL2
S4//+x8EQ+woC1vM8Erur6oa5neY8cZ63D4NfL2mBIRK2J/pkB/WDovbzo8Z79rb
5aSLN9dErjaK9F+O2BO+GaahkYEhHNz1n2f3UxRx5meW7xWl/tx23kFBOl82G6hx
XwRFW01IiZST8HQ+uzi1UjiydYZUTiFcH+mwOQ9lYqmTpSuvTN8liZ9Oq0iODekA
naxsCcrk1MhssMsJlR9V5lTEss4lxN0Qq2O/nens14W/4iAHPIuUypPFEhQ7el1o
qQf7cnVHMuiiVmgDCBAfplb/OLxgDmlnu5D3c8nKbaZ2pq6UQhbUiQeCAligsgDg
ORLw2dXaZjJGOHTXDWRNdxUzelKGZ9XQerdmJbogORK9XOL9FfoaKXd+mUAuX1Qq
zkyljK7nZtNWBm/NCCl/BM/nHytbrKGaayRvd3o8d7dFafeQrz3/PgDh1m7/jhON
S7zftMJpagaD/ePW4uIqSQfRBFJP6ac2RBGlehpT3sGbwGpLktvIzHYTK0o7VIIk
6BNJ9/hWO9GjtHh0qlNTcWY4olrOU5J3KwaA2uqJQYImnbVdwABjFBR3kAG8U0N1
uaMBRrFwQaA/4sZ9jvtdnrAo0CZZ5mPPgGJhMx/RCgAEci+yf6v6U7Ve2F3oYk4M
ZUiaIuACBuP5qk1y7VOpUuC2AE62eA1XHKRDPzCpv6wj+7djBgqxNPL9wFe26LFA
TS8CcxXlFRz3U7Be0cM5wm+0ZFG5EMjRx0TRskZ772xT0L0GXvWERh8alqoONiq1
p3ko5poXcKufvFrzGaf2EiI/sKvhqvNLEsdY1cnrh85eZEKwpZfPHcsQ25z1zw6n
cYIg3VkY7T0y2liQG15y4EhIk5gODtsjL3Qm88xlakxMkw8WAIjF1OGsrTmemmVo
o8tiEMVoFhnbzpfQW8OIbCfu4w4l1c3bm9byGWR/VmjaLB3ax2SZgxgSBdwP84ai
7NzHi4JEwXqir7BI6njx0jNd4rzEr3vDhBYKVerxIwNuqqbtvL7V7JTKU/OwruKO
8ifn5cZo3WMb6mSajIE7lt/RNbSOMatKihmaFzFviY7jz9jF+ZWzLOdi66uCdrA7
vIAh2mRTTgMAFl78By3CZ7uzvapKPUZ3lzqp0ATxm1pSmFrXwLLGCl+5EmNwC60K
ZX5BUx2tgu5rcEfQMCh/dn/yWFi00xGjgmRxo2hKN5dzMVO7I3v5B09l7uEykn3X
o7F2vSPH70D0eUI46mE10NIclhYQ/ZSxe37tpuuEVIIya0xVEQzMWqFrXoKLVt0P
iWIxii4w/mRUHo2idpW6HEDNzux2bkWX0P0bmTJqHVvRfoEMfHLYvEou/kI4VjqT
/tcC4wntBk5WM9ynlmFHyby+1oHy2norb7yyWyUB8Q1mOItQjfBp1vYmXldpfcJ4
Fu9uObUXEeTGsvljZRL+cMSw7N4m2YZoPfuKpaowy11DYTGL4G47dD2WeN0+firT
rrlOzfwDUKOWFGOWto4sK4vPyls3nAU+rgl30mP9qiTATfkUT8CiEOyJZ3f2uTYp
NNtLjab7HiLsqKft0Nd1zGt4wSBH/Yalv8zANpvIK7gS9ZOhOW3QXCb36AjM9ra/
Tm6TZHIfnt+zjbjWZIXp12Z+JfgRV+8wxojCCEm/5glLNiFfu8dNHUKw0KaU7u9q
8mJ1Zf/W2LT0xy2sKQ35OxAy7/cHv/OOUfToXkodqQlXDl/RwoXKWXE/2KlNQfxD
47B3T0QV0lErrKJh3Hljbgb7kaLZTEfrAZsHYSr9UjNL5YBPMHUlLbU9/5YgO09k
8Jr5YsZLVsxT5ycUOGUrg1Bj7z/kWJVnh2NAAJ6dvwtkwCLTqRBFRyeJoH5pLQOR
/UTjiHh/Z7X8X62u7nSPXGYqRLiKub4Y4Gc58b/qQPBZZEFB/TDhTPDx+vK9YeW+
jDuQhnA5wchP58LLli0b4Qk9Wft1Cj77m3aGc4dY5FxLcGAdhojOCdM1L5tKk0VQ
6xKr8KS4PvuCm8oYi+2/MEazD7NDrCOvzEf0uhTWqal2XXln4wa9kvIBO5qs+mTh
E0oa1DjuTOughGuhCj0gTCX1eGT4lwuRUsOQKG9p0wiz5KXz1EHC9v5s/+I9ebo8
rwn5axvV/CBoiUdht8/J2PfJhwXqSyiVJpesL2WtmRsKu8XGmmrX6tHoT9/H8NI0
lrW8Rsm/mpA/zwGMVDWmmVJuet3wQxjNrZ1CdrFV4wArBxSA2zpJpWGZDfvaEGqJ
clCeDDXceWgn03ULoA0R988tX/hJpUllScewvNtjExinz7/l49ePzqFzk6h3fRzi
65Za+Ru7UgQtrbdKM1ba5eRnc1OJibvLRzYAqpJLq/er3HbLBbPtzubrYm/EDwA5
14h8cLENLGr1AUOcH2jg7u0ovbR5RSDGHg2doUIz15RNWXKrKjOlI4Y6ZqHiYGET
hsDfm7SzZA4KUR0tINu6ihVVzC0MYE1YUpTuJa5JXD0NdSSF28LbVhY2z/Hcir6u
CKyUmK+rH1ofCHRVUvlFBTRATz5DyPj08yBsyulNgqRJH2aYqKjFwHCisflTTEYr
JotVoLdUaD4/Kq7EOGqi49cqUclVImN1VwANdaQbIVqjQm8HYRHf9akrCPvHapPZ
yvts6WD+asd0TQxvUdAYrQX/GDfO6QFMzKX2UX+WPC4QFC8U3Tl6O2sV0Rl4MD6D
Bor78zXdYYV4Gk98ABzrCOxgy5AMobpMf8EY1pFtE8AI1bPw9W289htXRx7T9MrX
STUzqPLmFo4ylSo5EOzGSZ+BQbZU38m4yfVUKtShrGFW+1Q46WILIeByPX4BKN+r
DOZIDFUMBPXYtNfEcUwHqdqz98mpwqx1WuB0wZa3VVKW6Pu6Tj2BrQrImqMbyFIP
0cMPG2sKaZAyDn514929UuY/NC8ccbSPUhoTgLWpo+xqdsP5WV8FbQIvagUeY2QE
5VDmIno4eDpHIutCWmLmcO4EG7v6swDZVlT/rKo7uQGX04qNoRPLeQYgkrN1+i8K
lS+Tb6DhBuTO/M2IfKXd/d0+GNDqVxHMba2nH/iKdpJSF4S+mOxlbzQx2Nt97Xg8
tdyWof+xmhU4AwnjSzGoe/nZynX/gZ6c9YGLAaquMryZ3ZsbC89l9k+BllJJJC5m
im3+Jh7p0g1C7nW0a1AGYwfX5maN9DFGBXjxHBXTWn4f2pOo8xHbBRnsXofZHlIE
PmOCdcHxeazTP8LrUO55QgQYlcEGxWFRTLy2noT6QM6iu19esGM2SCqzwDjQqMsV
dmrLAYsOkhwjHsoh11SRri88wv/98jhUJqiXm1xjmF5P/3Jp1t8xD5sqdgi41jCJ
xIe5Mdpy/PewrvOKPIJ3gkVHy0KI5JwQ4SFhVyO6uUPB89K/PawKWqhRKi3SX+i8
fqgQw0mMO+OmRV9rmjvMOHlcqLRnkVJfCGIKDDnX58axNM6FyzL8oGiwcS/hRUmx
wgASgPjRG0Xee1juzOgzVJPNENjDZxT+6x/fT+fCdIbFk3J+26mCXIP6sUytRIAz
CI/dInXiw2VXPMXhAjQ47Hlv4WFIo4iGVcIrB1kbLJ3dZ5Q8al1U3IzRfZ/SRVf3
QFkx/rv55hoyhj8pRZ3mqecBMET2I+SFf6lMejkKzeaDA6GTSJ50upxp5tgyq4Pv
1BiHOViT0RO+CpbLNULhxDIAWXa5hSz4KhkBGDLSDSnNg/4gnfhLR4XTIPfn/t2H
6YHfFVRPgFEkXi557n+r2oqMNFgpMlyEfHaAJVl7cpH/qJLvscTB8iLiDSsvdq3P
FMcmtKuE+p5lnX5KvBhTGmx/YYpOvvVs62E3nJ2jl4ho9Mvk6jCUkij0zlIPQIUi
mM7FVJkIJiiBMvnY08wsTwZ0WDqeGWNXbFetSHx/k7TCGAWof3I79pk5VAtinj4y
z7+9q0F78WEj6lZdgBj28VsRnAF4uqp01edYh+zix3jHewZp5J7VkgOdH5tJQPIJ
zNdp+8uao/01sRnBE6bJjdhU2pkbLRuapmpdVHpol+uOklY83sk3L9n1dIdjQ3BE
w1bl3WRdzK02rliMZ6dS9EY92wjGo5EM5cehLVNi4iEKl49W8awBkAZKbgW5XKUg
TpDnT36hCj1hS10iF3x5CUsRQUfEdxV62GBg+HVxT6K+38WScvHhbO1oHVwwkSIh
M6BjKjOfBZqpViX8r0QfT1Qd9a5vhWI4PAuyd7UyzShu2YkRaisp3ZMIqaYUnI8r
59CY4M/3AACrXMLAVdg+9SjH7lPhogS5J0daQcN4NSf9yphPs0Jg3GZP2nLq01tH
52ZN36G9EggwvkPo9MWtjpiRmKxetBxZpkp0uG/S1baum0He5JiQ6hmcrrlMslO9
6UKlVnMPS40ufqXt46Rk4uc9qpuvYCfwQxNJ4NjXP3SKD397wsSymF3XnMqRC3sN
5tupnAS3TK2O8RSHi1aNrUzYt2ze109X7Qda2v5/EJ/wGWSw2zeMqgSuW4W0BgO8
0uDTRAmoDxCcc7oS1n15jECAnFY6a0f0eKmfpKmVXKyD3nbke4cBT9KWofK6Z7AM
QfZLb4ZKeQCLa6kRTBbrbx6G1QZEckq2JXP4qyTmE1W+SVIoq8D4KKzRbvQTEXa4
HpnKMbzDMvrbk15cDM9oUip1GjxEy6cI3WHh2TfM7tyfp4/20af1kpOBFE9fQhys
EdOzTmB2rvfWbFnn3SNc1mC4lxa6SvHgTfaKHdmjSKoDB7+o2Tt+Z9H3ugqbLbG1
GwfHKIR79d7qPtOsYukWJn9BMzIojavHWrCq/2hA9fjd4OwHLKcg7KZf86hIdTb9
lUqJULuWcJsJoxZeekYO2fnLK0CUxwmFOk34iSLc/i3B/5Uc74P71e/C2mO53ZUT
pWVnpiKHMWp5yJp7npn8J1hhM6kOYMLBlzWYz1pVmz+WFchPBh7RFNuHfzGinFVE
TfmCqRVDS7dE6hz8Dth4MJrHEmdc+vImfa61bh8PoS1cgbd1FSJUohsOoY0yeGYS
y8UzTennclnHQRbYgujsMAJyqUh9V/7j+YF8ziYrbcj+6Nxan46PbCmvwzUFy6iZ
erid4pkrh2ypHlDLDfs6vLW5v7p7ubi+RkeR527hP4dfCo/Zwt8Db42ONHy8fL2m
sT8uTOMePrBLo/H+ZeZRHSnzErndNDMFdIG4CiHbGZNkSOv3MMCqha+xYHCgxEKP
n/63BQhXbBBb/Q2R4r9l9muB4xDP4Yh+KHreVaJclQdu0ZSpqWStgpMvcN0VkaJg
c0Bqv+FxKbE94rTaXGf9yB5tEF+ccVJ+h8Yxq2wXxxvN8Vj6qpM9jRtukubAk9Zi
0MSeACvDNZ9Eyz4zAYTafnD/6ceQYCQHQzCw+evRaP/7N0xC/m9yB9OU56PsHE5M
GaqdSYu9gQDd2EDgshdYFlO5ufstdfAgd5Qn+wh1efYfwL/Rdp0ccVSINhoEVk+k
dbFaTZR01tRTDC9sgdPNXx+NWvrhV9klf9x5oFyIajJCCNSx2PSb8WNzGYnGXcDH
846c2ms1XeCHBooZbJAX4au1akUy2vebz/PkqBC7VAULNaW8kyd1eD3qHMqsHiO8
t3w4rEQNSVqL4V+3jJiL0mSYAHqlCrUO9JBsqZ9iIOwAPwg0S4M9w7BIQz3W+k2q
5HZpNl8NnA8wpMqEyO7EhgkZhYmOjvTbh23hVL7q6MyUoRiViKyhh0JC6MbeM4Gb
69jxvunGo5V+ZWgNnN/YYmyRYW/XkvEloU3Sq4f36HQZqi/gBbwTAHXiIma7H55Z
rM43DgUqzPrlikY0mOZd8uIfbSn60NzCy4r8OeC0ocu+dghUSJT6FAzUKa7NY2oi
dJrf1iNvfZq9d4Q5fDN29zlX/cUj1t9n9ENtv7egRBT35EykBZvp32PEbLyQmsyy
XI4C7ZqT9mY80+b4A2bxvMTI188p3YpQIGtzVfzP/+obwWsG+Xegz4v+L8Rjw2th
lGwj0OZb6VHVl0p6DurX5vd1jFyOCoZdSuXIyr/ZRdu5UIROMRQSbp3DKMOoGN50
7U7T4hhqb8sx4u9pccgVIVGtyZM5jYXzb6szdEjOZSSO/2zTfPoVHRx+HdwbDpQ4
95+KIJlLoiZJ3oiFmzrnGBGuMkV8CJYPKt/cUraP0pI9WNqbxq09ANmuA0MEIz97
3PtlhKmFzLQJkH3GNyfR68EwMy6tBwtG/IyYyTyr+610X4PV1BV69l0AoyDnADyG
Egpvv0nKfS/Cx4QgO74Nr/zEep2nxyutSYDiuXDUOiQUrCz2Iv4fqxupkQZ5JLQP
fghnNTtm2PVTlVdBu1nwxcsDcDBriheZKi+iI6k88qODKFmPvxoNQqhEUGHi8nAm
LNgYOQehG9gaHBKptivnLEjs/bqL0ZPPmfNY1HBO63IaUKWAxVQJhgm5Q8RLCrPT
VkyTx8Jzcoogq7WZzFj/5MLg/zNGEOVkkEhqbQxb1Pzdk93Hb4AqbltWhORy3xnC
FjiV4ZMsTeQI/N9CTCztWDR4HdwC8qMl2CYQq67UoaPN4gfdwqpzK5qYqxLBy4uI
eXNSDSOyLG3y08U9n1tW83DGAkHU5kyI13llrGfKsaYipMKZ2IiRFNU8/VTSkoVt
rqxYnCwVlI5eUNfRQj0rDT3lB9kBjhOaKH8rEel3ou4+HEjNJN8THORsl0SHWuhT
hg2A8mHcKnxpW/JTuPfDMIPeR9HsMnojOCxQIRvgKvwL++gGcRJ7u/+qw01RLlfl
YYlWsFPR3iuWNd4ZisyRaoX+l1yb8rILMsUXJeZcD6JzzjMAXAH/0GdwdFQyUTnM
pFPgv7CfS3deXM7FlTgKLigSJi6YT4JheskuBzBSKBN9esGfgzI0crdVPSddyMSr
NvJihpwDDry3c02AHPVk/grJnNGAzG8+WHYfi/Q5ec5YY4KmdJnuwM73lcMNV0KI
NJdwm0QYYjom9XSo4d59d2/3CUI7qm+AKudco/7nD1T8JwimNIL20wcveJlvuKz2
yVo/sG97+vYycRAenwtNLDC4OmTU3/MpcbnIte2fJrvnlpmFkcyPC0ak7NdFeHR0
PcAYAjW/aoaYZll5J8v6+FMVZ8r6xw3GC5Z0FWtKEFuAMIooh692EUgzwMqN9mMi
lWhjpg4cR1+NuWuuOr3uaG0L0OHXxZLMr87X+aXcrvAWtX//eMVQGsa8+EjZKHCX
ZSsMJE27n4Fxy6btRHtyBLamxPfs4cwICCzScBzku50Equ+80/XeShYAcynnUJQ7
UACSlsntKYF+DCl79MuSDYnLKk8hgmmGggG46cFqm0TlmOiZSFkG3vKgINqBQJ+d
tC85s4hHk50dmUUDQpVZOQi60Ol4BK06vqvSIIUagSNOxNSQqn1DYyiRzE+ADrj2
1q+zeS0etWRj9ESRvmNMU0yV23BFNRzBk8Q53XnwZGH6WUb7TW5xOxzGsxyd7Ji1
ML0/ahrE8dJW1Q81UaljnRFq4bzyu4cf3u2F4SpDcSKri8o0ZcpBK5pMPIOmf9a8
MlV/x7gZ674pmSyDGg6AYT4QxYrFLFS4SwzGqVSvvTlhxevzE8eWymyigeQLaqvv
MiSP/w3nY0p0UTMEfBOBauJ2NJzqG2Y4CFHQ3J8QCu+K+wbrmFqnO4+CgUnrexzZ
/ZlqFAcQm7LeMqdDHudeszC8XWVkxJVfw2wNascbY30hAgZpdrH2/SyWqzYzablG
U8fckusWxMnLTPqLBFqr150pJFTIUd1HVO5RT0lie58ZdOS8B+lgnak/65/A1B27
NIqsgU6MsV1jz7bZhdoeve6liSab8T6NhXE+vHckSjtvo6Ir3rqHaosdvf2Q/1jI
+jqT+KkJK4CZThUn654/EHUguc+ayMazdjVzxdqdxKdoLvlY0DJy43T93qSmsXNV
C04ZzwIiOG+qtCvje88ZShZieKOpxW86lR/kR0ML7ndtRcqrUal+xusRdYMYt93o
plevJ1Pl39BC6xYmZ88e6g/mS4izncORCMWJyrbmpwoJDPX2zAUl/2zz1EiUhU0x
T/C1OJ/l4wTEJfsfXt3vvOnFBaP6qACNA4px7KJr2W/j8Z+UN85Gy+Bj4QsBZ37a
P9oZUvw/iM5BXBEYty41JMz5JI2W1wTsGMjtLWiENpCzfcrnIgQCSfp6lMQ7Xg6p
smBjoxEwDuXT7IYG6v9/e6n/SG2xD6oPaXkRRrGcPziPPwGo31bAuPmTDmQ5Lj27
Dc729OaxyHrYL2SN6H3WGPvN0qvQAfru7sKUAolfgWlqXicy6fZMJU7YBWnjyfUN
dAx8qgxEQMd74m4KRJw2vac/LT8Y4iIM2EskqGJmSnxfgPSPhnEjdAli8FZzMDTu
D/t04vKlsPWAGPJEHI6NupDGEtlChLnpqCUtFrHNjOn5jF7TRouHxTxzA18LzlOC
HSAFNx4mm3cmH88y0gYgZ58zr7F9pdq26I3dXE42XREScMEvhPVtb49/QbIRYsV9
ssObcK3u9RavxIccfmlu2+8eAOmg3rRyVyE5d0Cs8w9Xk8XJc4q+CruSoSzXpwl8
s0VYieV21bG+4He0Ii52v8TDxEfxYWne+Kzy/eCrL7VlayTX/xS5yFDMJN1h+mJt
WQYOU1wrHl7QIHqIyn0rFXM1OjVkOOHY3ZHtADRWzT5f5WEms2FrM5v6PhJ9/L4D
N0ZxQyzTdW9rFwXMReIxmEf9RyqQ5V5GU4CJ1M5xN9moMBGAzI12u2Dp0fboe60J
lvqrMZmfK190T2MCpxO0rt2Vyoq1im6ITNvFUChCeS6nQwadBilssWIi1mg+Eixm
YdcgbUbUUEeJMeXybB/KPck8IPlvaz1OG6KOn8GU88HKk58q8+jVH/i1bQk5vZSk
NNMY/7y2zk06zmmc+Sb9gaGma4kF6XExNY9HwUt8iSCgMsjSiageGrv/+3PbrXFy
N3awSDOw9PR1uz90iNT9/XxeYZucpAchkBFYnw+GGT+Xk4+wMm/MJZDOP4J9aiJY
irbwsNqHZz9v7pOnMA+1l6UJANoCDv+y/PHryzd+3MVA38Cl3UE9YINKJIB0Rgd8
RIpxSbmhFXLt48haVeEP2EmGA1lOp+morlSWdmL91bbJus70zNrizpnw9vI4JAp4
+bJ4l3Hl5+/7ihK1ELfnEd0wO0IOrfscuMrigURgE/COapEO84nSd7PN/7NjUhgf
Pizbr556xQSm/lyDnqkDZojZYkc06iRMcM/d2U9z+qGPbKRDjgniNcZ5lu1hBqN/
Q/cRFqVmKR7nKmDHZ7PZt/ospDF5jOyWcPDt/Wv5DYS2nn6gHMLmJu4tXPWpEAkj
qdDykha2BLz3U2xf8g4UqHNpJPgzVqikphmiFQrZRro+NnX4IRPEVn3IlzTjP54K
N/G9Tqv4QjKUuMbOF8Z+0dnjKffrYyBJC6pxAQJhipr32EaQyx4Vg9wyF0gqvZJ+
7wp9A4tBudXROyjVr3xYWZ0xCrkwnlkFBE28XNBptMVDZUpdXvT3slDQhRNs+d5I
6A5QvO/9rdMmW5kJXkW8YKwXwwKwSPmt3xWkcU2Y9V9Br0EpO6dk5Ot7RmxX9e7x
QhUuikfSJtKSx+NFV2PYOhZxzwfQa5Ev1mDX19xVI7/gnWO/mgDhb47SC0Pz3icy
PnSlwdLR6TCDeQLY6t2wblFb1jjgRJbttCS3XBJdlcxAAWDtCZpgA9pcLI9xH1jh
pwQMfB+jefcDeEt/YMboiP3gZ7frib/UZMMmBOTJMDa7GHLcO1hSpnVo75ByK3nh
uCyQ41FUPOiUv11pvg6kvhnoEa7oW6De3MpPLCT7kiOvLCZ4HyIVZaSX2bsxmK37
Y85Jgihmke31/d/3+EIuRoDH8eEgHVpEzz99j+1UAbqqtcZ1p/2Ra3hjGI49PXtM
wr9bI4HIzQJhSj0rnSPMfCXO+glcPD2nptFbCpOQ3T/Fel7gtVN6UAtLSxqbotcV
pDccTY9FJLatcoWYvD/E4HtSFBPQetQH6WLf1mCWyO5RP+BBoV2zRs+7FusCNDlA
8zU7Ep5YBA7Y/j8WlXJrTVYRsqeDP1GQYhKUpVVkq56axOagG9z+DvI6A30v3IWl
5OnWL7obboHVsX3A/J0ZQWOGzMDsJLLlOwflMHUAB9WmuytQcpRy23IMU6eN70fO
X5Z5M44wtlcMx6idEVsLmsl7+UByeXVq+718H+grCZD+v/OGU7KElJfkAOzuxqkX
uB8FZrOUjuWSVQyBWApAX69rjDV9+svnycmuif/6T+YHnMs/JuD8uGEs4DHVmsTI
QyzouJKx+tbD0TbLtRKNP4O9jvETit8hFWwgD8/uwQIoo3E9cRgAyGY5ObZQUDtU
hnTQRGypO2khOT2R8KhUqhtMwZ6/Kb1Arj4uZF1jEqHfXgRL5VlTEJfK+0iQJdi9
6PqCXlEM7sCvhsFBPXZ9VsxaVlKeEOiF0m0YhwWd9LrGJZDbsJLD6T08fqXatkc9
JvbShUOHBBJlzqQADZEYiJOCiHsHRytwHqM7opRmhLbSP17qvqcMD5MOd1ET9jzv
7+2lIkOmK5CXVVzCaDHIFwpWuxAMZFOeVVqBjlF+ZnbFUSCNr2hssM9h8jlnHpPx
U/2EKedqF3XBuTuSr+aNPeCHw9Nb6d7KbuKOV3AhhIcdKOCO5ar7r0vJzxAZ1lD9
tliBUaSN82m2K1vRvWq4H1R+lnn9Rm4ICaylrKWFdP6QDMvQ/U5ILNG68JrSsQm0
Wuw/AZHrWlSJ+gkb6/h4YiWIuF/jwnyNpC9ziwAq2z9kxlw9P537t2pngiIepnWA
NpCmV6m9l4XypAoeKKc9IwXxX+Is7u/ucobGETFATbXZA95Wgp4KgirWuWgO47OX
QMFw91KzoTx5hgCQrGYnhQ0joeLPFLXHNp84VBJFS0+EGJzyegIA7XWrCdGrpvop
TzQw9sVzJ6GX3/yuFn5jKp5cCIpgIn3l5vgynLpi/DY39bazDFHdbtTuw+TJYQUb
nBV26dcGjMvriiNIHGNs47UEyl/KXjRL9ftu+JXlUwxoLsc+2KU8I4KPpvidE0kp
CW9s3PWSFhU0UfAD5SMJL6bGme6u2fL7k4cu+X/oMNlCwM5K0sbAbvApegJK2O7D
Rp8b2MLppvdwkSxsUfud8yG/AjkDk5O+bLDjpCXjLiqE6oTAcb3RamC9BLtx5YqI
CEKQ/e5IJgn7IKP6rAB66y8tXHWxtVFwrvKCT6lz/G8HMQ7+HldTjqgDd+/V/v2H
9CZagQibyLYDWBFxdRQLu7qp/kpiWClR9Y78INK4E9Spkxl+Q9cryE8Om8lhH6ss
+bTmnDlGfaWK1kD2k9/if9RIB5iI9SYDnnlr/DaJFD4fdNZhoNkvAFzurW8nURBM
aLGB7wFnfnLJ5gYKDNxjsXVgBKX95tb4eKsAqwUEu+5sbiOl8spfMaLmp7P5o1UT
ZhBMm9JEH2uhEuoY+NHQ9K1o10QKUDNP0qAXgiORyltR5wwYZS+E/ve4Q1xGWHP8
AFMGCaJuY2evRHvalJxqkkSszpHc7RhUeXrmw0eSg+O8ABWVyoJaYosYAAdEH3kG
uv9eZCVqQvChmf/HF+CEWKsYVgNcreC7mWrjTM1sO5BuB8jiqrzABvUOxYrpEGnw
2141dQqM0IhfHM29sT2cO2h1jz0fYtUu6BhK6kKEXnctGsigUbZUuDfvnPj3RD0a
zQ0eb4Cmp0e8U4imSYkmdMBQ5hJ1vXLgAJc8pUPh2i3cQB6gbIgRc3OhyRehDesJ
+jHuB76w0egWbhAE01/usXLWgW4y+p0qNtGDdQzM3XiZC5zGeJTXWs83Li8S2f/K
QFdJX6PQOAq+G0O0zB0HBFGgVTbT0d/tfviFk9Xbf8ki85eXVV8gwPn5unPE9kpN
SdLajoZh8ElC4/gOxa5M2NIRqsaqwSxmXT4Qc6iHMfQZTkuyAe6O15vYgA6Ea/mR
3lig4tWNtOtF4el1UhfYiv/HPVKnjGWZUxXkAIKTqC3yotpW3u4uUnf3XQlPqp4K
K/NE1QevGLHOjWDHBDLB5hLuF358AHyiTd81lyVnaeeUO3uDfyXybqB9lJI5K8Ut
icBiPiYhN4H/YK74R8cpUuUgipgkdx44XdzH9GJQ5/1qEjnvuQV8aOKEYY60jWrP
4h7gcubMyQQAnWkCwoPkm6kDRvKSX0rkzQgYTGm0eMnNHOOAnf1YxKg31h9HXGA3
kDvV9Ns46L1/LxCB3F9ch6dTIVS0IfFoJAfay7PVN/gGKcJTlkyornBDxNEUp8rL
O6t632/OD2/J7axamWCuG502jbb7IcGuc5H5nWzGP1isglk3XHCLhZ+xLRDF7wv3
COQlKFVSWnLZD6qlGRRcoTmSaSnsjHARrxohXUWTshZ7S5Qv75VYdcIgIRZ8UEoT
aIt7ui9T4y6rg3EMAU3ilWsFBNOvKzslhT0PCPPADL3ifLYKr2zkyiuuqVQniWtW
AwdPSaJAAZCk3t0D6eXIK+/J8VlztDunSutk2gXdFMvLqZ64OYw4NAzaNd+sQpRp
EGBf2wI3NZiYRufrSBQ/PAd5OqBcGF3FPtapcz4XIbpxTSsTIWBRsU3VhjOH3keo
uI4IY5juqjefqhY/8EunXSWBmqyDlgZWOEXj/R3cDEtPQCMgFW69QNe2bLF4d7Ie
X8F7mwncQfUiHcLYJjA6X5f1ZcYM7U3stMfvvKdWquDOlAclJRF6o0q+T3fv81gE
K9EBrVLkh0joaKELeNBqguKedKHGYfVchAAOTS097cN59CyFBBE79GvcBvNIPxbd
OHKF3fW/a9wjWajtnSjnrFSMNqO2wVWaT9twgBDDmWzygkeHraVFQi4uxbM/ntUp
VHh84j5PLrPZlFB4aqbMmeLPOQKgawzO/oOJiFAtlAxfMn9hZCk910oW83ZQOPWS
1bg2F4Xk0Rrd/28XICzHO6gG2EkZN9agu5J0y35IFwtxYHntBR/Wp0RotsBMLWVb
pEe+YFtwWu/0WyjgPlnUeyCVPGC6L+Q5kPg61rNzbZoef8ha8rH+l3DrsJ9h8YgF
XJh18BP52EF0w7AffF7FB/8E68swnOc2ji3ShaAYoNLTuBQ5M2+ZGlguv3Z6Uic9
SXKEulb4tJufmLe3ZAtlF5hXMiCjTdh8hfHPvO4wCgXFJdEaNsJL/ZKX39k3pCbT
xO3cKQ58FC9mbPYIBKnj80otJmRtQ/ymWTUvT280nxDIoceDuB5AxRhr8BpT/luu
Iunw1KksFbE2dYwtTyqgVqb1kqQDv+X+k8EsrI6+0Yf+MeR9nHZFpwCtaMXMpzR9
7hvheR40NrOmX0Q2ZYGKYoCmHhP/YK90CPwEkpm4sW1YnkZkjLkWFQh6/Zp8DYbv
fqR0pdkCnHw3VmX/7hZM54TfdEWfIwMemeSJRp7BobCA7VqCWFyu+ddAYirsODnr
e2au2d4utd1cluaqW099jezf7GHhRbQc9s9/WjQm1kwvHBaiDLxJE95F3Z+ctzfW
Ve62rX9WNL8tlA2tUWo+fM9sRjD7Ady/Tu8mtYvaaVa8bElYzaRjqV3Zb0nDtoKv
Y8SvFJxJJwsfOiJjtPFLNuaiapV2MOD5CLl9lWw7LNmsKQnk3ogUCJ8B17Qi/PKG
lCXQV8Q0PAL7RVZzr43LBrNUQ0DuDL57TMWoiZ8VNzHVH4x3kPeQk7k7CTrkQL6X
Xtaciq9OE4UHZY6AuAldM2vIoQHzrHHVHUAtH/ZYq1do3b/3l9oL46Iq3LH1PAEH
+DYge4TMcEbfVPUhhcLJxoJT52k8IXaM0ZZeQIAOhi09De5RqP+wIbptOOE2DqeE
xnCGXUwPKI5SwHNWzhemATEpL+G01U/BE3T0OkL3myTtzsz83iuew+jcu+r3wjtY
DxmYG4lCiRqB/gqSeyfkwwt1262DrGwI24YLzRnTAfJJibnK2zplore7slkrTg3p
eKZxtQAqjZkto0cLlsHTrsssIv6x9E2Hqb4ZLfiiIBGUQOZ8tCrn3NXUcN4dHn1E
gdQZVG6/HthmZ9tss4uckiYYkmddBlQGSJcFZilEXDdbRGawZDbgurjQx0o7tj6o
oczGICibYTqqtfyMhBUkk8P+PRHKLIUrwByAsMFZoD0Kc87NEnKv+m7xSal/F9r4
6s551Ksi6lVje/WRTvMHJl7p0TdbvY2a/5y1gBXSrJMbllygWifSskLN9uiyUJpr
FHaro28YCOQvgeUqwkRyHSc4MX4YLSJEkw807xVkfYHaXtZ6vtQvGCV+mpSlj4ND
qRyW9yimCEQNwV4Xif/mCVxEcnpKDAvP5solCbVdyYMg0xWtU2djdXBptuDGkWf6
WVcebVVGQ/oZHKpCmmOdsPyW3fDYL5j6UAOPTZFOBZ/4aBFO3hn2RvZKDsWrfELL
pNm+dXfp3NeKVjJlWogICD+SU7+ZcNfCBno/pzWIZMrQPHQ4WeO+BDj8BL3Kh0aI
bwDHd2CIC6BZQKofpmQbbPdxg7ydVy27RIjrCRtTHGh1prgYhOA/FFAlZNR/pMAE
SzA8vdsf1seI0wTy8HI4DCV3rAeSSdRVYp2FPTt/xxN5MuTiKjOKte09VW+At7gN
2r0LFSrMZ69h3WJeG5GBYMfiKBEDruETbjkObdIyA1YIEsK+9gSsUWcbfAuFf0VM
M6VijngnOACo/gjzjJKw3X9O7wScpvF8VWA/wbBp9wP1GxZWitL2EfrWxu26CMq+
qKOzjkEb++bHGawqnrrhQkv2tYUdakKRTeLDoDc+u6wXG3rJf4oC9G0ycHqVucOF
zuyaIT15PHszd+YISmTI7iSu6T7BDUc0yq0CJLkgzWVgouq0wHltZMX2fdV+zzM2
vtFRSzGIUNlEkyIegn9sj0M164RicMucS8JFwQyQKMkA2TwMys6qM+k/bsar+HFb
ZFpDlEsntbEH039BZRhsTvIOHaTS6nXCIB7pTbFcccHd3UmLQCOjy3qhfbaPgJ4H
HWPmOkLl1AagKI5mkNNJDdsEwuLt1JFqaDvjqpcevXKrwd4BEf1+d19Me1RD4YTS
R5FIxvUZ/hORVKBzXSCwzvyl9Ki8t2dn0OAW0gPV3ju8dMiksiqMHCX9uDEv4aRT
aXPArXVHrFn2AVrAYjn46rz7fJQiPa/fxTSlM/sr+sLftfVxCEUb/7usBy/1MvdO
909k17ChmlLsAx86YvzC/DA1uAYwKas5ZsjGiz4Gcb7WeSThO3BbG8+lIACRus1C
8EKilKNSlAYa4vsmaZFgE80w4uvcFcglLuZcHDiL/mnUpIqmgCKuzzdUJnasdZkm
4+pNkxFceJx+xeiwBkSo6RDFkoGCWhirJZxygYZUmMoCj7hj2oFsQAn/WAFm/qAq
IJgH6qisV6BKKRNojeFAnsVJ1OPu1X4dekowj3e67eU5Z8LvCvHt7NxtXF10SAw2
sd2arDmKReEgiFt/Bn2yWfFFBN/hB2yGUgOVf6mpSWcbStK+zuX4YC3+469WPjyG
UqANLOAmxBj8/Z8HyyaZcMOx8Q1Zm9JR+dECTW4sqxOKgrwXKtNxWoXiEvFzbM17
1eFfuknPtuX0E7Fee+mP+1ZgxXI418Us+NqmexDJwwqJEnTNGx0li4sKjaYXCjvC
9Sf8z/R81XJe5FIThKtIiedOBjamgW/Tias7pkYecqJ8bPO+CPosRlhiMtn6tC3W
9HcofenagQJD/irO36Cd+PdvS/8jSDYYSJLFNdnAnQ4EtLOBmDofZX7+gqFIYGWE
E3GUbgXkcnhbyLAbZxEMC5w4HD9ZI2nAc7pukWqUch3ub1vpoHNN2KVWPoWoazwM
JKRVx5qiMjpb1xKQZipq55gZSZnwMCAzAmRGVanNr4XKqZhr+VIvr4nCONh7rtGw
6EIJU/t0hSzabCQ5w/1TaO6XMQwUhSMGN2iU/CkrXgIKGEcz8riHZnDZ5vC7sbIm
YO8KKB2svwILK6Lhrquye5uJgUbeLyMp8LZrjeUJgC+wQmXfWLlp7YBlabWp5uNT
4LncxPLc4nf2nlIdRrQ3lrIlLA8hu+6ubRVJ79fUR+KjhDtC1/NupqtYXisyrtoS
xxKqvLGbESPBr0JsNfTH5C4DsTgBCQiV357DtQC3nCvGgZT+/9mFXobiq5WkvfE1
37fgsoK4Nzk032NaLswOjmQ+vqnuuYDBce8zs76tb1fA9rWTiOubR0UaF4pX/ZbW
8vPiPD3GIepbICo/pxHlSpg4Mxa/uTBrzCs6sgi58Dmo6knjEUSiB3/0fO4b8IZZ
6hS11Yue27D6Jau8xzmA7zkEqFtY8ynYJVF8poV+IOs3GTuKHyXWgb4k5cTEG/kv
+q8JaXuvXtLr1b7eU99EVBOOi2wyo8CGHJwngT5b+QgN8nJESRB7mIJwMSL8cZi9
vUNm1nUCsgrKxZ+iMxYLyFlvyp7LZ0ot4SDtXdwhoFnAjb7nTKn+HHJzDwED1JNX
SzqYaYzqraoHlYh+x/+6hTv+5bCvfPdDhbUNvHL3l7Eq7Fyn7A2ZZsiYSqPepipr
urt0VJmJhhzAaQ1aYtsQ8H4p3P9ZK5n3nI+Buye8PYbsJ8he6IaylEFYgBwqevof
NzxfC4wHe6quDbXQH1I+drHuZ/bUa2hB1U4VnEfUnuDRR2m93SI6LW6lgha3UAJT
BeBsuSbZ+qCaCjNIK3ycxDqjGxrAe1LwwRbOGf2CSFpVgZcwGctkXKKqipxC/G2h
JQUE0xdHthopBoxcU+10aWmKRI26xhq0h75qQeN6j3cOsQk5BBVJXFcjzbnUWyHk
mS13p6mE4imi7Mw41rv5KgUr51LxMpQk73LLfZvBL9+Vd/IHQK4mjO9QIQpoUHDf
QciNinPeBhJQiaxrNLtIJ7jVGYdhbAaxc+qCqh+Z8n31M1q/+2szPAxyz6mSyHK8
KnF7JreguVL/97aw//PSJJNmDvZX3dNZxRXRmS2wly6VJu0AVG/xiolSMSjJIEIT
Nlhj/9Zo2mdOLsmjo8lBynE3J1+mPAUec/3yyAYR4301u5K0MkuC1vUgnRbwD/gA
P13R6xOuaj/w0/+QAnJ+MKe2hdobNRNT2F8VggOkP9MJrOaS2b7R9vRoLkaUg7fk
y+8nNWL1p1rnHADIHwOP3FMkkS78d7n7vZ/dv1888NaDI7PQdk0YQ6YQb8ye5JOv
guNoLpt0W0Pd2opcBc5b8vg+hb9HvOnPpQcyzWNh80pUBZk1KvWv1nK/lI2q2pTV
cvvQ42Wb7DLsEa/VXwlUQegLmjOtLpCQreBEwpGpUWdm3zxsV3HSydcZIcUkZ/Za
6qOVkUj2nCMuywwjR+bHaj+hBdxwVoilJ8zcWHqJnnHEUcnE89tGUTSfZitOvOYv
xFVQw24fI6fLIamr+j0dORG91jTvqtQAX3dkr/XNorS/KOENRggPUnAmVrNUaSua
abC4BwNlcQ7mhMI0ZbZafLY6ytNQyj+ITNTMUQg++u/RwHP01tr99Dq+EdcrpNbd
tUo9zuR9By0pV2Tk2zq8w+sCg+qh88BJb3xItIlkBE8h/m1DyuMrDRnIlDD0ikoo
WjOL4WAGHHo03HRhaLQX8xUgBp8snRo1mRvONjlMpAbYAReLJUCI4a+cu23iyLX9
czCMcBWe+ooK+nQPVylxFdsLVUnFCMS2mChcUoiguQuYqTerI7ABPWB6DzTS+Orr
PboBbiluTi8lQXY8K8hUnrx4xTlVQ5yri127VxtwUxeEDt4g2+NxbkI/7pE3Diny
+F7nJsqr9/sGrtVKuckPSwjKwAdY8OnrC2fnYLWgd78lbAYOYSxUXNer/zECaxW5
NQ69VMumeqUzV13JfgOFbuXzDp67y/o6qL/aw5bQNzW2DdmgFvuDeTxurkkC0mPI
n68BfVuc4r6NfN7i7An5oWBq+t3PYrQq9Pg80Vud/JKugNn60EkwWBHnXknKFQv9
26N+1c5RD6Y7TC8aJK6W6Wcng/FnONo1rf7rI4SA22mjsTKnHoME9gtcvdEAKlT3
moa0Nc93YHWrD2D6NT5LHlbYfuJHaikVQXg8JtGVhaNhWtPuu+MdfjHc/KKiKAv6
EwZLQYBa0rNIFe5URuGN9wJQ4OoM4yw+7p0hcQFEmILfBCsxWP9c4AthNj6HwVp/
99kVD6OoOKZKxpfDiRVVBpcO/lmTve+7yD8xarWsIHLY8zOzQm8a7XQ4Ar/raLIV
NyAQe9oG1g6iQxP78oImrVOcL/OpPj0BYKKZLNfoxIAqx0BxOWCvGr7e0xv5s3Kw
842RMg6BtepAbWId5VRERSCqk8zC/RQJDsj8PqnOFyMqOHYuzOU/tfIg3/9KXkuM
FKXw/aOy1yFRYsnJQgEO/Y8EkziyFIVmngyCeYGZ54exemynVXHTNfPUV2TimW49
xTJKfIT0yDzb9qZ2CAOqGU6dviXNL+SIoGcqjT4aNCdqbvqa89dc1ID9DAhD+dRt
EjKcQeVW3IRwH7LDyTjfmRzfhawfQETmZwiIe5q71YAxRPVGJT4A/vD+Na5jKENL
wa5IGv+ArUIgkXlcqYf3L+uCO4m6p41r0du7YbZhyCvJdHQfa6dGRO/DL6yLPoTh
54yTZZdkvnUGoHXEYR2a3pCqBs20SkxZGfcKmHi68kgK81W+c3o1ki3OV7do4AoC
6tdNBJAUsAozWl802o1DeiWeNbImLv8Q4lvQubXSc08W4OmrSVLgSGLbupWJndCS
thvqUqYJK6aMUa9le7OcFNDnDANIByc257TnC691NgC2lRTcOHVj/bkuOc1yqiZF
GUsvQT+sBtmmYEBXWYh6ASSgs57F1TVUEr6EDXliep/AwXdk6LOcm00i4+9EuHWb
gJ9Z/Yl0Lv0bJMIJCh6tVoruxi/M49+ZYnEu2HXl1TtfSBIuEqEdedxmE9KWNJ24
pUXCnnPKgjGtZXctTGKFm8QpxqspnqpeIJVf7yeo98z0CxW/YbjJ3OMoLgVZLa3d
LOc08BJpQrqnKkY7daUXYpAq4Zdw+h60aQgy3yUqLyQzuW9kZnsnEeHZsQZmAUmO
1LeggxH2MFpPNoJh/KpSOgDe64ag73jXWjXG1INqzdQ1dIRhSL4laLZp041wbGnG
2zjSfIS9h42/QtEOdJhFkkb4Bv1o8m3VZrwVd51fUdvrsdLd1H0JoSmnddsbPY3n
m5PlFp0mfaIiD1Yh1SHcm+Ht63nGuejUDEtJjryJyymb2uzgJGP7mMdZMwRZt6/i
V8JTtj6hBiYYO6V30B/e7eT48KpTSHdWU3tTEJcAyik4PWvxqkmUFAmprej15aK0
cSszTILBBqlkDufyKSQZ240MLzOT3TK3OPwrWTB2IsJIulajR22XVVR4qlKDFmNo
OclL9FkmPHt3z0P2FSNtp89PSYi7FupCGst3/XRoRb7fgG3KgShR2kxe4HX6nyQi
8njjwkz2T8Fqnqx2LuZsnpWUKIFOHYrenmWpO0GbtfdQbePTw3/Dp0t2H6AxXM91
YBZaGLNGxwL+0Cq/ScU93IbcEKB+KVt3/1CUBxtntu+ePHlk5XRDeP0s/b4adpWi
py5I+bcWC4tbEepRyhVQfZOrItS75+knl6649lmAawQSeb3w+oSSVgAH8hMpSLMl
0LWCgmfC6rb8OfaOrjyOrUbUzsO8eiJ/rxzj4TBAMeWp36SDs4k82kED7slbvyKy
WHnT7qp598jrepaLYk9KzgPL1uN2mAmQEB6bR9RXJCmJD0BIt9OTFLDURuwp23Q2
JU8XkUIKM0P2MYTZ6SBzCDTwi2alI+R8WUX8dQVIqzJeOz9B2LeRCGeNmJ5pOwLF
41CXpIf3KLc5ldykJeGDJ+BlvnNGOpi6B6I6YUXlkDJaAR0OmocrV3WsNZ8ei0YG
94Pey77+itKoqNgVpaisnBUloFPOiEEnRdIPcCmw20RYiriO+gAikodzDTSjgu+o
UknDXm9Qbp/plC2ZAYj75rN712zIqXPcYztKt8lFff1STzsGkxEL65bSWuSzHoNm
938PpbsXRnjOmGhle53zS+JmrO4wnnI3lmSkfzty2WDGs8fBqrTs0yv2nwPGon/K
f8uWv5c0Q7yLmDC+6Slt++vNx9TFdfFnSKmccWob5IGT4qWICq91zl14vxYkvGCA
bdg+qing8dTwyi+l0/rQs0QI4ThAmb3pdxjWDtuLf7zWcSd2VdBf+NU7d5iIkoDv
fZZjvv2SicZR+izOxe/6O/QjZCuP0YGPRtwkl2ifPy1qFaeB3HQAZh1QnKExCH3g
y19p7kgNXWoD8dBd841vWDG9kjkuUBu8uNv2y/HChW9cuTDpRLoXGiBisYuhJBZW
vln/XtOW/nolJSbaqRoKY5mDIgtJjVZSVV7jv3R63Tur9xi1I2fJghWskHArKI+A
PmnhCey+Vd+eufUVSvBe7CBUd8+/sJMXRSNo4YUAnobrat3QR22EeEYJ7jvXaM/S
m29DFIwRCduOq5Wklf4ZF169zA9MPVBLCXsYGgq4Mznzmq2l4DyxcUtlcIVzWgBu
hmEZTxULP+Ss8PqbuQVSJoObf5sSMiOOiBHta6OKnK8Tp2rQD1hMeUJfpefP61w3
n9i7Kjvz9MvelI2cp9hwBIhZBcJkVkmMN6fPG+8a3ob0OiWbrwGcq2x3FOYyTxXy
V5npcPGZ0ita/6qK3uMq0HseDgkkcIhooJNvX8T4D4iWAkGwZlfSyx1KiMwrcAGn
FCcltkYmVo3nLdj/eayGozCJKN38NJcHS1Fg7vFbMw7GrtzohWCuXYd5n2cFyHwV
qjE/YTWEi+pBZaFvByUYrs2pbITYS6r06GCFdGeezjY/9gzfvTYVofOLC4vzOZwP
vDxjrShWtJa0jIizwf+WBPHTs55PLLOwUB4wRm8F5cIBlI419BP67XM0T31gPJl+
qU/LQauO+GecybbvIXTOMlxNiucNpPBbXXWY02Q9zwqj9RpQWGQPGtmOWqtSqDqV
mY4SpEAw5JxEKGndPUEmB8XYUY57krtcW3cRRZ1cKTIfepGjviTZ4CdUxC2Re1KF
Apfu5g3iJmE0qRhbEOmn0CspZmwe3N9oKwO4UnR5Eu7LViUyfHGylpA7G45qpbUs
cxl+ie0BCnfkYT6TWxUos4FgJ0MilT1q8+Deo4BY4dCln0Uk3QTQXHQfmAcMIGhw
T0kp7Hqg3hujAl5V60YXTzXrdRnvnlf5fGKkL2oQZHckDR8Zb9H4p/XW+Yhmw7zu
hXzNyDMlHJKeKZsgESqFMhXzugQhyZzwoxHV6b3NOJvsc4BubZ3RZodwb73/4ugU
dOE5fwKg8HRUchzDzhY2WdNtXwo7MTDFkueSBdbYgZf/LgbKyRRUNyB/ysmPJwE2
jAlo/KRNLS5JtCiu8R5VtxRNHdSrThDNYH0sOd+Pms2RaG3JNaHH8i6zZjn8VfmD
UOcXPYtTupPOb6bCnb4+zdJFtNHDk+TBYioetOyi7rRkrIS2KNdGPA8SyQNVS2Y7
gB5m9i6JuOABxEpcCMTbnsjUW0DTHmYn4uuM1nX4PIOm+aXezqIXyccys8KQOA15
n5XIpNRyYerg2H8SQbLcQBlfVFO1l2F62GM3yzCaBmA+9VArrbI+G7sNCSrLzk/L
Z2vCrit8dPP1DTPaCFpZknrjWYRhEZ7H2DdjfeiMKJn7KxEBPNCtgoBqL5+FSFoq
EDPtgUqBal1TP7KTLg5KFplYLbuZE5nq8lph8G9ueUAI3oeCexo5iNNXVggc2t2C
Xzm2nSh+CZgW3JI7p0xCHFoeeIiDPGhtM/psq+vXrJNo+x6JjLl5Wrbi1I3T4fmT
iDNBGvAtelKz1cMd+gkpNvp3qdZ78hoVOnmiZbvHtSMc7pwKfxdfPEYhSxEHHrg+
vFJBXQJEZZ3t9Xmyizf7p/BSAC4OgCPEvIXj79esSAn+Bs1XRFK0M1yOCHSB2gkn
ZWSOpdHbAenG8qhqmYQUa4tuHJ9mVrXeqmJPxQ7o29KQGSL72reS3RKc2cmWXFqm
CR7lLUZah1waZ9i3ywrqnoy61bfQu5x6T+l3ou17kCGlVQnu9MjS7fQRI+Qv+DJU
cSaQlgYPzZROYjsawGWxOwgPoZLGpu1N6LHuODjC7xXgR4Hpv1u2hCZv7rSloeUu
lHLDxpYBy2w0zqnZDVYgWU1ueJeXnObPU+AJA9xhbsV4QmxVu9DZvjX3/4yUM6Vf
dPA84HQLCagyq6IbS5zSfmxF0PCoqN/rq1v+rZ6v4iJy8G6A0uD+vstGR7eh9Qo4
IiFw+NukRsTogCcF/DHaJl0ri8qdKc164HPzho9Kjb8VYaIrGPLxDolQ0L4TisGC
RctFeG+Ez6lbUUFYki9hxgqRlWUHGbupYRWrh/TQBftzOYyZD3W8YioJ4KjR8M/P
UNvvv8HjCP9zI39MoILqL+Rv9lssbN24A87vPt/PGfRe1W0jffUr63z4RKAMIdvb
3QG3kAkI327pWrFsJ/lyeT//GjpRY2rV4zarl9xaQ/cIRfNVJ6EZ6eY1Oiu9WNsp
2g1MpREK1QrVarxy2PWFGSRS4Zb+DevYuhv2aw2F6tuTzYu1+MpTvBR8jpJRcpZt
GPBQL7mU1wgcWTWIAlw4rB+8b7Z8ihzzEyOodWPr1eU+QJsqhgRorfgGwxH2+GZ5
LYRi8+cIOwi8xVBo1okTC3hKrXYhKNQx2lArSV4TgLZvE9ptS8PVzmmqJJLYQ195
c1GtcG5JlowMVM4P9OpcHoNez8KeIRht3X4Cpov5Igsyelq3yjw22XkeuWCZTsnl
Q5ZCg9KUwFcyKgXZribCv45aDAfIgjJbH7rCliaBDJithCMMZPw+FbE48wOxPzkU
CfcnOTJNOfhyGzDpOyK4+FV5JuM/kzfMxvNCJfMprh9gyw1ZMwdhvQgn/9yDAeBY
fMlNN1GURzYgIgPm5Hky61NMgur+ncYADcwkb3Gf5Ou4kM5yRX9ct3UdswMO3b6k
5LMyKa2vRXukcRwotPEHAdz5O4R4THt8fLYpch63vnAlJbPyVUFZLcES8kJR7B0J
r1ovW/C4zmVSFzux6eZDPWRINYOGaes5BwXRHCJ//W0Wy7uGTTEZGYMAQ9fkzLeV
Hw+sm9HRpsNUPd/G9ozJl0Bonyi2spLVBETb6/xy+vJUDdOTm96EloRnjw+DXIAy
Wj8/xAl/MQLjb/uUtOOhrRsbFSAPC1Ii2jK9KEtIlNcmDKe9u+oVVOi8dKFrjGac
Uazbjbgrvu8c2lfbzfNLvEUScLDW2gmlvQJ+t+rZFPoj4m4rKA6g7TsoqfFAV3xs
WD7Luqg3jcBSGSQSa6w8P2Y8GXRnCA+DEDFhp/x81xL/z80WoRbo7lsm7znoXUpL
uoOzcfTiBQJkhpVOpVsFZd/wOFh/ByjBcTgd0mifCUDqcYY1HqBz7arzSWaNWA77
EYgRFn329vAlyJzuDb26jAQ5Z2tdyYAMhsGzdZO8X0SVUUe0ow5+XM1PhcNt1jVa
jqg2pmryk9qdxwgWf4KynfyiHDgg8bIPT/dkI5Mv4YCfHuv3OcVkx9mELYDJ0DFm
kIWlgzB7wuj2NO45SqbLP5bB01rez0UBPSY4qS+vVo09/vziU14hLITRPql3t8XE
BjcmDpjSNPmWDNf17o0V1qw+JujinvdumuK9KRukJoinhtQ5lx3evYJqdNNYWJDg
WQEgwyo7FdwLxzShi4AU977/pudmkWTj4xr3ccmZlyASjtYOcr3+tS2Rdb6BRg64
FM22jS+pSiliiZqQbd8Q3w1fSnReXBm2Mi6P1PthrR0pieh7WjvhieZ/ZETJGtEk
HWAwietSRdxXxPiqI5LTOuRu0SPFInWGq3nB7s4nUSjGPbvdub/07kdsnTTZ2dS7
2x5nHfSQfTUDR99+N4q5wH6EMdTsRitFTsX0lmd42N1iXrSEh0zwBZSZBBfhQ6Ha
DquTcCL3v5rHwUH/5nXLMRTEbxzF86qgk2l2CR41/HcQ5Efr8+j9J0+DvGAaIbXt
Y6grTXqqUZ8ksk6VAYDSTg3QOwMMM+1s2CPNOK0JRN6k/vGAHPzkqGM5oJZ/9gUe
4R48IOBJ24rws/tIkfl+poUXGQZTqE2jCGzN6BXJUOxpcgG+I5NgIsEx857CjWob
RNoe8EXc99JRrkaFbdiPjpmZwD9rJjsdhDt6phDVGYPul+nB4F5z25z3lI8tTz5X
yQQX1lWfWx63JJXGCuzMnyuMXNZXzBk1oRHTNHIwGVru3/7XW3KxohIUqwysX2zP
/l2WxtOOuKNzroy5pyYwTFy+N35khv4ZzCtyijhLuZLAdXozY0S5Ij5vvGJijDEe
tfrQapxn/zUqHzqZ/a+psqREeJ3wNksmR29FwMna9F/cMjklDuzurcgkDivvQmci
IVkTryGNGoq4Yd4vc5I2PwSa3/y0fXhGv9bcYyaqsJenVY11lsFVqYW7xzGuUrIJ
kv8cQ8U++/7ANh8yit6AMn7Rlr4nJPLyUmrPyaLZBWO0GBQ37VQea8A/UjGOp21H
udXI4MVLMukIpCVhAbO1FcX+vHxsBJ8poz5ZkSbChUhy+RQkEeFjIC6UQgQ/9QAz
K6uZQPrZHKU8OZvNWJqRJ2gbO1pGsyn0F3InWris+O5MeVO7XAHUihJlDk2NCVHq
uYdkMvVopPeXZ53Oqr2L2Ty1VdrF7Qqdf1Ho50cosWe3pI725KU2KaWLWmukOx3X
HWSgUMoS8Cq2rqtxYTUDPfjbKuuZTdOF3wnu0POoKZMTlD4XJo4qlolkhCsKZJ7l
nuha2bsuz1fGW0bm0auDfLNQhYl/NLwCcdhilHzqo2bxXWhgvI2K//FFzm9cPqCB
9l+LmzJWURKymqnVU+SRfGAk/WmAyDdl1RFqK5ezEW+c6DyXhrzZ+Oy/qzo6sveW
hFpqNPF49je7Qq+WlM6tdX4Z/kKAb3oJVYO4Qygq6OlmP4K0v+9X3uxjfFI4DROs
MxDMz950275Jkp8kaSDGCTcZmKin/Tgvk7gs99zZpIeVg2TaFLlilAk2xDsj7qcW
CpSZvh4O1mKogAs/SGdZ++m2WDkLrISXgNKvzqmzl8c2qIwb1W32n5L0h/Widuww
atIAzO8MDMv0eoNVHGWZxW8jccLhnfWrBoYiIua5XNWe27kN49EtRU14yFsRU5Kh
O6y9F35jpQLrLTtUTcbw3AaA95Z6vRLRgzDdW8gYYWGr8BS6a90LsNrDwSGRKf6U
oHn8Csb4T74d+2G1pDlVzeCzzrtKxN8wEENk5+d8HYAiu9X6dxcKNM2CbnnfUtMB
kUhiLxG7lP0KgDYTTKugDNZlIMhk+iqCRBR1+UAiznw+UANdw8sZil3buAMn2MvR
4Uc1ZuKzx0gp683YiCgU/6Ims5zo3hCc+GC69RHV6aw/O0DdGofkUPhZCaqbe21S
l0bPAzuuHExQ+3MQXRbI3RywxNKsUeEIK5J67rPa6cFgOr/WVE1EYpheSwHEIHs6
Eu9lzotlvv38iNFbG88IHfqDgsbL19IK0zaKXq9nuAAkHur27udAUPsPTU05FeAV
Eie3gDL2rQht8Fi0CR+qYMvMOlbC5s4JkFKds4DB5hVUW/oEjSUK5VPkbeZp/aad
10Xc0s1xCfoT31uy6qwcnl3RXwzCuxuWT/fWGU3Smu4JxCWEDH/815tPS0cM5dyd
KjNJJ9HX9exLEO6qL+43ERFjHjC0bGBy60C2ohTp+pb7vGee8WrrXmqpuceIjVBx
uj4Z/YxJnUPWciIqQYibsi8SkHIicEpSin3X/7pvg2vD9143k4auuJToKOIcSWsd
WduYU6OfKIAWw6IVa6fmBvxoIeCIYym/81H/0v9t67F03b35n9luBP+hgEDghjsu
H6zHRij3socpZlYJwkMit9VBqILKHexgUCHJLXsy0gXsxkdD9Tr0Ur4BxNjTUGrF
nTxK9Y+VurIz3/lmjEaKEiWc2rvnBvHBjd3DMpz1ZfCX/rDAAOl3EEgRTojBRHoP
v6ceJay0vn3lyG3dzFSUs6nJxc9ebjrHQ1lS+0MOSKSCwX8nHcU8ygYHXxtTLkU5
ghK3U3rvxaXQxPtSVElDMyfpiPDj2+ZScypCPzlxDp68Gv+Xr0+dQKqKMKnlYzO0
Eg+fBNUeynWsREpjDKvXJEMEJ1awTuzZxIWVwxS+y1gb9ACnsEus94eUa8ZpQsUc
JkreIku5Ap+2C9KeMl/9LNw6WxhHLWO8TC/ftBCt/9JA6OIg79pHsSUiy0Kni8x9
NWEiwfoxhrlmACVE5CIOBvNMPRg3UcaBfLmwrYrb7ik8JvpowTEKcQn/dbTN96ms
hk2TyQhxQHncckI5k0voqK0pJRlkTb/aUNdtn2FoEpIG+y1SKiZJlCS0J3HkfCP+
3HwjvZd+Y6fhLUMTOQScIBvZ1gHEKO5DXpJ79yR75QonvGTWkJFhDXIYi1XsRDi5
6l3GvzxIXGaB4DgE3mdhkAOq1c31K+2n9wYGNo88f7c7k+mku63DrXLLni1MT6K/
7LbpzUoGj4+hyqa7HovB4iAvdtaGWAEnztQKF8gqtBSB4l5JSOlpMb+fJyMGJdYU
SC6ysBdMsrABLtFwghQnxSG4QbnwySwAiUlUOFDuord3kf96oXlgW3XeV5ikHPfx
8PK2GGxDrn4oL7SUAbo3yjU0XikSEgWAGyBl/sRsa2Ka89/6HgmZWX221aic9wIz
9SJRTvkf8rYpnxqwzumNEMh5RCvrWeMWP72ZKitqrXzyK1xxb7QKGEmrWGKMcvgO
xc114Akwynyc4Tlju069KtWYp1tHKt/sgb5ZJG2u/8H+0SOiHXXIl9olzn/+GLCg
s0xw0/oaAeahZXbjZPT3FEzmSlkV+VfUFHBaySjNFH/FmATpJfPKM3KyqZoxkl0V
sC1UC/6rSfCrZtUduxOBpJ/Gml4dNQ2qkqYP3GUEH1Pht+aqR8IL5mBkTRHh/DKW
lV8OKdn9Qte5YE3lB+OXbfQ7HUPA/lALCFGHPVMFetmEmRf+ya1s/YDdtQKX00vw
GUSxHmv5hq3UdwuC4kUdIi+gPe0a0WVAVDGP171c0sFCjQBwvrKaAgw1I/+K03/y
JhMy6JBkEMkG7ClppwWoeqgdQ7VHkwybDtA3d2Y+RZot0G+hZ8LGZUKKthEJ/KGq
5IDtV7Jav5uk+5Qz/7D/FfWegBBohoOkBOZqDNyo6jHEEWFM7ieEJ5+hHP3flvlx
V/8a0aU2vsA2tyeAY0fQRj8n2ex18Auffb9WRF7YKJjPS0ew7j23tSfQZzbIDU8z
HWDng6VRgYM92s4sXJ4GlKQNpfI6ao4E1RdoDzCSLvz+NDrokgvY4Cro1GHkDYL3
Hnwh/CdZxCA2nF+WoTd0mIgFnGEjtUQCDr+yOyPpSdlo+ve0/SWF12IjTsgEO+vy
52YxvvSEky0TnP7ShRKTWuguqQwsn1nnTu2Tk5Yy1wPm2k0bAA+sREWw9jizUfTR
HsUYUETuThBFtTxy26l2p+tpzXKk1XF3rm362g39PjTx2kDDEM2991WXnedaYGcL
aVsBiPaQajb2O+PQaLcHAPlzaYgLnKHF6+ol+THPPTD/r5Y9FhkXSIRQDwvoeRYh
Tkb/7L/krTUd4MLhn+s890kYd+ctz9jF6Zgai1jP0+P2sUwYIeWti4Rgy8ohpc1N
ZjuHTTIFj49+gurAI/HWoUrAF2Oh+qy77ZSHHWJf7JSCwcy4mT9KmeIJXnPbLqgD
JdlX0ge6JtFxBd1oIZGlbd/1G9Rdkha/Nex8YLJb0sY7naGEy4LnVPSVvFUT8Y/1
rrA9L3yIjj2D9isdgYL7DStWO0ynLkEXhwd3Vblon40mn35l0IzDczYRXXKNN/vi
0r1yV7fsmSLiwpLZveF+1XTsfg+UC8Mqb20sV1VR3hqxR46cdMG3FXixtkQaymll
S2dl8LM1sHw0IcipkmyVEEFVYXFnEdLxGHyWmfPkyAtbPBNe+wmunprdH+tRAhy+
npenwP+p3qjbGX1KkGnRD7+/LEElLSaIc01oh7Q1Q7IxcmLiV6IEU4jx1pRkMEGA
LeppI7Kbc5lQ8vD2oSam8PRhle3K+F6ExIFELk52oZ6g/+A3/zs82pPO9E3kMJt5
bkmqYk0tYhbv7dK3l/v4LlmsVYOcIsnfIrCzTV1PXzAhRpWpy0Ld+StfqHibgILl
AqNSHCwMD//9FNoyf96TlTHHMFggpOgST9Y899c2tfJ6qDNoK4rX9kJIRJv0tca3
tbgePdtt/CvOIUmW4HvEx8DaxTT6FPiDRFzqq0dL96hplJRTZZD7iL8Scp2Z/tTO
2wDbom5GQPTTRo8K/XlZv4bvrBFYPUZ/pG7kQOYJmUpkpgc0fEJuDX1kywjT2W6m
ec0YhvcAVtkBHWlN2X/2Qsk+padq4u6eiYJPms3HNxSkCApV2Rf0vwcP/QjOD1gE
UasFCswrTUmB3cimqBoF5q5W8pv4hirasq/+TprV0EJghpoUoFp/00ZBf+TwUAd0
CXwPHL9eoePojkYcGxv53OtMHnPhQQD66/siGyLRcC9ZS5MzuQrdLQZdea3eud8a
iToMFFtt6gB1TUnM/cVuQ6zO6vGHjr2c2WuN5of6IWZoDKUH34esDJ5fuI7hACNH
aiUtbjCAOAxShHmXgD8xpr292TQaIxF7D/NMRmhnHbZRfMqDr0Ohnm65GxerPars
zOEl4qtzos34eIJL5rUGl9XNR4Eyg2SgsZOlHltxhrj41wLm8+NbpPM6E+bZ5cey
d/1vON0F4aJX/m+jWqSBeB3X622bG3hEgnI2Jo6pIzWgGO0XXctsojRu5n9qt5Js
UwIirRxQ0fNNeyTta0NjAW2Y7GG8KgsY60QuujoPoEpEYHxcDjaN57d+XKLBo4I5
mtpBDmu8SPuVNoOmkMfjxz1chA/lgRv5tkaBOrrqqbU5GOHoeHqnKoAVcfmACGES
7Hca8sdyvLgOag7LwOuWUVqt7z/MW9KL8UvTN+MidoaV87g2cOYWD64Sv9WLjvQy
YDdO0MapDAGwjQgW6x3qlYRYFjXl3Oir7Iq7Y7qlbDfOrpg/Tika6o1IB6TfzX1d
xS+sjKDIUU/vxkY6T/hQbASp82s2v1Om49OWIfc6nrq4adL0h3CI2HoymhNk1c0A
CT18flCNXZjIAH7mm6AeC6iZiE/eu4e9uxTdERPop3VZult2PGkxgy/k06R1hBh/
+slN/qmYdnoArQhoyeeYOBencrGSCl8Zc94ccpFYEiuDXAXdl21woerINjxVnuOX
he1kHAL0yTsagFy566wbhqYb3C2+YNxloM105ZCwnt1Li4DBlFN0UP59aboY2/wQ
fa5N9IPRaqNAEki2IjwBinxBOLg+q7oAaJnInQTvFUgrKV2shzWysxl+rWrIWvET
OEMg9Kp9I8H5+wEPuiLwCz6k8GNywhlIXSRFQO9lOrTq6c5fHROoC0RnFLoKq08G
Hca5aTRvxuRZSNthHFtcYJMQPBeJgS+tNzwgsY0zuuuVsowQhTHLGcLeUPd7/5zk
miTt+KHEyGLqelNdspSd6wt0w3O17p/xi63BLlGDVwwMWOtHIIsO85ML8MiTL/qt
m9z1nA2Vl9pUu5nFi5cenWRaGd/m5MDf3evMr/pw9SSg8tCRMKp+s6aY/9Sl+oub
YDbQpdco7lOYOOK30n/12l0W/97OmOWwLVoD8BwljpNf8VhuEL6b0mGsZXlt3T0L
2MFr1aQYmK9n2A62U3tTGxS+iXx/VxMW+41BB0J9zRIKUNeRB0sX9t9XMTnzzgrR
1rCUHjYY8lIY3UN5xZaM++C2r06RGoxGddBeY1dLYkgVXI8dDFxmOQCocTOALvZO
auNVMY7P2b/dhxDg17lMpXhrFNsCOL+I5tKNpx7d5KUxdxvC2Yjp4fljbVkS7L9Q
s2ny7p7+nvaissWT0kIQe7Pgqi3xa4ApSgulNykuNGs6PhZhId+zlTjMy6VGqjx3
GVmF8QnxtoUeGsmQsIIvJ4EtOwa2/YyAE/SjyfO/wDpowoLGlGIq4x2YvapkSXBP
6PNelImah91TJ3Bz19CZoMZqfSB1/GaZD/aaWK64ua61hH9U+X5bmD1W6aILOLiu
fc1Lh3UsCxnrZoCqRk3nXD+ndkZ43tPzwvOiy6e1U4eEwV9UTwMgbmfQD4DOvWah
pTd+yrK19KtiWWUEeNVfLU1atI6cW/XOXENdTgBzrIoAqxfqo8N2TMgDCv9RMef4
WNOSp01ELXJz2vjbhblJveVil9obZmPco29d3te7ijVAUrzTVphAuwYrUv5Npmdm
MCetAzcw3yMwbFcGmioo6IF0nR8e9tMPNEWWhQIOJqe/pOsjkSYRp7a8EpkYk5DE
XMwuGrTyXQKq5QOxPBlIIP9TM1Hn5kAdc5+KSbj3Hr9VpBd29IDc0fACaICZwj5K
J+j35rhMmNlfNAr/g7nYLe7HkVKydy6WU/IlFWrVBB+l8GkoxdKmviaWVvnUbQzU
JyLkBXuoUvDF9MTANpjHr7dPG5t76VerIsUbMPL4HB+GSvc6XssadVMO8oe8BwZq
LUcgZrbbVPniwLN358GlxuGYNjXqnhdzyTOpLQBystEiM48b8iJcIb4pWNyHdrc2
FHTiYM1i1vyqkREtCx4VPpOaQOQos2N7GhFSnqqKl6uAlHg99zQp8t00Ch7XOU8J
Vuk3Hs6wL4Lo2+O83fnXcB3qnXw7rbkPsHULV+AwvUS6dF0Ri9gpaJdL5jpZKYVI
dkyh9OlQIb3ti4eilNX5/tmQa7w1B0tRnge0/6tIAdOovnjyly74R5PnOzGPzxlL
strMFROpUYPFHG9eVCLjwWEnFjiPPwwqZlw0rqgoQ93zq7Dreh+REcDb1K0Aq9Wf
J0/7CtBYVAz2njIEbaNy7DrQTc1EJkRamt832+22vnVYkb3lqPaxM5USZ6uJ2bX2
CivOOZ0Ro/ip7VUsQEGeRxe0303xh5GCtABHg+f+lLKaigrJ/bQVjFz4GAjyBLrd
ClKiki+hsGBfxQYIV4Vos1MctwriceEz19FrB1dRDB5gDM90MsIW8fbb3hoitstg
O1ekFza4LnRmMQZefPqzEI2r4HuqWXgU+Per1Tk1M5/3R8lzJoASoBWgQW+8gak2
9sbh5GUT1w6lBMwPGdCstXG+lDT4thrlwgFTrifCRAUrx85Hj7znCsB2funvYQmC
LwCcWlYoZrVu1Uzz+ROFpqYRMAW/c+32rFz0zn1/FQxshwTRAutf2uOeEb1Cukhy
Vj45Qo043+Z4u5DD7UDGuTraZ2SfdBbsEmgHgBGlop0KmcScocicy2V2TiczWcdp
wGzrr1XmvYHYL6Sfh/TccrldTBy6Y0PI8yqxDZEBhpgUVbJJRFAVMyhTnNXgC3Vg
0SQhQfX10JGobxfo/rtyV8n4S3kIU8LPJ+xJWw4yB1WtVVwSCNQeyj8whC50GCsx
zUVq8hraSOmLv77P/VSyd6wSOY8XrUhw1Mzr88BPAtAXN+pOXOpMDUtsQ27nWRW9
VKGpz01Ll25IWmLylqmFQ+Jh5Bh7W0IAteMGE5FeFcUfKvwuUSGOdiTPuxwdjuOE
7/dkdP88xeMWYJs9SLVDqA7fl9rBOiVMg/CYt+odWC0XTfM7/c/w3hlGnEoDu3do
uIUSRoGV3fCTzj9Gmxae/+X6Gl2LaeeaXomjIN3iaKeon9qkZDbLSnJk7u7ZXzgS
zcbe3VYlzzhkIhZPttUxZHCR8Tl/qXTHMk2QPzbqUEIJ7UHq1Xuf8tOUT43kWjZq
DH9zrHqlKwf1zP/8lGNgYToTt/9aEOfJ0eqNwOEJeXxNuLh3kn3XR2KZCo42nRol
mJnfyqWIVyIyd/Hbdrq06HL0kPKN2fLBXq0LCJBVsOjdsfIzgBUp3YrMr5beDUWX
sDwTJdK35+fsvdhQ1IbTCO9+DP8vZ4iL4vaZc90w7jkU0/nwKaYyj2wU7fXFUNsz
1n/pwmLCqLxO3Mu0H85bBixaLNoFc4/ko/8CEas/gPNra47eaPqNoRLAZ8EDu9te
WP9l1nA/GEtUF8LtSW7R4SewfjNrwEXoZPsx9sEHvhwTo9fv2yvPNOoqCa8MreXL
Te6EWYYJ6A2UV4MNYBAddUF/04ULl32AmPZqcfTbo8wS34juLd6koWpGyoghVVKJ
lp/BToaysMRmxfyG6g9CiluzIsowJMsV25JU79VM9Zu3/7bTulqfwN821igblZL8
Dp/+69Sc3zWNSHCF1XOfeIqn+yBeC8kVeoE1S13sphApk/pLiIDksmAcPcZRbKfC
irmlXN25/IpQMXBXKhgE3AtQ9emyCFnYg3OAH910JRewICaiA4hcUkvLeO5EQTnz
mUzVB8aHS7QhmUBZrrCnyvqnX2x4cXG3KsC9EzqKk6xExejhyTTNF457Uf5zlHwB
w8m86ycJoaXRzWJGVa3G4OMDF7cnJJlH+1q+pdYYh3AZSjtKsQBjtCtLPw6uwlN3
v6PMyN4mdEo4TY/61Ft4uOHKYCYi6IUCi63n7nmFNTSGFd/UuTou9Sp/PqwcKGo1
H2vGkzJe7ckPbGSC62kP6+B2QAOj+A6eZXduy9PtQ73IuibwlIPrGPY2876pn8SY
RmS21mPHsTSVkPozs9/RJo8+rMzDNh73DiIILFvpiE2ZZb3WOCcXwj8kvEM/xFhh
ljogEjvL1jsncAHY8mJlD7M28EKEDOk4WJFRniYUBx811m6NoUqtfbSC8JHg/C/D
kvY0dvc7nTIe9RTTtLFGPFCec73a9cDCBzbzif3xxKaZGfArY3tF7ZFL9CqNerdG
aGvG5ijRl5DrJiMIDsGKdqJfr1pUGeSwjo4r6aX+b84PjxGlaV8VVJ0/kVqc7Esj
CIh+G1gcHXdFUr5e3wt2paq8pT2GPs5xPWzyIlBkelSxKYIpoFCQxNXK0nd8uodF
N6+p9cIhNoYjcH8a7dcGCurU8CSmtcwtWdcV2OT5OwUpM79wpJxgGlNK15+N5rxs
xZ7FF9Rf9GpOHt/TYPEdb/xvF/t461+0TkSCHqq8NSS/BLkBWHuKef8iYQQrOA6x
6F3xGexr49yMavCvLFw04KEfKmkvRH/efLW1YSomKKI1AMmLYovvsuJbwAT7QHbP
pizc+wCGtv1SV1Lf92RjuLiRGuZPW/2bv9YMZjr2MJ0F0JgLF8qUUlR5kZDRTOPF
pLEfRLBby4WIEYdu/BSA27LgQdwuxyppO4eKPEFYNuNPa4okwOA7p8yT2aqu3Qv7
4VlXEbPZLC+W4j2FVPCxlfWicoGAwopLUP4z2RuwClx9MYlGt1Luv0Bs8Eg5q7mT
O77cbB5D6L6LZkGZ7NVUMJszvjV34PYJYGv4vvNLyBbN+0U7c1zXjooqpWlPdYzs
4PIwhhmIiutIp1LZMIkTXXkydT3oe0wwTRO6qmus2kknvh0QQyYVomhOojStrfoK
LTTifyubK7Cu0m/qGo2N4AEKja6Ewufg3JeU83bR8/tIiXhsbh7WWosoRVGcGodS
td7WRmDotU+fdSDQrnqJUHwVJVY5O30hfwI3NO6ci2/UAPHCnBiqDWzwPrvnK+S2
kGTs3CPAisWJagaQVrdLI8yIuhDsmgscQmMpsMnmKg8u2JSePr1VqjBA7+VEwKE6
BWStsDfnhlvnKqgxirpDuwQ69cdskpjNZcQ9tdUKjkIs2q3upucR3det0B2vkqaK
fYomEOx2jVOsVym/RDPgdKgxZI67NcWD0rvb98olbz9CEIULpBOZQPTCGhecpFA4
LHNHyciNs4/khWPCxrXpUurIt99rli4E/qpH4PnJN5IgUlgrbsQypO241fH36RI1
Wh3r6+llQsgj1OV7r73dWcGiWAoVezwoN6o8U5C2kwy4YAthELmasGxOg3vq87LR
Ta5UhZjqJuhy7KI8PbTlwrJHEiMkF8d5kNBLUF+dw8URmOZLJP94bCbdTg1i1g+r
PFyc5BQ4AXIx+WpQt/I+kQ/YdbgdDeaJyIQMctZiar86ShnBiVqNa6OjXjfrNoJb
nr6yJBYLb98YPvjcjCNeQ/6LzCUaaedyhBl0fCUSMaV+6vizqD0zDdpb+v474aip
PR3UDqPMWEWkeLIzDrWLTc0faFLNI1sHRKaa/m3Vzcj1ugCaIPufqwmGnibMLDUJ
KMA3wOtNztD5/NrjtbH7h+1OK3qrcgiK+ayu7NqSYmb+2jyaZyY0Z00jNuz7foon
vy0noEHGke1nNyntrVZAuH65hsDfqp1uWoL5WFsc7UW8af8fJ50zNvjd77TZpL8Q
3m8G16TTmG4a814A6IJ9DOfMCjdHODxkM25B5iHM5k3yUtXTGaixHo+gBz1r6w18
KngSm5We1UTgnCvAG6gmpR03tY+bXIkeKEFpd+seORyHqe9srxDQvVGZh45FpIsK
KReESxGF5YccoRH1744BUSZvAri76lhG+ZVpTO1KLVXcZ+Q6s0fRABZEVGhUnBk8
34fKL7E/eTSPEiJXiEq/lsDMuuGX42UqY2AFDbZHh4sQYucdvFUVv5AeJZUyhBu9
HuAnQcIBRdYEhHsW1UWVdKL69r9K8uSabSTdbN0LyzByebcEwci5AwMd1LiHZFCi
Srgj31DrDU7RJt0GkYhAuliY5Edc2bwK9ObKOi8jlHuBw0ZnNNXkpqBbtSUDrv4f
hb4xo2xYvobls9PZthz00srTT6R4jCogSAt3pdDyagVhDCmB+4GEJHi431J0+Cy5
xR3tTaVs+E9XO5A9eg5SKfXWjtsRDVaEK7yrzoHzikZcS8gmGr70U7ZM4JdNXiUt
OkaGqk8VorETh26KIUak1lasyiwBHiW/RDQ2EjmsNQUYVvSMnETbP61c1Y/KGfrX
BDilaqDiomSTIUZNZ10J49b/o0taajOQ9dwAB+wZf76rUH85F2v8pHFB/53N9QzH
4F1cjz/pqRpvIjexKj1+XRxxVZiWCsc0lO+X2y5ETy0UbaUZPvCTnX9BTai8WLlk
cXKRkeXKznI5wxz9uxGrRlib1JCcAT5quKIMSWdeiVLxGzYp4o69kNJozRYuv20F
QZb3UjJBx0MucBa+ylRbzocaKj7SG4JfO7KZ/InWsOKzTdvCI7Lp/oCKArbpgp5r
Y4FvX/M/s6vQcX01/EazLIl7ndd8Kz2m0GOilpGUtmdb9TaQcM59HsS9otos2nAj
hGakKAa5K+jaX1M9Z1XN4y4+LR4KpTNYi9HziSLTW0MDnIu3Dlu6USF5jaJSSVRA
WyKNYaWf7c6zNEhDVe1BJ6SGll/f7ZMcsI3LEdhKLt0fmAfQ/gIZmMtLMkRAds1+
BMmg/yMalQfMWXTLWOa24sxjzpMqn4FXpH7QG1wbfa+UX/+UQwd7Q8zQRDyctUhf
5pEkj7HWRm2TFrJumV637jxnnHB/nuK+OLNnUIyNvt9k1d9Qde5HZWTqH8yBDbep
8KPONtOkkidcEWzVGIr8HGUtMK7qHxRD8pY0A6IF30+OUA2gPYPMmV4/xo/aurqa
7DXtmPePNBrST6DITi/Zd9mXwejeHOF9XngfIpRU2QHE8A6Y7qsy3ybuau0RxTHA
YRK39/9tuFpiOSsCw2Q3Kf7xrzwxlqJny8ngrB3f68E8bbBpzYlRDAbXoU9HZvFP
BKos5G8bXrzIt6FTlbCtnrKAaSejr4Y7OFj5LfFn1dffQl42JjgOWdGbhO/PBxD3
CUQ0d7ZVELyIQS/NK1NxBx80VWtFvFkKf+pO+8Elh4/1UxJRSTUEMS6CKfrJbArZ
uplEVWsFAFoGGu+eQJdz/mv1nw/oWS38xQPtkKdO62OROPKbt/b0ymvW8L/TQI7S
wbXcJ1zq9Bkuc3h7vIUHy6qtrinjcyw0QOLCPXQptZwIhVytKRWUMknCdNlzosMw
Hp7TkVWZVI1lAA2bfD+eFKdkI8x+R8cm7v3Uko5QJ5R14X+wv8dIDp2ZXOq2fTyy
BSWNG9nWv3jRYWTcfkhp7gqD+8oSG584gAVNBS0UfolL5XHcWckIQo8DhwJ5I/Ch
hFqe1odnqZAi9gquuBSuMl8rNj97SoQ3F3jhoiQWojnWWpGuQJ6KVuHCqpuKzhnX
KUmp9Ggo0+yPE3/CWYDloE2+RCRtwpW0cDeWmWknZZ0llcUc3iBbliuREkr/Ekz/
dZIJ1xuofM3l96DB1WCm7TplxjgFi9A9uPf60bAwvlMqYXywzZoTwvC2RWDG+x0I
ULKoYgIPcUn7snhFRb96HocfiNnk9QVrvmYzI93/ewyraA+UxtIk/IDW7Ys0RuU1
a5jFOSbnVmWYqjHxwbnlitkheAaXMclztagLm1eF18ohBIY+uyNgcvtYaIDOAYnF
uwUrkRhVeUGbsFB7FO7eK8EFjtJlhiatLKwFOmgWorhbpi4NF3ATOQzDnwx9gLeE
ijmOfdUOWRXIpoyq42ibCnBJKbV8lO/FWhz6Yw3QXIvb3g6vaKyqguOs38W9uWWv
Ms8iHWp/00oJ7GAk1aRiVw50M1kG+uHc5j+RxKBmROQVd2Cp2kpAE/OcVEn0CojK
Ce2IotzXoRhGX9Cc0HLtVovNyKVoDheu89L9DkitG4l795N36cs73DN1z+yit03K
An75vVM2AlNcavhh0jAWfK76tl8/jQbGaYTBKaBpcN+uHcrjK8HvS+bRNjcOveqm
y7u/ufOryjF3tNWoy/C5aQPNZXPN2uM3dp/sLHe/RB8oeUNRC+Zvdu66hlHzSlUs
v3p1thitP1W3vcuDyH/gaiCt4yeQtqZY6puNCY7zLzBIfrBhyXomZ94KFtcL54K5
vw4+TU1scyO3dJAQesKcEal8ksRI6wvFqCm9bYiNRXalCm6ZMzN0M//CH9wIP6Kx
veq4eS3TMliBT2lWoJ8ttkffnwRo7eoGkmRWKKc4nS+mx7QP/pcfvRtLfL6WELvj
HXVnWNc19WAd3oSqnN3DUh/ZFa9PuH0a+YH6rUoYe1CrhikkTq1mQ3iGJAHSikMd
YPJgWaoxRI2khB4PQ45V+u1O7LG1bF6iBhCTZLdPeaPO3vpoRq+02w1InwsYo1bR
2UYa0P6UiPuwODEb9EUQmJGXJuMUoIs4MtCVDrM+Jcz3L0mTjpL1oLK/Cn3cjI3T
0nPKDeq2DxDoD5K4E8xgl+7AVLB0Ja6OQkNhZZfjMDionA1WXY13tSrnL90O7Moy
HILT+t4BOPzAOASGmFp5KitEBWzmgX4muZDpXCKDvt1MYJDek8EUQInqKFspPvAC
P/URDq/7pMtppcYyvwbClMx6F8Ze+NotYV2+OUec41wUHEYu7JVQrZoT8o+wSzJ2
7vmTpFO9M+AJT1keKXfotmPSI4kpaUQ8n7Ikd8k7oVKcQ/X1+OSpcQg2ajk/toYN
cwzfSKmy6xo/eyR7I91N/IlmHV8t5GrLLJ4L2uEVERloAtWbMJXmMln/UEco5Vwx
LwPG3Of2WDxIugWZBIKQfQ2IOLyauvphkJU2IMeUoc7uCEqVR0cP+II6eFcoJmmG
G4MD6ohd/yr59EFK2hjcbGHgc8NbRjHTHcJV2yC+vhLh0XQ4Olk50FkYWnO7nuvG
qD79Auo5M/bYVVdCrMzI2uaRY7Q6jz99YQEUt9K9CqWIO/1f64dhY75kJjRmXtAp
bp69rNZPiX61Y3oP90eY68wMNoC4hVwPqzwX1o1P6LQOeOUqQ58jTdHotswVcJaA
5+hLBDfSwmI6tVUacAmDvScJcwJzy+3FkY5r1s3j3arnceqLJa6jucgKSUmm5S+j
ulCFi+l7J0x68xM+yZMc0Olkm+DHEpFv8p1mhKIFC86B2Rqr9Pj1QkoyZ42AEUrR
1vsoVJT76J11nSX+paBQHomSBTvzaMEzzFr3JeGqYazsgskxBB5eSGi+R5ea6/OB
RT1OuYyw44pUl++Iq/jP+Vz187wkfO1RZ4UWz3cS85Tf3iWcS6r9MbcAOww+vA8X
suW0yN92wToppt/vmrzYRQ38tlSsFEwUyp04HhPPYM1Ij5YAKEtwcPr8tq0D4stl
OB6+aRZxa5AlImgJGlz41Ik5jD8e1KKusbPHBOfDsGZ/SPTvySIWD3NtsejU5/bn
9oLucXHeGb4MghhkwtZUB2H9oLP0H0+oj8gpclcmhPIWtPVvkyVCux5I3jVfAwXZ
IjQ1rkhh/utrbo+ebzwR4KSHwXg8QY1jrUCh5m8lXf7ZDGV8cJ1JqXj+Cp+Sla+3
zYzcenKwDPk0rc+dlfFP8Kpz9bgcW/laruhqwZducf2K2D/iR/4GimvXdqKfQei6
4DC/gliK1hGPdUVThvi07TozEloL+Iw09R9Gx+GrrZkXbF3R0W6iBgV3ZLZmK6Xr
8nIrAcc2tWTR6PkSxeD35wjaqigCuDym0Y3p/F9ktDvhNWLB+9TnBh4vm3zyZn/L
hAK9n7RUlYhMj4j+IyOBGPhSBuZxxcdJeVEsnt6homL7AemJeIhbshiGiWe5eadR
7R7NVOX9GvGEZW3/XGD/Zq4nFnVRwqSaq1CNtR8UmyNpq0GfmtCYRee7MQQs1NbS
CdQ/tggvlc5D8RIOoIx5IWcqAzWRm9ZSQC44pjBVuO0Y3vw3NAiHZnv4VCC7t0ym
42hGsniiEh9EBrdJuQm9GZ+P5b4W3oIB8irbGiNGtoFTgj7l6S+2E4p96Qtey605
tAgaWIeiSGqlRnrz27JXxzanSXkOLLRcWwENXKKWg0f12K/FpJKK08eTH6WtBCTR
sqQ0I7rzOPLebXwns8KKzxfPositSXUZEvTYh/RE8cap9EJJfL69Sxc8N9oTAwPy
+oTJfJ+GEW1x6evIJW4zZ+4bRXpLtrSWifLwp4Qqw5jdIjsQ7l/Y31pfRdiOlFYP
86Mj1+y/iC++7S7dA055cg0U7g3Xqaq1svW+sCO7dYCwhEisme2MyupqHRHlMhQH
kT3WuAeYXR2o8AWVknfFT/aGalr8tIuKlQR40DQmn81lq7qJ2986lQMkcoBJLVdz
JQaqTs1Xp9pj7mIM2lLyo3GHzafLskWs36aHNTTUvzsCsNeBtltfMAGPrVGs+Lz0
ULXRBo2nJAIaamBjGFBz0wffYR25mYzW0Si5DiASDdD8DyITa9NoLcLEyM1L5t4Y
A6tRmHu/SKgGelLXmseq2jUGf9jni5AFzDEXhPj9mapxelzXMhbEylk6L+EFtZ8a
wCmMQwIHS7/pJtsjPPyDpC9P/+gifhbwHpJYQNwSYWHPAyKkrpEuMA2wOu38Wm7o
NfrUPzttzWuXW0EsjbMcc4lpnZjaWq8nev3zbxIS1C12JVtz+g0v3y4heb2x1qMG
9ZcbBLx4XmMKVX2+KgGRG1Bwurb+petXGFmFr1QahHkAvagaqy/tVX4tqHJdZkgw
LKp93ThAsOpU+hdbagWTBjD1Nt7wATWXt596DTjTxUxLe41v18oLm5MRJBXx7p5d
tVxGJqpNHYbfOeujh1I7R3aszuSjzeO7xF4ZcGvNGDbVBLL9OJCQr9NLhCjmClja
yiCB7gQ7AF8PhoMHQHu6VufGbR4ESjdudEV6bwmrgsExeMIpq1J757tQHW8DwmO1
EMWF755f1in3LX9vmBRWpw2WB4ZpqHcLdecpucDOburBGSikI1aosbV2jK2omOJc
FpYuf9RKYFFTbrS2E02L7cX2WyisZCnQWCumbaewjntmddac6hP8kP8+uWtx+Yco
hLWYr923SKPdpg0kFmfYV+0WLdmw0krMFcBuAAfUuZnIxN4JSvv9+sVvIze3vgBr
6EPGWiLe/Tc5SzrT+nTctXpSxHLXQrfWuUccAqjOz/Jvvj3o7poyTSgwLrLfTnmT
HqCIPGtXAQ0fPaCFhbWApbDZe4Gk5k4neaJIvLrsCUQqlVe1gzziourNB7xb2nFc
Z/eqeHV0OP5BH1IZwtQG6Ph8AI5wdXUTaWBj+luPl/idN5rfd9n9nTenwMRYkU8z
cfLcfyFltRIsUNvX8uZRxt2pK6Z5ar/wOEK1rgHjpuUcGxSbQKKS0kp4wPyR2gWl
oGon9JpgKBRg5dqAhTfqOfZuUfy30Wp2E6sb0biRqWwken/8q5y+8i+HFYy4KhJw
pg0tNSjXThjSv8uvEXxzhPA6009zWZ8xiCOofTE1hWn9WnA2zClDS25r2uLHX2Xr
oaDHeQGoWrIRRMBoKYKsjtU4yqrWN8iyInPzzjAZKjcTJP3ScWEue57mqzbLog0O
eqmgQ1wbNLodpI74V7YnjG87w2HCgoID+Mtpnp9pFraMuEjp2vtuj22GKS1+TTu3
ygcV5QFKif4zTWwckaeSGQuCJK46Df5oefEixc4NEbszJ2diIMXAVJzQmDKec3Uj
ageN4TPHfS+0WhZEbGeKOR7ngoVUQLjDdSTAwrFuYfUGvQhWzn5ztsBLUgJwvIXs
tBWReQiyzKfgzP3eN0gR4AfTdwpu2aNZ3FsLEffHaSmm12rrt88PfneXtV59ntud
yO94TtkAh97kPAMxDTS3N3mej5QMZHpaICOD1NCv8XJ2m3PdM5UrMYq66ZBubtif
ODy2WeRmFbB47kWeejBhV8HeXklUB454lPvdjBvG7farAw0e8FfbL8ER1rf4E9li
h2roLDA8k9QC2fkST1Q2A6srhUCDmyUB9M7QPrWYLQrdASjl0RM/X8p5KRwnBS8k
QrbcDvKBXGUDQJx5vhT3WAC+579qLuZTvZfuLyRWJim2l8Iq3fbvPCvCJCKkvRzC
CKuNlvbAWYKrKeKMMxqRcHH0mQveYVBGofXfYJ1xVy2RUs3onpmtiVq9tWfGc8O4
zd56m6zKcyryMhJMlZFO/r+C7L2WCXDOzfYCR4nT59hWsDa+GgiPFVsn9n7pV121
CW8XIpcxTOmBpzR5ITVACUmdy6zYMqIIqhgw+mV6E1gRVn6c8VY1Za3/lNaTfbdv
2ynGKuOnqxedE5u/JgVhJ/HT5iwpju5iDZfbuLcpozZ7lsA87MSOGU81emHdBeLl
TRgFLo0Vnmz3mkmvki+u3iQXUd/CvjJmwb3yNeMrBgGkMmmEg8UoOzH1QJbDlTCL
lkUEmOZWD2cTdYD4RxEr2nrJzOHg9jweCr+AZkaIGjjlZwO6DpPyUAvDY3K/R7/8
c/+VNxzdbwnx/i7e41N0u0bLEsKRXpHp/tldBqgWxopWL0p7VpZ12HVOJMeezFXZ
Xc9oYYt/cAd9rb4disc6fVGcbWPKdL/EMhvBye+3OR7hq3WSElUWqTBvpOYtb0kj
igN8Tw7FxQvKdcttOwS5icaz5XN5Us0vJ0PpKnx/xAUFOBGjhldF6aXW3YFuluxF
WFaZoleXZUtkrjqeHI6hD9XMnT2Wfy55VKlXx8/KohQeESZDCusIi+tvbY2OFadd
tzDgd5b/3Xrj2BarX3rdwZSVTAIZLzr2fDTLaRxAodGFHc7aDcrZ9Qga5BNcY0z0
B7aMAhc8hQI3GM9eFaEfTt2Lza6iSEbgZolmGIE/aWPzFvrl9xdTNSq318B8WkRH
kYFmXzm38McPQs5iua+j2gQt52sioOpUwYed97atXddgTqMGozNJGUlG7hxLcPyU
k0Y3xLP64PpDbW8m46vlvGGycbnwFoIAYnc2uzQWxJTCBU1cyKa0MlGFUTtzRjpa
WJymeSs9QE0Zf2L79XDqQFWLnAF0Q3s7B8aPiFF1llF1LsvNcyVE59ON5DKRSNfV
qUqx4QTEABBTzOK7JBiRx8z7kNvmft+DnFL9p9zaeRwfQZoxKK/nYl/IyrYGsqMc
IRerDACCraxS/MZHB/xCvmVpPho0mLeewOYoGKG3BpaJ2OvFXxhu/12zubD3BfWf
JBTQuN6OgsQ6Elqf2IO90XedhrrXDcuKrXvweLCF95T6Li5XnNVz/bl53iKs3A3X
mSF2tma2xcny7Ibly961iiGSnebj3uqCKnmOK+znhFnhAFzE/MWhQsDiq7MscKiq
PXiVYc3+Cj6s2aeVR5pSOEZln98r6mSNGSaNVLPAHJuQ5P0qoKQkjjkRdFfy5nnK
y5GVCa4+rG6VNPtaYrV90yugvayDAIMVtrscgTYbLCnzMbV8gGqrzUnNNr0OqK56
IGc4/l82K6fM0uqGUJmE7g2f36dWx+YsB3xbx2B8LDZWfnvAiukSPIjscFoXxvLi
czFAeVkVS0ceJXsEarhrsnu1CtM9pxztOkd4oLaq8AKXACIY0dY50WVc9ss6Lszt
rWBL7a5IUxw1lK3FM/2OoqikfjH1W+LagENtJbrkaR7ehF0Jgx5KBJwhztRAWm+K
MRtpJ0tkJnePYj8bI/ZttppJWeJbPaTgwfbT4tbSUVOfH67jrqNR53JnMgo6yUSU
sGmLRfUbDogp/OaKiEVwAsEWJD02XFEEXYopN1lwp5K4pHu4oybPIUbOXElMY6rd
M70pStX6+yDGakk3zrQ82Z60sPWbKDKoe/xS7JkhrFX0p6x8OhnUCAyHWyIt2pzG
5s68XRs+BQP44Ovla2n87TKK9OsBsW6YEByFAJ1TZzzoOe3Gv7HN9yJ7wL01cpVs
u6u8H5tPP0Y+oQovcQltDJEK/GCqRNut64Ond/Nwz7QZGh1qyFCvxDtMYKFHVHYV
ZbKr9lJcxSX5ysL1UcsQaNZxFuUu9Fl+G98hTCUGbljBFkQP+EomnafOTqALWlPu
xJjll74FTfwgqVv07kvB88iX22s9BsWc+2XvnlJPxnrO6BZ1RTGoq1LX2Or70aX3
ld7NuRoN4aFfhZHMXK/PZlJqgcROCXycgSCrpjOSII3aV8W+V8GG5qyoWlaJbqL6
iybl51ziK4hYJv267JJ5YS9MS3YBgAn7lTrJ1cYOQWpI73QmGU4vK5bsAQ+dG8mS
NTHx4H3gb6pzRDV70XJqh0xFwt/TzRQDVkiMezwVrmluhvawRXt6vsZXiwDcFeBI
ZWtPAIO+478LuZ9KRJyJ5Yr3qXS5YgWUuD9wMSNOuNJlx+3+1qxRG0pybYIMrdZr
jpcNKJT/g/WVvXfanboHBmudizajYloqcu3LMOUMPiiFf8MSdp0mli/40tjOuNmt
RtOi6eWtor/0RyBsVEk8QhVzJSkNB/vxZ57fNuEX3GtLgY4j74GwQe8ml18L3CiF
KGLXcOtitMTvT63qLNFYeRRfzxep4N8TqXXZGv9Maxanyc/Fm3hcfRW8p45v7XK0
buvLZGskrhMSYepAxe+4RkoGWnUmIeJIngBAx0gjdsjgARvD/zqge3cPEcL9W/uY
RW0UdlV8lBQFuaGYC15S/OC3bz8AsrE30nfayyPODLZ2DqdJ4WMGALp6sjM4m93c
XMkaemCaH620hbbvfTKT+SygdKEcltNAc/eDz+niO+q8BT8rZIPKrIg+xY+qAele
THh72d7SHB+yyjSHkRvEc6faHQlQjYbb9LdXHp7B+1INsgdMdnoKCHejA1BM9rUK
Unbplbi/esb+c4CDg0ESi06ynEVx1NHVvNSI2gsNR53Z/BrJpBxRc6LOTGV/mVUH
VzQP5Xx9LjFGruQILaMTWX1OPlmqHN2hLeDJhwGSGqBxgLA/F45fO+690v//LhS8
zJFN3vh9lPasqffGvcL8yHN6zsoFlQ8do+9Vv2Mi7Bi8BRVXgz0VRr0EBLFSFotf
q8xb7AoESnKzbNU3cXnfx11WcaTbS+pm59tVYSJCrEeRL8wL7U4YocI0DB07BLR3
SLSScsmU+l+zxxmv7pM404xxaQgefY/C9nmSC4Jr0/GBRLKpIhOkubhaVOpl0vII
oUhxC9zeqgDF/0qG0HLao8o6X6z/hB8V5/weQQYZ6uzwKcxpc8WJ2m92s2Y7SOZ4
1d0/R1KsIDahAjuM0rgxXT0M8YXJ/hSHDBtStDtJJ3SSf33H/oJQeJagpW4qXDes
Ws2MWpTaQJIM4lmBDhf7HH+QHO3vYQUoPGhGTToQizH24einjW6gmRg+dkcubkZo
awDCUH/D/LIEvUVPDsAmWLAC9KrZUnPUchRY4LMCwV2Ui2OTh8Y1EeO3HDGwxh5C
NWZqH0ibFEXda7FEkRdf3sAMQV0pWPZIi+TypVcGLSbfFRhjIb5yGFxgtNF+R8XC
bDgMXy57/zNddJI5Hc0UpJShh5HkmI0fZQvrB2e8cvcfD7s0//x/5HefklxhGvjR
TGaRS9C/BkC4qAEzODrxV5VuHDp/BrHsEwNg7Z8v5UIQfqBE8m461w/pQbtYe13Q
h9L2c5LwepCwcWZSsmcPt3l+zZblvU77y2AQFaIj7MBbbUOT0knB3fBQYYM3H/Iq
MSNnsaUkN3Fl9m2Xgd/EnslldA5DlfQTwRKBu/TmPea0G2XGhPWkqzmtvF+DX5tu
AYOWvawj+gjanQxUTGy1EH3DUPYWJrSQ3aAn/ygbx1L5PF4Iron8ZGuxdC/cVvp7
1nmz8zU4PjNEgbtZThtmErcsD53ceu1OT4gTgU2J2hgIEEdF2CNthP/pqs6JYgqi
C+BOeTkXR5rVjGHYsSPYPamzlnoxKe000Xlnl3QIb5wE+soo16A2gMXSSXugyu+D
WyIFhQEeyFJau0ScaRVgIsJGyMi9fuGFm31t22yZChSC5VoDBZP7MzVw3kiN1/KK
zQAdVjtp56sRK/MSZYyaYLqLswB999FlQE4VzgeQgIGrU6drnKaByOi2MsewQr2w
xSlcJboOjjO8KOFUqZ9WSqAUEsIKrmIexUeTUWfxNY3QtamlHltCxKcaEP/TjLcj
3nq/IbUXW6L2OeJbs+P35Gz7r9wQow5mlKUFv2uvc5zgwNF7a730mKNI+tLGzrRh
yZ6ukpYzlF60QnkIxTTszRZn7PF6f6Pti394MXFsSE3TD3y5yZ3rpZUt3MWeox3l
pnPV5ZpjgkWxn/QUEXZdBly+AeAzltlLTCZwiXMrNVPy/Q+EI96H0Ocd77LPqr+2
ngbB+RZpGluzcHzzSMVXrDzQNIkyYJhPEg/7iIIICP07n8+kTOqmw/J1SDKUpRW7
p7eoBsvlmruFRgfzDMHvCdx+rZB19WDFfKMSoQkADQ6IqVlcmzIa33S/7jtFpA1H
RgLUeLhQNSDZe0vjJgQyCD4vdddeJ+VhEJhk/M1HvSf99QbDZPlZu8lwOy7rsVU9
HkO3pTvhiDXuCigqy/bUqv/YACLdFX5gl2xhJZekBdv7f9OWVBnpL7Au33tPW4F6
RDALS4r79SFxEDFEZVprD3SOvceXf1tHTK9TGBmg3/5rFLDAFAcucreaXm5IatZ1
4ZgU5gDUZ+rq0uGmiweHDbnntrt3PvlXIo7ZBqo+CsMzTEanTVX2OjfxbACcboWF
vauY0qbY7vti87LY1gln5TiXbD15GdI5/2iI8bXz9nCIsJCyrnaQxqM56e/zA2fl
HOPEJ5v9G6QkyTntZRC2S2oAwV7P6slgbpfQOPamYLRQCsyfZH0R91yxq9A7ay3f
JTBhpbunaULn+vmPpjXxOvMy2TAdDnHoEmYww3WrBiyp7FvinkOac4/gyyDviEXu
RL3ffUF4pmCg8cgumr5vXL5jvLBwGCpgXiuRq2I/IeAT4c2B8Sb9bB5iLHPFmCp6
1YuWhppYfgQcz2iDz1OBbDy2pGI4j12ltZ6ZadQwI0d04sf0WXAW3u8cZD5UCH7O
7FXQK9FDk7wZAwe36upsgDrQmzLTXUf6QY5dx7/xpn1FRBR771E5ONFJIO3tLJ2W
Ilft0SocIqVeGY+3Puucv56B3FdqEpxpFgIp1OGCSv35MbOfhJbPs/iC9nyPHNUD
GTknmCiR+DMC0tWcPzTKktRFexlHjRsClUV52PnJDjRtAjH6ASr6dJR0H+jrPRCt
YY6P9yZnI25DBfPsQhIhOmGlyhsDnhZPG+UKdVIIka15xYABdq9Pq28Om3eIyp+Z
sVViRQehGE9arIDAHL3KUkRTgmQxE2Hjhb3H1kzozXsEusgOySwmAktmuKm7FrFb
M+deSB2bOAGOdAlIVSAasMhUbQt9jf+NEDo2J94OkaZopn/5EkRpHbibkyobXbe9
2AoCtsK+4INjqcp4eNHjDIWU0U2yzAcfuAdleSvs1DjQ/NnXLOljhUpzvFG938lk
P1XuPHoG1wkE+Z0JF8hljlktL6ZvxNCXdOZ3Yby/sXCSGC51mPWOr5ta7ooaDasb
ja+iWCVXDQU9aUiJ/pAYv6V+UaF9Qh24QGhAA28R1RLdP0j/W2vuPDaBGv+zsgyq
qq9XxfXlGqUJUMzMs6c4h3K34M46aEGxgK+1Z+PjJx33NaItwv1K7uAFErzLFHEN
cD++tcg+tUo5ndCTRQhS1QEWBLiMQ1v+GLXeobMa12fUf5sZDTxa8NbbF8cozDD2
EaoYJINhiL4p/RO5yoWHxBwBQpHa+zdKTPFjpq42fS/sazixZ48qwa6vzVo1Ob1i
Sqwm4xv/5HBGVqKmBJ7yUiX/aaVSAroC7HEoaFF14O6IJ/nhYFbrY+ZJpwRo9wnY
AV4WS1hf7Amcn7MvqJeV/nMtsZhwhgPPiKM4EPAg/U0c25yv2aNwrC4T6LjYVP/4
5+NyA8ISrPYifPAlKkcsvwwdgVdMLqMmfeDLSeNAzn+maxEXqPvrHgaA5WsUH3rq
ld8KwVX5bC4c42DRn2UoUuYTJA3TcfSEJObjUvLCyvjeNwt5+TzISHeezAVexTJ6
mdBbJ/+qzfH38rccFO8PdIeT+xVrdQtA1NE3sP7yyO1kz1YwIIk64g/qSAWgWf+o
d8b1T1i/t5GE6344ni892btcbEB6J2Hua2O6Z28IiHI2FkMFydF6avE4g0mRFZXe
c5nH21hgBOuMN0wHgJGUR/TWZtG1LgzKnCFGRQOb7T15/HyoG99HNei5BUxvA9TC
XZPbrLuafk66XJr7RGVFqWBKqitGtfNBWnIyeRxYUV0+TDQdpx9Lik3OPp6tIUoR
WESkmCjQT1a1aCtyjAftWxu52aAbaTvLLuwbMBy6+UaufyEiP0MXAuZSlE8/qcW0
WXWMhxTu4QSMvvxCS71mdLjH65ibuXDZ78RgvtjePG2uGecVsbtEWX96MswXnHuy
RIvc0qlBz0WvpqsOEUdDg1uhXrb/TRZJcmBtckqmvIPTLybMHBHE2Sz409j251HP
IspwVsp17G8z1z1XSPn9AQilSX3z1NMnGBgU1meKf4gdIbkqi1HcKPgFKyjIqkOh
CC9CcoqfYM09vhTIIbQtpGaR5nfoNY9ioOppCLUtOfAQjgG2sdMPo5fy5M3aVtlb
jY4ft4BdXBBg9LF1zUggxt3n+HNbnKLuW1wr2p8gsA4xaGtZQSlY6tWjF2GDGYrU
41pRtkyaySaUmu8NNTULhS53zbRedhTKDSgfgqiTmwiONW12YxGkutJyh1n9lfK2
EPMyBXNYCH3OiwHul2bYEtRSvlA8LClu8cNmvM/fCRO+7U4PrJqhmkV9dvWb/3TV
Tti+eSZgtOwp5uCOAO6mxqHhp6xUEXu2ckY+WyKyS0Vbnyavvt28IKxgjC+eoDgr
3gl9R6lcm+mHL02rp7G6HOlQDjdsQ5iaE5noeHS028IsQ6oSlY/UW1mt2uomqsPC
sMcz+UCSzqUvMzVZ2Y0343wrbRuEznrNwrgZJmhUhNe2P+T5mQc9dL+1peObRwv4
CrkgzxQbvx/SMapFxPaad7jaii5Z5SGADWbshaVE2Ku7br5Msned8NeWh9NqpSiT
4RL6SNmTB/PIcyw/eJoHo2vKZFGwpAKZOnQ5QqAI1fBbF8EHBCcJOmEDpDX2NuaH
YMfkuON8ogO5TI16gtXknT3eHNr5GFQ1MTRI6f0ZHVOcFNOk9Z4hHqTAdHnBIGZp
zlJA4WxJ+GQDiw8O8Cg4ncKKPxfM5mohCz8KR0wBKvunoCoRoe0qRVm/CO+szuT7
/TH68yxnxNkC/KdjC65jGZ4Ir6JFWT0GvUfFRw/aH4BGAtLmgThYHP/pr3tsGDX+
f6zQcqaoc4goR1pDKBAtvYggZrtdZv4xk8VYxAAv7qB1nVmQJhZhWhYEXWuIe2Yx
tlgPlbOrhRhfYwcDTZ+ThqV12UDgIOgeatWmrmVm8ir+5TvChMKl3VT6xeGDfmq6
qyVfB+zLiNxvpIIfbjlXCMg+4DbFsvCfmGzetwtilJDvwbPnPw+n0hT8xZu+wgkJ
we91cDhG628ArFA0zHsC8ZP9TltN6i0/cqZcXL0i/8x/wsYKZzcwDG3Q/nfn2uMK
CKraHK6rXt62MDa+LGU8+vJ48L0HkZhflbOXkkxV0vIcXsWlCds1aK3qbKNmPUOW
50NIMayC5HvNxLqEuMAiUo/L6HbcHxbd1EEuOz2a5dxYI6dFhCztMwx6Ff6DqKFZ
c2aNVsOKL33re5fe/wAz6HILRE8kWHUbfCx5kzguII5WB/dR9QgxK2gicey6rwpZ
i6IACA7+z/R2BHvUePvIA5MjPRO2Fb4S2DKHPV4PCs08N8amGSbcZaKv91wzwvQe
GHw+yGJm1H2XFVkDFHtwmsW0XdWXWxZTLoS90lcqXdokCfOw8ABMnV7ODCL6YqU0
oQYnRqwAus2UD6oxkvG1XD0xSb1sa+/Q1jHg9VYt13OiFmQsVOSlBY+4OBM3V61c
QFhzy8Ph61pQeTuDE6LaysPERbOnj0S0krPxwP1Ub/x9D9uSn3Prr/GD8QvDWH+7
mzsGO1ketRR1q9ZikjLHmiHpHQHl6fdK6OkgpWNY/CMSuNSFc0+z+e+O44UyvNXx
a3ZQLTRVi2SpL0qbppniR7ySIrlkO/sUXAcfS/YqxN8DcstDAAQBQo2F87+GtjjG
VjU30sSVgSFm4bxbKo9z8twuCaHfdio/wkpenjDkxmE8is6TEawE4zoaifXACsIq
0ZZmD8vdm6CR2o++4a8QABTbzDFlK4bhl7WkfZXjh7bNzkISCOpg5Whz0GUJQjsw
xsgH6W3ovbno65+cxARxbQRAuLzIyG465KOyde3CCTfwWlcEYpEt6w5qW41l2AFy
zkUftYWfcb893PJkwYudP3sqxUYxth8PAiTQtIXTBtHko5O/48Fhiq2hDVPF42JK
p7o83gfk9hHF1Lon8L83cSxm8O+YBR3uYb7DfjMGhEvaPa2mIOytOGyCrn5sAMhV
CcO975BTHLm3Kmez8GuOnJZvLS26RzJVMlAmEQjvqjNcLakBo5mQZcS9wSz1nu4S
f1/NnDK1Gq0d1wPutrZuMkrlVz4hKthJzMQwoVisao7Wlm8JV1EejxiKW3FPoMkZ
wpfRAzH6TjwJhPFWZ8OCqRs8VMVWKmeavjkUH8o87V1RN2LsLyWIHIA0hEVIMmAY
k9Q5Pp0g21kP1gw567tHO9wTymJdhfTIuz1vPiewBdUKcopTzoPRorCdnE8oCTI6
xWDmCJzT3UmCu3gNkeputE7jHqoFtVCKNFdhHJ9fWMdEMSsjX6Lzky7aQsOXcyxK
1vzp3znmeyt2RrPEyziTyrPwWqHzTVXo5bdM8i462cAjCSdmK1G1PY8r3J2G6uKF
T3WKCcgpa/hUKKcK9VpWQifDB2nrcFCO7q6KPum0Vucvf9CNwB9+dQ4mKUhYtfZQ
QeLC/nww5Mp0U9JW532VjqNQN0cpgj429X0P2QTMJ0IaHkTj8HPzGqWHDzl7o3Ej
lsjE32cWkgq2f99xP8AIHhm3TXh1gQ7N+acDBWorXJhCkulqjTg0Bzk7/Af//jgY
W6t00kOJ1/LUnXWkr8gLQ7ZP6tvzNeRUX2ZznPRkVSVM17xmBMueTADvX4p+Yd0U
/t6Mi+7xSzaYXwSqZmGJODBv5+Ze9CcNbtBQnQ5yCFRj/beBj7AuCmysJ1tTBcNT
b3swbGZ+92LRB+dWsk0j1kVAGBF4z1jpfSdadYUQTFXC8CHdroV5HNEXIH7kAhaa
I2HEKVT5HYhMc0njhMrqwpeSglPloU3wpWXyA/sONkuYa3VaHOCy78tls2EvrHjX
xDdeCmbnCGq1hmA8y2zCyw7uafkv39Rj1VHo9xUcfY7HfHQyqZMt3aMwB7Ghi8G/
p8yoshsz6G7jH4rciW1CQOy91CY90LrYAkHazmmAv5ndrclOz8M8Y9QtSzmtuChA
z/I28q6OSqvuqRhPDB/FiNu5343jTr1MiGP3pN3Hj3jI9PKlnLwnuCf0k12kCz2U
9R/i8wLtJVCTt0G+CD+0LMY0BgfLdUsoetaRphwHBxQep4Th+k1+VhKfs5YTC20C
YTJCRPHmEpJ0C4IZhm/Q2eTSafyMsrmfXy8uKHAxYMN7vF8njIEZzhaySbv/kxtP
TFafhS+C0tTsFWDHEO5gS1HfK9XzI3OZXRQDi6c3EIPXhyOzSsfawJ86/pM9syba
23gytcX+BELobZq69Tqh/ugR6dUffIzRrH40+qcYRee8LfQzfXvVRx+wj23wJqgy
jj7f/H3XDmj5mX3fSArJ0F3clRIUk2VmQcqizVyq4GJ4lu4sP13I+mq/16nRVW3e
lkRKtdAeRKzdkSoVGTOFISheW84xk5Pd1pmpfj6eKNWfu2Zw3L3aC8di/smw3cis
LgC2MkDnSQxB/uXSGS5RqPxjpY9uuJzeWSClR0ClIHOWGf+voG+a/o+8kuyEbsyD
c5yzwIWBhMNMet7zjvVUX4PgLzwo62tup0JGWkwdHixmmMwYyYBsWaYzOPQW8Nog
d1Cui6YJLQpY9As98SgK681kXGxZvmGtc6LWDyr6PenQ8c4UBfzNEq6DImN2FN5M
tM4kfW0XH2RRFyvGIgmrf5fmDIAp/cR84jfnL66CRerR2nUhFVJweBkoEruY9t59
/B/2AAvXIQrYXJhu2vGsqEQIf/qgZVrmP5u4w5ihoiUInqitJz6Id9DYe1wpdYIp
LdrSB34hfP8Ovoj2o31VY5s7BpZL/57jrrcm5//RZ7LKQFqHeNAK5NR6iOgErhc6
H/ttxv9d/7QjX2T/f6MYYViOf/3SH91R2W9pVAcO2U/hY6SCT6E1rD0SrNSHAnM5
/nxBouAU4c0Kw6PCYVWG/aWkSyiGISAfgweu60IpuhE8vK7N0UXCcCCmdlHKGxdr
/4Es/RG25usTBWRCRzLTaxu1Aa6220jwt6ARAf6rF7aAjpJyujf257Ufc/8DaPQ1
sW2Rlb3S8v2khtYq014K3jsKzIxS2WoerBj3/TLcM6Z5BrGRxmwDokyIoM/Ot2PU
FPnGABb6p6VHU5ytJ2TKWz8+92hxA3+wEAHpJDZqsIjKK6pJ7923NN+QvuCb+I3f
y6y6RRf+WDgfW+D3dLWVwTz1RYg5e+RD6HIH573ZaIph5ftIuPAkw5MWa2vFoihm
iJaRWTvw4vkDS75ft1oCTSiig1mEyZIu1fytcTJKm9OLDqRwSiMzm1krGm21kfrW
dVYvMqOiZsRR1i96PUwdSCanCwyDgJ0Bscls3xF16Z8AIXkOONlmyK3gE2VT8fsw
drhvwH8VTSnBuxiOUf+aS9OSbUdO+ljsBW/ewx3WolPfqV6zFjHgX5aJpTMeK29O
wvUwCb9epxVj1XinAjR64IzGJ3U5bokcXi5jiH1u4EsOpG/RrDfgHJ6GYfm5fIzj
3R/rYYVWPMtZvCcM1aoVpRxfP83InBr5FLC4Mqy/wZkOZG+12xeFSYcr7pbI/IUx
nIq0Jl7yEPlQjwaqyXwO5ko7bDeFpn8afzpv1CB/2pKVeoPLisYYOuCtqpT7lWsC
6hLaSR8WV1ZDckijrD5H8y5yZuy4PlDB8asoYyD+0BvEN84Eh59+b1xEADS6D4Cv
7L5UcfFsN0BMviDxya+cm4eebewG/P5Jpk9PgyNeaO7shO7XAqfg2beS6Hxtukcv
pLysTa8y5d1bOSx6Qa0crAQPouJK8o3jXT/s/w9KYSDubxAjNNEwVqpcL9+xhABk
0SzCDRSEQTiggGzNQUyzT927onRhjEdp7XBIWrsh6BiDW4FvtXF52WsIDFxqfOWa
wQI8FCLBU2+JAJ0DirdROvea2eg0G6fIIBk3tHAN73AOK7/qCaRWSc3p4lr3bgy7
xoVj18EmhjUepGZyf1MgClO8abPKBJRNpzYptvg4cpCA44O3ISKSaUGm67sP1cuV
dQ5vcI0+v7erMb8utK6YG3EIDN2MqD8PqNa+4MxyuP4r/CAiyJ8310h1wI3Z9ets
D5h6SgwTyTNsEK8f4zSPzAuX5EVzCQmAI2/rF3bZE1K0HLYxX3YeM+7kB+ruCDu0
fq5U8lT1g4cAWr9EnQkKU+RksgFc/aKfYjKLpxDmaYU4KAJGVkoUfdI1tyal41gF
ErVNp8QxvxSVztIF1jt2NyhNjKFYbGfgIrSLF+NAchp1+BaoSvr7BNkHlextM4f2
INL49glRHwZ4IlUttGTg/etvJGXUm/SLxkx2S1Iv2cNpbIf59pXIXWLJaBgJCnBQ
RQvwzy7Xu5p8JAaq8o750aniAIQTfDRp9n1WgKA3cCmSqccC/MeVbO8UhpeF6xtn
2lwCG5EstSf7Es9DJddQH4lwNWfk9AOY9M2Iv2758xdAooNyk4Se6ro/4lFVKfGn
I8hJoS5oHw0I3UyvWSxZDSZ0UFGJ2C7M/r9H7iKTSnbmh16aZZ1hBQ9Gt4Cshmcu
jm85pQW1CKumxKQaAWCq61ZUkba5gB9v2XAsNmmvoeGXUjRiJJ4RA0egt4wp2M8y
pBXb5rCtA50iMHwbJqdSWGAKV9pWdirfg8m2Z4J8fjbabht6OApNgQ9PsSR9iKKT
Nm9Fvel+flvb4C06vgja8KFP5F4iLMhJgwXIDchFEvfr5tuGrTstL9D3ozYa//I6
9ABPsvCF2UxTOx5FXwwY2a5AZ+L+QEMXYzK9PUZuFc0FzKsrKK8tVFRTYIrLuxA0
6K8LF1awvN6OTHpyFfD+7MshMCE5vD/hFduIHNNL0VFNzqTEQ3IZ1ZqEN++Bj0bX
ayXAZ/zTCjnNgO9acFlzZvUldSkKvwECxyPLefBYHwR/xq08VdqgIjWwfV7ZBBxb
HSTGJr0LnadROHev+Wi2aPS7ufVQ7oBHSv90hkZGHbbYd3XEyPA0gJ8WOYHtRqis
9wKdfpUCwznrxuC/pJAp13WuAHDpPcYwMX+mrDLl4ts8yEETc+ZsYl3QtcT32/Jr
GkmYNZm9ilEWvdBucAJLQ+1b+6l7+HauZckdY3ESiLzjLe1CGlhJ5jA0xyIFbJ4N
aMHH/XpGJ6yK8YuLFXc5URNzob5mUf4Iw2jb5jdPrM598TMwIaajESq8B5UvUV+i
/aHOx9dprq+hAn4ot349BAF6YX+yqtA+JgxpCIWH/c81kL7efBfd24+Tm/T108qr
R9Ee6J0nh7mRV4CbJiIb5WkGVFOEEqDjOxIpOe+juF03qQyMkCRLt+lPBzNaojyA
VuHVxmGWprLRoieIS5f0SwwMlVi/guPXQ0DrjQ2d4GvVSmFg1hjo2SZ0A7rbWFUZ
0HgalrJ+MgWJeodkFP4e1b3bDD2sAwHvC6Gx00B/6yxEi+E3ajBFyLgfsBWwrn9a
Nv/6PUxkcSM9Il5Awh8dGlzzZnNC+KVCLnRYmlywOKnOzBIn9rncNbdwUEaqCU5C
ETv/QRysErhr8AuyGxkag8k3qMYd+NQr6BCTq6SAFn1IAlx+40Zhaunl9bKdKBlh
ZXVi5rq/6dlufzkXz6rDVpBaMGbA4XAHYVK+XJmCrqjYhgO8i8AgsAJo+iggUv3j
j1fhrAE4brIj/BcYgEuB+uNF+2gxS+K6M/HV5UK62bIIeldRwIMN2fZBaDaMmE9C
r+mBhKFln8sEFdETrjC15ygu8P9PdlXviQWlaaCLtOs1YpczALqihyIxEbLqYSjv
7hPmYyKheTXuUvRwgDJuKdWAYdq7/U9Hc0aIOcWbz+VFlOZH+BnlIaSMOJtUqDID
Ms/mO0XWhSi1Hgi8+PsS8g6L4rSS5xzrdrzCbLRqkhKN8TIWr0txEzQon20W44TR
0XCj6DZ2r1fkqOQ7niqAsDvz/RuR/K/t8Y7vNbyJE91kAjqoYDjUAObPJlHsJAPO
XR1UNzB/kt6dPfp9eF2bFgJY8fssEYDwOEEJfgwWdwzYwQkMkN/Xwp34XjmN1GpI
rnKLSoqTM5WWpj5l+7JK3AH0zYWWZTCu7RMQWc3EUdU8ovueTsY/eO9UpXPVTNgR
EofYSJ0gn2dhytIMq+KvuRc75KAhC9YlID3SlLPhGupsdsj39mLL4T+9lYy4SLug
OKoLaFLuY6SqhKNoHqDjoG5vbuPYkduE2+u6z5Fsd97MbR4wGDOcpozPzEACtyKx
hTrlktvxC7va0bizzJ4f1WMPDECC5aoUbu70nw84UOIPpr4onXunWV68CMvtPCFH
dQUhMI8GRUi5qC6FAncfKcbjM9oedtKnKAN/Qms2OPdmpw/WMN/tOxX1KAGcqt3M
jvUew3Ztwf5ZSlIlJHE2didHXMeMa4IotbrROT81FvgoTKXNahnc4rUrC88nx4JX
KUpdFSIc8MroCytoTPVdA/8HM8jbKkuI2/xDWRB6oOiK+HuwfSY7+hVRJzYqKkRz
BlLrEkIRJ578/6I74m+jUMKy0R0F7kTYL3N5ICOu6zi3Y8Jw2wpCOB49iOA6moqZ
7iiN3ztGgiT+envV9H3SqcqMuX0KYs8K3BkA57r+uQt476tMK7WEIAv19MhwrdA1
/R3D66Bl9KqJFm9hZ5ULYUbxoLlMZTY+LFIFTKmPaxA0DFTAxEY8N8HxVgXxoR2Y
q6VGu7mcHjYoYfm+UGDQq3bQHrsJhR6EA8XLU1GfGxhjG21hB64Sizt72xA/S64F
DhYnOE0Mki025VqEEdU1owCkp04ktYmTRQHqa5N+SRGQrnJuSgcQBCs4J6Xe/9bp
+JpQ/XHMTBLDC9AYl3t3e26xRPJ2fXKYOiuEOGaDEGJpj+8iEmZ5if+SYJGkrCHk
zcCgxlig2YJ/JJys2LUthfzRN6830rbK5FRxuCte3LkR18WGrqOEtKh3H5qHnwYN
qjbux1Ac/DY+m8n8MQGDsuVKmx82VfrgcpdbNxbddeCkaKRC4cNjQoFav16BAOSl
hOKCzqt7+REWQrIJtLce/QAv9FpJMJOcsVfqHiG8DddExi9rEJ09ewhBqpquSLef
pRCUVnE/lKQtlKKPZWpQH7SiofwgvXF7TAJTl3W/qRBKjkAPRI1HVE+2WcgbDiFD
ryzu4yJ12ewuay5bm5SPxvtrSJcDBDKCEHDtBnLqrhPqqC6ROz18X0VyNVwaXpAN
s2up+XrmfGryAv11pT5vZ/gtUPwMQoNLRjiLYYmr58Oq0yjrKf56YgJpfSREYr7I
erVfhuRCWTN/vU52KS5uGckQIB3zAQNLFw9cc7I2PHFW6EWopXOkRk8t6W88fzRq
ioBiRXbcg4LRrMFJSaB526wmI7kb7D61CpB+O9lqBamvA/n06vGHJcyMYjTaNHma
u+ZKEqlVlcM1myJL47AY4jrbeg0H19g5rNyWzPjKMgNaKwPTBG4IpA2lN18ZP2/M
XkCtnzdhhyQEktXC1VIYE/BAw3HEdOW1YMsPz1kHoyJ6F/SfINjqJYkuoDzTGcLf
9J8fpJUjewUbWbNjk+FzoT5AfX8d+2HkOfFG8ryL/0YeJbMkqgoCKVxU8mDUSXg2
qm4bXkekIuTK0wcWWuRoJVJdUR0wJ7S/rvOIcsBCJyE5alfqQBLTXUkC2JhyCwRN
T90JdDlz6pnhJ6g23ozYKNPDiMfe0RT5NdlTt1u8VrEuwlWeAQF/AFU/SboEChSx
ML7lMZEeSJJsq8qNoNXKe1OM9Ze36mE9ZFcPwKdB4e9QFOzwtlvZV28MgFEf8PUW
qZPwDzjS6TT14x8Tje0HAiSyzdeJdGFD7ugMEdVZclUksyYddB0nCMxmeHXG+Kg2
dvQhd35DLwG52ZeKXLiVcITidYrJ9jPhcaBu53a5+upD/RZ9ZeAimnbtb24wuytA
Sqw5fGTEU2GiIsuX3yUSab04hwzVYydIfyw21G6yBJ+HB+K7pPI8/njXqh/BY9+J
tcfgcj4uga2zAMvDV3gGuw10rlKGIxgEyFx7jqFiMFXUEr33dsEFmZ20SzUyhf5W
+RA9h69u9jdw6E9PJMna6gXWT1t+adwZBUUDgYbB3kQl81cXVyOdK1QB9uI7aX6m
Z9nNPfLiQskXSAzUJO53nR1G9xVsphzSn3q4MHzzykJp1QLasxHTVhmB7XSMFN36
LRKa/u3biv/U6Py1S4MfQWFyRHj+7bOeZ2xgfHweq+bfdLPXXNO+42tf0A/twvxy
iB166ggt/6bSxxvj/HZOUJQH1pkvsa64Mp1NL27fsp+9EoQ3K6XhfSByesrHboP1
/9Qf/vrZjSt9DSVwFhgUw2jD0gamry3fLArbzqmJrPcQZHHn9RCUQOXcIEhjYWKS
FgNo5v9iQvbjl89+bhs4knTMxO8GbIZ5qNMF6UN639lW+woxoBwHrejyflk7GpT6
8TGWlTIbU75XYDYXBNOJzHwJr34MYdkiteK0fWt8Wg+oTR16dye/10BwoRQbZ+OZ
vPrqAXAm6U9WlO6WsUBACG/g1ZU/1L8OyAhLaMhfO5uOUAuC5yWL4LQCvdaoPNHM
+PGx2LmtsYQUpJJSVTI7+M6JgzZk6NE4K1zzbyIDe1a/QXf8gcKf3T8msPe16ds1
wq/JM8epJ5HVCdFIopQoHHiyCsI7R7FEtDoOvvybwzw/5VveLADXgBCUOBon3Cv9
OARD/BGG97tkcAR6XL/o+XuJsHAXv4GV7MH2LlKqKKH2hKSEx/RFwv1ycwOT9onq
SpSD36CojhrjUT/ZXT3fzZZDM8r3X0X8d49VrWa2sS0tXQD0ZHDLBoYfwAL8H2FS
fyihKhUKWEGJ9NIN2VRzWxGcGarIzzZAYrc05kIFvdyGU7608OtMz8q4Um1kLGMb
vb9EPSUaQnVs4APsgrs20bfvys1BcU5JV66qbP5S0NsYpg3oOsXgvYVLLe3PWXxe
OtX9J8FnTLEFRgieKklwzBKBYRMb7k2HOX/0puebJiUFlEEdbalEkgEDHwweIvwl
5Q24lf9Oc6t6rRcD/b9KzplCphvKhMqdycKsy3IaFN/Tj1Wa9sZPGV+Mg+CGVufZ
ZGPLEA5iQ6CDjdiYnbj2z+p1IUVfHuJB5HlzsdaR8FXtE6zB8Dyjs6jCF4WSm52d
xqaf8MtcS3Uy/GZfP4aNnfSZhHX4jSoNAg+8Q4n1/NaqKcfFSMSyMOfTuCUFo9mn
VNA59jLyCZdOTikdxf60p2lH/lX/YwCbSnWJdWyRZWvUhmE5RnBQbFaQvCuB1dPi
iq3ft+uiC99sBJG8+mMFpkAqlfXI6oczKC3i4/VZfg4gaYqmL/a0xUIrkymsJGUf
pcSdT3LBP8VVYdGDBJJh/8B8pnpb8VhFIg321RRlkWNTd/SdaD860GBjSkDbGuHR
DBOBD3Rxnklmae5O1aE6OJYrJQVcPkrhNK8yAG/ru80fP/oh+uunLRpuUbj5UHe/
+iXaRsAhkRRM8fCiC9BL2ug2gNUrkFkfvLPvLxslsNv4POAhDL2ETemVv5qxJPYP
FdduMIw/5e57XnLG0NjoQKFEWbnqICv7KckHA7HVQPmcfTLuKShFvQ4ghWIsG89b
UeFjxQ5LKPyMr3SeOPHSKN0SA8IU6FhzwbXCTfHOfk3OvsxZ7CdQjU0aTyQSRwcd
UmpIFvAS65QhaOpFJsZoKLJwRdxhnXJtiyHjwouX8mQhwpoIrljh603GL7e/GoU6
EeIGnCdnxEWUyLKeNeGKlhz6eyMmvTLp0lPizH/k6vYmHYnbNUPiOphBWbKbY5ja
u1a13z0470fLMLS4xLgQ3aHDAjen3HNGoMsNXETT+srF51/I8KJHcArqKsPKhk0v
21bzG2YE5QdhzFujsnVXamcpQTL+IPSMR6iNX38mksu3jhL0ueZQsSVKz3/IixEx
etGoSoODvVTEQ//NEd/J4KDonTcmil7EXlFo2ryX4sU3FNrldilmi3kapiu/M2eZ
BsGhj4xbBLm0Zj3HWbUHjJ9P77ny4unq6m6hIVt/tH4DIX1BcXQVmfWed0g1GRJ+
VL/EdhKC2GjBUE+H1NcjaKSBT8bnllljGGw7SYtsQTr6VTDN/oAoZMu7+ulvJqvH
5zvRnxBUzxgJI0qgYFnym4K+mMNOtT+9n9Cch2SyquvNMBlXWLrvvHmT6+QELSlt
Xd6RkUSy8If5T9hPe4qoRtd8qk9e/U1A5e4mALACI5mQXh3qL080JFYao9LHBcWC
TyVTVC/9HscJ5v+q6JbFiWqBttUOvumLUdE0KkmJzYw4M0eS2r0gSEivwuuwMyWy
bCkTwYrCW0X13HhVsDv3g4udQCJySB9FE24gcEugakzJHrCr1kwYMEx+kAMiLsP+
tZwa1670009akdccl/tx6dmgjQyN0SnwcXam2cbaXQBVRGE/7yJHZJIznOp/jpxW
VleUfWL1q5VPGS4sXJDb43EoNG+Aj+yiJxzJI9Wy9Hcg+msZ3h/k1YTWJOhA7Yym
3Kv5q9j3HSjX6OVxHFkrzRcSi7QAeby7ct9HiNCJ8D0Ak+2Ig2Ar1w9+dBs/jia1
1MR2Y9BPxd6658WhzF1uoFm/HZgNv4CM/QuQnaixz49Nk/MGkeynozijiqEbKior
3SPOAUjoE2VQTFt8OZOTMwzsFr9X4oP1QrBCBs+JN2CeD6C9GL1KKQjYZkEXsKFP
X+xJ+xmr03GfSI0wrzQVyWksulJZ+yuH4zJ3Gf+SofF+DIz7b1axUlNULYkt1t9j
+4l8TaX1IOUJMhu1XJz6oy7Y6EIWucvmazOOThIHBZB/LjTjUfbmMbvd2x6YYC1I
BBhGl24eGuPIaLOoTnDTwAaRfQ7nFzKUXjQBZ2wFgajPEJv8oTNFYfcVeUo8vNHO
DYh0AVPmIZWK1cV/Owi3NtCnIQXhjl3b8cmBDAJah3Vbl6CbOEv2qPdGSnL2xrus
JZJbFZUE3zw/OZDmO9zSS7Hn9X8qk3I1u47hCgcTDOWny6nBXT/7ByxUvwrjIO0E
HS28gGhfCV132Y4zh3wCoasI/hMxR+sOdx9CuUmVci9kpngR1xBz5Lom86RNbThf
rtULdJtWMgM9cPGCkxEIqhej91XyTq78jTTx8hLlOD1yDrRA8opYJlzwT6m5YQJL
z6C+vfnvfdxW7CuLC5usdXgkjhl0D/f5RAgpRXYWAi1lFO1oHwW+w4PARVOisK4o
HrrNUZQyCQfn0rcWr3FEdZBkd8ygVZaMTshAXmqEnMjqD3hpx1hOS9KS1YtWQyyh
EG6Ygf+m/cTfk93ljrHvzXfeTeAT06NO+I/UtFbHpjdOKerpCna3X5eOtQD/cICN
phHcJ/ktkWnv2muEkAumfX+tUdLDYj9AVHQhLvd8HxCJHvcVw/Wwg1ml3lHgkvGi
qK5gQ2NASnVOjheeNF4c/DG8aN/p71Ghn5/+6pvfatSDUgQzM7DJg7eqDw5rPMMf
FDYTrayytT9UgqanRuNRu4t/P57/2qaXi50n+QLoqvZv7RlvdWkCi9HyC8ig8gpX
oGp9mVKH1s/A5bRTvf0rYMSSXUSZ5odalVpuwrGaoCzSMEN3r2dFqgAg5OzJ7gA4
ELP9oIZ19m+OAPTBipbYB+QFhouFZrY6QRXjXzMU8TfJ3Al2mKcHU9TLIbr2Y22/
hdzb0QpPsjTZBZXg+gWWQpPcVyvKNXCiaA0kIqjywvA+KZPjQTyW0dt/zS4P92Yf
afauy+H0SoCt/0Bu3GtveywfHBQWkwvT61Y3GnM6WddYmAnzIgGfoZxrKM7mwS0H
XIKuBqWq7VjP4VHdmVtEmNnTGUX6gXw5Tt/q4R8Ippj9OpiBjhJ89iu9K3pybxUB
zHlVSZGOYI9jHg3UbipfCgTClqvqje8hzcsGctwTAn3lB5Is7fxuEieKmSaVRTqm
73hLUQEFNHIEEe6eZJcByoTSvIQXiajW/L0dGmFORTZNDoujHGoBEnshIfsT8TUO
CDZDd9Xj5EkYX/THaB0GVLsxumTja0LlEQac11cDBFLAnc964L2uoEnUDRqd60oH
Ubfm/hzCluTxK/zdIuHnBHEf1NkC4snK0KdZlHCw00ngso8SSTbGWoKwG4Gtptjw
nVWyVMo1esOXSc8Gqje2gBA5+tSDH29OZQzHBfJJKwHtn03VYBmKKQ4gnyxyVJVB
gj12E+jK+kibat/sz0wwpwf2jKSiZhmM5kVoKK0lrDFJgPKVKQTZsVcwEh/GmDbA
cfzcu46NKEoyVcs9Qrxo1UsOlsXjubAnyeQwqscyBVKCg4/pvDLEo/OBxLzWvgX6
Dj6O2Am0Ua/wfX5yrFDlgvyhZ4yseCmZ/JldDP/7JuGYitxyDMHa2BFwyG7a2vWR
uNa60tG6pcgzwuAUpHH13CM1lXrLyPhA/dBlvNw33sCRfIcF8hXn5kpZDTePV+d2
Go07e2N7SxHNnZFsb5lB6R5hplJ+Giwj9JU2sN9IpVczs1Yp0vBkbL6Bw+Sy+afl
S+0pBK2WN6Pj8J/SwgwIChLr5WL5nQ2BrMpwi9Odj7tPpwQ8ujYAFiJK3U+LSaN6
i9GHPLkzRYdmFz09Vt/PYYWRZ4AlrPF6wpYapi0bR0U53IayowfGvYwKTxDQX27b
3lVMe/0lJ0Y/azIlM+QrcrNatZGxCwhahKTvLs+uAKsP1SMtuqM/JtUeXmbLJfcZ
VKVWaRsfSSrMmnLQgz1IBwmn1Q+uXabsKkYCuLYOAeUB6EVWYXmO7QBRn+uTlePr
3u6n5xduJgEDYDcixQ1FO5BFrSbSBxKAl8EyVJ5AlyIbhATEnef0D3+5nNVUk9Oa
jEZ9Ie3UFxdjeAtyrAnP5fvnHtPZ0Vc81jxv2AnoLefXCD+UKDlCEuVSVmfdam2n
oZutEJoHjRMxfdP2Zuu4wy7HiDGBVdGS49lA9a1nbfOn/bhWTOazjVTPHJBGs72E
O2fq07/L90TO3zhPR2bCPxnh52MM8Mb+lAaQ2/AMqtR53/oGtOcGe3au805QvNzw
31ZNgWw79Yo3jnStCh7+sI18bAKOqQ8VMrLgI1/la+vT2hv1D3xezWeQ/fLF9AuX
q41p09jzN2Mxk5pfCeHkPeNZG7QBwTkvCZVvgQOg/hR7vWcmUoxqbrbzAyKtxIO8
v0IzIUptNIYWqTCZasi9daggflwAH8svR+Ww56Vu6vH0LJV1nxc3Ie8xYNs1I4a+
lDLhddfHhFo2ZzJBpSb04xsjZYRq/nSLDvEdSExBgQTI24WpCGKINXFhjxQ9qyDr
B7UvKgAOsO1lEtaSdezTCC0IfEBmp40D6zJ9Vc4r4suS07JgLkKsdB5TfPfsugMu
MWWsiMDJdubGhyJomeT7f7Qrb9uv+/WXODfrhDiJNQe8p1iIfzYGOES7K6fwfTz3
aO6I2rgXu/faALXViIZJYHcLzgk17dif/P/7nU7Dn03XzDwShCmWEwzClIxUZJLQ
zObLVxpfl/7WXWIwGaCTt5n/+gZFB5deCkz8oCGMA78271TVxqOQ+T1Xh3qSmy/0
FfhPgfCyKea3tRPkMUuKfz8cB6VrbkF6wKf0gbptLpmEFXClkdaaoHfH6e3yVZVw
zgH+8/s/LD8ZTPvhfX18jSAUpAICnJPfFzRmgVfkOriZJBixTa7lbNnlqojzpI3r
J4PQ2aGHhTac9+mQ7s372FDJ3fXGDsdsIGI74O3ihhLlhQKuOV9SQ16CfR82y2w0
0tb2Wu0D155EiCe8SR7amsbJyLqiJB55GKtIlIw7uQMoVWobH2E9ikMTdj2ftnCu
s9zK+XXfgM62MFPaMM4lSa0IUQLbSBS6oVWXW/IRKezdBBQk6r2uVbYOKQulg38Y
gF7XAE+sGj0q/jxsCbfS4Bh0imBjSxsI5iFp0SAWSj1wi6r+3vh6m3/cuzW0Xjy3
CU/kYirSYKsvcmA62JWhXIztFgYCHZnRosLJTCKm1x3JIb924mB7Gb0Y26dhawsP
PZk3c7mlstu42m5Ch/OrnKereA0at4ksIXSK0MMQfAlIUF8Vum73l/gf59BKDmwz
wpNcPZfT5zHbNwqO/vhBln9eWz12SwA3hMtgUsk7kOavBIFAqU0ImvXfW8/hDYW8
2+za1GQYJmSRVG4hAW2GwX+7MERK/JRCpK4rbmnPfQr5sLYpymI3MsTihVUCl2wN
Rs8DjY92rOHR8n2gv8NsVAeNrc2tcJajpoVOdLiu3uKo/+8eI7O4e1nTrXO6IEwW
cKM4C8zzckMy4evQOYtYZnjNnNyUpgg3egGMd6fjkjnY6BpM8lGKUxFnOKqPKXIf
sUmP+39TiZvqm6xi53db2TXY9XGB1HoVv0mQDVCvh07Xip0iYHVt0/6+eteFwSwY
pusZ1efO0G7IocZH/+/ri+0wqhOND4EVVI0OtJ/9ekgEbY6lF7szsBz7cAbKzotw
DxvT9JbsVvoLYxn6c7Ynx2hEfSTSwR0SAGa6kKuzAtvr8oQFC1RtRS5ZUD7KslI9
bNT0cFEYa/QsVp9cLS2JYI0uluvr7aRsgSyeE0FMW3vFDtLIlOSuVdnXQTsNTB9h
381rZjrSIDQh8ScX5fbv2vYgrtWSjGkY+TRFKRCdQoZHJuyAoogsfF0FOj2xl3zx
CJ7ayHNsaVLBB6SmMxI3CLmLkcSXcKq3sJ8IB1Z+kHbxnGqbyIdR0HoPaJ4HD5Yy
LTJjRoKPyqBgjnN6dxb5VMngYZFpCq7x61tPesgixOmwpkwc/A9b9MWB64hfr/vH
CsvsgIC6lz1JHVLpS9qVqbza/lGn9ZyROSyX1NbCWS6e1RiyJtMeUTWEy7DmtSr8
ztxtMShu3j41dsi6Wi5DZMWYy+yNe3b2x0uOoQOwvI8dDQHy1A12JsPe6S44LhhP
CVeHQwH6I8K5sfaBT4bAlODdCXEu7sysid7ryEC6yezHIKTMQNi0SXZ+3bOrUWng
49wrmJpIMmzBtpNjThpXn/H0qUf2QikvlfIWixEgX/cA89jLBYJR7DnijvMBxiPb
ItyG3Fudw4eqmTdu5luTRyRmWasQHU8p+/loxbA+BpsaJ172E06rocEGVo4XAoJo
cyovfQP2/XECierBi7Vx/+1nKDRGdGtbQ1ZkNk7QvlIMvoJF5LgCvhSEpqsarU6s
7sbUPETZwtsXO5EB68x1SGarHd1ZtBCh/RdGFpfGnbouHA/hflX+8+wvDZfdhHKv
I5yGJtDaMmHvxl25pHhERukdtn6gZDJAy6l7sYARJMG8pku8HZz0rIDSBItVcOgL
4F2wiO8pI8TXbFzWEy/IEPAeNv1FRYvtpsynM1Ty6sUrLCQFDD2QWRKZf/YxRJ4n
MCbSNx5WFe7/f87YY7kllwZphhKQv1Jg+l5h9QN6hWoxdaAbxx+Lna2JpSHBEpJ0
R0T0Vk2swNposK+ik45q1UUr4FOZN+aVrWUFipKZ7vM94doZRg8h4eYo4lIpNTf9
2IBQi70nXI62cOwzGwSYmQzOQDcq6RD0giR/US6DA7GKrZx7F6U2AD8PDT0lC77x
upGw1/KGLqpH9eLYvOBzrvOp08jBMr+zsvVoJG6B5tElFQDD17Cs9FPv9APzU/LN
SSD7eTVSS/ie68ua3VEZUJxLdKMg0l5rhhRLHYkkxgHz4vLuOh+v+swRXrVjngrh
icQTxKzP/EqQUx7ZUgV7wt3/1Nct3JWZ2rETPWHecYC9u3zomCAPvuHXa/8F7BeE
QGZKnWsPxQ+aZ8R7CAsnHdby//EQ4EgCAkl1LcpseWeCdJBez3hTEl7cd4zdiHI4
Jq/nzB3RUSZ5hqNDIDyC2PCve6/B8P3uDHQ5EiJuSWfTN5t4r/4qWSnLdEVeXAfX
CIWnje804iDWgGm2M1OuWnDkqRRznmyx2uOrj4CJCIYDZmf6A43U/igdQH0JsV+h
3qHWdOuyMydw2EM3IjNakHxjns/FvkQt6kCEVdJlDymJGTMdHNAiGfr2r58fLrc4
wuSMtKshoI8blFropWvwbbB8eRx2Bw2tUwYhXB5lnn3FGpuNbMAPUbl6BFil3k+v
Mp1uEOct3DE4BYHAA1v8dg+nPX1ZX4vUQKJM7cKewFmyNGikbo71TLp4BxitRlft
SNFct1aizLUXcIIxYUq6CLzTkRbjE8TCgV1IYBzFYqYO+BDlKExiglLnGUi+dwI7
2M/tn5t5arWcJWBbv2LMM3OV8wiOfmWX9fh4TnpYZ5oH8n+Bi6ivyQFzKoaK0fTU
Z9+CYlhgp54mnnG8BtwgoX/wf8MfC3MZqxNtyhiRoyWWpneZ7Id8Ni/vmIksyYeC
5c+0c7QoFF7NtRf7PRbk/RmNAYo91e+4Pwj3jEVlthAu+iCSNagHSiG+XfzxduLC
PF+EireTs3glnmTgpgTwaRE2XDI4SVjPPq1OYl+6bOBDPeF5wUZCcQzgUZKKsh18
19R0+/XhBksXI7JrLK987mMWlBSxp2Ohns/t+BD0RzxyhberD24dqkplnhrvW38K
8PpU90HXsdQ/3mbSOOZZWCoXIb9uT+3MhhB0dadXSxpbSy3fszjCUqLH61DnqIZ9
4InOQ66O7d8OQ/DLGeKMLWmXXQ6Uzfd33yr4YwnHde8cope4H2D4bzz1xr+fpuwN
A5/O0C+c0lKpiam+G9VJ14k0rrpzWBsBobGAH9G5mi518Z0BVptII2HJmt77xwTg
LRjJ3KMxGYydJEPM/WJShCQXeR6Z/KAogWVbZuslbpSCDQeSncogvZNS9QuExR0N
XQZe9vPWFIPr6araYv769eSrptqG0dwkE/Dw5NlVKKc7VQB+yYJ667OSzdqSMBbL
Bq5Oz5gEUlZ0tSSX1bG+49Is96IFNIzF6/L2mN/yyU1h8SRqyO9cH6ioV64ScDoN
6f3FNQz3Np65nD8eQtptJL3R18TECNyS10GGFPrvM6C6kmQTkkv13uWlPR6n9bkD
tEsQK2wjtpwIafInyVpYLQb6N0exlJdLRZT98FdocCmWItP5UoVkIa/LWAVSCfy4
n/lPGUhJU///V0ITQldQqd0JS9Pe+yksQm7sqTazkZML6IJA+kUMYh6OhrpLrhQs
7/waSS1ed0quyuhgc/yS+qrRjVXGAPlNMZabn55puNsvNLyfv8pwmU3PQmBNn3vA
MhlKFSOgb1OYzAx981f1KW4yfTgBWwrB3ZuwTEIJisPwEnpB+SNS0vZZOxnHq9A1
gNvnLBMJXtaX5XqRxKFg1w1KeO4JONtIDD30me7R93PXRxCkpENKMn0MkUCmR87F
TrzI52hT0v1tVaKRCYJ9cI6t2fwFWGAA1n6nZbd/US/wFqSYm0yj1hKVY15nzYBM
b5MiBxU6H8GCHJUZDvpL1YoQYGrKx105nfTGMd+7i0CPbEdBfReLlRvS3k1PaDKo
XF5Tfv9D76X7oqTi39OpVn3nYPekNj2vBdz8T7jj2MnyOvxfv+rrX+gbGzMhx8MQ
UH21P52o1QY4Kl1ct+/wCuGIpRoc151CDQEZQ4L8Omje8ZOLANFT1iPbhf6yj1hG
owA/oNj+DcCmVp1nTJjacf8Yf2qYEjRl6wDUwNKP/yTJpWLCRrECEcipSf+Phw57
T1hBzTq+Uf5w6JLi5YrWKa4y0xVrhgkpB9LfPvxNzb8PsfMoOMZ8br0CH8L8veEZ
yzVC9hGaX4Ebfprf1dR4FFmgqTelWxLMzYuy9V08P4bwJV/0IXGRg5WHIzcWNsdf
y8nNaCmTwVc/Xgfu9NGASE4wNUKEcmnuvrNGPe05pr9FZf9ezeDOlbrggpEJcalx
qEcjmXdGWkgQswViQk6IprGpO5Ks0veUbcNnqYD6RAn17CcjMHCQkAxjjNdoGYsx
EA2/FOD1HdYtIxqy/X0ALcH3123El0UyJEQWZxHSAohh0HKlKaVSxyXbjGxqzoqh
xa/3kG1DfIUQyk6dfo4GihqSRUOdruIbxl6J0DNiMxpO9vGdmQ8e/yvMxX7IZoMf
fCGyuI41xlhaBNMz7JZ0sdmw/WIslZk3oTbRPehYTmEgPcCWO9DhwzW+GPaDTK9i
fHSXr07lrgOtD6QoWDscdv5KX50RS803aED/22ysP6P2FHb8H8dWnLC51PNSa7Si
4QxRLMJegoummbL5J9qlDohI8rq+PrVGiPerz7k5qhSUyqxFuPqrDzW5E+wfxh1D
VSlg97tQa/REZ3wSU691MacgkxGr65NI0pgkjdc++1vwTKpljzrC5gkjfaclacKW
a6HcyVZ4laB2VhIYwR2fozh8e49KULVAcrjRxZoia1WChQ4XcP5OfirFCRv5evjC
ZopL91pRSkPfOucEj7en6puT73MQJQoBQXf2RASHk6oLF0A+Ux2IQrbDxxmmuE/e
eD3HzHpUHrpQ04gLn03kzJsIhgKdKuuQL9zm90VevQPhXx0vNS6+jpcjizhg+7MV
liFbCUsx8B3J2Rxzw2xziRePo4nzAOaftmo/cTvVcDPtxCIaGA+oFWCzWowwnWmU
mEz5h7LEMmmbmM6re5OAGotdq8WuGbJj+NxJMBRr+h5plfVh3Sr3SRCBQ4Gu8T17
LM5Co+tU/R/S8pTjzlqjkYbwEQCCAR7CgfXNuxpj6ZqVWIX87V1/MotmOj9pFEAH
BDPtgR0RSEiHPKH0nlcSztC5ty6qBd3SQM3PspNJYf0zA1Wht/gV3IHiMqgRiFe3
t387pps0Lg09/C+XisAGrNaIwBrtAPu2uRzd6MUF8dA0793A0ercn1g4w3keY4fW
n8Xyyhs5BoyeVe2y0Y59H1pjVDptfxEqtqomWwN5HVR8rtyxgL5xYO9fGS/FmSfB
Mo5/LITPsiELco7nsvU5PvVegCDZsQGfn44rDM5B2EYFSqs+UC+fcukaBlo3qSuR
rgQ/yeisAuqOZgQzyyT5BEH4FXzDJ3nfish6G9x4UvMM0VegKW2bpSWprn4t/s1O
kLKuqM6fPQe3qemoAuoQbQeCq+g6nsFBg0swMeash4RJYm1BpF1ARX06tTAyba6a
VTcFnkFm5g8QNdtp7ADU+2P7Ku5reAN25oE61n6doKXX0XEgHw1lfT4xvIfpWo3Y
9KFKWY3M66m8NyfEp3yAIygMADuHK7GQCA3YH7hkNxa3v/A6iKNkc8VsTIhmKjDP
Pzr+Jff9mTBECI2jp4gEI5xAODX53kCtafbOtvfF6qpWnl3qJi3KxYttGBdPewPG
hIGaBwZb25bgtGSbpn7CcFoKs2iaBR0fghPg2tnu4jNJ9xFU1M8JGpRzrs6ja7Um
dvYuMtDWXA2VM9ah8IeMMx8HqhFWUCqP6yG3BnHZcXqeREjzwsvLpXZYt4R7Pw8V
tlrWZzt6agANVpxbzlKZqBMM6ShHpu5QtvaD2wcjnVzSPR4gkEBFX97H0bp+PXgj
afnqFG0Bk2pcNjDYLeP5kKIeKpLb2MDjrf+AxPpXeAP1FqIo9Pi4qgQuiazxLEOi
DgYA3idmxqDCijkO6n2YXvTi3JARw6BSv8jbmD0X8I5PVN5entblUKLVtekMG6fY
1qUnsXtOPJ2XqzXV+vDxZ7jDv5oPWhMnaCDrRi2/6giN82C0HXUvB5XovFbOxv1O
U1U+OCu3rlXbGkT5cTi/MQRDbY2r9U90TxTSA/ss+gob/tFkLthm3nOq/9BgSS5h
FgIL9XReEb7zOtF+3LyG+x4GTyVMPe8LUmLbbZuU8VQFRb/vAlg/MZZP4YRhpo7X
V2xNRnH72+SgEvxVWgpa+UW9C+XPnVCcza0rbqiNj6AWtEAOXlbKTqorBPLnztBe
jE6DakJc/2b4YG7BQVOFnKIpAwO6W8kQEy9HsQY4pLz69n5MS03Y+2YdQ/qiy+A4
ghdaHz06B/IjeotuVLrPpMRE3RvktifHDg6+Wo97hnySDgqktuTtJNe+ltenLVb/
qSo2xZXov2DK8084DoFiBNSY3mgtcuGU1+35jIu1RywqZvL9rgyblaf1TryxW1M2
6eMRCzkwjgSCTnEJOI33r4ipqyjOOklgZZfLNvehs5Fpc4TQoZapdXr116iNBMto
usiVbDkqiJETOiiwLm/oGqCWAZEZma8jE1kNXVDslfNVb/q96JeJ04+mnR5jIGBt
QITQ6W3nTVhfkJ/ir0TXQiTs0jwtQYA5LHD1shrsnBj12Vr0sBaufYkvoN9NuFRC
xSBsxb+BZQNJT0iqxu0HeWupxCVpPnnNk6+dkb4TL++v5yMoqZSH2N5Ld18EyxgX
KFguWz3toZU90Wj4yohuaeoRSMfoC+xsRYTLhw0qIg+GWaNrYHgxQK74PcZgl5tQ
BGMil2ayDhGyNIub+NnpeWYBx+qfqrucuugUpXxrCZlavKZlJXEFeVGbFlh5Alhe
IkDFMDwPgKeFkaWhCWrFgLYJ8nHXLH143jlB1svgUKo1F9TngZmwb8WxqD7zGHnV
wPdntW6QYRwr8NYmVqejKa4DNb/hPnG3bSUClzIV7H+HDmxU6VNQrtZGdj84SURe
c6tXNCrxsdnMSZGSxKqFhtsFgnUyVniwIpMZgsmH8CISN0pEiEW0TEcDuhZS/1jA
Kf4VBORKS22aNau1O2vDt0S6xJ7XYAY4W65U4cclVHvFmgw+eJUi2X1wkltNt4VP
J1OpuYtgPWlRB3xkdTZJ706cP0932JGp9/e0oSoDcrFRRWIMhjWk6XD5KDGxwQcP
NNNamc0ytlDOR61U+NZ8CJ64xx9exLSXk9lLNZJLM4WX3HA3Upb7gnAqCHMF7VjA
QWDZUVAGnX9Z4aa7uOcx61J36ukBAgfQOrkYbt4drtWjFPDCcs463tIXk6CR2xCk
l6lACQYpLX7hHqDIo3PNtdlcqXP6YAPoUcNSVML3sec5pcBQXqu/2WHOdMIG0ahO
mAj2FAbVzUoY9dpZ2idje3ZtxzmrcF4886FeJ49pDgRn2Y5R2ZLy1LFxxr8jJxh+
fv9VLI13B0twJtQ1PfEMQdGIGz2+TCxzgP3sjTJ4KYKY0B1jJw3kcKFBd43xlgMJ
zIs4HtIvSzy5GMgGmB7Da1Tj05hyeIoMuFa1Lgjz5R7MKWtAyDYgdcRn49o3LAPF
LjejgP0cIcN21MxTG6zE/jxgkQtx/ydm8XAq/Tx8nZwxjltidxFGukKAHdnsS2VH
AcgLIB89dt8HKdYvMELwxf2gO2NN+euoxoqwoo7Z1mKRSq2y5jDJRntkA1Yt9lyp
u8kWjmnFCVgmo3S8iP6hOat0JUvx0sJG8QLzkmdky+16Zo3TWWR2kZ8XMkLTb4BF
frseLUuHShwgz9VeS7TQFlfyOM9eIDSVOjvDFBejIbKW46TJOT1S2doJht98FVxF
ozrtL+7ghnmf0ftB92dyx7NypT5dvUmmtIH3bQTPTBi+4YUa5DY/bEiyhxCAc45g
//Jwmz9IyJcgNf77fYboWGg5c15ebtLuvX2rLVdJ3fKBQ+AGRfV58kax4IpPJU2Y
iDPLNQQcLquRI+iXNnPEFJhTW9gmjj+cww+ytHH7eMSjQotDx5np+QBXew56PMHt
6EiFSSQXg1Ly2Ec1T6VuKn3cgVnOVJ6bC/XcL1PRbsraY4Gtws6/KVFcbA9jC9qe
X9pt/7E9f/ELGXlZYu6cfF9lqPzG3Qdd1oF3B1Gb/I30oHP3aHuUJuGyuo0HUFVc
hFlaKcaxV3SUtbRSAZzqokY+bdureoAp6Y/OZl5gWet7dXvKlvpKdmYFN9E7Nqnz
wnbN4cesBFrvmBUf4Qz/g7TZDLKryeEC2KHpNLu1ZvU1PSa5KXWUVutEevnkE5fA
8ByCV4+8NMmu6jFungn4Wf2e17VAFSIIisAAvx7bZ2oVD4xB20CiwQlmgd366G7R
dyvyPe8FehfxVNDbvXruZKCcAAqGeb5Y213teDzI5GJsFYJ+Q9hPAj+S3rO0wpPu
MBaAQsQ930yU0PN8v8X/+2b6DpR/EBOzO5Y9ouSdIo17xRuIU5xZPu+Cyvoo7P6M
RL1Qz4Lq4op9seyD+Qmom4Ip4PdRSlI8U7VX7tOf7KYXQVhAG7KFZ91DzPAxskMp
JZlYaFQ7XZdXcZCpG3Ma2hoSkdUt2KkQQVFPyknQ0MkWKHem91sKInASRLRyZYy7
uNNkgFAQB+og+MB/UtJKx4nySfi01IVWo6W1Jq2LfNxnLUZP/JnP3fcYgBEhkFOt
Akhq7N1mMWFVM4Q64VOoX9OaNgvXaop5O5TLG+4uG6QMv3Lt1YWgePbPlDkws+45
ZDHYNWBJDhyMlwlaeo39+PEaSYdTqiw6qktSBW+o3oXWm6gBlNhP3lcEjUUbiUuE
hJMbLLQWEcE5g4SAJqfl0m+sIJ1XfgYVpz278+8OErXsvUZInYNQanyYITy6Dvvk
2Ku23KLoKYbnd1tj3QzPRtiVICJKsdbNfGbqqrBhSXWgml6hQvflRpngPFcCj7y6
3Vnb/1xq4nlEzp/gm+/BArRyKyqxRNrTfVulnOB+RGSDCHJuBG3hxeHIWHAiH68x
eAIzd7W8BVnRv6oBqXLTO2YRiSaBOG9USQEw/xumSXqnZ7F4+XO0oKJtlQgVAvxD
f9WhDWC5jWnyhK9YFlkuo0ftaiSzLZhFmsz27w34DgNM7l6a9Jmeok+d2BaR2X8+
Md68kHwGeWo1lV8SWOUrS8BUVi/tx6dYmGiGE26Gg7BtVYChDOhyQs76c0kT9Nim
3lULDs7awDucyhJ6/IviEqL9P34fd2MMLI6Q/kZdDjIz0AWiUXbmpw4EPT92F9x9
w9VXIHWgqy4XtEEq1HkpTY0200ukTxPGhYM9oVpAJDKDT2iKkPjHICtKhpH4b3EL
LsPUJv5QKNTBzgiVBIltWGXzeUIiUqpdyuAJ074Obwl3idmofd76x1hrQu+EOAAr
bOHNKdbI1B4wq35V3yT28oqHrpEisA4vb4Ty9MlCdm5Jfy9EsSeo0NSRm8kSkf2H
b3oYPG3/e2M/ChFZupJaerIaCxQlMoT6jZVB3CbWXjsjurCDDkjL2pWsl+hLWMyJ
KdJXlyBixatKuJ0LyQxXXgrisLRhtbo6BBEz92vY4YjSy/xTOE+evynGBUaggk+D
XaoN7HETsKh0JYUHYLkC3XnsFj3COZu4EBB1vtI2SkKbu/G8a4ucbxI+UjQnP8+U
Vu/fDb4I/UH3y87t1iT6c/PTdAX5x3UxqQM7j4XIQslxfA9tjz9LDIitpCJ4V3Vp
XQUo4JqTeFKMepwRNGzO6QTb0mw6M8+HDbf0xdrY054e3da8AZIsMjaf+VYMuqtB
mSjnO1dXxuxmnKZcMwQUbGyo1pzF0zXbBeZ+vC80LkPcN7ManmqulCI2Q9lDe/ib
AeQclzQJPgwBM9cMF/wrxDxW9xyLw96bez3UAv9TcdiWt3GRjIPvpHls5/oplIuQ
X7M8O1BrJoSt2jKPXs0V+sZb2ebh82e5da4/1uLqG3FwEctq691QGjGuolXKuEqP
Oj9hgFpD07gi1fzbeEqh5YMYQP2ULU2R8+X6EsFBGht1DpsnFbfDuH5HM1KDfR2P
RAw6aAbc/ropKiK7Wz/EswdtaeYiYVWQNHAxi7agoX77L/kBhFU7bXWnm72v4zo2
52SLNSfs9aOzXtDmX5GvplO8tAFbUWPfk5zJE/k+lPchKKvMnb/yMF3EDcoDxWEI
yqPr+TRxxnnxVBx0zUZYyFUG3HC8FrZ8dneqY5X6LJzI4EFHbr0i0rXAN+LH8p3n
6alAt4XN4aAWVaSSynNIEwWz+spBgl//uwDZwDeIiYse5IUYqxrOEfV1RgdlLysw
xl/BNMCxm5hcwMFvh3MetvBOTgW8ahJtBavUj6hvtm5nJDiDnghCZDpthX45+P8u
wLkjjj9ShwAEjzkaGZ1dKOxuubdZ13fyodnOp2PPrSXan9PkEYrDyaNWafN81h6S
c9aijIacEwv9SRuPX2EgE7oMO08BcybMLCq1B0Wt7zT8OHdN63+03nB9hiQtXMM9
K8wc8I52Jlf4KrFmDxNzZ3orYP/ByVq5aa2/1UopjQaTSQYvLIy2jQAjkw4CqCxY
chYQdqVaQyPIvF1ycwLtGABFAuZ5oN4GpRa3F+bwDSQvhHG45xK2Zr1mOaUFb4ai
hIQa2saKBMt7rruwTH9Wg0k0Kk4mPEMgUQtf/jKL0BUO1GROKC3pFeR+/4YzDqfB
fjW05G+utVKNgQJ608SgC8rXJmRAmx67W39q/yRXgYCs1yArfCZZB5IPbu4kd9LB
6Z4peePutyIZzCQnTRFzSCyNrRePaOmL5Y0C2o0Hptv300XBfRYjkJadW4Cnz3wT
0mN+PBGfN3rK+7jJMIVNl7tWJOrSX0CGKS++pvR39ApJ/W2XG0JuiyfOykxWROEn
grnx4aOpfOknIe+RgSns7EYe1ys2IgULBwmChv5dph8C0Rz5Fs0xHPYnLrHO7p5h
ztdRCbSrkpYx+xWvZ7jZ+KBQZ0Sy+r11fUTJE5Kj1SmmxMsseQR5SuXoVCE4VHhs
cDMQQNg6FRHj002LufZQAV29y9tHjkdj1LM5kIzPeOeaXL4OBiFkZIAnuQRmQ1pV
6qGoSHxArIqw7cU6F3I7i5HkMjfWmqyiOgkcWS3r0tzKt/YXlN19s9Gi5c5IwlxO
EQhBlE0o7Lc5deyZGO2Hh4XG1NcPFB5uE6h4p1/4Lncj5VodHydsEU7Vl0zrllGU
U3rVuK1Fq5gvPVES/GGWbc1bSTb6LWCpRAOjOlMbFZAcqPiz+GXZTWYP7pWObvjx
GMSTEBJfx3QGDHR7RZ92E/wp6h76NB74fNwA1bTF0/jF3IEoo7PUdinKCMY+z7q/
lxAjXyxcp+4NDmU7HZ/F4VYk4NDxcUjyCetHP5d77rPtFVDjFZ0tdVdxRFYW62Me
ESS+zGCe3VRf0EtYU/LsghPY2Uau6yUtJC1GknS76AUniHDYARk8lIPafjU4dNT4
H/x8Pss7jA5rLCI3svt9Qz5qhaDkfpaXFXpNFov/6evfiZ0RINm2Fr7nJZX/FaKe
yXfYRAqLwo88Z8LHT5twsHG7AAYC2/Ks4hD+w7Ox/oStnlVNUhnOxZwAZzWoU02s
VkqKf2LunCns3/X7ONRfBtWyl0jrCNJqfQSavbl6DFlKnUMbvT//7Mf6TTj3ZRlU
JsT4pSrxow4XJbqRNZ+H2TzwOWn3MT3+4KbmS867q1SQfcl1Nsm4q/sNlBHmm/Q2
iHRCe70tBf32lP1B2pNd2sdNRn4SVLXT8aN0Raekl1DVRhftgargDzPYOEK/c/dF
IVS+DY+Xw8Zr2Vd/+w2aZ5GU80Q+alagQKJvTMwgCXkJ3YNwmchzuJNr5nf8LW9F
hHaSiICs3eyUvTY69ys4WYvUu+Y2Qg4hZ2KQu6vm7AmnRhK7GINbTTTtHRb94x8V
kNJhFD070BYIB4LDR3e3X2/AGP0xkwMaN90xwG0MsCi6ybGu/rGhokHXy0d/ZwyJ
NZ+alzOucglAsgMgTxX38PfMhUOnwP02uBLprOilzdXE5/KMVEydOCyFTyNiOhkl
fRnvLWTIkWZ/IHuWAXu850RU+EU6tAO//PiQvfrIO07BK4unEt93Izn7mwWTskOn
4/2E6C8e6SivB4G8d2sojbIa4ch7w0VbMe9seoNuaxHdJzD2bMuLE90mhxBXZ37L
U2LqYYwFZmPfxjMQgXwgKlSqNuOFAC3+awU393AY1IF7jUO33C5CBkP4P7i9fqQF
Mh83QBlJSdA33/+F56gyLhY0bfgV7196TCGfHI3QyuX1ourlScmP6DUQgNM1aZTx
3fd/iYqUqDezIaypqv8cCeydQaM9JwK/OOe+Kl0sXGUHjx9irsV3Jc17CeHpoLvA
rWBdHsjfhQ75IveHGHAEneB3Tqrmq8UuQzq/OEWMUzK9v0dwzU8ZeZfszO4awdhH
Mg0OhbUT9uuOzzywAu6kBkRFx+WFxB0UYjs/UCOJAWWqNcLPNRHxXYCoa8BDMkQR
MKMgHHcVNAoMAzAEKyJb/HQJ+ZVb+jvRP54UszmUfJWq+0es2FHAszdaMA3iJD21
+TbSV4c8yEmwr4AdgQVR9ySmrzMdzB4RpHuy1mexe55vprP08tAwfZ8MQlgs3eUO
2eLJTCdfHzQOLDmr8eKz6qsAh2lzIoP5KJN5KcoGJpdaEgmCvC68v0z+MybkA4UD
eRRSWZa360flOwmZGIIgjpYM98xkA9ygbLx4skcWm6IdN79FtkcFsL09Gpmz3cnQ
YoUz678lA1UgaDebQiCZ2HIwfr3OKwWI/20jdX13oayEqHFl5JVA6fCd9itVreKr
6faupqI67DeV+RD6a1Itl6OGgb6xnsLFe3bK7bFyBk/Q2nKegZAS0s18u3GB0APG
1HEjzXswvkSHG637lzc2A+6xLTZc197zymD3XSeaaVpNqHL0c14ZNq7xNCg3kqBY
GBhMU07u5K9YqQ3TIjXpH6YgG8+iRHx3a0UtceMoLcGroFC5LMWLeCxpaSWHKEnO
4dqwO2K4kde+EKQ4dJUyeECWABAWk7oFNUoMZP6qnsi1hO50PSYckqHNJS+TptNV
K56rjF37EHnppYIOIUZm3VIvvk6gHF4QvF57ZSaG0Iau16VtGC8f5jucA91N6Yzg
jnreG1JxRrmRRQNxnpa2fXGOZwvA6T1a0HOPOlrXsXzmdx39IuxoH9O797LWZh49
pEW6mlndrh8YNquTXgFX1bA36NAboBvqh8afBAdG9585RBrGD+kz80CmEsv08Km+
EW1y3MKCPYbLDxWY1sJ+E1DcCwElMiPB4wj3S/3JZf/0c8fUNqCsqM70C2QTg7cP
YF3TkjYjTA1BU5JjuluMV59mNmibpeBQyS4v2SHop/fSHmDO1Thtg06VmPznctrJ
I1YXi809vNaa608PygTh16FUmiZRIDadvv9ZnxUj7G9WPwSJNgBvMR+da/6xdrKf
8U1QlW0/qYvTItnzGbUNl/G5W4NL+g/c10jW3tcK4uvDm7tsYAwJiLZT9lGp3wFn
P7Z9f+2whyX+PDKlLZLPrNpHzjraQBBycN1Ila7/BkjM9cPAAy7Gt6lvMgjxq5RF
SaZK7aWHAuwWj9VSvweYMiAGlLXeGe+AnN7QR+CGqhrZazJgS9zKiHo/wGrdCdLu
6IscZ1W3JiK7cQrKjGPaOwhNQYZoSh1F5B20gi70nx1GyvWkq8TxCIX5jAd1jN0l
44J/v+IvwdieGjGTyiliD90rZcFrE9r4D48uQ96kCqDQOzwKgh+mTsKC3vYVaTrU
ZUiyGtpSZWmtCCF0m40e2bMBUyi3fUwtxbDGjv2eVwg7Fqzey8Cp7E1hCPbin2jx
X9IUOYiBe5/oeK4KWRkEItYCVReQicLM33LMLlitI+G4NtaRVVxyU2pTpxi9CTY8
I48pBPXRJRwa6nyKYKFL81VwJfhQlSY+p15IAhAIeCY9gjQbnHK/GLylPZIPWdSC
V/8SINowrTxt5HZXeXrAz5ZzkUJJkh9E7I2eBSWylz28LDu3x0EB7G8mWQqsFDLY
6yXachiybIQeMZXbp8VUlT7TkM89Fq/MsONqRI+K6QKvIPIR13JoXYk7TnLdz52q
XPzAoa8FYx//KorngrHxmxFEC7tPjFHGtfcU4HKzB+VEAR4300jvRcvI5YzdQgOd
kVjvWkhwIw8jjDI7Bc7G5xPas7fUblaqvpyFwAwCmkXxr3wp5QVQScHGj07YG7o8
7jsFt5Cz2pyx4lA8FPRLtO+B1bsGHLc0vMBlYlf4KF86CjeCYsNXubtuu28z/r/4
X0Ndq3NEBKf4/hKoOu9LtVRN+OczCMXJYH9xqZbtYZOrr14slUy0AqnCO8QVQIUm
LhoT2is+nB/+EUUCjeukV1L7Oe8dVYVnTjNl7vqfpStVlQiq8Ihjcsg6pxwJfxoz
nFZg85VktSYFyPvP5sfFU2p6Hnyv8VlQEUo1oZJ/AX6Nfp1S2aEmXgERGdJqB3p2
kVLQpezKziK1IIXJ5fq7HkWeg7dOkOnP7p4ouhD04bTxNaiYyYDRc2btfQNnrEAM
Ays5yGiyfUh6wMW84W4LKZt4iZCnWG1dOmsBAArct8OwuuPjiC6r6UzkOlLtYze7
BnjxKNWekmlQPIuueDR50lzi3aEtD5c9E7s/prg+4qgBpRD+ySNfRXfYpfqL/VSH
y+CkpCCEYKAu3qVS9hp+EgpYQxwY9H9vxE1DAqv5n21vaoCfHq7cBwG8rssWR6Ju
Vzp/7pxf4VTH0lUIQpBO6SUbqIjwGYj7BR7Ux3wg47o742yt9Z79a2s7BNX9dSFQ
JpJEk83n+J9LlejYTFvw69vyII5j4abXVMwhl/BtYLRL8lOimX0FH72mOSXjVEzG
G1k6eh910RnxZ2iUJGvr3Ll29rxPt3QFzjFepDmRFd3P6msKA6ueLeRsj7J27i41
+JYGmZzUi1ReybhK3UjdJPVoE0jYkCXoz/n4OaXUNn3bmOeF2C+7MeakNM6UjGku
Gv1DlYxKxmVtqwTjN4XYSkhMvlAXBnVLSrAytLBhk5U6mNxI6gejOcHhPxuGCeVY
98wAND617GS7gaEviSvleRvQVjXg7PiFmKBRUWBBvz4G87hwFzvvAc/LeRlvqLaG
N5UKH9K+jzp1o12pRtGBoTFvtIEflcCPL64ft3th0IQuM8xG+JgC6NQySPSFz6l/
02t/pv5v+akoYRVajWxvt3RRhozIhS2ZXc7YU8Lv2SfchomlYddRw5TdeMOUsbFD
irL6gaDLSjTCH4ENqbp+XF3fyUAYkU5wzhrQ9VTYZcAckLkjNJ4OdGkvzPp0viMj
JUAdtTbDHPx4YZkr1rQ6wk0E0erhpJAgo1X7LEjJrioLEG7RdcNcb2amX7TQfMkB
LtXfhmFBKEe7bX1ukZAAEaMNHnQx49zJKE06i7s0pSMgnat6y2AngerEAkFKr2uH
eseJxbJdeamAkUzkiO5Vdga4rwf9yyZ0A+en+gszhbgG/T7mH0AOlU5lHAXXHCU3
mS/06UHP4TQe2c18Cu0qP1MCE4HOdSm0OMoZikUYH+c8T6vFaD2Q9o7qGn3D1hYX
UtnTjrXSVpKBJhCyTLHpTA5LSf1NBMoYV8wGP59jInofufDBB3IdYRjSOg6qIQql
VDJ4pWFezdvhruLuaWuGUUr+P4Tgza/nM9IiQEiCn/X10EmjIWGhhYIRmcMlyflP
gjExmgbXtBuCwdnEbmd55q4aEjHrFNo4NNLm+JfiDlnacml/dvxxcldMNNN36ziE
jtoET6PuD4NIPZ7FOx5Je2bX1A+EmdY/dxJSFuAgtsMf+Pm96FrTM8cMOxvKuTam
2LMMRn8vaB1MNGOFPdFzGNzQYYmWz9sRXq794Qmy7mlcXDqbycmUPx3e/UKuEJKT
v8c3mlEMaz7DQ+k20OMxvh036ZKmM/U01K+pOF9/01moAdmd9LuSDb9a1OgrsZz2
0q0yApNbCKEdsGYANWjIPxHQZZcRXHUGjBTCqEynMT2FJJ9yR7SWj2VDzFzy40nj
UFKWytswbnTaZDsporRMLj3mWe7+sbs92DFZusm6GyQoRtn0pqYFph5DfYE5p3kO
Us/gqm75by9fV62vwXU1rwcqbFpnEc9wQ7ZweJ082s4qLwAqBeBPqZeI2QCYXFAI
7HpG3OrZ0OErSckan3SJijAjEUVjyIEZBlvHOU1St+acxFUjYUjVWA35XlpalPyE
OOoz5BrKZqtV7VYosglDA63IJuJWL0IV9tRcGZI1EtjwJmE5rqZmfH7r3WGkOF9x
vu8QCsaLF02uaENLaLyqCyg9O5RtfcNxr2bC/5rYef8JSr+tiE/q5R8z/LkcZjm0
2XGC1GsZdSViWAasr53rPKwVzsIs5JT9o0vMF6qWgOnAIv3Ct8AguMcyzqAnYCnl
3Sso/beNSvrG7Ix6gXni9wD3MhscP9X6htVWx1BmpbIzPg+on/XxiQ40l1VUD/lB
lwQVfP6ac7XM7PrggqJfHOci+femzNrcPVRR+d97Vy3sMhrGD8Syjom8S7+OuwAc
3uOqhpmsG/RNfixuYZ//YENDTC2pQoj6muVsrftPQTR4FwRHXrWPoT1LfLZetkGx
oIZ5V5Uthb9sfSF91JAuvfuou4o3Yx34sNg/5gu4NwKi5rZPWrZe1/bGvl4deDcJ
SkQDU929Fijo/oimIV6/HlibV2sOejEVyFAaHcbKd4LdQQYy61nxSHzEBoc9Zkx3
wMoB9e6E9Z1wiFq+dcym2Nv9bv/h/X588cs3Nre/sK+tqAMjG1o2ZhG5lmCBO6y3
+8KH9n9dl70pNjJZGYxKAG/WOsBdT8seeoCcZEa9hCZQz5ou35AKeg4i6HUA3sHf
R6Zy/XSHrI2bcmE5JJ/uoacIqjmx0ZqOidw0PcCjIo8WIfLyu62B4pstHksV1Oat
OzuWWyvw5XvmWVblzMt+gova0/EM4up393HuM4mJ2QI+o26wqMGRDuoUvKY0rGm2
dvHa+PEjqe5j/Ju7NoAyF1R04ZlvIuTPzpgCyz+3+qWDEPAozq+A/xY9uxVqM/zd
wmTyCN8SJcj3Up0U+BWKXHiBWCk9fdtrNIgDGuWb2jCPYbfUC4zmEub08dz2EP4E
MTLMnGrpqndbsICh3x1D7p8e7+aFSy8+UR6WT+p7RUAxOqEt/9tbPQwWKxHhENAO
GIQOa5XGAfKmom6B3hzFpu0ETyaG/5fZhATSUQi2gNH0FfrMXoCrvgLngCYYYmL/
hfwurL7Vv346fSRIbOk7+BNYB5uI6sFbnr3kvVvO03H5iZakmPzP8y7VNPV0kvez
iz/o/m0abRpbaHgs3AJpWiim10+UyBbnHvaGlYveTDkbKal3aelm19v0/OEg4Rvh
gSCfX6kW8hVO5kJorxg4d4r7xGCKBbdxs44xU+h8PqVKhXe5NRzcyxP9SIXmyrNb
N2QGi/cLdNZ5Q60Zkb+sdi4yMEhq6z98bFrnAw7GHjmbzYg+93gFlkxE9rkLZaul
t6Y1nFxs1XKQ347AQmlnJa+W/zEPSV+jP+ity4xNiEs0pLPg3J7dTD8Gppa6V9zA
N3eC6DUrFZtsk+5WiG0egwd+wk/Mtx2sFdXVY9ihTcW3dvvFyUBEsABLO7npq037
iKpRxD0JSpCQyKrqDoIO50M5Rf9ggndkHXLQiOxIXXrV5MfeOKy+JpJRSr3WRIHP
KoYMhxjG2DaVzxNuKOWESlQFUImANOy45Lxn3Wgaau2PAqoVrOrFQkcRZ8jbxSb4
rvmO+dtkCVYS8NYEGPzk9OR+SicVXIkDJE5AwDCWIE6Z/ImijbznJ3U63TqKmS/m
pHit41C14uHndcbVftUMeoxqVnsOeSUAI5syCHQKD1FzHwWl4x3X51FeueKLKRQ+
MkGTvhfR6FW19lLZEmwGFa4CCNNKx+JssHIPF2EwYrh1FfyDoUXgEDVvFJWdx25J
L2dDvSlBQOEI7brvMeWC+T/qZryXZaYx3B205jdk7eLC8k3DSjw1bfg0CYzX+/Qa
9tuordGluoTJUCE+TndNpIVfWJHkOek5bUQZxc4wDC2aycbX759VaLWO/YdiiDiD
l8+UilnHzvRsFky4VPDYnwe7f39qOLKS0i0oL/cq/GIeWFGBCZeyJdYvzya9XaWZ
rydMOchsN1hASSRZ8b1FDp4LpVVtGcnevGW7lx4G2qyMBAvXoQDTvrFHmMsCbZ1o
zmi0mqHHr033dF6aLI1RS98Z7MJ2CbUGtxlPRyrBjy7XPpbCLtU1Af1t64n8CuQh
hMo0AJxoiFdGrUw9RMZfBZHx4l5a6CvlQR2wPMQrPcWhGVIHLWjQy9Vr1ajlGAdL
6rBJYY4hhKZat03RXX110qqr79ee4UN5N+lp798sJaCeSa0ou364ZMJrl8MqjUaO
pbLUZCQZIwsVAUQ0Doih6QDbvTZD5N97ruwzrywCySoZz1ooG0Ue8jH+WBo0r2tC
JeG9O6+jdn1v1Gt6xMHSJYSgzS/ego4+xFbpuL2ja5kMuuAY2zlehZq3mdKkIhPU
j/cUZxyj51yVmJCVc5CDLLKVUaft0Vtam1ySNj8CzDidQcCmP0jIPUvTfMdWA/pJ
gW71So1NGK9DtcdlxJ4o3LSE4rdZgb5aYLyMqwHFVk6s7Wbt4xX9i+jr0hiwtbdN
TYpFZchGkFOVfNRshvdxPJqZT65YjUizQSqZk1trQz/Gesv26dqtIbb95Wucc93I
SmLoUc2Io6t6pbJTdi+IZSoZxYo2/D491RFW1BNwY5JxEdfDGK7cd8qb+Qft+1+X
0b/4uIIF70/YwGQfbegbesiT0Oq7wrw8bc/S2Pe5wueCegsyVltbaxgXTLgwU6+B
f5F1HKiv4ymhAAILdFKdQgkJDoWIk5yNl22QMLl74U0XPGQqAog/SWBt/OUqRZfr
hwRaD82Xrudz0PvZuaPbFR5ICf5FlS716Ws8aD0ekHmAYqD2dWEfJwDdYeqEirOC
mSYd+RgIafMtjS8yrlQWlKZPl3KRFuBmHkFagY7ll83AlrpWsB/ZO6NL83Df7zoY
tyNJ3i+cDVfr02T4+JQ8Kq5F/HPORgULdAVm+giKkOHgDymY3AlM2eVyNoddOOW8
s5Ldt8y6v568Mhm7nXLDpWojvkmYxSDyTDtbMYX0ZbWuSz0S7HfBxRd8/Y2xwdSr
zoIZM13JG8wHLICRgwl1CYLCm7Lp8DEbB6pwSHiu5D8TakweQ8op7i/H6PAd7k1F
zlndfkesN/2aDTqB9JX6NqLosvI2K75Daixg431m8TeAf8TqkhgACcs1M2nSRRpl
xDbxNOwrqrfAmkipJpuBjl5yOC9nQ2dhYQFhewb2lW42+BwTrZFx8vRKFZUYynkA
bdp9ECtykmU1ReODO802utullzzLDhO/houGFqnTJEEEYcyOoOx4pD64EP43dy0D
97ZXM6ElrkCL2OYVUDa+4Rny0ikqHsWjzzrq4a7gkwkmkhFajl3EbffQYhg22OMw
aIEZEYlyLLTJRiHOHRrDhGjtERh510JzHbhojDWLw9MrqetU7WPhQ/lHlR0MTueu
0aajZG9DYjEafr8R2xZxCV3lxL4dP9hdIgvl3sEiWZ6/F4iZEG+BCkV08+quhASL
hB30Q6RcdK5521lTiO/USUYzaHDjeS4HiFk9+arHQLmw3qfsZnk6lgLNWMAB9Rce
xabMhXD9YkcTiTP7vMeEOc6VKR/FqT/vxTeI2JVB+aUGYjC8IrM0gm4OyjkM2nu7
prt8j3pKW3uE2ricIPnoQD5ZCLATK6mP250rnoHqT4yXMvgDJsi6EW4QMFf/JSjE
KzQzU9lDTpiKrnvc15UD2BIHqJSyUmilHYBG5JElskDZufqf7pKUjwKZODGAaKmJ
aIlK2kpKk7sawYfTrVLCp3qjjxWlwo2gbt2T0CetQIxm1xXARinzpwzEIrHJA5+e
zAIjavYBGF3Jzn71HxTzQ9bSmjBn5aN1uVqRNgm0TqxYZcaBeUeND4eqW4fBpZNS
aHAG4xkdmxtI3anXsgx3QXTKyczPJHcJYjJzaatc9pAyvJRlpZlhTePuMuG9/b4g
0+arzMX35bKgmhU0MfxsCbSXvD5DktN+jK6KGoBJuo8aMTde0oB50DwkqrGzuOhg
jp0Xf46MnXRUDPTqr7HcDvyGHqrJEdcZcsdRHKDWbz/I+2QyX4N0i/EKKSQ8jqMO
H7BbDQk6fJRZ/Q/mxTAIGiCfrAOJRjvj7VMVSmlhNabKPhTVEnMQK9+5TDpnboFi
jWVcKhQ/g66Ocbo1PV/GaBtfFF2yJ+USVT8HTbz+bYtsiPQ9G8abDeUhERIgZY7x
ShKvNcBAXM6zoP7bB+M/yjYs3FZ4OtOMYgnsHUmqqNCsU3JnWTwy/v91+jUhWQrn
yJA97Eo9Kh/VhQJf2DJClVb/NN2gUFD+ovqVtiTpa7yF1XAZkJDk5N8t2BOIhTPh
o463jI+RGPWRWNAXSWf51AY3yz8ImLS0zFraeFYTLafNseZSjPIAkllIOo2DtviG
H+9ByPWM8sgor6sYXccUNKH7Su8m8TVCQRTR+8eWUKJshbWzyF/NUu51TTnkiUMf
N0PEtBOz5YKEbbzBqezhBvHajBRVTARRHOUdewGZ1F3qIVEHiYC3+K3RLyQXNh4x
jfCNd2CXCz3tDMrSs71sbtIjLKs/fxmFmIEbe+KCH6dTr4A4Q/GPQAD+4l6LN8Ah
IHhfKsLAh9h5o60VpQja6KIDezI2bhW8j6RQ+nB6hc8sOgg6hFB6Q3UO4BR22qtq
MPq1X3xKhBqjF4Tk0OdpKiqQruYzU/7ole98q0LMVtVOz5TMwv+iNKI/GO0q81d6
ZGGpU4fojrrt+lgtjXhKsjpx791sBGRolwoDFKU6hJM5SDZ6wNMKQf4wWbz1j7gQ
oBCazFg0CJ+MMoS/eECupu/4A7N8F3zTLqtTQVYbT7MwPr2djmwXUL7mMgyrqfe0
UaG/U+7V0xIOMTfoNGoGIFQvTW7uc0p6FQdzPpkjfJf5EER/z/XNk8sJThMJzHHI
CnRmIX/acdB9jPyacpuEk1tAir9MaEYI/t3PY11ysO6z+3EIpZc3DSVBNatxi1/2
MFgcKIdp/2qNh/Ok625JctJnbHXX+WcHYREAKs5JiXviCywEW9ZDsvSFRUA5SztG
FW7zHG5wyiVww5wqUdx+QURvhrZQ6O4esIuXXVGtIqOcIBnfxrOjC7RQtsu5i+sU
DL19+hhHb17dV9Zh7hkuvPMHTyTesTjzwomsphqfWpyBFbwv4w4Bl3MCsx5Bc3L1
QNlGTagS1/b13DSO4p8g3fdQNdmJfQRTl2WBXQ7w7mxbtDdKK9Rx4io61Xp3OG82
XuEz9zNcF/x6MdTf5Cq7DOCDURu/FB9pLsdSSAJNTdhyLu3foUZF6zphCbMRGkUR
Z4Z6NLk0UUCcbDmaiPLfhKnyr0kqZqsjf6DSgduSiodnPIPLRf8A0BZ6VCh0lWPW
5xRlvr4F0giP94LDPOyhgt2AWSLgX8gyz0h3iqfZckiundJpvjuLPQSmChAQo6oP
8yQydX6vB9GUhiYkG2JCbu6q2gV2Sr/KKCwjLW3qHUe7sv9Tbr+kHkhaPHKHevrG
TRQEI7fYqwf68aZCudU+QA4V+wfrOiufdKPApyuLObicdMzFPQm9YfAvPuK5XCBk
lHddMgT0/5eGGjMQfpGJdZG5h9zd0AIug3neIws3KvbnXEv9EaYJCZW+orDT76aI
FID+LRrNGqfkzSxQGMlwNbVWvAFpAMV5bpHRdvnt9e7yq1HZ71eBzsULQAvW+Cfw
/ZRanqEcFKpednKq7EsxT63QLpb2SLTIMG7wT+ypDffaKPC1kUeJATGiOpYkgeKg
wOKtpWZ61RaHYJftvnA2L0h7n+FJOSSD0WkBbCgALf/XNLqurro0cMT3Xvctl3zF
jP2TBFLcFGSOJTA1wOE1OcghyFJpHvMKVul4mnS93V0nPkk7Ldzzqwy93fKqBSyB
qCzLFfTHeQG57SxvqzjsDBXE6T/LRVZqhpDSpj9WS3rH5zs1UYCHNcZCI5XBXj+T
eqxdBbBAWWcLug+Leh4SRT4SM0WnP206gvHVOcI9IqJgAdfZeP3ThkvlrRFLGSjv
sv0OXN9tRsaks5zESJfXU6iXNMfn72H/rGmIWWGAzAlCSSPS1Sb5EW1Nuxm+zgxg
J3KPez8NlrDue/Hup5rLQslVH0Zj/Wr51C2Ne0l41hDbxGxwl8rOkXx3kPAG6n+3
zL3s0QGczxlKW/5b6eDYcJWifuBJzGGs0rQoS5I6cxOBc0IUWniwEa9duUGc+L8f
nqJCw4B9FbV57k8De72v3A3XssTr1G82HS6Rlg0atwayA77QMqwlY/POx8eEqgu7
kgprlpXv7xts54kxZsoQglbT/96tLZF6fAOR37CIx8kaS5qT3PLF8kUI+c3pY2OO
y3W0SyeqLjzgQ5t+duV/UPcfsTasHdYjL2E3bnt0I7FNZNkg1pYNHVTWBRm7tJSA
9taAmv1mIqJ8rUioZWYjEpOYW4MgwMGtd2N0/Gh2LYXTxkGM4itr3Toilz0wNAVB
kYOP5K6++sG9B+D4sQOncnwSffzisIiJu0f4sEBiCkHaIhuBWcRbNXDNltP+wF3e
x61v68Ameb0Ds/Z2mNJS86cEhKJc5Lm5Wp0is0V4sReZZ8WsNa4doDqq81W/Q25A
kTyJxy2dGSsDUnn//pMyZZEw+AnppG/IC8V/trm/ghcnbfsd6NQy+q4jHVAcG7bb
DMMv1kv4HKGoOGGjSuaH39NjdL3a/zLtrXHDHS1hPSynKt1QnTHABT2x01CPw8dY
0XM2hHgfYjFPt05jHihvdzo3q+2rr/FRUdn2p7Cg3/RrMflkp4VipVExJ/rhQbOJ
JCDWfvCdOeO/mSauKo5Yx2XASF0KWnbRxX2I6nJzzwsfGPeLIUGMK4zxmcy8FFt7
g2KQr+L+QuiNG1nJ7EGuiUmGcovo5Zp2zKURVuCJsjPpCgab6oKBh64Our/py7rl
XQuEN3hWKAQkA3KR6vIu6Fel6lTZq4vFW+Vqce0B0FCc6Zjno/cSEQ+k4X5118Us
HiC3TMw7uFZW8n342N/UCfc8ssEE7dK7Vm3t6UyUBzV5VWb5LMOCIdQETklYzOds
HsMgA+0AgyeUCU77Oe6kpqHTKKccO8M5h/sZ2OpOJErOaX/lsn/EdZMCoFyzSv5H
KV7LMGh2z2jRI/44u53CVBGmWs2TqbUFm+u1WyTZblMdh6wyxoFpv62R1gEj5EkJ
9YfGQZLvK9Rs/MSc866WNm49bX76g/ezgg5AK6s2FyA2xh38WqkHmsESIBbCX0Td
2+mk7We3FYw2q3SeStBDeVhFSXNv/skQ3+EKzq5FoI6q8bLYk00FPIivW4iqYRM4
Df6AaDk888X/5BvPQMv0bwkongNTjg7nBRr6tp2SFwAM/0Do/+x5SMHXYEzvJ8xq
rEknaBfu7UnClRQUm1tl0T7h76oFhzYkVKVvcOM035IAp408BrexvUf5si4pagLk
iGSebymVXAfIeF+7daGgTIMAQmgJB1+r7hLb/cMTcnJPEWPc7saD1Qrm9OuAzSwg
785O1hUu8noHi6fpFKNcjSGQLhXvCRtr1Ps+ZtUnhRNKC4Yzzd3KLq+RVjF8BJB/
tNRpJHYtsgzENvvv5o/eaRA6wdnIF6e0fC3cm9HVePscxGTEBxCUbZKUK9+GRleb
P2kvCptzUujQmRT8/B0YjyHLmBNIz+wPhqadb75bWPtZZwSPzM1miVUD8GkEjTes
BL/dCVeVdU3rhdFdOw1F9MJPn9mlOdy9HLzJzTYaKdFz2TnFz50+vdE+S76fo9Kt
6TGbdbpJ3gSVs6KSmjfWat9pZTbAnKTEtFwWt9M07ONaY4N6A+GiI19YXmJ7cBb3
MBqEryS8csiHQzj4g+gl08yFBR+DQUWuB3LwcdxC/MSW50UEgUl3ZwJhGHxCAdf/
Jroqq+e7+gCQEF/Sb0uryMP74JG3O3FTzp9LafAiftof8/ORzJT9nCePxJXrqebb
yagt6du/MFjy4d9hXHUAXM7Rx0mavSWNqOvCptd54oFNxHhuIU+P0aRCYeEuU563
2VO9+WDPnxoLoNyiVei79AZWHh0xyShhb0xtHSSmXmzE4ZMUAFc3U77hckzyzg+N
34jR1Rn4DgoaME8Gs4RaMvQROmXGespOC5HtQVDBkk5VX5/jwjMnROTiM4aHI9TE
jCwr+Z3K6si5INE6pdB835o54K1A9apLh0XZo8RbW0d+DlBL91HCjv3xHGKYoHas
zFJbsA4NYy+jkutMJ7sdkhEeTuB63nUmG2l0kNSLQYAlamo3zB44JAGppoSmIf7H
gCBL9P6jL1SKeFhOsY866Gsfgz/T7/Ko5/OKukdiSk8ed0heZZhQYQcoICPyLRqO
JucOk3fdAp5S7CDJcXKO+cp3wyNQhFeUp3YTwuNg46L6YQxFa32aQnnGVoHb+5by
NYof4zYCkhe/Q7IAfpIWE4Wvd3iIhl/JZ02F1Qu1KIfbnlcg22HVFqKa9WQB/3dP
n4uDlFMTjPZRLaAXFRspYc1H6bXCF7k4aNkbE1/tk2f2Jb9HbDmTAjU7KrRmxuV3
rFnBR50Zx/LwFST2qGXtD1QJpxauYFou/rCSJkhXyjtUocGDmvF1CtBE+JlJGyH4
DoRa9jfnZJHdnSMYMyReL/YOQM9bdRrUQ1PVU2TlB7hwdBI7PsxDw0PUIzP5vSR+
76l6FBzhWZzcJ0fdeAJaplQK+WeFw/mt65RL103yev1Ve4KyXr30sCkYkJ6LTQ4w
z8DgnUlZ06qb/tt9JmnCFYRH8Kj1OybF5SCx3+mNDNQnHrxNQKsYNa8eqlGXUvUW
mhBahx3OeP0HwM3E5Ie4YbaIiDqnYYtYZFfCu3xx6CKnd322aIVpl27WkEnV1yNB
jYmuoXXZvT6YHHroPTYQfWoTMfMBHsLgKiCJsdASb9nkqYkimz83o3oEFXx8FqgP
6kXR7unjjJ46vo4i3bZRozAqIL/92h/xm7BV+alTAiLqm3lDaqv9FdI1AKQwqpAW
9L+sIvVHgVN++suztuqHXZXy9gIMCCripwH5SCgQ4lSRtLqS8+7KKX+NsES2BEoR
v0ilrv8xGEM4ZIEjio3nFTzpsjze7QgwxaaSHP1qRozFJG9xtG9N9skbKtLvxa9P
g0gucmlg/yndpVIvZw59Ct1wobt8VgyvrOBMHLWFg+ilC4Pds+1mRtCoEVlu9S5N
We/6ShJsue/aBr6baq0Le27DTvTny34/ZZ8bRPVkIvrvf5OIKl4TLvth7nmXNCeH
frI9EmWgAkX/pu49jSI9o6uLN5oeaT8ZH8LXbBPG7ktOE7U1PeKVQ85ufDZG6kae
olJTMp8NrDIjjdqpxHdwxi3VW/kRF1B7uiV9AtF85Be3TDwHJmlN/PC+8G4nOGhE
MGmXG0miLzSIMywatuqYo6EtoxYGsZoZ29OhW2JII/MsriJ6/eMVdOj3yrxRj1tN
uaJPrqFoj8Cg03fleuWggUpJh9A6jxnhJsds/qnsMaDw5ZtspZoLIbeNGCqF5Pty
w9utXy7PMd6bZSJ0g11PKKAe/H8ByuX7YVfUVS1VFy1TATIoKddfcajkYUKTtViS
QARN/WpI5bc/0JOlAdLqdoFBpngLofQ66EZ4f8kXKuknykJepvcxRHgN9zTfrVTw
dBuQOD5jxwwvz/HBkwBE3qTWw4XU1gHbZgY6Wv4WdskrkST953z/lJN9rUgg/V0N
vsVP+IEFO6DScvl+XnnGuvvEQWJpQDsf0p0RAOcmHx+7gJP+xwAR/el6dF4d51Gf
uZ4HxF+ssHJRT9aRMkrSmf3eFOXNLoE9SNQ4SyacUAApUZ4iqucuJkmjnXglkqRd
MzRtVGgZ+NVee4GohArtAMEnPZiMw0KBXn9PE3ahYuD56BDwMUEhDgf+VhcTQLTx
Qcgvq48WXe7yOvgf3Fi1MqsOoAzYYI8vtzIsHAABUghXDbBEU/rUXLI712alpB5s
wziFG3PaagPQzXeSnTEc2rOjL3gMoZCe6e0Xo0m1gHlU8niZ0O97mC98aCPlAsbf
9uGUA2Drn2mDPtB5QsdTMT89C4dyZTA5K49qxKo2VcjlwWx8EV8Embqq+iNtGqt7
hYwA/egtOfZYciYUo8/c+T7Ef0fArGwNQ+DRth+w3lwx60eFisWNvZzL94hHAOJr
vX+aSNgw4d2cLzyE8oUhQNYII2rPxl4Hc69epkrNEgnMdOf2u8cWG9UwcH4nDoyw
6UU0THOOFeV1kvkTMhSHscK3bOPIgklNgBdgSxeFOoAzTOAz9wkzBV6MKQGNoJA+
wWiI96Et9Gprmh/MIpTHkRLs8lvbHU5PGnWKDENJ5TGiFPGag/W4kjgAbXV/Dao1
Z3kbBXcVZO/3Ym5gxbZvRaz2AJ6pD/Ve4aZoTYjUXk/X9oOua+jZPSdrAlPJUMw9
AD7zjTp0b9VWwK9j9MTJFOO9eTQNLhsScbK5ANVinpfoy3GBjUYqFZrR+Jc+Akf6
U0byPgHgIvoOdclq3K6Wd6t7INv3ouK+CHi9Oc53PlzEWc52GhqnJi63ny3kiI8Q
ruCSy+qwLp8zPyFtL5eUsW6xv3lk2sJ/EUJ4H/Z+fFTHE9tCI6nK9V+XlKhDjn0u
pbAZe8f+klMYpz2MkzXIEFkkg1ora9vQfSAv2TMGtVKrmw4tk52cAjiTKeVLyhBv
nYab8GNB5pxgnCPC9o9pZmvTP6agHl7iKj5J4vd4wWQgtTZwHeEC+AnxepG2vEt4
uzYhu1zygTYjGzejlAjSqUMr8Iuun8sBewwko/lFOj/akjav0pyMDn8AZjfxw45v
ccmeFUHPX2T2GSq72LnsWSRQKqVsMA5Im7+VNGc316OWnaVS5TNpW8M4pyXBv99A
jG0tW/PkDr+gAuWoflfCCtSRCDExYHNAGFErrcqVXuOs2WaHz6QEQyXw1vn2mc5d
FezrYcJv7UNypnXMkU0hNcTAs8d5rgb/ErIEJeVkoO73onqASGm25HbTlYwkENol
7c5u7X+9VjUKHWcHGWu1Ibnalz0UU4g78hLeQpl6HAnsM/5i9bF8DNcXVZip+9pb
P8xMulc7P69o+tCcJ1JRt0mLoZTG3Z3UcQEAb2t/KaVAsBp/7i1PgIdP87RP+ncJ
yQPh/4g8q01kU2uhaWxPE0CLwK+0VgFcDbDcmmMKmOPYINR9gnRQ0xbxoKOcNaAj
QPZ0lyUp3K+A2d3/i/O1pVfzOU+HZPmdEM2RS0NA6bklKA69+rWRh/Hn4a9Sag5k
K3Md1BEK/TEusSMgHUKUwcsykeKCbVoGm6HLB/hBCwcJ4uA8yF0ZOVspPB+nzL1A
mi4nfIEnDPAtk6FYyjeULri2UOKGy53MpCJ8e/+dmlpUkvXhP3Zt6AqhGEjesIFQ
QvxGJvM4EFGt0cN7VFB5Dem7AqWYePIkwZChEjThEI5nDmwp/MwqQoYANug+GGR6
wuhFuq2XzoJOKHyGaHuLWvSLOXNjifjvSNgtYy1J/KEbR/LyYAGnr2+smBLLEQIU
2WPDF1v+YaEr/GyDWGSTgs2rWLhIPhHdKUtHxKpKJNtUbhA/DDNSs3dVkJ1HW87u
bYkGxYjOnOoxf1INrXJnDZb/C8hW7tLJFPRgI1Vc6YDpRn+4dN26UD5Vr4322uHo
vfwpi5T7nKAHa5n/U9I1lMVh8BqSlzZntCIaTSxkdM2jrEjPFv/yKFIoaDgpSV0X
3bE0mtmtBtFO+7NUlrkX4my/kmdZKg4KZgxk1e0N8KoMjYQq8fGcjfeczuEkDFL7
opLmnbID10ipSInaTg9PosBdRfLhH4dBIw2vRE41Vme+LY5m3RAT/IVpM6OvEM3j
L1d/SK5ZItpTsWgvvRxUvj30ipcHmqRb1rGB5ofIBqO+eh//5w3D5PWkK19Ivshd
FVOm7yotwQTmUU7spNrsAAh/PuxH76UqahY2UXp6eBMwvleLd8XdftzzOMVcvHhG
AeyVoVgQSEGRwCFPi2mTupyNonOIXFySBXHeCpdSHbEnlxDP/JH8Sw2etjWfGAJ5
bm66/nwMIRV870rakWOAYmyn9ebZWodOg7gEYZ6Y0kViBzAVKH0x5zouWJyZetgL
K9y2GXhcrzwev9pno5AodRbwkhUocf9jVsghlb7x4nssFPnOjbLjcbn/PbdAFY72
Y9EHu5/bfJPQ63urh3xtuSFZzE5VjWHwC0gfd+lhbpbBUxpOGSrUoAz7z0SlIIfv
pUpyIDYVUpyi6NzX1enPgUdF5DNlR3f8z3yqRC83pUvUgbCtgh/5QP3Y2hzqzgjI
ysQSklAMSiGbkpBDPZcIUtMyMHv5fE0LwX0DWlzZNIE9r9xyGSiOxDQW3CYmHt3E
GaqO00yi3TthEYgnOmBkPaZPgJQqnoTT6x11/KvhAJRZwIm3Miev2TqFugY4k/2D
Opf/Kw2tP4Gy8Uveg7x0l+lk0/B+FCn5u1DWbcepbQaUnI36Ui0Yle5LyJVmBtH9
zDciajIV9u/EI0TSIdMJXHMeXyqMnLcE7cOcXOnIMKFKzACRd76JPV+yUdUpNAXl
yRo/xja55bFqTMX9Ld7Q5P05MrmvVgAx9eJ7tQDBOGYzsNW1g5DHKveXrKx0zY6/
bLbZnHxNkyxhgXbR9s27cE5svsqUKt2ykZWgEyCl3ufJQzBLBO1Ef/u9LUaH0CoF
hnftMGFekyGgrREC05YdYtwtMQ1pvxxuxSZFT2rxGFdOBdU0qQ+FeezHiPJzMxRC
W3Smdwh9Xp0Jl23SZCjeLHhhsd6NFmQBWPLvZ39PKTX7NwxZzVTz4km7QeatIRI8
AeqGosPgCvUNP15WrTHwnj7xk03h6e5EMUSxTgCu2sqbxbrneRHwqaCeEZjfVMAD
x+QN7y7KmwwC8LOY1ZPPPZAMt3klzxbw8IRctT57DW1sFqC8uLWD9mxi2qE8Dt3I
dTrri1FKk3W18+3xOJ7VhI3bzuRFdjxWNJDaFQeSd2Uu49eFo/pn/vLk2nrPN3d2
/b/R8e/yEjlXwF9IVL7/kr4XszORMhJn4ZdgYMAftaaLTB5U5gmWzLcagzg5fe+3
C3UouE6+6nv6tMHWEMvzcW4MN1slNNhpb9S6oGuS4KrM1bbTzJcx6IY5+GOQ1G75
HmBY2Skz3n9/h4qTWmUbDv1Ws3lvHned9/mGsnm5HKEtp7SIX36JeMPIkzRxbPg5
PBDIZU7aMPdFzibzZ3HNw4Q0xuGZ+JaoOwJaYydCLgggS4c1WafymSV59y1NAi1a
l324ePdB303MLXOwfNzh2673TVNILIm4LbXcm44zDBz3sSaF31V7Fmq9BMhed8Ls
KvdYyFRNcjEWMceZjzVn7wbUlDsAXfLOKQ3s5GQ1AHhoqLz/ZHM0F+mW2vFF6r4u
es4j99qOXdwG3u4SprkkSu+FpGHvzDYonvUSqtT/NFUIO+2lxp2X19aB9zDWmS6/
ErthyKF9OlXO6pxmM/TBfNIrOb01voSgZjXtMaBjl7Go2RuJFsrOrcH7lT9BK/Yx
pG+kajCW+k5FnVJ8uLqt0rjU07Ol5yPu73hs4H8JoBhnUXS35q9h/Y10WFsD0Bn0
BUxyO0o7jfLoBa29A5vBBLO6WISFsN4H8GuMZ67b/52dBJYf5LyPOKI6Ab1BieQV
FZM0h04sGtckqCf0+03t5jjSgH+jN/B5cRdI0CYsmA9Gx6rpgBioVaIphUQL2LtL
vMiA0siNczPA8dXlQznAd6IH1zaJNjmUXxdwshTOpKpoWJo9MwlWKcGLz3yg5cJG
fBIYzss1gCHDePuHCkY5Q79c8cHIQsRRDai5J0K0fRO0DuocW1l11pDr4ajSRnA/
46Q/CTRh13JR/hWfZ/po9R3jnkuxafk9WIz2NYgsN4lUo71+jVSm6fHrlwHlXR+V
6KLpIazsTIDOLLzrb4DLN2dM9AEdKYN5/WZLC3/Z1nV88LsdVuqzW1lsex2UwiQn
4SlEiz2KboqIxzpkCHDR1o1D7Tzv8yByp9Mb0V/sX+yyN+PvTDhBgpbhFxgiGazV
Q/hmCtocshkOHVzCGUsI96kc3oypfo1uvsZupaLB9VPxmYVsmVOy+7LQP2TjN9mi
FIS2XAl38+N+ZR7vuOCVOgfjDjCxjsfAOsTpUe0ABXmXNHrfHcpZrk2aoPI2xvoz
6xIdiGixIAPjvb9sise8MHsd/mX+sFny6OyDz/AtH5qfBPC+qIjzJF/eMXmTvCbh
qVB+Peyd19JgUlCvLaN+u9OvTFWJvy5eK+OPCI1ftWtbYvC1pf6qEfIXyUv2N9uF
mRaeybPr8KaI4PfQ2jRRCsAjLHbwElVmW6e6nNaIf2smJiBflI06Gs4+erXB+4RF
vvvtmYm/8iqskILDnDWZzYHuNZgh/qqIUucbkeBKmafTNl+wQEoonZqoWnrR2vZu
z6k3fyjpHxbgrZab235N7tzBOGZQ6ASoNFXrIdu4V1BslqPffw00gP5yKoIFMKld
epB7rjSB96S6h4IG5xgrhItxX1CEeoXnJNY4R//UI6OwmABDr43esLJDgla3dPFU
6VU2FviQ6oAaWNZu1C2zdaisFJ6Zm2CKuN14RT4EocJlKKUXbSoEKcMcXeEcQmqM
JKAW03hB3ZZU1BHFmC4WuqTeTLS2AsXnRGrjQjVdFAFWZueBBYBh9awGWFFsW+/J
0Y3mjU2ejZtqTu7z0lGZwSm67//4gON4gkxv8ihC7L8EQ+eTfeg9ab8fwJQqC2Cf
8vdoi8+oPAVBGb8zjUdXfPr4vvVvnmq8AAEyPqbWJCeQVOnLFwckef1a3U1n/g6A
yYrs+Jdt3rSfh5cOP6qVWEbXRTK0yf3/XZJA+02Gfe9b+son0tInGrdrur2he9Lg
n/mTaKG10pVY9OYOHCQD+Mi7pnEcPVWFin5sTyaiVjsZQNRC2uWFk29bomdM8NQC
9dPyc+1fmuaqzhi10HQkMRXW/iDmy+iPed+Qf/cSXXCSjAqT/07Ant8fDE9R1RIw
F+D149aFEfTYOclaYbLFiwPGTKkv5ugKn7EC/+75IyB5JaWBVPqgiKRkmwzYzun+
tnr17RNtO7dS9Cw+OHLC9pF3grjCVJQAnGAO2x0R3QMYs+bgg1eTA742MZIgAL8C
3MrOuTfzBsQqQfu3opHccocTlLOis6ZGqbRwFdwE/Ug2aYvh6hdsgsMYKeA8l1q5
i8Ql27WQcMEGEeihuUENHJB90wmZ6vez8utXjImC9MiPyyuZOTig5Ln8l5ZSatjG
VO9+MMGKVgCUrvnRswsTSqlNF4moqrXrV+Ba+I+34gIjzfNIkBs74YGdVG0ApNVh
RdzA3/1hUcBbOFD4Iv8OwcKO9aUnzxDy+Nh7w0baxq+d5Ic+sYg27aHtERgVfDqG
RwoOs/5sh2NuZ5CLYyQnln/C6JrObvW/H5swtkxnfo7pxbJc3fF2RMAAz06u5o97
WmfECY92UJhOXGEysxH+WLeRqXkeEbTc4lsMJzUYrJskrjCQv5X41hEUaviXbFXm
6JdYyGNfgZwuUKsx5WXaJHn/eUtzR3ht4wOT7mWQEpr05E7z2KBka39JILP4Hd7T
D0C7QaJ+O+P+P/Wmk6Xko+yEfjRIT3hAhL5qJO45Q4EkRjbATqvVtpPF3CDLK9kw
5iBJ9Um/4KJ3WDNfF0QDlVjVjNY8RvH7a+orplrqjR+R1aOOSA3rpt5DUvrxcMpG
F7G/KHtu8WstW+XUf3XTvvbeFtO/UpS5uogRuPzQ6JnyRX+g931T607SMkc/27Gw
+85LiVUq6huAAnF6263CqJMIjK8yIMryF92qOs4XAyvRBUqDSlZr4QtXsyWeN/u2
qvZN9hqVpcEMu66MpdH1158kNmHyQXMKWAi/rfmHqd6MKHR/NZtmy0YRMNDbvl9D
xyZjuweAyGirxQC8vv/s70kwcgAvd55ST5ZiXqsDT/XjZvHL2Qh8paoXRRe5srVq
zRCYlAGXfIkQq7dZPoC3yzxTk4SJmHzC2+PXzf6JeloYh6PZ9wzdhRbFp2Q3r7Lo
SC3/21gWq1peI6+gmK6xExabwx0d6o1f+hG3+vCiT5D1JFxmBqGDA0/SVuzZnVCP
FoJ5KJGcF4dwQaRaqq3P42iTVqKHDT7DjSglRSIqwx3HPujKaRhFh6tX6L3caEp3
8GemB/ORFAxLbfE53mOPo5Pz8OvamDrXFiuqoflTSlvMVrgrShfpJgFP5jTPNkIE
8CSIMgAAP7PZvIErg5M3FPq1o81CqAdCNttGGmqi7Jit2eWj/mOI/FgSEHmcHepN
fzLz4/rqf9Hju6eMjrTOVL+tcrpJBPwLj1kA6aNCfy5WZoWKBknn/LmMd8pWFf5I
YWPFlJXjS7sXPwb99oT2eptxNDSwRdlgpIoElIn/8KY/E5CPRB0gU3x0m6TzzBw8
O0fgQDi45BDy3Tq5kudfzROi9DBcnQjeTQlUM4hU+eCbRgLN1CXvkVI4oKNlvqbl
L8pCwHPdBpmdc4avnMn099iijIlDoDr3KaL4ZsBy+z/rOF/zzfCm3bRA2Y4bF9T1
dyG0W8KqoomGqQb8MmwvURfrCQTSwb9pp5wsMzqOOkfeE3kLmi4pgHayTkcCxA+5
pj4foWACDn0G5l9wKEmp+K37EdvcHhD47XcdpBhGQeGY0fxHbKhDiYvq9xVbhrR1
BfrLnYG5c90UBNlSB5M8c1AMrgP8N1raMw1DA8oGtA67/bNbzUeWShMTATvQvTN6
v9uwmdmCtou09XbgXkiAIAVq6wod/imOvqimbgfUiR6hY9cyotv23dxinpyGdhBv
a/Aq1nQoUnkaJ9wdCVgOv37c6IoeeMnx27YFSufP3aSp3MAVRA23bdJrf66khJ65
Ule4czuqIPx6hV/MEM5Ku+Ptw5wjONafkGg4dDAhzJlp3y73O5lsS0fq2jnYh658
iGnwb380u4x0MsNGHbTVNneNZMuSK9MaXBdKIsRmGQuYQq3PAsGVslqH2+B0u1x5
OurkQxGsBs8wb1oO2Gir1dTmeG0Uv1tHHdSOyQIj6LLhQgPg4h7ijLi7KYrIcU7r
LobjW7LpOR771sSqq/sybwf/jGqM5+6lFOcVg565RkWS+cSGPbKOapxrqS5po8PJ
zXC0UajsJroC8wYjhkxL9XXpIrL2n6Jlwk2JPkkxn4g7SO1VDHCNckk1BpCZfK/l
aZh1cQDQkxG8CXHzQZIfKioju1jQobUEUuAFh6UN+3Dbx2sIR1R4v19jg3sn3ymQ
z1gZPsD5ttbAF7kI4PZpUUYjuTHeuM715c700fH0zHLsLGTbRABDKR/WkRdGza1J
E1yIK2Qi1vArX3ikk0tOSo5s3Kb479Sgtltw++XDN9nog7Hk3rararNsk7ed+YH9
vLSQz8MtZGJd0+4fyse3LHuIT+s/Hsplb+sydFx+0pEhTEunV+89Uf46+nffdOdZ
JUV5cyJNdAsE++vEnrsQIaZgJ7W1t0N93L3MAXvBPYCzljzsLOe/ya8h4T77gOmS
dXBOEjaQNcZ4FnPaHzF4k9sOdqntGQRTyb/dPnU8pGUrlr0VwBqUSw58TYNeShrj
wlnA6bLi16HgYPGcHK7zfTJ5qz0cWZm4NDwo+omCMorfRZFkKBX16JxYp9DbKFAI
9ECNR2E2TRX/nSkn79FtGLa+BYG3zavGnfMcYigk//FN/pWTVcKTOr7s6eJYpQwZ
TmRawI0nH2Cjb8PX53JievElp5PwVx8DPAisrT+ysjNo2zwGZvQSM8QYnlsZ3xGG
vY+euz8iSu42x/76OAXAS6CAU95pB9eyY4aM3hy+4BPVblARbr4E3ZaxaUr+HMCD
XdXmC0K6XXXkvk78SQDk3l3s95LJPOnIJ3mrL57/vfICM+U5Fkqp5QiUcKvMLmo7
6YKwEXX0j9XIU7w6qhZVKppZxHYCoKgkD87oCKYhOAKoCB/HUSMZapaiJBCwttfO
NtROd7L+Y6A19Rdrg90EIdUxpjeUs2sXhCSPB8xL0W+EBUhwbIiiVuYtU2dixxM5
+GE/lqyEhX2mnCPx0Y+FJ6mKCKSSMPBZKC8+xllq7P9JLpoGOmwK0DfCjoLabuEw
lQGtFF7xuG9voquXjicJhdmZu1J6SkQUEF5RjmDAzCMsJRq24WQUm+djUO18L+rV
504Yph0zIT0T6X8fIenRC/0j8YoidqJWA86nqxWqnNvyf2dVPW8ttqyNBLsUKT9D
EnLCUCsR/vK3pMJi0BGgOJzPaNQln9s2SWHo9A1vD/Er0nB0f2P9xA/BZXgZ0q/n
k7rgT3hBT+zvw7Q1M+v/n5wB49leeWepq0MFIIJZJ+V8GEIkNc3VjrjZPYO1D75r
vfVzMzndQByE1EtyuK79Gum7J+aqkfC4QAQXdrDIRAe+5piWKvlS+SeNLM1osy0W
11cQQ4QkmniD07BZ0BT7D5JSMlzESiOSVIe/TIspWTgvrcc5zAuzzyhtqk/t5IjR
Z8BKQz1eF0EnwxaJ4/rOxog7dJ7wrnv6F+tsMxu6LOKlx/neP5qElf+iqNp85nCm
qBGzzSiFkchp4N2TVSYZ2EiQrJ8XUUo5f+gPDQhN5Xxm83MhzKYR1nbkDY7XgzPu
jFHzg6zDvKaNFwNwlOi18XfOSwIjoW9UzJcWDeHcttGOyOi/GMzyrtcXk85ovvXX
kRvF7YHxVfwd3tF+sE7+FCzd3f3jY1XKc0y6D+MVEDjxVpzz2vXKIdUJT5WI3N9w
Txe/azKXd6+MazhpV+sQ0A9raLfncz9UvCQ0gP8Qgj5w/diUSTDLbYf3IHJSecko
JtYW2kWMrxvyCAeXe0rO4Czf/K7AoG+XtiX0JQuSVw0ooEQdfTmWcYsBk81V1BFG
ln/2B+f58zxrW07oIuPjT54zzYm/QuFVws21i+wXlLz375fJ0aAT72jEsGR0p/P1
EOj6vfwLrMYSRsvlMq/B5c+Oc05QA2DrXceI0h9Yo+Jwtp1i8nVaWh7a1ViZPfFT
/gPPxLSLpQ5gpSzQ6/IfOPKh2pUP1czBhptiJiTUDqlAI6zM7o/LS7usUf4LpMbj
SOknKFW5kZjijtDwm7vx5Z/sbxjkmy1dEPAshH12Zbnt3+Ju8NMMdQnbMmUBLeVq
zN07CQXQwCeSBx+Am+klTmX5esp9PHXsW8eRTaOap8lFUTnjJLzpv4+nVfwz9Eht
XjY7Nd/Z9lzWa9FGw4KVveuggvCy1mbBgtC/TB/hpbwC2V6kMynvBU+TD1mdLHHY
5ApRPyI4VODTpSReOHmvPgRYE01lEXi+GrvVF4dXir27DHQjays/G+8QUxVHlBbM
f6eMICJrQTlbVzTQ/guAuM7qdr5mMEd7DrocCZWTL5TAuwytyN6+0qRDgOxk+8OP
vifgh4mh3WkMPe11G9sRu1TovBQBnnIxIAsAjg4N+dltIbBO1MpujizGUMtV5XAC
tjM5DkXUGiFpiMAkibKf8TosTIEZmcsfmZ7df/MJcFl8sGnMtGULzbHUBj5okfnK
QqZkGtx2Lt/ko46pioIHbDOONg3AtAfiRnJxAdJNSuYssqno1SS2UoBWGnB1cHzT
AjLah38xnUxk0iGIMH8CPLPgj3KnpsPpUKtKGVEfIpcujutXp4Eu9trYb50LE5gi
SvNVEXTUq7zx23WFVPzFrpA1hhzXtjS8QK5OAuA8EfYsYA84yyWD7y230C/PCGdJ
mXEfFGrxqEyvQJJeEq3QHouvV3SWgVxZvC6Kp6YTq9NwlP9CvXRzh0s0J/OHd8wr
6QGZHGVhPxlCb85Ced6chCgjABh1K0kyxK4SzD5hVqdwRNeS4ddy7ynuPYZMPl1z
fiyKawP+mpvlNeyyhfAdconwnbocYz9BCXyuOGVgJFZEVhrD8Rf7whMgL847hDaG
A1HY1PN/uf9z1K3T5ZnP3UE+V3T0pBxErKObo9dnZjTYKbNCE69myhHmHlp2rykr
KIAC0T9H5rSVoFMkY2/nStRUytdmQgKjp2vnQgbw4Yq7AVarYxuyM7Fw2f01GSZK
BJ/eafFv8kVhCiT21cDLoHf7g7jhuoaPX61SlUvIVHZN4dyGmthYp4hdV9rw4tzk
ZbMXs/S4FnuBKm+uY3zuhALLukVyc8cnzRGrFJyU6d1W/W7nV+0aiYgmw5a0wM5T
6p5r1BgV1pQG3xHHRLEgGDgpXv3Ci97aVwV8k0V6T5klqFztvcNW+B1xw/vThani
cBxSS7JTwZURjVpNaFulLHXijBQMJUVSX7fANZFoY14BJZ0xpi0UynAFQtAzvUPt
nk8qQMMkgY+je7L8O0UtxWVGrUIo2YskR91Za6gr0GNmNTLe/vas+NIXONSZulXM
z5Derb6Sq5GBwsDPPs6fPdswvzPavn9wet7h5jhR51ty4O1iDxu05wIvb/bKZwlP
afcN9CQLZyjeRwTaLkv3a/0K5tgW6dGNKfR+4NID01ErmytcVHngFjJoM9c5JnMw
01EnSNYtNejdejCFt7IPfpObaXVHvI5hQPj4XSlvjrc4K6yFggmmu8YCwJIvGUjD
EoZvxlXKGjEmyd5whulCrLHhBkTw52wtwCiqfVaJfSsweDuRibjAsfyjxBVH4+53
uwnYeF9lLwj4BBze9AhM3f6Bg8QT+uDyaeM3q3xBgmY/M+KCGkwya/le96jrb+6u
/LVBJysD5lygJ+vrvLtECK1i8I/59+WdGyZIbCvZ2oTVMlSctOVO2FoSg7W9GiWK
kCK4z7AwZPK2OQuk8qkVs7rAlY9sCv0Lrk8IDxJH0oSmCAGuyBUYJuYvlLsi8704
F3GjAD2lfD9hwa02YdGu5bDL4dWknNzDwWQGJyMC/AQA7CZ1Cz765CmW8RilpC2q
coL+AK0kHsviy/YFx3BbwV/SCQjTVlgIaWLEYu0+uDn6ohcx7L8wUzB6dVaj+kUM
7Y+AaWycBBGVWo6bt7Nsob5envF1ogY2q5hCfTm+nvh77jfZWd0LLfC/qWJRN/6e
zbOu6UN2BozBijtOrBxLsfra4r4Oxx9Xt3nEHNXcyv1cxeOHO00BJj8zos9Era5T
rQBeVzZ068AxH/6T7u3X+mWjsO+xx75TIPcQsjEuFm0HL/GQ22YLkjSholPTbFpD
AnJ4Y3rh/+8K9NNESjl3Pb9q2a1vCCfnYxvuKdeqqihdZOKG+L2TQ5KbDBMWbv2m
yEkx2S+X5mlNNd4ugubAXt64Y5p43U9M4JvIZbzKtDVtabv4FkwDV/jWV8d10Nco
YJa/fe8NymwbtfgnTrwxPPIs9SO51lIGPx+mB57MuwNO6pdS5lURlljVq3cisuLf
Uq9ZXalvjdMP2nGiX7+3PSgXipTzXOGKnY4vKGPgBW7f/DUpqmP1prEsf/XQO0VC
nxOX6lMzqfnmwzB6vksTp0SXIMs/eyInDXql5ZBYyNFF5EDtwFpH1rPNC+oMe70d
QbYquSRKlqeN/WU1xzBK/TuMJ1wA1LelAS9ikblvnNbaBYQO5ghjRr+pp4uZg+ZE
ltCfzJJm21Uw6qi2bSEo9Xn93YSFHVjiT7Fs/f02zsEy1fzFRuGMKoqpdvvcU+uU
G6RqcBadx/ZRMa6OHK7xqTE3FEN+a+UfVPUXY8xIpff055f5i6MXu2vAB+2WAXE/
XgNauyWHtBouaIpehCTNKPg4nrv9rT4d4F+aMUG/R516kqVi11o2gBEQL5PqxSnQ
7zckI1C+VHkz83tjdfiMeGY9uH/5e/yCuEq3fw2VJTR5NJFzLSdJvEJFqmuzY6VZ
wYFpIr5E5Md93MFdQCuGHVaAw+itNzspKTzQ/x0jWJYye2+EIHN2Etbq8phoGlwU
7gC6gFlnwBN4woVBw+ZXBnVdG8j1DY+Ob9GK4H3WqMzLu9LuA//O/84AmCQfwcBr
aqtou5no63xT6oNhuLuro6OEXBMyXlkOCL5yQdBqiTIKYZ9YngZFR37dLcKWacZJ
JxruqtcjdBvWyofuodvYABhHmbZ1lWPsBQpJ5nl8DtzGgowc8v3h5B9pyXuJA/rf
A4BVxfL98sImTc8N7zes9Jb3fJuYoIrXv4RuZAa7iuoFoLpvgvH1fGPphtrAWxPx
b2fE8qbeF21sBoxhqiEtNM7+GiKbnzJ/2u4ZZ/NtilELQiTbK7w8tT6MdqWH6gv9
rBplv9LW9/HbjEYSPGS23e7PqSalSHInBmRFTsxY8qcEFnyRO5vau98LWys9Khux
JnHar+QWlxm9WOR90+qNGV2LP0OzR7tvkvA5/A+8ZT5VcuyQX7wUhV7FNxBo2AqG
ubCgoI6Nhh2og0Q9YSVI4bWOcTSMnbG3Cf73G/wbPRyMsDPRy/7aRJ/MBb0nEFUW
9uBzVPcYVYJs8RuKtSGeMYqwjiRN0nON8Y3JLvwpgrMDrFFZKcaymEmIhgmvpjWA
fjKoA4QwQl8GpCrkylyrZ7tKbAH5enRicPAm1kvVHJQ8IxWwqtWpyUCxM6eso1EC
VpoVyz3bJbl0a75sJuzcDI46xxmi4QZS+NCdbbK4DQGVaR+4z0BMp7BUYFd6QTaN
0mwfbiTwc7E9TyAlL1RMnU+rZRae/73x73//3VI1C74MaYUflgXYovoKs7RJ3eCx
h1LT5mLS3LTJ65o/3V4AVqXfM9UarcwsCC7yezgJ0Tj4YYK5W2vHpAjNWRw57xVl
d+zvave16YBDeb/kGQKWacX3GPFO4j1/F/a/Kb9l5qO+rcOF/sGR5n6hXA3vSh/p
q1WDfsFn/55sndtk+pJy/9JLjoo52PbVWSZXg61cpE++Nlycqb57Xk6F6f8L7CVP
Cg9q5sVDLax9SgC/tMZus7eC+BMp9XgAEZClBxdlPkOi8u+X/f7Rf02fQ1YZI30P
VHqSkbp6+EjQ8q50pSsEdXY0iu5f2yYr1Pb7h1YZ4qvsTprYQcIsqQaEBCy8TREH
Y8WVYAi41FKZPtLELIClVoXKD++Exj8M+RL1qJwU5xaMqd7pqbXN1cZa5X0oHGbD
av0wRfHkgKdUHnzS9tOKcCe0bul+5O4a9rVPZciad6fOLbJazI/usd0N1sIZJd5W
XbuZLwIhuC6lqKzSmfn0RwsSWIO2iB0WUj0/iN6qQJ0td/JAPzjSdl+izYAJ9mUo
hQW2imqNwMp4CnRih8HSvfG4+EF2sTj+BCKvH5ULM6ZhyFGunnYzNXeL5rbkHtfI
OQbJNU5sASg63r0Ke779qsa+6eG4+EK5EwmXhLBaVEYBKiVSigv8XD16WHLWLfiS
ykS8X3cfmPGqmSkHKv8TvrwLPD32AGrgBaU/eN+DQgWCuGMYt8pKnXY2aqsPm3LJ
AXy8q5pvIfVJ/ci0uxJQKrtWuLufwLSJwGsw2tRTG1xbt+TALHv7tw7butWITy8n
OB2ImCw2Xzg9DM/LF5tOr0TLv79pDi8yJDzrK2ukvETBhJfBKPChqFy7wL123uNr
oiaOxrBei2mJLX/02tLbuRWY+qMH3iCFjGUf2dfA0IEjdMqQ1SHL2hgYU5lWSmsj
cM6Cr0Fs1ukvIuNqbP5S2IIaIkbqStt2zdvfgXcjHGxhHwllrPLXrF1HmNtz7XgT
mAwdL2BihuFwSvUeCvO5daeOFgt4Tg2g5AvIXu18y4XaMhA0eye4Bc/a9dIto+lz
k4K0n0JXCWxWALwhazCW2UOosFTnA8QiQKNgG9ooOviWuyflP4SBl1iQFLyEv6P+
si226KU7CVUlGFR5WJhj5nbKMP/vWk6XBc+6KioHdR8FUYwxsOzHbHjS90ctkvra
OE2FQHhMt8WXE07eDs6jBMw1ALcl1sqiw4wsQny4Vs45tcPVogO+yKV5KNb387KA
17I+ZCr1/b2d0ZXZ/MaLwSu6lLSEJ1Xp3cQmp3fkuIL+0nDZ8QOumVWQQ/jONB9a
hBr4QKAVA5JBdHL8bczhPHYwjEPaerz5vx67aiPuCp1sZebjBC3jteSGVk5W3SHp
6Pz+LbYECJa9vjOcvWkpbfY31bLUxofe/Ep5Z51IAYqSBBpEAkbdmTlFHQ02VaTq
4vJ+qrIFQDhQBBd3ljkZNp4UyildRXYzQzTJZ4got2ridruiHnhoIQdOiZ2h20PY
aKXTDM4fibNg67w1P1AS/Y3gXaCC5dvFg6C0i+bXsrGmmlM664pw6aGDP+4vUxtQ
QoMzfyRA4LDgI7uQXC5HbSnF3zrkob/JOqT+yGEhEvDW94Np4I07co21uEuk8tm8
KpDW0R97FBPCrGskHa0mI9mHEAYZtLEdcGCuImnU7v+37Jvrj/VHF0KrM+5Uct8t
DYjisYqfP5uOb5KSF/etSk2ESB5xJIBW7MznRLhayol+HJZKcERX2y7L/ZC/hEkl
dANuL0z9YB9eF2QdjUkVfeIZ3/jIuVhjsMU678kewUshy+kEd7JgamKnhHMPlqai
1Uy4stnaersRPiJk/fV2vKI0benCOufOv3SignP0LGBAMr9YcabRSyU6WlDCJXrp
VsMNQfDcpQ5sVbYLv3zGthYoixhA91AG//ci9FjsIqVKWdT8oEVGisJkLqAjJvxb
WeSkzXyJYtfXT3A5ozE1cW/aAl8n8RhQLSq+Gb/r77AciLPNf5V3oiQpB39a4+pO
8m7/zw2u1C8z1tY0lt4TcN77BS/FNHIxpGHj0WhZDfMd0rXOL4911/SVkcR84X4f
6JyHioZrykwObodw+uV0URmNF43oCZx2eOQfhrLoGbRjpzYAPKXHX/RPTlQzabUL
OYxwR02AswEbpm+dsTBq1/qN8IMwrIdOrUjOrbodZ9rYakk155OXElPsnEg70zGa
t0RQcqqIzj3qxJVigRqAtbNEzcgmS10gu4TDqa1AgVesKs8Nm1W+i5XqZMn3pLu1
QUgNp8Kl7119KK/3yNm3m6IbRFGzCqpl7NA+A/gzXlO2p5zeNUINbpbnY929PKdC
BXlBTFS/q3Icq3ZBwE3lyo53PPrDWtYqqIP+h7lADc5sH1bXObPM8L9yeV8lFTVe
bI+R0pJb0NSXt9WOU4fstQt5Yk70DkPQ6/oLEJS5iTPazNZNqS6rV5l1+OdiDsMJ
iIlI3wAXIctLrP6RV/PtsBN7uGHjmK1a7BuvMzWfxfNRare0bk0iVHAYq3I5X18p
Nbymo2frtF9Y2TLvvc71npwDWybmIK2s+GZDuZTWfsH9IPfInAnzVuDSGsKatZZP
9cvV4xQl5Z3WG72nsK6rlus9QGQPJVY0I1q3FejMNMPimu4YXuJj7mR1UjJDqfKC
TlQ+woqKlMdll3ABgOLO78hH2xJHSXfkS3Ns3TWiAXLpAoee5d9iqYneK1GRR7My
Pd6qB6TQubHR6IPnptwDnr1EqPKggi7WPxjj8mdfCPXXr43cHv9Nya3f/NZJUUKf
r4DIWZm0411s9JXLbBRVU9lw7fxhIxXhmBX1V7Sw4w5dbyStiWdSg6KueF5sI6z6
GxXaEZ7msClK9nA64jBS8MYbqXrvMi4KUP7jHYrIou3pYp3zYs9REV0UFhaKNACB
f0MrhefFrrd97+4usJPZTP+pHiay4rsaSdU+WfKpQEN6wP5/7lDGyMPFQ3h9rQGA
pjppiXdwL0OyrcFMhp5HVrLkbbn0JwazNGecO/PL7s2AFujmf6ydVhkuHy8qMSCA
LlUbWCLHymF6iQlNX+9KYucLOzkTR3yqG7ZD7MqB+l1L5I7rhlxXMgM0MDdFiMb4
GQEEaQOKcdMYCuS/EJamZ+f/j9YIlb7apyLKONcekvdwx+nADlD8QVrS1YhevV/4
uBbqqvvZVO0ztQXdEdsyJLz9AGelEsHjYO/uOoxqi47XfJ/UaA5F8gxpTfLbRA47
vvIU4a9YSL0IDaQ7+JyChpz5Qcz2tXBd0BS8R3X6iLkmu+RSDvGoebHlgYEpv5+a
WuUg0CFFuhY3QMx0jGm/r7HKd3Eub6wbVCmwWGOTehqX63jeupM69iCSQbIBiRTi
ILgJ6phV27ZkgVwpT34jG9jQGzxi62q+kWqZo/lMmJu9pElyYhZrJbCJJkotBEU7
y6dduDVQPEDsmdyaOomAdHYs5/is0lUEHpi7f6zc26ixvs0H1DjtoEkLa5cvVZZD
YpID0f3/7kEBwX8Le7LbfbeRLOazrvTWdhq01kiQjhyUs6FPUFZDF8oE7sRpc8KO
A6+Hwl1/FdVYmZnCzhuP0X4HUi9l7MyL+aDGxPVFy3Orlb66BRQq3YN55oSTnisk
T1xTY1FSYM+gmlagz3xlPqb1sqXd8LLz39qDxgeKYsxiMl0iFKXBNM7MV76bSXCv
5tetK0Bh8cSUS7pT328Qpvy1D3F54JtBHVXOgXiW8yn1N/b8eK57aT8dxULDz8dJ
nR+GE/1kgTlAS5QSUvPiKG5FxBUEkxApnGVHg6UzTxSN+JQyeVngxoLUX9SdonkE
BVaORZeuCYDi3h6vRUicj90kiZRiFyZyKyUwrtLpxg/iNgbicM8UMJZythvV4sdr
uYSme44vB7LumuuDSah1wzv2gYXq68SsJyNF5DwI5ssk5+lMF3Fb+Iks9wDhGar/
6njiHVHfQ/ajHrQRVe8km2ruCipdgjJW67+yGvZaQV/0nJ66TchI/vrARtbuPT0P
uXu+1FU2EHVEcq6N03fYPW+2bKs6Rva33boaOHvEwZC408DRm5/9dcxF43dUKj7O
Fu0dup1nXQLEPU6LinoEC932jklk8jXE9w9AxkXaCaFQgtS7QMvXAyA0QnxzalmK
jBjmEjHauM8ymxCyNQaFryOoW3xcdXQh09YbOSeVVbIg8PJipfK9HnMmDt/qjWXb
FY8ew/m1YxJpQFse/+EjweH+UDEm3lij+V2gXmStEgcvbYMdVuOykvkgIs99W8I8
YLB1IW2V5LNwwixsfmyvBuhwO5RO3U/5mcrQzIKq1q1lgpRNz7HEtPgyuDlanBX5
FqKPTxP+ZxEI/CH1GL3GGFU5fx5Lu8ZvSMY+sFu9Xodqckwly9+dFigqNgLvjSid
VtxP+LwJjbV3O4z39Kjaloi9gOLR3GZCmm5hU1vMeakt6JXULl8JwWED5zUD8ZfD
rj5GKqMA2zQtbhT0TaVw7sORduFJ1xnLk//MowUOlVF3r1Gd/awnUlEOspTjQcjd
bpBmRHVi0Ig/6aT4hZ39AG9liJ0PQ/GaBoFMBn6BwjGtFWyiiZXpQ5NZwL0Cy4FB
omjFLBAhXU0m1qjSloTDb6xuxuI/9RXQn2GVIyGaxaRKnOTWoVNDPdkRFPFnumr4
ccWRC5GtHVeclvCLWaYHNWjdvTNXm/tYvZXLYK+x/wco2xzR8tFoFE037MG02jZX
iYSexYQLO6rQ2p54lKAK9ESbMM7KWdho5rI6AAvq2jDfENx45GuB2BUO57LJqAu+
tEDvQIGqylg9X/H+PG4RQhYtixWbx9xFEN5A6F9VSrJP9/CF70CZnHKaRU4QuJPx
jyBRDF7eg0JJWF6PqNljf3GC0wV6ot7qCenCnZphFuYn1ygvJn9ZAyzhHu/2rLwG
f2FYM9JTNp/KCEk1k0fQu5/KS43U5zh93dBoNHosExv2y+dApHloLyjkF0qdGpFf
9mhQphY6/DXn3+9njgaQnqIEPpdihGdAI4d/k5YCBoGLQrIjs/YyVNrL9djw8Esb
gelC6V5iuSjHDURTU8EaxoKB3Zt6FO2gnWWRRyB0wbK1LCXVNKb8/txMhXE7C57n
m/CAQs6NWyrbap1mc035AcxHlbzlhODpUCgLpaA+RRDYkHyM9TBklN6eG/sf6aWN
w27F0Kr6QKhJmKlgqSVvYfFvj/zSY2b8p8XrmdF5ChNmFpquWlh2S8A6Cxka3/Rt
o6ATif8TLIl9sOtM5kbPs5lbIAPfiIY1ls/T064gD6Ht6WxdXt3+TY+U5Xc99W97
8B3MOEIhLHGo3Jwu+zubax1DcWXGcnJQADVu/Ss/Yg637KpN6D8GdDxh5E3lwXrS
5NR8yFacoYrXfah81QUibC2Gtk6cXkqx5HTTYLd6dTQaBNfWhcbiV555eWblrsLg
tgEKBLjKSeFng8LinP1gneZ9aexA1qdMGrE9sfHUfYdsmyJl86Mt6TSzvByE1lgR
SZvUCP6UwNjC0inOL6M+3Gp5ry8L1/83dKxmYy/BScUvsHDiIInA3c0v3qaS+hwT
4/Zur4QWGk6svAonn/Is3sK+fdWV+XPNIeSjt+T/iuRHK/5iq1po17ugDmB6ukTE
bK5wRU1Z0sFUumJig+w/6RevG0OOE0TbXJEDkblNNMT7SvHCnkAceR0l4F2TNN0r
oXfBoGWvmJ7Z/+Y1rLyxTCHw1M/9ai8m6n+JNxoNPrk/W/kKJP/pjbzNK0XrVmpd
u37AFj9IPjlSY/RresBPGRU91XuvXG+LYxcboyx+9hPHe1LixS/scRmRphmLhdV9
k8hLK17kJsUbOk8T9v2rsF6OhqikrePy3IT5bVE3PFXBkBvmJqKkxPO0gYJxjLzB
E+LYWhgRxBtFc2hhTdu+uTW8Jez1n6xLPdNfjs6KWaMeKEk9XXE1lvP8P1CZ+PLJ
FqDmJlqPrXMoUaL+KE2AsqAgs+1uUtfPoqZiV7EAV+EjdhZ4BHqmuB+3Ly4T/XYj
xUpb4jskq1NRX3t++EhQLh8OuwbjPxhDTf5kTQd4Px+xCORN32rgO+svRdgoEmlp
u03gU3G3UfFJggmIzEcK4aBKr8TD1QZGT38XKQMQN9Jo3lva91CixNBWszoSj5Cf
mYjsfcrNKKiOzKg6+CTtuVgfp5vqYN8KKyvN7tw+lLRQWbTyP524E9lUrfIHd992
Phv1mmcEX6ETt/thC32bhH0gk+dRoxK+/FJ6dRGCJfS2rRJ1dcPJ560nli/wDFaT
QQxwtg+DK0WvcWf/4vXFFtMs/pWOFpnqxqy+C0BlFVJ0V+Ag+D5GejXnqxrVbhLO
YoE62Y0cQ4qsqET1RERROuhq4qjA2+UIyY2rkYPtIu4C6Y9NoUjGibRgsfjnlccA
dbMQudxl52txo3BVvIxaFoX+D6ptnXGm0Vz7nrOfc0JbLh1l+pGzNjuhpUPsjtKO
l8nF6qLVI9iN8o9/eYKWZ/fpssQn+JAtpt7GRsQI8lTlesphlTRz0LjTqMdc+yvW
FTQJXg3IjEHTY3eWSFtK07Kszebc+Rz0UdJ/lIitEXfDVfzi3E2rdf4Y6Orcle1D
rQrfohmoFiSJrRzzEA+P/p21HZSXwq3FhAajTifGbvu21IEFdOKNZvh+AmRDugbn
ObbJGkm0nnSxKPzYd9JngiPOeKDNAOP5GC2LXbca6sHEd/tdxKpr2yS4Ne3tYJ87
Z0GVKNCrUTk+fyh+mxx7YhgskpvW5WI2cLT/v6YPftHSzGR/LShNFMHsOjHII7+4
ylubdTCTgQBs6XPTA/Sh9zpHu7FyC/620CVmQJq35Xbp/ZHAwPKmbKtAkcG1iz+X
7wpVrXxYPTgnLK2/1vEGUKNYtzbUVYRa1kYlejGm7n866tp1Ff8dK9A42mYcY137
vNHuct6LHF9UT1TCqc6/rloPD8BDZMC7fB8H6I+4jOh6fe+PvegEt1SwFnwGnWwG
yL51TtMbp78lx7vXs942inyobw12CtBA0By/EfXDT6oJYcRGA0prDTZrG+CgY4N0
JPCw1DJzZdnmwjdpipTDSLBdfq7nc+uNB2d8pbIq1grRWe6ipjj/pHu7zOFdevI3
2nAn0fOMFbvuKYoP36wCSp1Alg5iXtqp4WbO6ELN6TUi9qllX4wLZ1KAgoTDCuJK
l00AHprLWwB1CofI+0ykrhoLQlmwm4WTOhmXiZ9Aoyt7SFovsqw/qgoVzqIvI7dN
D7V3XqEmIXc6bgX80SJbirANzEQJFohQXF2kSJm44qVwJ2tbi7eRcmvxmZx8Yxb6
55pPzx0G1wvJ1A0DKnlcRhvBP8VmyhTj0oIFPg4M0HHNrMpf10G1xTS0S9WdFCR9
MPEACdjlZQeZnQEvgD3OGOBLv+8CJ69kVTZ4zfX0z+A5vJYixFOtm8lUnKamSGqQ
FWhOqsM7bGyXEAl/RG1uw1wHQ4yeWIpC7+dy20ES5ddeqy0i0ATXghNslRxcQ5XX
Mpf8oxeWWhBTJmZMMAFdIx9Z+xwViezZ1V8VvHoEnBYMPZ8O5O8SmJRAahu5J3S+
mGSk+Q2q0kDOquc2X1w71WyDX/ubVCCMRYHFWxNpqUHCSB7gw7Of10t+ugM8Wi+Y
zjxCGD6uOu59cqTpF7lAOwR+bKImb7WouN0Zsi6kFRsdV6GHNpxtJr5reLgkm2Tl
t9H/cOZKBDSC/oEye7tPSLXNKIwKcxFaT43n66IGiLA10nxZ9n7YBpHtKaJaBYGo
fYteYAQ4T+ah2Xd8JRjlftjwSeQ3oSqTOhx7AxM2mX0UvPB7GtOOOpiYANgrBrYT
dZoRt2L1IFh2QF9YseYz3r2eKfAdFsYHX+yuH3U1Pbw8jX8CB2LdO9g0PPV3b6jh
EKhijcMlsZddvCztnOSMbM7upmsnnFH3dVu2Rnwkzm4nonxY/qoKdbdQUQXINAQK
Sojkasu8SsmQHnITty1/onhn+4Fk1KlyigS7PgeMhx8IG7uRQ2e/P2UiHqGmWA/F
9wUH7XsaENeHdxnhZ366X6mMxv3VwjdU7KXpOxv9pMHagTSYqCusPOAILWF9ZsK7
NzZwNX1kVBMXqJzCRW4xjCzJKPPssKZb7UZRZ5ZtMfJJym5A6xtL6nMpOlJYS9Tt
Z08z2sp3eOIOi2jeTqJroI6v1HVuDFdB6elfa+psg2JZ8NFkogVl3KPx15y1Vmjl
uKALByL34oGT3edr2lPaLTEGTVxfkFb2sStFPxIiwUv+f6y1Ek7uO10Zn+/2QqZm
BvipGkXmwAWEiXkjvG7VN2dqBvDK67TcTQqAbDlW5XqLN0dSjTfGsR++ZAPZwAiE
NYYsVqDaSMOzDN0qtq03CqCUfDZd/xRskxzl50loMJJT+Ex/Z9ARnIL3wxWZR6MA
eR1dKm+iL8SuGQB7cPP9n5pn5MJ50mn0GxQPGgT6jBO9qH5iZbOie8uIIJjaWzlq
uhmDhAbH396emjKx3i06CeeUCEIE2uWO6Y4Y3qGGsJcvVC5Na2xaWz+L2758l9Kx
VocfOC5YKRon62i9HKEzMkOWrB9JuyOcgS21R8roStJPXOtqWRZRajttNmyZIKsa
RSBO7fUFIzI22VBmvlgQ6wLavKNEy5w5AMx0C1WJ2P1aB1H72v2qtzU5Fb3HbrIG
NUmhEkr18pt1McpdH/aTraK0dmZRhffLTKOzdv+V4J2m57BLt9VBeHxLiAtKCuUH
kGUTf1Ok8LkV7DK08BgDZw0f02ZkvRphkit99VPb7PKksrgD4S/e2LTbA6PRXaJG
GBAiIIaQiftQfDoTsUqdAQ8v2A0GBlPs1RbT1YkAPcvbc5gd3UJnWeKm6jMlUTUS
8IBUbc1/bGRMe1YiiZ8JckmOnVPy5lSW8djdni0+UN+VjVukZHZTNJSYUTgjLqEF
ZaCscAMEua8CbdFp9keGWIR7pBHQRg3Dwb2jEl99d2gou4Kv8Nuq/xkw1/PgLQ2t
zTkeYuPQEe0ixvQ/TOj0RSXIedHF7Z8LsY7rshaY10oat9TogMWy80GvEwZpS5iG
2ah2bfoFFEy/bYJz5fwH9SF/iCNt5D6yEjPilzcowkegpJLWI5GoyTIwbYVdUZSY
+J+v607wx8towMEFmqCUPxqAFW30IDxORK/6GEHFv/BEvCwb16wdcV1wynir23uc
xbrkKaAhbx8zGcfcaKvB+0H/ck5Vhq6Ek9I4Bx99vn5L/1BgvpDZaSGBDdwTtRnO
k+friH4sfv/NN26m38gwj8XD+Lpf7jDhXxe6va5T0tOg/bKWp8QQRC7SurdGYSXQ
Kj6eeUCwZp3SHqtdljZ87bisy4dZ0uCBoImJQ1V3v3d2J34dkR1kH1aCWsTFiIHf
5n5KYkT9ai4DFRtapT9typcss6i+l9WgPYoPJIzQOjb/uA8uY4A7cIrpro7RAUWP
45/boJqOX8SzWW+oZ+W54TeWyx19GB7iWG1Z3lQYN/kTR0YuDt+HecWa0urJvWIb
vzHMmUeVAxZ4h44TOscHPIj9Sxg96A4tZC3jc9lD5+rYqH+CxSn+XB3pYa8PJaqj
i/bwCcZtFEtPeozISDme1ciq7xAqvxhbVrITvKMrhwJuW5hkNfWexfbsUrtNMqzK
4UGqoDHtzWJK0WsVuOju301KE+JldHYwoSHzaY+bYzJpt8NLD5lQ8aaDcvpRtDps
LRgVjRQc3FSKzW/nQmvlokjecI0AWMGe7LQdocDGuR8sS9A/mh2gZtamUcK/Tgwo
zfxY2VnVh57VrdU3sIKiGbcIbgPz3on3O3NUfufat5g6rWn6fj1ic0aszEZoP4nK
qRjFCIbbT8TnF0yG7aEIq+EwPIAFp/h5nIGyycDgNeCIU5JLrMqGbSRdy5Sj3fQS
h45CrCzHefHr8qmNuTk07PKHb3hpjSTRjyxE9dlh4RHg2NoxBGSXHZ4o/aunV68Z
KwIsVJZUtnv2Qgxo/xVFsnQCvUmzq2FyLCEXVeyTodrkmK/BPVAI3vg8LZ8YiP+G
NY+VwyGCOTCutfYek5Sig0W0ZF1VbF1leNF8uckisg7kFoX9dGhUrF+oID1KYJPU
lhInaZiSlJoy5NKWHhvsCE+AKA4Ezyu6y3jSXaI88FwCIFBDSrSbLLbLSj6ynDoG
bnoyDN5J+BnLeSKJ4S5bmg/dwcM7rwSxWzzIYxNP8dDEz6ouG3mI2yqL/wuGAKi3
Pmw1Q/CD9+kKUObeNxSAj9Mb2e9SS+Z2HqESAS8WOUNf/vwFyQkk58QR6w7kgUcj
eh2onUmXBKx6rNE+zXW/jsmM0edDnTvtizW8MZvYqwR6sko1un2yojZEo+CHeRo1
mFd/3Bx+RrdvIKCXSYpWTGI5AgIRVeK0FXpGvLquyWK3UZhHFZtP/vG+29Jonguy
HmJM9vvg9LKGlvrrfByv9lC3sP4n1nJ4XizFJ+nIaMQgsdtijdahOZf20NpmEjmA
CtjrmRk13V4dzgqQakzNWpVZ6Es8dG/5WKMyP58Bi8tD0X0VIdhZ5huG3aJkMC1u
WEr50ov86OpSUT8ZMed7pgExLyPt20QHtVMrh/95mNd3Ri8lCO8vrCNCq7gAAia9
/NBxGAFrbw2CRUWbNb+dOsblUDx4sOFrqx0d4f5VuF6Yq3mBX4aaftvO0wj5AUaw
zhPgpaYhfQxRDydTY1dx0fxSlI6n9dZOEEM+sINotihCPHjVIWHBTXAPCzATVDPy
h6fNSXIN6SkDFjUwhvoIUgUqNcWwKcMCWfWesRBDaR6vso/KIdlA19S7gngmWXMD
osahfFm8qJyAPNReoF3/ACV+sLMVNMAmn9HgzUfa111vqefzhEGyx1YWhznjPGle
X+ja+ncYLsfpDsWyCVbw1hgEaxVihIEdAyIf1nc6TgJ18VGO2lWbSp7w+L2UiqQi
wof2T952mAiALtJyKroLIze4h5wP0pAzSa6kyM7esM9hZeoqWfWmik8zD0giz6wD
f8OlHMwwXp5aVvOAdM1yGDmuNZ6bnzp6Y7zt5qJU/rFEOemGzYR/2+szG52J0lGl
3g/mxxatobD7Lbl2nv0ha/4HpGMGodbjwUPpxTHWmcAIuN2Mah58kTOGa/CoU0ok
rbLqasSpncQLCPaE/TlxFC0aZDeEmXQ+n+IbUKqTcn25xxj7XuTK97ChgXxiHASM
h/mdNT00peH/sY958/ymlDs6w6Cj86CksVCZDZUVsgZQv/Wsi8Xd/bnzDcUWN8Pc
Zn7f16/TL5JJpSArXT4o9jevyoVRpcxXsMMzTiJwC6k2tlS7xTFu3QCTDWzegyt2
MFef/8/SU2GMuP3pLZW4nDZ3K4tHzeZf/IcFamHAnr2vvWPgzG0zjr2TW5sKc10c
XSiOI3cV6MZzo4bi9lfRTgaRxbMM6/cW/LlCPKNvwIc7VLhUYqkf9bP4hcTEiG7t
4wf2WUG6jmH1GanLg9UllhFRGyDYb4tEkPRc69IjKurpRx4m5eaeC+vUsHm1ueRh
JGhs27VYIv5CDDfjsOc50qIdjeVUeDsodZywP1jVWe1iIlXe238J+AXxeEy6EuUF
mZUzSZmMMXWwZJJoXORJkE22vR5yibARwDOZK1dLfOP0TqYpvP58NWk0s4K549od
FnnKPvbA7YV2azmmNsQVLrxLIRwtRq21iY8pHhgExEvCxdpETfXsLvKICbmqhEYK
pxes8qo7lZfCLoqC38XYuRqoYLtUTQP4bGNHV7z+KV33QevwWkz8jfSuYLXFt7kA
LOutX2MR5mj2mFv2vHs9FBM5CxvUUwsAMV+xIAkHvhC/qhWS1LEKW3lZq2On+c4S
K9EXgResDXqN1rIv3LWHdrHya4CHo0fAEov1yIK8/ebX4WculsyIjFImNKynCCqb
sZxYR1rTaEPAXmiKFtH3LC2mgeQiJV0ZX4n9xlx4oxZ0azoDUCRZ8VtEVNswJP8M
schvbWkH8CQopTSQhpUd3DcW7ERAVtpQV/WmW0CtWetCu3c7XglL+V+P8whdF1Z4
lFVm7NCaWAzCSFsBazBHNWy4ggOrcQAklzTEF6ypJlpbpoJd1AwwUygDdIyXHm8V
/mqT3K/uw/FI+Ax08jCD31+aOmmKoTHyQlK7jZKRY3b9OraqELpymsW7fKToZuVv
Exk1vkYnBEWSuU0lXYxwTKr1QWiAsCusQlSlGX31g7ikQesWyN2irExlg3z5X7X8
/Sl3cg2zVHwfazIfffzNfSiBQjIF8JCVcewEfReU9rssnyfWzO1QTAhH3bTudM5d
b4kQGrRPU5GWs+YE8lyyZJaN+CxDCq46/fWX2oG3YTWad6ge+9Ugj/R204NlJZZ4
Gt5OV+VF18i9voNr5L8ovNBOz3jXg/7al5gnoZbM8Uo+wk3KUDN85KvyKS7X8XUn
buYPyo+IqLbeoOp9n3wIDfasXIyFMmxw8D1CL5mdr5rymIxaTz5i75SarQY6s2xD
/lYmoLkzmQFrzVVVAItQ7+bu5g062tj2DrEC40jHcjz+lIYMOTx5YAQr/kG20lHK
4dazAT4b3tMXhQ6ZvNT4l78dqy3PL/odDdsdQN6p2cG5k6/GwHLdKSJrv+C33Zp4
uYQfkq7SvT7SV4tj4O8Ybe/EffZJYoNb24tONt6FEgis7ofetlUDyIXkfAIhbm7g
oivwjwsT+NUmYiRKcurtjUvy7WCycshnQj48W0ramBaxXkjsp7ye/mfxORffTV7Q
JcecQzRNZtxhzYxR+OKwndZP4nchHbZbXSblqGetWywa0ynnWkFlaZ0yAmWBOYz3
g2RHjE1Ka+2Kr6lFKwS0KnhDgNaojm/zz7C4oRPnFv1MeJDVfdTKthoYGiHwH5bL
ZcCfGcLk3RiiGNCLusCegX8U2xcHlB3CIUyCKLfSfXwUnbiKpeL3Ww2OtSp/XJBs
dCaHDOgZbCR3pmsIIKptzGTs3NRJr0fm7KiWNr3MKb3CygrxEYfUmJHLqiO/Pyp+
Lc3eEouA0n8G8WNzAS1HGLAWAdiWNItvxHjSSqDqmb6b/yeYYedn9TcX71fO0Mb7
P5C5T8gnTd7mt4nsuDQAzUgoNlIpukeCyWMnEvLDCCsCIP54VlT3UP9o0KrhLOc9
oeSyGy9iqvs76B804OETKasErNbzH2vmZz0QLymWJ+sRwG49Wf6kSynTJBmcM8X+
ZzyzeYBSwWUhaNGrqvJq0QruO5G4IQnrgL2IaeFEVfRBdMd1MY8kXhTN8nkFKgeM
CNN0qMWoIjCXJkmmO3rQ4k/iLBXcFGvfhJfCaLiOCDGDB+Wa0JujKEZXhoCAelUl
/wMhfdp9bVqRp5tgHXImP8rrVFuVHvhBzRpT28pTSnzoZaWPafDu7Yp0RGgIWRLF
2iHXEBHJb5o3DbtBTjk1fo0//5uF979T2uzQwU6CJKkEat2YHFPWoJJpJCwXkKlr
TcOGifCHKSwh1s1/l+I6JC7C9QT8tBnLa0f9aHELPNxfETC+fDDR1FKC3svWkysP
O12tfMGKgdpmo/bsyqVMino2uJZPe5oYFfOnufQLJtAJrkWdl7m0flR5b4e64Mt0
PRa2Kh8Kzm7rgc50WfVnWRmKNI/gdWGNpuD5/ClDEmqvrO5rhu0o92sj0T23QHRP
/US9JRdc5QKxY0E5oCdmhMyD+M3unZZuiEJk6BZpdQvaYx439frQQlF7PjQkNZ8F
Z2rXbP7QNvSlQiWgf9svnKt4j6sPJ1it1nPhpiUkJvUwTSlZTEKHw6gIFR+uF/jJ
gVTJ55A0V8TikPjBcAuAYo0ltdWQiXsME+439PBJx2aPRpYoYtBr6r86tqYBthZF
AKw+6Je1lSiArX9yLac3EhSX1C6aMDNjxu9jCztevVkVcnhxMuPTVCcFpRKh/7/y
wbV6YAW9Bm8X8cSyViJz/XXepSUMGfKMI/YnH8MsBzqiYP9fbNzaqjMJmbt08keI
hsh+2a+AaFa5PXcItz6FISi5jUaEP8gzqWQKK9zEFDUQCV/0q3bWHnKBCirF2+Ok
Ef4WyTAkQtAQCwjP1S/DCQoAH9jM2oWyIDmD8KcJl7WEPYYweLQdI7lbO8Qayvgu
tzk/7BybWc7Qiz0Fo4ZuOFGZkqQzSJaM2XNumLUVa5fjMbrotEhFR17RInBypnnL
BNnnL1TKTGd5h+M1+EVrMMYpRgA/PvAef38yOV9L8VfbrmWrNXArovAjYYRY4il0
pS2dLNENBdTTG23y6OwKB5PcrGPsJO8ppYNqME5aV6FFhtG33rdx/t0iF7HjqrDF
UC1oPLCWJYZ2ThEa7X0ecLv2E72FdAmqtIvwoVkchZnnWYLL14I1Woom8eWg+B4M
61nnT28ZHYFdxLW4EHHwep93eu8VLjL76DN3hIuEUC872I9P9XKwXbd4soC9Pgpo
vADgy6SuoC2sSVkdm14WR079KZ6MDOksVtwRLjpNyYBwW58l8ejmE865thWU6cmZ
Sz1IHcpEKH8Bg9rwZijx/MtTJ2Xzz7FDmV7fc6BJ2hiizPipAjmUtLdtEoMNMvgs
QSKeUzY3EfXhqyxVf1wu82wuw6OVr8DjcjUKOPPlaDsffkCp5dytN4yN3a9I9l2I
nfwZlXYtX6fL9mEXfcTxqFd3PxfCDYYifq9V085aOVddY2WgJoxMPTt+G5MBjRyr
doTWbBUJtH+MhHoU9opK2MyK9bYSDSJ9EqRbnumMDXLKpNoMX4q1ylsI4Fr4JP4l
QJYWkAGXBz0pdj4O4TC9KrzjdOy/dLwQ2pIszcSTXW9hTL37E3ZLlO8Xtso0eEXJ
pTHEgVQ4Rby86DYjQ09VLzEU8WhUBtSmjGx87B+lZBlknRX3R7XkPRS0sXgxpWqR
xzzGdnPZx3vJzHPWS2nmeKbCAwlJFwwOLWIpOU25GgTlf0JRM5gGMXhzK5Cam60E
/NEx1/GKZUg6Hp4lbeInHuTrz/QHESUmhSyR/S97DEEVZYrZ9Xmd2s93OCqaer15
Wmu/VGpIiFm4VK1glC5E8BBVjdNfgJ2oGc5aAquyTkb/3wQUpu9Ek9RoJ6MKWsY2
A41mZLcDVGUNAyeKSchB6iLTn/hOE09gl+2CUEE8iWAPQfClHVGzqljkH/l8bgUD
iJi0cv1MPWJ1POLJvrn3Q1LP1fdLUfpvcrNzwUPKXALZRSEyzgHGklZFj+GXYODR
ztXMIM8h2eLZ9tOhThoRpoej+bnUGpBApWSFj7xeUxMUw0tcxNOlNBHYJlqCh2Rd
Bn45nalRv1Zkd9+F5O7HPKbUtQeHXtEGmFUDF+MBTHsLNgJGW7exl4ABiI9ozhtf
P1DwXuuzOmBw7684bTvdT578ZqypAxFxUEYY4v/Mbx22M3E5gIyKMgMTNec0wa7r
81NRK3x7UEqSMWisZ3yklD7FpK1RVPw3JeiugRpdOyh9dgg2SdDdveNo4/L1vCBQ
sF1sDiZJSKgrrVf0yrKQ26jEoJL5otbsG5BajqfUrrmFjAiAClng+SN878iGaLEF
nbS36bjM7Zmhh2rVWvxbg+LBz/esEH+WSafwXDSI0c4Fwat+LbR3D0zV9u1KKFPv
2fNa5IdxC/xBiZlaSjYn7+qHTq207vGYN86mYCyhMOH/XE4+ocC/RE52PvL22Mec
uxsdngoKnMbnTQZR/1hcbqirbafyC4H5YDJILgyEu3hCT3CBt5h/ZpCEMfMb9sTS
qqyD/WF1P3z1xLV+xFB3lnkww8k9zAhDM5KG053UjblID2L2HaHXWNY7m/yugF3X
3qIrjSOIkFllJX8VxIWItUajOavAbPOHPV+d5cdzOAxR6g+y5krrPY5GnIgeSbqs
W8zEUdH77yJX2LYzMXooAFJKNE2+eMOU65HKcwvcooQ211XsY8f5L4cKuC8mixpD
1VOb0Cl/xg/LlNuChL2cBKxHSwnH7p60yXOShwDsbrBe+budqiZZzppprnn8OQBS
lZmQXagiyjJ+O5AdV8lFFKlWrEYjBVTbvClcpHUjgEE3Eq+fYkEeOOdRWFRxe2s1
aqHdYzjvqXXs1J62zbcDTqxD811PjW9w8H7YW02B9ywsDQCDFhXRRRrZCjgjrgc+
F5kOlUI1w/wg3ZBGft8tGI6TTZDGef6Y3vNOLJzmagOh38bSS2Upb/YI/URGS5IE
XR8v/3FCEckdzgdRYl27dD0aqTAgW/Fx1dnZbv3zu6OLI10v5c70+sbZ7W4nj+8k
q25vvuCc7EblVffHx2O5aaYDtK5txPUWKXZHqFdFxlDq6gep8zbHF8+IFG2W1IYk
63toISThhWivoSKSwFhSbLPeqxs5Tig6JhdqZ4hbSq/TUeA01xJQDT3lqQJDdect
M/eaxSDgvJuq4q8ZBu5IVyGQul1lbS1JxPagVkryvGj+mZqV0SKEynssdE5A1EW9
DWQLjOu2qJlVm64SKxnPpTpDRx9Do9lTGs7C0If5RYc40o1PJa/1LrqPygduaDWC
Zxz7Vfw8tqgYDcBuTA2wg5OFKiWhZ1olbX6BxHCHRTqzMyBP3J/eoknnKNzRs8k7
LJTPU3FvY4Vf8cYhHksBYBCIrxjngne4CvE0/druDrvbRgqgJTVgBEY2HVFvvjE/
14bDFYeZSbUrkJYNgXT8gIQLrUR+daylrkr3DKEPEzCZ8ZqfeT4SXq2323byACV5
Usi6RAB6CgXawzcFJ81uQq03h+MnJ7snhs3kbKc2VRv+WEDnf3O/idcFPi83V/DI
02ZKYzVrw12AezqGjKOpGFqj+2Ib78NsSak4m6UFudIsv8xmydODCYzlsT5MYR8M
fSzSYJxa6go8yIPSFjHxMLDBL2O10jSWexCnYA5+OqYRLtvLCRi8bsL1hPka6Yui
Frrzcab2aQSZmkiZ3L7cLx0lccEo19V4O7k0oUH3ZjFHznCycMHuFf2P9bLOI38d
IQKtvXV8pQiKIt4xavoQTR38NblKLCpRAig2lhPzxMNYufLkDwqMfEPimXxH6Eb+
4svPjCC5RgyTT7kVkJAzEorJO+Ohm/IB8eIPtbZ884S2xLhtw6XZFOHlagvvRt46
aAm6MV5UcMCbHJ2Mg7yNu4kL8N1v9wDdn6gJ26++PompMQqPYNm//x3JaTBmYW6i
5qO3g2/18/Sygg9uEZhkw8C6avLFVUlYp86Zh16mdgv3lJES8iFWyi74+FhmXTXq
dP95qH1J8Y8zdmJqrEyz7OTIQt/kl9RrPbstpXxH3gcJl5i9wkxbsaHZONbC99KQ
mHxbL53XE5pRPyBhYcBul9GQ3T7Z3UQtZckuEipeCgHuBk9fbwdKVnN1cngRY9Be
K1lj4TPzK7Z5kJ4gfeColaaEvB9jZItFXr3PV4OvEHnownpWnF4ZCIvSJD4PMnN3
H7LlyPK9szrNZI1Cq2QkcsRyDixe37jsJsTkjlizJzRIMr9rlhhHqMk/lVAP6G3D
RKohbBy9Y946TomQAnAV09coTaFhSfIQN8H5ccUjollztODAb+mQTdrHFs05t/6i
kki/SOe5CyJc1TRgx2BGjJL2DZ2sAx6NGicJz2g6xWkGBbEJvdTG52a70dTw3LbA
ZKZPdA8LE2iYXI/ucUWGzBfnCHbOzb6PeFnBV9UoqUTcdMx4TclfInm/xdZB5Nax
lVbR0p/PYIYiGmi2V/UrX/7FzGvR/fApKCQs+YZA87V5cFxOk61i1hVBMOpuqWWy
OwVYqO9NowXGZqEDMyIum+hHY4DinAn72MlpRNLWkRXlTyz+n+NJW90pEMpnleFn
69RAoiN2A7fVC7WlC8JyDPgoDhLNC0/pzjwTf8/u1B9dxlGWNra4lSmuHJPsBPSx
2ahRaf0HtVAk+DUt5cOas/EvAMQHlHZRaZAs5xcAvTFZFKqsLzW0srd06rD0g0HS
szRgbdirYIkbLa78lqQihcRpD9XSQjY2qeRNICEcGklTyy1g8/dyfJpqtoo6aRax
aYQOoYeOmDMC6YRpIa56IWV0cP2o9xFeVAoQKWgEF0EOsYFXDYZRAisPoTmbJ9Wc
hdX/gNpdF5ZNoI1ddUhR6CBPyU85uWgh3fK4rK4Y5brWX1U9s+4UcXdyHq8R+gz/
ZLzPTJHseEw2IiwPC1PSO49rC4srlIRynNpmPkTHdXuYrOV9341rcjCBmFNEZsIp
2qPvyz7/GGSteWpITBPnwYtkMxES+6TUNeElA4xUtndDFi4vf2n8VC7EQUZb54dT
hXPWr9rC/stQpmE2gxs6hqxG+6MNnzl4I43OnCJ40bnry6Yvcma1OP+gE2leELyb
SyQ0kPoLoOhMXs0ICcgRRe0YiA5q2v4FSBD2a+ArdkwOtxqB6q7SDGzLj0E80gR8
lU6NmBx3Ui9I250znwzHGJ4vyNTMhRI/9CHja3S3beWnTQJxzUUGtpBPp9KUzn+5
lEaMqOkXkUtYpoFFlbKB9N8CyyYrsH1ZQu1cfagSGU4DkaC1NohSSmVIybPDvB09
qZMo2Kb3gwLhvdsc1sq7Fst5Ivn2UyYCgQwzlSf4aIZlvFCgjEU2YiLWoghQ2E/n
4q0xgkNLPsJyqy48RbESOiJj8EiyrrraTjCgZn5qpeSRI2FaKb+YKiXMByK0um+r
KXWvmiu+WhnEscV1XpnFesDh1jnfV2WNajTUeocLifjYQBnp9MEyr3MwmWiTa/w4
BqA8LvFPjvWqdnQ/hYqpqN437tNNd5ecEu3cSQwO2KfIT2rIAWCK+J+cK4AuH/sC
+7azYDDA99LVbHsN/SQZv1PknJbYkQcEGUwcwGVvBLVuO6aRuIb96gTa5m2emgjq
c+HCpGVLVVKyxHVekv9KrhlKSd0EekaQfJlxGxmCqHChxe9aTXTrp0lh4innD6Jj
LfKq7pSShLq3GNCBpk4xv9Z8oCPRvq4PWTVg7omGL00ypHc7fXCgRx0pAbxGv5sD
nj2iDkZCW8/yBciJzleQ0ihRhI9l8DzsOmZmS0svH8xyTKV7ztLxAWtmA9p6aq6/
pQPFy+fs4iOBiouLr/dPGMpbrpHesgHZkXxLua4S2PFYXUgE/spxLMfqURVEu3Iy
HAukXkMEdUmgLtgb92oEiWrHWkUcjV55WwPCiPUnjCHEc5eTw/6wyjDg2pawNJ+4
obFkL1d3RcXroiTu52AR/9nGce7l63qCbZ5ZpeNq7OmgTxCjv6c7MDz/En/NUKM/
FfAvW4DopytNoIG1E/8Y1JppUe2g2Tp9+eAmCiDfFmOtBXj2MGf8YFyT/niF5PlH
Q7kevE1bhElvH4WswU2eGKTEdCDI61jBYKHftFyUL3YVIUYjsJaqqVg0eLr/qk9E
0n+opq/6SddaK8nloAOO0C+FpZprvXvLnd9XX3NA6+Oza8+MUs6s+nDvmdKfXFoJ
X1aOKN67v3DUkygbEIFU4mx/BntqlNhjStA/Ig1vx3hDZhmRKKcoFSwsfLdQis+4
kyifOS9rwDDlaDzaU+P4P4ke0YTjHp7o0rg42GjKPeLrU8I/MtlwrlDc7t6iOOkL
EKujlYARlHdqBvY02dqtpI7G7ZqTGdOxI51JR3WAS1HXGU3uh1EW69SIEmGpiMnV
nyH+EhiKVFL+RxV10Ju2gk3PbVllmYmjk1NTPu+QkVehO6EZiX3Bl7JLzr1AhLXW
RuphvuOx+dS/BQdVLfVgtIj/6BthSH/2Tk3V4/EymQuA3M/5lTcS5nhtXgMMOWAE
1tK8qbPZ3Q84fVfrapxhv0iRnrFIsgA4KqGxN4MXnSJgzjBMlQhYM0ST5CtTAGjI
zWOGo2K6LV8cLD5y9HXR2upE57kTHLP6ql0qEQUrh9UMQgy8zaR1bMe4YyiTODUH
daY0XkcE5wV1pA2uyBCD+FG6xQpJypM9jxE+YZaReTNSKXYF7XpkWV2Dj+WXLQVU
Xg2ZB9YfjTvi+OEKRlA9hxL3kqVg9FbFzj6YDE/CXDOgELVz1EJlQUc0jeq9Diqn
7ikPzTB80Jveh+DicX80m3E9VKZ8Td4ctJO3dBzZu66jg3ulIBZs/udWUl3d8Icm
1Mvs4DetqE1AT6PGUBVLZdGlGofcfhQH2gVtPN0QU3qcSiW/tH49KCA1jsqNwg+m
oX0Lc5W/yw9XI6XgLEK1i+WlKq4Xkqes6nKFbxQ3F8l+cWQ1agDJQQHQo/uDv5tR
jlx8vbGVNPDztiXCe1dwbBn7/vvethbhPho51aHVX/tI5YbIpaT3Kj70DxVq3UxZ
fjA5NomnrgVLp6Vj1ufr+Wf6KU2Mt8wnFEaLcsfiaGIsLfvqjZZ+FQpY9COS+8Vw
XYOv6Tki6CrwFzFNC/Ia9naFKj1yilk6JQn8jkLL8NHyaffyuyivmMKdkpwINQ0m
B0mxEh95gXviPSB3pRKl/FE36ARuXxOh8B51wPkoNA9TrDlPSmj6KQySoJEv3NE6
H6NfrvBwfWvAE8T9I+X1z781LnPkIWygIa+Oc4ih5tQ8RbTlNZ1xL0bDssOxpIfE
v3UtStzhnxqgHs3eg3YQljEzOEjI7C5iqs5oStRv0tSoV4TwUCpYQr8yntrNrXj7
Sj72VwqIHN3XdQF2oJq2Qr/nXTznRSjl1iJhM3bxJaQWJ1S38zXskAqN9D+bTRlf
mSgrgAnNSAFsDuw4H8U+C5Jsyo8hwCFs5hJKXVPuy267r4+fQ3OrJskVt+IIEwmV
mgONzsjrwDH+bXOI2QE2JGK7Ac+zVp2icO2Zqtk6IeR2MQNoP2HLVojxfcqrjRIf
UQPisPDC5yI4mEFaj+fg8tiFUN9L7ZM+nWn/pUoddJyQbjHZ9MKc8eVau4A1wFtB
aGIP5HMpWP4W7OPFJ9QBq9P0Ne64wyffo2/XKPANaqrzsuJOBdcbyYkNaguvuRvG
R93znHI/NNkKtgemBgmnz8XPAziVHQXTeOvWsw0bDkkRyoHxf8wFyqgJBWljOFIo
9WED1yXGp6XFkfZ03GOZyknVEruPaQsmuqA/uP58pT4WTWl6K7CRAWhalz8RZkYm
tQIS/1QSTM/XELV4Qajl5QkBUHrZY4EMn9sttWgyVsxevxcmudg8Gs5oSJoAxL3B
XUqP2VCPyuXp3d8sFFvCd35ILRK0NVBXDD/1DTeDou60e1+goqe/wLNX+m2+SPyy
h4PhirlTqRRTiczLiRpAx96cJgwZwc6UeXtxT/jFjhLyxVpTWZ8jyDIosgnYOtSe
m6z1NtmLASxxNFyPf574rTMkyVJoNR4kIhd7+eCsQcfRYDtjxG4275i/hiO3mwvT
8OEitiT1tR6ZzwGdq7/wbGTHWhJ8wcJbpPJklYeBdzkm5KULpZP06xTb4F1p/cVS
t2wSsI+0pze64NnbtiPZnxPxYVVIUBaeY3qB+ewFqUiV4b/EswqATQX2DQ4BBdW4
2lV9qKTHStWIHb3ff6FxSWG11QF9NtOVUpIyz1r67HhfCS0+WzBGZe0jI4nQ17+P
Uph7QErVVT4GhE7CU0bk9omv1W0hRsSYFnY0XdLZ4ejefXv0s0F6JYL/QWxeVdq7
TkvB7FEMGs6v2JatdpdYATPIGqGCXOt77KQZekzOOuctjPA9A/2umI2jCfT+1YeE
WGd6S09lshs7jKWeMqF+zHobF8qCEgybSprqZ8xGfEObTt4EoLWuVKIVrotlbV26
CYx6fSDazBu5XbYQLSjPF9IAE628PrnUYvd9P9C4ApgWQNiQ20MUJxo9pkozKVeG
ca4mM4RXTfPkC1lXumZGESADmmwht45mEzUfxhW9eTZvffgSKLymGUc4D0M68+t3
Ab4LJeJ6Z9Zv7Ye8SyPkWxUSNjNu0BbVybsHTOHtP6pDmlPeoheO+BVaqsdGFlPC
LmM93Hs1IThHs9pNnOQKOeCLcNvJAMEwdiUJl631VODwj2bDvv8P54EpRGA8d2Xr
pQvT7dCPjYiqaQcMhrI7tn6htqz14JpwXz6axaZJqxZlAp5m9vqHFT1YhK04GXs4
3XhmpbUek6eM4lQl/bPDptT9xRLF01ojE9ciGrqSii3Ki5RlkK4IMaa1mgC8gzTY
ULSgfEpk/rgaQP8FhrnQ/+XgkoRPhnKcSUonZ3uHfFS0lQ5U46Ktl/LHVs3kogvK
GU1WRpv1nhA+V9VnbXRIAIDrlol4p5k9U7svsXTkYooeuedrXSHXn+f6Jx5eoJo3
SOcwuXrxfoRSdtOdpVP+mZLbkVIDAQLBnh//x+9xvXKVNhMEddeNt2+g8E3kyXL0
4lw3bcnIpJJn6mqeW078X1disMaJ2eU0J6CHK2KL++DtOk4lVhVdiYOzWjqqf1vp
LBaxVC8Utn0MNMjqTKIkuvdqLvuM0sObUbirDPrtsgVu0rQmQXxeoFutF71rdUqd
HRX0Lyom1sx25QlCnUfPTMH5mcoRV74sW5qZZH5JONifMu3tJDQHhF6DvH3rrRJF
bzTh3vBIW1pIWAyd7JIIMiQHI/WSmGdNH2fCchp0MBatZUrUeq6KTLbbAGCw9pGt
7NxAd9LvHdxzUdVhgugjyQQd/TqUd0JpAd30Ny602J6arccF2zSaMmTcgJ0nha9w
DnydhyGq7KOJW+dOsoZCL1PZdAOHZklGk6+snLAiZz1sfKD7xAcqn+hWMRlhJb2l
x8vItAknuxpQgms8yurCvlrpyZflQ/nXGidka5/WBJzC9NfGuzB6C2tqDhNyv8ho
MgPM2d7gPIoatW2P+/5UwPTzQmLCl8Vr8SKRbN3bfoaWpEprcsHiUf5Usd8bvLvl
OTBbAqJQzgfje6LTCtxG/vd55S7BtJxsqjcdY4EKSX1ugrvubv23gO9YkkltlscH
J31s5O8/izZM4QmGtxuR2EUn4KT3irwHJQ4uRIHlSm3vpuB79aGPwX4Uph4s7VYr
Pqj26SFpaVyVVOY0Fnm0wYrdiFuvAQFtOtHzkcfUzS6wMNwYb9Q89Wa5eduJvyMc
XWFU6FERiTjXN0QR7llPsAjyGV+IIi28fGsjijev8hFFte00kuvQ0WOupc4LPzwg
5M7AC5R3StPimAlTZWRNfITvyCN58B1xju8IQldiw4t/lPNNNJ8c/N3oj/JbpE3u
0eJ5GU2VnmlpUdxmSxfvcgzWL8wqoZQQCeHB6nlgeaawnBlFlzRwGzG8bETtE1SG
+eFY8YLwpKjDgrj3KJvcpClirfehNFXD9GnYrY0odwkcZQouyRoWPZHV2B/LTQSF
o/H7vLahySCILX8BSEp0fPlegiWzk9sfRjDtZ8g92ya78Xt3t4w3gKRwlkvxNzuN
UgCzlI2Zu1QbZGmHp53cUmTL80D7GzL077nd0VaApRtzJfLoQkdu3SJpu/YNiWtQ
gPX2MV16iUP2lekzedp7njDA0QaP8j00SIxYXCDSvgRJIDl0mkwc3Mvr4GB3fsE2
N1wS9fpHhIBccwSk/f23fZx4brw8AMfGZzaoOdzHqcokLB9Nq/WdoE97B1tJAfHF
pT3rHklmBBPcRj0MHxg4Xj//tSniqQJYr4xw3aUrKd8mqmnxLvFJES18h2uBDDR/
qAKUQOzQKbPDevvViLfiDHZpC73G61dYLCkjFC3rlGeQg0IIlFh82TYYlHo2Tfbi
Tf//VXpgTmGoe6pWai+4raXny7JYv65X2jGrZGlia1CHEsx1E39Zu2jsKaWNXMCp
EvhcTjFs3O65lHHlfPSE3MMWUIq8hlOXJZlC3wvmSfSR3Zk1TztGuiiPDvpTMIKA
Cv+hikS71rRhWXZO9wgW+Oc7i8IVgmFTLreuHEaMsBG/giz3ULlqLbfbwYLoUQ61
uypd4faKwjqYTtcXeFO+xohdVSbjzV+O8hByexE9BMmsJnXsTRENUE84Ex73imgK
hvft0C6Jj2ZLlwZ7fuuZOWLyOPbOZEwNV6YzxP4Q8e/aZ3QcGx/qWunypcAdnLmR
M5m79PinvjCvGOOe9A+aSNH5xpxP/kIwSkZ+f2h1EoYOQzl2fzLkjTS2C1CBMYsD
InxABc59BJ42qu7Pbe9WdjF9OoE3bqru7gbOfNMBJr+maxOzYjAKm+wPEIJ+FRwj
CTq+srS+uN75IGX/yLhfalq9pK/AfH0TY/QDlEQJHVIqJxtrH4+m7SkZH7oCzNKU
pkUgy59L1eAr/b+w9iaHCciRh0f08/Wz26Hu4+KQ+n1xmr6L0yvdUE33QSh1dRCV
5JF48PYkBWleJd7nK5CT4e6q3BUFed9AAAxXoKBs452MdWUC0lecpn/1ZDv0wSFu
78Z800hV/pc6xq00886Zh/041hdWIC+kYsyzpBly572KzkShqESQY1yFtM7n1o/p
4L+ZBDyBsHOL2TjjdJFUbgT4J5G6pB2BaAEIca4K3rmmja/4LwG2r3N9paaXEh5a
qDN7hxmS6qp5MkVecu4/9sOb7PYIp81QgfySlAV2NeWPOjw+32+fUTFvr5DqBjsi
4924gL/15DDeEFV4y+UGf2+Mqory+EiSdRbW1K698aL0sUtM0zI6RmW7ABx6Hfpf
HmLKOnqAa4tp23j4n+L6BxUTGKMDXHlMZ6S/QXQNSZIQvJBdrVu0wz04oaaS58OY
YOn/Tqlyyv80Nwp5TCAVWop0i5VbnZKwNu+YUk/P4TdSSyf+kBmgPsSQ5+yps2fO
uH0H1dVezuiHkpdw/rW1edQKWGpUhZwW4GrRmAB/mCdUwkOhKBMkM0zSvzQ1d+Ep
eaJGvT7ICU57PH115VRaqfmqmWoHl+WXonIZRTK91xncQ9IBfzJtNh4g8KYNUt8i
Q4tHwj7cVibO5AEVIlE+ikrOwS8/gbEXhGKQLkmA+/FwXN1zQow3NpxeMJEGLjDZ
/ZJyuHAUbl7ZykJb5ZNyyQKALVQx59JiOqutdoxhC7fXRtLWIxC7mhs0n6i7YrSW
bvUQLZdjfMdF2Lyt8JdBkFmmCB43rHdMg4xReO6q+lAWK6GsyR192NTuyE9SZnln
upu9OF7IM92SEfCznPrjStI4Vn+WnD4KbbN4JvsY+xMNn4ZDUazDu50XTZHMM71w
Myp/7FD3qirp3kkAhSHR2/Woumqc8Mxemrc6AxcWbxDIcSmNCkS+K4bV3U+DE9Ah
U/l+JpIm0AHAQgIYzuvYdaT6nq3to9eu0NLaiuHw3rbR5Mf5EeteNhMsfX8wkn/7
30RHeZMXox+Ht2aMcd+rH9A2hMZ3Qmv2Gz2IdzM75/x9EAI+Kf3N/vFSD0u/5vHo
YkDbATJ6zEIzl515ci7Jl3BDKUk4LdoiWkbJXRV9FmDOD58SiV7YxaGCkxLcTGQB
xDeZHTIwDFZmWSpwSGJBe4CXJ5jTEOvFV7C4UZbbwXoH8KUah1U9x5dSddSjkAUt
fwiKWlKhG2BIwDoNQA2SdGSvF/O3dboThxlGec4gKnU/lIfXf93BljG3f8xM4Ng1
zaCuFNWMZNlFjxmewbCDF+ZBYfqa0ZHw3lR1EnTCabF41/vsnZpBJtbf7aSntuRb
hflC5gsiAQ05RejORXf8AFqMZoRtCaWfvrpheefzDDyaadA91JNHMOAL2le82rRr
LkxzlPXH4AdH2uMKLiofQgPQtjHS7zxCnLybYDYFzc9sbWQrSaKpHY4HLGjvtQuI
PsXFxiDGjQWnJDpbym2HOvTHazQ+yqOdZ8HPOTAo1ANzOANOgm+N2Jj5KvK8wd3k
aNzk/YQv9hVrlZh4C471cNfL3brUzJfj2lNgTOTG95N5YpLwY540TCNHU/2lXz6d
p9bAyjfuyzgCbIj2OME2odyJWqW+yJPjjrVYgxZRuQ3W/6TlOfQQRf+jwYI93reK
64djW3eykSiu5uh+7N1+p5xx+1quYIsdIr93AS3TKsacPHAoybTPQDCiDgOi4sRQ
Na7TU2O3T2LRh+piFzBctwyFqaZF/+pE1Q+Q5j5hRLSSwIaeiJAaqsTS5yQRC9r/
NtJEpK1+u4Up4OQuqK01CTACuTKpvYb7RodBZLnYV0L4nTJp10KvkPQlTosj2xca
LI8o9vNzkPp0DA2hUzDTIo4kkFPe9gPNFN86MYNg/q/a5XQ9H4TnfxkqVvTDAQiM
ZxxHPrJS/o/fJAlwtu2Dt1G2UxgzixJRdbS7cSqBs5Piw70ShT+H4654KYk4BbFt
Lb2XzAoHe0EdLsTW4Yz+0FD/D82h/l2Zwc+uGRaRSzlV2cHDmJFeMZosx3TRau01
adBeiMnEQGi9lNrGqBoIb96yglnRPTli3W2oC679oKivrVX2AM3TXA5ncyWrHup7
KGt+ICmBzNoxnvabgY7PlSevxcD5Z7JMS7YYoYIrymv7UKRTrxMoQINn+Wrc4N5R
bG0/ucwRzDPD25InHb0uM/JlifpydaCg5mBnWTobLM9ywkn4tFvMIWa+xTnAfk9w
2p15nxXt4s8g3SSHPiktWhhvwymr+6isYcbPe6yu1mfzNbsw9i9/cQoi6xkPrRZE
s5tKOVfUQiyhoDoqwfP2w9Q7iYGTn3azb7FQsCYtNxcPBCJszL5hCq7yItEgkg4M
Ul1+I5cbJwsrWzke3DAKD7f5FWpJv2IXRxoGYC0pO7YHJo7H9RG5G6VOUsz0CbXo
E9lY+nO0hQLMPhxSUXcDKCybvnh3jR7x4psnxMlKRS2Z/L3X9gzryDwXhIsoJfHI
k5O1WLpIVMVZCTWlJJY7c8Z1k0qOW6EfgtPHlV8WmkKikC6742U+NaYk0mt65Qtq
ilhtmd2BhtF899b+/P93GJLuQEJ2E6RmDQAv7geNvnrhRcQpB1EUgIPGyMXDLRpn
hy7evlMZOmDUkamANk8dYapcN8viQzxy9NWISXdut+ZR/YoCLFpUjUI0CksY3O6p
l98RwXXKF2Ap9FRZMN5rDihJySY1STMiDtNMMg5VyewK/wGhaH2zlbTlp0oQ+eKx
/GiKqtpCkDPCp8NoXnJGpiY/jiG2ahx/H8ANHLgVw+uHDrD8Zl1aMB9Ns3V5hnTO
VfIOFoy0tud/zVsI+IwmhRwAQNzFFJ1zlhiKC6wEi+AGQHY5/qpCNh+h6RKNbCjX
T3vhsbc/9RL6bRsFaGeuxzbqy7+3618v9GNyMRTH/Ix1dFzB1v6xljEEP3BpAD0X
HCJf7OlZQziOoMKM3T775X0VWkIH46leGP9YkGnRM5CTmf8DAvdZm7RysSE4pyZS
QxEtXWD1GB1FbXCwXewUCt25Oe/RbYFe9Tu6425dk7awl2xFZO+4yxeefxfBMgIj
5XFdVp/x0dlh4ec/xuSJVkgi3/jUmQk7HXlhoAev8U8PtudsLBJm3+M4MH3PYWJC
8V0SDgRZXn49TX8enccFDKXj9Z5+Jif10rbcVgnkFlXX2tKF1qHcy0hlB38baBol
/p4OgKA/dysUC8p1QuSnDunNGe5AS+bzISrvIRrgzf4gqm8gQM90ZCMMUBuUW3LK
G1Wwt1U1y/DnKc3twq1RuumlV+D6S/7TjXtz7x/j4ppBehUvUjDU/YqxCtL9lnko
y1ogKVZrDBHAVJziR7Jj2shNQtUKW/dYUTQb40MrsEfGdVEp+uq0AsRaGSTc9aJR
Morm7sDjIZJWKWIiD29hGS1cbHBmtMCkUXEGGMaPk3XY3JY6rMh3y+ZmHo/jw4Z1
8+XoeXxUpj5PTNO3r8lQkvrAbGaMuNYZlJrnctlyow8uacebJVI5V4M/+niItcOy
KbmReOspMGHyEVcamDu/usOTWtQRvTQ6QVJBZHfkGmi1SUotEdWBjWTMKQPxaFDd
7IYjOW10BdgcKlVTivGELjJwDgbK21idQDu93U+PctPM0PhVC32Ociy33p7x2arc
vB8LfifdXaVa/VU7c7n6BYt9FcIOHWHbT+eNfYbikDyh7RTY9Vm7wL1LQa1fB8ru
1d7a6WEabsYwMT3sXekW0wHx2Cgx04ICok8l/u7dbC/fwXHMUidsw2iIy3xZW29k
T4CeKUvOy4XcBG2GLnBn6HbHcNNuvJuv60DnywAHWCcFUDqptVW+DmY9KyebDq4E
08DECvDWcrtX7ixtxRG4Cy6pL4o461DKWGTMO4qYU+r4nNXBZilVukmceRakwsSr
YdLBEGcQHbcy7sf2xGohZwdlUGF94NDzycrtQ7yp7HtuVNulpZWlVGZlRbtQYi+5
OnbpgBz0EDAp0Hl84nYw3QgoaYdDfQFDzac/Vt1EFoZRi6oAVZw92BnBUDoS0lUF
feAEjakj/SY06onq9tDnXRSLXLLks1Kbbm9RuJ4MiVWVTMIEQcd5OleJ8wbDXDWD
BvgyFvwOYEJ7Ak30v90hTgQYxnc9ee5YMFO6aC71/qEgv38YortEWmGsSupik3mH
Cdh9RtiXXkofhoQUyHwzEahwImGa7KKKMDdaubCbvAASuO1D4FXJsZE1OMrgdsZm
aLoB5ZDxAOSlYkf+qjDtUIGhKg6AnIXa0iSbw6OkZSjbKglj7IiXBaGT7JAZKrBA
c2sctLOvH6Z9h8Km+LIHbvV2fR3jAveDoghEv+Yzn/3aDQoSgm7NT3CXoUQ+uwEm
4JZA+jvkUjbvaW0+vCSBOzK2eqmgqNDNc1DF35lXeZsTYg+y9nLj209MVY//y3BO
Zu5BeUW1l+ikFF8HPAB+Bo8CLKsdjJGCTusJAyt4Z9o1QbHDFPT6FeZhndskpw9a
HMRgjgu2gRhHU9yM3z31gqhxr3y/+syqMWijW/Z1VwcM8N6RMmLZ/uuuX9v4Sgpu
YRLTK3SIxEUY8Q9d1YO/EUn8LM+jmBkaB2w59LakPB4HyNurhQot9ljIPEXYjDT3
34MLVc1Q/Vl19RBkcGhdx1UUuyX4hZXdWh1WGmAHRxY4Dz+sukvgSOTctkEfDqCd
HaOiKqO/IfG3d9FNTE/8auAbZ6vGoo9V8IAvWIbISrELxFW6El458VFzWKP6+tst
jJ7pCSLYmPnS39VDPpsGQADmM8hm2BuV/Pck+JR0v4fxNslmXbHKaAwfBS6fjkHE
8Blb2gu6LfYNMVA5fv/0wBprwTV2c6PEmpAxwQCsjnAp2FBzEJk3NllThtd1Mcae
P/KZREtNXlF7ZxOXXO+dvbOK1yQwhuo3d1rPpRivOzno8hNgu5YElVWs8eUHPWCk
H7Via9jpOVbGTcOgM5njFQn3jYfzQ4wTazrb+SZH8xU8VauuOW6kITczPQBzfPFe
Faq8lbXRwzVJ5zHqWa8rrCIvDXQgLalf/csIMrVj3Gi3FYsiS4rxD3DB84JlMW/6
eNBaIZbpnk9Vfk6Ob++aHM5gO6xxu9qc9qp7Vw4mF8tV/LHzg66Tu/m8O6n7Jdm/
oWb/F91FV/9UVkMbnXhpbs34u5MQ2wgTNox9U8n6WJgEUl8j3ewsUHU0VkypYn4D
xjLEbBdtEABr4tj8RDy35Bvi3LK6/Jhr2nN5787tVyN5SICRdHCOW+3BwKeS+2vz
D9DAaInRahrVje8JptzUFsnCPiyCr72FX1K0muGz1wcKc6padzKftPcqdC7cUJri
oSTnkFAV2rwBUFRi03hrM0fxKFvab6quOtDyd+whOyOrLf/0stgVnMTM348jhngG
fLLBRstHrL1jjljquuvmJL+cWIabjWGUx0UUQ6+AyGR5501U3YseyTkZ711rWpbS
ucdh2LqmA6kZzG3s7vmlRMxmsI/9VkYRDJhK/3wZa2+ZErspiWfbUDPgLZoa0tnA
QfTn0nfcu+AcDmr/s89S8V8as4XyeqK302XObGjgasLNgJCSlUr++00JokzeJvJx
OCne1QIQ0tN2P9G2rzzh3sQ5NC6mGSxZOQVRibkrhJsAHPeQc0zO7DhSC0uzQNB9
Eci7rLxtGH3aKUoCyHLrDhDLivhUE6mHLHr3uuRpiVgOG9zH4RZkf6kLyAUGAYpm
z5TD68As2DdH+c6SYKBbNBN95OdkPcTcNvLJrIYxUiwnWbHXzX1G7cHB50SgmktU
OVywvkaWQZqO1gQbIoTpssD+m4kztUQbwLbV6Ybh5EUbpG+RJEQLse+RwUR+RNOg
X1rnhWmeIKDSZMq6xG7c9402y3wu3hkkRYWQwsMhDJFCNYYTCkYrHlO2qPySgq8k
8PDGS5yBMRNasUKdMxJzvk8OpapAE5+USJ+GAf0sXrLbXkSd/Y9nYGXJHrpdKrc1
h+Je7Wx6td+X6YJdaH98GB7exK5BsfzbDaRWZZ54Z91KJGEze9e9guwvqMG0x3MI
AgeL+mqX//Jm8O+Y3pEZb98sSQUsQ5B0KWVmEBajzbPnnj1ql4WASzQtvk913kNI
Rr14d8iz7PHq4GjiWNgskzTCsoaWBKprPX3SdCMVidM7dltZpmNeDNXXUK9HR/wU
VyKGLLDTuBw/0cO5AOSJA6cyS24v3ZBumgEyhJrSidwHsnAA2MKj3maYoDxvM2mZ
3ZjOr74UFkGtzfueDWc9QXE/KQAgJhT6csI4i3vKlfi2C509Jw8dgt/unuSG4CTp
QLXj8Yz9zCu8zzbQ6iIGwKQemqXQT+kA/sfzmHi5HJvGxxMDL8mg9vT+CqrTVyWO
a0nwRyRx1MbYDPhn94h9N44m8zujOoZpSTSaHDf7KtABXSttBuJA2UotBW81W81R
9EMH8r5ihXe9sRX25/1mKy73VGyvfDIFwHdL9jV+3pVfnyfH+LJPwCFyBRINqOyV
BR25e/QY1Sl8gGVoo4/lO/KgPzpkMJUgwhclUrpoD95bjCK+nTkkhaVrGV/8BtQf
GbCZ8W3cbXhesxkLSEsn7Jj8qr5p0NG1/Lut2k9EcL7L+DgxoyNSNrVoAFGUjrfK
FjghICmIA2BHfcWD4xAJt2nx/3NkLyoEiVgQMC+/R4BVlDd2Xauv1BIO7yA5TncT
PTVrU7K7UVftE++R98eEHx705/OQmdUsZGjWE1kR86GvDeErr82GayRgDfHVl/g0
8Zl0s83z+erNmERII+ZSWOfMFJ8nwXnCaXe3bC//4zCXwqexrgO/v07Ny+gZ6HFW
bBLKbCb9gG4zvNJn5vDPyHWc5T9VnisrAcp6+pdI8ZJUgNUhB70I+nhCIgU4+kj8
/Ha17Wmq0+pucYlUBKhNOlx/FVkbStIrE1YZMSpp2cXKRYDTLoAa6qdISWV62mog
HhlFszzDqPgJb6+mJ8ZAG7J09HNDkFBsMeOsf2hxKS87LshWDPFdevioEVIZkyw9
0Qsi3WHPChqFolW+l5WZs3/LVdqrgHbxgut46FetGqNueAX0RpxEoDvrY0ytWhGC
oqA8FwcfJ6egb+uOlEIBMVbT3im4/Q2Whc6WSOyrC8rOx2McPm7AYfs54FR7th1Z
xNAlRXtwTHRLEXxtcyMUtUxm9Ja1lhzBhfBJycjg6aOc+WmClLGDLMav4Ho8hViA
LlkjnQgP4VofS6kVTgqj+UHJQXejfquACuP8CCLZp/xxIPWo+mmDbe2m/UECL7jW
57IC8N/w+7aJK0IeZdBLhQoZEMsjmdxK9yGgEjwhpjwIScGbESUjWpDvcgmRG7KX
EQi+2hGliFRxnqPAgkSC1woyck6OKI7bx+SvNKOFGtBe/9zHksir0ihjzIFIEKm+
T1RHQEEmeLpoQnwDsJGvLUFa5uWPh/W0d2gyoscjLX0A5sZBd0gZyhCNezq9eHAN
B6sdVGCmMo9bFXNJO3vvOls62B7VDT/RsqAspzhUAreD0i7Ac1tskE6O6By54ZZ+
ESeU6xTujxJPoUGTKXFPPfiSdXps6nywQLWpsP8ENFuqOyReAuJOcggRBNrkBwF/
oBkr8Dt7D8DamWGnZpmHu/PtEVa0OfgPNZPgfmr9asMMvEC48rZ4Nx6gtaQ0QjH1
Bqs8fB6oduCVLUIN/tNX8H/IsTzMrc3oHjY6QASCpg+HKbXjCO1435I6XwmjWFBc
nx6AF/GkrviyO0QzAGwj9lRs0dyV9qLqc/jGUWrJoZTmzBX32xc0uoCuyFF4CSRC
Kf2sTQI2Gy/26xfBYLxKv6xlsOkxTIIm8ZIr61Gyu1ze8/vKh8txN6bJ15kS9lTh
OpV//Vh54DdSqWyWDYFeBmiH4ErwMhimcefwzZuG0fSqudkokM/ygVxopyQA5nri
zK7Brmtiw+N7kq/PPXY1lpwt0/fXgve59BMyoyUGyHQ8JVFVMecGn5mE2/3j+evG
gARM6vmEIVdUXj3382+pAx9TFayEvkcs8DpfUS6O8KDram0Ti5K/NYbcjReBiQLL
rvabc4oX0JmveP061fCai3mxXdkTlO//y3jEVdrCy4vUcO108Lp+eBLK6fSHxbx7
z22B5kZ07flUCxVvIk8I7VF6U1cldx01fMUgqKOzl/jSyajSUtVtOS6EyheovQf9
CTIaV1nrFRNMVGvW2eUzRtrpcJRbgFwb0TWoWpRCWbtDa++kbO7m4+a2ffhJQ/jX
2hMHERT6D0ubPJTLLejQnB7uM2mErT94x2NufvHnbBqViugwyEeeaQlToLjdzJJU
ECPmrWpUA0unMJsMgnZ+5bWFz9M3YCAPvtXtxQ2L3ro3oTiv2Ul11IqAm6kui7Zn
TL7zGYRgc6XJx+mQOt3d4sk7suGdyy44isvJd0N/FgNaB7K5A24VReNRQJSB6hh2
ivOasIZUqtmSZYpQIJ8vogjRUIaDM2zr9S832brIRyRztMIiVF+kJ/kaBCMoZrkU
CzUo0XVapJhWB54XMV6RpHOw/icPGmk29GcZK+XSPWTjsrLy9CG/gZlO0KDRAHpw
1C+G8Y29HrL9oMXanxbkRPl8MQhxYv/jqlO5E1w6D2oG3bYrb6r7p8v/hUlxpNDU
aJQx/jp8KG1DKc0+mXWwQdWJjgoKxcXw3uNHUTEA9vbOgphtGPPyFftAEnsebBVN
nxbVUivCdU99AUEZZ+aOKh3l3Xy/uLZl8BgyCdyWkd8xR5iAT/GfPnfa/n6uCAS8
VyoJ1FMY7DuL5Z5AssA/BCOAEoqhUf9C3id9x4wgnxWbM6mEsbDQUQHpZUVJykgg
7QmG5bQWm3Ry7omP4UZHSQbM/iB6jw9jr9iVw1sBFzSRl4hvY0y48sgE8ipS4fOQ
j2DWox5QIJt4c/LqKr/LFuTLhLO1X7kFXQNb7R/VCJ3t/PKQjTlMPMql1DkjMAxO
9eeQxyu9ZiQ5Y/x24w9ZkXgMUjFv7ccH2NTKo+0aoMToSxzsIJbzRDoKEkTsnCyV
yF4B+idyRwqP2EoC7Mf+RAepWau8WsMtSPnJosPfCwB1OnQEzuBPNTe+Exo9BZla
qIt/rfntU2OjgQl1rfjyNpUbVIj+Zh66i4NN5ClH0Lh4FopZedgxCuYP0DM4YSPG
j2OpV1Ch3AVgHkuCjMVCGcQ/jmg6Z8J+MqS1pS/Nlk5Vm7VKV3XQDBndWah0pHzV
cCq9gQsEoRkiFamjuQJzQhWeURu+o/QwDbUScwnXQ6vqr+PDZdXjFy9tya5KG/AC
0woN+CPcTOAFslE/Y9Pdq33mBWUiruXdsk0LWhvl4WIYREChAtv6FsEdugtke6Ps
ZQ0Om9kREAAoXFepJguV4+OnlykdQXwjfHZTQU5rtz6LuyZGmFuUpxImK7s9eylt
BumDrCmY+w7uKvC9Jde/4YNBwyWQkNoJqc9uxPdRq1DlFfJ//Uvi37vOUm1TAo95
Qq7cYtv7vQAy4k5xiRnwsa/nE3fz7QQNg26uzjY8xy/JHrpJ7bARFcOulEDuFvTJ
Z80vvTlQdrDx+dDilmzwwh+ovpke+KNRQaLE1y4s3QrWgAU0e/8FeY9zxDhfRLj1
lR4XRjG2GqgfPTeEoetPdXUEuNWUGQgHr/DiwSiOpFqoqGPLerEYLCvwZNw2KwEn
4pDvsP2U37t3V2nMPjbWseEq6MwKM2HdM59klULG5QV47kgDTePAscYW5w5al6t8
p31irx6R1vemgJuXLZgs8rAgOh7LU/1BKCp5CphUQvrqujLcy1WD1NchTJlBmyiZ
hmVR8cRxLISduZf5E9fEW/uLw9iEzOSMdzOH7krGUq3AI2YBXqPZMBSy4GBh4rj/
8TjF4Q371+h6qS3ZAA3YexPuVAtwU4llDMpL+D+SRupZBqJCRcAix6MMgJTmYEOe
ELmAS91WN1MwQLIJdAcvOnzxzBf5eZMT6Biin0F0ccqn9zlpm+g7nVN9p/pcqpDe
SSZZl4n2ccnXy3tRGMAgYPHYOMexXPN+/xurc7Bm/TXU7OuZ3+orHkffy1v9ZPpn
G21G55G8+EVM6EPXGETc4Ru/O2k638sAHxeLZT1M5TazC/N96a4bjDnKyIYheWHP
nO7hNX1K41MUnq1TOIai9g==
`pragma protect end_protected
