// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fMytIrVxd/OIlKLbkAysDTIANIBElv761txzgUQC3JNmNBENVDnAeiCi5v+HZ7Rf
aaYbc2f/suL0EG00lTWECXEpvi6EOqyLOU0Glp16P+ogtM0jJuZb0l+nQDYz3Tie
MiXn/sPwtUcJS4b1yhqeic7q3Rw35RUOyD7CKLPhpnU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30528)
oPpQfgeFe6Et2FTcRPpzgQxXCk1RGQWxKxe6EJ8Rx+QNBwXD+E+KuLWOdHjsBMVr
fRs7PaoKfivqUr1rQHK7aaTsrKjOfWTeUQJDdmBM8mGulsXMTtpInBvpW7EDdSRW
9T9l3MNTpbjfSJGRCM0hluJitYBdJWbb4ylN4rDLoe+10VQ+jZUcgFvV/VqlTEVW
F7biP3/rTilDZtRSrNG1AITI8jCOAD3Gsbx8GLbh6TCeTLXrvC39BgDlo8GrAXoU
FhhLF+x7yikVebeex0iABYjiZ2eER92FP15RI+KBoNixRInvgBj5C41Gq8CE2Kmm
q8+YF1Vg56vAmXQ0qv7p/vqsbPECrJJdO6BEBGFh3BwSWvSmLmIjHYK715n3vIwh
xTFEeg1A7qUNyfLGYi40ajuV30kjlYh5axncFSRv4ADg7n/Nug9IsyIgKA9RC6Hp
/1hboQy85EHdn72f6/YC63IIyFyjb1NvOsEWY4toGZIYmj8IetrmdA/rT9ppH4qg
yRfN76iy36AGurr75Zrv+WE6bI39YzmJTHDzrfr6tZFleILm6z8JJ9b2ISbfH9ur
LeRfCM793aNavwWp3qmUNfrTeIbhPNHI538fLINiPtJ45Sj8uU0lih527tIbuQqQ
ldS5faVsrm0sCeWtDJJqE3AeQooXMhxLo7+oEMx9zbz6cr9i5K0wFVgR6iNh9T7i
xyJ3l+GThsU0v44/5G5p+Tj/rAtptZ/gf0txvj1v4G4eEjuWyevyBb8Si8JJaL3r
XqzrVM5m2OP2Vao9vbzGSOMZOp8Fv1mUI0RN/UyM9o8fkY3NUJ8ZRgHsfF9rkbii
kAoJJBT9MTMEjepL+33PO+9hyWlirxUerS4/D1U9DP6shMi88hj0HXuqr5Xkr9So
ZUZZDN5FN4fVW7M3U1rhhjGrrBckuFPV2wduM9RyIN2l0sR890/hI9sMYeaDAY3n
7h05QPqt67fUXn5PbgX6HN2sJrx8WQsVEhrasLEOslmW8+1QOKUoNpvdlomje8HS
bN9z1qlKhUIWC3oES2NdJ3w1hYaK6BPZFRh0yzgnp5iu1HWPGlkb5kcKzh+sCftD
yc5Zan06XdqSkgi7EkC+o1HTHqP+7MWl/39CScm/27uGkCkVcLY8RbpYFJlsMd2T
PvBIxIsvZBptU0vFTZGLjSV/vOJkruD2zh8mZGTK+1hcLhovBFN9VEGIa4daQL7I
PwTN1oeIJWLtU3tw8wOZUH6/Cs3zzweWzdGG67lVFadeYuxn3aL2tzmRnKV3Tqby
nJqyVo5C5m0nvnQs4n5n8xxlwXyqi25iRXKyBnnyKYmz4L3eCiWl4M7Iba+Tl3tf
El7gNvJOZlDF8O9rYP4rDr6mBHJkq1UuXp0FpX/TJjpwJl/4PtZv99KS6uiOZs+x
NhIScTkyMDPxf9ErcS30GVNzAFgLG96aaGXNAlO2983dnkGw4kbF6nhuJuygHhgG
6QeqT78mTADDvXkj2cWs/Z4RxHW6zZ3+Ue8uw5XrBAMoLFtAKh+Z0qBU1UnCIvMt
A0ME2fpbY7fkpHzV/E+aGaPwkf80V4Vus1B5B91/PEdX64xGuN1HXQ9I5Nv6o/hs
xBgndufDvoDgXF0CpLgZqR9NuTE+1zYzp5VDkAGsgxjY4eXH+RgrRCZvnYcvviwW
B6g4Ry3KH2TVARiuu5SgZLa6jsHYRUfoNwDMRElgvlUldSYcEodUR5f0gKu18YYt
b1cp2lX+OYTApQZB3SqaCI0ajfhgzRvjSwolS8gPsYwbvUWAsKTGIEAsm796/nmz
j+tojUtx3beeOKhMQxEFlh51Q4MvXgbkXaA7iafZe9GO201I6/F27r6QDGCYfEJX
YQdseW5vILmwAavAnomArXuwFI/hYEbHnIX9jJaR9AX32h/7j3UvPBX31WKiNj6U
4CKPUkq5NNBPcqsSXxjd2gjg5FsqDioSX4Fa3wu74bZq5KAHM989yYd9pyElCKa4
HpQcC8WYmjgx0/7dQuIXlF1EjIN4iofuT5O3BEaI7CTF1yeUL6xuJpCLuRQIfZiP
H7l/KeLOOLckUxspNDRskLkiFmEx6g8iJVoYFpuHHqEdOPtFMbxwuKP4b09UeTdg
FgyRbq8K08jDZCoSoZCyGneDabbwkPRrW0YoqqVit85s2x7hicVbmBSYtNrah2mJ
kufwHGZZhOzhITC3LODCuevy3Y4AXZO3jzM7fgCMg40uUm1/2ib/+dT1v3aqudH5
pTtgS+iTzKt1c/54izZc8u7z/kJmoXpYtxzwhshF7erKC4YJemH2XFfzZPttvgSx
YdKvt9E0FgP7DsfydtkmiT/IUGgGhbvGyrnwVj18M9XmKoEOwNrp1Tu1m1Q5o0w4
FDRTvGitK07ZKXtjjjm7ySkcsg+txawUASNs0RxkXMwZY6iwQGdyk48vtKTu5vwl
seZy2PntI8/T5OIf0gnujo1h1nM5PHu+yRuZIj1mnQQpdwXiUv42U+j9jcbLOq5o
vJe+ouYDG1vXThisDA1zfjBKkr5RfvmkUT5CmO5jtmTjbCgerZqbmBSU1vczwojp
1RiU6tJF3vN/hac9L415B1rTnVJ4nbiZuCcWl61Y91tvXTCtyPi8mmu/hND44c7p
k9TaMvqBkB+qsQyDjstgA9+cOYnq+4gz86dFxSE1V1xIbBjlvrJGCU9u3BenG/tg
EIkW0heGxbogLhSm6YGgzeQBURc5hDrNYVwj3RP3WSKnjw7MhwZQll6xux90tW0u
W8WH9BRbZcF7eIpL65744ZGOPQ789IY5B8zgZODurj1I/fD5FiBMBnkE2JjGXMk+
rqflkcOOA4Ho+fl1GzZxHsNLGrfMYkiNj2r4sAdqc2tDgC3CmGH540GhYwFdM0jU
lzknnV28wwUNkrtsuhVgZZgDWrIzk/j7CmFvWM5AN2bnMzADFEVWnNUIxCPKwNYA
22pnd7IO5mc956Pp68FVIfs7Hm8G9cr9Z9S4oBdseiO1irKYb0OqgM51ma5Upkjk
DA/Rhu03zwC1FHJN0JQ8oQOzKaWz/3D1KptEbts7zTIGuVczr1Lz0NQ9+AYI29xf
VfFghznDwsDSGt3rfRu1AtCr8nuKbdJ0gcrk9bowlpvLjpQnS34Ip03bmnqTJe05
4y5wIqEdl/kQ7bE0dZ8nN8oXlpXm/7iJuCnahG9/r+8o/olE8i0t4nlFzwtOFS+E
ykuvPyfvJwVSKEbgSkvnVk8nVpwaQQXx4Bqu499U6SxqWXXFTebKWM+da7c0rmfg
Wg1PRcjRsterfpphFtFFFLjzEjX9AxVcjJLu7pyjCBql367/dHu6lIr2neUYZe0V
O6Yx5MlMEUPtkw6mii+BpRU+ycoyYro4NWpRdvFJSVNow25ss63Xd3DRGNRjaArq
8qD87wpkXq5j+/QDOEN8Yej7kp4E5I0AtzqTu0I1WgB36Pp8AHn/Ec3nb+wEzE8/
KW9iFgCLxLl8Z62GVIi21knT6ROYESbWe4M6mCudzblKLnTkV25hx4LLF+Yt5DzZ
EFuJTw9kxHZEz3BoiQyO/TgOO9mv0IIFzSybiHU3JPbo6vmACFLflJH8b0Kk6hfl
APcr3tnD/d+/VicvveDQKXzmXzCsJFwToILSYst5zwHEJ1NFDD6gyubpqm8fa+3Z
InmVV5YQWZLBRfc2U0eFMum63Pzs6YnolmU7RSRlp0ukhJiDwM2b9FviUk58Hj21
DIyNQuvJ0k/1lS0OT6VWXjxyjpG5n4x+8c/AfeFb8gBwHRj9eeY+fS0lB1qJOeu9
SXgvTcV6Boa1hWtSp59xK+S4phMcQAqR7EDuFmJzRf6g2eVM1xbm/w4UqnnbC2BC
vAPdqP+6lY4P1K4HCsc9AlVosnj9BpprYhMOdX+V2gF+mMdVww9nwk0pjPM1N0kw
wZD7Ki+AdmpyOtCeuOtIVFt3erKESOdiU3F85ca2T+STOi3kntrVvILxYQ+U5xEu
qYvQb4vrWbOfQ07zLtlU0JgobEcQFdR3p9i+Hk8Il4sg94a+4ElgfHGxRcQ0g6ll
6PmWWDMrgmIkl+/JOk3BzJvHslwU5I7K3iQ95I/UMYlDV8Dm8Ph/jskLFtDMTCz1
n+NJIFe1xV5qmz0ouihPOELZO1CUbw/AzrswKJuk/LqQn+d/grjPyUN8vOJ4gnXx
5Q9nEwe93JqwS19OUKTY0wypjOTBKGEAqWGSs5c8VBYFcWkj7C/Hv0WIneLpuoka
HnDVqS5vT+YfmH0GNwaeTZZ2DOmTJ/Z5ysUYbQKH3iW4eHiuJicNG/ILLXZo4AJg
K3mbPXtEPaiXtec+p8kY8jfs9eh4vahsWYN4SZzEt18Idgwoo9M6Hzwvt0QufqqU
VNB5jhsgVFbvbn/SWjN4bai8vfq1XzyQa+ITFaN2Hmu0/WzYqlzt36RSrqai/EAh
9AbE9plUDwCVWNYCGDho25Zq3ssoMRKUi80aJbSNAjNrJvGidrS/wiSo3Mr3Z1Xd
GgSd6G4ojOAv0zla3jtuLQisqYyk/fbtO4N/vGVb38JBaJi5T40wfA0mlnw9tsKi
wnaSqj54nU9r2tIs7lwy7jlsmxgSaJJFsoXg5mMlueegWKNClNepO/zQiN/2XwQS
V7cGAaF6do5pTxiMxs0A9TwyqZ9C0x+KCPAIVQD/Go3aaDzu/xEWTuw8CeBcw4Sj
tiDofEBfnGQZ1PNusW4EZy4IeEodf+eU72GNK4kCAU2/BvsXG+cU/OBUcf1hnaE9
firzXDVwZFkI8qkRrlQYNTUvogTpTV7ERLRqk5/eEat90Nq5ZdnNjrAgtOWojq0v
9lRTjVWIXmvnVEsEJFy61Zz0YrYDfEWRuaJa9t0/jKXOevmndF1UJudi4vob0jvG
/JhNJ99+Vgk0eZw8AMJ+tBgs6eNHFzm4bAKWyw1hTKJTq0124yiY52B7qFZv+GUh
PGdcjnk84pvs3xNR8wgGcgSfLvp2BP1QdEmOlFXPBDBNMUjdFanGKOauvZGJoDpa
MWSAM67hgQa9Om3BdkBlhk+pFDaWl8Nm9JV2IC0A24B9s4VrTatHOCbflCBv2M0L
JNSKozAbpJvk22tt0L8LLu7O6WwvL9dEDEFfHgxIj8jgXMvPMEXWKYb4o65pyYnG
+HDE3s9xeh471YODLIAozH2gS0JM8lI1wjdp/776pvVZ7MxRD2E/girdzef5C8ne
4r35E5/Z0FVNsp/ioZs5LYl570h57McMXsk1EuBS+KJwr2wPLaW66etsrU1gpj3U
3F6pHkpRfjwQk/RE0Q0ww36LQXWegQYpbpKK33qX9vRejJBLE+ZWR122z5ZgiOxW
GykaMETY+bSqHMt6u4oTTgdmjv/W68Dt9Kav/LUJ+7DDd5KR4MW6OUHJ9/K5wYxS
KMBArfb3q8rLAD2Nkr8XG0QFMVHaoZLcMVaJN+eGkJRTYOvo1ldzdQw6fmK8gn7C
dVflK/EUNLusewD0PnMl61rbrKUuVtM0CDsXswynMmFxVWXVE2RGd6x8aaVlX3Az
/v4hKWOPvu7mSRMgT1yv7Esfw28Kvv7skaEt6FLuuGr+WZaKl19ZYan6Os9pGnbW
XXQL0GKg55z0QFKnHGUQSDjaFBkKbVMROm6ZcyGAjOUGqhh/hXUJisqtG+4N7Kt1
ZvgkM2kKkqP5Cm2xvHk9hZCzmCnYrzPd+17gCuM1thU11reJVnYKAUuYaBDj7rH3
ohTSAlk4yUBe4App859vg3hr2E58S8MVodKbuab0if2q27xvBShBz9Uzwx3VEEwB
vIxZguwQcxPi8LtJziFHx+dVX5JLNzn1V5m4X7ojPfgJ8K/PuGox2gZZEO83NfxH
sbFAWUbcJf4tGwqgpzd9zLbUrKJYxgY6NVt1QV2al5zbFA4DJr8v2g4p9OjW1WaG
qOKnKKoq3+g7IcCD5pOGw34SYJB9Um1K1q4EpSXoULkdIrxF4dj2WIGfYmHuefXP
vwmdODuX96kQC5mkKh397eQMoVTKjgQr9mqtoxx+FEZyYLUA6JRyBHdGgUcbBaCu
NBn7Kymgy3aLCgc0XcWIOTkREqiR0xvF/S4k9TKpy0mAaTnoyJq4ACl7cvnYd8PT
VWIyJOHEV+fQd8TZdt3i7/st5lG4lXUHr6oxyn1AS/2xON5Vf5WIZJDFQtwAPiiO
jybt9vQTNMjBs2xOEYVa8HL1cRLIBuJimns+6Jo8D1hVD0FIvhJJV2e5DNlKM+/8
ZTAXu+SrAfK+tR8mvVUypgDwrlxWoOLId8LqEhqbcurZKeipdLntZmFY2QKGqY7I
x8Nxis1NqY2d6KjsEj1YZQAvJFpftPdYL8Xejy7+VuC9dlxq0nwkqrsgsnm5YbK7
qip6jgc/c7y0cvIgcsuCXNFDxSW8A+ffH/J+RrUotrWEGIkuG++nwhL89o88ylVJ
fwTm4A9mwPGg1zTeCtFXBWngExEOVEQW1I81mrlMTM+g2nGQ7prodzz4O63wUACe
r4cKhT00Sj/J6uGz3WJI5nx2l8xNdGZgWGQKr1FnJrDsmKmtCws9rN1hdmsShKgX
T56V5MH7RCVStwP5cEUpQecsJ1JdxG0cY8SjqWrsXxYE2jyPJNHr+igoI3YTPEjx
N/h9yl+DYwA7a+4b8oZhC64zdYptYdm5XiRbTKEtQSc++e/PLxSba6VcZ5EBP+kZ
2k9vz5ORJ6u9WR09TXJ1gw7QrBzwoXvnQCn/s3gLlW2baneMd9iLJDW3JgPqTJHP
jySuW/BFIbE9URh1TmR6XwP7RS5maQgdFbKzN13Yw2N1cXOTtfP/qXLOs3NcVqS2
PGowkn2zFPnNH4bHUMJ7nRkzwgp+sCG9Qc/JYILUhSuezkuYKl6t0MsLH+8by/UJ
Yai2GzQWOR1p7DdLQ7COKV+gKIuuveVI6mCCrBFXK7kRlwEyyqQFMyx2t4BdnzCz
xA4Hg91ZsyDzgjiFw6415xvOzeq7e2sphpEjX3bdt+OTfQmPuVvGIsZEoykHPtTT
m+2YYp1clQ1Y2V0Xdb5ZeI0s6jyoEyAftkjLg05cgykEnY1TizXP8s43Yx9IUPHP
Tm7TNvJGw69aTSf6Nu5ttg/iPAz83n+B56Xn6bj71U8PV7Gz8fnHfQEUiBQnqu3b
lL7RfH5QZzK9M4jooKRNXSblLdkKKAHTo/uXGlsHTbeC7IMUvq6GFK18cUlI3AZC
EKMQOMD63hQFtNqOgkLjBHYIRAzhjrmehTY+RU5nci18rcnzVZTWb2C4nh2E61El
6KSyxPhl3pRcFkbKlDKOTDAAgxriMVJtcdf6ztYhcBzYZo+mnQ1LUO7HB3CAzD4l
Qt4a1R/1YVDzRX6cVjrow+B9TP5JB5R/KlqtTzxxbmmrl6CzYyeU1zKo5wCiEtna
zqXL/yPjHDmKKnuHdXi14wqQZuRIaIy8Z8FpwDSs/MkUDzDG13Q5T4oClry1JecZ
vMWluz4FbMJMmyVPfqyfaCKuLkKMTh+Gi5xzHqQFZNFA9GJHi7qcpPXfhMpDN7G6
R2tn1sqhDx2WGHY8jeJElm3QcgYVKJj5JEuRejvqaSFciN/iR6p1wZhFBDlN70c5
NKrnTWaDs6lbJf/yxTOF/yubBTeijqlczACrM5Owd6oUVy0curgy4gNOyMLWfycx
UZmxV4GmE7bH6L/l4e2QzV2RQOQD57kwwZmwHNq17NxL7n7wXEw1P9XyVA2kk8va
++MbJp0XfC2au9of/NHYwy2pMkVdQNCW2K2bMuCompvkyOLgW44/YN2P43/xgiuc
3k9nr5zm6JE7MGoeQHiIk8UpwpZ8BBqPoAb6xzZ9yv6ATQxsNrITGSh1q7wcFCr5
nedubEjeyNx7bpj5kMwPBPkyQlafDqtnvrKs1GhlPq8IKviFDq/N5Xy2LjMklLaX
MXAe51YX0WR9zN+ubz9vy/Q5PCbFD7QrOz+QuM4QR6Iop1rMGdApu5jxbFlUmL86
Z70/0HS1YOxOdGjQJ6Y6p28/tTBQnD2xukfacmwG8vMH5ZqIJzd4uovC61aqDIC9
8SlgZidccVAnMPKcH8elaQy8ku1tRaxIZYILd8TYX41uWG6iLBFp3XZl/MicHsXZ
SuxsZaMcnrWTkCIX070ZjknFjpfsUQAT+DryHdksFVL0EEeGpcy1eD2GSvPZYbS4
zwseNElnBNMfARXnCBJ4riV7oD53OzcMSpCtR/sFI0EGPNCs16ZY1+R3NTQGKxsK
O3jCdicmIezTyZnIUo9ZYwXoqfstvOWg0bfLDJx/Vh7oFp8RvLBfm4RTO2FP7G6e
BkBsgUS3MVRLdAhHBsGahYi0P5blgE5RtwODWXnV87E1bIgg8TmQTSC+JYJdDMX/
4Vl1Hr4vjHOQk+zNqHRhCtJuYtWxOAZ/DZOmPjILIwXGBRdKWV5/6HyMj+hkeYzf
UzCi34w1T7FROy7OrQX3ZsOZFyDzDVXXw9rb5CCeelFPj0uJZSFlrotLsWsiIPYY
3YOWEtN1YSy+wAOXAkJxK2zBTfq9EhhtmfdhmFUNwXTt8aDPj34rCpSxeLwLBZhQ
joiCzkYQylBt+wYgghOIbW/4iYsVe2yAwBn5P2Yg6EWoF3IftaDdEQnKQGcqsT0D
CjvOXk0DdUT2G6UQ/VWZpLYolRGEdSr5r3TFy+ah7VXAHTHTpxwQNbyKuf9SyMuI
XawhmJYLQxscmkT2DBKB/g7NLrYiEp4cHmpKTaDugOyC4oltYFNsT3wj3JHVtShi
XCazBegAE0ct/YQZUdz8kXbVf4190OVslTKAvz5dVMU/4ljBNFfZSFfaLntruvFa
redRW8QIgQRii5z0+eXvwsSiWhlR52rFLGb8LZwpa2nv/zIMmgC0DOsRcga+b8hT
WR7JQuC0gBV6ilYNKNRwy7DQxbwwYpM+DgfCxIIsVYFb9ZQKXVh3+bMMBcBdXtS7
Ssu2+HgfLo9oeW2pB0wjuhh/vG7SoBPkSmKNTdCGdZ/s+afkk9VNgd02QPbTvRlU
RuYF5rLQNLwei5M7PVg+IHZAszNcFik0X1a4+A2WYNJaIcLzYhqk/31HWTIRvZRG
DKOxz5+yWJMkAa7JU+kYccNLSndAzrRENY/u/DW6P6LIXyhhnE655Dt6V+3ATaI6
8nQWOUURl4FDp9DRa6MaJMYjNAdcMaM7koqiABfc+lpa9TNKarZybqHFtjyS55Hh
lzSrEerHkYabIYk+W7JvbvU4J2ds8etFQiaIW6CVcjMEqK4yIh6U4kf8FPROnGEO
cGFxQP7upKE/vhtdjsFV6xmoDqXY0Ek7KUM4WzMf0THdorDYZZ7qvO9uqbZYxyn1
UWv2xIXDt2rRgvZEP9JC3BF5kOPuNjMuN63ZmjoE2bG78NO34tFdsH5jtgeDRLxj
NjvYQFZiyhPESiqvFFZzkUQg6mGfeb+uuEaz46gCBqhCkK7g/AFhhRKm5Z2M4SdU
hZT9lRzi0Ep2Px6Au5SFepFhkP/6ONPQBmkrVWoJDGaWa4oYRl2ezmFoy73ddBxu
t2WNDIlKKD8XqRjqXd/v0EMU2H9J79WwX+pfz3AtGjmorEvUVUaKYVzWa+XuGhQj
ypaNfcFuDPWFqdhnGIgJIbgEsBU8f1OzoQPQyMDnzAPqzEpCBgwqgznMEmJ4Oi6U
YTwv1Xha/hshKL7WO5DOq+rY8hWkI1+J+CyXyIvchRWlwHIDMhkrwj2U74mvMF3E
Bl04a4ub2W35+b5iDOFJCZ9QwcW05VpBDzWJLSuChPwXVqcDZhc/RqnDw876gHtT
w9Qrs1+Sn6F0Wdf1ElvdiGf1sDYUbkFFi0PCFJ6r6PMlE9jjeiS1sO5lm4c9Qcy7
0ABbhzpffe/+p/IQsI0is/hA3KsXjEJzZY01cRZ+m0NbOXBxgmF8i13GhMrhtbNm
4pP0DtjIsetZQbocB/wuk9bvJDJ58cMTmwBgD3il0QAVOFRKqHJOsAlNYz/5YPY+
nx8Y73B4MeMDONWs/Bjlu5HzEWFyCeZ1KMWXmRy3xWDiRda/4uAv2SzjZtE0+8jm
PvjDIDdPhMx2HbcDMF6Ew4s9dtWPMBD8W8pw/i0ubFksgnfX2+PX/DDg9rPobFhf
tvPOS/h+2wItriCeMV3+YTnrNAULZJP/v7me6v6FTeP6QDnnkxTkoZUAb190mYno
5hbYDKEQdU21QW1+KNpWp7oA+pcpnfHJ39dPMt2I3wJn/VdRXyv3TAeEwqcYBoQM
rqoMytWX371oJZVb52ntc3pmhV/biHSxm5X66GHLp7snPlkaAgkl10AkOtIMTksV
LMCYM5JKv8DYESUEnYS2q5wCnakI1+Rz0QfXhXsQL3Hrixcz50coKq7cBixUNRDi
piSdFegh/Rle5FgUZpHRQptjfJoUyU48UYqpf4XsG4MchQelDtwgLHgQ6NWIzc+l
vTew1pdNBG52vq+pp+J+dT3R2PkSRCMt9n9yxfhbu/SVEme1OEjMzH6ucFenuyd8
+Ajpa57uqLOmqG8Vm3+pZv0YB/W8J7gJPNCjehfr9nMNQ2Lm9wxCSq+AZ5zl6VFd
tMxiV3KQmYkuxXeAYi22CvMxgSlmqtoMDK/Cbv7Wv1l5bMjd1oPm0iX3Bw5V9mlg
XR5LNH7T1KEtZiVvmJhnu6rvChOX3iIBvzymj7ewFi4qmFA/oCV9OPJCPOmHdyJc
4dEDmONJBXeubqxdf5259O+haJLAPUroGzBY0Me4Tef1ESLqA3FjGZ11CQtPbXKC
y+dixMF3BbH4Mdz1esLPlb6ZZs9m5VSSCfW2ZDkGC7mMxDRvxi3ssj35sjj/cDet
le05ahMTjeiECiaFry5ZRtCy/DQnFAEGleUiVyF+mrMxXe/r+iR/1Kf6OyxvCgBw
sxZhBmrZ+/s3epKywnwtlchTB3pxfKE0vK1csfKNDjMhUjNd8p7rvTKU9UUehK18
ExKTfB2zfBaJXrE0/0F+7/TGpUtD1EF+vywY+sJndPZ4B1V0poVkDfsqsgnpc0o0
PUeMYMIe9Zw+cYt1P7jiKmygpG1p8M6xoa6vMD+H1sSJIMYtW0tM0ud22vwryjgE
7E3gW2+nKCJ0b9+/5YuU+0319fpqXqfh81cl9aCLiVBQ37JfgXApHpAwFORRmREX
RohqgQOmXgUxNSyWjVEvQ9vzGsstk/GqfryNydJyYkpRDEqz6wIocHXDc626rQYd
bUfaFQ+Ac7zdn8EVydu4VCf2fWhQal3atkDlhIwmrgA80w1BEscXTR+OqNTJWXXr
J3oWsoB1QMJ5sWf43gpd/uvPlk0B+VEtcaZTUH7qhq6Vi7zmL3xzExFLkdi0mIQu
p4dF010u76+nkTl4ze+o4dMmBWkSjumT5wlC2/VgnDKQCQ8bLUjpO4SymFJhODJ9
xQwdWEtkBzlmoZt6AzofzWYkrIgEWRS/HKj6yVjchrbKiSZWQSbvDdfHLlI03x20
vt0g7TM3L4Tee9QHml7qaYMPIBt7YWJWCp7Mnd4OFctu6HAtX5CLeO1Y3MtIlbi3
2TK6fQ5pLu6Tl0/tufXeqGNv88UBg5FBr1OPa7mgkIuwTF44KXGCZxXUp0tTUD9R
4qnL8bBqvDKODCTR6XA4XqWcGFp3O0lCLU0fgwJzydNfMj4c5h6lulPB9HCUihoP
wL7A2jdPl3uaZglyNFqhvOluhuA1hkb1uY0Vm6ztKpQSamGwBBE4ON5AvSjMFC3Y
aS/nK12na942DUR3YEoegmzFvqYKVd9f7Stgmno3iLU46Y8OzZv5Kct2j6+9IAoo
JFUjGC50JTTTZHOUVKX/ocICpAzZ5VycfJpvh+p1bpKCJ9boaSGCPnggqVotehNY
xqW3AdgZy6x/IctwRzHD9ldFVUEomgyiSVcV99Br/VGUUcJZnYHeQSNojvj2imjj
5I0Ps6dBCfYFa5fBwY52yD6x7eRrI2Uoe4tu9kCgmceZw4oM3XInlNzG1N/aYu6D
rGHmgLCg2/dEPT63AbrW7WL08jdP71nqdsj8qAsonsb8HAGw0Zlz/O/DgaRLbJwc
nE/x16rUGQPsrBev5IOOpuarnDtj9m7Gv539DidCBktNzDirrj8YA9JYknluUPif
Nyeg2uvBBRSoG+8i3hEzq119S3OC9JqFEG1+oQvFPaLY3DAHHtS4YXauNbtSj+ma
t94UnN43I0ZWpC8bCvP8H5UeSJd82u1ee0gGMsVwZ2G4VDaoCwsavNiXvO9pw18t
NWko+xYnj9nTaecQHj/ve5ZHLE6DbQFQ4ZSqchLJcq++a3mJ15zsewgVPDcorbo4
2EStCUs8XjxWv8uDKYyWJQeTLajRKTHm43GAqdt6DpxHVTl4odSk5qq6JAq/1sqd
k6GKsSNl2Q7menqB2QBvrcOoRWRQ8CbL02RVYnoDP3oCSaxI2vGkvieGpIN8H3yw
3TwUhj7QsNeiTtwV/QMbcAzEUxyi4zhYAAmUrwJ8HmJNEji6swVBYMSAmSlk78pk
0Vs0AZmjphrLzL8tZLQCLnDvH3ZBuVdcVj1GWzA63jy4ZImUjdjBgUJGXBiEazjF
1yyBSRxZyp4TwEcrVaudYRFIeTlsB2eFouv5QxOrOI8Tl/X6THVg5nAv3r1lEV51
YcyjgvzMJlqKkGBQBaj6GwhIKHEypGCOhrMzBGpsvYbPrHT74LB/ndFSqaRszvvQ
izlBsQli+xqeO/Ui+nquKV5Dq7Jt8/MAKeHBoKMxBNPl3ZRdE+Wh++9TEjyw9w2W
MowBzG4aSYJFvAHQzxtfyIt4M8qtUVFqEvFj83jAq4uLBt4rU/A38agLYf7Wi7vi
2zzMk3UO9GqVD5wLHAMrYXKe/m5Cd7OR6M1dJvy6IkJjzUzUDB7NpSt78nrZV+FZ
MkuFAHuN0ashX+eCXjoGP/2nO3vefx4NJtSqeEc87VCPzyCJQPYC3NgOFtug1qIk
Pqv2SxyABWV/uqBdWKcYCO90k7REa4gr20NTG7tdyGnyZPWvyiTTeaFLU5lv4Tf2
rOzM7h83XwNWxr/CMLnnhHYgvgNFuv5doJjRzKlbaZmbbm2lgopP/c7GWPkyxa0M
8nqX5dbuOT4nzdarGWAZH6ijTw6dgIOQXGuU/FwhIPoSyceUu6UUTG8+/dNUtKMb
F4GtO0RTE+GFQBZIsWXhACxwMQSzdtSO6ECwzMgLUAwQCmADeVmrdQPnQ05dG3Ey
tK3Gih6o7anNq9U7qLWZnH/JONj2JT5Nk6zRZdst9swdOKeRju2ZtPBr4BmOftK5
yZxuGmwJAtfiXZ8hGseD2kW8llzMkP6o2zSwzkity/D7sNPbf8ZxuEb+p9DIKMLw
hKVTDeNmDrimxGL9k2E5cyT71ODPT8M/MrJV27E4V0WZOVWA7ZjVyxPf1/0iDXOz
P4c1h2yyffIMIQtuUXbbh2vtO8g1bz1zUOnNeLBPX32J0pWS+HdKtIhd4lYkE+gt
Nf+11oZRyTc9FFPn+qZ3RRd+iuZ4Pj4X7BGuPVrSnMJkS00MF04rcEQtgyGY8OW6
yXTRcCO1FY5WNZzmU5uJSS18pTge+4XB+Hnj4IMmw+8xkguuXmbKC5trhqwRRtSC
qnRw+v90siE3wdCo/VYGY/kBWI1UFHX7ZsswKNdgzT8TYar3k8iSTcfb7kpNZlGg
fwXKU8qLkk290EpAg/Er+ztJcXyqJNRL+TLM2KrIBcoob4jZKgFVwGH1EZs5SGoO
pksMMGkZY1G8AHIrCJ4BGpT9eogGiWl1cXh+I+CpGVktWM92jZJ+D9CgIc9ghy2r
gFDRavfGR2hHClFuEJms2Ly/rGoJ4D0TqLPvafLfWgd3ZW+ycI2IDqOdyroTQwdq
rKGCRMOS4xr240wjrT/hjXK3zPIp1AUVVNdDBDFPawpCvWd8+2L2kROiCufY2sBU
wEu+O6+PSULiJub8bnv8KPUh9YfZ1bBlAmY7JyYo6EYxkhCFwVEeaN1RxafLc9R4
kjSQesovcAnRGnZxfGMuG3WoGOf7eOpOdukwvj26SZFn0u8reFUDTX9SfG1+Dfw9
pi5UYOqRTlSkTNW68C669cYGdgbMm+KVF47UQOAkL6YCaSxwDAWSb9rp7enRCnfr
0ULP/ltvEQkqhzVuea5yusg+6em5x0aJkDh3YMre61LnyyyJYBYOEmh0XlSa6Lwj
VNnUvJkXgkQIKD1Kza+gpkcIxDIfbJHHIu+EOcFWjxsF3O8nPI2e2Z4cVjufZUyM
rQbRpdg2eMsJ+LvWCQfeZb+bKoAu4ob+ltcDG3AjQUvvBL7EMtC3D9qebJ0PurWH
u3i5pBoPHd7cXhnLIDvITw87avy2NwCi2dxrw2RPuMcEQAhQezyX4OMna2hWx6OA
suF5TBZO4QtdZ85quIL9OFMqgu6XoroO8xpMC63BH+/sOfFqzojVF+JNfzaCSBlM
9/2HLiWntrGBwFgiWVhbiD6b3m1fII9z3uTTB8NiQ9PgsUlY0UVkPac/5iZWGTj4
iVZIG4jAErkAx5ap9IG5f2AqS5x2oZdYLMrpPON9hsDSq0qkYjv5s5Sxnct/5GAv
m9JSHsQyOenaDUoK3o4KYdMVclDtUOLwuIi3pzG7v9srMbGp7Uf0+CGtdF9AzQ7k
Bpm1phLEvfDdolwJAusWDE8gcPdoVSAr6vecNTYdTd6i92zo+0n9vNBcmH5Y5aik
PER/SeRNS8CZ8opiT2aaB8V1/jU1r7pCcARWiBISGPBx0fkSOPLoD+kfgwuAV8ul
5GAjuvpLqIygVFPqNWXH8zURpFseHzb2xFWApaI+6j3Ayh6QfNl5z1L53BQ4o1SB
ksJG+JzxUoXYZELKNIG0sXw+mIaO5YC7cuQDM6nFJxKW+yAcCgG3lnbSSuYNEq+r
YxMTcd+p/GyMwjWoRVu0HsbUZC4Fo93P6zJkAqmFILujpbrkH8eGdGGAkXNix+DW
Kyns26z84HQNSlAxZmsykJwJ/DuiNL17l0aiO+GE1+ebJgzLSpeMiAF5I8EMnMvp
E1YEVzRthx5JkHcuyBGmirxieGWWqbKfgk2GPo/bGHkOKY+0ApbeSiKLoho8NLwh
nF1r5PPQ2yF4fODAw9blNF9tU7KB4b8RcF1LYdUmRYDX4wUm30OqpwDkqVIYyO72
cZRh6/bY8ymnv4kTwqx6DdAsOnhddIzw2AJODbV4J0nIVx7jCfHJT+naY/EuCZlc
qj+p+XV3jHwpbW5eDvhSw3jKdq0kiIgEyctoqN5vENCwZOmSBMNjaDuru0ShvKoM
9BWobTUHw5kZOS8LHTUerP4+ovloiTKLMsWzaOI9nyr3eCJM+1ymNVAYnTtC453a
t0aOpEe534e8E+Ao9yIV6GyKAwdtKPEX6VDEFAga9MqLDXM1HJ+zbCE+JLhs2xuL
Z/ghoIFBOfXZReVY9hDXHk7tBLNXKBUGF5IIGJGKBA9f8lXAsYPAC3ATGq85MSHc
1vWdfxFkyjCWcIW5PFPhbZrju11EygV2v6f32GMT1VxFu/8SJgvMvn44n8m54RJY
kxfSBoR1LlOQKw2MwDCnvjZyXXJps3IzhKBze7Zxu/MZOIhgkFWX2zoG7cA8aRgg
qgj8whbhrJblTxyR/wInaIfR5ISfWxCJGPxq1jO5K79ztN8LWVk1XEdHOwghtWA3
gq/FGtr69fMi2pDyUJqg3YsN5Wq5BiBCBvO2WdCNrthGA46eR5Xgvs1fjFajQhhX
AgsmiRKQIT7Zg5rNcLJvL/tmLu29H8QboolxNZnyBH6AJeh/pyhNKjskPhIMKTGr
OXtYZdMGLH6EjT21amsn9DIn2ibVyIT9EbL6kyK76V3btTfEWiA7LznTdzlnLtow
XLoa+CVS5Ge1l6WsjPs5Rgus4AN/TgVVcCIbd4LFCuVkO/IyaoXLDUeO2nTXfTGv
w70j+Fv05vTPADSpcnIAZ2Y7mehEY9VB42ONyNiRNraZOPRP/HNDiUws9fZvJzN4
z9Qb0iQ9wVMNXP2BvAV6nFwEOXjfLSGWt/NwBYVSkRBHygcIvUv+WaZvhAYH+TLx
tVO1moJ/Ni8W4lc2bp3uh4t4g28jwZTkPjeiboMxrFdMOqo1AosbLWs3MJOtWpT2
fhdH3KzEcWjBrUDApBZirkuB29MfOWrxLMKHOeZ5ir/WH60lbU9MWbCfUveBAkuS
jQMxOsEt+CUTGYBwnH1LAuInHOSj0oyEOSSks4Fh9ed0xp0nieS+1EjiC8OXIvTu
CXvc1YHzfkAziXurX8XlrGGB4HJ7NMDABIbXm3Y/CTOIPGnlCZiSelLJVVk4WLrf
avaOKH6ehldf7p8VW16qYXSc9uAfpJu42koXZWeBys4WIPm2pH+bu/oONVrBiyuN
ibLQQ1Jvpx9j8Z+dFSG3a/xF27xbght8ghdewPs5HdiBSrPy3s+X8bZ4ZX4VX/fM
OY065cCEv4+Dwm3aZIQCI2+Gx9chfMSWhMlnWbxXCck4GUkCqewa7LXmxo6TP/Fo
9siwj9vA7TRPJwhiFXDJEcbJKFVBB8gsVUBzi9dOrqa7gJaCMttYCQ6hHg8TEa0j
Sdh27WLUNtPSw7f17SzT9suJ75KDEwtjaYv80JgwKTI65BnyYHqfZ6Q7JnB7D0x8
Xh+dximVTGdnckrNS9MeUsuiVfXXZWC2i6wYaWHFTlX5Ome0NDB59WAp2K/dVBJU
kGRxIvPZ+Dq0AlNZLC0/4rxWkCdu+mOf7AJOZEiJpCMIqBkXpdvBB/wZBzqTV7PF
duZpej+lB7d3T8Rvxps572VM6tO90UQmHM5UEcDwCMqMjwV00YOEQyf0B1tgOPuV
Bf5OT3+KBFKpvukkwEfl1joR3G2G3cC4rcB4c2FXZzKh+Lr6dp5gu6KUGonrlwf7
ZgYltm3SsmE3cLt2Y7k7iLQXym1Aj8U4pMqzviyAbU3u3G0EM0kJekzwlYukuVcS
iVAg8juwCWeEEM0Y5prCYxHgnzyjctmqSnQstoHlo3wIZ/+Qcq7ofRSEBJ6OAv1R
WxRh2e2M922LtsxtmgNzJvNNX9QDcWrO4Zfu47tWB21RfuCo8WgWGDwnrtfqPNtc
T40QzhXvHZMsfD3g+7QUY93YQQFbZF6XIIokttWoQCkkyft16P2RJhM9sMvHXoEK
LV+4Z4VvX6U+TRlpOS2Sg4uKAHlIejbU6fx9aN9rI+xtPIJMBqmwfSAlJ7Hkmu43
lYCu/PzoTmEHbxvYn9w/sHNCovN5fqhFJ+ym4YJaEFetHQF34mvyGYhqTjSUoyat
p7QxAFYLTn98+sHhFiyZgpezzsiopgoy/a4VwL5Af7DhUSAUvmIIu4X4W9hdzGGM
IyVsaYuHiEKDkQCUbof+OTYb3vT90NCQAXhOxmj6OTJ2XCNC/6oyuzf0Feu+LvSb
g0rbPYl7Ju6UN42lozuuhO+ZQqfLTXr4jOZuK42TKcN2WGs+6TS0bGPNkwJyK1F5
FlW47qXXkRsVzD3yRMp3dcoqlMVNsSSq2SEnsju/iQDUVOtifgLhmoDF8t/97BnW
YljQ6/qsee5tUa8eh4/L2VxTDxR2JEWEptg8KGPZVe4hCrXnkqM/rlutKzzQbvzD
aHFM5kwmkqn/ZsNFlkiH5hpcvNlpiEPkBtchwS4kPd24Gy285bkuXf0SN++WXUIX
RX/CTnA5tZC0qqPlKUsFJ4SKg7Ss2swQh5B/kno86Yk+D4XHBndxBJlJU7wTx1yf
1xOQ0HEoWMHuyP6zfInAjtxiV6wpdkSb417oW74FNMGA8OCSQVehpGwslrRzktED
NkeuYeX0v1jzcPFnJ2UXrCMNPmLRQpwb9D0batL3P5bALx6VgZtZ3U98nQSfd5Vc
CFjE/jz3JeoPH8qwcfbooXe2s1hGYJvlZcXvc/h5gVHlMpWxtfKuRLhOrPGw1JdC
4Dy8SAq+ozVGqg7nvHdYbzv2uczvWDVNRdslwSCjt6MOxr0ClqX/dMTWxEuK+MaP
824nA58sD+alQFP+1i6T61iLOSu9mbDiHu5zz7fUavwurxs2UcYo51rLwvkK7al7
DW+cD+YcLx1WYOIb3GxpAa971Ku2hRmOQBjCIkPXVDGprDu3QuDdTvdtP43rwdoz
Crc4POoRnAEg01X052x8hya97PdtaSEshM376GRXaavQy6QDUEPfnSwbVm1mk/Qd
Q+WAlr2fRG35L/8G8TtfYwpUnmpN0PpVFoo38BaIy8guwTCOhxa2GJGyQc0QoUKB
KWmiile0OPlA+00tYGS+McNyyKfrMU+xBAi8gEOVRA/tdVj6iIjMJJ0pb5ERBzL9
nHHCqD0+GP0tCKm80m94UWcU3F7O5H6gFOMlkZFk/ZUKWGkAAg1eao7xSsHd3Emg
UC3gcKRmLqbCxueaFGYrD+z1zVRUAW4C3MThTWJqmVrxVNPAEs7sz/xV2/lcdUkI
RuzbbB+RoJgyIZDY4Pq70BjxAjzRO3AS6rbvhkXT29z56FZ6MHr0IjIw+1xiZ8xN
1E9PIusn1S7fxU0XUZWuCHLSez1HsIZD+F0Tj3l2dAQQ0xAjpn8QjtdVM+bsmrc1
NsyPPlnPzJTJ6lqMzSqJXp3bnAVWxDx+16r534twYkfATNJ4JqyqR/4VA7rZOhtH
R3pWgIGIm49Kw/tFt+eIfOpIOOzlyf403kzvEf845j4bhvyNCCdokSLoStv3o/H8
I0PHb303NtrQRyRBC+oOt/ZEow04xgX657Dz8/XOKJqdYqGK9KZaZblbg1LeVyoy
cT5t3GxvsOd0MjcRXMs2NWtqtHhAJ75zTh98AR9jNyPm+l2s/B9Vcxz+RwyOquQw
Lqb0YKQsDOWyNOWZFlexR8iU2fkBdR0v1X0o18lV5JMSf40cKPy0hKJDGXEAbhD7
598JrYjYiUev48SJdCLJmqEKMxOb8QBFDIR1yVeEF4ZerahreZ2eZmnTUAKzLlwu
902x/dSKJYt2vP1xZnBsBLPML5HFvjev/Ct67T1zqWFmnu4QsEL9qg7nAiS7Bu8a
A/8Y47zs49HOgX18V0q7SprM/NVcjKe0do9ajGkgJHGODFmm4dDw4IamWdL1Ny+p
uyQUgabh9PclPYoeniDWONp0Ma0aO3zSvpKXwMxWx2NXabRG+4fB6OPcOXKM6dQU
Q/X0hjaVYAdjbM+VwvVXt7L0h08A/l4OPkhJd9E8fTWADmQjz3+Tt6eQcA9C1lIJ
9yc7NMDTZyCo7u7yKHDbiOPVRbk3M/FiK5zVI9lqUZmJJE9jV8UpTvPpfUTCWa38
kRsf68FshqyJnBkGaXEe0gC2ypwJeQb/In6unie0LWysj6RO+heap0xXS52ZGiYK
Ge9PWFQrvSv/AGUn3MZdJe4HKAepYIyt/bICksnqnm7mrDXxH1HgrTXmPF4BjnIm
FCwemdSZMPlrXtbyfwUS1RUAnG5cjvw5HonfaXiDSoCQRL5qYQGupTGT47tIEZxy
XPuGvIQ9Sm9fe4FJ01qc71gatsOuak7wbBQlTKIz9Er5fm07dPlKLa/ZvMcwMkIM
C8KcHcFE4bINxxTGwxGGGvkNCx4HBJa88Y3ajHn8yJgMG8nr+sZ1jQ5GfabbGrvD
GNe3Hu+cSzlenfohhMjJjX6ShpKHz18xqMBQgAAXQDcYkz0DCJyp7al4QVnndCeP
ZQcS2jj34aZA1Xt/XnTxAMG2E2BJdq5bvz+9CtxIAsb8NNDKrWezk0GSX9V2lLNl
H9ANzqELqrBONQCkZPBQ8HJMt0mPCgyvyz20ermWTFouu0Mqim8wEDON2Rl+642M
L+CLRgDOEgCne+r4/YIhFYXKs2I4eIgfmP8p/1Ed4KhIBtL1NDB2aNQkaWpG/JAc
4S6ZM+osJtIaf1CT407iiBAGwEIwdxiNW3TmhjtVtSNcHHp5Zb0KsWQNy2VZKCy1
jhvQ1o6wEjgfRSqdE5yKOixYjMWaH+h2oDtnOZAFIk5/qidMHIuo5DVxXP8cnV3W
sHyfIf5fzcOyzKx9PclJ1k7UNoGHTOi4Q9m6TVD7KmBRCyE3CFMe89rr19wmEMfn
VdUiMu8EkTD2CRrccS9HCAuSQvTCpAZ2670JztuXyKuMP45wzY4+rteGq5sFIoup
42jf3/Qyq9lAEk7DzchLTCIhe8dgWxQv9o1Qm52YpSEhyx5EOeTRvPNS5VboCShw
ajNXGpE34LMfj7HgnFtZ3/Fi41Vm03W4U+S9aKQmDLMCUtt+Zmf8OJWaqwq4qYUW
7Hg4ED982GKd6jrOUp9dp9DYZIFW8osni5r/b5LY15DCWBHqoMnPJ3CGuXKF093/
jq8l7kxmfpZS2ncFCZhmBp4OAe4Qn0AWzEyKnFNxU9DMcnhVzPxiXx7KpM0pTa1C
CBkxPXvIxJC0Ju+LCTkruune4kNRviKZBvJKm6LuGYfZD5UY0TwP9fxyrjZvHHC2
iuKTvH65hcDt5nw1ndAT3le4VhmGEXWeZjaK91zwOQanfKjIwy1F/lIm5/lKfqRe
9by5DScGhHquPybUtdYchvZ+E2JxCc3RLj8+fKv6y4Y8Q13o7OhmXbvfWcu7/EVj
slQ53yc5NJZJrs/xgfHxZeO6eOkWvIPFC5MUjEVgHWUu73wx31UvmlbBVUCAqcik
RNsal+iu7j/G4SDG/dR0N3O1NqP39VcPl9tL+3aOXsyXV0FFdzn+784ZyCf9MbuL
YXNGduCMMiTTse7fzMB4q+P/gE90/ctrsEAM3g0to+HYRAYVJnuYOoWRYbjFj9nV
o9dk8NeTeZ1XLF6oC+isSq8BBlDjJ2JOM5pTQpT3dc32JePRyrWzX46VOyZXs4uE
IcQ4RjPQZAdpOMUoACvmWnqxHI4IMAufVp/IJVuQgoGujjY7qEMHlGSIuu83W4o5
0gbHlSE2PEEnE+CnStDIem4SsEyD+Wt2PNtgcIWQJahfVJiJGz9vJ/iLi5pdoUKe
MK0PK9n/hoMJpH/F62AUjht0RD0+w10NNqgHfMMTonHuFf7U8/mCBDldqkfLZWT+
rRrppZxDP66pXOgewbp2/s4geAi028KkkUFg/QXubRsEy4N0k6/TiSkrZ7LQSFWa
wvU00EFhuBh7Io38V/YU2V4XmfdVHzlNCWgKTyjjbPmKMUJllxC39rcwdFSYkHsA
rrdQXVEUc4OLqzalanZlUt76v9IaKQ0FF4//VbM3jh/NgLJ+w+82XcxF21d5gNMe
pbbOB0Rf/Ot3nbGUqb7J6YvFymCotpbj+87G+E6eDxZR/HZSYzY15as1GsOXU/tn
u8zX9bQAyl8st2pMwopohww8m/mVjJUwrS7qPTMUAkAAoVvszDep2V3wFWMXcoo6
FHlhwcUjS5rjj8yAzLvboTd3h33RrMnGLhzhc0ZywCKkV0vKDZfWCVV8fVEYSCWy
8j6q5t+19oUBxulfoWBaX59j2ZVL/fqtMtyFaMd0w+8Bq341zVYhhtstg4jd65Ch
a4z6sj0jxT+EfxFEQu2HcSIy8LnW5ix+X4PMf/z/LWuzx3BJ/f7AcWLc27hPqToI
TWvt6YCNPrPj8vI439ffoeLD4DKGxU+A613D9mt+SJLTPGSFLhet94BW1ORAk3+X
WTmQT+57NuRMkc4ecctAxu4DHGm3Tka1KvASTTjB9PBRpG/IXZ9NTaCwEA01Pn7v
/X4kbjy0lo+K7nAyxjIU5n85T0gfFAkez9dNRE+AqpgoUDLT62ONVWKCuUwq6eCb
foT3lCcjZnpgZDvNyyKhABskTfopxWwLXIt/G2bwQfwIYdEUKq6oi/NAnZSoccFe
9/EP/0CQ8EW8JSriDs5YFJJkN7J2obH011ZLJf/iLgxjFNr3+XcL8+vhJCfTZgrB
zTRNem/N9ReyjleZUEiDLR0knFeYUJoBi7Ky43DltjD1kL5AmZq1yr8R/YOST/Qj
q82NrFsCHklEAt8v7Agr+zgO7lVs7l3srY1s2XwRboEBJGmt72jOmmB5eqEVkKIw
EZ/gUq9/vpCciHB1ykCHrsYkVOrTkMRuU1OsOE4jHvg6eebImib8Vfo9MA9V5iH7
xLNVOEbkIo0ynGVz6oxa/t5I1lM9g8IoCR9EkpgghzGxAAocnh+lAE7OTMdNIuX9
4gjVJL5ZXcmX4U9RwdgAPuXdGU4DaxmHzcGgghxcf2I0OWDBN7Z4GZ90n6Ou/qeU
PUkBUPPldEjfhTaJlUkDs2D9IaeSgEOakzYAMCe1J3EqlYn/vjWojLkpM1GJiOVg
eHzzrsweZGiBqisQ+F7ZWkGL2u/nbiM+nUEkkGhzofvpU4c6vHJGqLcJ6NlM4CUi
VCAXhsmeCZO57rlsKNLS2K1UorQYoYI0YB7DszjZEbJlDuT8nNWs7GJzHcSm2VWT
qkMOp+0XITWzx+xxvAf+e0ABLiBIwldj5ub1r+f/ICpSGjGPgjk43sFKy+3UsNob
S03N2XXv/pW3r5EXuHTBNd9KWYuKkdS6OtKNAZyRGUmqNs0slbDPc7UcqvQSTeKx
ZhLwF2jSmgmw7uj0c/vqWm9Sc7Isqk3KB5OOn7WZ+yyfKHAQEX0NkiU7/ueCx44B
ex8pmBwZMxPcZxQaO/jupNELIAnYjw1RtngnysB+2JhPMPv+rJkTFB8r/TMIRrjx
D4HsoVGPktxsP4xCp7jy6+VW2cK1msOjR/wE6k5Pf2dkicKJar0ywrcjuz3Zjzrs
1WHuWeT7tSsy7wNbUq11pAsW5bqwePAvBlKYikFufVFUvdeY/BRYp9+l7ZWli/IM
0fLNXbBebh9Mo1xbzyCztO4n+7Uzcp3eqg1LxefGNZbgoQ5c0hkMmbjCLnfMnukW
0GaXQGhW6SIYwF0PH6tVHgwjAQCrfS2fMkn3I3NWUDQjL4PAU8cM0iA2bUNNN98s
kirv1x0lzc8fQ6TtH1d3PDNBmD6VpL5YOquoupdNZ/oU6ca1HCKkuAzPkFeNphxO
PljrAiLW8wIBWdQuHOwChjDMo46QXyLVH3Kx4+9d/zvLaQhgFBLxo9dWgkMQIxeu
GNweohygIZ0i1fwiBmwuFTffBhZ4+w5JGl3irpCYXCrsz9o8kqgma14Wq+1m7RT0
qT3nmVoaDbJbV/5QPayBfaKoJ6AYD5KTGDigBkAlHrXi4kna3nTN2plxLfOVY+rW
VVzKcNAMvR/prd4B0fSNMoWShDiWrrienMNEb7/U2reQ+xyQjDvsAEXSIpmJfjya
I4lziiw35bTIXFF0Fb5/eLxHXnLFcq7lLfbmDMP9uldGZXFYR3MZPlySTuDpWIcc
b8dVJE4sD2cKY3WnU+PLFDZyAeEtRd0K0PTwFUJ9Lpk03CQXwpPJkDhVOc7mVHC8
aiQNuAZYAiYosqr5D20LR9T56cvk6ZH2zx4KL2/c3Y8MCHRTzhOb69JhhS/t0RfA
KnWlkpZUyNH5mYPRGMEX8cmQfRnBbeWf6UYzd0RyH41rNCpp/b32cAcs3ZozYCN2
y6U/o/hQ2xAK8lYBQuEB15yWMeB7l+A4avcqKTVF4t0CyPkak3GMD7v7cpFFg+OU
DNqbRmcrLVFGcKQefu0SyEw4JsKELZWqWsgGRC5hyFt40OxYLxpemW9nc+gbjbAu
OLNjKih3pMM/lzwmtrmC9gEYgjUBSjlc2qcPIwmvR0fQtwDcAuj6RprxtSQdLt3H
oeRG9k2qGIWgRntKVtxsBdlO/EQoIWelZL5FiqkCTg0Z4p3LpbI9M2vZl0brQtoJ
tluJYpZ8zAgMUWF1loVmmuu9J5vcZ2tWqmConaKfqnyHrKY9v9/3qMpfDWqNmBL7
WA3WJ7Ri0w34ZK3EHaQUvsCMdwQZ32BdpIqTjH4ZCq3uT3Y6CorInf4LJkovV72H
RIaFzz61zs5fRkzWF17strpOekrdpv4Y+jyzYbZpnTK9nuWJy4kgFOlskZRdM14u
6PlfQVBiiJ4uC0lc2UpzZAaIk6UmgWj3O6rmGVl8Se06neR6fr9JuTxleNBsVGSM
YXHvf2K2P9rnK76kAZoQTORf4C4orQEE1bOO/RS1cywhaCmruzJa4mz+1uMW6A4e
YiocVeQgb2ZfjvOv2NEEAPLl0Knf38drgHqUxi3T++UnYBD6St/jf8RPrPBCDgmV
/ySD/3U6olL58Vu134cBkZKkZniC40ntuzw3eKf+DVxzLq3niV3DkQAr3LQsFspq
6d2cl8gmnCvibtRucU2sH3EoZofvcxcO07A2NtkiFw39ihgMmAlpWdE7B8gZISJz
MfDl3JxRUgy3dcnjFjNwN00/m/mB6/d8lajwZGmDoZjzIWIejbkq+RNwTi+PwaXc
IOGO7uJ9oA+QL19YL3IAk0gbp+/nWeNytz6c3PuFZKoCfYijUVrQi302VwKtyK46
dHu4Wy7EPbIozvH9Pq1lyvHo+WimgLT5OT5oR1TXwIzS9kM8w+kePNXiqFEFYxvo
OaXAstH2gHSnQhK61sfCCsUmt1rJf2Z3khL+1DihmFoKQz+FevyPhc5T8uJXiZHR
xMSR/0q9yxWEov9j67s+QCeQl1mcN43yBRJphT2reQXcFfGoZ4xUjolhBxONw64h
cOUTSke0JEoAXkR3CXk7zZ4gn0bxC0hbsF43KcyIz+19PJYLQ6CbUBQjRF5tRS4U
IdbCgxHpDBdStm8dGaXBWQlZ8A+OQyFaRe/waEPNBkEn3H+PisSaWFFcTHGmTFPE
adMThJeNsH+CoGiJz4chmxc85GYZYCCuQr+xko9rF5Y2oNlXixAK71tHMuCRSpCx
W0pqAd15ZZbECXDaJXXTi2sOD9jo3p7kzf3Yj6PT43eYe64L64cfXID112C3aSWS
9gA3S9DzSk8ZXjQJhgj5LeBUgwtc6nzlsHTeOyk2Ii8Fk+Hvc6KPntM5HqJmywC+
2kMPmBNBk6p1LVCItbuJSmFS3vQRL/en2kH7DRJWEpAkwwd2cd+JNZdNKfAR/2rE
lxs17MnSZOmU9mFy/SGTfdY431O62cR0HTney60KR1fLwycWi9wDIfEmKvkJGHzp
k7pA9oQehiqtgqlC+LdIcnB0/Y1tToEshaLlpmSJ/37D+7VJRRjffYTDPBHcaAsG
5y7vfv7yRL3bref4oeSp0NlL1R3cNPYQpu5SwfTEiC7RmGXddftQ9E3bfKmtSDiz
6K0tVySjXw02Z/BePz1QVUkrY3XOj9W4FofRUcmJjI6D62vmJxmcmwYErgXfCJW9
/tnrL74aUHciBQw2id38pNGrblQHLwPqQAzREp/hkmSNT4mZAH+i10LlV0VodEWQ
HHt1A/A3tHJSTAkywdNYZ1NeSD7vbLRYH9l10eB2M8P95jWzzQ60P4KNPBnE+KzH
ggClbbjXRtr2toK5MGsr3oKrH5zRjwR5mOKQGacNggKLHW6fZfo+SaPMG/bkpT8R
ChIl60JdT/hZdN22EOdDhzYM/b10t+cRfcdP+97xkAyHo6Uqbs6MZbmEH66zLCum
rSpWQapEQpydV9iijPBddyaj27AVa95z9NDV//mAwrxfHwf15OShSyv/bsQi2aUV
1ZStLCAs2xxppCRtaZRYTtJwZ2oKbJEKM+RXXks8l4pe8y1Pu/BEw/HMp/pJGDUs
9r826ixX1019xj7h+kW8J1+mMxs3Fdq0e07NeiHgcjLBiIhJsW3/3xlRr8f5+cFv
nUAcb2F/mCaaY/OXqZYPhtcYB3Y4ZtCAOFsriQBfFztgOggSNpBFQwRAGcK8XqKE
PG12FMNNK1vlAbnrzSH5CSTQ94lg/MymV2/wy73Fl4rvExjBusvLpDlPSmByO8GT
GrYWgSVK2Aq5PzrlGUJ+u6zTZhxbtusQRVVd4d2QrwA0plDcz3VUxov2cFx/UMbu
VZl9yiLGh5+LapS+XeaTWanaI8jeqIka1sImuisjQntV3VozGfyXZEx+DPv2S4Er
dmDjbaKlr4B/rDN4RC7JrFmbPkeu0Skwg/xqxKlxlfNTLFreQEUahAfuAojy4LHd
LtETAO43bPzEEnUr/NI326gP3RtYvVplgadq4yIdLcMbaehemmI9wwEsIBiq7IoG
DNbeujyaE48Dr8c3NiUJ9pZi22TW6L25gyaP+cwBq8yDmRtRqbzdkelo+6l6xEL8
1u6czbdflXEsamwaSM7/vMfcxno0TH/+NXEl40Kugs8Vu8SGKYoOEAtZJwgN67ab
0pLA7Y7SfC1WnOwUwpxIYtvERSUwsBGf1Yfu2B/dMlyV9OucbC4QvoD61Vh2ylkI
A3e7It5Mzwr01ckEnjtWL2pjTA73OT8eSjRZzodLjLbeQqZBVn5OrJa/DmCUzxBE
FecjfsbdMmXfWENzWgD7+VeSmwjSmLQMZbHVmzNR2uAsfL6l36xf9sY2uoQlL8qA
euNLcnybeUIJSx6rkfpwywLCNfHgrSoC1X0zmPFe7aHtCivfE6XKHyf6nv5DJkK2
Gx/Jry7Eho2sZViOBPPYmR7zUQtWRdesoUMWxXXhSpDebtHsdwMc9nqUCw29BTlz
si/eX0ByrwnPIoityZWiTWA/D2kvk6b7Q1qa0Pie+2d4LDRtVefkxFv9s5UXWBtz
dvE4j9yU6UmtmQ2YGW6Y6fW554lMWmObByMy83PCOV0RFNaJlnnQDNWOEG4N3ru1
KMwgYfzsfmu7maxVsOJiMueQsUnPraagaK7Pz8nFtD7+CzP56HiWDmNOBn6wHrDA
/X5pIQLJU/GVAjNBdDNtaTk17QDlicywYmm+bDwrYHK/WZjfWa+RS5X4knLyJnta
AVNAwqNNbagYswRvFO2/rTYaCaHcZUb4NU4iGOY1WBtNA9DQUbax6hz0HH4vxlfX
LWHxjQ6uHjFDrOFp5Asua9C5jqPs7o51c3VapK/50Srk5n8Ovcnb+wykKKcRv5/V
z5mG1xAi91NNNypfayb/V5MArnPE9u4H3SlMpsc3VNOoI5bBLI+UIkixjPLGmvEQ
6nlCa3/BvN0+ksvQojG9pIoo5k0JTBkPK4FlmpxWB4oTScKdlm5XoqrvOE1I9ovg
1QRHuDn6PK47o1jkKKS1dX1OhKxvN4NpSXy1yAJwfHQrcIeFyRzYnk3w+0CXDgAe
mjg4YNmwRu+gfTzvo8pgBinoJQJPZjd4Ni1w43vZSYoXyS2K1adlArtCw81Cf/Y2
CThcMoPD97jZ7HJk53TGnJIFjOfOUthpjjSkR++ecJHqbZOeI5X/EtwD5xHxlRu6
uIyfJ7LtB35izhUbzNKCk3ezt8tLVYpxLslRjlyShly/UWb7vcZRY0ORLG11PhBn
5Lql35cbrOKB/TkYA8k3fYSvi9kgLQQeD+Qgm1gPTLFVFOlqEu0TwXnp0gCj4yWs
0PbIFBxFSBjLBP3DY0ZZn7lMMiSd61TqmHpuYm4rA8+SAh8UcOE2UcE12aloNwwi
Ma6wkZM5Op4vyfis1UEIESPNlQXVFT7jLyXoHx4BO/Jjzfq9GdK/qXRBy5K01Qra
43+ykmTPNga1UD/9gOi0nBExf1YdLhOG1Y7L4J+U4DxiKg0EwGk7N52bfU/AAW45
psaWhXLojkDxSJXC7fby5G28j0sXC0EwuMVv8KiavwvyRXMqUR/KeyttIkst7znh
thqGwE0D60JLbuGSWmJlrQZCfsLXhB9AFPoomNi+b0AUJHVC9ek/+0Q8hJ9nLY5S
NutEKz0YN5YRjc7xuibFVyuAOtYq0Ml3d6XHXERdrcy1+fmhHmDZJCNby42MQFA1
Ok8tzCdEQNuiNsC307okNd8ebUtsgRg0mWqCFcKwVDwH0IBhNBxssvSU012zuYSS
MU8Yz700QLiV+e7Lnaj7SUHDim/8kVhrpHOSatcCw1ouUp1/1Wyxca9selR5QJft
BDKCof3bYDnOPjovTH/p4/3epId/8wHbCD6aSkyf+pMRB6B0d13SRXmvchBtQdwh
chPBYSUG1YHvld11mgYx/i0Q8B2/P6kYm6ZWsFBVxWusw/kzWxRxMUSb1G3OJzh9
OUskgK0+45b50AApWVJ6DwgJajD22lYtQTnCXodpUgspvLOo8KxjF2qNqgkRUUb2
tRMD1hfmWJUd8AmdEzh+sVMuXgARw3WroVD563Qt09V9H7ytYYf4hh85XkIezI+3
rAQGkai8Fn1i9JDbhxAa2IxS5dEptMYK1jJPOF3cAfWKt6T6n5HvnXG6Q87MLaFC
42pBkcojgXhUodek3GnQEQa+yQ4oswWDLBhVXg8SkV+R0GYeT5C243jk1O/7TTPX
umrZedQrrZ6eYxM4r+Kgd9PCHplxAuoP3RrepBcyO5pqwRZMR3OMgMmIey/etuDA
HD6CSGhQXwozpjO2a75cFDco4NvXbDvBBpN0brd79oERnu75wR4Kqcw7rD57GfPo
ZKj7l5ncUTzfawrv1vnKEcENVDWIS4eXPW/YcRvI15No66hyp/fwSpazfW1k2DDn
J/kB46ia2LUF1mwNcZ9ddVKmkjKqSO2Lyd5xi0kj9eCqdBYslITt+qXmy/Ez7rNW
JNk3mnPQzEQ/oIBk8Mm59YQ29y4MjsQFfYxX3JxAMTRo68Gebdw3C3TwzbVS/Sd/
yc29FStqTqtJki/a2/O6aV23FFmVL4z9NX8vOZIhAG9m4yr20JSxAY3PmzZbQYRb
WUofGiablsRqtIs67yLDcQHZBFbGOFzA3fyHJwg3I9123g7yjhJSwiOmSEXYg4CN
cqseN6qUcVkeGK11rDzneaEYkCXFEtqzkCBueL49gAbIqoWTaxaNs1sZ6vNUrvbE
2BI6pWhGCWKu8rUNG/O344jN0X+uLmvFkDWS+YFtg7ecScJbi2AZwsZl6aJz0YG2
jY0em50yHXkjSE0pealeDgv5gz8wYsxk5ysj77qULoMsh2rQaoV/6naJ8sCc0TeL
OumAyy5RvXgtB9nF8WNuRX7j+KJgEjQH3f80j4RmEv4Y+jOwRQHPb/8grAvQGOVv
0N/Q0WPsQxxWPZ+iZKYv5Hi8eDXNA5ZN4zWb/NDIHgwr02Tkc9EDmRfcSHdAuoIt
Pfc9G0Y6E+Q8ojQfXbeBadQULRr3fBotn0CIPv3RIafu4nXDmiiHk1wXL6tXKkum
+vLFFB/xWH97IKsCek0v8q6cT1ktVSlS1KsdhFVquSBOq0wtS6XK/1lSD9GNxaYz
rWD+7PSnOxJg8OSduhvbRNJr+jhwyy6jRZm1sjyBeZSaSCbWnmGdYRU44YnMFhRr
NzJodGoMHtZfuGRZ1PT0G3PJB2bFASCuXXv3mez5IDRiG+dEOACFeXjFtN/l5v7+
k7zlIDckOYrQsIktSx/KF2j2ZMhScEDpBkCqp3ADCs06qmMDQwe3NJqxOkYRKr9t
PMqVeRKiPyLC4aJT7ZK+SQ6AgUrYwED/jJwRYpkbn36gXSdFSFoqyNC0FsKcx2Zi
9Raf+fKYuqA/FXklahjfwRUgrMKp5hSgULWWDbQGWACYt40TLC6J+t/DvIVJmUz9
IOJmi5BPVSZzDAoSOxBJOlpVA7msDhV9iIcbkL2bm/dGZ2mdaKEAePgxDWzfCqrp
llnlmWyTwoX82A3Ho2NHaD0Fs9HgkouabuHeyceBRBpn8Uw/nGvQhPoAvbGJA1/H
i3GcwEj5nIkShcSMekbWnuOuWWcvsUAFLIjTi+nMkW5OkI3Qod2M0zyPLl+KGtkQ
i46pJgC8dp8lT4iX2lb/VD6ZfRbuba40gtlg5OoyCJlv98gwRtrF1MT3izVr7APS
lloyjIfrB0tBWjqIGMOJcizBTiv4rdQJBSwQORBs0kLvh/tUbnx2512lHASiyrSL
FhmuLAlUonAO+P2isbx4F/9BaN9jiq5nVSmb5/W5B/WvwdnYRB8CYJ6AmyvOTd8W
MtxGLZz3TmRcZhHG+UFvRaJj5UqU48Cp+mQWhQULhXvyEHHA8u+gbOd3J9XwMo9b
LUcxEnDhJiyovlHoFXWU0k6zoIAVSMFX115OfZjfw37JZySe7A+OxkON6t/oQsHj
V7rzvpjAu6l3iaHmRci/IH4O2mzvWJORscPfCxRRSQXi87NSrBQ9J6HeZ5XQWYNh
+FhqlkuBgp/i6XTvYVhO2t3+84E0JK499hiXxLqWkDuClm+5c+Yse4FGydNFrzGK
PIRiNvn9cq5Qn6O1VsCEiWJQnwjNqoTP5bf/bUPfRhl9WWFcv+hLNEUaQ0pmEoP/
JoiLEFB6iKFmSt0mNyNqeH1FfiMyyqLW15Qp4gJVEhVTNHyNfpyKYWpdSo58mmRF
Fg0g8VS/dx2iMYkdRqHmrHtWXQ+QBegMcns6qUu7r3TV/iMWwzLAFs8CPqV66ojt
pFU0VamyO2axYlIj4mj9f++QROL2ZkkTL49KIFhJBljuqcP7qOlXqhna0pasZdWC
OK48FjDOyVSTRC+GI0j+7/6WuXHE8PTbK2TizlJcRXpf6sRJabFjh0D4qMN+ZLuw
zGe0AC1J6/OmOLWwMdRKXgAxVI26HIsnQBS7ZdCx7ld3STu7gTIHpLse4comQ6p7
PPiGs4ICnYAdQz3Na3syMHlZwohILMedWgP1BQjwhf9L7lB8pWl0Qrm87qf2vejw
yew8TnUsmA9h9j4dFp96VQgCgAr/qoObOO8B0vVcqHYPi63SrWS8X7fkvUn35C3h
YENZU7tgUxII78IYhHFS+5itNfIuanhPV6agk9x1ZFlW66yJXkhVOhjH0yCger3+
DQ3Q2i2LzXEYzHdhNCyowYPR2PJ1N2ZKicb01a7g68eza+szZLJL4Ehxl1uLhUSi
h6kuQsmbNokhAQjFhmf/2vAuIkJoDeUQHafa8ieXGTy+wA38OwLnWsHJYXW9IUbJ
NFbv9yTVeyfPr/Q9y3kqgeKxPgJ3FLNkGe8oV/9L43CH5loEC+JvoSfyE74eUTl8
1rLA1ionfJWVFR9r3qbIjW7gMmD55MRxn6ZPf184yV9VkMeIbYpKPxdip1gZRsqb
5rvYIVR64Y78us0BptaG6Rb3VuvsBIuZQWKbQvNxEHnbiBJx/HaChRYacHVr/Duu
ksiL77gGTrPox9CX/tCmVRNyRr8KGbVo8+YTx9Da7pOGilJQHFGI+rorI9SNPgIE
iZ7Vw3dKITGJsGttcTFFEyDZez4LxqMhLr/9ST4aEEefO9bTqzfzZok/kq17TU3q
XlCpW54XhKgYV0tCiTJGZR7h8rigTh0RqwCLEzc50TjRLmgquB1IDKS4KpRt3DJy
MSWxESSDVPOxPsPSFh63u1VixtfvrUscSXhxz5SvjHZ+JzQIOWRDXT2NF3YOy+O5
xTsQMFX6wPPOuN6lrC2sf62+Gi0ctvw7C5x8DqWWnjbcjWsykclhV/JxRs8FJtDh
JK1LMprk95afX8VQONzpjICzuMaTfdL2jtuo8fZ2aIgDfAyYxU5bAcYrsDYtW5JY
BbI6xSy/UUVSaorztUcWI96nAb4JB68gRYZCMGQzuPIPwKTLlIvw2ZQ0GFE45IN5
nlov69u85S6Hzxxam2JV3Zv13RUWYBh2zQ1f3AJ1BF4LRLaxrP/Dl6FJvgapI1wY
Hj5tUl9sXDak8+AqldJIUm3y0XWPICEjSghIYsWHoYKxWurIdm+PmHEEyPakFqh0
qRqMtqwhngYv1ncfRwdDjhrJ1K5vdnol1RLQyul6becvK3FMYchswkrNkATW2IpC
7sFPRvhkOu1+OFLOz1NSSSVUzf1j8I0vsA7CrdHXTYMLNwbyB3Mvi1gmpgKreKqP
Oij+lFCu4fXZVwNex6QKwdHubNhNv+Au4rTkQiTCfhzsvBo/fjye2CPlEEnBpHuW
EBsOfoLgCOJxB1//qGTPA+9SOn1GjQARViYtJ1HUvoL0CgzCTFsACktOjrrMj5Lc
5IoJfihhhSaKoXq/Giy6cDqQji3XoXbjB+6WXoSZHJXOuMF5OJxtHo9fjQDMERyO
B7DdjPTyvTa/lfJjtFYK0kLqY1GBN/rr0oeYU6oH3wer9hpgZS8XKDuaodIY46nI
RzlHTVcuZ3bpQaVJ+zSSAsnvdDNoT60qEg8tb2cDAiEhCeTr04VUBO4fGScd3loo
u6udbWae0zvIi+mAkmcgMts93LLsEgkQvF/SBTTM4+eigDKIfvPnrdd9GlIrR5Gq
oZktXFx21XNk1z2MaZ0u5To1vCZQQ2df8ViWZD98/BixMDP4KLMCcMV2oF0To4PG
8iGFgstGV5wzvNfGNbPOO7w4am09g53n5T+jJURpwGvMp78+/z9SA0ZoQBy4canm
UzifLoJINIb5iC0WojjzCrU9WuzK1NhDGFru+Atx7F7bwi05sj3fUQjawffj8sbZ
8TNtKyY93KdnwscO2QB5+eRocYdzekWMXG37KtNju4D1KI1FSTijR4jB16xKzago
pP0cBQHx+ve9Ne9Z/75FkHYjRvn1n27G7QtRsK5XRBJ33yExIDVbZWAq2IhrC235
4FHypiO/3zugpHUkeXaQ8yOmHEAT9KtHu3V1+HSWMHcaR8jJzB+ox8EXnUJJelcu
9Fz3Az+SzeZoJ8loi99Lse0V5kEHol+LVmWYHFEuqXcmW7RXWLvvCh8Wc39fHp4I
RZegzeiHwXpa1AzSgXMZ+2/wQBzjZfIedCHapk41m2fk4nIC55T1B7p6CYDxJfjm
nQMYrnGpTN3oSXbZ14daawsYMfFkwFEptlIGDB+N5nOrsYUYmPPelxnG5ZNK+NX9
OnsBRqNoo/CP4OqMLqR451xRZFDJrXSxrdbaqWrkHuCZFY0MpHJ3UKGIKbHWRReJ
3boksQsH8CtBBq0JyCLI2h1TylZrI8WiIWqYuatfjtJv4B2VTPOanvZVEPKaq9+E
LiWjuy0+7aysfNbMSYOOqZq6cQOALzQmI7ojeMbBtQ8s5u9X7lpJMvirUBshgo4x
PTuR5MPT5C8lGWrrg5KK+iSJ/8JhS85NwOFtISAFt1l5MQRo9IBjAT03SRmKEZFV
qqRTKemWd+IroXmTil0EYJ7rgUX0cgszhXp5DMF/k2uiSJr8mk61s0y00zC1DMut
eetwPAo0O9PS9oeteT/BOpUTp9hR1RCBUQpULbTTmmNUQ7D9+9Fa8R8/ph0DrtpV
JLxORM9PrIGFoDQQh1gGiQPVezOHCD1yz0QFd0RqEm/uw4kgY4qPTpMbXhQ428Hr
Z6Fa+Tdflp0pUkB1aoI+YR++ZSVpoPULTTpwMhRBbKL8vSBXKKRG9v9PCHLtvmpw
vrPqI034L0+xAJ+tzVu/COq0FksJSQicshNYSP3iFh3nrUi2rOM7IKgqF/rZDAk5
pTL+rPw8zSovH9InWT0vvKRtLsaPmQ5G7UGOhx1/CykZYBOrKoKj9BKxNii5W+Wd
zWY+bR98MnFq5UdrvD+qYDT/xucTeG8EuaLM4vKhCBk+nwiMHQc3ZO937k30SWL/
CwHcRSbPy2gnSL6n+Sm9AnGpA+pTD+7mwavXg73bB5TaZVZOPNSUnI8u13of94Lu
Lwu7kOovKqTtS2XKjUIEMMAAKTzlY7emAI5sWhZ3XAKJB5bU4cG3fUH4bF+/PKuL
mYam6AZxZq00YQ+cX4j97MgzAo+5HbX38GZavsuz+M4KwEOwgVavJbPQ+OiL3teC
tDat5onV88Fx7SfaGkf0oRrpxIPgCNgyboSnvf5inSgDwQDWBT/Abl7cd4TEZphv
BGVfNDNugXMWK3Rp9Jd8UqyrmqiAtQjAC53sK9rOBPFQ7zVy9QzgBN/et9E+M7CV
b+nQksnGSL6JvgmNh8PIoX63hBqPhC+W2D7hKfYn/ghkPhr/u05lLOuYv1RihsUy
RxqC+wVgbsAjWVipDovBPQsjwqen+k5i9W6qDP+/hU0HeKRRcxzJSscVQ2MNtw/T
Fvj7VpEvvCdTmh/tGXs60l5yKvp0h/nGjq4L7d9VYZxUq3KzUj7CM7SYBykT8TOu
iQ6Z9b7EtNELjyVaE/DbvdP+pQZ+clHs8Tpwy5laJLKbM7XnYtgxSvgwo3ds8EMT
GjvrPnJXgY56txsiFwDqxMxnch6wHumAEcA+oyg2z/ZzdRD6l77fqHbpA0ui+BLr
cXc8gO6HLXc7AYyZQ2LGqFQV114yL+cJ17M5+aADb0EDYATfHXfyyHlUQrrGCyZJ
4mptGWN3ZEzDnJ8nrqxaJ4FQjs6/XSoJA/OxvGmP8ATrmd7vMtnauPbWIJZ4Ed1C
X/Z2OqML6yeVZIMe3aPlcju8a5vY7biUrCqvokT3hz+zdg2+BB0GazPPRAX+xYom
K/HA5zzbQf3oERwCX3so18BTCeUmOOJXNlci78H5vNLa9f+39Nu1yZVlfzAPSxlr
RoNJbSljiHyY6aHUOMsLjUH2bNbDMmEAcQTxM3CfaIpOYzH4cw41JGDSblZU0ShF
sAx3r4IjKNCpOZPzYIudMjyEXUa3IPcYAn0hdMzGqkuAhuWW2owrB3PydmXa7z9H
cGAb0gM94Mgzz3Q9bzw/8zafEhLEaunmW6sSK6QT61Bl5dxOXQm8/Tw0mXFRLEyX
q3uM1VZGWnvBNfrp+rQqJ7TJm2qSLrpAHAb1/hqQ/CbVnoRZwgLOZhel0SYLtHBm
UlbCiZxpoe/ChaL+EGUQ6XfXxjP04w7/yhTV4WoSOUSLdwq03xIQPdK0mR+n7NwE
Fi6FBUMWjhQY/ubq35zRhKtyH6YumL/3Ns5IrQ8GKgPJp1woaJGkRlNKRxP7K0fT
JnpmNy2LabNiAT3u5+IhgTENwLzl0Zsi/Lx54v1cFRvOxyKbsI4TipNSBl6zRuYK
U971NwRea743PBvZxLT/FQvOxktWglBvjX5QU8sv9F9JXpVz773fpNEPFRfq0DxM
/gFwoWV0AGK+0EYVnhQ5Jo0hHIAtScVqEkzx9qqD7Hm8Vf8Na9v/IXeegPw/q0o3
Qq5u6H3eR57FWh2bHtU5/nfo2E6WSE5YLjzRhmJnD/wn9yIkly/JqaFElEXtRWU/
WKolgUwFGTjOf9Q0AjDgh1MyLzLscPBV9SMukQpUq2nXgt/aOlN0zOxjDbJ9hjGs
cPL4U//ZZigHPpUtTgrBad7xiAKdpkgnTCywkvXMhIQLae1mCKmDpZG+mffeEMNG
6v+JqLFKagkCvXM98IgliWFhxE1GXhRYprCncdOfid8TDCo+CACUu77HcIG0WyBG
g+7/+FLs2sbXtoNTyW4ExO3Bgdi4xbSquNzzXmgc1BFGsIz052KU86iLdQuWj5mg
ebLwZAY0v4eFR4PmXpeeiyvJfElPs3lyrx1X2md2+e5AksCEKlJayB4F02TFNlC0
L/ivTmUvqLAL39htq1FPOIkRwDjQnv+PJ3zgoEPoOmryfh9pT7IwlD7gFWNOyUL4
9ZPkyT1Wd7FT3Gfsf1c0xl67spgprRGbo/js8dmh7RjGaeVuzzCE1uRK2gINN+Zh
DZBu95XDUEs01nmJzlh5dmoWy7SCGwhbJc2qEv8B2dBefMYwp5YRt1HUsw+T213r
ZEB3D12G0pLdDVDarFudNmlVpdJdEDvcv6jX/tD0Xw7Mx6BtJBuapvEbUUVJID23
sFHJ2xaAvYOt5PKnTANhRPk36AaCoOrnp8WDewSPxwkkDOsZSExX/TPdoj/LOCzq
ShQeyOPblHAUhwQF4fr/2xBUPkHU6S7LsV1C43R4r5JqD/wxbb5vTkcG71cS2gES
GIZWNaELz6TrkiPsfrJBQItk5cH+EWQ7AuqcMfX0gva0qW9JV+dShuGYWenBzjoF
SEf4LCjdkWDhl4QMtiNiqgeXq3SzUZ4wfLNg7rYpdKdbQAMJoo5NurcQZAe9bM3u
Cz/Hkz67A4oXVqUt/dFEYIpHip9oZnGfAz1c5fNWhnCyc0UNcv5/xi3BCBjETQy1
ffNXa4T9+PqJ7bfL4xKxn2xwFfl38n9X7HA3nCGtKax0xjA7wxM5+nCqYLEiyOKc
HooKIa+cYoI3NGuYdSYUveXar8iEk+AdfIk6mQruIfxZY08DBM2IpI06tJeYrnVW
SSBJAlxi09lIaRRaQnCMgir8l0c8tf/CIqz3bvXGRq1ke5EzzSZfkmF9nwqTCdet
r+QN/MbHHAFCc+5VeOPp4fjiHsbLfHzKAk8/uNt0Jmf7YC7Zg/4BpJLvLlU7Gvx1
mwbpkHnFdwxXeV3laWV1I+EtorBNcXc5r9MXbWPhVjG2fRlA4hYl8J8+IyPyxHGf
1eg8ArzjOGE9uXBTp7fa1CG5Fgcex2jacm6Qy9KXFl8Tfvwyu6v6Dax7Lu77Rf0B
n5mEn0RE64Ub+Y1rYgcbG2X/+NKzZvqSApdfUVOWHpd8pQCTfDEjDPXrI+BtVCmB
FjlZ0LpELtcLNqEtu1qDwbxv4XYYFPW62vduJOMT5kLuh66rCembzMZdHAv3nFwl
ZeH2MSBCWx01Fq7NGA8maXVMZv6XCxUK5eNlNl6t0kvWmbVV8zLavKNo2206F2gY
7FWjKAWjvvkj3ieVlNkiosH6oOJP386S7Um5099NlJb4qwfz8dPHHAbD07K5Tvzz
SMxgCbxY2melWyJec6b7UsTR2G6ROByy10+LBa9XRiV2Yk3RQabOSdsSQ01dnJk+
vAKY3dpmhR8KUcFhwbMY3/6HzOtBHULprO06tGlBRNpnA9d7VmSCa1j3lVyryTLr
QDkkl3hjNoLjOXCBO8R8U4aM59vgiUaHFfHm7sOfBeOOS4gqhe8MstQuYasS4lXN
QBgxbKihtseb9/ovfgaHFRd3LLAOkESG0Ql/cIX4PGYRmBHidaMCVMlT0Ydu7871
TCpj9697OH47TVQ75tPKStQUb0qwTLxD16qC+9hOU9Kp+7dlk9dKUUtU71l0GFYo
o15UFb205OprnKv9xsnrGp8v+l9wnb61Z6zOadmqxQBTKEqYY0WwAM+QKJSo2TbF
0s9UkJSZqKuazulZNM5sKigVdMfx/GR0sDImgP0MZOuDiqrJibDNaF4y7u2yFntB
Pl+P1w6fBo+6uJqZzF7dFDJSuUPRK4GYETAeyyWLaMlP79GedHDt6MgQIx0BDufs
P3qv4aavqB+9uNECsgw6mv8IyAqWk/cGVQ3J+Ehx5sEOJtvjpK74t6kQudJCxPpE
Vhd9VjqcggxDhLT4hcbhYAnzjm06q1I/e2rdpszfL+DKL+dFfv21RdgNMxwsbQ0Y
grufyb5Z2ySnN8atbqMcEaX4HA70dVN5QC6TcWx5rAqMzg09Et39kE+IgAPvPVEL
s9zBSbABhGOVyX1+W3K1M9SbONPei8j+bCUL3Xt+IXbOwGxh/NkVLdpjvOF909HD
Av/JNE4TYIidA8tE866d3T/kIoF5XLSFm6Nani2sG2oovy7rWGI4joXw1I13EyfS
ca2+61CH7+ttBm4hnrzsH0OfaJRORGVFA5IcmhjATjQeeb1q6AdXw0GrfgdmVlVS
J5WM1Ei0HACtneJBOQuUxUacn9ViLD6z6oBGxUxmcaJSjp7HfO700UY1yWezJAEA
KK5qNrYD0cJIjg/Fap0qVVlLdulkyK27lpDqehMNWqSJR/YL8v8zS7lEk6OlQfEe
bE6iokJDIWZX9Qsd0BpFmCkuJYrDFK93o9LlxZxpoH9f2EEIxvziNjNUS/MaOZ/M
YyJelLAYRsS6hvHh3ijoutFoqvjTQWWj2d+cB5wc9MpN9Rw/jeVcacWu1jCF32hw
oSGf8OoMcDXK37EtOzWq1t+7tosNKv+7ZoxUElYvbiFNXUcQleGSfnqA3bfIVRdM
gInctJiX9s3VnLDFFiz8sXqcE/r4V7EuRifvapMx326FmQWHAU8UZv1hlMIc+qjG
ck5Ij0/QOeSscq2S4u4EBb+1xCkOnX2zRBjIxbSx5LrbOxFz+CF6W06CPTly3Zct
ksfeM1toLXRiDPMI05OWGD1v3/nxRU7e3Kt+mkvZ6AiBr05y4a5A0rOphct5eAnD
Y4GNsJP4TYqVlq79B1w1PA99z29qGfuBOWZ/x2BoCDqIam4w10JRuGUFC+1a9Tot
DFl128NsiN427uiM78Q+NDQTJGrkDQ9mROUhOFy4T1cRM4HDi6iJoVsVXI4PQGYm
iB0tEzmue8TdxUkmaVJuu+mqI9ectSI46W+5/HTuhmOF3ztoKNUdctyePkrMt5H7
iRbJen68uBAoXSHLiSViiA3LXqPzF0eUWHeNzRLTHHuaa1LBCHVIl/QAd8oyG8oL
Fmag6Z9KYCwAUNAbq4RgztUpv9uUYbM6D1UR/e8QGwD8yvZRMmRHaURochPiTn1B
kou5Hhld2EuLMpTNmDtgp2XEMji7PiIfhx5tzUeWJwaN9AmRDPdI7nC6XOxOsv2x
W8huxOypiMBHOkTZqRp/nr+oI7eQEXbJ3ZfqUKxblONLc8kom+1OagtC90weQPnw
1kXc2FBJrSRfXxh2aj986xfbvlHTrTj/3WXsnVoFtRI5thhyR1x5btd1A7mx7ZR0
XHcTimviMim9y7t6MSo8MjqeVo+QBFw7r7BrPr9XQU36n41iKhQpDUDnSEAdASLt
I3Sl35Gx0O+uPTUn6YZ78HiXzTm0L9dxmC6E5CUu6yKIDnn8sGY4ipPywEQ2Lah3
9+T+6InpqK0aa+Yq8GkiN+C8+LTU8nFq9YpaeRk+QECo8Ca3fvSEDOlh/nWVkyrf
CwD0zAsPc1cUQgAWHqJ/QEEHWzeakRCbLD+/fCY1AQP9ijqOZRPQG4AbvGK/mUp2
wVbScxspUkafz/dvKKv2W/V6ph1H2UfmC4aM75IqVRFJZ1Ilf+aZhfz5ZZnRQHmr
IexNCZR1EOFeGisEXAIQnAKFL9fm9rRCqJUijhULSShe3ll7UBUZylK8WJuJQ+s8
+jtOpIcFHUg7XhboDYt3seRwyl+cGlDR0BmCwgKDX5ctbRW64ZRgN4jbxJKKNrzv
alcZnXGeFhBRtlAKpUzVwHQs7KvATTMXcrO03IrhXkWKFuUbs1ld/OnPiKBLWM8k
59YEJv7Rh6x2SK0yPr0nwexbnP704zowyEuHSa28tbuCxiLANUF2EmnBUdmckGg4
PJaJztqjOnEgr/kqU+vqqSvEmZPp0LL6yIczD62kTgYi/IcfA7h3093W7Kf09zOy
ilBEx8gsD6aW6oV0B8jJiwWO9jlWTj3GsofX+lTRd6DKikO9UBfgwvc/xDGgVZ4O
cwkMoj3eK8LWGfHu9Z2nAWJakSUWulAP6IkwSxVbEjkAmedEiSzTge7atV+RcN6i
fw1JgL5hcIGJ+7AUbDr3mecONh6mw2aBgqUO1nvAy2zampqoTkoSGWzxy1ua9LPj
0XBD49357n3eIOXuxjIo6/rLoWUnkoSv5+X1laZmVctopA66rI6ri1nylgSH0COv
PndIhLOQAoDAv0vkxbYKhKh4VJdZWgNuQHZ83sVPJ1YlhpmrCiAsEJyESLg6NlcR
VITYBXzjl7Xnwq9IL8RJlYV6BhMf/0VaNMS3YNizMuBxCmcOFpmd8sIs2mJCVZtK
LfGip4TH3Op6rZYBhkNhc4trEK6JaR9QYCl9NdA60ACrGknJJqE/LXi8bSPzsEc8
O4XaaeiZLeHiMsyCjEkvLKwZeQrtCfcALIU8TNC+vSB6Pxhc+pRj6AIIkRRcb1Nz
eRf+YkzzXs0BhcFk282Uuqls6QAgjjsIyAXxXwwfEyFY+QQwVdaZ6s1rAr2Xy2oC
MdwXPcx83Qk+9l77D7d5BWbWqrMPIQJlnrDidAHh2KSkNl7/p4JlU8OM6FguZIdR
q4ZX0JyNYw3YD4NDohjvuKh24iapgKcAqLtrfuJvc/gjflrDpjnzEKrOa1Dyu+8P
8yB7adf/RfpL0P2qTga0HSbGeaYDr3UW9Qp5ddeUCKocQndgB6PrlK5UyaKqDmit
Fp7YNEBjMR1Z0P8ggj98exkrYqo2fTcY6N9Oux2onznEwuRcNrQu3Xyx6ocuZ9oc
CeRMdVE7RJx7uyMOBv/kGXWRrB/+y2UZc3xDSj8i+ski8cu8Vt9Bsq8ATW3IJInx
5xmdKrTwCf0wXqJZqon92HqKsVwjXdhqMM6XFwmX0Wz/Lj6aGR4jzhfP4EgwLbzJ
P3RlFDL/HvYcprdZHkxLGM8wvqFp8FCrrQhkRdw0zNRZ8h1j0IvPFn8lwJbXWNpY
Zuwmy8PbN26N3ca9BEt4dSIgdH2GX+KSBvqV+fVTE+Epc5rf1S7F9L817kpVvp1M
9s32ZiKjRmBO4vq3VbNYUEIS9WzQwTS2u5+nw07KrlFEmGhQkcEWykQM1HH4spK6
mJmadHprARDTgGZkWWCtgd5sY6jZLPbSaXhxepO3M6n0BFnMVZqXArIMQuPEh+lh
uZqmt8paPnWcXS6cfM1Kpjg/5HoeetJwNO0kZqQ2R49kv8hXtvxChBfEavF6jiFn
8QDRJLOCeQ4+qnX3ZR8VsDSrHR1rPxXUyfCvhEQTqVhzzESEktnaNlYQMg18Thhp
T61j/e0cfh0Lplbz+B1B7Brpcq8fyqSgOB35fslSJ5iX0Q+jKcp61qGF7F7fs/zo
c3k/rY3kAeu9/IG0Eu5fyj26HmDLVkpiYu7JbiL1zmHyWqIJRbHblqccCqoY8EpR
vkmCp2N7NSK9hCEPgsKNgQyy6s1p30mHPipd3PUSLjMvhY9ySPs84ojx8YUxKxmZ
d2J1iEGYswhL+8lJ6LUkPB4E5EaGmpAmxthiSfINWtbF+ntDozIjNWDTyvidOlhy
14fGC0fEeJkncPefwVD6yeklIZ6Hrlea4Acl23n37z4OTA2M2IQfk3VWnXMunnxy
b5VpbBR4AUoE5kKZl/pA9sXoEi1w45dKE/nfgVy0g+EzViWBw4/KWtkpMZNedU9T
W6U6oMyHHN5QHl0AH5GUvCTu8AnMaWasB61tFg8HOd0adKLQhVUaywgrZ9RcufRo
GKDkFsDxHxAAHIXx2zMy10udzjDpeGsGlUOB/KlVaZoNA2oRELUZniB1Hu1N55nF
bLgrWjEqKvop0U54aVKMuP7AAKX2EYmUxHvo8mGwb8+EXhbZNnEEeHLZFSeyx/Hu
`pragma protect end_protected
