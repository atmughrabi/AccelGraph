// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ER67+FbfaTuwx2QRF9QFK1GxScMeu5diP2e1KgFXTsUkGmw2lwPodFSHoPpwlhyK
JG8xTTcsXjFHapx6suUtqN8p9QzqEGSaiWe/1u36Mn+dYm3Zym3j/c5nikShqalW
7chQ91emRPl9ZazBav3dUhQkg/8DhnVFrXzySTDk9N0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28016)
SkEqaxhhh47kJ9ctnVJFhgQrpfmMVvsBKzqgm7dWQQpshaPcX4Dd7VWlW8fO/E6j
KyxQ0SPepS9ayRTYh7sDMkT/tchjgh5y0bqvtw0XhrmK963qQESb4rRbz3r106+U
0EkQDjNgMcM2gszS399+ptQIgqFtbB1CANARJZmFdCl4k27fZPe1UGqkPKiOiXFE
wOraxmk+vnqs18uuRzdc51CuGFBmqNvsvP7e8PNxyinMMcOLNdhOVbOk2TFVXdmZ
NkDqxq1B2iY33bL91Pd7grZYUrITH8oir+r5fFg8Av5ZhBV0tz1xo7TpxW54HIxD
SHCnHi9jZ6N+sFmKclijYBE7vTmpleMD4uXz4QS05QaqnCiGCh0hz85gPXToIWkS
aYys2FF+0bP8XCDBYquBOSASKQOgsbk/4IriWFeTvpqC3ghnJiZ4eBH07PdppW1P
o8bfSNcEeCKnyeBF77f2GPL703K3bukE6TAXIjiyqxDHw/1v3id8OeHq4+FDHYbK
X7MfqAPSvSGS5DhS5U2EFRwECEMdufCN3ExX/zKmbWbVONxPMY0PzepaIsGaPomc
NtWI8wn4ECKljFVTHzMdgIotFDSq7SxCroBVmpBD+lJcFiPC1TEd9+oFslh1h8GP
qbxVJM0dfBc/FppGrYAuFNhlaH5iBHWpL5p3x1fTFohNLVM6WFXjpJBjYnN0mdCA
JOXFQaIvxunA0BCFmSGNJOf2erXY5AZejIBPukeHH6ua2bT9Pxle01yg9IZFKQPI
QqJDuftRSfAOM7TTaRvsgFh7vv/gJJgGT5dgdg90p7ZimjKFlP7V0E3HdsHjS5Yc
+FqUP1Jx/0E6f7HiUAvblGsQmkK7GHTmuFu178EoNbTP22lTMrBB0oKc9ZPS/psg
tMhIA+F0fmCtrqNxxDQ3XBAIKYFHMDMLilhf+TpY/8Fpxf0g0QZZzW0zNoEHfvOO
6/DFoEuuzVZF5OVPRwOSefezBfhYOZQCcZz+P4oYPlfeg+J1pqh+7oDDw9V+mpLz
jxqCOQvfsjkb/K+VoO2m9eDznuU069kcCX92uU48dYtpCVryl2QEhxivkrwHsK1T
J6Lj/enQJtMT6V7LuH9hVrgyUPJz71IAuSBc6cOa7p/a27oGJEp3MtVjzPqKO9S/
wldSgFJa/AoEIJtnYlLiAqg95NbrGc+40XysQqmDnVf/cfBxpJGmSRMaQa/C0Kjx
ZhP8ZPcVSY4+1voSOiIJOgirSS4ttwTKbXQr2zk4o+X4xuXRMrJavBld0KSFDYWw
pfpLA6vYV2eQtQzJnZaTjUEHeGcj3JeNJkAddBGpk/ykLdHNwFD5lTkFjdHRGkux
p+CuCIylaxSGEeZC5JKUCcVLuKhVwtcjRO7IM7B51e5zalqIqDEqrgrxNrSvutLB
Fp1j4Iwr+nYJiO3Uqjk15jt0zDyaW9z0ikuRbrmw7NsmTjBvCZEPtsZYRkOpoj9J
i8j/0xeqUNP52HeeCFoPq/SeVf0acc291StdLYnT40vB3rJ3OonHn8nsaWymNEP1
ahREJflNCL2O4sX+Y81RWDtx6ExEJ4J25cKX0fgmqDPq3kxJ8j9J5LWBINNqfXJB
l6+bb8+Juy2Wt8NF4Ooegz3v51BaAPcjeS4HoMcEh8AstCiwhXwg+moA+VFyy7su
edDdSF3UGX4W1TajVgv8fSj4LMys+VOMDb15+rExDbXERihLXltbVkdF0AhMB7dO
xi8pXk7bYFMK287x8BQ9dAMAaqeag4hghY35XDcnkePIweBCcrZ2sRWVwIK8jDiI
vpBL90wMYhk3CW5PYE8gU2fdqlIInHJSyNj2/LW2P4TBOlDhRATbQeQc3ptp5JVk
S1FiwOgLMMYxU9flsQegdNVnXmHt40eB6OhJb9Vj3VDk+VcGhWu3oZ3qoFKyEEUH
6ekVJMWBkLIBFQKVFIhdX1LWUjXcjMz44VhGEqpxetkPK/gye9iCDafQD9qxPOC5
oTMB2KbqvT0GoLcbdKI0E+W0fAnPEsBST9CykQQupaDFTxipeVyczPUoRnrhLlQ+
SGhov6K1zQgka85C8pox4CPj1myj/v5RaGgKVHq/CZzIkENbRgxZgm5epj8bEa/d
vMlQgqQBS9TDpFbmHDrE5LoPUtYpG1pj5HvpVT2m+hItpX7vY/JfpiCa02OUS/OP
nyKZpf57Pytk8pdpp7RXFIgdFlH5+9pDZDyU9g/37tNSC6pbywznR6W820yI1OP1
RI2EGyaxAUGp65An1fl7FsBZsN4CDgiIMMv9WvRO/hXbFaB9Wea4vzSOWhUjqZiE
75Q15dS5FT6Ld/xjLlHuzlyGDeRe6c5CXrcoViAYR/9svs2QYQ2JfWVJ32GoxpD1
uNKFQK2MsFE/WJETh37jujRoXfjptVNReEU/u/WW/eekgp6L+I6z96bTXbW0ezcl
n2nMDQB3uDKH9ah50CJn88HLQ4yaPSA5mezc/s684SapOU5s1689Jr17cZ0ysBsG
DFcaFLuF8zYpEHmwc2sG316fjWdv3t1SQ9mXYFN+j70Y9erhwxVlpYdjQqB6e5oR
kzkYNse5DwhJXvgsgpJWuOxDix5EG2ttg1rlO1+kFf9n7OqH0X8kc09Tvaf1afLH
fB5gUUT2a8IofJ3U8eDBepbF9f2NsVERZJpQcuumWbHra6A7WEeqUcRErYQnnWaN
Szj0vqkk29c9o2RIUwV/hw3oh23cG/0UwUOGfEiDlnUv6ZI+8Sgl9NgdjSlx3aFD
L1IkSvSlycbyqs9THnoifIyQMHcIAC0tOq76cR/Vks7fPXRHQgzRZ9cJm9ogAE48
pkULTBJcesGzTt2Mk+DfChnejS9UpwtOHg1P04RUeTN+7ti1YCf9UyPVCkqfOJWD
GDzYnosCSy3KmEiw93T9XOKiqozIvLk/5dS79Hg+xBwiZ3XpCGqsG6lbsRgfwEi0
BxVfEpOsbzMvF0hDf1Z9e2ZsiGl8pDuR6qimjfNhRR5v8DKM2nULgKHunJowgf84
FMfXf6tfvFhip5AMegeD+jfqG2BlyVr+Hx7wf+V3Q4h/2nvluv9xmUAVh+BU0Hqe
30TljBf2+RI0uT9BEC055qSAIEnmsbO+G1OxY+bSMLu0h3S1FPZw2dzwVSMcbSAE
fYToV0CBbVHN3tIei1MW4Cr1OndXiskrbxUO5lG03HwJp4IxYR6zgJ7YwIEOwJR6
rVo24megblH7rlngOsVn0R9svRPEzhBibBvmNdYE/dUc+7SuXmT/q+k4uIykgyKO
e0ezuYCnXugvOClzmtaJo/ztEaYJ3LHmw3oRnonvH/DtvfzCExSX3z1tLSARa6UH
luVAe5WCoEdtuY2OGJitHfnRouQiU+feWUDdn7H1LAboHv9Q2uj6qEoWLgRuI/2s
Zx9jRWVOYW2uZeakw8RZUAUVScdYDyVxxecU5IVbfRA3KF3qbsZazhIB5cE7HzOp
gRt4mbvP/5cAmhGwUI3GsysMJp82WX+Ac8MWoPEehdlpRv+3hVJdnDggtdnZswNu
Bx4ZoUOcfzVnCJlXQtfdmmvMgXQeyn3SiChRhnIAOAuSPVoj4mhhnGXRtHnHdNVf
NlSbTLmLeCSGtryZxqIltUGL9l76uTLP3dGWRrtnYtTqpdC46kSWzjuO8/Xdlu1p
a3Ysma2XIngOTTu/11b4Zvn6dtEJAPqDqN2/DugTUHbyEJhKoJ6/kxa4WKvfA7F7
qx0//IvEhXT3TKvIgGA6FCuayz89WW8HyQc0YxM0i8UgHV03uQ4Pm1AsjiRK+ehA
71SJY9isSqowRsUiltJvdKUkhIEiT0RJ2u93lFV8+SljmEizd/r996h6nhd1fQm8
zghqA5nLk3ngdhjqe+9WdHeNUZEVcYITtgqSJW5uwar8VhglmXjfzQQ7FInZpJDL
w5z1CCjZvPuL/d+E0OBRVuaNROkzz/SRnekIPIj/zRXN0Z3cSZzgtCINDmtjZtHK
NoLtgRXNpVgU0n3lu169gv9pinbLmcC5DOCnH3isHoFd4dGIi2cHkMer44dJL1j6
za7w2zvHrkLhDglikTBjk9t1NAepLzMahbHUs1QpBgfeOYgONk3p6dCTrFaqIlou
KKgifahYCxGMX9f/fd5mK0v4g4Ox/5//QmB8idWFjuyQNZsj0m14YXH4kQQplrXu
AzUS1YRChxr1tjN/oY3J4v4x2iGF7IoL2vKZ7dzdY6Gs9F6y2CNUJIoqg2VWjwOs
bjV3QxQ/GjsfPlwr/Ik55nHSC1QeixxEcR3SbxKuVG4R4I07QLVzvcVoU8YsT1z/
MBxawo6t++nNxmOWpytt+l1B2gN0Fcy35vOvy1ZS+omjFazttK2uKoz4ptptLrYh
gnacJ42FFf4J/ExVPO/aYQbzEIswz2H4te7xgfN1WSY3pmeod4ePJXKKKwSuvCuO
lmUEQFY2DeB/ICd4ORsqa+0kBPqfup4nH7bBC2WxfETUD5DPrVUcYjM4eVVBS6Xk
qafqfef02mHqbs+diYFKZVO4u/5/OlZ4eFV/AJymuWOqIqNU42HuVIPt9V6KskGT
IqnjGxV90HD/U0MzMKbpm1vRxe4B5MB6DazH/5U7axT5AHiMoQ9l6OYdqt4IuTIk
tfL+KfS+fhG4TnQaA3ZozboMdyQB+nLRNYEyTC0vDyJ/PdRQEMn8uVFQUUr5D7bI
gN+MVk/uG3tTfIqHlAnBon3BiNTr0zPqI5eJRlPJ3rluPPmlrWKsXgRvVWN/Im1w
z1WJFPJJEcFRn3fpGt10yYghvis5LcUhxeAjzM3tHuGYY380NpDtTQOBMc1P+Jgj
nRMJ2eOs+WnLicQNbLi1EuV9MYTteCsAAtGrFV5rMX3FUei+2otWTG7G10kGJFuG
WG4FiVOnACI/m51cMSpXr2f820K0230jd2lGuknmk7oFrU2J/m+lvYJvVszCYVGk
cJhjrbs/DnDcns9U1AjLf5hXIFt9iFftmQGUMm3i62taCucR5auFeIR+YiND1GbL
8Vx+Ie/JGWL0m8FTKSQO4irgBFDZpyVkxA4MIm8UhQq9t0Rhi/OfoRkfGPphoT0e
EvY4nbtQxMBO8PBpjftuK2W9ppXEUaH2PbQmhTEpv47eci1wBGUhh9yzMl4mE+jK
42t0QZJSws3RRaEvwCpYKVqK49Bp7lCA1jtU/9oIqBzPVaZ7VTHBtQKCRdPTiSkF
uqAfa5EZ0hPd6ZXkxd8BSzAp0RKPSsNe5L5JXOzj12o/ApzoBzeyb01de+1CJPFG
mS6uQk0MB6vLH9QEondE7iaZwlk4lJTgnHfkLWY2RL4I7GEaX6yaAFs7VRPiusLZ
OxXQzk+kroJVydNge6E049ihnMCUnwt4qwrFxG3b7abgtGHHtmoK3NiBQJCruOYm
mmGGC2+K7hzTpuQ3669XOiGXjz/2Hxyp23K51uwzA38Jwnge/IBKnYtSdJPNiVQ1
1EyNQgBC3xTvqgUaj0ta/phm4eh7sN+Q94dVx/6a4TXRHp9mw/UBej8v81YGpbSp
aGbypZqsSxjTEcC4uIUkdeB+oTOIrKnHJxiqdTfO3yNXJL/cc8MGxU2Q7cA/djDU
l5abyptJrJTW1z31z3xfzB5KEkkGcqSGCUeLb2i60HyMzk4g8JSKxdXLRwQrpHkT
7pJAkrhydrjkjvYf+TKB6Ptwws5/Twsu3OQmD3+3XgJnjtMTjasOOOUvBZZ7rHMZ
wfsmCoZtczY+ia7MZ8/6P3Q2rfc/Essae8m+n6uGLmWvr5UgW9RZERMUpNoz6NS3
RMxfdK5fyAGdBYv2xQMqQrC83wvvfywVPZCDFPdP7rMaeghaShqIqMDF47b3+Tqt
bpRuRuKI1GkOxHBisT0p4roZwLCPxMSz2OaIlY5ZrTKxlSWdv4ukPWA6/TxX8ZiD
hIf66i63lvrdoyJkYhTwxOA70IZ2p33LODWQ4lqBL718qROYrryqTCl/NHhVZEd/
q923DoWMJDDzUCb6miZFSq1dMdEIXPD7krZHQLVewYrFiWYPJ1yMwucATcns6BNG
85juEoKuHCoJ38gINGJKWsYrc9NZgGSRn9rN6k/S2TI4mXHACp+P0UXXUue0iYNv
oOGAQ0rF7DLVGroNITIsOemJFIvdHmC5F3VnswyVKeYWlRX1tHIRY/cX0mtaF2K9
SpWvJ3ps98I2b6vneIdKXAQbtW2YIrX9sSCzAnK+S/o+iPSdKoA2x4hJWrdioqCw
P92jQD7W2+7RVTusKsWU38vUjs6gEDepOyPsM5hqGRfxVM7ZjxXuDp0575POvwh9
zKyJnhckd6dALP4+68KoHTKq4NmYDKiaWUegCVCE/ir0SAXq2y/+2L9FTHWTxSNE
s6RgO2+8XxitbATUdxSVSEE0wDCx5/3Wz2wir8BgPRMnVMLxW3ZqhPx/+izjpn6+
PdWg+F0nEFTf+e7/4WftaxoSzXz/pDPQAbvgrYL0GoD/7uJ7ys+KOdLve5AhrRJg
6a9Wx45Ur/8vQKjrGxxUThx7vTZLz5kdJ7IVTWS58gBb9h+KlwxZfiMNZzTbV4Fr
puHhIQzmkoNi7J0ODUVjCCM6GfUtsc/ND9wz+rkgCL+lVB6LctZyRSr3juPbHZeq
A7V4wH2wG/0xybcGZMxp6PKFHyP15XoTvAz9FhLJPAZzcoPUGCbBogxIf0rrSgsH
MkAq9RRfx8DFaCaJ99L/9HWJPBCpCj4DENVISFY4dchPkJyOmIT168x4ah5OQ8Iz
Pedh4rRMICO77Sno3D9P/LEihB1P7kerD5SUL/pPj4T8pZBT2o3NiK4cISulWTp1
A0sSRU+Xu5nXPk6a+sRtMEdE0HkeTrHuuwztpIV80mLiPwDjWAL+ns5fISzwhqdg
YC4qKyaC0zAxHk8HbY3DEbtvTXJmUMaXHfgP0JQko0nUMLDYAq7++SyjGL7QgSbj
jUo8L4gLpZbpnWKvCOSeySh7McqKGAUVB3l3K3hq2Zsywo1qClMhZiL0o1p4lci/
buOqISMw6kdSUZLQXeWdlA0l816AdOCEN5G1IXvm01R7K4NEiqFDaBAn0UAi0y4y
zLITDrcilAVyth9lLUXd+I5NP4wBZybXkIOsqZr7tQ53byKSD5WnINtu7Pz+nktX
RPvM70Xdv7Tp/KbGaT7mMEKJ7JXnaZ8XDjjUuCvqT2g7lDqexLFPeI9JMzztfC+C
tHZIfgttE8B57DdHS9SKQNWbtHjsuV3yb5VeNcrWmvbeXHT2qego0aiDa8g979wO
ZXuTgu5MDjBa1fBRoyDHYN8VSr0bfZ3voR3o2RKe93XnPDpAf88JRWE5JtLWE/Rq
3f5UmNRds7jTEQzo0lVxxIxIpW+IrOkMjU6AZ3jdHBVlKeHF5aggAeKOEO3gOFcn
aLiF/zU/rg0NRhLPlgOhAdLX3IV4zmOjwnm6V6EZEulM+deYR4hVGCPeH6Qk2zTC
YumnSX2IopGxmAQ0ULYo+j6KiOK/dZQSApZBF3+KQsF5oP/5uXPGMvsIpRU0qMKT
t41bqPPe0juuIo7K8JyVTO9dkE5LC7aWz7QOFR4/tKHyjHfCe5Vi0RJe+FxTtClG
moHf9vj5OgccuNot+6qsSLvtpzAwURaJ5TCti0ge/KBXtRxx1SnR5MhoNjtGKPMu
kTj4WdmkiHRDjAII9ro8LZipmT8Ig5UOfPgPZ8Nba+iRuJSV5slfwh1BLMAZqiWd
+O2F7+k5o9U8qgKLmnp0Ebjp5UfyLEScjBhNKdWkA3ZwcoHtuZRrItXm8zYkl3j6
9Y656VBT3z69nCsvOiQDwQdFIfx+m9FNIbioduvoH+OcvdYR1yTN23PKXBxBSSnO
oJXA/M0q7+dZKzQ7NXNouwOl1WBB9zVol1OSX1rLUad+NlT0Ln0s1XXjqkxoPwAK
NF6DqY6iivhVmgR+3eYiDqGxYp2yA9TDmJC2mfUi9wxzY8BolsYuN1beufgDsOze
PwUMV6aEOHIK6jX21WviNrs6MF749G+xzKgE2NghvdPMyEyjzq5bKYk01gNxrdwo
qaqPd1+8O5etYgWX1vQKkwdfcMLA0ZRBk/ffcyp/BkA8Dc+iSIe/z3OYLqCUdsfB
ibn2oonrkRFvt9F1GBqKEgBP11GavFdgYNehTRG1mHtiKyXvcI3UOq5FkyjL9HqR
n47pjEX4MwjfghR/wbSxgtn3pPK1QVtC9Lq+3uyUT7cw+4Gr4qWyOKFpmGN42zFI
Rk+2Xgbx/fAd1wiRkRPO5boJ3xJkqwUSAPeCrXBceyz3zsdpbMoj4bHBlMlJFoyA
+WUiQw4O2dbyrmDU+l+VLLd3qq3y0EXEDwG29kbq1VlAJZEWZ6TMiEcIigLn7UIf
8P/qE/EHvuvzYYksWnUwp3QWB898veuwCQm7Y6SA5bHHiuct+CYPtQxKY/mAhYk1
o8fQ8xHXkouBjBAsk/QEw88G6ojOFMMPo+SVxnaIv7om2LabmWy+1TJCxM1TH98q
ix9IXijMe9OJxw/qJhBAIzmadzB4/8Vb6nYkic15/piOku9VL/p5l3UU8pzlU0I9
5kXW/kB2V6qfr05dXYTnk0GHMUC4iBc//IzQAA9dGg8SYS+Ynvjk+9UVCL2f1r/b
cFuUYeA04QA8rLhrItvnrVgTAqM2wDbNtsobJBPstPh0xK8NoYlwri+1WPretKRi
f7GE3Genj7Yf5kSakhj1nqFn6RDiaeBzTC3Mk8RGthCwe/H3uxfa+RessSyJwGY7
Jh91S8Kt3onVpyKERG5YnCnGfNxhLXbywe5SkMQestE8t0pAPQiQ8ngLtCrJtvMQ
/TQatnEySQs1w+QOYglceLxlKUjOuZsfJu5bhtwwYVTBPpnhxLguZyF9G1PnByN8
Fl44pYpf0qvGzi1ZwUORLt5Rk4Im1VfklLedMusIlQqzn8HkOzrahMdz+A/ryj2Z
DXHFuRcTlNVPRXumNJnMCKctgeViGHMAWeuOkgQNKzCrqDTyYSlq7HTVR9k5pE1f
dukkQ+vV64NHZbZ9WbZkw/BqYv+wdR/hmULS9LQ/gAM5oZ3Q/Nsn6VWKN/JMMmPE
N8chypz1XXeVzloEKbq/PU0vuH7eCZ3Z2wxDarRzP6CgJxzew16eTom+RiI6rALv
lcC/sz8jMxgoQ1qgxpPTlPu87HZxuQvkAgc1uDqoeuqU4h1kz83fZMul4HBtXli8
Aicod0KCV3v+TOqPeXL5toWwlZVw115SiPiv1vN1dtAx1gWxu0RtzMNMmu1F6II8
Mz9hukyksGhUFtQe6/LXX/l/9uT7uiPV3mSQKA/tv8z2k1SwBTPacA4UPQy7Nxoz
EEDKpwD+fIeo6R7Cci2IIScBNUtXL/btg/G46oFWQ4rIVzhv615u3eYG9l3m1YTu
xqzy2NQJrcjKIROUrz5DOdGtEbekxXMXmmljtkde5ZlyNCOAoA8b3v6gYK0Rv6FC
IwZF+URAnKN/pAsbPa97ByGuwWq8PSDHMWlrTWFwWSXOHdUitZxPBqDY7juNbnDF
e/bky8Pdtsdrn0OJxcMVqpNGSoO9SC8MvJp9t90pG27kC8bb4Nn7ojJ7882Vv5S0
cm9+ui8hOMOFXOXTBAaRXm2Z2ThffufboxiIKIl+fn0BFyRoD3GDA2VYd2zVLSMZ
2Ed3BAggrLH+6lj+HoJjHA6GAjyECzDSYCUV9F/Md9iS0rPutIZCbntIPiXwu33q
MGbzPnB8Xa0r5KHPEbTDXBcUytXDwPVFQ3C6xuq112XNSEtjPhhWzFbM+YWrs/vK
dENWJoRO7kFPOHepML5kO60M5AGgWYpR5NQomUqw7BvuXxfmEzFWX0qStOVCOT0D
mG6nkwLMztCmLimV7mSRTzWOAdW/wMhIR3Y0jM96TK+Ydkl6QAdlAomRlrvtffh1
58DQ7PJapzQPnhO3ZzO3r9HN+LVAGFVtBXAnh0vLyBrcw33Iq+PxhpwPVfkPa1f8
B1bNwT7B7IBQTSEC/G44n/SX+z4Yczzmkvu75Um7KXWR2GOGNlcsvdkWCIFFE8rR
PdyLljGhvAZ9BPuKM8iYPCzpO7INfJHx1Un1c//ATVztQjFZIRNfag9yrT+ys4Ur
csbA0OMLOsULUDwzYYtjNX/Gpql7tWdjxgo0xcS4eCFWd6RokDCrYTxxSLAjjAWt
am9EQtqg4S0juBqcQf9fwl3aNUbW6FErXqj+B4Ipit/nldlJpYfqil3CEwlyqUkY
t1kw9A6QtnWyMbDa8GQo4BoZtibAaFc9GDJeA0gxw6xPB92jS+MJ10zdLmecUs2M
CDDVO5YAb+BSrB/sFC7IuomOuGnqIaeebcztbCPdteV6oT4oDCko3+ldu6FVfmVs
hg3q4dDVxusvX0bjB7ZuFnnFrtdldkS7jV/otjR305QuGneIa66qC5zviybWF6uX
CwzKwJ3mlPI0WYiVxjwNOZKxGO7TCHQ7WM6ZWsgs3i+jew3MtfmXxQPSeuIknhau
++Do9qU7NmkYLGF8AcqFs/xFqcYmZchkI/TGJMuveavBq59rSb9bPOx2/DOBSof2
7avY9ebtAaO0o3nMchknIutxC2fNYcx+I2k63bLYFdEeAK8VBOBUoPPymDtVlaHZ
UPic93JGvbXeTvFtvow3qaMql0f+Eg4bfPqguvHs/98AE7QiF9KtpbPWCNhgCqWd
A9H7bmAntD8vxq6p1J0jcwq8fO1nE4WFlYtLbIMiAog32wyoHu+hp6lZjEAq/fkJ
+48wcx28QZ3P2agwJVo365iRJKE7FaScD4CWyXJ/JbqusWElgaRVNLtAMo+5CIe9
KYHJPDDFRJJe6K4h70fxk82fq1Nr47tDpe6Di+auhIYmf4Rs3NvT/wM0kA0fYnN+
e/WCjzRRFgsMuaVxJKKP+fqf1O/+BxWfwCnFrzqWOjMgo0vELOON2dP59l1x8qOI
y+LN26imxLJxbAaZzSMpNouuxzUtL1+qk0wo1hiWszCanOSvX/8sjPn+4CNvMDVG
HC/EMwLf9uqgFBozbGPvLVX3sj8stOvGzgzn8MPTzSPEGnfsAppNHwwRipljLNlz
u/fMwnTsxW5e/FrPbvZT/M6FkrnDDrHrQ7bi7O1uDX6D+EygK+itO4y+gg21LEjN
KbxrL8ul3ygtXDi9cP6/hiXQdEp+TIIGWkRw2i3WGoXBvVbCdGQf15Jp4+z3Vqa6
2m8UfZmdDdmY3djDGiXi4e8gdhr3DQA85mtQb+HkqV9ahMfCoSv7n8qyOPHUX6Xd
9w4rCLQezcBlrE5Q6MTiFVeThYeItyrbJGPb8o4LSubqDolQlFdQUuvumz1DmNq/
D5pSg3QtIrfmylq2y93BJjdD8acKtnje5Xg3x/gMOufr/YQMmXC+lnsQ6jeJHGoi
KrAnG1FL2u5ewSV5KEOQsOxcWSihvxg8KdYe08+g6/JBuChSqArs96jEDzjCWRWb
Apdg5hm6rGGHm6ZIp3lYvWgZQppc7L6HzQJ5jyaMncS73MFR1+rtaO9+wTFQ4EDu
kdGWxs+o4bm+W8Brpr8RgMUhhE4743rTun8wVlPCZeyG1ROiGmU8Hy009O9mDYE6
xTryLwXQr/D6JClPpSsqC/eXB/QwRniAjdDcDNSjcuP1NRBJpRbdp1t/nBOFxDtx
+zFVl6gSfFGTCkwocTa7cfeMIXsjBzSkRv3+ZBL/WsMuXd24AlQiLEzRmJQN0Lzo
/VVc7NcEoQfW9+WNiDCO17Z1T4/HAGSY7M/m3xfWZJaPHaxQJelW7vziwrC/f4nQ
48bck7NXqvC7f8RF4E5KLUFhViGYpj+XCxodha8NYKazcscPKa0A08kI7qhWt0Dj
s7heduUBN1E5aFTYhA5ar27zA1xn1CCpNLDmNT0jWYalHpoq9v/GBYRmRhMpRJk+
xCFxsp5i6H74H1vDlebBZ5mcMxypkreoOGTGFrE21xrixseux/Vj5OTmc63Aa6ET
kKUf2relSYJUlhcM9yG65FA2yukwdTx+1U+GaEH6y+ybmeoSOHyPuUKzOKNlo+KZ
Ja73u9LwH+T+v7+wYSj7e6AbO89DmTsYR6tsIIqSoOAHg6VeqZ6PjKB3P6sjN0uq
umQMBw0PC7gheBJIGq8NXPLT+YcWlGF5QXnkkVavj7v5voq5dpUPHlvNVKDjfNkF
RjxuQrcAV6Wi8Sj7sRPPk4HTW1eBlFGj2kntddNTrMo2IKz1YNMXLlI5hmm8glNW
//QzjYEqsJ+2z5T+Z+fd0R3MWUxsSVyMCh6o8vCr15wEwO6YLz284nJHz9hfRRVQ
cXe65xEZ1Yo8KYXmYI3Vgn3XYqrG8VSnTXp/d1LCgxHdl3T8EEeSD3Gh5MaynQ+P
kcSTbExrJXopi+LAhS41NZWzO1smSH6t67BindXZ+SfGcDnIobJLPMtNjJUuBvIk
c0rWOV70kem4xCGSskgAkHX2NbdOPnhhQdVzNZl1THXH/Ryke4rIF4zqMgFyRa9z
ajs1Lgn6v6u+0QAyO4jjpfhAaUzKPldu6IU/SJQpB2qWFsPgKahxzLell2H4XuKo
gnn+VKzODJwScYLTaO89PdCyFJSRWYjO9mUm+8QozlVka00V20UKHlyFVQbUKjr8
sJEetk/GT4QXjuMwmYRt8q9DHHBwO1vR57DSckO8kuKVeUn1eHAOsguj4dtWBnf+
LmXWYRPIWQHgZD5EJs/Jh0Y+bKSREXa4vfRJsEwmZ/79BBLpUS2jZmUtY+p29Jgs
JBQdL0tvGYmbGmExEW4OPspmxbso87GAvMaAyuQU2AxtqrTbSUEv4g3jEuZG49iT
b5v7Wq5qAknFwTeg48jK2oGy+1PVUoJirGRce63RewsIvHkZkahuKdqGQXpk5hXx
bEtvNNY1RGkl+IocZ5Beva8nvQYKRG7RHGM17nwUDV8HblGjNf/qMzAuUs0fHo1/
7h1yZI0ooKMAC42CYLcqYM+GeVkkPkDq3MwNvtfjEdoKQeHdbs8/DvSRfy1MrEGC
f9talJDcItcLH66mmE0vyIRCHqnn7aIGcjzwF04wQG5R9W5zXsSTp6olMad2LNuy
xNzdlftNA70TcL2/vWvZlsFV4sCfqDypvNpj2cm2WEQ2CU8fAGpgh0111Mg+oPqz
ebyGOC+xPtFr0is4dzytoOaMp+3YBheltp/L8IUfEYhIaaQ71i3R1fE14Ze0RytL
nBjhVWqQtpPMBYAVVMhRKHM6ohlc6I2WYbhLuiXqtXt5rh6J0xFCvQXH3iHtS0jV
x6gFXuhQLDDXAimErnnpIUq2Rtr+8uY+/2msD+u8kHRLIpURy6K1C5YajNRKgo7h
QTYVfMebnqDsL3uKs+hykB7Ch6rWDEIxOJ6zKaMycWfTwyvySNRIkwaRJN2kwqgr
YjMtk52/m19pQvPTNkvLTT4KgXea983PHIxyE05WLxcazzqxgoLOMXr2E9ssIjtq
cAXA2IRq5+G8k99N4OJpnVHxBqikCrHwl1+n3OAiGAaM/2lhZfFXPpurogrp5GGR
YrZ8lEIdot8R8vqpuhJDG8zIuTN8A+vNtWEa//XIGEYZK7pzYjujvg1Ljb1QbO5B
xhhHg44NpXcIldeiHF2TIeHPLzSLzVLvyJj4VFtA38LrG1gpoDw6GLZUQvHbW8Pq
4wPP1sO1WM96ktpG3sOuXYaL1CQ76v+6otB7rlzJOXOWyBevaSPl1zwc+gnNFiFX
R+VjTADudV3dzv3hJSfyoS1IjYRqtFX7Iezo4p4zpT5VrVumShFAKmBqb4zDGVYg
bX80WU5MjrQgM8L2nr/fkkDk5dAHwNv3hjVUYEOKFZCx8bBP6yZ+BrZEPoM8waoA
tUSf63aS2L5ZTrwkprieOQqDHp7R3NKvRdKKOdwQ733lPT2hx1H/XekcpHgfUVbL
WrYrBJBwfpQhrDvmBeTl9aFF/OHSGTNOHwdgTtoUga5OhV9G4aok6BPHjPkFFrwh
t9YJpjdmZRb58e8W3SsFth3MVYvGJSxoQNWrlQmix3ivQHXVwwlX6TUKKajfVLWD
43pyaBPRcKWhT8W2XaXlL0jXjm3lT0VD5zlIVm/OnbkJ+s9IAp/pQ6QQ1w5Hxvmv
bd0WP3YAKfFymDb46x5anWJ7+i/GX4Hu+c11LJ7TvYcsIX88Xjd3f6Uo/4tpgLQV
5HEstttkBFrtlKIAS+X0Nbcupg6cAh785aTFJEzP9X+Cp8HhJ3NBNmkTvUxTPHW9
Yyi6Fn3BcdA2W40t8QynnWAmavckEBdXpRo+T4HSl+eTRNzfRjx25g9sr+Cxxt3F
nWmUspY+p0Dff7hS9aLCSQ5uyT3tbgj4/VI4Pq1gZ2q2AiwB6K3WcRdmhvqx2sPY
nIgQZw5A02bsVHuypos/9j5kWTgT8klvrVGBjQq6AAc10XhWKxLnXgLe3EH1rLfW
jn7e+P7jxCPRjVYOWPUNf0JgXYQAE5c+Hmk+iVkzc6EIzku+BYphoXb+QNDIkk7R
E+CMz82ZAB4oGEPc+gYCh/C6G2um0qJB28hkZ/4av3bCfajTYFlc/aIjLHujIDRR
J60NFo4cr3HrL/Nk++frePpPEVwassF6FZ3FpuHANZoAHqMVIKnmwmfhJR5TVa7z
F5/SsGZ8Tzo4+axS8UCg18ceynwU8K9Ca9IoHLIP3NjhAiN/7ZGsJ7f2jbBIiz55
qdjGHli74pDI0ZLM0nkSwvSthXAKDNAoVuwQCb8fOBikJyGc7MW/lLXig2/u2X/V
4O5wV3Z48JjbE8M3lB2H+fJvaKRn98MwchW/mPTRYvj/cJbDN2EL5a0yi7RxaJl5
vDmb6ZbyRzB+tnmOThS1uCa8QfodGhjKOaRCyKdUNqJg3ldjSNTU3LJhwV64wS6D
v6+vGtCtCsf4ns9AGIr4WJuIXP/wcrf/iJn74SxQcsR6jsQ1pevTQE+LqBmrffA9
Y7iZrHggDLfj+UhauZg/2mmCKGu/HZUMIonOkvIOOobSwQ4BCRm9cJJ6NFPT1MXs
zGBBOSozvbLpqsDD7dDC2J027dUmVoGbZ4FB4/PvM3vY0Rn2LbmYAZhVr4musGmE
O/cIcPTD/oZSqov0V0OL9IMKGOW2D/YwMCQqv0nD0tQyOtEJE99iCYcRumd8oTh7
9pw0jCuMmQGiUBOcGLyG6jKvRCbbdZO6/RA5WAFZJ7ASaB1hTbUg/atHSmTejZ9y
qHO8hSla+HtTR9ihd3cSansaNwvEt5sEXfDcDR3vef7QbNkOJ5IkYmgTXU5QEVsa
7x3owx5/MTbg0YjODFQPEJhFkjrUgZG2Z69HNbCuYU4AB2bhNLLGZHKv1wMiXiqP
Iw8d1KRZ14zkVmu69dZBWw+VuQbvfFUfIAHP0aaMAH+7V54PxQfSokK84WzAplxT
tr6A1mYvQb1JNTjxkti+eKFP4Z0dM0CjmZT4uwOAW/mPHTWNEX7cBuib7VfscxQI
gq14X4COZE2N4ZBEvvOqu075f8UOZ6TwLPbAhQI6I10tKZNWUMiEjraY7v4Fxx8k
YQlWZb6E9niOhKaHMRFwS+gd+Yh72H5o1i9KJihJU9bTmSwLcBdonC/S5zLDUH+K
0pSAZ0mh9HACeLaZNpAgF1ISP0V+gtsyHC1XUc1CrHFbD/3YLyfTgPhSLY69SQVq
aFAo4xJAjBj3AOEjZqlWgBPsDdPaZn79d4n5hnb/NFvV9LwGJ6KlDeNIKNT8u/cK
/aTwm3ZUFYP2mLoE22we9IMhP15ptBStd8EE6PwyjLzuKmio3SioL1CLc8XDkGdX
WhJFn5H/fRlFeYjMxyo1jUy0xLNTBBiI/VICGd/ptaT9yWa7o84ZVQ+iFhH1mnfd
WdxFVPrrGbxQHdxHXHZTfXtAudGiYmRM1HpMIKguE/RK9VfDow97ncoj1PnKt/LX
oM7f7NQhp67Q5oGINXobpZLoG6gV9x+G0eV0yKWVzwO7Hwx1kKKhcByiFk/YFXS1
2QzX6l5yDGHtHnr2x1Lbd1XUNVvxwByO4C/o3MPSW7cmed+wifl07WtIE/GASCWz
8GHYCnSq8x6dVfMoE/VOSos+azQeyXTgpMRaMgmYKTE4zjSh4eyGPRTGAEwQ+wpV
GABIUiDjSemBsFGbbC8q6Re/UomJO7nfeYSXeQav4TZJtuI1VHa9MjvqSKzrtgYQ
Knm6HxhXMg0o6wZeHQlme9gY6eAKdJ8gZMSwwVVSNsjifa9yis5QD/T/pjSEzW8+
Xh9TZOH3R//rkkSWs5VC971YLhDZnT9/+fSIKZq4TNOr4dkYMLXH6AuNYe4avoZH
pM5zED8R4rxuoOjxIUmuC0FamK5YyfEzASWpRbxsC9K+EQ8f4m0vMAGuVInVRQd+
koDwPWw5AxnaIix0iAxGsl0bPWidDnMWAKwNt2Lwp20Ji+a5QNZcWoYqZ39qSMh7
amlOpDN4iXly3GSb6ZUPbuNBsfKj3oN98Aca44dV4pHhxJuJe935idtizVncxQNr
Hu2TbKnGeh1T1PZqLtTzmsNe8OlWLf2NJpd7GjK8qxqnlLxSFBoWQdH55NAamm6U
0x+BoA9mL5+09AVfzPR/WnW2/1Sx/lcP64144Gwn+29FA42WIusrKUT7eoQ658ac
UAGieUK068QWI/tj9xWkxVmEym3ieAySvVE+/9DQinXDuQAObugZ9DDTNpcngZ+m
0RHQ3qZpsOAVVtlsKbL3lccSM48sGi4YS13cY3PyrMW0Svp211cPtBAHFh4KoLtf
Fn6A5Smfh8xfIa/my8iVUeFAXnXgYU5zCLqhFA7z3+rb3qXMVj2gV5BjMI9nNq8P
D8SMqRt3EjTgxmyOIouFu9gtO9l/sePHGZm7wAuNqMxJy1tCZNea2XyA6/b995Ps
qnCPk2m6Qk99f1PMmglqXNcfpdbDfWyqoAjT92LvULLxjt17G501YyDIZkku2BjJ
Iq98LufbL8IL9+PBzOYxtQ91X7zBDXR9pOdGQY7Dl15QLxCrPbDgqUG757Y5e0gA
zzYMcf7g3QR3DbGqGBsTtgF3uAfAeExZB+DZR3IXSiVaObpWiOnyDzDkU9fNO2Xu
GiQ1Mc7wApJkMiuzQ3TXvhsd4bJBJOsAbU+HV8loyBpDAfAs9fvhQCei1c8Nel12
YKbeuCbwNuQ5D86XRRUqTMQ7oPJgcC9p3RbKOe+BWaEgbFNJP+qhf1sl8GT4d5Rm
39mmMwZI/X6rduSrjkrmV1AfZiY42y8FN5mcGTsp5yBOSi2XsqN9A+iSA4N/13Dd
11sIBlqJQI/CVL+D4LA6S9VcKlHv9CkDF0WLNVdXY+UE6v1ivVHzaLUNvH9Qlq8Z
rQElHJ7E5mawsZECc4jybykL4iRmlXIjbueqXf4BfCthHnFiZtI4S1B5qyjCGcVD
FBGCHZ31ZXhJ9SHMtrVTrmY69SAub8aQ/bUApzFd2vsXeBI+nBtHlrQmjUQ13x0F
6FXp9m2Q3tRMxdaUdmhP9kv4W0DaHI0VeO7d+3peU1Ajl0DB9XytMMT0mOtNCjxU
1bO6aOE4TtVLhU+7kPIFn4ON3q/yzFAcd93Zvzpcw7HHn5d2brTiIRvn1qW5YHdQ
VOe0z6h7QlrwY1rcc9vJtMXCyjzPCnYWI00FKAp4t95wOxn5NO2mA9ZmzTOHUSAy
RzSAaNmXe3JrkJnFnWcYZqJ9Fjwo9QPZtGXL8difIBcNO05rznSQ1NZ3nX4M8bFs
fLGeSE9G6CpcbR0brB6nY0ehW9wdrDVol5Ew0lRz4SXS0aJhIgUsRwASgPGZjAjQ
21ucplx11teBR/q5eKsuaW8HBQI0sIHBAQxIVDYRpzaPg6wsWTZFpXoSBRVddiEe
W04rAgWWA13MPKwYr5HzzgOU0Ic+DvKkXSW1qUGfAr6SjSGCmyszkVavyirYVuAs
vrVvaSov3cW8bKypH1rLN4VuBs8tJNB1d2C6s/6zqwnKmeHBedknlqrGv4x6pCuR
9VRtBk6LDzi09jo/NNXus1MZar1+NzOPz93jewEnL5d1n1AiThm1jaozG3tzKFu+
AdfB8TILG4dqsTTS4dER4bDnY2YamR5UuIOOSXFX5s+3hjb1qxLHOOYRiC095vYy
RdM3ez37Eztr+O+w4GcQrAePU/QGph0fucp09dNCLyVR/f05hfVLGmwahWVK7z86
yL37jAIx70PzaTpnEfDrcvZum+AN4UeApgne+HGRgeM/XNBy3EVRUDI0+gG3l4kH
uEL8EmWOfIlirVbDkzbmndPZE5hhiTEEO5Pw8DRakXdBunUtvfRim486EP4enTYS
mRgVjemOqU7iEEvkF0UMkSBgPlzAOYf15gCDnNttZhE/w8yHvScOx5+TWIUnjGvY
lkt0KJdlRC4djtB5bYl3fQ6gcFi+PtH6eGK0dD8BdbU6dcDzGBPRu5xj7lxyKQxU
scUghzQFlKU6Hmabl/YANp3DvfOuoffHmuB3B5a9KW9xvi9Qq3HNBkkq6uxiLkcK
VLP6XPBvAiVLC7Rmuy1u284LKl3120Z34Ua8+Iz8wmInafu/L7I2q8Himygclw23
dtk9dQS6NG+K5zrJsdPzh8hd4zzL2cO/jbRPskhSosQs7at1Iz9Neopd4ofRCUos
aR1TsKYyZs15EYhdv/6N+k8exMlRufoTQH+iVHPqNPjKmXt21Qay4rwWEJK3RRsF
ivkyJ5GYAos72cCSoy7doNgXwpZy30O3rn0OQpkLp2d1gcSdyHrKIlFKUVXB8UoF
8fDt7HO8DL3QMaIM6ptfyV6NBBgHAqhr4CCD/3qAKue9QKdyGHTVHMwukOIfomau
y5K2qBH4Q5Pxz3pSZcxG4AFH5FTfIPatJ0a92EofIHqTOMnNsegmyfCpvHt/6jR+
h7LB6nrctXmTr8lAjOUWhD4bEk5xQCVfBtc4UjpfVfE4Kw5yqh/LnY0ViEvubYDT
UUJxSMsRj1e2zoTC1Yuo6FydKe4X+dG83cGwo4exILmyjTYCsGI61YwPOEgpt0z0
7ThGnMUheYq1Pa3eFU1chDiJQl+XioL8LJLRJ1T/07soGUnfzZE1PMjltdtGP/v/
BpPrntNwjVRpDEw6AcjatWMY6jx7VSCu9R39B+vOZYJal+SlLPfdXQDpzf59OzWt
LZVw3MiftZ1GjYIaofa+fAcZ87D+/H5x9MMjQu33CzHFEJ2P19UwEWDgyJTqY0QW
CYLRHnCCDN94Kt1KDh2SuM+JN45fKbCmOT5tHvirrdbn40z8oebvAvuXs04XZiMb
9pjCIdFN5EKTV+AlnxlgS+//V343qdZLSt4pe8BNB05XfbGAbGRO1nEZkE5mWhZy
UctHPNAI22zhwJOYkIqSbGMv0MtedRMFZmme6fMRFob+Nmdl7Erh7N87kc/azbxN
I9MNtdmUmvn92PmjdgIknTgM3yHvWHg9kWEw4ouwc0zes33j5PEGR2nFg3gWE1/Q
vF5xFdeCGIhPuD5UWqVhuFf1hn4valhpwox4AApd0u6ysVLodcOpxEk05EM/PMtG
i+5E06hdD74umUSf9LXZi7Xuot8hmHtwYYBaWEseN58ETwPA43lQe6cdoDhxZXQv
AH28v+s+wh5hohh4Ita08ugIWKg4xp1NqwGE3DImVEisEnIMyXCrFEPjxsCS4rOh
xqrk4lfY0fwEJmxDpI+SuuXRCBICAqn060D7mdKWDjMbx9JEriV+4SO+z0zBsz/S
I2jnY6ETsHtKiZP0ipucPBlzrtEjQfLcWOJJmKPW0EylAuDjgElTo0IosnzTu1yE
615Xrt/vuy9Fw89e0lpo6H/l3m+RoHdTPdaCFGp0Hmk3cRc7ESEPQUv1KhHXKffo
NBMgDDZKzKmWtYrVr8s6XiC4c2W3Tpe9x3k5XNx+0VyFMyAKgXMpburpFOL4qMD/
jgwzvA6kbL5AX+ixD/kLE50bozzGqy1efRei2DmN8k77nkU+S5RMyAha4l5RGuYU
fZSOwy0YTseBIDH4mCDuKbBGbDNl/v/1PXoX2aWVwTrYWQAhAr+D2h/O9HleoJGG
+FyWtilMX8h6dTiNnxcFQfAW4vGoGSCr+tY6RV0Zntmysc0liDaWHYi0wYNlh5t+
1f9rqVfW+M7fEtS1vCgIGdIfRm55ZwEluuS2yCRwpTN7vs2lGpUSixiEVnofbe4y
LgOxhNPrmr6johyZ5z6ghWLL9tdiiydTWFjzibhfHsmI16GQ8joDCXfLPtpLZQBq
1WNpPDkzwmfdg12ARtOhbaYxOwQGQr2iUsHDFAn8ajlMZETtCeB4MMsOi8Goz22P
NzxOHD7GMGujxssbDNo471dfswsctyU+sIi202yDCkORkUfb8ZOfoZGs3NHJgdew
uVtJaqgAHMdLjf7XJbevwN7e0Ici0u1LfA4FBWdgiEF3olktuEJi7M4KprOOHYet
e4PbRmG2dH8tGPA94VxDCwNxrJSG64rWinbixzC536HijiJA/U4Pk/hCBUabSipJ
ZgRKne4vnr8Jkrqr69D7ymu3hUQBvXyTktgOE9UtWU/Bm/CNqwImsigYMmr4w3zA
j5mlHsoP2LTNxv0g4ad6WLJT3/5aidR0I4nGMJyZ4ycwXOv1361pZ392j63wa1Fh
X3zZQ9iYHl12PjUrMvcUil4nxA2JUsU2DJkGlUgXzIU5WDf6zav+wyHQ3os5Oi3S
qOEPZlD/Bjjes1FZ3vlJHsMT4RiUYZeAFDSBgspGL/SA2if6CnWSzx4YhHkSkadi
UnPNCE6v4cjQeoz1LRop+4rkkHFDSbRPJcfGDGfv0T1Dne4t6XMnEoaD9EdzpjWM
bVON1QWg1Os8JBr6WeHjmF+54xLki88xnTYgCap4WS8aET2qmARt4nqHQXyNtnky
ne/GQQBJ5zhnol/IRcZNJVnYulAlDHQUxCVY2i0ETPdiJZG9OiUFpyDGMHSySpHw
TWRUqjxZUfWKKyGz/a7rnDJ2W4CrTNqHB1sElLeM/pZj7zJ8tdyN+pOM53f7xaRH
MKLJmd++s7+7XEkFDUlxg3Z4CCpkIWu8vNywPK4rnLpZbFOi00R6oufJjm9S3PzS
T4haExGFvXuq+LqESvwSwWJ5OeRDkDrgWxTJGN6RR0nC8WpXmPIcda0RLOvhzCrA
5xJK8vsAGVm0cRSOooEG1ZxIvxj4qCGZ16Fgg0pkpcBcWp8b9p/sFQJF97UaDUeS
EQH9y4CpiZaNFyWqt+WWgT3Jujh4Vz/ckbtkuV0xw59lUXMW8tHWZHFRtnfGTba1
8GptkqOPpklfP6072mfatVwMzbfq9LqoOa17O3W71J38BcW8f60bnr7yIMq2lAFc
lWJsSnliF2+rfSOvQMlYH0vuksNzflVCAC4Lszqkdnl2XpCxGBkZ97/Pp5S0VsfS
K/EoJ9PtcgPe3ugoKbkf7MwKzQRMBpigx/VYXmEsPgLHm0Qgvv3+mSIO4dYtje7G
VcOyhDYpsnBIpw9Rvg0WQwpiSluRFZXNIkChXWQyT4Oq5ICZbiGHiJb1b2Sv25c8
R7AlejLxJosfRCx40pJaCZW9wE1EM3FoPzSeuqeQldRVw7OhWedGTz5I0B6rHHcr
c0olC/GrIZpjU9qNFoHrgUs9unqQu9itlOukeFUPOVFTjuqPuiu5S0llt79GDYjQ
UtbiYcaC1mum7qLl0J7CKWF622RNi1DrL+1vqQruPcubjMrNexMN0tB7nnHsQBLb
cJ0+9eoiIxvkBEYiTNS2XtWSfkGCjDKp10TBH+EtY/5qruvvG/L1kz4L3JM41OCR
Zk1ZFS5fCjXa+38vlHUjKJFPxzyP1knzbvZBuEX/99q57zBzv/xcqkB4dtWxQpKr
OQ8qzzR7j3SVUjbHgBlDNp/TRs7Kapmm6qeBDyzHzPlOUQiy5jVIFI+j0kR8jBPo
gI2iXK+1QDupcihSqMRhHDVQAkUC/ndDyBTVkmn2q4uxk3mmBhW/BSep6fFSigKx
hBiNOpvjoYpEZ6NoUWir2xXmHXuW6xNE7E5sTZ8Rl55R227XCbXh7OKwJpgahwKP
RurEABUTtrxgDL5OGiRaYswnCPsCMwwi4pGYX3+f+JIosqZqpSitvK4fjAHDvtEr
n1oVz/WeJNOQoJkIZmQ9SOyxZcls2HgUiFgtyDSZ33A6ePE6qHgifqY7iOfQxdgb
8Mj4rB5Wp4Nujtj5jaRKEcgNMRawjvp6YAfjI77BWZfer+2y28KV3MIYm06Ieh8O
MgCJqP158vFB8UMSNz4ytFMPIweEGR8v1+h8ph/47JzddgSaeOZ1rYrU0nN6FHDZ
5ENVDfg9U6PFxBgv9KbZ+L0jQM4z0GaDUXbyrldok82pSvWfW/yVZPvfESS1ecZQ
hrKvTryI1Q85eZUkH6rWWDVeqhT1hGpC6qB0xwObF76Yu1STtF67TZ8Ui9jmy2PE
ZzAENkVE5zoyY7AQ5xssHNxiUGBVAdPuFEbKKq4VEx7pQfJpCh/rLTI6DH9R8t9r
9bERpkQfe3pMLIBYs1J2+uXmnOa6xfgUkPjHwGyKrNuLt2sqgd/Fhh9dKeGsb2D8
pWx+p5zOI0b3hWT73XVgKEvCWfYwiBq3fO+l1SLZ4498MgRnD38unBpvvlI70U0y
3jg4BYg+s9COvHLAqJMvxAUxsU4ZIbPWUUKBxYVIbFlMSQze97hAUN7H6G3dqtIi
ACtvAF77T71haTTeqKlPf9LAwcRv3WaiwSXdJJLPbgNbrd/wDbfsZ3ZMABv/y3Tu
RGsnDLvV2kH9E7woBIF1CJRC+OmLKhlKQK+1zh1BogEhrzNMnCk6mdumy0nC/WPS
F29oIHw2T1fvVB8iz/j1OxEuQYL52TEOQBs+3IWUTG7pRYMnj4Dor98jJC1MRb+t
enBSm5/XrQsWd/IkCGr9kpI2or3Ia66rK6tXU7fPIVRijjePmQpACR/rwNBW8qOW
67zKwFZ85eOkvky3n2WDjhjyUY5EVKANL9WwguSdd3jO7rvMA1f8mEDvYHlt/SFP
WgquNe0kBYPuZ3lJ6bZTZyjyJvBLQMhi0T5MyJL0+Q3xwD/Ztp70MSh4D++Og8+n
URvG9fOFA6aZH1/oCMgL3II0SaTsyggAu8u+q1mLr1NNXsaSW4amKFQq92IUhkYE
w8PY/B0/x9d+3kxDZw0TJ1EQbTzKKKV1LPDEOt+KmkViEXaRsh0Hb8ESf9LwIWfl
tut9z4nslSYZ4enaXNDA4UdJI3qV1zax3hCtFKFbNW6Ao1FdaAYVOEi8THGFEj2a
TF8OxTVv3g5xJ4oSeOk3d3ao2x7MeirM+iBN9vyLKwIY/ZpEIg7nHuoH2vVl9Uk+
fXJovLl4gRjOPeabZDpE1V7MwJLxJpmjiE5oqnEmpyCT595IbY6gkliINMNtAVjF
+Ez7ZGmSDOcyUw35B0fz6zVjg+7B8bSRzu+Ep51vzI5rI+q6iEBu/PXZg8TWq9hl
JmXZ7hVdd4Hd1AyKX+mHN41CMoKax+xUO6DaHgxm+t4tnvpYxk6ras+5/ZpaTuk5
/xRWj0iatBWvepuGnKlsZnqGp2MnQTuW+PfkhQBXf/r+v/yf98F/yNs8iXElkc9S
DzdFA7hkV5mkPEUVR6PN/nrZX1+g6JPF9NaS+sJw8UYutCtIVjjOWq0DCwbVYQKc
JxAHaVeKiP2oAkhEx2rBBOG7PaUvyOgtKBb1e4+nY3bV/lXWm3YNH/79FPXE3KfR
UemwUW8dKzf4XTWFbiPxOLwcxoPqzGiYwBf/IWZ2UCo5OE6HrfHT6DfJF/fHS4fk
xQXYd1n33qQPygYn9qV5/7Hu09BpMTd3fd7lUDG8SCcuvv6hw0SZ3RlaZNfYxAdM
XncSpfu1UT3sv29ZTKIRpX3zHPmLwpeq4hwBoVGjDG8ZYApTNG60CrzumV13g4ry
NvXr6Y50nx6xUPCs6JS8vpM0wsgnkLQbkkZ8MKnHn3BtoOWVFELfb2EGYi3w0IcW
XiQNZSonAELWuw/Js9X7PzjLftK5JspP4ooGKQxq1IYNaeOBnzI44GsWYD4HwqEY
HN6NPKiZ6COEx2ndqar7w5uw6+UWwy+Yp0JY8Al1jy5Eki7RcU8Rq4H41/oxXyZU
e360bQe/8lyFFL0po4LC+pqcqB3R2RxjUh4tPTdldVWy+Zo7+QsmaHY/J8XT+jlm
H3DjgdqHBD0FHv08vIzItmOO6iBNpjlkClQMOqr7Oi36Wu/Ah+NVAlJMOJhEOw2P
e/2FtHOjucRRq/ScfrsAqX4InRfT8IvsTMRL3aPD1Sq02nyaHIe7O2UKXwC0D58y
nWLl1fmXOoFNKaKACHPDg/eMdJdViTZLvEtkUKsTViUxj8JpLf/0FYYrgLwLSqhz
xqgvNY/T++0oGqZFa3ZWWvb4HEoRXFCGs7uNrtFg+fixrvcBS4vhKmLmWSewCR9V
jtEd8UcIyzM+32nA8+poP1gJbC+DvtiQcoMqhaRsjDZHfr8hv487Hv4CDkDobUwO
ibCwrfQVc1X1xEDGXvupJTyB/s4cnghh3RS68kNpx9uQSDRxemVyXChxvJlKXuoE
/EukbbZLxCuypCHZaUn1iJUDi7J9+rLliyufnI8rQ3h7JUTVU/lpcH99fwS+6urw
LpK7BHkLBfQby2vJxWHV86mgdZcoqcC0Ti3dH0qV+T6+hHv+KRzo0/5Y2H0RfwDO
XXJ9U6zVuc5SkMJwVXjldXd2dl6CUxAMBh8N8W7yxrmXfV6hqLA/xjgBHV0K9XwZ
IX2xVKslKuGgBtXu9JIjfghJ86s+G0RfdoltNbTkpWidHH865Kx/qglHd1HS0KxB
JnwdKjBPYPEn4G6Z7Mm/q+hpeXZwtXZqEvRlh7/3NdE9+RwWuPqwADhH0ryo8olX
fl28x6fQTGbaVz9O6JHIu4ShfXt464W7f+n1kMGPAzZcsxqIdrPhsJvSWxNxktiE
S+1sqNv4BbX4UpejcuDfcIc+MIs1OYaljHorLqS30tdLeiZwRvQ67aWrOGkCUcMR
ce9wdgE2VEcBzsennvkOTRCpIzls9IyOGJTCLTeD1xIVTvCSuiX0ovskumGdeIrD
MhrvFQ7cnxnbSzb3SIe6jKqgOLSdsbC+F4bv5IoFiD5QzuTn4MXEjrM1DSTR0wya
3CUqpiVvYWg7dJIKGjs7YbmKLmw/JbEBL3GCUpg/R+bxzGd54Rgqwijjh6E4trQj
sAou7I7KW+ARGC4Liv+RZcoZ1zHcu+zmGnai8cn82ivLRnHBh5aAhRBiuKLrSnIb
9/15e6udnOxazcdbTtnggN1GURqgk4EKgFAm+DtcKxWLhXNQcgH5uYhrOlK6alJ+
wdvDLDR7hJ+0Tp5HhrYDQn9aJiBpmkO8Fk3cSQVFPZJ/2bjiUFXoR+wlLCQqh2gE
adzvmt3k3hd6TAiSPdk34Tr2xgbzJphaNL5EFYJh2oub9hOfeVzj4t0BZfbwJYbI
768r+NLKnzGTG828zSm2v7nblORqVUMxqolomxuuHvAoWhGZp6idzVyfXSkPBbcB
MWrU+pR1t1ByR3uFOUQ0+6T5psUDvnfmEPqUSCIX3GQrJeGSjYNDawQVMPQBubtO
Y+XLGqeKehpPEBK2Sc41Dtk475VI962cBQNYxYa2bYZrcQAznSX7i4yNMWUD8e/Y
/KUCvFIFQwnlXTBCJwJr2As5dwu7NwZYSaH6nBDwb5UMQ3u0Dj5j4J/E+xzslIBz
ygkfgmTBIlj1sjKBPEeK3W5T2ptTpcvdhR/iiufxjeIMaVevlJHrYWwJnYnFkieP
+KToCMwe6HaKHF3G/gwvNgwmTXnqPiA4NgJW/IOR7aNNuFd5xexwzAyvUWUlGLqR
xIFKWnIpwSshMFQt0VWyfiyZN68ZqzTpBI83ciJi1RBAaPoWFZ8Ey0tCHFuxMhf2
gRYjqFDo8EMrah2EPwP6c9+/STSrZuTtDPQTjIvKdqMnb7ddZjDM65HuVj++vOcv
h4sUhq76sn63b0NA9HmN05Ib3I+YMOXpThrhdm9YcB/ZC7MIUZsWDEAFrRDwRYKV
dz2S247Rc0KjomiQTnJ/N0uPpsRL8he3KLqWj4p3Rhm9Yu89x7jS27neRLXDzDoE
5r0e0QaMgutWcFNBcaOSJfDWyL9rjTiu2v1r4F7dbRqmWSTQDmnC0Sl2u/oD4neg
JXeaExOM/KlVT3fP0eUxjLgG/dvkYk62jkJa1vxl8lVBkkeS52ZkRwnxpg+We3Ez
pTivDuOUb0Dl4EpZmBWoEcC6YEJxTjbceHdOW+ZuF8/0VYX8ScK0vInuimCnV60i
ph70D9X1tRAoNHiAlt7ESEsLo5Zvku4HOyHcf0An+a0OSbCNaLGY52G003tea6vJ
+UWxDjGGzu0rmqHcNlJrd8ax+ys08d829G6Ktc2kqTgVy2hfjrJd7s4KRYjc7p2x
DgHn4mbUGSzz+V0yJ+s5RPz2mKSYE0lryR6iuRvXAX6a5/RDjkucugBWPE9PyhmA
IUKxeE3wQJiUWZaqvISFuVbM65gEQjIxkRFHhgA7CXXgvuWQgjYJEbjfkB0dAmgb
MFaEMn3bpTNLv06w5OAuehqLQD39OFvFqRGZi/twshI9HHQEludAMFuLTzXVKZi2
4EmenBtzTJbqZsKGWsHs8HkKo9Dd+35EBWc8ymqukGB2lZQ3Mnw0YYhmQdQiSkHn
xs+aL+0xCdapgCNnOXvDnCVE0xSVE9dsCo3Y31rtCZEkk1j797un6wiWjvRAM5Kg
QR7cH/wCBw9XjFk2+8iqyyqX8VQXDxYRDkcR0ejfNSrIUSlFm+NOF6Eh3mpcEeq8
ERetByZ6j6DJN0wI26yzZCIoMO7bLXH3jza0C+HbMlDLkWPowgA0QmmbGXmHsphA
T12mql1dVa1EYtMydO9IRAHVyBKTJzZ6KWoUAeQ5XTo7r2W9DatCU3KIGCoAjQY8
6G0GTMt2WZ1zvlj/LCA5/yXm8yyWxpGoo78QPxapndbb2AEm4IoXfDJu2BdEnaRg
bBxTHuENs+8PKbrdmKEN/M5DEtX2V9YTBukbNYOugpJMHNI6FnESkWf7u4n8qdal
V/IlC1rVUJCweGXjC6ZiGYIEP881c1vLAHj/saA7EzrJwjm2+JYWNA7sfuyF4+e3
rjDK2PiFr6VXOPs+UYxCFZqAQUsqYH7B1pTqB+CX3mD2boMPkGOKYkF17XFntehS
olr4bzngGYs3xnXDnIj9VqOS+xdG7SJDdHhD3YyX6fWHSgWLWESR2nus41ikYtS1
5fbOJABzZiPO6ge5ONPFrJAiEkYTOpSHd7loi82d8aqoePDMtYfd9dddEIClK4fI
01Outed/mNCFgkzUNDZs7IFPrRa6wvYwWBmkp8hfrxc1uBvgvNbd54oza0tqzZJt
atXFSXTbRyo3pjj8e7uBQNFZ07YqceY08EYiyRiOm6ty3mm5mwWBLwouxPgpqhm8
5ua02MqxWbSinKPIjMeBW5mk0QqM79hfl2xS+hJ+3rvfVSh14idK9r8qimSCrh9b
s/NxiSC3S6P3Iha6BwoqifDNGnTLVPmZ1HtWMEMoqkOx9NcMLVZVBVkUwS+qA/rw
K6NhGner9nU2Ib6lg4m8f8pwhxU9Cy6h6zUe4gR0hjuKZcQ6lrgs8AnoS73tuUDQ
kY96nIA4Frp7GDxNrficZCULk7PpaIsG7PwcP7PFLcMIsizlKPxf01eeoX97SBu1
Xkzm+V3zyf87Hpl1TPyCnrFmkjwr771mwhaeeG6FSkFlE4ZtPCwYIFALF76r66xQ
QAXyHncNYYiMMQNKdhx7jIWkisUflrVTAdewzfloXFY3l+YI/4C33V8at65+korq
LDvqeoa70AXIkCUliMg/YPYlLPAN5WY+VBjF8l0cfTgJjdzdFLFv9mARqfOXi49e
Pp14JAg5HGpFki6+Pb9Nby/hNqV9VN19Z6sH4uflR2qSZHovm9+8KEC4detzsvet
qJ8JoAUOhAYVMGjp9kdNp9CKJGGq/mvSLEiL6p7E6HvmzCYPPby4Z9H8G704SV7O
x8N8q30qm45Y5+Dq7QOhIFq6b5m9TkHRxlTfnmioaUJbYb1SrBQ1xXBc0YpMxKIn
S8GAEnc8oHb+uubKwcSmZ++3sX1b6uUbR682DY3st24pD9zGeb7gOj4dJhJhKALS
ykF43MmWDZ7QPgHviJPYeer64eyY0AbGVIUprovHvI9EnTarPRAPS9vrkWCfjc8T
aMvTzn4heWo45Tu3qmMvsLgK+79zl6JQxqAJeqQTPvrQaKXHfpXRY/HHrfgYBOiS
KBBYm4Ip6ctRH729qEYTwmhe9iI6Vp1sKf4zSlUYWMsQjsn9q8QtQUuDIFOlIssQ
ayIsuE0O2t52xrmh9jjBUlIS8TGqVhirHCzKJCve/bjKC7yPLzjA2rPU4Wvo7A1d
6lBz43mmr1h+Fgv/hVzbhAvQ/rYk1HzWP64pIdNKNJc5WFV5L34AseFXgkXpkLeQ
EgR7ZE5g8dfHfJDpyaECi9q2X6D/hgfpprHz0qmdi+ZJhKv3kSN1vZF0Od9MPZE/
Oh9ghnTADr0+ld/Jyqx9kEXI2RKbIqhZzGYzNC1rTBUMObTVhz/jvBEnkrTIGRGQ
udY+bTrQr8DLAf6BssmkbwwqQjMo6Qst1TOHPf+wmbylDMf4YqsQnriPfJKBNR00
uIsX1ZH4UCn5lvIW/XvMvhQ6db8kFQkinwFEUj4LCKatWSSbf8CXh9XldDIXHjiz
0XB1zAb73cTXICxR1YnTYcQRvNaVslnbVjsXBsL3IlQLFoE4tGgoCCmBu4S+zbFN
WLgoC/59snOxqDfBoh5VGg86YR8j9XTe6B8bjNU0wipPqU8EzTkTxwpOhDMrLY1c
QZXwxPm4ykgqEZaaYR6yVeP7an4b6jOazuqYSb1qDPSt3i0Goh5BO5y8llvg9qVi
xHOvxbAZQeJWpmdZTfKiBoEwZKUIUBfbQpCPQmwnJJCUZXZ8mzwV7Cj19TwYRUhH
39ICDXM9P4cCkOL6Lci9Pufisg8PXzigETg6Dy1EhVPN4nHlhu+NXGI7OzmgtxkB
1FNFKJeWhLurxbvCa+n2dxNZaLHZ63/KHadzqUmWhQm0zQ9ssdwQqVABqtrLIJpN
AUM74RBGF6shGePr1qZyCGyksWVTnY91us9ebYMzuzKVQ3uWBRKFbIpOMNb4Bnkh
eJU8HHIoiyp16jlyXHsSXCwbduMWZskYAG4h0Tvm8mCTAKWfUHVEJLhmPJntLTYK
RbZRnETTVtqj3BrdMeux+BbLiJq2VjPn119yvjYFlRyrarLFxlterkYFAJfM7S/C
az8Hg/1AyEHc4yoz5HA4eC2ecWjfGX4E9q7Oa4YqNWLEgkLe3kF2j5XkyfanQ57p
QoifbLH8WSZ4SiWkkLkKrIdT5XLTsLr1nRXbK91ijns+ev92TT2VKh2PUOLuNrCs
SpPRUBECRgcDIoUtSJ4y0uuSDo/gFlQPwZXffRqhChYhUO5FSbrtY05XSh7wG76s
mZflVAZuZOaTLCWZ+cIRMC2cpfyoZ2UL5gkFceacF+B2Wcu7mxg7nbB63dsb2Eej
KIj0R52iBr1YL2LckKdq0ABBL5vz9E9hsr1a7lvfHeTTcOdholElUx5y3AjYkVUc
EPIpAKBJ49Xw/lwpmQ3hjpUcVSmO6oMWFrcvScueN3DtKQof+w+Y9Z/DUAHocDrk
viyNyKcotwRs4WtQXYZuOJna86l1lf0KnAs4jVyu3r0EePk26A5vEKcQOeAqGi/n
rk8pIX6DV0Xr5s/GFhtGB5fxE/zXrvVZKx7s4HVa5WSPbW7tQLW7RWVv4t/FNmbD
vI2JOmNYB4wNn8d5WQHru8SQzz3UxfC3kzsfbxOgKJHDeiS4GRBPpegDnkgiBLq8
WaeUO8F1AQ/x+D8Fy0sYuFEpZVr3re/dTDMchKJvxC2jfaxQsLKkEnY4u/DEhsI4
MEZn08X5HfSfMf0Im5+vva3L5s5l3XbCiTLo4uTTHteGAmsH8a9n2dSkRey7dPoz
C6kDGF4WKIsMU50XvrNZOA9T1tZ06wxGvFnedyYeImuBHWhq+eTGnVaLFlmWa+Ib
r1NjRiZf1wH6lawWpZcLDVqelr0vXIUE0c8RfUzoekJe1ie/nzOS295ZhyjHclJu
QiKxeH54nj7laL29FBjr0Qi02d3xf2UUD+sCCi/A+gnEjy4tC6g4aRRjBqWrGziG
j2ZhCvOLT6Lv/ZtwytXfMlcC765BeR54ObgDyTkjUfo5pJL6OvX3wQtJrW1fDYeu
t7/yyRDhe7N6sC/Qm8aRpclbLBZ9NICS/Tu6rNk61lRX+ZkWB8sQg0ir7haqub3a
0DddRucmiDxVY22kz1R6+RaIkalcYtSJkncfDYA8hjDIgntE3hJIKSpCK2NmxMWX
HryxUNNNIBCyOcmBszpbSK8SzRnEx0G96bEIaj8knEKrWjHHhicoGYzDv+Mw3DvF
KY4DYAocNPKYJHg90wIdF5JhHcpOOB/SWxFFr0GTI2EvP8jpxaU1cP2hq7tMfYfm
iHVwiOj3Ov5HE3TOk9CVB6h43UVJHzmyJVKX9pxHoNyiKI+g6AYCq7Z+BPc58S0F
u0fXyuwKAi/Fs58nEzGIanCgaUNDOb7wXruQhE+yU2stN7/Vx0ljlArCnzv1QlQA
nbzfPCdya4SWmNhZULqNdAo6neSU/JstBvIrPa7XJuf8x9sKWU4BD6HqUN/JxNs2
AbxXKx2MQOB4OR/eCUhLhuWw5CSeBmDLf+qYk0rYLnw/nN6dmEMt7DRxb/y4Gqpo
EdRVRIooObdIEowinpN3dgvmbzsZwGXgzfJfzi0dz6dMv0LELjouuVVAGJEmTYq+
kpcP0VMUHlHfkHHUYJsBizNRgI4K9iaqkEpOzAu8bzlLXYGPuGIalSTAMZLxgxc1
1WRKYGkRDMdYV0KxIF20b9hoTHyi3QSsxXz/B76aKEFLKl8oAqwMfGx0SQXIFETv
5Mp8YN79zOSavA6e12OfpRxOLKJ8Ou4GILVXvOo+6o+2/Pp9GkNz8K2MOBKZScIf
NSMLVkmbcex2FhyLP+J+IkdeU2XCHQdv2j8+heMq0S+OUbXNkrtkcYRbnJPvHQ0A
R9ATYA4HqneRsSXcknv8BcP+JGgXsgDXZdEk0GX24gBClXIkTBdZ8J0G4H9eEVS2
JRf4XV7GpX4vchWndGsXeOQ/j+IPO2ZrD5C8U56A7gW/RmXxt5C00oMcZWb77zo5
XmACxRvOs1EAoO98LQ5inTtXTdjiLKAGCma6X4IT7hSCggsRpFiVY96Rp+K4KAlK
ZE0NdktWsfs8bBG0LaR2NhsmM9i/5iIHO2jZKS4bRtO4fB++U/h61WR/MMoMse83
WjnLyiteI7yxEKV6z7l1+tDdu4q+XM20D5Y7rpgOSzlJBwA4WErMO98kUE2IYFrh
Y79v8B9Azmc/NFmsBWR95HNz3PIr4FAqCIvU1aFTRwpVcH9AzkPOH56KSsyOsziz
iahUoT7BbOw8nboy1Hh2xQAfGTobZkLaDsc/bD4EbrhivkGHPwl3EGeXjnFaYZix
1sbXJA9BPjF1iBbFHPonlZebC0wNe3HdQisZtf3c10fMmAvBmCY9T4FEqe7IFtOP
edBElGF4Yu9VRIdmCAThK6OKqiZm/2H1QL9F6ld9nBBnswF6u8mJyLJLbeyyML7l
r0TKCi9bjUuN+wCXR3QY/3BN8cd8b9MvHPHVvxQLAkG261LfrBnIuTJHNLsGEi74
ooquLiwO77ynwH+XkWWAjaiQp9ErgsvjFuKA7Atz963BnRnRrS4TWHlJ4BkKA4Dd
cxoJtCJUpCAazO3ad740pKyk813clLiq08MukP7pcDIrrqTCNWFwd0A3RM6gvuiH
6wYmq8laaZsFruu32lFwT+qvS3lt3p8ozfZlomIkV10wPrv3c9Nrp4TJMzXL+uua
iNeNWdXZC/nXAN3hVA9RUT0hIOn+L5gCxK/GOgJ/UzUxcmAhCCUYJKKfjajOPMng
tBpzrPgghAV0Uf3gD1fR0ioIfHGV+NOPqPyC/hVepiPL3CkU8Zo931TSYJddhF/F
9LJJhHBM2V2DlqAt670FThk9GVF+xMZbgP0TY/yFx2tfZfz3UyMFQ6Mdn2g/uCJr
JtItdF8qu/2S68RnwetwktmSuI7UPrnCUb0T6m1DCg3QF5Q7Q70tp8EclZnBxQgk
KEURVzZkgQ5i7FnOy2bHrm/l/h2n73g48W14KebcfVYgRgs3ROgFFGhGDlec3Emj
QDncCMtihzvxhrTKRDX/hiPbulJC3l8YGXsNOOA+TOnmerLzLf3+UVjxMXHswoDG
AsbNlDiquAd15Yh1TFowo91J2WzvAiVbFb9o803Jv3uoqHfCChBNJNNp0ZlaxCGn
T1TjbgULWFk+qFDUp+Dv7bgUjKXtD2TjT5ZZ3XtoUuXvvTo0XfTt4bbBGG+oYZn4
dcIOMghQfyzqbFj0P9FjhD3Zymk+QWbc4Y7oOD1jvg9TxFr9P/dfkFp/vHLnUSrV
WM4ZQGeXCLg+gA3gZJr0bOv5jAQX/IFCVcbNljItVpKJ3knQw/l1U7uO1ZbhUD8X
bEQeEJ1Ci9bewFJYYiKy2XaZyoQIojnKLYrtJuZGY5XjBOogRoT/C8fxoRZBaAQB
WFkdTuqew9l3Zh3NeyZhyhtj1uPhgvrhuog7c145nPHug6CrxVkx7cfQSWr908Yn
72KAhEt42zPaglVIMqj2GpQTVLyZbGI/M2n17L7E6hwooJrcrsOnXxIsVSDlrHpD
NFKOKCZyL2vzTTeljOjzg9VqzS9uG88/JN++ddTRWzunzFEbsT7N/MJMJHLjQc/Q
2jM0OQ6VW+tebtUzLN6rt0wyFk2/0HKSpC7hvhmOA4b9ysQ1fAde0/gtojaXAb3V
5orkifcXsJcJHgj5AnAzWEezCkk5AAoy6uoYaRjonxuiVc3tFAhxHJHt3CReuBzI
I8VnIRcUebEhevWR7SCeCLFs7FXVa/gGgLTd5mfIFj9RET20njSlbAfvuGLbAytf
jsKpaHGnSD3DffllsAF7o7kVUvtbshNebukIp1PbEm72P8Xs57fi99Qu5Yl60MgF
omYsl/he4HleRt3ZHDcvZPvAtxxjGYBaGQNjXQpEPxKN8j0Zm8QR3cNf6QrCEzpl
pDbFCkKcqKnaEbRF/hsgikAeppJqkQZ0jjbNEkJd6RlyEHOLGpT/gNsYqm+5suWt
2rxe6ZjkvbPHUnY70YLRI5MQI3Dzm7ZRac2c2bLWimpLwMGSHzM2nbCm777awwcm
n5XyKwofFcVT5T/XsOAH39HwCGbFcZ06scBhF75T4nBaa6RnauISDZwrFhEmkrTY
FnpjXmk9nh0+KzeM+NX2K0lL6oOgps9IBN/V2VNHM0Gny2hwa7IfLEFU9UdaAX1H
CM62GmlQ6sSaVYhPvOVM356/bYIDHswEkCEMb0JXZy8/p9HFMQRO15YnsC5TbB6N
FZqk5H5PsDkOh2O0beIQnoBRsNNHNFwLBlgq5A9x2xXNN5msF3RdfcaeIZIyoe7G
YE7ZB6JjB0I8a1CGKewfTHFvw/S2R7p30Dtz2klruN9hUXWy3DE7oPtz4in7P1P0
hkI+81xIf713Kw4rB4yUfGKBO0iqvvJNRd30UeDMNq/lX/6Pbm1Zzz/qyPwGzjZz
6O8hk1oPKiR7VJ8XQNTIgJv4gRH5B7noQWp8S56c2L0CuCfL5Pspx4me2b93VRiY
PjJ/Ar3QM+fOcA627/812BxaeXtOJg8QsD/1EJTofI+ebL+5lRyfmxx/1kYypj6X
n1jSvPLfbIgtU+xqeJn/dRsv+YGPXwkJlrLqVgyvxXr267OLjrFkrkvfhx+A2zs/
DuzRNUG0L2jflm7zED0XpMRLRFba/oGP+gZO+DVYPL15lpBZsdsf89Dev+uecpiD
i7R+Z7fBsHujcfzQSekmQ1trwfwgTMN2QYMf8gRl5Nd8sI0k/6Mi26HlzzfXrihm
q85lfozzyGZjWS32rVUjAoCI0Dq6gzUo9mrE4ETQIAFNHx3y4rLmjeGP5YARaGnQ
lYaV84of+UdfGfXWJZaDcsYcsAnnhZWZZtQXxDFbqZRUseYwaQ0QcwXpBPWI/M8T
3GAXlf2AeF5cubP2ALHCN3BvV8kO9Qzky+5qDG/mgGXIWBtNkqWPmiZIP33NQTn/
isOttdTl2omN2jHRmp/rho3SjLHtzEk/93QB3HzJVCeWI+ZMMbQv0B9xRwtZgpYh
mxqah82gX7O5+hQ0DYTYf/2RoPFBjnM42GshggacKAhaU6R6+s6tIgOVwLQa4PLD
5i6zzPhMeLpEN02z0tkFTpMPTcW8TBDi2ELaArKJLtuat6g7I4LVcPCYl+C4JtlG
fP1yu5oj/ALRpOZkbD9kIsRs4ltc8vpNtfFL8q4Xa3s3LQgrCF0R1aS6cXjSDJKK
HbNeTczQpM4U3uSdPRJ69uEKTUdjUz+Rv5wisGLaZqm2Y2zMRqdTid2ZYnEEFWHC
XEvaTcelrE6+8ifee4KoHubrZmeC5UPOivEHTi0PXyYee2tYIrzmYF/fhYQt62tb
A629T6xCMPof5kecpdwC0V6UYi5NLopa4jIfrNfShiX0+0smhl1CXpQgwahc7Ouh
UZoni1lSb2wtTgwQYIrOQ70kzeBRGQj2Fo7WsdgnWYnwCBM5R8v/Kqhi/wNzzrsh
kidKmbK2aVpXt/tqTtgxcGYW6E/XiuBhMK9Ic72JcxzuQpNj4hdOqMtfMKa93GLq
HbxK8+F8VLGWyf0WqAps6v3bQ60uHckfNyCccObGl/TG1rd3SvooEqa6voa/SAsC
4Q7xF5c8bIK+ort+e4fUrgTEgycIeq7c5/1hYLLYDudErx2i7QeZ5Iy2tIRlG+E6
RAiVcQy86nbXnwdIHKpUa0pVMLpkPF10SOujACXV/aK1TgZHPFTLxPry775WzN7R
4WshMTHa8cH0m0C6GMAaJFeRpfHtEchWNYU5PSyhuFkxnKIAljvJ6+czXihBwCBH
ykfEPyIliMEVcwcbCHA8phOHwMWUcenjOM3ecbwwSiCIzayQobupBgCzBYjEa++u
vQkklYfoXvgXluAQvzD7Cw+it66LpQEttlrsa8EIPA5pZsdRHlUjp+8Eg85lW90x
5ik7Jsi+hwDo6sPxoE2xNbyHem8Zyyur7llG6tHBnn4drkXMwa0sXFwsVdPHO5A5
hsTbvGwrMjSJQFo3cG5KfxH3K6H7xd5LnfGJ6WI9vyPlei9x7tmw+/MvVQfZbQgh
vkClNRGXE+SxkGLPZ3RMhuwfxp60pJiSLhvrM3oi2heJNf6pR9dTMVSbONmRiqmi
4e0ZfSt3V8NxEalaAnws272trc273qBGSv6WiKD7e6Qh2/Fo+i5f1Ha15D1xxx6S
pLFLjvzuC24Zziwzlcl7iJdHfp+WXOkphCjXl5oWaXgBtyfKy/4TjKg5oK+dMfKk
9tLvzxGHPU8QoT+QSLtyt5+4xg6wiH04vYYur0zDz0XpXBQ+ZvUT8YEb4+UGK2B9
KLtwsnD1R5xYfL5GA1vT8qM8ICgMgRQdoLKG/22gz//lhYBaJiUm0DZixyB64OC6
HQ7btSrizfk8huhl5qWZEoWStbNi7nSjIn8JfQ2HEPiqmHEn+Bw/WzLWVjDGvn3Y
kkrt3Ih7se9pnp0DSssBVGe4dzsS5I97sUen7g5WN2ySKXcvZkHcfzgK6YhdDLAI
drjc5UhPRRmWmWkAZlCRx145MZ9xzF4on8HQv5Uzavx+Maz7Qx+F7COPpaSQCta5
gEZ+mD5koIf1PU+TXe8OtGtMPLwTaVomW1O7xJFNoXA6/jDkqFdfrefG3Kv194Mg
ryDVuzhnGbRz7VzOqLl/uuReu2dJuYPB25Tidify80WvpNCd1l219wDZS0wcrJLe
ErGv1nzBOTLesYc9j+OpkFUBmLuR0bDD7KXQXTmLEQvE8BB6vmhPyGlUfO0oXYcz
h+pnI0blCHwRR2qFYlRbXpVw4agFh/2hT9WgEfPG1xvqBU1Cb8yRuZJB/e0dYN85
pNXxQaq0PYhOzfQWSoeTa9yq+8t5IroPzFrpE+oHHREcHLTqNTvEuNAk4WD2Jrkx
UEg3NxcwzEokl/Z6gAncMG8ipyPDQfUiOFrIO9ltK07PSlJwRxTWLzEkTl7eXXXs
z9bZng11oznL4KRXPh4T4mTl9deLHPNvH4h3ExeUivmCDhUKYrjKEYPeqfJxYunX
t63K8vf1oGz0OF/+xjrwROqlimFusoKFKZmvOd10nB1juRAfBOD6RXCZXnfbL+Xh
fCaBwWV+NDJFXEWcfe1eEQ+T8vOl6A2RZZhucqzubLG4C0YoBQ7oLbOAN16U6S5g
0S5z0B5xWLnMDessFMADViEFyFyUhpVXO1UEpEsTFso8FCpaKK+1KUS1tDu5RVKI
4BZjHDtR+2pOcSASLhPpptSg2GehTV6kg2OwM6HtiL921LF53vwXGW5L2/3e9HDf
0JJ3kXWqUjTollqDd8eqjHCfKrUiMHmvYHwqBiRrrTXZbF1HxEbyHAplizDEN2pH
v6RNfPnmRAyMGzEV8bdXJsq8plE/qH2jw7+BFEDiYhs92d4YhNfdUMMEKYTcvc3a
CoJmmYUq3RlHgq8iysPfnLVlLpK356V5TuP4gjqCh26DazOriKCFDo/vUHX6eJGL
o8CZVJgS50S1s/X7ZE5GxUaQOu9L/7ZFqa0ybsFS54bNXFmb8yj5QiZb0pV7PWZK
CyEy91ny7sP0s9qd6sU51RWBK8eDuYVjJGXnRYWcMvR4fOGSSji9pnhnPpJPBkmh
pKHHVsTxVCUpQJIBDSmXKhoaH+jZX/RfaAc460og6f9nmz9u5j+9lmdzCUtWdsK9
Nb/veb7dMejdjkkGPDfhd1NxPn0WLpFUwzK/s5zaBvoMk6oZY4bwrzx6T5fYIIpU
pkbMym5GQGeFt5pM+Cqow4WlLuXlDXGn8I7oIo4LlHwVQBlRE6l47rsTPyrCZ11x
nP0uvzZH8ERzFRy+XW5a3GAMW+HMUJysVbBgrn0jN/WB7Em9vlYdZuwR8olXPynQ
jd1tgXr61Gnbj6IvCxHlv2RnQi8446qqMz/NvXOfxQTdEbB0C4OXy3LoyWK7+r11
xEi2u1DuGhQ29Eom8UxVeNeGokqG4J3fCvsQM6Ylg3DUiRlfSOgQRmhTN2hGmFfH
luC5tAblI5XuuNwre7Vn65rC3kMUVxqu5Hoih7DxuoTzNklqMAw9RMxGOi+FV/x8
xFVFYxNn1X+8m6p44ByIWtQYSFTliwg2yvn2g5eRD0jlNMQ1PK4NIony5yfLq9ir
BIZT+EPhrxmMHM0Z5j5/4VkvuE/gedODGsPTPC/jhWOUM5k8LeYG+2EEq7wAMa+w
OHVCY/wx9PnesrqMRT/yiE4QwTplSZE8fkSEZQnIfwBH/YQkbqAZt3KYj2I2RhKy
2OeYBFY9bd46beC2o6B9+AHeAd3H0xQke63vyRbjB4S+ylctKpaQJaqrShcwi+B6
HigGOewol2YC/qosJ+Y7ZDZDG2aYW3lOyE4yp7mGsbg=
`pragma protect end_protected
