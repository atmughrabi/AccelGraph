// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GrB5QXKHmr9BZZGxC1lyqua6JdNw5PiqBcbbAVXHgB/arLTVewqsxqt0ycvMLjTp
X23AtBflmSazZElYEdr4iXtxSbWWzlVATDrmvJ9qoMYDOnE9ek6enobax2mAei7s
k+HcwADSsYcUJ0A2XmHiaBgjxAZ69d6AimT+lSSlDJQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8464)
jqb/5Dhci/4r8y/XiEJvVYhnzuruDuZkHbDNbdgm9ttvxc1l/R4t0a0sav8aVPXx
ZFo6m9EhGni5+EHJD+oqbbxafN7eusHlw69WTQ9/+kwPT7sZc1EqeB94v8J4Njy+
qPEioVizPOw83jE7i1gcCctUZpzMXesXPbGMCktxPC0FPzUK81EIni+J7Kc9+pQb
+iqreQTdXs9o48vE5IDaORPRRzTOJwC+gc7JyW+7uqGOd7/Dfsb7y/DqnHhn/acd
wrPwQ0fEq2zeHTdCbZetz8WpILCE+1lZqi/NkljgnfOrqk/5y0zBAEHtTXUu435y
n9qvSDT8HxThXpCeexv+SHAzfErHZBZYer0Lz3Ed7SW/xbviW4AfGC89+SlnIIfn
EmH9sUu3IWe9DVM+ydb/6Y23qA/0lUa27dm0EeBUiCi96N2hfXtJpX2HA2R/4Bmh
7KhADH9A/Cg+uiOIAn62Z7I8JuJTR6wlkhKO5FpDRg8Rd+5nH8aeG+7TlIFi3EpB
0bSBKZNbBZQ5AGgXit0wOedseFzVIjKKqC4BirhlyegxwZOO9fPQh8ddttlTtJH3
osEKl3ph7BUQTf9rrxPITubbANSR8b3eZgvI5/3OKlLHYPeHufPbnxgJXlsMeqn0
wl4KNHsTSErOxCQLP2OMYadaEJXoKF4vVlCDBkGI//Vfll6cMy5M/kqXF9M1e5R/
sRprX87z3NFMoEtIQT8FOccp0UCFazy1PBY9n3nV/qTl1eGhchcH3qp1LZZEfA37
TxraxuBUG/ENtf2EjtHgy+3EXAtRWC/2Qp8MlP7wkd7jRLuLC1mRoFZ7i7691kYk
kV6Ei4i0v42v1hMin6NTLHMk9Zna5Kd+TA4ghDrUoDnwWMF7W+9SEZd5YaFrwWZP
/S+/KrxqDfbFWAblGNd55dudMrBFAJoxrB6eCnN5Z4am+Xn4KrHsliN5QeGJMBnw
ZMbMRLb98ovdTmtezRmJxCcjMl9mtxpkwg9FRAvlc6y4OxVRPg9rhMbrrGBqpr9A
JFLYBequn7ZzWbXCI0AKjJki9Npk2rRD8tYE6hBWyZZp788FSVA6E6Mnx9rZRnjq
PDOYbNl0aSPpHDMYnLjw20hELG+COlTkOYYd1z76nFDNqgwEbpPsiqumbJY/Y/5n
DRRq+dtJy2SqeDhFJSHeBzg4upTsrl46l0O9nSLsMY6e0LDPJ/6v/r8eG3YflgWB
Qt3LTBRWdCYXzH83DftRQ2nvQbj6WH74ym4pkoY+hCeUKNwzMFPsOE6ncalyX8pM
CBwF2W8B/1ekwOb5JIOQr7DTh1oKZtufA3JdUNS7k9RmeEIm4ztpabM4NJddDb7v
QfgQGnZvths7ldu3TEfjgHHDGgmNMVj5gNHqcvgLwEXFmXNUH9P4WXq1vWRpQbW9
SZ9C6L8XQRUXLzDwJd2aj4+qwzOw3g/1imm/aDbIbdTI6JeSTDqCjJzHjlKFfsOH
xdvfccHQk/NQMnZQSvMj5CBVnWxbBRGPCPcNL6TMIjUSqR2m3LjP3APqwLq8AJBm
MUC5FKKlJ0/rGhCdUc3yEHC/yVWvtgGt787Z0pgNNTxtesSVVMEVIdvBqDbF7mMD
WN5ZAdnSCO6zLgECnQXN2FFWOJfZlXUHNHI6H4E+xVjkfRYT9I8gTXGhv1WsasQm
kuPuyz6HaEoc0Nb2QrypValDdmu0NuMAYX22I9SDcd9/lV2/aKBBqcgPD2FaL+Du
14mUBAY4UmAXvCOEw48gx7ptSUYJrNoqBoRS7lf23Inx9xI0gkZVBeW8jHmWfvrN
XNBeCd7aFeUREmpkeGJsvGRClfe3/sYBHAWaSS3U+XMgFHXt86I33IF2NSsTmFiQ
ubq9CHya/Lr0nduxtna/lXZqrfHO6HW46oubM8QWHhXTknue6/8jlGyHcy/fZv/5
5t9H+Q9RX14jiQpWjJqzfCDK9QrpU1AdnG7v/T9YwgP2KD0k21a0JynwKAtfc6aC
uCrocZlg+L/3CYaf+sqxNrskfVIjO314H82SeZWd1Zavz8YIha+dHsVSbvruY9xw
hJKDn28YonpoXWL8fEH1XJkOO8J/CJkgTskFGnHAdAnmqGNkypAAS3Ab4M858Msj
O4H5T3udS67kV8QEjUOt1k8HSJMrRkl0rafeoepJpnKoJfunVrF6ZJErZia+a4vt
rYFJsNccJn1NBr3fresBhvdk836gwwkMNfhn6vz+gydYCDbmbHCDsPpW6mFv/viI
hzCgNJXLjchC6fHcWoUZPfT1wZGV6r5a5Uxq33nsUJMJXzhkJW3544RWFXAOds47
NuYq7tJHnX9pfcPoyke59MRkPjtp+vbLHqk+qYNCipSxWWvdk/B3Sqfe2rR/5D2u
qPfT8EtR23s0dMcX4MMLe0LAaQFJ/FdHvDkWRwJpGBjQXfKHY76yOAMW6JQ9lgKI
1yrWoF8Vmp3tw3rQoOAlsrpDz3MHSpYiDV8YSfPIh1/HQcvvasI2Sa2kirWevmvx
5Q9ICXJXUFsxJUgKaiqaXhjkr5bG3uY8IQGtZ4xUjwbK2I6hOEClDpeMnCqZRr2d
kPG2G5dDl6/Qr8lJjpJ3tY9/sXpdNAuNk+rQ1ysSMAp43CnQaqUvg0PvgUTIBXuI
i7Ov9KuPqrJnkioxYDmWSA+U18S5O+1bjxorWFpB/umERJ2YjzipuQdHs5FNpQK2
/0mp1XIXTIbavsSYQW8aJN4mdeVSf515RY9R3FfawjGEBvnoGbpuTOeD7DqJGk0Y
0oRr+3LLtk0UdWpNcLyRj4l4Gvdi6qEVDWXz5qTVgjsbo973wC/C/7yVGte23aUF
s8OIo1AIevwicTajBxAV1WxtaLUfI0OcaDzBleDo1CQ9MR+9fsXQbeKHIFI4/qQE
ZGU4DICwoYb56S+qO/EFhviAstQ/UfAAs6IF5hI6jFvwEy2/zoGlx+e3AW9TmCIv
SXUHJ+eN/ixW5mVKKJntCMMsSjv0HFbLZ1AD6I+jMFmMM5CwW0k7TRlBcgWtohy1
k9A6cseV3f0dhzLDwvjrGPpx4BiVdiW+zZoOLRg6/f0LAC9VFZDDGa0YyoYbQsUD
xZnsqg0gjyim0n9TnrjMkvA/M9C0YrblEtk21aAp4Af4GlKO2RfSG5FVy6rXiIaR
FTUoOFPVTzKKrqEz/72mhrddEKacYO4uvbZbz2hBLEQB9hH0CxyFwa11PSI1aGX+
+hXHQW/1m/YXa4J5w9e9OjN+bJwjVOz8o+dFv7l6XotHfHk7QtmCUtp0jP9vUXkU
OAzJqdux7TU8Hs1bW9r30ht3JQif/TJtKa9rFqcS2XL6iGpspM/5J9z6FSdc8Vbo
G+Zi0It7zRJRdfC/qHOmbQTAXLWtAUtnwpAJnEnqS12ETwyr70szU6+8OQWk9ush
Y6YCVCD9LPaemjkjsPa7EUn4XiXI/aGrPnndli1RrzY7YkdAbVCXacBPvWSGa6h5
Sh8c4xqm8eeFXdq7j6bNGX6A0rF/v3d0AlbDHCoPjRUeZw0MLJ17vLpnshpqPxSY
4f5csMnggyJ5itatPURcuwvw2ruFXfICa90eEaHFS9IhQZDPBE/Vw8jidR1+A1B4
XYXO9WRIyJv7x4lgJOBI5qJdeFhjlUanFV8zeIqIOn17RH82UrrLJ+uDJsazoybz
zs+IsUPaI8SXRylam2T8276EI3KSeTCWVDYtwR1ZTALPRoeTcFmNmG6WXPVJjyCn
6RItC9lpewAI9x1gXOePk+9R/nu236xvDfuLp2LyGSV6rx9PCcgOh9GjYTG6kVeF
1WuzJwiusWbGBVX5ZF3cDLJBmw/tZQIZSoH7T+Nt0cS789rYb4c8jcG55pc9LqFj
bBzjJA+63CwgajgfdO4rxQL435nCVGwU+tJqSxLfjDzeu+YBljlBxjaVcMCIbG4z
4wuoFIv4X4XpNLQLVTLjiNbfxo59mkLlFRE0ofBnV0/R2Inl7zJieMJINlhxTJsF
QW9lSmOkIy+vBZclHyeLaYAyu2hCsONlAVBYrmqU3843EJoettaALHJ6J8CNjkR7
fgtMI23WDrkNWmkoHMaE/uG9ljBm51c/S3zv+7SGYspeCJ5fh5VXZBLqolCQRR6x
Bi17ramKjNiPBygpCtUEff8kb5XkElRSRS5I+JE39Pgw1zItJH/lfsdtoVbdsYNF
PA4/JD9xc0zy+QFBiog+qSEWBUT2LhyI41j80QE8zDC/CkH7QkCKnFBCedUEjFj+
FJa+EhJnHFF8cNTlJw6pADzabSWjsKBK8AjSs7myRlNarQm0P4+fJp3dF/1cTAuC
Q9GLnzJuJ8iNaIZR6XJrGI5KRhjDsv5Gtj9mU14GdUpVW0QxGgqCZb8zDtttw3rj
c7Kv218qC5GC1R1xOrCeqr0o/3EqVXsokLKjsca1RqvgMoXddsJ/CxP1Z+r5tBK2
lQYiwIXmCFNnOMBytaUTm5sh6qFHLMKi5MZoxCGPibbMx3aWm8LogqBSBlj9mZd1
gRqB6mNuGPoZ5PKp44XbBiXXX+DzzLznwo8WjGMruemX4sXhXiVVVthzQlVmxAvW
dOp4RuDvaCX+mvOE2+8IvY99vXOf6csJ9uUFtzJbLTOsZKcws3ETb+7vbZLxYdZp
i8xNUL3ZclbNvb96SjCa14/vgINe0gRYWBE28JcJ2ybX988eRd5zQBTEVepKZc0c
LH0/8a8fyZeZUGWBRK6b/fmMl0XbUIBIdhZFjTKcsjKNkb9CsVooZNHjOVV/ciDK
AvwL0DyCihh8ZVXsAfQ7aaCjiXdTY3ch1nRptmfZpX385fMi3J7/dDIJ/aVmxl0b
5LfeWessCq5ZofajcVaTgXcRSHGc/yc7o0uPSACZb5B/etyBG7OAQOqAs98qgk6Q
6kBFa/WM6G7u05+k5wGinaIzx5/7ZjV7mNYJ13RAjJRmadhTHJTHC3/vXpzbVGpB
uJfNiw1V4ZXzxYN30q8EIWZACrcccX6Nbzo3h/3/22QllzWXdcaZ4LIqUKp4OanB
rTDYqsc/GkDCvZCdel1AfGj8XLUSRVQ4FNhoGrZE/hIqrh6UZzQo14eIAYR0nH6X
gQNVNSVhfbI0lh2m1h+iHY5SyzbGGRMQfAnfwkwJx2xI580t0Mkz9tt8fDoAfluU
GrNZPLXG02k4tGka0XBZocHK4IsXFqwQQqK/ca18z649fkRj7m0m6887XAubpJIZ
V7WDh9Vy4oEmhVNEj0KCxHcwhPH+kQYsfOiW/UHsP5JvgpOspzunLYscf/XZQjRK
iJeMWyG/yKhNLMyIod7SwVdjNaGMJnWRDZ9Hts7+AsNZa83fTYqCLJj1WQlrljM5
FqE6XuKXSTnF91idvVSR7I4rG0tfOqdC+fokTw1NxT46bZv7N6d94Jrwc059rbBZ
UECsAjWdvB+LGJj0+OR5K0u996zqVOq/Lbqmup5VbUyGmSS+iNJvU9MDSXdGn0Su
nn1C153Y8SdagDow1h1BN1IqKm3iydyKk8hEMicBCk30+ZYznAfQVYpaUW9QH+5s
m0eInRtZ1er0iKEz96CbEkfMBJILg7EEED45QvUmEXejYuwSPg8VqlAnvdI26iNh
IQiEV6ytaK7NAz5DkwUmSOzew8flLxclpe7Ij1Ef9UVR7gIIOIrk91Wg58byzJ3Y
Rjo0YX6gGc/UND12yEYCIdgHEgdbY1strqkne//2l1LYh34dY4Smw/inEwp4mM5Z
+MYt8xA2CMQBBspw6B6hquM+23ppRSd39dZ6Pab6LHbfUD9lmp8rtZ6yogHiGueZ
pFzY3/gUPbAE/BEntjwLvSAqYGpH11YDV2kbfMwIz11lSgs5IWyuPdzb1tqFHxJl
XiHhK0ojGEfIGiM3wSRq+b45AUEbiGdYt+WXhrILP802S6xqnfM0NI3ZJ8UVRo4h
5XXr0rXF3nylZDIQ3sCJ+cSbDmSx1FK39wEFYWRHwwlnSYZObJv+dlv8BLvn5nJk
0JDWIVuWloacmOwHb569mmvZRW2cENL/hDQVOXaDHrt6xMBjgaMW8UcvhbH1SgdU
mmCkqbOKslAURadurmf6dOWs6tf4rwrdzdoTRxYeqN33RMJTt3Nz5QcQ5RhbdvV8
7MMbWhQXOMgZXts6B8KfDcqeDd8c7zK0PaxdF5TvJW5FxPKmC5+4gfCHPybQnkXv
bbFT3WWH9nZSoAEu9O2fcSBWEGDFrwKgKtrzPzypuUW2PiX91Ln5HzrIzXAtL1Dd
KVNVIV5WaXOkhn4vv2B0TNDIOHrQTjE7OHnUBSGmtuBKb4srBCAAtWdr0Gp1IhXR
BL2a2xrmk+57bb06T3FRyYwzM1X55L5GSA4r7H9pZHb/nuO3SrcOMVhFBpFzlRXb
2EcO8CXtDneHgkpLkAoCP9tW1IpfnHrmZXIivNL8Gqc4ZShf2vOrXfyWW++ViA/f
Z43dWlXkRAUvSvKuYqVKAOtg+QRHa1nZyVlaE0INO4L2741fQvfg5HLuwmQHdsGL
0XXczAqUHm/kfDjO6dWA98gokqyrIYOl2VViGfxgjoxdGgjNrq17n6KCSEqAniJ7
INds7ofeeaxcOzZj2GernjgJcubGhS9k+bTALSLl4Yx1eLt4n5gxa2FUCt07fhuk
rePLITWA/V6UKLHrRMu/KV8HnVjWUcb/CU506ecavASX3dCLNAWGe8rWD97aMKN3
1npn+kgV1TdlJoGha/xHND5qKkn5bGrVPlCGmpikzP4BEPD72ji4QI/6BMlUGK+E
1GAgAk4xJzsSh37/LRRMUcByH/llv1uQ8y9S4Ym0rF7/aAGYYXewdy8zoKI2uAho
Pwr1IB0k0n6yXBURaFDX1aVlIikfFmrII27IeL7udoT8vXtWW51BnJZ2kx4gLpqC
Q9E9ecmAv4sQHKBgHTLUKKbAOjSv/fCvXKyNAv/Ad7yHvTuSqfdQy3jIsg1ZRVA/
gPO6i4p3RMZStpNKgjfLb9M0pSvf9TiaR4szRSJwSm1ojrM1DohxwBPY7MTB6qvu
X7NX6aD71zVHN8lcoeYgppmpnk9csC4Sf+yMfpFRDTFV9G5CUJe36hY9tayzCf2Y
qhD+eA1pOH93CpmvVRfLSacXzkAJ/HFuZxTJI1nllMaB13TIRhxXp4cF0dpHPlft
3rbd1zOiykcGgSXe92FLlvSJSbiN0A9UkoR4RSEBk6TkyJRA+uNv9ThqveTl7Asf
Il1EzbtKtiJgpo6lWhp6yi+5v5beuH49Eliqwk5+VOQUSjNYHV3ohnq1cFMzXefl
WHPcbTunAUkHT9RlpidDw9WuQjoqx046qtLzbg9YiGqgnFx2OnOg5YbUDDmJnR4o
fICCmMh5EEKpO1kHTSIwZB5PSrCKcSTw95lVChIxvL5sf4VEmBkcMeP7gsUmVOGB
PqznbZw8l0KHSfwmDXV1aYFZgrYDJTJV1a5PiB9gpVw15A8CdfA0U2yKyl6IyxP5
0cjguDPuqQ34K93mFMB9xm5h0y3yxKMkmFkKDsKPMYWpOxrP93QEicX0fLjp+CCg
ouE4jV2sChj/mIDHTORgC48UO5i92T78jelvkRtTfuo5RGVkqrkhRqLXQkwiUBTb
yRuV+cq5WuNzyV6IZsDuWd9YkKCaSSf1ley2qOO4gh3YM/uFamwbiGYrXvE8NYKy
vxc2u3ovqlRP2c0kl2zIvVLmCS95VkuTQ9d6fRmw2WmXP2ZPly8L6Y9E6vz70guw
nk+ETr2hBQUhnBfUkeZ33+PaMxcOjfSDzoFGbivfNyG57m08SZg9K1JIJdcNG8iq
7w6plc2sNGX8TsNni2sIb55BxHPwYAhaAmTA0G/aIhfAfu+IuVcS+X1Xxxu9IYfP
YM916T2s200cmKWvvsyYEjbYtxuya2luPGk+3m7OPof+Lanjh/j5j8Ap+p5T/52x
s59nzOiV8xEpcZgaheA8le0qXGJNzgMmIu6sG68uvVkPY79+Hou9dtGNdacN5rkJ
OlGJs6aOd0kwOMDFWsJQU6bdFb9mi4vs8ib2us6IweDw0H25UcGiq7kWP0e/YPX3
vPWstUMHjUj4Dy4KrWaW+hotqtFngpeOfIAql/cVDLmqixS3VIqb4xGm09fddZt8
6rPkW8w5ui6esBfDExld60BygNLsrfsS8MAnYKvJ5owil/284cIETLV9qpc+BxaE
pghvslXiGAYLsE4wDyZEQVOWSH0aY1OI8rysO0r4oPOKg4m0O7VHiI9IU/62uFuV
JMnGDyDwCyIUNs4kewRR4yMfNDu59DOdI5v0yw1Q0T2wzR3D9eUbMfC/M2gy8YfR
x1PX99GVhgOJqblmVFBA+2gSlhXxo0vFMUW9L2DpOzt8HWpdAFHdzqRGE2pJEpwR
2yUCu+3RC+L2+G39NGuU5Cezr0wUm8at1SPHKQ7JLiuuqwuiV/UXQ2b7B4Q2DjXj
WN/acuigzGLFBBx08lzlgJo982y+E3dR8hG+NDujzWO+eux4Xj0KCSeBd+MMdSLB
dZdkwIg4r54L87O6Pk+3549z7HP+xE+B6gMZK4Gv2di7xb4GkRO20Kzw30uMi5H3
RrMNWCZJL/WrcG2/dgcUCynd5tkaLNn1R7oW1Jfp5sZeo1uabyozkXcIQ9dVRDR5
U4fBhxBxJODWzawC9k0yidzc0yPA1RkrlwJmbCd5pb6QyxYNJe8yO1IoYlT8h7HO
/qphlbPEOaMX3wWnywB4/o2tMR5h96zzrhAcj2k21p/mxoSkNFcmrG9NwjtCEt4W
uU3a6W3Y+3yUCeJVrE1BYhYn3Uct8V+YUoWYUUCan+zc+EEEbVciJrneiDHvnK1+
4/r3ek62XFHoi7Vs2xSCu7Ocd7juWwZfnFN1cQJAzqRmzOcFGNRgyfe56zlsrJak
xSkmWzv0ujULngdB9L26q2NcTRewX32HzSmfTsk5HGVMc3UvlDv8YBSH40/Ns1D5
0fZkOMlfFgKFBZin2Gvq2yy8q32+P0I7p5EWs5qDHpP/WXykIyr04yV8v4DzK4nI
sAHHslTmgmGaLSVDvYiFHF19Z/lASPi0ulMTzvCGWCJ9vPYTvaJNHcyQCFV45M0s
7DcZC6J1R1lW4blswf/wq+m/BDZVu620u9o+SSYtl/vrQSOpxAWZRsqDl14JtTP3
catRvRfo8R94Z5vi9OUSgJgbADy2U5Fk5k05GwkRFma+C5gTwyydTOLcuIkwXPRn
lCHu5iCHGkqallp/NXb5KM3KUW/UAM6FpsRDovKnJTXNqBGxXR5LdbDDL//bg62u
3CZeecKQxmjrG/sGrDTawqfy9iCJNqt0AldQxRdksxuCVYtDpT9bzqNuRHoKm3WT
4TwqFBUY8GxTlVKRvKwnVJknYncjewszZhCgNjv/e8r/klaEpVExO+c1xtdIWhvh
6u1R8SEBDeLf/IRATynepOxmBrAe/Uc4mvFX6RoaLhvVY5rExBkKzbc30OG+rlXG
JXSNnPRmhG+5+AjmkZBqmTjHQgaVvMeMvBEitJ5XiXxCaaTa6tiKFcQ4naE3vD4A
tOXdY8UqMDJqedMwU/qwKwPxUMdM7KA6Lc1WZuO8CT7Ztsk4G2RCyGiQ2cOltIc7
bdzLAIY7LgAr5HBEWVfC0Fx/0vfmeJKYiMuzF+ty5mYSorSDbHUxjH7R2gI3STdR
iMJyjEv9+ofWATiGB879TNWRxGfd6mLMqPy2MAI0NDqGCpUvVEEE9ue6XV3lani9
nIdVxaw0hBqpmPpetlpL6MLq+9ST7pei1xTSLXqQAroz7qwVkw7IEBDRLphfUiSZ
FxxOuvv0tP9IzBzJboTJQnJI48mqmAxImnIh9UJE5wg0mmduBRivkfGY9uctr9fl
PLPpQGM4plxSw+rtp1Fwn79I6dRx44hETOEoBuUpCPcfnlQ8Tx/LVCs6v6S3HB30
8IktWwsiTf/GmloYAaHLiaWk7LOgKXGY8Rg5r9iP7hhKosMhKvtcCJXrp7Quy8zK
o47SySV2xF/8dbgQeZrdy1GkediO0hS0irKUcyqgW0ndqldjtNzbUo3CTDqF1ya9
zmv7mBMnd0t4utGwHq9iSuMuB9XJzotaY9tHCeYkvGxR40z7DB6KRffZMxm44pbj
cniyDAyKsUSYMQzd469+/PULvQWMrmyejp7dvKjXLUccM45NDLco8GlAaEUhkBFn
SiPcUzt/eNG2mygHSwqBg4yF6c9CtfGaenoeem6BOKwEd8DP3w0otlQk/L2xFOPC
s0NL6ZKeGj2/KopbCysBiKw1olGD65GlfekHxwI1gFVO8YqGNlIgTW73LZVMqzfl
uiWyYKEWrIM6Ct2SvNWDrZt3ynwEPicHN68TJfsvmTE3Pzy0x9ETEYlcij6PtvgH
8diR57zjpdB0nyhsHvJL/y9bdST3zp60Za6hHN7LeaR264vzFkojDGttxiU4464V
Cb3JSmKzgy0BFbacBR6coUnS1q17/OB00/rY2TyZ6BOzkLLhXtOoebI6nBoushZS
Z6XhUx886hKdT1rvETK+aF2MqsOfvxXJJEm6Xezxjsm4MLQ+Pfj7XTWFLQ/eJ0Ls
tdfCxY8YKU4ZyOh2e9ikj1dXyRS4c6+LEHZkGDrlK1TJr9c2y3o8xwXdagVdK6Gq
DlorXRUGta/Bypdev0/FWXujB2kAgrnuwqCrAhF9YDJ9+e3icUWCnaPK3yEheYbr
Qr/gfjpNqkz0oXxp3dNFqK8sV2FJsBbACGii4QdwumYBwlj/Be8lIn2hUHV9TgGl
PGUnFDIGsoFpuf3V01YtTPwXWk5MmEPgcF0ikubl5DuVCFRw53Ly0UI1W/Eydhg/
I7juhvDTEPbkF/1jlaAHGjfxUiBBjh9EQhY0SSxhyCLDPClfJL+ASFp5TuZ+o+Nw
AJHj3S63gq5xUXU+aq8y+O1fBxbrnwixB/6Dc036YUBo6mhpfzdb4IXlXxvJ/1PD
G8XyjWEGOrKUeOeMFGp2LraBGm8vnwlMgJNMHJyaj6HE59qMe37+N+LxbCpyfMK1
nb3rsUht2+CvI5P5gxstJZSK9gIU2i8/vqzK7e9Dqy9GRCRAzJCuM29H8dr6JiCE
pOwIS7kN+lCP7lPtz81JGCwfadwczvYTuWP275kF54dC6BIt3kMUkJVwJW5e0lba
NvoZyNRXjS52oLgkG907pTd8URXilAls5nyk+mKYOV4/NgWk1e1PZmxqiKpucYKl
VGojEDlV8PvYgP3ZbOpRWrA3DrZFl4ldSh3PlGXR//P2PvFCwiQm72TnH2/7OfxH
YRZE6aLnpcCJg5JBF/e1WSa/XjMGofeG0l1sy9Ih+wEOd8iEmdMTzp501IlfuxYS
JdHmqXOc6gFHP8IOHfExbg==
`pragma protect end_protected
