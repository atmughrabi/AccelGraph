// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RS1lz7mdd3NwjOdnyFm6CBbvmyrcY41gLA31TD8psK/i7AiTny+jUrdtqXyc78Dg
aE4pT/vePUk09ihrHrvz7YBMGI+v3nGcZoYUh2ejb8HTHAJHErm8Oo7vtey+FOuG
7rdCHe7zzwJnHgpVEos4d5cWaTPkfPZKzCiFgcTY70A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29216)
xBWiWlGPkmxGrI3IB7+5wDMZi5RVLpTzcdMr+rIeypg9KdAscn5HYaIkmWSBB4IE
+kgg+CtIPv5J4fwLjrGDbA35CJthGHxxjVKse8e1gXHUUvOBKRyY/ypXvbf77zFC
qKmBwzuZAArZr2LF6ZilI8yF3PNHJ+JuKry9zMT//1QRP5kVEmQWvXxmBi4U6SJh
cLvYtJ9NKdgXoNcTU2dPJsMjAfYGheJJbrB44zFU4UV3xqERpQNrLbkGsK/xh1/O
8FIbLMrMBijYQ+oefW0DxvzKTgITZ3A2BjjeMcHsdHeONTj4d3BJmnSfrlG3/FYf
KdC35dl7vpCEeCBQh971nYfPrcimbyGxpB+Z/MPi3E1egv87Iu/1CHwbKh1UTtGl
32Z/SDU+KDxBOIRuf+vsH9fIMQBolf+uf2KeZh21LOzkB7m0r9MOtBCevIdGR006
d9PTaRKyVz+xS2yTh2qjOxFJZNC+axju9TB+4EpEYEt7BW/BaVG8pIw71BiGiIih
lb6yZ1PD+bSDXbMmQEUQbyCwEkCqHQw+c+4Qqjm7a3ixIGSX8rZCo6/LiWpOwkas
MMhQyqZe7TxLEdSqVlVCTPkGExN04DSAnV2tiH2oy1GHvpIA8YuRvoV++qLt9GnD
AsY9ndy7ETaQk21EAuazQqnZ2ZQ1PPEmyeEYuBkGTobRXqDv2B3yblQ89dk7BMAo
LA74v8XBglDRZxXGv5KSuGJ2PMHFWjOnAzUoISP1Sbfy5UlErqOpMTOD2B2xJuk9
63mKb12tUug1ue4nFfTSC0UVfkxEpj2FYO/lQgMLhyyqTr1B++sN30UHO+RpAb2W
ih7dlaxDQv0jy/kU6a0Z7yrYSJK2pPtovRDh4pVRtAp9SRNO+KSBNHy4+kw96+D9
ON6ogwcLZM1Rsfml4hwzc/dKSKI2KGRunOQGZJe7w7ZnLPmadq2LTz11c77sklk3
IelA3zTlbyp6t7fG4dCUldnL1ao8He1gFZiZ6R53G4UgKtRTem2+8mArvSriQMQN
MDbk9oBq62fJ7/dTFgFZ7v30e+LSjDk3Px8+X3nuL0+KiyBfIrX8fBGvImaAlK2q
OGYWN189/VgP0FI57/WSkxDDmh1jki5v22EWoHERo4WDd5zfai2shGvdrbid33TH
LibwhN9V8VHaVa72IbN/4iMy626eiBkCGT1r5VJPNCMcBb2VTnfWlbhTk3aSXAGm
KeQwCbUbkIQ8iLAOjftG3JjItOH+yvqvq2IB1rLtljpwoLgedpWODpHlX7C86a4X
quvqp5PKW8hmncdLkrDAIAueKpWtITkedjYPLJjn/WVyxr+8seK+BmF8YF5XOBMj
6JqTgUVASwbAyg0RkfqhrYydX4kwAOoUruSddpP0mMOFf+opN1T06bCzVcwbug0j
0tNi9b4MRmj5wZw5PsfCH/ZCHPJR6QhwqXZml58XHKOs5vdOpl2Jjb+FWc7yhDUM
CGQi4S9IOtOSGFdHrcFR1gp2s+VNrL9efPzh8GcoEUCa89zwlEvuHT0pJnOsGoel
4Kp1aV9EBQylIFSmb/oxKwiq9d4I3VhLyRwCXv1l8q1BbbDP09KiH+cQz1JOnr5x
sN6J33JTi6t0KYKG52FKzjpZ2qKgieQ31NfNBskTzV9xy4gKyGu3aXBw0xmT3HhH
I6LsOMJu1moEMT+g/X8K3QuFUJk4R9LM5pgK43suy9OauNJA5/tYmlSvlW28CG6c
jKE0uuKvFD8Cv5q0q+9yXooYURn+Vg0zoEY/1+3rVgmUUDRRhw6+LSjAoW8xjLK7
GnvzRz76tDnxlo7Q4rt4Rdo085DzqtCh9jpyiYtcbnwwn1iBf5iZFc01hdhGKoPf
7CiKIJzIDWGTofdUMx7aNWwoneJyHMtEeTtBsQBbqfUbOeK2TiPqQruKMA4cGtDQ
n0cTE27MyvoZoEe6ANXXdU06rxHGeXHr/TLymeuwkC2PRcNTHLBmuH+fybyrctxW
DRn7nBKIG0kYFWeDSKRBjSkoKvvF/WiRq0/uCTE3FrS9R21rgi4rGZBu2/ZcNC99
TM41pE8Y2wPrk7J44RpqhVnizDQR26YZvXDGZd5fbKKr9psIDCxhgMoqqzv/IHsP
m72D0t4p25EuIZ1gra5p9Z9m8JEN3DvEaViLGjaFkpjO69wvQ26J8iUPfAjZjqQq
41tRP8cFznx4Mht+kG3nm4o2rY+V0lq1UGsEo8zKDYg8T3qEhALFpxJHiH4qL+hh
u+41aBi7VAx/W171eb4DK8TNLMz4gc8LCPcgx1c6VPR2jEkYwpDIYT1YznHfZc9s
/Nl141dfcrjdNl3FywYDebY/BLqxvoKl9zyagw5B2LWPZBL5kCkgb9mMTezMqY+H
40dyh4TfJNR35dZb4o0KRppzzC6YHWL4gfnMWdJNOXU+XrQn+HoDuXN2bW7Fm5xx
kR/aNpoI1e1/N22ufDaw+yig0mATrh2/uWmbi+yrcJHQe4KYt+RQgyI8ikAENuWd
Z75sd4A2y/9/Vzkc4i6F/hITIkMxDuo50mHCeHRnPij8kmEYwTW+6qmy4LZFRr5T
9KMrGwbnKzN5E14NvvLGRGVAC8w4GLurd2Iz4/iLEQ0WeWNJrmBBvgvL7Oz8EjG0
Lk5+wKTWBpdnLYRm5yb/qr6nWg+GvduRDiIZkgRDChXVSY7bZOofnGVbrUi2yqXl
wuu+FYBooKBqB7vX/o5KhRhOsE9bAIWw8MyxuAgcVq2ZFPVAcnEVDxMhTaOkIwFH
qQZetnKbKltmr3lSoSypyPcZxUMG+kXhIQpcIXQkkgUiS9717iCsuzRq0KZR9DMF
DRaMLiKw1rQ+aO7uNeQI3DHC6b8NF5Zu5Y7g08uE76R4h6ddhQagayjXyRrNzc3p
OaH0n4RE+U2QG6L2upBSeslcEvl5GJ81OzvzvS7QFIcyPmtEReD9EG/FeBnICX7T
XyTBMBJHKTI85DaLiIPoIZVtelypU63t0+fJQsbzEuXxZUGFj8ko2D8cZww+pv+/
jsmEazcPgitFxv9bhSc5itex5gY2/7dCqZS1G9m7xvRn0K+JpCGF4njUiPDvv3Kz
khWUiLzFPQiEM0A+lHdPGZcuqrpY+FiCIF1npryElXaTahKjhW3FyywAmfGwyVOq
DVt31aPDc1q/v4bcosjVjvrhkpkB+8eOEMfjoT+c0y7x31oeaWPttVdpq8qi3Ars
Fn56y77m/1qB6Xtgt6HnJQAFH4R0d8O+0RA2xptt1D/CirtXc9dptcdFZnD/g+ZT
8buHQwKvjSYyuht50oVJJLtuWowrBgU0aVbruL/7GcV6G4K0PkuETiMzQ/Bsfwr0
Dig9839iru17iOhG6PGBlVprP9XBtV9DlNsUkGo0H8E+IrvaM8Q6I9tI0bkc2jFF
PIX37HcM67P/8GXdc7HGR7MnIO8D4rD4/nJilF/Bb6/l4H30FXe5wGr4GkgauQcu
49WG13zEOwZ/gm9k8u4f/RnEt0H5ThzF0p5EgsQjyoNOA8Vek9iW1svqatFNqnhb
IQuBZyjCvZ0dfdeI8/7TTzHJWaZY9g9VYT/teiwNr3mFYNDPMBlUExjfIhQncc4P
+wkAgWqPYKl4P2R6QKBYcZ1cGjjSiVQSFp31B10CL9KzD46bgdVJOR93AFqhfRlJ
fxM9hKNXndXTDqtQmtTwtZZFITXXCqGFWWnGTUsRXHzMWpim4+LNKm4SOCw8lX3S
uGfMiejZdSgu3vvvljMgRcNAaN/M4liZ7Z2ShBKsVz0xeGSMOlUfXEf7bEejyBKF
eA8TMlUGieuehId1dRRZthfYL9SmFjXfR0VMwoj0mFBuRCeRvqHlWLwNlOWgzEKE
Re4nhKItLNwe8stgq6NXjLqVp6CCDNKLHBgyt042qp41QvxKk74gS+RaxwZYuEQV
c/P4s4Bj60JQx7ulVKSEHPsZ9UMrgz5ufv6KilZAkRJ9F1nwqjho+3HpEF2WSbIm
GwD/kU4OBAaJeyFZByoLUPKlI28nqR3PgZrU+ir53XRoaW/uOwlV+vpXzrQlPyjk
DT4kUORvzQXQd1zaNTf8ro1+LyBZ2PhvcPOuOr2JCtECDcNJLPRugmqLav9nBPzE
ZIReLvbDXWVJHzG8/xLR+iaR3pk9DwEBbYUyXENw4Rw1Y/gdbpyVIYYfOSuvGmfA
xH91ULrpTGefwcfjyUQQ3CHzB9kq3zUPBaSlC/ChTszLxuI+/OQV0AC34C+8I4pc
fdWfejVFd6CPzvRE9xbusSaJZW1UYgeTUSFnZESbYjEa1fDlvYVVvTjCUU+JN+rm
y/b6+fqV2R/sU6Xtj0Lsl0hxdNmpxPHC1VInehAZxBnMoCwj9aOzvz1947FYqgwE
LDK+KmxSHZEQ5zDDORgiWvZW8NWaatuRJU6s6aRfFjl+Xd6/IgvTIzIylYwy+Jte
Iw5BLobmc9nK1MlIk85P/8mZXY/84VDDwpKID8JM9GLcAxmygY4xJGE3hlRIqIYu
gqVRyeaQoyQ099OtYo+F+73xIVVAtnJa9E8maSOzzO3WZYF8ff9uOC2TvWhy+PPl
VfsVGh4EgywUp/GB11ckwXnmaDGKud78SLx6NjVyxYfEnTm+d8Q4zETBhRlW0reV
NBwX2dXSIzF25BObPJCGiGejOl4/ushJ+QIlb+byOlppPGdyyRQIujJAR5P8TSCU
U1+DaJh+MsfPuH9iP30HKiRyZjEf0uV5s1jAQQ3UPFjamAsaVbFbMTE1CXK6YJmo
rHueIAJnxdI8RqKFPmYlu3uk25V+plWOPKqbp81qGo9/LhBAd63TBU/cFtBTLZGB
p6JfdNlDIVi0fMqQ5yeLSQXYhGTbQ8Vi0xcnmEaK8hfCC9bEQl4HB9WXYeTyaedn
L22vpcljOURbsAW0YgIBo2YoWAlQyCMer/64+IpXSwjYnp3QBp6ow0UvZJXS/caw
ffVPIqhw/xYLt2k541SY+wp3BhyfreGFL+vTuwQ0C1Mz0ESgkLxZPh+XTI3Uxcg+
+CCqEkzOkZNUqxQ9IHbvobTsTA6XdVZ+CglFYk23uRReTrTGaaHbgt8ufsYKumQo
Gg0tCG6VPqWGvNNK6kCSUWXKYqLstdUcBexfIIE9fRWitNRebK8R0hER5hcSKJJz
hmrvcyenaeiRhyUu5QeoLJ+EbXRBJNdC8gHutIi3pZw0s690K15xiLD2J5gsFi2v
HmbYxJvp/csS+wvaZyzpbAvU701amJdlK1QNw7ahZqNwnZwzhEgcCXoUD86HWCci
s7kbBYcLrTsVxfSRNyKmc1UGNbbVkm2kewU2UO8euMsVDMEfFXKQ14I+6UA2d5gX
efpiS+x8N/adgz9Avf6gFhM6iE9gBdnv2rYtxwmzTEEg6J9rhEl948DTD9qhoaYy
XNO2sgT+8COGT6uz7XVysYKnXAY59NH3CcJETJPNjXzj6rrPxoUpStNIzzt6S1W5
33yTjEjY2XSrcqx/rFKCfhAVwC+lpJ4k+LojYNBOlZfvO9Ek+1weGHUeR+XfBv0J
lDrHpGYXDbJ0LrsewH7lC+P4nLuOlX1OT2AZYTQD1zh3pWm1Vt3gM9W3c42rW3uz
mxvCH2A38tx20ZlRupgmvSCIqELi60ED+8/rjmkpxlVZf46yEwcTxLPSk/2LfU0r
vR2ah+DFr1RmGINlWXr5J6NnZjROT/0KlPhVJPzPPg8+Reh8mkfnrtESA8BtKz2W
SShOXguQuBOW34Iz+QHJ7uPHs4+vGnS9i4ts7vv+1upw/eDkj/L0pNV08wAGPtIO
fACTxxR24XnpUqOXW2uvxi+uNOuwHVml2QD/eeQjK5fk7thixDMdpnGshaDxk7Fu
0YNvdSEKbPIqZJJy+VD14Ys6gK8+8vXwpl+DC0zMMI3A1uGUYdOcaxe4a0uBaIRj
hHXd+AXPAGr7aiHQ7XzNnU9x0/AsSR4FMvjr9tOwJG5xsCm6wfUEXzbUrFXl3nwN
qXJZPceU2S0HFpv9U8gC53QPVtmCGZkw5bYHW7Y8Ttq8wOnUMfXdoL8HtxPOCfaJ
xHVtuk/wXxEA7S8X28NO6s09PN31QGWWmJEuRKxa87beE22MzCUJ2XqBjb22z5QE
ReI9ZvdoFlTuUReZYI/68FYh+TuoL5p2YcBXm1aYD6K6ogAF7WkvCpsjN90swUAy
MsKnYTUYZ81VXjYmIJ2HMmes1u4uhlmYB5KR5vWVmme7Zfm4NY4wgIkul5jkAhkB
wA1zOvsT9PeR8h8ru+/utZSAEC2jeOzC0IgpTSmV2Xwe4zH0xP8PnS2GohpHuFXn
XDUn3Nf+wQPNTZVKV/tSFfj1npEzF2lmcgfE2y5OrOA6a/Ii/z0zytHGNwPXn6KM
bh3T/GAp0pPdptjVNqhMlPkOhYLt8kMITFiSvjbJct3GS8uH8EsUYM55JxUmAAqm
aorJslNFPtwBhnMqLyOVmWF5w3XdBk/gUsx/PZfDhMoiwWmqmymE7P83uBoLmbaG
x7igRbvfLRJSWmhFmy/DST4eTb3qYJXMpAmdP6DKTNMxg1baQ8RZbm3CyCRrtHsp
J6gt3msh9DBEgQRsexovL5c1lcXJxP2PTP7c6T0RwiZw7v9mI8JMIEUZc/3fp1o4
lRFqhpjZ1tILpxgsxL2gBmQRnXClzto96/VQuCFigZ+z1tzo7ELkYk8wHwvfQThr
SE0/Vs/0JRge+QWqsNl4BS8zFuV+rHaE0oQVBj29wkocQu8QeaTXoCoP6gpkW6Zk
+fVFcsLVwGqi3Wg3W/REaiTglInQGYk4w316Ilg/rd0in4iOP5iQehLlExqec5os
Rygz6URsN6aCW9rQstLQZtkz2Z1cTri/n0aQmdpgC/3gC4pq9mEROXHNr0Wg5Vai
oCiotkiCFdOecc69qY2Igb8op9Cs87Za7JWIdELgJbk2DNKQMx/NqN8zpqtE6bly
NzaCDaU+DVN0ibKo2Xsu0IGHfg2/vGkF6YMtSsbJ2Do4UHFuSP2qXLc3dD4oB1YY
S0Oc+9qjFt0vOA6xodBP4fBTCf1SWUyst+hjpmctB66K3wFWec+89GtNZt3D+GnC
RjGFGSOhw3Wlv/gscDGcXgyzy1D/Pzs/J2+q2AXW9DVNLXFtsipcFli93vmtL9K2
rvzoyEJc3mbN5+GeVvIMrkFvc8I6aGDvR5ecjg28BbI870y1ApdffbFJGTvD8PiR
4d1BfTz+kWrzs1eLAouni6Gs+w7cq9MGG2R/OA8ZZ5YMC8KbO40d1gQlZPhmSvVu
AmaR7MVYXCxBUTkIXPcF2gnPJXsNBXk3a2uwNT79CqAh4/wcFhj1pSQOH6m/YGGC
t97nWQ68mtFQYoS1u+IHEd2jc5mGflI20PAidM/uC3JN7WEh0rAmeqCaiM5PBNfQ
D+J1EOOy8P8xTKeqMMWmmtxzxSfNW9GE2Yw6vmDtThu1VDZZClMObVHEA5bMmAr/
/KH1XYm5RsKbcd2cxgJf34bfq5n6v81UM4bzZ59C5PC6gWhZ2TRotUDaYA9cTcPj
yTN+ukGWWmuSOWyVjAo6mZMM6/7fncSWznQMZ7lu/9KWz1TjbE1Ku1h/zxawLsxv
eP/l1YllSQmEUDFO+qLCMfLLqkAKBlLwLoWqPF4UQpAfW5e1b1aC0aM/vDD+x9J4
27kPnR8BA+Dj9sSr7lTY2fiBBm/1kKbTKie+uduEkNqIsL43eISmBsDqk5TokGAF
O/f1aKhntxPnV0IJnPYPbxcNNE2xTkjgP1Bmcsl2wQN8rub9FtSQQQLS7nAMixGe
6wX9zFKP0UCJRpqMhCNl90y2TLcVob35H9sv//NbG36zGCYis5Ad2igMZsfi80r+
O3JtMGHS1/+ilVQx3I3bQWDjt1YvBJFNX9t8fDdTdk9Xmg0KjBcNQtR6aHUjTs4T
aFecb09UCw3JWCSqmL4iv6J6ZEF1Dj+2PQ6BN2JU+0tfN1FZr0D9wx2x7FA4f9/s
SC36TwZZBZHcF3M+wN34QV5EY19q5ChhknuMxwz/CitE2kPkMEqWiRuY0fC/mnRs
t0bjZm0wNDr7X0voM6OhGd9Q8G+ucaKMm5ndJZCkkyUKcnTiIALIXRbQWaav91Hn
j5uLGAYFuBOeHBYmAiql7HwiDxv+nKarAYT2Dj8yWjuV2uhUKYW2VTn4JVbnYsHB
oOtcwRf3IbuATzeW7CuWquMyQeh6U+aHXmkyuJJMftBCS4NeRDM8Hdp/clBwcgm3
0o8uiLIBJHOYbttmsF9OQS4Dj5hrgAvNHEcVOKqIyCVEtjjw0sWtEy9yhQ3uMa0q
obWXBuuM1YLgCq8ES+p24vtTRkf6FjeB4m9FaRijz1ab68MMAroX+6ytPsG6Ra72
q1bsXG42hPzMoQZ/xINPiC50k7EjVZAKcJrfaUhtt0RouovzVOljYFE/3GDEHLiG
M4xBsZTuCTSX+QSi2uqmh+kXi9Q+uLyfah7FtxPUkn9L0WWRJ8/4H37NeylSxq55
xjY4dy2zu9/ulx72M8YlCC8uTGHAiVwJAavLHIH4jLw+Pq32Zu7ixAM/9XyE16ad
3z1Wypv6rhcfP43X+pSFgkWMwGw8iSmml7Wb15JxpFxw3vwhbtJbkDRm9k3K5m2L
ULUjcDKR/I1UL4srWeGmuAzWoQIzm4+XriDEhl3LQLPXrq0/fB7Vjy7QbdS1pubZ
44xrluA++MbjhH5knWoKNqQztxKCIFcRjahYP7c3tRiQVTFmQAXzJbgY3AJ6JrJZ
/kKzfy+0qQuIlTPbP8FMbEen1SnHKwJkak7aQCa1X4xqBDPxT7qwJsJyQMCLGdDX
I3o1FlYrT1z2PlYk9CRQ2M+YiZyqs+V1qpjSg1CPlyn1TWhNaMcEhuDcbKMz68IQ
Hu/rL1n/6ai4zn/DGuwy9bxfGkXoQfBaERwQOXiu8zOOpCj6/B7NiV4WopzRELp0
YUM3XAhjqqrcCh6dZGKdISK6TmJlV71mh2UjEMCHhewqHxiHe7063luyYkJh2Wqy
RWlqajgj6xE9ds7K3hV+x0mhH7W//jczwPFcyEb+8Zz9czkg/e8yrbHvFoNwTtXR
kQ3ODkccQhV+0ErXH9uGfjDnwckUnlABxVmuOGPrvTffQHM9JcZeNhqcIG6a8AbV
SefrKkduDHE8b9adaa3lzDWuff4SjeNDgzGswmf23ScmWAul6HImV2IL8HzQ4rNz
sUdk3T9+5+u8GRJ6PLcVKmMGkI4KgVb64JJn/twVEl5KDNQTMLgscFn1eRcrFk0B
HDz8VJq3bWObYLpokhBppVtFVwpTK7/Qgcg4d5OK0rMLzybLcaM/SJATsoPjhdgu
WapTtTrregL8QjEC1ZHUgYTOlmTLZXTos/NJNinkvMGEVhfoYxEOvmYGRiwtrhBT
8+BVV1tkrT7Yfm33sd/oD6YNEPA030YywdSr3HvaA6KJjpXH+nLxizN+rSc3529T
d9diou5Gpb0DVoWRxImNCjLn3tLomSQP7eyrjTiyP4hP0RgwMiCeLeSD3u8egs9f
GTUywpUmAPUjn4l+jeSe3Pjcbwdyr4SX66sGNh+3Q6i6xhMreMyg6roWQ5O5mKhc
frbZYJQEMut7tmWVLrOauWMNtthb7z1d7xXeDqu1qpxX2ekUuyXg3WgLWgWyYSA4
2zrFiYj5JBwpiEnuv7QnghjvTMyBN5GOwSp2a8d8vTs+hBU5vVoJHtKZxHws7oFL
1lnVxYprOpIZlgqz59GjBDnm1BiPK8pTF6Q/vYltpm7wQZtirrGOy6FMLBgb7oxn
tf1dbg8WuAUNHNjayd/KNfbm32dTIq9ShXCo7idBgZzyLQEeoudA0d+1im3r0XQV
YKrbbYlEx17dFq7vY4NoXNFEgf58kJnMd+5uV07+ADtLnAIt5E+pd7pZ1/DTp9lS
5D2wEP9kuw0dVIB+h2BOmVb/NZJp9u8luqwFf3vGODYhVgJIJnu126dGV7yOoGkH
6BLNkH52z47BLt4YsJ9x/joWRb1njzO9n91i+3nGxU0vlF/4WFu7xI3jUSKGVN+x
xA8mr76RDC+pKW/dC8H+A39AxnSngWWBA2sAGPeMK77i10Q9af34JIIBtcAvWT+M
M2+h6rfvS2657SxpF/DsMMgnLSO8tw4As3Puhtf4xTwqv/Ks5/mD2RImCRQypFwo
aZXuKr9g3WlPPMb3esESUNi3RGae19Vy00Z+7Zmdns2/vFA9hB4+c2bhw4oCeJn2
WXHfEMwIc2CFYV7u7hmQseBv3xVMTEDupIDg2exSKGL876iCCJhVOhRe+1uacmuh
kbJAMIhKOuVJnzL7pJC3eN0jmgfg3cm8GelN/Qz3mcTKnQTlBADOl7MU1EfGkEq1
AmFstINMgFDBw5+yGdKCDNf6VKs+oThEbE40j53kdnWL0XAXHwez3fLHdF2MVRKJ
nAC3EKmtqRQfnsP/xG6EI8eP8GTyqeCJ6isVk5nZA2lJthdD0/2BDojl5qWA/Dnn
j4rQuAguEM9wSHgqjN9VQ9QKj7Vu+f4buBZ/NIbHEnDhW+Z3qmBj4Z9OOSejqsL0
dD6amR876KHbRJW4mm9UN7q8nNR+RC/znh+mUH86AX0yn0IPr08zzd9ij/p48YGY
1zNEARGPxPXnopXauCIwlpbHE8RIZRPmaRn/+QoeddbllKih0VTfi0Qg1NeUvKAJ
Loq8f0t2gKOHpFWxM/1sg5cGXdn9AkORlKU1VxVdEBPIqJ9aYb6YJ/GK0tNUIdGt
ujXM3uPAp2CaDXmrfJQPADZAOBNQcBk2Qd0sA5IkifUBT6tPOBSuCR/N9GFHTF6x
43hx62NTbNtQijjdoj8likgNDOeTOjHdbpJCFX4J4WxNDIBeUprh0xtkh/AfCdS1
gjxGbVJYX8brY/Z9OP5JKdEBKKPvPxZeBKUv1cC7UWA9aSa3JpSvz2BYif7w+PLq
YymQTOKBDJM9EwP+iEcqxllSPQJmaH2uuOwKTWhBjxNLWj1N4m16aDindfsL/Z1z
axnX3VzqtAVfmnX1rpna+4YKGLQJGczbEel+TJIii80jF9lomH0aLDcRt6mdsSb0
FJ9PIdb1UAYmcYDbifYPWXltFQ3nfOJnb+NEaNFi5shsl3Nx9pDUKazjmaGn/sHv
lvEqR7CCh+WqgySM6hkZ0wGiIxpxkcBD7eQY/6gF3ipxjEEm7xn4LL4H0bog7QpC
jTfBJw2v2drxZPygRF1nWG5C1HPpW/s8K53L1gH4wAgZjIMsLlZ9nh3cqf2Mppwx
fDoJdHNTwBf5X8xrdWE3+Exp0GsXsLWHScfbNbCbk8Nv0ebv+pw4GPfGiOatvldO
Ga3nHWvr5rGAxhkTClny76LKTGla6IB547m6yG8JjsrbM06mDiH3cAgs0jh7IaC1
nj0qyidey77+P+4fb56SdGHC9vzfgiUnegWyGzrOUp8WHv7tD4Yttflen5PyQGci
PU7PNrgbDCTHyjfr98XUY6QtgohPkHv6mMEdqpTC02StZ6RFD9wzcQUnnSDbudFJ
PamiV1sf/JA8H+nDiryiOC481GNyK5grn0D+gzLNXLEearWRFNrRiSXyBEV+SK7x
Ge338hpXZAEtdWOdmJ1BOlcVSeZlk3DWbK73RRx+Iv/bbD4reSn5ZhY2u82RO39c
Hoz2looCrsGL3NArcVCS3vrLoRMslRtuaiKOU4+ks0Y5JLJhuuN1b9iLjZjWT7U0
ob4pJCNK5CuK2OoTh4Nky75//OlQkTBTip1wCA+tkDEQ+goicWU31qEg00hwIqB9
MZ5R9w5IaNG9FsUBrWNRx26ut3he4HH25F/QkhFnOa3ZzwHEFOXpXBW3HUbFLJIh
DBNKDJ0fns8BmEQrCD/oCgnz83rZ3iaBip6mP2Z/XLR4qpvzbqRQDtTU1PXFev7G
2wDfuePCX6/E62eLwHXSBLi6OViQCZE287hRf5PJq9zNFZvkKiyvHqIXqZDuEyJ7
u1n4S0LT4L+69P33zalnKG5E/7Se2WoiUaYY5/yXygxOBC//Gd22SeO2jRTeJve/
VcM+iblANecH7gZhJqh8tPVetkI8tCyoc+Uyzz0dL4NoBKAkjqymhSIeJja//RB5
KFOP4M5IwP66M8tc2QUJeM3JO7xYDXYV4Z7lMBFMSRyqWBueaRPzqRLuAwRLxkCJ
zqLXp/dzADvsqXVxJ+otQPB4EDqpjHXHSWHuSr9N2iBzDGMRUm5RdRaHsqKsdLeb
G9m1LDYTjovFjd2A+sTxSj0MIXbVIfC2yHWPeC0G7+20acH4xbZdywX9gUyqQ/I8
Pg0fgCfbMt/kEzOCOvPfH04ug4rIAXeNzsKOjlhZTa2GisMkg4dw0o6pHfzMFl5d
zSz2ZF8cokxZMoG/SavAit24+J753D510FPRYXnjrgiWd7pyRgaNPCffLW4OlTEP
oWpR7Bgt3HM2/sdHxBojfQ0sMPNt1vVfz1rOZ0Zwnvo2Zna8cCrOQ8h27sO95OVL
oJasNgUdsftIPgUaavnv2hZOBRsOG5om3lCMx9LFjbc1eiwmviVx1fcXsTRDDmbZ
KHSBm4YpEHnP236hvwy2Ui9jLoCWbyoAJR50qP4T6Qh7UMR6JgwrJcNdP50ot/Mi
9KHIYIivxJgTtScVqfUW8ygvpWZxM0fTfZ3AsdAL1yHfqrES7rKxi2G/3H0nSYwN
w9wjQart8gL27FuUlLGnsVkCA0l1HH1d1jm+56yGeTQOMBpqvJx5qmJ0V4IjA/Fu
qq2/ZxfHak/LMdYioHdqSXvqEE7a456nP+XKxuwPG9eyzcEa9lo+9XVi21nZUhCy
Vo+ET2lN08Zyk1AdcHExQQALXdQIrA4wuO9FazQJqRQ8yPwG7WCevLR1gCM7kioU
z7zBbKYJ37RHYDA7NapHQaJK+Pk/087YIwkRmtC/eecwQOGWe3/DfI0lHZ/gPI2n
pTtnMTkY/jNZHqWMQxCndemZ3RKL95nN1TCAoUijV13UtIU74ZwAnNyM3QICljfT
fBkl0e2+nTmjlBQYz82NQKuKwobsdgr9uJBxI64jwL0ao3xpXknGizPFsFYTnFn+
TbsUfR1tbU4dwzgEdSmN1sXhYuVdpHv2X+TbR9x4R2NI8f2Wr2Bfzqdi+GUZRSZu
+BdrOEA55Jizby2Us8CHIEt/pyNIYAUYSNLC7tX7Q24UV17g/BdhH4Rgyai8zMwI
CuKCqcPyXL64dKYTEDsJa6U8vuG9nrybRimXcGXYKjZ2SHtIA6cWMS65R4a5/1PC
748XWuarZDUiGVNEpwbt0fCZQn+83ulwtjjw2ONETThSMKtkkI03ozBpkFwzn/Yb
q4agU1ePHKduure9z70LYBJiHXx/XJZwllsy8MwLENXsdcb7K1o4LkVcZ6VyWnM4
kGvH1Naladvh9GN6C+mi1jP2uewym88su9sQjJbAp+nnBED4Hrg5R5emgOg3ZHb2
9B9Y5UGT2hOSwwnXZAXtbBgGUPTEP1wDr7lvJzDRISnzVzfbHAvMnjxaTPFdEiP2
jKJc9dkGiSItdkdFNQp07mkoZE3HsxUy8DYqDih567YdygQpRfIzHUbIzyyk9+P0
R+4PeDuCeVxa/domFg5dKakrSTIowETDEsgvkeHXf7BRvRrxH0D24V2jwtXapJsX
dd7n/KJwgE5VbtK5OaH78aKE53YSVhnLcwm+KIzsml8B+OhZzKCJPFz/LLXrRFRO
ctyEzMy9dLdsuWMPo9midZ3YgSlO4/J08rNgde1csMLxt+zxPi+iReG3wG900nZH
zeyYG5FpkA/logZfP2r/CnOySFS9RIaWIU8MTK3kdunPcqdu4ZMATcjH0KQVI6kY
gb2JoyxQ8ziYJbmJ0zpfaudRJpRYBv9KbNaYIPgZZei6dkn2yOZYLFu2GeaW3Dts
J7E4stvkGIHHSz39MaxmSc0Mz94c3yf8Az5/cdpihLCpf2nm6LxXPrVr8yeys9dd
hv9PHBGfr1t1jbXYOev2m0VqGH6QBk/nu5JopAhVDOoIm5NTECFihDAkzPisYl07
KD0Q3Y6Bcq+9NR54HZEnEHRbLCQWmmPWnGvf+QwkWk6tHE/TFDi6UbRdpRaIW+Cf
Rp5GePD9seLhLqWIliSbxFUNO8dQtlewwZBPVtKfan4WNfo7L16ayKhA6ZLnrd3s
bGBS0yO71TF9qd/zsAR5Yfxk7LBjEoIZxFv+plIxP4HI5hLxKzUEG2JH4DhM3fqT
+52RdVrzgaVfWTzrL1hpwRGwv3AkLRrcUtvPN3iIztFLd4+VyxxpkiQ2M1blZko2
VECSQUKb1IkI5od1pTw07tTPCT7/GC0sFCMVlFvMZZqwFkpyL+Pmg6/GszS0DBjJ
WCSr+yttL/mtGNCtci0DodENyP2I/EiO+QbhGmDLn5LRzfObgvTp0mLj+BsP/njF
tiYygEecz809toTDMiFdn93IDR/bM/GTw1rh7A5qkC7z36xG2fN/8Wjwz6dVrtxO
M1E2bq/eQKLRnmkQaNTxAcRY5MGSykObgNUdajWMtsMRYHpBTN8c76AwkVX0njTS
C0EQTPudG/CFypW+FkK1yqIC21DWCk7aq4cMlnEck6L1cc+mXtnBTAa7u2aQal83
ppmhWklRarpN/F75lwA9tix+RdZkbJCj/TkupisLLdjEzcMO40roNKW1WJjRsS6c
yhktuvRHayHZOeG4ywN1l+arLObUfpEOcDsNDvxZjn7jonBE5W8EGhQsKt7UI+ky
oVxGvZ0QEdUKMHwwGrCYiUeY5WqolLvjOsUaS1PDVtr1t4sDBgrbXQTSjPT5lkcZ
LiXh7JMBTtSE+B1pu99xQGVcHTq9TEDPx6OJqVkbpU41qylvY4h3/0XuJ/7ToMBQ
X75oI6sg+VtAps26Sm0y9FSwqa7x8rOr0gKFvCw2WsyTn9qt1/Qyz5g/KB/kfxfl
ARZtlkb9ATE8PyF8IDX6SZ8bJ9qICXKVdZSYC7P93QcNVf7bgSAx7r+T99J/nECV
mYsRTn4YfInINri0ES99pc9/S9UuUWLGsIwtNUg/PeTga+edvgMU3RY/jGnZFwr/
kmbcIfWwk/Bex1lnhhT6UDkHBohZohH1hDu2qVURTt9rE3luABj/KMWAhHkjTK65
5ZLdDc359hF+kLs4/UXEqklXobZIQQBUH86i8/n8ikD+Po2WAqZeL/CxZaz4NRB2
1xLAW2OKD28RasA5XLqsWTfNbtEcRF6L6YKGNpOht+sFTF+qcy3AeguH2+PaQXL5
QiGflf/cztJ/L0zXWEKBaMZhEOmCpeGvewV18Cescq00KGXMzklwG5ZSZwUTSR8Y
Pqo/xuXpfTS3Cyb4rAdBMSMJRQpPjf3bqVEmwt5rVGChV04c/gPz3f1pwd00ibAB
YOnZbGhLOz8DKjDyLQQ5oA1TLx22rXkTDTMyNvKiOPxpmKOJGCDgJ0KlrN6/U1pC
JvOBh34uWOCT3mR8AHWjLItX2tliVhUlCKWVQYgdVJa8BNvIHIt4V3z/pApv0tx7
/XlvFlYOJx4yMjDBvs91E4M7IHauBoAPdcxa4LhMuQnIWMK286psbdHH++AP4AOu
DLs9dnvTyxDRcMRLgmbYbEU+/zHrttj/jPJJhv7hwRaOtoIP4BouQiCGg2hHrnL5
nHeaBcrgu+x/s9tZVnXYWQ+VVWiiiyLlWv5oTyxItcozLmnOubsOco4kRgCsf/Yl
8hJBPp21fz6/iKqnGxHJBGJN3Yu+afoY95vcC+Bjvab462hfnZZdXqdgtWdhs/An
cFzbH4VYtoMh4i9zy+umSfAduqSSCsilTthpfESl7z/69jDLWNUxdhW5okEtJcHu
O+4kEFJon+iHNxTtEifPMaQgBrRlBWKujIcrZmj21bRgKAVrsbHqKfjaszR2dy4g
vytwUfHneAR1M9jzPST19CI7ZYzzReoETNcaOtQ2rXQOJgvO+mClMSX78sJBuL8K
Yev6jLjWZEWxMJojDSsGvOR+AKnAPfINA+CD9KpbyEXfPEYmcV8N1ASyC04i/yi8
QSShCsmGs5i8fZslCqVcqERXyJ/yoRZxWYbx/yJeF0xb4pp+QpPjLd0LGZrov0O7
LjsYZZrWac8Rb5PZDf+ar84dcW2N5Va6b9zZJ5snr2vergPxewsWp7uz0O97pPAF
urysqxtxYkdcFaECdtTQpA15h4D10aXuswADCRTDjq/UlglhmmseFxqMRlUOSlqp
M52GJ8kVAriD8LFdVpx1VN8HFMgm5pSoliP1MAK8OrSiUDydaNOmcemwg68bWllU
hXb5qmstoIEoy5UdZU6lgkp/GW8wIP6bvawFaMntxGu9vGpcvuOmewo5qJlN5TWY
JC4KVSpu7i9OgBfktZ/ho5Q2a/9zcY37ZgFvQff9ceNUMDZdRPbeV0Bcp7C5aINB
sDCax89gZuSLm+l9nCbnwdkWplK/rijziyT2JWwZJ6x3PwbkLPHDBgLeMwiEAA/1
pO1tnJPeUuuZk1FFC51tOR90wspTzJZ5CzmvmO6m2vjNWmUUIxQIZcRAudaUbbxy
t/XcJOFW1k+G0CYdup5/xV4LEEACzKVcsuwTnSYnehVEBB7lL6prGwSJkn+ha8GE
oOJg2rCKAymFsX8eAWWVPfvxSHGEHi7KIyqEmws0x0OZrwmyGqckupaQreeUBHxj
dw2eAX+2WFhuj3ziaa/wWzZB2U+KImyUpTqP/8aptKq4oQjha6adJ9UDK9lKPy1v
Jpa4A/Tglnp7rJ94klEqKQddNCZqm+plvvjOIzjGUSrww5IR6vWfOPU2LbEKUld0
t7gRmKuB6GQAsz9FFX6RwfkgvOe8+bLMvJliU9AiV9KOha/nw6sOiUo9B+G+xuO5
Q9QqL9oRex/NrslttdAcJyoAMzE5otvUJtTkjac9p1JpNrAjM4a1htIf7dSWKr8e
pwiiW10efxJvzo3BwoujwiyxKFmXy/0AhogU41mAyFj43lVQNL7PdLRl6YQE0kd/
o8fmTef81C6zewtL9llFx/FSXButaYeBvOjqBBzrzvgAy9claDo6lByIRV9xbsv/
7m4DFlBPtgHwHvL//WNtXZN++VHNUuaMpAHkYXaCjLtK2fliYtRTiwtL/q5Iu5B9
meS8OnjE/a3BooKC/C1OiuxacDrkSw8djn44d36i4vhT4uo8MJfYjhAKGJKgj/dq
SwQxyOs6VBXXt9xAlLBiAPft5BQegf0XDe6reKSaXDj8bE67E/A2ZyOgn1yWElGA
tNBw0uyHXczqyZwJW0zSCvl/Z0HWfkcxNPdgEg8TRUBr7h71mmMYYMCn9RvNzb65
3eEtfq1cyqWldNmoLKmZdVsKFL6sk+SKb1D+jDR3YerILazy4pMWw6K3H+B6MSc7
jTcGMOWbfTXU1BMg6p65Gzs/8UYSsUbWDXpreytXEXHSH1pkE5HKS4aSnZiwPSsm
ufT+Kb7XolY3FPjQdZJ0xRVrilKUVKNXpE+gdJuTMP6B/uGkoU1yBkAcJu7FqBQg
whYZ7JZUy8Gs8l5jEjvcAmqVlJhpiBJNZYFneYfOlMXpOHpqlJ+BxzXwTBEdiARa
q/DK2qC1n4Rzmv2rwv94QuWC7ZIbvimNZsX2TsMPl5ywnS30tgQh1DjMichV7uCk
OzRfPlHaUTSDreBdT8jQPOx5UOdqCQYqOKLMQ0BaSP8uKYd11TTbqbTaYASOuiU1
UupMj67gYQ25QlKDs4jVjbouYuMPIafbJU56pDA38KO6zO/7hgClGWePy6h9puLR
yh+qXva1/72t3yCbD/onfYo5X1BTZXsJpQ31SgkiZdA98VkpLQsyOiRoQYfpMapf
0xyC7WTsCErXMk1+zBQRRZlAhOcM6RZlRIKNS3xc4SsOGK0dw86Yz94xUpwNjKHy
NRj4+GijpwO4t2Z9rMRBjJPKh2L6PmODdfyujtz3+nZPkm2hqgei+fv0EdK6PkWr
H3u44S8fJbiH4LmmDGAnahHgqZvVPmZTBmBzvRFqAWiMaDK5GIJGN0R4WN3VA0OK
JKdAusXbJgyIvbSiQ02cuAVlwavnlWUV3/ey2UXW4RcLxUVIAylMt84Mvf4f7AWj
L8kB0qz3Z9DaiJzMOkCccu6VlIsmdiP+VXY63k1zV91qsXkmrH7lJ/zCtudFvfY2
z3aS33KI42eZCpPL0Xs2Qp6vg+pTjVfrJvZHlxuainZzkJZeQ9K/60Kl4mv/bOvM
8eNJ+15I4DRmNWl8oRIWyGj69GWcRc/6tucGBRt0wtVbMoOz1Wid34Wn+642r7Kb
wKBOe9mWRw3kFmFp79cdGUjLT3pdD1CSpDHEHHpUzaxAiGUYosNCnIpCw1mAZwJv
3ieAluTpHeuPNLceAsbBXlGavzZobYZFNbi8I7USvTqaqWJEFvJ2wdbb5w2w/fqD
mVlyLsOXZZ9Xzl3oRUP5sgp1e5eF3uPeZkqYbbpwxTNuKdWLo1GTRtAalHaetUhF
WCx8CYOWKHu4jtwPjH9LNoy5R+p9V8hvtKd9KWaFUtyCLHF620LY+bYXRzhjvR1E
ZGlDBED8F1Nf8NlprSdqq93uuJJGB6D5kP4BVK1ba5U3q25hmp0cSHUA/b/9RI1s
tDL7UHySqhuGLcPAN6t3A7GaE7RbaTBmUblxTNEcFOS8FsRzvmk50OckP+wn7vdx
Xya/4kdU2vip+oJcJSeLeQpOijsJE4q7ljboWTenL8F+688Rvn1CY5tp9OSpthez
W+hsHGVb84OMeaxWs5fvlQE0asUTCnkfdqbJMfvlKCQscfuD7IelO5KfN56/VxcO
ly5wfL4Vrmq3zZ36m0hOc6VPgiQXcxhSBUhQFNs5F15QUQUo0AkJ79Cu6+owKSxu
xhvee0GXRLL+BlKZl/07CwnOcswNgKfB+NWZQVHzPlCV9GxOqVMoQsxFWmTHz1PE
bEU10kjNqgJkPjHCKXj95LtUD29tI+/aYI6Tt9qmrTSdON+m6fljrDcaMqfSSMvd
tO7ymomMtzK4gGGzYCuXP3NyIucSl1m2H7PUPnOIjrxUSbJpq4y2mzuBr5dbwnOS
a5uMZ8gMLJwsbAag8lQGgc2ZeXNf6O0JzWBo+IGxSMwkuzjLWu91LiNz1plvcYP2
S30PO2gFlfaeGXnsH0bvi+GPmx+gVwzaLmoUBqRVjkGpl8l5UHTxA5Lx3p6Tldwo
ApjnhGXzWTBeTDie25P8SnEAONJ/UKnvLMDZ9smZdM19YdV78wKDIHRZhXaGEzG5
XLXzzr0kQ7sTq55734Qx8zYGeEPcDXIsHrlcAYNcmoB+EeUQw7H7Yj91UuBQpNeC
FouUUlfUbuWdEMIKURGJ+VgI6cxIWNwT4/umGUCENWIDlxPDL5YReSOlKNZjx+x3
sosfyNeKldg2Kt9w7ULRoqOowwnmW2RqHPDFUOlAUg8emJa9oyX+N8cC7+wvPmqP
yqjguKl+llw2vR3nVFV37dO5z2XlK+ALxMs+640zx6nZTSTWj27jZtDJpW2MHoGC
yvWh49KB48cwR5zNbMB6FIzFYHE70xWSWeiG98usMIe2I4Rj/QQin6hZ09nzlHCL
2O8r0qI74QnHV3emkf35aV3hOGNlCFUv0vOQuV3RWGiIzoaErsbUuAnKt6nOMaki
TffuBSPHqnEGvdQ4/59ML6NXCYsv3qiwU3x5c+CFnKva+86n3Jho7gCeIuVGluyT
JaN/mq/HRT2VLBypizmQCmlPnbOhBPBtcNjMPhjpmnnsXaDnWpaBr3NAR/6fVNqw
CTMmWIWcUnnZQ6zui2G+Texi1lvUEKYUC/ZrGIVbzic1BzZxD8H+0QSAN/mxKGYs
yJhkc1MjlXyBm21QWb0UKbIcwCJ3iBAVjX7r6cyTh09tClKd1Y0LtZgVkclcqNNe
2rfhnjPO/eT3KEAZbviRTkf18aZc4h1mC78B++wZpQQWbn50HfjjmUPZpCiPGKCa
j2N404/nZeRXGESJFstGbJjZOq9vnd8rCYQ2nKMYzZiaUCUyMpA/pMbMLxzy6DYs
PZy7ckijlRrFTJi1M8bzGdJXzFe/Z9tm6egf6prSvHukKAi5uvfCg047TbUvkSAW
yH/9CLSJSZNXRJYkKnicFd5dOo+WRfd3O+TDkcYrVJ5asuuDax2cA98OMaa1uDGF
dRP18k+rp7PHTXk3QFpdqNJkGMvRFhwsd42z0odLZlntwduW/pi6/hVy5uBdS+2X
+uIpu/7N7XThZZFy6u58aZa/bw3g7UqoY3BiyKESTdCYaG5+hn/YbuAPqyJN4UKw
ecXWHzCBVN18JskI203qz6hJXQUi3izfkJFcRktY38p1d8H4mnnyq4KYkBXaXzmR
H+OpyMStW1Qn+zZuVs8LGxnooGExfICRnloPkV/KnTAiH+RkN2r7m1Nr6pk8GQzL
6c1JrO7M94IAqwUoDAD637211supdovYPdI+et1AoGay9k1PSS2ctRj9yDB/yXAW
DW+eFoycKTirTln2jQgPDgLEE2xUgHfrJqi+CB7nO/3xgDqw/9wMRuXSiEXarv/5
3crZCc98CqTkW3Twhq4ZmEEA7/9NcX20ep0ko2Uha8gd03KcjMt9wDgo/Aubc1uD
8JamQixcMboyZR9PqMwzRzuLfMHKIZrBWohkHiVGc/lZ2vxsiYjAJY9S3nqHypRJ
fIM9MvafWer7u0YXxH3bHI9rKX/SGA8z90tORcxlw4BKWvbyR1hNrVcHgBiG9Qxo
yqOARBVcuK88VdMu081seWKz45Z0Qf0SLDFN1sYDDYdJfSF4E1suy+UGgXh9bgZH
9KStTWcAMD9DCII0M7lwjjJn9x0vaI83I6xdaNh2ufGUpnKpscZNxXM0xxr7DIFm
kKf7OmfPU8W7aAJ5uu0aZL+5z5+mhx7niuk7gOL7rPzC90LGTCDvFQSTQXbeE6jG
IqNVHsqr+RRr3sKUu2WUqY/O/W5BkOQmifdtujwAKXU7r/mjy/D7qDBMgyFXbjCi
BO4+6dlmYnjZVwb6PNqdb7bWF7edOqhiH8SpHsf7vgAscWvw9l0UYCpVg1NE8LxZ
PntXV7uBaL0HfjBVcZoq4PzRQgSQTTVZMhYZrsbySqIh8UFSnb+YAt0FxZUHh0+i
f+KP5fYuuh73yFyG8dceKaC2NJpttp3OYaqUf8CVWJ3yXp99fDSV44a/nnc6KkoN
bPNqv2PziMiVVIguAt+QLfJoRWdKjOHKkR6Snz53yFClC6Ga9yHRxHAqg6m+aWzK
g7AGAIDSzNtvdQ3pQKW3h2sidb4NmVVht3eKCZJgNapR2NBDIFRRq18hLNaGWgGf
6NOjqDYFMkam4pHEqO6MpgrDkrMIm1UPnqWjJ00wxfTJGcwLGbTHz917bB78F+WW
y951POz1L8HD2Gd4PrVCWjW+74xpGzevMNrJgFjgxes71a7K3gsEdHodIUEXsXMv
EFPWO9pusauy/fGhOyPX3/bqujfkskgf5zzEbLCxKiA2c38JHDmgXr8eyJNj20XT
7kadJ4ZiV7iqg/dwyKaT2ibkiELvD35CEDgqwDaXTHKdRIu+agCTFiXZ//vyT5vY
+bf2Yf0NyThQPg5Waeqsk/YatcK/knrY9QLfZv5clTEylHkDUWMMDBdfNDns9Qli
BMifvy+bpM+msWRLsD0GUj6C23n5M7rUsLj6idcglvLURvNPdpcn5VC+iXf9+oOw
TAgImqwzy4Ct3X2ojKwgCLq5Z3Zqfr+cmI9hh6FnwEA1aXScmJmf78je8gLh+sg/
nNIKB3yGFUFNOongSwLzZoAhpUZaWRaFODSrzg1x+MPASL4J3u3CuTwlm1L9GhLd
cefuR7YX2v4U0pK2ocggbpuWVImnyZZWlIhQjZZ87eC9Vx5Lr8IRIzfYxhi6kPC1
LXMxx4TtAuK0+TMzvUdiJ2s0g9zPNg1fc/1dzSQREzQX65k3yV8rCm3dDjhF8a7y
0t42VNezE9H/n+TrRynB+taPYd+4JiPISVYNesnQpxIEw9jFOpc1bj6bfzUvr9zd
XzXTpnB4OV0InPFgZVjmESX032B6uSzbcXzXgPvi4SYGq+AwR4HdNkkjJtYQZ/Iy
7Rxa267jfsizkKx1eKgA7B7sHx7kL7zmq/uIdP1wVPKYmBZ183hBteFtxxp0TuBi
Fzib2LlEEkXeluUAkh0+kEXzZp6chV4Si4PX7HsgWH3zzSaqbZ1ss1D78pCHYlwG
05QILluGUCSXigjej7xn/rHcJ7kx+tsmdmCGrInsTVdw2g2UeA9SUFEYxy6vXt3Q
sgjil2EmMRFqv/HJtZZVlgak5lJeennWSjuINVZQOH6LCguHTz6dPkkt4ex1/hG/
nNvXCTH8XwLAr2Bfx2pc1qWh960IaSNqrKqlQzDAcUbUnxjCffT2XA+SJXfMQmpv
xKWQEGhvBBsLkSql0HrNp9uGL+ZVFJI87yqadfkWL+rp/NpB5Rx8nkhj5BNP4Efv
lWkxjtGs3mC7iX7xzksgxIDwUB8gYBvSfzii2YwHfgMJBYRWjgABvPC6JkW6WrIP
M5Z04V//GNuAdPlxuPh8J/HxNNf+QRMW6b2kTYMWwexQ8ICuDoey3n3W77eHYd9Z
Fr3FG+Bam+OTmlHxZMmw+q2TiahpY3Sf/GnyZcpKKfad5ujmeT22jHZZ4Ix1aY+c
xhu+uobDS7nP9ZatTiH9mbC5/tf3wOfCgvIRIjk1v9BFMC005rcRijVKnqcg50rU
cTZ6c2Ddc4LSWlULacivnf3mdWcSr4Yz4W+qA6BFjj7oY/QXpRhSab7rYV8QBvA6
17QTGEjp/w/G2crTTNqAm243D0ty68yJME9Q0xPNKbEe0SeL3Y+53A/VjLXu/xA4
XWmdNRuYKkeg3FVpk2ZpNq10qcuCyzo7HBZ003prKhUFuhVgcx7nHGoycR/D3RgG
ZLXNfL1WG52orZAyTlf0BSq8uYS3CTEUOS4qrLbbPUCzlY2f1DMXk81JGhHe2gVF
/Ua3Qt7dqhxZU9dcs9YUQ5Lq5ojWbIAMmiXqOaIdKqGUSAnTHyRkd0W8CoNndoPp
lTnsmTeyvPgnMqNC0sgvgGeB3k3Wnbx4/Arkm3Z5Epm7YVchCRQozvWAaHCIc8Ex
uHoNpnaTh5KkpyRSffTUWy3gLWmBK47wTjvQQFKD2W1VPetvc1K+7m/zKW3Geg9n
g2yfRVP7Tj8awc+l94o6fz5yqSZyCVllVz4RPdWthAPYObm4I28lVnWTYhO1ws+l
1aBbs1If5mM0FJtA6Tr7A9MkWAu3vgy/oOGqXQNsRZ4WK7xa2NtSyg2ycaAU9SMk
MWDeMwmBxsqADk30sr6Ru/QBqA+PxsEbldN+z/Kmf+TnnZxIVCrt24c4QDRC6dpF
ntXtqZu8Mi0ITxNaCiGo7Cc//DKLfttMvgyz+yGAiJGt4dQjEeyNCOLG+mg49RAC
nJ8KylCWUfrQ274LtoPTa2mAluNX09UmaaH8zxKV2r4Q/d34Bsz5M/vZVtaQ22DQ
VZKv7gLY0gHZHaqiVOWHmjqksXoDDFMwRRz0zQI16P5m73Np2vvo7qcB/TzGdMN3
yjSSSbM+PpZQsOwC8rHNigZx0UnwLuYx1+AnxGIPXHPYGIVyYquA8Pj4rCHPw9oH
JbjRmUreCaLg7003SNHfSZfVJMBHm+aoVx0AI1NhHfiWBnIhn7b2w+rM3MmDGEvx
MQV32GT7yiHtQtJLaAP8YDt0JudrPJRe52H04WqSle8wdRLT6ny/HXPaxCeReoie
hTG9CRHyJYOsphug0fGzG9aAud8RtYq8IpAPi0yaGhdQuHW97UIMGsn+xhQHoGcu
u0+q1OhCGZUTATn+6hOgXLv/rU8H0EnWY7Rr8GmovDXyY4X1ZLUkWjKH8sX7SG1N
2IC5YfmIa2P+StaYAQD1kcUsrmYfuAmj/Yk6gieMywRGxiCAYiOABI1y0SOz+Bef
ZH7CM1pNh92cVn4nzv/dsv28f11afEBKEuCYAkbeBLIMD2VuXUjvk0nO8qrRUAbI
483KwOJnAOwtHYfnrPk++7QLBhJvW36VQ69hvhwyv6uyDLnaAPB9ybzSjhicPpzC
ltLmJmBcDpsiW63EcrpN230tmVAAX4BegehSQP8+BNJJqTVsXHba29fz3Juth4xT
EAtaaK31vbxUCXZS2GcowSrKvuoys7J3wXFgWRRCc22YZi8VbLuRrhavaVHCCWYv
1IzWUnURAqxfz99xznQCpI+o7KHye4q9ldCLWhMgpaWgv9TfcZwlefokOb7uERLo
Cfq1W+jC1DgZSrs+axJFxCkFsEjyAlZu9ZlevBtBHahqyJzFsh0eKaBcktMLwCqq
TOHw7NJEm92V1D9Dbk9zPK1SlnebrbTfZ/y2w5KNrVizMJVIswixWR0DnavnS2L0
JAUeVqUHf2uqLM67hK/FmuYYjAiksb+CGS9OFx5g5UsPV6uB2T4bblfMTL1+0Nv/
a5GRYyv4/SxT8jOqSwB51BOJNnoowI8rlNf98i54uhS+SSHeH6ElCZj8g1l4NAUY
V1gVJ5G4zNWJQkOC2RRFJMAAy26PcosTUjt2s8Y5h0lkd4MtfNZrtpeO6S73AQCk
p3cKmeIIazJwogJwwA7OyB+Xkw86/Eccv2Uf3lJZAt93/2E2CkBq+B6ziumi5UzC
QCOeix2CGDiHamVikPFPbpFkfkRK+x+EyR2OJsOVbq78qgdXUwBESWOSvCUemqch
vxE84h7+d3J2JqeGUPH4PMQpQEwPguh+8KuG16TaPkKOyLEYl6663lHNXObhY4pi
SK15n9fItw7VUgcCmrklNdH0XnQCEMRHAxVUUaYeb47d2UV3vePCqAPEhfmEgeqX
64J4Qgj9wn7/Y8W9QlWYn/j9udHwygqLej95Q4aUqVSWy60mQRoNdUhS6B8C7+V8
O61HM50ju9gOlXNcfchH0l/z8+4ZZFJb+yJyM8Xd8AAyycAEQppeWgZpGoCT2JyY
RwbW3loKHfeEwCfXCBPewohgGrSAsKt6KGD0d1uSh0ujvzJBdQ7oZ/fBHzB+3jFB
MVihaNfcR1JPT9oTaLYgQ/H9yVDHFQ5PGAIglEBDcdTc7J7UDpsstPCyL79LLLPi
VirVVNbZ/15srquUDJNjrxI90oDxw6B7Fftf12uPpqO8CYXPR/ZKWxABL5GbbxsR
nFxuyb8id7bTV0t9CXfg3GVW7e6MHrBUOhQnAnOH0Y5tgaRW326foMowejJLVauf
H17nECu72eZl+LuCj1nQ9t5EGM0qUzk0cbeNqd1cYvm4Wdy6M2BSfCzAtwANyfZk
b4hYQAD7471xP2hRTBSQHBjMBuKW3ty5uKuRb5loRZ0D5eceOoNUuDd65lIAB5Yo
lv67tUeRspf7wx5EPvwX5TB0WFhCnMwqtzMioN/HC9NOEiqttYPlM0b3FyseneGh
om2E2llX15x9TTz4qjCI2xr9Ilngg4Quse7ZhxJuSR2cU5PpnzdqQhwmgFFrf8hk
fLIN7jKFjOK+JLNxPF8EXInnnDyj/Qr4xqw+ltXKghkDseXFfAhSgXzEAf8G6HP/
glcNcKFeXMtBIN5Nk4nySKMTWWma7js4MWWc0I4kaZm2sY5SlwjYzPas2b7a0YRc
R26VgaSaoMckMd8WeDi2Voa65Ptn61BHUGD3zHkUhf33bgTFWH+DpWKvpRiJuuKx
CWbXTaVobSwhMEMripBd5k3SAD+ctPEFCDRdFNm12mKBc4IN1OfYooRPBqhWu9HQ
sgo33CyK48hWkuYCV/908PEeqWgDEEir8Y80bN6LUh9XZXViVrILwCbd0KNuSkFp
jPnng6Xvo6sH8NBTrTsq/hHwhIbRS1j5JG3NWL6Ni27SvYcW7z64C1vi1wBEir10
Stw/Hix/IC9eAYf//VloiDqx7VKAgWzBPgqQ9IXs/MUjTIzINDfLLjzZLqoirWEI
RzVtwTD2fSNBmF5CLHGWUPGDZ9AN1evM0cAh1oihMlB3kVNWBdxMk5lmh6Xn2nqU
joXPyPcAlmQfsP6KBhoTHHrEwlJ5pUgpY9kvLjlLtQtirBZ/jo01uhrgz/A8XgxQ
i8Sn4qINF6rJk02gTTBiOyz8j/esQ9wT++GgHxjmRjU5kIN9vpVljkwdxPM9sNMN
M15bdSi/W91skoUxTnwcIkflKE6O0b1KCO36e31IGi4Q//Ge8veOS1xzhMOJRBMt
IsOKBpxI/AsKmON4PnZc2UGMOX6eu/zmAaVv/fJC7qFcEqHoyzZNrZKlIXzdmug/
a4msDumJN4wfvsg+NCXy8aHCT2fA+LqO3iP2PAU98sCuIcUqtykS31L4rMaY84no
Dh44ozpyqBtz7anaXDRu517f6OnxBQO+xkK7O3rXY0MS7iC3V0yyjpHROXRHAL6V
3JAs8tJ/gNQLR5+AtFPebnB+zrPznMp97DWyEObLISW3VDC/iuAa3eXBTd100VXE
ABPeoO/kWpQtwWr6m/Icf1UlyWlIao8GeOjlNek395J5aJ+av2rkBe1WIdT8Jfoa
lJXkX7NZRlzB04iMPxziAG5GPO4xeaRiuy/azBWrvvIGpAnvxG1w7Rc9ECZuaVS1
/mElKmVw4B4YW+41oio1OY6YTzLp1w1spajbYwhYR6jPT59oV7Ito9T8jE+SE2cZ
4YdIljOh+jWVhiXO/zWO0cwI5UFvIR/zdB0LqGHrNjnHVllz/hBRUvDokgSVkpGq
CYh50eQrraqdF+fhEoUKnvvJU67Bn+fiexz7OayXX6IWflys3c69uSe2ABHorAXe
BCdWE4d6ad933wn71T/LPBflLlbgi+/N+ERqR/aOkUlO7wQE/FwOaFNgphzOLwj1
CIpsAZH6wPXMsX62Dl3lnmkfHMcTMCs4NixviDMyUYy++nsK4hQjF5s4OJxLpgjf
rfnOQd/1/A/A4djXr8InHLUHTLR68gbp/CNQDc+Sn7JEpHwbStwur06fT9BsyZdI
D2snG3xfwfo6+WNEO7Q9zlT/PmfW2YhMOQqQU4Enu+ncmOBhXsmwOrYHis2cw5kU
/WehsrM2YWWxfB5uDFQ3jua91PuEivleh6JZ01OKKL5tNHNI8wnMR3wi4yhAV/TZ
D7cw6YYDIn3L/42Ge7lap3jCl7lCmxS9cqRbsc1FzV5BU0tQQs1IffX9bjGN9FSI
fECLzoa0/rpLJ3nHZJrRqQXzAzab9x4R8azgKH66rFGiRBjqeYelwGpVEZclfWSm
Or5sMRU5aOP8gcTV43uU4JgS0G6ljiviqQbrNOUNg9XrLAW+r6Fu2zML3YZbymaT
2Y/EmVRqW8mCDm+c9oyUZgsZZExQeSrh/H2uXDDRCeAUoF2qEKJa6z7em0njthVY
zBGO2SIl+eDrakdh6DJIPe9tB04HpEfc5b59+FoGj9J3EusuiW7XxeIaiW3b3yxX
O3xICGqk804u1z8rdorQPV0eNg0KlY0MCOTQGl24ijCfSalU642CMfSSNb5dr6GC
UFQvdQEnWmBHfYBtxD4GzjeRCpZgyXodNy+vFHpfs9vZlbUxM8aM7jsLEEYNAz3d
R3RKW3AcdyFPCDdKxY9haerBXe7PPZ5Ybl0D6RicjzJxEHGlOGqJtTyETwMAsq+3
pgr3+vvO9UtayRtPqoPbpR8fdg2lUQzwteFwotZrIAx9hpPyxWbtRvEQ2bmaBuUG
RzWuwAQ6kNbI0YOPFTcdxmDYYRethGSfZ+K0/EzdMC7LOrORCKidllIFeMobBdQE
sC3nRKP1SlK/E5g+MFBhzIwpPggI70V2WgyJOx0PtO6IR4MeuyXF4Zt59Ci1r92s
2+rn/UvQp3+HrdvGItbNaOILIzqfIb3JiIbgC4kbYLOQDzp9oaZBSipxu3VCvjKb
jwv5m5vxqdpYS6DwNCFMrBrBmpAQzfPg4ZYYinSgVY+mM+6BRow1nXdQg8dKU/zO
BQRXwNH8rcc7wVYt7Oh5Qu5nR9VX5BNf4s447BhF7+vWx8RDcZrBp0NXsYU/MXY0
WPGyZrxZM7btX6Xmt1WTx+kWHOpFCB7IQ4aXDlzrwD9sSiKCXNSHz/QK5GGps/S7
MPDIfHhgPNyGfqcjrVaC9PvkeS2O1fV3W4qYEKveOqlwRuB63Gwe1OhS+kfweMxA
EKyIeFK25nE3Y8GgXx3DSfCfZhEy/ZX2vNvcGWVgqK56IkainpbIphVMo/1aKb7I
NqFJy0M05xKdnYYC0by3UKTTJXfJSZhe8NcuT8Ap0WD1XyMEM9z8i7Ta2kSVSX2F
vmmYfGgbvuI1XXrweVq2Fw7sPHVTrPQP0TvH55TaDqquOgghJjCfvFOjTv82ayaf
m5kpQ29Du4j9TyY0gHdkDVDj9lh7rpW4HeJTDIHikk1skz/8Bn74BYuYYTN7o7OW
Uxx515quTudN1nfByLGsjXaiudBEVuEUsZd347Mazw0XCKfZi8y5ImG1R28rLwRD
43kXDkZq0CAXhHmGNtB3V8HL/hYLUnmjk4SLAhKCmpvGR/IkBBeTtsCPhNIbqhe1
IS3fhvk1cCpX1CYmYISEcuaTV7SntzXFphqk9CEzKB7hEFR23vvO6iawUdggERPa
sx/pFcAUqASWiFN/cyjMslong/RSynOpdp5Q9yt5fg0LiecxvYLEDe7/tXgwcz4u
/yAy9/wIG+bZ6h7Z7pBOXolhEmcRzjgFg4N2dAI6Ym3HrMTmGp4tVu9TBMIb28BZ
guI3zs2MEmo4V5LG0xLaCPHbC4LsICU2erQlvgEtf73+UOcx9GnyfvVnpfhszpYf
KQjud3BuM+VOOnoBU3aPTkXf0v6pspFR3pC3HKDe7sC7J1rKA3V8WD1Pt0r7dIza
luOggwwA6ZdKK0zcwE6L9bnvDLaGzgw45mAcKubG6xrMvLkHI7Kxkk6wD1mkhS7f
oYNNZKfosWkEaHU0N6fr7j6voI6y/GdyrhaB4+2IltlG3r7T48Zu8yPx5XxxMfKX
ekhhVsasVIDc9Fl7G1qzOm3SfrIdKmPudjiQCXbsBXKcA6p+u8ivubiwiRVYEISG
vs3BSJddIF43TNQiXdCR0UHClVEB04BgmudsLWb6zh6G/YVH35mT7b9sAPDMBGA2
fTdx2qIBQi5CUkFPdke4ymyoWxXo6XMHwjNxpvnhF2jPfGnzcVAtQlkep9oiWdLt
qnDR4cQ3RyY0GuSgiON/Ibg818nP7VQgpnCfb/9ZS9UckhObPakevG8XoKeDSIEA
Wxe6NSqpdL6BGzMyN7JjP+4JdJ3dBIFQRXfDz1l5MUoMEGD5W8quwrpa9q7wzoLY
qH5oCS48FM5xA0cin0/mIjp7IdmCqaXQuL7fOl6U42ZIFUWHUmuE8FcwCaYSQ1Qp
TjVLX8UoxQsuxMrANhddzSrjU+RWZBabcWSt6GaEXBiv/zaj/VvrONHgWgUasg9E
Sq/GlbZGdFAat36X6TwJFYllt4p9zpBRaFMeDCoKzJf8EUSwDwDUt4D5CXkYtUv3
dFbX3zMUKjE6NNoxS+ao9L/U1KCTdYaKo+dRpEpY/Q2mWQ8jtuNrnsCEuKihGO4r
gbI/OUe8ofQottbF9tiyVMReqxhXDGZeWB7tyDKUQxgo1w4JULXDFJ+ok8Zr6oeN
IjwGPFFjzGGvkPlbFfd36foanFfhGZEJvkdFqYyGLtFlcKtqmuhGetrwjVdtoOrT
UIItWRBdoW9Ro3nZnW+BGizXsTKPdY6CChwE57zewLv5X/2N8/lp9UHO46UFMxeR
pqpmzHGD7e4egBcmftCK+RGp+lD2rh5dtWDsbhwixpG9jxpU+RjXfIMDxw+RmdfG
RAXtNGWaS6pTnQEuQoTlNnnVn0Q2em8AD8h61Sk+TDljInvJZxTVefVITOEqJ9Zb
iDAhCMqv81X59HnU4ayS+ONB/HU3HXZ4RyYlf2hMFjmAi9Sb1aHHk0/WdEWWjt5v
0kdMlnmHFMOv4TmmzHsVzczx0LoMJgCRygW3zkWV37ogVc6z/Kr6tn7Jj9OjKADP
Gw9uIR/6eLY0qn/T5/9pCKXvkezQMKcKTdRSCTHqTnJ4TMXAz99yzQcJfkUiYxuA
qwaxTWVunB5KmF7ZTZTH7QQimi0wmlpyJZlY4JeLq0mcjAh56lY1O35YWrPnQIuY
FKS2WN4zXA3Hdm72l2DPA9LAW+uZI47OH4QLJ7vxPyXv971DZXvoRp0AGd2jda5p
GGirf8wpIkjm92OhC2Farls4ZRYPF294KkKPi305Wgekg79ead8FBtQ+dK2qwzJ5
J40NilOOyACys7pLdpjFyol5twoI5v2onmuR98RgbxkmJfbJEri4pZFXk7QF1Nis
chsowlPwR/u9qbKw8YCHfwIc10/kieuIucQhs4sX12eo6MdheZGKUpPIONhMAc6d
7kjsdgbMmx55UdApEN/S2u8Ok8gjbXYk3yrSQaaDN/zov05uMEKEkNTlfNdrCDqR
Dp4m9gJHSJSA1h+UxhOKtQIMO8170CM2/XWmlEFVbg/lR2raOmmLahpTIfald+Ok
rqHZI49a+k1Qi/FmDOHtx9HCHrsjZZJHPPTDobbFZb6VSXLcFXP8cIXeT/WbSQi2
Du5dkfbiwpUDjgjN+TBXSFH1FZTJuxBYJY+HolDV6hTWXGG2ZMAkqqB4OGrRbiWV
4ulP8txsB2R+og+HwFmje4C0Y7OKkQvN0U3KjpuYppMDd9ZgXz6Z4xiASMdjKfk4
eFNXBEo7Yo4uzmeyZJLCWkZFqwT/ZePpj/GGVErASQNKAfIzkwuS8LCsD37eCrzm
M8DXt5IDy7jEwYVs7nf66R8LHaFYlXhXCgvbUs3JGcFgIDFF2uiYpybfKhnAwAWS
Qg1TSuDJ09d2MSb2s6jNPF6J1I/M9eB574d4SmfyqcxaenATRNqu6DJZ0dGx524J
kE0zdWrvcYxSLxOP1Rz0CBNHhGDhdgY260RUuBGPGEPzGMMjb33e1wYsoeShyISK
DOeLBuUgfL+RZVQW6qfKUjvhvfzn4uiCToWYyRyhgLeMTItjVPjp6jZM+YOu19Xk
leWtbc4D8L319MoOYydljF5c/PYYryrOHDOa4nBsSeBc0yVgwOxuZMeowzzWaqPt
redjTrTu3WJyTImXAkvSVP1dgu3poF5f5qk0QeGbiBL96/FLtRBP+BsDl0nsGKT0
KBmrGA5iUmRb5P5ukZKsvVfyhtVY/LTipVEh7Vaqw2isLFzgtQ9N83HeKJfrWkR1
pATUaSW4N4vHtitkzTCFjTNVTN+BeMdZHDrwt6hmCL14nexepTk66oI69i2+M4zR
TUdLwaIMjANooVl2nC9vZILgV6EVAV24Xm29QnNn+IOhh6hO8F2TvzGpUhPL5Wkv
pbfe3fc9rUeoBWycTqUhQd5BPRv1BPsUYzlDkVH61o/64o66fIpB+L8UZPGtDoD8
cDhlsLoev4dzC3Lu1i9pZhzi2g92EFxpAnXHuP1Hsa+8k5zz80yx2nVcO2/B2iPM
G38myZEArlZhDeXNTFHiMA2DXWFxGX1CTpTyiahx5fgZAJ5fX6ZrTteZ5mSdnPpn
mX425mhh+MOeMjz7//P28uDjZGLMcw9Vv013/AUq8HdowB9yH77SVX1NKHHpT7X2
lcLgVTYHtdFmRxt2HWgum9ZIEL3FM/n40cTwoLB9vzkDYS6KpylfOwIrWN6nDs/8
+igKUS/CEKeD9NbxnjDuxB2P06Xy81xkRN8kTsDX/OO/HeJxgU6TkQdY/xfK+ZQM
PbgRDpEGrSBXq8DROc7VtztS/VaCj/NQY6jywZx+XmSPLO6ipX0sFGfd1kQ2M+Hq
32Rf2KKW8y8A2m9yU1oPU8TpZ492dnqm5AuPdJBUI3r/To2wkdjMP60vRmECUOCR
UdXTf9dDZiDFAG6QImkMUcoxLzkuPjvI8nxaCH0JNiGCa1mukuEMKKeJvviRXS0b
ySrHr56OpdiAWbZtAMr4Y61EtkHTa19TDst7tuGB9htPk9BGebOjyTkWw0umRBW+
YFIwlr5Kwa+iYViQGOP9XizYDpiyA69IQB9VRLNz3sNI7SCpl5kZofRgejhpQGg1
yitw9nL91wPlTW0QTgOIha2BJd0pReosoKhu5BJhsZ1aqrR09tvVJFZ9gwka3h+l
JrtiTS7VQp3p7U/B+QRu30VUIXngBlGNV/T4Tbra7W/tZo/4mdbjMAw12WA8GIVG
KMGCvYgH3719wnd3tiitAUvPRRwp5MJZvw1Z+7yLe4JBMqA/NGWV6mIHTOEe/DLF
tqQ6CZuRfaGCFyiWE3n6km0uYv8sIA4A/CH3Aa3XdvXsFytfJriGIZERBPjjiD+O
LMafLFLjemRk2op0oZgawaLrFADa4HWb3LSBezwSjN5zqulfc1M3jqTIp9x6iXZT
dbOuAiguDhD3a4ZTfibLet/mXGYfrlEuEoSk9redexajpHbOGe9aOCGLRuc+kxqp
btmJv1UG2noxuq+8G/LmlvJNqcdM+ZMakNMkdtjSd5VxyKWN4U1lltUuYC+sfR/G
1lGgfIqCwQswQAiQf42ozO33OyIrSObPMfsmoNlB3ZMvxn0Yrt3Q5dfR5JXV4OPe
G6e2VBbKBAH/6LuOWnX7NKS0PV6jVbqsDHWLNwnNl8Rga1DuqX2pkBeMzXwHE07n
KrLhmlqdOp5jjWCersTFUClQQvbzwRg8Q/yG7eFyhYl0T4TnOdWNxd18duOOkTzR
KHSh2Jw8e00rMpQwDV0Tqx8Aq4kSHFVTVp3POzXa5Jz6tgb8ExWCpIyN2mnE6MWl
x7oDhzH0NJLl6cj7hxH8AshQotPQ9wtlDekVrUGsyKKT4gaJ27fOBq03s2zGg4Zx
5LqPx9zBD2BBqNmbReyFN+cQnENUmaLpYoCTXAUEYk8fjGd5Hf1vAhGTNNHaKX6c
yYF3OE++ZEXqGJy2fAOr/fJswbXnQ5WkAhgpqUBiwPgVnDKMOvnzW7vwJlLDOIkB
A/wNCn6kqF3XZuE06j/OfcwhhEhhS0w3pomPxTe70w1DHsIFlZJC0OBZVcw/t8L7
nUuwN2YXVRk/z8VvIzGVgCdZmfVIDBNYdm8KJByIvxXU/JLaLRbT4Ro11sqrFfp/
vc2tL7xtB6F88BK8MnyKoOmKVwr0JM3njnsRRyU6c5GZL+wmIGjqLqzLeQvpb8JB
Yfghi3GJexZT5tsoTXq8ru6m4mRWzUCiIhnhT6tx+PZo//RIx1NyQzZ9YCpoINL8
iVN3eqCW28a+s1lcX5ahwClz93piXbjF6FETv8bjiIW4PxO6p2U8lcDTNCHROgWO
5PEVgmKPQfP9jG2YA5910cXq7P3hhhbDNOqx1+NSky93V0yFT2cmbT38yx5hyITE
mWLoJHTBoUTpHGEk8tv9jxq6h9iDialPVVmrqiHFO83zEkqDCEGPSr3DdjkBTw+i
y7LwjH9aFNM1j2Qab2FCttbgCyMiIED0TX1xz5Mig/QGJLKHYF6sesoJPBscnWHx
EvCwO8A0qLssHlGMvP0qRlRhk9CY17SGqyigJVxIRuHdojKhemGux1z0BCLvzae8
mxK4dVOhhl4gyfBKZNEytyFiJTVy91c3IT5UcCDCTUTGunC1hIMpySSKu6ngbdS8
FCzQ8qMvRtZFqnz8d+eHR3qCpTE388C03uENiyHmKQzuoYHZBkVp/ZRKZaqKGAxo
lilbYd6mxa6DQm8bohKySBqEMc+YdtNmrhDayyC1XFDQXYFBFroYD5rXGFWFjdIR
l3XaMvCX5Y2mH/rwMjdLfXp+5F0vEyw2brILnAn1GxUFaqwAVVgROOi5rxATCo6H
Ww42U4cYQr7l/e4h7t3q2K+3KXTwIPXonMTYelOhRN6jWIGMNv1zhGZKhQ/ajnur
f14uZpcehyhgE0iCQMt/ili8YafqQMCkPGAQ8vr8M+6hdx4CgYYyUYwAI+Gg8ii1
oJrBe7zx9Sutu1b+8UeSxQf7tDFdLjKJhTOc/tjO1w8Gza4O9cVo8UL90D8J6lNR
pd2NZYuMgzFMnRlxlb2n3SY25FXxQR3H+N83p7Gdbdg3fW0eQKkpy7q8Wm4jtXEW
o3I46hH1snv8sv7VYzZrzaC+xDNBI4QADSozPUMqRuAlOH1Bw6AFRD4uqhHsza+2
Q4ArHshgdcitUlYIKamVwgvAI+XHQx5ceFusuIZ7lg8E7OstV+Um7usJjITArmKb
ww8BZ4AeS90iBU9WdIFm1rEKbkdBjgm1EiLBja8E8e962ECzzSHLDWmQ2DGFc8wk
rv/X6VnKXwmryXZ2z8/3TqeNyVE0c8W/9WwNIAO9gpKcjwuUdm+SqOQsGaVfRirr
BkdGlUVO2YuvIiRkvVYqY9fZlKRtCW0dc9I1tR8u4zesyWvA4yq+Bx9uk6cbcDnp
4z7H/s/wL4Tai5TMLC8rtczgyc2otJds/dYXQ8XQOfArgW7Db4bmYE5N2hQqqrHD
gOx6hOfQaNNgiIMm61TJvQlJRRu/qmI42Vd0BA+FKbJW91Pe8twhpT2qz4yL4K9q
f1hP2vRUeXbCeX8SzyiqYeTGLp9a6Xf52DmfjUtkR0LS90BgHaPeaz3/Sfxc3f8B
PbpVATMt0ImpY7+eOrBJXJ51c3nof3UXQOXVnnXnD7kmTsTe5hVUIi3VNsNCXc+A
a4NkKG0WSQ/nUxz7pINHkVUNOvv//+BbrqwmQ6AUr1RYvavIh9ZfmzVellpI9jec
4wnLEcN+LS+aDIyvoPoIZa6QgBjN3dqozdphQ5K8hCjYpBL+2y6y6NBNHenY9h8+
qu6sjo00ZFGst/w+7ZKJZFNDM5cu3TSoEDKHotuMspg7QREZaC/dQIxOY6ZClbvI
ZlCZi1iAt7IfRkzmH0is/CA6RejRzlnZz3utWhkAwF+t95O1S6f3pbr5q8rWJMvJ
wcB74L9y/RKxxEstl4XJtl6o6+j6pZ07Y+CsfISxP5ddbgstw4x/PxOHUaw/GvhF
LdpSFytfFLg1ysExCdO73UpilDdjz/qxwArKHZxaJ5agbU1h/LZxdd+A9L6gunxu
7oMZsTHwq/cufcDLV9UK5NrLEyhz4vXpMmM5uBiQELRhmuhNtv0a3gVLkuW1JEgn
r3FVN+4HaXESeNK70EjPyiWY85QO1WWFGW41cUzC5nzarC2pluXxKwQocIgPQ8Dk
Q4TtMq3iMdb3EWQgTppvDFLi7J8XzEhTlNN80RM8PMqYyaNFyrdZZWxQIAkIOTTX
+j1dZ6KA2YHQH3GQ8HymKn9zC6jC9WfVFOWpLfV/lJGFOX0jdpYxGXrXlVkIF80o
fg/zYfv52rCbvG2HASAMyMW1HI+qOUKMCqpwODVW+g6J97hyXlNImVvo7kbSswg0
g1iUZb445Z5xKM8hswM/vSrn4JUvRveS0YLchosrEX3nq7f6LmJsVR9PjE9i2+8X
vjC3kfUzgsU7luaPMrJXIGYGor46u1PQuAcXRiShgV2IrMBIqUiQhiEQbWEtpYxv
rUK4+JEALtOEpfh8tOTyJyYjuC8Xd07bqU999axgX4sMdAG2DGPBQt8b+1WYTGqN
8SxFJDSyfaGkbRUTLQYezzEOOX4t5GCYEtVXblHcnhmhaPJ7Bu3ZeTxCIMH6H6+u
Ef34n3mqNEu8dCtOXY6CaXnGGxxHUHMP5t8K3NRsRCS0LK/iPDFWe5v4WR9IasQE
Sch4GCm4eojzmhFSdfqksLhjLjgWyXQxrhwZtyeilzmPWtjUoIK3OdlM3QUWdP03
7B0CNPPYv0PfxOC45y9pMEX5Vz8qwDPyz0FG+uAlcSLOrIrumJlr3SIb6tSUvK7/
5rJcSjYV+g4c3mE6VqHag3BgZtPwWSZNwqbW9wB++PYv/EHzviLlTsMLKskLmFXz
Jit1MXTP2Fx70bG4bh4sckpwI3CFJbtetiyL3ut6ZcHMHMQ1h+QNuhCYVFsr7RsY
+M3NjXHuh0tON/6G6oRtBAkJZG2Y015VWVwXaQZVfQn3aesjsuPEoB/3SizEFDfP
F5Ou6aJTnPoXcCUchXanHEQZpV420UUD2qJHWdanSaIM+v2KY2LZb6/gP6GO94iM
knFYaAx7J/lvBwWh8/Zp5gBIZ0ds+5JK/n1ido45jSQ10UHNMTRTScPSo8If5fKg
GhhJMmX1RGd0gZELOVQiMpWPv97eYBHd7NbxY6GroS2ehvGOUm1EjChId2HSLxNi
GiQ1yq7B94/nHeyAaG0LXqK5YEIVbf5HAniC4BAzqg3DRZETexRumMiSY01pBQ0t
r8lWSSV6KaOCbQR/75IK1zVA5N6+Y98nF8f/qkPM7ywCyP6Jl//s6ru+xVmR8vlj
Rw0PJtYzWYZ1Prwr8Yw2hyWcb5bqwTD+Xd74J6kTvfw6CmW+IH2g/PDxCKe9ntUD
9iM0XVhX9yk0OaNi8K7ABw4O7KuBsozEiA/ATKx8eZBuCaHwNHW+LIJxmdX65izr
k87gKHk+5bN8fxIggRJEIGyIEIS7X4cdrqyrs9xXlaV6yMuohu29d8ZxY873UtJQ
hEPtGJz1HS8dkKk+zR/6y4W84OPhKgSph79xXyAIoCgaQlUDVxD8W7dBapqijZSj
pQmlVLjPHshF7r7TNwPFRrXnNtIcIsnSE7MqKWdSm7H+LZndxyUEYsLBVoPFDGfU
Zf2P9TelDzaPjxIyUR5YSw6dv6U5WJHnN7+448zYXsCAB8W7cI+OP9aZlZ756gmS
Y9nhQxI4eARW1deLobWtAkIEKJTePZiS3KcdJGQA4SXiq/mSqUv7ny2jx+7i+htB
hsxdpG2NgHI5YdA6SfMspLk6dN1ih/FEOzKEMfTG8mPT3PrQ6RN1yp/dFzQxHIr9
MJhfoibMIWk0B9yRSbux2Ci7WPMSuBNpXTNyJATe6GpAyQcamxu1RaTjHGmfoxJw
rkW40uf5fWz2OP13xTW8/5BF1HOBqlUetM++MZZL9KLXlrhO8gyCLgYkkoYJMxQU
G18Wdqit9T4htC30OcHn+tRrUg65vM19nC85qmyAS+fVEYWzDwTqGY6VlBcaR7sz
HL3qelHysCJwy9AXlTbUgLiG6Twf/QCMVPYehEvXy3zCWspKBXRNfACE1mNsb7r8
UZob73NbB+VIux0s9ddDwBhcVvlQ9any8Ignz5fFJBCfSQQv7xUZvyKpWV6fVvER
ka4plhAjQg1efqzg1KP8DToibnRK0O83AZ7znjW1m0uGf8crfAJyWVSoVhhA3S/b
Ti/PV7113/DdOPdJU2NJBDFv/fpOJhj/nPHxvggZ7FK+gZA5zQ2iLm90zmNImCSm
kEVhv7fotMK/0xo1dP8Cgy2i/jU3HgnORQox3kleAfplpmtCPwbNYAbbxpqJr6MS
WDKynGRR+4UxwGubbllng+RuvY8wgqO2U43IDz7a2ag066DWtd+bk+KLnk6USfba
GxF6pYevUmH5fXaaxaT26pzx1n6mF8xx9N6fPD8VuMaDx+MEwbIrmS0wsYUZIEHT
OQEXSEZV+yDunoBvdI0ArFSSy3U5LhaH4NY5caCQ5uJkQJbfwqIBB7C+CqG8Uamy
Fpu9ZYmc85WjUtwe3hYp1/ji9U+zUYCFigAilr9mFsUNJT611+bs7DGSBgJ+wAJR
e+u5C6WQtseyJETFR/SsAJX03FQ1HeTJQEM9yhuyIZMo+5j7WOVZooaxshW1GXCB
BW25g6NU4yNaGySONZH8q91R+JDjI0zpcmeRhAB00+rbmYgPvEh8tce4k5D6BriP
cozZMUKVfUB4iRg0+zQCywpZd1QTW4Zmk/+qX84jOgSPek3leb43jT+8JafQk4E4
e35f7O5mTqgqBFOz7eidp8ZEywvQZrlXj8PtuCs8O0FjsmYT72P6QPX3M52EjXub
1rC9Pqk/d2O1YxzzM5uD+HfiY9Ss347yvBwq4e9oseVZdimY+Fa2U0pYxp9dCml8
DVZf6N0JuUA9y30nm/PirqJtpjwQDk/DqUJ12DJY6uOMX39Wg0qbapRieheSsd5g
ph8TJUtK8TmQnC1IK/O7VLBMb+aOZtB4nbasz3hsIACPr0SHV2C4vdyolfZtagB6
15i5wLY6xANdRIXs6hA2Wd3r4o+Ih2kijuhqxsWA64IJBM8ZU2B4QRh031517mmX
/1XrhYPpOmKD/e/KqAuJJcyfIwvYi8mlZKJYYAsNc8rfEVbeZjb7e/u1GrxM1wsP
lA9s3Wsem/8i7swQK6gxJwEkwj9Z6nVw190oTqeMusQmUtH5Qk3/S91OWAhU7jDj
ZA9iouVggPiRLehsSK6WJEOgC2/kOPyoUzZ5Hjapu752HZHkQg2YZKVabpI5tIzj
nPWX1m8ABnn6MikqgnazA9/aK3r33a0V679zAT1nlEzsmQGE5hdxv9Qm9nqrVa5i
TXIViurH0pYlzRAMv7hED6pNmjfH8QM6z8BDIer66ToRgsrsNwp67kUVQPLUapDY
sqGKWJC5soBJWJ13nnQrWbci4zupFOeAhfyn+CDNK7Wa/FTVuL8ZR5/RDbTT2KGb
HcI94oFdRh8eSISpDLcO+41cSe8jcgoyaBDflhsuFKkDblzi9lPfBXlKcxxFpLV/
NDbShSSPoypSHzpHmIOw/2SIoO1HXj2Xa8VTckpU+PqpduktgdoxqFWxjX4NHr4H
8JqK3Gb8lwjzVbGMj+Vsd8xyzuExufePSgC4oy/hP2Uiqt+A0cB2LWKsKxksDVBT
/NbtMXhczRL6/TjANREPuwWkbaj9Dbw6a9+YszhHsRgbz+JflEJ7STJA4ReVntqB
iyNFEdq5HaWeSXApmgJQ7kduaTm2dMzV8mtCqtLyPZ5kv/QH4ysFttz8oMy2E5U7
ovgifdJmGQYOTf2RLhqwjPmK/eRJ0tfxp/bwZ+ewuoHsbrKVIJNHndImCAaL6b8r
SBwbI9h8PCxdnqyAtt4OrnT8pdMiUUEiA9U85mjneATLXgAnb3Ib0FBMXHu1VN80
EemIvEyoN0tifJYo0kNtoVd2FAKsWPISmgUQlx5FtY5yDMgmG1Q3iNduOuQ4os1g
l2QzrJLFLf09xw34jLgGRdc1TJewx0nU7AJQUZkzrvtYquFFQLcrlCAz1+3U/EZA
TetPjGk6+n2JcnH+v4HyS2aPkWprzEcV4MUJnp5SwQ5boC3tkAqQCW6qvu6jMPSS
ao2geBGv29EfjGc0R6g6Y8Q+UKOMGMNnks8lh0OJTNc=
`pragma protect end_protected
