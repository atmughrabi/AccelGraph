// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GFZTeoErfJmO+1vDTq8GW+n+gztSYxEP7Mp09NWlTQqj9V8khea+F96WM8xaHaSz
3lK6SFYyFY8Ky+IajmuyksvyPTCDzt/JiDzANXHjhf9O2yWmRcyNdG3CMS/CaWbr
eezDN6CqDWbmNHCcCcHeBJvzOC8JVYs8pmTv7gJOEn0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5472)
zRrQMOSDrYt3LZsS4GDKpKpSz8dIG9lLhpZSVvdxdQ62uxYN5JaZaoLyz/Ztw48t
Da/muvQ/5A7HbD2+0rElNMLnkaLMJZZSn+87lyMWDCPUL/i8Jao5IOxylk1KbEPG
5zz9tqci+Mt9nUYtJwaxiImQUJXLeWDr/4mvrr8eS4N7hFwn5wDw9yTrP5K7RKwq
vP0cUXS5ycRgpIgl2PuBN3GD56Y7YPUGrYgiVV9ZFG/4EzKFhEGoNgDfDq2OtHoC
CzIT0wMElG60+K4ftxq1UZnGWAfBYMq6lvOrqtzggQBPa3VEuaBGtL436pEps0T0
kA6CER8jXxzRxiC1Q4cEPf2Cah/a/CJp4BfWFenQu8oaBWr9DwNhqFo53LDnNSGD
s99ZwlgqbMKJOcv5QVDpbkQ5v+JNp8r5sd+9KXer9sPkLaoqTYsdG3hBSFoqW3TS
c//namZ1T5VFXImTcjxk2P6F2RLerzZTJB+nEberOaHcFYjW6qsdLIsDJmz51Nxo
XK9mmFhcPg52vQRFZLyCH+lUc7oKrEO2JoXtCF+FALpn4Z5gQ1/UjZiIT2JJEuWn
/uiD3dBj8rnXwSek2M8ZQ9uMJN5rci/SrvaKBCqPqQbXSGW9305Hdww+ELlkKtqI
r9ely5IYIkYz3b6dquz+Nfr6Mtn5kXgo2aljtP4YXr9VJ801+OJsuXzpMfjhuBnU
QQbF0Nqc19cLlch2Zb4TUm9+XgQLU3nQEWDqX4J9bMxD6jTLySihJ0W74i9ZRSmn
5eEK3pTpQILfFA0ioglIq8XaTx4Ll9pegQ2dyqIBtR8cVjOtGVhcloUD5SZeIhqc
B2KBUzrgrycEMZwzWTeWQoykVEWHvpV0i0XZsn+hjLlW8Nci+/FTOXVw5yDuVTVC
H96fP13nIbaHrd2uRyn/TB4tOlSmgVHis5736lqWur3+8muclOGB/cLbXzgYCEAT
o7IHtg9xr4JV6Sitlaz15VNADElpmyGxGouGT8vSvqlV63C0pdFSZsbrAQaFp+2y
ey9fxq1QL3iXY3CSXOvPMT1hFNKpjJl4u5IsM6IG7TsulGqaVXchyLB2o6uo0QG3
HsaVfQkRmtgspYq2Zc2cELZKri0ULlkObC/9tRnphgkg44a6uF628kTKEKJCMz86
Amm02K9A1xc/9fRbu5uIScDM0hYAVN8G6TfwcqEW07hIyzDmDWKdosUFGyJQ5Kqt
Y1Tm4pskOrRzhdotk6NbtS4Bpq2RR4A+EIoucehiz1lSfS7AHYtIThsj2mIWqMsY
k/xxx9OQUJ5UEVtPPSihW6ZtmmnjTrtDEXcOkeOfWs3gbCDgFyM0yZ811QGas6z5
U9wMNF1Dq4BLEVSlt/nDgluRePPp/SSNcJ3+M0JaPOEWTJvgnIRQ97rDa/6MxSq/
5Rx9Dsf01OME9/Hktu0ZDg5S4bui4lz/Py1e3xjUWKrxY2eWZ9q0FtoL/L9LgKZG
PanzDZ+/dOrgGIioAToVbr0DHNv82Q7ENbxIFnxi/suyCKVkwWNAzAoBrmiNCq2O
nI5Gh6V8tIyBM6NxtCFwuPAez+6SsPOyTt0cRyVN3crvoStJbZhYIFkS1D3hEeu3
z6JfR8T4Tb57RCMqtRtXq25szESXT0Tq62z/Xl28TjvR0xqhEBB34sIozDAyXrLY
NiAQU7oaOndENEbvlBb9jN2sgM1nB0Xtpq1e5BOGdwVwgYefKmrxdninp60H+QcU
3wEAwe7f4M8U9VQwiT/y+bgpQ7U/ACbj1w718LNuQUdir9SOf4qrLumOS9EuTOM+
UUWw0fNtQ8ZvFonQu+HPfajl+c9EZtygCwC2oOfDELlMVLXMiteAOEUddHUqRsL5
5dh1XNbgOxXoamGzcpYaNZKaqrzOT3iWTYeD8ujZ+b55nZuWlVDNNP0i3aqqJ7bv
ppwQHvwe6AAJEAUakhefspkKZzprboBHyF5o0TOgiUfMzkNGeofyryerdyVZfm6V
6XAplZcV+R81qRLjzgJmV8FRFdxl6tp7GEV4W/zxAel0DvmPWJTjXNqtkxmb1LZ3
rYUCmQbKOpkAT4IZ59XQ95h0k+HjHHVBy/794ZhfnSJ7QWSul+inreV/L48mHWqw
M4tp6W0gvRldE3VSCiVr7xHnbAH2l1zbYZuRcMTl8iFwbOyvstUoyUTXfZpem5LK
o5CShq8Q00XYnXOfdOUujSWrEu+1LHxXnvFTwx3g/0/eKsAjwM1pc/Y6iwZUIqEV
P60uDOdDV8Fx4oRDFzWt+eTtPXiaNdxEVUUhfCTdsPAocHkpOu5wiRlT3S+wd+9m
v3rTToqgok37Ag92RymB4UzuWqS504408udDnToCii8m9KYCANTIiCpgkFOljTlt
gOW+bQciT/hX8wX3UFsokNwHSGnwKGOmFLnRXQ2XeZL+9NHY5U+7d17GFbzyFZD6
uksf+Vmh2x1ITiym2Va893ag+lwFAzgDWbpp3rRUlOOOS4g92K9olTgYzQJxJUP9
qhmhE8QY2pUks2fpxMMBQmKpeOogIjZ0JOjrxO9+vdbr06AaPebh37QH7L92Cs1p
asQh3tl5hub7VkSKncaPeLXhfTczKIJ6iD53NsAEqlX5NKxIzsOqHKIk1Fkp0TRI
Z8Z4F8zTNlFYx9CFZNXdkCTe7RgB1BI2ObnrdOjJROmlM5a6eggCwC7OjGsDwXpV
/hPMv1GRb8C1EPbtorvH5l7KvnCS7mZJXTPctsIkfm0R4BUxE5mYoPMICnvfJiXA
nhZ9xcWCFyfGmua63lqko1Vi3JS2fEXmf/JjYOwkQbVCH+8YTu2e5x/r9xirn/O8
R73lr0lSUud2nNUHb4Jri6O6yfuFGzHZ30htQXq8fx8hxnzdPESsBLhsDZAUvgEv
QXrnEe19nssqOoLju+9n+n3zBMwOLESiPYiMyiSgOB4zdqMXScC4osXFAMfTif41
52Q/RUbRV6egc0gKdmKcx6e61P8bo0jpFGfVPefGMR2btQmj7oM6Y7R6PpGOgovv
8Y05Ja8ckXhtvFVYCBb1vmzFEALdtZOrVuFR1u199ZL7KD6qYpNOZN2d/1OOn9Hf
n3BG4EN4+c0GltlyBEDF30+fWcFBQJaZGw7hC860EAAMoD8J/JVrwwVtU+cDBRhZ
HN8Y7tFEIiQiXUVjBsi9684qK4EcgbqgNZTvLzFzUkoVAuL0wpkvvmESqi5gshMh
qFJ/ZBHSG0Ukn9f3lmyjkuOeThmKgbZKSlhI+63Y88xaQXflkQQqt4jE07XrZ7Tm
T9Bm7ttshfcQ0ODnekABHGFLysLcKAnF4ahkH7MNjIGLayD4XJ7VqElImQccqoel
8RWADnuEOFJ4GLtTiRIVDXjmP/R/0vWRTs7RKD7A3uXTWgtLrpXoZJF20/ayV1w+
bsQRxo2Rnuc4BO/fGQp4iJjZL5+MsWKdRb8IGo1p1Dp1Sv0OKT3kgCV2kFusR9K3
uGfD3vk4FHktLwShT85Qfy6oX/EwLQZwcV7Hpk4CHMltaS0DdVYBNpnapNmFgmDG
zk2Mj815h3S9ZGT5WeEq4bMR0RtMkcbwfDWNRzfrYTFforAyNciKHwYMw3ZA5fJo
Urod/MdfPOfc5wWc3JbuySFa/44foYvg3Ti9OioL75rWdPiEbyilAR1Bowb3wLz7
GxU2H9zHBT4SuVuxAXZcjMuQ7K6d9qeVzWXj5hjspX7qjQMvISFcN13vc7gSiN+m
/R6zMqhhf8aa9WgaFrW2mw9AbF59QNGDNJetyoc0M5l4UKulGnWZxY90Th1j0Xjn
aXkkleRTK4ufQSK2hiPOeANh5W0oxCV8n5j3mtA7fwFxplNztlfDjuh6HyMJ/sNl
DY+kjOH97yhedkmY/e161qwzMkn346xilDmtuPekDFgqnIv0PKBCo7YwAmEubTgC
NKlQYXN6/wjXDSFvDi47Be6TpX2jeDcJcawO+LkPEjKPWp6xlV1avJ2K7n2/OR7f
pRX0aB2jhdDabqTbTjN7bVaa701+JpDMgq6VjRyebYjL3HRbGQM+khPf7GkQUESz
fZcqgUSXc2kNfr/TtgGrvPOLlP8gAKiKVfyJUnCPibH4eETAGgN/ZvlhKjerHiI0
B8An/4xu144TIUvy6VhBnnD0TzxbAHRcHIeDKwiscu8pdJqH9DfB/7zntbj5D1lw
1dui41UusHOIa4t/qWeJGOLSF/O7UG4JHOBFzRhMzyE3PA8Rvv1R1PS9X1i0hwXt
vn8NvpDhNQmbqW14z5PvFcAfveezDrMS+Hbk4C+RrgeMMs+6WlsBS+cxCSJSWLUX
1Ycj28mBaTuAlEOqCWzgMoOp+bIXlOP74c3EBpELWPigdluBbXUlXGyFZO2FojgB
oyWeJGdUvYx073fHhYAqOuBXen/TcTb3QxmsabVQvVtvmbYY8EWvhu7FLJhSp6UU
ke3fdf4vr2QbxOzza+R4NWKamfYfBATF1ic9Zu5zvNV2oR+8Rp5xFQDh8zsbFPOH
FJEMROxGMpJcSmiNQEQGNRs1+UgL7e+y1+UmCrs4OS3Kp02Wa0xtVqk+OJKNcxB+
3iUvHQRIj1e43xhUEJkqATo/LwOLlPfziLIAhDIMgS5dwhYh+yg6ucNx1WuAPZsB
eQ1PMF4nkBED0489OIL+JLkorrKLrE8BE58dn+nUt00tKT42HiedXfPRVaIOpLGz
SnMTfa8X9YULThHCcq0xmrqjcOFp4vX+VITr+0Algcr45iR9iXWckccjMtK7D7S7
lkkQRZ3rhxyzJkgVyYljpjUkPQhbke00fYKxcVbg0qM/rScQ8d58+PDhsIOMRdT0
LHX4zKdXsmA2/0WJYe0+8J3v1olxdNLz3deWOAv1rOHlgJECDx4gT2wDB4ibSVAK
Dh15zFikX0ucJMQlkixcO9QezyrZt9Pywwe+5qmw044UAY7gjBqKyiH+qOwwedBF
nKPkSHSIyPa7tPZKr4dFq8bw65A6jbaHoXG43DjV1TnIgukLOvBBvkS+drR+4xFh
Zxuf2U9nQHrkfyrVxXXQqbabwhkgcI99MC9+zDJaMjiel1UjmrioDuMtasFCP1iS
y0ksWh9cyLR5RRaUSi0FF5fW/+jIKkAl7MNEek40fRVpjhOo3St5SKLXG5CpAnX9
Qm7hvcvAAwMrStBxfTK1cIRAyGWkTlvUsZjIZydhf03wqyVjLTwtzKtT/VbxKKw3
AkjiVIqee0L95qxRjdTffVr8aR8Tf06tM/jBIppT/SKMTGUkUZQzf+FdPacErWfd
hbYlE7Yig29osvMyF04LcqcRAHN96rtWdIo94Y2KZWEg+14/nc8Zc/HvQ26I+wUD
406VhbaFQBpW/crz3ZD6Oyd3AEQ/N9tw0HUpvYnjOjMH/xaq1U8GYp/1B+UpP7au
Q9Uzgga8qEszOg6sRSNudwywROCUuXWuhdj95g1mr3KE5p5MzU38P/Jt+5hfDX7Z
SYWjANk5wNbJ6IMWTOD+exixiw0RtboKL5SWJMDkWAXRVyXxuSt/uXxbaSs3vRJt
LNLVQPNAEyfJJYtsp6OrL/tHHALlPO9/lVuE3u7FZLTSGQVkNtarksK/bqLXgWUx
o27WgLXuB1txJAFQoccGnkM2EBlj1EWHGUlZaY1kjy3VGH2CbxJVqoWeNaBgo8jX
7h0jmnsiE73YBQFaYg9g83ogqVlSkynMXuT+fHhjPhXuYCb1BcoCNeTaeaSku2z1
21OaBgFXaA9g4/TQ2FPJ8+MZDVBSCEeuec/av1/zfe8jspbK3gzmvXyCuftsO/rJ
QeWL+kWqu6qAkIfisqi+NJIwzt6iQ8Ab3H67hCqd6NMICxRJTjPJjR5xcJaE3WuV
BP+wVzuANQN7tx8YqYA4Q2B4gJfn0oO6Di0TMwzV0EP6UOIPqZ8H9mrbO/EZ7W15
eH7wAMmXiTrACP6LAqdoFxBTUnn638aBFJoTp7p7CQOpyTHi1z8eTXRf+MHakYDE
gvrGW/JQezRTErJiYeh/ThqnUzDw5aMxUFfubE2hWFM9+efOkKLGShvvDvFmE+Qv
m7G/vMYDJ/X7ifDyr/fnbyowDYYXf75f7KuH2clRGweds3jeqvVkXqmaFYspm5A8
9C6NrC+uTqyaDaqtUDsnbJH2IQRLNThRgZUT8xbM9foDFPwz3tuKo3+9p1zwUtXC
PEv5TxeKkdlHxQDIh2OPJSRivNbpTuEIqp8N+LQvyMn1aueP7em3VMrJ/9NXPw0w
PChxyMp2fExpI8ztDdj70il8yAe2OUDGVjkPSEW3o+rjhpGNVzrozS1lwFceSnlt
2UesAhYK2OlPxIT08VRG4OxNL/3zDvRn1lN8IGNksY6c7kG83ueiocGzohVN/FM3
FYgYWCwRGYF27kAUQJDoDnTcPlYjCQ/xb6o11XK25AUF3zub9nXKNGSz+VTNCMwx
ESwxW7arDbxi9PpE+zPYkcrfJq02v+UW+WCEBNq6pk8ygrIUNmkTyfw0bPZIXYLb
/ILplQUE/YECnhveT4tRXCSQ/nJL4YNiVShbuOX04R8iUptakW3orC7RtRjQSW13
71/tUGORlQN6RXZtTbsq6Wo55GVAEF7HV8JHYqoF8So1He7FoBSBO/lXTlVn4L7A
NZxU1nWC1OTIdkVNSrFSlbZGV4ffDlIB2Y4OCCbuZs9KHC3ISNrMdQzDNAIHtEq/
FpQSpezyJVbcsntw4hOGGfimRfu6OoMa2HAxbXH1ad2kYL8AYyQL51CIYUkILAZ3
F+gJHMLV/Z4Ojs1rkeRtVVDLiH/m8ZRGQPpKxbTi0/oSHC6gddUuRlDG2dsAZbNk
CniIUmb6Y8+1yWa9mDjmZtbqITgKM97e60RCeB1iKuJin1SwsdLz01a3BNnK95Xk
Y6fquZW7kgcM7nxYbHesshe6q5EtmwndC9LmjgfqlwJq6G7jo0Tv99CoTVDbKqAK
nG5QLy6Z+0/Tx5hJ+Cpl2rtn1pfY+q4SqHDyq5PCdXlKWMjqeaMhyGtN9eK7KIX8
M4UtD0zRnwIdSu0Etnx1oBLpVErB4p8I/9J6Eyg6kEJz6CFx8oux8jfk5EXWyz1h
ue0T+EefcC9ry9iFI/fnjJIuW8ppi6enDuP58YV46x4S7K8SU9qAoaZsY3OWI0Rp
Uwu7izYeq0S3a6YutxlkbtDIkutoVd5Yyb1RDFJdcGjqBq2RaLfWGn3bqAc5n6mt
d6LuSwyqNrgG1eRS/ED8kwONqde5h3xOeScBlkMZ54LIY8BTJOJu1uhAc+BDncEU
tqQSt1PzXWxM0vg+9uSDGCXSjQb77zh2POD1+TAYu0qTvHVU7O7EOvXy7eOOr0YI
`pragma protect end_protected
