��/  �c�9��ߝ�.��q���Kaz�
0쌿�&|�{��e繠L����i?�!����l��`��x,&����i8�}��ŋ��N���62*���n.��������vm�� 2=�n�^�}�ou:g�-�M�G�8f��g*�So���Z5��WJDR�%��9߀�����5\h[n,qb�7���
^�TF�΋q8�~��������l!��g7.�c����2&��J�W�L�S��̸+�$;P߼��(H1W:X�T�m�#<��8i�l>F�����O�Jq�Gߑڈ`q��-�?�d�_=�OA�WPt&q�8<T�.�[e�q|,bg�8����1精���>����Z� %{���Te�	�]헟�﵁�2��Wy��(�mE1\��~����Y��Y�SC�P�&�p�fѩV�$�ĶփS�kh?ҷ���$��z�e�T�$��jo1�w�2N�c�QQL\��:,c�	����*L5��(��)���`�i@]��j9 �&�R�!�!���*�\�6����9��H�&o��[4�VҲo�u����?v�^��7��Y�2ق�꺛�}��]3IE�-6זI�$�oGҎp�Ͳ�<9mi1���*b��R�A�s�� {0�q�:�+�����8O�6~�Q&�eI�m��9Cm/��ʓ�f�V�� �N�Il�N`�I��p���~ɔ�(I�����B5��}1B��PL=�b����0������G�ո�*o_]3M���:}�d���T�,���Qbi��$���ۇ�ڱ���	��Y�O7P )T7��Wp}̓������k�|�}ߡc �����|3�ͅ71�:���x������%@�.h��R$�T�F���9:IZ~��e��R�ۑ�Jk���%%�XZbxbt;>���#<�.p��`��!�2f2B�bv�&h��N3�:`���I���HDG��??{�}��?cc^����=�X�����І0��������>�=��l��`��L��������BW�����p��ku!�K(ڗ�F������T8z�J���[���u$u�y�1�#P�yq/GϢ�r��vrY�Y��OM�L�ˇk��l�e~�L�~�Iq;���@3�)�ƋV9$ŏD��Jm�3�=�=`����\'�z��ъ�L9�%w�H�F�z��b��ǔ�� ���7���}����D�F@ک`���5�����^="z��z3l4�ĳ͌�۬�ϱ��Ӈ;h=���,&L�joҤ�u��{��1�Z����`I��	�[u�����=��>��l��&�C?�8څ���*i�s�g��w<!3���4৲���\\�mN�v��H��eͱ��ֵ�ӆiw�*���$�w��7z�����Y*֓+|�M�{$.R�Pv�͢�u���n��'Y5����e�w��30C�������v�X'�4�jk��4q�A,�GR^ʫ/�}|��
��s�L�b2$ڹ�L��_��c?��D�>�q�7� �\V�c��P���\�Fu�8�5)[�Pn��E����H׀��e����4�����g�C뀇bQ�"D�c"<�J�8��,F��L�@n˫��1�#)s�R4h���\���1�UWr��DwD�h%0_-5�#w[D���T����?�'j.�_�D��J �(j�Ec]�2ig+p�p�L�/EW��jW��n�Lw�K�k�F(�[�6��!U���J���+�`��}�����͹)�z#<"s�PX!�&W-��a�$��G�]s��I��� 3�=@3!���eڰ�k��q�KZ�z��>]��.G*�"c*N�:>�$�u��#:��Y�L���24�\I�JlN�8q\R~�ĶcɏR
���#��-�~+�a��oSy�7x�ˋn�?!/�Rg�E�L
ͪ���ۭ�w�
w6֮|n�1� eٗ5igX�8M��8��Dtu��%���]�N�5x�1s�F���>A����s�� s'>%nƨ��ՒAJv�T!��)="���/J2�g������X�e=sH��`�����'�êw��}��� T�)u,���_Ĕ4����ܠ��q�mAR-�n����ԜK$�Ν��a@#��0�8� �9��}]�����(��FO�Ơ��E _4�qT���c��f���� 3O�rA���S[�8��H�O吲\�dUU�����~���\�� ��B��;�jM�iue�;�A�����B��R(_4	�����<Gǭ�)�"��7l�|2�V^�Y��ٜ(?���[���%���<��{&�W} �t�M+{ �f)���	��Pu��K���wi�.G���(�7�g��!&3��*������xł�m��,�
��'`�yk��:��J<�K	RQ�3 +��M��,j��V>ЊH?��B����}jgW5�4u/����>x��~|%��d�?f�^��T�2ե{p�_�a�H�T�1�9��V�7{q�C�8� ��#k�:5�
��!$Uz�W:H�o�Ȭ,�]vs(c�Rfe:�D�a^�|�q3�xq�%��e��gsr�� iT��8�mz?����f-�'~9�%���t�Z����k0g� �
.�ָ"�n-� /�T�I���+�\;ԕ�̮�ʠ��
T��ؠ���p���!�#_�uJ�	���kIհ�@�猇���R��qE��95)�5w�pV�_:A�(j�S�u�lm�NԌ׵���Y�����;�ìR��d�a�&s�W���]�6��L�cޮI�����j�.�_�}�l�p���M �ytw���f�&�k�����[�ޅ�Oٍi���<�AU2�A�o�Ю7��`z�{�Gi�H�@	%��� �+1��pʐ�A\	�����^�*��Xwe���1Ky �O�W>�l'�����빅e��:/�VR�<ĕ���1���z���t�I����Fģ8|�<	��T�d\'�ki*�0U������]!��N��n�z��ξb�\@��#������h�t�5��Z6��tR͐Ek��T��������t�����r������R�|drD�kO>�*�@^�;�����/�������M���g(��⏡B�^Y�o�1��팫�����p�6���?_ٿ%�����W�m�����X�G�F[cb�D�	��Y0��)��':XƶDIew�h�L��<ٿ����b橀���L����T��Ѡtf�4��H�}�Ty��Z�T=�]���H����a�=pwk��|O�[�fi�R�E�]3�E	��-�͓I�c��`�6��[���E�*r�K�n��izJ�Ҳ���[��y�5B�m:�t�����O@�c����@�Ԟ��C��*��a�+�0�'Tm��������_O��dc��_��4�jjB��6̘;]�?�
�5l��q��n&u��b����+%���V p�x����MO�Ki��pR7rK.�S�o�x��fo����o͍>�������+;�5[�ZS^�����T6G� ��Ll���F8�"s�f~E�ˉC����&r[�O��$}&��ݷ��*������~|p~�+T$�E�	���{�<l���b��x3��S�=Um���nC�9m�������[��I�Q����S��i^ j.2�'�&\�'P�K�7��^��+$A�o�k�@�l�<�)�����Hb�Ť�!r���w=��r�]�[�{f�K�n[Л/;&�r��`n_��ݨ��OJ�څ�o�Le�1<xW�PS��1Ή�#��̈́�Y�؄�S�a�Q����^���=����e���/T2^�Y���\$����HK͸��e�ĳnN�(�{��?琏#��w&�l���z�#;{����pi4���Hӎ�+	S����@FD��$L�_���nO���-���k�O��3N��sɢ��,Ⱥ�r���/\���+;	q�d$�R��@��K� �߶�O=�Q#��O��t��eaI��[�����Uf�l��]�������?ChT�j�ѮEie���<������mB/7�[�I5r&���Jڭ����zG>猹���5,
�3����&�	0ӭ^	X��J_R%*�I��f5�t� i�8uZ���︎~c�L�ny�	`~LE��d�ZJqV�N�ʨ̴]\<6���ZӪS
A����.R�.| >C��O������@>U.-&ȩy���ag�rL��o��^K&v�=h�f7��z�5_cϥ�r�O�%d
��Ӆ�#ؤK��/�۬_ad���=����M_+mi���Y[X_*���;��K�:z�ч5�����m�B��5����^��Q�D��SƂ"(g+�;�U���X�����K��6��d�H���}���6�l���i����?��{X��P�� JNZ�-���_��ًОcD�&
'�0��8��m�-�(�%@�����H���ֶ_�Ru'��f����@C?��r�n�OW���^4���� ��?�[�i����h��]�fF����{-}]�҉�=�v1�ڵ�4���ً/�"��̅3�9|����Vf�:Ts[b��� r~l��Ԁ�@�~����P�ߔ��&�o��_�+8F�����1�Y���O�wWU��{�^�`pg����a��na�<<��Ǔ��1�r"���#����q�Hk���ֹh��ߞ'����Ս��}��L𗞯��O�@X��Ҕ�l�B�� ��Gx�����Ǉ�
R!��7aTCق(�ru��
a�rX M��0;�D�M�4���/b��I�����7r�a�z�M��5��5@�P".�Zo��aM�P��g�EP-������-%�<V-^�e���֍8v�vm�k*�v��ouN�����0&���	�X��S{f�l(�ܙ�����xs۩��'��[F��r�JS�DI;lP$M Z0l��^4K1i܏����4�69���z�&	R���j�o�M���d�ij��@ͥ�/�&E}�N���$[�C��X"+Ut$)3.#,��U���*��Qf$��Zs/f$��H�m�Ql�����p}k]��|&*�+���݀>��d�#��_�����HA[�r#�&i�#�gh���S�E�� ʩ�9;�[��w�c�僭�8���I�ޕh(����@�7���1�8k�%�78tq����y�67����q���� ������SH�~�4������V�"e)�u@�V�T��TlD��ugfY��]P��M�3Zc��R�c1�/����썉�w�+
r�ќۗ���w!�A��T��IiT�ܤC��=�^�*��4��/��5�����Xb{e�EO��lh����4���0��>X�W&�i����zy�D�I̺��y�#*^��*���L����/`T��՞4�0�P�H��3��Nn}��.���꜉�@6e��З,�	���52�2n�J��d.�FWD~ۆ��OlK����PU��d(6��e���/anc@�X���	˰y�G�_ˤT�����/Z��6=��46��Z���\CunKO�a%c��GKg��P궐k.�$+�۸ز�?x;��(��B���_��Aˊsa�^x�*�g�j�8��b��b�R��K�v�"@�7�:C?z��ǽ��ݧ�\�S= ���S@�?�Jr��5]7�ከ��=v+RL=(0��>tPs�� R�J}M�dR��?F�c�/|�^��`w;�0e<!�m��3�|v�TF�R�ɬ��ʠ��sT�P���u�Uz�F�&��RU1�6�42�Ibwt���	���ч�E�jzf����I� �I�߾�t�҅�0�OW�����?���#�C�r�ffK��Op�0H�@g�91�P+䫡�]�rE��{�Q&�}����5-dP����ٹe��ݛw��. ��h=�q,A�ӎ���lאCU�7A��}��p� �]&��"���
y0�8��ɝ��8�����Z�c�7I�By��9�Z��=_+>X��T�'�R%⽅o R����s`ؓ����ܧZ)iZ���$��$K���\��?��������^ɡWm8��NB�!��(A�Y��R�h5�^���[�n��C�q�յ���m0�j^l��2S������EV;n��f�<��^�	���O%K��kH7���P:��.�(���4�NX�1n��>E�6�:6*<!R��@�f����t�wh�t\�|�{�qmt�'�p�|���#�}P�r��RyS��ŭ���ƈ���T�=X]�h0C葉	�s�{W�$y6�������};�`{�m>�2b��x��s���h*��{��P)���*Ӷ]1oU��_�-���*�A>��56�u�0��1�\|\������~	+�Y�)"f��vYR�_6��_������*g�;�3�K�߿��o��Vz��@g����e6�+6c��3ZC������:#DbS��q�7�	����L�v�B��g��
�C��= �\��	e$����
���pum���gB`2�O_�y_��H���}��,�1�9�&����e���s�bo}-\8�ɐ�qR1 ޾N�:`5U=�Mݓ���8��=]�@.w�nt
�nя+�.���S�-�m��#qjY	G�Z�Sx_ծ�l��0�	Ⱥ����=�����h�"Hu�#NE���O�?�ħ�H翾�lE� D+��cL��T[O��j'�{�K��g��"��-_�h�
�Հ?��a �$�#��^<ʝ��5�:y���s�0���� ��Z��Mk���F9���^�(P8�6������S��T
}�D�;atċ<�:�?���o�zgǏuCj�b=�~g�>�I����>�0�voujm%Y�t�^ d��p`$�t�hlE'i|sHy]c8pC{5�eE�Y�&�~�A��U��oja�#����O���J�L5ե�#H��[o��t�ޓ����+���y���*`�
"�c�4�O�n  �XG��|>�'8g�)L�� ;�<��Ym Tdy)2\w�w��A�x���R|�X����l'df��L]�y�ˬR�OrYz>o[9�c�7h
��ܵ(k_��t=4(�
��v`�Ȳ���'%��>)o�¥��qMN��t���A"Q�gU�����B��@���&�2j�?P���0�䜲�Mu���C��)�X�^�/K_篑��%ܲ��j����<V-Em�j���WG����p�cа�RmBd���h���HR�Uؤ�T�0=��Cc�Be�/M���g*W}�����ː߮�/i(��%Q�T �|Ѕ�6E5�P�\x�扙PD�j(��Ҋ�b�9�ɒ���#骝����Z'3_Ϥ,SP����'��7�Hc@�m�徎���%�����o2h�$�f��Ʀ�>�?Ͼ�ݠ�oe?`>�(�
�g�z��:�Y�J|b
H�(*&B殐u7f��I�#��c��h�n'�K�ti���=֣��w�Y�Nܔ2�4@�v�&A���׼ەJ��h'��_���J�����>e�
PB��ޯL�,'���Ǜ�7���!~�Q��Bv��r}���������ew�M9��p��@<'#+M��B-g"d-��C{��>"j�(�n�b��q��U�z!�kݗ�/�b��A5� ��$�H��kz<�k,��EAt'�;JPG���_�!i=I�+*=O}�(�jt����E��/{o�j�;|o$�Bb'馸"�=�7��5U��n0@���߹�!�%y=��3��W���Bؒ=C�H���3 ��B�q���Ptu>ˋU^��F,>���c1֡@�H߾��b��.5ƪD��)s����0R$l�]t�/�Y#c�, �'�{_���tۙZJںCuQa��,>M����@( h�x�W ��-"@;�����9�ڃڻ��i���ځp�Rbn
9HH�B��_"��%r���$4eWQ�B��Bs����2�K��� 4�N��Ӂ'��P�π��X�س�^�
�����ۢ�n��G[��u(zC�iV�{��@�d�����b��A��r.�VA��d(b	�A�`�����:����e�ڄ�d��������Q��~���ZY�����o`������A�8n�{��4���.`Kof�,���|���C/��F�FP�1�!��v-
�ܘ,�I{�������I���7���[V�Hu^�����Tv�:���p�n���Nb�#�<���O雨��4�E�4�HR�b�^�<x�d�Ped�0u�v}��S:Tc��I��
�aR�5�I��$��}����kĄ?�J�1%�����?��1�9CǴ�69C{����
�t��lJ
��m������K7Q� m��٪\�7�J�܋f�gx+�(^��6 �J�j��an
�}�F_y7ă��lj.T4�Ks�W+ ����SQ�9��2�2����CpY�Cvw�|���c��<s�+r�o����#�Y]Ga�Q�G�,�^M�e����%�b��\��J���>�'���d�6l;$�����Vk������'�Qf�v�w��f ��ʻ%�2�޵Ave�T����\/�!��"o�P�d)NC��V�W�ϟ�B�@o�8^�#��c��E8�����?]��W�/���n*�5U�2C) GG2{Sݐ"(cW&�7�������'����ki�Ħ���-����Y~�(AL�L m�k���ހ<;����#b{(H�A|�~�߯( ���Qb�3#�<A~}�I�c����iٲU���(f��"��!i|�֑�l�q�{ ��*(���i�tQY��w	5t��O�[I>)��ǽz2L��E�݀�8����_�6�{0\cQi�]�'��+�[�������@IBc����WǕ��}�`m�]�*��u�b��2�+�']����#�F�Hj����A/�Jż��H�{��y�sb&8�f�u�㱫	�6��/&�F��3��=��9���eԄ�<d@l����_­S��j+��l�R�l�����YK�����9u�_�Wp�'�>��-A�6`���R�V����O���JmD:����ۮ���z8�tZ�9�*O��8d�.R �U]7N��D)~�B	�mDϊK��g ����Qy�_����_�DEi��p�*�2*��3�b�㤠����� "��wY���C���Ac5�i�i�}&��L�J��Ft��� CGFu@"3��~4�#<�A�;���gKx�Mc��P9GDKƃ���@���zb�N���E�+qjNB�r�\6j2��)v��ș�oF��m���W䎏榓�1*xK�޻Li̕���&\�^�K����7��w�L��s��=�T�
�qI�����'�Q (��Z��iqsg�6��N!�>ypo^�&X�Z�Ǜ����9���@�nU(���tMm`����Lk5ԭ<�ڳ��~/�E�Y��ŋ��N?�wS[P��C�#dJ���_A@)�Yd�	6~�ۘ&$�O	L���а����b
�;j��͚�Н=���f����Q	P��$��7`�d������i�z�<`q$�o�6��Y�,p5"s�\t�_�����d��4w�\X�{6X�a��w��pO$O�ݦ�p�a�Q���mxq����l��m�������Hܘ.���4���>Z��UR6�̹6��L�ߖL��U��F����A�3�����Hz�b=%��'C�ҩX��*ŵ�A���@B��D�V:���B�I�R���C����Ȭ�HĂ�蝫�1d�����gEC�k(����k���?^! �6��e�6�1���!�ĥ\T�cwz0�i�~,p�Z��gZZ�l�֧��J��5n/�RkV��`_q����ݺ�Fd�=ps����ݝ���!��Cy4kU T��-�G��>^��3��%�"Ȥ����0��A��,kL�d٣wᰧ{��I���Dlf6%��V{2t��4�~�m������H�x����-��� C�y��-�W��rǲ>�b��m�l�xgM)r�@M���r����}L)�$	d��t-4����ޗ�!��ܱ�i��$��K��>ί�c}0Ӻ��?�	��m����ݹ�]�ׁO��N�^�7�ᚭO#��sݥ�]�c�XI�2u ��%�f�L-t�AKgLee�)I�ODV����%K���"��s� A U�!������_����eYG���,�����ݭ�Z!L�ȋ�N�A�u�d��͵���	R���ؚ"�Z����BDѼKɉ�T���8lfLш�ݸ��E9?� ��$zq�-a�:�-NW��m��1�D;��Q
�I��汣�^$��H�3�P�l\��*5 ϋ�����݆�7��1��X0y��F��{�Έ���B:-�)�9���˫P�F�Lm��sG�	���ڹoʮ��~�mL��Nz֢'�D��Gh�2\�0"0��m�8T�{�p�X�Ǌ"I��%g_ 3'.J���<:�*����R�q���K����}�h����F���N��m�jYs?�� ��z�ً%�Ό��!���?�w��O?s�ܩy$*��K8�l;D�ȗ�f���^����܏��\ţ������?Όӎ����Nds:����'���[���^���6Ք��WؘL�M����
!|?/���{͟Z6[�Ӹ��~�&oD���~
��<�H�
���g%�D���}�>Z�È��v��^����ƆWf%�,�����n,���%ƯI�Dq���K�,?�*��k6�l��j�/�ݕ��-���~�R�rYn�%,s��J�	Z?r���	!��q)��N~>�\��'Et�L}?��������d�g� |a�n��=A*�� {��t[�]
+�&�b�nJ�G)Nէq2|A�W�|�lٷ�~ :��En�U�"p�7
i]����@
����%'�lH��U�A/�B���a�EH�_GiJN�<����ooF��Mu�[�����4h�7�D���7ɶ��I��&Q�˖ҕ+*�i�'Ru\Jx��U!�@�v��:AMZ���ǃ�tdm�����������_#��v�J!}m�.{���l[�]�e�Ӆ��G��LFXY*n�!�4ά|pK"b��f��{:ݑ$�3��?�Yw��eT�1���Pc
y��¿q��O$㠜�鿓5E�<�be?���;e@���}<�>^�4s���U�/A��9��@C�U-��2�o7 c�P�XXqi�T�Ҡ`E�C��8zܯx�X�g��z�ny0���nƛ/��J8�F�.��e���v�&Kx�h��z��P���a]f����/f<�����8j�+�I�MQ�zsE�,�*i��
>5��c4���\f���-�[�<�w��j�eo��7����;�].�S,���stR����uu8��&uY����E>K�6y
p3<�^���"[�I�/H���%p��|̀	�&x�$��w��ڥ����P:�[��/b���6��c��U����6s��3�����/�P�N)^^ Ѹ���31��:;�0^��^;oa�j����ms�o̠���N�,-�}��)��N��ܪ�-���[��Vމ[,��w@*E,t����� ���j��G>^���7v��غ���x�kiH9��2�+���c߰��.��*J�0���w_z$0A��r��	�]�.}Z����DX��:$Ä�tnx<`|�z��؇3�;���;`�G�f(LE9�I�	�Q��BB��?x�ϗ{M��;���TrQ@o��/Aʆf�8^WCS��s0,�`8O�H>x.�����C���!^�J��=KrKa�5{ �y�c�[�ʞ���_p�����goos撎̪�s�K�G�S]�B����1uu�,Z��8��t�X�>J*�Bcd��Y�Qm�����g�����[[�l�ff3�̴W�)v;���f��
������8��_�'�ĝ�y�6���N�E]�j�D�HY�^@�M��e��T ���F���:�d�"`G�$Y�i��<�mI0�*Z������^ñp�p�W�#Z��8�Q���k��A���K�X�G�9ץ��Iα�H6�Z��3
$�&�ߎHg��қ�s%�QaD=�ǨxfrH�*0Jq;���r_~�5(2���*N���w�k��|��z��E�|����7!�b�'�xt�^��E�0���Zs����`Y5��"��{4	2s�TA�b=���=KT���k�5�����i�(ގI��ϕ!l	̒i�-7���+)8�GUY��& $�R�Q�lHD�)��kz��2��>5�����YG9�	�!sZ
�����L�Vsp:���!Yϱͱ}�47+�>�������c�z���$#���Y��:��
�q(V�$F��|�f,g)	5I,c?u�1?��Mm��&�Ak��� ��'�i��,���[��݂�'����k�B��ң�*	��?��:_���/���j�X{����w���[���͒󭮦�h��jA�#C���-��63������)�\H�m�����.�wHK�+@�&:g��\|>�4��O��p����m���8o����`�Sa������Pi�Oh�s�b��l��ԓ��xN�V8S�r-�hFݢ���u��̃���B�0���I��6���>�M��lOD��U|�RD7(�x%Ս,��0����/�N_KZ���p�.SA�5�$-]�9��%D@����7QBM1�)�D;�bE|�D�'���n�@}b�Բ� ���))�3,�V.�#��y�����Ed�J<��
������sUݕ��&��r��� ������?U�*���B�Q{?Ht���0	��B�=�ع@���I(�3<rNTJͯކ��Q����Ym=[�芣)�y</�����Wp�nq�/��4)��s��n���F�8!�#q`���6���R�K���R��A�m���`{�s�r���hZ�~T���v��Mp%�����W�|f4ћ?P��k��*���|y��X�>o4�1=����y$�ױN�K��5$0-����xbF��L�]T��ƊU��"��I	���,ѿFs/t�W�\�p�C�x1T��B�q���\��]>q7� ����/Oa��l��|,]�9%7 /���h�������S���T��3,�:��7s�z�7���D��'�������sC�����Nm��)�N|%ĆgG[�����po�j��˹��R��t�ӌ�ߡ�ԟ���)���OF�ywճ8�:w�]Y�.'b��#V�3�!��1.���`��e� �_�����e�AI��[T�2���l|FE�38���R����\�eUc|tW��ʸV7'��]SՓ�n�Tި��󞯫��!w51F��u�e?J��Iwl|����]�fs8��3�ǉ�R��/��c]�Z��%�Ob�Bk�S�죔����!7K�N����N �/��#^]���{e�z�*C�K#9Ϸ@$^��yb)�6�t���A)C�\��
w��^>�_��6�l�+��t{��;O�����<���B�'s(/�SV����ي?L,5P!�>\���<�h�Y�[Х� S sOe8IX�7�Q�5�XڭV�A�� �����"��4z>�� �J08A��i��I�$�)�[Y��J��p���$LT3Z�w��X8���t���$�K�h�|D����}���$��������S�f�F�NL���7�%�E1�<T���1�Df�FL�_T=(h�,���xS�7���M`s���Dɭ��c֗�l!��l������3u�P|>���6�����m��YI|P��a��?��/7a�����E��o��f�]az*�?��[�y� �sۛs���.dT���V�6lO��/_Ie��4��5�n��(�;�&q�����Ek|F��3 wӘay��T��e��&�tW�Q��:�ţ�A��^z�.䘋��C��������Fn�E��/#D�C[���?���F�A7�H�����G,�&�����v9 W,J�XN6)A]œ��p���r�Ӵ�,meq0ěe�	""�_���YDQ	�o�֮�+%�{WpE�VB����s�l,ۄ��Z{��)���<���ot��^,��闆�����'D��r������5R�j�����3Z���~ja����d��7��ɍL�3נ�**�*�T�5�lu�U�?����	��Z��_-��d��$���B��_�i��_{'HQ���;�y����Ǉ.,l�~����Z��ˡ@���GŒ�-Q����
R��8���>��d�9##����c�3�w,�2�lJ�2�f�5	(�*��n`_��j�i}7�1��-�J�������,%btc�~�&�C8!K^De/���ȡx��N|{��_�P~�������U�'�IŐN�B�]l۩s��DhF�@pq�W֗?a�F��4��z��K�� r˴Y&���)o�n����W�U�䪙����cB�����"_S���!�Ù9R�����$j��N	LI��n��߽�_/�=v ���� m�S�<����|:�����e8��-C+9���[��j��z�=c��w�+wvO9
�ڃ_��2�>~�è���G��;�필��S�u���u�\{ ���"u�e,]�،�7�"1h�+5*����)sg��YqC͉�__����]�3sr���Yzp�$郾z9� ��BJ��*lE����M����yӒ�B��(��D}ZJ��b��\�O��/[�:a2�\�"����6@��֣b�(�����/+�n5�����zs4��l�p*�}�`c�9����J���|s����HК C���f���Q"nߔ�S:���28�/�����.P���ho+C��?0j��T5�8H��CY�|Y��2�$W}��eu��R�[�P~ ٟ 0_n�O����������iIwR��g~�s�uߕϊ~2��pר̃���k��"Qޱ�;t�aP����i������OF!�J]9]��H~$Z)T������}Y�䭨���U��h M{�R��tm��ɒ`35J����BG���~ڻv�hBD�_�J�X���w�j�5������{��[z#2�U�js
�]�����K��i#>+-r��͸�#wO	|L�svƝC�����<9�Ө��a�iok����gh�hXy�T�F�V�GT���N�,:�M�����l'��F��{n-���լ�sQ�ϲ����UMy)V������H>P|˝��TX0zԍ�~ja'�q�Ĉ&���9��=x3
tQ�|	�>���+1�iU���i��<Gyhҍ��g.w�ڧ�+��X�fp,4�{׭{����®�o�)d�U�]+^D���U����t���C߾V5Gk���e�� �N\Tg����	������<��6�̬�c/�V����p<�����bb�%�8�zӾO���hY�c�nj�}�_��5�Cz��9x�\ IeS$F�-���'��D���^i�pNb�/c��cqB��������&�w�T�3�˻S?���B+�L0 +�l~�r�Ee�V�W���n��$�oV�2���I��4�s;)�~�J�d̀��
�k}H�W�>�$r����/΃r�������w���wi�M\��$�Q���A3��޸��>^ۥ�ϔ�l.���T_�䍣���ﴍɸ��H���K2��B%k�Q�Xu�1L�wd82km��ϐxr�X:�$`�&���6�1��>/�B�F7&�bB��9���WrE��VL������b�o�͞S.�<DIǔ��E�a��:���-���HR��~�I>��K�=%M�=E5�Ǻ�T@��)�a�)�r��Z��Z2�i)�^����j����=��0%�	Yش=D�-����і�V�:ۧ{1�Z(Y��I�fJ�|��S[��"I��Vb?��� H�G!��7�����W=�إ+���LWN�
.��%Y_5�O�XWQQYo	]����p���Vo����K
W�%*��?
�<�C�'x���M�/3���A��YCh�
%�Ql��q�^0�h��7PgL���F>��JGf�	r��GVI�o4�.d� ���O��h�����2\� ���$�;w*����a��a��͎�,u�Ǌ#�I�}����K�t^"�=��Jq}�*�1χMz��34|�ٿ(�[�p��U���v��w/*=W��g.)�-A�������%��2p�ﭟ��ؼ"c��۟�LK��W�U&��! ��;PN��y~w�%�a�S�������.:��1��/��)𚰄�E���"Ӻ�pN{����ٻ����J�m���@N��)n���	
�eB�ԁ�Γ�:��]6���V���\�-d�j��=}��!4M�J�oO�J׭ixu�˳��Bfq�q�'Jݔ�l���'k���\�
)�k��J�����('Cݮݯ:����3� D�Wr�m7��k�����g�I�b�g��[�XDBa�.]�{�Sw�g����X�iO��Y�3�6�[�<�ot���I�8.4-�jmO�ۅM_[���a�&����3�X��M0k��gl���M�έc��=��}7�ڴ�h~���H7�7R��w�Tj��TD|�Nθ2g��cC��Yְ�Q��Y���Z�D��M�������R�SR�-B�;l�M�9ff��F'��	L��7(&O����b�:0I��o�x��;SS��������h^��3�t~��O`�b�!>�ݮ�D���(��.Ddu�\kz���XX��ڞF��l�V����W����+kܲ���+��;����EZ�u6��(|�����tMM�Z�o-�j����'���S���t:g���t�1y. �Nh6�"&�¿sR�6�}�ݒ�ޤ��h������>���X�E�i|q۳�.�
��GL��&X�Ib6��ܐ��� ҹ9q݉R��h ��V�&ÔC"��y���(J�%��Φ�#Rw�z�Z,L��L)Rç�Iω)��f_��L�Lh5eb�p3�$w�W�Y�X�UyH�I)iK|�����Ll��]�&�ɔ[�q�w�`�qr�@@�d��,�m�o�t���F.@�[,��δ�9>�� O��\qF1xVRێ��԰8_N�l0a�M����ɋ�֤GZ{\���қd�kfqz�F���C  ��h��-�z��Yv>��U��*�_�ԹCr�$�Yx���ڳ~BH���L"�)��>�F-y�g��Pb�B�U��Ed�V~��.�o��+�h߾�X`�I��g��o�%�X�/E^tS������L�]"A)�f��Id۱)Zɰ�+5.��z��ە�B��0�f��*20~�į�pyVg�ܯ��nqdv\��	 �GJ��wd1R�6̸�+��"O�X���qM��1F��<�!o���:(�0S��'�+���ן��ޔ�F,��hMއm�4*�h<�z2d��-�2+�b�N��z�� `C#�1|�'A��;�W�3	-�Ƿ��ߗ���l�
�~cb�ว�m {!�M�����I���?��<&�lK֣��D����M�̑��p��>G&� ��-�r���;S�3�ق*-l��Z�7~iJYЇpH�4T4!;��z*f�'���Z�1�n�ob;#�(�'�Ĭ��iS�׃�-�QJ�t龝L��8i��Q`�` �w��ʚ���O�\�s�ǠGn��޼�L�<�6]��R�أ���G"8���:�+
�9~��7>�@�]�	��M����Q���ϩ���)hE����� �t��z]�W'HD�m�`��*_�¶����4�2bs'LL�,?x��.��^�7��
�(A�n������F ��L�����A���|X�f++��#,Y�*Vc֌������ؔ�H"j��i�j�4r�[>pF �|��	��o>V��C�c�_���5��x��W�8d�zebx�E ���,F~�}+ m�M_|d]�����
���L?����-ԩ>V�/o�7�wwBgˌ�H���p����v;âM��s��6�J]z���jxb�7��*m�7��<��m��U���k �wz�����h|A#|R"��l7�q��tN0�f�U��MX���|�z1�o���o����F��~�E<��ׅ��/�1i'r�;������_B�)��>�$�t�;9PF*yO4�D�Ӓ�|_w���}g�ࢼbȤg�wh�jn������`F+��A��[;�i�}����u^:,(X�![wI��E<�_�V��bۇ�$
?r�.fX%ݸi����h��+�2�Q�,K���P�S� �^B�ɗ��lw����N`�5�-�h��; d	��(r9YQe��`{��
(D��6���#�Q��\'e�7�m��V<���Z�<6�>3�L�>%(N�g���j糠|P	�.~ruY�C�w��'����&)��X����;�n+:R���"7Dju;�qκ�$�$�օ��駃���ӄU6�H#Ӌ�߂oYk��6��ubHbt:9�7$�$�*��m�n�������M��[��Њ_ӥ8_Z��*I�cS޷���4�q����Ñg�VLg��!�P����ͅ�o�/sZ�!#|�.��rD�ʼR�5uK��]U�t:py�XL�.�����Cm����������0$���b ���.���-N�I��~�{�G��9�S+��N'{w�䆁�� �����D���8#q-��-[ �����w��Ǳ&�������}�Z�j�?��[ܒi�zJ�������3�Rz^��r��d�߱��Z�h;����uk���`�n%�Gɚ�s�4
�"��=�� ��{�ţҰ�Dܮ��G��Q#68�V���k,Y�����B:�B�Ʊ������='�JF�{��N��L�Ja��o��b���bST��J*�\��ʨ�d�z&�P�3^�a�'�Y������H��GZewX�g�ߐhύ�\'�4=T�=ϼL����^`�����HAj/,���KeB��:�����fd3��"#��琱��g�V�l	^�.�UEA_.�3#���`}������F�����]Sˈ
��в� 1�̬W#D�
��I5B���^	�j�Y���VZl�r�6�����X'i�)Y-|��^B:Êu8%j�*�^���`~��� A���~-D'�	0�p�!a[b��:�I�U�f�$�7�k��U�s`q?Ii9M�T���I��?S�mJt Y;�*�x&����\��B��ᝤ���`��VD}S�{>4z��hWJ����S�g]E#�c��΄᮪�1���)snX9Y�lX�m� q�(��b������()��;:F�L|9}z(�=[^cȠ(x�1��<�$���%�=9X��i�_+^X�T��+���V�Nb��_5��kF��ɯ�~E�I�]S��	
N��种tB����$m�+���{я�@+f��:�-A��F����a��Ў���e�:��rP����޿�|�|�f���kС��*�H7G6@��ʢ�Oj�N�7�ڒ�g�f�v���N2(
Ӑ͇_U���˰��"鼲v؟UR�ȟ�9(X��F�  �ٺ�Q�&�};Y�T'�﫲�l�A^�F+�ш#��;�8�L
�\+��գDG��๫yÑ�bTx��]�,�Z��X�9��<�ja2Y�����,�9���fx�E�m�|��B�W�6-d��S�? Wc�ʉU��<������<���יd�CHA욵��&�H6���+D���{6��|�#~��}f@f�B��'qẢ�@o��k�$�_U�m���_$���00�Q̾evd�Y":�X��:�\�;:�?�� x-��B���?�ilH�ݗB�YD~Z���#�8�vm ~O�Sά6G8������]�5�!ˆ;��^J&A��C�l�G�o����](��su��Kr[*Y�W�3b��N�f:�3�K��nDD���$�4�B�[�������_$(�y��0l~�K��_��b����0�U<�G=�蹻����Ջ�uP��PS��1�BmU �^�PI�Ǚ&�k�a�z���V��i�t��
����=�����s!!�,�3CS�L����6ls�^��GE���1�l�m�pzU(c<�����D�(���/�x_�7�ʋ"���Ŝ��:�j�)V��K���a\��C�L+Y.�\���`@�{nB�et��}��q����^&�kuX��!NO<��P(����x�1��&u!�n�� �R����:�"����9&Fɂ-Ż�#r�%nbbKr���ri�~���L�^��e��/n���X�Ⱦ\χ*k���3���p���z��r�оhD���!�x@��j3������aœ3��A�^�=[�h0sJ(�+o�;��{��#���}�6�6�a�qŪH������tG��|��)
�Xϴ���Jƛh���,`U�(F��P�G ����!mQ�`�b	w2s��~G9�l��)��L���z��4�P�>���Eyq<t�C���L�P�N*�LVD/��7�c�	#�3��w㻉Fp|l=L��1���bKT���U�'��m�ȓ�e������q��� ����#n6t��Y������x�-¸�����ѳ�mź]
�b5�)`#*�>̣�&XR
��$�i
.V��a\k���P�	�6W ���Jc)����_Q��ڏmd�i����/#`��E�8hu؍{��α�}�w��ym?ccR"4ݔvTU,)�@��i���֦h�n+��ٮ��񟎓��݆�G*�1��Rh�t�Sb;�jxvZ=��|�;I�B�)(2����[�Q����t��#�����q�5�K����v<ճ%He,���������]��𶑅��?$	��%���t\��}���?#j��F�����6ʭK��B��m>O)� ��p����$�FT���9�0?["���W]�e>�@�%�0�Ffp���,�+���wW{�����ocD�I�o�Ha�b��J&�51�J�����O��'�L�jjwc��
[�\�.�,y��7mM����[���������*�	A�~~z��r��{do�c.�Q@y��M7Y��Tнl��rr���3�3[`�yT�]���D�Ia�<hu��s��Lt��d�N��������(�^����P0�e����I?�)�Bo�&�{(�D��j`W]9q����y/r�)BI��'.�������Q�x��M�9�"��k�>��C7�~l4�©����5O [�P�/�q��B���R��$�#����҆O��}�;o���M����Lb�fj�\�+����{!�J�
��
8���z���Ptt��l�7sQK3��]P�]��%�bI��>Q�a�,��\Cڕ��V@�-({}2f�oe7�W�������uvD�Б@�X�&��L��f��6�/�
��|�	�H�]t�8�����f�����5:3}"�c��k~��\h���p`��"��Tm�r���U���-�%���2����7���`n��ql����B�\|�>j=�;��?�����a�s]���N�:���85�M�iUשn��-�He�buR�3���%����M+�6�
�E|�N�R]�.k>Ӛ�r��:��On�_1^gE4O��!�h�z�RZ�,��Au7����U�ߟ�J�� ��-Q��TC�����`���X�T5�8��c�Cl��L" �'����r[T�jfȋ��b$��>�3Y:����k�-̡��.�O7�$��Kƌ��`:�L����"��=+��>bМ0�0l�E�9���@x��A��)�K�h�A=B���te�$]$���o� ��J��_��~i/z�dퟗ���@���q��$#yo([�\�J�w
���ү�`
�?UZ����I�?���&�]�	�ǘѬ�У������'>�q������twP��p�D����������E�y��.{��Ӈɔ,a�}�`.��MԿ�{3;ь�K#޵��Y�� ̃���G��
QE�r�^�k-:%�,	lJg���U��9a}�&����1�2���y�������C�~X�la9q%��� ���������okT�"e���z��$/oM\ع���1��GyQ�ڋk�;��m�j�w�MyDyJ�"�C����C����(&(�3���\T�,�b_P�w��j:�f
��@�x0)s|�x���*����t���K>�
��~$��G=�e��L/��ե_��j�^H"|��8���X�w@!+j�L�7�/�Aʽ����ލn/[����C_�?����5�\�!Z�����"�du�;�A���r�C E������9i��aԀϰi��+ʙ����۪�1���l�q_�Z�ldsW&5$a�U����W�à�h�1�S%7�˲h5�X{_5[}�L�����Uވ�v���U��R�ɑ��@�O+��B��"�u��u�|�9���ь���~T�FB�:�����:b��Z��qW���-ˈ.�T%'�L�(9 C��4�5'nժ�ߡ����)h����PhON�^^���ȼ�!׀yW��T�-�\����Hժ�()����zT{ط��-���0�B�fǓo0���Hj~0��MG��%�,G]�;�v:KEV���r�9�G��s�H�����/�l�޸�gg���0;�5��$�Gd ?�5!�l��N[~#�c�?:o&�rfu~��	$��O7'G�u$���i��Ri�p���f�9'�S�g?n�.8�\� ?S2�	p6v��J~�dFT'�"���\��d�L2i�s�K7
xyz%�^�A>s���9�Șt�N�.��h�bA�[iNB{2���u�h���&�f[�eXא�
T
�f���-��(�]F�p:ޣO�-^a�c!Gޥ�h���F�t�]Nge�Ϫ0ʫ�q��k�X��f	��L>��%to)�V�{ '�A��[�xOH�/ϑr~LUm�����la��U|̶GB�g�!���7A�T���l��t}��Rܥ<�0�&�@���$�/��	3qW��`�Kh;I]�}榞 ����8�tB(?�ߖ�ȯ��)��#�
P�)�F䨉%<FM��;��~r���wi�J&2��aӖ�a�N��R5�f�c�v�\��(�)��?�C��>��G�@\�� �3`i��'G���s־�ž������*K����@��Ւ�h��@#�BSH2z��jZ�rr{��#���5Tk8� �{��ZR5������Q��k�N��S��K�,�H��@G��F����B�\H��r3���CQ�!�R2۔r	D�07�Su� z�6�%#��*�F�c�YI�F3.m�T��X�M-��̓�id��&��Պ��(�B}����@�W��bG}�5�ۃ�� ��e�d�	�����Q�<Я6!k�gAa��1����U�2M綦7�����:j0���U������IG.p,tO���n�5ԬsE���;j����N�c��f$����������o��2�h�Ѯ�)��[a�b5��l�4�%�-�WK�m\(�x��U���J�� 
VW큕�1�Y�wx�߯z�]q�o�_��0N9"�Eɭ�5�q��y� �S��5>��������\�����2�'0W�Nպ
i��-<��8\�j.U�f%o�-f�c�u/��o��S���v�
8�7�}�H�9L�� đy������azM�`s��xozyE�3R	F���|Kǣ]5-gB�u�S���yϼ������!�)]�g�����~X8�ɍ��y��Lh�m���ת/A� ������1����Mv׽\1����0�u��>y{h�zV�_\���!�5�����@�ۛǋ^��v��9$�ȫ���W�1=q,���)P�8-��]>Q�5��U��Ĭd��u[�]0�S9���q=� N��`�
ܘr�q�3j|@$�@����IIckI��Pm�&;M+��r�bq;r�,:��� `���׽���,Tw+�`�m�'�x/��Xiȥ�����n������U��u�I�]�9tN�mR<q�A7�6��}���I�i3sl*#���i^D�������u���g�+ ��i%���%��������V�Q���%@,��Tv�;�Lt2�C��Ė��۟���3�x%��D���Q?���̈�Q��3j �%�U����d�;B9a25�`���SR��,���%3z.�:O(�$o��_zt�@����@s�*��ї�)k@&���̋�˫o���u|r��|[Ȍ�A���k��(������qM3c{���4�ϋ,ό �2�Ί
14�����5�,��fk^cwGw̒�"�ަ��83��n�:|t`�ȧn�pOB�Wb�H��vG9�\RAuN�#�d����HZX�5b�m\�JA�VĩV������
���V���3���$��iA�+��k�s=�zZ�}�*E�8����m-Y��-�B��Db��v���9�o�D��1����?|h�:�> ��ڟ׿&Ue��Ƅ?�37�����jf��L{-*_��#ö�����o�pGǙ�/g��	B�GXH����0����;m�� ���<7�k{�h��7���f��KE2^������[Q)�s�;�l0���i�帷��jebiz�#4#��}�=�����}���mZ�2�::��^]IW�|Zr� V�,�l�n�s�i�P�q����X���pO7�r!Pb!���+`�H3`��f�� 2��?NʀjȰ2R� ����1�Z����?�����T��kF�Ͽ��-��&O����evn�\s�q��w@jt�mJO�-_|�����ϕ]��D���"j��Y�QN�yϐ)U���4��ﷱ�5���m��#c��BV·c!��i �\8�쉲�Os�@��O�6��O�˶Z�����K� �1sV����>�ll95'��13M��i˓~1�v��P\6�'�X��ے8�ezf�� b��K�r^F���~+�;9R�y�ݝ����8(�������NA#���[k!W<3y��Xۚz��W��l/ ��1=}qr}�O��źQ�����9�H��4��!��r�������\w%E)��T���&�
�=g�Z���]���nq�]+A�$�S��H�	̹e�^�-�2?�
4�oz��?�
�P������*��Mjal0�o{�3H�����qyq#	�Z;%��4�n�Q���AGt��R.MeN�m��S^�h�j�V��uǐu�V�~��J���͜7!)��ܚ�����e��m��S��b-�D�a^zS���7�o[)AH<k����ZZL-�+ �JY��hw�!-i0́�X�r�K\G&��=#�4��,�̕�X��C�ڨf�,_���Lϊ%�7��{?�7nϯ&�R2��F�X=���}1�肙 J�뜰�����K9��Z�l��@�[�b�;z�f?���}?s��!�h��J�?9U��x$���诇��� ��lÍnq��E��g�� �!?��	N�`T`��j�=���V��g6ru	�z+my���`$����Z���WA� ���WC���~��KiҢ�@I�5����2���%��J��9dug�O �#�Z���P��w��wKM��g�Z�/�0'��X���YS�R9��FuT��� ���;w�{`5~_z/J��� ��������Y�U��@F�#�%� �&-� S�>r1�u��N4@�}��t�����%>
4�ȟwɎ.���|�칍��lSy��'�A�K��<��k��q�j�U�V3�JE�~��LaP�܋�d��A?���ƣ`���x�ղC���*Lo�~b���7[Sp�_� ��m����ֺ�eⶈ� ��]MS=����Zض.	U2�A��������2\:Yn-�3_y��Vׄ��1s!f@a4J�Qćݏ9b�4䱀�v����f���\
<��7v�O
���(v����G� �V�@K��َr+ct���(yLMg�r���d�	Ll�	*1!˅��:�Z�x~�)�� �.����YV�͎���:�	�*��Ȏ��?��*�5p��o���X����v]����J�xs&��V���|m�čt���8-L)�m�X!�<aZ��?]R`f�W�]׌<q�W�t��Eѯ�\�����Ti,�9���pZ��\��͇\ ����5S�<�;9���t���Rrd|�M�f�K�A����1��Vo)���r�ىfQ��5wW\�Â�RqY��~5Q0Y�
6�g�g-GFA�� I#[�K�92%�w�~,��bL�L�uXM��a�ܚ��wuN�X�CC	��%�'��k����y+n�w~~G�t:\<\ݕ��>ƃ�g_��=�D�D���M�d�n��Ŀjr"A�T"
�r�6�x��{�r@���6��J��`��u4�$��)��E<�mL=5�{�O�h��#��
1�v���p�2k]�L�4�!|l������d��P�B~~[����a��6N��m!e��*^\Y�f���ؚ{7Ѵ+M�t\��wJǿwD�H���^�:$ܽ��`Q�<�q�i�b�O�A���T�$��Z�(>�C1|ٶj7<d7�b�����𵡋n��or3���R̀���%�n~���i���4)�ɜ������8�*~�B45;�	��\��%�\o��Eo��6��@0f�L�?~)K�D"��f��%X¡��bR�C@�@��Ot��63�~���7Re��qcZ�ao���a�,]Ý���z�.aEC�[2�W��}&���f�B&n����[]7����?:��7�c�L}���2ȓ�L�x�cBX΂je���<P�h?�ܩL��l(�P�ݰp�{��6'o������YO\	1����f;gK&�iPX��4�-�L�n��njEJK�CN`h����j�_�N���gc��d2�LH�}��΁1��ծ@��
S�x3�y��QYZ��l�\�����<��1���;xn�G�7tV�N.dN���ݜ#�!�`�(�@/By�s����D,u''�>$����2tB��5�e&L�;Űճl`QQ��o�����f��8"�r+�yU�[�d*d^�}�]������c^�ao��5���O�b��7�����E���r�O�`��<A���b�P��@�� ՘�:@?���6���I��l�w՞��c\r�m�<��w����I��m����SEZ����Y��OV~��̲c_��L,���>pC���1e!�Svȥ�<�NҞ�z�k�U�������㚛�`]��1��U��o_&r��,���#,�/�{Kd.��e�{M��}%��`g'�	oaJ�/��֌�w��:"���٬(a�vh�������D���"�騤$�X�Z�MfO���j_�g�QA��4�/��g�1�k���I���Z����y�b���U���y(3̕���3r��!X����4��x5Q��+&}*���!��=GyQ�=L\�<@�P`[�	�w���a��!�0C08j��1�A�����u��	dVnt�;%-�#�u�TxPS^��&�J�_���қ��4����:��Q-j��@޲sd�'��O�-$�	�{���U�_��<~��6�~�O�#еw'8��5:����Ggx��T#f�l��H��[T�
o��C���W,�Ȗ��9�y�&���i��ŬS��=.��\|
@���rϸ��!�y&V�����Z�T[DM�Y�2�8� ��
�)�������v���;����."�ل���Zw�hN��A�����S�� �B!AO%	
W�'N�Vq�g�#^�t��L�t��^�ت3ΛU��z����~�G��a#�����-�i3��?Qua��i���m��6w�o; ֮{(U����K�F���Δ*�[�����6l�E�/"��(�\�
��E��SiOK�os���㞥u� c9����ٹ�'E��і"x�~[ט����F�X�.�Xw�݇�D�V����`2w}����מ@r�Ԧ����*�I�N��*��)�.�A �J���M�5"���'^:C=>#���&�n�t�Ea�S����\C�=h*(Մv ӶC�#�U����ף/p��\}�'��V��6GH o7�gTl9m��{z?}��P
/ʸ/�#����].��82�B�}�;,�o�)�-�)Tˮ8��i�@_p���ލ2��ܬ(t�;������L]�%�]�td�L��ZofG�f��>�`��Zߥ$w%ݻ�5	*�=' �-%F�(F���� ����<��j�d�+���@�~5<9P��[���k��$ïq&Ø�_�?���Vt)��eH(��IM�&����G3�# w�P�g��9'��������\���Ad�U�`_(0�aI�D��+o�w����a�
�����:���0�=;e,w����a����>hK_55�'=�'rb���c���x͆�s��y��]N��macՊr)����R0��1$� R)�� ;ZZB�\�f
�������[�����Y���d�S�r/�06\���<L'���I������>2�n���|a��m�-�~�#Ǐ������0~曐-��,�qB�CɈ��6����� �3"�3�ɗ��L��ߊ	��\A:�m� Y�c��|Ɯf�غ9*ty�w}k2�=M>�κ_G�)=\��l� ����g_����~)������s�4W�¦b�d�)2~�&,��bZ��;v�%H�eh/+��9(�Q�Ax*�r�(�HLs��q�~���M��T\�d���nY��{�"A�L%@):����A����鐙��kF~�&���g��������h�}D�\5Y��L��y����u/�1ڴ�딽j!�p{UMr���'l	�r#�s#+-L�*Ii�}I�%�f��d"����%ޙ�?��Gخ�����{;o�Gl&e,P�I����6T��IZ��>�I6��:Я���v�Y��ش�0R�����E�J7G�0�(Y���!Sڸ\�m��1Zkؑf�"��,�����)�l�z��K�O�WCJܧd�;$�c�2y/���>�K�?����������$!4���j�oƬ_��PzG����M�q�������TeN /��>���;�����`x|�H����M<S�4����!�c�>����J�m�Ţ�b�̈�iJ'��Z�5����	S<��O;���y�\����r~�pقE|wx@�}�1�U���F*j6�-�L��7�P����f��CL첱�(=�Ϝ��u�a�1���.�F��eFD�pd}S�f�橿U��Ӫ>�kiVw��
l:�&��Fd�үݻ���q��*��t
����.�9��8����8eZ�x;�R��1h砾������X�;���P1ߡ���0{�}(o-�m�۳d��\�eF���$'�$�S��p<��J����d�KM:���h�T�|��n�~t9�Vz���?=����ݣZ�E6k�� -�gf�d_7����C�gXD���H�}$a�gO)�8�)��[�߅>�h�-(��m����WP&u��z����ȡ�(������L'��qO��Bge.4�X�茲�B`NR	`n�VGoe*��\rt'�4�sA�N�p5���#�K�~h-XO�ig3��2u�k�uB�������\&R}�p*yk����B��C!�:�"IzR�fu�M���g�V��!@d\�_��/����vp��F5JeH�;���x����~}mQ�>���D5�wV�,����<xl.�;�^��('���N:�4��Mk[rSZ�|��ԇ�N�Ndp�0A�4$�JZ95���㢺ջ:&��1r�b
9����9Մ��hQ�E�/�!t��O���!h5�Ԩc��ܒ�n#�T�E@&�Ȫ��k��5��p�n�C�f���kTD8�a������j��R2vX?���,;�WjDI���E��P%�j����$z�I��A\R8�^��x2k#�i���>�{��=lX6چ�ފ���H" H�>���21�M��1͚0��JK�Z���>ȝ� &��I7i��>_��s��<y�?Uext�i�W���k�k�t*�a��� �&J�E�vr�ɳ���b�]���]ΥR	�$��y/-CU*fJ�I��
7Z��C=j��[;���������leM���_L�e+��.D��-��#��>�
f��Ma�R��w��]��iz��M������oY7�s�
m��$t�A�7��߶�*��N��A�_!�9��Tk_�6'�.���e��/^e��˖o�	)sT�\	!��D|pٽ=޽���(��{��-FIc]��l��a:Ҵ�_|��ϔ�tː�R�@�����B.ˠP�>K�V��������f�DM�O�Š+�h�1����BT�C��E	(���5���k����I ��ט�5����:�-��M�h ��sm�B�&�
^�y��<�j��cN�5�^�!sTj1�
̈v8�ѫ��].��Ƕ�9JG.�Ms=>�7i�?�I��$\w#�Qw�r�m*rԫ.�d�y�$��F,ۑR��?�D��G�~3tFܙ�Û�.N�B�~�M�*�#зM���j���+X���ŵp{��*�b����z�@*�#�֕8]�;L)���Z������q��M�*��,b9$��,K��d#���M�� �v��ڋ�w�1t8��¥ _������B��o��^�����S˄վ`k ���T댇~�	=>�OW���[qFgY���}�~�q6��k��e S��9㨬�z�ȣ3���}q�T�_�wv�"]�e�1( �������g�v��>�)4�R��ƛ(���Q���2��-�!������a�$���ܻ�Q�@h;5��x�0���?�����D�4��gN4eϘØ��?=�5��K��m�-He�V�(��d˝�ҥ�����"p2o�f��_K���r�-uc+�AMm��t!�;������E;`��`�2�_�'M�p��LJ��a(��}�6o_H�I�^��(��k�]�De$���pf�q��I���S �w "V��ʁV�� _/�n�|qn�R��I_�~+ClI�?O�D��~�Hf�sC���n�>�YV�_�4�����/���,��[o�ۥ���`σi,�X�/�|T�bʋ���W���L���6v����f�;���[�e��ލ�`��`����
~_t��a�h��Z'
�Zܦ�����'/�b4z����K�[׉����v<=��R&�u��[�G�Jec��v�|f}�(SL�0Te����^]��������p�-�Z��"��W%�ȶ�kL�(���<�f�ҬK�u�j��X6����[Jՠ�\D��OT�V�Y��E�*���/7�g�JYiU=R&M+W8z��0>G��	Y5�	-����o��F �*uª�=�k��ՖPs��71�qA�����#fʊyB��,�UߞN���ʃ{�{x�������mtՐ�=�y�-KG��a�%�.Q�Γ_n/���N���<bb\��u\%�r�w,��>��,�=���H��������J�m��b1]�3aY�Ķ�w��)��u��[O�΋��?�GN�VVC0J��DA��
�x�[�)��c����Q���b��)Nk�]2�߭��P��91����կ�	�l �ȗ�W�~Zt�	;�Cj�f��Cob�	Q�x���ro*��(&�|c�������­=�E�mk 2��\X��q����Z��i��}!��AEPGr_�óA]�P��-:��[Z4�� kF�{o ��r.W��t
	���D���F���|bP�b�;�b̀z�(�e>,��7h�Bȥ�GL��"�=g�%�F���l����|�'P�o�m}%F*�v�&署Ec�-W��7�`��x`��KC�4y5�e�h$|�<L;�(Ͼ�Np�R��"���}N���(��ي�^��p���	������@�E]Tåj�����f���b�]��K���P�fԪ��^�_���d)��98�`�[��%�5y��Ǎ��	�>k�Z����̗��j�0����Ց�1O�����
�r.E�Fsy�C���y��bL2���I��qM�x�Os٪d�͓�'HSo�be�ҝ<8�S9�8r�!�)�q*Դb������sr���o�k����X^���ӿn���T9�S�f؇�	Y_Tֹ)��o���B�`ny�݌oB�I�!S��,q'��%�6)́�û>�q^G��{��	��GNvp'�0�M�MD��n���>zҸo�Y���!g�-"�Y֫�-(�{&�"�;9�	�u��ƈ�+>J*ׯR��s�ef%.��8�aOO�/%a�Q`颏ӧ���U��������I��o�z`���iF�e4�����@L��	o�0C+�Q������\2e�/�"�y����O�:��'�Ń��Ew�E�p��p��f%̋43!$Yt{'{�o���eoO����,g�����Mk�:�z˥����h�w�k���f���岃�����ڑ��:Uq$L:&l�� ����xH����#E���>�k�����8w��1��6M��H��3C7Y,/�ڠT߆a5ʆĔ�X�p�:��tr���"�G4c�?w?I����1���I�F3rn?�^E��vv`\Y� S��]�Bz� �7�U���/�Ab_iĘ��O}�b��Y��@��e�NK���I�oQ��%�x���v��s���
�X(a�r̷���.������90��'�H`�+��;�����/.��'&Lu�$W�R5"����,���G�@H�{��#�j��-}d���p���_�F�����Y�J=���;�
qw�G>����NR���f��6��<}�Ew�n�IQ�@��I��]�v�\����J�tnW�@d]Є'�eG��k_�>Wb�yN�C�i�3P!Vx����Z�;��_���o�S6�����������0��ZA��I����y��_�ȭ)�\o�/��d�A�-������*�m-�QqAt�+��n���6����\m��ؒ��������Ci����'���?-��b�����+��T@ꢕ>�+m��Ȕ����4���	��U�ȳWȞ6�����(ټ!���]�j�5T��o���}9ֈ��t�#G7K��4px�Q�'&;ꑩ<�Z��]OS�z����M��>ed��w�?�©T^~��P��P��[�ؓ�(��%]a0$�s�wRq�pI�oU��r5`0�*'�q����TI��	z�d���)��\I��Tӝ�-y���\��6�U{��Z@޳㢑P}�.�E�E5D,��7%��>�>�r9T�m� ���v��7�T���?Ȝءmd�D��v����4ˋ�G����^�_t��Ng1��y�=$TC���\.zV �UZ0A/�sj|�x���1��ڿ�ߚ��R�#W����X�4*�����g�Q#|�}��>iF���|��UM��f՜@l/��H�����"t��0��>t[���a ���>��U�Ł�����!�w�=E�p�K
u<�_�[���=�Bk����%j������*�>w��jo(��cw+��2��3���Ȕ-Z�|�v�?��OY�D1dkw.o��O��v�2fr��y�Ml4����aj<t�]p+Ա�^!���xuxEP�!G��¬O1������]�s[�4/�
c�:�"��o�UV~s���n�{�ǙoOX`O��7�jL�S�}�������V�; � Q=�>�\8U�4�0�&�0����+X����^���9�t`|N�^���zH��P5AG&z%�,��[�q�G,��I���[E���,igN��T��s��I���6 ,;���o���6�ug�[����@��7n���FRs:���q��ǘ�/�<�%�a�0�鎧��)�A�!��?G��	�S">�����0 9��#�J�\ �%���zsj�sgM�ȎoB.�ٶh~��6/����FƯWӪ����ȟaK���%.�Y��.�C�qP��!ɨ��=�dQȳ�$/D��MI�ga���X���v��)z�'�wCtȆW��`l�8�<l�P����it�v�6t�aɳ}l��(aNi�Y��P��^���������w\�H�%��@,m������$��J;���g)x=I_�����6%��+��x��/�/f�c�!��Ϲ=��ȿ��d��PAʋ�M6Y|��vɰ�tq���A=@�qCee����^�o[�'�9Ҽ��A"	b@�3T�WN�<0��1P���slA!-�����e��`m�Td�ȉ�Hx@�:�5I)��V9�P"I������J�����9$椭��ft�2�����1l3�.�N��󧌂�hrX����J��[�X����G��K|#�Izvk��	}�T�/�E�s���$k����	���((�q �]I'�V�%e�fng{�w��vB�%�ى@>�rO˞�0pʄ�ꁉ���0�@��p�7���^k��3��|�:����<)]q����k1�]ja�ab��;�n�+/4�&HbN�ѭF��P�8#���c���'f?�$"�\m�u$�m�6�2��4�	4����L^V�s��IX���\�Q�4�oD����8��4�co�TD�'@��Nk�z0���K^&���� \S;�ڧ+�U��I%t}�`���ʪ�A��u��.>P�[ o�vG�ԕ��t�^<}�tc1�?q ,F��J���6-��������η��eu僟���v�W\o�0�e�� Ț�Q�H_�%��S�R���w+g��I�h�-'2�.L�}�V�[K:D�$�&��o.씆F�inx��ļfd��:	:�ׇ��vƾ8t��_^;����'����t1�0%fi�U4Qu�����2�G�Ek��$5J�ht1�\�]��:�Q�-K>9��G:u��9��F�����t���G� �!Ӆ�' >�7��Tк%i�e�A!�4�Ú�%c6��Ts �s�A��735��t�'
��D]�<21U�4�e�md���ej�5�5Y�p�$I�R-5M4�BQ��1����M���o�Q�0���)�à��'�S��+��߽�4���i;��{g?�_�ns���4�^�tC�`�����BT(c�)��T�Tb��n����^�8�W����:C�����vr=7t�LA���H���@��J���\�$�ա_=�%}ң�\C�Ɍ�!3��-s�%����E�-����Jm�R��h��_,\%x=Qem���'���])@����j�6��k�e�9���=ů�7܁�щx�b��[��-��N�d� ��}i=X�m�9��O0I�~�o ��t+&�*�����ע�l^ke�Vm(�(pmv�&���otIha5��:��3Oo�k�]}����6^𯳛p��ܾ,�����xV`L�=���ȳȮ��ؑ�ƣ��mV̜P�C�awz+sW���h\��d�aJ�'����G@��R'����<�Cn����z��n���.�x�<�N�Ѻ��6J��\E�4��$���p��A�������D��-JN��@b��D~��#���H��{�U{���`��/�+@���B' ���`�­]��,��
�$G6�Y]u����5!G�̶�����h{��{�a��Cw���a��[�yݳB��5t�4��֛�&�6�6~�$�������iF1�jQ{W��Iq �m��f���:�-���x�_�Hw�e4�@-�l\�&U�2JN�Z��Z9��8�P���g���������	#7��:Rt�-e�1�T2�Pl�{z��}z�.ᮺ�H�,|�Z��#�Cbi��g�2Yѥ�L���E"�%�������K�mG�}��x5I�
�2��#�f2������saǖڜ������4��S(e��tP�b��&)�|�[��f�����G(A�U=�C}��kD�� 1i0?|@�z#�d�d��C���E�'�G�x������#$��Y��朅2Z/&��^�&����������#�p�u�	���A$�,����)K̿�9���y�@=�ԯ��I=���Y76R��0_>;9��H$�����ƽE��K	i��? ���sȑ���� �2~cV��5cs,n�5Q����v��uQ\���ǧ�rC���8�'�zPb65�|H����O�FE�e�������X�(z�<>b0"��{�lmբf�?��I���<���/롦����q�pt貧&S��Q�8�&�؁`F���#�f�;���/���Vn��ac3⨵��8�/�v�I���B&0�;<h��D$�I���jO؆Ư�sˈ���;T�c� �T��߰�u��G�Q�sM���Aó�X@��ĩXo G��Ցw�^�l)
�T;@����l>n��v@��m�_��N��^sc͇����yb���R�>��3�5N�w=|�vF�I6]?ۥ��e�ڛ�55Ӯ�aRQs��Cfܔl�v�������NH͉���T٢��M�!��m~���*�L�I����3�����������!,��DK��D��b�����!ө3�W0�}ɱ����L��	a]Oٲd�@�@���ikv��~�(x����G�Aavv�?�Ne�[���x�c"�秿��l�ji[��6�e�����6(>k��ʗ�,��D]`%�v-�Bf�܋apo��fF~�ȱ�7�wGw�	��W���&=\h�b�P��NX�ȖeO��	B罌�Ҭ����/�BWJ���f���D�1���k&ݩP�}e~���	�v*ˀc/�C�J���\�0����g��ҍ��3I�|F/�J	��g��7�@�}�Ny�y|�H��[�)��Qm��Tl��N������ cS�|��!sͻ�}eii�wݲ~$�J�8e孴V��n�\��`!uE�	�ށ�t�a����Sq�▷��G�y+"B������7I�������<����3�q#�~�X��=�7��В�?���_WAr'����0:h�G���V��y��>��?��.S�\����Y=�þ���P�x��!qp��o)ݥO�������#��t:L�ja���X�螊��|�%���`�����vs���݆�t�M��:a]��|ȭ�f����\�+R'���z���0�g�>�,s$E��t=+�$@���AK뎵��W�+K��r��7g7P���_��ZkTsBjnΣ�h���>PF~�0g������\��;F� f��� <���Ұ@���s���|��ꁿi�g�,M@ s[	g}b:2��;�������%��7�Q�=`�l�!w9��G��>���,�q8T�J��y�5���$��_�
}qto�����N�r�q����G+L �`�*'Q�UB�PK֚�8g��yJR���_L-�Ǭ�����߈u�@ ���R%K��%.���G��\Q=�]��m�i��<�
�N�>��2iO����]��ߛ��G�E��� �Ӓ���zO9xC%E$��[M�>rf����:R���y��ԫ� ��H����~�3vEu~/��k�cW�� ��?�������GB��2�|�g�vSx��,������IY � O�:�����Բh�u��l��)�ZC�G�ܫ�:o��}	����F��p�����J�[�G��C����y-��� ��t�:�?�!��A�CQ��z�jl�v�}#�'nݪa1q<>{��]R7�էo��膈�g��`g���I�lu�_���2��A�ؔ]�����T��X�rز5��%�	���ox�7��R�tcht�낤��^������|z�ÌaKfF��	W�|N��q��Q�ߴ?��p�g��g�r���p}��d"�7��o�7�0�-g�=d{}w"�|�9ƎY�깗�E^�f�K���� �_��ct�0σ�v�����=�TQ=e}�,�k��YK��� �K���+(�p:�L �%����NnJSƿ֩��	_��� �����F_k�i���:���{��V���g�&�)�"��|j8�1������ԯ�Q�kvAր3�����7�*Zt�Y�sEeggB�'"�b�B|Y�dC���0��W�\z�?d+O�f�r�Zí�(z���h MY���h�����
�U:~$���W}�}�lxL��* :1�Y����r�#��h��� �'D�-����-س���'U5��4�`�J��+� Z��&�T�+��|<���93�+��=׭n��V���Jڃ�%��A�5n�n����.<j��P�.�%Ցb�b0�Fl��9e���2�ޯJY<Z�'> ң��ƀ0���sj�a�GRo�����4g���x�EEc�xwi�2��>u3oQ$���be�׆�2��ԕ9���������-�	gF<<u���]~c����0Z`�OK��@��_&�˫d�;a#Ř}&Y�r���xy� ��ջ.@��~�%K����U_&��E8��<W@��þ��M�L���nT�� ��GV�71Wܭ��BLa&��d�j����,�d���G�Ȧ���'�Ԧ�ܶ�Wޚ���!�	N�J�
���,$Dc�>f�w?�[3İ���ɳ��`�ϋ�{����U�@1wW���eoݪ����C���;���ꈛ�H=K�~4@!�V<����R�\�Z�׷�8��iL �o���r/�`u(����'����ٛd�~u����0�B���8�:��(D	6�b���f}�/ؘ�IpK�4 �����!<f{�Н��M��r�@}��5i�B�WA�q�V��v�X���5)�nN�R�5��7���j'GI���ً'�@��lG�Y8�Y�:�t
�b�ŇI/]��p��"p��5d/wM��W�#�sz]���n�du�s�v�]7����H�ʤs}0��Ab�J%�`�YV$��^�����k��M�'�`l�&�~�lfו`�+��~�@������E=<<3���[g��!$�׏m��F�U�4����]<�0���R�{X4ö�Y	ÂE�0\X�ۮ� �ٗ��j�e4Bc)W�DQ��g_��x�Z�41�d/s��j����`�5��9�#�A!|\i��"V�������M��aAq�ul�Vb"���d�흣�
<a�! @�]�ؘ��`5s�}����P{/��bG��M��l�+����<�aƘ�ZM�0\�l@\r���;��j-��o�
Uʹ8���F�W.�ڵ?��0n.w����̿�k��T�D������I�`����o��?�8/i����YYHF�U��B:�;��AY� ����B�����ٮ��c_	��>E��"�}wH�<�o�pa��˷��.ѿN7�����t�L��¼�3k�ȾO�����6��ե�����ɱ��J���4cv`�~�����	G|��j�Iu�i��Q�&��
�*	�A�7<J��tr����Dz3���>��kv��Xc*�������Μj���K�Lа��s�͉���L�q�̾]+���U��i�Z9�-�ҥ�/rnu�A�S����Y��ǧ� �01 �R��R��'0�0��.Ka
!Ws������%���c��&�PPc�x�'Rap���T�e���\����Q:�3�.E`���m&�}�h�5���u7�A4�ߔ���}�4/�:)���c��'���^�Wʾa>j�C9���LV��;)B��bw��'#���M
e��T�v�Y���s4�	FJ�P�� �i���
 �k#8�0�6�U�gm�my�T�$,�{-Bδ�����mnH#;���P���N��,��%x�JܨJQ5bFQ��|�)�Lx�L׮X�k�����иckӏ*�|7)v�����e��e�3 |��gQ���$�(VL�iԩ9u3�N�($���nc|�(����ڣ� Ҿjp��ǣ5<;���˦���X�9ԩ�8��ս*}�Eʌ�+�UhQg$̀�OV�q�;�Gz�
��U$Mϼ��@����OO�*c�E�cA��2;� �;��GD��`����s�\	�0[�p0^^�ʨ��F��eq7�0��1�;:�bbr��x�l�d��9ұ޲�!$5L�e���+i�2)0ax���d�9�^ ̮_���#��	�XH�����2d�oZN��7r��W.���������������$�;�Rǿӛ�KK�:�t��i]$m؋^�{:�M3~��B5P�a���A�KGs������>�a#��8so��iN�����L�.���Y�z.cp�:��!�0�3��4$�վUm���|L��:	�5�<�1B���q�Ȱk�DYB��ӑ��g�'!�pZ�P9��>䜶��M����~I��Lh⟝M˃�C��p�SY[�{+v;�BX��2��b��(����p��	��
�Q�{~vL�T|rM��<��8$d�:3�7�	B��
�0l,vA��*2c[[��'��R �x��lBZ����Z�!��qYC㼉k8���.$��_�(`�

�M�&��j�nL?�jvv���`'��T��mx��0͂��T�Ӹ���c��'w��I�y��e�̾Q��5 dm��ٲ�/��%8R�|�)�F��0s�(���ߔ�?�#�P�4��x~Bly.�c��Z pk#�kL�^ ���Vj�A�:����%c�x�ʆ3��������C�X�X 9�x�TQ�!ﱥg5��w��e���T��C����U�H�R1O%e�;Է��p$�DVc�ի��s�P��SDjG'l��c�7&s�.h���I�5���ڇ��@�1`g���/�泸(�~zs~�sX�k�FV;��I��k���8���:V�5�"��q��C�̢U��E��c����]n���-FMR��l^0�9��+G.�4�k�\���ҩ�Ǻ^��2-	��Ĕ&��Ss�6m��Tt����	�d,�`]�`�"����H�:��$QU/bmL8׆�������� ��/K����Ҭ�a���x�5X은�9{�ߚ�bTL���NiL0���� GͅC@������[l3Z-����l�X��B��jiTJ���qD��IA����;M��R�n�i��H�p��	w��;q3�٩�e�YS>:�S����ϟO�\0�	@|�����J��UG���y"?��!�+pD{��K�:`V=��Ϭ�V*��m�~�-�v����e�u�$oi��ؙw#/�; �tHS#�5d�^�鹖)�B-��P2�r��d��_-����Q\����$h�4�~�
ܡ��s�ݐ4i%sM�V��8S��wO�fL����[����]PV{�l���q��
g��I4���*p��Z>n��u�����rtot��I}��|w��)ac9l~��7����$D��ӿ}������H	�.�TXC$��?�ˈ+�Fw�{y0���svK����_��%�\z,j
�2�NȊl,����1s��ʹh)��t�``����kB��`s�_�H���(�n/j��2,�s�}�#$wCc��x�}���1��5(�񣁐�;Ķ�ݶq��h���9��!8��<��0�W��i r�����;p�E���@:�PC���qy�:k��х�J&�jQ;VT}��_d<��!IO'a��6��T�&�L�n���k�&#��(	pB�Ѕ���Q�a�����*�?(%iu3T{�OB�ХE�����z�ֽ����ҩ.��:� ��}��V��9��}}\t��J�&�zt=��GZ݊��g�
���P�gH7%V�TƢ1����������pW-�%��+58��6�G%�{CڐO�	]�l�6��J��4�Ի~�M�|]x,z��	�a�B����,k ݑ�v�*���Ě��w��0���
->f[��v���}��L��ow(�
����4�P0��1Gp��[���
����9_�/���t;h~G�f��ꐌ�dF�h��)
Bvlڄ�@�&g,�0I��fq�#�b`Z�����8!ϻs�3<�������	�����w�]:��Ȑ@�A���;���dMa?�\'�Fj2��#A���]A��^�[�W��i�ڜ�ܽl��d�=0�0Ӊ�1iR�ņ�ʈu��������:���^�&��ȷ�W⁁���1�*u�z��V`6"��q�𤼲���"4!gĜ�o���>���W���F�\=H�C�e�(*�\p�{�:<�%����2m&��qs��������e6��"�/���gI]A�VD�v�j}(�6c�9*�ÿ�T�4�:�N�)w�-�֎q��i�܃dh$���Q�`��6��L �d+����U
@f�P�����${���UH.��h��������'�-��}J/��cf�����tg]�&g�G��f�n�
a��a~��9���2�4���)%,a=m�ě_��WƇ�M$��[<���T��Jv'���Ŗ2Њ؟E̽ۖg��"5���ԇ��O�\.x��L�� y�7KK<Mb�H�]��6͗�*-�Aіc�˙�l:B�!$F'�V�<����c�{Uz�z��+�у�� U���)F�V7ǊS#NB�(pɯ�؛�6��.I�|ձ���_$���P��g9��+�3T$��%>gZ�\'��Y׵-��p��t���*��;Q{
;�ʚ�sK�p[��wn�UoB��@"D@^�s$����7
���.vB�����	u�ٍn�����9�'NQ*�7�F�q�XtG���)�Ld����[��*߇�έ�Z�d�~� ��@�}ʹr���
:�+ف)E��1�|&T���(�ڷs���SI�����a�	H��{6uev���o^��w˗��-��m�F4�)�p��KGWu����P�`"L�C>�����F�"�%�ؕ0�FێI{���C�����W�# 0̔��F���d޸Ь��h�tQ�FY���rԺMH�[��M�̽�O�۫J��8�dם��� �,m�����)�x���mq#���#�>��y��Xe�։�?����[�V�t�S�/i8���kk
\G�%��N/)rveä&��W�[���h�GyNece_���UgVp8c�|��^�k(�l���%9FL�7�G����X�[�~���+���R�pEכ�԰,2�D����y�u�/�ۦJp�(�yp�a;��A8�f��z�Y�"�����`S��(�kFٓ�-<�sr(-���*0]�%|�$�\iC�󀧯&���u�9�R�lL��Z#.y��q��0r��T���~bhA�Ӗ,m����o
$�FD3T�I�fGi�A]�mѷ0����Hbb�����vq��ϫke��g�����a�k8�-�Q �k�MEZ�`8�4X�Uds�D�Z��X��%�Ge��x�����˟�J@2~~�����ɥ��+p��[^i#�dkJmWV���>�)a�bgN�!��C��`��`_3qiЈ��F<�8�)6�[^Gɡ젵z�I��@�0Y 9�H�cP�yۋ$+H�s�,Ǖz<�O?������&5��I)r��&�6�{�~�.Ƈ��^���j�a��KT\�!']���|�d��C�~�@Q�b��O��W:�L	�0u��F�9sp�h��3D]J�)�7Vg`K��[_�+S�����N�q,�˓a�wr���bp]���Yi�;�پ�8�6˵���B�Y�z�Z2�� l7�6�J��T��A0���,N--��r��Pq���g���ӕ�=du����G<�7M����$S��~��M���f��zJq������U� b����û/�|����;O�kHN$��M䙏���g����+sR�ɲ�������8��̾��A"aV0
~��>����=��<;	�u���ì+�$����
�v�5�EM돿v�?���,L�q��p�xnil�Pݧ2Ә��WE���4 ��-T!������w��ۇ	�)�!YO�1�Jo��5���Ik�=+�����(���:nBk�M�Z��@�A�[��#������y���.�;��Z&N�b�b	kS��5l(��ڲ�ӦOZ3�K~1���$?x9��e��l�xXg  ��8���%��_�|��2�Ѐ�/��Љ�O�����#K�r 1%�J�qP��CJiW���e�n4��\!B�Hј��@�2������,i���\�b�;���-Ę��=�n�\H���Z�Q�̤˔�����b�����ڳ�Q��F�ͥ��'����a���hР��1C���Q�u��V�o��Z2�3���������$��n/+��eC�<CS�k���f�o���|���|v�X�xRH0�*<zVIC��w&(it?X�g^���E	��
��-W�(�Hb�zAV��8��A��M���.�y:}ٳ�/�Yi��ù8}�.�����n��t~|T��kC}��,eŖfR�Xۡ&��+kZ�z���������`;��Ḛ���5��5�H8P��Y�=v�^�B�a��N���E��Wd>.�fm�L���r����qy85�wR���o��K�Oħ@[�G9ZT��9��\6��{qP�?��4#����k�:�����65㓰�Q�wo1΋.a��V.��@54��K�%���.7�,�F�P/M'&�҈q��7N��pM�aǰl"���[6����x9�d 
R�_�[���X�&��;�;���4��;�^Y<�)�x��{�H=W��r{5��Pi���OW�����'��[j�]�9952��فP;�U!�q�\��\Y
��hXj8�D�F\#V*}��؄�϶8ఫ#w�w6"K*�
�_R��K���������o[a�1���h^J����������X>���Kٵ�"�c}��x2����(��l���t���K�J���|-K:����B��`6iW��'�h�SBez��OV��CVaz&��L����H����>0dݺ��v��yt!0i(�
>��u�=	�Rs��i�#�h9	�fݝ���$���n�����>��0���>>%P��~5���	lQ�K �̨�:�N�!-/���ާ�Zqi��b�dR��������E���wꍼ���eO�z�<:yXj����/`��)��$���.��AX6��$�[_9�	����v��J���n�ǫNl)�eY.�L��d�E�n	0����S���k�D~�A��0<+ی'�p=J���,+������JA��]�,��"}�]'mZ��S�x�A�%^Z(���-XWɚc�Ж�}q��nnނ<|Y��<)ė�9�cw��� ��<���F�:�ۺ�R��)?�{^3av�?�	۶F#�����ύ�|`4+ie�>8r�K
�9�s�8`�=,�++#Ȅ�f�߃�?���_0�&�aY� ^2_�W�1��f�v֚r\MK8�F�Y!�Bɢ�gA���lUZ���+&��P7,I*|��ϴ|;'�dV7���l��%��5;�;�(��P|֞J���������Ԗ�r�.On�(I��On�`�&Q��||��aJ�72|�����ѡӸ@:�Tn��<A�0�I�UP�혝� �j�B�����ɭ�^Sgg�-��_��\a�"�,}��lT���k^�b �!�������{O�b��!H�gYސ-��<��.#��8�]�]�sY%[?S��u��[Y̅�So��)�k��&SN陮�������=�����:�!�F�����/~�'�m^��u��b;jL0\�ė�߉��3�h}Z����0��A~��O��7��:�ڌ��2~��Kvn�>�T呅��ń��4�w9UX�`A��i�Ԑ��P���b�2a��b@Bn���@�L� RnqY�w�����mH�:��+޿������`���F[�Q�c�U�]�!t��r?[�r��\�?�T�B���1V2���2uF�wo�y�&�w�N^M"��\���!�U�Vaw�_�C�'���J�H �	6�2-�@*BJj͵��!��M\ka:����P���|��k;��%R���D�ĸ0EMx�Ga�6}*J�ŸK%0���fkqA�.�M�����_��HH���1t�*E$Ԕ.0�:�'7+��I�ח��p<A�DD�'8�&�^#���NE�1� ���+S�7BE��ʗ~@��Krt�
kx�|��+��x �n�~˷�5�������1�G�EЗH��mlC9���/��,�1?u� 	�ٖ���⠌h�=t���e�-S�S�6�W���_S��9o-ng�(V�Q�zV���+Z#rU^�ӝ����N������-a�"�7��7刘�/6�����A���VqDT̞�T��c�Y/�ni&�_��N����>���4:Ԙ�!��9&�JpO�ߏC !�v!��&ٵ���Q�鳘���َݹ�=`�#wsi�a�LkPE����	�|��n����4�:�t��}�_��wD��|%%A�p������X�R��(χ��:ua�Y�xkf�,4>)�;^ÔJB(�x���0��U�P���=���P��cr�1[�KO,5��'V���"�
K�������7ICA ��	�a�Y���e��4 O^��4�ԩH#u�3���sn�C��˰Y��Xih�~�3P���11��/��a���l@�x��{���u� �R]3`�4+����Vb=˭��.��Ue���y��=����Y	��u*lS����F�F����7�*0KI�����MA��1	䦇��M�]��0.8��?�Z*��ho��z��
	K'��W�ʭBLX%#)+��`��	�~�\3I�p��ϊ�;<c��|�����^s�t�Yj#Lh���Դ�]1n�>_ �4F~�|0� d�x���4�&�4�`��ZD�r�$�@�^�ĥ��*���r�����RfL�H�4@�:r�b3��� ��L
�9�׿W��uU�]��ֵ�5B"��v�d�Q��b9�
/��S`��9���},j�Fl�T=����
�w�Z��W-Wxl�3��'U�K���u �iy��e�-�0ZJ�ҹ��x[%ɫ�1i�?�u,"�q'�`��H�I)���5�J���Q������Y벉(�i��
Ú_�� +R��I$�o�����w��9e<� ���� Z=�@A��wk�,����4�}?�>~_`�0_�CH��T;*�. �gO�mu�ӓ�+�
���%���D��S&r���ӣ�]\
��Nj.����� H_���$gZ�XD�M�����q9���Ѐ�ğ5�����ۂ'�P�ML��X�g�Ф�7L�����t���&C=�Hd��&�^:���1�7�-}Ө�U�+)26���_I��E�̛?����TcD���f�U�t/�m<� 2�����U�Z�eSww��5�w��^po<�`&��D�{N�N�"u\�Lc�4.Se���H?��~g���M�2���wc�t�
�������6o	��.�_�ٜ���<��:���5���=�u �{�����D�����"Ԅ�����*r�X�K�����h�&)k�����V�X�یn�/ ��v��d(����^�\����U|]�A�6�]�d�V",G4G�b�=�n���Z	h�<���	�C0�������G!J�R!T���r(&a�E�Q0C �'0��`��>v������ ?��4�O|+��<~"�ϔ�z��Hn�V�Ė�v�q�^(���M�%��/p}.\�J�-\�o����Z��1vp�����+�d�������6�<縁�����;��;���[�vB<Ӭģ�ž�W	�,jjIJ��CMƐ;����-�U����k.��|�lqh�W=�����}���G�n���L̃T�D�WeuUX.��l��<!����v��%�sg]m^�(MP�!���;қ�]H�!��iz;{J�i�c�YH�XYz�d������s�O��������:�(�nF2g����},�0x+r�W��m$/jP?5-�v�9��q���&(��� �)X	�{5�Ċ�$,�`���[�3��l� )��ہ*��Q[m����\7S�l�j+xU9s6*��v��]$��s��a����C�NV���.?��.��)%����|��u��tNlt��\0�uLKV�(Z�/�2n6[
Lؑ���~3����$���7+t�"��?��/�Z|Y�B����9ƍ��3$�GFS&�T����glO��Ug
$��0WI��p�es{��ax�?j�p(o��gV�+���/�b"�p��л���t���S�S�W�m��r�'#��Z�a��r�/���^X��!��lQ�߬�|]�^6�J�1E�Ѡ(\�n�s����MK��G����'[��
O�N��gp'P��#�b^@r�t��W���+���c:�ԅ<�$b�Lwp����Oxa�� F�*hЕ=yo.����-a��]Fqs.�(-�j��#��@�Ue�����ǯ��ʦ���rB�p�T���of���+"�hA�������Vs�Gɝ�9lcy����iy��E�Q��jEP����Oj�f�hU��Ļ�EnEu\���ᛑ��,I1=�P!�t�1r�(EȐm�x�)�<��½��Pvfbj�* xM���FO�������R�4mw�����ǳn QvZ��/��]x�E�,ӕA��	�������f�+���A-��LJ\�Z�QY&�� b�Y?^͚�֜w�J��l+.�L��j��1C1,�ϖ���K�<��3hNv}s��'ZN�!��E�a�?�닁���J�(#�����&�Q����/���u-��Ftp}?A#�"M�+��_^�%����J�u=ox���/���8�NG[��9����E��e������ڏ�R�ՏQF8����5�9�Ag���Yu�s'�A^�ЈͲ.�e݃?��el)�R;z�V}\��X�+^��_7�VGd�@a�~l��MI�r,�?T�����
�D���~%2��=��H���\�s,��ZB)d��]Rؿ%��-��b�yӃg"�\��(fܢA#a���x�U���?1g��}`L/}��X�
%�R&����>���1T.*u��c_�)��
kzz�:DW���L�
��r?k�܎��#ʔ٥��<����3�p0_�ີ���q�i%C�=�j��(B��r�A|�X��$�*�H�ިt˟ȶ��/.��H��@�ű�
��y� !��0$�����nR�Ĉ�3�r��z�O���4�AHP��Ů���/-��Eq���^�'ϳ`'�������J�6��<߼Q0�'6i��o�Klҩ����H�����nb׽
������(������y3{��ÿ ���1��˹�Ԉ�&�ە��ʸ Q��g[6�C`42@zg��_S�@C���������^d�i��%t����}:�j;+5��g��1c(a��`�Ti9�n����$W�1=`v��hD����>���"���KgWA/H�K�;`�����@���]1%7݅�
����l��Z9�!&U����[���M������Ɓ_$3�����K{=|�'k�#�UO�;I�����"�mQuu84��^P]��IP]�����$�5�ʩ���lA��w.��-�7j̅%�1Q�s��1^�Bsbir��Y�OLWx����M����uā���R�e�=y�OȢ�#��c��S���r���W��iZ䈣��9�7u��u�]�X�E	h��j����p^0G<x*�k6���O�O��~|�X�r���@&[�&
6	O��N	�'���V��8�{�&�U���|��zۗ���D[��{�o)�m��(��ȳ����Zh�����cR�_^�FH���l�t,y���vCf��_" ��u�Ҷ�$Th��-p��� ay|�� �˸T���Gg�ꬌ�5؇�|��_�V��� d����� c���aV����K�v��gK~��JB����������[��.�B5�ޤ'����G���i$I�0gpX�E�b;�p;քKc��d����Š #���n�����/�y����g�!e�Gͺ/������Q�A?@
	&�U"����w�0� �YcU�B����J,Ր�9�����y�L0?[� h`��ѧ�e��y'J�e���7��U?R��gM\Y�9�f�,k������A%��}�v��2j+���H�.=�,�Q���s!��{ťP����r�!����}�U�OSd%J�6q��Q�F��C��˯������W���(d:�m�`r�1���	����J�+[�B5����(�D̐q�VZun!mJ�D{�l�B'p�Ъm&7�z�k�i���|A֭ò���l	���ћ��(�в@��{�ٕ��ZT��g�.�	R�[��Z�d����@e�)Gkx�1Z����v�ظh�i1�EPB��~�ݱLKSV�����݋��d�et���rKp�v�1����X�a(k�_�wU8�`�h��Ֆ�m��B�VGb�m�z��3{�������p,O��n9f�^�����}�|�b¶tҙ�������E���|z����&������9v%���(�ڶ
v"�>������W������[KM��S���f2!C��7�-�V>d	&���9|Z[g�i�j�)�Ԝ�~�W�W��i�E��i-��9�ò�{|M�܈��ޚk~��H2��̳Z�^�U/����T��yhn�ƅZ���O����Ũp� ���	��/TZ�;�3�l�Nl{?�(@�'�h!�:2�@����	�|J�
��pŅ+s|N��oc�!iRgzu��FVC�Ky�065�9�����h�����/}�6�H���/N�-ʬ��G����ܩ�HГ���L�}��Z���Ǭ�����C�����8�^\m���Z��F���ƕ�j|?�� ƅ�A�[�|�����.@�._�)������Q	c�)�4p�־�齥�f*2����� Jb�S�{o����Umq���\ܲ1�%�L���**�E	�ېo��䒞 �7��������IWЪV��Tu��Nͧ��J��Q�v��w�,P$��W-~����=�˛��|��;�+�P)�W�ԲS&��W��������H��sQ6W!��ݣ|�Ü+� C2�7�$;�e-��oM7V�2�c�Tr���$�<�a^���$�[�0�c�Ӻ�ۆ��iF����e�/ƅ^�\H���wJ�bCg�9.D$>����~�r
+���ä�[:�/�"d��F/;��?�v�,�o�R��ݠ:�a�\��FH|n�94n�}���0ʠ6�R�G��r��項ā*�R��V����Vi��!z����t�]�|�+SY��)��>�Gb���J�6���l ����X��T�E�I�{�
����ϖË|���`����r,�k��/���S��O}��4(:u�\���J�s�e���������z�L�C�����5��&>��L�����T䎟�	��!T=�d�o菧�kM��k"(yK���C� �gn����zG�Sƻ=��M�k�&�vǷC�0���C�ה�'��?wu�N�U�ҫo��ԧeQ}|Ǫ�7�W�UyM:ۤꥣƉ����6BM|c_q�|oI�"��i-�K<�"������d�+�����>��D�p�oưG�C5�=8��*'e�6�Y3�	�<TPB*k1B���4�W���zh%���\>Y/E�Ā�uk�A���.{
�>�
�
Gi�Br�`W ,�2����� 1d�Qй��V���gݎ�HL:B�(��:�T�CG����+��ڠ�d�E,�J��jh�Vbr��+��Q�Z��D�g�|��>�$�Sf�+^�~���0g]�cB��{�*�5�Ȝ���8�vu*|E �nՕ�O�8�b�!�ЀH�ڶ�ւ��e��ݚ�.<���a�� Qn<����ȟ�72�z�^%�q[-L�4G��I�^E� ��(�vQ?�mx�E�����ލ��J>~G�3S���g����P��2G��l�&/�~���}��]@u���y޿�pa_�0�`���7��ܮ�B�Τ�^d�XDD,��V~�a;�A�ëߕ`����c��uWg,�u��R	�����t�~�-oӞ�w�gF�9.������*����3�]1��%~v&�OQ���8�sُU��ߌC�N��si�e�CD/���f,��R������;JH��]o�!�셚����sH�:p���]�9?C4m=h�I��bP��>ս�%���}=����z �\k���v �h�~%#5ޅs��׆�C�������<����c�~�A⫤�-p���׬��������_įvRT���K�����2O�$j���.{Ѫ��Q\[P�;����3V��Q�h�9�v���Y�$�6_0m�/O�t@�2��2;�̤�i�\mX>b_������aL�`8��Ÿđ��0����(i��$}��n?�H���(Ļ���Д�a>s1����JH*2�=�&�2�*0��?��o48V[���	��+6Ze��|����ll	R�
�YR�}/g�O����C�T���Y����v��+4�o����f��HI���8���k�<|HBי[,�zt�g"�2D��pv�y�����/���z}��j��-1:.��K�>��P��\S��G>O�?��0�m�L���J�G^y\LA��ڢ��mp�za�>"(���f�l�{����B�t��oD'>O�Y�A������;�wh/,�m�#=�0�_s��K�a���#�=��ĺ+ʹ���J ��Ș�v��	=�|�֍# ,+�AB�q*y�Z$OL���f�b	�[�ek�g(��2�C0�y�CS�7� ��뫙�>����^$�d�P���V�*$�ܮ5ٓ�u|h��4y�$V|�b�z�K ��Eh��/�
?�����#:����q�``BI��0�r�|��\�+.Q���2	9Sr��_������up��^L�,���k��E�t�u�ά5����:�z���R:7�PG������YP�A�3p^���-u��'#��v?�NEx->���}����Cs��R�Ep�=����.�_�ٱiA���N�ҡ	
�[)���L��O�Ztc��zzX�v��\<�7\���Owj5u,�M�v-�m�~��%��c�^LcϬ�se%a��b7�Ǩ��OAP�9pƺ��I�1�J
!E:nu1z�f�թ׵3l�����i����z���&�N�WI�Y:��A�]Y��M|����q��ٷ +(���1��0�K�c�-��W�5���	&�kh�va���ɚ�8����#�0��{��%�@�:�\�ɴqv+˯�����~�V���<Ԃzy��A�Į��L���f_�n.�~`M5:Ҝ'0��g�vt H�+!џ9���Z�6���i��Y"�'#�䄰���l�?q�k�����MȐ��$ٜ3��}W��e�]*�h���x*v$6n���6y�o����⵪���������蕃RM���\��Ł���ϬFP��% �ƽY��
�f�CA���ia�S痹�	&a��w��� ��`�Фr�aSURkƨ'�sDx�q�����m��8�-v-��w]g0�
B$��zN�qߥ�"��qS"����'Vi�|��g�5�v<�u�)|
��'�{*x���U*}ڲm��9���+���A����u�
hRZ�j��z;�Q7.��.�ӰƉ&��c�5F�6��WYئH:O�����Ԍ6�����HeK��%��+gl� �T������r>�y��W�Ɓ���QC���C�Ṩfh��jI��q�+�a�2ʽ�mj�hҭ�4���@��6}Ǫ���O��`/�����y���zzU�,W"�e�q7k��>��}s��nm5�JX<j�JQZ���Ȗ�~��y	\����]�>㝗��������0UL��dX�P�5�D�$u�+z8�4E���K.W`t
�i��Rp}�^��7~��5'w,F�TR�J���i9�j~��f^1�H�o=�&Z�H��:�����J�������f��Ɣ��c��$��ׁ�[�Z����quE�b��H:�yf�m����-�mz���G{�%�[�GHF�]�)�6�Η���=����ا�.υ<���5L��'�QǼ@���c0�D��+�۩�ؑ�n��儀�s��{q;7��>qBq9�wB|J�oӖ�Z9ׯ�@	���Z�g�u	���:	�
�R�*5�%F�� Y���^�pbh��9�����н����oh��;�>,h�O��8���]N��d����q-�`H��J	=��8�e�k����	dl�]���E�[�4�y�b�,��%��b'�$X\��V�*�v���Mf�zQ2�N�\�h6��H�[�5��]ڤ��[�r���b�/U/{�ǵ�`�=#Ɗ������%k�P%��~�;�s�^ϒ�'!�uL�J�w����P�R/Ap���<��A�K���5!1�ty<d���/*��vI��Z$	�d)�� ���v�wl*�%�e�k��-��1Yv��Ȍ���
?�g������)Z��!������������Q�n���/ugЩ�Ǭp��:�M�W��e����t�g_��e܈����&�c�Xh�,�Ӑ��Ҭ������N����L5�]"7#8��Y��_Duu!�&8i#��fu4UT��T`�cs�7�ޭ,p0(k������F=x3ߞ��^ʴa#�^h���x��G՛X�{n�DP@��T>QX^_a9��-x����Q4�:�G�����^<t='��K�zF�gq���>�&\q�2����}R��N)�Ua���e�����sY�N���/\�z���{B�~ �G��^w���BQ���H�^�I�\C�ݬ���	@�w��g������ Z�%�x�[!�!��^
��N���p���wX�V�c��f���	>��a��;��'�����<���ۤŇ��#���1�:�>g~�K)�jm5Lښ>
1| I�U������E�#��J�P+H@��M�4�r)���UT��.LZ��^�?�YrI�Q�E�h����I��=n�ok����OSɬK���#���0�L������^39hAtc4G�-D"����ի��奈��]�C�.�����ǥ���k�嬄�p�r�V���,�붊����
$�'�=T`O�]b�D�Ŏe=�}C9B#��< �]�S~Ch����H���(q�>
�#%u˷���#�]���/�0��,�!QhyKS&0L���'+��E�z���M[�vMGB��J�[6[��������'V�Z~8�їP�컴uݶ0�_B��eD`����;�
m�=���xVC�.�?�\4�=�V�=�ԣ��yo� ������%[�E�3���t���r!>*�2�*�����{�J���������y���P%8�k��;��ģ�߇!JBDs� Ј���������;Ztk��D���Vb�yF�T#�$#=�²�{��H8št���[	~�nM�N��⬱�~�"#<�S��J�.u)b��<�+�x���\�"A�WUZ=�t �V�o9��VT��6F������i�vBk�>��G�
�=b~c)���d���e:U����͙�-��:�t���(+e���?+����V������i4��F��3��mēE���b��t�ڃ�և+
�@p�����:�9�f �E�'1�B�Л<�Z'��L��+�>�		t+^���:��'�mX�D����qZ5����w�l����4��J��5��6��i�!8�4D�����C�{�C�#?��e��oz�ݶ��î*1�����M��7�R9v`�,EKQ�/�i~;=s�˝Xv�&ΜB+��}A�p���L�1lWF��u�����/!Y�ȅ�k�4Y�;˕��Ok��tye��`R���4_�=�P5V=!�����j�Ÿ��,��߂=jU�Xc ���(��\F%b����~�\&�b��tF���2J�v�?�:��Y�IΑ���/�GP)��_5[�Ql�����Cu9�����k߼$��_u#9���÷
1^	��'�b��>���`߬�])�i���T0��j�EDRm�VҼ��8���3�V���)�'�4� �Eue�ym�m��@u#s��8�05�}��}٭l��Y࣯C�A8ʃ�YƐ���y�#�1���	qG/v���	�+P��w(3ŉc��gCQe��15��������n2���#�g��Q��������<`'�M*��s�Гrȥ��������%Ӄ�u���?��19�sA���5j�q벭����y2?���O�����G���2������,�]<4�X��.C���b�ܬ�?��°�����R����g�~�:W�.�w�*V�$K��+h]y��%yHCJwD��e_P��{b�/��/������ʌH���`��(3�x�_�ɮt��1�v�]8�~�/�i*d�M ��&T�@�l��*zau����{G0��C�~I�V���̀��x�Տ�i+�ј�52*��'�]���<� ,�h��sg�_���3�B|�OMs)�b�QQx�E<lsc~x��Nk�s�﫪�鯍19݋
D'@,�!���|�ۭ%��J����l�S�e-ߒOgyi���Z��y_�S���1�#u�Q�~{�SO*�J��|�;���2$w2g|J�?��S�0�����VAv8y�eSҎ�����|��ܪ�ИH���`�3�k ��̽��@v}�EP�>�/id�����>��U��'�l�?�R
��L�o�I����E*?ǩ[�3��j!B�f%#��[ΰ3_�L�=����TZq��4�&m/�yw�����q7i�����F)�*[݃yy��\Ƭ�)ƃ{�J(v�i#�iV���}�� ��c�~s�cd�v���&J��J��v�r�ʇ��Ȧ~8�+�>6��{ g�@��Ef�r��j���^�&Gg���r��1,C:�8�VO�ī-ux�	���铽sM�����MDjY7/��.��)�BHC����j�m���ٶ���X���=��v'��ሪSQ�Zo@F�=,3��GΔ\�0�8��[*�W��h�r�ɒ�C����o����^lh�.�%$K���Z���Qǌ#������܃��Q;N3E��E����A[�dW��P-�u�;Q�k��5L����>7p�ҏ��܆%Dt�rC�T��<�)��Ca-;�@7��w7Q�C��ί�Z���&�i�R�pJO���*�թ[e"��?� 
�=R�g���uYtU"�S4[p'���D�4n�A[����˔r�#������5�k���)"�:3V�f�gzE�ࡳ=K%��\P%����25�Z?��]���pdz��<$�s6�<�i�� $?Ca!��PT�͎���p+�ry���B,Kj�I��i�Xͤn�C1���CZ2��K��ř� X� ;�i�<nZׂ{0m��[T�za�emP���D����C�n�5FJ�x!&�mܕ�_4�F��z�&&D��\n�z�UK~G*�����)�!M�v�������"4�s�	�C�}b�EC�Gs�F�s',��4�r8�����wU
Ü�=��=ZCӺ�-������ǟ���GՑJ�jf��v>��e`f��
��j�Ođ0��05x���R,�DI2�s)�&�x��I��}��/���Z�L��6F�ӈ���+w!$ ����/a��vڿ�92f��!X �O��.���@
V7%S�'�,�Ť.���x�p�OS�2����3��T�����!�.պa��&o�RA���OVi5�?����阂��kNm0���-g]����Bk�:���G�lϘ���~���6Y�e��ڒ�q��2���,�D�0���?�� A�>5 p������{�N�,�O����̂Ah�us�Q~4��aO�	�"�(܀�Kq�7s6Z�a���kEb�!eDz�w���Y��UPo���E��4�[���Ϡ_�T�S!EL�s�f��XYC�1BE���y�}�vR	:��Kb�+�[���jZc:�������w�	�I[Z�W��/�L�%���K��JW�=u{��@M[�VJF��g%�>��{���%cL�!҆�Ѫf���2����2���D6�#@��S+����Ŝzh����a�d�.�����D�7s�T&c/�s�,$��[Z8t��蒹�KpF�gɲ�! QK:l��K��1f>�G��r���w���{3.�dX���KLv�H �;�ew%4&�`8�t���:u��<*�7�����F7�e��'$��k��A���S��y?BK�%����"E�����wؠ����#L(
t̖
D5�7�'�<Z޲��@xUM��ih<��d�9	:��Sٌ�pQmӥ+��`|���&���fW���*6���	fb@7��z�x��D���.I��W� �O��5�<[_�6���z��R8a��g��e$���~��8T*��޼q��K����o���L�Z�?�#ZPe�{���UVv�K�\L_�:����^�3��j��� =��v�Z�K���I��W��H7ӚD���t���w��!�JbX# �eyM��:��W�61���w1H�S�2q�!$Y�;E���m�S�u'�k�K+7"ot��~kN��!��t��	��Z_�C�'��#"�J�e�*㰞O�g�$�E������''e�z�D��ٜ��Tq�f����v�h���A�n��ۯ�Ҟ>�!Ã����w��8��c}Vgq�$0}�5+%���;,z�?��~IcCS�t�����|`�t넀v9��>^I)����F���;�q�Ψb���a�A��g'Y1��:S9C��z4Q]'an<�.���N�_KF���E��.�`O;\%��}�ԟ��]Z����:n��[�����UT��H>��ip>w��(/T�V|i�q$L��{�_���tU�r�8Tt�!9��nܓX%~�%;�@y��!�M��.�a�A��V�߀y��Q��.E��4��z ����&�a��m޸�-eBS������5s)+I"�%��X[/�ە��a.�+5�Q���v���"��v~�I����|ؙ�v�rO	<�48��$F$`D����:ez�'��M���<�,,G+��>P��
�<+=�Qq�^�m�8��Mޫ$�ۼ�������b_^D���W����;�0^?�ۜ.Tq�~l����t�~�4Z�/�0���Wᬬr�����el�m��T������v]��!�Z��&ASr��S�T���m%N?��@w�+�>���k:ோ����89�!oGs��tJ �Z�/DX�S����p"��	Q�JN@����_�aI��:�]Ǧtܚ Q\�lN�N��J�ۓ{\��޺�s���zUEm�D䉸���⻦M�4z4���N��s\f�T���9-�f,���\��'�&��/P�D�b	�gW���y�c5G��i�� ��$�G��֎E��f&�l� �z1X��ɭ������>Sr��`V�D�- R����c��2���\�7��j���T�^X,�}�>E��g�(�Z���;ord��͒�i��^Gb[i-�|-`���܌�\�ŕ��lf�fۇ���+�	�!6�`L�Ycc�#�ї�d�4}K���>�'�E�o.0F��\���(� �Ⱦ@�NEPc�ز��{|�w�r��!~%,3�|bsW�/D��r�}Ƅ��9�L�ZD���k	�4.���ĥ��O�S�����Έ*�@w�_����x~��6!`'(���]��CN�O@� BQ
F��=_������_�rO�e(E
�2���xz���G�Eu��tk���<4�i�_����b�zM�q���FԷ�y�����G�*��ݸ|m ��\����J-���	� �%$k�`��
����r+�q�`*v����s��ɕ1�U��q�8�D]��X.e��t�C�F;�뿛^�*/���s$8��9��˟�_$����ck5inR�����-Cxsȇ��߱��:�V.��W6|�~A��nxt�<��>Zw��6�(��\�<��O��: ����=e+���xvFmr(Gq���'(���{~<��c0v�N����OL���"��`@Y��{cNU�����kHj<S5�!�K�_4���s�̳�������(�"��"���Io�'I�_���������(5PRH1��@��-:i�w�N˺��F�Ҷ����θ��c�K��}ɐ�d.�~,(�;.���tiD�S? �#����n�S��ޒ�r�!����i��s dz��|"���t����t���S���@��������I����;�:&o��У���А��GsI��jd��vBf¦�A��ֶ
��x��I�h��/6"����Wڑ��vq�w�*�W'^���K�Fz|�+q��� b�qf��W��eӟ<��[�;��k#`�d|��*�̋�:�Iׯ�d��V�հ���9$Ij�����q��k!p�<�S��9�YJ��<R|�+{Qhcaf��*�GS	=P�o�]��P5�=/�ҋ�wq5�L�q,�#�k?�%A�0�ڂ�LKi�����ٚ��5�l{���������r^�?G�����^-t	��ԷPY����?LJ%p0P<sp̄t��׾�7ߠ$��D
2�^���-Dk^?�[�ܤ���+�,�B��0�N��\�I~}"��k\�J5O$-ż��N��U���T2gɼ|[�Ä��:�����?:����x�-�����`eM�W�df|�����'Ǟ�����#<X���[�/�α³�q{ʒ4�Ѹ�@8�3�Br/��Ocɔ[�fڣ�#�^H���^e?��$2�҈��F%)`��n��8.�k[�=}Z�B>���
����S3p��$ߟ~�����T�1�Pؚ�A��2���&�1Ɛ���e�`dR@���>3�n�瀚{w��� ^������9�p&r�j�$82˜�b`�	0H���34�U9��y�(�Y�/C7���t��2��]
�0t�p3�X��02�i3�ԍHk��n��ZN'.�<l��$����wx�c��}�9���H>NW[�;��ڻ
��:<���
:�@C@)a$�@Z���O����;t� �}�wO���U} FZOQG��g~�B����C����IB8@�g����b֟�	a�M�*ă���nV_��p�c^���@?�E�q��o�
��'�����|�A�YЩ��=�ɼ���(LJ�� ��L���p�$�����)ެ�TY͞��׳!���.��~��V�hq�z'� ���(�1N{؉H����0a�qi��_�~�_4e:�{�P�V�c?N�WE���;r�/�p7F&[P!��3�@�*�lX֗Ո�&[X���e	~	R}'	ї�2���줎2��e���'�f��ڣ�r�������'n��d'Ğ�-Rwl����o�9�[��̎�w�9&#�Uܲ�u�\�SI
���5�x����B�lϯ�=&���o͘P����|	s� ���m�����%m����d���Έ\��y`��W�%T�b#갖��ļ4�&��EFm�gf�r#Y:(���n:6u稙��KC`�w@��ʻ�t�=Ľ�L��n�{ �G�ج��v�B������L��HgD � ��:��L�ۋ�*u��D�p�P�c�H^4+P�P"
q`DAr����hh�Iuqi[� ۰�����))΄6�w
s��_���\}�q�*'ʼ�E��j���Vp���(I��V�}��x_;��Ǩ�G����=H���*�������R�^L��^�Q�%�ޛ���"%��)#uЩ6@,�a��9��a��NkNJ)�e}��#�s����:"ta�p�PF9�N�0�`�\1r���w�o�d�N�{z�k❺�7�ڜ,����#9�=������[.�̕���|B���B*������?D%����?r:-��3R}�ڛ����D!�<�5W�T�����toֲƮ�3w�p6D�u�/qPqC��i�sa 7���{�>2���I�y������cY���`u�[��F�0q�ъ��`��;J��tt��\;7��Ke�����=�ư���*�y�s>�ͅ+���NXZV9h��onu�[�;�4�3����D�~���(����%���e[���i�LVǋ�f�2��W�9ir��\.@j������8S4-��ui�`Ǡ�=�+���ϋJV��N�	��S��蔆�r��T��`��䡖`�3��N���u��HLG]�B�L�je�3�5��C͎;8}��ǀ3FZ��L-�'a�L�WU��b��t�wc�1�x0���'Dg�.��<q-�������*�օ�\���gI* 	{�ͭZ�HNq���맸(�����00�Nn,�n�A�2�2]#Au۲���J
����n��,OK�G@F%-ATr�.�з0]c���@��E[��'�`��6�Ch'��u�/[]W5"Z-��>]�7Ps�B�Vz$�1���4j�%T��c5|�)�h@�d?�4	Q�DrE��Z�&��,J��]a!>��ö_L��^��x7�t�1>X�����ذ?��79�JKL���|vn�
�&=H�j�o��[�]0�E7�Ȑ�\XM����I�y.��z�L�K��H�r ���2�Թ��S�7)a��"��f��R�g+�g�|lݧ����q�A:#�U�c$����r{�4#�ڝ�˟xI�u����m��P�N�
f@)��{�-3:�������0�
�J�����n6NWF'����@&�Z�v_�������2GTa���S��M볌���;K�T'�û�=v��M��@[Ӳ_�X�>��a:��t5qW9�ޓS5^�4G�ئ�}����o��xnf(�Y�g��Fz�#S6E��O=4���Oٷ�)��j�O%��V�I�t�l��"�_�/Ei-����Uv�;Y:jiS�X�气�dJ0�� %r�Ҩeꔧ*�>�N�z��/���@�1Z���d��ꇉn#��^�x��]�y��^�35��&���_)�܅�B�)�]�>E���"?i�{�ˑH|��1�d<�,���'$ޛU���h�n
�C�6h̑_S������s7ŋ:J-�8� �.�{�K@�4��3@"�}�c���P�7�8���V�br�0nmvŦ˲)ɦ�bD����5z3r$CU,�D�W�N�F�"*z'��.
�Ԝ�**-ޔ��"��I_Pq��u��4�����z����Q�� � ��á�оt��/�<�8������&���!��5�Df�)t�>}�L{7W�?Ek��Lkx�֪�.a.�/�$@Ǭ�"`��������B�٨;%�f�VJ;Z}r�	��dK�qX�K3R��$�	

p/�mC�I�6���,�ȵ�-���e���r�nM�k{���o�3��(��R(I	�d}����l���S�G8�F�oj6�ڃ����8t>D]�8:�G����+9Tl��%J�Ũ5�	_��J_:-��}�1�R\h����������+;�qI=�>�pl�O�:�_+�b7^���(8������{#I6TO��(]�E�?���&�Wt��g��|�G�
��1��E�z ��
ǯ���w'T澪*��D`��:��w�
��u���hc�S�-fɈB,Dh*���Cս��ؤSߌ�sp׿���+�
��&2@v-��jNK��͘
��f�n�ULj�I?C�8�\'�d"p� ��f�M����q4�s�̈�5����.��{!1��5r�XkP���>�� ���A���-7�A��:����� ��c.��~�x�1!A��j��8�����co���]��sq�k�c$���Ǌidc��
��%�����qj+������ߔ����l�P�TU?�?�m��1��Ei�:-����)�9˾�1� �_ngL	����zf_S?����Iy�M1cc_���=L>J6{�,v#�z&��������;av��`k{�kJz7��s�.�����f�H^Gݜy2����/��k<ճ�&��X��.۸�NƲb��L,%{�M������C����MO̠���q��B7�ǹF.�H�)o�n��b�Xz"m��ރ� �4;Q�.�y�g�e8 ���K���f�s2Sn^q��*�
;�n:p0KZE	��o��wW`ÝM<�T mx+�(�a����@�t�G\{-��U 
�*-U���z�� ������7=���.�SI��I�y{O�o�g��c��F'7r�g�ӡ=3 �$j1�}k���2u��47z�:�5�P�u:ԑ�����&�bD<ދ [�M�qos<�t0�_ �`#�x*�P���f�*N���]��S��u���[��$����č�\vI�$m��ܓxM��/�M�ԣ���i)=�+%�Y�6@7I��m7�3���f��Ik�͂�6���uy�m�`��H���D(��g�"�+S�y;tO���ƉHTf)���d�xE4(޵|�Q���`q�ܐT˂f��J[���|�&$o�R_P�1AXY��,:�x��R����W�ӒV{�"7<��|���'�m0-i�y!sDLX3�1�;S7`F�7G��5�z�[�����O0�O$4���&��Y��0'@��Y�i����;Ynɱp���(�(��X%��4�/��FX����߲��Nvţ��]n��T���t��s���&{$w�i�g�������e����s��l:���'E,?	�Hd�*@���:���v,�PB�V%f��	kR����z�#�9��^BK��ap�e<�B]f�U���w�>V��ˁj�Vdb	�̎66���m���c��A-5!C�%�}����˰�v+[%ǋe~�h�34��FD�I�����8���Fh}�E�t5�Kćr��I���2|�dK���h�P�᥀L�>��hK*�ܮg_�B%�00��6v�ti��4�ᚥ �8���,�(�+��υ���i���yjڌ	J�F�{l���=�X	�'���3
����A��dש�-���{�Zy��UJ1o�. ���YI�.%� ����6�^��ΐ�>:o;�^�R�B��
 h��
N�j��V֪�)�'.J��;��i�5�)��|eJ�(*��� U�a�S>I9������%������w�V~9|
���ya��E���%۵nT=�:¸�d���h�l�(���	������Z$nY�������Bv�@��S��w���O^d����:b�6�"G�@s
�1Sޘm|{�^��		c��8�7��r�1��|e�����������Sv俎8J��#���r��v���PӀ�{(�=�Ē|Z�	�����X�w�d�d��f^9�Q�Lr��:����	�~�bݭǿj�%)����k2饵�����iD�:>��ME���*4�u�V�r]Ou�����UרT��Uግz������hL5-<��Rq| ma��n�Fn�Լ3��/y�!�Ģ"�{=�LHA=8bn{xQ-6s���z7��l|�$/��%;��{�hq��ϐ��"�gjsA@Ĭ�@�^��zA�3����q���1�������u��<+/?��+�q�5&�������j��+��c�TT�v->���S�.w+���5��%�Ak0_w��̿��MGYҴ~��jݠ�u"��z��t��C��ԏ��<�\������{[�)�ޗe�<��&���X|��cRk�I�U�� �ۘ[���ܕP�{f���u�m�?�� �G������p��F�N�������B�೔��(��c˻���
[����(R���>K�ve!��!����S�8N�C��?m΄9#!�X�&/�N�y��"��`&H��'�$6�4���aPc�&7_�V����m���t+�>$�M5�C��H`SgUN�\h�UU�U|#���8SQ�)�(��c���&o�	�г\��S$F�-�Xrg>ғ]����Xv��Z)�Mn:�4�.�f��,��������W�_ ���p/�g�D��ir�K"3������0����%:7o���+��5s�.V��e��(D"�j�6#�t�e�v�F~EW�L�Ӎl�^4I��sƵ���2y�������Ҟ���9�P]�)�7��7*�{���٘� �i�y�k�c�u�%��ֈ����Pؽ�0����`QX�wb/f��#b�/�)��%XQ��{!�U�^�Y��'&`ǕDl���$@WYQ]�kX�/!z�B�$fGcK�74a�t9Rm�����6�O��؛���URD@iI�҅�yB�v��~}�ښ�+mR��EgF�mj�^倣�L�o�OO�틸��b���(���xAշ�������9G�*.���{�=%�ɘ�k��蒃q���?��)%��\�����'��'ium�����$�"O�N���Dm=7���M�RLF���ŷ�&� �}=x܂0+n�7H��x+���Y�B� �W�_��^�PuA�ͤ������ro�-pR�V�Ǳǖ�i=:7x�$�~���� ĺ��%>]�{�Ѩ�X7��t�f7K����<�������fW�j�/�e7��b��alb��1�͚�b%,��V�ڽ��!lg����2�9��Q1Q�gk*WĎa=���p���xn��
!Q΃\�z���Jp�
H�=�O����LG�*y橔�4�ő9J��ʷw��D�T����ZZ��G�_��s���y��G=�����_n�7h[M.�{�(Vc�T��/����ׄ���^��G-���4cʫ�9/KO`�%�0�n�>�O7�*Jv�g�|��Bp�:&ݫ�[�fRĉ4RV����%W׺��ו��c�@k�]=�V=���/N@�D�&_F���r�<���-�G�V;�Zw!%�MZE��.����:���$�Ƴ�ݘ:�����{�ݛÂ>�n�q
�|���rp�� yI�0�ȼ�BRA�o/�xT$o��5ڶ�i���PKW\%P��� �|"��T��t�רoT�U�2PN���^�M�iiݤ?b65k��e�&-�x9�e<�Q�_|#�H�=���U�+ɜk~��7�~¶��Y�2�>픝����+�\7I���b�S��|E@� r����ġN�W *	��n+�n>�5.��/��ۊU�<�gZ�l�Q�*�`\ΞO�z�A���Ļ{��&Kk�6q\z���	 ޙ2�nnXa�6+���["q�����2�( <����[�������_�*];;{ #��,�ݐ7�*���JV*!뒹��I�`B�W"4j@C
63HL7�s��ۧ#�����֕s���p��m׈���:�*�:�q�E�1¨iuok���\��^2����|S���Z9�w�E[��b��BD��@��'�*<����^P%oƖ�3G͹\iv5�5T�[p���,�RSi��ԕ�Un)�1��gəU�Inw.=l��� 0M�٘��6��Z6Ӵ����V�����*Z��bw�ގy�5��ⵤ����*y1�F��O�&Q�b�̃�g��{ai�x	���3�����=8�
rm���]��%ۮ`�/8Hv��=��O�/#����{���S����T<�F��&����Em+m��sRq�y�M��o��C�z���s��`�"��:MD8�bH�r�ݕ���>N"]��6�ˬ�O���^����W�:���1T���dG7�G��o�
��h��x��*31���N�i<���t�Qn|Q� z�՗��l����s3�(��ԅ�:��l�Wm�9�<�l��P}E����JV��=�?�N)�A�rV�-�ґ̟D����JЁ��n�01�m7���90�h���4�0r��g�#�[��2R	�v�4�b̐zo�Eo	a@�ͯ��'��sJB�x��T,-�15%�}_��/c(�$�T@����M=�@a��6:F��T�iժ��S���B~��M�ɞ��l��h�bW8�D�A=��(R�*�]�{7N��E�s{�O	��vGդo�wl���۔E�G�~�$����G��/�x����]x�a����:��/O,7��(Be��!|o�!W/�k������p�#2q�V�dN-"r�"�	A�8_��S��(�0��v� ���D�m� F,dܿ�!l����U�DFӏк%���D>����R��h=���M?�d�5 7�^���LD�i�}+#|�W����`�$ oIg�'�u	�SyS["�ܛ��xB��*����k*ֻ������SM>��!��3bBp�&�7~�t+S���&����7�+��c�^{��S���|���r-Y�\VR�U�4�2X��fN�Ip��kz�Ѷ 0��wx��sV뜠�l��݆Lր�q\��Xd�e��������	��7��A2�6-�}�A���Q��x�RD�<�����G��`� ���_�C�r��j������A�);	�q�r��C���"1f�:�5��ֶ�-_ɷI6�"<��`�k[L�k�5�$����H`������1 }��4I��'��koa����-�!M|�+���9#.yV�����a�d�kqB����}�ygJ�{,�'��\*ؖ��T�@�F5⭖�S0��D<�zD��Ο��VH�� v�@� ��ADV#$��a�ڹ�Z	�2�]\Hx =_�z��CZ��NM��t��<'C&��R����G�Y�����9O�нb���u�K�[�޹H�v\��s���.�C�hlZZ��<�u�[��I�Ӿn�BV��<��b�kP�s��*�����fJHa�cN�H�-`��Z4�O+�e��m�x���Eڐ�p�FXyH��Of]��}��Q?>�{O`�s]|+��[I�f���U)6�.EA��O���<�u����M�+{ ۇu�<�tor��[�Φ�Xϑ�Ғ�J6�ͩI�f�����^
��CS2�F���RJAfQ����;�ieG�V.-{j� �`�M���ud�ľ�h�	T��FO?�{G����j�m���e+9=�ua<áN�M'f��]��#�	���%#w8ӕٸ�DW)�F�u�M6	���#/hJu,]a�A��_�N�� ~��CUT�����an?�x�@�a��Vs��:�-�QK\7׾A�.�$Ք�fb���$bT�K�t���g�
E�o�t��%~��|#e����@7<�2z��R��Ԣ��_���.�c@m�����zw�^Ȩ�|b��;��Pv��\�a��s�`Q�iz�����Z�Ӟ��Z���R�W&�`�9�N��4U����w�#=�doKh)+��3j���({o;��ܽOl��ҿ��(wg�7���ӻl⩁��P""����~9ܔ'�A�"U0:��%�;?8ղ�#��nh%�юd�ʀՍ= H����d��w�(*��l4�\�p�o�r �vT{1�'�;���,�hY��|w�_|�`���b+�z-�L����O���!�����~��	g�S d̂)F�K{���@�\K��C���0�K47dN^#�3Qw~��W���۞�2�|�[�E�g�L?��\k����g ����m�3o�fD�i�0-�U���oLO�����](���q����3�`r��.~�ozb�zר�_�4���� !�
��M�O�_�`�r�LN1eDZ�,��1�X�é�˅�x-�I�W�s�r�$@i���
�W</<��	4��T|�A�|?֟줽J(ޘ�M�H�1����L�t#k�
SO��T�󳚵t��_��Ot ������Z�d�<�5]r�a����M�DS煸)m��ᨨ^�8�n.����N80�g��A	��Z"�w9:�~�@d���c���l1��"�����`�3���Yvu�S]f]���O���@Zb�m�2�;d�d�b�NU��ն�H���Z�A�e�#>l��A��`Cu(\XQ�\��'����[�Au�Dk7��򆞞�E	y9f���n��
�=N^���������?�)z���	�B�]|��Y���Fv�%v���3�P�������ܺ��"&W�q��E|$��%��~l�1c~���W���q��K%����W���҆���{�z�G�)����YCz~��];i�-=��5#�8-�����n^�/4o�T9�(�n(��|�n�O+��;[*���˟�ȟL��?���_F�S�� ����0 ����
8wCKG3���;�4�j�dv|X*]��,l�U&B�*
����se�u�����#7�=���wC/fL�zl������t+Bŵ��]sU���&�03x@�E��<��u^V�s�v��P)F���~yH?A<0{�l�;H��D��<��=%7Ԋ�s1Nr�+�
m�UD�Zi��t���QNrsR�I�'�ûTy5e�G'~A���ӳ��x?5�H�b����!䥨˷�DS���ҍ9���:��<�����i�pl�����]&��a���I!�T�4��b�Y��B7�5�/�3n��1�A�����Z��E \���hE��?&ߌ��M���]�A�h�N��Ӳ���0���A[؈Ề�7��R��Mcr[ITY�_����u���/e�̴�5�pa���	��ͨo�u��-�����ꑹK :�.}x�'Bև��+�|�'F,eZ��w��t���bq;�]��D��@�f��sj�4E_}��;��ķ��%�6�עD�َ#WO��phm+��e
5���w���MYnI:sTJd��d��TUY�A6�s�LG5%�uL�����l����Lsh	�'W�xYLK�_7�?�� �Nv�v��^Pƀ/����hs�#��"A+����B�IMJPV���[�4���.3����.�|H]d4f]@�WV&q��r4�24J�u��Q���R��=17k|��(f=t-�w���f�1VGd)�Mdy``q��[��=pb����ZEИɖ����]���1�'��� �@4q(�@���=�&�@	�t�������̦�8�,b(w�0�BZ�|�k�����WZJ�{�3��KP(hh9S�<Ej/H��u�Ǌs CA�V�~hY�7$�Lc�D���4��m��L#ٍ}�Ml�{dj����$�_��q����׎�K6]҃si1�/i��6@@&`j�ح1� �1��rt��M�CHd52/�f>�.��0�Z����i�8���}��5��;�n�Bp�]���!���k��L+�:?�ܒZ�v�`w�j�!}�4f��g�&SWL�����}���p|���8�Kw܌k�:�$�U�8�M�s g�.^���"�T��O3Fz�͗W��^��_Y���%�qI�d��K�q��
��Wg\VRP��zLG#o�;q�go��T�C:��R�pb6����� ĺ�h���~�f�a�ޢ�ó?/)|(L������T�[��X�H��h��1"��z!�[�t�a9g���&-�N��ڌh$�A����G��D����ö���'3��D��Δ���GqS"��
f���6F곂�����I�W^/5&��c��!����<�b��V	���P+�#D�2k+�����?�ztع*.���62�	�|��?f}Z�ر�P����К�;C��Գp!���ݙ�@�,aye�J� ��[)І�9��p�����3�g1c�D}�55�.vH�UД_6O*�QZ�x|M��m�=��"��F�?,�P	;��WP���&��k>���C_���}�A�o��C�P��}O�������e�v\��ɭ�_\x�I�,PN!��Q�Y!��}���"]\ш1�Kh�Ϝ !0&���3_���x.qu͎a�.yu5|�0�/������N`Zo�O�o�8in]AqF\����޹���f�KS���G7嵻�d�� 3��Au�t��4�{Nl�S*gZ�<DBRHR���D��o[e�b�!NΫ$��Z0!9<V: �ܞ�����d_���"�4�e��!;Gg���?��3�3�J"LG:�	p��Bˮ����?A]�	�f/�ǉtÍ�u�Г�p���/�)�b���w/�-�]�Nǟ���B�/��\�� N@:y��\K��ʵ?Qʢ�B�4U������I��w�eѴ����DAQ+�`��R��(�9-��궶M�:�#����Qx�4�tS?%��� ���7WLyJ(�E�f}���\?�P�"χ�!ڈ��U�8��_�������tV�є�M����2��F��gի�5���`����%�7�
7�8�mr�rX�F��"W�4[���Ϲ!c��\IZ�:{�4'O/!*q��a�Z��Ϲ�"����@�Ȯ�G*�H�>Tu�
�=Ex���x���0%d"ߓ��x�^03�2�H�����7C�0���N%hNR}��W�UP�������	���Q1��JtZ�w�z2�]�P��ER5�#�K�G�D��N���1�kTMu8�)�B1��sR�/5uA�m���B�ղP�S���@�� 
���k���:�h�xpΡsK�H�%\<q����s��;-Qe����]��p�5�r�q���=;�M�X�M�/,���y5�Kh5O�I���)Z�s��
Q�V*a�>��/2ܼJ7"��t�nx�N�X�wu�����S2����`�k nLyt�V���H�x�MI�<wϖgN�Pl��{x~=^e.qt%NV���PM�E��Jԯ� ���s_v'�lJ�?ֆ?À%��f��}�� WH�a�s�6���]El��q�g����UP^2 I;]���o�w~xj<mD�Uɍ���Lm7�#��EESOcF�җ�°OC`Q���H�F����#z���#뜝�G����x��J�A��C����k��oS��2��b܃x>�k�s��8�θ��.��4�h�jd�H2�<R-��x}�Ɖ4�g[�����1��G�[G�!(�}/
�ɲj+���|�C�d /�K���Ɋ���Ÿ�Y``Ə�C)I�ۭ	���4����w_�~�\2�m�f�6�6���\�R�Qb�{i���Ϳ�J�7@x��\I��#�޶g'��z��#����x�����n�7Tb�ټ��^Ip�,���R�al<^�9~��Ë�<+�i������|��i0n!������ݪ�A����|?�����Ÿo��v���̮rAD�Ud�N�g��Z�3�� ����&�p�.k;�D�N�J�-{|��\4xLxc��6M��ۣ�o�1m�U'�Gs���/'�����)g�0�x��yIM-:��l("pe���w�v���SIZǐq��m羥6�5���Q6os�;�w���w��
���vf�UC���@9{(���D�P��v�R������Bڻˎ4{>���z���7��#���>�¶b��c�By3���~e�\��A!Ĥ����1R�昅`�ގ?�3��
�Rm\]y�o,�H~��$�r��w��Cp>$�pz{����彩�"]��Xg�_�6b�<%O��Bm�.���.��_��(�Y��y��s~,�6秒�D�ƀAhb�v����.��C��-pݞ���f�Ƨ�na�b�X����ȷ:���10V9㵜���д,
��5��;�Td���,n{�n92���Y��hT%.ut[�L��"T`hI8��R̠F׷ͷD�/��m�:ʜ�<�M9nA�j\�1Ĩ�����P�6���8
�,��_�h� ��H\�$�g #B�d.!{82Q?��hu�&/0|��)��!(�og9�A]J��P���^�N�WTB�4��	����?rI�%>��͔�z�c��xX�5ӂ�H�9Q��`�qL�f~��[&w�|0���������0\O�Ң���RRU�J�}�0,����82��uF!�%Sc�4\m1�}i�UN�QTd=���d�����(�5/���By�4�)��E}Ĕ�����
 ���l[3�*��а�ѿv)����_,��xN6��m� 25�����g��E�6��9��F?#���oC��qڑ�	��DpS��wOa�{�anYۊ=�C⼲��b	C�� qF��B��_����1#��t�8
�����P�3���e�CR��P�nY��V�Ԣ�"⮔]|-�,.~c��ìq�bMaS �7`�(Oty���ș#+�Z�5(sc�)�%g��B1��@��I3c�,»ѯ!�v��u�B� �r�<�b�0�[I�wDd�?�*z����Mi<ٴx_JL��k5��ٖ�y��������[��t΄?n),͛@6�I��o��/N�i�J�8G�I�ܘ49�P��-! K�nbrW�1�Tpܗ�R�f�H�HB�K ����`c?M��� �ZAK���Zk&O�K��I�|�Ф%.���rŊ\��\��������	'j�c�ґ���G<�B:�9K��}f�	)z�'�ך��T��'�lr�X��83�Y2'�b��;e�ț$��i�^R�hl-c�>7��L��;�]I�xCN�ݛ</ oB�+l��Uiy��O��W9r��/��fl��9>����_߹�'e�R<���X�_n���wȜ��5��3T�H& O�6�o���rBYZ��x-��GIU��VȈe:�H�#S��ɽ��g��ʺO!A�/T�#=��]N����ݔ�9vI����sfXng%\����JZvT����l���({���l���7�����L�� �WF*-��ځ��<�ƪ?�?�uh+1�o�O��}�A��5�� _� -�E�iY��6L?�E�>��}��	����I���iTm����|d F��P�;|$����*���otM�G����$����,�� l�F��QKi �_S+� a	8a 1cˬX���I�߂�qE�f!�iw�i�<Óm��V����A�#lp�
)�;�<\��W_���9�~��2l࠮�1���.�r�|j*$�c^���+�KG�|�Mv$�MnV�.A@�q��~=O��s)�e�n���5�]�Eh�U!B/&j�����ȉvUM#�t��7�k��_�|.$���{T�<U����f�n��YЗ��<]�N3A��\����4*g�*$�5?�Ƌ+6P��-y���駣��fGXN:�9�P�,!��dq��'tG��>��{$_6��v�ҁ�=j�Ɲ��E�j��D�:��܌�1	�+[�!*ZB;���ԛj6�[�V�����"G�����,��� �vzo���
.Z����{V�&��었g��V�������n��ݝpە!����ٗ��<:F��l�RM\��R<;�ݨ�ď5�xj#�J���)"d��J'c7���}`8���p>�KԲ0̲MO�ׅ��.�l����H��;ܼ_�j�PY�!&zYO��X��ʻ��X�2�mro&��tҼ�����ݶ�VF��T�I����3������l���	l�ˋ�c�Uq��cjmey} �T��im�K}lDmlϊ[�"4	L�o���Q��囚�H8~��nY��d����3���T�#�'g�������~i��D`ړ�U2��&����)��)_Ԃ&��7?y,ᶈ�.(��զ�B��j>�'��s����YN��X\q�:�!�5rT#>�����[�������dQx$�L�8t�n��g��29j�3,��3�̅܎]F���;�Zω����՛��츐�U��L��̻TZ�r�������
��;ލ����)�b^�����֒Ҋu&}�
���ؑ	������?�S�<p��h�e*������1.�2R��=��T�4���(�]�����qQ�A?�w%X�xg�����w��/�CF�Hƒ����j�**��pG�[T�����u6��ȗKjnS���,�C?�� �P0J�|��dFϤ��t���LvC��!c|�V�@�2�_��>���C�v�O�p�'�=�W��kY����ܦ��1�^.�2JO������J��6�Lf�[�mn��9��"�S�,.Ր�G�����D���{���5� s
̕v�x����GDkSr+<�lk����	΀P2u��~��ډ��N������1����"���?�[���L�# �;	�_�U���5c�d�:[�ݏNߘH�ɨ���;�����U���&�������{���������!�Ud5�QT=�K�����v>���Z�3���^'�����|.�a��А���Z�\]�s�u�ݳ�[@��3�S�M!��t�Y����R����������0��z,�t�d~�b��r�%��y�[�SI%E�{i�>:�EČ$���]CQ@f����>#O`2Ruz�E�Z�g�k��h-Q�jP�*�l�?>+,�d���F�9Aw����ƖB�7:�K���ӻ�K�*sNl�������ˠ��^Q�j���Z�kOw�����6�5�rۋ�o���Pm-�V��0����H����{Z��n6�T�5BL;t�SL?ܓ�:%�#��z*���t��]������X+R5캅}��ͯ8q���� ;� e1w�a�uV'�UL
k�[���I�T1�ՠ1����6x��?�� �;�䵼6c��vD�+ �-R��P��i5�zE�)�6n	�{�.j��E
�e��)�P��~M�[^���)I���l�@����O�/�lR�m(��O>B�=s�t�QEMޭ���(���� ��b[gk�@O��
���l���O4q�
cg}z�.81����`op�`�s��ޡ�8@|��qM%��{4�&���
� ��-�A����KV��<l	�*�*{�#b�^>��a������ &��n{�:�D4�_���:=J���}���o^:�1ye�
��K�n��I�!ݟ�1��g	ߔ�4�L�LY�e����ڗ�6>�a;��p��e1T��,���\|%i����WT@�<H,4K�h�ob@0���l=�1g�T���d�^�J�aٚ���-��?1y�Ыy�B�;ToOeU��yt�7�I�<�L�̄����g�ε�X�w���f&,���N�����X4N4��$��z~c��U]�z�iO������Q���;{0�˅+\�v�%u2]q�A�Tj�V* ������Pm�8#}���&��YJ�9[��~EU�E���t�kmi��6}j濈q�|��'�L`����*Y`�΅��t(⊛ۻp(���re���\7u�����R���)^��3�C
띶I�	��B����-���^�tCT[�s"y��ãً�^���y�{h3w""�P�����a@��p�P�e��sd8�M1US��g_;�(H&ɖ�������f�ZM�gn�/�(���A�i%R��Cx]��;�CH֊���l���h(��u�Чs�7ؠ|�]Qn~f���|X(�sb�ϵ�_u<��AiJ�|xy*_m
vfNr:e�=�� �&~{٦�I����߽����pAO9��h癮�����G��Ĩ��t�#�lj�GM{�BTJ2�82��R(w�M�f(���Z��������S
;r�(�-�gz�-�r]
���˪������>�;���e����)JՅ8ƒ��aϚ5���E�r�o���d.Fh������/���8gz��;�)a���f2���㒋�8f��p5� �zX�)�3������}A2��uA�j1�8�v������#&i����|(�(� 9��Ú�.ei2�9�<����3r����J�L�H���1�,	�������wܝ�g���TȠr9��a>�S=	�S
�l!8���0�t�
���hμA��i�P[�|[͵nJK9�:����oଓ-o5,2ɜ�ck�3a�θ���ilHE\�|��ŦlP6X�JT�^�Srl��y�^�p�m�B{
�>γA�I�|�q^�oN�����}g����W��c�1A	�������9f����M��:|`DlȒ���d8����I{تH"Jr%ڐz��$b .>e���/E+p�/�M��#~6����l� �7�r��|�f�h��'S�w�!M��!�>m�J��;�E�p�x�>�!@?z�p����:�H���g#̔�Ӳ����N�X?�����XZ��M����K(T�$}'H���A��U;4o_���\�c�`�2�wZ�����^bQZR�\{7�$cP��#L ;1̂� �W�M����Lk
t�9���Z�>�H[��sU����[g!7cs�Q �s����6x>�,;�۱:sܾ�ӛ�Eu�ii�D/VL��wGp_��>i�7tv)Udj�M�fn���V��?�n�
�3�Fٯ�02���-������ӿ����-3}`��Z��W�a {�*��E��k�+��k�W�i� d��?ʯ{h��� &
:�ў�{����(uP�X\��#:���E�2ń._݅�zlb$��˖�0ie�v;Ds�[T�� b,�o�)U����ct���.����(;�
�&�@��OU��0W>�zSi]C���Z�:��d��QЅS38 �s�
�~��n�����j�E���I=���Q�?�D{/z���t#Lzr]6%���50�%E���W`�@"�<ո��
�*�)ul��er<N�fn����"pw���(��8����G�kL�;E�����2�����:�J*:�%��;�G��}��]=����P3����<JþF��Mv���c}�[�3S�Cg����d����9Ips^,��-�E~f��AS�=�2���Պ]1D�Z	~y���n�BW`ϠqM[m�g�;$��f�����JFZ��R��[��q�ث1�����H����.%:n͌�d��w]`_π���*�����O���ס���W&�����gN�bݕj]��g R��\X]�+���r��T�@�EnG�0_�.�C�pM�=q�~ω�IVDs�T�����>AGħ�M@��3<>����B�3y��d���c�ڮ�}��&���|�J|�&�}V��}v$����J�=�q���h�8���:zD8����7���)vgA��o��q���O���?���k^bFosjdA�X.�m��.6�t"1�%�n�ʏ�k�0�W�/	2B��B�p4���&�dj��yuA��y�f����Rv�,�mo;t���3�.�_���"Vi�T?����n�<z]<$���e܅�����ⴓ�F��B�&6�t�L��5$�ߪzs���e�a�.�c���������"� ���Y�V7$s�}'�H�v���9\�R ^Q��5h
N�v_�,9y��q�R��Ρ19V�Ox>(�hո 4�=d�x���	vvQ��~}fg��:55D���*�Uo��h�
M�9�<�A���73]�ꇓ�^��G�Ȱ��1p�Kg�*b_���;:�R�H�M�6&^����U�9\�Kbݢ��8��M�#����ր=LH�*t��w��g�� �p`U�"J�G*�����p]��Eɑ��j�]+��>���&	�^1 ��Ƌ��☴.3GG�r0u�8`�%U��ˠ:q��P$0�yv�̃��y�La4�K�a�ޥ��\�&�� '�����[N,m�����)�͍l\C}?~��u�T����9r�ET�EF���Y�Fc�Lp:geφ;�R��y�AǍ��(gV�2���rU�W����oӌ5�o�*���& �*強fy/��QMK�H|�J�/1�YdO�K(ȏ���Q ���VCmM��k���WA/�b7�8J�}
���p>�`�����T�����:���w���V?)|�[l߇��4~�`��6���K\E|�5����}��vP����d����$�G��e梶]o�U�a�u�
�l�(ϴ�v���Rj>EZ��Y�W���ω���	�������8c�1�g������N����ǌ�3�
������=�z[���SQ��*vJf=qq[��v�O8Cץ��R�wt!Ԇ�,�k�\�����~7,��m<W@gQ�\�����N��J�Y���qΕ����U�r#����k��.҄���x���#���V�xG��3}vg��
����I�L���_�!'�7/��F�W̖~�*��n�S��d�1��9/N����,Kh��e��2_�7�PJh��ō��!p����Ku�A���[��ST�n���Q>�`���|RTR����}�*��Q�l;�"e<n	�7�B���D����ʗ��m7<5��S(����53|ۊ�,A{d� '�.�򼙹:p�h%O���\��q�&v)�>V����q��j� ;~�n��B�>,�TR�=J{wM�n*�*�Gc��=l�0C�sOl�Ay�q
��K���!7��۽6Qpa��������`@Ub�����b&D�æ&����`&�ԣ(�ק1�SI�|��aYWRK�h��S�U�ơDZ�(s%T>ɶ��ז��N&�9PXL����:L{6���V�9Uy��Ifv�ןà %�M��v��D҇=u�!T���A�I�3_����b���/��[��̌��Hw~=��أ��8|z �
�3ء��	�o���Z*f�43���i�v&���(���7\�7��9��<�MzƬHM��e9	�<�
�	�����䱪�\�?GD�3K�6�A3u T%�͔�ɂ�^Z!�ʭ�I�}�dP�����E�J��r|9~�Ѝ�4ӣ/v�<����;[�5��w��7�^�)˟���D�� �4�LECdZ��
�Km����w��A���]X�H��!����C7���d_�G���!�!$�]�(m��(CD3��Fr&��x��J?T��)g����=�����ۉ��d�uYe,���|�Į�8�2��wk��t�2�j��<���:����[�w� �l�{��b��W��HʉR9D&Q�qK 嚾�&)W�*[{;�7X��ٷ���b}�Sn����"m&7��O���,��h�L? ����"mBZ��[��"������;>�Dk��LB��mե�S:������{�jGmw�t>H�k�T�.����A�J�=����L�����P���n�����}���K��b�AxFq�x1+zw�4]��֐�K�Չ�f���B1L�7
�%�LuH�����VX��9jKV�2nڼf�13܊�ߖp���]n��%��r�,��Taf��	uN�ڴUM1xdJ��[e| 0"t-���&#�Bu'&Ghc	���S�E��7�v�$NX���<��i�,�u��V��ݯ��W]��JY���(P{��g�i��iZ����|��v3�BJjN�v� ���W7tm��U����G���=�M����a,(K�Á��OE�o�z���[U�2��Ae^����?�yo92Z���c�VR���3���<���B7kh��5+|��6y0�|hK�����!C�Ji�1������8c(�y|��&$���� d�����A�@��;������?72a�j�pi@�/�1��t��3`r(]�~t��X���T�Aw�^��(
v[p�Pm� ����CeU�)C�W��+j��Q�W��-�p���\�yz:ą+H�o���f9�=FԔ���I$:#���N$+
V���#ӗ�����2C^��$�J���.Z��d�Ӑ�cR��`rK����'�����2�p���xߝ��`�ʈ�����̠U�+�QjES����E��R����ſ��m��������f�LÒ�����fʍNG�����SM�-���&�x�h�P[^��3���gW��b�=?<�*с�X�ط�&��g����Q��r�4y��P0�;K@^�5�:��%�<��ɱ�r[C�TP�(�3�۵��ub׋��Q�ԅP9#���ǅ���Y]C���(�x3���M��ç���b>��@8����C&#TPxo�o@|2�S�����GO��A�Y�X���̕Ӳ\�m������w~��9�3��*�I�@�+(�z��o':)�="��V7�s?G�[����NX�*c��?͵ѝ�.��x��"�i|������u� ��Bm�na4]f�d��2ί�-YFDjb[k�g$R{��e��v�$E�=�#���_����o�*����FB�'��	��b:�`������Ϭ�x^��}���(	w��?v ϟ��=V����#�>$j�سcN+���oO����u��РS
Z��ʒ�6��F��t���,�9|B2�"Z����D���ll!�	7yWQ���Yv����f [���@/s([�]��{5��EC�x{�kd�#����}���,������t�0Ƈ�O�Xχ�bb�lW�� ��:�Ɯ�M_	�_?c8�����%��L�i]���P���A�¨�ä���Y�<#d΂�3�������U�9k�����4ک{ '��+��R_�K��t��h�/� �C0��3>'c0��ZZR����\�/jާv�fzPW���	M�M��]�%���g!Z��@�q���']�m
��i�aQ�o���>9�6���S��g?UPQ��b���uj'�z������_I��$i��{5-.v���ǡj�8�7n��@h��H�h�Ѥ�*3����Dd�K�p����)�4�3�;���� �fʩ�D���ݭ�F%Nt�x����p�>Ѭk$��J��r��o�ID�J{Bs�L�&w��rO��~x��d��xD�i[��+<"9�8���S��F�>�=bpX���ʬ�5�#=��M:_. ��#A���h*Ps�wVa3�����Y�e�L�,{r�t��!���;��3ڿ؊������-��57��N	��� 2��������FE�CJ� ��od�,M8t����/�Xyx��H�-�-F����;���Ya�@��p�Bv�E��Sh�:x(M��(G�tɋ�tH���e[�i9'W�O�Q<�{���s4Oz�.י�m�8沖`�H�=����"M&"fw���F�<��:X)�j4��Dv��fƇE�3��:ϯ����D ;>�*�/�E��]�wf���H#l���z�N�'���m���¡��>�m�؏!�|��Y]��+7}�Q(��Sw�0q�g?i|���nG��/DD��A� u�u$��8 �V�Ó�6����V|;dgEd`I�@�`��p�m���\���WeЙ�����3l8-�d Ŵ�v���BZ% �;��n�#��Lo�!��Q�"Vޝ�<7l��"�5XB��p�,6�ҫ+�-R��������?�+�C���Fe{��.iX�G�]�&K����Z��=�
�E]	<�Ԑ�	������qֽ?)�qAx�Ì��|��A�|ß�r��)Q�-����O���p��2 ɂ����V
�/^�JG�B�k�.���}�TɂU�=%�g#�~/`L-3�g��:z���(�u(�dfG4tpz�d}H���e`j�����⥻]���l��[�6���jf��9s?]Sg���?�(�zG��:����K��EG� K�F�ϛu���%"���tEG���J����{th%����@��Iu��u	���=��P�-�����c�kq;/z�`q,��39I$cH��P��6��M�y�/s�,zAg��nv�������
�p���61�|�F��B��**\;T��w�!]�M��L�w+��m�����LiO9�9�p,���*�ܸ�ߕ���VnxER�j�J�l�������,�?"�n"í.���Xr����#5��CM��\!-R�!��r�uʌs㤔�![�o�ª���C���
yg/���n�޺ICF$��6N�f�W)4׋��F�f�W�yۂֺyu�Mh�W����;*��&f���42��4:�F�F���K�\�Z�e��2�;��%y�8ߺ1Jz�yEl��Se�,Q3q�,8=�^o��O]bP!(mT,V�˩�3)�'�L��~�&�4m�~H�*fǞ~�ܮޚU\������K�p��ָ�|Al���%E0������l�M��aق����M z�O��O[�&-�%ʉ���:|.ARo�VoUrh͜�e�D4�`I�̳�!6UN�/�P����/��ɩ���VN$M�[b�mE2r�{1���X�[�����Q��L���=�x��x�C?���k�S��±7Us�r��0�G0x�݄m�Ի,Qb�� 53{�09`+l06��4{�z�M�m�CxhX�����-
 ;g��$l��K�ǘ8�~-&��6xqӦ��UG3w�����(ju]ó���m�_ ��c�=ln8aa'�sX!;ɤ��{���
�n��V�����7/��H3�����R�2�U��X�]�(=�{�K�x1�k,k|d�J��@R�џ޺�:�	�D[O�7t�T�V�#�����h��SE��1��4m?��9�"ڗ�⏈$w� ��g�.��裤(�̩�Pmr�&~U��"�H�\�A��Üw�Հ�'�~����������d�_��!�q��3�ل\'��0����8��^�K���t�� �����P}c��#�{�?�@.�P.��AK΁��ܽ��w5�p]���"mJ�0�S����Z�S(oq��Tf�1�T1U�.���0�j�e����,��B(P6��L8�1�y ��!B�*V�pT����ha��Mv�'Qc�$�OB��	���'�B|�O���ڠ�v?ȉG1�����}$�3d������=�K�2��PX��������-��j��@��1$����谵�(����]�=-��O?ۣR�D��mg]��)#i⍊X��>��?ז�y��W�🆶c$wa�#腛�S��Af�cU�duQ.x��m�CLK�n�y��X�s���'���(�ŭ+�XU>l�p��pDwGm�G����Pw��{M�jh�Wup�xN&6^*$XPe�5�@ ��ep9�U���vaODQ�+���wr��e6�	/ո�����gD�-;v�;V���m���wڿ�yv�!�]�v:������| ��T5g�{�ad��7�+Z��#��/ �3ջN�������@��a��l�j���^2XE�m�K	�;B�7��Ck�ZE�����#VؐI�泪�����ܤH����w7�w���� ��kc*KV�U��'%�*�왏<��2L����آ�B���J��O���h��!i20򪉦ߤwg��Vw��h2��$�̾0�?j����7;����6?:��j���M��P�\	�����M�\�XTwӿ���u���1ڐU:������f蘾�~��#��^f�F�����]\o'/�j�7�J�����û�A�q�Ւ��.�ڼݾ"�@#�H�?[��Ѣɤl��K��ъb���_G����W�]+�ǫL��}�@��BBn��j�)�t�!-:��/d�t��=�J��ax��߃PO[��ha�
���`@UaZ�8��r���IV��>��P�p�0�z���ɍ�u=��tOج²��.�@/������|'ߑ�0�^������j�qzq`M^�@�
l����/�R/s�+߼��W9ݪ$�
ü1�lC�����p�!3U\�%��[�{
������+y�������c�jTR�j��$5��_� �s��:Tֿ$ N�y�6���=u Ur�}+f:u��6'o��S\���V65�[��B�Ion�*B	I,XM�r��qp�F@�����O��x>�	����쾥���%��U{�
|g6c����2ըV�,���F���r'5�,�`�� �����>kf���������4h��M򞸡r��)7!XS�_�i�>Dսx������<�l�ة��8/O��;���_UB�Q]~�1���}��1�UF��1&rNSC=���	��\�(�}�
/T�i�t�b)N�LCF�J� <�`��!�B��ۡ9ˋv���K�b�b�4p�aD[������1�}�y���d!���U���N��g�^������"��pѹ]ߠ�Z�(t��M�e�P��UE�u�Tq�����V?2*��,�$����@x]�c�0.��=����w2b[��3��%?s4� پ�Ń[��V�d�S�V%$���9_F�ig��(��
� L��|��x�P��*��JY�m�K��`�>F�h>��-a:sy�hds.����Ț	�n�xP�%�~�)��3�����sb�?½M*tF��i����j_e�M/�K�MɱY��H��7�.TO=ܩR������{VeL��u<"#��"|c��	�̷��X�k��ů�����d���B#���3<əCu�<���:�[>����Е�����~�c���p�0��ƥTS5<��C����`bc�ҩ��sܞ#'���ɩ}T�P��k���A���> �l	p�[�&9����=�
m��]�T�ۍ���0=�Ȳ� �)ʙL�ˇ�7b�Z���� ^$ճ��ڔ�6VDXZp�����횪�C�b��T47#�N c��.���~0��`�3(�q)5�}2�pT�Zla�#q�X��7h�T�n�Ǜ��Q�0�����z7�,�;+z�l
�މ�d��LL��|,l5Z�M�D�h�QiL�?��԰��L=�����6��v�b�1i�Hw�K`�H;iy�` wE��Y�pn5�ތ�m�o�\����jr�,�tV�Ǣ��
s�̈́�6�`�x4���@�`�(yW�Z>� <[�b��7W��m�u�v�I���-ta?�J�q�Q<�:Uř�,�IǊ�k�T;�M<ݚ#7��0���~� ��Й�X
��9�
�t����6Ī�Wl�3���ڏ��ŉu6�k#�PПZx��O����0�h����S}�з���t%L��6�c���~��#k\�MG�ˌt�#`چ��X9%s=:?��Җ��z[3(�}�{��y��,���궊G1�{(ؖ#��vg�8��6!�T(ar�?�nN��t��Jם^s۝נ�v��'��$�7E�<
S}G�A���	s� _t��G{�pG���x�%��,ad�I����v�ɋ[7�H�i1��蕆�9�dXyw0͟'8�r��5[n-6{��n{�NL�D�9��xZs�@�*�E�T��D�2�T\�s��5Ճ#�h��#��D�0���.˨���@~�BT}5�9�8p���$�8m��&T���SF e�-��ddR�x (�9�����>�b��T����D�/jؑ�a<J�O*��7.���5�)׳r�ϴ���}O�\ݪ�дl�$�J��QX��D�a�3��$�](��mV��+��]�6A���8�?���e��1A#ޓ�8x!��� e���Ӏ����Q���-i�_ִ���ո/�N#?��zI�N��\���/�,�e����]5ᅫ���N���������0�Q���)M}�Ѱ%��O�fI}�3u���_��'�.�7��΍���������s%G�D�>���O��8Qs�e{齳�� �<��?i�~��yTE0��#�p��V�(�Q�����_�3�P:9ؗ�Ff��;l�zM�K6�����bM�2�np�1�n�}��0H��ԗ+e,kS~���Q;��y!�ŋ�m2�z�8���4���ݓ�&���$��z�z!��PJ�}�ge���@�%�G1���ͭ�y�Pm�`�c���s������aw�EL���i���6�8�h(���N^�,��q�;�
��1r2�ͮe�7���!����͆ժ?[B���SCi�C���gviIθ��M����M���ג�����K��{�v���O�,����ZO!S>84�����o��m{Ȓ����U]��ai��%��;4la����o�Z�a��Rd&i���p���W�]z�j���V��o��D�8��d��j�ux�l���9������-��瑹�&{��'dP{�.ˋ�'g�
���=�e�_	KD��{�|��/�}�O'�gx�gA۱E����d��΢-��^	��.��X�ʿ
�P���^�7?��l����􍯍�}.~���Vo.��"
�A�]-����[ɼb��cn@aA�4�o*��!�R�t�\�C-w��8
��4��$̄�]�ǉ#��]�S+r��,�h�r]�����"-6	�#b�{��R��;�2�E�n�!��ށX��jH8ѐ���qDp���ͺ��t/И�f�x�9�ᯡ/�@��G�B��._��$".���!��P�pߛ�5�s&�@�pKr5^$�z1��ݯ��C1��.L>�_�)U�뽼�6K����jI�%����E�{%��=���u�
~�� �����L�݉Wa$����Y�F�͹��Q�+�y�e�^���E��6����?c0�������Q��P�6xI�v�D����mY�!d���@�� ��n����y��Q��	Ȩ��$��H�({8C��K]�ʢ"�x�3�RYc��p2����Kw
𞅖�)L�慅�T
V8\jp2�o%�򌒐لM�[���U/�84sۿ��HH!8��\F�* 6~���1�k�ĂA�!�Ϫ�v�dgu�5�zAa�J���4��^��i�_ �~��a�"n]:X�ߒ�Ծ�4�I�9ݢ�>���{�c����
T���T��aĻ�64}�烎�"\�2-x�M�!��#\)Jα�&<vb#rb.%��XP��ѱ�L�T'��EQE�5A^ڙX��Q�$YǸ���`<�g����F��(���-H����;�? u����*C�8I_�ȼ뉕���+sH�D�JYu�Dͯɬ Ǵ[��|�J�p�1T ��[MaX�u/����~�_�
���>~I���5s�
%�jHs5�z(�gQ~��k�q����w�˞lt��<B�y�Q��eJ��t@+�n1Q)B<�����ܱC4г,��\p�5��x�n#O��O��'�9�4���ԇD��S�WAK�J:���/��t��6N��R��OE+δh�W�ph�;wq�ƷCʩQ����{�*nku�[ZUO4������f�����c(��H�y�*