// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kkEI/A7DczI8rM0ZXgNlMZrlfcyNMwE8r7jgzpwLxCKaqsdMrhrLSZx7pOFKWW94
D0aEuZTj4WfTfuMsYHIgBJgczj+nGWobN2RDMjEKNssp6tSGCwWlWvIdfwB4cDZx
2YplUHRFKwt1UonIgGVbvGriBMuhxKz007VU4V+hddY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11248)
1oWtXoarodE9hsJMyk4IBzgMzhtAQRDAPt+62DmoGBYxvhKHAe4ZsDoo7joJdyJZ
Z6DMrkDIcLKPE//CTcHq8urlSAH0i2QOt/E8gJNU8cRvKt0NnlsSlVM31ei0W3Gs
f2F7O2AwBP9+56wh0IEmBb/rfprsVU0JzZn7ZDJhYF0JToBon8XtthK+t5D43bMo
bQiDtoN5Rq5HePKnEMiBFvji7rFBaoM3ijAgjTPWjRcY6F6F1dUujwjyk83uuZwf
+XiakILGnSsi20OePlr4DCNT3JE4IjkyjSYQlEeNRVhhZfGgaXsPBOk6jufQYDbI
F09nZWIcijrcMxDTf80QAMHbMRg3QJ4LWpetf8/4GsaqWPQnT2lZxewUa+2QldP4
Dp6G5jNZS1fzQo1lZQRCJVw3IhejKUyeVPKFdPxGyjOeYoyF7KvnEkrT6pKhu+ZK
2WdnrvsjkHCJr1jAinlQ/thRHIIVNExezZTRKjnetMlj7hKi4+zVeCfXsvleOdqH
qrNUuDuaoxV08lQM/X8TQaTDjLZO8Xqn4btEnEBa63M2oxjl0Gow00eN42KBmCCX
DWUmRBGmb3lAK5+KqPF1gbX7zEGZv7N0Re47oJcpMQTOqLRhJamBdeNm91eTPfmq
Dng+lRB1YruO4JVYxQdxANKbhMOyDihlSeI4zlZF8H9oyqm12xrOm9Sl9IDn/Tl+
EUdzzT+aHugzlWCM0lFC+jPfVQXhMYcAqZq6BcMS0nBCZH52xZsXlmWob0hdg/5w
oYovwo5vmjw/2eV8aaKRl2QweYaQNVGmCInh5NJQLMj0f9oLTFELX3uFqrAQcbjj
rRFQBDb6wO3+u3G9wVQ3+FhV2M0hLS/HAP4Z1liFwHsixJxcrxeUUqJ9VwSHnx0p
eypKJjJH6kJ2gXi+8R7+Xwf7QVD6F5Ytf5S9VOJjQAmmVh63/4oAj8twAhHU9qHa
WBEqi+mUoKd1qH7FNmWcghJ8hM5D5UlzVuUVj827VUQ/MyyI6xub7TLGhGZ9qk+2
hvHoKztFIe1IMkbjoLkLFNgyTMZry5CKr20YnkuBu6iI1gc4zhjVv0sXzSKX8YlA
gYtS6jik14gxHpeTkv6OFT7449WAOojGzRl27ZEwOU1MGT1zC6Xx1pNFisXo/zTa
E5S3SijCICuEnQpmGKoHfA3yTsSiN3Zbpe6/jp0d6Tt6uZ0L2gfBNUyCzRIHEnNP
k46YUCeJTneARwYUTndD5XlFbFJOaV3FVfa4rPuj/SbhjnI1i5ebMP+luX3RdCrO
WGKqRHchukGllB3i2BFe1AjAIJX1mRbsroMm75HlxAgvkXyszqlgDIiFPb9jJdFk
Kls4a+NiNumLnzTakOwgczXpnN+g75r3fMwsuUQ3LtmFHau3+IsKXIfUpkZbs1TM
RibFdIKukQ7a8McuzMDnWQVW0PCvsR5L8j5U/1NShIzmaJ/UkCm5r6y7IjOvAUvi
lldKRJB+usQhoNPLPJKNzYVZMCJD3z78uR8WkMeiLwML8o1vWJgI29jOCIpB4ILW
kngUa1Zvgm0oWuvSWtaQ8Jy5aLt+XhCUPkfd5/MRxzcUGkXUD9hxtl6S7ZHAE9XI
kJPTkqluCXuxyHH+zm9FaqFTR0xe3fAnW5NY1AriKA1RVlW+jKZ9LR5jgXm88rIR
ZrIy89R1f8kCe6Kqdz15eLr6+uH1YGN3O+3Gp6mM3ywywWSvOFpWm3Ao8fIf4Z8W
VqFog28zCwOByrWSkFT/+NG3U8JvzZJ9ZU6fK8jemOS3fUTAup/FLVlTTA0hSfOt
9mD2RdMDIxPwl8oSnmgJUIKcb5ubP+mdi/AJdzk7KE+Im1mQYLKzM+H0V6YLmF9s
1EUHpxyUVByd7xd/nClUoknBg8z/cfI8fL1eM12auL2p5ODbXiKGtfQyy2XD+Pyg
5/ulcfrMErqCH6shGVQQZheimgIXlnwHDQDHMs5th/EQQu3LBMO3sjNQi7kkA6d/
6ZUksRsiEptzfzlQY03SvURVsgP0Tpn/r7VjTkaL5OJ/mjyg2dC7yMGXCrjjpbhD
IgU6w74o7YjFJPHxKcmDL926pVuE/3G9NV457QiEOu9DVAOol1SdvRxovJOtFVND
3AUA4v+vM9UGOgtX747K/HPuAXktWJ6beIwHZe6kKe4TcS2x2bk4ex9gGqq3NrEu
jDWMbtW45bTCJhLnAX38brwK0237EM+x3g/Rp2Ic88ztugD+ZX2cpxSQNk3zjCbT
UBewwS9rniXu8bUsbQzEFjAdApdwivzor3Fhw7qCBlv4lan5u/XiEHwa9/Ok8Ftf
mQevDeVEHVO0/xEn7du+BAl4CNMTDQCZxYY4zZwufLN2pfg1HTL8yq3344/fpee3
5+FLRBPJ8sEzSvq9Cu540Tsd8B/O3uUX+NHrsZnttzbfTiCSsrBzkfjy0OanUOMa
LU3MXbknhWFrQZeiLCFmh/U422rI4b7tT5edVokcDoC28QKDDgXmq8R3FAmwWHhj
pHFYkGiRLU7IGp7f2eLcun9mjWgik+RamD8lIoXwPpUkKBfBUsKAziBDmBzpcQWe
6FzxlvSNJ5+7ms6H3dI5a27HEV6b5lDib3ssSK246WfgDbwBdfNbg77vIAdW3cVK
Uzdv79t9GeJJhQ07Mx0KJFhhE0bW3q6rpT5m4RMxk/UDREzhLiLVvCrqstY9aeGx
foTVmdQ/GJ4xUCt0pJJZSNKiekzFMXdr6O0M5K3RmPH7pbQNMYGRwuQ93L+5B/9S
shoidVka70fNxZb2flF1wSuQdldYB7oDhEl6YsowuPhgKmcTP3N8Vg4HXc68Hpdg
YVrsOiTxqv+3pZYjJTznmS7h+0hJYQhVW2yEJtPwkSqJXB4FVrRUBoJtuUganzA/
c/GH0Yvaz8Yph2FeMgN/TVqe2hBee5sOHCrTq8tblnvcLxEnrkRIyVcF9x757Ugo
8FzP0pVuyOKWuUWV4oLRtOXXLz3ALnNMtNPxLPhbMST85STeVGthENRhOSE4ASFl
H5PjOvi5tPIUJvQx7bPOHdRBwW6nvhrsHAeTTUmjulOUoDxjwLYoVgSjJj255DDi
asTepoQxgj+eIExcGAiPhueCl+WgHQzUdIQMLDFntZHjIsDPt0N1mG7EJyPlFezx
JhbsYUCnY1i8P2caPmdPAvFryGs0nSAPl39S4W0Q0tIuigCujDbZfEv8j6dmuw03
VrLKTcZGf4E8MtqQwrEaeOIHV9yAx9ajitANIHFWiXfbJo+BEDakB71sRo8FFv/1
EvlnnzsojZXJNwWToZgDEeKPbfyeW8LaZTJ7sB5YYW5fQhwGDiEz3pSah9dopDa2
ndr+6BMXhDX92lsX0doCiZD82sc+NoFLwW8FmJHsOW4sehCceBlWy6C+5Sp3E57a
Na+Vx0c7Pt1M6V9IkfkjK02z71s2iBCxnqqHlVGaDLK0OWZC7DFqjcHsmJE8tTXp
xvmYYkenC0lwyaf9We2zOS0xWWZTUh2Ik4sVdTkAUSPrFbgnbmVmjSf5TrKZvNYT
3T2v3xAA6W2K/MDlGLBU8zGBlpsmqeSueHwtiuLmgws2H4ayG4a3HYY/t9tPnmJa
H9MgemAFMP2+nxSCca4gC9+EVyxBwyMTaTI39D6Zov4vtqGmfUkrOFJYj06+d9Mv
PffPmQ/2S/0XBOyu+P0Souoz6ctK7vMsVl6sQxL2KRPkhSuTK8YpNXoBvbV+bwsZ
Lz5h1wSFt78OIom8BokAXU0Wh5pdoIdD+YXjJNDO0rTiNblxyJB4o3dE5Yhf9zuO
GWSIbuH31xnFEyJnzbneDZJM9Vmdp0n994ont3YckmsUDozoFcWXfp+RYDE3yO4x
rRWJDurW/+MYrvjytQYOCEhBp9A/mWscvAsyYGOGsOiQwZuy9nLoSStOImRWhLgn
KjDPCDRAhr96eM70MbdJ2r0wlL/YYBRJr7vZ1FYldQImm2vu8U94U/ASHIT8s31m
fV0om6DyJCYM6SHjsrZChYMS5DOkBsG8ZmApXNnSxwtWuQmfs1sIJy/z6ydFwsgh
wrQPdD1Q7T/XMLlBSfvaO+/53BJCL/e7w3Bj3M4oBX0z6kxF2aK57MY1bvTzKg2u
8sQrx7p6kmPEX6s5U3w4vswQh6mIrYwF2fl4oi71bQ00gdD6zO/YRthhnRhxOixy
VKKYAQsA1JbLeXwwMlyLdBWs3paRjMaR+m4hRn8/tVqv35VtVeObJCTHEWn8fWN0
mt9ySwJDrQ80s2qcMvIa+U51rE6wKrr9BH3LkdeCFNnnp6oyB3zQPUagBr1vCGHD
qiKrpBJqyPvmu0/DXDVFl2AGq/aPxD7T+9IGPJkvsuYq+TEvx1LtZ3LX9N6HH8Ku
KV7Za8THFxori/rVB1WzrVugk7ZKbvUto728q5xDHaE6/rpLKAfmBJYT62M2UVAk
Fo3Fm0wWoGTD5VXkcFRrnBYifaWOV0jE+c0Dgi7j179HwClIwBpoHKa/KebwVqAN
Nj9s6IvfiAp8q+1XZqY9I7iInY3T2CuHTJP3BE8LfAnrIdACBQ7NU6Vhgunjh/YS
ZulUfFZI/u+Mbh+lYgkPRh125NWwwb8zM3X9euT+tgiSqwfG3R6XrrvEe0eENNM/
CHPS12RFymPmixW5YLPNWLQpuVvy3WlZXK+0Uv2CpkidWPetHK4uZfnlWdnMDVyU
rvqQhYAMD3GBWVsBDF+L28IP4Mdo2bSLU6Rime7+52kKLjmroqfgriuVcjcDUuEr
r1dqD8uVFued2WKGp3iW79hOdHXw8RYDPCb/sGh1YKSln8KIVxZY3zg0wCg0qPcy
o7JUokMrO0M+cDWOYkxQAr5Fe38TApTcgxgttRqM/TrqpSaj3VwcqPNHvugl/eSe
X5lrIFKuPjoicsiVxspxRlW4cmnS3y4uwMAYdUpuqBz8wsFx+ttT1Yxsq+On52lc
xOolcgFxaT9zLx3b1acZYW2TFo09BzrTmQoqdX/954wDl58tKUYviXBtlFkymTrc
8KeTOpoloGHVU7XUVln3ICPhFBJ4lGDv6DRYCMpFZbb73RB+0WYid4FQdUVF7xqh
gv2v+q166ropetu61yXb3aO6k6zlKw6U2SZ8kvQCnlSMX8xFtY4t1xxLFCBSE2Uk
bjnHmdgE5CcLEUh5kPHyclYXOX6AgNs2O6TTqcencxCe/Bgf+Focs69IGmd576Nb
N4WaNWSvnEXM77ofIA5fdPTayfAq+JyWjomk2DrzOrooioJP1almbEyaVcfk1oVJ
uHSb6Deuc9f1ExuvP2S8wI+6HxgFwhsHjASF1M1ZVMopOZEIJsV6lHPEK+uvCOHt
Uw1DNm2tqBhfP4Qm6CQNCTqDrUtVEChhMFkwxAjyTuxSfZM5gqxn7rX5/FBJzPOI
NU8VxzkGjA+U2k0LyxD0wIZEfmp3+hFZDgZBje567ngsT4tney8+/DdDxFo8jefE
a0OabCOJRPuRwr8n51NBAV8WNuwfjkSTNGSOrqndmGj56GwEDvXm/QxuklYLzUBu
rYhxysvQnvfM/h3ns0RqoqY7J6hVIFFOeeqytEXaYOa84gWYF/gzyDVItdPzpSs0
8ZQ1SpMBBmLu+f4/hoX+sLW6pHV/rpn7r5l9KDlWGVrfh/B6pdH/26K7m7HL3IHo
RvdrnG/sOikz+xEQphR2TZnaVYY8L8ZCRWMz6IqMFfW5pQgeJKCGa+GEPxvdjqa8
HZV0U5uktQh04A/aOmcBObVP5UmuJbachOdz9SogCjTbGe0LLHRhtqvbqy0MAqvG
KdjN348uwCwBDQu1tDGRQDQu/slNuW5ilztNWbeCZ0a5Qpc7Ev8+OpiIUIQrM/ki
I9VgoYFN9Pq1eUMlrT9CH9WhvCugWKoqnzcA8hfJtr98NAEa+WdFVTYorbusijTn
d3J0ElXf9uzOFvLvEwmlGsLnqLIGQJhGdJtNStqu/B1+hTfpR1BqYL8VnEw6DfV2
lwQ/S4wgnxxMb2MflAHnbR5qwm6Gq141XW+EI6QODDhl6ftrWBRNcVeZgnhh/BwN
Et4MTdZ6yVyPdQUPY2wOj31/nSkXjdJQ9NZLsHbxi+tVLo3U6AxhCUItnYrg7YrM
6Gtpgb86Sr24ShbPq+MEajz92ZOtcLREkBUawQviUxPk4HUmavTQJ+k1EwueBUtG
LhE2NlfTjB/9KnTb5Moafi969QVmQW3OkyIjUzMj47Tjm9uKXTe06UVUqGGhhjng
mceGffPRRc1KlBaZNb2mWIL4V763gvaEYXogrnht8xiY3Vtnkr0nvf0m5CCLvJ9n
r67uyNWW4Bza6Mui5uO/lnLyQMnNeZ3BhWUl5m/AZrq+ePqOSzuAFmWhOH55oRiK
rtWqSGrlTHTuLwJFRfhP53Lto724nXkNVvvL8i0Jq3o4z8TLQ9wKDiZKDGpnTsu6
kPByBJmShgKOfCrylmmMqA0UNTe/cNnUyJw51Wu5qtsOWkX8OCp7oYo37vwKwuwK
1WwiIzA9IK6dCXb442q67FFVWLfiNtBYt25hXjjxl8kAwZo/tqJY8/RvuzvdwhYB
c8YTnBjL/Y2QhGZzNvWRWq9MWA1j1REF8r4ziRTiQZLgSJxdYoSw8BY4z9WvzrJw
8DoVB36neSXB7+77gt+Rbajc3ZR7jED80DR24dRRcUOO1vGd0PGkAoD9E55ZtcKO
Cz0KtH/syDGeuht7QXA7zNkgH5JVJtpFy3SnvlmPUerPmYVKRbwdW3Ji2K/kCbBm
1MbHCWyjHVT+6dVEgm1QuV2hwOTMWvsd5/y6/roFAVrKqIyrtcCA48aVrZxMF/X2
5ZH/+X7w6l8Roj7EBKbRBYBU3Qa/tAwPpScXIW0XiuANJuQLdwP/xVrBvKpp058d
Zx0/Kuc79RjMBdkY/eOSWe8JeSSUEg62YmUQGwaI2MZTgMIFbgpU6zgmUQHzY3fs
GKfEj09SJkPGZDUXoyt5ToWoH7/gemcgpUCV7pGYTuuSq6YEWw2T76zuOtGEx3aY
tMHfD5f9vS2NrZV8sax75reobiOVYEQAlAv65NYESmL2hEc7nDWWHu1Tn4h9qbl6
aiBfP21mXtf60fBQXJPKsFvSC71CZrNu6JSx9ZLgtpDEnjya6o1+Xy5AX4pizi4q
HgNeFCg0Mc06+5ctR0K4k7+7DIKFI7A9lZx+vggX7AAcXAJLXsJvtItaYrVYKxy6
FBntvdYEzIM1mnDR3VimbT5fsrPNstbXPZ600nnOdCCqHwPRdXmRUNOUmb6rkBVv
C8moyTbh8kwkLV8vWRODtTJO082tnMNY7Ad4Jej01G8SxdvvzLEB9aCDn40Yos9X
Ah+jeENnKsJtefRFNAt57Xy4X0X/pwhIb3876sPpoJU7Xwfup2nPBCC/JH30kZkU
9oUvbqljx4fVDSTol8N/oNAvkS/dENFUzNzvdr8OB9O//xN9LIEXK/Pr2gFt6CP6
F32dSSEyReQ/N72K93360pa06rebM3UMjrXPzYIjWtN9npiEYJvqgcxN+y4OaweW
u9TYVB8DJV9/HmH6AhJq1tm9tj2SIcswXzk9IMRHceFOW9RdfCOwifTFQuMhKMJl
S5CXnYU3rQCvqu/F1QIRc0LUzpr47Igv8QnTji8I+5PP6cSkwiENbW/hDzU+ojMl
HbhEDnzrV8mMJlo+fo8azxBsmg7PIMFUOBTk7823HbsQj/rUAdc2JFb6uU/9/osT
LLyabZ5ZZYBdFkeK66U5tlnryfsiEChBfq0gc7Z6xpbLzsDCJSiEZmwvtUXcG6L1
BopaJHhC2ua6ewDXHipWRHEMDrY+Mh3V7Lu3eW9MBoSJkW/5HZEqroYH5Ft+5Mja
0SiQGrJuDtKoh9YbHjH0dFIymGiWeiWhdrqzaBzTYIEbg+cMY0ZadjiK5yYUOrvI
QfQDlu/QthcPL5RoTSGb7h8xrza/JEn56mLBvJjfGBox0sWq1BnXhG17qu47DiyI
HRHDUEnPtukKzO3JZ5OPF9rbYU0eIEwvtPqmVaMCxTo8v/WWN3lITYJoIOc54GIB
z/CWBfTWveseNCgdms3++lPudwdcdqLonedje8LgBBtzxZmn1xDQL13tx2kvtPDw
HPXUfKcssZPAXqW8oc+mju494IiufVTjn+CLWoXs+9DtoKzJNDfUQ4tSVfBlRh2g
+rm5DZRT2KpuG0qJPm8HljFt7BEv73wmj2RIjozkC2MDQqOz9t+UH1OS+eOs8C+d
+ID7QpDSqxVxi6UB4CBex3Q/3ys1qNRKDrn+J7mrZNFE4/nsZ3RHRSZcK+8NGhRk
+cCtWJDjUy3YUhOeT1s7Kg9L5sHVBLliNIeJjOz7VXyYVNMM8eroP/xu/5RlZl9M
7wC2T0QQuV/Rf2xK+EzmB5OTYlB+kP7gqM8LG1ZGO3qveZ6QHiTpJ/XTNdKOBfBB
Lg481wy9KxijzFkNqJwGkx3j7P6GmL/TzbHGH8wrCcKYsodOlM4zhmSyF6nEQ1Yv
M1BiqVJpnu+iZsmnH2J32baqnkqFq1jAExu6gzzV0LSSqX9B8WoIvPFMechnFn3z
SUe/QJ7NHF8S9S0NucKJqfnT3FRhvEhaUXf/GVmUCusdfX1i5XZx/bi7Ggk+H16t
vqXrDZ9IgGU+FIluYY93JvDtMKZ3yTR23MwtdI2jQtHQ4+lQJl4Uou5BI6x5zw6V
X0hzwCvLrz8tu+1Ln3RtS7QvNHTQVR9QbZabl4w/C7KRtem5Lpn6a5Rl9KaValVO
Nm9b0kgHL1iD+lYycLzBhtCrSrYV8Et8nq99Tu0X9jUEASmIbkrK0KDpp+WHQsGM
3zzbonOwy94D275IRlPtVXEcHU/xlgKU6E8UoXsokW3ixLoE6oisU3EaxCqArYi5
Q8pl8Eib/EekgCmHf0ykhV1BbOrYwMzI27o98F+3YRIJH/qcbO4cA8fmWw5GE/vQ
hJ6pEtqfHsGVUUYbncHTy9YlckZ6zEUDUoigkkfo85+5j+mjGNf0IM+j4SlpdPJx
WGFVLcFCRuM0SZubK2Qjgu9Yh5dqOxaibrDGLCyBq0UVeVTURbt+C8bFbAlDtOoI
Ii+YqX1v6d25pagF2leJVdJxJFrOBSYK7qvJ9tcrW06b0B59oKDwFIR36/GL94w+
lY152M5ajyWJDSJtvU5rcrn49ZCEmBKSp9zzJ3DZRqLs/9zikCsajXrqsXxPD+eq
6AJUZN05wLhwWL/OhYgPYnkRSyu28Nc9ILAXcwvltiL8xVk1hQZ4QJ5Q4RDlS9mP
lxZpMO3ZowBemtP2wLJf+hNmMvwsfz/2eQ6dB+YyXs7yHiMDqHvQxiJQqcxosrbd
83/IyWVWgZNWxgU6nYAVO01/9yHWLRARoLL89FeZbO/8zZ/aDMii4fm+2JjUaBLA
XpIpH11qIVdbudRXzpi7hDjLlLbRiN2WH9CVuinof5kIX1L0VoAk8OlgLP28pBTS
d59Ym47wQqd4TcC8gJkOesNC1ANl82eiHOR/vo5k3xNXFezZuowLmRBtlHkED9Bm
/tkjbdj/n0K4ScS60d2nS+ySR6WStndfdnnL8BwomOkJhrrJP6LAC+IAXOC7oTv0
fzH1C4hB2mdiKhpNRBvYT+R2Urg5xqy56LnSgCn1wvNTyGF/pg0D5VlV0a3itx4Q
29/88m/7XZGsWmgAv4sdaqv7O52lSCJEUJJBFx/2WdXWB3ZxmU6cSRutkDpK14ds
OFhQJ9Vi/CZ9qtjrzUduzS2ozu1yJz/b4GJLejLsB+rZdxf7QgtWdk04bUxuiJVy
gUTtm5I4J0JhOyjE8herOxWHx7cqEI5B3X1YSc810KvhcCSyduEoixgcVcPn8Luy
kNwf2cO8On4MrSkyOgaOG9/mscS2podXz6g6UuAsM4zYBoLMw5qML8BFnAtVYFMz
cWHBtQ/cnxeytf+MywW6/LXIHfXh/62QluOvocwtirl7VWU4AQj9PtO6JjQShFpx
dEPwmx6lY1B+eS6aR5t1k7EntEsPVYw+593b+0mqWSADELCZfPfdAF1nyBzrIrYm
2yGfj9ZnGR03Bt/68R1xLzfQ4qKe9UmyFeMIj2M8KjOh3SPNU7lTgGuDlIdUbJ6P
Du+CrWs1oYOx65zh+omG2Mvee4Y4axaLpZzsNvOE5nJzo5IzQtiSC/T3H87w00KG
qgdNyGQun/9AHUq/KlBZB1GoZDdYOjW34ApBhxuFS7BMf9e7LTYFqOTttU6KVTCQ
QBN+Dvw9Aj46DpPCno+ZuocM3c/S6+SlHQfjt+o38eIr9fMxaaVMgkiIrl2HZT6P
ifqz0Sx5ERrEA6pPkEaoGuXCqxQSc/9Zhf4GYT4bgsjYlUrMF6pX8nS4Z/j8rvNc
FSP2/UsQRkRiGoc048FHZ02IoX3tvvNa6ih1Qhxpm20GDN4ezfzKaGO13TFL01tv
ykewjMbpi5ErXF1BRMVUk4cORAti/9OdLGYZNVAjBNBK8FQBld+Czi9v30R+Os/H
YBmB+llJ2oAh8VAXEiv+rXDoQnBx3JPWefjZUp79TfKf6rpsuvGb2awiSOE7lhWM
1Z0ZDW/xQJ2zpd8fvb9/vTuJQfaDPwkOz2YtwezwRo4kC5UyatWHPo6AWc/nKRxj
hCGagCIn09819dBkU7/R2o5LYy2Nu847xlGix+59LqQHzHC5klIM+Bz7+PBFnUFB
trDLgHrF0kwZ6kkdbcOJzlzq0HhlqDgG0375s87vEJtV+Ee+R2Sza1BGWA1NBHrl
9WxmPIxgO5fYf4tppt2luLhy+Jb0X3tfwkqKWd/4hy6JTONTR/OBqOm3RZKMnjrI
k/RvicWZL8EYoTjw0P/7tSFqMVIBGFLt0YJWE9wmzjI7SjmdJMBhfJZ/GnPnh+uJ
j4PxQ0UczMdJMznddeiJWvIa30R5OWg6SazifF4z4HkCOVg3CvZVYRuwkeyCg79N
z9cf3qQVLt/4QsGNn1dvtaM1y3GfGLyN3O35G7jC8WttJYUkjAW+tmcj3lHLIDsE
e9serQa6hK1Hjstv4HuNo5xF2Ah9ONTBMnG+gaQK5pUxvKfB5M5P1BZSQuwSvDSW
qIrm1S2Q0q96xsfDWaNB+C+I9FvnoSye6lGz2E7ulSrlFySwHyFq9TVPf20CORcJ
2sZnjrzRwTteeF9f40OSj0+EF8s0W+arvZfuKtKjDbnOiL1FBvK9eeBLnzltJCGp
BBYBylrcER+NbHTI56w3k733vWQB75P/LsI/ygUegWf89Fif5nJ8L370ygVc1BfS
+YPHsNBvvFZkeTAbldQ17hkQACaUogEiHlAQFc+6yyP78dxVnVqyOH8h7OErtoHI
WJ7y9ty2wcNori/OJyFQS8aaTib7TkobVPCZ1Xl9X6B0vsBHRwqDWZwZE0tit55z
9I5n1vw6h2RIJvTLh6Twei6Lkw+Vrr0wggymzVFgzfYWtiMOD7jmJ68G+DQO2iBs
J3HxJsi2KvQ81Hrdo4OJ+j6GEKfgzl+vigLVL0HgOVQJRXjHfMW1D0hb+UOxpp4o
9nRHXFz7s1KPOcFiLpt+4OGZCB+OyF4CajIPQRWiHV2iq0G7U9Vtw1pjQZl8/BoZ
eFvtYXcOnHVmBbzzKpW7sI/NY/67QxKzNz+fOOFj/RJ5gx4Vw83gIv/sTXXHx+ng
CNNXCZx6aeHqio83MSUjzGRy9xSFja/ltenfjQGfiziBwu9DwFlt7H2lIqNV79Bg
D9NzybMQFqcnO+Tk9mBJJU5QP8o/8Xzv4G7Rvrt8HfydmXHJgQiQ2Zp1FSzPQoJk
61qbN1ko1ufl1UOZ2XUiNa30rn0EtSg3L9FHy1ZIDOH9SFtZlVwOsjd4uwMU7DwL
kf9jBpgpyexyTk3po8j9l///GpUILrzD7KSPIaGYNXTTpY7pxoMjeaVVxVquGf7f
Y4V1x6oPQ3xqNYaePabZCWUV8ioQI+uJMo2nL6xnogpHCIiH8IJ57+IjXPqGoooE
ObX1F7+3Zaq0pTW604/tapfCHq08hcuzI3WQhVCHYmTTom/pA3eTI+ruYFsMaflH
RpQ7+a1fNRQ7liSP9Jo6757qBULa/+3HtpL5TTccBfpJXC6SK/j2qfPa8igd32ys
YtXdMh7nGL8nomSdBLy7uay5MkolYDXi+bg13+JRu5Z2LENfVsd6zbddgZTclfVs
kPEIwxlas90DiS52u0F1S+ze8p2JlCIS1WFfCv3acDT163STJOFsznDy4saulI8H
bSwwDDi1dHGAs7xArV/Mio5Fv1QyYqmUS1K/5+qKOmdJjtbPwQt5X+jqnSX/pB+A
sV91b+ccwHRF3f+u4bS5zFMsXgoUPQVrCcBYxLef29ov7NiCeUS2+AUfMD51mKpH
du6WSPKH7A27aLxwwEGTlvRM1eFgi/TMSAZnhx8J9Qmj0c5J79qbQTU828LvkFSB
xyqpuYQFjwC1qLw2AjZeHrF2MM7XKzG8n72g++Z3725edJd7r28BkUFTR6C6IBBM
AgD51hwE6C5szi1vaxu1Iq5h7oL6BCGwFrjaIXUiso59TS64QsZ7zRe7i/l0cUFB
zhHyVSc/pdGuZUO7w3CXGJzpZoK78M8gqQKmjpn5QA03GnG2Ub9T4kxrvTKsiWub
gF+W9H3/X9uXYh/GviJOAQzDvm9E+Ar7Ra4vsR6617/Xq9IROLOW+UjOtAwzUQw3
dB7ry/mLJ9LSAMkd9Gd5jJlQsxKZpLyT6HAtWcIGDVI7cQna9Yu0zGPCvoq+vmxf
PdFr0P1BxL+w6PqvfaaMu5d6t3RH03UyJdxf8lr4S5pYjkzputlOcKuR345oSeBM
TAyMuSwAmrrPLpMjsJ/aPxG86Vjd9qgWASQcpqM/gki4+wjj7r/yuLJr4chHM2CJ
xuIYvfVu6d7joJTaw+VNtqfTg514J+1r7bYgCxV+IZ9OONXmR7OPmXweB3Vb+iJa
DIuZE0SUDJI2AFwaPpXQ//ltcKn1KKMmerXK19ft9QyppwH8oyvDVV8WWvozxhb2
5EMxJEkENwkBHDBQ0p3AbfyAm68qyTfilz2Yeisw5J0aE9K2Rfqg46k1JeyWZkkf
ZCAv4gnPUJXqPEzfr5FOA+XxNxoaBZVWDXRE4o7uP3J5tiFEHBXUFbZ7Uk+fzd+p
gPppS0lDoeBQWakTzcT7ZVzpznmdZPiEARfbaC5eL7YkqVewIVJWFbOd7o1YJaJS
YtpkviJZ+B/dUodfrqwZ61b0ofUtOH3bgNmswAs+HiGk1axEhx4ZiaCIcuRVhJfS
QjIyQgIqAJIwpKQeO3JqV0X8pynRBhFFNOOfjgL2Rvu377NQ6v/rEIm7+hse1iWp
C87F3BE4nt/Dwv++Mzkoona6TwB4AuqdlZ8E5YCs4uvuac1EC6IJh9uKD7Eyze/9
gw0xIx9E9ZufA3qTA/3HnYLvhGI7li1UJhQXEwf7heCb9p90SaQrRsYmV+XQr1I+
K/mto4SVvkHS8d+p0w+awKqtcM4XSYS7iUYW1ZuB3Yk6nAYY4YE0Dsm974Oqj1KH
DlntNeDcKuBy2sSQBZz2oQxys7zVkOI3wbTjTDEgyTVaTZESZ3G1aH6OoySMm0pt
1Y66qHU3pPLSXmGixeidyoVg/u9H7uZrQJHpWMcdWAHdNbXLoQPBCjchLDddvt9J
I9D4kd04pkpEIuYQ7+mwqvGQKvb+sJvZYKH/LMwaK7AfqVizOIUcauYmMiTloMjt
1N5FOYGBmqHWkfnmQMMffgbTpXo3wyLr/79n5oG5GloxOlG9JFG8uZ+732A1xCtH
MBAiTi9vVzb17HIf40nueJmpqctddLYeoSjts1lNSgF4LGrxjg1qWzrmDjJm7N30
4YTh1Fjv+lwZm7OEcJLbo99uKqrLmUE3TiektyoTAGTFJYE2LFgKTIhK62xObV/M
vAsFlArI4kmp2fyBE6wudSPQd4IGsolxGuDQ2HvFDszTwk7tMHoDZF/wIOk2E3Vl
YNt1flZo4RkdjMPsRqIgSDjHKpecJhxKdEzQzF274wunhfy61IgPBETCBU8OX6jK
55Q5sLclrip2rx8Tv2/as8VF+89XDLnTzTv1Mbm0tZJlJuzHocZagE+DBoSaNjGu
Xz/lrW7AMGy4c2uxWL6vY1S5r5QgAV43XxtlR0z7ULMsO00hu3cyo6+A3DSWBQoR
bf1GJD4CTakskh0DWWhAvI+UErz1ncVb1zM+3oEec1ByHk3tRODOTMmOcODeLhhn
m0zC9Aa2El6JbeNAziA65mrdextKBF1G7oPm6LJyk0hceUrUrdLH/73NY9ZhO6If
+kP/RWx/5z68NITAMBphxxPpkdB4CzMW6VKpjo7CpCYmE6hEBrm+zofbvFHFG02z
VKeP/6tKEd8BiXOOuxiQ2mhsfe8B3j8LtLQK6LMvb/7K1Y8NiPIZxpP4EXcLGGdy
rSCBH11xRIfyI7ZcQgK/lhbbaLDQHdwUH9SH/fH6ARjkcZEGSj9jfA4wfSueyeWO
1ki0C/gto6G7lLABEhXuFtOnQKicRifRJbf0+gG5peatjH70vejrgRfGAP6BI2oD
obfhTBlRp0Z8ojlxAma4+L8so4xVtToS7shmT9tkdY+WaGFtgC0AeLV7Svo+7/TL
CPS6C7NzZKMYCbJmpZVbDNB6AeYry7Ysvf3GNgluhne9YCzs0KufZI9HeZJeKWrY
YWJU+h7Dlguv9K1yb25GK2oTgRiT3f3nsMkntSzYm/eVDE+OpGsoCq9y62YaMj7E
Y4ay0EkprTIalItyNMk4zoXj6irN/+C51IfBqOrhK6yXcX7chDtFdrNUJLH7f2uB
2QN32j42JEs+OKY9DMu5JXe0uLLltricQfWpN5swopiyujVxsBOKzQGDZl8Ryd4N
CQO/zHM4hatAGLSH0R64dAXCef/LUq4bn41f2OLKv9TZXzZLaO0XZ9r2DjDRLgrt
Y5gCA2VVUjrrHfwoygZ/guK7J4w0JlAVM3jIzxdgMMbbb76DsYuUKudW2iuAdKTK
oIrAbKHu6AWuiyCHYDRjQ1klzeW11DFLjuMD5/ZpIMJhmViYlOKsg0/ONwRCqXLl
oBYP8g6Q6Azm1/d5RX2tTg==
`pragma protect end_protected
