// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:02 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kZJMqHBzzCc5UjG+TM+JCSkI19dNdLVmq2Vb8dtrj+DIFTKxZzeLXuW0qwVFI+SD
T6/U3bqUPQVQcLYDLLNZCsqhR4O7D3zb/0y816Sady3CUyNfswoNszbYlR1YLZ3b
dGAB7DcqE8D7jn6AvAvaXT3TY+LFr2W06aQLZnJzMvQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5664)
m+DKqQ+4Pso4VzRkZ0909GiwHkxbNFZB8aFW/ArqS4Esbl6R2PCTQLk0CG0Aik2I
L3xLJUG+4uhx0sQYiqQLOrlqVCCXEkaR5+dCrbXhbfQVzYY/uhqusntKcWYiY+TT
ndUzqa7qwGlcYodyJOGQ9ShVy9ioUajCevsQb3H31nUIOFQDeacogLoErA5UYjAs
NJrpujMJnH4Bt8EhoxiqxkNq7KaSsdRM/VQDOTROdAdAyO7q7nDJOdx9Xm97oGIB
2hunxiu0qMcthCvEvLDv/913SafY6jYM54XxF7MqvBf6HAH4H78ajU6/qKWonH7K
ykfDIrmNiVJ0UyqJPozSGqdIrtgyoiP406rJI/BpH9UQPUbHJBX2qjWbiIck6FqX
WHnffYggPoOQwEBO0RSnYu9yFk0Pc0kBLqHiDpnPRC0/d90pkVbmkB0Ue+wPiri+
u02VzWbaO68mWg6deEDrTdiH1CmcGYgPC03OM3takv4LaOQbSiUaut0huzltOWXt
koyptC05o/ZmnT9VsxniIVCPGRT1I7mvWVX0WZLM4FydwQMTJFKVURl8cm/U2dph
koDr5rIzvZFfSMHQti489aKM6KTkNhduwLJipyZFCoUovG50lFLHUt2gorJkeRPb
kLyg3oAQ3t0vYIFlT/+pJCyOu2yqRx5PeXihr/dZi8Rw5H3YTIQJaZqbz6lFBKm1
TdDDDd/88GHQF/BI/cVsy806Pqhexsr9bEmTdgaUuPvS17v0uyQAuF0lERo6pe6I
B9LkXfCbkTxNIK40VzV4QWAdHOGIRhUuuaF1Pek1MSWqYQd0mafug0YJSMrAZors
unIvpubVSiriZHxslRDi5Q6RLcOJNxJ4XGXVWvhACXPEnsVvB3I71RSX53Cd0hL8
q1sxT91v5RC3cOiadNAcSIG5xEusZig9dD8gPupppJG7eToE97tDJLcf/y5O5JCs
SeLGZgOpnvYoXvsvhUu/lRlNcQ/l6vHeCPgU65QMXF3/zor3FHvrafBH5Z2VVP9h
wCB9Zg7oStgezqN8ueCEOxB/GS5jTo3F/AZtBBsA6/w7boI+peOfLYzSMWHPTh01
Z/me//JypHtTMi3DDtE1tLQUXYTaWhcqBidKOt4lQoTvBNSKaJ1+370TnuoUqHRf
hNFxboKqU8ios4FJpcI3qy0HrnFnqbqOH1v4wleZsPtHsimpFgz3bIy2Eu9GRkjv
4K8VOVl7IZ4WNo0UviaGRizNq0uvbJ92jK7kXZR3PuIhYFAsOwMTx5MdjSbkxt2x
gHLnaU3zZ5xeEzKQA+/WP4Xk3cpVAfnu7fTZ2RUEzfyqejbDXruVWz3sudZqqMBr
3y27hPFORTezYYBQVG+2AJ3sxGjq9Ami2cF365muCYym5I3hi7AqH8ddXsW33gX9
K/+7epS1omZ7Xd6fJZuwC7tjlNLX83xOjNAyuzXBg2r/TiFNoJkaihhd01LRnhj9
37iM3sGRn9QIC5sGjrG872mIc4PDUXBWLZh29ectxZ3Yo+M10n3kgf1SUZFX7qT0
nNChVlPYL33+SijKSNj+ARfKoFlz8fCnx2ksS4MwkPp1QlNC4CciymDUVUcbysJS
+biF/JkLbkOn9N5MjNNT3ucsKoFLL04V0U6BQSj8lsIIZqEiTrf/uE/R6kAU+iYv
MlYx/h0o4ce5Czs27QJW2ukSh5kaLifJpQH0a1kzGQwb0dyASDn5G54AKjf4gQXR
GaSYqIna/F2uqDeeR7o4hjeFYwf75FJNMkolB2I1d4fAo235YqysPg/8UuGeBFfp
cTTcTDgTcFUqiTL36ylTC7jN8LFJPk3h2zQUU3dLPTb8JJuTwj/HFeae6snLnkIT
7iYJJBlwpwVJFhBB1F4FmaQbmis8Qa0AxaEkTtp1E7l8bDLCWkO7dlk89X0Ysrk3
Z0HeWxUT4AB/gc64p4MFiXMk4ohAG+CDXlUoSvyhDpm0UJbMLfwX3gxLK1D0EXOh
WVKPq5b6EKuoMlFaGyiQsLuBnr+iGMb3EZBTcsV8GFQYtaBezyueN62OOJ9XgkTi
INgX4kxtwaE5vW8D0uTEIspJskIwk9thVHL5n1Ahz7jb2XJv+5G9HCzTeMKCCrfU
SLdGIyLi6YGQ8YDxTC39aIidy7yD1WUICPXCywClCykAmumXFjPI4rD9GBu1AZ7M
r5C+89q453vD92A3GBNmCEygyU7AKLCptTPx20vsmJwL8rVQ0J/3IaN0NX2FxBqV
7Yv88S6L4w8Ak3mpZ8aRA6mLkVIuusW/3ZRtd6TUEuDmdw0RKTxvB39NSRZwciO8
qvf802qwhV44yg7yisLLIuT6h0BMueGodST2Ls1VG9WwEkdcmuGOtuW/sA208Oqg
C4Obb1G4aGlc9JHMcPz3TdXUuAB6Lz6edUFQCNccce18ZJUVVQ1m2nWvJ9dhV7Fu
7aydGoe4Is5/LQvbHE6gP/T/Nhq0vqTxLpt9W1zRxNRgwIzC30BpaMESKNjqZpN0
c2dtjuyqjwnnaaOlKYJbvRYrdKp63w2cA2o8aZbziMA8L86MXC5+B+73uOsDCdrO
FNWyIMFw3PkoeoKg2jmrw1F6BV9xKpmg8CP9zG0Z6oUvo8lXJfJ/rkWGgCe5NzHe
vCTyU30wRhEH9xa7OaG31Kz2b0XFGF9g/bsrL2aZwaWr9wV6MdS49JmgzNxdFUs3
t0fuVKwRP4jv4do5UEd8Lppp4GL8EB0k/VWoa6G4/l06vFeDuR1ktNsHttiwpPPU
RG2i8mS66M1iFed8KrH0SUksCyoabwsGLROebRo52wsAM8Xe8GCqzHxFwtWzhU27
80yWw9Nbr8DvMxRHp2Ea8nltu98kQNmbq6Uo5cFVcjQIzWCPTn+VENcYU6dqwchY
6ZlIn1JQuwNtSHxc/hfktcgcFxFx4wt/OoBbwMaPQUoTtbXA9ELaCHMotrgJA2R6
T3nsHUpHRXJtPOGG90mh0BTfLfkIOuNlR56Ab05FasP02CuFwesCKWnuIUw1wEVD
Z5hj2kr/u3kyyWtqDW8sb7xZ6mPW1dflEnq5TL+/OuJHwS4i4PJzkbRgd/0HsD5e
VndgJv8qFy31WAdNc3lLhNpXLYjB0HABjpNFvnLZquBqVfkZeZ3yo/CbzttkYsBo
PPt6gPlhTeHNVYsabu1iW10qNpxPhg/3KNHuVWVVE/a2b+4GdBaL1uCE9zSvE0Bm
zw3IEt9odOmygz8jBUtW5imhlhaV0+93OEoNQZ8YfiaoxEDqtqThSdo0eLwqVPgF
t83BH6EnWeRJaaCJk8RsgFiIN35AAuLATVknAZZPeIRTVTbi3/YLsu4+vqYCXWV5
K557hSym4Dbu4QwPAhxr0EXUcecQxbVb2DRDfXornfaQndenraqJowT8zXWwpoC/
upjbdEBTCmLJL+/mZyApw6m6WIC602GiIiOhjtBvIND0tRWjJvNKF7ZJX7E0p1ci
65yBbpIKomX43cFzUsm3lWNtxYzdih2nfyN2J6oKUeqBEE9Xj4Rjj6v6pJtk1vUN
0d2tAO4sYd4Ual5ufhzhbZDNP19SpkpQ7Ygam23tthOFNdJP+6cKpfsvX8P/o5Nt
/d7nJsoMWNZAAZ2ZNoDQw0xziVSlETMe9wuX3/nUd0STrswQwHnVnnQvvKab/N7J
ouWCpsYUfSFV60hBWpK6Knk3VpjLF+76HJ9fWbtB+lZGfK8oODb1fX4wy5aIHVJw
u5rMtaRY3p6vuYS2+2SJBXsr5kTOJfmWysmrSmtgWkX5ZQYrK+9O98bNwBilImss
cXmQbTrjnpLPeHt4QZ12IRH7g5RrzPGkoInhXZbxCHJ2X8W1mwahWEWLMd7/tFpr
72qmIklXxMatxfbd8hLeQCxznIn4AOZKjXsp+d1jFX15FE9FY8fVdZANkl68pBiR
L/gf/JYX8zUYixvt1NvJbx7lfsNlNHmYc480tS6E7IbMWENlTadCDLMA5Tl4XMSN
51dL2K+r8ffHW+jvkhiSvkFeT/a7SS0ELWtIlYgjROiSPkyQXcUuWbDIAORdUgwp
yxI5o+jC2E2MbNuXzFn/NwSS9NOGhwNhRlN24xNh/zB4zfrx2Yk8/Q12CE+OiKmp
CfFHmU4hAv4QQviQcbFzC5zHpE2sNiMqX9H/PUuOxNiSOxxpLOPUQfTToh2oVN7/
iPfDTdtJ5xsH/I/U3KNyHqA43DSPLKIcQJysfq4g8sVkBFzJv4KUgkbhkJjq5cdf
V9YHP8kr1Qjks3m+PDs8Sy9lrXSUknTE715l6abXt/Ufi8giLF4uMvV3XuqT6P7A
ou5dOrBM2XuD82/PhzL+iUrOHFMWw+YEejX9SE40zZlFHwO2vW8C7J52eoMSTYQ1
qTf2PcV31103oQWDTAoM6FhJkgIV3w2fx874AEtHc49VTWVeKiu9LjQblnX8OjFx
vJGxr1kaJqWYfHRDtpm52brr6AlUqSpIzx3vCSk3GcaTx5QPgNiOcsK1Z382Vg+t
XaFZlirqIh2ZWqH8qLvkp6SfY3mDObNcei9Z7FDIL+9V5Yz+p7enAZ7fFBu5ItS2
QSKY87cIpgiiKREIvRuPF4yAHJCV96nO/tykxFs0qL5stt+c7GD1aSEyVy2xm0Bd
Np2oIFBU8Fmjd47toDonc86dO1r28Iie5veaH3/rDzDKuxKJnfQLnJPkaXPhBgCw
FCbq4zwySzjgIV2Ejab/IPtY6IwLpKhM3baA2n498aIdHamvN2zNLEs/i2f2JaoA
Wjp3eqCfqKkTfJDZwlblxUjnZfbdLZbX8hIF9M3L8x064dB9GTzyXs9Nhyv3IcKH
Xr+Yeb4Y06P3Jji7KL9IK7OiaEUg2ODENL66ND/2hO1WQkbsqC+VjYanC0rAwMW+
ScnvRxuidjcFohtHxLZv433fr0VqaRf5uX6sr1ITHobUcriiSBzV2HqTawZrStTP
AfsDOztRRcP1eYlRcRaymmJHFxzRiGrvzwPkfk5GseADqmVJAcArQ564yLK+nVwf
N9RUFv38M3pHCQZF9aBqsgG5bsTWF8dBpRfh1Laq6nFsciw59OL9yZcz+zhyL9tt
FqtyeFzzcj9jHOPedEBlm7/6Mw9sathBm4UWAHmCzGWhWATbVL93T9CozH8gZ9xb
b4ncGPoE6UqJ3ivAeCHX40CUiUV5ofmxUhmA8xBiOUS5flimAFKomIzxcGkQtIyK
MXmMSmoeUkpTfQItW1zcz1n7S/aBN/iFsvB+wP5gpWocggyXSk6dKkAw3vsE76ER
BjjrUpwJUHOSRabU7wkn9zIOYirJFdB2rKKojX9UHrAJn8qCFjm70vxoAwAtQk/T
naKW4a1h0Ox1ZAIz4HGNdHwCFjN+mzGj+XZnNVOMNQU5pN6Zkp6/hU7HZ5zx+qwQ
bNg4TKjnWL38horLa+JsLJ4o1Qlgfc0MupBIzpIgtsihtKZgTP9hCOF0LQ5UA6LW
zEcEMHH9QxIloe3PUTQYfmQVxcrA22s8hgGv+Bqxujji86+4jf9YO0RbiATI70oj
xj/V8uHSPY7G2AB2CZg7YIA/Y+6arNGyPOGJRBoOp4DfrGpsYutHVNTYpcGNKjK8
WFowzF3S9ml2GcZKFCnMpprEhv66L5BcRkkFOHrhewnUIRlYhyNx/YgiXJEY7fy1
KMj86m/n2DJGLRw1raBpWbkR/VjJ1ZrHEXZWBAKEFM9gdbELzjNS1yy3jyJeJetE
isFE+r9bpqPHrkAZIi/WqbP0XiWIMz+hnQgelgakkefh/b3eLgHXjKx32grHKzrp
DqBt/tR9gqZUhugdotWnQB56GD0HRlgm5zFNSDVseVBgSbfswYlua3NpujTa2jgr
+B5rEoSHk2CveMSCKL042xMU0VlrF/l7PFSpRoIZJM4a6mRY1g0E7keaNI5x94eH
WJAu+RKdtfORAC1cC3iGCozEzR6/Yagd/gl1pwSYUFbdFlW/ra5P91XlKJN+QXuz
aHEUpiyrHsu7rUjkWXtqMBPnG5DBNhIC9F1Ar0Df8tF4C41LmJ1H0Fe9LoeiOOr4
rlKarpqzrbClpChLOKrjzo3jt5R3mCOasGaCI6mfEatUSozD9ajAjgi/RqIWVvu+
sVCe6UGRp18Q/CwywigLS7IX/087ELhCD+p1U1ot42DTy4WGssdp07nG/+Ieqbu2
Z8/L96vTm3pi3kQ2B2lZfcW1XZVjF/L2Gp0T2XgRUO0RIL9GS35s9xen9bQtCrsU
29QoSZyxe0yq8vzIx37xMb+uryoE+Pp+8tMBJkcjG2Srun7ou41+la8qZYWbmwpp
DSbFVVBGtWN/in3I1g3nqRT6xX38gE3CDksHcmFb4YFi2C8zV5TgWz2cS81Az6SH
4URqoN9HR9H1EhqLmP/gJorD4oqWv3sTXHU+etdJm21NqoUw4W4nNgZiFOSDWCm1
5nIrsLETOqscN5Mb6jj4eQjSicSe9WV2F+2OXfwCO58p3QISmp1YdQpyeSFLaY/P
0GKgTlpZv/S9uN2uKzMn7j7GbrnqVTAiTcRdUgkZMh0+KNDaB1mVnkXw7HVYw5Rz
OEJK+HR2ll64E26OvxCM06oRgGX8UCLZnqbETfgDrjaHRQJQZSJp/DD5UQ9AmUoR
EzV989x7MRNP+bHq18AyTJ7cEDbPlLgNn+z2YigAmLHQdcizbQge6ZNAWiqVPuIJ
Gs6xdDnq9ZNYFCuoWPSebFHFHccSY/xyfgEbsA0+l1kgKasT8bxEesAD8i1JHC2z
ouiLL+ogz4oJCu4kv7DHwi4mx2dScHvVhsIGJj7G1OTFONpV3ww93l6YM0/W42XG
Y+P5VZDhqAdW76cL0YjqjmvPJsJ9mJoZL1TfQJ9QY4LtYXjVz2ia+Pr4CrkZPgvA
ASWFQ1A69pHb26tPLSZXpSFPOZDuYQkPijtuFhHlSKlH+Fxf9gp/ZRTygwVYSnL3
Vr25t3YDtziGiD8u/s0/VHdYaJ7v3/8qUlMGQWN6YFAIebREkqmRik/Ekt1M+Gl+
d2lha5epOM5hnDNPtuUeJVGduYF1iuXkBwumE3Vy2AJShAC+HnWg/qbADElDivmG
CR1bOqOqdAScGLGK/VdnVDbce73vl7JY8dpFIkNK0+dvagGhL8nQzveVxjqaSR9e
zSPbgzkGdhj4cHlta1a3LLXXBM0zvTBE3gul95kzhMwwulu5oEyqjt13t75gbrDa
UHKfQNYGXzs7dlewJJVf0rXuTjMs/vSKr08eYOnK22N84ZxxUel2dTc7VxxvEzob
z7z2rKnj+m0Dkd71+eAAfsYI4kSUh02CLOorM6JElKwyGjkmICHu+iHsR7LqGHtX
Dge4YizA55lQIbHMDZk7Ru0rVCB2qrvoM4yVPPLNK+v2gqMSGSjor1YTZmw7kZ3+
gByGEMDwtfCsmv6ev/kvEMMa4rlbDj7SkTUTA0L8MCvAPkXVzbbSeYdH0xxn4Jq5
1VqBdpvX3FPH8Ao81dIvHbNDRrNt/O7srqix+uA28lU+PYj6k0jRBFzUORB7iY4z
lyVehnUSMZuXk4nYBvbCtFRrp0ZZRhbNRxyHuQIHdtK4M3GH/6toJLwR5j24AQiE
`pragma protect end_protected
