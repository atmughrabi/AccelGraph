// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U6r9lcav/7Up3btmEy/qncKSdHqevyFerqnS58/WMZWH1TU4JjHKNgD/VUNI+Rqn
4QEv9mE5bMaWxqBiU/iP+mnOoN0T5yEZCHVjuKswVxHTKNZCafUpAD8kUTl0wfJQ
1J32oE857v/5/WCRdXyZYRMymKxU0BSc40TR+5LcqEo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5664)
roTP/FGTcc0UDTWjWGNDH4o/ym/SXNunkfxvvnoqXlSGLKbGRIyIFr+K0Zm0ErRp
yEmiBYzxMj3vviiqo4zdQ+1NJ+arsUWIdBiOSylJ5zg9us2zkR+9GPVlTojW4xg1
anjfYLRL8VMaXeqTAyCR8McUyKqSV6ffhN4AgPzcfxKFUxnrxtDe5SUO+sovepjc
a4yHbjCIMNk43gPeIPnWFvsbMjIsUbklmoN/NjHLPAK1rgxABPidQl6BLpxBaOQg
xdD+VC0XqmnB608Hlq3ye3UDjM3YEp1PP3WPMsteFxV+CQY4senVZVnZI9STUVyh
Cuy6edvh5u0mmvkgCUIbWXRGsf1GWMTfQWAxTRLOHcvDHqLSWXR7UPe151U05JYB
sVZNvaaTGSF8UONlM3Fpbp3RkCaYv/CYb0wjZWC2Y4t4U+aNzSH35Nw3lcMzPe4f
W2y3j6bsUzI2kWP+gDvpeVi2vvQ14jK9frRzyCEGrXo8H4flQ6jZ+HS10LIePfmB
8eFqSejtLrSJO7eB5NHQI8smz/RJW5qphjWMWbB++YXis3cIsmLLgUGtzv+5dQ+I
s6bZHo4T8SvTbuZlR5r/RYHnTXmPhHCNGF3/8ASXQA4XVn+qP+5LxpCSSQpCr6mE
ErRgC1yjasiCXunmFFopHlzPtl/p+1SRoKNQPPJ1uEtcGjlYlGI3SsSDyke3gfUE
Ov5H8ZF/+Fl5vnnY69t6rc4x8SFsv7dAQz362iGw1rm4ONlJwgxHvBr4CByjKyfF
RA2Ud0c7JJXWqZ4emdlXJgdOEL66ef+r76ZQ5rYy26K5Pke+CMSpNnnuDLSHpyY/
JIKLS+MtZ0UCU4JAq+d3DZkpDTkr84iBS4HhVRGtqyqMGTLLI6WtM78vvfrtKMQO
85+aEzB0co16gqvNw0XUXgov/mKtOS9h2WTBK9m4e60GaaBeuoSXkqGxwWPbhWhZ
6M1RCZnioMmORDHeNSNvEiOrgTu3H/gTNPyKSK1kq8Ktd2+w/yj8rHyKuS1n7NNJ
uMeoQK0X2yWnWIRyRdGLijEHKm8/elpG0vY6zqzVqAquGzurCwI4TtfBJdyfc64d
LJK+PEkjbda0xxdztpT/Tzbyty0UqzyLG9kHQnX7hg6CTXZSJ02mUzYRcc9XCbPn
z3j3OAkZ6QKoPvIVjLfR7HnExiI+1w5k4pc48W7ROZSb9/7mXRDQHrZfPqE6GGEK
vMhi7IHDN+p1C8YNdgEmpY9zGjHY/Bd5YGSQHNgBnBZn7K5XvXoqgMdAVb8GlTny
Dhtp2Xg+rgdcds0uKvgJ5P79I22zKvaj0LOFwPIT6Ct7TSYka/TpxtHz1ubF3EuX
Hq+d4rPJ9pOxTvaV36vJPomWWzXwo92aBQUWSoQxyznGK/ADLDDhlXJTvb+zJO3E
qMYDwLLzpfy4NBUW3RJ7I3cj9hlDS6cHHspu4QH10fgoDmRmRHLSYDgO15+/P6tE
/UeUltMGGhyOGswt2YgHI3AXhlHMyDYcGW8H0MSvMyXMUuHyjXq3gtEc3H8VP5HR
cS3oQ1DnMVxR3VW9FnTTfi3wzALCTCVwGA49hyz+B0koFlEwXvwD3h2EwpaqW6o9
36CD9XlANKMiyYn8Y8Oh9q8klh3/g/Vt9U7hAxzOvkjOSailikTDvPnMHTq16J2u
vRXVepQ5a19NRHw0uJnrjT/c0csaEzJw+woj3mfAwv2eqwevLv08CgEueQ83scrm
8e14aYGz93tjKSUMkorr8Q0c9H6nlgk/X/Qz0gNDGZKphanhFYk6ZPxpwbQ6YKpF
y9g5YW2tcLla8jA/Mf6R2yc0EepzuMo74apYmaZwk6R2T84iRzCybAhMH67vmc1x
O15L/jrJqw8VXZgChClZhvYneE90c8v4wppiltg4poNpi+BqEmwJ2+L/BTs2wX+M
zLXITWELvbHXYusZtl/zpQUxHfZWtTvmLrRsnAlsOdDX7Z4R+myLVLU5urdT+kAa
aPZd/FoN8DnK8NdLHHyajCKuh8a/V4mAt2TC9/bS1LgdQZPX/0U0cJkfM2ofzltd
oR9KFGBqeIQH/nK1VGJwj331Pzh8JhM21fz8OYkQH0ie9XW9BKL1DjAKXFCjV/xS
TURKCNOrqTtxKdH1R3HXZaCOJ11seANSpuZtvbZxNHHe3zfeo49ez3YaYAZsGqqx
FioJgHYCpJKdY8pq+LQJ46zY7X8m+glEBkQyiC/u76QQK7/35PX0rqOKxVVKyQrM
azTTYTd8iDAIhq6/M0K2KwMLxNtTK43XGxHTFir9rQ5j6A/xesLUwgQb9SGeD8l2
Otf+Pvq1fKbygFwjmKdMaSZ3hdYR94y0evwCXLSVLvMrETzHb5Yma113su3tnvZ1
1p3TnGHOMDrqF2wGEXkXVyUwrTE1wbFh2I5yWThzRH6+KYJ4n7Nf/AGudBBaJqVi
obd0m5+0L7fRqsa3ZMyWYbjLPSIpPSRG0rs4hzQLwViRFt1p9d2r8Jyn34akFWlX
oQPeCekeUDcc5x7zoebsXT2cvFjv/YaGlFCfxQouVH4iHbG0cUB95oAjiruQztiR
9A5uONc//yvsQg8W7+1ygob5kfjc1kv5YWrjqlWvde/8tyhxGbjcox3UY54ePEDM
sz8YGKHTSpSXYxOFBN3gn6FlfzQsTIA9YFuBI+sKHHYm273iB44x7HFplKmuzh2H
KBuCaZ4vJwY/97W6oxL2j62VElQPUlfQo73wP2P+uyG8rioB1PiZ5ABPbldifgmv
Jid4Crc9sqqkXTEHLzFLnGMDjFsCMkt718Qg8ZVzh9/pfFwmaA6LZ1SqKrLvfq2P
JoyOS7MnMC30IdJIkhJKtvquywls5mCBnIGj3m5J9mNSJgKSMSIeMltASTbO0Hl2
CuEiTVPn5eyW1F/WPf4YYVi+fculc73IZ+vgAcR+O0E35gtoSX1tJ7ZmVUVIjvxP
X323PrxY8SNet8DNckV8tyOTy9CNjvN2UnEuFcX+wEMeRn99eeGQPqoYPir0w5V1
Ix+s8AnZz715/dP29nFfkhmLob3O7wt33rffQp5vGsA1x6KfmfcpY4IZPNlNVqN9
nptDEHdhlTdN6HtI5RHLLIS4TL0m5mtENh2gDBFFIzdSmUxvDaCI7sBRzGXHDFss
mPrCNRDsCSqUnbFU6+rTek+fJ8c0YWFE+CATfPAsQSvZSOYyUdUyk21Ut/tX6/Uc
bXFcPuQ152Kw2VZBhp3qZDzhBX5mYR2akysj+XxesB/RmcK7vjG4TQv64c/p314I
cP/rKkrf+KIsG3InQokC6ujuHPC5ZpGnYnbz1nLEpSatFPySStJohbOnvvPOwraY
hGSJBxS27+eIJhj7cwYOPoXi73WUo0EH4IN8A52hOSgIVwXJ7UDQ2Mya3OMCFFxS
kLz/jC78cA8bn9/fEFFs7EKN4h0y80ZSmk4dUshyz+ukqme/lyrwPPgHe1CrA5af
s/fh01taAVZInD0mG2qyNgGGXgKWe85KmjSgDvqqhyvQ0La892pefd44DlRa8y4s
tk1Bl1DJgcUMXqQSJXh6WrrGZWpRKY8dwMRQI9V8yxziLFh9xJrQ6PJOFHiuJ3so
hEJ4TkHigHHpkZfHs5Aiv2N/kTmI/XyLK2YDXOGQzHO2HUf5OFvSgrpd5Y43tb/4
QlSj60qgnJoKWEm2kVAVtRWCYaJUZ9wMN4NtR0D50RoV/o8pEyamk2xCKRATSiIH
joQc01KH8mz2ygTyM6jKmRxEivrSEs6a+LHhYnJQ70VVLFwZtXm1Cubajr+Shvfs
0HWKRkpRQghheAOoH/L3XFoGiwn5rIYYxuxZm1yE4hxBRK6uLF4x2nssy7ZzZuus
s9HNbnSFTRnxiGSVYLFRSKrZmGk8bVUFEL8h3sv+ZM82ndJy49OgBA1cNGrfGc9f
YJsdTs2yBKm6mPPJZV5J/RYoh1m13nPXaxXh1gCFs5angtTHQC0vecJyXkDPhNUX
7bvV8n6tw9ZNgC3iLf+EpmZXyxUAw/KNLNBKFdMbjMLhlX3qb8hKyxMHwk8beAv9
YrGTc4VJAc1iuxFcTH6DsjkcuI8ZraiMD2u14iLnR3HIZBs5pDJQjAKmQ5gxuDnK
i/RCPTsg9hicwjxrcwx/sAO9VACKnerukX99HMNHObctqIujzyHR9eVeyFQh97br
vFSzD767+kmNyIn5MtcgRvcny6g03snGue+QIY1mvNL7n4mUQZg1oLHeU4SjSj2u
AwQSJvxLgn6T/hrSu57GR0CWrthDtgn0677UTAoPIBHTvscU2L3NUhggXnnIdTsS
bDk5NlLWZRzQqnT8SYcX2CcB71fCThDhAduUW2EfNL5a0MhyZjKZg2ymwh6ZfZVM
r1rVTvNgP91s43I66oGohewdCfwU7OS0SPeBTzCnO1NLG2KhfNUnqtwLy9csnxqD
WX3dwGAwmHCiKlXK6t/hi368oSa8JOmVHY5jYHJm407gpwxitNM+jw3WUU6hfWra
97jwZyip+169AU95GUbzhwnNrqt4HAPhb+efqcVho1BqhFZKpa/TfM91u9Mn6jqX
S2DjvPS9BCQP9eOmIHey8JkJsVNFysP4BlBAxjEip7u6qCnRmBmuaNUoq5rgSu1y
GGAA5lBz2/PvScOx5rE0x+1jjH7t2fZTt2pKsb+Q14euWVniACiRe1yM2jWf1ZLs
4KVHis0f36t2CYrDmP9po6wWYka2uVZEFx+cAd+6HPqEYTGQ1be4sOydW8i6FjGG
2dAxYulz5nkiIRq6EB1rYpUrcLGPihczwr+bsvk3m3Ymam9zdzUb9IZxWSIeYZfY
b0o5CczJYpKmBKhXi1TgT5GuRjSZPkevR3+Fx8AYBIMFr+4cLcA9zNu0emU7Uyt+
IBze/T2ZXj16I3QdJVaG6RcdatBtC6Pb15mVeB4xSGZnCPM5Rb0BbKzWn4zuBBS+
tEq4QJXNGP9/RlboMXHG+jav4mRteIs73oBlKFe0dVrADN7yi02RkBMk0xyd2OZD
QjtWF8HjGPmWb+8YXOTo41kGh44EqIoWLbO6od326a9xIKJTelLx6iaxvbEJ71kB
Lt2OEJykzWDGnPsXVnBHGadzkjF1mMXIb6junz8E/TJcWuBRiSdzDOcLUfj4jdjK
yC04mxCvGO3LxrHhybK1RyUOmogRMpCc9TaUnH02LrnrHGzMbTNjT53KoKU4eQ0F
t5ZI+mI5JqHAm5CwnznL8NO9h1kvdmGe/Piwnl/nCNvmZMfl5ny7ETZK2C0mFLhn
BGoUYa13CWAsBtvV33qCSv2sLbzcvCXkJFDqzWBal2ucljgpyUjve80h6t8aGKFj
jJS46nca0YgBPP+ia+Ckp7A63WTZyhqtmQI995bgRSZ4ve7QRgaU+GMA2WUoQu+x
ySZgyQGqbvn/ZDABjDy7a4BrUCfDU4Iu3goTOfnj9OqGXk0Cfsd8H1uKHqjbgLvS
pMP/BhaGrnDGTnTUOdam48reSHacGI3J1jS3q0swjojDSjzUXRF70CawrwAvx7If
i6exPdfjEdBLxKXaWkhHjbUs1uMurbBhGT2tviSpLXcX3pHVjfVkli8E5wktZ+FW
Rz24EnwfQ6qWaJHq2MKJJcXoYRWpJG3HAZiMO7TViaguy2VsCbjbHADfNOSMUISP
njXWYrkP3DGnsWszP28GNzyuQzz+nQ3kdCalGrw52+U7GHq3uNBW4Tm/CkFd2mMb
pjesAhNlYv29fGt8ZzEiS2ESGvNTJP6GooU63yxgYVLG0ztn6UuOZRjXSVQMRgyZ
sbxJ3J10bImU+ai1ukLHwOunM82sbuZIU5SLBMzN2BMeGVwtshSwXkebgR/8NCsZ
RXsJ8jYTgvvdAT4OvzUOUHGxd3TO+/FqWM88sLOVer42Yfw7zgJlCxQcwZ87VVyP
M9Q6cJxQ7Vv4pOiuxcTwhbe+few+RuczNXWSTAEdPQNJ1k2WnyKRuNc6MvzvZE+x
GSQSRYPBcWn4eemwcGLOICvr9ZXxSgaSWIathUkXDjQF0YHo+kU9eZaw0tMyFtFC
N6LLckORrbRzBP6+MN/iomeFf0UNS5B5T0BQAHPpUDvwUnlVsK0Dcht5QMx3dnPW
AVtlyrp9bCAi2Of6JnEOxuHlzBzmoGYwc5iJ8T/se3h1U0RZOoHRtN6YkfhqsoGV
S2nCdIG+0518FoBY44ACVoKwKzn25WTDsOxO+aignfCiE4VRrBvCl53JESg13517
93T75xnRo+qxBMBnKB9oscNEd4bA/JNtAkCn9tPjyGnHCSO0GTVVT2tEspqvEHUf
izd3TAc+iEjywusAmErk8Av4w6o1NngYT3oMih0zRhSqFMz+GZJ6cDT+4Rr1/AvI
wohcRegJDRUYbWsgiqN7E2RG1RDr5DBfLKMyRkHemji2azN7J2D1eDPM7UZckFSX
Br1AohsNAv+NCKRtDePKyIrIFYsWmGsfQU7UFHlGlRVNj3j2w9xaM3ALFEjtyXkk
CRObz27Krx7mmgaH++X4BPYA+gTMrawDKVelxFkWRY/poL3Z+ESphLce89b8Zvcl
GeH/uscKBqRPsvzs7H8SK3c05uQQlZUOy0h96wtPbY07Vh2xfFGZkNwUnK9llr/J
EMZxQIwYfyRXgfQ8KLRNjrr0V/RloPWwUHXpSoIt1aZEo1EuPW1yeKPmpw7QVpOX
8POcdwmfv+OjyzowcaKhBExV9ohCae+jCvBW/NNOOOYXsl2rIAOkHMPUP13Cxqht
nzkt7rmy0O+4Cnbj+0ATqDR6FzImogpnqqo1h0RKMo4VF1NPCNzJY6QRRsjFodm1
1/1F5ZHHzWHvozvewvzxmt4am1y5lcy0JJzPc0qTuPZwWZGWYnc0gpHLK1iA39K1
qjXN+n/8JXRxirUz6NEfDG1I4xl+KoHYRwsJ/R8C31AXk/UoFUx+PAekAd+VCsIl
mc6qre6asMSFXYR02fpwAdHS3u5WBm/Jr9mHgwdi4ixpuPWT/SCUP8KxW1vTrcXc
zH7KwxdPoOAUuAwFe3v3une6qK9mvQvkwfAVBI1mA2hhpo5byhipynATuwt1voDY
aHmA8PP2mal5xqb/0X9THsg+vZQawVo+4fsUXdr5s2li9HcwlG5Q6dQ1kUnk74fi
2NG/7bpLAICKtDMh5C1BbwR/zzIbydBDH7vj0BNQPvdIGDDD31COZl0nqhvZEW8v
FuCGw01X/5NxQs9dmN3S5CFeebKxhrUrV8zF48+VoZgm6HJ6yhBj7q4LxiidvSwO
kz0wqoUlfWh7dP/Wn8gs+hD5jqubOJCHjCxrCovKDEmMiol0soAMw5W3O26GCTi6
FRqczeYkxgLWFrOdl6wBM3tj4gSr1Cq0KCg3MhMf04QzcpWjllxe3WtIwGzhQx+7
YibkTjMqGirhEn7K7HF5L+SR49S3tQSDow946Megr7lr+OQZsQuuSxgZZ/ULW0/T
BN6nlz+dCA2GlUu1fZkycRrsap6pbCuUpAih7joc3nHYrgRxW8t7aD88tvzTAlXf
KKFnuIj4vi3dBGo36JO+5l4PM9ZFWBp6ZIZ98JWNbyzJIYUbzy7RvKZj98pniP38
`pragma protect end_protected
