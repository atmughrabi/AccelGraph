// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Jwv5FDlZAqGEmT2G93uourMT/YG1LKd6vgGUvlmHH04XPOon/V4kRRUMrTvTeepp
TQ2tWYj+Zk2x33N/9Z5VSdMuN8fszsyN/dxEjjzPEHIAzNkorAs+fXloIaVm9ZZr
N3lisXl4bkMHv2mXVjyIADs2/SqQx2uSU2P4uy0CneE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11328)
L9cim9Kux+2vXlOMptV3SXvPvrRKVGJW8zfxGLokGZ9EbPH15Thv3vG5XQp6e+RZ
X565s+HRrXZGxGNLpHHlvW4HtexP21bOv1jInFNTbLMPK/9ufA+7nPohYyz7iyAm
L/jq5qmZGlMYAJNWldfWPG09ItlTgC/sdGnYKr6cV+IBzOehQvrlolkWsj93C35S
j5PBD6cLQMl6tquS0WwWSNWu6u4Qrg4dQ/+4QGBJQ3Q1zidjdnL/fyjA88rCSYQ4
IGZoxO9etbppT8CSrYyIjJWEtlze0KKmrwuuXkZfH19ij9BAWZol20il8Rhbax5u
lCEQd8UQJDHKCN/rxeqmZYlnp0jV1HtK5EVj4SHZYDTvgIgbOddsfKZdiLnkU39j
jG9iuSroY5YTvVJMWl7a82kKpP90/WTB4hghdIHGkMJoqwKSqPToBfsrkT0/NTtp
uRF3MfMCJyU829ij3iGAF1VWpxTW3lF4X3948hBU86lBgXuty57AwCZcJJvy6bE0
z+WMpIGlSkvAO0k3+Fqn3uN8Ugg/TOylbaqPJb9S7O7fS6waAEXU9I1NtZ8i50zb
hwIBpz1ocowPK36+PjXn07ZLlYf+cDuzU7iaTj2tVIZb62tl96u+YU9pKlmgHbWu
cL9ibTE8R7gpweCJYi3yvUOJ1XzeN+PnJ7zM+k8XLv/L8foo6gfYymaIwp4ZdZTR
Qsac8qlypYOtQTmwthQPR1Y7AsxjBeybrJLFz8RcI9wiyMTZe6JdTOk1EtBtEm0W
n7F6OTbUc8KjDlpN4ccBhjtrWjsKz2aol0YSp4vh3ZwYLk3eKgkPza41eRYtQ6TQ
od45qCnn10rAmdfqoL3uqzx9WLAD4z6ppdpoUMSc8ZqiRNfUOBVMsWy1erDX05M9
9JFirXOyA9HLWxYiP/ryzrRSnvDu3hC1LPx9UgLa/AquWcnHOfI9Qr/pJvFXIYGm
MUARNMwm6QVnQt93pTbkpGrM6OmYQ8VlYDj6C8+oZPpXVOj4TDJnRppSQI7YAcEU
xm7fu7eQsmX62QFNP1eqkQO/XOvKp4xoSQ7MkpfMYrrVjJS8kyvEmfWH+Xh+aUUd
bxyMDi9eKHPDCMjAwJ0iLFe76DKMdhMNDI+XqTYLAiXXrDOEpMCAR3/00or4e+v7
KEqaLDDDqIMRSu9iSdXqkcZpvrmMo8Wak87D1hFyWtOFIFNZ+h+03Q6JkHalAnTR
dtY3dG++C9tSLp4VuyUC4iZ/xrDoKP8llZTtdCeYk5yrdM2iEy7NmATTk7sPlT9v
76HTL104Ps0EV4p0YFmQi6NkwwTKuyU/P9pXBuQaGV4C6qU2LvidFgvwc9vnZVeM
ofFZTwq54jxuIZLPWyqh21yvkGeT17H7bZTeJmzikYlt8t9lPhry95HICo/ocsTE
81sSQAtMQu9MgOa96THa95hcEVzb0bs1euC3Fytq1erFeCgk+y8LOm1hC5f0oJ8Q
+EadZpBcWHT9XyEdhOn8+nLz8V3C3b3Wv3Aw0ruemB0aU53J4eZOSzGwnJVuAB+z
BPVpJT//Gf/xzADD/7YKjUEh5hDIfRnMYjkZoBzEBpAl2uXOoClZftYREe18PCpF
nxIwx/Y5gjLlpKC7fFza/ZFy5IDTHFUGhYktS6uR5KM3mYa6+ANv3+DGt9GvnoN5
HMiupTMUeOE2MoSnoMSuRg++FCYmY5d1CU2jftT4XfKsYSQQrZSrQ7pRdxDg2EsD
xLjUed99vVAGVcBmbqhXUqu9YbfSmAh7E2AQMEp+qVFeCzyJArSYZms0DdvIJmxI
h5sSj22DqouncWT4qjLk8r8ELTY+lk6AUT2WpzT09qq1uQzTRNx73+F4xVq88Ez3
e8UUhf+L/2VCplouhOxNe6oAVLydPhc0JGjqVsGY0olBg3G9sDA3prXxD5yYR9wE
G1KmqVqAKN+wq7AcPt2wD6MmbNBW/TlPF0Jo52fUnoxc+wfPsrKf99Gw2fVLitvX
l2LIgFEn9uPjDeWXVDBNhDMSYA89gLiTI0tqvUj5Rnsv9uTyWJx53YUZeyFhehJn
/8uKAty4otM7JGflsL4O1OaTq3vKIGHAej/kWce61r+jK+Lw9KH8P6v3tuAW0KFS
cWEpoD3QOHzg0WekSqtkfaq902U4o0rENMRpfmCpFa5EcLXmrwQl1DW6VRN7LYiH
UJINzsFi7HLpnGcUXfHBvxix+5jYSbNJtAgWIAazvmB9gA4T8bHuHjW/BMiiQbpk
F8u9EOgtNlumBb12Fn66yV2sFYJOX9ZvlkWVaZrVJs/Qvsuk4N2TR+0Dw9MiDKs1
aSfdnGKFcfnY/ROeT43oORtiIzlscDQHsE5SZIqSqLOIMorRi3luGn8KxHqp6Hty
D8Rd7rb6kc5MVMEx2sMO7fL0nH4vHqkjiCl5aSwmosasUb1hYmXR0nZ7mCGRYWTu
B74ZAqi+tE+f1ioX3nUHt2i0Tz9wZo2Ru8y03wO6eDINFfdeuOAg2zyqxg9oIop3
3Du9mV3Ux/ci8MWD6bDN9U0Fk06A2ZRpeIhPcnnAurJHyHNpr/VeGverijXd9w/C
ODam8pmOg6uqTs7i6l9qq/dPSuwhevjdak2FnBc8lwH/CGtiWbfk0TM1CW8Aqov2
rWe3x6GVpMDotu9u+DYA3udM4yujH1MBMWt303e89Gmpg1LcE/2SKX2w8Q8U24cp
hsOInBasY/MY45AYa+24YM9CiqWC2YevSgUIGWWRfUi604BFa9mmJ/nRs59YdqYU
CD8SS329Mp8FUdc5ht5i5+5DcjsU7+nUw+Nf5VPgimg5o35So4ZvLzwUysmeQlyr
bNbuzoZlB1istCqMRneNHQCvL6VMEz0HKtn4IxZyWWNi+7Ygbpuqm0LPYRBcmax8
k9rdkLMXQiOM+Lcv9UEvAPSvfkIgGz0+Ljrn8XYsTmL8kPHPrsJHOF0HpfzAnZ2d
i4E0vSAxv5K3fwneqrh+lZY+tkwNW5oPd6pVfw/vsLvNrf3jPIn5ccCMH2lp8js7
ZaVQWlsoec3WSDrtEICVtpfui/uG285v2avqFqkacw0/mSE7ISplPtqn2Rziwqci
PxW44I36ONlC4IyrkUHtnNHZ9dlezsTXCa3vMxEkN1NIhh/pLA2/h4tTvBihC1xQ
itrSPoU9drQ6Hi05/lUZ0JLQ1zZHIQwNhwMVHg84nzMZuk6PzWgDfPX4XLSa0kOy
nmaUwVgGL0luPvi8yBBs77HMpY+OdXC6M0C2jvk0cvTD/JqZeA6w5tjzW+C96C8X
v2NkgVOaTiSpkfx8RcYul71SdISj+jZP4jmKUCwQulbPYMr7opORahZ2ReWeJj5l
9japSBL5S5bIp0tILWsYrsae+Tpy+SFTRWtcPGeN/DY00U6owpA/uKavLJBsSth5
AzcuIF0qCwZHdcUjCEwUZPEVR3KnRDnIbyzLzSeDu1aHEYb4Qgo1In194b59isSV
UZjYuuNGN3qgONbE8Vh72H3LgFVCseo46cihOOrFhHacXAvjh5mMzlsHPAP9zFSG
2BxgCeOFvAiA5o8Z14s9TxlA+oeOXe6PVVmyZiw0Hj0dFmPZfm3wqo+3+CuJDGIi
6W72RZoPUIHZTR5DH9meNn3AC1sH5HD01FMYcdIN/1Z38tZEKkghq4DMBoeesldk
qmCcVKNfIz6roo8j+ZCy5xpEyl4IwuOmlZ/8GxtlbY9UrhFIhH6G8T5H+GDwnzeq
2voIMLJNKWg40IIEe094C4gTiyqRhnUw2R//AlYc62BA/x0v9QYCxtSXYtczLKWT
xjMJToMRmLF+Aq4FQKcG/YcJNhS8v1G65/b0cVE/tw+Mz+MFK3keV291e/BcHLvC
uKjZSTDVwWUv4Piwd5dh6xssmgJDM+YALkhRVjnpewX4ReZXM9xGaoMIYYcyCJls
1ZdlOR5yBFZwtxLTJoQzWepxBeVe7z156YwvzZA8fjf2BgcBr84eNbPAaXABbNDZ
Aks8phzGtYd2I2wBVpORDkqmXSUFnyezenqt2b/U3+v/FjO/4Oc9yY+7b2OG+I60
QapXnEGLa9a0lH0CJkBBMHIrB+dlFy4RDLl2zTw5Jl3hAgQPAhfHDnL38nrg1R8s
acCIKuyNlwmedsVS+KM8aShQbqNqiXJ2p8xdNSABFqp1iaWuM8BIN4XNO0rKh5JE
lerZV+EUgoYA4VEz2rvVLbG1oHVeksoEPKADU29U/1jhfKYIh+jIMyO2RXoMZ7PP
6uhn4upnHbx7q+T3YPDYQBsi8GJ+qJEqiyFc7jS00GaraEXWGWnUxcV+BkpF6LVi
L8+5Q6tBO730VbIF9MZSqYjFy6fG6uQu63ZeBO87rbESQ0Fs4abTKAuwFMx9PYwD
MBQ3zkQG47BjWqTBm2EQ/z63xL/ASf4Mf2oRb01PaLnj8clSY9ZwKsBiZw5SY0KC
0MUxBFVuK/2U/wcpIKoD78wRjX8DoK4RsIJtjfnBkkC20X6qma9bf+U8FXpt7PC+
DHF4XU37OWxBR7VgbSo21k0526U7H6aDO3hf9sbfza2ZWAO6AnbWbqNKB0ePI7Yz
iv/EK4ecoXiMGJSONzgeFD5YuTtNykvo0ALKGsbUhFWrBSuS/t52HdGzHg7moEbp
0gxdnEgPqOlgZTj3f/smhK3/Bw5st9GYOILHjPDVsPmjTtvVSpXb1yjv+mhbgNIo
03Y5fxR1Ryi6LArXt+7755b7+x8VQvV6GrobTGV0bUHjsr930JnDPqI6krJRkY7I
R543KE1eCigTUf5FpH1Z/cPnvXRFARShJ01eNojZfbdrkvExFQPPOFMw1FObQdyC
3zh5sZFyb/x+i2hdyfFY4NmVnwt+Y6A9+6t2EBkW1RkyhcbF7lINTLdaHzzlABbZ
GgiFSZCflu4emZj95zOddlbm1BZaWdii8p1XPuv9G1ROlC0uUyzLzOmzsHMc2fKi
uZTxWyD9fqWaXDQrjPRR5HODuEZxoDk2h5G4/XkrqWtrGkcBbTj3oDv94oZAWoTY
8HGi6op9ZIL55MguzCEUS6q8p3aPArs09UYCCzUXl6ZxHPs03pyjbfNcJ9+DBgKy
CZ1MF/8yHTOO5po+hr4wuuBCseUEmVMs5mKLlRSSjIPSqoeoY87FuNV7cXqPe1RW
l41Gffz3+dk6BPgMveMnPv+uQESzwgOHZ0GPKnKmtlPd+3dXme+gtVwSDN9mwhIo
RptkeKiQroG9gyZ7A44/IZWP+Nczmmz/HfbOVjifwiYyUHs5IV+SkK09u7L/aB5P
fwiJ0HzU+1C78kRKQ+GQLU3VznZ4YgRkLMC3/eNh6imv3WLufb8zW+9FQQrQBsgf
+trOZ7oHmqs3c9ayzuToAq6bF0sJg8ARUBrJdsrCKmQh552pIDKWAziUxZrE0Rd0
/cz4KpRQ16TVurKbIm2QYKhtyputCvq5QM7URqRBASUtYbZ0dLlM1qp000WgCZ4U
ypGIwqaS0oYncHYOAph5FGRwzzfMD83m1GCsDstTz1KVbkU+SvjsN7MWIh0Y0OD+
4VSEpBmogCI5qWohCHVBBQlJr5PUgPPSlRFf1IIHkH93tPyI0NTZ8LT9gJJ5l15u
1sGdAt4eea4rnmHu53K7as6pkW8WbyrKSaX8tuGe6ZR1y4OuW72MrE+6hPBfoag+
uVDzeFxlJsP2KNoiulv/5DA9gl+OjhTDvRlnsvoLOQxfSPAYcGVKPdZ5adivOI/d
BlvuVObv2I8jFSVLYxUj+1NpMlbojYp5Tw3hlnM3uYeIgUGItE8H0iapcYEeVV34
7J+UVJfpdhgLl1hOs4K7R1bzbrPoJAUZs7PNmpBWXQBSt0TRLvtZm3K1v2hOIO9D
EjwimMCiv8EpTM99Of4jFmf0UliVCsoCC591kRheya7Azj5gEJzNiihnkSYv7z7c
esGa60UICvAswsheTyAgfidWttWtyHq0SLZxeAGRZdT+8jpjTZowgoRSG19KOjw6
0xyxU65KdzefpATn5rKYqh2TTtA5NqKpekrXXHIg4k4499I6jnQaEZ9JGbSlOqaI
unupL5DslQ7ktvyn7ZUzbRS/lo/Q5hz8rGav3J132UwI1mA4kEh7mmvklGPLV9BT
TFiEeq9HV8Pky10nDozA2nJH0jUlMX50Tf6upmiGkv6gpPHUkDzlXZDdVmLN2YNP
SCXs8WacpkbRjSK2p9frTq+7lMCE+/theT+1r8ldIgdJ8dTqPgqaO05J7B7XLXiK
jfgD4va6jvMeldTMlE1ErSEKRBZBNsqfYcuFyAiEyRTF3wku8SGXvgBuvoX8wKIi
A7u3M3M4IHh+Pt7BnZyyVWhAgXa4ILzpS58SqzqW4zFhx6r05RlO3wWd9AzIdJAd
fQo/LVxlumaa5bccj54USlPwf4L6ZTzRWta8CPwUIdS4wIxpersmHV2h4JdahXFM
T7yfNAI5nhZBnOwdH37ojL3Tg6wDoG3DAOscrg76aD25DlBWBSTmNVIcI7ZtEyN5
AJs6tiiNUtNcOqnPastLoRhRRpbGHl160RUHZmvvwF3mtNY3Gt626AjBxaL+wNaz
MePTzgZLdGP+ZAm8CfX/2INkNmXxAcc4SZSSKp/PtlHqM03xO/uVl8d7j5agbxeb
cvSxwJolhDhMvbcCBMfSRkPEwbx8dG4vWrv1LXDhrOg9lBohl79uQbwfezWrMw+h
CVIrlCyhXCGvgXBbfnceKJxLJCL+tSnQ9GSMswJ3HP+UjjO+WnSqfoSLIA9+WPZq
HOfs4YnhlnTMEMWQ401rcOCCiCb+udgG4iX7abVMYc/LuLYvTJ3NOQoMvzIoLIJF
KREY9iZPEb7MWWg21upsJ5/zhi3zYesN8EpYTc0YySGaELNsAgGhtf9+FqxUe/ME
EuEefsFzTefwsQ2K27cJxsdIX19G/JNhtpySxkZc+sFlDHL++3cistt/adaaSuuS
bGdD/TFBgLusifaWSCnJYW0o4SCOaoBfK+TzAjBaW9qGwMGmGLV9r6nEN1upYin6
j/tXrvrGCWYWpBXLIYlcfGK7T3geH121U4MzItRlzPQv0oGy0UYGhjDb/hJvV6ME
DJVI9bUkf3HhlMZZLAh+UWuxw7oyseMksxGDMrpWvS7yqQMAYzwSzuRw/NLg9I8I
rUKHNbqXwBnf53ORXZyTbIPFixoQvNtF65BUTRttQqdRzRQ945F/TS+2oC6cyS7Z
ctw3kFJXKjFc/L3TZDqcPM+nemZxKA2uH6CJRO7w8w6S3QQuJ+MmKBNzQs92cypQ
vraSKw3dFmBIjX9ExSK/WVPYaxnbHxZXtIv7louHIz2l8eSyktQq43HGlT7N1dRA
CCby0g6oqONFcP3XWO66TWSt5DCl8i4q54bObf8X/V/KpJKhSWRlTqIJ1IFWzCk6
vF59QrvLcw7JfP7Sax5SWNFg51P+cqQd1mQeSUi5ovvT0Al/UR2pHPeCJ9evbZY3
9A69WloJp4EF5cnPB8iesrgfchXqnlpam71KL4aE2Tznm4arjM+jgq5MXFMj3Pl3
0/xutw+AsyfY/1vTwtCmYDsbqq0Ihk1Jse2w/WLdAaUwNtCH14LqrG3e1kxxCHjW
u7Xtm7lmBUiDUyGEfzDscm+TWMvf/Xr65RfmH1gcGBq1NM/4UWnutb5fXx3GS3FI
nyOfs4z464/IC7blzztt9n//mDMLoiPw3i/ywFfOZBZ74rxOUK06MIVr2o5MxtTF
Lc2cfl+YZPLXqkKeCJdTcFSP1M/9dbF+aNUMQxjl+5iAluDk+l4XTk6RgEX3DBDF
8J8BKQH8KamNjAz3YmSQKOaY7JRFzbIhj/YIO9IMnIPRB86Lsf+0VAlTF21iFnU6
qDP8ZisywvXwoeYjaul9lrayoO9yTvSjRTp0OOpI54nddLtTDv79WlOugqQBsPiP
kE3QiMKSocbf5byZsjGvlTxxoFTXma5QzVOoaRIcXyCuR79brulJeSDQwUjbQbSn
HXpgX52+6USTzTs/aT7IQg74mMuvQVvt7ZNXt15h/3iB0O0Cw3cFyeuuGsjvIn+z
vvXib6eiC3Sx1jNVYU31jMwSWSKHTROQLPrU/i7lFOrIwxFkzthZwGPSHbqvPzqa
7el/WN24IP7NrPCReYbmq/2fRMlWFS+spEXSRUBDdv91C2Ctabet23BCeiTvt2MM
veDReLxmVq0jFaHf28NXQCbwNZGGC+SUPO+eApAT6iBFUP3I0O+bNLcWKqKdcTDn
wo7+/5H5udtdpTwl/pimL9DWEFJZQUQweSlyUXjH5Cq0YjvCveEJU56N38A0z7+t
eWVy5i0U/JauMajk87Thf55maPrpZDCBUxKNWwdI63TFzLxqJNfCSQwkWbtUPmN4
6Uejsmj8Tnx+1QCMU4V2Hocxp3NaDI/bBCBKBpG8tp7whvAGLaaXs9orlU0Ac0ne
WLxQ+bwHU4IjzKykua4Wn9v/HfGQVIeV75HJwMv6IJn0Epd0uxCyJClLGANe9Y0b
xvlv5zYfj4jbrQYl4JufLjvn9/WAwfGHggM++O8Qib++zMt4TbOlJl5b4dVkw8Rz
eB+aiQnxw/Wp3zFx0VXri13ItvYG2veeCxzmIJPrLfQ7I7VPqvvWc89rc4kTJ38K
sDLLsUX3N8bZLkt452mmw8C4oJO0BZhjBLHzyKvlWqzm5Ls7PZ8fmg4qcPGnmEWB
UfM/95iD2Xh4/Rqki1fzCHg6dNg53Cfwo+Y5dYikrv/ZRHO4npi2RYHiA1/T8fTj
xOrGQkAkbNVEE0fvzIUaq7ky2yG/kx/Xthcw1ul2xwetaW9xhvKyX1Pm3A3u0W/Q
oXVh3QauPF3rRQNnZ4bWQxmjoVz6lpqWJfpWUPAFj8AUUvhFZgjchCJX3E/BPEj/
2aT7FLtLi/UrGow5Oaspt3rFjl2LOSfoUEAIkWsaCDUBe6XbWWEWKYu3TG0uTM+1
tUAZkPgUbw9lqDYtja1jZ/G86UUhadpHJ+Uh7uiohFvpd5Wk0wTZR0TbcPDArJcU
v/Vb+Vz2m1M0qlMHQ1iGCOq/73srM9FMhUsa0cpt2Nq0mjeq5wmWgQ1ENA0HRC1B
WhrP2Zx7+22xJCv64NvUNET3ynNFHGChRTnptHKlVv9v0lAL1LNgK8tLHERxnxtU
gLMVRI7YudW8DjA8/eIDPjbx8DFKOiX3GEsQwJJQWMT4NxMXWQ8ofBjhCdWgI/lp
g9unjM+IUgKsJeL465Ey2pK4CHQtakSrFX+8MgxQygRTwcSzUwgPkT9kkencEkHt
1G+5YnJVFkdcQJukN4ryynSnT084FABHOcbzKeo2nypY+3OH9Q2tKmtaf/mvjpnC
sWSGEQ+u1JJghuI8tv2OGUQKt7Uk4tvAYIXTOkQNeJil2ohKr3rWZGEGuQjhAM4p
rk+JIb6UKW7WJMHTk4aFmb0YN3czXIq4MSQ+tsh4jGvSUQe1upM+qE3tg4rWfouH
qVmINcpt5ruQPtPN0a7FVVDv+2mLSdOEj6GYFzdpQASZzKCtJg4B6K/IkCVoW7BH
CKXjKxWtElqWEs3iGkoQ/1fShGJ2nC/qo8PGXK8nOFrc2MDm2/e+6q+sTlvCuyTx
mvbxsidTraYdmYhzKkzYQUjj+48HcBSpmNwudmH9X4CZG1CXiDR4lef1lvxNL6QI
1xg7BMSgNUj0U49nKviaSmcNGMTlZjYBNP6ZK25LsUL0rlLNVS0PwtHbe19S0r12
xVoYKEqZeu6o3SGHizE1Zwswjc0g/tRWquNGwwwxQcU/uf3SaA15JZr8j+k6H9RP
pD7oAYkIaiG8vHAXBDjeccwgqkcXWofT6po8n7j3V2mNgnyJu60wymgkDNpJ1+kp
bKr5u1iPUQcwtOXgNjp/Pjg14f4xW/0FXkL21WiGHuEKVo5OQ3oOKj0Z2d+FihPM
vIqzqZU/yoSAR9UzwxF5xouDKFdGUgc8Pl6mwocANP3WgqOoc5TslSZUJeIx5FWK
Ni0dCbLW6zhfyZvs+QTQgabwXkc52Ji6WbeBb8wtONujXlyZcYiepGlzUaArRgPi
yMu3nm+5zxLpKeM1xBFxWL3/KThn6B5ab+2XbVSx2uS0vBAPCNrk4juiX6TZBXJD
bCz0w8qjGkIviODrhSO66Yxai9RyAzB486zap3tvvPEeYOocr/tVdALthhiq75JJ
7QcfLX9+x6cYb+/q3j59kmPNGlVvzCmRuCt/M8mHPlhtgox2P4TTRQkWvJ6OkJbT
1RRhO5HS2DUKQPNBnYxmlU2lD+AyfjEribkDqdU2+AyzQK4RhUwBnrZ+/BSxejDc
dGBB32s85rr0EE61ToiaAWDX1E7ssWt0n05VZ5db2NGbRtkOoYOuEaF+nt+riyVR
cZvV3wNQ9+HV2BbqSy9AbMQU+mbJvBnn+YRLgrd1v70o3+ngcYqAa4FypmHNNym5
NI+ffH5emR4IIVoSIpw3lnnJs7rVLJRtLXbPNGpjANXa1B7U3yIHcBb4NabD3v6v
R6CEEqQhdidsiKZl2ujXlU+VLhbCoiMSHZVH21mcavhf2FeDWHYaHBV1Agj30uwA
h6tSH3TfK6KBtL5EePAJ56KV4iDgkvUXCUefXwmDiT0F3TXTxklD8Vj88fXOuzEz
1W87AWBX2pklShzWWWkEohNNM9PS0C/ipvJJzw6p9fXMk0QAPtaioAgs/4z1WDj/
apd0r/cJHsL6Q8jpDKem5eI5/5SJNMDNzheYyFVSExNgvTGmTG4OnUhjV7EFe4mN
aeGAnFFgBPG+ZUdols1jpT/Yahz0Fb7oJ5h/WF5m33L1nzIVSMjL1NdRrwbzBKLi
ooJbuRlkTNxPlQuSbse8YZdzTijpRQQ+OtJW0Ec4kR6bM7gOlDGJF0rk0tdsf+z2
7JTd+8J1yUjsLFLdTOnz5qErRs1WzIj25RRfJQ9lycWuvnG66ov+C0ikYlSPSDTu
Yioht+nH5o9UE6+ZXUcKI0JxrhHc+3UYN+DbsqN1HhAeNoj6MA2y8YkhMzSlHROO
yITZ6xjK0+JIT59xJa5WMFLcJwGKdo1yEjNnIJ9MLnXnoni9/u21kPE3wVGden1r
LyMQHa7h010DfOC8h8DVYemefJOdzZXuPY6YfBHmXFJ2b4I81zrlIOgE4Wx6bVam
ByhyVThned/rzqC4scrO3L40F1GtuBUCe7EjhYu0xErDIs2W+/PNOIM4DE7rdn8k
xtbi1tue7bihR0D1k5yBf8kSFAwx848p0P9kgWKOM+2tFyvGAMw8ZHQ9aStsvD3f
pVMO39gqGpyrX0w9vKld72WdTw9zQsAdfDwWNjZUvEyDX0cVSNY+4yfqdesawf7E
iMPopNSMAs9ZNbCOZqUWKdpg0Gtyt/MVPwVGchj4k4uPZzV/560EXb1jmkQLGhKo
0jfOZG1Z1S+KKvK/nKzwHhLbKrfFFgVLZ7EvfT3zATak/pw18ZpynMg5BKuixcLu
sjpcgyGZI8ARzmIuPjB+f+ROoqpQooaGZsRuu51aKPERcEYyCTZsI526tgVkAzSE
XUbPJxweEaQZmCrURMFmfXcrUFnWKMc42f/b74jn++epRDBxSq7kvkyt/pzUO9NF
tr4zAvs44beUXGp8GAvi/DXWPgnqgrzvznhk0ZxOkdOycgosWVAkypA83buhTszq
TY8HPX/bDh3fKgSZ8PswBxlPelASVrs7emxO4XxD/qU7y4BG+8EI+hXqYxIOJQBU
Eo/KBmJLMPwl6UMS5cBHR/FyzpBt+Mno84dcEIRgTp59ZLWYv7twQXT1XWYfdA+C
jDZtzZmqkMJ3C3tpZ/gE7g57oQdhLX1U1Ng4DA4wchfqMbuIg4WUuDa8kSNFsEZB
Oh4tzP1qQS/+I1dbccBC5fVRWMFdQZiGIh9+SGsDi4CohUO1VdLqDEMGHCsE4192
3pZayi2gn/o9to0o22f9owq/O65u9KhpRjAgk9h7FDbewD4TwjFBIsCIMXMiXIYv
Xn4QA9pO4RGxGzH5zngTdIeVUWGgKhPXsvytwwPij4VK9Sd2xuZMvlAGIRPyl7rn
PWOZOQ0OfWL//5qfvIxnRrpfvT2Wmv4Lzt0qcADilqucR9iPCDV/livXny3gImvz
qs+pwadTngU+RQZp4IZrIj7PDt+YjZ2vQnpPwOHMU7/LA5DDfcwFBFtxuBZZdvXM
IBC85A5ouvLY+QyJJDW3Hh0wxrFDUP2Ci351B2DLvo1f8h/XIytb5akuEF7QlSM3
bveZO3xD/vHr7Ua+BJ3P0N5XuQUwZtzAzugiHl7ZipoRMQowm3+s9TrIHh3ZJTNr
/qRnzeL4ERZiKXVcyfUmYA/A8QYtvoUrUB5IjXKK99gXMCsv9gHnZo5hIdGMBpIW
+royJQ+LuFqsjo9v2k3RDtpnIUvzuJYDfHuL5KDlX2dQiuaGHSXDdUKRcn+ubrih
pnhmDoX2XmOJp51EZXM7xOXC/l+jIuu56koPX7LmSfKx5isM2QI3N36VnAkS8YT5
FZWwFBqSYTRh5UZnR77ZTRgQwDqWA8DgV7Vk4HexQEPDg/mSoFuX1jmahrq8nsV3
G+TzoApoDGAByckBXTHBBB9x/V7sSsWJeigWQF4W8z8KVnhaDBuOOSMZdnGz43f8
z8eH+SPe3WvaYStZiFlDfHXRh7QTUS5jpt1FnJTQ/RET0zYyldgsRz+nCzlQF09Z
dbf6JiD3fVCFHL5ko7NCJEaQb3jJAMiuQDLE04U3a9vd5szdbUYTDPXOEDXKUGTz
XyaIPXaBiO/z3RC+PuCP02/J9ahpfK3d9LCOoBge76ttTR7rpQw2VT28ybMj5UfE
Fle8m6ZbMbfUCXyUoTSiTwP0aRQlgryMdnFAUIi7W6BAF5F/5TGfdDhA4FTEROK+
HJmEsSlf9cpkWVX1sLBD/1bII3n1DfWEius5tcNIGY0BGUZ8Yz6+ruheCp7KFImk
nE23rh69UXTuU9LBo67pDJw/QOqdW3OzufL5Vrxm+3wrGktUsBPvLc2zS+HOiFoz
lf/J4cgbBPf4SvE1QjEC0RcPwDa290NlT7V8RBD0Bf8GojHj4MnEB9jPRNkB2pz/
3U9CA+NapBHIVJ/1Lnq0BwkgOfvy1x50K545W2ZR2/nd7ofvbjXcxH8jfGgRYQA5
zC58VnJdZ/qF92g7mYPDVYfpdOA5uzVMu45zauUsjzmfVFT9KjMVPY0qgSmg5g2U
0FKfw73BdiHVW+lBgUAjKYQ2mMH2YyVed/GjG8IsbzMidJ6FQ5tpFDBeRuSYXDkk
8tJ5DxfoMUcPhJTG6dVd0XsVenZ3wCS+yaS1Ek5GUF2jYGcpJ0UN5jx1s3G8qZ5I
0oYZTVYIYgcEhouApBdfLQySHnNyXXTbXMQe1nN1HpmL7xqRgzB72HSdywnbKz1k
o4YR9FV0dn96EIJE8srWSupZMAzlcJMrnDflNLojlgTYIXlJQIwpQWfJQNp9KCqJ
+07b5zSWIWtnleD6Ond7X4vCYw+eSTnDgT3viaDtDExwHR8krBGlHTlcbqxiG/91
6syGEbbaMp2FwmAXY91EXtwkUNgnU/Pdq2QZ9J65rLpKxDUvzPiKPSavkIlJvkLi
QUGRaN0D9Oiesq8mmQL7cTuEi1PYa4LnmD+erVzpxmpdBQQHBKADNLDe+CpANFm5
MZAfkp/lDpEZaxSsfup7vTxQVFjRqAk2rQuIO9EkMqXjVMzh+nEiq4hd0bpHgwW/
1KbCg8R60A5ohz50etAnxoLK14f+ENXjOr1drVsWmHkUTa8lQSgl2JlGBXcRiW6o
diRLheWJSMlp4MyjHoaCci34uPplmiklbRuujJCFsPM0+pG+/txgSqFf7ZaGQX10
14f/JQY/axsQ0c6mhl9xumwZXub2mIlIjODfO2PL/027VX0i+b0olzKiLlE8li9m
GZsrEeCcezhyq30PBympN8c7P4aLXXlXYwGxd2cTVbTo1ORdyYBQ9ix2FcZ7Nf5q
luGPrbKhj/8ub9OhA0MCiBXmZ/GdokYN83Q03EoOcUP014adFyQ7UhBNZLNMhn4X
T9F7G9Im5ACZEmL+ss0veuVsX0V/5yoQRLmOVOW0vIC1saTkuBLJ0RDAaJCwPRxS
C+ErEnReTFFFUDnLjfPp0bH8U4Up09S30MXlDcZFcn6C7JGDmfGwaZsUOGOnNAZJ
imJZK3ihgI+aZjd9XNJezV7nBpwOXo7llaZDSMtHHwj9TUu1LgHYtkqPRQa5aIRJ
F+ev4H89VLGeOPaoAGorHVEJfaV3vgkgFtzjvpSm5Y52wQbCj0WOfVPpRPDHBv8S
BsdSvvcRUNbAdODl1ZWoigvr6hyN2TnDjeYWAP/P5VDX+qE0v5698N2MnxlrMuRn
/3cRgbt0cWhZCQaTeDlNuY1E93aUj1frHAjDTSTRNsOdwjgsG1u4ITM/J8TlIo77
QfihDhyoy5S448Fw0ez+EMX5e5IVoNj6KqOp7hWTxM2f6vJoV3wfiae9naROp7+f
zZ/Lh8WlOZTs3O5ihBLrWaxWVOnVT99+XCDTHrgEaUbyCdqNSzFuizW609ZjG/rn
D2WQRDr3AumY3GDWojgBavFjqS9eTO4wix2fZ0nmswI7hkM5/e1PnJN3oT+xx/Yj
kuwxSx6cUdsVnZjjn6LbATL97JsUFN2U8yeicnRga/QvSkWbrRgbRi2WUW5O9VFH
H22JnkTdJjEKoza3QwipBJNbD8RuHvccbdooSGNreAKpne/Un8kXNW1TEy6e6hwd
PdCLrsdK4MS2HjzjMGsHaZtln8G4W1sLZIIeYZ6KI5ONeotOoml4063CCv+00X9F
5/OGkhzmgiz3eH7edyq/1rYrMdF8c5y0CocuQwLIMek3ea4nZxTDMVwVJkYSQxFs
8u4k+tfHm8CoHqnRUKIb6TFiVcR+XLbcbJxW7qCgxxkbA3i0pJiewoAOqltqvCVL
lQuFV8E6i2CQGHcJmp4yfQgJ9WtcjHgEThrKtetTjjMoLXLU6WF7ViJQaYP4S0rx
QtpJpdF9dr0fj9UaK/BhFOfKpN1IfhGnOxe7XtMUPYKYtgUlttFPQ4hdZ/3PSLE6
BkrtxL5m+B9MniR1E/r1IUeMZnec8+PBY889afo7XasEp6338/xV/yMrnZRxVXf5
ilqqZ1b+XF+VPmhRAEaJ2A2G/yJJLvlx/ipt2GIwa97+UMtWZLQ79j4AHfPdsOqv
`pragma protect end_protected
