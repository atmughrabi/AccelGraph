��/  @9�n�4�gߝrk/?\'���b(����%%�0{��~�� �����ѢYɡ�q$�N������َ�qI_�K.�l������B���@G��H��6�41M -���3���y_�b�C5<Ol�TW0��et���+����HQgV��EnZ����E���Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9�㑴�7e����P�K8�Ʒ���inB��ؓ#)}����g0��S30$ꨔ�m=�:�&&p@>�ۼ��p���38DiV���,�_�,���Q���O�/��R��Af���K�Yp[�ƥu��������a�G�����j�GF.5G�whR�q�u����o�v�]?�➘�>1a�h�G�"MS~C�m2\��5�7��r
�\�+�^(k�Q��gS�������F��XR������t�wR�kd�'��?ق`l%�=,�y[E� �ܪP��C������a�K�D�
������~���|�̋�}$���� ���V(���J�Cp�:[�O���
�J���Q�6��>����}���K���
F���u������;�m�����K��ɯ� މi�P@�&���!�k���eS�{�@'z.�����h�"��-)_�8���c���G��ҡ��?��;����i��GY�#Ϯ���[o�7Tt�/�[���v�o�^r[��\x�g\��f+��#���#�C����1{�c.�L���9)ĜY؃
%���e����-�z�؁!�C��5?{����J�%�=`L�r��d���<	hR#q�AY}�#���Q�3и,*�RM�g�Sx��/�4a]�|6:�ZC-",���l�#4����V�$����nVvO����
~���^bb��;��_ ����O����'�Ί䧤~1(E��,6�|`�*N��y�{����e��e����0�1�LV�F�~AD>��W�{ܫKe��U�Hs�5����|�	��r;yK����U��^�h
%'9�%�&PX���f��ב��/�1�,dw�]�JηQ�7��,2s!�����J|Wh�t��%=(�]70�m��?(�>��� �]�������n������ر���-:^�ݯ�˃Jt��Ԣg7�6!������[��7Z��'z�,>^������d��6���J� ����8:(Z�(�qtaFb#�g��I`�~�R��Uz�0
���.�z��ƾx�ⶼނ)��5ō