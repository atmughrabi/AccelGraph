// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OSpV6zmuEkV7U6p423PshzWjrM7Rhjb2KBWYmxRQLqAHu7f8SRKED5os2XiiiD4f
R3MjvP7BxBn99KBTR6eCW83MVFxdgWM5eSn0woQcOgysS/nC+6Kh3IJ09RuFjI67
xnZmvisNsrW72VJ8RZFC2b7omFC0Sjt5e3zjwnaPGg8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28192)
Fd33t5BfulcRcc5EGxN2kcJcQcsRAMriu6EkNx3mQQEKWGU09tl8Baeog5YHbJxs
vp4ANtCjLx68HZYUvMZqxknHjgoNng4xXFBbrCCv4aZ5y4oCJTVuaDTzXXLPwRxN
laCcpU3jiXpBTCeXicilJJAr0RfijT8PRtYTeXmngMi4cLClvh7bCDC+bgAOPfUz
2m+9UwXays9I855NqEDep5pNqPzCD1VD9e49Okw2DjhxnDLgoMtTKIBRyU3YtUQd
mLsRD4YL4vIfVSpTaMJpUqAzj/d9+yhMSz8zVQc2I013W+kcXXMd4UbQUYVIhZUJ
epZ62gt7DUcNgI6EcvYIH5MZCrSXt1b7e4sL3TdkObJbTRDYsucpGdPeSZuPQXzv
G0oHSkaBEYyJdcPVvETwlO9vF1sE5nt9GZkci7QMXiDo0ra1UvWPrEKZzky5SJLe
q7GQtAC9pPw+9TR7mHd1k+qRS2YaoOlqwdQ90+17j18QAzyT6CO2jqK3Y+xZdVK9
73LTNLUDoWHwXXjK4015IJABA1eQDlOWytL3RBRrm+TchIgt7cN6FRfIb2f/2qYL
whnVaZNMrk3hUfPim3kCyzaI2b5TetrUArg5td35snvW07XeKYPTi4h1zQCCZ7R8
oldilwRKkmArB/QmUDAUYMSK2F3Ih3VkNw8S6msPiMxSPR3UO4zcgecmtt8KGeGR
gZI062I3XYd1T1cidaOV+zbVal8kHMdhhLr7xhLtDD+w+eC76hIep37FygCdmBtH
GSQsxt3393uEAAV12TvYzix7tKB/RVwN8a+oNJt9FGpQvb1ZvGomVyZQbEIdAmFt
cec4FdewELMXDYYBNVh7ArVFb6+5QlSOnlkKKEG+wmRXCewnqfIb9pK+vPEHaWXN
xFSTvldo5+GGUIs2094nB9bWzO3yizJ5kZLBqWziURtkkcRzo1lGc/OvnGbjlf11
a2Dwp6ii3mOouZDvBNQWdUe9UJv/a3F5Dna7HeBGQumEmilsHkuPCHbhl8b9Hgj0
TZMCtaB6jCtlbtLMQXvRbGuwVDrrGQyp7sLwAdhBvXKoS5UHu+HW6onEgPS+oZ0C
+alsnO3jodN2ad6jrAAXFTISFzwlOdfHTGvbnZGwjzH2K6S3GaxbCA1WfYi5ysX3
GentlWtEOuMbYmrQWFKWnm45sc6jw/BVUkKyyEaA4KN/VqWFv2ZvPh1UrTGStoaB
+ewwr9ohB62zkNlrUZb549Q4JOOv8o6sOdFG+ZaVOe9OoCp7XCY1AW3/tnLYVX1p
adEbdaN0vCiYakCs9P8gskuFPUP2UT18ZFD2V2uBag23/xAwJhNd8dxXYaBzSKaJ
VSXDcY9WTAg1P2anmTsHVUJFkJbIJCJnbGTqcI8SdTKss0Ww8ASHVWSC1cd3n0sb
2F1HNERCfAiOQHqET1aE9w5YJdtXk01y19kYw0bDzYeYpPkMNnRyrtBMWz3I0T4L
LlGhyCVJOTMOgYlxX7WSAlLEPYJ/pS99P3uWGKIXKn+o1RG2j4oiz5F7MJdVT1Ma
L1Wcx2TSnAQ3Uwq83sl0mRos0MNeIgUohh7BrQ2j1bMvgYuLGm57l0zXD+El5Qsv
9sNM7VlbIh0CDynOYWFMul7Er3PbRYaQIl2fs7b87ULtArB5pZN1IxtrzOhw1GpR
80xqp8V2QPTFLDc7vy8RaxJKsESdEF+dyO6KrZR6jSMmzm80dmj2AxQqZm1+XwNT
rh9L2vOMIToyBoBrHYyv9NR81OVA5Dk5mFs0plK7CRUvqDcOiilHaix0Dy/PGrF1
Jm0QIj+xp2yVclAOFX+H5n/vG8FoXJBNdvfZHXOKbIkmUUFmgCT+y9OnqYfVCNSd
J7DXoGGHpUJWmqa+InyoUXrWNXo+bz9TvNOgL0I3d4kaZ27691vYqsVRdcwh3eL4
2IyBMMi4fc++sPbO8i74F2TaIzyhjLIXdcxa+neoPvGm3sFmXm9smYqgJOYkDg15
2pLe3Wyp50SaiCGt1nve6meuzURhg8PMcxf7VIQPxZHNfLZovjHsjX4N0qLJBH6U
GY6q5LRnHpTR11G67eEAPLgzCl0xyZHfD9x5m477fSmV8XUDfr2EVuPfAr5h/EWg
9XgLHVWdk5Jwv2LmFBdO+Yc+UVhdZf7KRrOA/JZKrXPveP4r5Qhv2Df/T5zMifsr
2kvzq/zdj+CI7/lz0DovMjeHlyTIG0Kp0+ndJvP/nbB8AoIxWR+rtis9FCg4msRQ
s1xMXcwoRMSY/ExWR9lV9tHEO13iPuugGH3hdfBEsyDyiqMtcRstAYoZdMfU9grp
f8cnAYKgIXYHu0UeuVrglXMmCDjS9IOvLX6ROzW6OVGM5AyFRxaKTwFlpa5DfJWY
tBfteJdlwzg9lWdVBZsHc9w/C9+rSv9FonXW2/QGiLyBRFOgEGixONQDZdIMckPw
08swouC4ObDHRq3E0XYW0qAGBLH877x23ObPBnugoBteyyDZRuy2FqABiAPsS74V
anWtjI8xoWIf25ZgT7mov6bsU6tuN4+OwzubiQQMj2rtIDjLdzwY/jZWhvZTCSa9
XLDB91syvYFHLGEIW2s+q7v6RhhPjSbxXNq+vwjJh6x3HnvrrS6Ek1CU26d6p9Yf
ZXRICZpyA7E0XHK1ctNaheE3Yhm2FHuoDhLK+d2xt2QYYGNM2K7Kjj11N3bEC9Nd
OrPVSYbBVp2SvQqX4mt8lDTOD59fC3boLExq5waivjEN3X6EWFk4Y0MUFWL/BsbO
pw5+pguF9SFP+fBgBl639vWiT6O+B9u+CT2K4JY2nFvjEx3bnc75yElSN3Q1AoK8
D+L6/VW6wMUQCXfK5aojnt42GsZm9D40jPr8vhGvdUke6PmWxsnoXwbKWK3vaekS
VAJIMInQ3RpMYbUNF1FxnAA21B6GrRr78h6/lpdWs2n4ExTu6cindA4GGN7rHKbE
8yyolcBBzQZoB2CB+scGVwLMYtZYio07j8Hd/67luwwfjP65babfGftnru6shz+D
xYXhZwq1QU48SWjNZqv9RCN7qXT1wyHxmaAOyFissXnwGgXbRUcoOOqGXhW6oUJB
c3tdXT0MvNOGRXOri6m40oubXKB1GYdkAVEHJ7aS1wuJBReHjtLp8CdkyuU+zW0S
j1vxoiWMgBJOW/CrcqL5qGEBN6khxy2hOGRphIAEsLIoNXqXQqaICCIU6tqOh4lE
B0DQxyl6mRFdhzf+cG5k3qlxsL1oPe6fBObO6Ca2Fl2A54Ax+0HcACJE9gjmgjpL
8PlGDdY0ZgrpUExE78DOvk8+IZeMFS115IaRi7VpV3C7311aJBHVkejD8W5OgB7P
i17d+7aij9r+wTXJ3aK9TJeJSFV4a/F1QpO3dDyU2X3qhjv8dJ53OcbXww6+RGlj
poussEPzmbcvGeYSpT/UCDvkfv1mJgES1QTPjVnTGvB5V4w+8czSd1AoXxQZROYT
OV2DhHFRcOI4Z8SUHK6VMjspssMHsaJq2IxoV9yWtLhNeqJ8iHvto2MYUrDXCcTn
Y74LecyO/XyAYEo+P1wEkBe2u60Cu0DC6a1IkfuhKEaCcmlD7Co69li2QDEWkvke
Bsa2LpTaIYCliTUKH/SXgSKOqdgt5Z4q6LoLlltTiXO5027PoxDKBm3cLw6UtM6B
guTE6guLWimcBW9TDaFPtOY4WVo9L5wO7QvUWd4T6ZCdEZAPR1t7oatgpreQtzyS
nNLWFptdGSVkYmi6sjCmduRmBpqZ5g3EQkKhqOZ844daTj6Vt+KPuH4ZtiqrvyTD
ngz+7RgAM7ijXs7IhexZ6ND6qdAUjhzS2Z1bJc7N4IMzjXn1saVRhwKWSa8SvfvA
/GZSdNr4RWVeY1cV1kR9L/grLEoBNoZOBcvQwZyAT2TJyD4h2GzcOtU1uRLx3fvG
ZG9n4upGtmx15ksGkza3YkctvO8x2fg3NGbvUDd8Crv1grpzJUb0V6q3PTOzZIt2
cEyPvFVhwxPDFP4i0cIL/h2zCh4xdEDfLa7abu3CVLkTZo8lwtQUcKjkK+qfULDd
tdfKN1IMydFV8XcJFyz6LxVImHWBDYh7jIVuMJDsjHaFYCP5MfkjblYxuHFz2bG5
hdgmxCZMs6VY9ixfprVgUj+FE0anQobT/S9AjrWzAdafK6vI3fO9a57Bjsy8vWj4
C0TIkpPkkUFP9qoJW8vBRj+zuVRe7bTyerOCXuqM6CpXejO4e4tFf3yzrz5K6jtg
yfTHPHobvarsjrvCtW+gpc2ehdaEe89snxeqmSVIK+taC/ICU/hiaXct+pXc5mkn
15JLRJYn6hFtmfPlqdH53fz9OPsvf/MXqc9fW3Lmjdk5ptjWk19zM1CE/PlPOu0J
dAk847ol/KYf1fN/MD9OEcaTchTylmGj6MocwodLoL279uclX6Ay+X+nPyE06l+P
q5kOGxYmDfiSQb8XgxGCGzvKZoRBCNskGQhVkE+Bmcep02Rg7RYQkOKjsM4RnzWF
ogGDq2m07Vi9AGRWXEJujYmRexMeSAEJ9LR4nT+Fccl5jVu4o9ZPSRYlAqkDzLs1
gaIPyX05xw5Z9p0sCsUVUisCJYU5Paf03alyPfPNXNbSqUCa/NjPE2lBjT3rc5de
XnrOOBXKL8y84QLJ016aJHLWW0N78Hv5xuiBCzjW7yN4wyALoRKbXQqMgXGumjto
EzGrz2dCqf/tV9NlRueRsxrasZfd4EngdZ55hTtsLVZpdFjyaIAQF77SgDjXsRIM
L5LHU/mKzDcm5EfIL/bNAsEVEo5j0dYAETssnZLr89tC8zGVPHSAKKumeHC85S3N
HDkq5yE634m4ztSBGt5PDoRijfM4sQ0yZACnAjEyY0BwU5ButWjWxeYpyCGztkU4
GpZlu9qpN6NZPQItEIivl1nRyIlUwfzTRh2242TEYWz4zsovfJK6igywYhOTp8J7
NTf/zZlMEfD4pyWIXMPZI8EAf+X31jNHHsswJ1fszpQVcdymiiDEpof5Pu1alEew
KbDKDJiZge321GvI3I80L/bBdbaKNn3KzQU3075A7iJFGLQ99v9g6eqEKFrw8upF
r6APTObRkAK82UsSv/eNPQc5dMrxRYoF70TwAVfHvxLZF473Qdcj9wLFFZvTNz6U
Wd/WRGMFpYEPgeposL+NCo7a8zaAAnvjcRX/cvkSiJcp59yUsFt6Si9lwAxTjMTY
6c41yOtosGNmIIjAaV8+xeaPlOSKuCxjAnpPnEgg7clew0xVFpoZ5dS4RtGMKnUC
npXy86CVzdemuop5Q7B8uusjaZt+JUeeKijzd2adkQPp9SMsaK58+nRVavLVEuIX
q79iUukPaA+44+nGrxFdEHUNQlvFgANBlQHGLjaab9mZwQCHoWabu+QvW6ieSXdM
fL9j0ZAGjVx/u0YMk4VvnHfgiqpXpmPiq3KHSDI2nL7ld9rq1FKxWYvvrnRa8R3S
Jngj2rNfFgiqku0CqVV5zfZIfyTPiQc5wHVVkyKALHtQEhzDS8OoLZYNvodNzbzl
RBBKSTzGShLvIa9JkJEKAOMiXiKNpMgNrBUYDdslNqHcLZLOqLyabGnoQ/HF+USU
nT9wFSrBmfUxIeNmPNj9J8mFMnCLFePHrMQ5CNMiLIcVGWAoemeJKHaZ4J5p6dGQ
halJRM7VsDARi8phvFOXGciSyLngNeiM6Up2ySOb5ZZIWdEUZJlDTqxvWeRQaUl6
EynwP6ncUMlMshU1nBSilkLmpP04MRpzifo3oQm7X8Q8Ktku9WtcVv2HSPaqOmZ4
7jUh+VCJ+mcokYvUP7Bitb15Pton1ZAsvnJIJesEKbRsgeYp57v+zE7UJX1df0NI
oEughlF7wXTIZ/peInOsFBL96eccz4yDd/I0GZ1OONCbsCPcgewaVN/CBma17esl
yLiGnEnjR/byNc0TPpZMS94KKKXH7OdciNE6buG+f6n432xB2vNIsblmDzfQ90cr
H43wsxd+SB7XR8wxS/mv8j2OqrX7GhJrLfV50aiKDmMdT43OeWoVH5H9Ztwgbaky
eGbH1srgjEdbJdSnf5oLnsMKmC/JcVs5qwYKnaUkmYCyuX/sNy+HnomsqGhBxji0
w2rPn99dT1h/e7AB7OhE7X8Ent9dW7dOaBUXqEu51c4Sw4WwsDAuTdjDV7Vb+lcc
VoFbpVjXOAK/Wqwg4hDPXOfzFvR9fFhIK4j8eSZHVzjbzSCJ/oVn1PcCqUoYpi6o
5pKeeabrW2Csp26Tvxsft75vcSFAPBh2ZUjeYKvBkKojlFDcwy6B+tm+COO15mLA
KQE/m5WJGI+fk4vqwagldvLflBQhGBCSyVJLcuRmaUlaArXgUKFH9YcqWbIR8nsH
Hvvvxc9gzPEchUGBlJQHvBBb5hacCtDLg5yuP8VFoQtF/sOIFjZ8X4CnbuieN81J
Qtz27B63GXdGdIOVhT7u0Q+t1wA7v4tHiICNeSBAT8jq0xD3DsnYXRExCLMuo+ex
rb5V6hGjjBmXMlqQz7xQT5GNgKkPru8pB0VykA6/C6adEnTmgQjSBXBV2265/DCi
4h0AxH6yoD+XjzFDUHGwI7YQ7LyqWyveJ+fuKsCQNp30SBIUKIcIZt/STy2SkMmq
c/H3YQeU0mUFW4GlCUPTbtEPc3pM/XhQl8eDD+yOK+6qLkom0y3eQmMC4zXUZboQ
xRg4MBZ8FR542cuGDQRWwV+xY6GE2b3tXgO0wf9zYIE5kb4QtwFeCrPzUUIMy7QD
BeICitqKkmJzjbfb45717xgLare1esyZYF4n3Vv8Ows9LhctmtMTmVo8KShZKxFd
S1Y4sPqhc74ZkBFTP/XXQxtUj2uPPwl6raUxQw2yt4y4cuCuLaXor7rlqoHlYCZq
i3rKlAALiuJGkHeMYCqaqoxNyYYaSVMyttD5TeuFL5v/I1JrCuWIxNaZi1c/tfWo
wPOFDmsp35LFi4BH0/x417l+kQEDZT5uPEvj2Lrtaobsqs86GdksUoT3F2aHqGSd
5QIlPAei+w6MX3sOWh2hRGjk+DnJo7zKmlnLVBoIQ6vPt0syWwtLJEHA61ELiJmD
s9pzEWxyEn+g1+QbXiJk3vP91QZIFEsCmXiAtvp5y7Fg46RTLUy/Lo5z2QEDfYeD
ozzJysHd7C06ULP2sqLDEcoT4aiPdIgfhC9jb/VDvR3o6EBKzg9qG2tygAkOI6fW
VxCV26xLbQR28ks0PmsM09eUyFlpNzf4aVr3g+V41BSFJz0VeNV66S2l5ZtLXh1k
HTuDIdJLjZn/4UohkOK6JHM5vjlMwq1fwpsIJeC75NsTap3wuHFxZDCH/eNI8Zef
Tdoi3/0LmnV6Al0xmqu2Yt7YRmKofydXujdkxbgJAgJ+jYdu8K7sOpsbLYGqP801
zTMfizk0yxKpmLX6ObyKsQPJHUHOaoLRKqWgItt2MtU8XbautiHqpPpclUYSqKzK
MVukN99WE2ZlpeTusi/E0H0Q/g51rIAot7UZ9RDyjb7G6p2rOxBbngeEUABYxMAD
g1d/GX8P8hANl0hTTkUfF6djRVvppL9H9/etzSZ8JwMGL7pRteyKdHrkCBpznigR
Pr4PhGFm9OnYLY985aJ7Fb/5tEv5XMIzfXjLO5rvId1nsTeGPdy9DMMEgJj26eX7
yAFV0HJjZVn++rKsWoD2oI1Aw9tW5tmMM4SazwszsDcaacvis6rKonOVISdtKMo8
Fkng7kdglTIav4pdJcJrCi6eSwQE9JtBnvEL8Jukl0BCG5jQupHMRcd9rQPr5cSO
LuBUDdUpO56h4ciOOa/jAOTR/LoY3Rcfn1REkPcw+dOySRSa6R9CsqtxETvsTwVW
/NnhWZneEikf2KaFPdmDAq8lsYBb+NDZWsL5z8CzAoywjz1eUct7CkiucOte2V/9
W31JodiOIPo9ENF7zRKIl7MJDF5Xh5yr9sQ/Yd1+7OVyy9QWA2fi0ct3XybgXAH9
55oGfOvrbwoyZSz63Vsuk6vvP9Ejci6EgwvPo4+SsrJMDhVNjdFRcYHBw+UWj3ml
hPtqbKaJwxlxJUeUJlN8WZkvby9yRCi6sfjligkGGjElhkJdeLt9dieGDPhgnip6
iLlADaLlLw0NCyARz2NSJI4vemgV942USixlIvppoeP2SBai/WaMUa4PjTH4P8Ex
Uz8ZnIPLdEEyVmzIH2jNlqomaJZVPmFuImi5bX7jaXuVeIKKPYTW/+TV3bJkm/eN
q7V1ycTqRMPZcthMeKpt+Yck7DgmU9heIqRxu6KIJ9Au9Y4QgAlurDBEtpEB6lV1
Iakc214Yuah0Jx9+k0tg8CiFBSFZSea9L3TkxQMPUUZIUK0D+beqL9kv1P/L5rgr
I3lGPdVfRu3kvV9nYq8SV3PfdkAtNHLp1gGh5pGpX7Xlp8WHAHNZGGVvQVOcRS3a
lyuQbsTffNtzDtkZ2uKk2ybuCkr3eurmIPnloznjp1vMhI1wx17RPdUhHtutFhGV
xFGkMyF3GJjyc618Jj1IybibUQ0IXPaVV1P8dYuz++1IIlLqvlpriha1li4Bj/B0
Amd2yJ5iTPMByUBMDHTJlN/l9N73Sr7hR0M7kUX8ptwiLLeSrKk2FIdmGA+CwLGH
5WT9eH6+Tb+B8K1E7r9AmL0PZe/qIVPXzTcRKH43FgKX94TfvrAwa7yZoU/3b2hy
vsOZpPqyUuvmPD152D3z32scqxqGTcKCQIR1mPdK2bnrKaBHg2sD8TQJu5/2MbO2
CTuM4bmXaHZfJAvtjQIXrRK/8Ii8M8v/PGDRWGhgK+34SMUt3nUCc+xL1tWr7cvU
ZM3fklaTHGgbr2N5ZQgk0vx7zGN4qphIGdN7zGLJqsFyqAJaPaT+MV/iunaUkFhJ
reZeCeyyFsrkekxdgXqFSvj3dosV2zuTeLVdAW61ikIUTqyHMuYEmlYMQx3LAgGo
j69/kFpdaYTK9YNBKjUNqj6XfUDhdVftws1H2e7g86EbjpliTwDPNswsn7seVB/G
mcuUYz5c/2pWzvYqcKLhCgTuztIpbV4DmNAZ/A87jJiY4sCgSL8ifidrTkrbWmxi
se7iXP/AVITV5kNT6/n1jU/IV+L2jbA4FK4JF+dU+BZhJ/mIcJi1xPCwUtvpd8dm
YPo7FFhbqo/CNem06tBnLa81XMx8k3iLOpzo+7GIZZjW85uh8Pt/BCzM37HM/kgM
NpxotdINqml1iNtkisYcSqJT6f1zl8yabTIyP4YKZEMYhiZQkqCcBWu38D4ovV/0
q+Gobrn5nig7T2WRufKOwX0uRC954zh8kzo+y16iPIVyQiVenhJGpQFPbBSBiZ78
UOBvfQv7hocfj1YbhRyXq48FWqu2yhWnZoactX4ReU1EHUYOrK/squ95UrqXyLqs
bJ5Kr1A9a8T4I0WdxV5GEPlLkvA9e81kxwOFpEq6Bjvqt4gGSjtiMtUnxkaMHpSv
dFcNOcM2jgiq2jHTcW3XlfaUFVwRofHIS5kbLzO9ZSK2uqARsNt8mw7e5rh4PpnN
lDUdYjrqan05OzGwYbYQ5G0+qYZCEQSzSBjmDwA70IETYaWw1BQ63KseVFCIB1/O
1bdXYhn4I99REGq16hoC9ctp224PMId3iTkZbD7WRmr7U/qDoI6z0H1KYtHhiA3b
sXsVXGTovb7S//NV+UHx1OVO54AZ5A5YodOb3I2dS3/xS5wcavrvrqPzNQs0E4+G
l/nOqEPIa82fJHsgVaxIZ6ThA5yM2KAYg0dJX1zy+8jMe43Whmrt9UwYHlKdkarN
Be9HbzpQSPedrSRiPYIQzM+NNsf03FA/K6eZUZ6Rlo7EEkjQAg5K90PUSL7oNx2B
rM8huckaJ11wm0A39P4yp9+D1FIci9d4xSuSv3BMUH0/2z2sS/BD2DKJO3cIH+iy
sjHbbKlY9zUzjXslWTZkWW6wJCOIEaL7KDVkr9VhB0rw2jo7O6Kv/1VS3SCxtSfT
zIe3/lPzIGwgUA70fRb/5gsFuPF4FMCMKHu9zEOQLnlOVRzryCu+nZW4iUIAU4K+
Rtt9adpR0biIzl0sRvgp8Sry4Tf2iIWYzu8KkFHqPHQvO/StQa4KUjbsq0KMW07x
m+99eNP/w2s52hiKIVW4vDWQDPk/PFyI/lnRRp2fsGCpjk1kGX04QZgMYBmzhIKs
nFQg/mfGYEWqw2bwtR3ebxG45SvuPoU3MRoMZaA5sNhSiZ95rOqhMyyElc7Tf9LH
Disz0+i/H88pHhkkQz7rc7EyP2PgTSPdVii6PxnHSrz/VckFOUfBU5jG+D0AJlv6
W5Z4+zTqv59w+YFayXIRRwPm3EimRrXwrAGmGYzRFvMEkibpKFMQqYK4VDx/gGDO
Hv2/2VpPfUFkfQCEtlVxY4Bl9urxk2DQzJbvwLIELKDKzhN+DA+VLJw+tzBmP6Pf
Z6VinfFrtxiJO643OuIZrtYnGSqckmiZcnL+uhB1mJYIaKCWHuT/MGhfLYpCnJD5
UBvDsTGKKEF/vGotGKzOKl0RSH3YrmXCXOrxQlGizAAD45r/8e1zWVylTWU6VPnL
SRYr+gC7M250JfNRSQk0uAhCBYE+qz+AclXtPXCg/lzezXDb+Q+FzYcdbv18l387
ZNYClLDGoCf+XAyqo08EeQelo+OU4pIIhPTtNHkLLRd8nX7X4iu8ICa3W0F/LRGY
E/xoC4A9OmDcnXhGDBqVlivcMWWxZnO3yKOg/B79z59MmnPI0tn+5giJz45k/TiN
9OaS4CJqeO6gkS+WfExkD/2E6T7yLlyf/lpc8GAJp7XRcF72kUv+7RtRebPinTve
A8DKmP31Fa7QNP/BSW1uzDwvtScQ0TmaUa3f5QqeJyIBRSy0OGubgebyzFdGEWFx
Vc8LFsmHAN/TyEGLyV+K71+nIsK03ZxExzPf+fkFVoiDAGUiyPPptkmY878Gc72C
4jl02xn9lkdEuDus18z2OFXyy9HXJlSEwSXGEm+glmfuJjHDwWXYxMiPCRcx9PeA
TfVPjvQdUQ+16U0FMYZcfP6L9DvT8kibJ2Vsye2kSiiqm2g1lMHj6ahSR9yfYSKC
LuLfTefcBE71HE6PmLZa0LrPtK+jDxcHnrwOZ7pMhKAeAUcvSLx+d/XoYh/gmQ/e
CnaaTfs2rqTV/x5J1TjXbNSKSdaHLsKqBftCm1xWbbyhLhEC+u46TzayAGvkcSZZ
xJaMqPaZIu+3K/Z/1XAaIIx42F03zxx79IzyqZTR98pRETrkmWhnEvFLnAWQIIrG
iwJ0qtkOlnQ6mmn/nQ3lE0U/3Le/4Xt3e3mWojrKduWzpq5LV67P2u+lk+sW17/A
PJWAmYJNOBTAm/0t2p1Q0xbjCZjvk0/1WLTbgfDScStMsgN8JI/7n2YYhUu2x8r/
IeBedDmUpnHP9oeKXtoonFg94dyXKzBcgmONQaonWJz3uN0kmAQpmOdWaGX2ncu2
iaxYNRbK8k+UgIQ70xpS2MSh7f6lJ2f+8JJP6Y9kAKiLkF1HtY1b7Pucy09ASjzb
YswrbTtBmAFHe8vzw2N/gnc0eaSi9wU+0IcB098iaduLoCruT+rNaRLjJWRtHHqj
JdyRGV32R+BBUrzRqA60peYPMv462ohOP3p+7/p9vmIz45RkBHGgbxhXeZ2b1W6i
bdxZjkDMGMVogq03sqjcBAZulGQW6wKHgtYxRNZlNA3c8JAbrNCEapXDxHT/qIkC
Ene2JXjpdGNg/XYroOleS+8Kly1exxanOBdkVLUh2vSYbJwuLInvWvrmjyM0tgQc
GjawIirPDJ2ZoTXboHspaUw4Kq3PvboRZG9vQDDYUEeVjuS3VwZ3+hEXDLsDAvo5
dvsKsX4uxSwvz/Z7YclkQZadnK+locbFwZ6i6z4vsSt82Nc8TquctqKf+wWIPGSM
tEdBmF9E/5mA18CUcekA1FeQHERFWYPBOevbaobFrsP/XZ6zt6NtwAlmroXyRkcl
DqhBzkgJuBQYQnoa7m5+5pLxBl8n/cOfnxXLYpm+jdYQtm80L0tBGfcnmf6fyWNq
wKFKB4tMm/oRKkQw03wyuEVX3BBoMmH1nCvH3tCJ+kwSZBuyOZKqYScterovSNXM
Qg7uvpoKkS8mQ+3dQ5SYJEUbzxrQrZzUNjtTGf/74k3/EdCAyvlrhED/HX8Jt9Ao
m/GKPfcx2zbS6woK5VtQSMOWXkPg0XwErSlMA0jQKaoKfz2LWp9qkf47ZIUuGfYe
5JkgypNEf8xkwxFd7KqYHIzq6muVn74CKU3GLr9mhuAFd9F5SKQ0K9SSBi6EtkcG
KvfYprZvxfvJpZmxTcrdEiyoQgF+HKKEGVu01mMZ/6ljsnFpGqIyJX6J46plr1cF
cffjIBVG9sh//r+CXlduVS87MiOwDJlY6agzgPCO6umrOBHPSl/aGxYrPSI7/VDh
B/4IpTnbIOfruCsflP7MIHDz9aAC0/wumzxXNg++PhA7M6y3tNH/aVqEiAXey7sK
dKHk0FEnLSw5gbQUK1YRfMbuxaPRJTOOsA6HC2JXr4EOMubbPlUU1D81GAVeur0y
gkuOQStdRkskioxEvD9bisbUiuKXK7wvkW4mG6ZoYrLI/1EbyqjP2hv93y8deJ7R
TKfXzwtWlB0CT25PGzFmVcl+azoA3gNagfCc5VSiaoZv0unYAf6w124ZL8hiRqu+
Kt3a3jUDe0aMMpF4YZv4FWCcGlu/my7aGdvTNc40bOluD2ygB7XroifyPhe+Df1P
ShVCbRPWE3RnrcAEysabgs/dwW4CHuf8YXWPzG+itY/IsHVePs6etm40UA85sbbt
ZzGEuMVzsM5Flb2JvLTX1GIcK6+U1evZgIhygy2FaHZbkoCb2yW6yDArW9qkXPqk
l6Uw3hODnwpYuuCV6KmCJRk/Ya+I80vdbGm+z3UzImMo1YjH3/GeGsiz1bj9KNbi
CTJtozMx2FSF9GA5oEGaclX5x2sMRoKYP25RDtemTB+HoP45DTSWl9bxMyluFfsD
yOie8zulSF+Mdg9T9QYVdIKSP6HF43iSIWsBqSYoMVs+hDPGg4oVRFSV/J2pioQ/
wHApbvd7zXeZYUENrmaabhyo6B2ecB/F5vrbGmRNJLThZgVHTIddYq3pP5LwASSQ
QK22bu2NpNqs6SiQc2426vkvp0Q/kXy6iWaKSUeqJ5WAC87gVM2W83kwYkfVEV4A
4UXNBt5Mi2f7FUT23PX8YBNjkQ499aDwa5+UdENjlAHw4YjOC0jQ13EKYI4Q9UNF
QCZDvc4KdSOIBizi3ixiB1T404WyO75+8fmT5Upr8uPMOF62J0Eb+97HzWtBFHwV
9SHtawxfdSqDC/+UW/ekgFQSgEPSPqEbMYVC4c41dVOg8z/pcgMqlTOimxKZxopJ
yxV91Ko8hw/0taiBthFI28zM0BkC8BizCSTZY9agAJKnxdjIRzUSiKVcXh3pk/iZ
CwX+S6LyQPPME7hAhnvMZfhyk93hDnpL2ZRyf0D9rXvhuLtr4JPQhOM9IJLPZNt4
qJSGLGw3MVlqL67h24NTuOk+sjMf6dhd93SiB2SdaXX9hclJo3ZOBJiNMdNVv8Rn
DE4elkw7m5z0K6jfMBIGWLCMRVWUjxCi8BrS0X6lYYDy5Yl0NQMx9xW67zQE/YH/
+U6n8XzCCqFshKmhHSOG/Xopw3L2uJUddr+fgKl4MsV6KD/ICfqagYUHDFQq5rj9
2h08PQqu99D3IFzqrVggGYUudrINZAR9kUBAiDSX4YkLDSpp3o7L4MY3kY91pHhi
MlPkNAAVN7StD2abWW4lM98tWC7lQRPx8p0C8agntGXHZXhsoBh2X2i/wuKZOhvj
10PS2+cjw3HotnJIS2ygGftROMi2geLu7GLxN+UlDX7QE3sDVjfBslGbpMPy4L6P
Zr74/Olp2hreqtbaDMyeUiz/Pxw8P13lc4Siqn/KaMVpzb/uSzXqJ4HSdd0HgoY5
Bev57LYBz3R5xmr1dnVf3oYYdYncg2w1fe9RgP40RdUXVLyrHtr0AkxJkDZLZK91
2dMH0P6OsdJzyDuzcxfxWgfaYyo0mvkQK+zDI8U6h18XYydlV2M7JN8UjEocve/h
v/4KDw3QsehHDRpq2uXPFKiJF8nTIfNsP8LxGb8GhhaHZQ79zjHD4f0W1dSvd6pB
BW9GrR3nqAecHUIwtjueWf0v9g3islHChBWC8IsWG9JtpPSUZeqQMJ5DVLw2yqGP
12g/wp3AfPSn1z9s6SQ52+8fSNUlC1h2u777dlKwdMBynlpaGrH1lP18yx0Sto2E
3RAyQKHsiOv1TuGIdjql1AGsKAWQrZaVe7Vr8RG3jxrxmgPM4tDaHxQFj00kzUXl
P4rE8szYuCXl9RhKPZfuz/+rZid6iwGG52xFR3jwrItu++4Vh28tLNJmdSILMT3y
n6qit+bb095eoz5MqwP7mwJS+3H5ah9zps7uaOPWZ7xAWsmlPUPzrNffLC68i+jF
APK4KjEBzIMPn3Io8I7Rz//thd16yuA+nuJGjyq4aUf8FF8V4xLye7xcN45hvaBq
hSHRUt9yUIz7JMebwTgBAy1MA4xX307b6GuRcuriD02JLBHJQ1WzJWFdVm+3jzOz
Syg0UshqjYC+kCXZwA7wazNkuFf2YCtnzrmsIAn9p2S23AkYTSAToDk0ujZ1jh/z
c997YgSIo/waku0De0ie6Wq+x12D5Y4GT+ApysVsTdyIJVBzrrL6Htnz1LSPKUR2
1lHKfBCwHPalgI7ksyOxkDP/GOiMCEgiWGKAOmJ/Il3izsQwKZTStoGeYfd7k98E
ZMcCt0gSgiOOkFHJktVzrUhOGGwsSDLEfsgVCJUaQORcYUUxepSAefIBrM0sFgJK
b+/BLF68NAOt+d64+5ITUy1GBePbNWLtyFteM0GCADVPolIAclq1X4iwQXIiUVRL
XEdSS0U7I7JGFWQfcGnra6xvfjuQVipMtycDuKuGs4HVH1mv0lRl4M2t/2NfsM33
Hljb/0DtlIeqPmmTk6dAKutwcCb+ae/8smXvQKGthVQ7XN/mVhTWtlFLTuUVEyWM
71j0qcnvNjsGOidDMMpzhSwi9vRtP7mZv2nfuMI008RuLUzjLz7ci51dyTbhYzpA
NsVW1lKv4fCw+6jntz3OSI/9DI5GVgdgTXjW0EiBP3h0/guONfaS6carYvZgKIXb
ilVYbLnwKarNcjORVWaGeiCdR+tBILq30/mPp/B8TDPtaNhCXmz396CKFtdoDNRm
RN/nCVL7eizuh6AZ1bKBConPfPiKDvBx3EdO6SDfr7hHMWm0m7KMAdS8jsH9CnhK
mJFPFh5F/LFhPpXuftnuiuAjZxOUsU7aZfq6eSPA8cCy3AcFVcwpv93rtNLk91wi
aBy1Q8oyOgli0pYL0VskDPjOFgoTUgCe0z1WAKzerGM/mveerzPA+r0fr3wyVTcY
d76CEswddv8uEXbMtRdua60zRVYE1oY8ExaNI2/y2cD1UYjqvkyLiyHFZTLCJMHb
kXNlCzgKwhi/LR9r4AXrQqb8BcpiUm45p55sK8TF+HuGMk2EexO1v/YjgTdrY9TR
VmbWlhmYSqugOTQ/rescn09JnkjSBrRJRR4haHR8UjrGqgyxEWpQqqEXoDPkngbG
9bhtSS1tDlZzmf6law/uj6dtWLu8sp3qVWIZHtW6I/kN7TcATmjK60aQOa3O+TV/
fqelXJLFpma1j0NkoXUAO8b+CSHZO53h38T1Ig+vaWVblj5dAVxySi7f/CDs8zvl
svWGAGP15nSlmn1yi0/JtnF/MzIjGS7es1XXh7/As6jzJcnWzCa4Hvl9SW0nONGh
01fpVl6qtzoLKOg5rQDOL0jaMeWU9jbfP3YOs+07oO7VyldGKlJ1vomwVJWk4eAb
zS3V/wvD3iEdgPio203dJGdNSgiD0VrVGucPETlzYgD4zczRGKt872SNcuu5xb6l
ii2viYhMfM2oIkGCSdTlvLjsf1St5lWcar5fEfAw2UW7nbq0tzD6cbQ/SxVyM4Gs
o1cQ7vNRRf7LJOBMJ716aTwn1Z1bWa9iWsrWKp9wBslKdHPXcZYU6qNj3N6dRYt4
knqRmd2bkJBmFB9CpgbkuWBvDSEJ5eXY0n5xwwqY8ZESTgNPySCQdmzD26hR0loK
TlC24XsRxU+QRTOhBAlYmjGUeIVuELKiFS6bqX5jceCWP085TIeYIROcNLuDEFWr
81IXsUSSqBRhxHyj4P6HF4tD5+nhBRjZ/QpPmG5im/E4hn1ZVPni8a1M2KS0F+jK
Idw07Zoq6VzWDceIBKJaXDDdAA8EioOIqHu+zESiTC9QCjYYX/u5r98+wbKgDpNt
4TZK+Ozcu6Arjz8tzPChoekW4gKjSpDZGPF8Q3Kz6VJzDf0cjCFWdEIxMYyS9LIy
ZvKr1JOeH0zQGnSQ+LgEDBU4x/u4jedoEySwtBmNwlmqBdJVGrYSHOPBnUVl7yQ0
4LoNY/dCJIM43c/6myviUCA7yMO8zUA7sbMc71uZENiFYNAicrdZ71JH+84Updmr
d5jh9PCagqfsnS1JhEfRUE/QGR5OrqMA9GQU2uJkxLBK/puaxsicAFQUtSuXnhNl
vaAJFzbn+5SpT/AJxZwhiiKilDXb+X2xv/jp4mSS1MsDzw6Q3C5Jhh+4GScWtWjw
g5S/u189slbwc6NbGfxLkDGtbERIll+1Op4Q0bwAjMG6k3hbNQpvnn71RpEH6wFe
evKewjbRSsBgoIEhomzMtR1BSUTOS0XrfzwPykLo/IbSJDs41/EvjvG2uhtfTV4S
R7sniliGtPq2vVDwyX7B4jrgBjggJq/LJhYz1d/cVRHOq5S1w84FhkZhORhIEE7/
njk2Ml9wTJlGiSB09H/A3ZSkqPAKZqp5QAFr73vjZ44A6EcAj3h1a2seUnCjjuu4
Sz9ddLmGWuQ2ALhhwKsLc2NIqmC9UMsVu1YV5NNkVC4ttnT3t9DIdECXi9A127pR
OY84/2cdGQ5FONUEAqxG44SSWTYSTYMTWX2TGeKG3PLnaMalfUhPU5SJzOXFAYy3
FV7YZTzvji+URQOwf4pPKycHwt2vvbSzBY0ZFcFtmYq7gAU84fPCPa/nc5xj+LGx
xes+pwibU5v0L258S1yX8y4Tgp4bkd5g6gNTRpTJCP285+jjbzL9G++z5xO7K0a5
aPnGz3ILFmbbZ/wU5tGsfkO+HmMvKzKbF1LpZnxDq0XVzCwhF8Ej351K1m4lhFc0
zZ4w9dDkChJWB/vBNjrHcv3wAI5yawZ/SmAepSGyfekVM3+ZGGaMxnHc0YJUWGIV
T9M+PwlP/oB20hL8x1cNFCkiC7IsJFh8NjDyAFGO6d9tv/elnp0hi4LoR5DogGZH
w4c+T66Yoi+8+Qjot3s3qs7J/aeK8ORz6wvM7KXKJrm/Q3Krg3tGE+UFoh+ZvJ4n
vw3CdtqjCNtWnA5cgmGTmeDbI0gtKtrXqVfqboxqZ59vrzex4XTcYWxNvhUgbPGT
cWWmhilc8rD4VAO2P+fScIUU5UmqqDySAoIb7uLzdoc+LyrEAM3WhCSeUmrFV5y9
qlyrswtzJzhqcSd/2BQly0jUHT8L0fSGrQs0Vl+wJCmqCPwC54Y7Jv9lkKqdEiJV
nbTBtdMllvV5dghD/11qy/TYtSNuFKipldOY/waKxaFZAZQhylffJsrSYSY5JZ1Z
SBVuVg3AFDQsDtIKDfB4zsPackrY9chdZvllobygYhepptoStb9Yh40eAfpFbkV5
4lLrFfIjvfuxyoLSQoL2Mw40lRvfRXPqbjJMzbAOB21XaSNwdeq/c5xPw7KTMsR6
d0f+gxVTZWJtaCgiJ7ofccwpr09WjeBUA99TP4qZSUHueH2OSJGd+u5xSB6B6dm2
pzQ7Tf3KwALiBvdHAO4SkKrSup/D5m6qRHPF0dQtiMD4xEcdsTyk2GmNJrSmosFs
n2BqY7HaRXNPcRoWQWqm+5x5gSfWxWJLoJQ9jMjugFQsmWJvcR+8WfJTKBZPVpdk
zjLk8uj//PWdRo3giv+tt4+AxykR3Qy0Zn1Sm9zdyDEbe+JiO3c+uxhAHAy/iuC1
41WPJbbzr4HxAdmAyqOSExOwqOvwmLmssjv8ciKSE3AqsHHlvRdshxsGkTgc6iTj
LFqGdP1FNdIqdPvBz3zipDGhweH8PebnK+M1P0IKaQRXH3FZ+ZTdbfb7Pna8+vZK
KFzGUOyVGIPMFqLBH/IpRIkcKrihXCZjCD5BrBRmhfuf8cDhnXeUYl9D+S/kIwrX
ge1S3RcWcHkktYCBdyyvnBW3JDLcBQFz7+G+3fWvAqVRKXsdtMRRDESe2YZw/TCh
bVCqx4F+3bZD+FejsG/5FMWV95MLMq9jwdGYqYmMol66DaaQ45Y1N6Ww7RByQ4Jm
BhBBJ3LHHIW9i3oGl0vMTDcw/w760PLLLqmvcyrO8TVRcXgggG5zRM7p8SwiT3rw
8h4IFJp6+6utev3sC8QM5QafQK7PFU7HdGvMtVi0MlugIaOOR3AGzURBtzX/f0SU
YgsAU+EF+YsWNi+xjzw2PLQIJ/3ZGRu9TfMxAIif+oYNH5pcsZYCUXA7guxYZX8n
lbF3d6YSYuE1ldm0a25vGEgwsuVUROIuDCUZ6j20x9Db7WFZ+2q1+QOAqgGNgIfI
t4ETLkyezpnlqDSLnzEGaiie+A5nV2XZWv0V9QL651HLd43gk+07LA7N+76lo2Gr
UbDM3HAXR6MJXX1M5Gjzja7vW9nZ+wywEl1ZwN5QLn7EX3KbC46mwloicGmg7A+G
Ul6q8A8kvP/MV8CCageOzdRnwAy4AeDkCXzh8UJBfXZN5pczwNBM5CL64x5Pt2eS
B5EoR9jDnKyaXYawZWlT7JIP1ghJ5Gj2JmJojMe3Bp5IxEeD4TwRPMA90yTcI1j+
ELnuTARmVYo5YeT4lnjQem/z7DbUvQ9+O/lbG4SS9V/j5JmHJWg/9JX3Nxw9Ku6z
HfORJDebSsPdZnPXZXeAR7KNprEsdmeeRx34ISlsX3jj5a2kzUsXq8CE2mXxmW9r
dxIC/4HAZxx999gcX1MMZf87GzxPWsBFNinzLod8OlaGTn3/LWLXBWKUFTA+51GL
sJTogCUzktPfvNfVsgf84oY1l/TIEDhUZ07SBG7DqHvpFWHOQydnrB/kao8WDeiQ
doxCntHd7IiNHoESd9lJbOMgcrx2slyqOjEZSzq13sWYv/R0zKaBKq+3hPviHr0Y
KDpmvcqfNc7yPZDuh7BpzqrFb5BVYUq59Eg4bEvTspX1RXE4Sv3busmXT0u5FrSU
DJqPxi1ctLDygIr1cC7rcdId+A6UFdI2gfB0wqflZi6DWdt0eD9TzM+GXwRV1so1
UK5guPJNR2dJUXrBsOSFWI0rbFNhq+WuYUtJvs4sdI82uVSBdEmAfoIWNd4SF6TN
5fu0UouTTh2hkDBrefwwJ/zWnECGZF9KBWCvIFUP/9mxbpTiMiWOYPV7SJMeS67K
E/dCwzM0UQpCUfY4oBd7nwAiS9DXx33uHDS5uOGKqITt6XM4FCZVdeT0evnQ32Af
8oXA5gqFvwXhYrZXR/Hzf/vFnEhqUpmzGQFezMtwKcNzvlZ2xz4AWa/1zIstM3R5
fWGwwpGBTlmLm9+GULy0p36RU7zFrzWfYH2kBQqbTWEJ7UDaUVnOluXXE1fIjL3T
cmv12AOFJdkTdWQQY7F+DPiQhwFH8YjFBmN2M8lqx7oT1/vgH4dYfbya4rptJ1KZ
kuxN3qUWO/1+moRo3L0nLzek7iHfPBLxen92FIbYSNrcH4IoXsPztPaUYVJfwmWQ
T73hHLyzYC8ItcrFhU84qIAG5vXyOY4BO3HljYYbW4DwGXWF2IRNluHkYRqIHeWn
gQtyQflYfcBZyAZwy9lQ6BHbPZglNEP0SGnORnUVre/UYccmWtQ1pSnjkB+V6bQj
BPRg8L2S11J7uchv2/i21iM5Wg7kQgghXr/F8rzluvRHlROF0oLRfSiHP8/8Flkb
IPOBPdjNtm9jFKmoT52cIIV0A5ZZ/xXJG2+D7HCSuVLCAOLcFoM0Bc21IxsP1d6h
9KO7UyFDXolwgCGS2GGcJF64lLQgdBePdOHTG/k5rKOPdaKeehzAxNyGMdjm0gRQ
8nhaj4RQcpA4h5sBVNJTOhDByDIC1+ktImZDhRSeyotrKkJmn7INigqFvBSgrW7+
PyYLelkU6/OHTVyMLil+oU/fWe2By2IHQ39CfDNuvtSQ3DG+2KoThYw+p99RJgwi
jPFrc1YZ3hgpHLdb9Yv+/on/s7VLLoz6pl1vRWGeyywjhEhuvvjMUONDSDu+jYME
MT2LbymjsajIl29rB2vnql2gTloHumFddbFP+TYJAyRG6ODOrmb446VAmFNUdbC0
hZg7mobyRoLwW/CdDFAmeCAC60Ot638BWlOS9MsiKWCozRbdknfLuJP/lszOGZ5n
u/M9GfQo/y1d6bEd0XJHc0Z8QnhauoQ2hF1BnNbTTvIDMs7Y5YYPqM0oB5Zea+IS
yGpYu4OcltbIHoQGBGyPbNq96HVa/kf9+SGzuDcX+f+uQOpg9rfd/tLWOo4E6knF
4cBHVQYbj6Dk5Up5BBuYBNxGIDiGYt+6ON0PvyBpElo7TCebPImDXx7uzezwv6mb
qfd/E9wzox8l5y0Vv5kkGK9JbBGaWSa35NpfvwFeEnmTpa3JN7lQtp4+7BJg6jtl
fAYJ+R0Rsq75pJ2m4iwBTuMYNyrqXEwrVaoHvfQE2Wew08kh/ZG/nHaMlZ99kHmr
SDvZJ5Y1Jk1kZ1vQ2SU/vTRr53CAp8hHk2xp2KogobB6NCnZzmgNfJ6yXRpvQ0O9
MZ+elMgLsWHfHRBrDRgkFTPHEP4nohKaVYqTiOs9DHHejmmcJsmdwPZUoX3JsI55
ADMn+I56MVkEtZfuOo8rI3gDwwnyZi/NlByHntbh+DuXVaMAkyKN6G+zZca3zT+w
fLkawn4+srslwOzHP0yo7vjEKkJlMKYgC6inyUK4lt7B6zFoVoxRppklKf/P+yRd
x4ZXxa46sfJZ3/r+YugsuJIQ0E840Z5M8dbp3Xi56g2OeUHQ93xE0O33tP2/2w1d
VF1xInSYel0F66MPy9h9PSXla1AccRV29YBxA7TrxZLdIz3Hx+l8q2pODjUjl9zv
9KEkccAyt3a60gd2ZnVEuvmRmm45lNEYg9RhZwm4AEG4GFA7cssqg+VxHe8eVmD1
2TJe/fGoGE0HshReOEXPUn6Kqx43ihQIcYWTn54uTm1VbdywFWmZYiPANRMfAmnu
3yA9qB50X985Xa/ouz6cux+8qfcsRWtuCfwdiQNjqiujk5tYaLTYMJ41mVvWEotT
faMjVO65ZsT0cyaagfxMboZ5cNkPz0Urjr+HS5qXa46V4U+c1yuaeq65H8f6VTxm
QGYFl/ydGC/648pa2Pa8psvlkX+NJvR0rNRGYiuP2QBPUmT8REG7CC84PVLWOyAt
1CKnPQMTGQ54DBFppF95agUdk0ofPWtn1yVMRWJ/DS1MRelISTzu2IYdDJH3C/WZ
MXmcE4QjJdNwEgRDjX16WgzE/xvYn8qjKoDP8UEhJflg4uuCGBAfjo4RyGbKXnvi
N2Ror/OJbDdj97XmefjjOY3LUgHYsgfyHRF1Rie2BaYK5yO3qgsr/4+o0jJE84Jo
/gabTzBnF5iLOPthjp1/CQXAPtNb0eLnM/njNcz2seJgSASG/4pc35YeIBH+TB4X
FSbJbLkhO4Al0rQHQ06yHosWiHDyiF8yUIEeUHl/beSSYUvRXRqrfiW91qtBwcgz
vHvWna4nHWsaNXfUN9uImOwSe/Fx8JBFmZaMhPvZd4ErICQJkqNZrBOg+uqoncdG
xx0fMn5/ccqDRokaDpNUvUMG9/hp4f5XwQD5MehAIuriBgGZm9zL/w7CBsr9IiDL
L7d6rlKBWVykTF16Ogbybqubq4UTSAjD5N/hXnWKJc6MmEPzwz+I9vN9/AoJ9oRb
xDuIR4H6OAmIgWqO3Pq7OaJF066kX0QLowTtbAtPT93n6wtiiienex/EvjMVKTKd
pIbWfTzd17dsBRxmP18mCxDuUav1Iny4i6q3XLYxFhI2tZH5IjwtHSnb0pJFPRDA
usRBuJLzhE2U2arXX4PqE/R2nJrEaeYUv8YuVOGlPLfi+Fmye7Cn10oVGZ7QxG5x
NspguIcjGMElESrtWujo0rIW+YHR+FAXoVxy5QdpTzn3XLpO5tsYRt9QN9sle1aP
9l2MHs2LioSoean0vEgDGpJHwKNbufNjbMOkElp1R1xzzow5wXnTbubZELxEJa2L
W1K7UWdi+9+DxNxHqzgso4nKac3hL8sO+OIcXg89WIZnP8YwHINGqlQSPpsdeBQg
OYiMRT34pycGy4WK79T2fSkLHCgA/IL5U/1TiFGeu9K9VwlcprUAlDbXsGZvY3WM
lWD+zpO/ZWpExTwOMOJU1Zuf+a2xO2yPKXkQ1lPe0z8oH42wQ+6NgmlcOGzRCNjl
qKRrpXK3RkHamuPE7oxmQ/EspbFVvngBLCmkBvTGCLSBFHrJQYduYhgBaUjXyfHr
9iaQMv7Y2m7M7uMA+e0w+B/7x7A18y5L6RuuSk9GWHK+LZlug6Wj5bQ+GqqN0Gsi
hfWXQa9/Sz882Ev+l77vBANvLbLdHuYaDJPNWJESwANruzj4A9ohwD7uybN1DKH9
1bFsyj1bbbOwvdaYPnzXfTvZQYHQEf7FEt0/1om0HfbU1YvEYaMJ43PySArx+gQw
9iBAZYCQ6JzePB4dM6Qt2vhLdCiVVkV/l+wmPX87FaTOnAdHe5WnQkuACKze/Oiy
SYcBvB8iGORsfrDZGlDfH+31txDRJB7h8QKllt6H+jdLi3iYdrCeLFKSj0vYldoX
mnZ0NkKmshxtfaOQwQp8Ed8F3ktSB6YlRDnPQkFGuATeXu2LsKpuoRMpFmsrkzm+
yk93j5un8Ak+HaQxl2peaaadC7nEPAg4Af3QW5Pa6Q9HSeaaa1wY/vNzt6nlANKY
dHenp43Hx7yK4ISE+/Tp57B70IUI20U5Jmr2lddgjZnMpsQdQJKXVnWCXKMid8Gp
ufY3PQ7fNy+QC81dSkn9Tc5lvmhAR15OTTJ9uNymx5u1M6k7ifp64oHxBRxmsHyP
MNMhHZ6DuS3AdqIge8zph+4Oi4RTLRfdsmYa85J1FiuK5x8xvLa6OMRGI4HG3OSJ
yTjsKjurpGSdb3qYHwKNDtJOLmGKzZhtCn6bcNyB22z3maJLDVmV7D90t8sGNFOq
nYivYsv8dNN6CTnbstD2mdKRnWiHmr2UvnOWVUrx88C8yTO5EuNG9z1Ylxw9xM5m
5Aw4NkXkmVifJxCc1o3/oVyYGyF10mi1unOYLfBRfpKW4iwfusv59gjGYIyVT9O8
gcaPsxgQtP4fWkO6NHnxprZ0weqRtlvPmh45vZ/JHmajbf9caq7i/qsjV+6EyPXK
Mo6Z/ZPkuQZIze1cKBDzwm/0IT+8V2U1pBju9gJEyB/H1IkolS4T+zmsNllPDNLA
Fh0z2FDWwk9ROdmOjW4bEOagVdHanK9HCh+rFoC19XCraLc5AjVL5UiBmBpgE3l5
PP02ek5wLWd1dXva7vTLi0PzNeF/ytUSOtSG6QzigHI/wuxozehi2YX34VlQyTsP
/E9wddXv3SVVMsnFygyOzrrh8CUZoW8cOIpC54zOG3EmzyVXnmeUujDz/0V2vgSK
1SM2sg0Qy/OFYLOFy5jLl0T+QexW6xQU2MwhnAdejk+FBy06qyqPIRkxMfJELmW5
RhY5wfLI65ix7bxak/Zszmrxlo9S1UysJyiuzsb6U3BOB7Gqoy8gyyU/g6kz3MQq
SShyW/S65ZsqAgd+Q2DJ7WAgJ9CmGTefNiqp260VKjlDl6Js62Gd8pZLtCfb2Ghw
rPadi9+trXIXNskag0xN22UXfLOgpoUQCuocOojOnDg7Xfc/cEmqQdsjGYlbt9Fu
gxITG6BvH/RpzudPyphmeq/AmnhxhbjkECdbNi6qdjzIRbHPh4es59OnSJfxUogh
gozYGnvIw+r4YZO4Rjz0BheP3mMf2JHIX4Yn9FSt/lRzuROKP9b/3vUA/PVF7bdn
6eWUuI21fU+WZ1uZ1CWV+env5nZ1fMRcQ8ljWGl5AAOwFqsXwci1ETqubrPfjAvj
3aezxo2DcVa6Ml3LPGG0OePVQtJ/JyoThTJHcokYHedfi61ZmKEvlASkpFxP5gma
qW4JO1oOEGuXw/Sym5nlJxY/jDrHKG/SFPEqT2QBc5ExMAYYIEdXHd6xOx3hIpds
oTBvEGj080VHGWm0JIZEHWBEE86f1mru2aRKEr5xAO28rQdfgbtFBwvDV/xZ9buT
zZnRyUNof/nw8+YQz3F0Dpu6OzzpFDj10Y8mXu9U+rIsmavE0zTZnXH/xCrXj2xr
FqhOJYTdIcVHt+1/Q8Q43MO6ff9PtShWjVcmKps1Ud1D2Ojk5NgCqo1NRGuuxugR
lsJYzF/95Os5hid2T/WoxAQtwA6lD8KcYiK0yLuTgQY011FTSdcAfyyPbCXVBd5z
AElrmMDS8IPbnEzwQ5UIWSNnQ3nzWKB8aw56EJ5eSQUUv1eCMy4zHaYmakZz1fVS
A0Qk3zNE/gK9wGwUPLtm7CQkNk5u17o9LjWYz7rcclQk9UByz1HR5isMggAUL5TU
8Mz0FRw5Z8ZRBkeB8lWztSJ+b/44lmIXDC84xoBt7ZaFeOeBtxTzmZG5v4jczJwO
zv5Xp+qt74IM9T6JESEL+/0HtKzM2sQ7xXheHDvMglcGAk4lsPJgBXSbfku+vtLg
kz6mvni/ofPjnh1GXr7bbTHhPRFMaQ7qNNN6Qengre937Rc7xe6kVAGXb5SNY+mq
2+uQJU/IWaWoVzw7ZRmYn66bM3UqKsXgpcQwZiDh2UENqgEqbS5KQVu3u+jH6bmS
AjgeErvmIcbdaddohqOQ02xKVPsiN4TtnV/AzFK+xaXBsRpBvfpInjyLQ2S0gREB
1QFqxDhFaRECsw2HDlcZWdnLKaQ56j7vwcDOAXc5WGBd/UtFxU4fDnnDn2cFwfta
/Z3hY5kEZaRxG+M/Shla1yYdySYJ5R8Hr3p9GnBXOk6CMGJT+96BmT3HGwC2cC6u
2kYGu5vGYeSiM+/OeQTxZtchC1pM+NQwipXzNwj3WRm8GbWqbTSzZg76HfKXehQv
K2r5M8Ue4wplTlR+DO8auGJ4hVkDn3Qj3Yk7G7eYKsHDWZlDXIv8v9wc1pS4813K
h+Jh1cJpJI/QzoDYXrvTG5XFrTgTU3by2TsgdfQs5ZAvYHmMshXtzkc9/HaoM2tB
Dq8nwTjPpc/rt/q/2ORYtTH1uobJcxdqHkEqWbGc9YSwSxOpLzgx4aFnPeVAjf2F
K2puBovxQRDnNwaf7GeSdQzSwFhAJT1UxIhZ6IXN+g94m0uoOpD0R9SS+OsQzwpA
NbUVjacgZ9aynNcPOaY8LEjnW2tppkDxrBRsUM/bWeK1jr5mY1j9vjpmCp9hzruh
YNfr2UgKdiO4PVREo5D/dzOiXTRWEUMbHDCoZXe7J8RZ+YPWoP/dPnGNF129ynhP
jYPGN92Ym0bcScUO12N1mjvUH9xS1kJTRz2NKOE8+7CJcwgUub70q3Cr+xMGgFAy
X+53zxiMd+xevoECnJH8ayWNmCyE09gog/YKwhQa1PpMvup80gzgnlunAv5gyqiY
99dvdL/9YNsk6KVNOCT2KxUuhEIZZm5aEwkuyFwS8h/qCE44bRuwcqY3/HxdXzpf
rUFJlRMXYiYlzp+fSImPxxdj6yYwhEh68L8Ape2Tck0QPAUa4XvmuLT8ZdAiLUlf
WhAWab5U1Jux+rYiGGKYECctaWAa0U4zg4akU8mA9s4fnPvxOsBGS/Wz0/hZvxzG
yL0vGjvLOEHmEccRTIoBV7tPB4lvmIb80auITpwgTqFtm9iukvnFUrVp65iL2ZlS
PYe18nNXGIZQUEpygyHZG91iuu+HIBfVfUezPOUykHlI/NVE6FRG3PK9wGpis7+l
6qgxTNrAIGzT5PNZj09gsIZLjj8VcKqLaItGo13o27rel3WkiN/JpggbGJKUdXy5
ZLKb5J86WN2vKhytsJwQemNWYfnKClIhD5mLReNbKsqScZw6iXJ4lC1hfjwgDYiR
XAyLRqgIMUQumsbwNDZvbKqfzt5F4Ss1FavjAPUwlRcKl1BMfpSu7luNWm66eR2d
m5djEyIcgsc6USPWrmX7nvIc1IRCfDswZnjiSNSOOiVgWmkmZcHR0K+/fCy+hgHJ
OX1Ayw/5xMYlcNa+gk+heB4Mj8X6dxuBh71Er7owQFdyzqUnPfmsXyb9LwoAOKLH
FjPbln7EKAWipQI0W9VDNZQdztJiQ3Jiuhdz7mvW1WPKTSU4ZbP7hz+AvV+z4OO5
1cFqtmuAoR4ZqYj26QytnQvptZ/arwTLmE0bmPDvwHBIDLLEaWKUsck8qpdYH2+0
rtTSobzQ9nUaKgelKU2qGg9dHtOhJnvpkbZ/5WOxeCC30KDxlAj9mFUqU08QuDn3
8CYIOxJg9gm7LoAEkQk5YPAlI8iS8U72OTd4DHqNw+0D1cOvdAxQ5aFv1tg4yhoq
vqMJ0dc0fdPk6IWWa+vNwfbmGpipS2luK4k6y9w4A1e7mbe96oOv8sL9IWJwx/8g
5UygUfqIVthyWI2bgaCqgJVqvUrxm6NriPSTSaJZuTCLq9CcUEmDT+k+E5Kksk8B
E2fA2LkyBPMyLQzFC8be2UAq7HPsj2VFjSTN1z7tHgV5Tx6ucubFYYUNKIUmgYML
zsiXMespMP7tc2iQVWRXRdOYmITNym2asJvaRztucQ7KKYLyIFdxUQGva73CPtGK
oxwoea3GWuybVL+NoSUqJRkTs65PQ014qSW9O5p7vCTj3sM230jB2zoRSSDI9j1j
Qf/yZjc7DndPqzZRwLHge/Fqs4rTkpQJJcGrwhc3px7VoZc72r3aIqM2TgUoOuH6
xn+4/r1uf7DR0ltdGQ4ozAtMgSXSWEiXUIe5+E47DG3E2vFA9UxNZVipZFY73RBu
skQnbm3d4pB1xIJwd0YIdI0+ZGt8Zeb6Xp8oriG/zaLXm9BE4Cw3wOo7Fp++X+tJ
lqw+9nES9UmfcTp546kgfcxO418NyZWpBLWvLJa3w/kyhkA3HG5thlk4S2yviDuR
t5R8dyY6ThPidCZRrx1oDl6PLo0km1426YQ20x1bwXe9SpNqZ4mRYu8ENJqDe9WQ
w5KN6aBET0TWoPCSyoEhFHuuwYt79d8Cef2xRfaBUHt3uASbZcc4A0VRNLWKIvql
rO9SoSLSMvMtxw/yv8Hvbjlna8/nlafNKMmjhduHg7pB0ligGCDnyd2UCobTuHao
xmg5bvtHmXys3QGDhQnZ/tApwZOLIog/rBTW/lCMbDKpimjCYatm3RZZol2MfyxA
LG2vnOKLWhSMsJQq3depbkgWbvw193PgpnLWXhPcPGxEkVQy82T3KSPbJHmJyd4K
BrhaDKHGeUlb7F0jbZh20V1gyvGG2IuliuGw06JcnHi9w6+JMkE05vvmo/8Lia8z
VWU2dXwET/O80jwHNaspvLgiaL1KkXGsg7CpTgTBgcKSNN4lh2xvzzbvxFQiq5Vw
45FJn7URG7a9QHHaSWpGm2HPb9rIBWFPESl8aOdscbbuYJWgi6Aj7+22IbA/EGAP
Uq/MGiWA3n4bvCKSK2ieMzSPgXUGktnW00PM+eXgrRRP6zQfvTGv+ZpaiOau+Ucb
clNNpLWnjRtzUm0G/0VUrLxpBHAiAJfwcgSg0Z7/Nna3IAmGghDtj7GkTEQ9BWQx
koMg9dqvDHfaEmNn62HdTL7yGQdrVWfLTwfiV6uSD53nb3Cm2+v+ZPjBbLx/eFeg
P0fJ22PQJIb7C3gdsp2q+ZYkmjTyLCqDXu5orsL1ctFJxI1GEBKrUu/sdVtALuCj
ahWCHLnybOTrnroBzdq1eORW+nBuI7gIakX1tqgxniNSCv7n1PcnongO2aJvhTwv
kWUsdaH17Em/nK24pd+SQp1uQaXzivWMhhjjUX6O/5lmfcppz4J/QoZB1BIbPhyZ
8fLmG7EC9zbPvvmD7lLVs159+NwxTEQoLouue/wyZW6HyuGj2BjaVsQZxhdZvIHY
U0kRW+A/QK/kRZmwWDIXZcL3wlEIMGc0ycUo0FVPj7ixZOcydl/9dcxFX34AiQxQ
881DqCssS/MNyy1hR5DpWPzHzKYgIU54zuF2df1WgA9ioaJHWQJwQenvlnz8fG2W
Ses5z+fN0mCx3yVPE+TVwsJLK4sUujm4vM4lopCQfiH+NWMGzLvhDovh9eRPuiRB
85x1421DLO/FgZv5I85FyRqlgetqGp5xyeZ4O1eVsmoYhEp03V3Ic6pjVoA0qeJ9
0HdZP1zytRoHv9jLYrNK7lFNRSoLl0J1CcvO7FuI/2h0BG+SGpdu3vf8AVLlyEil
XPP9OdWgHAmds1/gKnjMPo/VIzZDoqhcl5lUFvIU+0UbTlQAKOCnkKVw5E6F5MLA
zfb55H2dxaWluITUlJP06lxUjamsJk7tMp/nCKu1yNTf6tRG/rKKNM+zMdll7P+X
NMbYOi1GVXixsERXW+PCXRvNM8fMrjpjPwfxDRHDhZjf6R1XqmWGgdkphIlgId5t
YyXWlzGXMJMnnd9NcvqCvH1T7BSrebzLTzJO+ZkHUnzYKhN+egeYU0NPMq83YeYh
zoxhYyuekSEfUHoXsdU5Pjz5kRS74acq3iFCsX5YEiW/f3u3sV1vew6H9rMkp2XH
6gem+IqlKnf2hWCBVKSeYtHoLxqpHgxUmZK3crw0mYIeQl6h4ptw4ZsXnIfP9Kfy
Hi9u6ZYaDAUosLyyg2xrDM3K1JVT6th1TcRV/rdkUfYsbv8OhIM0mEMblNzDtZXc
EWYVegkuldIfJ0Czc+qEJlvtdEIzAy6kL65q0YGl5lk24ZERPR8mo7MsqIark3+y
N0lb8tWnOyHqOH6utI0ZJddbIYS8PaRO/Xe+l/mLlxiiYxq3IWWeeqpwrcmYrIkJ
P4GsZJZGCYRJwOA4qCKOhfJJhi6IqHh2ao+5ilvoUhakX16CQ/hlaZgNgP5pcdrK
fW41aF2KJ7JHTJIeYqYDytSCEbBduFBVcmHyjYf5nyQdphhVErMXImmmtZFAJPtw
8tS5A3Tzu33SLNfUCUgEo77uKuxuJfef0GbNLAOfooWLr1HFqiYvgV7UvBpS3a9t
cDiBOdpUW0H1zSbzR98EW1VCv41Sbx9B8bR/IDpupq1ZMVxNfsbnruKwMym+FrO5
odRzyA1gg3FB1P83rK5SBBvdJPj/hv7UZ0Rau6VSTtFc/1GwyOKQZCZr4y06wLEb
ZQa4tf3HF47BtDGWLiJXel/Wn5irA1gu2TpNB8AS/EsooJ7BFlJEGN+yXwkLX/45
NRwzt4yaRqF7GkwRI3wNtojbGa+UVHeYppKfFQWhzNUlS+OJPfcyQhULKAT6LKmm
RKxX2vqnoLnoDvESwcaoJ4pdlr8tPOSAPHFbHu8A1BNvpvpEI1sxB7vTwoL7AtXD
Y2XKne7fdKmr8QyH8ciXFeoV4Oavm6kVxnhJPPRPQhq9VeJVOO7nw0d21wsPTlTi
MNxpMw0Dq2KVhLQO7UkpSksEf2hfus250ziQFj5i++l32d4Osvgjv2wUWXyekhrx
fC/IfYXB6zTjpIP+7aEc/8GBVv7SPJ1LxItxNweY7lSaEgg4euxgYxSFcREdOeVv
2AehSBq6ykIkGBP+VkJSKJJcRgj7xz6Z1jDHiRAjc9R/CzER14kEtfm4vxdjTBcn
bdnqIJUbD10OjS6lwbajoc4306aky9WGPYIfFGa2gNz5p2hwU0NKmr5IRnaDmgMF
5JOy9J2AsjMDemqzoVrUlDONJcNB8qE22NT66efti6nhY77J1dRWloajEJJSQ0vX
+pugyLn2rYlvCXmaV7T2SfmZjKRbJQnniRet0XK70Suylmj+QjStfoTyO/wMimMC
aqwnpVY7epbGU8G864UXCHzthsm8OTpRTR1QNLHd0LibjQesHGEBuM4wSYO4dCgG
LOYgWh513FPfPRwzPtyDOF4PRaiq7LN2fZiUxWC72jBy5pu/0l84Ox2fonrB6cV3
Xtg2R4FHBvt6WIWOQuYN3qpPqo7mn+9oUwVuHKP8jqGntJ9VmajzGF9flkI2MuM1
cg0lNeBGKmBZuZV6MmQWAYZVhwj6bllLMDrcREXvFhnaQY6H4ngvx/KIv/+iYUQ2
doP8SVbr+l+KoJSqgS5BooaxNurIm2UKeT5IHIEgNscjC+4FTyXtT4nwY8AQuiXK
qcI1hQPRK2XAjKEZ8Yu5LkO96sO+Ny6N0GQ0Yj6U4cuEP3mf9ARJCA+1AAJiOqkn
jz2QPOyFSqjDH4Rzsx05NMQKpvHbi/JZkb9yWVL17ywTEUHDlTr6R9pniw5uzmhM
U+o2FWppIVXIMT7EyT6LUGSURTzfy+nrxU9O4qHYAqXu8zKa4U8aaDurRlAGBFeV
M8JRdCQOkd1+eXhIilosmL7O8KdfpzsxZXzT399O9jvfG44vDNzulB3Z1JvdP/Jc
IV092FycK0Iumx5TAZdj+AwrDqtftHK9UvHpctWu1dEOI/jFLKPWPSzd/fynFnCi
MziREZxBOou8mmOO6NUI+8iWhKsXY8hjmXWqDwsIDiN5CoOkwGUZcH+fcyA6NZ4L
XaVCrPWIHJEPQv/uvq/nkyhudYaApvJWT2QrdcTNDqdvjpOdTT/7rdEdmfkcyYrX
EL+o4LExpYF/khmoqHYBevtfpf+dAcZfm38vDKaRV/H2vywsU9nbBqCINd5Aen1Q
Ku3pEu9lDFM4/YMA61r3W7PbB9Jzyx7sU4p7tvfJJ6wj/2JVGlkq9dK9sYczCM+U
/gNhMj2DPVZ4JrbcOeO9xZ7JkGEZYgnx05AR9GwV5uWg8+oe3qx5HCVok3jbLUi6
1sF4uGOL8bXMCOdSWeEjtPl4AkNBJcsdoKhdNyA728Q2vnIkSWWBLYwKTJHgKBM2
8tnNtk+3sWzGxexEeMr3gGkiKXtlXlX5DRDxba/w04rNMqteVLMFbG3WicyFu5v7
Cw4ApQBCXqEuUGqUfeslC35z8I8GyjdJHw5qvblpUyCc0fMnK/n6yoHlmvHjYe7G
6daFlSYycObznKrvW/E2bEgjtVhDkkLEXJIqK+KgdYpJR11Yv/cGcJ7EjXIq9mdz
h8TBdClJD4xnl+4OhIEmT8K5pi5t/oTkPtdSw/ig/N5SC7VNUeHRbKitfYK/pQwy
vqUvun0719qlB+KDFNAlMGm/avdX1hPKgtKxOgBxJJrPOsuZ3N1k8UtWHOD7KVR6
xYPNS5KlEB9wT+Ed9Y1BGVMoFvPUrVhMqUAJNGuLedmVg4sTsBzy6nOKC9F58zLj
37JWQUmwdJXYb9cJDv5C2Sk4w7lskPfme0wPOenULmvzUxHxH5YDPTBYN4uTFcc7
23NFbQe5muGwkjTFRl0/lrEEhK2a/l3XEZJ1gqc+R4ZiuGmpG9zWKhTWiiqyKvtt
pnS7w8+GjiQ3HbePVr+Pl14AvR1tmn2ixhBVpMsKNJje+CtpEL2S2nS0nYaiwdPL
dXK0zIgNHg8T17AYJArejukNsHxjSwYB0LVko+Kv6KQ+6n6fa73x98HjvxJZv/y7
FUguSk0aBbVTJGEBHgXNiDfjFy9ku/KeESX5hEeIWj8MzYJbjgDrnqfHXwq02u6V
5aFmRQqs7XmttTYGmeTjTDpO6F3LXLMfTQi4kP6t7PPLvVCIzDk43Xjz/O2WGxNf
4HUMfkjWbkJ0XsYpsmptm8OL/Fv7bF7VVuiTkd2pGUUytGrQtOG+vZIwzsxwdSK7
ZivY2j/Cw+NGgdipQogFJMHot1Gu/Ivg/6CXm4pTrlmFeiPyQTwpLFc6uv04JeuI
p5S2CR2upiEMH9QaJPfP6iTdmr/xg0nWEw5tCJfbKxc5rLNngO7yiU0+TOOrVWZ+
pMPcdPueq5n3fITW9yT7Bp4gmC7/Gh5HA/HBkqHVc7SElWXMYdU+QztSXPhc43qx
FbbpA9ilWRCI3tIZAnGCr27HV/RXDeQAJ5uo5Yj1LsCWb6eY3Rn9/SeoXroGk3gd
xc8P7gFzccYS8xPYw9cRDGAicL5VZrZQ2BsSV3tDqCr3RNaoF07X3O9FN3Vnidnt
3Ylr6TaOSXvk/AuVNpmhFn3q4eBqB5PMlzTHoiKWgY2Cn6N6NLj6o9eOSZC8ttlz
fcw25b2gQYqvE1QN+iXaw6AFeE7CgeRdx8tfmK1FonKn/DAiZ7SYJTk7JEwHdPx9
KbLnIKo7YcCwLed7gp02tcKEBLqnTluA7D4Z6Zedco6wH/toJb6kFF1eZXoexNON
qEQ/0LSrAPjdBaB3u3aU+2pI5QblW7h557WkZMhZ8jEoJRv5tmR9/0wJfKMdmEmj
u1+6XrndAGLqijzvFiigDEQXKfYcH/DCpVXIpIgxfeBn1FtaxyXbo1b1jykGo4Xo
sB87n+DrFoknAGOfbNI9OSHgB2zEwIHd153h5VmevfMiBGznpL1Yv9tEJGG9aUpt
BgjDp/oGvFQ3TIIdBDC7pEJnC3eL5ia9wUbTF+AVaXTWUIE847tBT473TMJLnPoh
4KPWueN0NvorzJyl7FcXK5BNsN/XV3Jjf6HUHCIc1vxO+9pObHVTXUtCdBq+ovdJ
meTUW5atf56fKQBafmOudB7L+KnNHgZMA33RvRvrBxwRdPDWsGsF8WyO/tblrNqf
xB2AbpuJx/CPu3ASV4YK2WCLlfypsyOVAICcZoUrkYO/F8k/SiQeAT89iNPx4Nt6
qvq9yMTzpn/PlOgHPNpC/cFL/8JdIPE1PWGnSEneYSEIh0sqBgWk5snUHYUn4wSc
L4Y8Xycu9mKb+c+smCCju3x6jwr/UMtlTKRL6WWA9Bcu9fywaltQEp5acpOhl/aI
hLl3IQK7AKHgeLCXDxZ6AyOHnI0l1jeV1ua74zsCSgGlo2V2BkZMc1OHQUwpTeuc
jzbm4q/gH7iz0gG5CNzLeUmvKjAb5da18jicspCGFhm/VlYQD2N8D8T8V5ocwy7F
R+O2ptYm/j9JO/VoNkuPAGcv6R44zariGmf32nGDdZ1PXMjo6mwNJEaAFaqaU6LH
xtQMPX3fsexluycdTuNgwX0GQfF+j5aHDaGVlaAnrMq53u3nsMNSK0n9HCzL3cEA
OIgN5XxTuQUewJfEufi5on1TqkwcSJa5LJfSn9AS25Vwtybubc5b7jSOAXoBdTkc
HrjT790NgxQoTDSHURnaJ5MI0JWsNMfdn9Hw9wq9cy2lURt8A+IYIxU6W8BvOojP
9pXplQwbYYRqcDXUQLISk9w2XG+DGaXK/CbgnR9I127ubiXMoOGTgWMzSNw8pmh7
2+s5085QUaVZ6gCD4Ae9Dvf0ILpXV8iKGLJesmVGrBa3/ugdhVeAOCZgslCsAXKM
g5XVN5M4l900QL3KCQh+q7PrIXLEwvz52GG1xevAUw0gUp2kUrVM/fg1rcmZEZ4v
/e7HoNAK4cEU3/esEqcPq7qETCj3T8QCv+lgtRL+CrtLswj0mte+fx71HJoHXJpH
GaCzDU/xlmxA1zl3InNhzhI+ibn3RLXqOCSAmWrmBoXcIQCtN9Xen20l12qHPMPv
plAENBeyG4f+pMlRzI7NG5lVYIBA85lsWRUGg8CgEtfp4gvKMmjc26wvrK4U+MZw
c9JlI1pkcv3NM1cIVWuaIJkY6/3drHOhtcPeVn3dL3N8KtCQV+XcJD0szUT4KtHD
qXl4tc2ztbE5Rb7ZfjOLcmEV94UBf3RSnPWWuiDKM65LJvrgg1m7FY33s0bHmrLR
x+t/aIPvqiISUoyY+3UdqYqUzq6X5z7pIGGxhT5W5wJi3nIFinzWWXzP4xqzpLnU
NPeYvwPwVBPI9tKGX2vH29kCYOcNVNUgBLgCqPqmi9Mh9kzCV+kvnu4jT0U6z3Qr
bcUXCQATcwc5gEjIW5DOZoshYKwxMrgaBz86+0VJ6PP6/zRLHDt+ogLMRu6jnWUI
a7a0vBfjprUWfIlbyA8d3doBOuKrO04s94RMq4poCebYnKJoPZ4j7EhBGbXwaoeT
NO0uH4h4d1mRS4Vc2Vc01LbpjsjaHlb2czfWrYS05TjgTQkhnwpZSatQpxpg0nhB
bNzthqgZrjn0FOOjvpqwp5nlTwvoI/mvOizudynJDliFQxOm+EIUk54SN6x1Pb3X
hVj6M7w1Cfhwlo1sHCGV8zZciNvp7Tdn9gaxLBMh3VXZ5g9UmlbjHSrPNHmHnQVc
rOofVtQ8gAIZZYdgfotBUh6jSPijG9I4ZNks/YzetOvhAPT8anOPH8Vqurzfy3Ei
35lI0+X8Y+L8cXcGBwZeTpWBQv5FRzZbm1d1AUsFcrAnQQVT2fkjmkiSBkPLWvXa
0ry7zY1oiOH4grVy+HJy4kRQEACL2agQKvTTCEbalWCJG8DumLPt4HgOZP3UQrxo
ODhC/2FsutnM6R8tv/cKy9iBHmZQaToAbGvmCdB3LCsG9wnbcsAaGZIkRmrKBZs3
NczU/ClrXqosibeDRt0fC26/WMOHHGekrvqTgV6tGLghv4VXateqdYTPcYJhkQYS
oBsVX4u0lfJszKFnR3ycCGCNFjv+rtpvjFSARWljbsr7LFw49YByjETNigKioo7Y
5I7IoXfV3POAty7EOJHoZ3nE5pNGYwQ0QLFfMQ03O5Is0wkiE20Ap3Z53nDHrGS5
VuzyfOpKqTkDsdAuzzNpCXN8vxYMow3QCu4zz/9m/U0aXHBzdUqEZOUGpIjhFMAw
ccuCHkHuz5bnpOaldzQe9sZagbBl6mN0dj4sFe7/HaIPOvCTSLsKiRzZlngi39dq
Veif6hTIgvqF/0XgItJ/6XNSqifcj8jrurpBp/J23cMM3AVwU3WXguzO28DldKTK
LIkLyvfNgueKyvIN1NdHvx2jRahRV9A/GD8fuqNciVhUxlkUjMMByvXHXn9HognV
Wur6LoZAVTRH1eYZ5hIMpwvXHOm2QwcmwwiLBxsPFS4wRcAY1u9W4mWWllp7+MhA
UqdghB1xypOtAGDt5orj86RbfU5Z1pqFxejSysRTV2QfxrAqmrUSY7M7VGnRE3ja
ZzzChuBeAsxfidnJJESYtDn5e2CQh8l7wZqjLJSXIQ8F0/OeVmPmGupFxbTq4LwY
UaR8TOYvcRlFIhoisUmuOXMchd4/9dl16g29E9fzXyWwdnB9xhjXk4vOfAhSyV//
AO08A9ijpbUwAxgjs3aVt3+6oDsu1Dl/WcyOR7vLX7cX5A/wa+gb1lFoYOoICwpg
s4Zoz4Uc91EjfFH5m2UZgvHYBHxJI61sXvy16fiME26lYfey3p2OMm/8LOBzt98J
ga5RBPHQj+EYJtfZIIHGTrswqpKht9uHyvn+Ziy7nNIJkksxn1eEvtSCpqiocTbj
BxTgRS+YGQcIMPdU7LJ6swt2vxamh0yuGgah3aVRd01a6oZknMs6noYHLvt4qKn5
On7z/5FGusbjMDFZd+GihpeiHdcDdYRd1jxwNkf5aV+Kng9ObhE94zYAb7d/5aE8
wAvPgl1fyXIcgoInRyoGfj54TBGBiOaLKqZ+QfNvYzBv7Gfn2+YoLJvz949g65ok
3w0lfyhMBxQeQmUc+dkbrpa/d8FcuCNMW78eydLzyOZhns1ctt7NOtzRVyKMKPHM
4dtUIgKKkvNVIEtWsgBgHBk36cT3pcfGXw8HsjPUttPrX0HvvD3nvxq8XahxF96I
E6NJjFxhXO9llY/Dpfopr8v2JBg8246hSM4pEfFEK+b0xGu5CIW6UNdlsOiTDrtH
Az/bJY4uuLy2I3Ah/4DNkaoFgdM3OXqNCqlgT69X//jQXbTAgAO+hQlENNRYtj4V
3RULFqlVon/uxd2siCtvDA59s8I/zL3tv5Wf8qqVb9PDOVueNK+kkbQ2yA8FmlyP
VIdL5WhZNkwpdbDDw4UMmSlrR37eY220x+qLu3rZZFHXuWBeEN5aUZdhuGrnNLfU
XAqM5Xxkw8rNaXHKls5nP5IHDQ8he01P8j9cvu2r5hg4usQJUuG7Jm1k4Af0NiW+
77V1l1bIVJ1EUjACJ1jRiOB9815OYJ87xpUQhJUpZdxsK/fudhRoEAvCetKnT4Gy
eSgjAwoA9oC6QpBspCU4XstFHTnVrHnIxkD8dkgA0B1l+RvctmwKOKqESK6q/v5d
UbkcziepVIvWSdXUkVJBJ8QGoTFJVlqtoGckHzgpWQOuqhPZ5Bq7he/vV3FykZY1
KqhRcc49sNBfg/9hKGnQku/lVJuP8Bf/WzoXkMNeY0GO+8Rz0R3NP54OZmonvcrv
Pmpl7JK15WtOxGHitHRTZzQxN5p2ALpn2U2Xnku5OehVhkVaeG9e5r3T9Yg6ckJD
M0FhGCE3srZoq3r1G4AhUX82MNppGRTJISS2//c0ouT2qvg6ZcbatH1wteysuYFn
8NGQZl/sSaORQdwq+qKc4iHW/UKW78oFxlRzQQI7cZDoEgLASa+ogp1dQ0fRduyN
2qUVzpAObJSkZJlKy2b3vaIoHsm/ku8ZWNtonnH/H+nvM8hYVfVJkvQepCKwMpfH
dR7cKyCOfqigO96e9X8dT9ZyfYXZ/ot8X23nUAwUcGEED0wCxNQ14urcwGHJyHMT
+h9aln9FtXVkwxr2SoeUHGhVdFJwBm3Rvy2peD6Xjr80Cr/P5HZwlLCQcZfOSKym
Ep8x4RjIoao//VqUJSmqC1h2lFgUVL6RY/AWhWxhSwwldIhzVVDuGHDGwp5IR0OH
wMwgHSUaEj/4SbfR+SYbOJ2zoCgwjny3ZWuWAgQ09eqMtUh6tminG+ZWGJg99fPX
iiu90+u/JKjEz9rax+Gt0LuA1cmnd35NgYqP/sMBj1uQMlzGd8P2nE1XYe1ypP2p
Ag8h75CqTG/JrBiYEv/YLuvV+wIMUBwQ0+n1rvuWqTQIXkhfB9b6SSUhRij1tO5B
5OOebZeTWJzw4S1jJOGloVxr64+wLAhKL5ruVB7QISImdPPoojkWhPOBg6JiqHTF
YZ8Jp84igzK/SKGmwjAVH6vBDVGqNJL1XaL87P1Z/51/d1nOWmINzkFbZwednRYM
ncuwYV2WBFu2h+DWidSW1b258Z2JcDjhkG6uJB/LhKZ+5CPFD8Ubw9TP/AhWFCe8
6dWsYTJUCq5hIAKEr0zB4g9vP3SAbl6zpQisonpQbHrYhnS57tHZrm6TZt7e562v
cykpTSMs6i7fgQfjR7LJkSwNntYHdpdaCHNZ3fNUZBdlJDF/eC3e2WuRzIa+yAAO
DuXiodknYYPVcqEzF/P8+IW+qeqoLpuAb/e3PfcxUSA5JNxK4pf1IYoIpV6QD8mt
USXzmsdyv60YOjCQari24+LLaKqsjin5glnnpZX47LzslmUTsuXig+JnIHPpeEvj
xiOrwJV/HCk31UzFpGp3h4JoS7Zx5/10Q7Mdas9BnBPvm8kwInuCpN6Qskr0hX9N
XVs3xq0wc1Y78TVSAXb/UqRx/B/2Pdr1NMXivWnlQKq7MQUVSGNKAJ03xBWjnrgW
nXmVZv+InFLT6jbcVFqtOzsBBn3jXsIVN/CfaXA6MXUWMhsVKHkIy3Ce6RZWZuZa
d7gbNqXvv59iXNBFoGxbAKA55afthxe9A4bh+sMw04r7N9UVQb5CJ1TC8HXO7gOm
FRDJw9fB9dPzLtJBjK93Rg==
`pragma protect end_protected
