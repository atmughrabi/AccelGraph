��/  �nה�-����^���@f��	�-�GKQ/*Ѽ�Q�*�
���� �bY6��M�$N���A��(�<�s�Z��o��� 7���g�)Б��U��;�LW�ͪ"�K4�y�~�� ?��T��,�=�"�b���~;��Gk��gS�&��^�Cȭڂ���Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9���w0��m�KYpp,"��\�j�\��:����Z�X�?v�}]v#���n��RJ���{�7Y?«X�[�e���N�b�6t�NJc���`���t�[��[�*�eM�=�G9�y����p�]
�N�	����`���ú9��EL��rQC]r#eW�`j<3~�~���ARh�0���B��>��,�t�0IĒ�yy�x6�'��M��H)(�b$� �\�x]�@���^y�8��h����?<��tB��~�/[�2�Fϰ�ਊ���c�$��+4�ϫ_�H��b!�j7o���ZN�ܲb{0cS��$���ر<ܛrP����5@�4~i�����j���`+U�}��y�,`~�g��_(d���6r9�mi�b�������`R�GΥ�sAۍF�F�(�����\˂�zF4�IU)������w/?�ې���$�=L�s��z}��Ն<9��1t�ܷM�o��8�Yq8��|5
!Q(��-�S�� >�>l~j�T)4���d�Y�O��rDi�|r�	G�<�������\&M��tۅ<�v�ܯ�u�Ta6j�/�� ��e����W,��JAX3��GY�t.����Đ:3�v�ݮ�?w� 5������t<-b
"�ݴ1�q�VM�B�=����I�C������&��y��� �hճ�1Rc�����Uf�:L�Y%ب��Y1�f��TM #*�>��-"���KJX