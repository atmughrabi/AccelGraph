// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GBnBNfvFmebGoWxHEVgYoAfbiByBhvSoG5OqheZEVKS7ngOfh4uHh4WqBkcVWjok
xcjDwuLYJ6ijqnV0hSqlwZAy79fbLgtrTYxTOq+8xyWARKyZByaGB9aJhrXFk0sx
SwEvjRvyboI5eomJeyGuPLeSAEYcsVl2hUq12VSbqhk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25408)
97A3XLnY831rJKlP21RukjDXWlDIMwNwMPZN9C9T1Z2j1JOsgqPR8BNS50zOIFK0
suygc4FSVUQ23C8WbzmamnamgGZJNF7ah/0JcQtRBwyLUkSq+WMv2iZGpVelvafp
KxMidwYJWFj+K5z+ZdvYrUFF01lB//qiwgt+XXWzE8n1+6W5nrgDPpAq5oUKr4aU
EfxvlQj92triU2BVQ2u4vnLxeWqJm1eTn4+Az7+3ZgTo5Dug4nuZZtSijb5kYvYF
nweVZaRDcYq/snSEAP6eyCKsKwf/Wh/xBNhPN5wDlcweodVXP8FJZF35rG1bi8d9
BO1rNS7xSDoKifnLGXa6uqNh8qopLO9LfrtUDS1AyFXlBx5yh6xaR7hyQccxV0ST
rCuJfRYA49kWCYZAB5VR4Of8LaNeS6OPiy/hfidZpAEUDEewyrOxkhkCWVop74w6
ZZ1+hQlZwi8TiCxKgQDhvDN9rhXveAB45caDO/hxLRb71YyUXp02r8iIrGpkYuLP
Ro9CnNebY0+TrXSGqrQbLcMAEmJ9Hxq+Wus53QDWnh/xGIETx+UmYLpULYYnIoxY
DEQY9Fk391+x4l75S7YDweRxAl2qSo4FDGw4A6GojVPzXlyaXpiler5G1dqEng6q
kx5mRfdnmTCFi/MCTNI+9FrNaRubRKHnpgg09aKkT9Mp7dnqPAwGQgX4Gq1/iJJ0
Zqgza11tkC6GujHy1a9YKtSfirLDA+KBGlEzSXsXmbQluuV5zmxpSFymOJOZSzKC
StArYTbTM6V/7LiJBhS8hgsHiCpVh7C9V8XWMs+Vm7vhratxF/CpQ0/XxELrXFYH
6Hbi0lwBwlUb7PJ6Nnd+M07npXEpqIuOUIng6SAc8+5ZvksNMXWuh13KZeUgntQh
zjyyLj7VchyCCmlk7FB6+Vq7Jw1cI7ZDo3CnYdkf1n7t8Ubg150V76KrJgFqVdmX
eWoFOXgp++d1BY1R0GkXONkGhgFFz/mz2Al9O4rEbxhRyOHkHUFJ2XL2lzQRJ/qb
eo1iFw43iGqHssAPx0XCvx3Z8aEwEVwhe8H/3pfgWTp+mNuDthxpm4K+QtUl+GV0
kqYy/FTKZfHagJJy+DM3qM7fcjvRSX4+ag3uoE/jvY7bzuycqJSUM/sR97gcyeCX
gJ2hIAEeiPcD5boK2ra/LRW1l4vzme+L1rqtnWuxxk96iGFC72x1fv62ZPzT56IA
1UzxINaaDwx1ZVNgtTRm9YJAveyjBed4K5Vkso+Y4j/+ccQz8O6xrjihZo6OVVVj
iBFGO4T3K0vquhFgzx9oeaVIXcUaxF0ibmngcPFghH7JKMuHLKaes2dHJuPLbemM
zavK1jOqDCYK22zdKxgNpFa9pUsF58Dk1p72KbgHu9MT3WfhBi0ATMspFeI2AM6G
CcewXnD/yxu2ey5ZhEULLm1g1FMVn8X4hYhXuX8U85XPRvXKxw+yg4ODFYcmrPC1
RYYBviM+gOSBH/l52KfU0XQ0g7ui1gsCDmw1P0YZw0zlvWwZDX38Q4dciAfXf4Q2
icVE7p9LdeKyVpk2eT4u0JBcVBJq1z4+avqJN52I6ZTpeIKRrAA3fe0kyJaHZ9Aq
BuFe5exJxJRyGuUQMQvML4fE4RVRGf0JP06HVJLzeAqAHfkL5AE50OgfBmNa7LO9
w9qzI3+SVH0tStyHjt0doudZ11IR6Ds3T2r73CiAKMjhIZmKiSctGtyRXFI5j33I
sl3eqdqdU7KkmD/pKw6Yq2deQwj5lpBgXLZjDRudlXf0mHnM/6tWbjfGFOsn0ck6
UlRxIWpYlYaK8apojW2M6ycwpIUpM/BzCYZn0Jl+NFNqiN3Iz/hRCyjOJECjop3W
Q+Arxp1V393evkjY9COM3tzXxV3Sdd7acTYhtSJPl7JghsmeBtaF4+6CARK7epV3
Zocj0Ezpc0YuyLGuEF1QYIOZsn+fuyWeIeG6YsOwEkS9sGlet4kuV27/+AmO2SeQ
z/qioF92posNzTu1ogfml4BYRPlvO9FTLvA7oWhKPd9bxpG/Dp/TZM2adWGz3xQt
N8nlRzTFK0nvJ0qaA8FMPN2paxYczN03YNFiZ0KoieJ3bmwqWr1CnSGww77KVriN
Rjm0vjZzD1AErNiWCK6g6PZ6ZEqZ/Gs1IgVWg0lQ7f93nOMTjR6R278RdBbA8umx
qCSbDkHKksPllqFNQzBP+SRcaQOdHE28shfPNOpiPXa7qi1x0o2rFbOO1x+nuJT7
ScoPabkWwwh+2N1wKEfuqw33eN6skPzONDBsds9HbLv3V4dL8/CqJY4M6VSNxjIo
LP6Jf2/WjkwIZFb/agAJQ1ww8N3M+8kichYZeWrAyfNNJWc6zaXZrKyCADcRfnX8
URd7qep+j3ZgM1c5R/Ofnlxd4QrgktHUb6a8u0J52nzBvotagVYXyhWjkmWaQKmn
49wOCIZdppE1JUn8B9+YJW2zNixHjoc2X9lpzQkAk0l+TWZB7JnLj8Xn7cxRWNmX
pnvQM/oN+5aPrjFbvGmhjJ/Mxs7IYE0Wu8S7556s8INCVv5HHRR+Qs5qDaASWza5
SqO6+yM0WuY1j+zHAplSJrg4nYKYbCwB53pSRw3lW0ySVctKTCzWob6sDVXBe0q/
9nGht+0MtG1APCIR0/xqBy8GZHCu5zluGsAPCEdO/lRtHuwdMMhoWLSSkDO07qrK
q6C+L7DywFXrxCUwO0/phHE7se0hoQ9wRrSYRhYmRYIL+FdLwWObG2QJHa8P+BQ9
avqjTtizlOEbhTZEUEzk85QUKZHfjhJd63b919d0tY+SbYgNhPLOB5nkYn1Fe1KW
Iu3oxZPwbDG5WFMlHHHxVbt8Nh7Y4lzXIB8SLJdf0HOYoqCyoNnv5VMrA/zltnEr
8jWt1ufl7bsxpj3Gv4zAVAGXzxJESVYKrqqxqGCsemXUsGRX6leRKy8f4kog3MG6
TZ/sNxZYdJpADFxXpx20KaryI/FEVIJ2PyLbdXEbZybpwlput+NnOr+9Z2M3I9K+
ejbzS5Whn38CLpsakKEpXU5rqFN/04gi6zkRUOGY38Z52yoJtLtilnvP3BjJjlUR
YsNX9ik4l9GNniUKXmbGz9058XG6OlylhwjziYqmVkkLwmALvYQTnrQHp/KIeFHx
KceeWiU/ZaxWCalWjGhlsiD42VtJJiUhKH/LgLf/E+ZhiZE5L03a0fMzG0PWRZRU
2fXuwPUY0RnXc2wetXVvIkp3cypNmBC5w03y/MMBu4DQjI/g4eYPsvQo+T8zOvld
fxzUO7WFagpP0Dquei8O0/FpgBmDjSEKYn0qHxaaj5XviDi2+GAmW1Y61LCz/4LT
Qq5pW1K4kb89L5mbAfgID5WqxCPA9uJbuEosbMkOil5aNz/8vZp+mdpZG91hqo+y
LyDIvgyuE7p2WJVuYhZT+GUT3ELVJqIwM9mnwyyPFzknEp2f6TUKfm8FiPepPTCV
cvAjkYLQI7VJ324P05Vy5YwoRwio/kC395dkW8xsevEI7Ko0D2Czg/nc2w3Rp1hG
WvnT9QGRrh1HpUmiGVCtr++qeK0WocBjWz/PQL/WKMFr1uc3FiGaqmYRu1SmIcAg
/lXBlmEeat6lzcY0AlBkAVeUhvjusJokiLYNTrWW2GW1LuZZqroLb8H7uSXHaMXk
m3T7G8gUIvj63DlRRTYP32ZJxQNYMHn2yWt812tfgcfy0NLo9NKWZQNavjjkAI/C
cwKa3vmKWa95RjyD9M+LTcA8UqWS7eshF1AMfLJAsmq3L0o2l+Tk7c12vM2SiPJt
SiyvQioWSENz9GxDjzMk8ObDbmU4vy0rrxnL3lEJT66NaV52LwVNClO5FL9RKQRY
I6Cg9G82AVfLQJy5wnVir0ycXRrwGRGQG+k76XKiKk0y1GE8IBrGao+h3XxFJ1u6
JyMX5lyxuo/hOCOpbGBGzAf0S1OkJIMzRoo9uCjMzz5Uv4OXrA4WTBJgjWapxXyP
zD+Td/kzGGOkxLcEfj5r9uxQ16+m+yigl7DHUzgmMWes6C8SAgcCr6Y+X8uEndJl
oV/XWt/IOmF9F20mjA62aCfosIVAyZf+hltIG8HbVlzL37r9pLTUVh49yFJeSjIL
DiPyEUQJ8UPfXXg788SoLn5lEaBI5rxJiLVpCjf/hrKWBGB+kZbnNzPrgEMFDFEl
0pT2W720ybf0rDtCYco5/fZ2izD7Hqa0haAne/rIVO4/0P+hkfmCtin/dvVklnoJ
8BfRDoNlcY6/dFDp71sMrJig0hBfREDsZGPYt08iYDzzUgHqGZgV5Y0pJOQe9pYY
u5L4nmE3scYlxVJGJXV0GuNAG82KY3DaEqhHv66XB86a6xyzsdwtNE1uSui5JnfR
A8vCG3oxBQCALtXzHd+DoL72luXJehbrvX0Se2dV/nNvDgKiz5+a4h3lLuHc1Pj/
sa9W9gaCCVlNFMyfV6ISxB5rB4v0L3zvyJ1c/KeFUB1DrZ9oJauuqWs6aSD8ZPn8
mkiZt4MgxnZ33iTXqu2IsKtk/qDXFfrykIwrMwg1yMTsCrcnzBXqOC0wWrFEFQM4
97f4xKZTAaJMxQ9wmLsLYWXr2g7G3WFHu8TvkdLwq2wOxbyOCwfZRO4pR2eyNHlz
mF+PDqtz7JGttj1x9Alk/HqB94oLkrGDYPHhBNESl8EU35s9cNEyph687yVRIeu+
xjMqtSCG+ELQyhZzBdJhFxb7P79AImMZ0qzs/3z+qMJz8epDfm1sFGTiCvdugN8j
2nPsp20RqcDdBxXERYCu2WnpjfkhCQPfL0bMMX9CsplqFHQtJUohCYyHQohg1uSS
h+D5BPFUWBkXx4SLeiHPJVCryW5IpBjE6cg0aJ6MaGg7pq9agSFEyPb2kcMJUkeI
8iCxliPU1Z9S3Ncex9Iwc6KT5mz9Be+J2N9Zh3t5nBARSAkeHnPeWXGJpGazPzGE
rUM502VDmWnloj7nUCq7i/gCRVf5tGG3crU0HptbSO2E6hUgtl7f0ph04oB+wnbc
6JaJ0KAS34i5S99xTCQEd1eP+0VyFmiTzMcHcpuKnUgP73X3wozrB762qHliqx63
N2cwCjrDS9jmLK1AS2dDDZjNZz2wJ+LjCgHVRjucymyPfREl5Zn1jKvhtFUW1ine
pgIsepv3jjuxBEOFcnn8ykWO/q0lblPyIa/UxdAZeFDlHhqiZYjYWtrgghSaAKzv
EPBFM9+ZSRwt7XifYrFstnJnTZ9ii9JdRxWgfdkSegjuW9CHT87vEoUaOFnBmkV2
ROqXpUOxM2YUwl41PKJyF9TsQXJrzdgeU59Y0H0KLGzEjadiFyzhprCqECs6LrVa
860JmrFNDz4nGrB7QYE+NWdYhpQOXh+6EoI1EvtVVK0PYwWcH5y8TP4DFTz6tQRG
MPTEsLTugNw/CalO3qgZv/zjEn3ajaVpUENkS3JHehH8TVCJe03Nb5hcxO+GjiJF
a80Ve3q5XKqAcKipTa21CrrjOBhxnvNr4+TxDy/t83xTn5vxxIojBxswBzkL9V5j
JhiCi4Pmv5iShR/t5/RtPGi6JxlyHtWhQQo7phwSaePTm0FX4rDPTswibE6F14aK
Na3XpINA+PiTUzbdZPB4sR8R0JSgxjxxaa6PQag2+xACvZ7rkOPbBnQsL07ltwFn
/zo/EJLK1AbljuzofZRb8qYjtxZAo8nVPBps4wIB7ARJHw0QU4JKUXkIGlxGz2KP
KXBD03QhViErggbbevH4PPZ0KWB56x5vp3r0tY883sljqK0U+1PW8rYFEVfZyBtU
wHrv7rTgX7ULnwAPrajv3iubLr9rVm+r/J/aZzKu7uAfIsAcGvWxM8G5zZPc07/Z
WENV+b8C/OfYxnhUemn39zJV3USLgllUN7qAMpXPj8V6mM//JJXcggAgPHu77zxA
ZuFV+4ztWb9O5MnbOiOIjzQpv5JKLLThurqUN7r3hX96zExqEPQHa/XgmXWlNN6+
cA7111toeVwkj2mS5dQ8lYOPu+SVF8gGYFR6ILQCaiivLR48qgCFylnSiAPQJpZF
LNnxgQzeMKZEWc7x++UpZeQklja+XQsh1QvX/GK0JTuTy9nD/3gP3/2zf/3HzLNI
k1Q6aSUHJtt9KfVeVusODUOQ/cairprp1tJK2FbFl9cLagQRGdwnPCvHQEsqg2M6
cqoMEEZj7pBO6lcWrn8EJWBTvCj29xVu7ZAjDP3fFPjt/i6RZiETrSsKG+FwOYkM
41gmZhm0umiHYobX4f72EoaktUBD+fMz6Y1qwTTHOlXPFZ4K8Z6D7LLPxcOSTiPn
hUsWTbh10fMxBwIrZV3biR16hv+iZgShyGmadeDZOlAdBJ1chIo0WhPjSUSE+zHT
W73ubNB25665ddOJh4PTXZSCPsA3Q/FREX/88IVdXCMYJE08xsMuhsKBNzICmpbq
tAQ1cdZ5QJh8Dty8pQVN++eWknfL9jRqGrlEsPlE5Tmsvc3wnzTV3WQWmVDywnb1
UnLy29yVvsQeeqWjWrkO5Eesp/HARy4KWbJCowZdKetRi1OwWrzkDZ3SNJm0lcIF
Vrn5edQGOrLcnnr0ojSXaqz+skJP42s0bOgr76GUOPfWUKCBEnGXhGvvDiZYjEwM
DmYYtZaRCnb0+twO+6pzgRb5c9I2iX6Gn1vERfD+HwR+jBN1cMingv0IsIXyjrr2
uNMCsB9PK6nAxNMIQnN/0++vP1H6ksVl9UGcuLQZuycvILCBy+rKkoTDjVu7ZsiS
Nz4Sawz0anhC2HuJrNfL204HkuMMXS8r9usIjKk03yUfcFMGSM78OTPF3/+V55Kb
HOOgpBzszoLR8+8cii+SpylhWc/H5zyX6uLj9Ugqy5HukvoN1T+45UVUbabwapE7
VVe7jR3T1z+s6saJvxLW0Nvlu/MyeghyBMbZP34eP5YtZBLb1UkO9VYxibGIngM7
zY9JAInratl9T/y1z0mwODGemV6PX3CTiivIQ6k1GMEAXSBA+j849vOVCiTdpHS2
+8P+fzlnQ6PUfEUoSYCCOLQ3zXVTRuMhgffcJEUJFK/UDW7HriihMz/VUK28vRCO
6s0CN/0qweTVkSfwX97Ud/gFpBt+N6g22WrmCuUsL/uI6HJurRB2MNa6gda4M81i
0xhysnNtMstRvqK1zTxH+TglBd07Xz8kU9L/upFNER6k4YfMrvo09W/is5mzmpJF
TctG1JyWDOevT9Hot4rSj9Jkf0et9VAtfg0cL+4RNSv3sNj7a+w8YwcC/tLPJ/n0
vBYHB29Fc2Z9SMnbfhre+OX1ryeYAgPgy7RrMDbaK3o+S2WYr2D69DzGrb5ezC49
29x7qiLfGqj1nZRFg3whtLhJuaZvNc138M87YIGeCmXL2AQTRyqq5yd3Eqsji9Rf
vKJs02ALPe2RuCw314S3N+LitQAlVSiTTi9cJ4ByyOWUurBWXrv+X07IuBcSmMGd
ar6auoUxI5Gy+6s4SwV1oLH8gDH8AALUOn/9ensSMbP2Y4p1Mh6N4AEJWFG5F7RK
+M1vY703n3kmqQ9XoH7HwovCEwlrUO/4xry8Ce3N8CTwSe3H8p8NCWpXgNlatwRf
P21GRpksKn3+o91oaTqrR21dHMQrW6LQPVUEXrHyFxK9wcnLjKHt0AXDp5o5LPs0
851kEEdEucpZuSohuotmLKAouruywqN37geTpayDrxV/1g55HKeROQXJGb2E3qdy
vK+OMZkFX9S4P0aWg0sQp+fav6KSI7aN6h1QyaU1hpsIHz6/2Y8majgB5NgOs5s7
wtYtwUopNQXavQgivC/GSaJKfnuj29NjhDQRNVLfuvvJ0Ft1eHaEeJ0u3LUBy4Ge
oJgj+ofV1YCbvKcUm39lLiIMnZ5uRjTo1XHkVMViweZy4P9Mr2ihUqRz+ITuV/4F
YcpaQfD9kI5GKwXEx6+rsQeZHyYxnhz/oK/0tNSxN2Zi+qFvaWRDbUx02VYyH4Bt
20itTPZ+ybTHSw/pCmzCFMV5Qrk2M5jPfEAI0AlVSZPCEmT4r41HahR7JPNBMP3L
snUrl0CQEdueoNI6OlAY3c/KHaaBTJT6J9MZZckl2kuIZ+cg0CIhzfcbBOhRdnSz
mipac4hgnwlnquTA0l/gpAdlyhSw+vvFO6ARgqf2+uTxgjC7dL4e9LdLgVwzhblF
Qj7gcKW6ptTDGA7zbwN1vkxB8ab4rwmIrUF10emXiXsCi9F407eHoebwUnSebueS
h3fACw/eIrI99v3D5mAH6l3/f9hjY8QDTfC1sJi904jURueG9KJgYLqXJCeGF4Yq
+4SQEpElN0c76E2Jvtl5lhZbK2wsVS3MVznyryPqMVqrcrIH5bqBGYppHQ29OY/k
MAxIxnx/bTLxN+MV8mkwHnVodSfZWqYSQX6P+V579+4CQTpcxBuF8hS3beVLpXI2
V554SZnl2wu6Z2tZ2Vu7EY0MjOLjz+AfuCcxyZW6Fj6UE3J68gjKqe6s84RYDa9o
O+MIOQF2MY2J+j3MoDLHq66d6BxiQSek8R43uDkQTwoUxe+OooAL/SmZY8LsJtDM
F09quDBrOwMB656DISYQVANIs/cULuSKCx+6O2Jb5GCTNbspS/CfCi8XSsJFEAlh
ymDe8WF2maw5IPiOf4zC7wv41gYsag27j/y33J76X6Ln84oE8Tig7AUWceNm9gF0
NtyzhBygUe2TeUqVSqIVYzvhi6uPP3zzoT6nF6KRMGsrr5e6t8csua1eujqLxGkq
JuA7k4t2gSCHjXVJCAAKI2h9CcDiqXlWLtATFICNe18QStCL4i+LqNjimt0wVqHv
xGOgt7v2We6lW3x6yR4jYSsmFsbd5KXScJM0nsTrMkg31s2y9yvR8MGqHs0TrPYX
umvAuCZ+2O7nA4Fb7S3KT+wK5XLFBoxOzqc4Px2pHZDvOf4GGpT/SNzCrrVG3LVa
XS9DG6Qj0SMDAX2bbH7MsOOW3QG5UycL/YrqUxYp1XzYTo7NHrpTNUwvImGXTlKr
CReaRECTyFw9omDZ9At4+7/oFuXkfw9v1SdB3orbI+SGMaZCfZCAZYKrQhrJc59h
jiJ+cT2wa/j0DW6moFQa916lpijxlLFrJTrqbuG0HpkSM3BLIJx9sHLzp84L2uRk
bUTEum2FyKq0rm2EIOhJj2eAAy8kwARKLA1z1FEJ+B5+AoSXCEWiuL2K1dUGqh7Y
7Mw4RlkFN17/26xmyH3JxVi/nJxsqpUzVDCtzBrtX/5WiragJFaYnluKFeXV0m8e
2cASW8eHC6J+jUaLGYgJaGFWGQdpbP+/NijmwYy51HXhR904nabfLHRWg+OeDNyX
SiZS+SGXQggMuaozC3+GozXEbtZv97rPnwnYeqwPVRZFx3y3Cra+gZMCH78iDMLF
Oc/4szWhxxJWGkBCHa+OYrbGdNJtlKg3D3MylLb8YoeUfrky54gmzvkG1WL14z+0
jIQVvWDZpBO0iunmP8hdGCgwdCHTxg+XEcBwd7dDoYIbEvKN1ekO7iE7znIGf3xm
brTFkzWqmCuLrtbw4wphm972QkJEpTuu2NazoRshr4ZHh2szuVmwntHbgxifl646
M4IfR4FFD62qrcmjBv7NOeTZAylcMJ4SIv/QG0DX6Y25RHh6gDwgrPCIAqCFxdyF
hGWtDVTl0SoESfouIAvfGBMnjCi9YRbz5fTWVzogGUV/K40KSu6IATjRGTfUCCuy
A+DogUUEU4jc0oOI+ha9HxNPv+Qg4Yo7As5g6WBImXOCd9NDBJ6LX3UAK3PG/Zjd
PtgF384gX5cc47p6wcXcfKxXBD07IdJG+cbS5uy4sZDzlUAfcrGlylLR2NNVFdg9
JhlhfYMWQximec9wHvlpow0884Lkk0U3onx/px8zLnoHHX5ZEb1LzYNHbbEOIHIN
xZzIJG1i96ZbJHMgHfKHOYmEkUDquUMeSj08uVJ8Nord/3xts+AUMuJ2UBojGQ0s
08uhFO0NLHEsBQu6MU7FXrFalxl1m5jxwC5Yc2+T7fGeE6AIkQC4UxQRCsn6IlOT
LggQhPPYQsxWSoyBI1ps6YxY+DnW0204uLAInCe0Qf/7XUVFmJiXoIKIa4NUuI12
ZU98XV2xdB+y1qYTaO93Uzl2uP+5Q6ASjVf4ORyjXCYrb4BKVSe0kD/aHPb62cpT
6MBRdmt3trLX7sgAauF00aAd7QK5onlc3lMVGyMiJwsAWWKvwBHsyDBHNfYWUrdB
VsBX0tpNj7vfIYFBPGuRDBba4qsq4PN/9RSJjubVd376yTwSkv/pTwXjAlYLKJIP
0MMMu2/U1bvtr8V3shwi+IfkMGmcrHyO9kUNrkL6M1FVQcIRbutOEr+/n6wGThsH
+N8FnW3RRJi3Djk6Gb0h6jFRDesHiDElQQFUPXjyM2Tz8psbKXeXvrAZQpyE1wkb
LQkiybGSktqQ/U7lZXOsGDXjztXpVbuW1WjEmsHMSBI+rKwytD6xp5HNyQUZDY1v
wvCalJuU0YrtuZlCqPb0Uq4EER6R5zBEjTTFeOPSjpoUaC0SJAqnZuNfbDZVErNe
TeMHhd7VHoWEbvz9j/Tke61+f69sSb75Tg6pCKWBojslswFN/acZyTd6dLxtHbLa
N79tdiuYLHHb9KdCxsuRb+WYMs4oZ20FQtBVKh/WmrJIKZq0npLo5zuaVpPqag17
N7And+C/CrVsdEF3cZ+8xyjExVX8YGC6JHDHGEUVg8qN5W1yExfocxUd+9wTRtuH
YGWJIJ7HDGlqR8g0eIIZSYmaA9AiJSqwaEci7aH3crO9OzMZMQWbJGZXVcxGv010
E0C9iCJBOhkeS0FSetgQo2ieVr25TWCcmBJaOMsWEYBulLH7iaTwyeb6lZ7Q+wOt
erWXZJrIdovYvkkj9EwhuXZQZxxTr30DBrTzUl5aVjBhbu2QbI5Dm0b7nbbOPlK/
pVvcy+WzOiT8DNTyGzJi4zS4qJB3OBdINWrdBtHO5P5aC33fvRLUtBBbcR4HPAMA
2/D2H2uz1jd1RsGLyWMWVk+b8Dz0wzNi1xYRU1Uxa/Y7BBb3Rx0XgEa8ay0062Es
gNTjrWae4HRPoTgMhExTNbqqWa3AyRRLsFcoAHi7kQf3+GL5Xd412u2a4nS0niYc
Hvq2lDixyK/+Q3fgfbeSknk3kqSQ5rZpZzGRpV4VhmpB0sgD8tla2Y75/pXn23wU
4UE4HA4JhzUnhuHpmhs/D1pC/3WM0O8OWo16q6PWz7QYTRBXEKnqHea6sfhKoIou
CamY0BvQo1mh3GhXKXZ8H04RxfhXUDP8u4Oiv6Z3cf7amtQ1kHLXQWASjI6+SvEi
lNtwXXnR4nllG3QDpgYDJR7t4n6kiXk3MlU9RLb6mmeMf9F6jG+Nfat162kB7SVt
Uu111ySTUcfKy+tBv7gxGw4m91NGpUcuxUOPf7u/EFdO2TbQSyNMuTvKYhCg0uBn
J+vQXyy0ENsRe3qIi5jqlMVpVZADNCVGT0X48uy9dgkx0q0FqHwUF86HpTDtHlNa
n4N5L7G6yHkADGmXqJZYpu/PLqWvj+65kUdKimzRjGQV3YU756y22L6or2Y1x6z4
3Jfw5QgIalJVSwHMsaXWEZ/S+g904D/2B2JI0M8Fw9DtiQYrsDm/hzPyhzsy+zt0
X2i/2sPOxgsMwIiINDCbv64IiX16xzhUP64xNyK9Vz0h9gwcRwupy2C7KEYHolYz
P7lWDo0Wrh5I2aIQoAQsYy/RhAzI7VjUkY625jfO8wTYZzGl+bau/lOG8b7qddyb
o2a/rR+AhlFxztNfFQGQkxMoQZZ/InZHkqxg8KWP6MHDnEeEgGl+s3nzvgl6tVZV
MwVC8jOeNFti6awnYRhE69MnHU2uEujoA5q23seFgvYe+o4RU2rlU/5UbXPzVSns
PBhBlkQAjanKU///irA4U11YXLPlKa1gYJacwlIz/w6djxvc9hHVPaXFpH05EVfm
fDnoYI1jgU4h/noR2ganmO4kseYrp7zsLIOy3b/+6aD/X9c4jrDBiDLr02nlcsnj
AgzOMVV1fClM6TOFXMLS8bDJYLGYL6/RL8P8AeJU6FiDgDz60vyDVAxwRMq+Aogg
yxm7S4/YoLJwQbOJxRevfbSwCGTI1FVn7sHz46vRaYAaz88rxC5efTU0CeIQfF2H
i7582NedZp+gB2QmuJ5XEXzObXRHqpeK608+mkatQzltfhE6KE3zPumCKqGtCM6+
RWa2dOQuvzRHUMJ6nPKeIZw/Z2oMw5QHIN4//FGRQZbC4/9TvsPRZOx/rZr/77zM
j9wGQZaJCtNH0Rse7+LPwy9o7ZFQ+PU0Ywtkbm6kgd/EEyHvCu0ugY6nqiG/cke7
uw2kV9xUq+2ey7HIOCn554XOJXwKV2vGz6nXsYQfU51X21458R6c9tfRHZq2PWxF
DtqqP+puqqzx0Pt8WAB/yHtHB+2Cd8YFgb6Yc3GiCoS1qyU/96p+3rgYRfMiDSfZ
KM+ljngMBgbGlhT8f+a3n1iQ2AJIrnaw1blUBd/3t0unwi1/UWBBmmf8qrVruvau
aLRJRAr3g058HX8Kg/i0Up6SwQV+muGoqFZu+0Ib7FI3A2Pgdgxs5uSF2xq0BlTM
by3Bj3o9hcUARn/l5ZJZjIKGMREDLSG/h/nLMjVvBB3JGgYoUcKIK4EZEZaqKDj9
uJCUBdWW73Rxy/KgZrz+RmEC9UqBWIi9YxyQeWDoEdAf8msT99Ovl3l4/iAVO+U5
3IFDTkR4b+dXKqsiOMRF4QtSUm8thdV5OXyz0RjSSaeUBxphVh5zPKhkWQkXUlye
OETNvHwQNZ8kEclbFettuEzV0nHZEXD8Kns7Fd09W1J+HrTA8i7zfkbS1AdeXrZ3
D4N7XCFobAVfSWbRh4IaFeiX/tUuwFGnjceqTZP+em14KTKP3Cr0E9p2l955R6aM
bWrsdbnWqttjPJ0VRCwfCr5JU7JAxb/Ywr1S7aCTcz08WxDRvCycoSQoE+bcwrWv
vODEFjw1zjFMm0euz/itNVAdYbsf/x0+6aEf8XjYsEPi3hhjWvdsQ3srAIkfdAh4
wHyylaqaOJEO371VflWgghmEyGoQcwutGgdq3X/zh5HSvBIFKO4Ox4RhkyCYR4sw
hHA4m8gjJZZcMz+cN0gqEbyXadNLLGxQ+5RwkP3hnteF9vTJca1tUifCVU1a+bXE
UBTl8K5MrPjalhovVOnI0bu86ferzLjdRBFXyp9K51Vn5zpgeaCnENLUtANV7vI9
5ImIHRDL97Ox0oTOikKZf4d8zvgMZCc/A9ZnPYPZoDcOvMc/Jg+dMRGrTrG1axOO
gUqfNJvlUEIGJcQeDetoHhWEDYpssXwE8LK4O4Ku75B2ujjSenCFFpeGqLBZkdui
LpjFNNKnL/782Cqz527BESqvFlKtypN/DESeFDCMLlJfIF/Eu6fNchMseB9LQd07
DWW0OJed5tuyxcihB+lMcE3ASenJ+74j6qlHZ/BTgt4VszLjmDkjSPIvffC4ZtkT
o44WvfcHiAIc8l3zPMQOI63Z1oUMKVLt2DbO2MMphzc1QYKG4kGdPtubsO8DpHhw
pEJ+bbczl/7/xf+fgG9CeKJCAKBYExLQZEH7El8zfOKGpf+GuwABlu7L9BPTJHvi
dWkCFkkPmbmxLsoh4jZU7DpxWShVALZfyxOvJ4cBLLHhy4q6YB50Jy0H7+j+IBbd
KllyLWixZi3RqfOtLaueL9wmUOOAvsQw+S11Ii+u+PEuCob71DQJQtJjNKE6AT4G
Xh3khvNBGYNJ7jJloecIiZF09dveEyFn3rbfNZhlWBQFYM3FWIAkiKesAS2HI8Au
LQLJlrPIzBLLh6MIFkcshpQRZ6q+bZdBwOHmNZ6v3xNTCk1e9AENzhKnst1/pQD1
GuvrQJCnZHwKTIPYNnhokJoI8RqNBxPJANZthe7dB9c4w3snIzEnl5l678Nrelqe
7cO04HlonUWM2Kn1YtrAQPMJEiQ6yNfWCQTGKRg0/v/P3SOfrqjmbG9OxCCP90fw
qG3WtEnV+suag222p8chJnCiPQvuplkxxXjsa7hxeYfFLmgLbUBzvAnaUEObAzb7
/j/myqq10aQrrflPs8OdPhXTKu8u8bTn2ktOe+TYH3wtijAVV+W1z6OOkUQU/Dcl
bCTkeEW+U/yJk6H2jn1deV00guwtz/4v4HeChL3uP9t94Qel9ttnk96jyqxDXj4t
mMNCBVy+CqsT1d74dbSjsUs4ZIgpRmTb1D+wB5dqEgkswsBi/+YU9itCevzLvBSk
o8wkgvDaC7hWeVw3asaOOyyKjpCgD1/oqllgMbG5OEOBbjvm69UW9nYtnFXrQz/u
gG4r5l0SwzVY7nUYs706sj117y5a4OMoNlnr8TWZQBTHMpZ1rS2qLaaNRIsUhx+y
22/O1u7gLZDYdSN1TCV0/LuvqNQ7U/08fJiHlV6eGz+pMal/4fEG9ZngfpxUuPsB
szc09/b5A54QeLQ7x2xrguvV6dIc5b/it7TQC0weROHvjj7bS5CjkN41dSKxjA8F
lx/fTfPLNOFoScNnPI5DZjpqBdCYZ0k9kWbdoH1ifd+asJFN/Wst0ZvP6GSJfxkv
nudW7WXOa3h0JCvC+trFxCQ5faUxzJkWWVEt2pDkTonD/WDCqeS4+JuMx1HQXgt9
zS8JoBz/7Yb9SPqhwf3jsyhKHnPVvhwzpVbxYtQf14CCAEfnN7rQ5IeGrDebQMwI
Dc4r5FcQYr8t82qLmCOagWUI6pCJuqcyUOJ42qxLG7MdFypwVpo0lRFwDdKY+AXq
yxCn198gQ8EqCGqiqxWyhmQzP867dwqNivWpGieeHaJQJB7vcT0/noB+c8NU5uiM
j2a/OR6Zm2kgvF2eq+lZLzpRFd8+u03ujG3TPYSCmtsue620fD5sdnMyYWbotq+/
0PU0LnBchs/ka0Fi7MBQy7RKZe0OH+M+GLsvwctQTzLQ5Ad40blr9vKP62S/py2d
k1yS7OsLlwf9gb6GRk4ciVVBMIA1bNcCTFVHAqWIZJPLM9iMZj8QyJb7K+UGWxYP
SXw8ez3eD0qzW6XYdUIogjg2z9eScSktHP4v95BB0E8c32vJkDasyNdA/p3YWqKh
4thGdNKh3qb7pR5f20RSwjLkds7X/Auyl4+MDDc7wXBuFQDrZGrXlWTv3Wh7MF6e
d3TWEIPNhYIwHKeUc2Qkd/1yvLpql9Eakj57RkZzkTuBKQYZWXJXaBS6K3JFuQqC
/dacn93ClfmgC2dfSh2IOmrL6/res6MWNHYkaJFPycPaU4Kh7LSHaZFryYtzPK+i
/sXNVMbOZqyFgzThgvGbA4menq1ELvddwGXhaS2Er9DxhzvC8aJlE5CgHRh+FCLM
XwbdN0sn6jOS4nH5VJ0kLFGm2mrnFAyhtnSmbjoNtJSqhk5HRh02ivqqstonmVzJ
Pz91ij6oHfYiuiQPW25c1pnxYSK+t1jOkhmmkRUvrxEL+nvxuh5Vq2smOIC891+J
v1NjiwqbQ2A0/KOeFura3ZvemZjH2fhGGgWzpckdK3yvHZ84BZY+2KQmBlpjMJVh
8IvDl3E72Pf1X4vBrh0faQhoe/vLTXBZkJxbVm5YYEcZwzOXWIYPweALffN8gnSJ
rhA8YJv23MxD4QRI4ersvKx/5M5LY1E0zkgsYRTV4Tb8EhwSf9PS7RsAleoisGrY
ar9UB9d2c9iCZEB7uavt7OFeXCqVCQwayfa87l74TfWCKTTpHgKCMunkVNCYxPVL
92EfY6UXKaR1OOxb2YZyDP9KKcZaN00S3T8sRWUEh6nQ5wI8njv0JH+Y+FK3JWDm
OxNq+GphBT6S8//PuWC7v69fjYzYg8zcjh23x+Gm4lis3yOn5RDIVGmgWjJP9VVV
Y4V3DluQnR2kRulQUhGbdWfnLX9+WVP0nfnmLUpigeNXAT3ZwZIlAU6PuAprbPWJ
I1aECb5ky/2p7QxPgOEj4/Rfyl8iZcBebJ/BREQ3o+sZ4gKlsQ4JycaCHMbGCwIW
RufNcBVJmnWm4CoeH6VVVDOR25Snxvh6bELdHZj+9lKh204H3RCF1ljW3u2REHIF
EFWgQY7tj5Fzpz5L8Hit85+uryZN0i/Sl823KScP4Y9MZkGdrtDB50gYDJFoMi3j
//wn81jJz3//MtTV/eZSml5aBrlGjBrZzG4msSi+eWJ4Lvfp7vyPgxJTas9Hf2f7
0V769ZYsOFSXlYJe+Tiao5Mkf8dTNyB7XynCUZWcuStVRUOgpt82nGQRhnzF1ONy
GGdFKazbJYroXB4QpmoxgFvnA/pN9x9tEnqCUQQDAtJQ1LCvfx1HdEnh/ljnnxJT
d9PE+b+HzOo+UyS0SePHPsVXDdP5YPPNlAMkt9FWMaJOSzRGVPW94uZ1/Eff1CHS
PV7Rapge8KA5okA3MhDak7t13pHLQ4RfMmlIannVjsTThoceHCGK4lxNNenagh6W
4O5qAIsw6VfDaP+wEJ+IFGC8pErWJqttOpnEwe9SfapJC6H52JDjMCKzDIAAsBAo
HBmwi2Q3eC+xuoVgSsQT6gXgUhA/Qe38n8w5A7MRa2skMfNoYjuy70pYzxs0KfQS
0JvozMZZF/r2PshoOh9Jf8nYG9aMmI2xMyIKJZq5D0PghE7H2DIOhDaDvaM/G41/
Ig5+a1xBCjlCbFEtPRCKjNDWs3goKedRUBASwqXJ9kG+d3HGKrYrTQ7T07dJ1LIN
XyMRFNnFuL5twgTmG6D8Hk/vAIG65db5MakTW8EZ6UHvvde1FveG0Yog3jfpObN1
e9IA5kciPR+O1sZddYyBMXSjipgVZjepc8xVcWCDUKiJh9Q3mKSnyZSNGcjicOGC
SSLgJrR/iYGwinPipoDtdapUq1PNmG9LkQO2uTWTpHKmgI6d8aCAjKSoPbe0EAbx
lP9NFt24IBt8w7BdzlG9WOs1fSfMtP4KmJP+K/pdnEFhavDMtQfBzQw/40Q8CNUg
fuOSK3yWo43DAuNRvLDxe/VzrCqxL+MdL0BQXRxNzQqj2eCOUxOauVqHgucvFhrI
zPP3sOnAWoK1daR4ZpSFwkXXG9C2kM3zs8+NfBvSjIetgFT1g92cB1CAH562tMEv
M6u5X6ibT74Pm8VUSEfndKA5SRZiIv2LhPnx/L8FuHuOcbH8uS4ufwGaHF1ByW5K
SlMDQRkVQLXpf/WAGrz/+KegH1kLIT1ZtP6kmo4RPEP3Hovxbmrf8Ks9CJwCyIhb
/a+0NlAzjuecfkgat4jtijIuNWBX/5oaz2D0Tn5mdD0nzsyRj1W9pBVZN6IsY3oW
aAIoYyat11NQaHqAFOUh7h6d1bsrp0I4InZ28CY+YSH0jl2TR55/q/lTcoWBhwmq
FDi1YLdWyKiyiCVojsjmSK1sl8zhFNhzFpMqsQPdT/mZ7NxoMbalCMvI8OncnU3I
oGkci/9H05XncXarCGr4u/pV5WEA5IE/aDM8R2PowZCa5mX15ZfkDvPB19ukHL1W
ybvE9d2iaLcPGH6uDDITmgEKJ+AmvoxHjSfny9Yu+v6wqrpyryiYp+Yx2YdDKreC
q3wx7AVYXEShfzV/P25IAq1KiNt5yyKR733BWh2MbHISXTDS/wBMrmSXdUQkrAKA
6jIzsLJwtm1T59IX65BLeaqhEZWWK5Y1fslgsl9WdbCKCoiyAJQ37+vqZ2zC01k4
2SPz1Uh7ylx2leGdoaPLb3J/KZ6yKn7hukhSPJdZ+7LHdM7QkeUgwRq3+blhvWWq
F26B6HtCNIdrT7HIUWFtJZcBxCgmY13nA4yJTcKo7B3lQBJ1VWhrpR76ZLoFteoe
JuxCv37PMk9Rj9wtNdOJ41JNdc05O/SDe6IS6nwY4yUqDC7Cc2wnVtZ/p988fLv3
rk87f6vD/DTC5HhiKOqSC3CwKvE+jOzAJ7UizWSbWiGylavGq8/85mho6zYk5CTU
aKQ3/2JykSS1BkHjW9s0UQNoTPR0qWDrOBAIRb+LWmdVtjR0rpvmgWq1f/fU2MOO
HNq1VVRKFTkyQ5yDJoP6WnhIPPGA0A0cvTuMJLj/HQBdsBXCn3sSsqBQPgzmV0QF
Z0UAqiiXzJHnVRc8S35GZ7njqmiwHC4ZOgSDchlpZd7vb4pDVwMeDS3clQr8Nzxi
9WWn2yVSA8+6t1kQHe98EweAuy6ND88H+Mgze4nBz4olVcJmzBETlHFsWZgz51c7
d+caFEUAUjQwFqtiOvAMtp0t+IXoCoKuxuxrU0Hrxs3mD4TtPKxKBvukLmrkDMtu
kv3/LGQm3cV7t/o149ohHh2EaijfbtVstV8/ZuhXtRcoQOc2PDz0/cCg3XmSXiHQ
WFHxrDxNGABDNXKjM6d2i1v+Jinyz3HYD35EFwYywNHosvmm5EffeMfLWrQaByVa
OFldum0GgWCUqh89bVPPgUYSaXKZxIZNMuWhdTPwnBmTQ02WvJl685z3m+QCazYR
AsiWmi4KqUQVqRby5U0a/oB2ChL4nY+LonXaYWK1ouj8WjFNC0RlEsHIQbdpi6LV
11ZgKZuGj0efUmzadL30Qw/Ca2fGiUz4EBJIpHqOhTWSRmQtYXqp4nZsGvOfiRdg
mExmswrCs21SS+Cq+aC8kTBi3owWyB5vRT0TzaHomq6ydkZFoEYpg09osCXxzI43
mUkBfB52mPxcEpGvXj2zAWU939CrFYRTPJojHOXxg873XdTQLptzXZhMITNngSA2
MUnWHTSVc4so2cOQfsKEPmgbDav2kPikB8OjiXEyXSF/mmRJTqutX0DyIEEPmOEF
Ry35ikpLYd/4DuWmFUdc6IaHmUw7btJJgbxHMg4p7cN5xYUG6Am5so/SGSrpZHH7
oUIfApzrIYkM0Hhf67MoreWMDO5PusNCTC4XPOM4V8LzuStRXpBAOolvsuDc6mWu
/SJYQ8ttrcY4Z4q3Sub4aUnZvl5UbZ73YHg3YDB+bs3rGXr36x0aHd2MLzsI9by+
H2k13fOVeWyp9I6M90+aewvCdZyqUsimTnrQptbXTzfuzme5HO1/iw7EHvtewXBB
9oaTh8IvGpHxixkygL7VqK//FEHKUkMNEW/UtaThcwlaFzCCrn+fuX23ltpQXICW
RPueFa8SFpLgf/c7ZfFttr1xTxILbZVuJ5Osamk6H44286OIqUwIOF08LEBJyDEE
EoGhBaRtLbs8SR/cTpoCn2/f6hwiNE4OX/aOGMgI/6nmw3oZhMG9CB31Akk7cDAS
KoiRRUhp0DN3zEeBpGW+0LBgWaO413zd4UQr5XezA5a/pfDJSKplOGeWv8TqYOJb
MYEJqsEuqwldbPg98NaT0ngCrfyDlazuszCQ3EBas0RacbGzFyux5QEQg7W2GNDZ
HmVq162P1STe5FGegF3uff5UrI56m066nam3Bur5ol6bbu7U2qM13LEAxyrGZ3s6
+cFW0jC5TDsaBR2BPTI1FYrVL1PD9BsqKOSZ9LCt2ipEuErOcYKFurmK+4Sy+2UD
UT2dAzasMUxWeuAJI2mXA2B5uLMdzJDn6ad9uOUnGKik7sLdlzKu+aFpVzNxoF0a
USpbVtfzMaXaitxEi6YzV6PiCv3olJMOQuYFVSan5TcLKesuf1vx/K2lLreZt08B
Mcq29ECUk+DR8gIM1GpYWaCDWWgOuEDTVABHPp78wENd8StMwsMOQgiMHJ0u5Ldx
bb7KEg56JkkOiFpBt+iKG/YumgWxYT6VLJVETtf6+CWhFA5yJJfhD/iKDkYDgeHi
BYwW6hZu6mSOIVjx2b5uSNl5XZ9cZ/f9x7i4h/edy6P0/0PiEVmuSLDLIe4DljUC
OlChafCOrglFhzsm86snc6dDcw1MAq6X4Mt1eEOOUsh+m4OjCgD/KW+9/+UN9Ckb
gDY5BaA/dvi90HlCAHUC3oxAu/wBBhbqxmJ/25FA4BG3gvFmlzZPej4YLOBiR1Zc
JpCSAY3sZvwisTDsfA8nuc/2Ab6Z6SrQyGdhRs/p4OuBVloIBUO4W0xpWTemO3X0
4T/DY8gx+FK6p8hEPVofXgMn1MHX+wSImKiPD85Va+Kd7+txsXn2jAIM0OdbnKzB
4sfthYAR3PCGLARQ/c4B7X0VZQzC5q2OBpXg60Tkg1fO9HvQt/Ht257uJfA75A4f
b7a1vbf2Uho/uiGClrzN9jWZw90ci4WsJlNs5w2Mf17juPc+tUm2yJNkJXIObW2p
laTAHYmqTxAex3+GjE6txRWsWrwWpK8BRvuANTCJVmgERl9JZUCirDvShbhTAlCE
FficUAqcYu0f/N04N3m9+q7DvtrvL40wYdF29b+4HmNGpMC8eIsMfR6dehSaJGPH
V7fq7y6wA6WBeRx4WnJudduj5ylU+xJ7wFBcoLw0ZzXIgxsq5bETUMc7fZ/9PIgD
lXdtPYAArqhTqk282I1Pmq0s9vdUgumKNHyU6gCJgL651jrPjdbizEjnmZmRL7Ut
Zp2itJc1HQVwuVXzTIgl2nVGhOZA6gkAm1xgVvF6e5Ree060aTvggfdKxN/cNvW2
mJ6ThtjHl3jCx+u2NU+4+HlgpmwkJ8mDFgUT0T459gEkauvk+eT/kL1+6dR7Oahw
fuYSa17v1w5WxaOeXLoNrlzSi+MdhIslcy0wxG0YHcTb8GAD5C4Z2BnkHBQgdzHG
d4sSRzcVFAiOrsAD8On/sR3z1JQ1oGCQ6lYofJdFHv6Dv+03jjJoL5a/juUTPyUu
6jXi8pTXK+XkzQsbj55mFdLchu6mTCTD8YWfcmgkzzvn0d0ffTksbvGUW9UMp5TK
fn7KjyZGY+lvx6Vn1kbVZlEXOMfmfZKQssTUUFbXbMiWZFRYBBz+WiWb0slMzV7o
SnNGk4FPvMK7pMrHvtlo0yuquojOlyW6tmAnpgV5iCxGGWZPGMT2y38RxFRi2x9x
TwARcNXasv/D8fdyB+64zAI1NB5T2mMj4zTcFizcAUWgBv5aZSmdaiuQ50mqE+io
rlz5A1Fon6G3b+k0iwfvN+QYlZTkddxKuPxFSNQFWACvhvf32Sw9w2bfNoJnR7Yv
t1gZbIc7vm21orJhL+4HhfgVmvXPmhIWMjb8KqjnlsD0Q3YrKYtFRurrByGItbbk
qN89m5pRm1IhnH9+re6PibW12XqG4wVlZ2pdFCN7iUj7Ov/3g716nl19uzKCLLnR
3ujsfut6PTY/v61EAe2rh4eqsQrTEDKUcEzjPg17BCsDpy5s7HUfrs+pZL+wzVQ/
LqjuI4lCdGka+TFqQbcPORiRBC0Gu7LUaJ8L2YwoJbtnWmyQF1q64CPmGaMRcpT/
FSspDFiKfHy1j3sAUj+muB1/neIpOt9JG8n78leC883c5e29IE1ixI4bRTBM8geN
Um3qdbj2nzJuxjTZoa0RPoVz8fn4FtZ6AYDz/ikPNfYMqkRBx00FWvbytlozcQzX
yZpAu6GosPjV4Ytj0ge4PNnpFNWtrupgAuN4wo7OM4kFqNWIPQR5Ekp/5E4X1i5i
r03MddLHeVpmUWN/aOp5sW+WqBOoogYGqe8fO9C1h4PXqRjIvwkO6RGj+ph3GaYO
/QC/YTwn0NlX/+bj4wxK/GR6p7dYKEOgFg/2QOwPjeeR2CEikVTvMDWvo44IphDY
A5+XwBCQ5ymfEpjzQAuIDmKHtAaGUp6yRmwoAx7HhOQRKx8u9CR9H8q+m0UZwKq2
+l2APBNH4dHRTLxh2Sn+G8jgyAvhycDzL5gezSfYjRSksfp7DAjVIoOclvCBVaTA
/hMu5cRz2pnx+bZ/gQWI/5hmGPNZC8nMNEHOuwBfr/7wW4soH2eI1Vcb4/zlyTI/
irQwEGVZNutC/C7GJ+TSwCnCqUj2zI3znnXlllTAvQAx70Ol2Q45HotrN9vF2nvp
v1BlJyewJCjTY2S+RcQ+i18T6IhXB5/XNVhkkZlWS6dkt3dJ3iMuie17Sl9VQ8JF
U2pPVNLnYYzv63CJ/6pEvmI+8Pqgi0mAolZI4pied04Er81XpSPTFZFXfvO62ZQQ
UR1vAxu8uuLkdnddHT0JHUVaD26qzQfzHmac9mD15vXwh2zRityAz8vbHN2VBFV5
2Qct/iGwSMqhZo6Fii9rDVSW0PEwZ30lK5xk8Y1YdcQlOOE1HD4YMbsN1JarP94o
C93FG9Ybxetha1vEs0j2qaECWsSKXhnI3b2wvg30/h9Pth1gTvQXsvuTK3WmBsjt
mDvhH204c+qwiqUeXcjKsfLWZTurrrGJ5KxtvRMXmeUM6rP9j7QgOJkvOIRouhEj
dYkh3TSKAJeq3BjAHs5quGrfaQlc/t4eFhqHboWKrsq+FLESpkn1mYPkIgHvkkVn
7iYJ3+U3id5QOCK/YRTNLOC6nuh9G9fTAepjs+rak9swyO9kEi0tQ9DTwalf0Dt9
CfGLeShm0+QJ9dIL+RIaRQXdZjxkFiiVKDwekWJ11+zos7OAjCyRyVmTYuiPAvQz
rSEfz7uJhkpkqnTMRJ+Xy1aIYT/WSf23/lWa/P8Gx2V+9YfxnkpOr6i7p93/7Moa
9BjlGIoOvLuWiyg5E2tcR1X3wEEOnTz4aZ0ozAnwtTUAyoyfWZvtHbJSzEL+gx9i
p4krIe8vXdftDzQGB+46WDUooHi+sEplTzMo0jXuAIaBfsWmd9kA6ysOLFj5sf9X
6qGTuLV5uT53Ibt3Fr9CGRf5YnO4FMMFck9pD0oLSv1ARVvVBCeCGIUwUivhwP9I
q/jBooIgTX9s4uK77AM6o1pXasQBSB4CmJPdWzw6dndxXd0cRPiuFifbE/wel0WX
6K+2MFuur+p3nn8oPj6OgHtki3vgITXc0aW8gjd+tbwYxVoFjRduR3M1/1rc75OE
REyhPrI9Yc5k0mxVzTDlYS5E9C/NsWywwGz1pv6dKBkCB3w58ReaypWu5jjA7EPc
S4Jn4TMcWbVD5qQR5baGH2aC2MyUh8KV9yf3YBAtESkzt/pcza0UMVEt1CDenV9j
fblxCT7Z7XHQxQqatM4M0YdRpYrsp7OfCf3MY/hfWqZa5rFXDY/N4+7YHdvfeGEP
bZQEpd9oGSTWKylyR/gAmH7Ch5AGXVh2HkKZCHHBZWgLXlM6gUo4VQ7ay1mifqaq
xfS6ycFuIyQHNb2EeXADB6Q1o0YYFNeqkEuF+fLuh/OKWyhBh564yPl0gCoSqQip
t9YtHT7wkzoTk2OjicZ14fxSGTCmLgAdIf9sHXnpn/hdiYobgkuhHKCDy0wJ54j+
jqgU8mMRgMvknUlayKZirWAlR1S6aMbTCQ5uM8Z+Pw7eWL0BMoo7JzgD2B9bKeF3
fBOCmj7zp0Jka5Lf2rgMCaicug6C1kRk1Ha03v8xjoRB3flCT3dCmwOGFCNMq7eb
pKSi+smW2hjRbY1fw9JdyCt9ws9xcpyNi7Jx59najYJHVQzYT6MMxc6ipRotE1zy
NkJDvW7H3+kCOn8AAsAzvEQaPFEXIXB/AycH3hBVojHgl0zbP19ur0wesiUBNRZI
dalECdzl01k/Dw+U2EJzrANTBVkCHVj/BpmqTVLD6mcN7kmZ9esoufKLhsnn1ERq
kks222KoHGklaIbL1jARN4CI3/KVSY6V+v7CNE+DOi9D7zZIQAP8P8/6igVB/zrK
Z2okUKHVdXbQ/Pzz6ViYgw6hyZvw0nD14WZAdj4Cw0LXe8pIfRUuxp7lK/29FgVz
sdD2Gt9NJA+sJQqJiEIfVlxQpP910avLef4TDb03/P4tkLC9O5J7ic+xCEGZEkS/
dmInYPMns407LzwqcINi3RJnh0zUlgwVY4EVgWaK8qBCG0roRtvM5XqD/5kE3ejd
9b6o/tom5xgiwMF9HjTfps+1mUm8ZoqyaU4Z71XNDOSv1zfoRFJkXmb8C9XKmya5
A6WPI/nlVHECfaiBd9/A+ybbSQxqNmEeC+CfR5EjR3AHUdyLEEzhczIPMlgBB0qh
7RIKNZNzStiXpvFY9B3EpKevgnc2fWKazkAun5Nj4w0PkJGTKAmB6gq49DNqvedv
VSweFxJJ0EBNaduu2XGiEXSr/5Etfn0es08Pa79QwiAukWxH4oDNWS7rskEuSgXJ
9kOSHN+LkTBtU7Ka2fFYUDCmuQogLwue0Qbjb0waPY7/qoXnVWh0cXYIPK+hIDau
ime8xuFwP6dUyP69xnRbZwrrSA4x/5NmT0aMjJA/hNSqc/3sc+1opLINe4gupD5z
ImxGqxs1dsr828bFAaiUWP9U8oIo9HLLxAbYZPG0cqiw5tOUW0cRmo3Dn/DgSyd9
T8If3WaWCRtJDoBhkhPLLbYtann+BWcZfP+pnj0dmC4fSc+m3nsPWBLk/qK7IVpp
sx5adtcaueak/BV/TA+9vtjVHa9hkdZLoAUiyecmIia0m9Y8MzN2/ah0x81bTk7k
O8WNORWvJGUoYUeFx5v5Ghi3VHtHuWcw93KNoshI5pBaKTiklR3Wfq8+vKS1jGdE
9sBc0xZKFbYpN3j/Glj+Y+lsfq18LE6A56Vt8CGzYWVFcnCV9geq4x1fZ4axg6eo
s1xB1nozKTTqFS8PAqsAQizDOjySUOG5W3NMiDGmf81wv/xDy+2mcPOXpJhRMvqN
n8lm1URqdTn7Lao/UkFWcOQTSpKtzxpRPTkn1hgzZKd36lCbOp5JLKi2z5kVqIkO
bEqkGPAEBCH347c7f+5pEbDeQSXXVHkzFAr2Kg6dTi8P9Bw+df0p7K2NTzBAPPm9
G+UcW21WJH+btL6TtnsqhMxyGdQ3ZEa7+3Z4yB9D6EalPdArPyJE0MUnUThy1Q/8
6MXAQ+Z7msH5bBDSppD41XWdCrRUJ7AXF0+QGiJG2MVpZcHJK1n3FLmlNDOvh5uC
Zfl3rMmysH4P52epDd2wmrmrNjaY61rCkWpbp0wKtwguWD4sywgx+Dww4qe1fvTj
wuFbEh4vCOscYiVVoInlvDJNCOlUTzl85Z4i5DjWxpF6bQU2l98isMfncw8Aj6ml
LH1V/11tQnlZNLE5o9zjXCyBPe1MKYDt0iNvSlkC58wgR+w9+pt8+PPyy8aLblHU
TGPWyLfAmPnnAUelTW0mVLJJ/Ppui4tzFSMGAxt0vP8+uKoU57e/63ZRcSxyqoVa
s++/ntDdIQ1LXxdppEJu7Q4v/8PcgpZo5kLI+j0NNlN/WcV3S8Vlmm2NnmLuzmnr
h99THp5JTrqZPYabxrnaLn+afgupwm7Fz/FhTzRBpzFARtzjWlm8CsyoASyrR/M8
dg4bkobUt4QjS8w8Vk8SGNiDxrI1SzaaCX1aidXzL+iBgQc3kShXzphYUHmcZ1n9
hTfs87pGZmlCaayEh9Sf1NLOutNVcLK4hp5N07IHEm8OKhDv1EW4+JiZ1JLZZH8A
ycqVH8ABe5zIz5W1fpTVsGWCJXLEGyLzoWbacU6dXP3h0u6nop41SwqQ9iyU4+/B
eZpOLogTVEQo8x/tyMUBh7UYmE/VNxuhPhiDXQCNer9FvpW5IEvWa2ae4O9JFUXp
VCLM+yjy8e2o9Xq18NcLBQcjjLEtSz7xN2ufcUE6GesOtBI3iD3UsOrNYqQGniTY
wcNSn4s9iaqQgUA9fzLj35dmRwm7+2pPIexzC+w0Jl6D6znzI7c2yyyz1ieP+p2L
RV9fcUf7bobW+FUb+c3gna+wpCZs4aTKG5ULtz9xC2UoXg40YR4jh4I5FsneNz0n
nCLUSOITsh3tCYMlVfVCcgLqke5ZdNFtDxmVnt1ITAAtptWJ+I70r4AbWzagNqpZ
+ExNetpMWX7qX68L+x7Rh5UgvezqcpXcjSepC09dGytRT1V3X5yhSXE97sL4KMSN
9aIN7/5ALgcqo+HbsqYuQ6SFzVqEEV6sk7kgrLaEN1jY/c1n1dsAjh7zJvCP8VcX
Z0l7u/GnVTHAcLWoPFxzFN5cpO2wSN+6UgeoWrMF2o234iF7FAt5svX5yf//sG+U
AWjyOvBFJKAZV8EdcMx6WiqOgeU0fNsTHHmbUug3uvHiMVvMmMgDO6P+rBhzMWh4
T1Z5ZT5rLRjR0P6gKUEcar6q6YY5mxZRRuZQ49BNllMWUO2hwsvKQIWPnZLnWjbC
KINqjrA1tTujNIneuDgTx6CMo6OeInnimCVIooW2WquydDDfeOcJGU0gmU9dup3g
CD9+GqR7MIttSo+1O/dyC7JU/9kxf0Q5l72koRxnTgnWYg3vf21s1eJfMYhM1okj
D+pjCvntj30QabNxEjtdyPeCeMUiLNuYcKr5h0+PGNxriToSkk+yYN8gp5u4G8mN
ahYQgpCc3/1Yikvvt9mycN6xcb9etJ6/vLE75wK+kun/6mpvOXGcj5mShlAGPvYF
sw8O03CPvLuIsklygmWrPPemwhuKQreJqRVVn4h27Cj0w4BpJA7zpS9XqqVqjHZQ
XXYcf/kkxoFM8dVmIw68wMLUCIO0oHsyhdZbHS34tzubsSrvU6lzPN7yr6U/grrM
XB4qM/CUKUWIhNVu9bLGDVPmWv2IL/w6oJdLXB4H/82GJiikauObGbkXudBwq24Q
xz+8SDm6ij4xT56IF855ZLjn8dPiaxRhOJyU20euJAMTUH0W0LeOpIiDq0tiXgeN
xH4egGV26ECNH3G7h7x3pLzNlYL/gIUQGllAkiCjKfZ9iGOUYd44CzzC6uX6TjZ9
Gcx0N63CMhRzKjGZjieC7qtNWci994ZPU7l33tei1P+7hp3lQYAu70x7wHRVk8Ve
A3WxtbSTYeNmH7a/FJ8RcCaRg2hPQX2uxINUN0mGzIDjJ6TI+xKNN+o7V5cYn4AV
fqxNQVnJFPjXmCZsrxnamLkveRFd978K9CLeGSaAPOLVF/Zph2h/CM12OBEPBSam
vrRopH6kk5N4ZhhurLoxl7+qZltVYNsSGgX9w3Fbbc5sxDL33BNC8ILJhW/FG/Jf
ycgbXLqXQ+OKgo8VvqcXLu59WJwdSG39FmT1LD+WkWnXMazjx0pmGRd5vXLOml51
qhGNXaBVEaFQKNXnieM+492GpJAHcDNr920he0N1rcAh9piS4J563kd1RWMYxj3R
hGaW6l3ovbRz+WpkHooxDFZ3wJoktFRdUUanCaSVHWlrv6qhtRIwyxFUqmPx9Akn
JlHq0Y7n2soHA3n/X04qrQDNAeuWwjYZWY+1p3I2Mlg9w7jVuVvJ01b0y4XcCXDu
dhtvhsZP7IhGzUjbeE+P/FUWBnwgNnuimBIMdok2kPaVNLbtqJRxHmPYzYvSNcHx
zI31czwgzdtLmFBF/vOR9NksCZw2MzTMlJkWjDZ+mGl6yDasQqCO1mSpvTjyB3+V
d2ireXamZgluVtX7nunN4484vwVJMumChQqanz1zcvg15xGwweEVxE4X5Ol1SVIL
ezhlbBSpn0WS4QxOeu+PTg4f8J4iC5syFNPLlHy802Go2aj4Y5IK6OmA2cp3eb05
/tJu3Ddf99I5QqhkrnwDBgXpeQ3Q0m2kAWInfhnH2JFyu+Pa7D/lE6q1QFuDe5+P
WPlSdDUfR0qq8LBrH61XFdOXgvuhhwVl6+sTWDlxEOcQ5Ntm+zr4zZAxlBI4XOlG
IxS70EOq3Z4HNa/2XcI2YPSWD+KPjelxgnPcJuwGpqLMrQ1TO3jdutDpSCmuiMbN
PgxL+Ykt/oTkdLfEfaWlJ+/DAfV0MY6qFXUmJiCpeMPkdY3gD96XdSSo/cEp2nbZ
bRferUOeASe1piVsSsEyal48uXPeHQFHByIPkNYppHEVzuT6aT3DaSPxJHnza7pC
AbH5L2GSFIDS+Qt45jtCIJRVrBIwtSw2QyA/9BhJahP0ZJ5JrkZYncHSe2tw+VdU
bxcy5uLm+unbTrEDmBpw69fe+Ph72+41zRwhKo68+0Ffau4lGOxQyh1CIzEwW/pH
tn2dAP5ZE4xyFzFjJOLSNKjy/SbcNb4lcDitgoRJd7i3bi3neVzZwvB1FBRSo5iD
EIS1NSyC9TLIMo0mecqnBknpLd3yAtVlSZfEQED70U31+tv6YE702DWUbCefD2Ne
DBN4/krCgFUwF/zU+Q8WVPN+HzjTV8LebVaMWOrzlYRXxqWxrF9/y67z41+S50bp
PulDDNRYUTl/SZy4mNrIXFnk0Z+JLl7jQksJZCnYtW5fKVjl5hzXHpRb6/r+7I1y
T1r2b3kSlnT7MbdNFh5NEiUjha0g7bOsD8Q5Xi5pJzi0GoaZmyI7U69QVBgVmgBO
ZMWxxYhSGy4D/KBiw342A1fLDLjku3UZTj5MYRTpTXbzFrMQPrCs5UkPs/76flNw
3dQPMQRncxfmFPSnh/m1iADZYcQ6gQCgjP/2a1AbggT6lZHHwqsYfjI89rj6nFw1
k5jkjXbPWWX3tfQTFDx1L53qDVFJKkRCDBl5yQJ2EDt49m+HJdvKJ234mU5QWxqj
lH0mv9RA4SmA762XEzCJ8LZqkoGnspQtMLOtGhXL8mPt7uJicKYWd1JjYTpZYsnj
nF8Fqm/1i7JhCHdPfevubvRdLlLyvOjutScA1cxv6EOfDo/PFO7In/Ju1bpa9Z/3
/buhlecq3OC2nv3kQtXBCZKJ89xs7j7JtPDZAI3OSNQjhXChGsxOP+vzRzT7E9ja
V2CRuuAychgrNqnyCgefNCIpCm3rLjOdy/AbwSKh1nv/wHM76osf20haBswuBwJi
U0cJiNbZgABD/Rd6YotH6VUQ34sYE4UHLD6kLId6NPQ2vTAv82qKrY9diVyHrc96
Ne50XEFIbTv7Tr/54Am5Y2Rw2a6zAU5B3m6JhLUy1qHsB3LoksmWka637UZiH04C
yktKUZamDHr6gL4pPN4ougYS2xwqpFqmuH+tVXNMI50rmFsJFa41cM/cdHx+85Es
E6N0qgphRLAJX9MKVUBZUoa7Y/yI9CyRJRncUljp6ADgJpCLMvWOh2HyNRVoss+b
z5qj68WgzkW1u8i7tLeFrC32YIgXCIcjVJnVCF22haTHIYTAkD4dHzKe1x/wmofc
iaJybNpJlnfcStMPZP01AOis5HV+B4QdRkJ9WgjLl/vpVMjbezS8HIuuz2xX0I1f
T8a/5NTRl6p+CUKnl/0P7p7LY52pyIWaY8MAE+8OxpuKaae4A/sR3zGlMt2Wy3eM
5YEPLyt+P/NNjAmQDrnHkrzvGryJb7cuuhiIkWhjM4zupbabKoGpBklhi7QGWYLv
la7+U8ia5i664wG6vmZqAJfTGgwd9XPVIeP2VJp4FtQUb2Fy/Ox5hLnl/SbmdS4T
02KCObNqEpW1auJkanHbI5x2/pjbIGxXHHfLHQza4KEoTuOLc5mCSO0QAlDsXTDW
g8q5vzoA5JggQnllM7XwqH1iudjiwfJbCg46/5t9yC+j0L0/0+9N/XiDtJNFvOil
l2DleOVu0bYaiA9O2GcakY5nkZdNrJaPQAtWOds4SPWYyU4gQ0u85Wnz0PHvGudi
4MNTo2/o7804M5ZftA1FqnB63E+5F+iQcP4s8ONYd8KJObrYVrCBbf11TbCdYsgD
S/H/ZEBUIorIQMAg36m7NkkxuiwIWXh1kSiyjKDJ5ZMy8gkDHf+F06YgdI228vzF
5sMs3/u/xAjBMcOsO0Dznh4FHrANsLmVY1oyB1syVGHWdTerUQP3Lsc62fOEIzla
TRG+KcbVdZvEzJMPqjOLNkP0101BrNzYp+oaTHiRboFIZP7MP+1IYXWYijbXUzNG
J5w0SWfEiBKg6pw2Q2Kn/Tp7THAhhrN5emBVTTX4zWo+dexXAekCmhw0av5vQe7t
fvNiVnQ2XJSnNcUHSrnpmwXHr/IFnjh2M4HDnORAFAE/XENxcec0iaIqdA3cCrg6
whHNtgpalhzd30jrSkvHGIHfWC4WruWSPRfkLRVf8LP0sv6tv4nJRw0fUgk0n7Ur
LkKz0OAyJkmvUFfoZVpZi2sD/tLpmleHOb9JnKoiEq7LCSWl2q08YelB0be46iGb
znuSVEXs3lIbpZ1q0fJizF6XXCx5qy+t2E+gd/Kt7EDBCIr2VzFNB020KhoFqf6P
TBVK+63koC4221HWtJk9aiz36at4oDCPOTqqv47VflpO4LqTZnq6NTHSD8zsphSX
nj7lswEwGDmvM6KuxCOYFoLzDVRfLDAdbpHv4FbD/9CLliVmQeLmZDsshbz0lTk3
uEWHHpxuQuIOcPUHz6rWk+qDIL/ieo19aft4YEuFd9/c3ckd2iWs0DfXAUwb30MQ
9UTTmIxFANv0dLIxJFDUvaHxy66j88DUG8wyd0tcz+Y2CUW/GvzJ8DZmnRa69532
1foIIGjEM2hLaGXjzq/3zedcNSpvqWf1fjKlLyhgiWVPT4XxpZBTwRb+C4gM6DIp
NWZ5KkY1JcU+ZesVMv0tnvH4+Q/2YJo4U5pQI9y4lDxKMmKX20p4cgvXraXoEbo+
TJxpJIeF4drMP1b0J3MRjmOuAlBj9Ss83zvCQTkB7nVc7FdUrg/Wd3h/+GRU3xyM
YfJLAPRnNMg7jOWPDGYbnde8rIslsYeTTlbedLx64P7y8aq7b2Gm9n2SJlZmCg0E
xg8RVbOCzTajFtuUNaXTXpDic3AY4ggNd/66/nvLq8tKoARIoR/BsaNM0VX4eQFE
4Y3AYJ6gLiOAmoO6QkWMc0yy4TDwDDelKdV/7/RPkiNhm1oHSr5M5YPmBXkFi8x4
vmGQw3lHhTHUzJUDb9gKb4CnSGqHJXikfTyRivrMLf3M95xBwc5DSQ3cNgfH5KjY
xwEsc9GbXNyi71DeEUGKu4ZjnqzMNe34HA0OQgXC2K0bCUuqWMJJJuI4fhuDVSKh
46Q6Nbq5y6GcqMTlLR0Xm4ljSZypv9Votah4d0vPWphFmh5U6TBej1FNPUekiwSL
WvAv5zYXdCA28L7YJlDgWHuU+tVLFT9Up90D4XOlXzcp4tPSh0tyM/Me/ZX85V4B
rjGlfIlHiyZNTeVw7aT/47p+ouvUUzxvy1H9JJ5DNbjHzUzuhVHh7l4EBqEjAQfm
KIxbq1Vamo19J6rjAz9nMd0RjX02nrvMADBoTeE3gcDagJ7VmTigxQDvxxDuQg3+
vK5Hy1iQziTXBQaXffbHReUby3odUBTUVSV7oOYYQXcIQjDYy65p2WIbHJN3xwNs
hx/6Lba6it7YWy+Wpg6XhyMGLU1XRxUgSiqshENAgl5btPh1jKDJkiHXzWj3dx1B
x8wIbhsVM0UG7qC6PIntDQgm6NlR4gqg2dfBrKncZCCFRBHzDuVS2EAvfAuVd8E4
6qg17GmlFdfZzAKhVa1QSUFFJaaf2NQA38ubqKt2tIGcUr57YaOZpBk0Vx25l7l2
1nlo43BwC7yaWxspBM02nhlwmH/zBKuZG211GrLcTyFCskeUL3qKzPqGQINU9N/k
5obN3PgDA0sN55hOA+FAiN0677rNb2PnddzYOw8udi6nTYhMZTXwSSQyG2Fy8OJ/
UMWk1x8g2mVg/ZuECtUOjbYYqcT0N7FvlWrqAJmOuf6yAfAPZpL0FP7zlvXFeG7M
6GSRAIM01aY/RbRnTTrosweTVtRMWYI1UIo98tRD940tYO+I9VYFfgI0WdAQOGeY
dzfRD59gEVe5eMgRD2ByYOxRLZZsw42GJnbuwVRd3ygA8PAYr92lZIotWGLxoZy5
LlsQlK9/FYKJCRLg4tcXANYtbJwpzJQtAecLFIdKpG7tdIBG6gGs9PVVpSexskdb
gZpMLWBiD+R0ON1ov0jdVolpLtudWlQt9gicL0QH9GCkr7hGp6L4uEuZXC6PoOGe
F0khiLOchWeTXMMCFXmvJBkKtGrI8kXaE/v70TYPJouJxVXjc1JbvoZpsE/h3jCh
8mL9NMpSa0mCqoId3UQjPGhcAWUNDLdFIEQIEfZk9os1H/p24at9ZEj5xN8J44pl
M5PuW+aVGZ25vJ9j9yWaO1ZNDJcZQFOeCAm12BJ9HHwnQTWW23oh0PtiJzlRrvW5
umVj/AQY7T6jtk5kdIAMuPOfij2uotmpS6qzsG8d3CofIZnYDAtDOCS+5mvYj7iL
ncue8GUS/WP08li4xr9RIj8dvRCaW3HseF+4fFx7lDRAEqC9y8TG62yrfVQHJjBJ
jpyPaPMHrT25tjqMxgSfGRz/WBCA9lw/8LsgfRA4T3zAiG9EPbl28f+rAO39IgSA
y6sgTb5TLYVKfjhSIYJH7YU+1ACBTU1iSxOiWVScKPytOafZn5r5YVz5ybHLOWsY
GwvfbCE3vAjLdphoJTclfSye57+Ut5c/hRSGVxXi//iRi2DpPpq/j95o31Pkp60f
IyWbp/CKwhY97A3/bRm7lQtJvNGy+/JHCgVO5YRMNVtEV6Zj9wBPFLuGbkvUNNND
nVSk3v+6ewx4c+8fs00CwR71hDNMC0OmNtGQXi3Vw8EJ+SUjqegAmXsKUd4aZ56o
v4DgXr5U5NplY6DVhYV3GOYhCzABfa931W9u/NwxIw1Y+FwWpi7wNbKqYRl6Zs04
rACcRWWbbmvHfJIYyiDzP62XBBmMXH/dhqYyhadcYsU1pkAoPwxrML2fe/qLvDrn
wq7ZGcWJh+2MHAlTdEeLdIm+1rDhvuH7OW0zT3H2Ecl1Wn7UwwWxboeGv9eR+sMf
lIBXmi49kByfk8wmvxIdqn03hfcQczVlDoU8GsLpQsWTstPHvZcZL522G5k8upmn
RRSgQw9c305z+goaNThd6IChZ2zgIV9DY8og+lrm84C0fz6fNnny3qZgZ9/GUBLi
xZwwtvsXTB5aZ5wycLlLUfSGzIdeojjkYa0vYlDiOlAO+vqwA/X+ySHst6am4qEp
SOaJlc65knKPIh2La+f/h5HlTkDMN3FABPCLIsf0VgF32HCflaNznQ4TESX919dE
4zLvPxVRqRfeapg6Wvy08bCXuCRYCah+n9EzJuGfdV/rfxXKGon3fQCa0gctZ2/U
boVLHvaRXdKGxxCzHhQEjQZWhWABnzmdD5v0yPpnfs9715Ps1FESRjRQ/vI/qwOE
5J0dYlIwv4P7upDv7EuawzBalMDetVirPRqwU45XGvatXyHY/Caz9OmGIHL56JEX
vCUo0V9IqVeebW4ebGchvbFxPSfmtsM4P0kcL90Cg/SRFZ9x1LAl0CQXkVPBob64
WpneNfw1iHT+hJr5HYvVXd98Ue8YkhvQGXzgShSqXP6ulKEtOy2VHkMor/2Qu9PK
ob5TKUyvw0RfnchGIehRwBS3llzZumO1TQGyEkl0Qar6gvtnZEdrTWjyH/ICKUjG
kkGIkTdasb70gRABOifitRCqkbRZ8NZEFy7Aih4HBy1DoBG+bYmLbHRLYLMoJxnt
1NRXULty1bbbavQxfv9MpeqzOKH28Hf6hunoCqfaQry7yTJAh4+NqEkR+al2I8Sn
dlX4ug7aVXslrxJUPkWbaJo3/JJfLfAij3yr2Xvm3E+G3KHNB2JMlc7OXeLIRqV4
zt9j7zsU0g2+2RbEIli5XjxnvQe7gX2r/TycBGD5rTVzcQSIUzadSBjL1sRaFNMN
7WKZNu6sypt1T+KX3aJAoz5CO/rcmjwMRtqdew1/dcIUQwaYUtb7XMsgnAVKheuc
m2rKT4pJ3MIw5pNKXfjAaRauXSNKHdcESIA1wZZ6UcNJoUeB/6Jbt0w5Pz2Ejkb2
RjRHSte4+cMs5DSvWLoOCzvRVd75sGsPRI2nG8rMttLcmUjFhLN5KlTItbChm9mM
/7Q7LbU90Ss2KFk013OMXoOW7+YEZVSV1B2ms22JO+NMvtZRGyHKyxRFPlPGpQBq
1tMSerlrrJl4Hc22KwHuwa8e7sU7Axk3mtVsUlk6/XmVuUykZrsrzht11iRYTTLB
x4Veli9BD46jOE49dovbdMCNgkO/lYYT5QU52ewWM1EnrXTPoIoZ0vbit4ogDi+H
gnoY/H1MtHrD/n9HZ+NAROA+7Zej8rrmiDrWtsyFJM9sTpZ+OB1+F6AqFUnHCtrT
bP94ginGv9eVRS+lDenSAhmXHQEWn3dCjozT/6H3ddg6vtSJTCbOXWdy+7nQSAJU
QPcmswEnqp2RubfKWXVFfFXXFoG84z4muiKEm1PLef2YsLbUguHwhxCuCMuhkcEC
s+uNYigI0sxSJMirU13LHg==
`pragma protect end_protected
