// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aby7n75XBQU3yowewmUJj0lZB2a72PY9Pt7gYd5lpHIj4P+2YTDL/M0Vr2zZwb9z
ng5eQHjdS6ezTANNP+P0NyaKWNU6HcxOHhRfivKDCQIcpurxIvRH9jaD/K1eEBA5
GTQlEum9BhSiNhF0BjZYYD50zqNaXU/tqVeKjqN+yKM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6864)
VjGW2LA+ZtcOhu/SzHJqmchtlBFi6rOC1PdeYc5rLNOfTTdXtYjA1R1BQWD1cXS0
t1S9wTEJL+kSnRKlAK/JEI5eoVwTAtIc4bBx5BX6IGIzGR9NcdWv8DjHrEapIdAw
B7Te4ZEzUS0who4iU3Kr/rKX+LGF1C3pM/rN3ABKywgCf8zJJ6Nqz+HNYtthOncF
HwzBGtNRvwboZ1Kni4M9ghObyfUC+8gUzHRvIPkKvGIQF4JrRCnevqzYbvSM5MJv
ZrqeaKJT1LZ+UAR4+bR3vjAcfAZkEW6gxP6CgyOSpTKGd4NlW8hu/YOdyxYMCIj0
c+dPnuByspqhoa5m9b0HhLQoh4uavT7tx4DxVkhx1NX/QkyFkWjbtINTH7l8Yz04
aXIFmxhD+BfZgMNmUkY3noiHhklEn6JTHrAsD4fNmnRu7+bKS/G35wkTQkLgQnKX
jpEWDSXuGAYvLhzrqkpYQHCkQ1CyfhdxSsS3jkT8cxzf0FZ8FI5nbfoxicYYRcrL
L1tyj/LTaY89vWvSIwyeMu81V29UZ96DcxzHxMXhhw+zRMPWdbpw/XwDodtOS44e
e+E/hYmTxbbZlo8lzv5KtT+Y398c17yAoiVqnFEunyGGaQ1QC9q2+BZvCjIHPVeM
AXJszknIT1fu9wMgt2XEUkhf01kNXoJWgU/ao592WQqbBJAgwn6+BbtwJCnWywK1
Io88iYD2wymmxz5TwNycHrE8DEGj+6Igg5UN5c4kaZKhqV/OxHeZ42e/nbz5/Sfy
u9YTlOh9FSxZFS9vgs9BwYCDI13WY5MKzBwwlDPtRhRmsAnr+OWOCPl9N3b7UqYm
GfVi1nStBRqiaBOGqskc0qfMd2GCKyEA6tGDDulShY2IxfScCgxPw0S6CoFbr4cp
rlTeo+uw5bL9FFfM7E8/KjUathyeU1ZO8L9/JzOFujeG9w3yTJ1UwDSafgbi8J0q
HPXxgWQbCjiTWslh/bTwaWTXyXm47KNserGyCFtVXiBPcOajN+QMuiRg9nfrh4FK
1OV+dIahMG1jrq9EDdCImh1nnnlb92iqgghyXSCGsUNp6kRyXd+rhrSiZcmBKuGs
NkbKjujK8FCkVWwAKFB6C3AazbDiW/ijDFOAbM2o23d3Eb5i8ikWTTeisJ/BVsUH
nNyjoCqJ6YMBzhIRlj9Dj9FhIxfLNWL4uEhKAKIbIzyium+4anzgeDQV6Rxz6/z8
yoCpdJX3j7t5wwf85zuxK5FFDcrKv4pV0tOOy7zBdIcfqSEkAFdvtqoIZSJIUhXM
iGlTxyCmL8eEVne2XtQcp2yOW8FpheE//5auA8Si9PAeGg5liAx6zrR6gFrFzyQF
ilNGbLyve99lHlkfvYVjsP+s/53/bes3X2g0srZZnGJOlqqe+Q4rMCSpnDZP0Lik
WVuIj+UXQcMWb3rVObdfv+Y3N4s/PhdpoZYVh26yOrwCXTPjqeCxpzNimVN6kQwT
jF0x+7DRYuwMMRqqSlkNnfa9D7saWbRCs3OetJ/wNVV+ZImfdw+yEhCEbDbLtPIV
MudDCztCe6+dJXhlQfiQUK6Q0a2QFl/19KncimDdy/T++RZIxcBsIhMiUaKNsSoA
nPeNRSEgQDt5SXZ3LPzt4Zezb6djguKSn8KuE2EaOic8aCt0IKCgbplHEPgmc16p
zarDU3xocOU6Y0et2QyOeiTGve998nrSfnA+mXLokN8/Sfs/o9nGVbaXZb+nTBLi
piVJvxy4rNt9C603Pp29jdZbYsgRHclONhlCnBOYqn4lGPUHPq5XXoIf3aQ1wJeq
SLDip0ZRcZnKXnMqu//+LB3hpANWEyWjFX/WoxjyxXd6KssFbVIoim2TAq+it5lk
tHVajdUcCb/ZVGpG8qTIpglqk3xg0okYGVi5KRYuh0TlQ1+yaD1RmU52sFU2uI3i
MT8Cg+59b9PZKwaa3gAseUhT2mLzDNDklFWhYH08NxVgSiyiY5LzXopl3HVixJVO
pLXzii0VeC12y6P5zFtD6cK+RTEeJv9o9m6eIhpRp+NyzfEK4t/JND/w2w6ITHsp
5O66q0BKbrW2wC2Nkv6kKlPcqXlVSadmvvlhYprM/W5I9y2NH43dNt22DAq4REyK
BfK+bwBN9Cu5wIwUiaTGhlCGTHL70VPDHMvQc1RhVE6RVGPwvqB6+3deU74l1dab
uU4cP9v4BJ8MLorQjS0nf+xmf9CJ/Wctob2shvUrlN1ommwbcSxL9oJexvXmgu7W
6w2hiJ9AL7MasU7Sl3RUceRKOb+dIWn0AnGnAqkG0G1d8/yMk6JmUT/UNuPDg595
R/87kM7A4W/nBlItv6yhT+codPIfIf76Tw3SknyAs2XCGRZ5J9+wIZxhcUaJMb2N
cJP1h6ySp1Wb3wM0hm3zYVC0a5JvuRZ9W1SaTcXZVnMn0cdWgrBGkM6bbpGbvDXr
bkZf9ZUuYhiVoPTFvAZftGPXFnr2TRIopd55cy2vOl5zWNW8e+qQcm5PgOODJkV1
/JHzFYyTm2edJFsenNtTsQn4Lar26TM8GPUb1UcXeqVLAyfFswN6HiHwIW79Zcz0
lyh6Edaso6GRqjp/K8A/oBPyz1FJ6CnDzB5Z9qAAAYCtZXCtzkl1sDRJpRaKjIxP
TIiQp38SO7uf2qsofaImUWcRpoaz2qDMJh5dYQT+x+gdJyJmdkIi6vxok4yGTAqr
/nPmqbH2CMwu/hG9bzvQbY0O/qoyMj1+Gu6UHPhRPtiEeaOPXewc2g2e5Jgc3bfm
FxnsUXtQiaQLc8yifnAbAq3h31EJRlpm3wPp/iMEB4DSHi2MAUqNIL7VgKUH/LUM
zIZ50t7AoWBUi5ZTfR2qwo5BtaVyH8ZjqHMks7iNSLscbqzBtcpWFIVyxW21REQJ
Z+mgYYELC+seW1qb/INsc+hvsjin1sbAOBxCerEreyY/DrQFhzZnPWEqHerRiQRN
GSgbg3XAPusza2Bmd2wJeUzTKGrwWC0fViX4AtwInrgHnaVxziF6w+Q28Gi05A2q
npXXIQaAN/dVzjkrRoCGU+ryhy6lGCe+qPHWk0o2PRnN05YJKNaSFtgfgmLR6LIF
oePN2Qmp/2SowqgcIrnUa4FvQG1hPOssqyLS4io8mEB7a8iF6Oe7sF9PtMeRS+L2
jiu4j4ME9aM6Uh1jO4sUdE+duy5WPj+bv/oSRV1i+fL2CcVKtFua7+1lXgtDoSG5
jh/nzQIKHrqnpK7HtppvsfJB+/wFmgpWN4k83RSNRsD9yzG/9P4BEU2k4XNIYVuv
WnyeD66sY6QLAJ3ZlHGT94wZnfqAaBsaj65dWcqWNv3/ijSM4Q42neIwYTsTrkyD
No0ehnVcxvns0QuUmTD9yh/NlvLRiB2J7Y9/o5TJAIGlIWPX9eXj5fwMILOHJgr5
Er6qe9otSoGuDutWhN9NlcyOPtiWWyxINuzc9vl1avBoPtGKTmOdDlFyRt3+SDOE
02FXDjgpgF2+SKfCE9O0XmoRag1xcDhTTVX/x/hfOme3Tm85PgcfR7JvV+7ltf3F
qD4++pUewv6cJ+25FhbT0wZumodBheop+2LiosdqFzJ5pLZE5e3gH1gmaem5jo/J
WPSoxk9T9VZGdcR3LZlBTfPhY8WKZQkMqkzkJQ6Rj5yaucXPszFNRh4MBRP6pgND
fdhQhNJe5SvdhQsvSyh7TzxeAodhVjXSNHjVxep9c/Z4BtH8uioTYoRuLw5QPqW1
2MNoS9WUZFgDLvBnjZxn1OTs2EVZHM6UdNFljvMkn1IgmyAz6p0pTE/xJ/GdpW4I
RZQ5wXsuQgd2Hie/6qJLMnYGvSXPnM3SMtwaAzvc1UoIEfTirug/M8vruYFeGRpV
v1EKO2I0oNHGdKZGuBqI7NPagx4kZ44O/9KmgZ4CrUKqe+ZQJ4hgkR+lk9iE2XJk
Khoi40n2NktIDdpakeqNpndwaWc4ctcR/yMHy7BHfSs+BJnqC0nKrIhY7cce4sHn
Rq7oEJ2FPpQsyr4/HP2T1g2O0JZnYAOszK+5FFJfNNl3NFdezvk4dFkBvCnC/4rn
KgLqJNvunP3OZC/W2Hcek4GdjC3sDm3iROduR3ZcS6s0xs6a+KzXwvCE3LrB++Qh
CcGmGMmInmE44Kqe8u34LMiqt+dQBMcKU4c6KlvXlFTEgqwYLDrq70ZCFUHX8jGn
TLC8pdMMRvA0MHhEWaMhZzDgMjWvA15b7WxNmpZ6v+Xq77XGppJaYx/VDODdboAa
H5yW9ShUWCcA0D6OKtGUlo72rR0Hcksvkd0UzFYDzA01uISKjzei/baMe/6jOJtv
7Vf5SX+NzY3Liy41Bx4PB8ZfgXGKnTlGS9cD3Rvx5dvsrQ7DJapc4Cpa5RhTw46X
772Sk/Eg6Xq1CLOPxC7i1dao6hVL8vmBuC9m3QANr23SdOP2coX+azQLgAD7dLcg
rAoLdkckB7lyuXafC9NUTIcTXbxXybuEw4Brl1/K1nDm+TQ4kz7n1GR6iuacPtGb
HwsuEjKOTxhGKq3MZMMksOENjB3owbCyRxqQdiskoHkHhPEWLwYg3ds6q7HVT6Wa
DWKdPs23xceMb8xn58V4nbE2YVteD5BYP3VUnpRfWddjmDdQ4ssTsaytazFN8F1c
qgJ0jR2jXNRMUC1dlAaJcGDZkFzVSey0HUYreAolRmM0YKgMaRmF1bZ6uBwepwHV
UaYtQGNLfQ/PEFYKJDTTkUEDIGJcXMKjSahOLulSUtFV1A2p2p0upcTfs7S895KA
VLWt0b0RsexIa3MdkonsMNPfaZ//amBUVEgDbGOiTW79Ha/3B/7XJW6gPvBumXPA
5crLxS0Fd/w6dyvyDrdFKhNw28Skfws90IG5hZ+C15EvjpbiSplKvs9K440E1GCl
Gh4Q9084krwUy3oc8zmz0frSFWI5UgvQXrsyrSLULoXPWQVbYGOqkd2NHmQ0w4oF
ptX2c8U1OJHBtN/thjhr2ObWqUOMIS7xUGiz18s4D6miuaBogTHNH8g8/Z/z5JEA
BpIqYQf6I2BP9yHFZ6bHd41RIjSeqRdvw2ceOt2gjlL8JhqSwJ0iKFG57eBGRK9y
Di7ygMz7bjl9/ydFwtjGTO5AXpZatjQ1Fb3ibo+5scCb2h2FD8Ao6BaAmzRIaujd
b2K/W2Wk/nAtZGD2LFjjJrHSSKKO/HNxV6ZUN9GyOceSS0xSBOv3lxhCm3zds7w7
rXANX0QcPq5i8/sKXlumDbKIy5IFe5J8hCj4lZ55q2th/ps6P3ZCb/zQzJ4KtLzU
UUoBt6X90c/FkDpkhSX+7YxwBLzLzJSwMrbJ5LEFEYJ5xx3MRWRKFrUp3m52RE5G
240ygBf2u1UfdI1d4WWsf/Ja/Tyi3gPgAotKfSYiDIYyaO8l0KRCOCc/Lzrk6Pyf
m+bQ+TGpjMqr9TEhjd7GLsVVPnGVFe8MVNDjM0gcTChFiFlJULM+Kv+wnjQM5N0w
95E8BZtJnCzR9AnDNC/skfjhTn7YMM3p9h75iXFijwSXny8yBXYmquTeeu2amKXJ
hxDBw1+XYZVPM/e7tigyjab/TEHwUWPrLC9KNWBRfx8eIC06cWo5Etq5dPpsAYg7
TgEKp2CVJqOoaTPB1kH07GAaX32vWV6kMERyjBqcWyESePS11O49n4MqytwMYjdM
i626R+n0urPClKoEwV2PVs9t0pVSWsNwwAGwlO1CfjAuFZyTH5jxPYIS3Nx7UyyE
WkG34F5gXVPg9nT9i9TjjK8cFtUeEYYWR5UuaB1I8yFOJFVm/vF398qWyc7TkMl3
gpTaUBsPupQYhEAEJPB7fykDMMN8jNSRLY9wJWrPqR3KaCijBFZWmIQTj7FCKbLa
3PUEjEI0lqdWim9Mvr5Ws+Yza9U2c23K6/rw872zjko+hZyCNuWckqy5UmIGCVnk
GBmpEq4cv1G7wiEHDKHa7tsPecjr7QTttN80wjZ8VapZYeY/UhGh5OzakFPYASAB
nZzX7xxhr+tzZESci6942VpzrnebiUjsQsvApOTQOYBWA/g1IYAdGnsLCIZ6rfym
awCRNHRZXun4nRfgYc1uoYWq5RtXHArfduG1IcVp/PnSJ4Q6bN90pRf2PJRewUSy
xdTwr7wJ3K19QDItlzGRZXNY0hTCMwEO6i0yffsDUoDmx7RYci8W+tlUL5UPgdCU
hN5ETMgn1cM5LHEz9DrLWCk0W7IQ92PkOVuYa6PjM+aix7XKgw4lJW0mr95Pe2nc
p3Qz4UMr0KLpT3xxGBtRcnqcof9rsk6As+BSlqRSQQOu9sUAz5N6fOOYeXQonIKi
1nxcxjCYujNeMuOZJsXixUBoeI8Nr74thWbCnMqkLvskeDuEGkOGVx0+ePZVFNDg
jYtOfgIutiU57xppVTtXN11V/gMYxOBWJsWGOBgVoo/PU8V0MTtbjt/UI3yuASHP
sptJzKnmU8RKF1IvhGwVQJDspwF38ZFhaJJ1syx2CXKka/4ICuaSDkEm8ZviE6eT
zBEW2FiJS13ltBm2R5llfS4ftElX/Zseekj8pcW737E2cEBkP8kXXBqC/N5x88FC
BcnM6U9iEKrrQzB/ndM71uCDS6bLVJzlCOjDE9nTr1tTic/Ukf4OdzqTCtqNYoWA
lGKASznEpiT1kmLHGpO1JhdXMFpgLv8SfiROSElnfNry5D6mDuqkajSzPG07oPmo
9wzmru75FJT1sI36Vf8oBv/I2NGrAnI2VZLHF+IF2tAG2WV9P3UzefOd+BjIJrIH
6spRW65m2XqdJ+837TapePB4usrwFg6YYFBFC7+DoFKtfsEqvrbhd2GWLaUzJnK5
/G0atgXaVIpeHztMD4cEJxLRQjxYLRv+DRjiGDc1vo4U/yXjxzXSKL2e9EedHtY/
SfsW7ybvP6cMU92pKBuNJ6M3vmlCHSvSvej2e4QHNJKTvk0GKiFtHQ009QBrsY41
lj9YiDh5RkhBB02ZdFcx0vyGNXFFfzBo0Gc93xVR5jCP9HZY9WCxNSlJ4coVnSEH
pwii10z2YiDVtC/oIkVFy33icc9OxitwMOwSMY8s12W3yL/Rf9s6L42+OBame6GN
XEwB5vjf2dkR3tYDmvrwQlMBh2QMKnz2H4CuyKn99upys0JfPCmmBQC9jaOtZ7Sb
+ea0uoqNBt5U0N5EmDHaLXn3OYmq8lFNr7jrCtaECv0J3dd2yN3j5IOOZEEsCuZZ
42SllGT4iH9a90IcSmwNR+p6bvCYaM53FxYxrltDFyMc4NNvHCA2zVwimA8yuR7W
uHv3uNYWbnkv7dJuLxWYwCkVEF/y3WZYX295fkMhWdiW6Aj0S9ftL57G9ApEnIPC
bACNe7zNMjmEDHYhblbaDqiTOwivxaXBPoqVBgSbLY0Tm5PNNSZRWrRXPax6kN53
dISg0Qmvg14H0bVB7P2Kla+ciRbeSdNHdmVyWTVataT7aYB/gIFZbI9DBnKtyHWo
xRrL+rVnjShbYqSQkykbxFaqqEscfGEpn0M+Nto2P+PNV9NaLetefsJyiETA/NLR
M2VT1Jb3BnPViyzCijrEARHbAChmtS/RFTeerSD/6tdnAENYRRWCP3eVgtj+W5xk
eWlCpjhPk8C9uTys5OkIF9+BNQ7At6LxzHeYKSfy20SudCplQd7aCrgpjWEHbdnH
yYckWXfX27XT54dAoLZn94MGXESZebhaNDgQXL81nJo+XSwOLw8Q3X2Wd8yx6g6l
MyWFrLvNLryOldEiyDH9xdMEODe/GL5WiAXSRoxRSsuTJyzYDqnRYg2q4BJHpqvZ
c7I/3D73DRQH0RprMibIopAMGI0Upicaunh/nWtUgpcXB6ypb7w6BGI2IZCWZxNu
wDUj+3HrShBBV+gy3JB5tyErBTDiZWHU9Hb7mHMkt31nF//k3M9xC/Xp09VAD2b1
2eVouqP+Y//ItQV58QYrvWA22hhMvRnn5713fy//9xcH6Nt+1KfQPOZ6uei5JW2Y
bk7mCht0aaYvsIjh0Hxb62jzF814nNACp/IaoWo34/jNm9/cKDreA1cZ4paSQXHd
PtaBDoYlGQXVW3izI/w+gi4Ws8Gy24OsbnLs2Y+Mb+AowZwD38PPRGXFR2kPLnnV
2ZpWD+eZi94FtW+Ju92T8fKfZaZ8BTKGjkb30CPyG+m2s0rhGfQVsQUtobJwW4RA
TT6Sv3ywkd4EaBoyCrAkB4lFVJsXiqk9yCmqy2UeH7qu/K4SswVOu9RwIUdtj9FI
PiMrX/iN85AZLPlHRTsFZgsAvqZRUnuFrCf66U78t+PpmqYgQ6uniEM6gndAu4aq
y9QWDjZpQk8izyxzM9j1wqwVJDgRDMft8tmUdQrd4btXUdqbiVzxU2GX/KFSrD1F
vlSu6Mzk18Gys+qpnFlO7sdigXT92KiORHCuKz5bKUmW4eiQkXyCaZRcmbTkqgbi
n7eQJD96Vqyhmwv2jgMSE8ELWYuJxmAmCCAijfsNPjISx0l/pFMb5xbOE/YslYll
6R51v06ZQKaS78AFfqPwIJi/O7+hQxNeX7MOUb67yOMcQydA3z3pn225u7NmF2f7
N63Ll4ZNr4B3iby9WS/CkP2Kb89ltJ5pK4nUmecKbb85cm37k9LSxWyrNXqg+LIZ
gGhr48VK6qumjGK0L1P6XPT4lxTA5A0klISWl6F8ZB5rXTPdKYaQz39P/0JhdjYV
zhHeatdYKLB2T3rFDhm04lnvHdYrx1LXawye4h3wlEDeAgtyLa1xKPnBcei5aOcE
eLJNNHEtydJRZx4tqATW5N5Mpb+suf0zZEoqjNK/c+iOldI4yi5k7kaYoEd1tXrl
OwXMMjF9+jC0cvoLkUMD006IrTLj+iQ5oVDDdRqBaYbokrJko5FnwuDFDNSHdOEt
uMwWNe4XsNfvZ9deviNdXAwxG8tiiNP65wqXj42A24ykHkQCKlECWSZY6TW4kR6G
TVvBnS2tN9WXopepix1PmAaxq2QU+StdbYLtq+TKRLEwSuDDVjWUZ7EHc68KEpsG
jdqYjkm56RYO001kX0TXTmSvWS7UuLiAcl06kXzaGnQ7JAGXGKuH6KPDMMg6+wFR
QAyU4Td66hbVAeztCtuF3VXL6mA/BA9g9tbbJIHLV7qSg7Ze2vBiB8h2qyd2dRL2
LcGUfFRxpvHIbagqVd+5iM62TvQ9s9wYG3JYdRO9h+3Wd/IB9u2tHUVeQImrEDFi
`pragma protect end_protected
