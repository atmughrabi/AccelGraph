// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rHMPjJDza+qFkcdQY08EzUislJdeWTkpZaVvTUeupkG+7xywVs7Dl4UkctQWGefL
XD7Gfu56Faqc9PLYXx/1Mi/sDr3TGB2Qxxg6uyCFkcoskQ0odbdA+Z6pZzsViy56
dtmzvtetlwZsw9ZPh/vthIkMGTJCW1jc0L56bfl80gQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23232)
Kw1PLZ0M0+78kl1GwyC3kw8x/EMrQ87IWa0zBuSSCSPYB4xySjf57Kzh17yZFFoI
+7Hiv4Uj7TJfefc2PbbRl8mVX1U0kqi29u7508fe67t+S0BiWUsPFu86+NKXNNmD
jxaHLmrT8NDTyeavMzx8xFeA9Oi+sdW3OwL7lahfNCeGSlX/sJUEU/NlMV65ktDU
pWNAoLKboO6JXzydW9m+sjAyB2+Md+BwGVdsd/piiJeSA8DJ+TAko/quLzFCvHK8
f8UW6OEIOnbuVS1M847ZPYJSuf53ian4X+beSr+ZDGT6/4tb9+MfS7LvN3fhGMN5
Y1+OLmWcumwEe8W/1c8UhHs74yg+I7rkewIrzD1sr+gSWUKGi5P1S2esSiZHG/sz
kGtl/2TGoLPeUawTe0PIXoHopcve39iKssaWpFb15o8WpW8qziWrMQczuARczJdi
XVuNLM02rlKuhwqoGe5oe2c/Uu3cnBFHDUQnnNH91RYruxJBWbI9cJTtSEhlwqUh
gm4zeEb70hpE16UQVeKZQrKwZb9n8UamcbuZCHR+peTCfDCViaMYiVnOa5CZE2Jq
udKykAqk6NAyWd6nq1oS+y9kB6zFS8rgAPbvxubRT54CWiSLghVKTeuW+JXHaDwL
7DwURkc+BVV+MgK5n1cZPdQ1lrhJQ18NQHfWa33RTCzwS2OWsbXP6DZ+EzCm1GX9
oxVa9B8j6F3cMyrhMoopetsAJDGufVT7STn51QA0lrsCIf+RzbmlGcdC3VeJbanX
uCRGuK+HbtGafBVYUJnYzMYev/mhyaTzkv8sz8EgZKjgevJEHC7t+zmPp5BNeVdp
Byvia4OA4Rn1Enf9bg+aJZJCgiXlWPIz0eNgxfm6NEjXBA8zgfuG5DdyZE6s540z
ilZJW1qYX97QSJERyEM9dlqgBaT+kCa6b7oP3tq2EW9QkWZeLm79Fp6Hzr9/Q/8M
9KrWuMYWbrW1Rad4JMfOvT2Mkw/C9nsmkfxp2+nGjb7d+Ud1iJUmsgZAtQ5oVGPE
c/pnL0dX/24qKkXakyy9GpGZIfiyTruYqyWAT3UdE1EQyeBcC1ibdwHZoh0QIN/e
DL3FabQK3D01FpeC3Xr2CZDhHvlOLf8YGg46rUiKCgDjyjR9jIyEHXsOqQ2A/RE6
XWmvtK56YIFP9/0icUfBXYJf0ttcXM1qBl9PSyK+SLCJGC5DW6htma/QSYLGKBYx
vJnOFZThshn+j838PD6hnqr8wUeKjsEmeX7UAwmmAPGdAKLxuc8ahbFU4vpfFOf1
BbHc8NtbBewOEbk9EdGG3lyUMIcjdg7rtuCXce4OpZEWyI7H35jGNxd/RI3glvEQ
yfoXB0R7kyBlNDVoHM1GlZT5VYTrWjaE2Wn0ERfwxDnVWn3nYRJpGW1jhfKnnjUu
2Vz45egnqgYKcm7Mc+escmS1UfSxoSV0ZduOT2CNdHikeWSQpLjhgYgo99CTFKUT
ERij/NDqb4Ap+Y+m+GUGh62OskzNUHdlgWpIaOEMO41FdRcMaQhSkOrC8ukFuMQD
MVAD9SZaT6ew7atabtphhkwb6B4Fx0FuvsBp98aqJ4+JSx5vRx6GSGhWmMKlDdlm
HCbVtJz7w0WOASC1PFESwnzlj1Oe26u2X8nPNzt+Nb1pkwRDuJYVUiTdjTlBDkcV
c6ikfRIwpGICWXaFpTFI+lNckM3icr/aj5VqMkGzyERc/hAmGw6ZKns2hMNuZEyf
JwLfwjPxGB5cILkEdzVl8g3wtyhOVONqVgLYklE/SfvNLWfF1gW1en5TB7G7erty
wxU4I2QQ/dbl72ggPUe/EhevAkMhE1bTlobPmTXyS+okulub/myTpq9G67rakzbB
jJ6uAtLZFt93ygjhYc2nZU8t00GG++c2KKdk7gZvnFPMPXE/juPcGpgJpj4BP657
PA2ff8LLtItIYN49XC5empEEF/aS7BfE2UL3J8470yjklflVrveYkZlrb2ujoh74
fhnh+HUIqqZLx1/JpoBRIH0dA6TAimd3wxbs3FuojQsRHQVO3YovgRz/1y9AlXB9
HODIVWerxJwN/wKMhuLuTj7eyrZ+5piGa3MaG8QgVNMPlGPR9tJXLuvn+LvLDY3W
bjQfGSW1Tdz5OBIQmfO667gvgXDUVA9jhS+BGHq1OhpjiW+IiCF+7QTQXpKOLNBh
JoRKZEu5DPuriqzsY3/KO4pPbsCc+RD7XQQiEDjGcTHckY4zvF/XGksDgVPgwSua
eW025yB+9p19wec6jktmx3ZG0hNCfHGOi6ApCEI80jiOKIk6mJmVVVUXDcjDz/Ag
19HY6eYcy2JGfgxKyLrztwMWn/pAmQtFk9lINlBAhIOXVBGGAQUVCUZCUufxrulC
S6s/r8rO6ySiFDFD0wiTniIUcO554RAkTGOpYUvW4heMcWv2eWC+uM5ngGlFVzTz
yefWWG1UdtvQINFLVD30ZwJAm3q3Z9IKKT0B5h0kHa50fYApTpFA1GJlCFfOouy7
qOti6TUh7AP7ELXOXW2nnYmTUVEAJLvELy27gezCR3pxdxKNDsJnqMxg55fveb7K
say21SdjHrQvsYhvjhD1ptMR3lQ+0TZnYs8NqkfocTlv1++OXDwm/dp+z9n9C37W
IlylXJRwuQXPUJHtA6sciRXCgnCROKp8Ks6CQ1NcrTqJr7dbOZM1XM25onmDqefM
j5DN3ZqnDjRxx/tKrpni3Deio+yncebCETlJxFO2Zt8ttzdpmrKkaiaeFwby/m1g
ES/BDBczDEc9qJle23bM2biSXqGpcTcrQgyylrYWRy+7E3Z+Dj5ly1jYbFrPiYD2
kMKfUwhAfQzNAuSsNmQsQo6Nla0rC+hAy1vAL55Z+0khsYOh+VeFmLB3gmSVJZmr
HVhmPUY1pH7h6r728d9krsdsNUfFnYkoWotnmWdD6qIzGtwhTtRGJf/ohedgtF4B
Jot4Wb+XuthCzEYK8o/rHIzwBBZaNoHMfk5icZ/lH43RAyFKt8vOVL/MO5UTF3FP
gQzr00PX/bHTBCRZOoqDBNLb0hVV/MbzoQ8HYK+SESoTzs06ZPbiEktQ/GNNLOrI
JUEWP7ZoolQZGomCx/QLcMZzOEEuVWs7GVbXK09lmX6fAmNUpEOOT3Yt6sduIyOE
iQoXy9jLlr3UcEhsEwJvgE/lgBXIRUiv16QiXVob01OhelQ8s/u+klVynZ9N67oM
FebYNNP4mpXpc1BlgBPzHFgnbbxvmD/4eF0sUfcfpRSfHWZ8pbK5nASejKI0dTHQ
ZW7Kz5YElrk7lquBBlcQ3kTF3QyljsJvyLqDR+php3CAHpRCdX9ZPf5r+6n+bSgO
xVP8ZTM65WZIau9slblk12vDINgxk873/dKow8e3SkzSCVa89GQU7eF/gf6WfD/Q
D6tqNLysp5zCGtXmM/H2PDGvvy5JgXqKh0wqqNpLfX1pjlfpRF9TCcnXWqtv+Gj0
q7A/tBQkr+WAeIjIUaxuT1gUKt+13gkDyGICrKpCGa1QnJVrbS2FM+L9UUrceyrQ
9QLOK3PXbInrBT0OKBH8nzYzAHiXYbYB2X9KZDw/MCSDXv+66g94SvG00wglykbq
J+o1luH3I2C71VC4xpgg1+3bcXJhsg62nZqFahWb/05kPh0zU5nFO/GGjU0pO82y
7M4mODj8UQcmvmf6UQ+b95PPLOzv1adnlwx/UpSHqsVxHrZ0hovxvjTFDaiMBjea
nR30YI53AuABlsQAk9fTROlrVYdHcZJAS95pSM4eQUkPO6GyBBGXj9Ib+EUVfHAF
o8243x/eDNCKfOchsjWz6tRE9KKQ9jNQw5JpXSUZ/DtHxURNbhXeQxLIVDNdR+Ru
9zkis2cfCrYCinsbnJgH/Wp6GGrurZR7ujWpVYhvdAl5jNVC9yEIXttPhsqROmmY
oaQI+5ptYl9M0ujP9ABF7anhdKmCBTAG3EJvxzsMIsitBJZUAGkC+ezGT+5avx7C
cFkjI7AQ+0Y7n3UtQn+JgBG4p1e5yj/PK85wFM8+So0ig8KDBU0pAfNUaaJt5nGn
hvqzDop8bzOST+c/o5a9fmzr4w22Elg8X915G8B5cOSHlaGbNhDKIdreFhCKc0Fv
/v8xKbzm41wptpYHQmL32O9DAWAtsSqjiEViQj5/BUGFLaGCzzHznMJyOhBCdxL7
cF4kynBxbjFQrVmuqM2F5UCfOfm0kR2SRkTpDUGBNOXvjw/FgUOq5rF6ugXflCwv
4x3eV+xxy/4cgN8mgW6SibVxFsTu5ShT0EO8VwXFgD5j4w9udO4LkhLaE11jXBA3
LErCcpPxf2f/2IaziSHJvTflaJmRPiXYswoTF2sctsVIk4DQou4a3umxV9dN9CSo
cggfvEVJgucHLLdpYtlzHnIIuHOjqZ4iCmN3nu4h2lvmH0xVgvMvoF30RdINPYSc
D/6jOdYr7dJo9fPD/qTHWBBs8hnNui1iCKegiyF6aLzd7xfu9RaXbioTwj7ESBWx
tqHsEj78KzPQYCt0wYvMqiOolhZfH8KPcny/VyINsJSTkAWcbmt4s5r0//Q4M6GO
qpdvHJZ2JH/arYSTPQDZNbT7iHGszOFHDQK3qvZ7tf7sBnnGhxDRYbZuzy58DfHR
iSExl0l3nIu0UG3v6HZEqL1eUJn5z9iNqQQFiRTLA0qi/LP32sOob15vWnWFxcdH
Azy5/cVx8HBVDanB0AIhQ3/+Ev/Wi1EOqreZ61kWt+wGO8eXWmhU+FOxu1P8fwaZ
trPZT5x3acGUzXBWBpytX5OALNuSwTt5BOgNK9fze+NteTxiQ4CRkESE9ajIZ2JS
RWU6jT6/fEkCYbTK/2ZXkEVV00YrSunkLX18jsN7yitGNwEvXhQfzkyn6ijm2azm
QuBib1OAz/0DCvhmMGjN8G5e792sUd39NxokUTBahfUkctWXP5h3Ha9kb5TfKFYE
2ZTyPNT1OvArct+KzDsyZhGbZFSyOW8SN9Z9FCC6MMG0miTCVEsj3HqGLNwg/EaO
2xOfdcVEahpTgt/BnwKiJGRJFjB4cvQANcNc358pJZu2Uay8PcDhIjHnSM54a0hY
S5F3G5g4K0YSvOi6qLD72CwZiW+UdFs8w/NBdUt/4LzykbTXzlUUc6kO4dWdrcyH
w6dD5V4gwGKkye3V0Ikz+/PUjVXorW3NW4C6kIH4QRZrdn7y2b/AfBvBRfYJi7cD
NmoPKJBngibGpW09KvUkjPbIWbHV3htW8UdcsWsiJnyzVFJtfndFndxHYwtRGTmG
ZjFUlbXWovo7AqogyhmpZNyx3gxRmdygHanepaHETLBD262CR9i/ku9PKSt3e1AE
pM9GbiBS+mLwoeZcbB1LxxcX28DOCsh5GvVP9qW/FXAEnoKARgGL53IJnT+rgYYB
zw+2aVahEjoNUn2D70Kfux5ePx/fkwqvLk59oH4YiPby2Xfp59Z9+sxeIlvxO7um
gxx6ocFrd/6ESo4tw0sR7x9rr4n0gG5R0buN37jgKhqIP34/4oB8MWeoU7Fqsh3t
joggs4ZnNDgTvHmnauQSlddlazN7jUtkqJUVUkw8XJq8QXDST/ZNGhRJRYBX5cvT
qddArAsCrJnBLVleeU6sygqWyBnzfEifGr5+JgUv1lnSTBGocCv9j3KxPhwwcV2c
1A4p+Hk9fWmqHaw17JF+izvSygqkA3zs46Qr1meHPQOUUVRtB5GXi74H3Ep4KyPT
agrbhe3/VN6FUY6MpcBjT1sflzm6M5vMyYcymrX76M8jDmoyc5L0KVWyMA8f+kn/
FxwQdxCF/9NtnNvMwrgqg6bDOClxZC4vZuZVrHIEZ9f3mpr6VSpQYH409nDBAlX9
y0afu1/ymBJLUH5a8KzAfz7n4Jsu5wMQZlIYRE6CV/ol2SBe2SILlw5fxStehCPb
PJZogrfiipGkvUInnq1p5IA8HD4JpOYwRuuGhSFoD4anGUmIMHOmaJ522C8JGQDE
g9jaXy90dxwpVuazK3/+VnIFkL7TAi7SXAQ1AGmmHVjSNXY0eEE6FFTnT2x/51C8
+oFqGdGAj5jZ9nzABPbbG/3Mwl9vtu+Tvp3TybBnVD3qEFOALKjD36QT5AyKFdJa
fXceaS6kv65p/lu6+c40ceTpm+SakxHXpZiTC1gm3Hp+yOVQDx6KIprAtQcmh/l5
W98vzBeqhBFe53ezt3GyQd9xnbClro2VSNDHGlLrFug1hIRmjr+L4fnKSoQ36/SX
8X942pTY6S5pH5gFsTrXsrtPwVJVUrG/tF7CP+fKqWY9jTzIX1R8r6hEgMIKAilQ
07GXFaDO6t5TwgooQ/E8wwsb2CEpNFow5yeG8YT7z12Em0X9dohazbH/9zmpWEiH
kSJOTap6FHTr1rZZwQ/2mqr9dAbGTySKLoBwwyHsXNDZ7dhD3dfmGtDXWRo2MGgL
AVOARl+p8QH1sMNY714Lv54VjIhYxYm/nJHS7RMop7kONQeR+Yt1cRbEjHAJz4yb
F0aDe6nxV+xwvbeuUE9s5txvL1H5Fd3WrC4rLQPKPnOW1INu1c8NHDNNn6lfWU7V
ckRFlC9HHEyBJG/k2ZNXLfGJBOp6nKVOWDBk3JVilMvzbBKFm0zD6DQMtN2HM2nw
AnpDncVt6l/JSJNab9fWYIMYMrJQxIRUNzhFhK3HyaM8ya5RYPONFrfQdgwItUXA
HPiBlV4XCxbjMVrrJOhmtWS6+7CwgVtjI1TE+5oiIsGslG2deDk6kO5d0futrZgG
E7rbUm771oFZF/kY4hB1n0TQXuX5RqPuBwwYrG+l1DX2a/5h73R7sv3v+V8GvLiF
FTQqOqaxV7d6tfWaMKB+nnUXh7YjtRfddt3UxNVrdKOtBJn9taK9UjHMITR7e9Fh
RE2EwO0Sspf1NkopL78zHEVRPLs9j799XuMt8kGDT21GQ0RmyuXQoEH5fdJqmHrc
L0O4im7owfjlWRRSiDYn42el4TjzAjlqOIAWTHItZbYkEeVARc7prN3JiByGzcff
/i8dukvP4C1Tsb2j/s15TRuMtzM+5+ahGgkJem6fJvI6QIKUpOJ9aCxRJMzkjF6b
nQhblh0nePie0Sjl0ap+T+RBial48sLyTbNcFJbK71OhQwkXVG1z1YcRZ4nKTwgT
0E6Qv6z7Xww6VRenBOhbvyqD66BvMNdakT/3IB8CPaT/FuCmsx2c2U92NAZ7W0yH
RxxZ0kvSXgkI7V6cVzxzsXi0y1fQxRg9GAdaYz+bMlwL6fLn5I/XxWkFdnmqMWrd
gF5FeRwHWrD/mo7do4LVarbDtJ/6vwlf/r4YMX1ZFQGrCnaDc6jIWPvHt3p/ZqJr
GlUvoVXG7ea/1X/5hSchumbJmuNKm8Rax8Z55wUWowECZ1Y/wjbluNdzPA6sWgU7
DHIwVvC5dAPnp4H7So8WffM5B5PFVN7w1IsB+2JsGOGw3TMll9zWN5/2R65ttuoU
jyOVmxf5lrx3nWadfOspBwkcG1A8wGDeYsicogpgBhvOdkts6KF5reyBbv/bh25H
e9cN/HrrJiXeopzPUrrPkY+yz0KE0JWMElAdfczFZW61u0JYm/fizgeYlsK1IR46
kDZzrgSunjtZ4vD4psc8M6VHFDwM6ASmDmswqnUMxFd97oqFAfK/A5EGag62Cb01
4d4+fRQU8uhfRnpp20qS1gXecr5raJqIoBD0ohg4bXXQL2fS5TQj5TEi2slGTNV5
Lw7ph7OFlYazDSwO1OZa0KjdAXLurFjW22SnD+VAj50ofmBHaJzlYr/S9NVADBoJ
n+2TW6oOBw0holsPxlakKDrp2aDm+7x7mGsnUl5xEV9vYmulj1SOGtF0z+nAs5A8
qM3eHifKfKW+Z0I/+/ObNUOspvrcAKThE1okHtxP2rBfXHavhStmVd6hAwcMWoyu
Mpux7UitqmWEn7wCRBce0ofKqxyUSCtzAnQJaWi1GD3dFfFYr8od5fQrlXKaAFCI
0mAP7YXxDmdU4vgfpLSULPRzAjkT6GHsurGxnTxKFAN6g23yV5E8emz2pZ2DgUII
wyFy3oZPVvpqcH/oaKcDJRjTfuVjq+dGcfDwLEywP7+aqBrg9tmaEzuL7AofnFP2
5p+PhWAx67CeU2T83Q45ap+65sCWR7bIcNBcHVT480v1God1tTl6mcgucvO9fYZ9
Guo/pCCY0ccD26H8Q/26f01hQWjQ77INuK5QY1a4p0epGj7tzeT9gMiN7YNFWVPm
4jh1uHTkoaEn10trqfY5rMRnWOjaaNWHubNSne4dBu66H+My4PAv2RWmoiQTxM9g
o5wcTd8CsltYmfZE5/lsV226py8pO0UvFj/pDptCjDkfbrnwgIFhcZZL1Ykbfhg3
cS4fBN5X74ekcg9cihn63J64Xz4F1TTJGILnFJlSO7RhE/XHGYxBxSBJwp0Ge9mm
y+H2WSpsBLtvGpS7ikMyccpYrvJyZQeKoUsaGhpLZXKZ1EN/eUut6Bwk7gIKptWc
vK4lEE3eKdGWAev5bmJ1Soh0r/UPCsCJNpswIOvdvmFFVKEyAx5fEcFemSucS0ID
A4kmJ2jmvLdCwGSTxFEvdsYAsYLrJX0I3NyhfZJvjaxbhbxJ2m45Dec6IwpXrOxT
1qvueHY0+cfDpaVWfbaR7c3/pKPHbymQiQzKl5PQUivdjLWrH5H1dPLMHTAl0Twk
xa+5BMpaNsPlsg+CYf1AOluMxPjaEkR7dPJlESxgwmbHOIifdFaam7v3IILMJAwi
ZCOHDxhq3G4aHSZyhx/iMZ5g5GYjkuqYhWr/krbB3vayLibef6b5SeFlUHJy44Xz
I7xCKtAaEY29GG7M6U3SdinejmxJF8F24vUAj52op8WUKoGDdOwM0DlCcI1CtYQh
gRDdsbRoM7RKmRtjHGP4Y4tL9R+AIdPLeR0LzyHt5HjToNteOtRMjz1DOqQ3orXI
aYdPD0cdVpW3sIMYMmWZxMmBcwPU3Xas+ZtqXruaqxh8b4GnvCk1zzdDTTdcblBp
ontugtLeX+bOYKNsCEfO/SFWWpjSR4tNIhPBxamEHYEptDEuuc6ctMV3+OVJoLLD
jXhjsbsvFR1j4HLje/UU2k3HU1hpw8oWmI3G0S+odctbKkPq3caMICsfQ3Oyfthz
VuNJh9vSor8S5ynxAcw+JmF8Qz6kGspwbmD6J2m26d5qwfvo4O9B8IUn2CPBViYF
WpDLJKxrAGjWw+9oUdffUC1tjfDAf3S7Is9KAR5Ctko0+zxcJb0T29MIUSWWSQhK
6TR1pPbHQjqO5RxKXbSeq0p1cHtJNbgYoEKSmTTL8bw1L1B+BI5NQgecfTyhjBgp
xhDslYl2e3YDAr8EDf3ziL9n4VE2QGn7DpzNqeiqtNlvh6YM3Qug66BCdfNQnpmQ
nRxKcs/4SvYporQ5+Va2aOQz45SgA68smPMlLZqa8DU35OR9TTwiQUpa+PLDu2r5
8m7mcTD6wNcyLyFytoyKTBXo/2KQ7gSiIBAAAB9Vgwa9lT9MSoLCBtkeLDa9KXaO
6WR/c8bk1mDs7lvFEhE0jvEGky83jbdONXZBg+OR0HqIgOB3SHO4RWSf4bsHDci0
0kfuxc43xvtTvk7wUZIL/GuWN94Zp/eblu0gsEi38m963TRjgpxATdBAtABec9Yy
ohz/6TWAFzJ1LNH2oMyLLNVrrZXeO/8ylnx0eS6hmG6Ll/DY5fKDSpS5B3Q6F6Dt
6mLEFJ/YS15Jj33gXxAKtPe9WYLzfQ60KUggI2c99H70YAzDwP2wYi60Wfuyl5db
elPV6am83coCpiOP+elzEmFGgF2zcOhCy+HwVRlP/M71Xg7l9ErsGP/+dhILA5X9
2+qhoP9blsmKwZ36vzyvND76y8w6eQvnP0cb/GMyOCWN6Enfdh4JmM7fIt+lK4a7
SjLkDv4tOzyYLOZdRS3N9Q+9KuGril94M0cFeypwILuNgeSWEEfBjT+nQPYG9uY6
GfvIF9spwxoyRvv9AI/BhpPwknGEvB03MK/gylNNWDgluQi+iFG//ClBpdKN4oOI
6wMRbmv16x9hyv5Vhm5SPDhmMoMLkbzctyba/T2XRcv40HEHFS/WCI6CnxothIGT
B+MeB1A4VFozbtA21zNjwfCC19hNVMpnzhpVNKw1Q+wWFHzkSbuCtgrYSUIZFFMa
ZuMpS5ploPpm0j5xPnP/0YvpTlUbXmIITYiJJwMDOJPrlSxIbZaSQLAGU8cXHsMY
wqmDiyzzBwNLRrSrfzO8HxwGp8vDJBH/TdNHSbbLTgqnex3XyQ7qj8mrstjlDLvC
8cFJXdnGic3EBKh2oCUoQ6WaeTEsNeKHAs86mJBMzwsC/Y4sDREjD3ibzYM5xMZW
rWLf6ZyY+VzHTtuyfWzMucGBw6rAQPsFGhse5DGIxCjZV2Z6ZK3jaJx39o6GhjCb
FFkdXJe6H0mM4Yk7NGJMTY/vGQi4K8rRk0HGA/LXY4o7fI9Qk96yh/XZwoygp96G
6E9Oum0scrmR9B6bE4fjxznyKSEAaSvAptHbZPTv0GLwMai2j297LLkCyed7iZf2
OCV6uunETrYCqB4L6dBTJs4ls85exmP/lvJ9yUT/W8rc5TLyyrx6wh6mad9RHw/A
eHBKg97gWFw5WSScy+MbenHcVgBwm8djhfXDvdCAqVzDfIKO44x3aq6ofVm7tCZZ
6xuyPWaqOtI+5ASVLsNMFU1p1VUJPQlp3jVphyGJln5Mk322Q3wNuBXSeVFJkcoG
62Nnf74Fu/lzthJNTwkskPRrs1amQK8Y53MOxUZzPByCoGCkOob98k4gF4oy6q/7
g84hsm8XuDB6ynk6F0wqv/o6twhan3xCNaZphxYNd6gSr8PnDHjWTCdezQvFgVw1
8uTVtI1yXq9tLPjaQLOk3BeWzfA2A/hmCx9C813eEYwjvlLOyIav4wN/+Z863m6V
gmQ+ODFREsuVnRgWFWS5NnUEL6vZDpFCOMmJdN9MguDt3eRbC4qCmkBazaQ7bJLI
uPv6Zs+fpeQvvszmLmLubFmoyJHYqhZZNdns0OSIy5Ior/f4fl1XNOkKkW0cTRSE
ZZJgzp8fXegPt370syXzdAu3zkY7Btm/WSMQaa/3bp+YJ0YlRlBA6fbaGOYGY5zk
uRO3z9uJLFjPgd9Y2qLzKylXzpjqCaSzui4FW9okFZVfOxv+XPwRa/F4VIW5ghaq
03ykYcty1goBoZlg7/ESXzfZESOzxHquWmGfAGna53kihCkewnblZ5yJgP5nVLjs
F5W3tGxbehEAK2gkUMNlJAjKoDa5FJF2+P3t6DN3K/HrNHdk89aKdOEQ/Oid96D8
pTljnI5T/QJUtIRZ/kped1wiRJJ7LCqd3fMeYZVbGngS2p2Pd3vottIzFe/4Wdyw
RNe/kO3JMFMzBuQgZVosFLXGp5kfiJt3bna/ITIu69xcFD3Mn9OSNdreuYdc3Bas
eFxJDpelpcaqkETgabmFUSoIjWTNd8af13hS6ek6R/lMsIqo0fDe2ZmcHXk8GIlE
is6LdjGQPpzXqmSmhTOSPc13heor1K6sgrR1t7oY+IhhJUw1HabCgjWswbUwn+F6
ol/IoS93djX1440jJkUtJVW3UrRpHR0xwIcY7IHHQu7pUk+GHHJeNCs4RYvDSQ76
wYAWbCtlsRIaj1yPRinUQaoN15cI6wpcvn9zgLlqFrgPqnWjN8fWQXw0YhSj2e8h
6G8oz2/rbS0OdeOCjYC0TkICMksBfGwQNgnkJQY7O3uCl9FzdSBG4nvIzd6FKurc
vLkA0KrbqLzyBu1f+pwvoCL8u6E5RnODVQglbc9DZihF9B1cfrRM7TfHLnO73gcd
wcOU28QbAd/UHib2ZTKvGg9Vi/f5wEKgNTGkA8pfGvZsbhRCVp8IOXD7w/+eo1au
dJywQcGPeCRUBNpQcBy8UlPvfg8JiR2Ot3RwXxZGvjmiKqbKkvxwF2hXWqihJf/y
Z7ayIsVRzTpHVqNoyFb9XwjKzdStpQ1WAArt8DdTTKUFs/rDWESSdKL/9G1gALj/
Pu1w4f0A7sKdm2ygurbWvEkAXkckWLGkkdV7M1ajcI0CHlrVXYUr+M+Hyhjlep4J
/BcfycHbfHNNSAP4Iml+4WcqKZ0HOM6OyBCBPyl8f0w92PiEGL0GnK3/OWUh+rzc
tsvRrN9DMISb6XFQcmsIb7kU9HPwOuNJ+85Z4+I5JjFKaxVL1aGpJ4YBMmKfEFoL
WT3lY+pkc+/zqVxPBzNdEZddDrqIA4uV5YfRCAlIh28V7a2HpOHwVK5yCBsSeKYq
bh+N8jaCbMPRYp1qbc2HqaAJaw6SWzr7BcoarsYqBqkQ5w8SicTgfCJqxzfzI2ew
Ik9oGUhhdzXWMxPR2w6wNLjIZUUMAgVyjRz7q+MlNrT2H7vqMSo8hPzziy2JENlM
vcdA8Fom0lTf/u6YKI9dNmjEflLuvDLxVKfMAub+fd7U2Y6BV6+U904+dbGSH8+U
xQgzJpJKHIdhUhTtprSBkWNNUxlYa+Vp3LZVFIam45tBQTOSig/ITFeMfk88ZrUK
+kR06rFgUXKTe5JoGYqMYE1xDACIOVGpMEGCersAwTp5sHHXaWboniZYXmHtDWM1
vIuubqMI0c0pd53WBkBt3iwL/tS1+JuN40Ydn7IacL4zu0fTOFveW5Nz4gINJF6t
etCqnEViH1PWLeqghwpToppkylh9grU9ZpFbbbIRfiZgMtYC/u44EJyLmCVW5b4d
EqoDePawBLAanoRDWkuUeC5DpVn1itGbB+53/dB40zYwjp1RrlB4ie2wLTyhw1td
dgHZoiTVUOaM6JLKQMDoypM9bLfZHKN77OXIMt3IGQecvhhVcS5DXQGl4Um6jrDn
iT94zsHkr1YgbE2oG8zrQnCVk1gKnFPa8HCXzjQj4DxqZVQ35t+bADLezgxWcz8C
QtAyeLr4WDVQkJg5RNor8v6L+pzkXgy577R7s3uPcVVs8xv+rHnQ6SJN8hQBFWYI
a73w/kNnhneCyB1Uwmv6inxqCMui0EogyuaM8Gd3mIhGHYarW8ClU7etmcCRMnwL
NfDMuTowB6Va1VNeRub/pon4mfz5tlcW3uK+EE3LhwrvYXWVtt8LcVD/V9zCiL9X
ytkCVYdWhag0b4D//9QmxZb6y+y9Dfq27UO8/9a/F8arlK9YX+SdtJ+fymIzXq/Q
jpjjimS25tU9bcCBdEWc9zO7aWJqOIMkmk79PAdFWeluLEqF96x4mxN6y8FCrlPZ
EocJIYRs0oNY4Ol2pYnQo1+or0SVMQW06zT0y0h5w1roBvy8IT9IgotqtyIxLBDF
c5tHPZMjoA5VhtCVJ9NVn81VYJm/DamHF2fg6D3oOeiW3NJ2eG1jLguORlP6zcUL
TD3qXegBiB7GiaybMr6uk9uVZLYgxUOPj4AHahbOc054B/Q3T7RNwWx7+Lphs1sy
K7XtKP4IqnEMvBn2ceGmIk0tdYtllkcCRSV20gl/LX3D6zIfctf8SQrot7/n1ePg
o6k7tMYwl876UPUDLhyEFNt/O+KOfw8JILykYcEd8j7m1KELqHacqpYLpV8wNr/4
zSg0SCc7F2L/geLIvFW/PghkPQKYXdzeo8B5b+IJ5uOo1JaDaBXsZzoPBo271BdC
iTW2HS6g/AdQLCX+QdY5REICTpuWqYSkIXxZfmmlaE0eewCZJtSVuJ5I5S1YV7Ey
0oMN8TzG7u6apqiCACUySUqox7VB8xYQ5Q69iHJNFJdIbfPAQEkLhuRMuJu4it52
FITLEGQP9pu/++XTlHpyYPaXeEZitywZdS9sPIcb2chYRYRqjmzAlYtrGH2Wp1Rq
FreygYe4VqwJFPGyqF0/J/2nxzTqg6mjDLtub5S/e2UYGOT8rdQkUzs1B1fS9v9Q
Ws+8Fp1tURq2mQupKBAlemnFVKOugVmOF0KDIknNcvr8GdSjsBSiNNNfvOxVK3eM
4KrZD0+gQMfrRkyBf1Q4S93RSn8F0/Xs1oUc+Azv6/WycsVWNemkLeFYyDUVmJMX
Yr4tGUchtRf0Ic7ld4oLMDyxsbWQUFJzr0gig8uEHQuHCXEcXllaVbFfOOJleRGt
bv5slQiIJEytgx+D88bwGwZBh8cSeI0+YsrYFRYJYs6dyo2dJBwp5uavU47/Xg37
bzqF9gJF8lu07ljhsKt6T+3Sw85dHGTK+77C8lQnm+4r0qGx+sU89cOaQEee0tj+
TyReju8fCckmjzgoUc62NoKkNEByT5L39Q7GiYGgHjK02qx0nVSWhcL4ej+pBKJQ
AgPfuj1n/wUW/jmfGlqYxZg5P++8cR1zpo4TrIu6LqinWzQ2PyZ9rZxf5rcdP8/e
TN6mJI0VMakPpxuBeTReH2VrNuUXcx96ZeqgY4VVfrc/uLaRrSYrS4iEMypZVkwP
hsn758PGkB8H9TOequuCnzZ/mFIG2JSSs9L4cjf4NHKO3PBO0hdiG7Xw2MzWEzh9
0/1BBFO9R3aVw3LpIZp2JfLDL3a/UdAACZUbzWvb6ggdUyEqHJjJQ2enV8UADdAJ
JC8lvZTKEieHPRsciHKrU5Pui/QfBukx+ra3AEjllt0r7nqNtE0Xeq1YMeG6sf+z
sZDFlWv/SCgN2GonEj3s96yzFbkZiHXMXkZ9howB0TpgwtFVz/MIsAiV26GwJPG1
P+GENmtBAEO8fR3yKwlNfCsRcd1SxiYrFMlbZ17cLwmyKKFTP/HKe9dYdp1/PEqA
yFqniiBHKUPscyyZ75TZWTOSOnDJIu2hDvlhQAnHiB4a+BiRwaFKfsNaFUSalrb6
Txfe7axBB6CtU/UAjjEas23G1Zfnsn3ZYMetAYTdJNKwbfu+89ovh8gVyaoiZ7N2
r4ZENnOG7kWIiSAVmW7VKyeLml6mY3Dt4yB9k71N8Pu149Af0K8PWWJbcrn5t7/X
wSk2UZsLi5WwiN0fnMFq3oMVYsDPmy8nwa9jRX352ciIZIh12JaOWyrBOgtJ4M08
9W+ssFwuZ7BpQAiNgdFag3Ie23QerAJvc7ITyDruGgZ7+IiRiFxIXBXh+vKpJVXL
hWPOPD3TfuvX1IOGqh4FnEMkX7DOX/rfUFcF8XqZSk5etTSJhFIk/a00plC9OmcS
q6PCLxKzLrt3DeufWIdVcAZMZo9cXq3AYUPPjt8KCKfqPlpQdp5EuD+FxEUrj98p
KYR9RlmIt+wu2rvKZSWv9aJScRtownjvUpKbt91CUppMz1N8BoD78ijEW+51aUf9
QIAWTDvjV/aygVOToE7S/oYBGjEtTLQFOzcJ7NsAJLRTdh3w2z3TNi91Ve+/jwmJ
TTPSW98m97GNltP+GAxsHfKHI6gH0vOLoetXQ/W+xUuQgUzqABeWPxSmTIeNTMes
UNFJcnVlrG90kAuJ56t30uJ5eTP1S0XIq27rg5r8LNm01mjhcUJPKuYbTmOL5vNE
kpAqgZfhhM7wI7z9QakAqFr11F0laIm7b86XMFL6Tvif6UX0wjXH3ezqE7WnT/9/
+YPfxkXV1A46RooqjOfwBG46HpC+Tjo5mmV3wxz1kxPTsSDVGVlkHeMd2KSuHzFc
GbQPXMvaJR+8WXSnJFKPWYqHa94NwxVAQ1aweAvn+4RUGXcoKArhxebrgMkw3WcI
ppZzJB4WLRanthIEP3r3VCep/gjQwUQYMpBcgsvUJmFNSkuBQHeWvKR1FYq41TQX
ezE9YJ+b4dcsrdd7hh60GgJbl+gZV7SuIABjE8UUmubNoVujqIRayfg76ZMme9Q2
GuSIjNkXS8/21+3mYphD1uG2lD2RNUrwHNZdHQ0ZXdr7v/QXA0PwCWLeNM7p64cL
Rs3WYBFDLzXaClhup3cwlSZBYOFdoT5RnmXpGu2WzPh4pLa3Zscqw82gUKtCfUl0
X/Gm7RS2v1EBVtUdgv3KUn5ovE+YaT0ZYA1z2JOtPYittnFdWfD0guT4owarqqHQ
zRGndjx4nj11ANTTdN+yw300vOR2tB4L2hh6u/961aIbUk6THCqmKlJAf8nc8HVj
Q0qr+FI5cm66wUSr5tldGRjnKoKMN0fn4muN52mcEQVWzklqyTAveiMJ18fxLsMu
VjDWJ4Ilrwpi7u5U33WsPr6vwEwCkPEp2dIN4S90tcZtAPH7PKLA+rk6eFZDB+Pq
oEQlpcpGPn3kOdAauOL3Qc+nMDeQv+09mV8LwRlDo7aKDB6gTGIshuzsZlJTLJVz
a5S+qqR7cDrVhYzQQZiSzk20tc/Tt8Y3eBlJrnptU+aU2n7HBIn4BCaKdtbhekUt
X54lYTruFn4cobIBCd3E+Un5MOGo/t1fB9HKFYNOqIEBTGPOZPSq9Mksb/iqRCWt
U3rxUtxISHZCvs6XS5sWTsQbSLlfYMzy4ABnVSXNDKyXSRju1/a/zN3LHSRReX8T
1D1f7uSVYSTtC9XVrq45Wszq5MAMb4ez1blaphsYDzH2wMZEIMmkolVqLR2TxbI1
+u/UlIPvqcSRn3kT7S3aVHbXI3uh3jiCNmg+QYn23V+nJ8VUjNQ8kNigEOUSa02c
aIuERTzo4S0d9Z01m+8kMXrK9VpMdkf4xK7gO4QzalRkvT8jK1OO6cDxyR45aX79
KpdAxGRKNj96OqVbkLqdvZmCiSsdDAni576mGgOpHb3ONeIxUym1z8m9q+UgnSdW
2W89vx3B72zXaw0uzov8y8CpT0j21VIZqOEOdBWUeHgjuntFB68679CHgqNcEdoS
wQKCf65krMWlrwtRZhfoOoLPKPZ6N3J0nrHM0yAOoKTZkJ2edGZFbAQG3P9I/CQl
24ZvXm9zktrAHWejWD7LWpRGn/HlxBqbVLEgg03oW74Zqs6a363BtllGWhvWx6l1
pf7GfhoWA+FVH870FOtbWRnPHt7NEfBE95gBIIbAvPaCKrgJu4H4gyyiRhCeol77
1JRugBGwoiWPXYT+8Cyq+DDQzdNJILOlB0AdazpLtas1TybRnZeMXkX+jZNWPbcm
Nj/abnl/qq8OoZ66H8v7fFt+ytTlW+/Vvnj/HzFEoJU7j5vW/JAcvbc7fD1Vl4Yx
+jZH1NaRyi6ZedyDO5CfSQrEukMxW1SAUjRV1qPicJsVjhCZSCvF385xg1yqZDcn
sE52IqM3ltD6wcZyksn9aCmdN0PPxXqML6P1W/WYzeXvPWfswOYpMnprx8okzobV
/u5Nr/wSfyiSEgr+28OPRdNR56LEt01lZIfAtcSImrCyyxvTOLoVOIDlllPjfUeP
TRmNPJjQ2S9PppBLVfkcjgQykaiaKdEQdcySf6x+47Yqt/x6v2joEYuIQZXezmPw
wC2+LXCDVjPhW7hDOH97pmRd8jOz/3K40KhukFQC3u3l2dsB8kgVgY9kRizElObE
wKsFDykQAuwpu1wG6Td2GTDsBsrr8AcpU0klHiKPWGRbGmC8BukRgfu0JtAk0ze7
xPLrqYPjaHREogTn+4VbefWjxEAHKFbEfI3kb7T3rAjkjcZWoxYHOIEVMcE+YmTH
FC+1habyq7Y8BRyLzgB7bXfa4cLBkZxkoazyiImEzCrtY7JGlAb6nG4eTdyf3DT3
kTNRVoeijD3s85V42MXsHEDRllzfLMkTJzssowrqmBpOxrH92VDdxlSoHUG+bKYl
spBB+fUaG0QC3GPwkEMUPWzMwAAQQ1nKZiKGRi2V43HpSaE1l0blALZPKIiA04fT
Q42sljgSob30qYxll8ODE+smNCtR85zTFNjcFgG6TAJIaTXUyzkuoMlbSkhiLwUt
nuLLkEROLi1FH7YewbkhKVoAkBI9oHsD0KXMifJTWAEic3tb5Nw1VUPKE1oyxocL
XGpuLf2QTl1A4W2mlJhHTpLYaLd7Tulof2h8QjBAhVieSI+ejD4tjwLhOSJmw/AF
ZGwXUUBrCnZeSQggA8woYRGMBjF6P7E6sfB1K5sc0jQ1ItLD9qLmBAkzMBrTW7LG
OJ6lHIvRmbY1ia51cboKy0MLi3yidQT5o3p7cZiCievXsXTRF3bbkFxuSEmi0TtV
LuczeqUQFgN75mHiFNXPyzP1BOihwRBBXaFWR8Pn9U0h7jUJeiHpTHUVrCPSyksD
lydwsSRndMt2WpyPeDzP0E2VflolHrehbQx9Vp2knLySbGHf4FHyQR5JB46NYadZ
mZ29Y+ZGxO1Cnmp4SmZioenQkZcYZz8832fBDxlvMnrSSaYnr3Zn1TggYvZUqE4L
E1xXSJwfMclwi3t+XYaU//ljVWvYrYsxmxLfLMv5BCgqToJHub/h1scYV2HsMijx
KtQXOTf+KWOa9RVCKb7OzpYidRWfFnBPNJn44RsvB28mfclJpmY1u+byMxJb8xKT
M7whm2I0k43dXIazHhrDBOrE+kJwI/kdP/jBVRZQNtEBrQxbb7uKh3A3IFffuP59
5pqUtomFgA5TYwg+yAnABxis3HD+nYBnXInezv8tU6pfG+XTI8e6AB+D7obtZpS7
Y42q4XqVtGZh9hzS3K+pRsugQ0P5+SKF+Vug6nhAYls0XZwY0AlFLTORRNC7Mm0f
ToJs9mA4y4dDRnOuX9ASRM9m6cOFVib7TRRducrACyDng92RMBkkFlpZVEIoHUZy
OfQh/p6GCzkorCSWlwMZVdMEAfSUdMzrVwYMkr3xjNY/ZgbNkbOvNMmNdbYWJcrI
WQq3xG3QAYOCEDLI5oOnS7Hcx/9zw6/B+dG1B6Jdb6fRjyQmIKUc8D2uxfX3o/MR
spZQML4yWuFXsc6dsuqduhcfSOKjFv+EsMFTn7TLkASHYI8utUcpG0Uycqq0laRk
ixj5i13b7YQqL5zBv1IMgvVJdU8kpD/N1Y+UapjGStXwylz0tpcEo9RpGhfsdEoe
33wm2P+4coXes13A9NQHcZse/GglzKdG4H3gog/sSZBffj587nC/cWlpZGXwRGvr
gR8IMXAWNKpaDbXSWrFfhyFzFXwTaER/veTdQZS7PAU4NQ9YPJHIokjpPv7ToNpX
aMUo1V5NXee1XZJ1r/+FsrhHtN8l3Kjd1LaQznkTHkKgNiJpuv8WOIy10vlszicx
+0evGiwbS3W3l47wswYKAJuS2E5fcRHFaIqXUh0POdu1K70RuAFd4GYsZyQizAx4
UusaaDz2z/jl2xtDecJVJ1qZAe1d+Vs1V8GMmsZDkMXQ50SZzglyR1Q/s1dS8a12
QyysypZxjcxmSytqAppPgoYklgaocSdJ3y2evmV8GSGHUfkYlneowt/1vGzwdfPm
XyfA6VQcj3Xt6KL91ttvdeyJAHSXav9nIoLVOt4wWudACgpNLg3friAjxL2adqJ3
n+O8sGEOn3vEeGtVm3xe3XZOc+eTYllhJ3EiAVy6nFrQW4mdBTejZBtP6nnNd9K5
M/kjYVa9BxcDy1l2ex4qbHeBv94NxXyy45cfbhdykoCAZq/fbZadX9eTBxBuiYf3
9PbvidBRO5+0b/sopw8L7Yuj88StQdJr3M9GOVK3qNcnSN8SSHhtzkZ/rvg1Lnz2
KO9jlJktjzo/Ofys2T4fGoKc4LWnmxPme0AM3cuUYkPTCgI26KEyr/9Pm5strWAX
V1RNSDsiike9s9CI3ILMn7FSAsROE38wXWEoimyrOjm4n4zXpdmZsGfbW/53gF7M
S2icS92oKbYVFMgsq7xjx/x/HhpEJTHSbcXaaqderNxNVfGOnKZGhXpgWBdpih2L
X4JzDkipKqgcUDuNYbciwGmLMsGnRaruJrhPH99OJlevN1AnrhLhE+p/MQBu04nT
YUXyIBZEaw5MmBP0J21BMO5XLX9y1MeSXRX/Ub7dSSyOld9TE5m5qFKN63/jtqJx
OMHyjPGz8lWApJf3FEQ8WMbKbbdRJWSlSoNrIvQeS+pzC4LvwomdcgaSZArqa5R2
FrN2CV8TN0DkpAMtDhTANgd0Smat0PdthmMQ6SeF6e6zPi93W0sV+9PsJWLmrOqx
3ZtAHRbcE/0DL3cz7ZLWydzi97YikAy21RvrfeCQ9fTai1/RYq4+1fb7fKbIgXwe
jasczn7QSA3fHZFUKTe6HnmCY6SmjdrddwSiRbLDPG4RiBpQhwViVu/UMTWrtQkU
PyRzKx9iFf3GPpFLh1W4Yoo3iQ32adxLgOK3fup3X8JQ1snCpSTVxa9JydspwkWI
tPkOI3cGYV/Q3mPd9jHfaQHkqXCNAwUHqlIXAOxSkTbytQNzop2PH8MCwzuv5olk
DkfEqdfInREMqlu+L5nVNsFa4kvvmRyoAQsCxwOttuLd2Umw374p/+tDkFPBAcDC
qtW23favh1ViuDyNZDmf44/hJx5c7Xv2tTFiBc2TcTOiP/EETdsMWu6nE5aGzeAe
hdewo2cBYT1SEazYFDikxVkslclvYo9iOD0rPGYGnxJqLZoYFrqzaERwV0OMmREi
PH7ObaE6y/csUhqFmE0XE3+LSz6sITWJVx3K/GRz4p7CYjK4D6LbChR4XpdujeJY
YJsWiXL2vPGcjBnW0kAJix/d2aSPKtTBMMZOutNcjR+/rNe4+qTmWdI9SNzf8rwH
85ZsSfVQMOM/WHng0zListshwya6x0ssXeyDyCNzo2P9jHiw0Ml5yVSqo1tXlJ03
1lRBjq7wkMdYABgNfG8+OtUqGm7CFgO3F1kEXZtldPXnBUmNN7k9ZUHfS7rGBuf/
YPm0eJOt94RdAnYow/gTA/KTcJs+AiaZ3UmVleZAg7LMMgu5jFpzWb7Tz/6STjH7
Giojw7ojSb1QaeZHCu+oKTZa0NlLSRdGIF5c7pC9ijMsgp9pb5K+Xr+MT5kj78X/
JnhUIfin5id1nderCawkeP7pytoOeu/s6yxlTpiXi+yR5MnRTRBjNlTmgBJm2KIE
JJ+88PlELTixB81OhXQL5bRuE8HeSK2oDUt3i9sZSfhfo1WsPqI90toSUErZXBOP
UCaCweNJM+f2FfbvCbu1CQaHWfjGOCV++4QsiscxXmTarIcOi/f/oJvGoD4gFNMU
kr0AXxO+RT0Us+D44oCJH5/H7M2UOLx0oGcJY0KdYBA98Sn0QjhVHYxHqxC9+n3F
TuGSnUfcAV/aiBo1fqgl7YBUttQBbtqKfUlqzMxuxO4IwSKEreVAdNQT2UiBhImg
twGL1Y0E2pUb5MvT5fj2Xa8/syjii1yUivW9JsgMa5p+94I38o6dWHMTz6srmpJG
WZA4XsDXnwHbbBhY/1oGmjUhVISDAFg1t8+LZCJun9/WZzAW/UB4eIn/5VIotyFU
ZjMH35NPnwT+3M0xpwr2aOu7FEqwHeTvV2mb4gyQmthrUwS2+lKlP8PFYeaLIbvT
miNU92RqiWKzrGFP6hAQP9W6cjty7wzQ2z+zsM7hf1ZWO93bymJDRGFkTT1cC44s
R4EDlUZpMwGC2slEG+V4ttk2HJEpTIUsfRYuifGTW/AZM7yrb3DQjUNLLANpHwCl
AnlsU3ovrODYz4AQMmG5hqAqjjdJz1VaDeBYsELAM8QPExkuOor1oCy0UGUcJOtD
eLrv6Lt9kRGKPFBmK6ID8q7gHeH6MJQ8JE2KzArP5EP9kvv64159BjNYoEWshOz3
l/6ISaMZJXcBnFSr4RXLc6/GtupuY6gb2XZ8AWI9ak2aj7AbdGODOgdNwTrJ/qVf
nHOz7Vv47dSXp4C2WIiq5srA3RF97GaXTonTi0YUwGSoTgjQYYQyp4ewvkgxC7iD
ByVJ99HOFQS30S9BugH8msW+5kD3ooxMEZf4q+yop5JgOHLaMKqlIe1MTQLFhz55
jGzzu83Iu8Pfus7aWtR8JorBHFDQXaCGeq9MPloaVkgQMAP7KpYdAnmqUoq0WeT4
1v/VETkQ5SshBcAmAwAds4E5FaRglq1puwPxtUMOIle5toai1HjSGDOn+mVwWyhR
5Uq7xXhqQPEMz+GdcMjSWaQmEMzLhYVqN6DM4M6O9fXP87tl5Pw5KdESoj/Wu5l7
2EunbSALYEpV3CDeaFXjUizZQrSX/MlOLGmlGYFPQCiBS9ZMEpz0SX9d8c8fg89b
jANfAnJxaWS7GXxnCUjxJ+iEG+ohKMcf/yN9NLfOJ9T4I4YKcz8lOpbjLbomPhW5
zJFKs1To2mNhgjhQPK8RB7vPNE5DVgVMkV7RPbw0lbK7hPwvYnwsrHI7nuggdRex
61/gXdvTE/Z2yh3ElcDtaVUMkrNFiupot3Oi3J+fPWXkhmduTk/GmiHg9zbZ7z8y
alAVg37EIkaZt6/Xk64edaz5mr8ZFzobJm26GqHyDpDL729bkifItXXtEV0CKp9t
7OkD+fFU3IPHwNfVp+9wBeiP+5hUT8KFcdlIwuWwkRX8vDBCZv/iVuk3QhEdPwIZ
FhqnWPnF0vc6TdIEUvdU2mu+EfOyf46HHp8X7vPbYXfl0vPRIfsdQNC2pXB3r2xx
+0nLdaRZ+wumVnrQauXKPp5j5INUJyI4xqVBi5rshZ6b03Pe4QDSJpIT3gZOU5Fz
8s0p4ysN4QlHQnl9HFGTKIz4HbU3J/J5rWhf/P5m3dfGXnN96d0Hz0IRjwN/Fyeo
FwHLJXu6DWF18fYLR9jhStRFclaGke3oai57ilPHx0HYdATE6b+V1JzXzkYUwCu6
MoGgbHBwe3tVih0SiuoZeBwQEFlR9LEa7DV4vNrcGEWkBIxZFRYnsUmJUTeNXGYm
M298TSUncA8tB9hYcf+qTELMprZ0fDrVHMHBZqDaJh+WjcUhR4v5GvHuDCNeVrbG
sVAgBygg9ojtj4q+yRaIBSlcZ+zVKJyWl4dAp3zDwbg7w7Kw5BKCH1agfEy0LGOc
c9j4moKvtzgysFjZweib1ejH5RWZQT5iTwf8ku+V2fN2qIUdaebp+IqfVGv55Kg5
IbfbkoOtt4AKx36By0W6Ayuuvu9RrquqxoU61e0AjyZmny2a+rRJBjeR+d34Q37l
hKuKJmPqRH9jeZz09bbfV9Y7YfakaQeiAkTm7FUqK4UINlzEU4SY1Lp8z+HxnIA6
wSTJTSSFtbF/vCatJipgymC29eDghFUYzxTGHFH+OQhBw9tzsOSA3zyqUAvLIttm
HIzEvprvUHVAMhDbayT8pMfr5yf351vLhiAj/d5BmON3WtKyNzwHdrqSnkNot1iD
RhGU/Gb7nKaCy71gHHHOJhhJ6vH3Qc5xWOpjAY7WMseqMJYB4WlIiiX6EKLPr1P6
VF15q+T07zn9VZJyteYv+x1OY1oJBuUC66XN9DgJIv4pDqNo1v2JFKYCqvz+cMKg
DjF1Q/SOH2YbidsRPbC4lP7Kxs+0zJuKiNP5FcZuzjHwWjMwPYu9VeCoOrqourPN
jYfSKQjpH5Ggt225nQEa7vx5d7NQz3YpyO3STCB8tHPOPZw9URDORkPsUza/V0ah
QrIE99aTuu3Y9vfjmvqmiaD7Gi/mV0reYvI5qOYWcf58Szg14QDw+TwQpP5WsIni
jTm5neLZ3oDbJpbOauNzO7tqhdUHsFTLog5cfWnsyI6mwyC9LVdUG7N2NHoCCgFb
g37wctSg53TS/fNAwJAjzxSApUv9pNGY+hYB1+a+QIbsDnPtoKU4YVSaw50A58ne
aM+9v1fpcq8ZR1NzkYrjmVZuQauDFSfdKWGhx9ZwEqkvc6gWVh+sUlF30YdhzT2P
ZJ1fCUvAtoSfEG5ELY/wrlCCdp2h4WSNXaKY38y1Br742kZ1AAZ3rsNPY9TehcYg
Jv5+8QmBf1zyD7dBKLuro4LZpaS9LIOBd41MQ4XM284Qm38cKxkmPwrVUJF0aMJu
a76ejtQEScrQmW4wJSfJkxZrxMLjw2/AB5qYZLtuqN1HvornnRTN2tcEDsMqBivz
7UZwvld1zaro3DzlA0tDdFoQ+216KFMsau/1y9qk+7D6sqmv+oFsfKIJ5ckbhk9O
3oi/Tml16mLxjtDT8/1eKjo7qaEzNIXjye+2nw7AW5gfKW8xjVOwwG1uLV4BKyb9
Vb/pmYJ52xrVoBgl113btCUPrw/RBKNvuwy78HVDLDa8ulHFNEc2SU+5KcXVlH26
0VczvaxdcwSRxiPH+jDdOUf/9scSllK91Y5jr+t2CNrnFSNBWz2yH6Xf8EExBNgF
5HyNcGPpNkNJzRlw63kdbfqQ9ZK7kBfPHdQjMQ6CrbBzTQK4L56ZtS8lPlNcLR69
5kCV0tjRcgeBrpODzlvMm6N3sjRTUZi3IbBJba2QpW1jEkj/9HP8XxeJyJLALrNU
VAG1k+ni+laSBRYzJcfGdQG+LmTQMnyX0YON/xMHwJDIKiUQtNUAyxAMBJagyDdY
fVMPETkc2CIYcECEGF+9Gvs0P9EXZP7697io70qy5Z6jhDD1nJD8ltyd1STGIDuG
Bk1XCxD6Yer1rJYq+5NV2O0KBfPCkcTLg/9U69WWH2FYEYIK1ijPU61lgBGYZgo1
WD+V0d/KHZXRVfv5JaWJy3+43zgWQsQGh48YVV0idbRxTPprKqkGHJRC+SfsU7dR
wohkJT9BiulJDdUcRnlycDdXYf9yTRcbprl3gg+LVqPPh84iQpvKNgB9VRRARJVf
H/zsRM1J52EAgazPeFeMy8avm502km+9r73l4/aiefbQoRaB3Odmlq1+E6w0tvJL
Nnxa8bNemHt9JD0HWRJ+/vBb6YbN/bGn0vw6m9TPPvCU2y9f12+WgreZSHq5u1Bo
28ZyDsHCojB3dgrUNU9BRylfanO+Jlk0ehuMtPiVuVyXpu8HxhO4EJWEDHgYOhrG
hCgUzhczZ5RRSPLk5rPMkZHWvp6Ken4Afg+afjlGg+QvW9BlLPXYGKYg7cAPT7oX
Z5izdXINLr7T0oaTBfyNwTrCVrgQP5D0RfHDmWXwdaULmuJPS4OMS2lbQnKnsNuL
b1d/FVP13xKFkFeCQjVM16G9/aDRyxAwbgNpjIIFeTBBdaT6P1a2XOD8jHaEs9Yq
qdvl83fJFbpbC5WW0taJ7lvwu3ka2XBifqhnty5qeu+5Rxp9EmQiuWOZungj36OD
L2SlQbgazb/Iywjw7sDq3qxbu+3FqI/BtuW5l2kxFLxQMuarvZFbTvIetWig0b4t
umvrOH3AL1pW68h2dx5kYE9Jz5sQlbLoiPwU6xc4KDnqjBlJ9D4VbycqKrK96QhO
4ow09IYMmJLPE0AbCK+XPNLwi4evfw4/z0g+0lLz3ITBFv3GNEmc53CUk/9LtwD1
j4XKxb+GkRYowl69rtoXEAZI4ndRO0xMOFhfEACbRTpEhjqgkfo3ACUGYJJr46BB
AAZy/df82IZqVDdwRxzRzzN+2oEhTbHP/z3UvtO3eO9v8M9sHtu/h+1x/x7sFPlA
zZ0lFF9LtyXFut6tvHF0++l787R0l3xi6cySNUKTQwF8ShSwDEeNrBqStVwlkTnq
p0Kp0fx5E0py8PJw6ffd1uuc08DayR+U8Zb2h4dRYcSdFWR2ynTh5i8XtAeYoEmK
EEWfOY3GcKxdlkj0QJ6J4loIwXntrGNCy2dxEtGeEx++W2yjHAN99Urc9pJn2aUB
HNk4Hr0QXOBOy4ASAIRBOqp3cnERymXLO6MYn2e+t95I8Qjcx30Kz+2XJ18zbhJi
NJNVPlRKA9a8+H9lmZBRiiyZ8/gr0iyOZGeI+mW6OkKISZcazKNdrnC439DDC8ks
igSpk1R75G5OU38zwZOnHlxXRt2QkTTFW3k3dJUM/CQUMA9sn4U1Lin1SmTsTBlv
DoNgZQl+exiRgAPIGIcALTbFUyuLYG8ZWn4GMqwD5KlJGOqUU/J8f25YI4FkQMrs
r1ALFpom0x3x2N18j/fD/TSUA8aumXdJfDMg+dnvA2EuPtAT2ivjcpBSfbucb+u5
C2Yfe+nBDUjYwdd6qJUUwvh8nuDvZ5hfqK1Rkac2aopUi4Z6smxYYCZXDCIMvuik
OjKqfAVHU9PUIQUWMo43gbPaWqd4xoPEnaxWZQ6RefcilYSwkI5+S/yAOZWt1rgH
VqZ7XtGUeT5lOXwrys5LG6ab8dVLz9+oE16PBxCLR6GenaRX3imt5+5meOOAlLa7
34PB82mUBFp+Uwj4HDiJjVt4xhxSSvvztPcF6LHVHLz1qFWjdSJ2fpv6XyfHo/T/
62jrX0CJP/0FHaie0iFqpb7Z4GU7/2k3CfvXPFGC+nCZqbHm2G9J0ve50rP4VZll
4+4bZG3oILnnt3BFZnnruPb3h9iLh+VnJpvLzeyobvctqCx89y256oSvx/bYBlxV
h+atdmOtsutlHHvNzoArVl+87Ev6+v0t6zKcEV6tsq+CfXEmSAkEYTGFNKJ3/p/r
5HgU8DBHHJIj2ZU2PiWsk5RVtMn17gYa32aPhqW3DJN+uUuYliyLrYND0bh6hJwk
aM6XygIotYtsuYVwgUhXxmu7nCvCNLmaX9tjxK4qzZqRSyqpigVShbtl8zxYfO46
cmfAILXVBEjEqyivIMdyZfWe5L1xLljB8yaYthn7zcb4VlHBW9enNhClT16A6qHs
tW+DkiBVClXLX7Om48m+KP5r+x637QXhIF3SIKsKjnPMFy3qyWD46nRqNzjGSawn
o5BtC/oaC/1pYKyqm53LoxUxyOvMJZ8tPelkmWxF+v8ddR1IIwXwj89hw31KKdhq
0T5LAN4HGPBTP1pAmWANg3B7Iyl4YDVRbN+gbcDvw5duMgRCz9/UwyZzPDsQHoER
r0TMfxZa+uFo1v5ymtmEJpMcj/qDzLoAMjZmeQB2EWf4yu1mApz8RRMmRREs3k5l
kMO5VkOCEvyKRhASMeFVDyv7GNkRjZvaB0wkKr6d+teJ1pWdCySj0ST9SQG2eti8
rBGsVfjJfgfGKQ8mIFlLVXyScO2vsyx9GgnDTYMONQ6RJrTNaNWQ1WIJ3rwS9Tgv
MOsSbDHES2M/7QqjtXpCgDFi45RWlfpWBf1whb0DGTKmFXMCRQ95us1dFaCQS1Ql
TELRRHJsm0l93b+xFngnqzmLy7D8aJuZkj2okV0dntIVMuMfGaNYSRHqVBFDKQCv
w00snoRCrP5Y8lDzZD41hxiuf/Z5SwL0GC3szSzxTLyQbgfCq42boTJ0rrX3S1bF
nMJ7m3is91UiG9417XmaCMBpQVMUNa06roBdvrxpPgSIDsdPO38GajzoLlaBYIE/
bT5M65NeL9UjAFN27mH+CNGGVwIo0CyoBCq6EXOaAujtT/s7TQ/iIX1HqWMrBr4O
1YbUJ7u4tytdkIbjFgQQrBy2vJdRYOPzfXmrKIma1VVNfUu1G/iSwLGJpptJzSm/
hT1vTg1iQkHZxlwMWTqAi5TwG1HzQU9taSd92nycGU/rOWv5Zp8bg5oXNfNhlEgu
aMoVjaWXg3k5c0tURhw73FuG6I7tdZtnrTMupkvIX0ukOZE72Ot4/UrB5IonAI+o
cxUUWCKtOcvN3dZxz2c+7VupyrUd+qmL6YQr40wsQBXhHKffpxwyGkO8j2wSNRnA
IdwrNz7MNyC3RFmSaQYKBO3y04euepC+vImF4YJvuD/DftDayL3wuJDrhzu++hvw
3s3IYIns4pKoIn9hrE/hYGCDCbDq4Un2w7DfGCGxpX7fwTbFfdUsXdMnbExYWOn0
mERA7BZoRhsiF3gxpsVV415T0U8rGO8aHvoQeDIStVzd6a3G6kQ/WhhKAf6SfwQL
5rGkB7nJfYFJQIlhqNo0muCS875rx2gIJBxbLZscDfSQ4Y9uqqTCbG1PCmYshTgz
O1Qa0x/lYtuy/vnot7uLkc/x7gc7i42Vu7n3j9ehBBSirle9asMZViSoxINRL4cC
sB7BltoJV/d70pE3uMa5wiXS/xUm0epQXZVToUpTTNhaU47uq9B1zpPuV62YwoTy
oou3b2pBc8Z7ef+wHxDx1H1HjIAYPNg0rCxb7zrxfVtDH1Kw50zE+oczOlHKc+3b
fqxWrvuCX0Rmz8oqbmkj9tXjQn/3xpJSB+ln/t7PdhQo1Ac2R+XqETm8Rd//iWMp
3x0LMD1rUCHlxztCYyG3ZjW1MIKvq5pirAnh03XKTLstGjGZ9bgNWhTFlJSxqe2L
Ybd4sK0JFNSPiR+ri0zpEzJHXbpyZtM6TGZTJDKjuYoSkW7XEcg1fCSQ1hGwLO/N
4QS8Oy0fEZ/Vt7cwlfAy9EMZqqC5Y/ZZHEtwYvHAV3xZcSBpyqrdnTYGljQ3eP3i
7acJo79Nw/+91q2jnTTu98Rzyt7+D9TQSyNsPQc5rIWfeaPKKWSKFVJDL3JYiLNF
OPkBmpU9W3bH48OWCs8ogAkYDeH2CcbvpM/hwvPaKrAP3puUZduKlw+Jf8zQpr+j
wQgZkW5sWtNpe61SoD3istCzDaregdTLPy9H+rSe1WWTxxlNfeoN5uoFYI1yDzjQ
SDAASc3lGC+D7zVc0JdFDQbArIysK7NrQWgEFVHzyzfLOtGQcFg88Y0eXvWLyE16
1Q2KjMjIp3hhYOxVVEhaskAaaDg5WvHmKwZo/BsUEJ0OuMgF0S/WQtn24nEqChmy
W10snl7b8fH3fpqKVZxVrXIR3MGCwrw+HnY8gPaIhTMx3IgLGSAQKQ7W9layE9Vi
Hcpt9+mwO0b0dSUXOgN1R+lIMComMMXUNpcFC/ySrC7FloJC/nZ22Xp4GCkmx98w
iJ4/kbXkENmmSDOMeL23Don3gDKKMAj1NIdRCZFfnNclW90sexrF4SMcIQTAMoWO
WfFmJofBqeorpqknTxP0IFgGUpSGhwZR0p9RWd/WZI8LDL+8T8aY/lx2Ijzl059b
QvXtE5oydf/tFFCJ+JgkmqRFethBge5iFO8v/YweHrEv28NjO/a19r4RVJZlbm9m
fGk94iylOo9LrpNtzlwmHyryobUiVo6mIDRkKOHRAn3wpVNYgTncoCK6jiE29ZKh
u2Nly8IZelgwnta/10Al9UyXJJJbsBk9w8yJLSv/UYmYGogvojqXm3ey5AzLvoTw
wiPl423WuYOOb57EQGdOFxhvKfGqBZNwuBXKxfiTS3guVuI1YSLiGNh6c7lWGIPd
8VsktRO3WmLuzAt9zc6F+xwRC8MDdVXa51Vm7sEMoHcjSXMmmMwJKwX63hr/P2Fp
b0jQIM4soDCy8exTZZbA7QZ3N7oLDBuKfXoDixjegdUzXLyojyK7W6NTqIDO3J5s
+YNCI6GTI4u+/ICNMzFkXus2lFJ/HPYWbeUhNlhlezgMGMfos3RlVFu8KB38BRGe
98/irF3yII9bi4TBC8Bj/wMLJfLVRnpZBL5S6dDzcdCGRljo7nX9fWqCrYlZ2nDt
eG8BoijJfdg3xZ0mvqFYRls6bZIeUgzfBynRS8kiDGpvGMgmH9emzhYCCwrfmN5X
AxAOWcAFcXh2nGIZnpd8wFAY3+vZ2gES/k8Xgb1H8lq1d+Vxe+gnp6eZ10h9dtIg
39T5YVfGlvMmNWkXXmuFDBLo0DNtp371L8dMN5CCP5vGi3fiucm4VYc2RSHoR8JD
9Tiwfq76OhNRqfHlMxY9EupRsrgmvQDAiZW8MLCUYX/4sPmoY1CWNXODhgJ45g84
MjKICUPGJVOKZtlBJHOl44wg/vGz9Nu5aoxq4cNq5djUOTt5g1FpG0/3bhBTKZH/
H28CpJ8Cl1qtsq2FCNFcBVRxKARIwLpvXSNkZEWydoa8jnP795hD05YkyPixyHOl
By9y1XiBkPbw9XVTyggb4TBKBhnJRqpoZxKaCsxvuDNaRHO0en5pNWBG7yWz4sTD
17H/dEqJ6V+GlKZd9XDs9q6VPDeYwm0GlPwcU9fypd2RcZyh/uzs0CZGFhRd9Z7r
A98jH7TdOpQz01JVvHAfd+d/brcrUDAZnczmXpwj+i7THT7uAW8FUw/+BD8ixJpI
TPjg6MyCxxS4Y4MO1ygjLIjuFNUlQK9QAJIj0TPbVxl/yXFj49W5XxPPDyu9OM8S
HRRxhgGJ7U1wJIodiovGp2apGGoJ2YuD2iACPCLfp14VAehkRMOHpfoa8HzuoG9V
uvQtxHrwfOSE9hs6GNp9zlwG76Fc36dV0lJ+0nin0xEU2Tccn306R/P2+uSf+ByL
0Syp858DgvTzNXzFBams9CCHQ1q6NUdinmpUckTUwqVli2QgsUIZFLN9OzrmqbDL
IWHNabg8Omqae/TX+8j02AQHcyE3CJYRvbzpevDDVEg+VeFDDJrdbZb5yPDTmT/O
ujyP4J/quM4QlQ23utDN1K+6GxR04RXXipydXrYVrv1b7SG11IPRSy0PpDIzGgVl
urejWJeqWm1Yp6SL2XNp46zAFE053GHvD8spIhP+yLa68T7lM4iT4YIbc8B11b72
wCERfmu4S6nJqukepJ68RyQ4t1VW9ozdnqIslRDJJB/OY2dfTy4ewHTehgotImpx
ZzKhs/yah6YSg/Dcax1PhJy37YlVTu4xJ8Mie0BaHW8Eu7gD10pAiY8uAl6rAOgW
2XjmW/LcLI+ELoSz2UtpaGSNFuvJ+fe+8EJKO3pDAAgmntbnNcKadx1rIcD9zheP
QgCDz62hNtEE4STH/SnE0EbWMX5BvCsBtEet/nVTNcL/Uvz0smu1a8SS7gY8IjLv
nOv3rur3UjxwXA1Pr9Tns5WFDy0BBRfxxNNWKjFY8UkqWt2GLKU+elL50Tk7Ct1B
f2xfHKMuk8dhH3eDxQokAPoa6Lz2sl+hgpSD2NPsswRLdweHywCqM7RbwohALGcj
xdCjt4/gozllV/5EQBJ1KsASbRuecIs49ugas/R72Ov4t1ZQ1AMb3c9S4n62kHT+
i96eoj+z6n/NDeOPHb9NWpOz0M964Vu0j8Zm7XRhr1MkK5izfAJz0GO7nhJvG0fz
lqqzwXLpHdzlvFb53KeXfDhKPTWfOK6ftDTXaU28rHP3Q+CX0zBAPAB2BoJQvCeB
lWWHXs0ixrhhKEWYuzKtj29eLUBaOpRdVa98TpavYbmNudvavLUrCsdqvMeOjTwL
hfscD2QueqQSRycNlcrzyRMXbqrH4t2sPVv9U309x7eudXLioTsnjJP5DD9W9BaC
uwbgmsExnTHRF6T1bOsgnraCQuxBKbDoq4qYbQVzQIAfM68vnHTbprxrptlJxGAL
DHduvpqUWh88HjI6cc8PvJdMUB1NjF/95eKcNn1dshQWoRbVHLS/TPeqhkfvHda6
9XtSarhllKKhfWN3YNYGW5DxGAe3CbpEkmo7qF58jVNWSo7ibyPHlF3G1vge/Ex5
`pragma protect end_protected
