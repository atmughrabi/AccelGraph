// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:45 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CFGLojE4goamgcg1TIFP6P3CBEYVCl6aIswUHsja1A1A8zcLkPS5BA1IN64pncjN
DOR5Y0rbkeu+pTZilfX3CJZ0LMRH7EoS47F4zHG8svuAp3agLX+RLssNOsyMqc73
OLrb83KnnRP4GpJyu4HPwVTY++DRToJoHKeufo5apCo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5664)
NTejFdGKlqvgVxLZgJWYiDNnjm21yIa4KdRC4BWep4lBQxD7K96KhSns9JDtlTpA
/5pmDZB4PLASc7Cvqv6Rll79Dx6QDMJ97qPkTLEJhObLmiL5i6bVatIyxSvjlcCd
siu+TZ1Y2wortg3tv1g6lpMZ+VWdpbq1aGrQGPVT86j26l1An+BPKXByQUOf2u4i
AKi0DwHSla67aLB3WI9M0Fwbo41qq3gY5qV02B6/F1y8wXzJcxXh7ZS6GkMz1ioN
ShlEO2G0CTG8LuNYwuVn/+nl5AtO7rVTD7fOxgfyA8w/S8lJXK+d4j5b4KNULcWn
ST7bR2NPH42Chbs0bH1VHWz/6prGlm+YhWIc5XG41e8HaZvt1pvRr7QFRlT4wBft
7cM8hjajzCeb0Cb3rQioLdstabxTaRPvYEtEHcvxmT3B8qght1UqcHdyHqITVl4p
oZP+Bp1XxTzc+TnPRlFxM+Te+0P/nZ8cy53iwl+MQnE9Gy2h5/VuCMGpuArvsUiv
lhDXqgNhWZMmtxgiOisPYh21G+LLSL9b0Z1EoJWXJZjKFDMfsJfGAO+uENQUncxj
tQwLXPcnbC7sflsDCf995l35rPgj60EvdokTt0JmiPlfz09j1Agfcz/AoyD1ySAj
9PaO93HpLlqNivJ7VkuvLTfYMR8NHCAwRSQ5ksaAg/WfUmSlLFybeaiH389+jV9c
J39ppZRxqF44+Kiu7nT4hSexL7u9IooGsOj4fz8R2AmGgBNSHiLOKi33ohEcf0uy
I9nlmybizwwFoIRYpfnYGlzkIz/eVBFyseqkkgkt3tfKf4IqDvSUz3qpSxbpWFXS
YZrg0XraZEG5heTdLnmr9AoN3L1Sqxyftz5dlZ76C9zKK7Z/ADH26WyVKB5HP0ni
UD8+wMV34N4OwLVMgokQDi0Y0j+EeoaF7N44T7INBKsrXnjoS9Yfv7q9xJGwuZie
Jt1p/lDvcvzw60JViXYVng1MbynC7leAiDs1gENWK8vHC/MkRiwLWveORb6UxSPF
9GJ5lyYxu2htw5siiMNhPd/jshDsD/XkRJ50qq5feuU4CQH1cHzlPh/a8lIqieT9
oAKUTufr8yBTSdE7w0IpT66EJdRSSg8jqNFzEyzrcnJizVjDdgYWFRFT9/ex7G6C
DTQxiaGgLCEtgGamx9uWarAkViqtY2gtKOS+QsgnBO/BG94J90mI8/vUqRtdtcM5
SGL+OBmLQbLcg+1d8mJ7Y5j/N0F7wiyRLzECUUgPK3FgP4auwyYafMe3xaXSpOxT
xuZLfoftQqiO6cAMyKL4SmdX1Tmgr737/Mj/b1/NnAD4hj0AZ6/BvZBhhoomTtO7
ivTotAZmUcZ4MKTlODxXORM6Gbfpz0LHwrR+IngdR9vAp1U4z0TqBGvxgGI+A68f
Dr77Poaz7zaaV4ctpvhfsOYeIU2+f2HTUX5kTtqEkX3V3dTPi9RCI6/WOJISpqTs
u0QOjIyiDqYGyP4bXfOZzTmqaXkmx91kFCHqNmrgAlAWkd550oV5w7wqpW3PaPrC
HQZF3Q5TH0pqQ9lwfzltAsy+m9X+3uKC8P26LuMxWK7zyY4xaCH0be1aRw7EdTRe
mC2sAjrS+q9uDyKmRRFu5FspxJV0JiezakhhnqVACQLFQB+OzylfIpdeYkrbaEBO
2rOCIot8DPfG9VSKORXWSVacen5eVQO2YmN0nQpRRa47ZMy4u69Zgs652OEYsrpR
nETmz7WOUGOWf0iCE79IWeY21ZZhS/ykbFwwTqOTvNXETBxoaAxoE8O9Zr+tceNi
6r1wrnKcvQvIkt9aC5y+n36Z9nyDlxHEW9l7MeqvGQmNWyG5dAr8+pEzqFesDGjw
S9H8Zkft9Xm7QShiHfKI3nlN8AVyCsIqFgF2WOcewNkgirDT6zWQ5cT7dYREkMni
UHEwl5LO9U4Wk/u/xQzQk8PFeJj+0ZnewT+H+vl0Xoxtsi0PCz0I+n8M6aKR9Gvi
1O/1gmX1cxc8XaITV/nJjNf0N5+Qp/GmRNLDl38F+NU3xRAOxPz784zVr4yJSUs9
VxwxpOaU2NQcCh8Dk3sVSNgAjY1X66J3vQP0agsfte+smMB4Ya0IJJ0gNOO8Bt2i
7ZUj+akpl9H40ovxvHNuptpmvJ0F5EIhvspA7Ibon/+DgyjzUUAsOMm95x+HjmT2
KRohrmW4wlt0oDs84Y9ETr9n+f9fkSbNiW63LUquPO/IOfU9oF3xSNddKiIU+WpJ
qBOf3TdK2/4rXclewUGMIdwbkdWxKI3wyOX/Qkb3IaDgj/BE7iMKKj6Y5uxyeTMY
Oy5FKxMGQQ5WlyLv+IlZF6MQkDkBpxyRWmT+RMaGnRvNetTU+8XDkpL3Xb4X+uQO
bA4wyh/zHfh8n2KnH8dbWLhuzJYIujsiwGFlo7Vt29ZXv5ebJQqM4MHcK2ANYQfo
+p0HMZERzlHoItQClZ3tm7hpCktftFgGZPqKudoCkXNMEOw83VZze92CW7pk0mBH
mO1tukZfzyraLPhqXXWZcIkokT10uyuJhsq5sQ3vfB1wkIoXLr+MkYVRfEVyuRET
ryDgz4vSAU1b7felu7yV/eHDKhI6LHHQc8opNYB65M7b6JjX2FW9L1NX6CeflOiR
VB0elxcFrUXKgs3XowXQSS8njD5IRnwdF4bJy342QrviZNjrmZ2tirnTVl0Pk33Y
XUOQ6s0sl7dIexlCQseap2LuuosjV0xYGrhAkfjvMD9TuslFTMq0/CqIua+LZYIb
NmY7UNvSwsQ43Lgklng0i2QXe0egQFj1YDxwN54Ch5pGlzmXdXlGLqSZ5opfSu2v
9HMRGBoi58Cb/ldTiJxQotANkVRNzd7HNhYVmr1gNEMyLYVFMsmLNlHqd1tjTSb9
HrrGVJNZWR8oUMXnXyvu+9aDypL++2RlfWDaTniui6M4ShK23VhNCFfqoM4fvqd2
FeyezKjF4krX2lvlG73QZ0HI4e1arJRfm2yPgEubnz7/Btfsw2SZYL6kXFTDXg8Z
lznaKQtZDBqpUb+tQslvX2uTMyXOF/Yjg3Bv2QG/ZMK/Yz/IFZQFclCzde8mEzjU
dNwTFVfwlMDFkuFxkEeKC2+XP0+FF9xctr4f58M1lB/xSjNqScXiUgUdqOVNu0dM
ZQ2HGYre+JpGv5PnCynMJVIIQZUi8tHP9D/6nWNhvJfim/CX+H667yeojNoMzGkM
q1Gga/SJcAmvrj7W1yMJgG6npGjQx8EeaCL2PpGjWZROxDSob08tQmwzCQi71dYy
eXXnD9bvDRNPAtRy7q8BH6Gfb23GVRpEFtLdDUDlLqoxxn5goEt1H7/flQ4cKEZN
Zb23WXO+CvA5/T3tt2mtqQT4bbSw+tbw1hmif5tCU9u7uPt36tgvPHQelearHE5p
cVzsWCzLFTzhN47YFvEZWUytfi4+PI0MlzBZiPKsjkiPM3kxgW8/hKzNVtcATgFG
TplAv3Qskk2/qjEndyJDQOnQ2mUi5oqY6ZTrpPIhQ50J1RsPWnoicczDDSyh2DvH
ysnpJ0ps/FxDHggS+k6heR00izOFO6gtMVPzw2E2NFpqZKtW9PIDk7Zf4+jwXURb
x3HiH2y/72D6Cs3y8IvkKCbegz93KUnk1BebhKvn+jWRKd2JErY0FIrzbLbz8kMa
LPJLuf28zma717Owm+ttUcDxmqc7Jm4soEc58Lx6KrBlQljdwFBgSiaz4OZYMCOT
AJSEHl9DDid3NcO3iSzyKcuu7QKx2kfDoi9zEFOBVF/Aq+cRFKFU3E4FCtNT/ND8
77ImfEhX4slKG3fapBgkF/VnhdZZd9X1GgA3Q8obatQjEETr92eWmbBEpKXznrpS
XzwgjkV8kh/n2CzH5KFiujw9Xvig+iUexYis72vn+p0ADtY+8kW6VZLbHj/J/lQ6
qlkq+FggeAQZe8dG9Dc4g67C7/wk0epL7LBXvFCtgp9CKNgYlCQdfcIceJN4ook6
kYQ3IyMNZGI3lHBEmsEl6NJEACom9k9873bFs+R7qmYEWymLmSqQXhyZOYmNI1Yl
EJATSgQ/tWuaCpF5OeZi9HTyEUm9UDGgFBL8zOXVGFoHW2f4HJTYLLAtP21EMQd3
FHyvXYwG8q77SQ67W+0UzVca8BhsOFrru8v9pf0G28a7F4yMBOkmT/+2OWT0vmWF
mqrYGAlpSfM9cG+kccsLq/rWxZhO8drXO6E2LJxp1oqKhVZ1BIqEwxlNbZORiVTH
uIyxoj2pUMpjxjcEEKSOOfRy3KAIa6vP7PQvHhONQ4POmH0dN7icDl3IKUpmBUO4
ESAdNus4CGNkAudHaqeiRwC1RbF/ScE6JPGEh1cTrxHisNYAkpAg7+8/9mUD3OM+
+bz8BZ5KrbJjkJMGNvCvzEV3bodzR2TmpRR1Iq3luWOEYEf1eTfZSkXO03Es8g07
Q73rsPDULjoRlkXkrKbyG9yRoPbsXT5KFzfWSg22BsGjkmInAuifjA4p8Fb7yWQf
QRUx9Bk4f6sYmB/pQSxbCHGRdgRd/6wsfT//NcTvCiXM38yth5X1lDqSI4H3+l67
vafeTxedOkoUKRuKI3RhC4rKxm4bb6QINrVHG4LlR3H09VgzxcB9QOxY5J6lPne0
zJfsHh0o0YvLFG92NLbzxdXWl3BDuz5LitulQeekmVym+x3FcfKdcw+G2gptmey2
cvCjZxMSebj+foKl2CvXKTRf5nWIPFk5Nxj37JTxSYs0Gs5q2FQn0CMWYauoKzgQ
8G2uYGDoAuiQzS2zt6554AFELL5rEas+9rut2pE7kf4oGWxjCKHUbwHyFhAwoZZk
HHfMNA34VntHpb0BcfI7oPhv9XDbl1To8b4bZnGWO6tnurwpvDbi2OYmMCGiasIR
ITZz4BT83qw8RbJ6aL/6f27NnRQFidcqwfZhzxvum7llkX7iHzay28NMeHig/EkB
SlCkxI3Q1w394ksG/N/vAUR6j+Sz9SUc0ubPDIBW8YXL3LobCawj4iIPFQHFDVEv
8Xe6YyYZcvtvmifhrcWfIOKbs5hoCSMQeYN9hj2EOh89+sef2VS0mDQrjtRPryu/
/D1keUkPZOIfqOiQI6ubvaFf8MhGguyYhO5qVf3V16eFDZvZ/UBHs0GSovUNAEr9
71Rugw1cRXf1lA5rBy8P8VzuSXPzHXQ4AILckB9GULBVbjHj5dgYtfb3RJpWH/Ym
KPDwAJ8cHWnidL63+LHT4vI0Y5+hEAD1kM+C3ycmJe8x4T0gx4hCnbfHQ2M7ROIU
eW1e+AVYas43rUmCTwbuTqtwQqYaocQ5R3xf8yQpEAevBFimO4cdXdORHrLoXDmZ
D3BRQ/sUQlcqm4SHkXyBVDeqhxU8EGz8Kz3rNibJ9nufdAwhZMG3fXouIRiyECY5
knexOZ4ejHX4GHCjN0NT2WVIRCZR6Py1X0whEyTi1IlPBiVuFmsw/OB8MKM2iGUp
PZhlfvAscNaumizBtnoBDFWlD39FBZhVv1AJmw7YNEXzOcY1FPg0G4wm/K9Fm64D
jUoxYt5XZAp8ejlwzcddccYL43FRGjQz4zFp/VZXT5C9l5reuzqjftkFX3guaWkI
RO2YsHyXruC3z6HHe7r086n2ymRWFV0pxwt1P8OA9UPFjB2ZoEPLMzrzddPUSl/q
dB5O6tvdv7dHHx35SpACsEgiJLrEBe/khKnEQqF6kJzmBGzfb5qlam1ZbHPM2G0o
GXcWJVTI+nbhCTiAeeKiHkwFaDws3akyFR2ZSwxlgHA9JSXlRY34tvPmLXFY7lCy
apwY6SLD0QYYCKJBZemza+sGgxI7xHFSc8lh/6DcVcyiUVd9zlAMKx/slyJtXGj4
J1lN8KjM+fH9sVk5TOglgW0soCWC1zQvkBEpsrJJ7xynvdAlIPR8Y2ybWywoUtTl
68Shnp4RRl171Fn8CPM8efpegi7ma2UJbQSKLn86MMt+gEE6jtAdSom1Dvq6b/Hv
bw433earN6fiGkHCZgwi07I0ZFoufh0fjsxjOTcL6/eMn+tWFzKtQk8ViBOQ1Q7S
l3cRpgyOUq0ricq5771ggkCXshLF7O1sIM38Ep5Sycf3psCuuemV+iEOV/+Phqy1
krtXHzagrHqu1MI5FBQ64SaS+w4Q52fDsvqQnbHrO0ZnK9AEBw0t5n1ExMMpsRzs
I0T9E8jewo5zYKlvzKF6+ANYzQNunsv1boaaNVtaniH6MUwQyps2y3djsQt1UmFH
4ZEGuEZvhyIyGRXJwiisIr8faKPctPt1oxJ+5rRT1cROQ10l/+TbUO4rymLPEhgZ
++RFOQ6MsIN6IrU76VhonyYvwxLb6QRyN1TSPgQZ6fmd2Km9+Uj86kimxxeRTDSq
GX8uXRkqhhz103MLt1rsI87vUWtlT8sjafg3KrWUThST/mDwpdtb18IB7eGruNS0
IJXUYI33ivgDqOkSErvihVoTCf05H4kFzkC9FEZp5TwR9hn6ipuqv/vk4QF8nNZA
dqBj1BS82VYBi/NSRopzqXf/rrFgWiZkTITPbtlceNipHZ2AxOgmLmjWjzDbzoK0
myoW2pWnflWPP6/tC5AQ1z/rFZadPuuR7JdvcTeAsJDkGmBjlUyi6ZWaY3Z0QBMI
U+zt1Lmkp290xgerA1R9l/ATNU5C7XwgNG1KAjZd6kzg8H9b+WL3cfDw1g3kH5yp
44fTLxPZXlyBYXeA1vxuMYsOPzIakGAYrmBY4ZsbXOogBCD4LFZrPHr53pFMjFH1
rg1mUegrVHaiIncRxcNX7FpjP46ESGz6cudjq8lFdNE4mi7hkitT9PswnMadplmG
sqzI9SCEilN636rUUEwEsrmbV8dBnvASTwoWOCZX+MLS7lkvA3duGZegsuRmvff2
X5EMK7czGB+ioeuv+9srswkF+VuSdfuBUZ2ZXeXO6qXxuopb6t1p3KI/qv8oGbve
9ysdFsEFLExUUWdhZJb6gf4WzueXeLF3Nrm+tvDvrl2R11MJpmYNmMOvWnZ8Jx0c
aBs4ftFrNbqiCw1065GxbjNUMq9+7mTi/0tBKWCQ02bOPnAmHFLKDx+DIO+KHkGs
/2taCTChFElAQ0mJbeOaVZyDblRTrH6PmbtV7d/GGkIBy6r7D+7FsFMm2iavbOTi
i81YPq6yBidWkXaZUB69zu1DCyuGNC9o08sStLWlEMU2x23Y8DW8RREwF2n1CXg/
TfJ2PAoqb2jQFRdRSkKTHZ9lmOQnJUp8lgknacGXbWn3dc1yutubTctk3ZGC4rqS
tyrYfhFihxgbNMAi+57xxLN3cXAIP61iFtYQfqtldUtmYRwoDK/AMsdGZ4/vtWFq
VWsLILrdtmCVeND/MXqX3tILB8sCKHHooS6CXATmdQmhaOsOaklZvw0ocVfn/I39
1AXT7su1IgLZ3KGDz+XQ/t6T8rjZ6Xo0wOc2ebGgfskU0Tycr4jX/2cT3MU3pUvp
ZqjSbpyqJF4LkH5GfgJYsnSd1j1k0Gg73V7yGzvtp7/fDophbB62vXDP2DZrXTmR
Ul2JbHp9lxHK/kAkQTkwn2h6giZSpHNVN+OtgPcfFjzMFlBoy7EuX5kleQblnKAT
`pragma protect end_protected
