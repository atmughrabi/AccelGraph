// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BTHriWTisFmwg6avfGUak1Ef6DymeQINyhhTYk5HVXiCayrm71M+jnjzQfOjt8NP
WhD+AZ81IqqMzxo5KINEVu7R1hwUHACzUR4UFDKSe6edU0elhf//HDMZLlLV2s5N
taS5VoSwGOoIHOqQ4QPFkEtYUYD+qblGfnLg6+RyxJY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3232)
X7wFijqdXJZDtC2OzI8e3HctHHH7nJJW+37HTC3lVffLdz79BBwAMa4EKS8OwPmq
+yv69sO756ouuLmZkuInScww6Rud3yivvKUp/rr/gLnlWjyBQx+09MLIobIyHrck
BTLZew90U3BRUb/9LRdChhs9Xc4h4y1Qr+NOstzHkIG31av8GzUSDtQds6Xj1aec
paDUL/k8Rc2zPofWrw57fn6pyC5fePovOb2H6wObqhUDRzZzSyL+l1tMZdmQnOVY
HeS4lkCVZYXEfwTPYHYFqExWtSGGLIRS0GTbxZM+q0ODIc8mRDZpotf9Mz0rwRhg
nzQMSnl4Z/VAZqWIFVICaGZyACQqy7XBfytDz62UEUUDw9gj9Q29gE6/i/n50I0C
BKZtaPFp0Xj/Pa/cMJhoVRigF26Dtlfsxt5D1SZAhoQFp+mJBT5EcP40dxZBdWIG
cVZvPMdA+IAJywZH/vdzIUQ9kTIasM9EKsbDyjmcJhow99C4OUFB2QSiMhTgaeQo
z+DWeI+k8bIvAXbozznHxo42oq4HGMXiKQMYcQnVoOdwMonaEr5Ry3nCyt8MwFHy
/dzoiaCzyspEnb31pXld7qGmFEvilo+odwtnjttT+q/Dw0u5F4tDf37K0gYuwC8B
Woobap8PBYgi7jSECKiWaFwp7ssGHPzoabhlM/AIt7C3Mpqp4HUz98inJf2a1w/J
zUCLAvR5+4kAyMikYzp4gEsNzWLxRkFm+KdEWtJFNXPyx8c1/6MHIKh++6RO4STh
TIloQ3lKUmd/nNaOVupBlI5q0hcChn3x2MjAZTOZ6653pIC28HNGpV3S/w23pXmI
DLMXoIZVkYK9yZCKtD5E7DCqLNhOVw4sBHzdQpCPHrBz54uMT7TLeyxnKE5xpjHQ
yCDyU5px1z3Pwb962BUOuPTcRn2YcIKiJgRsL2+9kqTcBpJaFqoweSopVPSP4EFe
kwPQo7fGlEO0ibGHnQAUxcCJvF3JcFCFIcqQdGqYMpV7hVOFSTJy3MdXEfcl13gM
0xVcq38pszHfu8EvVRoOk9Cch8ZgPfFtwZHuGOG++0cgW1yClPwLHhemy3bzX+04
pwJmMQVoZTyl5V11a+erfAd4GirZfH6yB15PCe8ujXj4n8DEqINiXcDoLBZUl7V5
XcMryBeotMeIX3Qe6wzrKLb7569R8k6rzkpegv6p4CvsuqiI6VnW0Lk5/7i5PS0h
U4FCZMHFSihFiR4c19RSmyAop8mSxLO0gWMzPbaY+ODZd8n9zFTMXOiq7xpbI1YT
SpupF/udsEEDKPlBl0s4t9QVMC+cJreK8bgPyW0UMKkzgbrPplszKp3GwtOfMk3d
GTX+qBq5NeGYsO9Y7m+kOLpSAqmh6AMODJcjIEYSaYPWy5XjR+hKdT21GAHeLUS2
OHCvLa5SGYtz0KnJ51moN+XfOfZOnFvIDpGW4mzKcrtQZSHpp69vBAvZIcv9HHGw
ArGVhC002ju6mHipACVgSjrcGKBEmG5Xbbn7Vw0vkrOXXfQOc/VjVJ0UNlrFjSji
QEP50ha1QXjCSloJ2XwlqNh2HKSdjwmKuIlFV1d0Fj8aWREdTXDtLPHeidmJa9/5
l1LmvWTXAg3Aj6LwuranAOHk6ks/oVmDan1ImhuIv+wD8MZ0G0eSCB45VeJVydqg
Ez2hTDtThhjf5drMdWNVnqqD+8W1lvw3BYbem6FZw5YMCnwc38IcwWLEOwTneDLk
i42KUm+gm2usPe1aYh6+cOoIwJXbEeE9F0CeomW+qA126fFCIKdDKNG8PZtcSuWC
WSw34KG0zeE83nGzRi/yMqvZVYnjeDI7hmcsxw8Z1bHMCs8knw0lWhDS4cABNuZh
IrNFtXZ//H9xicwHQmBb5pG7r+sZzt9lKPcfi6gemaHL4gUR6yfGwP/rWLyMG80g
9Oliqr3lgxfACpUQQsPC4Rd0XCFAbOVx6P8vLJCrEXxhxu60/ZWVpbvAj/2p00BY
OdS/BCuts6fSOKsXZCKqKqVX38c8pcJpwM3bnHD9k3RJUdo9FyK0IynIgVIX0Elh
5h4alT9NlIhdpHQUYvLdbyHxBvUmxzSnXjc7l0p1W26l5nN5YNqcwfU90lNLpRdw
9MXhlUV4Maj/hdX3hCSrP1EOiCRBN8sfXbUjsM9Q7HXIeFkNwr7Y7D0otRCuhJJH
xgtns9qkhCFYfJIuujd/hWi53TLcILmoJyaiKu8pqRgM52gSekvRZF9aLZZHxm3Z
JxgaxXs9fBY/EhIHnKH4rwDXjQQyPExYfI6j6AouQ9wDhdhcGqBI6JPNJg759M23
w8sbOZisb6RUvScVZfDPP18TJMGoPGRO3/S50yQj5SsUnuU0gARCU5XXgaaLLvcb
luhLoE9Q+AXzWuCj84kxzVgpSwJ3pw4LiuJbw4fT4UrCuFbUF0jhv5igvyzBpPU6
EKolLVjGNqp5RQCE+/QGFOuWn/eAaC2oKKoQUUADyIv0Ea3PzP0168Xs8/Bxjgwc
M72VAzSb4t8swZEOW7Lo9J8eP0ww6EBdxpK7zq768U0mnJevzWfPcTJ+DJw44ESz
CMkFzsj69pCc/xorG9bqk9IutVhYXIhWjwlQjjDMw5uNjhL+l2OVkRuI9GKwFUQx
D/OVmcl+1ZG2Dp1njJEbN5P0wdzgRt23qCJT8GBdFQYztoz/xSw+gg5ly3OYVDPg
IM/d+/SJ/dekojefXh0cWYBTGiqBmZ0IDw+XZJTcxsRCAWTvH1MEaGXdWeZj+v+j
0SYOUmrCPOaiRxn4yiZRSTQQmbnDZjamL1fN1hCIdGy24RUn9ONO0UN9+OeZQQ+Z
Oum14pm+Gw2MNvBQxhoN9aRvMPty4gnSB6aTgs8mKq66DXV39Ud0mXi/neh/pICO
njeC0gHry1vG7JCwAE9iwgcUT6WAIStEfefvN0/rGW7HwmBbT4UolX0+M+mF59gM
h8+ex7CNujeO3QwLEFSSloTlK5XvY3j8tDTE8w60l0oqqJ4o/AHTjd+lIzgBRbAl
C0kp2GgMGSyrLK7k4kWY8OCCGFMLKcAPVy7zZeyu3iU3+Y4Exy8bVITcvPeJ/iWA
wVbj8e+0AgMQPJGK1uAJAFUeBNmn6CdTNXSQN1cWIEmMb3bCt1Q5oQ77UicQ8E7s
qEEZi1lr63rgQ/Nk2iM60aLDvstqI0ML5yTG453hBqQwwGds4opmQn9akOqecy4L
1TFFCEcwAFlXTYi/uo4Hh52n2WDOZvtYT5Ef2rjr9P286gP4jkPXqNW4NdUFLumL
iAx+pNE07JSHLgq8SESmRPgN6o9Ml0KPUdBYFf3qpjL7tV+BCHXilGXk6TSO5rNU
p13JOQPKp5ux5qa9GRz4rl7+C/gIy16JIYbF/MbRxJAK1Ni/AJ9LM5C6h+o6Vcc6
baKsoJVFThCsr1Sb5KBJa1VQtnqgS0iUCgXQMTTN9vkiSQSNRZF/mlv0DXq6gqF9
KY80hVqkiytGAG3Se+yxMPb4IExT8wzLEg+L3NOaX2UM9bGW2KSU1cBKzbYMMAUl
zWiP9IW+QgMqq++JXmGYK9fPI8kXcd9tqViwKOwyz+pBpA+6a7k5eeHRB6Q+vdUK
sLT6DRq0I4B0n9y8KCxcjrNk7VnMkzAFaycI7iExl3u7IjAR5xpPk7OdzQW0U9um
zD3m66DZnICz5UPzggoUOiORfoLF18/tfT5Z+kpO14/Zn8ja+ULTu0yABO5yEvf0
H0ijxUl1fmjsXe8wHPVZK80Z6vib/yalNUaZ4NQ38+/I3PR6EyiMZN9mIPWAoGIo
IJOUZuMl9VXSSW1cZcgv6QuKzrtmtjZKNO9XVk6hbLGUVPxdyR9hSCRyOAKrezN0
A3hgTEPHfcxyKJYH0GxZkE0f9skBMmEJwpboBh4KnecNVbPP/AugcBp88Op+VwNG
hF2TbX0cUr3C409J4YMKCBEtOjB5TVB2ruAsxsiKQi75gHp2IcSNUitEio5fm0pz
8+l58qsl3OVarJkiYarYj/GSNzWXtMe02tDT6ePc2N/h0q72FdnOHLrsU0sRl3XE
gAVvByfh/QfSXcee4xDOB7H8Jf+knOyu0ObjAc6VJKv62xrGaPKLnNPMLxBi1OeZ
ZRWz/QlFnaPnX2SeKRTj090fuPChZYDaGvviP9Qf0eeRomxxcvgKeCQQftZzxPZu
HI5m6G4c5kE9DOttgATzZJsKilycJEKDWxXZ2YJzAFgxqDdJ8Y7Wadoow5jLYkSv
yT8+AZWV3sDHJ4lE24veoj9zSMpHE18anuVrwQOOuMwU1j6BuQu/Y0lE4ec+xxcN
sOrskDnEzk8Xx7nlnF4AWQ==
`pragma protect end_protected
