// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
heF3UiryKgTjSmYfdXRnxRDUc5ITr2TYbeiIwOKYhGptOOlsBROyzSW+giH7t0N0
279t+LJLgY5NfB5m+r+ZV8SV84oz3S9ZsFsses/Fu/Mt2y0ZXA1HLCdhJ4I1x53W
vJF+04h6QhXPpiJCH4GJ4X4UUCSMFm4HKvP/IUYDT/Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5632)
IBfi+5NeuIhaERyiS6Hhav6PSLfUyxGMaxU0nhG/h4s75eaK2FSpoKtIKdKpWno8
8EHj4fz+90q3Z26eBmS/DiPWVdQeeG1fZ+tpW1EiazwQ5VSnMMT/gB8c0dAlfTPp
mr7EmZmysVBdqM4x3otIz7dQiYGYl9aUSJ1R06JFfnSheVcS9H5qRetBtKQA6E2t
CqaaOsfqgM6Cp5UBId+7vooVUBkUk3PWXj/8wY/a9Asg+WshuTb9i5gFB7owcHmF
oB/VIcYnuHXF6xrPsY96FK5Av0tNOnz9JSw5F3IOH2w61z/NjcTz79uk24R7pMQq
94JFIY3+6wYpcYIZjmKrv+DYZdXPWg+UFnDS+9sywOiDL/ieJTtcKEOloi7XIEnJ
4AzkKKsyWRQZ2lJBl05TTKz+XZosAd3+y2SkyatukIWx0993jtdA1samtCtuUuOO
FKTBF9O3gen01bKaqC57sV7e6sdhcvwTywSnzP1wR7FWWNMVnScWfoEp67p4MdUD
h1RU8oM+FyLsaYn0liWxVVc4gRCAXXctoiiJc1eTzUo/UdyVgCq5Eff+pAeCwqJ6
S5y9FphCXuk+6OUTno21QumzG2Wo3R7iuf63EAbsTsvBek25z9tR86hspNCTNSKB
PyzmSiR9Q/2xlMEQ/q+L+kWkByMoFmYut5EeFQGjZ/vL0q79imNBa5il6Cd0sw2L
hipEiL5s9XOOGmDJn14xSzlBKuF48WLQgxtDmklsSkf9B9KjqeitLP3VavKbJAAz
XV0iIgTWrQYle1WCNszWMvWwh86XveFqglOIeJW2PdhNAdSwhlE3I6ZWtXARxdi7
pe8YMUkrjGuI7+2o8SVjkHrnoUpg8eegK67uyvT+fRlQHKgVJYJ+HM7dZnIwhhUz
3a7HJD75GBNO1kbVP0gTpQhhp/dCFRzYtu2rH4Y2Cih5ItFCdjAH3ysEv0WT40Cf
IpbrQF7kRLa8K5SSfdj8R3iJovjM8UPheIpRigMXENn8pqmpqjyraUePhypSiHo9
APnREVfLwpvUfZKYzKM7ROj1CEFE8tEyAwtc1JwaMgPJYUYsV/2UX8hV7IbUZt1s
FfxtNPp82QY6aGwlOF3hfBBOtbA0TWV+099MlOtGvG+VbKBXge0E8JlPajPfy8WW
FzU18IBrqYdtGFNwvEbkIWMjyq9kI8EHvn3MD8Noa7RVxw9DFWwYuzjAE2MsQAzU
lMZxu37TSTNbmTBwXFMmMr+S3vhUoig0nd0cWq23o1Yb6ixtOPxq51D3ZsI82vM0
VHzTRyzx2DXTS6zyri82psfZ4q8fvEGpCKfkkO6nQ42NctubLnxvtDr+4M3gIumo
KnNeNjLcbWgC8J+boibKciGf3tJU++23qmRTGgbxQeA6rg8RDYKv0mycsFDK6RGk
n37pA3uhgl3KqQfoo+0JfqIZGjuFClwPinj4kem0RjhiE/zncRrScXwnUl77USo7
9uSOuphfecNaNOcbctK6gb1BbagPWX+DLKh6rMMWtDc9177DiljVglp1IG3aa/j+
+qqb4eEaW8i389QrYAP/OgdmVtEreC4HbdrRi7LASA5JbfBizIbXQbIi/BblTUWg
6N6R2kTfBF803yr8Q1+qNbAWOFlePHww3WUGhxBPo32OtKe4/Jc65bYERNrtbpY9
1f+bXZXJG4yLArwr6WhvjElgT8ZdHa0A0dPmbNJAvoTS6t6FMWOX7/YcUyvpaFfB
r3lpLQu5M7MGC4WidY9coriNMKy+KrMKw6FYL/ndGsMQ7Q+Eg7ezjaATVr9rBJuR
jv0b/oDxmZ/O8bsmcP4PKifP2Q+Eo40YH3YjUJqeISSLcVXHVOAd0l7b3YDvKNwD
hBKZzNpCji621Hd30ED1envaTFxZ9H8AYt1+41VRDfe5xqt2jlKyWq5VIhWHSqIq
TYWqjbEnzzXyYFybN/kaLzjnsNgBTzgXR89cKaA7FCe//WASz71JwXWG1Jz+K3xw
ud8MRuFN4UAHSOtlYBLanJua83WOxiqez/SpV7utWcJSjlVNB9mAnoetio98hYR1
OiOfePWL1N8S1hyvYYFq+VXNY1GkU8v6Q/SrXpovcQbPNcuvt1TjaplytaNWzqMi
ok+xuVjzUOHM4xbofZ+7JtppuJdkNUst8SDGlUYdAoCLhyMUTffn4o+LJSUdfOC0
qabFD3eCqVydnAws8BiTHfjqyHOiTmCTxW6PHKaRixNxMTX9+xx0IbvOIJSPQqFy
8g4BkO6jlT/GPchAzLa/xunBKjiQwKqV3EyxZHrdUyB9DUJHbe6eK303J4TfK39u
h6PzNCt2Q6u9YJKj83WbYVQYt7OB4saBJVso58E8XfIB4ppJOjSBMDYTRESp93BK
PK0VJyqy9PnwMkU5M4tcCi/knWzOZRCKG27YhXDqukICjMZ2220QOT4/l0LANhCS
oe1LYQo1dcCXgHBwmc/3YYnW4EmGB/Jov+u8tH7FNQlwP5OiVX4Q8VUMe81gGnKj
CwlNOLs+NoTlIQ8Lh3s78zWp/3j4Wz8KQx637ZT22M4gyXVE44C1hMdcuUqEtJIu
YsJbpc2TCfLBXh9ZTIwhySwcDCrEb2XaxQvpVImYJnKCDThu1tDqTy1DA1U576G3
A23c7J1rChVqlDgrOUucaJieZRtc2HlmprCrXpRA8Aj9f2pU+Ru832B9Cz6NEjQ7
yBd1pCtIEwxRxjOr6BI7Wxe15IfNlf7L/BY6QyhuzrB03JIiWq84ugrxYm0ygL23
IAG9Yd/a8MTQLyKrlB64UVMMRlKkNmqM0/mrRIQxBAxFIZ3BU9rhQRCFgRCHqZ/j
4nYohScRpuMfU/Ylseddl7HjjhDkMnie1REoupacaOTPKbNNtDEPU81lVhKyHreX
fozWrbnbBm1ULx4PB8rv5GnKmD5P59aY0rcmKixCZjnTVCijcWFtTkM13RoCNHtE
Vyeh1p0EpWtO/ce5yzk9Qn7Q2KTHJpb9zD06CMn1wSkWSMT1uCwIgEJDWEqeX7gK
BLKCMXRBuzhVvLGeQBHzpXC2AgKMNsHBptIcGvhNXV9EPHswhppHkP60bNuc4YL8
W+sXoKu8FIpgaSpVknCtkO849LlDUavKEHt4NqNUb4nN6CfPp5A7AKHwtrjHW0XY
IOfXc1TyJ2pD2b7qWvWaA9GsxIYn7UmUtKILYQsvVH12YMx9vjvYmWZeeU5IIf95
JarwO4LSqJs7oF+KRVniKRrKwwhl2a8fa8ulVqNlo36EbsuvQLYCMkZlYsZDoy2r
AAtMSRNflTd/OprDN0QsEAaeSYGlPl1KBmDfnIgRfmO7H36h1yDhxLYOZ3yUapq/
Q/G5nzg7rVjp7m4BANlhD0XJjXSroexDeXFAXI6TOfy9LdddctnH9LfD6N5J5AAm
RGqCyjJHkQmIODu32r9l2DHWdYGpTa30v+Vl9KawNxDAgc99cmUaiYwh/ifwhrar
b5AbKXoSASc+i4ycFtfZCg7V7PxubBQ0fatMsjoyuShuT7rRCmmI78d2nIsjcGkL
KVPmO4G6B1YEyJJN/yKmASd64IIN18Lhw2A8ZORlGdaPf0uFJ+sk2WtZGbF8t8v4
DIQAmtV8fzRt7eYhDoxhtlp6khcha+IbnfZYDYVdqElntmpVta7bCjLioFgzdKYU
kwqWNr5+kiJaa7A4X6mq4zIsWst+m2r3fgSIxEXvRtrRhO0Yjw7evpTbRPWMYjPk
Fj4wRGowT8yf8eRWcIVW8SJ0Cp+RAPS3ZWLwd0JTZU9K/vjpVQAbmRbjKqmROtlj
+esMyaRwX/pHR/a/i8UA4p9fF3SOokcBRoawTEoc2pnIf/xSAonrKV+Ugdt/hktY
ykYH6XLryFByFuCTvnODrA3WOWDKvOXsnYfsxdWwLHbYbi8uk5jOJDZNWuyAeihj
cztIXno5Aw1l8Wf+RC6HjBHR3IMSGR4V9Y3a8DP7cjRNZh5QOBHIXwvFDMZJYDOm
v7ILfJj47CvBLy7TfP+n5IpLkOlA7akmc3IrWL9s84O/Yl870F7hZF9cb+Q9HJLz
neWVKHZzlSYeFnrmfzGZWFcpgyDxLFPPEFDRxls/RaEAlJuHAZ+8YHjOkZ9XhwIy
Orzw/AL7adG3NkozKpTDVQnvAyxJMyreFA2w3VWqLn2bptJc6GQlw6gYXvjy2yfL
wZIyvDAPCHUmBpQZsIym790yZtJo+FnsCGZDRgeD3oj8TixGnvsX7k5ArPVzYgtd
psUMSuxKfs5eo8M4QGMIjOHoMEB5HLAbVcRic1dJ9trpE2Qmn42clLXhSSmy/dvS
aeKm0+FH1qZnrj16Ljatpu09wkafJTn5OQl8ya5TK/zXq/isnlshY6fl0BW0z92J
6/5zFNOZmk2lF1hhkyMJ31nviGHeAoMithENnvB6Y5y9mSeboYkGzc2TrCyQYTng
2lc+0YhmimHvHe9unQWAEHwc0NxBRjlfejgluyOWGMJ8SDlLcC9uAhNUmFXgQc3O
G1tvNgxS1QVO/oTiq/dqn9PpfxfvF1Px7we1N5bnazM9/q/0m6WctgAHIt0cG6Sk
sBzN2jRHL9MjHIn+7G1ctSE1FcmV7XSwmgmDFk6UV3GG1vmpMX5xH/pof3hOBgqe
N6r/ds3v3nyAu4vX8pjc3ArP+2gdrNAbYw59jFCGpmS86ye3UA+ed4RFIY0nniPU
5mJ56zqdPMuojS+GlQV6CnAhHMvUAG+ErqQYrRYIaEljMLspXRMaWlkJTLHL8xwX
Ny2zRH6NJLoOuRq29dgK6v//3Hx+UFYUvMSLqbRyIL9907ZhA8OCsX1e3/Y2Q3YO
zhxTlPN2aUThSX5aDQYtLgJRR6tzGlPGIHdMgs2/5z6pkZaM1VrwGPBHJn7ZkjnA
hD6d7rxkF8DTb4Z1/SKfe5hYdW+zcTdtvH1PMGhZmF4tzY4nASRTag9IwVH/zkz9
9wjl+nikJSjL0z7DpGooRE4yX6805bQsiKuPYWgJqRpwWGthswlh/efjZ5qBi9A4
Ss/6jaayVySPfn2NoM/+Luq0E1QUgKBDnQhrI1LgzhPQa7v0s4KwSP+1IQd+zj9R
7ykMM3zvR9k1TDH0DW8Ckk6Rq3/v5wvLS15J/Errw/90jcbtUeAqTUWGNuZ4H6+q
IxWooPJOCzP8+MmVm+F20bqcSiqg08WUes+Cy5MsuKV/zWhwbVt7MzzTOXfRnLj/
R/ourndFUKLAbHHHViMh813IiTCvupE+EEZ9uELpFNw2xBumQ8EzSX3j4bqXrQDe
Yr2FFjfYoDZG3tlERuUnmtf+IASzRHxbvslqJ1Fv/vXSFlU/dipRzNVQJk9zadb0
wzWmyEJTXgMq96LEaVLrbZFVqzcdc7EBaO5imPanncnt05XTWs2nghiKyXr6uNvB
D+TTI3BFT0X9Kb8ILXaIqzdlYEUpPdy5uOH/POvXs9bA3Lm7oY/5iEuvRhZaLe6x
K35WLP5XMyDTDAu3dmE6U21/w4MQ+Fj4c6ojksd6TEpYMrZ5IL1LaS8oafKyrtTj
MYJtQslfsvFlG17gKAE8/MKdkDjdsSvd2VTRMTKIl9g1BbL+PeGXE6dHxFkSEyUi
TXsQkkAHNjL1R6MUzGF+CDlt6ae6IlsMH8n4zDpmuM1DvBxKdl7HDhei5bAfyZqP
21/7yaTNrMG4sufjkvyW+VIIGRDv/ma8to9E5Z9ELkgb5bXyMTzSJggpoiCYwS9l
mpPZN//jwl1ny+o9tHQlzyGasTyFAJdetPlVoRJ5OS+QMsGY3cUyt0ZDeRzBnpJd
DkpbmvyjUcRQbrKqTgQ+mwxi2MNABfOZ6oVYO0rNnY6XtL1WRfvCviA9s/Aew9vU
qGRF6fCdTKhQm9NTKAK/FCNf6ycB8Qe0gBv+yzowSXqsKXMUYBCoQ6UZNAMrzcQf
5bMVZuel0sc9jIwN57zUkTWqLD5oIM1foHDG/nt6xl6mbfkiOXTMxAb5fbFas93T
OzV0IboSayFC6poy2O5Og0F6kFXsJHbAC0cBJPBqhQwBwTOxA60VfHL0WrknN5tp
HCh8UfIhPD7vt+zbmIOEuAKVdHvObyrldYG/ENiO7MHyKeVjwpEi+77Hx5shb+Yi
AtYNPPGn5tWIEw9jR/2PSkOwiqQLgkSCCySNiWHCt5D78UdWRfbKJy+cfarv759Y
wr+zjzdIc5ix/MnC54RVdlCY6cfPR4qWXWns2rbygguNN4TnhC0ccPAISRGuImuU
oaos9UsIrHbq48ErfIgElCO/R9H6RpBfW4c+vgPQoAQEE6w1/jDEZerfhD4MXuk7
A5yv6WxA/IVpxb2Hq9VpEuQlppwtlCYm7ZnoU1IlMtXxK4J5PZbfAk3EDt4Gsoir
Im/WBCo6v7vje72BK/NxZ9+jnudEV0PDrvFWJbUGPXB0Gd+AN48DuIGOLuvCdbEp
2/o4tuiSATP93mHoZ8CRlsIjh85aODpUhOVcb8uhxnrt72xKvApuQV0lQPE/aOBX
PLLhoucZk6cbqS4EYD98uubMo5bqBGUcksHuofrTH4e8srnaX7OSghsR1s4qom/T
SbcJ9H+x/W9gw7J+26AFKMJdpObmDQybkyaWiL1O53DDz3bHyg+GSFhpIvk7K5eb
mQRrXjG8uB7mqERU+a/fjCk5rwLkJiRzI9zm4VKZqtdITpYhEl5Ol9C3o1z927wh
aStBu3cRutyz58ecJnpOgu2yh4qubTeCopH7vuh7QrWzEOTFwopzkSHzRQaldhwd
HS+EV+k8EI1y0wuGVeeW5NnB4R3hRgu9ipKfEwgZRfYc1X7JjNQFVuvl5opuaUDd
w/fYDK3dM414W8DrxDcdZ9bi1hQHX070F4Y5SzvdfPPFIlZyeTPvyzZQyQIrJDAe
orK6a39MRUnMAUzykDKHdzMQL3SXfMPFCjtRs7G/DwaDt5CufOLUCECJ1N14MKxr
befmXjXKsyt8p2oth3FtAlLg5wiCf95SmQ/esrBTfxXHfBme4ft9oA2BQJRhIyu9
dSW+eWwfJ9mv4vHzb9Wfu6dubklFVZsIGh1z9u4PZurXAvWAqqn2iGS4k7lyDyog
RM7aAM7qOpt3aFoqo/Cm82cRbIj1G21hKiMwDzvzoe0m6xdb+kmTryEgrpNijDrO
PFlQou2G3CZUi5tjaK1etRC4s1Pyh3KK3vjwxoTi3qnG6piJFdJ5ddt5HD9y+nGq
CBOeU9KkZQxspjE11xVHGlWqFAu6DnGkWlOEFWJYFTuM8t1t9F70rAAklhApE9Ws
72sDH9pmZqOD9DD51SxqvyUMKONIR6ULRctGa0f2IpI8t7A1rJhNTfkVEi4/qUIC
I9a0IFv243BwpMXUGRYX8EuJPHidozDO5NNJUIdwcnizNHBg8A+beIqepLEM6dmK
0VKob7AdGEFZbHOdJFnwD9rEB+6/hrVRRJcTEoPa+Qzeco67kDoP8dJq/Mh37LxC
+Sq8mgGuTe1iyi9YnJYfwyvxMRpiiFAFNcdV0RIV7UqtBt9wCCi/aNv5VLryghQK
HfDwOAB0V5VeDAGWHXjCWQ==
`pragma protect end_protected
