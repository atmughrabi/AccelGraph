// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:45 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Dg9mSRfljBKi8qV/3gzKnRgdhG0KHBflRcO4ZyBgXofdDjxdrQ820o+ILUJ/zfTF
kqDQdk3Qu5oqdBQwBaI2mPdx/i94SfoeeKZVSjQETgbyruF/r4ZYKAnEshGJ0D7+
QCa9B1H3ABqvTKUbkFy5KMuNM7xAEFg70QrKbGy8HtE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 110208)
e1eZi+Op46yjyj9fuWcoO8L39jT/KOjrzcVBZ9l3FH4W8fG6K7p8He0SboxtVAIa
LYjOoR2jfeuQMYug2FKuyqyoGsngx7PCgC/w8fDIbXrXX21NiDLO1sAAF32m8KYS
N/qjwgkmECcxZwxK40QJ8dbMwIzaFBpv0rNB0y9vE1ez1ozwehd+kJSfuGTfAAfz
FKtMV2UWr4HpB/wZJovcLLpRs/5FHEJYQfSi8I3zuy5PiRyX9LEkhzFdcWSKn3HL
Jazufq/pkaGZnib9rtL47MZGWMgooIZVEITDYZ/6Cd+ZcBQhnPQbNI9iJF4/uakT
PxdBL85mR0I8x8Uv1vOelmnvCgg45uM21DU2zp+VLcB97RlpaE4nfxhkiSib1m1u
5ANTYJLjvX4gwIqwjei3Fy0DV/WEYX5nl92PTrrIy+rJFqu+VBN3+I0y7Z6n2UI7
VkcABZh1OsMG1qEWLlQrc8myyOga/DJus7FMRY/0XkSwHIyomYQ/u2935j4sPiQX
mt9M1TKQebvPphbUB+g8/9xVWM3KVwJeg+TsSyO5zxbQKwCKD+vMAMyblwRfsBBw
CQbONOEvvEINHzIDtAyVESKEzhVlVIxlkymnWsZ3hoYJdpntCGeo2VgA6XWIZt55
DfbqjsmIhA9iuESElIcI8ep4cbjz2PjoHO56cYWhhGp3Foeb0+SvAOFAvN8e2Err
NrDzC4lio8czAFpHRYg4vUD0yb9kwOQG+HeqvThqiHCngMn3Wku6BS3uNOY/BuKs
ODHkZlO86dNffqEX3s3GYwuouVBPTRFHM626b1PUIz1cuaH7pFcpMryeIk2hQO37
c50BhL5+Xk/7TqVMGiYsDdNl9z1tneuavWJMBRmwWBOoFqfFSNU7ibScQV38gQ8Z
nl7NEMESb2iclkeFP4FIeBw2Hli0XjzJSZipuUgkZqn1EgYivD5Ci+6t3QEjznWs
f6FuJwcFds0csKR0MRUFEEWg0btv4AkgvP5qAUbOqXGPqPAjDTf7ZAmuyafHhcVC
xzmoGG/d3yFwxd8UOS35/k2LH8XLaTHj6726jx8CxCs3EyEPGMJw3PPz3GWNZhqO
tUg6/eDcZ+ALSzIHKQ9gSM4DBpE8OS5Zqi9o2g+6tBghURVgnZ/iEVE/xQ2cD6zu
wdm5CNl/l3G5Grte9n4UisHgq8kmcPn15EAuL40pfiY+/e9GH1MI6mgebm+wt2Z4
Ns8gT/uqExnA8xUl0u0XXRg/C8GwRLMyssbyln9q8R4YUXfAJa6S2H/3S6FdY/TH
kqeGia+ssNNXO6R7PzAzBEkngo64rxbojO2EwcgrGLFy8lV5ykEniimL4of4rQA2
pVvLe5CHQlI0V9D3xmdRd5QD3Fg5uX72aWMa+2WV/OqCn2EEbDkP1zVibzBwSoC8
yYFdEGRXPj0AcKdcUBg+ZnpzyXz00o3G5b7yfU624lX+5LPq/TI8pgY1d+8NSCia
uPYqrNV9UhqhjN+bDXeXcwStt8AfIebAKc3Sx5znFF6PuURpJg9dMU67B7DPdYUN
Py3OHDOGyORmR248Phmsp2ioaD46S2uakMxka08uq4ZSRP/1zkKXTeM48VNgUnU2
AzMTQKuH1PYdN2lofRQfVaVACt6QjR+dsXYqDAt5eGCbNEQ3ryqZR6dEWybjLe37
8xAh1Z/aQbBtQnlZ3kU7p15tmvJAxnghV2jP1Bjs35Jt3oZ4nu1N+WxivViARsLY
/fBgrFz8iJKzVhg4ror375JYqPloslNNIGmF40cV2N1MXBsHBvggHW/jGT8tb/EY
HzTHfs8maAmbYKeZoo7M5ot4II5xyUuaRLhBQZEzUOfOS9n2H0n3uglU5PjMztOf
exH1aVKpfdCFmARdJVg5ZAaPwH96HpaSDzCPMMBPma10k6AQRFXC8KSM0hXQP46Y
+DKrgaTN7AyEUsHzZ8570pCkpwBarEwmuAa93zXliJo6PcyF+MesdYVdfNJSANGJ
blwIIab/rzyDsixTte6lbcKvhQq2ulhXxrqMwqdPWh+qYfsageMGFpkrS07vOxRC
EKRtXNIR2auVbl7ubuBeUQKJU2ZaNKLpCYfrRUFjdeBK2cDzVtvb5QvYY+L8dOmY
MATTbVUmjQ2HvxUfIZsbHcm6TONqjB6HVAKd+//21owmkS5xL78BbX9YqddGiSgF
zGzFeKT6trATJn5GX9wBmMtPUCMy5HMMQdQ6O7bXJMUMGiVzMffLyfviPZu3vinY
SYGEWt4puMOVYMm2TS8yDFUnKO9AzYqQJd+crawtUadKjKNyu7Hi6xl9bOWXjlP8
YPyLDWhvQkI4IZuGCyYCVZAo2plavXPutelb01tzScKQRc69FUlWkk9bidyohhn9
tQPSa1s60g1oxmch9ZRsWJy5lQOLubGztHzrZ/s2Qmpdq513R9iI5QdjA5/Rkxog
mcgu9SkdrKMHFhxKfl42nqPs9/853I3wI+P7odJBz8ElArZ4EpCm6CCjd5gC4mS1
/GMmRs6nOtqVOcTqNnx/RstqFhmFLUE4BquRDIUFeeEiW2SAqL1Dpe/yn4DyNqhn
grW1WXIxECTqE856AVHfxrW4fVuE6Ali6aWkuMBKsrljM0xlPW2G729nxL7fz+b+
lRIi6jGEPf+NZoNLvHxnLPQG7CXDhkfXgUey36xsnURA7IHZslpOjrSQGQQMfW9m
C38bmPmZj8FRhxpbIWnImCJMqKAnrf45GCEvGyrbc0YucP56C1Ja6Njm+fbRSF5z
rNFuYTB9Zhor/PzTUnMRxGgbkeAmf7hA2PETc+kSC5i/qHFbICrAlYZytEgpCaFz
TY89Bvy93olRxZZlNrV0enKhUl2XNO+zGWWewlUz4LmWcL8+rM9HAiG6lBufGfGG
apq6jHZRNg814XhKyHnfVatOR64zZnzjenG80A/3GkyZ1oqTULa4wWlfEYlzT224
Ou+IF/Sbw5n+/dX6uDN4SpZJh7Rrj5Ipp05J1ydKvwhxf3EcGnC+5VjUAPudAJCt
K7rvCPlQ0UqNij6iXfdtBYJ8qiuN1dW6x+PDvohRAnUqT0vNZeDAcpgPYI76IWAz
ofU5eXNjKz57oMPv+yns6sKYeayoCb5I1Z7YxwkvE7AtMMZMToMhjL+RD6G9cAIG
GOr1Pvxw20E2qkXGFFaLrIcwHTTV2NPE0I+AY1c+tGqu4PfPQFNWHVnyb2dKXc6V
WO5PnYdRy62phTzYec0LNdklBoSBrxQLATznHx55ykK7mNXvj4cBtPyaVarnoVSG
HvlM+HNEpBnik64U2MnZNo744Ek9OGQLMy4QE1GdTxeLgVZqg/DlbTgqzy2YMYSq
zW6SJ5a3bL+1WAat53CA50UYsaPbMT37hmP15fouJRaLeMclEjvvRRpuk1VrjQL8
ahMVsjtoiBB9INg7Gm1XV6z1k9QCSuSKjxDvyq1mvTDAs/XTeyk38B3N65KTzA5J
NL22O6rcntEWK3bKWDd+5JQXY8vI2K1UP1WiRdtGM7vWBuOLSJgLdiTjx8HrIIIh
VTDyxzm+VhxzlMUfEeRY52cgbrBb+Ayl6D6XlgeIC6HbPO17FkV7TzKB+8E7PdSC
LqjBSBNPS1Q/SEyO9mkZM92X7Ro2pvivJcDMWeQRiaDcL9z2CLKtQ+ecRw+s3Mpv
HKj1TIb6/NhRKJmZKcafvsJ2iMFHZ9rFV53v5alh3IRAYIMeEn7QakWW5QAGwAWl
ZWESj/k3u++PA7SpF4kNvOXOJJ8oA4xi7JvJsBOjm9ZG+R9Rg9PQ65wm5RY4XeaA
8L5mHaVMdFT4733ya5enn1tKbIBjk0Ju4N03D0aNuz+noV3lJdG6zrJVaT1+DmaA
VLReYF4z/OPKi+jARfmyXvHMJM/T6+fltT7SWiTI08HgP20VTPL1sD7Y5wJyk/xQ
KYFOz2S3OTpUJyn+tOODqAHoAtByulU+M2trzdNGJxNHV9QzjytBDv/L0X2PkFfc
Wz7nnEX7q5O14PJNNa/4jWXRuBFJBUJ+z2GkoFm1QRrLCe85f3Cp0msxQCIJLd3/
cbSYmqMFk6LX+VRxn6dfTm3Yiag1R9yIVADBKWRniGyL2z5bjUroZa6HUmanLomi
DCfkIqRUriNlVkDTvxsa3N1kDbIqpz01KyhsKtAuFQEWoX0uKU4d24eBJRaqlNKv
WZbTSjdSRuc7gZJvWDEj1IEu2jpXmsky/u8zwazH7IWi/dNB5ZdAzDuyQUccKx2/
Kk6UsmS6TVVJtb5OFKWp/oyDtzPr/xOXq5Un+LG1ycwA9VllhgD+fDol2M74BbOl
LJNVmn2Bio5vPVEV0sZdRVEPqBW7y0W8VhqPxH9AvCIDwlC+eWNkkBANnUk8hq+B
FsQvZluJH76vYOVaRNwfasOrAnbIV3F/UxfH2n/A2W7PMQN7xHyvZ63vqRFH4Gg5
LLgepZqyYRJmzHSSSY1LTSv66tjX7utx54Z2rGrlQwCQGkToviyE3iNblmrPofJs
8JXJ73n7M1qNrPSDS+3Tnfe6QLcf/9LL6LxrMAmZl7HjJvBK1iOng7aDIqkS6Iix
tE87Bj7lUz9X60fHrt5V96noMgzKQLBSAB7tnBuCv1b1vKhaf9DYCJ/daCw3b0bC
NXbUNbpVK1Psr253b517ekfgXcUHmhqVF+VD0iMCi04cLbaj6KejkbfH2m5441Sa
6fdLgxRN6TXMWHDqz2b+cvVB869TTb4cwHg87hsBcuA1JbHT5H+93PJ0xXdXBM9X
SWlwT9K9tDnzCe2jyk3B7CCbuDEDV20W7k1LN6cCHnQ9hNkL6MNv5pvUu8pUVqID
T/3RfP2eN9yRpVIya34cwg3MysaVHdeeWdN++3hVNZlgPWm51Woxaen7PAHnAZmO
TQasg0nzc4W7Hh7CnEspwVFcCupYb/Z7WQmx11gmByUOlwTKNmhzAbfcqaEzvScN
zZGB8DRlzUrZsoGfZ8FnMnn10h0V1eYcxssJwIKUKmk9aMyU7hkAqHQYVZVnHcN/
kCDNlBd5Bvz6yymNn7FXnmpUwWCdgtOijfIt1FMhgKto7FOYs2j+I/NOE/sQHCKJ
RXaxfUqLB8xmEphM1zpmdjvT4QI4TyUOvQG3rXrP80Q+mOxQYaB6KpvRpBtuJ/R7
FKgULa9s3PjDgrpujfpiknKPKCRELxf7jLltIJFGWY3zVFgBsuLP/MQO9xrKrmaN
5h6qtjImci1AbdCiA3JaJvLEbYRAGt5cKbfnnuCFZxHSsMLRam7eU9A1TBYPXQje
sb0XiYkCr36ko0UYq9qf83LQQoe+jKSVo2VbpIHUGMY2m2kLBrIqhan5gDF+d98g
E6rNtCTCc6YTvjoMQElNrhWlwMQQxVXD/CuDOspTIvPGhX2yDxIjc9hlFK4hKWi3
E5vxIweoq9YrMH2zZRGPJBCmfiD1D+/L8vMat4QMWhBgYaDO+LWQ16GSpPQSCWfV
PmiAztBoYccJHy8c7lwkYvvZgQ3lak8GmZw9fzFwd8SdnC9EMNUgrPLX4RscFQt2
JtX8XB5lTVW2PquWRqthj8/u9FlUQvLPHFhR0Tx89r/dqEuLqrsQ2VWBOQy0exsW
7ehapfjsQV3PSSLIp1xG93ddMBkGR8rgb9MHSZDPsMovywvdHBTD0FJ69/CTLlxg
tjWMz+IFc9M5rqmguTXlSlU9HGdKBFedA9rel4j4QOIaAwgFdCqPakkiyuusXq78
q3pPs6THRySEov68tcyo+u6iTvnc0fzaqlb4HFv0ulOy3k11womY+E9K3krFnqfd
ynmnrtYvJ9PAkZQEiMArZw2IX/R2sXwkZUirE6hSIjEPJmz6uO4jSrX07tTRxVNN
632wYZhIHczKJPZJsXMy9PV/2Yosu7D4aOIsuwB4D2URvGxOPhHnAR6+Qm7qGyyS
XaoRjQAt46Xdm9nGj1CkyexskQoV+R64lDzR+Kmx+rbf247LalV1EedYvRLkNYAf
xJY3yavS2qLLMF85bK3SzpVC8cMD3z6GiKlyO5R5o/yuS0gHFwPMqLTrK0rxkDRU
Njj2dYHxS05V0ng3Z3fhwCTT83V4A/ixM+le1ySPWEqseX7lYGl9VJjWpf7xBv0x
Ntpt9n2is046vKdHl7qpMZ44U0MDaxQV881ML3H5FOke0TBwvDli6+CXWx9uBNoh
Lecng7HRVl1RtOUvWY11s/UYqlsyZk+yBm3YeBpfYZy686udwRdqyUXLu51FZdu9
dxav3FBsB7YYfZffJa2iDaC53F7UZo6y9tM366eLx9RjCtD8LoaPvTX94cbLvcMe
wUqoDiwpheIQgp/ldZ7eSMaFkUXXQcSLz3nVN9yzFoytC9PYcHQB0G/iI7kJUDfM
s2pBHA1VNefjkPka79AqqGphySTUsHJqmJvMPpAJUxHW1YeYzChVsw5YYdZ9GXXC
jcgXYAahWn8mWHeSApBx3jEhjWXGrlrFBf020lCVwbbuU+HBu7ivQh6vPK3Lrobo
8mqq+R8ZKzT75mo4TvqpjiNcw4bx/TrIcEjcCeu7S9zRyRaj+b4W3s1TSMAGXk5B
IvubQE5aWDk/u/wx0L6Wa8Mg2IY1GS+jG35BQOO0V+5cJKvub3km8Wjya8Cuw40S
If78f9Grv7aAA+FPKmH2JOicW7DPHhpsMjH0liG9/gduPw7Zyjmbhz6cRV+/38Jk
MHikMYMEkBztd5VeYQEAWuklwLVizvrkRrDz7+EDcbjPT125Wy3zeLfy/AffPYd8
pG3MNv9ZvcjSY+auQZ/IPWtVkxJBIgyuKqEQ4iKax9m4Rm/RLshPWtefIzJ3spwM
LEPzkDqw1fhgGdhfotH8bJXHNq5vhLHzstii40r7FdZ7bx/JYpj6qbGc4RYN7d3U
lnBaTn5pxQgnZTkIhZF3o0SmAeKmzyGUD6u1W+lu6YL2xryxeFZkV6GP8k7FanSJ
7HJU3qHABptW2tGD0J/L3ozNUQr79bMTTCfH8PPWTPEyLGvZgPAL8WDqTm2ZWZYW
RMqTqCwjUsk+RyVukkhVvL6wJAjwHBPHf03DGYyvpQ47GqHS+KjIHVcSvQAi9aJF
Hj6v5JC6frgoAnGzuNHAW3CLA3rwrbF5qSikeo2/wuurubEIKFN5VJaaOnPrnlUT
3ASSRPibg+Pg/Oz+PLoA4yQ+a3f5UnCU+TqO50L71FvPs16llpJfBVQJAGanleKT
fha5nbVegpWoiI2KKQyH2A+ltKu+J6K724+uO2CcaFgddxN5VatBhbvttVqU6Lgf
JzwdnG72JcEkRBoHc4nCqDO8tfOu8OEByiWGcPKRDwUdU6OTri5pnCUWpZWsCpYN
e/8jEaCoTt8fGIx2HPgNMcfR4ZpLrWfvOhe1BIoSsoV/LlxD+VQF22E+/teeCC/g
BEebZcKgULDsDZWmWCGwP9B7hOHwi9AU1OL07CDUHO5xMYMxQgWwGISki9316N8+
jYrMDRhcBS0ByaHPDP6ckEeBIHKzhlSlwyPdNEGKTBrEPk6/70L04vrYHB1QkBMR
tEVW5IERVocCWyL8OSEl1BZTR6qjs6e7MWIwHPq4sFXhL/TnYidNSNGzL9ksu50n
VEk0RU3hX8yqZfjwVk/gvud7S5AIqjH3rdPhBNfKXp83OnjFlzPfquf+/HBCpt1b
JqATXWyvGuMzSoE/ScmuEYYROZF75DeKBUi5rp7UF2fck9+LBa9Rv9sfU7zUjLGx
+wUs/0znJCYxSzI6ftXLSn/MBYlT6fijVIPPdCSY9/ucinnnECalu1zZyKTECPGy
kEwW7zrLDKqQfBDP+i6bzB44PW9I4Q6eORfhIQyoiwAEGiPMGRuVo3tUCCzzBURZ
+884T2RgfDJcz3mOmsczvf7sC+q6ns3F5x/DnSP7zmy7z/w6ZfF+E4RdcE+Bn1dR
VQBv0g37Q6FA9H+PU3KRFV+kivpJ2xtTBvzJpsI4pL8oU1uViZZipQaCd2PTcirZ
hsTRAI8J7cfsD35fHU3nvogJ7kz4gmE+y3h8abk2fubfZT2SyP77dF/nFVjDSKqn
L5KGDa0H9FNunXDYJ4vA7qCv1ab77KwEWRudDOdAWZzgSgiuk7CXFXvnuJy/hImR
B3jGJzmh78PlFoT6TeQkzLFWRIDiO3Jz4dokC07AUNVMwFWGnyQH/R9OxGPxWL9e
OT7cQR+UGl5z53pqzhBTyiyIneHlLW9y+QnIvoHEksq2r9+8RQBl1Dyl4wlPmkyb
OUP1JL3Cr+M8QqzLBlyBr+x/UWfENFYYBaSjAlRja6+ZY8CTB+9qJ4QoIH8yulLE
/ribFRX+Kx2Ygy1wG8ak9fMiyzZnNrrV/sJ2OITZ7kclcGELRew9MJ7Dve9zWEcn
W9Ru3KFMVIHTtaPOZyMCVPppZzomRfYWOmP/2jyVVeOg2xak3rxEsNMNfna7wquN
A/JhJFEuf0mQJJDJhnkT8A48P6oFaanXy2Y4gJwCqHfCWZALTlmDU2JAEl23Tamu
oOmlfd2uTDZa6Qf233Dv7JsK0W6V6v+4LRGcDueVGLSbMWPTtz0GTPohMhUjl0Ab
syze6VujTuHvvWgIBw2d6hhV/k+cW3nPtehdgteaUOvvpjTA9HX/mASGdKKSv9fg
apjQxsD3lcaHDTLawjqvFSNyX/OIU8RsUtg8RSOWXDaPMvd0v6liDQMmNECbfrfl
vVRzNdVBOwNYfFvbqT5uV71xe15P2EDPzsqEx6S9qHA+hLW3onwlGCBJ1gxIQR4k
w/x9QLC/VqS3JSyfBkZKGDV24aUnKxBj4N/ADNw2/mKuCfm10qBehKb0m9kSP8g0
7+5mgifvQwg5vJHjFsPV3mtl6Qi+d9CEh6oSLyLTkVHW9RC1bJgffhqVGMmUvmy0
Cn5PaOwEPO1hZy5zS6oBGxoss9/M86Ul3faEzxnQODtsR4jz1J/j5vXzUiJGg3Ba
hJijF5BSeKgr2gXfFE7x4IiznnaIfhed1e32peMG9H283BMK0PHjt8tpsuJBDkuJ
2nt1WIZzfj47t85K2nmA1Td2oEomAUPhPPVlFUdOig/rYsrDUjIT2Jo7KHEdtHgZ
EEdTfkKNdzx3euXYCCWk7awgdYAxCDYzmDVjsLWBFgVBjTSdeK5N6bkVUtbUKrsg
+IScX5diGnR/KE4tg98Schf4gI/btzqK7Kr6s5ZSpRRqg0hLydb1Ejkn+OpQUR3d
kgvtgVSUcvplk1aZ/d3P7xb/2hn22V5pju8R62ElCcQS3g1n1sqrbfAKSGdpClCm
6yAT08uLiYnb5+QvYmc/x6oV1ZzwZ6kmYYighdi66ry0nxWeT9h6C5e18+q1kVLi
6+bzyb7F/oas4qpRd3TgktH4o3XjUs01OoaoF2CTnEKIoFdhr59RbN2bh8Cov30V
g4irKjWM/a3CN2ZHlXZDYT9m54eN1yMSriraP4eJMdvfCfdLCKTYXLQJYfn87Wny
0L2Red0S6tTCRN1/2nAvnso8T+CmG7pyo+iJKQXqGFqDjUFxuW46sXb6jKbtm9ci
cdmhCANzeaLoDgAkAkgMhGOsF05lp0tqrZMlYsakZmX0ZACxmmvJK048nEFWLJcO
hpBmFObMjYqJCDW7nfJ3UpLCid3p6l3gsI+SWKlX3Ol4hMKKaTAuNKjL4uFdyMPA
m8H20eeROynqwrQ3SprRnctKhRILEn5VXupXdK4dNJL7VYx25J4hPu8o7lj756BG
I8bpY5922w/cx4syMdQvmfYLi07DzD2Gl8ItrOyeTzoTFWUyIO13J+3MbphB3CVC
QZMHT1OnlLzR3ET8EweEmp3bgiR5t11i+KtJVqn/S1vPZ/0SbGB4exqLDHpgb/5j
qORGkj3K7TrJ8NZmMRPL8365xJ1pBHrwNnOaFwJFa54VnZ0pUG02Go5ezN94KEbR
I6Fcbloy44NgL9aJMeAktEgT/dBbvfLkZCOqSTlKiydklomjlIllSJm4BRKz10CM
p0SLJ3gQFX9jyP2wUwY0LhRBux7l8KUCj+GqyjV0aJFyjWTw9xDuJUm2GUsxuSq3
dSXAGvyxloxTOLlcXVXuZ9HDEyDHO4XyG//R+xbr+FMXUdsG7QDezoLgjf5nWv0W
1bMYeLOvGXdA6+JnZEkb2J4SPU6CCZkr5ZisuzuxKZ4X4KBa0A2aoDhgXLvAkSJM
IX0p46GhlMUhV98D644t8ToxN23f7/QFlywUR1I3EhCKeJhRONMEOxm1/IncXtv8
MDTHMZAhI4hIz4OeEtu780gYSEA5pE6sgon+MYviASE0jkBm+1KqTHa0nqsn6YQE
SxWaZvwsxtKhyQ8/g7OkRXARaKxV0YVX6VudK2/sonr6l6uBFhuIKuapxuPV/l2z
bT//j4iw45/xlbJyxKvQN74380ketl08ftxCk4Dj2p/tA9DT5bjnHqtGTslYuKk0
QCMv1ie+2WvRom1H9BhVXZufyFRKe/PK16jzFHE5K3w+DBxjJYqTFpS/7XFZSCnu
qVXOKsRF10KXanvrJnQ4MypNYCZtrNYiye94PGJv+wr7uCtHKSm0MtY8omaGiUuQ
wA8PH07zEoL66/QhwidDvRgQKtN2+zCpk6/TXCj1Wk3NGU5dXa4FFDcx0AbF4ogh
eLudMWAiWvbC+yKxVVTM8sKu5EDlfe3cJIPfB6vwDU9aQoVCr7Ode8nLvwoU6ra9
KWj9ajYQ+h2iKDcvIIgv3TrhgwXoXtpMWKkIJp9GYAou/sI25t9gL5E83QiJMGaO
huQcXbXwaBiZ3Rnnto+WvCQ6AxRcGnjMhZ3Mr5eSoac6jQdhApAHw81ur2O51hTA
jwzEdad7gF4cyqMCWfpyNEP9UkzWCZW9QPhprmTjYDGD48abqhLPmpi2nBvSFK0W
MYa9LljCMDjfWAlrjT4JYXwuIVI9kGAK96DnzYTU3wNqtcnNo0r//7/V7/VlD5O6
OYoF8o0+weSh5pmLINg4qZWla6zmFWupylzH9fBwzdNClPDwMHlzG/YqSBMx6Mck
Y8cxoNNI6QkNIjN6q4aJRoKM5ANrECSKMuZ4QwMAETWYi8a8yk2mKbbdunTKp2un
V4YtG0ljaEb80YQwtL98JOHH74WBPZzrgyWR7+iAcEMIFvpyAj/4LA1SHbTzCv9o
AxiUo0TAWBngBFa1Z0AxwQszvSgag70AEhJcjP8mYM5KhbcWxHTb1j2qnyF1tZOI
iAqf3E3osOGMM0TxKfBh1rJbU2b/SllzOE5rCNCF43tWTkrRP8t5g3GxYB8SYdBR
RAykXUidtM03ivEiFFBXcENGa5nMDkZlhHsNr85gaxoaO2tZWmBLeoeU3v2jTfIQ
Fws1C8WfK88+sbtwAxK6Io/XkPB/mYtMXZbC4leE959iWIkCLatXx8bx+7603YdZ
EzArGJ5aUyLaCIMKeelnRk20kyeu+exc1f/JgVB3kmVXSKKNJC9W5tR230Mb5iRQ
0UdglHubmHsyKUIMZ6BcXpo9I0C19V7mP0sWVyGjfyEZO0cn7Ez7Oucd55FoowHt
ydZhKCbgvn2w5R6iwRem4Go/BuLarFSZiKcjSJSEfZ4MQeGTMz98yTa9SrMuotrx
8D5rd0XeGPv6/SFt4vpg2FA+gcPdJZwFrQqie/PWukd+ZgkM2r4GVU76HMw08Q9T
e9P20tAujaLoOO0wajuXpl4Agz20KltinlYKMGkIY1z7ttuNQ7H0wBdastLKreNP
tYVQLLhJ4C4f/UjCHUEOwcPTfC9c0zN13Nd6QlljN524INBFPCqIzqXjgc6FzNai
pqyHTtL0/LjfLQA8wpX0J9LA+TVQ02B2cHe+JXju5XGtZr8fq4QVMSH38CsrkuRS
UIvF5hI8wwBpTAdPms+J5W3YdjwRdKgR8gZEzyLChLZnMHJWTsRaTPqG0eghEXMg
YhTqyIMMvJcgnPEvLDoacE1N/sV+5lI3UoMGXfkk4yovNxStySHss876SyGNzMQE
dQkJPKdhpgORVdseL9QoO0/i3Y3Q4pPceGbo+WNaQfDPaG8sLV5uY7H+szpDI67w
L/IUBmDZz22oIsMj65bCk7ELzqA1nc9irJpAesTayxjHbgEdTxuHksS6ysis5+Dn
/JXXbbHCMA/8eja0n5YDcqJQ9Ol/P3L1JWOCB/1jb/aIj2bVpptxFCDkuDaCofyD
vQOITnMZeAsb1wOtIztjqx5smkzAYojg6fK/MTAzfmcn0NyRngX4RhhBX8UW7oGK
aQp9+FhC8Pjs4oa/FAEVDu/v72GeJ9RE325SzAQYN/Zq9ubXgOi9AGTPX4kx+XHZ
iO/Cx+NH4cEBbceROdQzwV0i4UXG1jWOzjyUmipCFS4156LCzdPltkUrAVvV7gZX
jTXtgAsVXJsea89/l7vUxEfWg9HxWN9YVrVdI0tLVcyb+GnHPNImcpi5/QL0iLpn
oc1H17aJJ9SN+WLQqtKPbJd3nNURdt5V5dfcgL8lKw9z5hi/Up+3ZdUw+GzUpdjH
xMmaDOJy/QG/ySZ55x6N8wygVU2ZUcIHl9dkjtLOq3FUNECYeFgydxI41Ng4rSUp
eTPOL5dq22dRtuGSBSq0C5Drw7NSRJQto1uWU/25aFPQZEGlWG2YB03VXiqajlS+
nLgCtJWKS733C/h9+JuSWRQdRDnDYiGGWvpuzH/xyvN0iH0ZhvkiW/clw5UGoGUQ
WdGZO9cwT4kbjUtcogPF3i0543syR89K43U4IYomBBZ4Vo5vKDhavlob/c2szV1k
M5n9LZJrVDZlsXaacup/CxxdR1NWJUh0blo41DI+tNXonMMRHV4hpBVOp+oEyEr8
3DjdRS1pegC5YB+eP9i3qlyNHU1w5J9RSqcInLLaL2XZojZHRlptj1ukMTRFTGb0
4EYcFKPVNceNwYDgiumcSIjQz5bAd3RKp3/Kpby4GySmR2fJepJ+PNbG8DGKQSAn
7SjaR85AX3xL1pSvXIqBzEvs6Qlu1ezwJWjhOuVzD7TN3RzKepVU/m9fYUCZ4lgp
teFylx8ymeeqtrexPxKP2CamOMNcQ+Xq4KPA6ie66bjXS4hnKFycfVe8Xka94Ht2
2Nok/M7VH54tWgF0owRAMj9B150RolaZ3kgVxJt/nJ5M+ij+Q+8BxgIJf9vR3BKv
8xxe5S1stWCAJKvdcQtXQ+Ta9M8K1NifQRJrPqBrrITy6I6sxnzIx3qOHRf7ze7O
gkil1SRoj0xtlQ6mHlq8C54I0ojhYSAqip0Zdz5NSmyu9LLsAJCMi7bULJW/FbqV
S3lTv1XJsiYm+CN9oFPHNjPZKiR8LKXrbo4UOvBCHXu2Zvw/6fVymv3vgtq1jgtA
djZlZ0RyeU/vx7Yl01VFYY98uaF9k41cbU5t5a1v7JyMG5/3pvyklqnnxc38gbF4
UC090GnHiT9MrsyuPiKTyxv6bkEuSqz2rNK3h9USmbL0b+aVvKqhgP+ATdfXm+VL
Xqm0fkrTtUrD+6juETBhoykIc0MgYqLtlQBRUR+CJ1gLhhKuIBhtxmDxWpWxpmQ1
6+CpdE9uIegULhV+hPqCOSJaGenQws6nPDIcXj+xpwrCAUtDJ73eIcwrMN35tNI0
kyiTF+1qkKtY4eJeFBSRJiG7ly00B2VQWIqPapaVTNUHAqJC2PQOiDFpgQJJkr+F
jQkDzqkkwJYgYMl/E14N2GEZEQdw2fje+b3ZOVZikiruSs6nw2mvdCJjmVv7A4hj
qmrzZhMHXUj9UuQ8ojO6UGABk7Vjf7hkCFvtb4UkHu7AVKi7YAwQFIdi44cigkST
puD5ymwjOQRw8zC+/AXi+H7FAeCgrHYqB8BcD1xPaQktPwTEtdZdDAZoU3iDgWjB
xPHctrW7/B495VAWvb40bC+FPmTZAfK/kixE5jM8b1tAJeCqsVXT34j2coeCf9IP
bIknmgaKKGpXdKHDjf7kUCgH4bFDWnr/OtRq0qnoaB7qxabkDoKyZ54nXsCKgErD
FhBf3XeqMHlXyScPwSCr0kfaStipESnHhRTVuMw13QaWStauRGgvpg4+ZOeoaWqT
v/Qt/6aod7nDizNOL31Quyo1idwMKdODxiex4hzy7GJdNc5HgH5f/KXOLBgI8nFB
m7b2CP+GfhfMqdV4uLyG8MnblYFxw8xOZ6Zegw8xt5ND+ggHILMRWNp+sHVjnGts
oXpM802m/9pkI4CJaxanM9eiSNYYrT5sYs7qSXGBShP2kbkobiFK+MTiJlTAr61Q
VI4O/L7g3p77Ka7NX9CGzvoGbiq3LoiawOeD5/EsvgdaBUT+Xewi3kZmP78KszKE
5jg36thqWQUoW42Kco7gb8FvkDg2zRFqLR32CbUnRwAueha1kDklXI+PwazaT4qP
N9Bj1SyFEi7HtYig6x3UKS5a3uBLPEa1IH4dXykjTkD91NxJSTU5u9uMXgXgATyf
Ec3tNCz7L+xve6v2B6qr17/SKvTgT/iWVqQLCIlJxGndW7rD8WF/SvuTQruNFqyw
mLICYdgTNnZlAUrgwaELv0nSorj+LyDZ9YAp81M+Ly3U9x52kyHD2Uy1jxxPXR6C
IxxMUy97Gl4HNw8y2unTLQIM/b1iOxcUr7wB3st5pc4izsXFinbMAzfI4h6/aMdI
vFsR+0pzNTNktFs0N8AY/dQTfUB5MAbehhGw7D3HLik0blWx9nhP/ufWx6WWHoe6
6Sewp7VUoGmp3u5Yd2m7oK/tJxjmrqLs1VjBBfIpW0+6VeL6cY7oAifEi8FefXUY
OiP3uRzSpQORfkO7mPa0okM0sGUMuIVpy9txQSTkk+UUu+efAmnCnO9BUZ/0EQtT
mtBMkD3GWQHMfs9tYc9Afiqf6OjhewO66iix4sCdh0xseMPOsfkeArJnieF+GU6S
15n1lsXuB+1ywmDTn6Erd0fPICUnb4kphv4F4fTzUMS0Rh1P2QunW4fUvjgUS/le
EV33ZoPAIhtCvOdcNdYdJdMYbGgPE4ZlznBqFhCHbRPsWeIf9lKu7mg+QaBe59D0
uBy/ZSUQGBybFLNfcjdR2SEGhZfCxI83JjDAuxhqWyRWn1y5m8qsOLFFXpdqMpNw
WsDtD/TlZQ1xlTLiyLdW/yMbqzdICEF08ssvffD1lZuJzhMnPIaeMigJegnmuPJO
meGWZ41vXcai9tYKXpFxTqlVUUyzRCqOu9cbKCzVZOP3ueIj8vBLhQaGp5jbZzJD
GtAnoZYZe1ZVl1HJ1BJHOBysNO0X1zFt7UmVzRdcBvBxR0c1MI63EOQZWU0IwGtk
O3FJTHAd9GMt2OVHbwRN4Rw954rJXYdEZgEg1Uf5ug0VRuZLpkXzjZkXE61rs04f
TyWVGHrqIcxhOjNIc+y940Ho+89abwVznWOTUwsXUwIvh8/8HTpG1Eg7SvDizg1w
dJ37asAhR2enMGCjSzmrjyEbEDeE069v3tgwqgZhNntgPQ2WS1XY7vlc1NfZshZt
i4do65CNGbkzqV2K4t9wbOunhpWxNd7TFaThjqCjNaQg4Qlq2gIsOKhTZst2vyaA
K4dyYX7JfYCP16RI1iu4Lu904glEx91ZI3BYkjntMClOeZqt8OYudQS8ywL4PQA+
qF4k208xqEbun920c7f6IPB4ybGDCoqySgjP+rVvnbjeDynxT0lHwO/jzNG96lMG
oMAKXccfM8eIrZG26gvEOo+Z5vPrvMFk+CUSWTPX2EJQ3P6esUwIe1K+wC1Z+pWo
RoClYYOraSA2C4azF7VE4BzvtSTIsTmAST8nHsvpv/CWYbwFF7x1OlxdNgDYLcFw
ZdtpwN8ug6TlO2x3eI94u/fOYYoQZd15cm/CvOMB7OO43zn0sJOxdGAiOD6hw2RB
n/RorJECuM7Xsom1zM1l3U5DYWGUvOB+oX8NM/8UkHjQO5zYl+VRWp1E+Nu+OU6c
ke809eRbQkOk0drDLDILpbig+5Q/sWFugcZpoDRbLnCW8rmzsf6lh5pVEfYK62Pl
cyOuDKjlHAzXFt/26p9hrSTLhTDdfyOhLjkMIOIh1TkeZWtNEt4wH9MFRUjGWcuk
kqrMuU55a9V0jgsqORXu5xR+6BrBg5VuSI9Gg5tOqyl1XppYH7YkDGNS+lGsewbH
q2keSNGU/0FWBvkfyHTKzcRYesLOiqEUaEWJZ17AwVrZW/5wF0+2oIFC6TLkXeGl
Zwh/HzvaEVTONq2NAWyvKryrH9D9FZKOTlYYH+gYCijj4c94MQi/zCqj/2t7yAnB
qJlrfT99Vh6rKeyIjWvtmL77Mk/vAEsiLh6Mk1NZjyVNVVGo++1s7+sa25vmEx86
GGYdz6i2aLkVGRR0dMXRXhcffBzkMwrRY9IIb8kGYVZdeT+AJrXHh7SXmsSg/aOM
3Q8aJYr7Rf7YM2Z+x66OoK8qaO1x1/qF6Ii5/Le7S3vUfBk0fbjSvYWP0QVog0YD
KqQIUVG9BrQ3YVZKmOge3GIYpXHXbhO0WWdwsHYIcYdAH4zjKxafQA4kcLUGRQrG
M2hjcYn2Edpp1Wo84dsaXkEmYHvyNnYDxAkm1rPXp1ba1CLPwc7Vj+pTYsUQmrVG
jdl3E3ZFUbHzmy8zA0xOFY4yjryL0cDXW8Zt7mwHtK7gSbB+eEW3vyQeholwLDDS
1nC9YmDFZtOCYNiIecXz+159u0J+OQgjLobo4VXiUJMiigZmQ7GcbcjKw7QjC4Uw
5mU1poR0nshzuOVrS8+1X0rBq9HcO5NVaXMltiAP+DfG9zop7hTBtCDPb7wwwkBj
6kGvFASHXgoMv+d50Tm0fV28ajv7Lgq4aUhH6cZ3/da+7a8g4+wHU4LhDCeEoG94
0H0vyVdDYi6lN5b5kYxYXNGfYnxrINw2tzckwXrX8oaeIpPtIxXtwodyFtDZ5coL
LDsbt3aQ2BebBpuaCtjGZ0xC6V2gb54YaE7WqmOXQ9aXg6fP+5JWG///vT3IrG6n
hr0kjZ4DGoaVOAGOZ0YjoLJGMDDDO54mz31tPv7KtR9eCW42VhIeD2qlxaQnxxTO
lFE4yt7/c2d+SqZFTyypeheMR/rGncVT81YnAhOln3E/B3hbBhq9Ioa9UN0munIc
yG5SghYDheNLskhCiV5afxqENCtEF+Y4HmWXgAUQvzPPNtXviqvkKNFioSirJ3+4
FdiaVmyLNzcOCJtG9ImiY/B0qj4Z88GKi1xzl6R9Gh8Dji18qdrPqz5leIqqJLAf
QNd9rq2/GVUiBIze3Q0+d/rzQTQhI/DHrMcDRa+GlaSZVHw4ZijKCjCt+/6CgEJ1
FNNdhwKTkCPzcp/n10ZOMtq5THAeur8jSKfQf8UmzuMC7dWYP0HoR3/AkY4ZDELz
bn6EHQYGd0i82/DofD0cj3t+WbVhHLKvlBn/jh9y558z+w3YVHwx2woYj2FjGTDL
vRozk4EG6y8SH0KScWHcRrUsdmqlTJ2KDj05SPMrkItghlSHUTmE2ekFmeWfp7EW
T32NaAGSxsGAT9FqzpU9/Vf43kpiCgpJjP/KVk4p6tEs7H3LVE7xRDSKnEmyp9Ig
ypxft2cO+5Vtltu+1NMyzEmhHfJo4BXXHj7jw/rIUH20/dNXFSMW1mDmyWh4LLwf
3RIAhbFdLRwTjjfzsXugMD6Mq9jhw6yWSJ/SucrqU9isBrug2ABvK1a8rst5Z0Uh
TMucLMvi6rTBQb9qQIGfCAxL29sMhgNifH3FSXdZV75ze1iwZktXe2buTOCHSSzK
WQQuD3QdD8CZOb1leeRxv9Ne+Iw5Lbde27bP2Bp7hhgDqO78m51/ZKHHBd+s8Uce
+vnqiMduH+wUrsvoeZEEw1/HWr+QEBj6XvCTtVkyxIlFtBO6mvPq73ZQoTRKnpvd
F+WYs7O9L+mRjYwxmBPJMmvgb6HIUUh3vXtZMEPV8UdqIf5pGBTVZ4wJ+HExBpCO
q22iHwJgg9QxkNrReBVDUWHQFs0Y0mYclj+PrbMUtbLALDSM1lxY0XULtT6hUUql
3R3SwiPLwBzXEQMXNNwCvY7y5aXB5BK4iDGR7jWfxpYla/VrSYaTWXH2G8vzQ3Qm
cykytifNmo6YN0ccn/tPdUKHM9zCt8ga8KeHw3mVMIDcCIw6QrQU1eoYnRnIXEcl
UBQHHfSftMhou29WgGuwSki6OIPRatbSZGZurolIKLA2z/JAs5vhaEStA4HhJ7LX
McAAhIyBQ8kmy33FlEn7lN0FR+KyxhPT01g+7G7UZqs6Ji2wvn1/nvVhethxwuta
TE8gTJjMhqPjI8+AsDb9U7i7mDRmAn+IIRx51qvwQpNkYLUfaGLNLHSXVDrPNmwS
1o67v9kkEaQAqR1Fa+aI2E2cU9a60CI8kEMR7rl9EwS2b30gIr3uioqxQtnyKaJt
fbwFhrRXptZ900G2kqyuDSGdyFraua2lzyFHcmfwmCxvCLpUwHMXrJRtFrNiAQzf
yQwokrH3x5VjQkOLTxRqdZj9YfTdPjkioHjZIP++CbFK7mvGuk4RO3DpxeW/vbxX
mhLYhgX+QguxhcatscsLujrnyyE7hsRolQvhG+Aw/ONtIMo/+IWzr5cbMuwQVeOo
U0a/G8PGSmW4/Jw8EcRQHAtnJ61McZHQTkpFUGjG9Dd4z3h3HA7f8adR4iaFc6sB
MyvQvNxV7zkGgqDc5TEZIj+mkUyfdiLD/Rhaxj8s5asJCd4rrKEiKFHKGYaxRNdQ
/3DqqTLankh1m8Xlv5pTh0zQmb7GcIeGBOrsBoRUWY7LHrn08bFj4Uoh6Phlniet
7xF3YrieXSsoW5KvpjV/Nz3zCidbFLZu+WqGca0joMsJgZ7HnozezjmSLDWKtwog
+fO0x9Nri52oaxzUIZzt9cuI5Y6kzysB/QhYnU7Epd0W0fZowhq9+nzmv7kvADXO
8CHBGdIuwS+ddzCv83HwrdOnINnEjZLx4n4YVOdlmYzFJo1gmVYOB6rYU0IdmXXD
vEl0qTsG1yK4ZpSz+OMRPEjjHDy9zq1qLvReyn+ivfwCID62HfCo+9LCLqYCe/9m
eYTc3Ut4tUz5QUVt/zZzCC9stD8Ya9eZE+qkaq6+fpqGrnjxghChmOF79yXJm/b4
YR3JHDW2qQupPMbjjP52UYrDB12kja9jHi/w+T8HYV80fiorWEH9i/tlj10DqYDF
MQ0rmTaxVixBoumRma4fn0QN7ok3KgQfg5bwumOSIsJ/Cs9mT8GvhQ8QSvGAdM0P
fUHP59TILmwmY4VaZnwHgWKYfSSPu4aZa7lwKn/2UU86Sic424gFbOIZPJizTV96
QlTvOrJmL9EC9XZGboEI+HpcPUi+bC1JbOaUFaAomfmFBNnPXS+h0nd8VA7EqNJT
ouG/fvj8k9SV0sDbJmzFRzrfkUvhIYoHFtsr5BALZuOuzbPZZHwobiI0Pl9ZVNex
Bd+0ytG2G954AEuJHhe0Rb5z4WDuFQ0Xd78x2FR/AfiAwfmL8x7pLZvZDIHGYsgr
0TtC8Mj6sfQRt5d0aywlxf8YvWX2pMO4FuW6m2kQ5aKsNhJ2ygfalLP/Oi0VL1/E
X13Ze5q8VM0oFCw8bemz6P7642a7DtzS2XF9+BpvJnANaeoQghXbbOnUcXTY3Y4v
togi7gEsLPtS6OApFJ9nLPTZfxk+7Tx/x8WBvECueg5sxoSMb5nQ3F32Pn2xm8hV
m5BSnAzFUjNaHLO63vf6BreLRlm8VAnKd8eclKBc5Ytgyttu1AiXR417owZZnae6
r3KlXgL1LSn/uN1Am9se2SPftY9RRiFVgPx+t9JeAzsmMhQfyuFeruq73U+Mt0K+
6SQI+y6g8OqZOahkeixiN3KqemVhkvnkyduBgaAYPD54bHL3HT/T8dAEmcvKe5KC
BXhw7ZgI7NBKNFVhnijj5zapE/9SOhqDccs7JBAUGdVOP66sA0tgF6WuyugVhFLg
/5QL7KYQg+vF7yoJTMEl0Q15ept4jNjwIsNKGkG2lXqTOS9QiIz/eekW0qqHkDd7
dih7y71yt4N6OtpvnkDpoLTnTA4iDt1dH7YqLw0hu2DktNuNsjtiW87/fJhDNPBr
2GuBVGJ0wreouOxdiUhv/NZ73PTiqIRubovUuEWAWmvOme7KZUMaRbxtxWKqN8hl
jJ0VAx4U7l0aB0sZfn60O8PWPkU+MMGRyCfrsO5ZuKO69Apu3BmkDWC+rl94Gi1o
dt+DSiEG+0ChMuyE7cHeMFY5wlCCgswShSqJOu9kuHxscG9upXm++xdvJ552VLsA
AOIc0nWlP+tAXDhk/t4x+LW8GeURWgAsTCsDpVwQKMxNWy2kcgGqO6l6nq80F6PZ
WFdRPlP+7xhzhOyhUkaxf3fZBpI2acvsSWjZ1mjJsb7Nzm1AkNrT4vnzEH4NFEUf
7sWmG8PtyCKC2+Zjv5LVUHfXklO/5wYiUOI+SIBoLy+iNo0r871xApQTrHhloRoM
k/eNCvcqwfxczSB1YTlbbebXuq8GJMZPKQ2M+Ukg1wCisg0J3uk09ESqGtsMc3vY
61tK1QZAl+8xcPg9TLsGyzZso6aAeNLXs2PreqrSAhZQfJLnJI8cCvqt2eQYuYNW
CJ/rHvVtaU+HnH+sFzpgxWB0d7sC+MJG1RaIMEJcQv8LmTSgKIIHSK5fCphoT1HC
oc3fS7zX+R3/hwY6O7EDUPsNR7QEYSyX1LoaN0PMZ/X2H+nS2/+tI+MJgh8MES1w
R996VVTyvOh9LObAzdvLZGYgUAf++u5c+VmEQwwSmB8deru0vJaLorIMHZ0J9sTH
mUZij8LPdQ8L3WY/IV/s8uV1w12ePzbC7Yz0+zdwmypwoQhVGnAwxv0JYouWcPz3
UadrIIxM5SDpWwcUHwkYHiXi4/JDqEca2KSuztgzaxk0U9dXEZPf03b5bhAVehti
jCydIsLC13q++KKuWf9ddic/QfQcEy7Gmx/Lqm/8KHXzzWUwEcmF/EO+BQWlcDBu
Nvvo4OMtu5QOPhxcUrJlRBgLIQH1rPNb99i3J/GoUdhKYtvHyUMXPINriaVFXV6b
5R+WXEQVjdgFEq6VPJ90Qb+I4m8gSGgOWHj6BEbZbSJBh15fv0QbR0Ok5vBdoN99
7FFByOLlAzxafnZ1JPAjVpMUWBw8KkhKNSuwSdOkFtbYEYbo3n4cSyhajZyjQcQu
+f440uLdFId2hAsFZgJag1+jB9joC3r4eSZW5GGA3IqRe2f+iGONA9Dk2/V9a2Sy
gz3NF5upaKz4WI2NKDoAmvaL8W/bn8EJpXT5UQWPtJnQDpjoxEqh5lPxTK+HkavQ
lIwHiLFBlfDJbEnvQIRl8Nh+5P2RImKWBP9DK2OEXYKIVZ9uC8zqX5RyVeHZk/cT
VNkpS2/wBcFYs08sZ3e36QUTvWdQZydJcdQVmoGYPIy/fMQScprFHuXsW5HhZdJ3
KB05L+6zaixtAonqqO0wS7qAQ71xrGxC3ZhRZdB0x7DSB4CY5FN/lT99pNGM/uD8
1sm2GUc49ubLwS4nR4qgfLP5xkLslY5FPYe0F3GUTBWaPQxaKOHEZx1U1sT588KW
J5wpbReNwlwJ8gJR2e7yzHyYwIcAF8+C9iXxN5k9v7oafAJ5V4Uq8UR1fEiofE29
D0/3ULPecp/nF1j3aFpSIXrzjCY0ineW/5JlNef4M5Ocr1viQ2CD7PzohL/arm70
w3G+RruOnGBcXXjL+0Tz0SICOSU3acxFPYBjVNwZdQwADF3H/h9uV86DeVLZ9ylY
SiNz+xDQ4gwfvmxVbAL+SgpWhzx2h/ue+vIbfky0JlFf78c6EXAb9djBbj7Jfolc
Y/TGrDQB2aLMik2yQCAoaiVjctICbfZ9N4MSjy5fH35QNfRj4Op9FDQUlnfh8src
Smbvkcwyrz2YdAWpoWhXeoIIxGBmtCHwYRE5rkjplq0P9BC61NWoKGHHxgCBIzHX
nHNA4IdXrCrUW5Zdqs67e28UhPCWE3fiBIAkuY7NCqElS0L7Ch8ekL74qaZgNMKR
GnqAVRqv4H4waLy7aeGwZKUP0MmCIcatThIt+RniMcJh6dr8URGL5hReRVBjbUFx
tLb2tzazGKdMrom8TB1pDFyPCyTa9oyAmRNWUWxCXwclzcJ4wac2+1/iUgyUEmv5
yeZPhuZ2dJr3yqPbGgY8seg5DYoDCXhw9yeEEmGDnUUU/K+1EtoY2uBXMejWj8ca
SbKyeLidBIND7yEy9USLkv1aceGSLaMPXxYMsLWKN3peQ5181I4CaM9LRTkEhCyK
qB7r4gHZeAjk6SRqo3FdYMaINJfyeMOMiwZ8Z7RFza0AyZw4xoThUT7vyMDevWWT
nbzMqhno3s3YZcrX/hVCRXWm6muqkQqY9DP93ZWRp6IJVyhm/yPFAG1RXutmQDOK
+HZt8XZ9uGAZWCz/FCnfaNlZQG8Y0y1+23xCz46YAL9Dk/Gtf4oprRbKQnsXDAum
RIMFEMczvjAadS/6p+lOQ7twITfPsWMxkhv8WQksgAfbW/3qbe1CEbru8GGbNn0t
ifT1GNTtoUYw/MIAHrFjcBkCIzp9xCEHKQb8hTND5f+inScUByohjX4lvioC/z/g
duvUtzs6h9D+gveRcOBiVi4bEjmn4U3dLr+el45qDyl+fBLvP/yQ23Ie/a/ogG4m
ZN5u2cDwD+rEaShSD5ZFD9T5giU1E9ptUTjNl506/0SLMDR+VQtsLoHZgqAmS9iW
1kUYNfKxhnA7dM41DSNMUnFhUakKlm3/y7kAuTA0UKdR6SjKdXNBzXyI8JnBnQZq
4eCXPly6BcOqnOab3oi5N3OcArVUk8bb+9ihgk3reTLz6ztp73b2eWNEbkkHsLcv
0Kv9+JjvhcN1XccMMcYIWkjnDWk1dmiTb0TMOQsNzn/TYSQ3B46/lJFJRNmOGpBJ
EHC/aP2ukh06fjjYboboDpcATECjSKG8mqEtaxIofSchZt7FSASWgTHJ7aXiGyGz
SrMdCKDzNqbLBGrW0piySW+G8d8G67t0MGvL7jVvkSTOmsg9Lj7ublVum3uE+yQ0
9RtZs0hyag1lt0/w54b7UnOezuXTEjCThY13SW+qTJGoB7DHtyY2jjsJNW/qOtjd
EvCcbc64B+qk64a3tQI5NM1GvQl7gf37UqF0SY8CyhpTNxyvDU10tovF8ASdLLn0
G+gn2gM77BkDfh/5YSg0CMc3DLk3BViuFVQFFELFOtR7GaJiaIVRl2thkBJhQTKF
cbr+FRHWp63OpaHSDoWzscVYiWDQbXGJWXHRmCRzAH9jYrWl7tVAp3g4unkd7qpt
J6eq4XsiLTk/3OyN2u/4L/nEYjRxZMNwGkAQHO1M36N/+r2v7v2gJQDDSA4sHQgY
cdd3H03cWl6O1I79feuu9ApyYpgLPUDy4hDCOhTR8ysUHxCVogi5IU2qmfekXfzI
wDzeXGwEg7OMg35SzXfIhiH6qZx1wz+Mrt0/te/LhKOItXyaQUztDYiHp0m/TINx
tqYrgJNTPXulrV1OqldOUSgF+Nio0VP7jKGpfGJj9Ra5gVLHxGCiUM94oY7gINF7
0RaCr9V+uNKy5WWg3Ce9LDtRgn/xMZN/oG55Y8wzHvgJLkJZnehD0y2nWZ0QC7kU
mZZ6uSJM99L1VyqV4/fLDLpub1gjMmXrG+UXCrcqe1QE5bqf+6VTpguDOf5yGcXs
W8d4CGFuashWM+HqGYo2hM3EqNiHi/qqmc5YwvaLFQVDgFQwG6vRAqh0p7/4APE0
wDqyIuPV2Ty7fxeIVGSf5Kshy0a+GjxTF7EgcNbiAe6zsSjlD5/9mhudtklCJyEr
5myEklNe+hzkg+Kl26QSr/Z4xoE9rzcrg3FV3O2PwTuuJiYIZlVdtK7I+Zgkpbw/
9S0w6TJ5xTuWF3yYlV/Le6yQLDPCYLPXEB1nuso9OXcjxHxckhk8Zx2pfPiyRctW
h0+s56IgID42HTkszXjFJBNbHF56bUPjWAWJRoW93RFQ7WteAzxicVLOIvGSlHtf
P03pVMUF5TpkNm5Ze+FfH6DXokjH89QCdRFv20coZXaGBU9MSD6jJJPMtykV+Zwc
jugr5DY2McvyHpFEOg2NhKraFIRK8K2xelE6DR2XmVjRSZbybCi2iF9cYwZ4EAqr
cy2ALycdm0UUX+ucxN2ZE+m7xZH2YfFQ+eEUa9F5HmRH7wC4pWZvmWfB2QCX+aKM
y9lVP5h8/0uZfjB44G7mFvewA6iNT36lf07/fz4kHdUzYg7xn+4dorocBrBk+jKz
ojoe1YrXdB+wq8B4alSQJObXoza4QaGQiDMCKzojuuLZnquslCAIF98DxY9HPe/M
XpdpEDG1VLYuuR082fAkOOzN5pm6+CFk4bL/7JrIeQ/ZiL0OINKXXrlsrK+hMtfi
HYDKbwG7n9YEooH0qDIKS2uUPZAcTdTNplV/xmgUK3E96yfRC2sMOTxwc38OfnY9
FuJ9TJ0pZG6nCJ8jzpfna+AJgiUWf2HMjrIQphDJAH/LYzlSjHRWdTpmlo8BPgXF
G1HBiExm47AF3bNhY/HaDZ/FD+Dr0cdy1QLd/nA6wMHu20PvTvD6iIHphZP1xVFU
ctkzvZ1lI8T5eVKg6c5Cyb/hCRD7DawxdGtuGo718+qaspZwEiupnedc0gSCdaxg
7BNm2ZGYxnep5adgwy/1onIUCBcLX0ZoDEOGOemZ8GBARBGQ12+9nMj4YyLVxJHC
QJNhH0ZnYDeczn9vENLCmzc7QRL6eEhLMKKWiEUAAMyQwBzE1NpkJnBIOMEnKMvv
NH5wcADzUeHp9a8SoTSIZwci1hydgvPEhiN5p92aqACtkXhNI8EOMU6n+Fro2jvz
/cSaUxqjKaZvya0LsRVb6KLnU+34llj/IAzRtCajtZxzsSCPmjyR6AMGgFYY0J8v
gywgMofE39TZvscB6cOJ5GeXEXdtrD6XfxUSzA0G/48iAWzzgVb+35nY/5HpmkF5
Vdok3CYh5adHHkocMOn2TnrJoyDgo+hoj3M7auZygoH0oKN9y6lRfsW8lTOisyQh
FK241ggkN/+LlXISz5mSPxIu95HBCRvfoE0Ow/K5V9722mBWYecOEi8w4wMLLJQB
ixTzg55Gd7uiU4bbOMfb7WIkQKhm4w2ECAE+euoCPXK9TUCV2bmR5hmg5XhhKrPF
smTmNoNvPt3a2/Vkt9Un+2W+RZUZ10/YvP6ePG0WZohu6BAmTj5ITVL4V1hpg8A3
/tWsfyFsny2MXBa+p/GoWF8hN/qk2W+qth162r5anfKqAnv//n2bC6nxFbiWUp0g
Kr2NTW3C92ebEQiHTRQt5DwznQEgVPM4M/TPzB4ezchKkoNBLLxKSVUlkJaH1v+u
n3+OA6kFyL/wVgGCAtRnukeuden4FFeQbdqSZP36STJVJ6jLaovcIve2hgwxxlbO
2JBLHKZe+p7MnUfEfyGzb+CN8nIutkfM7lbmsS8mkGuqJ+WXhgcxaPP1pPPvDoIv
tjCwI5LCCERbA9Qy/JuO40CjNWAHRE3YCW2of+pHTqGO3QQ1Wk171q8f65E1j4Vr
xLU6s0SPA2/zNpasfIQ1qIZYVkVQrTi6a5+8YC07b/pWtDbHozTNE8Agj2+NtStn
xiRgwiedNee6bnUP3GCRlGOKlYRiir9eoyZHYXuMJzkRxPrIiOWmZzXCmzX9heKp
0+Uuq0SJZHIJ72YRH3Q7+iIb6JOhMEE2lxR21ubz1i/fgQXydH5Roq8C/rWOf8Va
fJnm5ZyGMzw0EI7dL4+nP/GwpD6td8lSuyEoszzdvwxujEJm4Cg+XSAr85iq8XXy
4Gr2Ny8LoLGVtVL68yBH/DPsnINQpwKNofN5otcWvfoENHfjNeghSgvxVlfdKdEW
F1eBrPUcvcflbBM2qFc/0rZ09U8URSaCWV6c7DOdvxFCE+T3LeMtyMf3yPfr7oU3
B91DeS+DRoBPHmSUH7AacmKUQNNVjfqEypa46q2iNfayOgThOofJkI2/fsQEV+8v
PRH/WN31ue0MXMn4ySm6XZnuWiAPw5WdX9bTQbMSHOts2pFOMJ833Bp6nU2Iw0gI
k6fiZ73VowYDOy3O63fkQJEevEIprXSoiWY10fVCBYWyv3D+zs0BmSeF0wtoCG+k
Z7+iNDD+hEfI6PwwLtWn5OEBS8Y/9iXj+l71SwVjzLSpSDH5PtvBPBn5FHG5YDLu
so1pSv1Z0o41b46WS0nb3QARYl2BgU3EFe3K9voirB1D8EN/bkYkkv8rLmnPHiZF
tSO0ERCUG5IZX5ir2AxAPyt1uXo8QgrDHu1AoT8M+oroI18xuXmEpHp12Zoz1gsX
hKjaw/J6ogpjkTSylyRn4Z7JnBh9ou+vxCZjspXyOjXug0iN8qrA+UKyLKqAukBE
KohT1aqiDKXLn0DH5xNiezZKgG7euSEUS9VGTop5i33uevxSri9Jzkqfnv1MF7ir
C+om3ejs9OB54QUdqul8IUnYfD1MJRGXfDn2tVFP2sRtFSBnXyfV21KiaAg/hzor
slQpWn5ae9jvh1vOGCec06O4mTJNhNHymkGUC7VFpvsHz/Oc1/Z3ZXbemxBmGR76
gYuLZhvLgRChXh4evAkZjHUT5SPQht6p06ppzek7+egIgieNGR9VUBhpHUb94lC5
rA9OWwGOLDfYDQAoxgSPybSSNkeP+gK0Q9zz8OlHIgzDIIPbRkQ6aX1NVFtIVjm4
zUeAjo6Gt7BhWbAmiaesxlqYYHQBZx4ulLFN2AKVb+Ng1cfx1p1X+XhD1xQh4DkZ
Q6IReXqMVOYJBTGvffL3wcHG0kbE7Ig5RX2Ge4Vp8JJCHETzTAn9mRll4FNI0pCn
Bdf2NRdBY4nmPrPsCYfaeZcBJsWrStHV8RxrFcf72HH76sxQDt5vOfToKJp3j5dY
XO0L2RbZEcuvevXhPapr7NVhbgfudksgUA8sLLii/eUw8B7tkle5CBdceJhkvRss
SkQgT5Cd2Vog7XY/7yPIF4iIU9XZqQeAOhrkkudpTee9qFKGJeMR9n+s2jlSvZ16
2RKZfCJxAMJufZy68UMjGaXvMKFtM0gWXZBDdfccgYLVAmja4pP7aDJAhKwgoVUg
w+xAcp/Ua+OW3uDJ/GpaTd74rQ3v6CebV5t9lWsj4pzAR1436ObinN/9v8nE1hxl
ry/G6XPo5adKWYAxgGWvJ5Qc5zw6NcvDwoOhTNHmaAKzStAtOvAKpKeZ+6SXvMi8
p0LuMYV7lL9Swn+MmpLoJYSJMyW0GkV0nKa4LQHS8elVQkA28nSCRYxjWWCjZrzj
5cxYWwkmU9EqID/3XXARJL06y5SQnAZKhAwnyEKeVMcNhOFQYHjfXbwnMVOzO3D1
28IvCbxq3IlMtvtFUSbqOj7XPoK+V1SOoYXM0q0umLJymBClijDEg9fqlfh0G+EB
G4vyT+KL5JYgeSzfUIEY+fII3pJkxO/GGdBML/x790Ev2DXkqOsbFR1bsIZlqbGJ
eCth1C6QPnMDRkfhEwh5D3d9NGVU2s414IyYqbzwZOHrzRPaLFT805rupJx1BdeJ
u4jLF5i/jchaXmf/kv5rNBndIlRGmb4x6+BYpKKDHpn1J+2+RkdPabV5pWa6iFSa
c0V/EWMr63yIJ9l/TrLOIRsMJmDZCoWX0XwUSzBt2oCRKKf/FaZvQVIEIV2rEfde
uMYiitv9UdwJq8oiLFp89ksxWmIR4sgrUb/nXzWgoKJP5DMj0BA2Y1/jCiYiPblH
5bexmZDk0hab8jcyCDQXqJ/w4vl1wRV8Kvlht3W82/LVmcr2Ha6fbdotbpSfI7Le
//QBfOXYjqoPXwhxIDr5ImDN5QHCJGpOXg7vI3yUkkBPy76ZXiMnhI0D/u7vrgAn
5ZCl4EK06MpgmKvGH6aYMnfDggBq8NsNPFkqqD4QgDoAbhLsgO3I1yH+6WibfdEi
1KO/GQNq+3FFkCOG5l8i9Ym1q0M7YOp5aqcHbfo5sjLFa9wiA3GeoWzvLXSRb62U
OgVmURxBkQ2mNETZBlTgPGNJEIiE+5IDtp8U88fn9w3J49cAMLtzVJGgqxwUKVfc
qg6ezfkaoPadK8/n0VAcTSfur4VCcWS/IdIiicn5hw6rV49M3hPXoSH9fQ7gXCQ5
QMI3HSAyB3b6x3XJjUFKXATehOhinWie2GjvLRj5dwEawZP+56Yr46zrvU3qO8N9
4lRUQtpEJhpbzEdkz24msT232MXrsTTFaBHSydrpy+eHGYhCdlCoyrVMytIYeV9P
wQl94dav2ZdrFNWJyLWzo8j4Q4otOrEyiHhPvj9byTNOUIYIyL+qQ2CfUIF3UtGJ
m/0M6C/HrG7fNK2sfS2+1VhUKvEYFAgWX8XsaXmRtHZaOvMeHwlItDXrRROdL2yZ
/SBjy4u28r+C5HJn0KyxF9zNwarr+jw3TcdkgNFDb8cB0sI3u7aTTQyAblXKdrrm
Yia6T43sotNP4Ja8F+yALsA53dBLGaVtxkhqH17kewg6+ZylMKky8Nej+eOptnx7
QETnC6hYOaig7hxUtg3osc0x+IRJ7fJnoSeeoPX99AOHSaMj3zzmtqjGEp7HqkVF
d8KM1pE8kXcCf5F4Kup6b8nTzQxBlf4I/c4FnGSRkjOKnW9l+1KVpP8Jb+iWvvNu
FM7Qrztxr+GGwFMjHimb47pc73vPjXx7ccp/5J7ygZvDdmUgeZs3cEXeFaKe+6eS
UMKuRbfppC4vzvTckmBmEnIQQlnRmwy0adVi8WxlKicTjjQMCsK/P0q9w6OR7IEQ
+qSFT48HStLzs8RlbeM+xHJlaPNmLanSVQJkw5eCZ/14tPP5Ty5gy/IzC+U09k6j
/EjNRVacfz4hiIS7IWTLZ6iave982cCM8nvb+VI3OlsMkB/pTk35jgufMT2q2cwh
CmuKuZTdLg1LkFqG4RtteUS7WLRzhbt+NHpkUWTI2lYZLdgY00Q5TRQcKLwFp7aI
rja2IDVMaiyTdN83un/Z28rFvvYD3Uv3IYApjCVTOTo4mMoC2n5+froUCdUXBz/7
jHE9H1OhEzggaMId6QCmXYYszSwD5GSy5mfvJpat//yZrdjzCcqQC1v6DGMfk0gI
gqVGh+sMjfd5GDVigTw92Y2FDrub8UhAvMNTifYXMgQLT0/PzmTKYJJZkRv/E7Rq
gNCR0600+TvvTYB8SnAET2z07XKx9F7TRPDe19iy9I5w25eWgBYQvgHBq9qEpSeL
HD1Ge+psGpEHMuh0tB7giaqB+gBIbX8BZPXdlYWqdRUln1EX4aSgUURABvq0Jupx
csf9T27CGCQKu7Fl/0UKL6zi23J2er1rNL5TEra5sYQD5G14XTAAs/fUgQJHLtcn
NB5MJwU0RY94lUyhJqr3GTyo1RXVTpzBNI2Qx8iUKFyvYunsboh8SU4qZhBFebgJ
CtHIyNWh7UbZg9S7s5h3/l8snAOQE1uhm9nuRFHXsJvA2A3QxJcMVhoBNp5UD7Qp
MSMpkjBQDhLJW580X8yz386LtC7ueMB9VTr2UrXFgLU4uvstNiPbKgKyR4DkPJGi
9KdZGH/SYbIIcF87BChA6Pxra3SREuczQ0bvUQak34BAt+F20LGIde2K4j5VBy0R
W85RCWOQSzhhu8c/P2dOP12FhnjmN4P/+AFpCL5aSR/nLDqah44XP2D6CgdjID22
MLmqyOZFrulUpq9LmvOIZmxiuKDpnPGU8pyRbyLPIHXKEQ82p8ATcB7i4c3gF/Mi
u81KdNQDrU2J8EzSaPL3gkwR2SK5yLVq+t0nR7CXfk6Juqzyh5xkXRGWjJK4QTe3
4/uCSToqVstHPbzMc7wubP8pgCiXFZuuTFdRSv7CuSe/uXcerQS6zxy6wpaAncrP
YSFqy+ubs9ewlT8sjR2wg8Ech37JVFBnhXKDnEKBDaOhOQ2AbUrafBDs8UkmhHr1
nCNrQl5XtC/y9H6d9Bn3F/ubztS6Es0GpD2fCasfXrTn/VJbloXI9Ha2nWMZuTG+
N/9yJYdiGMHAP9FoedfjjoaYDEAMwh+Um6LbMtAQGb0D1NzjBliXNXMYMX3cauIH
IiEc4LsAmMYGRXstLbowZ9ZYYaMs4+xlFzwz0wOzEZbek0G5dfITCLjsoFLecqqT
Kab6Civ04Op3kYbJGl4aotXUmCAGQePKKhwP9qdOJSynW8m41c1BoOV8mIxWCkZ1
KLVQDXOu8JgQxkKb4FfkkXpji9w6+PYQv8+K7c93qTw/QhLuqgyelJNIluqga92s
UseghtI0QtxpygZmlLGzkwVUeyYPs2gFyaPKr3sOHhD+U8QR+Qz0tO7anltXH469
0h5ATV0Kvnon4CghwJN2kmNYTdCz1JfJwhMc91tbhqHIUDk9F4LJn2MBULg/w0OS
hg7Q/m/Pt37RSKj0llUjF/6z8R6OXHJR0hXO43BxqszFRctZTJKDRlYjGHOybH9G
aGPwpu5XEyYaSOFVFJV21I6Zu0cw2I0pdQkaMqhetMMAfFE8r6CMWMzPWmBJ1K1z
g7VcyH9AqOlXtZQByE30kNAnoDsYfLceZDPO2a9pNYq0Op8gTMgobesOvWTXI5Pq
T34s86oo6ZGQd4b9Hutu/DamiGyKENO/pFoRJ8xhoTIm3H6VXp7zHW/TNMaejbXp
a8E0vhAcr8QVmyrfOCSaJ1bTy12gSNNiGSOaYxCyYODzoDlIfeaXyCKb2cfYl3/b
pAOKy7ZszADwyfaMRNV3/ZNJlLzyJkSb3Zhoxd640klNQWdatsy4mZGIJJ2cLFyW
PNi+j2ycowN4LpoSR0BJV30EhZ9LLQrKRgsQvWc8ytuER6J8xDVdCgr7IYTPrORa
PtGADhwsvhyanNerbTJTByEUlfiUqrWVHl6GfZebn3lfL4Lyck/6iua5kv/XcCdA
Ajp/cU8fXDWjg8JW97bqMMh5EJ824fyZupOy++Fl9HPTytqo9S9tJEZMgK4/NuVl
1LAyDINWmvRmvp3U0KAfq4KDj4qgYkMA6bZFw14U531K6vF50wGWhG+D8dpOtq7n
FXZMJLutA6K7fXDvfystF5rJfXD8JH9Zo13eHPT0kLQ5AN2Eksle7J9li3iJh385
iH2zATQ3MUJONZQDjizfNL5zTdA1S7RYi+HF46MwNHV09KbPQughYvKxAdmzuTAl
oDcqa1zRayNp4LdklUCEt4+P0SkSB1lxtfRPsQAc7ullCrVXVgS4W2m1E5U2nYNj
1Lkl2jjJ7/glqD+mxTbwlo/YDLjQXSQLvwlwFuXicNWuhnCrG3xf7FHmqLGmQz7j
jFwIyewhXiMSOr0jKAqU+MuhlvF3g9CkexpflQnWIgfHwiPZDiwiTfET/LXWteAB
4mubLT9vaIkAbjSXqxeW+8O7zbNCKTkjN0DfmUQDuVr5r3qGjpTJhey2iLD3/x0M
UkCvUbQewOnpeLJxG2kadsUIEQAda+uoIfuM1liyo2ktqC/fH9dYAQBmseO2pj0u
FiOydaYQkXffzuewTX/VHGrhLZ69FMREnmxHbBMihR3PNYch7sEIgA8htHFSD0rC
8WBXkrmefoEs1+U8UKhYkywblSz988Mu7zcptdC0kYjbhOTjII11F60H4iFTXCiy
+swsv0lm9pMmHO3rKQFsXeSH4+hvcXHGPS4lCor+Fcyo+m0gtnbAq/5o0xajd7il
l8/j4gHXex/GIjwm5MLvPvDLvBF9k41y3cWWzDe8clu8Wow4dqajFW9L8rWgv2aj
EPwb5QkqKKEo8pMRHuFh5Ohh/f2kRqB7xaj07WoBgj5c8zieGxTQ/HRBfmJLDLY4
OtwGtZpXmt5Zplt/hYMvc5WYjwkwwX7dd0XxqQ7epbXa/7VwkZAtqjTtU8dos5KA
OYs1rlz8hJmKmNAolLu4u2+B9wBPCb2UYKJGQutNaSXKkN5/UVgeAHusc90NMhXW
N5VUO5sAvKRKKObslfOYNbyU0bKow0quVtlWH7GVTQwZpfZ2ebUJnnDXDV2rOrU/
el9XmqY8iIMFEALSzUZAoUcZ0RBYXuseVo0dz0GvMtOgmoafdplCHKULv1FXcrU4
ZGcIlIqNgE+eli9PMPZh1gNBE1/p5fJQm07qFxmULfpaiwfhWzXTr6DvNgz3a+xJ
PX3CJrHjUg4Q56GRlDGTiDPjMkMKwHzWRYfFltF1t+sA0T9Y/qjlZawthcgic2AA
8x2WwJcF8AoFHEhZL7QlxzGraAd8bai1vBYGSs36m6UgMmX5p5HOclMSvGherLUg
COhL9ihqL8vYaj3wiSOHYT6fa4wmk7187AoM3mZ3BxEJVTSsUx7jv2fdhcPIrROG
lHIL54cc6pccS+ihUf7DeEFfjyE9tVLlYwLysK7DXaHQcroK/orhGOllpFMTXT33
tkoY52F2YhxOhcPWuF50Ei6T7fAPtFkHjf0CKwzcr83nOP0oKPZrnO9or0H1XGDV
txzAhDBdiMXZ0Q5ObVIoiVTJ2FA4AwbGZUqu7XHOms/rgKLUtdRqqhO902e+O17D
QXMghYyIxqj3aUZ0WuXWoxbovBYhlFnWkWrqnv1H4y+9HXcefjhjLdELBSszRQP+
fKqEIQsn913bT2hI9TlYD2vFsM/lTuH7BI2bCg7JuMWPpz9+Sr6LEqF6TFW0AHgG
Y+/ugUbQ01RPPFpqx7Qw0cLgPrZysUIpQ7mMQN/UaI/OQLeqhfyhUg6MSPyibcMf
Z+YyDQtOL0w9JxPnRRjFw9jYXxfWy64csJSLIZrhMDRgtt+7t4bdkrpLOm0zxsxe
OEKiOBt5V4ZpHhfZ3nXEWa2JTv0uf+TzkTflDslVkMe2udnzF6Ina/ybWO6lIS+S
WwnUS2YqDRehfjx1aqvXbMAuGGVG9WLr7pwhku4jP7SUjTqVjsjqqt4e9PwKvnnN
NSErKd20wpYibiRtHHMe0UWDd6sLdPVWQ2WZZa9PCDXcPdaNfihvnGzRmLnbqZQw
CtlIOjC4UZaaXXO4NZu2PofFTYNmgldT4tJUI99hz/lDIY9/aHMHtdugwJYWafIP
F1zZyTbSRue9QuaGWEcJ3t9wKbfBltDmkoWMiIidTEHm0oUjsX2d6SmwvAqOE47B
IM4lw0Kx1ZCLiCLeiniT0mr7VP9ciu+UsYfGHNhS6XDdL4hgM/xUA+GtsnXiq74r
FLtB46yEJbACiXimv8kTctjOOs6+XrZV+VmFfZPPbLmqGsY464AFpmHnnSXvZgXs
MBkb3vDI+ofnr0FAburK0U3VP6EQl5DcEIqCOeSb0KxcW2IAFD0kC/3qRQDR6mIK
7ll1TDAKQlboZ2j6yPmrJcz2eI9KXh+ida0xwoqvbKSmRmHjHTsfd/fplcOQONw/
JlYnKagkJ3SOrU0SWTRxbRkMgGPjkGSy1ABMdxxVAg69Wh44aqRxRIfW40CZrryC
9RdxM2AaxK0qSScIkFsLzaPqyckYgoLbMY6iwUjx14yUX7WE/A+yPhSCQguk7ZFz
+SPyQLOhDZc08LIwf2X/r7dYLTmyvrRRifdrzrJrlJmHzUV1/WFMhz0SeK3NtXAg
ZQvrek2qruaD2oodS2lKv0JGptrUv+jHRuPRc4huikDjyXYsRyzwhKGZAmuv/gS5
cnw+O/gNhvnkWk834jDBVgBupVoIBXJ4XjD/jFx9Cq+BVULmsghman343pqW4ifQ
CCMX+8Vl/6EqS3uX7HGjwH/o58LDl8U2VEorHz9WoSB1NpVKyXLkOgzUHD6iHMDx
zG4teV1qUP+F8GDXt60qxcqp9gMqqBVsu5SQ80Jn/rtrX7eYE1z/8p3B8qeCME9F
UhbSjJ/jKtHeBXve6U+wiCYBz2yboSsu623G1YhpdXTCbz0xCYXJt6mrkuJt+MiU
9JWJrfXY6DIY6lUjh71oaVR1TNhrPQQ805Y+lUrXUZYKBPW2pRmUZU1f3UyX4pi1
ZAV/Z3cskdHM8S++Ehvq3/hQQEGSv8Hqd5gA8+IoVfcGN9lkz0Gzfibpimgx7+rI
r4atwhtqzOSH9PCw9JOPMyiK2JQEzRFue0lH7gwKcFnnP/Betg9GreowADwnXF8l
ImaQALJHbezYf6ggZZSSiw9uX9+477qe4dS5HVSsO4OrSRsOf/CMhP4q5ShA4DOq
aCAHqlyBDG28aRnrpYFbYbq0V65QHi1sYn8oAcPpgLJIO4rCq5mPodI/nne5M7PM
3SxviqCz+uMeEbFUfTvhyZdpyny249wjcCDNmxhYYb2LZgcuoMzNWJaNlQ+BMIki
rgJlW4cW1ut1chYcjB3Hr/xFKnv50TfUEJYP56iqita0uoF6GWYHcFGNdPTpVd55
uOAo376ohNsm541thNkgldcO6Jb/5dTBEvjzLP2VYUQlI2RwQ0ClwPsQSdAVZ4wZ
HWkwvqWqlDmlDfBhKwzwifMOoofWzRZLGxVbUssdkwNgw4ykAenUSGWyeJjzEeJW
olm3d1u2j7caznpeFH1WjqfMQqV2G6w7b3LsFWWEBQSJAoZbYiJza+SvCm+OIddb
EI82rtxuVOVXwgJjE9LFh4AzG4KWC3qc2Hhx2S3oPI/v5yOXqAuaHD/cTe2G6uE9
A1ZO22O2In7cbmmPtGuFDts/Bc/rwvx1E1uzIUZigoXGbZ0vMftEo6pBzOGh4ni9
8i8SQR7JbKuZ9aRjaFErq4PSpqE8rBaG/8clWU4FfvYroVTIHZcBXl6Xk9FKds+e
gf5qqsSDnPLTuXjnZpVGcstcwbVfdUGzKaQw5zjcwDm9TReVJlaMttlBMCR+Vk8L
xQEZDhaCAdTBa+Oz+vcHfOuRsCREEblGEwc0OXzCsEsws6vJb6T8MLfKVfEvnMg3
ytzkvB49COs7RMsvhlKk+79hO7f9q8CCByKJ76wLu1s9iq49Zhgk7npFhJH6otNs
xGZD820KyCgvABiTe8KF15pFsDnqfTKqII+MtrnKeSLrZ4B764Kf6w2mfrCv1FS2
O30QIaZNvqlznLCykWv3Tu4z+9omor+YXSHfQmVdQj4QsgDXnppFw699cJFhv82d
j5INWQYQ2b3BJZLAUR4gZ8urn+rQbLd/04xkYZm1x+er5K3yCweBvSjmDOGGSxTk
sz7Ng1yGZz3FKFMm9wAlBQONn7VtRrrQeNEHbhZO4a557uWib64qVrL4Zl1rq3vs
QleKDI2JwKTDycijFYWwqUPw7c68AInVjmHeHqeUgrdDbTPvLU02I18ab6fpo8OQ
VWbWoumHBKds5LgCECad22X3stfLj9GIvEJPZympRpAZjjlTlbauQ0gc3pIlA3tZ
IlM2h3+A9JFUZRZEawUFdW/oaA/i5aKKW3v9DW/P8Ac8RuSEVUt7/3Nq48hKnHZh
DB2XpaGUxiT2GSdeKszBQQc1vSjIapMaoAyAo75bQtjTwM0LybfwDosraiBmZ1N/
vdCVruRlq0Yf6JLvBm3kZZpi0a9idZKl0o2vAArhW6HUlSz6FmXCuMszJ5qMhG3P
Cj01RfO0XYv5rNogYmoZ660tmw8MQ+s7e2+dS8Wg5CKva/AYOJTNkbGYmRXLlH0r
9Y8KO8L72wUea3m/v8hqbIU4V47RUwhPmr8PQ9waVr1/gUjZ9MUrMndax0SKt9CD
m1OdTHE1LVX0qSZyDIIFd2xtQ8/p/IitvqUmMR5PBMcy8MymsENIQdJdm+Cx0bwB
ttwxhFDJPRjV4jhWW83PRvU67ljHHd937TfWvgjjEO5nsb8wcC21/n1osspu/u4O
GStVJof+nUlMF1Ue5pEgXsaqFmAKTCq7/KG251tW1BWwlXHWdAtyTfAW0zCcfM2P
KnrOR3fOHn3U9wO/NMQXjjLsZJ1vdfO94QBjKtroz3NPGgOv+rwYcxdEmgo/Xx1i
YFQgswEaQWQPt4geAsDUgf8r2TR3I5zR6BNRW4lA/nw9IkR6+KKmaAl/vHsiu7rc
jcA2pjMqGuKMtHFAwbA+bntcp1vUjIkNVo1tLmwZpRTvnFZKwXWnk92vOsEyNW3f
pUee2j12xb4eow6RSQh8w8zGubY4BVfFGVibEEAKQtLc2TDU4QL3fQykWn6SzA/4
S/FjbfsFiKqxQgmtbeQpcKtP0dQbHyetnG25skFAX1MZRo2eIJDf9AcpvtoVqgoJ
kQlxUXmAN2qhNuISRq+V9M3YBbwwmjtE3l17Tsya5F6RK7yxMVxGZ4CeF32UbjLo
jZidnMYuSrXUQmf7VWQeQetHvLuV9yJhWpHNCF796B0bVnb9fSN2n4J8RDWu7wJc
YeGTWCMWU1/FHVcRV2CLoRLjS/P2/UBFxkFDEc7cupGywbN0DQEMUrWV9IXT8wDC
W73hy8tz+otth144sfb5lXRqneOD3+RmUedeD9Qaag3a2az2bjUj1SuLEBuYXcIp
CZOEer+aeJrHh+LIsgr6eRKEVdh2mQ7Ad+1MYLeupudo2D4px3x0OZ5KlJDcyGXI
+o3gYFlD20W6PUlDuCDFb0Xw/IC6uXo5EfJS8v9l4PJ7pwgvX/WOXrwE5nWpxaCb
Lu9fdhmoYhqcpDJOj/hKfHI04C2/Hn28tz+hDQuOqx96o4pAwe5bCUhvJ2G3PEKN
G3Vk2+XW3nIyQ0R13AxyVx5TzA2SQVLlgdQHDJ2XDdelPWEHvbHllklwzDhZnWAz
ECj0YubK7F2v5gCv7LS5W/zHhs/tNrIGDUkwOuwP447WqdlgHQNMIuB/OMq7yGSB
3d6xaebu08my1oAOOuRVnVELC/7yPacJUZ+Ut2aje4nUG/2Hm2mD5KNskPT3cgVf
Y6BwDq050oJ9f4sbP8fCZSd7rMZMSoUNdhXP2F/vuXa53eRa/il9CrlOArIXatdP
4ljT8XMY2V1csbJJbTXWecwAFTiMST9pZ3Tu75AnnoJPAXgaKgsVmWaxWpQnCFky
XDVmIKxDeqI+XBqF255pW2C8CE3FCZKr82mvAoT76LMLu2CFdDnQ+xnQsjzvfF/h
YVtW8FDy99jpz24uG0FyeoXMJKjxSSuloQ9eVMPXSB4ge54bsjOSrivXLznvY3Vm
7NpDtNYrD3jsOLe5FB825ob6XaujFS63xh2RjUFjQbh61pMJQglcfGJgPTSiNzWz
Z/yKpR6pnIxqeIhqP7IWWsTV84tCf0GpAZ54RAIyyLWADRB4Z/lm+tktOF5qcYWC
9P4olfoXUlZWNIf+m5GWvL6retXMEP0qfiR2c1/CHxQg8bSBgv76P+g3ZOTk6JqS
hVpJLt2CLoofYz3hiaXN9xzPyPwE/ruJrvXpxJWMlfIHGs3hppzUngRXjuSkl9r6
CmxulPqBKDv+u9oL8HWLIe6Bc51pd7T3pGonvW1LZLdp61ectz2B3tNuBcqDq5By
6euw3ZGs0BDQ1GBo0JTvN2pLaxW71tsxRBsv47XoyHWvKXvlCWatNVhRF9JbW0qb
NnPECNMZ8pRZLeU9Wh4oRRBhY0fCmBzfikUVdvqImV4t7xXG0ZRGdVrunTfmxm4p
0zfByOusWhSrUfnWl5wnNxRbLViN8o7YrLuYLeC6KwRGey03qYT0a/zVRSY6yYgL
ibrk1JlbudmCxwDScs+4j4kYbpco/5MGJf/hJCKqDe5bCsHUy5bUxpcp3itGcyWl
YzTayf4CKObkgDIT4k9gRw1XwoBiA2+H4OxVHx3lwph/nSlrT1CC4yvMHLgV+83p
X5iLOHrf/moJBEq7nAWhsUH/YzeM9tRgLYQux2ZOCIdOoto0VhC5G4L09+BLFli/
h7fpjjJBY39WUH23tny1bH546kQ1Mspp8nKsurdtz27PkyRrN4ziI6oIkO6jvgF1
Z4X4uoLPe/C1wQteViPbnQMChx+n3s2qktvQqAaw7tFN6RotrvTRpmBt0cPeDysZ
rEOzAquOGjF5XZaXaVkJv1Fu1KlmefB90oe8dpYcqAEJunE7Vlfn62VgmtMM7+sX
p85tPQSBCKEvQjfwOrSDSOsEe2OPScaNnjyOnFKdm6y+q9cK5Kq5Rj2hCzfu3XD4
Dj0GzoYErOikacx+4o1Ax8t4JmHzJ0kheL7MUDiMIUCL6q5B69fM+1tdsov+DIKh
zLL56wGQuhEdeU249QlZdtJzt1FK1R6TMdafQOktOjwD0SrtqbV4ULCxNoVPGiLg
eK1mPGhQj/o09sVZ3SsVZIpOp8t7G1dzfraP3qtQDC8ycLcN5N4gTxF0Qmq84ww6
tTNDiS7jhpvS9uM3IkM2HvdY+oJ80wiDH5HWZtIdxDhp2Be0zR3BTwe8NgvCkESq
Yj0kmCXv/f/mwtT+xaXbKA6EzBtalJYte6ckWigz0zwErblK5ulXVYfqQTs+7DUQ
RehLuTbAEJ4RiFmCNNaSReIGJxWyACu/kvXkwd+MrQGfLRdlCb3v9kDzaA0tRPQL
wnZomiDYBBKg2kR6mSjVQaGTjUHf7cllpHlB/fqjGKxYIDdhNZbVsBC/00xJ8Div
2Pi+crU80+SFgWgj01n1rkQFDsqBUM+Ig6QYS9vhiOU57A9zuSBskGjSSRBopiQ0
vpXjGy0YyGOyQW2HUZz1T+9OC9nhP+ex1CnXMYNpwdGopzix54x+e4W9K7GaYlUD
204TxGdxL6h8+weLkRV1KVM4eW3OO2jBUdZXx0/ZN4/3ixXgkSN3Kmbf9Gfg5++L
MUswM2wBpSEuGzw425HmKnrBbnvxGPrlgqtRnJw8uJyl+G5hPhW4/WWGuULB+sqM
dyoIDHU4+nYUYea8L9+3S2XOTe5KcB1UIZ8R92llfCIMkMnsHjVacKDp3M0UbJC7
4nYev2pKRAqwvDlFSeBusLYYvVv8dzZTg0U1gk4AkN47z5Ol6pq7UCHLymnG8RyR
WOguHQTo3ieHPoyiJnyG6+KTTVLyY4L8WWw5K3HnSquQ14yqp5HVmR9GD5inDKQj
4iqN13CZkJkplMKf5jccPfPPZvYthAxo7DN8srOlom4QfKR/iQ28bAa6kBZ6opfw
kY9xpNrvQxPrbb142IzqWhR15apH0JDji0efsMXM8Bj1k1ggAesaYXM1Y5bOtNdM
IcVnuJowcTx4/e04Ktt8EFmeZ1THCrx9YJJ1oo9iscSwrhZR4ThbGgtKVnUeislG
ahtbRkerqsG/hNIWesAqK7XjpLJr02KjfyNyeuCMYLxu4iey1kkNXFoD9ijJBo7k
Dkh4inHa2lspqVMNyyV8A7l7NwbSbFmRschgiZIQS2YMuV+EGW3K7h4Xoe7uDM8L
OoESrt7NepL8uS/A9Arm3mpfWF0/U9uz61xngaArYC+beXf2hdlIs00syZIm9cfG
KeDe+RvfZ8qmaJCfAIEbfK/pxKcXxV6JxU4wJPHJUejVXomhkKg/6vAOOVAOmpoD
94A2E2qAUIH5kg3r9AhGB6jg0S+Zsvw5wbDvt6u1M8aCsI+uMFy336T3mRvnT717
IdCbtYy4gSSLfLIReASwR+04/Fq9MfRSSoYy3XSGtinuSFeUj2FopsZGEa1ROt2P
WDW66kb+h8bry6udlfX0gj9zLs1Vcblc1WMLd6Q0tsZ/Js0Shpn7CjcBzkX9TLmY
FG83byyDOGTclTb9wWFHKj3mf+SrRO6ohgNND5h1k4MFtUEe0/zGUSmXYdUr6dTX
F4c0/n9swNueB/hLFGolHAVXTiEZZfSUpb5jKrJmzeSyfxcKryWg+NXB6BfBan5W
Td6eKjBF3utkQnPHR4fvQQNXMggAsfVmgLYf9N1dFxh8+y3Vnf3q2IjUPCQkTXYi
UMw5dUSgHkS13gAZa/0fG308Mh02yD/YkhMJ5CfhOFX0ZMz/5+6+c3qCx0t3kzxk
XHgRG1kGXOapv0gkx7eSWiFsOuXthIi+/0id9gQ4GT1J7vXzeNfWMghQb0sqZgCb
6m+ftI3zw7j8EimZAH64eoflxZGc183Tw3VX0G9bDk1+Ng27oml5+SOZ1XohV0fE
Mp6fC2aqRkv91eGc0PWrMzPxiGbEVWOTxLgPHcw3BKPoA1b4Xwolqr7zzquNlxT0
H3CyXJ/0iO1jKVIrgikOB3G5olH5kW0cHA3rDR9fzMaoNqDSZz2udTgWtWI44Z/Y
9M8QYzDdu9PWgF5FVNNnxLcjzOWkIivPEdn4AexfiTImS41qZJgQfoyfOnFSay2K
sPS4NADuRxNulK29Tkq+S7YdBDSACiWsjBtRmi0XrX2BEY2Gk2CQJ8HozLwVqFSc
DNfGheqJ69aOu//4bHbjalLKVF04fFedkAuR9y6Iy6MMvkoBMePmOOBiaJ7LP6/G
ZbUxpjo9GL5MPo91S4DIAe7UEAXweeZY7mIMk1685WOdEVZRreu3PdJ7YX9AkV54
LP2hxQJSoVS8yiJ4CTSHtweogkZYRLFRWu6ZR7D0iJ9M1L9hpZ+gsR/epdoVhN1o
YjCotPKrYT/oygutwTPEOnZrj10zSSlCNhzJqiIYPwiCgn53tsQEujdj037QDDD/
lIxqyVugsbB0Qwf4a4pQZ7U/OUWbUUrW/+tXLe5w6XxcA2RXm+sOBwQmdDcuOQ1C
P2sECMl3hs6Iss5zvTem4W6l6BpAoLbOyk2S/25NcT59sgVhE140b8KefynUDhx3
CR1+8x/CHbryuzVLKOMxdw4RysAy7ceNjQ2DSaFCMu5yl/B/hGAw0ZmRIDMCQjRI
NjVIT3hOWxzcMDzMTwHZcWQxZ1S4yRzF9+yGiJB1+MMietug9yV2bOnQvKYl3imB
TeEl4F6BmtnJvx/zZfeMMQOTfDWLSmG8Be8ndffDtl2HTEdKlLiFPlA1QhGq2Dca
zVYezS1sMAnZPYPhTmj+80dVfyK75KEdiU3q6N0Lu2+c2xEmVFb4a12Diq1Vzyyc
J9L3bRbRXvBtnIhvWKatNNcfs7vtTGPLbK6bmPB4H8wF7Kqf8IFT/d85aU8XHjKv
ILUtTrmk4aY9VTQRUcFVIrov6A0eu9MN4JEiDpgjc6kdiVzUh7gGyg/43kMhd990
hzJ0x5iA4EjAWyRltFOrs5Fx9v/+8LpiKXGJZe2upDqUha95YJvjnK+uN5QrNCSq
P3p1ZCdcQCfoyyAOFysMcHek16eP27h53KCX240RD4HmL2cZwbPT0+VWaaROv6AF
gGTO84eUSCve8maVHVg0tGvWbY01uyDJljOA5S/zURHXQGjaN+UTM8qgvNdOOvz8
AcyVVNZZBwitF00/ZfSFs2nA4u+q6NH+2Mrow/AEPSAi1As1o86WQRJiThhzsZ7i
nPdrmnw6fklBPvUdGWqsBYhR9br5kbUA6WwmGP+WQ4AO0fHtuLG7NOvr3KZJFj7t
8bt911VYAgcbMkknLlG9Dpv4szdXUSmy4iaFvRv4YrpZ+jQDGxYNRiAvJ1nRWQ0i
wS5SSK7DHm+aWpR4TwWsCrfVclSIF0Xrl/7sPaorqH0hYNeEui/zwQnTBvwi8aV+
QeSnlqhrxWTXt3krrVDIhHQWtq6pIQqTbXdxNzuMTkLYN2KMUYJKtWyfjtijtd5V
rNLum5qVuXc8pfbLph5tyLGygykLj8PukmzENQ4oNpEBo/xZ3fXfbBFghcioVrYD
i6jGK6pK+mnNussCQ30hXDIGQ/y9H0dgEKHUyb4gGQtzrIfJ0XwsnUmSD383sM09
nnqlSUU3aYb27AdRtvI9NKkW2svKZ6NKVni505NUpSdpzmKw+jOBZMkBVV3qdlcU
lcdATESZo0PCUbkYGBeHYzpYZWdizsVuxCzJPmDCyK1G+uXeNG3LMUSQMoZnScu2
/4BuvV3oxvxejpKVR1lrCptnmDBeDAzmLn5j5W4m1TUWTj8ZPmhT7JsYVkWcqS2/
C2lGEe1mcLaaST59Nh/f0MQgPeRFqegemdEFvdcr31/0e9Iv881lh/g7YeGUYvW6
JWNDYmTO/fi1MvwQIFdbUl6RBw7ieUcQWXt+mRWYbC1aGHDVET2i2goV8BpBt0wQ
pP6o88WLCHW2+uZYxzvdP1rXG0lDBmPuj1DbgeSGCKGQR3NGKtnezNC+wSlpEfs1
7e+lXBYUaSW21S75xPcgYkICsoSvzd5zqKukB4jHQSksRlwugWAkvLCj5sgq1j4c
9JUvf1zEEUlFNLYt7Hnw+BAYIuB+6l+w1RD34TiJgQoVFGI01F+XBhef4al1gpaI
q0JFIwHcOlDnyANX4P2RV+LGwx8EZs6evb0KVqQI7X6TsC0Zx2jsDa4YwOsxJI1B
1Yy6o2M/o1Z+cfTR2grQcp1jXKjvK6/Cf4VOYPvpmZQVKMhDgaSmofl9w/Tt6jLD
X15+SA+KpTcPdwh14KlOJGLG7mBPMkveYCIjOVe848ai/JmyivUtBT2Cs6nXmHAQ
QaAaVp1T2xF+PqBg1ypJ8oohKvbspvSPwXrR/GOJJReKD1iaH+yGE42LEiGvsX5Y
yFvY7AraEcL+e1lxXtzBd3qCG6hIkgPE4FiU+IVjm5zJ7KEj16fcOW+l4fJj+E1o
Vv2uoh5rhd3UaPC9dQKXbsgu9PXHfJQKPco6FOWkuUB4z9N2Ix7Dv5fV37xIQbqA
HD2oFFZNpF4rkDCJwcQvOyCEUY5Yx5wNxcdue4cusUHwJJGTx8z0dSXluAygMb5R
PH9Gw6XjkcLxxt1RzTsEtVsDIyp2haALrvhffs0sJSsRsM6fS1zwBCRx1hKfsPVX
+mHbzD9Yu0cmUWiqbioCIcSplybktLc4ftCPQd6oAqYA1FGup8m2kKJ6vOZ4Gi1f
putya9kLC7p/iWxbcjLIqOVIsxqS8iKhH4KAVhxaPweMR6xW6M1o/Atr5ZzIvblp
PGQnx9gVTWtSy211MzF68aVhwAK18DZ+jIa/5lNLUb92Z/SDV5vJOoQuYFDZXjNN
obJgs9rXQaj4+Lzzukh2rOhHz2d43tu7A0D4fObLXPz8eT0919ceBp+BnSj+fyus
xCs8u+IQPbcvnHeyvy77q/1W4JY6liXVgKIu9MDeU46Su64mwn7n4Ox2As7ZjSk0
1zJMozyIeW1FPdcr4czEcVXRB67dS4X1abrmd5bE4J7GEThs/IvmA/cjRqPBRdqr
tjim261leetk0SBTLPSJBakuCBYKiLVp+tUfZPKRe+MY2mP5zH8Cf9lpDjjvB1gI
h9HzC/8AihUHUjEw0lYpgWQU6RO1Ehx30ELkC5LnEFkg5wLYLivn9/pL49igM30Y
8WiDyvoOt1w63Zkx/VBpBJQZn+BffxFhLqbN2HQUWH4LSW0RvEt6f3wXm3VZyvIm
0X22OApWK2UoIOvvLqwxUgEDrRAgxPqt9iHiUQEBpiL8+B7ruDNIbOefo04ECAeL
9yxq7eqnDQvVBxMHD2uXZI4FD8/dt3e4H1aEThRu2mYHIXNY2UVGjGq6FGR/E83Z
Mlhnau9qW6+0sTJ/SLc4GAb5vei4cFuueiFNJcHcvOk26fZPqQd7fJZxMgdfewYq
AXqzozVRn2oJiGd6m1fC0/tkX5p78v/GF+Cl68ly6NdNlgS/87Iw8osDhKyNaq4b
Xr+JvdDkwZFSdy4u/oWg3QIivoxxJRfn+iBzZhwQMhdP/N5lZ8nvtNHPiMY5Q+BX
0b2gHGDh7JcO+F2XgKI8/lqiC/J2vvX6pYqghsD+pEh7scfjiwKYh2xNBpFWN1O/
W5s03fHyYmrvHLMzhXDOxJ+i7XARlDlt8ATM8cQjJVEIZGBnGSybCuZedavWJD7H
t/m7Cdpc0IDLdmkt41yvtVO5tjoJD6BBhY/F+aOjEGNDsLIIn3VVfTApzEhtLt+V
Mtkl3QWwEMPsaYiNc8hO1Rn8ouXQvyTUSKV4Qo67VPVxh7llPeoGEccqnqkgFOb/
SkHeF98FN6z+mZVuXn7Wlg796AyTYA0J6DnrTPBmKdfjiwNZMyXXo7QT6JDCabFk
i9Y803onazgfxh9EYnKxm6VrrojXRLZl6MEjA8LXsYf4GtmLXAhtaNlAueTfWF5y
xk3Moq6CafATxlhZhCFNFqdb3qazWrfeLUztdJUCgEDypifB2y/W1aqxAiGIX5AE
AgAdqczSJmfAZBngtRpL2fhGbIaUugJ9ta3bSmxe5DgEqcHXgdWZcL6ptCtyWnN9
2FfMdEGCp5W6hylaKYIV6DmYyrRDQ7En38nFAJMfXyheLDs0cK0EFsndxesR6+I/
Tt5US4Jb1RwgJmU/HJjK/9pv0l7l478kba78mwjBXIQdO/k6hphBoWEKoXDPO78d
JDGvGXOeAy1o2T8xO49FtCRfyYSBzr9Qyj/UZPBtUlukAyLndZ5Js7jAV5bVUii1
Q+vUHfFQWWTtBhYbw6MTST28Px7JXAZAK4qAQGoGFocjG7gihjXjCVGd9FXEMB8v
OYrW62uypx+VSU5fc+kds1lUAHya2myFjCzpRiqsNvahPqaUm83jOZXK+nvZt/mo
yee7FTSp4rDKI7dkRcPA5Becwr+IUctjlkXbvYZWy6AlGE8n8lI/SYf+xHaT6bpr
TT3To42cjHjI3BTxb+uqrXtUmD9G2OUpwDZIqmT4IJMuuY69/3qRitt4rkke+J+j
ar4DfrmlFAfQF5MY2SqhkkOgGnM4iyI9VYIIXO34Mb8fKw7qN3HarCzldxLgcfq2
Mqey8vWit9C1lgwfALQXGrneJ+rDgO+0SkV7LwhpOC7TgPPR6eE6i90mMb5TSPsD
W8AmQK9FrOTmLNfptGI7WEYHdCypeGzeLSf3kLOqf7sA1FZl8R+kT/1UkaxWrYUD
/q0svL7k7iknt5PybEA5+37eFbxRwuwKmdYPU/xa/I4TElVr/EXQHVPVYcPXyF7r
9in2vesNr1b3YtS1eHulMO7pZdcLF4oW5KczK+UiM9ICuHPF0CViuIknYQHdsqwu
JGA/4PF5m4i1dG+JJMfM1PMQ3IFvg88YDM9uOhBv6NgoqorI3j41PXFIfapiow2i
UXR27ik0lIoRfdgAwBQo0f69qE19zJS6+PieW0pKX4TTyxc6iKiGuqU4M9Ut5VH6
Q8JYxYhvWk/3aLv6A3+1zBaH3OvF35Xi4easPk85UAyHPML3Q73ZY4j6Hw4lxMJ/
poMhx3q4B4ThPAE016vvX+nAJQkAthPZDUe3lRGsWkRTxSLtjqlBNLmVTiXOsRBG
OWSMaX1E64+WH7/NQ159TsnO1NUYLvpFP/D9Zz0CHXXeLbH4SDD9NXhfXgufJi1i
3ahXeLD1RIlmX4jzNRmrm9av4BV6mwmQG8ddIm6RBkH5IoQeQ8K2hzXVYMmw/4A1
9L+p5ZN+KzampO+fXmm+eeX4nodOko4XyO8r7yQGkVtx7nxuk6zMmWE99Qf2q2wz
pFPI9rkaDDPEj2DhQxt1b/0ePiE3MPQMMKeGIeihMWphOrqe4IlH+NVYzn7UZCUk
GXjhnW5zGoLVupXGNaFFvo1re2gqKPRJdNSIozskDgIomCnKMTxWL8gxjesJn4fb
y2YsJS1ivdi2zWp1OEsDuMsFAjseyHVKsKfH9hscsZIbskoqYSrHTmcK5Z2WlMXZ
rDGXBNMFDCHvox1mgg/tD2w+RlqkWzXwhOg+Q0u8TcAA5uWXuEdXznKsK5g+0OsH
u7HBhWKrDhZtNjtrv2Jo7mH8+YHGq30c8n+r0cJeUgTboxil3HwYf7TEdu4YvEcN
bQl1SPMwT2Z+X4HxbXtanzR5mMuMA3YQPqxulT3l/qnpWhuWUwtOyuiP8tQMwJAg
R+dqH+xORQBHHii2p1pVcA1GkI+2ni1xWdAZX+/czDUzOewGBw89sXOr67rlpYYx
eLE2wV90NbqRvA9kkP+I5LqXAC6YkSbW51hRVL0cF2O4mdTzEYHMXc3szVWLYgtU
ZuZUfa/DHs6Tezd39D5vkU7r0NZLOIiYYcm5jt+4FCg5TWMKOvmmkYcum/cI2i6Y
WOm5Jj5JcFQ+pCEC0kyvVXhABHT8oHNEtDH61h1NUg85CKSvZKqRCtIO0cy2mbAp
FGkiX3WMtuAGKSmuti/k2crbPF7DdG6pVADSAl/YQEHcpTuPDgiBRl4PLtbaQQtk
92Y8Rv+EovTz4uOt5BG/u8l7QWs0ajVg2BlozB09pOAPpO8yNcNB4tL2om8YPoYd
GUgP+jFeseV5hPWq9zY8xLCNMF9KAhTros1UaM7a6OA7qw8e8Iql1g7bgirIB4i+
JCvwKPxLM18lqgYgnX31KJeopiaIXAJv8uu3AhmXeII+gLlPPDPYYDyFHCekWfCW
O9VBd4h6m4yEwAqav8w3p0DWVWwZWh0ogTnTQo6Xz7tSmsxZf5GmJNn+kJ4bXUIL
yDa2DnaISN5j6Ow0hF2Y6CAb6BNCojPoV6kSNw+cevC1iW99UwFqu49mau8cmWgC
eoShJfvDgnCwdtNl3MGslpa8UAig1Kvg0EAYGQXohEEvwhtLh8JLMf1EStRpt51v
nX8XWGCF7MoPDwXvoDMpbBq/vIZL0541zCFV2iGpvCwMzItIChF0yK2MKOEseO0A
ilRC6KHDgNgdSLyhd8QUZmArwkaWWogqChG4QCoTzvWNbuCydTmp89wKfucSdq9n
KZZJmvMqkssLlEmNLwHhoi3ibA0ui3QkLUTLeNqIaPKttMUidyvw5YBZwm5PDvRy
Mbu+ip0o6zN4m2O1w+IXLOR4gdr5DDwaC/UzVM35r4stVbbYn1S3iAzMBwv/l+LE
TTMf/Rt2u9S0ivMvgIRVxyArtztS2jU9W0nwCxt8EzyQ8H/lt1eff+advzcWluz+
sQHvMqtGx4qAnN6ArhroFgdjZaYV1U6VsB1XpBP1Gyw8FpTTIdqswd87da1A3Zds
l0cOvKo9MlWnmcQYL9Q/ek/f55Cq4OV2sTUGnvSc2L33Zl14fhMWLBUil1fb55rl
wIIC24lV2rKTsrzDJoCbxEnV9dnK58+N8pEA0Df4o0pYeyhh39vBHbXqcNfSmVbY
ojh8tWiI8tYVuncW4HULzXH5e2KjhMNA/0rQNzlIY+5bbZLWSnXuuVjMmWVaIj/H
wuMUuQTTxkyW2beWyFe0NoJPT6gK4hRUC4sRBjetmf1gX/ZnEPXintbiW/ITjpyA
qVcVLzSUECwNXvU+V3GhlrrOjaI6Sv6+g3PRRSeBjm0hwwh7C4ZTup3ryq4Az7py
vr+QD1ItzCfAKGbQ1CQW/Aut7H9w1of4UXWVoIgkORloemlZCIE79i3PaTm+BXvb
n13tnmOeTn/+8tW5bS2xo+lRD+DK5w2O4ccHuHKVJAZmTP0mAN/0xoug/iNVMauj
OH9gbH6mgVllZXgtGx2HL4ocIk94dGIo4u+AhsLRbqwtJSeZJ/i2bXOkSlXFP6tL
fATNUWcng+m5oaIBrJcVZ87GpTRcIo0M+5u/T/0c59v7uJf5ED4lKksrHCMb3ktV
iwEE4TLTYqo5WVvSv4+lH/tD7LvLx+PQz92Jv2+CLJiL/6Tt/9aEvLRnm1Uiq2Fa
YU7WWqra6jgXO9KQ3xYHNLXd2ywxSJVK6eLJI8Mb9ElE5UFrMN5xRPi7rwK7qr/m
PzKWp2+R/nsbJ11OAUtT3NANoy5VZrp+VJCA7d1N2N2Rw8YCHpf4pUmaNotzLksa
bxlGgJLQVtfYZ3p/IsvjvTr+e9+szSHodyOsjb/6CM6VQZDvD2QaI9JmQtiYHOLK
jJGVJRDXLsubrPEzRVTP5ra0Fnsl8somxMB5S3Mr7i+mQogdPpqv3cAbd2rsHhXq
opaachLnEPIcHekwCWNppUlLt2SlzN8c6eAJtmsrHKrFCIORoOaMeG5hLghlQKiz
hesHQbFJT322u6d4NAgLlRHyI8AvX1DsCat6nEpZoFnQpuSl7d7LIlEfZgqcItVS
fSmYSiusPVXBPT1E9X7J6tZFxnX+ndCKudqcy05ZMGpG+hGLZOwksbFPP4v1Rrtu
LxFeBhdZv3IORjlzyR+9NLDa6prDYUFnUJ3NfNANuwiTEG4AYloYeFc00GSQDCji
sMZjfJBCCCP+giEpnQHV1U8jRveC+xGOVmv7t13OGeSUbsTqZG21lv1DKNg3opub
pRb6YQb1ffz1zoxx+Ku+proiFz/3DcG5+PwLinbxA/JPVHvR1IX9Fmns1PGTh1Zh
5chCki0e1sO4UuwAIRyDBFcTEGRHqVY7WBpZKfmdagdoSZgU2lPfL0UOymb8uTQW
U4MkvSoxqJj9CtVV2qTRhWcq8ma9F3dAo9Ful0ByCR+2ylNyKzCrSa6fjR23owTS
a4GtNVuWbfAl9e9/xN8tOK2P1D8izs12CvlQnFZTq6vuyjTW4fgjdAoiTtQHRxYD
Y8Ep/5AwC644E0u/mKIZHPedZMld1n1NFJuyWpIA7OFYGtOC1k+lF4+gjObhvWLT
/3ZfooAGCpsbP3i2nWRvff6K9ilZGheMIJd6HCTaIosucNJyZtL02PS4rHZA+mEU
3mkkeTtw8k+TFqsxZiKzy/6WAtRdBCUm3kAXFVEeKRYi0Qam2BPAdyETn/v3J/Qr
ogF+rTYGWsrUgsB7osbLZdTqqDlO7YJsPbFEUFM6I7CjtEiaLUw6ozjpLzIwvIUL
hC1jK6duVz1iYlAynb59yikJFRjIR/zWR3UcqziwKKF6PjIUmEOzwHEUM89UoQ25
w5HbxBMHLTJCw9GLfdnQRNmSFh8MBhwn7p3it2u8mwylptdPVNBHwmokxGOZ2RUk
TsfUf0OwG9pMfk0xLbexvEHYRJ+aHYn3ANIbEcw6VcjOe+PeGBdvHyEU8y7ec9HX
iP7f532zC9I0iSyckbrqUp28R59fuYuUjH3ZBG3SxM7R9zxMD+KrUb7OHXAyzS3P
d6EuujDTSwo1GbFJefW8dzhgpK69qQBVhQqKn7+MUVSQNfDTLK3I3OWNqt7oCXn0
lUwu23C+wJPX1TgeyuhcyYmXjvtTz/nBPeYo6ImZPBH3WrUXjGLgfLvTQTmIlBup
pOvif9bXEjyxEKpuOrezDZBnJtGvSNcROv/+bBrcoh+AekF1OogpQ1/z43yibY+U
zasWMsVy+tOHhsSaPHgieR1YrfzvMIPlmzORKp+NMHElAGg1w0Wg0iZzf4/A8d+C
XpdoeAr1vqTBEf+4KCdA153tzGvzxzL2bwUVqTypCnWj+crg/ICal+XBkFXYdurZ
vZb1l7jycHNZlJoBxYOqP0UWqYUGyIPERo6HjEF3G6NcBNyaKn46sJuLhiClK+uV
u07++3xHuWcbyVarSJm0iBp01IMK+KVm/+MxkUSpbUwNOM90Pzh7pgtiKlHZF+5T
3N5uYvUXXVlOVL7LET4CpBLCr9p57D5gEGxxPIDZgyA5y4j0H343uiFoEhfP1jhr
sVAkG7S+6P0Ts9n+XPu4oTKdXtFXULrrEazo8FXoYsLXpsFWfYvkw1JLoC0AXIwD
QLkFP5ES06EbOI44+vWwYK9HL+NbIpRagMccYwUqrZHTTijhzjjv2PzR7gWWNWNp
g6XlkNemc+aU+lJuAy7XLqK9L4d4UIIQ92e5jQ4PpU3pY+RSQA8JEuaBmv8nMGEU
siZAJtgVYFoMOlOby4TWlSzLpW0OR+UFTsoNK1mSnRXWf2HfiF2TPYS2UHZqFM3D
4AB0076hDtcDYZ3vZOpKPtRbiPYgoh4tE3TsF7ZoPtTjUrwIeENBRFTYJTTNXAnD
5H1ugEoP0GlCC0LcA3fMGgSwOjrYmHsHv29A+k4bswGWBw1rg/M6gqDPAzMkWgLB
XrLANh4TWMGz4ENQ4k9nRi/3wE3f7zBSn4P6ROjxiQAzn0rjgGHilW1EdaBd/sM+
CP6DrSydk2sMQLk3Z5owSvz4fydJeda7T7nWIgPWGujyjq5fUEcroD7ARoNy3Myh
5E0ptQZwT/3/70Lw3oglJW5fqFT8l+2FOhiZKsT1RAwxOvZwIDUMXJBfz/xIlXKc
n9p71DvG7kzgDU3UXwN/Cl9HLzSbQBrpvQGSb8hqsLtDSm2fEXawask1HKg1bAs9
OA0Ok1Ddo/l2wkOOITmG3c7uLOXL4SOmgKY+KdIKp+ysMS6lRrESVIBJPqIAHQzQ
Is3bQ63N7UEDEThCFlK6TPhpPUjQ86kIQqdy7r/aHLM3DvKJYmuMPuJGlge5ix0a
r28ewoSxkNMzxWbnSqzKTb/DxBWLIbzkQEi/NqypeyTTsQ/hVX+qj/iQzebeG7h6
TnAJ8vKL5XIL4Gb7A+dELnHVwV6fGniapmOG9WfgyRqS+mXPqurrDjxrgFAATOgS
u1PAHq+CsZHpuw8vNsUJAaRnsnRju6xQD406hW8RN2wKIcGFPnjdmFCUu13gqawR
mHoAJc0kZ/N87n9BfGSkMQyauDglQdfJrpsKgs2+GsxqSwdqC8lcI2Mlq1Z5kF99
HvihW0db/zsW4CNEWd0RsHRJvqYRjT7iacW0btarQzkyGBzLUlSU13qal9+WDLFt
0PjeMYWcEj67iRIBc1+9CQGrA9tAsrCNQR2aLhdsMiUiqyiNT4hkDAZb8bH63wPE
Wx9bK8XSKxMFs1LtqhdRIt1+10lC3zPL9vHuYK4byE6H9xVwlv0SwUkjhpvadQtQ
imVcHBIPOyWmJ1qfezjXI2m5FYYbZ4/B6GGLysq5HvxkqOdG2r93t10/Ak/hMPOj
8ilTHqp7fsTYZCUnIdX00REZKS/+LIQyhKG9z8YPfSBNobfESXZu6GimRXwbnB+z
kxfW7PojqQvvrb3IHSrXRZyQUFil3DueF+58De2RA+O9hOPr/nNWWjPG7ZeHN0Bk
0uqGnLTa5z9tGw7IK8dWUcYIMJzH1VE1JqJI9EtxH4IYnkcC4EkdQfIjSImjm2Up
bU3P582uRyQo62R2ofjjrKwYup4PFvtb3Bcr/Mx+IJH+ogeK/yHwMWPE/t4jNqvX
TvrlFE50gAdAmU25nSx+Q2wNXUzZMIPJy5qCW80eC6p7ulXbx3guBQqsI/94bA2B
psjqlCiR5S33Yx6gdEKLZsUIa7vzCh+uxlQxuIA66c6wdrgP4at8kpAhGrYWj0mf
GOHw7KdGQclViZNvQZVWykVfRkCYsdJEQu7QDJTi6oUXqNQLhHMzqsvFrk69d2EK
k+Bn/ykYZLspg9svqWrqsojrVr5ly3oXvgX800SFMDOyRAMNo3OLAts30vb/wg/3
J7pq+3xjD3+GJjXqc29tj1avHe2CzW5e6U5bAkCWY8DQPxuKW/qKXWvziV5kUts1
aiTCj1cM9+RT9R+m+y5UtyjlNlgh1hhAN4m9429BtMdh5LxQIVigwz2cS/UgXIAH
jnJVHVwVCXjzFiCGpXoIs1BUHEr+qBso5gHnhoslKDlV+oOcY/wsc1G8eI/F0W16
BJzXXis6h0tE4n1MiQDUBlNX19jOnE12NDRo5ZHDcCQ6Jf0rHgqFWdWLagUg6S65
ZOUugF6T2k6Qvi0suXJ3l/Xx/26KL0DS2P6J7sc/iFmrVZd2bHy50uQVmHwiYOtq
Nmkac9TqNyzvPKbxGpFUDqtCG5kwL8FoOPxfqvjFW74TiCtsdu6IdUcPNuVJ6cF+
59qz+41pQnUZjtAPbxBseCSCwpm8ToVDUjsvhP8m6ZJKnjnc+9JUWJR+AlXoDBKp
pbSmFozK1uK80N6r8ZiFgTZdX2DRpTnMqAilN1Er9kossm7N9yRQvIWd/zoK6Dzm
zkobF49gYeylv7OF7UrqQbWi02ow0dQZAEpCoHKd+yD+AkvGMMO6R9KvJJDWZOMY
h/bvdox4A68f+o0Y3hG0hCWftDg0UgqwRPyvaFehtEu+LXSAP0FScN1TvAIQKOKY
Rcnv9W6N4J0V+/rNpZgr7g2KEAsNtmfutO9FtEUt+EQ7+xzj3CnzuvLSJFtlViGG
ejTKm0jP+pM3fKgj78ZAcSprnfzErweqflzlcWJN+w8KmeH3K8zwBiDnTVDZ8nVa
NY5Sxf3Ah9UpwnVZ6Dg/9Y25oj8XS7YADn2tqd25aAxkG1aMOMfU4t+6P47VEeoV
dKX3MMUdExCaKXhgHBGe35yKiEmSKO4Ur7KTkpteJRTfpF5XUO1bLV57g7ZBO2tm
Aa/vzrj6dmQPFzzVz2qAvfyg7cUVeFLfgLlGOtSmRw+QH+wWqUNJzT/4hmyeKEY3
Ee0JoNF8jXbZuxd3pgQzWRPR0LaNGMWKTF3JdToJH8AXCwFBdtn+cYvcub48dlQg
4Kc4O7pWpChD1McRQO2QDcSYKgOvD+Fi+JaOhviMeEzzGqLMnsYo8Xtt/ahHbasE
QcIluD5QbXXXlKtEanKTbB+pCZ0c7g+2FCUurGefWX8yNT7WZL48xQfaqO3N4Ie+
rngxoWRyK/RFCrjtHsb4MrTJsHVCfmKDZdHKoJtoodrMAdP2PSqtbN1xETYpFQB4
pw8ANDZiWGz26bU9IPqg+LZmM9CGRhXxHl7Wun23uxOidfbG2zaU/KaD0nWOa8Bv
uVsumcZIjn5TDwrxzxxC8fLIvr6dMdBbEkT9yjVcA0gLvZWvIT3fA04BAi0z++KH
rJlD4i8iDOJUYulcufde4n1Uucf3mgTwyFKWQC1wUjsigXJZUkbw6mLgweeTE/xM
cc+nrG990faPeUUEExzlHBHCusv+ztFE/rUThctr/E2LrcjQX02VkEgXo2/E4lKh
ucjNY1x4yAfYbXq4FxGK2iHlDR39tgbJ1C0RBQIuhwirWabmVUZxvjKIB8vEu/ut
8lI0VBeO5EBNlC842dH3QkuGkNsuS1okfF8F21tUF71sXbqHM2KD5As7D9VvGBPP
EFFw2wAgFb+CiLV6juExAingGe1l5h6GU/dYC1NIAZbCASZSEpWEhSyPK9zhyJ10
valYt8VN+W/hpEimgUY1WNcBr0FKuroVps1WuwbL++Y4Q3qbAvp1LS8VmQbwzR1T
WbWcRPRg3ZJ8IVxbjXXMiOz1NeqQYHJmVEL95WcZ2Jv31rj3dH9YvFI1qYFKzo9O
RotnTw3dEMCXf7dfVnpVQ+Phpg3U7rqTIaPaRZ70vNQAmOoYnkLMm9m053QEZzjq
YGwnwggUo5kozLizLLvIqGuUUI+z4X++3TJVD7MsR9kEsjkVLVpuHQVwDewzX0I6
AuoX3t3m37MH9E+BIWjZdUSJNeDEfGgJbvGSjTlsuO6BgO7BmFC3GrArIHa0o440
UCacaUEJ7Mk3Dx1n2lKUsv4TM3ZZANW0XkBUKaOQzXKAt80xd6HielLvUYuIM0nM
44VOu0mIaMCCHk7i+Zvd76arknxKMgh3I4/WjXfNRcW+iR0kBDrjBcysdD5bShfI
MFu7cvz7wfISP0C5V/7W9kNquEW+Oj17IO7owrNY6WP+fGWPWWf80ozGLCVySqu2
9Kmyx//nZ6GgcTgReFIIL1LgN6GrIKAP/jNlIq6BcRx1Uc+0vj38wUN42fRs8rTp
5tXk6USi+cj1eOG4/qvherHVN7n87L24Y/0A5HpB8AhNzSQu4R2+UevtrTApHYjZ
u1nnTGozPPd60vX6vFsOwZzVzSy6PR28bS8D4N9REjFqYhGKNO65wYaTobeCHmSH
xZkoy0qfxV2zARpZgf3ixuB+yzzJ93ITVaTcGF7iTxXULq665QQWSls8t8jndQdD
K+JmlofeUnS6jr6eE09hfD9vFrnN38h8MhAD2yXXL7G6pKi3mP51PklnWTRrT8xc
MtnUxB5LHE1rTpYPnqAqMlKS4Uk8KdnbpAdJKfqi8djCLitNcobpJYusE2/1beyK
/Y8Ayg6d9DMZmQf9/9fYtX1ogSxkTzkHFVc7V6BQA6XahC//mPYCwqVcFOENpmLj
FxbAesL8UXik5iesHk6ats2ZCSf/j2ifhHqGSJUDE4s+5hFzNzlGjZr23JoEEpXd
PzYcTb2HNII7aEn2gZRW+YlUKt1AK138N7B5Y8K74rpF13EogP553eV6LlxkDid2
XrgPefuoex+thuNSHbYoHF4Lji0HgbaD0kJiulJ4by/xJon0SVuIP3jg1v57K+pA
tlFHe4IGEKHmQeBKDAIENdvYDu/kNQYSKGa38HFRBFQhvmV3kR6ehKTxmaRDPIGF
2X8KxMWwqOSiL5GYZOchDsEx0ddTAHXDEVEOpFKT+3vvMd2JTpupx0+pTNeQfeGu
nI5VIWG2J8qyemVne4MgoBADSp3CcpOQX1JGksbz3sREwQa020wNwklvScoTEl80
D2WqEO9/auZlCBjaPLXjAnjUyvald8NUFrVKVK1DlsgcNuF28BTqTNFBEQ42hLe+
PP8qXm964efcfbn94kaA+I8gihjN6LooLvauqPtOjhtR56nmXMVMKhYfmmthCiIy
nrzKIRzjqguc1Solouvas0i1/L3RXIdXPJyk6uVUX9YP9hmm21OJpLINQelmx+WC
gwKizRD2G9dH9eYHbePXwxa051EySfNHxSANgELAHdzAIChCQwffRKaU35d15x9I
kJfx1DHUJTavUjBUbUuwyWzZ8n3118QvF2zWsunMUCMBlDgPl4HPALve99HleIPH
iFLa5+OlRiBcc2V/zvXRyaF0JdhtXeG4RRYh0rtB5OJvyfclKFSuprV29eEe/1Pg
4ug24g8LtqZybkhbDjBX++7c0ZCN+O87saEXUh04h44I44SRmvp37LH1T3HRaZur
fq2Pp6rthrMTXkt7zocRrxkiH/cULkImXygMVFrjnpQQpeKcvXgFik2Tt8ZcRzH5
o3uCQOW0CPek/7qqnIFw1pYxPKO62Hgg/tyqSZoSGEUhn9udYxvQEG2U3jCoafpV
eYZ+yOxCGo11ybKO/PXL6jfbukRvdCWzWRTI4D0tf1p2wnWQmbceOvOX8qu3qwQm
4c20KcTRs0ZnuCBursTR3S3aP8ZbSbZM/oAOR5Z3J5xhAymSbvaTcXe9FLa2Hnwh
KAeBRsgJxnePErwbAZ8Zxlb27sVx50wmVbNC9ePs5ZIFP70SeIqZ8ji55aPVn3kG
4KP7Ju47+fZw4/9bEMUUV8J7MB9FORumOLorN8V3TWXmkqV9P8zOAd94KiTETy4V
9KiEZIGtb7Vr/Q22vfNjSqujMe701OVc5WGGp9e09h9SLlLJVDNN3NXPWw48AdhY
7tpC9rhna+XC4vG/8nxUdOr2tEinZOLos7BO0tPV7gKcw1U8IoEK3JnI8sRtyAuN
7G08xT/kUlH6Xh6+Tn5xcjhyTPnUwZ9gLplshDIIRwOnD4zbihplHgY0KeFfu3d7
PneZkMEapkMg1dJX5nCQya/hZUW+uNUADlhLUAicY97deDJJEoyvmKDD3IEDkrg8
gmi4VhjthNKf8MleNSgFQlUf2RwAaLZmZnPxeuJqVk8AsAt3qf4Q+H3+YXrDvfAS
gxJgSqiQl0YcVjMGDQgYac8NMREupNMwLjOLEzphVsP4XQ7WWMLitlMcjJ02rfLv
NAVqwvWqv1Nft79z8f/q0CtRtKJ6iM/X0EEClZojFQQhjF20VCV0p71wSjPZvAAL
bC1ZRuoJZw4KlJsP56N1aIujNlMKR6U6FOJwORoaQv7crMON9QdF+5TOZSMowuAJ
LugGZJgqf+ufxGNHw5KBcvO5t6UPaJFwPycpDxQzhSb6CeAn76u3ZXDab6844Ksd
BTj+Q/G7mOeU3uYR7bI9AgT83OWw+Xw7jPzGnnOYHkToCBLlCAhq4UyZzUUuAnDe
n1z1scAeclw846ivFuavSbmoJLfpvTMXCivzjMLKlL0y5TTkfNYod/iFXIeYxYwb
AQ+mLht+w0QGQQtXV2RGrQjnL7W+O+rcQr3vwRIZo6kw52VK0LoD5IIDyy7+7p+B
WJ1hOWuGbbornshQfR1QIgqDk6cK0xaM95VodNf/jjhy5Vj0p9TrRq+xf318Wduw
DRBtXHBa+R0h5Z+dSuC5SheCUyyPcPeltKUKVcG8/TigcHeCdXck/HCOgG1I4QqZ
wfsMqty0IPw0nW0jwdJrTu9uUmjzdf9bhj6KP79etU063DTrtxfToZd67ZJIjN1n
GOEBRyJpdyp2CEWGZsmCgKRUgnryE9aDKMrXTt7Bb+2oCtaN4zqBuThMozrks38U
RBTXwPW28Vas6XsSg+WO+jr+SKnI3TIgIGFhUpcBT7/hzaTRcv1c/wYtbENS3GjS
odvkP36VqXXHonXV/9/9CEUwFYUiHjYcdX6bRomQbmNBV9yFiWnOCSBVh+zDqSx2
ZzsrSIWuvVTvshmt9Nmr49zREFI6mbEq2nRNKBS2Ssca9sOOe8n3uSfZGlelPt8a
cv7fhukEOrHL0DrQGr80Uf/DNztdDovuK/tq9Uo7TyErMTHQ3gPruDsy0/kOwDkJ
4zWRnOtqFuGUktpbYXIg9coXSSo9c0WpscfwpLNi7blseYnT1PcpJzl3cIgCkmJ+
XdQxNdjs/AI90j45ca/TKGyYbfxN6ptpYxRtS9ELNUUIM2bUrqClTsNMQ/2gNT5j
dV6In8CMwyic2fXsCnk2VIRj9gQ1J4q2j930hT4WDwop2jZdx/289lnPrKQhlfAe
QNj8qWkMrNfF7EkI2zGsuho7yzxFddxn+3I5nu1P2PTxD29AoD+U+4V/HYKynxHd
t9OcetkruvD+oyQyFlZvfA7zfolszkdkxxcURFa2ANhnOovG7dTKhjqViPepXGtt
rF/8AJvnxuZkiNvyyIzsLNAbePaUItGi2iYZgJaGKEB13VF37a7O04alZaODXtHM
xF0EQgWz9PhNr9uox2i7+u6/wF+Ts7V8umFPFn6yMJDA5L4rsnRyhel8dxUR4SbW
bLFjHrm8ftvMQNRUcmvSoff64JyKCKucZuNfKcsbBFSXDrazX3+SmedFzoOdgQmL
N7gCl3MOPtgir1RRqpX5vZpeIKnbxs6jvResegnAly3yJRUgv2UJe0RhFA3r4ctH
hQ3dXzh/ZzNq8aOsMVqafz+keQaS2m7VU3f7ah32gn37We3THnhh+Grz78wctoiH
WGizbRbrmyOpYCN5r6h0E56AOGKUdE+L1gyQpC+PKtFqWRYFdeAra6kirv1X4kYT
1z4oJV6OfEN7CeFpeWfnoJwWC5Rs+HD71r3g8oTr6RDGk5pXuz1sARXQBKdcPfbk
hIy3UuVwrmGaEzkUjdHO4C/jmKHjvw8EIB2wSSj1WvMWd7QZV0BQWTnQ0/K1PDNu
ZZcgPP3WS6ApWD8dr4n9+MMwT3/oui1JsaiNmC9oXPjm/Ra3PQ8n9rZrizki4Ua/
lxsDtdVSreKx1H7EyBBe6NWG6+GsrQO8Y+mVFk1f2LM/jcRPiCIuVGRwxN0Qt2TS
ti386aBvGiscnDTL77M8BuzonUHapq9I50W9yr5+o302P6EvmqBlt7WgfeM/VDUy
SLa3GonBAhBK4DV/p0ARSg3IoOizSdUiVq92D+t+RfcRF88ek7Fm5y+syNDkDQ36
3JRvkaTgWpww4jNfFpm+GSYWL6AAepGb1XbKP9OPTVxJQfD1Rfym+/E6TzcpEKzo
xgnl1QL2KInb9NHBsTDLnXz20XrgkkUTTxEKESm3JGEfA/xkACC8r3wbFozISBNS
adtAlD+dSb7FClCCIMOud/tpIzjI/Tgdga0ax1zPYNjfTRt0vVhkBSkuFqhA5p23
kf7HwuujckE/xadmYR5vxk5Vw99el53XY96ZwbSczBy3d4z95/s7+vcIaHpj/8OL
2HjfTWt4FvNNb0atWK/8p8Y63IQ++1Bh0GWkLW31NLCESCiXni1UM8461pvk1gmX
CtvV27n1a/wtQPckf/lCd48GhZO6ge4W3Rj6UvdcQ8KXt3nVcSDl/HI4aibY42zn
49HI4C97ihowFkNOzerCzba1XqpIezM31ineStHMUZJNpVqPBeciSRHD+FcTRIxy
knwVc3g/utSL1ZWCL/2dVmIvHDcs9YK0BxXZKY4/N7+8iPu3S9QuULH2ABH0iH8G
7iA4U2fe0h5VCmAjybZuiii3Bhr+j+b6F3r2KlU+kTdklIFcUfCtW8wca54skpdj
Z6MUMDyJlEq5oeH2+9lfiUNXny6bMIdB45Q+xBhf2Iaj3KdTZzT4yZYxo46AlhAK
+p5RVcQlXs6fPRcL4J/mYaV5ANt4+qqvOszmf6dnixSmuZmsxINmVM+p/9uqJ7fW
ZKIGvHrRiw/SlhozZXlleC5gNFftrDz2kbCg/BldUpIKxQTBVdZ72EvP+09XlaTI
2wszyc++LOm3uJJ136D3IA9uvVeESuz3M1B90o7+WenRaouHKSyYU3HnUH+7X2IJ
VQuRk7GyW8sxcU54ZUUHhW2EyTq4GIVVqTCP/mZ0ap7uXlwCgIErfVITgADEOPqy
DNd2YbzcupP4B1rBuIohME71zoRpXunbxmuU422vRhNb+tGBMoK+LhNMOv9kMqQ2
V4PknT3zY/b9gFSoFjhkW81cnWtyEHlvc+6jFOFveJnKXTQmpBSecdZNRmrxscZn
uA7cfaolgBE29u04QLjm2ebA/I3JDiA6p5577aYdUvwEJp3DTC7p/QcHj0drXFRR
jupwRSHoojlnSjE5UJ5+gsHaY2jSr7+qjrM57LU92d3pJ4jLktWD9D8098vLbFDI
2Ctx3FPXsQBmEO/RQ/m/DmPsQqSdlGM7A4eTV2LXvC0qWnywzJ4u5QbWOx/Wlra4
d5mj9eK5qfjOcXWmuwE+by8fWBZGdVE0vu1Ic4u9DHRqNXiDyPtgmlCaheGCRhy8
M51F2twlOTOwpl8OybH5WJWXuf2ezrfIx5nBG6BThZJ+HeXClISFthNWfLjWV5Ry
64EMniK7ZpydHB6eefq0sBuTNwywdV31pn5oHsgDoS2PU+Mr5pj0DVRIVkq4+roT
5tD9lS6g6Cr18HUbG0pEZ7LJ7gkerNuvz5PJZOkiNyUHzNu6Cy9ABkaWCJT/wSeb
wIWSKo4z/UhDzUamUBJboG3m0QOG18JkW+lDCKj30Z21py5MdbLQjZfEZjPTV94N
JTNW23shVnDdPtV48mBoowOiiP4DNi1p+x9eEnFnJGVkA/om0ke6ytpQKAsr81aE
EVDFum29yyq8kezXFRbfUymheVEjnR0VzZTV6uDBYfoTS2Y03WuooBXDhEWll1zh
HI52Xyth5CKEEuUXCMaNqeVijWkE/CbJrXFhpmp7PJX697aPs2NBBnb9IhOyIGHN
d3l7wKPtu1Mg8Mnw2+RzdtrYP2TtuSehKSR0tMI2aVlzbwzFXFe8XzFKCbgfH2uW
YLKbrR36hVmZzaJRPaQt6aAFny75j0ObJVP3u031xqBf3ktwwf4mW9A4jMykcQM4
es7wse7mM6e7CHIveu7rvgFTJcvCjOtpufkqcU8sQ4H8eEceFeIfURH81ys+C3X/
eArS3VfJHfxJdENHD46c6VO1/bggBv7cEDTP7QcefqBiHCsgFQqYZZd03/HXrGIu
RrBoRMm1NJnOZFrpzBHtFEuOgVTanSJ8xQfZFMRh6+URNBomeTfPiLCLOjy7Z7nZ
e+Nx7WD0pA/ib2iM3ZocKgwlSxUVOAH4EtN7PSYz7uilWUIzUgz6uOeHIHGssSZU
AWCVsXW7TYRLWZ108oHPojxEntHwaZasjkBucVk2RtAFAIvxav5hRwzJW1vB1J8Y
iH1zL1mSqeZfeuuDCPYFfGLPLDOOyalE55ru1nMwHpHEzk5yVHo5udlZ49q+3OMs
GnceGhDHkpWlJlZFjxdj3jvV/X44E+6M2CuY01gPEdWt08Pyk7gSPqhuUAnnb78J
N2SjaQmrDm0qfv56Zo4j0xjK/jvlroQdEeZbNXCYFAm99caNyDkp9Bco7ou4W2oa
i2oEf4UK7INMeznypO/uAQnWcFENiEYCli0Eb+TS0ZkR+w4XCpKr7K4dbaU6pQ64
uFOEqACUvPcNeSW52MTnw3jzI0y/xn1t+cVKsTxkK+A7jIZ55cCoW9VYtsgo6kmS
w5a4AVA4G4hU0qtq5xVdiST78b2AVYUzJLHzcX3IZpLohNTdU4eq1uTB7JXM1xsx
AXVOLaUP90UCrSy/JjcnpvLYzkBBaTA6z72Sc2DjpwKtj8Yvzj9E6CgU8brGXcmg
YucYOrEXvBG3JUkdYzht8Wu+iIvUHMaKPEUo6H3IAu1i6wT+zpCPLwcwpmoF/ycg
vX0bYrkeKx4IS3ii4bUIW88sT+RPkAzcb+2ePEfx2uTm/AhDwjXq0nQBX9KYpwP1
fvyRZW3uvpnwyLfMGZzjm4GU7rKSXQJQhXDCGOENQbIYiK2EgbOKEnyzCNhXi5Qz
3P6X/5s2heU3LnTelZfc4mPGwGeKq0GTwLnBZPPNpiTsEH/jGszbtLMxAUk0GvHq
3q0rTuZZs0soc8TDTkwVp8g9ZSEGsrgKfh3HPgvQgPSmFNM3JqeK+ZhDJfj1jYsH
3DHzdqSrUntYb8kz56tF6ZLIs89918UEaKnIu80Gag7FpBIVCLwLgv/e/GL2xjA1
6l+tuijbdHGoOhZ1BxuRtZPRu1rmd1IXEpaSSp06YSdfDilDvNlpF2q8/BeOuWSF
zgsKoo07b6L4MY52vk5tfSUrW4wxXUSCbuiyVTx06Dbul1dsj9xA7yAZm+Am1u8e
O7QHTExRHo9rGmJf4E4DnWBHhKNgcfphk8JqlfyeoGdvpuHAUL+bnj9RJnFGOLPC
/MIhvBd6S76dL4smB4nWQZhrrNqpBXO4ofDIbkC1aKowSn0fdN+BG476pi5qgwX5
yB+5K3B3tYCEgqVFBH9BUUE0vT5OrKgiSl++IG9KwbQDULbPVC0Aqu4M+iYJ//7L
ndjgftD21kDIr5YT4qTrBJJK8vFydMDfxAEQcXRgPohXjzDoyNXv8LUwfv6Hk7L+
bFn8kaNU9rXca2BDH2ffNw9PyHM4m5XEtEYuRHm8/z2YDf7pjOi2CmJNsAJZrkF9
lVAxPtLIvlkTwS/5p4I2teFnC9UiKsK+kin4lb7FhoFi6YVTRocwqVagIynFZysM
5GTEIy0ZpRqed8eJHtyZ0lfYDpZrTEM+SJ1mtImC3+ZeSJ1ttueouJmpKUOxT459
CTJhFy9Be8YJvMwBZcfx+PF9Gza86GgPcvoWQbwvQoVEmf468GfMlYtUh2+FhOBS
ykUkxUafOXR7cFSnhJSpEbDiQ297OT76biwKAWaTfqE4pb/odTG6gy/wBrHp7wAC
MtK0cBcpeR95uCrY78LZRI5BZugMDIH+cJvhWoczHZVlfSmZJ4FKyHqLglKst20I
s+w6x2ZD8zKbSD5HSoWk/pYFE9isX/RfdSiV/EM9WFEsq9PDd9uwxWSl34ol5W4u
nGti5fgkXokWMFY3e6foOLe9ov/0DoUMF3AnnqYXkQjdHmCou0loo1XeKt5gIk4Y
nH8R3Xeid6pgUxvsPnjY5VuArtqLDufAxAnlubrbJTVKUfmXzrufYhW7iU3uu0DG
bJCGpXzlOi41TTfzM4DcN4uG/dGDi2Zn7YyE20Po16IGLjYgQmEc8Qon72Wq/8AI
EpABTLKHWMmQM+381NSZfJOv7pTTKKNrnL1ZXh1b+E77Y9UM+nz5p0J6oKaU0CVw
XFMo9WJ1HfU9LMvxHVS2nCxaugNZ/AyiK2ODp5WB/ZtBZ0Q2+M7QvI6HQuesTt6R
Dc9mtCMKn0LGlnVprc2hha1D3yVmMzzLDVPWe6ULYEEc9nojs0n1pu9/bzrJUraP
P9ouK09hqmi6tiE7tOsi7/bKAQ49LshgZkU3tdZzLySUDXU/dxnfuYUE9SKnhj91
7zWjqnQkKKt10YKIPTPfVyGVZkXvgxwwuuiPLsYAaPUhSa/d93aNCFJMdg+njYvw
3rMFRAILu2N2CzYmW9ttSGGMIspMJ+WLlG221IAsclAO/l24kH/I1/BIk43wSQmq
X+wsw0SzyXYt3Bcqd3AWA/4gx4orhbXjSaz8Lo4B8l1Ihv+G//yRNt2Wppg+jKEC
TyblXecG0wOkwdDDd90J6dA7JBFqlNacG50Mw6v4x2l+rWHUmmt8npJoQO07Zhrc
37q0GngNxfVz5z5FW9y58jCNm5QGHF2M0VDyLwrWIH1Fjbe8ahHdl6LNhU1Qf2Fv
bKnN8+u3WAclNxRa8aRgIBBz3cvfOQ4yHtPipJXCAYQpFrdCq04rVw5Vdzt6hNY1
sXCfEHjGLrx5z5/WETCZl8AArswWhgI6IdQ+Rr+MgWOTrufkrmX8v99NpPjeEjot
+5oWDB9+Ayz0RfEd4xse4DdgmsqqBGEyIG/eeaZyTn3aXwtitBCZylhsCRhQuXF+
uUEWdimTcyrbLyn9zaEcsIzlYCCOTkh0B5BkRfGA2TgrrKmvIRthRhYSmDCKcMjs
rtKhbQm0uBttxQwOwlmVSF6mGVzngccVXxbAaPXaFO4Yr6ULQ23nM7ztDpz23WdG
rdrKnYRhr9tHlpH8f+FH/XmHMdquDlxMg8o+rZpWHL/unYi4fIiQtMNsOQpwbYIB
pSwOETaztBhIzlPpux7+050HT/J6qULYStNu0pB/mdi2+j3vIc0PIgThhgAzdTjd
ySxmAYqgM+CZ6hFlX+IP9BVvjX6cppFBeZZb6ig9w+Ss55C6YIkXnoHybiPdEtf6
MS4wyZ1T5fscHJaPUUjS2NXkCA5ls/ZCuLkF48OSyosVB8ldOvabNzumnM1fQwmw
plr3GmKXneSS7XQANRYcNjwBZWpn50+z0UJGIvAmdbwhy+918kNwTCd1pwMCNmod
gV6iHY+quSHZ+Zrtyhz4rvlEyPtLR5TVPRbxfll8r9IMbCnSpQmfUeXeM3Ij5X9+
DGdvzhKkuyp43hNQUlGRTwG1Oq4scGNNX7z3eyuod2JqsuoPI6GjmAMG837iXdFy
S8rWfiqNO3UPyMvuuCUJQEYy2cFlFA1SmnjqwTE0kp4oSqdTBFWSkmZPY/GfF+MR
66GQSsdH2n/ZVYnVcuFAsfPXN7T7r3t0hvB2p3hhZDq0QOT9E2EIJ9iqvX/NYa1s
yG3X6kqhItABzwXmdejFj+t045GtvV3XcV/nP9SIiCp7TYAn3/myoHJAKdAbBHhf
u2k26Ni4uzuZGJ4h6io5ymUvODcNKGW4AIuWcib1uu2PsqAt5qpo+lntjVBGHBGo
C/Xt4qJyP8+bJj4UWzPhpOzcaz18dtFgGN4KY2zdparfgCZtafb3JnuOnmb1ZypN
Dpfkxh21ynStcd1Nut9vRPx8qTJ3bRESC67D/JIGC2DkyS/F8Ebhslb9m6Jd/B5I
WuIfRAMUTryO/6qGPHoCSnUQrvvlCCUEGnrbZhBCOp4KoNQnyXVPSBI9h0yNdHcx
RHMh+vdKomE0wfqaGkXvOGBzZ7JPe0QdHYV0qj63oeQ3eKE5Mz1BlVfbRPidc5Ud
sgpzQK0w85hMeDRklU6KJWzyj7bqUNLuEHEUHc6HRW1PLcOAOPLsRe/AkHvCW/4j
bzSbhGQdu8jPfU6XTaodcFde/4xfwlR22UwKb5JBHPrTVxvowePtmyS36YmaBvHJ
uVBQ+2mSzMVjxFPUJz0DENQv8O5o5zx08YXV6KRmgMGBKXJL7eQltPPpml+0g8zt
OGoQlfFxOy5OrVdKZDIPIm4+1JRhAzlBNza+RRxSKmyT4ZoSRLcvaEj+/6zNmYog
YmKluDkLvbrmYJ8LsRp4ZThR21QI5IdChsxt+ewf33p5pDSZitJovqsEbEojPmoo
Xy1woqPQr2/uvEzJb5PjGwVnKl3KQz75RLi/LOF+0tMKlPSjQeZe70kNVXetRfJt
8aVFh7MRD3O4eEJfdf3Z4+F6jHIwc6zBwiZ4+Rqby6KJLDWkZpp9KIzsBy02zDsL
G8mPveiqz2J6Hhysex6/2hwi8Bf6Thoq/q5xZKAeaB7ArFVnnnHcHIFVf43Oe1uW
CR0iVy2hqODeakotQ+EdlJQxBlB3a/U5GzVNPrcXdswX2zCPsPp3zTLTXLsaWcTq
GtIUKF2i/CKd+xY1jD7ZoF3SfPa2BOmHJLV3hW7fV5we3CYHq6EJxJCmb062DfON
Ovmy0tBNZfbXWKE/2wCaZHT84ufhLm+bdnzJRdVPtGOUaWNtQKMVx8XaZlqrP9+/
Oe5+SEZf+7fWX9De3y5BEta/gOhhcO4UstHZu33U/eQa5Kz9HIXnKwzVhV5V7GoL
+eKp7p6XSugVKjeLISsdSpOV/jZtRvtPZKXkSn274jS/coE5YQHliJf6rGhEopIX
LNUVJ6mbLhB8xC0gdW1KlBlfiRCtGVt896S5HD2FDv8RXeU2hktYIzweblGcU/NN
mIkCyTPim4Hb0pZEop1e9xBNyRRj3zyGbGnDu0to94/RUOEPSXf/xt/U57bhYSGS
cyT+mkgVD0YiIQAn08HIpxcNs/TircW3fWOm+CnnqUJg1UCc+iVrh2oGGbY+zcTM
tTud0GVKzS7RReXrq4Yr8Arz+ES5cR3mjue49scR3XGS4Bj3IGDmaz1xKzaziUOn
XGW0/dLWz2YSMIO3y/b21oDborDBaTcHKYHdxqsN+ZgKJLRyDHQsHM/9q2PCsaxz
V+8ea6wa7bGrfvLZVSIQGG96dX0WuDunDlrDV9xq+pzCA99aT3eWkvtAFsA8GpJ8
sYEcxLvSrXLsjVMREDHawcQi/muNKKaDO+iMWkUp1eW9MHuW3x9GHVsv1xbDp/xm
7mJDn0VODmt95cNUB1wV5/vIUezHchhn1AytT/npumpU/6n4APSutPOv5ETHN2BH
0s70MvtTjQiKQs3t564FXhxaLxb5F4I4ghEZ3/FBVzZF2iFo36a5h9KqKTcqIf/H
dp/F2rTJXIZ1euTwOE8i9toDmfoo/8Whj2pxeK1nzlwB7yPOGglM4vEGEuwTzKwb
/G90pKfM3yeijUzmCH/EJjPtV9ZEJ5l2HX0b3vrKWxDyoGduuLkYHDAu2UH+4BEE
LVkeA9c45lP85y635DP2lwK/itwD3gD0frxVvl0juL9UR6Q/94qAw/5ugWEIE+1r
nCGfkERfVEgJfkTbHAr7/YeWfgLqcFpTQsAcuBnYzxGluX6UEwEw24UBHBNTw6dq
6In0ShOoBmW6NK0/vIDYeVteo+2cGB1duJvenGsfph7UxSbwzpp2pVd6AST/3Y3h
fbRB2R16lTbfcV0OB6NqdVoIuh3Ikwv47+MIFDkxKaRH/FXmhoQ9zltRGB0oCiRL
V6s292enAPsJc95RBqCWRX1K+hXnc7eYPe9Ys/dUgPdXkNV5SF9xIhnJxuZteY5l
DlOqf+eC5fs8vaSlmXxg9EIRzpM66NqFc8Pqu/ye69Vixcvo2oiPH2lbE2vWSfbg
QtJAFHgvzWiUcbZEsyIi5kLpsTBdbCIII0GsXWr4auPFAazXsInk3hQWyTIaL0S3
ssB6cJn3KtMs27btgcCKMn3+vGVoxUmzfGQVKN4EkC0LBXh4AXeQC9Mc3disc2zG
BlFRvhzAMlHS81nAeyJlp6RKFjL96BkUlYRSz+bu/LZQc0pArfd4mwXcAadS+SBl
ZNpwLhJzuR/sSVf9AowfZvJiZBn1DtI4hzC/sdSMkBMXGvOYjntCyL3SKT7DD8Gj
Hj49L3YnD0W2KWfUChHw8fgLjmJXWGhrTgxyjSDJGXhWazgcSihjDkx2kTmnyFdp
WJeKpEVOw2GFyJxXGvHzmqO4eC+hFx9ziUxeir0OqprVmp/E3fWBESwZHQFbbFYP
dol6clc0Scy1f9UaJpkse/wLaFIdq8OJ3NZEoTcRSB5Z2n9cnHF4TVeTEfoS/kTz
GeUdkvarNiqoVY2uKylep9hciUJw2xzF3INheP91GKHeXnj4Vd8Zarq4ir6sGC8Y
0L1IEMoI25mna5o0yBte7ZlUp3bn9ksT/bGhGeSno414BXamR6/49d+8ZSlO/akG
kfvU8F5+r6jS92TqHSbWPTwoUTxEQXlryVJ611O0NysBn+lYZ4Ezrk3F4J9uhz40
Ez6wcJ2vZ0Et8iwDoXGD5WFUsnhWh5g51c0FyKqc/6CrFLJaJmTPQzs3p6cb4Qfj
4DgElkSxuCAkTtsMTbKLwJndEtrTm/TODNJXHTLsZJVxXQpGTpvEVMQ+ieYrFUGh
/2NKef1uOiG6W+fwwiDdMSDY9lWz5jWhjTcThTH+ede0jJ7lsJQMQ/UHISqCgdfC
v/mGihHIIESty33JBBLGRMXkoR9Qp6njlUz7f/dUGv9aRbh4O69IFBRXAF0b6kfU
0Yl1a+jTXmtmpaKxFv2el1Ju/rAFf9L2MgHUioY+AqEPSGjTKL56oxNDww5HEnJk
kxKc79u+t8RtHDVow9td5OCI7ICnR/fnjlwkP14TurXCSADQkUzYtdmxQ9uiSQac
n+VEtW9/DF5bbcK/WC9gI+UsdBfPHg03qxaoqstp4Vy3CntCQhq2TglLvSJ0mUHm
OxY2EzPOxdyfSin14GYGlXOT/bkJtwL9hOVLZ9BSyzEte27zZbRioZap13M8nKsO
ZrO8e3CoXOOHtUsdH5RQZvkzixwojOlqSicXoEYIIVVhHADCqNHSIqw4DUy59xt6
xqiK1ynS5bGz3Kg36hQiWcp6hYTfXoOFAoEEvZTWQ9XcTtIzAAiPk9mDUz1JX+nz
Gybhhvh39OhQPhL3JSKVOg8LlbZAqRkjXJsj4hw02nWA6EymXSLTyBksF3tYXnY3
1lc2LjuGewl45W5e9MSBvGR346GSwDy+ZsXDXoanqudU8UPYhyoIVh8kbAd0Uyz8
SnM50onTC7kKYHys6O4iVcoXCF0aQBbRKo6DX8TJPZs5xRZMIfqXjYUC48UER7qx
ovi86NNlmadnFkUab/rg9V++8rivKunx1Fsp0HdjS/rP71PKqn+noTY0UFLjr47m
9L42GHaA+HYD2jIIjJn5+hP6B3InBFHnVuxlrFFZrya+3laqr110MLmhH9ZlsXVL
jPWT++YRGJysPAphRXn8LEmXPIsRoo/STJyVbp4ATxzf5UTDq4eOt/xp3ieYu+HU
v9VaNtGiDjPNfGeDR26D9wN7ywjM0s5Xn4UVcTugW7gWhTvpd6gjSMZdb/b8bgMB
3wWDo7KekCeK0EN5oZStkZbK8QbMsac8E4r0//APyu8NUY/JU/wu8VZ46a63UPt7
kGuKvs6LXyne71IF7+r8lQIwYM1K5Mt/2FqgFtcap5qLYzzA09cye/S8VX7te70b
opiqv9F41492IVKOj4a+pWluDJ2qzsV8ItFC6ERKa6G+cKHG7HnW5WmLJJs9baxA
dj+5Bcr3bnlXLh77bgWLxlwsdpzFohkqhN9CYjRroih6+zWhFDH82TiPIYKzUJmS
LZr3tC6E6UY0yksWAvXOaJNlMpXoaO8KaqmaYp4uumg6bxGJCavnMfIIUI9dmGHj
t8JnNSuNaDCM7Wqv9K4INNDuU/GeeOCn5KE5gXHYkjLrqjWBKOMOBuw21NIfJNX6
Wgs0PNwoemgvuuYTOC2SDdSth8Yv2sQSQFcj5k0iXHXzMhqB5qLC5kV6Jm41LCYJ
0U0q1TS6zwNEG+LN33CkjkNXs7GSKZl0l+KdWUVwae9FxaycQMUTLzq5sx3vw2GD
xmq0YXpBPMXDDksAZDbIWgY8cMzEi9SZFPyQeqY0LNSQbRRXdxEa4jHTDTH8rUU+
wwNyLrhzwAFKnaivkYjDngRGRtHWY/Oip+a0hwl38UT87ztkILChNJM1Nj/m8BNe
0euV1qf92WTYqqZzZ1lRdIX93xp9p9eg+gzs+/B7m/55ljnJcvoBqNXrTQm1uk7d
XsVDqpZdI249bxuioQnhXitcRPc4P81tpUh4AqjhNVb1a91nywUwkMsYAugZWmzK
ZNnxM5G8VeAGTNSOPQ6hfPt4J5VNbRp0uWlY/3/BhrGRT6Y/1RQIp/H35B7q06mk
TQ27vd7MNqIjUNAc+W1NaOkWQDRp9YWI4YUBBctXFITbS+q/qb71S3ILpi8suMXb
cbk3tfmBlAvthHWaJfGBnep6AOpeHhPCaZQHNgJKRi/KgZaf1hhIM4Uc8LSvhvXt
N3A4EzdLmEZdgf3CuEZEBv8QpVFPVOK/GOkhVawg0PlZaHStfvHsbP3Vib38cjkj
bnwHpt6ITSRISG/kp86pTYb5I7nQ+ozNAGjRSAGvkUnxYQo12tRbqu19de0MbUaf
lVLpDoMUn+In3FKKdc3wSMIUliMHEJqdc1iY1hVEaU/+Cwf7/XmN64CtCH2BZ4rA
hk3km3O7JwQyr3HYV8d1BM3pxmd7qGfKTVvN12/G1RA/DdNMQ2aMCQtCbTGSDPhG
Tb/jr0g3wxa/GnkF7M+a3EIPewlapgTYck7B/Th6KJZW9m6RUf4FtHDZCmqLgMK2
3K2N369EuHFlvrlE8hq2flSW5owJUQtRmUU4nvZpCm58jieT9YURLB51y4/dVj/y
3ENDqo+NICJH3/2909zrW9Y7J0TnBI1/aT/sZvcB4CfLTwRj66NWL4lnSNjHBl7Y
8/H5RAuYvTVFmjvDzOP7J87ratz+rGL7XZTgjLX/N5NXr6V+VRrR2JvXdDPpMivt
IZ3itXv2VfE9w0SAVhbxsVNcekmHaLZkfJsWO3qyvDrFR5vGn2wfYMQ02FH86KxD
gEI+bjeaaRsiEfSO7r/lZ+8g5UVLWA21AUFNMPAqj3ShWxeZdFel8DMcuaQd7Q1T
MWt+JW9BNU0aNYTWTN6DpnvGAIOGmL2hppYEI3Y/wLFfSfAy/s8uCnOkoRrbVKDc
c/wNySGTDbWL1MBeuy7bf5O28hLxc1p4Ne4Aeu4Q0MujjEBwmqbSz8WFTTVsx7Na
PNWyBUSG9kx7nS5wiYLvF9nQVLmByj2nWhY3G2YahIZapA2RuQXS/cKpngPbOm+V
iBYBiC6uNzaRuEB0wBHCm3j3lVSco2a/r0w2UFj1V1pJY9YmyKch+e8tBS1MXM2w
Jtp3WWvkiI/ApHRZUXzoIwZYuytbCKw1/7/yaZB9tDGs1zy+Y8VIXZP6xzbir87k
I0WfvjIKKBKlSeKahsSPl04700r+VrC4NzbfYNSJJxwZr+sNUiLTvbitOopP/w5u
eDQrzx4br3CsaXY4mxZjxMloKrZXKxa6egoar1qTAGsBwOlthfaQM8xVRSi17AB0
Mbs5yDQuVHtF+OHA5VPxFqfl6KfnH/Pto73Z5RO0boEvoZW9YMEHeDfphto1CvnN
z3LurfZXkMnc5w8AmpUgPQrfMHiA3bxo6p9qzyNE66AuNUptiZyCnUQPhbAZjMeS
NCpmkdTcZVZJiKfS1kHUHOWxGXu8rK3++WTIaecjAat9aiwg3+Xyz3/VpDC1K3Hr
CdNG80GYSBtNrPbK4T9G76KUSxo41dktm2RKsqTmRLsVSTKVtf9AFhQBBARAgbB3
T5KSo0PdGKb53Sw6s30LCNEh76JQvIM75bOIur4VhE90Eoaj1zB2ihWDAIMiWgG8
kKdifrj/dTwNcwRRuOsC8+nKLU6/D3T7DwGmq5ciigGbvTJ+okDnivSq8HHybta0
iFKPfLrIQWvS1UXzk5frn4i8Rdykpd9OjexkdMCKoVxU9aQCh5NMZE8NnHkcFbb/
gQ8hFxWQdvGVobx9jJ7WSU9KxLZOI/Pvp+StBR1pXd+gFVvvyaMWfeD4306MnTI8
GTPbl6f8PvDAYzlNUhJEOaYfpfx3FOSXezdheEez01sDhIk08/oP8eyLiRNmksM2
jnDjFmKWLcQoRx8Uy2cURgBLcEg20zGHG8MysFgUAlqCcc20ccqJLGZmsPaida7k
nzB6nAzwVXLvWYKPtZd0gXUaG2stjzQzO/7AOk3xhIELAa3CGN9imNWc/pGupV8u
hG78UfkGh+qPSS7tDwsBsLhBk8Mk0W3E700sQiHJBvt83eIgjHKKTA6XWhcHMJme
8QTleYpRZ7QVg8ROcKum2Y6bA3h249l/yXFscWPEcJcjDxvK31hNZtxCzYJvlL/+
5foNCq/ycKEXT9pTlp5JGvDY7tO9mNTkMEpA8i6VOxL+QS4XMH0d3kqwR7AQh+/w
YYVt19M9hplfCFF536nMi041SljgqrvykjtPJOX4bib+pScA2mahf4YKAHPIlg4e
70ON0Ios54LaU+WQhljzi+FZsp7hFhakQbIspwSTIaYc25NgUASZpR/9rO1ExobP
dWV2jc3eECjIFyaBHe/fnIwPFnlaFh/VVuGTM/0ZaV4cwJnXg54Y2sFQyND6FFNP
zfYsSFKaUK0ZAG/2qjCpFZchMfVHYIVL2iXIbpcGOso5bLtxvvhveJLhIQGg73xm
S+4pNLIFFWv899ufJEn3xCFWSBfPRmRFZypgjw4L/1tUqESLGCiVuCBX7Gh/45Dc
mns7/qo3aq8wzXeaakNmwq32YPspdVvZqcg6V2DhNQ8AjKeaQxR1lS6LwZP03t0O
s8pE24YGNqxqiOrF5ujHfMe95cKBAj1cgEEJgkKUUw2LD/xqo3RwG8gWsDaV7nIh
nqbydzieJ6U2bojbY/Z7MROxn9kbmRmpwV2ReoBYMSCLKyhp+eX5M9FHW1wKiRrn
OFMS69j4q3kIuss+yZPi3DCvgAQfwzh0Igx9y4b6bSMzQOYqqd6zagfpHlq6dJQ7
MA6SyD2s32rvsNbyxrkiNSdEn0KQzHwdWU0e01O6/jPcf7uQ9nCuLNEyFeEhKb6N
jWU5pZ3NfCC8BvazL7qutXP1/UN93VwfmLvipboK0yFvnJ62aasC37X7O3ra7R/i
W2hWq/BXrq3uCEH199JagAwbuQRlJH6XVam3mpRkQ+hZCcGnM+6UidoQj1jjj0Rs
V65X12XoJXU8gS6PXkYm7yIyTqXitnnesTSTcLV4YASkQmhSLA5gUZzUl2DxrlzO
uXjIexuDHqUj6BPUDNCgRNNuYBZzWDZ6DUWESuDV8vED1sSLWO8/xFbmirlyl01j
DYcws8vneJCDNZ/26fpI9p0gtYlLmp7g09uMiHuqv+9Ur9MeEw4C6r/yBiUdWfGc
I2VF1gZKqEeQHwOxJ2qUce2EZdVqzUVkTdG65INPqD/7tqW8ve7KnD0zUsp0NM5c
VLtey0QaDlZ25mph4gDfnrnro5WZxcLBkTFBXYMqsnY/ipH1XzoRnx0l7yUWf4fr
uTE23ZlrI/h0fNFYEvVFmB+tFv0erDTQ9B9Bt0VRAIbHJNfAlpp4xjqa+S8FojrU
9BLR9i85vdapDx2gvPCoH3MFtJRIWpvqTMX3Psjs+jgiGFS7LD8a0u242ZKC5jvz
04bKiqd9I4XsP0ujBDogKhHux+wTvrw9Wwes7pm87S2d7BCwvH68FyBZ/GlRsbCD
kGXavAUemIuEKgVHuvzq/kmD2fzmVHLcivTc56qtlsg6grPVsSFGCW7ZlmgRVZ99
LI3ipNW7Tmn5vHm2dFp1NakJHz4NgU5ma49eMQl3yahfUuI1JAfVul9LOKafxRCn
46MfqIrW2vS1E5gYrFiRg4bBVlBKZJSilyObfXqFgjwH4ByY0NViqbf+16xyMyWp
3yihz6K3z72zLslO/axL4jGvlt9O857XRj9IPCZHgZcAyqPafzSXmiQtDmonOWTZ
N7xUP0dRa64qixjFmxzFRdFh/7wmx/5A+oyF6ImHsoTWDHZfj22NMmDmvpIQyfEE
SR98ECkWdYYu+yuWd4pZOHXMS/IMy9G7axymMXwynSby5yJIuxHwsE5PD0fnxOqU
dL18Zp5MacCIqdhlG9FllGBLYz92qgXUlBmK16EvvwwqEiZU1c+PH6EreiX9+Vtw
Y0umAwQr9t3AeL53EUp7uin5YI8zWzaW7DmAjUBNNMGlxaSNLV8oUn0TI+bM0lVl
C1TVF9NRCMSObMcJ6d4CE7ZdloaQMBfOBW2LRIc47nkJq+zgEZUndEmDYiWtUAu+
yR8xHq/4sx3DnnxfGP9ZCVnhngGWkcATcVseBreV7QMD4E6887jN2/RKmHuB0S2j
LZsMlYuCgpE7/z+5e99k/k03iVsu5NAUmohnGIV07j0ludM67PZRIthKyKELt1gw
aXWxRlx4XsRQ3/VXJy6Cis/m1X/Fxrs+plMRSicHgkI/sDjtLnS/RHsX8H2mHKCe
8adu49ISSyLr0JJ2j6uDih+QBrWqk0Yh3Ay1nc0bpYVUJ1PrtvsSBHShGGIvNZ2J
XJlgoFv+DjdlWihDFSKlS6xbLcc0IBqe195T95Fm4QPB+5BtvtNwMxyWQFZax/Hi
QUSxO+O7akPAyysbSR8R1jOCCVc2ZebeydeF4XH0OWwAVa1PwrH1A78f4zA7arwO
p4R/xMdyQysc4ykFN3VZlOBQG8hLG7cpU4idj/NiPIkOHddf1Tx0eYipK0f0JVFT
tnr6FiH1MyEE33jvxjE223qVbj8hDFhN4WOl6C58OU0vxntfVA0mQvbgWe5jHJ0r
HadcTopb9ekL425WPGDsVCPzsTxY8+/p8FTcoyNxnz/UElA1+NcI7vnkcyuytGqP
5ggKdRV/21tUQsi52R6Kn267jr9AWkoS7dVu0EDYXNYqydj6MTf+tvRY12kuebMT
vlmxMnP/JGfc1EOOuwqoci/Lm44BrkNXRPtbSsfW0gA/vnwmO+OvCk+eZPZPhtYG
fvkB292XYVgWnMGhydrcjg1nME4nG2zTsiR/P02iDY0W0HcgZLTmqvEBTu0tdNwy
5Nmqbjzbojpiz6lLLxbse0hqxAliQQH64sjqQ+ZiFn3XnLnPJ1GpSR7GIvO7jgQm
SKMCQ73gxvndH+BcyoUDL/agVJJgLiup19qz3FxWL2isF+LlAFpAg6oBL9AYT5YJ
/sXmLiSohuizd+V824tcSdDBq1uu+Wr3Cq4zVpOiIDfRD0CAJj5p5NtT63p0DdnR
WHmcBmclnS1QhbY0JSqPJ7hv+WXum76/2qtNuEUlvTYO9NXR3jeAo+0TMMqpEiNu
YA3Iug3hrTowh6vVqPT/ut5/To32PTg3jciPsbC1UNgwoezPzLWoUEhixDXDcC5T
mEVLMmRUT6r7XvqbjlNFDD8htXQ5sSCMR1DH410blRxKxWTY6sqLQk2PRVn2by4t
NBmIcCFNFNxTll/Y47CIN16tK4zCuW6lLQLgbS+9ox3sUslQTYEfOGr2R96rkzr/
V7K3Dt+WQxX7A/06W2FThGCpoR+w3U1wEizRInxwfy/Yit0GTwLEST6SmQI17SFL
83dqc89oefQ6y/v8XhM8Xg6LiV2snGodiThpD9gce4Q8cnrg0ETZMGTwZpOE4IVy
80WJq5v2o+zdPPNkPIjpZVa8AaVXNwpT/dlNnlDBwt38+AG0KhY6yjGfgz/frTg4
Ij7hG0VYDz4/0HEWqCzsWy6WhZzfjTuNmqeZ3QPcBKJ5Fv0S+ZXGd0VhIi01Qrqe
YbOC+Mh0r34e4RnjKQcAh3v8Dd9cegowVFNwnEjXw/PCNycpS7hsUh6No9l1Xht9
f+rZVs2bKyQsW9TnrvChr6L2sZ07odVevwEsSQ1FBalzHGPkcqtBM9dOty07wPa+
+OQ0UU1lK4qAbH4650bdgQSk2kGQ4YiHZ9VS0G4X1k4D5217ke8P7T99oBXhjLKQ
v+jOLtVyvF7qhKrP1QQkKBUvEHBJ9W9xLZ5BcbbUSficd/JQjSKl/gZkinxCY7O0
U7wlpmocJFXFCavowqaOSSY3yqHNFeQNnTwO0FIGORrzLEbHOiAQnIImCSwVOouY
P089TtdcyrsiOpvtn4S/r+vezDDleHfhX9JBjfI+XgpalAiY8OWzFDy92AgDbjem
up92r1rGG9IbM6tdXk41aKMEA+KkTMk1uwKkWbG/RCNO7UgCGUtl34K1I9LDKk36
AepRZWsIyuUGBZ0XcyhnmpAVvXM0UNCMWfoTrhOPtICSF6tapQ3FQZGXZlwmKDKh
Q5IygGCmgTGlIt1pTk3Mn6si0Zv+/bRujIqNP7W1xXo2CKi95k6Q1dD8amrTTrVy
QNYBa/8/msy5oQ8WTsH39V0GvsaDEoKiAgKv9SVpaYE23O5U1MtQWH8/AX51FSUa
nM5VbPey5QEU7fcjSoPaOhcgDKcIqR0zCXLN/3Oj46RmXipDIPHWZRfYYvRhuRoF
PfDXbiZWOMyaO4m9RbvrDZKe0OXrxszksUmTyHn+sRP9iSslZml17N9tpFd3jinL
Qqmd9d+WrbQPBpNvlkWjVeJApTRI9lbydwzeX4Mneh2tJkX29aY0jxUnD48tHFtc
q32CVkKI1YDaR2R+NU2B5K7uXMvQN32+8iTLImuL24mjEw4hEGD/7V5dHA/iL/N5
LU4Yv8doZlKfMvzqudjh6Irz61FAm4JOTUqzi02vwEo5O65j0d0WNxut5kvWVYod
fvMxATJra1Tp6DUqeFn/ujg44/+Libyk1bX/KPiMjjZao5PQqlwIRQDpoGake6Rx
L7fN+mHNmR10UuNJEoxggj9Sa0M+H0Er5cVD6pjofuuoHyi5Ah8xTU39sWC+BIhc
yDChumrSTsjPJkf4OLVIF2/BPQAEmZJlOi11TM7+wBAh1RWEnmerUFN8OcKKuXku
PmUKgs/jybZu2SpI6+vYBSKMNyPvc20hipDd7GXslq9bp7hNkkqC32XXWSk80UrN
ecgla7ExaDwHPcNy0W01/s7n84mqTeDOo5SXhpwLJgFYhL/aQ8wmITOEvYjMtmix
JVa8B+Ts/dLcO14rLYA3LGWTpRqcZsnWQfNECsvwvVJYfE6g9za8AxJDSZpV4tw7
GdlQ9+bDYU0hvakiQoKtXpSxpwGhqjjA6rt7auEQBL696pTHL3p8zfOStruFBAdG
ehnSN5EHu/ndXyfgwU6Q4Q8BdIdUvMnWX3OMT5C0ceiCVy9OEyrW7gBD/dvQdjXi
EJatM2Jvu+/LJQPvSH7GGGalicwD581sYzE1Pw391nuGYu3VpdEWmWBY96SM0qb8
vRE3e1/YmfsILRDPNaxLHaQqKbEnLJ376eqSYXuoFCyb2Ys0/BD94fEXkMoKRD6i
42h++NhtJlcseYY+rdDBLe69tUmyDMLfenbiWFELCuKnIP/D3MEr7LpfENIssq6y
jyKWAQ8ho+y2UgbZxAE3RzE5JPhgiaCSAOeTFFTNP7UPSaaypHw9R6ie77tPeQmS
TkMFyikj7fay2dv0m+miPLLatfS+o58cTa+p5bw2WFKSNFOmKfQOzBcdaYU8BHR6
ATOphOb/NJ1KplfzQuXwxoI5sHdczzXLwhQlIQZOLMRZX/9JejB1Qrt4yy+0z4mF
YB6SkNstw3fPQMF+YjxHx/6qN3O1BDxDfmfVsUvPKe4tm0rdNAQ4jT55UZFi/ejm
APjXBk8M1sLiTSByVntjGjFDQNFvdecN+At7hbIjqLddHuRAvJ+HkBA5wahwYxK9
44d22ckaLHPU61MtcvxNcMLdVJ2mBicmYIf48+nJpUPNcMv5nU60OGI3iu+P7NBX
A+gZn+UZeUrd4zzePkHDVFYd4iZZIdg21kshGGhI5GIBNHFS3MIJIsUAmjLCOZ3G
9L0AxVHvE+b5eBFhuEbNSPWonlr/XG7XS4vzvtTX/7grWnc4Mxn8IhYFdCoZPpej
WNp0iWf31a8OyI4F/+psivn32Iv9svv0tmzB2A/fa6jiPrKlNyRDM33i5vKSlgn/
qByNdIYnKnbTQDSvd4CY5aZQZCLuQt7HCfqEjr/bnPjv7CF4KCsFGKbaojrk/+w3
Vl7wdR7VDQfl9EyQGviMWYbYFY3a6o+/PLEEnPMZO1xefqLi7vuzGYBNUD1atVni
bLqky78Oeo8q0TaG2XU5TUF+79cknE26cJX4uRyExaBwksrhlYX4nvE7MZL3GlJl
xRvLFImt12tUQWy1E3M2UKoNC0nJPTCewX2ivq5oKPs5A/7fB7/rIRZPo+M14Mma
r9KA0Nug0gS3cxk4jm81PdoN6abiGWj5TY67rddfVm5y+iJ2wu21PnurtpBACy7P
4Hkd/guaI1/OL143miScalxlrPGQnkFFWttNrH80t9LAsWcQSib3im9y9j9VNBuf
AuzN7R/nJe6Pa6IzMdHZ69hum/E2Flecc5Cy1+5I1qm+MHezYnv0B7NNEa9ADPnP
GCSc3aXW/+QTZUPlSNyIcnKbYMFpmFbXFJK/qu1XUt5sybbaR3uEb3zeDNYgfJxH
OQ/QjV05gHzdAsbNoTZfPrx35vUpPoN4gnKY9KLiJNqUIihz6kJB8nkoikwNVPDb
mSPm8DGtZ2Mpvxlrtn7Lq9Z4IOosuIju51kkBcj6mLnH8R1ypLhMERbHUBdbCJ0T
+8lBT2gO+UVIx/8/fFPDr7yTOurXSqxzysVlQMJ3FwEp3k3eoivHq7XPHoZ3LCrk
j85ukljOO4UGuUa4BpvgbOQpnXH0YsxthP2DV3QF0fil2QYbLfhTJy2ssbIK+Ioa
eZ9oNPtwRm+6DPdjrIY52gBY+ZdLERwGKgvrzDKXbcxxzdfIafLuIKFjeq09mjx0
2u78Ypck4ujRxtWmnb3NQJ7iuiM6AVfWuhV53k6aG7KzXvK/Kc/DIlE/BmlWx5A+
EZ3Upz85c8mHjNBcucBY+jVcpnW4EAEJMM6CsugXXXqs7wnAR81C4L7KWzkPCnS5
+HK6cCbCDDV18Z0z4pzFseFfOlbbt9xFttCIzqOY5wpElFo5FUjV19TUC7+RrcIE
Bdpy6lgSX+iE7R2PrrYrrTcaB5UoMPj3rWlcGl0tYSBD0jlctrHua30wXlfCHNf/
xF2+pZGt5cOGxRePrr0dchxuEdzlIedtT77RNwybyZ6oI9w0ucv7OvB6pqfUo/Cs
HqztECVLh8EGdrUEICd5nZhX5xnPIC4lCpilfw2LQ5LNtZhjuM2V4PCh9h6YNer3
dsEPou+RxuOQR5Wbskx+MLgPokqQEXLpoIXw6UIrCS2f/N5TUi61R0nFmABX9IWX
fZuoTlq8Ms+f8vKs3gCH6gv5y1yvLkSaqH8W/4Xkji1QNYRwus+P9gVGsVKFvE+3
yIcyyG16LvdNOU1mZZw9NhQiou05zeNs9yzEoFjJiOn3YXRUhM063B0oMvFhNFIg
KLgsstifOtUiSN0mnYkKddJi26X0MS/a+jnNlM3hNlhiw2G/cSMdr/ajBk1adDcB
VQNRkBmrHTDoEWaU5ot0U6LF8WlWAA/PtX50TUA7KiA8hXWfV1Q8BeaRpm65wftj
2MK69Cns8ftM6jUI3uO1n9kYr4D9/4wl20J+wuHxGthJrqAvtOg7pTUEUHVJWJug
a2rZg/GAFmmd2eF26dC0nZj1jIfIqgrYBV9SOugbuFkdR2iJIM9KQBugGQffwyU0
SPTpr7SugIP5d9rBI5xtqDEceId1bk/3diZhshPLmyEPuVn9tWeknROfn+97MInj
DBiku1fcZPU2iXieOwGZIo6nDTawpoCEF0idpv1xfD/+9tLQfDFayhQomn1up8+L
he2U2uBuk3X73fnRFY2XkcljqUu+Y5XCD62Rf/ndfCL9VjHP26es8yLZUVoBv0bQ
PTgmY+eOwViUkyGCDEQUi3tlRIuF4WNIsyAb8857OWkrH1w8MYvSM0r85Y0RTN4o
IC115NdKLxfM3A8cRv6W49DYhlP3nW4EEBQfLX6bYofl6NkFN7cS2IS51GCk8nIP
Cev9HvcE2F0iauJm4wSSIgl+wqHjijN8i5nnr9zxFbaW9jYhwXJhpVrH54PYxxB5
X3Er1GCJ/CHQSl8RAi3Exy/H60xrQ709m92hXpykpzJDQvTNVD7e2wnRLQRIUS4z
OMmfIDYo7Pu3xtj2HKLAu41hHwJzmDetuFumMkWSbOqbe5KWEFxBNppX+JA4uJGX
4oElZnVO10JGIp9ub+yhGyoIm1uZxEqlOvvV1U4CdhPGoYk31jKQRq3WWGNoZElB
dB4KrQNPk7BrtAwA/KXUp0YnE7vfiRcGUwkBwR6IdJZK1GtZpb97fQiF5OVp/lr+
vjMxvuieUOE5oRB7PvBaFiGNIlQNO+eqCAW0u2IJ2AVLqKpw6AS1Y6wQEgPT7zeG
w3hWHKfANzAHVoRUU3DgNG067oCrBqm7/3XHMXKlB4lRbxtIRQsiubWRrvUJadje
w3RLos54yiDrsph8lYAOa+I/QtOL1r/YbAGES4eeeUlj54edxqrkae5iA1Dz7D9x
AXchZHXaDnyBVAptw4aHak0z9DH4wZJQV1C3eYXHENHVzZO+bUFAbykFWHjrdRUz
WxaUyJIYUPUzSucLu0koh31YWV8L0Qos6K2dG+DMumhAGHGheRLCk6XxGND7HX3N
Qx5AhlQMqTocwd2CNW+7Kx4YRaG4rYXn21zvxD+hVMW97dLSkw/sNXkavnb4DQK4
z3WNOJtN+u/KiYvez0q0kRdrOZ50JPCCyBPs6zBbth+TLyBnkvaAGCCzCe+Bx6ck
H6TANRzf3ReF3nQTqtmirwSUczDzVkXO8a96BOfqGIaXPh9bZTB+GU2Vcce4hknJ
FxAvP/cp0+019JMDpzhKJyoZgT4cFrd7wJ8siPniDC84MUrv8jFLr9HXOKh+x27L
rfjYBYrasDH9JavC+F0hR3BxvxGperRdqFXAAJXTLMrkj8EPUfuhraQZtYf6Tekv
ur9Ufhy+LLYVu8ImIy7PUU66N8Npzbfamew4VOF1VUm1ZFvAnfJxod8YJaSBdOg7
mB3qgst7iJMRow11XKxLON/T42Lwvclt/F6UlGA9n+pKESnUo3n/gOucvPH9FK6t
9ah+QbW5JrALbR2LtwS/nSexho/ZACx2qk9J9nofE2QjYRAVmh3M/26GIxVHCQvY
junYcR+o+VA01TvQkaMRw+0ekVSuG+tlXdMGnlVm4++Bjkgq2WF/jzPmDUViw+3r
jdCGZ6EzH5SKJRjQS7Ngy7yvoBDO6v7h8mesDbdQnyBU4Cl2c2kpoIUcxB4lqVR5
VVDrdOpAQxb3zDA61n9+7BgO/XcWw8WFKhjAvICAgmfRvHpBENb1YZUdMm0/Wjf4
9gYPHwQCFLMPKhBs0WQv8iQ5AwBOSrZQx4IHkE70g208L4cGRNKl1r1zA40VpF1b
f6CL+wou+8WET5HOQSUtqwKNSZiw0oL4WZULAnDn0naumjFVFsS3+czv/d92R9dF
VLwJ1ElU6IEb/dgfz96xCsoTAaoiNk63PT/wv4/slZEZVUgkXsCBzoZTNFyOEdxJ
DQf6dR01NLMyVicQO2nSBxSzJ9VbdtvuTGKeFleylFexH3nR/Cx8w5lCWHOCWVwZ
tGXvj0H6qnVVkavhMEZ7tsMhEv1F8qAz3lt6qY7uUmcybJiY1rK5Kw0znXMbC3ig
prxaGMSO57CCMdeet4MwuT3IZLzCLuOLg+cVeEk5DZbNzB5B6b24wUFaOc7QMi6/
wyq7c9arHqOBNjuI/hsFd0/nFs+NFWZtDUjh9fmC1Muji/3De0CKyNHFxuA/R872
yRxq6CtovpTL/7RJBIgn410qnlD4Hcfp4N2Sk6pKACcY4AGZTRmwyUSzzvhdwTAs
jrgIWyutl2OD1voMAYXiDIg6MZbTqjCnNeYbmrUK3Pj6LQaKAqyx8m5ujoU1tDz8
QmIJANLqS6jPrCdHH9OsT6tLhM3nYE12QGHq/+IEFbBzeaY55c4RHUe1A4PPqfVF
fIxpHYCcm7r5Btr0AxZNfdjFE2PpxKBELDxsYv4xNLIm+STWU87ZfdiJWLvyXzZH
XqUNMQUyn0GB6xt+mUJh7HZKmkCTyJOcv9XhuhudgnweYExJ2TFNh5bqY0t0mkec
ayOz/2XjA5xsqYYKHMokWWT4kYlhQ3ipEscmf+PdbezL2sSSU+4Kl1d+GcxQZDP9
g6qyELcSeA3V1vnF+5qY4cBoqjNE+Ni6JhEtoUaP2v2JI8lwb7fuGGfFKWGd+Kd2
gFH+eYg5aHMdM+mZ8FPDIWQMC3ickuH0bKTxydP8Gd4LJdDH3Xsb9MPBmrfE/aTN
vEw0vqmtJrokfbv7SPilkIHGUOeGiImB8Sws30VRZ+RFwIey9TfpgoplF6Oc+c30
PlrK2zPAXGrgE/E3ZpFjhS/m7KfyXqP4XNNhp8tjLNA+gyDPF/lUhNfdpa9ltFx2
Ce6JeyBt4a8+x7LJjoEsqjwv+YQBPDgZV8Q05h2fVn4wuAyWTj6KBJmnffZkNgSY
rxgM9gcYbf59mXM3YDjHTr+Q6J6IxKzN/DBabS6sFTXG8z396Fh06M882puGSB6A
lWGntFm3tCvuCos7zps48zWBocwfz3CTL2sLMV0V5lfyITAAu23/zPQWtVLyW1dM
5z1wzB+KUESOheT1UmiZ5cesN9XPQRcNNDVnVZ+eqpnD8fQEh0JWqtjf2/HstMhW
yBn76K6PojzRUVgmzeADfwTsm9sH3ccq51uqpIQlzI/9/UAf2qxaseJ7c0hSMOL2
Bjs8Q5tlB8boXLt5EwZ8UsNz/SO7qQmYrTuyRMAgsD40IXwsYfw/pZDawakiGrN+
H6+izL+IyBLlYUfi1zupA7K6YEC5OlNevmUXiIw1CWPw7HZGQLv1FKzIucU4710k
bprjHfjUeb+qLr1vo+CFGLU/YAKfjQson97xEIieP8ZKh8lMC13XuKSsI8A6viS6
PPKk0n6zIv6F1cjY6ZYveqkYl0U1ynRL+f2sUyVxBiAV27cjjNqMer/sfudwBziT
tY/njvRrQZ2gbqOmKHYnp/JRFPw79uHi9KVlEL8VALLKhkzxPUCGZcio+8Mp+HQv
QXb0E8ES0gd/8wwXqhw0rtX8jhj1GYd8qC8TWpBQzI5aOOz1h2KuuVv2v6Ini+Zo
xTQRFCZq/rkjAE9r+SOr4XtCiGz1tHr1mC4AlrW+XvAInHUwYindQqPZ91z2fKzN
piSTCwhn1nTQ04V4Gpclqo430yIweaMNMlDtsjFfNT2HLV35TpBrFaLV4b8LNYzS
scDBApVrrBSsxkYln0Zgh22fKOrOVtzUuqhdTs0Vj3utr7ckKmmcxcg//RMpWxmZ
Be4dYJPcwOggiQqMnsdRWrZvp/WMcrA6wfKpth2ng1pASBthlPFdknxoV9+ft0QW
3hmeV9mz5/NcjZAPXsx3flXNFBwbiHaqCQ4VOYxxyH65psolIV+iOuwNr43ct2KY
84XmGw3ya4TwZcJbPBJ0SI8Nf5fL2aAh3o+1OIvwQ18rPoeExh/zFnKe8V9eEh2V
NCT3WU1/ThSSmCFHMXR80zuWGHct8/Om61gaFZP/xK/KAmcUKSp4kV9yRC1MswGP
F3gQbYm/4tj9CM9UMI8yxo111P3mm8WyYVxdXfCodzIHaDFASSucmwtCv85rSu+9
QeGimsFx++0A/YCudX+Y3t1KTx7B1SjQylJrmsNnEuPGOgPSG1USUItRhpJj4Inr
2YDOEXmCPjBVPOjHTBTGqksPvesK8xRCEwbkg9Of2ExcvRrDPgcQs3+PXoP/7hta
2BYuo8YVPJ6XCUe/80Bf+e7Tonq2vrPEPbncmo6+QlDN3iwPWFt5hpy32z1inQo3
u2e3fkDia9D3UALU4IFvrc6v3rghjwj4Mf37X2oMSU4zIzRdRbJmpxQaBUZlVwMI
SJVAeg1EPf3Ye0Y+ssqXZKWAtRh8ikL5j8/BAivZv7CtJq/DTPvWAIk3Mcu6rDKF
jnGQz1OjbFf3XprLkZaaWypRXm1fMRBzJ/ly+nE7dSqB+IYs+2MXlMh2GuFErnfQ
MIYYm4B4PLor2/1P16ZS1so3QkEijC1cSLFxTsZJRDt7nY27mvJ5x4mP4uLRhKfm
kwCbbDshB5GfZizjOs2/epzgql219yPyYpFwlJK9c13O1g/XMsKIo7IFJG4C+WOW
j6sy2ms5K9wPtUj/4B5DSnlMEfeF4SN4ZyUfyod28D3wOE1/6YxB5Vqn6NCxLuHi
NtyMjsWgAwt1d6wDurEjohopKIaq1CiVQbq4gCAeln+k9IV1eGYmBxli75GYvZFD
+yehQQTrneubUhMy2iERRZftDojHjd2Iaucvsd4fHFIgPSKXvr2xIqjEEIYi/PO9
ivTYaEvMXsCUm7sc6g26NEz+Bv6yce4r5ZHUBVQ+0x0UfXlOq3rONd4zjciuHXRh
mjQ1XfAqe09BLepUgAzjC8Xl4Eyzz+aMiUCTZ3FS7RWmNP0CbdG5xT8xH5gsOD/6
3rINxdALO/2WzyZoFjj3DBZmsY1DKt7kMVtSWdrXhsy+iF281PQ55rY5RTiDK3Mm
4CpejEZidD1vgUZyF7JgDgLIbXlC4WL+ayFq1+9tMjyqBo2BK/haOxrzO0+qEs3r
CkJ0ntTqcNVgOsedZhwmrU51Ozme25K4iy6TF5NgtaQtoTsF1o3QrPd+zDD/2BND
05hBtgpPM8gPyWf637AiKU9lGfwz1Y9ka6Wl3P+LwRZMmY0HM/xdSQHVoggk4LlS
cDIwW4lfuayo6Polv5n9IfPsEDLFnqeZQ/ohW2G220XJncYyHTerd/tZXwVNW5Xd
b14LULWKF1jizjEqt86ti92WihcXCl6gOPDOqxhfLEUcMYgYRjfFRlffZ4G1ZaqS
fuhewiB4/5JbaSABUnG6kt/M0OL9xIc16tIhFW24tlPQ+9YCr5ULAcAj8Nu9m5Lu
juSdnzoSKNFtqHHSdpv1mTEk+LS8NYnsdRhhwAEUaEWNSxoZSADfcoY9YJ5sKqIB
Tju/0xI1zjETuIUAffkDZkcUVsdl15izBwFDLG0kfmTyjuEJmKbKs5vcI8YeNXSP
McbAbDz9qDra+fLXeQPHljEXiTsjBhTS6caqgpve6VZf4BJ7V1534h8fT9qOXu2C
AxgnXX2envxzcTFmh5k2uO3v6bxs+x1LHiPKb3MkmZ7Jxu/VTCCfhAXZMkLhHmtL
Yjd5bceSR1X38EK3KIXx0P1t220m8gvJkZWqRBTnirOHiSuJyoMnHw3PD3XlPa1c
pO4TG6tslPnqkm9wEFE11I/wBA3L4N1C1qivL/irQIn5F3fVyoSc1bH9WK63bUB/
C+ksiShFBxLxG4wzXSruka1BZgdRUI9EQhSY6f1ErRjkJbht5z/fbWeL3vTrdJzQ
umWChCAba8/q8Oo1YiSTtWQxuQRRTLfc5s8EJMp6LqDE2SCDZbmpVjsgxQrI9dFR
ahv47DmPgFaGSnZJiBtTo92m/PNCc8h0FUpg3qGMyipHY/xJCP6LR7wX1EQoyLCZ
RhJnTRU9yI+pK95FEmiczua3q17CBJEQJOKgJb6MhkqzgK1yqgmtYybvjffVtceu
pvHoKmMsS5XmegMHJazgpfoTACbS8KqWQwAQNa3xddiWXWeB7qcN/rnMpZ84ucLc
q8uGjFjZkXP/dAUClKwPzsER9ObH1rcBxYbvhARFJI4AGD+WryLObCuyJep5dSLv
wl6o3dQ6JOrHs6hfDIMzA3gGLm1b3T/2EzqXhGrpKSjMfBXZjqOQKuiiHWyBezyR
veBecGWmj63e5IVXEYFUlYt3hbFPIg2O5mL3mNL9t8fB+EpCYTAWtPVzV8USOyji
dmleICz2IcRQ+kkD8+GtRRse0FwYMIQBDayIIljJt7ygPKxQXZGVvq/Tb0gByysa
3K/0pSMv3ZRcXskJgcyNoFZNeZdRaJTHG7kkJtkh7HgogHxx0ZwHgYS1+bKdPKdf
ccMWO4COvx/JAHFAmBhOGAyEPHSjlSErAMhVCVzn1NtwY+iJRmYJuWEm3Ta+1vxv
l6quUx7Kc0vV6TQQdCwx/DDkR5BwzSeiq2BahrZqUc30HiAS4kRaUGiZBpDkjvoK
LPzqpxy+x8+NAxxTr8DXV+yH01X1CJoAybocRkFWs82ZgQVU0upUJEduk/JPKzkc
d3k8mpmy45LC5Js3ou03WmPkjzAsz+dalzBxtSrYjuKqYcN7mGGCQlFfgvXpNaIN
ZjRforWeNxgn6134vcXQBcL5ELWc8jdw9FUpBaKBMpIGLODyRYT4dHbMAVoc1n2K
kMPVDtxDy/GPNGi63q2Oatxp/C3keYM+NbVfHoxdn7JRFnCt7dDKFZEpCix/VTBk
3USxA7N25MNEvk4GifgQeAJTo/60gfCA5GJmeDygYLzwqCzmCraG38VrtNzDtIAP
5WBMb1fuO1eraCH+oVb0UoTfz0t3qqxoIahFpKk6Wd/gI6fQ10fXiEigbyzF+oir
qxFOhjTNS8qqSWjZ0ntzbDOB/Q9bqFfVuOfcA51afClibjRMymNr9aV39tzcT9FO
yNPp9z2G6MnY2Iv0ieL5P1IGw4zwwaBC+rcTy+/74ZFJgIFI9f3CwIZNBDF7B1VM
d3UFclP2zaSI/44YX5y+UTSZSfhj9NdcjO+G1NDvv3XcyAGxhJXXClJJpf33e3PY
2UaslMgbaTbJge51yErZLR4M2wLf7t2Qq5K7Jn6wFM3gjcD/qJjyrYeqBSBLccJ+
eTJA85FOEo0SGDL1U6BptYt9CwcSCk/Mt7Wb5deuKOKY0VzKn1QK7yB9zxm00pIl
rGS91PQIONJ4Gw/dmEzqHEBx5l6/6hPAIPHl5gug5ZkkE4OaRNiuuUaKjvf7ICL0
ddqoeVu+Oym7+CWU8Rvqe2M+uvtPZiZLRtw54OuZ32pN/2NAh9TIt+8Bl4AmKAk7
saIlmUq2bRaICi17eosgILZJTbAJEuFFt+zoW/GDn1l0/EKUvQJmWfxpMQTYPgAB
qcxb1iC0OExefKROykIxWHmB4CKz98MxtGYJ5Nmg2Tq3MfDD5khP53/n7nYdFBqL
SAv16Oxujo1jf9Ihq0de01DBQ9S9rmJKOc5j9diWn2u0Np+aAQ1+SElMvSzHj+8K
3ShJLgS09xhhfRW8LRk+IJUYgjmNXLik4nwEqTCKALxnxYXN9WyqRHcs1UXuiYSH
fAQ7LCEPFUNAMVUkhVZV0AZeHjEddqGS7qWOWqr0b46w73vof2uspwwX1CbXNBZR
149x1179mKCS7M/r7fk74dVsNRO0innYqJR5OT1rYBPxMKbzNHZ9j/+9/n7uekzs
yI4EKuxHgE/RrpuuMDQdW1PFKJybtvYTftvIDYhXKGtk5UHumthK4dqtdduXnVZZ
g8zdLctyDXHBMU6ggRAc2um6lJkcQO4X8CGKv3F7QQeaAO1CkEh9w4054BHnHrrC
Xov33VGxpiUrV3ExPyPCYsqOXUjjbldRQyO84Vwcc5Sc/CDE/VxPYmAXuYektkMG
GUz2a4CqyMipfi9ZMzWaADOnea7D1G9aaP5xQqGX3oaEq2ymevwL/6ovJiFDcTQJ
NA81GkW9qqqf5+FsL7NYspHdQ9RQvv8gd2/vQhkcUxn5xuumM71erTl5Qf0Mqjgz
T+KtxjDmUzYdE3vqcCb1s+DdhMveD+2ureccPUVo4zZnPJGf17pkeG7Hv7AB+Xn2
TxsTWZbQ8ChbjQvN3rXV6nNsyKsRLD0lBlY40W2exJZCXtOmsrqKBKw+AKLhpCE8
9s1woKrNjgR1UTNMklixxFXUqdqOtqbjgiGQPrcpJEwS1QfP72fkfZWFvhpZKh+V
S0V5LR6gl3ZQ2ly41OKEdrri2UKvMhtP4/T3gIbCKI38MTg0QYpJJTUICjv0ZlJg
gEBE1DFhdiKhnr8xew54p4bOJn4T+Slqo3DHn4KQOQqTg210lU0BNJKEkZLRgK6N
JHRoWqc9xI7YXEC+f4eeUkLawrNYsXL+mqxhIGNjQr4Sq/1+iO9/vXDd8yrWQoh4
yqDeo2ZVKD8ndVQT8f3UeOMKikTgNEAGTSi9tL8rnGpoq3Fwmb5u9KoZozfgJOui
rzWwhTwOMMRtqwKjndm4bGuhEZBMMlA1kI/CrkSSlgTvu9u5jnGygCRQXvH8V+tq
EXL5sYBfBJlNMZ/b7Gfk/Uq1FUebv+DqTIAw30HtR0TV7jKEn8R7htGj36ZC/2Tg
0nizxipE9QJADPFOgPXJJpXiFk03y9KWtYpFx/wO0mqmxioorhIQI8L8GEm1nFi5
iQQz+KwOpPkkgKhwOyC+88j7p7kwkD62nQd0L2P/7lWeNxyAppLLYqXKhH+yKKkP
PNg82bPDhKRh2l1UB2PIeFe/f2GCRWfE93s2bGt3OFTvNvRJqISICQTroIXPsZqq
sALBO13tbQvbWCQe4PWgVdt/Fv7IDIHubrv/cSP5XChUWPA9AbQZmHK+68zMeCQx
UFNopSSsg/VaM93tkaShtvTPyc9/scXqhtLS3GOxh+jfVpPetUsXq0RaOE2tT8/n
fXv7rLecZi8Dy1068awgLida7HibRLohL7eTgSBtp5MaXIwWv3MelvRL8zWteLMG
haDq3qu/StEke4y+D5EUX8vTrCiIZgo//msJ6geq4HXxL+xVIXmNiv3UctKdUQm/
ySjzJTSStk2sAXtdZzIVhw70dtqnB5HfKqyILCObL3hfmlAWTZSXNWphLNdiKo6i
oAP1kEv3qophoVu+KqXPTbqOpSwELuLmJoTCBcdEbn7pGd48l1NsPYim23AQ77CX
59wupSpDQM0TJRN+5cnNsXdjTF5nWljG2HC6n1mSFNT3yZH40ykOT86KdvugUVEV
4ZDbCLBgEhKa7EAY2gT3StrmK+8wg8wwS0r/ODWqfCpx+EAbMB4uvH8HSoeXjPWR
W1YVBpuJW14UivTnzbUnxPPm/0pAcYXAjBV6k1zhyePbdP90S2aO/5cKCKFrRqTi
lGlnpXyuH9xpJtLeu9jTey0/zZx2+/ljeI31qPj9rhXBsQNcoc9/bcRm5vEtHIRp
0hlWdLP4sw1h/fe18HBtG3u3G0IYuKr9qpEnPrHDzJfGGoH+9MhFfJswMheKMYP5
vEKHXqw4mkvsig62WqFfxuCi1nQT+odtLPUPvK4bZ8FpaEYf+8rjJ1z3KPX2Bt+S
6UDISzf3+v3tKVcQzLPXslQ8ZpIKY3ODH7pygX4Z6u7Wt7EmjLVdp66585toLJwx
SGz18plqgQaR6uZysZU2HpayKDox5Y40/2XUst5zJbpCnMORP0IxQEfj9mrriNy+
S3tEeoBVpzqrjvnIoq7ie/sGjNF+1Hct1C99Z3VP/QNPvMBmwH3/tx2ofaA2VunM
iVQQg+fSEW/7uP0ihMXMw66HqBO6CGptiTFFN4Mj9hAMmzJwIEtYBbuaUioR/Ufy
1WhQAJag78qTfE1D+xl6acVjzhZ+83wmvFZ2736TJ760jFNjR2NP8UNJA+SGcqa/
GDFypt/GnxzDJW6+W3CVlBfLa1LT12iMQYZUMJSghnECjF1qY/Gg0h6hSabNg/+A
xtm8et5uLOH6DQ90QKICfTzM3R+BKS1ZXENNJqEIg4ScFNHOs27qo44N81Tq+3KA
b4+ihVjo/OcZ9g9jjN8sjVAJQ4hFbhyypuwRMEBCeH6aU9uHQVL3MSzZH3rrkVEK
z9rkFbUIFmvwgCeUz3KRY4UnA2PL2xLpU0x+VWEjhquQYnaOrczfleMLhENvlwT1
TdLb9wDTGKMVvySZz1QqN4Dcl0b6DtP/pKdyEcSo6GmgK8lEJJj8lXrRUq8yMWmF
fR5DdnIZhb2/3J1dpWDj0Omo01U0XGHEPQ/R+C//jW8ETg8hwOZSfmOpEjq4S51z
k87sQIpNYuZP4spAqy4ybAJOdKC2QgZfrn7eHexHuWrcn0tXkMVvRFd4HFLODvt5
itc9Q2lHWsHTMqx4Q2bwFDMze+ktsIrP3MoDjQkcBJdDuY2zULkP8MCOG4oYRpF3
tV+rEK3Vc9bbqST2l7rx9rcfuqxVXwQu6XD+nsII0eAepNH1xs1nEGqAQmnCjblp
aOjrJOVA8+4oxG4pUC+Zu4KKEibwMPnpPWBiIyO5AEIXvSJkv23S2O+1BLoGHZPC
fVuPnwtCQTB6XgOeq6VjEfv/Uk+PLj2IQ9eACtd68oJ2/anhIQ1ihgwAMhGdsd6D
lp4Qu2ErsOw17r/XQ+EO293+b5+5D6o8pHJK0G0sRo8YGIADEeo2rSQslEGsBbfR
sUqJBq1XK17ANuDo72VtBQaotyO5FyT8LB9ko91ozJhfUQEOWm9o+JRwwSnSY6pF
xo4rnz+lXrAJQ2mLmJY8ShnWTcODAKAIBkYRYjF+fAmFxl6H1QghdER4nOLkxrLo
qMdEHRqjGIsvi8VAnEm8wVsFxCfMe+XxVpKkgUr9FeiMFihn/WEnlKE4MFUSOIWJ
QVVp06lKzElj7lZkdH3QzJr/JSW9XwrC84b+l9FTMYntpbNjbE/s2NSekeDhmkDJ
ocx3w90e3GuoxXQ30U99ZG138p05fQjpNGK5Upir3QYlIhASYG28ITB83FYVQhPM
eRKtDpmGpNg2gtFfUDs24dEtX52MXN3HazoYi6aEwhabh2GQcdBp5xbL+i05f0Vd
6GRHrvmNoyVJGoBGA63OCUWavyF0XSO3/jcQZNJ+KKMnlzAeHa7cLzBoZpQ798km
qqDDMxnVvIIm3tyJU3mq33ACIkcB9XPtbGCTK+IODbV2qX91qde8bZzmJMgmVUjj
AYiG35LbiooJS/xS63mfJ77Tx70/r6fCnQAYEuidJyI+22v4LkBlMi98aOGlUrhk
mXQr7SS5Vx9KrUzfsy4w3hXo8720bNxdV8FgNzlOf59dPW/gHtVPiqWe0efOEHrH
SKG5tb/wqugRKNsOoRS13mA7Vgy5jeT3z0hvL+lMjZL/uqnRdBoVNOrYLpFCtMdc
6ab6a2r4fKwPFWsidf06CmaJPo7ePDS6e3fpuB6J+8ZIl6QwLOEpypbvY6jstLw6
Ojny4zTvkVyBhVj+2pBI+SA3Z0ijB6JKhsLvR0T6HAr3dWDF8s0sJiVIIkOAruBj
8nzzF6LPbIifWLM1WKIObY9HL2hSeW+4Nw/w9DRPYqG2ctlyPLkk33kGN9/44Wqv
kp/4F720QJWcLjlTjy2s/C2ZmKzCEOHg6m8f6RRlQZ4WKWpN30AyB5JUvrdO8XU5
MXve1LaGZqbSwStdlO/5YhMX0SwUG4MQIdmDnZoT1p3DmK0dDmi4/RyYKuMW8wVn
Ux/uwjWxhybr6CYBG5iQNfv28lXj8pqsWHHPxo7SLSynil2trOpYKTCNIxqVVcQW
77+0vCTgXxUw94j8VhLpf/NjX7zNH5wMLlmj/4u4atkffeLsZV0AYM0FwWX84MdI
ZAsg09KmO4qNnllyv6HfdL6/2hIKbnNJ3v/jkg0ZWRwv9xx/sRQ44xXh19lQV9US
eoqMfR/sTAR4xrhhZkhN8jRd2nnPx7yTipZd6mkhTU2QutcCql9keJA3Ww04yIJv
BCPEhSCPxufeY7cBbBmLUOC8bU5NyN1lBAsq2XOB9hdwqDk2opF88W19m+NaXbmE
EG+jgIj95v43WpDM/7pAJL7USyH3HxBO72J0X9cElWn9Gdp6fN4B8dFZxWulOg5i
F2YvAz3K62umPQcbjxcEvIQwJG6rPA/7Bob5FhF1pQRa+M7cPPt6zvDTNfW/kcWf
ah9WG6vNLW5d63DGGB0vkIQx0oz9CXTcsxJ4H3ddZJVkJSpeIJcIrcgdkk8QLuE5
lBZb2qDOkm/K1sNYvVfQc+qK/y/nWDlRS0cDU2qCHEnZPexGS/RW9fe2AcHQgYaM
qQi99Hn5pZ8jdO/JHOc0v5yGpB2LAIK6NSdmK0GCE4Ur/zp3ZQ2LJjuB4bflpH3R
8eojHsuMHQKgWHPee4+yWaV0OvWOvyDW4FCTuO3Tix3YTPAGwoEGqtEGXdmPT1Oz
irSgJD9k1W68kEkO2/jVVz/M0V+InseO+aNhZ07wIP3sHuw0nqBGRrGF14u2WMrq
TxuBKOSbc52RjtaizemwZHHY7BCpq+KQEkNDjzeu2quxQh6m1UWhGe1sBtOLF5kE
C3/acjUI4nztH2YaFjLJCirhfwwqOz6LyO7NaJlg95dct7BE016WCcY6NErg138L
6COlWxY+zf1XMbi8ow068Q/ukN0io/CcsJXl3LbIJ9ugsN0rUG5cIzwtpc1KnHl6
1Vww5wmW5yH+xrscZsEdj55lZ/woVu8a7ikVEP1hi40YlWxG7JN9degzPBeDenct
rw9JGvDv9Hvm9s1/wJ28glauxrh03ljRlFM+zCok4HDlSX2zk7LJC249yFnxh6vt
lUH7cdMmak8aQQ+a01Ry64IhtA7SGa/bRr8ty7MiN83804rXYK2I0hqMY8Dn7qln
a/3KhC+V5cfZ1UuKuxpIPpVDu0+2e4oruKKNFaKtZaMD/HCi3yJ5AhHHuZ6QI7FO
OeM3dqndW9YqxKkDGlOWZV1kIGyogD0ss92PIYP8FTypyCihBSi0gVLE+4hadXFq
+tc/HLx6dUhSVWOX3/VC9NMwYVd1IcjaIfthZwqRYjRyyds9es6iyRwci5gBgIYC
wmI4QduHH5BlFCLhw43ffvcFDHFgY9cPjkuXhySgUNcs6lDnxGpNshXzwlrjmDxr
8gqRY1tilxMKEN6mreiCZZEVhrxYpcTi9Q79yqXrBTP5ZFBu6llkHwG6Fkucoiqe
PCaMHFjKK/m3G3oQndMOtQItnLnfdM4HfUknsFItyOtFAAuvDkboJzHnUdUWmwRd
5qm/i57xPhU9vvSr4i+aNZig+4p9zdp+6k1SjrpBx2/wXMuIoYixvFsoxaA+cWce
gqraSYysu2aO5yV26DpI6vkyM83W4AG8+v8nBpKFXsDfKnDu84wfgiW/PPPFiQDN
cotW4xTsPAz0HJ7i3kXpej1qaC/qE4UgCU7quQbTJZqFFRzwnzrgSe/5pB3XDJ99
Kp2uplSIgUFAXZAew98c4cxswuhLf4XBMQkT/gfMuY9tP+0XfzXpn9eWTVwjKrJb
MENTIJarbXoVj4vCj0g9ydNkOkDMtp4H9uwjEpQJVH20jcgOTB41q0Cor1XCUEkB
QPPkLpL/vFjXUv6JCpeRP/7PaGknRqWx/eMDZTPcm0bYwafU1NO2OZhwqPobPU8k
cR0MzOfwq3zZjbBXVUUsDhWWkoxPS+yxh5nooYsZKJhgWHAaedthJdxvUh6wA/Q9
k4yRFk4c+m5Ewlu4n5C6Fe3E+Qngj97x6Xx6ZDrr59rJ3vkPW7mXebUdWB1pq4uN
4oVkB9Hr8SYN7FUCH0b/BDKD1VwV5r8a06tEW3QwOYlLOn6F45we+1RyJ2sNtWe0
d82/pvGA4qWZ+o8kmvEdzFHs6fqwD6idHZa2rncFOdE7Cd3gtTyAVukSufIqExEP
GgoYaOuoqosLqblkNeKmBQiQoFx6PIPUmI9Fu1dDNs9gA+KE9oxTszKuQf1xyG3c
lrD359Pucz+eb/Jv4/zMDG37I0gSwj+mmGJIeQkVknWdol6rCEiWxPVPLXVepYJV
5lY5HODxSBOJWABqqLNai35//QnjKyGQMnX/8nEeCBYSsNv4hgwqN/IUPzqsxi/1
XYZ3pBCweDWeXdFXN59qjle2oW18LH/zUO8tzM7KpI/2BOO3VMRmxo06CSHJqr8L
OtTc+lfhcpLeKFNb2Y6sfTicrwESpKMrXeIvsh19SBw81cFaMkfqtiJhFctQTrec
N0CZfRQCw+M+q88H/87kzl0sfo07lFLWt9LeyKo6z7VgzFtchaFXrQH5r7NOjsmM
xOWhriYDW7xnPgp/OwcbihlTSQctBx1S2nH2sLvpEft6HW4JmlqG8ssN9tPTTZrU
QygRkJwaKPZcwxbCe/i4snlzK0Qs+tcNGOwFto8TAdOwn/O5vgcU7lAVs9Jz6IYj
ArF9lUXOsIitCxcCR0r9dFjClPINpT8Hy38GC8tPZLqwHw2ZS3rQvM/+sLDJ8fe2
xZsUFHuNu4FNLtM9GYSESxe4cjIyG6Ftpt2V2SOyDMHnQlHXqaIgK9xP6s6OO+GS
hWf5/D+IhMOt8JZnr/r0zAIUitkI7ASX9g6w1/ECR5H8YZj04afTOfpjCPdmWqne
rI+gAtpoU4oSZOG3m7/raHh1biUtnUCyvdiMACmaprjbUAkHq3u3T1hyJ5khspqP
DhpBHbiHWrv0BOLfyaqR8Znre4h6KB2x3AIEEuwMo36SfH4XdJwJtvXQz563r/LB
AMG+uHYIPeGEw3Au0x15srH+3uP8PYlGDrbtKggwQVsTILi/7r6NPPrdS3cnceEI
SKMwCcwPRC7M1XBNprsuyDucQnC7+gqpnpx+/yS1qqk3ruIJDTdh0BrFVk2Y4Q2k
yeJYNIPjMxEsBVA1ax03yscYB9oQYunroXHbQzK9jTPfClriZrSD1mvBLtq7XZoH
mEi7+M1wx/L+MmeThqtPjbbe5qkr/g3oGUgUzo1fNgAouj/H/nHYk57NBPz+Ghh3
lFJpKEKusLkPXv9CYV2KodXsb102AQooCEitrODy+35Te5dZ2JyGo8TOUuI/60Zu
x6PqTidCbHTb6eHf7EWTWIgFYiHtSN1+SMmaDiIt9QyH+6dBtw3cnYPII7rrHdTJ
AJbOI9LO5A4HdKB4Hv+zJNlSSRqNxqoIhneklr4IRL2YGF2g8mxc+mxtJFYGL3i4
8POF+I8IzmYFvpwlmuZ69WX/yFZm7Iih/2VcbCSyFk21X2VsQJhhRmnSERXVDu5g
jVxlAj6hfrtwGkS7AGYfcaE8wC5PSk8vgJiZ5/gvl56Cv1DMDp9Pwg50FPB+hSTD
03k7dML82RHm2h2HrCSYVRGmoAw0x6R3DBe8t35I7d3dT3pJnvvP7bC/xS6jGxZj
AASqlqpILQmbyaME1Wx0exX5CwGvyeUZThZ+kqNbCl5kMmE/BT8vs9N1V6UIJHiC
ZvOaR0CRSAgQAi+6oTQqTm4TQZqX9+JtLLuHGXcF9G83BeWJqMTDq4vrUGOOGOTn
Jr51cBUidv3U6+rLz9loK/ZVd0RaqxPn8rm6FjHizA0gB1LWSja+CTe2bRgXlxX+
kwirfhu2i5uoKc5h8m2ImKuAuWbFTpKKVrP89WvtiJn0Up0Pp7Z1fidIRLegzSkB
Z0fzp7jpsx+2YnOKy7/0MR2PUHWdt1xkhLrsV7H+XTONX54zlTCQUhO08/lLa/F8
lBvVg+BRDTE0j3qd1V5+Z8P9AnGqL5pHsStyaP/C0GT0TWCs+Glod41i+ZsGvO+F
hS/Ni6pwH+o2ldLSjzKhUw538JM+AScn7SmoiL7RGhKooQZOuaS8IfFDqzkKMyZT
a+4HHYitEAHnwz/sLbEXXMcQJ59NpWgSLPGafnE2vOvK/zvEQnnU/i0O4M2f2gdL
874sIIqwkV9NDh0vQ9m5ZIiYWxmbEfOCx8yzz0W4fAhOWaWl5EGsTCJHqukbi/J/
MA/D94XluqDxnVrEYQBjb8/r84xTlG5kPIS9LXRhnN5nD5XkOCzI8nnuQaPquzhn
VnwhwJbPeFiqD+sAgN+4wXdJcJtXTMVOt+U+/671oBP3W94+4LpYdyd3rXcHxzl/
k/7ElPDb7lXVA06WTqFQG/HooIAtdPrdBUxI1gAtXgf4JQ3JrAJizJmUBuSNrxCh
uTdvyNiyoB6LiwIVp1HgQbFSp34/rf1WOlAwslvTOfcuE7NgmQxSHJE7Gh4czwBn
z4iezthmWnX5Ahm5G4DmDmt2x2emBdYaDP56U25qkjpKNDVla1QjSHqNF7Ic9SPH
dZoWhsP7rlkcSJff3KQ1KWW6CS1QdKLzZ/uJ8VnQj6cHYgVq+MnoGsJUVJJwtQ8F
kPf6Bwwh0E74FiWYHcV3B3URnKFPXTRKP5qRFtWpnmC/YGhiMECM3pxvF+n+wfrY
JLbbPaaGdTfuz6k/H4LVwtO7pR+soboweBhcB+Y14bvXR5VY9yVUnAccmED2BiRm
aG9mHf9VoA1lQ3gjgOvGHVR6+D3aKYDErRxl5fPbIey+tE96NdOnde2MFBIFuo+T
i9euquOHw3GXlCkn4YxwDpy2X79iYKWI8jKMCjk4WLCboyYzNkBvQ4QCENBaAixK
P17H1xDemoyfJBBtGYmJmkejuBaazUVRjsv/8sYHqZcf0UlQu+ZZW0qtcFTCvK+K
b4misMV6oY8jsSR/nfQdXxodpbCV/kICxmquD5ml+hlVJojk9QJ1C9Zd7UpLDEAy
/jAcZBTYQxNjyHNgXd/O834SdGzDbw2+Kd9kmpF9cpIDg7wp6dt8/AFM/iLI8QuG
l8e2RDGhR2zEix0bMHXrslbjkCQvJNgcKTpgu9iGgVEpZNzEUK/SS5g+xUQuJx0h
yGgZxjNsZmvNbo6YMI/twfgjZwhM1CABLwxK8TNbuRsP7/5bLO2KEgqa1SfPwdlZ
8NK2uDbnHscRGLds2bB0l1Wug8XGL78RPePfNDtbWspKRbIBctymmTLM4nbejBXW
qzr29Zcl6xpEAb/EI6+K6z6JkxWtxq+XptbvQQ6T/98i5exiLSRwxr05Nn/MfbME
ZKqnEnWUEbY5Ahx/mmV4/Z+OHJVAiveSggt2WtklDQFWga63blJdV+q4VpG7BrdB
GE0oXHqkeqkMzlPMlXdLx0i1Z/4Mh2UnCgeU/y9zbgS2SaSJqvpzpTaSFSF+uFVq
qRi/3+t9UGQD8me1OkfchLkvtnosaOcPWfoA7SpFbb+wn3Kh2P5hRvTUiYyZISdd
Yo/EpfMUaw0mpXk0MNnOvXjZVb9lKPFrQ9dUfPTlps3sov4mZ74JqMNOIM3hqzCP
56UygPpykbi8/9AwB9StWABHlX0lcJDnKpfwGybk0keWnyK0vPkWTBrfE1CED9Ab
odUWFlj1Rq40zOrTJoWvv3H4DajGHGIRTk24hdMMMUGsXLajLZTbIK+g2IhPyTwU
w8j27QlZphncYSY7pLx88rPoz4HMYimbY/XsK9OGDYLrVf8cTsojlIvhp6D938wd
J6GHoY4o9AAXp3ZhhSwvL90sJc9cZAOwehIVq87Zx4jFJkRvfF+30DnNHzukX4Bi
Q2j+yQMhRoZ7EfbLeNiwD+TWp45L1+vrpOY9RbinWywm9eqvRffoIEGOIjFYjDgQ
vw6gRON3+0dsx17ookuIh1NQDGwhw7Zg5JQLRIPDRVh3tUGlmBwBCYxvf+0Cnpl4
g8kV0IuAfaxX9hrAS08TNwcG2jyeWuYlfJA1S1bbn0pdvo+tbUKnQy6ssH41tfog
39QXJS4oXnkKQ+AQAOXpYVfoMj6pVcm7ohP1Wl/VrUKWmpRnF5vqPJ9RmDxEeKp7
PTtZ3egd9KI/ox3XfZFrZkWEvkRxfVElBXtXr8mkrMFy+FRsnf7zItyy/e0Je1tZ
BSflwg0fESRByviCe190UztvQ8UhblCU92w183VUy0TUwDEND1nEtJ/IrFZHrREo
HUgrmh30byrp4aPhQeqQkS1PdlxPu6JG5LKRbl/CwHqDWpZotXRV85XtIKojWQPn
88ritfpuyIOG1f4NrUN6+nF98kdE35OMRsmqn4zm1WHjtAx7cSZazkcz1ApwPmBQ
ngscPQZZ3f7Hx4f7lofhSJ+7h1fQ+mLnlxdwJPleXMdaadLURQDgLVumlnNe8Dzu
NnMa+ufhFkj/8xLM+AaZyGgbLuYwgZWlOvIQJS+me55mom03Ai5c6K6HsG7jaXu4
p9Ftbp+3h2gN1z6tDZUfifhXaD3nDz+5q4wU24pavvkiHUhHxSYzYEmWCZuqlO4T
whjTnfjjfiTHyt2ug6NiKHjO2B+EukcJadU2Lle0nOd7o+iedzELmkQZbmRjGZP+
T5/zKb9Y5Z/QUrjU2X6WnfblNsO67sl2PPCdZZ8RRayfXB9r6xo8sDJioQhG+yyX
0LE8fUwtpPQzVzPLwrnoUxEaeQ5VfzD1BdDW0VfYlJSogajmTAqO2ngzYa6uvN3/
cOPla9intw3UjRfOX4muxAGCzI/KI8AeyDNreHnIiIVfURQMu3vBHyOey2JJcTwp
n0iaIh4f7enbWFDAIIbx8wiaStFaUtOKyFulqsiaLWF6sDY0j/fubrW7Nz2obYVH
5bzrKEkQhuhUI2PuG3h1kTTjt9hnJNJEYzVTI36jnLS0mKWUlCgP21QAz15n99PI
q9ZBR+3pf9B1BVp4bRI/QC5/zpIHavUMEU5dYP0OH3r35DOWd2ScT5fB2R3PfHCL
zeG1umkZyoBFeBgC/pOUb+YlmtEQZGOBHO7y8lUCN6skcKwl04Atp4A6kJk2jQxJ
DdRNe5yyNqr2t83+YMIJAFqKUIcSxbeOozKTubD28iU9M4HK1oSMQr6zryFzpvnU
430JQgeo/UzeWOv9gaS4XEeH23uHNML1/tqf5pJZRg40TWp1fi+cmc8tP7f1izdw
2oiT3NI1d2OEP1hp5NpwEoX5yh9Vcm5KM9PWkUemY7XV3b8jGfwGcHddTuYGkT+P
TFtpmdm+UemEB3ALkp79josLmLMzar5sKgQepY1uqoBSzBynRtN6RsuKxmC3IPEz
qOhCTNp+6WqbR7Rv8gP9kD744ugKLS9JKC6Et3pJFXZNBj/Pz9grOGFCZNk1jBZC
IEQduIogR2vnSO0b9sVdJfCWRsCTNopfUU7AMZ2kDoa6wDPhckH3v4iUnHGagsfz
ZmPxxgr4JTRH7urc4+5kptyhmWhsbVI0dJqq061qdd5OgHKXIWu1WgJZpBxLAq9e
5mi4J/kLsAhEz21dBWdsghjFmoKsigJIv6ieYgtYljVEV5LvBut0CYVltLM4kS4H
cCAD8pCRdpwZUr9ZjTlNBdFpE/7IPgul9ztcwpk3dsuz04ze8o5wP02LcrQmluNi
zx+we0RXNJWI+jDY000UwegJT7pTCEFnbJQiDisfqmMyRiND04rDT+9c3LDKULYt
JB0RPU8FSE7O874BFf4JI3ByihS/PY0ROsI2PuhEy7I06jGb9343rsgzuw5mJfjV
Yhr7qc/Yr5RDdulKHteb2hwoZ1MGbrsSiwpvmWim8qUcM5sctYHfIpNcA5+5qVXT
M5JQSl53a7Xuhr8FxNoOVF9YYAmDYJJhd4AJ8dZ1qQm0IzTHJ7SS+xY4LFbQVNYD
iXAR2JLioeI6qHZHHeO6ffo1tD87bH0QI9gRkP4f+i+hZIWFpwXfbsx8KzC6+m+d
NOaMp6VaeGaNNysQdbBXVLZJJPuV2fuBjwqdo58zX8wVs5tZeDVAUEI4H3TSY5/7
0RO0dDjyeSIkgPb85Pa0mX/V0w2n3dgLGnhurOr0YP3NJfFvpSqm+GiVjzQf8TO1
bNAakNl5SLkX7M6kQu6pfqfkKwpfFhGTp5eu913SUHjPI0BhPYl12MKWlWmNvuVd
sV+ZzCzEHGFQYgzQFaBG+hOF9bo6SzHqN2BHX+FjJSJo6K3GjMAyEmkd3RdkBHl+
jui8/Hwf/LnJnjVEv1ZETRoJK/NE48dAGiOxrTiotHIJ3YO4P3/f91Ni/n9Esw8u
O7qbH5Fl1qaI4KH56Edpd0vGeyuyR/NavWxxpBBpIDbXnYptq+ap2K38PcnAT8N1
y4HYuPLjDiLZBAzdaPmDQf+g3EQqbBKurjeuEd6uQehjbzPEz6GYSkSH2Jbk1ZNs
h8JuGYr63ejSz9AfX8HYGu6HXTV13KPTD48eyqljzfNgHu7W5v9A395rLf7YvJ6n
rpNd4ZQUD5zZKqYMThYR4uIvASToUgEAV0nqbIm2yVarC2izQIwtTtzvoGZBrCIY
fe8f59cRRK58j/fCOW9iuvW+HDOtYFcKYfBIoToB4x3U8mFnBkUOKjqsOMLNnr2R
r1sVdeDp/9gGIOFcRWgI38IlQb/vpMqTDWiwUnN3t6N5sMT61VgPwobB0sYGLmHf
9ftu+Oi+3cl1kTIXReJ9VLl0Jl+dPX4ujEHp82Q+MVwOI7Rxy4HqOTriphL3ABEo
Qpkz94Yv20nDDaKIzRPmOm0t8/Ix46w0Ytiv8OHpdcs5f12ZO02QmJgZLTiANlDZ
sDOoElCxtzh7R73R2k3RmBqMocpsWtnjxlw/7NI94vMyelujm0lYiA/eSPhiH1G+
l0R1hWrp3VhwJ8Nbh0YRiUr6UU1qJd3BEEqLc4RikcGk4B1cxSrfs11Ebpq2xhEg
OIi0xza0PndTiflHdnkrKNq5jey8xt5U+6eunOseqsTUuNazMmTv2LPmG+l5oxEL
thR3pp540sc4jSQEs6ogJ0Y9LBbfJQUTptn9pWo60HsLg3DbpAor6v8D++excvyP
jWcafdsWW+EMKV7VXCCKt3ftf75eTkp1e3rmnuaP3jmDY5AXqqtyZFXxpwCLMCau
4zzkD/YYduI75oU4rOIuZJcOdJVv6LBRmFES5lfloy9HDcZv0b6F/Qe8t1OtTbNE
mp/xLM1mKuf5aMHxXA0va2IqcS9GVuYol7KGmLXkfVJgE4GUVVyn3gONrR5CSjAz
xB9rK+KUDQ5//8CTLUYKjT3zojwPBRRDzeGiiUFVQbp6eu6Q+M2CFfZdt3XpbOGi
Fs5QoCHgpLUtriKdmE+JSiyINo+9AX2jCOEyKl4J8W4rhjl2dH1XdBBn9ST3PS6X
l9TkIqVn9glQ2AWQnHm873FyQEBORvlg5KgjuYdC2PEcB9Y4AszXXZj1cft+JcYH
pliO+E+fXdpd1q6oSwizkVYXfn5vXHg5rEUbDzkBSlbRFSeIYCk18h4ymbOzTrk0
/BaboTyWvcpyuZ2/FUvQgKtvssMjSKcVbe1VhCLbuRZMJsJkGXNAjEkXPOMkdPBQ
Pu69tV70PvfCDWTZ0U03h96ifi+IH1pIfAZsFK26+9LHvAn3wLX8q5bdE0OTT1pO
PkkzB7/BmTldK/W0bE0FpczfPb5oikUAUVhK8aOX9uMUCLETDsGcZ+Bstox3NSWY
dUZ+uary+zb7tWcysbT4lXM+Ix/XuBgX+tnUQo4xKQ6ZIjkNh1NpdtAqlvVBrLko
xGmOC0vCOwcID12Fi7ZdjhuNkUzR1PHuD6TolWnsU6YghrXWxGordMY8BR2vcuIE
+zy46TEY09yI/W1fJ3lssHZOXArbDz3Ky2Fa/MOGdgbh+JrLxnAAAoLnWFPEQzEW
U9rtJetV/uQF6/svDiUabnNKPB6xR6cHFtpAKQx1eh4y+Q4/mgRdc5fTJmrP0NBv
yGkdeTygpHxtpAlpaiCSpnk2RcSZ0/4b4zJBvjtinBzC2s1AHyktVfNrHr4ZCKOo
Zixmuo+yFsFgwZ1NDO0ByywPQc1o3IwgwtvfF7QNgcnmv/N7xtTAbZ/k/CCG9PlE
TW+i72gIMLWPpeSh6p94uDyH/PH6mWn6AtiMFMi83gd2u3pMsqqVOKMR6wiOhnuu
5bF1yxk+ITHDgEtmn53zzu4QHTiQpMcGzXCJsI7wtcYm2bJ32w1XaG1B0aXLwEc+
vBpgCLm4JkEqjU1kvU0ouOWa+3Bf2CW7hwbXWAWKoGqQPBWQ2BIgwClfUmehdPPd
d71QqPCbJjzU8uVXpfoA4Dt/m/dQWL0p7TaviwKdKHHUntm/aDYRG5+DDy9G9w+n
OZpeHuxaQexrcdG4bMkjqcANVJljf41brEyHIeM3nEjUpXB6TnNtipkh8rlYZr71
57rU8sjV2NDslMR/hYxFWJyL2CSuVs8ERsLdxHGWjffqp3k8bHWei42EAKfbT2xE
81ovEfI4rRDBk1TIvHx+qCU9/aPfMZgQIf5RxYNIH0oAYpFY0tutzeAGX4y6wbsa
Vp98zP/tEpZzgkv0TYUUrDNBHwzfMXM9dCllPSVROfTirtLQpX4YiRhcje60mnxB
FXQfpH8VeQeakcJS6WR1ZWOC/34TdAHpBnjRdYTGbBOYt24U/Es4n95zEZKeR4Jw
k3oU7dCskjpoPohYTCEo+td9r7Trc1m/5bdwVbKIORsGeJT9Aayns2Yd4YyuNp8y
0tZSaQYT2cDGgK4ldYJIEFn561cdecX+mjRhC0jjPWP8Rk/VK7SSmKd2aDkBOyFO
6AbHDYLXDGnuzXEiBWc9OIlNCzutl2jBKToyGSIKhLdu+TF11rs3vwU9dPLELYWr
6qvn1jw5/5qEZj6C7FHI0ZMFZKO35WUzbwT79T+xvsZkyhTJWmJkr5rrymr2L9YY
40PcdJAJyG0wHgvH7l1UQKIhfdltzgpDIYYOZNPlLZaXaamX5RZnTsslIbi9itLO
0NIE6I9pRnSJAyWVUL8VwozYP5SHoVUYEJhltm/Kt6/r/hUgTtoOP8cv1to4qREQ
SFUPaLXp/vMEr0wngQUntOAljVvutECiCQAzemsalcPt53b5ylL0PEVDBfqcOm00
Et1FymFxRKuGXsC9p4wo2tk0/1agU8U9AwGU1+i4M0r1revXut/d5rDxJUsSE9rF
5LkYDcdc3D1O8ZsgPXMUG8w4ot+rkTW2nRqI4WLW+eV1zuxKuC8fApnOrkw99K24
NXPw1cudIbLHNIedhB1djA6xHjzawgGgBZBlb/dpUdNhLlCouOaBcktlI5yZ8NCc
I93JeiRUcF/J0jQnAlSOpd8EYEL5FCDF0TOGUAbZVlqyV8TnncuOVEjwlwx2fF30
KX+ds1ADu/G3ABS4Jxv1k8WR8okwDbHjCY0OeYhZvpfnIZFyEJU6vQYp5CjO7cmm
317D7gK9NxeLgQX7DTLGK5XHH50E+WYaY/fHI0/95BWB4SCmYkBUdHlWuiJWvsbB
JNx5K6GZ/G7GsK4AxC4TlLlilhCaeNrUuonR+DO1dt44Oa7Cj7d5+6Qs5pwD2BSd
wIfCfklx97OCyjAtxGXR0rdXL7Qa8fQ7IXavXUD+jTdft8loiTGuuPjZFPZpFl3N
Xa7WP/FAHSRqO+lugHxjqh724rUPoR3+f1YR5cdAI+r1nTQXzalOf/MMUih3Mu1+
p0rZLW0oGCkMkzLIYY91u9UDxo1iKfAVY5bFNZPdaJx7dja40rOi9rEi4IP7OmLQ
GL6zfxTTFfzjAAOpLrw2a3I5E7X5lxzreCJAq+lG9EX20mgO8Ocj5P3uAPVBZD7I
sinU/qko4f7r96/9VPD5jhYRuOjh5nH7K4GcRncRyA0XOZvS/jU3vOsef/SX0gkk
wVniTS8Kuuvf7UF8APteDq9Gv9wPU+kR5ccQQbK5s+csJlOll66HPUxwk7BvoCAP
z/V0NMua+hJa2Vk4qCVY9Or6AWIMbvZPJX7eTNLEETc4D1xtKrFKKm1+pgcyZVt4
HZjMOraMEGg+qJHC4Pk9pdIU/HxdqqwKGTc6/LdYjN0xj6T01NlHD+6SWFoI2sIg
0FfE/GL7UQRr0h1CDsBEpDRIVHCcZYtU7xGikluCbPA/Sf2/WkXvD4/B+GWtAY4d
9ISZDJ6SMqWJwgJWZs2clhJ7tqQmQbaGrRQe47rxJg3mr1Q1z23gYk8KDd5ngy1A
w2m7HbJZ1Qi0zQzT9idl1t9hvQ0oHcwha7ywAq3rDJ+RXpFgs+SWbK1iZJ4YTAyK
MKT+hH2ZLd9l7nJ3/axCCBuZdGLizRHexvD5X+AHodb8k90AG1pQ1Sr8/ZiEfjBV
rM6M0eZdtHjKUhZjL/BaNquxg199W0kR4jq6MEyb8zff5AbsmHw9WkUrDXRB88wp
+IN9zid3QFyIhIehQ71I46AIwd6SvogqKFXkVoWo4BwUQjnmrdtH7gilJYLEhdv3
yj2JxLnxFDf+QAYoc3WOmPkxbwnkl0frIrsARYrf7p/NUSyonH/WI9E/xf3CLiAk
88+ynYteHxiUt6Mt0XnrdyQbhYaeReAyc59RRcL7yVN8b84AAHRZoEC9vaQ5lXSd
vgk80fDYuxuVxjbUv8ls70ebsMQmZhz8Ka1+i1b0rUmkjjgplEVlQ4n1S0mKCKjD
/mZHhD9iDbJF7YD+mgQa6gOiRRumNqdwFmrFhqJLyPalZW1ArSoz+RCRYBNwNYtw
OJGwxYOS5tG73NKqDVmnxjJD0/1yljnk5EQlmA9Ppx5XdF/+tS9x8R614fMa6GzH
DChsXmUaePXE4JysJ90AeHc/Brjf9uzyco7DMxB4XzPV/dGjJhFPHoN/j7Z71vNm
chWHmYlSbUQ/Gbf/5Ja5gHg1MoRSuGRBDsxYpqS9Xnzu9go0K7rYakHpl4l0gNXJ
rnrCnesMSDmoKM0hoF9xIxtpJHCNQ524m8f3Vn1Jh+aAxggIvceSAAsGOjTy7Rtt
xiAx1v9vo7VbOa+Ff8uKZz+6EEIXXYKNpNcFGTB0VWCVfNHpuqhVODEimXs9qca8
n1T2sRp0mmonrFbM4S99DWXigoVcgNFV7cEX4lIrhPDExi6FyClUvHs5sdw/GXBU
Q6j4Ul0ZMl7nvo72bVzMliT9ibcnWbDsrfecvGSHAQHvdilILhz4wiq+DU9zVofB
pMTEdIJ04nH9YWkL0Dy6rD1VlQsBWunSU7eDW5L9/HPg8lFrO/MUs35DY0IBuC5A
gDXmjtz9e2ioS0CzoajAIz18Gj4+zzRpbfhf3js8R1Zj7VH0HT1YIDPVeUVXfSgs
j9t0u92c4Cjvs/AbEd7UlIJHmPEdlMTwXwKMawzrejX0q8Y0pSMMnc23MIc2fu4r
+biAxjMEHgK12Ux+A9XvxlzheLzL8ivD6VQB0rLvzv20P/QCSJjFnbX6hKFaQUSW
IBLFPrsvKVqCl0ke+fX34CHS+ZZ44U5gTvU5Xjj/taNfHr3aMKp2qREY7kVfOh9v
fpG6BVMEEYmWma/Ktn7iC5lXENJ/5y94VCmpX8qv5C9lt2f08HG+3CSLrk+Uvv6O
F1//GVwajzxIQgYZJefkChBgWxtwuaQpvqa8uKT4fh19zH7wQNSS6oa1dt0ZZVyf
Vf6Cwt7ztgfQxqDqnYUIqJw0VVY3cJ98WSZphU+lFPcfZMF9e5Skt0t7Hdqoz2RU
92SGvLPoBEk3rAV2m16wOucptfG+4g7O3WIUSlz2cdlxduIuFZsoi5JTISFlVzl0
xBfYKqL5ly/k4NopvBT1iNi6Co15WpfuWchlnfx5v0zJkj12mOAUq3Adk2db6MKM
Gk7aP2Ko8gWT4q0ky9eAvGYP/6td1whIKU/PM4tZe4W/x50u9N7+dhc2svKH8RaV
oGXDo2MoMp6fq3qr6tVFeG8MypOBMbsuZRvxNtJ0/Ff0VoQLA8i4y1EhNbYiYCYB
z00WBcUSd1LWzNtIl9LPieMFPr5QRmTM7eXPr+QBO4dGdyM2+cXrpWGFM88Aw7MU
+YiwT5+DNEu9TPpLCqJOh4tVmc7yjY91I86Qm/qpudstoza/heEpm+QMUVUG7KJ4
Ns0N3Vp63HHI1ttm+u8fqm6+FhJYOoQB761MJOVt2HLUv4+Aw6x4SBQuIlBm47EC
ny4/Ocp6qWe/dV3xwLN81PoOrlBODgXD2wCXhqAWu3oHeShgQFL9MsQh6hqRB6Xs
CbhkT0KYl4YlOVTLGH1ZpF+s6wzBwimhkYZNXt4cSiib6maWdCthezqOT/ejEfDq
+9+oINtllVhhQQ2CZKc+kjnJ3c9mJ5Lt6iYUevBpN6chSqjTsupvphzHDJLZg6gK
fEeV8syK55G7RycS7cTws4T08smD1BICuNxBNnqnHiUYB/I6lUBT8Y4AEoiE1O+x
+ZFXQdREviTV3GxgLX3KUsUIxTmc3p3cWn2rEe5nVr/IBrmjs9DlZzElQNEoT14r
59wkLPDvAu9RVRu3oRGYRM3zofOErYP+Ql57apIzWXPq6jY6aJBiNpE7pFwbNTqn
2i7j9AGiDSfmMEderjOmooxkwRwlfNlMR18o9+vpponHmOx7FvbSZ9Hp+iRNDF1J
4PZLr++FyoTIRh5Ri3GTtNpPpPOPkLTVNEKpgIUN+M2wHO3JEgTl9Xv96VmU2qBV
tOrIjVD/J6+JFmfconq4AWMM/J0UF1ELbHWELdb5gQDIJHW2TFzDs1MpPr4H5NVh
4dUJusXAJZlfMiLKGk728ak20fzjtJcAkzoKdpiNkaMont5GVIpPIfTgMPEOJLJG
PfRT6eHP01ChUiPX1hx2xIOqCc0VsMbZC2ZaXu07lFgKb4xJD7G5+oV1zw/Ysoji
pTeZaVf/WKtfdEr6VUVAbddgVsgg14dee3wWiLaBIQLNsfUWO/ZGtv6kheHwpOuo
NMgP7EuDHUvSPqVenZmxjuBwSgC02BJ4Bn4Tty0V5cA0U+mxw7KTXWGrBmiUaT8s
sSOHLQpT/A08Ri51+Sx44zwpWTGTT3LYfYfrsOQ906OH9Layw1SgUgdmepHy6AYO
J9XtOs/8hg31DYPMX28g2pdxr+HP8MnXZmLcX4AXygQHDcokUX2h+FnO/kdaftfk
PSo1MDpgxF7oKdNdtU4EftmB4xFa7DVEYQMS89MLsK8xqJzvBLKgJ+klcxSdLGRh
E/phmzsj/xKBFUhxoMSZ+6OfKc1kILXF1Cy8WSA6gWC131hePRcOJWPyEmQoUuO3
gqZwDe+BzxuPbn+6YaiGRSBgSfnoHg6Ae2u52n63WT61oZjQ/slH2JC3Ov6QxnLZ
myyytpSwogQHqkcKc7bZsInREBUX81HXtxwWSb9WYoHs8eScdKJdcvzeWqo27SUD
81NkiWO9sUHx+pXgTCBx6JT9t6yb+EjpeX2xobeWOHmdMr6Ka+/+McXKecpoasYB
UQSB2ztzm48CFMyXc6LY1wDXlfld3IDuW1C1nG3pmbGbZJ3cDkJyqGIuNC1Wd1+A
q7CThFRN/X8NVgKuCbVvFgRPCZ7iLeYBPGrYp/AW3wzE+NYrJzkPta4kYp6PSczM
7c+zPD0tQAozwfJOQdz5kOjaYwr+jf7BWPd7Fi1jRGr2NBwy4mKdnbSIpZ5yAaom
8/uJN7ZwdvAZ3JYcg3/N3XTIRIqTiWAymk8jgfaQhAcAmbiPvqH8Xjtu87vpIS+3
wR/zECA8u8KgAced15U3JVc0QiCU6J+af8MwwbPGEUXrvHmBCIWECXY3AzrFWm1d
/0rTz1+htpTGkNZm5osFZGZUJGSFE50MA6v1NgLtDynlhPzHAWh9RXRFhLRSq/dh
RKFdX+Fh59oNkfkYDeXuKbGFRkYxWEEzUWPcBDr08kshMwNmISa57lT4PxahMe1s
Z8UkktEF9Ufr2nmwuGfabntdWv98EjVuaRyQskux1NMAAWNGLJ7Kd4nY8wXmzoHY
QxIcZw0UKJkwwACMDSlFzUdafw1WM9HguC4pUIBsGEgi1bEKcPuUZN9QVDOFYtkN
0yHAo2RBGXt/+eiCnd6s70kZ3Kc2jCNeixMixAlFpFEori5fRSkLAEwz7eEX+Yux
+uut3hPyyub1m9NnEOA21JTQMgxL2BXro/PKV4GCqqa+/7EW4Oz1j1HmJkfSIM5Y
+b9wqNIWxNY9aYM+eTEhY/3zDnSqAJ0dK5RVXdSr405yV7lE+yaEm7l5HyZTgZ1s
zXVkRRGNyHSzwh+xrmETg+k2aMMD4NJWlSt6yM40JwkTwtC/E6b2AonbtkISzZYQ
s9ly53vfi/oOI4jy19QAljBdZwOSrgSlDB9wsEFaw0FWdtiAu6oTkU8ObmIOCnkw
368LQ5yP/eml9qvxcZT2SJKqsWbJ5997ae2Z7ItgSQI6CxZgrirJAmIQUE328RxC
1+CYdF3m4z7nbh9lRaBMKxqWtpVfhCPD4vZ8c0+7XRC04FJp5kLW8O89rh6QBoU6
wcMuSR2SJpDbVK+4EqkktWzAuT2fK8UWsin0wbmY4AkjIj+NxCZaslWFf5ugCBS4
gpWpw1B1IVzd43Eo4MC29RBrNtADsBJ40AM97LAA+OmyQoDoDf9WPnvQKgc7m8HB
jwHKbnKj77lFrwApdS7AP9VLvR0aB4yUkmPTfCntRFca+CEHioVWGqAnrbU8ZIpi
sbkjPH6oLM4WfJANh40SsaY8pH7JoPjqk+syu4SY/p+/3vEgJZAzIfSSPH7wVMn2
huW/IAjuGRIglghrQNeNbGlscy8G5yJBAHSSXRNJAfo4GCTKa3xa8PRaOF0yUJnI
nwXoucLhm4DZa4rzIZYUZN826jh8jjoZiRCmUJympf+MpNhgL0o/amHkt5NhaVFb
KwruyW55DZV7Ossr2o1g4T8YzdPbtB1teu2Cs0dJU0mocroBXFc5fiKuW/pgAj1S
0A/Ip4RHG6RV3glWHmVIiYfrsLeCC08Xmwrvx/kT0xx+n3JOiGPPltwq5aOhJ8yU
WZN4zrcxzhZX89/5/IPwU2d+0/LWw53m2rejD/fzu6QEeYXcOXQzjTHy/oBDkvqM
FCOXDi2J858Dc0jcEnNLmnSViOmuY5pY7tC8q/x/y+8W8bAmNifX6+uBSkqLYqCe
7fYRRnoe8Zb3SW1BOG3Px2MxncWtmlVYZyogF3oIi6B0mw2yvDxhAjMx9+to26x1
OFxMd6g9+oRuyta9lo2ii3m037wmqoW4G+Z3y2IvOagP1p2rv+iWQG3l3AED1O5k
cAQ13G3Okjnl0yOE2jXL8klkzswdqi3pkap00vv13zsvwTzCjf/eMEWAlHF0T5H6
RCLZVW+f75mjIquPKS5ywWVBpA9/GC31gHY+2ijueZGxd3lzlxyQtX1Yh+JJhlMJ
Epw62+SOWFDpdMgDqEHYek6iwEqNCU7rn5es+Kjq6iOmgPgtJ2sgboKE7VyDfbsc
ir5d9OBYYZdSEhldchSlFYDzWndQvzrnZQICVCHsKp32XN9V9khHsOJxpTqngCSC
qmKAfzEItw67SHNYp4HW1H51JgJ5zmW1XiAW07ifw05GioFVEPD4faY5DOjxBPuD
Wh5dy5lAKoUl8OLZtRtOJ4D486MYizEEQwAkfT9zRulXANz3RlxOLAaxLEC8UxTG
4hpT3jfuaOmCBs5N+FYAlnsVts1e1rQOBk7DEDI6YwvlovkQk4ysRf4ctBoU/2Dy
y8ZRhYqOsc5QQdO12LBA/aPOJpHysZbm4R0yMSr767PuMy7y6aIzpERFONF37mwk
x7+mVmUXWleVLTorC9/ThJuFzZwVvHeVgGLEuOe5fRZqHR0P+J01YvKu+fAR8tW0
+9htjXqj/ZKI9bHBDGSrdcb8EGin0fub1YqNvkkdz4tAyJbPG1oI0ujyJlVIttAg
DyNBg8xdNr/SNMz3GKJU72KH5ryFaW1lOlPgb3/khdGx48CtPN9r8PvRv8C4WjDm
lq4/B4CQVba+SML9LCyN/DmxAmBVxsgzbZkT40YH+bGqTmK2l5Nuj0DNWNc5V9DV
koK2YKdE7QZrMIJj/ze4YFQoXgu7+ZgHqf0PGhIifY+zIHBFf+PEesGWOGLHqkQX
Y0aptwh3LtjPxW8jrlstSvYc2XP1rIBnHm8foVxC0I+4K+DLumzb+7T/Q85TQ9rO
PxS47oq8GUNagl9OfwBI4b25xa/gvCNEHagJl6017PWJ6NwjuIFYij1rFgiAZ5n6
xqtJRuhN0YzhonNbOm7xqZ3Rlww9jjiqa4eNV8nYeBBFcKQf85aYRtWirlQBSsp3
0Izk8lknvhF6rK1YkapqmaYh0W2Nta65w9nlyqOqhf2SB2QiBR9e+WXnbLZfPzVW
hgaIKNX3mBMqODyfhClj/7Dyik52UPn5INLgK9YZb6xH3rSbpPu+GiduzGfWgBpZ
ZnYUK81Q0Yym0ZbtMVcrnM6IYgf9bjIbiwdzLq8n2+vbO9k4Eq/4SQa3RgaXDoHf
bP9sQRxn8gKDLKPOjcJOGLrCgcolK+3etOAR+ALStZjyXpBK3yQMA4V0fNShBWYJ
Wsg90nw4Yzm4vLRKvJlZpDiFwpU+Sg1uzOd3hCNkJ8k33drVaY7H01e6koj4f9Tv
WRPZMAXsmQV8jCi0V5ouw3nOeW58JhkKIwcYshIJ19C/FxKG6uUi0DC+l7BU9JWj
P6bSnr7V17YKmqePxfqkWIZIzPVoUB2WXIqGMwA/yFWQF8Gjw9/7veSoK/dwxHjS
FtB0NmGoYFlxi+bV1jmnt/xOX0ftok04mIvP83Z8h9yJUBykpBqZjgQtYNZms8+0
HYZJ8ip+vrLGoPr/Uy8RJinNU0zeKXrZlFSErx5DXNHRrWLyPc4/V7uGRaRLu7hh
taelk4JN0jfEtpcSpRycO6JO79zaDn9h9kCzfLqs7Xeph8ls3mJXzzaBgc7xFw25
Xf0cyaUasMBGDHVQwLuGjxa9hXr+lMtj7Nmiqj/RT5z8gljvHHlywGfZjgwyTeL5
iwxUnkmSGaPFDbqaTNuuPTttBNY/ORzNGPNKOvLp3El20Io9asLq4rx7AXV0+seE
GYD/8IOvPp0U1vYKR30R9HkWYuCfu+Ps64t4uXpwsGpvtSI+hejXJ4YbQlH+yVbR
jlBuVW1t+3uuIrz3/Xwazh3Ibajsb1ClEiQuz+nynPERnB2IRDLd7KSsHGZ5nblu
rQVdMmPY6iuSo3QcdTBBfH7YTF5Oopo+eCCUoMkx/riE27P2jF0rlJocS22gn0Ua
j+r1WY8SXe3Ew8l3qmrKEtUJiZ6tZ/zVZCWx5BwtES19vEl81HEy/D3MbrZtm//x
SMJBZ2ZLHObQBuOTuLQUSsLz3DxQr8LE1JqA2BRknfS3Gqgg/Gv/YK5BOiWboL9+
gfurwz0uKLYf83/HU4GVagOAPDY9Ij2Y1T/ySF7ttUtq1YvQShoSHb1GN+GXx4Bp
1I2r+bSEgJcvG6Y84PrZ9rURlcGjRLk6TPHNkQcft4vBJDR37tbx24qqtqoE/H+I
lMfHcw009IfKZlYOijEqAA7D1tlaBDJ2NyUxAZQi7ua5NpjGtAlbkd+uqdJBzpE4
TNMmyY+a10Aq1xU5j/ZMIZPxo8PXpWZHUiDFV6HOZlRwoMDhntvk7ORzqD0OCcgw
Tm/IHNg4DcCEH3zeGYIYg1O7WTu8JTJDglLEWoefdhwhSWFBgn+bXbTCH2sfMXuK
JYbSfiqZhwAsORjT5GFqgPxTzVR23T4gmnj5SxVBD+REa8bmzTAHlpwHJPOWuHaf
K0/YSBP60ZSBbJgp4IITIoii9tibHzktO7uAID7Zh+8WIa75Vy/yeqS8mE5GB+Pg
s/yv4mfEMRLvTVtZGrYa/vxcYfP/jBROjt8nxjMyvk8iERHuJW9d/PzurrIcE6jH
AB3qG6/6wWhzSUCeA0ohvXXigwdBk9xwQ519f58E6VM9O/EyKDWxxd/tzLGfQoxM
skmOC89JdXLjMBQAo5HiApcwlcuMijisgbLwSZTTAYZdg0vweUBf0iD5Q39buMvQ
FLYP30zSX2ROtIbhwBsZ5HHDdQRhpLKlK6VGFXMy6zAKPSZy5lk0I900oUhJcMIG
Yg5STrqNarB1EQMXbosDBzDu1We5DPeox7CqA05zJOjNhDqJUU/G6KOneA1ilwjS
uO/g4jaudHE5IVayxKE8uHU0Qlx8RRi2ufSBXCBNobCK0eWfewcOxe+n4bKE1umG
u85OTkVr7qI+K97vAoNrt917+bHJOtmt+mOnUuxSnbaSkMENBLc+vK4vAWjSav3y
/BtEnZvYuLVUXOgUWo9SeA+wL6l3/eDVEp/CUsomT8WjqpSGL9Bz3j444IRAl5oH
BEQYV7EdmQ9pYpGu42Kl5h8m5wnf04C7VMdmK2+RR+HIXFI+M5oDeVv1oHbjdbju
sjMiE3o50yfzeALqS2FRTNzrMdD3t4QwuchZ+FzbQ7bTaQAqwmBhc8qLySSj5Hm9
1vLQjp4Qi7zStawRJ4L8a1yAVtboVUubIciAxyYL4oBaFSpps+sHqlzPtBAxy1j3
sBhV65+90ww1yM0JuY6aeMWTNBbcSlMU9EDlltN7x1HD4NZv9wSUe5xAm6VVg9ZT
9PebdG6mjbJ3zwEjYQ2JWJoc9BaNwvpOc44Ft1vF5v4s34ws3qe7ujsH9OLS4akx
ji5phewCrL/X9otlq4nSV4AFyAXFxD9WBvggnD5IU18fW9C7Cuu1t+ltSI1VIerj
Ms/9WR0jPiXygVAcrFmp1vMlGtBphayLre46oujAwNz/xvA/74pkxjiR4knZJfqt
K+Blvdtzjj5PsUzcCHyQ1uoevosOr3dNx7zoBp6aMTGZV1a9P7cIYekIAX2YlHYH
zGUYmw6ul7uCLQjzbQwi77LrH1Qk9cbWDIlIeYZHjjTQcVyUQUKQpY1gR/SjjlQ4
38QlIunmes12jR0gKur8r8OTKJZS/198WqzLwAS/4vgV2/5m907edsYO9+1FgoS7
rqG6nx+C2E4CBAhrgRQ0E4poW+Txrj1zzbzB8a8VsGwEO/VE5s9w3LKxDupXKeHE
BCgAmnwTKeNJiC15eqGYTmTlIr8onhHidyMLWCc7LtAoi4+Xg8JziC3x6jhvXjOR
zGuuvzsJZLzUanfdJSvaDcfDQPu6bVZRho2MVb1EfksNhMgzi70EYhZQGfY8kPuq
U/Rq3FRLFeMEruE8IxCLEmhcFWgmuzMbqLD6TW3w0GdTkpD7X8BHaOcbaViQmETY
gGEUYHZOcEbDVinzOtD9vNlKt3839x5p8V6XCidz9QqLZ5Y5MuKyz4ykFkgD7vW8
mcPbP9IheafbPUdTz7+/8yYgDFItvECM/sb0ulIZUrMHvfmXK3mjGQA6gl03BJKU
cMz1g4tlB8JhUT3P6YKLDXaAGdIlTceNv739JNVwCSSXSqOeBxEUGi8B6YaDjl9A
PjZvgxwz5N1B+v6/mbivQhUIM7S9EtBDN5U/tRF8QPHPg2D7gM73ne0JuscimvtW
TglJhhOgLmyVCV9sNKPcuwrPe+0L/csRQYmqihIENV+c2brMIS5rB4+E6s7+DVah
84R6O9Vu5MupvCEJ7Po7wxDg6m/fSjC+tJ/IEA+uE6rOKzf4UpYmLiyM80dCBWAm
BOmNflEkWdc2YmB3YR3QtSrnBLsCFwJS1W5OXAdMgQWe0eckZO+4Zh9iWbKD1b5+
AoaTGuh5zRafEGUJeZIJLgULx4lR/CMKkJQBF6mghDLtmcUjR04x8sJk74P6zYcx
Tyl6GY70Mj8FXZseWaFygUenbkf2pDgVe0U5+g+DDCq/HcPd96dJ239as4QxsbFS
rWywUkuHPKXjk1LrO8GQzFoHhLFq5KGhXYXCM/FXbc6CdWkVfF1ROox5rj4DfneN
HDVUVSA6z5qc+5BElRmlyNHBRPTDENsQDgKOE2qcL9Q/DeLpfh/1C+vK4nh562SU
DjrRz+vFuIsYc9Y31wzyFZWLF4vvIc2IyzxXm0ajkHSoxynqvFldDKDA7JI1dkF5
QL64FvPsZsaa71Gft8oYx7pCgak/mUVdUDbKlAsvPkNxn0/f6buwv1QbPcJX6czl
nlbglpjXFtqLeer6KyqB7ojqCXmmMunw2zpy7Tn9CXglbaSEztAdfoXTw6rk5IyE
Wuqjxd8yAE9PB6G+QfUxngjzXXC8bx1qMqdHDoBASkffHMBIgXRgoIt5q4exgvWZ
bUisXQ2H2fJ5w7GT6h7mQFb2Y5YlxaMTmAeN8qAmkeEB21NMbX1SjN1gx3NOong4
S9EnxHOFBwzjSMyCrIR95tFKnYIELG5T69YDckHQ0aQJ8JQEPD9K9KQq0mN6/+uf
XJmlO3lSi1ThCJABEpvct79xKkGD3oyDKJMkS2xA/RmieQgBgXrAN6rtTWsuLNtJ
ObCisVF6dlbSJuWk81RHr1DzAcryHWXrLGCs1evZ/FQjsTmB2HCYcVP/bjH1ZtmZ
HQpevcB2BOKJLul4Zcf8Bb9t6p/TqcW4POjmfcgADqDxv4cva00yQy2je9JWVvxD
zXeKORaiPFleWWVGPRvbUZNLzAFTL3wH89bJOlhYAlKiuecm2El+Wn1mzcuRCMWw
NvJOMn53gr3JHzDadpzkQgYswUQT9sM2LeZlJbuk48Tvlp9KqI//IRwGQ2ukR3Xg
NA7ZipBK8PCRkNAHEgk6e+il8Z7Sl6Kszgga36qk1vHHS6dG0OjqU23HCvcD9D80
x5XtL2LDIo2a91++Vc/Jk3EYl0Uf+kSPmNWXuAWHuZAIgSTVFAaMGX9UhtUYgeEF
CwamFYyx15BoBFrWhfSm7uzDtZCThiUI5v+qWo7DW9COXPagrvY7g2Jqe7KZuZMR
wcm4Lq7JY6nCniV3hs6I2S1dYst/DcRlhs5gObdAVy5BeWXiPeIv/hgEKyeW/oTU
XxY3t2JQuhv4Igasv5elPX5n1rYPkmI1C7T7i+4Aa/ea+VLkPsTzxS9YIzIymin2
XAwJA5U0PSPOp3+cuCmPPdVbWLKXt2osG7Xe2W5y9YrkjmsbvkHgkM8WPqhp2Np5
ME+9q4QnqFivoeTgHHgm09yXbFlLCR4kkP2qnj4St5qt/OzlK4g9pZfkwERkBndy
r00ghvKaoKl3irT93MgCPCtmCkQeyQUSRQMPnEhfWKTOAjMjsSZeUk5cfAtKrret
HVB9I4q+egldZfPuQseX/UIzqIHityrh2sDAmDFU5SYdz7Szzs6srYrM6wkaNBxM
lW6ApPM0XyIdC7Sa5XdwpOzzYqIvzodedr3vlard19PhhVOx4Azzk85m+wfM6NQn
I84gfRm/Id7Ga+Cxe7okyjUkoITqMnoUYWV6BCuhUO/vPnEmP0LmmHeUicg0k+2A
MrT2OVMxi0O4iDaUUZ8QqU01Ni6/f2k7KXuXK/2npayUeFFhQGBY0mirGA0PfL7e
hx8ReBf/ZRzhDi3L15PQjEoTqwQbAFXM6yaX/V3iN8CwYQLRKQglVG0t9OcZ215X
W5vOp3Pw8r4Y6FYGT2e/yOK5yFW/zjRYvjKUCY3l1mRPH6PLbRpX8H+LFUOt6Ssn
LbKHncuy4H/J+P+B6ocJpASUJ0v04VFvhP6UOqSOWjrSbWCDXeLs+YQFk0tPF3Hu
pVpZrKMaClFZ46bGZFp4aNBhLy82RFQo7K0yrZh92XSMAz7K2v7cvLLIDI1iWLwt
W3eCVJBGcmzBsz5LNy3zQgKPptKNTMp4V7Q2ge0pS9tF+I5q5MMx2bcIyp4KvlvQ
ir4+4a2A9OhwS33k+TqGZ9uwR77qZ10wWrPNF5XnYkjoPLfYfe+tiSbHUeIUUvSZ
EakDFxI8GOcRagcybQO5iVCyxzWUs9zcrsWlpnt+XGe2elo25Z2dKoK1qjR3dP3K
3AUeP4vBdid/j/jBtSZagRAk8GxXppfZi8wps5NI+dIBxGhqnP/oUuGMcvutjJAx
+HSHRwkIgNZ8bsEdxjk7B1f4ZwQ+xMyX5k3rzgz33AQHU5ckDHtIrZT27P6H/cUY
cerYvxyTLai0vyJn0eT4fqkwTVZONgS5Hjr/z+Pn4kE1LwnVN86bvJewxxMdvMyg
cFMSK9R0CNOCeb5haW1qL1kQ6BJISCAfirEH1jlUof1AyKyj04VcSVHvPlFCkD+J
vtaKqiux15aeVd+zRDAR9p20i85udkA7g9qyuXNXzrBK5sKW3jaDH9n6dLrx74S2
fzxBwqBLZJR5nQTG4OoHJ/IDJUulklpKCG0feC0kK3OBVlwc5gGVVbMkltbRmbg+
P0aBhbyoT0Ghg+i/z6bBh1g5MBavdEliyEH5DY6fNxk+cTF3I/1DFESCSRB0g+Si
7ayN/DlP9UCo0joAP/GLbTjM6ms7lBdFDYUrH1qxTiY4HAHbF4mgoX0bbKHiP7YM
DOdf9KtVrpDqY/ZQT6YOYdxli0NtpapyMciAyhVq4vnCLpkuLnDbdnOWoXJrecvK
cUQhtEjFFfKQvY09KutZvlqXRcLXU1DEVtsSVVb4u444a5vVK2PjHTnW1nCR5eqt
36az/jy5JrepmZb3oNjKK14KUTEUV2NJ0rEJuABfve7kWwMTGKtMl4sjM1OSJZCA
0J+ak8YR8TBel0xLnoUMDZH47CL61/t77HCl0zdLV8vwAxnDcwsBlFbaZUiO92kr
xgOCKSbnuJjAazcY+c+Ua/FKFzE5IPSAMT3/z5IEVkcwmDBxlhZBBGPqE9MFRnam
h4tW9jXO0AkXQRYzdoJcbarJTW9ykf0McLSkXIqW8ncfvcrNeZBT7Tzw8m5N5ixn
T4QQSZzFIemQ6aM0tyZbtH0lo0p2P7AtH7okC8plGqTFpCiUe8n7qh4wRtxhSKWE
LhQr0Wc1GJa1EmN5IrfRrW7vK4HHscyEttBP0RxVC1Fbg8ju3IbyuGWOL/JdVFBj
lUjF5Sb0cMuvWLTHwiI5BoZmLcNy2YW7YVXdZ0+r68zRo0zfQjx89eV7O83351Iu
n05S3UBQZf67nDD02Sm+Jn4+W/FVoKSJnVK/+opSjrhL9xt2srqajk6/g4OqbXJ8
3qdWVt/nwvdPUbGIpHgNrnYB8nQg2UAvWx8SiKVBlqrwo0yzbN4xjkze4CCLpRue
p8EUr/UYkpao6b06YEwfseYLAeM8koLion7qHHgAVxtOWHXvwfgFqy8jfUWgYrOM
gvAaCrZut4L+jnI/x6/ZWcgA1h4l6l3byK7uRXqMLQAlzSbAQpnVhfhtjv/Vloik
xekr7GXbSLgYsRIPR6AR4xghobYEnpv9nO/e/iHRba3KtC9iOh2vtKUXWTb41VSs
sLHch+K1hkNZhhbeb5NISfKU+paBLrEdXrkBCNUZlwgd0mLltHjfvvNckKXmC/7T
iZdrOYOQUW+3lfbhLyQOV7s7leUBQABzvg6r+I43QMaFLoOqO5Z2VZ1RWjwXNcKy
71tVRAzg70k6MiIY0DkbRVE/bNqz3SSSxRptqfiFLfX3SyObt/ZfNU0IddQnA3R6
36n5sjDI8uMflT1J0ke2NHhxuG+5RdnRlKSrfjsFiAiUUXb9BnRFAEP9LSMCTC8g
/j+t0TPIzdGvxpemVN8qcm/YZ7EwJC1IGwsVDg1OV1o/mbZrsM9b0RDFTQn6aDKp
f0VUXXqPa6fppJEtlvGEGIpaC+7SVSfKbAoagWEZKEeJ6Ya80g5yPHg9TsC7Dv2K
CnTsEc7PJyd7ye46nUo18V3FsvTzOBN3XFG16BX+aLbj3Rn4pk06OL4oiqI7PnbZ
FlmmJ7ijY0JAbtI6oRHtqUvdwFkPaXsp7dPQcXe2HQHlfTfvuF6Sx4X5YsXlhe44
8y7xeDo2ZTLIASwy6PkbvSSDU2iGhTn9GnyHmHY+mM4H6v1NiYwHhVLz/3OjoYiM
+kT7DmV9jt7pWxloWVlFQHHIw9QcUeGNE+2WCUMv97wzZhHQ0Gu+g+F7YCYC6lSz
wqyuAXUNlVaF9FK5ep7zahIVLHNSAgUXPnfBw9xQdY5ay4sowaHYxA5hle1ZkCy2
UP9l3P3KHurDjbRkRqmYXP/+xMToDf+n6CbCUN9UGoTsKJx6otsy8F0T7ERXmXGl
H7XOEgi52Y1SVAC8sCp4FjQeHFCy6UYVym7iXQfWz8fy4/JlKS750dlytYEY/4T2
SoJeElSiXebM00ZdW5/kBYpUkWJAqpxlvXOTPQ+effEnzfCyM8FMB6kHBBZEI44e
dtZo52BwYQ2O2RgAbU/eHWZGiS3Dr4XgKTFf5pjp3tLGC//4ppxYyTDfpH1g9iNM
RKw6k27qzKFlNh4oeRvKytGHc/tfWbJhU7ZjkdJN1aL7JM5MzTD8tGZqcAs8HmF3
ox4Kgn3DMXnPQ8pfv5V5Rta6JFxpgiDA70cvZGlblknEF8SYER4qbkjm5PM2N7Xz
Cmw0Y4RPuGFsHdXqYfsWzbPSt2hnH/BZLwSK3my4qdQMREe3j+6+cj6Syv05scSB
+03zmeoiJ7LdqMLflFBatwkM8KzO3I0MXeM0De/z++Y5F0TgCU7tfsshwJns/I3p
0A58S1qBttYBoNtLLteg88j989hhJUDv9NqvdZvf4QUqxC7gB3gVXeMuwssmDj6J
sZ8V0y3PuPFMnaIYtZ+BwaqPX4O+p1ZcIhWeTaCgzrbIz3wJeLQW1h4uWm955SB6
1kg8KKkYiLedw/e3OChg3MeljADdi4/t7G0oVlrexA+OoPzm2AOe8W0rD/HcfATh
040h2h7AWagmGxJRw3BNljFwCreBCwoBJsHlVWBrbPh0aR9Zs9/1aEp+OAo6ELBF
bLVzWC1PhVOIPwG7azcNsPugCIR0gy0KK6PFhbzrHHpEjUQgbuhrAK7col4qiP6X
aXFdhjWJ78kKqvf05r1kInytDXG1mAfn5Nub94hcW1TOKjC5sLeuIo/lEfWxNIy3
2TfTxK+GORiMz41Mo6zcDxfhTrD+GljnDAaov0trY6isDfMB1U3h5JnMAiQe1kbP
uiBRVorEqebvGU1LxmhQoZGX4QLWD4oBbFYM1/akkvqhnVaXB5QwGeNieAI3dWWG
xk14KNR3yxI4jANxOevj+tdCRZZj0FRHMyek0WCgUY9uZ+mafekR+2IZ6lcfIhog
bDxAjaTbPaMtU5cbvy5G335c/ksuY6/8iEYtVVFCwkTSyZ0tLBhuQzLZjiWHiXrE
T3SNuhUyuxlloXsRvuE/3Ij5F6AEe4cxv6kYeX/exPpTeO1nwraeFowUrN6rz130
A6XB1vKJslBT07BLtsu3CdeeA14xyv+IFMsSWQb0lEpzKUgAr7jq/CUOeX24Ctu1
/rtAy/7rEsoGx4c8sgcdzuaNFdiDk32A+uESbZkuJLJ/xE6eNMKdGKDcRmOgI39o
Hwk5Gq+VDLPqPGPuHaLrjhh49FdgKNDFRz5KHXs64pd3n22DnRATyzcxS/ZHmedF
4NeuRVGGY3aI4HIOIE6ho+lNJbfDS7SfQ8a7gbrck0vdFENaqE5+y0Oo8tgt/a5s
d4rs0nmOYu771a1P2I79ZPd/ShdUlDYxcl6Cd7skGZu6JmtEpxLgJgDADU6irxMP
RyO3hg+gw/A05kC0//F4dGwJiISlsXEAMYPVp4oOnB6Rd7z0svbaWkiiduZI+NTl
Zo//7BHS6iJ/RUgKR8ITVBok3b2iMj/lUGyfNciCg7xrBW8lAMJr0s1IdgoDnizx
rcOrg4o1nGCVrTbHzp1X/C7d/lpTqRuSOXkn20EiIfzEX9RP0TJEvv+0Xqw6N86d
VLl8orSH24Ue47r3T7tywEt1mIbQXfLtMgtxYD2KtYgTWpRx9nDdWw81ncHPwQ8I
01p9crnUrj0f1lg1y9CmjPikrwYJ0iY7bl9D/vo31v8cbJermG6EZodX/I5Q1/rX
qrL2FfF+gfmhYz8oVXFgm6xBbhu0mM9wTp/WedkAsgRcDIvrnrFOVARDJaCYfyXh
71LnyxRJbJSR4kIEfNN4tfqVDKLK+RqGX8JropERrfWQG46ALMDsD5ZlQKbBj4NN
P4vs5s56mDpqNOtacVFHojKqT7zZSX/llufY8DUyDjEuCyovqNAzhE5hn/1f+JRI
S/Ekwqgp/Owd9wb3RkiTJIdn19vjX+Z8LtT+lTq6BmxKFy9e3BX+GzAQ9oYz1E7a
oj2Ic8EIFBclL45wY/KfMfrwtOhx0wJ5W++8XJGgBKEq63FXnUyjbQIXr0C0A5xy
DK8iuN/LUxqpk5ytvAy8WKWkGAS6ZrqrV7DxEYfmSNSbJtXZzc4P4cvi5STNwHry
qMoh49eV9jrxDI7R5T8MUogqpdfAz/IYx9IP4fV4nFJslFFzZ/+lW/a+tXEdwLKb
Sbdc0hRonJdO59m5M8O4MIDE4XaQaWrMhuaxm2tkSCp8JzwjvSYrKKd2AZTb+dlz
VShMCFLBkj+PRSphez9m2ThpGzht3aL2JN2lLS+Ed7j8hv36N4nIDRGxt7MhlLaO
YsEaOb6da8yPl6lqdDkGTyIb3CRSzhKmGuzV+6Ch6hkbWDVpq0J85h86kTOs2Vyo
bShEtvwMIJDJa20RHSuV9NUV84hgkVan/crstijBgYB0gvx70tm3OHtGFXrw9wuu
BTdOTXvhyqrGj3xWE2l9e1Ea28B2N2kOQGIinSKphIJSaWrf6Twgmxvlp2eI++u9
WQdMrboELvSfsuCH3Mj/E6GIFbLP6KxzY+zOO//xMyAUVtlpRcNL1I24rhoRyf3K
Gzf8My4/fQbfcuC+8VRmfFjWxp+Bm6vzTY9Fe077nbOHAiDLMRW0H0HsbPS/yb+F
bp1u9xnI+0qzOlM4QUipXwP5r7Ettyh+2880YYlA7HCF7mwpJ6uRaL3s6DMNZrv8
x8Vu7d5ctDZOWJLk6sVxxODtdhHDoqL2P/FIDnauGsbE9LGLZ8FC3pbdse2Cl9l5
+MtCBrn1Yc3UWT4SfiOePizoWnGyps1b/jnOjcu+YhIOwtTLuzutf2ZAod9UwLRE
3S6oyH9sPzdma4c7lV8Ch5mN1K2+AYuN7/T5nYGgHHyVGlxLdn76oD6WqAUt5eQx
Mh+8Kc4x3PVEnX7UbxbV1lz0RdMyWfbyyyJNi+SlIRhZ4oki6o9eBvDqpWWVnEF6
wqL9hO86/Hy5FQhtR42GCXYuiDq+l3ruprmgtmrUj3Tjsy3dZeJJratiz6HMxz/O
qjPzxXVAfWCv2en9eq0nI07grcwuEpzKLQOrtDL3s1hTF3yUnAhHgjtEh6ty1pbn
z9yxXP7JQJTPJnpbRkrbtB0TOIat9gyANkjIVgKMBIOfFfha5vE0IX01VEtBcISc
ZLbzFfgajr6BvE3R+bCky5hZUXEYGvd2AYs/BwOWUJ9npBsMUQIyK3STy9+I34OF
twWCtYmLMWaYBcLdXmyGPfUGbQsC8F3sgC47g+jJ1nYVZNFT92l260Bk8+Rk8sIw
8ohPOGQHG9Ih+YowFUq2lDwlVy56DALieDilJvGyGd+5RKPdmEvpdZUyvQuIW8KW
wJLu/4tBceAyfdKLuwL/FUm7F3LAM4orpH5vZ5hlIuNt9td9r38cHdjg4nUgb2i7
38rXBhaHVfGT4wGVYrdxdtVE69lTNHBM7MIAQ/oCPUd2MVlUJi1mIWsxREOdyjJz
2lR7j/ULFb0XDATEbb8yt0FwVkBwUkEUzpTmdQMVJ/Nark1dforXbS64Z9cNbhpO
5Cu2p3uSx8SJXt/L/7J9pREM6KPhrB3xOycBY/BpUFbpBk7oj1+BlSy9JFET259K
/PJu2De8NmKrmmzmqUQdaw+JsnYX8Qtx97BtfCc9iukq8Bpt9c7/o4fMfTsMkydA
hK4t2Z0M9ozKyCaifOdAmc5gOvIalSZvAafdj9TpZkcrxJxbigbHq2/i+7YJEwGb
psb0mOatIflzmbkt7T0twG75Bp/8r1Umt6iW1/B247f36r5Fnyo/2eCmk8+Hgn4z
ycza/aZZ1dpB555ynJmw1R7eDaRw1lr5lFbJuzzUWxuwebcLERo6EcOKWud1Hry9
xxkf2l+orGJrTstkueugt9nmI+a7+wMSCdne7xbZug0Ll7F+zZFrBxUV5Kr5INNd
1XaOziFY/aucAE+Pi+LMQ1yX4MggLynxzbbzOU5UyaY94ZZMwYhknS9OD//124oj
Fxdk7wPzKHJ+456oDJ5h8HnXK0yrsZHZxc1BbwG7+2cpAALdZTLqseN0QuTnOD9+
DzOa12Vm3MYhzV1/6tCPpfjpgy7kNLlHfnU4yCuMc6TOudyerAnbmDUmixsJaPy6
5uwXAf/N8LEWcX2c+AB9ht66LeU9v5atpcodSqPWX4IJGpNJZZfSL3cfS0YWEJUr
kzb7Sb2sJ6go2pP8wXAwmMxIW/0oYlIw3YRjfl9DUVwcCu5qzipvZXXebdD4H70J
mzSMRpPtBWMAbCWEVHTo76oj39cOA4PvalOb8kJT42dZJ0kSBTS/1FpzWD24FD+W
r44Pb4/W1zS4uzsQ39bCHL4NY2gru5U+j3/laHopI3dWKAAThHXBqC6vitZmWcDT
l0ZaHNTVxUnYIyZyO3quZf81axFRuUiwGP7P5VctS5x/K3+/DeRmZjjsTNl6UJva
SLZN+OhD2F9aCdqqjTMJQ/T0NdQmim2alSLcCMrb+4FqChk1IQTgbY98tLVumMKs
ehH8sxwBrP97hUtadT/KaaATOWtVPV4G+TTwKwq1TvO/52a19GhS0FY/R6m13Blk
pnGnWqgUGBZWV75pHvsPN6WqCRNncy74a+KO9Bl2G7dWEJOt+OBN4RSqOHaOmo/h
8SFrXLS5X5tcTyrGG441Jc2T53DvkMDdyK0hkO9/CHLmRAauxLKPLaZko39hVgAQ
FemEtwEP5pcOfaLk2+5aleCgkpvEy2Rpg44aQ0y/0/QzrpZcuor18Z+sUIofIiqu
qFPkce2gCLEcSW7a/zbCGb+aS8Vc5GVq55NogVeVUu6ILErT9Dp0AcAlqP5eo6R2
9OuI0xT8auX3kyoBjaEiHFpS0aYjfihmj8CfAG+W+b/ul3S46rAu9A5jWpUJRvT5
6CobJ+VyXUSjdlNvPiYLE/SLDE24LAQtb/B1nemBMHqesfMjnhOzXkguP5Vn+RP7
U8xe0EdI5Hn3AjSYJFZpsOYXC2YVghdhxz7Ny6AnGMPrljwmQfHk+ZMIa7XxqxiC
GNTd/TukIGwolg+3zF+aAXmxhBAMsE/P5HG8z555EAPq2EJXb3ny7sIlwtwaGG9n
rPw6w8GwLsab8GDk2QoqvCZPMGOxTcBOjYhxW8xwOGvd35/G/Zkwu5JfKPI5NlpA
vo3TIAx0tHN14ojtdw2mDlLXIrV2/RPZs/kghrP/BE+7GhBWI7wXLa+R+E6LWX6N
kV/Tqc4FwiSldtHToqV+mhbUDYHMOuUN1ry92A/s681zZyhykUPwV5s2s3mu7vib
EPNfuv0tI6iJ6IOK8wpeLxK6o4YIVBIQiVI5FRV0b4kXzNJgM479gjdS73fSzIaX
KuEYQbEkIEfX+vDa+AUmG1jgzjc/Vd9zSje7HZBxiDYFUGc61rrficoAIRxiXjXH
x5UdbN6YfBWjvcRTps6P9m3T6p5vV0zlKp1+gjvNyLr5TvPq2RNt0cL7w2YZztRX
a/Ib1eslIt3j41nDT+9+240ZC2SSCy5DuSul36HmHxWf0+mLttV2Qt34Lr6kBa+L
Q3pZv5i9na3OoSHfTeZyJFH8MIsQl2BZL8cbQb7/aeBNtwouANiTQXBaz0Ta0Azl
KJXbvVrYPdqUaoRp7lSaL0MxXJCnQwUjDv5MfifsWbYhPI3YUdYsClWpyNHJcYyO
Hp2NOszULfCi34IPfhwta2FAIQ8v2HX+XvUKWgKET12Yn7y42RD9RmErmVBCyquQ
CNrj5uu+coaT6PiWLbVhp5C36asL5yqoIOMKroTMKy76WtpUT5j1Zr01F7MjLGUc
cl57xXzD6c2TpLwGr+43SdSyL7Po45OuaXWhYZBQoBzLMUB3gq85/X826TUrh0lp
C3e+fUOqEwP4Dnduvxc8U4+gnCNmzf8Q934psSfEc0/rzZGBTnJ2I8uihfJuJrCJ
1ZfULI5JlDbxc6pnrKl4XXPcxUTByuC8omjh5t/c7nZlL5h3VICvfnmLvazeWqnL
MXN4L7GOCtc0fxXzh9sko0wOlV55m8zeDDZK/CioMOsFQ20k42jPfavbKZagXeOd
IOn/IrhNN39Ct0A7AocV+bRNwDkxLVKhTb1RJ9rlQCGqvdvXLA07y/yZu0iSyfoo
gIEGKRTeIlCStaVujtNtqVyZZjwpTwYpM7Jl2c+LQdeI3tqVPeOZNOARFNGLEk8k
Xd+V+i/KKi4zY1akL7aYsqd9kiL+PgHnANSO3dWfTSQvRgG7alMSO0z1TSmKrx8E
7XxDfAYJFaz2GDqZzR2QxTBA3WbqeZoCq2eiz46xxREFlZlfG1L41tzLfZERCZCW
zH3QTJI7u0/2C6eqyWdG8M124gWXq0jeIfx2W3YDqoCbaoq2GgbM95jwDRCDvp7T
nQtT1rP8wQO2K8mteEn7XO7lY+CaoOCpRJdyYHyfhvR7wLMvcR3mirUDcBb+6UW5
KTUrcMTjdCV5UzLi89onU7Al7RhiC1DDZFzDdAhhlnlFF9+lW+Dkpxp72LChzX7h
A1cz0jJtuck2bdmx/QBgEMp2zS6EbZGhy2GGxmdanDTch7YkZsbPpsI57lN0Rqtp
JNFnduk752p3N5wzURLLYa6DVnBy1MjvD9qOMkocClkxZlrhgCdoL65YTh1Twcq3
wIEIHX1yX91nZBeb6wS7smL7vFfOFcWkT7g5kMR4NYQljN8PPQOo87kM+PazClEv
Qwd+iMzehtgjf8BOmBZme7yKNzeYSG+JW5KtiilkNG3Wwkm6SaBX+TVsu10dE5JS
ws1Wmn506yhPqYYc0ra3jRHLNI/e2qbSAh74XWqJmUQ2RKG1UtVIAU65QdmojqnQ
lJThpFGclf9lfdrU8pw+8TINiiRynZQsib2NwhqZByXdYyo6T4a091YFlcc1B5zw
w6jRB+4pRzD00dnztO7mZSgtLvvNlNrBaKaXDnm8HpKYDD1Z2g1zX+UXLAhccbhZ
uw8cSdcvvJ055eId9l365wlH05V/hVEASjH/9d0ztDp9N0lp90zFvF9WuTFTrLra
Ibw8eLLpSWUoLLZn1ZF23ZLQB+im9AwRJlvIcvJLpIx1uph6E3nlHLOHn1+Z7uUN
DDkkYfgxCnq7i8xUvJQkRC0EFudhQOoBQsXM5SXaMlDED+ZBOjk8uTOExlyRJveL
vrXdl19kRuc/nF6vILTz1r7lnDN3TDjY2Z75snN9r7V9+rIAm+w7rG7E+rvdnd95
lQG/eE4Fsri9OM+tsUoh7iP+0vlxlPA7qH8qejcx91KFkmKF6DcbqEE6wIc8yRiH
uIFCoAsA5ZZZENihspqhxhbtAY22VkTefHyBw8VZkc8VkRrCN6DQWOjRDHl3DG7W
/OYrQiRud+fPdObEd4G90pucLay9EMx4ibIgsgmBYePKQRu4fl7zXNAQ94o7FE//
GeUz5z53hPDM1OiTbuzzsBy3nU7r7x91/33TuV8k/vPryRTqDip1stKTEUWxlNSk
/4EziQT5rBDFHof7+HWGCQonUFdtRb8lXUV9GzgeRwBSws50nd5qGIoDB5rg7Xtx
C0Z4Iiv3oz6u24xePO/FPQV0N+/ApSiCDnfEj2KvSD3OTWiwC0wl9a++IaBoCYj0
wM1iAktz+KjxpuzwqAlXl36ri4WDyp50hXpnPE5pqEwQ8gKtyDtvYWWoSBh8GDvp
nb2J2odgG1SydJU1M1U/VIskUsi+Mg+HLLcXD0KuLA5L9AaRFNWP6f5K6AyM/zmV
weh7oVuWk+IAHwI2EMxkJwualwb+4F93vk0c8pgwd5V5QjgMMvREK8B8XOuB/AHx
3w3yl0F4zKB5O+UEq71GEYvsMJpVrRR86wRKu3+EpVscAAa0LYp3Svq0PaKSr0rC
SlXMJ4irMdL1qo0ciCXaYslUeYnX4OcT60G8mSqigCdxsKREctmglTQujAfdLAUe
8zGzIrdzw9wK5TkHaK4KU7e6o1txpsWquDZq2xlZwQN8twkL7KXWXJLKiUYjhDnz
UaLRhy6Mt/LV6gWrvU+LArp0iP4K5K85ccidiBrs5HTDHr/rdA++liEwXzS/lUiY
hLCzxVrywuAJmhqV2X/axuS5+5+75d/RpWEeygMbFvano6mr9toBfryiffMK4ZkO
TZ8AV+Hf2/8/jTtgq0BITTWOYLh8hH9807k3C3EAxkCCsn3V/bImYMGAztgLZLwC
Dve+0CSLAdTyu2Y/kh63hiwBNHvpnMAG+6VaBDKLkJIkudTxfctl0KQVC3xcNvFw
IKzFIzfp6DQdAaFPSMscsA3WlKNaQQvhNtJTFBEKJDG5RbWQTyJ9KW6I7VAamqOZ
hqmVfs05omGmWYLiMJIKlhi0MdeFHpyvSOjkd7eCfYcWijGwLLZ0TsXj1aL7Ef7J
1N4L4x/z35mL6o8Sr3lJd3/p5HoK0b5AjFj2Hu9j6aQ6TMuBovJ4LJfkJpJmwtIL
k7APWHiIYDGVLnGHXmyR36VJy/hit00/EXgmCYR47fAV9Td9aC8jyZPe7KknABQl
2RlJLqrRHvUEV4FWbk1UThgKGaxS0dSmrt7kUNKh1+092WDO7eVq/7xUe9F44hTE
EsNaFYylEwOP5KvaK2wW+MEvMFqE4iWrJEeFjDeaqKp9BZCmf/5jAjeh+ECKKB9F
zKQ3yacuMNmBHQP1BSuadtUaptQ4D+w72OPlQpXRTFRMY336IRrv/vK3xsG8wdhK
1OsOHUlpse/mGtIZjF+F9fxtfgMi7p/OTN+Jn6D7X2gAqCewtv31+o29ElAGPiUQ
CSFBaA3r0mMMjxG+FVDJQBgO/xFxWPTZjLRgZCcJ0yV2NjQbrCivC0ZmtIchdCBg
uscd3aNrW7qySiW5fdETSMCHj7DdP78h/FmXgNGc2hSuV8QrB1LVfaqc3BOMr2HC
QgsAHELx2datC8VuvaWwPvHKXop13vauH6GMas1hFzAdJa1LPK8irVeGAjgNBqQx
vEtRKiJ1JU7Mg1uDkq/WgUCZe6ScSfeUqOaAYAEmh5C+U3T9nWi3DBGbjhWEngNS
AWhV1X816mAEfAxCdPEmjjDVPfHnIM1T2LGEOhEO3IQt16J3LZgC5cO80a9SHiPI
AZQNX+FHOTFQoMgZRUeRg1UCMYVki0kDeaKA3p5qjA8MhQZY/AAaE+vrtNysnJJV
WiDQJML2dajZfz/OJuRYtP02duVGBoaN9dB1PaMqRxKn4R7G8n2Vjjk1BmTJnlSy
3Q97pAkcEo0GjpI2m0aV1cxZ68ZAEicd04/Y5NG8mRsWSbBGQ9pjYdSm2uRBQ81u
PhsvEk4bFq788BNFruKj86JVgtghy5zoBIEbsw0ye80dYW8/K2GG83sgz8ik5Aml
dzhfciMYT51X30/CHrJww9TNNLF/BU7Pi1oOG+IlQuuR8EeUmkV2QnN+5bkyBuAO
A8CQ2i4YdHsge6hrEApc6rOfPp3XJgLheU38iRUnnGxlEe2EeeEAPRnp1Bv7b0BU
E6Y2OJCXfUZF1UHG6bp0ZhTDB19jibTTSniV6BnE7+Zhgm+jgrBhO3ffVoqvMo81
prcQIMZYQES+v+RFPQwDB0SzgKN0FHikCUWczMkn/WScPHRLEdpRy1a2L3lCclTc
Ty2S4MODBwPBhTMYxphT+rr1C9/fOhsOg1wFR1q1vcptEXMC+vH+ZW7W7vUbc1xT
jWxiaXPcbGPStZVa4pnidbhxWcrqy2O9hy9IY7yosAMNtqRw3YJj54pPuuiWrScl
mtNACEFFRxKCvO55LOZl4ezvs48iqaZ0Mz2WhE0C1XDoHd9/YkPFijEtC4ttC1U3
CEs994Wv9K4FRZQaMmL3TWUorSYUPj9cr3FZQaTcFkj08xkXEq80f0L3ds6ll6FC
o9DHXkNrKpaRk1lGa1aAiPVyRCrMJCGgSF42it7dKj/ZhbgX/r2Kf+SW+r7OaNj4
QygVITiUWsvol7FLz37XX/ZHDne6XsVkzn/M2qrqTIJFG69O3f/N4TuMg5AWe/E8
TdVs5Lss4Mo3y6CAd4PKHCkN1yuYTe0HB9UE3d8O/WVRwn3dlHfWJ1Ro8D5z8aJR
mwmc3uhFO0efC6RBofbKdOgKstDqL4Y8vB045a4EvRZofH22rDFO2H+TlfihaJP+
JdjYdJ0d8afEPCukokp1M7sE6v/5BIVkXO4YNOusPhCFtk3uy8Vvn9bsZIODDcC6
ax6c7wOXcGwQscpiuVWwQGUIvjDGhIGeZgKGptjAbKfqm63zYcrspx//f24e/lZG
zHrjaSNdnVZVtYTPkRfXTozLSzBj6p7fLdB6U4VEv9dwf/N7tc1QFHzpxAridMLO
CCNlbg+SptPUBxv2Mgy/PzbRNtKbCmBRZILeQ931n6eDa5UnBgKPdMH/2/8KlvTD
tV/DJJ05XCYPyWuah2oWvkMlhpOMS6wIS11frwBUpzukXtBMOu/Jqrj2kYpCDGsE
gCxTftaFS1k1Ol989MtWBx+xI789f2mW+ChjrCOgIfOBvyZZDjV9r2m1Bz6rlTlY
vEPMnoO07mP9syov+41bZnhiB7//HqDbO3jF66t/5AWTWLLxtQHuVZgZb3ptYqif
Imh0o2HlNy5MqYiutApBLI64jsuNzlQtKlD//UZO/orNf7VOU9lwXme86V+hArcZ
/XV/+3xscTbKX4XcdT1I+Ac24yYUmpiICSi+FbtAWbcArTPmxyzHPIf/VP4LjCVo
R2TMvg/sl8Gayo1dpvpxjkTBsMCEzUcrakZDd9upe8KkkjVVdoF4NEC9bZVf3mKY
t3ZOE8POzzI5hkh6BnO3ANIcKtcaAa9UCkfbkJ14iLtHPJ32KxGWEAxSiMHn6r+k
KhIN0qbDWZULLl5IBmMudi76cUscMDp90/QElvvgXV56nbmtltSkH7nZ53dKgdwz
FFXKG0qp4kwZTE1diMOLJ2rKV2tgRvZ8xwaM33VmB0VhaeCy5xWbPTFAYGR9zJjK
6GDcZEOcSqBNwUvkecFrzuoKcEQo0oW+ROz4XGdPoVDj8HD2kLCr2Sdk4gjs2HBJ
FnbTLi8KO1jH+8z8cn+usaRzUhe1MmkDPaRDuuOJaQxXbv+ZQlU6JFdrCw3tr1rP
IhRLX03dbkiLOOaBobcuRx5LomXrEM6caBp4fRUvkdQyPgmy94ViGGlQxIyWplMo
Wk9TFK9IdlJ7+tplgZBk6lBd6f4eXda4wxFZ1qi2zYlld2kRXoL17ELeYhPoAGEe
hGCfi5M0rx7bZfSYBUozM4waKWJ5joiJVvrYpbGjrwqPX/+V2OJ/wcCK7Az+nFpz
p0qkliYZCJyFi5uCXhKsUclbNtYlgLQFElRbBk+s3EwPH8reoNWj78bkLMvCvcK3
wD8B+LuPIUZhShYJ1CoIWGBtvNVzHsRAG14bE/FOdkSSYCsKry9e12ZM703B1OhU
pxe8EIvqhUo6Dj2O7TQPYrrViFeXW89RqjQQ+PINtY39/xVRYfPxdHuaJ9rny3Yy
5i1zM0IThgkr6T0fhqjPb+tTOhMOuTJYsPqYYajUfDSdC9fAzXMWOCOWRZXl6GAR
+P5gtkF4bUT2spj4ndC90Dw5WwfwJO5P2dlw298qYiInyYEE3YWcQvYSYcYXNpvP
LVTRgbdsZ3TzAdoNHl+OPqZcOR0Z1qfKyRuOgDg7J7pwpOiQQYZ6npNTD0ceAYRs
3gcdn4HpA7Gje2vWWe71HT5h/TOli6LA54lQB5VHGo95rEKdOZ+hqsCnWBdr8cWq
dqW6gTVmYqc7aTCYiZ7JLU5R6NT8XjWq5USwbCr9YeqNosqthssTy+6onEOQphnc
JQRfD4EB7YmyhTeViveGy/vYOtSfUWbsBrkF49ttxmV9MqIQPnETYgM6/zV2ElkQ
VNdZexkr7QY4frwXwkw2+d8Ng6jgu7X0I5c3QQ+z9YlcVAX/p2OC6ndl0WinYgd3
EoFrKda+JqaTWR+H2lRcU696/iaMVNCJ9h4ltH5i7timoNEfgAuzfwgxeQKtmOsg
O17miSYhjWHSab141ZHggjrKlRVrKlIFc83Nkrutn1HCq0XzvagPdNRkow1PoUDJ
bmdf1P8OXYNOJJWdEv+Uzm65puWY3oj//JRIQv7xGtKp/2UOxfwHoDTLbN9twaqM
BcbJo1aS67Bc5LGEtp69BCQCRxhLV/HTBvBWtgC2gn8a3J0NY87wIcujk2Rbk7ql
/SPIesPLY8OUmFoGBT+31EGfa8/6SgW9UlH1RyMYNNSvHJe2+aOh+FIzFvNgIDa8
ZxTVxoLxM34C+FcZRsxzPqCrm8ZyCZdxF+e3E6eHn9UEUBe5eyr6ztdLGjEfHSEl
cb6OsgUO1G6fmeqOMZffS1SRgPKd282ekmotjyz1X2n+9yFBDTowxjI9g/M+sp8c
+fZFcYV8MAJXfZ6XBrggwvCTjzAuKLjQokSj2withdsrFHUSofd+ruCpaHy04kCN
CKhCd9LtIkEK9xR+4uZk8bC7UGP8wQu3d3GOu6jRW7oU3uD1jUX0uSU/cKDMuY3Y
zXsDTkhuZCAC/HV3CSvluJRhu9Y66LqoG29VPaP3NRM5vBTz//jMfsDon3PoXAix
A5RPKsNBytm+TFXw9d4jUegvhbs5edDuSilT24v1VQbwNX4tCYKyQozq94CtDVgp
8nZP/PUL9tVK6Fp1xO9nZ6EZu0u48KOBv4+QBYIBaT9uWqGE8bxUPfGGsp+l+YuG
pqwMsyNHajzIB+CV9CJ8MV331Cjaoqyzf3z8WUmvbMu+y+ncfi+sNdwsnWrbmHG1
opmI4a8GkdAbydomyyF9iE4prb6WFCeJvmj2VCDk4iKMlf8f6yq1e9r4orTUOdgb
mgE6MEiFZEaDG6BURJVsl/NHleMA5T0vYV5G7G/kTSWAuLW87TzP4QuI1WhMKGIn
ACmQOXpCJ0iN62GFQhJYR4wnCPPZjq8/a1SfsFhLWxRsQbKGl9xJ4YEk/fMeGSw/
XkHmGa740YrZfLaqfUUSIwy3G6tz/StRQT09uyCbBFAI1SGv422EqYeHQ8UfAGYY
KkMTYp/604ukBsGCt4No2ouytIl8Lhq4L3oNQ8RKTXANAbLZo+B1CWk0Z3u0GtQ/
cKT55a/08iJxjVXsjSOEE5gPMlqP8cywYie2uBbGy4OYtJ5MMsa5xZ0HtCFTgjXO
mr1/AbLGFJh85XzpgN5ZPStiLRpWyvgY+W5ukuXvQnI34GZgMHS2bfRN9vqFwDfZ
Xz9sambqR4ZrtD1vud+dfKoUrq9+1RPaas35NpUhyved35rHaw4JF4G9OjQEx97l
EHh6UPu5yH7kgzfcx+IJ3lGV80iaArC/KixCSyBAwS0RjX9p43QyvxujJ7/aD+9q
PYznplbFeCRc1IvYKCngYDGQQDLIoGoSfjJfsQmxP9IUITmo4PcUs2AlMdX4uXIB
IoZwTqC512aFwXot73Ry0oo6BPX+IOX+N6lUu+X6tJrwdxe8swOsFSU8o2Xk+G2A
ShMw/AIEQ+Sy2WgYbltlMHc9PHmjKDkrswheNIT6y5jfl9zQm5/F+tr6gZw7jhIp
i6niUjPh3oL6m7mFOu1c91SjNnH3rYqXavK4G6+wkZCxjwHZkibsSeAHqDgHObws
7mE+bzwc3nsSqDh+xYf4FG2/chjuCVUFQ9migdpcYLfzxw4r6WdcSAcUzq8NjkCo
mJaQqAWhPO7I+YTh886K2iWa4ui+wAg1HZdW6GYl9qx5TMraKD+oAgJdiSBPKnqt
14pt5ATvdEIJgXjnBQxwSaIWcMBDuntWDrppiNPA+sOtnuTvRKT40o9f9H1cZWt+
95tRRx0UMhl6lE5FCdLG5/JsQUmfffSykE+ho30m6w4AUUaV/V5pNSgFCFgcmT5D
imI3iHwhCroW4ZP337wlA1nQuiTUpCKoythbO5Hehm5MgBM9o1zuGdlg7zqv4tXa
TmDW+up6MKkfUwLFbWf0DH1UXXCdlhXpM7g7LHWKzfkq+m5tuVBGVtNQ+yROtH/f
QsJAfwnoWh4ZKr1+9ogh65wUtfw+looyRAhUJoKu+jZJDzy8RiO9pcGTUo6Cy8x0
BANSdOszvN4rXOOuljXH397EvnZBOGMYXHqzRvhjltmDzdJ74rW3j3St1HYwzGq+
Ih+7ayPfsibew2IbEoRiTYM9Mbn9DProp0VrSGXBNi9ycVuFkL9UlsEud30pOjpC
xnIvyoQNbPofniUM1Z3KzX7m0TkHuEeDWVFdZimaHA42RdVy2gnZFoOmQMygNr0r
Ke+5JDFZ8yunYQPkZZGjV1GLmOPkOlotU7OIXRXkkYBzZL8zehMOaFrw9qibI99/
HVuqTnV0BJ8+R8Lb0rRBO9ukcXBPrttI6GAYHWN0wzIhujwxQBvA/XAcrr9OyFp0
ASnB3LxtFA2Y+7O0Z+VYnAksGg+iVkXM0oKtFiNBADJmwTJrj2zadzN92eXvkvBw
gu6XvfI0IkYFYsp61zp/b9NsKLd96l3fYoCdCM6UaMhmjXlFMMSV5uOZ7ETWiCIF
0Humr3RQ07CvTIbYLGe+52KykMKInsInzlnBd5F/OIkUsiGrjeFe4EWN2dK3GlD8
lAtXcm5CQk5eI2kYVaFIjOokNuQSLF7BqTyF5fcPUCe/kpksaFdZL1fQAi+xATlz
brTBnlurzDC9AUu/uxuF/HyDKQv/xbpzIXTZ5Vg5Qk+/E5guRp7WLa/dEA3IVXvK
o7WLPlgHTqLSYNDzXgGFm1FIZ0tPY2D07T0ZD6RdTfObI0p+iQRYh2pabgupIF14
wgQRA9kQu6s4IpwObmLubRqanbTueT9hlyHXZMPl6c5Yf/TuLPKxLZwv6rq4b0Bs
Hu3jqtp5SkszTe5RdHjcxKqxjeC8VlRDvydm0xgqmV2MOKRm1gIj0OuxdtfTkbGX
E5jy5ulB7DYnM4r93wpBkeQAteMlSMo5CeAQI4VrTtzVjX3LDCJEF5naVVck+ibX
p1vxshLrsyEm68wy3zEGfomkdWg0zL3nYKvUOt2tgGrm2I/jd0QRDXKAYVwgBHLs
Nsk7wq+Qyk28Es8ALRRuhly023/CkN12kHw7f8VAjP2scVUY2hDXl2Je9rPYnvJR
NIX6GOhmKYFXxSG5X8TpRYihoG2QyqkF0il1AZ7GpWyYNEvcJWriRQuWUWRhT69E
ZF//WzoobO6epieNDIexZwRTM/lxUkcD7uvAIGt0qbxAPBIUo0CGY7GIOQDKcNIM
k7G4ddAVbedVLcLAi/9K+z4PMC8xHqAxMPJyPqurR5VMrIJ9jjQ0NzKuLzj5YuWY
sZxm1yNbQdNcGFOfZYPnsYNTb79/grpXWMEeqMpI+YFSuB6PZ9PWAFK54iX+BicT
SVoh62OLEtFWbRga20IbEn7QxWfm4P16RIxWU98+YmOmAn7eAj8iGi7nWNBgHU5/
8qXSRRoiKnFtPWC3rBcMEPgbUh0kgD0U7Uh0pW+WCSHcaoHBicaONzpUdzUNDoUx
RT+xtRdjkPXCDcIifTHQhc7q3Vk5gLEcXPV31/rNCYFkhUVOAbNBiozYOas6kEhh
C7CqS3Vuj3ZV3IPGYyWnAipsmgdTR/G7HAa8r06DSSgUUio+DGZVnDa4WbH5WENN
od3rKkKTP9TsO9U3c23AelsrZS8BZuZ8CN2pJs9VEUeRlQSBWG7IcJhWg4SlaOpZ
TnBWmBCl1edvXEW5wBNXJJnfQo5a3le03bdeY2tpE/OJUmIxXh/TufIcE4UqtQWW
2niKtZbX47h5vKtC+9FOWFBHwJGC9BL6R8LGvH/41gwIzok14c+u6N/60vWEF0Zy
AEbm1uOKbLKNDiN+FBmlOuLsGuXHpmC7ht6vGaosYZABPDJvtR8UwT7wBHIpTzP/
18lPNo/gL2BtJfQ1vQrYnpreASFamGtCBajgoMgH/t0w+8EJvn3UYZuoXt+5NHjM
vIEid/C0Ks39nGKdfFVZ8u7u1RIIWmBV9gzDDMvplgY1hDnVQ1qeQGRTisvAuilA
juPvdwJPZ2GaacEazKsH0LFpxrU5FH3QZr13/UGExrMQSisdaK5jyMDHURQjitHl
EOymwEeVBHiCd5XsgZNIYaRmbfPbgPafbTnmrKfzItq3twoJHdcb5rdd8TupfMs0
a8fT+mdyRlGKyetgEy3l0chLNrd6Hwx1HQwwWOhBNlVWN1CDkKIOplwXk/kClaf5
AjNoLHU1ZkD0RZQVFKIALkthp9JdF+WBWsp/JllElRJA2lDMjiY2LX5C3OsfO1Mr
lg+BWLwepViBfKy3TLVnlv7mzeZQuPlR/rsoYKVY3JTs5p49y5RJUzutI2y1qhYJ
+LRX1nLCD5l7Vh2VczfEQYp6/C9S5lIcLWcqxkhtaXEAGrejNxURDMBpwR1jDxgv
RtNnJ/hfehQvCmXUcR2DWrA33V55aQaUdf+hT3jWtPOQsZWgXUmn9K0DNAPFEB27
XR+JwxCAIzugqtsEf4S8TY5FY91Ro4Q8GgGQ9JTvxytTt7ENkhrb9hDrllJWxlH6
OWfzeZ4EYeBsE9yYLePWbrbKBn2mAknM1rC2AuUqCUGUUNp7YugMUHCFzy6kWTWw
TCSXDEFWUxh5qIQwsu8q7wdvDT/1t0tFDa1eNOIjNMSFeCKha7ZF8qklI3nwA9oQ
d7vGceJf7KWfw0xVAd4ACuQ4rfaY8BipAKKzTkcGdspYBQNWA4qYtSjO+d5siq2i
D4m3z7WWrWw3EYoDZYx6bWk8ykiz5GzTDkM0+v8iX6J4VtWFuSYULR2Ksd8rm3Li
chHhTrYht/mxGu0E2re9Wn3cVQ5dtUB3/Bo/ydQ++dPqpx8ie/QTT7F06L18cEOE
fhcul0wJctSERP1foiRErO13bOIGG4axhocYcsG/p+prxWdtakgbYOhPQEgGf+ni
F9DBvLRT7eaYiRYXb4HJEXBpcnxBf77VpLfmwx+HKTAP6MLRF9oKhrYUKM7WX+uR
N6Myyd0MnaZLMLvFt1C4TEkjLgBzbhh/I/4shAFpLbWa08oTY69dZ7i4J1s3Vixh
cB6vFculL9bkZMLpqIqtK8kp1aie8b9C47G5DL9IlOsWZuMclcokwvtL7C2v8sB1
JKuYJDds8KUZRVbVSzOW/S55n6JrEVZ/CT5DrEkswgUzAKUP6ixavmLNVjFPqDg9
JAnc0IA6dQJ3oYpeQqoWHnDTOZVkPlT18tB0ZqqLyV7Bc5OMoYSX2U22J9siZ2WP
dYo79ewNdJIMCHMFSvbo6naxrp2kHSiYaokPyKbn/cxlmaMyhccgIa1oh9GUZ5Fk
posUAwTvwE42bgwO7f010Se7dHTn4cVw6B5MH9GUDF49bXYueExhPWXDTBHsM/Pm
uixjOHkKEKR4rjNqZ2aGUXieLNNPXxrhEtKP/7gg49yT/3cBZDjnoJvs5730enEC
+jdhOZ7CZ0GrNTpTPobDZMAIO8tta0d4n8tLYin6Eo24aCqGexBeRS1jSfczqe/w
qDusxZ9ptL+3k3yuzMsG47kK2Bc+CCiVn33V8wfOEzy3TRgvh66UfVJ5bd+qeKTg
zsntmgZFMh9Af7BIBX7xi15+1y5CSkvGyoWWoAX/sbDbbJtTaGZQzA566kSBNYvF
LTuGRPkN3JinEbxlMg8pTc7sP4ySqNfTyi1SaOnWXfkOFiY1aX6o2uKzOaHGqhYu
Dg2q2HNVvGtcRHg3lx81vXV1ElwWrKow3kCXhkUrKYNti9Bkc/rkTq2ngZRyrb/d
d2LaTYCCVgK6R5OPyUkvCqzRaKQ+QDP3VT6lz+t8wNpIUiMKH4Zxhckhk4zYx/WB
n4OyTUZcrUB4apGft6ePCV2aSKowIzLDm3qpmeEn1et1fbaEZ80Rq95kWsYnoU8I
FCrSx8ak8gycrCYi/r2nAPq9wj683HJaoHIqfiw8iB1eeLjt20TNsPnjp64indmk
Yz28eIC85ugEr4w0V+yysJpyO5XhB11QpWWITomcoG3N5FducoGagzopobcvOtr9
Nn0NUxshgquM9K/2dtE4f4U1ebARim753jP3RXQo1rReZXh1eHqGfexcH5ktr0Zc
b+1Q82YMPO/WGmETr376YGXZ2s57HhIglL0hS6C1Skqgj5ljcG2l4v8EMhIOxE00
7Fxx115k5iq5LP4wdlCc05zRSCtJYYAJNLoisgBBVVtfvO+Ec4FOuXg8ixRM1hMc
iIP2a3R8YdCr2Vrv6/JdeB6rHG6emf3ccu9ZZsRFrnbKrmc7CDw0b7/5nV5AUVsM
5zwC1XsmuIS71Rae6Kq85kSfuZ5BAFPiBQXTxMzjcdV7uywAEmkhPcR1cioYSGw5
3sG6O85svtqbRYy+FVYWX0Lg+S3Sw2S/z7yVyNzpFfR+t3OxrDy2ed8CkmS84dKU
n/GydJbvtPbip1yada+u0mAnzz/G6dIt2dwB/Zj8QFfdAqh4+onGe7tyBAYwF8zU
0eFL/BubDS3YEtdB9yMYeAqbkXJ7nMREDSZy9f/D3nAQNc0II/AXAJf5hfkWtHFU
ts4DoxV4ZTJd+5wU2T12P1K/tPJiU3Yavc0E6bCwxjy3EUaX3wy0OkXX6Kw2t1PP
bs4h8enPPJxrJ9dvnl961yZ4SFBBfn3DXN8nQrl0mMEpTtjsXGgaJtEAIp1cr3GE
qW6KosD5MFeStl/zgNhUnHFzOYh00yw+3Lu6B8MZbYJJfVXNe8snw4ujA0t8KXqV
2IBlClYJu3IG7YX/hhkal29xvuBvS0pABe27yRF76YIPPCs1TK8X489WALK8gkix
ueCBTd30u8LfbpuAx9HzCVFj1SruUIWaR3QnO7q4LqpWTCqgfu329zVSZMRmNWuP
SekehREfLCDwjKsWB+rK5mRfu8PtkgufO623H4jBjeojufdT7jytvQptQ5XldH6o
swEuVk0Uj7Ob6mZx1FNkf/3gVJ5A6ynDIu98EyNvk1zQc8ncd5jinfCJLvZ8c9s7
Js8pJSUj2NT/utRsisuaiq2DjBDDWAXPQWkLQTX7dMamHT/DQZ2M0SRNk6TjQNpd
3JSmKNJ2BONBB8EaGauGkvgs+3I1B7kSU9/BfTZBhVBC0y6H5QgspO5JjP1sdxYn
Dc2MhldG6kvMcJvqhGa9oEWgrkQ/OkmyqY7TKSC90vluIESdgWVWOg9nuiZo8dy6
SGuVAt6GA48zeq0GmrESm6k2zmGfqD94ar/vfMTYmdwUy39e+wTrD2riSHVE715S
2nvLuUwYrVx9XYaPXkSoTBGlpHy2o6naUvMCc8e4WHFCZwAHUzMmTz+8UuPoVFHJ
bFTs3z4+KPp7s1n/MlM8+4hT4O2nYxWtkEKw1TXeLlihjwGznYc16tP8o4vL2UXy
yxqnGTQOkQqoY+8ZqM5QxAiMYbn0B0ympLZFduWnl0j3x4xsbuQ6qjlXf1oakgvW
wcNDqCfkMsvAEEGUyN8cbmy3wpwYuhwTi5QVbEKBX+XQzfFEASKfU31weJqrDzSR
M3gKyhO3ElBqDKydaa1aZmQbyMgdZU1BQmpAJXRtSYdGc2pKof+MPeu6QSTbVtPa
G9bLUj2YPJv87thAYsZuPWxwQEgbwbCCUl2oCiiwH6ODj3rd/Ywa431kqriiF6pg
KiGtNStwjbNYRj+DDBs79IavKayAme/+dqyzc2luHpdzFurl9td1unCkreU0SmMf
s/hZnY3nABmciH+ap/V2ujjG3NzNHeFSf4i5I9+1125wzGYPmN2xUbSx8clf1vi7
BGKrSVs4rm1CQIRmJpFtCT2VnG20IiP6t16RyDBVsoUk/7/qLLkTb7wsIc/FmaPI
crw61Upqm2ti6ghAV8VgfvNa7suiimbz8a1nCWsm+TKru0fnKeCtGdqgimdGFaoa
fZYRfBseG/L28dsUNZGgKaoOrAoKRR98oVhSk9uUa4gzVAU2LlnH+yVPNkIk+X4O
+rvh78iFx1NCaXtMXND6GXGZUpYPwaHPhXRuPpYyaVhwCbg8VdFbIQsCrTqx6k1A
/O6GuN3qEhSc5WnIrz6692QsdwV5lYyE1c9zy7Z1aNn6c0tr38EwnC8alwcs6p6C
QEtNWmu5hgCERUhnasgvbdcPIfeJiycNokLwt7N/xl3o6XBopQqx5Lmn0Ro/tlM+
jF8KxBEiLvZkn13jVrufegoYxC55G5YQkMt7kWQQ7kvuPSB+KEsE1eZiadyNHesh
qD4FN3BnGqoxRV4V+LZp6sC1hkcqfyjI8qBgqvaDZ+/I7aUDcSGmUCqouWB9hacO
BL5YKVMUwy5tP0pwodz0OmNBQtmZoxIBItX042L3wuAOBJLChFUZkSUElIdDT69f
+EA9xTDrY6ajXKVWt2cEKVTCZCiyoZwBg2t01s/+z/4N+zMMaDFBzv5BSF18eslk
CSS0bi5mE3KM59dzHIDx2qn7kAUtG2sWaaV8HPu//HU1A+KkVJOAiMchdaHCLPeV
qp+1C5Z/AryxbHi/PQdPY3d0kdMQOWYSNo5H0bR4b+vWUordapud60Bx4a7KAQOz
GNfDGhSSaWDq3pg9hVqQAjA6yKgZI2v2WjSTq3oFcHpOSKpjV400a+0+Ut5BPNcS
43tnBr6RSISd7yT5qIrr2ibF4Jz/TobhGg3OCfa8aRPkTRZJs4KdOJ40TUTqNGoO
+yMGchmlHQrxvBH86ye5nRupPS5rRhuUYkovn3vMYGX5SXwzO4ghj9JQC7/vz+xJ
CfR+nJ2vLaCxCDhKw50pbydRE6VDzZ6faoQiiypUyefSMzOzNsiRufTQOPqfSPrw
9SY5CgPWlwO7gXpvNzO9y5xX6sDhA+6x7LFVKMh0tqkHLr7m82F9XcBEagfOHE5X
4oQAAP3e7qx7yrHvvq4q5gEhDHltCbQEG3x+0d4XsdP+NiCFTVO5/X4AMhXdNwOS
FbkSLLgGcYFJEdoR2blljigJoIa845un8daY8FMT+86BwzDm5S4zatxdiNdbOzu1
8yYxam2DGuZhuuFkaOgm5lkIZsjtTOK8LdY7kcsBI13gcdOe8N42hYMD+IBcd5Aq
exijqv7rFTAR4RcPvfX3LD8dpjSeY6JjX8k90Vye3gEU+qbiRa8IRzvQNvpyEKai
ZPYMkYcYu68+LrfMGcHi42aJXNkkw+cbosrwQWS+XXiza6qtLKSqYH9EOBzT23po
4VrvcDwIXSin5LLQi91WGjVs2GAakjswXp41F4G55dpizBLr38fNnMmkaasyiOae
quxOgNUELDRo70oL/NA3jW1HjtAxN6yJDGMugdmjNqzrsu0v3DEQn5lGdFs83Lbx
tNNMBFXbK7ohAnskT39RZfGzTYzu3yysm5g0TGF4YdyR0jIgTWtJsPUZ1nCbSi/Z
qG5gZw4cl+tZEeXjcJamIpibHmPYlLVqFHtOlkLXlVykWRvdVYr290TO0I4ypMKF
VREEkO+XBj+gea8W0etADjJMdlRmGLXDEzAJpVerrGXak7Obdh/sAYyXDiqrRp3v
ebS795PiTfSbJ+vpNiuC8N2QH2IQIrcoAYG01d8Njd5LNJXCRjMCC6WC5GilyAo4
3P6QTQNLq8qLOQxTEMUgPEnxS2UVcyqEMltPql/fcEKcDT4Yf4/UGKu7oHy+VeVY
bBYitl7nzkkHyEAED+byxSgtlE/aceNDk56lkg3GehDb+3l62iYPMS46Hu2fuXOm
0oASkHRvXRRctxBBHQUTSlGFZnXpizn9wE63FIyh4VJbSfNr23eoV1wrwjJZ7yW6
8TMVh+UyokrV7wfQ9zxyWOdf8moIF0wpRaLHT5lSC9OqyD+Ynw07EHeIgsvLebYm
UJclXRSaeM+Rel7VJBQLsrk87SScTNaHC5827/3Rmga7l6f6/UAXGiy+8CeKIgpU
z4vLaiQWB58/vYIiaAIMEnDi+TLRE88sQrjXwG8gT39XwmwtqewZ+QLTDuCTMxkG
aYjyYwv1nVLffBEhpuMAxa29TEZZ1LOL1fhPbGNk5w+Q4F8KT/PxjjJdr+zzElSH
XNJXTjAVdcjepjz3/9sXa/dRq6v/TdjSLeYEB5IKgZ8Cvyq5Li5hI8XbL3VnYXE+
pq+WkkndIMGJMKgZeDDAlRvVXGP/TfQEHL2dr7Q2XiAhyED9mTuX9K8Ky5WDlwl/
woq0BZGITTUBjQPY3IEYnNaYBTkRuH3x+lOckbEjkvH51L9JPXYMciRGyS7BaKq2
tCZCOOCQGSbNc3WvebI0LmluIzjftltwrBDE2wskCLnwrlrJdu2djQ+C2BkdceXr
0JvvkxgjVOkY+rDaY7KxZR+Y0DCYyvKtd1++CrWHbEj5XmsIWDAERakh2sifM7u5
hsYQfMojq4WLIuqLlv5tVFoYC46ozJ+bOEjaPUgeuI29sXwCQ3Co718x56yo+qnK
yqMj+OxcugDp91hM51/C4QlhPT12xpqoekw0Uxyy5mOiiukYzGtDjDsXBsJ7usF+
F8qCpzE3XJyN8uVkVBH7QZjTWVSD2Wv4Njmnj+S9pqHczLKzXaXgwIk3qLOS14Rg
x6uHzbpXQPUXNASoa3CrflfdSyVaVPR7y1k6gs4GpL5vrZc+R5cSrkWEO49Pbf3H
uhrK1+gQMAzId4R9NZMCezToanfVQgcHoewbbUu9K3Knur/8VjpLXLKqziujmaT/
Hsdgqu4iTBSmTa21yicHE9gVIl575s25EZfVYuTX4RD+5w3A+gowtR1YORRon0Zm
fWnfbohCOhd5rZPu1y0BRhubiLPB2tDVF0OhyWbOU0laavKrF6rbV426yvE7UGRc
uqtsk+9hQUcVYHRBkoaITZd3AqmTyr/TjAwTov4P9YpoUweh5Vzzwg/E6Sc47t/D
OUiAj7D9tDARnkO6EPAI1gvyEhodH6oIeK1zzTZfPkRoLZw97RAdQmGlHcUT1JGN
Y+eEnIToUsbKcMm/wx6J4qbvp32QuljmqKAYTpTvWPwr+CoDrmFxLzerRoBkfL0C
aKm5VT8wF4w5Aj9aismyfvysK571b5zVQPRJqFvhe2VzFQp2T3gg55inO5bSVxCz
btzzkmj/EJa9KnrAtaD+82SWNI0nHrLoqzdZxYVP/8Xw/Bgp5EDVguae2FhG5Pt6
mhC5HTtLwMMjXzpqhg1ZzKTtBQZqUNzxngyKzMnHCIWMAqay6xl/hYNd16Arv5dj
6tkkAE6dzUik9UTC/cFrsrOj1kimqcH4+eWiLGHbBfbFDWvi4LWJWUlT1xDsF4ZO
jiwxKTT+T1caFFVLkgmfbn4f46I9t8BpEBYQamWQeCxfheQsuQNCP4C+fjdpKNam
sS+3E+uvRsEU2lZiew+smv/oxdCJnT0hRIjwhJDC+lpU4Yn50H0p+m0lSfPH4dTW
0LDxmAfaahhoyq8mB/lZcrmKRn+z9uEnfgbGiHuECKrr7/OW3do0F16wObXypy+8
payUq4k1rJKIpb8DogtDVTDfvCjakFeEGSqavoMvXVDpGt/tXVaqoAFW8uZqGNQ9
cuvjmOhW/1lovQ9F+OA7JjVmFWtQxlfOuCxx+hfTAKdxCk7YhY858iA1RGE0buYX
XktAMavhTUpZacnHRn2QVsefop1eU1dR6HJRaV+oplcm+TFAJ6KA6oZDBU/UUQXy
cYanVZhCvr7vMLZhuHHytjZMwt5r2OEf16zx3GAgCRvYfGmInssKhS/Or2JkiHBU
wwtL8Y6PEFvxE52Vt3tMMefS4gtuRjpb3O3Oy1D0neYAurINuGxmbZXIIHPf7SpN
jIt5RdgPpFF4esKO03jVinkIst98/WxdUliFuLF/B5V2HI9LGk36959N5Jj5VDGB
OlZJmb55uc/mrcFZ8QWkLC1dYnR7PbJs4EGvfh/+9KUoXYwe2/FK9ah8b6D8CTcw
FNaJ+NTLyojx1PRXoTAlm6Qm8DD0jvZvUoUKlMwQyN6yCeSD8H8aawenTwFRrAmS
NRVJQvtE03tjJh+QmBs9j7HYO4ornK7bvm92SBPXCP5KuqwwkGjkydJQnfIS2o8C
DUMePx5deTGuXW+O5dJ2l+jveOjNEqFlElYioHNJRZ83jHfYQzz428QPx6QO57eP
RqQcogOlUMv7qDOFFJ45/i27MjHj26bIsI3jndB41bGaf0qGC3dqNfYxK7uoww79
siSF8qRfboK7S8a/oNtu933I1vMaVIR3dHkDAZnPCPEo5fmsUDHOhKbUfuEvzOga
12oI5fWIwasAuMc7B/p2WWwb/Hac4kc38G9GhA1Awt2Q+lwB1GM23myhn/fCd+wd
2itrSpz6wkXYFQIeQ89exMNcXoApbWfarcE1ZXGQpuy113lJc1K1pXSB9G3Q1ycp
I1nQQvjYf44g4VEkPBq8VIrPUoEb/z9pcMX7LJIyFnKmiDaYYLh79ofukYLtxNph
xV6v0j7WtAXE5PcurEqQAdGeCODTREMoODLpx6PDDVhIkVhDjEmwgti9KP5jDhEi
Yz9Y6lT5fOPwSnCvcv/QZy4rFsQGxKkECdBV1pSNO0bucBNfVWGrYpU1PRUlG4YS
Ijr5Qtrpk1JzQfaLP0Ju49UwyvIqahoxBvwWu2vD4TYaqEwVto8db25bKZFltc99
39eoI+72kxsIY64E9IxeO58KqSXh/7cdCAdcLE7WoUAG1GPeVkceh19DOh4mQi/d
hhIDRktkTuhZd3+PVPGlPK/FS+ek3i+2FUEuLkpc3/Ke2/SkUoLHIvm6ToSsXGAo
6YxIx1LToVv9HNqz6SbxAuxsO3pKOuG5zmuwDGLscHlbfVTk+BOutHHfqdUc0U7N
Xua2FntDE0Tq7El8SIAutJBEHVnzII2v38XDgI29jl6EAcaFnKF8KSii5QoH4mIU
F5oCeH612jonr8w7bNbrWsZ9AdfMC+WLs9iIwg0gs2hRi/UUL99F7OxC2F47nw46
nxV0zWKxHRisbyHizuRjaax9fh4Gvro30n+fJFRpPYEyUwxMvO5O9UdoWmm9wV6Z
XCxL2n/N2ygBAqwUjR8CZ7shh/V+lDTNu7PJ0kIPDAyWDJ33mJAJ07qNC1VjvEg4
XpzNZAaX8sfIAQBQkqtkVfm47pRjm6VBTpOXKcmZpBebjcjezjgwemHcPjcw3xYl
uLCNI2uaY0DnTl0wR7gOpk+OfIQN1J1yCAFRA6G70QJjfUrWcSouLHa7YwF8Hc2r
H+JiQ56LP1nexYMPFtsBMkgmgFErJCE/TNyJ/U2ImudoEvULW1nreM/8+a2l+MAf
lzWKkqBsFSf78R+0J++QSISsr11xmuPsq0eqZzH988vc4TrgLHRyvhdbh84FBZjl
Cnb0vuWeOtGfeTvsu31TzfGNelR911X6Ohue0fdetCw810TfozJCJF4K0XwBwgYR
DHhzOvZSLaZsd7BMm8JLyyw8pEaCtnJ2ORr8YhnP2C9NuPb+cy2b6MT8jqFiUwSZ
q2ZC5uKMb8ubUjHuGRRx7MQcfsGZqgYBl+uNWFj/tQe7SbMTzjkn/aePkKsP9IvR
fd0zVgcBDp1htGf3bpAXmUPOWM2BIOONKazqF7mVlvKG0al8wkM7pRmxNoS01c+k
ItDwHp/Tp+0L9RkdW4iGrIJK+foQ0M6/Qmgj6dOI6gtYwo92DRX5Y87s1oWsgbYw
+60fGauup6y0vr9HYpO9OnROU5nXrTeBy8m2FkqXsm0m16QaZh5W5+LHMCo52y06
DZbgwG77RDJnEKFkyKPGGBW2RRZ2bYAj6sMo5zKPSIiELJmPQP2IxMJdjJjdUEGj
sxkBjGADn4eptbIb8a5D/PN9YUiN0Vsr0uOJLwvI4brczd1OY1RmaFHB0d0BJMtT
k82HLoRkNSsl54n8LrGIvgKiPpaxvaWElnZ5v7O10DmDfa8Gn1GSvbcFWK49ix0w
zYGXZ+0L0ahL/4Zt8QXgjJCGSiwWYmwMlqQa4zbRUVptoBl8iUdj8KyvjE6+XT6y
jR0oFgPV8012gfGRNmsjQ+K1gUdvc0Bty02UDvhzqA4Rfm91/5lBLW8v6+FcTcpd
PXhmOJmXxXHVM5Nay8YV0WHCQrzRCXBhkrz9dzn4lEYOlwwJHcLYB4ZycCwpjEr8
x5eTXD69fRfZt9v0u8g5dzC0qv4VmAuHyJdm8sXAhtMNyiUPiwvsLGKuXLh1UJnZ
BbS1hSN+81bdl9IhF1U30yexwsXDzFUODNHw/q1DrmZNqJC4Lq01Ql/ZY4hdjRqj
fM+Lu/9tcDhS5rjiY50fnJpmO+3VIjvCviyrgehX0m107L68Wx1FYkye3uvP0ORo
NVU7Ta4aFARshuI1avtpxJHXtTCYHmxJICFXZFwrgLBl4pN/g5W6pWOz5d9Wsw++
1FoNdC3KOFGoE9RkJpJMD079DmTJ2S2YgeF9cQIjPJd+st9TM1yzvdurMyHjsZu/
RfMQu2wG9Kl7EKF1xfeQwIMH/MB+znQBPJThKVZ0+x/uV6cXvpDbGweenQyxSIp5
HDgRu5ZOYiVZgyMgmsuf4KWCGeqf5MlgPOeGXQlQ3jjj58DH+eTj2v7e/QWMFwuq
ZHGIHudXFFmaVOI01SJjRo976TPZgnOboYHRkcWCQLzXmVbndWvc4i1ymv6qyjG9
3xxnalMGhTr5x8G8SfdS5H7EPr5wxrLy72mACAFB9v5WOZudrrR4IWr2xOoj7Su2
DWlHcEOdnT5q+5sliJ1mqwojhjAdPcfaj/jevjW1KosJHTzxZ1eWT8Qf7yHRKhYU
TttZDTPD4Qfm+KDOIvmPilqXTcxrz9FUCFEQKU53x3YUqt8LP+S84dTfHOyflCqY
lhd7plH3c5pVdIaBJv8vlUTXHFF89Evm6JYxqqysKBayLcdBKU4PtHvQ04tLgLfW
gw92imQj99bZnN3Ys4aNRhsX6kFuEd+5+3iDpsfpWAXhOr9TOkcuFMtQzQwQ+rJG
0znHmKxJ4jXfah5SmEuRaAtje4d63tHu5jNR6A/NW5m7I0LlL/WOQAeNICsMlErO
Lh/G10A9oxrLCxKsFzazKqUuEo/6v80jwRxdFfe7fDhqGO/Nh8oD+0tTlDe4FXrl
J2BPE3VIDooWFnB075RyCMvhglPGH8Cb9z6kuoIk9ngS+KlNyQ/blwsU71eKjZke
YN6TRRCYyL3UID85uXjQCwCRfj5p8P9A+mFEL+oA1tg9HfQwu6R7hTKrNXb2KrBy
lv8yXQhO++954atNqBZWDZGAawSPmcY6k3weqXUq+S0TRb/5I6VvrxE+ecRYmsGU
cmzBKqvFUQcxJfxMzvp6j3BTZzyYvJ7k4HUsCOJfKbnAhWu2oGk4ndY/IQ9QjL+Y
lbxX2bYqNpFnjcnPeQrLalaR69UfKxcI83GhTQSxvmjwgrBZyyCNeUJp0RyedAaY
ato2yQNfpXtwA5dLrTihtOW4ghZh35FfQjrhfzEarTJJ3QUeCqWrNT7jalM5pBBc
yu175Pi3N6zeOcDJHwNReLI2IS7eyANOIgjjfK1r4dQglHl4bYJnRFMUSr1NFr5X
ASrn8LY/MfprnzWNwKXEy5LwPxQanp7IPaIuLR35fZs70q0f9mb3tAFfd0j+EDtV
5o+VS4jGq21cWhBjvXqHw7lr4yp+jsrzV4FPZ4D7Ec6IS84ZssX8lAqFyJOmi7OP
bE378MvkfCLyqxwErfeWyS7t1UNX+N6h+yCLP5QhuagTff2sYL8uFHiNKm2HiZb1
93gUgFH53ngRZfhBT+cU/jJiloVL2H2qi1kXgLMl37b28wv2aYy+DQuDgl1amTVO
n3N6BvwY0lUNdthQe21cwoGa/D4eP66Tz/TEscZj/dyrEpary8wQCTJ6z2tp9DX7
ZkJkZK4BCK/GR5QVfs0zuK4d+Kh/8BxiOzhT/SqwQRdRv42ifelRCOEXlziautuZ
d/kg95Gz1xFSWiBh2VteJnxbicRq6Z0iSMHB0VnThz7R9EnJSu3wUFA6303UwCau
eeNUd6XmKmRx69uafj+6Ipdt8XumuqTgbxDQFmuI7fu2kkOQrBVEvvHwVqo53O4o
9ZgyQF17QI4EdEAo5wkuWWtyCoCD188aVJt9ADikjRaOuHmZtr3mpGPXd6mTJZRD
FQ5ovpfs0l7sxkOBrGtmfGE3RaQvAyyNi3juBwNM1hOyQ0F+KyeKtbrqNY40H3dm
1Muy2+L8ebgiK/6e6Fr1j25rs+ukjy1aEMxaHjM9fb3lx7CSW0fvn7IR4J82g3uN
pykmOaurL6sr4iR2gnyubmqmyC7V+Ft6Nvs9aK0c5J3CzF3s1pc3iWEJ9LeWESwA
l1g7RXEbINJD33bCmpkfDn51k0A7uLfDHeeLWaUd3pKjzgWABLg1TmhxrOgHaMVo
pH6pVX77ehGVHf275B5qdRISt8a1KM2vuAIdqBuIeyq402GHxjwTWCS/YtKTkCw9
Bo3KXBHdVt/c0bvHEON0zakxjfRM63Epnq1qh6mYbLvU5kUCKKsm8FstP2lKJlV0
lq70Xb3tXhKNPffLDWavSvAgqP6Mn88r7TlG8mPaSzbnzTqgl9W5L5VQyv82I1Ea
IDaD0qI3RKDcysEkCbFeA2OnChhk0EE/w47AChKVophXJ77Pfeoh4Uki984nTNrp
5rW/xp037uMnkioeYY4ahEtnDDO3d7nBn+VGuAlljpOEI1258Rqvlu8NUkd9MC3o
NJKwg8t9GkTBKxNokYyi+2dNO8ucQNL8ogw4PAa0UbQwG3gkNsnY6FrcfmfXO+y6
rzkTyqtC30B54HoFEHQGJzaHOx6JWoLEwwzBIw7bb9zbyv2zuvF5taYQb7nRWMLG
cuhnc+/Wy/Dg352ahx5X6FyZlu3XVqOwybH1a8+iYFqwHN8h2GekX3ndKVUOqbBK
Zexz2L+TgrBnMoiWWeWHsSHH5kFC6aHpHPohlp5l7aAPa2HUxhIsEJ7d9A7ScER/
zF5N2tn2W++n8FGL0S6ZlRs2HGnf+TByXVaKGfwcWcXlN5/BZlaTlpD+XAQszq5e
OpsEskC5Ibq8P/+RYeVvmkSpIbkaPUniyyxPs2IXGEDU8HzeNlURUrKKgrW4032q
nheqC82YqmJFY1e0pn6kqBdmyGDvB/rizjdU8K+RV8qnJIvCpaZ1GXuBhJFpS3/O
l+ZXsrmBP0Z7Wf8aebuWrehhQ21ozcH3xh/T3sIJW02Hj+VFLWOVBHUPePEHGfrV
4D6z62vzoCdV3VXFMtsd0+iIO8i4cjhxUny9jFn8w0StvMt3aWCrvy2GGgmdlZo1
JKezNq9+p0wdRWQfis97UcFb1LqYkb0MnglpTR7EWn65KCA0y2caoagDH0kLowVD
s3g0Dn/GkwN08gAMpa0x5I/1s2MkhWnDGfZqwi+ZHsu1vWFJiF5wwiTZ52CIm+lZ
Y7tecc22dgnyJ3f4iu1uWPhf1GUs2rT7/LcpUTfWJHwPZBtgoS/7cqCFogjkaJXd
wONxOFXa7la42xV0zZ6tntfAEdh/ATTQiFnOvmCvTptuQLOwfI2T/27K8c0UQ9e8
Dp70+80AwB2+fQiXRiI5QSptV6kTZrcI5d3SKO3FeIKpenCHFgS1TSXB8CzXLVTC
+pDHn/48j8qSy7fGIzG0y8qUk1zZJBfV410ZqK9xMRqepYMXoxoUhU1TlCNLfJGE
MPK2Q35+mvj2oxbp15PngiTA0tSu6v61xIKiKfoKvyMvfmqM1HJBFZTSieWI7k8U
Vdw8h8XxI/aZQ0d01j4/KaUFcjLQsi6/xXDnQYXNOKcnK4S1K0mxHivT3wqJ9oya
kNAlZLSxhbhsdiZ4uHBvqnDQdVhjOwy2WbD3HiiGRCZf/rEmHFZID8yfLxBFn044
3w2lOL2ySzOoPb6XPUHEFtxd6tSUq9E29VDZcOUg8MpxhZ7NS92rTMEoLWZgstMg
c5tRm+OB10Z5EhZha1qfNeQEGNj5q3tL1mRgvEnheX6HcAiM3LpPAF8UULUlQcUj
zI+n6rHhtSQKMBQbzX5VIz5CcNRounM8WLYarQNx5/ENWCCOdL/zB2eRvuZlNnU8
TEThWB3wa0FeXFMcwGNC1jlDvOTUxZ6vmobgNYpk5mEJQ9ialNgwiBH4KbO5g/Zh
bueYKOlfXa7wP0GioQXUpENRPhnlFu269CGNRj4aJ6uvCwgTbZazMB0jxVK9Qx0/
xK9bRRHYIHLqP5HVpVBA0yNy1BndfeUY5EqpflRx27Joo0tp0QEMDstMhpIPq6hU
97rIbHZLnPQZEe4P5icTavakMt9jubsbOft57rehk3QUNWMjAvjupyoGSf+0JqqG
1OgArwhTGZTDymAEFhJWEcYQ5rd7DcIDXhyq1TfIWl8qSm+1PR29zbj1FNW2nCrO
E6+CGRGptMxE2qax3cclhC0nzToPqNZZsPs3SNqgRxjudpxqRVuQW8IOie0+SZ9+
7C1EVI9ZxAt8alVzC4ZwMSnj7z/liPjiUPQxi5EArtfv+mwtOuFSs7UA/illcId4
sKI5T8netcecVIbHuwqVzgZulZZqbPv9cFHHIb7wDjtAU8EfnE0dVnJN6bkd5zXB
oafZTQ468ZjHg6QOK98jT0ob3+LsHUKrky1ZEcx7lZfiCUBdvjqIdirB0i0cXaM9
CXxEfCbJYHJVPxRgxZHPhAg1FkYeIQS3uDHkbqzLlqAWdqpdPrLPOawRKjdm3qVG
XyAFC9jKkUG1jIeiB13jFDAGJbg2Ss/tx2E6sFgPky2zMCE3dWjwg37uSAKnYKg7
l5opVVdXVe0mce+ANvDo0UskfIzlQfxY85KTCp6w2QIEX6PtV2UoArAYA82DxQWU
CSWTKgPAxge7popX+CX1aQyVaY48bQxNZMkVm+z+d8Jeb6Xs0SXnP5ze9z5o78xO
+UtAced8qNGkh5W+OPRpxab4KTEfhK6xaC0MT11fNmV3bRr9IX3jdhrOszJ1PUxU
Jcfoxw9fugWQniqhdE4H+vxPdN4plgvU0o17qc5mDqnZ/6Xujkt9w5+nvW+cGSYR
R34pRSD4IsUy2xWtoL52FBC9Aho3NcxB0x0nNQ5fIZIoaTeVAahTvWl472HySR2H
Wddcbw6ORdCpHWptFRsLOO0GZPzAZ80gfu+hv4HBkk4g8wBXDJ7pYDfH72ibutlx
i9hQ/brpfPAG8vi0LSSFmAkMuy7RRllqaC7GSc6cdbiUZDaGC5pHWRGYFjVAG/3W
h4FP5QNUlEn7J6Fb+3EGGrYjx7U0gaSLPtx150AM8u4rEuI5B33flx8ASZX3bzs5
BYKYdrngj+2cJk8Q7SU3Y7bsz8bmVWB1YvblO9cRwHIEAl/ZyWCU5MH24g8AK+pb
vhYSdljecqXSxng/LQDnRKsVhYBJSWtRjW6YgPFeZDT/YrlVdlWitQ2zqz0xo9xj
N0AFyO3P38iZ+U6j9nJhauntqtK5KgicHmKAKgOISfMXmRx3jFVyJbfb2ziBpeDL
qEatVnNfj/qrjqT5IMLngyaY606+f3YK+Bg3AR4tD3LiX56CZ/DNSHLUHWEVPYKZ
CV26ytEa+PX9rbdOZTaKVeiAZ2WxJ++r0EB9O4AscibOgC50Pxq/oK7nLV193tMm
ZaVA4CgtuoRz2n3UWn04eCV9MvoTUwCtm0kOloHX5/6sSTtR04jDStuhkPRrzpYi
7j6Xc6AqJLtbWBYd/YrlJ44gvpx1+9rOrXr0UaReSWgt8e2966D0qcTEkJjBDVec
byiaJyv1JcM4j+cDQ9zK2PRChXE7Kf/V/rfGr2ZjhNxdxeIOkmt24yl08VqAqFSe
7VIzRp58IHNmuF00EhFRN7/AozpTUObqdG49y13FicX1ndDkfHCaekTmCsW7gvQE
tlpDkcl1CqCdmN3ZcqwixZNOQUm40/f3F8GpYOQeyieirxR2KwkZX7msB9llJ1dC
yDr5oQuaasshrJLAehgzLeOILQz5h+DImupREtqO/KvYPJxedV2m8cDQ+ByULDrH
yc4d9MvhxFWk9lIWYhDAFrUER3FZ2uIcHRhSdQ6WVHWEZusRN8q63h3rUMJR2GnF
3sog63X+9D7I16qRa+cWV4nuettMPaGWg7CgCigxT/boYQLx12cFzERve1hVKRbh
yzzlEmn9TwPcz8tyHlsQnaXLLBQ5sXSJothUCPP/V4cafD57Q6Kd0ZukE4AcWkBM
OpZwILbfQOzyIP4ZMRN7CdQoMiITx5N8zSYI+GFdkYEAN2ee1BRrscZsO9+qDotc
q3FPjQEWEi933JGPgEz8h8Au4+7zQtPZzhr+5Ob4rVSRP3DysUALHayWf2plr4L/
aXm+5eyIQTkJklhnFcBAxmDK86SYcz0FkwYqteqWLcKG+Faa8n45uvFM3guWnAZL
RL482ws44n40233JKZP1yb0fnYMeFpvOprWOig7mpJAIpkbHlwjNjZ/z44CkAc5X
l8vHUwZkhIjAb/QduCw/1pzqU0TQ4fV7W8UZOtNlUn5DxljMC9O5KHYHuUwpSY/M
NnP3oQRojDLpnqysL/kk5eYzTMEBv6aULrUXXVjuvBBs5HBI3lXxpvg1XiVg3Bov
vt+cMlD+nsXq+bnfcmxeVJ+kxAaptYpeqtYIQ+GlhEXvqLlb67e+ZYSUi6eJ0vhh
mWp0CnE6LhCLa8zAmdumY7EJ274BtZyFsg6PKXxyVsSH4WmKlBg2Eg3ZIqLCET6a
38oxT5THrDZG1RoYpSlr7KBHrJ7eVCw+iAfRrkChRUSELuPI3kYJRmf9uB+R2umI
Yb0oe5EP6zynbcuFYJjSHxO3mnHK1xoxfvxpshzur+WR+76G1LL4P3vrDfalwlQc
jJHsqMRg1sAod/ANlhr9gf+GfdaAznlawE6JoW0F8tHAPBeeZklSqb1Sn+Ro7Npm
pDCnAj21x2JYSw6hwHvsUbnklfFhaLX7MjN0LAhImbPT2cKA11V3KiZ4edzbbDS0
SpjnzybGpO8oL+BfZ38CrUcO9dIyDJFshJLt9qiLdBgToQmlylCIB4aIpFI43WHL
86zOnuw+9YfMqEIEIlsFcmw+YVJce7rFb4dsWPWnFLzEiPL3VuT6ODjujsnRgFwV
`pragma protect end_protected
