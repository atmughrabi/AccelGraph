// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iMWfU61DPHZK59+qNY0vjMLgoajO94jVJnUCsHWspQ9F3nZatgqIRtO+uNtoSG4i
255qtcnWcH9nweR7md6Agt7kiMu2Q2gM++W0VnNSv/8kTBq/ZRieZDcz6YhV3d4j
j4IwRC6tfKqTj01KxjSFpgsKkxRkYf8Ia3K3ORb+rWI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8288)
ynK/jOddIZobjLWHmqurxvRqaLs/1s7gKkkQkpCriR++mgWS58vAIDCXvPZMovm9
lrTAqyWmMiKsrKpr4zlvSQCLUlxNSHLJb8zKYlxFoFscGu57vLSfuhWaAq0ZAbFA
4JhrhVQ61pxbIzaZLTvIgZoWHfm53C3WOrmAGwBoYG36yD7kU7wYhjTydaviGo/Y
YGz6Z3pyvxKxHY6xphuXbl+lBrpkg0+He05g3/PDKsJGRjp5HLQQBGbQngR65kjL
Yfc10mVOXeRGV57BtVIjRimREgNkGbfeWo+EEDEBSjA/ywsxouzXmD8t80FlY3U9
lKlRxL+IheaM/3RYsODBXa8Oc1Rv46y3qiMtu5SVgItHXPE5ZsNumZX3UVyzCfeC
TDx3aYHGS5Msct9ObDG+G+H3GRKXkG5r060DgZkAQZMS8QtLlfVIM84mOjXydqG1
qjCmB/YgLroQsuFkCG6InF+g8Vw975VDlOZJTY9XgRJzP1uPYAlXCqGkErEHfa3C
W63kpegbRzPCkRS9EL7onDIj2GOlNKJaVJrURuubIWzfT21aTBYkHqvn7tgXuF5K
dIZfkOqpsm9SRQMg/riS9XO+EvUHsqnKqn4CATpVlGbQRrVVeviWNYuQoqu4wnuJ
bzrvMK6bfM4R8Ltt8sLCTnTIC6rq3fGE0R1sKpjhN5ab8z+Dum2T9AIJiozj7oO1
CbBVf7ny5I3vZXtRkdKiXErGIlL/Z6RnbCGgfO4QGix1qXjqsN9bDEeVzu5GHI1l
mHF3wiugExCRC/aIyOAWgQjHVe3Qm4Jt1JCssMPi8c+OJxm/4jMwXxo9UtvNWj0G
lw8dlrXoR/q0wzELJ36S2gsmjk5EYg1kG749wlRKjkDT3ucSIzVfInYJyZlRYiQN
PPPqr0dMVCtLh5DDgBStq2QGLlgAicFh6S0TBvgHvbtHL+9v57Xo2aTnaeULO4PI
oboxMq/6yd2Rld/dO/awYMg1cj0eg7sfHN7mZqpEwDjwDyH2PiLGpdnlKyAdIW+j
KBbMki4Nfo7xSO81197WrEo0hpv4nMvpoZxvBYcuZZnJ/Re75Q2KIGzBEb8tZnfC
deqYbXmuClx6bUGjKLIetHJE/GaH6oEeraGmTGYk9uiIXQf3K89FPU3GFc+DTzc/
eXEY/Gq6/PQ+S4KuY8YvRRsZU7KorJ6pqzvljO8vFdfycgiqW4t1Qm47VT875Pwi
2qPGSJivQ4q1e+TcGOoP2zBYuZyLDpJOW2jI3Lq/d6PqYdjcN+IDE/Q8fGoIXU3u
djd4ZFSX+Jh8wukhYidjaZelsgCnb683n4j916DZN01a1mdDlTb6Eo48OGnx7rAW
QejoSAQp+jzg0rJ0s04MulM6Hk/2kAe6+LbnSDNR58PLUikoFf8onSphUh9ck8ox
XavaVz4SeRMwBx2N9ZVCa7YUfc/9UKtAkqaBhbAKFRth82a3EGNTiZhodX1pThPE
Ib/6W/5aS0aFzdV/OFJDQLb8ebNQds6LyEsSVZxrqcnu0RehM2LCJ3ZLAVEeGOoD
p9M5aRXNQtvlD0OtzIPq4FtZ6WUI9p86ZViCq5HUJ11e+bxf1urC12WOfg/yPJgY
XM6crCfrIJF8p6mSqCb+5AL9qNRdQDPzAmyoNQj3pTrt3sdH5QL3dPUFZkoxkjYn
9wZ03vOpApgNboJI+mLa7thLSaTbIam8b7llmGo8DnUULylCjQC3VGZ9s/qbN1rP
H2BfgirsBXw0DUyYimZSXx+vhnsVKX2+tWGtCUgZMLy04LjOpO1UgdElv9o/+bj/
LuLG8MHxdlUwfxYIp2+4yqqy3QyStwC0jDZU7I/1hrrVKi4yQ+KCP9agEU1l5ZQN
nO2Gp57jeNd4fFqNFc8DRTgK9Fd5uyPkH65LuicSb8cTVXy/Z2JPwDb7jY6FKdaN
SWfAFVbjv1l/1bPJWTNMpA7922o9XRQJgJCwFku/FYHJtl3RQgkZgCNfLofUPgne
BodpqIYVKZJx2Dfpss9m6aUbN9Aulqoth7LGHViBcL71QssHDK/0lC9UO05YDF04
SXiDO2VkNwvHFIXsSGj2U6K6Z0VbuxtTBS15paD/LdiXo5FqDCOGyQYyFpvtCQH0
XOoETTLp8dvV0N8oaW1wB2nAahLi8RTqFf5MLu6GUclkP9thvIBIAca3a4U9Iv58
9d5N5z/Rh0MS2MjMFuzWnxLm0ySaVP+QWOEdhdtYf8XgMnA+elzmzneO7pXoxSkr
w9edQeiKvNPyaCmf46psIcF9zTGv3HPixqjrBDydLkjQsdoxl/PVqoiSCR7uInoR
LFUFS7JyisEMOnNFhNBsSPB2mYw5KYfL9RtCsLqtCqmubPVjh3q+ueyPGbwSR9BH
Qu4jRgthHJZmyHJsbOXwD+hspz1YUQVtWDu2ButaMjiXUQev8bDEHB3L8vChLQ+2
wqB58ku9V1wkFVKUgK/CdLGHidLb+42NgLlc4FoIeHArA+Bo+y+TgYkHkdqTUBNV
lNLnBLtlqLfsPx2fzJsbBuk0ffgFRfc9zDAq1u//sKGZOHZw1xwJhz9KLQZWrOnz
IfUuFeWzfhxXItypiXJRptS/unfKK+ESSp9qx1ZMrM8NB6CI/t0W0bOb7ZRwQg5u
CB/G33e4PcEM5CHAQVT6A7XK+5s8fHN/hA3n13+cYxAbnmixyCdyTkXQ8ndgt+My
JP9nXLmWAgC+pEThVZYrDHLwqCljZCM/V1dHANpByf0jTUYkMfhbVDrTn0o/yeu7
HeCKHauG8SpGaiFAyYvVnFT4xQLOIfSxdVcBs1mUDDZ3JcHeoRIFIiaUkN9IzEcU
EzQTTN93KvqPgH8P8MSm+kc3obWOAw0wiWXX1fE5dxseOyFd38/ua1fm6rSMrcwD
69dApebQz7h9JbRWN5TucFYv13Kuqx5Iy0iZj6kawH5eVkUdWaiL/j0lXA6nLkGq
nftBqhFG4/1gSUcav5BlOvzq/T9joduS8s/tatoU5hkqcqX4lNQ3nRgF3HCCrNLi
lRpzYFMsIcfsPtgiIdsF9uceorsHKphmZRc6IUE6lFX0g9LyWVs0N42J5WGr5UE3
JzofQLAUHjY8VFOn+j136YGmhCPEnJh1y+QVVQnPqKqqgZik0XdmVixZN8MFvOcN
2MepFwZyeyljoYwxNvWalz23DUSSf9n3LCgDsA4xWNJzGddpxf+rs9e+tCJjgtNR
id2FOBBUIrB8m+dYDabOOTmrA9FVHxGndCECT+2QPL5ufjJYb06H6vHL+8WbDn0b
tkuhrTuWvLRDALLfAdfi6TLoumCXmJENea1D5ZRkbQTMQdCKx8lGfkQxYkQSwQgl
Dm4dAI14MfKX6YK8xfcAYCZI9ZT7GMnmdygeE52iQeToisJxBGoZdnRGY4V9h/Vb
aCfxw4G1QLlOqPy2uGYJufw34IglhspT+FuvDMUFK21yXqFmHl0R3f1QFgk2POFU
rDAyt6uWgTmrsEiyG2spjE4Mdb0UWjI7GySbIo1PIo4IIApBuzirqXUEOS7HEfcU
VkglCn53C7FcjTUrhaGOfqX3f3umkHudLjQPf7Ncp3dSUJWngl9FEqjkJaPgBPrn
TflyPBLGr647kDY8+/yJ0lOZIZIsFvZCblgp6FS6/U5POF9r4OSUJyse4bvFzc9H
GEDPGRRRr9N1ub8cgWSNRCLqnK9r3h/JG4Dde/UOHfHPieGQldxKFkyeZ3ZrSWBw
F+IM5GMFUwL5Dcaqbo8tcQDMtKs1O7Xi1EVdw1QPuiUCVjGEfneLj2C/409wrzQC
bGfj2ba4pW0HXAeozSh0H8WR+tsFm7wFHw4s7IB100txPNocmjdYO6fyEdrG9QA8
JYPcsUbMSbGjEg62gsVfuplq4Lcgh2Hwc59uoaTl/q1LGfcoKCcjKJEe3vY5RiK0
RGcIJ6a7QWK6g4FsOlwt8njbo67G0MKXQpPOdK4vjwPyCin33nm+Dr5/8FptS6VY
e6ZiOfC2qMa+fRsUbBRcbrFLQU+BLS2wcMqVjqHcodqf3WtCATWXTCVjQ5VH16ip
sOUQ8Dgys27BRAZ5affMX2f45xCmehIu6jt6v6vwmTMn6mJq23NeXxE2pSpYaNB8
3OGA0vGL16Q9+SYJhVCKx18zll2LMsuwPtBD74TVqe3l06jiX1J1k9DcggN5IVZC
QwfevKAf9P13HsW12r3eDRY4NuKkhM2+a+Y05/rj4eCUwLLS6jFyq8H2K+6paq9b
wV0/MxcGK6d1B+rMLd3DZQD4EToTC768YyVaPKGYjjGjEWEnjvj4nSOcFwOk7hGj
ZC/ZOt3gO/g7IZJ0FIcYELj9PCFwCOk3/4BNId/OYPzLUu/yA7rEgpu5eGCSRkZr
0UgKQKICFpeej+JutmF4JV/qgL2RBJLlQRIViMgPvpN8/q2Wmb2XzEe/TcKFYOGy
kGSir8a/0aw6mvTVLkxe+5NIiu/6VZGWLOnOAigHNJm1Vb+AotOiEGLbbtUBxbvG
uk7JuVT0SHk7u/xG5iQmNSX2Drc9jgpabvFvHlZ892HriXr0vaULLfv3GqVSo5jE
pejfEMOlVuEJS9cKNppVmIJk7CyFRjXKlY840HpDNW8KebcjIZwI4Y+vjbHyBmIt
8GheuAu66tuE+G2md5/piOwjZRXeAo0+jjw/uHOm/nZtChwuCOZ+ki3uP3gr57R1
zeg5RaDJYZosmWCItC8uuipU/uT4RmBoQ3w1MxqIGfMDIg9BJEinjT07xYsy7xqM
OYXvOkvDesf09Qudz0U4RGbMypqoUR/TgtmUqu/kaKs8Bec3uVFGnqh1byY8wQn0
p4eOyDOrkR/gvTLbiMU4e7q6OKKdsED7XSzmgqT959jl8c58CMhtldjmLH23NuB3
1eJd6zFoDY9dIDIG/860lGwPHUVeN3lfCJS/vmieOr53r9vC9EvLf2QDZFcRUyA/
wwnHog8Cpnqs3XPHt5yTKEb180vvkNZUaa2vc8t2cXcEuxTO9Pts88KhhP7rE2Ha
cfgQ6QFCTju8i/x8wIzTAw+2rJkZKk16t0cEhELdcqWlrQ6APY/aA9zn7BypEE3I
ghT7Sdyx4jzHsFKnRIkLyD6QA6vdLvB70ZIpjOnLOi/J1ig7hsvr04/CJO+h1CJr
1pZ/pdnLkv9wOjdz5YXQFNVx7hEMp4RhFbz8b5l5c2tn0H3LnvqeiAc0u8tfh3gq
NqMWkIl0hAL9WPIewC0GWhUfQTxVGtO6ye6FcX535utGHj77AKbpp+fr/M4UOyLx
04gDVzhrtEnEGn+XDwlhVAXUhi8HwpKbh2wD46c1OLrlfoiQb+D872UgUvvCQn0P
AKh/TGQVf134hG0i+utSSNKD3r4U8fpbbGQw2Gdddr86gAivABYH0rJ6d8ZA0eKI
/LW/aQTQJIJJQJkmb9DXdD9eYX/A/RRM8IC5ac6Gr3ETrwZHJkQRg6YWql6hoxRh
J6uc9O5n+Qjt4r+ySpJGaWqv/vCQs3Ba049iMnrzTA1YeGB3yyzrHHESMKAX0Ecf
izNXOJYgUFGfeTacv311qI0V46ZUY7qmqPfrey9APDcAW5fh2o3aVtb14x1e3Txu
yrpHpfbvoc4b3ZN1Kx1E38tnmfhBnQbGtt4OURBtow8q33LrMQ4qamVtaypxJQJP
1CikGeLLgJdpRLErOI4+C3jqOTCHZnc3/QBvHrLnMLPio73trAXFJVJESVIIA8js
L61Lb2OBeHsTewihO7PrXrwe5zaH+XJZ1eBdgM/rTy30ZutPt2qgA1bkwj7o2ItG
g4IsNC+UotBaHNPvKaN5aGgufKV87R7tFYPLkH9QwYIxAFWWTG4tC/Or8vQfogpU
DWudXXOb2uhbEW1BspNXaO41nkFEbvC68eD8vadD3V8Bl9qLhCcnu/gvbXnZoKeu
OUF3I88Jfak5zjk8bAAOZq1n0rf72UEcxui21o9qkRJLdCBs7v81bLv64uwftN/W
S2C0ZKfK8Hrt/x2hlVvhhEhEyOtf28EhDUWLu4twGiDIcjlaLO6TN+P5VKlNkr+i
oxHknZcZkkig9vBxtuFEbJcFoie3BLFXjAyy6YL/tZrbCUMXLg0AoNfCap7VSfQb
Nlp2slVeza4JuN2qX2WGfdB3b0JnhHhTNfnFmO5k8Y6TqAPQ1JpK8VL8/l1oT3Nb
3p0lHnR5cec+sfvVK6QLV7/9b8PggDjSw3KIXt8oXuzDxQYTNJHxPZZUkgiryLNA
KMa3bii3Nk3b7zrZ3MpytPXFL+OXAiQnxbP5r79IMWqBcLgztQ/K9cCE6Ryj24tD
X8HlwONsQuesfkgYIN+jOCE6tC2Uc4MHoKV0Or/6D57qgkW0YUtRGREzYB3mBzEu
tGrbwbOK8uNYgnmDliKj4F1KXfKIPFdSF+fFsZGrsIQDB5VSzCZTD9vWk8c/HxR9
KlimPJrl2agEkrXL47yAKAcKRBHdPPlKLU72BQzfcU8wOSpNzLVIpxv5HG/JqGl3
cCHaE21i7cJC448Yh1Dyv9nuij4yJuXCb8/mFY8vANAYkU3EPYG9PYOYRNHkwUQs
ukVzDnUlJ2Aop3Yhk6sxrVyPM1eEmODAtf6VAWeZncFh2RaJx9M1iOsF05BboybQ
w0p3gkUAAvuxa7370dMYh/l4n2Q4f6C9ZedrDQMg8HK20UJq4Bb8r5aSES4QTtUw
c20fA13Sb0AkTFDB11sHE9qP+H0KmOH7BHVQJpit9TcQHbPTYLO6yGBsgRhSeueH
9iVsV6LBK6uRzfKf/nIhVji0nAJGx9W14znQ1/SR1lZ475OtEa5BVRNfeslsxXsu
GlUuqshGGh2sD8xmfn0YSpK3jVhcG66FcvmQXoCKE/3g8+JvWxQfJXYP7/bARr1G
QMM9sQC//KS03oMhBHa1GqkZk7NWfxs9xqGzMzrBaS4w5iy1DE+2vndmSF6aBoWB
SZL1meZ49kPl1zR1VNLZm3B2ghrhOdlFTBZzJyV7UmBl0RiehN2DF3zyuLmOuDoV
NZkFBvzE6ugJ8wLHAfAbRK8VKtzKlG3udEcv0YTpmnebVqgsr/tyhaIAEjYV9HUN
Wbp3Xs19OEIaq7sTmK0wuszt/Y+ScaQBEwy4F4Cc4x0+dWvQ81Z1AnT0L47IvoVp
h0yY/ADdxr/J9xneQI6SnW2NFprQGmcy5l9L1tUFTVUrp4iaBvudChcm83LzC6ko
PacFouQ/JXM1brWSNqRT91NoyjBFC53peAQIDVahy2D3ZF06FgvrSJdvZ4DMCcmM
azKuqONE6y2GCTNHoT0mHnQevOHQ0bat8XkoKB8uvc85KRVWa5pc8PDURn50Myo/
2R48anv9EhgSmk3DGY7fbY721/kwfhXh8RWiQShl/cT4ipUVo1yBy31FNxHIsfbQ
vPv2XeUqINmJ8azfNvG/fsJgN0Y4OfOJB1W2cYlgPxiqs+aRPoY4WgV8Tf/uAg6V
MPjw8p2iEs53IamjNNDiJjxB9F8Y49mGNVBDyLnvTA4020RuY/pAPoE335Pfel0F
p/brGctPH0KaAIcezCj1m9RifroKtdgLJH/I1LFQNz76CDfl04ukb/KzqSQvXX0g
PUuHxpTMvVRVFqW+3A596s7g4sRkFa9xJvsyYV5qcC5Yo6hYGAX6glWC8DGnzoSw
EiWvZWUQ+4SvXXBMLaTVLzmzshwQN4rR8nwGpCvMFe2lipFcUdoLHbYzAAi8/oxJ
KPqSuv2K5hkNv5sowbZLXkaTHfMr+BneW/SM2OjY53wRXRTnRj2CjPIrbZzp7ub1
1U+I6Ss4YsqX/fr1rHHC5UnhwgKAwGtFhtc6Ro7E5HhEZDmkggiRK4bzWi/Pce8/
Ee9poP76CarEvAdVpD7NUVXm61rSaCzMZD6Udu9FeTuE0+NV4ZE0O2psQdsYgbeN
S+9AUta4+N4oSwD8QmmneNCKyFGvMQ/pplLdxgZJQOi7Bw1Liqkyron+pNNua+Sh
CEfGa9g51YC+NjuA+rdq0yAL0tzr4vxwhQ+T5aWZpWcZyiYvxdupbpkutIjVUFWE
Y8tPR2hkpvsKB52+8h2J+CX/QsE7P2qRKVAlKPLQQCQ/E/WSEWT36FRWFAp7TTA9
N/CitJsWUbVGaWJcqUx+YeQOAhHR95vCTEHklVSKOyXDad9owTdy0/D30Y5gzXjs
lp7Kl6ri1aPS0RXvziBMaevYsfOnet6rYZguBcaoEQ7UKz5ok09qXbw1X11ZDHyQ
cRDWQKQJQ9pzOiObARjiWNFB92pFr9jsz04Kh3rmHkamIHxRHQ3fHFX4GjD00Siv
wKJ5V+3sBk0mTmOYjV5w3oVrYSqXph+e7wuQ29JtuXpAvNxxo2z3AnykxaKlBDD0
uaSHSwLcpO9P5Zr6YUxlpzcc65Kj5PvXeO3cUtGvdleDVoqiH+b2yf1pdTWhfAwQ
4Y0osuxbao4jlMyOnXM2ZdPtfuEH7FlAkgi95xzJkJcVxqNMAzwn+ZVO0wuJhpBx
hcNJuxUeW9zxDf6Jf5p/jgZq6dyLZLHwxBvxm+Dsel8+R33QS3vRfMEhM+p9Y7zt
9yqvzEha8In7OkJxWDbo2kZnIPq+uIuPqyi55Mc88yab2KpzR2w3f7On4Rx4StNY
C1L5DaPH5PsGnLS9A6OF0mVSZMpe+Aut13I9qDr4NXCgzsvmLmsVidcVWlgiBaJJ
ccOHuQE+j1oik//dKtL+A7y/PZZFV1Lqzitp8h4La4cVmZ+y4mEOY0ytqB9r5ZGZ
7ToohfBYN4Eat+wNRn4ePGNLeG5sAzln6BLGq8zg8e6DZaqUO9V64QiUBo82A1qQ
TxdukG9BTJVuT3BP2a+xWnGI7c8Z50QI6C1jKiCRxpiEg7mHHgDaAFp2BehgPGtW
qvTcKvjDMn7B66irlRdiQr06mwnX4l6PI0jzMpOdbtPRcMbT8vQNrg9bCORck09y
x89mIkM4YHx4PslUg/zU/A+TypYnZpOnp2DqRSOs2mhC2fzEuDzqXmHaWU39eep2
brCrvmKWdn25dx1oEWHIRM6vACf7aEVCUXmtaJG6OwzqYiiZI8sbRvg7udJqEJxT
2KujSQCl+TK6q98LGJyL7H5SmtmLTO4PE/qvas1iznP4DVsf2456c2UWICR+J35L
8jyqLkKXBcMCy7e+AAtCqnroN10wKXUXFXLyu+OEiAFLsBjdw3rT7UHo1ROUAwXr
L6Mm3dxlXEe2t6YzFK5eQR7u4mE15vRpzGxY0gbTwvy2OHXE32EMmytW63evwThs
QLXYJMa3AAY67pjD6Ga35vxWM9kFS/ZUdIqnCrAp+ga3QpZMkwR9mBeRzMA2kjQe
go/pN1SXd62K1oAuvcN33jpNxhXwyvi5YakvT6lEuxgKY6gt7/o8qHmE/d29oZsk
EpU8RloYMXTZw+R1Xwfc4sveJyS3sV8/uU01hv1gQfK7jGXoahPlI0sIz25im5Tn
ElefhEHXyRW37E+kBg/Tnfu647RK51gtq8Skz5zBpXZ+PYCn0kIDpie89HfqmVDl
z4p8oPys1aKbAnMmg/ydXpLn1muAyTpAlmnlhcsMiB7aVuobTJfQStEf3nDxPSGD
IX//YBY2KQGH5pea1lBGbgAZFQlkP8xCUXz0bub/iG+OBmUa2rtUMMODWThUGmtb
mqg/3cjpeuiwWvhrT/7ZUPSksuWzohHqLStufSlOWJldhvh6G3RYbeAaK0VTJqDF
A5RqlqSb0oh7efFWpqrS3iEzzvMuah1I5hfaTt9OS9hUGthtUz/fTNI7ss1p5N/n
hkiymwxoLnTur1w7C+EbwrqibYRETsYziFHG6Zc3AeltNsfcs8TuqjrLQ+Zgk5Ls
ruchi1yrqhep4xW/zEZwrXEnlaRZhML43njisHD8OETwmFodzqWRjsMCOZza3vZI
cGUAh0GOy/b60Ln72+QFU+fKIWrHLNpYjPDEZKy716UFtvETW9z9pun6Apkz1dlU
d/ujtjxhl+eJ0Vdogkd9EVok64oOerqU6pC/yMj+HQcfZckKmcvhscZoDWSdJIJm
f7GGsQH2P4QWac5Y5HVXy8qV9/w1hsNxwJ7j+S/QlmgdWoXG35MYdx+Vq3sEnn6C
mR6I/ZwhP1Bnsf4NHQcoC7Uk4yY7AZTgKiQYK1/VmGBCN3gwE2ahoGdgLCELM8T5
J4elVeF+ODmyakoxB/sJqjzWKIy+9g5uo+U4LNnsheR+Vo5VyjU7Tdg7DVJPUf3j
39GI6F5dOrf0rIoh0cEKeqHfDr40mM7eH7iNsdTRV8J72R0bqSAnnO6bkZQIPjWF
WEFv3SY8BbJcn+7pYOzvHDolngk5Xquu4Dt1ecWehgs+rlpxTiwGXDvAEkngiPbA
1KlIwvm5YbVbwz8dpkn4VLqldu1mZa5hKQdrQqqJxjeKeoFp5DFw+hFTlBgxOfIf
CkbcB5rYb0PCJMEmgzRcIGqOsJAjZDph4EiVgFzP+D+7RSBLx6BMdzdxCAakEmzL
K7/ls5uqBDzwtdZFieEl6SqaZujRl4VNxTax2IyaLezNwTQ/oHtn7nG8WhJFPkHu
qdIdgZBxLVDEIwnw9Zok4J5MAbNTPDCiwaDAP1B7bCsOMXNtCQ92KiUwvZBxJwfZ
voQUxLw0hwvV/dEStP41hD33Guej/MbxumN4JQf6+Yt8uZKZQAtsfAzlpcbxkyJc
3BTR95P27jLdGXkKd9B2NCrmh+lNjJuKcphLVKf8yp6avRBomelUhjJAu30D2sIG
++ei86G5yA/9xCxRLstpAweo0N0r7tPAwe2UXalLHZuiCk7LCiw9FRDrEzAY2htB
ioiYcTYQB8jhV2Eht+ykXf0Trip16B7aiPs273/a2mO0N+lRft3XVB9Wd6ggBzem
41snySMamdSl7MuQPR3KSyYbXQmJyh2U7p7NsBKYtE8SSGQu5DYfM51sZPQea5mB
teDIwlN3DIFF0jpevf3eQacgtOqHOW7fHEX0va3rsfPzYseCHfLdSSB84FE5Noyv
SQkMaU1AXdoGidfvK2oNfMlfuCHB95yi5X+BCqNCPWAdhm2693GLrWkvEY6XLPwQ
ifio2qrJQGqsgrEXBxvVTl2GGDpmyKtjvfRmNRBzoVw=
`pragma protect end_protected
