package CU_PKG;



endpackage