// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SSN8HOf7mAVm7mfQBNVBhK0uhpTREcgWpgIsFNmTOyDFCH8fQ0O7JBCyk1fg30gr
G9569qHhMzxWB3z8zSk3zXHzVewzOegl00KXgEwypYaJ7D3IYye5mabJwkhyWpEE
g05+wpjqhf0vwDV3CYP70FRa6eSyBPRE0D0fvnI8WTY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2240)
bGZnUnfxGix0whPsYUmI9CijeWKd2LYhoZI/zpF5BD2MdDAtK3um8lpD/1ckoilL
WjDbpWiGVbyilyk6p4L+LJRHWA5TZkNz5zKz/t/v5Wo7BFHirSj4NhlktUEABZVT
ZQq8HWlv0FRJmnIguN7c5b+EivU8UcaYNJiEHEGc5tJKr+/9IbM4qFvNE4WZyfOf
3I9fKIR1IKAr59OSgTRaVm89da3wMWTJxxy+z4lN0zF4Fh4RrIJc4dqSnkn+S7iy
QmRoMsU8JZ197OMxTjLB786jKbur3BNj4ZnHLORrvDSgCSsjhfckcDSLjOWv2f+0
eGtOG2oTa+N98k5Q881KUopSNHNUr8uQIsXsU/23Jkum+cERcTPiMbADZAu69Uue
8Q7Nc1DngvbuK+xvYs9ackGPcEtsFTO2I+kdS4wW6kWRgy8igbM0vXme/u5122N+
IZrguiD12ogU7Bjf6EnZqgM8Yj4cbquavwPP71ryf6MbbH2OVBiWAeZvm3Tk2igN
ADG6eb/8AxS+oRQx1ZdH+Qj4gqyuMrygRgD3dQBUQQ4ssqMq36HOYgwMYCJkMHfu
qKou3DDbBBH0KT71EaK/1yefBPXmTOJD6EayprjRVvOqPqf4wPoIuCGVvBEkUBrU
Zsbl04ZAll3MosQ/MhRvLiS82NdC92iS0L58J2R5En5owt5GEUOeoqhBaOlEXNha
k6sdVgvxXxT+rmnCyI4WQB68Q0MpjnPt/PsObReSSHT2Wp/akwbmWMos9iB8+AZ6
x0GjG5UspTBL+zRWUNPenyAy80UUDBPgUpQuMswhMmtpSbntJnOX+wxIHoOwghb7
Kybb8Xn/0ve8sAnEWzMFfemxAJ13DpKLwzXNIzcR13RjviA8RAnw1rAX956nxdUX
i2ONVJMesuQcMAEeSHVAPhInSyqyaKHyr1RFZluxXkkikslRSU4/3NSjOX0KHWV5
qJnAh+jOfsPXL7qzAoVJ0fN9VfqS5ZCrTIpRL6zEdai7u6uVY3P+XUdeePZ4tUqa
4vCQwjmRk/PBU5Vnrc02fX51En7mCD5iIWjWMzNcW4gEHvzbLiguULZ9qrF6sDTr
pDG0/lsAmv7V/1A1r/yIEDoPMyGz8eKXsV1DE4botOM80R1tua+9yMu4WYYffeBb
B/RED1fLjchMx021GGlout/+Ky89vje1WAaMmLiZ81oqvONL3j1bMTcaxn1O2Ftb
6hA7wq72KFTnW/C+eE5yjVAAyzToa/xq01haAJZ5bE1tsFeG/iyaGwwLi5o8M65Y
WGxYDpMYX3LaOYLeqxEpZ6rtS8fmc8cu1JG+NiGcEnagBkkIEadF5RulhBD0Il/5
IG76NAyqhIeKWETtf/950H/T5U2rdTi2XT+dgzcdsRNhsmFIqeAehIofKnfyLOd8
O7NTrp9Y7S0LoGJzKMbvm3UFYs+Zb9qXy9wDR045eq0IrQ1/zaTpCogCbjY+vSyU
piumlMj5ey7eqa35tOX4jbCPJb1621Mjr9QgS+4CJC7nnQOGKP5kH0aB81qp3YUY
Z9881rL6N+g3VSyQ3jayrB5TFuNLuvZg2g0u63zcxT/QYaVtqDZqrHgULu/Udj1X
/uXoNob6JasokUXxQ+ysMCFOgojMNN4T14IOrRJPSPEQmfz/ApJ+0k+nl/fhKeIW
M8fAAvgF0S81Z6QqSnB6sLEujNcKstkRJvhVnoiJNin4StymPuPzWzmymGhz0H6P
4iGD6lAn6BgWa8fS15FHlkM2LERnwHdE5q+T7wMQUR+Tug/J/i9Q+gFNbl6HYLvB
3n+8oqEQmgkpfasBrtxsp2rpoql/56VYQDoK6yTD8rRkFnXzYktPuEwFkMJSLFuo
V1suxdiyzdg33vXqWieiEWWEd/plmkakW/XeyyL76IMmP5Br8UVjl5OLNiqOrOp6
lv3hmVWI2GGpj2eueV2wTI8Qv29wLDxkujGhsjVsrTEb1OP4j0hXBNx+Y7QqDkW+
YJWYaB5KIWlLdSQx7FJ4R5SZQk6c7jLKx8KY7GYIjVoGtm/wMQTiiT/N6NuQDutn
4lWh5+W+NfTIHPZ1+XWBXFPMh7ZNAZX/dVPSOGTM5nN1NrCbqhN4gd6ia4o8o2Ye
NcfgR1V/aOjXk6RqiBlII9LL7hkKyzcqMTYvf0gZ8czwecSkNqyEazdy6io2JCZE
VarRgATHrq7xXraES1yyqT6PnaknVY4OfciM2grH4M1TBd45FdGf96GYvwpA1yUI
ZA4qdcfLgnfxWfEwzw6uS1tPOwqNFNP+cKjSnQzEPh5qzX6PAJPTHvyhGAWpG6+v
Kh0sqKGLPQ0KaJnI1HypqXLTk2kcs/nabjuty6FxSGSceEAPD7kWK0P8TtgdEniT
q+pV/emaWc8LRRpyK+UjHcq2hYw7Guywah9HZmGgjdggw7wSu6LQg3WkBrI16FIU
Q1VK7o3e4kjl/4+w3E4Go04CeICI87VOuxvZJEBV8Pq6ODkrV7tGqSLgMD/6DsCy
1JMmFBDOFVwQw273fVoc5xgVYM5uazP3GvXISvCLVme8Lhp5rRdxALGyOziB1Nx7
sSppqfBUUd5rFGaCnpWS29iyTldechQGidpiclrt8nSxRQiGPzHJ5ic9a2KJz8St
FQLfD8WH7ujIndXYarLj9nvwCcYlNs3cpobNrUylx5aWy/b2DuBSn3dRAYN+Agpe
CtNV93HLQTsd9ZtPuhgYPSSF0kt1Zz6GB6PozVApi16MVg6RTxtIRyujpjdpqqGG
+PhQo7+v9Jdhru7eNd0I+knj7Y1KnJq+q6G1Qz8e3kFj+9OjKuUvCt5sWebWkUxr
Z1F+y+LZqDx0pUM85UuEyLnnJyTYNPNfupr79e6OjH49QhaITKW4psRgVWb2iPkG
4XoaJST9MrvXix01LsOgZ8MJd85ciIIIJX+HRU8dNemFmLuVUnhXyB6Y/EGPZsdz
J5xQDgLO8sI3HRM0Moh9q/nl0CW2uVyugERoYsiYWqs=
`pragma protect end_protected
