// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WcbaAQrHZ32ie9QEoez1yfNB9fhtI/4CcjGyg/xvaLo8g7FXWSDWhIzJ3TSXdLeq
ZB04+LP0lz5vcabfJPx7/mptb9h2ATAFqBtz+S5et+wZ62e0C8YPNsDSgySMjGKL
b9eHM2HKClb1dmIdD0Dt1spVgWAAAAGmccU7uljLsvE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 45664)
BGFPi+ZIzh+G02ZZm3uLYZSP0HjYKfGW7PTGrOhW2e2Pr15SSo3LeoXYa9q5D5cB
e95ZZdQ9peCY8QCzUM41IH6vcoJQcVeeO08a1JuTsSqMlcCITLY/ITvagxLJ4u/6
DAFtVkob+i/umd20h5xLP9Pr4z3SK95RAInA2nmbzqOMrgECFBIxzX+RYbwNe9bK
4uA+CQAreVhrpzxh1gMMCk/T6QDVe2ZAUbcbtsO8I1ibTStoOD+FAU7PrWi+bOym
KeQHOteNh2zpzn5mz88vpFIh92UYDvP4eBJ4h79ig2Y9Zis+UZio9QcRXmfBjoeH
zeFto5UTJB2qYX2Nl9Ty68g4ozxYqI9uBSlu8GgFxVYDOagfzl+e2ERDAMmT9xQ8
t6lJC3fgoMf09mnAh7BiNgoaCB5sSy3i848853v/IdBJj8CtMB8VsUkkLkG93Www
pV81I9qB8ngjGxfWCUSNsWNqCo+0RvhVYZQtqN540ENaGazghpSS+EA1mjOMKY6C
EvNryzGvUZDK3GKA2EwVZIy88S/f/04AkBXxBgoM5bpgQtXWjnzYbzN0y/31j5Ez
wz99aeBs5M7y5lW3azj3MSCJYCH04iU1Jy6H6umUzhMTRora10TuypcPP9Zg5jZc
ncThndSyRmSNHWnHFcIjZFlJDGpflDsEpEwM8vaafkePS/Ahq790GctU7ksFsRrD
xSmIp2ZbnnoausdZjC2A02WBGuk6vPJyPdETuovGbLBZWXz4zjTKSvUqXUAsipTS
w7CtPREWiLYFjlVo68mdd5F9vipNO6J+HCPXN29K0HR2DDTPprVELk0kj6MXAPR8
Y1qYVbsqVWHSzO8DXJPpzvxOho4rPZKiHNEzYDLvXPX+Uy+uNWu6U4kdra63i9g/
lj/bq1PbJWrtfMJP5I9bEj2OS+8cShDL70S29USjECiW4RBQbgRsTBALfILjlMdS
zwUar2lQNPvoB63e+Fc5Mj10yUYSCbuih+g1zHKPV8betJ3aro2rqnApHFvbyyCx
RlxDB30SguZrmDxvD/C1OhyjMeWBrtVDyDDNfTXN+glaRNquT31Yekmh17t2pCtK
HH+qW6mxoiIvC0DzYjX7lnD84wyAhwof2tZY2jN30Pa7Y58jArZI8M8Wkwostym0
yIHYGRwIjFgbXFqKZi3KbBwSS1SEPMv/Gm4Nf1sOfmD6gXyG/XqPZDUU/+yYuBjR
Y8IoMHdS9xmFjIxY4t5nEmI2ZkTv6PIJZ+43g+gd43S1Ws/xi+o1CgkUh6nE35hO
Y3++Fj4Z1tGvW0RMCgd37wimOrQc4YqBX2jkwpHV2ork5J3FYrWn22/b5CiLh1ec
IAQINUH6X1V6wvsy039vDoGSIfLSeMs6lYhg8LO6AudzCmk5vKHE8B7CBxEXVmGO
TKfV3Kr2OFf6iUTVE42wH9pFdr1IT4AwuxhYPdkUmBX2r5eX+nv8IYfAi9NZvzn7
upLpHccN1m2hiNd9nycSvj5Ml6LfWDB2to56NxJkXwLAY4h4q/4fueu4Pk0fhzq9
g+Kytq2uC3jmfg1USlsWHh5WSGeBCl3svliCfzd0BPBfH51+Kik4YpLr3iGdOQUv
OLV0SEY1XLV89bnaooz4qhedFuNwyDtv3an0YwEb6YYijNFKYHLbFxNOFV3+kgN0
9fjFiC46tQFc/J2fw6Byj1Yp7zascIstvZXAnjKhGyNALtfgLcJLrhv8cCgG8HVj
xzrjJvmHu1qi5ADwLMn3jCd9ftb9QoWoku2gH1U8hZqtbU7h+4i7ikg3aQrs3GGR
/4HSYOn/jKE8tN/xX4KroP39ogxBGuaUJius7KEjMMGSj7aKtf+u3/3KH0+VODHg
SPWuZ1mltbMBXFdXwjVuwe7BLdhQHGrVzTb2z686HWhFUwuGn43acfdRuoGbMW2Z
CqdMOp0XqWZRHPlSXE804ZnmfhMOmRODN7iEUY2Rtm2Z89YA06IQ8BYbeKr1U+oi
vWNJPuT3FKRvDwqZR3DqCoYDVWkI22KhVTEgSbnyB/o0riK45ipWRNCIIvzQthGi
pv62UqVtt00xnjt17cguFQXqhuUEmL2IzHnHHTN6u0b9toqQXWV17JFzVbMtwc3l
5POmZgRxr1+oTdNFgcgT79eLt58ZiXUvxkWDX+2VFiolvUoJMb2yKnjevUrSS4qw
MEqjFcsoTeqpNyrMB6CV8XtkBVmCctcpU6BmKwLW/1g2b1OK3jb2juVkiwKX9FSt
mci1ZsCTsi96FGZMVaGGAkSj0pWvXVPX6/UIhLz2FkTtlidM+Ilhv55ggUAWwLcb
CExR8LuIaxz/3dBAi5/kGiC2eUOlU6vklvYkgh+2SYbgrUPotBRMutOJ3Q0Nt6rm
zc1cCDAaHJDvz1gHeIK73WhbLaaicuViPBEnW3LeP+Eeac4YNondYdjZ8uD07T+B
0Zz6KiCk8WSvRjRfUHRSATQcC/apEFgme+fyAvOaA4D8igLoI5Kx87foiELvFiwm
+bRQeNZN70pdeBLqmyoxLaw5wZmjtYyYuzTwBWvn8mTMmfYPiNXxB0crKfqPdIHB
bs76hk1BqcF4R+hliCcyxW87iNQbBDsASkTNm4r+H1avVcQLCSptjVukkuplOQD8
HVSVAwjPWxh+k6dENjL8ppo6D5ORiK0ehjfHpXyGMFeOH7YXiHZSgkyCduAoLzCW
UxTPjv6EhI6HGueAov8aufDn0NB6vldX2qoKpPWkyCIe8W8WcEV5Az2jmVWgUCZ5
sWTMhFsr9FbYxXVOpzXzYyFArxl9BngiLmVvEsvQjvJ0kwk8nzQmG5ryc3NpjP5T
b5+0Hq3El6VYGTLdqEKMfL8WNO1mC567eHqS9cVzVQF3p4jhC0sAeguzvkwftUjh
ROcACkPBNX2ChLBocyKiNDCxe+g2NbVEizVrTOHjZUCi8fe3NFJ43JieNkF4Cmgt
/Pg/MIcaebDugHZbmdHn6sRQesNsqS0+FKzmFI6E76NOWmdljqh+LV26vctjJFDg
6UIitLyUHkl7cIlQEhKamWW3mtdenxDuPsxk+NlJlz4Nn46l9zxYKE+vs0XoXwLE
z5jCm7+o8gemFrdlqnXhgY8pBMef+VmbUBLLLr/TkAshzTkZsiPlc1DcpnaYq0EQ
hXLN5yEQKqNpaGbL/JGnQy3I9YuXg685NY5EPgE8PL5erN6ktemIVNxhfUCX+pw0
vtsgRZ41SPjdg9NcH0go51p3Oonpd5iJelihlDZJIqJzcfKulZvXsN3h2E4LotLT
gT3DqaVtyLk8F1cL0bNCKewz6c+uP3uWpEeoC+xQDqJ+5u8ZJn8eR5Szo/ACAiM7
OpBQy4rtZCN3mt+XzwRZyR43+oElVCLckpOKKAj1MxWWVAx5ZsfHVnzDofND1CPy
NZ3kpwdqcX2eujTudf+WowHyiPi6f9EFEVGlYhHI7AaGCPbYz5bGaxu0olqFGdBP
3Frr687MFhPhU/7b6mtXg+fW3CRf6moqI2V/vx3rFRWr0sA0SGdWkJZ77//XryFB
9SBuQtpaJgnZT6Czzae3V2fifEg2AZC6u7SFkuCnUIdj1zaHIzv3icr5lHRHoIXj
HUmmx5vRh2+9YfilzPwqwQ4v6JUcJYGQbMpO8hVKf9vGSPf6aIblMMT34QW1HbHF
2LVH71kD4ID76q6Y+5ooehvvbGK7G4Gle0WxDV/KWprlRJl40UVR6lQZMGaqf4+3
AaXYsDTPcQaZCNlcaSQf1SKj0aILAhGpXyFGHK3mTIZ6dbGjEb0ZA4q9JVURaEwr
o1+QIB/BZ7PODaD50VmiXD9X7gcFqncKPMq7eX/mrluzkCne1Oqd/26ZFTNjF57W
MJDwDZebwNA9Hmmf2a/tFv/jWj5OW6q/27StyR+gZuWQv4JIKC+VfBxCtf6s3Jyt
e8IxlZMOJ2hei9GTznuJlcWpRmioCQ9KY5d+cdH5uzVZ10LGHOf6P11K5AE6ub+e
N5zqbjqf5clSoVK5Xid0rnxDf0XDS7879e0v6/0a4mtiPWrxobQuo/H4suthzIAc
tEZOpF3yy4lr4KNfXfzCLmt4nLr4NfpSz5l0FdCiQ+Vrj4QBkRsUQ4t0171EaLFA
tUEqYnZH0ZcCqaBQrqEUU0Kx4xA3ggWoV9X8HefZufRV3KvcnCEXFnJusco5ABVG
0zacdptSFhVBT271XGjc+sMDLoqaj3eDhdvLzSBkxxo19dzPmLyPfN019kKdfXWi
ftIcXC1DF6Tzg2KR5OsXXgQPAAv7ysM5gV+7QOYKnBzGncUdhgOt7JNXVbTKTsED
cvfPdEHfMVvRp7Ib3rPiXH9qHyDTKfQDY6/3dTObBdprKlBIzKG5KvwiXxbgCrVc
N4XhlbQPHW7hRpGLdfcX79RFG7aB6Nhf3uzpYCXpNW4/dLchLevytnSkWNRFJSJa
YbRLU8ztVlk094Waf3EKkpYcZyBsCV/iNd+6Y1rJBfAbQxNzSS9w7Nij9XdjA6xz
OfWXvGDCFD1offQz/NVthBWZ3nOYqL2Ir/sEDBXibEay6mE+/PvJ33F8pVA/nBcW
w/vyjhLabA5nxu/hlQRWn1Fbntux/0qIZ5Wirr2ZYYxxZmEFiF9i8ISvDmVO9zNQ
CG2cQGhiME8wQ250qvIKBpwUP2EZIaxJUIpOHcaTwtMoxdd3r2YoTjGlgrgJw6JJ
x7/LepunmJOTyHB9uM5MgQsKwzS8G76oVhigXyKx0uiETrqlCSr39MbbOC1uysQ1
SvrdVTXbQQaSuFRbIx0e7NiVegR08f2GB65O5wOo4x+PTo3GvXM8vhCdEli/IgKy
vkK9QqqPXYC8xAQ0L0UXYGwe+7a3rR9ifjMH7uhGdXO5xXCBJrrt3yWsuECnewzu
KFfwSR0AFGxmTAgLGt9zU7MX9+nCgN6TolCKk+RJGS01WGKeXEsM+sKiSFvXRgqH
DFr6eu+p+8F2qcRFJUVQDM6dAAakqioy8vnmrZfb0hNCictFc5OD0dfXhgCn1vSM
x/8G1nqPuBTgRP2wjYhL8KdYwEde914KNzJ4HwkWIds23v7qc3P69GTYTc0MPNlW
INGCXL4DTtv/SifoO9l3DCt2Vxr+160mw2U1mw/fUFDVMQrveqQn+Wzaqfek8rVe
JT8sez3Dzf7/Sc4vz3c7KOGMVEQgKqhFEuXg5ga66MnoCV4M4B9ZmfYnBYPP5LSL
mcvi2gQDAR72urnC4ln+eSR5XsH1BhyCCDL6awZXWlj1NaKS0vVeTOoxQlqysZFc
BiVCfCXXbjy508l75bGKgd1Ol0IaNXfTrhxTy2/gkx/ugKNQ6qrSzXzb6oOlJ1f0
QJV1h4YhG83T87I4k3a/0X9QOSxy3nT14mqsoTqX8F12Ub8BuX2X1ol0Vhrbxi5n
mxrg6m2wt/8GjZX8jJj+HUge/MD6iZEWogjcrdWLr0VZRRSt5/EucCgjFf4PKn/t
V1TTO9Fw3TJVqATcjNlGyTvH+Qtma+lI1XsuxYQ50putiDsVv70CnZl3x2KohcDm
oyS5wP+XiFrutEC+S0+LFJySXHG3fgQf8MckGD347NytxT7CEA5vxSuXqtKJDQxn
+DqE+5vMYEoxmSsS2pjkFhdHgMg6H82lMH+F7psZ3IvxrXnA419GHYy2w1dU4boe
1GaxdwwGQtgCo8h5GoQSMGVuUlh/DM3kUQCgcK722urUmyKq0VCnGy5xEwXeOQun
/7BIPv993cUNmTSYTYPLZv+x9rAHJ4kmr45WfkW8WR6nH6cNKC3CRIYwAdatt1Dg
1pcMVolaLl8k0FgfVOvLAb465WOKcXoT7x0aIE96R+Y0lW9oPWlhrHwlDbfvl2Xs
x8Xiu6plpp+t2VaQCXKXczvTg5jl8ZyPFCqd44xlGWqgDWFuQwN/MBfFP2iXhf4U
cvHVfk9OnmF+deOpL+l1zWchz8wM5PYGtiZ3d2p5TEXZpwzVOGlOUFHhDXYmUrul
21i8a6J28+dtRreGmbK6W3MhrDrBKXiSq8CPrcp1WoZmzWVs8wmUiXN23dCpaEFp
0VgLsfXr0qsQy6wKBXh6vY5S7SrxlFQBHDmr2779ZwPbBWCWv7tKWXCU7+te0BhI
6lqcTV0pDBA4sjuxjIYIoOfL+Irei7Nkk3r3+tsjk2QxyD/Gfp5SaTavzMi8jDfe
5wjf5PLRwLbOGfKF8WwpsMG/gxTx+ctQDx7E656ADjurfhP5JnuU0ELTMFKi6sw5
ud991Irnl9ehbkcbIKSIDL0FXUzAO2DH4Em+VyS0douQuSLt7KoEZ94NYAslbkH4
pl+Kh8BneUWv/YL00tZug4FZQVfdgZfGZjWl0ysQqqtlnyoTtFPLN8dgIthAXSME
9nQ44W2IJCfdQo26L/huuLD3g5PtLiOb3hIyNYfuuEXHNmEl39rtrHJnyRbceP56
5AkZPf6eWKBxmlIf4a2tkDnbrvAET8VxmbuBhZXWjaFKLoiDdj+jEXtfZyoypBYU
X0GRAgLClYav+AkdjSQuOCqknKnRWbXHheCnvr4eHIK3TwAv7KQQCvAmxcGQtJhy
SL8w4M4v1uXbqC+DDpb/nLydEtPuRd/1CYG6OWXaQ8FW3lCoy/tMxz335fq8PNIJ
Ib7vqAAaD7emyribIWGp1w5UTG+tgLajWB7W3cQoyeO6Jah/prvSfH72UNrFCg0H
y4dXdVNHZDnx1jofD8vL/xtZr/2zgG886/fhH1zUMGUIJjkRl8Glh/QcfLRM6eC5
sg/SH+BI3WXJUEuWKstiDyazoH3mQYDtTt3HLeSjTTMXnr0zqhRlSXm/Q1vxU7Od
PPSBCoMyLGDVL6r2WAm14noE+HXHmj6jN5zA2B5FtZLNooYHYSe3e+6Waz+z/5gr
YoQihq1rMIVkakJPN4PqakcWm0vcEyHtH+sEm9BKCu0rY+aa6j9IDOF5rszs6n8G
QO1VKlkMLmkIdKz2Lk169qzA5dvQz35G448IDXdqe1joE0M2FIMyL0OMrdwjn0bl
7OB+awEquj60VzNFsGDmhX2tnpTdFNGNNAnBT2fTTMWnTJt4ieHHaiXy5c8YItZO
bexFmrXzZQEMNAyeuZ28uq5cTnWpmbqTUSodiWl+cd350/Vf4tHLd6l72zEdR1P1
8Cjpdwo4SPxvz6KCD1CcFARy0UlJd1WHUPf7l6+45ei2V4sWNTTQG5zz50bm8Bqt
dhsnEoaFn843k1iprkEdO2MK5g1jeC0RkufRZcqP5ohvXxUojMraG4ln9r+AHFq2
z9MSlWV1GXiXXl/vSd5bSwFcV3IYLuLpnh5KfnyQtZiVBdGSBOSJsalgiu0/wG1L
qRV1FdfbPl2xZ4wCppEFSvIi7urvFPmMXZQC5ReCpfeESABmjSQqu88M02RWguRg
tLaJwwZ5y5axWtr57domDq+tsW/k43EflrP9B8D3XKF9TqHWFtV2+/xywbVuraRd
GGU+JJAckCgi6WX69g5c8Oa8gAv2K3r8m9v2gHBhXIOdxFZinmHluNNp0us7w3s5
IlLZaQkUEMUoaI92k+kfTrKW17O8J/K/GMf+BUeQqF2oUECFyXz2jaCio3LAk2Mg
46IxHxLNnDBlgphCpFesZxKydRhLgWUqIoRv/YEM2/a4Mop7q8WIRQHnpTKomrK6
mjlteg7QOtaaUD4X8UQ6XAPPRmz7P1tQF+KojVsQg59aIx5LgLRXXap9ZxVZPzRK
GfAiHKQDYFrtQB6iZSzU0uq+wQoSKpPa2DDzYyCJOmEsKKmRc+HlMb1FOnsFKm0I
uxNsRbL1P4b37yxFuQeO0C0CGHMnHlH+l0El4D49vJjKM2bBlh+WHwDF/gHZC82l
7CQyTeQ5TJ7wsDwFwD/BoYj2U0165sAemPdON4WaW3MmgBO3zAsNCVyjjD6Or1Wi
Q3K0k6CcL3pCu+7tvkRzyfzWE4WReUPzIiyGXlrUOova+Wl0wP8cdKayUkIkWZFS
3xYpkKoeYTBFV1atpWApkiNNYrneJut7wrQSexXmD66/+WnxYf4FTgxL2y8q4sIC
hdHWmmW8mbJ++iaTzE9vWmTn5xBN5aK4kGpBjuelkPd7rBpvkHLaLpoAbjCm9tgR
7O6qtN3vAOKdHB1Wq4oG+5LMzJlWaoZ+thCN0S+bFyfwAhvop3O0J9w0Vwd2axOO
prSgCxDFdZWu3YZ2myyBe7uM5+G2V8QaBjHUzZnWrY1Qyrx2sojaFCWA5UP3XrH6
iwywgwg/JaQi1vuTi+6jhlXA92Ovdx93bSYRi1YwhArrQgLdH8P1YHTmvk61sYAU
7PN2Dbov6u54r6bwblcSl6f5sVYvMVkP690jx2WQccGlfC7Vuk79IMPA8Y7BPUFN
mTQPuCneXvED2OWPChsZnwFfXw7vkLi8SffMk7wvhjSCoZMyV20wH44wws1R8YVn
VlN2lciCjhPIcQ0Exxc1Xf4BSCpsHglm3KgjzyqFjTqk/jpKpobB9iVTg5TFkkhr
Cmqgb9SrEsuug/eWiS0a0vbdPre0DBwOHVFPUnY1kngv9oLIShVxH5CocGQDJE17
DynrU1T8HTw4XctS2p1jz/mB5kUoieoPDr52u+zAXQ9wT9LkwKZT0ve/r3jmc7up
RxsF909+qCyFZ8kvuOcctdfgLyN+bCoJOjbot9HTMrTzNvm0Hau9dwFTLd+XWguN
KBpj7DvN98TsP0yogFYgDLk7/Zgvglinj1Cdty+B01MzuQ60WkvGs2NO8q237xOo
iX4fsXSw4aC7LaJXY74X6j7MQZqECQHEIr6orf2etG4fdD9t0swWe3yMbW1a+keI
acaChuVZriL2ZgF9unPAhpJZRaFG9VEAqXkYC2Z/DNH8sYjvL2PNo/YZCOawMUkP
a1v3y68/pqRPaSxCnFPBh+5nZIHLqblEAOwnJdvMNwzysX6kYDA7Lwe5FslEVy2J
u0q72UBn9eFl1XjZz858ftiLw4quhBdVIvGuKnaZL/EBG+uDdIOcxz5cFGMPdbMU
5fvyRue4S89Knczf1cmNhGjU/VR+oHEuYghYp55UxP/gpgMNWV7SFP/5qvPiPzGN
jVAzYHCOVBrvVfjhEotcT6PDOxzSnTZlGsccESK/EKVauLYPWvsZjrBlRYfKs7a+
FLi0N20JJJ1jt7dtLSswOye3UOR0I8FuH9C6bURd5UOfwsq16IzVXaxtQjvtOr6Z
22v3jAvUIEzb8ssuHDyMjozFPvds46iDrek/BXtOJRiuUj6gT6pJ468Q/HUYLVYW
vfF9MKNrpwCmOoVPvrWdkC96T49S9SXM019TgUZyEtUpyzZlxq7UZ1lrv3OulfzH
q23nmJT7nqGPTbQASoQP3QoYYYp+UJbuwSe/7BSgVkz0LkJU7+ZRuoYOy0aDsQia
Woo5jQ77c50fUR2OAqxJAEO1RUA8Yy9GUkbYMqY/rGcT2gHTj9AiBIz11/38eO98
aUB5qoETK8V3su1IWXgxowX4aSCaAf+dXHeAxTG7SRLFsJwRhGALRu60hr2y86ge
Mp/hzaW5JyDPwZ3kVStE4QJjM6A28YZew1dmB0RfH591dQUjMIC/e/ujR/Ulyn5P
AUb7J1DMH0L8cG1NMvYz7CBQly4rWvVYlVs1tpEzTJTfwrj2nnHHLi5fLczgykSu
e2L1NmYwKsHK1zm9OeKbfqRFrzngvtgM1M1W8grPcm6MVPvPNhBD/kruAfBVDNsM
rg5r2tl8S0qlUtfdBrgvUROWx7kqul2OvkW322FWRVatRrOTg49SLcBVHpFh6rqp
hBxV374DZaoUNUGP5+9/CP1iqXUs9a9y/p3gJUY8/26QYKQOnWfIFxIW6RrhbwOf
66882b9l5LiFS8n4lMHmK82Xb2qh71NAiUKwFf7+mZzKZA/SN3WdLUleOoG3xH2n
fv28zBAFOMRQNRvCJVHN7ROGQdwpnhh/2SseAOoloMWt+4yPMUcGjylq9iLSkzZi
uLW9zaD/Ch5tJe+59p0XWWDiTX2v0VebSQdf7SSBcugSSVOdHLAEk5ejkVq/Llcp
kj1fw04Jt/g6/oBxTGHSstZsDXzG4junxpSPDylsYfMgUyk+/d8dgSk2jmn18zY6
urKiRriDJmdEXjier8unmrpr7lDMw3SvOJSiQqDyHYnPy0Eu2fyTrvHJwJEB7+2L
yRPA/vNVc103AK0hDe0Oug+RmC22Oogct4rLlcygv4Uf7ZQm/URJlL6IUBMu4yyv
3Vu2l2OoFniBE86YmZioakj0Xge9RoJyA5TuCZE6hhYleubO7NsJB7bVBtHyf4WO
vBPolCq9C19QjrzDrMFu0E77Ne8o866KuKAy9NBhFHcTERs9MwToX1ykWqdaa3yn
iNc8fTVet9WDtHEto+UL5NzYx4UYCRoahviHzsMk5Flv5Gldsbe7RyXO8nlCJ4F/
7Lly5E7FeI2kNLaLMsZR5C4OnqlWDw3Xhfii9EXh858qB8SftEssp4psArG05Xrt
vXgRRuD5kS1b30fjc2QLAakXRmwfiHC4N9AOuWBKw8ZEnTPfaRltpONxgGwOkFcR
J9ByJaLkAl0y/ESDzEhzwcknKcOk3MiJApK0r+nq0i2LABKj1e2DsfVgAM6wWN36
hG7z451XTsC7m22OIx0XuMrEvyYASV2mlIex6octzwnCI8Ys5mIWHE/Wu4eOirJw
BpTAXyqAI/qEDsbtArGTl0viyD50+44HIbpQx0LxCxXDOwBvpn6+QNBK8rp7F26s
QAfDvXfxPva98wDuTnv/EJ8U5SmpUcBD7VZi8lMdR7wxYy41u5b7x22TpjoMRMe2
9+70emmJOjVhHmjP/94rUnCMocfz2SdETxRHeI0exbSrplBvJfrXgMFNoc55bZdu
bfsYJyBBxhDMq2vjaYa6wyRdiibYE3B8hvjNuyjNqXsukOTiohwFo3TS58L3x+0F
MVefRoLWP/DY7dyCc2MJys0oXOH8vvdfkWn7rvi9gMbsLOMU7WsXyRZ9Qy4KW1lw
NTo0V3vHJnYfeI/otuK4vmVTGfPtaYIKvpXHQWaSg97liHkvBEo2hHhY0O5X8NJa
YUPnbS/vwj2ljzdIXHN7J47+l4gu83roMNvunsvTCeYwzoUjaa+Nlrlg4AbX2oAz
vErY8Z8Nh7Msr9wpVDiVq5s9wUge+jowBj6DrZON2T5E0RUPSRdSPBzSATGoDvt/
n19mNgymAToFSUk2X3zCA3hYwe8mit4MGRX0pc/945S8u7XMh2xRAHprRbAoGFud
Wdk43OA2KentVcfj+76nLsyp7gJMjykiwdcuL8gKr8Mn4ye9b0MMHCKhIwv9CLgf
sZjbrA38oyhRA8ke3ImrS1WdTC2Jb0icXTRiguhXzaENvUpEpRm3wXVRBMGHp0MI
615P9iyS2WdJ35MGjO3J/kLW1yFOzPNVC7OcPTeONcYxs35pOa7IWHmXKpBM7BUS
9aldyrE6QsufXBWh32nt2uRPqmoT5TXcBta7XbGVr5DWq34CqZo168c52YWzjwA/
eJQB0VGvY/2M+h/xpLX+Ls2QPRIm86mZqXg6rUgNqovLTpz+sY3AyQDNqr+wyWfJ
+FXUSg4GohNsi38pl240Huec7NXvlL+rhzzC+0vaqFpG5FdhRektmkoRbzNdJvLP
DYH0f15CktOlnUTxDoEl9Ia7DZXALgy5jN4GIMTY0v9dIVucx9XeimKF2IXocGMs
cLuVvOQFlSYc+mgPZNvkGNFsrhLxKEzbarzIxXmm2Sw5PN1pTP7l8bJM6n9Mpn1n
8fG0QapfsmJciQVIMSkLaoIo9O8vC4zuIWIPJCuE87S7wodu2f2Nq8fLpwEqtB4+
djfd2f/PSpCkmIpSW0h/MED5i9rt9d+WipdlN/wUwEMFWcMwt/x3qYh9Kb4CSkV1
6DUeD2zdh3fZrtzS+9DYlwENntWMxD6ZUdhlzlP8XVlgPNMkSvwiblAQjQYboRft
sCU+TwBFBw6LDJfSupXA5rpd0womLrYQfT/+PvIiy78mDb2D8ZqazC9qRV3pz15w
Ts2zvL263xlwtuV3iBBiT3JGD8ECh30Zv8GrvMdHyU4s6s6ixoLEcy6DtZZzspZC
3RobxRaXK91A60kaS9+lmiqOTGKJMimioM3h4w1GtGZ+fwa9nqOFMdGQmlsOl7ia
lJL5I+668AkQFUBLVFq8lIotNuViVYGC1thgSrdqMF+/OITkqlLu4bbUu/bPQ8rQ
LtYEKAdLiT5fxxIY16xPyQGMMum2JM2WAvmvMjjV7FpQNtP57xjawdLENsXDjyvr
J56o14xNLW56XtV0JkccXRYW5lKNxg3TIolkqnWFWVqWJK/KBC4F6vQp3WuQP7nC
HMLQ3dNcNyhwpVjEgaDfuJkQdAyuLGoGXsQ8ycdIgRglCHXsD7nypWdzp1k+/Vrh
mHBo77y+RCsuKHK2Q2cNYcRz4VC8aeJUI21DTL2ZYNlRIIQfVDORJPAytS0Edks/
mmyE0ABoGxrVWoFUIMB6YHF9SmP4YzAA6sYjzRCF4wlQu7p1mxfMwUv0iJvSou2z
8gEZsFP4oB7GN6Wg7xUYoGZC932CzftP2DwPWyPzNyhqpn/tri5Tr4YEFMfvJz1Q
64X+9igfW0a2K02AQs+eMFMMuxv5j5HHcXzLo7ax4fuBl9NkyDfKeAD+ZhLXF0ok
Lrhc5uT28A14O6PqQCYUakNF53gp+S04wGagfPKcN4MkmGQeEc2Jr0X8RgBbi+I8
prkc4OJ4fIHV25kitw2m23ISfxyRkJ/CM3R72/8HyxMcRTn1OyL1yKbai5hlPnwQ
3+RN+KGVEGDddfXyPVzm5WSED4vJ50YDQnnOyP0YgNerwMOKZ1V6XKhtcgcGc+MN
/wDFVJ8K2UpE+oWA/YPtkvwvR7c0FDPtoEblbYlqLfAkD+q5DXynJ/Ekt4WWami2
OZLp/gPRRaqWMFNDNRZik3ISgW6+m/heU8p6IH6ArWvmYVh4kgDd8QPYLYrFQBGD
sz+JbnTYJmf82HErjYQm+kZwqJrVw7aq67IkyDBNqBaEOqOpaIvfZqbjeZYv2rVD
xDHoQv4U2haQ9mh3Szx5HENDRT62isjQHBtDkk7dWzgSCo+/z2sTlVHxFoxCp+HD
OuSC+T2Qc0/5luYUo9WgAXTSG8l3kxGFbbNzLFOWIBBWm5I7AQD7Ou3JjA7KMNrQ
TXDr39Inq8I7Rs4UrOaxAEqNg1INTvz58JJ4+FeM46+J7a/qF7LuMmgEgDawUDjU
v7HuzzrYYfQ8V8HiM9ovlEBOawhQTnk2E/D76GEiNFIWwfgU0nwqrcjFRzhB20hB
OzcQubMarBS7DMfx3JkwokooUI7xVeYJqzKbhhXrBQSVuk2MD4Hhiu6H930ryjbc
DMdfKG2Ag47NeM2qOZy/IMGdMBspwmORU/hLdUMmHEvGyvbaQuNlEqCPRc+Ng8BH
cvc7VSGDYgp5AJro3D4i3nbTLqeXFRRcWrg9C4mwPeSvgsJ0oaFGn2SU+35cq+GF
umHZ2cv1b7HggAHfjSvZb/t7674t63fO1ymgv/tqeuc3uQuBV2D93Pd1DsGqvZ7k
/2YBdYtjyXy3jv8Re9Wo/OrKn54WQaF4fh65+I4Iq1Rfzj8RHl38e3FjhA6HVMiK
b4RFqfb9+IyWmRvQueyNkcHddB3uR5BxOlvn5qTSGIVbHsGc9nscTypauewtEghu
vYW5hb3CrvvMJ9tNyPacVcYoIQ8Z/DSNpiqUWLDRaK2PC1IsaHp15RaBHw0qvvNs
XWNYIbK2+D5Bgl+aQWiTrNkBt/MiUOARPWmpD80A/xgiFDjtsjU0PD0p9t4kSOyc
er/0MsM8QxtPJUj3p/g0EaYK7OkIiKBT2edO3BeqNu8wndW7Nbn1fJDWXvBQFaLg
C4MYyOuj7iT4a8XJ+Meyn+YlnbcpCmpplzJ4nzsTv5p+LJVIDf+co7/vhHvD7+Ts
cQVREh+QIKivl+It2aQb+SyiZvXwNdOt3YRHHUY9xT7vMIXaAqwlsa+9YK8IUdaS
7Vyd0ZIBrj9ScCNjOScpYiU+mFQx+4/3trbuHDAPi0sCDjxTt60pSLm89SSJaZWq
eQZjs2tseYWoLh98/aLbldA30FBmoe/wNC8xhFCD32aYgqnOeV8o5zztiOyE+fpn
kwrZKCaOprPqbHUsTPM1+Do5cY/7+PC0ZbiZ/U9y1ujpvO0nf3rkRkstHIm4n8ky
ZUJrI/ux8zP2kgxBwSb1ea9NOnNDDFQJOgYkjatV0S1iXVqY0hfNl1xww//lBJir
yj0MvelgMV1PB+NqrArqWog5pO5Do5AKZiB2W0s4j65pfsjEwDL6cgrGqQzbFMmb
nHcpzKpITjz8rqd/rrvEywnFzX2GO9jgtaPPhLR9E5fwg8InvVYl8xuUa8CpGLlR
70ZAiTgr+EDXRW2Qqqd5f0YGBoJvy/mDxHJtkaiGERuuPKQcsa0UGVQ1yoA/5lRI
IBgITzPA/tOfLUloYDPOhvL9RbXvb4/ns3TmBYIrfJg0weXye+HDIc5MERTEJ0/x
+0QLU4PdJFc8QeKjH4MusK51Nbl02Vq9YJsgTJN6tTvvRF4xLyl4KVXIiPEYvSA9
xWItpNX/Sk1f3NOI6IP4HuK98jJmS2kqOKe0X0I+q/49zjmHL1ecMjEqT9FZWXPE
OCjEYtA+x1p8xJxpdo4wQ5puvIrfJfuvlwCUpo5E2QIEBujVDxAFmR5nCxabLNPL
J1QGjrTkgd6WgzdQjvVuI37V8xoZaCIEjkeO/Blw3O8DGeUTXyVRzqWb0cy+m1V/
TeF2xmt+xXRPmbovIl1UUhqMwmW08ABcbbBtbb4m15pjTUBuVJCpN/LyrabOxqPA
K7QyjUaFUm9NUJGzDE7Pt6AsRObq7fcU+o0PZbxiEAcjMA9q2dhXxiNdN729jAa9
740ftY36JxcJUACMv2y7i9EK9UAOE7inM1dS5xqjD0YbvWQckvxwcuLR/ojWeLFP
0Hr5VgyCse60ibY4iT1GG4/83jYatrcZLr25o5WI2sOVHqg4h0LxwqKhifU3W4/W
9XAEs+yVU9u01HpXrgLDsrHKOzLw6AxIKRbpx48itzTraNe/mnr2KhTgvDHe/JVN
3ThqAMwvwjVIVxAcxsljdo3aiNm0C0Q5T8aF8o1Lf4VDvj1s9HNCJ2QRJsb9CWy5
t9JD6uYdtLDT3UVeKwT5iJDde68CgxJKb6egn2Frg8n32OcaltgSic5jvFmEGve+
8mZU4Z4lf6oFlEaZiJlt/hUIXaRabB30hwoMLPyoqCktVJuqh3wQH7i3rDj+99dB
Il3cip/1zgGlF5DYtfiyyx91C0iNvESDriV1FcCzpSWkK7JShxfLFRFq4xEXBDDY
zyv0y8991/Bb+6s21B4jRfPfhHEnyLa8BT/8he+JpuLA33G6EPE7EZ9lNNUyDOaJ
0iDOW+Snhm+yrlgAQQdoL4iDZ+qG9Z9/9lclFqbrA6hZ4PK2ABzRO7czod4o1XzZ
jDCzU4RZYQ6cBwN8XTEY1Ai8cKAEVH0FHq1iUyQLxGodkl8h4B2ACLHh3a81i+FB
iSO25gcK39eNrl2HRo8GkLGz/VUqWKos5z06CzdLEsIG4SAETjCuFBXRZSV9d4hc
tdMnmUFX+e/07qnr7UoySGM5tDwjClYKDEMdegmV3sLVH8s5q1lpQORP/ixgh4X9
yYhhw5PNlmZMv9HtumeklWk/U4nmdjVajETHaR5MOdqxZLfiUVFGVWJ+J5qy7PY1
oIxo2quTaWrlGWUgOzEknpAwOArUSFlgGHf9U2QOmG2HPcSaSchNXjY22Vb0yACl
WyvyFbF0f7DegnM9p2/uGS8bVVvEcsIEFRkMTMa/RwjBKfCCp0Irout0nXDUqC1E
s9c6CN6U6mE11jKouk9Ff1LWKvy3d31umaTIhRC2u2Bq9Tf7BFCZIlaSn2wQCDRn
CaN72U3SL104+7k4TMZAmNNxfdIZ0YSDB4SCP2tfXsKg3pgiL8PUS0jZ+idyZ64L
bqGaDIGAchR65RgjH7cQu3kXBeZKkwy9iAtdWmaAtCiWaMb2K7flK10a6xCfUeBj
ETY20xryImMZdJczWBokJtf9ZHTOlYOpuGDtaTRrz2n+fhAjKeZedr2O3d3w3oOB
0YIZ2LgYIIUiNp08qaWBu0PeolgfWTPq73AzlAV8XPtA/cqkfHZGDFaj0y+0sRoR
BDJrmo1Tcaweni1aJCPIDBfW4W0oH55mx7X4HcDv5ZzkzUIclbK+m2VwPI8EuyV7
xFINNKuvc7NZqgbFJZ5N6CqKcDVCVZ+axgPhZVKoG3NdbRlf6sQb+3ZH3VtqRM/G
TrBun8GpWfDikWqjJzm7LDXqJed2tAL5cA3LtZDsCwvRgwKDDrs4MxBEAyoOIF5a
THhAx+Tk01JyASElPKFcxjwpOLvj01igj3m/jG4jPTBns87Fmk4AcV2roD8t12t0
04dd5PLKDJ4u2nEfL86HbTP/ZpueslHvM6wrFJ8b9t6AN+NueeGryfvknsa/vgNP
7UXvIBhR/W2PsFCOthBAGADvnCfz9OTthsEUJNrnTZisXFQDalQef95EqCEOTcJ3
+ojsdlmdMmAYtYyrLTtPt7gBueF8K8lRu+IfgboQ1/+HYdsb3k8IyliwKpZeYWP/
hODwpT0pkzPMl5USASioI9w3fWuKx8vFOBYhyjWHDftggaUemCzgPGfDSTSG3VBP
lO28PxGTYCYSw5zxQNo+S7IqFXE0F/MjAexpSIbBh+Oj9Roaa+o2whJqFP4UYNVU
/XOT2nMQUE+DTyN+l6soeSOKWo4s/0gSvIQPA0gJ3rYjIe7m+iSI5+6N89pKVIgS
fGDnkZVhd1XCphFooGUKJxguqIaoCYmBofvQFPhjNvT3xUjqxcQ/SKwmwhpv5Nvj
MfeqxeCeipGeiyQIm4tR55NOeQRsElSLC2XM7PFJxWM6v+tzb65Jy6vaTdQz83lt
wly9VXGm5zTxKr6Gy9U1Qqf2zBV3AOpkTb7UjY9gaVTKLcSwzOKzSztkUVAlLVty
mCIfGhBDTYgMW4Ej2YrJZ86dywhHVcyEnhBspyExooONapH8Zi1J4pL9Dy7iKtj/
b6VaiSHR5rV0BTqUDc/zfGgxJTljmxqzAaYic5R22FV7dOuOuvXnQRKD7JJF8KJO
kz0reZOkaDXSRNxE5QyrBtj0AK1Zp8qVtwrgiilKOEjlFt/jg+Wgas87Ks5U8pzP
NOmWhUXXTNohamPNg/SBRm4HNpyTYihOxbwC5I9uUNec6g0rZeayns0HNOV1Xq3z
QJjxyhUdoMx48OqOf1BE7RQuasgBZlzoOiEuSw5s6DNjaf3vaC/ZpBauo/tyN16p
uYsILBIApy87yp3q59mmIJQIYKtL2l42xmHM+SMd8csJlWkJ7CVygsg2sBqAnGUx
atY6N9DWJzfPxOy4mdvo8zxxy0C2RT5oJQsX6/BTn/O/dTjJL8RwFLfDVi9pcsRy
uyyx17Q1BmO/pHs+FLqqduD3PhRJgsJFgXC41CqD2KNQP8FXQKgWsq4FN/1tpYzg
Dv3DkfYj1tunKr3XmnRmUW4sxc5Yhrhwq7aOz952Q4QEHUc61yQcsfjhYvTeNdHE
qFnj0h6Z2WlGJ2YCT+fNZW+3Mh9tfJdfFOM+jZxRI8JlTE2JHr5msXgtJ+FlynBd
W3rTZ0LUnWBHBrDOhsGoB6XlW7dYtMguvYaxY4SHQ50sfOKAMuDY134FCnQ9lLFY
qw8vy50RicVZEcBHNBIn07zoDkcekSnsQdUFynEOTMXMIQ5Ra+FMEOPFiKS8CIRM
0DRh2NUzIP1ecyIu2e2zp6r0+f2W9go14BMsaMU8EP/EigoZn28pafLJHAVB3B+z
vuLkA6L+eHm4v3k8K/4llDE1YvGoGYstXU/+7GGawyREulLCOZRMJ340pSVdtFH6
A9J95N8c1MlTtsmyYXYeAXy2JrQtd93kdEbjVQeas+tsbfined3OBra2OBccaCkN
4q5xW+VGD2lM/ae9M9RtSxJcJ4fQwRE0NYrUo9jFidCtnarvlDAdfsloXEFK5Grj
TfIKYAiVb+KERzj5BjGilY0AlPpyZ/aEfLYHTTZ1/g9nyo/s97r99Rp9okAErWof
HxxuFmxh6DhAyGdkAN3Au6yPDHQD2MAeoKJQS/qPqKIaHf1wsq0xeFzp7V1OtTZk
jtZg3rY3JhP2yjxl47giYWGohrnhYYGb1xAAiy6eDhRa+8dtkLKqmC0rtbGbE1nI
cqpqHHNjqEUcy53+fBLVYTArepA0kQFt7aR8kkfC9RcMdrKOoKyEtOciYSDjWIDn
jMW4xQhNNR9oA7QAf7AakTwH1lkllVFCx+rhCB8YgwQ6Y+3oyOOmJZkfmNwaklla
DXQDJlHmSSvgcjQRey3wnP2mH1hs7EoSB116/vFiyLh5kdu9z97f0t6RA0GoJbOd
S6dpMSROUkcxaQqjVSl2U60mTaSRHOtMdbtwioq5ULgtMcFnYCW/KK+yqSFzPVPX
n8Iyap67JOpKa9si+TWN4HbL0fjY+wKThMvkNNbf42utq3FVzZk4OJOixTTJfdBa
uyilt5pdHJDmQwSvSqrpSzr7vMjeb8rrmpb9kisW3LmqXcXVTVXdyJPNJzONxbL0
D+VicmFdMsb+nsVwzGDLg1zThrGwijLNujnMLSBzqX3mcsgUU6fgktzMdngjTNBJ
8t7u+iRn3EshZv2tcsZRTqCX4oPV+bzmWNPTfkQ0IXJaIvsKSynFEwiXEeqd+7Ek
WDJHzq5Uf+ZMGF6RjUrOlfjE8glKLBIFO5Y6ZUCHiz+/k9T0GAkeGWO6aZ1JPSdy
4/qNJtkYxhzWJ8aT67jfsCCbzTyHoeRinmKBRu5GLNYYrGTInYKbYiQh+Cv+b/tK
MxW1DlMW2nAkhQFOTZuSeT8hPvs40JQT4nbW1WFgqCNpksAVA44ubOt1sRJWPhb0
WiBv9iJIr2g9ZAFTZ3bovHvckaBmABU4pPoqhUzKrujfw6F1MZ3812apWPaulvQ9
CIm5RCvkJjgfeQcbQUlUx/nekD0ecNfBkfAkAtW00BwZq/geQmheH9Du7a8jXPv2
59tZhRKp7S2j9/EKkSNommgUfcRXSjxE15qvDGnSXTBySmcjDxIOjAojWCWnG+eF
CA9l31zIGObRQ2REAgvFM7UydZMT9Jsmjutl8hdCLwhM3iQGbUqwzGF1m+GS2ycM
I6Fde/ryTAeG3WIrBP1erNye4Hi2JCwCOu+avyB8KRIBquo5pfp81ORkxjR8ikeS
JHUdBPXN2pXEqfGyi4h70lWsqF7rwEvMCSZG0TnSitaN37HsQh52eAxMEHqc4yRR
hjPGUJbyIlSs2iOyKE1Lf+WkyFPBE/0A0V71E11bnpfI0gdCV5JtQp4DEniRyAXJ
R+zJFezewx1Z1uCaLCKIUFfNsxYHMRRDPpAVktNm4ps/tsAmOTKFFolg8+VihSkV
WoYNibUyR5Hyg1gIk7AnuXmrv0U4mBinMSWA3eFd+vQqNSXwcBMD3dxY9da2i0R5
NhXGFRj6Xq7jm4r9Pr8/lY2i/ANmdRzvOMtweyhaePDMukAQyJrI5uuaGKdzRr7b
hKWyP1uFHpYgV0Z29uwQS2ZS0a4PXyNLX/fTThs0oAJ4ExRIFBvMT88PTaw5l1D8
n0P0jQbEhRIA0K8ZNWa5tL8rXKp3ruNfYZ36AzRazy4YtlAuYIPi9d4r952LTLBN
Pm20d5wDYX28AToOtEGwLaERo2eJmhUve5q6SDTNhY61MMiQLTW2vG+mWOzaVnAS
29pxHmwUIthVh25K8n9R5K7trNIzjoPUeUYtLhDMPlTUFlKeQ0sG4RL+pIp6VxAD
IImo4qu1RBnzniiYS+eiBE1OC2DWo8N/AuSKKz4d5RvWKpXGbwuv7zQArg66sVR9
w3J5no0bGOj8AMREf3mTJXNWj6CrUsci00eqlRVYy3qs+ENCKy1PBb6+qVyu4hqj
q3DlgzR2HE36VrgVfZHG80haa+liVplhZWo7nf9OXMSwPIc+t0kXoQ4A/ktyvJwI
QrB+kSEi0j3XISHQ6+erHTldBdfn26vrjO/qdVPu6GxwRCDSKyY9JptgEVrDxErt
XHOXAsscKMZnrp76TPrGj0aAO6qSEQi/ILSgPRAgvep3l7llWbi9KbohDx4aauL1
+/XwmaFeQvzgbVGMUEMmpvfb1AvJl0SU45FFC5rn4Vyg6E/1/ej8sU/8zsEp3Pdw
AieRBS7Ja62NYVVcObtphIOlOUgxzMbAWIbW3BQRbrbnbKhq0wBcoQV597AbTz8+
rbChYnanrYSSfRxps8FH9oXo6ez1EqJ4tp+xItm26gALnypS5rJ2bFYKrrWuqjF6
wP/4ept4W86jZm/dW7PLOz+7dP4RYe91eKBJ5JTPOudmRsI2uxND0QGs+KDRTDFa
7li365QDhFHMOUNBzvjjQ8P1YVUarqbtB5QFqb65iAQ1ZdE7KOGH2ksy/iAdwqvY
1PEDpxRQPyNYNzUHOHlk2GMlc8Ap0Ag+GpseWPtR1zK1AU8vuSptVe9GN/jRxgGW
Ifsj3cVHSlVrP6n+HCWk63I9TvvQcCNJ1SFv314bqAamMtzJoQhs0WCsNlVzwfu/
FSVy0tCp4+2ubsm27XWgcIzgBXCMmdcK+tjydTabvRCntDmCJ7z92JGLkVRb4ATf
1XinweAqM51fXWyT3dm6ktT/H4c1bCXsw2so2sLM8hjvYMKopvu9oKT5HyeahP0D
2OcKLhRu+mczpsCdZtMietuKtjfrlUGgJi8l+vFkMHNT15KYwtzmxu/mjoFBgkII
tGtRQGlulh5nBDv0nBKGLAlqlfAKIg7k/fcXGqBNyR0dSbIFh/5fOpAccAFWwWaN
rLQ6bNwkQiCRrEFUBrocTIdLyuzRoY5q+ADGeYIJjAyRZUWJKj7LDDvGCfpZaAe5
KoOF7cGhiaKbHH7V3IUCB2l0k2xpBG9dPhVE5jn8VRIWUi18/iqUPJ89NepxgkhD
d3KS0hNb376/VxxSlUkcVaF+qPnL26hPvvdVOLVH8IhxpGtGE1D5RyUvDdqekbn0
C6uqC0L883MTx1WkrFxeOWYY2RFILkt5Gm1RG27qOI4TISY5uBqgoQbyF0NFRG03
WmxkGjNlW1IWbEXS2bebtC/mpm6Xcs2Kn7Ep8UAmDxRQXnXd2Dk5K97waqdctaME
4v/d3k0gVYLbgTANk9bCZV0ygELZwU2Fo8h0ru0SZQJYmrbIlHA4m8cHme0GxPdl
tzXVShllVSxhk3TB9mKE2PDcPqmodTPexMnWAZeKfUqXs5ASs3FgrTBAwAOUEH58
gWTq1rDx2XfjtgTxiUTIVLIe0O5BqiJScg+Z7CkZLBan99FgUO3Zy9LikH6/8zse
dj1HXg8FqBmDAA/W806DJJcT/OofiNP0H9U2Ov872y8No2vNZcOkcQPcvYoFYkU6
3Y8GYGSlWlr2A0o1XAAHB9JQHv0+zcuD6O8/rhbcp+nmn9WcGfp79qDlb/vw41rF
Mg7+KDHBgHEMZQX6FDQLi4kzaWkztRfue1ix2ewRq4NM+DLzWpL5jnU+o1kJo/Lm
P/+5+oOBnionxpKokK+q5veRnRii2vAYCGgwuhEZ2RSKQuxU/U3gv1/xedXhyiyn
dDwYcDMHrWhiCZvhQ9X8X3K+dtKngLsUOu1kcgNoXd8KtHnGIWxg0rjTRJYJI+s5
GKZXADwle85R9To9jnVfU1zzFOEEh6xBFfzHq0FWq1GIRpgpL4+pQBvivnBSNIZX
Ic3TDMODNe1UQxJ9wHXeLoui6+FBIfJ6ifaBryd8uR+4d04Vi3gaXIL7hc5iEqtr
CDUlcAJK6/xOGJzUfn3cKMkfKTWsCrtg602gLVivbVezzI/KyC4sATurkrwRPkkF
Z7X2XK3pMG5rtbqRGAvJD0qUoncgz6U63oYpqynOSiKP7rWtPYDu+jgCXjHCHgAR
ukRRxdm8wdC/VsJVj0Y03Qlxx2ut06OD3mQITd0UpcqNtnDLliewZkaqO3X2DJuq
IjLBNRsvkgirxLPOztalOloDbcIeJmR56bmgqzVQIOYf6Q1A2u4mhlCfkSGMUxAz
hEervtJLP9U6EmAG1sVEJHGOSUtMr6S6ohGa9L3cQ6JzdEf4ZuA9WBRoJ3NjFy/Q
n/EeSGQtSYdE6GNB98i3zitS/qCBQLJEgPCqv2OmPluGjaz3ZuW4ku5hrpysJ49X
FDoZWizbSrnLjZzwIasygKXudOfFXegsiFoj/c0NUbzFKZcL4KoRDtBkiBu714xC
M3RzpjAPPAzWTT/thz7w3zQCxWCxzIFpgcuYyA/Nkfqv1HWrotZ4fnDnnsHZ8+As
+osn8bRuTlg6xDXJY0lu1dGe71CnDeiO53Iqk9paCFvATjKtEm7YnaOBuajy39y/
SASkl9+nRHsUH4nee7JW1KXR2vZCPF6FWjp9noB93SSfdYkSbxS3GMaCsHeKCG6x
NDulFN84z2aZCsxS179jdE0WV4HkhxeyIJwGFBbA1b8m9XaMJ/odEPPSeYGlbD2U
Mj5PH/aMtFZM+BM/6iUBsymW0WT+k/grW9IawGKKuqOMillzGCu0a3Ub0RxnG/L7
/N0tLsA3d3I69OLV/0UPjUFUH2TfYa0NNZgh79/fiDEH6cptntBXI46mIACV6AaF
AUZP99GcDJoKi9CzfYWsAKqNV6SCnqhLSRV/Gvo+1NElxpfOa3CzhXQZZcR3gBiH
CTZuDPfvn06+vszk197FWMEYMf90aseuHgGmVYU/ajQsIKyov0zVTrnSRDus/+qx
GUbiyFPT0u/C44AzflNBdbviQN4myDcxUr0lmOrJnHV1khzzTD5vLrLdSsBqWibh
ctLbiB2ogvkQox1StfweTZZLNSEvtZLzLQTzd/A926/NfiqqL49ZwwmF0E/K9Nhg
TbrFZNJZo8ZlPAippAJfYMaBEZndBHtJ/RyU5J1/e58Y96z/sYrleLB642qr5I1M
nDU5+R2LajG9cnpOfmirFkS49Za2BC7TVxTnpsBaHoDwdpt9GXoLLR+6T6pQH3ic
CbY/s+wMQM5pitXIzhzdzNEVq1+TZcL7T55d5W54GkJqAwMkVH5Le/7z/zvfCKjr
v0GeJrQBd2lWSc5RKuw1qJX1CM021yzYxA8SdKrzHgDysAU2EnvgnorWaeOQ3N/U
LggfIKbz7wWlHhipiRbFmoHpW74+MlAKa8ZFUM6wfaZP/G8AoKb4M6eBELHQmmxe
kD/P5zXpSvclj0qTSBcI/KViS08DzwLqBRflH/NkrKD1dTePSPJ2tjrCPH3jYl5Q
6aLl47PTV+WDlXIVr8GHBdcOE344x7nFOxsyR7BF3TRR0ZD9FkKH7JHlWhDfwtKG
4ZPR71CvcnjQxUfUk+Jt//OFu4Q2Yn+I+gMuiAgZpvqjuWPHFN4fZOXYx+ubiBGC
FzrBEF9TZMtK929XZMwsFfwbn2XZqRuFgyac6W+yVjh8CbLflKNKABuT0yRentvo
j8FrNJs8NT6GvvlUAOJ39BvrgRsGF//NbZkODXJ53SoXS0/jIll51YLlcRjX34Me
eLO3nzD3YgcTc+mD3zPsK14bTg+X2dwLcvC4/VvFaMSuPuYk/FrKPTTU9KiCFezf
+va4AdJeUvBPQdf8EOKo9yjOLBoBXNnk8GUx67r+zvaJlAmXBkYbfaTcAFpwM7ZH
F3tjg7M8xuD23XOFpujWJ/6Ba1SxWw5cBoGOYGFYsnhEd3RtICa5+eOBKKWGeA5T
4oI8g7gJwLa3XrlGjKQevEwtz/pbuOvglLP8uLEabdCboiUOFZOM/nK1Lp2B/LsP
DOnkXHS7R5b3EgBCVvCc2k+jMZtP4w5gRyXeJ5ATcvaLIPai1EoE5JT2KE7Fmbkk
sv3lEQ7eKR6Y+hV/ThjR0Jtp5TEn0FRQO/YD4ejPnEAN8mbjHn7mZ8gm8E+vWzQX
Phgx7uyYY/llz88Znh43uC5EUpkFj4Xsyaiq3OXQHnfvUXIhkyPvUPpKTJgtkOPe
CbICWhMz/gtet5Ksy56a1Ao+L+SHFnTXK8GHcrEUSetjy5pOYGsz6AEUBPm4mRiN
AO3vkTCxOZG170olt+bF7C/Ir+rnGIvZO7A4o9p0ws0sk/2Z3cYdv4ZLGfUtkNHp
reJU8CcXYVqOy2/c+VAyBJZGab2Jk0MQEFedXb8EIEo0vAhS1Xvqz7xjdGcZEz/B
/1QpfkurVtuvXGCODjRZyA2vYur+IN97PY2fvkF7f5p3tH33BiuG2+ie7gRCwnqI
xLk3Im7NhldY5bfuyD10NmD4DQrXzqtQ4YcFuTNO8/0F4hyDwuff+5+LLHBHYSYb
Er6iWm2BIWb6dSafTuWhAE/DJiglDNfQFsSkzXLP1ZCzsvLBppfg9e3I43FVZqLK
t2eqVbvfZLTHX4FbIYa4kilnuU8ULE738A4TkV3LsqrWMirwBDkM4Esm9lfJavzk
dSLtstQhyq8CuK5METLQtxfRNrzaCi7rCbTDi6dyhiFsq9D+bFMwGlE8eM+8k3Af
gT7DkUx+KRaOczuMhNuTWmpcjBTVdP7JQnVLL2g9H13bjT8na1LxW/E2Wc7m2ODY
zOStHdhkwcv+auOagKb9mpKd9mYtG5aZthoAUjtFdxl5oLfJbIJOlr4Vm62Z/0L8
I0wGVXAxRSIx2QP54JwxREF2XUSb5dytRRmswxn4N26xkWHv43BZU52eUYLmTvpy
qXgo2Qllq65dSt1s0YjNOHsq/zJ7r5nReDAcyukwVQOLl3jBpQAI5asvGMIzo68x
t2rTTxSleSnCzncpvVku4e05b6KhydTm7eWTgAx631WK6L/awVU50+OOQlHn08Cm
LXuueAkrd5VE8KczP2E26SysN8yuws7fp0YgaTMx7zgmpqyzx+vrLkKD1WK0mbtM
LtU9E/Rqj+SUlORN90aPiLW206vaLdEnToCfIq+oz/iKCo1j6GJMka/i+yWTCEsU
rVrqo0GtTTvzgSRZshGtT/p5KEtjzw/j9IRdJ6MtVx7O/C7A1kpWYzzypGYuUwH8
w6bmUL3Q3s8RNmMRCCVG5ZTJLVsbpTZcsVDjyEnXDzVEt5zbI0CdEuQMdTGLDi3V
+VK726mdglaDLbT78oeWacvyPRrEKhMwmtH20sPg+/lTFb8zApWe7W4eaIexoiEl
db0IjLIrfq25IEqHkeM6aG/l0hJnMVS/6v2Qf0JUICalLZbgD9fUbB3f9mAzKvJZ
8l7HTMoqGHvhfVHSFcifR2NaE+aygRDT0zd6Cknv2wQka8JWFqXTlv0J8lMwZMlZ
yjn7lM7SCgiLKF91zgjPuFoWSplnAtwtVhda1yhJv+kOaHx3i8aqWIl+e3wGA//G
/rJQegQk9wBZd3RAZWUZGN5xnjRcGTM/NjwSOPutjrt75qkkFPnqG04SOEPGSxYW
qZ83lkKdcxR+kdCXPAxOXIT+lNbgzFwv2dGz+nmSFwkL6lbhjnbNK5/cam0tGO4h
rBh/JHcvrhlP2K/RX7KXlbc6pdDNyEbwUSpfuoLY1/y14ABL1hkk1xdaf+ucCG8J
7ZehDngtokfwKV8CxGqP+VHvXIWU063evybt4UM8ABenG9P9ELrVQN5NLompX9xR
dyuURrXBTstvwfsTyz1jrvBYmVqgPntCBhqoIH/LtrSntnFyystgSxHT/9vK3XtQ
/wEwI2zVag2NPMPfoFcjDTluigZmDLI4vM01K2PUux39HuN1SZMsusb16Q2jX0fP
+YLBGIWEMiovIqktTqfr2NoKfBuvZ/q/wJMPJTyOouR7hAykdY3HjXY35n3QbwQ3
C3JBGhXfRKw1oAKo6hHVJt8mB2VzTa2kPFwDtripmtdhPnFmRK+WZmM3yczp6NFx
McimM0Rn4uV/l7Yq7CDfR5VWk5XqFaNlxCsZOIUKWTOsw5Xm+OvVxe1Sru5MDCwO
m0QmAOMtBKIQObohZnW+nyTRM5L8RHfM33v18UTErcEUG+j8uKmlIKGbwpX7OuEG
8XMae9gb/sjqumQLyePh3Rz+wyvjNXZnXgnt5O/RZR6E2J19WuDssCZJFqmG+Wmg
m2qLjaPOt71RG9khye7MdG8ccJZ65RJ+f+MpG/Z22jjuHMF9vii7dSgYpJTKMHhK
uZJwhFtOrFazcP4xYCUqseRwI408TaGFg4BVN4ZrvzvGKTKPvcQcSXXujcCXpdCa
nTvMPrMCbz+Ia333/9pfBT3XP30/3yizeQtQ0BWT7dtULzMzI3G9Kovu0K3vRubV
bmM6DyfASouC2tLQOemCP/VDjCEo7tI0Blps0+AI4Ck4lYdCFHxVRA8eR/LpPB+p
rbIE5Y31bA4z/CCqNpS8x1etF3LSCaNxjBT6CQl1Q0B635JZeqmJwImF71si3I9S
Fu1GkHPttYiAwjP9w/9d/1kF0uXNLr4NaXcoVjJbDhtD9q1cm9APlG67gxGRDMjE
neBH60OJvWbzu5ZkbbA5M5CdwB6nrMBNZb6Teihr3C7wMfgpKvhR8uMY++9E1doD
4VfC6wzM0kq6MJ843SMppwEqCQJN5PmwSEnU2hJ13X+s8gobVLywli4XMN1rXByj
mo7o4FWMfp3j6xptLoZMsbMHSivkwysN+HhRDGtXUe/oZ2u2g5jsQeaUH6aSGrHJ
iRAzcIbGjKG+yTXkdDVt4E7hTlj/0zQrB1UJw70q4MZApBnaRrRNNkmVr6EbRRjf
9zKjr2NDSLKYdcMaTSvlOXBXHRSR0GwHuzxJHdubm+QIzq3Yae3ejLEr/cf9Qc5z
bEK3r/QnF/Q1mNQiiCMjdzYbw4nTqUEjuEv/OI6x0Vfbu7DRu0aYYON5bZURYawR
cUj8waG1hCFCFH1HYce2VxSoc/0r8fCgjXqgjv24tdf5wg7ZLPiIa9oS5yr6nK5c
/af1UuXtESuYT6x9hHuGtn/Aw01uMMmBVoeqYhaol5UiaiKAOayGwSDMitg8V+ef
m4wEG5/aUIJ7JyraVO6zxYCHhAjNYkK7GI/hFBbe9B0mPAtGv7Blx38RCAVvG2j/
HtSMaIICosTH6ESXGjZOIssWW9g69ZSlnBA8NcBwFN1Lb9WYq3cUOlaeRgfvoJb0
/adAL9ipk1OuWki5fk4JJTHqAkSSSpeWB8sTIVMhyHoQJveEyX2swihcDiZLqQm4
jaQlEKvt83JUpGbtuRxZG98vXUeaDO9zc75biaJbqaHYRuLkfq0Is4d3PpmrdKPm
Mqd3hHhWTm8qAWD3th/ZyOPNa42oLni3kM6+x5Q47Ahd+WSBBmocWCtwq0JOQUSW
QXG0dcJup8uidT7sMzozrV9X50OsYa9kTFIOTvBRvXOyWOgHLFGOxrx6zZQNSvdn
epWnvYsdDgxti0EnhaQ41JJZKtsq460+s6+aqQv8PYuyVmDcx2sW+EZLj/Hd9lw0
o7NYbkGhQWXqPkf+aE4qZhHS0oAqRlPbvFh74y6Un70Pij7J2zE4o5uhHABqYrXR
dSiZ8uze0LNJmMQ7TJfaTByW3pFzdNspr9hBw0pYvMG6dDjC+Ws+U5NW0A12Q3nr
21WojNh5uND9r8WGJ2Z3Utc2bR+Vu9syvkisSG4IJnjvO+zFjlghDQN5TqKlsecK
WtGAhAW8ECwdBjKF+DLme/cwVFFLgL7gZjCGfb9Kj7z/KWSylIQ/2+vjngTLGeC0
9cjys8+Tr8sSsnbToKjarV7McjNTlLxrQ/3PXEek7FSpxqMnszFAAV5WzXTL3WGN
PZjNz6PzVmlCIa6Obh+V4N1JfEqAQ4DxbnjvIZwJg1ImWD0HS8lv7TcK7z3Q8VTC
XOhK+jpJkGngQF7wZo4wd3foJMhoYbHCS+ifHgm7N6tCsQsYnGCjKgN/JfJTyzyE
RQ+kJeXtY8UINT1Uo70vyCpN+pDklWngDmAaTbGzgIbgcRibDQibrRfIKqenFWav
VndB/WlScenys2Pi+apwwGaIu97YEpkYXFxIMrWwu6P/VZU0uAvRHcDh2NkyC8Bi
m4Ign4DpvvE9nrdjpZTfvLtAfOU7ZyIiCA4nblycJ5yAobrwdeO8WJZAtJLFOQrC
Q/e3nrcWCGwJNk0pKL2paP57taEPm+XcZ2537C/63N8guCCHHlLheFvblkWu+pfC
k8Mg7wkg/DS0Ubh7pryFCQHYipYDT4PS6DWdDD30LDEFVRWObkM2UiqYQ4iAhnsd
cFCg1773Xq010lah2lkkvM5f7HhZsiCXC0Xtz4C0ogUi/LS/HRiBhMB2AKRH2+wX
IpQQy5475P3dFgMiYD4492bizL30LfF8zeXFlfpUIWR2npuRzwLs9bijUJNrUDbo
o36XnrYaujoQjFypWC8t3w3l9V6Q7gHBwQnVj06jJy4p0SnYD6xdMWq9E3oxIa/c
do7MFOQbIoHAPhwV1GqOQdJTblPsHATHxBtw9KHnpt/thnrlYJ+jP5hJBnOODiIi
yqcL7ihgTYSCWVnJO7rvSWbuf4EHecgxgMcNMtt0wCUZIoBYOTp9XQ6k1FPtg2fL
xtLqIli294QGb65nCtwJBDOfHL8qqtbLcD4aZ1aFAdFm1rdZQxe5WpFcuJpDEKcq
oUfOE1iP3L44lg7SklnGg6MNyPvJzgo0ujg1+p+VifcCIeneq1ORxMqHs7RDKI9Y
50Axa4+df/AIMcevQ7v1GQUdm7RP9lYpDTuy32qLx1lBHi1w6IhtkPizsoXi534M
QujDVR34tTt8HsrL8sOkidC31M7fjwbQgLJLdltMsJSdwSfuAJtxsv7pyTavST7D
ome+yn/s7T9BYR0IthJtjZ7tBDP0JNxd5uQcOfa0/U9ZnapbChgQnaET0d4Og8yV
YpWIiASaTNi+DLl/NjLa/DJ98niKVMh8iJCDCVEb2KjK4QcCEhteP3WB888yvttI
9TP7GNDYReT3jSE3ox7cExe63eXxwvjkxJu5uwvrEqVBvXTP9aTU6LGAF35dSIHJ
9ECJZf7Z9TBXBC7+qR7PukvxuNKkCdlmWck8D8pCwQCMCXGC1C/bBp9VjaxcSQMc
E+F41lUU9iVsJ1wGVhk3c8benNWqldNGUHJZU8NoxNhYOiEZH0cwA9H3z7hxqYho
c1KNAFcHV8ziRi5K/4jczwFkTQrYUn1h9XrB0BcxfihbcJGyB+BFiAqpqm1mnnPC
g+5X3rI7/Ei9LEMbdPIETYJVwqggjOIYEegjl25/gMkS8EtNay5Gt7PQ4LYF9JnS
UfUrsbOZS2xVs0xhAdG8hCRK/l4RiMqrOHj3bZ4dzZnu33lOfVBx9II6rahhtIy4
WziPtUN972LvTweYtqmJNB9IxZvb+8pfc+edgSASdG5++ndpHfuFscGTMpgVsHlP
yi7/z4utHkpCGi+fdGzfwEW0wETlEHkwF6g956kGS0gYMsQl0i1s8ROKExzrmUF3
gQgx85HyKIzp3U9IoJGxpFba7AUY0ZfYErsWugMiw4lggKUybX/XreIxwzNORgP5
LC9zio2b865fYAajx1e7F3u5UDkJC0fmxSyP9W3KZWtLIBE0jWDxXcLnFtdVLTLx
mer/hc5F80Ss7MC/oBtBtZkGJ4RM5UZN1b0HG/t4VRVbDgNBodxt0f6wDGeZUx20
FImaTe9UdO65kwslQ2VuCXsPTjjeElnGeTHdlLqwHngJ2sqhrfdy+E29P9p9LX8G
xZqA1Sj6O4fkT7STGGd0Y5j4e0ROwHRJQ/O3DaG/sYIICXlYCMR0cia1gVWF14sA
Uh7MciShWCZxltQNRb2KEo98+bnK5/2kPGto99XQKoCinY96+lbqx8V7mF/toyMI
vcnUq3KOCe7nUc0OwpbPA0PesnxOObXH/BBrr5Cx9zTcNiWdQAJnYjpIVweZsC8e
gPus6ay++hI1ucW2bKSbZHLyykbkfbeV37KwuzPO1wbwoJUU7mZyQnR8gWzF+bmO
dV9lCAoAJqmFLo/jW7EV4uhKbVoMlpZX0/pkJU3GfsaDG108Zgu1x0g1Uzk2K+gL
3aVHFcnF/U9ULGt8eix3siXWOAOEct4k14jseqDFFnIwzZdjzyTwEtcJM1QvFJQg
kdg+qGENfmpeBI3T8/6Ewn/Z8pI0Vl1wzGSvI5pdblWwbYyWNeJ7PHLvrjOcqONd
Rdx1uIJYwCTOT6VAd1ql5kddcFxyGhg6P7Wgy5LiAbaoNH/aDfikxoF2CkvCNvwO
viWPNFJmPx9tLm86UGgWY8CEGDGHPFATMGEOWfiOTeP1N2iL3pBVxbFuAJJ5r0rI
L9F0ssbq9YzbgL1eCZUDwvU0bfbbo8MqUhXRBpYYt5KsHOp3nZS5MqdryiLwYfJS
t5iiQoDEGjobb2+MDPBKeU+ZTJod3u1N/b0f2gPNdVCPSWvqPlEsCsf/CThcOfPP
Z/ne7LOw3unIlnNiw7ZmFpN0yI4zFQbubj4aazMOJRlu8qBoPOyDUXTL/VlpefPJ
uz1hx/kNGBnn0znvDAwC0mRW7jfdIOGoQKuPDdErTkQW6/+/uXkFi6rNsS7lnl0/
AWSdHkv1bqV/wF3vWbyxsbpU4dhQxcnNhCGBTq7cheYJJ2hsW6Sgr0l1ftn9HBrT
WcaIFvvxrk0bGz+OVZGpoXjqukU4fvXZd0Q2RCOr2Oizy1DGnHI7SvIx6wEOxeaA
6dKmdzcv+1TA48OAFJK0EOgG2FM1nxXvnpk1KZn9NlZ09KP/smxTUNVsSlGPm3P8
KDo9L9F1TRdV/wh5EJ0yJ4ABy+YO8VcWiWQGurZpSzoKowiGpuFaPBNUvXGcONvT
0Bb1SfHgR/t9mRlvB7CBO+PYaTlUVkLIlcRXiUKezM7VJx+iNDR7Cp8h88MV8CsC
ScVE3kI7lk4ojAXFSEKdhfNDex1e7xcyOiCL73IoXmx5+18q5R2NooY9hx6Sz0az
I+VXCEiJVDRD0F+b+T4XOh3p0RN/ktiV6sIZ4f9ePcKXlzdqiTIQLDY3hmfePLLE
atDIMtZwuX8xoTWLcj/EzLEOHLR1KaV2iMsrF/yk7V+U5j3/rH9XZohfpQe49D6H
4pUlDNrTaDU6Zzy8o/u2qthF8JKgFbthGS+pAsZOXT+klOJ7cnUxIqAIER90xc46
+LhPwyYwbGyYMJJqt0qgY+u8rsSEnJ5LF3fg8s/zKmF46Gq8I8mrCnp+ysxOSny4
NgaAZFcHakRJxgDgM6VLUtjFIe8h5aFAXaGcAtonXMRW6ElVVWxLaBuc9rfPclsg
sXYUcTQvBKC/OfkFccyYuAct4bAWtPiKBY3Jshhz8/NoRyltpByf0oYJrTanIfu1
5QAcZrjWlceUxh1rwGmWRCYLcFqv0b9128DpmxwRjE9UcoJnPstcwkLIXTv0xqMO
aGkVQHEMuMvtOuRQMgKP8qAkQePfoiJDvX3oLGpQTxwhOk+aClaTXJKpsmMMuS2G
lnSgKKak2J7Z8dbSUyit7HSajkpY6An5q89TltRTa0EADJd/EzmwYIVWCYTRvyO1
2VYcZQELQvFlxjYlWQ7uN3IK702T0R6wqAixF2iT5KR+W6vpKatXNYYzFfffxfgQ
BrLHRjyynIdlBh543N486o7Pybu+aUMq6tl+KEfxv0cCfIs1JTzIvntnt1yS3pQr
TK/4zR2KNMnz38SXmI66yVa7tUHinzssJ9is2hK519lQ1Y+fTZSRPfMm/MxKPgxo
+XGsPzLhxgTOmIDVUHXHrkqQLFFGECh2pqSWKWZQb5XwUvx73riKRAgCGuk3oYIB
jw3dSzwqzO7fUh1j+CWolSPwPdnCiC7crG6ftsO8xkQW6r3xDSGu77fXL9dLUDiK
dW5k4+vCf5xP9Z9ok7JLgojKwL/Nqm3PEoJMnu5F03Jbvl4FRtfpINDWcxJEqn5Z
P7qgBoEoLv+bagRYjWRzkdrtVH8I07IZni0R8NxVHipfDWWol7WO4gHwlJeIOvVY
HUmEKlKxkNnYrNLUWj68A6/qeaMIzYD/+KkqwvgkoQ+ozyccuh4mFvaI25TrOp58
GHcgDsH15ZYhUawAPAZozxDuArBnAcgWEWBv5gTB49u0I34v/eMoYwJ1yJzTZQS9
RqdI02y0XukNyMsUstW+4QF8b08lb+V8acifPh+JdJW6e1Slrs2u5+pp0HNDlKZV
d1koxxoD/vYrhC8g5BK3sGJfCye6FWlq8MI1IcSHPIa3UYFbT+felrpHwr5v25ax
3gLNACp5nF58S70RRlPQ33C8b0X4k8gaSyPrxfhukkgW7sh4Xxy2ExiLfbuFT6k+
/eKByIjbW8Fdc9QcDywUVWABO7zjbqzFuz0aDbQducjW8zimuGyD0UGouBLq+iMG
o+6QoEuPXMdNLdWhySlX19VAkls63H9aeUcYMSAb1DBwFiHH7FWLu/BlxtCWEWqY
w4DyfNev/KkIf61Euwsq9QVUYWODgCPu1Z7MSY9BL9buuAhx2wB5zWPIhtT8z/Ae
utpXM9ObSM0FuJgYWv8Xlqh/VosB6yl7szsQ6nDdR1gS6uGPtVhpgNfM+fL0vWgs
rK4T4NHLzdnVqGFiQLVmEXeXIEWTpuMecYSXMp3gaRpZsmLHLbUWL6pLsFbF0uYm
7MM8ClRSSlxjbNqhN28vLNR2yePvEtoRfgmknjV9XbTLa1na1LuI/95+bt10EPKN
T7u3zPSvCJJabZOeolx56nblY/YFnhSfN8LYD3AtpboRc/kDPdtZ0asTKsSzrJRZ
e7ZkRsB5jXS/F/A7H6EfmCA9nu1MQMjZVBR0o+8mSVGNmqn+Kl6hhmMEXI7gKf1u
DeRHIjNX6QCPK5KEisSX3IZuWW3kmDjlBg1crJ8GOP+02C3GQweOKSTxIwru/X6N
dX+C/BSIStovsyis7DoyVRGsqONgMT/zjFBUETB5BKhDMIt8VnqmDYGpU7D5YrSO
J4hA+4z7BmGd+qxNywxXlZd2ylBRjggbF7Ctbnl7BGq/r9p+QfXsR685VlL7ugwC
LsWOdJjiubO4rzPrzKL9L1e2wPMGW5ltLGzZ8btgwqkzCsbw0g8JTlBuP+BsO/8C
OhIBVyDPgldPLYxf+3JQuoHWiQoMBKi4Em87JFEbeMDGMNtrFnmo5G9B6E2WI1c9
itYn6agBWGVC908vYhRYKKCEtQRXt9BmfBqXZXY9aU1dOzGxRXtAzsDFsRLil+rf
sGeZr0f6iDrWskbfKSuN4uNKpO/Gff/TpswrQM9w+0VauRfWFWXpf5RCGlt69qj8
cADLRWJqt60YLwSg1k0oLXX3YNHSvSb19v/YvbfpdBZlg8FLsIj1XPYw6qS2SxW0
U1P9NglLtMhKN8J4e0THcT/3xVBRouo7dMJ8b/OaIewKPN1IOMAbTaBP+HXtNmPI
VYvpNoK7gNO2Q20sbIMa2TepruDO3MfrTvwRzJeTwPWlEth4OGNALEuRzoTx1KtC
9jAXyVLf8R6w2S4nY8HfpbIhsd/JRFh1EKbUFP/hdjJfkmsCWeQp2HheI+TR3QXz
YulWJ0Fz6sBEvyVN1LoqR9JjnQGm86L2O/UOpJ8qDxyzKvOxUorXaMXdzfvLeaMG
GDUySJCzi5RN0A4XxJQbjokWOZum2mBW9r6Bi7kZUDVytGUEADJfQ2pUfJT7f5lV
ANyBKd14UoWep01My+rGa/swunzkyTdOxEWNmyEYgGjjnJ4LZ09ioXvd1yHoAWq1
bcmvh5ApRGGdcOw/p2MHEp+egSQOrpB1HIjGqr4a5zqMfeo5hsP9sQ1hdb9sJw44
6BAq3pSqaug+3578EkE5h2AjtfpAYKXpO2KbMP4TQMRRJForOv9HLlPcLQ3BJH6U
UGdRFTBU+pW0Ezws+s6TRCMcjyr8/1vUYy2/IDCLOxuqY8NLoNB/VehbO+2uUMeX
EC51i3EC3MqclhDs6W2uviB2D0JvGX9RUg+s4/KzyWQjhxbOPt8dT90+7qDMuEfT
shOnVSOHTUN17HTgJH/R+M3f0qKOAtdBBqPq80do8vXYmcx83sNz1EatXbAQlYdz
/8PZcTtrp50jon2z06BcrFCNildR+2RDAQQ5MFdWMTIXgq9aavReO9+xdcGZb4Ym
zxZfvTZRswhpWLK9AgJdBNcKT3dlzfGz0aa4XYaR5CDbbJPxKWZLBsXxCFsvNLFh
A8Zi1RxDOdgBFbf7e+O8rJXSAa+agozYNXsVeYskJurcV6g8aRszxq4NLUhyKSHD
00rEer52N+EhsAITgGdfX44e2k0SmL3/240wW1HHMGZxFygBu79WGFoRdVPYZB/W
b3BxwtL0DOAHIKIDkX6AuyHzQ24AEfd/WMqP8ZLTl2x/tOBASr3cfLvYHZDaPoI/
oVUUq2H8yF3stJYSEcVF/K7XYjEg1ce+KOCuGFQByPMxcWT67b5HfI1+OejmRT5H
D1suZFMlETJm/mbJAw1Ncpi7XqtBkXUGJC0h0dfVt4yBGJ1C39x6InA5chf3bUV1
oo4xBgt1DF6hukUfL6hXHQ3fOBLq0jZmJuA5aVx5p77q8cMGosKk7nCupOmqUT2a
Jc/Xh4Ui2DVaNJuxI7AuyQVrx1mK/40MqZfEfLLtvVZZ/h1wwew92d47jIWapbwX
2/7+pr+VgUEgp3GxIwoLHG2xsxWQt/HOt2IMK6zdEbn1hifqml8WKNLQdZQaa+rZ
RLcyVjdgSWauNSAUX1ZsL6oojojhRJglp7TMIQbPoBASuhyLDqpOjW+WJjhYE+/Y
w7dtEMWuBMiZyjkrU8mmhrpf1hV20zeaCe+DucEw/2MbxE1F3ERmpkMYvHItbcZq
Ey/fjtjGQnmUMT/dvRE/qzULKA5ohkz9uHlFE6qiuPhwusIrPosz94deFGUgtNFt
DOAuLxvxm1fMEqgg2v5zX/TmMD5yiLX4w6YB5hBI2PUFgIhSEeMXT9okX38n4iQC
Pr6xx0MhFby8SNzi+aBaKcWZ76Ov1487vp04FTBrwVDIueMCsjjT/wkGeV8bPGai
jRViWifgEiBCL0OZXnJxTH7k12efSgbyaC0UGVcLU1MOiO1dfcakxC4zTeiz0rZ0
uWf1w2iQ5+53c4lZUqmdskrc/dhjzQXHrYTS4JjJ4P3NEIOiGj+TmGLqPb+OKE6C
+bk+gQzE9ggK2ALno+bWWUSDelKpOz+UjKzSHLndVMWTew1XM/1/wY33Vjex4oGS
f0ujKtoTvcQuUqHC0gvO+TspyCAEPxmL5XtKpnDurpAHfbyaiiLN37PQBs/RgaLx
KvbfUwjom9SeQPWwy2q1MthRQ60BBGkJaHihsWGzjt8+Ic5t8IS8BvkLAcW2vKTM
ZRJ+cuKVSPVFm8Di1C7Q6bdEpVmwyjO7aZ561HG98IErRxtJ2boDePzTjV+s4y1K
hGOflPc0uBWVw4gkWu1ckWoc5ZTqLNQmti1sd24mbEoZvhqqKXoQQOTSFTeMaaC0
US+1DcOJZhKGLkcr7xbxv7B9suDkqeh2et6R/tiy3Rjpn92ciC6q77VPJL3ZjVja
kLSQfLnjhu0hN21VYhtxVk8ehwYsVAK8/TctHmiEfEAKRabwfWaEJNjguawALvbH
Rv4s8xnn21vCp7iFMFa/DvYA8YUDDtvre5+IjUJPY7mAP7Ao9phzxUGjKCK3g4n7
Ztf0rNRlhPLg8u15Mch4UPdk79TZUDCzoHBKPh/1oJkIvezmmwZRyb3Xc0V1+r54
2thRDVU48tfkDhNrB4tKBW9kFaON3pDyaXsHcnFPv9Kat3jXMJzwd5O1UN8dmDa4
F6hSUkTY8aG5y28Y9APbgACXjNvCCtaWxhZOxBxtZoyoGlIhJbzAJVTwySDeiuq0
gAVobhqOPAlNK8vTJkSKw/fZqawyzJ4PJXcAi7TNAnqEWQZt2fz8OoEU2mCQBp3l
HY8DDYdkHBoZcEScmHUjW4LPHr/cHVt/BmT8OKCHRor2KEDKHhpY+o4cawVV66q0
16oR7BzaKXEqdcgBwlEyGhwhmcnFdokU4CURndoqoyQkKxw54/VBDRWTPmQYpJ/D
t5FuMhTZZ4jY8xlMXLpXxJi6nN2PJGKDA88eBfi8pBBF7cnRuEYbJqjkl1IZt1Qh
LpDrvT4aFPpNJfOE4C2cR47GcEbRrkswfoGTIglOC7gwbctgRjyYWv34JiGuigaJ
FLu8unDyWcHO3rJ7Txjc6f7iUa1LOd891JQ+NZEOKf2tentduTBMQmVhv6SqlsOn
53OppTvKS58tZI/mMElZoypHLMme2QtESThuq+QvdkrMRjm+WberZ1Pne+RfD1y0
AEtKvBr3CyUVXG5MAn/SdRnmcZ7maV01qdkjGgjMk+viWJbEGraLzJd5OEbGMd5r
c86tabpQyP9Y2ks40wOGQE4Jk114u/gJAmiikVYoOq4pkAOJLB9XXGNQVM1GTzeN
0Ciu9fD+WjX8Jz8dIRk27w5I0NOtgQcHmX0FpzJ9bIrBekGXm2dTPgnBe9fX1Nat
5ajlgIWWU+obt7fm4tH1PombgNBn9xeNV6VcDP6RPxM7XIbYP/CDbUaHoXeIeM24
lhzETF9r8pMEnAya4icEeck6OrFOKP62OBErzKn+qKa8t+Gnzvnx21X1Mb/QyQEP
NGQvSXmtGakUH7lDjjUSPsewnu53kxf7jFni+xaAUyRHEoo6Jtu57On/9fNwlsbr
ULZJRcdAJH2L2VLn2mlSaMMzFHP1hOQ76utjAhFtkX+LKQuFiWd22R+Vc03Nb4jz
zgv6KWZuy5XnlFykNUC947MUFf6LVHuFF9TBjBoKzDbevNYg05KzKC99c+cQFrLv
ymHRs93N7lH0d0KW3UF7iIlmPW5Dww5r8t786XftcUXqn+gW9nbuGINfTwIzkMSt
E0jO6P32KW/PDsIJDBJAjxAIakycSb8TIqjbesOaILZLJmi9eBKXsjeYAAzFpp8d
ikxOuqgX0ddEV1pY2gmPfkzyehyftrCg7oWE492h7Axjk+JcxBe/ZGHCoRJpGmBE
TXxM68/kW32O/pP9CBfYftGAZcsmJDlxqkInFXrb2xMUjUr2K/p3zbde/x41MlIZ
fdqS68weGYRkEjvTn6OjWrlm9OaUckKUorIkcHt5t3LnibbNbGtQ5XxXdMycsPIk
Td/KGcl+slnrRQsZNGtOTZRCtEuet+uzkeY6u24LvofbVs2Q0DAD+N6GcF+QoxJv
W68dzbcQFZlPVWrrsiUY75S1YEur09jiWVCCZmAQZCcv9GPfU8aS3N9Jph4AYoSY
VnM3brO8/rQojD73GNGF1lAWCYjrJwAA5+5B+eMUkbJx0zBz/T/cNNkM5kjo8Icp
5x3Z20Df9SDSE5uEvxEXHklrtIzBOVs81HrYwGOkcPwW57+1B8eMnlYGdtWMQ07m
L3fxwfufFgnz5gUwkOEqZ6a+KwcxIgjb8e9q6rFS5NXknr9i7virQXPJVkjmkX8/
C1r/Swy0yxrZbUIx5FJsT7K4eljT+E1POyKQJiX0VvJOqXzAzSFF9nkuAu2Y8SmV
R1hgpeAygDe4Hdd9AKX8smJvVyMBkCCNvZJSgE8KRqoUZ5CpkzrtVFNS0fUjRgZK
WvQoSk0ha9WL0CDMtiayxLiFiblIMEW9dTmL1+tGxnyRpGurjpS0uimntYfBzB4K
tX8RJ0t9e7dPmbal7SViy1KmVZ8cR4hlKj4cA3PqjqSNJDA6gN9L4sKhOsMnf2Pa
ofxkixlKDo41VvoqnFxLkIDQsDxqKkvKOFVikeyXGGE+2LIH8BCaRaZNyukIB47Z
xUr2WR7SHJ2n3vRzbE4Fdg4AuMi32fbMAMqjIHJ65ytdswrmgQe9i8lpojKpjNtv
P6ZOcHBKlKiN705lndmMk4juhlgDOKA5mvLbjHRHonTAh6GJIafh7HyTA8qFh7zH
VH829BvMGD5f5POqllYrxSsGMTmNtFQ12xRS6P5NJwHVz9g7L/2EcoA6B8kdZcRS
L+xgwgtFYX6MI9vjL/9Zs6H8NsZglaYo6HCv75/gfT2NkTo3DcC6jJ6qKL2YYvB3
zu7QPbg8HFMr3nGoO6c+bn316JPnO4Ot2kA3gMIaUPShIpC3wm23gSRiIQeUEDYd
//mAN7QbySExCEUzig8ZK1FWVVSPrXwKkGrW45olJnHigRBy66bjRWaNSU/VJuS4
Rv3e1sUg4K4TddbEMone05FhvwgxlOL7wkE7D2XocoY1j/uw5loZ3+foFUtTlfIl
9jRpPoVz0dpAwwGwgv9KlYJ97nhMdSWNHrwjo5hUNsDqQQOtJCXAmYwEQxCNrHUm
D1JkAaRb8PRUlKKrNKVim1XzSukZaSYXRihF0zZigxGhRru/8dbDjlneXvW4laGe
iZCbNVpgiRoXAXC327ViFpkAj6pF1OmVDmPSGgk1S6Kh3HAVh6BLilN596AAnXsa
WKkw6ri0GLq7n41pdB+N/wh/5Rivy2285P0TI/W+VF82s4orALPpFf0CFgrboI/c
gOfveeO+kSe9W/bNXJsF0QtxV6ZgvITLU8wQ1E7wpkWr/MlT9wEgpZxLfTghrbig
plxrOTA6XWyZ+mU7F/MQdAFR2R6nUgH7Fg1A21xs79b8/lX3yvH1T30EBATCVOyE
YhgJ9veCttXaTXuJ+/cpRcUBlY9/lm2a0u5LoiyOpuVXyrL6pHggk2eJxDgjkr75
Z3NdlOzbTQciiMZKLvkL5tkwYXZmpyPbKCLKcbZ/t4BuiMxXF9Rbz4YEffu111XG
j7Erx0MVneAEhsoOFr62E5zyweN7NGqjyBBFFzI47F9ECbaNjvlEX9Yn30XtHaAg
oTQneW5OxW2PKhA9W4mXLm9Hj41wnmNaB+lmmjL5vpOmo9Ar4lBmeisq0iFHtokx
Vzw3mjf9creaMU5ny954JsGLCtcKWPrkQ7ERtW4M3y3Ugbl1eZX21KW2WFujj8AL
qAjXKGRVvrr9M8qbJGHKdNHI9+njlfm9AazX0lbUCBY+sAtfEsBr3/a/BRrMKmSa
wHjxHw14H9rso1xegYn0rZ1UlpetJmg2xEIc4EqqlwPzhfp5KhNYMSglewU3Tozv
/g7CIvx0ybQTGqT4mLBD9rDlHNKsE8BKEzPXHKcDca20k/yE6pogQ9S6zQj6khCv
tBy+v+D3rZMldfBZYLdLR5bhQn1xAPsAknTJ+AycgQikZnWPnW7JoVQRquJyrGsh
uyPfN7m9Q12+5X/k5KYk5H5JLK54vURcWRnZOYk/5wYi6SwxRUIRhADdpDzBuBEh
07SN1hLE+2F6JrXZi5raHaWTSJV1EddHLfAZ8mT1aNeo2uymgq0HgRFymfrULTiw
kbvAe4T/x1sFTjuTztVIZMp2AXf9hrEVYJOxsBUuIN2K/ZtCHNmojm5+jE4+RBEt
nTv/gElfykyWjm3rrmYahcRVTLgi5tNIbIQfH/Hl6Wlw9QSISvWc9La5rKCMxrol
ydk6o0/FuGB5eq2FCYfuN+dqc91Mxa+9pvBLoYeI3apPqpjaCVt+Quw4K9YltyNW
phFqAZ7t/eLXvzLxg73BfZKquAd8Pna6GgjaZvlnO8MPKIGjVADSlhcfyVcv2QQQ
KMiXzC0W7PkwL6fahZZ+Aiw84nuJsygr9cKHBp2PXSheCuPfFiGf7HbvdgNk3lNR
bI0ZqumO3DAOU9COon4+Yo9b9q6hNdhUrZCgGj97Uj9WqqydAfnMgtKhWU0f1NUp
430MNTIpx1MwM/hYlJMdkw7FLgx+T0383i61OdXUuQRRYKKBPI6I9+7OsL1p4UTW
AK1quIQ3iu2jWsdi/R5GvL918WeOTInbLV46LYqDXAz/ry5foeJNis/6B2hFBAAm
rblKh457K9dV4pQAenZzMXyDOFk2tMTqehuflyrtVcp4C15pk7qM/MCpQ5iOT584
sbLHyB5qYif5Plvf1wnrXQUTDlsua+MKCRYhOHZXkk/wY50eDER/MhrqMao2HZ+z
Ci+4RRasaCurfC+lnQ3BXI5lurZL2zl9HhCibwDiEvDnTVCuk7pTKUXg4ei9Q9xd
jjoXDTYlSvectRoQeKoQTSMUywh55iszWqcUS0yvdyGGMGAU7uq0X//14173x61V
azMCkkWiLVUNBZu64a2xnw7Kdeg9ssQdI00RY0iRnVby4rQmghJGqObcSDkebl7U
JFj72xgMmGhjREvYmrP3/4cmD9TNGSYvMyraaIT8W+irI+alrG7Qqmpm6PIt9kri
Yv1C/BlRguRhaK35S8KvaY0nAUHT8smYsmJBWAYI8a+QxLuVBfVDpuU7Cb5+KwoM
TcjfMYwcXBs6P/8OwUdKHaizmwVxEf39MpVZlQOcOPbvbPVwVjDisBspTukS72cT
yEibEo4Owtkwuqzw8RoB5zaTqrOKY5wlD6Ovvc6yq327ZjmgFx9L854FuRXeUKl1
jfYvqwO6OpbEL5wOdVWaYwprafNz94Z00NKSabBtFV7kIkWWkcBkH7I6Wvyxw5PP
fDcblc9xXTQbcPjxsjl+++W4butyu8fBsNJojgk0mETIh+3iUYAfDrgJXO4zJ0n9
Jqq1ridxkALJC/M06dJC2Wgzq7e+XBiFtqr8WEro/1ALzcWuN7V0plCT/IsP/5cl
N6Ztdddl1s4LINTBIaJ25Zuxxu5ga2XcEhmJCW6qIPOcVv+ZGBKkhKsSK2yog0j3
KSL+wRw6D+ifJiTX9+41B7Pmkdn+Bn1Tn0PxNDPJbiyUtuAUWfBu41V1BjRurON6
q8xXNYHkiJGyjCrBgN029FARpK6xHLdISlMr8H6jOzui0rsF9l9mclhIbPja7z7i
/22mFJDlz9hl5/xxflj50DjH92gRvf2iANV9rZl9GPrknEulG0nsmyORtV/Ox+m4
AJ9e89PboB2rNLeu/1LTkZFIjaQXugAxAoeaz1NJ4xwZ+cUx4Jkk37mSLJH+0tiG
f3GHG1rfEyWrOKnIaWZj6ixye73z/wFwu3wQQ/vBpS1JNHngGl7PPaLbSYxUiP8I
ML8MnhoYC0bOhuTx57yhKfiD5DkFK6qSI3IF69sV5ygr+hP/vbzU3JG8Qm9vdyz3
Rj2zzDfK/vtI48xYHfvUovULUFxoN/ZJ+pHTC9vvT6Bv2MqTXHa5iW2JbGEDmWKw
Q8O7VoG3O/5FwrnUOou2WGROf9bxWUl8PDvu5VVFlP1schQrcD0louaoRYcZHaRM
emsPWk6c0Kh+I9jB2JXE/IwClsNg+rt77hvUmfZDgpNs8UEli8Q37EjrhVxL3CH4
qLsjeXxUXsTumbtsIxw03WOnxPZUlUhewSC+97qlvMpcJdkJhN/tJzladvG2HNF6
jyB2dBzSR4Ej+0p2OSZFu7Zyt8XyXZCB8DhZ2cBvhDPy3YGfVEqO03sus8V/eftQ
6cX96Yb9xLsVgmQH1S/7jvxQYBsHevOHCaPne8mF+skFXb9cZqmaR61oCgfIpxdu
WAiSEZc0TfywjrSZmztIeWoczPE7Xa+5RNTBxGzMD/Cc4s1c2GyIibmYy1sygAbV
gn9733R7qZjUY37lZoGlNnSMgDycXQsRioH2mzpf0uM2yXLO3COTbYE8igG75aHK
SgRUYxIFPXc+ZyQxYEYykT2Dc5sSVrti4SZ2bDnr1DECZBYMcwi/qxc6avIR6e6i
AzCfDXI2BZdtyLcuu5DS9gl8LokYvv7P0yr9bNfd6WN39TftR6eIWNN6gozeGri4
h7+emX809rC9UMX21M8cLR979ES7bd2hP622Mh/ro8ANLZibsBiJIYkftkcrT4qd
AeiaSCSBX74pgRMafSYSgfnq8lUCmvjRBwopSnnfNjAINL2KzJYJbAB+TFbVcFU3
i3tWd4df867FgYpxoajomBxP+RdUHX2VNG+QaVQ/UFLnEVhydHH/t1EhMJ1w0dDn
BAuD1+4ib8OTZra8k8xnt7wiphrtiC27puzH/WMt3Yf1xBX4GcdKa4UXtImz1o4h
Hpu3Wmv95J86j80Wems7cGt5PcMPRXgrT47+zSuOn3FhlqIDkrTZDyiZVpm82WJi
jrB+FgbCC1aQoz0E3FTEFvOURMWPE1ovLyzKwKgxZAaN2GnvecSkyG8vA+G7teUe
Ukw0KYlj6O13QRhIffD98yfeUIKC3WNgMWIcH++4uEO92BWA2pdincBxLchgqL1/
2btuZxlhnF2YyqPXCLTYkgJ6omBnCVjVACgcxUur+ryES3/ZjbzDGHLZnZRG2bdz
+O7ucjjXMskQv/FPRSKtlCbboNFzTa++1EKkZZ691556yIMA1pNhFaiw6v1tzlqR
od6BCNJ8gBFAogq241nJjQPwvnXNJz4DDc6jhHmxQfhX0WQr+06fubW/KHTsndqB
F0UxevBUlOjRzvFo5hxtjaWpl7NqhvvES5lFM9Tcgi58Pdww+oTpiP0UDOn1lY9X
h/9LZwjGIzu7V66dti3QakwePrABP7YMYuIBY+ZSiYI/O/3mAUWaSbKnYsQTrGz7
LUMLwAqaOsTmib7bw6Yhs2ICtHaX2sHvKL8ua/D2Vu1A1yMflIJ1/56o9Y6sCO1B
jQ1NttN6hNo1DLWk9ysNgWKHj+7Uc/Bw3Le8WpdiifgE2XXXUC8Yjog+B5Sjs2/o
ir4OTUdy38B1W8QLTpfLUeb8dAbc2A1fczmQrJnwfbc4kITbk5nTSKe6ruI10GSl
aXY/TC2Oq9l2OrTYOPXpjgfUpsRboBnMOltLE88q9WiQIzdi3p72fJPsGzYTz3Vn
Osm+tuakIJnxa/edBNxu/3a0kZqzjgCu/vLo/YL5LeZxVGsRv2ZX7YWIrXwB35Vn
pciBAfaBjRULBo0tAoKOG4HgijpY7zFsbFDOnc3j/VnfNU633taeO4cqE4VK62wn
hGXfYMGNmYMNirNCKhSid+6wQ6vlEZZIpfUTv8o1A0UQ4fe5LwhGmXQ7X87Ebw1O
7WsQmCd+p57dsBrkaKCj825nt+XdqkbK+cLVspgLKuowOfHI5gptBnvPv1BZkGxE
omf96Kfai8qOZ288UhiECDmzUHzEUwK4WPTTRA809l24fSwNG3dZM6Mpn/v/WkTG
6ZFyHGz9gtL+JfHRWsuhA7KC3XKX/tVJFLPkksLAlLNaAjzlZbqeZgkkw7pAlBnz
Ezc6T6mZ1BLfKhSq51VCuAmbK2h3tIpLxRaOSinnWOLvw0kcko3z8SfIrRWvaZEL
ekRKBQ/zzQttGeQMfIrccm7s8XHDPD5bCGUp4LWMQoqobKZusuk18QSZ1/Jvjoh9
x2RRkKDFcJpY+LkLE5V+iyLyhD3na64fcR0xVTGHIPw2zV37jg/iXS1cwiJFBUZe
SwAvY3s7bNo28v6UsAnJRtNQwuFXAY331SQ5JOwrxkBOhiPxAkKwIhKMvb6QRWIh
pcN/EPf0BenI7g+BJbLv1Y1tNzocuuiTrEfl5nnMmkpRUt+KmECrxMkjkWo6LWs6
G9CRbM/lFQkLj0xRnbcPR+mLaBjrGoYuFXZ/4rJ+ehptbv9isl3K9vWNZtZI/z/q
tAO7DX4NDpgVFVneqTQJBN6NARkyYL76zBC+Qnh4KMkg/LkJ3qBFk1ahLNcWEjnh
m/xQO+GYfCjK98WK9ZbU1TDvPfl0d7Sg7IBsuvKmCPy68LE9ZpFZA3R3PXzGd8wE
fdsAXD0Yv1VzbZ/04g5iw4b95Uo49CCUFrWl8qn4sp1pmCsP/nbyDS6Vu9DXyaJk
p7CkfA6bhMeozAbRuIgh+nsErwcbYRR+cvS9fytR69skCCz3eNwyRcbkz/ZijBHs
PG3EJYahwgeflAuMQpsAdyK5MT7e/S9ge+U2e+ZMF/6rxdjUJr4SRBwX8t7T4JBY
pTFL/Ee/kNno+cBiqF0z3rjwwmaQgjolC0FSn6HyrBh1ZVbJdddinTYygWbinFhh
dJUqm2POj6eEhXItdFtBf4MddNpmQJXE2JMaFd509lxQseU5u2APQKWUG0YhRtJD
86wfssZ9c4Mad1kABe/R5hnSC4uxGNFKAr6Yui21OWpZK46C4uj3iMl1Bod6C1JX
HQMCMhXsG9xuICAzZEKKjGzaYf5+e6aXlsdJKAUNqv61UtDxRq68YkU9W7+kHdf5
/nf4QCtX+LC6sx57TA4VCMpEqOfYfPuxGl4lBRKYFbF/2L8lc9Ca/e35kvbH8e/f
v662/sKWF0auB7A6W8SZH8mXUlhdZN9tSYUjyI8lUMCIp+4gyq/IlDuIF0pNDvk6
xOZAOO7pyHuuvf462oU+O4Fa9GEaBx7pm3PoMKVLb/pGL6K822WBwF1zGYCTVE0b
y3aNEMWlg6I7/o30WxYoDF7CfxXDH9buZYkdCuY5msORSets29pODckYwQ38q8zj
M7sapz6w/YJNNptNnCZkMOjR8cHarx538MyLn8Z1fG71+3MCzShdmQVVlHm0Q0OP
MghGBciQmHY0KAeyGjBb20+vktzdYwzu+WzQm0iNZ65dHe3F9DqNTsUTTX1DGQt3
sY6QBUxOi49Q8DVuIKuRD3l/nTeXQfghb9B5UBX3uOKlnrwMmTets0XtbEsiarx9
zocef8serkWsdCHMPLsD0OQX0mV076hZy4AmsfDjDeZ9ZecGSa+86cSifYpMOlQz
iDeU+pilNMdfFVU3a7OnRXsiw9ebPLQhl+ZVcvXllFZFG5IvuTjNdqfjyEMS2tP8
/mKkmh3eN7U2kwMoZNCYMOqwMyrhVFhVdEw039K3uo6xImop9dhLxxmVOZrVi8uI
8v62cEvLnVIMxOTAIcajlXU+t7gxf87n+aJWeRtByxZOazonxRVN1wRi6ZtTfKs3
/UGWbNtTtZVftzIzHW4WEkEU4oQHAqZMOI8PWTCqOIprAqzGIovy+HPd+MdLKER/
8/rHHyp1rG/fy4kDCaGy+i93r4A0ffrqSg/1H+c3d8rXFy2pZRcOenJurAvt/wxk
4I+z+Dj1V2ym2S1enWXbjIl5Au37Ye1Ru8oV9pdz6vEQMDfdRk+lcXoTdiGjoyQ/
9fUpstlwowukza5Vnqwkuj99Qc6mIbMkBDfdAB2e4C3EpJ24FKSELqm3CEA3SLAR
IJpD0yuheD4ndsYDvwKYXYgLUR8K8a8Vr/QDUQW8zBHfkEMwxgDJPdaEwId2/TI2
3obx7yDxdDPVf4Q6KmyuCoJwoqWbgm6AskWSwNLn6ZSM8fUOD2YTvhznyzArY919
g4mYSZhmtPjVutj3cTk+JNrK1AvTfS9L5JDLP9ZuIHkrdDZGpYwMvSxWfBytNrL/
69vcVSF67CqsscgkqS3f+qo77+kAKvdib5WAIuLmGHQf03nBEcQvDeVe4St3YP3S
m4o2jd/6X0dDwNirdjmn3vJbBFtoleHAF2/rtTghHZECAD+BnqYkCJpxLJ/237sP
A5RkXZTfgk5882JXxq6gjB2esA9O4AeggUC4SzglshNatBBg3TfOwDX0zr88fmnE
EZjqNkvWFPOW0WHmlbLpcqa6iIXyoXn/cnJzqEyCwwqTl6z7egnlPTY9nBRurH8G
6TB/y4hSJV8YcHor/k6REEJkJzbHP08IhStdiMuI9bZqp67EYhkA8574qLqE/bX6
cas1TJ4YpQygvbNd2zgdJMbl//5yBTXUvcuAwoT8vBhisP2n/CIXRfpV0A84dkIH
jpzGBO5hRjwl33aAfBClp5nthBP5zJ/OSiS4fkbaovns8o3a/07S7BWHVoIhAcrD
xQ85tvTaieHjmnvpoafmDbCCQlwEj8mDRGA40NfZFsHyK82K/2EPlev3q+zWjaj/
4M/MCTDm0k37d0XF2xIV/DO0WxTjGlKx5y9PfGTFNS1w6ZjczinKewCZ8tvMKzmo
spJFjVKYYX8IJjvSEPctYFb/s6U++liAcJq8w0d+nLJXSSOKDkfEARVyz0/aCdn7
izwav10Z3a+H39nrF2LOd9cF8UTvnpFCgoX3CeYnj9OZEK5DPLQCU89KtU3CvUCF
KDpOpEqus+V67VEky+n6EiZs31pkvTKHNX6imQeoCiXmSAalZVnuCFuiyEP4Q4lp
QbNked6KF9edvsYSzLn+qilcxxJoShbuW8Mgi7cNOMDptoQU4SvS1LUo4SDTzG6s
VLHR43tMSv1uFkvQnaphVqBZfbtVUkvLgXw5lP3Uf5y18isBYUqzSK8OPqdOrEDh
E40f7af/e0QzusC2VTkAIGxq5vmO9i0lF+uaDhJQ/C2PNeJz/d7UY+q0W1+DyMZf
7aD2Yf5EpL8hsJzQcQLr5U5J+jLOedCPY+04ArJBTqPw6XhyaEaqf2EBkj2DDE8T
zaij9wARhyx1aBDNuPt8Vr6jwtm+ocTSfIovpyB/Ygq+U99tfaWSug5DGFFpfdA5
LJveZXsd806w9nfiWrrsZsMNJ+MrxcOUmCvjOX2erHp4MaUaFtuaMn9XUNAE7tHb
+51N8Rm3n6e6UvAq5pu5q94Ffl6WLUmbkw+3uVp+TH4DzaJiBd/G3uJV3x/z4F9Z
Nd7aNSCXHYZSazs+hdgOXRowXUJxfx+CtYJYp7Yl6LX/4an6jc9QQhov5gpMC22N
pYV9pa8Q5m8WE8OXIMGZyGANWQzIUDIazj2jFHMX2EVsC3epS+DLujhRYkNCn6V2
eOoA/B8e2kOOpVtKydaBUP1Nxgej4y7tINoW/WNjzkHdrw7rvxvGjeMaaT9q9jCZ
rjIDfu1c1CUUGVoF7/iumqhJ0HtVK53gxL4lSC0QkpU0O8DeDwwLzSMwL9LDgguY
TRol0V83eSdPqgRtBlRYbMPExBMSnDXWz3OEI2hF+Z6JOZVz6gQyGqoF8D0WAzVp
4Rxp+U+RTUSu9UBAywi76xrMomHpCL9b6QrwOAXYTX5lD4TH4yeh4vebJ62b835a
fqHxWA2hKFMY6ULJwJzFMZ/wccLksOMzanAwqK1zHRvlV5GVoKv1O5VO6kdSNzu6
HnF2SEuVeTWqX3yOjsqZ4Grb7h6RnpNGajagg7vvJRf6p8K5YF0JaZlDFOSdedbW
WEKI+qMEgLlQrdpzd5qxAXhWE71U2jQjULXvmgqJnjSZNCSmGe2tDeVoTw5YyV36
DNGt55Pu5KEvV5WRhMwUcxYxTNc8H4geY/r9KWVDcAnO7h+vA7sJlP6oBJk8Rs2n
oKEb4Ihdabse/b2yrMXXZojIuM+vw5sNyEiL9zvthtBKbW/BKM+VrVsFABkVuD+m
37LG+TlolKU4vp8kv0nDFCefzp9PJWkytdNuOTGTBglaOlIO7zQUF8+KsBgvyvKz
Gyc1An1bWf1EIXY7pOEa1DXR7+2O/BstLB+njdUvZdU7wD03lt4c4AW1gyrzEw97
P54spFTnLNijf/Nzv55H7WUWuJpGSEMLZ7v2APl1HksiAXGRlDzb3r4UJcLx1Xx4
S0N7fKr07BA46y9+QlTh8S7NQgWMCGelSKxfQiukssgf7sFU+yY8VyBEyC+7NOuD
NWe7YvG1KPrOflRpDYtFiKf8vyNFeX36UmYuoODdmOgn3YeFh2X9W0sX2pFLy9V+
sbB96ZwVga58DYKnrqnU+f0CCgi8CqXpo8Ns8w1Ux8DyQBXN88hJ+vhiIxbN5Re2
78w7fOCQLR+n0tny6XMwmtGCHNJHVv4esJ+3rPt7RmqL5dSlVShTkT11FRIbN0k+
xeGuQ5fyojQ1xN0ZZItrpY9oAY1TMl3fTMzWR+yhXgNc8ZXvdW+E9Lyrjgd8csk3
1Xrenm8BXhPbjl7+CTk1ho1DqTFcSlczfn7Eo8Tr8b5y6XpPgzGsPjpHi+KPzdvQ
wokDbMTj2VxteoOkOaoQHa7HMuexN71geMnxZDAlQs+j2C2Iax5C8YW+zEaw2AXl
aZt0Rcu3sReDHMmcnhVPkMAk8WMAC4Ijhf2AzmAUe5RnXmC9wVALb0JpXuV/CFyF
bc+COBQSqBehN+V9wXKGPkwY4dPvm4xMnEOakJ56plXusFK86IJFOTFsc8Lf7sNl
m8rENtsoyvbonLWzYC2wa0QJy8/Ol9NT9SpaCOIqBGXNK2MXxHNNnrWy2/HbWyn0
jaF9s9f5nLgjzOCtb2I8tk7NHZZ9NmJuhbDUANGaHldl2Sgt3Oph2c7VRA/0S6so
VbK4dJC5IZooHH3RUyLK4wrVt9oQTpQCXWaFm94b3xoWl1F4S5cdXnTdu9jXYdJy
rmEVZHG9l/23qJSaUcc943wr478AAz9fkntMzwZRsxmRwLgQdZnfGVzQ1CxWBgaS
5GwfXtDNn/Sbf1SjLubq9kKWGTfI+XzWSSYtdOcX+BviKJAnAvGRQSc190NtWyzu
BCfcANYpTRadAGe1TGhEbE92K3AIp4P/Lyd03Fzd61U62uolEFHE60SPdjg6G5Ev
yHm1DGfISAPtPuYACpKYM1DN2Oc28yiHiF35ISl8ixCmrUSIGb5YTy69wqpu3Kjs
2lgyR9lKtI9ZQkACyfyN10aJ282p4WtTouTmgofqU69Lrb9iCzq7sFVBwaFp213E
+fOWfZ1sVKA8pvPs+TYikolFFY9OkRy202qKU3cf47tVhooRYqf5G3UhYhiR1McU
dtZjHqmKz8FftUeJ1N/+DhzRug1CxblT5UZJ5vzMdwxfs9D5vY71aAlbW21NRhBz
An5ocW/PZCDJDD0A5MmbHFBKkfMtCdFZ52uHCsyeYyGpwJBQPpns2siloF3KjsHX
riB5ryyLn4KzMnsyCPkUf0jCr3fzhZOheO6yR+00V3EO8OVmjreT2WwYMFcVZU3I
pPrWnR2uAbPk0/azQkCBslbH760TsvSpyjLQBL22zEXcSn5W7pElqRuZoYhl8gAE
jkf3mnXmVc0BKl23p/Jq60NXGB/cze0USk5eQZ5cic+dpXTM7E/8arUgZLZEPiZz
BARlWrKB9yOV7KKWF/4cd3yvn9fitgPFJ4s9xFw1gxtXokwZcgvtXWJFmFY9o9py
fyspb5Cfjmndotl0Ev2OHrVle1L0nlh2saU5IKuXMO1mO1pga2+mCipc+zgW+CUF
20UqR1qt0GQtWn7tjbOF4Vh12VuwgPDaSeZIk2AwproDX68HNHWPjh71KHYJaN6k
FK69iS+whE4ZGCvhv7s+M20QDnu0kKSjlxMydvdNtop4S0VUy8u3jdFXNQ8ZI3Vf
MTuS1zdBMX2V4w/Gznfz4JUqQbvKlDjmtvGB2Ahc7feb43aDMK+98P9kP8sr3cIq
pcnmhiE62XtpitcrHFWwgOdYQcdSIZddc13UrJ61H/B+CnI/wAp/ItFJ5qcL2oPg
NmnN6meIGOhOw4fLNptynwp7xR2Ingb47WIos9HdN18qw1meU2hJa36H2syvp/Ha
vfV9eLLAEQRrg+5Cx4baVS6ttKjD1qXOIcrHfmxSW4T40lzXnkfruCAUPKVoPJjy
YmxES1e9m64S47r2i2AhhRGWEvhJzfXx2kWEw4fSAIRkCHnbn1nWczM22woIUG3j
wSk/fYwbvDBfGN8OxMwEaaqmQKFlx/QgPwl0lM5KU1aV38ELV/MGfQhMRO/pAUFs
lpb9sp1mgzV/nYP36gcHgScCJov5mplKDY2hu1mPZcDvPN4z7pRn0LlIY6oz2ctE
bxJaJcoljaVmgRIG6QPpombRJ5qF1SckBvKfpB3wdcMM/oU6KiYiwjfrJez881vW
HA1oxT6VXjlTzPdoLMxjPf+xuNBCRyvmtGyU91MBSy0OYjZqd1adKfbR95PALYHe
WvsXKVDkaMtffnir7WR/tqSZfFYffMrQ7bx+2Uje7wNV0Fr2OzTWfZgk3hGdziDG
j017HRSNMQIp/FA96IanXf0+SDT7byDXWw6uZGI76/8vHgN6AYtxDv8fw+K6BQsb
/rKWZHT8CMlwXb0+ZLONnaE0uaRc8ub3hmjtV/JPGIF91GMX0mKYSKa9pmTz2zps
NdCHOALHm1rzOC4Nmj4MQP1tAqN5LF1V0DFFjLxo6nfaf9RvVM17RPitFOd3BNJU
H2aYi0rUzY2Eu/GaQkUvcQXIEZxxRdk8ROuD8MscbLZEVOfXXgNqB+AHgxKVIXCr
atMhCQhUyLjOYNiMJzzJcRW8cdGKhUiTJbCMYyKotSfMDLs4Ch99x8oaZeylTqLt
vhtgCV6vA5kXaYwC3b2uLcj+kdmBNNKd+OMcZx50Gm9osQC9x6hO6ANDS4c8415y
nr8JFiFFe8tnN/sjfmEIhBST1SOkgSDXizKSPTwKQsaDbFzCqivXvU0bw7v4gz5/
a0o46rF4Mf30jtWu9+8zM/E3gmw1HS8j5JFpsAmNWAQPlKiO1UEuC7qsflhX8gTO
3TvbQaVah4QzfenzziOg0T+O/k1gsg+A6zxSD5HzcDZLpkhUCFk/7ZOIcPdH30/0
E6Ku6OW+AnNLUpHrQJG8BFENzFP/N0UxTC9cb6Rs9XaYORKrzE9knhR0/GEn4FAz
DrHYJzMWaKcMDZukSzZ893r5KDCARXhQOZA+ajRnCliuyBvqE86USKMSdwzOqjdQ
FU0p6QyvmbemumDuZ9FlCO0Iw53BT47aJL3X2+QBimZCHDsonMkOB+cbC/qFFsyK
rTp977NBvGNWOyA1bEvfh/1lfMtapf9+tP2JqPyIXDA/4iqD8dulP3LX/fQZLEyN
Wgf1cz8WWwI35E8Q1mF6zt920+MJFIQdzWVqBhShyKqUVvBcgHTZf4bwC/jqpm/B
c2/mnDu57DaoON3Pk9hgRTWSGw7YOBZ9f1Y7wQB8eSZoIwGJ79+AUXAOOm+GDxIb
GKXcf6PHjO2pqxtq8XbhaJ+upnIup8B8qLGqO5rzgY1LsSQXoJlzvLke9gjQt1z/
WlhwqMFAJ99n+xOVeTt4dQaZJEqMU5dMIPLUFuh46jI73r0d3CAIiEt4Iz6jz3Gx
2DfKqThaIjo3aJfoMEtLtgjkvNEkOTy9LjO9fGBjPdFbP02DDxXrFz+Yhh89s2d9
Xx+tg/gE/VgLrSKjXnkvRvQxBPLhcrkJ+IRscg3WYbZbrQdrJ2YOlTZqjymLPmZG
CsAcxXNrr92hh3fYI9euVFQPLxeENK0jsu6Dyel7R964VflOiw0n5NOcS/6grGIS
dbMGZC5sjuZKhZ1ZygApSzgjukpsQwiiGoUHlyNBGNsh/xfwxPMYkE8f9AA1H2xU
kwstByS0nacB+ViKFTvCr9hQEGEPvMtjUydiomgED6wnXkoANKI56W7Qodm3PX/a
gB2ulory80QiBf6GST11Q5Nu5rcbVwlUK0rupu8joevFM8SHa/qTvJ6oBW49JTtP
R+0niM5caUMAetJvb21mpW+SKwxcrzKPFDkRdlu8B1pFc7PKv03HCHSb8Q2wwTdt
ZUMVO89bf46UtW5rPcCwjEXv++oX3FLZ1RnrrCrpg5tlcMlbWUxQQ00dCGS8Sd9r
9eFc57BOG8+qTECfFerf9sWg1sh2xSO4zh826GteNvbCwOubImyP1J3aU4KsOmDd
DVHvr7CiRxI2T51JQ8YS7XnggaQ1+bhWaSlb2lj2K2KLLOByvYBGIBfVIGPFP/V+
E5zBrR2rstu1oiPDy4k2A5t0oca7n0HTfnYAymZFIZtwAC9WRw/JqvuErW9zonh8
kLV8b3DxIX2De3GdsrqyAW5Vp6pEis8LXIi14i3n4ULkNsUswDOaBl+rXgBwpKj/
/hiHSBCJEh+VgkzKQJ2NUsBeLIfVfu3FBIoJA1Rf/+GY7OCkuF0Dd+nSNFZotH9A
tu2nZB3xSpW9Tkc0vGRaamtpPsKA0HUE4/XNia7cdLDevqMEGMgrA4xSm/zMZgU6
S1EpCp2nF6ziQmrRe3lF9fI3iLQwYLZYK/N8/+Jip+eQyqrNKl36j3oD437nk+Q0
GVkOkXZuNcQ438tBYYz+N8aULpVspKM6ESFZQi7XSAYKNiHIf8+SM6T/oDbtXL+8
Ni8jaTujH27DwINm9MGmF859PdT1EP3yzrSXJXzxLRQEqosxuuqY4NHJkLVhbfvj
uHijIURbIryl+BbnxbY0atniYnuwgZW+n+Kv/V63HpkL5lXgFdE8VlccdViYgMgN
81hHBqX41YgpHB4hvRyFcFyk3iGNK7Uuh5z9qsewnzpMbaxsrV0akzYqT0QHaM70
OTI1GhZdcrp/7uORebbnC1YzVI2S2aAZxejx0k4cK8YGSkjQcBq46AoT9gF8uGir
fnQwtDu2RUMKIsNSSDq0Mu/EixLFIr0J9SSSMNL0ub560bERx4hXwIav8I7/VS5O
P1KRGz/DkwCF+aQctOae86tWIStpafuysBnrECk/w1EeCreJ6vvCeU6RQEJ6lPCc
h/BXDcYe8XQi4iTV6pPY6N1x3sWbfS4Josq5gT5XNa9G3ucOxkmbMaVrlpHUP0Rm
DixJ1RK4ik0asjlKdPn4U8fpefuh3RUzo6GZGCfXiE2B6HPk8h5Oz0QwieZNAK5h
+qVOT7N2oOdMZOdEF7nzf6d3UXaK2v1uFUxW1s5YkymYx2dhYoyOgZVHyQCHrwhk
H/rYx8zpCUFqnRhFuYI2ts+FtPt2/w4ot/6V7YyPfK8TnV9axaiiWmqvZ9l/Yok8
vPiAQO9LVhNWx7bDmBvkyFYv6c35UbNGx8TnooFMKVsf/NpyWCcmx8tX/5/viKqx
mMfNfYCPraEZj7DrNpQSy1jT0G6YsI04JaC8YyjkL5jayOF9RwpT/PSiSdx1buVJ
v2XNLDtldIVz7IPuapj4DLIuLVvMw05gAIpsvhZGimwBR+oWRdQAD9ATC/zIvgRS
VX40eA6KFebE8a79alMe48oUgeWmG9nX5W066Og2xuQ271za89y81yXlbklYmVJ/
uDelo0DVDL1hHsfbcI29CHLvN6o7ig423rqqoxyuckT+2A/iYR1mRrrhc/h9LEU5
JhK2fV1qDuvmsT3JM3B7Bnu1QhWd5dQXKtJQbFCz8b539+i9SUR5OR/4Oi+CFKmV
mbnWp/Wx0HBm3rDrHHtvdLCsZjLbr1kJbG5p99ooI+JKyiAntjKJmUVQ7QqUC/Ee
pr+2sF/3O7IRv2XhgbLJ0f9gQ1MKj78dY395TJrJtNaNie1mco1mVkvc3ZIrHErj
DJRTFLZZ79qbAB1IgvnrSNPTEF82NLbrQNPeI7BpdzA/ry4koxEUBwCXvuKOrgTn
J6MUe/OMpB/wbx/v1llcmZmV2E0JvNRoA5AcguZc/uyNrv5/7BwflwNk50CcCLvd
/OJTjnxyxI9VIVvjAV//yjUq/EpUvu+NDZhxOkIDGLaidRoAE8jdWHNkML6crrkI
o/W0pcptTHaSs8/rGhqeFhde8HEMBTTUUTxdEmeS67G3Wi5u2QDNbtTOCQBlLeku
IPVkuPKPGGL3jgbH0gF6Li5CtH4vZtF04fPK6BHgVG+fWmsZPP534wGgt0BtUnGJ
BJj73OZRomXk4P1Ihk0mX4003XxIkSuBh80NCn9tizgeH7vb4I5+o/wGFte8I3hF
Ze5y/WtjWbfd4Gwrtg7QyoWfq1jCgabr+40vPwAx1jD0wcDzUNp/VI1HdNLimRC+
RDX8GydoEzmJpKddKp9cs4q66tWrHPf3sEjdzncqavlqOdJ1eHQmagr5C5eUofGs
vAzbI072yWzHE5GIk/0K0YLCF6DRNFApZwNdjyKKowW32OpxAF6fAvOyFRh5nPpM
YATD6acgSI6OB0Hzm1hcl2O07AerTe30Mk58JC9TuVbbo25yJOzUuXydIg1sDMmW
JP3DmU3w9luzTze7LaL4eI48DL/k4k6xVpUiQrckinNJFx9t537ugwnWww+47Rkl
1uhTjpjLh08X4qQpLfxj+6Z6AkpN24+DYuOfVuXZZBQCFoMmN/AplMA/S1yT0CCf
ioG0SQ1dft+MdEv+gYiXnJ9AWVf1Ji/YD25W3B+TQxKDhmUYPB+rRIfV55ykqLwX
A9FHOSKJp+kAJ1Pjvq+R6obs3OYbvlXgjRzD+hQb4wSTOUqn31cD2dGyWPMZ8UZc
rL9uTEEXGWM7us2p2TuxNqlaePgisjaXl0LsE/M6nAEDmeFPspppLEjaCDfOS23c
AgOTNfHes5Cu7aTwA1cyASLA6s+eUcLOOWr3SrmuL9/5dwZv4scY7pb5gKhYKNcM
OMjmwt9x31sMNduOs9CWj5erHB7E/oMKYDj8wvO+4O7603PIFqYNTHcAdxBWXL2k
Cc6UfUjOdX6KTtdKfHwUYlHw9rpFjbSPZmbvKbS6i73V8KKrOGf7CstHXghgyM92
pTCc8wvhWsksJaSsPjVQEi+J/e3At2/vzqBrdAa+LeoexKuhDmf5DCVwgOp1SdBy
Lm53byyU/kMSWcma4jXjg98j7wnO0wiXurAOFynKrH5hmStmqgLz6y4UeVxY+oeY
MynGB5EovlPdx+Nk3rcHiyui22p8ZSCmub0UY0ces+qVzTQ9QL5CrKNk8ZFFl74r
f+g4a/YQ0PO6VsYI+YI28hjq+TI6eBlIB4eQG/HI2Hxyf5aDftWrIJXUGJyqNbk6
nyvY857aYgUJSwAxjvHYovi+4BsV5pWQxIXW//3WnZvZqaLE/iRve/H0bYLxjamv
rcXDRAGAQKyhBrf/KkRjd2zRqDNMiZux3bbQVNENfzLfvzQIw/bZMsNkPpZgVtma
6/37L+leykBevD4ksfVNmWQEiTufs+1CfFjGBM1vUJ6F6WxbaHrSsJsv9nrYgidG
/sDm/uQLKWjBq3rUXRNK87iaSiDSbB5ZCWDjgNO4ZqUB83EDXA+4t5LPsCXvskK4
ktG0RDHXBEKmqgBR6qJifzf1ncm6tyltGEqowEjKkOQCIsH5STSOpoNNxxzmMCzT
dYENzGDOqv6m1mND2qTZhCjVZUE9+cdmOY/Tajn3/CcuBKTqyBOBE185MbD6wsOP
8RgPHgZ4i1GUZslA3cneYoRPcEeTNqxfuFNHnSTo1nDIsyp+CWcS/lKG4uH8A4hq
+qQQRWl16k8Yv/RolH3+tbfnIQ+wCRBzBiyGV8Y3P5QK8seZgHBHYUd94VocLzNJ
ZUTOGH1iGvIES8YQZduVGaKvHh24L+S0ZRzYbbBM9/h9SDPA4PLzYVYmskEH2EHb
rtBs21QWAxbwRUrwINTon8xn2fqD9y8knRJttBjbbhlNUTOJgm4uhcvCDGKzZ94m
94YNHjPjrLSiiskD8TWlozKI1qnZHbf4roc+WFNDSE+JJUWDSI1wTopr+Deq3WaA
wt89LBP0fqTj4doB6I793xP987yTBQkyXVgYGRrWCj2y/hn177O8BZj0MtJIKmSn
DNgwdS5rKYWNLuWYe8a7X2p6AJA0GcI4ons/36wEx54klBL9DDxXVw0+Yn5tVFke
iyx2CGTZrJXfLNTbafpg97IMWu3fkOyAFYMvGMcDXLi4hdL/EGmQmK6GR1A7pFat
sGhDzfr417XdXBSl/VM5T3ovjTVS/065H+1vdQLzV3KaHO3EvXU2fYgMmALKVgYv
eOOgPbVjoiGLik7DKgWOdehaIeLmjtCM5K6i/tBPdpSTFNHJJgB/AdwvsmPKTmB3
ybCzvTZhDWov5YUgrFzVPMPLaHWXSKwNod17dHXnyxfhJrec92DRcHokUNquz+yk
wKyeIp6ShafN5jpIzzUub3XMOLo1Mb/x9fhYAIRu59FB3nf12S9HOlgp88Zq27eK
QR4XNAi0M8U3+DSmOLmQD6t7ECFcFdhN6r/y/NbzZE1WbFXDoCVdO8gK7wMN8ou0
uIhU+ik+N9AhNTFPLrtUANu5ADqaq7PcVLRVTgLP8fdhsspJ95ZAiDlTU7Atrg7Q
RO0ob4lv+A9qhzMCFCeWNJuSdps0XiesVOj3Cy7Vtnt+vfHV11pk3K2UL2gTC2fn
ASVb+mBTNRezNeaerIVpGuWCpq0Vl3rWapFz+xXfsQAIpq3YoJ+XVIPXk2NFd0wK
7DrHbFWoZXoSrv9jtTIGCS7XfIWgh3MRXpTYLl/3aXv6GnmHlypKOREHldtA9gy7
yX0JV9qxNzK5btsShUQU2A6hzlemIHTIvr1Mslx+XpwPyUnRaLNrwJnMOv19aImB
n7vNE1k/vez7g9ZXgNfUUmmdrqChX2AAfrVpjKTODm5mRimQ8jN743kGTt0Mgd4m
Y7B5CxofDr5Or4Wp2UA7oI9s1K3ywLi6sR7XvaPHau5m6itQHBKKmW4b4ctJhEmh
SX/EQwoEE4KcrjI3YqmzIVZkBsSpya+HfjmJ0xkgbOJuAfnGAIgvFLT7HMqP0Vsh
KkLuWjWh2WNW9wlyZeKcS52t217yAkZLxrL5uAlNcA3tDXdnUWxb+Tt0LH39IpDV
5J+gbndg1MKQr/GTFtwFCcWsUUjK6A7GxTSX0k0bBK4Xe5/ZJxXtQFcaBKS82f1i
NyGibN/hnoPdxRVqqTCA7AibgFxT5RIjNOwv2CGXNsWTOxQdE+inn9KbKbN1qeuI
JjmqGusLj4iYFsUs4LcgCO8IKTnYCYUnA8MSfR98wqSiVDYSGzWI2hMph4ezqX3x
R1pjk5Uxovtk5T16PNrry5KgYWpMznvEdiaWvQSloE28z1yCQLxrwt6Hb8I0hlnJ
GqX3CzjD2saDyn6/VUaaE16NtyvIgw9JPJeczHVXVXuD5oMDoBDFdV9l7IzzZFgh
WgQ+zIAsm2b/D5z5uv8G+7gOw88JfxkOJz021nOheSKzagW4PXgi8ngdDcas6Ar2
aGAIpfCm7V3lrItwwyCeGVmsYyFhI9fKeXH3pDX39XJHN2Di2css2tMl42ftBYin
dtDwT/do/WYh5I5CSSd1J83t3vOyXcW/tYNmhY4QbuDg+HdnJ7317ShDLrOeCv03
solJd8dMyB1HHZt9BDObe/Ov9AIz6WBSlRS07uRSFyllXI4TH5BJae3BfPRdmecu
Oelkc2jNt6rLTWyyoALUcqu6nkmJWTlMmH1Ik/rNTyl+nYzvJZ2b5PaLsU+7OmOM
DElNUUL9Gycia1i8qMD7q0opY3fM4YwN92Vu7vlMkbEQjEEUx8D3XhjD2+0g5rAb
Uby42lgxl8aVSwEYaUuufCP6Tl/KPMeYi4+SUaGThld00hYeyODna5tePi35k+Zl
QigJVgA5QUUBXGWg2u+xeKVITHrrmp/8tijuOU4+hS14/gZNT91L9ojrnAPVgHjn
eMAG4EZuDseNgz+2cOlkh7YrP93b3S6YVnJzxmso8YJt9bNhVSxb2ddHoYdMIKwD
wWKjGQ2PzO+qWxZLljU6Xi/qk0vxJ5bcnWtwuX/giEIgkO5hliiY0kGgy7tLTX2a
ovNABF9okqnb/AYnXC7OBjpSpNV+zFYqT1ZgDBwxrSjO4MX9CV5/Qyvrd6Jkt1iz
v7Pq6MzjgfL7ADUll4ETNFkausTirqFUVE64Go/3L1s32Rl8SSdEVh4h6oKHkBjo
6lDNgCepWbtSDfHY4+xZg7f7qhv/BhEZ+gts9OnPKcAZbluCs8HWYrQc5G8SQr9t
277FMJAtmXI0QKaPdCXto3FIjo8OXIOl5kYSEMXE/3xdmsvPZvXa4lGiTySX4TsV
roV5bHfwfxmrTgwN1socW+Lv52BTsruqV+0han7n3tLmgUDEIqREHxQOQMjL1EU7
b3+C+KeG1I7KyxH49AOvtJeiRSSnaRhJiN8ggUkqysUT2nh5z3eibio0IJeN0d2U
vQH4fOgjPHMJQdZ7nOlnprYQ8GqyxlHAu+6K0Enn5vJnfTjm55Hmic2p7bjJQ7fQ
/6FbKBKSZ1gffkFWMXpVGUh0YqUilfsSedLGBZpZLwFO18UjQzbq92eRCVgPwG6S
r5v2M/dVaVCuidGx1ilzdFnhAZOoRy1hC0qLpF+g9mWH3TAiV94O4zJBbc/PEhTm
7CsYHWs4+3sx03hTj7KZpKcI8TNBPxk213ViOORk1cTii9J9caO0bDTETM+53Bwh
ihM6IL303bq6nW89U7PQ6OxRM0pI002w9s6tpzq8pcYl6KTKkP7dKHILqDnEKsF2
V7OOudRdnd7MVjMA0/XrdCwWrK1lL9UfgJJdg2uKCHoEdJtOcYd9gFU1jf/U4t9B
RKkqfsrhUfOtrAVaOC8kKMkGzwMoPe/DAnaUSHtpaMs1iQgRU5shh7slrhbie6LI
7oYulWUlyT0NTol5/UK2a8HD9asmYSm3g+o5nQtiYMH2scayfjGiZO+juOrunyLq
eAUQt6KxTf5OVB77oR5j4VILDeH5975iDXpPcxPgTKgsQZzV2Kxpq8MjTWBUBtQp
WRLIilG0klB83xlyAxAWJmDSQZchfePCIqWcBBKTSRMJPnCpmZN/z0xDJKU9xbf5
1pk+DVoXqhB+3siagloywz57h8kwIczne9jhOGLvblcHb+scXnCmE+w+FClzvPm0
L/nq5TnyB7qeT2vzt0vVDfpR6FgJx8pnEdwCD4GXjL2lQ4+9wC09TKl62CN+wxkw
eoHj4d8pHGNkJ766h34nNRo/HzsWpg0vt0HzMQM52SiXLjjzWTxSd9/ajHGxY6C9
30gGfGntlOflbI6hlpTs6WIhfT4RoRT4raKIcsyV0OMmVAvH2bR3zaOsWIFSfHET
H5+YwLfxApRy4h8aPTChEQcF2u1ufsT/h7Gc8I6sjYXRk/ISsq5DHxuN7CwYKaEb
XhJ1jZTjdB9SSw1R/x8yQU2NMDfoJACwj9NUGYDx+tS/+RNfozJZPKHMBF9zEg+k
c3R1XLPThg0yheo+DK0nQaaCwbS4jG+ebl+l961pdUgFabBUTR/gwe1INvCTYW3r
sK/a/FrmgVlb2znSCZw5DFBJ+zeETAxqZRG+b3jgfckAOgMgupfpnrA8N9qR2HTC
GY6ADilzhAQDIPnCjy0ZkvKHn8Ouh+SU0kuGn6ivO2KJHsc7seOh0fFqm05AqxvC
SwQaKytMngDa9lfwnY/tdc+sx1/C5BqKME+xWsApecuITYr5uHFWUjKmuNAejK7U
m98cHwko9i0omIXrU2Lb3We2v4he3DTpQpAZ28PasBWcQmvZqKEWAb5WNJu/GRE1
DW1RyYu6BhKjKaMCb3BdgL71j4AsDAvddfgH9cATmJuw2JCQxAWt01TaHQQFRLLj
XVSVqEJtlYvFmvQpaOTbtgoLUDtc4OqTMszgAGs/s9LrZXSdZGePAaM5fqpEY4xC
7BLaDlkUBy4hqvGYk9O+aT4t2a63grGIcF0RPWAdSdBZEkRE0axgQChGxzKnVw4d
V65q4zQgIq5g3oTcNNi6JN9GuYjuDHLEGNFD7PTSbFS3+OT+2X+tSjZCu4tL5GKH
MDR9jgHY/isoH2deXBrkffvAZbwAD60viuW8EY5+KJrMt8YRXYKXJupnvWisAANQ
jOFJZ4yy6f6ni0TEjxXXodMVlu9i/GAws4cARI95Ey4Up6tdFSiQfCQEPq89pDaq
m+7Ft4TtWrbwMYu2BlXcgWbCF5tDmZVl1gaNiPBetqXymE4ihvaOTOG0Q+Vi9pDZ
Ku2vA0zUDBFTkXK5e8SO24whaCLUyM0nuyPo62Tc71cO/NBUMTUkguBfLeQH6kr0
/IlCTZ9uv7a6lzSKyIDKK6nuOwPQFRShAS5JpHT/ewnlelUgLdgjJWYHKc1XClfN
GCnlzOPq5wisgR3aBY3Agh7LjuX++MAHT5gBOFK3rM+eZuQ+QeJhyFnGeASdSnCt
eMVMndDLEOXD9jKdr1sus4oGxflttIZlX4Btnkk9KzNaa+iLvu/tBzAY+rJAFC3y
RuzzpMfbY25forawOpKn+SkFS1sPIqh250OOIutKEf+DtOavD4vljyYpKVE3ilQW
4VdmTYIX/55mAt2bcp5dIctMixPGVSjaeu3sL5jKmPKGthKxRMRZ2KPXpCKsHmdO
x/bL2QaiaTM9oDZaEmWWelePLNYZGH8b9mRO3o8WtFov/hOZIew5X16W68RPi+aH
Aiez/gZ76otqEqV0pHVzR8aWywW1R/5Og7WwURpECmJj8BXwXM3mHewCxwjQXM5a
p2X0JvxJY1lYg0nKEEGgT3q+gVpEBDNYnDWdpqmphmzzKlB0+UqI7LlttSrBVY/s
UxEUhbAWGOmLGPG0aifDCE6OrM5OwQCHuTY2eKN7L57IxsY924hJdSaS27Hfy4D/
d/1XvaLWnW9BzJ04oFC8XPmqbWbgz+0qAkeR+kKGK5kDL2E2I1ZcpNoURs+h2ane
tQlJQtsIlNgxpX5eQgC4SZzHZqjHfOpC2bIc0w1GaWlgPn5bOhDzl4/xOrFkE1XA
5EeM7gEBi1hhldKS/LPGgTmB2sXoTmUgWMxVGJnowxQXG2EmyuctVINnYH/0qZ4T
AqDrHSZ/z6BoYc1m92nnDyeqXjfOlNJaHTVN/C+kc4ORBLZrCvFzGiU8LJZae9cS
+T8+zpuLX1/ujCqkxRtoDJbtD7kqQclgoEALsRgmoDFQ9kwTdLmOjOhdsoEJJ2z6
z7KXpdUdvaZCq7ABqGqhY1A4siMftheWSxelYhoO0NeNIzgYqckhPRNAxNTTTDgi
fZGRnYOLNNJJdr9lItxmxK5/SPoOZ2EygzPBLq+p0LUkWAYzLAMdLlkNBQa7kAsr
O2JLz8faJwmfMbJSyGBfz0+xrR8KoafLV3IoQtrmM6Ny2nGyHAmdYRk++3cZfnzO
21Jg0g5bNLvVx/daf2FvqTYA9+jXQwOUUJIuWJm6E/sldnBM5m4wX+lPfG9Yr7ra
zpNtxOyLayS9d1mCRvo0fl45k2A3CPNskJCjQ7Op7ZpEqPKwWp+0iKn4/331XFPP
AhCabGTLS+joeMxI3XWARkkVA9PIFKIeJ7nkugHlkDbCBVENhNqx7JZu8R9YcTF6
R3G/U94jPXiNYnrgj1UqPmFCzCZkqwZH8ZfwqCS639LMaPwf5C6Oo3u5Ed78+FDC
sOxWaP5Vhk1/O/ZE//mE+S+C8PtXFJ09a3VVlZ7hDCO+9Pkmmstp+84MirnkcCVi
x6NjUkrK2Tdxm6VvbbPqJoO5xsxcgUuyFs/xajrhCsjefbQmhmuANSnwmnSMu/Ig
svug1g6jH4andavcFYBrn6tPS/FHdT+wWvq0/fP2ELl6YWTVSAs8U/aaetVB36OK
T3LRiuFv4yEFt9NmPgZBkbYgFCaUpcrXq90DcQtxMazkbd1sCKWwztyeEoR8prU6
BtsF+1XJLv1iiCnsJ2EfxCL4WkbP1gCJpFukunOSi9xJXGmdB4zyNRJWlJHkBxFE
CHBygZ2tMV0dQxvD7QdrKwmo5dxCYX9XW3SlP8FsH5Y3dxMY3+U1R5IiwNxHmlI+
G9Fys15iQFJ2lZ/SNk0kzg==
`pragma protect end_protected
