// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XDZVCQah7hz9kukQ0geBdg6vcRg46dU5wZrcO8VN6eSeokJOv3ahJbdFSp0ahdfR
lgcdsoIk6L/VrE3NaJEtNxBd/orsnprXvTDSFPclQcU8OkswjCkIEmGSf/day9jK
ROz1l4GvTMnKLxxIx2wuuxOhyp29Iuh0REPB9P5D3vU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3104)
jlQv+QV08XrsVU+K9hVMhbg1VsJznJyBT1s2hvaFoflTWxcA4x6OqllAr7tSIee3
8MWGGpNJJ6ZMb4/6pVcnBjpwOFpTJqa9lIqCYIXTsyLpj4kDuKmjAgom1JYJPwJ+
zq9Z90xSAcKz6i8vyKglLo6k9EwSLdptT3RyYGnCOphb08jbrfjvbxV+LN102ZXw
HTX+YMTPhjmcJR3VFV/SZIcvv0U8DCQYkFmDKf/PnICyy28iR7q2zo8yvXWXaZGt
5KmVbk+7gh9Eih3Hk/QzgtrlndEvo98/WboBnvbl/2xW0r6gnC8hHBiLVeuWGsu2
oTxZ8FrJ1sLLQ88x6+Np90xg60K3ZvmIC2ygs1RerhuNHndFmXTi3Arir7XPylAP
SmxkyumGzslQaR9zRyMcuG49xGsOoZzyOac7lxroJk+Fg8RUt3lEQOr0PTKQu4IE
CEAALoSWDMMW4OwGju4yv990Hlx4V58xVQFEJOkZeTejHVjEtHbbSDHLAxfrx68h
4LwIBntXs/ADjLyEBqGVr42v5dC3XfqwP5o0YLPbwpywf9MFvO5D206hJqB0FZR7
Z2QczmFUdLNPETyFr3uakg9cikAX6dnmFFkoSAbGb43P2tdRdTcY/ZW29IELmxcA
dXXY6NaowTZV4BDT+fsqTouOWSXU+h8z3ZvSg5SIrlBhp6lzOjBtTD8pYCAM93Cc
FkoRltVGLf9ST3aWOkEcyaUBu6cSYN+GqShihbowHe9+L1yKVYJfhoyWQaN17G17
ouStpKtjv2wiUmKERsE6tvXXGMr39ORz4NhpJdIVGrPVb4a9BtjAYJIX69RZGLjQ
XRcDO/UV96NZUYMZeAJ3VDtYGMWewjbe2g8poqHqpjTtP6YYPhcbaE7v+/GB4etP
kOsya/5yz+Ss6m+sbneRTxA8vNSRQZfbxlgX6is8WLCzfT/7dx6CjraY8Nyc9npm
iBaWIJbulUL+0cLnKvhWyjw/AWj/Z17UIWPfJIqezxkduRTdYLH/eVxPmVXqXvOC
oXJbQENg6XESVOaqgiJptkJX+4LjqS6/ygjf0TnmXkH7PLbSENgj0G1mb4yHydrf
QxaaYgcMRBq73jQenORogyR+0710BS6i/4ntBmXURvB8+mbE1FwVoFSCIrZc9FTx
wlA3AsYqsZFbSPmAGxdYwoIZFhhb9ONqsAdpz5Pk22R2OKAMIAqOoNFgEnsoxhTq
8kvWSoeFpWXzbNKyPEo0tZNGi7VazdE4wOPDBvsRydS7bXoWMVCvnyGfWYUOMpYm
k5Rzta5vvsneP31LltqnXh1MCME3l7ADqKfRzt7Jqklzg/GJZE7RZBhB1vLWbZUV
4MOLblBz7xC1mhSWosFz93dgVK/wI9T+IEZLvNii/LQtSPr9/2NQ/22lFlU2OOvp
lTjkB38Iv6UOnaQb7DpVrTKPTmCJXX4+XOOKeDO/ANFXfWActcwsVeq1QJYTL8hB
nibmuRycP+OAo46skn5e2/riPkXhKhr+XU5U9toTuLw807GnmctN5jsUYkZUpmom
B2jYwDMpY2gCwLHnUwSk3b34yQ3oX9iMiSO0pP3yeAO7RydFfXMJ+DtY/cLJFx6Y
yu4YObSQAeYpov+uCovsOB1Mgokc752mrs3LRT93q4E7RTz5xYS0fCrFtwlyUxaz
WpW78VZfLjsZCg+iHe/4GEtJKiw+fHAiPRHZXUKa7OgwQHQyBvAX0p5uCmh17ujJ
Wgs4B0vWXMlBUiSkMlaJhhAuFzm/2qNFhl836Bu9hpzUt0Tlv6O9rx+ymof1ViSe
toly5kUaDMOAvTBLLYDnQu92uHUYF+04gC1i7Nfk42d7gQ8f17fTlX0+FOT58+jV
XSYHSIpMeHTUFRMsNny7I0KItV7Z7ia6j0Qqvk9WtREeMynJzAUJiemmxsJ8x0wO
2V4Xbt6rDkc7ymmBgtEAhHXLthgza+uEogpJ5YqWbDObxVfh7AcysP44fsE2UjCM
k1Gk7pPL/v+wxfccaDZi7GciKoDD7Ow/ZXW+ZdfXmq1aLuzNBr/oTGgauyWzrZZX
kWJ4Dt/bpnWP1PJB6Ras44ukPCIxvIbJjh3O9bw6lqshd08/hcHQ+u8bSuxp3YSW
uehWvoVSA/z5wa0KjbNaxFVZxMsOcxJN3HWwCP+UMlRwTTuBMNMQtHGJa+gVU8e7
gUzPk97MBaysaZEurvAjelnCqnnhnN5/oF4ZZD9eJ2YaZXOjwfECCTjJBjyA395f
VHtNxq9hRfiS5k6AFiAftI0gSMGEec9Zxcs4v5qXTUDF0KX+0ScNikNCt9/efN51
4djicIdmXUZoD8+ya/CVaAM0WaQcmRExS8wDSA78/FveB/+DdhtP+MX+e3CEJkZs
Bm3fp2evQfvILWG+Q/CLkLVJa+qeohlmbbQcnhE/ZG+fup86PWaSdnWI7kpCXbla
xf8LZw820bsbb6Om4FvwBTErzXMAbpBvIKr3WNAETyEJAN+Ypfu8GG8/lS8/vT0K
v4pTvI+y3m5NY2Wb3b44yDJiQptuF43MdzyIOFvOZnuLRNmNJcx9PpQ5AvWG3HAA
9AwLabfWnMxu2HgbXfr/ynVGlSv2kWueB+kokIxblh00JD9vNWPhUNiaG78x1F0U
i/6LtdGOIj2C+mJ1tK8rynXLcnXlZnp0Tf8K4XXUeRqEJ6zjLCj8cwybWfPr+koW
jJhQcjwRIcf/BBw/F7mL+Y4dmFGCh6j3AhOFR6UGTJ/uVfnrZm/xzcELAqrsqHP3
oo5VXJ977Q00PgQmFDm9RnBwTuwhOsjhF/ML+nkgirMQb7hfNh9XMgzoeqkENVfJ
1S7bP6Nzpe6zWsPT9lmNygGiYIKyRDJqpanF4aS8cDm32FtTUDQNhALmoOoinwXU
39k1UezfYxxerUUHWjbNlAP2ib4oxAympafHWYRao225MgBlgZ1FauAlFcrN/bXf
HWZqfDftV3Acoue/+X9VP5JvguANraCI5v+9U1wlmS/emnv3arYZFtKahuimzxRu
7q6cERn6H747AxBtK0sXPf1AwdXgvSsXEDHTGGIfbgG2+8q7VXbSyn5ppaKmUoBh
dDhN7Qeo5q5eVY3qrE2o3N48krgAU3ZaSN1no/cfXVshIZlgxCLlBLth/xDz69sb
bqR8j1wYoy55EDJXynNsKDYh2oZtwtA8nq+UaLXHQ0bfpBMvcKkM+sMJbEKDPNr/
RKI7kz+hVbNhgTqIvLPTsdqMuJNp3MQy4GTT0PvG2Wic47X1t4GKi5qep/k6jVvj
ZVn2TFQezxhrskxgoIY1GNILJdrdDITYken5SCelrg7hQixOsfh2lfJ6Uw2eIPFM
0ZekowIAIm+Vrvbr+G0xdnRJg7RaDp9jHzjU6+8m6XirfLs1FfbhKG37cKw2jmLI
MWWMadGZTMgaGcjSE4jMTmj5xouMzafFmSz0m7oc8JV9yJKA4hbx868v7doqDRGK
td4LQBh45MhBDuRApHpZTLaqaVDzPT21VPuURAA8kN2i/3IHgMmysoLx3k3/xrB1
L9yTwSS2K/qWeXe2LTfpcO4o5jdxmlguxW021sa/j+vUhQ3qDYji962la4FJkdCD
JcFPKnE4aW2jdafOl7IHA9VFbST5HD8DLCfWQAFtzcIwBXNaGSC15oNz9cL8MGBA
h1ZC5ZrUIjBc4/KPO/jtoz8lHJrTDNBJAOWIlKg4xjJJJl8yXrUYoZjWgzhsjwr6
VK2NxgDrSsvlg2YoKxS6dbQr/zcU1hTJSOymkIcdoiEmavolaxD6kEPHj+cmgg5L
pRj8ee65T7f4xNFMCATc+sEeAl8EF02Ph+Tgq5LR0onVZt1qAzTn35r98fHd6Fmu
jRFCUL0js8MudCLXTMnn9Kyf+1qVdRgOV+VOTghONPeGs3BDAnI8QMePF4T8CCE7
CIGpJtKOARO2IzUgPP7U0RY3ZDYz6o62UVPZYDgEuiJ8HuZ8OKBmoBoPjnbCQnvM
sh6X19DjnxVT8uFf6tOv2SHFlTmk4/95Wy5ngifv88LB5qk8IlyJEcztwGE8DI3R
UjO3qOA/2irG6AoI7vJX8vtVKMWI7xmiNuV1ZCS7WFX/xbjWg1mTQhfJ/4ZbgrRK
ZXcAX6fPCjo0LVzQLuKMtMuaoUHTm/w5q0R7jnnHPlY=
`pragma protect end_protected
