��/  �Wu�ٽ���
�_/#N��(��Z�A�n��ݜ��O�d�ߎ	�Id�)?�5Q�	!5�%�P�JRw��w�k��5��ΰ��Q������z�i}[�T��M�ڟ��f�x/���+������������h�����u:zU�`�:<����Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9�㑉���f����^ӥ;Ǽ�Y�O����~�/�������uy���7x�I���\��R$�i�|2w�j��&�ކ����ZF�f���%^T��y
*�\�8����qi,�g��?����6:�sYoϿ�� 6��(|�iRnzș4�O4=�IGVڰI�o�so�{�Q|�4���fZ�:�G�%R�W�{���1ۼ^Q��>��I�N�ց�Ԑ�c_n�Lk4s	t�^Cܸt�}���-�X���]�������Ei���8�"I!s��j�hE�+��A'�<!��^t.l���(�"�0$�J �M '��7�G��(@���V�_Dފ�}s�Ω�A���cU�1�]A#Oy�ђ��mwxɌ9�?�g������U��*B�I���w�D�mrasn"��
_����
�'\:2uJz�O�a�si)��x��"��Hǫ�ɰd��]�'?�aj"~���Q��@ޜ���)V)d���s����"I&zp*h��M&��?��5��Q(T�����s<�z�ޤ��j�?��Uc�]������V�8F��#�m4���Dd��&(
�/�Sx�KgN�Ѽ�I�_I���a�p*L������:K)��T8bI�E� �c���)w�`�:@���6���S�<k�,�/�Ԥ���ZѮ���xE��~��!����4�A�QH�h�U.#���^̊��=�6f���<��Ô�rW�I���Gŉt>֧es���㤩rz5�\(�H��n�z>���X��`��8U�����L���%��)��ֶ
�n�pw6��
 �6�bk