// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fVrwwxuVcDBX66c/oDLKfy15J1usXomDlwOCDWMDBWqpdNavfBwvEWwBRHOPfKCw
BEbdeQmk5T2uGpzPkav6MIXt5uoNaaWIpC/FBluMTYMLbZEIy0eS++YqSLHdUktY
Z6tGPCq7N1Rgbybi3hfyv4t45l4xv0O4UAZei0SV4+k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8160)
2m33UF2LL5VpSFvfigvwM2GEXq6SB9q/qiN83dJJx3xAdbSBP9VKPOfD1iXGD52G
RA9YbcCORDIN4X98yu/lI4BJouqGnTyykiJkoAbRkWB5nkIF7v3qj9Jg8SAqePEB
dtvaemKNpkrX/q4YJ43ZqyU8FfoPROzR6lq3q+nnTX0mJMtoB+TyXmIvm6xE6rk/
g/SCO+27Q3S1uDDwhqTseW0jpTo42jkRCE2rotHSDIfoW08C9CfT7mCZ+vtHByJ0
l/ukrYqrtwnPKtt8ZcE3XpIABMIIJODxxSt5WX8hUzP46H7FkOM2WzTmwTmyElO1
bsybs7YHZ5WfupBhNDZROwF/YFz1u2rfQh7fJYTTPIWXRp2Wkq5AkOWt80QbHz+f
n2Imnyaxgte4vHVgrwDQvIhle1aqgZGVY4hVv39oE2ABVJu8LBGzS02dfPuxymst
b+85ZQTriT9WsuzQLO12KRCjE8JeFjlE2nuSpXSmQgfHWKgubf/eD4cTi8X8vXaa
4xY6Y5KwIjVNNqewp+r7NKlXw/hADiscxaBSMMD9zB9oTCeXm7raKNt9ZqrEv4T0
AS9jXLzAs/QpESGEnp0X6DzFTIx1qmX36XoDerTHYCn4q4uawA5MxLng++gsV78l
LGVU7QxamaC4nMzezNWFV+EJUj7eypykPNqFuWE4hTb3D2TOrnKWodwrUp1Ztf2j
aRgscvOeuG1HOIn+pZTenMoxOXZVeOyuDYY4d1cR6cEN2NC/V4Z7HU1fIK6y8EYI
6kq/nucsVSQefmxwHcYCbJhOABwLY5lT3OJtrmQQxx4NjwrimP8NxCLRprBjbvZm
8ZygK4IL+9FFZ7Rx0j66/QLQONdgp9qPr9jihm3c86Ogx2XRFOz5RKESLvj7X1W3
j2HNJKhqZGZYZPa5dX96yJsNvaM7qZPAlpf0w+hE/pNHRHyDzGJzvfk7+n/yjyYl
TPe3MSMUul49dvefcU8N/OIaHRg/zT0Eu8qu8iIui+ouGeUEQyNK69dUBOndfgnO
I/CikQ9NVMflqLWzBRik/w4WcqnDZ3A1S3zQ+amS04Oz7STHtc8QDgJOdCxrDejG
NBKa+vZlctnsDigcl3uT0DGjgZWpg+zBwNf87xr9G65X74kLRoBJdjLlhGcT7KDU
RodqZB1K7s6x70jv9/nQiXHwP+06q1eDBBoDPLM5dBfjL3771xLNyGV+3MWoH/Sc
QNiQVUBaODrd4H/Hq85a3IldJvBzlpqJrJbCCI3+voWwv+XRStzITUyI348qDsbt
ex5jyLYD23Uu05sVIjYAGfyZcM2XNKeiovQi1+Zuf0PKB3FcOL4kyOsgN7JbdumM
WSu0/2QIMn/JZAdvLnu+utAlJhiD/+ma+jy79nhiKHSHt4s0dqa4pabdOkwl+OgI
Nu8XlDWJLIVGVXVp+CYigItp72kTytEaZW2aIjqof0xuJ1UnRBNfuYzTeTZXfpac
Etj9JjlgRhy3EoDBvd+YFMKd3HaNx3n0ESopzzZtXazwaTvxPBdWyrTZSzYApzDG
32uo4y/S0chdFKUI2Jn0P5IUngWgz/zjulFje2Qe3beZdrIvhYzdqVX8kfhSTaMA
6UrPQkJ7v+eCpD8ZbSLR51HJNADAOuk7P3EnRLB2q8x9Q7s9E/j0lRo/FFxJeAoA
LJZPCkPS7gMV2gcSpaHGbM4U2mr2eRRKPc6XK9fzRvFXnO9+KYvTlZnp0ii/mdTh
+dH4hGBLWLZ292Guo5ttWWUb9YFTuWPYm23QuOe/3juQK+keLiOzBvtC/HuDdO4Z
PwxUsAkXOGkcGGMzmugECjWGg2LVZnVQwr7Rwh+eJG26ai6/nEealaznU3KkOdxH
fSYqOfUHXcC3S4AHmn/p5c6x/rkcQKUF6wRB3pC588tfgqIVH6rKsl0sCjrnUuyW
iVdUbxolZjdB1A3WxUNO8eiPc0NraJ71HZnyM9nzeXOSAGPGxhHwiplaCpi1Gd9u
f+oN0WUm/QjQwSgxO2+liBNOODn5dKUHWJELfvSlcmzu9igAgdxJH7CNm0RjHF6P
L2h4sJOrbEoNxEOWSftp1dlRhHRm1bY3PLZ0ux2karu/pKIkdWUvoGeY0UDL/OTz
BSpzQ7gCo2aT30eADZ5e1lntiV71IUyleny6bf44tfSFUjNjjKF0goNfNgiF05X8
4TrHiKccrHzLvzQP/A9dF2qTgOywooF4iesi46jB/QxUjCLnVlbmeqkwxUyASZiS
8+T7cLJBa7zVIy1H+6bBAYOVCYrrH4Xd2YWr2Eyp6V4tF2r8d4Q0vk5Ucmx4KVLk
5ga0zQQfuKLKIHFSbCRsN/jmxHtGHwJQJ8i8xkx1q5MMrZt+HMnOrOfck1q5Hx8V
gQy6AhwTcXmJvf6lR0DmdByopFYDCvJ+LZMgqozkBZ+78r+bvYaEKzepJijtY5gz
ZMlUyvf3G9IDVzl/G/qk79zbHyGznWz4jDjGMA1gsdbd/s3zjIiPh/UR8ONLxFkG
p84J3pwdk2JK1FMIlDRyVSwj/vwLhtcd33zDGgtduG8ihJrpOI8XmC4aPdlXAtOC
urhyKVh1u7eVLM5Hp2eJodp7haMytGemH2zjz8Z3YzxPfMqjAvE6/ZHg7oa1srr3
D7LrQEl7EOCeqT21j2uCINAdEqHikF+iAPGh1TnGFVTe8IrV9DUHIAMkRpDT/4oX
4nqD8MCbsqgkMPsqwJG8xTbl1cSBvJUliF0Qi/h903XQ27QX8bXVARv7dm+DLX+Z
Cxn00gt3Xs7WV5Tic1Q3g4a1uPOAAP6CMGB1yf0ugcgvo3kIrHaKd5fDgBVE+qx7
WhdcT5WKYS/S+sGloAsXcDrOQya2FttDq4ChWJdmmrNwqwGbo6ih4tSKOhVtJDQX
pyglfDtGgB1Flwo+tC3yV+6R6/bt8HKgBzlYeoE+8RizdOOEkN8FAi3cWC7ir9pY
Weha4hFVAgewsa1zUvMlnYtW7mOLdHYc4J121so+5k+3Gj4F3PR6r/ZvH1FK3v4G
59vLS0ulbvjFua+JKv63H+8p1SX7S4YwVeD5UXuy9tR2wd7gCt36cG7RUt9f1a1u
+1eFKmHyumJirs2BaXrBCnBGs0+klUiltV4P0h3TkjWxzwMrKvmoN7XVvL/OthmO
9syIRrcugKRfnS+v3x/qZZfP5GHPDNI2PSPiiv2up8EZeUcOTFEz12jxOrQrBJO2
cUgxYhZ9VDgKpx7aXhs2na9GQFSbbAugu1KH8Locdq+9shsjHqf8F3S/WDmhLeIY
Qh2mPi6T8WWua6ZkSBpgBaLsw95iNTGH8LwxQzuLwQbKkuHivqOZj90/l1O17XsH
8j89xLgxUn8ctb78gXjT4AW8owq7oXpeKdPn4HmjzDJmjL1P5o8Bue8K9qXnhgrO
+h4W3Zwx8Fd2eFXKtQpnNtvHZi8oApP4iANWrOgsXCEUI2UWBhdtAj3T++s3XWGU
2VKUFPLrWWdLyAnGPCRksTugGjrYQmKKDVmcRxWeWxFy70QLX/0Q4Ovz5wwHlIcE
7hkUD2QxUkmBS7LTdZ8z0XcnjVlHsc6fzaH8tNOZPdZQ5QeZVY94CxKW2uuK+I/b
WM5mi+gHNN0e7GLWTYft95h8/QAhOAF5XbhnQbd0lyVa0UK+dyo4PokBt7p5b8tH
C82gyHCvMuMQziNytwFfgQDU0NlQv+CxHQOpQ2QoUgpwLlrABTuv4qDx1pFx+k8k
jtx96D6qKc4xHG3ePW370pHz/Mts5B0Vt1WmjfYEeFhEUeA5cNZaNjvzFyVgHaFH
c7AvHR2ZC+LRR3L1QBwGNeCtGKUKtWEA4HsD0rIx5OibsK1AkhgVtRbNdtd4zNB5
jIBBNcZPkFMPDLAcIDBm+XPpcv47jfE1jEEf4pxxrOGdLOATt8n+M8pTF3m4iw+7
pax/lfBaJJEx7y2sWyAE6OIEDuly1QDO8vBDl4RO84saL7jLtahoZXElJ36IAbSY
/+Squ3otfS/2n1bb5+MS2nFSewcbP4+ioniGoVrY5hnH18Gn4pCHUjut99Ldeo6w
vCFohIz3vOQtOuBcdPlq9splVIAgj+zT3sDc1w4u95uoL4qxRIXAnqywWCMg72Gh
WPQ1f7zC9FcCRSfVBVrHw+OWb9XyZHmiY95Ds1CXeAzqoiaTEKcYUXF8G0eQ7bp5
O7Pd4Ou9SdiItyHcAOOVKtW0S1Wtz4YTXCKFixM4GN0RKaK7gJ24yOHcD8O8JWfA
38LHOVAhdDMoksQkCGDTKjeNRsF2FwUKGKGrIePIaxpS4cgKFRiZvLMLxBm5iOpg
8Zj90MBdqBsmVHruQJqJQljpDf0jKgrn1oAS69gKg7K6aGIw4RO4TemTkakH66u2
3URzu2TNbDBy+7sxw0kssKc/0icizVyBXPWzmUmIaF8ARgXJqjACkFTxvhDJhPHQ
7WTzjPuSoDZxhiSWG8saHWkFJ45IKvV1RGeGjiWBlhs7mGwmOvZ2i6XXuwTJRMM/
Fnudheaes2XfpgVJ1ponF2iPxzrgeAIXD3RavDrym9AOx748CGCjAs5PoOZc2EYP
cZLIFgDJcH2dY8IM5HetedgRcrR+6+EbKHedtGTQThMlH+10a1k7K70K+2YXxeH6
DpDLwhYH+eo2/x6N01w/iy6eRYxoPr999QoT/HMDbFb6gl3OaOA19sUQhX1BErfq
aemFGZWfdb0K2eV24dOLm5qEfg92Zl7BJTEpiRQR2rzhUjbnOihV8mnZ8267ekxy
8x6W+p5ILYu5VEp0GLDN6D0fl5/BF+uNls31HCojO9kYxbBdytvV7cTmLbepQzsn
KHx2K1KDUvf4wINwWOvQ+BXFOsvmRJpnYJiS2GHMAitNCB3sSFUy3KH13QxknDCx
Nl/iv5PKk0Rbumn43h4ultl90oyfT7Q1eLsPhhalGgInJSak0QqAUfpElmKHM3BW
wXTVD3DuadDc0t4JqE1zTbrqH2/rsl4Pj5vzMYtTaCjihCK+kaJqgJ863kqhmmkI
FGyR4nDVbncyDhYZJcK7VxzXGFuRBuvXCpB/CRZDbUl0BWfjkVn8dbPQ423+5kbi
lJCONTBxN4zRvPvp9Ha12vYlQn3htEMg5rurpIVDkATtvesTX7mFzQB+eTFIfMI5
t0UV9RsRysx579wwE74ZCqLpzYd56fCIv1YrH7iEiE4JgtG4kSkymlWXEqruoct7
wRROePLS3TJx7m78ml2g+M6EDDgx1V7aFMIIphYunWM6NJafvBXWJMO/SeuLeBhV
u80qf2/Y61mM2QxsQ4JU3SfUHAguJPADRwOk2XpJIV1tihtYMgZ6HUr6dMF3LOqU
UMbEv0A+6FubqA34wG0ySF8T8gj0B25QsJKBPoNf347SCrG0IVr//RBBHrboIcDV
VQYQVr7Z+DJVbDAT6ZbjxbmtqIgELRhw59cHgLc6QXgebvXtBOD4T/TKhQ7MJ9VK
SBDYopbSkHubUYWFXBcex7dT7TJw8Na9s77Kq2C8Upt9VvOD7qIcliogindQnelg
BGtjJMT4eEhMGjrbJn/aNrxWYd5QLCAeaZyioPAVEHN3RPQJINhHuq046bxkpav2
C6MPSrlSOfs55va2QguP010ZY+BbLUfsHqqKlcmJtasvH8Q7gNtok7ZENX5W0tRj
GUGDIfAcTAEFQ+UDcyTCiEJmN4i6EwjvDP28yjcL81kis2TH0qBHaNzXPEXMT3+x
tEQHR0/1cev/Jqul+P4GdygZ3pnqAA5sqgUvI3iWOkLX/SxjB8flySkbWLCTBTU/
T9ETKc0ttLiyanQASw3tphz6abeiuEtigzQIulLcfatp/4kOMNDovK1eD38nmyy8
R3iSQxjPmQOIe0WdDpUm+UQ++dUZKAvKFSMY4MPudxeGGsGmmblZNeUFITps2gfN
MZfZ2FDgjZo5vcW8mtGyzIcSD5DYg0mQWT6fNVgXF5Zu96J0VTpAfRkhPF0ACOTd
cZATuUEu33qbGAp8gaCqliVCGc5OPk96DeZ0Ati+lVQkxYDYu0iZPvaDywo8fHJr
nL/WCSDrV7d20DtavUiGMBRaTKlck9ZcRpDdbvc6VO+CxUPCG7Ke/fhf+yhhJ9gm
hIK5iOsT1ls0aCAezM8KEeWV5S2XfnoezOF33l6Xf0T6rO/f4E8YHvdJtRX/7FxR
30mQ6BZIPVJVFuJPfjj1QVg8JCthTiGQTjV/MVZArzZEInwrpc/qWxD3laI0JWXZ
K6BaN5/LY8Oxk20u0CAqCu0MNSDCsTzUvDRtmKg6ovg5lSOWpJjKQM6moJvuVK1D
LOLlYCW2M8TsW6M7WwbQKx9tYpvJaN5nFc/LydmwDxTTg7m8CCXh2lpGMbRVNtsu
OWfo3fc6e34R1ERuoW9byNqGeQUXzcLihpWUO+pqIgrbUtCtEa6hVersvK95/8Nd
snogp3JynMGdtnOgxwEO1qpe1A2OyagRuELKeLR1aCfkEkZMuYdDq0t5GcWwW7UH
ZPVK8bL0EGZvYwz+D630aSw0Gk4v3vhWM/ErFlayK0HYkQmNGJgORyrK9ZXTqi9z
MjpG2zI+ApRZCM4orSPdfVgSENGKBEDADhqsWB84mZkVcXrDOAEpC9AeteiDFKPZ
cBhXEu4DzqbTmOFxW364nvffPOLrzcCLoYAj9+9yN2vQxcXdoP249w+sHvqSyS1G
Cq+pWUMwiugINBGZf0Uqpr2f0BCBuy+Mhv0409jvX1ePM1KamnhOzcT3oWT3uFpx
4Kpj6grlDWk7tFMJLicM/4TjHcwKnJA7F85hhceHemvnLdDH9q7g146R3tkEGxsP
4yAaDhMiYRSkLtEEhTqhQoNGRysG28gcPU5u16qtvJhwC1pMpEn9cU6QNIr6fGPe
IifZAaJgsOL24ikrFhrYZ2dMgECJ3LQUgiCixeunEUQR3AHh3m5DWZPaoOf73Wdr
ku3+nX63wE06gRUiJvMA701gnId/jUcKpG/nHNdNFkvE4Zz0Hq0E7YUp111NdDdE
uvOZM3VW4ixw2Fp6oFFGiMIyNWq8N8l/QnHyXbmy2cAtzsYyOuAGh+IanGuBqSQk
5BksHU9+1jjI5sfwvJXL6dthPzLc6NEPwhnM85aH0rHJdTyG/jQEVfxyr94/k/+L
W4SBtPdZQhBGeo9c+SKEanY9hlv7ngwQzVPXBDFK73QJEsuqRw0mws+wDnScmqq2
LeZH6hTvjgj/wL3bPGea2xkAwRUWzfQHyP97nKBdGVH7A3EWKzPo0UUWKMIXEXJg
GBQ0dKFvy2jn5vxj+bXhC4V3xIWPpvhmdfCoSMMESlCBXJkrzwbZv9itvHA8An68
v0g2+VEezRYTGWQyn1loogTCOA5h0gkxNIEXNnueFEKj7Y+F5RKvqg9h4OP1Sj76
VF+gWVVmcbQv4RJm18qizAPGr9eiPiBKqpS6zDdkUAdlAiATeY59Mqndz6kBUdo8
QUTI7vbD9KsvZYX1cu2zCfiS07gPSBu83ZXNx5EdnYCi6EIl+zdeUyBLi8dL4Nli
XAt3wjhXcs+/X1HjJnCGWuoVJOrnVbnYIT1TGW4Fhj+cji7Kj/8da+4bmTH2n3wV
wdSPg3Ve2UOHq1g81RGB2i2zh4S9YUr7oXgZQcpwfVKb+nzSv8OeO3ei8MT7S04L
qn7qw/1zsVk95v+/ruyH95rq9AQg55tW/ml46v0vtdeIMXsiT75xKciX8rJ6bPRP
sLOV/N+q9IJGJl/KoB7P+JG7qWcwdZTSRdIkxObvZml/72GLYTEB4jk0C8uGSLGY
L6bK6Tk9T2FFeW+AZj9szv8catlY+N7v/eH8LY9rpUbTK7gd6UreYAmOJe2oXVCz
tuYRQxDNa5a8r9fP+YEoxGEdzD8u3q75DuE4ODIivRFwhi4V53WbY/WY5px6QVQM
KJP5p24ZW1XtusBJXzEhoX6RYRTmtO06eYvsZ62/E/A1us8MlTysijTCUj3de0wl
+069hKIY3LKq6oNCfUyt4gjL7X90cdqeZt/C5f2uo3VBA8URsD+KNxFY7P4F1mVW
hugwvTGxTQBh/hyqohtzyDTzu3zdkQQYxJkevKEVf/nxWZiwfhcSvu7IDEHiCSqw
G/5bIjga6uInsWhhoGTyLyqnsUkT1A+rP6+FCtOsFztLFsJrKekiI/qmdUGNs+Ru
vGFvHS+ippXQoJxhxBW8NBtweqCm5n/agrmtc9Vgb1kjR0wvFlbIcWbbQY16k2DR
MWRsRcwMRMGnbI3EiPK5Y8jLojt1iDisTPPPtQ4bFrSppow0PXf49mk/gOhPTogk
sG9Q+7MApgrd0xtF9kJNp5Ktcf11fNdz7OSK4LP5ExmRYdV+R/u0FVLYu+Q5Mugo
KtgEmWflfBibqog3HONYorALcEQQF1DfspE/VzOBSDyT1iOo0FJWRyrULy+ezG40
5aTaM4uJqCiOsAr7fYCdKd+ZjQ8C5gu9AdkFRqKvqA508CHE8i4Gmu+D1yAlgAfJ
c+4NcWUOQDHynxP6FxKNBp+7zcQ7nZGtDKQ11D3dux9CIHsefuxZetsWrWZfQK6R
cQLGboYc8dg0/D4UNONg09Gg/mB11yN7ZlT9ObrMo9HyTJaANJfBH91TSKzhU4z/
Bq32GD8mRgS1URqr1ROfqt/kjrNe5FJMP02E2XtzF1lJK3V+uliWijjV6xn0StSj
chfk1QikrDtyzIGkDJ7ofFeqp1RsydeTm1errGbxEbAtRINseO90Cmoc7sJeEccd
ephUInEZiklWu4PepM7sIvSID0FovaiT02Rk6sMC7K05nTjR7gSMmzGutcLjnA6L
xqeLgnlE+SCprBCpz+GLHZUvEyfVqLx4YdTMr9vPGXhuEQhGH5K/zGr/j2OnrKlD
DV/3+Hc8sQOUcPqs3qfjINc+QnDB/UMO7/528Fln1FxLGdBk4clYQ+hC62hP4E+r
vjcQxdiy725OiminAfa05pb63HpRxgKoMxgq2zpz1E47mT4CiZdRYqYWwrDZgLex
qe8aAMzzBxAPQPMGlzlpvXFxoPJ+XXSFP6xH6a0/E7RZj8bcDKOgHlfH17+SWo1H
7yUYPvFBGpoEYIh3uN0tS35e7yO5rLf4yiPhDw/lKt8GniW7tCbK7QL5I0Udx7uK
jDBugnEio2TB/TNIMoTpnm9P99iuTVp6+tvqLYuj871ckn99r5a1yqATS0nevDKa
0A2wN6RbfgV8OphIya01/U2fTdjQbhvXV5yrOp7AARhj4N3cIXXdc2/cndbxDi0o
CIZprFQHPM0r+NbsJZ2zKJyLry9yQTmNMKH27lnYQ0jL98JJBAXDbKD/rgMjS4rM
XGB77tsYCWb1mQ1Oo7t74wFqb0cppsO7UC5dSJEco87yk+f/KVUVpSHZgXIzZC1O
ek/2mPtUe7sUVV9xcy7dT14NaD2Yohl2GwsIMq0Gtj8II9QjdEk7E7V2J391835k
CaUZYAfJ+8zZ81d+EyqsVrvW5nsozCSZ90+sJa1YAClQXFTSxZ6adJKbn0QpUDqc
b1bStq/aOZVmuhpeI5AoLX8pBbiZ8aBnI12DjVzUPS3yFo8552F9PAuIh0b9Gk+r
s2c7H6DxVsBBaOr6s++D617Ho1V2yOm/rpsfaCozR/EIlxl6eBzqgK17GNv2Y+z/
xOU32EO0Ei/1qdlaMDfi7nhMwJ+VKPc7RcO8IIOBhFJlErOWoW/bHQj9Lnb0ssry
EsMqfvLAXwQSZTGko6Yr3AAOrNgLaeQdvXav6GeIe2WbHNJsZFDrCH2TBRsw5mEB
alMvT/atmfYvhSzrXj4MKPgY4P9oUH7BiNiW0oM6Y59SKpkumpCKX/b02SzVldsM
LDn3HdhxFnpHf2/S4U/ze/wYVs8oJkXwduecgl02ne8X7Vno87CuUUqtRsz+zWTb
yL1e3vfIeIG2Ad1fHn+1EMf8IUqEfk9Bpx4DjOo4eaP9c0JClicMM7HgcpixZThS
8sMEFXjcjGvcJtf7Yu7ZZn0CtfNH7H2NNEbUPG2DOxUSav0tKSQPTTl9I8JXZ4q9
6fbSrkhn8MRrZ6yjyuk/47DDDFuO4hjODiHDJwj36Q15HZf8rkdxINo6JE5eeDjI
ZYA7SoBryw10PmAryqC09AzRVdDO19Im9usehL1g5RUaAI923kEvUh8cztgcCBer
Sf+57muhEF4sVB0b+QWqrfmZ28n2y/Rz0d7ir3CwcGJ4td4/9fxa0lsAFfMOmQ1e
Bcwbl+3sYhgobwmQvuYKTSdrqFCTh4+kXGrWlR8j33Jb89v90OSj2nOBVWCsMBXU
mls/gHtjeDLRNOktibyPRLuE2fpfQTp57sGcqvSCzhVlmEuGHCvTwTJqo4dktmkS
lYFzZeJ01Yv3t2FzeDc2NaDnCpR6RuY2hWjhwujgzlMwMLkJJNhAaxMG5qtiSH08
WD8Y4XMC9gyeLS7ww4NH8ElyUZST/lyqUrrrMFbbfDxYkFrZaQ4W98f7xJ3Rz/vm
M6BCMXjzUDcvAlqTotjbdUEMs5Um0VMWb/llIO4pEwcvdRzF5qc6OzD947ims/Ly
ja0dzAO3GQoldz8V+tLN4z5gXD0YfO1w4bgp9REvbg6tUQY/ixvh6vAVX4C4A1jL
eikDTsSutTkiX0M2jqMF1zgfgtHeRaHYInoCJjmZlOCpJEe5FxT/luRtxy7/o318
WCoMeulkPTti3jYRHVeuxxPXWqt9XCN2hMx9BRIp3R40nlNEdabERIAQ06Oon39a
MX/0zk9Zl2t1uvAhcecnu5MWxSdEErKSdrx52sn3plmGbtlr8teADF+ssY36GOJA
3UcNOmyF3B1wZoV+6Aam1zryGyar0lvCPa0mrHeKW2Wgyly+3Y1C1VY6lGVG+bzA
G2uAgA/PEP20XADIQ7FExEZNEi4ryy0BGCIY9RkGoZsslAiXU23JKeMB0sxeggXx
`pragma protect end_protected
