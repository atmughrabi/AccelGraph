// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VBiAHxIlvY1S/OQymOooXj2lB+SUSQaUeWV5rm1x4nIdmofQu3s32yTvbHQCbG9R
nmFYDdSC5lE7Lv+vWivSV3eSYS7lky6pDhlUsZx+Al0t5cLj2WWD+lLVqce9foBp
d6t3gw28w7K5qMptmlMN6Jeb/7CQRq7Zb0zm5bkxeZU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8064)
htRZcunOGe+yFXvXM8wklaqdopNgHDRo3JUuQEyVYS//ImU1S6civDpHufD7it16
HLpkuIqmSLaM/lJgzfuw2oDH8vju5tUg+3oNDEL18G5bMRkWec/dnpfzuBJCxCXM
YHQ0qgZuFO4G3JqDA6TCjjLgalx5ga6sn3MGRNhgnwaHe8f0LEad88T/CallQw89
grITvLfZqb0FnjHyZdzZNUgowybijqL2OJajKAz076AxkyL6OdCFmU1O4lBNVHsW
ZwRS0iVrwP4jLjfXCJFoR8IzKAHelFlimUyuaxkdihqAvloLgbiGo50EE3un25Qd
o3o1rLVbFATh+LG6MnznR+mAxaQK58u/eIvNv9jImmui+l3jDg71HjandxFIFxA6
tWc5VlqbeBWV19PRSwqZI2xBwtWcF+KxicYiVuDWguA1jKIfUocMLxHW2aPozFKs
MnO2llRWOVBnDufI0/V3NGol/VecmqqU5qNMkGGF9K1v/VMlU+ArKNOCNNBIbc5k
F+0/pti2XpPRks+lDuVZcKMssi9WEsP8KWkXx2BMm0nqyKGJ3hQSulIkZf4DcV30
SStj34+hyvrcLNVO8ihtr338r++ZJQ4jV44t8Rt1hnn1BBY6wwPFml98yPxQAuhp
AnCu+4PDyqPZB/z6DXSoqjfy4bhZ4rixrVBy+Ii8SU07oo7U5z4q0iSlWpDpRBhv
qLWW30Kn7fmB6MT8fEFKWiM0tH2by9VHWSrMWq1jY3SmLLKnzgyhD3gR+e6fjYH+
jGtuqpXbndzCNOsSDmiL+bgEHBYU+Z41ZZ/gZ+S/RhqQ8fz0YIwPBKyXMVMK5rAe
Or1QSqPfhCel+3+n+KhKP5aKYfB4WFZO9mRsZyfUVQ18ohxYTpNb+VVbCbGDTaEy
fYmaY8+ji6D7J85ow8MSn7T4mIwvqFRwESjo+CkH73JaCfNNIWoSJ7npQoYpve9u
kEgv+Wls/Anw6a6tT56FgVo2sh5Fi6aUmN822g8eRYqVpZIAmqn0EEVpOOWTA546
Ier+z/vZT/uHuk4t3HNRSX5MbGriyLYYKeLRUPHn6veC/tWMEcdrUZf+ST0ko10R
tN1M+xRF9USDoE5lVrYn+ngK/6n+6/yr+DMghAsWcTTl0cC34ryPh5uMX2699/YV
c/37KgebgPHVhbEGt1ds5/Gzp90/002TPVy31MtvfzGH9GhDn32J6atoOVzlTngI
ye15XgnN1NYQesPpFEhefUFcp/U8dOpcm8KS2+u5pcdOpYCAgMJD3nkaeeQiC562
CoCNjOKiJsulh4WsRBW6gJ4W/pOj2tolXl+DKU4vknMxm8WiRdi/seSk1kWdhfaJ
5I/Mvbke/+KWXZMAtTr9yMsNcMk3URirBmCxRP8b8TPRQrYl/dc9ey+bEHvZcxqv
hOA2Nu2KOKx6AMiPeoaGSmUyDrc0oPQqXgmjnnTXCBpDhpGLMl3RMCAT2DSEN+Ta
FN7aGWCz0Dm9H5xJ1b9ydSSagbhdanCUJV5SI+es2pZSEBQWyylZzroIiZaKu78P
iUt5xBWMJrgwJzKNXtAzPCdd+dEihkWTnhf2qfrSRcvMSx+VkSuM4L7gBHjia41z
0MqbVcOEk6UAB6GpQSlAx4r76O6HhLnBq2LdCORsR1z+oK7iBO9hxTQBcKGcj4Oq
czvbcFjpH8L9G06hXOWiL+bSvj3kuGqqZmgM2eG8LpDeLk586CHTCby9u/O2C68a
lgFL2yeSic8yI/Cd4jLi0H/VkyjyXXf99YOdvBdOlRJ6u14ZdPxEc2vvav94xgPa
YvJKKdyDxPLnTQ1fTHxaLbGf+AZ15a04cXc2eFoJ04Rvb5hin1E9C2qOpEuyl3tV
9T4w25Hv40au5pNrmtr2RFi4an9Yj3jl1ExgHclrOaZTUP8C0q5qOLg2OwoJ3Fci
tWScW94NR17fRxQBnFw9PE/+A/RheJNWCEdwL+BmJJyYwwrQ3g4kdY9wXeyAI2Ta
PVs55GTQGacK3jR8DA+hohMBxwx+MOeD6iw98hgDF/xzmH4Sv8bLsqF7DiaX13IY
dqwwhd2dSap05iadZOPaTECgoct6h4F+h3fqT0Rctcup1/+PuExhkGwJ2UYtXvIo
81JqhASlC10nAxA6h3LMx5gR/avgP0PsPjxvEVOOMjskjCyGgUty+ndJ0yklZJdB
WW+hbgzMzNTTg9EeTa2EbxQr6qpl1B8z+sl3nQhfi+A8TD4jiGgIb42YSdI93ca5
GcEMrLsKfKqkVoD6FuAR4nKh+hk6XvBp6eNSjRPm5YomOx7jDjrtzmiuSyunprvl
dK0hATe8z0qe02Pt9REXheelozj/O2TiuvI+4AIX1g2NQY0pCC+R6LTG6R0Wworn
xHBFxd8erALXCLt4oyis8oGSOh51fFZ9Wfp+7IuYbAOrInxg+4D3NhQrNoQiNWHF
JtR0iHcu0S8VidBUIUl9GoCj0FaL6IGjraYV/eztjhoUCDp+jk+32j1YoOsiSVOn
2BVNu00e9NGO7pMowX72bHfv24/CfS81a4be6C3+uoM5C9DqYLwXFLDMzUbMUX3A
4B9shfc+2AQXtXtNS9JQKzpNfOzFk+j+rdc/E7DXCjI4MlNY4OJ9J8xAF2oVobG/
sNeiTcOWsyTbyiBGDpngtRIxWZtKep0C4nMReN85TokCtd+AFEnGbhcvaUzZGIIK
lli7OG6hx7vJey0MFUrPgV4CxRiqhAQ7qAn8DZMp0TdhN46e3vfzjT1N9gDYtDIK
m7DN2tDJq+r2elrwtMNsD34AqDTxnAg3h7DN4WZ2TDUYu5Tf+mDkWZy9At/bdF02
70b2sLCs7aPx8R356S3XkMIbMmGQ1AK9wS4ImKWfzbE+vlbl2E8UXi9KXvBC00nW
35DnPXS4Ddrp2ci2HX94f7eiGqVhqt1KPhG3NhtyxELltMoracDWlNfMnWNhqfHh
hI2ZptMFd/I/WG/NtbLeuFv4qq85oN66ZllzQj/eslaEKM1v7aR+77L55CamxQu4
k3PX3kxUh620KbdMsqRTqjW+uAAymfu8y/lU9QRVFLh8OK17Ykz5hu+S5JP/+eb3
ITP6ZQqcgsoB+UR/e9qxgs0GXLWoBAjYIcgqA9t8ts+8jwJajzVPOqA/4jvpRQsU
HgnwX7Uims2r4mHH0oZJStKo4x8svPVybjlkTJTohsEhbCUjch+raJ5bF1fBwaqu
WP8jkos3hLmV36uLYViEsEdvHAAWQnZ5JWPq5JO+2aW/oIe/Wc7UKh4a9YWrCNXF
MGEFfbzxi9No72JlDpq7VfeVZzbd6FZcrqcB8LLJeJErCE3qe8qaLlW86EkZu8pW
lZUs7uPfoUsaOQ7mft7UbMtRoojffeG+r5Vj0SvSmk/xKTeD1JqIYKcf1VFUx2we
btLdKMFJpnf3IaA8eyzDt30nxzstGAxNo3ILfy56WvaMVt505iyF276Kkgch1a2J
C1+Bsw23os+lrTpYoNv1w/kPygruxecEqvXMPJdA3BsAdZ7JFr4OIztzFcfsH29R
CC0J+Fo4KaSbudR4xdHucnmzq5UeKamBEmq775VsmTdINGzNf8S9lteVUfVYinTJ
YymxzJplnnnEkznc57uFZehl2nDpdaxEBDMiui55Ww7lDvSf1eyjolBHQKBEkW03
1N4R9ThHqx9J+MUmdZ9XbOc+X0mWygBdXl5S3enQefhydfOIX1n/deWkjz7yKE/U
HObVv6Vhph4wu4gKNsd85YGXdReJ8+ppOnOJjmh5Q3yu/9f5qPSPKvGkG1Y6fvJJ
d+CUi3K6CzMvF6z7NfR0U4OgD7Cafw5ZM9Ykaa0bfFM8vJ69998RTmGvs4K3VYzQ
oEaZ6b7gJttEnLB5x5uYPMk0MbWjd3TDFknQJcIDNCBBGLJ4gIk37GFsU59gQRIT
eF4ia3zuXMS1FCNFMHQCHskl9Uq92BS7/37mMg4woTPMxBLYLSWphoK8IScNAb2B
ab4z90jg2FbrJiW3eaDKNFvJOWg16u57rR7yKQiyege4KDoUvPLNp8Gi2JoIZWta
ebo1PQPjyuK80VBjGI/msXbWMZyU6rbseqTbSq0N4l2Mo7Kjk/EFTsegJLVZ8meA
qUY020rCub9CcpWSKCHTO+52TTQunNXm+glw5m2sRNreOvbp2DSjE4KBx2/IVYRD
mScIUVmkiiEeajl4vwpQLRapNyVEeFwPtIt7Luok/UZbYOgA3giTsiT8gmeGRjn9
GS9tNY/+vI8ea8TviWb9HHdIhxNaBqCJvJjxpJoP92zERkSJDs0TX3rfEHqfJQUY
DVU6m47UMpRbRZt5q8yxb/o7D1MzmTs5LLJra9/fVVqSZjcbQ5Rlx5jF2Xyc9ZRC
g+55/55I3HlDVqVLV77OPl/sGC2FIUmk1+FWIdpaIdCMXouu3cRG540cM0PUd+fw
cU0gRe+24c/ybfkslZW4N66ZLv9T/i1XLhfa5EHTaQ5G13URVPP0UFP6mIT3fpT6
z9qxXT8hHkaHxu4la7oNS6aq+d+qYVpzn5dimvQrRGnR/6+IE8Ybl8ZFtLFicAX7
foHoZyIVmoTQeaG2R66LFcgYSVke26jUYOhxPyuEIyz+60qbQrNMM5KHMM0CBVQ0
cGVgCFOg47W5ypBvv9mZL9tTMzb7NybGdezPUnU7ZFutWd6TWow3aLsN7R9LWkYI
a2e4WASVFxATWa5U0ZqUfokfA73/Nrscckm4o2X7MUFMpPbv32sJkPS444D9nLu8
lx6qyXrK6ON+bO2ksejg8Ybf1CwYOzfxMny7MrnSB/Xw55BKV+FbXu+plAG9y+Yr
l0Rah15i/a8GPmDzU/6YlmXRX/2QKNQD2zYfQdwDzFPpQD8oovCa9a7GuxoftQFx
WntKRl0ZMSFU/ieCfPDpPah5B6ffh8Ssn7/9dzn4plhwlMo9HunXWNnXNrbd8cAx
4go1gLdn1pCbrI9bpqRoDfT3U2CJf1U3Ub1/FwNX8FJn2jzxjF5mfvzllJP4hwyP
5uGsIdH355DbXq97aR7Mv3WFQvUc5hhd8nOdxoCXKD7II2DGnRRRXQu2ve7C7is4
MQrEiie/xrOW0aL+s2MRuaQf6v3E7VWg/UI/eUtvwXdDe9fFRbF/iOYDsuMu+6v4
2hgU6aqH2baZNEZrURKLWnkHBM8udMzoblxNy7sygK8+iMNFn89s693P3SQoFQxZ
sTnUkK5T1wLT6K9OsC/ruzOpVHiNw+ifG3UiVLKZV6Q41xx3et2qbn73HxVwV+6Q
ksZLmbCexcQoo1DIOlzOZdfnnFpCvc82eq30Co54ezBQOHCiRWHOjiACLOIeMb/5
DnuG2qT+Vnad4QuZzy20KNmvWjH6NCeg/P+JQbK7VVSTxWs/OcEmr9uluhZCHftQ
y2r2Y2ygsuVmJH/ePs3VxjtPK6yeDGJSvR2QXJBSv0z0zBEMqYPHZ4aLo2bKH/af
4QgzzxwzWO0yPd+QwvaqMDflNzvWyuPBOoxSZKozvRsgTox7AdCoBTJfXncdvr81
PKXti4cpmBZiw70qdiK5DVoZ7sAnnwb6JORciRPXRWMpG+FakMlWY6wByysGXpfu
FLh1EVqi+ZVSoq8CI9az898hI6GlBB/A34L3GNPrlE5MgKaINdX/xjrBNQpbIbun
12yjscbWa3R0OFTInmstQXM8eaLg0AB0PjzclZYFQPrVjgerQkmUlaqvrOcyerUq
SlHCYwieUQhPCTIvtxWeg7VVS56fC6OGprF0cdxxSpayPXtvJzp0v2BA1vnhuwTx
TZqcwVLbKO9AlAEfN5h8+ex9KsB9xXeOoVdkKUW26trXzj7JK+38YeXKI/fZycpB
b17hMPrUxojVnlHN+mLes3gt1HvHI7XEbSAqLqxXpXTta3i3//giXhXfskyAhqvg
K9E4rhef4PZPtGyd3zvorWzOSGqg665Pxh+3YR0HgpzV7ZPL8c37JQ5FnZfEPb2r
VU4ug7ms/pG7Yyprs+nGwJdrFyUqdpyaI7IMRMe69PF948BoQcqpUFbjrSXjAxKm
Tess6H9aUrWpGPs6oEqz9iuRSc7C1zyA+Esqb/3QdwTQlJLvFv1EL9SXA1mwkg2a
hfacfTRn6l0/yTsN3OYfryIgPqZ1ps2K4EKb4qjrDOEzHTE5TUgroNv17/jkZb+Y
x2YektH0+kyr2pCBVgsrUmdkAxR8kwfnR6vlTbXpNA/+HRBfx4imozVW5c6B6GNU
4VRgFg+0vGb/FHCDJpRtap7ZKoSzYgJp3snrON3DswkSvkAQqayx0p5tz/VQsXfv
Dqgw2PmlKLBaugluRlouF5FDfKNxjBtUvuUaYMABcvyPS6fld0S0Gn9wyB6oKvXh
/vfW8xLJlZHm8TQKVHxb7dSyRrBfyvWlL1VeGcMQ3W6P7siLPLCHzZ4vZm6ujkhi
ZeQ+VMfRYeNXq4EKZ7yRMuJqiSL/V0rsuKLpyQ62w33lXyFHUPZDNRoJeDBL0l09
b+VvV78xrMZJi76Ld0tMZ9EeJn8USX3ei/XcTVN9P2Q1lgVtAHPnKQ9qEj+BUZBy
Xv7xus2TQrakVGCPZbrlBg2OOT/mpdW7Yml4UjmlHC5K3085WWsWosXou4B1lCy1
9cNBJgxLGq3WChJqKQj9obQydWzx+bdHG52gzrB4x9GhpyH/eE+frUm10eqx0HxM
gnQPQumbTGDCTb1l7kuzv80ZmbKkH+Zw9PEyBCDiGagK6qAvBMiOu+0aAYwoNR9I
S83LbbCnDkuwhL63IfZs/ZY3uOFDo3Wicuf9sai8TBpsm5Dt2qo6RfbQHvEK09FK
f77b4yKbLUiz2f2aBvF3A4OYlJ4eEEvhr/iDthLmduYuslDyeViH45uL3WZQc6Rm
nio2h0S7CZm5iZxknHghk6WTQQmjuK4h/k7cKorWsKu4qEpIxm2+1kVR201/YxOE
srVKmUHiI9BNwD4F8qhcJpUo06UuUO7k0WoJ4kbNytnOmR5zx0gCVC0brqjzpBMI
Zewlj5LWnJ0O5/fitEtX/tqcQI4+NIYarqWUyYB1uO0V80Pt7f3YsKEdaYGgYWzp
HQs1kJAb9CJsanTkEnjXu3sph6VdsXZTOPNF2JLzJ5gRTH5/641lCQNMuFbD0LVP
fYqhmGLmsXEulEKyMmxqIbBlectPuOF9EJPRDDDio/6UikuFj7TCACU3OuoVx9/+
BYJVLBuxLYk8sAd9FeriJmJiB5/Ru7glR5eliUkt1zahy+sVoaIhigE6rsr0AF+3
OBTAgd9LtJovpxBh+TPUMZdVP+fRk8z8BZOujelor2ixd/eju7Alb8Mg+FosDGh2
yfGRkixQt7JM1nUjKU04JYyh4785ooJeYW4rVpxa8pfr3CyHQ+v6FM2AYUijGieV
oTXs2u3BQNS414rIFzVNccoGTEclSnHw36YS7cwocvwSTxTYoyXijXJlKuOUcFZa
rVvlZa0LP/WyLorycmQHgtAsw6t2n+rOMcuoEqjWvkRY0bwbtP4hqvqj6Dy7DfIN
pxasRuREBaf1XwdSYX3oC0ckYvlCUXD38Kh53axytwPyRACUMKmraKbNLqxfQm7U
i5IygprWoYrXb4bUA5x29MaIUnxvJ8Pw7Xv/80aT2pLClc2mbqgJdQDDaRm4/ov8
LnzmViSwbMmOH6YEAl+vIBiPknbYtmCW99EFgT5wpoREg9L99EM9bBw1jLS8cSPJ
2CanN+3Z9Wh81FH8PloL0u23zKEbgYv9CquN4tDjOjIwIO0peVE/Z7OvsyYUSppy
5fLv5hs6jsQlaIh5rAfmgUY7uyO/Gv7aKyWCYZMz333fHRx6rT0xRZBJJBOIqfX6
K/+mOLs3mXyfVsLYwjyjXDd9E4D22o497isN3WNvDyzjz+EE6KgAP3I9UMlIhk/S
/+Q+dTgJVLqRB5Lg6d4EcxAQCjAse+Bvdh9CtUvxiL0dwVYVYkGdZ8iusW5q88kN
1lvFuOYQF9rvI6Mtyd2kT2pwoN0cFWe4MnkljUmMd492LkMPEskESQcfcybs0/Fi
e27vP+BD2y7UGx2zY02NXHyysoOdw1fOIZHJk0GiCFdTeJOFwg6EmOB5Ye2kN1/L
J6kU/12aIClboKuLb74n3aiUU+KSk3LOPMfxUDJkoKG72PlR/YPWJWhAO+cefG/e
Wpd6gaOZyz4b1Y3pQ6YXKzrLHXgTGHldUbf91oexQKTrOdrXxckey/H14ss47IpA
gvO3sN5PgXqsaZnIAuUW6RCtnOmFL3yVJPWcQJaMozs5yym2UHZOGqvPJUZEEySO
+FEWeOGYw4Y/7sq8vtMBcxQcUExckIdKsh+T7+iSQjM32zCOXy20UUW6Cv/hNiCk
o4tm57eLNQI9jlBr19w0COOhh0uHhJ/K4is+bDMrHiz1eUTQJuJcvT0/GBzCZhM5
HbwsvfTR/NGu6UkoN9zx5uDVd2TrC6d8GNbe3+wgh9YVnh2JSaHsdQ1aKVyHpfqB
6yQ4N2wh6haF+ZcceBE78Xv9GE5U+XeWoogeYuoJ8fvmmpuDHidArKN4QDDY0DEh
w22h2H5Z10GHSeQTkuRpuQeAtTM0YtybaH26eUgK8sJEsGrlJuUqt8KGa7RbdJkV
yV2rpUzgYBNVLOV8nV+zx8PUdDaTiifEuNol/rEPkokyZ+4n3FsFVaR7IxK3SbDN
QtCJxEfURTcLzxw5HnHazeGIBndGrSr5Exdd2Yy5eSnMWifz1dpPEgj8lVhWzIkQ
CSDd/b4im8Cbhp2GbZNAnx69N9EZEJmoBVCq6FVQ0EhENTRW/VmGt4LaCCUEQHC+
XVS2bsGGAybv0DTA4YIFNf2GupXixgIg5tA3/b3WZu5Zz/p4KCRdGLeBcDjtg0Er
9sg+2YeLsr/5iFVmRXVK4yDId7HpEXJmEXL09envKyNPjQtcg495vZ62qnAH84el
cMTm8uN4RZwRdRbneyJ5NSGO8Hvjo3/0bucYZiKpRTVuMk93ZPW5fs5RcDK70hYa
5ABoccMBgDw21vtW3JmFX+nIH3ZcJIKIz3f55+XpsqvWC2MPpn84apC+oy6OYwhO
u6pa2AfbNDXxg3kR6bAUnIvILgujD4pUHG4fYm7LEJb780J5dcfEKSqHBvVrcOUE
X+jFPcZIWEEQuuF8G8GPJB+e3SxU1qREK+u3D/yN5VDwCLU/nWK85drTOyg+hAj7
WXDXtZ6fGeztnJ/TgWKpeFk6JCI/WXyt2c2E/PcAq72+aXvBg3X6vHS7M6V2pj2n
V8YZmzTxiLfjD8gFf2KcvJmTZE7rHoSHydfvQH21noGEz2461ZfnXnD2AXsHuMgT
LLfgddcnUece4ZMeBW2Hc/byOX6qvp6IbTnJuIMRusWKZQKvX6OmxgP4H3GvE03u
FTB7duH3LTGedlKNuWLPJSM76sczmg1m7WT2NK3E+Ifm/6XJbejFy23knx+LXxo2
M4pp83Yff87qVA84iCgPxrTlkSWE70wQJY5lcqSbQ7MveBNdFLKdASQX4JKwos2k
4Z1lqYu8tOqPPKm+r9i5VkIC+EDB0aWocEHRyLIrcHd3rZfmM3vPnUf5Ky1aEV5t
w+spQroXK5vvc4bZfuHbpLQlOv87gSBdqzI87I9exzrdJ2c/+HhHpaacQ0wtOOJ/
F5cqh97OpHHw8239ICs28EjdMe/tIXK+oEmR/DFplUKHcT5uMhFufp3JwUKJXDww
d+BuKBrs5LW3LCUlosHFazTPz2P1D2mpmsUX0hdKJGs4ENjt43xqGbmIw5zcIi9r
E9Wv0trxausHiDpKIRO05VW6B0Ef5Sml5kglg8VdyPEU/pUHS+hUK/AelFPC9acg
GjXUnhzO02dkiPwYZpkJtpzOeYETDorRDmk/8YOXIke804L04BhquUnSvqYPS18R
iSdLG+Fg5alqjh8pNa8vBKtmSuOQt8GHgdcnxIXVeDBUQy0x/Ss8yb9TSptQAlO9
2SEQjakugQKk67YYeuPAMf3W9jvTWvpJBS018jJE/0pASaJNkwp9zl/VnFLbU4Cl
tqWGdTul081vJC9EzHQwkcNwoNhv/CbUiAxRoGcp2f0ywpMW9Z3h9bjz53/xHqaH
Pbi4gWr9CZbJnGFDM+EqXZXqonzhKCFEWtBZaJNZD+j5DlKEcynhRrDRcsPf1b+/
oNzlrgAZtSWwGket4TR5HwYt+05+uUVll29zrrIRq1bCvjatk+ny0xR+EB7qmuxR
CWq1y8ITJwSOjB3kLqY8uwmlWGpbXTN79JdFzqTgl26dDmwPH0Enmc0G82caZgCZ
CVJCFz+feItIUzgJMtNTb2b+2DH11CvBpNF1IkkZ24Orr7W5px50THoTGE6t9Zh4
ZJGai+14262BA6xFBzz5JLb1qXxDiQBtI2zNkyrdnlYPa+pm4BJLi4dwrNlSeFiH
gslu6qjMFZUf3jCrHXQFQqWUuKKAPAboU3OTR/ljdpqtdZ7cMeum12Hwp29jQbqy
C9v7ysc27bb/B2dxlaI4r6VRtuwgqCcvC+9KaHs8ptmyRb3ewZCUXXw+712qQVqx
g5hHHZVXwCXCOb/9+BoeZ2c+bUajohEy3xQwAZocSEbtCVTt7aE16Jybi7AjJSa3
+/+Bz6WhfaC+LOwUCtEhH0P79hX/evsJ3uT4whIBLKFdgHpUoiSvjKKM6mQrmvu6
XsMWe2LZ+60CnOfD5eZ36Bdf3ER39iI3wXdZmaB3NhqhyTJ8ukv5kJ/sfpgNDxZ0
ff7oRQDzlIenxXlxWD6m6apVT3YDXM9hHShElWhE4QtxnwcG42/xLYbpCAlqaBHk
`pragma protect end_protected
