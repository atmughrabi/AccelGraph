// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qrqCIwVJGPObAmizd+rt8i0gUvszpkTBWnD6ksr4CZs2K4/PKnZdkCbeURE8WrqN
PfJ1c9w3G54Cdd7bQu6M38V4At34xtCimRaZsHNl6tw1eSca2UzKjvZQaj1Y88Xy
GWrIGqRiyDyPWIdoRde+YblbP/Ua2u81oosBPWwdQnA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28160)
DkkCu09G8Ne0CKgZghDy8RTg83FvNcAvPLl2DUSneX22KtvuRmNmTs0FqZIbbG5q
MghKRD6SQyaw/hhlXCBO8zFoTiTYp2xpN4h0ZsV7jmicvYWX6OldyF8Mm7KqAYK9
O65ckOtFHUiYtJ9ZRqxF5T8Or7R/boSGfsfScVAw67xPYv5A12yJIPyQpFOrt7Cj
kI9MB223mjfWPvKXRbHyMjaFRc1spToJSFzcvGZNBEAcMqKpg9UKWaO8X2n9D+Xq
gwrEktzsu6hAs8BG0bDEZK8fbCN37EV7JkaS20TDZ/wvY2hWMiVaPmDeXms/YuIS
Cm+emL7jOLSHHiTwh76iRVGbSqFVfy4dX58F65vLP0IE7cEiEKX/wdE5eECrJi+i
F6bcubCiqw8vujfnAOsHu8MSJoNSBajseclL77Na5oj/btJON3qAg5nvtSVheXyX
exgEb2g850XmrZYLUku81d7MvO3h5ORpjXx3eSQxjCYFTaJeU/fU99c1lfhWD1qb
/+5yA6h76u5PyPpbF7W6T1C/cWSkq9uoo9/MPUSfJW//4dOtT/Fesll5mal6P9Ur
WivZAvkzg9uk3CV7ySZyaEMwnHc46WcV0F/LtinrLuR/3Q4LZPutWKbQd//UFDQJ
Nz1kB+Xpx18RHUXzokcvYjyY5AcHWlfCffufX05Mc/zpihhPNJj7ShbO1bcdn1sC
W4yzGqiSZbuwJk/8EZfBXo9yzqeOO+b1VQnsRXyuvqE0YVmiMMLq+dsfcJE4oaz9
EZ5ATb8Ye4Hdr8oNt5AG5VT0Zzl6kzq6ODzNYhYOI0IBAAW9qWikEuuG1duQ1wf3
5kEAxNujzujlzyRKedBudZHhtWTc6Oe/BFZqBMNrPj4VFmS5sSB2YwOYopTOAAB1
YFlOCQX0oVXwz8Eh0JaXxZx9wdgHOGhQ15zSg+oymthJ67QKpZX2leuWCdPcsdmM
20ArUsp1/x2TpjF1qnqT1w2s5AeuKOJyxS53iV2Q58EwtINpLRRdO9eNLoHOSWk7
ktoCetgHpZkh4tfo1uWyfvJlM+srmOMXnE1AVJNLyc+2OfqUVhxBbbQJSZ+8E6AP
riMkebu44unbDpLshY7JVUchF59Ij8hPYNbpfd8IspNaHzJk1kRAE2w5xZfwuUzq
9/hcm+SMsF02edlMHBWQmo3AOayZMc6HrgEbtn7tv1XGltlq3sBuG/eKYUhHewjN
f0TgdmPMbKz70um0fRfDxp0Pp3p0jOy3aoyy/+DReBIU51CJhrV0XnJW4OybIpLG
B4GmYjrjc2GU815xj1gqTDWlmq870GnxYL08N7MlgHg3ZVD6e0TgY/5r10kUjnKC
6dWpiVZKTCpQ8zBq/DVJSc46A0RSI66q1iU88d3exq+OF51+ugEO9WXmv7yO+zHu
gBRGMtLFtoRQa8UFj4siay6nRS8YLq1I7b4hVdU4Mx5u2HbEUZBWQ1Ul11M82V3n
NBh0JHzKsGswt6a1K25rA36FdOSOHVQtuLMhpr8zJOqKFrFdDryW2Q+S8dYuGZ6m
8bPyma/rAdWaS0Z9UX/EmghuOkrZahLNW84V6ViO6jD5XAZa0G9gFKndKOkZh4aM
ABTJeoy+0lhlFi8OJPhd7oK3IvtiGOb40RiX6i9h4FlSwovMe4anqGEpur6VRbBZ
UynXErRSRnRfIrUwwehrdmX9LtLuLswWPa7+udXPxxSD1s0Fe9HQqP4R2p8EW8a2
mcvBmPVHq4OZ90PPa5mICDKojLHhiGhZ0BXSgfsfcn3SOWuiy+P6osbDUOTEkRLC
kOawTxNR7/9sLzweRxYYUmQxMxklmR0cOmKsyBoTxiXV4TDqDBZmMt8grkYRP3jG
YrS2KRfsBvMe8ERuNkB0OERFl6zg5s1K1R7wfxwSqYQFYErd+XFsNzSlaeZMRoj4
TikYILwPQnhHMZUkBrt51lZ2Ndl0NzaqMpl+ZP+CPRZIyJZXqTmsrPWGTomlxEtJ
cpptAEkYGW1D5TX4L/upQ/OpOh23TPJUamTBkH93pv9G/yT1Q10ea/BsN1IzawgA
5Lwiyhg34O8hzrHgnEsdAQDf2tBEtf/eOmWB6cF7QWVojNb7ZxYL1DedITXl5tIx
aRYcuSTLsbSqmQT4Orpw+2TAY3iUkOHJHYIKriS/mcY+fQJxjt32+h/arZkQMpG9
nf3hDqIoT4cWzpORLpGtQ54w4F/iW9Eq3eknxwYfwAqFqY/HrD2BakZvB9W9jhPl
Xn9q4rq1rRlJXOdab9rgqGHzlFTAjGsmwOpr0RtE0XT8SOLmh0agrtNvwW1Hm87Q
9lopn3Pc0Pt8GSs7VK5QS8vgRKjFJZxhjYfwp6pMwVUQRTDWzAnJbTZoQBgRcIUt
AgZ5JuFKbuziZ0dLvIZjQpCX671wQ3XUQQ8GwrdWneU9Sow0qFXt4EHbcbikXd+E
+XfxrPUSQktoQ3oyfr72rVY5AdyrxfN58kGmwOxxAJHKVraCm5LJY4nSjxRcnCM+
sOegOdycIQ56Ttbw0VID3psGsI+1oE+f6iDSeKZvIzZBXVxmtdAAsiBiGOzSl2hR
f6w3YNAVsk3xkBsb7Fi26tYhbzswRsNyzUieKicSTg+I1pwrRouabXsiBxbf5XLi
4gtnwVUwpVNlpo08MsP2UMDavsGPDWorLWnUslqww6YOVFDrsGypYUucVnYHQBG9
cBFdZZBbe4J6Php68B8SqHBW2V/V3yqxYHNKJBtyKDABkwVIfq+3/m0wJ0x2JnjI
3/xG27r2OlWoMg+ifCttY9qTrZcQloJVI8F97deWaLvRQKfrdNf8LZ9sbfZfOvpD
77zcSJzHcMr+LhWq2LY0TwvMjzVXboIS61HEoBnV/VMwryn6d4hlhrc3cMehxPKr
DtWFDeBegPcubEGxagiiuqll/Q6cS96VjqazUrk+Y+N9WiqNBG8OQ6NvP/z5hbgw
FdF1ZLfsiYkw+GifpspLaglgp7GEaVvFpUXBMW0WxPpcgcpqjufhvd5Df7sSi4kC
v+PuG/FOqxnKuoK3/jqUB0DSXVUhmIv+X/eBwDogYWZJUobTSFt+ESEXB3XlD1OX
NQ+9T7FCQgl3z+BsJFS58rECgEiifcd1vNdt9MFtpzSeLLQeUgl26h0rDoJQ6ovC
wijDcXTNPNOoAT90TnRjYkOtsbGoM3ayFx9VDTVjO48S8LGf6wsI3bzJRB08nTRH
mzMiw6zyyaJNS3K+zcYBiloree/V/tZquowRV2EcsKIbiRyCrOZjjfyIYIUaDSD7
04B5CVLBTQGrgJrQMcDqxhJH5ARLAXEb5s36eErV9x5iD2Gggja6ba3Joq/UaxDw
uE1RiHdAK8r6SEMUSZk9Szsx488SlgTOnFXEYOz1bWnU6jNnVkrd6ogfM5GDzKos
ImO69XWkJ9L0loZw2u7RAoweTNI7GFtVfpDGukWQ8jy0Y1DflCh62ZbKg+4SjW+U
ECof76oxVnzPIIftvwN0Rn015lIfxSLzexA/w2UruuGk7+uZkLW6z56D/bvJN3sz
nK4gtxZ5Vyy8D7ynbs/hE6jGAXMTZRDJkdiJppdjIrc9rWbcm/MuVBcNEFM3AXwj
QzUuImVCmRZZE6Fg9XUH++q7edcS0fUGKNQqX4N13ZV9KX7UxVREmo1ccChwfUHF
JtQF3yX0mJW6/75GDWTXPiIahWUyz+YhSXR4YfAlV8NhaBDd9CYabG6oEHeohgAR
cM9bzkJr9YzjBtmMrlgcZoV4Q0XD0gYEPoeV+e63v2yP+RvBIuLRFrRVRDr1eFEl
cFQ1mDnfyN0Ow8exrfKhR6Uu95ISPp850pHnDkRMGiReerohr4jdILEQvXAVx9vU
f6Tw+RI+3W2IW/SIQddjg8kV0mL/eBmy1bBLFrfyu0SH4QVRhXg/IGNjoZRZx3IR
s4sMo3iY3TZ39uAkx6m6bsOML58ir2UadXixtfO718ZdocUeI3SAhyRPMcVyslT8
LWrjuh2TGgkb7uZ1zUCzVuk1LFm08TW6l+pHGOHoV28YoIlKOnlnnSxrUGoF5D3l
DYZpxgJuOyxerWv/xBDP/BxSol5KhYkaVw77FjLcUR5uNlmPwD8OLtRQbGqoVAex
iFXGi79UZ6k77xWONAKmSyPcLEiiZ0vsW810Cb0oMf/dv5spUsHZpSjPDfnoOv1j
ToVJDBVMu3GBSe0mHzXoJgxmMa88Y02H7UrL5TdRZSqqv/AuRGpK1jJYbIMKxkv0
Xj0uuigFLMJANTINa9Le7SQobuhm04BIt/MULfGqOM5j83K4E01GH2sQxr0V/1Yl
VjngmrqTvqC6UOBUQxCJRIyluWAby8QoWzaieNntqA2pIB/okNn1yDjzE+h4DyLp
ZPs/0A15TT3bOfWZS4XbCkkGiTeDgXDQ1whIAFHGz/8T27G0pfsF1eWRWe+xc9St
mOPTtGJMQ1DVEbkHTRC/9rBy5zjbITss0EXVPOy0moMnhWOIPpse8NyEG5DG+428
OXQJjSiQ/HHv4K2vWK96pkKaexX9i7IIh9YHUz2TL8cYAlEeD21yqjZmyBlepE8P
GFnZJec52l2hJ1xkmjJO3B6B0jDOGnKW8KDTDQyi85xAnbqiBpqzNhU81KoVD67M
q3ICJS9juBAR6UamK8fKTa+7jTh9b1Jp5AYPc87Yla5kN59UPTnlaWsK4RRiGA9x
sAply1vsU/3gRhHeASLY5B+1UK4iyT5LNY00KdjPVhl0GaaCTdxuOzETHWV9Knhw
CW3jfgP3ckdc3oM+cWqMVcDgnxLfeOME+sKFAwHEdEIJidjmlowt2rvhaTIBUOCF
iCk0jF7tq43p7KPAuOPIC9x2lFt2pkaGIT3Nx2IoHpH315wMnlWPDyEhXsNx9lAO
CeSOLdwjAXIakpp/ZMSwn65Y1IHCAe+4RX3nL1DHnU3fEwTVZMNsJO44Z7xdG1hI
h554ZJNilVFAuKxOIdas/lnJjYCnn3XUBZcEiN7kzGv+JtfSVcTtlTSI50owg4CM
Z/1EgAGqEI5e6g3/HjLKa1ufBYVfEc+O5npcxFIwUj1MecKOVwYSv4tEma89IpwA
TXfhPzPRdexdbII+Ib7WAbExTz8Nbfm0pmdYfQzPVUCC9O44h2nxwiP1MqeEn7Gb
yhB5rGzUcDBH8vP1PTArY8opgHrC8oKW/2naWxo5gDYP28Uhkf5sBdOm5sLuRz7q
UZVmZasq6Jso4awzNPVFBpqQPqr2sg17NJgT2MVuMB0IIKadgYIB7o6jp3XPJ7Nh
U+3pK3W6wCwDeCIKwjhkFG8xLn4Li1phqsGCvFzb0gCzZvg8MfWQNJL/k+UcBpIC
Fod2AkALkE74iKwqNfO5d+Je6Hi50JwfqGSYX/foDNo5OYggmn27QG7aUcetoYGO
byZCDAGaxFhl+71bL0ndvpjzb03V99fu3PVFFmnHDbds+tdXHwIHKe4QCCms5vse
AcbaopDQ+82cuL/18QgpkZ7R2GeiI2MK48ggj6LCRdKHDsXrzlDr997yD8UlBksb
dtHA1fs+acYCA4GOUpCt0Pn6e6MCBtECBr5szBLZOfVTUl0Rldw2lhEZwQkE6RLT
lfJnjWiU79i3xsBFYnCw7twXdpdynHEgnKhNqW//ysV/OD2sdfdUdNrwWZxUQBw+
QFB6mbqO///1ODBCjpc9hxSCZ36xFiilomX/Cy2XSTFbjy+BOLjuoF8aZISIWucN
H5NNoSV1pTbNTT6ysO/jq6VO3iV5MPa9LOdqzbv7YzrhrjfC8w0v2kHYyic7Z2rn
/i+IVR+VMbaPOU/AFuWD46aDFWOY/S1Vsy9j5eRgUc4xQRl0FHLOmKEsC7Y/r2vA
4JllWx2h64SdjEftbCsC3jRRDZpQWOs21SJaSX2pVvJTX9O5N+r+zU6wTkU/Xqvf
ILxEVOvijAG+BWJ/nlCQCLAgPbyhdSgyYG1V5rpaLQkYjth7mskAWhv9HlzjC9KV
/+D9Fv+X8oJchuYaRwOHbgHwPspfucF0sGzU3sxl8cwTVfOjzQ3mp8juu6cNoK7k
mMBkvw2F/AlIYd3h7N/EHAgs15fiOg/7fk6EpIFKFarrHjMvVYICdGAcXsfNkJBd
xO5w/9KolOCufUqZLyP3L8X4Pj2Tgj4Vpj5hkufzx2dsew1VN8OeJWwldSEoGO9o
yoGdxCTa1+cctBSqaBjM6nv/q0bwUuzOIiKVdj3WX/lsCr6NG6fzxWe/fAA+o5ht
XL2odXAE5iSg0Hj2eu0vqTtcRpXgg1sDE9qlL1ZPFq253s8mZrBfvCimal/6YKI7
qaeJpRLyBs2MmIpumdKz330oEYz/Iff2sRGHoGr6K6tQ+X7HvBFeLvVqiGVGGPp4
P3Szt9xko6lcDPocK1na1DJxj6OhYHt7xGctBbJ9D9aDsRrZ11lBFQgfKTEIcrKb
qHhvXFrS5fMggmtPYzOljumPb3E0Zo/JpSzhhidpF3ZHE+xcRuHi6AXWOEhEhgle
Uo0GApUVVR5PoVXkgBEir6WbiauAVm/1iP5OdXJB9ieyqUGfwRfAXGRAvYIEp3pu
ey9gdqJaxslDDPVGqPnTFq+0nlGDo8ZCkI6qXOv/QWEMbphzRKM/Qe6/VUhfhvEu
ml5Isr68JJ2LVcmdhik77mngJhYiu05wRCBlTkyR1u4PsfFa5oJr8lsbm4rQZc8e
7cG9x5s7sc6TsjQoBq+GlGJAWvpETP+Uds7EpgstPOe+hGvuqfCbqkM9SG2du/AW
DzxNixefa+Jgg3kuKAV8q+EbB+hKwgEv7x3jVt29Sx46MuwZYV1jRpjqDESBQdNx
4eUfExWEzQ7XWxFV07JcZM/zWZj5UYn8MHoIXQX2N7NSGkwaK+5DMADR+z5GR+Ww
6KgDY+A2C2elL7cJl8rfZ4D/29KMxpKEv0CkK3Hl2upToCYCoUDCJqE2/QY55EQ1
l7ZkOzmPZ/Bi5vOyTkIiGDbA9l1LODeaFqHVCy3d5uxRjKmv4r/d6KnnyuS2WFHP
ldolsfD2/vVG6YQ/pJv5+h93bYu/KqiRsd1Mxrj1M9wKvzx9AaYAVIFCtPBlOriJ
UZBL574/QSw2HQbJzH6ZRoXAhaOv2xkJY4NX770NNhOywx7DB965voRsXEgtOWQL
Zfj0ulBj6Dcszw0QShg/tXG7vuWlcUqgJQOmVJph+/gpE2q3mRw6VfXrSklO1XAm
kY+kMiF+lyMqk3DMgJmzh5fhvGopjjWO0mK9VYkeRrrNl1nsht9AA/EL4ItydKfJ
uchH7Rijbyw4EVagslV8obx55q8gs0hsrvOoKj6TtUB13a8O7QYFauDu2ALS/DBs
Jj5eCfoLxEsgT6/ILNNu48bR3rWebHc3xxhfVGXw2DIFbzQ5yUkN+hQ/HAY0Nc1s
SvsUqgOKS14Jl08SSlCtYqUjnc30A5OvAKkMY8rT/n2LYck/O95znNu1YWNPqnNX
5V5FUspOP1fTkEkLH/+jna3GuaM7/NT6EI1nH6TfAlfZrlp4D7YUV1ML8Hhpp3f1
p7dORKjfI2L4rEUg+w7R+UR8Cmp/auMdJ8aiktqJwhbH4eoQlKHpYnfrBjIlf/Jc
Ia4XR12sgusdBwK0wm1qxgQFmCvWR+RAl5Y0m8NWS837YMlAbI4EQVQ2FGGcBZKX
RyuXCbsAfFRPYdHtNQedKRcEeTikn1kUy623T3zpHlaBeeEq71iv8TOTSDNzZqlE
aeMWni8z05ldQGVEzh4hP2SloeRBA2HQfngqvp7BxS5IcvJNM9qjo0GoRuBrywf1
D3CdgDx5V+AfrROUElYSxL54T02PBAkrZsO0L+SFpUKLzQ0DnbMEityK3vmI+wrg
5Ws+1biWRcak3qu85VheR5VlQS2Njj0I8NUOIOLjrz5VjBl25TsQgXCSUlQ6VOQH
pAnh6TLgBCmzamp5aK6+9BJjfW4SNHzgYGbHK38R7GjWIxQktsaWmlPjOSZUnUHb
RyTxBV9fDG7soOmqE1HRULN/oCGhE9n0MNgIdbj9Xo3qJ63wKOU3agP/atX9ASzl
WorRLzIP6e28xAt1jd8LIFhWb5YkE8i1GiWwfyh1ccINL7W6ungPP6zwZk+B2T2k
n3tV87nILqXA8lON4e1sBF5/OEUp9/r1PdfSUCHbaHcVHuNpvpy0vr1SNZw9xQB7
Yq6F6CY3DSgTnVyJsts2xplxOyHIT5IE5A096M8ycPCe/iZy3GZDy1CXa92RLsSa
bV6N7Hcc5e4tTStPkp5nYW9UQSkLmhh+aJgtP1LaAQANXPxZvsNJ3CJ7whQc8xeF
gNaJrRR71Q79eNEv5UMvNuJ2zWgloYybYvrC0SjS2/4b1lZgsxmp9hs2t9v+pw7k
cPfVn04UvkMnsj1eb79gdgs+jmN0S6ZWSMF653AkjEHzK5wFH8YrgoDOOwDSfp/a
x0zxqwx+4XseEtbzoWckqUDevLmYPXEQ2e05UVK7Kl7BITx92H2hDoOrBs2ZA0AZ
+53BUAjOoCkZYja+HNM1wwqc23qaHirwbzaWzeQRjHNfHjOt4EYI2AYtMv/GsEBK
JAdRHNO8vAAqaStrILa/3sckSh4aB8VAmBTg4MrisokTg8FXVrrin1CpGF4/ZqpO
lHKuZAQ8tFvd60Hm91gyyICtGwj04F+XxKJ/6g+M032LeFhFcDwfUnT4pAdWmI2C
blukx4UR6Py5CkbgTut/iSQHQvyKnqOpj5rbr/YVv/ELNWX6vALl9L21VMLPU+td
RdAqJFSCH7sj91Vxp13UsFOOQPEL5KTIhkaW+6p46cUTW7HdfgMZHl7mhkHPCjrn
b9BwQmodX3bEhOxMEj1OwLqEKKL+Gyd5iid+G9Ehu+29NWB9TgoWHkklY1xHeIeM
QVQcwNTadGRWSgOF1Bd62NfPdyg95YC3e/eVs8z5yFqQryuq0UgEVm/E0p9rxvxj
GDMwKuFJK+Yl+U4o4pqwgM987g/icRbVRjEb8GgKrWjCEy2XLSdAdB/Rk+ZXYtLZ
my1nAw03GsRRkP+3nNSIZwaFao+a0cqABA2kE1exwj6sPYotSmqUjV4U+m0EKkNj
kYQ/ctEB2vawcZtatKVVRDVyAwScQlaPxImsqnXJ2fsRmPDjegOJB0Xy187Dh3mS
HrI51pvaZrx+iZCMm/S0XzXD/Kv3FS0N0qkgglyhVv5tqKR9vWP0q4Eq/D9hB0HS
JjottBe8EAA91OIjmC9QfOate5s3rkmvfA458hN/fAXjyoiVHXBljK8MbdVCSOgu
31xR724KLWN1ebkC2Hz3mgAzYZ05EkcMoG/wDeobTubZMhU0/0QXdqVMo3sJPsEW
chCZUph39QQTK6cbFCGbTPFF5pbJXUic+jGoHBA/Cmnt16aF9LAm/4gf4t1M0VNS
94RRC3S4DkSjcn8Z4bLCPzVWT96RrURHpT6j9BqOZIdmk1PEEdtXS6xnkKHq1xEI
izsnz5UPDrQ2jnPWB6bRCZS4FgVoQE3QVkVsXlFCiNYIRaC7ZCY889KnYkDiO6Nh
16Vbbx+DvlwQAwTDwm/XKQVjKE9kv5i3sTr39XTx89FIfzKQV+xcqx1QTPw7hVqT
oI6LArcd/euz65EQMZBaxTOeDK4OShXfumBEMyc1fWWdAi0Lr6RpbgVitMT6M4kd
8LtwYxrh/Ju5A/jd9X4668XrmoBCTkUjkgnNw7GAUiDoU+wE9KfztSvcgY5VdYBa
ctGfdCGCRUT7s5Xx5SOG4yHYHj7mvntTkFB8pr7foFwZsmA+j+BoT+oyOjNGSO8g
0hVaXWL77eKFVMJTKxopfwyagNJNoj2Puq8wKto0EQt7kkQ9XMXLUYRSU+TD3gCu
Wo7y4FWgRBkh6vxVQOxZwEyQcSV5K24qXDjmg2xLOf368diksmzJaKTjg01z/ZII
DRG1+zSsOnSajC902UevxDxN4q2fqGLazSuY0XE4dy+hWipHzN87CWhHRBDDkbRR
NpinE/EZHnCIxXByQXlO6zyveY/PST8rJjBfwgKd+HYRymmeDu8ZD7wp5wbMSsFy
aa9yBLLVIPxcRvkcz+mjRsTcu6y2/HCUjw3FB3JHqW5KihinEZwsK75ZJjnmlvwR
tSp00xQdoVd5SuXa8hK+UUTWDLF0P2kd0vjRKlU2XR8J6MH8zsJ3joraEVf+PQQb
55pYuY7CjLEJ2ckywl16errixA3JCbIwCDi42/k9A07WnGD2ezLTQVbhJU6YWv0Q
V+JDZDUEyMY6Q9EMf7HpahEKNoc0MKr4TRegoo5Vi08BAmhUHOTT41yO6dkRhlCv
eEcCz1Il0IVDm7EKTfTii5x7MJdQLW7IktrjHJ7wcdOig6296At7hATcejSqTgLK
PpPymDYQcwG4Td23Dc1oIw3IMMxgUdjViZ1ISlWPMyGIt3irOSBOR9gMOzKoPsX0
UgSyJI/pT4o4EsaeO7nAuNdadcN5pkko1rse/CnoK8iXM5cNGQ/3Vtvf5b3+RDBA
yCtqsOrb2EOrzVy0ogsTyD+DLDVq4xthKu5EKZlnQ9xrPnS8KnHdnLUfTz287xAf
HV90p5+JPBsgT4OVUqrG9ygY7vpqRuFF25g/UhjkhPVBGeBojOKnHUH4ZnlLk/aK
uqN1PSNdj/PwmTbtmLZx/ZBHzpXTOu1CLDF/mYnqmN8t0TerNsZ3puYb202kU/dp
YZXcoQICW9kBS78wIUoL4EKQRyQDmr47ljMRtM091Onn0UyvAyeY7FoR6BtYrDr5
asV6deN1bKyVWBH0Hw1pAfbUJoyaWJ85BEdaNb8sB1653p2x+gG0BXScgFl2wJCq
sMBuqax3BM4XLYL9M0TjF/PrLCvMeLJWJZ91f0Al/KxxsGdj/3sFjbmiPcM+jn+H
D/gc/WAvwvQPumNIq56OQT/MAuE1ZP7p+0CMCEU/y+c4KrP6a8W3EXqSwfB/nfr4
bkytAs00pRxG33SKyykNLmiVGCOfXVMV6THT06cpolcviax3kAM1uDKRcWxdu2c9
wFg90iykpoolEmDje89AY6q05MZS+g355g3u81pekJGTSOHZY4mlAarw4Zjj2gIa
GUm6DsXY1Vg/pap15s3h5R08SQD6oz/B97NrBOyBmFawq/oPzIiOskpFukFzI7El
pRV5QI/PDhWob6I8piMbuKpu+wFKd5UTLTWxYmMvjmHnUvlUnWRTN8zzEY++HBOl
v9TfGJKJmt0ADFvjQw9hjWr9wfLa8/BCMgM+SgGxswFZKRrIcv7LOqhngtTssSPL
ZyFLGjpio9hNPzetiY0PB+zeCJpPviAsBgJKKO3IVmTaK+XFY4ug9t2jp2ec5P0G
gfr7Rl2YKxvPbSrJUREFH0z7UxxieMOgnIW4c0B5KjxmHEce1zZrnmz6rnD0pyvI
T0yAhikaCsHiqtsUDN+0abt12aNeKeb1q9xg50ofCvWFr8awVBpL9plyLmwqRswD
YnVfOrfbixCDBBg3Ot4xVG/z8CqurR4LDBQ2H+d0R3DfiXsH7LlcuFwgXrdvL+9Q
bvAE5p08DcVQMSbGUEPqsKRAs+ps+TOEtRBbT98KduAqcg+Yvb0cFoOndgx3ysjZ
XwudSe5DV8fv+AX1aqYoOPkqDYp5TKqSvBf2PuA8Bqp5mzmJ9ZKTfh9VbApZRWzz
5bnKzJjQDnmrxK6+F0+nW1SipBHDQ8WWJ7UEECB/4xUnniDOXBaZKsviLI8YgfCq
L8fPNFt9xtaf73O7zT9YoZ9V0v+3p1B9OCUfKDG19wpJKJodc2BafOSNAI/IfbK8
MKacATEjUTgD8uiJnpNuOiX4n0bIAjPQI18d3g9pJD1QCjz8nfff4dSMpR7OIsiX
uGne74hLSLRXD9dhrx6CfR7C2JCK7JmDrZeQ3l2SJYB4Nm1BK+Fp4bsSZZ5U5tlI
CiA9JYs13nAanYUYDedloHLxWNyc+cwHW0hnPjFk79dZW+94eES62dtEyCB2uxxC
Ob5B2fQlbdYsn+HbDP8ZPosnYqkoo+1x5gUv/b+64z+8sEBl2SQSkNy8qCDwd7L4
AawlCw8Wr6Z5uriW/aQUQMC5w2Avp2KCNdMAOhAXG0Yui8A/yq1Z+q4HkmxXi4cQ
2CNZP3AtEm4+R6FwDndH7eT7SlJgO02a3qCD7hEddocLq8fTfNLdzqmS9MWBIIKo
CzoH8wDQalMbZD6of4lhAtLKUKFxMWHNd6lfN0te+VeBXjE5+h4f6XmGDr7xj7jI
14jMvsuFUgHyM9B0gA2pdkhtgFVJoHiAOEAoF4XOrDdvgTGkvE81aQUElU10SaW0
ec6TP4gqhUL7MNLs5vDzouXkMn9ntHHqEXckJNm0HkCg64hc3JEHKadIXqTxZUJj
sHRw0dEPGDC/5knK8uM6iHTMM64xcvLBB7RYOQg88+JcD6H+AZrkmZBynlJnUbc4
DQnpqH4kW3GqNhtibERZ2aizYcQcyHBQqGF08KBs6hsZZRrUQXXRpquHXhlvDXwu
4dc3QLBOovBXEfRRMj/SaXZsLGj0hDz3cQkd9rW40vLPaW2tBBJ04fBaVOTm118D
L8uZyNmSuu+fsIZhSOgoOWsk7auplnXRqn0pcynSfOQ1uiIp2jxqTDEse1tpYP5h
wAlzAs+lEeTl1e7VMlYfiLF68GO48LyksMWYH701J3a2vySA2iiBkEJeezcxnwzT
6HlKsCx/DLJQE5cq8GwwQX25rKTOws9D17Vgek+XfpUmMMp03+JqMSUgsu9o4GDc
OFBWkaiGkDfgC7Tses8kmig3w7uzYCRkDsY3UdSRvqOGAPzqn0VuYebo+ohDgLgj
WRPTHuzM4Yffu/tqABaRRhPWF80CNess7TYwdzfvnu14yCBAhKqxce2JGecGLLIq
taP9qWLhsJlQycFqtkebSO1nwFsTzI23Bem/6s84yL/Xamq7jbPxMqMD5dTLZgGy
4tCKf/zAOBvWYmTY2zuUl8fyvda8XlPBme05GcLzHAhptCDFeIMDpzZZjjmefftn
lCsIh7IYmMFrGyo+j2qNB9J4QihzWvBscVKFYrSe+FO23Rh96uBGA8yVL5ppKKsX
t4mKq3W+kPad6EiX1t1GY/6BhL+a3Sids+kVLCbM1KACN2Dm+oxV74ymkMBJRaVO
5CKQeONHzot7NkwVWs3TibR+SWBwSv/CSM+ccqZ/+U2Qnzgltu22ZHJnLKVInd/O
E/q18vw4IVg7aAJ5mMj3IzWkXoeKJd/O3zmSHV4IPFLnV/O6tpivHbx+eFBZ7Yg2
pHq3M+8V/PKOga/33xbw7cvJlyWHMfUejU4q7GImzJb1O5oQ1040gaNn+4uvfqlE
BcXwIhoUgI1qN2KrrvT32Q5ABlSnFxZY7LTk+1Dx/fsa7VqZPzOyyN6aDu00MBhU
3tJi3h1DEfWMUwHHTHk0rPT09cocoHphdYQu8CxVp+i6B2riiX3gN0E7W0cSMtH9
CmpJgC5ath1LH3ywgdw7jUQQUVwujOwcJoiefakVjnz+LGS4XRm/AJSHSJwA3ISh
bZ91jiXnxkoWSdI1lrs4SxpITFW6O6wkKSN0lD+dSwvkML6nf2r5seE46JMCOx9y
I53YulDDA+DaUAW8w6maiSW/NjUFYIQM5X6GISyYdDql7qHLdvZ22ZXRZu9qeRQ2
tQo+QIPRNOB9qbgjk2hA4kwe/ijGP3z4jGTbJwy2/RNJ4/cQguJGKuwyURPj9rJN
HPNk6wzBirrvLes3aFggP62LeUIZD5zjNtZIwLunaeiFqn0Vrb9yBtCl9+mu9H2c
/vLU13rTE3B26aWMgE8VBcKFblk3r0q0qiZrz8ebOSjtFbuyCjrismRPQVA4ppKn
vUriDf2lvOlQJLhkE8+l9MYEVFGtL0k67zQJ/QcEkCBozduRIjI90lyOZg46H6ON
L+SxFuZ/jvP+G1GxbBbhff7FZgAJ9ZHDuA54qn6p/Bon1mIG3EeVLG9JT+qt4MgR
NOPxVv0a1/VOvELoXxUyMwGIg5nEFE4bXH6N0SKQFXlMAv/aortSPX8Xlqp/ObYI
F3R2v67QGW/GkZTSBQ8HiZ/kdqw3GsfY/891e91XcPK8oCrh479tKfKGdd9MHVK1
oBmYQtW+L1oYF9dD8GHHTRXYiDsH9bhZrEU0IwFObyx7NdMyvvrPZiDoWLvd9Bu/
83pN6wGdKhaamR4egjZPsex3JKR5Jtg+HNkETGmi9yH0XiLBqqgtLGdv2feVMNBZ
rpOfWrTENp+EE7kANZ9yA3biDIjVdZpcykC2ubqZq+WRaevpt7W/BvaqnVchzY9R
6EmBQHIc+TlGmHOu6vN6tw/CmVtbW5qfa+GYkkYiPXe6hQlLYgs9pwv5JQUXCRSq
xxVEC+I5slFwy0413vw1xrQwoNpHlHCvnfK95iJ9QBBvEuqwRkORoqYSGBUT3A/q
24WdkD+BkrzXUy4L+J2nWr6kiefDTHqH569wYC3+mJ2Vy7zsMx63bZeyFOVYEgig
hF2Om5HPs7fGlJf+NwEj06KSRwePD7QioyqsLP/B1896MlXyaVdeZgMsM4HWewqS
xBu3eyDoARs0KOZd0fQznsVDHAikkGpxjXZGWWv8NjQbhUyxSxGJ+5N6MLFCgXQy
BLYrNznT13Jc8XGAzHkubYj0ksB69kuYSIVWnoDlCWDCAD/pdPT2WthDJEbyjFNk
+1Qi9jBvRkigQJYwn1byyRKkFtiZjEcXC4sqig7HPWPsMEHXvCnQxrUoahsrO8Sb
0ae5Pst0w0Zp0/EE9EibQskHlFa351vjQov6giemZxqV/+kOyvLVgHbzAoOHnE/B
/7hEf7v2jIIEmb1rtpnAFW+lrrKcCIHS5+TvaqB1cQocQ1sB4WtiYRLGBiMk++h5
dgVnsZOeqRavSH8kdlPZaHtNl05Hsb/E0ocOXVWmFTac63pUG8VwH5MNHXOPlfuI
xr9pahTj1tUvSstp13vZqIDU2tT0uhTmoW9nwzgJ1W1cqSU0Zq5H2cHTFWJTCq2m
Qvoj6BIun+ee/WxL3Z8k/UUqXHrzZhs6GKW3MueOi21VBmetKfsoKSh+VsSEOnDk
gBgp+PN+SqLzxv0zG+kkxsOq8wtc4sgGGDyrBxSy6h4GWmT8s3Ab8+nIIbmiwq+q
v6UUK9fglED6UzdFoBu+Q/4IXxQ8saivnxjoOca0/5X5+rwlBhe+u4S2okDF6J+S
zdUXmG1S6oBHa1EJ/Pe1F8IuqyGqK2j/wsF5dQd7YggPqeR8dhWUvwsNNdMPQCeC
n3F4RYZGm+CBhEu8Wdkan3jkbdicniqHEZqBSKeaBKKeNeHLJA/18/B5uRO10ZQ+
CMcFZvrIbSI//kNyxsEUyoZBZgT7lNKsKWXwVdCDfhQZLRwRtP1MeE6zzcm/Fzpy
l6ma+XeIZWNOg9640j/pHhenF7Kzn7nheahCD6N75VHdMhvXrBREebuiW89nZ6cH
IrTZF6nFerKRZyfY/FNIK4QGxFDDYkzaS5mKXcE/RKiYy76tJqJKCoK809WkiPXO
j8FlTYpPvmNiUJMJ96pSd2QcBsQ/uabHH44uoLJ44fj/h1OLoYbnfMBiCIXdH+Bm
YX8BM8GfRiHGVrQGdYfHaYW0ZwkOj88TrHsTCyqSEQnDzdBiPIWbd6R0OouxwvZJ
2kqhzpA6C2TCRTOoy9Rg24pU++U2wu32i8cB8fiKWiF/bGDR0UBuzkpkLFSWLABt
iEV+fxtndnFveeG/NYM5TrCKIWS+jDOpzObVUpjCnqpUJO18MgAI4DmZI1NYxIlZ
xedmSOyeRBHxXciRVDlcJrbshcx7IJOippr6b1Wf+cFi4sr0uTh57ywggBVlFclS
nRvps7VUSuw55hNXOq7ThzAG1ekMJsRiATQOdrd7YORF9U5zf3tPYk8Iy4mIGL5X
8mEs+M6PLo6D6/H27LNKyg3WPOrtmAYmPPKTJvfDPZgx7h5Qmw8kVsT0xBhZia1+
tamw1iNMNqfUf53QsdOsHYByXEyri8hP1bufdAB4Af9M6N2phLYcrIEZs0zNg1eM
ogKBb4PdWJhcr47D/gGT8idW20s6Bm2jK+LWmYdTHz0VotjnQpiD/0Q95wKutww0
uycPMwRmdEV6rhyZhvr+Z5WEphM/JSH3XFFRMdxoVPHn5H6lfB/5Geons4A+sTtC
UC219HDmrbw1YvbWBg6JDR9ZifC2CgsizCoPaaZ4dMcDBWbecP5M7y0oRE8wUG5m
mlUgDiKVfBb5lQj9D3VKTUVRaLvUBTcBYcTXNdb5YXmn0Sd/y3o9BiVQBgfg4/qp
RwZUXvPH2Z6jNL3034YKySruR++crzD5psTCaru/L7h9qsENKYpF90P1XInPodxZ
GdXcnc+a1D06M4J2qYPvxjfDllqAVUvsZffyUKFBrhka5x6xAGcU9tmMPkzdl3L5
kdciIGl76V8SHPCCW2Qsjaf6rWcrog4PsD/584b59cjmfqv13ebibJUMOMUYdJ0I
eSWSk1UlRKHUmV/XhZZ0K7/CNUdTx9E8CzwoKSGxCX4xw7ho96wQZ12afvqnMnju
itkEdKzIJEfEcXWbT0wQYKHYvJqabH9fEAkF9A0d9x1ZAD9pneeUmVhM2SDvy2p3
BpP7JGyx1JGpvNmR7PwDhDizrWFfefs7Yy5aR2ekcWtpMUs6D4WugDxAJB4jmjyT
/oJ7AHGlFXe4pzxj7BODQooxnBiz1xNfSNN6QcLq/XYoykA5fCTTfM7rYTQFHv0y
nl8VLIcOh9DR9V1nO4g2ZR9fdy9rMGM2Rzz8f5n1ua7w/0Yrh2MtMyLy7q9tH9/y
BL8xGh1HII27ETtXdCXbJvW8bM5iwFChZqnEIKGw2bd2HsI3WEg3Ilde/O2Eh/kI
RF4atzhduk7sy9P1zH7QapbUO/3d9sPevpe/Ui2+gl9JL2PMaskQTm5oXHNYx62n
iz9OpEOTeJHuM4loqzY2oHH1ASdrq14aHWUSaHh4TJyznfnlklETbaFnn2S8Ogl5
X3pkk6AibRnLNnuvARo6tkh3astCODD1vaCp6k0qzfWfB3CHe68OzyMId8T9rB5K
yx7iypnMtwyPFfUv8b2NbjAcCzkn3O5NmWJ2fVYGPJ8KVRdE49ZpDRPMYPhtnHnH
Bk42RK4XxqN7OHdVrihD1bzK9rD31qp9U8WzcWl3E01GkOAtU8GBOEi2byQOzLmq
w9++/lq+l0sgli8yi5YZEUskW2PPsQV9kZD3iZ71M41YH+SQGGNBs1cI1XW9ltW4
dwmBIUhFE7zrzjOrJtZw82n6maueLNRvxDlIQ+JEQ4BQSCdywpmASUqEQa3YhNon
DSvyu+B4Sg3NpDjtzqvB165R0PAJihtc5XR5CFw3qUVwPuRryUQlz3y1kXJHzncM
Vm9uMcYmUMCJx5TKPdgzUTUzJ6mU06YuomOrNk9KsArt60j/orNoOB6h3IlO9Dpv
V8UlDbvcv7ZGaMQiCPKsKdcMAx+F3kziFTRk/yejRf5hwhAIyGaz9NbkGTzGi6h8
rezSBOi33U7WrVk5dOu5jK1o7dp9V2C2rpLrJuG7oPS9BbFJG9LvVLPUAAVIvxap
r8Ec0Nz2hffI4Rm9f2kIoXNGkwg99jCQSTa8cK1bO/my4nPnQwilK1UiENEfnmL1
jLT065f2IRbfRcRoInrw9FZVqSltFyAYgSR4ZwKMhvz/rGlmQ3hAvm8BiPclDrUR
6aDFYgBF8Vo/Uvs1qrl4TXvzgom2az5oubk1HvdRuJPZuXW6hm+VGK6fZtvZprzP
5v3fVjITBLDnwkQlWpKiLnq1mhh3fe9Csy+nuqZLillXcsXch+3G5cJhNBRFSVOe
i6IQ3luntoN7ScvL8bHl3WFQWLs99zhJ0PygButwf/hpl8+QIC6tAoxXiW3rmnFQ
Q1Ne/P7su9CFaSF0/nkvuqqOURYa5c1+q4N9G8RZlST9Lvb4mhCEaY2FJCYRUc5Q
ho1D/bpXQAeNgI1SlXjXWsUDTus1BPetgrmUrM8OfWW7k/4OO6T3iQO9yiHFeUzW
zJX9RBrWTSmafWosZliEPLRZRYsnPHTQoDWrDycUKY04//+DZh8/KbL72Dq93GuU
fo5M1FegOLI8NvVW7xgWiDYgMJbfyDWIHsaZr11v2AxgANdTJcqBnzfboxtNMoS5
z8x73lmJE/FmY/HY/CMP5zi5IOm//+H+LZnVGv2KN3zPeCpISTVbUGK2GLzz2QBc
0G5q1lTGoCNrB6BUqsWLM0n9LiHh1cqoTFgooHW1we/E7cOGmf1gEk2AVTkXagK0
5Kizjcu4rPxGFgpDXP79htWo9nBWjhpkARQHbCPkFwJJk958LH03pamHwEaffR3t
dPy1sbOlIHvyYBkR8TfK0T8lNXtmDdOEzf8/JT7PgEnD44aubvcP0CRIzx0D+Qmc
qF3HUqtahvlZCdo49rqmgbyFzjgLi9ZRUS3b/KtpwWmBpecV+jCwNU82QVv5RBMd
Yjlj1//Ljf9Bej/Ysm973hD39XJ9aQHS319i057zon/SKm1+y29SU1bBKbax2BZb
MCY6xtxcjhXyALwlGo9bfUGk2K2MSRs1SQDOx5BSpKupo9Noku5yMXT1b/PnPhZ0
y8JLj5v6qO2mJnTzzV8fyIY/we6jFjCoaPxpTbhxq7R7V58uR3XMMhWWDlJaOjZG
qPDDROT964srYKj9ZFVjUTD3/9qean3oObLKIlns8QkkeplHBKLzlopLQdDydstf
aJP3z4WRASjOdNEpAGXQ+ML4MMwbjI24/WU7mf3GoPdvfzFN8xWB4DvOlHXFct95
jLJWsHW837GKzBDrgm0h37SlTkwv639JyK0EGUPDX+oCwfZHCkmaboINMxRu4jw+
EqtuhmJA4HGii81BRTUqzVA+0bHOL6gIxvSXOI3Quu/Pasc4Dzk0GCuqDcdCXZ/f
44u0jgb7zytYahWi3P0pazVXmbeZtnmMJJxlSN1dbhomeJhjqyZZAw4IZeEcDnK1
eLktbEBQaWY/JToSnnBQdyUpwGkarY22TD8bZ2mSmsVu1METjMf0yqvLBtk9PO7X
50b42V/n5xxVMgPzh3eiQqm1vjSxF205qu3Z20qBxzWeBKbLdy8U+83aTmm1tchA
5Kgx1n/GIVh5v1we02FRjIDP1B/esnPsMQebpBxiN0ldF6qmuPOm2ax3gLt/fnBG
o3VeBX3oR43vyiTBTepwqgIfEXxgQPzNexNNowgdd8T0A0FfsOF+jQMS8n3MRBVw
4xRXXC8KT6Ih1hOHh0gpFoNmwpqmkYpw4EooUhhg4fDdyPiM4Gw2lXzu4UrvZVK9
qsVplv8XYLlwg96a9JWnb9aXeQRtPDtMTQj8mrWGOg8c80XjnbascP8QxB6+ICQ1
CQiJ/8cUpFlWo2yKMqyA9v1h3bzOU8cLGLnKiZA77iO4XVk6UeFC2f/RZzamlbL+
xYXjF3yingu9tzMUTbP45CBWC0/9IK+pRUfKQ1foj1fPJWz8JqnvUOBkO0pYgMbM
wvYvzwLVvqfmYcJMPiHK+vcKSmy+iW7Z2S1Aocb3UYScpU0Tkt/q5RHYwH7V5Zj/
vQcoVKbZksxfPMmta0PuuPoFMpKUL2aWAeVHRGe4TxgpwuoprSggeA+fSlDGv8SZ
H4guepdxIwfJtprk0ANYco3ybYDRlP/sf2mh5I9kz1dzfMKBKAUlVqx+7pnieTgA
J1XRLtkVAJ+LkHEpkoTxlKUBq2ptVWEQSFJJY+B1r28/4k+/tU7Z4MtxDR3lmyH7
FMWQbqbS70TNG9bC7Spgs55c4mNwtKQ77648DLXUZ330uKjD5v3Kdc1n/TQqif8/
yHXKjbbV029MFhZW0dQCE2vvXmb8jIKYW4FqOj8XJpFk9KFBroBCpEKONndS9Uuj
6LBvQNcWIIlSYXSs2t/zlw9v3BVZajWppw1P9KuS0ce4clQ2n1ixRUJh9Mg4QESm
BWN4cOpDIX/yQrA04WtbfSiQ/BYpxisc/P3iXoA4iP7LFzL0hFiZkjsl8V2Ncd7v
iXpf3wvHXoAK6c9+dV2c/f2oU23lhTSDy1yjy95BxAzfGZgAilh5Lqkk2Al115mY
iNQKU0x50Cq1Rt7KLli4qpDbVsB3VX+3sjDWzCzBwjQsiAfUjVDC641M16+bp+U7
Y9rgU3MS5OUvlupgqVzbzfE/cbI8/2eo8O8r7wLyPaVzyRf0RpAxIkpuBdxyN6xI
JtzPBOPhRw+VoX0rAYCFaVv757TECuotRq4pGePuNcsaZDXGdDbR03T4XwVmZht+
SB8+XqAvVe0FGnvo1yUV0JVlS+PFcFuxXP4Gs3NV9ZqsiDtBGbi2SYh/Nrph9eXk
IIDo8PZ0o4skcNQg0ou7NaiIoawDwetqXkWk/d6tHufzrhJ6+CDhtfFGZ15bpT4o
dJiMt/OQi2v5WraJCG0OAXdDv4fCpTGjT6AxUY26/QeJFEX+WRbpot0dDbca505p
JrnwiqFndhfXvckKBu3oY1aUacwBNvPSGcCeBTCeV0nRRyrFoPdCnSimDPQb3XNk
X/6j/NsT0FvF8/eZOSc8WI7Q7uN3/rahdWZFj/W1gogGf4YMEbTYOtQ9HmQvfDWs
T4J9A/UPqmnyDsf/0W0l1WpaItb3TdQBZ1perVhYvxR6Zi+/R5Nqndsjti4foJmk
lG+H3l9vx7q/vJMulPp3NemOFKwiVjAVAZNGHxbqNxwTDH9U9MOp/6gv6E5HCfcj
OxCdRYfzdSDmQDJ2nj0v2BjSHzHLrGhO06QTsseF5rVhQAAOHg9C7m/ed97rsaOi
B5MkgR6dnQqSDbAWHdc+6h8gNkj+CUhGnYD9z5j4M+iAvKHaS9apF5eeCTyCZnOG
yBYRQUCKp2a2UrME9fnUgqhB30XM8ffw9P6rXc96YsxBww/NeLzorZn4RggpEsD3
iD7q3p9F7dAk6zYXW5ov1JhHzmJloQB/44LRs+winbzmmn4lnnl4fmIxrXxaqy3e
j1j6ZtcdkoPrjMU/3/pZ0SOlxeIf/CyyKbNJmkXE9fN+03nRHQJrGYN3tSLPe9cB
bpzR5cQXrQvH0QTju1X4mAZclh05SA0Bf9J/sx6tjtT7P5oSz/+eB8KHEdfWd9D6
x+5nZoqkocQAxvnf6R4rE8hQge/wSuzpTD4khGM6N+m3yhfY5GzQes9FStK1sPeo
RMZa5/T80hFzhNJ21WY8W9Vvk1gHJZw/gq6HyZkRUFiIeCKYWB+LA6W+5ZNzduTI
lAafODwlNGyu1h0gKT9advc4773ci/PTp10JEE3RURApWvUeSt4eRl8JV7O/C6gY
xNeCL3uEKyLLClRbjJFrgTyb7Za0wPpjMwoQfEtJe8awcqH1vcLkejdlMj+38YL2
0KE0ZygdrilIMBlvaZyBdroTMZgELU8DMahlzhXv/yX3AjHW/0dZesEOxnP9HPA8
GG0HOofoBnFoDapSytSL6e3jkEjbROfGTTtw0aDI24Ev7yrcumB3TVw5HatiYZkQ
rjf9x085bq99435OruJ7wKvtYppQisdlk0suysTbHODDimhPLExCE0eIiQon8CtP
pOTTDhmckASEDqKuYU7AQXckAoKYsS3seI1/tJU/trAsYPdpUvzcwfwt4PGq1r2Z
ZTM24qm/0iwrwI9Zcv0xdfdAd0jZ9o5JbKd5hS98Hh62/0N6NG9yJ3Xz5FvT4rxE
JWva+vsbskU14X6rxRp5U5SD4pqDE++ExDGnTKoAcIWfnsF3/8wzLmIPrh1zNyX2
JhZyA+sd9MNPDsFxMbE6R+ubTMx9H8B1BB7Amv7ahQ+HQKjmkpWU2/TRikhvFkcj
dELSrWvsLaWeogFY28GkOlVIV7Vb/pd4tU89se78sa5RgVUJ1SA1qeSKNM+s2D/1
sCJ2OLp9Yf4khOA9yE+Ix7JkzH0FQuXFklNsBpL72o1CFjfaE5ugssGyl3jExm1o
7faDUSvtM0amINakbpnVgiLKmLPC7ID40wPIkPxZPQbFIyyysBO5gbvsxaFZiDV1
jzWGdQzct3oQmDUCFw5Ig2U+Oncr759kWnpLXpkfOiVbyXKexcqCfMEMvA9aQ0i/
4TZ9dfC0BQDSlGLqpREmR1frN5RomB0DHtAv06K8btUXGq606Gr4ZjlbAgNZfHg/
G499tN1uWz5MTDOdLfCSrcWF7Z891CWKy75/a325Q2dCXUgOusTdP9CVRuvxUdlC
I1bSKRz8fzkxrxXC1c2CMkYMelAgWfF+OtvwNLuEg+ZrtRcdAesRc52+CEJOALbS
JUc54MRMXvrJgMdW/15L+/E4/w3wXENGm2uO22oQEG7EZpBITd7HhOvvlnp+CKWv
IE8bzxe21DmkM4gOfZxRKpHQ2M4gOsHM67Sx5WgnfGQcZhFUa5gxevqgUWQKswGs
4AeO7mGdvdo7Pactx4XrHn/IuJo6dQ73yqKomeKOkjn1by5A8o2q58yYM8h5XYLe
TLNWMM6XbGzGv03GY/cVW5aTejkC1yN3MThD9xP//Jc7Ldd2EY3EzfgIDVWcawZq
pGlZEDPSrB49ZkiPc3NkLk88dk1+nwxRWZxHMaFJyNiWpNu1Y/csp/srtRoY4yhH
Go9TYNYXhWVUqdXR4yEQM0GVcIFC/5EpP8g5ZPX4n1fIliuCmrirtV6dy4DwJfte
kSjMqE4+L4fEOZNac1wdcN6zzCke74Mpr32J7POwtEAnOQfdUuIxSriZIRYhe6h2
+PWxpcAk1BL2d9EZ8bkjrbH88+8/A3M/90fqnteeaQ6eZZd2DrgWUrZVpyxtXgay
1KhfvOgJ4HRM6017F72zFvmgIcUagv74HABi0+NMk0bzefjm9ub8Z3Pzmc+n1cyq
rgx6yCClVixAmBtYegH6dI+hJEUq1zxoc22PnHi+8I6xT61jqctfwkkHLjfWitVM
lSNPLSogPR3LOxxiLTL6FVKKf626YjQmPBZLb66pzPGDTrGARP6VNxjhtBnL3BN0
Ij1shYoR0TkEiOiivBJ5xGkCKKVuGf0447FjgIHPIfl3EX4wJ9EYMfm9vk1bJqaJ
PObln+BEPO5ED3gO0O3JQCu8PG3nXbSLNbXVrT+QqVDVgCkOSaaV5xK4pzsH1HSc
Xx/i6vsKInsYCSyvYMOUFcjrs/TwRAr1TEch8VUQP1w/gJSxZDxK0eGepihO30t/
MnnZOT8bk06EIK8l97phdafOzynIQO9eZAWsQTSaZW/vyKmr30IlVqNQMorXdvRq
cV7qR66Vf2dBPSgUf3qg3N8SgsOOAUUqPEtYEmHwst9vfvMU7q8yx6gJB62SMmZH
KOnTqmf6B0KyYs+9Qns/fki03YHJukOPfSAmFZiytw3j8tkivuXKf6nbXFm2Ln64
EE7TvW+VR1ErWWyUBL8W1+4LnFv2mdaRVt3xBr9ia/V+aSw/6GVn+iNzgfmSHfvY
a6jJvF4rXsQdUnTc1/+ZxSU7yqmx0Un3VQKA2j4a1Q14QNY+0AI4no5pA8cUBDo6
R47uF/oHQ/EBU+pegQnyDgR/DHkpUCMXBsQ24lwZKHQIo5UZT0CcoOgqgUZoX5zz
ZiwO87Vdby5w+XESEW0FWA/ORRuAPWxczfEar5s6hlb57HhyTFya20vP+tfVEUMT
/2hQ5EDEWK9bLq7xiHV6x8CVxaEewQOcS/nH9FwOxs96BIh5H1PoN3RbBhJaAafv
Dw61AMV8GcjWkEKHSXao9QdgXIV6Kp222BVmnEFK3M8oU3evhZsyRlAj/NfHb0Zo
qSTWqoFVuOq6O6whm6wDFlae5irlb7FzTFuKRtXUUhbGsRNbIreufKIvDxolOVjd
mDOy1zSFVk+oBNiI6ohi7dpfLluJQrJuIMVscDInTrNGhhov4Fob8pybdoqxxKsw
l/Wb6Na+bfDJEauXu0s6qbN0brR+vHpVemANK94iXR+iZk4R3zxjSXBgl9X6zC6X
CGhjioWcdK1wgpWurZdJshweO5hC5TKyH3OqJRa8nG73rUthyi5D9WXY8+jccUgj
44mO9B8HYcNPwh9annjunep+vRDt7maTxt51w6IeiEciplV7KCiox14iPyagergb
7BasOelzrV5QTRWEpzeJ76PPkoo7RyBvwUqMnQGj6XA0fmuKpuZsA9649mwhBGrT
Vh6v98BfbnrNgO6rPIqGJ4Iz8+wqEH698SLL8SLa4dZL96RN4Ca14CwH1yR50V72
hhu7RwJx7zt7DFlPPlSbrIJD3HUOTZOwBzgz1s9MW4BUU2cXGELCzjNK4il8NxcA
OD8T4AgziunrH1Dk53OTQHTizWlAOt9kvOuw6J2CnK+TPy8wbr4PLbr37xxx2igI
EOGzOtmPUEndOxEB+8jo4yekYgtL98RP3lM1PUF+5vBAe8YsR1m5DsjLl4N6F8s5
aTlPWiXKh0ZHJ9ylBFIHi714/W2cYpHkm928tcSADU6DPdipsl7RJptTXDWqt12K
eqjy3GmHYZ6GTeeLhojAdyx32413gvdQUU/9ZSutGLW+fCEgJBW+zdW3ad7WvON8
5Om7lnA9VA34/IF0MHZY7khFddsexWh2JNuaYMh0JrV32K1KPaH/8MwX9K2zmwmt
Nl1YUbJu1b4Rgc8WMtaY2A8R6jrLochTlWFayvEK1ohH1Bb4drXoWEszpNLp1ED+
ggFSXPAOdpbhDT8uU8wBaQGhEDY3R8kXKABtmVFfrGcgSoVc+NGuZP3TgbO5bFwu
pcbBrupah8P7XADJVcWX5BsRc98AAg1s489JGXditAqZCZ1UNj1Dq7gyF4a33XSC
nFOZTeK/wYYP/nmVpKzQEteowO1+lUxl7Ez+LGDc8M8aVOJy/RRiMFQJQNO3J3FO
p0SVyH0Gh8bojF/iEUla+Pi+pA30T+T/FF+Q+MCiusc88Rrja1mIYCJ1xO18OBFM
m52wfnNMTa9iXJfH/XFVBz9krUJt1SjV0E6sfyAVvdzuWl790uVq41zQVGr6l7TN
HhedAvuTrHRaP/u+u69WePNLkn05XbZw+w+KLs+c1b/hMxYepgYHME+hlEkLDdI3
Dw+/qLQc7zX5un1GmMTAsJKI7KImoez8OFqlJNuqiwRL5JquzQ3hxBmCQceGruY1
XlwSfBvjD1Aa/oQi6jPfEboGdzW/fpUT1Y9pKx6kN07f3NSHocQsQNAhfqHrR0/3
C6KKJMvYCOBFpP53/P3oVasHHSiZ0fdepQOsQfZ4Pqp/SIalARQ447KJDeDZkefW
/GphZZu4gIBAW2sFHxIO8a++BNSDyhRuHYy69z/wY8GPsllSb0MuMQMhnNDx+6Ux
hi9IH5zekkF0ywrfb0Uuz4pZ+bUjT6r+6yfhSBxDc7UV50V2/m2LCiA96mFRyPwA
FMafCbanOenXeXNZp7q4fSrYH2FRzfLPeKcTRYoQOcFaTHWnmYG43ZkQnjGmn9Si
3RcAo8mvM3NQkjAeR6Zbtgz7xVHRWe4F+x6JjSnZevfB6ueF+d2q866w6PcMkpl2
Nh9Dy879lllQvEdpM3M1HDxBqjSYFWvZu/z0hq2az6w8nA77bJi8aYkTwy+yB94i
R6y/rCa35w8FSHM4TtrODQ0Tm6g+Mal5m3aXe/ghe9YURJ3ItePo6jO8AKlnNEQD
E2w1yYGgneRGA9fPc5p2mPAx8/t8aL3O8yeiNxF1YdK+BpF1+Yg3u631eLYZ+wZ1
qCOtcPwI4zmuOzPsGWMowRg5fbf3hUQayEykUIXG55XpUb9qKjloLQtRsKE6ksDC
XvL0JJcI2FlEawHLLHSZqeqztXB/MXe/eNeS7GqNbWudJ7F8FsCthk2kBqsb9O9U
yqY7B6JjPopuQ9MV7U6sDUD82DI7lBu7e/luAyYejh0Gq3SU5JZm5vvBh9ldNfYp
DFbqq73YvklqUgIFIWdXVw2Lsx8G8h3TxT+k+jTAw6PFD3r0dwVkjYAVeWxyknMw
VcvXAgEgxSeVbc2ylMp0NfD+YThQqcajUw2JRav3TSinl8mMQU2pwpkXgbFeQz2g
itJ6xQTpSrtxoOUnFofssL8cGezf5vy5VjN5Ba3HnAz5bvxjotuZaTteL6azeW6X
0r7Gaw7YTjNRrIiMj6h6nZMLLaS/s4UA9e1z4yDUO4LTHBNdk62EAwMsudN8Pl9y
NwiNMTlLzPwLOYGwFAR4W0ppOfxJPx7SpKTkCNwkKR94gln6zS+yTkooRSlcfztE
Mtk0HA99bcqEocZeo8cVGUHnji0DA15yBp4OlhNK+8Uh85mVgR12cNo30Br3AIO0
hO+Ro0++grMFkI64frbvTKDHhWw6nHySG6MAkZS36PYwcTdkEbZPcYq3QZt6He92
IkMtAg45qV2FGfVGvBB14Z3etlp5bchM/FttUjYEBVpAVutB5U9ge+xetGLN/ApB
bCJNhfm2VFVOBZnKA71lEag9QjFp63cKV1sItHrrozWfTdBc2TvNRUfbN3ZxulkW
nGAzz3Of/MlyVUp2hNPVKQswuLNXPEAqVKwvNG7rtE9ittwKuBYlAyAycK60PGjJ
onOimAw5XL2DkEWl6t37TWDwaNOHYYWvlmVSnl1Qb0rA8nwS9N1sj2WF+9aRFrGd
bH2TRf+oRhuxmOObk+xUmLZebbnn6PLnxToSdhqbuQ1+1eyxgM9MhCQ78J6YVSC+
I5RjWLyv9u0fQGVNT/PJw61AIU9JzcMfbf57IKg/gvwsrppZ9qqxKIxSKrDCPTTV
skGXwGq8ojGRpQmqnyIcTfFkIGYe0zizRHjd3wjNrGnVSvy2JyRaru/9b8oMdb+4
Ltalq3znOkscrT47UZPYizO5cRyytzEnxiB4IiWul1Po6QPWugjxLFku92WWO/bZ
47Sumc6pPwdf/Zq0EpOaYx43ip0+l3ZqPq2k3csOekfrGja/3czpS6VMbjZkQ3di
DX8HtnvFYq3uiL3DXwzQ2qHvZvhurT1kAeCOjFXxKcSpm8Ub/hnmxk+/wLwt+hHA
o2gd5mFkpM1e9i2x3FXasw+IJsLEgCDiHjZ4D9VZUt86G8f1pcRC5cdDtsTbm5wr
mU5oxAjdDlR8/+fOWaWfVV7C4+J2tyb4covxG0fWfooxr3a5jYoOSLpYsahmkXf+
MhPM/VWKEbAQZ+NefSym5fzWvvzaFZcst5yoghXURM2GFA1qiZNm0wG7YmvAFa7A
tDB1R91h89TFRPVQwyDurg4aZPtoVau0TPPOfDw+9OKM9g5XswfwIQT9UApP3oQY
UsB2HqDeiz1g69vBOOGjg38+gIOtbn11EllYSO+HZ3td3hM60s00AqIlGjewOQvV
gT2eWGJVkoQ4oGCcwdOSYmupHu3OlqHa1RdqLaxinWGL23YdJkscMpBpwUcqAwku
J6414eFLDkx7XSJqcH6ezpUGtw9s+Ky/+hUI7vY37MyOzuae3/MfLAKRo4uD9Mke
wtUifwFDthiosERnDIj84aLJjuMjpPMj5JDnBQTL8X00fliq0PMAt2mExA4nEVH5
fad/+2lPBXkYGJPWlwkUu3lBE+l8UhiDwd7+te5Hageveu4n8TPflJ8qPBLgCLPX
dPftZzcsRP4EsLPon4bVDt1797UZzLQhZfQfWR4fq1FW+OSYjQB+YYSortf4lAu2
ZrxP1PyasIKdFYamyNQenbqg7vquqADX06wcPColxizbOv+Eu81Mjaeq23tMcDoJ
igNsuOraAeDyZvp0+oYUhMUiXQKq8ZkH4jup5jaBSsLiKyjIrID8WTmd3JvVrKSl
zcj9ZbOuwq+xRkZAQ5DLfLPdTRdSdE/3ubuCw96YGw/5rb3MpBLYApNtVx2sjlk0
Qzy/Flxtv14HRxsmtHMhrFZY1KnvhU9l+KJDuAUKxfkO6rORqj0g68srUgQeYb5G
fc1qVjUhwfWK9vWoroNF9hKLonozBULsNSQ/wcoo9ApBZJjgRVrMSQXhEDY9Bz+P
6UMIsaPLUO029FtVe6jiq3PJMy64b9peWruRT+XQsSeCj3F4OtV8BRCb3Iw4VGqq
HD5nnht8topjYk6ZhXbGI6Bmq2HrOnYQyg40/p7w7npGqaELKjz2ZoQadICGj+HE
8J+/HM9EOIxOtlfO9PZdO32iOhs92Mu2xx2KtsTEgc2DnxwZcZ/xzP7KYOHvE0ji
ud8r6J68ElDMuHK3+CSEWnyGmJAHKA0juHuiOE99ELfpE1pJKJXn3wDQ6NG+IFnt
Y2iqcWJRhRXJxMDztdcCWPhmjr6IG9IOhlxv9ltU+saysBlKxTK8d4T59UhoYHAo
CkLUxwdO4/nVlsFGwdB4L4QX534fS+9IVtKS83ja9KG6tNf5M6UxZUU5fw08uUfu
goyTmdPaYvJAO+SslsG0Bogqzmrxn6G1H4vGY1Y82XoxkdIEppyfIxRrIZ/yoBS0
JQQzDxtv2pOZSpVe3z1R9tK8hnLasKZJLqh+PQ2d/s4frnMJcO2pfmb49u7JqGry
ezUSe7qROpw8rktmGr3YqF8WAEcTNZWCiqXdI6+FqQR+zwdK23pSiMkEYv4XaabG
FAbP1jnnndDpPPWOi44BzvMH0S+c7+Cl73OKw037GWi+jv0eBPk6o6QSFBKPyilj
TJtwSv/Su1uUKTp0uvtfYAdQsQgd3MYEhtXQLWM1LdE9BHC455+f/Cm97Pud2Mmk
+OOSKRFOC1mKKsPHoascnv7XFGawhcI4dDykM59QHF7NAbppl//L51D0Dt+vL7xI
oBs7BkkPAfRYE34cw5Jl1YOBJG1nlhjgPIjcwsxclxsk8qVyz+4Q1UPp8dqYwjqq
x8mC7bQ/iQmcTV/ZwqG/CI2sec8XPAnoLzbq8d5tcTUj6F6wYsw2PSUpTT2HIsId
J9SWxCOV6R0q098hXPPRnR2mmW3udfN/WUDfGJIFHkBVdsZOP/SdtqziLvAITjVg
w83A7rwcqCgEzkYLmje5WGZrU1tojqmtOTXv/iPAIhhg6kLky7auZnyhsNKI5wRN
JUVflpTb/BRkAMNYq4RRncvPnbysd/5ET7SGfvLaF4vp+grgkzvLPka3wenMeQQH
0UvF9XqiL7ZOzMpC4PuYaUCR0xlbeeifJtrj903qoavLLubPY71tARP0J7ZHy9nN
+5uLybw4rcaMLPxcjOXmoULR3ZCDT9Gh41h/dG/qhG5gzh7tKBsMxYJqLThsap44
nSy3YpxsGl5KPRTfgrBa6Hew9gzg1XSXp5REE9oBdnLhaeHIgng3n9wcm3tYizOq
SBAPSzie/8NlgH3RCrqWPDnApMEBjirivoBvCdvPkEKphHRqS9aBD8nu/OII8R0T
g4RQSJ1xowkiukow3o+4VM/+gLOMEn+3zHGjNCjIOa/jSw8Bumv50ZsjKRpNJg4/
zxf7dM8KO5e4tsSBXTwFD0bIAdLDYpbR/vFbkrUMRv9YgO94HVXpecEpssNzoWaX
t5RjLZ9lOABjFTUdQyF9TydKkNmETpDGk1WlrECkSbqOyDDtTudK0rJ5oeEn/+Fk
ZK95NrzAatxnOj8EGyCkdYPkJ/t/598Wv7WkN46aKimyg/hJ2XSeGBUagYgjYEOk
TNh+b3EELhRz7E2tiIDFL/ZYG2eliSxvVugSpqIcqwuc8ugHYZ5GOejz8icoILLG
+5qNW1jylRWGGutRTAjtvNq+Obx5OZwOnJubTlchKtA06RQBHvZS6fDHso9xvM3A
lptr35QE9eIpDJDm92wlmcJR7gO/sJR3Z1kJIqppCSVJySarjHsb0vgtkaZAu0EG
TgXDmE1X7TRfm0v5o9fJ25uC8JZ8/mg9+7EqQjDPXl6lp0X82nqhTCtzxyukOTeQ
UGr7sThQZymvzTs3t3xrK80jq6sGCNY+TTOyQmsLtkfCBm9bMLMjVoV5qaPT84D6
lDuiHsMnMPoj11I9tvr/tYvtJz6RTLrY+9VhSPKH0xG+EQ/K89hOoTjKI3UnfUuG
4wqxkmCECnoKyItvStK5fZ2vvAWkEkYeiz5zT9HMFidegG2UPaItl4ODcMA3Fwfo
rgx/p9NdPK9pvyFtwks7wZfMu/A1aAap/RyOQi4TUP1uzeVRWaj394ObjrE2NSl6
xXFYBuAx4JLfkRg/voGNH0uvYIW17Dav1IG9AydogQDRmKAiclXtDyDZG63L0cVw
E+w/2eKn3uwC0DfIjeSUQ+DFH1OniXSQziMqmakj06PWHKDMGIREw5ikG7lrcTSq
i1PV5olJGrALVrhrWzcxAiPvZrehwjPSsnchlppwsnr3jGIuI58VN9+bo0grzlSo
9BIPB5l6a7g9XXuKgxJxaLo1CLmHiztg/AyFLZ9IbWlGabaADpKXTCcL02pHLXAw
U2PpMVIdx6U70k/Z+ucMKDd1ulebGzXIbHNOJoC9j2ydITmvcvFCbp9zpFpSxKEy
gthfjqmbqL1l6gakXlRV7tfi/TrVpziLfrHfX25U8hwEh8kcWtXgMw17Wb2roKCj
o93MWrF/2gTplXl1mByKjVh2T7PZR2VUS4HFH1WReIpY7OyhcEt9hgvB/MOnbXM0
oi22mtMD3Z3Inppb0iAqzmRsInK2N44NTrvmJMa53gTD6irk6pGVNREbuqyVLEez
GrFK4oa9Kl0NfAzH7yPkfzwAJbzq1EnfnXQQXHLxkk2INuHBmbaz7oQnI/gUzQbd
Bz2yf6p9g/fCtRewlN+qt0Y+yGO7rIu7OumXTC1W3Rle0ipg83gzsrqYt5h5Lii0
1hZFMWdNXlkDtY/kLRuCEiQsXvNpxneqIwiEnArEQI/Yev7GDf2NaGKkw6vUiAGO
KZigM3HXaZLclm4Rouoh7LzkPU3+718HTPtoxvbXj4oILjmuxCXE47hSpymGXqmV
OJMy870gnrALid8tnuA8fVayWpl3CUG2xeqKnt5hHRiv69XIiSe4ue8HZ0klEm1+
HtvvJQDmz6JSufDErwTBawZP2QKj8IwzHx2kHtESzZYNUzcCBolUdAkkXRGWiib7
56zT7wYUEiupMK72FTmriEKO8IcpajIE4pJUHjZpvaqH1iS9BD43sPr4RJ0lh7yz
NuVqnwPEdBaAVwPXePR/vxCs53AcCv/Fbq4tX7ZexIyC1aZNS3EYJw/1N8lYaE7J
iMuioQKc5z9gRJ5KsPfeRMP8iRCGo3emAt+kQ+sSFgwR/L0uY7xmMjMENSoWhIOf
xMtuE9q4qmEWnrX+I/x/8tukEi6ntOBjcEzbQP2q30qZrdliuIoYFIA/xotf3F/6
/ot75dTMWJSvR+74fb1GGMKppOwsjElnEW5mv25tWN/sJ1DoMqVdivUEP+HbXxgG
XWxB25/iSWD36uyRdQ6FOzicxwTqEdx/Fdt968ymBr2Peb3Z378Gs611Jzr14Mo2
hZc5LUjSOtBmY41qg61u+DDuudNKAqRRw+xPUW0w/Q2LLOm6AkeEQ8Vzety4m3R9
h5e5XuqNclgA4rKDEXHJEUC90tmZ4YdWQ66uxueiIWeTaZdUrGP0L+aYmskkRp16
1hN44vwDLjF4Bim7pFoWp0bf9lz/ix34wcYquWkjd8f16KClNDh7EpOlAUGhgxL7
BRXuPViuK237aBjvJJ/Fk1iCv84DkTkugSU7n1aKNCMHa1izYOb2D3YtP5HeeEqG
rcuwl+j76MenrPnV+Wgsdd4Obq34Y/g0Hpth+/Acu/jRtVm34+AnXrYi4uMLfoOo
3nxAHaWJooHDUaWzivC37/0zmWlQLe4LuNZ153kBvIDjHckTYPhnd6D4I8nzsCka
Bo4TTLkSLmdhosyPcu+gOy3orfdPWswDiAQRcqvgDpo/xtVGvgEmWwCI6YJYGCaJ
LvknNgkWIXJopst8wf2FbWQxYumxnQGPqBrmhWhfIBLFlE9WO5VDxQhMQkpP3JWr
4iGjmR98vHFLxRWvIYohBWNF2GaS4OJAA9UR5ejdx79MozgsHIbfMlKRfOr4jk6d
LDG+FB+3C2MYBUDUtQWExum3Lh9PvT2kE+U5iungqwDIS416SIo+Sfj2bBb7dld6
JRqjvLgN2F+S+EEtd/mV5KP4aPEx5S7zJJLE7OBMCuTMQlc5iNOvnC7hpiNLeerZ
cn2uUc19uxykCISYCy+xFhhhucaVIzmQK6hmL0V26PBU2IDLQ5odERXuSDM5GagV
W59ayBZWHLIOp/qkj5g+7vUJ6XtjRDgWZrjNCQc2C0Xp4eYR6lZSDNkpUG1jjtrI
tGUAyC0bHi3q37fEvAhrmOqqMoXauXH9UzgiRtFB3AcqTH6iAHlgfTR8f1A841S3
lpxyL2Z36eFpdsTd9QqNZH9pIsoQeRjfmFCUXgqW6m2B/EH5BYy1a1iA4JFnh7HT
ImFA2jv2cKsHhaZ8b0qBRCg6X03jPLMNMtbRdZOsSUS9bzUkYeoWa2m0j4A/8yNN
Cb8HmS+5x4kxKdfFo6tQ3jme7Z0pd32jWgUbhpUTa91paX4uN7UPVp3K5jUqOEwY
0pCgAKVZGTOphc0hIwa6ajaWUmTwwffbBj7A94DpD5tRWk+S9ZVYVjVT72+MnIO4
VrQEPzHiEoiSgawQiNaF/iajkK0s5+9B6a41nzM6P9ZvNE+gpt3Tq2fLPa+P4Lmw
pId+7NVj6Jp563xL/+qY8WTQZT1Wgh6oRPh/xS6v7+8061jW8m4TZUe2KOc4vWeh
RwSdC9tqwB6V20mDmI/8FAg293ONs1nAw+Q+DW7SP5HxzYv1CfK2vUi/PVDQKYRu
Kc2538Nsshzfs68LM9Z9hgT/OILPp0M7XwbscXtnQnpKUG5x6Kv1bnKfwcvwzF9t
0m0J8u3qHNZSSiaWuEz3sIGSS0pE3qmNpu0SVvn4LKmSP4HZ7+UTISnTKR/rjrXU
GMLVpaaPHZtCPzmc2HkjiuDHBgtpLRoFrHTiLG7eCtTmYpqLj5dOAsdF5q7OyMdw
qT0QxiGlvTlN0znXrSlD4SAbtlIVgImYQ9v82iNcGo20MTzhclEP++W7++/t7+NS
mVWPN779diMLzrkaTU3eNYvKN626lXcKZv9up1vFjwhtJOkb4MH13lpwxamTm+eq
jwBaMI8pkA983RUxK1updLdFAyjg/oMYCpiSoGjj6KgSCOTwDIpdruMlmUiAWQVx
cO42BDLIhANtfplSNdkwvXoav40R6XTqsefWKhu5QJqAXPhY29kkzsvGvBUlJd66
xnu47ub62p6UhWG+9zarc/N89oU3sfL7kMa6w1KwG7x1h5OI5KPliFBE90VPvk6z
yPnklqi+sopIKTddWFKjtoxtZPro9yBiYNCQTzSwjSbWrqgZB4hrlKLJ6CQRKFDS
9PXcQTYEAuFHhJiTJ8r8IBE2bq2XzAyFhOMQgtsFxZlmldZhFg+7APTavRedZ8lv
X/48rvVXjpppgyGG9YL/tpbYdqgK7mV8uPNtMDYufCdH+kccuhdM0i4Q2LzQ5/TU
vCeV+bRhFurXsX8a1n0xK8/dme/wuM2k5x5PIx4CO/RfGc9Phsy1izbQe++Xv/GR
pOgGE6bo0Z/sed7UiYou7cYQftELVqvBpGRMvQMxi92StuPb0zS6/Z3rU6sr2cty
QbH2JyDcYtkHer/CTesEj51JI+MlCZaehsBvxcoObOBoWNJ5G6madkXhiHEsTXUL
IUlrkKBO7rtsbxgiHyyk5BWHIpnpYi24uK1izR7aLiaezTw54ZYbVx6ZjzPkl4Wj
oEVAbGY27ZiVWdSst6V+q2Iiru2l4VgA5kSH4hZeOya88LXxC+HMTRb3+T2NRXoL
Cd0n2i0x7C+VPJItEd3IqvPNSBEBHcgkLcimLF9t5pDorVBEMOFZtz/SPW1KM3sw
+B3Yru87z3CEYOlc47aDlEoH32gS+Zg/A7rwqVKrtKBbKO3Z0nrE1XBOvaW2gmB1
gfj31Z/QUHGRLsiDiqjXCVtyXbvc1wFijtQRathaX7uDSe3KClxd3f/1SIyKckb5
rt8kQB8efOx4JvAVWjR//sWMNicS4gsTY9lSjPFesnFpMTMVJ4q/Yyw7HUP8uNuD
zN++c4Hm9hpXVpw8f4Yk7N0fHi9y75YVIx9Mf0vgy6FMXGh2TmARKqXqZKtyp2QH
cIaka2i4P0kd4HN3PyEWxcN23WFh9oWEg5PWKzucjrqDMkSC8Gc8dR/gaUD73PIV
qNO0l5HWSKYMbbxR3ZXYPIT2JCop5TtSq+YKnDXbRP1l525lfeijTiDH7T0CZqYt
vT9Vizd89IeHmTk7ZfdAy3AE2nG/VBgIACZnQ2tamwiNgxUORC580QAT5L141931
991MDjKX5X7Jcdeb7lUXHG7J43VU2vpf29B8vVMOvb8/b6vYKYGwa+g7JzawcJDn
597XSAtWysqxJTR5YFo1VA7YowPWB+IyxxdIWwEbDAnYx6QaoGKY11ALpQioFjm5
0NNuni7SkQEOAUT4H3ke22jTjzL1ykKR/0Il+hnUXqEC1bfzHf95O3phFRh2hPkC
IFN9OtsUeU57EaVt9B5niCYaE8mtNkmKGQ8wiQVDU2iYS6ohqv0/+WpJ2riUqX8Q
ByiTSUvcCTurIXzodngqrBOzsasvkZ9IezZH4hZI+wgxPfQifU7hHwT5QHzqOroH
REwLUnr4ttwUFFXzUs7PMJsScl4/QQ55gWxFoo9eNMGAbFogKd1LWplS9NP6RCL6
J0LSQZWopBXkwvdCWeZokk3s33k1xyH52g7WAqFo5Wr+6Cjw8FpMIHlTRM0smT9V
ffqwW/vvj75FsLByu5F9IKt9mteFBsxzWOBE9uftNzC28i+MIynWHZxO6xUNO9TI
2iNKg64+jLWgF05jzCq9iOUDyIPGeTN46LpiVAyV/1JAZP4AiyK7yBzlIOygb3LB
f9wAzPM5KMk99eRZCpvkmeyumBNHbV2hsUr287mRmHbjsASf4fAo5teVRkER8iFZ
/MoN9umfGgbMjJRGiHUvPd8M6RAyibj9pmO5pz+fvrrSqi0smw0HN3m7cPXZ7VNL
dSYsat7eHnMNa8EvuqeqIf8CWEAfJ2oIJ6c9Uh5fGI2CPL8jzZeD6vfraOn+ejtx
rUp7rWwh1GUYBt7mMVMb/nkjoGFZtwOWkUoM0m5h3bqPn+fiudLzlHzqpyTS4g0X
hr6GL9X/NyUgLuHQxiF27HbNG5P6PzA1SGJsnkJhiCoXbL8E+YXbkNd5BUMO+dIF
a1wrfDcTcF6aQc19hif5ea5kqR/9QDJVQZdpOmC2v593wOLxPn4EtYwjL1VsIpta
9lhhFOJGjfjJU1pfRZO2Tu3atb3wNVJNMbN9RUGPT0PE/pm04kcPorHvJOYy7qMT
JrrFalSWL/B0GWAi5YYUFmHVCAvuCwvQttwww4b0ZMny8DxTt4jVnmJUVUJVSSXH
cAlcsUW+/j+DwUVf/iZrf/DNiCtSOL/0kX4XqrZ0T05UL6B8/yAu4i3fPV/VKnjm
IKFnuiQenKhWCTc1Cid7aZ+xQxGLiVUeDVHOrRNTfyX6PwRshGZmQ+gjH79ND+N+
7hAwjEzivbT5kP2xbfIWOIRzLjb0RSxdyuAa4addmsgNjkSSUVsAYY+Fe6sUdeGh
Za5uNMUojEihWCRf5F9yU2F27C0w3Awgm9cD81m8D8CLtEBfWamvT8CxagNbBQk0
NtwTS9aNiMmNFQ5AN9OOuptpLDX30cSnqEmP+6Ei3kRCuE0XQOkbHJ+aysMsnx7D
KUl8h2w+htrn9K1uneMg1yne5ddelxrMKJSm06sTZo5uFIdR+JN6ZcWnxv0rYzbr
k+J0Z3GwA6U0VXVXoKUQlX6hhDkwOEvSt018T2zWCTEvlHd2WNqSyVMdKDXc5MGW
iSTvB/xSGryYEExOOjGeb5snutkuyTRI7lOUvhRqvj90AtS+pOTrfjZgMgOF8XuU
HwQhR66Bl8hpD84IPwLmZ8Wivb0IxpWoTx+N9D47FtljN6etU95lbictId6Egm07
nyppqsEZ/ax+3EH5TqaPICgZ8jxaGVocjEd9ABHbA+/Mh92H1VlsiEKsNTrczN3o
yj8silKqOHpisD6Rx8vI0HUK6bNLLGD5v29t6V4GBpJbp55T8dPgsESVIsf9p/7W
y+ASMZ55wKAb2+OhBuLmkJfvxD2xK72XeB5chUgClvAkP/UcGnocuQmwibkz75Ga
EZr0pl/EE4GghWiwMQt+tN/J3FP3Kt7DqOgVloygx1A197bcz1SlmMc4Pq6h+lTG
1KtkhLFPPFmKfkvKfn/n2VMVMfmY4QoX2W8vkweAiaQqR3ncIHLnGsCSd5inh44R
tblgLw8sqfkj7ilyx7rNfycxgnvfHYEe/tf8XnT9dLW3K0zTMKT6g/iDJ+PdMKXa
KZecJ+zIXXz87D7AHIFueqH5Z1AGjq1NK9QiluA+EKcMjy8exbY23g6BWxcsvhfI
zv5xXrdhRe8upilzZso2LQL1KFMD4j9jJbyUMUNMMWECnw2s72WPhCIBvuqYAdUV
CZZXguezLj60Sqno/wzCxhNzRMcP9yLQDRQ0HICTa6B8vRWlO6NveZOtZcWqkNwt
7eLwSg7cRiqZm/7ZEBln8rbJx1neXPy5WHW87f2L7zikigbiugWmdmtOMnIiHKxH
Vaozem1f5WZGt+b6COa+IIQ1uIQlNj7PDYnv22jQVoN8pHC6oyqCykKOerq4TrzY
UskYL08rPsEYz5kUMEE6zZYP4zpbXiSJSvRcwo4dEbUdVggAjfcM4FicjxJZdsD8
u/V98bqvcoaQpdvTy2IWnVbbO/yxPVlFBiql8S1Nw7T5mpBAdkRYz/rIBnhAwKoa
tq+JNPiSv35AnnHGHyvAu+gBC/uNLB49lCcYWsuw6m2LmbzIxjgkITHZssWUszoF
7mOq4lxgR96j3CBQH2/LK2JprVB+YOn9N8HBkec8IFPESJ4BO0d8Jb8fzmcibnyI
1OsTYLJwqzmjX9FWT6N4ZJeZ3qveWpEJOyr0exM6+bKbFHL0yoTt0tRQL407O5Kx
JgUzvuUb+7zqUtC6UJfwhkCCFZzprQ1pbJrXeT0JxzJDFr0umFKsowzYxBx09B1J
VRoNNEhp8R4T32hc9J+2hKl86z3LDqJMZG9LFXZnrO9Zp4zwixeB7DqdeAbQ75vh
YmvyCHkudAYIUbXJNtVyMFVgUdyC80qmfB8m0D9pnxeZTcSaJ9AjXYMFfa2wVtzU
aBR4ySvdL3XyJ69RZfv9THKLEBubWZEzL+sl6+XLGDzC8WSuOV8YbMjhDio5uw/R
3MyvwJNmGquyGDQ8GUlUKM8jHH8Ws7jIIgZPvpT4beS26Eb8TkutEUY7zfCmwhbj
9QIZB4odpyx78Km3qPtawBxBe1TCXIq9E57Qsxt4pyTFtZd6PtOQtwNydPiiTJ8I
K3rQfsHMtq7O0lmeroumdp/jZ4eYKv07GWrRCTSi/xKoNbSToPWThPW2CSNt+ox8
xQBs11qafq3YIR64q4K2JstLkynkXP7tz1CVI4oWK+dfvyKN1C0TlttmEHHevpSh
lMLOT6KhBeCTxz4Ffc7Ixme8omOqzyEj38T6UeGpuT5t2pghpfyR7U+Ch0SQRxue
Vchrb8z6p6sXX+uoMlq0wsKWHVawAPboyJ42tRdqRGshRNu/fm/O1CjSNetSNtHJ
Dm6KP//NLRnXMNdka/wvrbnnQ1B+yBmM7/dmXSNBxNvqZjGWmAvvQrLuDn2x+gFE
O2J1jZKW0yZwnIA3Moo+aEOpHnDXpbjyU43/kBiaNQHwXJ5HAND9xANe4fSrDAsa
zyipvuunfNqnxkNHI1gBg1GycAWl31Lwy+5CplQNVig=
`pragma protect end_protected
