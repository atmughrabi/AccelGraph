// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
I1/U7plIS/5eDtulWoNo7jUAp7aFKtTazIM+SVDek17oSEJ/P1Gd5X1TyXJoIpa7
ckOfUArqyiAD6GPvJ+Y2IGFrJP8f74N65G7pjQ1kTab4yVrwrnria3whO5Cxh5HE
PiDqPAHHo/zeaZ0sf1z/3a4jtaeeiKB5fXB+OsEHbNg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 193728)
0OncLNGkUWvqVx6RqVFjMbA/vFPJkrbQpq3J6fXryEUl5JPWiCddO8e467mB403e
HLT5szFxtGL3VIPx63WloFGLmzgoiXuwlYrUacdi9A40MMoN9ayvmf3DPYkDowAl
ehc+Akljq7rTssrAFHqh/Y0omEtf2B02J2myxgbZVt32usaNwKxeM3T/zZwMm/If
tmO1MAM4UfuRv4uNakoTjWeK5bSP0BtJhEDCUfGbu42EzNm3+o5JakoARgCG5LjU
r2bzkaptlw39afCIBMO0eHqHsZ9v3apjrtIl/cGMCfi59WKpDUplb/QI46XaeAWD
i61nNBP6+0jgzByeTT3ZoSM/VCw2IK4+FOhPMAiZUrXAvFSfOxiuGyxp6eMscrsW
mKpwmfZ+oxuugLzdWYSNRUVUWX9u3jXjSrQ05i5Mhfcls3QHQWje+gMGlRCxkikZ
zaw28iJWo5Xfsydh42Dp3KUuAuTdMXTGdlrjTSQepewZAF6a1Y9LzrshwSIMxqaV
waqKRJs26WobqEvbIiLPzU2tc0oS0xT8eThAqm20M9BYyBw0Sp7+pDiBop9pUmEk
Yi7djglDMof7EQZ0nSXI7Z/Yzq7szHYQ5oc6NmTETlAaBukVhXw+YMPmwh5qKPT7
eVFO+ZpEJK4g1OIrkfLla5wizkwzXCuKmliHnn5aRuikVToiEDRsupQtxejsIR4F
l5w4fvCY3unhZEByj1BcZ54w6itpHJ6FR54DOK02Bakm3G6yhSGHH5GPYYHe8Ec6
qQ0oaa3e21QA2XDbtW2FOw7KEiZHhBATgsH1454YaO7u5mh8EK8u6SFMNzuxdq2n
A7+JnZjydmSENM0rkuVhnVvO20Ilpmusv7WY9r8uSwM4o4Ga9aZXANuCIHbLVcqE
hPuz5Hz783IRJi3jTgXMB9Z7vfvZbTPCLgJrF69tEOUveAS8/pOc1zfKrSnA7i9T
8JlKg0CuJ+dIOKknW1m4pv3UsUF6AuXJMOVaMoBPzP5nrVjw7RIyc9pwMciq9CgT
GmTXZss3Ti6hczeAM+UlXP2PqTcIhVDB4vMo9KhG/RqPjcTz8DNzPVWqXyqKTJe9
As6xJY9sUfC+apxzZg+NZ7yDPb2AlSaJbDtoBmg3WzgHAZu3brHvMu75fK69/6LK
YtVVqvlYq9qcJCYjzAY6iHmrbFxa20NAj3n/ENuRfJN02vfqUY0tN70YRYiendht
h4eoFClmGNsPps7I6/dCLmCNpneZBV5JuIWq2Vji/akR8MjWdqVToKK01pgn53Wu
Nzfysyn7986LQ5cGcti+SQbV4UdSdp7WrVBzHF7A1Vo1HdJGwrd2fXpivjk07EBe
gTGoqV2iTz1l3wDDY8f3LDKeOTNkuBKjmHqYDqhjxet65aVuxf1dJmDx/ao9FHFH
UxIe5M+eRGuV/GcrG/sVkx9qvLvW9uPYviQ7mHAkmJetfmbgWVPOR7lRtnr6KupX
nkG2WJmRN2Z66AYtrHbLd79RH2JUUpVCGEmRX7k48joAKhlAg4/97sUiRg47hehv
GvtEEvuXPyYxfhGG/EpeoR0Q5r5JlbMLbiaBnEpK2Ia/xj73RqJyw2HyZQpa/8TJ
3UivF9vXN47Q5751rs+HZtCeDd7QO1gP+5PrJYRBY4HOBIcGhznmuoxCBH93/Qx2
RS2ZOxM76Te8aYCZ2Q3PRUkFnZpXIA9v13M22EfPtnGghSpYP4SxOx3j8Oiluzyv
RFCDbuhIxpo0nyoc185c28o0WZm1eXGgYGVHrYZdlxzKvl/Y6hK7j5dTlPv7noEA
9mVnjsDOdPxmlXa08rNUhShDhDJLI8UfMLS8tNukqypyy2p3y/RdKMXfRnwn8Ydq
n7bnI+3ajn/RUcNf8/t3dHdJN+B84oG+V0EKV58kGY9lJFILrwqz3utrylrZxVhd
qZxZ+EBQ7fLRbAdz0M2cKKB6v35GMPjyioDNwNFdzAVOY53g7Tq1Cn/yygnuNbfC
QQm7hOZpCzwiJtjO0cheTkdVIgsfljb6mi96IZGT2KWpdHvYj9F7u+eGYMdUv5ab
Cvjyol1hcLVy/RVj80/pzR5+mIyaG2ntsrqGVP6SNkpwJL7oqWKTKt/JaoY/edIV
71ovft4Wno7kdTg0rOcfF64bRMYiliJ9cF4Ssp3rkxPH9tSEiIdy1Opd51q6ohM9
kkuJYbcBBGikxknbL+esiQSVFNj8vBXrI8v3DA7JFjzCcY4s1tH27DGUDjVPR1xF
a6NIUqGnBpaP5utti1EdDqqGUUM0clFNGrWRznPoitkKAEd9jv0ZZuPKTxFyBUlY
ow93Nr/5kMX6IwRy/Z1G/uT//SvN6qskNbcYku/pP4BbPHES5mcnR1dR9XfKL3k8
qQ+9vHMrqZ7hHSO4W0hsl1P3uk1EB3UI3ZZxBu3ecjai3EKILXispspJYEUZ2Qla
bo6/ob6ExbZbVmnG4Z9+9QAJ1OR+61XZGTvgL4ZjsV7Ol+4vgfpSpavn3RDaI9tY
9/C3WENHQrlETrQGBbhXYxEWVNEkujlTqS1DJJOYb/e2W2/fvt5DoIpBZ8H6A0cW
/45PNWgmFwNAX3/OawJKPKRguP+15PlHkVUQDguJ8CkZpRy3XgWeRFSCX8ivK1Sc
NyEaVWIWUxco0CO+JMsvAr0CLLSCJLGj0hWwpcTc12uhEgdnmU+wocT/ByIguB+i
pCxZP1O49jbCi+pC70qkiQg2C7RVflvytF25InD48MAqoO3jmTSAHrjPfR5bF5qo
EkGYNcWeMrJz6AqUh18G3r3TDvpOaQl305jVUIGNwt/dOQCZPfEsHkL2dL41MwVy
mmy4F5CHkDQCvYRkqfcS1M0RD/AlE5TiNl0XSim6UfjTsk1CpgQChnkEn3hulHgJ
J4UPKnSRoVJrTwmVA+GdnaHbX2l23q+jBwdg9/O/Dz2rhTPHbeUfRDRuVyx/gViu
8Smf5z8d+ogsOR59gXwlYJfHAK1LqR4d0uloyFhh2/eeEvTlrNcquLzQZawP70SN
Oo9brqGgi4w4KcJuRb4gAIeADh4ZsUBqdZyUdGVEFsUyCZ8o9koNE02UIVHKuYr9
zuYKLpmGkJQsT24M50zty+hP3nyDUehNl6Pexx85AoESMmCBwnc2B3HPWKb9ZRs0
VlTNnTSnHrZRX371ueLmbuZg/XtI5iJAMMRfeLCiPwkFF2LpRnKHEPuootORBERv
kPufYQ5nvlcQK1L79PVnFVJxCXoOKeQfJmWVOXRtiq+1qXVuI+9XhM5S7rgeAVk1
RbncuUCZV8dcB0n7IX1waeNwm1H6Ab3GzlKKdVI2oBMOUvdVSAJIJlsW6H2R5dmR
hj9RLnXcQkePkAFJIAP1XtsxhR1pRpTM0x+C8e4qYpCN57ICil3ioztAtQiNFeKY
C2+eKnT0nxMh2tMiVEOXsOWfkhaeWSnRUB9FWODepoiUzgbTujZcdLXj5Ln7OK8U
RGb3x4qvJwGceZKT5b0KMpo5BQnPiu68J/l/gLWgzKov7Yo2O2saZznALwcc5B1+
NlIGtm47vFFPfnQGwrk4vfheA7ji9fsA1JXa3FgQwzpxJi4SGeKuwozeZwtOeqRO
q3J6AFyXxbf2a7+g/nPwnuFIERHHXXNNY6RbJACuaRbqt4WfWgEBEkpsOIiALN8u
YJw7+zlYq2g2T0p8dCCdE/7AKGVW42obg+NatjbrMw5PZY8APfGZrY7gYZCMcWbs
gS3Ll1R6Qk9oenmlEfO85D9/DbwHkITBOOluphGpU1bZj4LIVed4wtsRWavwQ6Ya
ZbAZV81OUWLA0vijj70E8xuA0Qbh6gTIFbes36AVh2g2Id/oGzPCLPOqSGQ2ZrKs
uqeVLGJxcU5OSea7XTgUOjxm1+d5W9mtutLAwHBa2E7IgzEfmFCtsMWsHcdfx8P7
C3DzSiVQ1M0xQHOe12op1/3tPG7UoSYHE9dhd9tnJ1ZWBs9PM/o+pMquS/5VkSs/
mCV7H6BQc9Lje0TBuwdRCMpyPnzwEY+92Grmo/NMNwmB04EBIjXFssMR8Wbx8QlR
zGH0AVb9ymyjnQ92u++S/MrTvFgopBGtsIB+DNPklNkYnR46c3w/xZ0tJmvWCmjx
tGOCgF+8l1KUP0T8JEBABbpb1Cvo0zqSZx0M+wq9bVtsItzaghbJSkDEexPGjMwO
KvDU38RjRAu878ofHOyDZCjo0ZwW06Y8QqdA/ZkX7fHnsIQDsp4bXoDVmjXuCUZZ
t6Wk1FnGuyDwk4AgpXDm4Mtvpv0DofTbzRTkQXj3MmijwqFmAnJHL0Bxgthf3HH2
iguyrVHmAhBb920yEE+o80dkGDO0s21Ig1rSqRJsnILxyToXsLlQK4WRP6+lOR19
xrhEq0mDwlWjF5iItT/HxVlfPWP9WmM09EKCrVxF+Xw3OeZtD0PzCKj+Br4CyxkV
6rv8RVD17hnjg1S2eQ1c4NtgPcBmbAUal/MvESFv2HRNof06tIJlLkCyjyh7WJo0
d3RzHQtNAtDX9Ap7rG7iOpjB/UY03xb6wow2IaJk3TPC908Dsy7sF8xb+CidRzD8
2a9pFlOq1wx2rF+wbIMjC+NlIKcIi6R0/WlE7m9TDHhsbn0u7WB7lQylJAocMsBo
2Ex8GPzviKXyGpQ9hVTcF1i9E9b5QXwzCr4hTVJPhyEZlq6vMCPi2eZPynzILsUO
Unr0HFyccZat7ZQuoLMWpBLGXXs0eqXRwofxUYE05FPpXe9WmlCiKn9P0hSf61lq
VlH3XCPPrmGUvvmLM27RxWCPCvlltMNuYwBNWtC6/Lq56+j6N8xaclC1FGLglr2z
J8hFQdxB1ZQigKKGHgnOMSFuUKfeelDe/7W0oNCjEm+A/clNYKlndRA+ZnqYqysd
svTHSWcXHCz970MssEPiK0DIlw1DqAWmzSwtuJNErZn0c1nCt+Ki5vgoPGVXnJwW
E3mr5rJKJ+/po9NZ7qSIGsvCNta/YtvOW+pJyKE2zxaAnaKH0mVOwFyfWnyDXNgS
SMeRn/rqfCB4Vs6HxxZQUglFX1TTy7G9xA2ZmFkoxU2tUDIcAwduBQfDnENuzGOP
SS2S/idIT3ZGIsNilG4i6hWG3IFmFubV2W9P9ePEZrraKIUXJWd25ZjRdubMUNO1
B3a82cKCJsCGHhdPFNvbA7f/NYSVrXNU/cURnW0wur7+ONtlO2ZvXfOaFcBNn4rU
3l5ODbQwjzJqDQ/c0k7NI4kQcyAtOFJ49eqx5TnbWPyEbsWcA9wp4utYTOVldLFE
Oi+WI0rr1z04C4QEqvJH2KQToJEPxXNtbNA420obC9xkw+c4eQfdAD/71nsnBXNy
SUf8Jk53ngYsAvao7ddGIc37AyGDKkmoC4/9LR9a88LdZxEwDychkDVJPsUjXvBn
rUdItbxxEd/tEE/O6YJUTlmcTg+hpluMLKvBhslkmbqM4cd5ueDHLwFpai1aVNMZ
g1f9sqFUGwUtZhcvxyWqAnv2c2nssuvUBFOkFw9JP9I6dNdL40mn4FueQ7gUSo5z
sljuCIeE4RZ3QdHOBA+hLj3cueGwz1KaYNzzBKA/kjiV7PYHSIGICJr+WUPdI+3O
NbzQBsJun+z8+w/994lrqAc5U21PjWbc5sQfdSIehBKV2S0Kb7zPQrGvuYIpCGYV
FLcidOhfbU9ouDIAmwoW1MSriK33uwyozJVqlpNaeNGIgjt05kIA0xG5Yk9/gHUA
ldqS4Ta8+w3p8ZMA4CAht6oD7IuypzZvz7ILwwZXZmKFjjGARjUKQXYwmEK60efx
+su/no6c2GdAJcR03nGovfp8NHMyMNq75E/fCo9/bNRo+YjuEPvroYQ6fSh0wIG/
QrCKmNAqpGdVezYbKVLy/rm0W2VfIK2FsLgnfjoG4gVQAnIxoO1koCKDabWfvPtF
nJxJ9nqBfBaiT/4iCw7RGlQzyEP+i4uA4fWhheKm/rDk088RqdJWcE3Bxo5BVr5T
gwZ26WWU2KC8C+7On05WJrS2YCtZW3skdU2Vdig9Jj+4LJYhWti0C/bj+aWG4qT8
NalYdoCzxzKfXpXNwTWHmwg4ye4pYm32IWRuI5CX6vm2OJj5x/o+HpAOolNE4Ugc
/JoeBWonptHn4JS5tLzfpmC52a7ySNL+ftEMyZTQLqvl2vcvWtyF8eUTs8iJxW5j
r2jCDUdrFDqJMU2hpkIxECZ9O2YGTSoZ2B/omIz9IfhlleBprwlXT56mcGb8Tf+g
Se1CWkTQLM6fmogM/IyT8ZGoxNMiUzUF4HoNLG/FEmWcxyygHynw0VZV1Ve6Yhrb
EtfuKYJX0bAE1XSc10k1Ks8nZ9U402QOmSgxmVAuh3LaNn1l6nc7qn0XSehLhhVQ
rLM/KGTMX4NJJsf7ttPD/qPwcPFeYYgR4e5sTliEGwT+ED+Mx6NPZAcoa2ZNCYoa
LUR32vHUYIUzpX0Ej/l7/5jnJYHzLXrscoRULC1PhJeTa1mnRaO6muheinrU+Z4T
ohrweMHU+WBVr8+KtHIqqO9A/+9sQ6U0m20v/9l3WsmyRh+4vCc2kFkc7/DukUVR
enNCTPmsRmg4C3weawovGJ+1MzhM8Ko4JcKePkwqPwZuaTq8/JZ3E2toR/vXvWzE
u3dTWA03X0kNNQoSB3yq/5w9MaG9hkYmeXvINlyfnHR7ZBGVW8Hzv2ABAWbVthha
XqcQuIJD0XpAHyY9hKestugLOIFjZGhXawNdS0xV8lsRrMjuQDSRC7NdAuGAIppK
7zzEaIsPfKM+nf3zZClAsEkgAkX3dWa/PTKtMVadDEh4pHtV3RPrvWGma/i41fOc
YO8AocCy4bXq1b5XZhp0iEw8s1vInaherc1qJK9a5B0i6Ioo9YxRcKajplDMYNL0
IqeMODaRB4FdNNvhkAr94G7QbZQMM0NwNukKk3RpmilqwhxgFF2d2WR4GWRN4RKP
DBME++Vxcgv+y6aefB72TzGCm8uN7AU0Q/vHDA6pz1yrl+9im4uQvixcWjUfYe8M
Wln2tu24kABAjsfq/zDwcPkBP6TCHdvDnsuAnwjTz3L7DxN+WAKlJqhm59ICOu8A
X/3Mktl8KskcjGE6WW0c2N/hGhg3mrmUq+LLPcvCfivSCJ072CQYRy3Z3hqbooD1
sy1Ptn/X7ICxqljOeMY9ICgnhFyFuAM7DN4h2H5yUvuAXwKAKiHXNqDz871ugThF
6nEPRRVYOEs28+tAK37gvNfvkonM9/BWc6FZnvyko6QZZujxXGUerLo8lh0YT86H
Lxx6oKz98yXDXTmvVQQmvM99CVkOqM59upbTp0lLRDtit4BNaUMP32ci7ntttJmC
K0hH6oUcN8Ju8AzhCsWwjRVZEyCTLbRnDswVPScdKIdiXwyBsedSgKzapHKJpqJl
jjazPeoh7a6+883pXisypo+f7OxLOefwAWNSLN7C/a42iTLSGzyBkxU2HZ/IAMSg
6g+AMfBmVKjB+83MG5mvQoaTDN1BXeK4BDqYN2nsbki56RQdeTVY9ZQQtfQDKeIs
/lpGeh0S3VieKftRsCTdwMk9eqP3iqfsUaznYPWtZwuf1qCbaTh6BFbN0sVwh4/w
8VtGDFLKuOCtD45EDcxTR77vsaMH9UoQNMzk2b3o69tLQHDnTnmufC7mUzEj/A6k
Y7GuIvE3i8fTYO6ssMAECJS4ie/TsnaFsjDF5u0eHyrExA30Grb7dpweWlnOyqgC
nirFl50QCzXB4tbJzXmKD74GXkeeqh3RpCcpaM8wG0j7n9Qfgx3zsubyw8Uc6xmn
I28Ik0O1ywnnfDZ+asV0we7LArZOYzg8mTHySt038hXbMK0rNwKwBa5DNqYPdhIB
YT3aXCJxLCs/TeASdbxTFtBf9ZsPdZX0U9XLHj1+ctxOJwe3KaDQdLdr82+7Rm1c
wB7GHGdA/ffcGuvKdr2hz8keSFz6eT4VF2uGoVIg+W4PiyxB/yY+q+2dl0JXNsMH
hP6xutRCXwtzoJ4GP7jxJq1ewg3c3lpmrpyyfdYX0jai9wdAZVRFEQjZpboKOOr9
RlhGB4b1ZGNHRujdNZUILeuTxMW42+fTJ+vZ4B3mF4eiUKmHy39pzY9yzcPFdIJV
+uMoVY75fn9NUiCAnl2ZVyJkqOz/2Xyon/IHhIJM7YV/7z+oqQJtGvpi74XketEg
k+hvQczgh0G8FUTl3YYKX44bEKJovc4UK4eddwmV+kTXbRIDpX2p8sCAyLVf59V3
DDChhsd2QO24LRUmKefJ/J9LD84GTM0ZMqP3H7PDFeRNPhkHbQSFlz7fwfAD5OMa
bcTQ4IvoTe3o8EYbm7AzLW2uwgzwdnz8XQE5hf6+yDXGeKB7BDXr32m86QPQBsth
ygjzi2Axa7aggerIhw2mjwwJ/CP9hDPSl9VC5ppAE6ZuyfHWO8Invlj4teexGe1Z
jr+nG2nKeiy1P8MqmC5fIv0qwhuRpMusOLSw2s0goLuuO58a8ITpCx4+/STHhRzc
/Rg30kmsbaxJ6IW4C4OjespFdvO+obJX3mQqPxkWX5RFBBD6LGYddb315xorP2YQ
SPFzGVaD7N5Hul7E9GyvmQ3n8yRfmtgLlVv87QzrkPR49NBhLPHS6E0w3lK2wLce
aK1pvjG+m+OlYLML3xWyh15KzXDZSz41x8aSKKeT1aybzsyrkx4c0RqlieIuIHQr
LRW4G8eSW2MhhtkBUR65XxpbQ0xI1bzkNDQLzWdcULt4AFUBrivRFNMTbgV57OGo
WsAUgeKSLpTvcMBsEJGevvhrrVaWmSfhJWb+7lUyakV0O4LE8B+rU33dZBwrOkS4
bBtb9/0gY7Y/AeE0t0lGeFAG+knHAqzkojRhrZmfQW6WULTDLKHY3v1I+q/77+mk
89bJs3e3Ihj1xbbVHNctJFkR3KfgdgXEAz9Il6aCj9epUSIxtqMGoVBaoYP1cqdx
/2Zr1i61du8UpbrbrsGy6H4o2BOSj1HfSKPridDmzSeitcxm/9cYZhF5Ae+vJkZb
1gofiTDETiMAUdcmm7aPcuxcPJJV+I9HrE/ZcMFHesvvHmXU0X+pdKFBHJQKUBYi
GETOsE589K/xtmceTrSYqpaFfnFqusfnWerlR+dUlA8U3G6Oog6VEuJk83/PYK09
8Fg1d0QHE0Ukv858uqiaL7JB+2+E1IgkMWOGtjGJtDCSuL8awpOlkR1q7dRUtd4l
wIOnPpolEDzpEwCpTL/YuEQx+QpEZyHbItWzEtFu2wt09ytgwWjc54NBgUjtp9lC
r8stIhM/jeSSB5AP8B004D4u+s9hadvgda3rzOG9NN6oUcbiLHNsrIMJB0OYoQQy
QCIlzGFdnCAd17ipVbMcbHWqxRMUMVy+yTYnZBt7G38VjGyXEbII7vhW/ATpeFYk
OzrnwyO7qZoBPWphPy+PCQkiPaWiYHB24GnwnaE/vOw9RXWMQ/t9/2I582FiKgNy
jbIAPAcfGAy2CuWyUUc5usSzgEyKk1gI8slBA40N8WO2lYYnER5yjHI7/tuYun/r
ifVNsa4fg452sVEYvMjvzU62ai7N+JpWZZr408r7P8JANtH0MDUscE3lXUW3J/e9
p1qUEUoVvjsnmw9rOKinArrwp19mq6hsPk+IQFc6HADA/Dm3SSK332QtG0eVOR5e
ZLfp4jZToNcdLRqXTe1Iv/RDjbjoULWNZPUN/o10pC3zFSu1MPmS268GLIMGeBv5
BghitUu3A/i2E3o50rBbhKH0lZ1Tuz9ODYhBDV11PbTIIFW8JZsrujAiLlGI/shi
QgjjEfCS4uoKz4Iknzahqy3LTtjui8zEEQ35CfqJkt23pZS5d2yo/G4MkY+ISVRD
EgLeL7IyogqPETOEMLNmJE5IZI2cd3hfvXO8pdHJ+gwCDREqRsEYDuW4lybwSMUA
Y+gBNAJYWL/+0K0ip8bWBjt9H984qiVGOm4tZWMZzn8ikGyss3MkI7EWWuw7MofY
6Mx4vddgWDN9Wpl8oKUjdM0O+hSW3VMdvD6RS3E8al+zqvZ6EsxKICJ45OYb17A/
DY0ILyNiYjsbqdOeg6b9B0on9NXMV/zJ4BfyMQhskTv1agfhlQ2GTRFMGAMLoCoa
DLOn5pdcKp4yuf3dejESa6MpaysFzDjmak6b7zOysVgZ1rFpNH5lHSZOnvc6nPBU
WcARH36JWMkgfjNL14DgUYs9HqASi614yfTwYo3xFOlUMC0MIWHFSGXA2P7GBQUW
BwhC6zpiiS/S3KmqgykYbs/6kYYhjPbM/Dx+YUqIFA3wSgM3QU8Q1nNB0ZBC84WN
IMyuBo3WCPFW53C3QXMMOKfAOdk0C01+6mAx6fdFL/HrR4FvboGxRtvkOy7OiTll
mRQlSD13/mU+ympPaYg0xRaGAq744NbbMAMcHGjq+3DL8nzoE8Pm27jVEAy7GObB
D+tXIvmJCg0iitcYXZpFqhftg2feUApJn3ZPQAe0FKrp68reRgmaiw/0UgkXGwq0
YCvXd+VZFlCW7ch7ZZaigJe/4IYwSVWYClG6YITQRwdALiBaXGaqi/FIQ24b5dCB
rl+Csq0LteTyxVCmlfzcgW6ckytAeBq+EtaQEaeKaJG/Zgo9yGX9YcTxU1HS1LI3
cyCk+J01frh3xGSeeswuFm/AC7eXxL6HmgxEoaZpmlDkKFwaosCRDYCyf2hKUdu7
wR6mm3XydOM5EBKnX8EMQkQ9eZg9v9FFzQqWlMhRlMMVkISmN2SsUmZYrq5cwhnb
hr8rThRXqK0n9HWGyr0VvLmVQGmjFW51MitcoK9G4bQrwor23RN9YXGro7+8dl+q
ZyhlGgfM3CiLTK09tWY9opQCnvZ/IRA4Dw9lAlsf/a0JUH6cxbj2RQLilbXMUuwp
jpzmYDeTuGEthAtsc8Xj56Otc1nP6ap5Z0LeNoAQNE6mKsOAzGhFWj06FEdL3g/+
+lFEoc3YzJQKLmpKQkXEkQtYXuxrFjcuXRA/AFQLXUsVGroNG0Mzq0t3aqnbvV+0
eL61a31EsuoDBKhvzGgsnvSz7q7Thze3SqjWklgyORCnATbAHtc+/lP1XzaLJOAe
nM4Vz1+zBOQQVz/eg3Cm3OL7fF4LCnqiF581w/fCt59m4Na5DpkE1iARKDa8Ln3Z
/UbnI9/dP2NUy0oPeYCKjO0cb1aNwkTqNg0QGAK6GVsW0XpEpl7p8Qbov1BEJdlt
fP7Vm6aLmWG+J5FFs0H8AtK8LucXcvXp0hXoq2dq4rCWp1az6i6LRNjLApFxHuxs
E9URvQRr50xI1gX8Dve+txGLpBYtxwwoRHRfzfnweIo2S8dDIkrpcIHIKP8Rwk8P
CdGTWgoITmv88E8GTYvQuS9X6H8U94NiEjGt1CfMPjVoFhV/eoyQ2cHtTwVddPXX
EV0LJwLx7GJ7nETiUsd3FAWos4Q1syzOw0lvS3cqV6wXVNBNFnfEsTkHRvx4C8ut
+mL8srOsrvEPPqrk1VczGOSwh6mqx7jA3vrWM764IC6e9YEngznlCR9U3mlJpQwb
XcvAu5IipVEXAZ0ufFBahg4MwvTpPo0tiS59CHYH8OE7Xg4MMo68N9G/7pLveKBK
39BKRW3+Y2sRqWaE/Yxg+PPEtG1Bftr1T/SAR5HrpCD7ouNejkPOAkGzhcMLvt/V
O9118LcOBspJY8M+FOkNEOq8+f/ZaUZcxKd01vB5clte8rNuwywx9PKiSHvnSc1H
Yt8BuF1ROGlpM+F1pBjJpTdaERb4d8Rm46u4JShS1BdcDLEgSmmDuwVNPHLavlxe
F3TF1KFn9nXpPc02LrimTiAJ0Dg4tjGUr4f/DcY+FGESqIQmQ+a04gmwXFYpNgI8
c2vWOVTaJi2ljl9tqhYL4YsweKYABmSTSbZYYlv787YEXWRvZgK5Xg1wSuy5RdwO
HUJ+e88o7laPX6ecarC2JjNFhMvoItKHKormNVlQzj7iuWHHk87xUub9DiUV1Of/
ADNLui6DK0fpYDg4jKuI50baETL2o2JT+KBfbdwGKKO8zqSb9qkNUz3c/sXncShk
xrNobRWn9i3WfVNX/sqL35pBIJlOT0Gqz6um8Lv/39SGQAn45zQNM08y6bN+Ajoy
myVWmoI3fqxO8EbRSD0pzDbEypfbQAaVvZwOx57hrrNHTBX6g6OFGB9wsmddwvCh
v8O/gZBJo7AS6wn+6IybotA7JnMjYLC+CHFgNUS7aAUgQOuq/75gsF2qoY2S2CQI
qOnIy/uY42PNID4xM2dZP1W63I4GxIxzO09ioQyh1uKMrPXO5yYdN3OvZc4giul2
vd7lbDVm2nrPJOrFD4htyuvjtdy+tknVPYmSdpWlZJKOmEZ01pMuZjvg/T1RZ9w4
XK9O4a/9uZRucW768bAiMXqwPTzla2ofO2Qf3m6xS20NrosPvEJU/FXUC0ZkE+8b
NN5R83PQUcnnxIqlTC06fytGQZYoLLd0dsarFjnysY0I5NLSfhZVNP0hu7ZfFGBk
IKs5A2Kx99t3DnDmH5dRngb4PfsSE3D+HEj7lQDVrouyNRterwhbBdSGgQjkCI1v
5o09AtESURyWM+vgPDYjEODk5e9fInV0Iq4WW0jW7Y+u5UPOYrlTPcO3EhnAnpTl
MEEf6sepici9ADOvCA3uVmbsmfUdJiow0bxcIXtGn36Tvs05SqgT5evjml2eq5QV
GCyqrTPaPfVhBq4mX1OuScszgif1A6aapjH0Ug68XVjk7SOrd3D85ohO5FvMNq1v
I7OXK22MQujEtYBmAekMJiRMu7utTqV9D1KelpWzK8CHIekebzDUIMaCyZ6EbnyS
XjZ/4x5LeeaX+I/8O5Z0v0fwFlciLpglmvtlTIXTDD6XosC41kbThrtxBlxg+Qum
EATqzNkBhRVXR/lY3SM1z7oBuedL5imqqJZmP2bB8hiRkqiPWjCiN1TqkpcvP4GP
a25GU4XdMDFtz3r+Iczzj/Vm6AFzIXFyu9I74pUk8zCzGB9QrBJSNOLoNcbAsyt/
ciOpN6SZJeUVrHfzOkHXQJODAYkHzhpJxsJS+Jcja8ynRwp8wUprde2MTWSry+Zo
eYfSK2a/7ToKS+bSpj9zX+s55NyJrPrXE0x3CuKGU/VVlRuAEegJjndNUrH86FRf
nmPNzqw+RPeFmI06g2Gmd7KzWg/r2+SbP0uROokr0eO1J3dSOb3Irjky1VrC+pFO
hA9jTAF5uk91WZnAnG7bMKfBQrsfmZQUjAqPrnwVpZnb2LI75ELnpp0ZimDVAGcz
PIwIiPvnUvj0ScTGqO+cogL+Q68x3IKnnM7TQyDYJAZ3KGkDOVmxP83/qJDNqa6F
qmaMeMaeWn6LWYFu+Nc0UYFv2wvtxEd3A5MXxlNNNqpW4DJRHwrpZdgeOptpKOT3
h004pxXtCQTG1Ekeug9W8V6zCrMNFgooXrZseDv8MzGBZRcMy7ZNy+2Wpi0wDT9o
ZlJkBF0Ctech/fctHfsGMBJ74e9TAlJKdAwiUfKMU9U2dbmiD4A31AKsEAOuU3Xf
gCLw3cgPon2Kg7wPdpE1jgGkYpU5J+QOUceNdN6eiN/+/pTBNBODTb2wTOI5tGyQ
U+7z2NXlKtj28sP+JLWKPLxxKK5rEnJJ5TrSLevL91DdTscjgfIojCWQoCaNmiMy
CV8/DkLQdacz8JskxnTrX8dvOk5T43aTXQAgPzlvAOiJvGk0o3PiQymjUseZLUUn
SCgwVoPEU+gmbKaLGlbTjdK7ICG68rBYceT93NUvV2QLmzRCkR3Iw4KYni+tZeYW
8v9c7YiZhQpm/1WOM5RTZqGV7HEUoWifgEgaXPP9OKDPbMqvIHng0iJqfHH70lPs
E+dTU2Vn6GYVVwqnwTyFAQM+JVDZHNfhHrsDXI1J152dxy+w8N33GiKu9gFBWA6+
Jbrc+nk5Wt0wZpgtcIfyh1JwgnQDCOt/d98wmBKF3FTozlWwf3OkxWZFOQB66J7m
jcuHzELvUm4+dAH7ZxlU3pQ6DeFcwdTJl8Pwc1fy2r1+RVfKWzvH+SA/n4HGPuJw
Bq42b52EmRJQzBQ4Nx3LgmX1x00/yaS/2jbeM3pb5o0buGoMtTq5S5O40ef4HfaL
//sC14IX2kFhWq11OmreR5wQhADIr8WzKLhPPrjjqxhI23U1lH9kSrB/v2wX6doR
LoiUlNp5rlDArTyPSiXx9KJCSisDAUzRy3PvUZnUJQF2e31dS+rrTkk1fkv5gvih
IxgoNm2KpZGbwvaRalurQ5QFwSA9PcN4VC2EPbOAhD7LRmPcZP7IkwRidUr7mBSU
IXKCejh/asb4fzdYvvbgpbP0o5V249SaXenPU4AlcBlMNhYroZ0UjWnCPjYzxdrb
rfanr2idDJvpn8KZylV0XJFTyr8gKF34Gr1N+RUWWZU4fLvyYKBzrYZa4uQONKsu
r4eTQhdbuMvVLh0Do2hw9jTv/YQy+tFH+tH8CfPYzrTzGxJQqxdaIgEQufAqiGA4
NzSWfgTplifnCksFvLqAb2dsDK5FciRab7yoyQUL3yERE7e3hFAJsPzrbYCWWO7Z
AciXM3Jl4aOkcCdslcPPj1dnoilBZf3fRZ5l8v19Ak3/fwM8tWfo1aJ5HBEU4aaJ
zi0l5Oapp8OXqnhhw26wGkm5QYiTK/3y1CGu0T/xsFMiECtCBNsWrvSOLdqyf84k
o6SEcGz0R2Atai3pVdozaG614kUIxXcwt8x5VVAGdiFi2OTrn+P8Par8T+3VyOQ2
NGrIH3+l6ZHn5mqhV3Y6yjkI1s9nkvea+r4wcW1AEaBKiEVetEU0JS7gSFLhGNio
DguNu1wMM9aT/cfzRf2gynKM7SJwmJ4+579nA6w3lxivC04PEzr0dQY6jAvBu+gf
K5lGehWWiV2VCl1Gq9DkItNvpbpCxUA3JUgXM6VY7ki/ynt6MNAW4VydNESdle/0
Lf5eSOHKxz1ghsFRbjz+ivYDeumD6r70qO5T1TIts/cy63cn7iD0F9agYNJpzvvw
j3DYgUElaqpZv/Hu1GPKOSQe/rlhT8JPKGy0z/vt3gK/lh+yknyjhSDri8NGva1e
303tLoIHdSCfpDF+4SPX7rzsWaGv6k/bvPyeqDO+Sykhh5hYQPDhc6BREDZjwRT8
kny7tobfZH4oXzV0ZJyzgDiwcv2S5gjUZW7LnSvw17PJmZdzG3gFrV+dl87/eRch
SMcKF2YjxPwE2gf8TY6J+/vbTmcXwjRiH4SwP3c3MOpGhRhZILVal87i1wDqfsww
jZDMXY+o0a1KDq7zM0ohXTftBqMLFa7NQHb2YwU06oxlfZDOT+SVfq8tvmGwCAQN
H4pH6w1NzlhKJabvck+dcrb3nRvhZLg7HcG306ZJVcuLLENDxKOwPvIr92AFZsiC
cWdgcBedDTBiTbWXwG9dZLq8ndeqvtf8vp6xmZm7fSPCR9u1f2MEbXAnp7qGw7Zg
eLHhi1SmIM5pVAfGLhGTD5qm5oR8lneE+A/r2atAQylMzQhwTLYvv0TqjWI4l8fy
SdQVFLs79Jjy7jM4tWDTi4VY57r9YEZio6FeKItr9LRm2aBPapJsebAjGORuzAu4
OT3bdrhqfOuvGyUodIAR8rr3Jo01Vc2U2r+VntRNWvSZoCR/ko++zuSk/ri1UMCg
16C3A9eV3/xQLo+8DROdrGgYuXx7w8TsXdNIuezHNdJqkEIMg0vIeJtPbfu8vlJL
wLSLT1qyxZQ1lvf2bunzuxgQ9RbHDjgbLHbRir2IilDLa+GEwlquZW+pNcjT5Sx7
CddQ5Xi9dcpY1fyP/YnXF+mxLwPz9QkYeqb//rUNvG4DiDjTPCl7u+xR8n+SiLIC
VCz0bQ8N2b13f7Ac/MD5e+3qq/l43qML9fYSuvahVBzegdS8tOXDRkZffkw3xKUx
zEtpF52WTAZnKztIy0qk+bO2wBYXQi2+n1qEKlIbysU15Wk3Xk8UmsBj7kC/SY9C
XFMlLGhmdNX6T+wVSWxyWYtP8XK5LElVUUaONp3KadEu5IoxOg2UVyN1HrsYzVeq
lTcvy9418vrkyrWLAlHVvhF+PHam7qNCv4IGeqw2VOfoGa2QdMh1iMy2hNhzU1rV
nTm/x7is4Lk1lqcsX0/z95H3VvhIZupLsuIiI9xzFMpZhnQDYZxTOShoKgtVBTZA
NyPv2+2Rbmk4LcJMBn/+OvogHIi7Nq2pPUxxdAgzealeGpGCAup5X/cyOBnoe5vJ
CF2QFID9dZ/DeLznodTq+5vwjbPrOKnan11FGgP3oR/qgz3uP6aGU92jTb5z7n/w
1/DdWj+/ip4hQIeJiLr5EBv5G+vsUkad84rfiRDPAFLCfMpAjU9Rt0Mqj67MGhS0
3oAXaDGSGI6LBtEc/b7tAVvrthm1UBUJcrxhrvak/LROrMQggxsTMBYoK4f5HJK9
tt88ZeYQROZA49DHAUwLybU/Lq1c5MpZtXnvp1VRk+HQWdkWh3kg+fQMdnRanNYY
LDZi7m9NOjw7clzr1Dq2sIKg16ZYJeSWW5IctPvYbO22NHc8gvw+B7AUvotTDWeN
91LNHDnLe2SWermX6pBhYoSlF8qWuEHJaPy7e9YvFi0ikwYii+29U62uYT/fI9Ab
x36NIefweJJyW1jew0QGiSAeiWcIMFql+q1D1hFH4Ds5tRg7XkFb74TbGE3qi1Mk
ysnbDFO3iDyzaY4VRFSMeLysLnwoLCFqwBHUHqrWC6+5BAiedeKL/LhuS3UVXl2T
swPsNscDrUowYCDNeDukSnD7+DaptfizOx2TbF6KfeD0I071AljGyNYcdvto+jHk
MTIuJLhw71fZzfz0MiOnheit7VU8kidbc/+CqrnFmzAC2pLnxSHc9vOxLVSZfoup
iEc4E5wPiWak9Kc2xc2xDX3Oka6RmDaE5WYa8kYJwMhgBbZTFg3U7rRzJwvLUlsk
daJ8N8t+FnyobcVJOYxD3ujMUwFSgW8Mu6VjpeP+7iLBPYzjAhwGTkSz1ookUh4m
PcCDEmTXpscoFwWTmJl8PduTJs5sbe2Tb/2jZfB6j1t401J+Ph/Znqdnpo4lMFnN
v02U8Mk6YgvDR8cPc2ilvrsvieE/3OtkO6kvmyo5CwFY4RJRwkm6qQ2zWjtcUNvR
SWorpswTVWWgFo7U3Zqxn0q2CsyB5eVH6X/FT5UMCnODlKE3+j25eI8IhojNIURl
BcDISdQpil9YEtlFWGl8zHXgvB5CSTshRXSQrQL6D12Io1RxZyWpxsUFeGwjrDir
aixWiX8e+pvF9R/YgwdWrvnPtwAJ3rD777OAEBHkmHf3851EiyOZPYKcwCs3oy3W
H6psUr0fRUhNEIJl/iOxYiDGmDQVQyxaoaCQ00uGMTAXQLzRhOmp+I9y65sFEn+j
SuJU3/ENUnQ5b9BCUcgdegzUNAETiqpijxc3+DfmImJlod33Qb+TseOrZH5SpvHy
xlb6qSHKe9S+IBvWVqh7dJj8rmUHi30rgPXNo9k3NIO/V/16BfyjQ6aTg+jUmFaa
Tn4KvMqKXg738nA9/rUC1Aux3W4rysMSthlzFBvSACaw7aPKE9tFADowx3M9kGRm
5sSI8+mXp5Pi9DXsWlCLQ/ujkSssW2pWvfe8T/Lu0r9oepGVEAw00IjrHFN7WjIa
+24X4YVFUjm/q3uOWH/GkQ5hMb6u6MM2LCorEUZx52rEJHE/B1Urz/xWrrz4CD4D
oQurCGOnNKMoKAoOaQ05ySr9/HhnL4IAebGnwwGbsCIjgEluUFqztZv99BjKlEEP
SHXOwWYHCd4v6B9si2HcaiCXkU999XOV9V6OxCKfC+YhT6+ybgyuIom//IeaXSTR
Kb5SwfnSkAe40mi/85ksvOVDebvL4kLVx+Dq1uz7TNnBZKz96g+l5IFe4IIc6h32
c+qvopMQbKyHN7QosUDJ3knfFHsbNog16nOT5wetquuxf4H+PKSn1nrTscK7ayvt
ChSpie5DX5F/JPs09dIXr2pjSBV6h6Pr+MOMgdVXEAoxD/X8bLaiSu5xLq4xmBXi
tk4RqDoXX/OySa3eMjdOY8YbJgGrG50xEIF/Q7UpI8nCpO02AnP7HR/VfHvbMvFt
LQoiB8r7+rc1rxI99sxpvlDsqn/isW3TtEFlBzdvMyRsvL1qWYPpJOjlqAzx0W+e
/y+bFnc5UkxP8r9HRC34EUr5HjBaVZCYX9WZ5tpXPQJ9Lv/T/WJ8OLdH1Mvo+i8t
rYdxVhriBhOlcHbv9qDQCHYfO1nbrP28OC1/O2d5qCAZPlWmkrgMlp6nJG17olLL
OBZCMkk9erKXQOCi8QZ3sHjXUWVxEkiYdiG2IpQ7ZuqA1ybbYh7xUpQFIYjIv6Tt
Y8RhHxMsCiHXVeLGDlwXf1jWwX+B+FyET2dKODfcueGSgZrRwIQ9wZlMZ8FfBH7u
7FReb+CV6tG0+zESdyLpxX/qGwCVUPvzMIVT0rzO9+2g/ea29ujQpiC5DkqS5M4K
JQpiKqmCE2Mozz6btuJNATqHPjMYk892VzLik+QD0rLwkBoqHkcWlsTqsiE7FsJj
jU6D1SipM10t6KR85CrY3lk9+wcx3q4GUla1bBGLssW/segSInp5x276QdILaYCK
WshG5HwxhMVlYelexxPpQC8EMm6lObLnCQ43BaNIYuW+z312NKR1GpB5eV5F1cSc
kF0qM4fU8rdYSuq/M2J99dpyB+lCA+cC7yktZjWRGo0sGgYme8Mo1hAyaJno2dKV
Fhk3r3xNcTUmxhjuLplSZ5A6YcOsA6t8JVoVMl93XPHJERQCuMc0bFa6o197D/ON
zcAx8al+AAICXDOoejENTyf6v9BA6lAHHVPmENkI2m4i51B37W98+j2DwMnEu6/v
id3cd8DUdhMscHm7+lg3sm66iQpHIFfo1Oh3ZsLSg6WfG6Hq/7v1rpM+PKmmiQIg
HPQ48fzI5pG6M/w5N7MRbbprxZieB2UvbQK+u96JlWNVYzLkeHVCaAZmw09M97mk
S1pjTDtcfboH0NJ+cS0lEryCvHjfjNfLLj/p6i/G/2Qho5SgNKGqRVSNhvlz24IH
JIF5yE6K831JBH3UJ1v2ryoCS3jTxqOOktbcqpwb/5EaC7II4+W0T0+So3f0C1Bs
7TY+VoYvsf/dtVfWx2YD8Euj2e++vMBAaGp8K0LC0Syq7gx+NRWeFg16B0Tn1Jdc
vO29fs6Ial0Tmg+P/QwlXzQkWLBoNlFbAczRsUI44zree5iI/bokzwgcxO4KO6MD
/lhAVU7F29WoBpY6QkDL9+70tH3xTwQQ9wT0z88ABHyBgZujSAu0znrFpY0dGNmr
TZWSKZgMhTecOxkbQmZ5Ii6h7UEJrOGlytFM4JysjZmmpXMp3b9xunfuly0NJJzH
YLlk+9pws4tuH5OrL7ZxscTcrAZoeMg7ooTeHxp78YyKSn3E6ofYvNmOO6jBX7eo
9NXizFjPCxTYGXQl37ydH/6Dt9VnJvFLz56zSJ+pzpbPSrMdL3cVcT+ycyCCWl/a
W78zj+qv03vwZ7uNes+KjW0kzLpqtwPac1aOxh1SCIMEM0ArwVXvcvtrnAy9h36t
mPp/JP2gpmyZvzEWNpuL+LTLQGKASaJTNfNv5yP+/LSiftQ60PwifJP+uktQ8Td/
fj0HAL//O7t3RT7EF6thiVJSCEQTimPewHV1r7E2mkOk4tTMtDmuC0cEhg2RmP2a
oIj/ssyntbG3mxzv9Vd0WrgKb2ZiFbC2uNfXhKmxPx85UL+LFZM8VtvrRX/QAZHb
x0tWK1sSikV3GPZc1x7vB/UuKgxYT/PE1FBeLc8imgXljuG/1voEDBdUY5AOqgix
ggLB8J1CxConXqEaSB8hj1zsQGoo3/U9ulcbB7KE6uNhz1GGCfCDROYndlpS/Pvr
9ZhP/UZSeppIOvKitXa0m2U+Cuv6OFqQl3iaBJQBZziml9DpUINUZ0yi/3LVbPeD
X0hwTV1u1ErlCvnx8FySm3UR3nDF9j1zfr5nLff5jO7JN44+jJ5zjKPDXXUOHWWJ
LFmwAgofXZl0lF72DAKBOV9zqjRhB0uu7y1zoWP0xR1DJAeKy476f1c7DLDtIntp
8Ij8nq1jX07FQ2mijB9cf/chiC/7EWsCtZatnELf/AASdjb5NFlNbayHBENkA6wF
0AU9roBFgAddUEQYFvipG3BtFT7+vmtdCZxNF7xOJ8nUMi6lMsx8q+z6P0WSNXJW
sLOTE3Ki5x1c9AbhwOi4Dub2kxn3oK9DVcklWaxOH8/L8tzlrFbqMxmZX30uyAm0
Y3+tBz0uHLa1LxVWIGFQunWcmXwBtkN79s+hZtzhY+oQz/YiH2cS5wluVWAaiUxF
spRrKYhfd5/QKd5JnrtXOm43jKSj2FKd/IdujhgO6JSPiOtmxGEWiJPZ+DQOuG6Q
XJwhfaFONuwFShr8il/pPhEI/Zir22fE8uZycKzjgTzqSB36SmD874N2Kv0LHFL7
Geta75R+P3GanmKLxKg2uGGYkE2aUfcS07OC7ztHbZ1+sytNtvcZwkIT55woVDSJ
IhceT94CnsHo3NjdYusMl+fyIRUMPWlORGhQsYbd6nXDIRWrb8c1Ol0WItof8wfy
J+QSQ+1cEGvU2sdp+UHvJwcBIhOLkYZcM4HfAdMSZ6J+CFPUjCRodT3A1riwW9pe
vuiN8BJYpTj6MzeUruytDHW1vPOu5bFRKcwcV3MsHYBQZ4uToHAAyryOn9I9laRj
BEuG5L7Jy4XzrPoKjciMPbFf5E5HdOl19v0QGDZX5FwCgvCsQrWIhd8l85abLZLJ
AymOKP/JFYjya+t+1gaB7AUqM8ivJnWqon997Di8h7PoO1jJbN2MEkX+sEVFoyiN
Gy/U6r1dQxPxUuFA4kD0/Gv5KMfq7gjZXZsDwH3/lTKj2KZrEmDzKipiyttTE+Xt
Jee+hy5b+Lfjf1pyWRjBsgge+v31PTYe+leekCUuyMo9ECGYwpLTuCMQR4R6cqD7
9naCCyQfCcDV7On+B9ZV0oNY10JEw9KlvBOC9qk57CddMMV/+VDNYpfxwBIYA9pR
cpZ8fiOVnoTNWtQKabTwGpF3p0XSrFTe0s8kI7zKTkAOevAY54Q/iJZ1kupDPd6h
4epapgJg8cqoUnSZ7857x69/9Qu0dbp/P0Yb5EBLQCR6UnvgIyfBRgLiFNITpNoq
kjXqdIkkM7doo6d2QlMpnExWL9c/L/Z4N1vi/yhQXOTr0hqaeGl56rH+7AErowGu
GUUI/FVqVYRHoXw7i9NNs/ssujCXYFDrtbkO9cXha+3483coedHTI+NHaSvvin5p
KHtMqP6lACP1fQSvvuKJSHbgI0IHXyFtdxpTQSgY4OrzNz30vMUAkxxNYl3TmYW6
EHQfxh39faNM5nSNAB8kmwgrG9GY8Xl7LEwGLO9odLzhZkEaQ623ALSpkm6EgOPP
lmHxQtrO+cjAELZAJqrXT8jank9ESqU5/+ZF5j2QdCUNxYTczROmARJ0ZdnVZsVT
Ixw+B1C+JoSQKhNnDckcPm0dj3fZTmL58xG1UaiaVF5xMhrJa8AlSWozyzML61EH
YLl+QmUaq/Sr4i/aASdEGd1r7p+jo5VN4RI0Nn2HyMZdt/ZqaGsEpMMNOlwWXMfT
Oo5ppxTeYWnz3QkdU8zWPgPLwYw7HJnMi6sUh8y3kb7iFT3D02L3TdOzDyEX6PH+
wLfk+qnkQJMpXnABl34zVN+Y5ixsB9uyWnwY9bNIeP1HKPayd3JS0pE0Y4JNoBgI
LWgm7zne/PcAYIj+vLKMtSDTXSe9Tw7BZqDGMnfZ1D1aV/fH1LV36cU+MbMbLRxW
1vNwEwsHUAmXt6++uiIxFG4C2GHzB/bD2STOnFvGyW8tP/spcZogHAUTg6ySEzl+
x3KYfmoMf/Cape7KhORPSkQAuXuNeyD8HX6mHCWxs4Q1PiSmj6yDvawsQCEUrbJD
6nKNGeoiFsWgivSHthUfQSdgGAwcyUVW8Z1X/aNi/J61Emj1Ldx51dgLtJ7uIeMk
l+uDxM29xL9/B0v//HkyI/Ys9kuRrxgyqRR8vOCiazXVTutbVuU3Vp4vP4VX8no5
kWFuNAtzpjD22pt2aujWv5RodvQXV4CFWLGIxCmR1qQGorRojHuxugtMHzunxKDb
cIz+/8wPPWTUzZTZAxWYXFgfCQrMMwlcv1lwKhmjnRhAC9lV0tVOW+qo8zjLnd3H
I9TamN/nxuAIOxOVKjn2xxfR31PukERRj5rV0ghHJ3OvmznduArQpzOFvKRjyO5W
J6iOcbrHir+hBpYsxZiLxzE7cpzrjaF3pubACEoCzUpm/Og3fesHvevwVuJEy4iG
X+iiB8npAISaOy13mndg8MQ/5PmqVCGXxB2dE4DyOHhylpo1Pv+jR4+X4qna7DLH
Ul739JIQQ6YtBtxP1kBroZEjZF70ByHAG+BjDP4H+FbhGlfyHYxkDG+BhpsdcFYb
pm+4zt0jfQ+Z/pTJ3KwS42rbO6IZ2iUHkY6xjWQfH8l1fpLemrDG3V0hwhvwOOHN
CqfiN1wAGkhsmMkg0weF0vypKiG6oV8PjilbJEu1X5NdBNhOBEUfxl8lSkay8rft
2+eZwwxVQhlgpXf+aLhREZw+pfhWgKgKJ2q/kTSocOhBaN2mizsE+H8gXTGXnX1s
DzaOvGd9rTqumM4A+TH7fynocWqXL5MglodO8OCMeRlM+D2KC0Xk+aZFBaK7Xxql
u2lctdCAdUjuOJREWobkQTozz82eG4wC1mhAdqzcgtbtlYM6VwQXkiNYevNlNy7d
LlhIi9fOHyDxOt6qEChhKq9mR9kaYBKaunVjZBGXldv77luIbEDiP2bvhqKUFcCt
1QbkvdGGSJpbt3qTD+p+tLhKkuCLwj+zSGsA23x81JpqLePLfTI0mh7/XEduZvBV
sZz7h3KSjGv/3HuON+5QoOFgPWa3UTzESZfog1W4RKw10Tnzf8w/teu+T3xe7M3h
w8njEHqdzEbSwyLJDvp7MHK8c0P7A6LmJcpJ9RWpNBUp6OVZkfWco41XieJAVQg7
Qz90CNZID9Lagm59zzrfvzoYPn/89ihcI0MuVJkTqogrrzEqsQHDWnQulCgoWDBa
5EzshFdd9C4o535MbYPIWSxV+ATf7Jru3Vpv5cdnAkz7taSj8satHd1vsjAB7qM6
ab2V1cUw2ccZXuFDoFCtalLHtp3ywgE/IS66OHo0sjbEhU/tNyXERrfGC2Xi9PPm
h/LBz8+yCA6jqwhSLCawuiFRf3mbLZTN6HesVyEuvgS+Hw0pBvbNPHgRoE5dgAyS
VOWI0A6k9I/spc0qV1rXeKF/QSHe7/7wNqx7PAFKCBdiz4eqYypHel+2iJEd9SDa
UDeFFXqTuF9FyjEEOKcIevgvrWkKcKULdz79/0lCWj94xGL3hu+2939QebMwLRdL
v0I5kQR4eaZMLxIqxccDavXWKiDkQQUteKov/fobUv6ZRy68giEfegMP0Z61kXMc
EBEl51X/AB3UA4DJeVAw0XA8WfLpS1YiHLH+y+k2PncVm1OcIxED5ugcyEkuXIp/
W5a4I1jH4zeCrVvDdwK9zcbWEEKJ99dojM7g1S5UGDABRnqwm1kL+5dJBG2DTeN2
n94r85k/ODhLVrgJC0DJbAhSoMpLbmngF4NcYytWBJWgLJUOLCLy2jhcBXvqsH7Q
o17IkfKIJXACLh1Y1DsdRrfrZHHu9WAVZNHwUJ2D5oXdgKk74BwvqDfwvj8WSAVQ
x0BUJx/ZW7tqieBPDMcygrD8+ZChYcFTHjzGLsGxyiSSubOYzDcWq0P8VO4f0EdR
udyfID8slpCMQPHU9AlZATTBENo0JFdVHtBXFLfDniLf5Co0gJoj5CjuqcfR4gmK
dvL42qMJgdCo/1rW8/YxEovztwyhQ+MO3wDYbDnIp+cVv8YCk5YcurBUhRoDFmuc
8b97LJuntdAJArXS5izS99GvgLF9Q/7/SQXiEPT4B1KsMsuaJHV4f5Y+I7c0m2Hp
/h8KnndVCvk6b+4toyq2ML1i74hQLZtzP5qlbEzUHDe0pJt3YU/LcrqyKDuekAvk
ZwOtURdAw53429UuQrPz2gPahLKtkjC0RRY0IQmJgTsq2kZ8i7JPlRNo0Yt3DLqY
/mHyv0A3hj4ycPWvFOTEtp1n/NH1k8ntEPN1mEqD1eexNhyON5lnK5fOiZboz2vg
VRoDA3hc8Xba9AlX7cz5EOLoJu/h160qZ5OwZxxKmE5kSOHmcVbNikVWdCMfGP84
UZNvFvFnhN/Yy4DTbziEluaz6QQenUgIZy1/szcMrqOhwb242qLhLVlY5rL5pBpj
5c8k/hbcMwtIQM+b5j9+xRardf1v+1n/AG8USFpQvefRUb0rIuUCIhpWFgCeuOSo
12GvgYg/23Prmq0zcxm0p9zKVllAXDxjHlN7fxeI5pRGdsMbYvMhlCDdOWMKZDUo
oneHYsnkjUUULZyMRgfmtV+bL+Jk1EenM9Lq2dIOwgNFT1YUaKLo3AajFFRRIkg8
S56DGdoX19BLQMyAACPyeKdBa1vdh7jBGe5SHmlwEpKbBJ0P6j08BpOngMmW7IkI
8I0VECc/Eq8uRoeSOZT1QFSjUJYIaBj+3urMBNeMytFosj0QLflqdgXDi18ZGND6
auV+nN4g8ILI1nOZzZ/aFh6C5u1yZ/QX0ne2OEdasmSBIDqyJ6IsCL6ptkL07M9E
+s+eIT9JE0MWXggUCGsP5IqhXnK9DOx/BDabhDJs1mjS7xQ7wXjOFC9UwEuQfMwx
dHK3cCJezxNG5vpECYbzi1FOrW/TCaU1E0KV4I/iPGTPJCzE1iG/iVsM9vi+35AO
IB/Gk+4/sSuzJDdoiZWRsb2Jsn+U2dd+ktsyRo/5Q1kM7jmQ295jfLLpgr8Bt7+C
GYGC2sPL2Onby/jfb8/yfm1m1R82BpZHKWSeA+UYc1z2OOTvuVfk9rjDhSlZ80ON
Slm+Eph0vTPlPhGKZICr2gSBAS/WDtElfE9h65fF2uMn3Bgw5zo1psglN/SuKCxx
DTK7tOuUEeACAGVFG06R1ubbhS5ymBjwQOxpPKj4fj4XTwt98vlD/TUiG6lTIt9y
/oj/fmi2FeAUOCuz0RLLudYH8ffRYLc+k0FehHHS3ozhL2FnymJlQTTlRM5IGaNY
BYiTJxofpdVtMJMl76s5PSRs4ix1bmeBXbDKuDIMNGpmSI2AcLFBAefcgf6m+gFx
YsGyErK2LQ7lWN7akwembUMXHs8PSrUlfJvYMQR16jl0v1PVia3iy2PGsYpBtG06
m4nRzCpJrvyCSOJmRLCoQmZJaXxjoPcsI0Ry5LLaKEXWDRvfmKOKwFfUogyv3Xao
VBhRxxRCM6xwcnLe8URZdfsl98I39XD8DHg8ts8wsQZshXr/R+m0Ktl81eZdQ1Wn
vJKBm42WxTPDeskJn3+92JReMYaotSHUEPI4w920763vsTyvBVSM091NMpWjhqPc
4etpu58tk+1FYVC/kY3jDXz7TA6abIKdoRrt8wYiF7ypc3VR3Wq1WOCw+1RGqNBx
5OilSXSitz7eesraaWVbiNh/55B956DS459sxvUtf3RlBIZ6jULK2wq9tp24ZnXw
nWbZlPi3PzdNHvxmoG28e7Bn3fFv5YqItR0pWaT3Cx011GYW+2PDzU9cmT9GEWll
OlCEMJI0lFv6nb0Mpnayx5hFeeImTdRZlU8Dpglq0O2xFxFQzsyGid+73e9Hv1Wj
Myw4E5Ion4y7opjX1kRuNa+pUGDVY+dSjSctyyLW39ZZXFLz1jBEppObsYdmLe09
vjBCpO4CIUWRXoM4IsoTUicRlV8+/Rm34jba1mneCSJHe9rzEYL+OakZV5V6UyLM
h48iEy6sGKUwZ9i5iqsY1RNSyS4p0/akYxF5W5YwqpnMz2O6UgmuOVHU0GQc/tY5
rcq1dKRGEkrM7KxE9Xf/iFTuqKJiuC6VdEtBrqWuHwvFfLbxr8qa9BlYOMDNU2MA
XnP6Ux1ddT8D1p06fgm/VxK7vLCQA8UMUb54hbqgtrk14jYRbSZ1golN/Cs1mDyG
wV0Il1j00yBWYvnGNpglpej8NUHYZ0Xi717PsaKeN5zFcwThnukkiJpYv+jr0fWW
1mTgMsueDSt+tvhj0AVCB/IMr5NRqTHdoElUzC1TVrG3WB+cHLGZBlENXqphVnkl
Q1z5gnue2edCuy1Ckz1XxaS2rODW6ga4zGrgaHke0jxrf6fwv3AleXXfrFogC7hl
niqmonNFFSWo69aSXAq+yXzE0usoiNBCoLRjQP8ObbK7eX3nnr5zh8RzVI6HzM8y
Q8dhaKqtoWXLGElug6ImP2xzlfMreNq6ShRHFMQKOIDjy9oDPx2bYW5UC4Tji6zn
fJLVPBhkrIwpUzQS+JHUz7Atb5gFw+Wnb05S52gisKEj8KyNrtaCWdQ89zy/cY6p
0CNod6p5MvDrZ2osMfd6TrZp45qCAjjkPI82ZMopprC67+DF5gQT9zfbOqyHOg8U
IjOa1NLw2Uj3BidW7mplH7nk1Hc1DT2Lw3kFhJUone3rnh1ZHVRyXUww2bqtCZrQ
Nb6RlZ7NkXsmVxtmGmDvZUxl2baDrgzTxaQ/fMPcHKY4Litm+8OGrOEui+TyLsQy
q5bKSkrZmWEvIZQAUcOUmzp3x405T5EWNvNH+3Ho4QNQqBX4By/WmmZEtdtPDvtn
m8CD+Atk1vNerN1Zc7GC2ThLD6PW5Nv1t+XB1q6Y9aT9rR4xwJtbMnaCjWpK+ob1
zDVmCIAysaQwsTri+k0TSGfyxfo2lZwJCxpr/wccc3JDubuiR9x9KpYE3/Bv8Fd4
QpP6/lNTS9PDoB0mNW51LPJ8EegitZ7z7QF6VMRLvV6GI/VmTd53DWaswxM/oiiq
/4Js9Fa65P6C34u/1QNf1L8ikziZ6HPbOiSiv5BD52heR57xgNe/+PmzRREL3khh
beusnabd6biUM8qxJClHr9FhhMEJK+37hZPJIrPPbjc6KykJGwC82NQU5FPf92f8
4rybEjXevu8m6Xp7W+aINzSuKILMTRSasCQLZkbR4K9Z5DcDm37QpBXGYqidNNY0
LxZWVE8GioXD8SSiffWHFpobFWdqrPMwvPha4Td9vlyvV4haZ3Xe9KCOHCbP66qY
aLrEKAWlPCJbw3R+CNdri+SC/7msTHy8lCkZ8WZ1rQNkqd8BdpsJBwhupSgXxXef
uqjAOYP1WQaSuocrJYIOfN4bgnTHtVwMkBd44V9Mxu4HUoTuzcYlxL2vCkcgH+5u
u53DpwQ7M5v8SNM1zu+5g4HTPcaagPmsJaD+iLkfjO1oinbNZ4rdD1H34KmsqlDU
6/TPUWlBdLK4Z5rbMYJIY8P5U0mhZiWtP5OsTjda8AeLG72Rv460WiioXejhxBNI
iH+Maexi3xZa3N2jwZuOfqLtMtGP/TnJqGgD3BNf1YugqCCqsEcaPlSk7g+PEDg7
ROh+vSTHVE3fUvuTmVem83gi50yHl0LyZHhyfksJYY9OfYGxAqbMEHKurvMOuaOm
IK5PgA/TZ/v7/+IKeAJO+3s+dmkNZtew7yG8Bv1vvd+S+oFckmbMiy4Xj/GUeL2j
jKPn8ILzg53TVbusIa8QmDy7fsfKQHelw8p/H3Fxl8uP5tJuuCppAnW9LO2WE+uD
iwjuekqC5GHLI2rIORLj4yFmopGq5eJO4KxUNK6yOj4vug6w9zWE1I42BorzRxaj
vbfE6wj6O8gvdPmL3zxhM6IZbkIzLctcqZNOF1F4HAne16JJ1bXQtBIObFtM3J7y
SFklKWpdcuTOa2x5PfrFUi9Aarl2hA0I6lUTEYse2VKlZCLaKD0Yv4cDqB4q6zyk
AjhRCx1hK8XgZKEOuZxoxle0t96xX1OSf/tovHQ5BJzz5gIIIba4Lzn4I+pZnTqm
arKvMd+O7MzQnVTk0y4tw2WIiELxffy1DsCKobkYhRQ1dX62Q+rKj6MPt3poDP1N
QuYxdwyjHa7EiVDOBOIwts1ruRHUo6NZfA3q+SynCRrUzWSyN5dyYGnyP08USX/I
e7BbWiQLxk3EPY/A/SQhFei13hv/1yredKSqnyBN2ecIES5FsE3/7YQtjjkGme45
u9efsy2y/EojQvC27aJwa2rRJBpjsX9XEIpf+5opzqVfw7X8JFc0xTPHsdcYX5lU
uInovMME/ZlgQdPcfHNM9XkcPMzm9ev0f+aR1WPTUabhCQP2O2cUcYXA0QdRdJEZ
l0lvr/p/8J0l2sYMBL0k77M5lsubSQ8T/PLp1mZYmM+Oaamphv5DLZ/vC9uArqfr
Ug6Iy68O8ZsA3MfX7pyao1K5QaNXZSSii8hPnAswq/hJpZrdkxOMgH5SSTcL08C0
Xxi3sElwkUUG8GHSPPeQwAVKA3FHFbAS3Mm6ND0br1Vl9WRrE9ONVdj4P+NwQZah
0ydIKLhJkb5ZAdN8hGaZU0ksOQp/Y9lYnx4dq4DdU7CVxQNKnzeQERmC8/7SYnOI
/13qZYqHIrK8IQ4gYre+LyoSEs7qHJEZ1Zj/+foRL68CvpW3/Gr2+Of7wvINeeQ9
tiYw0iLJtsd0xXp3XPzMBWBfkj9IjEjzBcHeshaVP1S6JtB+Avb6iERgi75L4sUB
5RQIPGfjy5e/x6Tr3+fhbnk+NMBSong15X1T8EHAOhRPjfB3FEipwuTYTXWChtKJ
CE1144vNBVW2a3Z92w/KfhtCTozlupQ9gXUMO9X8jgFFG1BkQu93RY5H4yFHoz6p
flMjND1s+eN0A2LgUrXEl8L1gcozTMj7CBIAlXb/4lnsrBi3KBLbOHgUOs93DkPC
Cj47RATYwuaEJKgYSJOmMeCBkUmkJusBe3GJWTCWFoHo9vlvBNNi1cC8S8WcsWXM
daFc+ANDnzqaorrxzGNZmyNFIDWWJI4c4aDCyUsVywCkd8VFXQgdOdf1TTAlMKbb
+7lMZ4qp9jfM1gEWGEiTNCiJvPb6UPZa1jM5r6jQpMMoTR/2kO8rO5ontKDC14A4
VXxW/MC3A3GMARpo14uhtDBM672Opv4SOno2oleyeXoB6I9NJka2nOX3UE/0PLCb
kqY5tIgE0OoKFYwaat0uvaDnZ4bPJrCmQ6XmkFgaVhYnahVF+EgODLB2R607dbJF
JfP+TAAkhVG0X8eHiPnFlsCMyekqsGQRrzffetGqbvLt0nFY1eKhm/Jmwct6ex+Z
7KUPb6qRA8zpnZecb75DmZwJqxyUHno914h7BVXzqq1v7IhhuRyjRj8ii4K/uZar
g7EGXMzbmy7u+ApIbyqN/21bsINI92wKP6CbYUG0iTVYRoSWp3oNt2OIQH03mSi8
pAbbQxnDm25c+AFD9UR2tZZEVxf3Xv40LdayUpDwxr9FnbdaIt/Ea3bfkHCJGLrj
lGzsftRUU7pgWuril827rcWZwNB2HBqL8mHwQXVIZU4JbX8IHI4gXPFCYoSs5+La
sQPvVEUV8u6hBgkdoRxKINFCjdi58Wk7wEYPTEieD+v3o4w1c08nwhswS9ED1nz8
v/D8A6Oll/57ZBPtpi2GdMvJhg8K0rgdIrUtpJO9IK+KaJ5klik1o59cFMqzZzwb
Z8+e1Pxre9wz819oNNCXBSBt7a4+wkWPFWUNSpg3E/IDNYufqAfMotveMcEXrWeI
SOFglfoZoJE8YNBPYnh56o4tabmDg8iBL7TcnN6oQAnEjVHHlKNPadBOJXdpZQ+n
XkRf+kElssqX5FOS007VrA0Dv6mpVrl7SegrHJpolTJynYDxVnEnISEkDfZOq2Md
nUiNL/kYmHhYi3Y2fdDXGhSwNhTFN1tmOePea1mnD2/NEbvbGYMDaOvHXxzU/bao
rjcByBl+CjQkW/D1GlqkDL3xonob/deJFm7qQ2OFEjiNh12oQWbg2gtJsDA3efDm
4ep8GwNSMJmmepfQmukNComDHpUZ3GzGrxRhbwCz6Kr3fYMvj4G8jZr27cptHGSd
V/XYpK3r1msZ/w+QTzqymWMTQq1y8h79CEQDxnlLwdNEgzVWn1iD0DwRajYistM1
EowEZptWGiSrg8w/Uoda3qOqq4yMMvshY3YKOrLLcNunW59WOcfweHRz0tPKh9d8
DRu/Xr1ZXUHEPA3bg1vRuLBOIIRvjLtfWKMSmZ7/to4fRz9Qiw3kKA6VtsjtM4eY
xcz/DNimmgK0KLxrs1/OlkxeQsKTjoWE2Oh3Vm3Z7/A5opzIc/xyX+o6xwRYyO9a
gd03z1k1MKR1/QYKv7BJ5p9R/KqdluPqc47qCs9D1+/m53MYfY+Coq6ydqmsT07u
CVYC81BwEw+Vy48KKLRev4QL9Z9ERHLSL3mQbluJxjsP0/hkTo9QDNnBA3sSUpnv
1bHpQZo23pm0amIXECEWu6FiQbcOde1XMtJycCZnMx5caKznN0E79QfYMPwRQeuq
iz8rLXdpMWgKTQj6FNAdXmlzFdqQIk0W3VrmsVya43px02HjDh4ElC/CmSQi9dfw
6+tbZyiIhlBJNX/wmUdjMYLWyw1Cmp0MF7e2kGbbcDqYyQJo4tR5loNaUBsGSSOD
1+z5/kV90G/s5WnDURTKrfZWBrNZ0gcFt5Rw2HkAwUUBdcptNvQGAVpdJLD6I1x1
U3XcgPqdnrsWL8dXW0LiVo1bBxrb66TJFVv/2yJpdYq81uIEbdV3lb76bVvrcm4Q
3o7ZgDUSjvZXsRd88bqBO3gxiOiG9kKNJlQhX8yKhdM35DUmH3yUTO7ed6/OVe7n
CpWKXF/dDh4k269MYaoj57SAuAwOsDidouBNNwvmFoynMgcygVdx/4AZYXVVsQjX
v8sa+YNS/SmZr1Di2CBDYeanA/hiaZQqVldbwJwEr8Ih5GjAStREpjn/Gp+SBHSJ
w+SiWxW1zB4EUlPdkswvOm/jCD+MTSDvJ2Po3VEthNr4ljV8hj/YaJ8INE8mX7zD
gBXkB6Gr8kuoMEZqWQr+1vgrMXQEZIdOy5H0txSVqIBXt9D09/Xlwiz3S0xMSYwL
V3czTpqUaMXFrW/CKEtDhjLgmDvoMLRrnA4P/Quv+6rkvZOVxz2x5viI3n2q+4Nt
R5nyDxbSQ4zEHne7UnZYrgy3dkuKBlSnEi4CJD6TC5IQz15CBKH+7oI89ys5LXjO
WGKeUIzK9udyZKlGXKhGmEhat6iaOPNFuCiYehaEw8014jMa+92sNpBesx0nFQZm
3OePkisMiYPZWkgiYJetRH72VxHv8hsrSooI1g/O8TbAofoLahGjh/YoFdMfYgtI
hV2ZgtITsJtdtZeLQcuUszkiA2bajqJ8vyAQ7/rgVnQpTIvQpIA4yWsKBaxnGsuT
hhpD5JbL1mE8bmMZn75sTRISpTwviVhphgiKh5TojTn0sSD52c8H+/vGBI1IVH0d
SPD0a+ahXBo1iir1n9AxpZw16a/EhIAEo4YeiJC2hIv+JZ+2mQSmCxWMGlQv+KvD
ieLxduP+v4+Zc0vDHFQgHyn/KM2UpIlOnqr2MRO/JTQmukldEVllt5IEHa/MTdkz
aHEZzcI8/ENeasfQ2e4JNibamquoFjbFa3cQ5OklX35dlatomjFL7RzJEQFNw57v
wPysczeQHhDjwL+P58QHcIzaVUr+sE6wlRGhCWdTDCcrRtdydA0g+ZhhDWK/80uP
uOGFKLiKj8B8eKdbM7XDwtx2ao2c0oDqZUp05w7z2VAQ0H5IhCQ0xT7ssymgPG0z
8odjhStvWZNTwTdVcquG5FLdCy3JuWV0CwoaPKBYdkqSegRmEEKhoROIrAhWgd+j
wY/0s177uEyFz87Xif7o3Ta7UfXlDHWOMtjAunGB8YOYNiq2xG9AvkovH2vv7EtX
7mC9w0e4HtdN9C9i4EMUPG2YrKoUxJfeVwDJZG6eaCk7MxZircU4Ue6mDw0d8tmt
kHTD63HdisFlQNEpr1RggU8wmCQVpfBt2IH7PYh0d1LezlglwhHqT0Bev3HOQcqb
1pbFUukjkpdj/FvA8HeGPo1X09zl6EHAUCzsGAWP1l0JIHSaueArIegeNasPBFK/
JNmCwDNQtRvCFc/Du1hTrNWjQnPrycBrRTs30bM7r/xjogGNvShtbfgBOBaK/GYG
W/n9+1847K55WzBiQMC9B9Yj2rOgRXXzwo2kQM2YTYpJE4Jk4xn0dclFz3L1M57P
0nXIoCvny2+xxK4CVg2FczRfa7+MUmnyVUmygKtCc9PjIuL18C9En7GKFNLwZEZ/
cpafTtbaqzTdkZOssA5oepweyGEZ2P3l7vTIdg8Qvpp9c1KzviGQMWAhlQ8+RiCE
oYv0zCggLrpB62hrBDLYvSZsNxhWVKoPhJDgdo6jzJ8YIlbaZwXKdNkDcgghddBh
8v2o+9VG7s6XNriX7wORfRNSrPf9LiFTCF8aJm0T2yJvdmz61zW1J7TJOD69k1Vw
lHSO1WYGIiCBLKlI8A/oMDYw5gTjcjqP3UJABslXUDpgfr3l3IWi0a7zfNpAIvFN
WCdbnMiLy+8B7ZiXyOnHNFFlX97Fk4ae0fP5YKkylfyxqz1JJZgaYL7Tr3aayFkk
l5ofWIjrupTqvnauPt0QtyTKaqI3kUInvD1zKaR3q719KxCzJMHppM6fMDn8OKJD
vajoLexNuX2I2G8DZ6bqP1aT+5bI+grd/aEq1XTi9NexwN22WOfb7gAZRccQUZE4
Ggl3Jar19Vj3yY5kgtqVmaX5St8jSrDVmjf3BNoImremfbEVbmKgxKX3YTITQxZc
ENsSB2RvO0UzhMC4YNm3G+htjiBE1EFzt6KJBfWfLzptcfff55Wvz4+PBdQjRQbm
2W23+LbNBJRfxEMvPQVqLm7CBEbfzf0bBptF4W2VKBdH6aVCxkX1Xy3r2AS8G4vW
ZQ9AtLsWxsCrR+TTHLgTeHzO4zE1lXtfDyXeJ9OhM+5rw8yKb2YoLkZxwsKpvaxo
SSFB3mOddMWC4VI0qSxxOhmLjvToDAQ9zJq+XbLTmxA03aLqCz5oexogkPmofnCd
lGRyA4tvPB/TahtTuf5gyVOt2XbIAuE+bK4IBh3UT68IKSOje0j8KW+2j/RCFoel
C5k20OtpZk2FS29ZFsuN5gPYkGDtb6lIy0In0KPvLZVY+rlWdMfavXa1/R2CCAwV
OmKKa9vVAWKH9rz1+OacQ5ezl4AgmxelmgLRja65dEulMuZucFBa1uWYH7Nuz1VQ
jCfcGiNHOuAy8sxMo6Lj6xDKj1/UjL7y4lyMRAi3NwxtwqdTaSoB3O5zCRls+kiZ
TBZdXbtRSPmdRXiBBfcO/YXZS6/vrhUjmGbNIu6l2pMT929PsQNZP67+1u/Tbuh5
cPqhRAJdcwLiLNahfH5SqrzWGAUdWXt8gv/fsxJK/EoZ/oOrNEibHFzSAqhkhVgD
0FH2PGumQDeCMaRAX7Wh97UX9ewDDc/jPDGJqoZOuxzEtBPCoR+Y8pTySQlMeTGX
PLRCJVPgsi+ftV6FWtjwOaodGjqA8cYz7nqX5b+hedgrOiyzWdMB9xYFqNAzs48C
1LdoaAl1NOpRu7fBEp12IeZ1QcSqBs5kSeKSjzmNBC6pNX4kFIb3DKkqVSTjSSFp
EH4jyEI62Ii19iHXhz7x2XOAuYw/oY7QPcxPsPQJlwY9c7yaHite8DpeuyKPmGQR
q+ITya5hACdmnlBCaF4iH0nkTtehqYtUjb8hh7eikuCz8ajdA7qbfrkuaKJnMbq9
1WTuo0AhCO4CoOd5ER4nKmq2+TBdS/95FFOFsByO85xslfOZgqYWulJNEHhg1i/S
RMw+T6Ln63/WGBH91pdi+I0wAqKxiU+/O9ys3e0HyRO4jz7lVkStM4N58vhiViy3
O+dMLa1WNDspTPXLhwO52grr0NwFhh/ji4LRWncjcNYdlVmc6fzXSslY8/7BRKs0
+/RX/KqKcV5TW0t+8gFKQIYjuFIDbWA6MM71h1EZt38gVXwp7+4WjTeuK6X4PQdX
krmZsMkxP0Xl35id4cWBaB66NM8QGeIN0BGM2q7un3eKBElcGiZe6V2NIFQ/0HOK
5taCoYXrH6rBbQXUr8OOrteGEVXdZguGSoLR2FpbUhCtXWbCot6KSA/poCZUT03b
0N0B8wIKgkQlG2svGXai26WQeKWKy9BLShCdBiet7X+XmYyfkz+VW5FqJ+YYYACE
R1TEpWrbjWa6Rkb0cLZ5i1CzraZaxPT/YuyOaxnyGzSjqG8tSCTJOvxg1ii6AhUn
c3ygly4WAGtZK6krLE4zj7uqdGy4HYQWA0McFFB1iP5o3cLGexXlrMBH4da+gQ4d
tG/e0Z3q+HU1joLOg0Gnf7rZZo+o/mPcBVg1wHJTlqMaIcPtUQSAv8JAkIJhohPw
Bwf48nNtbJDK4009gnlhXe7KHtkKwoARhAk2aZWCVRoa6Yoz6b7Eids2MOEeIaYZ
Q1CR6loWjw2g2ODhh7PCSlA2bPxSxesA7GRGtIlAkzrnQdigK67euabcchVNsDIJ
LpBC6Rw6ep/ZTcPSdwf18+AsiiBV2viRqKGi7xpSOt1HltwwXObcPoGhVfc/yK/S
okldtPS+tbPscYKVAMj1uKPrcLGPKtp6bnPcgvuIVZQv53F1gxdXHIID5mlbUUVV
FlDYzBDthEh28cOnw9DHIi/dMMm3x5kPbVgCjFXzMCQEURI3K+q25vz+tFcm/5Md
/t89/8tV6mWy57XtsYKdjaJi3zGcFY8y+kU9Hu70Ng60qnSCgDkPi3JZdvPKdHGa
aLoayK+Z3FCm7ZemrBlzGgRAtZ99onYWfOpG+KeGJaBJEYU5mlgVCnZlS+C/Kc4C
UG6v9l6LMFV6edjuXtW0RUOnZtpmZOQUkUq7x73tDXfUup3g5SaLkMTEUu4QzPx3
au0jFi0LDC6hDuPdKVt3nBtrLdVY/3kp9iD/jMaxuekEDDCq3V21+v1fBXlgg2Ts
7PM7FB0rHMYLPm61/DQ0MvyIb9TxglZSZK0rlH6nfmMfjE8la35qvp3a2HgfQK9B
vF2+mevjAxaxXwl4szbPIUUIWRMw9XHNA0O4TeBjWgLknu3dEmZXGQazH4fXSM08
pvwiK8fO3kW1WruOJuvqQKHAwPX0YHR8aaIJhtvKCQws3Kmizwcs3kDrQAOM10yj
TPUG8PblGVKPoxGiNj3nVvagrE/Hyhhk9jk3H1a1EzjEw8SoomBDYJRrTWJfSW3H
Tm7M9E2DItRZMArOZMyXQuzwejm76IWI4jLuGH/NEaTeGgSupotasXobHe8Fh8yr
UtWe2quOLmt4Rro4gJ/sZHNacujsT2zLgLfEJ/dBjl8jAMKJ+9IuqZrLvuAjYSUf
2FV8n793V52HlyUi7A/g7UEqtpd/OjeC5sXLEakdZ8i87EBOcT7cTbsdMwbDs//7
zaXdVLbzHQNiR6lQ8P2dE+FyOyDS5Pq4RP8EeVe5UoCI71WHeYHHPndW9+8DsahV
aumuxtfSnI4LQhfVic8mjqFD/U84F8ToPYGHDnqFXe0FMZ/FTHywwvveIKrlkTP+
u86psfXu8T9Q+be6LvmJFH6WoWZ2SucY/Vr/oZHhJE5+zUNgBJMVBPYBuYy/wxdW
TLc6JuIuszLaZ3alUv9UK+4+UFs8P4cQESrtMnO6SZaTSQILTFwF29weuHUWJx43
RZmhXYOiiuHUhea5Xke754RlQLa5/eMlT88yr1Np/moN4m9XwDkgsmT+OVF/HYYx
k+TwGJ4BnLh9NzRXys6wauRAnhPpji0syphSl1EpJg0iwSWjhpxVNR/4I1Mx9Stc
eTPcV32TRKv5+2LgmrYIDdeWW27KcmGpjz0ysZiPUGeBTtxRyiEDDtiENhoVf71R
FmVnAi4vKeQJ6c49SFj7czA1vr4m7M+7LE9Z3y1xKmy2jRT9N9JiWrGGQeNtW1YP
Pqx9vO3svT9eyenGiFxnZQuFMQHTaWKZZaIRrDJNdhTLQmiR5M4C5M6SiWGJIFK9
BL3VBUobdro7XZh+bkO+Q1MLWDZmrVVIRaqIenNqoL6F5fn4vhvHSsOASkqD56G/
P02Cpix6TaNe98zQhHvrQBsnLkbcaPCKYs0hUIxHCv9eNA5xy9Bo0aSlLuhxGd5h
A83jxGASF6S9R+05KBRtQEcgApEaek0dStqyQRGK2tLQRXMFDCq71l4Wug3rl8Np
IGqlS09UrrtsCxxHq1xHSWzFj0vvXaf7PijhLaEQyLjvKbIfvEs4ybEkdrIjIA82
3IJg7qCtxmyZS2E09nffgfCa3YjYxs6Q2z4l3Y3EEZrq17289b+wkM8JIle9/RKf
zmxCfR8o+d6faDLXLC+CwBvdEhrvTAlh/Qu01mNPcB2fb7ihIrGfd9vCXh/YBaWN
kmRFwNLZrKVT7Mb34IU1YzNlVZ5OuTF+KAMBouPHICiNoczlMNY6JC4bngC7B//H
7w7jjuicEuwK27kxydv6YL3sNYIHj5G2U3gesKnpqgQAcaRhtUFu05rN0ILv+lUm
zfuCewrmNjvZCDG7wVLOg303BrHmAa78mtBvevKkDNsPx9C9DwhPVym3YjEYbvE1
FkqVgAS7md10OXQAfYMSqRD5xjZq7+W8Ez3HNvd31lljO1Et40PDnH5X0MuH8U2n
cVy7ZIwIznugzaYSZuYZjpDA/9gWtVH6gTW3Z/pKKptfS+gMrqYFjQRKeufZWtlC
Py78/fjXtgAFje4jy3CZh0lWO7gkIFf4GUitMzppCm9WkqRh8dlmDqL/P77vcCDS
vpn5E6XCgXu8FXk9BI8JT4uv6Of+FTBr3b7RUWosDnG4pBQNYZiivGQLg9ACY//a
0Cd9MmPFUNuE2riCJjD3/T5pl08nbRKY95xAcgJfO9xo2uKwU6FHAz0Ahd+UFVHc
98wHlr914CDvRb2X1ywJuaEPK5SyhdTK1b+sV98C3/YtdcLGzX6nlUty4f5UiMUn
0KDqA6PHa6gVLb9Z0r/YWEtcr+uxvkRyKaPFgx4tCI3G3Q87yzvsoPwVoGYLMrcB
7gZtOJysJvkMR/5C9KX7EXDRtcZBhErl5snAWtkgIy6haFQlHCgWAmpdFUPtDLTF
CpeUPmYgZDIkaazV2du7VueSii6IOyzKrCjjSDf+q1vrKq9zipJBXzQmYz+GmntR
3Dei5E7M2/TatQ3RgjrCcFkMRaJk/aZRHEeI9zu3HBZSkUuj5HCBUWPcChgPbKAQ
ZVBniovubKL17C0t+RBFmunURH4rswKVHOSmGCQMyYVt8yNlmdomVX1I3TOhS1s5
AXPGhM+rQn0WLqHvODhfPs1dlRb6rWAiUeKLAWmdX92q1UpcTrebdx9SoXtMIcQn
A/KuouXHEVvMRiSibvLdch9o36UyZfDae7UVQeccKSNBdzOIDSaCtfEV7s2lLF+t
nwSZDwn9tjYIC4Huw4XH58nzTYDu56NaTqvtguMZtx87GqvT8TjH9h0HUcxooXI4
R9I0C5m+NOBGquGuQIJJ3oRnObfu5BZscmafDIwazr7gXx0b2NWQbS2RCQNasMcQ
ohCEMoXQVeh4aDF2TwMpZOB5hzs0jLo3lGcbqlMVQhTMxf9XdqIpRgYtTP+tXCVB
rfQJYitpx7i9u0B7QQNA3q+/R4O/p+IcLTCcgOMYdf/SohRGVc9JEWmBXHNNn4Sj
aHIw61HwAfost+z2ZlnNAlRikWuuIKfE7PJxR7cxZ61Axv8MkmQ16cZ+2SrrlwrX
jerJ2nhBr7CDL9ckMH3sQpSXwgoLzgEYwu3xxHlM5KOdhRqU9CehPVKZYTGnLdP+
6GTTmFONr9/txMJLYbXWK/urmTKz1ceZOu29b8UmH5KuBbYKX6mUeoOEyN724L/G
q5FkL0wx/KamYOwkJtslkpksuvOa0ojW937CXHotggjv1jIe8na0lDr5FghP0Dhc
UTEAbyqijs8VWHYsmvuLAsDokSi0xS1UnzT9pT5lVgKsPwtsMnGkpM1uA4+84Ln/
H5K1ubGi7O0czczA0kLIWUkx1VQZ3/eRRErkMLsIcM1iDhof36/lBM4Zyer5auLz
Mr9DG9q/iVECXgfk2K5nWqMgapWS8Tss9NCmuG831M05J8yedLOtwFK7FH03IDvt
6lRlfvfC5VpmCBluJjVdFycPmrHJrJZo1TzQxe2Riq2S3V7CD5ltniV9MXKAX9kE
tKLIYXO2LwCC8QJjJrNP/CP3eFAmopjDD8sb5S1KLYJhdky/P3NVB2H4e0ewt3qz
cxN9wnIVWJclqrJeBd+t20pVzEUCDsM6/R6S8Djc43U02XjYiV3Tt7IkAsb4P7CA
oFXiCOoHENQvyQKTUWK4IN712AAfGhRa7cDlz9w9Gp9smGq1Y30bkZ1Olxvn8Rug
OFgDKxln81TJ4oln+5SRK0Zsu/7Yo864bFpguvovqnzHb2b5N67jFzDNb/THtlLW
yx29GKziYAXJF7sz67lP3HS9IrCeOXYc9L02/N08yB7iHTlx8TG09XTmiV6BipFb
uJ8eK4Fx5DkbWsUkvFLiWmjCqsdr+tjKJy8UTlPw3ww/k+JsCgX9rlFQEKyx4vAt
qpZuHVLgWYnlu7sfPyc3Fb9zUy/+GIcg2IX2rQSllrItgJ+dN0XWfWCE2oWsxGt6
uLYwJDoeo5l2I2l7veVN0h7meDPXd9oJ50C4bLfQTUlXXxgYqFbW0efVlWLHYVRz
MGhZbEppHUMPauJCW6tff5ROfgvSykoewo4XWZNaFl8g5vBHaR84VvWLjN6uWSa+
dQoy/bUKpov3FFn7I6XfMtxUxccaSKIfTScwuP2h95Kfjqoc/87erVZdDNGeUi/l
s6KWpeqPP5kolr1AeWVZIeJSO5/J1JS8Nw4I5QAAaI3Yg/jm/1rv/SqmJmxPd1XA
pk88ArVSVMMtQwSNAf0XAFwrrka1UsvsfirtNR8BtsoWYLwWLdI7nLqQGuI68n1w
gBfXqz4+0P1LTX101hS43WWvamJR4kYemekFDee0wHwJfbQdo9LRjwq0fqXs9YRa
hJXii9ZgyI3Tww7cdkE1LlSBpQ/xcE44VbCDXOmopqgMDVkX0jKJZ3CuedAbe6C7
H8RRokS0z3NaPUXPUXrI3FtVBGKzTdYFqu2druI2lUwfaFS1y0/mzR4tmC9UKIOd
DsGpJPjifL6TPt1PxIFQKwJDXGF8Y7wY8VnlzAQ6sRUdRJ48eF39qpys93/g+fpD
G92Rpq+AqgoNhrGJYRKFbpXcvEj+K1D4EGPDXjoPUdMnYGbzqp/sRsmVu3hK4JC0
lcpwjgJjnstxSNLqcI/2//rtWX0GlMTuorAArPWGcWkXFnHtk/cLAJINO1ctYqoD
UPBmfYKej/Ys8zAQE0cgMF3LZW+bbl/x7L4siPxuu/tI4VcWS/GEapTH7qqDgu6p
0Ch9kUw/m93Id669ksnJWQ02HvRntMc9KVnRFO7subDkNU9PQB6uVHuG6xSRwTe0
+zq0Y9WqQ0NoB4iSt95W4gmfYzLbzF7+ASGUMdlcFX2M6iFrzHNOnccFHihC6JsS
kK4OhQ4c9c8CX5Hbbcsw9sx9HUvjCbm1IlWYoAMeEWpFdj28I3v9IYOjFoyflbrA
yQoQZvIhmIo0sdCuQQlaUjCegGsfcGXwuuo6H1hM7P94F6xi+hYO/mErTxYaK5Tv
v5lHHDt3aFmIHsY0Q4C4B+6mSyHJlJODZ/9MDGtUvRoWvDbpQFY8Umo6VDqsXisy
+77vZ0TN7BHxMZAaQnsyFr2lyETy/O8yu0fIxJjpuESwJWIFZVgjMYA6S1WPnSzp
SD3yBrIZ6dsJgbozCr/OsOIxyViqrngmQNMlSgnTK7Ky0QkUEB5qlpK5/kMuDR4g
oQfJJN20mnKn9CfZ8/f9LRU6mtH8K9J3U3ev5q/k1hvO6E6WK+PiaDVm7EgXWequ
HleVh9ZZCIQZaWbzlW8RJRGeE/U3CHIcRN5BQVFWYexFz4y1uSLR/8wiixC4wicr
Yt83HTovmLU1dhj71j27XyKlW52Xge9M44TCmFFhDXPoVPfsgkPmOvQX3GhxND1I
u5lUjtwK4bsE8leqM3KTaBupj0LwFuWoix1p+zFkeooPFo4fM1wN0pgsJfus7jql
C0Zjz0ZtEA2NIl0kzqRIQLAe7z1tbTag+8JhN33khCGbjQihmIHmyrscBmChC44s
ZaccJK1SHenkCQ8izm2kAY4u3pzPNcP/QjC7awNISkkI+RS6a51/RFO76k8bN2dF
vp3xXJAZ9aUFTVc5E07gdbmreUdGHVRIVFXS5ZLJ5+hLYnFGMmzeSS6MiSLWyyZs
lNDayA7ILsZY6ng0vXJXwKROz67jOG8e1jQ+GwKEB4qMZJYYOEZLLQJHB8AwI0ka
lo4op2FniwqWjCk/ZAr6jhaajzjUbrx6JONg9540BktMKvj/EG6/pIppsSWoAuYw
iCyFdUWFncUDqFAy91U+jD82CAN2D5K5p0blLgYRt/+8jaXd8VYRDiZ3tP7bsHSH
enbjWhoCYf0FkLG/6saUlVKD241Ucbdp1Nfj46tWksSdtRpj2YgQwMEwGybWEuby
0k6PYcVAQnmtmw3NdDx2N/NAPAFZMsjqLnRklBqBQvwASoxMGUjhRa88wtspXfjE
TcvTx7jHe+0rGYycHNZSmInn5KEjodY04KScFPyKeFb7kFHoQ0G0OZEnNzGC1dKj
krjFN3ajCv5BCsdgAuozsjjQe9eG71CWkgOVyj8ZTVLZ4OXrqDuOlMOepYwAgdd0
BQe0QHxCoxhdVkY53wATCsRu/bTEsgJhDEh8XFRosCMN3JqbAU3inpPSNVbfyinD
R8mUSuIqx4TrNdf2ivPeiitOCF0g0GlkMTk1ya5ww+gGKtxuxHQCeMaUAQseJuKy
P+fIySSVlXWCIRZrAQ8xiD4Y9qwK0odpeXTsGc6f/nJc/3comuCxX/4o916KGpHT
tthWWMTIHTJh0gUAp2RdcEDdyKAfjMydI8If+4DKmaC17bLLfqnQc0XfqvsEzirz
nOhFdKxHkCGfdVX4mJu5oDKL+w6nMEEnvVtJuYEm/IB8+PttfqjV7Iy99hoYsYE0
itSg4YKI8s3Lir5GNS68lX+bz5Pn7X5pBbjW9vTmIK9z24ipD16QxuFIaNd4pyyh
oyN/bELdOeSFyjIBoid2RQ+BYUiAcKf61Z1fTgoT47AYO077hAmD1/GNqSlnkTD9
7wj+wGqZ+wJ9YHeDTNgDddRTpn1enRqm4eqv0Ejod8g0XYe7aVA8UfiOD7+WZagj
UJcBlGsJa/PugUGytq3K90P7E8FlehyRM+af/UK8eacppsAsCrkgoygl25iM51ut
1JMHzMnY5FCBwFbr+puY4d9Y1XLfEOrGvPwYiL8P0f/1M8B6x7h1UPFIFrcsawpa
ndtiDgl98qvBYDBtVqL05EyJCOIzsqiVhYf/Sh0zYnVazHju/wzbm49IXj9EgF+F
y+MXrTx0hc4WElMfuKAvtP3GU84U64WfTHhOkms+s80BVqPm63qX87rK+lBkTVzU
oyWvoyVSpAguglAX+JzLCTJMfSFcsWJgOg5G3kYXvfnfZ5k33ZvlWk/3JInMiku5
oxBNWe/QdhTHqtx4IqMEabTpe8ZrWTSIQXsxjI98yjcjJE0EOaTUZZpgDKxGrryP
lU9H5rw1/2utlHlGWgE1GhYyoj6DQxzEyuov195iD1QhQcKMQSJ307gjMJNWy/Px
JBkmM25wXuFpi6HjUpvCV7L5PGrEulC7n2g3o5scIxAIcbr0FVbtVbiEhHqdwixo
SOX3XQRgBe1g3vFrf64B7LDrFg8PzWn3DmjDz7sFsEQ0rCzZxb0917fONV6GQdOg
kRT54r6m+7nPfwTFncpWWenZgwIGWE/u6n4kqobhEm8t1E0idwfRjrYiwRNeVbX+
eSHUprK6wKF+/JCAmSOzI75DL/wA9ONPM3bZpWU/P4n2V8Y+yKt7vCehM5uYXE4e
gJii0sqqZcKNs39GBhkQ41Jhw6/qchLTn6huTDX4Ine8kDAmQ00gWVY9Joaaci3V
u1VEgEElgyonsfkAsfawAD6GjB7MGtffS+MfqnrChDLPF2e3JggNb9tGXJQZZcLB
IE4YaVsZjFnt51LTmboJmyvlaaoxxEg+vLuxByLXRuoicGsUklYi45SQ3IB8lHfx
JSW90y/tjxwSPtw74fIpOphD69bhdIOIns3fZSc29Nz5zr1RKp+gc2EDMAKSl5eG
nT8yyKCFLNJni21nXJguDp+ZoaPG5JwuQ9el0SLSSDZOuAPtxC5cnFGfjfh3IVWW
1VlrJFAUPG9VVR7rqtTvORD6F2vrNkcyOplMdckxrtCBquebfDz5/jVVrkX+x2ZN
rWnkF21Q83Trmo0Li/L9JUQjE/w7vM2+Dgb3XhggHLLpetg8HA/SKAN4VxCit+q0
hUzO39NliRvv1asN4fWDKKKI1STNfcMNnZbv356GBGPtLS+9HPa4uRHLnz3iu2Gh
4Lgft44NqQSmOQoISQMP2Xmxb2pdgQN0/OOjCcJW9UNysbKVmCUOWP92LUMm//lQ
vZZvdvsu1CzONSz5wgYPM+eDOPSqNeStpPJaWI1BYpyANj03N0Z0l9kD5sMsPYAm
+VbSZOCHAT4h7Kj/4w7zFDTCsi2BwmSijoZVgmO4EgeiFY7GC5EV7EpMdyW/r0Xt
lVuBD/zT6xRebxJyVbfPsEpWoU+kEAl2t5v+tNR8cDtQa8iqvyaJLZDYwWvRMFc1
CrjNNsg2ieZJssLs3Pm1rnmsFpUs3H7UCEv7CwSrbNusXmyTj4UsZO5UxfmMUsYp
NDft6JoL5YXF2dzzqmL4BjZiqI9c/AUd9VLohaeko1S9chDaOXga0S3yB5+f65f9
Pl5UH11/L+ByWLW+hRrRTbQSNKU2G9rBrRs9Gp/7r80CmpvAqrQfOLBdOFUtWV0N
IRUDqOhA6CX8PKkCyYMeU1oC/fVw9Cnj8ChSzmF/uEjqxCZPfpAyebBG+T+zpgTQ
mPPT6r3Qnmom0nPJr2A9khKQeacvB2uqOsDTvCAmnsm7jiuTGYS7M5YezvUebOte
YpyJoYUC4uLk0bTzWe5SZNYU3iwYwMFMQWChyhVZZx9HQK2PKicdG/A54exCIAwm
0ABxHaCMwM1PdsygsxPijBjmCMwd+t4cBRT3zT3sihLvc63eJXD6yFzIiIlUp5Qz
gIu4raNQ3Q85i2/+8sAjSdQvmD884yidMnuUzYd6fW7ylwZGOE2haGiqkI20/K+n
3cKu78j275w9qYd6lKS2c6XqsUP7VGcFUReDTtbdDOBCOK0hkkNSeaIa10EJIPqz
1KrATNrWxdtZ/rAwDx35ohORJLFnOh4WMf5EDTIKrwpr4plUlQEbMHXQ4wSUWV6O
VCHHsjNiVE0TWswp4VcI5vlRBmHi2Qio7W9K1t26bukEIXiibOpCj4/4JEt+FJBb
uhcJx6w/AL31Go4dCzlh/1jQuinLXahXUV3/HCXj+GFb/YLBjJzrPtr514FZs9v9
frzvzxQglwsiaEs4izqngmmFUv1ubAzkAVpwo3rZ/3rts24xN+ftOgOLxTobFLw2
zfiDfAaKerF/jzJTtiTZslJvcNlPvilvQ7kjmZMUumlf3spunlfztvJwJ5EPwORQ
7rG4Nm3ObAOo+MhYaqS+T9CCTtnCbMx7frhLJUAlZj+TNBPjUSfI32hYAYFX4mY6
3HEmZYUqQFHlnItsfXFUS8iYSKXBpCP7DjrlqpnzSkOvMN5J7qmI3roL0si0qaAY
q4cBzSMMB891kt9/7yft3Wxy5BKdx7ukLG1xA9UQsuNNCL2SbIPMk+hJphiPs2MA
pPa84hNS/o0n392oAP0SnkEaY3zFWoxDQ2GSRg6v1FbdugTtipb/I22aUyLBjTbl
8Ci3hrR1TQ96vrkOSY3TBCcVijVseIPMCHDMQZtGNjl+WAz+9WqK/tY/Ja8HtLyQ
vEPltmdmwatL4rqR8kyYrf9AH/bH51YZ1O6ivSHEK7ncj0II317eYzFDltwybgds
1oJGObbAKH1NACzcN5iZ1uRre52Mbev+uLgLU29lBiRqmvQ7HZOE+H+3VqTF/6Xx
qmJWXA+yMv5Lr5yXj6MvrFwVpy6vf/51Mgz/SpAOh5BgdQ0hss/tqvPkGdRMEXjI
Q0IWny8nB26iYiBIcZ04kFPFOFyyFw1SbRU1FBt1Sb/1nm4AuPM2p+yUsdHahHxF
lTGt0p3r9WwbQKpqRAuDZ2VHoHdJF44RykJX8W1M5uYhb1VcSeFk63YD38RGkZni
JOv2nq6zB/buLZjfvSqpkHEt4NKH6nm1MrSQVdu93xnJAM6lx9AeK8/Ov6AOpW9P
xaBAvRc+XzUCj5ARdJDYXeCjnuot71o5/rrE0oD0ZNmvPS1RUkppTBQuZ2vkLbWY
s/0zP8DuY1OECQ2Tt9Xvwgyi0+nypyvwpIzjmTBvVW5V2JKMBhErewFgpzG65OQC
VkOE5k8xyks28l+AJ3ttFX7Iwb9jeJX2uuV+kkTvocDh0WqN8du4Cp8umkN3cOJt
j3PediwtsVcCF6H9Cy080ZtkQaXXiOJFFOGWuDdJNeS9Gc0/VaiIILTZIqcgMq2b
gibKuqhV53ni3lcrtEziwu4uVrIqlRSi0ROvKtEVsfIEHbo3Bo34UpV4EyCq6ufN
CfAka2vcQY/5D00nqUMEZ/b+CYvmCG0N6Z+JoTIMXrm9uq/bUoli2sc3G0wFdIqg
6x4N5gffCWxep5+o659MUwAYnVW7D3oozMy0N/XTn1NPhuBVkoHv3cZ9jRhJTQ//
wt4uApL9Jhxj4+vtmYX1QneoemAkqBBDmkbCforcdlflXDWHUIkcTGM3LxiBTmeC
gwtMWX7SVfFkedgIS8K9/X6pHsdRj6SdU2l1VrtvRmlKyA4H6Zwz8qnFWJCDt+0r
aCA3KMU8t+FqvmxYCZ+1XPId7nUz4HZNpcsME8OPvYW5pit9KpkSiZm8z383fXPl
FzlIm3aya8/thZyui9OfK6h+ijl6hdaNhbhquIjiZ+/qXobwr2gGoIYV8toJJhbJ
cn/5AncUU0iseFOFVvUFTsCARK/ACtbUqpRXe5ObkJJ/hnpDJpZOiC+J/mFnzokW
EhZHRacswkTlrjSJtvQ30tQO5TIgu7nRBLi4rG476hq9b28RbdXToE4WwUZnHloi
PlR989R0ROv1401LSbQsev4ngsmn0832tw579DtpyELMvM6jXR1Niu9sXiCJBmzX
Ko84Lkt/4LHSeO6anQCWnzt/5ieLeOjHsqKTix5mmjQGa6//QCFeUMADXRr5XHon
4kKqGIBxhjfGKsR2u+8wOpXRmorC4oBPDk1cDVZv6Tm5xkllXnjSjyYLXAP9ZSue
fogyvCQJqPrPhqodhHS7N1kHcgqj+3GvIPxl7rdVVdL7m9o6SBLXp8H//DKmfqrX
LOPck5gNLY9a/6sbZwdKeJd9H15IaWpDyPXsk2xOwcDMV0pPktTgFmE+0VDggUjm
FPdTdEhconLWKg9AQw9co8yUnsap5PEYFIzPa202qVwOWcmfhYS6UG6E8vwXHjOQ
rxFRCsWCi3VuwGk4dLu68RoxurUNIFlD2OvMe6DSf6+F6mUL5aICS3NNnVKNPAzC
tF1fCqLiesq/MQcLMDW84XUHnPyfYZWrwTtECavitJEUQF4PCsVfTxPvXzbNkG/J
kg3gMB0qR1TJe1PNq+VXWBaDXE8Gzt5VKPfTX9BJPAvsmZw2WQf8b8lVeNoC4Bs0
rkS7iH4Q6UxnIg/vgth7TseJ4WqAJiLDT0EWqXNVWz1ZIjv9rkWRTKbTvuYLKHIq
KSkWYN68n721Eh4n8OJxm39S4UP55nrSTiNWD8kKo/km/6GxkLHZrsBog72j34RD
rKTxmr6/Bpcvk5Wpf9v78sNO8M5Yk8520HDxgBIKLHlmWtL+M2tQbxSHLhQY4VmH
rGgA6HSqga3XgDeagfZsdvG+JsOSA43rs5qHUnZJdnnpj6n8yrAf77C7Y5jsdiKA
KLuHCB76mtrgyFCBw31OBQQ/rf3TxIRc0gvy9p9NBXaSXGUP+e6Wit+RUAOBjeQ/
vqu8gLQFknDihqhcmH5EUjhkflD9vlXK8BtG4kyz6BIt2RA+hhvPG4O2Mf4SDh1w
4vm+97msHoRDkfB4jgUQCzmQ3f7gkYEpREqWAmqFNsPyXN07d3ZoZQWptn1nPo6O
Or6ITSe1QW8Y8yccPdVbrC1voffvlOEQTSoa9A9GMNBa9vGRH2PeR6fWu1ePxw8p
zB29K3d8Xc/DY0yfthXwUYSMPCpq+Ipx0do/2VdjEIHYFJ+TdbcokPe8N1SZskoB
YTghd/WAnLgu6EwnY1hvuiGnlUmHihoFWdJF2gdJk0bzxKBXYZqs1DeK2MaS0JIe
BtrV95iSZwDOj0AoDvVrldSMllmZHDPYobjuqWhVcpzvkCJB+rPQvNtre0O+3VuE
RNJwlWI+SboWBrbbXT/vkdeAV3ludSWqCnckswJJXp7Jd8IPnmvBMw0NQ7vmUCB5
YjNf8I0bFBMuEhnNvbbEuv/vj3zn5Vxr1kPYf2qxC8BfvSpm27NgYASnWYPQyYWB
SjEgprD+cPsnjFETj1YfoGFtIoxBoe2ENq4vnDO4StNxtUcrdUXEqY21j2fErd8x
rnSn0Af6KNNwOZFw3imqpIp66g7fvAKF9dbCaiD7MHQw3vrmUZXzFybAeWg5nm8o
krJaNirObUkjzhdFvsAzthyWpaJbi71C4s5Z9A3JwpAIVs80bfosi+lcqBxBOzOe
/H8JLJkSbRgbahY8G/CCBHFWzxVQR8X8kHb61FL8js8XbyRHAriPfuYtPw6huWQJ
kaQWcePF1xNYDEtbCylHAdrpazbAcDqK2N0+A5Lyw4Z0V+G8re/Vf+fmYi73nNCz
2mPVMI32tBU7u1lopXAi1XyMyXN0pjZutZLKzKE3Y9euK+sZc0tDVpQusM3ibidI
1IaUOd4o1+IOUCjvmSlf4RJdQ1o8yReC/3y5/iRvYfQDpmz86aHM4ftgCbnKrryj
YMzfb1Kl8UiYlC3WO+VlF+686UD1DNQVyuClR2glq87bGU0N//39Ts7LSLyowLsw
Ed6sX6ppd3B3mINc1hejqI+eaWqxtw4hAVLnh9kfB/tS2XHBpRdSnG0YeVTW467D
Vqy4sJnlOJEMc2gBw9EVKhTDjCQJ4imunxdFEpbT8SaWNe2drA5ZX7QapxOMy+SJ
fxBbmvsHexIB3fkg+IBUtt7cOxXGMHlenAd7ju7zzEJ8uejyOi3XtcpyfcJOh7eq
lEIiggoYDkqxuF3NCZT+qTSVtjH2piJz6NIiDx1qmgIi9aYkErSHR8BmYnfM2+r1
20CMRyPrC3IIOyL3RA8QIL7idesXmXQT1Qs0qJ24dD1opt+sKagCXHJnUA2IHU9P
ts2DyX84YbEmRQuXAk/hvMDKWMKuImHMEz4Dm1gRTZBp85S8x/8BNu909ciqZXMS
hs77o0qVOcE60p5B8vna5RWub6A4yEMO83qAvHmeeeVkGnyjMUeQ8GmFWrEjFAD5
n3YwohtAaIZidRqIT7udlX1fTkD3skHfSIwrhF62uazJx3TfNfMDcIDNu0j/Ji2p
1N1cFgkhDuovXG/V8VOYciMsdlqTHeRpt84GN4wN+xM/m+BgQ15mrOC0akcs8X4d
HRr0otjq8VKORYfN+v52kClrEEOuYzb3OLNPcfOd6y2HhFzu5mU3CyS933l9dyxT
P6vwaEZU4kH4cNYdUn4on8FSguUrZqRluH96IQ6Bxoevxfh/OzRqysyLziTpdlyg
xSQwnpcFWuO6eWrRCKtA3d8OXRp1TLq2651mhZSfDxpwtgyIpuSzLZ9aObHxnQnq
Q19FEWqyPTcbV7cMoNm7mfa5KIM7SHhkGZdmaYChtrNh+DWlrXAK1kJJm8RF9Mf1
POnLXi0009hywjROSTDUwJvZ4Zt8uPsOtUlxwBhleV8hIMOquRhRzT6LPVH5LGp8
OddxEWKdMxp7twGDJ8gJdaa3ILIm4ZCN//7RuiKd5NAQT0M+CD1XYW+qM96E6jIh
ODsWARLPNgaPPdX4hTe0MLTAb9pSX6Tfb+NwRufT0r+jLJ/2sJv3KqsieD7z2lr7
VZ8PPnYYoZDBXDd2kknSZfXq+6BWajq5rA96JocQaYO8HBZvON4C3fcTW3Ft8zEt
/gbv49nN5vCTO9UDi5VEqjhB0Md6G2c7LfKVSpqkBWstiOY4567u89+VYg66wpQJ
L4RZ6rdk7xYESIlvFp0VELPBqUrwRIaLsywprffJrfx6crN3DGY3xIZ5AUPuxmX7
fgJuMiOwoiSyRDs3FNGbL5t0cSk6OxxdZMmtJPMm6foDUBtb71ximPKsDNMwBKti
mYWGez+YwdPlxfJoW7VCGR2MPil++0BqSbls5brpxPp6+SNZqLsQcIbrdc+GV3PJ
IVk5JsZGG1iB7kxtghr5nh1dzcRDGlcXk5q8zzU6n4YLHlMF28qvj8l6Xv1yrvwm
h08mg6GYMzqKptHLiVOla5wZ34VDRza9UfFVl0w5AnkDY8VGjH5g7hdZez0ld8vr
J5YH5GB/85VmafL/0CEJ0h3F+ZTdF8Zsfq/74hfnd0jOKDRCBVN7BLIeQYtvjFq4
jP+twhqOWVF2xYzIZ6QkRRlYGGb6D/Et7svxEFA977BdV4f5d45aJncV2WsLgIGF
tZ2+QGZCoc2n81AbJt7kFINtQMqsyV2R8O+QgJJi+HlFSaFbsvBUASd98iJQSOLh
uAa+riWZ1Lqu/jLHR6IzHfHzsvvV9uJ8aMQ9GdjriHIpQaALllaUtH+CVbWe8m58
YC2xpdCTpSi8IIXv9+VV2tuwfgHLnZtk7h3Yc/D6kiUzEGrA10ZwLgVCPiObiA6Q
bazUTupYNwLCV7hrMLGvDg/XVUdGg3HgLxMEOv3XqRLbJ+85HZoYv7/f980LtzWT
Qu13jAhAk6J8f+p5hDSLa2JUhgB2umJPnCYyFnU2pjW+vWDncA66ZcqYM5C38e1+
bQ2Q1Y51OxpM4mtyiZr3hguJgjPN24yqA1IECnp1oNqKlKpFvHo6izJl7Euiw84i
9uOGgrzcWe5eq7lD9BVPGFIEbvW0GZeDekEI2Usa295OfxNi6gnBQFfxXPL5w5Th
zWac1TXThVQ3Wt8HVzutp+NPepR5Obb5VotD+HXIkIeJ6r57pGYxghEXshKjGed0
OEgMDOJAH3FZPf06g8qUnPRyQ21odgpz7aOtQ1m9yYT1UEs2nBxllUvzz0fa0rgx
Kh20zEWMYm2Xmx5LUyeWt5oJOPGIxW/GQlDFNNgg/42bRB10orBD1GjYhmFrsQgS
IwNu0JRcKtvan82UhO5lebm5jERO+rVJ0poSAaZyZ24nGeQXf+iBcftFURwIUmsn
AK1rTdCdCj+epDoTBy8RWkOOxnyVQJop7Q2cOpMW/3wXAWq6c7AioArb72evNpZ9
EP+7QBzZQnGeBnbkl97Q/m9ucyPNoYnmHoa+ERL9og3SILjJsk+OLv11uiZcfVO7
MHxDaPWj1HHpQ5wsRCQ3X04dehnCfckRoX2PEUnJJslxo3V9zIDvIuEV2WPxfJcv
nPAlJLKNW5KRDMhkVd7LFJ2gZcmT9jO3MiDxex4cEamxMwT/cC0vi5GfVHpqzU8i
RQLbklXR63iiLtQviE9+Yo3x5GGlt8HlcoF9NfjttmAVZuccSJdspJ7GpK1fchv/
L+CY4JZXjwbz6fYwC3jjFp8Y2zxKOeoHIviZKQhWx3CzSwy2KM4sCa5cxAGUVOC+
rciVuKsfXDtQ3rhPQ0bFGpfPeEEUzUvU4DaGYofJ+mLeqxf5hrDQFRG3w5Tkj+Fo
WKT6aNZkDj/kIRxWQ2+vwJxOooSZBJKemfg/edIOTu32l5cnUrFwOoirowuapwHT
8lG6c4fggqtbCcpGJXlnVbx/qP0lJNN8/Pxk7CpO+03UsAdgDduG6gcYiiBf1bsK
LGEmsnPtaD1stHGr2xUMeE0K4LR4RTwehMXOSP0OIIsmawfGggQYF3PLli75d3AO
foue0nfp6ifJlrAH7AWxK+RGnvR6vuXpjmwU/Lf9tC7b1TTLT39xmvnYoeDM+6MI
2I2hVTJeoJeOF/PY9lJNF5DtwvdmX6lP3Nj2+ykPAlz8TAYahZuBt2UIf7+ojNM4
Fhko+6fpqI+IhgtGqmtFG/qjYvn5WTqZy6Q3DD4xHfhxiZCxLpBM/1CYXqEY4Bfy
TfsUYpSF9ed/PR02wT3NgdZQxz5vtm+e3RM8VmJlq0QHElIJMaRXPWSSbw3ywPOb
l42BLvWZ4/lOh7WmVstk2Y/MR0wgZeG7UHbyRhvsyaasBBqSd5pB06xZmslHdycq
Wwu6AVxk1r9du3yw8BeN9RjnfrqvNkuLLqH9D5nvv8DBW4vXK0mDYoCAKOPFAiir
8Qmwu+ecuG05zfi+0JFiKMeCMtM6m1a+zPLEUqP74mdeuJVkYgBuSY1E7mMvYzZ9
9+R3YjldxLCW4qIbr5SNoDglv54kMEKrNmjUyncI693fdYKXGD2bid2rInm2VIpw
L69u5dK58x2v529EOwLMY5sJzYeWHlUPsICSAalKKhMvZyefk1c5+Gv6BkYOdfiR
ApfXVgp/aIWgXFM1+1drdWaeWNoivulg41LhhwEYp3yYQeRIaergQlZuVGU6A2Zb
p8gFyEq+egzCCWmx84dfu90CUV6J1xgpzH2Awg/sjL/FO1tiPdgeSeFUhZS0Yy6u
5UVv2HjsFbXd+KRZHlV+7g6xnTL6W298HpK/+t4jpAx96BvzXJ6ic1Hn+cSn+rLg
5VWTJVYVnmzpb/UDkWlWcok9Pa13M1z85PittqiAVHK1I/H/C5TUEMp6DXnAhm7j
v8nqonoXZdKDfd2NOtRiqL3PiKCAmqZqV10IBH0po8C4KEF5Iq6sbVwZ8FBGRrTm
ckG8QSZpGS1Rp8RikWFeVvyaW0Vqr4hHEszgjpFRNKWCw2+KGJK3MRBWmoxFgYbF
b6UIgPMss50fU9CHle3UtPtWPLwU4UCNr+5ln58eGnRaLWwtel7Qww1tnhsvbzqf
VQYEALpAlDLpuGodEAYLMGbL1Ho+ETzSStbpbxHTa8ccEiptW9scWRxsMlX0rqY/
Lb5nuEB6bn6el1lMNxqGndkwdVaFHB+rAjdWgmVpEozspsbHd9JpYOLFIZ+RDog/
0B+g2VFDWEZOC2ZMtcO87YTBm9ihX//cSetfyoVyHmYZyKqctHKSpns4Z9NxX7ji
fXZQxcoWlhY5RzJa3EWUgC3F5PidDe0xNSw7Tf9ozaoGfNh4DIF61iF6ZcCTd0Yo
wdeXMZOy2VlPZ5M2aRHhtVIqu6uYQ6XxPiEiTAa1p+B8t3CzlsSe3euLDMzzH98V
tpBrZUYgT6wgWV0ifmoSuo0ZzjoDgSneHJ5uMkihfJWxjh7DCXGq/gKGBXUmOQqi
kAc5IWHqmzuTGH7sJBE26Hb4f45BKJoFVHyF2lVnrcDnQAaDN9Gm0BUO8KI3iYVl
QtnNBCkytF93C4d6ruvylDNAgZsbaJ8BEX9H1TB5rfLveq9Rpn4aDJ62pRoTH6ea
87tyIgdjvFit97/FhFgHXwsUw6V//58m6++pXv2oKcphzfnYsEzIc9v75JMZKyaG
c5kYhwPYWkXpnS5AL4KParf36bXM94lK6S3rS8Fhg5KKgPN73IwmJ99GzOI12N1I
7MXxridmuf21owq2p2/Stt1aoI17Rl5bUZsCHIGB26S+TriSQ+lFeEN4Ea/UjPWd
TlBLF484e+oUqoQ6JZKuiy8YGsV3EakM2C8KcPpmZNXRAzctlBoHtSzXV5lZRF9r
AOk8T2xNaQU539wGF22fqA3N3136m35Fs6zUGkkyFnraLIrnZHSGw3CqKDEH2q+l
2Eo7pBw79S1rNi0ddl+k+TWTQOw53MwwQfqucrFBwqe/O7u5nf1xzI+lFAkoduYz
F9ODsqFudzoBrc3FPWEstQFbpSKvxK+4qN//I+mLTL2Kftu0eBgvbRcnTExq5CqS
1fTT8rwljj00hw6y59CcuE6ZUn+ztcSiokn/ZA8ks6fAUgns2tP7moIzBIplgY5/
WCKg4t8/M1pzoIRGFMBi7W8PCupK6aOlwPaBizeBAq+H98rOgDFYLBOQfVmggYyN
/KhI0iCGcwOzAPI4UHbfqL7I86bznUcS+BA0AtSk7VI1v2CmQw3MC9MboG8irkry
yBuosHRZ7VyYszTsC6xTWNf7BdsCIymqMAPZfb0AM8vtVwoVeD/r7te2t+tvYOWV
s+8fqXjus+KSTXPutP2m8tpgHOBanwhMCw5brnaMpMmsrIevf2SpruqHliItzA82
gPT56phPq1F8vGmxdEQ5RYAKHdHV8sPS9mukNNV1gl3cXtXY+MhzvBpFpSRsuJoZ
xxjMYmkU1s0Zv51SG1wHiLFh3FdT+Ce8yDGAEv/y3UWU0HnNBiyqIFCWy8Ko2gvz
uY0vO14BeGYT5Rx3Uw5tUojR3lHi86/PuzbBWtK1ivvvkSQa3UPLAM9+eznNeaTg
xRKCWj9QVnhpy4p+RBf0qGBCL/JZNDr+xIsunW76lVtDfkp7eM0GZi3TiscqIq+t
CLNaFgb2VOrdTPpumAHqTsYuZs7MWmpxuw2xZeVuh64ja2V5Dey3RBuTa7QtkXCr
pOvTxAC+LjdvpBA5FNe9AHMK3GCusbbGlBJ1yvYNDEtIjvjRuoUDmDjtSsQLt64b
yOy/EI4C7ftHin5W1PTxWFkxRgnJdcEN6cCUFrwQvTKIWqAdI1F7gxq30lwuULKD
hvzVQTnrFhX8CX+8obfzTXbK3FXJH06LdlsI4lxRN54BGvtSm1gWhMCIZxbxQ0Ga
JPS9XCiCZ8HXlacOyXpO7cElGSW8hlp4vgeVofH8Bxd4EhP9U6P94CP+npbFZqXH
iS9ijDDzjy8whTp/9lR0P4jmidV0G0JgQ1p4pfMIxd3VRpafF83NaeX33M6c/D07
dVYoi6Z7lYVVtg9fIzrnGd19LeeJQHLd+ya0aye1y/vAMcDWvTWM4Voozenm7shf
kEGaiGEIBh8qINrPMsClM8GH2WDtCY7DR5wmX/yBHtZdsE9ZB30IxBDy3b4+wigs
s//J6wAtamZ2Occ0PgHI26M21Z4KtWs1kvH77G4Rq4DNV52ihCFUa1m4wfpFOpVk
eJrDgFrXxInkXv4zBfeDCKAibINHtL4d5wBkdytdd2MTRwrIuF1Kc6pqFAQgz7fp
Y8gVh/6XTP9dm9bbnSfgqEuL6JEjlGZytTnq7yS4fbLOrYm5Vnamhgw7d0Bq7sWM
EXO4vGKNgqs4GxjRjrvTPww4XTktYkue5paBoO7TDiwMrY0YnLgZqSHbBMtJk6uY
cDtCGIcdB1pfRYJliCvCRekRNc0uzhMQEtC5GcvJSKJkKcft4UecH60Cxik126gk
YndFUALeD4kGBZ7FRrfODA1v2gopnKaPHAuqQ1SXDBls6TwxFS68m1m/FCQhICCl
ghPCgkQCvCfN+XtfsPm7LBKM26KP4P195KiwIOjqvYqvVIb34clP07pmbifCZ472
JFd7ArlawCLDsPRFeIWqEA2zb6m9thLjU7p9Hr6ZxYwUGa5zpYQSRDKysl5PtIGi
LFkECf+RpQwKjWE870Zxd+LrLU65nN45XFhVfoy8eo4I7pKQhjQITGwQElm4T1zg
/23V/dxRdaLVWGfj7/tq4F8MsXAnuOp7CJ5sQ2Sjw3dkfcAw7k9aiLyHg6iwbjyo
3XSspsJuMPFwtKZk/1rU8PzHVeZk025DfWkI5UykeGoqx0fOhSsp/3IXOnCwvwPj
b05US0bjDGZGtzMFY/zNN1p4Ab+TurVRaNmh03zE714FiUWhUczEgGnsGBegn53C
fGM12s0DH4hb0rBvmD6SLimPG0lwApmBA2rq78vpe2j5Zh0SJbAzmFTng06SBndd
1UXqYRN7fRLo/sCFINN0oBevCsGe6vTwGZHKFIRRpRguHntSNwUVuEZE6yJnuik2
S8IvxlAPhQJ/7VucAf8Kplm9Mi6IeZxhhdn1nrhy2EEvuePjnORi200Sy+zTfwet
2KzMsD2CpmEzJDQLn/IV6bvWUHdjN89+VkuWDE4cNMRx7K52PXxBASuDxyvfbwBo
CDC9uFUFrwNV+QTa1K+Go17Ruet7fvdt/YHd3mlC/hJUGx0DzXrzk2wPr97incjN
R3sOSpMNVWIoGllY9ZXT6mybPI36+jTpB5Xwgu7pG1zS7x7fHFZYUjRDudmMXuHN
OVe1C47lOL5on7ZBPAwfMcEJD6ADteyhB8dzvpv6S4fIgGE55OeImuP4qp6hNYkF
AEPWsKYENPOCLDMh6VwmHPhAPn+qcg+YqiTZrQheYm8rKkHSD/cBNENFaCexVrd0
yKoWgYz9jA0V7W13QAu+0Q3wGe4Ysi+Tw9bvRUh+sSx0k9zSdvEqON0CIgCoBrvJ
xrGiL68DkZ61WtjNeUz5qbqVue50lqj4VZXBu1KKfgYSmJEsKDzrLfmAE2hSIh4b
b43HegZhS7cRCjqnkdxExQ9aHjAI7BWPxpsPKM5CUvc+Qxh/UBq1pf5Z/CSFSdxv
D4lEUTl0z5u9tpLBtlcriGHnfkjOF0wNYMQu4U6dt5AkrM+HK4xJKg3nqoMiohNm
I3V7Zu2rTS5fbi3kdbj+QpcfocRJ+aMwLLdoG1e2G2cSLqR3X8EEwONFaycPp2vR
MPaenIEz1UcC/qxbKLK6/nVP1EOWs+XEiATEi6PzNnBaIrGQrPVRm0xWOGPxXq8O
IypgTcM3hG7FWen2EQw8G4BxtNTo9nT+WiQKq59ZoVSzPLeKdaf5P3eLt48MJR0z
48qhpF0DoorfJyK0IgNuEBM7CWue1lXVdQocHkc4dn8e088liHNf3dWCsSyLUQuG
/NPkhQnQ2YTMrfWPGw5VXSNdjIVn8E+Vp0lWHoOT7/Xiig8KTxhV6kS8VflMr2yd
onS60y3Oo+U3wEOvnMt5dnBj4tex4L++EaaHsH6GuEO0sH77Aj+buO4Y2FRwCoUz
7B6BKaBtog0GXcz/PX+4cmANkcEs6/bUAnwj8g/l5WeiA7VGkiLuE2MFkVfADbrk
0IfJ3Wz1jPdXsaIef5jUp4aJq2Ltb/G+eOsujv/BqcFKfot1qzQH9e5pCGdSj6lM
o1D9kig7tkA6Kp8EFUKW3QACoSexbsESTVYLH7to8kQ664SqppLKuY/PAr51iEvk
AKoT2e6kohOl/ZtRVTL1+V0p5BAaipWFFlU4sqOvAV4Oi4cbj+FtI/vpXhZog+a2
K0hR+K5e3GEqLIjP5AqQmbZvgvp5MO2IKlkSbC5IA7lUUPhchMpNj0ONH+bYSYHm
B2PxGvk+ZLUbdwcyZo8KR2UIhgf62EvcFyFOifh5espna6ry6LKoA/fokbplixWY
gIRKPsuLw+7KAPbY8pPptySC17LnDG6Wal5Bkm3Lxxs7kJVcCjfnQh8EOtWFn04H
43TIxtTZ8gZpC5ytHyUBBClQDFMCV+m7lFNpUD1C3Uq5GhzMX+2G8NUqeeKPJLjS
wfSLGu5AxeHgXvErof3SEOB7frMjk9zLArNcqOYCcgQzTGq0OhFJznkfQznOkB/W
QKEcjSbuTDqwGADw9DrnVxoz9zC96BElTCHBg/UIaSamcf86er2ecpx+SFQW7x4P
VvGSCYQi84V2WR60A/fB+qiZmGnA9/ZVrdA3uh1v2qr2058kj+MS01+XGCbpQ1J/
7fRY0PHTfeGMPZ9IdzbWnqgAFBOyd8yA2QMOe+LENjsEKndyNFfexpPyf8tWQr88
JQAeR0YoRLPFM+f5eDv3wGrpumK+z1yGm9hFlbQtlMFyR5R7/0kGcwlgeKlRoK87
BL9grY4nalxMZMg7pCWkyWHgLgdxNTfTjWMErsWTs+ff/dlBymQmgCc8bg1h0nK+
Ohpfe8EFccN4lXQgNu3sO52RJ15Zt64flFkr25Do7PB7yKgUiWTPmslNnZQzSWou
OI+I4r0x2e/PuG8vJIEAktMIcAB9yf0+ZENq6Hy0dZ0L74J7bS7OHmGxYYbC31e6
DithCp3l1IncGjLYbd3VRLRmi/f7Czwz5Nrg1ecb68VtMWhciM9u2+WpKSZDv9BD
CSTi8BCtAFyUvVa119ovpnPHwRrhheqk4cH6VmsmAnlylnA6fedYunoHpckh3pPq
DUAp07NUvUz2cpbZhnDQgDrt7cu10ZJgSsNHI6gi4FIDFu9C0pCM0YcXGLXXYv7N
1l2gxRtPdtIl8hgGwmiZ9yu4qYkrb0/UrbH8EArZPItYy9d/ORApdvZK+OSg06ap
rBFXrtfz99I15/jgdMJO+0E6GBmspz6j2HfsArbVAhd8aHTRiLlLfhXLDTUnR8FU
grtM+XeZoSkHcZBert9BHySIVPCfWFfr4mcQc0e0gnrhgAkXT0q/QxKZ0rP7aWm9
2/JdgN0Hy0lybwTGFZg1GyGX/JS3gp5rM7cZQNqe3z8LEneBHC+HFFsGxn570HVx
pVPd+nZEd96HzeQrtrh+a/w/CRFgtLZLmIhovyv7gDbpNH3TjULUn/VA9cnEcg0J
ZoWiyb55vdGrSogpy8EvH2Q5jJB9cUzGveZ+TV8HdeWP/w7mvwCvGdSfi18WfHBL
xTLBiyTT4weFDI5urzjFT4ZrH2VeY7mzmi1mi8gNxazngYWLvmKjYGR1aq4HANk/
4BtRGrVKZ1ZSoK6ORIa3Iv4fmJ9RoXZaoR/9VDEVn+k1ND3G8PU1ZkVI0vhs2SWT
UxK0S1scg1Xb9glqMnJOvE421eRnj5oqnDQMARQvQNqYpRMkrzPr9UJigtm5f/fW
RZWVmdW12uaKA1mZp8bfg67aruYQWXLcuKC3/H7r5noqcdoV/z6+P+4zVm2I1sDY
buobu0MBNFthMuWSAaiej6OvtLpcgtf2M1MO6DqnXr8PQIm4PGyswFDE5DaQXgoe
P/E+54YTg2KLmQQ28Zv6ljwxnuIdvBDDIKiShM2oTJy4SFtJZyQ356/dhtA8qIXs
mXHxaDs7Sl1EzMA39uI/DCN2u0Ab0KLbLZ1YX6RvyGJVaJHl/DKPDeGl3CBiK5il
aHGDMFj463eNxvWu1c/TXEeAJxLiROTHSnilYbtL0WL/rlVABXiP8dh2f1P/aiXY
je2D+0BdBWWNpgs8Dfndaezv6fGyAKOnH90vicNXGh+4kMc5fVuPZcP9idgLYY5G
yUf1UHbQks6yTfnN3vqHsMEAUqVc467dvoMdJwISzY3HHy//iluf/pfKqOLtokv1
XJgdUH9eza6KJFtGJUBSQ2C++c1cXMZZ7rNzLPL3WGUZnbyotAdhnQMMjP+CGjJ3
eLf668X4odb4TfMmN9LK6uvHRjiPVVvwqGifoI5zZnnvnNw7TU6kJr7rV2pBWQtq
VgqrK+vT4d2akAuejhkDgTc1j4QOdjnNTQSyt0qHN7ZkVipfOzj3ZrPytwYukjlS
FoJDy5+iQ7zVjcQaUqlQS5KK97yKrMfD9r1ndWC3A5w1UoS9Kn4A15UUtBulAFER
mEqLBAG9KSfDI+pdiTrlj43l3GXTIstL22ZtwxX7RN5jJR5Acgvpb6n1TPmUsYfL
09TeWQHXESKFLMlyXDA/blW6uPUtBFUaJ+D07/d2kmqPNC/A0A7gJ68+fpbpph27
o/Ooh5f90FYCLVoIklOEirw0P6MK5ql9G97EpVEIZUShztH+1jqORRYZlkUF+kGI
CfF9BMGX2Voherso9cKO6FbO7anUPz68o/2RcGKl27mN9MeD68s23k/BRzspx0Uc
fXfi9EQ2kNq5A2OIChfyU00OCtTrJ22WSkYEGxD3PlTod9nTMnHfzwIAhopk1g/q
0aGZnbuiwMvy6W5mNXXK+jCf2111EdF5IGWEJJ4Lc9eZoRLsrXmIYvkmJWs4JCV1
qCfE7vfEcknJMmh/+7K+rcjFiqsej8GXPAoggexroi9Vg6X5ZsUYKizFf7/+j7OJ
Haaf43zDibdMBQYg5DWNK7qDfkNcJm8K/mJh/ZoSI5N7wZ+P0G9MmOkJYL7ChLZJ
z4/F9T8gaMJQJS4fzl/c2fQG0x7+ji5pho9UGCSEwwjRVKsU9fLhsY6Gn8bWgYnW
J6owo/VcxQr7jY3zcO7W/1ZN8Jc6ob48e/JiB4EFpuuohK6piVMPN6UA4n27px5A
DCgp0CX7HC0JNk5WY8gCrN1suPo/gFRCqNCGG41szZbv3qpX5FsG/5ZY0tzX1rnC
Kl/9YW8+N3NnhV5EllbqATx1Bd6bMpLOqSRalHqDQ2bYxhuS/pIr/0+pxtuA6MxA
Ziq0ZDRMk783bMRSoerJOBPt23ntvL0wM09gbYB4yCyEx5coDuZstimggN++jN0F
MXJzr+4qcoJUnvraOHl8P0m+bn4eGjfh2wMUY5Ik5fITVy1KBAEmc1yyLSymS0EX
CZxEIeECAKaL8OdvvN/jyMLmItkhJHJCeF2BNKMBGIRpNmzWGYPq2Tu7YVsweJWK
L4GBdxvjXNwJjhlSFX7F96j5YHLO5TgRGas7YUn8yM1DNvgsf6i6akCxLENSIlOm
sX7kybMrPxYuDzAA/a9+zZ2XTuMkWzq5C0H/qFEWzTJRl0klWlSXDtE9dIxSWd+N
5poUbHA/4bKffkA3zAy1ZhMvf+2U68tsOlGHMtbpbyN5s37QlAmprPcRWr14D7eW
Lg27/fLOm8sk8ziF5ZC0UnaRvfftJt961k7UxaKx4UvQL8AZjcF8hs+G0gwKt5og
+0mlCj5VjLW+8oE+soHRNB5MF8yv0YB2YA0fzJvw1oyI+ck6qAbfaU9BKj4BLgKx
NOa7IiUQ7eQf8oD4Z+U7MH97Cch1n5r62n0NcdjhOlU6TZEsffj3wO77tsFCRZJD
V/p5WnK/2Eiy+jPdLxHKlK/IrWmV7sSYwWPylYJL/0EsumlADTWKASjvKsRpJmQI
db9ea2naFXWPhRqL5w7r2AGTb0cBUWPb7E7KOprjEtDOCY39knaGnyYT5PzLbMBn
kMWRaU69yimJh0u6ss37/IbfAUfyYOoj9SCibeBVKrrgIWXGIGgBMTtvtvF3AGCs
cKtncSDQG/56lZXqJTfFlEmuHEe2PIEx5mrXvgORe2XRAYOrn9j4aZ2YEwIBJdf6
EWbn4h+yfoJT1e2sVTh8TM7ohb3pqYEIksV3KAGBEVtWSY6pPGdIXTEinN9GWVGr
Ge6MjEmLpwB9CKZEZ/fHbIiAVoFHOSbv7YIiY32N/GsQOIXUwj/zT4QjOgXOSiaA
dQsCm3XvxbrIRvJktrNG6avW/nqWuBNTbot+oS99AoQNAYAQwDAm1GcgGtMiQ+l5
xoCeyd7IwpYTzPOJCOI8ozSy5A2BH9GAPGNKAQhD2/5i0ohw9ehmbcItjaeCt05o
ilWzgiPVCZ5F4bgilf6cTgRPXdGa5wWT/ZcUVs49ngfS071zmCQWgu/z/JHJxp0d
EHTh4sX1yVOwBjnpGvoONThDU4MgfOrXaLSpRuD5dVbZUpZMN0XqvcYeSyu2+oJk
93rShaBkqKtnzWrmsCdRxvSbj69cGh7XuSkwKvjTjpKOCQlwIJmtFf32ZU1uFrwj
LcUXuxlPpD0zoh7NXzjg1HoufTlKJpdqFjTqIot6dkE3Afcmo/E30ZG5kmGMU7lF
xXeIzmhDAypl8rpjW9oOTfERKxeq6hgrIUejaxbsKNktrgQ+rHNuiSDnnWGmv8QB
RYq+xLfGGQ5igd5UJIhsBGQxTKujA+GNYAMMxpYhAeT8B6M3tvIPcdfLQUbfINM7
iDOWZfrTQ2D3O0DLRsOsyjX+0YfN5bMfz43x7lwTAXc75Suf6+U6m1KJoBXxUfDZ
i0mRBsjwapm3YmyzCFTZDz8KNeCF2z1ZW/RZjIbM3NabOHezH3/zHaDvADHMYdrY
gS7FegvJM1q6Zew87JnRPIwvXeo2A+Vq75ncdB2p4H/PZf72uUT6t97DpmwmVJON
Wzulzat6ZEuCauCPRQTC2OwJGeViBonmURXpkGWMI394u7QdvC7Gnfu9mgHNEbTJ
xqMivZYV47MBiHi531XhZZqlScOV1oRSUYOdV4l2jtU24YHAA+LqBBXAKlVtC4JC
U4w7z0ToVICfITWCQZCLBSLCxLfgxNu5Lh2yK0cdz4FuMirigy0PkPtogzM8H307
XXqtGGnYEo6o/0+O4+0J49koMJHOBZWOX0PhfobKkqt01+U9tZI7MMTHSHhK1C7G
+Utt4FceqoF/FNSr0B5fXcxDwYIPHE4zgmu5FksS0h09BxUyriznZ7coaqr/k2de
ZmBzgxGOhDWlSZtMouafPnEoI3Nw4FjJr56o+nnUv1b3wL1jim4V/rjL0pfO/Mmg
RN5uzrrb8Kvy3HEsB07wJN8r7r60bQQQKjqKjr3bz14tfTECy6V9IPHE0NSqfUPo
/Mjc2Dc2jgSbQtRvNS4YEvrYkXd6TvOWP3kaM0tD387C//QDAPjAtH8pm7ikSgG8
wc/2RA4zvwj5GGAs/Ovl3IvokBYAZbAdj3P8JUAEzQteglSQ3oNP7NTkruc8Bhvi
oQ25MnNxEF0gtETLIyRprFRZgAq7R4f+CX4fzQNppp/tEdzLogYrAwAlsWVW1oK5
UMU14y7g4MWUYPXjaxsDSfF3EUZ8K0HqeHKePGJJTx3jWGO4En3OVwrSYazsUZJg
58Wtd3azOU661y4/F3hAzta3YkQtfGKcozS2narXTop6qgNSVr9XDkXmPeDdyEHW
Y40Nt7eVWDvySpFtCcOlme+EziVwwvBX/+/IYfv2f/Qb2naY3wF/lk8QoMXriwZy
9SEdcn6GKY09qxXeWADMjDrWRC8sSipzP80nOdv0BXsFittxfKcDH3WhK+ZJj0+O
93QxowpkIqSDYf+wVuvuxKN2z2sDXJl2bPfOnzqzsu2NaTRvATCPvLdTr3jAHW1I
fxQ0yl4TsVoi//mR0qIRRHXRq2ryq7yznRs3bKeFGccMWEw8qQbLADMnqc1RPhXi
kBN+mP7icQv5h9QbAjg1iYQMDQHPBoaOLnjbHI2gS0pHHz93vAtR2p4I5hXRkHxX
l6i1cRN9qNdgg7a53Psu1OHSQj5Uk+fk+RsC8nqiKWi/FSD6unVLoMyL8pzZ8l1z
Lwxx7vQS/unfksUNFevdqOGn2YY3JMMKJwHJGJ7aeFjpCUr/JZo1ND0Rxeb2srnA
I8xD3IQiTgmpakV8x2Wy+7Mat8l7U4oSEAzhAopKcUs2v6XRWC925fnJI4NuuO32
GHzrKtiAIYb3E4yxQPn0Sz8B1Ugium8Y9ewLpvNNhUzfCN+3ddAR1ifRe6Am8U6y
8GvZjq9SK3MtkUdRppXD20sfk/4yw9rTgq3SJYSupFnFMYuSL3jlgJV2H1atguy1
gVP0Q0cBvjXE21hytp5lDVvxGOp/cq/hgTY383bDLi3X4A/epIAql/SCfuC8yFIo
RcaJyamw2Rj9ywIyTUN3xBxJJ0JY2+tvlGYa5UNr/lPdZ9vf+QPUgqSY9zgDt7Au
ZeRrTW5irOCamuH/RvXE6iOg1Y6Nl5WbH16DWN1ixYSS8SHcCyAdBTbEscDpMcgs
3EUfg+yPMNKEK7IqUQNw2Jt/RnP8p0knWEFnuxJMcXdUwB585yer2lSnT+T6YSIf
rpcw023wtHVRjzZnqU3H8aUFieEE3rDPk6i+XoLdcMqp/KCsBjCYs1cV3UZa0RDU
gSQccNNHdCmNVrEQidQ9iqjdBi3tAkllDubYObCJeh4WYN+169MxUpZEg2ntirVe
OqBnq5kJfYnzEOpced2Y3S/fDS+Td3FpbDaZgqY/2tYLD/nFSGJZMCvZNkNz63J9
EFxpVjyjiH+pLhEJgDD67FhVGtOvgE3hUmrXFpfWfChqTXOpu80h/UoxLAgFqtci
PtMiy/C+xMwC8g0smotzPKNw3EFU7hj7iJUXYy9vy4Ky9asnhFB1FB4UR3TSeL66
g838oNv9s6GLEr6bHkP27liI+pqlIHzZTzG2uMMhxsc3RTn5Hv0RHOt3FmkxXlEs
tE/VnBqUinNxmpe75Jnf0E7lioGQyppbLIdRzPK1XzF7bfUcddi8zeKOUV5aK3Rs
3IQB6Iwcomvy53A1y7OcsFY65A5J8x2HbJBAlbAT3UdAMatnLWazuYY+qOTpzVPL
ZoxeGnrCS+FyvgubpFy3J2lW75NZWTW/7caDQT5YjgckrKEE/WCQrrJZc00Cwq1P
mhBvPacba6XPk1ruL5xgbhHtJO2rQNJOAl1Siu+4pY6B5gFv7JkwOyHO7+70EX3m
6KGjTp7rEfmv+eUeOFBUK9Gg3dVLD7uBD5J9YhD+svfv+gyCqYYUSD+p4tfAM3kh
k378uLbj+fIDUmj0nMNhzuGjTK2oyYbBt4KmIKTO9oYVgxx7mUS6/OkgpPInmQUh
8I2em9xf0lBtei4CTUPFwpClShkF4EsVTHX2alGAEYna2hmpkMGA5yHJJU8nGOsT
hPgev82rqFAuJOb2jgb25fGTbUeVyhzIXRXwYDpa9h6QrzLZP7SoCnUXXqd9j/St
1CSg90Hw7mM8Ot/54CbDiQw5ARFgmaFS/jt+33vH48wNRlxBl0f9PlwdeDyA+J8H
CJJdEvENrucMNMbksOCo84vomNvDMijnNFsfbPx/M+VM2RFDQRp/7G9uTdnQuSdf
mjoff1mRMy9BZ48eOazrhQRAI0npXY/FcHnodScaN79xT+8DxO0WylefxCkRUedd
asPxf1kD3Czsx9F3dUjm+IHGdx/obeBWcFxnEhyWwl0ZqpOcUCtirDRU9bqM3hmx
OwcWQFg8dNQfvxryEYFoUfcGvGvrg+lD3Cdc3kZYDXkEPVdfoFXYnmdS07PvnW2I
GN+fQ/2ejuGeVckGJT7quSILciyFVOP38YdSd4MVnr0Uzy7KZ/o6DNdLnszlO1xm
oYE9H0g2kunKfVAKXluqe3Cof+XyxDvxzHRl06iczInRWxzea7lGEb6rZGQDv5LZ
DrmIIfKpqmwG0W86viKK5IDOQZFopzMULNt+G0UuTPfDyhe5hFxMQhO7BtANq1hI
hXKa38jJEzww7BQN0GgYL6URKLl/Jg18wZn+MgowiXJSHVA2UPk5NWXe6viYlhdR
TnbnBWjNb3l/fBPgZGJXIUcc4PQI9JXhSwCk8oODELeaIaMLSbj9ZLVhmKS9x095
+8/gF0+3orZhX53sEGIPVJAIZYKU5UTEMgH0cCZOyqQWMyOaBmEq265eECbfQ+sy
raVP7xKOb2mrr8Db35xYTsObQqoQpk5RS7gpnoe3DPwS2P6mq9t3h+oF+DcN9CCY
JqSDDgbD7BNRmLtE/sXppVwh/mCG3zP70pMfwxqodKjjeoV7qwmvlCERHoXkvMWK
ZxpdPyifk1fIXgw2quse5l44D08e+WwkAJHXQc/nK+Khvgi5hhN2X8ReZqdy4d6W
r3I8RoA/I49qypv+1X2cdqolu5GwBVy5yaE7X/me0K8OxTSqxjJXkj0POj5kF2Qe
+U/rdmnLbgHOq7FuKlF7KjEVP0UeTx5HGGoB77pPA4lwwimSZX/TwqRhhvVb/wO7
zRt5Tqr7o2iHegiFEWJ4zy1iom+LKGIYAEy4aDU+cFut5r3R9Or3uCy5Ta9loCFY
6hRcjQxk6L5pwe/gAAEcEU2Y6oPBcOoyV5aRTj7lEH7NUkqKnEs+6ffdktFTofqx
6I953gd2Bom2rnxVS7z/MzNtOpuSTLNKTm8ie28jRC+mgHeYeChq177Zxx9UeGlR
vb3imJJkFOtzgElYF0Q5r/DPpPHCO0Cb8jDv1X8aVThKwuyJU81ZAbrlZXiu4wG2
1JC1w1F0d4sbrpA5vWT9Thc9mG+STIJOcI0DIkQbI3OAioNu2SnVVjJ9sTI4SDHb
H2K1aug1PcFXjhrz1PKkV3CguNB8JSfqNkoebz26Fw/WblbuwXkUdZLibnl7UXQ5
1A6P2pOmqYLVc16jUtzIEdlC42EmLXrEEZxcbe+U7d6otrtOadRGoK0kzZjGIZ7O
VIPj+pgo339t59OJZT4qUmhXHyfjeeYT4Vj/fdx+Zaom0Qyuk1hNUC+5I0bNuo7o
xJeugb9RCeXA3gAUiUAG//Pc73FVSNRXHpxtlc/dcEpuFylHvNlE7SfdxmKYUD5z
dxxup1a9ZuQOmYubSnE2P9mO4uORLG5lMuCi8VYEcddH5aHIjm1iEph1dELc8o6R
yTP9VmoiKfg33Z/uQOgtjmciSpy0md7Q94yw5EV/Ta32fBTdvQE6Bl6yDkkLxH2x
jFT7MarkMXndsm/RQwEHcFg/TkrrBaJ5xpUyscEr19g/lGN08sS4TpTyDUlxmn/0
VwkoZZgru5wB568oT9N4nkGq/mC25TFNnFrAflDHc6FKWvfTN52l0HbzbQ4iK4LX
DJra2xKSNiOpyn4pEY/FBm837AsK8RtEP/qPEPinxdammcmPANA/6HkSeZEfeg8A
N5/7ojSlRtdeJD7qjwmaHEhLZcK5hwVUEOfegybSxNMghhJAWfGYB3jIqRd13Snm
3d6c0LwGDoC0uXBdoXfGDONGlz68Z+79+2hk3FXYngP4LebaUT/sctylIcfU9aGv
z2IAok0DdGxXIZ6xnqM/augF5SfSrO4eOxxY/FNNPD8/ezUIzk/12pDMP8eIz979
x4pu3QTBLaHSvWhPecZM2JkS09x/QKRuN/rktZd+mMmuhT7k5yjAcpkInfFm/kZW
NZtZXDjVHFI5rMP36028QQrn1DspeM9maybOPtNlbRQtng1A4iLy8kM3UUmuJCYA
mIH/Wi1TH8B6jTqxLPU8Q2ieZ3ODJ+WhC0Yg+oDmHLbysSO6pXpuObqmGD76o3Hi
ORXE6cMp5RE5h/GtG5PKdatMRwv/tipb7xRU75Czguq1HTlDdJcZAqHcJ28jcA1O
V2T+QLbJEV+1+0BGv+mpqg/rEhmNenAym/A02Uuz5NDUR4eC5TrsmfxT0ygS2pBx
xUDk9yaNwCYSjU9f4EsYv1QNstOWucLiFqIdnOkKkacJtOBpEIH9rdUsM1JmQ/XD
/9i/U9xAJICeeeLiLmncbnjQmglCOC4LErPOBIuIIzFIcyd31bz1XXIfSyybGlfo
SpXVTaabRiCFCtH+IonRUp9AxoJxyrQeNx8dOs7O3BtsBuOlVooN02E1+uT43JP4
LIZboLnyAslZUlM+gP87371fGPYDs9p5PS+ko/SViZLEazl+GmZgmrv62Td/zY5t
h4qGpKRSQCsJp+pvO1DGS6SzGV9XLemoocdbb/wGxegTS942LUNBIZJx8u3TT0Wj
gfsxGjSLcBHlGq2+HHaDM5uMc9CHtPdF8To1gBjQFM/+hKSTdneqah1to4MANjw9
M5qxVEOvI68R/Bcb+E/E1Uuq0b/ecwB12/vWifaJ2utC+j9As/P+VkLhQ3g+ZT0d
bf095VoHkKv9BQSjeGQjPYlwjxoO/fZF0lDKxf0/uNXZjP6NcDm63mVbIMUGcC0E
588AcYDJOI/PPD3bRJntv+kXrEnFkCqKBPwi1I4R+7JQg45292NQJcyXhlp20YfQ
BL4Gee0zsh51atBlRM5YDvlYQGE5EskM8zRowf3uOT8s/rwv8Sq8I+CVNfMAtg61
WSMkcGNJnWm/M0PpTRQulZ8DPCe6bScaK6aMBgTpzI8I4hUsSwMrvIHHL8OwdBnG
T5E2C4tEZjHXtcHW0b4A8qaNV7HurZvtenth+l0roAj2Sneg49H6e58L6eBTqzd/
VqSODnoMp1OohBWsjLuqL3O1lS8K0nu+Rza1ey8bMm/EGMEUpG+nWmgsDIKPeeU7
lVc6666tmN6H6+vgPcTygB6XtXgXjs/LxULjpf8mc0Cf1XphXtu+2e/dX5EAJiYf
HYunuTZbnq/nE5v/ta+jVSCaxQie0Xj8zWgqMJhsi7px3VNBTlRAATYtZFlx1izd
13nHGgni8dBWqeK4pUlOwheNq8UXJ1ebXymrDQx0bIIlxXontBI40FJj3UctWFFY
5TAfrzh4bZWvpMKOeCfAj+tnrJCAZCTZ66VipmIOf6EVQMTXzswPIroSiNLEH6CI
vr2s+LT48WL0sLlZifKsAHb1LHg99BwNLdRFseLYhDovPtzwysub3GBfivOF3z/h
gBytLtcrsnu9euJSh3Aze+goyC13HOFoFbEH1VdHuU4dDROFPq5V4m4t8i5SmqK6
2ZIzHrkV8dI5IIx3it5ZrCuBQij7D7BNIoExumT65vYrGR1T+QcDnQkp++1rbfAE
7CCijouzcemnmtDezUJi7OwtdngVn3AeBqxg0Y0bw8hAv3fFkh3RyMpE9NT8nkiD
j7G0Z0bQGlSXfRyTyfPrOhPyOwlVn6AISavG8gJ/MUxGxZkN4yWoOnUQX0QCDwJv
YfOoVnpEFGFmBIUJ4TF7lV4T4eiwxPyGqyGt6+1ZTAVV+plU8Wkc4UfU6Gh/Ol01
/lNLIGm21QnXFBg1Iwr5MQujbbrBJGQmlKnd48SXbs0zSbr5+F4SsSb8fBAAH6ec
utANK5gNPyu9cwpaGpc0HVvEeBoTMbdIpd9Toe/5ESDFCvpgrvEHpcPrsgWMxZnW
iIJKmHQlj2MFcwCiTq7l3eE0aNnsmJsdhsHDwFVxUtI5rEOj5hgjlhQ+ijrrNKI8
m8COU5eKvECJpvnjyeiueCGHwpYlvZu72Ox1qEQ6T5iJoaybQ0JSlJzLeoWLFkys
vOTDIBW5qMGRzjI+sjUWwaz6bQrVyp84vPDF9LiTDW4E9YiJaDv3RXcYulds31cT
WaMBHMAPigyJMxPvxN6/Qjn/Tk2StOuY2a7hBITX8MXnsTbVRTcyEYDtTeEzyHFw
pKwCJ+qzP0ln1VRMsChkGG/hb4oHAoBLYLZWAzPko5gPUpA3Cr1fkFtKWJcsdwFk
rwplfiUPzcBp8SZuP3ydA6A1lplw1TeNdzPPYT53xqxrs5QKBld5HSlqTCa35jcF
qxWYbjnbAGy/zpErEl4jwPLesgDcIjKfX4FIFyJifWnLKPMpmn3TzRdQdbaVq0jS
Wx/opy68x85zXvd1uzyZaPPnheDTM/LigD3pBC1Phzr6lIphNK9+0iv8FqKnNEcm
9L7ysVeYZxCF6cIx0YQm4rUii7t+lFVIsTq6lIiVH6GgncsNbyYvWFNyeDdmdUbc
dNrWZNKmiOUUgLNNfVcuiXYNT+tcVAqCObGO8rucJ/8b4dW9tumq79kb9MgmgZUh
tINlIA/BtFmxiNxJuKG+L31e217H/g9SbGcHTelodyLQr12ZZqpDUJlmpP6tpqh6
DiXcyLomC9FdMVkT54+a9uUzBhcS9eyPPDj+jVcqxGLXHP/cs7aucXWT3hXBEvxe
k7FDoVHxxyaE/ecK8HtffA9uQ+croouAAlDjM+oM/b59xO9z+vYvrjPk4ZQQIwVW
YCU7YaEeMw0gHTj8mazPcdJx8Kjnf0/QSI7BwnqCPVey+vcz/AAQvyRB5hKyhlnj
awCkrB8B+cxj4KNLICVDxzIPhtVYWkVQohd0kXIfP8Cde27WGuI7MRWvtTA+w2JL
hag9oT43piabjkZ8/HuO0SgYCpFpczcDuS4ZuqjWZhCKMMZtIMBdwmnLu4qZmf2a
YLIMweEHOsHPhNAzPyibtWyF6mg3u48fkDXynBMrq+IS8iebHh9Ykr8OPS6uhqmR
uFv3M626zMIY9j/C9F5fNLcromeNXm+WSI7FcHrxzfTTkj0uTEiZPbCGSbYKar4u
l4h8Jl9iyPbmcHrQqFNWrvLE7RGgCb1Cg0O9ZxXF1xv5bB/QufFWJy1XvGG/QItM
0bY1GD6YIJG4f6USSW3njW9SUL2BM7rp8SxnpAll4t/NhgumnsTFsu+iaH6twkr7
c1wurPVTrboxHI73SXv/sSdreOV57lyW9DfRBdTwyPAgbpxncVdWdL3KyOG8K8G9
ln1zAOGxhFHOaB5Y/ysMOelcCa9oPjTFdlWz7FW2z/lc+21ke8/CFMwZAg9pWcpH
5uAWz2gUcIHIUxivqnSrUM29Kfk+S4HBFbi57lTjlAC1DZ4yumFpOchzgIiuGbmF
y0TPv6UDST+H3eJHJGx+INmAmyswkFwVwXiqNJ9LnYPIbcAR6Zh6EPbOaXJ1N9Tw
MLathMlVY3SXig8uGdko4QV4FFfOUTYVEN4ZF5+xyXr/N8536An+/WCiEPhctczF
VLwvQsExIPuaOzFoLS2CJlx3qjk9FRMxcRtynXEi5KGTovIQlYvl6I526AxFJXev
VabPd5EWiN7598ckGSA93lJew2voeh10OivT280h1KYMyuLBgzcDFA/cpUYZ7P+N
d8D/sAMtxTFLWvvVBZq7YAC6amD7nEArUMiPH4hEOcPKu4+gbIWuxc66Zpk4f3Q5
Shl4tQud9bxrV/MbThBGIjV7QWfbIYwfN6euJrE2rHGcHlWEIPYt9ijEiAVq3twR
MbmqhTmHRojx4Jx3MuWNE5lW50nZ2e8Z6T2YKBHRfjtD5484RoqFQejCk6bfv0rA
iHnPse4tiPkp2x3xC8G6SnsAPvfOGEX8PgTI7mJvcNYtS6+JtgkZQfjaows2uMpc
129JKTP87XO27BNR+x472GOKVxmdzmCxmDGNkAUYJ/4KcMLLUPMGvP+e6eiTqD3F
BKTLxY2qEgr1l9/rbJhViW1WzioL95cWc66/tbJEel4EadcBpcasa9p6VsEP9eAv
Xl+NlMtXnLwQQTuvxR8UAMqD3JsonyJaJNRX1bHNSsKCpSFm4CeqlFATz6z1K8vQ
uvjtWNMpXvUsQF+OoYvagkBIy4B0xwbvqFfFe6CnOOl81RoDdfqB0BJTB0SkLhKQ
rYrcnaiVGlTF8XjVXZwIjOO1+XuXRL/ZkOphl5/FIDWKnvmG3UNxZZAgUmQiYRTY
aNHwnVXyRsC8JZxZyVeQEg5/lQMdgSKlKq9TWWGKDVfYdFW4r8AQlcnKT/c61v+Z
6EeF4N/D4F4RbJK/6FPb+REpkodT7cg0ixxrUD8whYP94TiM5LzHdt35wLMOFSDX
MNdMIuDitdWuxn7rlZJ2obHm9LInlRhpln8pFsVW1GxKN8ilTbrhl7g6nuVQpTpu
TbCA8MtPEFF6lDNItRFu+SRCMzOSLxrReZOLHxNGSVRD/tjEvqRIaLiQvj2rUr2b
u2ZH5WV8BCmV2lO0/Oqrm11DRCehnS0sh/z5dwZFlgXIqJ/MMTT/YevZ6lmHK1MS
gQlzYYomFmidLJEGAi09dr6Acmq5nRhUvwm2l3HPz+a3arnzgRpZcFoGR3YpgJaN
zCdl+jBDVdOnpiCtlA9/foworiL0WI7/GcwzEf+DrAwjunmhvP8FCc9n9yJyCjWu
EPnAWR9bqddHnykP35HdHeY7yjOqPBMyk3m9r6BUPcSjP7GaVqOLTUq2OQbihhBg
BxuJrQtlniUWqfMwMaOvfZ1Vie3wYaTV179yhvzjUKGxDZoSJ6MwziflEyJHPSsE
NAYd9WY02Y/phgvGUwxuCaYnKqb06tL7oiV6pyIEl48SktloTqjtrvwrZ3gk2pN5
c2yFtmzcVbS4E9N1GWm6KwtUNTJ9pzKspYJ6PzEKDAIJIpJOiJCbInaX1P0OolK8
dqzRF/OGAqFO8ZdakhQpSCdV6jYg8Pwyb2vMpzhYl/SU2egfX2GVXIVHdbeLmqCW
8nSAYJUZc9wn3SjbczzHnTA7qPU6KSZf8tOoWX1n5kp8DkigcOVJ0NBzkWL+ngMN
djYdjarJ56ITJk9kcT0XFDiAVHZFSAZg3ZpZNl7kXb8uJHtoUaD94Ef2IME4AnFZ
nsqdWAxNGvGeUSMR+UoLRPvxTFI0fcyJEF23ZFXHT1IQg0K2Y4WiKC6Tz7D40St7
sKCQpaTrrVx5AJot9D13L6m+qd9sgclOYVJn6Or/vNRan4SYnDWjOREaNtTEBR4S
YX4WFrOuGMw6+MrXZVD6vwsWnoLXdkePx5Nl3j/Y4hx/sSZGE4MQLjyaQN2QT9MZ
113dznf3cra0OQ8BBPnPSQUL/uk6gktXUZc314G57SvfWDfUTcUZfjE3HPtB2mrf
AKby4fn0PLB254kMNN3wCqXiIw0/6US4RUjkzf0cKqxF+YZ3ZZv89QOHRiz/R6zk
D1m+pebc9hh/erjtF9R3TLNLQnSnSNFc8sx3OVdeKz4pvrhmTyBnBin90bRIUroM
K5YdZYdln97rE2bZ5WkLBdnkhIiFhk62eA4Jd2sK3WeZB6y19HJx/0wUZA3N7JBy
oOhPcW/TBOnILLEdN9RtzkJDr3GP97tKZHdFjUW6EoXTuMvHnNMUsW8tN+8LA3W0
1d9MhzcwmKSqjJy2CzL3V6Gs+JoQokGNdyIz4BjMpj68ZbQC2Y7rD7NhrgQ1ZUU3
SFQlzw6JoZEhpDwhJ32mrRDWEian6HphqlPfMQC2NG2Vkag7qA6Og9XAP4srJw5y
vsNxglTkkDu/216Swb4/QPp7c3gM6+x1C7Rt+/WyGBD+uNdRP4SNfylqybgNtS2l
QtUdl0j+BNFUgtypahjY8qlPEZxVHXQNUGoJXZ8CUtMtKHjGi0Mm0231bGiaTQk6
SngeccNPIfDUtJYtDAByIlXMaBijop7xECCTMjsGH6an+Rdu7iSo21Hkp4UTkFp7
Uh39rvwkIEYYncYdeMWYB5zQfr6JGJspiSxZqofS6lx2Kxj3A4pfSIGbRm9tCWVD
SjyhML7t626FlLdtHkU8ty3Ypawc+W4tioOHp95JcsUWWf0rZUtdfR65B25Z4wMn
l3dttP9mCCN6TtFKzquJKQo9YLhqcNJp/W2hu988K+QDkUbo/dspULp5BhJGSYD/
7zGjN6zj0Xa7LUVHfZIJ3c1DV44VPvnfcGZSYZIvX/pTcKHoVy3E3w2/QmKirZe1
3P39QA1kuu9FwYC4GQlPWxlbto1lTFStzFFwnamw+ULHeUAEsv5B4/uRa5Te3AjC
f1r1MmNsjjfoAJbEiYXt7xtZiQT9ez2n08T5YDLhU9FbE6odeMxlo58IING6NEry
XXg5mdHFDUY9znEFQt1SlKxicniwq9R0cmY2+VHrkewef+ogesUCH5oXmvWYl/fd
L2nArnH9G7hSnZiPPpZzlTLz0FlML4k7RWa8dYpUEMv6b6mb0wFbt1U+cUlm3mKT
pztWsY1hDVYvG2h6h4dPC9gYUECXJDUVWsmDCSVo2PNxi90hWBrX+CCGboOIOzG2
wJxXvTx9RpocrHRXTVIgSo4+WyFdtr1Mk07wQCIB/XTzZYLsxIN0AbdmkUOTy0Ux
5nDsi2FFMF8bQYVjYlzDr/A6NLLHK8DixwBjSctbn/E6Sy7larMyF3O7uUGOB+av
BVx8NYTnNN5NfsGH4tTHBFnOJp9rBYO6jReRzrb8Ldq3W6U4JbTyqOWrmLNUgac1
pM6z7q8GA1V9aBALPzY36Ks3N2N2i9qAwpI5/yD4i4mT67+bq28pRS6Zki+CmD5l
7/1VkrgcVtGICDQivHYrs7SBjkL7jcHdGxeaIG22bJvnDVrWoMpqvrp7DBFjhv24
PqQUya2Au7NFQjG63y1xQpFL6uUHf7XIkQfKiYzpwXcG+RZfb0jMbS15XAFuLD0y
VpiLyAVDlxfvCbZ3KNQxJorsxPUr2wOeJBtSvY5mSSHQk+ZJc6wJrz9hS6tilmon
I3XU1NISSm+oZik2xpOeEKUlDGE18JufSu71BoGNG90KL+fwZcU39lV8lhbVVB9H
iWonkzmDxPhetwpfZSusn1L3xEa6hMI9SCVgWoUj62Yy0L9jowvtnAw3M0IMghEp
0DZBPWHePHu7xKXiwOdkRsewL90XBpZiO8y5WaGxV1YuAKQjqUPKsufvOU5i0BNb
XtEeuUMc3IM04gB6S+kx6I4aaPOOuFLcDm1+3/hHjZ6sTm2Q+cR4HdWz8NZqgyWN
8RzISu+NfcCxH4u1ktAUFpG/6rt/xR4X4D3eOFYxKY5h0wWtzaW4n02Yriwu1Xru
lSmrqaObLpyr0teTqY04EihkkZnmvw+/7L+VFB6HF2JVe3ph0WGjEKwW8odk25ev
Q0PG3Ws7g9VjbgFcKKJzkXdehmh2Wl3rHIiBdx8gXvWVy8yBMUxQphncFE5sxZCP
XuveSzkL6P5SrrxmiUFhNoQCm6nUAU+xJmbowfo7HxS58ld8u2/d4lWY4iPm/at+
MEiOOvhqJ6mtgLJLwBESAsLLBveH+pBb3jEJhLqHYy8Xxct5r8XeC53p2P5B2AhP
ukiyNyu1x+K1Tak0GOWdHro5BjCzwbZwjJJi0i/PlxKWLM9rEsbU+3v4b5/Gm5xU
+YPSoycRP1FHcddaa1c7Ow34aT/wkw9IwMjbmkRxhVcCGS+SJs5DUE0N46bGQdE/
ZQdLANEjybSbzmrnV9UzcruhqtlCCD0ZpdxGuwC7XCNOfkFRmZ+feuWk2PR8W38C
9zGgn0dyVuKwWajnIxytcLqjtuas31BwyblXc4BATfoyL5lqSX+PlJRKicgMtz9I
FlyPdLeD04t/SVzL98Es34kO2RhP/PybMF2+k2jQ0Anew2Lcb6pqpBawA+ZTfdQ3
cDjnjxxOLAmDT8Do0p+yG7FD7zKnl48Qcy8Aq4i/60QryALN+TAdZBqV5esUDDFz
ItWRyRakHQUSV8XIHbqTQIy7k79knaPf/nZO2aaQ4VCyDBoisQ1b8uShKvNRTnBV
E+/vfeinHVUs9J/Lc3kJ/o4/iDQ58mM23f0ozbfbz0fYOn7sBjg4Em2XhmL69fHL
uYNHkOFV2lSD23kD6MXEI75njqpSlJC0amisJzZfVE12DGslG0gXk0MlI3t8U2tr
vpMkyAXmuySGX60HWJKvatx0BYLg5d4nUyZGNIo9VSLlqFK6Lfthb+S9jPG2dqeZ
WCqll9j6M7WkFN4IfTzThSGN8rKJJp5m1QHOBZt3rALxvxD10+w6orsuQhLYhmd/
jrn9E52XOVYA0xOaJqZmY0iZLN4MvzDUpJnByQF+yOVr5MZCDfrMIJyrGHkXoH9y
CNmmeo24bcwzbfei5NMkn1Sdk+reveJ6InwmVO73H/T5fp/jq/erC9/FXHvrCJch
xvGZE7Da8qNWkE9yu90H1MY0eY7UwAPQEMOFaBUQBa/Vi6R3l/N8TpNVdvXPETsu
uR5Wmqn5Todq2qrA8//SPhumfvSNtQHdU29Y18v9y4L5ZYZJLjtwzEf8iOucnBTR
G+344IeoeMSyTU2TFzMB77RPNKHiiOc4Ot8C541XTUcW6C0wCELPC/xRFzMjsoww
MQCZIYh3O9hd1gcDjaokQodSsx1X1LWj6oF+HQxRQweT6A2wqPtSZUJqguYDwYIW
yHdWO1F/VZGgXZ5rSKMCTfB7511biLZq8+cjaAs25LCJZ3i/DnGt4Pu0z8cSBTn3
KuP+yC4PtG3XeWgx+TMbd4T7JyPBstmbdLmgNucLH2o0rpV9Dmq/V7HN2/nstNyc
PT9S3FfLk/mmB8nHRssJ4tCWLkXCsMIcBe+W9/iJ7tV39BADYM+OVxh8vruPghtc
L7deu30zIgBjiYMhYDgm+l+p+GtzSpN9Y1mXDE2XPFooY2cBvRKEheqJoLycTIJn
yY/aPU/zs+VBBvEpL5Aa/qpg0BSpeg8EkuEw7ZZe1oQo0k/UrJthhs69qyZWFE1u
kOYNEexEvbFSj9BIxkQe6CGF1CAa3SpBtW4Cu3RMNwRXoWPyuEFMH3BqCE8XF+Yy
wmp72JsZWzytSVf8p2ua+wC9JSgrTOE7bynnSVkuqmVzabxyzFheH54cklf4gJ+k
MY6s7McZstNTtKoZi5GGRJYaT56lINPoQbhWpQuIs8VLFOHKNcCGKdviXQfwO+mv
DvwpbrxvhwkGiRF1ja2xa7mBdAz8Ef0zbCJZgJa293ueKD1LxuZDHEOmLcV+e4dK
qTXHdGT/4aCZtNYBmmjur9oU1WVTWy1n3TiNRW95FNNrL2+Y3eXmL/ssUTKTB9L4
seqHtRbFvrhVd+qaXON8DaN4Qp/BpNMaHsMFPCTuCmWM5Q9THBM+uGrUi35vd3PS
izHyCTyaRvL+Urb4AeTtb8QxquXuxuxTXyx6S/JHkHSPE5OtHnhi+gAg/MT7ptZn
gYdRZ6YdZddioaCJhtnHyWP7Rme6aEtX0GnwutWVKemukW2zldjEUgbkNkRO79+S
BvI79OjJnpaZSe4EkFGPtNg7FRTIZJTU/Td0qLwFb3ehDJkrn4yvXwfKWAZ69k/p
TfuwClavWV8/ln5OQHQVBhE8WtK9atAsy/H1P3A5eZHP+sOPog3WZP3dOEMrv3St
xW1nw6D76xDYkNraXQnDEKPB1jj/Pu+sOO7gChgPuBxlK2TtAtJLf6cZFJD9l1hD
4P9TVDnLOhRcjelm/6imhdxT5emA8jf+SETAjSELvBK7Kpxj34fCjw9+tOkBRgLW
90n7A79e8DE2288PrU8p3L1wcwcYnZYQQ5pDkZRVclQNpess8Un45cwmIqA/ThH3
kxUPql9cbb8VY/fK0TDZXMYR8yQ31lKtK4M9CtXRWxR1QSbihmhxSP//8hqzXAn7
55FnbjhF2deLWa+RUcPAaXWwLd0RP0ZOkBHfXhTOz5IO/idIvgcFKaoQkmqshM4T
2JHU4dpib3+uvFBtMKfXzOMpqhA5tIDCe9M7Qn6AlkkcBv0sk9JaFYgKlv9Ao+rm
lFnFKrKXYHT5N3WGbddMzvgKjVb7QpWur3FT0PxbIclN3LqrsNYfzUfgYXopbFcW
BUNGAJO5nGWHI4hrspKpPoQC/qxuneLVohyW2Q4xOxQ23Cj4ZrYbm3VfI8UvhBg0
LxLJF7+v1NoX0J1qWhPzgSzOy5u7ZSg05mioVyF1GYQXNIiqV+uKdri8vSVwre2u
6LAdYQRMknhZrN/zTXzJfPgncU+EXpQO6RZqgdMz5dgI1iK0gZXHDnG6uEaYBqIA
FU8iRnbb4Zzf6zH7T4dl/CI1zKSEwtlibWcCYpb729Cc/knwvvTmuc+wCIpMDo7w
Wb/jRdYOAwkrV6SHcAu9CxGzjIssarpLlBq0A2OaS3jGmVidq9CPt9XXJ95ZYtrB
gqJMsxUTeqfrIlizAtUa8ROmr6svxfFOYgMDLgZjZwPZTeuwOwCacfNs8kubeePy
+7+dXxg5drc7YLsQH4LTDvxVlg2EghO9uN7gbrLM9atTnOHo0JCpZngqWyuFBF8a
uBbfodFZGJgwuIZXPiYCxomBiLGAUDkhTi+Nax0ZVY2cdJjTV2A2s+l+CNmOpHGQ
dFbHsaCmIGceFIsX1jvGjuIoEj8pBRI5gYytc7zd5zkKVD+77awT7hjKFuP4pmoh
2OJMKD694nmCCYoospBagVSScmaRkRpJVbmM9c5VG1eAV+wUqI1VFxi/Bgij1T5j
10ba6xW1hggX4GITEV+zRDYei90Iff1kKrYer/MlPFK3v1UcgbIfkzheWA3hFssQ
daS31nvzrbiqOzR7besC2L9ZXXsAYiS0t+tvsYTqbOo1VsjwnlMwUVokvl8X9xqt
oh+i7/C/s1s1a+fFaKnY88MPNCtYeT0HJjJqyRHcfEpajuOwjU2O9kSO3+ROe8/W
pvteAFFkliZPv/h+AefeDO4Avz/VU9blf+YBboRFtBZVquJsbzLbh8QfEzeLR8Pg
jMLRAwoxaY+KpdtjCPceg/DdWuDMelvnAMx9JirqpyL0YwDIvRhaxjwmt4PZuosI
I7beKi6w6kVgKecHf111blTtaEshI3+6LJhoTAxQmyFSh7a5h6HzcGBPWAKHdEVi
ilIFHDqbv84UdDa157RK2JoR+IwbeYxOVmerZ3H4y6nuNpByDcMDxVUg7Iswj/bu
e+kF/5jvqyHTkbEMJcHLKXwhc2xRXJDch24eCHd0Y9grzqLxx5y0eyoEL8WhRRgK
Rr0yYVx0briiLFVSIWNzIkjow3RytUTsakKntdaZg+kYYYZ69xHqB56QdCAWnmWo
c5j6gMoJgS2ZuYl/WKgPswuK5JCvNWNgV9qxMsUjpASr2FVSmuV6pPMquiGo312q
0fiK5xPI2JMDqzwGherteWN29r8KH0kb+TBwr2dmRV3s6LlH3IfLIC/SHluQES5b
4zjuP5Zz4Ban8lloIbShnPg1jl1FFtIQEUrbG1AZWU3GOCMNv67Az88yFCLuJVOn
U1p5UElJal5lobsFvFNzhZX7RBir5STJrrFqapV9jxjUBlv8WXzSBzKJqf+fA6+N
FkmN93OJHPU5dg+lvFE04LI7+frxcILOihsOhqijOcWWv9+531vpetAkDWNFyoU6
cSaih+ADI9r/3fuVt4EZ+vqKsMcf4+u0BpKLoXTqbLJz23kSm+a5IoadZxgOBxql
AumIhcjzOuHG4qFKnTEt5s4+pfSwk9GYeagHsHWVc9Q6ypV3iuWiE8dnCkUJO6xq
SPMnWyC4PNUskwsUf8Q/xNJkAlbRBkZ8ez7j38Ud7u7BMtaWgBCIHraFKQJunUBf
KNo9/TxuVc88I55pYVzyggQ/S0vVCC2AbcqbRWMSok9O4uxYauTjPRVtWMQ6cT97
Gl4eHYaNkMMnDyUF/nxiaGaqrHPOSPeWZrAMliu93dFtNI0pPqha9QW9qGv9WcyI
Q2O2ciuBb006fJKwizCXy/1Qrunx5aT/ZT9ABck7zSfM4Kr5Xe6sRqmqakvh8egU
ISHXEvZPPP6YFO3YMLxvQGtsfGM/SKUhhbvJbBTfvrl3FVBeIVa7t8iADS1/wWbu
mh4J8t1qJi3U/q5/CNnn9+kzP7w0gBVxrQNbmceB+DmcUoX3iZO0M0nBISG5XWCs
6+QXPKW0GEmGQiPhetvSixAk5JLGhWHKA0GZN8BG0LjxKepnwDDKE+OW/wIHWvzT
69d4LbP+/GRavoIl3RolD8XJN01w8d/svEFDVCVFU0xKBJo7BjCe8IUnS5HWiUrn
xCvle7B6eWCGoqXO2cFHqY3WU1FigF2rj7fhZAIASjeQ6QUe7KzoYPfSNFpoDjR8
ei3Xh8lQgbRTEIGVxoRLeRrxzzvE9H1A1ZAOiUOhol/gP/U4aoiT3btMa27hrIRT
juT+UVJy0g74CXU1kOlXpDDCkmUh5ejcUokAYoK1Aa1xtITia+V0D1swG81wSEUh
g8XNDAIXpis1eMzSMwnas/E3r/rqgntQqTD2o8rkr860glN4s4OFnM6+fOuq5J2p
CHdWaNVqJ0rd2HDJstyRUZMpG1CaU5aL3jxwTxJ137VDpVpSy3noi+6IW4oO+EzP
xWBOcU5KiyRfbcwqdLVTKtM3d1hC014ENYdXa8p94jz2b1rH/V6TbYvb4Fmj3UdB
3giKSx6XMxlzUKzYNZ8Z3nG1e3sjTQ+0RXBtlAiN/NWMPL31TR6oCm3qK0udkIHk
rj0XE2DEHc6CkyAhXze0FCAG+N/Tlv0hSF4vt1Xc5E2wxhrsBx+J8hH6NszmOJnR
frJfuNIwYb9ThQsztfnXApS6TQsl9Gt/M5H5oUMGkFrdmiP5yzoWRYYbS4Sajk06
TVZZ1IyAxFpxWaOT1ICsz4NDqXcXRn0YBJPLbT9Q2FzgHRpE2JChfOIqRl6hIyJN
l5giSfRP4cDjS8VYe8AVApN/BziPns3HNjf3H56gQXv7CrzPmRA52UsRsQwD8ZQP
OJ3VrRM2QZReT8mHi1OIjeHLlWMfkePqDT2FhRIx7+THJ2fy8+inTtctHJFj0rVI
HjE6vgbs/pNKOwT6p8b5a7t97uo6iM2zUojWkIfQrMQt8+vV2KBiYz+ejQYrbS5A
zbs5zXeVLOYsUWZ82QgGnpOVBDoOvDH8DLr4h7AnmezinLsGgqcbLHpE3QXOWHbj
HoGW/i7TwVukRB43/fIU6+noIRBJ3GSDDwg7L8duqVybymhnA29NGDaeIUrWyu2W
LGucko+XK6CkGDMAOAfCUOhTFlhUc6KydlqCRL9wCDqx4w6R7+upsihp2EwLnFBN
Z3H2YOw2cMU6zylkXzi1wUAx5HJ/glT+Rrg1M4Ibt+PTq9xRBvWGn1Sh9jaZQFPP
rD48mmapFUIgVbuB2gBgGlOjEx6Opoo7nZZh26JzQqK19S49nzuQGoFNaI2QuA2P
V5KBZYbpbjXyGaDuF4/+Q1ossNibozR2rUmqHB0QPFGfSF8zEYx/W0o9VaCXYSus
lu+CTj5D0PZ2fiBIH/gYeUqksQ1Iv3LymnvkP8GMOwzBRKMwNuZ++7ZVCXWPJGOU
OMfuKbYXcOg4HFP7ZBfKSIx888P3x6zPjEs1yZSFJlsoEkvKgbslAICTTrURf/02
IZsvTFxfumjn0bt0N8oZMduAi42mNc+IM4bhinVrOL0c48RBOLpcUfi4/OJ9g+e5
53CJW7nUCxQkNz6Y1KFmOc6S/G9LG5GRetUW8dhVVE3qaw4t43y2KtHuT2Yxjdgr
iHHmno02GRadYgIrH8nJImPQXYsLeulg1dzjYshgvvJ0DBynTIozEfXfMxA4KPNY
xD1HENKvdkP/LgEYPLQedkYS2It5zt7/TN5uoJNUrV4VtkxzeSRIMAMUdTzKSC8j
A8nKFtQOueOATCBz5uHe5Lab+pPQcKPoiBnFT9STUE4QBtNafG/OWTY0Bw0iafdD
j+Tt8imrHVOq+pLCx7AATkYHIQiFyiAyzMLha779lfzqY4MaS2hQ4TNv8Prk2WES
Y0iDNFiP8pfk2opeCK+OrFU5z0MK2ywtckv0DdszEyBaWQhEJYA0RYOH9d6znw5V
QiyitUY/OCCHG/LX5MGFdAjr4T7A46NnmuBXpvm0WfVtJ+PeXjIdHvhZcV1qcbUQ
Z8+ETADdBUis/rsQYMgAa1ZWA//W//MdeP3JHK7570+hMZAoV4CRYlaX6drIWxx2
US92B/tW9CgLtPGPEetwxzlzb+149cVmqLxd4Axr/xUurXmaR/xEIw9PEqh77acn
Zhc1PQwr8KafB1NSNvrmEaxajmlokdKOCK6pOV3uputZe58ArSJLDRURijHmc3V3
lqg5NqNZdoaQpxDBFJj0Iu64a21NbxjNp+u2RG+O1f7eyf/0UdI+T9iKmmoSymw4
RzMXPCZvqsgF/QJQ8CB82gQrgnUQzTCYsqolhlgemhAjXIGwPOB9NxAQWO/SOf0B
q0cTvE2JsTy1gT7f6l6KEjnPADY28toNH+uB2ng5mOI8IGqKvBOKgRGjFoIPBp+W
NXTLJgIPaz1xSoUpKfB5kIsPcvTNo5zZB4d/YpK4H/hUOTRXcT8cb4f+qVH433uF
gBJdqixFTN0EHode3JvusPAEdxr5rBZdPIAsn3Qc8n86SMNRpLjGLTLjiHLzDCGU
IYvZqGy9eMfdPO6p3WxehlnV0qGSntxetIo5DQwGrm29df9WQxlrbRpaFeNJJf56
hNBzxCNLFrRItT8LzxJ1dD32qrFAuJ/NTHOlcgDOkjj9s6yV6qsI6irn3Amun+rp
pKrxwi3noI5fyXuL6Jg0U1WKObzf3j5/0Ftd3g64vBFJC0FtJ06UqUHKzmFZWxXp
H7ML8WVjQgLUvOl94Isy34Ix7gYI1V/Tf6JVRNJvL6DcRqFUWNRUMc4U025f+Kig
XRy2RLz9ko2b51q9FoSMXm3aLxD1N8/xBXeMau3e6ADHnDAoXbWBtzpxd5Y/jFtJ
jHsdUbi/MFKwZxrRtkzI8pJSNGvl02aIjCJ4gzXRtC3MV/SMsNao0fFp+kMB98+2
NrGemNfu/l57IjGBeaLzU7EK9Z8y1rjGYgsETuA6bIT/S5THeyWoMqTZMbNwDaMP
X8xZuynVhvZHAi5p7TWb0dITe4KPoGg+HiKoKSzZHG8VFDuSgBjwkapzxI73M81j
jiWlYyxUh3ohbAut5FGGWkuGt7NzLKMCh08A6Q/8WXouBiZEI6UorMaWS8LCqnZt
RIJg43Dp3Vmoxzav4k/oGsjxXagOqUVfhKI+giyi/XpKhqo7hWPOqXzF1qpgmUYO
hsCG4rJ0C4IN8DQyFQlWnvLzHPX4CLBe+/O5ZCzZkBKxAKZOBYGEuHxbG5VhshRO
rr+bGhWZarwy+qySGETkjXtU0t2JPtLp65JJL3fyBskhTNLPQImVoaHYwCuiPXF9
MaCr+k7QrffVlauenJFr4d56ORYxnXTzL0w6sh1qOKqhlPXRMplDPhQp0er/M7N4
bHv8dqzbCfzXB/M3kH9rkigKLQ3n6ei7IQz6A/tj+gHFfcjaUHRsK/6agHAHm0M1
h4uZvQ78C66g0tD6kMyaceGuMc1y7coxB5VvT7gvcDxUvzUndNJAKKRNbNZpW6fg
LeeYC8Gd1CNSFNwixIJwcyXk1EPprlJ9Nim+JvZZNI+3QmT9PZUjkF2yNvO7Y5PR
fksy4DTwTJZAVZO/WMYXODShhdayHSpf0SmptEOkQ6Yzonex6Ilz2ubDJ0Q2Kjl2
sOqY0yA94uPesyuAt9pTB7Zh6tqhaXIEW5+vnXh7g8zifLch5q7oEmvE2eMcOsv1
LGtJ2tyxmBh+Y18f6Pabqz7xdpy9LHYewybPilg22dETBEtNE7dqVs42T1a/NN/Z
U+p4qCw+4EWuLkV+xj2dsq/ZlCJMTqpzykk6PiRZ3tE2FB/CGvYrmWm1zfHi0rLR
RUzgGMNKOgDspOUgffPaRNtzkKrO24C+J6QabPZaLnBYe9wFgodDHQN3eZrLB5ar
+wewOY55zxn4inMhsvh9XGjSXe2zVWgDdb8L3iIfZh2A4xU5cTTX/djvo92PDUqp
2pPD0646vg0VY4LB8s2HWlxhAzzdOsCo+Xj9ShgEpQOoP+Sg+RQkyKTSCfffMqn1
26ZtWStMANHLNgAipUUyaE9w7cT7wjQYCIqBf2cK7vs+IEFGJc80jZh6E+xu9+DN
Teh5XllLWsnBK0r61SRm2RFF9+DPR5A/3xbyGH6+rz0nw4keQyBxCRoGorgh7TcO
op7sEWm4hYislIKrdbNB+1/dBZMIPDhngZwecxJhdS3JFj5UNEwEdG1J44bGwd45
V0K/8BXrY8vGTRmsoynCAXA3w4l3LLkirkXivZHR+PvdbBKTEBSsIEVJWwR4KPDa
w0eKgkcdEfwOZX+5R+OiLIjVtt3RU+79KwCyinAU3Z6ql0/CJqDGcT5jthlGg4SO
n1Ev5fKRo5X69v990E7+GEMMKa3i7jsoKg1828Yr5X866NkyKjWWKNPXcNwQcpC3
TTSLuMK4pKCJxNrk9FI0t0uiBAbwbBqAW5mPjAWhnSuH03lQImkuSo6UWCSzSFlO
RSe3C3zS8dIeEgHadKsCTuRq1u/alUTjbo8wLc+Fls8yv1VO61Ky6OvgkQH6R4Dm
lmHlY4tORx+e9YYvTZiD1h8NbKdF9K8G8ebbI+JnmYBc7UmukxmA6jmDYG4Ggr8a
pAlQ+1FOgoTrHjPMPEsXtk6eCKkFh5I7RYJpsyYCwrKVGt8tONqSgLdfKo/mvcRs
9LjYN8Tkam2s2KkowUoTyMtIBADwyjcX6GzRVaaXmsmb1CniGf6PaIiCtT5JlI+E
c4BEeOllYNpcoWUoA9MGNaY6Up+IrlgUkDj7zXV0RI6NS6eRWMibkRAops5dyYN3
5WQz+aRL68Rfbxo/gKtsFFjgKZqAZyzudql5buZkEI7iU32CQZbc9vd7oRPgvzm0
jPCXEzBSE6FZw31djreY0CDbcTzoXh+BGOum5zsABfGmMnATctOzr6YUHshRz8X1
FiN4U4qXb+j2Mgb0pmB3hb8u6ar58P7bvi6DPrZi6yHULWfV8HTXhmcLsh2PB3Ye
xXUlvtaP/O7Hb9Z4iQLhlS9dAv7d7aJlg1z/P7Wnx+9Jk6bUzz5TXYk2VoN7nRU0
Ua5UIkjHe82fQUlYFfANpArdwcEYnHxRUMYThvQohxFtajMamWCpx0K9h9eJjh0w
nssc8CDuGy+vX9Bj00ZdEKxuqaUcDFROcLxqWnpwNnwDkzArT/5Vu8tT8TJCo/zj
6wckItmPrHmGJ1XN1yAOMWkvBM57pCkhC4I1Y5q1IWy8now36T4w2LKhNTxCv9uO
3+5lyhPtdMDcOE/XP3kipNrfiGeW6itdTbQlP+fXwG0FAOnucRaygveG7n/iCsUW
q0J3mnd2J27AAtIb5plmADdMWhtAnp9Ns90TOm188GcXb2pyJnDrTjJ549ctNbdU
edG6eoi9CCjXoOBvRAudlH8fobo35kz6KyVUqzoK17z2A6cqRhan8JDDXfG5VLpD
RqTTY177UyZnKrfZJqvpAjBhQSO8OxxST7D1Ykv3mhAe1rm3KQHHpqGjSqFHlk57
S/a0HayalwJ0NgzVMe/zczHq/ya6zHg0oWTcUVmBj3UjDXwtVmAUujweOMjBJG03
g6QmQ7VIAs5mlSSbkPbS9KPlivDMuH8m0gj8+FyOaLu/MeBz2YhkBjoc3y5dNGkN
/KHnZOaLPhlEecytxvw4iO0GV0MksX3odyBO0s57ShomyqIXYwg6xe/J9A+oaIa/
XC7BCjoa5RsoZEtdc//shZEURWVm5nrQr4Fa/FzniO1NPTGiTMc/sabxjotU+ftf
KAL1tcJuM+N+q4dzV9K5rc7VJV0gK/NM/YQpbceelmEJpcTDkXeuce1AGv4Ei18R
x1auSRnnWF75J9VhMmrg9YwZufgurKbPWdr5MWyAS0L7IWfolU/MOv+gHFMEWW5I
Ki2dF2thByrGvj+NLlI5PrWHTMea4bJlHRgmbCI9m98EyZWQMi88kTWAabFS2Be+
eYiVvFGe7txLeG7qmyBj0XKwroNec4BZJEmBWV8AOXB4muTFzvy440u61H2Q5GxZ
WTe61aS1nuWfC+Cb8r36DJqDntYQj8VtJaJ2thhDa0IBLJvfdaLY0037oqQfOqCQ
XxRMGXYrGHP8kdadY8ApsgLxb+/Wgk9gUCKyCCD9lkpSMTMD5cLyEQQUu3kicYIQ
G+47L7Mz7GIt+1Kotb/7dJuOtRMDh1NEKLSYHNzzI2o6FwViDc1OeLktd1dfZRvz
b2RopUBQTZj6SmgiVl9K8eSh6Xhyu4aVGQNh2IE9f/btJqyvEit5FQ233BppdHol
M55gH5LUF4Otet+qsaOfCLm4NP0um+x1LDf8x25ipH/j7ZVDeKZ4krTf43z95IUA
XpflyMY1+R3R7eVV6jRQVBXVJmjOi3d8FIKBCU2N35YNTzvOJ6U96ygAmHo4EWV5
+b9wAL1E5WS+wnBVnB19DkEKZe7nEU/znlIThfir9VHyAlopXbj/3DJSSJUNF8Rj
CiUvZXuqMOtML0U4pKnaq87ee1XVv+qGDqG8j5kFgNZsCwFqs6takYHVzml+Ilol
arGplcdVzvfQaVZ6tg/uZLBdcVjd2pnOx+21HIowZrUx+3r+KCB6JGP31H4UTIl4
2B8eZGjyWpkrAvzH9c7BJiaxyqNJQDBByU/QvGiZeRajtOGYC3hFx+FEltv8Q26w
/rUeoWGmkzBVjGJ8I8LhOTt+MxgCTdntSsSXtv9sI4ialgjkv4WMyVk+7d4n02z0
7hAPA7t3lFeJULRmTQjVkB6j1SXs50XY494H4sVDu1ONTMHPzDW7rE2qeYAvO/n8
tkjeRjh2i5Pm5meT+MRnDpFkLMt7OkGQfFtqNf83anQoj3FzECpeecAXiEvfZ3JD
iOj6d/OFRax+vLPz+chAmwSFtQKyfLrbDlFMKq1ZPUIN1amJuWolHq+FyfqVeVAj
RThQ1QidmPambl4/YqW3gtjZyvNucOlXb4ssGS7AsLMizjiZLoL9zufL7z69d4F5
biJC7B/Qh2tSGc7FjEnCZg/+R77ZrCPLKkOB+hHtPK7Z4lFuk3UOa5qqgSkcPldL
MZQBhqWbBkCHvqmUQ4Hei1C7YhJK7ZoutjfkgZiBT6toi79QoFGj2RQE6u2hLU5g
AmGrHRja4agsDBsr9P70ZoGbDtNatOYZ1WIamW/txXSgctS9HpRKrnZC3RaCpsMi
GWCn1GfwKn6KFctR1jlJYZmIZKhJiGeUeFASdMS64zXQFeGwK7+s1EJZXHEWxctt
ROPvQEeppIE9Ye1ZrDz+5XOTn1LgSM+QQzRxGPACKp6rWLqT7Rqa7+fKSr2uDLfA
5V3Ws1tm+gapdeyfJW6yUy4ez2O38+I1OuL5wMbOldnC6YgcBLbGCf1k3v6VridN
TgAjxqdaFbubalu1hrO1BWfYKDRW9Qqh6iMBghepVdyqItMEmB4J/RPGC9hJKCnl
MFfRwbwSyNZ6FW5Qh3Mpgy91c4lExWFEqzhdiPbjBFFLfXDM/awNQiFzsG8gIf6W
FSYq5MKg+UnxeQx5KVK2Kz5Z+1bjmgoOLDMfzBcf7zfbBY337lvypH2oCk1x5wuk
jpfF7TTmIxV47ylxKodG+CPpJGvQg3yGJa5cV6844ylPawV6iZDAr4VWZBnZwieE
mQv73Pf/0psElPjjAUt4kLRTf60ssfiW2xkTlioExnkFNQHcQP0OwCnu9U6REBH0
SGW6KqWhp5IVmU2ioHi+VLVWvu1OLc82gk4cGyYHP6aqKVSc5pqhHauJWyOldQQJ
t4UaBkqz23THLYS0a7fBqiWWJkfxUvur5+i3OQ76+NJtdlSUDtBfr17qo0VzaG0C
yHeUqCQ8wgjT7ogbMJXCMnj/b2OkOWidwTaa2IKz8yK1mq6XsLc9dQiTP13phLBQ
wCH2ft8c6BkviDBPKgHnVY2uzUiQ2rvjGp7P8EY6O2VZzN0Imhl+C+GAdAWFSZvt
UKKgc7WkDkiBozwrXCQVQRPLEfrz0Inj6BQx1DhREN281NmX6HHZDdzhsC5Yhn5F
f4w/e/fRrNs6mjjC73CiN4EvQAqj5EK0ly047cz1DPxR4WKmMFc5YXa/HPUi3TD+
HiZH0Gfy1PhxE4X0Q68sLFFW50uRVtx2IIZEUkBv7jPrp9WaQVIdnah3GVxxcRA9
0vnL3tUFJXLvQhME8WCZrC7fjiqD2D9j7z6Yuav14R++g79CLRo3RPItZBygYDWw
KHGXJjkUrHV9X/nTcTa2oa9xqxR2SAuXvoAVJiz1GOrqobN/8pz1ZMCoq8hYMYDD
xRx5EkKsNB1EFecnIq/nTj/fwLizO9R1755G+uzke0mQ3IIc5EdJkKWW5bf0UPJ0
IAOfMXKIZx6INU5jedSMOQ2qxkRpGbE63RbgWAPS3MxGZMALZ17cSfVa3EXL4eWl
QRoV15KSKkCJOAledmo1FXvQqp9ZP5XHNFI2Q0cmn9Rcw1KLC9tjGL0jAZJQZJmm
rJvghEBaZ5o69rAvyNf/J3Tibg19vOa/LsAJ0ipCiEQ5n7fji5E2whXKe4/UeYzH
k3gplLDQeVk+4ciMcjIMEaDH4TiLR+muhuubc0f6IpMfvhJo8d+DLylmk1SPtuAR
UUjwkS7XLLuyeZC1rTnxYKFkvvwLkAuGMsjvbGzd5Sapvww9eqpLotHb97du6vcP
8GF9UWHHitzHg5OiXIVQJLq1pMH4YcMKFGROw7Emu3GvxXI38FUk38MZOIcEHS7s
lXiVbdTivDs0q0fFJnTDJZZ45RSRGtJEu21Xzd9LBLSDqzJC0wgFg9lpfzxVzjRU
+8j+fDIMi931Y8mvaOsVJgMgRCZTme7mUH7hVyXIpCdSaLF6q1AjYUvNeQ114yI/
WsbVkJlCMrST89AqxoPzhHStgyYSJ4da0yVLGkTY/wybFqaOOUJzuRY3RvwW/uvK
tccpuPG2FuF3LelH5e8O+UQ2uh0FnrecyljsAoCN9l6+xrQamJMdDm5tCOJ9JW4/
x4crwBmJAW21wsik4dFIAxrorlDyJBCSUMPXeUzSWfWoPkQEXUM0tT5Hke+8L9Ff
BqQzG9hjsIcCbI++uF/Henh47Weth20LLnFsfeNjuBV4q/RaFerPCdIwQ6itQVcC
9G46deOqJfYQpC/m9IYepBCIxtxuuB+Lf34QEyFh0Yxqz6sjqAOFoEGVCkvMzecv
OVpyVwFBHE3USnBMRboDceQSLkriKWKRrSx8TF+32jzw0mvXIQ2tjgayaAT3HMt7
2UDZNqenxDbaf+UH2aUXsWGxa4w7oDk385v2gsAYosQshk0WpBPAiKsALNVFRtx+
d7LtHP56r1vNM8SHDdzjPxFAVHsAwHp0FQ/eh13spj5Qy8Ol1wUln6smkEf1UnMn
aAK2QtRbaWi/PiNXTebCCeq4F+utENq2pUV7mdlh3+U4djqpnGMNALxCicYVVfso
na+8SGNw16xcZIwIuX2htTSz07fWDMwrEuehir8LE+9Jaw0Henhuuyyg+g+yTXuh
ed75JCcQGWfNezlbde+WZkC2lzdLD2tVszrUtmVDgChmDHmwBkVLGrnnxaaSBFDQ
j844T7qbx+BMNUFc8hGPh8nWSk5cyP5iy62ML0/OGlmgFA/xVVw9tnhypYblWJCp
Hi3Y57vCE/7rBuFarygHq3znXzfi8FWlOy6c1kqcdjDqrkKpe8XnxJ49TOF1dOqf
cbj4PfXIeXhchj0//R1zEqehv9x8FEkvjjYbuQFC/SuPG391pb4oFUARBPLwmsz3
HTKc8pmN7CteXYdHpOhrakQ8ApRiO2vcCm8rVsR6ofcRiobh+a7nxKZ0yilkQhOx
SJcR85LiSYZdep87cro9lHu/Uid6VssQjFtTzPz+cpnrhmhX8YWqcPWrYcl5C7Kl
qETzZdl04M2wUPcaDESX0ACID6DW3BFZ24/UKVbShKSx5Y1VTi61VoIa0Ej0Zt7q
WdUK0KJmTNH3q43rrr5uxCDlP+828vCvqt2giBJ5Y44oOyTqevihWwNFZ3FBzBLt
a6V2kF/g36Wtw0KhEmLNsuhIcJHtvrginhbQFkG7b+pmVAUuyu14dsVNxiyTD3KW
BDPQVNypm/3xCvrA2g3rH7MbAYBaSUYQJMrYmFQJaBJ++2LF7pLwKEvUKRVLf2D5
1V4eh7RNSd/PfoUEqqzbvtuufrlveePy9cwS7KFnFReOQmnoYvwebfNFsTXj1cgu
Q3Dlz7Dt5StJF9oge3vCG8ZCtIvkSnEVnY9+EQMK68+u2GoLfrSobrfYHSYS7PmX
ieWZO7roSFKJgmO0glzAo0MUNibsJidMNFf7Ka1JKWc4M36o3CUQzglw2ZbxV/SW
rDnppSVbrprqL+Ox8jHPVwL95oJ6hj3uVgv7dC7wtRA0ibgRdyZYF3BZQSKoLbBy
6g7zHG/sreWnb8R698LXzVBDnoAq7zWqwObld4Gp5OjNdQyjPVsg8VBJQz2/nb00
wMaoIB8QMrxIcek0pJX7KNQomBtlE20p/izeXnZNBS5w+8cxpq3fWFR5mocy0SJI
NZeEKRo2tSBKZi0FJOUf9hQXfcAl8vOlT5BNYne5UZu5wsMYx0CMzM8HROxsKIpn
zp0+SBryci9Y7juXSD5ko5k0aMzUFoaSdkxktllELQwwXappKgdlLqqe60ETu5h7
Hok3710dxV8c6/PN6UhmstAyWFD3L+IcmXEBmjm+O4vLsUBCXLwtbaKCu7GfuMw6
8pj+ULBIaWYpDRXUQcq1ji7Jv/apJzeOMh+vqVBoe+nSNYP35mCOTnyreI8hMx4f
lCU/pyntWwBh7sY+JEvbYwf47ZO7R+ZH8eG+/HRNQ+HQ92CrXy9zHN1FdPtSie72
/VIGKKetnGj0HbHZCHDgwwqW2/BLatj5c1nA7+q6/e0Pf55pXJp4+LDVEgPr6Z4V
w3E85ly+sFwPzw0fHfIVLQayArVCLFwFEck3JBXm2VBjGtXsBMBLiL4DJjHDRb9P
ljQdEnZM15QkD/KW1vASRQEpWaylDpL6O361+ykZLpOJMYRBvngHHGbX+H9nvAg4
ucVdZm9zsOsXym/zxMtL/Fc62CbNW6S+SQsiakcNLaPVoIcuJkdX5ZUNiD2zCH5K
AnV4yP59+IRo7fHpEzslYPP3p5h+WhSu8wxQjvc0BUiHMRvfFinK2mcMo/0FbwoU
Xs7TMG40EgDRJ+xaS3RXeYOjQTet28l8SmdGFLtNe8Yul16I5pewgjHLrm1XDi3u
uKFS5EQZN9JEZa+jaDffgROui0jCDvawCBgz4m7NgnxiUmbgR0R1mdQM3FBUd+gX
2nEKIGQw8S7Czue2uI4i4tZNnmBoEJwfn0TptIif27B0G8VfYS+uVLN+JF/pVRXc
vMnLvzfM2k+vFP6D4AU7Km1UV2MG/A82BqumpiIPovNNQcI6XDJCT8Ze2GBeJrrn
3+sWyLm8oomc+Pr+nGH5jsWiunJHl7FQ9ZE4jrRlIO66UvDeq0iwDDlLMFupTdGu
ADrE0Eql1yxQ03S+I1rRllciI0whiY69nhZy67efi60xjkhGc2el0ObqTkIJ8sLk
msQy8c0k8hGB5pCmb8QGfsSv37aVs4lcOIOvdopAeZW+AEYwQhMeaDGpM6iZ4f6J
up+0FQ4IGwQOttZ/gEqMF3V55x1uFykgb64Gb27xOJFttoNzxQovXRvhcm1vOg7d
CJEydD2ASBu1s1PBBjQ6sZG+wZwXFLtaHZ6g1gcLH5jhJBY2hsHOD//L92YPLcg2
OOE4cIEvtQDpf5w8oVumK77TSNFW8y7WZRo9umHIqJzOZrCRd2pnEcMBFhC99KAb
tdnYiJUMI2XhPhGTM5ndJLhXBwodjZssZCxquAfSyWUpAajlyjQ92U6IQb2GoE82
AzBhm69mLK25+HLHQp6CoKYXR13M45sNRLys/KTF1JWgJfyauxzDxXF4GRRWXoSh
OvRLHOsQFXhYjr22z2bnCpHWD8TIR2vwq2t3Hh71Rp4phqangxXgdB1q7Ed5YSNa
zA3d/o7n86KrDicHITwxgz3XcqkddmyDOb/g04FwVy6k9UKYCTmY9z8IaChqUssg
QimV9Z3f/tYmxXKrKYAazz5isMZS/8z5Sw2WUDwzkwmDT4Ez2c83mkMQ+UFvnM3s
Q9jE6g50nl9H7Glclu2DpCYj5GzwMQsYmDukzJBh3526uomOKE17ey1WpTk7JExC
vJF6rh0vKHZe2+X7tR26ggMsU24ZwM9rmzVQSXWQyYsHrpDdAqGx6xTuas4DKzLJ
KbVoJAOxeN3J2Gfi4niEdZphgN8UW56IUBSykjCuVwSD2oKpeovDeDHqMpaay3qj
VkdaSuPR0v+9TrZUZCeiE3B89QcyZ79FuRini8NjsenNHT3slkfurREK+4sUDUGD
HCNmIF+65oVpkb9MLSnL8/ZEJ2Hgei66kOvBF1ohL1vcqOLuAUwbE0oj2TewpNuQ
zocBxKLmJI9Z0U0lH8wx7lgq+HQQqVcmkdVG0T4sZQfV4HnGiO6GQH7cPgmZjpp4
5fhtGLZFYNJ31A2axqEqvg7OYqeCnBRVeYyIY4hchC3v86BF8a8WhGcHEPDj8ony
5vSubEyCm+YPqaaU93ZB3X3puSfgXhVumFjN27bAxZaOTg7HJXikxMHNTqJOfWO/
IdjI2E+5LFB6VUE8GGwivUwCBo+1MLuHjp4V8IbY0CqvbUj6bcWXVUEjd3JMK5l2
maB896g1AcXFGDYviVPu3ONt4AMa6LpQQG8yz6yS2meykOPrcYEiYWi5DYVxQDNE
IExiimuOeei4PGvbogN4ac3ChHVIFogI6zaDmkX+SPDwafdO1eafIRDX11xDxbZN
3L9/NPneRhtORzB7WztN0kGhhmZvkgydUZTGtYB2KYFiCzHz9oHKdmeUwoXZqMrN
wPTEsDFCnW/yEo3diX12zXFcaWXw/QtsOCiBqkefbgtH2J65MAiuj4uexSV2Bz3D
R8+J6MTW58o4ZJpv7iusCGjlsjvswSVVF6zC3tSDDTm6ATjz1VnMpuDrZ/yeMyVj
T8+SG6WeYtGvbnYjsx4V3HRSeJNsVVP+PNoOQlVl6UUrnC+p5Ps2kZYk2Gmf5l+T
53Nc8LlymSQEavZWYvWt13MWw20YHZmjYYUOUaMAJ4HO91aH5jTRzW103LlytSVM
LDptKqM7BWIIWXEWyy5MOZ877vZb4zxBGCLKwVRMCSjqt/jkhIp20yp9yESRbPq0
vO6u84DPs8RknQCmeB+oK+tCxaHRQIMdrvzfONx0mS7j4fZl6cmPDqdNO44kOtip
937BR2xg3n5Z8SkFzNKm4AzLTFRLFDY3A210FluMQ/1UmIfv60+vaJbeRi5vxkAo
uVvX7DuoZ1RDxK/KTA+ab73avFfRrVakijL2roEQWXkOmefehbb58TKDhFXAKPh8
PKjIIlP83ZRC/mISbNkO8RBfZQ00doae1zO1euq4CFGeO4trdi+FRU+2gJlyhbzI
NnXeW4mqXb1JpYV3taqkiqgaRpv++zi68qTrVYZEddXHA1GYAYK8D0GT4prDvAsY
UUKXpgeZvI7+Oud0wpzwpUlKqGD3dG7sxjHm9qF4l0qGCua/8LmlxqbTdZpvN8r6
FstaFgD4KImyDrY+R1oZfdJtnQK5vLnQ72/T3/P+/evS9UnMtacsIl7wG41cbiJA
OcK9NDNZJvjCw+4y31IygdOr2jK0DqYanre7GkMI36bZt65Zb+C9Akg8GzjREWYF
JVrlSOegXTzL3KoPvbKXupFcVzDQXs43UxttIGC3I5xbLVvNTKjxcXN+gsLZpioV
a+AgrkWtOY3DlF/AhZu02w7cIkCsXVupOM7A4AlQXML6DjGs4JSaj3mLRabXm61+
dFVfN+Ng9JlqpFdq0eNG5zFGJ44bHPI2uU2bSMV4pm+fQTKLUMMMls9UJugQTMc+
3ZZdbeZ+L3uFsfy2DfszDAl4fOUWsVup3f3jTukHuKMDesbb0+sphZSDA9MOLJAU
v1lRnL/qhSynOqFFki47tx+odMKoSruqEyo5rbAXHitMaz5JCRZqs/S7VN7bzIy/
iJQUzilCE45nWsI+K8wqh4kW+xkugOfXuOE8OtpbIlac9/8seH1mHh8P0G1v/vnI
zvWY/VF2K8KJPX8LQVDiOoksbVQtfdWPOrv1D0z4H3Gdn8bZP9szAhpgd0RDsxBw
E6TBqPb/gttmR3Z3SH5VEceBgZyzV/ZqelUlTw8wxEg/CvCVhfjvD/Krn/AQjs2G
kXBuUkWnz2PDhah7Z8hikNfRFZkxrpRZHFZ2yunHIm2/X7Tku5RgK6c+vCzfPqge
+Oc5tWI6I0eF1cwxXvlUDuuFUsX0k3XlQMYt5wXzCcW6/R6Mr6wAs/W8aLul2UUg
9HUh1HhZfojOrl/gHWyYkRDAXmapYeUv9MSYpezNKWgRG8DzQ4DKNHMmhrrohChk
1X4T/COg2lh4luIxa4W/N5u5VEPTHL8/pG5XGoX2/DVuSS5aERWl4p42Runs85fC
cTZOZ9xKuuMWU2rcuQp94ATFqvkX/nOAuifri4Q0mMnt0uzbsyPA59wYH1qwDT1N
QxTGXgPPFhNwmG0YW4UfSaVPElnw086jLy8fhzAe86ifMWG0mXYR71m+E8Wy+bwh
7falyd1LxlplDVRS7zXm5+28RBuRGZNFH94IPOaRcXslnNVTeOACOTh2eG1xjouF
gVVlGIZCeSXSNicgnXNQl9YTe3NNR0iQ0KapvyHWSlIY92upmxDNZakHjHZSuElq
XMGk3v5TI0wOJEqfolNQl5fkPQbNY0zGUX2+zMUCY79o0syTg3Hq7pFj5B2PFYm6
KlcjYz5qB/kUqAnU893yOh7GmL1Ksijl+OpzXvlKkYgHZmd6Fig//OZQNpoUIUKU
QpDEANL9SfzNWYPYgqO2WewYxLwbJRx+g0YuTxyl6Zu9uALA//kQuCqaAu35S7Vs
POCjNy9w32fk/3yI4l9creztJ/LvhBwRhuSBpP2RlaT0aaW/3cmwbxo0G7h1xl3C
giVxMk/UG4vPtYR810uURYCr24D4cVb18+q5RCW0+CRlV9e0YTE302L3HfOJbCRc
t4el0ZexEzWeq2LikYgcoBA6vUxOFSPEhJrKPDdZetipoaplZGolcyhdcOqBefW5
Psc1N4gu18GW3fjpAZc5JK6/NIerpCCh7pvIoG2sfJvX78BYsio/IYtJYIvpEsHX
ibUQZ8uJa8LBJeHpBukR7H4S5ysg038aJEqHu+D1LTz4fPPNC2HV79HGw6axNA+8
QvT+g/7hgVzMD4ZpjWro6G1ZUjsM+y0Foo2PnCrbujf4wLiQ/PlwiBHtCr7BpDRC
MS6nHn+QDyvDSpg1/tcrmEWBnQnynWc/mzbw4CmmlC8y4U2qXT4Nh4IctOhls5Ab
9EOh4rgaZmrihir0aBmZEDM8/jenvBQ4rS4YqLzI2QKE/WoS+LChVPaQFdkbJk2O
iUmI0fZ7YgtDs5RVnrYiQywfDK462cJ0vcu42Nq0fqYXQlGmDed8E3rm9R6RnI0y
SPmKAduf60KzotO/HaCDOL1HtlgbGSpNdaoVc5aS110JST5HJyghg2fwcsSopiN/
Hefeg229z6jVkbpyJBJldfK8FOPolbcvLARAgB4nmrSoG4KcNRu+3sWAyq3owk2h
wpPryGd4MsMWVTi+hoPAqa1AX8h7fmi5H0vol6tNTejKNB4NkQMBDm3Yk7vpBYfE
poKXC5PyGgOWbgLVZUpjeoTGrNoSh0zM23pG820+8rtWJ+6c6a+6S+Wsnkps+d0B
pC2coEQcZ9JNnI04KNtJeEnxI/kJyhcNbnzoLV6xWQUOxSm14R9ArQa3gLmI2WyY
egYQLZtLeqeub75dciD6pP88ZGpF8UV9M3ZTH5dFCGvDN9cz9byayydRJTxXXoeU
TTq/bXsH+DfjbsN3XXkS83YQIviE5tVkt+vGRExKv+5PwB43wRKeHbRZScK3FnIn
68/NGRxbpC3Qv7oxiD378FSwCEUlSiw/Dhm7CYsk3MelEHcvI//N7GjjInwQPsh5
5G6M2PV98DduJGEJSmvYRsAp9lbnGCf+vjgA8A0OQHmYUb2jfsdKLaD/jmNca15P
84/rQRgcOSnqZwlioxpZJWbdI3+SfTAgPsNkekHnZznHJOkbG224kcfpF0ansWlh
9uYUUQ74U7SxmjOwdykua2WRTqxL7Hc/RQgw8+HzXuY1AK5wYqcrHZjWTEo89gpz
vxfMwq0k58ZWJa7bm+PPbhVUHUzLtawBh0NEgI9ImVzc4RnPGVYEiq8jfWMdFaMr
+NmmqU3//aCLyggByR1JeTXSGQsHzONOvNfVnm2ng9YhXvjykbz4DUdY5xxyv1vd
YXK2GcHsXXFr5GaGOfKNuUuFbvfotHSofsrM7h+QFCGnKEP125q2Uq08g9HJ7N5y
QOvHLWfDYKmczedqsYVzPvOePkfFQdnTJSOIaG2JwJlQHPOsbw9qYzfjP1naWBWd
hMyKZnVgyfIQOukh2VicLUnLDKnrMFabMCez23xDrlZb3CSBfeaCsaMA633vJeL+
T+dDQ41VnXViZ9fr03g6NYVGLl7avsH9DVvYKpT1cuZssU68FC0hZzey7d2jqqgk
cm0C13VK81bRXSk0aLHcVbHBIyleQAQTHUT/4WfkP8HMCRb4wg5w36qMXpvqqi4D
uGEO0q5/DJ73m2qSKYMAOvn2TM0SiAy28fk340QodgUeH4cvsUnI1BUgxF50xs/V
09sEFf8MZkFKkkupusUnZaWD7LdYvLmuha751aXhDR0mUGccY+IvDGQpvrPJ4g+2
frxunN2MCm0dNS6kS7/yVLPF9XWxcukR5gplPArua47aRhhJ0FGGxoTt2grqr+t+
gR7vjZ4KYQiSWpTIH1ThLTo8/F+SdsvWxk0ob5xfMag8PtvRMCqItZjX4RSdOEqf
bvPu1DdXZO2bCMfN/Mjl+XziDhwb5Mf11xaQMGhy5uAzWONKfopQ5k7xl5pQu4oq
bjtpLmsY7AolIZSWFTstrsQZ5sIavBM5gbW/+7wzHfsSy+l1cNqzSBdrsthl4ffD
OSPLk/wFZtaPdVzbdiOg7pqhLMd5WCqzBZM9gEVY+oJSkseMafxwWK2iVSzDsv+o
kpHEqQ5eWbGUBznrZzu9panki7lmYObv7sXKAkyEq7tcZwzK7/Hn9XqFYTkQVeJH
6qohphWD2CrwcwoMNpDRFKuoA9qVLOU4kf66qIHdD+Mz+2l7tHrCRWvtOga4Qf7N
5mDFrNZ4jGGC6ZhPtW9vQxYL/v+HYJ2H3tdxkYmCnFIxFk1LkRZA0J9U1BBa3qox
tQxBGMtqXAH+CkOjtgm51TuizuKU2ZbaiIHYbgho2Xc7BCkx8X1uFFw+wH9IsKRq
9BzWTuiQEmEfHNZOqYvdeTDl0b95mja+ufHSU/v+YLyIlUGo8D6j31Ssed029QFV
1ulIr7R46n/bBDhJAEx7wA8KJYDRUkC7nLqELWLmrcnksbZBomjdxIuwYUi4pACP
Z/kqqa59acx6kJwlEzcXJ76xDPfl8MLusBEtusKQVIdkDcyL1T1b2Jf4uXku38ij
DiPBUXNuRz277/WWTE7+kOWBRguK/zYwu2Bf9KHr+dkeicUe6r7YgcmZteBg37jV
loLd73fieIX76bGC4FfVaERR12rYiaeA5FJLP3m+VHBiJGJnXaSfXfwZ5JBuKy2q
VfC4sbX9gh8v6bKxTa/l8+DvyE9LW08o5K+tPUS7gBeNigb2c3nd3fzGc1j4zdeH
yeZcWJ1ozTj8DIfuQjQVBEnBHYpf5lQmXjojYE3mi3plUdnJTt3leVsvx2FcWX9c
UR8hOqs8rCYKiPOlxRJnYQQ18RKNIPVhP4IISLSt3akq7EJMHhOQRFh5VeRscQ+P
0Z5TF3KtXSV38wsiFdevyyPPaEAlW9grvKkQWDm/YQiyxCZTvWsrQB5GuMXAUAWq
tiucyIX509luO2BN8WZ67R/sXYth+NTF5ypAQ3IHlzSHdn3Ob1Pgppa8kxzZhdHT
9u2lTFn+hNUvoel7JNnXfqVMTzgsQhyzWQlfFgK4JC21S8R9K5bxeCZKDYm2HHAw
spWD/2Adi+xfMCREvnHU380BjvdcH4Gdw7XYJEkojzNrG2VJ6OvlUEY09SCd7W41
wQN9jtqJWiCVANnBViu5Cp5khgeoyapILtNmQgtiz2xxls95CHIbzoy2c53wexVI
C1YJCeTjNBjXeJ+ZYt+tPnKcLMiA32sdQSHQAbbvlelu9Ty5sGkPo0+awCQjyusH
UjFVFQnFGwJ4ei+XU2k5BPoUo4mG1//Vq/o+0TFuqw75S6W1WsQPFyXSFodA50NX
7t9xcYmsKIbfKwCZXIvgMqxF2MN6smvm2s6UdUioDJps4tkYohMesFPt6v1TF/G2
YrGJFBj1x0u7seOWntVAZ5A/QDSdAnak6P2LnD/3lHK6yoCLf7uLJKLLrKt+STIa
lzv13zq0D8svQxmVXlM4WSvno0NrhGiVIN0/VZUWtCyQTDik2+Lgma8H6z8goEwC
9YYWCHLQHUj2Y7G/bG9K836aUxCUbxzStfL9blRzCYGtE1vtqS7yWxqTJQDCvU7h
FtLTjXVt9EWX/qpkNSZ9hEUJ8UjRvy56M+jYA53vh9p4fqp6NJk3ijWAgjxSF6pz
NDwZ6YGWQqPo+YwrvkwJU9L/iv8Bi/AaV01cmU43MyjaaZVwIoz7ZMMSDauGiETx
Bgw2T3ViZUh7DmxbXzQJzqkANPd+U/6Mg7UBvQzoCYhhojwfvDuAYBjkSfvNcVIw
HC6GSeO2Mjp94d44nbExF3mMbgWHgHkBYVqzBRDZH5oyRIuc9X+vB6MMIxVRSmYg
eKai9sh1oQk41pOBeXyUT0ujatoDsLP8cb/xH/sNjv4M0lHJk27TqFLXlD3aqB8w
nUTOxi+ITOlQ4Nkm/qKWD5YHbaQjS42hQwa4koc9N68tBz6UZ0/s2+at2vBfG7Iv
jXoQxoGE4diQD4iiRS3GYoWxfSm30H/OSCeBgy4D5KbWVv7s8kV5/PyP08wD45Oz
wKkbYWbkOpKkgfveR5gOJ0xBwlBaI0Vo2EXflx3LhUzgvhVQwIA6Pt6HRLTBvHHu
AM3yTjG6EjEem13vPFSi/NsDoQn+BYVT96tTpYMxO3idkxihETQNzwHLg/iQBH+d
L3sZ5rCFzb+aU5iVtb76nMvkVYsyW23BsnbkL4U5m1uc8d9YMip4yQj7HlOF2WgG
Mg3qzkSo5Tb4JyxR/uBR+6Kgmyozf9g27/V8hbDSaFBh8fRX6FrAIweAb6bYJk9F
xBXZRimKF7alStZUrPuyW6embFygUOGAL/GqLAxMjJqlqbufi0kkd8XCgWN5d5FO
lAfaCC7Qkhl8AhZ3hPyH+yg/Fi7haVJgtf1ptiYdkjbsccrROTOj7ZaP5sxxo9e+
wC1jcKeCR7NjPQBOku6SiLk74hCRKJpmkW5fUm4TcFffeKeJN010TR2m9JwVt0bk
+zY3FYYYEKnNe0ehEeCgkHEODzgafBorsEbd8HjaUfAdzcOxR0dt+hf32NRpOhb9
6bFUdVcoLS7tj10bCyNcvyaVnU9+Lymmm+xIPTsNjxQ3D2aGrJ/H/xfTTrG9wbFT
Q7F5yBzvvJ/PWHyZfA0d/Au45oPoI98YUQGzAEhlXeubctqACWeyE0oNi9lMGVMO
vUEM70bMEJ6MARD3y5BY15JUoOD1vRR5/3CXOSOqE7PffGjER4KmxABwhL/jPGXS
Ow5gj+hbcaZSyC76sm/XY0T+PPPWJzIAdr1USSDdB3+loV8kN62gEhQuGnsR2Na6
1Loqcv7myKVfmC3Qtb/lVmryN5l2dP+i0lDgklnFq7oQSJw+3CyX639hEwwXeFD6
S6nyibIZyyOZgQsTjz6arqPlk+Rck7z2hMcxsZkd7w9SjRyb4yKn3TWSlFisJjjb
rBZ3S63Ih17n2Jit6/nY4u+AdZEf6mne2rnzWvTI/luH5ta65XFB2SwYbdoMC2AG
8154QmF+Ob3nWWmD+jOHYXR/mVWDaZZE2ke13xKmCEsTANfwoLDKSYNINgyako7f
+SoVKtWT8s1G4G3FvYPR+2wReB3amqzIPKrzwRtep4amURzOvCAT1bZYptjWB21G
IHxaX24IOcb/xtH9nlwEv748UmeftZFKJ733hsdwRdsYbDu/a6MRymP1BTq6GlFw
xH0k91DDA8TAsO9sr4cE+pj1DH5yWy/0cKpVs3crISQCp47L17VnSbg0FtoA5P7U
Ul41S1sJsccwbR0STlE9FiM/xI9jmX141i6S9RIT9DBY0vCPeqOnuZ6GeiT8GhYs
mqyJAseizFMZNGoBvLW+JbXRSRFr9wgmpXmsmySU0qOxe+A90dH8TML1defRf8Kk
4xP5cDxAgOkFZQECoO9INxDH+htEEF3WHvrJ/3IeEtaUsabNNzPbYcSkT1qJd+EZ
Uqpry4QeFWMkCDohoAbQ+A1cotYH6PRJjYxYB/S8spZeMOBGUBpj/pOYw2RnpEbR
SuyfiFeHL89CVV91GaBVjoGQ6JT4hccY2I0Wwh+qf+DjKiTzzliJ1J6n9croTAb0
Qf7MN2R1IIBUPZ+emNNJWu9Eb6RxjIW96dzHvHDXBgbVHeNAVy6qse77h1BFVWzh
OhQdZJQOaXOOVjYst22Fv1Rk3N0jNm3wqlaGI7wi5g9KNE7maKRBl+0HoyW69/4u
CnxF/TIjtrbRRwa7FIZkuf3Qf5QZU1BooVLsNEbpb+AV0wyNCfasyOXupiEcQfn0
Ack+931ngWcwk8wxOrkPmdirv2ydbgQF49+FCA0urG3HwsaQImNWRU2Fc7VdbRzf
hBmXaJEJvKyevLUe9PUQvlPU7CsPuSpgXynWDiPO35AR9ayS46bslwhxhvU2SvIV
fdFgi5JODS1VtLjY7zsZWZ3L7EkBGrJHOZ4o4y8qRyA1j8QxeKki5pMrxAbgunVz
7byQ2hVEfV+Yh5Sz/fXscsMp0g3eP+OAe9k30Je9hcFw+NS/EObLgxWpGT+BbvIx
em1xW+PZ2wrwelIXmBs/odMaC1zo8zKi0OGbJkqEXMyI7dG/SWEdAYuzYsVAuLMV
1e6iqVIo38r2VGUY3UQEsDBZUw0gfsBoFPxks4TZAylgkZovmP3oN901YY4y43ER
ATDfrL/pilqdVb2Nhv7iC6RDJL7WwbiWhGfhXglBMTfcI6xqV1N4QKbLLxLOCF5b
zU4gJlnLJYjwyLe/GUvnLc/vvCSiSDrmELMDAPnuI4s9a6wgbavS81sfM8WLDXF4
xMyD3vfHNLEmL/Mf8KodkskJTU9e6GR3i9YdVPDXRyAcv8e3JQtd7zM06VfBBQWH
UhnpznIy9UvfxPlmCBw1kNamitrT43RYFN0jdzeLsIIcuNT1HMbzDt7UM0OvYzcD
eFes57diP9ENQjwgeRFc5dU5Uza51WGdT60lM4DeWIfXUgd2bygmSyNnyw02XiRT
UVrUF4eeBr8D4/7jzCAAojJtiPoTas7IhyiNq4wve7QnMVttjbg5Ty4M4Xo1GMev
mfR4BbD1li7/mKZuKh41WAkYY6O2OqrOw1hXgeIGGIanIwdpO2f/kk3gBWvdzHnI
U7WNZ6rzqViQpb5bSkfVSdfPJQgGIBqsAtY5Qp0j5MWsF1Q0GQsDxQ2pPjSPwwCX
ZKA3hOUN4M3m4iojKVyzAmfNLwHo88zaGv7xORxrfklVKLPBsEqwBWqJWzkwPAl1
NEN9fG8uAGiGaRVWyV8ExVIx/KBd7LszvUtJiUB0H9SVz6HcZ+pDd3fX3UF1bzyX
E2DuACqIqb/RWiHW97IxLJGtOKlU3aGV5ja/adsK3cbTDLtRA/3MEk7DdLld0SJj
7iT0jodH06/gub66g3pRsmQCz8jEwHDIUo7+g2EZ7QsOC48nrLOqQRXwceKEo4XG
euzwAUC7ieJUUjugN62mfgU4ouhsldTm0jJ11vUAiiSBIu5qX8ZlJksQiyG85eSx
C87CI8zuk3DOYuoqzy/mBUQeUy/1qK1DzV+z58tOYPJhdMpNS0VMAN4yycREsk5y
tm6RS+oF3ahxTEsqD62N87/E20jZ9qF1+RWwAM+EEc3A1YT9QxGSd5oWAV2KZO1P
MgwS3XTwcufkXGSmrXIUcIuKm8VObCJzfBHWsDUcWlKemomkpwoY4D3IUTyZDlNw
1xYKhw/KCQEC5cXr9PqllNAYTm/z/MTNAnXt7Xxx/s8VEyjO5AhYduumfp1PQo3r
pzhwY6BPXQLk4+Xz0wXsv2b64InOww8WsT2TGIN1fiB2vg5SFsyCAxTgtZPWm9WF
7MEqEwJCTt7JMYZCO585M4LR9aRX+4NC7kxMNl6Y84VR/zz143fcuyQoofOF4VDn
IKJMq8K5Xn+9FmN/CaEjL2+pB+spXOvA7TzkvbSKSpx+08c0QLYwcX0P2RriWV+d
BQl8WLuSzdfsMu0RGskv6d0W6a1zvNy5+Ny9+3LcNWmRbccMgCA6rtLZS7SAf4GA
PK4ZmbnNVBBAeuwKh7ywfXS5GDVQKQvvS2Q0JyLPevVh++dTfBPDqkuAnJdJ5Cjd
Ky58PekC+AloUJ5Zu7JH1A1FdHijwSXYCZIw1OoXH8vpMcHgLmt2sZ5xkGfKle1o
3Mkr1KDQewzJIW8NuD6HAhcHskNCEjzPu1ayM0Nf4KnEXpCA7RNDeSU4r+2aLDa9
YBXOay3dJfKcrUzG5RwGpxLmNY8bhSuXckqJBZI72GmpsUtInAVUFFBbbmo34Wvm
fgusfej7/FvxgL0wslsBV2zNYjp/UCULvUFYZu4f5LIC7XQn6UxkfBDyPvg/mJ0m
ZihZ4vuJfOVKRSVSg5gcOeLOQQiIgmnzaguLY49aVaAl8p6FsOtZTXhmL9XHnUrM
esUMPHGRIQfu7tkLr3xIN8dBgnaFLF9C9CUpLk02e/faeFqKJusW3FTZ5KsPDTyr
/8PMIHGYLc88yABlKfKtjuAvBWcgUXKnpELJY1MBZKWEyNpbQiXCag3gTz+ITFyG
BTblrbyjgFyx2aN94a+gViGR0G3CmN1lnUNwHfdssHFj5vVh/NhpwSBzjJijDu95
PzZ55a/w6r5Q9Qng3zbcp0/7GR2avQq5VsiwxDm2PRayJW/oItBV0LidlGZETo4a
2tZHDOwr7tWqHUbih7WCQZRXOAzfYLUuEnjGCRkhqGlrm1+3miAY28pipE8goSWh
+zvEhegjiDAA//uhajgGKneIjJvIYUlWDn120PmVkEhwPauDsuBm+7oAOgF1Grek
ZTsGryCUY/27n5XtDJ/lAjoxlLtBTTR5CP3UlFCShO8EN6gzW0xxc0gs9aT6JMPs
H6bdK2cUiU9vQibgQk6EvRCw24AgCtJSysMf62nv33b8fEC9XS5Bh0LRSCHXtlwM
2ygzjv5mNebvhyBV03Fr5xhPCS7eN4ia2VmQxBod/29Tt/kdvZXaEeRCwSmOfom5
VL6hffqSUQgpeyBDCW6Gz1eBG7VV1YxgE6+rAp3ASg5hc0J0l1fOcp2ww8MAQGEC
LZa6s5ipwInd7iXGTlF2/b2e7DgGSB83op4kU5+g3ukz3Q3ODLuhG3VJgPppF/Wq
/SVnHvPp6lbVQh9hJD+okAgP1IAnC+DPvbzrVEg5JraaunFwxlWC0EXSEQEStnTs
QwijvaXoZBs1J/1VUKuVJV9xc09Ism3AgIEYEZNcwjTxv+bWuKgf/yCrhVxdXtJ8
d2YCYbWqVCUJ2meVmoxzmhyMn71DBTStWUjIhGfYHEwKslkxuVZ3tmr7j/FEGYoN
QI7I4lB42WsODHkQGyWWgMAbcGaORTsrBm8eae2zXzg90oW99WihQ2gVrXX40lIo
iUpyl77aPa0eUTNElhxkinijYmVLcwoUH+TBTQt3OsDuGL/kZfpGZ5ZnQEgc8wnN
6dgJbC6agl1XstLVsqNaIgugP/t82i74avFmqkbZ3KCMnTmLFNFUo326TER8n4Nn
LPhnwTrHTuppXzeWKn8wirnnZMOa7CuSBxtxjFNPonD3D5mjhXJ8dw/gdadMDbIG
/tvvSz8Hyl38IYrKo7/wYFghRoX/fNuoZ1olhPVW6HTYfZ2u40UKfThSJZEFQUMa
mMZ2j3gUFEuwt/9WX9z3e7xf4eGice0gUp0mWuJegQHpH2RJCBOFNi04JGp7olDs
TmdSDUpGdYgRpYw8M1gGVgWgrnRiYtXC2k9Xvb6ZXxaDmvIoWQtncdbAa7DUtZCw
50JKAH8hzeGWRVQ9nqenBORdk6NpCf90CaGav5/BwWDbRD7EbPQe52iOxlHxsC2M
neIV898OHYyOyBiF3j5vDmwAF77Pu+60MweOnv3CPbf4AKjdtUxa9d1GCgX2lOx+
FKQTa6DvGyKSRJCEHqaMg+xjGi4/S8BmwsW/6kK0UBWs/RHh1pUlDXe4Wz8WNDIV
5gK9JKiK85zrZrtdt7H/6YawDBAW+Lv0EUn03w0hTW8QyX3QlyZqGPiBE3dSn6Wc
/cJ21ZrYfh7T8bWICCpBDI7bHS+2sAtYOhmG3vvC7C26Yx+2KBbGOq5h6J357o++
lVx1A4sGxjAeYsNm+imEHC0IAHQq/dV45bU+GaDnEceIBLWbGnlrQjpMhNHqf7Na
XvWZx0qjZW7RXyGHSEeCX8HUau6lvQCUkz0a7oPxGJbdKHl06O1y8N5oR9N8OBuK
MMIGeFcwiX5DcZxZ3I32RtXOsjzN8nQVg4ugeSWdYLiuTIbzdOwNqXthTEzg+Cps
aZQRAuZlj5rnDjgD5nvghzdv7SIwQgOGUwMA6r6ZPqF3pKu9zswmcaYliNcl5R12
02QeUoEhsq2VvodkzPH7veKnmsdMnFgqBchRuiyEGS4RcrrsdJQ3e6lVJjptyewZ
Rj+iOYcuPjh1HxnEiC/eSyDcRSTcd/sKdG6iHGNoRwbpwpfxov41TbQkHOOJzcsc
HA3anfSa394PPUS3L5sVYhs1cyTijOBF33EkOs9ERFIdWBFLeQiI0y2lBPT2eepk
pYv9nskCYZlbN4K1DcLSmpbcrsbdsZJjRwVQLuPa0c9I8SouhInMxZix+lWudo3i
BqrXh24hDcVoQgAYh8ICrwM5FfmuZ8BV01tsKTqC/7hDpLaGqBHYy0zdc0zkjCFa
h0IJofxGw7inakKP2SU3pjYpJIKohqlVwNbSo1wsA872Y/jGUy/WXHJYtTaejyKN
1Z5flUsa3yUUy9GMNr24jwKahH1pVxXA2fE6lSsZ2mG5FFaR4PsVjwArt1abzN2A
nYLqrq4VACqev5ravwEPg6M+V4GT92tpJjC7utzbY+m31yGUKiXmv8/SXcF6L6Zj
MR5Y8iQP6oeWJhaQC+Sv2HOHJ74MLKJKXxVhBlSOYmisVmPBc6L19aZLJAJY4inT
2ayGldUYfkHD+y2nGL7FFuizv1zGG3Vz3FT8mqBzKHoKQt2e43tTBWEaJK+khNYY
v8iqGqjp+iYX0Yz2J38qGCXQGwrQC1Yf2JnJYHN/tzXmzONWhiZ478+4nhmnVW1X
ZeFBYdmfYbop+i/Bq/RJzL62wQpM0ISWdcPVDGntQgOVL86t3a6ZFRgJFcN16/A5
i/55I5xiA33XclHMzOqgBGK++omuvHhTSYfyTrI5G3Ypf7BPtq9Gzbjusmh/Kv22
p1JPm61FwbRSHUqtQBUwWDYGJvJ/xpotU5sDl8HdxDKpzqEas84/ZZiWHnnv8wvW
9NvQI4EgTCdTkT2Q+gjn3teyfizGh7p3sDkzXlutAfUyEPpJBjMb0Iv8Laam8n5N
3QO2PzmhI7N/4DCQErO1/lIGnbuoAoZgOQeiahyIGE3jeXvQVrKuQ0phRI8em0iO
62lp3k5Hg0bEKQ+jezJGWhL8OpDJh97RRGLg1nCDJYdzMOt1hnbVsMv2ecGf9k+z
ctmmJcts09eH68srzSjEKTYqZq7dc3e0AxfJO2UsY8X15MtgpVimbXpJYq37Uk5I
s1yIZ+diFcJxYeEzQ/toOdCP2GcSwqFYTvGLOTV1So4x0ulpmyVcODTqE8AUVy6H
EHfz4nVUpWqicsz1gHjQ2zgGk+53YaMVm52pQIwdGBEgrLQN3LpOkkP4+mWHAvPF
x+ZVyzcPUCoXI/QQGDHRiZloDbUvuPwb0zKu3NvJJ59M3NFvrtP5SkevDZRcCfuW
OtXegvNYtruoaK/hL/j9V3A/F9EcuAwkjXjHqjfB+kdkza+uv2jhENfoU6gLRQHp
NRLvexqw/aVZwxr83lXM6WlzfQ4Vgft1ytW8zLmKpoaD48Awzo63mBAwFrUVynn6
04u6DbZxfMcptVk4jm5AE1oOcZhg/7XPq4kE8QJNGrjyGolzEyMmTVbjwec0ZYrv
ZyftYfBVM3fQfJI265ho63d9yxPfRBL4PKJW9aJjr0TrkP5PgGxZpLGXFNBKkzSC
POVtpSlmdujT93XHkKcLUbmeKF1xKY9jLsO+LrY1BfxVYiTHA+lMYRjD3fKiZsMB
leUxQySVB/Mv11J5DRNWnDaNyto9mJPRNmQtuODqYsgEIALa2Wt4/6UUy1BqYGUL
56jYv9fTDDIOLUHKAFags0+uMRPBeThd80vs0SRhHC37hRuYmaK8W1LcB8UFKzsb
inRZ02muQPiZ1tktwuo/sgOW0sChqL/kyij1KtBhQh9QPCwk/ORJAPRUckjweyXo
uLFykPwDYBt+eEPt50pc6+4mjES488PR+k1JEz9DEb8BpIHyQCid5MH5fflWX4U8
/IjSGDhBSInozBoLz/Fi6dS53HftLQSQKas6YyVFV2PTBl6dq/kjlZyBFodKukdL
YMHDGxGBiFCBGyt0K1Vrj8dZcoFLuHXwadGOEf4DSfKDRtO9iKisu+/uCM6kWAPC
0VjjnflcX+tPmVesRKCYZ85810/ezFhJhXnwWz0Y0fL+882PT9BrPjhHsa7EI41k
xMZPbVh/ZuUyRH/uy58gGiVWaiYgSHnld9IPoLVqW4CqyvqVQfB4lTcHsoRRg9+v
swuIy6eAzueDGYqyg2CSqsVF5+9D6RB8+mcaIgAd1D/1KXvrF28q4FsEKm1ZMTxY
FMSfjSxn8qj3wEnrtngC+yfKik2md/A+wxxF09eSN+GP8QwKmJ96VMMKfS0qLRfL
OuTQGQtAdlRkO7jI1vJ1ftDSdyBao/8r4XMHZoVb3VYbAfmhjf5CLQNVB/1a1b76
PQdVExaNz2M5NDpbDhJCMSUzXuBzoX3KN0pL8d5lHB+EZH33lPZPe8QzulnNBEp1
sW+DaPEQj9oLdfonCJMvQK16IDhqRQxubaE20S6RuJQVax1Kmlko7hYv7BaRdROo
MMddYgZB6MZz6p3nQJIQwj8aALIvY+Vd7rXcz8s3SKr4fJPWzEd4Isv8N6wwKlVa
HZ5VEt7+r3LuVaZuglMEj5ZVCIbx+7vlsvQm/kgKK41DLANV5J6POFFGUBfADSTF
u3xMEusok8RedxO6VerJ26py+a1kiV/Si4mXC8049rvI0t/LjjhrN34G9Tnn4yfN
DtMljrZnpfJwJO+npTzAORAA5Etb1MmWvAIXzYaOlAK6qvBNyeDfYZTsJoOsSYcd
7nP16/81aaJztCmhSSXziDZx7p7LXIcgA9HzOGSFVTxHtW3AUsV42R+rt9ePRtet
LqrLVNvTtG4T5uGc0iWhNvbEJxaHxdD5TNaG8rLHvnfsaLrBPpGGnaD07Rw3tQj9
D/mdwCahG3kZd9PSfqj05oj9P02IZnrVJrjyIrgWyNxp0e10coJCbPNTH5yxzCc/
4r+GFdbzKkrhQ2Aa0p3MgcQRJFlkUJ0j/HkvaglJ+YLnMdPqLuWM0dezbiBu2jU0
DL2NKrMrTro1Ch/KayddVprcQNt60JHy4mHa+P5BfscYRIi+4GVwiA8GZ27KnV0K
VPF1d/KGZcOIX+/brDGfOwsdTJoRF+0U0HmW2AEBdMmOc/sg1JLq9kUP2dFrcnMu
Ht2m7PBI695nJBNRnm8U6sqxJ8ZfCC9j8osc0spdmPSJFB84jFb3Bw0qXWiuTmCY
tFbsgYbLKsQKS9HlV8LszI/8jCsKUECAOFPDxErZdIUhl5v1hWlwFtb7vURBr3ID
eJ5KTKS6/CPXEs3SuI5SB+NjEvq/YkzdssU00Mzw345pZQg9v0C+SU97daG/Lx/z
Za8O416YlCR7BIcRZpjwjutEnh/eBDGkR2I/zOYguV9D8QD6oOx6v4PGejL4jTIA
wHPRxXpMHK171fYXdV/WENqGHYFq8iVkhNCsdZ9ykU8+khC6hDVZSwVdeVlfKsOO
KTn516iHnkhB3r9YbX88t9/cMYufngeGib0woBGZ8Sd93sPt6203m+sVWB+nzv5X
AIQ9Jhu9BdnG+Ex8lvGqCRG7u5tgLnFiKdSuAODigMOma1gWndb60rvwLPIZPwzS
AyLRH7VaA7nyM3eDOHzqfYLPVSCsj3J7BvIQevIpvlFhtE7TqL5gZ/nrN8H8LypI
ycXYgpD4ZO1uVnKxF4ft38pyklEcASbLn5nVl0ZpuMDc+y51VrOw0kkkhPayEXXJ
WrmL9smkG4El4ZXrLITB45tCB3jYqp0TCJaDeJKy3eTV3SiJGbBzaI/DE1iWljd+
l65V4Q6ftoE3OuH/GgsItdNxeTQ9+U+geQa60WePv7lwtyebcjd1tZAvXD8UlE3W
397ck1ZaS8MjgpNxqU/OdqMm7IB/bRdrxOEWIuGH/M/fw4SVfB7X3MHSqu59nDKq
3mFQMxQV8xf2WWEF/hdQD6hWyzDp5454ZeGgJ5skC16JXfSL9CGo/kLZ9EWl21YX
HAHESTKsjY5n2UkP6EXFnFII7GseijviOats66+S1EArLmyQM/gxib4WjGNWzDBv
M4JyKsUYbFFut7xc1hlop/Xs1UC/2Wo3PrUv51gzC9+0h175hDufcKoJe7yCzMAv
g4Ftb9mJ4B2PkCnMPRqxdVLxVWql0e+Qgp/LckQDEs5JD8PrDID2iRbDkSOdscRS
qBgxx7OYNpsOFPWx6Fx4QykA6OcQ9YeAs82LlN1Db7gvNidsowh1GMvvN2HNUBqT
912csBOCBFkh403pR8vTU4vZQNSpsvn3xeg/v/oWg6EIC8nruDBqFsTqir3zWpJ3
Z2XmNfruImEYxXtlQAnairSoctzcyw43N0H3ag0fgxFX840KxpQOnWiD6oMhqCpI
50PLYK0KMbjqVhSbpQqegtWzGPQ7cuwQxXRhReT7QbUZz+GJ+BcL4Et7piBJG9VY
+QWiGqKUidOG6z5b0odbUgkDjuJgAFNyEzETQyDzcAF6/Q7zIRtWetHnvroYR1by
/bemK5p9iLgrE44T2sWSj97zS+T6VgsaTnPp6w9bLvqqyqr5LtvIG0ZhnPAsvASp
gSu/LSoPlkpADZ0wtDwNSEudrrsDi5tCsljUAqFlS7STT6xwX9ah8pb0TmFAJtWd
G80KmdEF4+i3rDCdfjcE1hDRo7CI9fGC2X3646rZ6eRC4jrh55scspmg9QPIy1Nn
njDO5iuTRCSiEUj6KZnpUIuoSOlTt/uEOPuhDHenfsrpkgfu0hDij0P9DMquWWS1
e8JE12lQxzIh8TnDZJfONDN1/IlAeb9HmF+nqFx3sk9rkfXWJIsRmj0UvUB48Wvr
IZwHFXRsLQX2Nm6tKYPthHlZ6OabQGkenjQISSyJgMfH7Xqv88nrBsRmGso18CP+
sJ4d2csPRZ9Sojg+Npbo0d1Xgi5EMM6E21JhjTJSwGDlwRb5JV82n2DrwxrrZiPl
KJLST7VsA1X9vgZ3aGXsZjLiR+ZhoBdJedV/hAW1Jmo8cYDlLV+Fjf3zLkKAQkSR
28v6EihEgS284/rM66Egh79VWZLrm6IVTHqy07cR4MZ2sfYOVGgd6ejCq3YXf1wd
8KBtAdFIHw+yPLpfdA5/1N5zdm+C7VWv0kzvVaUOVepIPHvdVpPPWueiBL0VnrFr
U1MdcbE0e73kgAoSfCJTsMNfbhyhEVgiF2n2gRUhJ/UciHhUIYVLsetORAsGpjYE
7015x3iU/Qoa4i3EvJ7lekODzBClLzLJI2nuim6Cc6PN/91dVblBwLWLsVYVaekt
XHiKQGIyiSYnZtKXkbxlXh20pTqBsOhQhhkLli0PEgcApA0/zqgRGCOtEokkoLp+
aM86/Eq/3mfviGZifKjJO+Jk5Zd5D+SZsudnePXWYGGsEo6yJ9ShUo3kswa2saA1
eK6phA0/2QP/dCS0hlY9RktKUxJELzhy6eme2LioiWSEw22+JDRRI58FD/U6gfsd
FWX2sYI+AARTRGFYgsmXEy6YVn5y4ViKPtk7jp7lW0NSXMRzVjskdbPL/I7SIPu3
A3pbRnJDWix/ShUNRogqEXa46dnqUyf3DXjA+ShLO4sj4wKK2+GSzOXbqzJk2YSR
UcTv0EvvmH+8Q5CdpsnFKHk87EIVPd+uqx6pSUQRw2gks9fyboTzsy6Lz6eUllJM
Bl8GI4vyzQe+CjNC6YCGfsHvpeS3bgOgFRmkHkNvtgni5QK6Wccp7jaJwIhwg7yM
H3QJ3rk/lze9ftqhZEQhP22V3p3C37TWIpxcDOoGV9cevDIr8cTO63l0kwD6FIyi
pOdOrHMJMCrzRDDk0Jmrw1Dz5vMiMt++36kwTtTEMmyP1SqbPZo3vtYMJ65aCNV8
sH/sKr6THxh9CC50k2vCm5WSC5WMuk9dJ60vqDWQZ6FaDil2LfYUEiDYiBNeMgq0
xGluCOO4sc2SBxCwzVfQfWmhvZHB0+DV+f0nrH8pQgTs3AgwWjLDzQK+laILrRom
HiExUOnQk1CqXPvPQnoMDzV6eLAJRQhbDH/Nead+te4exbPqE8KrXm/10dqYHGHK
gWY0ATzN3Cg0Jcs6lleE03Uus6Z7WxJiRc1LnhoYa+x1G5Lm6RmZZuh1N1K2LUjb
AAi53v47drpvWduGWAYE78lmAdshon5MGRoOIGLGJSuNze8vlbWq+0zWd04gWSeU
J4bKQIy9nSf3vXRZt0O4gjIsu2yIBPabu3NuKE8zRtDqSmbi0rK9PXk8rom3R5H5
br8a/RrQQ6lZEtPMfQ4wHdqZMDr8d/rbZs/S8pcuTztiQhs5Kf1BLB6Q7w+6SsJB
QR3ycKmSbEOuFR4TE+gScQlbIWo9sVvUzlk+/NPDpXD+vCvovogMFjtNO/KKcUeR
6tqvgeLPzDfTUHBokD3ZX3mOGViHri/vQP3CB10ouIyho1CIKtseX/ABBlJceSCI
T8HM0+H6IL53OdxQsvNrpKp6xCj7fSneH8pMdKpjQ1ubKyPOJZSfQg9N+mRlV2fx
r3nktYNCuYOIF2zBqofE4NFD4mngoyiLbjA4D3gY+5XzLVs5O8aNoY5pH0kzQyTN
VheAN56K2VbMJR3J55VGyh658m8zOb2zmPXztypBt+0z2TjcNctQL9nGJw+0A8iQ
ejf5DPlHWLKb2edFjbEjY3oG3lLqle8RoyxKL9okY9E00XkwV84L09MPIlNdTP3u
qAgGJ0C1eqvYenmKrov6cnpPfXdRVTQKu+JNd9t6EsOcaz5dJDTt7i0EU05aj61A
aS7T1P3e1Nwg2YrSqqGOjH1YN7KHabRj4YYh3ragS2SRbFBmcoKjr6Gcmhd7w0JA
XrHGUsBQICUN8kzpBJ25r8d3pDA5TyKWHvSlDYIYvF2kz5TxGuUxVuYZ9ucdCM4P
4oJp7hq9mfF7l80RgA0MlAhHFteCmtaSHs4S0rINj7OvDLZUipXb4DbXeMw27g4w
y6kJM32MIqaz6gNymEphb8qjwnYZvLT0jHSqfQIwoe63s6fwJ28QDxDMOFLlMCNf
npdj/A8FAamW9cXrnWBJn/TRJ+dXceGcefTXx/8kPnNIl6TBmLKJh9ZkKzx6IwAb
IXxgZFjD/i7A/0QaAg9h3w3WjmlSl168TvXi/BtHCLmh/I1iM4nLxS7EzZcSN3Pl
uQm6gmxiuNU3uiQZM6GDSnNrNDCIhJvzusCKJTg0cMN6cZJLXmPIs/A0tWApbB36
aKhQr7bFR7QolBZa4NtYiVwycXRLXRFzkF+XD3bYAG3AaAvokCZtP3GIEbuC/4w2
7fWVHCKGGhVogHikV2hGjcxCD8fpp56p20BjoDo44GTaW+TVbqytp4k/OIrvueB7
PS/H5qC2zOgQiuoLH8ADjWEHyBjLI8GUxrf28kyZ7qM0F2xx/5HW+bVrBoMU7CFu
roow+rV5r85pvDR6DrIGSMySZx6dD8uMQBiMrCBhYqmNGCZsmz2oQ2FGT0oAj3Qj
rG6+ewR8YhvhWWiQsq1G30RRvHN4wEWeDv+i4NZEOS3DqclUIYuNoL+if0HrLtHf
GIei6gelcax3z8eWLGnsbfcbbKRMQGilnggNa1K1a2v3j7rL/iiSAcEUQ7wWThC5
Zl7bNmSOMS0euy7CmmrM/fMFoLtspgxuzirXRK4sR0yNXhcedCgcXQUzNSd3I1Sz
EIoGOE8KY56sC8NAunmqhrLxHAQEJSx19QxF8Lf9PbHVsOrfs4x1zNkYasSP34o2
Ar22W9hmrw2JiW1nRH5DY22Uhab2aq130G4+SCkdvthUALJi7wuywF0OFh8d9Kkz
jkhYULnfON9bbLm/dWQ6Hk79isRlFhOsovg50oF8hDAdyddJYGFNztwNfJB8zr46
X44IIryzyN9TZ/0FoyET/pGez/G8Tp4sPMA+Hov+7gkXqsFQu2JgNHcEwVjMGJ3o
fGnjB50rwPFcLCa/GH8LzyKcHcnT/L4gSgbKZbCwVqvDYCZROzK400TEv2gYKZ7w
KyLdygB7xKeCUC6KSJFLMpyEtZsBwHmBO6Ju9RXvxGeJ3yXBS7vWidee2SQy5LWI
y7C15cALBsgqGU5aW7Pk0WAWx10rsV+s/P0imnc6wZ1/BCMapONcWk57DbDpuhn/
yudA/mdjtIDISS1b5M8bsMYb9az47M+64nIaG0HsoqWJMICsQwNMzMr48yya5oka
zUK5Beh4PFxUHUa0ARnaLkCjZZVZkxqFhTCcZlTcx+htKl4MP9DVOOx+r0DUEYvP
9WTjBH2NQgFFCXnzE4hN4nS4ahGTP9ryHyGqA4Bg5npp0Bhm8OIv/40zuMfRIUfE
hAxkmZWbGCk2T9NOuFVVYtrjarfbY6ZY55DuvYgRbcuPVzauo1e1ZYr4j2Za8BI4
kcCojHG7kVC3R2j7bAaOrNuUTwQeFb+MighDtjXp8HmIwzbJ4mG1oUouZNqdW7cz
9ZXrGgHH+OkZaAYXaW8H65ayYvj0HrY9CquX6uF24o/HSyg24yJCV6z0w2b9giZq
65LMiZG070l8UEEBPRI37tJg2ASiY2nfAFSgvnJcoW8a6hCWo7PJJRbbDCXYcPZN
Z2AVrHI0hdHPsIu38bH+esIhHQwKvpE9bJ90QFsgo6ALBO/xtVoRDuDK3HAHERsa
q0VLjQtBA3AlDJUeAFq9eP6uNGsbDyeO9jm9lGzHMX9i+RVAPvdjlVOIL8onLIBS
WfMiZuZ4vJqONoj73xAFyYQNAkFT5kEJ2Xf/QyTeUdiIxp3ODTXLh1CGlzI9T7zJ
EFaBKRiZVbJXnwe72dFrgiBinzbiUQccPZ49eds+4SqePK6ziP1U0jyDTykEk9ca
dtUTKszV29/sVIDRKJMsPDYtIzQ0pWYLk40Jrcn4SHdjsNiRNASrvugpffKAJW68
e0FIRjkk7iDzl9Xci8p3aTDKHpkQOg85RrUi7HxGAizmyU76U/RsyxIOy0mN/fpK
1w4DMSil696UYTMdmtLiWNquqsz0Y4LNpiPWzHRKs2EjaSdJz4kzDpnksORQuhkH
fm7dlR3JeE/EEjq+3mEAYWfRseVOdx/o7IIG//VIytmZuQxK9A8hFf5EQsw33PuP
KaP34H4m2NqUFsV2NCsAxzutBIszFam/U7WtFxdkTIoFOYuKPVhXMKtPRv5ZGg46
lZSaZXg4wvvFG4phlfW/gRe5vxlhwEXhEtT3HpFLncvodJ+BGk7poUdG1qZFvPDK
2eMb9tYjFi3FjTfFjg9+1oiK7fKA2V1qEHyC+J6JkjxeJOFLgbEoooXjYiNDr6Nm
lSOm/jINF94sqOBJFRRotOuBcEiCAvRFmm0v8dnTZeI5nKewOdYOt6xQY5gHhy/I
8oX8gPZdFWH8wVl7WZhTfO2ibqxwtMTQfQZq0wvEh/xeOJkXtwTUwMHKPGnNhIjV
WfdK8kHEBBnNhHmqq7nyxgIg7XpkQ2pjBJRb5VgB6Xo8L+dqmeXf5k1RWE2Hbee6
AIX5tLixt8CfnKSWU6hb2oLVyQgAP2LpDvEpiNSP4YMT5v0BD/wJF81Rney/hDug
79mzKGjUPBCbbHE9bgHdFK0UKirhzSg7JJ/1lS9v2tC0Q3fpqYMTTOov01/W/dmO
Rp0cw7T6DxDz2UACSbDr2GAhEEMwVn/WpcPNSkd0wFgAtrgowQv7V7+G6qZYRZl1
jPYpUm8OkKA/8EPRj/gu5IPhgoHD6ogkPxnVlrcqSaxLlzy0Ns/8OBOZa4Q3M+hw
oo8rz5RU9qyI67H7KPLkcAzbiLBgO+a4d++e6+bnY2CyEF8QBqd/pNPPXhfjAgKy
hvcYsqaY3X/ogGZfEwgH20DyoIdr8iImM/pDM8SfNFfUlFI8f+8YWIzgw39koeBZ
hTitgPVmrVFQhYTm9vqo7GZCUd4h/TadjYIFnJsXgxqfqWhowxcJvHkURbAZuwno
LZN3yYvmnNQTB+RGF6kmRmM4mWsRaBZhPHIMZil4yqo7vBTJfXPWZfx7bvP40Qj7
aWbSswILR9MXlUJwfRz/LGuTvSRu210avfsgogiDHhsrmlMs+MIKB+49A+W91CTv
QDySYiPXB82gvp98+X1X83K3p4Wu98YJ22YDOK0rwzhbrJTYi+QmYl0+qT53/p39
WicOlaqdbTmqWWhxseSEmnIKltQSfjuiU1oIxdCeb0HudK+g2CCfuIy04CVaICqE
3gwXp3hejGswF7qLBY/iu5uTOYQLKUDAxxN/Uh9ReEHLxPnNfJAJ1S+5WBMBNieM
chym4ghW3IYokse9B/cwxfpV9X6fIRZrCDu/QaytJ4q0XEa7WFuhqU98IySnRr1d
8yN87tanBvS/mF4wU9uYwQ/3QiRiA2qCfdxcbTwsfXn8tyWqQwP97qJkT6cqYc7K
xqDGwO4f4bB1oiaw1V1cjZie83+EWg4cTyJFcb9K/XcKOoo8PIERrfcRSZSFsNIb
1VSpSJSTrbB0hXnPGnlnNzqfOSsxNLjBgs1vtiCYXpp7ts25R7HMeDHfbEYtk/u9
Idr5qcpVugVHAs97ZpzZcAL4hJfMPhHlnUDnyyoI+jAufGtTw6sEX7nYyfrvrx42
i8X1Cqmky/C09jX1/U+Osvu1MKR+KfTy6fs86kVN6/6dL9YI/JBPl9Y7+lYxtNlJ
zJUMjOkkAjZGF6raIbJPdS3thTLQgCGIHmrpuFhCubSd/vzdiPBF8gupwN6/+hO6
GFtBNhuBkQWpOacCYBgDEvSfzfiYB/bCjBjYzhTBC80Mbz4uipYeBxzEXoVxM9/t
sJMiS0hfHfKP9conhsoO/B1Bk8W40UQh/ej1TJscjyzOsEj42HgeszWIVd0Nhcv0
t3rv7u9Mvmc2QACczxEpFjcIIRKvmEujhvqX9KWhAhl7i6CclZ3Iqt6f4JyMfebF
eEjH4SEGtwv/9Enh0EC7sHAPEnaVCR/Vxd7EPP1v3FCPXBjVT4dd79LaO49DIeck
njeULjlrEY+D/0qN4v/Et1/giCWiK3TQPsQymFAG5+7ehWnoksDIRW8h6/h/GPuz
+f4kF2eJl+Je/ys8gCM14LG3BER53v8XcsNtOxYMcDxvVfqljHE5AeZyBJ0kNr2I
Hg+kEvNeN3L5Ihoz+Zgh8449RthS0+DDpRoFK/vnbQNqoBOB2zG1b/sulvZHDicb
Hajjl8A4z/9Hos+UtpT1An4uAdfP+fxCNiXIpzovMEgT3N7V+V370oucPy119z6a
sXMi6VBBurTgSHFNdn5Hnbwr3XLeaaop8ylqIzMORSgID/SccCQLd++JtQeM62rV
4Vw4U90jCmj/YzG149Xf9R0XuHE066bYuDjvQzSGG2siSzg44KvTEWVZnaVpjwBA
cuE6j2IKAGm2+THTS5nNGDBj6oVz1jwVyoRAJXL2v9IZPeOoHxdD4k19uFxEABIT
bP0dt76QmriPEIpcpTXuzWP+foV/R6FZ/0ed+Q6gcnU/USIbMu6iZI0l5n2OxcyB
3fhUAUGUTmCqbxLHky2KPwvov6lVrZ+om2KR/8ZrmxdQc/hUu4TKrxwIzPGDMGzd
8RmNH1hVxcvsl65mkITK/BckyA7g+sMgpaogVlJC2KhPKBmpq/DFpCOWkrxAD34q
q3geauQE6GVfgV63y7nWLJVyv1RlxDwKAcSi8/aumndcB/yTNpKnrmYGlSxaPwxQ
kw4xcreH3JnhnN/8b5o55MYsrxzmcFEYE8oBZ4jQGaD/LdJPV6V/tSmgqhrJYavv
QArGHLgA5tr709A0H1vvG1X70r1dQPX1b0wDHnhKoC86CLtz/RuUhtdqEPKqp25Q
6GeLTCMDRFWBhMpMSrFZHcrDPTTRRI99UCIqzya/fhb+GcKI938h8WUwapOjaXqG
psbalbTPLMNB9QJw0MUt5aq5R1pZ0hkBNeMqjtsXNqbAW+X062ms3JzMrZqjxLfd
CZ3IUS8FimL7f+pvGWWiscoPXpSUY0K09+HjtL3LmSxviIz9p6HRnyNFLZZIlLWh
EzXE9IU86eO3MLebf0vOHAaeGJUU/Jum9iXNOJN5ytIRXTBF0MGc44yF0YO2vKCR
RZlzK/QXze84sb1uF83p6tWgcClhdWgvQCUxGk8iv3TCH16RVdJZW03JDbOHwQS5
DLiqoZKUzfqL2lIwM9mDNLrlA5Z4CAapzJmCWDZuPlDZz6DOHJuCSjuGelYI3lRH
HBqnpANV2fgEk1ItDiqBpGJOH8O/85kPc/g2Nfp1ALOyRdxw5JUzJw267gAGc5RA
wEbDZvIfbrrFw6Z+/BRBewlCqzRZwat+yxXmYIYXZoxa0sCZlDueUpV/Q+xRGOrW
/ZPY/QKnRLDxeA8ohUXDR+uRsNgaN6WUoYeiYCdQ6AYaG/zheoYoAkhGErHmqN29
8fI8jisKnkuLhpPdIdzyRzO5RQfemXtFYyddWNiQfxXf8bvf2nxDGCX8/djMx2Ug
ceFgW1oC+IbOiecR5YKoNuUHtWkw3rPUBWJds+gM5R5Fxnlsn0l1h0oihE23c5h3
GePBWWW6ni58UO4bf2G7calNeC7cdcpuoHK4W4spia57hK6zKTvaHzqx+8VHTVYG
1yp5JDtQ02XIFhzsjgSDqMTh2tTEf3RC5pzX8l03r4XpRdAyhhCOmtK/bcsy4A3i
a1tztm+FZi04GBMk1VmykgVhJrjb85PYzcgiX+vZnAJIHs5WiV8u9bfjPy/PWeUn
rmTR+gWIPssu8YO2PdfkEx9iPjFCHPQdudBceZZNlFt3eAHdtrcILS4ao7N5y/E+
BQ/Ev6vimrt5QO1dd/Kh5EiTAN2iXg4o5Oiv8TO2hOyxj6clWrLHMmwWvyL/1Pk9
Ux9TtPl9qQTmtSE9L3wOfPM2JBL8p88Ne5BLE1fzLeHN2Lg9U9rSxmjJKB/m8e8t
Uvg4BY0GKObwsBOyoEMkQzYfKDdULy9UNY1GCR2GyeZgXCz4pkdNxYMjZNYoez8q
gM0VspkDjjZ8bR/9VyGBhOMDCkJfNukYZoB0myJC8raXKsdw3ZOn4zdtipz09aZG
mEZdd3WWobMkIPSoYpIq742QHBJtV8SyySP1v4LCITgm+rF7G56VFIAs3lIpUIYl
VCXZPxvw/Y+bVSGErKY6JK0z0X2+baa4mUws5p9DM4AceNLpg6/NXUXL1FKNNJWS
SGfOX3nMuKdFy14KzwAX0eXld0E1MoDOvYTx4J27gQnkk35uecs3ffDCu9dDCAx9
KkjaGGq9v+IfY2mfUdGtrmiYJBkU++V4CKnVuBtKV4DIO5ynAVq7tCFy2R3kD1gJ
ZN1EQ+KmfoscGbvzh911s6b9ee3st2XPLuNuXI2uUyPNHD4UTuXXxgoUEawh7RaS
jeHsh0Anm3g+WG6m13+B11RZPZmWyQ/vzFal7BJ9bhSihO0PdQ1lElg6DuKKXdk7
yEhBSkLtPw/08KxDZG7pMD6zhSHoCL4U0MLgUH41Pct1S5A1sGdNeKKVTIGm3Qht
U/4UfwBNVZlaskx5dmIJAvqD1pBAZqEDkmEQddIYChyFQpLhOQ6Yf/1sMSX4xGHn
MbRzEVztij1rSTl5sjCRT6NC/g+xNWbfNBuddlq/BDe+r4PaWhXJR+3Zz98quDuZ
Cqih92Neu6NhfcfNuvllH1Vc3+C+kY6Im5A3MNHwT33G6WzW5uRKBTj9ur8l69Xg
SODZZsTLP1PV2zIyBfRhQQ8Lkat3Ep0cbd/iye/MA2RAfpz1iCbylbhVQDe8hJ3g
NK7jY8m5b7T3OqQnk1dhnoFuZj73IFxmFR2oYdqU0RokWH0BxKQDBBayR9Ul8XDf
YXRxW+vmbKdrpGdNBKAshHpy6UR1oFCS4GJmFqU8l5batPvSkDjje2brOgLZD4rC
Y/pKXalrczCre0jUml/Ay2vSCajDkKaLaOTY17uBTebPEwo5mwQzSycEOAGLFpaW
GTMAXTJ+hCQmmdoFCJ8Ttks47EPdktFRzYCeHpod3LSDlYD/GcpETCNcdIFKmHGW
/gTqBXn/PG7f2c9Cr9qHNoPQVtUilGTIocNeZstyWQEeBkvBMeLUIvPp/JXRgmpF
3Wa+JeSMznDcmQ39uqAMVZFyiT3gAMihvRnMYxjzs7HS1xvSWdbu3HR31UOXa8f0
tbc8CNeBOuDvo8VuyPDZ9gyDiJqFXtf/m/mcQDNoZ2yjRPtOx1u2BRHlC53P7/In
/pPL4OQjC7+8jDydrOVrIJ06WcjUlbefhBSTZoSBMl5siEabvvn5MrBHWtpcd8PN
7vzVUdxveC2Jg/zNe1XnBeRiWlyBsIOgU9yGoNzs29sskXDbIm0mgd9UXI0GL+ku
X/YbWDvVDkvREKyrSh145DybkR1XjnUnFKDSmvgtOwV839fuO4QWna9594V7AkPv
R4nd2iGsmE4tVlNBo7cq98kt0mzt8UHsTvM89VtsfoD7plltEKyP3T9PY+PoSvIW
eiNRNZlHLJcKkSS0QO+vRYNfevNxC8P/snLXmEoDITnBgnGdG5DyLbjz8VZv6eu+
AWSs8u+tkv1Jk5SsUI5T4AnBAEIXfd7YwbLo815i/wCmODiHnUVi6DOKyE3BuBw7
lJ6LRwHrsM/i30Y0c9kqN2mnN24M8TBkGvnUL5QYyrBa4kxxcqT9IXzQyYDBBXNo
AjpkRjKF9lj8AfPYGfFrI/MGk49hDmJ+m8oqbwjsZfn789biHI0wVBFblFFOLXs7
5t7yQ/r0DVX1XEURtlnqoS7cb+PEq8wUq/s2DsecgcTH5vPMMorhbCb2ahkEKb6o
TgLTAWlvJSmclxYyS2BFU6Q+mNXF8uEkys0SrF9q6+htcV9UFDkspFh9ceX24vmU
tSzV7/QrWwoNPK9utoK7M3nhTVEtdej26kigbNZEgK2s2TAAV13dIJwP47Dp6UY7
OdhXBVdpPRjvh9gB6xsB9bwo2E8eGNS4sxs5tFnsxpmdiQ7n/SCrKUlnaxf0khYS
f7OzWuQfA3tV9O7pWxjs97WX5f+Apf6jW7gK4tvaU4V2CDAIMMgJIZXeW13Up5uQ
wNPb0eMbzU0LOOLQv+3UMoPR1QDDr2zLwYSOiZyrPhytMqrBZxQKK66wlO1wYwJN
NK/rWAyErIyEjLQzeW5Y80Vq67HeqTJBOrAXL8e+NDPvDFaRmpt6Bs3JNpDl15ot
n50RqfXU5w1npW1uKlxuRPxMt8CgQUUMPiAlHy3kq3Mjsix1rXPm8sEjNOMizTrE
6Nw2snLTk45NuhMAL9c6C5721thUrI03YdcDIp3OPt26aSs0WWBz1gceqEfxAhIC
/WOGAgYMkeRE3BwuWHbi7ZD/Ky1ZH+0PrbgURKR3ci+OI3L3nYAw8cB2s+ZT5Wxh
0t7ghtBmLFD86E2uwRbeXx5hS3BsFeSOPJ+qxXiCAa7jG/XQMC8ENTKulEvWi5ig
dyXTqgCN+ucJDeKxprCGMyLXOBQl14DWCgwzdnrtkdG1l39x3NQr2SXIwEmLG8kC
C79WyZdu1vNP6LnrWHrgVuyfMGUQ5qLD+MwStH5RUZWiclcrNmrVV1OlsLQ0CKV0
jSbkn1QDo4yXr5aPZBtiQnhJkOuoCdnY8jlrFKVhXncUp/bw3IHr9PiJ+zfbaosZ
8oYD7Ry+kgNjfp3wKzXAcW5BmlSlDPReuJoLN53SFbPn01auq1urCAQIcO4QjS7g
pkczcdBNQ8wcQCAZ9oCS2L5FiCPykc6BSluWPlknDty0KiI9sskUCnDXVddAvky/
5sPpoNCupKL1pJgww0ihYEDTm/EGbZZQvIrEVPj39EVeFPZ7d2TmO2alQSVsK7t3
u/aW/Nn0KNwRT7fZuIaObn1oqrazEg1RekpBkcwelBYWeUv9L8EqjGs0AJcQj1g6
BMzKd1+W0rJUWNjsSufDxqucfhBNv2Ff2JtsK8CnpqbmXJzwX5aNJRx2cIeLGGYb
xOhGCAT+FymYbz+YzOc6SQg7V1aeZkvyYAwl4hCWg0O4a18/OgeoB7jF9OQ7tCvt
90dwq+YIQrk1XXgM0Cfq7UEu8J+ufuJc8UDe9NB1dp88Wgo7mKZ4tETU4h2jFp9U
s0Uqy70MGzbPnGB4GFhfVy2RyC3jaDiq4POtH9rwrjgqxvG+HuwcrYY+RtTpeJhw
P4CugGXKx7BrnJqplZh8ZUspCWne+rQxz7bKHLyEQNN37pr/0PHUZj5hx9ZyFYtT
3Dxp4UiGME+Po6MOLr5bicEKM2RlvvNlNVPWSuELQtQQvl4haqdPeIHV95GmCuXK
h4/IYKSPAE+sTHZWjvRZbbwJ8PWupbVCvZhyyveGUd/T/U2k2NsI0wEhS3ux9lRD
fp4c6yjBCytcc81hS2B0ZqTnPbjLyvhf6OuF2mChpHtEMdc054akAAJvKKOO4H4G
H87ZorMyZHNyddoxxpedA2MeRvuLFci2DCYe9QXd5A4CqimrVNwMkKM65W3H6UCU
7VRKzR+0JSw4Cxpd6LNxWgHQ1csXMfNcKn81ZesqDCejJC+LXvKVWcG7dc3z9nib
y5CwM0ipym5Dxql3A4Nf0mXnVmgTiftF678sW1OjL1Mef7T93Cjz6NFmjahj8eol
0IGSsvCRhHZTsLje9qt4dDGwYTT+0tdBgrXLVQER4OmFo+EybQEqqI2l9AXwbVTU
m7g7rgPaTcmeFcocIOS0Sc4r84Jp5UH//QtvXP2be/E/55CngLpF6N/IlV+zN04C
Z1r/Li+Epw3DAjvWpEAPJ3FdwW8A+vaJoqBY2Du0da2x7uXeOeXw7uSFe+WIgwYK
K8HzAubrrAuv2WoyYxYmQXhmugxEq5tljrfDnrwuKZRhnYVAuKM2ujxgHKYBx8ji
o/e9tK5iBm2nfXCYrPGSoDnx0M+MxOE4qTjw2ZYNiv1JxJisArt7Qd1aGIxM9I9m
ha3AC4O2MCNeomdipnI81tdJGu50Fw01yjHitg+yGzl+vCRet4HlPcoi2FGJ2H0N
ieTabVKjxyom0sfCHoZBp9Qf4xPoDwOOLTie+6whxm6W0F2wx8nELCF6Lbu1GXXr
SRXQs8lrQtQ6fBSc3+J1V4KuKmP+s/zEz/bka+QDIcl7pxHizKCu2Prp0nkXK3hh
N23LdIpJotujWuArHLRZ9ZnTO7T7Ufj7CAKc1K52ZJzRkfSeM7eKsBTUJYCkRdj2
LtRhsMQDIpPk43j1XIsAyZVpq4b4w3RzjE9p5rrtFYEYl4PJQqOvLDO0OQIYYuP2
K381U0EzgG5kYrrb49wWvutEdaprbh6A+Op9dTWz3y2rA2g+QDM8bAQGiH83pyMj
0HFTfotsp+7Dkm2mlklIGxWKeGGUCA3GYY+7Jljbggg/q/ipcfWlxF6X3PWk+S1U
1d5GLFF5WegJ4VgdaHhUIhVaLF3QItqqfTM9NIYCq1UCqXYyc3U0kEagZ3tDBYc3
hTgi/kb3vog6VQdCkiwFC9ho/fqTvUfLlrd0xZ8+88WKBP6ssir5VW6d1RFL82k2
a0V4MKBtmST1GTv3922t00oQOyy4QVsFJnlfmVbTju92exD6KqGesNWKISnnxYor
+W5JTcWqpTgnHzhLVpK4WENxlGTtUcpkSNJQbalNg6cwQQjlDnwTZui980xotRWw
wVatIFJ1UXBaMblsQPyEhdZLUcnNV5rLJfVRaGYMu5Wq/T82et66S853FYrYymJR
a0oH8J6Dy8ttFnWyEcTt8k4cVuvk/b9K3lE0ng2xw89CR65jVKbRDkwn9sfI4WPh
KhvVypMQuWQWYbsDfcmC96uIjnNaO9wUkytpOaEdH5Ie3jNUS6vTXHq/Yxwj7zIx
njYT7wxvRp8crEjC9eLDF5wke40r610tHBhZauXKLGvDKSgkQ0bq6ldnqNh1s3Tf
cLYo9thHezAedfEADiInOlRD1FxFAUUJqVA5A+seqmLgHOxXlrLQfPROU9+Mpi/N
3RzKexx8Pm6pd/Esucj159exhCMyPc8jrPxo43ACXeQIx8s0Q5Pel6WhlW3ImPK4
fxFIcWkXby2aNJJuQy+YndaFUCfMCXHGfESCm4Lcn9SaJqssonlGgAJxg83pV20g
56f4066LtNjh7opEFY1zwONkN6B6AKmn8W9iTeUj51dUefdBd7YAGDHlnjOEn8Xv
Q22sk7RWMLcllvjBgL4n5FdCurVeh7D7chqVJd19drXmgoQDclgZPEnpQDvcGyXC
rElPZe+eXUV+DXfXMNGM5MGTw7mFQU7owAvpgbAOc96dOe32GadKpgRRbBvcQllk
ifk9tuiOISIQ8J0qbudjU2XAdTHI78/CCRiH9eddY5WuxQurqMbkRZYcOXdfnWB+
hQ5tBhK5bwx6iLYaw5ZViyg1HOfKYnQfUhXAge8u3Vrn6fYBktsEWG7YvCyVfYiS
3OxE3/6wWCV/2pbflt0Un5B/7fLVhPrGDkLz7hPzB7H3qCbhYjrJ/FhS49hZbsSj
R8hnqp0zgXnQPHTC9bYnaRzg6s4lC9fJcJjXbLe/MzT3cMmaUL9S1kpXrJqCoLzF
dm/ZbwKvCGu0L4RD/MVBtpYwh2tDAj8XRo66K7j7y6NeifwsOb2JglobCzLAZHBt
PhyVwoyaTxdpdTKIHbJE75j7wuxsSZ35QHMdxawLPISV+pM2M9u6BBdLDGJljPtP
/7Viy9Y0adxw90k6f6+3TZA7ffdkVhYSAEQCkRNR2Eca38C4onv3orq93NMaBtwt
J+AzZK216SisyKhPVOHWPGnovJrN5t6oPDwxed+9XAKdd6C4YNGkDF7QWk3YSlUf
g7Ehw2oX/FWVIJtjwidt5FeJN/BUhLESYc9u/0MWNFpFrxpmNUkjfMf4aWvYxMX/
bQRuowS3aH/9s/dKsYdM9kgnzhvB6C2Py/ciZTlj7CWRhY2NvI4UOOGWtwRvX57W
JLaC4VTI0bsKzutzrjQx2p1EBxDAS25jT0YKyMAHmXq2KXE2tFisFlBTQ+TXNa66
O3PHuknyRUTDHohfVzu5M1iIwJGNRNd2sFPrPxl1mNq/1nI5paYDeUvGukgYfEXb
Ura37GaChYT8PWAOZXVDVhw4MExPyWN8tSre9TTpT+EUYXHcKbF/im1f5CbGTkRJ
yR+0+8DeVBotM2EGIMMWTdBS/MiYJfvDDcTF8B9pAk0POo9pbrIiB9GHBJWeBLj2
vKtKc/yThjwbhP2inCo4nwMtNnbBcuZblf6OXcCduH0YhKIcLEiDnIQJ2l1hNJJT
ZI3S0oHEw0U4ZB8vK+rXFvcf7dmAAupgdlkH48nBq+WRwPkNZXHYhXoJ+t95rw8w
PSC9qhnzofvdfow7ZyFKbnH/cTcAo7LIutzWviaJBg8ro+FSjmgEzgzFygB1m7Nq
AHF2NoiPCSo6V2oe5W+dCJ5mfVUh/Er4MiL1DaQYbdUs5CZmH7tXV0CrZQXWqa1g
SnT3pb7SciKHioqJBSiR+7t1/6IBoRV2TwQR8PRm4J5z+iZH6pay/HdwWBTWNDAG
CacLtiPg3wxbmn8H2UMS8qqF+JZCssMWAc9cWEIBq2qDqS0YYX2QHzozSf8Tmuza
JlJ7teWZZ+RofZOBREYO059LVIQNA/MSSmloglwMF1KheGX+4SmfRV/ENuyFDkzx
X8LBiCQaIZoHJokb0GyyRWG0UEiJMsGOBErtbOu1QS5ViZnrAZAuIc9FiwrGAMBQ
LFwtzeoc0HyyvfwQMP8PlQchkzSg6PTKyLvjye82kzYC6hOMByLwNTGqH5lUFOxY
bumd/iJMlfPBcpX+Q9SYg2if55iTy9TAKS/Zld5KdpMSewXwiyPMKUnNQyNbar7X
WJqcZUOgSSpkPsCA6d5j3NNg1Alp53KM6XUr28DatTIVMYe9IqwVv08ljiswgllj
K0tdSTrWSqUFKHAdAk+NugNpKqKTY0baySMkslHI/vpvHMactjc7XYRmOi9QCdGZ
P0U+ES0EOIQXw17r6RpoTyggBbatvr+pGwRj6RGlgoLUHxNfkJANsP9E47A4IGf4
yn10tfxqXS2zngSOENYV+LQ5QsRBISRZLtUFbDh3GGoRJKgHu9SHskcjuBH6gCxo
xSIqZ11jlqYk8g9afhUk1IxKj6BZ/oFgJXgYpMykFPDj3mxUfyulowXeV3JM9B0k
9XRSA/9lCNH7Vaj4SlxmVyj0Ycazw7KXFsshiDPzF4m0pdOPFBvflFgu3mzoN/dj
lIuAFEpRSsZL2tay7mxuYXK3bX6nMm6SpsoPR9gohlmVgU2RDe96Cz2oLZ6rL+1f
9sUiLWZtYJhJMMuKu/Trig6O54UOGkFx+lk26SGUXr/qwBlgDd6AkF5/TlFntwTQ
S4pdyJaLi0PA31FYG0Lwp+hbBbyTLHd5XsovossKObCbcfTJ7NUPbySZhZBYBmEM
xZdUTw/xjY5tC4LWoFacM0tDroAmiNM6J+7U3K6fiWFQ802dU5n7O4ROQuetmlQu
tp/nKa70PDkH1P9tIojlpIl2yjzM4SHW6W3S2T44Bylswwtb0oRmFvVQDXvG8hA0
TOZIsK13hUYRQphqnSrsn3eVoNdQNmLhbSFLe1sefJFWKosaUAJaIufONGWzDwDN
jEURwJb7SgC4cZA1Xyn7uBR7nm1nNofJ+C9j0RXM5nVhA9bSAQbzEwcXZDc38DUe
ljpievf6k7+Mf32ef8l25qVqai2eQi2DkFpBg6N+0Le/t52KjmI7S+STzzCt8Y7S
AbLSaFJONUitntDGvYM6/FxilckS5+gLnxjhuhJR6oZc3TFK9Msu4IMJ3rsEg6z1
sGJd6vUQOaYOkEDQYvvaGO0AFoKRb3D0ltZ5fSESI3Gk0L+jUF0Kz7F9tg1ZAi/p
u8MoctKbnPpX8FcnRAOXAfT8UvwmfQ66alhIujLr2lxiN9de30quGLsgAmFWQxRW
cWW/xN5ojisorjlOCE9V6mcpho3V/JfQUHDMfTsVNDFSwrh5N9m+/9FvViuWHdlX
5m5zUtcx3sIEKM8U30QkKWj8bwSbbHbd0Z6JarEOdam7rOh+4/R924OmfnOGd4tM
jbEFfHiKPkDHHtnfdQYS3HxCda3b8ryW5kM7o/xCKfRwdc2bNiBsKjDW/gODM0Vt
vtUNWvvUCAB9USW1X+M5oKChTKtplPeF2edtoF0NjCt0Lyq1LDkzGTpIk91fy4NV
Z2OQshbuAoVVEsC38oHIZODzx32s0N3L9evYG7pXNl1UvO9uK4JcPMIdKalhJJTQ
v3HYRQHHLRfmxCXOb4loAQr/dq5+0gLumFW8+8P+gfn3h5pJDy/ipRPTYpkWJBPT
ZJmeYSDAtOwRZjINaojw/BkUTVu/b9FIt+M5IOzEZJT0YdHoupor/YEkanPj5WsF
bgYzgmb84SJQiZIz6ATPS4wJa5alLOfIIXCj6c7DE1R8/+nwpIpgAs1OZ79yBP/Z
6CJHydEy33GvK13lBPZdkTN8MGCU57loJ4roEV5O56kLO0rfhysw89afBPpQAxFn
T0AEtS4bCmocuqO6AQNNJW1l8tNqKB0W9iKsbroCWiNp2TltPc3b5qOH8iR29W03
tLSK1JJ6FF5xnnNv261WV5R9wtknHT7vxr8Gzvb7eJP/yKBPbz0Nktvxjl9DQIbb
epyATlIt7nbvAQGJvTzRgV+VqrTJrmMc2nWqQImjPgaYgapmwQCMJenWU6aUoRA9
TmcdNna9+22tLIpYxaFZuXbb/t4n5f/4w6M8twfIpL5CxXJ+cM4pvHrcRS8hnEDq
t5xHgx6dzsEXBXNhXzgEVLUHrbgKxc4tFMZxJHanefZcl+43BZEbhHcIICMN1kHI
1oQSORv6l/PDZvN4lbdxmJ0P2yslUBp1V2N0dDpNkXRHa76QLZ1HjNmxMlejM+g0
Eqq8t5yNVnbXdtOMhH92nnTi6ZXRhS0wLZ+XAol6mPkKsqpLzWdPafpcYN8e30qK
oml8kkwKQmoU6OT6DgueA5kYrBM0yxbxYYxqZi+BU3vQxE+M4ILqoTmxwSficzn0
xRZg2d88Q1WDlDnzV9YDOAM0J3ZJbV3dU2Lurx24lRkVq/1/Ik/ul5CmQy9Ccxnk
Ts4IFL1XTY2lGnUcQppJoNwAbhRGvVJQZG8FfjCmWMAgP/LK2zDulVljMEJsy2BP
2QWgTHPHiLujZjfiWP6T86nZhi589jfalXbP9zokt2e6uaIl1wOYMmVU3FaqB7Lh
f/oiZJ9FW72CFgs4iw+OPtkWaOIW8x2aYZTBAt2jCLVpblZ9ndezD4Fp+SGL3r92
xtD3vib3NDh689BVLNeqLLuFDrLm6ETvHTxUOE2uoPJez94JQq0l0vmLXClRSJfK
EuLWPJ8MMnzTudv1XPGnMy2jMap0tMlAxPDguK2Xagg2izkiik1Ehr4VOSGFxDYb
R72MkyLVVkbB+prMT9CBWOmq+y6RNPcYw28MSwwz6OaisQ5CWraO0AVH7EhDrnu+
6l5El+0cGCrFYMA7tvOW4bnAQUVv+oe0iRCK7g5wVoBAGyN7iVYb1dOSpq7hQ18I
r4fZdbevdthFAlEQV4G8xA4ioNwRRJhMaCJ8TDKo9CSDqImQ/VjD+vwgEaJDKGF6
Pm8G4TlMs+DUZivAd2of23MdsyWgu1mwjGyTlvNr0HrVi7z+n2EYBcBjYhQO3NDH
2gKj6CvJU11CT69SE/bgoBv8a/Js08fzW0sTuOaLwwhdgvzZcPlzLPTYPH034v/p
yng5hMbTPB27X7ngDFR5rw0rgRxVuaGRH7LdxziyV3zJchqvYGQmEfxoUHiil5Py
/MlaGda2zwKfL04RdGTFcjvckKPKDr+ut0x2PjO+CrzNn+aNp2kMn2nXg023vB3w
ZG9vlkXmW3X8Ai3+s3CBUiY4quuz3mRwZf1kpa/wzTqB4TcfAd1ZpTgiQRw/31xP
W0Pq5afjB5y6E8Tt4n7iOwkJNKfgfbkyoDwLAPi7wFZsYslaACrQX+Wh6P4SguhX
/NnQMPwPp8lFWfNglDMVg4afgpxwcy7V3jekBbG44OJUYNAYtihz4UedJZa9Laei
KAqifvsrqGMuWQA1Po9NEwO1pOo7T/rCJ+urPCW+HV4lUNAj86pTYVuQjPpHHmKW
O3jhKihsMHwIOgTFjB5BROCVTuG8uG/MAPDOz3C/odSA4soDS+ActelUpjTnhN3L
+Vnto32wP1F6D8jQfw61Zm7ZWPfHkUyLeMsIp6T5EAfukKspG+OqQ3Ejvw75YvMC
LRnXR7VZ9AJ5C5Q5mUGAw+ttHVNPDQXsPBBwDUh1X3Yf5fudrqIMG7MwJ0Rc4KZh
CFK6S9rV68jIj/TxJLTVlvi8ZwD+EDAuphM36mHz2bRxThLvE6kS9vB1hP9KcLc8
2ygI59JXRZX6+HY+8FJnMUjY0bD50ZrOD0jTMhbCoAaYH3L9MJ25u5GJWM5fM3Ux
UAT10+AuUq6ID60H3s1m8hSifU13ByZfZdskAjitS5su8kgL2xGq9uHVt6ns5p5b
ZA0gnY9wVeupF0vX/L3C1E93FtZMNHo2aYCu5Y7J2vIQH7N/YnqVppcv7jRZvPfH
3/9h0YzBRd6T+SVoQNnQnWYTKkD207oAQf/VwoZHKRwRlOsAC8ZPTROwYT6Uo3aq
gxvC3Kh/hidhzRrTKeJTtA6WIa58tVt0sTvkEhziaVPI0MIdiejrfLFNJeg16QPW
mG3gUqALD9JtoF+6fe4zuhImzJO0F/d+aLHnL1D6NIdbVNhfz36aGtiu0AsUHRGp
M5muZPmb8IxZiDzgoRbkGmVCcs67kEr8MiNrGyv7VOPcrcA4siJuYHjMIb5oTciG
j1uQ/bbU6IKr46lQc54wfLGUZ38KDZESruTAFKNuzBQS8ZnTOMMffIV67kMbl7TV
Vfy4oWSCiJTIPsBUXewtD33tRx5NQBc28DjWV+h+DK9Um+ZrJa3ZbVKJNtL/LN0k
OmToPlx48oVlqpV/qUzEWlYY2sk/xWF3VRXEObDaUsqWbSMVIfW24FCAzT1Omp7X
wCrciQzyCbSWqIeVTiXijp1NrYuvHd+jYcprRE3oDbo9m1LH7aapU5yN2jjim9m6
X+vkqGvIEZ9D7TQlmtGwL/0Xy8UWtzZTEFoLQxW9UCg44BOPgw4ILHGnlTgBDIx7
5U0uGhvu2p5FjdATeMOPYych8B/5awQT9CR1X6sLVR6LZWRUhOlEeja2SXyckFqQ
wJuD42HP3lOsERkOKVTT0PxhBOVa+6cHID6D9Bk6Pm15HWutg/JDdYBOiiy9+QHR
dO55TTUSzwvJuEURs1pFKwwDAS76N9ejqicHa8vWBt03KabqXqFYuj5bIG/be7w+
uh+nii1rQKKAACpGSTrOGzmTEc80NFOmV5K9cViw32mxBwZRA1g17bC6VOXQkPjn
/vLUs63XIUjz+8XZskQIDG94T1fJiWKQTtyRGdTTClyBQDs512yuVhtN1V7Y1NYi
60QgKjgltneZphVQB0H/iW2K6L9qKYWbvIYK8Uuss4KCopQEsIUk2eXonQR7ZUjb
pwy5DBbbMx8xzQE4RyHbOR2jnCszAjfzUuY1Y1SOtOFPkRcKAMdgYzh6WMtX4yDg
NtfNY1UyMo1MrgJyBj1HpkSLMfNr3vqEVpGcrSi8/3pW19CAC5UrnZYuKZ2END2P
IRct8VRv0KbMBDp0ZbB3iIKAyH/tYh2nlWWT5AVxmQqEFkwPYNlLLAibVbRGee+1
9bq3NOjBoyNgJ1rmDAOfe+xlHgp97lZnM4smJAVNnMyGvhenuxGEcXaiQ+Ms4O5A
JPSLPr4G0bZmLtIKaAAtNhaBarg2ie5cwgAQuDntVedwoV6ZtXHpF0Xws0Qcf5W/
S/SDMSKihaT61RtpnI4/pvzPUgbTV7unIRKnotbcCqNWr0+AHkD4u9/wJO6rvlJA
F8tYto7N8YSXCx+TF5m5BD2FSFoBg3qZM3XpP7MCWiY5AN4MQi1mNLPRAQbLQ3qM
e951Zbt9yRF2l/YDv/lrlzR2TPn/axMLgczRMVSx0FgaEhrjAF2gooMEolfk6ASp
nA37oPlkr9Ehb6+xMIMxbAk0MziwgXbS/+msdC4VMzAd8N1Vy1ftdRn6+rwW311p
V0aekIOdzpBwtNyAe6HzcweKfLyM5mTzIjhdh0SJghOQSvWHTuCZyL4RzDuv75s6
M83TzN/Dwh5//EKaxDXvADD2TmMCCJSjTqaAQEU2GRiLIPKpdD98iid4N6v4iigb
HY0DdYfcSD22LwkiiarcvP0VDpXL4eFgc9qApjZfwm7CjX3nxz+9woZihjmPHpvP
FyxFSFm9o43MSE5n+BpZQmxWgImpsCiIxZ0Ba0xEYQcrca+HNU5kx6J9ZLTiP5Ld
RfN8Bv84BOyeXcc57l2CG4Qst/M7G0Xz9+rhpNfeU0VLXJhYfZRrKZfrG7wEP1A5
lN27aIb9M1DlBiWgHpoRprKDtLPjskKTFeEUsqMe3pfYh3El5bJEgxUgWRnGUuSd
Ox42pYhBCq/WqJ08kFfTRvF69RNZpqHaGTVC5TsmTCDKLak38ebCNI//tvgzXNvW
VrcWmFXIxf0rzy3WJbD7htSSN48Jf8EftAZaPuUeEcTcuGUdBVrA96em7tHzqTIR
NYtk4jtG4y2tJxRRHjTqc6DUX7eamvAf0PjhF1F2L7w6Ss7UiBYZLj4KVeOmnF1/
/zuoMSr5GBuGNJ4XFDEav78iNV1cvTexb9tw4j9JnxeUpx4GvbCp69Koj2YL0apW
yDarTDoMBpZ+9cCmB0phGupLDcmwbShFRRnswqz+sXfMXJe3q1UEiD9boT1l10CW
3hwT/j//BxLBFbJ5jbUWH1F0oxtjxjfGdflIvn3ZTtGJtMh/rW7a2AawFF0KY+wd
yAIFIFtIAO+a6WaNPEHgytNC7/vVmbIlGi073eyBRmQ0kOeJW59m6QzXj1vni4Eo
WA0U6RDqp88DeMrbfKylYrXsRfH2JLODeBnyIaWx1O6x2yYJmptuJbNNjwL1RBD7
vuM32IhfmiDQP+DSXXDGaBEbrr9pPV6tTr/KnF2xH/p6Mxi8hgaIuLcrmG/5JNWs
UK+l355hrKug0ClLUYvf+pW2eTqxj/r7UfhW0ph/ArGNwliGbLiUaDHGMmt+Y28u
TgJQJpHPNkFP9Ng4/abxgYTYSntc2jSG3X4Nuhn0570e6VkuOa0vF8H/a3NgtVvw
zF0Rj98QPciA80OcsAWhDiXvRpoXpxzWqiYnKwJUIsm5cCYGqYqIgWlKV9HSQnPh
4B9E4Bdw1q1QA/85v5PuVRJTly2JGP2Xpa3wjf88oTvFd4Wud3VM+p+uQ2oPF29q
sV7K3RgUpLs1r9ZJ7cohgg6XmRg9YTK64MTiGIv4akrHtC7RRBDBtENk4lXfLd/1
nw0vSU0aoXaY82uLbcpxAWyDn8Rjsg+7a639ZqHi22TsXXeTqB4iTu9IsGSRVVSq
94sRZ3HTn4oO1WFU/cwAtq0m3Dc3ROFPec3R5bbzSJRiylZhoEzoA1LFwvpnGneo
C1qk42+BJ+xS5/XBZXEfYQZuZ68IofUjEmuaN1n5wZZ0ed7Rkz1ltDWWR+dp3OG2
ElkRugZ3728peFfMsbHJHPSuwZOsq/qYWx11qSWqR9H8T6JynI62q4GSAs1E05nl
3ec6/dJxhAIhrpKNNiCSxXCOLzpFQIhNlBFD1b6dfvN4uZjF0BwtXxV4X+0R+K4Z
KwOO7Rx1EgRk8FeNRi7AbOB7OROvWgjLlUMyFgFvEqG3MmOM04u5uEwZi95aAqfQ
gqAyMTlnxieNAZsjcndadxMPJoNqmmYabG4kBNgTBtS08RzRLp6OLjoNesCGMdcS
Uo/Sxf8/6ZPZJCaVPqrJ0qxygI9xeU3KdjiC8l4ZrLgz0K+QmyHq2MhHIkDtgRnh
nNt7tl4HFgx1OQqQXc7UhLCrlu8kb1yMFGrSUI9gDUqeaCL2wJbGKcwcY4WiyK8c
ihE4YKfySxGni7rCr79ryHONYDg8ZhDT2RR+z9Ka3UiboxgWT933usmht3WUJx7h
hLAir1IO4kidy0131BBxWtt1C28TLDVrm80bYmNKtA38tORCl2hFOYzHYjkpxo/j
AYZTidHQ+1hnmW2j8/dJR85VqNSvyRjN3De1ZZmLiwnGHg5XEVHr2VyRkRNSIzvf
bBu7iRorNYxA7p4UZr9F9DrUmwfmKqr/1s1VS1Mik+aiK8X8AZf2FCRqEAdgUaUR
bBzK5xnay1xI9utOLNYPU5/nwGZxLvp/M34kqX553K8B888uk8ii0r56XFEIGmV8
9oPOUICXp1sjjC3Ukt28qKSrZCuMza5SD/qZgIwsNeo2QgnKpwBLkpLA4gW/mlcg
/tz7fS4mBMyqyP3W/TPW8uXrjFYZjtGH+wJhYk7ihIQ5fDdyYZbr2gkGhRx2svk7
vokeilIbLrJZ52NYYWTRIYc5Cy50Z9JIzzxc/3cWu4jEIL0+Q3Yoip4BHy2imdKz
CSMQggvtIz4Lel34U/FvQA4wrnCoDixDaxp20ermRxSuSUoRg8YnFaQEvVsN95RI
StzvOkw3riUP7u77ANQ0n2yH66zK73tB+RdjjEA1IRB53/MqsbWaG8E25R6uOrs+
WdyhJkyZYhZBdGmQddrajJoDQMwj08gIg7BocigCzqIzd9QTyiFkVVyEGHqT7RKZ
IcNYwsXkIGxaZmtx6e8qKLntmMVVwEAH0aZnqf12w0V4eIgJU7fqbYtUNo0EaVHr
13bbTwcJ3OTbLrPMvWaUodhOi5FlzuR8R3sz92rai66HSgGjMYj5yglvBpuHHxn8
LnW1FLKp2mBgKL1qBpfCYS6pYD4KCDaw75T2XPXDcAEn2Fs4EcyfuqbYESF6CDj1
x8O4UVV2jq3TtFXL2Q4K/CdB3JE2L+01bcjHxN1MQFnl0XD2+M5ddk2FbaPxE/H7
hFrGh6LCMbwbAIgFtg2RsMDwAeZ0F5jLbtslySKSO8p7Ka9fafSz8uJVi7gZcaHa
F2CVDaAFpsK6pJztjXxX6JzD3SK52dLIa2BNTUGMZZtWDPojMZyD0oFJMIkPUH2Z
JcecS1ETYPdwRZwKZnKnGgCvO+49PStkXk+HJoFqUzRp1ExzlBZIX9fT2PE0HVeU
/yk3LJ4InnwAjesX5yZTWwiokgzk/XGWb9r60b8UyYrJSm2EhFS8YRuRVOUMoxwb
7YpsO70Y3VOTbamD2OSNl90xgriG3fJ5xQcLdN1GsGhOI4ai3jUVmCIZVbZOrcAn
stafGd1KcSeVQFeK0Xfr4Y4tjGz2mD7DIqL6+NyNyuw8Pwwudi7WUhtqrjYtPC3f
CHQPU7/hnSWFGzwvaxsYFMOTlQ0vzqRuJTfLbYP+kVNEn82WMhnlfKfNGQNJzwT+
M+qntN/Pu7bX2oouXQg/pnSZXTsPlb1ODIhD+uFmksEFEraJTaz3JYZXFlTYoauB
izL9LDZplleSmhKU2rJK965HpxoUpZnbDNiuQrPb7ZOSX3/EStqfUSWKI0Ca5obo
U/w/SyD68O7KyEkM/j32gzqkeUThb2HSpxhbxsI1aDeL5Vj2itI3DhAoJ/bC4sHr
vliNRUKeiYNDm9rf9EVVKO5PoBp0J9wJ2om/T1txYWqYc+ELKQvuFz93yQQv7F5x
Uz0rcqnzPPnIEqUsqq9uZK6sXOhfh2kQF43YiJJ0ee4WIBcCQ2PNNXyhz+oYNbtd
5lZUshIkWQdDbucm9NDt5gHKT5JoYF10FITgv+QnfHwsv3w7/snsLpuQJWQYftc6
ziDXOHGa1otRO0F5ONVIRnxJHhwsQuyvEsyIfJodyVcNPI3ERbuQ/STd+FzxAxcH
fLbeDHWHKbdfCBWiXRlI38UOjAtmhNjqh6sm0ZClIIfN/G1eUr3mcZU7FDguVZfH
IraWPvcL9SKHvqbjoi99C5tGG75iB4kruCmWLXcV6ghzbl6ZbzSAz2saE6T2uumk
yYpjNVZNOfzRMG0eYBLJXEhojocl204GbVjFiV5D2O64NIIJObgoRG+/OJyNRpl5
hXkRAS308G1zOg+jz9jZOkbh76xlBwNhIiAZAUYbwUtBZ/eYdOyTZohirccuOEwX
Aac6MotjiZ79CPjtFEgNcCdq0limWbxtZcZqi8r/RPa12K47up3Z4aT3ZXEmz18a
oiabc2bhY13Z3MGa6UvcwfvQ0dX9f68dEeZ23HvSGqUqajB/z0NfEG6vm1n9fenK
drhIfRSIfXxovKaC9GFtZOxi51Qo49C/3+ppyVP0kILOCqvXvaZDtd5hh19oUue+
bRxHlm3iZ6gv9wptugnCNSaCrcPj9Tfu+dKWSlDqj8W9hjltYOmBebsryAlcDtWi
TDraVCYPC9AmbSAwC3f7OyQI3hFIxNCreNkcEBZ7VnypYWG9pyZczFUo0UldEEgw
dEkUODL9xb46te3SG8S51efgKje4M9kvi1FkxeAULYW7u+xi+b225WOLq5uaZpjq
1KjTar9JQU3IUhIpMsW7OO/46gR7ZoXbIfHOC3S0IAW0M4rEwvO3qja0MBjfrmxa
kX8+IY8WoDTnxB7Gj7LGggfNqf8Bx8avQg/6vCTwoXniGtBj+JBIXmpTtYei+Kmu
m+P31cvvrPq6uoWuXz0zwjRmKH8szZ3LdIWtsnT7ETJWJWAS3Q0Lk2Re/Ylu8gPu
/ALP5w/HNv3VDJktTlrpMqGC8wabS6jxlksV0tiU/bEsPr6F7SINJFHCAghxNeGk
KQonCroBGmt3jCHEtZH0tNpjHlZbnPWz44CM/D6mQC5riUVuwsWDl8gEK1/u7z3Y
+L6+bfzafyw6EnT1V/BjeuG4vGrNFVfNahHH3c5MGgCBUwfAEW9YXcm3dUViWuWy
prrh1j305LbCR7ZDFx/4xLOW0ltPZcHlaLmh5V06xYfy2Pd5BLqjasiIBdu8S5m7
mnOur7o3vcV4Pp3Qz6T8Dkl6iIx/5aL6aSVX2xYP8WoAa+s5cg9R6XKl2Nz3L+W8
BkBqn3WlxLAMF4vapOaFo/DRhhhEAMiM1VyQItA8OjqI7tpI98y/6a1UIAZ4P3RN
e9RLfzCOezKhrUO8IV40DwjAIv7MUkmSjxSknBWq2ojrwstyF6s38Dy30zSBYt8I
wgVk3oIqKQBVPuOWzk4UfV5y/WBrcLeKkqQHDAoaII784uUbLxLmunRBh68Mj1XL
gps4XX9nqLPsHqjqDyynHgAHWC41sQ1yWXd8yiAUIj0sMMTdyZYV3sr/UknNXMqU
SEAoql06fk5vFtBs7fLHwwaMLMAbo5PO42Ib1ZhvggYDVgULk612kjwsJ/LSSk86
b1rPvVcbUcE+OU+xddhHA3RuGlOFYfFsiwfNiqsDc9BvCT9ex4NR+1hXU2PK7eU7
AMlptiz4MAsuLNbmQ2EimVU52Wgyibe3spaj5DDSh5eCDVBuIVjA3mTVqkRXaIgA
2Ok1Rn6j1ROrCMMq3aI6xTKmcemGeO1NmvGCCHhBtVbXC0mVchIo3NonlKC6ovIh
mNPUVrf89VQj/MhMEhHMugAMIWTzoePjt/jcTeqEAFfzj0J3/2X8H+G9bJz9XIqR
38wTQJF33XVjgExtCsYHLn//0mfSF/J0Dz/MJFqqgXXOaRXCnidjq8ZBMRUFSfzI
Bu0RHA4IUKiLmiyXLF/RlVBzh4yc9yALEPR96uoPYfTQB2+GkvFTyVk1KvsuqJVX
JGNqZ8Vxc9pAOp40J40kvVw3vfwRXgulZs+GjK8+ZXRNODIq0mzuViNH/nwCJ8Do
RfPRYoxwLRLtNLSLVSsFBR0PzZq8cihZsMYdvPIY/T5sgHG72cG+cVuuLVJoutc9
2f7Qe40A1gvv+Nrj5x6vmZzkZaHPE2jppHhgBexvq+nkKvVrug9iLPEmcAS4RlSn
AohQO8dj4BJe8ROYxhLmAm5U4oGrb03gX1lxn5UU2/iWLJS0kOnfLqR7ochoO2i/
YWIKnGS3Wls9w2zyy5ujGCSTtCDxI2kjhmqFGM7xziGaORrdAcXumC51i4ownAcT
x0BRm9NYoAz1XmfrKTIQnFg5XXgoeqSBprx8PpLI+l+rqVNPbsyK+TpU78jQXJPJ
EuMMccTyZjtymmGPrGZQ+N9YsrX4p9VYJuzOiWy8nRVLdaQ0PahjHmELeDFvbBEr
6VWUcQyDp2oe5lemjGUmcPN8smoD76kjzLWanoHjdqZISucZzt9lnqSTFfmpBu+O
3vbHEcHtGnhqOrr6FOjQroWRXi+RY2oWUlSdWT+w8jZP2WVWMQ27ij7NduEg4eJ1
b8tWncMGmK2baNZ1ZGNTWY8Bm+0Di6uKcChLWZ4D4fK+8piz9penrlVz+e12+iF4
2Bjh5h79kYAOugbnpWCuSUS/1d88SS5I/SCI2fAoO1QMB9jncRn+XEE68OYPQllP
v6Jt/0mg4of/XmNnuz3sSXFfYXH4f4L4priX8L0KANTscGiCY1kv7N9b8zdvuABO
ogJ5P6QEEjHfOm095QpllbSsBCpud3yJWChX3cnucYQgYqLcjz5CM7SB9ifnkfGI
In14x6FpzHSK8gy21Z/q5ykwV9sOFR0m1fxZOenAFSugjVyKbHGhdUh54Mlk0ign
gJN5q06R0eA2ul3U5cM0kXgsrVjph6cvjZrPH07IUQ5wBuU/EA2CQU8oSKB6taSo
irRLaElb5HXDZ1R6oGHU+hrF22zxexwgFAYscxgySXvu0zIxeQt2tAVEWeT5ERtb
ONRdUbQplNF6GiiPcK25kEk9gnrTbQ6+XbHVT0KsZPj1ucORoKffZeelCSerRIq2
TSITn2ZKzKKpt0s8pt273XvHCGiaM4wC64HpeDHUb9sn+OCcgL3MrI9pXOy31EVW
q9HNH9FLs9NFd5bfi+QSSl57hGN1MzYbMojzXUTIox7P34B7rqZWerUe7C7CKtKV
PozBaSZW8qfmK11MOScpIRivdJqua5cd+3x4B0iacINa8oHZS0Kaj+ZjRJITPlbA
wFIISikNcetmAaOdw1jW8NltsvnXu1CFO6XmVnInw+nvYC+ivaT3NVCCouW9LBgC
Cmgas2FMdiE3Zhbc0d8WMi+vyfhxVqY80MZpLfYTkIEPMCjsL3jYJsCYdl87xaJj
BP9IFVXKZvIH6uxjSscAqR8RhSz7ssOHQbwajwAPBUgqJJs6Fu3n2kI3YZVN3aCC
zO852AekqUtFFt0N1+qiLBe2O9RGSdo3UK0cdQXojSrsjDLtEk2Vuchyw8x2IjGM
YxjQRS5ekVL6H+DFROslgB+Fu3JN+J70rA2POA178kEYl2p3Yi2X5BbcPRM2qXYQ
nl4S0QXLsPZ6kGurWpcNmadAPu747naNDidH92NjFq0mbUkI0tm8UyXGszSR4Fqm
16TNSaxzNTEjLB2BHPDAXO6D3fTLE2Xkexn+FeqVEC2KYwjV3WKFkoQQf76Sp2en
zeSa77K5G8B/Sqbcc7av/Ta0tCiolChPFv0e1GeGHWNab/NgCin4x52VNh1sMeZZ
0yjaLPIm8RgLQpbX7LVvY43RrRbSHSFWDrr+IUA0IjvuSIUdXlVauPYRGII7vU4R
9MTxcKBwgWIzd7HhXHvoiWY7QUgkwoad3lRh53+R9gh9zvJO5+ymXzS/Oty2tUnS
xD0x5MaEMugHeveztzPFG9+CswxnWfFcNng7UCBiNKYnALkT6TMAW9bUTo3Su/Ar
Ym7uPly5e9vjfo8RwMzfNDcUNHVrDz0ktNtZHFyhP5F8kYNA8Yi6G4aJjMsX8bU6
jq6swTTTKz8TwcYu29t1oA6xSpvmNaVoYHkjj0+jl+FF6m78f9RNuxVR4POZvToB
I6adtl8ug5c+jrfaXMt0zPWexTRWpKvEUkbQBUi9CZQdf1AvDWQ5oGNI8ar0inw7
b9J06dP9z2kQEV+0vdOfm6RBGJkQWNU4EM89RmGkXK+sK1BL34civxKYtprUYOgC
ryjYX8vihckaBbfCuawup3SpUIMD1334LWqDC0wiNckpHCZoSZHFj25L5q0wqC/c
5WU8XVuZ0LWxyI605pUPrHXkdvoqOoCm38tvjoHLrOmnqik0fG43WXtHrNQQqu9j
Fy+xMhHKPiBcNsEd2XpxKAUg48MlWu+wnJdgj7zpRtWRXG+6+6jt8CI91MqAsZfn
F/18xNsA5o8VuC0HJ0gttazEUYFLuO3KfFhRHHOeLSpIWGwFrpMXRf0uCIsK5vOl
HNaL0969FJraeCBsHaoPyZtQQjTUzdY4rFxxBZ9Dk/3e1cYeLnWgGaeO8JVikwCa
nWxzDvs4yxJZTAaXO6VdYIbp/gFmJQqxjSSz0GoCOuCBeususpgd1JYvfYD0IC3c
adQ2tURvTZvcRBvDQ7tsWohUQ7adeM0uNhL2iim8ryEYsEcfS8S6Fqz9GksMHg3M
MjP+pW8SghhjGqLT2/IC//qTdfzIrqPR6MZjGKtol+3crizVZFzJQtpgOpJ4c0I3
Pjvk7pOZVM45C9RTZxqxqtAaX/jY7q3Ee2GYbBevqLX8pY1sHr78zoBz6QFYhWe9
JI9y5sDmWhXSXZ6ovlsAX+9/in32Vc7xmoFRGt4ySR5YKkFAc6RIWyr03zJujWyR
c4Gfmtoa6IPqkTZiNdufrgE8WjMO05nYLTIhRhGaVX+Ee5VMAM36ukLeGfwB+GGS
p2UZJegjelDuId/xaiv8DEh+dcqvDloIOJX66GWmd3g8TZpmrLFYqQayriMayKHo
kr86XkSEgkCFRvWCplHOBHpwqjsekB40wj1eQeUp6rGz8CGC3F0hc4ggo2G/H7Bp
g5+9RHcz76ekSnmMVwI/pu6FNwijTO3L7dG7k8G4ql0hmMtTm1gNEAsN7Wq73YoY
X1dn0/lhr96eh2IA2YrpLSrP1Lo/Du7wQb/JTX09X593RQHOiKGWthzhZZ+uDKS2
W8Z6ZgZMYb8GUZZJml7gEk2J7i1ckj6teM8gZgFoa5czH+iNak2cDpPP2f1x/iJe
vPPc2ZpnCYs5UKcVocpIthvGmp2ZxyavVjeDPbliN4XxCcZUTAWJL3w39LSalIn9
0R6Kzp39Koknqp2OZwa9drCq9Fhs5DxaNAbo11JtrAcRxiq9eoMps4EfcqljOMdo
pPMnJXUgDG4dmQ3bw1itujxyYr/ixLKTuf/S459G4gAZbDdRN/HeGXVLv98xib3D
uWhYbXXzkRYLawz36pb2bBOiFUP3p2pthrGK80hae5n6fFMQnwXtC4i716BYQ5+e
Os9kt5J8Ea5Hp47ZQYnyi2cxzjuAhBcTsc+A1Zst6qLwk5Nk6/6IbvjsMiLOES92
bWPMqWs7rwXn2wLnpPAiI7emuBmLxrzG72bKkCns4HoURDmgFymddQX3COmuZtIy
CwCnfz9+IRdvlVPRne3/S4JZudbZX2Av+0RLKeXNy7y/NLtDVZwEd+hQgQww+O8p
/VsIwcg7gGi5Ogn5X9XdH6a6+j6/xjuPRBmKFnFLqCGWivNXjPnqJ7NE4Y/DlNRO
5do9bJH6SKFGQcqu+S6bY3A3H4RdaoXceLDWl92ZmMOhn7+QBSR2+o0+6PYgKQu6
jije52oJChIyS9go2/Rzk8fnL8qa1YhI+WEeOUvxMRTWr5xnkNREJJ2uPpAW1r5m
pEJjuOHOFj4XA6lGT4vQMmLaNQmYEh8nZBEgK00BXoK5au27L0/9oKIWIC3Xn1YM
LZrrUAydCP9W8PKum63/oJGMu62popaDaWDJbwXR0DXM5ZekYjSAOf0R4rOWDjhi
0Lex6myQh5NjQJTj+MhAcBqOsxPWrIaA846AIUP+adEDmxxX98o6jVU28DTp+bnC
Bf3V6t58NHVCUfr09Il16dQrX6JYy/U4WCG6UAsJ3nqp8T0EukmmH/UZeATT+id3
dZT90o4suxpTbSlinfW4h3jpB5JfzIsZlTTDQ1MA56qqtDFp5EU/ArF/w1s9cTKr
QqSs5Kki9NAZcR4Tk/0t7QAPLY4D+bTt4zh2/KkDyvNj4lzfSgmnyBb82dxcI0e7
d4o+YEisuBeHEar4qqJt1KD9hKRrGOJeA8bWAyT2JGmfpjmIBwooIJWIvb4eE/B3
mQHkOVO97/VW+O6fenensKuz/zlRjpqCFESUyg40xE59uorTnhy37qJDoy51OHvR
c9M/WeKGQHYxpVEr639iDjg77zGY8m949nWjcaFJGD/mFxm6Mzj+/n82LE3cMDnv
MGuDD5HTLC/qqgWluKw51jDKSr0gn3Rs+pu4YGegZHURg7/faURarKFayWqttZPr
5UGvca+q29rJ6wEoMbmitw9P/BgKtiKmogPC2wNKFcq/xtESfLumejFtNIRC67YW
LxZcSMMVJAyZC2tccM8tVqMAS595UmBHte7oO5sdq4t0kZYyWAa5ZW+mY+I7W96G
jSkt52b3XodYJOXmixaIbUuWNb4C+fJAlv5OMHAsbMpH98fwDgUeMo8lgJna93k+
JYNfskcH8NInwPzNVNeWStCg949CnqT+NHnZBgzuIPNBo24NFMxL8SUWqk+FaJCQ
LH2k/dvi4tqcocp07xJTd9QIR6qBotB3zmHiNb8FDMYoRMfsBxjS9oiFHnt6dWnB
qjMsoIuVIuyChzAxa/5oZEkds5Y8m+/4xCAOyT4UENgPTteXJqG7/8TkUW5FKEXO
yTSLnsAjalTBWzl6kVVqa0OKOg4T7FvxIpIiE2PgfNS4jC+RTOGBPJLD4R78KJeN
Zo79vwt7xQ2FrGhYMRpjMFl4EVCPzE+/CUuPzkfZHG8RlIwVa2NzMcOfwL90/d57
hqloCrCspnT16CZ3oJ/zs/nF2Z8JX69lGBOQiAI3RxBkRhiEGgoEBNQgJ204VlIf
wsRrD25S9mvI63ORHEAs3jR7spauFeErl/YCWLyT6pz5Y+tc5GnBUgyJ0UEqjS0Z
evvsIXAPYAtpz1ooGRPoldByog/KNhFz6W2WyAo7PQx1t/Axp1Wvn53/1aOpxCCB
2dDhQUeGW1tSecSfDdNpZHOFC1dTB3GB348PYf+fJHXBdXOpJTq7M/FkaKsQ4g0j
ch1Eie9wN1uLIKQdvu/WTOfyzpES2O8c0jSmX5a3FqJpQWvLCMTuLOD94wi9SDbI
28d2Dm/A0foxq7+Y75T8RwVLPyANqDVJzDTJdle3ZOioJqKXpYYjR9qJhPnsdKC9
/Fi7AyhFj1D46rCP82SrvGY11wVkOBpfSIfr/3YShX+yyN65xoa6w06CtANZOLTn
aiq6PieWX3CvH1LYgWT3fBX3xfiwPi+io3dQKxshjAphSNvK4+bXJwiJ/L18nS4R
GXNHVwgbrYPoEiYC9SXLr3v+2QDjPHE/VRUQYF+mYVxvjoyfSsva1qm1/P2NoHAP
ph17C8A2N+zxcGZS63RTQv1phuqF4CQN05GuymTwCs/nFd7BLxuvezjlC2X0jw1H
mPLFqU5p/ZK7CCjud9po88Ves/5v9WWtjn1k93Scf/kQbioJh3ZzF1EUbqyDZ+rc
435mNtNWe3GUOEPAzBoOcDiV4QHmhWM/T5UiZIZH29iFKCbW90zhkG/Xd2R4H1T1
5Mt0mX5ZRTXlFYNycCn8E7HYKUSvi3bo6NzeP61rTUd8fyN6bjzbpGP13tegkR9r
3ibewffCXMxLPKZyI/EjXzGSy5WPCTcg5RWa5K+e0Ou3hmM73PbZAmeQJp9+J3WC
HvSQxxf/32gbjoXDONmIUdWJOgas/+DUQk7R1g8okvKs/8zsmOMIlXRhEvToNXxF
+lWAx+mAhG3jNkasxgWBC9k/aygkRbocGEjaVV1t9ZunXXe5wOmivt56FWNnbbWl
22aj8KfU5TK43ZrdgN/E/dhwp3ZrlP9eCHRcCC0Wl1J0tSUloAQ3jN5it95ZFdkt
DGUS/RZw58Ln6MpbtpLpWNGCEPOJi7ElulcUX1nGy9+wv1XnKfG3Inw3tGqX2Qxj
IFvoOMB28vHIJaaMNwenAIzN6Lq/JtYSw8hjmt6TXf0j7NrN841na+s0LvHxpKt4
Lmx6w+KCgayzK4LvxKc8SxMbGM4FQV8MqOQb2zixbUm2XJeeDCKCpqp53oMZ93CB
oSUMoi3RWkKdsJUbAwpl+OzLtfQHTjaKP3SKnzX4hDX3jbu/TocD/o6+92DIvMY5
5ukjgWth7LIr7Q/kUFeuq6rU7uRjSfL522X5I+mt3uLReyB1EXyt7DpLUXQ7HDN4
GQRQjpdXTbf4aHiBwO9C6Sr7JsuGiXR6b4vYYpAttsdMJtadT2dliyVECzpKzuCG
p2j3Czhpqw7hhD1MZJ4PVncGN85yThdyYi5881b4ynvtzh9GZEq5rTiAYCy1ylat
Lbk0Ed1kMOKxr077iA5oLmX8FdK7ObsFO7TZXF15EwLfIuwb5/9Olcgf8O5ZRdBf
d3vgEm+NL3zvCj6cwMD1fplDVzFU3EsSoNF+W1ZZBaAUlE8YieY7AOvfMV0dQgZ4
Q2NQ4R1GdNDgHNfoCmt7as9lRmCQoaq68RqVzKmzH5qn91CUKG7+HW3vPZp5oOHE
8rGGH7A32jBzibE7bCsTFc9e0qCo5Q/NqBG5vafKkcrxArkupGxRXqhgGGJBrbwS
42YcZxB9SByAyQ7S2X4RG486Sk7gB2gLLS0N5ZVLgEnl8qE4wTaC8histuem1mYG
WR83ksEQlWM8lawCEOL4Xm8S/iGNHEh3JteFc6eVCmH9KCEUT5zZue8wIwYxWCUK
3gT1mHeZu4JW4BjkWoIljhajA1mnOBZNN4mFpQignGkwCXHHO4P+CMVLfWAGrxCA
7PQEiYUh0K9mgE7iPGZQeugd5YjiO4p5KER21Sj9kJoiSs8vQ50UFAJ/HW6QIQfu
8FnqEypQtgghScCZH5B1ZO49vCenUQvoskdgFQC2hvsuvOgnJm7+OI3Okflt5r3/
TA/7+Z9dkTjjWWLiPgJi+FFez2pth0/BD2QhtPFGYhZLrl5MOSX9ZdsWnAAZN+qq
sQacvHh2t2paQq2Tv9HyxjZnEt5yY1+1N3SHtQXCLA3aE3XjPyZOZFeR1fEiDfLl
75kcYlWiUTVF49HdY5E4086OdKvPSBIleoK4qrMIOdKUDRzWH2ZaB6P/9y9FS9Lt
y8/JvzGUWy0br1htMDqQkNl+eZ3IiJfNBuQ9Uy0Rf3wSo109SeO2b2EUaHekopnY
SvA8vwCvC0MQUIO0cP46vnTzOzEnZX3uVKcY7EHcZ8fOrj9neFjywtph/cGb275f
IjTpsoeVtWamhV32t/wlP+sx0y3nLTot/5eNhvwAEGAaSoURVHZYM6Q5QkBSMw55
yZtXbEkA9p8jsoQewKBrMtYxCOJwhAenJZUZ/mv5PIxsN4yCGqXveNlazgmVsdce
/Ijr7R2zjsDQ1KR1hfKUYilBf1zorJF156aNiRlGKbmntxRkhIyLCo5VEs8PZxJD
/RednmByaJ2pQo2GQefjOkolo8eEScNEgP4vGzBpH75E67nDea+WEt1/WnyHFISe
Sj8B6z5o/xOqulRiu3AFxkL1BGTfnWOKFyfGF4FkMZzpbVq//J4fNGML8BkDOyOs
9ntM0q2+9tMWUWL3OeDYeNVzj7ZK2mvP3fT8GGmYlvJgB5BntASfOV4kR74EV+RA
564v3H7aEqELUcVfzjM8BQF2j34/Ccn3tsUOQASpyox3AB92k5D7fj/k+cUYNZ71
uG4mBrH3iSproH287RSS7SQ2NcF/+U8UQYz3oDYYBTv0iOVTBZSIFYpo/mhjVvB4
d5X3qfJ4JTVFIKWchB4NHwwXukdRuG2MwXygzRKqiJ4oBd2VBJnGc8KRqF5xwyfR
W+BCIH/e4cstIrIR4gU+5SXvQew/I6FmrSN4X4x6LG7Hy70ewQVthrCcAOI3niUM
DXKPtbkND8gqCtpTFPp/tz7/skgg1RxEwr/FellG7Jm1+ypq7+NQtdPxZ1S/aWQY
21e08SzU3qXUOXIABIkIz4hmP0n8nFP/sZMJDv0mmJ+47wOWHpkokCZx7VbIH/Y/
IZXdTnZmNGxF5Pr2XtFXiqk3ed6WObCnAMawALWUa1bMaTjA6x7PZ9W35A9Rp2tj
bNxhUxLWDUX3B9p+qUcYwzKoBql85CQzwKyO4yflYiEvMduYbWXCtIahOp8nulSG
oL3eXTYy47ChQ7ujTFt1j4UQuDk72ZpCbXhNZsRo7nWvrF9FZaIDLvM2V785gaYU
FYD6zERZzzg+506BGSEzfEZq6KK2mG9DDMA9710swg6zRnHQqeL/6ORbT6O5v5NI
8pkMF0mZzvthm1zbPWHZX7DHwtXtbzr2GSDnDBbTgihJnyYA4UhGE0ESkDumqvqp
znFp8N/II5+aS5FG4r6iVypdNiLd4hW1ZUFgQw6IQHAjqLbVwmrkHh276SvGzhC7
5s2pWstQgaFymR8JabSueSZzHAZ8FRiSjuVC43jDtADmJdKUiCdZ4CSThc3LKiAr
aFPDjtvoOsQTfb2rGqTMGZK1gcdbC1f/S6ovVoiPZSLU5s/8d0IjprhCFIchCJ2U
RM4+XSxDWHEVA8dJZ4uCp67fH5CyqX6Sf+Q/Lf08moEere1zzIoQCpDG4nzeeTfo
RVUekVoHOb6cv/Cze099izA3jW8LY1jhxww3wOONQyA6uTUlq8nTvYLjMrR4cxQ8
JobtvHQQkFHZAN5BPNuitnGa2Dhc/3/tElgp69YUzL5wTYZuSL6LW4gH/bbnPZNh
kJz//DhGF06FGLK4/sK3ffMhvFMgMeC+EoEr49ZdA2Lg11MWjvQj4nBJJE150Wjd
VU+CwuPG6wSMPdLTgW+bCyqKMIZtA0acdx55p1brjpJTChFfHoASgMBvsBjHBB5T
Q0hgC/wEf9sSghLZ7z7cs+iKb6l4FuacIBxp1SZv7gZuIJwUf6ZH5Fm/xEbGW7Zq
N55lvldKQ7A6rPfcR48sPAQCSUJr0HIe6Jz9PK0yGJpmi91esoCR35X6mXJSf1di
V3q2cnDj51GqXjXsyoH1+kugcz2KaoHzsi/ZnB3fWlkLv9V4a6ZAR4QOX04aq6gI
js7AL2tJi4ryPOrkxhhAvUY+TKzGmKpf831FPtIp01WHAaAQU8SGwCj1aXcyrvvF
7woIoy6BaB8baGRVwfnkULXrY39+ICGPF46sepYCcPjRZMlYCcTzOj+0HgvsY2RW
RANm2aattY+HVvKDPtp6N3vjAkKRj/ZE0mebE3wF2Ze0fpJ/bZ0XR9MYIcLxiZIU
+/qY90vxYHNs9+5NwAp29mu6LMpH5AK8NxWnC67M2umPQMX+RbGK/wCaq8sUjdPQ
0OXdnl4aZa3a7GMgPDITMWLuev6QN4889mIoSTCFevOVSv8Mz8PKiugJ9A8gEiMY
tCb7GdSyY1g3iDah45+/bkz/0LPllyo4EZ5NSF7BTkrl209WJBkSb3WrN8ANXN5c
92SU7CiadIMfL55Xa0jzct7dwYsM7RBmNtb2QouOtEz+M7KMYzuDYObcZMOGcuqU
bK53pW/csXuhAKrtYeapRmr17vtwLk2yVpAkkyYV4zdkbelpAHh3ys7Fy11/Kjqf
gDroEznfPeA272Ofo3ibCi2r2tnbjw/byqdPcHqzQD6b755dqmvyWHRLjwKLlZ4V
SJF8vhdtoQLTUVj3myu73mZgrssNYN1CPkJ0I2Gd18QqUSsBDeRI4ux8cddo55J1
75ZdB2a2AcWklrpeqlA5T+0ce6TXq3r/T0vwn2aCnEhCVFtPZM9sbGvzcf7ByDI4
G7y4hqCrk+jExv+0VZ67BHXDuRpNh/m6F+P1fF01goWprvNaxBYLV7Y9kgIlakcL
ExFBtjItH9Q96fLyI54qtmzdIlfQ0th5+f4ENw1LfQAt+TnFtmlYsGqvCTOn2nSF
K0e9t2XHC4jySg2TksDsSR57VZoHIXCq0zFb6LN2smwPyyLnVtPBHwzXGjfqu/gR
jM1iPtDzjDOd9RRStAhKlWgH8EHdLpYPoqqGnQp+J8BQQRkEgKVIu9zYXe5Khcvr
PyG/h/wakrvXxNLwZX/UjEU/RQ/MpQhjCGdmt4x/BCB/yc1vj6wTSmofs/+EEtWr
NuetTSCKyfuUbNVBGjj1PqoilsyUIl/ceG1U+ImYzk3iOxylyacGM82tboXLj3U4
9YtBa+a3Wgyx8dMjAtiVPWf/yscrn6IZ49xeNl1+1xnTFfEx1GXXVxNl7J6saVIT
E11oC7TqYSHWIiWtZ1dsXdudqARaFgb0gXK+xEatJGZbwYttd8ENcIemaCikEu8Q
AEmGZiEiMPtnxJv4TE09Tze50bfjB5p2gilEnnSrx51y6TUjVcU4UwFrECllOS+v
TXZ1vUyAd+4+F2O+oSZzAiMN5RCU4adJlJGHV2ty5i1dxjApqj+RLO781vj+rSaK
xnFmB1xhCsEQr0ays4unVgKU0kFwWyMcissYJZTY0+F5sq4Vuug88/V/J9dxfIRz
+s3YrcNQfG1c6UWiCLiB7Tv7XxyHVZy6BUpyMBSIuRYHVLSsn2dW1NiTQg/oRUW2
HEAGMHB7m2juvjrT8S+Tr+CUnffiG1PpeS+5SErtZOYQncfwrX+rPri3lLbu67rA
Xn4HeYOMYWUxhoUjS8cFLr4Vm2Uq4I4dPLZBo36t1GR+hq4QsjDa32mlRqgMmrI1
MRj1lH3hGzXhjEqVSq31c8j7v16y9m0oBwbpcbzjHxx24vqH0QKODuUy3hg4SfEQ
bchEl8UAYV+lu5EbgmZ7anxzuPsdJkrdfBvwKzPFGzLSnm0XEeBGIuVEPn0djtdK
0Rp9vqZh11RCRRrZhk0Sjj2ErUyAe/HRMplk1RlmW1ufhOUQBhpoBzlMNxiImxYv
0ufe3qrPg1pTj8Bn/JHB7+W2RaKMHSUIdfwWZfMN8UcxLgs0oqIAH8tBDSwrcrcn
JgRo2aaIn81IgDVllmcgh4NlNrII336sC6fw9R7t7Vj7y7vj91P9sBFxeLxefavI
xoOZZd/Lewt81O7cURpL/1wEcnX3K1qDDcIR9OcfCQaMghrbYBVKX1FB8xi72mYS
9fcIx6QFWpnE+6x67v1/s+1X5L9T7Wv/Wr9PtTFlKDRWy3nrfcAk4d9Ge9qOh97Y
HCUEPxWoTur8aeyOEr4VY3xZZxzFsdY190L+/a/v8h1ULsvOPjnDQRM5vthFwNRK
ESEH8CUtXU+S5BmHw7ZpbwJ11eUEi9tB3Dl7FUYIz4OoP5lGaN5GnMw4WqAvSbMh
uYBLdn0NI5bdJ3/AzBZQSmpwMescBnjKmvAs75dVOWMFYsOFr5N8bi1I4FzNjm3e
kQrTeTZ0PKV2cCMOLfCmUF1udSP5zDmoUkowTDVR7mYPaG8m+u9Bsnix4lHI9c0K
Agif7ftQo7JnHuZhSZZFU9l2AM3KfrhD6Hq2eMgIEI52p1YMKOgZfYXxEuMOyOx5
hO0RQyiIww62GpwQ6IVfe5oux/tYsWWQbbW/191c9eUsH8mHDDehbSYEBGK9MiEE
LSRTVf3kWVfw3EB4Slze6f0aQAkEUmKP4NzkEr1PlXdKe3XTXPw/rBwMjDVc2yjK
Xi+spTliZRcfbKFG4ln8b4oPv3rDvGdvZh+rDc8lCbIP7jOl+Jy0sf5z5/RaacvZ
jQGpMahkT0i3ZB7LxKdwCAtVvVvjiuWzddv+vl+CXeeB0Zf+2ihZXSSFxiFJuJUj
ywB5Fq7J9Kmk8RvOiy8LnQQZMl6hduHZVg6Hh7bdEkbB7XKKg8pBGbeoJFIUg1qV
9Fmuc64O6fpHr+BuycY0aD9sBgcY+TnRnuhVJLz2p256BQxLrL1gbpmShjozZQbR
HsLntUzUVBXjJtyRViQYUjyql4r90Qzx/bqxn0w6JfT1DfTeljLjfceRfzNO5k6v
9z+bWRebikV2I1SDU6XgT6d+F0DwoyD5jtvIhXrVzazhrIa9MGDYgS2vBF35PFDb
S0jmop1mY9GCWrJWphjqlJrWUe5AoQS6Wt/p/W7KxVhmIA+e4LAVsLQVbiZtMwj4
bJCvORyoFshXCfPsz+s6yzIVZBSmfSHxz2CPLrvGbYI8l7lJD3D9kg/jsrsKSWhS
gxJuQwS4SZU5YzttwwGxwJMMdka9rIo54nV9RKELgITv1vAzo1UN45gObYuecQAx
k58RlhJ9fGYS6gO/xcAPw4QhI9Nw6gWEK57aCl637pehv/iEOHsj3YAXmy5fTCpY
BwsjjZtzRqZYlfJ2M0WhsJx4a3G30jGKECY1U+R9ueTMS5ckJ0cs5zBS+ySYOARG
WQtMkV4ILNPSy9D5WK0H0u1Bd5FVZ27y1gj0Dt731Df99im3CDCg32L2lBRv2E7I
dBwlcVHgK+e9rUrJYklJ96CZ9RDAys6vWSMexyj49CouLXe3hwXi7SAiMz0zVa2u
21S3DkU4/nh1Q5FF3+Mq2WWXIEvFV3ThWHHUw9T97AfcM/WkeaizAm6EQRynwDN/
vRlWNJ4fosrWqFF/dqDpKZztYazr6RmzQOjsucFjp42LuXSuBE/pnaYE66Z1pLQT
jOGl05kVmY5lxqgTpo/S5KP5bncG1ujTfNeC4Phsx9Qls5dJocGDvAOcOCtAVmob
IsBm2SgfLnRXlW8gXL6zGlzwc0espV5+WurmNWNaqGvGrZwNQNsuWlUSzWE1x9UZ
iAbvTkR+sM12VLVWzIq02Z9J7DATjAn+C5X03NTTbeft7oH81nwjrqNopTxuhU+5
eCSHTlhyWl2VG2Pj/U9j3ZtG2v0PUEdccMoPsSmpNi4L+Jj+JaoNJtijCRNhQzzR
2FWEwGVFAJ7CZwBmyyUAy0l/9rY4OcXW5lPSk1pbA6nXXVcH5NDkLYa4sRn9fgRd
/PF2XmQUTugEzBDRWsfz8Dedh38JLHsnaRQX1fZSrOYKGpcYb3sZEix0lUjdIJkl
2+N4HQAEHTGfr15DydhbqOoRFXhXMS54N1NHiXVVlfOqE3e5ftTmKPbSVBRlg7mt
q/bK8kg7DmHoiQbRHa7uzsKcuxz8sEdccTIAcoXz2sU6A41jiBN/YVzkeW+v8AO5
+yIKWwFh5sRQMuOi4JpI1CMbVJLfD01O532I03omyzsHP5499iBtBKIR2UkpXmdW
83DT7xcOeG/kiUrdVvD+g77nIOGRwyL8ytSV1Fp8tNPsh2clGj9vgWZezYmx3mYc
m03reUR3KR7nhMCvRT47zjTzx9Ctrwo1oJhg6AcoG+5Ib6BDjP7/LNopigNlkDry
pAzreFBJ/rGoTedKSidqLfd6VwIsru4wN1lBGYcWh6dpihJrjTrNpqptWsR4RgyJ
JFfzmHmEODCT12gMQ1d8kGxwHwWSluHlEGq7U7r7XhhVeozECV9QCayBoAJJpsLw
4bGFHQ3fc5uUIsJPKTv7Z2eyw7VzBKtiE0RyZSyj+ZUrQfyZOYiOpOxt6kJWeuHM
bSUL2yIK8qaZmIWSbXbEQO6yAvJpFile3E8ULfUGPHJLYWPjtIWcEM8CnJdDYCah
4qhuaXkp06TlP5ChmnIfLknbD61r5t+Lpms6Zj03cyuRIvf8ywUhX16NpyCWTbYa
TQBXz4+104XvDLtwzd6efiBYtWv/knN/BSBlevGHuCER38TSeAD6qLpuMpQnvtgp
WCJ5tX2Bc5FoN3G1Ex5i/d+J4GivbbCZrHP1PvCOe3zLWV+pcumWd4C5q+53LDts
Eb9IMACkKnDIltn6IXtqUXM5w2peSFxRPWGghRQDGfxWf0JvWe35b0qtOM9AIiny
F9ACynPqdQn7ayhYRPCud6oOOZyaXKQucw2v0cRXGAa6K6XID5i0pBM9fUgcWxaJ
8rJVqSiUWxpog96RRkJVbw9LOUX7Y0kwLAjJ8KfNVuHaO+/IVuQx3rk4pqKMpl1p
ucz1ENh05KvK7I7184DecmDvb6sqRWI35T+D2MDcQ5/4BxXNo7thTY/fCNFnuO1K
EpJMzx6y96vNVf6cYErDfoeVbaN0I64g3tHBTEK3HFEsdMF4tt1YaMzU8WyGXn9W
8+ApurSvGbxiFCIsgAFgpWsa+OJCnSFg6qDPRxjAkJmG/XVTOYF2A3nOIsJ5YCU2
S9aCkzYozWuQg/wvqGtNHJRPi0N8/UuQ1bF25EczvfRoCeeG7uwvTtfNABRI4oEu
ZpTfibSDffnUCyvs8bQ5WyjLKXb+8UekbSarzE7vV0wExG8OtLA7wujbfByvYv5B
/7JCt89pT161XOC++H5qXGWFsnvo9Lx6eae64Qh2qfqkjxOZvGCOy4HDlPdDh0tg
JLNjar1Ht1DJQi04jjAHocSAndNonotFMwB//ou9erJrTB63refnuZnp2JlALmhl
jdRnYSDB55Y1TqttP4qsFsKwqndi4rXe4mWGq/ScwhwGkTyhbbG0oKS7q3eyhxPy
81GGe1MycxbLoQXi2FOfhZVNg/0AeHclVSmcYfCmpuOqFVfoX9KB0NNmdWlaj4Nw
S5ruP75dXHVx6Im3fEUfGj6zvfxbpVXKlovsiM3RIoe0jqWQa+EH8W7e4mQnfPAq
1J/lH1Mm0P3jt+kAYNKQyF0LvLDyj4CrCjfHnRGP9lR0eDdgh+PcES5p3qmkEM1V
c1yM8nTOe2ZkVtT8CaOEsnyngtK9NyU3P4L9bf4F/CLOBNbDSB4O6tEFSa4mVBU3
/V83p04G7jDfAH/Lln0j7gu0TrP03m7k/PyS0MLbwt3pM6OdQYFOQwQEbxFVPHiM
HPsMDfqc71JHKXbCMqhiXTZpCPT8xtqzH/PPbHFBDw8BHDgM3dDYr4NKg+A38t3I
OPeXNBxbb5ug4B1DcJAcAD9V0+FvqKVygODvvSCF8bTWmQaTe/1OqHjISLm3RhW8
+R0x1EeF8l0vDitYtfixHnl3QOBny3Q5VVRtvQOJ/ZWYcBaR0MWvdftKgYHUOtyk
BgpZFWH2n5Ip4VtX/iNF0R5tYvpNMZbxtj9u4F70OiEjZlgNLiCEN0hvAGFUHr3x
zxLEor/cqIl3ZXuhV0eETMGYvCwM4OdRmSbS3X5H2JHyvBHWhuAcIdXGckPEiBWZ
+5nh+mkqNOhwSkGbmBVpzafpODdA2V4K9VVoE9zsEXSZal7oLRkA/taWd0ccqtVC
ejQVCaejvrXuu0l6ObS3FjNWNgaVqIDCGAz7sJ3ldoVgJWh46tfQTLMlzkBYPRka
Ce/UvCmP4WmiJxK3jrt8E+aVZoP1JQl4VZ1XmEG/t40zd7xdiq/ecI7J1AJ3LVBU
G5fWSe6GhSnGk3GmQ8OjJD/LEwxJlj71zIVRsbtYxQ+96PDKowXtg+WVjB+yhRjs
GcgC9IZW9UtTZ2rkv1Rr0KUwfPuU7jVfS6KWSEWDQWXadYLg69Am/02nvfB3aFov
vp/z0BZTxcQknUw1ZMxlMU6mRWbH3Eipt/Vw1IE1NcstJcnNWgKW2ANcl2sfAT+A
Pn9LgErH1UWgFSlSl7o2bnJJZ5ct/4QM5+mggrEx7mOBuDu2VfqT0dp89A7Ls2OO
7PgMtTJ5ikPECEQG9N1lb9HqPgwYntMtGy/CpjqdwzJyDPkz9f5GZnVhul226bc/
iXZnjxDdhDF4wzqczq1a0tn+zREqJ6NgbN4knug2Zv20NGaI1kOPQZiCtt1YUONd
ZFHBSAM+ZIPzM11G7b/k7Ah/SrHxzeOcnv+F0b7imfdY4sDv+tE1fg0a/j3r0b0t
IqLMFQekS14wKzyJa3clXsDVocL6TUcIt+TBOQOIrKfenuUqnTu+aGbLWov2m2Zx
/vgH91Cq9iTpcoCugkVHBP3T6rw3SxcIIZjFPb4S+26LpR1oNFymOqzmvndUEXEQ
BijtUjOcUpZhMGvvCeWlzXN0zPASqZ5auoUU/UzgV2J3BRxXUxfISCP5jzF3o0On
sJhOalqgFPWUcm0kP525KuEOztMRqozdKlWcKbBbvP+JE6e0zZ4tzwcW3Io7Dv2S
zMtG/rrNPIUB/7kP0QG2u+ty/iJrnB6LHEoKk++K8eu1lf45vz5yUKoI/x2J80Br
xmxvhMCnGpx7j3lKUG1pdV9o3tk/dX4ROYy/LKN2m6uISJ1gcMgEFPsOgQdUGC7j
MKECqAfrQJSHVfwqGdy4N4cBcaF2egqM/TaGs87XzfxgLqKpPHnZedquUthNv+WH
77myKDgdYl5VSmCO39lfbCm3y+AIdOr8d2VwGUtkGpuhqklzeo9QDcqIz4SVwBSR
Xt/8lppk9hG4N+qyU7TRpHJNueiY5+rQQC09+AlfQacHdc4GbOYaG5xEofEJGesN
yhXKzflPHi70uE59r+AtExIYaFyQ6GFpyLmuX2nqVcga644ax4FIuvPHnF7eJTxG
yV6zIRp7jU0ZzIfv5CkCgjcSGbsFLoVFrV6B8GwQH3TOBIGEfAXgAeR3ZKDkRD17
6jrsb8Uf/2hrEEMRUmg0QbfFoU1dU83vz+ddFb4c9ZU4y/wdAq2a4F0HCk8VwaRq
fe2+kWsGnO3v3kYDJh1pzsBPOGeKeetzBX4punV9WVGWXm3GrL98CdhmnSfjA6w5
n9GwIwxGGL2/o+K+vv0K/WOOFjdFKPkYG7ZF5gsX0Ft/FNkJQr8pfJRhKfC37BTL
FSfCWH6Klk/yoZV3rtR8TRmdjsB44pabtd/IAp2veayiJS2Hs9vzfSbxdYJPQHWY
LSKMn+p4GZnd1OkJGOcX77ZoLXbCxop6VrMn40FXzzDGXLYVS6GSPVMs42WEl6Qx
MysvRhJfAo5Y0TCwIU2AApXDONwbsnsBZ6OAJE8f9F1wv68aCcQUr4KxjlKNRjIa
DcMMKJdEnB0jlmauCZUJN7YjDM891w9F4fXYoGEYL9tSGQFdhn00fBpry5Cxr0I7
A5foXPxoyw9RhSeSHm72a1IdXXa+gqbvWE9SX7suajceCujBycQ7q5dDoYVgA9xm
EBUTHXIF4H3Eo983HuX7OndzUlGUwHziXY5ccuWynfY/WhlnAHOJW0mpMeh3MfDU
oxtIMJdqbkISlhECAZJFVZLJQ23H3n/JCAxAwfv/jvrl9IpPtDizwA5/4SGLTc+V
pw/kJLP3j7vYWFlMb4Bj7phPea7NUsmDazFQ4DCsbFfr2yV6+pTVZ+2OVnVY/s5G
sX9NN697jjbSa2bMuZnX5UHjoQPsVca1oh80C55+O9VnZwap+j+vCRGdzOciA2fE
GzLfCxEU5ly82bLuYr4iSjhWEvs1xrQWVYslRp1LbM04y2ol38PyozerlA0+lIR5
k+Mc+fOXFZwIG+7lavxaVVmg+2TlvDc1kmSDv1RWE1pnqRZinXUz2p66nMgwg0GP
h7xe+KewbjdMPTQV4k4Frgs6vGbClFyI81Ca72VhXg1pHrk8+bMDuZe/+43a8kxs
+BtzvdmQYgCbmXSdBmZgI5rmkOd/4ZFXXIwWMwMohKjO6Q2Y79WOdrhKCs7CgNvH
KWSKmEHA5lJcJT1jHrQhHw9ntlVb2UoH55XtWeviOWviFBJc0rRme9hNaRhDeoxy
vL9005FkMV7xPyq55xcgJOC91VP6WzIh6nErCFV1THmk9qHtk+di82z2ckjNEstx
gg3Dy6/P7jp+cDohaZtIgUAg4BpSVBVGYIkVfxzpOhv5+BOoWrWJPJxdNhWZMtuV
5rpBIgQv+9wfnvM+k3Bxa9hqSV0qKG3XrlQ9JQMtECEpQ7G3d9xg9c8wfkDh5I60
E/JVhaYvULd9idpCMTktNSjwbUMVe6lOqP6VtJmeWvk2GQ4HLV/G2TAtftQRV2U0
BYMFxUsAfKfYV94YgALH/P4HxFwHj6mnMwBbkGFNvO+OVHFhZfdVg9bCfKoHL8WO
8rTHCeL8ZEMNa4ArFRjeODsz6LVKbH+CCkDblVoFU70aXGn8Vu7EFIYbuBi4FXoP
SBmv+xD7hWea7JRomAY4D+ScHCmqVjvq1kQXigawZ1jycbVlSnYb5eWO665NkQdw
kwa2lH0/yRIKw1G6S8m9DlR7Y6y2y4R+S+j+xEfLDMeJwHzHmDA2Tl5Ro6TY03e+
ggJmhtRbOpS1LqhHmIWjuFUnXeHcR6UMvPymVnU1pqbaDzTZHBel4fzYbqe9BxlA
4aney3WjM4ZqF7kpW1ayQAKKLnyEcysTp/7OtRsySJMgePu1c1PaPKlMqXaNzDap
CsINI+Relu0PerXmzmo1YHXB3eDm267tPcpcWwpoY9itwipJD9OE58X8Xo+QaCO2
FZ6Gy+6p9PYxA2J4cCYtbXIUcTKzIKHH6RMlDKbfIjWDH8LavslUWEcNZpodz8Ir
XQLn5nov46sSNtHMUalUVhQyEK0aGxvo9SaqmCnUG4LWB0wcTfrHEYUmSj/r/rYp
lW+cpAT/9LlUHC0R1wXCKC+RicM6GgfUwloHgo16xixGiWrNg2n/EBCavVM/iAER
LZi2Sa1jOOA09e/DpeXgf/y+Aa16YJIuFzNI/CAov2UBG6ajv2NI+ct9QRbCvUoG
7ZMEmRX4u9UjwlsvcdDNlgIZLZNJB09chfUr0EPz0iQ3R2cuWuQ9rwu8S4UCKJu8
MemRjxRv+g7dDV3jHtsGeUUiwhDSGWrSjDpBjvOzJ2rjjOt2HrfnkYvmQ6jJ1wST
nRFdVrjyi+owz0uBphjdmZsPbHfxkQnvNjoiSBDCX7UtweZxh4AOFjPfxAMW+0iP
/wiwFx7UCaHpsin7Zrjo/Xsps8Uea6Rf78UZgZInF6SmPu9C9I34RNioBvBLvHtZ
XU0FTja7zdfqOtjNO4rtagyF5ugZvKpcMaHsipQkwR4pmS3VrLfJrJ/jMhXssDfF
hG478Ea8jMczQP/TVZKyn3Y9j05GlPHe2fHrVFbs7wz0uORI0XyWANraVobkEk4z
nY6cg7rkYkJKejOztmbxSdXBtOy2e1XtAsvXxFpYZfQ3CkGI8j3+omiCVkDJDui0
0s8xRZUQuyC9IDPyYw2z1vioih6CLTjT2V3N86AIac6Sn0bhnC9VQErVQ/3TMzqH
k+eBbFpn4CnXeNup7fkWaXrnMqjUx4v1IXxDY/AqdtVIsRJqDEwOGIaD+kn+kWZs
5JMtrHBBegq2VUeg9uiQOU30eTpiWf9wOAaHDpulUiOs3hUEYgneNzeAsiHEukbJ
z5Va3r8jThvi8r3fvXifo5of17ECr0yq5DQO3wgDrTXQKbm2kQTdcivlbDAuRfSc
F3ZIN1vLLWfrZZgkXuLroYdDiYuGKHOSwrUl+2q9Q0dmm2myVwcIh+FTAeEaX7jb
qckmfqhiz57Pdr24QGJzFHX3BHCKtXsIpMJZPZrGJ00ulbrZVqF1TBhQqucq7ZfP
1df0ksf2s7JrDbQFh29BPx/pxH1x5UPKLpx2ApPXRGN4tXrSoUG8cUMLXiBZ5FWh
2jaRWK5h147BozzkFTxRVKNbeCu9BbZOenJTMzibGsNgl9DivGVLwQk51Ij0j+ga
946MAWu+hUiNlZBE5GojhJ3NQx3xGjmsK2uzpOISu7jynszWvx/+nQ6iQ7+SaT8V
vyCjJeZ7zmKfZb1kHLpgheJb4Ew9uJkDKpY5t01hhQO2dvWmQtO9uwroGxs2jn7o
BtfiySuZZlzSscnxhV9mmQRklyVE1yvPIu1OqFUbRtlBU09tO5gUIJU9dH1kvu5m
osOKPi+AEXiBM7r1zeHcnI0wMtqz+nkjWGO7DvVj2V6u8gGjaLBzdJEbCDGGBrXT
kj8Zg523IzxMu7XYerx/8ir91NLnZ3EwTSm5/A1pe3dP2OAxOWjC3ES0luEsyUzr
ow2p7svAa5eeHoaLBJshFJiayczcEKrk1isr7Mo6QOfND+fyRTA0BVBmj7Pq1U4R
VhusJTBBN+WEY5lnfgex1DxekQB2IHMy504/zWzoqu83tolBimissdYmnWQXc+Y6
NDqOrTwRZQIgouGAvzaFK8DUDkqUlN3c2xxu84VmQaEyVvzVSguPq48TnMN4WG6e
g6KssxYce77BqLyjIEItHttcJazp008slZ4BxUulaawWm4Lhzz4j1t3MlSIMpwHa
GEjdXLqc2NLWzvAFsx5/GAUXc8Z12vMGRLQ8PGgTJad1CQBwMvW2+QRzH1kDAvjG
V1VC8fizj/TYuBqor06SsdFVJMyVQweTFkMUFslxttMj3n1fGhN0yGgQka7Una+5
zCKf9K71gWgC8kobB1zIz06Y+K6SzwnwV1vItfc84Uu/pbhZ13Z9yr4QTrVot6xj
3wvAD0ZSo5IG5cP0L/IEeVh74WvrBCXMDdSTNUSjUA43hDhYhqGq8lQ+fb16t+On
h3dyY2k4/1V6QBjXVtjVuv26l5GFPBUZAS7LWKC59mWgza1lVlBsUUPTTtwB06nJ
j9liscWExwCw/8ChOz51AWN+q1jyOjM3dCvrr5Ld4tak0aHowwpQQMhiJV+IjIaP
71utobcrpvLCaPsrcHR+UP/rPC5mT8Pye4jC4GBbhPi8CqqZ/WWoxcAxWjhaugim
oPRbwjeVXvPmWj+LLxZT/S3IfCKWU0mkO4tLMA2jLfv+RD4H0pFlaF7QjkMzNOMM
Q6J5dFqXvdH8PomQ/Zrk2KM9xZ/VSvPHxdc7Ej77ap/+TCNkjcXs/PQ2FdZyXpdx
+dE9CKTon5Zm2fIsnf22Upse7gzpTZ0RL8FEP3zNGzsSqQf1JdoXPvxh1EGFn6yJ
ScooM8p/eHAt5iEMHNHzskXApH/3PLTvoj9BtZxKZolOlEqWS2KEvTmOPcq/nN4F
HhLa/P+0oSjqxCt4gu5xsSEtMlpKrQOzjT23kHG7yul4RvsVy64AQ7LVax28dK77
IWa7zF6Ad99dlk863UMXQP+XAX3tOYe+Cshqp5PJlJ+0wzHyeYjbr6kZv+3Yj1Dz
joDhCyKJJsM3yaIwyasIKqDB6xmfCQPtQJCtt4/vgHEr4wSHhQR/QxGmrF3RDOMM
r2c1u3zIF/66/Tser9qFygRlM2snJ4QDPll7sGjf82X/lLflNHfzOLK9+xYXP1lC
Mc1ONZWc/eEpck9kLyR5Mca/JbZRZnEIVpGPJXziY3ytG+y2+G4gvqr2Tq77eO2o
NYJfnTSqmnA5H6OPmA9+V1w5yG4e5pIEzLzTEnooBTF18nWd9P88ZDQIG7UcZZ1g
i8YwK8uBmK0uMNJngEpZBB7r1/+vUFUWpC8W69lQiNl6w4RZcBITQ65sAADsF5eK
WmRLFY9biWfZcR+/1WsfXsMHcemIy18uSs3EzoMColcbXdBRdTlB2un/VcN9/Qfy
fYTvThJwEvy9S38LsHr3Aly0RYZMTXqdheUCPo6LmMsiCTUwQOVIb8xhaqcKUFXk
GggDjbaYqcevYCkDkn0G2kyFvTJrJkMjLb+7V7IZYyaCfA7lQ+X9CEIPvljVXNSI
QU3gCivcIlPL0/hIyd3hAtmggLilk/A0HVwBtRdBHekO4+F6NSVsni267jmm3D3C
7kWdrbVlPMNvm4vW/NRtb2+nDMKE6t1z/ZTUt6ewM86U1X1F1APnZiWv+2G9f3m+
nrEiMo8NlJLgaOMZKgFLIWRSdIuHwExH+nDK6KcpuV6uaCYhO0JFsfMW7NOAAta9
1l8x6Gk3evyR6I1/Ngb6bOdQiwzV7JROnSm1STsjCTRVJVTz3P2TOOW/Pgq8FmH2
JDdXDANuju3BkqzcIQN3CMvKhSMsy81nLXR2BKpliE6Rb/jLrsOkcaXApgZYeSQA
PW4NaRyALiESFQvhypkSTtt4V/YD3I4bRMIeAyphQvjJnBCIiYG3sogi9QfnzXvh
Gf/377uiVMYwRqU6gLZN0+tzQRJflL/y6T8Zr0cvS/O0k1reuuuM6a/HnfBw0DIm
bx0WJqZm24Bs4uP5Oe85FjV9DujcBnE3vOnoB910t5Zhka7ACjOohtOTHfj6N9Cv
ACD3sakCBaEY0s0NP1wUlqGQbTAaIvgIGurcJZPNTcbvGnjPzxMSMfFpjtvvLrhb
mmAvuWl1FgrXi9bBh2WIP4BkRGNjzUlHFKDN0cdGnkAVqUQkPS3NzcMlc6EEsUhf
Wjhv7WD/8n3mhZ9fgg8dJB8dEx3om0C8ASE/s2VGhTSLn+BMyGbBg572Ufvum6ol
4/2R7ht4wq7jmAAa/aDBDOpz1/MsLxYqagFZXT2RyesD97QDX9umXhsRbjFLgu0p
gtwDqCgO2d4o9uYupfC2OIWPJkhZAHreatLAHJY7rwY+MLIikAYl0FNHBH5ftL4E
z2IwBEMcgsSEdLIQkbuXyDN81NesEqKY5q1dUspViS9sq9AvYHt+swb+cGgiu3E5
g6BymDboW/ICbt37o9VIv2EjjTxtPM9NXfibrZTLXC/PBcN7DCbs9aAl4wxSwPG2
s5W4joOAom/OJ2MOkhwfZFZW1kjK1r4TCd+JEVw3XlmRcqSFKGJHaLMF4Igin2xt
9Oqjl2dbkjCRGJTFGlLToZBW1oOkfkshWC2ul7lJ2hkJdWuRNHkkuiTkW1H3M+p8
0mMsPDxXKFmW3y66XQ78m8/EwAEKByAJV7XyB3qQEyDvWAL3rQ4IEYZJ990OdxfQ
hNQtSOA3C62my6Jp5eK8X+Mn0BrCU/2NJBzzqgEUHltQXwJ1Zm8KKzx52J9E37IS
p7mV6bPo/EyUABgwwPOpBwqI3nL/dkjsdwoTqN8d/Z9fbZtD9zbOt/2ZCe2RV4RV
cm3ACHq1yc5DvtWuKt18sy/5HXWrjeNOy6uQa6Ot+1xwF01cVhppAxNLWtpAvQnM
ko8iHq0gRlNn5K9loiPuE9lz/EcJcK0ZkmVsWOfvWLvchmgm4E8Y8woRuAI8dV76
W2ChdZrAg5MTxyfvpskDiaStcAuIG+Q49ZscGNb52xBSGD68Cpzt9lr6/GlJdXU2
a5fE4K/SmaBNE/ml8tF/5DLkhf/mvN+IyOtuDSfPs9ahNltQ0kIWtqhLJvTA+XVc
M3KACRSwnLuELyVm4m/9UzryaIVgJ8fSBpe7Sr9w7W79WM30gPbuPl2tSu6HerSo
Cw5Q54WdTDhoLCJiGJmagpB/EloOuP1qpS4XGi8n1kxTv2J0fyvKg5rxnUD0GGVa
Dm//vNUrhEt8ZhihhEV7Wjb/C5s+2TPpzUzgupDv1w5S9mmYGdYx2L0Czde1pidE
bb3Q2TBx5L/t9DBv+MgppNHnexvQjOVQ0e0ovWPSQGCVT5UcGcNquPdG+oDq9IFa
xqPExKGwvU+XQ/v9ljYfFlFZ5IoWSLIa4TRdOLL4DlI9INfRGgt0CCBl71XkbspW
is3dISbkxdRZZb3XjvvKh9xSYufAdzZo966IJE+sH1KaSjPV0tZj8lQ3mG0SG7wJ
9GPOx7p2yrdQ1FRmVcE8aMI0qCI+OdAt39yv6AHBP4Yx/CBIrIM6m4DQVQ2qXPuv
/Nu3+pUyKTK+dJcoMiCxZBPlq51lsnJNsCkrqqViXK9/pjpF+ddEj6pMRP8XZghC
/8wXo8I/eoxKoSqfXrdT2+yqTagqR9XJ2H0s8n1gbwxc2Ajp5UITJqEykw08j3Sc
Lv6EaPTT/tsKt4//mJIEG1WkvyqPuBnHvS/9afKwVkH4YIWMmL7J9KYaVMOcJ5vT
Y4UmIfgOmlSqcGsHKhUkYOToYeIuihscOBlcplza3LEsv5PbmVhTCIIoO5TddQwB
ikgpz2cbB2wKHyX8yqRNukTaWU21oaeoujjY8mBa9Z8PbL0VWknO1IL9//44aIQY
yXL99tF7P2AIFJhZho/MIJf3b1I1ilt70G4m+QAKbKpDYSfnIHL5PoqEf0vWdkUo
RcyhqiadPZVLixFggqpA9UCq4sPYKVrMRJp+kv6f/dtF+aAsDTimMBo5wDpIQZBs
/0XK/QBqOO2FUgfMLYdbHr2+twwMNN8+n6SAzi2lAf/fANHcn9Nnh2sgftVPo12E
JhsHVGhamz07HH/6ZbnwWgK7K75DoF8bnK9NUpusLjw9RrZgktPs/jeHmD88ZTM9
P1riKNHT7sggpRD+jib8dNuG73Rka2Zpj8ho/B2HLS7bolaYsI2z9SPX0PHB9/pJ
mdW3LLAWY8xIc2btaJwywtJwUpc3sPD41A9AysF+Otw7bdW/U3NYl1B8jf7zf5Uk
6ghhSpsXZG2n8WNB0tZNHLPOaNRxFUtAj+FdaqsxNg0WwBvrW3YgthQsiRg5natq
B5z81Iv7VDBjvcryiIbtOYzgeQVfbQGnovxVKcxaQH2ynLl/7gGdr7SEzFfZUn3R
gMq47OSvsQBfaEWnNaUxyhfwKkrtl1CiEJx0bbc03BNoL4mjUBMbMRr9Go53g8xF
NHpDPmflK6+EVm76vvomCaL2XBk8PLqhdlIWrYIRj6Ky9v2+xf5VFs5nNkuGSUiZ
aIJrl/AzGI7rLRIOD8m3AAWotZ4Dg0T+Z14Dh2VBlH4NIUU9ozo372btUd6+7BLj
cKaAjlsZr+/WwU+wqw3t4SP+RimUxL4qxhADt8gdvVlJDqHyt8uXIHOiIFBymAlo
SgEVGk2gVf6QnE7z3ce2N3MwhpL7UZS3chauwff9pRK8LO4oiGX1cSyE19eGryVU
/CPNdy+6P4IYb74jWqOivTUoaGKy2zWkO+TB3WkMcOucFm0t0Xets8bDfWPUBLfc
RzJGV0uQNXrte1wne189JS3Ck0pe8Go1Lp823lN5kHXXB+YlWEgr6FCV6tIgkWT9
WlWEUP5vsnenD/LaGAWPzDti+OncsYcSXqgTFHB/uxBcIuAjDdGOytxXp+BQdlxN
MDstU1Rve/zd8O1qJTatevs69S/8XCLwVGOsZ++L3IgWWn1LDdGAwA4JuxFfkapx
EtPh9U46MC2+IYMKJPNm/EVyl7F4xR8ZighX8Ts0Ve6e0Sl66DZtkPIjKqeX6CP2
FWY/A8v2L0Y6v7+MK9FAyYKNeXKFPVP9JFINkkhdGulCLCIfwzCLpFyPsxYWDPHc
csA+GGNEODLI4vVsDu8hzOWU0f6i+wC+5CrDJnPwoWrI8EkKHgp3MFZcWT2cow+I
C3N6PYQSGik6KC3JmmyHmhaetizCSZMHeBAS4MM7/J00IfktOQLPoxf1ZzZOBw2o
CVd9dO6wliYhsfUouNCpWHWoSSV5c27bhpwh25JSCNrOLsWbR18S6+Dfs0OPv/nm
m9DJVzFmglWMrC7rTsAeVYSOaD3PyjMxNTbxDhMi7mJy/WwWU1cBOoODwAN2QnFy
lBYgogJkGCHW8YWvvV99frTBLI1QUjtYFgP83MF+jFnAqrvZrxk08afsn5c/nG8Y
4Z5k8TZEQgU//cCEXOZalAIXHdc9UvMCE4ypm6GMoAtrkODzliEA90R7OXjecrzG
aB/gwl7kszRdWMzy9HfML1i/VS4PTwKv6D64gy6J2bXuLTzA3rUQniuTeDXfqj68
xAD+NvMxz+U5U48qxye4Aq7fYphQEA8Qa50fv+LB1YcxgRSDY4YJkGqt5uMQHTau
Ax0FqKO13D5ZpsFNp+sEgH5/M3n26XZl+IDmThWasTezlXZc/mBZWYhl91zy89G6
E0QWnzBVBiWG9rIIMDtINuwmhLaHWqv5GptYekVamqojFHA5h8uB8U52dUV1DCto
tisLepdZ321DIrEBuBXhjiTO20FE7zln/AW5c17yGtdUI5zTiv2PSXovyT9kfwGr
r/vEAZXJaDrbJNIQjwoMNqO1uvu+xQ/fxWcQi6zgboUWnG6a9J6JbYxT7qW4Jxwe
AWDGsqHvnHtD3dhNtHXsUr+bqkl1LPf02QUhjyD/zPiKH2fNmYmkkhaiWEbb9qTt
SezkVEl66mzpI9FTy2UDkS0yqYw5xStTTT6O0YEV+Ae1TS6agV5p9l5t7q1Y0tFo
9rVq3DOD9HGYuMQS9YI7IxbHlixMIFZQ0JL4YG2nc7FqEucVPmiUltFjOJtD+M9E
VukZRZRf/Vn4uJKbbEQAv+HtxU6wBq9yZog++XDTwSTAFUV6/4pB5M124Q8RxNiL
rHcLwNdkiEr5KkEjcPvfHNd0b0PNeJSw1Be/9FhCtiMCrmqnbX08ZfwPY7FXX5zh
PpXof3+wtrztGj0mhJt/m6lV6HPlarzjJwBQPnJ1DTVzJ2U2R8Nu5gyT1wZd5OiB
G8cCdJ+xkh0oIxBbiMx02mRByKJl4zDq6JS4LnoVrXpesarE59QJzZ+HIOcZ8C8t
YFGRItrqpBg0K1RhE2wVFYMVN5wS+bR2sSMXf9wlQFvD+zqFWGqcbZo8F0hh3zgQ
1U/mjq+za5u6JvFNo3Ae2A0jvchc4cjXddMWsDaEdQTOgku83jDKLZ5XGtC+M5mA
CbKyB1bKPnr14B+XYtSMF6cPDu8kntHXA/qCxpF8hTuNMk/JP6s7h82/7W2o2mwP
NAAPy6OZaP5FtPDE+r+x1PpDNJAfEyxTGITK93pURCcUL6V8M2my5Ezl8ncd4ASx
k1rKYUctXIu0Pp15yTKEKc05qT9GieZcQe18HBseaGMf81iIja9/FFZdTAZEShwu
rw/K0boLDtWbjNxqpvXhY4ucOHITHDGyHxs+Pnwgd4kMXstK8ussU6AHzVEXBIrY
8zTTZbhG1Hfao4b83SKtUBAn15SQLEoMjU4dwLVh95j+3soUX2Qu8VhXCT/cE9I8
vzEs6yonng66hHuRIvjeKssc5+Nx/iiowmv7Xh7EL7owuKp6dKmu5kELdcugRavJ
fVKvx8VTAY0JGXVD1KhLk1vARw7sSQ0sTlce8B1L0n+YIAibjGjAZ+7sO3bPizxl
pEiTFdOJSgCB+gnBSNvnw2+d8ch8o9jsgMiZ8/kYPCTHVOGNeq0BCmkqVOe+7432
K9SZAovxyJGeVz425rQsjcxyJsx4asOTcuy2owRd3ejmfMwucA7kBmI9hJmnHCqC
XNkzxeJ29ePUZk0vDGS3KSjBSJKwDa8kn6dR56QRQ3nTOtPQ1fjRDT8TelzBNZi/
fqFZn/8yvXiG7uZKkPFbgh66YBzz/Hp6EGtMaTY/s5hZOftS8iyFmY27oyxLeZUH
kUeDJ6TjfjLk5u5+Vv69h/X6/LbkgsEPwN5loY1UQRYRXnzLItfW++LKNJTFFeUx
HjDGmYo7Yq7MZE/mMBwzkQZHjYSwgxxLakmWHPif5mpdHxXhnWh7v4Ym3stAxSbW
/EUWA2TvlGFR0TAzQyIc61HRqu3ccz6FwWPPycMJNRBD12TQC6vGq5kKx7HCkZbV
XZp+Nb+ppFmCOfnwGY4Clu0rGLFvDEbkgUQgHmBvo/LQjPHQSm3rzMU2bfwcjSVU
+VCvkuFrJLHPHmbDxnf8OTGbwoJdNUdfdawj/wTN7Z3X2icTXudR3NNw1RnIIXNJ
mWFKJXbYTsgcQ9paGS/4LLCR1KX6MON9TpC9qyxxObFL9MvHmUx2Vu9VmSwzm8QH
1K9dwwq0GS3sQDebvzXyEMvbsln4oWibNiTd6RItKI5+l4xzD71TKd4t4h1h0XIS
5UtF4UtJrmM+KpNBn2f5izU3yu8cILGIZRJmmJsgdjN5HS9Jm5lEaWqzdCHkfwG1
cBPmc7EpHaQbv+8cDw8JQi01yjava8G1qf3bjZivHWdBsRVuloCnROod5xl80cVl
wTmX6tHqRY9BHar4+ekveSOL4nh3amO9nfS0yeBHqoctTlqsKKhd85SHRUTcaT3X
RHYrbVle39zdVT4634LQZ79elCaLyxhED+NTf17pUI8hnuRn/XsR+laK6ZhNUrUx
un2MbUGIp2kCGYMoMfYMHHF84mI702qLLcJi08VkZYRxmhyxjsv//+3xjv2I7xfQ
ATN4h7HeHzFDf2n42UseHtRCyMhkQMrcV7t/m7hYKQchRr9jFJDIy2WsdSMjdrhe
7BUzArctD20Gk1R1IgXu+dLAsrCW3m5o5EsjLS5GUo4DY0wIOm+t9QMSeqCziJAl
ZQVL/ke3YDi04W2qhCPYLtKQvR1+YdiR7RXz5WIRxTOPk0tJEngWt3i0gjVsVCY3
SSr1vLZ3I2QHjhU240LhLWJ0TJse72cxuXH8vdT8Im0GXR3EeHKh4iIWcJxBbgK5
GTKN1+gH+WfW+Onei0LDZuS9QjhxnyTQZV+QI1+ANjsxQHC/2YOAbS8PwtqhnlBI
UzwLwgfTh+RLkPQmbiNcDyD3AWQ9dlk8jSrrvQsl4fwoexSgFB42CtG+11qYeRt8
/J4r5Ixln3MQEd4K5AS80vN3vbMqjxSB1EGsRRyyfVtl36Dmwz1cknUtre6ESjkO
i0H5OSa5JK9kYMGqMR4dzaP81z0zlFl9Mmfr9EKBLH/TENSExFSSZ41G3FmAsMet
uv60hmUGD/UUtNm9eGIyu1pDtc448ICLW8kG6xm0x4eZATMXzzKy/SV+1aQb4jlh
7ph/FmAbGgv0W0ld+43H+nfXObjd/3ytpZTRRZMF8PajZSvXz/DPudlVJ5RjgMmo
znvBbr8fj8lBi/A0QuXx5+Pf8uDfIO1q15KfxkqYi1JcN2lOkNByUpwM3vtJrCDg
lsP7P1Xzfym8i98POzqquartofCdZquedHZ1wKGsKp4nzUHRZK03NgzuZS4KOe61
bCd7jJFiALn4kedg4Bfx1n4xXWHVpTdgOQqUV5eVPI1gHoohIo7I3lwmvqru2+lo
RRPI4x89IabT+a3Q29dAoLg9ZhK7lcTC7FXSJACx97e8kr1N18f+63uSJcPTj3zA
xyHdqt3n/efM6kWWvryPFGRtD9DVwXHVlxxq+43vqo05BbR0va27vO9YH97eT/0p
v0TUp9xLaM0QR/7lccOk0YbNRYUWA00b/h883DNsbp4HOrlFV0UtxBAIR4eCjLMG
BSBT0oXNM2khtKYRInRxRhOSFl0kDldvbRld5htXbY13xLYxcBRG+I1V6fvVIgnP
HSLRun646gakLj4mDLfF/Z3hSmY0x4rN3kgXlHgVIm5qQmeC5BHD7b78RxpWoYs7
L1AO3BGjMNvkRMxzS7ckR0WnVA4VC2LoRyRknc4DgTmrqyOn6UMooT9eJdD9P/I7
MSaASxe9+3aJDRaS/65dxCnS4Bm8JQzVMQiZJOXkhSzK+FMeXWkQBhM/Av+2YzqJ
6T7aNFSB4SKTN/QAUf+Tqvy12O8Frv1HIcTU3CIaC9/O6DcjsKp3j+pyi6gdgOYe
z9/Zc8Y7b7G1q6aikLoRisAg4zTcwA96S0PayBhm9QO2q1ZZIme7bN4dEfPU79i/
jBQ8wD/2vAw7sBbJjS7i3amZl9zofzi3LkvkvLBCT2rwuUnijo0du8bgL5Q+yF9e
R2TYAKH58XoAzj7ZwT83le3tKgmU9vmqpVkOluPmYqpzF1iEHrZN5pnlV8MtQpkk
b3J9JGGZCWZwrYhJuXw8OBQl739oRIkilrUDx4V9lOiAHJhqf+rgf2j2IhGBXXAk
tO0CVFRvxGZ9aA11lQBxd6cTMt6agWdJvJd3YRoRH6JCcFPwk/NM8Oxeut6QEfMj
lN7N7SKjLYmfhjUQepmH4oZ9JJKfN8Rj4etaEIMKmWvq1599ffxpluUbxQxaoh7E
mD6a1tK6cPPvCSv9NMOFbPnWdFVEvr18HNnEv6syW+nxYQGB1N+3E076eBUgaZTA
dsQSu14z4B1xse1iq4RP0i3lT88Kb5qXzsml1PpNFO60yQUF0riT0U4hq6dbYnBI
pgRR37YzqNf2nsAt9VUkgpvOKnZzZk/FeU95bEbJ5oYvs41b9qBIiFmv4JxUO4ye
T0gQGYGOR0ZYghBVzgls84SbV0g4mbYRdpTfG+zjLgtVScQCwJmbIBUVD9TbIvXk
tCj2A63xji5kJbaBFt5V/2YTAVXzk6Bn2GfKnF97VLKgWcWZQd/yLc8yOGrHxoMR
yEqllKZ3CZSxBaurTgJOy0Ef5kUS9s04Dhfa2nuuaJmB0yZXayamq+4JD0jd/KJ5
T/G+euIs7uA/oKX6JVy4GESifd5PHLOUVadXFBEuzeVX4KHbzLIPu0j0rYGYSWZG
I1JmQ81H1+eiRgIBIs1MKWNTgSzfG0/+Nga0XVPV4/IQGb209DQja/q8baW98djy
L/gVujWwC+T2y5wRqyUvlLJGd9SrWej4G4H6xPniuSXaZVCB5PMiQZFOuF59qyJy
UHyDsyUwMWW2Kzc50hIRnGFpY6z76kqF55LrTHlX6LzE/fzJRlU8vsUhNrkz3pZ6
Gq73JPRqQxJXZuZ8xnJyIoQeM+pBWp/owIxHGRdjz4ODt8STAXNgTxpGBwtlQ2+L
OhAjLfrWwWRgGd+l9nHso+GyHiRv3GZOzfe759X0krYamqaKooXrwRsY9Kg/m11b
97dSfT2ULI3uqkoqKFM1hsjFUaWRyoCSo9SYBIkc3aiK1h6uLPUyIyk1uFnGOuHC
ZoTOe7A7asgIsZQ/uHNSOmPqX4iofEzEbwyCdCIFcOvLhUeb8AdsjDa0gcFlkNX6
WeYLFD4MbIwDPKdpxgBY8dgEkQbbc6sj0EVPQGJBuxq9zsBZvKvUKzqU9FoEdYDd
hTSOYeyqyUWSV1WlZkk/9g4sRHhCYBJ904DpaibJZY0E/rr+1enSc/9E3KJyOH9e
ZYToe6xmGqZnqVrTzrG8KrTFCXdI3WirBjl9PUNYDKwkd6RTtJeS4Siuo6Q+S4JA
bFXgMRHAHDTvaZwGsUYbPQP+HWbO+1wDH4xHZUqfdhe/XLgYylGdWfWI9mT0BUhp
+7EqGxqGcrM10zKBZOS+VWHge/Kq4awVUu7hwbUo50BN2pAS2wcq2hM22UzDhT/f
EQJ5yVtkGBIjG77M8OuWPWT3MkOFh4geB8kFcbulgwvPS8kRQInqr13PJTZqtTsz
um9Mwy7uOlZ17kkBlFBBxWxLuvGcPcqIp1on1J9RYO7bd9sAcfLz9A/aBFIZWBcm
u5ifCeUUIHg2y7Oj+jxJcIRXWiJQMChHoKBkVPzt3WtFh/S9hhtFKNwgJp/jK5X3
N58MRmr7UO/U5cHptU+QX2Vyx0kbN535hSRBNyr2fqzcyexTzLEMtpCkKRLrluaK
dUWNr7iO7aNagymy3qx58PJrDzO6VUOlaos8TTN1fpmqimR59hOdOaBZCuxT0S29
Vnio6vsbvibYN3dbOoI6wGpf9UN59/VV0G+2r6872Q18qet1/g6dB0wvg7G67DnF
dpxnxYOHMdxtpPgNHDNI2Hgg8q6lS/o0KPp2d/HnfKNqzbPhhCoEmA/Mbh4MMZ1J
m6YlOnj96NRKZMfnS2Dg/crD9y9boIt+xnXNrq3z4JgT7jUw0Cst22eaXD9/v/KC
jfXnFHi2C1GO0mJdDPwSCDNcV64tZJzQSbV2JfkZLRSciTgZRNeHFWKi/NzPeOXs
X4A1xeumdx83bXAqbLOUCmUoMpdD7yQWTNnwh+6Y4xIOnvLTAYIigy7o85GcqDv+
K91tirnm6hhXuVidQfMCYVqx0PUVl/E+iL7SJtrh6FWnNjdCg+5xAFQ8ZtUc+9t7
7w8Y8Lm6Z+11lxt37fQYxYD58c2h3emcvpZBv6AX/NX22aZNJ5sYPE3eRFsNY7Sj
xu/fho2P+tq7tuMScc+DUcVjH1H+k/VJ6FMKCnqO3Uyjcof/qDeUcPmPrUzdITYW
BvuDcWN3pZMHs6AvMWiQGTQX7CZzH3tB+OvNrfWRemtIeg2+bz4ks/Q4LqAq+Woc
tMz2c5eIA7FxEIzGO6DxCowGETL0XoMh3SSRg6RFQVBkbUqnGIKnf95xK5DqQHI9
PN21sUxeZTF3x6CL4iJgwuvgz+/7Qojbcv6IBXxZyuevCcPMsZ/GmCyO5VDOiIK9
f/WeFZsHg4VOtV2HdXG0crNcu0G32EmQk96j4G6eG6z386WZAUfafGG47Slx12IT
LPbml5BvM2/CbKouMt6KLh/hHP1oMTrZrBUogc0yWgbqgWo7QVe3XPENJapQiVIs
HLU4stGwow9BM63J5wh6IW7nBwRNX26JI4URCIVrNgtzvVGEyRPwi88hX4k9hsDF
/qHBfiaqj5UTix+w666HgE/L2dQlfcSf4lOU90t7GXQiG9aHWedOqFPFIfRp3VBA
TCm0dW5jxYcQKEhrje6yi5dFGloTT7kFRex12DuXwLNKSSkRrRxjfBBVayuxenMx
rFuJ8GO95rt11m4FgkvmTKC+bLRbCNfp6Y0YdVEUO5yaGqU6hB1o+zrZijejRdvU
vp0xepQm3vVwCUmLehVaY0xHHUxK/aNv7R88Kto0B9dyiWDKbfThokox82gCA0Ye
f3pF/CFtjGsWYaAJhLqAuqjAs1438Wp9sDkEEXeAkXc/le7VOfUwILdY7TRRnI64
pd1OwFESOJtFn/LXqYvCvBXVwQVl6uj2qB9EYqOm+7GZkMg/S53HJjF9GKNzaYoV
2I1dB4HaVNwaPkIcZ28AYuM+PB6I/5pqyTaB44OC4MGZ417ZME9nkmF9kju85Apo
RPmUpP2H+wb2/KymWOEuq2KFkKphhaTcrHLDdg4K7xgkWyXPsDeJI2o1ftZbbgDa
iiuakShy1b/ES3QNBxPmFj+MJ2OXrQG851GtNPJZqkpLdHHvqjuUxuhFgJuyhsXC
zuaOK7Vxqr6HkcRmJCTMAKHUACGf8k3uwlDIzkfZeToLOwNlAyLA9J6eIfDbRMTJ
33ZlxxdsIWGQZbBKJOnV1Jugn/Q6q1vZSSF0xyejl7+9LCyX9K0BoCRTMUl6y+Eq
QugIHVbzllL3JH7sqHqLopfxfcZbch1KNPHzgJfP8dtvr3DHCjhjHL1GAdvcM5G5
4YuOTpwmCU3O3fKHZuEH/tF/uH/4/4Qn2V8vKSN5UodUyRoy4tow9ovALLHyOV1f
cdHDbmN+Zt1ABvBG9urUf6OGvJUuewwCCtgLy46ePZLf4Kq3cN/Yukezl0tZHhCK
90UVRAyq2qFVn87b3zqhC3z/H9OOEZsjoLrkENad9mkH2np5/Dsq4TPC39X6PPvf
1sTheUN45s8ihznTSJMTULvkSqdRfbzvei05VHcN+YTPFjePNE6mucCoL81l5PBQ
IV39Z8VXdP7m1NgqnvuBDmyjTpUQ8Gp4b/sxbabZkNO2B8Tx5KK5q1U2Rhl03LCM
T+9xbWqnoposcGEK6ids+cl8pdcH6U2SEav3S1nTNhb0bN3ZFKQEvKy+rWmUaLyZ
yZVJe4svZ156zT69CwpjLC+cajpZwcB7n9ezVrd6j0F8pHV6WdRE2Q2rVyvvdYnF
fM4ZGBfQ61qAkh9RHA8i8xdHsem2F0ukxc2dSus3HQcDlFTvg1ewVf4VBDmur8CE
NU5psb8xsiggKIzNAQloV29NIqmBhFVvHZfrPCX6Xxfz/DEC6nlU6CvUNymeo/L3
KegQYoq5NM/rG2ecx8xQWfnandVGFnMCW9Hgj/2wCjWkNzYdgsNnHJjPuRUASX1S
tFqAavUB9AsbZM9j/X30cV2fHatY8fo+CV7mbRjr4uzvZ2HPUkhFL9t5wTWyWqOV
fx3qjla1g43lP4ChnTs2u3xe96C3yloPRtlM1m6/IPMFKzKccJ1kxeOUHXIplVk7
S7j92rNRcJBatLLHF8pS252bX+B0Q778oPMcExFyetY60u5yATCCGr6P8cYBIwZ9
0Ko8qrCsSxrSzaJjiZK9HdJNmfDOTbkkbYjcAZlTgv/v3JHKmS3vW1po4LGoUMcs
jKH5iFSUGJQyzJv8hTmo6br7wsE0wwS7oi3Xb0aydtZf6MHTrCAVcyw9fdGsBizy
zoHJMukFi5P6mYjbGiO0XhupVEv+JnxiIA4ITqXLyov6lJrIQUdql3MObzLsTGCK
NZbrqmJHBYSENkfwpOdEW/DrpmU1Mj/J97w4t3bT6DG4D0yCCAavmaG93owRqlKk
x1AF4SAYnBF9SByyxYXnoi2zvbM7E1Tej5KnarfOuaTCOZVzijhugux0JzlkxYwj
vKqDG1yRmDf9+3/ZyGLt91OsP79pKnfMc+Wz9yUcBU4BfASykOQrnp10UHb1sOCa
i/8e+kYfVaPJccoxeF0ZEoF3GzRFQPXt3gcqOi9I4z8KERy8vqKTyxJbLQO58fSy
Hy82z/km2zE05OyOWYNn52Cms5uHoe2WTBpFHuIZ3/SMSxq+F9d+sM0WSUSgWubB
WtKTi5eNy378cU2thdllHnSTIEmYE0PKm4KAM8pCj3RuoVQFPRY/CNMnXGjnh7j6
zUi5Lu9wLFlzsuCqAXuDll5cHN1/kRSoqoKjW873qtq/BfxyeNMzpB/OH+fK2v3l
KU/OwFwKNqfXkA06SnXqm3mO/qDzpI5IDuWiW9IrcB2FcJnoDfzwYhasBXPeju1Y
6qOEmRJobBN+tHlM4xPn1WTtm0R9jtZ6bsull+q8lAOSyvT2U82QB+pEyOSvQCzM
H3HaaGg99PMRoGpZ8g6/OQsEgSa1jYpdUV7rqM4j7lnOiaJLKhT+QVIEl7o0/iUE
aKa2UE9sUQ6H6DicoooSNAnU8WvhzVbJyB5GdhTw2vOMb7ZzZdS2284lhy/j9mQ3
3va3bLm0KMtfpY3JRofUqaFaLgODVJHYj21JWSTnZzQ9wvnzueJriOryKw/JupVN
VZEDhtOgvuab9seiT0HdkwUewa+/KhrKBzqeCuyrgmoBYjEJzQXaKn6XCH39XgRz
pkMAgIW2pZqPMjUX0/MzFjPpuLAW/dizfezftPuefnnAPU8dFFOZVwLJSqx3sLpD
wos052QpqvUuWeb5N9UkfqG0BLtoGJSgD5gRkl4sAkNgMCV+aQeEr0X72HSOOwIg
bkNxWf+GWCQySjGT7MKThsM6ZAXDHRBho73+PVUwzOpVLO5VuuVuuJxgZ1LC8Z2Y
N3V+6cBPj8JyeiEqpB0GfK+CI1uRDou7vsJzU2UGU3uM7KWxSoM7w3XNxGJdPeDW
6xVGNFUClN1o9z0c0R/qVlgGuX+djnpWkGsy55r8Yt8rBtmLFd7JWxh2T6XImjIV
QCYMqxWisYcMZNEfTRSTGf2eDw9sknSgv0IJC7JEW0MrqS9IUwOsimVJtP7oSu8T
xgo/ygFAYVfzXxnFHm+GycmuVWenDhEys+EOcpD5ZJUiya+mo3DOT4+YlM/0zEYe
JEHNtddojdEORM9JMMOZLGR322325kUynaNpb14lVg5+SlokbNqgH/XRTPoIvYrF
GEsHS3OsCGtZMF0nYeiJjW0Ij6xuUEqqz+P8vo5+Q6mDxInaUOcjcsF0gcR6YMx/
NKgvOxOyU1iFN0tpx/1cVgVOpYH877Zvr7kJb11lzdZZbslAWUmspMOdAf8tuCjU
U7JhUi7G51D3RifiXFw1zFITrHYDZhmrQCG8rGH7a/+5EMZ7Ijlu8cJnIGa8J11K
GqiOUHvT5uYkGAK4TG44TsAgXjkak1yMr9e7/QznGRPtTZLsdmul0+Ive761WSza
J7kHwkMzfVL3ejJ+FJ39TOU0UlYAGZXJDOIEeT4qi8a9X0pZyEuif408E5LKrL6Y
3wvClTydx/zJ4HOX/HyNiSxpwN21Vd3mAjNm5svsQeyLMmTt/YGsPaIRoWfbFUif
lVUps3aAzKRqH+Kbe2wu3995PyD2l3TlNOKgnU/FHKuNzkWgmQO4bPWqOLmCTVWN
7i9VPbN6LiE5AxutO7dBjWkY5C6Yw85btHhnmFHoFTTC+Zhqikqwi+43+Kb65Aki
wdMEo76YU5gWFuPkxXWZry+wYxtw6bCRXA0cS1k0RJJvmFhGnNeBOwVeMyo+8wDh
umDngaIhRHjxOrkizTJ3WKdBqe7iL4GA6a0zPn9MY6X4ykwy3te4NLKi/XeT/HqW
LSUvbWtye84F09MB2IxG3ad8j/+Ex8aoKwEEUJNqaPFeF6BoGhoJOsSYtcApfct5
eSz5p/78xT4WyXHKfSqmXD/KFHJGaWARXLXNida1zTv+69AhAaVsGkQ5hRA488N4
RGDoVg6Q4OiWvuBfKdAcRlNBSk6oxav5EY7MEZp3mSJQczIIwEkeNip93WAzksVm
WgVGl0qkFIlO8mY8XS+kBoD3wqV1am1OxQOUtbCf1xMBVUEkq64gxAb89q4BcS5h
qlKB3aUJHkDTkaKC8LLIFG8T8bygKw8TeqcpYQDyOGj0rDK5tVwMve6C08bZoIXR
wJw4q1+kdorzIHJizEE3NOY9WzBhKG0lQZ3vJYq0jEoOzBlQw0Lkh+2CSroNiDmD
GYgSE7AQuaoJ0pe8kxZEkaGbD95aasyRxaThkKvk2PYh9wTaQUNrDM3DO6zWh9ki
TshBqV/k4MmuO5WbAh/5D3vIxlaz94qZ05Rr6qEpfydMxNLF8B18ryTTAajo6Jfh
mLtGaU0q7aZ3gqvcMHi58is1c7Aqha7/luPGy/yiHuEJ9JAxHeLW0AQITBLwb/iW
nrByi17KPWEqMzOEXuG4BMTYaIe4rH9aVzAYsH9xDkzBo5RjFGTjGg/+sO1rkWb2
W3r3ql+2Il693wH+HadqV9e4TPldh77FKqlTTMGUpJQfhY/fV2uytMgGNrwhMyE5
T4cpgBm8tVd1+0j9fkcxHEgvsQktCmAPk98DOC13JigNdaUyTaJc8QyidOeg54cF
RQCoofnvedEVaNrz2WHVLEOPGLIb5TbMSYI8WBoVR3DD6Vl3dW0XZ/VO8NuRF4HY
sNDwjQT2BvLQ/wrRKFnrq79JovIya4U51bhU4oeG+B0Qj0J0nkrJv9S31NamVmlX
uXrF4ZrRst68K15Cm8ZUxQM3Z5A2eg6mCt7eoLHJBUR/IocI9pCakLp0FuTnCtVc
zkeT3mN7q2TU8X48HW1j8mcxdW6GBt34Neo9lb5z3v5DdsfRKQZUvxRMeT9PRfNX
caOfr/7+dz0GGEoQDAb89L/jYCDRAykINk2LzSWLSzlM1lIIySELXWvGv1a/Wtxx
9hZndJ1fArHLE8SHE7OfGj5xpgaF7We1MJJgx5lG9lTdfPp4BnK+9V/rgfhHZfFV
WaWDAbnV0Z2oAk41gOg2lqhx+VbLeux1HuNPQHSA/WvyzaQ0eOKt6GLgAXUeVw9t
8gv/ByojJ2OIpMaW2u4xI10zM0d9xVgu0wqSDkTi6j6i3D+xc8y0T5bssbsOZOji
ZXHTKxdn/rb0/mv8chLrqh4ypZvqwyyXN6zgoRkOWGayvCuouZUPv9pfJsDhL76P
gJi39p4+4RCuk0PT2ENzQVSOqS0IdfojrVs95LO6M/I7idycn1TWvMEIx1YbHoTe
MFTo3dTQJ92701cT/gw8c+JnPWu9Gp8J2VbIwdQnXNhJU9+k4fpfBEjX+u9SrFXr
2ieLP8MuRXTjCZyJm9qMYUeZDM6lPvpJ6xMMFSkivqmAU9hod7b8Pxo1zHC6GGAz
IcBm6Cyrb5Lv2M7gp9Z2PLohDMPLZQNmeuEumrZwW3f0FUTciunBcHbuyPxIIdTc
uhQN+kPg9yRIZvavmoZ9BJGuvfAtDOegw5/+2ndc7WNrdgpw3mwZ+oPYwK9x01c3
ylEHCz3QiMpYJ2Unv+tMUaoqHoVgo0GqY53gPHPZHpWeK8eoxqYVcWEv6sh0eNUd
gfl9RxyWZx8E8IQeAilmZDlo1AJcWqA475W3KB3RbTbpcbjhdoTj1Y+R3aKKvTrB
P59DbuB8nA88vswX+0DjUTtXyMyV6FkzEKZHYqW8Vf8emBS/OcVJItd2mCprUKKs
AZ7T5CnSPFv3CZVFrDDZAXo1tkmm8AMXlvP+bPafLMkZoCRcMUVHBY9Lu1rDUHcx
S4tr/CJHHdxlr7blZidvNV0Gc+0YqoXViIt7JCtu6Fn53Kk8MBJ2Mv1Zcjc+qdAC
ASJQrzeZfqG739s6djF2yAcelP4R9FW7iFK4przkomdEisWS1am55mnX3aHrvOZj
l30r+RIUxY7ysYWfzOz0DQQEViz6+ku6cLBI22/DgwNGTV0zSGbGZZ8AJSsYp0sb
UyiNoy6wVQCR5p00IwU+klCdhvLuDaHhHOjn3aO91LXXE8tzImlN6q/+3On0X/hL
utgFtLL3LNeOZ0g0SnbUG/AkaEdbOilgms1D1NRY25edMcCa5luF3aiE5SNGBWJ7
SOrNNlkn2/bPTDygAoYfefoc4CuoAGBcJG1sCydCxkwslMtzLbyXdvn5ZoFLVuoc
WVoqoNA1jm6VN+Ye0ffOrGET8AYqHDY2WFRqRwgLKsxNKbi9zzQlZWNi4J6wy2kH
WhUjW+QHDXjNZvo6KHiuLFUO1OSRPpdglV+kinHzPaUxH1yzYRglEkfRqXljKAsM
Si/6XHyYdFu9tS4FB3X5ZjdUDmSOcDufe320ONcoOnLmZLnV/+jfYHozYH9TjsnK
bVVad4GZmHdYWJaM/pPyo+8bcWvgKYpVCPKkvpQZ6fqG2dyqnkF7USYbqrKaTZuL
DtpiyJux30bkVG4azdFvNsM0DrvP0DnryGfENoKGLu6Zff8jb4S/6sNvLOprH7YG
Ow0oJfzNenEezsRUgU10LmO9znjvTKmvJUHqYhxZHh1lX0XPr8n8kUVN5g+4OgHy
E5a2CnOniU4N4qE5GIosVDC9y6ZY2v/PZWeqNkzf7PTcZL7aVy0T6TBqzQmeuh6q
5S3TZ+AtJGemG9LExPCBlKbdMdnntfHELguzINsCUb+bknZmjW92VFjGFcV4A3a6
g9IPBDKC/k8Zrl2LVYnG8eGa3gZY0sh5V6NYxC7telkmvKqazT/mTs9XNje8lzu6
J4jG8m5gsR1B58lajHJIbyyXlS3hKet+NxCV31AmUr/tTwFB52dfqhU32aHTdJkb
hTAXHe2SED+d2/qew5kMXoR+ikzcvEkdgPPW8gzQ9sjF9OZIk7VUAOJJtHRorAlY
wRCLzFzdK3610URUVH2cdpKyTwWPE+g9puQr2w6hKmIK8fG2rbZ9PNg954R0YHTx
b7m+STWAPT2yec76ZTv99SIAEZehkDseBz93p+llGNXV+SSrs71Et2wrlVvat//e
Gld+Ff6izrfrVbqPrJY2QgIDj8VsU1Hj2h6eEu90CFUzq7I9+Ep2Nqi+jGmOg4Al
qFd3HescLDSLjn0Rh+MmZhEcqfTmcTS9I/FahPsUenvj7DqNcu+xvKuEtDAj49vh
/3ALOWw3FcXdITJ43+g9d248GUHH16TQgww6JOXydTNBQWcgvP/PczkiI9Qkkdrs
pFhKHIh9EBkM/Vd3G8bIeaMbkWalitF0T3lwoymAVfCdJP8G2g6YlqFmutIZ3yWV
hy8xUQcrbq373j51Gi8UthpXk3X/WbFzRICI+kjmNxaiF5FHTSB+x3h/LftJoL7k
XTf7uNdQHY1kY7J7JwS9/EBYDNRpUR1WCpQcpCcrTSCDYnJv1fJVVAYwradR49Po
EAjUiWXkN87Hmxe8YJQjJzI5+2KinHCehirCo0qI61ooPg+CaWcPntUfyizjx8II
Pg5ONsKjzQTwCoY4jY3C4iDNZLuI//xRtwM8qyXA4jArMLE1QtMLr+GZBTBbmzJQ
zgbpnogQPOka3eWdKaui1VEqsi8avYz2Q7f3ANJlOZYYy6UwbtAQanYfdXFLrC9b
oM+pHr9ppBbbW0IKdOtaYa7X9jlvSv9AqSfd+O7kV9eOss2RTpQjOkLB9m3P+EIp
tA7ZuqPVpeTtSF2C/AWbfLl7P+eZJEbJCY4POSoWcckBYjRBp6jU27eSspHfE64M
xoHiHI5a2FvmcBSUMd8s2p51cH05uZ+R8YbJuSqFpjspwqdReuCUS4PHLMoDb8gx
tuiqr8HvpIMbiAy2c9gaAtOdRJ9Q83EJC3nK1PhRArtLZe4bpnmLO0ABaDBO7w8z
Fja72PPplbjq0Yb+/Q5koVW81+qjOeqINN8nkuGU+ArpzXzV7QOEjHLsSAoTh1xq
WmRxP1hrLqkej3+AUq4DLM69gwfcAgbIo53Ivx+ubGwl+MBXe07q4velLDc90PMf
x/B4fZ3t6a1ugtMGe/rfmiWmL/0enEKC3Fc36fqAytRrebBrSyBM5gh7ioky0gri
rMXBioi8wtVnx3g9ew2R8qdCmKcc3+PfmHNSZZDDf2sNfjsxzOvWdenFwgA1UjVV
QRpYwy6nlqFQMR+rV9d0j5R4IHbUUDB5HLLu7gRgyRfdhIV8ynLPBUimusWcQIPK
U5VjaqMSIfVKS6+Nrs3AcbIL6xl66eEv3+TqH7bsZGwTP2bqydB0dIZEKHAFDiah
ZMpZ9zm57ItI+Yj+LVRd1CzAS74QFVmDifC7m/YQg3wMVja3U+HcJbvvUNOu5luN
SDnD7OgI7FlN+UuzLrybD/X/4y0ot38J3RuilcSp+dS0xvxpFgrhc7TPlWVruZ2u
mUYGLbAYNv1sgcYociQnrjZ4jHhtHs6AN2WZ6I6uAiCWBg/t27+GAKm49hGlga50
U2ebGRoUooAxfzL97c41hEDl5rAqR3o3VPde6w7o8V3ZsxQd+6xU+BigO5JR9ie/
9AEkVMcq4JxBQ2Ph/Mu2NfYM7iHDCD/6XseO5LenzmTj+3GZ6r12+hk5PeFeNn7l
c9D96qf/90NrbAmoTghUtN3Z8EHrBRNy3eS//3jqoeFIpj6fREfSPwWQj9vfUuer
HqjnaAXhwW85bt1FSgkKsJgPwOv8NUG0LVuGsb4gYr+IObSqlfwXF5b3kAFkX4U0
yA/xN6siO4jh3CkAGrQzeoYWE+j++EHtwTQc1EIWKNgJnyQ5Aj+fYxO11Dau7Ubx
k56iZobqRxf2Ks2rDjWLk0AAIlD/12p9WkqeOMX4YJD9EKeIpWAmCmu+0EToLs+V
i35146eDQKrg0AMJ0lQEdYQgXIgnpSasNGlXXUw1/NlEbKoSEsg9bwujPga728tR
UBtcNeCfUQTHkbe1TSz4qwCcSIXUoGXvsBvCOvWG4hLfq+LUqp7YB4tOeqxwyEdJ
8zeb+kfVFT3tExmwUW+cKjWixTpj9bHWUHf3ABWelhAVY0ApEMcVjJjl9gFrjz/U
P2v3uDpt8kt+5yHdh4W+kcs3Bz2bxg72oNRgkXNdxjEfTcWA6TdCQuGaRJe3y5js
a2nT5kbL/L89D5IvGIlpIJrIjhOoDvsYzdtSSNBXNbirsv5jI80U8Zktv2AjO4n4
wxMzHMF2gnJoRTAYHfiDQfJRujUEyYV+n8HToZCsB5Yu1X2rmCrgqwCbJAY9/2Y1
x/0/b2yTurAjR34eLhlnj5Vxs2N5IoS7O5T91iNUn1eUjDgGvpU/PmpY9yMK31lp
a6ULP/htU0OzUHIiFSSzSNwe8F2dpgG7l1jgIPNLomYt2ZbY/3CfQn9N4BREJz8p
XwhlV+1+/jQ5zFFNgG2b+ZKd0zbNrxhky36J6T4GCnQg2yDvYcDqO5+E3F7a4SFL
NEqUYGSSgLj0CTh5QCv3GotmbADtRqofrXR4X4jUqOaP+qmuJyIzdiL1vtWQJlHk
P3CDtZc5a597xdVTolaNwQrauTskLD1fjNr7ONfJf24xbCDWx993KA2IFpT90+0Z
ZNqCkiTa+spfX5PW1lxJL8zzIGM8qP40Alir0sxhxQfc+8uTHSa/SsoNzcVcdgoJ
Hqem5gvgSX2akVaSXOH3t0YK8pfh7GYK3SqQPLHA6cXWyaAVrK3DeAjWd76h96mp
k6NpU4qpR4F5yH0LtvQwNi8XHMPSimUTxsm35mQ2vj/7pUj4VyOfKOwOre1px1ZO
15zIlrbekWfhQVH/7d7jpHPP78yvQ0e7oK4jwQz3CB4/fOjp21pRBC1b3eZbhGR+
6TgZAL06ntoxPojc/hrmvcWI16BGwRCRC9U/W+tSDkfzCbwjn5/KopY8manaMI2u
ZSnTEl2CzUyQ3zeDP54X+LNScdzs4JKtEfSu8buc9FcfRm70J8yKadoISwfXhfe6
WpQQ2PNQo502wuia8ptXsvtL46IkSN+z1AAmDxfy56l8tcexIuDAJv9uxZhh8l4s
vL0sU7nSQ+a3X3+ZF6Z4/raiUB6Dd3xZwoe0UuGfEG9uAyqI7lB0Fnr3xdExuUQa
thfzi/ylBE7SpCNUsTLRBr7jfdo1DuQBo5ZcUcXF7S20aal8r3LWTrifiU7M1thS
f4HiAfqdRUoAUDzMzzf7oj8NgMNyUFmYtYBI/r3bD4UsHVU2WO7nBzlP61OMEyWc
yYPvNcyYd65a3gTIPe9f2C9G+Bve0DRjzXrAkWwGgp9dWM9XLGPVZtBOYi0h9qyi
MR2BFh6n1pr1Cw7eU0XoZeb7/BhlqjJ0by/blTzbbd7pqRTR6VpKQuHL4k2K079L
WsT5Oy5pFaStJ11kZ2/s/3BWKmVgYbd3RUspCtZamB51m3FsOUYEc99KSWFB+avA
spi1BeVcOCiTXQI9oKpH06h3bRR8mDx28yS8wI/HCAE2CA29I1a4qBpTV3QPuddF
jDOhQ8klI+I4/55GCfaP8fo1MlD72/KKeZoCzI0InJnYk21xPoxj974KbOnN6T4X
YYrx0VAax+bTfbDeHZHbJ9NRns7pLlYRMy2ZbMeVFeAuQ2+h8018r1ZQ12e5qqA8
7XE5vs8KvbvRcaQrygCBDO5sh+RzbMMcmo15g0sLJHoT15S5IrYkZ/bcvXl5MNDx
zcl95Wcm4CkdEomFuhlNYbLcstMjml/3iXvdkAfIkCL/cG0pGlKrZvtQZBPqBjTz
ga6hpeDvLR7X16ZpW9V83nncqQsQ9yOXF55Tn2E+tStuetHxFrHdpYKwOJiupnVK
d1e3OO5NeMVoHdSe3rsWiBAe48l7BLPTztU/1vOZsj+dsU4iOhYe6EIkksfGOkXX
r8clmMMhfhKbO2aAdbchpwFM9L2neWKGO0vHRBfBgTWxXUk/IbPvGOqSeFQThJek
/QhvYw2Wi4SE/Pr0m+bSqPhf99G0GSJF8rbIw7dZJGd+/WIwqiAGmLmGbQC9XtKX
ygS6HeGUn24stEtsJtcze91eLOT+0DSgo0kIjEQgRPrucikK0gNNALNm+fr8VHFS
0MCOk9KNYhq9ewUPrOWxSvnRgoorN2KXbieEUlwB0HTF5b0GvF3R6/E2cVBca7vQ
dLctcCn+STNXk6bRRbzqZv0RIqU6hPd8Cn/CYKvtYrF+06TXXYkN2/Dvtxx1X9hI
9YeA+cU9GHAxH8/KE+2aVp5ZO5kboDzUL0XkFw7m4ocvRdASFaNC6icW1b6JMSCP
sbpLe2/6M4EZIa0A4/yuH4eFgx9ExaqjuOuZrZqajDLAZbKOA8HmVdbsT79VtK4S
6h6lfT/JV/UVWCe6ZHUd7+ImDbXUe03NT8hADvCnqmajr3wDMU96krG13gtY6sCG
heuyFMeyQSrbSy+RC5htqFBfK4p8Ou7/zYUvGhSJTNFrZT156SchFSD1ejWha1dZ
td4h8T5dHV40fyMOH4aPV5bB29WXFVB7BPXkYit7lXv9R27tm4zEXY6bcNcKW0PD
HMhOtWW3JNiw4F1kh0UBCVbIfOGCgbxQUh9NoaNYqCvZKNodH/L6hrMA4GUehHc+
4wlMY4aobBFqMeTasz7mWQVgRDI/2b4qOV0itu7KV1PB4LhceyW35AsDcEH6bBkC
t1HOG3ARXrkoR4EjDkAJff5h7fgKShEnf5ubvWL74Cm/xD/eIdt7gIpGEuIhfxgU
ErfS88MJrGqm9Fmw/n1J6QwL/eZ9KvYRzH8kOaqy5/MaFaEbxzfCMK4ghAnhU/Da
s535KpLOX1VuA3IaPDowQDi5ldSAvFijyjaxhY/oAEMOp2lnRVIgbRmrHMrB0LEn
45nAlfsilWtPWK6Ei8sRZUCNGStR3aKrjTKwIvmsliacJb5qFw8Wh5zJvmWRJmsG
lD9ri46DRpb5chO5wrQWg3BWRAx6uSKW31e/5QJZp/+X1DryUh+MJIP7c4+OeqCn
U43iwwTIqnsUAR5qfsn9B6YBG0ItgpkfogryUMozCyxUYlvsGkCjs3sOfplCA/UW
Kwdug6Lu7an7jpKgjqgP6kZLMeFBwYx3UNaCaCa3mqb+gCL7sF/N+SqxywLXCxxR
hFNCrh9EJyfzYQuJWkPyRBu0pSuk3CWULxiwTnVnSdBxREduQ47dYrHh0appnR19
lfHC33i0C6RPNDkZDo8SAFdSvaCKFY4h4rgXqUhRKjAgK0wqCdH62wdMrnpbjGAK
mdt6gZhXDrCToUwB16yYya6jvagd+nJ6prS3lcLwIu/nlY1ugBFT3klP5ByFCcIa
7B38WKdCk2Cqitzhr+xiejqJE7ts+LcQZhsa7wNEwPddFYnPR9LsrWSngLjd3X1L
tDVPumsBmgPDrwJ4Tr/nJZXlxtmtXIUAxPIdmN6M+tPNiM5GR76/Njo+IGQXBk17
0aeoe+4pSA4BBuHKTbnVhTA2NZPusqDc2LxSj3nj3D7BYIu4HE/1gfBfCLPkpTyy
MLAo2yhUeYc02TZ6A4eyTJDo7hTqE3f4ykACt2E36m562HFhLMNqs5i/0jtxmhHT
dFEH7TSx9nHrxsiC72sifpTHRh42phsXSJSPyNy1cHsADmp3814GvF8cFiL3ILO1
h5h1+XuySYF8yecT2cIqTwhIscwa2KIwVpcbq8ZsRc3pLIuuooIWWJQ+FF541gQo
92sSBktEmhts/iufoQovH39xBQDORUKn3lVBKtiVT7TRqQFQg51y9VqZU0SfqFAg
UTEZASM7D7kAL3D8/RzGSnaihKtPRse1MEmxLY/JPHFPHTaCNlwJE8ZEN/576M3l
ZCzrjjx91vwov1mTu5yHjA3VIREbS7cd1hQdexbvkqlCpHfptQeKDjskW+5N0Ldt
ZfIOqPYl1tkzmEYrAbngIAmwdu3Mgf26PG4j/+imLrAeUEOAmG1z9Riqkidnbmdt
aav4SMXMb9XTK/jxeqss4TMrto0opps/b32+ND97rYbH6rsa1to32YqGlMUd5JTF
OnKei+urI5Xgb0N4mpOabOo0EBuGjXeEvDCpjLaUQm2bwCYJ74qB/8m0+0blBpsW
JYiGUIfUVoC+4iUc2DR2rA94Fjrqb/DAfemP6KSo78E6PfprEU3T6AsmL6ii3qtg
7bHBDzPjiWUMtodP8vdAWheavNj+mo1bfdXOkJf9C3st7HrysroChN07L5LHDTJ7
KPYZdMn0EaJKWgrr5g3E5A7Q69LKyb1nQ14kvgdhdPZTAxDI3NOk54MiVtw58qLT
tdNYM5bMrzOauixmpW0B0Bs3T+ZPa40IR0r2BrxcVPZlttacd/R+gkbqQ9a0GLbj
qzzVRtA9DOhXpE/h7ivo/mZhEEobDbFAw0S9x+2XepGPPS57gj8NrY8oFQM+0m3E
x0F3XQmqAG9FuPdEky1grVhpFvAWzvxknqU7nll0lvTWEKTJGIsT5ck0g5LQq0m7
i7yZNJkOGCl1oXx/hH5X6AoFtPWBDMc9hRS/izRA5gIz7mn6+mlG+xHwnX9BqHIL
RMc1mrfID2yYjcqFbodh0rMicWasEoHdWK09eozaUY5fhnqEg+Pg+fKmgT3vkp6o
1oIdVfdYq1fqk14nSZWlaOPxt1d6J6DpZQxZzNSAvdZT7P9/7xgAuo56jFAZtQLl
I1FMldrjRR7UylgaGGtVkp29K8QO4k83W5LDepamV/+uyZSuCNgbBEn4zYU4SV8L
SmB3Dnfjp1RJNBsmlRe6Bi2nF8DTg09g3sMKqjdcDq47r8Re90dO/FmhybZEpDgS
SZ23ElBnN1A03zdyEYYWSBa1OdDU+/vj8bL7yUdCG9XKpRbYNozhiAj+EqsR9fJ+
R2cU3cNiG0pHbXO3WOcz5UrAuEXt8dXnNphHAqYGz/SjCUPezCKON+HPlrJ4Nts5
FQGnbSiHkiB3d72n9DQhgcd1gw868iIAZxldYpBRAGYMuPuzPEgooMKGPhkj+b2D
0bMmR6FdvzAK6vB7F3N5ao1TVH1Q8pLyT5SsVpMHTaD4Dli+Saja7iqMY0iNNY/k
ePKynKwEw9FqWYl66rJhYtQjIx7Y6GxEn4tvoDccu9JfJ5WSPNUR7D7PD5vgl6iZ
/qMsGfJRTHx4IOi3ixnLmAs3ZT7JuZtUr2+JXMCO3UJOWoT6hteIM0dosKUHV35r
b9UE1xET6i7y1+guEpqVLqarkZb5lxCaUFBr1AaXjgRNW4wvL7l64raxQ2uMI+RX
ohm5D5et02bL4qSu2B9KzQwO31VXmp+YsHcS7Q/hMwsaPKXZt7MP8lem12mjYJk8
RBAr0apNsG8KqwNe+ZDcdIYXAMIQZh1JGoTGtW2Ff0N+/Znnd+YeEDLHlhrcncR8
2FI6VhZtWpKlx1AEh5ZHjduOs8bIam2B26vaB0QMYnBRl+chdWz6EhJ627x0M1IB
rzMa89NbVwnbhVF6XJznfpYEMTWx5eKgwZSaYgRo7C31OW/wLx+953Nl5cgC9l0P
bA2oBcqqPOmB0sG8W1M4SJ+juhxVPTPo0dioQF5fysmsi58fOTRCqCfjFqqMEte9
62LKqEHw+5FQgRGTM6QoOB9haf4/5lACD6AaBBbNKNqAuGPjl6xHpCbmTFpI0tLC
Tv4WRlU1s1Q5xGwnsAmRPslKI2XyH+0MRooKgly3T8GBKjy7T8K5/omfN4dyV8+d
GRg8Q5fkJC9TLDb7IVssuikR1HQWwiVEa+S0IgatSPNIDq7F/UllJt6Vt72TcuhS
vhhlV/l3DfXysWO7yIDDgdKgzrQp4uxc/Ko1Lk4AfHTcfx08PKG3xypCZ9VsBBHe
yMZTDC9BNPLU049ly8mE1ktS8ofDS4P8waawbSV07aE6SAWxwK6X1NxeFN3xQVGc
EGm7ryMZiEhXyjL8Txcg9pG7GTYMoRYF+8T2nHtPQuzLO//qbFtCi3oBbBQ3p3M1
xOsi8apqrMEs7IVktzccxvKbpt+1Gl8/RYtSP+Px2oWSpeMOzqdq0Ys3an1kagvw
8fCiGkQC8fMtfX1ArtSu8sZpkIZGrqTia2HNlZjIZ2IRkIw8S/5q3IIBaPzKG2c4
ZyrUoZ+IpP3WcphunaxDSN+A//V++ajdX3ZkggM9/hUn4y78eYpW/YELDRTQa+y5
9XGkyss8W52zKf4M09Q7bikNfZK0Dtl5zICZQASBGwJtJpJDI1l2Kf1Nf4ni3Y2Z
8uYfRd7LLG1eJ5IRrymnNBPn0vvr32q5vYMaQlsU/o0OSy+mFaU6ftLcrowkNb5B
sfIjIS4d+1Crq6I9jl2aibbqpMdrROveTzKpyNrvjNjHoHOXJG5tN2jQ2zvm6e+7
8fIayW7JPSPd6Y7vLgz8p10BoUsYd7QUzrdN1LlVt9n5JlYnZmB7Mj2ZBE3cVafh
uD7AKs+eTJCtQZLWyQPN8B3gw45HqfJHCxGWKwtNxX8UplKx8LjCX6OkRqblHe3c
ASt4a7VBP+v3hjdttt3XWH0nM7zW63j6hfg9K/aSvtrl2hMUm8M3XUEjluoXi1NZ
93GUdJm37Zpmhpxk/YgM3TH7URkKPJT82t7YTNW9Gcuiu8qW4G6hI/QHizdn62e7
QKaeJDFRDY5uID+vMLL/FR2R8BhHO1xmuTmwXNwWtjL0oHjicVyw0eYM2G6ygz8T
434dUhPVSE70aK0qhUgBQFIQKyQOZOMaGq9qkcYOceLqOszEXOsK/RHC8m7n1QcI
eFxu6OsCyoFrwZUHhu0HMUPElYI0TaDYMZujYzrW3DLtNncooGRnrjonBFfVgw4S
W8PQUViY0TsCwUCg8b6ksiHVv6hSP1xvMwJ1t7Crn21uQC84GD63cL2+ZOE5ri2S
TSazse2TNQOILjZayP74XvyFTXUWEEY00TrJIt5u00F8Q0pEQXGylC7RtLn7HsRO
iiQ5EI7CT6/kCK6iqreldldMI6xFtLDIpbjr2mMLvLuK9ujgRDbIGdwBEWMzyjsA
EE+7XpjhYnmbqnRO8C18wvn/8ww+FWn2ko7fu8ze0mKxfI/g9hTDYN9AV/J/kbDj
l8cH51WdaFKSBbZw7Rv1X8JZ69j+SQQFzjPsuGFlj4FSimToSof94MpbRNwTv6/X
2VTF/3IcxFDI+rmNkZKanm7lG29hQSYbIWOEXVAnDVHg+AlcuMCwFaOcUwPxPtKO
LIg4aFc2DN41MCuPolkF6zI5SW41Y8j16kiAj6wWQg3kewr48++T02h1cFIzB3rw
FFyQpqXETnnHB2FNuOiU5JTAks0rxY9gRcV9hnTlTWJBQU4p2r614LcV6w1dcR1I
/wonDV+HuNaYSqahYWEbZi4PznhVN6U6krriB0m8U6yzbTJ78bf7HJESOCGKNQuu
1s3nzah5sEZb9fKH/LJZUDfn4z48suUhNWlA2pSBQcnKfQkDEx54nPjyI5LTnysy
EW2idUiBTnfAfAe9ZQOhddAAxmfg2FFMD+/zB/o3+kEDRRzmGs2uVi2aWqeymZmJ
I48pxykJ+uDfs4RGeaP+E4RhQwivpX03v5pQXd/Ougn4t+3oyKkpCooaLd5UdpKf
NVfWUSenjOwkozwp7b0BK+isqAZ9z+m2nL8Pn30Ta4ASRZDb04tnlvEbdAN+mTci
IRXFea8E7qQM7uyycHALN/5M3k8Obvpc9vGQ+BG3buCPRgXHvKPyNFhGPkbNzANw
u1Pu5UuIyFNlrbdePPklCH7wh+CXPeFDBbqfxGf7PqWSILqOWswnbZuwvyuBsf3v
ArJH6YdezN01URd/LXzU+Eh5vFFDtw3S38Ed+a2ceJJ/yXN2ExXk6688Zzmx1lkf
FyLKDe2l0R/ZLl9NnC62nDu4woIbGI09LzVwedtho21b9li7G3ZzG1DsGMyYJYn5
hKDemTtb7OkXcCerQ4vSttbVIXtx/Jo0TCTwY9HMhD/DbRPwuftgadQ0E+gyCb2w
fwLK3sFVQMZ7d8ZsJ/hAXEOLA/6Gz9hxgwagGaTFrZqmnU4HzPaXjlyucusObAJL
KuHLFi8Knq6AvSmrlOoPRrNPd/j83eLuYW9NMSZMsMAA534pkQ+xsbIwGsTm3ClF
KbuppOfkWiBib832yCxQqXUSNnKssNjYxK2bOFljqV1fBS4Y+pvxBUEKPvN/Jcrt
g3+9Idf20fFolVchzCEX56UWS2eMYKQTnzo9e//zYTnRvvIphuzi+vrBWCop6jWM
f4xbnW2KR0R3aGNseknFEJHCCzrylZ3Spc5ZcUFF1E6kzRYrCzHm6kEpv/4jF6Rc
LIBF6bArJxdIqMfVKnHpiMSZHO57uHELnE0UaPpUY8776bIp+emKIvg6WeYWeG/E
ejNrSYLyt376tk+Mca+T4aC0Zh2MEMds0Rqi4nuLNUJvfFdifplJeBN3XT/qhR4S
7K4XPJdtKENeTBKuJo066RukJWS9zQkDLP67ZLYP2WxndLk715+2Hg8t4gbV1EP3
oR1G+WTijlYZQ76n959JFQ7L9jh/GJdLFwwRMQfQhKPqFzd9uGpLg2/bIvcoADeC
xPzNtH9ibTX+2MARmiiMWlITwdk/FFkEyjvNqRlWKRHRWd1DToJosXso1Mi9+Wcg
/lzy1euMU1D/rTRfi4dSbyZt229w/pbAN+pgZ7YQPZwVumfmqa7pM8v6z74O0fpI
T/ZTjTVo3EIpBtR7I2xArCvYy/zD1azFdCflU6sKruAE5aUoy8pxS3cQaXYyBe6f
8ODaK11Xa0evQdwzoMgn4gAnswiNYmxkF9CT1nfid1b6xMJPABxI3qVZyOkF5Wpx
oLymDMorHTvGIyfCLnWYua+kS7GMs1NemEJIZTYhRyBuzGwM1h9PeqimiDYP9EXd
29Y6GDNroiYG6N5rAOC0yEh28vjcp/rKAxjU8ey0/JK6dQb3XzSn3V9/6THzBzVb
tdmzVHKR4/0r1n2Qlq4ao0w3B2Wqm3QY9lqDmxkigb4MHTdhOpQw265o4suOwvVW
Jberi49rD2hPbOBCsit4V8FAPi79rn94tWM+WZk9g5LsfCqLgIFkFvwFUABDS4Qp
BjcNH93pOc5+eMGTWTxgzT8NZWW+0sAJfaCZj5+BAb3UZHRHpWsjBHMzL11+aOhQ
Pi6/Lra6UhOvtpZBxBd7qFq3KvIrUpJJWQqTVQ1JxpidwEQxV6DPZNYCwjSnKg0o
9A2u/VWaKsgRHQG/ilq46WLBjsv8geRNu2WMTLMVEx2MxfpjAsFF7Nto9eZrOqgz
fTGpguY2NGleQog4ZEinf3gX6F7jn8NWMskAKI/7b6NmgDXLZ/iITYkP6YNlIGJ/
iTjkWP8x8ufpGJS5q9k0JmWNjVOXmxpP2Lj2drla6XFy4NCvG1gx4v5t9Gdnvoyu
blBs2fXO9lv+SNW779FIJCWZOd6qvOX2c0ojEpgxocZbpmyCa4pmb2jwILT1W4iX
3/RMvXCsF2weaXz8r54if68xZ+aMiOefN22vmN3wLZuM3Iha3fDqpaT0xqCS1Cj7
8E7QN2/KxW/+X93+4auhMlapSzJ0oTKvte4si4F5zq9Jd2Q4X8qYQvICXfGxtl82
A9qnJfoiJnFIsobPlxXYVET0RfbIpkENdmAzBzOeeeWwhuFDCfJw71vReJxvwEFc
KXtsV425tWWzrVz/bwRjtx0LPVqU11VEdkfzz5CP6zwyglVQ6wjjl7S5InwZdmE0
PrzE7tk3Jft94f0oNPniwngFaK5NZRB2t0AxXLwwN9VqRE2dQiFEhiBVWl2JI6W2
oqU7N7i6lQfsUYkp+EhRG1n4mYKKAW0xysORI2jvTBCXZU9TgQZYfF7qd/IFKYex
GI82c7wHhK1E7bVlHZijwibLI/yHyDIdMDotO9VlQ2/tSBeWh4F7UlpX+yv3vC62
8Mh3OlaVmjO+oDYKQEHuv8P9a6mhTp08rmJz/mFtdMgZSCaxJHYQvDMzjahE5gRl
I9OhaAoOquiSZpr+TjvX6Ivo441QkXllFTQWYnRqZutrwCUom5CJ6KHnOde7OL1k
F7cd0caXJAYAWD1FIuOpC7Egbq8CjmUb9OebaljfEXTvYVSRaZfxprDUriCN3iam
tMC0mFZwZJbG7WuS6rzaCbSpfjHtapGhW49PJHSnrjfOhikSE7TIhRB+fD9tddIx
Ur1vNHaezhKcs0p3I+TZgsA/2lqpq9yMpR2WmM+wsqtba5zF2ztvWEaeNnbqImeo
wqDu18sXA2gl8HMMfNUzGeUIS59ThrYtAfFhXNoxzh+F9KGUZ3X1A5uKWoW1mKTs
q77BHDinkmtwR0xGf7MiR2fiD0YSVganht/8QomrPCBmFSj/7R4fMXV79FowSvyE
kTIwkZg8+k7VEaKZWu4HaX165kS708Yae2UujQl8DMNyvVjtA/FwNi/YF3vHLVX7
jVbUt3apVRCCg243g9f/hwTHJCqZdZboFqjVGcrniXsHU7XjS68hW1G9uTvylC/4
JWUjMxNF1/NN5SUhjY/S3RzZ0pQVTKqzqPxU3vxHIrR48DA7pwts+GLoBZpzdcKb
/fm7DCD+40W29dCjvxWLLNiyfMCmgRL6FQQzHmMe6B5XyHwi/2IApagsnC5wd3Xt
RIxmz9VoCuBOHU+7ykUVrf/O+d0eOLGvhlwhHADsoU/6MFxFlK9jCyn9cpiNy5zG
cpv+XhEwhwZ9dBf18Ll8pWkJMS0a+mbuJfAUKhRnkpLx9iUb5Rf06yJGneEVOFQx
aUYHLaJj3wv3Epz9eZUhEaIzR5/PGex81OopZM9Ea5lx/GxujaUG2YbNKAlKW7QL
1NzaDMyvHhblxImeRj3oZYI3s+VWJcTJSdDvry+Ge10KPxS6lg+5kNK8GlyNfu12
BzRzoIcyzUwXx1LcbFzcgsz/Df2rnEZc5aW7d6dfrGuirc5k3QEAFdGVzgBDQF0J
J6THI9VkOk0UiRk6XXegnr6n0JDNVVnh4Xpw29iANIlttaisU8lebdpF0+0heuDO
rJLivTkw1ZQOEzfTZEWerJF7QaADWl+3Wy/+vSHEFChx2vK4hdd14krUU1s8V7YE
XWXCtFfMImCZ9WYUORxE6okqskbB8qZxX+ha4p71krQZuBEvKX5zFeBbXTv5rMW+
QrtGVR/KoSWvI8BPT6FFdBkzTeEs9XoEsHmAJ1xGqqXACI9nqheHTpC1MEJGQLXK
/6YtFryvIUaSOW9C32cFvvjWkpjz4PVnHrPJYP3k0GVhHhmPmp1Xto0tnaBravvr
Ss+fKtkrBtSsnifyPoaqVidTqBU6C0IJndVrw4YPJjOQ9g5sNO/FvEbxW2v+XuVh
wYk8YsuEpcnz4CBfzTrvpW1MPRVqVDcGWtBEVkIitD2jAHhz4ULTTiG9nkWH6BKC
xPDxTdF6c1Uf46nqbxnjE4D9q7qdKyPVTHhJ5fkxBImHyjLa6QtSqD+8O/HPObcM
DQuAc6uPx1cVMwLUCs8u9T96oWsT/ZcmILdmvy4uP0fXVTwlNDTsgmocJlpv9I9c
GSRQFY/F5aYtSnwpOVwaNdusOaA8TCBK/7gSHMxjoKk7BOMZvpefI3XjQgyIIysZ
zDSe3IJKNBiQZjwbT+ypDPwSVfDTszEfWt7/TSQCFigJKFDyvzI3nbRGYeLeU/BM
EZtOYINBeJutwkhFECIiKm1TD+a+qYej4NEkAu0ncWUXySkxrSluVVQRNVyZAioV
SaoBvDH2lFdVe5xQYYDfVvmkTcOYGjUlQ8f05HcNexpVtyB6NPXEmzEo+4yEYIkA
ge6r8V5RITdKMERHl6a6RVdQnmHck/+wN9iMMkOufsEvHmZ74z0A+ndP348GJMh7
NQOi8XEmKDdl2sE7s0lWVkz03c5/xuw1Z+tkoBD2oXu2I5WMQiTGV80IeUVD6ZEa
mRW8rsZsf2pcYBdvRfMX3nLrVEH0mPEf3zUrjwKx7vRezMQjxReIdn3sZzag+IeR
TggfJxzw3nC9BRbwOmjjaXGVBkdB1PAqxiNDqOBRJaSwWe0Rgiqrz2Q9j7gKfKUj
0jsqtNNOdod/kUr8FUBzuByf0jBtEyHnxuUIrDWsQPwwgdFh8PscktPgguNNTwiw
EPwUdcY5yj+lW8Jmt+L0bFsEMGapGAqqpsFW5imRFtaBGYquAEQNUN+3sy0VeLbY
nIwDTG9uJPywPPW+OL3B49/bB4zgAmdCgGawhyqQLwwNJDAwOwXB2YxjhH9ZHz1m
3vb5tmnDrP8XLi74L2X32ATjGfIMrGHN31gzZHYWiZY9nINJa5d4EIprzuWXLEk3
66Njm2CpowAxcX8YwCkSd/LpiDKBLsKrqCjwsMQAb058iKy+VP76UVtWpwyc1+2c
hq6EsG/4SE6z5tQeJdk4+oG2tB/piL+1WAxDXV6i1nCtHDFX6sururZ4g3mXZONA
WQ41CABz8lE2kr+Zfhx4gcsevw4oz6PlIfWaTdd4swOEgCmZPHdXa+0bHr3069AO
8x8nwnGmY8O1Pe3mCA0Rm3o3Xvd33nwXiEsSLUrOcYv3Ayriav0KMIRDuaX3r+RY
/yTfzYAMIqMcBTUXEj1D2OZ1rzFzjSUjg4rA06qVlLZKJvT1OqJfraIc56WEszse
oha65fFwyyF1N/jtMET1CcuywiwEh+q3zQB7+jbVkeERtxKIfaP45x0bUOfo5hXe
IPF02tXWBQ3ESUCMXDvEaCdKsdvPB4I4TXcZ/00b315gXzwnWbNmDTAVgvGP/siM
iNr4Mj34devEtoIGWX8zvn+iTnnY3z+NRg6UX7qlcdruAzV7UOZHpH7puWyoFAlZ
bB4Spg1dDWl7U1qZOFzQ8UZqJbqh1VsVbS/JgMdOUzAkCwXCkU20m2okLIUqx92F
UbAJx0WeJ16SpnmJAYGA3VozOjpPCh9jhFvoSrSuRschUBdBYJ3szWQJcsUT3U4l
SVWj9dPqDP6zD4/TCCWvwi0BhesOboRSI2DjFOKeKFLvn2/1ErOM+DssLKE1pV5N
Sb0KIWXaG3WeihffyXv0a/XfbxhMnYYi5Vg2xjMuytAGRxlG8TPB+xRz/SjDxZ/6
UTd7/Q6gp95675koEw/85WGT47uCzI97ETmderM/aSkDJ794RUYD28xTdvqfvhHq
qIAWp6cfu8DKYsGcUs9hmylu7ARFnHhezDeF/vPp0ciYQKkhL/XypZfz2mzyI75p
rkaGyBtYESvN9mCyGixa+l+llXmos8Wl/PB+AEC0Wy5y6Ptp8ObXanF5Mdp4X4er
/nsZXlgFlglAFXcV5ZvTVuk7IWbCU9YUKSRjHpKvsBIRY+g0gFkpCKM163c80qVI
Pbgwm2p1DTVi3xJT0Y7HgJ2GaVmsCV+VOO9/JjgDMBQkJh5biUiMwOwYVfE2rYI8
2F9DuG9XW2JIuxegVP2svkhC5jpkEURQ+6MfEXpTjVOKE8ZxVUsA+RvGJsxCclV2
nvEsTYNfpD92aLzkuHfVT+CJc7xiytEpkIEWdWKGdgWe1OGWxiD+8OjT0uroPosM
r5hGwREd5iv5s5BIqSBmcP+hBeAQzVNW25Z6+vcKBJYonT8uyWGL4Ihl/sHbjwNO
4kbDyXuGZmWKolCIpCa9uADkyEQYg4yJFRl9GCQJv07EMaizRIScDMCSQkT/AAEk
XkkiH4Cm3jV5i9S6rpP00gJRwaGQ+DWAPkqfqd1LJCVLEQ73n5fgj6qO4l4Uw9yU
X90tU4cAfJ9GjjjWi9OwiAqh29BcfiMXkNZoXXHFd3KHw0jLFyFTvFTHwct7hRuX
3YUu3m0v//ndqDFC0xE+W6Ojw1YszCZ0gXW4Moakg5GKAgtxl9YHE4IcP+EZocf9
RI2JtviWyIPf9jIki2q4CBzZXAV85rvs4R+b/JYc67rWneNDriGGOD8y/+MXngRL
n5t9/VM0mn1uhUlzWgj+EiIet/yEYihzp1yG4HrRfWX+OnxKPv+DHIcTWwmo8Srn
wq6dDdAebA/cSJ0puPsFYgfyBXnVxKLq+MUfZtmmWJYq9LTQ1C3xyQMeMIOnAKXm
ZBq8OlUbECOI5GDiiW/UYuL9ggImwgxVec8u4iSBsGrM6eMyD+0NRGhiUHHasKzA
UTJyOA179EpmJxw+BanIEchEp0VxrwNISoopZZLRP/o8UZK9ubBBIac/6wHuKbPD
ed2crLX1tWwocxphWov80JqGRrktHa8hC3X3wlX5HDEVdfBfiASySopPqv4EWRam
tC1jUvAMsygFPCVy8GfJTgyoYV+c7XQgpWEmkJKnpjy734UY+W5zB52zNUG/ljUC
o8KklF7lFrzrsNqcgh9vFp0DOY4ACxMGqK/1s+Af9sp0oIrPOOaHPVxv0VANYVrw
bcVICp0XHy6HKiWB73Ctevdfrv5wmn4s5JbLu4iYu7O8agGru3yfDvZ1668OF/0Z
YUEfeUJiiO5MBDtjp8F36rnyu9D6xt1tNiJo7xBfyYzyXsgD5lCKx/I5Qr+Z7Z3r
thFF4VsKq4q2vx7YTSvabHhcR3Aw9qnUvzNiENUqqVnriNAqEAEgrmOa+uG7GWnv
48KSD6W2WB6UrKey0mgOpH50kIcwPB1porij36c1Gdgu+QWOIne7uvHBDbkD1Q7G
VdHHjV5nzWnl2Ip1GC8fLr+QBEwEey4z7/2Kc7PvusxZiO2qvxRECBN6HcFReFLX
wwX0pP0aqIuNFOapyij5JvP2tLZm/3EBV5ToR7WGAX6e/hIWJQUKianUpyoy2kab
Rmxn6bI9Kkx8d6SWkKM/HrW2EtqtygKjdT/ESqI1s8Qydj9NdY3/zNNLwwfKlPMT
iORyA1pJpQuAI0kYoCfr6kSnn++oum6fCIcoDKGexhAtWFoLU+qPCt/jkAG1VI5C
v+9BAa7RcIOH6GYrHlv8tpB7rfzGZ8n1/A7itfeq/VRrsqETvnkL3+bQWOWwRG4o
rQmQY6j1fiFp1zp7SXYVNUdA17pANnd0TfqpxU5CMVCkii+LQ56NRw9r19bSMiFg
k1wItNyDJ+slFTecNQq1KLVXT6tV6ocOMQINMMPykYjmFQElFDj9CoX2Uq9uw9XI
fJaX89WI3f/oSn7sDAIIae5Nu526g1eHsa2jJ25UXkYogUb2Yi6YGn9WfenjPHqy
EsAmD/O6tlKB2NbeFN/ArtC9VWOHgLWckCnCO2LNWoKBMzMXxnsOebgbAsrDKNud
bbLVQkKm3ppvbB3gtfrUwrtBsIuvXObWyaX/JnpwxGdJjlXpz0wFTeBCylV1RucR
iQED6F4YJayDO3KmyxePusb9izDF2WU/ZZg2hkjk5AXHn06oNSRA08P0u5L45al9
8zXFECJ2v4RGvmVSHwd/zdBOfPYBNLnwccN4dQVoCX+P4TpjrEle/3XPtN2XqPkK
63478JKf97a1r7cip/mgsZtVG9ablnrj8JS6YFITpYXqA62zQEfwtFTMKkN3jVG0
U1WBAsQQXsod37W0vD9gc0GNjjJeFF1gEw2O+2BSgp5UVeXQNg7lxBN0I56p/ONB
prQ61JFsfrzTH+if/V9MkDtwEN0Jb/Eb6ufz7NbzUZ4uOZv5UyzVAXg0GcWCj/9o
VK7bkylEog2MGpnhgHyUSaKKZRoq6em/B3Ut+3tgKsPALupWimydB8+pHDT2r+Vt
IDXiH8suCeGgtMFwjGfpLbtdbJ8koV5rapaIYfGHMJFQVmV6hg8jk0Pp7njCsSLE
csqwrbQ62NuzEVtQN9mE/yj21F5HPx11fLJCvvu5kx/YMV3RVrWoZEqt7sQSAZzJ
JftWzbHmlzH6S8vAwypRMXdDnKK4y2cZdh1bhNGAVhm1gZ5LvYmUQmdyAXb6/gWZ
/sSMohiJJZlESv5p6VzDTBkl2YlIOWW0l2WnqvpRkB3eJldlCfw35JoU7O0aCcAH
XCZxoSJifUz0lx+5AZRBxCytTqUAyqQaOVMaaDTwGrEpMTQ2O5FxTp9vx7ZKxyVu
Gg5+GCiwwJ1uYFhMeysRJIa1/r1ADHMu2i+XMJ109/Y8hMahb8iHtZyEiy7u4ovz
NzVbjdwpwh3yesL+cankOcMjQRCJvIX/sI/J0/mZwcxNg9yMnnyHrn59Keivuo4i
WMbiiEweki73h8ddCtmBoqQDnZkpoE8rMrUe7VCp0OSV+GSVpDGkKL44oV9MuFE8
psxvK3gB/O/f2xd+Q5xwFbqyNNVTV+LyDHeld1gXR5z8efqZRVMGUhBLv9c4U0rH
JXgmEKUwlXjNZIteLitVka0kI0FAtKLG1aEkWf3l3x/CqV5smqw3FQaw/brOqO+D
EbD9fa7C5PwoJGbNGHLAUU/ekjE/Hl8rSIjMOyb5ot3heDTpebnwt5ULDlF76aq2
JV306ZU7lxRrH0VEF67ZO0zJUpin/POWz4RcNw36OflFGYnQLEnwe0tlpFwt6Jxe
/kxN99ck1H6ANr0dEl7rJ8sTQSybBvSHyao71BJLRE2CwAZQmhSII0qPoBQZkBSg
qWMRhOknGZTVoGzW9K86CPLiaf8DL4Ut9r0uktAAU09fqqkX0r7lruPqeeQPRJ62
gvgrFPHX1qP0xbxqooPyZ2DtGPHV3NfkO4zj/DTTENwLCBMcK+2wlG9dAhf8qsPt
Wvd6G8Svgcrz58RakRc1Tk5NEYsJ3NmYhMqnoaZZDPrmmuU39Cmg3FtIPt3GwI/w
D/NNRWaA7iKN8X6OStqpa4etUK1cMhT4ob39CV9dBo+YrxnR+g+kIBsT+KQpKwNM
yLtlL/F8R3F/5ia17Jfk4aOYOXnKpIwSGtYq/99fPhhX3WxZuOpAKpi2XNk9W6Vu
5oMJAW2rJLbshHslrsKE8488YyowBrkkiuNRmrNksT7s7FXoi8CSheKBb6U+A0wh
CkFYur7tynPvD6Mk9frITb85gEla1//qNyKrefgLyo9r443n4MK54QamJ3dszeYG
AWPdN0/1ouVqzuvqSiRtcXtVzxRuIeDOztulrfqa/XgJFlxjnkpmQvWAmXTfmf9j
QVUE3LV5ar6UsbpTieb58QD77gg8O077o8DQGCUQrtSnBARJ7JPhSofKIi1R13cA
vnIk3d5LfAVU5q8Kg9bSmX4e5alers5aAkbY4Bcze4Xh/kTpP8ifyI82Gr9tzfzr
iNIn8w2oPGr0Snh0Bcvbd4Jk0PepP/EmGV+L1Msctx0BEZIxkPdVLJUZwrBeQPHK
IqN7EVAdj9UeKy+noR4jfEaqbGQKLpkdIL41/AEKJxOdW9V7G03FnocXzwQGP0Ww
MLElvDHhkSyuZUaHCBfH0YcFLljoOT24SFqSPtOZSOzkQWSqh6LzIZzXDFxT39yJ
UtHopYDBDLJwvbSx9aRwVpMqIpqHWu9bh9p4pzFc8wZcmfekbgGj+hRiImpEJh9s
WNiuWD/CkdrIzzh7Lcr/xOQPiqr3bMA+0DrbBHBy66kz4qmW96MkOdw2f6oDbghS
RIWbK49Ky1QTMnHG7dFMYbHqgLdujYVaZZmETw1LT45s4KEHv4AaBN7bXHhje5Q5
6CtDch8jf9bjkfUNy/+ZVOeaxAG2Gs4HZ5SViANKkrb9qQGulJlpAH4kQ4vk90ka
nhPHcMO3vjUfgpSjBIXcnzjR4XRlXzwxEERpOnsHao1p7vMjhpjEq+56dKSxDQhM
LDyZO5sePaeV5GF/sO+GUcyXKy8y41Nw4XJgBXyQsDvZwJO9mbsEsunwJCvxlawR
vinCu3qgtKND+9wG4lfiXlTs43UKRupSVW1GB700anat84Pn2BGEVSbNYG7ONvQA
nwCUmQq/IRS2uOHohaDWFNn0hLo52idUQOMPfgdabUy2zXimYeFbmcQObFLrs88w
Y2qY86jGtqdRmFz5FTcx9DvjUDRFETuRwjEG0VXpqdje4YXMsGr2v1FwngVXXNGf
PPCrNlxKNA5AoHM57gNR9fAO9HS+1BbhZThUBQ+Owbo8I9zMhpRwJKR+XlNZPg2g
97qmT7UwmEVwL7t0Ti/XvAy8PtMdL60fRZNtXolmO3NxUifaFGoWbVPWfh8BCH3O
N4zc6/LUOMs02WpPC6LaMHvAC97vTNzjl2BeVvQhcErfGyL6x8PMaHKgx7HFFHW4
7vjrCARCy78bmOb1JXiWrgwD+HYEUMXQn0F3lq7v6MA2uBOR4HvRYY3bqQ+y59JM
uAWzhANzpVfshnkoWqbeGJriqX/+FmTTeuxNgsQDN3x6O4HkVVzRsPs02Ccb+5Fh
XkeLqHbyLXNBVfGsHzYpD1ARAnnUdkagEbI5+OAXVEoGSZMClTCT/YDAjz06LZOO
qbTIGGYhu7yIYv5/fhQOWK42sIq3bKaKdFjhsCz4GrggJSvyTRNOXEAdIQEmWtu9
xFRvxZrrNKiNKVS5ipwjlSBbhotG6KsQxHF+Bf1eabFC4M/YM2a143Dlws+nQfI9
5wpq0yqEB+Y7q8lDs3U/QaJDmDRwdURqGFrnW5TkIZGWBV7P7mCUqJmbVaECfuci
g0z0nh7V5uXrzaAyDqqaRweLqwzg2Y6tneKJxB57hDYoO7I4J2uI86GSOxdsBq7L
GPvBEGV1ID6Wd8DJ3kWLfbZc0D5JVX7YmbGW3/6GkvLiogzd/w0Tp67w9GJ8So3q
IjOXyxsjjGJsXK9ftRcCYq43n0ecX2fIvU2x/XvF7wsdH8awRidVIJwgG9iD7+bF
N/nycIzAIVXksrH6qdKEPOlcS8MkxfoL6CPOppMoWegvh+0SYZ/skKm+wG9EI/9I
eKZYzLjwx5Deh3nicnm3RWkp9YEj0DmKN4pWM6FOEx8j8zDF32s8Ja9z+MeO6zZu
7ehTTixqrxv5XWchevITEqbJf8Z+PwE4dBqBQB1fXNpeYScSawhtbdLr5+2gVxF1
Vx3q3A1ALn7donFCOLXExjeyOK4ezS72ueWy7i9nlkbJrl2/txibZUWasrP1oWB/
zdA/2elbyF9VUtfci8n+1FP+ybm6bQDZq7gVhnT8/fDiMJVUbMBTq8AcRlGltYIE
VSdFY/tEB+h4pGESFQOSEDPp0lu90GSuNbgsvLNMZzk0MBbqd3DyU/QPmYgr8z/4
2K4uXcW/jCMuZhn54Nfyad4yQzGwdzGInTwE84AQqY/xBiLjpBK+9YCuFSnSiJeh
U/ko2Xj10tBx99w/kqCwhXFCXBjQOEQllZU4ReciNpO44r2frCIb2sCaUCul4XmD
MI2+gdrF2Xmr8rZJe1VM+X9i1bp2lOj2h/YPMHghsptZg2eRcKu/iwBpgmbNo/2r
3CTy9JNhGlvbsZxvkz3y+CcR4aKOUHmWLEWVU7Q2RqCbLnOia2COTzozxYXylwxQ
SHJYjCoDTlL0Jx9ElARvdqai27T43mvLrRMIFUJelU3DGTStWl0eq+3sSdBehb7K
wrJLsHw4rjAtghDKTK/Tt6dkgFYP9Eartr4lh8r7NzMxzxF+svFLObVU3ALEE/J6
2cz4fLxv5cvB4myLImKX5d/v5ShGB0JLgbSyclCbrDOeKOzatKzmlfv4Us6fJyfE
PJ1Bl9Ye2VOq04ob1CmQ+7OsPpNYKMPTkWGEqleL6nCvekyIPo6nOHUoxuIAmzy+
iqGSDipPJG+g+ge6E162KaztM4UrB8IxiYAYmSmm+GB37xet6TFDo21Dux6OU45o
JZnv1lzBPoZ1ftBdulKHq5p5RRLjxJrmGfvOAjTSL1g0+l8LjoxNAbXrqp36VLcg
UJ9rqVo0kwUJEd6SUf+yzJVX93lGPXESgGJXLOQHZYQUg0BJo6pPglKiRT/dzWAy
ed/PzKYGo9EjGs834i5wb2YwauCbuDWyQq4ZSvSAXVNzwKu5JNEDOfsjbXc0t7/r
9HNBrMaP0GaIlwNFJusWwtCLQfmzq2MTfM7l1q5pCKuZJiFUAno/8oLzLif1UugA
C9/4AtQYRPR1nifdsfdbpTu1WDI2orkQamSUKqRs6my0X0WtKdyKtZx24rF13xlw
+/VUPfBFVzHUBnF9vw7VCppbDOEgIXGLVNkbur2+yDMAb6RFLb+lDAztMn/kSUPZ
Q8zVPtvl0XI+kqhzDJRz0+dYvFd23y2+wZTm/dDJ6rFaqv24bTgsrrc8UVA+2/be
98Kl00bxySlZ3KwqIOd8qsupmjw2YbBsZaCPB+owuq5eHd5Eqw1iNIm6e4fWRQ0d
WBpdM2qMUI+acX/ELc5vvojYiBbUSSDr8eKI6C2D8Wb1LDwShQmqbFn5nUfv6pSD
hbj3ay70lDkfTuiNd7AVldCNIrO8IC8d7YOmhdthTObYbzth8Xu5uvRlNgrP4RnM
Dv6oDOyorf5230UUtFAeM1o4IV7r49it7cUxV4xSmLMLg35BBnqnY4oXWZoGixZJ
mAOFufliJj8PhhJnJccooggekieAgqzUw5aJ5SCKF83utvLN2kiX7RTbNyINMRux
KNJdmPmc5MpZSgE44qLc2mMCg2R/7sRuwm+0y/nDASC7uxNCASFWceK+Ix6kHwgx
IyQK4xm0C9H1XdJgWNAeDIyO3U/CogpJDpmH+cNLCqkI+FS08kgs0p675Em77O8n
8uh3ip5CFNjxTgtCyNrwUesNKMMfjFPj1cHApe5jalZv/YKQuAe329dchlCO9WnF
pZgpU7AlZRx5ssMwDcQ3M7eAkvLN3qCJ+7wE5lybXgxUzRuk+mUSDWI6nqePOCRK
MZyzpaHU6r60VNyJ8H/1LYa2EAZkSycAQ5j0pANLT3bVEJpWE2A6roJkIh08bWyK
CCm0+DgH7fDWEawkcfDfG7THoCsDUXtL4clulFtAeFSdYo5sJ8IDNF2Tnk6IJKwf
t+HO6Qjl4Lsrs+DDD0aBkO37GHhE/LTDt3DFIg296nfCH7xWkzm51mIROzbkf1HD
sd4ki4w9uQMjQzkltTc20TfuUKC5PkdY3J+GgG53WBBZQRKb01BCaF4Lwk3I5Z+0
O1ZzZsnJU63JXRXztxpEH9bxoUs7Yd2RGP/wihEle3LgVGru22mTdwmYQvStX0M+
2dlCaE5ry/3X6Gd4XrJJsoO3bvB2KL25WxJF48ZuIPPSvHHwvmjyFOG/SbN1y8VU
+cdlhEP/jWsdyBpVyXoVZHryLs+PK3AUq33DKhrTkD/59Hn95zgfRo+7ClaSJQ6a
QRBRgtdmffXb6roEu9m6UUyGV8P//AIWLvOeuiCwzeBiGxhDY+EGg1zYMOhH6qpN
ufQRcfkTjEwks3LWDIHvSTon8fnxxEU5zouRb4Rh3/r57kLD+15ytROH+wPC/WR6
Ld6J9Z1AJ1tMLJNakZmRk9YLaIQaDWbPN4o9dnjVxO7JDcLRHDmKwABbLPCNv8i8
wFRLMAppbuLWL2Mprh/76wAMNh9PFj8O1/Be+4T+LPx2XMPlYDF/LrfIgqTR6ifB
aTvtPwTeH9PfYONXY/9omOEOi4ZB+msEr2vBjpbMiGPVK1RSd5ttxlaKh8qa/41A
x22jm2hLjCsIeN0PatCTFXB3QfSdV0X+yTgy6L6X9k7E794Nagql6RD2WnGxsKrK
S/3CyQjYJUkUx3osABR0l6UzM94OxOv+CDy60Yoi4301cXK1XV6FvMvhIglcLouh
F/lKZ44GT6M+l1YDC45+oxXWKOksWHU/6vvn1YIpD/AkCLGjKPNPpZojiimQGUwV
RS0FIaati8rF7Yutmu5MzEyrk+wt66BDDyy9o8D0Eky5vmlV43oXw1ZbQbD3G4UZ
utVbm3VdxibBG8UAiMe61llaS56AR+SCVulurro7oc/4ncadBP+dUuwKmHtaCXWn
j5rHq45hywYSwItz33O/63z7ZKOx6QLzVX4TFpm73DWVnlERX06+WSZTmghr2W7T
7+BOlNoFXTbTVNB/JE4akOhKOSSvXxJpDMroWYags87CAl8HRmdtXSC0sex1z/Qd
hA9bOtHhkRVlTBWt3A/OAlfh7PSK/zqDLDJtOmEocBh0pDdYllFaHvPxGHlNL1xP
8AaGfSkj7YKYjSFp4udexyF9ipjhMlg7JrSxukqSfndnuE4XiXcnUOVjDTiuUunQ
cV2O2j8kGWJkKHQPsha1uq4EwLOpF+l5WmaWFzGPCVAgTsKqeFmtzbWujtd/YASS
wq1lLMJHdTZLI9Jna3Mr6HnSMzrKJilroXNI7BLc2feUCbHl33OfpobeJOji7pr7
26Nkw+2goa4eE6QddUHLH/WVCAkuk2bAowy6IoQGVyfo9rllHkwYbAqnfBSXUS06
DECHvKaRzaGE/JppOsly21w3mmSF8jrUVfAZWcApDVWh/+63QDjaerz1BUoKp2Y1
ZKKm0NXrymYN3gdfMnL8F1UsjBZTpbVscnIOxVKXF4gf/mwxO0Y3jyItKByBSTX9
Kw//cW796rraI01NmiOSwjHmI8TGOIws+VG9YxFYvVxJOP0iehPAIOZZXRVA1nnw
ihX36KPQb5l5Um0vDNWKc+W6zleoDLrsHDI5iq1vpVCR2ZPG02XQw10LirPk2iCP
HMwznJ5oB4Y3bR3wZYsRwHq1FPPm1kXFxLnCwYHNToW3LgOUuHp1XYBT6nek3JOJ
CfmIz7Yz4EjOQBsNeYYDt18GY6LnLGMlfA6xK5C1ljlPMqxOkk8EHpUmeZEi/M7l
eklsUiT7ghFJlKljMub3Q4LOyv4o2Y5+fSgE7bN5JnHyQu5CMwnDE/Mz2/XFm7J6
tvgkZviGXth75538MzCfq3j6wzd9p46U8hmq6LkusG0SHtFrjebe4cfakWyapTQx
1Yh6aAJDdS9FxAhtNOIhoCvlFaj1R8YsDzpH0w1hYyu4zsr7djQN137nEc34rBwv
dDx44/QioYcikdNjjHyjt/czpdmHq00bFr3aSe2taCwjHXbVegv3E3U7eiCGac3L
646eqVObqKzzZiCSEAHhvcS6bxUH/yQT+vDWxdmhbuCBNNRsOl8asyvro9uDvBWc
0dEB6JwKATNLtAuxTxKYgRQqW9/cHZEpuhN44kBp9zkfDm8N4ijQJF3iHhMpYB6q
Lm+lJ+WjepUHgXPBvLfNyucGOy9+6opR2J+il3ho/YOJ05EFQG5qqsNLOEvR7Sg8
5NmM/MRBOGWQZ0C1my5GBLLUj/S9J8HqnAtf4YcUv32aF4n1sgmkVWlnOcKFfBVN
x4s4hGZcdquZfQSGZp4G29AQBFqEOjx0lWiaAC7ARRXM3w5gw8VPb0GfZRPggKeQ
9Yk1MRMxIvIx2CAhAuOuKEcdX9RwqHMDCWeR2kyVGHN6BOKjplPVtm0LfjET1USp
KHjnUrHFDGzfB+Zw9GVzoQy3iZjkbjl0T5cLbPRrQIiKnyUGnnpCdW+vpbBsn8Qy
gOPpTWLh09Qe7B2HBdz5DNtUvjMy4uNbqC9wsorLhHuIyTabDJJbURWevvbNG3eS
XVzfbAfb2GGTmjXba7Ih8FwZgc5E8arJYE/R4Yq8DcCr5ao8neb7gbtRdxHtWa+I
S/4KsQEkfht0l98ouW/Tl+MiDfWRvzbvvjFaNy80iVEgEvPaGSTooPyfzRiit0mY
5qq0C9f6NXjS5he83T3kownRRKmlkvs6crcjSLvoW3odXVrmDGWlOrucNRWPvzeO
HD4rKU2E+z2t4gnrU0t9rKUtDVMvGVCPfpD/8Nxr2+7PQyYOLtNsbKhRz5uKnrUR
PrQqp484biHKGRKvXdanL0ohthqsmdJRuz8Ay/WzInIWOiWJT7Wk82G+tgQGPw/G
LKY3R9+NvnuAIlErVsYFIliKT4ekRwOHkuJPu13wGQZVakwRvSyouRymNkDlLF6q
iFUTy0nCLEbmESvITFd7w6MEWOTPQk0G9D7SF9hfsUHo1mjpAAU2vaQgs15TedCP
do026Tojs3n04JsDQpiQ8xKhn9pDR2gu8yVdK6BZ8itu1oqTN7d4atnaHxdwsAMZ
gg97t3uS0TxDOB9PGOMzAiCCNTIHqk8XtV12JTCiU6OL1gqXRP4L9e8pWnGtqqQ4
tRl6x6emGa1T2Ie5qaLnxZqiyhEl17jsK/411RVa39g+F+4exBVdnc0pzaCh47mX
zAL8a4M7L9Hd4LPVqqI9kftC4AUNt1iDfkrX0cHVEiDm978+xNifglRo5gDYsLhz
XqNQlhsZHWPNac0bybvL9shbdlH5jsUt700VZsX6s3fcXx1ZwWWZCAp/CtsjF4r9
7+K7z7a8bOdV++ZHW+yoH6/fS7Ni0YHfDmvf7lMW0srM+xAkgjHKK2SjTMH3wsXr
zTjA8kpxKbOT3HbhEdI/vbzTgVGb9c6SigTGh+1uUKIo1fCYDiTqInG9Kns457Sa
LOw1GP0Oa1VKAqpYxtUcoQm57oTrEVR42RQBXgQkqbGZ18Xls4xkTO0NPBsKZDB4
v5OTUyqga/aoip8lCK5Jm0Jd347pxddANOcH17qwwHOEE9UbpOJRZ9NY6fsRsGS5
1pEV6C69w3JJbh7wIgSOIYTKJo+NjZRIK5wUhabkM3t+fejk+62qR/dy9qCeY0/P
tWyHW2nx9j1Z2VjzWkiU00BmMxGw8xrWev6TQtWvLk3NP36zJku3BWb3YfaFrEy8
oBpV8/IbIk43N2PL7oLqbIt0iIjzQub/CLvu6xcaShM757zq0cwC+7DDB+eFiB5U
Qn5l6PeKJ8wvyxoLsYNzvpsIe7a2Mw7+6U8SUcdTMxJJdbOKbarH8ShyWbOc8BTW
BEVNu23tbrh4ZzohMhat9TyNjLTzfKIMzyb7Vv+Z6hLh9VUVTBCcNPH5eKIi7gp/
C7PwfHDu9kmvh3XvZZclJfTEbJHcBCepgPs3YjP1sJ0fea6NUyvWh3XU9Kag2bYQ
MZ9gVKkbWXKwk2eQrH1ZlTSDWnl8SLez0F3dUanHh3YSi/c/fVRoLld/aVv7Yt90
WH1I5qp4GSVMwWyUTyCjHAUF/ZZuHRgOylI+3O5RUbUNZtFvQwMuCiXgRPFWvDwg
Qo7th4GujXxdno2NNf6/ejAiCeDZfYKX1PvSQGCj5Tn3ryG/oHHBsgcyDcoU+J/h
PVio5CxaoJEEuoxstFMvv5PaFcfS7Clcb1b2dGY6e300Av7bL1TIgt7kTkpC4Wlh
plB76J4ADz6IVlXNccaiZH9yam4+Gyj/R59098Fx1BekKS9Cx0UxyIrDoNvusk04
nu1y8jD/mAG3Zc/SyCw7XdH7mRXWaRn/mD3DiBXcHhJtz8z1gqf5RPunkQAQCmx+
c5GmsmbaUYvkkj5fcNm53BYMQHANmST1G7HI7z/Z9QY6y1MFG5PMr+HtrvNcY/wj
8bv7gxe0fDdf7er0xtz9QP1oHSCfx6CW/aUGGCxSuNYN7oqfvi3KVfQT//81lzaj
sg8d+VuQS2IDB2RXNJwcsFQYtzwvWz6W0EDKN93Pfayjv7eTkdQp0c7/V8DrVhdN
AEm3MLnrqNiYqDF4kJ4MiMnKMbjiTYvbm4+uwjbhX6LfumPxMj0VxR+99tGKT240
sJBnXk1GBssLaGpqe0YOoVWxQS0EPib2DG9hFoJh0YaAAT+VKiYOiM05mBxSqFo4
1eOrmFveNdIm/TOzpnVhsx7XNkfiAoIUaE1CqypkYqKnmf6mP/ZyYR366/9IX6y+
brojLCIM7NsfRhccAw6zctL/tADSUL9DFLkQ4SzHRnw5E5zkcF+xQXGcN8v66YZB
OiyAUb46BBCBLbJv0+8u/2QDfZPXD4CIX3+4SfXBPRa2hIuoT1eEhdzretkexlPB
9LAl0g0eXSOZOG7P2sULYPtQUoLtOep/Y8bfFWan9rvAegoXINwEi1rsOl6Huyrl
LWBQwLTLqkOSAddyCQLKqK/NZl2jAEahyl76ygbxK0bETwe3glKMDASM2Qr/kvh0
cJlhjrsqFBs60JlqC2DapnTWa8XK2DRnilE30u/KkwkDRsqa4TLxiu53Ih5/YPQq
9l9J79KU5rB/BEZhOnwGYGLSuUgAsp/5lGMj3bZLK8dSLNGIZ3gK0LmYfQEd3Xy7
wFVLtdUcVhgG7ku7wXEoPst1+2K9NhOXdrj+c4svOBLXaJMkvmRi1cmRKSGwml9X
ifnNTc1Erxj25kTcYWaR30i8E59tTvc2xZBoSWe0YDw7pYCZgNKsVaHgRcaxYDCV
wDyPePvEvEI80AeV/gOhfh+Fa50d/ZeWJDM+LoIktBKspKoqisn/sT2vbRcRmh6u
vPOYCM5/tvRSn7BIj9tnbjRc5SZs1RcuMupFgc4DMjcU8vqQGmZWNCIy85x40fgY
lhWvQqY2WeEDrclsZ8V8zV0EZCkhtE9rQveBd4zsoOT6DC4BYiLh9HiPS+Lzzsbh
0I1DISmjK7CMgc0xHNsMO9clsBCh7nYdYrV31EGnnyWLYE25MB61zle/5ho6vuZq
KB+ZvN75rRHR3b59uayhsTwxDbMqG92Okk7vwY5rcX4MUuphIGEkwHXa9x8DYSwU
CNefdmt6QH6OK3Zt+Vz7Ste43kShaecA3L3X+w59ISKbCUlPqITN79Rv9LDkExbO
rOEWu1ouT7inKxK6tu/c0juref2Ukq9/NiElCcFYWGllSxH9N+fG3nkovgfhsY3K
FOhb2L7OnsQuVPQzn+mMww9R2TkJwgjOwHDIj31WZ0iI+kWSUnIcI0MJwM4G8WL9
x8bmGkoPhmpVtKOwcOPQMO3sGLESnVdagI/7k9YOFtxBBzIWgtYQiqjQkNnVpTJc
WtE7eo8cavZXY5msEGc032J4By9a6dx8qUneguFHkb9gshjbR2YWXnvW21AFKAPh
tWU0j98mjKDeaPRP6sc4VEdxLZNqznDeyCipEfiGpnxbYKZ24I2IOxWwpEp8e9sB
9FhdwU9cbGfVCA/4sj5xvnVL+BkfB9cxtleIR/56f00EZQGIVNBiFom8Q5QGcBP7
367fQo8z/QVGrgE9CQIzuXX+cbmlQHM0wRZ3Tixs58aQIHhLw8L7ZAgc3cF04z2c
StWppg2N6OmGEXV+51TDqpowP35VGsHV52Wv7bzzvx61/nTfp2YZ4so7D4WPS8uF
YVXUYe3qMCuFuj7JmryOewIZfn97Qmjd5U7rxz+i7izS2TKd1q46228Ah1mk0dVj
VABDAybVPMnbD1As4P7Dl5+28Mz9x0/OYRmS9ghEkQicais68OIUU9Nd1xT9/OHh
8KZLdjUgQDPcvXgNfe+RZOTJ/RWAzgs+5vgf/9IgkBHrSPs8GzR3VwWLkYc/wczs
bT9GuAi7NUtsQLnHlpmffwS8Y6Hc0nxKYIxBBNHqGxFOJah0aExXxvKMNbxJcSHI
Op3LfJ0XJvTKso98NQfJRTWo6MUpUAKoZH+xFWdBqwqIxi49l4nom9C0Txw0OnHP
jy6fQ9YU6T2vfWAg++AvdVk99HPWfb+AhH0PLJVEVQT9cBiPiJeVVIudW+Qwzfxt
CTIj7lUUysMo5lSy2WI7FQO1MDHUes9ovzISpHlg8BMZHtH5f7Ylhj/sXBje9U2p
nUq+PHWPxG7vyh8HeUl7/SnMuKnTzyfnik9fQdpzpY05J/Sl9TSAnPkgnHNwmBvR
IWdhEUNHB4AFZwOcbeVCpcViVhafnEWNJhBOrzntLkS8veKeam4J2H6ih94N2AYa
zOASiM/HuSV1TOsC4qJDmiFi6kJX47fL4b5TbDF/jp7HAXN0MffS7foft4bmztkA
Uu1y8M/2WrHyv+E5DIaeRiUuFfb80jG6iG5YkDqYJ7Hg8Ez9lRV7//voR3tcDwPA
Zqg8gZlih/5HH/YEiiAxBj8zcGMEKCaopSTaoDpZ3aWeRimzaCug8PgujOKGHrBk
jbwj8oOea+SqjTvrITWv7AQhImc/qJ+OeQ+hor8wntwEMvdLPmnNU5kGneMEbGya
Lllb343xqqhOj+BHS1C6HH2NIWPk3IjTN17DDYJ8WvPCIq2eYSgfVZ1DKn97PlX+
PyvmsKpJcVTG/v9k8nYCmjQqQJFTWdV3GNFup6olKbqyA8FCxGwS0+38FS0E6Xhd
+n8oIuTAaF4RELucmbOmB4c4DZBCAVSLdnlOpphmIJBPz58JQD7YWU7ApOyGfJzK
5j4FoWGNUhjpb8G1tpoSTYZr4HIEWU+R2mjzbLlHygVRwFpBwKG3sw9E4aAwrcHq
Zwfesvag6u75FngyqVNT6rFif46l/Rc3U6T0doOoniwRyXC+DhMTVFO1/Nwd9NRS
r8VoXHX8AWlz5SBnGjVixcC4MDTKKlr0w0pk/wk4qDT8J8VjfldGuvIXwi542mEY
6LirqSC+jLEQAx6Ctgq7ljL6/CoruM8HbnWMPfx8Gssr0D0QiQ/5VgGBHM7XIX4M
Xgc4R3tmLCukQLQfgmzRsWsK5q1p0MtYjUJ+kmlqDxg0tHoV9fx/wXyt/RQ6n6Pn
HNcH/oo47rq370KXU2LnR4Nzx4AVrZMFaBPE/ymxsG2VcdmqtX97wbNrJktKzDPa
zIL05O7A2X3XFyQaGYtdrNfDlPkSDDigw8uMOJSJrAuaaSvHrx5g1gSdykZ+7LOs
ZvN4Jdxm8UxbBesUc4s3azZTel+zzcndwgdvelxpZcxihKv7FifWM1f9LN3cDNdN
VoNrplV+P37yQ4j20NpQKz123Y3R5Lb5JbNUuEdM8vFwXfIgENfm6FOBo06gxC9t
W34mnjxDW5rSkmCFQl2opcDLDqgvr/3YOmzbaqds4OjUPFfH124I9EHd2fLl1zV2
VOXrngnISiIrtz+m/VKRRyLeaw08qztOynNQz5N3YmGXU8OYhCV83jcuEAJhwyTp
G3Wzxw2M8Elt+ors5myGZXDnNGYT6D49lOxkUnjkqdA84lsoDMXsXZFayoVRnmUX
q6T1utETJVvipF+Uw3zT2Q36dhBI5NkbPffwrggxPgzKJRadvatJbVSZPhibZg3p
5GZQXmXj+R7lv2CHM/MuawH+orwT1eWv570Uo8voUWQC57VLxEETgCMUPVE8ptx6
ti5PtpyRMfC1uJe5lKduV59S0+9jyt7EIZuQDhuTRa2M4ZbSjlNaAK/KButQRWqT
pnG2eNtk6nu6dsFnTxjbBG6GnSq3H7xH0THvQ0NRxohM8rWXB74VBFbU22hEEL3U
P1HRMcSq4WyELD+6vYXCCbpazBWrd/UIMn5zfdqulw+aZs1Zsu2tXXuIzCLvBR+a
KJzJeIFmEvxyh1u1UUTRXCMkb08y4KCspjTp0jIctZ+8Jcx1yNHDVLQX4CiLBFLt
fKGMPwj++rh/Gm4lsZ06otz5JF9nmNWheKSNBnZOrB+YEWvgzoLivCPGa9/Lx1e5
3GfU9GBZ/ts8TRnLwEQLvLWu/rKJa28Gddx8eYwrf0Efkue30TxTvnvIW/+zuPff
l6va8vz2/0jKF5xQXiCi/uRSS+gtKPw5vNEqQ1xRiosncVf+Wy7enD4jKYzLY4bG
qmM6JN3gNRJ3FJfRZwqMl5ku4A5tagl4Nj/AwS9GkOdaiSCbPYlXqTw+5h46vhBU
PgWDntQYBwoNDX2HSgvbNc7362t/l5gq0DihAOosZtToNzR6zQ4+a2IoShJTjstt
A1XvViSDIjkiR2y8KTERHGthRDdTrw4uDlGz+Y5jtpWx1puiA1zS2g3DNOjX4Rlx
UBtHBAYHjkXOMcDuSiMFKYj6wRyMhBXErn46GWpQKh1FebL3kfjm3Rkf4bV6K3lN
jT+MAa6Raq3Z66+qtGhCoQVit2mG9KRwsIuxBDLZUjGVebzP0uuBIKDepLX1hmeZ
nFc/aoNY8g9MixiO+CZrE7X0sF9AKg/9reswUyhmyt/tGn+VjP565Dwx658q3dW5
2Y42mS8p6ppFcX8f/1PD6a4jbuLNH9VskievS4pD6OoIHVfZQFaI/DxNOOMmxhob
h+1+CKvXTEiDmbggdPndxYpxNsggXaIxiFlyb4gAcX4cJs97M0hjQIL71GpimQs6
Y1Nj+PyIJGA9lWmDj5LRD9YtD+3cma9MfWnIZcpwUAly0eZpSbjRnFgxunKQOTsp
Ou+lgSVA/jkEFuE0xy/U8eTUCzP1kCXegB0tupKRds1rjLUe66g41St+K/OXQyau
Qv2vPkOH2RV2DPM7lPODzagqynG3jrdFqy2cE2grgzJfuN/QPj35eKtuRLwzTXWJ
5mmgG+ZoCQASENoE5bfpNgvKZTUiAfkZenyBl7P+e4I1vgOsmd+T90Qyj+ySv7gE
M84oSTqiEmg6L+m1SBk60baJ2f9wOeVaS8BOq/VWZ6NVlXAkPSqkrJJTcsLHZa94
IxLJIkFnIWawlF96m0ijabNJg4jIgCrCJVmoaYhgd5HoM2sDfT69jCOgWGl9AJXX
NbxDfRd1USjsvHmHLpwgd9zUJwiYt0XPd5SPTEN7hjnKA2Bw1XAkqhwpAqGW5Z6k
A12tJPgLhwu3FBygjQ4gpeTwcX9TxDDekOhmTUoH2kN8vEJCBhZ0oJV1XMJYLLvn
kAXkAwNxiOdv+tGHonCIWlsh7mraI1MOpa6w45NObW6sGb2PwsWNjk3DZc9dgHcU
uDEivR23NFDf+P77hdIi0dAxBSoeJFsqHfjyk/Z34vOJKcLYgl+7Dh062z3U8z4s
AFQPD8y4B7CZkMArcYrw9uY6RC5qzpo7crnHZ/6nMCR1gb4h8LBLfd7M80dcHnxk
UQ2Wg/xTNxXW9OjMRtruhoblm7DShJpTKksqHRUVLsj3iv480raMn2DTIbzCztFp
TYNnRx+wrTJcH7FVIPendURIsD66aGuf7UaH+8JI3JMez2MNVIBPmooteSB/uZf0
Oyb6KIDihq9I6GDKWdTmGgUpUOkXkXkaIixng9MEzCvmKt66PUmY7VxZg50zCHNQ
YUZ0DgK935ke3XbKAJnBZh3/SvlR02pkSd91noEYcDNdcRHP87cvMhbMoPUh9oqG
sNOYLgNipV0HozRTTIM+fmDlgxsNIYl4dbx2PgkzJYdxG6YlD4OgPpm/6u37eXZ8
4k/XZgpC9EXoj8LJV4dut2XdSNm2hsh8NUEKzqi70MgXkp7sYvruKugNNbs2gGcq
aDD54UtMkJ7Jjm5Vj6yoSuzl4LJ/INLnoUcn0t+mwKvWWk1IHn+YYqOtQbZFqwxL
r0bbqRD8rC4Ik6JO6uRIEEmSiffipxS7Rpfasr+jwd7Mq6QEvtfvcHurj7yJ8loJ
u0FI93YXeIP8dwGrJ0/G8Vegf3oyo9fWzbEPmJL/evGY5FYB9ZBB320F2/qwcZCT
J027XrBzWn96ChDcKlJv9Yu5+9V0dS59+Hg7D5NTYKAA3D1TjRNsMjAqHhpBaiNu
UPfDW0MCqSqqK/IhyD9Oja9rGBALGVyArmdfrKzTYZNrtHmDVCohPHy5GlQjQc03
lqWqJ3e7mfdhUFAWE5zaLa2qFW0RlXClJZpZIRJNNhEbSzSgzYo/GUydSD8R34FY
+9yRtbcbi2iqsIpxDR0ZlB7c2NTwMIc4s/wjY7mKsSHSU/hO9uxifnrcXh+qTRQH
j4dPVxrfHryJ/t+H8L8W1XxDkK/svNM7g4Do36HMfcoBGSI2oPck99HJTxvryN9r
MkeNTYWV3mnJs/q23Rp5t+6gxEN0cStt5+YaVGpE3DAotmfLLuZtMOwKRvYkJNXv
l0W1KPo/gp5r3YrR2WXk88kmkd4GCzxVY5Kx0njQz89V4/Z1GHYuo7RBNVc2Zi0o
+KRcnJjgmv9ll5F/F+cxvHuBA/xUfIv7PG0U2WuztC3Dbm3sml81UJ8vWnLVxgM5
O6e/grINpgNXoEXgznseIq2nRYvDtQXOOJxHsxj+o68N07yuLFhF1VOjbQ85tJyz
xqzUCWl4SxT9827qfPcHg7f+l3wxpx57jnqDQyte75bQfgcUeiEuOjT16rz6JASs
Q4VJPOqzfGUkCYptJSMwgr9RNUyYTrSGqaUa8Fw0dL+yQxIAAp1d48POY0Z9HAAD
+on35d3Vh5x9ZqVwlo7kZfe/o54vAXNJJ86v9ZpkD7WXxFQLM9vMM30S8Sv2cM85
Ziff8Dk301OhUwNaocKDb2Uv7HImgNW+Ct3/KUJtlv6Su0a+VTo9WD7myPu9HLz6
nqROxOwAjs0vQakl+Fmcz3cY/VruW4+9+marw/6+ceqam7S7AK5SKLxLIhDLXS8S
RRvPxzg6W/C7LZF5fD3WPAVMm1P44tswt7BU+PvDM7DeOE+VEWjaeyQwSoxSa6sP
mEwLsJCUIw3xxoskl8tOr+G7O7UDxzrZtsrxA56fdUZdLjXt56VngLiz2MUSNY3O
EAGmkUs8yZ80ka2dYEho6JkQxZerIV7P3uHyFgQBqQ/dEISSRB4GjrliCK+MXL42
Pn1kddHIN7zqZnXkf2UhFTJdD5fsyFlttvn82n8X+2VBJqAb0H96aPYcL4HHEJX+
/O0KdEQCdE6ijFtOAG6fHl8kYgu5woKcwnD/kaBU2QCxpUSfhwkQkFpBQJbXAZ8d
F69xy1EB+NyXkcWfZNK3KHlbkUYjbEaNwTqzd7xI5uJ1hY9gQpL7D/+xxwfwtXaW
YvEMl73VTuMXXrQXSTwisQ4tzHKVtZrjefSUZJbPGcn1vSOr5z5Vsk5qk3VuF6/B
FUWI3UCiDsTOwYGlz2naFMZtMjkb5X0ImAw+AWqJAS/D+9PEXMvf8iGcQg4+8Dby
LcuKO6tAWe9NQVUpXasmz3AaT85hFunTZ0kRwyMWRXEec2U5yYjGQBC6LLL/ULhX
ku31Fp9nmg0ObEV5tWkhrtUkhH90o/3NASPZYvx16J7aRHDOMNguUhhyUNFnXl/8
7YGwlL3g7aNCQpCEceRHX9XD7TK9HWV8X+GJ+8sAyHJIYj1J7OWD7QANRkNUhz2k
l3BZM5VaPtjZRfOb15G7smz+6Fp6ZHKqonJGNYUtRVFV5b+L9LznH/3e0XUjAnpS
G6ZIFXUlnxvd7l/PTy0LBWb7MZO6aNp5lUQKYiIBLChjw6LaxWYJ/f7B20/fT0vI
RjonNZQG8tN+g4Mb/Dce7Gh4BcSReGJRIHUlMrft3RFgzfm2vH30He9GQiNlF0vl
eUsJQdq29nv/ljTK30X3dA3K2qN2cOF6e7+WyYRzDgDQD+Dge99T1OhkTyDlonRJ
hwnVF2Wz5tfJsY2I8bh7RHzQn/C4mt9oqVOT3ja5CumnSdTC+or9PD+1B6oB3dwH
KR+5sK5eX1hC2Iax7uXayes3PwwQd7N6sFVplBPgvod7TvM9ouAFBy4XOhxDpcVQ
c6wl/HOTdTXJutLt31fEv3z6fuO2EQy+Vf9kLZKNo36I2pXVfSmbJPRtZj0sfFZj
xPf1rpbW90CsI4IPxImy5xj2oDUXcjwQ3tn+9++q/+u7bck2WeK1xdYlPWi0TFcr
37tR4SI+degjIZwgj9JdEi03OPO1Lb69HDaW/2ofBEYvY5+mSKzTyRakQcZJpdch
Zfjxl+wgfifFLyK3WzoyUrYJNNTcpuc6lSk6pGnhwC1qNenUPTAK4G2l+kWFJRfJ
RNgYMRtT0P57i4sooJ713oS3aPJndLm9fvzzkb5e0NZkrkeMB/bjTzMu7fr3ikf0
NDP7fMUskbGooPYfZfawCVifTp1+G/2JbNjhd4iNCIIYbXOVPTGzSbvYqDH2L29Z
njOt+uEBIkMN6uEN5PMoz9997IB/HawCg3h7d+tv1f6VqeWPFgaTmdjfZhhgPzcN
S65GKXsQcaJZqOaBumFyUi37U+plD6ajSaUNfFX9/NsU7gx+kN3BVBSCImCvooOV
Q7VkUUgHw5zH9aTLduvM7fna+UW7JgY7SXUkxjgN/HkXr3z1lx6m9635LZDxdxgE
795mU6/4BMTJpapz4lbdmyQ2PAAXYvnBc1tAyoO4Ri02zFNAyOY1CF7C9X06ky/C
AhPwEVBT+zMvYFHIjwNEJFQVJlRnQZxemBRHCNltl/TeSt7BMC44iG5SII28Y8oq
WsOIlQJ1Jxkc8yCLwU0hTVZAFFHvDiXWHAX7uHGSR16jiGBCLIbMFFerzG6UwjiD
oJSw1uTNULUlQTyzaBRy7gPEdxBP1LpHJUq7VZMoL/DYcffK8pIQ+dlopmnFqhr3
v2hhk4O1SpUcHu8C5O0HxJ58I5s73cL+0eU043uWcI0bo7rPf92ee81GBnh9qMQ8
RFwsEciuva3fk1TCcC3X916CGWOZWvD7jP9zX/VboD+1ppcOR5cd7fqAsK+84yzS
kUubWD5kZ/V/DGdu3LSqStvfjcUu5GI4Kaisg00B1A8R5wv2J2sTEUw5LSDnIrz0
pGD780BdkWKlGEx1lYFSaRtH6Lc8MlNsd7MHLetp7B+rse+O6GUtGqRbjqQieNzZ
kgJ9Hruj1Nbm5HeTQL21M3XPGDHKaLit092Qaa2nPjAZt049m4RQu4MVSyfB9h5J
mnLFlIDAhQhVP5Lo/lW5w8M/m+4rLWf7KP3tfkqTSR5J4s/LWmn1+vgqn82ooIzc
ASDPUQPiHiwMMof33T3mDvnNNyaw7kQEDjiG62K39bm801hGrX9P+DaKmNWsh5AB
5fcAy5p69ENn2ee760vN0wm2AR/U3VYuMJtVhaxFj8lH+5L2PqZR1LqT3jX32A8l
omXElbfe20HekvW3fd3QCWjkoX1UIrhdWxvvfwRlP62ZRd1Tb+wP+SSYvkK16ZR0
DDJW/Sn1IISlja7yhVQvYgbMrgm9KoMjZPBatCKmdo1W8QG+ANk+Gb1Ui/Lhbjf/
mqod/3+u+wB2YVZL+anmis7PIXxS25gGdpp3IM6yL6hW5h35raJH0HASFzN3fWq9
jJVuUHAg5LhRDLANRAUL8ohC3zJKdGjgZk1aJxOOgHAFc9dIvLdz6bS5JCZwAopu
LdQESCyeG4QD9baad+UYIArY6VhpNSwRMaycdCW4kpqttpGdzeXHInOcKln3nbv7
5xpvN7JWCbUWnwdPVY7fiVyXvrecihq7js7JeRXzYaxqD0IhgRxfxFF4saa63HWP
mKlHy3Y5vAz0UD95rrjEvUGbRM+q6SDp1c3L8RSRhCcnFHni+GB244uKgOX3AVs8
sRGhumLzveduM5c3rh2S3zRLjHOns5WrefLIPxZSaD2vNSiazvvzzybgAb5YSPNX
BOqC8WUwssEDkxGFw5VzC3164dC9jEt2DAJw1Hx8ryRrZ02+KeDkIfUqlNTyKF2O
VvobwZ9mAzQY85NaooVzCoKdur/IrABPSYQpyjt/10n08izBsP90nMaRiIC0x5co
gh2hAwu/ZKYPCpy9X20zj70AIHTmklRF4uv0s0KhpeC6hV0fOUWlI8+wJSTaE4EM
DUzEb9cJOuadOCvhwF7hjCVPhuQCLFWu3mQuTQ9ZrqC1TdkJy7Zk1v2J+9cneCFX
wFFg+i26FdKizKSCNi25nNQuFE9zZ5w3NEC1uwUWEZQguEi0FUIAAUXoF+Ht/rwQ
FxmCFGbbReDTZQ3r8k70gfldio63kWyKAAwQXKAywRoYtYvXbAy9tBfEWTY8JdN+
g4NCdve/PFmYeb/fuqA5tr5+DQR90i28k3FhH9ntsGyLPw0z+8KYelvmS7teSR0g
CP7zi11JMZEBGR4qkZasZcTow6HL3hhBrZqyzK7WnY3V9kumUnW17mqh85ra6RAN
e6QP21EWFOQY+VunIMCfOtWkFOcZWxm/T/OD5tCpjq811D9fKsI7tKkA2KxGGLIg
CawfTdcI3rBFiqjOVvKd6XJq78iGEkX+nOthJM5oSrsJyUo7R2J9U/0w5B+0yI5W
ersRoDBlzmBgl/8fTvavRByzULawuhH92A9goQcDCDWBoL8xJj95PafR17C9UJ64
jiRd4pG4XwxjrUxuuTC379Xs3YNbBB5fdqvf1bUdsTT6G3Fg4mkMwAn3kmyObP4g
00stDgJ2l/K20dMxiqUgwZE5SSQfexZj99jMIWWgNw3ujxMD8z2FlRXSTyrEaVsr
gGwWzDvUk1j7IqLUuWUkpnJQ4g+xxOYZIeDJD/jTNCJ2vmy0g+tTAvI8nCIlzWUT
54FXsCiX8+dEFasz//c0+JxzfkS5awFGfhIS8EqYzLY+W32AxiCsBdNDiQKYlz2Z
e1vBrLS771mSkTR12e+j1lXm8kmNNpUfB0apv0h9aqwbnwihb934Uo1eAmAOKsQ9
5oBgC4KjxAdl6GTk7b8RCPghHdYhfP++zz17qz+59nhKu/QTsrim2snraGP2H7Ia
ytUKRxxCkNc2IYBOWGsEZ3XeL4uaKmrByAIngJjq2F0R1YHVCw/yU1myDo27o/ed
KLg0R+8xl7hFoZ3NdnAi5xsV95hwCiAnHqjcBzGbNdGmNHuCeSOVEKRxrvaJq0oP
EFSn6v0GmHlHgQp0IYPVpIbnMQagziGh2+W9mD6SsR2WjBfNJ8mpxDBjPfYo5S64
LQW5rORvARItTikEQZF/L1alMqBquhANYvZXgRFt+yYfG8uqn4JSLKsdiCPRwb5b
ZK0o32BExNZkf7V6cAVw0egB2LBkQFYDkoo7q/GUusS71yfJBccpOHjo5oEr8oeH
HvkM2pZk/N5wdZ2ETHQ01crQTYnKr6mlRmblAyU4z5O7Bt1G9ehZib2y99HtAz11
HJsKUJdgcq8f9FDR4eSfrsV42+O0XbLbe/FsiWDlMYN7WDN+ZHLlhsSsztqkfroS
eNEHI4Gq6yZwHIyTQ/iScb4smqgbK0nofYjCUDAI3drNqAZRWlyqXi5WAtzkQfdT
QdUd9hPG9JP1fOuJGTmJIU+fLXRiQ8UbxHcevz/2PwP9qy9DacHptxx6+BnY4Y1e
2qujErZNy+PSlSc7txYhMV+IuVkgIHUryzsseaMcryuSbeODaR3Q/qaT/Ebf7XHP
cREu0vdF6rDTBOTHIIHz5h35TPFuRVo4AO0kxG7Z66klJz8a/DFOSmMX2C5H0ms6
su7DKvWcdV0zPnaJi2geOIr1iqi+MxkzFxX9I8mgDyovF5dTqjyf9HoiQ3alRPpG
RK+4Rj6fwdn71KzaZt/6XqMzCAqHGcm/rzPgWVisElcjvagQ/eSsJ+vZ4SqVyKYQ
62JmxV7kEUUFj2gM0q8DEmAItm7WeprY74nQWRs2s2KIb+IfmrBdvQ5U5AI2j8X8
pRCxmNPHs4NZGPR/cSi2+X2B6pW5cIDyGfNquZRjhquOoE0JMnObMmqtCywdUQaT
q//fED/aVW3huUpDQNASAR0jND/nn1VBvHsdhDGmTgJrjNfxzlLMVBdm4hr6urLU
Y42wco2yJ3BHNPHuX6IwQ+C1toQLTShqWUwrlrw3AjHyE4U8BAmBs7qc/IT0wT+c
+PVZPgi8ZOhPlDRwJu2bOhUY3mpI3+FCUZqiB1gfX8uaaqYy4MGen8DQBt8AjJPs
mx69o5cW8qnvmqzVnr1AU5FcNEuFqpPhRoLcvUqTry4QcIPoV2fI78tDTJWj5qQW
oLU/8CBy/yymqS7ioH2NzFo5Vi2993+Nggshd5SffzFCwmNdi4GedwI696vqHURD
qXGFza+ZKeJJRti5TaWyuU8yeHRlE7aSTlMVBZId0+6VYXQXeb2IQVakd5etHL6C
GY/DVUrJ4fzrntC7Uzr9sXh6LrfU1p6Q6qXeRULYac3+tDtzt6/P8AiI9eOi+kgz
k3mtuYic1FM3/k2vlrqDP+Dm3Eu5qI9z9j2J5LV38scosiYPI831wulUXp8w4h0O
ChA3MTwPK6IIchY2PPuJc9RqHfbv4Bxj3SwSbV5ZzxHaiPzXWVP4jG6YdPq8Mjxm
3jD1iXYJS+Z7LRT98GF8+5uJ6upI7tQjnBddwrKa2SZiq8LEHD9PHcvyjdLjXvGX
Bt+0EzLai6T+mLreP5sclhXylfO6ccyPBEPndWSlrTdj1VI6gZOqf+TfGr168NW8
w9TKwCyUKShMs4915Z/VCACDdimpWSmadIUOiW/wvsbZRlWPPJwFN+q2yC9Dfuj2
8edIIKTEM2sIwslKZS7rGFzX570oEfKdTtEZioZhQY5LI1P3LmSHW8UJX6DzxO8g
0jq5WhkTzIryHbyEauBg1XktmVYQ64nW3n9aBTirmRfSmlMdY+5RKhbL4jcmNsYr
Rn8WOXhy2NC/sfCZQEAh+ZWzdTLq4RyQO/rtekEAXtfZcBtCx4tFYNk6Iwes4/UA
b+lHcZ70RKHejsmRFjmMw+ld97piEHKgxnw301L3/hceqn0X2OvriSzx3w5/2Keb
4dtJf5wIAKY0JvOhv8Ku8MA5tz1MCioCDeLCoH1nfz6NzGm+KHqFxU9z5sM83Xn/
L+46aPdsVqkQWi4NvXVYp2G+MDNTlCku3oH+KTEIJDQBarCeovHUXEHDoDmaabmY
l2dTVoX4c+aXr4Enni8Ll/ZAL0MS1MIogoThT6z2dE7VJjQL4PnwZXXis242/6Kp
DM+k5XfTD7xcwG8x4G8wJBX7M8DO2F238m6OA+qvx3JiDRwXcBl7nEL5b49USR9R
g54xOOHRrIdaMP8t7e0UY8CSXNS2n7/w8s7xk8jAf9Ksdkjy7wH0PJWUOAaYYNrT
/Ig1/SnuiMUCSWfFL30a0OED25DhE3rh2OnW2Tx1xUeckrUUu4V+1LRiaDhEAYNf
JbH76mhNbFG+P7xQeT5dqgHw9Rci6NIkmRoWOMF5zNLAUhz19oalcFqFjuTnsOo4
NVpd0FSV7MFFuX+qZSx6h17xUS6cF3Qbcy1LeLiSjMac9E/NcBMUcecOEwXVQMHV
iGhydXB2k8LI7RAIGKhVSuICSHSIyljVVZ5ans32M/UEooNMUJwOhaHHDg+9db3G
/wV0TOVDt8SPPPKC/DHL0SZ6i9amF4M7h+rkQuaZeSHqwJ4G7XN5lTNCPC5G0Y1U
Ci2DxhHcF7SFFEGeKLghmJF5pj76XWCne95xL/Sd5TtWVH/YPVXjgmr3fd49yiZT
tM+2lhsPIjFprXK7OcfJcAmekXizUNbvsoeL1sgonc8zbNB3NoPcJaDwtTCyL8e/
hDS490xnQX9uzdmUjBkrEPY+KQgcrTdeYXh4uyHaMOEVJPzxF7Zq68lAhP0fgFuO
xD1XBPpPQObZEdd6Y3gOivLSqlZazyrUUY1xpaKAgL23F8AfkfhSc27+vGlYUJdw
MAvLLDqlwylU3HTKTNLi/xstj38t9CMomtKsD6Bd9Me7zbSLO/pdai2KtEXrT2d9
qO3wNURg6ZWeng4OIMr2ssnoOTS8X1cTIixwa0ebMSMbySkXSiJwVyL/GMBuW4FX
tQeQcCCIGAq+7P0HG5+WgkLR1HijNZYYIbKHe8VA7/U4RfQfO/RlzqqtJzG+ezjX
HDUkYR7IQ0Jd6ygvVgTUOTukkV7dUb938XNDZiIIPhQpi3EMBGansCKOpe+SAHQf
dzNs4frO8Xs09bxrOY7YOAfViQAN9dFMUlDJExaAtnfBGPQBYYrVyjlaAc4OOFfv
fOj/wRl2XMMjYr5vfLhL+1OhdMAwOm+vNjnDcRh3n6eVCtfsv5afq+25uIIgmwXI
Xs0O1Ep8RFJKKMVpKJQZSMLpNHEA5YPkfvKB9vyDngTzrKiJ1/GLc+6XXMkUAM/s
O0OaCtk215+aqgoBZiBvtM4w2sDkZSP4VzEExw2IVAKsOlnxHygsIMchA6+GABlN
8WVQaV63Ioz5pYLfZym1Ex8sCEWDWY0ovkpWsdZQ28wXjrCEHTLo3q+bvyeIvDvy
4mAvnVAgfkcbkd+zSbRC4TvtSUzwYIw3j0kqIoR8LeGo7Tn0dN4gUSnrruwHFWcY
L/pk4JfRBDwaCgoP5tsm7Q84wODS7Ah02AOP9jA0UzcX/ymaPrlXpsd6chgitf+C
6sH0/KxfD6KlDe8vQi+G6Lng5lyMz1yDsgvdvSVr7YU2R71cDAQ9JfQKNc3uv9gq
CKyxiwa9PDrYsF1skf5ym/UrfY8hAhuI3XDYWdDAozWANCz42ZbbMlzAJmeHPka5
J/eRfLKUTESN/jioKFVOfgpDAvbPCb36kq+u41v9hTCLj6BV8peh56uplN4v4OyW
4dngM0J+sT008bPeV+gCyFPZWSKHOzcv1ojz7euuoigWYw6HjCa6UFlw0QBKRqWg
pAsIWLkU+M3SMTWMjEujRT001e/z8M3+7G+CQ3Y2v86ym907GhYCxNbfTs97WNxs
ZAnxllYC+CxaXLRzB0jLh4vNaMGlNyzU52LyYmS1b5zoC2tK+yVe5sZE9mFWVwTp
0BMYYA86uEa1lYEeqRicn4bjIY1qT9M6P5WnpMtSXxXzGQOGiTo9DWVKjZbfq3RO
aqIPz1uzaqibCxrYCDU9T3wCdza4Zwwr8Cx8amWgOouStfAVdCKwxBR+4jhZwZGW
V+Nl0P8JgVz2aVskM1NbcNxl2lKs+1WRxWg5J77vVBZ0QXf+k4C2y0jyUkF/M9BN
7RY77QweNMBYh3tm0Ogwz+H1do/VEkq6dOx8nFrAaHN9OwINlTiV7WXkSyQhbGQC
7HC3ojnKRuC27aj7QynK64TPzjORAhzmBiEmojxrog75a9I7wlkoPCCMQ5N9DCe+
Lq6F+U3jVT7S0b/1j2wiW8NjWwNZmZ9Gq7dC3mUo7osZFrrZtNqwpOI8knPHgKH6
WJHl9MHGiKcUCIr9tn/dGZv4m0hP2icgCvrUMn2NDl3kSO3Yz8VH3gZpNo0XuyRp
0+fuCM1dDoBY9uvcDlg2Q+JCj1/KI6eAKUPZZmK8lydBs4kj+9RhGDXYsdQ3X8t2
yAUwC4vhTmqUxNEcda1POJ6AVDLTE3TTcAZWdasrZLau+jsFKSzWne9+6Anmo7p8
d66EJhKC4KqkiK+ZG9iRlPSybrzO3ouXpa9JjRe+0WJ9+4WzpXs62MiVYZTV4fQp
TkUPJ26IYIdDzX7JRKEXPpxtY2R1gwGHuvLN5zqj1CN3vNSBszxpurwLGgDGuW3h
58SjD8PNu8NsayKJdhjCDe6qdDvTndUx+YD1aUIQ97GuMtgzjDTKmIa3QH/X2wDN
1gKGpQhIjZQpx+XFK6Lxrpncsr29FbH6J2iFqgC0Lg2onflhr7j8/GMarLiWGCmb
NEzuZoK7HKurcr8Gzojv9+4ARYkJMKOkOfMo9h/AX6N5VHgsF2Fqv3dGF0Bz/Exl
DEn/kJwhWsKs7I4G7O5RNcWQ7G677FcWIlORcU9N51WMf2L82ekm9oUqBWYyTmbt
hTscnXFWpJ1OybITAWEa9f0WX4VHD9snBqfE0EX5KZq34/sjWHOPVCiUKVwnoOvY
UBRcuIIA79YNc3r1XIxhIdmzw8Cq5IwXwthLYggBfGTvN8uyzrn3RB9P/YRhv8Nq
qjnAZN210pxbuGr0Jnu8SBxvtfwtzNt+br75GIl1XdEKA9a0B5JecBWjiJFE1w65
Fi9VvBFF0BSUEnWiWr65tJN/PI7421kDu8Zie15asqHZba4yhAAavlNBuZH5k//W
4hxcWLLFQWY3zM6fvspdKNTkwxvcvh+E7YVFwe5DiCYzB1i/25GO0T3jRtc5aZt8
Rj1C7rRwuK14Eb+jHNIEiPddzG9fe/4S1fd/4/dmG9ond0IT8GGeSS1AtvJEUELP
5ynsyiHL2pq1iRZtPmx0HeePauJzHuwFasVzBZb5CWOvqwAwD5oXWxwM2hv+XRWe
I2SxuZKHykcL0AyfwhAjzEXW5LNabRimmEd1pYVM/Rh8QE1DH7O4OYFXNNZejpxx
hUIcW8gqs+LR1fpoHZf9vMB0gF2XIYVhMa55IC94/FauYGQp40liySbsIEO3YA24
BvCWCnzR8J/OdPPYvhHs9MBo5QcKQ4RLqx5T1MmwaozatYCtOEHmcU6cDLwWmfaC
xYFFSEoFByE7CyaVlNiNyhjTkafcWTpqBgWM5f6IbuZPf56Ed/8l1UJcf7ez54cT
f2wTkp8yBJQaOMIpiYm3PI+QRaCv6nPF/wXix9Gx612O6HOxQ5bzYLDdmoL0MiG8
HROyzblDDcfI0Rp1nw6b8i1jrVEdL8WsKz5p+HtmGb3mnp6CmW4yyQJKx59ZU0Ko
M7VX9F0UB0zBEzSDhoPijl5imyOHbsgfrZeUVeVgw8wZCO8WyQTfWCvYpvNl79zk
9PcDk6LZ4XpWJAyXb5dXsF9V4SZ40OI49iXV/KyPl7JhI6mDoR/nkDpkMVT1CkHq
2FOHn2eHDfnpwyg0VwSgviYXQ7nsG54TM789ncWg2gFywYi9GFcwunGSn5yNYJq1
aWK5avCLSMu6hFnWWq3udD4p9IS8857aGElAooJMADnTpy5hUF5YTpfqVmdlQR5P
fD+psn0w/AIqQY41fEOPLnioNZ+hKIaFazo19/CL/i+ZznMgOMrvOv1WxGcQJT8+
K23Thq1OM6lRbaOCk4YW82PHYgl02g6TRNy5Rmy96/BxiYfUSzzUOZqO6P/FvGTH
G3/nycFv0kPSZZccjkW9lGySH9xB8WkA0lBNYlPykFo24FIC9KOh/DFmBTiiGI4k
KufKK8U/lWBxjO6gE3/CRYBPqCv+MPtHasfj6W93ZecYGi3gea8bh2IBukHzSNjQ
vPUFd90+4iLxjnenB5YnonH3kcKQV3kBWG8fY5kSOMyPHyiI5U3RDs7nhZqByhvO
AMuOQ2sHtSjeCmF9UtgYcw2bAH9jrZJXnIBKX9BPCYg2UurhrrCWBXwoyWniCWKa
Y+RSRPLAlGrgOkj9RczB6JkL1MK1XeFTIkOGoQxly8nUbRZ9k9ROnDca6cb5Lm+4
nvOJTRmbe0mGimPKxdRvFgyVf/OgSq2JWg0sh5eoSiuunvMrCl96gkSc6Tp5yr1J
a0RBjXbis4ZcLV+5Aab7phIihz6HFZbKgJlnLjsbg1hSz8Kp2XrvaSoDLD3Epr/e
DKuTARFXTzOtEHal1n1LUUX9qIiOH7RXWDQxkNESrYvQDhV4LIt+fRB4C7f63Nzb
kgAAMkRrqyBmvFY2HIYfClbDkNg4sSI6PAaeLBcAYPSmm8ds3updcKfu1T1bc2oR
7r2gubmyqGBVWTqyGeQwGcrE34crr5SAvDzCGuD3s8wQJ4M8lYBpwA56HF3ChXTW
BpZdQ3YewCL7LZfzJX5f/hRI/CDEsyuBIJeI6KsVsFeGeJOPZjSFpuEMVehBRs4R
F16j23a95UT3DXAwa/7no5j3X29pl+a8FKXgU7fKHYMspyJzlKUNer31xNP8hI5L
4ErjaJzXQs3uyQFvVMkz8bGr4hRJdM7O8dnJloUlIt/jU4npmxXbsicmlr95RQi5
5f5ST4BPuya7dkH5S6MAf4ZPwxipUEmL3QxKKpT0A7IupaE07Ea7+4dAL1cHIqd1
jzmoGmt8v2o1gCmMtelgByz5+3Jx8YV0Bg/XEpCIgbpVMOOjvLrqpLpQJM7L0D7b
u5Awdg2gKJfd43zgOItvMulTeFDkZChRo2Qcq1RBbtFJQnd22Pxf017W+DAd0Dwp
7Rs0b/tzNDBAjkOIuIMgZfG80ptitaesF9FlsGYaxqFG+TQq4mPcH3e13BWT/aXU
FwBxtaNH5aGmTb9EN08OhbICt+JzbmwzPzfrYzvMg8OXg1kTVNeKcdqUjz2zbFcx
cSNL4N77ltc5WcWybhg28luyhVqGX9DgV4XaD78s91cXwBboAYCIc/RNAVXu12Gc
ZgHJqVL0HRzp2QIZxnwuEDXeWp7xRjL//lfEuvkbCclOY+tiI06q/Ko5aKfEVKMi
SAxOsMfr1hav+b8wC+1jKl+Zi/Z4ZikkKIuohzh4VDEbFlJClkG1KQQaiba1JtGv
APbMf7bywDUYzxb5qs6aDBEq2UlLU3HnNUml6Yz5Jr90D1bslFlRFSg4mADuOD59
1iqhn2lX7EglPKmFwMKsh4J+7Qrw772CicRLLbkZAm0kQzBhR4jX4soPpPCtS6Lq
5Cy9Zd2nuBodC3imH3XzSZbo+UdSPHOU3kO7oh7yPg0axHaYKisle/yBR1zY7L7H
4kdSJVGUfHxY+PFe+IzK0XKMtu0NEeFKULI4LftFW0Pw0Y3M+Qq0GtXspy1kLEgp
Z6U940XMuQ111hUF2IhYqfPw3SUxRXL5PGbv8DRH9kmYhJ/yyPWM8gHwshYXNrAR
Xei9V2xe4vfUzA6iPh//g24v5Fm7DZmPf2YAHJ6SJ3ygMm4QO9eGK46o71Xv+Z3R
6KxV2giqlGGmIrX5fKcZjr5NVWNquL9+y4Cyo3lhHX1iDR3EqIVKuDTLIYVESg7P
3WlBvCchZTYWMjnWRjUUaguX5mE5a93H3Vn37XnDbNofITWxWAm9+ecOe5AHf+Bp
e+5TuGYYaoVwkjWIkZetw7TG8Pld+ezSCcwTIorAIkeDFvF2V9Z9Iv9gBiI8Gta5
oasYDtE564nWfDZsQFeXvh+liZyc2iU+U7toiJxx4rBveRn1wqv4zenQ6l/zJU1x
RSWvpzI89IZyGPeTp4v5tNi3EYuIFkaxeJGtnozVQgfygmWhpHdHQggs+zf1fU58
xYu5zEnNQQ4TmhD5dFkbnmgtyZkAOvqMxsvL5ozUlPzKxuZcUaxtZaRclY98tT5b
UfktjLh17W0WuDYKTzSD5GcV4vvfEscTrslG3WRqqLT0Ypxjh0ugG1uZBcbpn34x
4JqqnsfOezmyqD5KMujVXn7pFGZe5m+4Fe+cwumsYF1vxFj/7XKZZTaq1+ppoq77
I+Q7DPqUwlBbmPV9814q7O6amXjKQIjz1ehdn+g4D3+gms+Mu8wkln+u/nslnaLI
RBJqoIjQK/L3akTKHXzo6ybQRARnRZqAcTxPz37eB38H4Dv9hexKBoPWD1IKBO41
PuZYKnKh4zORJFizWrb6ELth6itrqDPwIXg3R7yJUKlGvIIxCKf39fkequPVXbV8
0r3fnW3Yme0dtOGpNO4j5IdRzAKxKE27KpeGrZ018HiDHrFjjAaMvFL5b9oXnhK+
sRaZMiadMERcWWHS2Hk19B2LDAI6B15+D120n8/sJs1gMrXslRXsxI9/7plGA1f5
TXdR+L2OF568GQhM/5Q/Ep42rz7N3VWnvTuBYDUIV5KHyT89GX9F75j15DqxIOow
qNWMbrBCnAQ3IMMS2BtySCaVL+W2WatPAg4MwaS2qh/3k+ZAy98yJview9cBrSVi
isjNrZWHq+5RiWwQrX5nPbGa/0y8wAMu1E0Vqh+rsdijHc1fSAwI2wMnJzJig02j
OIpTihstvkLwv/KD9cYxiGhCEALJrwnLNqarZHD7EOHcLIp5svhtacMSAyy5YFsr
aZcJ5pAIvvJB06uk8lAEyapzSw72gM+bTJIwQOJarppTncCm/+mcGtSO1GDjOuDZ
rcWmVYepbdytGINlgjMY8xVqIrHdLq0daXPmTO+sJVUmuniQR3LVj6zXCxFWbdI1
qiDRtROXY+cZ5DekQaI5cuV9WVM1JeaCad+f9g5oodulmqcRP9HZsYRTyihsr+Ur
Gm2kO1VRqWjGS2ELK2Vh+KcRfuZ5W176XKOxwEriPnI5Exnsql00ifklM5JrIyfX
4R0r7skck1f8/mvJeIi10H1w+C8IZaqej9BtyF/jBstRNvMO4vcxJJldE86sMK3O
whI5fqFkzjcyC+hqbtn7cmLIKWDNsbFJQbx4hDyjwG43lFvbeEck8DsI7ZkFZaLy
GRUmj27isAzNRjj0kFDkJdT5pa1i212fCn+w847JM4/VIYMWCy4nrAwb1rAd88h4
PRLGRPNUF9Qi41Xfy3cJ3UGBgbTlIdn0FzqDKe84SIyFQ7UavCxakfYjfiT04IN3
venvdf1S8Txjr/+u5VQ+azeP5Hq/fz632v+YdmAZxMlaFbwbQI0UKklw4st1Dn6X
cfMYq97x6LwqDrd9cX0aDNoYh/7X5lqyY5u1zqhfWl9Nu6F3PO+1a+hbcNnGT8kP
6y9ZQ5BB96DwtBwAMar/inNZ0Wvc8FRtJbGczKk0tIVECpOrFjRJetKqMPAJGctJ
5XNjUKAbKO7bhFYGA6FFOqWRf6+F7QjnNsb703jzCU/GtX5jtIk1SZ6DE8gfhSCL
oc6YIMBB3NuG2nAERcrFOfeDUkZu0s/iDdEwHufV18R9zF+zxOVujqN/ppiPS3/e
Up62i0Gv2RTYlF6sEyKxW2IIqtTeB1efloSTDUshOCmvxZ/G5VSbpgOMgFy/gAjq
ZSPfjtLLRQUS/2+Ej+z0w6qge1Wvg8/UBdWkmESNXhPG/8xGsExiXTekK2xeePKW
0rqKady6+fq5raEyb/hxql+EEe1wyVXhemSup6NLqsRLXtfqHb9xDzZT2faY9FNZ
xluSfdwJsl7NVQBKw7IYKt2ZHXheIsP5IpgtqNCuuRKL6UmtUalJUiB8SdtRZskP
3hr+Yn8IqrfuW7CAGN18xFHXYOcTSMgnzTFWXKq1V97323ZHtULnE1o/Aga4l2pf
VjBKTgNSLy7YCb3OQY3FSk3zGV+2EE9o2xmYQe+ni04t0k5vO11ubcJNx1jvhySd
XLh9V75GIH30rmypiSLNJxaJxEji6G7wBBfTMeLItraRe/CnKvzGv3mMat0cdmQc
V1y6iawMtYrIri09EuSrTyMvEP9c/1h/Y/bb+V3fdvU0Q2IcY/2VD7B/XwxWbYuu
a6aiMAdKxgf66/7O0HAnRwveLPpuKt4svfn5znYrZZbhhOjIIE8kHsNvjxefoUwV
3URI3KJ2RYqBrX+hKp07iUKDUz9Rg8s/AtYlUwsSu6GPMGBONnbatzp0AMUTl8Ue
KjT+X6B1kH5XgFEOO9a7RQb1+FIn/c6nzilFFnx0580GwekqRjmNRVWccfXkrwtn
88LiwqQ6hAwiNn3eDLZ8vRQru6vO1HOM52kQrZstEyV7M6m9Jo5Aqjx4tUKN05zh
HiCnjbkseIehsX1R/R77f5CfCvIeAAcLeAEu8YnFnDMR1k90pJ63O7SKAq5ktIw7
FKK2ynhP5DNfVonnOhZItBOnSMJFybcDX08Bx0dSfZUWI0nDB9blIBLfWAx5aR/w
+iREFtDos1th8pUj/9cr2Q6d7jAHNNG5N9g7awOxLue0i1fzF7UbmONhUI8sZROm
qEapivS8ivd7DWLWaeCUCEy6dQpr9qg9M1Qdlfh0U/7n4ytotqd5CJnAkA1k1nb9
IpEl93lpYkKzSJRYZ6IazNekvqt27+/IeCp0gotj3DK4NDxAOsaxODjp6LTAcgTJ
br5R/aBAdmL6ONC+tyoVIFV03ZRSK2JxWwEN6YMTUn5QgIbhu7pD0uEmREo4MfYm
3BeME9wzm9h/XbdvXQpiBw0N2FCsoKF7lMBZiqG450Osb22iFgzdLgD58nLfgFcw
ElE6Y/zyiaxf3AZlqTHObE0xr6gcNTC7k0fA9c0oO5jOmvw4n7bnTqztiODrsFFR
Cac+7CVnbPU4eXYIOfIDoygklhKr3qJVzXnRjwv6x/JQo6cRq38r8GCqqK15xDAC
+Yr0cg/00T+CZrgU+/DKL0GesG87U5dktzAu4ysfRTPmJEdaAfAb/PdyD0X4xhaw
eodL/F/PznHozRhqb7vAsVr+xuohdGOx49V7JqMJoILU3jH56lSt4FVh6xUsy+F6
MJaFXnEfKPDiGnWExlVkvtMN0gEP/JefaHAb1pkRR32lVxfIB7H7rRJo23hYcBzP
cVIi0v6MgsNf4m7Jptg1RxcyJJaRhVpbyUBh80ZfpYLpwK6WKWDZorLZspkcsOr2
INfxMFNLnHFk7mjUYx2Xz6GNpO0Cv1Mx1aYn9y+RYTsqtfYPK3js5zIbW135Uriv
8TFHclVIYMgn71ERiw2OhLBt1E8zKZETOmgw6w1zR+qgrd/Bqh9TYpqkWA6gYoeF
rzslMnIjnlfA2SPPqYXsLwkD68gx35ud4bwiCf7U8HhRDehK4TKCccSa24IxYsPo
+WdLUz+OsZ9SRKxuOSKx6b3bmJAEWFivgv8D/p2GXPhV3SrJfdDxuOz5+L5gGerc
UnL67CR8Xwp0mFVvGwrvE+KKWFtJfzJXRnKvuHnuL9Q+veqHt8vWyVaAStoZV8/8
XhTEgALADyZtZXIKqFhWRM61pM+OQpbhpGDvRznqiqTAH5ht/DKDmtekI5lZSOD3
UlrhY217oyRbZSGe2pg4S/0NudLZzgwcgZ4caRUw/U7dQaLL4a9dco2E7Z4ZBG7w
JZbdswCsUTW2kEtqCkdXAe8eNoyHooBVxdULJlIZ0DaUnKO4x1nBmxbqRSw23c5l
Q5gtamQV5qxHYZ86UGqGAeedeUdLTEOE3B0ue1oig26qtdib10B5ClrVYUDu5ZGW
0ZTouO/6lPTSqIQZQuTfVRfbWos4oVTxT+hMGdPzlaoXAkM+k9JJqBU8txVsQRlM
4Aa3O5V6z+urRE86VWM0vzBg56KNP+NMhWIFBtshA2tZRJvd6vh9YKnJGMjSqMAs
LhsTpF4r5jFVikghLKJEU0ih25qLAqXM9PmeUV/tNbC11JWRU8p25YMnaAuSJ6TV
JPH36LwigjKk4PM6cD+VOW+pCTQ2RtFy1oFdEmTJ4TUk/1LkRn5libPJVUZKNduM
RBcdQQr38N35KqqYwsdEiqRS1BYoORVbMm4VG/MaQcBgPCXRsDDhZ5RGUbYn+vf0
4K8CXFVfcRZQQpuJBlzbovHfO+Ru7snmka1jAaUvpaHWYF09rmiKc9cN0C02YBVZ
Z4FdAKLOqCIe0uDV/s3A0dUXzAzuO4yJQbG1G1pbcTiIUub1NKJZCL3XfF0jsvl5
2YxYnODxATdBRXmjMQow9cOe5pHTmsBYQduqSw5ltHv1tpC9yPgQW0vNYpa9vShG
AI1KPjE3ivO4xi6gho4LujKY2EWrpMJ83gykPaiP+j1MspUFsNY6VFl3GBySzKIG
AHu/u+yc4pbgEsYFwpO89vS8vPbjTy0AJpJX8FYpREk5wNxsQYRbWdrg5YV97bST
fnDYL5fxKeF2E+CHOwIyLJG55m+SQCLIJPzSHYGqtLYrNvlTClTMgMAfS8gmthVq
UcV1Q24Ana4IhVdvIPjN+vAq8C3F+4v/r9zNNZ2q402dn0ezMtJ12yVmAtcUCBhg
k72t5H4pgFjAnwN3vLdHOTD6JIg8ddGAV2CMNQscvczTtPMDvryysxMjHl+yuQqs
fECKjSngKFU5kXfHu/wr/YyGbQWCB2w8Ls+ucHuREolx5TcNB8IjVHuSpzClqqPn
ZlMIHFaXinyRM0Vs8+b6Ud8t9z3SL7M28i4i9escggJei8IdfJhbrzFf7/mcSX0M
/olxTkq/RdVyE1q2yoX9RoLkk2Ny7fYCdeHibwv9XwC8uJ4LMFJSu6ocod7SCSy6
7VVlTZcJ8GNzegXWRAdnLcU9zmZ2NE/x5sDPKbTQUYRng+kxvDg4PIAXWbvxZBbP
nnBV7zD8dnMoucgctFrYznLE8S6xW8nSKMZEU9NUKLiuLkUsyxFR/O8yfr5xm7H3
N8ACM8L/cZLalwvHqNMbl0nr/m4R6hKDIlaPb/ZNcOi83ivIcz44BMSsad83UbkU
tCPbSvJz559hYtL38Eeyhaf5CHzyv1W9ZleFNI0XaJZ1R4f6E8MTI/5yKwcGUlyF
Lvm55yb612epqFtZfg8Nlb9EvP2995jFf3Hai4qM4rjrXFZ9B7Ody2X5WTlrsYWy
Da2HJw6JfHZd82O047R4vvC61VyCOxX/WJQ58TYk4AsNjUKzX4UPQqut14xFx++o
sGX0HBOF8Kgj17bIO4xPohZsuVVFY3fUDpQmrpo0OhlWwGM2hER+W/ERJVwfC1aL
MOzRd98lP3vrKgs+uZYZP4OZaaOXBLPNXSJK1WeOIPPyDmK/NxJUFVy91jb/itUd
6zHP195FO0N/g4DLCLPjSkei0UtDO/HPmLVvnzdOp5QR4ppm1MmDW9IsKxAg48NZ
5MrPTDGHHUwOFpo+hHeJiJD7ubWM7b76R6pchYl202ZIqW7U56hooNwA3wkbKrr+
vTL7CFT8kODGtC3SVSA6PlX/rAu9j9BV+B1DFgPLca35sW0/a0jubP96cdyyVx9+
bAZ20hL4N35tJ1eoia1BVl1xNGIGa44gaQS1hQjk/O60gAjzwSRO6z72CR/NwQQL
OciE5fQh2bMCnaWnxqAO9CllSS8gmBEcKwGdAEPS3gAlfNKbhwvKGeCkx7DQlz3d
5Cq8Wiz8b13VynZbSiTkR7SWeNt4xWtiC/yenVACslhIXbZkIHM8syr16h3knd8k
SgRt1+ivluErOOsgkcmP3c5pskFyM1X7MQCjey1VYKMvdHfbtmhy/qE8B+narANe
CRPg3FnC3NJHDYPyT4zHSI9Hg/ugwWPdtBKTlyrtxuPLvQnQnn4Q0WcGCFwQ2wrW
ZWggo3lwV0ZBdCcLxWXt8skTsvEsxQpzyA99cQbPRTAGYZRihz8VZxAsLkmgWH4C
Go0XH4EhSJJ0Xcj3LbIUwmE9IDuvvHkIDS5TwQ9g/KsajVMyrfVI4VqxRpjTYYku
okrFE0eXdLf/YvmJibuGFCnUdDZO9tHgtBFRRKKR5bCZWpXMlqYFvtZoliFxSgmD
Nwvm57SgJAa9eS3kU0Qfl8B5Zm8k7fUHY99JVdszWXAcUA1DlR8DpVtvWB/WmCxU
VxEr6fhmzaLV/Vw2gQe+0NATHeYHCIW+sxdkZVaAy3BL7SEaj73WcQdYa7Fmd9aT
J7stx9I8rx9oAjFDhLTW2c+d+08QUL2ySwreE80lklMwCOXQdUb4fnveokZukGek
uoqE1kMSb0lbqB4iG0SRTMAgET527FbOYxyHrVfn9nEV2KjCv3B80Fufxp2OBY0R
38RJGMD4rB9dbqY80nfSD6bokXYlZYZvCDubSrlhcUBW+3tH2tf2YY9UZpNeQcFH
DEqSVGxGU9r06Y+YV5GayC68BQpjwL56Hsbf6PMStwTWcU9P2RZyos9KnWvbGe7y
NmH/pEuXo48GrA4bJsxNmm0WipQOlpr3BBwOH8iZIvy3rhGB2HbK2Z4wN/8FUtjO
+nSXgMAclFHMeE4W6JvsqQrsDSa479Be8Wc12KvF/rh2Nv5JvLlo/0rdoh0Hbdqq
Sks4o+4hSVyRPqn6/t6fezDRVo2b+7INhVNbyq+e+YREe/XmrgegqTfadglBuan7
z3UawP79//VQ6BZvcTuGLAJ5I2Y3hiekXuEBzM31Ek2opH7ldwLHTrJNr7fO5pTO
IKaJNF3kf87bbXdK6/iAFfIkN0tqDqrgcACAMTzKXf8226quSFvIDAgKYdJDf7ie
cWzKdNRf53BCAbGFkMqg9a1wbg6uEQocwaVXT0EVn1zrOuyiNJY+uVgkO+S70Pa1
iMH88jBIv7aDebfn8ICQRnIECiEMaSUadbK16YAfkZcPcf49pPWJyBKxjY0D4eg7
lEu9XVH+UvPx1pcVZ207Tv8MeyWqz05ZXYjfEE1i7X7UsloJEL7Yut34e36pR+mX
zqLRTgqOEiHiubkFf9ptWNTOlo6WhhLpMOeM/T3+otwLKxbxRjcCQ2+Ue+62LFkH
ZMYfjbAFA0mlOj8z3deJG3h5SMLdCNqrLKbV4YzD0GOqKdc5C+AdJLT/qdKg11Xx
yUobfT0gRo1U26anDFyCYa+54RvdbqhsvJcsJ+YpfUhpHahHZtFbOlIOJLyfEnVA
EaxHeiOdnqXdpV2z8HRQYHeqapkn3DdzYduDmhXG82L6wKyr9nFVW8nqSuy7fwMu
FURJZeo+WoS0UfoxAE00Cu+pEjbd44DETqU3v8YsZcN466wmRbnuFRcW0zpnX1g3
y+eEtdhbLx8yyz6h7g8znj+sGOL/dFyMo+Pl9E+V2JUX6njF4qcB4wpG1TBTNfxl
6U/R8HZMLi6a4PMsCEbbyCp8eI2D66iw0ZIXb9DhLzEfCyKVcFY5UVDl0Qf883Md
2vYVDkj+MVHgPBs6BfLUeKVruxtsjDkwB5RLrlSMACnqLFXn0rGG0wZwLbO5SOKg
a/FdLxuQ2XowKnPUWqr3/UUPMJoUROfmrCTpuZnPxWRlPU/aJ1um9UIQh7rwQog8
17dZHrNnZ/Af5bWSmiUef9Gl8Olz+2o3ZWnUvAZWhegQTq2ebFIv17Mj0LqTrbNU
KsAn5q1ZmR9hW4H9fuC1xzgggzqedSWIZ+ii6HnE+BApaFSWwUopLn6Fo7EwrP3a
YwRX4TFarMmZ2zyTQiGU7Poqt9wVbUhR1RzvMbGdrSSPEwtc9HmHeNvMZFXlSADY
rcs/7FQDFXp7HRHWVezclg/lpO2rtGAI/nxsoML9Qt0yGo03fM5/m+y1+TROWtz1
QzRrUCHpYiq/wTZfPM3xGCPLsH0ykBf3cShFBTYpv5+6iNiTz1KnZ3CMH5aYoDKx
njowwyHXhQp+NY0akFMB3U1v3A7IPVDFTqHsSrktAtDny42ow7zJqfNY9mhsy+eQ
fSbs0HFCLtEPhbiVWub0CXFs2ByRTNZLKcv/yqn0uGnrzgPBybPg3S1CgxOThNmV
lmqTw2XODYmqqPUKaAOa8SdS7lHdEiA4IX28wSf967NC9wF3WdDfmTi2vd4Cnffa
AqpmqY7Q+aKiMXRVWK2UXf7wZy4Dw87kHNRiOA5wHu1siaGS2kgbJWWVAXNKMpal
kPUPiVE6Qxs4g2nT2rtrxF5zjo+b22buTaqb1KmVs3XjmvSJH1apH+aQ7Xfwb/Ez
bBcPfGvJi4CzXajidiXmXIAHmmfs698Kc10FLVLlTEE0QHt6svkVueP/cTiFBx86
9lmME4whkq7c40ONs5j/h2HmgM7Yjz1bwx3i4BPbD9+KbLr9uSS40dkmIbkpXH5/
tUfWSiIfL2h3/nbKS37wxkdyplhZk31pqMEBdof9S5g3xKQXSqwYzC5M0+xUSQ6v
WtEfU0m/I5NtzAxjYrh3IhxXtW6enwpBxSn/wyQdUx3coJKmmHShicv0NimCEy7H
7vJDp1/eH5n5T0dp6iaqz48xH15hpa84VwM4DiU8XqKJe2smVCa39l3CaOeQa9TO
kE1s+lC4rDLlkE+c/YE8iIy5OnfAFww3WstpJkN73qWBnTMNPFPbW3nH1LyGDP02
8gwEwHmZoE9S8NeTWPzyugc+RwnxZYP7zpa9w007pSR87tPl5FzypoOLst/8D/ct
uLne1SjemDZB3vlThcAx1O8tiFsMXVK7odoeuU5IWfIGablCQF84Tvqe2Xesf+mc
Hca72P+wIoRwCyN97ZNq55/8n16sVUW+ZxwB0Tw3JW3Fd/52afIPzV4j1fqdosUp
F8xI7eQfrBUhWLK+cjqKq6TrYWuwt/097qx3ssSBweAUSOC0D1ygsc1r5+uH/3VV
fb8IL9WptZzndOm3bRd6UkjHFnwKVsEso4P5nWlTUMcU4j2jNqKadPLvH6ymKHJw
0uduzObvtw8F8JgyQHIphP41z9q6J1zk44zBk5XvqNyKLu64lijtj69hPoF5Cwfm
mltFhYtdE1CD9LWrdHYciJiCQtYfEf39SpboWkGhvPGPoifk7Eqi5Kp2qr9rJhN0
+uXTQmOzehcFW/HQuBIFVCpGdbCSFgvE8u0RRBugAgE9DIRtbhjT7JkuUh0Y57Fw
Vp5Ei11uUIoTc/QwlMdPtO28qx5x2uGN2639eP8KcI+pnE56Mgq8cI3tKHfjN0Mj
6TtymnFT2YSoIo2btaiVt42wjXQDJV8rLEMcaSiADcn98pAPWwqctVqg4PF2LPn9
VE0TXVr//66HtYLIcIYWWQmeGx0gvwc+35J2D1ijHGtBnNDLTusKLnMrQWTXOIfS
EHKgmr4jlqN00VOy+QvAMxRUH+Ipsp2QVTatyoQXPjT9J1dzuDZTzViGo0kD4LiI
Y2Yt7z13x2F+wugZ0kLylAsptjvMYBVZ/bGPzrJaRqDu22g0114+EKvVKOzwXHK2
fHCqCv8y1JvPAAxzKs9WRFd2QHhUacWqaA2Tu4p4Zzg6t8PjUpNa0Ux9HlAqwl8F
T9vy228GJFyIHR3uyJSGONirBEhc2BIs/bYILIc1xxEv89xC7zNKkwdwPqo4hS8J
LpyPNYW6RmWF/nv6NmwvkGYoNs3wiEsgH2e4vEZE5RsbJnlIVRy0BNiODse0Ld8m
XKyEIECFV5bO8/a1JBPQubQn5n4LZROiwyDMN1rwWksWRCXs2XWLUfswLt+ogquX
h/+4eHOIQBP9XjO0r8kOGwPmrbAm/o/R0li5TgDunk32/hn91HicvM7htCh6z4d6
6dagulCD6B4EMOtAY4xc+y+zDJn25hk6IycHHMaILnbwML/0TbK9spIjO3o2UbHS
3lTUreHGnho1L3laEAQao2kAjYM6RmnUFodkgtSqb1Cr3JYpI3iND7wAOn+VwWt1
IlOV2ZKOlDQgRbTbB7iVdedf8bb/4Aljc0Sl6sCGSSkZ6I/bVsnzbLlfPPxl8mQr
axWy2J+0mo19yRAPm4Q9mLJF3THCu7YyH/h8AjZeLbupXjt47k/Enjbo3Ha4rwbP
2A2X1OSVZ0n9ZpaBJUz1q6b1J8Mk3DitZ87JcKpoUEGMdG4cOb3z0f8qSbKW38dC
pLzIPBUfhxQWu1y1DSrhLeRxANFw5W3TGED8XDzLOV4ykjP3vlveJjzGJGA95MDd
OvZs8/sCr+Ov9lfThjh+FCPNon33yHy7TTfLTCFYBqaso2LMlHVYPGDwMNAxuFny
it3Lb62IUQbFVCXnTjLnXTgGdaW7XlfgKySsiDcVxVB6vJalUmrLHJ3z9cBuLkqK
lcRtYpv+Qd/YKTs5J7W4GwdNjm1FjHtJRjPnGO5b10sh4m4tXStN4Q+R+KAivFPt
UEZcHKSn2/aeYx4qC6RniHwOcVlZIibkz21l5gra+idViAVlykSKxTXDi7b/xEnw
+02d0ENYQlwlD23AkUMukmNE9sD7RrFL8iY8IWj6PdO9R7HYL4n2aQT+O24L2+sv
HdwynMaOKMIfpyVVaMkqHhbMFzxVrOExZfsV3MusH3kvTVVunR0dzSuaxCiv4yXU
jd9HCgfxD9VTrssSYDnoC7Zh425KPLr/V9iMWFgSY9WKFfGBpYt9VqtnpLktkbeh
Id3oCx7jSqTMBrrTJAZHTY80dzR5tASr70v9RZfR6yoH0zNe7O4pTzlZsHMAEfn4
lfd+wHM434GGKr7LktQVaksWfqzblfKyPiqvvH7KB3KrdwPUaUgxCfHxWA7Uouzy
Q9m0hTdJHc4QN/F+tvG+Uy3V0fdNJ/3c/g1yk9VEmjAXYq/mXtbCYv+nUq+0OvBt
wELBHOGh1QT1CRBH7PptFqOSbJ6mKkTG7AEuIHzihCLlVSd4WsRj0fARbeyGAeeJ
vuDYY7xPF/nVadFKmtu1W7qcvDte5kfIRsrJf2ZVRzk+qj5URFSvoq7F/FkvNrEC
zaiH0h0dngnUt2RAnFmklXCFBTBM2qlca58R15cc35AExfWyDSKz+M2ADd6tYIuO
II+4ovqZGvJ6qPrusa8VZfdPiyyrQCFnbrVTvsJMcKS9z3NnzG7FMEkO6BocEqs+
Qr+u4AS/8Mda7hoB/lWfJB2hhaBV/U7kyIId2JiIbbFvBik3re3Zy0dJnj3AlxDh
eCRewvlocVvO+lWCGo9jMJZtF2V7FHx6aDWRI/3TwXF8jD4G1RG9J/uu+UYGzkD8
oZvbKD0EpNtVfgu1HeQOWEcxgvLVyHF4dDVTrmTJtlZSezxjfLM9fEbkP3VxDgbm
GKKn4A5ak2hSlnLl1gumwZizjOGyBXci4n+QPpD8WslhzMYWCuwnSiLEJj1+XHWa
ixFlpnI1B7VNiooKhzWYbHooqXQlICHlyqNDV28wUFAN8Aip5GADhllw3MhaI8bV
dcRbnPv6JFxvokS5Z6u+Dqao36FmoLaQdx/6Ll6oIeVjb2GhP602RdbADsftAVxi
MX3r4vkOaz2yG6FpltiBAYVo1mpfioQEyg6iDbsUGyXEQRiE8BMTlZjE6QlWimev
+r2mSm0JcWiIhTXyXxe6s78l8M8ZmpxcjeC0a4A6Bo5edQ338+HTHLNOpaGt2ElF
vw4/MkPLuzNAQUl34rjGP5asgzgiTHg2l25qIE3+78dJ4KRdKZ/Mcs47zsklqMI8
Mmz8tkSYZAp7Qvwib+vCkZZGu1RVA8RYaJOxmVbnvJhuSnPBuYeASdiUA3XcjQ2g
0AR819QymktqTZPB6BNixczcJtgJwLCXO0/NHbip7XB3vdyosYFwCfl5tYpcdY7O
rerdivy914TDAUbW+lzHHV60872gtzoXbdgqHTS0mUcoO6RVQAfxMKrF0+XuWbmo
LAo6cdB0WUWeKfcdWjJYD4YfyEnbDb4RYT8kkXy2dLeLtABCSDTdX9YhvA0U8817
ay3vRhjO8GQEGCh20uEBv4dTNPiADNQrqVdNPsVsyO5kWi4Uew3qwqq75Vr4f/kD
aHq9xj+hVOikKrU73Z8CZjR7UcXrFpFVlsqbf5weO4jP5T4It9b0vTro/mfCEAt1
WcucmOrvwKIlsXUmztFGD2+KmpI8Dfm1KD2Ep2Hiy0jax5JpvmCrWuS29pvrw1jw
x6MwVBlgTKIUaYqPJgO39He3WwlSPf82CZivdm5+1rLZle006oXM6ixkCVqL3MX4
FNexGMaLwziM6G130PjpxaGDeTSg6sPDvFaVEozOVoLQLXjW+8B+2EGjcWYY4y6q
+x7RS0WHk6YmTNUa6VUp15594HkyVItyzLpQtkaBA1tt5ei8msrhSUkdFWffo23i
slJs2PQe6I2XbZn+r9DmgdwroeIAsqjeJej2wJLp7fflLpQaQswiBLMJEd72zDXN
l4JRmVMP6f1Vaz0vkEdNnEtHoyUZzQMHrpfzHKM3EEqNP5NE0j4IvyPOemIIIX1r
cIwMT5pDo3e1sO+qW4cFBbBpTF2CzoE+1pie1oQEWlyLwO/lSmuPlBmPEZfTQMdM
xIDgGNF2bYF7jxeu88EWog4jfkL3UzbGpyzBDGoyVku6En5w0FSzF2VGZBAvU3rA
4ceCP09SMDQeYCrvwunjvveE+BNP+nOgAcNec/ROSvZpNoM7NwYQtWAnTvCHGtfS
wnTyQLx0iTwuqnmVRArkPAx9i290idTWEoI5L5qg4xs55W5jSy/92zp/8rTez4pT
NtRrNEmV3HmrzbBTUYzFTjemysrW+WDNO2IbrcN4vl6LjTvWuoXoOHJhi8FaTsu/
wjXLCe3PT6lsJBl+yWAkQZnv6uoAqyq/pZ67ifI1MhFEaAMkyqDEK3l7ja2pE0Gb
13cVojFhqUA1/VTRJ4VQk+GTfiOeVmArLK4Iy0TAk+bq35YtA8zYuS7AVEK6M0L4
UambDvopuuJckZU3nuPVuvDRcZpBqaDvLLuyapbRlVOhzR/2jsKWS2UwMzerTMMh
yp8XiNhowjgODGThYJNFmTbrJRZAt34HBTnBxqJir6qVwTtc2DRD70SUQ2twhMDD
BSJVcg/9ps2sX8N5fXspmshRVtDGn/qrq8MWGyxdrG7EF5bY2fSiP/IsDMeeUU3o
+Y18AROCLgJF+27rSAZHeh5Q8DxQpgYgqLYcVJ6cRTdp4MRljW33/A84Yb7ahxaK
Mrn9DnXP9O1UWeNPXLZCNj9prK13zJdqLFSsm/Cn+/oqT09aR0oyNnV2OYxU6ca6
SAK0LDuv6QJvfawu+XbxyxaKllajih0bgot/B8bK4AXIjC2IvnGQ8Iki2Ky5WODa
UdiqC7dnmeiwHvZiYorHESzLEy1MaL6TVA3WJ+Ea16rZZgkcON3Gy4BoCUUpjJXP
T7Qftg4IH1/OBylVQhfBaCqNl4AGiM9T+8OXFPsWQdd5biYJciInHiKlGG/g2FSj
ecB/nFTbZGujdTrCXsCFFRzSkkPCjJKgYL3Z12ebbYW9xaoYoEPpod7KlDQbqTcM
psraOHQzscdQ9OsrQuyECQizaAmTL5JjcRLv6MH72T8UU7sbhPJUrOXlttcgL4W4
8VdUksHE43zbBxwZv97xGU9rUble6ZQYG4DN5O5dd2b/qXt4eeIUZDXY0c+5BTkY
PQzDu3zaG41tdUueFxoWYWqPTYnjdsfy5rZQP2q500+PDtp4Z5PD1S28grIGfB2i
j0pQlKQIiaM5SUGtbWOY8VGNVlLyy93JSvczU9diSFXRNai/s9pRO7FFhFrqKLFI
YrhWiv8Ax/LQsLNormLMEdlwAkjhy1HjXylZOEiYqdQZVfD1umYpNd0JMlblWESj
u8mNdFCfEHMnFojd7iQ2Y5B/b7KNQfWy/0djzUuyi5SQzH+oVO8Zk9iqTF58moj1
+PIPTdHpqnGIWtrGouD2mVgOv1YO9qNo6Ew8i0XtaxbtvVPTId52yuQQZ9TpADwu
N9hk+3nVAWPAMIHLZTDfpkeHezh3DiVb/dOrPN9yHl2GBwdYdVDavbdHJElEiyYm
9LWaS1/x6QTMdh+2bVSJTsxAmULdiCXnMJ6QEWmsX69aCp3fGPCAQmOW0PvgggiZ
6jU4JdYZQTlHI/pbDjiHLoihIt3AzAxmfHwg+i21e7Zi1nSJZvZ+FklX+GCCLCDc
kKmnbgd0GAxf3v5N6+kZFXntM8N75d134QzpGfEDvqqJM6TpYiw79Lz+vpl+IXpj
Q/CDq4oowPhCkjhXbzlwHLq8jhu+A8MMviRA7PltyAIsMKYcvzTm891rw8gOZqOI
J8XHajel/ruug5qUzsZQP1OW3Vmy7MYM3rSA1e5ANvDtVlMFONjqQ1D9ghrgEVra
icChDBcw2s8sMKcTvqkQ1KsYbd0aadjtlxXKaTQYGfTPgFM4xqjwDTrY6mIqEasT
7rz2tQMkEXnhH6icD8Js+FAcgHEdr0mS/HZqY1UKaCqRIIcMxzXFoU+vU0OcUYxM
y1KG/e/IxxVWis/E9w1835OFDlNUqeCW+lx5nlmcOCsMeqNvMxfJkOVkpwpxgDrP
yb6lHRoCtyCwHmhAkqIE/0y96hVD+pZN/E1OmL7V5+1Ove18/yemBM3WmWPxR3hV
SkQVkhMAJEG3LUjtbScr/ZthnGOc14ULynQmdv1pxNCShI6b396VJufd3fhs2cqD
M7lFwl4QMjO4Rigrx44iER6zeT75TaLdW0s0epfapGuJTLdKXytzcZYarLxDfHdi
NFvEgdun7sY7vxgb1+x79/jnSZwq9xBPDgLbFIKmpCRu8RzDK6Zs+ny6l/bVZd3a
Jzstnk8RaN4IVDthnvXcDqQk7iuDFYiqUfBj4dQgcb59r4XGQxiAgTwp+VyFnwDG
J5VOy9k/8dUPA826jf//jQBTRadRCh4Yjl6xk0Fyf45dB5Lf5j50xJwnlrTyUoKF
vzzy+dNAniMs3noeNHSI+75igbGYwxEt9UhrF9oOWuTvkOadxwBiNmiMyr094wl2
ZuMap7hSXu2KNaZBRq+8FUte4j9VzvH+2TsQgns/ugnD1x9lqComXHpJ5ylFzDZC
0fxiu0vSaZJUhF9k92K8zbQzMQeFEx1y9DlGK0p7YDnKI1pG0UEOqvFPpTtdyJXK
2nz/xJnnSzSJeu4mbjLpLX3nvFhW+5oSGVNo1JwsSHIw2/zTf8MktKGj2ShvpKpY
OtAITs81ZBtuGQ7bGKRzozP6QaYAiZnh6qvBQzzeoVSzeBAkDcaJFtZsEPWFBkOl
GGcMNRjeLLXCPNSARQ9yIhTWchlTMQlDIHP/VDjiER+UNFrwEbr/82zZnQ83wfJj
XB5zWN2GUgSrr8L6HLVkM6zWL1c1u4OHPB1aVCBcU5zkL2K4tAme76k+S2hk57Yp
WQtLml4KOwUj4WSAPVfLUST4/jv5v6K2JYlDiut9xMHxHm17N/nYGSxfAyaH23gR
v4bymhI+XrHS/5D2AYMW8BWD1mi+KWcArEnUFtsGlWJC3Inf5d0KxOm0L6eqnjMS
Xb74T+S0FU5hNVj83DtUXNifGACiwNPbZSyaYGySvfvL216gLyWUbdsx9rEVXzbq
OFuOPTB3cAryRzsHHLN7W4htQbRV9E0Sw+lpDJJ+Q4fRtvq2drGhq8d+0nRMsJuX
P07aW43T2GFOD+uaC/MiztFmLcSExp9MuWQInRtCOiQRR90jQ+cEpggZ9Ch1k0Y6
vyeoyMW2Utk5wE/NNopBNZRb3TMQ5fMgDNiOark6FcsDyogK3DvxT9A+Cb4jtv5T
urL5HHzCXBRA+R8jNTYIKfY4yKq3ZzSbM9IjAR4NGykRvsp0d9XkDi35m3zFG2zu
fddf1fUjnnnhO5JhQNd/SbLFtjIxpetlLzhnsEhyBq7MmnCWBtoeJxanHWv01vvg
D88svm4lyKeirJTzQHP1gvu43O2ipblXk/RCVLNYmRhl0/eQ+4lxPshEtoZ13yJG
0SGkZcFRUT6nPalsHHlcYRZrkD7yXfBQsea05tsLKyBzlle6mPeobzFhmae2IZt2
ftNpgQPLynPItEJc6FXzb2D0uILWDqbs2411xEX/GBQxAHQJdCMDG+KdNaz+1auL
ZJulMC49Xu0hiGCQVE7Q16mtswyooJdVJR5eZOFSYUg7QfTNuS6otLF+gwM9aLcR
lU6fsV1h9kx9epEEOUCivn/2huaqs8T5TPZ5HcNw8y/8iL8nC4lWFS8yb+Ymrxf9
zlql76EeWePBIOF/p/FrV7yv5UUWqkunFBDuRMrlRLznxd0T7sLZRHAguvfgVkm2
cEtziNFgojM9lrE0SBC5797v3HQiKQnUSUk1SSaSwucJjtGWZkfW/kVcYKo8zw6+
Fi+0rnhUT9oPwk7wBVyyJ80FtZbtXrxkJMw/rBEWd51nppYqqKQrQ8sXrcQbYr9y
qvaIdmyv9E/er4tG3NbRFhRgQGexlr6wPvs4phj8504Lrc7GjteQznSqTdFZW0pO
MX77HL+imHtQSFqI7yK6aFnnR3yXxDEHoJ5wJFum6UJT/nP7cNjZjk/I1lwNv20b
upTXNvlEaIYaSbjzQxITqLrPUQZHIbJDdx8Re45NZoogdgAjLKkDsoUjLwUPGYy/
+s5yzqOtWKAXaHdU0zrZAVFT6sgSPCVlE0Yo0UJg4S5mX/Q1ACKcbZQ62AE7cVx3
tRHzWTUYs2ClIWos60F1wYulX6H3WAHf3bCmlKvT1tAJbo/neuAztUPAbNSKDBs+
csLYVRHnQ1z81HmMSp/w+jaPXgeKjI2F1ssVDSX2wmtNFGf64I/Yb+SLHyzltQiR
FOQG0kR9wkwhm/wlTEKsspZWLoYBXWjl6k2cY+if5ioKBonLbSL8fZqQcmFZHeeD
AguOGA82/XrezXnp252x8ygKOdgjLJHwf+UvEDC3BrI5rUfRRgbrmXQMJ/9Flk8V
Lo3Tw/kTU/wSeVNslRI5jf1s6Jg9iEpfBAXRU6dY26HPgQ5GeEWiq64BgS77G3GY
MW8yaHnVvSpCXn8qD9xCRQCvCmO2vA3j3fUNnCUvQZIqsL3HW4PVRFwnKpiFbb7/
b8CQDZbJ+hon2NO97ub0QIuL0YAololehQCNIda/Bk5kDAikUYUdIdxIUWdUaa2l
34FJ3jFkJVsk/agfRn1aMdcthqWL0Og/SpflbZ7YA7HmsxrrDisOlz6to7AkjZHq
PeVOioR6wVyflsTb0pYpKIRwk2k9lAcinq/4IRoTmlFmI75s4zXEMdy3cugzexCb
4qi5T3X28k/psochJSxim7/cTgS1H3qdmyt0A9kw7i4XeI23UsEkzgaLcxFzQ67y
HndFHBsMzNkWUUOh0myWi+QIuQl0bRG+kxv4fh6wfQiGjSAsdKw5fcbb+jNe3NJ+
WEYNhVjsCbZwgDMoO9/3qfEXmPmvXKRd8WFYMkLpzigB2qwdp76PRoERlYv/k46j
1VrzZfdEbilVRqFCZuJeKEw7tnNnyP+fhwu3q2pYh5IyPgFtH9DiyNSKGZr7id+l
VfOMWYNZqEs8EV7nfPrkRWBXGkIW4QM7SjRcB2718cCEP+Zxvy24XjXH8ZoYAtQj
1HI+oeHTMaoJG3cUsEMHKvhO722RlDFy7gnnehA3PFQ65stVaKCZCO4TYIKy08X9
XXO8+MKH1UKs3bQfBaX7awF2cJu5x8A3VaM+rsOEEu7M1vEtqiA9bSylIKLPWmYM
HW2hdSN7AumEd/ElHto4DH1rCejkjfZM1TXg3FlYoxQnLyYZ8qayl9dO2b3mT3kf
dRAh88j9egb8yczbzERDnKPa+KXOG2UPnrujCRti+tVk+wzFu11YkqvyfKfLJgU0
wcRTY5TpuJrcQPlejSY+8z8O4Shle64jhn0jOdi2sz6nD/F5yAEz7yByVt3xYIg1
p8T1xsRdsnk7mgeAwcY0ICfE3ls3Bj/nEdLfrEhW02pYlUgeNSOq+ZYZg5lCCQDu
ChjCWJVFI1v1NIFqHzi9q12uTmHuFsHGeF27F0yCdcYUVJwt+yjbKnm5TbFapr4C
kiN/GLAYJ3i/2YTigNl8e1kLZeodRzc0Kp9wft24mFGwgUYOPg2kg2Ev6kx3Ldnq
wj2+xM/uQqOCzZJHB1lLzV5WY84V08iS/WFfQUh/2uqpWIoi+jCSJtvjpD9DLZlI
aUduKqoR0sKFfvncP08KFMyq3HcDelVwo0GcNUWthz8ye+HRSG26KRr49faUM3Yt
+3vlw1E8noeCBQpwT8zNr09pMs/kxAv3SObZOcd9JfUtSBGHsuA7WNdRGBUgpr/0
nZ7a+6vPnr6MP7TCPcFN5iA09QMcNZ9hBHyRXH6j5cE4M/cOO896iSFWseqfgs9R
d4woEnMDqXNhotCWxX0xT7E2d34Asb35OdynqD1Ff30ycipi0wIdrKP9lwsHeuSM
2EG7lDau6NO8Di7dKqJEbO8KM/PwWA4aKVcYuY1ceqOtSc97x7nxFKZmVsHFQ+2s
WI843jkad3Sxiq4pE2pTNjghJpbGf33Ua2TMn7XRLYNUvcuUZ9oNWC+CDbTNJtcM
g73OIsX8xTUBhDepIXrp8oSPo3I+LPeLRGOB6OwX5jvUxroje6akqT+pDLAabq7a
PeAvfo7BLBzKBg+VQEuM4YWj9/OHBZGBAf0wEiPKdk/QbiBFbMtXPxuiloVYhZkm
Siihquc9iXIpNoBZRZy/WA+fD9zn15y6DygIEM9bNin5Wkrtmmnsjz/7tEWZhTTu
GS7xuv4SET57FYSkK9TjhyzKC9uPNVHyAKNRVmSgEERrAYS5k53ovPBF1CLnyS5B
K248RsVVwL0UIDuYGQrLXwOqyaWOTzpI3rfSQhD5gjt/rsLeqhNAvowj1BqaXTuI
R0SKG2ZVBSD1g6OIhnGmuyo5IZsZEtoMWExLwVXiK/kOLZdj9E2VAY5SOQOXLiiX
mLfUtqxKhdQwl0DDRxuQGOPCPKJ0m30/tdmAMT+zvs1O7MrCeGNFNEl/5CACnyt6
Vs1oWvmEhi0zI4sqWCI0u+gYl69GKdZBV5v/k2SIparzNNH1ZXY414so0yBDu8D0
V2x8NNfFa42LhbMXVcnnO3iRx8ZQkvXmdjf7wZVppgUkYClqlUrjGRxtJUzOR7OK
4PSrWvUtLlhfyJKQ0lVO+GlnNowWqoOyGagJi2MnbQKPz/macRvUhEM+WDDbIxlc
WQJkgFEehotftSJo8Nxh0kcFyx9mn/HFgHTsUM/Ni/B+e/InxH8Vi2SSjELsf2BU
Ymcz1Q5MWhYeAxaZR0c9ns58iyXGE0TiMLW4UW9IX8mo+CiYoTTBPyYH4W2IRDc8
yB2j++Hr7UTONdCwsrBUVD8ifzL6HYHxmSShAM575DGlqVy9t7hfQ1AXtS9hq4m4
vtY3j8k08uccLiX0iYw7D8DZIulVBI5ONb5oWVGt7e1fxAXSfMj/+8JdMFWQ1oRS
WnIQ8LNoSmm2R1B2oKbyhf7KDXwVLJY1/f/nzYiAO1AOzR/B0wy28ZhL1UGeJDM3
ahCfqsd7IZAnmlemdEriQZZv9O/W46NjDt17fCsUUI/2NQC2mcHuYewnTiPtNKNl
ef9Ssm+CvSGyCz5arfvUYcQmk2BrvpR/pKMGFxNXPE1NIdgYNAAIa1h+aeKX5GYs
jcRt2zAV7kZdpkIF4lg/rncITfmLI5zVZR9WMGNazmiRDvg4xpTcrc+4xDPDBVIm
SngDCJgqMsQIJ4cr1tA9G+mZoeVTHt9VnrgYDlK3woDd6i1pIe85n/d7Ya+cxl7/
qrhTqHULAbUaS3nWtbNQEJXCFwIr0Ty/xZLOV0eafIEgNtLpc1QKXCo4f3L5VUZI
VLMe+dBFiIiMw5qc6ut/+70Mm0+BjhdLKggOaX4DGnWiv7K8fl/57GThMmdo5aX9
ljS+u3JKp16F854yVq24uPflwHws2NrZZYOfDuXciJAxpfWvmtmXN8JSwAJcCpI8
rvaROViu3dOiVzwV7ssPJxRgow/WojxvhNoHvVPjbHhjjUfWFUx0n7QqBM1AOZ93
i0IUGyh5A1OBDktF47FT8fGqPONTkKBC14DQO7rRaeD5XQKMRkb4Xs16jGw5ZjFC
kDmGHCwg/YtB0quBfDimiEwPG6+ccYFMQ2tJTJ784KrgOKcJM2S/9ch4vrgKppGw
4zyrx0tZFLAo30reBPXGGx5VWlEQMcVaStWuLRgzIkH4BV6ve9WQ5Uzez8X+lb+v
m+3cppgtTA9eRxYz9oKUl1rZb06Vs+my8XaBoJ0J7oE+2zNCfSclsALpLcmVwNz6
1GCzIXgOgrzzvHBjGLE0GnnWuY0516PmzAFrpG/rSv6p6ykBAbugpTuW04DoFlJZ
8M9OKxoOEFvhBGnUkAv0FG4Kip0yIsZvmgINr1JuMXtF7pgZ0rdgDt4tl0RaIaeM
K0hSpi2d2ci1af/lVFnoxMMYy2bgcAdMfACGiUhwmUOTOT4myvouh179xG0d9Y7d
BtqvyqDtZMNBq5veaw3abospWuOArNRE7WxGd7zEz4wYQKW1UDcn8fxblM7KfUiS
BZBLfNBbqJ8YhInkJzN7Ip5aQnk0eyrHzJVcifC4JJ2Gb/utU9tSf+PAUhjzpe9g
GGMoU5tfdAkbiOj1qhw9G+TbyrZT2HcAcOYn+2kJ1pA1b95RMAhwawhcxRxU6hgU
7sVsW2LdDnwMmU58Z6FrVZaJeK0Ucq5hgWJqJQ0XoJ2gvDIs5rAVvoE0+OpLUHhx
S4/qb3sk3+/Puhgop5/MsQbpubYv5CM68qBZPVeA2vDlI2WuX/zm09TjfmLsBRNJ
eONFyCBOEpX8AeNzGxWfkG21a3pNTnB6VldZ1mAyocGUVWI76nsUGUwwFzP6W0lx
ROUR+2d8DJXC+LEinozmqAem9CLND5D2yDDRadQ73xglLzWmjdzi3lNl0S1CxC1P
1EC9Ge1SIgzI8vddlcBbxQQQis0CpnKlXdHIycPzCdHc92T6Cg4hzwgdT0gadAI3
IhoBNbvzeE0Ew64l62W4IW63DMS615NHvNPINFgzhDl+Z3OiWzFdoZoi6so3EAme
XaxwIhOA9zRt1ECGd+oqjiHpoi0gBsaZxepn0NzBV6Vk2wWwvBSS3XQqIiItbtZ1
SqH3+NAkeS31F/mo7GRkUT3sUdbUeBJhHzROphVR3QPxcxkGStxSKIm/qIgTezwt
20HHpnUmzbwZyIw590kV6OQV8m3uDE46P0Tcw6RUYUXvwjLzUg5Oxr874CKjc8xe
kxyO+9KFVSiednuZTz7gQWmf2yOUgKY+JqWnxKaa+9iX6TrmY8nI5EWnU3nx2NuI
+AQ2t5UiDqvpKrYhn5HZT13/yHXtqf1JhbZa2TQ95jDDoKehb4fTkjb8/ZIo3G1W
1RWN6Y1+XyDat92sxVgcr/WXNukERuSd/RMkSpeZpbwiSGbAH6cLBQVHMLiHn3Q7
pxcsyrgJn++yPcLimVGYOkKqQcxplwUi7B/MQPmIL6yuuEuiVrqn+BMlbhuVJG5k
w11vg/wckrk0ulfWSbLWZxVQRQZLkgZFZDRPlFyLz6wmR7t7DwYcpCarju9iUX3t
CzvWKnNBjloBgady/3nyr0x/bwIN71Uejylax1V+eUzULIGDct9cvtjrEx9ztn7K
pLbx7+aDZnjo/rknMCE0y3wqioBHwb5HzI3kGbfr+H4cc+8qgoYK6wsNRjMoUPE/
3DlcQ2jIPoDE2estwuiPIm3VFhpdbJx8AUt/fZEOCc7367GE2JjyL3HO8hmh/eSr
YODnyyfRCgxuNyYjwR6F9y83xqODCnWmPL2kapxQ6i6HEY/Fm7FeUH/WcW86pRBJ
PChyAsaOuBf+jr4smuwhMISlw8iEdpzdwzu+HMIIQoERSWXL7RUctySPL3FA/t9r
9MHundvrhGOMQE8Gm1M7FdQfDfrRdGCuDr25Rtumc/EnDDUCW6MmDClYKvtXfm6q
M7n3W61fqvh9Mxr0p/i9SUHaD3+MNG24kBhrvS6llnwwAh37FIpop49Ab1SbpumX
E0U/bj2WvD8BxHff40eEOdTcUelvNo/qEr9jFfRHJPvmtZsPsYDJBWawTaNfsCsc
/kG56ZEYMPCbCXjPu5AlEmtunU5Uchf4LMTwUcBgYonoMxQEfxkoza/xUnFtUPkK
ttGOPWAkcq6D3KFYGcvj4X8JiyBDMhDV6jXKR0CFHB13kVh9tkGJrlDHowkfmeF8
xV/8+ZkwnJoU4jkgahn9EhZDHf79f62Rzizn71SvgKYih+MdnDdrV+UrqDTDk20f
ne6gXXNCZwwzzn9NcPHQV6cs4wynWtO131USr8FLQGlLiMbqSJIywxNDuCoZkZIm
gsTSM7d6QMWQaIxpDQ/ISqS9Z8jyX4Dr3tQC9VnV1P6GDmdS4ozSKLei0kFpT18l
lRH94VBEGApnwym8gHnmfT7+fevwT8HLb46w7j5EOCv5Q4jOIRdHLDkLbai3oaGX
4tEFDYtiq3cnQ9LWgevm0P2b7X8P7JQCyEwp1TDPPiG8HJZWpr8EIAfxcZVXUuun
VkNrlR1s+lhq/Do2QTuLjaK7xlDw5mVpCjgOrzI3Lgw/Q7JlDPa3hqr9TweFloAa
wduSBbmynsTW0dcc6wqizls28ITW+llkFphtPDAysVPjqcizU7n7jqP5gU0zPjW9
AO+NpMfzzxZi+MKMkJvY5poOHUx9Qz+R3Jul+C1t8mTKz1pvfkVCIjAC+Cd1NVqT
rjbCqUpf50uamshTQrLQcU23mR+NHVeKkLQx7/yeNh6Qc2MFxBIbywFOh3r35m+L
on0VIRmUJ4JjK88c467q6S9xLrWJxYnkimuI0NQ89mxR4jtlTMGD3/bPHgPUHyTO
7hxL7bDlc+SeRIEnEGHW7iePOD5K7Mf3HIu/2FHJrIP29/j+7c8JSDnS0NmwqU8A
BHK7/6fEY4IzGg8dAO8OCiK8JsASDBezxJNa9q26tb3Ce/2s1MeUwfB52WHR1CJW
TJuRV98ZwGupnEMXp1vslBYfLuId9a6zP4MePUEoScAdDOKDyudzWsrwMsFNLYWl
8IbS5s3t6IClrzgW/k59KmbNd+sDpH4CSqx3D4OGaSV22rJfZUl1hHvqZqYDvGRq
vvqkOyRLiFt+43UmdDZJSDKN97vnAbM+K0J7pvCXvYG3F7f4JPrPRjCmqAEjp5rP
Lt23OzNs5rf2/HURsZnHN8LW1JC4w7gtRHYIFCnnqjLr0U5zl84sJpWsdhotffdC
4mVpl+bavi2Dsxxk1kDvFox38aBKfeKLKo5gctIEyIQykiy1X0MxbgWR4mA3AY5y
c6QhLxZnPFStrP4isp5MYI8VNKXIOvJx3aztZy1Hi9XtfALttVuhEprbj3kGkDv7
hiHYBUaHzxjqhlliNoYHP91It/MfiLp2jDYSmgab8xkq1M67tr8nmbmAUGuBPU0X
mBE4wERhSgdwI2zyjiQ62CSSyWLTtBaDZCWtRT2fZS0ZR6gYyxZ+qWNg9qJ28h4x
Dl7PDg7b+HY0MqSQQfz0BgH4yYfrGsnTD/67ixKGpD0ZJl5O+bDn/hS66fzLaLQ+
O5vqhYRb9cC8XENq4w799jz9x0huOzev3d1/TgKPDjfweXnqyrJo1o4014sH9hUV
DiymIbWqElg/FfaQJrTQX4Ovm+UYOcccMuI3bYJUy1t90QERdmQokMFHQLLDd/SH
aig9cbYZv2WqKk5dg31qhvh9EgEOcLvDiPC5xqeadry11BNLS01icyHi+ajARB1+
Mtf2qQyN1tTaDlH7DQ2cSH6PBFgaESzt4ODa13joXNtRlMVOfb41oLTlSXtp5AwI
/xirDfDUu1/onTX5AAi7GLzfm0XqBzg24ymclQM2J5bIv6y+5Mw9kwVj5oUWQddZ
ydmuMUZpTa0vXe2iKhJzpj4QIjq7dvLQGAjOiYYg6n5kQO/aKc2NSY6uscQ9GmuW
Ril6htEDF2kdq1U1iNP/yhyH+4H8m7Uw9Lr7ClAGoB9gwCRZTTOx00HGyAH2Ci5K
Tp4zjeFvytni1Vw1YyIejZktsONUtzNnddMISvOnKh62RdW3RrkrgaygP+hbynrb
AfoHQOINKhcDUzhm3U42pM1gaBLvIyq+wLASSbIxlgxaMqdE1AFGJ44zsJQ3P4is
u2bli4tRfZzVFDmJi0tz84EShtISkvOcVTY4Ij8Vdt45xi4Kai463FM+UBFp/nbw
+VsqZTikXeOSFQbVKGX+vDMy4O/NY3Orv90uaySXuGVrL6eXUp+SNJp7eS95pFvM
49ZbNAXTR7X5sVX2Twt7Tt7OJi5QuPde7ikE19+jv5qgM0J/ZVVIMH9A1VeynoEp
+puWKCS0otaNlpj/TBb4qW4VfKhdf8ZlRBNbayOm4kzeWIPhq+aRjxfQZcydXI0S
TTdJgcHQZZ3tXpMGxKc5QnHY+8ykolexjWdO5VK+8QFgEA7kAHBXKJZV6P32aG06
sIRvTAjXCixLMJGl70zN84tumSXnd05iaPYHI6iWkrZbTu4QLXFXiROj7OnIkH9S
aX4wfibfPkVZPkHfDnTDQ8stMxCxF0yEyTiFBIggjSYd1Ytp7iFW4vZdVTd9+XvM
L7oDhVjTLvGXM9BAtx/i7dWZBg7g3Jb0hO8kgZttXxZf/Zw3zbGlB1X3juaGwYto
Etl6GXvQhxdFq/+UsX3hYe0O1ETu0aiYQHpwaT5m9K0Z2yZkXPbfaRY7bURTTvp6
h+vZ5ob+dnBwHdjxNgicUbgRoNWY3ejkq/GqNkl4p9VoLdOLcA9VHbvJjXw0vseh
bNzvxhx6p4IDGHVYvJ+Az8IdJ6FXMuUc79Rjdp4O4M7JaCaMXnKVRbssFaT1dHqN
juRsCS/JloZk1suWmYvJCE+hmbTW5UMqOnzLWLCNEai5jBIdkFp8PzggHHlkEStz
/ge/PuqtPcT24MnTC37foKxvEstg11pg8PGlxNIkts8uwS4IzchAuvN1gb7fYEBW
+y+UhoFvWJJz2D0VmziT3z0z/WUfjWHl3MHQykRdBNtQfiGgR/K8OPHmqSYukhxR
bcHRdD9au1LzHaraAspkJdAWH8NXF2uyDOAt/yOS563V/CJx9awAPFXMHLh0KNN/
Tz+qKIhMg7P7U6BRGbvT1j0kyQ1MoDIWJJbr9DL7nHDE6wC0TSPqMzZ9fQcNED7I
wsOojFyWmUidx3hgRgnjPXVfafcauiMnM+ZAQH/ipUhDoB+zNP+lbVsW6hZUUvhW
iitsZ3+1ITiaxZUXsY7ERUOT/e8NibUuefMpZWZeH/E5zGMWWF7SRDTapgFMeXT0
aFn3i8yjln1JypTV2eEGsR4YlLlg5sUifj+N8mvTIMoWjoFf07j9jPfF36AGHQ+1
TZ6MmAmIZWQjYzsIoSiHloh8EnShB0SIrNEhENUlLLtw0JIiEKjNQLO23DakRrvU
Nq2FZc/It+ROpc1VmxHX3PcID26vDV5KKRwcpbXmCiuG8ZW01nmfUy4dI9HZIqC/
uxZ8fpBLjiDd7loz1DGuCvkoFUCNsrNaA1hX8kT40T01lTF/MT0MRiYd/GKwo6vd
k9zy+TK//M27MkFtuhwUwo9JzuFmkORuzx7ASxvztEhfXIItDCnZfgk1p1KkHRCO
VoDk5xDfdGmS5AGIl54FMPgWAjR/XW1SIC9LzdBpzAEbLpKNGtF0T/W6wE+dEFBy
M6TKWQjDpe9PUqt87LnD9aHnSLlhuYr0jJ+cRXNIuD9q2yUmqkIem04vR8u/0IGC
tYPSPhIVDj6d1ytAkWDOXAGXMAJrp18JdgnLYpzOW3n3qk6jlpAyjevdocXmOleu
3DzQFavyrroBrIorwIXkzIw4KrTamwWPdvhZd/9UN8D8AJj7hwmxby0BzPtOC+wY
bRUeyv2cA4iNSmd1rmzNYlMn2TO5jYULRe45gtnyzzQFueacO+0La2WWuOP88jPG
XJ03wo9vDD0Abk1BrmvgaNYs642Cjqfp4fr0cFuk0vyBdz8StEIq8P9d5j/EP4RM
nSLn1BN2JcDU16lDmb1PKnV8rO3MdpCRDirDyvEE6GdSIwh/SDGFeCDOqGI1unTH
uLOuLg4TgRVPmdewjWHds8uiS2gCIr8Ajp8VAWpiqc5Gyt+YNz7QfnpsGDluJFCk
m+ngc+D09JJBXVkQOI22iXOL3DkNmpDFazM7AWoI9IvZFvYpJR+snssjXNfX10Ur
XdMy3SN8LpPksUZGqlSW33YKHX88gpxnUFuTgVZkTSUm1TcBCy3vWdqfuMmc35di
CRfRHRrG3lDYwTb3T+KFtsvMJCnxVpnaHxhPwMstSQ+MldGmxfJMcGSyyssMxsyf
Cxgb/TY4kpOC1vi1RLLkryqYSe7dXhXqqMazKLyiP1e7Dk7EUHKNNjx7bQNwl+oe
W8hthDc7cr8jeHQATLd40v1kWHDucnQEzNzlSrngNraNxTE/+S0CXHZNfF0YEloZ
uHzUym2QYlU06VYunBC74qSoDWdHZP6O0i8VN6jbBKxi8zKB3seX+mNl3Awt0Qvx
TpFcNl1Q/mgtlxX0dNrja9ryK3zPc+MxogV3vbOpwISxDFg49ZQtzALHTHRmCh5C
/yL9TjRXg89RPk1NK2GQCs0F+hxIxVKa6/NUN838qnunPbHgDTW5yrivPt84G6qL
yyvkUobcuzMu4zjVnR6KaCq629nQYtEy2jDAh8VAjRt1qLwUHHyFGXHOoktQDpSQ
4Bt+e2lGKFu6PUetNWTBHLYdBtqJxq2p2DOztlFcjogLXZAe5rHZvKqzsu9pmLK8
2vjXdVuDohJCn1nh9kYH3DqzU3G1mhq3PWqQdOZPBhXmg7ReyhslfvB902Ss5lLq
BJcqOFBdk/wOtDMhXnWdQjvG3lZOz9kLabu4CLVfAc3xeHDLj/Jps1iBdTeGQjSV
Uc8joAL+H/K4i90p8WH2I0u71slai+keqFTATh/wdvFtJuJ+NoXPs2IZPQBkZB0K
yT+TCVgc0su+eaVkbIPMI9v7JyBTU1SHTuh5/EeZ8DANp9rDRsGB3cgrLWfpKQMq
piiMYWXk99PxjdwE5sUeN3n0p4vfAXwfrk7vrEJxFfB7vB1jGpcBF+1cjFYJ/TOC
MqvsMr8h8eH0ySf5XaN+qF3y9qCdgSZ4cyOajNxaUFPswT+j+R33mGx4+VaDvM2E
oV1Wz+4hcv0VawKJMPVEpDESEAO/NDFrhmQ+sEHjn/GDwRZXdIMjD3WDvgZICRHh
5+p/0SM6YkRfDwTlVR0efgFp0qKYFOTaYNV9R9fxBz2m8zY0am5ngCxn/HHzkbLk
NiJvw8SVMMHfsBs8xAdn2ORlhoLSviKfwjKL52uQPgZfOeW0MxQaTQVY6fVyc4CM
XCtWRX6fzqjA1hio71r1ce7pq367g4Fl4jTPLZjXgmVeIhw7/AeZXk5vosCQge9c
4uWeLqvHVenC2BEUVWT8mH57fpGzWiUctGLZWEylnNI9LBdt1c0z8A8GhDPXelRr
XI9Bt9b72PBaIZuPryXC8lzbsj7JxwUbl3GqmCtqcCrwR0UTdq+Bz6PtjlNch23W
oddGmoNPXC56nI1P1j5CdIekG7LzfVYKG0s4t9e6XLmy+JevHXKKBnAc2quopUnO
2KhVS9lfc4O6sR+/jrClZKdr7/eooVxoj15QoK8bVmOtJrT+ncQzxQ4rP2AWVkTC
cQW67IDP1gqHtHQOSNFNdahECHCH6MKp1blgB4cvVaChVkgdRTqq3VlNVAd21euK
OsFc5msJUuLjlNLvKAjWHT+QclMRz55E+HcJole1F6XVqG6czlTqTh6v3q2ptMjC
pZWtbtxzba29UOJ+iGAkHUgLmEsxTQZN9rmsSwDBYw6MRCGZ5lt//EOQNDy+8xfN
mPuJa6doIe8zVgYyWnH7K0Yt4qh9BaQvDc7LWFjROfaaZG+Btmxn3gL2QT+cOgNa
VlJQxL6ppeJJgQbsUb65f+QgDqyDE8CzoBRBZpCpWk3rrsWTlOwjeCek17QqLGjS
/f64zRZKY05OchATiyNrt727eaVrnDtkiNTaYyQRhLicMA2MUaEeZ0YO4oxFgZ/v
nF0lyRZGCCLcXXAUmiju1Hffd94KMI1VXwv7o3gKyk+qSOMWQr91M71VXLKt6Al3
t1TYbLd7qkj/R/DOBMNjIgx8e88PhyubocbLcvPJ+WQ+nenN7h7aoOl0MjLBAOyg
KNJkPfYUVRPcdhmV+SBrdPL9R18Pvi8yiGYgpUBzggibX7oedpdWxNir+D9ubhMH
u2XKoT4tXUrc/35h3PvRKTwFdfC+bnDpmkQ3hGSAWFRt9eF2uqpfPC0kpp/jqA0U
Hr3EK8w3Oct//70Uit5sDGFhvhBHj5pnipZpMhFr19/+Ag4/hFL2njqwH0b2kOmh
iQiJ7l8Rxa+SGFNYH7alKIto8zsmBV+8gPWMECYHtFj9cWWWjNWIlD7FY46UKS0y
gxnEWbcvVESn0eR6itWeE/wEq28JLYciaZcSMK7duCHGky/CG+QuV5GT6T8UDCks
qSzwE8iwoIf0+Xrk8yAnyaWpoSphGzt3fDicp5BvxY4Z+sF/t5gpPvMgA/91HMou
3AmrzZjhsnEsTRzzSYjuPPRwSlb7AqOtUxNWadb4MGBrFJvEBsD6i0a0DylROJzA
RcyMI4Tf/TrQIbiFqAPbmUIn4XFh0Ih7vGyv8OhPLEALnG06tA/Zlhuwqc0VJtoj
eNDQfPShpQwdv4cCLHS+3jbG2uo0eGeqeT2sOuAQpHFLhNR1UCG6pNkdFERT1vJO
PTElub1FggcWgpCozkW83oCyoUPp7KTY4NqVlk9pnItzZ1F4XGDljfwWiSa40SSm
p+XcYf0sAK3bpwgUMpufTEcvhiEnrKl+o2g+SrV1T26UfDyhO4qTGr57bqE84ggx
o0Emi08TzS2KOqORcWGd9drwK9TRDAU+KHfwRCo1o9cO6KksPaVeOKqv3m0En1ST
rZHLPphM7ckCHvvxtk5otB3HKNDb4iaXB6uQBpn0OD1dhgg/A7S5kLmTPuwXIQSp
/O6AzLNHdRTGzn3tMi+2px1s+5zzMhADnOsLjq6A9pYERjJgiGeBDwSOvDOa1LEK
Y8/eX6OQ0A7NBMWeSc28QRWu25kfvw4nhmU7h6B2WeoY7pohA9UUsvghm9PM/6NH
8SxqJ2DgmMvS5JMx26Q6w91PWFOAdOsdFOVwTED4wO2RasyUXHIbkcNh4NEgMKSc
6cho6mtE9RSD/jjt1f21iHO4fhujDSbmEDDfSXvm6Jq/vNpmHdR+6caLjA98y2Mf
L2yxejG0H+VdQDecpJoh1X85UiVap7kgtJveGd0gnVMTlpfAPA4b7BTYXIJpEW0Q
Ye1myO/M2l9kdvB3ntwL+mhWXwrgG7SwLM+yLZm6G6GLmdmzGnuPX2H8qv6TUcw/
xK03P/89vLgUUZYtgZ8XMjT4HPX/P3It7zNw4vDzzafr4oEGmM2fK8spoHlsnW2b
tVrg/DvdA0iEy6x78qXOy3WohkNpLN5AnvXaT12yvfQtVBkaWO2lFJWUOnIUfW7n
Hr/LXW2TAKKOnatXkm7NVFGJYNZWVU67nNS4jLQk+ABFo4Q6Oz24AiV8YsI2cw15
GxbsL6iHPvt8zzPyLKUKZF83gobsqG42Tn8+LEzfqZEyBQMYpVIUvUTQPo8/RnPo
G2R5q0BuGLxQApdVg+XDK/g2gEVKcCSMEGeg/B1eYRS86xCCBsK2HqRTpbMMDGi7
esj3xsLBs8nxCsRrqtq/mmCiF5kYeWl+q8oB4u14aoUm8zp+0txZ1SnDVPq0DI+g
DtgvRBMf7RYC0auz4gK1ei1maxYZabd2ekXin2s9P8gAOWWtnj5J6rck0i2N5zeE
V/qYmXrXwV+eSwEsBnM0XgeHJa+dgsPPqjogcUXS3Fj7YBcTlZEGT7/GBfiTSs+q
HuK5vPn4kWdHwT2KYTzm1AepjvRaJj+5WXuU3gFj1JeXz54laniklmrZFk+jLpYZ
UELVXxfq/iG5ue6dvhSOnK7zRBP+SvvUt5CBrB8v3KgDRPq739nfEjQ9pr0HeO7t
EVBGeZ4t75ErnvbGs98JLOdkd6L8396VHniVVAEE1gw3kBbDEznBPiwsC+LXBLxi
bNwENHr/MxGblsWCJJy+Ih22GquCbU06O83YqgKL4OK3q/3hOrkfmZxeE58bDbsx
zPJvB5tqe6WM9ShUHSYUCefEG/4Cvproi3UlZLViiOj1Pw+I6yqJGqdPw+j/QLOO
6PvilTD/8aTz8l21PNJHmjRGV5gKL6jaA15T93Z+L5VqZZAmf69jT3i+e/G+1Bv8
WDimE6AKq0Viw9Z9+7FGmFbqxEgEjJsB5A+7LtEUVzKiJ/NlX/a9YmKDXa4NAPDB
gBTOGLbI9Ekper7i1nffYmf3oZRpgFg7JkqFEdsDMrL8Lu3etJDQiPCf/yxKf411
1+S8bue+7Uvz6e33swjU9fDR3nUbLUhJHy4l5kgZ93T03yv+E7mppA9qdZ6nV/Ee
NnxP4FPclapEpT+qRAYkW77VRpcgZkIEsIh0vkki7vQKupelt3/BOBr6aKdRbXV0
EFWX0vvbCNZGPfo0tr4s+Em9ffI/+aGNCcFsScrw9+AsFyDipfV51npavGCmMdQ0
2cBdTj31QhfY2nnbm7cYg7tEiE+oKa/8IR0IrurpLzKbXfOvuikJjhJM1vl6AO3I
3F7fTQGkPgTJCSwfekM0j8CywYInSMLlahLiDbHYKukdBDJNkSx9rgtOF7vRJ+Sz
RiqpWVXfog+JHyFyReQqxpSgqNZ6U8PlxjJkcfoF9aEDIH9xL3RL+6Cwugq7x7AY
2eizXlDMkSwyy5eYlyImmKSRPJLuxRpRcXNCvA3utdybUsuxICnuIXu1PZdVf7NQ
8J9qRUDmX017HnJWJoPSfQKac9R3xIm2/pLvX/RPeUT0pj7DQW17ppGT1WDLQpAX
Anr40S8s/sLMDsY5D73xECxMYJ1FmB3YOzacfvf/9ZC+4dSN881fnxzSxQL5ag80
q/r1kbXy4/v/tIQI00vcjUexTByzMd/Ly+NyHPGDeHxYb9CqdLaqYHWDeJfAaEUb
epQ8uORfrftH8paxccpjaLFvJwBgWv+bDp+2F4daU/XxgprX1LP6UBUJpcEsU6HP
CKkrusSdbpo2SlZS807pfxYN96NCY2i98/J6CvYXCOp5F7nnVBwkp+ZyRG6GwfO8
043C98DebL1Fmtk4C41VHw5sBX2Ui4fqWbkiWoQo6tOe6EzK6YdM8INg7gXHzSKA
6PqNfF8XKRUnfj7fGPMO8FONbnpVmhjYFmUt4eYbq/TwRQbuUeBvbI5nAUheuSbz
rV9rlSP6nR6J6iNgBCO2Dw+HMhb44o6dfh1h8hCJ5q7KddQQN39p1FB9wh4auUyP
2pO5KGPiDox1BBKmg9T4Fhst5fHg2O8eqxfvZqpAggUgLMV9rJjgUUtL4JN1pqav
trtufvoT7i/qXraXX2BdVbi2M2JGjnGhGNYUWHXP9NJRGzfmofQ0GRj3aOPtdkLL
E6LiUu+keLpLT/WzhHApaGL0+TmWlmFG05/gtb5g1+9xo6ndclqP8844Sqn3sYgt
WUdVPHXtKO9zbZFBkBp+vFyeph4f3fM2we8PUEbubMv3tD+u/erKRWu1wqiUn+KU
YEZpN6lQJfTQLL8fXK0OYPbBz2ZM1WY9lIZuNYNPkUkVgd6BIH79V0kbYr0hT7Pa
ppmLpFppc77mkiLedRciD18CD4hEtJb/BHvS8BFSL2L2eCV9/QpupFWWocFNO61t
soRYiZz9UIgcGRaCF0EBK634Mf20enCh8M/Qzf60tD/5ytRXGBxi81GQKDUGvp5P
urepULVAZMKo0upGbUBCkBTMCqYE5e8SdqGl27ofBYd0eO+bpp/x6EmxUS7CnwGo
A+D3EwVEITQm4MHEbnFs9qbM0io4T+sDKeXpAx/e5+S/+nZdo6xnw4afBEKpSQjq
E6vUC9dDkucHdVF5NkPpiRUwoi0MPO8sbwMpPNjPY3c0A60z9vMUIegS0e34MkhV
jrt0LOg3hf5VnQxIeJsaHqEFQyzT+Y68v55E1zcXOKuNIE2BihLm0sdCKvnUPnkS
xcxNdP0wsnK2NCtW29fVArSj9x4hxfMdNv6aUfhv5idsiiNWq7nRtMGK5NM/hmBr
ZhHjbHpfu/CiXOtV/tbejDRVkq2kfYTldzURa4Md5oKDQ7832bmIXgdCxU/0pkxM
2STQA7g2RmHMBClsRDFa9ND8Zz6z41o03oxKtB1IBniwqAoqWMm6d913kzkqWQJt
m4/0k01EoitbdO0gVmU99LivdGJ988rjlG6irvHxB/XRzgkhlQW8TArGFp/KTo9g
NtNOGQ2jzzwWjTG7ICLTE2+sf4G18lzmrUj0+qe/w94nB2pum4ZM3zhAwlUIfVgl
/TsfksuK1X8Ssj7GwGSORgnkoTcr7Jl5zHIeP0h90YMZwxQR/yyHxPa45OH4ahMQ
KFmVTI5+sdy2tzPx4HHignWmf9TpVKk9zz6/Cc9bCh0eeBghtDQHpJ0+dPJYcqRO
OGf7afx/+KBYDLz6Y9mX4A9teRSjp+OXRi8Up97fPX02ZmeRASxclaRqPx4PS7Sd
iRTdAYds7lKl+roTQk/js9ciEbgikHIvg9E2kkWsRhTnFotW+wV0OwmuyX32xwkm
Wtm12HGv8slNzmx0eoio/C4vHhuh0BihJXIkmsuqdDkL39Fp8eQO2MLt4OYx5hxM
ajfmg/MPhV0Eswi89/ujuaMXYfRREy9uBGsLFY8Z4UaxZxtSzeWUpMS6BXxZu9l3
kYyWfKTJsHQ6UpVQiQApc5UXRg/KwiXqeDT0e4Tb3M3QWR5ED+w1EiDZWhGvpWcM
pqnRoAgWktLT2CVEnaXrdh2SBIotIx3XSnJaIHuPeEWwOGRS0FMDqKovILNf7qAp
Y8xizJo0Sj3pEcZ+DMgfY2aXGVA2G6DhQGU41uKQZz76CXRh20LQzlNZjnz0Y901
0CKeYKWo8Y+TnbLkUm7KbzIGPeipRVrJGuBtb+Jj6f52ndgF0grFizkrpe2Z0kTK
Ljer59GiDZGLcO0d7dhTQi5SGb052LzXGFkwnHtIP75fRHnuhJrpRg0xfGOluInO
D4LT0J6eR385xEzKQKIS/C39LtyLO+Qzi/qIMaTr57n4NXnv1uQgObUaH3NIy9B9
zedXl7YocsK2kyKg1Bqo1FYVpOuqIj0xR32Pc+nEHHSlPHfuUP8eSlUsGK0LP5rP
Hnjklvq2JMNgxNQoHWITNnwI7v5QT3awClZZPuOnLq0VFxt3bQmQv3RyETYyveDv
DzVpzYitAfIa6XfNNC4mAmXa2glEWtdga+KcqbqcNQwoN1skTFIhu3fo5yYbcwdX
/jEN0RKBiIKXxuqth+LWjmF8IrCad3DNbVwh7ifTi2r+Vs3NLE1ZlYSWOV1uCghL
ohrw/wKdnAnXOXkMsUFanTrdm03wV4B0JKXAylSwuGCsk+bTKWotWEdSIvNBJKE9
D9GazLhaov4FCWgu7pTQKmawoXY8qk1lBbj8CsLyY+mt+6crWtu6n846UPwfpII3
YUEgyqf7cGDyjGMeHdQGfA63GJic6gIVxouHHy3zEwxhAbDgV7zRy7clcrSPvUUB
yAQL8v2D00da2x/o/O8+Mfm6lLkfKjWCHyOzlqxP91gOZvxTq6ne3yr/eWmIYUYl
yG6jzz9J/o38jgtME9YdZgBJne5G9Wop6DkKkemWN5M4r/vhSLLJLvtHxqT96OTy
+DtAobrl/++4CbalX6A4moFr/7Sq16NEQlcz7e+UqXv+uIyFc52MW005TnU5jKLI
OV/84hQsD11Jz2i1N1skGFAb/ZYODYv0akTa9LhDcEe/CVAOOGPc+n/J0/tlodmB
PCqdD9yHltRPOCv2SmK98fa0mucQy88bMoGqJ7I0iVrB3OzABp59BMn77pXmrktQ
bE0Mg71iUmSplIiKD4DO5DM9mxyO6DmFbvhNIatCClJsTLO6X5MYbLYToyQuZB5I
TXUAgIKu+rIkh/R6I0fZ7nBibzg12neSeZWelOtYBz7/i3BuyyqdvbwGEd9VKzKV
cZiNfENeoWZ90DICNVgqhhiCxOVNWpRDCaHeQifDpsSUO4oNJw3UZ7OBkfvCxsk9
ZU2gl3qwrSbaRTZP8q8W1id99ktl9oVBKMlAqWbgSFqoAAe3r7enQCKTYE61p2Uf
v5yNZFXTDbpZUl9pb42+IdNjUjjSLknVtIbVABe3nCTP5QXMODyhv+59PDQmMRcl
S9GZt6HYHx0k1FClOeE8fPVenULY4nLgmcuuco+oJk5k+Cnbk96RjkrRcQR5GCkN
1cRbsYJh+BVy/2EhXYVpdY4qTLPQU0He6XBNxAJHO963KZ3e3t8hVPNvx5l2YWsy
M2C7+0RCP0yEK+fSkdP4dpSDL1zLoFGUcbQUpGTFc2LhfsPCEdb2lOK9BPpB3e51
cpxhLIm4oogKbNxn/PJhMflm/VyIuem3UWzu8QTI1quryX4vnbQnGouv+q77tLds
ZXbwxejcObvyUDIg9Te5C5jCfqDg8o2wuCFUFj5AJePoFQirTbM4yIOR/YQs1I7o
r61NNT+BqS81CwuWxf8TwKmPtnUokbGgFT0tqs3G8wr7FeuNRGYCfd1pCgwce/E2
HGx8S5EZ1a4DyB4EEx9WmC3/lGa7I2tph3EcQiEwNP1R/RS//Z2cfozQM/cOI/2v
QUpy72e3Fkuqh9cdo+Y8YOQDIWY8uDvHeQTfPaCBG29kZ8ZryQTqi/hCXxiHxcOQ
F5E9y2qcT29dM2L5ClibKOS1iexE+Utx5cABSpu0RG1JZemh25QOTGvQdeBDou3E
uXtGz267wxWeluYXdY1rRtp6g80g/wweNpB/aOkM5N7sxAfhBy93u1gZeGxwaCkL
Z5DJLwF0fIZJK08euCjFuU7uk9x39nKck/8h5viHZ4bF7ReF+ZPlXzlHGJvEtZ3o
cteHxVVSkNJdfhvSHRZ1JsSApmSTx3Z0v4ywjbAeD8LKdnfmKdRYTT1ubEA2m4h+
9FYOdd7XkYuXcPZBmvLLq1hH1LFC6RIRGMHXsrCCRpHrLwDBmJvqornzmBoBYtTA
8rtGjd4PD8hAdvVVNJBXMxQjG7IenfKqJfMr8gPtk1d6epgOdxLM4wrg1S6wNluz
FMELmFnl4zQfJrUag0JT2vQgYmYQVA6QhwqFs0MzV7Up9wG2xwyGaW6wC4LzguAN
3kMJ1z1X587beM4zl/R8OOYSHlJK2mE/jV34XytBm1rPTWu7JH2TMWwRCoDeE2W1
/wtlVbRJFbqgsq+HuZrSsN7L8Buhz5KUfPSli/sYqeMMi08CFsCn4VNluJga3Gsa
ubQf7xWcBNwM90p+KdoeUC6Bjj2r2YjMH21EZw+Fr8XI8yVzln8SDe6Zqz/KXZ2p
USe+H6lzMeFTD8Mjc82aTNE8kCX0ChwqBZOSqR544uk4pY6Uyiy6stIwnn2nwyzz
MsyyURbc1o19O4B5gKmxaw9jjadYX1uItZdiFFhf+Jtej7VZCt//1ZKr0YH32oYA
Gca5WMUVBmoStni4z7WeNqTENRHFctVzTz2iaxv2S5KX8cU/IBoMUK/i0REBluPT
USXwtdY9IFfQlpGjm/8+K6obnDjD9ZJL0pYjUNFv7Sd2F1H072VPOtL/o/GzjdEG
s+we4xbIVk3A18RRKEkwBfEoS8ucp2+x/mhjKsh7s2yYmga/zYSdsAlOxSl11g3s
mCDZeF5Hvmkh6e5G3Z78TMl7uxVVNBfEZYohCg2ZqG2z7hENlw73lr6EDTvHcj94
QbJ1qFIfxPaUEw5KytqvWrQ/Yn6y+DXaxUW5yMIcSD32cpjB2ibrJNhSuiSvSfVp
nYgMkPnxibMqVBky45nb7HT5ULBMCh/lfFaW8w0ZmSiE6XtUbInjuxqUQQALdtPB
lhfFGIdBDN4YVeWg8T8M2nX6X6xJc0k7uKc1m6QLtvRTcQDRBykE+DSt7XsogCrT
x4jR5DWuEzU7Izrl/i/gNpKcxZLyO6meiCUwXMLeL3e4Absj3RL1cR/+MihUkBTp
j2XwNcYoIo5qbR4JlZtRGrbH8WFAtqCO7w4B9eReDMQZOSpcucQedW5Ktck5AJ+q
2Y9wwRH9iAwTDSjI4mPfV5ri8XUUvD1K0HL/Bj7SjpxCWiOtnLhrvVoLdfqK/2bQ
ipc5Y5YfU0BBaIGZ26szhME84914xQdhwi8hdNkZ9PTj8PHUIjCsIlQt+yHBKZpW
HDwg+EmqlXxR+aQG6SSYGraRQHk7ZXFAeNd9wlqANGzq/Ry8ymK50+seTzDVRqr4
Y99gdfiMMdd3mG1NwX+gIJazP+ravoND6rPRvqRD4ryK6w75Xwy9YOOQxMDdxHOw
m5pGKIfPG+QZtrZqg5zoSRbSmz4oa6vCly0VL+2H+GmBqC3owxtoyNQFHfhqXvQg
tDkBRB3pvTR/uM3ROt2pt19MQBw6DveesfTsC1lMc6GZwTJLlzbQwKi9T3Q77g3Y
ZwH2XZ/mvKHGsd5DeDsTuqlfa5RvScqOP+4PhQl2QpzPtfxrwSnbgC3c6hsZYczD
iwwHPyJBCEj45rbvWnGiiEHWAc3vQTQwGsBOOYQwTGGaKExFORfHisS+1ZTrbvrQ
DzNVDdZFcJT5L0VjZgbAi7j7L8W2/MrnWDE9pv0ipZHJuqukfP1Cb87RvwHOQ1F5
0q/TAeS9j6TcMZCJuETFjbBJSvTctYl6Am4k4xACgHjWmX3FZ+sItxvW9vmZylMA
zMgY+1J9HT365jv1MhOjJFtjMqFn53tLsGJsfz8jiLxBjCeoWlASHkNG/RhT+ibQ
7lndRZBHQJ8JNCb2Swr6u0IeA+3vuY8M9ALQfXhdfOTUZI4Rvn1UOQKYT/mS8Xu+
K7BUivd2jLW6qrEes5WblE3epKabifB4mlxVSMFy3D4JTaOPOJbSj9fuG7xKnRuY
ifbkXUiQr7KnIYK2XYmLDQkrTwF/t5mIalAXVI0otPwhNnMs/f06ElXHDw2IyOmL
9X702XPIaFcVtOW186x4A1uhfPBnnNUaOUJ0jYDEmGTrW7ba0cwdBno7xbPQ/aeh
CfRVu9tQyT0ipPxg/avLS8jKNFAuiMfadYT6W5pQsxBb0CHwOIRGsF/NxLg8grVH
63P/mNuO+PngHs45rf4/dG5e/HnS13U1WSY+zsqJNWzqqVjvd+eUz0NqPyI7x/yj
2DFuvhdRyf9fVnicuzZoo98apDDNjAtMTIJImYtJRFm8oecByLIWs0zdl5Aank5e
qyji1Z1FgYfkKJ9gCtQ7ld56SJe5psHJHoICdxC9bhQZsVU/E5XQGgT8EC874PDK
6yAMJo3ZbUBXmturrmYroFvsthKDeae5uMtn6N0RkN+6jbjwZZ7+W2HOBn7VCVkt
Vj2QNrsyP4DRBrxA6kN+atU6EOxkMIryq9x1rTQluB0YhwcPiPKWA2O97JFmf5kX
1cXk85hXwe35nQCffCHj1U9OAmSG4B9qJLtqa69eOrjSL5DtfPDwcrk5CgiERqAo
LDBwtcsQ71xvnOjCG2APqLkEo9cmmXgtvyF9qLXPfDU9cRGUD0ATyJ597VxnLvE5
6ep3/VOZXi6mVJMxwAGQso4RSte3PkIJ80+hQuVu0kHJxN/VbRCi/BojkhP26VeC
2+i3G+GLfZNS0WL74axLj5LsEevaBLehnrMr8LP1FFJL88HsYuFZHA+Hq4EmZPS5
FGYVrxmny+t0iHwAwSTMj+k7quQmTs0VnwTpn3MXlRTuAaGzZgrYUAMc/WZ4Tpxn
l4dt3F/lH4DsYy3mj0EcE4/wEdC8T9GueUUo93SfaIRQSG78rgTea3SvVCO32mgD
SOFPyYO56J/RLt8Y4o7gaKQfAcYbW28lz+6bqEpDOoMKxbnqp7fFhthQfdg1jSIg
MQvcG6Wt/wMsdmxuDMH1Y+lpe0A/EJPnEycM2XPvKBBdkB4kCt09U7ZvK+WUY5zN
GCWQC7nkE8fSLoJ0qEEeQUkKBPVXmtPyX9UpCtU5z8TEEvIRouTFjGHutRgLYxn6
kx/M8igMKwNmkLjUXulfVPHu+hijL19IuLX4N8jzNLLTxsfZHEjxoVtRsKbUjsrj
o9l+bwGeqHXga1GOCHvtmTjOB4c9NeFLYb1aiIvqnHc0RzRm11dUPVIj7asehZ6x
MoG8M+Z/G8u+UJRsqlz044nc3cpgEWCYnUdkBz8gm0YS2GgRaB2pk844qLDRUtQn
g0w6BxNbAryxa/zKhndk1bQw20wPBG7NBcxfS5l0YMlgGYZ/9VDxA6PunvV1JTT5
bplqguy92J1Js73fP2Fuvkea4Xm6oGOrPqhvEv7JEMWj21Mh8NPZ3L9yCwXkT1wz
7vWbXLAwVxgUumhjDbIkIwwhsfsYvYJhFUKcceE11eyg6z6GejB+//mxV8fNBbEl
YubBPfJqQNuyqoDyJJBHKBNYSV3vC/xBqDl18+qrUDE4d4Ohsxm+nCGcda00/KcT
aY8WxOsN/YBrCgEDVxJq6E0x+WVPmHLxlsYjygpxjpAOw58zoVX7PMhjDHZpDoRL
akcnn8EbZFGp1tIsVZrSTGk134pR3lSB7iy+NmAN6JeGZsl9hm25kgjY1lwulTlC
ii6j3MDR5Zp01L6niY9Z6EYmFpUF7YJ0UEUeh4JRi4wsBDm1g4EQ/XPFKNyZTEdd
rJnZ0E3zw1aqQ4nLlq5LjkljBgsuG8BqpAN4tl0P1WI6v6WBTuaz9MZTgabg04NK
J8mD3ntQyMpm5Kh4Biy8+NkC023sx5JvsfUQjS5ujvu2vUpgqCrdvQS+s1S+pAoL
vY7UIBQ/Yv1WwZLBmuziORP/NhhDOgnvgnAro771pbf+TbToqjKWrptiQdVkMIpM
IvOtjGG3vlDBCoaWR4lt+xH3JX22kKCCCS6o0WCoTIwx2f6rqVpwIis8N33Y+78F
zeKm3g2cVf0cSNvlmz/zPSuams4C759WuR1DwcmqWjYh83jldG8ZRdCiqE3lAyDY
pFqZk/utJ0BCOHgnYuxhUFORTQNw15qFM71lYa5Fpx0HM5hzShF+n1tJaNejvfMH
wIz4VGFQgxjrfTYydv+w6dLfXhGg1L0zz6/ciFhGk4mE5cpF8mJGxzSqQo87I+5M
GZWisum1aqkNWKzEXqn0jazmcP446vCEcbP4csN1QMfNZEDruW5lxhdPQVWFQ+oo
iR0uNbGb6Svb47OS0QQVopLrMvbIWuzZMMn0V6DpbKokI+ajQe3PDsPXbrWAYLa+
XXaZG89MRk9lXkHT35AFw6/jDpw3+qs1FBLV6A8UsWqGAWw5cBijCOjGHlPxdUoM
dgInBWy8X1+pmZ9i/N+Bz6Gjy/k9sOTHWsGCKaCPuyblWTz7zVoKhh44Rl/GfCKi
XREjnRFdOgyEco8t3KhSPfh0VBxMQO6wbHtmrczlh/BuQTaQ0kp+YBijYq2Rjayg
tpBRv5mAzU77A7b+0mE/ZyZo7wwV4K+ECUga1P79JwKgybYKrlkKMV71KDHIhDCR
X7ZDPGSndIpRC/hzqN2ceCg6Q9IKrMfzRyGMRF7qmaweuBK/mJfqJWxzRQlpZE/a
yaJEHuHHUlGvwhs6O3xuzPOzziB8kqqT5wTb0yJtbO79JjJwYSnZyCAbIBSo2bgW
YEUIiEOaHIdIHzhGpg5RJNWv4241ElMAteoZXLyDTv3UgZmdCjF9tXhJil4atxQZ
yUQztT0mFLSOcmtLwy8OhR82lCueV26qJvTMmP4Ivmtgf6XWUao4crcQxtQMvj3D
lMPkhhBlezgU/4dyngiXJ7Q0d8LZnnKpTOy7EVFMvyyVMxghJre7q7ZdQwsW4kKz
RvqJuHaQMhSs5nWw3bC8Gr8qE9MPyjbVmos6oQqmfClJ/Llg9cqQIlLtGgMqICry
ilf62pOQroptMmEdDBKjR14aa8WXDfCtiOu2a8HgZSWyuGNIm41UU7QcOPKB8vwO
5bJCiM583VJNvZEG5ZUE5WGYGHgWqxbmR616nAFXUKAYSoVssd1bsAYz7zBGIWZr
HsJlgZDn+KOWieNGPmYUlP4DLxPlySQztfVWYHuTq1d5tHg6s9HzS3tdQNuWltR9
xcaIXGRopsXZxFEp0gDJXGFiPyasQ7hXZHrtNoklGzyeKgz76/ehb27Z4orY40EG
BZGXs4y/5feFgbIsUDP9GIKCcd2AErjCvKrzCzQ8tJ+EhBop9Y4W5FlItRvXX4yy
zYGClpkeEcb7l/v9tPY0NI7HtX30WSumAxgfP3CQKoOM0KkNUrqZ+kwySuLY5M8t
mEI6xmiHVTuUAGwzoHg74Mamj5Xg/ZT3WN5IADPgkejH4tlwahrCLCmCpQBl09xT
i3ktY7D5bN7iKZM2kIPFhzHwhLaCGlZR7h29Lmlx+/WZ5cfJGBoGBK7w0VehvMj3
ApnPC9rgEU5e6F8DUi8hazFOOZvBpRtthnjSs8XVm+y21ZXcq2n+8FCTSip8MvFd
xjlEyt3RAzuCZND3wVakF1ESudWTOtoqtZ49AXZot5ddwYwmvpAtPOGLHPw+0UQq
jhF/6dgCJvNjl6a5M1M5HIxn4myunLoqK7zDFdWsp35a+pJ3D72WiJCSY8L8S5NE
GK4yfd5oW23temeFEVQOZJSW1W9FGgL8ZLZDHi5MFHJnpVfd3iFF45nK2OHFauRR
shfNy9esj6aSadpLDkrBaVaQ4OxhgTzSTO5MfBfBYvGzNHJkXSGmb1od0qtOaIkO
z84IC9TTP0XJqo6LmYgloSJRf5ehHZOyB8jH6GPk+tyfj1qfJCTQdV95xPzBej1A
eotTrLzM3HqXzyiopR9Ek0IvcqFAyCOJQCF2VNqM09ACi3h21Av8aRr6epVZ94T0
DhiExy5lDodoYCvHlVuIBFkPgHmhSpZBjSklCV+jQ7BkXq1Ubqah7aXG8gNaT4kf
a8f/c9umJL77tad24bpqINwHf4mKmDDIV5FG7tADNw33Fw4vcMWu1Lfwse8btJgw
RnaKjv2AO6azB5Y9Ks1yKIwg1VTYekmpFBUW2N6EbadgfKqjBmW3SUZQp4HqmxAd
2rorYVY6FHp+Cb8tK825qoOFJ8kGEfEcnIUq83L6TezC+eCRsu8ovNp//kNCa7UU
4mVDXkslPzSFSy8gTyQsDSsPUruw/p8LwculEm+2PlZIsHUbPipNWkUhy+dd65vJ
Uwv4uvSox3rNbPOSsQlfdJ6RaLHjdsf0IU83iGypbzijDb/Iy4WGsAP0pUQooO5B
/WqCc/g5Lezpo8iLhIBD2M5KmikJF+Zf42vdUYGnL6j9480FxGe36zeJtNJTS2sk
x8ViyUhjo2KmV4SPNEJLf0M3I5KsNcyqmjc+yGCKGF/fOZTSWXqq+q4OlrNXyn1K
V7Mt0d1jysdVFGUoHs6kpqmbDHHUkMz2TdxLkNWeK+Bn+3gEaOH3efa7cVQSWVDQ
bDmHehIIVfhPmLLghejUiRbM2C9M98/000wd84aPO/r8m/PvN3ry0uI6Wma6jp43
iKVVhVyMHBeHitpFRrdI02Rp1dW3aeyBWuIgDtpGUFynUG+x74LW3gjRp7oRFwqn
hk42kI5UTVt8toE77azLjgGM6UwYjoPUflizD1Vx3WjwIj9eDCeO03ngOJ++K9ED
BhWW6XFJP4dzFzt3zuMVJzN1l7U1FBRoutYgu+BAJ9tzjP5hu6EfjhNEiBN8zQXx
8K7T20I0/ASfVM27yIssG9vmGgyzLT4Y1WBYRPOv+Lb5Zc7F8N7eNzDffaY2rxlF
JXd8i2cF5Ely/FbOSgx7WKJWYgY50ObZT/cpDL1paijepltNKzhwQ++4W1IbYsKz
wypXvfQM+SSa10sMLTZFdNNinfijIYnVL24lwi2pL8KDX2kcSX/TA1R3tft2o9/v
yevnTpJg3B+5uOVWbIVFSK0k5W4ovHPvskRlxCptZllOt93wNG0Oc808Jl/dPy1p
r3pkVAs/6hmY2ikDkqxQaHuCSxRDvg8yleJS+qgyeugKZH1ZHT+5ZnH7ciFlMvs5
SBNeo30GPTcAUp7pvOzCWHyLG2b3o10bmBXfP4Lh+CMSCndcpfRfDA/KfAlZ+3dJ
`pragma protect end_protected
