// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dX5Y3ZN1cZYC0Rm13FT3zd/zS8nWiqe8iqWvZAOKDyQQjJOg/67UUZjQPfgG2VWK
VGDunlbCejLfrmaximSQZ56BqeEGKFJJ40zxJ26UtO904lGdBw1kSj0vlYSEjJAe
XfNZFm6e2AmxWQN/wJhWnIsVbZ0cUBdOES1q75SIuak=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8144)
IRnKmP9lvYk6ukWX0BSnQf12Gx5gt2ILdsCM/XHbmCDtwq3nPf9EFsvgJC4SSJx3
obBJt9t+cCTSPriyF/AF6fFU7Ueoh1Dv27IowrXE/GK6tqNli2h8e7clUix973eT
qrlMUXaxpODW/sQVecKkHuCVvzFEMwYnGqltgs2rX9Bbdlf7VEGyRFma853bKAgz
nt1BoX8qlxwGcX5pKFLgt0JEr+O1/puZ5AOOPKWyvbcqIQgePMu62qQhu4OBvI5Z
+BIOEUGepYL91Ne2NSkeY7w6ycvRijtm46AzNrYAZf67YwOxqwcvDFtfDqnPYGnI
2akmtJzsszXZa2bokonzrrswmMMRYjJ+iZwg47568EWAMETKtRwTAGFueoCY0Ouo
u/Sf/E9h4oVzo5LKaS0vyDOlAFR29Pn64r4wz2TgzsEdCm5xQu6TZPLBP0PdeOWY
cyRoR7oN2R0EkVIWDQ1PvhYoXvpwKMAnnjDTyIwk7e3EBch/w7qqxvc80Y7SrQOU
GuqX1NouYjosXPspUKFx27tL0eXOItVW1vHzYrzC+NJ1FfcGcANUaIc7TS046dmi
UiyrjJa7wjDlq4OKhI4QDP3Ora7lWvvQ911m2FCMBGvsTgsRa6tmK+ZUPyUVtfNH
n0PIz2VG4gEGyyNy8pNeXPJqq+4Eg+Ij5xM1qMqYSFMjbzstPmRQ1JM9e4CWGZUv
E1Dm52akE/QH8vZOUg36gGUM1rwIRrEAV62InSKXp9pSXXmRb2zG1XhLxA6pGGct
E0oDQOMeAVK0IuTbWl7yFiPDcIJvn8B1kOcQZjcaFIj+dkg2R4fzeK37bYSoMWX4
yIyti3RiaThbYF0jhViXFKFy+50/iJ66g8SKbyU7B7pmM2Oz/IcoLvqjZNP/cqrm
ipuK5SrCG1cfD/phpD0numISlcdhmqsGjYO+5DwTyIt6lYjm0ec2cGsN/tGrQOEi
zKjyUL3L6LnTMAMt9K/51ePBVw0xr2sH3oegmzubhTke5xdHc8fXEVFu+vlbdxoG
qyZdtheJueyE4/DGzGEir2upzpAQS2+er9F2uKVAn6qRbp4lOVulpeTPzjvmVsDP
ckwLCNyCIuh7Z1chrVe88shGemebH/aL6xhEksjQq56vevcw/2dA7ZU6Uow+AC4S
4N2aW9vycDcSU9I2xDsVCrU2WEmAbCwNbluc5e3YSM12LzZQrq7uCbysOIyERAax
+HRXDSB2stFmEK/Rrjcej9TR2HzXTZkCPqRQq5eJ7Q1Uv7CvXt+Vh91MIILE+qV7
eBg/KatL0q6zTvoaPC1rSysNO+XMLKq941nBSXCNqU2q4KpP+WpQm55kTx/MgqeH
iAsAkBO+ZS5gQavdjdGpnj03WLBrKqpoeUROcYn20T6NopLx6jAQn5Sf7I2JlRwm
SQsxnFwF92/hturWNTYSIc2QDcBKR83eNmyOCKcxbgpNY7gYyiTZvne+hyMD4dDr
vcpVXibz1eW8IIUMQ4ufDCAoe33UDhEUiHVQFRZxeIMLZqaUJNZscc9fOeQVeC+s
PRckeGSITB603xVn/0VJm+5YfF4d0BDjQM2rZDQ5GJ85ywmow/VqwqS7I7jhjEek
b708ChcGOkrfW8IOATrANbrKRhJpynctIFzUb6CX8HJhIoEhfR+WBYl3szqgYX0Y
HQuJVVRzbZrBWvuuLbm+TLJpJpEKrV8jLls5zfa81FF8AZEZPqqEI2F5nQ3ONAHU
WLtLe/ig1qINVSb2yIDyJ/42gjpfGeVfzlNzbfveyPMHkB4ZBjLJITckUQM2SyIq
AxWzGwKi2yt096rhLBzPiRkmVOGuEhDI6qftn/vz03fi9r2dhJFPrlSCMcVK7mbq
UUoonVj/8cipwa0Axh/qF1p81P3Bjgqxro2GDpRrSArpPaaLL/KckY60GjijO5Lc
3QIfP75jq9HGN3z5aU7L104B3FU//rD6a0at6y+Z4m77sVMlG4HQDyC2N79c+yCz
KF1bQC7ApJLnfvh/ZxiewljpdJwdMwfIeC57Z3pg2nZ7AtwomGfdPZSUBDl5tu0M
+Xsp5q2FY5TTxn334m8Tp+pudGapy6wwCmijs5NzODnKOLsQhhthdzBSr85sgO5U
c4uPZWbg0sX6w9dzDywBqodhWpMo+CmEIyM5eudOtG2wTpm3FS8FkHY7L094eybK
DcOJE/yBBom06ifWgbHj0cCkpG4m0pU3TthVmfdz9C3BX7OkuqLuzAKgZWyugz/r
CcKRwRCHhOUasygtETC+Ftc+OldC9gNw1M1qKT2vhJ/TeNMTyU4HgW6bspPFKZed
z9z/ID2QkMPUU2uoUJGwyMbjqBWtdrwKBJLDLEtJTnwuiOuj7DsJKu0tGMuoi7Hb
YtEOZtFnqinqHR9P/hcm1uqyx2sw6Pr7gk2zmSkUmL+CP5u0SkL0NcfXLeDLQha3
8GaEA+0kiKYGCVWs6wq+N6h3KMwaOvKNlc5l2TZUCBCtsi7bLNpFO6aXvmv11yvR
6Mq6L6j+oSucv8Fd/zJ+stkaqJ8QlEPdmjHN3RmvsiV7PPDYjltOhgowRBAA2izJ
+uHMyWDetZqqE+Mouh2gWm4fZaLRV5VpD2h7xYjZgD7EdQqQ1v+v/JIbRwBYDhdO
C4Wy5a7f+36w7avQtLM31u/x3qwYEC6oaShnxsCYD9WbytjlSwviE3sBmstiBbGw
NmO6FNrresvb+CUtHft2FNUlsysdVGg4InH9/ldnZg4bcLTyWaGdpHOj7N28Hba8
vOd7TBLX0PjH1AOqq3KqRAgLPV2nfQTMgRaA3Fi3Rv+J2b0SjUvwnwfRf1fUuJ6D
yQH5SJ9qKyj4kyipN9DsgrJP0ZwkyKt0tR6V1trQpWV48PYS2xdIE+uu7E1itYr4
EU42DneGn98Jettk+6xj6akPG5kXDKn/jCNvA53xMcG7i4GqqJVkGOFrsjDHtpJ6
X8FGi1RP+ssKlvn9aRuZegC0NggGUAsEfLCyXfYMFhhwcuAPK+6k9X3TFMDoG+rK
7gCvWj4+0mb8OUrd08ztKyJWO+AUFfUmHiDn6nILV6HSkBXQ93yZ6+rGbB5eo9oU
JCfAMgGXw5wYGGyaVzQ+MUdkh2NWiLLn8rd188G7fRAhVy/jCg/Ey0nM35aIHjJC
IYnNndCxgl1TWPZ+aVX4g/6TcuiCPFqXJXEgSgdWh0a6juCxD44OEcxCFzSIANe2
exPlEHbuZnMuqfhfqRjfH83dQVxN89ws2yfwBo/0kQX3xDym4XDzeVzGbi5a2Zeg
rKc5V2pbg0NaWiZ7GVp2NvEW54nY6VbgJf58F3eYZf8zOQF4wonhTPMIvnhvUTFQ
NdAtReUJmEQi/UpE59uXwrxLWBAYLZJUtCoeAeDCuKL+uUnPcOsft+sB19l00eiS
F5BEUb9hdsFhvLT6pPUqBFaY6vSOd06MInr5ObcClGuvcjQiUcY57NraWpklAtjm
Fbx9tdaax/ldn2E4hFnscplyc+lp28n6gy9j5k1OXnJAGd+IGX0WzH06tXPzukDt
qy/ac2R2okIc0N8sW0QNelB1KLtfNygT+A8oA3B9DZHjIp0YK8wnIlNnG+yZauy9
js94YbmP6PHOJ2R//6ilK8VixLq+wToakvx8m07VSoA0wSiV/D4KApbIZy0W1Vo7
bJSBbxNWCRcIeCbDb13GX0daYVvsdLBZADRq7SLREF6hCtIeJHfmIuoPJ+yGmq0g
LFf7M8PAU58g/ErFSvGxoJzqD3YniJln3CijNcmKKT1Br7M+ty1B6GghEeFtcne0
+hFkuUkOnrBgfyXMEVJAw1+6/5CR99n9XssLdFOol5ogJhNUt26OqU7HIYZTUgHP
yHFZKR+CQ+6eUUWcw4G7oPHVwf49RUCfahDQkMhi1I/P95sNf9UQSOTcraiuuEY8
OJoTK41Bndtai84v9xKYbgoPdhVlbIEr9reAi/ShKWSAqQGJempW8ZB54erspWAN
ddrKXiIaNNTTnRStrfETrHO+AnLxx7PbOhtpX1UQeaO4OG8BX+S+Tq8zHH8sKAHM
zbcfJTcSZsQ4/m9eaYRqtZvIifuZo8m6L6pKpTk3fPzASqF3Km9URCBZRAsUm4jj
sazN72yxAf+pEG/xuIiZ9IH9qsxHMITYL5rdE3yA2RbxmTUx6SAjSrmfLtMsCL7u
XfwV1jkuNc/MkmZRYWGmNNVHLVNYpeni/dj4I/IXV3pxqmKDZ46rN0xdgJIdD4KK
CAfR8Sc0EH00x4j4k17QBV0RWhcj63ADQWN1RBcyI9zUipmKkx9uPqCgZnaolFnB
jJda3HPMhWSXGZCqjQ5w67bYcqhsuPbqSYc6U5CWlR3Ogpm0pIWTGSSe4Wm6UQ9C
0tn3B7hZPUIL6d2xJ8ZzLutAwfNnvuOOAEEzP+BiwzQKZFCGgvSCk4HOccp+Za84
So+uM9yG5iDMRb4Qa8XcozDoZUVY7keNnRUqXS5IrXlipt98tfzdfTxmDbUn8Gi8
PhWgsXQCNHZfp8EY6DKTIDDIeNkiqC41d2ZPcan7nX+FOdfSpGqe+t8EmU1yef+s
6D7uCCjfhqEcGwESc49O93SIDrAjoExqEGEqGzbMO2zROOkKX+VQvGBjw279W15a
r7dpDSIakhZ+v529Jn/XRoq7H5OchsKk2QdnZfDIAVhhwBuAhB63E2xLDP6h6ZSO
cBFbZl9+bhExQkssEuXesl8ebtZZevrCcU/cCiSt3dFc507a+6vtT2byWV5r7WQv
arGBtn0PmGuugiF7nGn0/MhcVIIPhehk4eepu/sK848vhX25iX0VAzQOMK19Fgmx
43o/8UqQn574fafDvEdksZdqIzbLICa5ur/k9euJ+qFUGfOU/76KJeo2BQ4RQgvG
BZcSirOGzJj3/FyCdAijN90yIUZuPnZhcS8vSM7X5+gGsLEPbbBbiyWVEH8QFAmd
u7hgAU9/M1qmplPnDujvKCN06e+oPjyQIxFd/oTAPl3DTCOmUPp+O9oyRqQSehcp
KztroLX3e6b/bUyrOzYAXXze6OZO4EQivJv55Ioq7ZRaBVcvuEJGwzcI2961QFu8
PiIcVKuuX5NbXI97V77xbccWYpm0TjTzZDW1LmuQAV2IxfMRGNAnHNVPjGfEvIrK
iEOFgEc1H89wnmTDruwz/C6vuRl6puPAybMUxDSV+KnWousfomHC9GoVxxxgtXkZ
0upZQ3T/wEQtw342O8uZUuDOWlmBFhhHWTGUS7z4V3yTpsU0Kd5ZCCPpD4/ZhQhm
aMnAnUnXgAAQ+bP9NYMknw3nhhoxgDeCvUGOjFYS0qLyJkAGuIVR1Ix5OB4L7poW
SBdN3ojIFR6VpTdzTaC8Uxo3EoYklB76yz+kEiAt/yGbL0nWQgs+bYvItuir4uwg
VFKkCnFBdItqLfN8OwkTCWg9skEfMI4raGnXVTr9OpsbOFlfLbntMHH7cKlBmXcl
2bHP/TCli8+JuIt+ecWt+TdZS0Z9/oynaEwBLCQzGunP4mzgP9mbtndA82zCyO3C
sbX+E6UuesdMp0LlYWcDeXg49z+1Sn7xFk2KQ1uTn8CCGDmOpt4LkWWOpeirzKgu
mx22kMFRehowlL7l4dAXx09aYNLqmEhO63JN4WuRI5f9FDSB3jq1E3s47MVdUXXF
CYRUtslBO/BM0s9bOZpYBSBNuQ9EVod+qQQyfU3ZRQL2RC1+n3FIq9o+gNs1ZdLV
eQS2z7JUHEjLvJJVZuRUwruhZJe5GliEL1/FONSHSGA2rawitCwhSRv16QFJkRvc
xpIjrjLzFUUsi2dhIiTyvMhAXRrzZW3UoJ7zJlZSvt8eHb42o3ui8gUorgYTys8j
EHcPVC0MWjuWk6QkWyzhwnh1GloeBKULu1yrDQTUpeI0kINNK1dMdRz50CJ4yUmm
9dKweNXyMVT7YOhZSlDb+2QUIbRa2IH6XZIeYUoRnBbNMoO2pYmLWctIJBivjT15
TsPGZiCg537zb+3BZ1tu32ldGe/nvmzQXIWqr1fG81zVT9jYVJu8GKH6kbC1eePb
Of8nnCFh0NSZ8Kye7oxELVLECNHCfttPnUCvdFvb4sJNVLxYhQLWsPk9F0M8LFZv
XiRji5Usxb4zw3E51McyTprj4WkDDa1d+ape9EiQJ+UfcrNuRetKURIj0I07AALR
4WPu5guTRQlnjqCHslx+vbcxuxpF0tf0yFVcWtIFDlMzZE1oZTLHicbGqcUFn3uI
TzE8f3+IYOlJhIqTIyE60TF8vYYP+AobdQ0XHPnBFbukmWxdKac+iDi/d07umhwK
VbfB8C9hgFmmomP3J0i7egxiYhHXsvSdBrZ4aV5LQMIBt2kvGlN1pP9juHXxjzST
5zfOaah2B08u4984Ce6c7dW8+ffHBTfBaAbuk5uvR/K/DJeQsLT7L4vfI3wQk25S
aIuwznzu0gJ/j+IklrL1thZkMMbNUwBQu2WNCFgAl3zTmu1kzRYBYI3xGDBh6W4d
riBgwnTCMynub2u0zH1emajYZc1Zaq8vdNfx8vR0+5/0CdPfJXcS8tMHjaXSzo3P
VJ1sQXQKmu+AO8eT/JND0zD8q21nPlKWqFKkIfaMFTWHZxuGMscYpxGDezEhJg22
X2w/g8xaaZESYfzSj9ZFfm381AlmjgGDthxZhYA1LEgJsFS6fjzz9PCSkF4erG1I
ioFiq5ht3jrseFU+Ft38H3Gzr3uo4QeDUcATuGoLk6xVCUcYkoUvj1cJHgJwnVB5
gIUizAjDLi5M6Ib4z6PO6nM5Wm0zvmnr0Vne+CZS0LU71yxTVp2o89vbz52ScgZh
KY5HggSwYObn5aY0B/5CGOu/LEJ/3XCXhErUHD9XDFISx/CizBDrChmnlNY5351Q
ZZ3EMArNLw3xWG6hRkJYiXfPmwr7UrnOTC0mKs+y2t/6Qs3NC12JZFj2pCoda6YN
pBuSAb7aPBaAhTAeaoYiZsYpGriAx2FunzDxuQ4R1tee4JS9Uq4oUcby+2T6zQgn
oL79CmRWseN35auMdcuCPY+VMJIr3gad4lzHsQQLDQiCV7XbyWveaAy/7VNbotfa
i+3fDSa8k8SmfoiZuNRKslBq1eF0HUOA08iCrlMLnE0IYOMUK7dwsl//kw0WS+p/
f0SeW8BQPriZ6N7g19DMQ8EANjOWPbLqHfID/W6OIO3LNt31ea6XQfs+QQ3/Btqj
MBBOuSu4vT91tPI9ZpvqsiqLyzTg3uEH/2wxYYhUpKVQYwcLtlYiUXCAkVaNZHz4
66gC28xw5c2IX+S8drhQZumXWS/YyRaEShOZjVY7hTEKSTu0r6ZC3rOu4c5kHdJ4
/PbUAP6k6/t4Vh5D7K+S9Hf6lIW60OIt1jBsI/u0NLkC+1Yen/FuaVvf+BmDhxE3
vfj+U6tx2a88Ue2EnB9yRMWXzziYWPJRSc+AYl5y/zEnzGyGkYyVpl8ZpCxbmP5T
4BZ+bBRSDt1j4zzRSJR5sxoDq/6VRsWGesKjprIeIY1AUSJnRnhYBTEceKwktvSq
ddyts0duL8skpDnj91Eljmw/LYHq1WA9FO140U5C7QXJqO8YIHcfGI1N0KxGQvJ9
sHGryBFKzjnx3Sm5Ox4uWJlKmQAsLCRYRp2vA34xzlftEUd3c0I/OrUcvhCxG4fb
uPcYDyhNH/cCaUy1jwqeOoiCPzsYQgdMYSCReAyzSH8btZFJ7BDFJmWKHjM4lPdl
fI85lxsEUThXLJJ9kzrSbNl1DhQqnybsuLiDWbD6N+51MNGXQJ7E8qyUFlVsskrY
YKXFbWG4oV9/moh9AGcexUYJN4QMVz7w8ct21k4kLXtPUJg8L5+5FoUzZ3QRAR8t
oSqNLYEZoNRnhE0RXmCnrQKLGFAdUowvx/hu6RVYoP/YZ4AZXNxyjgocpD99hLWk
JSsjV8YJW5Su3X/S5YrNktRQdc0IlxE4Sa0oTEZWPqruoldpkvuTA0XFTQ9Vwoq5
swGon7Ej4wH7FErudUSeSfd2v9EzQyQcwwMIyNt8yiODhtThltyYxuy95+/tsa4b
dNCvtDiiSRKoMMW2sY68pbUw1VQtt0BQosQh2lnX7V5IDm9DvAAleCVt82rtJC5e
ZgetAKHudYNz1wOYlDcSacDq4IuL4Yk7jrqVlWpZzZB0n5uf0LSJv+I3lHRZQ1h+
vyu61DmWcm9jqK0f6F+MvOhFKpnn904vNfoGn8Kasks6evoR/6ewNs/tZq3Zj4rQ
b2uVYw1MtIMWOwcmDL2aGSNC1jnCY+Ij3vqG/jv2pVdkNEaLHX8Bd30JHuQNwG0L
z2WMDV+PwfWZXfTpY/RhdpuyUbpXM/S86v24uY/6c3BIn5mvk3l4yH8xcuntXVPT
nuyUNj6eLb3IeMmlsZ75wrpSN2cuWLG6lofxWoA6GkqfkbGWTACjiOwuubd8M6No
7CHyoShwyxPIbxdAWRXsnkktUz5LSgEWRII/sAzwZjUVwQ5xIg4XqJNW0JcMWB83
YflSW4JlLH0YVk9FIN+s4P0aHfFSwfT57Khn5oylNekfnyUIB6evlVEvB6wohdGh
QriBTZACY/2HNQLS/D3naTEY4eXKofXGfQMm7hbzMaD7Wv9hsO+YIOY+A4EQKWzB
H7K0KWbVlWzYVHbBW6TtG9OhHCej/uQxh1OBX7I2poQkbue/QW3C66ztLoS+7N3Y
n1m3hfLMFlwxGHW3RMv2U+0JvLfhMx1TOOLS8P+nDMLsoqeWTEx09BblllUzH8sQ
IqPl6SaDBWWX17gob0PGnEJgHLbvgNrDPJ81fb5FjAsDXcybO33t79zgom7vNVR5
uOuYlb1+8NAsC7KyPY9nOagl2whYf1ixbHinnfHIPzYoSar/3zdQlhUA6xOerN2B
sStN4i0yoyb62oqXfY1c4gYSxJhLm5odULI3ZdVbb5lW2qpL+uSNuNE6OVtWAzhQ
8j/JMMQ918MrBocLmgMk2d4FfCtZU4Cd0TYGaqJJpTkxAuJAiO+vofUNIFE3O8kg
RUhBLEqSjYmvxOr/D4Pv/yxzAD5vGaX+kPf1Zp8TjADEL3xG7FRUxkXbeGUYQFh9
8Ych8ZLRvYaxkHja/nSuPX7NDKye/SFySERvk9jcV5VSPq85vP4vIfoPBGI5MGsv
z0KWCdj7RP7fLdOQew1vqVlC22BvJWisJNHhAFVrIegehgKinHJ4yO9a8DbvxWAX
76CPNznnCvtIJJMrVZVzL2cfqN6jGcn9H34wBMgrX2dC7rz1eAIfcHzUQw8Dduar
ZZdq4diVBMENj+S69z/t/OLsgG05Pfu+O24qDqA3LsrFlt/sQ3MbFDNZHp7nzaEM
YQ0k36DBYfvOSQxSq3LyXlYzEICGY6J7SHGL8oA73sOKFxwtoTWWaUew5Wuo+1iK
AWwzNu52utlsudX0g/f7qo3pz4RYzqvhbyLOrAEmokOCpiowFTXvkjK3DCCpVcec
7WGkwPu0M3XBNSH0jUgsUyMYCuFLcZjdI3caeekp+NSl1ARpYDlPvvr7azHpGHGF
552IuG1dLfFLISn1n71jMroJIer3Zel9Mnkd5EfCuhruV3h9gPjcu/BvOCzj2KAj
hd9zSKVv1Qk3JCm5Y2n2Zscom4LG1JhzSK5qSnTXwXBMZCebN0tn0/DRQwtcTOT5
YGVUkQ4jv7WMr3giM0fyeWzWkkF9XMHLATKhMqBidaP5D/TMhbGIaQblotR8tN+g
niuUv4kir31BR2Tx1db72PPLPSfKjHgLRu8gZhryhmUWVHa11OLMLiqzavaschWf
fBXI4f/G/XWqJ8a3LbVSMIQK8cEltRBDLz1rFMCw93q68u6lHYAfPTIkUTjLIaRq
TruHZY5oUWFDXiCdCmMR5wt012ywdJ5XdNNV0hKpvWkOcRxA/NqI2Bq/dNY0Tvvo
1dWnSa+x/2h4PCbqLGFi7sQcDygdUpaEv2g1W1E3C7ye1Lpqe02KVbAvAWrlBRbd
7RcDVJr0IJEj25oZ8gm7r9ls0MGAfeRdf/otBgW1hsb7ciJ9RT7GtZOKP+FaYYDT
4SxJBhxChbIQRO33Dxq/HRG316LcM8o2Md8IPxnJXBHQ/GzqFlwpg9Kq9+JYfR/h
N2H3M2136v8m9wPZ13+Y2BwSmfBSmQz2+M7zzdfummwEl8mGAgAlTSp4NCit/M2Y
jjMF+AeBsJQMdZTJ6zjzefcHlkCgusaLm2HJ7VQw/xf+5FNhcmYWy5y0qF/S5Sg9
KhSmnM9gjiBBnKgD1eyB9JqNrPLyvOSc8cvI0m+klzbx1ouqj3UlJXoAISlfs+Ij
2alT4bjE1K/cqz9LdkmangdazO9PjCWJyg/nDRbOcwYJS/x1vyGZqD1ENCy8zP02
KeMmQStsn1FGQNcCz0Y08SFVdiodHh0ciMlYd6VC0cqs89ZgahUWITe38dyBAUXX
kpjeaKzyePiBJO4aFQpaqWZOv87QJvvNXFd/JBJeUT795HR83bxei+6Xo5rK9R0M
e+i2Z76YZDSsG3CB+JXH7XRlvJWy/8lm0qZ3b2kH21pdaGL9pT8ZlvPS85mE1r1v
f0h0/2rMJh6y4ZjTfbu1IKR62++5s3fMoRTUyv7SoqWFHKvSfnue6iNLSpRoRSAK
UYudM8kaQQNb/U+sQCl+W4L9Iswxi2dx4/heBE4SDAdGYHFz4TlxP/l5IOoBnFmx
znZu1DZHSIUrrpv+HZ0m/b6xG94MVyxx4HN2XVKzXGegBVNx4KjRw/XF793ZPQSb
dELnDM8n157alA0Jfsqu7xe7YIEOXuW9QZMXMxqgt/iREioaa8Y/iCFmOecJIsJT
3i38sNJ/Zv52k7w48Pwn27nDAkNGD8DJdqNEKRAUXTOgb6p2Pqjg5HQ0oQ0q+4C0
ELgGssfd+vDZqrdwyzr1SWgQbzm5kGAuA/KN2QiLjH8=
`pragma protect end_protected
