// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:01 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k4EZiZBE7J9xw4fO+fbs8J66NGZRfVDxFUVZ3m4NFp6dohYy1sdBuTaA/8x/eObC
EqDxEceMHLQsHahnPRRNmveonXUhi0HtsG89RuvN48JlwAHLr5Q5DChCS0G1aa2L
r2fp+YwZQ7liNFOCPk3z79AYa6VtRygqdSdnN3HHq6k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28304)
IXsvVK5vIm4m5Pk53YxnT4sR3vP159S9+er2O59AuMQnurLeevGWqYB6xz1xZGRi
7aHyUFBEsgGoyTG1OeYP1NRt20ipNoQN655Jtgf+RvUDJwYuP29oWUQm0LEGE2Gs
0d9Khcz7XuUFEtkX2CMjsIzidk410hOhypIwWL5CoUSaTPYjouenjdzUZxg1zqTx
YK5vWj3K6JIlmgUYf883NrfQ5f6mhfPzpyAQysxhUaMyUs541+X094DA9pshN9sv
ZiOPqa6GgAJWwPQXel4vOrtv8tJOEYG/V/atNt99KEtaVwMtgzjDWAbJDDIPQYoh
WSsz6Tae9ZSAZnzpRgY8iWKgH6TE5DWTiC3qZZEeKmW6ytN83wfh390Wdn6Ekv/0
SnDNFXDXPXtFcl2zqBswEmLuc9Preax7elYen8y1aSo5MvqKt0wLr5gKBrb1NAaj
tftmI69UM6w9Lz5ZSozAeoNfeDkunaUAmmkgIYC1cT7rd60xRCo4ecpm0atv02ZT
tKqcIfurCe8ZYo2DUoiqZJFK1TyYOJAd9iPDzttsEi0QWlD9wAkU6CDNDSO/XFQ8
09RIuhkm0GP80iJYjyzIQoBgkMvRgUiN151LfXD79oDFl9KmwvJI6NLSSnMFZDks
AGmUKQeJlocOjQ4JnM9MkYewAB3WxixAx82RgQIFJFY+QvtBkrLjixWDX2YI1svw
R4nu2Jtb6b9Qaa4IPLH7lpCzEe0J7O/LWfBjJXVTT0fOB6TmOxMoEG1RM47IAHMb
BQSnf96cupxYuhUi4tZYBhJq6jZM16N/haUJI85kki0x/nGisS/6t2fmbQeYYZoR
yaXBJ+kMOKDf3pQ9833Fpz59jiIx+e0T6jnxbWPAAuef73bOjMzdPZyUowMwZDYB
qJRTgIdt/+6lJZwSiEOKluVgnf3itJK24KUQNE3YBQyDChhkAQelJH7D2sEOhHzu
RdCyKr9GJyaM2HTpCTdFuOriRnUUuTLmkjCkf32YNodESmnc3nYbjsPvCdo5MJ2L
BwB/WSxO2Lk1Z0PCJdWdYyLJfErBH3sEV09oGsADW+ZBljiDpXy0t8y26jK9Q7lY
X5kxGH0hAMXY09z1iEVgHYRVUtaQt4mCrHXSepmisMaLtN69BlIwuHZKjota3J0G
CC7IDDo5IUfckF25Czcph7Z9KUxta6mswSwegyZc7vOYhPYhseB1QcLhQal4t+4U
IFOsaFNGnuP5V4fZ+63nGDD0dhSey/aCJkI3KFQ9b2N1I4iTPvxpISOHrVDVlK6a
xOABlzC7TQ2paqhprIbbOO5DFztYGMA65Lsbw6zNxCF5/ls2iWpmSGWOL52NW5Mk
44Wxq+5mZ4E4EQM1oBFFBBNYgeHHO/FMxfaOJs3ta/lM2CFypfwbSkSodwudDn2M
zbh0ZvvpupX07MlGg5nII90EXTcwosAHwXGT7Xj38y7fwGTEOzN3tiRgBobQTZAr
dJFGKvwIjTHO7uUI9/B9Dj5VGF7QXFNFRwFJJifxvk6CKUOWWeKQc3NpubTchPEu
eBbOwemNaiU9Go7HKtj7OL1eO/MKiX8g1yHRdJV4ba31EsVN52VfEpX4AMn2b/OZ
cAlFOMFJ1P0eh1JFsd5MPCdfi5wWjnC+kHh6qCveFABRwaK16r/mxJWlkLxMiADS
fX8J+0qiTRsW1/pXBiFJ5dvlBoVrLtzwUPXLXXh3gZFQCcGHMnCIpQoW/WguYf7e
UsqspPHBfe1Rngw4NMgequjIfOpRdf+nFUbCfRZ9QRzYxxFd5IZ+5YU7tyj2p5vy
/1iyBzpj4z7XQoOFkOiGIvtAFpvSr3TITq4xavS3thPce4ie3D33wwirz3lkPtK3
R9FrcUe7CljbPDbO0F5rFa7aWHsi9MATu/JMYW6cpPNh0p7XoF/LHJXZz46Zw7/G
bcIea+V3dFH9/W3z1p8g37Q1JdTh4ne5DFxnsjT5uKuCqV8l7QFxMgCCyEuPmvEP
V2ofj1YxYEexglcO9kvZUmUOULkBDVWXYTJw88YefCGF5pi+yCpkJajRT4Om+ztp
DJzRPSNoK+5cIIv9dV8jfGxieFwOOnlcZBnx3BWulkNK5ga2fQhCF6jMUJWTXqUe
wvwZowGJSb7qUPVhxmEdOsD00zrWbFGjAo0A66MyDR2lHGz2spVHzGvNTAWtmCbk
ElrbAjLZQfQFwi1gRiNi4DBY61n0EgYxrTac9DzVEwv2YSY5YuHVF7T/4AA70iC9
FBLOl8E8L4kB/qPP0QUy0XPl3V0xG5+SkGyydPZ+Abo3TeRurBgIBjUSOHzvIzbE
0yApTHyV4ppHINXXEDYJJr6bTqVuw2TiQjZEvjWAT8BYJV+B8zWY07YWNsHHbJRl
0NQuccWjXQ70AZx50Bi4Mc0KgIfkWl07PnpJAXkBjRfrwJSIbrDx0w2LlcL1xxWm
M2vKu16tj4iJhaDY1yUu9zoojtXfRViUKQoM2RAYFD2+zRkskGegdeQYlTwN2bzZ
DF176nVx7hcWKyEp83YxYoa2hjaBQ/WeFXS7AaWEZkH20r/tR4xIm6b5/DGLb8V8
FyF6zqgSOiOyIsQ+yYx94MH6DgxHYGGtP5OmdcBfvhsZ7Xd1h/C2+9OgWms2xyuc
0DFpMNk6L+xyYHpK9nrE7thjzxBpjj/Jm5qLqeRvjSCuLIzsBkQcrKRKjjFwQhnc
lWPVyzD47TppvAiak51ij0y/Ln79L7C8pewc8hLhgHfolH9jjZc+nDIYrFDv0YG7
XgV2iqJpNSjpPFQGsZZ5GmoKtNEPYWGYR38CTDw/HuVbYXWOG9ZAjXF7zXhr694h
Fad9vY5FXh62KdhW42o5FwVOMioMIvqnSNdBK2b1mdciBgUOYXuRm1BykdcopADA
VgiUikoKWJqyAK155wdg8AEBmjgwOLGjxdg4+AMHcAEnrALCLZtuVbACPDs42vco
QaxMHlhB+axi3LsatyOHD/YmB+3wM0eQLldemRUaAEpCDlaPHpdNYXewWgvSAex+
wNZv36YFosybi0i5FER3qh9WcIAGQHt5tCufDyrWxM6YJM7fnMyrr+ayzRy9hs0j
EH3MOsfRj6rcVtJFWNm2a3ba9sJXwhqE1yHCAYJwI6DZOW69PO0kfjKVrO6XgEuh
HhbUr+JcKZ1gXzJivN6NfBYaq8gTLmUhSHhsrhsDp8vTqihhhcaXm0kOrBFg/UKg
8IUlT6rA/GroV6eZMepnmKS2JS6zmsSqhBvSFlTBRCZqU71rG9q/a1XNlsvCjYdB
QVWeo03csYSg72vGoYRFLq3Iv6jA9qV6DH83hcCQEUe8q94XgsIYpWefCekBjVfM
heaOodyAuR8t6D7k4ZMX6stHy2O7Q5iQk7ngSrmjhogATp1A2E9fkT9Ju0xtTMgw
JLEZX+xW3sC8pua1PkwWYpFxUCy8XdmDcI16gnzgSNINBhMLq5R92IRC/t7QMj56
RtWRhyWqAg1qQ81rBphITWShX5X1+Z6dMu3r50g5qxKbIYWKKIwR8ahWt49AENM5
ofCwAOrisME3ss9oeSr8ZBeCPTgz5WJuOOADekaaXEd3P4+g8mRi3VDiXAdcV8ei
xwFHCSfB1CpgXC3sjbfxXvzKUyM8BLPNJceQ1Z6IF51fRACHlHjhfzKBI8KIq3tU
IntpWItYdP8NVOg5dVSghzDRZSUmWu46njK4LzhD6nSR1fGSAlSbP584iC0J48IK
tviHClKQe7Z1yQOrfZhejZ2RTfPL9og61RpzWvTUDoe+RkIOopaa+RJl4SVBN40u
zQXkHmPjLEJaX87rj5XEbvgA9kBNwF2qCJxqgW1wCmmyNQqswrrZ0CMgzcy0QF0Y
NPPWKZ920myq52x0gYaLO1AD+Fw/twLwJP3aCAAMd6YCS9B9k3SU+Ur6cKGrg5oO
PoIaycUqrSpQ33qopEHKEHc3XGKyVint39yr6pLd/HRUXUXlULaGpXXSt8CHMcFb
GTw3iCwi+t+hXyetxkyfeFWPhBIxNRcRubCBdt0hSig+LhIMPMXDHC80QmYvCagg
AYRPb4kAjtUwESr4p1sLjucm3mJ+5oa1nWf/jDvo9LR0oV/Cb5jcEb5+Qz22XhFJ
aMSe9EPgl1H9JUsc4sEoHhaHXq6woFF4AnQbV4u9SrK1na7q2qR4F9o26Skya4W9
69hgyOTdgaZIuKIqH0u+jkO42DGtsZ73OdK8jqX+oOaEVbN58zToUEa5BVfqW/EJ
GVrbS1pk78c4GAA6DRp1bGfzD1GuWcp287yNIsrV/Y1ODOsWt7gtU/nu+6bD38cH
oIoWAWndc746z+OPWNB9UXT5iiaSvbEEfQTz9r93oBZZaMJfZJ6b87bLzxTokxcG
cEa6hGVeXFzeWOp/2l0F2CqbJ+2CsqpXEClT0lbFshc71pGJuJCmKBlFCrxTOxBX
hOXJEPv04YsQyYDHzeulSdTsDCJ2r46/2qKcSIOkXQ0YuIoN7Ui5sQNBKE0pZKsp
BZwVKfV1TSJ+17f5IepC/zaChF94kyFJqdw9QX8kb2Q6AqVUzgNP2Zft5/gz6sgF
imA99k94AvFk5QV+gXYFUfDvZ9dRX3gLS+bq+Diq80L9PO79OpxdQdgYZTEOrd7m
rlSK4VQfbtIXL9ysQDVFr5KKScdIQ8tMMWAKZKoUgp0FLeoYQoJkGonGQViULThz
eOdiFZ7KkE4LoTCe5gW84/gFs1l7OBzazYG7DIzqFY2PVX23vFH3UyivS6HnY5po
75dT6l3FlViGCF9UpDTKMJ7aHnTQ5gevCdXLWoM80dKRzpu9vtSCxT9z8X4zyY4Z
c5AOlyzxwI97Ctowvupo92uByXqCamV78F3kkPsrZ9f9c1CXYHw76O5POtZGIrGN
i+jMmGiCpfJONyStkFMyD+gtWEf7nIlfPZY/h06B2pkhia7t0Bvd64dO6UHCnopI
qKr2FtzsdBKkbVM1W5Nt7Xix/xfa1uskusOZaWPyEcefsYb2eAwYNx9rRjW8ze+D
aYMJV0pilIw685xh1Ztwz4HnbwxtezA+mXCd8fJYzYsGz8SrDltw+plOWJreHldp
MQLNwrvusyHIrD9eBv7BSpwwCcmFlPJT+CyUGo+eRMxX6Sjqns83gkrw1neo6y8I
eQFVYt8L+6+Xp9n5uQ+jurTKz/rGKS6wAayK+cnY5DbmujvqDR0na35fKeM6vTlr
P1qBMZZ6LoJTYSKlAxW4yGBhNS/bRVYPK0mqGyvT11+XSVoZeDFyuwKV4ZuEEoBQ
6J56Iy4P2zVQJpUC3ZDha656adY94GLAkFdBHUfb80ZpfOwYUusSYGuVukQlKJE9
f+4j3HshejKmUw3Kr2fe51sjhO/M1EhSzkJIJz/d4A8SBHV6G2vfNkNpb72loTmg
QbYWeB47EXDw3PxE+AxiC8VR6Bje8BpwxG/qsBQOb10gRYieIlEQ6fPmR33L1PuV
49agIduvwwb/bUQaAzIJNiPhwiVDTA8YUabRDAYEg2ktFokgaroanbi88zPt6GAJ
GGm2OVaDqCNMqG40r8uGYXjsLRBVkM8Fp2CCbo08EAGqc8cC/I9MKk6FsJ+wniEC
OWDDVvp9lhrcIj6I8ZOIlrVVkGFCkdgSg9AIve5JlGPiA4RYKBOfRPeZVeyOltct
fuVOXlUX+GirU/CxZEcIDNTRrJQGpwnld54sL5KukuZNIFY2M0goYIfp3+03BwfK
NEQ3X3WuLWUspaiWcDUGcwrKrIIcY+pJ7DkOFGLBlORIrNUMC3IjJNAMaXZHkGjI
p+0PjFn5mucNg0HYbYD0fLMqU13LgacNr84/mUIm1PKYhUX66N5DN7yt4vwBQP0K
prZVZb5bMgHJYY6y4ae8VjiUgF0hQK9+Vmf5yD16FWgL/kdjocxT8t0mXxgJkJ9H
OsoskpMmLp4/GmaBt+sF/HrHj+pPY9TZ1MaiilDQ5eLN2hceyTuBH8W5RurJvYIe
REomFw3CeVL3ys2GpM7llwAQnsXq5WUMiFPJZojUHr96G0sp9mYPfHvXpQmqnl2b
18pE5df2nRbQGhVHFeFz9Pr6jVBx3xhIGmYblfRPnEMoU5ChIdOEQWdYtBCTTX7r
IHhdpg/YW2Q7DURb3bJeyJqMao812D9skJc+s4eD8Qy9fRjauSAFdCIed734XQL7
PB6B1QLmyHXx1QhdmTwQ2Sq8do+WtWrftTphVLmqPvunMvr+YSJ8C0HKiHb8+S6V
p1fUssCyG19JBJAIj6AqzPQ/CJUhCI1NMCHgLPm+5etX2LVbrLO7Y6Wyp+QekgI8
kL07K76NpEZ5aI74DDqgZ/iU+tO9Rz5Mm3i8hCywCjcFUXrhG1cYPvgCbt2mCHUa
ZaU2ksGilWSNJnM+Sr2ihcJQW2BNSlgm0cNX5BKsAuiJU+UXKc83fWhFTDbnr8On
+rd50Qd1ouWKuoIMawzyi/Swa5T3m6leDCyr+ivgNuBgl3tumrGyOhqcLbgLLAVI
yJUrimTrGCqGEETz2yZko+/ryFlhyB7H/ay0m6sAksTK9rEkykx59KZPFd76znsN
HTGIHiIkQsWYsFhwUBUanoDkUf4Ctq121QVtKKrVgPaS4DeFAeJa/wajOLKPcMTN
uFCXqsbIklhNK+apS1GLocG4pU0eG6rM5xH1ESEXr0mPpXABBeVh7d3t1hYRADqA
LldrsRYRruLEcPTqOGz7P0Mfj3doHAeZvo+TXl5cQ1azv3p+Nq5z6/uEOkIj93DP
sLbZJkpxH3AQDJfrlevB/xvK6F1kLfmoQ7qWhw2zMfhe2mSSv7QHqHSGRdTZyMew
0RODJXfYpyqpAkZYsZOW0mxsYcil0PG+hq5N7SZvIcrdB864jMgPvbAT4eNGOp3u
5qv40dKsFNA/Gjam7iXxQZwIZxi+KVto9VzGfVaj9TBNeJanMvqcG2dVmjib4gGA
ChIyeOf2M5sHZ6pEEkrJxM8LlU3bBjyuqeeuf+xs7QKu5z+Dk6Whv+twJNUrIz9T
F5kn235np1dG3heyBJdEPhRaTudzDf8oFL+G52AsVE/TkjeoPwiq3t56wv7khqf9
UevKmYpkypExihYx3N0SJYAXTIFaJqvAErK3nmseDmNEhnP/g4SmtS9bAqrRuobu
o7ocF30yHwGgoyaO+ZdeRbQn5LmRy1gPxTSkjZG0smyaI4qrxheLeQm1gJdOr1aj
n9xKWJqBq30oUmaFXz5b3N8UG+KaBfZ2ApLxXkFEIPM6ksZ77ag2uDlQxqEgtPXh
IV4AEYnu6yzylTyFwpIGpiM1Q0CL8J01m2aoE8AaabDgFn0avm7zzZaxDSsyMn+C
CL28CmC2F9KaSK94ph2RFc6C/NDqY/BCjyTRL7JEFall8O5vli1/pTkaIDYvc96l
Jg25cdepxMiwbQEYUkKoKnea1fBRADBIwPsmGWciCQwxSiFSrCuCR7UiZ0yP4/2y
ZfwMRy5oWUjtnbuhoOpy+l2msbrLM7m5ISQMIOCrSaNta+JoeF8nHem8GsEI2SoN
1yhl+RJhmqjozr3tmq3Cl9I0z0VEtjaw3W0IXkT9po6nzY5OO++hcN2Ej5nPhC3r
2THaMBs4H4f6nV9xj79Av3Og6LJzmWkSe3E2va11Vsx3GIYmxT9U1VF2/TOC3gMS
Rj7VE+EBHxonLyEgbjKNYb4vLdy4haS8cUANFB9h09G7BmNa3RKS7dSH63qBILh1
bPpqGwou3lAr+UbfulITsvPxlzBbE2s+Ifo9F2Be24r2n/aj99U44oXtif5qL6zd
fJ7rTvUfyL45YmwRCNCqM3p9hM1nTAFL23sEDSD80hplITH3Aamb057A1w1X4Yn8
TvXZp+QznBA+l62tSYqhiw4RL+29uxP2qkHXMOSmbhsGFqHqzqdUk44XP4nmTeNR
8094Cwh1HmK2DW9St1Jq1YmYWmqrMd3Awtntam1mYbQC7nOANvjzcA7qQJGFtg2s
PePy8fkeI0fPTVNNM6CFho9Gv/VSBMYqFqkpFFBD1Her+cPN3esjS6D3EI24IOdl
11x9Kkjnfidx4r8lX0t1ZwDtTkACpADSuMOGfnJv1FBQ3bW1QOFUuMQmevRtK2kt
mL8STCvy/EEMB0/yqMPLQJUQ36jGHsXJxYVPCErO42c7n4k7tHY6rY7cjuAgAwj8
AdkOdqU1wSk77s6Wx1mGXtrfTCBbXH5bK9awZFUGTiqPcCMQ8OOs5/iI37tpjt3I
5HjByGmjZl5cBrf8nlYD4auh87/MjEbqUeI0Yc6vLIliQRCP8XW9+JXmnOLOdHwo
MkISv+F2tet655PMQHRIqIP00uVZPUxV6zyJiaxWxMAXVhyYi1B2VQ75mc0PiKVx
iVvrpCI6ByDmUFLnTiHNkbBZ4wYdX1ULN6NU4zbAyDrcZ7YKCcPMZW69rf6roM1p
y5UPPX7vgtEAvbuX8e33Ze1lRGkURnIPukqZg701wYIqLE3Gc9+NzKf9f3yS51bV
bh/mEQszU9yQdyGrD22yZ9tIrfnt+kqY9uiQ//hX6G6ZShnbezagQHYDxkG/gxoP
6dDM01viogX+i6HbN3vWVggXEhqPZfmkfdESmCJt+7rm5JOXnMZsWS7r6y0meaT2
OvugQoHAmITIaJCOHzQi+3K1Cj4y/CpnkVz/SJd9WnX31+kPO49wClAMmJknCXmG
eDrp3AAAB0fW9+LQKj8qifZl4sFK1ehVLbeItH+OGVPjEfLLzTqhsKACqqhzhrJe
ADcOTYzvBUqYSh7S8cd0GOKVDYCltz7CD5JqqKKdhtBFQdkxiXLC51R2SLMJ5e4d
p/f89SnY20xjIK+BaayFkEICKesPzHNBbFv/t1yv9DF9ybDhH856BYY0mABPW54D
7sqEtm/imp9zeiK6wZ1H0RlstS1MgwO5IROhJIY/Km0Ig0EaRmne87x/ZJwsrPuB
VMbzaO7torVosuI0LJvwiymBVzH+P5N0/gBedvpJ22vXdmLUX30CsC75qohje6XP
Zqco+00Eyn0rbTwYpL7HDFxni2tr1tQx+ZD0rFYQP4l/Jk5/1G2BHkPeD6HcajZU
/EFTVxpi/Gj0IRQTiUfGlsxTo9e4f7U+SZ1simTdZE5L2KLCroCv+20sLOPu1VIc
xKrMQs3OtIxJ2CWQgN2uAb3YQeEswB97bHWH4WfNIRNIEtLFM8E30x+hU0I8d++S
oZ+cRLZEVTUzrC4KddH384nr8AiDHCj1snrzBr9tL/5ZyhxZ6rVgelE54Afv5Se2
Znv3ouGdeXDfIV9v7TAwjYacHODrcB+JTULtaIFCubFPnms16tRoKW5Rfd4N2wLS
juGQfVoyLRpkmZrf4+aBJ2AXQvAph5eTcFKFNd0z6MCHaZyYGwhB9jSMgbXUQioe
1VJa0GgYAi+uATol8Uxg/SOiXN4X6WgUQh/r6u5prYcY7IsR0S1Ki5R2c5QV/bha
RYLJN4UEErNGBOodY1uo9NQppb83pAZnoWFBW2Mj0O5kQ0ado9ERPzX2oNuHqnOe
YWGZd8u3EWoFUTvu7zfJjdYfSeRXo43nMp8WMsT/nkyGatjjxryBRWoXleO25OdU
X0fyGJ6ZRyVWDArMVVylYvaTAFpXbf9Gh8Vo2npxdNOJYotbYJDTMZYHXJV7OMs/
Y+HBjxyguNCnEUFg7wQt9qJeygIqG6dSom9Wz0RA1KMg59lBbNVscZqHcvyQsP92
kMY4S51v1yoa6kjfbF0GF/HJVxD/Klv69FFMVEF1PKCay5IAitTSr3p3Ro/9Jpe1
8eY5IHueVo3DLS9oMS99W0vCYHDkjN28Twzf1Z0mq3VmLukojtL8hH0UAkH3YNk0
EYMpPc3JB0pmLxRtGEwEeqF8cOyo0ANyyDFMjC36I1DlXs+zTsj6DPzXCgwVXIXk
eMOMOKViQy9r4AM+3v/sm3VAiZOrBlz54PWx8IDKXh9y7A75iYVSXzrydAnNCXkj
FxceZDIIZGQZee1G5ZkIoMRgMhsDwIMcnEHF2poCy8ybhtaLZf6xanFEqt/Z65ep
JJNlxR0AjExoCuwrUE4ZRiOW8u/EsvkFnyhfQJ4stIjrJ3+wsXdafl5Opy07eQ0a
ub7tmJP2roPv4r+e1joW1KaONvcqeFdSl8i8ahFe+3/IObambdrZnKFByJaEHWoz
4J8JxSn+rh9fsVp8nOVWJRh748N7QayCJOTiy0fX3Mu6ljLoqOTAyv2l4fEIfNjK
62zewAtZrBzvBBI8mSMd8MZqETcibDO9CR/Lc2mxV+G8ogSizccTtlBJcKAcgYSz
+B+k79K8Y+bwYCs2ZSYRNB1J42pb/PIxHVQ2tS8oxFV2QlAwohPNid1kZyXDIHzC
7bpUXeb8/C3C9NLcoXsUYYWQmAxcp/RC9hCgjoTvPntxqztRiM3+pq+0HxCEgNVg
mz7vqwA9sitPNduv2vvnliUlk+HEarCPaNkDg0ivpXfR0ttXJnMCMVqNPeHirxjc
D4sk3qeFQvb5se+G7uvuk9aVUt4Yp4JlLbtG3VtB662davgSHOGsYQM/8NNCEEJd
vsJN7oTN8upIgoytcu1sXIZXaYEs0W9PEtSR9GtUF1knP+hPz8GkCOz53+ERqRJJ
0qmFA4SSXjdxtbrg70N1AG71P+0xcRQvDVVFzPXmTu/3xt+4sOwAVaoY4t8RRkvp
TIxQDK65b7k4FWFYZ/lOxoKGm07svQcBZ4z9LS1nYTpM71aMgRMtRVwRCkj3cN69
21UI5xB2TXp5EsPvLHJWmLVNZIgYAn4c1m/hwuEQirFGFLYdkgdbTyzvwGll6gLP
4AkaLcM8wVGI69kqA9dOsqeUp7DsfY6Jzq+pBpRE4r/EtKChC0j/iof0+Mm1wvnp
O9RQg3CijWCH7ePQmewAag04JtlTFggf8TvBCl+x0x7cZuJeGZ+fb2fx0ICiz0By
auekrJgum5AYsvGEilgRNoiVRYsR5yk+sSl7wm55C4Jo0Igx4gkIic3CA1o+F720
OBZArsCUIKFTmocQ7PtJjoykmuDieVMguiAYNsFt59d2RkuMnYm+xtLuJSGFpFc4
unkY3CR6Pf7MPc8HcMede8l+EeXOSDvH9+cApQoAjd0yEkfPHuzjEHUkiuoNz8QY
UwrRWEPDC3IdWfd1CaiG+MDqnwzlCdbYR3zBcbs2OaWRRHAN/wj4RrugBMq/BGuc
5MLiXUvmnmt7gHzu6Wvi4HLumcm4FeMQ6O/GDtgXD0XE+kWsNTN4rxmR9CjU87TL
U5CfALW8W5F5758MDhK00JhE2RjZ27WUTMVWlAOLdXjuiZKxAgitUcma/H13qYnc
DyLGXaT8n++8nAOJjs9iqvZXkRjDxnGSGmy9X77KP8gj79FxIT/AW8NbuJqhid0F
X9eM0PSR/4j8FUPlnG7RswVxdo28ckF8sAccJvtF2PBmwEa7sQTJHuqOpESaVVNp
IrVM7ZZmDd8WhNo8o6t2swK7jhl3Rea/NiZ/eWMHq/aArR2rQTzARd62YTcaw+1B
wjWQMkxiSWQZyGk2kIkoJ7S1KMwrwGgk83WcsAiW+dCZjbaVZ9C3io1NDV/M7bg4
QAqnDig6hgjEhyjK+nX9iToj+8DwD5iI9QpnTA8IhmHBH6Xd7DR3QBZxrTKrMYsL
8ppQ+IWFB2EIFaGaZnBNTDoSnzGoVFSuz/RjPIfjX1Mr9BT4FjvE5AzbgENh659g
fwwr9xz1i/HzPF8wvzIjQ3wROQVbFD4FJpw61jvOk79vTMz7Y0lEiGmg9vIOdT/t
n1C1E+U+R9oH6YdvRztndCBR4DAqG07Izq0f2EknsEuE1Y+Vt3XiNyw4FYGqlced
VVsz0itn+V+elcj/Ko6Yr/ILJvdLlXR7gtsLj5xf6UW6pYhzUxLvpsM99pDponeF
aLSrIDMrC6kBhZDcXOqDAA5EOnenK0S4Wl+r+EuxCE1yA9QHxmVwgWXUHBL82lMY
MaO29Iwhm2+r4Kx08BhLFoQ0pkN0xd7RDH4nyw+3dgqK7xBstASI13uC4PAPNz9d
vvo4n8fITk+dFTIryQO73ne25CQXvTFtd36CcEL+XNxRBFjCi5yzWGxg9ZRxlOgF
sGVl7yMU9HXcTf2rB3zZ56SfWyL7DLZothzP2wmXICfH/D8ScEh1UNSNC9tTi+Bf
7ARNVIeOfpMTd1ztkO5LSjJOG97rrmpSbNxM4W36p2McfWXeRj30BnLs43hQc9yD
17AWlQ/7Ub3ciU1I8ws0K3Ptpr9dYKntifx+Tp5yjETD9JTLaCoj0s5o3l4AsulL
KOm3OfJWOiqBWLst7Jn0ogZdqIBT+WonMqneRwBGnSh88Dx1IRayQbkF33mXrvOC
AKZJVeyc6b6621MdkCdTFHnIbTUxhObgjZsF1ZEd0k/wBZoSgygbsz4ggrN6ihbG
8g+5hmrB3YMWwJo5YJ/cKLf1p7rrSd87u6gDZp5wJWTX8Pb3zN98b+hifP+5raNl
w98Wpno3f1X+6wG0PxH90f9/RfvXMQpGxCSlGqdDe7nUzS6u0TJieO93IIKTQ2lQ
N9tiMW6/obhTiOxy17bxDnGY5kFmuaMUUfmC3a7ynBDe0IIQm5vyUrUdTygPjNGK
L515PAkoj5BZRQI4zCnSxMGaRAl+VHqJLKtp10gqtn+kXXsnaiY2I/BGySzmpUCG
kpkXMuMiIZASWXpXe1P/+3FNex/WrIxMWrmuGPk+fP145hRDTr3xG3bqo4h3zQvH
55cHHGfOvRwPiq+bxhzqqIGjARAps+RWfTdM8JpivHd/gi1ZY3b1BAON8czfI2+R
cGjU680WrL6yV4N44Qyk6PdDhwA11lROuJ3dnlTBtmJTh5VoqqD1zaly6EZE1pCv
5+V7oucjlfivLLxxLml3kGu1y0uVikZXy3pgrQmRZyQU7ZVudexJTRsbGSr5qDJU
ZyZQ6w5b3y+K0Q9QKv29PC7kXRU3QhDbDFn+D++aHohppkC8VPUKAYlJuXGxOun1
iYBgZSUX44bevhE5KUnfbo37XHtLDrjjjrvqCE6rW8vaUfsBSjP2qlr7m0NukktJ
BefCUf7NlqFjJXjA5OaIKn45KK+cix2xGIfCoFF02tyJlfCgQVWc8XgaWYPibtY8
PjtsiygvjbB15PbPkfMFXu7lqRHxYaqRk9r1ts+FfE7aCEMrpMJguL5lP85FS9MX
9f539CcxzRkN/VLKsCk07MV760HgTHXLbTpF3VvuLCE7kICzeurfxBXRhnCrdhhq
UPeXkHyysSkFD0eaDGrBrt02Deg6lb7xtVKc45cnJeIzZHNLiaMzdLouY3wEoqLH
DzFKPt9du/vP8+rwL68g1kCtjUr/9kR2vWKbS8YwSW0ydvHEaIkA1GaQt5q9Zf7o
peaL24NQGU0wmIAvfi45NNssTBhtLT6ZtWfapPjMBnowuP3AxyPRNGI0UMpWlG46
3Ud5ewgGui4Fqlid8txMttvIEzYAj7svxsg6HyaVVsUVwrb/DqFjitIJfmwAAm9E
8slGENGJP5Up2COEzId78efCZ3uzSt75YgGDM1pEm8I2Kpv36trIa9kZdML2UB+2
73vX2eH8WBevS7uW4fGSI64wb1bOk4GWfJlbOz6mJc513RdOG+n6AAQyZKB4S0bS
Oym89cvO0wyBFqn/p2DEXenfI9UHGohNgkeoTPJA2qJNz3jSYP/fybqLLDHfFUNo
05Gz6SUtiMu4hYNoj9hb5dKqib8AOc4ktcG5r1m4Dm16YTmjq3Fy9wCe3PqyHd3L
YTxdvw4juNvjIRuQgcOMgZUv2kr7W/63lSW0ojQQ+59Ejn2bUY6xF2Kgadja6jiL
3mJXYO2DAgW7SR0jl/pOg72UN305Hoj0xVl4zsxM4gJ6ngX9R+wPsxBgdrUis4B3
kVh+pNyGXAsMQMzpTtccQC1L0bWOf3cZ+yp4dKdVtdLNLqkvudlmLlFMCLu84PeE
BBn21F+s4eTdn4HdrLD0mpd99esperukBcSpLZdXtfRHLaOKvYrf7Uw0ZHtpJdIM
+FSk9SMycBRzThMx+DglW7407gEwqyvhQTH7aX5hCfhlh/8dXQimEXIqm1Zmso8c
ripAvVwZ7a7U0VWvzrIZRS+HWYxEc5uJ/Eio73RJHF8+BUtvou2l8S+FRx0raodF
akJowei7ovBYfwfxNwCFIEC3jRL2pnLBLD20bpF4aKiJnJAlP9ob9B/7dazLuo9F
Mwd+sZizfrDnV22hNM7n/vvtoF1lVO6irlhBkrvmVcT8KRWFZzYpuvkfGFi4HQ4g
kTTYsQRSqM0OO1NMV/m4zjkDG2yaa/vl1PCKN+ItB+xEGGwvyS5Zq/ZR92e9ZgW5
hadYB79r3jbLglk+M1wZhaaLJV8jrui2QObkvZ68oHKk2wbTXhGgvjhzFW+JgKzj
Q0oYME6FsPZIYl2vNigFVEStSVPh8u8cWuUqj1QnmimRRAesv7cEuIs5veD4cH5u
hVX9IojKgmmypHtRyeLcyGIjG6nyoWy4bDDSdhX/0e1yKPwlyqbPNNVZ6cSFY0G8
E53luxUGnNnt8k6PFH2yvjR3q4Y+hWqdnhe27i5NYnJTM2PeNI87I257/6945PMw
OdQ5SeVSu3lGT4oDLR5KpwF51tnpLK5fxXv+v/yDPfZvILcpvWxi9POJJP5ApCL1
ZuObpUQdUXi6OuojN7c/AA9bROgwGoycquz2wpJWGyLDIHWvt8337fgivIal/l0x
zH5bMSiVmc3egBuY7s793F8JwvHkjAkE4sf/HHDdbq6QcU3j3kOOt0uSj2ziTXQg
PWGhBHE6xZX1oo4/mbyOs45UBpnr1y2eYjasVt5Y2sexOEOwXWRPs72Y8sNkQNGn
gH30zrt8CdWNYgCT4MMdlgwqIO2FVdsmFSspVza8bmp2A+Xw76z+mcWyBLL1yApc
nQNsjyCIoGQ1Y0W+nwMHUK3gO7EmPteweyM07qTPJgyjY8TIF0Clmco9cMoRMIBp
mOmdW3re2P9jaBrUXb7U7VdhErApMHKf6u2TkciAeVJXipBwVRbzO5QxnxpJfZV+
aAw+WSeNoKvB4BSP2AhKyu1x49hr/H8sDIuq9no8PXIqhQY+AaGLkn+mPiXybq6R
BsvCibscsSx45J70vWXd+soEHj911CDG9JXXRNMSsJ2XePxSff+ZNEmoa3n91cyl
JIJkHdo1/ot61bqZ3OiDKQV5MVkaNKck59OnynwYBPGk7bdyfLZ76zBUagqBlRql
jABCv2CCb/po5Wn0i0GCtQSgrkmdfMjd7OG0SCoenrcdFuu5xBx9BX7LKkgZwZ4u
vdszBPHqkJHQL9a0D6XXlRetDGE6Bc+sVPQASmL6yt3azbZocDQqP1RuVeNnOjjb
Ec2ZyY6hO4F9hPlsCy97lPpI1OeCayzMY3eOOXlg4zBRMdMW88onCTvweMmOtbUj
6UnBtGlGITN9GE1t97LGBOC+093WQZQLHMWVEYTY+1/+69eXBp8Gxp9AQHZJbmkL
Ytkx5N662RoEvRXzrXzvpW+jQAQI8a3RLNyl4zgA997AMIJAeGq/rp2NzUu+C5GS
kxlqBWWJlsnQlUQ4CzV9L9A9xpQJ0EDEMx7lr8icYnGSgIQRDSIkDvkXPrjIygzD
uFelDTyi1MvnoqhAKO2VxXDxdsvhW4URd9mgQqAn1ZsPIBnE1IBSMIhRVZX74KK7
rMXGT9UlnZsjaubmFIcDGBt3t/bUuO52N6NGILPyzYvbompf8TkYjHV2DzWu0VOV
+2ZfvgvXhMgRUv+zOJxHBx5jubi1hNxY1gxujOr/wFhi08LEUtnnz56CGjHUSrAh
svIJQcZYzOJKdWfoa4xM3eAaPLhlKHAC1AD9sJJ9AV4mA/ZweWy4HYZBuWCR7PiP
sLgZd5vfYQn97oiVs9SrmehRrmoyNSCq/V9Imjlsw155CWntk6NzRHiB4cVv+W6A
hmrQWYxGixYsN6FCPQrtlo0E2KTSrAP0/wRpVC8W59fRWr/TxCwMRznk/Qz4ZmGK
B5lOnKVEb2cMtlDD+DDQkRe+o74ivTD/QOmIsXTKlktZ7FtyGKlYJZqDy9n+BR9Z
p3WRN0XnPCXxsHU+Dmq4rLbKTR4YfNimDZuavnij+9IVHQiQWj6wVLWBHw7Hq2vd
w3E04hJqQ73HdCjQ1A3MILLEO9BxYVR5JVa2XK6j1PuGmKQ6pxZlnAALf3DmBp2O
xd5FjGC2HlEEwBQg/RFNGLepi7U3qD2SCAS20KdmyrKV54epl/FjBXKTnzHardAf
1H0XaI4dk9KKs5wJ2QiGk5Jp34SVi3JVVFek15C44CKOcfbIXdeGG3pNWwZU9kgN
5nbNrOI+2R82bu/u0Lt10JtwdCIv/kde017BQ0xX6U8z4e+Fn1Fv1xX1lEXcv8bQ
kPVc4Ltq8ZCllD2c6xJTrmk5sPbCdsPcklqsCWPE1c+yN4SLB+cK9buNB1k41LO4
3LlGa38VA81nl0Ev9UGtCkZViAhqnzOdQUOoPuHaFW+iuVPuM0Fx0XcKsoMoqCMn
O/qHhDoVv7fhnVCFNMalLHENWuyWwgWcbhKjGvQrcyMPxrYvJdPgfbECKHBcW/5q
6kdu04zOT3BJVYlPzBZRusVGgYRw3J8vlYacCQSzgRp2Knc5D+mTj34OExtpTy4w
du62h7POjDJ1MYaflnYozVxfJnQcs5OOAkfCYHvXNIGWqxMnQb/pfqFUlhE9OSnJ
XklXB7cXXtTCmwH1CuPbeYq0O5TX8ZCIMyTUCqYwHepxfyrXgfox4wvXpzi0RfoB
OdJfqHu5dlKSSjDq962r3b8UhLI7DBkyFpDPOI54SQPMJlyMcHeOYCChqnHA8XvT
xSJoJ3IcnhK21bIpFlTBmsw1JXXhtGobE9Cvvl1tpMP06DA502kyCfcPWcd+YZ7P
aL2+Yl1Pbv5XS5h2LtkyJxZFZu3agBu3Ye2Ni3erfljKyeX6in88nrzZsjODrVDK
wjdJqSSQAgf7O6bR+4yTfzsIIuRLepSYraN916FNU5oP8akFpuKKF2dmA4bY09PQ
5S8MuKzlwInXxE0hAiLHHYPkTY1rEJ32m0zbhVmRBDOuT8opxYsSukjHyi+Rauko
c7ZDXYfcrXCnDprEhpkh4mChqQBy825HEcnZ2A0hm75T+MNEIf5ySYTWopz7X3Ga
YtEmhNUbMdYl4cQJDbyC1OOlfJxcMlOR1OFuzPPDxOhdC4iLyzejf18pjAHzpR9S
QrRKoq9SFzVO2Jeog0Z3vkGIDI3EuTVWfkKDmDN0hvd752m1STLQ+S7yovIkSILy
9YCh97DKs+pKJaLcS8BYAYwFjNmDQpgXjRg+MabS29IfiEuAza8cX6fbTRoyMpW4
MTjLBnO7NqNsSvxiHVpIKtN5zv74OZf3pihWM8KPp/XBDJfFjbI2TAJWF9Jq8PVn
d1+AHAtKHbBcpdBiLXLKVucwMZmiWoiJKsmWGdQQlaZum+QlvRJeqEdpb/xTzUwZ
i7G6cs2WGowgiE0MhIvosRmgkY3iOHl/nTgztSO5/QMW+OPEM7hrti9qgO+Y2dvf
V3UWT2+EDaMq10mSTh3HO08gbdtyL6Us72oBzwyOZ9gjtf8bYW4A/A8/uBFExQo/
RwtJgD9CTEdo0tn1Uuyngorb274tqb2cL+65oPBZxc6k09Dw15Qx6ayHmuirBLdp
aEXd2OJ7QJj7ZEeGoAKPEajxNoX4RCfRe3kESKsLZ8DKAmN5ACz0hB/53d4hRp59
wIrE7C6Ub024mkDPgzxPrQOhseBVLFdf9aJ6NPPeS7Hi7naff/mqqlGiiTl9eYeR
vX7NQzcdSBvfXFO10bLjenhhmH2OiMG2rn7biNUH67QeegWnlqiB8YwrXbeH8+HV
sTumZF3ApoWRUi1EniEm24jvK9eJUuYsQVLT63ni2V8+vLZlSP30YpLOBuqwKpXu
batImaCs4pe+A6epG9OiioTeOXsKOrLRyDmjlQOkT7cbA1lCYxMO77PQVNkbdBM4
BIut9nVnmFyaUdUwxxQNMby/lkreidr6fzgMiNxForn5bzqr5dTwyZm8ct5pHkg5
MclOD0P69fA4UULAFdcb7M6kqgYzK/RoTDLZ1T2ha49apdOho6kXE+FrsrNCkc+U
2q9ZZR1+eyjbYFo9N3qSnh7JInjFeT4tjEDW7iessIe68DVsrPl3loE5WHkj96dI
6X1s1N1eASLK8GAPSsEKYdnkknd47HW8KDS2JrSA/bUQPKBooBT60M0U7Ti3/n+d
EszRzqATQBhGmB8HlK6j4XOzeUW3dYHs//E5V/vcT7PhxNAFw+OhCSaNwI0csya7
M1WCqrtNfxJKhkJDd5xWywAMATkmOSoFAKenS6r72ttrJb3UJFecB0FR+0IiZRgq
YPZ4CBtHwipYxu+l3rCUUGyA59MCiY1FNwnGFFY1zPudAYIS6o+viJV9xneRP/Ib
bdOM9NwAz1pXcs8GsbyzLPihT/QEaHKfYWvMK/5/QIBkMOe0gptUKJAYVvo2fUi7
u5OiZ2pn4bjls4BMXzs2PPSBK2PiyEZxnDfZ8mRmiagEaXhTyS3SOAwuFsbXXNKe
RSt91uO+1yKFwG6BAQw1XRK0tBdL3jkudaYlXXOKg8TOKw+DIC+Xh/zNKfQs/HjF
VZo4t7qNcFR7SgYAoafVnW3j9JW/jrWItgJZ4TFW21sCFRfBY9Q+cWyaNMyP6ru/
GUTpNHF44KkiapqzzEk8jYzohmSlZ07oFAIdKHJImvien2vsU9M0LkY7FIry3CPm
3fRuv4AOaNEDGVUgp/JzddHWOX0qcBPeBGUxc+4Fes06h3qqzhYkI/qqnWHpVp0R
kNPPEig2JjH6DVHN/zBwwoLTOmJG/fa1EyltydcBSrjpdUekAEWC8AXjFOHYWtdJ
G4fS8sst9FCmTUci5lU+whdN1wTZTseIL7gf4GzdomrbT1pI14+8lWdiqa+ZxJ8/
RMSsJb5j9dWbxEmnXtQjes0I43ZrZxHWSkIao+RGJLzCRH2L1v9G8ggiIjok2K+B
9ee/ac6Tu2gqRhSlRGHQBc9DollfD3MHe2T3MXRGgNLsdPn2TpeS+ajM4NEwUVDd
gX5OcFggi6TsysGdqJi0Sa4G6MVUNz73tfNkFNHqi5Dx8JOQJc53aOM/RGiD/sQC
6SlOKBY4j9tkalBYt/hCSNcn/xQR8V+sgvQzX9i8yS0kF3r3kJoAcuYVJe5j5gTS
TYUdKrRGfyPFuGrjv4/76LR8y3eCjn4eb3C9K0q209APya3gXuMBA8VZHDUZM01K
wxrveqPzoS9UXLyfXSDlenuAABDpYfwlf2LF48UOVscmNH6hcCA0nn0uxmdo+qhH
i3mRNq1jR12HH+2vzq2Q+HtKYW/MEjAhlz3OjSldyoNgfAX4C+xkMF7/L0qq4aTf
NEtJIHYHxNZO5DkCdcwr3DVd+3OKMxaq6WlOeGB4t0pQF91fjquxqkY0UKtfonb1
5IVm81wQUNckJB6990LT8vzNrm8kzeHYIvIepgaBn4sHzr/pM3En3mIjl8UvrRLZ
v42yK753MkdiyG1Yq2MKNWfvyPBug62gL7YlaS6O4lpSlYrcXADrJfh4DNjHfvru
d5jJ/P6/8MbrGJDB5mySAncWyp0QOa4lS8eKA5ieyzyYUX8hjvwE0jQdMsKcarOI
cD3U0hSUj4jz290w0ktjVlGLHothguZ/yZtja/e5SfeyUqGGtIXV+j3ET1y9Rnkx
ff+reQm6jbo4wcjzhJdRDdkGxPLpRd8e/t1knQumgFjv3O3VVxuEI8IbIZ+bLkqy
zb5ZASeJ53D0hSeH6Vy9ZoLnzxCyFcVOLOLBmN7/TvfX0V22ygavG7NOBcYoxRFq
1Y1oLm/G4zIQmctWYiKkQurRshp4/Nln1ZiJmyMOSKFEPvRIt0gH9ZwjehP5CvYx
M0myNeVueR8GuDz5MOttYw6TB7cdqiefT+8eiBn9JDa0oC+tviQjzzl6RrEHKIna
Y5v+6X7aW6R9ZwaPzCHxN+N/epdX0FNl1dAdVQdgpeD4eSAfFW023/Y/95SKAXGt
fC9XnLLmLU62fe/I2mGBToBCTUfzUKMlt1QvjjNmxnbyNrEd75ZPWLJESEK35uWJ
CTsoGixdWhSGKKq/o+8VHJmmm/+PcoW7Q3G5HUGTUcj/v4iKnqJxF+abTym9rdaS
97/2t+/FvM561L62H6H2Obhd/dXuJ2BTBvaf3tYbpe1VaxjPl9rNBGm7HT1K7x7y
kRGyorlzOqbGoauMSgfBjwpc6iA1zGm2LaS7QaSnA2yFBKTMrAry+m9r2xnqPGcF
WBgrKR4jzXnzwMCPQvNyEuZXXjdbYCyaajMMU2RhrtBAfD/t8mq4H2TK3ne5o5p1
gIOIBcpiSrNg6iJk1PhM/5H+GgeaBV3hyX2r0tb91lrbbo465HCDM8MgHH5FZAVi
epGp6fIH9ZjrRTfaccmZYkRUJ/u4/+95vY+RFlk5ktKV//n3ggTMOYyYRJEjP9rl
INJ7Kb+T8EEWwY4ufVBjvcszxC/KQpK6rxsnkyDGV7E38a/JOX0YjKmjIFSHoWnz
ehI8qwU+vFBJgPBwARCm+WWYmhNYumVWvJh+0pMcKGJydRk24aB7Oa9/fqapJuTZ
Z2WO0qaD/kT2Myw09o0AFKW9CpxAnGMIjh5F/Y86owFIbYvfdB9ETB1g/M69RYPk
c9DE4MZI1pMDEPJNi3MVZXy1Nq8kkKTYSO+F6Iixk9ANetfTcmUxd/7STX45ss8J
TNgzXe8vG8bYbj7bD7LlH1K0YJlbHhF515ou463sSoAEEgr9j7RShcaBNGPHOYjK
qzMBOCG9nlGCC/q/Kp8TgQDaJ26rgP7a3uXA2+5UlSVCv1oxtsGoRcWmIYcRo+po
Xee+5DtFr986+z0OCP5ZVVDH3wm+u7QJ0EZxkUcbaHJ/5wBIhI680Q87zvVFnyAy
g4Mul3kDDH/8dMvmiOhX0NMv9YlhTYvvmjcCSUqmk1En3GfTBamU22UNql1ktmMh
q7zMhSClJa0PDnUuQ53qjGDy7XegfR4K08LuSZWO5Y/DWAOZROm5C0KqcevyerBH
0vLsRYQsCeL0lTkZzCPjgeUMi/O4LNYfHoC5fgXqQxFx3AvCgrp646IIcRF2L2Df
nTaqIYlP3c356qM9TarGIF3ORzJc59L1dOLEnEvxIXJYyAdvC5ycJtUcUyq0P5YD
i26UO2OSVp035Qfx3j873/E9PrOYCXzwBlLefGsb0+xLUOi6+9ieP3rZym2UgylO
9xsA6NZnLBazANSP0ZD7jbHscn5oxfbWG6znCWIk+HfYwrcfZcVp12/P5eFBniA5
q5lJJCnmUZ20ibaAqy5pSyB9XzKx8PB3F2AR+xmzmYb1ljf3ZCCo0ymBEqUHVR3A
zSPBZvN/BILSeFscTlshesle0Qjz119pGcS6TifEJdEG+n+IWKA/TljCPbc1zceT
/xtjWkhGrKNYQdmO7r4gbOTLb7b5NNEJ6c20mq35he0pQ1+eUZiK9r2yuNFRV0La
FYFYXNq00AVLsfwiAxgZByrQTo2o3NYyp1XzhpOQgj3RRE6lyj9o18ZeuxuU56Kq
eh9G/jyaA4GOEYLlBFTiPtYjLUkn9lPaoVPbMxud7jgFYXeGmDHnbMkAa2HCCWp7
mZbZJS6bRXs9++6aNPg3l1iwbfJ8gAZ7JXJLQEM1Ba0+SZOIScKKa8G5HlWCFcij
+69bKcXAQNaoIj+Kn7XFInId3nLZWgXTUgHDdnx81aG/B7CFjk/sesu/TSCc86SL
nxNafl2rkrQCQSFDpQy4o7FngoKPVVsw8MRDzWdFfYL5KJuIhnYrgfJl7Q/qOtAb
cly5OIFHRaGufucVaenZTFkjprY+MQQTy2LgzYaaRvTohwcAJENdasjFDDy1Mhx7
nQqak3ZHxBo5tw1wpL4TWudWdUEx1SeDdVYVz3TlKioVBXElTD36kJNXrRNA8hMQ
6sgofpBExST2fHs28y01UZAwYwsqmPKvvJc6qA4sqGAnBg2YGslapiixd+kZPSOH
LW/EYSWiaZtS5mdQ9l1/TcijoehB7sdIbdw5z/FoJaMl3yYTEq+FHTg/lkeRt2Io
cERmKdlZB/nryG7Q4H0l9YCdHDK7rhSJ3Su5w5DqexFS/QQTiTsaMZyuic9NvbGR
zSyrq6/SzmZK43JXN4b6/N9Cr4ih7W0WTPhSZdsOADOpYk1cVUVKufilw7L6zBNN
Us7WNdRpbQGCetmY+qoO3g0jjp6iYYSb7XkGO0peg2V9Jn/Un3m1JeMmLnd89dt4
ZjmqvOkuy5b87BZfL2w5kbJJcdc8QH996g5ZAPBvmPSU+ZLYxDhQ5D20EbpIGSqH
2J+6jia6Pi9kpKufoki0KR5So1RxGv5nR/bD2J1R3V/0UuMbAnMBlcVpE/VyvuGr
PISp3M8hHhXwSRK4pnxnCxC2lEMZ3hqhHPcDV099ki2Z/EOS+3/p0EhhaP/Xfl3g
SM1uXxbDvxBw3Ms/8X43ipgTgoFDNiiDFArkkOi6uq8siX89WGS1lTVLkoMEJrpv
DSS4AsyFx3wbGceyUjXq8xiKgeObNiiAnz1KFQtJ+3JUXEwjWDcxOqH79qQz0EJb
PWprauzC50HOyXMrrfh/WFs4VgNjM0mD96N29Xu0rHvh4jQbe+tmRJkEFMEk7O7R
FCIVRme27YRawjT2wqAvxkw67jf5E9XFnAxe6mqynq95rKsTjiYcPsZ4WkNsCB1h
QfKpo2zwpqDrRf6zhUKEF/STxCbm0Hu+2o1ho+XWS9QiDcQoyJpqPECdvI3+yXTB
ZE80F1u49gkg/G6+GjpdWwxp0pu6KPyNy+tD4rWxNzFEo/t1N7On0Xi1d8+W9Lk1
8jktRBVTQcPv8xXh3yMP4KrychIrYBz++u1DkSmmtgNHhP7v8ucVWKHlAKoOni5d
QB0umPPkIgE4Fa4+EM6LBQfJwZ1SzDxeE926gw2mpUlwFgVsUMCuzbZ8bvoMDsGO
aEfWhVencXk4fcIkcyfHjILGBee2xwSGRlmJQrpx3Dr1qrvXfpnZMk61u1u0W2oz
8I1SBO8XrDXeo78d8VR8dKp5qJwoZ5ej5r+VwobVy2vIedmsc7HrDOY//GcBVIIO
7GO9+FyOHW7/AiqC9NFypIVo0XyqWpsfRbqqXKu/A+06Y2+CXmJ+vak8z5PXJrkB
+4D5F5pT8NEZP04ZRcGFDaoybDq+cYdCKBQ8gS3aHYeE1H1sv0naEnJo/OxHMQF4
sP4oQiYglfD1G5FAcN0G1f/Hx3pDQ4ohuIQk3a0MOmiaHM4ZgXIHLowSsiEEiTdu
zq/SK2yy4vFCt+it8Kd37l9WbuqjAo5pSqixw9Ujd9lkPTavsMbunjfzKrxURjvU
PDKwA6+NV0yJ5qBdmzD0TlZHV2qLgY/2nfcpjS8a1W/NSH42O7T3Zn3qbONu4CS8
Lx8ms+rbuVJkzpe64QfWQDkOpUgj+uezPFZ9jjW4WYEAzXEW0EcylMxwO2WmNp4T
jQH+dTdzqwKmf1tstre5g/Bc23bdCXk2ZOt/yLuvXb3u4vuzenSRKu3Jk5SHsi+e
6r3/dy8HLzNQJGEG58/s2/So9gwCIgtqGlXFFUU/uuzCKNW0tQDCltEjNXl6ThvH
0Y0087p8pD9JGEE7LVBERKMzCktPA6oevrp119htYMVehNDjz0WKXoXWaqW4qXCp
WuhbdGu6mJqwnGVWvfNS1jCewNKCMG/QtchY7UEl1hL9eYPzUPDkykgZayA908tU
s9R29zBiIhoKSV+CoGQJWIv6oFCintU8aGZdp3kA3bFKc+cK0fEPfOrOU/LbIkGt
zZQbBW+tNmTD96xHoRk8O6EZ9/5+8DyGWG5ODHbuE0g3w98ExWovWFyhrWHTb1D5
XbWuQWfcDNu/Gdlt0RfK9n0cWVZQbk69chz2zqr4zha0zmhVT7ZRjaxgmqiDCXS7
YMaKRNY46P+abUVct449ElEQqpAEeprIwWYA9+gBxaggEzUosDOv9DynN2c9TJyR
cyKeE7eOiuACDpMoZUPCEisPYxkCpIY4aYeEW7j0DszqSykTPhSzvySnf/QEqbPW
b4uXTVRFXaJ/1itvWZEJ97L487LoAiX2Iusmz4w2VVusAF08VGONIaeDzzh8Iy6Q
wPWGf8AQNLXrYmVLH8ryLWcsySfE3mORDN+eQ+s5ECjs04h3AaaQ+jS2K4cSBhqO
XA7BG1kHclyA73CzBdp7qxlYrsEtvdUX2QfXEuahQZhg4vvWU//ZiPm2W7HxUsPC
lVTLti+eehGljZPU+d7PBfVDgOLxY16dZwxEvzj0iRhEE6pDJfFrftazi9iPo0T7
+/v8m642TIq7UfpvI3UUSXF836kwtUsz4Hczi8KGKPG9YAd20D+pC4uyefFbm/Ot
OYSglxGMAbBEVBRsQbioicA5Gb3vmtQcfzhgnuxet0uucJ8A/yjQ+udMYam2bl/k
wmdL6ZdAIhZcL9WHZ0vb2VnmT4Mu7nqWef52Kc2v81Bnmt1Xh6eYbZduF7iwjbuA
yehWOj26AfmdyhVlBhzQ0Nv4ouyTxP/gHDA64e/YT1yfW6Fx654/CKS7fKrg7nCr
TMCl5m3iDV8oIPBc6fg/hNXPPsVZszzha17YullIw6CTtL9qgQ1nNWFRbdX2Yjt6
boDNBJz54Qp579XIfJhhUMrw1KsutRXNfC0oeVzrRSSwIsIYbK3RX4zHAd5fmCUY
wqHqqmZr3viRR8b/7I1561pBM30ktgzKTmQJIYlmBMXgQguVKFHB8G7+pux8K0kn
oh+oLItqFHQkAefTmnPnjKrxcbAJbMIs0M23JzuV+rKpv0A478X8Ke8KRB+28TEW
l/NbmyrXFLgQtguJX4u9MEwln6zuabchEQ2M3lPn/QJ89moE+LTFic8In3RWKYEQ
osFWEM3LcwRase+LLRygCrEb31kEFmpVPXC5a+Aol9WBJEWh+vewh90toKXkUBZC
V8CMmvEbF2gyKfd6Oa3pLWyb67gZwO3TvC4xm0GpiQk78gd4jBHrRppyHXfVjCvh
96NBHC2obEnSQ92S5PJOG/F8jwRSlpirC8L1rrUALt+1Ztiwsn1YIn4T8e5eUTJR
lE38ZLfGnpEeASAe/sE+4ijQxGweLA3ympUXI+dDeE2uIxxelyMr0qKhHklVHLuG
KfWMUG5N4zCWZeXRrB7WFdaH/aMIg57KT6MvKphBWwUKDqzLKGYS6KOW9qasdoun
f+i+AMcunmK/lCGpHHYkebgSq0fnKbgCwv2LlZY7aG3RkCy9WyP5xXiJotMpjoKg
2L8UPbiRu72wVp9DWVYHbLF+ZZJxv585XjdZd5E+tCf1DRzQkHTka7H/8enUo+WE
6af4L31YENLmp1lB/LMRUCpCRASZcbZA5uGYUInb6UxTiSuTNNH7J3gGIUdapfpI
eiFGkx2ls/wWQy6hkrDAbpSHD8eoNqdbgnq9VllSrFilrmH8m/A1A7gSdBpcVPv7
JRcqaJj6aSErDz1J7QY3rwndMXtdwzNnmMN9tk458MryOCWU/2CffOHyG/lG1lLN
DQqzcPCtPWypbG5Qg6tiskP1SdPrRQm1cBkFXMnuNxnjJohWL/R6Wff/siuaw7JX
w4dbzuzmV/gu09d6qbPXj0jaevz9JJFK/XqsiucdkTC6SBqOD/dTgoLm3+Hun3gO
T/nng3bz2bFM62wq3/ZvXlb6EjXlQPXpW6QojnyzO0Xq54H+Y5hA5zSg3xuJoNfa
ou61iloOr9XSyA5mtDT1tB2Kw7sFPogAAfog5EaRxpj3/2QyXODGVD8q2zKckTUq
vgtLs2gzBAThalvwVHL7bb2Ju4mqz6LHsyLYxXitNaPECMX6KViasvgK2DwX6Q1x
6CbVUXICR5+KrmNi1j1cQSo61DpKP+gP4+UXzkme1b09owOktIDaBykc89YUuzE0
OSsakjbtvyIlR0vBzmf4xRWIi8ONdIfwTJTW/teOqTTVVaiMPKuccVuhe10QcBfV
4t2csPzAptNe6FGX7mzwYn9iTpw9WGV0a++KSyqb1+xtj9NnYaYXXrtXGWNGTnXl
ELYkahGAWfHGihjjrxh5lfttGbApffSuvW1vrl0hO/B9m+QKt7Ko83xr3ureTrbM
PczKUEsCEFWi+dfwcmkdAL3NxFT3hDpTcleCxVcDumG+a9GxF/Qj2n89o1CfUdTT
rewAjXUtyinBUFD/tmZ6M6NQbGcdR6NvWjwdqS2rva/2W0eET1uglNMCw3Sthixx
dCt1YVHwBJ+tyql51y65FOGrm6o2WSwpveZmmxGLCL8vMAxMyAbMKqDwqFXWAV79
V4xkKJyC/AmhYQnPxlnRpLJMdT2ZslENpJOgGKgS7kFYXLqlYFP760qUhUS+TMnX
15H5CRkZUGAq+Gth6llk+mwXE0Cdh8gbPL9QKoR5qdfUQB7uPg+bUHcgzX9iX5B1
T1DrCHUfc1zuKITA0TR4zJFuJQx6PN0/DX29aAuuNUC4lro2HL50IgJ3+8S4s9Mq
d6zSryd687rE/moxuNMe9DDFhP2q9fWkjCZOCqjS2bV7y4UuXYPEFLIi1gVPDK5t
IMuPN215KFn3e8LTZyA4JD51q4lIqhEcbjcZpRKKqElGYkpU3rO1dZhn6mh30Pkh
zz1Oq3DkAALdnts3BiuX2FvjHyLmVnvG5/k5Et/M+w63eF5ici8dKUbtb918Rgwc
Z/Q0bqH5jpqbxB+AEMRJNa9JgBOl6MOcAmAyuXMliaE5zdFZFOVuxOpQelyud0jR
yw/CaLu7oJURu+1aj29TxcTmnITzJe540qj3chJmzK3UKUBcuVu9dYHCAL8LMUAc
h+L4U8FvPgxYQLsVGmgPZw0y+h4pkKZ5R6OM2z3dMgHvJ52kc1NBsgV1p0Rp5QoD
CW17OJ2LJwFqKkXkTLugRMwGvDz6n/3aBloYlioy41VERDq8P5t9RaTIlVseNh3c
l7q1kQSQdfsXmpwZnnljSz3cUCB2l9PI0nln3y5ArNCJnS7AKFKP3cXGl8/sJDEZ
GCmp7/s+sTr7gLrVPLiV7sdJwAQfbzxYzplx8kOOKWAwWOlwFfgAaKCspLe7yQ70
QIgeym1larW0Jmd13mMCqqdgayMbMofy6fF459UP9Of1fqCDYsrn3b6CvabVyyyp
2ZS6EDLbsZV3e5uUTtq7+qv1FmySRLwQ6CSKcOMGXnELQJvEAP3lbOQrQLeZoYoh
cGLVzI+d+go5zZvNSBCesEJgzn7THTUzS32U4icDdNhXqOWlCwem2G9fuNJ8mgF0
+r3djkx2qb7zS/ZPriasq1bhh/uwcEMzqkddOJSi07xPgtAtWgAdH1CaYAPx+17l
0Asn23aSGwxbFunYLQ+lUMzqGbFO5cLYrKeXdQF52+kTKHzaOhPyid+zqnpdz2RH
ey7SChry9wphThrAnLiYwlupSkuLeIr9MjZOhI6p58JS4aGtGnUIcr0yO2WakKD7
LhY7EALGr3pLH6tf4o3RCFDDH1WX3ItO6Omg1h9582pCJpgv2hviIbU8dRcRzv9A
p6QXPyQA6rN8WFCa9KkUmO6hNuCCdYgR1BU08b8RPoRKpeORe+9mosi8G/pn9nu4
hSsR+jatcI3biRq1SqeZip1vZBFb1qUoSxNURy1bWJhuS/jw16Ej7Voczgyv0JGe
F5enfb65QCv6369x2FgTGdqqWgSyaVHTsFd1jrrfx5NywDTP0lP8mHWXVY2bjaX4
CahmJF0TgKy7Luoi1pceWX4Nork1HWkUELs3Up2rSM4Toi3ND/k6hfBJoz7ah9+J
ud4zqwa0jtOyPrd0KKu03sa/jG/ya6CetbO78lpY1N7VI9Gn44VYf7GQEh9Yhx8z
v+VT3+o1ShKFd1JwTPi9Plm9V2dgx/hDIo4yezXrWeGMIplX6PUOunWkWFBllxWN
+J2SHg2szehAZtU6qGA2ZSsvVKqKy6p0QRMtWGw8BCEKBm0MtBqSZ1DnSmKj1jjD
zAXnDfm2DCrYzyyKA0KbphylPcsYBHsvmnDSXy0lRfS4CJ/gFwSlsQ4gHB5auLhH
TZTOg3zXngsO/leUTlF+X8K3M3TC1LhoqnV+qEyuxGLgKBX+rgvv8QiQhNzporK+
L1/WUjJKUFZ/XZw4wfREBzf0q/e3qtmlfeZqR+SiOQIBqxOtM9XMRMe9Bf6pjji3
POTfV7MAJ45N9vuoj7iXCOv9PNnnCzRJ/1omiOYnYehzN2yylWhi7UQBs6b7AOo9
ZyQFSdIwKja0RxL/Yjw9y7Lh5aznYSS7KzMKuKF/3nVEwAujB2iNu1ITYbTNinzA
b7NfeUvkH4BKYTFX7ls9OfvLkB1dd/NT/a5/BxFt2G/6iCpVX0l1CrwN/OUz/hUw
00qzQbcTzfJ8YkDZEu4S6PboUmE5Ylrm919byRbUkwvS4rkVTsZpiy/dVC+i5MYp
z7TtrsIetdj19SzIXt+rkZW4PS/VTkA9tQGXNd9HMkv90PQwVL9su6HuTXIVyblf
73Q6ITf/thkoNn6FUUchlhXIcGGF6LN+tIm7BZIhYseLfz+gMZHW/brAiqxDRbPr
sdF+dxZ65VbFUhbMOXzILzRRJJH1P6GwseWQTzrzmQB5CdnzXeF39NNss+U7ID0G
qG06mOOxUqlTHpFNslofdmDfpAxzaZeY42mPGTXXCB9O7oF1Ufjpjwy+f4Mkj12G
U//29B+UsQyq6XNM56QYxyUwVk/zRNc8wMk8wbZxZdZbOa5+bDertlbZoDVBzD3F
ZNUrVcXGqQxacMHDDZpchXBbNvB6u5zjrm1Ztw0X9g61FpkorVl8IScTa3tUT9LU
kpUC3hAQHnU6p5q7+NXNMj6xlXx4woDEBxMGesMHMIf/VpSkY9HIAYEgC5lrW90H
FBU/GSHPIvunQFrzt+ddfaJMe73mnsjTGErYEphrPo+7bVzc6oTFftU6ppIClQLE
bg3a/rxcXq6/hoC0Yw6XyaPBc8RMZajPhHNEm7eam8lPDiolezYAlehDw8jcEcuB
inhH1abWuCXPSdY/wHz9c4UhtpRz1v2cZnfJravfz1pr/vovRYLimdH7TxcT+QVd
cssK+r1646mcJxdA+UPwjiL+mOoV/pxnIbu9NIrDcIZY1424ypa7/K65I05n/aWU
nZB0Y+6ctzb6DefcpFGxqxfN5SjA5uVxgeJvMetZfi+eSUllXTWNCOhMxghYJphP
MP/odZlzIyK9vMCUcC+Xwwnl5FCLcH5/I8B6OyqggWEZYRL9cdOraQs/0MLU59E/
b1yZ0QYFwnnEQN1v6qyXxYxx9s13hv784cMpmxQNyHozxi3X6blO6OFKTNrLvqSL
2wuo5Uk97ctOJaHU74YPXwPJLZJOX8axwumoiWeLaFZhmZYHia2Nyc8DSOlZUz7n
lLnS/l5y2HBNx91tVoHiP9FunrRnKBkrV5/s/tcnbNjH/UcTDR6Aco50OOMeRB+t
OeWVecBrS9y+pklS943sJXPCBndUV9409I20xYd9Jje+2DpsH/YcMaqBt/8McHS4
r0C28wBtqz0Mjph68U1832PzJL3be9w8AttKkgdZpjO+i8PdDGJFxSc5iASvWug5
ZS45Zjj7dClrfLOAJ0xsOuJEY8SUWsu0UOHHTBJiWhlMyC7raRrtv3bbIHt7mldN
kDzhDegF1MiUQjukxndu0Ztle702JcE2Xe99qeOrqcMLRVZXQj2HeAE9KeJ07PZy
PbtJRuZYUvJ7ImfOy5yWWh3rSv16i4r7/9vMqDvh9LdyKpfOvdGavLMR2r3KR0n2
Xu/zSK/wF7xN+jBfwKQgfaQeZmxSUmM2FB7t3B6RAxOzjMSYJ9zbj1RWuyikJnaB
2zDWW/uYst0T0rP13/y7Dx6M3mKOjubN3ZscbXW8QCBHEPaV3wzPBZX1qqfxcVwy
wbJ0q2tbcgpAWnxFNG82Jp9jgaOiqQnm/RKIK9+tU8TKGW/Ic9ozUzTTpPGE0grQ
+Lvk5KMmp4Bi+lq3N+fMYcKzrHMo6ZhKz90obv7N7xI6AXpJrhdPfFy2FT0Ut1qd
QxdCBtxH67YaxEHWikBCkSxv6H+VSQbSdzugM+pN7zP60tmELy51tn7cE9JqIw96
W+zG0x1i1/xmgvMdV16EdI28dr3fqaLfeIFDSf2lkRSJsRspuQpfEXCEYIfhES63
qyoFL0C10fgrc5ZXPCr4vrsdvO4IEVuBVSFhaq+y8PjiOIqz5X4fFKeJeXL1/FDR
oXKCU6AWtqloMRTzUM7SYL9UGqBT4rDfeCWQFzQ2zILazsRktBjpc/vnT4awI0Kc
Ouu/OxZlPbfexR7cF6OLSOqC58ASSEG1FvssjXArnJ4kkCarFu93MqIf5fycERP0
E+q2iqRDaLIoKtm8Chksa06Mx+2q73mtPYUDreinpRj5m758Q7pz1L4oPNgEspyH
S4iI/KF7Z1ZhYGlEc/2UWAOc6jZMdhqFubsywIAwAQiZw80jaKfqD+D/fFAGqmu1
fVyQkQg1Lsx4a67XI/sdtue1ri208QN40XpFNYvVlJUedhKVgMV0Q2oRV3xGRbQ+
+1FnsDyke9/wNZQ9SLBnc8g43Gb03JZCdoya7+xX4mQwK2N29CpLBV7u7IzveKhN
crgz7kZwVMZaUsIk5bVCmgmAUtwaoKPtgY92WYPHV7MMNsQYiZ6LLy9GCjBgfx2E
gfzbObzmk4f9PFrsH9rjiw4qLIxTJWzV7F/QNU79qyCXHgNoPvdD2NNZRoE5aNSM
8N1GW+kpySUHQ6hm6mzEoKI807VBKNNBob2Nzldy6Np/XiCuYZaA9fHn/gdL8bJ2
sGGZ777qLXrps3PFWaIuU6scLrzyFDjSJjH+1Xr4EPC2GXDH4PL8M2quy4Ahcl8j
OIHFlT7SixhEmTiI040iQYE3YlwRBeTmK8Xl9GBmbeIHz09ENgaoVD/af7jDoI/5
v/HOndGw1/dUOrYwLlPsDX83HrLebFSZXdVhqEn+M0P40TJAkI6zuhDE6rDjV7/k
yeRlX6AXn2h60Tuh41rhjtEa4JjaFmUX58yHSn81xojpkDPW70Q2pS/yu4wZpADi
a0l9AQLmmR86rojSJj4BjRkoPH+KbWzCA39X6sRtBm2DS87Y7WZ+tM4jEZG2UWJR
KCRiov5S4i+ZViY4VsofweHsvzuR/vFUGn9MihpjWt5++uHemlc4OyiHqvoyLev3
Shuxv/wp8YobskDcSLAgzJhBJJHHUxcUagLrxrqGK0J1WIIf2Q7ij3xuIhHLIYc8
UdHdoG5y3WLZhwEIpwhvCndRDfCYpXdnohE2euR22SwMBWVYxLQQ5rMXh/LFCP8z
4jEHA+EFNf7/aJyt+AbScaNlR8fPXys9Fxkqy66n8tFnkVGmqbdDjccI30f0QhnS
ApsYTXaDdkJZ7L2D8kEnFWSCnf7f0vj6WcbrGQpYntceCFhjJgh+Gi3YafyQuLP5
B5Fk+h2cx8h+FrKaEq0W1Aog9yry0J+Z/gIu1QgMU0yzcXjE+lHb1LsyKWcJsR97
L+eJpxTTlojTSn0PiFyhWpzLHJN9QUZPeQRhC2cDnMU8aT2nwTuUdGL4EFFWRRKB
VKI6DsM6l58sf0PNBta19+CCaCRJrX1gwPzx4rxNY2n36TXRSk9AUJ3VodhoysCl
b6zFLBvqbj8D7gIiMp53nHbUHhT8aRqcDIQcdbkfRos7GCp64akhDXkoKmPkH33Q
7LXqYoh5EFT5jUK+eN1xEf4sIAD0JIL5Janzjo37DEw/vmfHCpieX5B0/JOE9b0A
SwCvsZTCrMkCU/A9dldYCpsIP3BoSEuSsICRRnj/CCu3gdT/OEkBQ9e+lo6hGD9x
ZgkYfzV7OEnYK0FRIJT30GJ+F55fYUuYC2wRCFBw3S9g5w4396cUXm0X0CfldjLR
keJoKEGj+oC6co7IMr6pa3ZX9NkHzqYzEhCRE183bV0h0DJR3n0A/xcJmC1j7F8n
DI3tFGL9L4A66NxZ4zfrmbVbuCLAUDjhG4AK1PR0QfouQlQiicqiWoHpEu5JXu5u
yTPm0sInh2/zoU/joyJKZYiEff1Wf9Wly/TvaRxN6RvEkaMa+80Lvvouk6emDHru
9m+YgBswdTooHQZpEt0+nxwalU9ONRGYPxId36UsCcdOhfLm+SLiO9VluwmBzRrv
IoP3sGSDaf07IE/jPb0N/Ap2EuYK8UTWOEQBaaWhpK8pcr2cfQq1DN6NYvqQNVHW
rAOCYhaYPgm/MXPur+6IdDi4YzbDKr3DHE/EkU8KOpuOJIMNeTrtf46XIG4tkD87
TRbin43IJi1T3irYrkMm8ATb28uJtoolNSM57yIBO3cspNQbOX6KE/A75gC2JB7d
wAbvj/Cr2latl/jHhiXs6JGl2XYrY1BHXhkhjjfaPMSOYArDzjEL7skfDg/x2dmF
gP6XUOut9UF+s+emS0KoJ8CIUUko63GH1tXhGsCaX8M5teqD3rCTJr4fAKfX1Jqc
bgAg77b6B9cchWdz/Oxpa9nJz+XQa4DVPfqs+OYmnlKkp1qAXiZTcYzG+oR35zwN
KP1HamKFpGSORvv8XL1nmBigu/k4XPNRWzu1FPGxOcZNx01MfxlfI2DjvZa0833h
WHQuvesLMjyhBBnVLaHhBFubYIqjUk+MaNg2upijPPs95Yyb7WgksOZtYP4XV6LY
WQDM5MNCs9lJRAXxk/0kMpHwsK4eCiT/pomj5/MRBzzKJB/jF2yPhkJHE6OqeOAK
+RA2AUItkPimqhlbT1ccnmYwapN/Em7riuysoRT2M0Mke6YqCATIFb0eQREHs2S0
lTgC75CsUzXdQCnMhXdBUSPefrjNsMhXpLKlf5mPsbwnTI3Ee65EbGwKTwx89rYQ
4+Z56bz9Y9+14IfSPnFdIhhqGCJZFjsS1iZJhsCYzCfWq1reTaRqHvf/hPBpBIb7
0yQ6NTKUbj0q63HIIrU7gVayU7MEwI+gP23VgNQnmQKGCQdTco3KBIyDp7ykil4z
8Snnk0u9WEP/8V3qQtEM96TccuLMaemek6OcKJrQYS+SqKjhSKq6ulo0G4IXdWU9
ydfDowhEYptF2B6zxuiHmUdcaY8yzmsuNbM9Hgh7w5rT9bNysGLQPZdlvi/nTQj4
rrW+bBnhjj6C9fLPz1vfybTt+4VcncuDTnVsHHwSYWKt0fiXyXpCJ8t07+F9gH9E
n9d+np7SHrOWpcrCdvF2zKp3gsZS5a3/fIPwd+1MGVEK5ZwJgVbLy5UDnHF5aui9
hwAebaLY1prmXYFD9Zi4E6VAog7AXGdtqcs5VkIoihwLU6IAATceUJM738V73zzf
6s4i40XB7O043WO+AYeryzQb5sSWLo5m1hLSl5qOht2dsVOH2lVX4bm6N5C6/zjl
7JR4cG/r3z+N/Gi3s0q23on2JFTDaiftmMqkXRASLJqqrcnUrI+fgl60YsKlNcK7
SkdqBkvo7fcGoIKVz9HJNXrnB9HpJvFzSIJq5myhhy+OcZ+tke+LhlodkdV3GYbV
sOIxo0JLNwu4zc5VgocV7mus3DjlUbLhWFfT0AO7/BxHprVquMlNRoDBZOHZX09v
/y29YsZNoTZb2vsWOVFea8alcvctylrO4O0O0O+WGdKCzF4RpSJRa7d2T5ttTzM7
k0vWbpwHIRICy2w3kB6+X8n8LqnfL+HfbOdXXnluYhUSJKOewdE3hIkNobvXQ190
Vt+DnnW5A+unUT3aGc6Pts4KMKmXueOwZESjoGI+6ogCEn4gXkT6uyH+vyNbvyrY
ty4jBPSEg5CuNDb4IzcZLNEn1WbT4lj3NweouSNloEEI1OAArQQRnXkRqfilHlLq
yfXUgzdRY5NCucqaL9VZq1VjKLCO1bjUUXGvlaQFpSo6Cg2O+mdlY0I+iRGa6OLC
vY3ZR1eL5xkpWDu9mE2RZ1qoL4m1Ib4ZzCWyMzXec8h6xe5SiHVrL3Ibv2h0eFGO
tOJDF4cSWDVloiu4GxBLZ/gHgBw9Cs6GDfTIMoHD5U+WyWI0kP9WNIVdvaTlPogz
L8rWSHFcvoHpGsH+9ODc57Cx2HrjV9HBjJytQPbvx9vEGbhumDgB/Z7iVtmo9f6B
/ewBhgDb2D8kOO7GMqC3IA/pWha+hmQUYbJALNJpyzAGXnKCfdKmm9VEnZ2G4v1q
Q5tvJYGj1yqoVnuZhrWC4Tlb/fjJf/WPvyQPlVhAJ9nerpZRX4J7c97D1deHWnAI
/aiICMAZJTI8nLJUC2bdSBw7DPiOajCZkrTtqoM/TtTG74kwbgBvHKgOL1G9t50n
0mjjjAKRjW/6rRZDxGv0/UtikJx11iWRgal3Xi4MRe+Mhmw4q3NnKw2e2TLJgK/v
I/HXVImnYZTPkCHeGgEOEtlRgWb8kYm16ABKct0T7yqG9F3gRDR8PWK9V/PhaC/G
ZmCo+tmJ22xlWrcPmfmRaSLWRJMk5jeFha1r+BlYfMSm62KNxocj+cMfhQyC/4ao
NFAHF54gZiCD3khB71oAIpN8u/gmuAZoM9VqTQbuOLuOL8j+BFbyizWpvuqRa2vh
bvzGwe1biw9HsBV5NTFNJ3r8U1DGv9s1Y8yGOnl5HPZB8913mJdG2PZbt5Zs22Qe
XkeGutOrwi4IP4c+MkvphKL5mHnNpl8ficRA/rlVhnD6/VtkXK5Dnl5xanex5CWw
5GhwKfFrSNTL/Mzn/seOppyX8AhkOYBd2C34PF8ahQ8AoutgSaMKuBfu6UbrUmhU
R6LHBSExEqpI3LfTYLUTVHwMKgENJVXQbCNCRfezTZomOQ6/4yGvRJb31yS4qbuc
GIrhPuV0li9MM6/NtOrolzWSPIFW22VHszZyJZt12KD3qZcf/0PNj+bJy0EQ7rbT
oWZazeCEM4gf8oNTGQBdHyBORmyRAuE6MFGr+lB9lmi5hj23OJ5IW7B0y6RRMKcf
iLH26y1J2WWOqOZ07Oc5rd2JqOyXY9OPzXNGICfcOHtwHNm96N+GxlHy9VQYmC2p
BreQXmAIkjYfV8pKTUjKSc1phdTHDmrlZD4haXwVg5W+yOAdLEnlgBuvfTo+Zn3b
DiRRDAoOh+2JjQoLZUWG1Q0+kdT7Ly+u1EcgWVJz7j/Q0xyRfhPixwr7qDiKf34C
I4qoIf5tuE9tonxHJ/xiOLwgUo1XbnfpL4nJzroF5IVJBOYMpS8o72Taz2y8q5De
BKEvO6OssWP1lFZdHL2w/GOF60GfgFsOSam/pX+j8yxVXXArpXqhb4NLu5aoKVA2
Ozz1jG6MM0+bHNUen5AGm0oM9aHYo+edeUSxXO0GWGR/8Rj8TYyk7PXVa7xbUhfr
qPFluzXZU/dSVmH+3AXfk6zrfHwYNJCJ6eU364blTWfCrFHy7HAFL4GXtuf8d67a
iTMsW6NSpgxpmx2Sqp1tq9Ne2nLzbVSZOON+vI2G8W+g5Yb6YllfVYU7iOOazlV1
JsaBlog01qyUgNm0wShHCQx4tMAx6fA9tjc5oku6a/SSM27OIfwOkD3s4fRMSx2X
ROHjnzPCdw91OfyCHFQ+ly4WSsW4Ou4WgumOKjX+HIqH+MVPq6AnH9fYOtwNJH6T
gLZ302NnzjdquKoy5pUiO+5ki89IdPtFlFoNsTM9YbvW2gafkT/AE+ist4yoSO4y
l1qJSxfTXuMPh8df2cuZC/Gt2AO/859/OeSSAvpKUFMPK0NTAAeedYt0BFka0mch
ctcV/KhZFVUo90Iv1490DOCa5NGOhMr0XTnJ4P4HLjBxaImXvXKN6UKv2rcxjzhJ
1x0zRjwad08k5UeC+qpF1FIZ+uSgWdrRBSENxJLhVwZ8An1JEBtXms9hQuGFK9V/
9qS1kUwFpO2U2tf3hesV6frRPaCToB64k/p9L5g8TDjiS1QNAgawRSxD24NaQLsS
w1hkqY9fbb1m+0b0860F890U3qdEf4rkXDzw9BbxuZMJoju6fIkY3unHDCPPLBDk
7UWKmMLpoNMtVZYZdfUgjlQH1+s8Y/VJBgOzNrdn03mzjAOz/yR0BN6QFNHQCvQi
0OhxP89fIbZi8yELwiWooP3S+mbK83nNfq7eKhOkp2s/7I5W7fROGBHf9RR274Jy
WZQJoPB6IAjW52cJiBxSl3o1G6dKKdVdvmElVdfuaBKjENEtgWy7D1Ewcl9/FAgW
8a54x0mMQ6fTPNkA2fJVMmvTIY92kXl25Id3Vfl25i19f+TfL/VSUfgRfsTVSWL2
3RhyO2M7tq+HeeteEjYDBaw1lpchPurKFTqKeAOtM0FE7hVWzCF4UR+TN7D+WxVt
e7dJVxq02za1TrP/mbpBSfg3KUMjeb22/Zseoo1D5Gyn8a6aB1cQoejip9WxMWHv
k3HglsjUjQN6Qqo+6oQ8gUB6ASrAKllnRu8r6OPc5+edbcp78SDidw8LkCTIvqSI
2+n3DzWsHPTMakw5Cdw4GUYBQ4OC4mEx8U3VT8Y9xTDW3TPHTEZ7GvfEFBxrQQYO
YjATr3vXOCPinCSKZb3TbGVTl7EW+EQ31wo9KJGm5NV9hRprsT7OfAcimxU2Lc9j
dQ95+QB16ETWfTsuFLKVeYSsw3BGylQEGvpybadWvjNpqE4MGr47iaSHFwOniSt7
11t1MwaUOuMxvTIX3zQH2DDBYQgZqoqLMSe8xyIl1DqAcITSFmmkr3Rb+kBt9EbQ
Z0tAmAqouIe/n/ZBBmYP0tuC4xy30LDiFWMbE5+CQmCgzC9alWutFPf06T6co3nW
JnUiumniim3ZV9piy6ovdWHk/HxCKP2OiulCz/geeuT0iWnpc+mBRBk+OoVm51hz
/37MBQv7+OwHq8Algn+880gsCkPMiMaRrnbw/tyvPGq6CCNogc4ge/nt2G9x3oVU
Oi5qEHUyY2gEAzHW+LFdGOjBIb+EcKfVWqvx1avfEyRJicE4DHaOsNhnIVlsuIxz
nYKWHKD/2vcr5ghzZypzE6a9YOd79lFsgtSYA+rtM7EKrM1DPUnlQrlHWCSvcAv0
YpOzX7JOP+RZKoKLdyoJwo39PTDbVkzneif4X+k0OTezzq/WXciUCT861xDcZvNZ
MBFuhXmcFLHrrHS5Uw/ec2LxpCGhZYUHIN3v5JR5AiQm9B6UNVfpglKIegaUHzJn
W9I5cXZpkwd2Un4WMCjoWzq+1CkXTPRZjowLAoohdVP7zm6H8MXlVCQBkjdupdsZ
zr4IetqOnvHJU6YJJ3zOGmQfM/efyWUkw7yvKpdZcm5qgLXhzCUSKYeVxRZ3NnnU
kMXasZXdfTJV5Na7fQXEi0mchSdIIaTtMaGBuycIXB5YKbPZkWhAJDI12CTPsO5y
pnS7aRI4ASXWS573jtPDN/1C6Ob4dNl9RgcP/QHr0NU1Ye5M0AHsg/Ok98QEIvqw
0cIwS+cKHmpwtWyaOu7YdBK1k5FEwIU2eLttE3WNpmQQVBMHiq/mk9D9lmtR8IiF
EbS98DjvlCludYKql6OR3GjuTZyzC1SvEsh7eDJ+3dwoxxDHGLwWTQsec1V5Pm/g
irbsHzaykzjKqXPHqyMGORoXaFgRhChCpIe12xwvLxTvX7wpLDgg3bsravsHyKPc
TpfyIo9N1mCShhy8yWJ5cbPsgOC/xkLEeBOlkY2QZbTHwK900abKdDC3bcC1z5+W
TcanaS81oBjwKkpLNE9bTa/TyuHyL3I0d5jGrKz2Iuj3KClrnvPEUfa6ndMqg/X6
08gre/846VAYXfabilqb+NKm3WLUNPBAh8VOAfsG3ckyGaeuijGwcqaBaNGqFFhU
xm3FaMYO6gs4U5n6m2YJP/htUBhwO+RT9kN1VR33z9alXCPNN4FGHUCH7GvnIwzK
2x5qTNx0jpPvZjc4bjRFCynhOyn+2noqD+9j61W6D/Q=
`pragma protect end_protected
