// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jUFYgMw1dYnl5Ai3Tz0fyKDBdFwJeg9H3kWvRpraIVejBnLlifHkv5HQjVSQc/s1
tgiKjYWrrHftFu9HIWF7BBlGbE2F8iPdGzsnWkqjIUBZODTjucAUGHipxJEDNx7Y
XH/wv/2xaIwBL3W1k9c7uYZTtY/7pyGW8Tjwh2+6KpY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9200)
Y2G4mDpA9yl+jrB2qz2dGtei9xGVk+TnE50mwJY9EYTLmRlD8P0dSjKG6jO8PVm8
ZXD/3SHhneAy1WjPLaHCoa1jUb8KgAmtMvF/HqqOGNYG6YzkPFuY/Ug/GXLGMnZo
hRg7rr+URN5xXXw1Lu5+aUbyR/umJaDTV/g+9Zlz8AOPrzWwexHdDW2jboM/YlXx
1g95CDpBTQrLyt04KuZgdH85Jkpbt+3tPV41Rstu/mfc2aJpfjbjvd16lemrVECe
8i8SpcOFI73ZZFQuF4dSpm0WycCDe8+/d7lUSipVImRDT7DP8dAmMR6eUJHpCtGu
wccGaLHEHsyDCClQiuB6pb8CgVpyhq4e5npj5IhzBqjEdwdLhQOBkh4mPI1HL1YT
I/jUjUKf+h8RhIAdE7exvkRNCyDR0go3r7B3Ax7+pewv1NQ1PoTuHGFgUWgTo+Fo
N0Bv1PzzhwpsgLS/kVtERC4oX2MqiTT3jlq5dET6kVdo9rCkJWmkUeT+8bRpN6zF
P5GXrYwJlEsylvwz7vX554C9QbxjCBZqmRJLA/frMtpEHsDjXi4lFvJw7vpD6sfm
tf+6Y29tEjsm2CgfSD9iQQjlR/qKYGuf6yat1buOjIjbNLRWeVeqFiHMndTCo5Rm
t/XFZEjmgHbMYoOBF+9resRiiiGXSIy3ABv85cQOblD5TdRMYb/45ifQCEVsu7YA
2BREL5FdOMeUi/2HzOQGEh2lAks5F2piQUqeEyGWBeFuBR4EKv1xOkq9ffjBH7Tn
3esY4cnGp+vchrkcoU74F2uLnodtPRW46nkY8RlkWY7/js4tb/DGBBnEpUlYg/2C
mNJnnrOR1Uy5D6Hm4YbFsgorICfsnTZTOpRfaBdIHINWWvTHzJ+beDPtKDcxlvLs
c2UjvEMnBgGn9aw2Ai7YLgxvTfSTRI9iLExrtl+dkWxUWeed+jDf6dMx7OkT14SJ
AjjvSTdvTGn1aBiO4BBBGC4N/JF+ki+XewdgfhRAwfWOWsp/zfuxlXSxTmC3wJ3T
AdzqKgRy+h9VQaRI+mCihgpCVq6fAnCZdDg9dx8THTi7HO+NrdBIe0NmIzL+AA8o
wmU2FS8hlq5KWtQLRYBNVYREkmCf7Sg1abDzsyQCeMxfJMexpINw25KpfS5c7/23
EoOkUugVpGuKnPQZO+C6cE26Nqg6A8HvpPE/by91DPdYQNc/u3TPLCnRRecvVHDZ
+t9c/tCRvCszwfp9CxkEsj5r43CQ62gY/IgzLEqd3wDhGH+Hlc4Hyewy4UWCm8Jo
tdVoHsHgoI1Naq7+XeOOxophy+cI7QZYhOrN7aFrlMmjszsJwZ2QlpXB6SSOlQrx
UwmomCNwnIQV5J3TnpbsUP1TBCCEjyN4T77qGHt3hTGlAUibyD77OWkRzN6wRkUS
yFc0zrVLGYXNWJEvdYYu+ZmKILOX6nv5FZrTWv/iQhCKzoGEQf+w+Y3SEnyz7rj6
1OVZY2qB7g3Wki0nxzDyRwforZhm/TxTv6E4K+5Znc4wYeZBwUnW+Q6joJdmjte9
2R4Jn76kSC5kgUUKpBojbCQkN85ZcYmvzmcT5K3Sp1eeO4kL36gvBu3V7JZ9Kw2K
Q5GUC/y18DevoMRiWqhfHFtSIk3BrKNwo8mfbzUUqYOPw2HAo6Ngy6PklOPLhA5g
yNwTsDTf2WSAJBYiQgHgdwVmeL7XcicdcOiazFvGFfHpZTRpZOsHTQMHBlp42bev
Qb4mO2D5LX93BT9a3KwJZI8ubmCCJDLmG6GWsHtR+oyBcyCneMIH4u02P6Pwi1du
be1FChEGeyrvSTqp0+Ncm64ULoGADGqwsp870oDQV/Nmpa/Affq0tvck2YA520v3
45bweYVkaKI0ugLHNTAhqnt/VShNwyrCr6J9ocVKBtd1Fqbwj0QMny1Z1CCYI7w+
R7QK8YM20eDjaELsOjzfmNV7DNd3g9sAegMSXic9lMkmxC423naBp5vqmn29ig1F
xM6OGdWR740/FJGk/PNRbuHC667lbNRwQKfirh3Sg+P2+xPRtr/rc1CBqC490RC3
le0YwupphDFwfYcSxLWqnTqFGt5vnoiDCPwSxVs+rne02S0HhjIYF6MosOIUs650
jYnMqFM6NzMhyAdGp2x5WgquQ1DN1CsPLIejzhpdKZOp3ANeytnaC6/mqg9pHqdK
yapoXN8qoHCz3w2kMkVSt7/py/KR1pMXXRuPUBpqGFW+kRmXGQlIf8ZnN2y6nMEn
MJU+a6Uk1jS+hlNPywBL1cdJK/rJnRR2vmIBrvd4egHTjmERj3YijOtBpuF+ILXV
d8TpYdg5xVXelEKkj0aTOyehADizVm21AvCPACyeMYWNjaKysY1lcQ5Q2e3tU/C4
dv2ttGzHur33bdjCwVaIYki+jHJVpZPkfBQ6MMSh7hf9dKmnRQglCKd/7U/VcIUq
JQqjU++BnukPB/tEAlsLdXjxLRCXLZA82HIBZezA6meME/N3Qyvfj/cTJGPNCXX3
J03Q6ien+vqnQFvu3HEvN+Y1Gtf3UGtwPZp4UhgPHPf0nA9Kz8tfcoeYnkNGcdg3
ZNuuBC/81u1zrB+W83heHePGlYJjIwwjjSU7C/ZilLOAzDWy38y0zuUfNej8G7Kn
EfcO4nRTkB2EAAkCzZu1KESBkjLtkHY/1dUQsUWB/W/N4uyeahTkRXnIVd7X0tyZ
ESGcevP98FlnUYh++1YH9zBi2f/EvNS19YsuWWKocWkc9xhGv9bF9jB//FsH1CYZ
tv2MFWDDnMWXGblEIFaBHFIHbMVFVUlqkQlxlKj141NHf9WlgS5R/uCXQeXaTls6
j2r2CFeavTR+HF1iPxXAjMxHatNkR5JGVcZp5CbBpuRQDl43Kzf+zCfbE3EzxmgH
oJaR7d25ncB/+1LuF5JnMr/t0l6MXy5n2WregBho6p4E8CkBdWoh57XZ9p3jW16B
E8ndcmkz0du5XiTrEV4G8yA38CaVTwXBAsgCQzkPRdly76olIfJnDxsyDE6oAQSk
BE7fdI3Ms91/txGDERnRXMwfF7nLofMzQmXC4hPFlQ5PJntrMazUA4Shch9N/YNL
cGSkencw9bPllVm/Ev2avDSiXnbiaiahKvIhMIiDdBPxEcla7fpwAKxuhg/wpcI8
8QK3fZ/eb+KGxA8M67MXM/tNHrc2SJLP3vKO2BzifbwL/IcnagNfRqdFsBFksW3o
KXLD/NTexV54xeivn7YrQDvBD8tYAZgQnrxqvilX2jrKZR6HNgFiL2ht4z4L+DK3
ZcAC/E9G6K9Az7sMsewWpRFx6eDELOm7xQGHfTiAPnxIcJ0wkk2ozB031OrmdhY/
IGIY5gsAk67Ty1zt8o3i8Z4e0bkQ1xwOxxmqUKaXuC6AmnUv1aKmKvWBdWwCYgF9
EyQtfb5L76Tu7lFMsNjhYsuLrJ3CTRfs2MiQbZN990zjGVbrsmh8rryH10+xDFsp
k8XbAoFgDOBrs/vPKGz3+oxsXczbh+k6Bzpfhiha+8gSw2sJNRoQzUiDrvLCYjlM
A3oXB5oF3/LEVlNeN5K4fTyG5Ho6P35dXBC2S/Q2vXvmPHKFAMtSsTYKyJW/Jqyg
/M20t2jB7pCQRKfAss/e7brTku6nmBU1wMlo6Ipvux3wmTk0Eq44ophc5Xub08B2
0cKpHs3q9cX2g8m6fi9wz/vUO1slwaDLsRZZN2t2bH2vDvJY0SRrAflb+Ep8xAvo
nn/3ppP5q09f+cvV86GPVQPm75CiIC0IMMCUuZcm062hiAe0zsAWEmGno7wgt0HJ
bhGOH+0Zt30GlPTybUo5/odX3BwFbW0kuo3ESzn4Bu8hN8fM8eIdSFfkUQHbA4hQ
0hWXr0bxwVDHfFdhllvFtdP/WEWguYB7k836UkX5Dovbm4P/rtaDQRXlayQoXWPJ
ah6XS7S4DlfHE7sOJxra0Ybka8kEsORXIPNRDlN29veENV7i/LCq9xvkZsWBLLtt
ktSLmMGWrOWzOPG3Gw/RO1/DyC+BfX1acNV1SkJ+Xs6unb7sJpFfuhc2FszgYk+z
fP3LuIRWXSk7L1FMLqUwExqTaD5+5i/EDBWkjGl9pq9c3vZpSg6i4QGO9IAJ7KvB
dw/UD6Nyg9COg1LpXRp7g/uBMcVC4aNzWQmMS6eK1c5aLf9tT0uTEPCBBEBpIQ3p
DuvfkQUQWZT3t8Wlia+I91trlWBzEQCjLk90E34iBLlAk1TJ87ZePkEuCfIuqj2s
62ReFeCzarsygmbTvw2yBZKXxQotHM6LQNKumZsqwjMVqRci5faTxx3J5U3qyzEF
6mySwV3XHuOe5hWoj6K/kv8CrMRxVhh4DmbQYUV0IERXTWS0th5jjhTzbMS7cp77
Usgbd+7i4an01A1K0D5xrfbnL3+cWlx93oH0X3mze1BKIC3WljMukCrKPrslDNm5
EdjJCp39R/Q3m1Fa9DNuwdVNCU9/1S8Sr+OpKCsMYIOFmAawXaqOJvaQ1aJOu2jE
Pmov8JKqPSCFKLIMTTorZMXKhc+NdbVRwknGJGmKIOk+4ZFe+qHK1X5IKV6HY9N5
BVMXqrrUDr+RyOGeTVcyF0yNL3+95RlQEvDkUFzTts+cOPdnjOlh2BDBmrrtW0IF
icy0dL0QH3j9fZCTHVBDT7+/YHGT8ihphfBVV65T9LFEkVQNNWzCUojIl+3pEfDF
trUulVVALc9ilWUnvxAi5oYjGXDkbgxer9670lDX9lqeJWzw+HlQSvnTSRY1/I59
uw4w05t7aXYvcUlR/rwV24DxKX67Pm9XU+jbANrx6leyr6Nq0rQPfVrlnhvCjxTJ
TIx6Ofi76dKZ34NGm/qIDFVRhOXRi/Z9ndAxSVNUx134Na+1U4abTTvebI7KPTlu
zqajNNT185NX8gGQeEcb1xMRejAF7UJiYvN5SOOAB4FfuZDJDyM6CWtPC5Odzkdu
zQwFHw3195+1gSJeauYaqfOoZ59EL2v4XwsSSZRxrBBpte1a9VkVFzD648mWnUh/
Cld9Grul4Snf4jasaIsXv6Co+50O6XXd+Obge9r4fYaIROwNokuRXKkGnZUxuwL7
agsYiDaQTG6zKaSIyEdbR+qidwajW6rlfKFzwa21PJQynJLNrf59t92mWDGmSQt8
R2lMjjIK/Kk1v6VrbRAyhPIPgJ3OwSfOyI7EgCXFYD6I0irXjRB39klYAlXXzVir
noDOifaY2adDiBHuWB8rBkphYts8khGPrHApIwm1EmEoWTtfYDPicN2Vm0LT7pqr
vZ5exPErBm+52LZSpS1JQLeGd3/0awwTspgVhxd9YDnK5J1FUylGAnk397h2KniJ
tymghNsQiczgQRF+xvQarWPVtUikWak1/Ub6g6gu+rBhl1iGcECC6fqceZulpWHf
2Weh+zjK1yWnI2u+lEVTwQ7D5QgKMQQWn+7d2q6qAD6o1RkPG1jH4an7zJmJedSi
flCeNA+3reLdi++OOzvdapNoo+tCCxHt3Wf8/Ez9mKZ/l5hxEL6oMVJVfabiw++X
aovlQBQ5WT76qlpXEZb0I9GN4s4Hv9hyibo8D4dntaDbNs4OlCI5tn1GLJvb4idW
0vHne+k5HAdhx/yGl+rzpXKL1BWoPlQXl3AvJUG3ybn+oEqbxFciWjotSSHzFPtV
kfBvWIIXn/KWEUUD3S8Aj0XADbAs5p4qltBEMneKbdYGqV6JJK9WdGZDkEQX0tgq
Fu9Ie8BSsV+sNFWV6XjkNIMbN5au1PM6d4gOj0JTWZC6pkIHgYu4hXZ48qa99jD+
rkyDvqmTXzGELO+ATkd+kH1t7tca1qQzDY4mjhpPEKVDVwcPP8PZGsNr/0TRjXjV
Q6kQkaBHzIFF9xj97q13jgTWJ9ds8kJ3yB1NLGehxgNZtwL/UJLbuvwKi2mxpP8b
ICML7yjVT434G07+iH+cyiAZSThFBqsJLgo1VVaWganACz2SPwXMBj13aH+kpA+j
a7Kc/dYO7TkT2rxvdoUkJNZVOYTeiZKDSTQLCL35Mj4lqujhJv2u+I3oUaQhIdZi
/F0T3s98FwdVsiU3Paq2REIIy3qWNboiQknlF3zLKfdrFZVBGNGf+jZ2QI4sEtCf
bV7CT8PtQFJ8I+GD2XWT7G6nL3Ry+vg/me9QWdnOThvVR6n8wwlm8vbf+B+w7L/0
WxK96qb5duriGgCYCUOPWwzvZ9o6vyV5yxDqWgPr811rqocQSMnuJFLMpJe8wK0M
L1WWg2PV7lcUgowlM1UAOo1T9B1+vB7dd8Mn2wbLSd3r1mOmHg1wJ76IYErfLghw
sdeFKIg9ynxOWZb90RinRgOm2R64xUbncf/SyMDj3bJrnojR9KMmrd6l9KJ03lX7
qhGClaHpA1Ytp/FU1tJNcS/WGWRmz82idDQKYgD99UvkEHCMB7FmJjh7K4pmFEMj
oZwb3p7u2ZqE0ShBd4SItHWtM7g/YvoZAAvipOjk3Njg2xraEcdcH2028PQWZa3Q
VA/3x6PfJAM3ebRfFpXsZSkW2GtcJuJx/3zR4V/A8XUHPhAmUrsFM6WWfoEasAXt
iEM7kQ4G3zJghIE8jEIJwQbkjMsGU3QILFkx61xMS/hUtXYt103kLraJKMgq5dDS
cOn6fxTqSSr+9SbOLhBh2qLz4xF+xs9CUFMmUd4GZknrthuw6NfAYsuBtrEdtyxX
SL72bQKKS7b5eYt/fBuS3Uv70Vnmhr8cs4bBPkwIGdmhkPCbTnyhUhZR2+/9Si4g
VV4kBMbUdUJEC35R2NMPOhNe/kBXXTBO6O4zOC0j3s7GrguQEW7MR8cWxtbpH6tF
GV6e9bNs+RuNjLi72nUoF2Mg91Bn2q5pQyCU7oLRtAMPrB51WSPycJs8YAW8OJ40
TmoxZ5T2oTHDVJMCKx6QzXIGbV0WLv4BBeBuYqqaK+qZiFYc6Fx5pJj7iSs4IwJF
bXVxxmPmzg5qhAPJXvLsFhgEMLW66Ox2Kf5BMZp6VuRHgt9lMd0y6vVkeKXPQx44
SpE/C2WWy4/MF+DQ74PbZ503Qlq2X4lUz/zsUSZpZH3VKbhzUCdN4KbFTdkJvIRx
DC5UKf9duk9xbrQJdVqwTbOtpb+PZ7vZor3UQPPZLAav+ItHdAvZJLa4EVKzvvBd
fE58j0PRl86PsrT02UxJIkn4+5iI9SKjqgoi/lJmG3gjTW0SidoOhVlWVjlJxL/R
0R+PcnZyGswpO6FjKqbVSZ51r2IzxoKs5laY6XJeL3CX1K4kwuVfUKC7xzz3wV8G
ZplrbkyUWw74FFOp2mNuRBIWKhQKs2I15cGUkcCaYf6hAVoh44OIF4uhpp8/P5FA
0iuV9gXJUDJkS0vGtbHSCNaDe9BofB+sx/jekGc8GWzirM+wrtKwR5VkJBTsxqMf
E/pQz8n6lPvOi1GE1tDJTI5oATf+MjYwCw3Wc4BwhWrqjv85c16lnLgjkkiFzG+r
O0tyvEvVDVldq62CMV/iDScehuEf8k5KKxp7PivwiusJ8sNy74PkgNjUX2UaMFgt
zw+s+BHu+FDJ2+UvirW0aihyyR+ADg+UEImafhJOC0N1r75Ni0BZdbFbGAGTpXwY
A6nfvh8dwdwc6imunUi0LZfq8r0bgS8/KplVjt4spLtwnwwuYkOWbhZ8nbekthji
Kem1xXjwifCXhBTMetgmX9Yi2qe8ZK+8MvV/7mGcjXwtmPXhNP8ZcoY8tyrqKrR8
wLxkKfOtr6IrnYrXx/zxynWwOojILHKZiNP1oX72xSYONljMclBEa/xJjG2WvXpL
2ChR7QNi9IuD3T+dAkPViAy7TjJ58F/hUpeb7eBmIhrzExVCwUdoknk7XK0gv+YS
58KfDm/E4u5R+dCA0NjoMNMmoR1oYDhfJiceIVccIGQQzxv83w6LjaJDry5fVS/W
wWUEOeEvwXxQ6aDjTyLM7b/99+N0s1gOXLV5BHrcEKgjE0xgqkA/iEXaXFHbF6Ry
w6lL7G51AV/seFAmHiZzA91VnTgb1sMi3dL+jGi8Pv1mSvxhN5lPgqxLtJRx/MoI
uCJ4VKn0jvThp0QDVzW5AY6CIzLfbJanECrSTouSGYxm4QBvuRff3a6bnnIJpK6k
7fNKZ3qAHOEZEmf8v/IY70M6hXq0kL1wUHHcNTvbN/4AiQ+F1KKwF1FY7LemQHoP
0Rnl6XGHRvA1vADKq70lB8g1Clgp9m66frTBXL2EmycByOuNnp4HFSk78+L8uBME
b/Cdgyi7G5wZO/tbDlph6RfALOE8LBGedukHa4t5WgXIcYp51TVoye9yjHfzOvQH
0Ciy5P+Ec9cimfYSSiugIZTgAA2+MbpCCJPDw/yBImMMAMisdWTOT0jMXxUFK9qr
s4SRhkrf6xkSQUQyAxE2EjytDJj8XiaTfbFuuzQgt/GSL3bP3iOUJIJ+ETjxkybv
iHWLx9ng3dx9Agq0MuVsMaKKU70rx8xIowdml9Vp7spcSW6P/hObA/GqjKAJYsrd
4v8aXW/NYkHFwKLldm6zPJ4FoilJVAAztKKdJ+oftcr0kEvg9nqeQ0GMdKpZMts+
F4Pm7FhNg6/thnJwg0CNEGDaW3lB7UhN+2+5nzRM6+boGVYFgI2tI8SU9+KZitLe
4LadTff6TyGL8jm//eoTj8olNrHKnfOr2Nlb4O+aX70aDcg4RRFuPFjvxPIbuQfQ
iB1DYJgxy4vKE/fqImWnxVKRXPXoNqqK44dSp5BxndY/pd/Gb/VdMTtU0HpGExRo
9pKAjj112iTv7abvLr0U4lrCW7ptOfecWhsKwJhupHJWMi6sK429bBgagzrlpKfQ
1sHEMtqvIO8U7J+yAa0V2zUbhmqqUeyAEH8gNmY04yCK07QZOewPSQCLXlP7k3aR
Ky9V6TAYxRzSl9d110W+WUW4+YkwOhGZTC05ywnVE4QTCMZJ4kFYVkUZCI13A6Nw
vV06GnCKc+eHTWC1gPLAlxP3zuD5YfsladCm75Tuhw7nu/J5ZHigsLIatMvIh+Q7
E3hiznDV4JO/dxeTsUusKg2DJm9WlvC7ldhS8E3rZ3416alzvP2fKZZZz2FRJUIh
zW84kVtwiyr0/qxDwKkAEA6eHIcZF3OCWzAi70sBI0y3XDrk+FQxi6LHdudR4KlC
cTptz/+LNi6GFkG40yCBIRDFkXygtmAsXq/1r6YQCfjhXSoFb3B3ESG/ydY98T9j
KCD/6ueGaV2vgK2r0aNXamykrit7RaVB2fKtTIRKwzUzmy97uG2DknJpdBgd61Ag
wP6kJnS0hVUrp9rtGT2el/627Dkhm/LW5hB7pdh3ewoBn/oe9BPrOQlJlw+pYA5N
Pb6/LYN5jJ2ZVl4E7YlQ+4On4yg4d/O8BjtHoBjDg2OCrfgteEYrmd3WU1DpyJoC
OliqFd+k15Yb9R6IBa8o1m1Wuwzw+l1tHmPexCdYJJTUe9CNEz2dOS5aDNyjLnf7
/l7LWwYXIufYDSvvOqtw/ic50Nm0ayi54vMpSdHbw4gNAh2MofF/aImv9/Q6ooY1
BsqjT+CAIMHCLNYNHGmnVDPQ2G79v6Z3Pj9ZMXZgeON3xx9nTTkdqhDqTGlWRl3p
kt7mLlWzgeklKXucXbcknY71MQeS/r0EwQFs10c1KMBJ9iw7p6bS5NtGHfeb+Dmg
9CURH3lgedt0duJdZCi6RdRNs5ft/RqYfhqwsTu3KcqZp7zloTgOtJdfCooMEzYr
pPC79O5RH6nEW6XSYQ4n0DhZ9hmLpmKbrFIv5Ee61CFdpi4b9FICzPMNWMF9kMR4
WtHQrUqHV0Hz92YTG0RSKs3MOQMe/KjQMGlu4tKVmNFcFUf10ERqmu+JHjBdSF3M
QjtrPlnGCHX/rATxZglH2/61y6TWk0z8rBedEoi+hKGvqZUym096CYPWMGqxemkr
mBanNKO7+mYz+nP1b4PQD/pUZiiacUyjEHeLaEf2AeWV0vYrpoxet037YJ0U5ODc
7lzdntMyzDoomhaEFnt1dZh8VsVVN1EG64d7czfE40Qsiqiq0R+OSHbgoFfpzsDC
7EuiqYiRG5LxQWuyXU/r456GESn1e0lbCe8F8o9DJJp0HaT4zBMMBd0kG2ASPdDB
jri0frDFgDwMj1aCeNkls350X+KQwU265R1rsZgAzhtnSyyEPypTl7I0kE86izfW
FI6TXnhr5damngfvEBlVhtIwoMdwCm/JRfTQX5xMMDu4TFOXFreyCYvl4+P6G7pn
xFK+G9biwBd5VEs7NB9q2PxECtUaFTqrDalS+uLHBogpKsuGecSt0UbWedc/4xB5
8syu7vmajm0V6w8ulcs2cQlvd/6lOHs2rqTCH6tL5Li1kkyvM4sfOhUeCsJQjhhV
+qGtxhUIzZG5Ip9MMGdBaXjyyiA6YQn7lhq7RsrAKfD9xmWkR2FPUPOdJPil63RG
vK8nfuAyuu+OodHZXAVRev68RcMyoL6TJxO5w8q7c+o/VpSZkbtrUgGD3vqX3x1S
5GHP6aw2ZwXswhZJctgBVygZxKdvvHVFhuyB6pMkD4mFkpWbEGv7bpsBWzNp6rcn
PPTmJ7NB7PCMUyx+D8EUjveLuwh1CNKd0xWDKQCURovZ8MnKBO1mCw+tli80IwJH
rPFa+poXRoziAriZFnKspJ06HuPbSaUe2mLdWdSEtYR94zrOJH1eLE9x+W8uJPVD
VcOOiDvvK0Na+9M4O+wPpfRtHGIO1mv5eXZsAX1r/NSivozw+ycYFg9Ao4whBGQL
lfHfErQXn2Ilxob1L5ufnakWDtFCJ+JLvp+zCA1Hiqh+YCqVhtvX9TZcnoDuPEG1
74Sd3R/MMZuw2Kbjl3kWAELyADLfvCP7PGYQKLKfiREh0NGtP5cJf3B4l2EhNqLT
YmDsafN9jVGdpoF8BlgcpTkCgTLDFdECe5hHUyBhPnHxxiU5NtTAIifm1oX59fgu
oeVZK+FC67KwbkHQxTyX5ws++BbkSbHekjAaLYt9UtlvbwOV4th1PIK+QEeVjcdU
hQ35OQQva2mtaZUceTtloAuI3wTm0MjS0y+H1yawZyRCWdemRpQ+exz5ISpx/Djb
Sk4HJTK7xQwNImc63fWHhyhB8OFdC9LLsLak6rjGEi9lpgZywiQC2quIJA+hkI/p
CHOGipux+E0jDjFc6ObpjBKB5D9Z8zCovHW5jldutK3Ap9Ir2ALn/A9Nd5Dt6U1E
XrBytT/xmWIoESp9bDmKUj9KP4V9fMHdIQM4aZKeLWTOnRWV5Bf+7KeMuvKniFf9
Oy0qZ4dOErvF3eRkt517ggTHK1b0ilhq+QG723M7Z7X5D2gbDOI5BN6Uj6sMOo0E
fZNcOXTHuj4tRhEy+qXlOsQhdZrK8QVs+v6aO1sFLFvBPvUOL7laRGCwhYlVyRok
GXou4GsfvNNHXEvERGHKpuQo2xvgmMVmGuPC6qxQMEPU2IohBkRzu8s7L1G5MxR2
vFoVeRgBTSftYgDHmXyoMN0PiTW5MgKhtMSCPOifoBfXlkUtZFxZXLP27KVQJJfE
/3+ez2LpcJGSTe0OMD8+4XIw73XQqYhS5Iu27hfyUBfH/90/Ko0tv2kmObJH1d6v
Mozy2CerFzH6g3FwNynLm7JA7td+goPSQ1+9PSu6ZlwKOwZYU8bIauFOjBGyuz0E
JXa0YXjj3Bg04VDJEcl0+KAHUWbDJO9VRJZ/UPQ0S282FgVZuXKEak5SJX8Hi6io
PIrtZg6fLfhbcLnxOaFsqAqzLNjWkffCG0ThIkl9h+iPJTStO4Kyg23VLwjFPj3L
HhkdcJxiJ7fV97iu/AfWwttki+TTBPCN52WMZdbiNlsFf/Y8qYk4QkTKxlKxqwrW
whn+aHherUOBac+95Rr8pTSaeFSp/MuX7TnUTr0di2HD/bZrlCBZXeHEwFCOVyQr
Q/bDHDPbyg3N7lmf1ODh6QeMVzj5MNX1Ga5SDwvKyLEszSCQO+Dg/ICF3u18S/6P
V2b63YaMRT0QL1Zol3jIQcATtKeQ+3GX9svVJ+RW4hjm1aJmkIYa3plFZXEmXbDN
oR+CA8Ky1t0nq6BFk4e5DjFPpDmTSFbbN5tEiWFcGvnOZcLQZtUrDLRo0youOVNh
s6T4c/cscnJ0UMsHw/dKT+aEFGr+1DNuWx1nYdAe1nxfPRFNXgObge9/qnDzBPz/
f5rwXyQwntMUXJS2hbKdX2IOd/1uULr9blzBXtaMfCzZRSEQtQwQiUFrGrSDZvm3
OPm3+FZ0/qzeQ7meCHBdOJ2yvjq9jygMZgDXh79E3A0XryrXQGj4dtlE8UsAhOIP
kafPkXU9oz5wcdkcqmMdqLAb6+b+gVzi/yIB6bUipbQ=
`pragma protect end_protected
