// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YPDW7OGRu6IMgF7Hctfoc10fUjTT6gmU+Yav/yVopen83EBekRUTBqW6w+5vYki7
X4yoK0hhmAN8vSn5G2KGMbY6nVuI54CUSf8lp7u2Hn8VZHmEcGmkNTh8WNqSaWgi
AQJqzNyK+HN7fzSPhgc24BM4Fad3zXPTeqO0fOryr4A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 126720)
PtOlNwI/cJO2QDrN2qS0dhT5OeDRQgVMeE39AxAclOpL3DaK9jLh4KIu0vex7Q99
2TuxzVYRfXxsdd6Zb29ZPOMxGvXzOhFaWQ8mz/2CPi4s6cRL/gP0h/MEOPsJ/+z1
f2Caa3/hMc8PKWEbBEciPQTgOZIF3JT3nLZi8yEZCi50af1/V7VOVFL4AB+g5v50
8B2cfE6JFN4c5kfVvv8/oUR5FxdI/cvpfttwunapM+CjtKcZHq6N8vHVeF3BrKzq
HdTaSgvZiXNU6z/bhj0A+bfXdZCEWXds33UUosq8CTZ+VG+MuZ8DlCdwym72ULVK
R42ME7k3AN8QgGlz/kHT/BnIPDo5yPhA0XFjdTGJZ90m0AYnxp3t/rNL058PRbP+
+THkrZr6JOpj2bkUKiOXkZ/bYOOZYQOF2jrWAXbtnsnDSWSxb33wFgnglhbRaHLY
FOE9ItMJ96pZDc6WwJ4pceKxjKUyNZHzCgX9VHHpNEug4nknh9HEwsgeNgUXcxJ7
ElYfW2m2PAhxuQjCSLy0NNpeylCdUUHz0HIw9odFEOzb0UzFTWB0g3VZITjbfLFv
q4fCsfqf2UVD53U03Z+p1a/V0HWQOTCHFxIHc6oR5YaOhQOLASD2BTR6D/60O82e
c/uRVfhM+MVWfp5lnWY4gtaWREeVD956DtsXsQ3+Kt8Mar8kqU+yjI6GytJVjtzz
kv/0XquMO6DXyvT1QafXB7d+O6qNIYt8w53kxAJS9T/y5u1eeeidBm7pIvs4QM+l
VVtbt9WM8ko920skUuzxF6WpZ9gfdPZuLpaOzCxl1NMfnQ/6t79d6Xx1Pf1XVJPt
JHiofv7GM4AUZY6DlJt2SAhoS1/TCNWrjTWE3MiYWHWlqpXdUctPYWPEkOaPf1Qd
PrMnBUcQHjHqAWj1ooJGfHhLO23e5A/Vf++8jZsNq+nuZm5R/v0WSsvXzMyU4VuN
CteFnHssFvOsBicgPvJcj/kJPyW5Fbeg8IkUS/yno1ZEQAtfDaCpTwswwqQfH5b9
rDuDxaUSGFNZeL+FzlyMuqhAsmVKGHv6uzowJkd+lGaZ/a00V53y/eYtO6WM36zH
Ie9iL2JWAuy/GYQdGE2ChnQvOvR9n7LrFNwjtrR+4qU1Vt50RH7yhKgR/BZ5SOEd
VrvX72YQOHP85AvuFdVPacCr4v1dZzjy7g29P/Uno2BIOOGDnmb+b5mpJQI+IBRD
6229l/Sd3G2Ew8siGgXD6cv6gG6f1DeNghUnrly3FVgjiuCYLcFoRLa29OYTR+ic
d4VQA9FgNI7iiXt+2k1IwAyrnHEyBAgcHG9xjuAEWF5qZRdKZJqzi5h6XQlUO4AY
PnyfXBhY0XqVuoTaCudwLg9zVY6TDyPjfmWFFTq+5y7S2AQEBUsw4bkXzhZG579s
e5zkMDAh/IUkfJUC/5pf0Le5B0NO1/BNLnBzzGjoVDtaUXdq5stUxPqHZ5ZpkgEN
9SM9gyjEvgHrXu7exCuZjzqiDv6BBa36xXZ0H/IQPMInEhX+3HXnd224wwGwmtNT
ZhquwpUkCV/EEVD10u0Kt52137PrHNF3FOxR9danFr8jGWc+zRWloOzdAIZP/DF0
tUnyELD6foAJwIT7xZWVw7rKQoQXNlPw8lbOl24iurD2/IgyhNixpnMPIHm1ApE5
s6U1JjlJTJ3vfG6IX5pChMHJZWrxcqM2cqC8OC2T0rzD2YzUJc9YrWVYRNYCQFsH
EQmXIsb+8r7U8oLlyECxoUT4OatRb3MSzhEov+hy7iEGbJ0gubRzv7354/Is2mIT
sAsZWCtzbWZ8AfweSy/vKRQs0DKliPsIQbjMprRfbXxz4LdJrvw8hOwdBabOnLDq
k/ug4WFsot9SHl0Sai69CNK7cGqxfz5M0apXd/Ajt4YJXkYBo7y8Y72XUyyRbDcO
hg5MV5VJmkZ8xN1bwfMGyfY8HJOF/dlBwfuh7IOgQF/AuvLIlnzkyXTu2ngzZguW
y3EMGjY2E5zrbcZ/XYsbBIiSMvichRfPrq/edbvuBwdESAyrAM+lr2o1jA9M866Y
UWKylnkDuTNvq3KID+f0nXmzzmI/JUBYtA4DZSCa2YLl5x9bNZP1PvZGJObnVuPk
vmm8JP8yX/Pkmigg9ARe/8BtsDptK1udeTStZ9zYunChHMx5oEGBdc5FDppF3LT2
1l6ibVgnKJE+Ubq12MPHuVy6fs4L20Qh/aFoNiJ1fjR4srxfwCtH1RLM2yQdaXHC
bkF1LUyA+azUoJUHSbaQBd7aA3XGNAKzCYLj0121IoZ7ZKDnDmmRZODNoMbDcax1
fm8ymw0dyHoZM44/W8yuK7t8UAX/EaSYG4plw74H4smPcqFXzQF/0TTPs8q8uHhG
a4r1ou+fuk4cxUFuf1L5t4sqVqEPaVcQdgu0VxDO0249KyFwD3zwY7kqGeVu+/eq
aRmdpiMYe6Vvawdk1XdmURcqyCLLHCNc0BpuC0BZuN7gSL15FBlK++6DhtiY4jOi
TbWmj1XvWASmbYufKKF5Yd+iZ5wvoJ4U04snypCqyRKE7Qjw0Q+MCdRa28KayQhh
t1qDopCQxXxNt1oD3wkWdcBDrpzHCzlz0JmBxSQmdiRLpW4j9CPMhTn7Pl7Iwk22
C08ywQCfTpFSWEjQ2XF5rLzC4KMQme+8PYKenXFmd7eSSexX/oc2KeMoQ+z7sXX3
l0QkTVqViT+nA1Yp8LiJY2XP4uxQfQ7+kZObuKnjzqa5gZvOz1n58pRZ+g3rpQzM
0qpwSZDIYEyNJWnd7mwV9ELbYR8+tM/Zn/HfUUXyR5DHFb2JvCm+vJzf7Eyy7tyh
b4HiOzlCpUsCQskwgZ5STmFb/6w8TFSNYKEJCFlyQFuFXr3687OEp+ndkHcnZ2Kq
WPdP/n1kyoS5JFP05XkBiQdPfo7AP3Ddrj1yKr2koNcMzJw+vs60sMP0x+oULsgz
pjrkCTXFtep0eiBXTG7xvifC0nRYjfhb7IEBbA5eoT53V4MviYD1KSuv2rVEaUox
v6uRzkCn61JeTzaz9OnpmqVBXgsI4VaL6mG3b9MtSIdX65dH4WXUyGz9wx/d1zp/
hrhka/ONN1WxOKv7CDu30hE7tNjg8+cGsBMxZBd7f/6ECgXQmmRpLMS+SOeFAyuY
a82xPwR/PbsvHXc3MtIEzTCW8hjUC6Xn0KFNjhmmCK5/HCwjlEKHecL8d3F7kkEL
6g99X5j/Wfn8Fl/vNPokJjhAvgqGYGW5fE2NU9pYgwU0qBSVVQouYpYCpkFETBqc
R8gLe79v/EOum3KiLNxbrRrbCQX3BffzGy3I9jYwNCBvgAZrdHZSFRoGErPovACO
kfjcmnCv4obTUdJppuWEAnCTotcnm/ACZ9YzivT41pne6hETdO2q4FJY2/EMB07F
0xrrKGvV7iNanx0mpn0NbWTYxaahaod2UuBVfJ7lekkU/PKyDnafzecbT3oyEBVX
jGSBumJcp33zQEVFQeuqp+vvwAzwGV5664sa6WxXqmm53MTWyafHZhtP6jhXlFHK
RjU8zQoJICrP2RR8pgksDAnmQaJw0KfvGwvDCJdhRwcZRDT2QxNYfqf0Gevx/GLv
A3+4E7szZHMpYrhP1VZ0xmr76OISaqNU0Rw58ZhnBvtlrTQ25gWhJNpOiBcgVz5h
Sph2RFQPrVRfzjLCqPOuqtHZAplNMj04phjk626dWulth8AFCyWqA6eH2z5Rz2eU
uJVBX+xWelYO1kMI3/vvWR0ZHQWAbwCLFTzZSHe/fEBZtxiFqWKaj+F9XdkFiZGj
HV2ivC7VFH9TMC7Ed7nCfK3jJmgodaYtrAuMRmgXtee15H8TNl+GBGUWhOh07v0F
A7pJlevYaZQGDLZH+8sN6sO+ddinXbWQoN/rS+Xbqup1nRd3YZ9zVNX2OpOeUtLS
tclmU4/aAi+Tpm+R9f8C7qlzJgvXozHneMIUbijWcRo02g/wvK7enE+2Ug8msDpT
HwXJD11e5ybOIzgM5dxt6aOLru+LYDW+5yGckugT8TuSbzTybk4+huR6C+mMA08r
ZjZha5iBpk5a7wfJRFYJxFj5emJPv2GA2DBgxEbSuEjrBWoFwqyc1tN1JBqM1ufH
vOeFFv8LK9Ao/6mRMxhZdSgpmcETE97ie483lC6qZdJm5vGB5g760ph5iPf1epz+
7kWuewamSyTOczeI1X+zV+Ew3Zd0cpGYjbBmhKIZqE8Uu2RoVaxRvPcL6uH5hy/L
eDsEZZwxx0CXdGeGS2zNpp5jLoMY/iF8mzUe17HDpOPvSZ0ws2CHvSIARZcyqvm4
nhi15pGCB0nPUiCb6El4qj39JQ5JE5v6+uktdtOyK7ERKh7EuWEnIV2xwsbTQ4s6
Rju1HVPvDeeYU7EnfFGsh/SVBa7Uyg3TSt0p6g6DZTyBg/UdB+u+zEJAEcuBgbwS
pNoPQr1Oa12kadQ1HUD1K6gQffn9gVf9iuDEcy0oRmq1yqR3xTxFlpeCPvDyMXHQ
2nmbykUwtvItsakEM7Oie0GyBozwGqZTL1w+qVchgYpItZzxtiNBbEt7pXsf228j
lPihBm/Wf8vRLLpdc2c7nDyKF9yxtViJhgN52Ivi/qyHEGvv/3J3hRJXMK8oukBf
HDCazpqHg4KCrbQQNOAxS+Eh8gxhupLMu97UymaHMqeTgkIoWBmlhMKoQPoLtO0P
KW8saCdw1mjLyXG6h2E93etrMWA9hxAIJ+q4ev4AH8uNnVEbDVyfNRcH8zNm4dWm
ir9QKV7Baexj0+Dyu/x5bRRI4LSnoiY4EXLqO679rUCEuvRgXHfj9uiJ+6aFkuvo
x9/QewWqr/d26+Rtm6F/ovD91U4Xg7qsXAKo9kftH74P/snUEKHgIqUSc0jyUPOy
n3WhwggqQjoMJ43hU98qOceUTG7Yux17JzbOWr4KfJqmyQB/67foOtJoLAqNk5Gd
/yaX8eS+N1lRrosY7tRWn9gdWmF2lYZnTFV6oILOgeDKjmTwOoQJl1qie3VmcCpK
RaPhKlvQuQQCT/Z3IDLrQORVVT8rbCKIPjA6hK35OkpWHx8tsQ3wGdRQCHSTBHtK
eW5VSMb4ALTonh6Y90G1ddfSCBC+Kuj8X6V6EFcHE3l1y2zAEbhZSK63r+cNikmy
4ap6DdUVgXLFwVq27CuokbNPgqA+q6nur0yl7XBC/iUVAnmEhn/edEyDDxKtEknb
I8B/4J+qssq/iRZHcEcV635ay0/ukAFUd/oghTz8QOqRS0lKKHCNovyxi4ayJBnM
Fck77g8ICn4NecGgTEUflS3zH87ORbiZn8R49Edl4yghqK6kirPFXirYwuQUFhlj
aTHJLFvwl8cQex9S3xFBCvhsQw4f5l0Px/RQSdrQRaWhYrxdzGLbsPNcQ+/o2uxC
ApojD3n9WaCdo0ksIKamKV/omKAG1EhSLQLfw9bgq70vtT7P2t0m/9653gLlWS3C
l0+2/dMkZixDsZN7WYdOio8wXRAVL6NMAO8Rg6esHwbZ4ej0eGYLDI5dkJGC5YD4
Fxd5zqTNBhrbpe2slh5GjV0lvfDzAgZSBrkHbV+EMbodSs2bO879OYtGnkOdiUNR
C2/jSDcNBWSa01vroa1QOGLISDxUjlTW1BmoIbbHkPHeU+izGBth1Z+IIpcURHY2
aHA2jIgFqcteLJO02O42igFZc41c+mtbq66VRpob+oAo1g3670CzaKcNTJhFXWk+
UCSucduXv6+4kF7s/9vhAGTZJS30vnznvk647m16Os1yBj8+s9RWpZk1Si7mW1Es
UfruR4WZlayCJ6sGS48QkvqnBJPAYHr8uF7D4MxVXxBzAJEIsEXzHRmPE6J+Kc8j
MeCXBuQijVq+meN6dp168vT/MkrGMtVpOYWgBKO2ISO2G38mvWcHX7Ttx4VKi6i6
sP48uS1ITRNKM+qIZzxlF1/dtWmS9yJJOUkqdQBEjWc+Ol0ch0Ql0K9bHw5AYQbx
fztxu1ZMaI518AbB/X3VjPf1RH5pvVaR+AsOSpjrlS19ufqArgRxAhLZms7OBGJt
aFjZhrfPDj82WGbfi+OpFK7um6vYBnluQEOE+f+cyebLV9MWWKTfgCrlHZ+kAff1
vJqEYcvdOTobU+UAQV29ALFV2+qn7Nq/mcPAjpxzCV+YsyAu+a3DsIgMaUmXQLPn
/0ZdIBHOJADuHsNVBSvaJ1z1pMt/+Ey8iUwbSe/7VnireaQR+YjlVoBiUKbYbN1E
m+GJZ5bb7IIu6NB0RsJ5ClDIjbMkH2nzL0DMnKWedQ0ip1O02YJnOEE4zdB1YIEn
LYp17VbGjMWal/qOJ9tejQ3lw6qeX2dGrYBWQW/E3RLChqB7hT2B3zfT9kZDro3F
nBEN4950oDc0BnGm6hPi6qyFqJpoQu82Nta3nmoKnOc7nTacsvCRTI4n791GY9Zt
1pFnv9+6D8u7ZFy9+d/7rFWQmUCmA1dAhzVAzpZxVTy+L5hQsvldOdWs7bf9iK6i
ZfQG7KGsvZfwhlJ6ho7ppJLWmnkHokfzMoU+jTzpq6Wy6FrQPf4+S6Sz7CbtdEnc
72M2ze7eWFcvnQFOZeZEVqYxpgZ/0Fkw6nBkMrhoSlNpSkbav66YqdmpLyiTibhB
vydsaVw5BHPUpb8o7zr/dcUlkBBN/wJSLPnR/f3UiWay9p5G7j60sND3r00QJl7R
ci28aa1ZiH2VdruwTkPP8DfN3b5UmvSRSscWSZpK3lGzZKyE54Yf2fCZTJk7IJzu
jziQS48gaLWk2UYT2UtmDsVY+uO+Hm1vvEQS4ZUHU7GqqTq+pUTdkgo4ig0qXjWo
HWWPxrIFMspO+lZtBbAeWFWMXtL5qGy8b7t5G75683TPRYK498it//eM9BQ6Pf1m
kyfWf66hkV+YC03XVZQR2dv4dO3yfyIVbZxvTZ5buKrETbc+VOjN+E6OyyBVtlNb
zM0i8Q2maOivwrgxgVH02EK1EKCDty9fzqYRyMtE+SxraGL4FJ3ju176wUUau2FK
bHF7YWlN60f0tode/cFWiEKwA4opcFYvpH11s6Fp5BAMvhbTRCQEt4XYE6Ss6b+r
fueicM6kmGCOSdunWFNJ6WL8x8wb35cAT8iiuLitUjhYZ2dJi3FpOtO5jz/lUyHO
oYNYHPLy4PpSbM6YMMEXzL/NBNf7PPqCgAq6A7UnidcwpGTjTf/pJLl1e8Derm2p
YjTNrE1oRIb1EEw/6WPU1su++vS/6nRyV7wM51VMOycHVT7TzxTHaXV7qbpZRPDx
yT8Ygn1oQUuMdcW7pgRtgFdBcJyvyYYrnFUEV+0SaNVDpSURgQ64GBFJSpNiaGI/
6EOr93Lf7vvgvb3RJikhlffltVRMDz23Blt0pLjBIkgpPWUn5xaCOLNBJPuVAxyr
GaN5KLD9E/3tny7LdNqtKQn4qeDyVTBweo24X3I6zBr6UK4X+ot8+PLquxdP7F1j
Dq+/7TX8k6cwawXodQI8sX2syVX/J+H9CQ0v6TxHZaxvdAiZrf3WKiJhQ6TM9J6G
EMJ2Fse5US0C+7NCJS0eDkmeuaX333hoD/QOT1yiDmT58ZiTcmf29ri+87hSLz75
uK8HM9RX3HUHizQXdcnfNc0kqdHwjvkLDUixBEOIqdHFMf586yfsWph54SmWG2kL
prQubeBygSTuN8O9gCQwp57l1q+Srdbhe4rGtNsKIM+AyP601x8LCszrRaokXIqt
GLDjgGwg8/RXd4mbgfFA3PD5SzItDAn7WTNu34F8ChXZ6WL3qZyh979Jt+V/HUOD
BEfUGCWl4fQmhWt3fUVgcqdlA4+agZyOQsH1NT9KG9FjxsXAnLxRYbsMSs1VmcaJ
DCc8QHMOySHI3UeWgzWEPoJxWChefl67/A4U07J+ge23cjwukzgXdEld+S/+IatQ
TgkMHYqNOiNhuglph41GaMmhWEKFwaXcKzQeesaV68DeahSoHSHcZh8tSpoGVE3e
culhaJUWYZcERWv2TYPQU3SuyzwyNGSN9gL0td+Tg0vlOM6h/yl7EkTZVOPg8Hvz
nvB2AaRVsdoi5UwJLDkGh/B71KgdxiwtzKgoFjDe3ih7oLSKSaemoLekDpcQMfXT
oBxrdlzsOm0RPtbFmUhA0uXEM9Kr4wMLaQrjSyXyKLbPwOIuSH0GkFgSNZjJHAeE
9DTbupEl3R9Y1GIilC9UMbcKyDEh/5NNnLj69PbhI9tdBVC/MHlEYuT1zZqrbCmP
jtFGRErkwYSjOoYA/Fy9uSh1OpZRWI+DheEWBUAMM+B2FiimbTFpHnEkUH5BVg65
VGYJhUhzmwEGMZzLfl4LOeTtueLwvV4ihX0wPw/tuLgdFoMhmKdnFhmG5rQE7ymS
c657elm+xqrcz3G9yGsdMGYwBVaHQbabvC2+5ZrAbtz+2AZYZDGzSEbEVeRuUbdn
skb9Hnq7BFAl6QkHFq5CyL6V74XjYtNi9ACZYQOdlp2gqwjHTUXtdvfw6OaIu+8H
vjCXHmlVm00PoooiNDWYs6dcbK+w2/Bp5G9lcrMgRCTuFjHO41ZpSbSmo5S9r1j2
VG38m3AMRGu+JjiFf6hf19nVWSwv9G0FbLYM2t1Ulgl6R2LaPxjxuG2yqIUFAoK7
zm3DuHG/jwYgMUzrk8wp+jnPnJeQWGFRbpT3WCYRcY5/6TU3PPHSIiwS5elN+vKr
HF9t6D5YG5aTZ+gzFb4KvYXAGbgrirSeE+1Cyu+cgUap4XKmkmHUVpsACxg00kbz
HSYG9aC2Rxj7VUnN2kB8EK/ljA2y66rEC/tykO4mXw7bZqUc5Htr+1rPDEIqUXiq
hudtu/jqry1jZOFKMI+/QfejEiI1GtKzlGnf++Q26M9KZlnSqeJE7BYw3cFDWqIF
Br1PVD9Qp4c/v1DH9dJbuNEQ3VRC8MaYMUM+i6x6/2NhGw7fRB9fLLL6yF+QmS1E
gULxBNlU/VHEIfVusjt9K/uMK7Fe3smQEaWV8HgH95mHECcWiBBHZkC+B7qWHGmk
dhUn5U6yPhVsGpY30rtQnf1YubElLB4+OuIeCjyVqIM6dPAjGU8S+issE1PNLZr+
RvfeET83c0KeqnWwdiyZweP5lFdYzCTs3LaA+5/TTYHEmK0lLLTtbsJiM9Ko1l3M
JB4E0cN+ppKRXpPZxgfefJVLz2hDQJNeoRGIcYjG4gESmFpHV9ymOcExhJ7Vngyv
ZPKK9dfU2Ewsf2s6m5C0tGxUqXHVXUGfqTefvvZURP0yiCUF54cRJTfb7KZrG3tq
6hnnwoY6Tg+esHI2TFwGdX2Yq+2ekH/+O49c2TDpSYcpEyLff5LG0Cr44iaCxFpo
YirzX7mldAQ69juCTeUSICYrWaBk8s2VOy50BqheD5IT8m5pGM0AUFcjN7nomVSv
SexgBDjjrDi6h9Ag36LwSGdfAWuMC4i4Zq9ljYdRj54nfM8bTUc/32/hIgMHCre+
ghXIHVJTVSk0xiUn1T/YS3UnnMdzPV5uYEAumjse1B4UXDnUBIYBDLWWrODd7dmT
wQKNbeD8bfDlXUSNAy51bQK09cYSZxsQRZYzSWxj2/6d7v2MOTzNsVMsj4ePkQP6
G7f2eqJA90KxyjHhOnJthrhn/93RW7xYeNTBp9qNJGUSVvq63oasZw6cXVJccHmG
cwWRpanPg8uXrOJtpotKzn1VdLWvADCtdZ5aRUKpchk808C13VRrwSzkkXEW+75A
1ruqnA9jD4+k1ZNlDPaoR6oTUZwt+Eu1npgM4II/witIWcPbJ/72FOZbz655JkxH
AQueAIeZAIkG07NVjUu2LiTKpJlm19GskmNJTXBrqS0w7kFvLwKhVWoJ42JLDUMi
MrQoVtOKJT598Gb+JSigvBp3TDcI//4hkdBdCo0BcRHPSmTLfbzch2XLXlGYZfT8
/bcQ3hKEBrR8Fwn0y3zhwKlHbOQ12HAPr2SQ7+tbFYpiy5Z08/kGKG84UXbwacGC
ms8xfr+w2iRVRDr5nreMBsFllMz7c6o1KoxKJF1t6ZnYRV8iwPuzU3KdfTADUAdK
iLtSqFRyPRZRTepBcqiTLhC4zbWVo6KMuC0mvTnpE/yUXINSR/13f5tbmH7xMuWB
q6gDZ+rQQX4fZRmvYB8qRYoFVkMbFIRm/bQjjdHf/tr4qeDcvAO+YX536VtA3VXe
BmsphPtdbtp9TSHuCtOgiWsc4NAZyM2o4Xp9iXG8YgIBrPMA9dQo4q+u+uNrRwCX
9VyF++qgQmy+FjOSV9T7/g2Sjdww9PeLyP0pyn0vMPwn/eJ0CZ1oY9Zh/sluiJX9
KSF1R57kVgsK1c2KPn25fQjRrrJuh7aXkaYIyq1cxtjKrptHr/Q5VG7a0KuVtnrq
JA0Ak1MrlU3OLI4tx5bVGWgF6+O6G113SuxnCBJskOaqIklVWhV43MgmT35VVreW
BZyzEV7NLKtl/o/74xMHfB68WPWAiESsEIWsb7CRxDkkf6PKE8/uXKs3EvbV3mfT
eV8REWRJ9famdHTm1se+xtgRUz+XN7VuPCzI4pojzal6zI1+Mabr/fSYJvr4u1e6
EbEmqXfQaQDv8mFl9+qFf7E5UBy/8TEkfL4N9GqB23aw1VxEGEzqyjWMNFBIS9QF
gzo8BLPRZcTI6qg7+20V7Bze+i5FJsuQ/1TWcaxygtzHGE1KWd5kFcNgus+10RJ7
wneutxerOUmbLzEILHKpxcZdP1AEkZkZcDBhBIvS3FQerHF/ggBqWFSoLYjWsg0w
sdktoEUCuBf4JU19hb6Br17w/8iiS3pWiTfOy2bGNb+eVkrUk4k4NxHTz4CD0rJ3
9MVPzcMtpgLqiMcGFsv3OEBviIDnx1wMvwMS2GwqagWQ5jQ+B2m0aSPSeY/ecRtY
lMuL+xPHpr2xyjI4T1ROCj3w1EtWH+q0uy8n9IAKrmJdsln7MZGvuGKYrBAF/+Kt
3MrkJkQm/j1J8QC4nxCyrooB9nSbaQf6m76NWsuCUqj304hDNC4wQNquEnnHQ9GB
yhtUM7RDMcvc0DvrqzOqMQqFt7NYxQbwVNMyFLZj3+ofa5gHxci7f5z5DMaD6b/n
GeTzStVaDKqyNjf+SR6aRllpusbIp1ZotVPJ6P5f+zCSh6H2vl3R9JDmNi/LEA82
8fQULTyuaK10i55UEiyK/kablY4MkiFoTJc9Fg/08iNceCS0Ge6qxZRCKNN6y16B
nQX2DpU+Z4Q8jH2Ig74wbSftzFCmF7ln+A5YEK5GvFDqcnsfVfuKrDTzKzf8Pewf
Vxd4Tu8TTpxydNhwiFyrHqzpNUPUptV9o+mNDFffr33ztD3siAnggV71//Lj7409
IKhychpdPjwYpeblVXXIEKC3+N2oguvx4Bu3/rMwUlZSduv+QOPSN4bfN3CX6RHc
F3gUiFlzI4KUEC7+QRfVEtalXjA1Fi9aeuJCMZNCLh6SBnIM+Nta+BlfFvfmyG09
sr2xHCW5L0fnjM0dhzalpmOnMLkiX7DCUK/MJQnnqRA7FuVASTgS+WMpEyWaGPhf
x3PNhUUpc9TTj+H8Pgyi1RG2PRqGvOXYo5M7U/EJY5ORE29SZpxmGvRobtY0FyWM
K6DyuPSGui1SPX6OgOtpBXixTXBnlR5Y26L9VFLqio4TbnF9XRz1UWCf8rB7ziXs
bvR4oQrMRwih01gSyjKq0P9nwXwiO/tCyA7UDEiZbrLpQor+d/i880DGsqnf3xRU
oAU9Ja6eB8Xbs8VeypxMCd/pMX4dA/xe8skhz45Erb1YthhXKeVseoIGF9RgAaEd
oIJ9BZKoozjT8mrDvWtv8ZGSGEpmkNf/vdo8Gj84ouSYcAurxPRqE7H+tGLniIu9
JAz/rqzBpif4n8n2JD41QeWyzzvozjrr5JgU6JXXl9vRglSQaarm5m8Sm8RU/AXy
gSzDUscAxVwwgfMyb2fENXlORxnCy/+MxVr3WhcWLczx/nEqp/Z4/XcS7fVmkklf
cS7LJWTaEnCobxDe62kgeowlH4iY5d2VP+8WBM9dY25vmf/ONQ6N3fKJ1cFJq91q
QPeRDupT7I+dYHqjB+c+haprQHKMjpGFDeLw4QVWJmoIKigh7D1Xd4x+07Yr7bGq
v+EKY7zHIBwnoPpw2jln0OQroB/C64E0/rhdD/Q7idcshD9vNUGzVeeMZZCXjOul
LorC//ZPpiFkt+pqPLDOI9rFQ4wt0M8FKhhsjsSZX9h22V4jqTHbwF/jfM8w8n0V
WaNzl69nYa6KETopirhHIThBgki/0z4r7D3GAPCVxByOkLm6lbfi4FZ5hYi6xQut
cV7WpunfGB+4qkOKz5PQpYQy9s5A0e6c4tb5HkbvMpcqer0rI7RZQivHXxJizw5w
oMV2rk59gx7N3XgP9v6b/0Rzevfs1nFt3hbq+i4CPpW8Kz8m2oo6F3XbAOT444+R
/hC/QQ+CY3d4VXNHHdFEcJarErW4MZkmpekV4x5CPxJTQFBkZKQSdm33FdzUQsAI
lENeicLEUB4Sf8ZerhNHYZJbLlOQnytwtUGWtttDxv0mx6cM2tk4430jQ1vhSn5e
Fdrlp2uA63eVhYVTAW0Xhp1n6sYpHfCLQ6NIrik4k4MCy6Gld8SCjTVOYinsmqvD
6IAxymB5HTe02YVUpEyDCvd5Ui9pfpDLCqBuUvj7BHrcSJKrxvyE3beg6NQdNRkl
d+43IPu6TIo/9jGINhd3GWTkIOxzkOSPYtXvrEhMow4IdTS26Xi8zB44evWgZIoz
xfnSJ69Dl+wqt9iumSJ4VbenHQDgGpmrabLHjIAXi68z0syQeNEmXqOd3D+GbbOH
wpEUFNkq8EDLVsZX9Ap3FM2mh/qtXk3aHbiiWu+GI9GR0updkAWjWHWzlP8zI9cZ
tiquBYCqNc7VaoEXbUxhH/Gic4DWVvznwS+RMI7qpom9bSjmDOrCYMVPx13JmbgO
aQM3IzXcGDJoUIZ23y5vohR+jtEmne2RWxIM+DOdB/CtpF7dTVXawhUSLTi+0PoO
B4LBiX4JEkmeh7pEYkpQelZOdoNszFrM7qKGTrv4H2nhdJOhRZenQCmO2cLfxtQv
/rEntENJR81BQZ1o/iTL7PWIkcrxyLpyOBtPB99Y2qp2JIGpEKMdO5oWQ5c2i4Ul
UqnamPWqr0YsV0bNcHlHfIDZvKX3PBumuG2oX69xUCQjOLVwA55ea38yaPwZu/1n
qFT9qkZyJa2XNhddSn+B1ZT1/eHyYxEMWGBkYeb7yDbc89QxMmsZDLZamFGde4eG
xXNYpsLRiqAEvE8MNn5jIfrp4APwdyjjfiacrO4tMGKX1Bz1Ms73HOAvvtjP5Fy3
4lvJ6Vr/22OkZM9ID/SCwqfzq0+bJcg/sgTokrNUhwb9DNAIdoj8xbFS0Xc1zvyg
zjZ1EIPl/ahAP/iB3QgKkiRmmD0FWcUZkR9rZJJHGYPKjwvz+0hW8Ug5iQsvZQb7
0U+nl09Q5JOPMEg83UlC3xA17ww17s43DxcW1JVWrrVEJkAlI++F6oU+4xJziUd2
JYdkubv5Wh/CiuXGOSh6EtkhqGw5NTHIPRR0i7JTCh+VbTzn6Ml/9RIzH9prVY7p
DiZ21bis+fFP0B4CkYexXs0f1bHV2SJthOSOa9yTUNvhWaSLlyDOdG+rMd8mu0pK
zfxW9pRNB6/fFV2W3h3KENPrGDkh/V9u9yGawywgw5m/0Vf/zREksbZn5XdrLioh
+ABM7BQrXo4vKcteEE/WasGWxO23urUhHUSeFuioREKBUUSvfgPrsuAcyeuqJiW3
ADipJBe5/He5EwJtGs9BrdM15w+PKYgHT4YYnlqfxHcCBfZVt1TsRa+2cpiHfcUd
EasGo6dl+PJImd3bWnqW02YlOftxLyWPvj2CKv6moQTRVFuiUjDs13+rVrVYMQiS
FqJunTIvWwszMrRlibOMBQORviUevVuTENuejfa4i7+/+tfOgtjfDCq8eR5lkXiB
s6fhynA1W3vqGrzABAPSlJ4b8ghaY/O5rtihmWop0X0+U2+JBQpWaEyS+gudizW7
M3GcYDlD/aN2tqfZQtBrN7tSnKnZ/6KHBX/13U2clstvIMrxL8srGaE6xUV0ddTP
VDiufOAAeFoVjuE3Cz+q3nNR/L9tpD7DEHf14BL6f7r2zk5Buc6df4QvQW3/dAi1
GUYMMivghqzMimNfcgctjR9LnWde/vYO+5rSkQOmtuC4F3FaLNvA73MtBWAMGpet
mwOyugJScQy/dW7SPDTEsmBEmHSMQPEIMWIAh2LyAp/TpWbD2yT1xG7/ir/EZf2Q
kjCu9yH5KjZaEJeZtmECAFFbr3gxpq6D1s/d+W/3fU3RPvMu8CuUYNNDaeZInWrQ
OlpGBtsp03NeTQvKAFaAfOhF4li3ONyqZzb2It6Xxw59CQ8IHIXe6HIFVlx1hImR
3PR9z5cEAitLiJc8Jvh1yXACx/Xblkw4JlxcUw6oOaesgTsD+teAk3e2hEk1T8De
KBfKlr/BCQW0SXNyrGa85pLuU5K1qKH1gzLyWetfADq7pnUSfO+LFf7AJb4ADlqA
R8rzY4ujm9GswtnPxg51RZ7w9E6kPQv1zvUGhERBgb7C/iEOLTT7CWgDH2LCzfam
pGM9Lv1nxUXWqCuBwoo+unchyAYtoFXuwkCqwNr3/AvvSTcnKrfIIybVeSCde0kc
jJ3JFw8o7ZSbuXQajVahAkPk24XhRGmyfYe6+ABxLne87edyBHNHXa291UoUH1hX
8a+gbMu1MkKFyJGWzJTrBfKWq1Kz3vrlvQ4B9Z4HAI+N2AMB8oyzY1LFoy9TbLzJ
hjQbQDaHWnnltH/th/DYdGRdWtPoID5VWYJI3RHIXsURJLJUO3eghEPOY+M8R14D
ixvcmbZWUDYsJaEYi1KE2moReKhBiVTrST6tBxyGgGLCKpBpToEmwkOUwAfVMETZ
T24/walw6jU8ave/LzYOeHBdr7gavG+CJUK3w8o/y72X89xid+x7/xcr6z5DUNQ3
qFf2Vx37UupDdkULGfDVMW5czWJCE+gQ9/szlIumyWW6ql0+fcTZZXLF+6sAsCbB
wa2TgHAtCg2u0n5/Pdrl63YKo0ssQC+MJHcG0nB6CjMIfv/RJsVYG4KV+BBa0V1K
etsc9u5gBCYXyNT4hYCEg/XgU3V5L/Ibaeot6jXh8b8yh0YhmhJBJtqJzvnQs3Fw
ZGyEFtH1xx6Qpm5utb3U2JVIsZYv39C0GyIzJR4hwiGDOa29TxDnqOBDiBMiFpKJ
0ilp3dJO4f49cRl+6IYXUdrQuY/dlPg4gv/qIYiKcj5c8ZTdk2ChMe8yICRRH1qa
KRT5KtYiDaC3gdtBKf2Hka7upRr5AGY6Vxi69ez3bddTBpIc8bAA8qsOJkMEglgO
6uSPPxFuurZ/Gukcx3Hocx61Io3b+c6h6rrlz08R18gmlRjlqz0wkWfu66RkCAjJ
w5vr7sOXnSPHevb9+fHFa4I94i6do6gB4WGbXd0X6t7LYW38gy3Ds8K1kno9BNC3
HImoHy/YOtEWndwmJwLvpLINSDs4VRt1Ia1DYJuOSYHs+c46EnbpAvRkT1n01Ljv
JYL7Ia5O1Ee9oiHyQVIcbGnSHBVSkZRvJQBSnj2C2DsAcpJ2aCCrUlpChKLYpkfl
IVbwNFQF4Er4yFE6c5T+w2GeHzR/7S0wfYJyDpBLkab5bNhzvByQCbm7tPZq0JpX
sF/othraZ2pce7m6TO6ZbYnGCCeDRXUp+33oExhRunHPbNpw4YlrTf7lgTqc05/g
C3k+t9BpigTDYR2caZfUM4jazEoofB46mSy9thg0VmCXKB2/XX/bCuX2S+P3cHas
uMntSq04dkalrT8HCLqnbLesQ5/8GaA6X9LMgIRCDizVtjqbHF+9zZ0fUrE7wTii
0hnQCuaUNTXwoNzV3tcXvJiJTqdoV4iqQ53i7FcnZH3RDb+JQcEQl9SbBbBPl90b
q0Dy9EDp43XcNu7bJ8S2Fg0hulHw8tvvi5c2nwvKqUPF6J0BmgmXPdVJOrZjBHm8
FKvgZdzn5ElfOXBSxmJFZ5KuIuGB4ZR6PedH5cMuY1lvgbvyh/A5yhb40pF/wYj+
XMfu/vgrSfhjOTccjRLGqMX6z67IVb3bQvir4ji8LorF8iHX1TMaBxzA4T1j3gf3
XfrAUFkQcmoISIQR0e70HF8RndNU2WfYfJYLHlXWbKoUs3778y3SeBEP+Do9likd
gYzUTj9Ydksg/BuOaPdvi8UOCV+sUlhxhU2QnvyVk15KSu1afRpVxoGlp7WW/8oO
Yyhh8pybKSV0uLOpMTYrs0ajXzKYaaG0Uo86l5XDgggaHIE1nMMkGFGCwX9jxrO1
tP2aJxdZ8dbmKDwMuEECZHowYw2BetEOBXN3EO+YBjn2c6+avMCUvEPUE6v7tuV2
rmFhES4yH5SI0HyhejUWMRLB61PXdA09kRNZb9b1iW0xI0tggE020RG8dt3slTqj
GNKeibYhwk93gx+D2cPJtZQjaF1hGnBJ4ux0P+2erQUi6YNKEe4Dl73I2UJcoBl8
dcrH2tdJNQL3ljgfKN6bDYj4RJbPBtAh85OQIlEvWFvfSV7yTg2u6OX0y48pt8dZ
EGho9I20X9Z6+useigCeoMu5HKMP9wO4dwzRvT0LJyRpaDBrcKMg7DubI5/MQ6co
RU0w3lYcIDEM7mnhiJEn3WqPvQzcYxfgXwoRC18fCnH5T4KVWXfl2KUD1hT8lgsQ
eHDUFN6Fa8yswXQAg0WxXSaj2w4xvK/xB8+02be5NBZjkBIUb0OvdhRXw5lpaKrt
uDhjDngIvgE0OBfMYFuNBIa+VZuByP5GPJoC8Y1caS2ExHn0W5DZdYYN9CUy7IbS
BVg/zPuEGZtCxDgCee5sYjcPg1cW601/MsZZkx5SHzDlH/w1fzBhaZ0znKWOANRJ
9DYBl5Pi11hzSGzYHYVH7/m/lxGQruADshq+hgzw6raG1QErlgyyPla8EehEedWe
dROnOC34AyVOIYdrquM7FrxpljYTB+Li8UueUBi3S1M5iwXSk22+JCR/USsHZ1tP
hkXntzcz5jLLYSAwzkKoLXu1xXeTZApTl5OIXWS1/ILoASmzj00TSQM4l0mT91pm
N5r2U1/1PEIEUd7iXtVx3Jf7BuhomysRkbxdlGpaP+Yu23ahrvRO6fUrE//gwJXK
msT+YVqrGEG1/HtaSY6yCizhuYrjNKygd27FKyOkL7yTI3+sqgWHu9wWwrCVfe3d
5sIA7GF7x7HEXwxQ7e1U3Xm9mZa9ESDIj6N3T+9PovXPk/+k32I+QaQ4ngon7ZiK
mdDfYl+UMSJwoK8miNzrtpbwgVXVRusfkYfGxqhGrFMxfA2vmJu8KP4Q2gLkc12N
zBzZlI35/Gghs5eNFxo6aRA9vZVVh64lg6/6luq0pDP2oz/uos9HDHfp6aPXWRfD
SnJdO1nKfmChYhOJkXTzBF1zdboyZAN1ayhSZbq8cWpi8kYIn+C5CwVBX3kKeH4x
e5ieOmpZgtfJjIhJrn2z2iGxdOsPJH8LejQ4e1JZln3YXs7yGqFVllb46soZ91rc
6D3DRKMvvegI0dr8m7Z1mCrOaqboMqZwuOal6zjkhMmr+6goi/xE51Tv8Vw/koFV
sDoUEEgDP9hKgBdHz5iJwRe0VuFTCpaCwCoXrb+VoUe3GnvvRD0iBtKP0u2ui563
w0TK141fCgtfHeIaFB7504V41YbgTfyXDkuiXwZTlmzMicqF1OBDx5qWOSSsI/Ed
RWNS/YTPseMZSx+KXObyCYyaBz7l8EcbFjXbDPCRAElcPIsiPKY2vqnAychK5YUP
JYEvqVJVkt6nqpDhqwSIyLrybeGEYpEL7/o4H3Y/BWzJjQlPmuVoLRigk9h6JK4+
9iD91OiWkYS51pnjl7N8M0mT5Y5xFBnRoM3tHQ+XUHP4F7htMAOxjBqGH2jN/s+f
p35570zkfaZ1v/cioaCdH9IffACO97Ris49DkAY/FIwuczfHUeqJL6pxP9kxFuoG
y/JgmkGeubZKVrf/XDnAC+GyJHXjPC3HZ6Dz5bFLvMeL4kNyNtPCLgejPDiESuSm
7tbszNkSSkAwNGeqIz5NSbkKtUFh8eR2a15EfwIktdSBsla+GMFpAEHAT8NbQw6o
Ps0Tp56n8cL7+zlo6Los9XP6xOFLov0Wak5yK+cOA4tXZi+IWX60ho3mQHqwGVfg
Qf1FB8pTpFdK0FV1257S04urrbgQt+tSwZXKDWhzGp8rTMwdEF+eBGodzHCGvxOq
wQvqxjVQLRWaS8uHh9ILJR8LHnfn3knOyL6q8PuHf/sszD6d9OY51GsQRa4G+f5d
m5LZnAWa1jUrvBQKuJvhBDW03lm1cp4TJaa83eoSRJY+7vBcylkeHGbchLnP9J3U
w5tMRF7Ljv/Y4R3rg0VgfiWaJPBpc1wxx7pA19OfE3ERp9ysBcdETk3JJQ+k0Tko
9CnfglCTVS5tDl5J5bAeoXogBXHr0PxY1UEj7J50kFv0Vz2VoF+aC7YW11WZ4qTz
mmWGRcNKxfmCb2oOG0x98LSS4Zm4/vf4ZXJdzPhNZZt2b28FqqFGgAQmnnOfhk2A
360APbSOhC1Eu/N3582Jsfo0QO8TAuqbKd8M6jDqAzpommDMBpM0Wd30Zg8Ajdgs
iYPRh8xmuYaS/ZYiYnzAvqzph+djFX0xbs2ulaGfnIY+SKbiPUBXaHUMfwOYGLdM
aBgOX+sFdzJP/aael8PakE0i1wshdsxyMxounrjw6OG4E350+O3723oNjww3Y9SJ
iRMp2drMbeAzKepUqLRxPL8/zNz+UYKZ2iMWbYz3jTxdsnMhZtbKjdXUv+gONOZX
M7mRtO0J0d/OZlL21Agw72nyRwiF2/8tl180vYixxW/DztPWtZ/DmoVYflqOJenN
lsn3X6XQaQDq0fqgkvMdZCsRhbxZOU/bYxKC8WlJJSfq0fi1FcTh4aGsAcaBqFAs
bV8xrQXmxY0j+MKbQeAItk4ID7+7akGMm/dO3zllqm89jo1V/89hdGS+b6Vb5WxB
ptaF2Yyw9MSNMKPUOFLYBNPD9Gzj36qMJvr9WS8EtSD1ZZ773hTEckp2KmPBF+JG
x/HH3r38U2NIjsQQ7nYy4mTeG/nrviis2n+se95GaXh+v4741m4DhtJg949WWYPP
BBCW2+Ehv4bsIcERKNI4CZo/axdG8ioytPrjbOy65RswK7vpegY+hiruQqbukouJ
LUpoT9Bsp3nY3JSynz2aM3Abi5jLYL0qePzTc4Yl4Bp1O/WL3XI6QUtCvjvXECM9
mctCEme5tPnlIbIGK2pd7FDDboRmwwKNqkJd7SzBhE0/L9+Lx0Qp6UDZh2Jag9CE
LBD4DRLOkQTFcHwAMpjK4MIj6UrZBDgBIczfBax6DVXkHL7GKoqUBsSIQV+asyY0
Wmyw6psaS2X3on11yJvT00r59v9tD+YDLYPcg31ogZWnLrULoFhRVlCjGktYh6Ui
BQx1X+T2fJe1DNlYGrNYRkNfNuI1VMEZKqpCPAO3hJmcJS3yDRHA6b8yDDaxinOp
u+I4dhuU4bfpchpmPRrJZX1u6cJj2dZrg+ScV4xCc/XaHMzjwW/PIoUG70v5qcVW
fK+Ut+ZnfmMoYhS9Hvu0U11OFKuoFvdSIlzASQWCCZ1cNyoPSKEpJNGXKWTId/vP
WgBtEe537d81a65ugp3tTwOVc7dF4sdSlpVZnLI7cPF6DvWhYm1oszq5P6jJ6G8w
p2vlMn+XzQQ0dpU3oPnAPw6+iNInNZxCwts83vma5cizR+lyqn/RIoEfSH7V1s0J
nJgkLE9CdcFgAQTs43nhYnm0QePyKFbN0BmAB3VYXZ9fSV0+ICvxysrtCaGgszBM
7svVMcUNG9bXgxbf3GipluN9CfrcBNYUAH7jaO2USv7AI8HIVr+P+oix35FkWXuP
Wc44e2zaPbtHXiZD3ZpEFa+rldvGWKqniAeT6wHK9WAfqemwiDGRuCdJt8q+lBOr
tzxcq6Z4zA6cgV8C2HeFnUuKZWjfyeLholMNiqu+SfSA4opJN/Y7MxXo9Yoj/D2Q
yfV1F6vMgfzFChtRPdq3aNGHBfHkl9buNn5srhvaSjiMl0kCN1olXBHUc2AA6EsY
Uk5rdDBMTdzdN1Ty1enw6rmjraY9gJdQguSF8ltwQBGDLcigfMMSt7Gss2hYNDDk
ZTa1M+hOnD7/OKsEnJCkRetg64AKKc9GyPnH2KKXfxKWYi6LBoXVcNR2l9tGXOcB
h0q5N9HtvMGU9JQxMddLdkp6GOo/jXtWKJ4lZ7TxYmL/cRpSWy1/HXy6uJ8o2rab
LkaooIKmFYn+V2kKXRUEUB/ytqHpV2ptWzrpMUGUw8U9z9X+fbPuVxYREnnivCoF
TZ/vepzsKQvY3Xyfc3R8hrDWhwZgCm28PoglByc19pEq6uX3wfLO6nRcGO26q964
np8EvCLTTQ4gPOLpxyrkIRp2xDuzhyObb2xisPi/T/tLHMA6gS9a5IBDA3svp7Fo
0xhC+qKnFOkzO65It2LBZVpt7B+ocMWvH0V01BEIVq1012arW7iq7UPgCZQPdmdG
YK6ntEdH3OouGow+AahUosaItL0z7Nm9MPqPAAz2PI3S9nZA2sGaCiAQQMbWXokJ
G/vz4wEuOSfQzDnVpXbRQhE9E37hl2moASFYa8PXBx4fv6HRUSSVtCoRNnAWrXyI
EkIpIEwy62qXVyNSEy9N1Qo8pkfEk+MO+CfgbwgV6x2nwuUdK91lGoqBDQ2C8QlG
o+D7KtUTi84GkWwMFxlJa8aGVtfqa/kvblNt9Plt5/rtY85DKvW6eUErZaWlzVRq
07zOnms8rS+e30D4sL7TA+tM4yfr7/QEOvu9Hfi7+3yPDN2NMVTDs7oJDAhjRIKh
fgYL+nVb2By45ro1JeMvnIGqSwO39Eq3dLiiY3iMPZhuxvWZsCYUKEojwd5pNNnr
d9nksa5Iiaz9ZgBTIFt9FrkQlFOcXtSWuyikNUvurleJ35X/SY0hdGjucAvH9hX/
ADZSmLSrnpdb7+4z0nMo/9l9SiprjBc8QQSsAfNoaTRzdhGJYliijwrgDkjEPe9O
P4tPjgCRD9+ZEVTV01Ri7Td0nsD3gdXk1aFdcrapLVR7EOutewJV/ifwyz7YaZvR
iStZw31SFs7EBeW0IGnDKwRBTwjHWlDerST3pyEMCn6/pA82Rt7mzEPoWiXF43Ne
/kbGkHW75juP+JFrQnk2uvkvglo0ZqhQ1PFKOY3YRWJXiHnMaMXDJhvcTDQcJwrA
bkziJURrF6X5EXh1jFuAY/0XiII2h/U7zepyTY8xmSneRlxtZMre8AwJ3DNRUCdO
lrfBISg+qOjchnwp3zs+7EDAxv/eaixlXO3iXAbM2mKUnZn+9V+F/PM9o7hV2SoJ
CjCfFZmRHLMuH+Dbnk48DgCVDxmHeBTdZ8DS1NmlZjerTbBY1cNM1RLIX2oDFw5m
8Qf0GWrp2ED2G8zDXBF8bFZ+j7dNVMsRuCZoSWtjP4d4VO9k/qvzB3B7N9/M+V+x
jIh+25s8HKLIkTjiw1fmhux0iRZ9IxTlc5WUsS8lwmG6/QBIWJ/bE/MQZwytTX1Z
nVtBxJ/aVRo2I5yscc5uI34Pz0LwNtx2vndRMujOtCzirLzZkTyZpUtq8iSLRNWh
ilfJFwmQHuXhMa0OTgw5sYBld88eWMvDFdgrk4Hr/eQmDaBiiZml+9VICEWRHjcW
Hw6Od+Wv+USYSnQRd+lzlBtINmF+LgOqVipvKUIYjZE0GNp1dGtO1CxGdC577gv6
8wz3tS8LrJIuKu2/ngsWEHyRRok3rd9OYqsAzTkKT9SMxvknYSWAVDNdkT91YeoU
6teYWVmDhdAXL1nCSaVPyTOWIGnLC6FbuQR65onGWLEmi4leBwCQaND+TBFhWSy8
Gh3JzXFZnlJApL1X7v7nxclq8nP94SzzcvURMXbfPtGBrdz5IUVaMwvjNflDxInf
FOinalb37HPFldsX3vSaBU4UEb4IF6XS9hzWUkit5kWbSiiDN27sYk9JMjHOLO7X
mKMc5kUAekzld6Fzjkmw2211ImQt6oLMGoiIgVsZ33eCVdbyexuokEbm5Umal4ew
d254WGOo7qZTSPvf7CW8Y6lgYVSlTy9TClwbA5SSaR0JE8wbtWqKfKzAz2EqFFpW
CwkSXSPvhk3hpYQw1X8jMoMOlfEESQjVsk386yHEacaYGOkVL+GnJFZxkMyEY3ZU
ifqE5J/FEH8S3DgQFBtk9dKpkWIh71jhL+knOWSpQvUFkj7ZhSEX4GOwanqxJGRs
nS6zOlbhMGpztrFhIIjzJRYlviorIi4XtlSpURG8kuVC1Kgb25P8mCcGCocxh3mZ
JoHlsR6bE64/LOuFWWau6J0tQKJoQYQ1Qh3OMKXxA/OjMI1FRFkgTjiTb7+uiRR3
YvixlIoVQeHJsvmuJvkENgyemvF/RFG00IwHjx09pGB3coS3JLfxHlcwTRDutQs/
rd9LgXbAcfnyjvMpLMowQIiDac8fWtakWUSgGk4jtbGie27z1LH566J0i89PY66/
I2fflnFPXwJcAY9HuVLRGST0ekVN1MOT2M9Pu83Tb7SZPU7v2/UX/x1GF8CNNje6
y73y6vxR6uVAtkXRAVM4226yD/z7l/ejc+/57IQUAVYzeNVNulYj7fE9A9W3GDcL
IB8Gs7vMSvY40vP0O2aHtEptDlVq142DtfIxvoYXykOA3DTcNd2yl5W68C/kD//P
8EvBD57Ia4MUhB6Qye1On3kKSP+A2ilxqFcaUiEyHpu+RGC3HMiEBeaFqU6XARTW
otlB2SqKK7wH7PHTrOwDQwSwXhMTcR1LSMrH8+o+7s4YRJJ78HZNwzqHx3gKU7+Q
2IFOY39kNzeELPvbJm0Rtn9qpCVU2Y7M5eefzPdG0QRDVm4kWQNX37R4lOE3BLvq
zJeSLEw1m6Quw3KcD8j5s5JfGWxSIrg7SowkhMym8HylMGphc/3feAW5DO4FTWnP
ZxTm9g2UrhIQq/xu5IdbEROjQeN6Mdtqyg/HpKB2IpaSGAsKXOYBCMyQosFl8yme
P1WESPnsHKLG2pqoyg9fH/btmbWkIXbTwqFAH/t+rPi3eDn/0IjpqWIPojHavDi/
nSrd3gvMSy844oYB2Le85wQwsSbZhwYXCBM3zrXNM+A4zpDubFD2S9bszJEkIupA
LJDomzDq19H0omvP0JtV9lgqk3k/yPNZWKIcyk2J5XW1RCCyVsasy/zRBZz8pv7x
5MQY+2KUEUk+u6S39EN6LwCIDzA+EAYnDtRDuFg8vozfRVboWyf5Rk9dr633UqBG
Hj2aRm710zh9WuagQFlR4WCecOSCA8C54/WpODv8Jpue39xDPNZgJaoNnjkgfmhp
YurzuuoCqNlg3ZV5TFPzWUdKrQTLphiGVQNnhN5HA3dbUhJqDAzNU8MY05fey3hf
Qe0vO8FezTAiiYyZkG1GPaLIQ874bAMzNF+nHmLwDF+NSMwsLJxudwiplI44durU
epq6AJ7GRkEL+V4fCOQSfFQP7LLOIJxOYdyD0KhLWZeWLgHFG1GlQaLBL8PpyGhf
BtTSmtbPqPjR7cbhkJjvltyXRCG/AfOllqBeIiJs1pkmvITXwEsMtB4zAFvlV17J
QPjuCo0MXV7Pa9LXXAAUNbeCaDWK7VMxpQT9Z1/NclyWlhTjAaILYoQlI8LFqsgg
Q4XNLPzriJMYjTn/w1wfnh0B14GvB3m424xZFKArRfINVtW0Qz04/V0fu2+d4/oW
van7zR92QmMukENriTrqwOA++f9VPPgerhJoZdIGr2MGesqH/RkAIoE6oc4RWFKT
dS0mPau4gCk0LBS/bWys4JcYRDAc9xNgfkW+vpoQYQsij3IIxt/YoJr7uT3ngr6j
IipgVA2Y6pLOtn7m2JOXHCgMWCbwSSsgPsP6iqyAuh4s/McM/L8x96+ElUkyVUVf
LXLfHW0tfZ9+Ve0ZRDa/VJbT/jI9AJgP4eghXLdQS3l0IyIVn1bF1lK4HIrEVi0K
KOXr2H0T4e1GgSnvMa85G0xmPazo289BvnsibrtjRxuY0eAQ7PHvfAJcZKNygB12
taksKThncxHthLMQmGAHk/Rxj6KCVgZUvxQ7BvJO7rNGHthe0WUDAUW6rIVFV7S4
GDesGUmfsYHWDAflcedClu7lzjVLFPrJmEGQnnc6xkV4fcMCLdStVb37KoLwsP6R
c71qQBlFt/Jgq2HZ6UBWGEyhQFCpaVX8r8MZDTryB8i75yz4Hu6g89Q0LrfHBZ7J
5fY16uwcZQGz2vFN93vH+re6DsZcp76ONABbVAzKPSRZcf+gOZb9e7lqUUyq1t4C
vgiNjPph0uMMIO59fC+KCIgopfelhjriPfGACZW6kk/SBdayEf5jBzgHBBbX0ny9
SuePNKKERnVsWVkX9QL/9olfZRJ4JWTwlXxjFyGF1akm7hjSrK8DkKDW18kntHF9
IktQclWklY6UHZO2qNFZuF/979/f6m+VIP14ARNvgrWIstoZ6AJuxhSSeosILakt
72Yz/wFXSmxkiwrpejZ1pRi55IJ3UbzWiaiR9GNnTRLuNHYBqShvKUxccui6aFGM
QbM/Ox6ec6JitHTMydzm2PVWCpjLdRMoNfBN39aouARTdCCz5qe97a7NjRoOVPaa
stX2laZBJC5SY/iRmrbv7KauSrdtwVYuuuxeMLEHkHcSTomGw0ZYnY0KZ0UFm4xr
w0P3didffvlM9AItl3z8awrLA5/NJNSgWpOSh6MRTYvx2eshsppusgdLLglwSx7O
/adTdkxDh/MMMysmF03FMvM9DlackkQFOMhO9bLp6deEE7C3BZEc4u439RN6LQ69
gvb39ynQt3haCGtxbkHgPgj5OCMTxTzhcB8GjkAoYgLZgTA8b7dbTvJYOyYbtWvO
rwLXkciZXnh2AseZ11/54/LSFNFtrkdm0LKY2bAROyHWzAyC8lwmDsotQkOgkbl3
WJEFCm2A0uTSOHRgf7bzmRQo9zLtI0o04ru3GhPbQ5sR7ijMlcShC9Y6XDechqYX
GuuEFz2IbXGMCk70Oy7FvG8QpLyjb5wgqM064d2CH+yAYiTRzx11XwkWn5RnU10n
0kCAGLLCDa+h3VR/HQmwCD1FpEETREkATXk3hiK+LsvPkFkglczVN125yPyLX3Rg
pB5VSEOJrRUBYw7Qs7iRaent9z+lM9bQDcldyur3UI1wCGcPpQyOSRB8av1sv8Nk
zRJcSAFkLBrsyfJ+QCeKHI7rkdX1Ei/3oIcEce/isYsTXuFCcdgBBpLAs0E/Is54
VzI0cOaFngY+1TVKdee5mv3YpZv1ls+PYW5v2n/nDVWlBTFDscTNW3CfzycmSoMI
7xwKnzQWABi12kfMHkqrGw4r6Kjsx0pT/e1kMOPbrybRtsaF0jm+CL7gKFcZwSxC
pjegyHm+A1EBNLXZpYqB/6r7VSL/Wj13qlEgMcOeADKLagAH2YVj+00JRtvIsfdR
AtuurxId3LutVQDcw6t2uQFsWtME+SZ0AMa0Fwl0YdpC6U6SgV31NG+mOCtJBAtS
rSPPc2kUdiRia2/mtSzh3Vm2YOy3fQp8HK/QbFCKXIcbvE55cjGtEQqcPr1w5pGW
rnncuINZ8ZLUik/Y4kOYndQ97hITV3RiTQ8a1fdAZERy2l5+hQb/Ktjy4NWzFOn8
ovSRuN7F3CLX5OlCxjZW/JErQtwwwg0pn7NYd1HbMpCF4+0DadG/ws1F9w0y1Pny
+N1ckLzOWS3VBzTiU6Bn6J2rHSmiqjpkH4KBdCAG8sPW87pwnemlmrR4xRrZtfS0
k6R4jv71CdydzaUnJqwJdP6D6acudZlWgersaYyIpjW8og21cTRBjyInrIaode3c
rz7pQyZBMTZW9EiC28FT+YDHk1wpy/Kvof7MyqsmJaynddrDbMgcILgRM4rPpenK
v8NCJTikxN6b3M957f5DmTyNsFbPhjGq10ppjIr40SYj3SQddgbJqONIeGiWUm1K
TQ1ZseqsOx2lGajb6QFnxvhc8ziBX2a4YW56yn1uqhbnvx9U04LnG4KSHCcUZTEb
EEaWQBGUeMLUmKROjGGRchKaUthap/PHWyCcBFve9iziYXf2XzdCdGYA9jOqdl8O
ElZ2Woo5kL5tnOooaYZ6plNA3FQPUh4JcBCEXTDWQqXpFGQXFp5uBENO3xd0nZbb
VNa0+RIfm70ixpy77siiKx40z/B46BASo0KlQUvffq5BN/e8Z/pV0PwAf/6ol351
kP1EgGv6/XwTTVZFceiSQhXFYbOZ+AHGwS2XNtOSBI/Gu57KpFGvvzU0cBhQaPSL
kQI86fyCJ8UIDEQBj1YjnbPsbPbYv7tbtahpbgV3nLRvu+MCHgTPjA5AmKPCZ1bc
cNArecWMYYvEVrKDGamVgfyTjpCFpPzT2zgAxtj6lFsHidSLmpcQjPTq3hh4mQGf
QNolN+ofBh8n4rCM8hfGbwuXCjrwou++3IBuCmK4l3qDJf6V4YJPyJSHRO43uB34
NwEhae7z9e3Mu/NTMPdHJ0oCsXzKRb/Ak8e3PKQ38PUGCXsIshairzPbxJ24zOdv
TAVv20YoJiQYNviJHwHkt8vbJ38gu4m3KPiCis3NwGnLarTpkFZLLe+gRtW8hgXT
Fa4n2QtsPjxtItXeTl87X02ihQRGkJOMkdfQaVlaIXJ0vD+ME4GAvFg/tID1ITEC
CigEKJsIjZta4RFdCvQ5VK5QUyZ1+DippK93PdPCme91ho2hu5AsKbpXEf+a2ohm
cPepfVHU9CMtjyoGE7bxnS2IIN7Iw+2IM7uXkofIkgVynj4ekNkK151e77+6DYHQ
N9uG9/0Ef5g+8i+X/g2mjjrW3vuUZjR3KDGUQpdBihvr8Der4w1SfAiipKzrGkFn
lWC0QbeuJp7LmJa7ydIdE6jJ/rbG4QkWZ6s2vxw01rSvJ+275r9v21ucuzSFUh/2
OkMi1VBZJiKUHaGtAOdKr57jhcBKI5v+Gf9LlAQEEfebvVoDZbCIT/JJiqtVYwC/
XyqGgtFQnKdoDr2colZ7oSzGDam+2eSB2uXl6yCxf34W1CjUjh4Kpg0X+8XICUZJ
qog5RKLw5CkuVqRpd2QgYKpjUhjzk0LlN7xpE2Cd7afgEUMR2BFpqgy0+vIafKpB
1FFGtWqtjwyxzkNh5yKToozmHrJHYfVOMTgti9BXXvENy05utCJjD52GKezNfQPI
PUgUML8agkM0L7WsH/LjqgBffoLh6Xup1z6LrD9t/DEa6Q0QHKK5US8VssJVb3mm
NjcQRgHlqaRQsAd8wr3qgmWMKa9FZzGZbrOayY6lNbKJWFT4POzGN8kgjc9Mwbvv
mov2WsfhQ1uEgLgJmqC0OA8PASCOX4LUJ11U5lQOqsB5q73yutXeN9XuhUWuGYAV
aNVTLbuYxcGKKa9G4BYG4uS8gs7LUdkGMEfPf8kKLHXvT82ydtT7vu61Wa0U2Uhr
Oie/bTk6JVJFCQ4c8oI9KhkC7f3GMaodPFeZlKOYtHhRw1Kj0FZnXWeiLJt44GeR
Ix0lSAnM1oHOYNuc+OClQdxD7KHv+Py/dCHChKQkEfjQOhLBFJWpT1yWaGk/xjt+
npuS41+TNXS+NgQspM5a4Ev54olpTqdyx7PapHGL6+zkV5m4IChGrAlbqP21xnuU
MFry7UD6EJXpNq+SmjlWzINPQt+OsVLqjNvQIf/JJKxvKHCq0acGuGY7ClEk5AWq
T8dTMM5/dUc+a2po3D62V6hk22UtW0+ec+MjtK7W3yeECJAMeBj1MYgbF6sbw2Rd
tpjASeVB4OoShuIzwy/mAC1+JJMGPpQADVqkF/PrtxuUT+bB60pmlr9ctR23WiJl
kE3tek1BiivUcKFFWTrPbXxFAeOi3ZR1e3eIz2AVKXQWruGCva1Ol+sDhUGG2Bh/
4a49gYoSzBA51BZJ3rUVWtUxg3Myku5mxZlDZq6htvcGrLPZN+i793Vj6hnaizLA
QPeO+vk3PyI19cS9fw+xu1WSU5e6UugD4bOdHGTLcjxctbze+Sekzy+LWPNs2TRe
FgD1abr3QDwWrJjKSMvrb4MZjWHEQDMLgQKiHvIYK4Ipm/L9l2myKwBvbw8J85EO
DX4HGFJGBjCC215ZR5mipil+xclsyPxBFGzwsWPEQzotT9X78prpYC9wmegZddgO
D9xQICz+VkCAJGKAOHgWIsi99s8vospohbfiJ7UNpOaWa16fXq1Wo9TBu7yWJCio
cNz1J7h4P+l0WjhSIAhTKx1DZM3QMy0Uhkcy3W0DM+AQmbj5GPMsiazh+qpdMxyg
psyypXeV4gh49qAGpowMcez6ctyZQTNQxU3zatTZM/A+RKLxKZ/u0jjKP/CHLePU
R8eC0llBpFvznf4eCSPvYXXIBiWVgfXF1ci9H7EHi96D9eMVY9b+VzI4bZfCyr8P
trhgKMy0Xpu1M2RdxA9r28LQgiPbBolenammuSAT7QV4Xssj/Ys0bVSyQQviiM6b
mLViEzE7guD8Fm/DbsZahUlBW/IulTcLUZ4KBxE+e+AmalrA49gYuj/RtGw1tdC5
MxCm68Y1erotOcjHb7dAFllHbdNCMeQAghI9N9Lh6JYoFV+9hjv5m/lLAvRmgi1z
uUvVO+4rW2HCsGmzpdesCnTjDWfOTyFkaMU8WCCB1U7vsAkzQ0fEunqQRtCgDKrG
fly8XwlYxFcz5meXGBRN6r2o8IwGW5RC+XIGOxjCEnYj33gs+S8xiBEAMshGbPMg
TUT7Pw984omGt54v3LhAvdPJP4BK7itdiOZlvHUpexWTZSG33UhdSxsmGwWrI6I1
Xzn/EXx1ZwU3QSPwIKKKOXcSsequpzpXAHrC2Dkboqx7vN7KpTdOqrhQwlcE4KXv
g9OBezx3mKO2coAKQybxBQ2waj1ETOkINj5Z8mUfgrYUAHek1j2diaktwxjCsgm3
keG4/lzCj0zOpg9fp5PMQPqnj0LkT5mIHmxxPi4Dxv0CMUbntFcejimNIFlsidyu
WMcNFcNDKAm057EVI3NFQOlghFY3K398m+dg54cyacW1U1Z2hIU3xo8bmmcKTI3D
ii+MPwe8Y7553LFf+THgDrEsUj/YJUbrCdEbweiTgvxFAMiLZw+ark6rllvLhlyU
iwkoPOIn/+HL2WqkAfDumvwAqFkqE3TiXvo/pTtIsEX0FmXhhDf7mNjw1bt3YQL5
qI2QgrBZTeebOwu85pkYkwqqrGZuFC+6eBM3Yywe4mwEAe+eZZcMdqyw3FihkTAf
YFJBQ90wQUs4jpk8mQa7OXvcT2WOLdbOYKdoibTCq+njEmnuNoEX61v7I/jvUFzI
h65dJ62hxMm4zzL7zfTLeEBclrcYRas+Ahno5+oid4x3VhJh0kLMwaOlmIaC3+DG
mmk2wikutyVVkS8gECtuSaZ2EoV9JzYhzIKAadpWAYQ37zEC7fXcg9EvtQ9bx5iz
UKKigZfMLPQtl3LTRy9+OKuweCOoScKjzpK1rFTayWtMkxRs/J3pwMiJ62qvD9on
xh0NkPZNzIwHdUzoJVj3Aeci+chbyBHobXYFagoI6MzoDr5Icf06ZN0J4eR679h9
n0U5njDtLszgHlDiiwdI+WD/Wykdy1h2zu4kPXKfo24mVmK4QpdleZSAQDlpaqHc
WfrbT4gaYWS+/1WgYiI02oeIfPeNlWf7hEjl6FnEN3Pg3vCZSvgQPMkaERPCG31d
MOADThYUq2bO8e+TLxakAsRX9zGwgR/qe/gB4HdoXpM3MxpXANbed6llw+uEzi0r
+ni66pgeAxpQkEYLSjrAE9oPXHhB2f2PDmUzkP19hjjBNa72omJP3WiRRZ3jvvqN
JbI/mi1v8CUIi8o5l7TshHkXhgQtLjZEileq7vAsmxJ1BVOx9jUq6WdXgkVHYFb3
B6l7zC4LJMcys5sidT/XnJ5PVctdPVjB1Hd3V300IKTJl/C066UbGMk5xzuQU5ml
EPo53GD+ajyIMpFesbu32flFailHdfDGsLUgSojGA/1HxZMCELCr7qZmS49PuYMm
Pc3pTbZVZIOl78XeS1IzqF+zTQYGV1d5aDZNPZ/RwsRjcXLsyY1uBzt/G5bj09tG
4L/MBVWsZW9V2nDrOdxukOwuqFEwGef0aNF5nItKVJae7XUqwDEr24kw8+9EWAx2
63/I/M72ZXQbtYZktHP7YwHdT0oEtbdFnnVi/tLKD2/Ty0XzgRcvhAgBXV4Zi+R2
LAEDd0PWKK2ato56zSkddVqMRRwWDnfDproygOdKluuPGvpPaHROCZ7gZcpv4lSB
kuO/at4j45XvwA9/5T1HqEzTMuImJPUk9QeemNu7qPzZt7meYvM/G1haFvXOW/X0
3Kg+CGsRF0xtmInc6n4ZERg9UCaOp1SKOxNU05oLDKhMhr3Ke0/YNfFTw34KZ1bf
Vj8JlYr0Xrz7nL3xWQkBzkeltl/dqyVOWsas6jeb9PKLWRbLN3qKd3hbRHkm/fRR
hWPocu6P8wltclx3tiWMQyNhlm/7ZVDW/tKhAFJNw/G4f9uQo0q5aeSh08gpbaqc
6ox88As7juPq9rDjLsCavA7wDIjuzQnQQChMlfYnJBXxSwGas873JS/RTF1e9/9T
NyrZM64N7aZDHhbMlvPVoOQu6M8jGfiZF4gz+XA/xZjqsegJIs/436lzgcm5pLom
E2mlgPjAR469pWP0RzFLB/szvXa1F6mNXcUmldtXf1eMw7dDJi2V3VAkPd5ZfStE
Mx8jfKX6s9XfpJhj3MJtKiNmXmLnO39K2+GCL4IrZGR9wTB1pm/kebN8DcTgymxB
bicKstZ+F41na9b/JjE+k3rqTgkQq64CKRiSNZTcQG1b9JX7MarfdLt8WGjunSIt
6UevHTwXoReOb9iGrRvvZycnjnJ1b7JR1H/OwX++dRqt+rH6Q+FuAddJbxEemiyz
TDX2mOyHdeRyAnbztqUVLxv8sIUfch3Pw+770DP+E30/ksYY/I++2rFV8Ljs3CMi
VXAZScnM1vMYf6G+jfDb19T/TkHLGfaHRbVeF2X8uwCwM5tT04N3W6++ja6We7gE
IMmvgjum9wOQ54PCswUuXWGs8/0dpDc39VI+/NpNsW5/qeNu4r9McLK2LQKClOKl
8SmUUp3W8sPxhBuycasuhnyyoUbUI5xyBRiNdSq9qZwDC6ssloSRbLHfYMYbxzkn
UOFDq5wRdwCuhEasMPb6n1knwaJa12kRgH7nrfWu6nyQ1TZhOYMUEvgvY4VZ8C42
/fnbhylp+W6Ys6lXNd6+dwErXkiOVP9CQl9cEK0YYZO4I0RKw2ga3VIUbQKLFWXf
WFBQk3IFAuIsWk+kCCVrU/M1w17kjlGUBfTCvLqxIUY/75hTTamBa/19PxgyvDkB
gZ2jIGkO47DKh226qGTB94Pw7PLVelAZy5ydcsO+smme80gcsyKgkWGeV7X2ljMO
kkmLOzXgV1cJwl0tM2254vgarkHFrCqjaIIvG1GQxGNLxgW04LhbijzNTt1tey8O
iO2zU35vS8j/DgbP4afnYCqq2cTUZ6ELgRwFZbc24v49io00muZzdhbkUYZ74HMl
btf6VfTUE7pIolys0APwwNjxEMctM+kF6IkYHPUwftTYoC1AqMrBHWLt+8w7mDYI
QeG9lwlQDsi2JW1foDnEsaYLGQpNaUHpTkLAr44/vKt4N2zGkrF1I7DdfuWcbw3w
u0I1huiEC0r+EaQTfKaNkG+4Hu1/zxpJ8QKCGhxKqZLLaLIt3NtKnX6qg01gWukG
Rh7SKCs4NOh6bf/BpbTQRWJ4DVdbISi8Soxr9BYArjh4Qi1VuXWf7KKY2J0p3p/s
k0PWVPHydiIKXKS5O3MuH4iWT9idSNbDQFB7qyZhCSm793+DvZ300SknKIXns1Qy
rz+ziiYBwGv+RDn4NpgxaSRyC3hafZ3PtIYJeDQFtU2Cm4rnhWvftYtm0yoDtjUh
d/tLP/C9XSnhgkylEMRXu2jcIbg7fm8zSHeWXfHRqaTFKnEiwdPptydVwORfbFDc
QyhIVFGbugQl/aMUL4hy77AxqYF1KFTabrKklSz2d1O1X+xdan3860PDXmG73hee
dYmXZX0V9Ythkw93PwXcIzwTPR14UqX/VdCXeLY1TVxaJm79bWrZbTWbiZVMtRv2
6Xf/82FNFY4djzPiwTzY3xIXsVN7qvGJwTRPttiKGo1qdx27OsMcWUqkk7AStT2Y
fJbqN08a9rknkC5RA5bPs+r/0z6zYps/jjr4I73zHWkHLOLyciwuBooOoM8HYbRf
WKk6Reb0Be/xoqWFR4nBGllHTtEJMCyPF1LmszGhd2GblBU/RF2JJczCEwj0wCUa
peGGtkrV1EiDYzlD79Sei1EhLLxbHmQ883nwqGkwA7BtPmP87iG7IXt8yNR9y4ve
/vJpwH49ZlzbmN09wwkzLq8vO4WDPPVk9+yKikggPUv4OVb4U52QXGNJqMAKyym+
CiRn9RqKejoPVMldEKXhe+PRi1jqqAok96vFsH5SvdeZgy98czjub7UY0zm++oyr
Un3ZeLWobo7h8OzYB06WbpP7wuopX5cwQvkD5BHRTRz7aR2yiOtPNV0onSC4Nz3Z
rp7Wb+N0zM9NvPlF/xqgj+FZxy8bXyTnl7oqZznzbwCBpWXQEYrglY5AMUIFgLrM
h7JCax0dzBeVxtFtFhuEBLFQK/+TDnrRTF9x0q9FYtAqE+Qn2N7r8YuiWl4JEZ4t
Ml5SjoZsoDE7KMu6jLIUyjUAcWyLPDM9hKBgqvSAediy6Xhkx0cXIyedYJqIF4zY
zH6uRTLrq6BNOSSx5kmdAp4ZwqZzPIglk+P2LDPVIyq5fSsqTXq4/BEZcRNcnLvn
Fse823AnR0LRHr2f6Nlu+R6ajb40mtFXtP6Jc90cHvOCVTf7nI0MiFiyQuUF6upD
zvA8O4ar0BpP4IRJ+U6QRksz++RaJmHwmTsE+qcX/ONKwoPv+ER8BljIhMr5ANm2
vZfN/8u5zCfXqtaMoaPu7E47SV6iQocr9OUWykLHX5agqLqB/u1NVA+GRFqVcKdG
ENlQrg5H7Vjkth8hf5gdXGw519QLV7w59OS9/k9TQzh11oikffuUjnC5iOiqBG9A
Ssg0Unb91iEnpKXVnlZpaONWjyGC8D1L6D4tmZuosa3HYlJWyxDTilhSimPpkKEv
+PO34KU9EtYSDKwPDyvttft2iE/9zXRPSrww4YFNkCbvMOHIJJj4fqZub5yhE4Fw
ZEKdzdFjjyFM7WbA4pTCh77C+h5H9UIKHlPPQqCVI2RXyFRa7W1se9chLeS0bQPE
BGPnez88thRZH8bUkYZZfppkuk7fhH64l45JxPx7rA3bZoGxrshffRBkQNcBrkJF
8C6RSDVNTAqDYXqzWjkLMa/g8akrmjhWC9OCs9tN/0ME1UA55XCkVn5x9WSOOvjq
rrFlF5MkRaXI9YPU/fFB6rFC0J+Yy7Lu9j5+Xr+OGyNF4b7Imr53a/XECUxmIoUV
wzqkEJiA/nXXthHBQSFNvnDeRWprSo0uVc9tv6abXRsaDV7STqxkwFLppO/r8whW
WcSSPqFBhKwBVfMoppjXP6ZACv3hxTynBdpc/NdHqwZS0P7AhM0jDa2YS0ZqN4z0
Au8pSHkZcqT3Zc5JI5ouv1CPpupzW0OitYtZ0Ail/UwM2Vo8YcWgx6asUEvXAelp
hzR0wbKJozNqMvRbPZNjW/pHwjJzX9plJz4//XSjsfqJ/WdTZXor2KrphZZLfpBE
T5KYA96hp5BWhIhJiO5GClcaaeWR3sDAJZMsX69lYqcEHbz9dzA93NJoG6buVNIB
ui7mhwRsmDpDZZ04aMg4slp+kJbpflKsEEpNJ5Nut1ixziZ4d6+0oF3RIDrH9art
5rErSm6NndT12W9XTVtU9vM3zAixQTBXdpg7JREJj+7gs3XnH4u0sf5lLiAEmDpQ
BNY7tdVQaNhRS1whxAu4ek2emDGtHW5IW265DVjfMNpSrNeknXRumghC+3vUWy0Z
RjXCqeRxjkHp4h5CIZmhcjjfhuXrlTh3muz2sj+rc4jtUh/kuORi8+P+gXRMUIfy
SO51Hhi5r22gnrAAVYhbXD8mjKviFgzqmZONhsdyNckXhExwiuBoZ6B4swOCbrvo
Hny7ptoB/AqhkhaP7k86pBnUt+FmxUKxDu6HKPGSFSVfxmjk5pS1GLwDlmqgJMXn
i4+y+KtAYcDs40FenXY/YawuofpR+o1YGGDHCxjydsntEixJJ3WtUVGP7PNLLFy1
K+qP6wQCQJyYpdBOgYXSB7Ue6zjQigQ4co8o/lF7nWPsset/9uccNSX5P2Bz5lKt
m6h/oPxA/Mx9QdCEuTq3FPcb3kcIDY594KM3J5cDT8wYDIZxCA9xXGJwFJNa5HIW
nVSWszQNiTW2bAUN9abSi2FrsEGL18/+noBbCNG5NzpByBnX35F9+DFw+banfLhg
PFQiKg4FInoTD9vNGU84JpAynONChcNgr2UWUJf0I/gxtKZi40IVBmVuE613buJ3
iENpAPmcd66rjHhtqpe9UHexlxNQcumOhEH+qgvAXm0D59tUZFKE/yusYzpShGoX
6pFe0W5Eritp9YObFEeRcoC7XNeSQtUlhy0dA8ZZi51dink63CJBx6ru1g6Dlu2B
+Fnd6BVZLreUl4KCyPEZipOTtZ9q1t95EzLr8aT4HGQbfQxRzn24BGhiwugWLEwc
N3ciZ0fz4YtVvIJ3tW0Lew3FdwAtwnk9GABxGH9DVPo6yVanJvejXpkONpZqAr4Z
KyjJGX2enn7ItZypOQzK2AuHbUQy1KtQcTe1cGUYFCjdfTfFS1ssBMwFdSpgO3iF
4pOVkYo56k7RVZ2aoN0+ciVzDDSnd796lDgosRhN/9AXDaUpBLzGYCRlbFDz/Rd+
ZuHyJNroTiqDql9Z2CHeiuPELK0fk6iTnw6LGfRTCCXUwO9KWbR22sXC0PuWQDZD
jgJktWgqeqfQPOvRzMje2LA7OG+nUtxoi3HfiIfKirhpw1SbuYhQn/2Jt6sV7QO7
Q7H4BONnErVdP51KdiXrVDWPNVU75H5NWZq71JbMcP4BpJDoY5n1m7RrP3vJLxtV
8r4O4HjArMiHItXcm5GFKOsihKIu40oTP9qLOV1y5jK8n+nVrk+yPRPW6nAI7Cj4
w32d+BcpiVokDbcF8TzAo5M37u+x5cqUtqX2tPMd0HBlqnF0iBQtFl6AYQ7VfIVj
NBeYgMdu++iHI4sTyii4Go4bG+HTOooOnVw5q4Zd8jfF4nfQtdIjtg6XIYt+KJb0
woEdsd0tMLDxyfwd6kHTdcaltWC4cwv+0oaZ5HnWJcvM3sUMZQWUDAVZSYdMjVdb
gPS9OTofwaVl7blSw0plGH25Ua0zjSoDw4wY5tClrmsburUR7ezYgPYkrLykUWHO
ndlF5oQdQu/hdF1v5cut0kSjwkd0IbP+H0oPtjfnO86TWYAEgZwGgIEIGB6BiDGi
GsPzcxfRXpEFwn34DlOv1gqBVRowind8sKTqsGXD9R7vpMg0/Hv2fu9pKRrdJQOV
4tE23C9KT3rkARIUh+2bjFXqEctvbLjKgmz5VtHu5U1SXk2Y5GuISPNGBKKXlAB0
zLzCJOlSwPhT731Qw57wdzE+0iAfycbLZKcFqQ2IqSVduEBoAhyo1ZSzsE2b/Rpw
FYkilzfPNvxe17NZxCaq7JDQ/QtB8OXogA+3vp0hjw55J5/JaejjEwd6YrCEJutF
ym9ADkeUWRKEt1YvvVXFOmOc+SO3U2uWQ+wR94UX5DA8Nx79HJSv6LVJ1X4Tb3hQ
qmoTg56Y6bVLuFScO6e8OiWegCrmacTyPvGtxjVHR6iE33h2Q28G3O+iR6OE6cjC
aDNoxIRtP4UsZ34nbfy83eeutNuzdXclvaMp4v19pWaKGobB8Jhk85nuL0lh1lPc
ED0V9sBw6X+tHib3SswYCYQE1SB9FsRE3XArvUx6aB6qexp2zarjBSetjqYN0Sx+
t9uX865zBzYAjTl4u2P45zkkiBQtbPf+TgTj+V4ZsBjOLYTMyRoXaeXVeWcPfPBK
nkwvDxQj1OJUJfma7Nd7aVp0hrrdqueSdl9wf3e3kO+2+6c6SqDI1kckl/qbMm26
jY+ehvbzsTr9D5y00lf/zIOkjtyLM9B1eZMjSYkp8Dq6xORG3EejSkqmjN46M7gt
92CL4iXdhM5ApGN5xjxeHwrwtHiePdNYz4JmJWZKnkwGNVa9oeQGS8ypZ1GfsqiG
NXE36Ca1AaSFBk1ytglvSOXdW/S9exHolzGYW/DdzxndmfZOtNMWUvvHrlqwmwHR
v1Ir7jAmmLC+h+MO0gCAGkvAJVByJE1pK9zdJVP7CQpWpnZu+Y49PEcLGikGjlbs
4psAjv2mBlvbAhjiMEIXkg6a9/C2wvfFcoQz+04sv/Q7CO5YxnujO+lULWGS9Nip
M83QRn9yWrZV8I3mTFsDubGGo+MbkbSaMvJNopXl4+4LQwZGo/b0EOJeOIVFx4Dz
Rf4Q2judmOeSXj2eU1Yzlv51tRWeR5n39A8Bxh8Mc2zc95VmDBEcmCb+oXc3ZLxJ
FfwOlzKHOJ1O4GV2AOOqkjxmiCPAvF5pANNgZNSP2fIkKx0LQAUumK7+vnUb13qD
/0HMfXcMe4YeiM2GToTsm3+sIs43G9vu2Z2p+JFHxiQ4IpDI3RmIZrvVovzUD+lq
CaS9HJwZuL7K43e4vnfCNuAtKvJxHJWsMDfr8UyDAJWWEbDbo3+FWcJhLn1RLBuh
UkiyPPEQr5TGoFJ9epL/9gUMGJH7QiG2FxBqM27NFl5ZV76WfJeUpABvE+ZDdQSp
pw34thYdQB4w4kWQUV98iDZJAqwkWDbQxrovPTAWoXzaKx6c8mi3qYhitaJ4sJIb
b69dK6JrQCw/9MfRjgTaNs1xE8DH9fFVshaVSLCsMtyQldc0IBFlq5pVRhj1/WtS
S67TSr3PuzgrJ0foN2efM+VQ/wWJfOZiYJOv/kAKRjdlstkGhsS42Kmw4b25Xu1w
BNOUKWsSWgnIzbPjLX6PMZgwWApbPlVpuZ4PSFNrpc4U+Sjem5DzoA5iikEAivn6
tdWn/T4oDUTlB6cnrZpjZcIULjNg1RpIkNzSYh1K2/MGEWlYDqYcV4eUqdgSbLuu
Gv1iWYd8Oa/xwd55y4/o4Ir+jLtUP57ppRYY+VJPfwpOgQyUUXQDPpriTErbmOiT
sd6Yx0ZTgwiYgwcayoo+CcifBH+FbcCWhTBFeQbtQ9SMP5d+Rnid974LrA4l51LX
1qHO/QIe3ZyBe/Xnoos5ALcYSqXpY00P3/EIUdDvEDv709aXKuMIt0eG11TElYZk
f3aQqlm2pwzanpBWp+jrGPZFuu+EhFz8/UT8xkTwiU3tFL6vcQ3+Rmbi9fyFuj0m
FhoFUHCG4ewRVbY6t8BR89ywaPBj54wC62S7b/TLrB733vq/jgD3SE3e54FPcZb2
z7bvxuFeR/FbEZ9PoFeBiBmrDbd2K4yMAtP+XcvpS+rrJ592QwPkQGndOi29nsDF
vtEt1IQieFH4sy345f1a22jZ4KkHdenvyU7IDAb6+FNjMUQsc1Xeumb9Qp2ndZ+T
ar5oKo8vS3b6ubuWDgEiFu+ENS5OPTYsABtM7j1rCNdlkSqZLilK7dl/fCnFqAyE
qqMvbQfK81AjVPUMeB6KMlHVcFu3h0eO9yKFuKm4r55b3BmyUPV8h3fb+lRpPB4c
ZWwpQKS7M9nkKcrfkgB88g0mPGV/SPUxheSKKMaZqt/iYjiz7OOQzfvL6jcO/+04
wjYHGIWWugexcUuuLVXgdddI/uPXU6mKcLLxgahQx8+Lr7gDiMH15aQd5FQbz8YQ
14wNoH8bRHzYOkmMeYMLCQ88F2qf100FnzCcdKcKJBVl5okqFuyzDGRT7cztklTE
ncYn2E2QVQPM480cUm1bSFYDwokaduw7w4o7RerHaO58aKt5H/wPW8laFdnr3/Cz
2JyymehzLzF/rZmfPK0Fss/r5l8JAkyVRAyF0pZe1iF+AfYYL7hUmIc8fvVd0c+s
eopMq0mtKpICFh+xUaugUIvUbu3fmy75jb66OCCc58JvPRe9d3ZJjNuVCk19iY7a
Y1xB0VQAzvUlloox7wTxR9LKCwwW1hijL+F/mJQIcAmttpNZqRLHgj5yumQS8ll/
Z9QmrV9Ckr4xL4i/MkqiRsdJx9PM7bfXUjS6UHFvtwhrdVhFykoFKfnT90Vflq8q
VJhItJctYAYvny6e1qoFfJOR9dgpYSrNhtFFmrvWdQFk37DZeV1Q/DMe/sIr8Xvz
zfRqoer4hgBFf23aUNU3ndBH9wFmtkVm9ptV2nFz+1D3d2TJKjTPmVatCoGlqHbC
fAh5nnSvFGGhKMqAozZdslHWBDpr1r9eQ0MrAq/MLFbZxYSDb25wfK2+MhYYzB9w
A2fZSNlprmuwN9bgODYTD2S/JMcvOU7WppeAo+8/y7ARdLzAVp7XAwmzC10Qb1ER
Br7eQQg3EQ0S4kKlJETndTzvzpxoR3SEXgSJsBY7MEKF1kf6T5DF7sjEXaOzuEy1
UnkIvQpgUE82jB3TeF9cGmLJoxi9sUxYoBNFVS6e0f/PKKB6QbTC5g77fKO17gX1
WyDpbkCHggo5lbkCYv40eh6w9kJqt3vsl0Om/5ZIP9vCA0C4bkXjavPwwsEb5p2S
+jyhgDshSyL/xjyGidnBZuysNsNqNZ9LnuBKqo/BDW54d+668BXyPgE/bAQI+sYh
AAMgAZmT2LCrUknMv6qlyrA1gNvwECtNM98/yoSGaI8mClzf4tI15u+K0X5WG2CH
RMo9cubFuDZbSU3Eob6EGtIYDP9zMNIM078wdsxEmsoXdOCeEVu7YPl+DREVCYIX
w5sDcY5fjj6NkwmesyOscq0m6cq03QYOfbjPul35CzR6fXckqQDVIYvjayUaw1ei
Jfyel67SlofDnBwDflLvwdgWPE+e4iGHPpBvRuHV724DwRi57Sr3b1WSVpUU+fgZ
09rBHE8gUoxtly/NGQpUCy8iCzWdgopR1c8pgUjd8K4JCsAnOy2NV4asRIXWVGam
WyprLVkf92nyGDtdYY7p/61+t38Tfh/IugkqSGWdk3mai1X7BgNYA51dpzet25zE
Iq8/bPDZ60ttdVvJI+U+wbiMRJ2TfcnRf7XTQ+Q7I+ESp/bTE76V1kACVESJPjAY
38rmWsy7/x0nspdsRQc5si2WRQufYzaa7XZlJitPDyfhoZTycyFZt8TesJttZJwE
vVYrymhV1HzdswXk9BPpbn3ExMamcZrj5s77/hChcn70pjr/rTmS729naawUJfFt
xKN5kZzn7JV/tW9YlbEo46AKDC8o7PrDDboXFLd6WCIBBrFWKEHGVu9izyg2bSBw
LTHvBjqiRx7QM3ykukUzETRCbNSpoKjwmq89Dj0U7HnV/RPRVWw+3hhLjr+rGKxc
E/Akf5Rt679xX3XjXXYHQkvuJyedCNH1W3XVpqnK03UOPUBoZHccRZY6CNbOn3ij
ipC9DRDHeHR0AfNDmYGR2zjk/k/SQmLTFjIdcS/Lnsbmxx9tsGXvjNgF7AwBI9Xf
cxj0lQB8Rk93tLXDkppH/5PyOubaokrDKHrle8nPIE6le9RZFur9CV7jl85cGre4
T1xFNOAElHtK49JwWUJ4WEj+BKAbOKo8K799h1Z1TrwhKvQhX+QbVjdY+pQZUUVD
bJs3tcb0ar2iRWA6+Ci2iubquKZE0f+EyHu1SfJPxUpUbhE79G2mQJtSJfq3fjvb
cVUYdXU3cHKRClPcYJRSa2mJBoXOhcJK5np8Ri0Id13JUBLvUDLLROLxrFNzQZ4s
HmOnUGZ3RCPWbwYS72szvHrA/4NQwl1G8mzlgSY0Gjq+qLqHZUo7qeiHqgj7uZZs
E2y6QdMIKP8mohmId0ApbjbxMaCUa2bcgSRrkhN7YhVUR2VvtqeCX8pN+VMV7gdt
YpeOldoUMkG4ha+axzyQVrxEryjoqny0HnBCzJTdAvrB24w7STESucZm388Gic3t
2VdCLZRvRIESRRjBHylLYEHCHAlNCZss4TVb4XHjQ9IAjtT3yvrzRoqvjELYPa9K
5vgPJn3U60W6rhycfqYXKmQ0moltIqKbuO1uSPP+Y21zRxkPwm7OAYxOcL53mY8i
NKGdha17IAwHPXzQviEbr4hXNmiSbsHYhfftROZzr8c4sWCEFpo0IXL92Akejmd8
bLGdQd16EgStIZp4C0UUwMR+Xg41U5YgqYLZ9sbNktk7Cm5dpsy/Y3XSIsycEQUk
KCQQSxUM6w2/kB9RcHcy26qgjL9z54ee5goqiUJ/s8nakGXfi2qhnkoFcLMwqhaC
ucHDIxCXsUncDJIsx3+vVvcihZIXqN1A84kuumhTZF0XMEZ04Fqtv5mX4KdE2Vvb
2q4mJfF+guRnMMIX8bIHIHcrxk7khDyKmjqtC0Cughcfylmc2yStE+z9jpLg211w
Oy9Q6JdP3Hi5qbQ73ebE3zPtIX+3xaTqjnhR0cBIg2GwFDnniv/c7sBTuQWznkxa
pZdlMCZkqaQNRrJ9zfTOhXLAxAvzXRupFlC/tJj8p4RR8Fox2HzUhjxlZ3qpHUNO
/dvsn5L5y+slCZUToqj10NiDonIhFn5L/RAThPfLNoBpQpiUpO7nWRK3fEYIaYTH
BCau10PW9PG0z7Dw6t6l/ufSWWI6kcJ8HpA6++s25v9hQDjPCnlfvR1NuX4AuPnC
bDHIypxTy2dF3C3RhcYK9jHZiHxUqGvHvtfni+ptCSjQTotwrps511ryOa/QIvrb
QatwdoxEeTSyz40Y5vxrMuqClA8mGyGKr4A7SIlB3iHyRYBsoFphO/H36Nr4QGmv
pm7CsFFXEiJS1xX+1x1wwPp7hbDCc7pZnZWbYDQBzQw8LnktL52AGnpJdXuyyPwP
Jjm3oUjPAvS6QRSIA64N0z7ANh0FK7PPxMhRZTSMMc4JVU44hfSG5nzPYnyK+Not
3WDeF4noUBWq2xybGkovgyf9oZMQsgvTutXuixLIHUIZ/s1ZS07JyRMjYhiD4Fuq
oLaZKUULcMsYUo8cRF73Kj+ymTlCk2GwZIyxtGAtZwcxOTRxOJn5qRYN4sJ1h7Y7
NMS7lEC2lGmyyNOCbrWdh53W7GuAHWcczmcgUQvzzormbQxrEV9a3nv80QbdDIWb
0p9fiUp999cm16d6BOFVpA0L2sJGjVthvDZIZxlaMapPU70vueKgYEFIdIVm233n
ALQYA0DeX71GL2zzDdGEhy6hpFOLdWc7OOVxpbxSxGRBqk8otGHO/XM/vQ65+sZX
JH6bh4LhNnT+Udwk7RvyzfLw8rbr7qGnHEOip7a5EP0iyPWRWJ3yrsLWhcEwOq1y
Mf4fqOLc+5ldeuqMjCmDpJ1RW5OcochahDjUOleDazpLLV0B0EzQu6va3C3dLrye
O53/OH8FGrBhikZl46XeoZ63u4+KbEldM7r08pkrXdU2g/ufhXn9bvXaE6yvdR9g
XjglLhQ96H35LwXYMUFpsbPi7+pkwh45Ny1U9yJNX4BagMAqLn9tLcPdH3AiFwGN
WbMp9z+KwbCHrD0CWmdmm9t07TFUFXGvrGvK35oFBIkjyxFd7OOGPhhtJ9cGkTWu
Oz7rZq/hQdbXcmUDTXYkYlp4cTjoDS/sn6rEdqjZmZz8iV8eG4Mdqgpx7zAMSKUv
pd81RkWNp8GU6Xw+eAAGPKAbSmI/0EICId+vhhXSAleU4QvMvKr45X5tKeOgqrPM
8xhcvACnSKvQyD5cYrueVV40RpUSq5Z0dFTFMqi2MsElzjrVNZSLt1rTaAzhIdav
/MuhpMbLrtnUwyNVtRiZ4Kbm0zjzmZKjQVGvPxcpi83tZkvRFvq6PrYKEO1w2uPQ
pZbObUH9IMhbZ7fEsrp1801NVzK9mayzAB2ZlBXCN/9/fwoojc6wdQcvASaGnrml
268sm/Exa+zRJElt9HqCp1h0FoLXmwz1YU16RkGZaDDfsjVZMEZ1Vahi3QbtgIDH
uXSjPeOKfv3JH3KVfCPvjPf8gcMxQt5ApwwEd1pXfPK+I+k0/fc6+ZWrDg2DyIz0
K7c/mhy+O6PrYzKBAJdpYwSgPp8v1YoU33hPINYqPftR7H5LS2XjmvWJ4RfCMOQL
J8PKIeuksapAVW1PHcdoSN+M1hxVCpMgH7NttEpQYxSvWMaEJel8j6uPFePbxqHW
XC0ebUUKya9SxTftTNnMZiu1zmUWYWXgBPOIGAt3jRP15V5ndToPVrDq/s9Phwsu
xUUhZmzTTggWWPh4J8V8jEDdjlA43RNu9zUO+FE/PSAmjG0Hca8+qDyD91lxx2/8
7Bf+ffg7icTZBeVDUSikC+usLHfzcnMb+/Zfi7gGivEh1M/WSr9oz2qsNnwsjylm
YhPTq1VILaZCbTmg8dPjzQgM2tK19QyJZK52ViugozVyg5oOw4Ngepr2Y3kCtbl4
UdDvCuQz/2B+PNN0IXFtTrTu1G2yqTtTb4Y3wDsvPR2Zn/zG/pC8cg0o1AwMhgTq
9d+ctUGAPR8BykieEOWfjKr77gpp8seV9hfD0aclTG0q1hnkMatnYl+PXUFiP1d7
UImdEbUzjjm7AaNsKkaJN6KUPPnwoukUTCQcZmV2gSmbA7XFpxrGmKmUwkecgTOp
/lkdNvqkh2KVSB4oaaguCnwcxW0K/oCjY/wDIqniszEcoKInqX3COf+l0zUusJvF
jXkCg8etzC4Ri2yqfHMLGXPGAT7ujdYjLYS482ZaVZW8aGTxGZdZSPnQ1dBe0/S+
UT0HPHgnbWLjc6R/Py9OKod9N0PnBly0UjtNkgd4f65nfMf1cdbi+ctOvTvvjg1k
6BQ4sa3L1uGP8fE514R6dDRXXZyKYoaSg0S/uz+aXoOls5qD/xB9ZUSqJh+J6TqU
1o5boWWyp4KosBbYFDqxASioxt6/wWCzado+2K4kaDltI10MIm9x/I/BC8l/gmb8
GagFLwSETJrVnq8vMf3wlb+RyE5k9ETos+JInlhA3PjwoeUHWVfBjfz3Dq+nenUs
vD+suGmtEVeeUOGWlniWYYmg8INPaaplsH81b9hRpBdPwRdRwpYaEjWuWryBsgxZ
/vN3pFPZQOSxqyhHNSpSEkTPC5bvUUu0mSWmapmQ7Z7UeIMAQudCkBoadIV/A1w5
eNfJXtCgXw2OH0UxNfKo1zILHmzBw41bQAniklI/n7ImQdnQd6ORfgVsjh93U7kb
eFp9FtbO8i0FNR/t9kZ/pLXuK44wrGqo4kWHc5Z55di+4TjZaz9XRuiUtMQRd570
Dzi8ahFkG8r/ZtYqtHdVWTdFuiQlo15inM8f7mWYwAwuJsitMylmGI6r7eDBMSaw
uUh53o7bTpdhx4E/du/YnFwGbAQyB25vRu94jDFXM6wX+NZAQy8+HG2sANC0019o
VEorwXrifN1B+8gjOEpxbDWnRBl75qTsM35TxThqKljTCP2bTe7jxwVni3QUzY94
CHi/hDWbqbeUIE67jQ00XyAko8pveV3Y7AgYJpCA/2l/53WRFhGcZ9KMeZbcqNMS
wNtUqBk9YKmlq3Uccgy0Nf0XjLpQksZIbKPrrzfiffFjL8iSbEVwJEx3+bT5oGAJ
O2EsCGqVb7EpZPpeFHk7mQ1O5ks21EcBWKuaGoV00uMFgWGM8LoBiSfp6UFTkviE
jRGBQ4kxAjywMWWdsV8r/h1FASiCxLun+5xrRPn7VGY2BN3lTmsvIaI9GRW1NlPY
iab788Tb+LisIwke0j1gSZ8/GiFPdBZQl1gsCgiqnBQ2sp/ulwZuoAxEA0ANg6y9
xma2m9a/VHiAB96IYcABsedfowEMKtc+xICngMFuFl2dziF6DDEChLMdQH8/fZHt
SIP+Mk3byGwkcPoE/pGY9dgXeeiWA6kn7XGsrNlwWLijsUR7tiYIuGswyCMwnJnV
h9kflemA5XFs4eFM9mQB+MNcNQV+yvFzJ45WCZHWsiN7mqZnqdHiTRLZBokCSkAn
t8YKTYLqk0FzysqWsmOhC/Dm9xoD4eFSR0cilz2PjCHyTkBScKLUDxR5/U3FoRuH
nnen6rd12xy9+S6TbquZHn9kSo9pakEJwS3XvP4K/rpK5TJzySRZyO+rfdzOlGXu
U4SKRztAxNxOzvRgqihEM0xnwFcpqIqeetK4mJvSkwyAR4uxSY1AkY9RtUh4nnmA
1RfBBWLpIAguQp5Dj+REhJqNnUpo61kNzf9rBzNFKGAlqeGJ27bTRiYLZDjd2/sY
3t/ZL43WNckVl8dzd0uOFwcFDV1WstxWWVy+eIiVV+yuC2O3NH9U8z8gRQR1puqy
VylZV3qaAqye+t+rqtwyY5efVs3kfCSe8iZnPjg4TsnD3bcI073CmSNH+YGVGK3r
FSS8+gvgfERN6EGH0e8eJoqVtQqCopPejw8Z7QFa32hK5GAF9pjBi/ZgW3zFvIiJ
BkhNSWvTapm4ByWMwL51eLB3LTp9F+RV6ZNq0CcuB5vM13JN805rbBRp+WT+Pfg+
v8YvoOCnN4ddov26cstTeMoFrzuEZOWOhjACn/ETucg6TDZ+jQHNSFfy+xASAbxr
XbhVN0tDtsd5Bg27tQPm9ERmwFUyZExkI51C0bMjd2fYG1v1ZZcTgeD7fkyllm2J
e8BoLTf2t+LHOjLsnMYosmYOBK9D+OkSHQqlOb524pblvpqgD+Js2ccKNcYxVeMo
KjDsf9m/AgUa2RJO4ByaHeALfLP9u5Bed+N45/kMpB+sQWyrfVq9hmSybN9628jm
mz9LobNKoPvEattb4OSE0ktSXrcmK5Qm0PqeKT3S8/EIfQIQArSfm5vkLH6V0b/F
RvG/1qlUyJUmt3IhRwEWLdNoMjzMoIESWyERstgdrHJ1el+uABBarrwDuFWwteHp
AeX05+2ybIdzf6AH6TqetRJATm1RFTIJvY1w6KJ1WO2TUeig3ST3HrJwNjFk7S9w
bM0PIjzUSNsMj+v0YuOYOxXbHRCZ/GU3BnFZOgagQebg099eLcnj0+EfEzzoxK3v
2dGY4dqIhwsMM+g4z5zyUIDNxBQpJDzy84VfVmlKJB/NClhTcRY70SFyHgB/1u27
1ABjWJact/L+AlTTQPGH8nwspnLZzkhqN8tpFPlzF4X7z0c5yyv8GXV87C1HY7aP
zMAVyW8usqVCZHPFSiRz0iN2s8URXEaJgX/n52edih1FqIMZQTmXqos1veTetd+E
zn+j/Gviv8dONzl8cgZqKtJdQSess3W+elV+GNb3b/8xv8DbRaR4yOsEk7VsMIoj
dhgRsdmrUmOoRYrrBa/5BRy+asdpv9eFe0JLWCac1xWAEWALGjyM96PLaSmjuvYS
zK92Z312MKe782d5hKfBcOJzhb5rNHEivqOSOGzn5QBi6Nk6IFUzuGF857MviOdR
JxH92u1w6nOEX96vl6naZAbNVsS5DW423RNkkfr6MbrrcU7yjNFA7ZvLoVg6kbgo
ZUpbU4U+FnEsiEwuu+/0eTvIv6dV9PvZ68nX/bxPR11DlpCPbzjFYgbPHdWevXmq
5P1LkN7EmlvRQ8zEWeZFaGRoHeVI4PM4stQXPImISrtklHEf7sAIdtP90RTVucLh
0zZHlMvYRtlZOH3veshzFL24DhoXg2L8jZL+fG+Y0crtRKtZ0GYzbk1hYFDQoUGM
W2JTixvBGXJmP2VezcHYKlUbOZbwpI0904nZDYEqsS29ag4KYqz7uN+eJLYsb0dl
iisvA96nMXqiOnjrTcmJ7GnULTrGQfYs+qqV+KBuHDG+09u8VXWIO/G//M+my5Mq
TkqeJq8M65ZV5mbozEglDQ3+q6PlVM0RfEm69EJTCq493xxXV3+V2g9THpVKAaaF
wVN5ZtMfQ7dUWKmePneB3kPuUCTmFHhZ47mS2me06nh8VEN7+VusOufP4I3Co039
9kjBO+eEZN3ZATtgmW/X9F1eaIAu8foSPd9GDbCyYUoM2R2vKjNvuhrv5pUXa21b
0ORGaKkf61Y80Vs3ZKlXfxrXDQsOc7HGPJsCfpuhct/vZMpWIOc5bq/zy60w2y5P
O9Biu8TNTCGXkzRqa/dg9/6+uEt/Dxp6t9wCmn0S1VU/YU27rZwWL8LXQG2eFbS1
lxj3bfjZug9uopwinip8+M/hXMbq81Kl2vKKeY3HydU6cGeeSPe2bscGcxoa+q4p
KdxBjm8tB5wMKG8xXy7mB8YGMAaQRcHZB67wkIRmftKYBF+9KQ5qnHscFX7TRTaO
mISwWm3NdNbj6/f2LhUqrdhYMvMYQpTNMx3oyBUEegbf+N670utIQfyM7uyAr8n9
FWALC0b1IQ6hP4HHoWJdMdMG2xLynFOWXCc8aVbOFAWWVpVtCncMhStd2k0uFYSc
MCzjPBJWv5QvGfwqiqHpBwWbJSU0bi/+57un6RkWoUGaKQ4VxQVTd22sh2bGCFsf
qCzUIGIW2UD8GOn5jPmh0Kb/8GPi8u2WCBdQhUak2s6Sc1UAtuSN9yz+fyPiI9H3
ZqZ8W2fuzvxluj90HvN/iveisGIijopJnnQJWBUyNLlsafCwHvVfgOyXtVgMm1bx
JxfLhdFNdKkQqI4M0jyUiYaDzMkARHvr3k4bzA6QomjJwiAoJZKWjmAHWwwQkElm
sX/dv2vFBIdE1li63Pk1PC+aHgR0qyTQ/bRHIafdv/pcBJdJv/n4G3N3eo3L/VDT
9h4O1ZcxFpwoykJEBAa4WJ6sUgMWhFh/qvHoi8x1iU/nMQWQNdWZMtYMDunt2N5W
lunzIi2pdO6D3Njh5mhCLRBzMcdG0gf1B5RbwnDFPxL9DoUR2HPMPk2diPys5N18
zA1jWbUyxWvIdenqW5Fn3LT7VA72yDoVSkkq4BW3JB3jM5w3C8eZN/zVSsXGIaqB
ri+GtygF+Yxmex68lVXlNwQOiYiBXnMdCPnvhdmYdQV3hP4EvNFobj9Xv0K+9dfe
B2VFlEVWxV0tMfsi1YEHYFWWxnBV3WgT+sw7q3vp/Rl2UiAUWTN4xHQyLtnVJr6x
iS/jahjSAXl6YzzjO2W8Sq5V1cWopz4FQScckQ2E8jjVk6zvjVTEDKyLH8jnR1tP
ibIDzUN2CE1Ey/xhpy03upQtEvRomGCdopASu2T7VmQiRcl6biBl1IDT4awwDe93
Yvq1mqPjEhAkK4Vgap7l2LkAdmKFerVXQu3hpbAFIcmkhDt28ydu1t53e6vaef9J
EdF+s4tDsLU9z4TvkXdIi03DuRd6iZJM2wqPG5ULvV08LfkcnrN7YKTz7Ogj/XZd
2T5BxbQSw0u5zGiYUdD6OqlT67y7WYbUqoHEKHcda69MPaVgzkL/JUXx0YS5tw2Q
8Tlv2/Y7f8omEQqVIq4HgvkS2bsBB1/kwq6pkSsZYNQjj9ob+BDx1F/BkO6J3Dh7
h001fnMyges6ybmXkIMfgxXOCTiG0v5QCw0EDnjn4LNBPd4omtKHXdHWb0DCyY7f
8xHHTJjMsMEeb84SdvqL27o5m/eLHKIFD1BYfFRg9GPw9Z329aGnFH+znzNAoS1w
Pl/aeqbWKYqsW+efK+axVUHRZ73jmH6+FLQ6/LeZ+JMsSxVsfE1YRejlE4cwewzm
SYiNJAuBAD+0oPOVpqy1BqCxglmuBP1tqDUxlrHNrXE7mja+R0Kk7KkVRFMqZ7ev
EFSqF+OSkNjZuCL03Y5vZSjAm6d6lkUZLwW4pmUD4uJutUU4Q9/aQZW2vHS2r8Br
yrFAXbdSeRGPNECoNWBRDisjgRm79KE7QHEPlwf5/8O56/HKm/Aaec/VQ08S2Gbo
NCQ1rpUTWmC+lyLLqlmOAjCmneiJolRWszIG0FZBP6Ecqf7VStA3gQH2U8E0jIob
bMEYnsosgUV7clSteQSMJH2NjiXDCWZHF2T8iNRX71k99WIKbc6YbTxKMCJ8waxL
WWW5Hn0VwNYXMZvDKyYSTHL2cF1Bi+vkN4qGZasPd99kEgxyF+piE/OmYDywX9zi
kQZ2Ik/IAVMELIn1cNSmvBoEsKhp9TasCIIwak6hk/4c9xs5/BWWeBtQxtkViMu9
oMLMQiveVTaQST3KPK78+cBE7BMyTx2iXjySn2Hg8/hKqk2Bxvl445hjs9Iv75hU
nKvsiM5Dh6E1BMa3SWHAnwPVGf6F3h8YIjeGXwK0DzEMvIhcLCBPqCNZE9AzE4Vo
0zKKHNdGGYJMD/Fd7BykpJWxksm2vU8on8W05TzdKk4ypo+Sn5j8qAkCWEErvCw1
3wDAXxf3IeVjiaHV1uuRX1P90eTyIFUl7oO8UOaXE0I/ZMSv8+Cd3Z0ZjvQjRUm6
soh5h+pqhEu/wI8oHRqrDYtL/KWaNnL74JuDtBwSc5lhQ9UMkdotPPJiGB6o8NUQ
tSgFv5UemrKfBASn4lToysexsDyMrlWDNEXvd3w9F4z7MpVsHn3I6f11/eDIVY5i
Y0idV30rLttJLEgtd9V+FK9fFHK4xlcAjZYVl+xiTTHx+jdlRk0uAc7XWq/mx5EC
ozCEQOWqHOBs8PRY0CB4GhPk3ellzYAfgWG+j5GayveIP/ad6LYys5NJ5jukaqiX
HaaNeOIWOZS2fPofGOr7DtsareFVyyijcnORS9EahMgm+3z+d7Zbc4FAjuBUoLv9
zIplprEOS5qZGaWAnyPLtiX5JoKEzncJ2mO56yrSCepniQcnqCMdstRd6Wfa/UTv
798B657SqqIsXBIhsnvHKpdH1TAn7tW4+uuECT3U1ES2yDwTXfVNst7BygnA3+8a
tfILeUCCvRPTwIbn4rw3gTZboF24S+lJRiutOErKOyTX5xv9tkKrW4lZL9aZAKMZ
I1Av3ceZL8Zwtk0+0zEMNjiqYAuxf5TW5PcAK9viI6qgoO3d5393LAPP4W5cRKFB
cxvGWUz0u8rKxG04FHz7cNpK7KQZnh7iJ+0hLFdxBqwVWpWoXHi3OccZfaimLBRn
9Exw278PsHTIUyy6QpXMJiF26+rXHabnO84HxyRRrLxlrTiN+jOXB9ASjjw17g3f
tamn1Mx1a5lmYrIlAQdFdc/XaOAnskrLsrto5lnB9/OiDX7ilm+2oipasLun0dcL
71KWW9ud1kyqqi9R8Hs6UgnXIc+t2o4AfcIz8909+Lvkv5qGqT2dmLlhEuNpo76U
e1pAa8NM7kEwUw8DHyOFPFA2xrFI+ze2EKG/eVgeO64FeAm5UbH1pVUNRldI8sIJ
24fhdQpekJGcfVa7sn8TxxbpYVfNlNLPsIkwxqMpqAEzJ8fQrAy9zzLUk6aE9XLl
mB4Jxvcde8VttYz9W2Os5FQbkrGAmV2JE3wiyZTIJobvcFOPS6av78qRDXnd1ID1
JLkb556HwvJxlv0g20ESEC6a/445CW3wRlWdSav3y23A7tgO7IfYSX8+imVXdTUJ
gT6qY6GwOKpZQ0VYl9kz8A8EHyonopirjoGT9kBkZCtHzXbK+uMOswAI9n8Of3Cq
ZeDdGMAu1TCJnv37vsfwmhPWT//TwsuxHpEb2JxHxFoM2nfM+vH5FqfZgDCwvQ2x
gtRbQTzX6EGeET0f9zJRHObthBXMp3mXt7tuzrSwQde4ujd9rXHXM3qIN0gucBtp
BO8XgtfOTmZGTC529LFYyKPuH1h4Rhcx3SAAfWFXzKIUJfadmZM42ftIWxKGs7kk
Y59MDvN+x9Ei3w+eXoDgQemw1nUipV5U/iwfT71bNCrS/2cSZGmSz4bsnO9NBor0
eaSqHCkOtPGeQUPNYrREV2rMfIJa1riP/bQ1vb+UCBiPlXWPl9D/iy/Ak2AkgcXv
eWzQ9EHifFbl6szO0xnm68sjjoenYBiVaN7ugb3W8Lnc5/BiUuFarTx7D6HOeDyw
w2p23NAXA+DOzx70a8f+4g/R8g0GB5oLCfCFItqk9hrmdYvHb8HaNsDOPbOSwF8l
b7BFKg0S0ZWp26ss5FDuITWrv2qplgk3CfHA0Q1S9BkJYVlKRObADb8ZcTJCQ+G3
gY913wNKpoWhp4s42TOf87y7o3jjxZO6XBqmbDParIzp77tasSfEUThpud38RPC5
Ia6BSQ4U+2iyBFwKs8BgXLEsJrEYy1nE0dxi5kSXJl+YTEpvHT838c/yxWqDBwTl
LyAnI+s9EfzwLwjx5j1F+y8rFMTKJHwHTxXgWIfSXQp4o4jwjSanrBSkAXfj5Y7Y
+X4bp32A9XA1uOazZz+vk+A92qeBOag1LnTpk4voMsxWUvk3ndJy2/pHyH96tG1D
Vf0eXYwtjpuDK+1JK8+Q8URtTCPoCrN0r0PneEpyu6qss83Poez/tlNngP+KGUVv
aM9eJAJSVkmcjb2IMWiaONSJ9g3Kkc5cHfj09bfa0zwVclZMFoAgrc+l2K+b8exb
zrx/OuUtPQxXCDAu6+aotXjOQu/+G6G2YPoZ9q1xvsAPndzNHVwkG5NKnnXa9B4x
WfFwIKyAl0Yyj2vbpJBlwmL/BqPEnPjtiBHi8qtHrx99xkwBYQcu9INFmzIJQHGq
nn4JLgoer7HdCP69ObJJRWiEwFIS1vEaB6nf9/br2MV+fxbV0DSkYwYfnw3hPTdn
kDqTwg4SCEEyE2MgeOuN+MJZ2GvRB6t3fkDdr9dqIADSFKEiKXOpp+85+In1SIfY
8usGrdf/65u3GgGQG1htzx5DvHpEFbr2PEaK5KwRSELo/sfddG7ijZwMdDtNO4OM
Xt0WA8dQ/fhj29LiIMGhLYYc+NBSAmi2ww/nf7WMtk+eFqEM9Nuaimnu4XvHDdUs
POV/KNPpBqZ3ne1Sk2XTC3UCNDBigFhhUD3JG2mFqmLN+vvNphknFLV7JeTNmMKI
HzOGRWwoFdj1RKS+Y2be1+6xaaYaJZjkVnY2RNNkv50i+DzAuo78JHjEAtMdA5u1
iREtV6KzKLY0cuQlzAAejJ3Nx+03OW2YhQzGRi1KvgDcvPqeFdjWYg6uBN2kdXkT
lVLIAA3Cgx3gkjKzqiwCSGM2hsa67DI6Dl5PVl4z4Gd2usZBpSBc6r4cCVC3UIVJ
hP4vZqc+ixXR8kiKakQJ19Be1az67mPytQ4D5rLBrYaA3qrmDw69SUXK7i5Ja4bF
N/a7OYz/EoXVoIf0D7qGQsCBUbAr7NkzcF3PPGtFztwl8sr/XIIjmRHonPg2hwCq
7PbpFDu4tYLtYGh6E11jK/5Zs1JNCLOsa1OdQeYCa6YQ9b4zPiERjFMXrKLQi2t/
BHxmlpAvJKbG/JsoQ8FnCk86xDMMLCn1VvS1Vtslfaqw7XBbGzP0aR7P3neTy5lN
nRFB9/tkX28kEF7TyHrQlklJI+JMq7j4zgGjz00I//QXXW4NkllENQISofy7e1bb
lPjfLj+Xj6TWh5JuKuNUlkt3oMLdfaGsV/IkpucUrd83KeeITvHR5AN0RF1njazj
t83CB2Ba7evWHBEMc0thI7/lA7FghFucbSOJi3T3mRSgCKu2/+R6dPGH1gj48e6K
Jgk1JWhrnjlSwQPZLZFJ8Zf0NsVt03WfT0djCwzg7ln55KHRgDNh+3f+rQWrOO1l
ztLnUsKa5NYUa5mQb2r0XzGeo8//6Jt5y9dEnxe30mRTr7vUAF3dkg9hFzArZixT
whNKDdWKGfsYHjoHkgI46b2VZZuC1xZtJCYwzKwrEmLEMIDUgrpuDgvfJXDstd8m
BbXkjiG0afMnEtcX/vtrRQXpUWUgbCmMlAP15wVcuF8FfHmwe3Mk475DPEhjaike
xjfpthv5eeym76o1a0QCDg+qwf1hG+NcpXIbo/CI0RUf/CO+Q4IzSQ/16KUY+a42
ZAlBqtBA1s7WeXFZjIbeXmNegO07vq6MHpsdrULOOezVHDpnQpSsOr2IUdEFUvbW
hVNfYbwADcBpIIoiiOFx4ndCzExLNcTV/YEWYRp2AHe6WOHYgueYpthpzR1+/tGq
khqJYzMTXIMTS18YUN19lfSJqf6xzf4lrb0V0NbmirOriUkY82hV+y1Kvwi/orsd
3tfHvxm+Oq63p+9Nis5Smc3E+26rYX28Imw6cL+dKj+YyZ7d09jAm0plNssjGekZ
9Rd2L07JHLcZmeeHHQXqJtKWV0GmYjFAlcT45FlOWz0XJqR7A5s7ZNCIGJVEu5lx
9Awaw1VxNKS4EqydHFGrsV8d2NklwoJdGztHOny/SHiZHtfQNVU1XWbVyNqz3PEr
DnMDpM+gDrVENt1jtla3FkiwYpbyD8FG0rMIBp+CanbpXw67FxuWytTaTOY1TNJW
pCKPXmB6DhYZnqIbAe5OmWllJ8ZosfF6TwZ5N0lkdvaEQqchcdU4KJrMIcKvq6qp
nsQUQv6krcySHQMtD4fH6Up/JzNEbrrsbvR7OGnFibMqrCwoFs1F80SahfjyxiAa
NysUTR9lekHBAfGTfHjZ/vI2dJwoZOsGnE8KB2Ptc6M9Lr4iumryCsWH+Ox3C1GP
cztD2PWRdK8V9C2fQgXE9ieRQpyf76eiFl2nX5T2TZzX9Du/FPv3tYT2/2J4QmAZ
y9DqN1uWh+EZH+006jw2BfBjc3a7A5eWCDLtDVJA/Jv1rS335tiuibQwrYpPusTI
VTjivakQj4OYd2Fw8p4L0i6XnX+ywrXoBpD6/jxt0XxDeejB3gXhisSSx4SdaT1h
I7//NYXP0sz55cvLd+ykDBeTqVupyrqm0C3HdXbcBI59TZmpcoiXKE5kWPf0MEaL
gvP0skZekEAttCbtRjOZH6kNgLeEFWumd6LnGvhnOxLRZNICu0KFJQRItxX4mHbP
NAZiUgYE9yBjz4kIBFDEVqqGPjCxLbPVqnCPaMuwian5HVcb6MsPBc4g/akxL+aV
7/z7XOv+LB9DEV6dP1cIx+FtxOFykqj5e1kPrq1HZj7k2ooS1MkDaQeongVodjMB
tB7Z7SF3wMBJwOHsPWH4TAK/xVVHEPJw/4VBYkhM6cDS+7ECPAJuyBV2rpwpTM1m
26733KmxVXyvQgMAs6x5MEuQA4pPbYL1zvyKhLhu0IFuV5BI71wT92x5lfqLkW2X
pnbopwnBZ3lb8FKETQlJ8Li51zbrZBKK6/mNXe5F9v/3NusExtvFCK9mniuee7ee
v/pot7TbYOLLcwEaYhB72qTn0ccpNhG1DAOStzpksb80ke31s8ZJdLT7ACk6paXd
h71Uq0yv26R2hMk8kXWe517EB0SM/MdzjhSLu30ILoEpqUZnxtJSmwlZAVgP/z9I
wIYrDcANedz8C6X7HkFmpVe1qGY0PLpoWbI/nvwjEU/zRNUE8Gpfq6K7MaqRzT27
PnldlfTAVpPP8gqS5W3g1RP9sRficL2wzJ4Fekx65AdQQCqTMxQkAI0kHdgs4Xza
w655uXbt2dAEQvZEV0Nz+FTHMbiFG56BRahxHaxz8JXic7avZwHfCpv4Owh4kVW5
abVP8T5qkSkEsTr72TO0DCsi3q7FI4QOikUsqxBIErGFWXB+VDEhX2qaREk1/MSS
Rd1/wlX3QFN9fMycvURuIT3Hbs0vwsaaOzVTvG7Tqc/CaKF/fZ8SinApV15p9KI+
m+y8jkB381CASK4MmF80pNbtdDJ2+5KbfLugryKex8pllq0uZXkDAq9lT3y0tG0/
RjM3aH+qulF/hf800Y3ayJ+xvLDW8qKkhjevZz6jKQOOb6RJj5xABiw1h0db3xy3
cvc7kPymZUSmomM4vq7ciuMpGIlc4/VUlidCMdB8qSE/FxVuYh0iRFEADHOY7AtD
CbcqU4dHbfEZSx/nMQXAb3k4OstRbihr5tqfdrm661kyXL6Y4XpE7ImgHCb3sLI6
reJ2jmRCLHgnmvnk77aYVv6F9CnFr69GBAaGFn2py7pRDTDV3aOAteXk/K7WJMbS
vdiLi+YA97IkYEkbm5z3DoqvwvViKNGjM7fdnHWGJtBrLZHY69jU6RcbV5eVLJNt
6vCIfNn9vubbibZyUPuJlxMvW3UKPy5g6TCXTNoSPL7MKiP+jaSgeWw0fD834bsk
65UDe/88WLwZWv/Rb1S/OyDj2vn1WggyufKLN9DJ8t2ZZiC2k68WjkbmaVWXm2Ow
KfvjI1f5fNKEiHn9o515WGEFBbYxSMukePbWkwPnfzXOSGFLyZ/Gj0ZqhYfRGr28
iYcTsKg0HzZgbOgnsIggrYWTk3WShy8CQ9vVXdPJmsQ/Udpsrq4W80wadL9B6GQ6
k2VZtQC5pS7Rb1Ga5tvMM49s7NJ0afynX9v/XKgWpvoffCp5tAm+crEC5HMLq6oe
o7BuuVt5Po6AFPwV1JUN/JhbbrUFpDSEBPQu0u8keHWdsLR31JN1LX3ZADf8hvP3
CuglWVBiMRg4RlnjntICYH+31PCb29DkjN3wo4uHUHTPdpyS1zkQcJZhuJCGhY+8
ZLjNsP/ECMKPQErQdf0ci/Fo+aovJr5PPQ+6cWzQEmYePdNilPMMtizCUb+E2EqI
CSwxH3/j9dodUXYFRuFnRvFpRCZHxnvK0Dl81yesO5n3ZwEuMzICkpBiK3EJNVjZ
Nx1ibDMsUH84DrtSEun7Ak6NoRXdjwfuWpHrQaFhQHDxuvTNCcbPtorXPo4UrOPc
q506Hl/lYD2Uih40reRIRHomA3nVYaWPsCoG+NTqd8SImudsFzI3IWUDMXYHys9Z
PJ5lim6HzucP+rS1r+sJPiuUd6oM3/ZzRzFwEMrhTqijryvQ7BPz6iSdmzYBYQoV
YDNb2ZgBqDT5tjE8vBzhgCXUJnwJoUcg/NnfNo0CTv4cjhL+Q3WMps4ibAt7JBOF
uRGX2bmgJ+7ctXwUt3PeSdGDxhSG6k46vLSmavk1K3rAptGndpfpfKwbUEovqYwY
CJc6cJ867S+euiv37dvV7AwRNH/mpFa1dq0QWlgxGsGzjRlQ4wxefcYI/oJWs6WS
LaGZYn3w6RFqT5NGUw59jPl3eUJ4qNIbFkxXZed6UyauUwEGsbS46nCaONQM+D7K
mXtdNNTY53k/oy+jF7ygOD3DnP+s/bYesKLpYSY70uHQiHsr6q67nAh7LyWSiR/t
KbCdxtWebpOaxOkyION/oin8RqjpYcQ9WWnuqCD4jBvISBNABTnqPqz15y3MUhby
t8JMI5QP6RURCVGvQfpCdEfjNqNMlPUBjcaLgqson0Z6Ld8GfhKGAzU97KZQiXD9
mE8IigcCibaE2VyvEb3lirxrY6Qo9zeqtcALIopjbVhvQ2uRJ93jmhSbC6HhVlfE
XXA+gkY2zNV+c3lJmudAM6Y8I21hU7/XLbYf+EJcLVo+ZxQSJqe9hQTSuydW9AOW
tGbqaAeFec3mc6oNo7r+Tws5E1AAM8YsaiwSoD84cF4qUwtMq0sp88buQh073Rwa
uDe1yYh/7ClDnjmWhmyKFzpJO0UKJdEKQ8yXFHl3lpPgD2XCXAqYxesUbqS8l+t5
HirwQmFOYXUXHbCQjmNzWAu96WwPR8Kj/uwHnkVzosbnM7gYWoJKJznl1X5lB3Gk
rDkjB8J8WjuQnPSVCGPVfH2ybesJdlDma81UqDhAN5KvEPbSa2EYPfGKJIBlbA9O
sood9xFMA0g35tqrcFbSYtbFUwP+Y0NdX+xzgHCKFM6KzR/pQDZsd+8G5a8HEphl
fB6miZBGDr/EmWNqXITQyh9gKrHVUdrBdpUyCFHY53wxvxomXMEG9G8uNPLTFIye
u7dxcK6T6FQNNOy6DsJ0w03LFYaCtPDtZmBmuH6mDiy7MPzqNj/2IG0y+JJLIYAt
1z8D+H3IBSwyuXWEXS+y6NPhIlD94cipKXEWcMnVqi6n56T6c7th4o4ijuC8tsbD
T4TQv3s51rCTnQm/mhSyVe7s+jjlw5U/v4n92DacRTtN9X7f5V/NJCWGGJSnqpfR
ZBzyCpY14q6f7ia2hieSsHnTJAjyunrq5rdj1QB1wPK5dfQwxSCwWGP1QNu+RbKp
t7yf2d34N+Zks5gXZfGSm3FlD/70niEVmugjna86LhzF09YOMxFWn2n4CtJr8SNZ
EUb2y4+iWI1Ys3RUWZfgMgk3aBQrre9Xv76iWukV+WWSlTBziz4NEtbKKmjphpF2
iJkPeNUL+ME4I6kJYaPpMMQNMunT9ChMWmIRjwTf/O+cfLHWeZ1JPSIieH0IEXBs
zxLS2BQI+Jy7c0hpV4p583azxUliLt5+M8YqS0Q2+/UW3wuQV/v5F6BI+X1CwCHc
aEjlZFHJkgoNUZCcKHDkP8wg6oC8swIrA4Niuivl5elRiBJ6Io+ypiBK2ZTE5ULT
bPpTK9j5pX7oeYjG2ewF5dEL6nSXggjMO66mZi88cwXBNow5evGbgh8tAGqxZx+H
qDhsEK6OIqMZxcSOUQt9srXbo2eSYOBe3I1zAS3z4cFvUx/9UsEsYhNTmpFE8shM
VbfU5TlKDAXt++5gvSvlvEPUY+IVyZFpUy/ABrMXwknHONIHTfscXpDUgHZl1MHO
8vU9h5zFupk0Ytc0wADMT7m1Tm6sOL4N1C7ifCiTKOL0EviNtr5S9Z67d7IrEZ4S
NJjahpF4s1GPQI6JDxRPHvOLd4zkyNIq2yEIZpMa8bBrWAel0k6AEU1b9J2nqYMF
bs10Y0t1bNx4i6VEtQDz+XktPQjVfIapv+WbqwArAkc8izu5FjNq1azmPOmb0645
lrLqAjwqVR8c60QxZ1bR0l1avautlK/btYN83DIaoqoNMouXtaHrndOimysegOIY
P7UOwfi7WUfHnwFDdk+Zzx4GMcRQ97P/hjomOxPR782P5+3aRBdKj6cb1jM1+iPk
uH+7mC5pv9Ex1ERoC2Ap7RvLjfDb+qzPw6P8UvB+M4ymo+j9pdYRabJnkUN/2+3T
3qD2UQEwURZ70RvneHBqh98UhVA4dfb0XBA8TX9XIMyKY0oLen6NSSd0pAdmpwC5
g3+IT+JPQyoWi1TooKNlI3h7TlQjjYaYSmTWB0/6RmJUGH8qB86U6K+PJHqAhTpW
wfrTaWXSPxWaZdNQf5yigVDMe1nCpXeyJsGtI1gr9TQf9HiXPy8Y9wixcJSDLSmV
xgpXbCS0aT7ZJySLgxzqZaWxMOQLv894FVQiMBAkKM3/is703o1JVuH/3WGT0Itx
rD3O4FPSMXXzal/HmYGKanaf94Czk0txks4D+mYU6e3C/DxD7RCeaRNlEJ9dSwTL
W8AAduweWEFz0DH2uLlfLM0jtL+cNmWcJWvjgBwzSUT0tATCzMxIxwxRI2v3I/7+
OW09WbE6cP7Ge2E+BhVp5IYYMBXO/AvV/dmmlsJc/rz2B4ZFdvu/VErNknkeE+o5
B/IyqE9NQ4H4g6Nc/g7U1gxYOKbJbT71x/7lEI6PRP01HoBZm+IBSXlufxM3XOhp
lC6htuETtIm7RuFKw3bJxC+3oPn8Q3EygTYWtXnxVw/pk2DAfE4V8ceGlghnDXu8
A53bzd59fkOeVL+I0ibT4tT2GrquKnkcrCM39obuPndhdF2b/wLS0gvGkBgTD2SS
vNumI8utFAK6cpRlxu4v9T/CdlBQcv/jQaf+ywXq80fuKc2dmM9WKlOa0kIUE+IX
O/ahOHqK3Z3sgRADx41HxGuNOFY/ZKz/pL7j2HlvWp9cIbNRR/LLi3t0MdYumSaX
3uNLgAvbCZm8jOgD9G0Jzyhg/xnrGH6tmmvd//nRSJyhuRAnLgc0jCaJxXa39woX
wL+efrKaFyGYqra0OB2ybd95GrH3KEtrbCoINuHbG7cij+JrsV2DY7SR1zbJgkVp
oBYWsX5sL5nr/NP3Jnh2LzsOuXY3/nmtv1tI7/dhNJ2iI5cqLrO6ZCK4oy39dwXZ
EYwrQcJPPRlDWd0Mwlcj6HKlb5piXLyyBnZ8preD2dndJy6/Nhe+wyrOiOSzBqrv
7Q1YBtxDiQjpe1+z3Y1BfaSy0CQDOBdnnZp3GX9QXwaKwP774l0Ny858ZCWEYC+P
cDqEE1c8n0MVsKwyajP2ErDUPAngg93zZdn3uLk8t1/N6EdKhzg/ItTdDHLTt8Lu
tzerPr/PFiSmKEsHwAUY5gCcjC5o96KiN49Frs6/+b4SBsqrRZvgiXaFIbSXP1+s
XdgEfQbLn1T1kqwD6CiWwhwjcj/6cmZwdor8HetHGJsGOHWc9uTulGaiZ9EFW/1+
Gaz/HUgv7WdZlm7YcsvL2mnpMBW9yMvvmB4hDNcDoNrULVAt07zceZJNfqBReI+d
YyAM8b2PmM4xGipRpk7H5POyTLwT39qRACl642dSB8OSWYG+cNKaiYTaBa/W7YFe
POS6k5sl/ZDYaG9mVc2BuJu7aqtgcf0brLEvUGMOAWM49AOHRaHJIn3N4SE+eEXE
n3DkHhjrmbKN3efBxxd1IGJq3qB/sxGOQaRZGzCgDViV6iQoGJKsQHGNihBTIZiA
a2mu1OKrJhP1x5AsIgn2d3F9P3EqyKWvM7htHawI6qtlZKY2EdxA7MA6qED35/og
rCmQy2Sh2eR+aHagryUI3ZPIXS8vSQmKsZDsjxrzo+kahAwNV6lzhM1FqMW0bsSf
sfnRtm0kOJUWpgiw9+BSOAQvnvVLTeFLguP+QOt5BC1xbdkL1/+MySTc7R2KnaAK
P/vUt5SCwOn9b2H+z6HwxvWv5K1ksfSu2Max6PsTclAC7kQu/zwApc+nvsM7QE6U
Y5WcOYQYPRzu4msZ/oeHMm1zcpsIWI8Pib+0Qi6dS4Hvwf6rOZ3w/Sst9fitFrb/
KEhVnemEf3BDtmk3I+zMyzNX71hBM/U1aue0NRVIf6rtU49uQhJIoCQLlrU9bVWO
Q3fagLm1ITEAs5ZL7O+p+izjTECqQ63yW6ozqnkvsKZM7S3YOqnfh2l8r4ZAOEQX
rvm2His3t4n0oeoAwutHcipRvwuN5Yj+PnmBg6zIrOtj5ods3+QUZx2P4RM26HB3
wEqIlUmHEiHj6ZcKwKlPm1kjQHC0Bemz5XrY3LbJHLSTtybPKn8h0eOiTt7Q/k+0
48hpYn7y20oghsJ5Dwr2FkOktxOgNcUj6WtDA4ZmpSckwnOuZBHZHdh7DWL9PX0d
aCaxQ91x3l5snLOqmfzQhpGOutFxRfYkYUE7O78YT7Q/PYoEBlCSGTqKWUIZaA/q
qedpi+f27X91aGPYutuktZ8/+VwRbpMWW8W/FhVCUYhYurStTIu4s0hMhyq/n7Qw
T1jMaJqd6YKbuycTsEIQlE9V/Tb931Ka1KAe1GZHDwvykxSEIvADQQTd+O2vrymI
CtCXy/jr19AoHjy3s8OUGaHx1moK0yPbGenwHHwi0FAK0TbpD5AXDJUFGgRtxmkk
+INbImMcCg8o1bs/nrjxWCfCM5PJOV3zg3AjRoV6UVpz8/47TMl9rxeWjQ6gm9n5
jvQ360T4HG/xqwy8pmjP18b4a+0Su7BCuZtrJIxlfb6lZMbUc8SN30p4c8N8sKQk
BQWPL+i61scgh88vacGsckAoWlb1IBElJziha+MK69+OYyoctRdQwUWS8HGtrJYg
jDw4wvmSEG6rD1YnCE7Mo28jot4pZ56yjzHfULUhlFEMY1i7Eu+QHYMNSJxxpAFh
9BjLNzvhTEKRf8ohsad4NR8wqBv/vgzCXzrFRC83wOE7aQJlejjgwk6bsPlNy5hk
yaPDKDplIKv0xuoc0H7Qgt/926BWk3rzSU7oxAtB8KnEsJadR0Zv9Ip0ZcKLp0bk
7er0wRmqZbrGkloYK411Hkp0F7GQ3UtGhC0lhA4VfMhPxSVy5BFxfqmV91jdE9Z1
OM7lnsKHMYFRHlssv7YT3k6tS9MLqL5xxb9e2inghJniVOoXqC4a7167uJ/AZWaY
dw39lCra6X/EeT5chkbqQB7twnAqvAu/g9rt1ltfx6tb9XWrBXk24CYdvnLvqzJt
ZB13oIL21Mj7MVLUDqZbX3ibh2aXWij/OHpq2VJmTAHzPj9ZuYPq/oKOToAtbKlK
IT49mXeOhxglk0BrnsYy9eeJS1ABeEMFEMcjvmrWs/lCqpljmuItOsPwtw2aeMQI
RwIQLhGFFgeO0B3wF6vhczsT+6jyid3v5N7ak/Vi8PPlfqfHOuh3Tmrt1yVuJSLJ
JNvyAKTML560JXXJvrPMAUVUrJQiXXMmtEeVsCZigIZzzgkyZhGUZxVR2nOyDnFD
arMlJfR/RnCymkWqctX+bMf+BqKKz2UtHZ8mxOW/+HIaaB5KOfS37gsceJATSrRx
qH0fYmC4nkhWEyZz6UBnwZ9ZeBZuAz9tjvCpmMDBB+lhBC028WcID6BB1UW4Xj4R
31e9KVexbun4myBLHmQLgaCNBUsE1ccTMe0lige0kWJ3y8QBby1SV+f0/voQubU9
i9jouQFYOZwrWVmX2RhmouG0+CBD19ZAFRhQyhg6pvY5wERGMw9YAAeDof9zH482
BCJHWikGgxR1YkqhrtIcnMmBXXDL7uN5d+7HvtNAErep+PnsfjrwzOUtAJslAObG
etj3/mYXP+7F65ITvPJdOlMHzfg4DQuBQXCPCCcEkPgMZ6ZnAtm3aQ0VUuI+1bzJ
+RMRLsHOrSwgFFFPller2xtxl4gk35qaxV7rqlAXQM/dGwS0Xi/cAv49/TtZ6HOh
cBPMRFbULaXqvQCwKO1WJwnApwmn9VpNzxwSDKJmQHcO7c08qk/yOdeSW230rOQA
6dNS3Js3LxCaykNbcZ8aAMudzWF/pqfhH8OzN+WmulhoR6S1p9+zbvqCAY1iGiCt
k/7weQnOsF7WLTfpERvQV3lFXrJY/oZWlErcY49c5IEt7gevd1GMFJVzGqksqPN5
MnWAClIKWY6ZaVDe2x9gaIvKe6pm3lP3x1MyY0TSR5VufTW8xnfrvaYmNnX8aLVr
1wyQnA4J0aDhhmCqRrfguCWaFC9Kh/8k/1eE8sC+XWybywk7i+uMJKTcaYXnelic
cCBJOByTPmWKYd7i/Lz6ojrfhxmgyVYnwX03Riy5FrclUs4/PVmYfQKqluqx9FxE
bam6KncSu31VM5iDRWBDzoy45jPUIIBXYxDDgzmE2XggnbiN4uS973mI8Ofy1LFo
GJj2jjajFzfZ/tHHQexddry0Rem/B+BqFQ4erOMdaACtPNWiD0yXh1hlpbtzXMdI
iyGNrsW6MVQfYuYlFvtXTgg4DYOytE38gL+HK7+aRqXO8V7f0CHhaT/PS6IhtZs9
gGRDJHWP50b2YdrHltES6XpJ13Rh5cNb3D82ERbtVMY1jt7IZc5uDWHSsvZskjnb
1/Jdw05+qPnBeXr9+5SYrOYtarJ9QOgQ/rjFUC64yAAkglS5UCLzbcZ8AlSLiB5y
qBuBj8aVRDHRxIVw7XT1Ovqf//OP3zBgnI/wD3hocDeunKxRveGRvhb2C2/3GMZm
5qp3S4i2m1cVro3XdOX2OIg7eITcn/5QgYr5wUXo+I3DJkt7MSjSfq8eIKP9KVlq
GYA8rssmC2hRXn4b+t302P1GCNloMSFvZ+6lPxLoQK7DDkjOJY2R2Qf716lfDx1r
KBqNhish1XPeE01h/y2eGJJjgL0fw7IwnxWlodvBAAT3SwxR3c9s+YvAci40F7Qa
/DtE4uJcDwUoRMTL1+XnqBu8H5Zda5oShKh8MyRxVYv82y6eFH0NwBd55KCDMCUU
OQU9pT12/rfi2fCcRVhBBZzotl9648Mbwl+2MF9EYwTc5WlyjeftYFVC+UH3OaNr
mIp+4iIsjVHomeYgX12kJ3rwBvykkKawifcB6B+DTZ9prOAS48X1BLmGXi0qs8wg
zMspJ0DZfWVDVXKwjsJs7FER9dB+/yfrtWE/xNBbib8nJjAtquZ1KB4nSFwzXeAS
2YcMAY/whCjaMrcK5sKK1xRR+wvPOLllu3gou12n35+aJBKCRDfLnyIuLS74fZmU
7a6xh2u6hNLEeMXgDcIrKEuNH8Ii1QmK40Qmk/EZBmIb3Wz2JJ2KhNUM06s678l0
AajH2z+rWl08wA97LqOFccWNi9zZMvCAMoFBD0f0vULGoZofD1dXwSQvE9i5ljFr
Zn6TQmX5Ws2zNgvnvvxpe1O7zVFtyxFfU1S5pGHnEleznZ8mI0j9G1jofZWge3Sh
3JByC0xigsRR+gORgg+ZMUEPF4S7ovXkCO9MUODJfmUJHF3GmbzjVBaBVeh4BbrM
jebhyhK6WJu3b2f9gua+rbjezimZs1bv7e3F4NU22obS7deMqrN6bnm14u0VVPXP
Tf1M8rHltogGBofHMzPxFP7gG/PXq014VIHu5mdhR+51NJMTI3Q4SbruUbob0Inm
7dvZWSWEgYDsCqwnIxst99gJXpZpsz9cQKXr3bgvNjYcuycVGN07z9SI/FtoHwim
2NgNwJ2hKr78yZ7ZEhRMGVXXxesVBralR4O97bqciD1fJ5MEN/vwkXEqXC8e8qUm
PLxs06ikxlBsPadB6fC41ZmgOmSM3jrnt/PaBrhN15pxeIi3vn3d2QB+qEy0pYEN
dAWk5SEE99OBbGz+mE8xaBBBAhso+TKwfzg+CiazQwqngcMzI/jVQ1/TX8P9WCQT
+gI8CvWjCf7gSHgd/xNFKwAYewWB9mpZsomWirb0YSBJ5MOyB/Y53mePCJLERb6n
huijldm4PMMmxuljoUqoZwve77tJSkP1KxTHUE/DL7hp9HuRMqbudc5phNOLAVtg
SCivFxFtNhSTksRatUf72y3aJW1w7WL6D6EOKsBluGS9btDwBeltb0Pfh+D+bRxC
UCYmFDLbDK1H40b6bdTwNYSpohJ/12rgw/XvdXQn9PaDwhboFAHVbIdQ3ZQfYuFS
tfKzcH+L0Am3FZSrkKIDBxgtRq1fH8q5SMAAkWVWxy/ODHLnmq6ko0ISonH3Xxvf
swa5vbvDH43S8DM/eJaQyk0WIFwNHV8CiZgPWWCdQufP5h4ra0UDSUo0Rp0/sLNn
xMx5eeEQc1fHZuaaeV5NwcnvM0/iSwsjUHv5UB52h6vZUqazGn0bpMnVbKvib+Hq
UvM56n57gLSznD6p33ym/5iUn/FLKVxdfD6SIVeHe5Dp/AxyKvrrtB63J7DB4rRA
IYrpWIbDYe3x9nPERa1+cwviz716HLr0KT7h0cmS1aVM07+onN1lud/UL08/47iJ
MnfBGJ1XLlgaCSUfEPo9bO2W6w0rYteMQUWVfJNe+cFpy/OyaqoEWlQfe889iEoo
qYAGR+qFjADwdY5EvGwV5wr+go9G6UlMqnav3tOlPe+uS/48AvZ+EiKka2DF3PGP
iix1HdHPYZXLPhaEFeoD+EkeV13LBxeGd68JPT3RLjTIzBg6TJtBHRaisr8Pr4fe
c/WqfmbB85yNYBmyOaM1pwEsfEE9zVGS4Yc1s/uP+ljjo/X2TkIlI+euz5rmk85O
FOqmi2redESgUVOcjs1dcjk/AvrFQr4KM1iHmxRqejy4SCV1+9/zBPqYrJF/+DWP
wvIC4DpbmG/9M7i7Yar840n7r2E19oWNIHzzRbD2fhbIaMAp6xXnri8H8u32kIDx
gtBAe1swPUiGDLG7Rw3SHYa1HLmLkEvKGuFQv3y7o6Mrrt9Dog9NUgKV1shLo8Wv
WrENBGDN372iChcHyEaIAxOFqLFvrbQc24ZDfPaucck+wvtQ8bc6ywJxePogbnpp
hT0QUB/YOhb9Qe1oRrGN+WxBe87hr336lOhfTIBWTgf6wbU3VdFBOxHGAixTHE81
wAf6fHZIDfq7Tp3rjdR5PTTe81IO6lmLUe1oQyvQKIkjhD8aYhRqAVTSotcLjC8L
nKOq23khqd0WZx4PRUD6TGHaM8rkuvHZMJwkvzknBUzJ0jNkFET2MaTXQumaRCKx
HMBg9Ooqcyot9g03Fmg37RTCZGZR65blGeLXAa9l0UPc+Y2Lbk243lckehwH0/+p
4ETApmoJITK35fPTixFoYfkvmkJ8cZbYLtlacMiPhlyRkQk9eYpu/Uefl9CPsMil
dHVoW6X5HDOm2ZBUc31c6hPgHz/TOtcg6FI0izUSVx55r8JTp43lyegvLfJyfqRG
DxLVSzu53j6OORvPFJqG+Tkr2ZgioDBgHXNG5CylhFyWyzVXh/pxkKrrm1ol9qWc
kRtoRN1aHCxLlWozCRmwvNIowXDm6V2DPoRA/1t10HREwZe7syp3vdXuqDH8A+pe
V4mQVZaVqRlinaUlDRCatHoHpK1FmMCLN6+AqLPt64IO23AI5EOw8hZ7dOrASsKe
DvPqhoF1ULTjF12+9i0DIg7AWzLhRJvrrgIv3lLFNpqrjZY3sd1xNSy8EPkDwkM7
rprpi4cfLQIGAsDY0xPfRCyLjvGwl6E+r8/5a9PHgRnSDg/eVtWW/V+bc+o3JyeM
X5Qgo3jgFDXF8kfkcj10BPJaz936p/KMTAzju0DDkizJczo+/UCkmxcWffgUd59+
9HJ0609yoqrSSPbiSmW71vohmNgDoyzbNHs3BxZoFvKZFK+IceOK75ZEQBgTa1cw
d+5Dl0+6xAPeLVNxsvDZbkES8zpYCEswrvUTnKRyu4st5AuPyKVRi9c577cjsZDA
y+UiOttcsKt2/2Lyb9d2s+pnYHH8S0FVVK9wMlx8vUHxvTXS3Up7+ap4/YYK3THm
LTLRWgxLn44RPtAoTZWyNuiLHjoBOs8pQWgtNLcppubbrOJTyXowogp6JmcS5LOO
kDQEDpJ1KV/I4a4Bbt9P6eD94mF0G4/Cc0yXdD+nAaqDsnqdAI6l+/1/XLEB25c4
ecEEcgSPVQHGnzwNBgaVJPzkNWGGnsoOO/njZ6ZGTmp6PiBE1rih4ObFwNgt6A7f
WFHC6+xRpvxdmEE1eSoVxO8g1CuZpXRJUTuoSG+NYqCoLZBbWO0BwC38Hn6/Hl1g
zM/o7mgRtevgqTkhVegA2nWXa/ceHVdh5rNTGCKgiaoXtLr4JjcbqoxB3QKSIEB1
iTDUn0rdWmODiW2CZU1I3h+gCn8e6cA02YDNtyBwfUWbVeoBp5DJQIHopvyCiKHJ
zQmBVC5bI8APC2Eu0f1DUk/xjej8GFg1peym5dk+/233FjnfzBY95/cJ+c/SHraI
uz3ASZgFfS6XsnOsIR4428mnmBHcbCy6wmyrYtQx3wj4R6rrVB3kBj5xUIpavZ8+
XrJHldNdDVriBah/RCOGc01PV0BPvpVZPdqWFYflb4I1ZNk02v1ZhRpv5WdZEPjB
aQqmajH533MENihl8acSQk06NfpK6U/Jn9JVjrBZUYjrDaYkg2cuenh+mT/4zNlD
FlGqexxv86GUNdxuIj4w8xROKBVZyWCZq3DNOyJ8+KBPfonYw3Vy1iFqH6KBvIHl
UsgMVOJdPZg+ne6fXlTyJ9b142AaMtzj/KxAr69Y4pho2YlTJ++1wbMirg4hBrnC
OmWW3avC3R6OYGQdW4hFuUkXwhC675UoEqj83xpt3ZsINoppBAEsY99JKJ1nQguz
+m9nRck5O0+oE5HtMgMI5d88T9DnEPeHB7Nf0a3Cg+OfMKJGuJ9rAlemlkJoxIht
iIQBCMQHZU/SeP8ZZNMviWIO7/Mrao7qc/6ZG6Z+4n1Ov9Vwqc0SBI3W/O3rCMq5
RvoaGIW96B+0uQRY5/wPK8RVHJBLonM30jthMRCi/9sjWk+OzzWNiCaGdiK0GhCQ
5GnidEh4bxZFjf0sdCAXZ9gLxCY1fEYf6mHRJWwQbvrz8GM8afCoO+6ECKSGPTi2
LHTS3giO5kTtQEjhJeWLTI4yX9oEa3bRNwpyvLG+l6xG3/EPafasQq0EeMkAUTh8
zeALLfphE/YcPKQ9Vj6baMiciBnN2sg3cX3YLlSE5JgJYaT/vELcu99/Li9NX0qU
Apooa55r0c+5ackSr1N1JqSYo57GkQ4S3CtSVoZDPNUgD0Pe7hRtL5QmXrfRGBAx
VWuXZw0Jp5FdqgD/DWbYVdVV9nGKt0gvcRDcAog53Ta6Vs+xzyk8SzY/CyIbNtbB
L2NwbXSbzUmBJY9K1HdcmOnJyM1YqRWDkqXd5eCnz5stjcXi6qQw374iERJWWCfs
IakGXjFqMVrwPjoXBFx4r4ygnLk0P+mxVOxZHH/nMlcOuyf1Q8++numRu32M59Y+
vcXZ1Yxck0plXLYbwq9fBf0+fQ48h+Nbc1kP1gRf7kJaEe5VyuaR1CuB2omTKsle
eGgFImBBd5eMKV6S4CQxj2giALeAnA86MymSmirlRw1Uy1S/LtNRkQdg886eAkgR
fjZHoOtM2PiYg8ZOxNNNQ0zIcQAN3WGbmvIpH7YHKN+1Y6DtVvtjOcUVOmlegAfA
6l3+EWzkAKWkpzIqCikwD/JhHhujf4H48yprfMa9KwMJiddHPg8s1+s63O19jq6b
smrSbcqas/0d4Jk7FJ7o2VMSWFw6RRL8+sN1XcqA8KiXnpREZiyDcZdhjV5rfbH1
8Fpn2nDRV4CnFUhC0Vua1rjJCQ346QiNGjDvqVLEYou2cAsfgBCc2QDXZeqFdfBu
9ZSzlb2Oj9VzF6pnlBk+JoVLxjYVIo0TJIHc4zN4cu58HLvNhUf5DYMjwxni0Ai6
6kcJ9k4WwgppkbrZ3Qv3arbkpupBNEMKd9nkRi7VONKZ/xfjGVms61AqCRzbSHzv
aoxdM9ree04p1mLK56YvHExFj/pvVbvfDKSg/NGXAd0kn2JGC44mU4McOrfDR5bF
nBxnmHZFzeqeKZUaf/dtS7YFrIRX7M/FWicOK3NPz5lDymXkZ8+xu6HySKWWzfLK
AwLYpCq285MuVoKtvB+mdvYGY72D4iUHSwcOzCjFIpSqPfGf2cqQeeSuwKnnJDTg
w3pP5VALPGnuB9e3EmBnsD2lupQ/mf6JSrUs330iO1hWWigrikja0pe++IZ3Bl3B
rLY1k5VPGkJP0BqBnHXVNU8kqDdE8dDh/csnX8D6BuFA1R1VN9edUUXoHaSA5dSf
W0ILr1FYy6Yte1AJQkh4yk731qs8trIzBVnokqOFLwhwL3pmzj4xi1GORwfuSKaa
GGzo/eUj5BcvvCcrCjo7BNik5g5O/FYvtm6pihm3oV7a47AX9setam90IadF0b+J
laQi+4NZKF3C0OzvfAt5SP+tpLZslJjPzbaOe2/B/5pNSVn0iohU452nv2bwwMks
YTKW8mZENAN9/cGfKNKhYgSdBrEPMrOE1Rs1x3I+duR0hiv8o0yHkmYHTlPJUZpv
gABe48jBQNJ52mZ+X1Auq9Fo+nMYrudHPcdqzpnpkyp7DBYCni81gEzUEZYLy9tH
kH4QWZXrl6zqqwM4lqo6NESnoOP3UgkAIgnmQ1mu7hKs6GChyABTMkL5BOjgviPC
XgMrOKJlrCWBQcIonxDLLjY9SaeO9nMqKMBn1mQqSynMVSgYG208R8SqkveomdAb
MiX+KaOiWd7id93QY2TZBD6KBjtUSH+/DJlKTl3ZAAMURTkctsWjcLNPMLQHZKii
2Ypx9DGjFRh1hugKnUxmkcuj0GxQ0iNSeAuB7YOVW9DJivjNtXWtbVYsmf5bP5v6
/UeL0w1GNpVCD5H86mxpAxknffiGvut4t1B2jGNMitGSI/Ostv+XcPh3QFmRGgSc
SJhZk5HyIMbAP8u86q8jRhqlgTntfL/xAHhnbR6Pub9x5tWcJaAOBVianA0++u45
EHM11Ml8Pb2bA3nxGBF0hnGujSkG6wJnUntYGgvZCePrVHw4S4wlyb9tF3z+D16q
5YEFaEKThSzKSZIcVuD1vhBd5+E1RdUXpH9b0bV1YnP1W36w2AvJ6ivNnarv5CMN
yL2UcYK576MTVnBmMXhhfcOOz10KWwfHF+P+eyT/r9EIS304QsBaAyGu9nv/Vdql
hWcxi/6pWXmcNexIKUffF9azZzLJoEenKDqClSxdFQnx4vYSXmrDfkYoIu6iPQ79
YqAL3k1yur62WVXKxSIhdJblaKHGCxSif36x/TTo2Xv+aUDQXM2C/pMTngoMT3ml
nT4um8mjFvB/3SJYqLq27XLfzuSLTn/I9SCgrhCU6AxKvI6hhhvj8htQJcpPIQIj
JuSWE7HI99YgH0tcTWsNDs6wC3AK1Hw1Nz/qn4ibrjL/yDC4DUbdb2Ix7GxirNis
xH1Boghh3G5ZhqRAaiLHi+pLA4OB97xahsxrjg28GjGORhkRUoRpffyC5Pn8Jyux
SxK3rs+79eERxB/fR7haB0HtHOsB1kn2HhWehkz3GiRN3beIvvWLIc91mLiv4LJa
2A/WzvePgcf3kFoG+eK7GOWMwJDgsc0X5VapyKv9vUkC2GfqcsIxs4M6oxuHOWkL
m8q0DnA4q0CvR6pJbhSMjz+hWQhCniBvohPKAbBsTfYRr13rZoPBXXM37noWXqE4
yvkkomXWg9/TKnUjIrqJ235gEzKbmEsKElEH8sqN9oDM2zK36YVuiMvKfs3PPos1
Y0vWM7dGWuuh0W0dIxaGmmO+U6hGc0h4CmZU+cuFJyVNsnHDVv4loHkHx3G48zTa
l0zVglsRgHRcUZMAIAkJFzl5wwfnKIUCOkdywdCBMz4EHfDvClVo+2sG/dTRSgBb
4ISqCWfeG55groWeKiQ0eb9jzlUpgVICE6jVbUm47VMJp9mR00IbFudfCUMWwzgG
MK2BdnWc6u+JIPdqVpwVRUMtIT3v+D/i1VJyJ0KqeEfNWP6Lt6Ml13tz0rbCHoqY
FSG5ZEod1RF++xDEVgNbqYsD0NGA4ZnEkyloPlICm49FwV5gNxxDcnD+e9KEMR2f
RRRIul/p5wjqUPIUkS8wicDceNSJ+EHc0foetXmtZKCcjMgjmHm8yGDZh1ZrBLxe
ikHpKEir0O6Grt2zTUWvuHo3p6LhDBQjppPfmkgJE7+tcAW4TcaQGcU8yApGBQ7c
d7i0k9TrbHkoNG2dhWeOlU+w4RV1EOqPgeFPeGebOKYP0RGAElayKjBx5PxwzRjO
fAH88jPMCFfZ1wmRBD3J9sxZ1Pa8jnRQ5xkp8b1kzWMn/X3BwOMDUWZL9MNvpJqS
J0BfViFqUCuCE9NRhXozqQ7iv4dUS+B0tgY6Ux6OfNT1M3+s8ORwLfcw49S/O/3Z
xyZQ0mTkVCEP0RqZwm0EdYW/dLEsxbUCkXqBSL8H97LPPGTfkdJSNs/Gm7GyeIi9
Zcx/uUIxzN0pBD75Ld+DqN2uFNPOlWmxiZx2bn+8wcVqPT0V2H9HlDuLEEKluVeh
1gOQhefr+vXLntIwRTKv3eLGlYktBMyPFKdf7dfOrC5qL/uEhXdaW3wQYCEVDInk
fPgVtAeiynB2ymC+c8uuYCcvRYmyRKDXGtpKZqjgBdX4ZoYcPZIU0VQCgNxIfrqL
zMBNv9mKJBrw96iO1K77EUAblgyadDCBxTmHE4oEmhUOjUBeiuBWJREz7gETBomg
4RzW+kI157nlZsaFo8ibvnZX+ki7781/beBKX4XCsUeBW/jN6ns+lCQuItb2vSKc
Db9UzvkuoFMtABrl9FJ80CovEmB93sJsCiteIbCWUYD+mB7vGDs00ILOe+Y2ARSW
b68dVuIzL5oU1M3sODJVXGDPmBQ9zMDZ34DF/jKybDAwXopthSvy/BLjXl1IloSd
G3FzYMYlAKwrE4XlwGSzzNT3vbTi4hDXeSj+sB9k5y+Ai3SWcGe7QtBTGVgao97J
lMJXuexCstuztiQu4KFxXYrtVmHrebA+BIsdZpBOcTmPg6Ywq4abvnEocyAEjZJJ
7kf39OFna2+IPl274hkR554dNUngxV01BmTmHH2uaMZiU3bf2jdvOvywSr5bFuZz
q7upeJBgsviDWkcjTs7krqX2IiN+XCIVy2xgO0K2v6W3x9qwaz5A87wSHGUId/z3
4KuXzfKQ5uExZo3HvQ9YA9g0rd/AJTxaKc6OZ+DkQV9jbqRO6cxDZnjR77ZKuN2z
P68OC+tY91x3GXZEi9aEXBovF9DLBVZ63vpHSc00CgwSReNPP8EqeIj+qqFo/OTh
C/Q/BSnGIY7TqVjk11T3BvXEl2a45noxNnUg2Gm+7vo35edq4/LfAgsSuVWLSbqU
bFmmCpxlJW632Hpkv/Lcg0DYLCl0qkB2a5wA2NbrsLTfwGKc7k1Mx3RpHt8nPSGG
TV6LvUcok5e7c/vyUDRfZ84n9lYrsHMPNB7TSzLXBeQErTJrMTWuDmWFiRCyYRWE
sz/Pcnr6km6oi+C2w6kogTcv8YP9thuUg2brwKWJ63wkAWwJV1WTdaA2xSv/0BqY
RvFhFkgeGsV/6CJcMeChnUQQlQkDRMYh2j7Gf5eqUhjMRjKd6fRKLv4OuqRkLb5z
3azWGG6bKZlbwVAXZJsuh421IoLm0Ig8bFDZGWhQQMSWGehh8dSU/GiIJyC4D1/j
1d6+AgL8PdVjR7E1Gx6MEpUC9Da7pdaf85YFXg8X1/CWCSIKYfkjbK58gXLgcwdr
FdNsENeJi/bg6FHfyubM/cAweAuI9Dy02pjWDIiQ0w8Z8yaZ2o2O+d4VpKtjI2/O
EvskkWJ0FjUKs1nyHRnnquTVKD5uHnFn/NVcy3UBA5fpI6T5FQyxPukvhau6Nbwn
pl58TU67BH1X1KcQPwPlLXCdnMASNyVFvMW5E58P6yHHlNmvaGGkke6gl8SIGf5n
ILGpY1yQPGdOcQb+Vql3Vs1fp/mAbbzQvv0COY3gZxOsuCupvrJF5hITRUpvT2ya
guvJd+OpL72uoep15EPGNNW3bhuvj01FQS+xUgBdsNto4lqWh6GH07EieDdJ35IN
OmFjZyY3h2m5kLfnzOJNyFqGdlaLNPiYIBD9SMPbVVV6eorfgOMEkeSTGAWnGpTh
a3PfWaLPdu+FpJpqr2yJ+bD7Tpl9oLZO29zdQu3TG3r3lW82i3vWN5Av/nPzIggH
ICUuS203DQd/Kvj0Kcz9hJoDr8KGeLvA3mIqGMlyMFl0Z/2UnUZ6kUZcHz+2tZ5H
4DmWD4pJmJ2D0gPJNZ7t8n8KWqHCj+oQzegw85xRFFuxrWk8HdiKFps5mHosqyYE
+NSjw1asaY1dXSBQ9eojZ09iRPlHA+0Y6hWo0edQVwj7mDiDNfw1IF1ni6Gvm4NC
Ll/5Wek61FKeMiPJXBOSDNDUz7paCOq1x9zv0TRzqzlr7aZM4+SAM1DZjzGZAaQC
cp1Aogwxlbt/j7yMxQH4/vS2QrdTBPIbj/fisZc9mnIlttvBVwgr9Vo9LYvRWCPb
5HFRXgrCgNQK2SPFH67YDGc2MkLhPbDKIe+UjlWHEM+An3ZJqxHYnh0j29mkLinC
0BFk29WDRVM4rMtcFWedKi4xtMSrEB7f4JcX2hpIuAsSU5w1ZYcgG1eZNu/B6Uti
CqygNaAmqdlCZhPfz+sbXhCgtpvLaJV9luSup4MinPosJkEfazOVB5rD3qlhiesa
wqz5YD8MYxO7ElsZkGDYU39TahZesD6D4GaIQiETct8b0DmyyazReNTDzJ8o6NRP
07P3/Ruj0nL1H8NaCW9OhlYy98zD8Vy6hui2t4Rnxdiy1wTOAwpAuimn62Kc8TpB
AmRgDg5WgF4CeD1VPhXHmTrM78emWFD1ej7uSf1A7SJFuogoGkEWMc56bvnTnDca
kgho1Xgl+aiI+bQlF+i4hT7uv9f83C22eODloOGluUipXsAD6wlw7gDzL++Djvju
ERmSPfHghU6XSKF8SdzBCK035wlbxpL48CwUKUQx59q66Cm9ZQe+ji+Hkmjcu17H
D5aTwEVWdqEcdlzXqTkmufCsvmp0QXsvvd3TFXW04KomIZijuAQdWThM5oKcYCOs
aEBr2Wsb5gO4d6e5P/XSSjd5FdWKAuHglgHahRsvBIH5n8/yas4apEOxwkWVd+UL
+9fCkPCQPILJmN3ALoHEgrTt1FkpjoyOqovFMVv8oncyUoyZcxHBUSFzj43tFC1o
A0rJg5gN62gkkW0ZeYnEXunAGUxv7ERPs27dIJ5VF2WRs8+dO1fduDvr4v9lE80B
ILKShrerE2y8yhz7nUZlhNwh1T9RABvoFHENtjyt1yQqwKitYyta0WzhtRgtduZo
GnksEnkeXlxSuHNIPSR50aEBFjXQAqC5kHBzlF5BQP07mGlI/pVL1ilUoBpAOMuW
m7WzuTIrwzT2wjo7aszac0+zqtWxbRx/jZ4wzgA6Kx4ISDf5UOYBcLZubv1xzJeJ
DVDxKtbhnY6pFh3Dyk7jN0GEhFy5SIS45LdwLo1sJg+5oME1vNtNVlhr7zStryzY
yoew+7YQubIIuUSk1m3FhCgq8J9KdHhvSMUOTp8YV2FMws1lZqkVM9sNcS7vUykv
HExVBuwSaaxDKhoeU5DBPWPNhjs+gPyuKTC7/5yCRj0rb/IFWFxYIzC89IRjx87C
lSL/SQF8Gt+XMU1+03Mjv4/OfQhXgEb/eIMBefhjI17e4DanReeVPImKMrdWIx+/
kPA/iXYPHXuuZlHtmhTmuxdGcWZna0awr7TZyTnZpyQUMCRVl8o8nh9L3yAoV9tm
CS5cpea+u1JojwSdBS8RaNLulovAyQQDQ9SrW02Vvl9t2nr9+iYR5GFXDHswSsXX
lcd4PDBjiqyeaJXhweOt+uf1yY1XXDIJT+RVY3rzBekYovqDe7+wb+uKsr6jN3Ta
84l9tWBq1ffq4rNX5tR0m/ToAifk1WbS4/Qeiv5jjPw4/IWiQDXUC79GNJEpi6TV
3XthKvFOhCWI3d5+Xm0shKzsWm4L+BR6vyHmk9+zoFGIrcvqB0ZzzqFK6GkMQBho
vP0CF3FWw+Xa8HlKSSxBIKaN3phc11f3YByxa8j/XDDNsFwcQCZhqoMJXTc091yH
9hrre9gMogUAn+2Q8IM5ntaQcuEPa0hqdsxcSvZPXH39KdhICbrPi9suXhmKB91g
eQajyvz+IvR1ZV6BAjPrWghXthqLbkbYMViuxld3eA2RDXoZeo6QGvOJQ+uhRdjs
aFXKInpJGDfgMmhEGC3k1Yt0+H+LvcZ8Q1tdrV1Z2gdnuCCJxKPlYPsSL3U+OrRk
qj2+VRqzQMpXaTQ1aqTOOvAvh95wMHkEo37eJu52WfYITU15kST17l2MukTyyvhW
c6jzgWo/4CN5/oQFTJkZvSIAhGR0DHk9YjhRiXdiiQ3CcrHAu6O/lcLRRpnx0cKw
n5N33RXQ10861vFCKK/PKs2n7YEmRjZGKKBJnYF+Pangk/zB3H6a9UDZ3lBPBoX9
ds3XqKnkk9tyaUqsf6WztUuOzL4I/L98KW9zycpsCRyG2pAbsw2iOxOwUI0LfioB
SlPEPr6XIEASlFLZx8QfEZGJ3i03Mz30HRse4Hwuofr0TrJO+VvHdwQLdNDsZUJZ
4/4HRo4n0PSNuhDZD2GmrM1PSmdkFT9I5EjASq4+dya1FFewD01locn7D1k9fs6+
Ssaq9aSSeCoplPHmj1JpIjiH9GNA3VuhcJprazKChz3hftVuO0kH7ythl9/M2dsa
bK7W+2misin8yqk/WAlHLSd872f2A4FlSiElm9T13hfAmQ3Vg+f3DliHBYJdhCic
bmc/XUNApx5WwQUp/GPBmYrywJ1BOr5oFoD/cJNevHGtlH0pKEEERCHoQa19A29J
HFiLRJ3veNQS+aACtaQeNjZAVQBb3xR+jfA8x9ThtQdGDHn/6DcO9rwvufj5KfyR
/NTdCSHCyXwLnpiz5WpzF04VmALoe0XWO3WEKbRFlM9yERnlDyoFuPeFVTO04ckb
rWV8eJbUwhfIUUb+AFmtWHtz0/DYkqSDTFmrtZfO6rXZsQoGzDLETvIcQrPu8YCi
SjoDB+a6K32tTF2U7SJw+/WyciChGXnlrBzrgzUfNSLDxkPkKYS2+gA8PyJs3Fyb
loKWyvzRUxhpuVo69n/l3QfepA9dk+XD7UlfRUtOg+UAUTRhUCK+5YI4ReNS1j6w
ri1yUMmO8UYm3qZa9Mjwe/2cFcEyho+XZde4fEiHw8HJ03tFDIt2eDEv8ksl/PpS
GL13szZVMplu+gnYmaL7H/ERjJ0YPbmTj8PYITCUGhqs2UEM5wNjs5jp9PxKMZvH
PrIQ6aT6ZJIS4G7xSJNgjaGZuXOMd9Cs7CSITJv/HE0c5bnKASoVB6YKp+NX1ezj
mURHRcdGDN+qpTqVstJzkOP3ueyOkaeoc+DncuhMSKqh4oLnsbbsjwdq0NmI6ZB+
9JVxnhifNnJ1jGhTcyji+5baiXxLVYfh9YkEWWp07cxAUPJVjU+VAbKbM0raH2zN
lR3jTKUhb7MuQgvrGcfiht7b7XIDOej9ByFT/R+bbUgqmwBF3JhoiBwXnt8c6sC6
cFsjcbyI+c3Asm5HkeFyeti49hurkSEsRhAMpsvFpnStgeBVWhmcRhdj3p0PyF1L
F/1LdeEn8Eue0o0YeRcT5GYncwLBqon7bEQsy0SdHcCoMrFynYRxOcKwRCYoXPv/
CT1gG62YTqB+RCAscQrsDA2i1pyFL5zy0K64SIWIE/bXCeaOC9NazY3brYb2lzP7
usmHPmceQ/Gl6vkbuynQcPFFYjwtMujHEXhg+1LV3scX6GJqBwmOD20xEds8FD9M
CwJLwe0/cwmFrIDop8358X4AKXJZO8tEyWGNw93ZMXkCC+IA4irMBIS7TjvrjAZT
6j/CQzq+XW51UavbCd7DJz3jkWWAXNsAuCO4aU2pNfj+PN0VRk6kUe+ldOqGse8v
VVQBpy23iF5mrk8Kjj31pYJy6LrKta3s9CZaEXhVi62AcOa3uTvbE1nDThCy3XQX
LmDIyhjdqgfkngIVsCgj63C+IPy08f+DlpAUkbZ+izBKzvk59aoPcUsRsgDBfj4L
lT9nALv2eNs2v9mVv/7A/19/6BEfpwiWsemzarxx5CoMHP0nUsh/EC5aGtQSa53M
0dp7Hgfv3BWhGpezcoMvmrP5BVRYkmglhB/U6aXQWKf6ap1rQY0hBq6HuU6b9faz
ld1DqfFMt0DN4PdKTfyb1nDHUUgF+a3V3hvZcKEsSdUA38O/Xr8XezJpYjZPhzdn
Hot9/LybWFlVMon7b+bafU0Lg4RsAPkhiUaMYVImz400BQWXwrdhQsmZzwp7PFq3
lT87G/Ei62S7kovrndEw2i14Ol43r+USlRwljLVEAEFK9+0cT85WAlbduOhtIRpz
l+9O9o6kj09t6RYZQPxqx5Rb+v2H/yu1TbpgB8ekasfjonWEPr8WLaKA6xp/xymS
LCUglNgKrBWzkiZeh29xm0o/agC7L8uEJ2v4eMDXm7CCccs6BfAJ439YaxKNkXhb
OCHpHpBQUWy+ntHhM16Gr3zTzE2S2g0uCKRX8TLBGQRXzBm/CaeTgCQdPFje1u14
kDTPKm3lFTHh9t9uxJCiV/Kxq4McVSfERaDQ+F+4j2aKfmYh1vhYZgfTcGH8Bkzb
R3PSztejl67bH+NJvLjwMar44CVO3l9EDIwMbdwuMZYYW1jTRQviblqzvm9Y6J9T
KDOVjDKwFo95zJrq8+bdcSbKm2eSbjDP6jLnXWlBXe1/VRxJVZV99JqYYu6HNOh9
6rJpIGtFglnT2ug2pNMD+mt49cirC95I3H3iYN7ePNoA5XC9VhbCFSdMzTWY9naA
BCqqduiFlYydasZ4anBm7yjZ25UL+FM1lNioJCffbQ3iFhHXsH3N0/p57/okbYf3
sCpijTPEfp0enTKAiVahuZCtwf9GEjrhSQWasW8ghzo2yWRZ89SMu8XNhAQeuv3q
lNmbGrqUpY2ueUV+YAFWcK4aaH/8VJi966nuZQwSOBWcC59ZaE0YJzYsVqjS2R+2
H9LR4iYJp1fwc8+WoKMwEx5q3rWvNasiObcn49JnCDFWUI0DSd7fVzXGFd5SjTLs
QCI3QbNzuS4/MR+kd0Vg3plEIDg9dSaGKU0d+P4ETyNMi1Fu7h7LmOTF7i+KywHf
fOjXrvRtyxxgWSB9eK8WwhOlAbw7Hw+yW0QbdFJ8GrrmYV2nT0RgS/0vU/aK7+rX
lbr34q1fvDO9VxIekbP+usFxMgTuHfctDgtzYxUgx8a2qUuqTxlNpaHXN/8wYmDf
36ZS3NbdsjPXLMqpndXY+2cAMCz5s7zaLt9Q3UGi7eXakAxK30qj3Uk9MNP7GMou
bAlCZk1J8T0Nwgc2Fo7n4+k2fnqT6fPZZfpuPd+ZYoMzFCOg/OVDfVUwZUW/N0F/
Bs2SdW0rqgReXCEkvOIstBcAYXpbHj8Iq1DWHNFUM1qLisVa4T8lSAo7YEx2jmBJ
/RVBowJecG/QC14WV8WgaHoPF5XzqaHKiJDFZn/IPtFRRY4XRoPxBi992b99bitL
a8vSFH98UelUBmklHino++KI8LNh920KgCwODObVQzlqveN0/1t3ggKT7s2JLxaY
K8YUKM7T+e5WOxe/afN3DDw4RZ3mWpWfQTGYMHhNpcvZjp28FYViIEwNgjdwpXnh
eZaPSLdyp1wuvZAqp1AiIFf8vewKZ5QCwfqJ6hY4+Le6tRmlDqF9f0j/ePtJkIrc
LRrD2+2iPTPq6pkWKfY5nCEORBB04iqa+3ewda2KxXt9zUrnmAiMiALBdB+gb0C9
Y7M8lqPwxHYKLff/ABSWThBovpZ164HkxN00EJEGlHBoiSHISB0gYTN8Rg5fIpoK
NyFI8mjr9T19Ce812xHBVygyZmIvZl7xkyvKfwbVf+MhniMFsx3FSue1w1eyui+/
QEE+WFlW+pRs3p7g1YBftLdRIlEAoAWRYnzhOTmsKREasX0cHS3o8xKtt1RwgDhU
PlukkmZmN6JkOm533AvVOAgT+oEEHmlE/qArSd4aPr+sSMTnepYCvSTO7QF+fPPi
qRu41xHkjwMI7AWHVdsvoI2WszXcYtFzttaMNWMpIQwcKYZx50qMqY0pCQA4k/Ts
fE+h6WiHjZewjQvhajhkP1t0pLP8/qPmnpSKHTTBI8+Q9N8Fba6dZqqDy76XjlCY
Ss1yWOW0+v04eX+91rzN+X3OX5J47nDnmiFvvLOx1JyQsxryoSqk2zrW01Qxfedf
1t4BpWaghd4Nw61KnZSa6QFU4Ef5xFHu1mM0ESPP1G0qmu53wCkcV+TGLzEmNF3U
WBrvsuLVk1Hkspt4hSI4Ibotx1u2BOwwin806XjTtOeS7DRcl/FdCHChp6eMlDUW
VLJeIXk75JFiL5aqPsagOEp3d4k5656Kgbm2kfusq1VGLNZxLkoe4YJ5PhtCFq+x
kLHdf5lAGW8j1jFJXr8TXyvUEfq6V4w9UPd7tBXCb2E8Odjk5laklQW9ytVjsqz5
rQlbKtxougP7FBud4jxpBGkSt9G2WtTs5UHIfMHOiw/hRfo+cjTL9Exila8llbEU
qjRNw+OZaC6217rvmM0QVzof1xN3Dhx3o6TwMLFJkeAtglhi0jZb3J5UKekHWrCd
RTLBNeaLq+Zu8vs0B7JGPrTeFklg4n+Mwb+//SpFk6KlqaH8u45Aqj+il+q2vIce
BlE1xI7jVV+wC2Q6qUNPvl7GWSvHhptRoMjkjrXCDv40wcJxRpeJgY4OdAtefpFd
1dwzU14N71mAb7JlWQm8Vl608JLe/sj0ReE7N6bPMUBFa1NJEQxWHZimnwnJ9r72
bEE3yzdQbx6BXzILw9Nn/IUoNYxg+h4i0DI84N3IyTfl6qJ/09xatbUpSO5aLLf4
KeIllxXtYxsote5FmKTUFZnj+Ipy9wREr+TKW0k72lGABKkmk15rmNlIBB7qqdy/
FlmFYhNGt/eu6Ic7yiY6QX21FgHazC7qGgdvi3iUY+AmDyv97gUZH5dZ5ZsSK41C
zs2aE+6rWemFj/pngbYRZSu+9ZMP/fQLG1k6oewI2jYr2i//Bd3D4yesrUiZRk2l
Feb858Vn8dbXC0EBMWoi/lJCZh9p5TiKNQ/qSa12N8kPzIIXTNKLtvfBO9Z6lvib
xccKOn5JYIpxGUge6igTbfC5tzfLazNMogi9Vjt8mEVqpjkK1F0NZSDGgF95ILha
wupnuwI1X2tNVO6x3VKphrmqPpZCJi4mx4GcGM3LzTOIhHjb+3Dbn2KHUsXKI9aq
4BkTd+Q3iti0geVDV9QoZ59vhrTxgyyMcf6pH11cGmeobKpjR/lEPyRmh2l4h8b2
ExSVNwx2SPx1MNh18WPT1hFJoHNEiayQgRjqwvJGJK0wOg52GNzv4vLPHLcKLsNH
tJ4Nm+zeloT9VzgpRzs38oGvMyhfPS9wHK8cxUlUCd4XzfOGL5G1zaA6LWJCKe1W
2MzA8od/vS8+CoJP3+daGt/wweM1yJpw0Tb3B1/XKagTSkIXkF6RzA/hHwE261Py
0IC3qgBjGklEzKEdQ6fREKUvJNiUZEgMY3InfcabX+UgBZN0fCHyypSdmtnFllVo
7o6DFMHNlJeewQnOT9X6IbK+2V7XErDMq2M8vbSWUSVNnWGfan96TxNnw1CNGaLe
jp2iYnzhFDH22xeI8tjeRDMyrNvCexSmwBdwbFPMv6uAZmboWox8grwmfkSQh/cq
N1ve3v5D4NAOo0rny4b3gnfJsMmn7O7IOK2z/fzpEmZaF/K5f8kfBNihxhfMtpnx
JbcG9g5Viw2f9AniXkVcfMJvJJ7fcqunDfaZFyyOSAIxMdpgHo5NTT7qdUIwXClJ
nSoQGJz6IFjxi3qTS9aNm1UFiAKslgwivF87KzDMgJG5IqYD4hTmkMXOOBig/WVy
Urv8P6kKB31lkuJ8o7ZYt/lQPvKoTQ/tNC4JoSpEQZFkxeb6T18ZwoCiv1r9lLNQ
bt2Lnd5D0Q2BTVGpudWnv5gFNEeEQm6Ye5Nn2eiVAqv08wqJLzVraWMPUgzKI2iM
bxJb7YOOqqhaeT5dBkg4yHZirs4O7stKlN6Xz2l4lDf72iq2jmNkf7nJSntPwRVi
e4Kul9JD/CAWLRCY/UtAOBYsnr+ajrWVXmTLGMpnnR4+z1T9nm/f2ZR0BGrBPO9L
bgGbrpJDuHfjEslTRRfMYTvScZbAjmI10FBbSMEj9qZ6knXn9D5EyPZlQbdZH3us
CcoQOqRFbJfqHDXdLLoPns/M6bzkXrLUskMA03irW4Se8oRmuEugj2kyHeFGryYL
WxPPu+8CKcHcusxe7ElkNo4Mc6omwW5mJuY2ftINi452O3ATTrsGqLhXlRR7pK9n
hbkT/Pj7LB7vcHb8ZA1SE9fHc+eR/wRSQah+NlCs9O3Ujq49BgOxbn6Oiy1PjtT2
iQssaj3aXJ84MojfdyTdv4iOayRi1nbuPDbvX0CK3TbHiPq5GXoQJAqrBGSpXzJO
gi2ywyzhrcMGDN3MgAxLbvFXCsFylXp3B0z9aNxd9DKLN8WmuUs/WDfC8sUOSF/i
G9V66O/MixwsWtV6pyLNWDN4j6gSSpJ5KHyOfbrHSDtuAJU6VuM4i7Yuvolt8qV5
mTDKK9yQAuLdUu5ozp6QBLBd/iydKhiqa4LhFz/2ZG0UMOXPCnM37QODizQxa0B3
PETXBruS67kWkCxAlGAywQpW/Qdfcm9mEDajLMNJ7jaXFiTx9OWMMLFv/CaoVoYH
LWkNAYJSWQ7F3IDXNYFnyrQkif/fTSPHZu81USnEtyhckvwGSRi/VeeGJ1fo8FOd
MSkORIxbblZWtevOBsoddbcpjUbpoXOi321aqWz9FtAkCPM4ZijoGLiN9VWJtDce
m01EvYmm1NkL/ZISHGwnpbiD66wM6PAges6xStaS8DY5qUhiDHQi2tM3wDu6XnQP
qWEY2QbByqg9gUTkjqiSc0inD9VQG95HqULCTpw9MubIqxirazw2RZOoNGmPU6O9
K8vjnj3NnNQ5igRDHoqJ0G4Mi6HhXYTmkkuHPzVeXHncLPUWl2n1jJmRq793s9Ow
TsQQanMO5R4UY4hsddZ0nRRTMhhi928SxoX0deDDiET27N2z8D1jF5QDP2GLC5US
EgilCos2Ws9DrYYSkpWnI+AsZevATnJSC/jyqJanqtUrPpkbtVcO6LAx0uMTFswM
vs+BpJ94dFX9tbwYMiCuAteMzhk5jOis4Tzx0m2nyT3YVCaOShvt2i3/X3LBRUlf
XthxQcnnCH1ziaTY/K0Hu0ilskcUhi2Rs07J7uRFGf6bIglr94S4ZeQDRsDD66vJ
GsPCDpWOrDG+Pg8Q8ETOSpPrzX124Wv18wFPrDVXtlLK5skSNG5dVJkNosfEhpGr
QOby0FLjMSEzOlCD9TDr4cHpoDLOz6S2ytFX/3r4NNqwiAmR0us8Uqc/yciGnrjt
MBcic8rpZbsEvPLjqxmsEiE51D5zc2UnTHWVe5ddw2Fwtk2pKowgvYGD74VuaT6y
M1Rg0S9XEi+/bVMCvx9q+opgQzDMM27EhI7D6Xwxy2wMOOMjVVZA5kEjROYLMlk0
7OaIv/KBNN5xmW2jUr+xzfioJ8lDvbUaCcjp/nWA2bAJLdAOj1cB2YxhbPXu+Dcr
wDuFmu1mH6o5v6UenudCkJ+GhSPfp86f37fxYuETx96I+xQB/kQhAwoUFM1SVhGl
fXTXOz0GvdzKaP+VT/qqjIx4QeZCUyzrE+TsKFtsWzl9nRCrMTyu6FP/QbjA+mkO
4d0Uab2Ra0gk0Mb6PSf/990mRIXlNAzqrglerTVmUaik6dm93q5lhiwcMd000/wf
c/Q72yaTIkEzlu9KZzkg7CDh4INSywt58BjRa9gnVHu2BLY5Yn8kQZezby77kzI6
1JrkzCiPBFBufdGc2JIERbMk3N1FueELCMMjc66fOl7EmvYuRVcpjvs6EUtoeScZ
CRnX/bW2uuSDSIN6Xa0HeET/9UfkdglijETEu5pOxisNvrJrlNF/iApWgeUQ+mdV
z5Kq19SXU5PP2nRgSfHF1vaiY5x8fFuAZ3lcdQ8gAuZYFQH3lZx4c+XbxVMU+QV3
saH6NwG8jCgA9ktZdRDKOxfzovOJOBxzqYt369WP/+VfyrWmMj0+j+khwyPny27q
I83a3lpJvgvSC97G/x/aNkQDzkQ+GnVtwOT1jXO0SSCRxItruqg641KWM6jhcvV7
zQX8jgQI8/2ZWeAWHMJR3tO22ThKK7EW/9KLgH+EtTwKcQGSki3RKjPltDubzA36
iPgFN8vcjBQIrDf9DadifY5i5u1lip6ZolvYRIXwkJb6jNVMwEQx7khgeJx5178v
vKRJSZ7bU29suafuxBJKvuPqRLt5bbJ4pakF0bIVqN9fsvqwJdPt0t+cqAGvzjwH
0rPd2rTpOHn/z8eArqgAIxnegQvV1NaR7wTPnFCCOq58HQ0/NwP45VvViJukYhs4
wJRcBkXLvlr4moVn8ufcpp0MIEpDfNv29N6pu4eHCCeW/F1GP13wJuzvELU1y4jw
jslKgUfxc2Ur5bPkGEI8jfCBfRIDxiOSQysdM7ML97BrEgr4FSRqJFgbP/wLMvb2
Z8H3xxWz5I2czcOj9d5GEjW1J4gk2sXLOeT+6rGW5wsUM/ev0aec5Moqh4UGx8dl
uAbLooBssEmxh+hPXnz6LoJk+H5GdoEOxEu7jNVJi/HVer7a/vd3b1Xct1xGUUAK
iGYjcjUVwLGzj34G9Sm9+OawZL0D6vZn1ogPMVYeZrPC/Rtm4hvqOAXgSCMCMHaF
jY/pOSliEScmbIG3h+LDHeJMmMEIphIsaCtx2hjQm7h5jGeTN/hO1INLNUPPTE6x
+RQzF6xwL+PJnQ0OYtWTmas09ouF2UJdLY7W8nquPUliBXX/C1Nxp5bce1fBeTzA
/Y5ZGKujhQV0XAz2GHHNgKgP9bcfKmfY9ktE4VLfUJKu40c+fhOvsRRw1SJnZEzt
S4DqdbFqagcbdO7sLnqMLjVfgA/qAW/dn2QoM6kL3rcxwlrzk6Y1QUakad2GXXuj
u1kTodw5CU9+x6mvn18/rwCvbSryNHgE7pUPjfhq4YbKPUiw1MAzHQ50zvDc1bkm
g1mWynT5RwWRTmlM65gIFYUK5vQxUuOIySsaUels5WsID0hzTv4oTV+nTOWp3z2M
P72x/D2W76PuqqA0shUq02I/yLHHoWdPmqCGUBzO/VxNUwTB2H0rKl19JnP0n9xY
dSpmnfodba6cxScocJmtUApHbZI3ExkFK1QMaPpyOucVW7u2tbztn62TZjzE7ojy
SaV4pEQcT2ihX9RzFnJp0BmVCxzGukw3XL/jYFracI2NAa6NUTRgEPYT6BlwKqkS
2wYGJk+flDm+IKajEPRo5JVkAoYmyZvXw9yz5eGWlKDMU/z9gEm0R6pBu3F2ZZ9K
KmNSChK0n+5HPilZbiJ9nsyFMevIqOXFVKsi11HrMqy1Jm2yX8KAp+xXhP767X8q
OaMCT07S9Ck15sQoHG5lqXW950I/k6PDSziiv/TK+d1ssNaN7wXQJ+qIHZ+u5pVc
0fyBu/R93fP4OFGHCmnNSPN4Ut0wxXc9+4vPyQWGKVQh/tvS6S8UG3xcECMX5ygX
3F6WTSwBipYiEbIMbO6GloGORoTJNdQAgSkVbehNfvKpdGZmksoXFzBZTjLXHfSG
UQAKfSZRL38IDzxaIHSDPOUWi9wZ9C2CZ56tpnP0zohaKfh1WXTbSRA1+wClCWOl
w7ikGx3imedZtDnhkrDeLAZ2DoY/Enmk0rhOTZO/TC6FHUFaRHhFMi/nz6K98bX2
5wZwhAQBtCVyipl9TF594FOIA1zwiGqipMtt7Dr3ajos+6NkXnhwRFAyq+6+IpPM
39aEwwmiyFiYE6Tor8cYnxk15kKi4C76NEMSITJtjvgVONTU/F5wS6GO006Tgrrj
Kil/mb1mnBLVlUX3h6CMLjESASFffnsjXoc/QlI8uns3oYS+AizwENm4KOQn0w47
KSFRaFTVUsZGm0XU4DVAaKmXjuS6ecI5SS4wnM7EcsSYaqsvF65LIoPGHP9KKBmY
6CQg03wzaT5AXE33R1F+6DHlQh9OnRPyi0dZRfg74/gvEbmfyF2zNx0ym/ggLObA
GxA8dLeciClEWmC12Sm7BFSQEqWrqL0vBN47N0PN+5kmmXUjkAmSpYf5P6gDkxeW
xzZRMbHo1fBpFiztYYccvQT9QAv3iH/ZwtVwxc5ofwBT7GfAXNmdGjvsb6enyl46
TGPgc1qgfm5rnER0S7wf+7C+Nqo0uR/f3VVK5MlnIJwtygI3jKSCcedUyTkV46ai
vmZ9spOjXGmYrismCK4f3LxPIKC6xZ5l+bXWnxt/+vdZFU95HequcitufO8Rhd4T
NRsYXdzj6rVV3gPG50MHwmWSeNjXiMD1m8xDITDpsfdNqIkQ3qVn1/LhxKfivTCD
/P+V7tsRfmYMHX8M4e4LGw8TDsIHbFfvpUp00MQBUu4NYhjOmsV1AXR2vK+4c7jk
rEbJ4fcbFu04M3YNLOuGaW/fvkpL1f14z2nBxlOnxcx+GNyp9ichQpCclB2APV1Q
e0SgeHKqnJjzcGgdkKB2hVtsM5OupgK+yUON5vcR1IRyn+OJetaQt3R+BlVAtCE9
C6a3DT4RlKWdSGahd9zdim03GixC1ubAAuXZiUCa6a+AXl44EgiBnvHr5MQ7xbe7
49DMIvqCqN1iO96ONSrnYVHexMc3RcJblY+686wlEp/1FVjUsyBsPbsBx1suRyQV
yoQQq8YkhR0NL9dDPCJxxnLVlAgHs67WxsIXQ0szSi9kJU1vjgV+KSXr8ZMk1/xP
z0UCs4ngjcEKlCUE0Bkwmg7Q3mwZfh5PY849MLrzkGrxyZsuTdv1+4UBqr7fN9JW
ECKUfYU8zk5umecIMxqFi0XH+I3M3zCHjMqt22RgqVdI24UZqlFSs44pSHBtXYrr
afmjpPNIkGIScRGmybNnuv+VFuklW4O88kmMKNs1GGAAUnw+gsfc1Nf2VUKatpwy
Oq0ino29rOdYNR+qNDSec5XVDl63B0UDj94Opnq/zzzvEo4CohaDfKhUT3PAWlKn
70Y7k4b1gBzDKBSgxpBSi6fXsW3eryN6sck/UKx/Vp42qlFsmUHtIq+7y0pIx+fe
G9bgxNAoKFNc3L5k2NzeqdzZP0xlQL80lbM91pOU2DJhiIAKwaY397mB3ge8IDgL
wn6xHLgOsUfzj9mqz/vLnnXxAnCKpUqwVFt0f5nPTGfdw3doF/25T5+d8CjTefaa
K/dGtbcww5gcpG4U7EOZHjo3m/uPR2m0lCk8XHOJ9F0fe+uscTRzQ4m5wGkP/kx8
1eyBnOWeorIlex1FyCORil0XdnnEOhMipDCTl01o+R3CQbLItKhExOUWS2Ru1eBi
PaXixtuSwn1kCR/4z+ishah6ZmCfBgdq3cnFNs5HMR4CDAJ+Fwgt30Uqxfmq5q3I
WgLrNk7Cxwxs6m3T9jrOrw4FNificPNe15DuHks5olOUD1glwcbkLDiykEiX3h1g
cRrDrRB+Oh1vLmHMIdMQ80DghELcBar6ws/cXkgudu5+e95kHtxC5w9P0y16NG4Z
NpX1vXY05ANfAQQDSEis66TTmFn6bWujY75IVBC6CoY2n0pLJz7tQ3S/fQCPc0F7
BbFfomYf+SPLj9265Mp7Xj8tcV9uDhKaxjAx3cYjOIvevhm10SZ+VvoKSkOKvlSb
1QWQHob1c9Gzbwoz1INtesJGXfrHWxWUCz69s91KKVKZzQfV6C8py5WVww4NioT/
gZ/q0MWzBhyfCLdXSpZgY/EybwO35LZpkfNnfSR9p0KCYGSBAKBrM1SAwg8SJYVJ
4o6dh9C8g7qM3u9rmNx38AVeKbqoXuDAqjy/qrQypaA42FvdkxwFFskKTMguuLYJ
hs/g4O/C+ruk04A1HfeOIjH6HCItVugizZYUnjVupDg94Y7Ue/wd4SXTlID2F3DK
2nw6QzQhwgncLdzAb9fIJXtEOmzmYX3BdKhxKVg69d/pa7VUtNs0khjnIu9FIKK6
vUWVapErvjQ6kItsH791J6l1k5Iy8yv06YaN8MMFBe76XFRyqh1YbvOh1Ea1GthS
1BoksWFq6/NhMhMywEb4Ch4AwSzufn5MkV/G4N/hAZHdITK8E5uThJsbz1aKR6Jz
taraWMup631R+YYfumvsJ3/EPK6Kkv4+n8Y9YFmcMbs/8mOZAj/kmoQ8/wsEn1T5
z6Lj4bHxLiED6p68AECALpmK4E655G4EbVOSW2WkHZsbozZ7wPKpO0t+I2PzcAcp
0LBkzu87kg0Qf5n8tN3qoeBKvxrC9T0kbW2ixlDC6rZK4W2iKV0BYUXnB4xNApUk
3oUtSz4FGsTvyczUL0OxhY8FTbM4oiK7HrShce5LveUe4QOnzcRtd4vKfQXrwwlq
dk/INKKa53RQQgviQOAUhicvdus64NNws/KA12W/7P1bU1gdFhp4J1cCsjIbPsqq
6TL4FVQabFN6sGq/KWQRt9zQnBE0wzH74ZV9HwxVH4iWbixyGZlKyMj3eYmmM8PQ
/d5KvLPCMU3yh9xSA0mYlLFfkUIwxz5MYaQY4EDjsYNeoKTWXCTtvbewVRWIcyoT
ZTFPSc9bNYtDEgxC7nG/H3/h57mQXVgMkzoasaOAbyVW336M1n4xQPebet5IUIC5
P1e21+ci1mbQKQPYOgDIfuU1rBjsHDPujB7ysfYg6YdjIsjDgR3SqTCVswBixbe4
bq6fSnRcsJnogaFwd25pp6nbFNTsJUAZr9F6/eYOBwbW128wuDauzUT1/dNxsjsZ
PiIL48EayJTHM8APPjpLX2kBttjkEr/7S3ykf6yBvBHPwR1lAHc3ky6NKvioNkCX
fwVQoEKBuWd5S8IWsMkKKkTxByqeq+KZ0D3VGiynN6tkIb7er+Ie2TWDLOXi2dX/
c2U66l/NMfdG5jvpHDPPfQoKWDnJwvpKlYCqsdgqvcmzROBq3cJQuupI6vymxQn8
95KtvSRtbwX193OVzwGjZ/ibM3r1P7Fft8NUeOm8/Whkw/B6QA3w6HXvzieYsDVn
NDOpW9YfG8mnB0BmHzqQYieeFCDeYmQ8Yrys02dY8JMJgNYS7hic885P1nJkczYt
vv9oS7nQbYQWhgc/8oEQ/jUJLvtPKIcNJZvuJY/0REYPtZ7pz7YRDGYGX9BE4nRQ
15RxqAZJqhdoVyrh2Tvh4brHCcrn5INEe1wWzrGm4JpYjkTsPuJwZ5xai8dhku7R
u+5fX5h4IiYki4E7BbkdLCYMZjlIHFxr1kIG/Vv7kf/wjZQfivgcKCyv13GztuED
TVqQIL03ydBke2Uq0M92HQMMIa/G9kRsa0+wkbhk4sq+XPIfsKh+pN9SbR/IEei1
qIPGSgPyqckipE5kAgO+GJpRt1dGHLG2254YJ1q1eTcCfN10hqZCoCeBlWT35XPb
L4/VXi/nwRwkJQGonxEYx0neF4TlXStC3UcHui42oqRf8zNaPZhOGQEjPEwpGWnx
AiUMluvv8sKXJwfo01g7Eg82perMOquvfRMwm0aLhyxCwXQ8FXYinACZuR0yg7WT
dROvxs3GpoYo14ElBbbD0HFIx7SnCA84pwPcL4yNM9HjbrDK2I92yKpzYv9AgoVO
syvf78AxqOzzH6vimLf0VY+ilH5b4XmJPdz1noRZNQ9ttj0ub6WsO7UfJd3e8Vjz
iYgpWVf2VMlkY47G103sEtLiTkwksyVQ8azYUND2A0OC2jfA4n3pA1fFu5UGEHvU
XpVRAXxGYWUg0L8MzRoIThk6gK79DSncF/CyV+Sd+JLfSlj7l2fbm8itF3rE2RzN
ubbAV6bieQB5zo/0fSAzaL4WfZfKSEl0QysAIgiXBOjUYkbDyyd+8sH2zlkeujp5
dLo/D4OBTAgHDXV3mt76BBKwSFJ0Aylpw1zELQvYn3c5jgAh7QXCjLSIcwDcAV2z
rrShFmIyK1e4ex1lInjuabImxbnjWBAtzxBO3t+hzM5UklRrRKRmbVCEipPkEr68
VE5KQ2X8V0RryPbJv61jbEa+DRvx+SKtflIrmFBAzWcOI2fdE4YJKb6mv0QZXtD1
z83JBZlrhxedOJYV+tiobdGGon+vjyS22Iw/uFNQTCjQrJN9UJbExkCrxtrmArEh
ihjDM3b9YtVSGsIaPgShlB2DRcVHiCQvUqvuFrnIYuYQFEEJc9+yOFCYYIZQ5VDG
WYxRHyKSbcBd0ZIH0e64dJKPpGfi8xRkPIr1r9nQB03NXVhwUUzRJSk1P3cSwM0d
12Mjpj3j3CG2FfqOyaPb53bKTL665f+68RLzRQgqUj5qcanoiaAiA7ZqAtDAWwlF
Wp+cUqMB6xw0kZEMltOPE91zLv/b7OTqeToBChhIjzyf++7VUNzMx8mrKYOllGML
428+13cXoFUoovP11wkXPojGjslnm07kcaMBJ47Zf3FJIbuznQyQPhsfeSm947iv
+0OH97Xm7Q7cR9P+6jDIxXkN3IB9JLHx7JnIsnUTqZhs+z0bWlijz0RKDMMsT07/
73Qf1Je6S0X4fJR6M6eerWMH+MY3WLG1bWzsZGF1vJaHr/QJ/1SrMvL0cu+Y6H/l
9uEH1BEz1XGB73hXzu+qN46mhFTKc+htV0+NjnKyNHqsryGGi4VOQ/zZVQbs3sSR
/ogDasXMPpnOCtU8tY0Jh8/ze+caadxYtRD+ZibSyXPV5MZLNHdkw3x2P+N+R1XV
lV+67rLpgXxWFyjsE8TbyFmnK3lSbQqu5yxeZNxyBZd3HXIaGxx4YT1LSE0p7Ccv
iTD+9OVDxhwIgpnaAIjG/8gHyWKefUifJflkB+4RxAHQ7AVgcNavuabMnigckdqJ
RFceqKUyugIXMVL1C7U9RsND8TMkQxGktppLMLy/Ve+xiJikn61UNZ86BH8DE7GI
VieuQ35qUkAVrwrKOBYX0RMA74F9hWKb7rR8V48+Lk6atYNxiZQhVtEccyTE6X+u
2I1hHQ6nrRRhvBLyWj44HjKmpX1DcVSkViMgzOPUNnwaxGmzB/m8ueETpxgVuzTn
WN3/eNZap+Uyi95rQJkI8hoOL8keck1amuhK0VO/7IbkvLVhthca42EoAd8Q4oz/
UhYiICWuVN1CFT8peGXYL6lXU+//fSUy+M/JJCUbIg76eltAsgQisgxs6rw4M8La
mkcFkXd3XQKVM3u5saesp1Vp7AODGX7A7blNUB3Eal8U+o8rqfxMD5Z0aUVRegkr
uHddmnW21CEB5kdkI/HZCgc/IhDsPhpqz/zbqq/RlmFr8hj3z2ln+RdsCQ1HWGpG
50hly+CV19wHv7YpwGLhYcPCctag2oO6FnpTNDDBTKfLBCIJvdfW6WVjaAj1wrrF
wKckVwRF2UZIk1KrucL4KKDqq+jzoCaqBJf2sWvvWHrY9FqSszoX/mLw/8jh2793
fhSNJjYvsDHzEkDThH++Iyp1Jt8VENDbaLEz5gBeeAMEEIuC/NWeULfqw4BmaJdP
m0H0XMhd3TAbjvrj5eCTnq86P9JWqGn52F7MlyfG7GOgFPi/ytGLm85MvIPaUpxZ
eBvset/oHCCoHDrcPIKHnUX8wE4ITE2MK23cTVJ1VL+wR7AtQCCNToyq6LcxaY/F
Br2cy/LspK6ZIrYvydt6kmn/o/Zq5lOmRDrz0KdRiUa9/8YoqS2lz0K6FQx4By+M
cGbMRskd/G9aA3TZ+tbnNLqzJB0jV4YrUZnD/ChdwiJXtrxoHu6wF4dsCNKMdk8+
lHisj39oUxCtr/tsMgIG88Jca0whnvWuiqkIbyGdCSi8ghgCtiXgvwNW2k5vn0Gu
vUqyiLCSehqCS/WtE14mj/7GVuQGlHJODU3vOwDqQD6bNSzIDHfwiz9UR+GhkifJ
wc5Z37+p3BRkws9DTd6j3VK/IoMnjtpSisU8i9NP2EiQimaOdV7F2bSxur2xdY7f
6vhM7CRtdYOVCBv9pLfYQl9qguL1fcyeM7hBIC1lUpIno2J+A5zDtJucoDbHHcQi
e0jNVoF4Yp3X1pVSsn1aKsyBMqizMzPX9Z70NvQUIO2KrRx6ioYX6VPA/v/bIf3A
uoy2nHpbG4yOKYUHYhqTY5CnvP+Jihbdl/vDfuX7REue/CfZF1HHXHX4jGm+xDsa
UwE5As84PxK4xYWpt36k6jKaKxuw+xSvLhNb3MVUjFE+Tvyngh6S5XbqCPKAqObe
TD8RccR2wJ/dbmq33XLDEvZ+Z74L3Bekw3bzvHqzCWdUUYW3xwfeiQijL3WNoQ9P
0mxmemldLWXUwvpmVaVaPRanogZTTw1kXA9u86Npa1lfeDsoyoylwUaWU2ghOKCd
EpLDvEG8zARbRIbng2qFDz30kMP3DdDgskWG4PxcpMoDqmLix5bsNGOxfAY35LQe
cPV+dUqZoVEEjKo8/MTdJYboNzBeRBmSe1cXNdRlNJf7p/PpbtPqNVf2XXDt4yWr
bWr9C7pIfy1S5aYYw3JB4FLRHmgC0XucVgrB/+7qrGikCFsYJmZHc5LpNoe21QY/
TAdYgq/inlTa8cAGNCabrkvrtzq2DcR6Pq/nags1oU9LKXHvegSscwaPw+iGxpi0
hdrfxsECi6UyAY799TTKyjQ3Jhs3fyg8YkyQQdiNNrPDjGEA0yJjqrlJ2cIr/00x
NDUu6C9aBYjWUSK9Bah4H9qlwMLVdQ7bHInTY5BLkGY+UZO4YoK/fzFArfxapX0g
KljSsL3sn2Ro5l4APGhvkWVfDMYR63LWIfZ52YCItb4yUWaNSBXcxThwi3a5/O7o
ZARi7mNXSm6tEpFefZ0RzWB0iZdAyEw8c6X4xuzKswl9n3cEeaVgq0Ss5/sGKPPN
Ft1Sa07yOfRqsh8e1yb+LTjgcwaEemvf7bWwBt3YniUOMaYckM4e+cYwQJmOvC0r
89sgkCJxi9N+MokQTFPyExWC7d/uYxs/umeNSYjRZIFTggH5/ChiHimTYq2MeO0H
lg6sC8ZFpRaGzgNDbis3gabiRsiMmPxQaBk1wyefRKLvkfmstQTUxMvHE/YFli09
uT7A9wrMhrW7Nle3D2q9Y6S/CihabsN+IqfHGbn4qBBAdr/AqXKa6mxyMqxtlNkM
fgwwmGqwlme8oAZtMbsoWPpggzHO/825bOk5qz0fMitMXxQcltmnV3anHvnL+qFg
VwOP6bEgX0rl24sqcc5sBd4d83dlJaMa3waYbFXPPP1QlA9r7vR0D/5dOb12towc
W+eaeql1NwBpqeT/jVFq2NHOahwdodOi/UqrRxlK1GnYRqQ/UPa1l43BxHpMcwz6
V9CbMIsjGNvTQX212nePXxtYTYPpSrM6Vu4x+8E0ZmSCBBmr4oB4mfeFnxCR0ohJ
hsRpL+hFngQt+mGijWL3bh4R0zGkcu5s3XxZ8o2G2ulIMk4K7rSVaKEOMRxtXMHi
ua9P9/zuMm0IuZ528tiWWD2dmUmMK+aebqp7Wjo3PuTdj25aMWwkvet0t3aIShOc
HWVFXcKc34Oe/u5IzWJbE4MaBB0A7/yPZI9P0CqwmHLGd+VhJph9HnBeVyM2FueK
4OQkxkThnAuFuHqOSODRzoHMm8rwUJvdNEoaH0rxC+zLiyZyFRM8fJobhf31Pfai
e9BQh7Xl+HtdYHJ5avbMXwibBiWLqnBZd8/o35UZ8rtppDTnfGE7f5faC7jAEn8n
KFuttvvG80Ivb9Y2MoWUcyPk+7M8i2Maan52SgVEZLBUgJn7aOdgiZB79xVQiogP
Sxt1UvWihXY5p4SYrGk1rjkaMmbOpme2tvy5zn5VTLWi6FIgL2qxGkxweEpiMrb9
9GyLlPTA9T2kbHmt7M4wj/bjlXecvdkYkJ36eMQ5NqMc+GuWhIdrQVDMcaXAvH9O
V71ZBoR8BXdrIdmiCaChFoMy0HC7El6ydDAFBJWn+QvINaI+KoDdORUh2ysYjqYp
XcZu9SC/7YVJTylMKVuO+yFsDD3E5YWmRj0dKOKPWsxcOWbhELWaqbhcIAsuaqGt
xY+c2qmIDFql/mS1VhDo+dGyDGBzkqMwwMO5YaX4y3VRBMAhNRC+nDk/6ahLHQie
9vOi+ylN0XEgLLfpq9LuALnLZrYr2olPd4zOv5V8q1n9q5QfLoIIJUh/hoxYN9ot
H0j1OnA2+7R0621OZSnODVbf9BHKYsuVkiCl+vZRkfVe0N+KE4QTRoDp8HgNmnBL
oc7q3HaNcecpwhnWThS35XlkskKDWWebzP5N29Nj2p3udVA8zNJfpIeKtvObv6bz
4HLIF/n9hX35q204G2GmzU4JjGK/2mGmPGwLUB51w3zgPwpCii/cRWp8U044CtRI
lx/ZqVu6c5IdwuIdWtSRGHByPaknfulntLfG1e9287Q24qdcTNnqCLZ+IOvrJ+8H
NiRVm6Vzqm0+5IBty6VEPjkWTLCoDpifmHVjTcOO6r38YJRh3kRhasl0xYOHidOu
bN8odrdXeR2yJle/CcLo1Wkx1Nie1vMv+ugQaEY2HRoqy4DdMtngDQa39XAfrLe7
MeWnMIFNwQZZRUVDB5KjD90c16RxsmlpIoGeUzl9+JvwkWMmZrHdxrzieGcBUrZT
VV/LHxs9OP1rsVcf357Nz/C8h6dt3HXvdGX41lsvJlLj7vPUawAU5AmH+wp6iBWz
qODbwyiNRPP5TxnyTW45FWhfPmzqNGr9qbFAdVD1SdXEoGYWYfdMfPMTEZMO2lh/
Nbi1mgnlx49GiH1Ti+EHh/yTBfEMfn+y6CIcOcNZ71WUSuzCQNkpYaGvG2IYFps4
MXI0zZqpGVImpg1hyyU7iMVbzz8dDJIalqDxuADz2ZgjT94x+Q7qD9avqpTTqjiy
4GZgcWBaDWZJs0qJeH/bBOyDALf7n+Lx+Fydu/OoZHftx7hQxMsIyZifdhjfltdg
sIHpDrPsDTznuG7sRlKMTELIjKVQPA/9UIsn2Y7VCcW3TPynij7WZKdPn+eVjz3Y
szLAeVtYS1rNZOzBoeRe7IMGNq+2/ffGzm6ToWdijqj5T538S02kPLOK+9EXSwos
rMhEAedmwoo5h6+2/cTxLzQKj0raKkVBN9Y+qw7mzCALo3R+ritjaLuCjrBPjEP4
4BgF41ly4gPh0L4x0Hc3Q0SxxfweqzOmVe8WfW14ER4Zoc0q4rjBAyZ50IC3LmE8
heypkcQi9jRuKOCsrRavqxqm2/U/962sfPPZoQ1P3W5r6sL8ntgyFDLNnMPuRIQ8
zjl4rSl5Iuc/Kqa08w2ns/UCxyALeJ4dF8fgerVEQEaKbZrjeZwwSocwr/aiWYZU
bwkrnx2SeOpt4wRUsenTyt5qE2g6o+1TRsPxUM3QaZ94PJQ0yBqL7It5qdqEtOjW
pZ0nsbHutImcXREljfyZi26YDX2y6WAS808ezkcxplBZ+kHuxXDNCJd3jgiVx6nC
DgYC+pILS5fIIwvV3e7070VJygqwzCg9qGlFsIq7j/Va+SWBomnx1tZjMchLtflS
eMMRsNA7cMmn4FBZAvTyI6ViTKywuy1h7YUxn/nX1qAhofXUvpRJGD2rxb7mntCJ
36XXizb7qw279iXnmLnQHZj5MjQmixWMxj2A3gA8I6fBW4EZ18dSbm6dtojtnIkj
YW5uzODJfOOBEowo0RzAuVTkez4bHuwUC1LlOdiXwmWxQNyCDMP5LdcT6Cbemzjo
DfXBPOVZqh3NhGuMenfEhDNEo64K0JOLGh2XfEMKQWOSs5WT0QPD/yUs4kBSmhlb
/JXGYPEtwJq75D5YdEh+MfSaH/4gsFJupS130GtN7kl4WyyGW3jVVVPEo7RmGXL2
TTvLRyOE65FQL9w0bGR1jNuRQXpmad3npkGI5kgWdzhxaoQMgkCutOxd4uyf2fD9
X9d80+wq/hSXZQWpSaycY4JtmMTFEMyrlN17qSPrPBL8pz0mznbmrLtWbtbgaiN2
EK+Tck1S5lS2P1B8ldN+a6Cx8DsGeO185RSq32fx5jBX8l7HR6GBRmdab09AR4/F
otgTg84inN2ReFXGo/as04IT7oknMIqrKUHxKOrXjo3cnin6r2kaxBhgvYA9dpIa
/S+sOCrh1dmN6+OZ0gnR88CKhCI8pVbygUl11NlBqvNsGm1iam8gzsAL0veNdW3q
CLX/EhWZvri7e5AP+mhcoC6WBeU27Jb1BE78fkwofhX0lSBEaIZ4/KyuJBn01DxR
ktEl1Gk9qdZkouyp5SgcKIziZ2aNIyTyrZuIaAVuJE9g2TBPEOmPwaXedMiBB7/o
FyYtk8/CDW7EfHAtOMrcAW8932hbSho2BiMUr+gx9RpLQYJ+3WpWxXGZ7MuJByfl
VkHsESbA1BQtR0EfeQAcwva4QxLJjQnEUyo8OKHW1M+fcIcJGUN7EIa9UYzpXcuD
SP0Ir9rtV5b3XU6WpcLNW9xkFBLCXILhmuu3b+zkAAzpOS73oivpx+rp3+u0RbaS
1iwdMPw+bw9YEPWZ228/FHebSbkn9rGk6EW0q9m+/CuyEJK2NZNjax+adPreQutr
3jGGxLTuEUdCKPCHCRIoLEJQDnHbCZyLjdgEy+K5bCpaKDHyH8YuWvjFec/qD6CP
sY2xPHn/ZrNpAeV6MHpU+5GYlK+6pt+6hDEHOoMiQSsU9bJFQe1eFNQGd0l4kvGs
76r8lSveMxeckMho3d38MiTaR/PXbGcuPK5m5H957YL3o6GOMz/rR1WESroT8KxT
7hoD+dup4J5a6US+2/KpAW7RETXPQBijHvPIpHag+js5M44ayrqDayZlbvWe2w7h
j462u4QCDJXmDdB8nkUJkM8FIJnWl4VkyO/NYPCHap3C+McElc+DHiFfBE+u+lVr
dwKX3FQ3vvG7cDq/j5qb3IyszOcHFK8vUPXqKVTry776A5NZyM4/tE20f0AuTRFp
pwD7+47Iw4vgUQ/+dkx7Kn6uV+sYNj5D1sQ91t7El/kqYlHMgsNzREEMO0ciNYEv
51+V5wRiBKh8rVHrKJv++FF/kV2t1GMtbaxrPddr8qZG+X+fX3vbuLLfhiGpFAx/
TR/E+NyL76f5kYq632mVzlFkt4r4NiL+i1ic+ww9sGfy1zmDN6IgR/MbMRyUXWoP
sWUCi1H8Q9OP6Io9IK+SVdgV12tqPdD+mBkzYlWtfqWO8c6yQ93fu9OO0DxP+Dca
LaWDumiKuAg5gS89ZD1GS2MNP5JiZFALCWLObTxxLu+YpbiIVFzVoBPLSl811HAk
9iJ7squHktlSnn3GerorJKeuA5TYAsVOXn5YLdLn+SkI+tlmwf2feJFP1QbPt/5+
3p9QUMeHNPzRfM042JMqBM8/tXuEugnoH5i4Kutrvb0LY8NZvsHmsh5Hk91qrCIp
ec08ml7vFCQ9a3SJiui9cdh/4vinyTEKUpEu4krbjc7TtW0BaFw3W0s4K3svNHDB
/Fxo7T0O0NZ3qqGGHSBx07w9dNj7r8a36sVY3aLFEWb9sGDfVbwscemTEyD86QgV
ePDYjhcfGabxfj72CpvWCJuNHEDtCXmX9egUMMHJQ1e1Sj2riOaFTytzthzbH4lb
1UfVXrA+Hp5FDl2OQcg4WgPdl+62DSmiD3574nMZkLAFX6EZ2b1Of1NuLzSXuVpK
VcCEf8z4+vSybxCwVnsv9POucyrWdtyf02AbxyzekCrAdbFEbqlveQIno7TUAHGm
cCRVvGMRMXGpykFSQGD5tKLTdEAwr/fNB4UFdYzSwJmheug9uckSzxkfVnCpSEQH
lY2LEnYqC/Y8Jsq78W3muP4grG9I8cZTqRkbnb2Sx3taNgLYv3Mq+1PktJTKaiEV
2IsJ01UaYhFIvMEobTMPo8ynjdfxAuybv7mwG/IlF+a70Z3tvp79isVKKV1Snllw
Y6Mgelrw3Gh8l3G1R0HwhabBZhPABEXzRMF7DOGF4jS34BPQEIsXP3dCpoBGeT+O
x7tZ4r5daOO29ffNlqzXtxSe3Wn8H01A0ei0imt0wDjcolBMoGys/SX+XYlCK2GU
OdRQ3TpqsbksRD7gO/Oj0OHXt4FN4+IAFmvtQMYvymf5jFWdicFeeMaiYIPziWY/
hJYwe0x6L1LOOPBG3mnSlfMrvPJ6duHRahVH99oMSlf0hJUFbqEY4JCvf7s0ARgk
yEtlf4JN9x4G3Z0HYCiXSgEeOMklBVxNQ5PVp8zSo5Oencxe3tdZHAifGqFPSvMZ
FnHopGfy1S0AUbPLpDU3pEuP6RIY9FOAnmkN5I+bMjCCQONkURv56Vx8wkpEeGVy
lgig/ecAIR3E7k+JoBCEHCOAOGrnV/b7Aq+DwSi4phyu73RahWPoF0Cr+hm0hflV
63E8mImqh+Te1dWrwK2GctkdbCHss6wr6CeCY+MIZuWtE9Znc3SpKHBnxzsXB4WC
tIgN1zL3lqI/q3zfRvvxtq74uaiin50S+GQGKVRIATIpyjfNJgekfzXysRWoPI0+
xRT8jZUm6JjjAsAO2F+wqexdhgf/tqdZ/HWlPRNzchSXEmgKPDNhSKklW74DMbe9
NX0jb4oD0KkLXbxUbrsII7Ls0OSVjCoX0DnSR2lT6me2NOrgRJBIeupDnjJhQzEf
+fvRReEVfyboXfoVqtdkOAaMiDLyjqEsIDtjjXd1Moi6rd5fdLd42a3GdhAL6Z6T
P42j4e81ljZ2PtaP+IOB4u4QhsP+hOYNiP6nWJ5TeCTCpFMB+3PkYUKP6MejavMC
9d+8/5bzQWHu/zTEEGTThV9qWe/hnrl0KERyhXEbvUh4qgq5qTfP1SJKKYuv6hsq
O6EWqUEURepniDO6cjH97V0o+/gAFhFbyQBWBp34i5970L/oU0UqVmCIuNFQbNGn
+k9wjIU8ZQFQ/vWhb4ILpTqHMWVQCPZHYX6fzJx0x/4XAr1uXULWY0ruksBCRzig
Ihg8eVF41tNi19H0bBolw4lmUsM6PnIxtq4b+VGfy0DhkTldB0Kknc7+AG3vEZAo
z5ACFLDqGHeP3U4WdmMXBOhXNVWAwVDr6UfEOHcAsjiEDp9A+T0xoKrNuT7ZZtIU
JwILLyoIn0BZIxMvTTxcF9sJ3rwrFWHHduKtOcU0Izv1nTSmNi1DtaKNSgIM0F2W
jzBcvdJi10q/twI/2gkjYLt7VHtRWDJKEQtdXJAffK0Cr1y9KxwE3/nadXg26K7t
QXctE9l68RdvDX71NGd4XLPf0r0j+Wf8H8Y6ecOYP/j+EgZ5W31NckQZD3aHZ05M
2BpfxLuXPL0p0pj9i1+zrK2W8pfZGnVDt7Z7haTQNbEGmq3RuFJYtvoTyhpC6/LZ
Xo4+i9/bm9cHcp+NKJEKayhXJiNDzBqSfQ2ZhOFz5+ofVFRq2VaEcCsRQS1rV5U7
0UG4/sVjeJhp3L+fZNWoRs9y9/HGm5vmSmo4vaVfIS92dpLqKNuADeN9L4AsPn2s
c6btRyYMQZ69BMR88C8Sb5Geh2DaTNf5uypiAtb2KbajUEvihOBnH4W9WFxJ/NWq
ORFBNFDwtGhCHSOQtRL9O/uE3FwrS7z9vfpHdUCQamhud2gLBYB2RzPWTLenRnou
v2A6AlArXjDBw5NI16GXnOg6JDNSNNPLSdsl4RnHyTO5igjDSzrmfhpXQXGDy1BR
v6Bsh062k42n+V9x4Xmvfk13TKG9PTuDiG7eRccpSwf1452Wodc8FwtH8I6aveF+
9qM4uxk3qNdCXYvbPk6ZXObJ/f+wehmf/HKSu6NB2cRJLshutRgilRI1147p79ki
wLnkoTZuC0grUc2Hw9QMw2q1+KTt3FCrXjwH8VDehQyZvRCUpc3bgPgdp/AutScv
QyylQgK7nkT4j/WgKwjojFkpNJiKy0S3eByoV1Uo57yJy8Q+VX54/87VVIdbYuWc
tEV/T1pwyLfeCox4MRX6W7r3S+b8BiWEP1VBllXRepDung0+56IGqI3BF/Eqd1x2
RwdEby65WH2/GwGVL0etUWKJc1ifQ6dx5I9esgG180GUKQVHOx3GBNcYSOmp0iBb
1ixPMQhRqorB3crzNeLJToUbtKxxSrtwdXJtsYgjGbHpDfZvqrnScg3m7XVSw5UZ
zXYAtwNIUhs9s5jKiieNA0PowGmGQQ/sfV8Pb/uSbV+K1nzELL+s4jIrzZJ5ySNU
YmeHBfnSJUYR6A6zNnVylxiyriwJ8PjpHpW2qHM9D999l7FV+tQF4cv4g4fQWmRL
efrW+YDEwIThZuP3OmucLAPoHmn8C7VXK5YhPbTasGXRkXvG6nrXI9zy89yxQsdX
Vv4h/IKJdh1lSZdDWo6KOtWWVi3Eo6KfqAlehxOYvjm9bwaJ9pRbr0O6R7kXljdK
/Ywa8wV7v4jmF21v8I7XhnmTsBJb4HgRNNzjsSFHsAuwYGELgg0OvlTWq537Ce5y
e66qbwXUhsCTm+X/3N9GwbRMbArpvB/wghHiISIExuVg2py1l/gyjqLEF4euK6FN
b32tPe0BIGCa9zgxM5/fzjXDzvJRyTHbSHpltuT2kZawZXn1pqV3DTr154MieNpK
WtwH13BcYiLATZaOARLrFNmnM+jUrUbTvi9Gn/Ony61hYpWHs6ZQO3RJrlOaV7ab
oCvtPf5ccH9R1E+I+rLGwcAyFrbCm/SRoifdc4X3IiFZxKcQ4hz3bMEU4zqahGtB
M/g/pGCboTzJZiKf/uJkzx2/ISMszr5yDtiO6Kru4jAxYwgFUi1O+cDeLSjAllWn
QGfcFzbO6cxu6l2judohX3dRx3HAoH+eAi+K3DaW1xZjRNFDarapxIbpIaYq+kUi
6ByIontg8WWivWVHHtpGnTvcQVrMaemf5bzJnhRvspRPtbZWFTLU1xqrnQ0gbDPL
/IC10tWbAzuCNvajenBuR9wRbizVp2LIiXA+EJ8PaZAl82gws57SauubA7ABNBdl
xzhINImZB8jUEnqiXdSiLsaSf7w6AkTw4qoJKoHWJiydoolZDsohrq8cs+aRQCKo
kNFqgLHxY9b231B7QfzbdH+U+5Eql/YozUdDaR2Fkxgii5gAqE3JAv15620BIxvF
hJcv4aKeRm4PAk1TjxPcv0zRi6gCpZ/tIwsID+Yu4hBSflpvqNI8tbm6yNkAWZYd
XWu38NUu3CTiXYYI/IbmPqB0OMNoQKqvZoY/sRjTul4zIfT1SU4pkBWlKCocppFG
Najy6yZFvHuplOK8IW8atdinoUUrqTj977tR5l+/QjeI5YTLOAR+qkuy9sRiuE8z
tHrEPmB/ftGmHb1iYhM3LGkXrW6AFMfuN2+fy+MvBl9jks2NO+Z0LNpj8+V2FBLM
bBs54E2FZjin0HsPNWQj3s83AUzUy0jCLgLQhLHd9f4CDhTFIkknpWL3t66L3nEX
Qw3ztlpF9bmVjX8pdtBzEohBlMMG+KLPLLVWySMeUbrlExnbfAYioVC82PLv1aMB
cV+sUkmvkPsYVdFdO8WhlDfRSwa4RY97zcnVbXmDZEuB4XKU40sKeGd1/Esf8PXa
Ge2GtfCT7novTe+vcpLDP+4V4LuJC3UnQtS1x+J7Mg3pL4tnMmsirGvkV0g2S6ZI
nLyRt7CXqEKRwCmr+Cp3z0fI/g7IcojOQV+Ydd3XkfL5kleN6oNOXZKFsrfUd8cn
0Xp3HSNJW/rCOrzeKQub61FbgL7mb9TvtR509QHE2FzoQGLD4XWWqVNwwgZVTztr
N6DZL7Wx2n6gS5bo+sFUjYvTU689Q9FR7VcyxuELLvPYt2rohZO4TUX54GlvhG8M
nz15mJKo2ODQhs0YUyHRM2jCxlrxG4dtFynqUYt+PnwC2XXP8Eew2AJ2INsIZ1OC
tBQwnQ+UUYufMDeE0Kc0QvwAVy6uUG/cZdc2anQbBcMBEKceGLPtlEjndYt0qRMv
K/xOugwTx/GUGVgEUAC7HzmVTkvY7aKLFZ6uM5cdM0dWWzCurrTQzDHLG+z/0YdN
bcSDZCbSujbMhpvY3Ilhmr1Z5i1mlMw4t9iWqa76kdewcFBYwc2cYpekc6ACHDim
YFQOaOhYIsj/ynZ+7K1HOTwpiAXoV3tmju4kkKui7qRnOwkWt6hH7YANySfKI52R
6WrJz8iYU3ayS6QBKnngcCe/A1es3M1hfLK4XqeEjbxqA0SVEmwoDkCt6/Xgov+S
7hdaGHg/KvGa2XUxG94W7wRFjB3Ik2r7n2MdiqnDJGCCdFVqQA0ps58fzD7GZRmI
Q1Y95jWgm/3d5NV7DEAYgeuvbUeJ7Uw85J6exl/0NOkpOBq4GrFeF6hONqYR4Xst
wlEVYvHzPvFb8bAazX6mAbnRmAcy4uJqAUb8J34WqzNPEfIn7Zg06o0WlgBXfHAM
+oidJTPKtrSg8Jbc5myYw5e0ADlL1HcickV5fBeA/DShzyXxcl2iuaTnLJ9nhNme
Tv+lvXHLvq335bw/cz7XSDG4al1d9dJYcqcCpEzVv8arVdE/7LmA7J1uPHMsANCK
n8zQvzq6YCE4350MjWrV6qk5NM3OQ0j9u2AN+ZT42EHUb9AKu1Ma2NiHSCYEEVd1
oVULcvD7DGAFF3osFkkAutM+VpbA7Ax3/pR/Rm4Yek99MoCdMEa7ysOGYZqq7/8/
7/wpdDJMASa61vqMc+M4QglII+i+sf8/o/pEJ6j0tqIPdpgs65po4hJA9D4Q2Qmt
1mn0ZS+UMjdHrr18veMj+2uF8/KVn86WhRG7RfOlRGd3vV1QpK2RsAV3EoM8B7N2
HuOjXw9yysScibNeuO0/p5pZ5hClBwLeagZW9pOD7ralKRWZ1ItwqsK+j1ZejYdi
ZV3g+26W9vP4/zD4s1SR1QAKKZSScgZrGSklxpZKpkuTaGCvDt+77MevjmDvuUL6
GbFh++/vyvNPG4iZPo9QNR8S4mOAcVHKJR9NyjRq9wjvOcGngpL42XXw0HYFHsQU
yfogLjY2qvrv/uX2jLhjfwA6fjI82YtpqTo25dmx1jF+n/xvxRZj2POFqQJ7FBVz
PJWt4yLeM5aUOlKZ2IoS5xm2FJeckf5XnVNuQ3i1qYv7IBHv8GeBfwuNsa7vTJKj
S8SGwol5XmoO+fOdZvT35h4voNkphpU9XyKytkl+Hwrofo4V8eL+SbX9cJGqmlhs
krruXCm4r6hpvHTShutKtvJRKz7TTfQEMHM4a8Uy6uR92w6Cadur+wWHS+PkcIDq
6/6VoXb/1rScmgtVOOs6rfTKx9BPYtj0didUipA47bBf7OGbQRnu7kbRYHkuwtKN
MRuCxCUVnKlLHZs3sPx5ozz2vBa7ZFdroTl1Gjd+Wl1uKg1X+FfZfz2eoYNsJEci
9J+hHHsRu+SjmoK9AMXEjnHcL+5U1eKoLHXU9h1VGznshZ2PqbSMo+DNJ/Sv96wu
7/pqjq9BA1K0jQozzt63C/jmSSr9NOE+FTtAt7W2a842yKLAJ+bNovYlkXoi5zbE
+79x9voMQlXJlzQZmDgnSkwGESsmgsm8I5qcCRINt0wiINntfB7cS6JHhUYAN8PC
Tc9Z/o0/UZfVoh1mgrF4sOkwlp8ihynwSJeNg7AUZ0RPsyPf9mA03coWxRqJ1vvw
T/f0C+U05EPDWiebbHwrKLuhtNpk2cMnKMcxbZ2XsQawRheC2/63NfL9DfIebVni
lnj8eXb+vc/PEd873SnjQbqBY/i8n2sgEc+1kUElSkMlEyPMDWyOeZqATLvCIXE8
84zntyd00Zd0pJsATqxb9qruh5ArEaJ1qERQ8nbiPzkoGdH66HVgwTfkyuZHCBO/
0KRwCAsdjEf8PDbhB9oMqFssNJ0LAfmX7oSU7aC3nh0oeYm0cBPFMEEqH6aquyT0
qQRv7SShEu4u5bA3DMtLDK94b2OOso1vJdcJTSwU15tuw7Chi5FUgtMEhIfm8SS9
273wcGxL/A6eN+mKDDynBt3O1MZrzBO1TM/S+Re1HAUzy0/iSOkag1JfGQ/WLTmR
J2KyBhL5XMEhZONhQrd43UGxTE7wli5B3NHGOKgPFJM7weuinZHdfHv7byxdZk0d
68SXlUQ2YlhPGyW2p2plFRZYF0Tkq5685TTrwAqRkwKtINBszbb1dc/AxME2UZ+t
dwGWVVkzzlbaVhxkQWB+qy57SpizYHqQIuMMt5lrHT06/DfkSZf19WY/msn93v6s
UunEus+xdn597uWq3u0Jli3bb2iT+65SKKYMqs4zWyItlx2bDJ9yWA56fEZX46M2
vaoxYn4aQir3oloFFqvyoUPWBe0vBbp02zr4ooBVR49KC8xc70GqJ43LEYrxhuSb
3r/RvMYFfsV2J0EdiQ5EdSmIjHXvjRKzY7cgu0IZrjWuoj3YMj82aK+wcBIDNLVD
a+8Npy4GDnbngDK8Z2X/ZnZOEt+qGKN93e89jjmcWwwkjEbhKAUH1nTOrI7sWdHm
Any1rrVCvqYeGZNvoQ1iINQTVZUZ/cVnOnMwAS3Ej3Xc/kOf6vH/JkQCZgs/LhlD
+pjx/BdyZLoxwMNIEz0n3aY+0odeFQdFx0cLmab6rUfItzLPLnug7srDlbMinrHW
5Nmo9jH/rjxotRhZta1WRzRVehLB1fzVey3/0AiwsQuYZ8RWGQBNqeoS6kd5YQZS
He8P0qdAs2NGjjc4t8LXGt37LatbBBBHf1NZCPIZGFcSTu8tBTE2VQefarQMbx2n
lVJKC2GP7+L5714UtzT8kpT9xJmghjwFZKuiLNjSRIrNep1lMSAFrdzbM/RZJYLd
MsyqVzfQTDdvDkAKDLLGmtgACvqGRvYoxB6uziB2VtNj2kY89EnYq0mnSCOIGnzk
YhgS2/E7/5GQf2hVGQzEE3SNHPbn4iCpmsDYTEa7ZhBMpv5utmiXfBDrfVtb0wwT
K1IxZtzY2uiQLWzlg74jv2uxRsbMkrWa7q3ua4qhv8rgdEDTvkXxKBRisVJf+zXy
7sy6P4FcSA5+tsNgfcGh7Adm8yFUvE+AquXSyjKa7aep/2aAuBcv1wh0+juyVwD3
CxzmUTXsgtA1KDPecTeO86jqKt2+PTEuAGBItBhqSoHdTwK0dq19CnG76pvfYMk/
zKe9TekdUQh9fl7izI+d3VyoBMP8ONGWDt7QnfhNiwcpenN5xlX046QSVtbsWzv8
pZtcAseCONvBhnX8CQmxh5BQceNlRMNDoG+LM9cA2r3HjvINJZsPCSLvp9paJOUu
PjPNFZUkBXsglWgFgNYFbiUtDHfULF0cRY9HbOxj/czsBxeetXt+lV1v2381wpxq
PFKTT0TW+BrVyLkfrzmayxDJwmWflpOIu4dg7m4URUqc76PqZ88gUCB904ZzfBXN
WzGqTS5oyybhiVttjrSEiniohqutfBq8+WBd/RaqSm10lw5xbJ9n+ef73rD0+3dO
NcmHGnqZIT71cN7uu1be4JSns/O/1EAXUj65xmTQ4c6ahcpMKijwY6aKUHFVxGw1
5fmL/LQug0Lut+0eNlKVhXIXI4n59Lcwc+N6nEWoWhs/DTVaJLIiaL+f9B1zz3F1
5yuKT27beAPZo2Ch9fSWkKKJ6EoD29U2rSAqeFagbtMcBzYBOmfnKFTrGoqGMqDI
BA5xgjXFGpX04FwGDURl9LRzE3avvWS4Cd2grxiIgxJYeCkpImS4lkW+Worb2DPR
dnAUgEyrGECSoD++36CLmIqYpN38cK7sqMosA7AQ4+6H6HCl2m9Uzla5QmZonIti
i8jrA5AJV5OtBjmk+8MXuT0foX2SX+YnhvY172G2PIaVl7GyVAYboDdleU39fose
sb5hJfxXjDAev4LT7O+3e/RFa57Q6x/DBpqka4cgxANZUdTrlQsI44ouLxeu3TVT
oSxPIDKCct61obW3JZQZagX0lqRYFvNYTeACa596aP0xP6ZmuB223kL0IrRmEDys
sq0e1vCmtI6nDvOPUhBwe2sRADO6vWxx4ks129zXGOAGeHk3SXp2y7dS73tGlcHm
1emGpCE9jJTEnT3htJ1U2l2SKYGlXXEEcdMBzRv8JTRvUMw96WuMutXG/AVeEuxQ
FEzUOWJ7FfX17nrmHgtk5ollxk0L+JNgiuANHrMsi14MDSfuPCuFKbqyHovCzj3C
RqAolviDhVttK6c3PZ4oj+z+Ys8fnbrLo7Cfe6Dk0EKBw59kC1apQYcpgF5S5Wz4
xfQyD/UTRONjvFw7XyYepeiwYryeafFsx9sllEaraByFjPAPh6DnxBiazq+mtr/a
kSgvEocclWWmelCRXVp4LQlLPlO9n6+byZNEa9pW3ZpqEOVN1QRfxRxiw+gOQleO
m1VP+iqR9pHgqXd364Lrg2NY+F/EjXxhxlZU4UUz5Le8x95yE4Wx/JJLbn37qv3l
UvecSl2G+nNQWzcLZwIl495ijD+hzN0DKVHr6ngEqbfAy7wL/ECp35JfaDvCoHt3
RynD49DEPV+fKtI7dyYb1QBOdK5/e57YQfVHndjqXrjLTZxX2HXikNoeZTnAlPBk
wPuYbxJAfpSy1AcbZWBFAzBqTwFhTii+t3qOmHaIzqqncoEVFtnXU3uEp2z4wj8S
l2TyOKaKctUi6Gc1Gs8O33f8sNDcUdx+MhW13eORRt6HNmY4l0nSTA54YHaA9pYM
XFuBYl+TJFv8BYRAHLryh0SocxW91QQtevSD3nT0ov1++AsOzLkHbm+mpYtJ58bg
CBMtqowSMvid2pO9wBr5/kGHCHMolVOnE1aG5YdH+j1d0FjV8xdawhrMLydupQCm
KYAdU9va9thesORzdgLt+Ne8YssK7aJNkDIbX6PZc3jvCGPg0QSizL11hFTURIz1
Edw/FX5XCm/HNu/YxIphwu5AD0cvHUUQ+JeBvoQo4HQKCWgvryJRd+W8gZjTPL5W
H203QkEosbfxtve8MwQGLtUyLzanuPgv+RwwlNFSIwYXKwvPGG5gSoqURX12/BIG
nkrw31D/9tNdYMJ7JTbeUMNuRpJKlou7g58uN7uPCfvYfTh133PoT6r0BfZ7tzX1
UVI37VNdhIDWNTh4jkNK3r0DwqL0++b4wbwPiSS8nkfofBsB8YA1dczQag19hj6p
1UGOV+cjYko+bTLkave++twAWwvirWa7hLHZBhUOrma3SrGufQei7Rin/CYOXrFH
DN2TOKwpzXyPzPtvVQpbdAIBevyDs/pGwa2VGWl4GU/75M+cHOUaAfmHa9kNdxxu
SAoi5JKdmeTzz7grvtCoWah8zWN9SOnZONHHLHuoWcXhUh0UQnlDIBhOOzofSn5w
b6vl2q+Uwos9QsKHKWPKqsZdgKuIno6pSkT/EkaeRu2kkA+3+j64xjyzL5jl3GMx
QlW1RUiBPZuaJHiMt83FM418Dio6O5DZs1sFfQX7YyTDgE9mPnDs7C94m4e2Zp4z
k6xWfXkur3ZMCfbr9gaXTjZR6/G+R61m7IRfpJUgZcCHBZ2Xx/5pSLPASosNGIMt
jnJlInpouhWQOdnYelA9+ZeF2At+tY9DrQ61trS1vPI2lMm+2Nx3bIymJNKMCzkg
awp25fyS+vHJZkmtcFgJAfcAcqCt9+aNyOIRu9eCcOwbYCi1d8qspp5EnFC7zJ2K
ow9p9+AdWVx6jKo2py/ia4FsDGMzo/rnqMbPzlLC2Q6MIqnpHLALfQyQzvXV/rvB
3bl6sBPCnNLaEh7OJ6abgKohK03ewk+yE/Hubezn3m8qEvJOSdAfJ6ArLMKnjyXz
GkvzcKR2iLOBX5ju9sjvNkuzW65rwlEBZOY12eQHig2u+9i+S28Myj8VuXnUFVLP
7/yrgpsC2y88IKtGX8VpPM1zPKSQVfkumKX8rm8xMJ0DB4G0I3jl61GXvRoufDnJ
L8GZ4fcnbYSHl/rPnXhmbZ5PenZwKZiPt954lLHfkYzByrXlGVvPgRR8AfSjmy6L
VD/hC6LNoYAKsEimnMGQUfF7S/FfR3Yd/yBYbIRBN2f9R8BUPiQH4DgUkJPxZDWE
XdbfGNQ66yVctwxhQLCxtiRPmrp1DkRqoaGp3Hb6bFXnwxILN1EXco8xzo21johB
rfz7tkV2ZYGLEYW34iVQ9S+jJYAIdfsoYiQzRfRKv5UB/yG6ELzq0A+nF5ocGjvM
geRbdjjDCj79tZvcjjkv8KGiAj2jJmF9BtZHiFAzh+TTMHzRU45M6SjR+0s4H0B2
VHztsLdYG4Db7itlUSF2JJtQhLLMtpLgcnLiZfJazdsP1URd945xSX2yN1WT/ulm
6htsx6xCoffl0z2806+t4sbCfUZA//J65zsz+dpkTtbDZ7UWgin9X5KmIXspFVv3
2YKMdnftuRZ84nZiPMQCDTbfiU4tHr4eEzUBwRvR2Ph/3N8eUmyrsex54Rr2sL5V
eLU3b7UZuC/xl4cdH/d9acRXtY2xBreey8FprYkF8gXD2pwxsUqbeW3ThnmTMCrs
Yn4hCSZkSkhZn8uN6LDRc6s7qDPTBNc6wwWFpMU0crvqpJXltPHQXG4WwrrrA6b9
P1kKXfxDo/LBfG80VXRHdrAfsY0OKyw2Gbl7qXKAeZc2NIqN5V4o0qiQXWF0VAcW
CXtK15YfHAVknty1drU4h9ThPq/AOsiop4tkvZsXRzVe/63Il0j8wKbMvIYDbnAA
ZsbMxuQx7gdU827kQWRopk7d22qH7H80Msxn345IwmcrQh1N+af3OGpJb4p9oDzK
DF7AtlH0Y8W3kUJ2hvTFwfXcK8hTn10HvHnZRJk+Oxr2oucAViAKHtw/wRp628wz
6WPJOrreSHevd0yT+5LKIHpZFbgB1/VZMnXX74N6VybyIiIKNR3UbX5EMC8vd6jV
8xnPFzeM1InZ8OmS3kenEgWhtV3ccjRE8uNTg+pm2WlXt08Mi79QANl559wq5oS4
LoyYcPgBNtPuUUODh+ath6GVvXPBLx9EDqFXplw2w0c42A2Z9Eiei9P8l8xj8eW3
TWoVQzuESbJ9MOSk879TKpDEItNhyGK/JHl2m8TL2I+fz6q1JKl3n5CNoIhA4o7x
qfbt9CnnbBHACV+tTaTUHDPtveiEsOu8tEVM6B87FZ0OKRwTmWIpFCYWnAYXdNZb
DAhishroloohy76LPdnGoypSFN3RWyRNvRPRcRj4p/WHuZ5fldQEMIyPWIyoHTte
0cvz2wHdAY6LtH0So0tKoKhy1NlQNvQsW/DSvdfIgd+1IXhz5suEBsNbWcAXH7zN
bC1/DMzKRlV8I5lVQAfIoY2vZL2cK69Cav/E4mF7N209GmUmdyDKvJhhCIDvfnfy
C4azWn+UmXB0Fq07e6YRlZiDhMq5umUSwyW1P0n3NnI/2WcZrq7HBWL+RpRhzvLb
8ImtaiAtFFRji5lWGV73EcAyjOMb8B12gptkuczvWBz/Yj1DTXN7qkPj68tj5jgx
IiD6g7wCTTOoDXkD4HfzoCR1MYuyw73SXUEXcPqJ8izJ4DCuSk93vC36zMoLIHzB
sQLYf2NTlXVcAqUnzuFmNyEWBDpPbWGRkNXiQbgosZi6/6HFBzTO7xo7+zlyNGEp
1aAQwAlmqMZciYPCUJcqX2yiwsfxrQ5USlFHoiMSMkVcGmkcEKcTiABT18zx5jYZ
bbHVyw0YjxFgimrobUK9zD4uehf7ucCBVUcFx0DdK34Ack19RfearXH0Dp6OrbWW
2gZ+rboU8Ftx1rk6CHww5iCsqMJ3qW8ZxAvRzruvFpAiYux7yhRbVxMc1yqhEPXS
vE4dfnW9dEDB1b5+VUDdLwDt5G1xenikRk8P7nhQtSwwPafx6vaVovEThRov5N04
JLIUbRWYSXqZtKT8hn5hhdpnZRolqXwBlsY7ut67ZmGsH0ezs4ZEogcfLe75nDHc
WJ3kmAk3YuzNKrovw9gCeO+FEZFKDhhgvbIu/mwghTIIJDIUnO2w47ODPNw6A/Rn
8be81ut4174iCz10g7Y5fuGuKwd11Ew4T+GHLULrRdkIOHYyGFu65TjZJXAxFm1M
EDuYHgbTm5j0i2FQF4ArZcnGwsfgazz1tp3/Qe+EtA1fvEl7/bOAm/bWN7duf3vL
X9NgZWmInWAH0xgVUKQuuQCGRTEsNjrOODOJ4ASJc9V/uZwx5EDtUJVxz0AQUYmr
19doCUAQjJlUmK7g++olk/MrtxsydzFAKtaItCTXZizVK5NTqKsCYUT2TLzNcsdF
P5otBJfK0e1RmCe6n4t9rY8bAWkJ4cGvPp3DX4XZEeCU/CYYTMgUREuwI+xcBE02
ndoVQhR9XTl7bFWVtFCi0l8LdQ3RAKzYoHVTN5YcFBbgWCtHhUnRPzswLufBPgOX
WjzUgwN/vq/r8VtXMB41Sh8WfSefZMWc9Ol43RSSzGtFL/CQvHuv3F1ZGbadWu33
z5pl/lyqFflwLxv0s1LoLWd/ZG/WATcwkxFZikHbXrwnX9yIBDKfhAyUbOrgzD+3
UrYA85ebiz5vFjBFX7l6Eikv7z9BEL0hl0ojVyb3E+w410ZR5ZV6LL0q0hWu3bFm
uYMHnd/KeF9YtX56Hgk+IKpEIC8G4rzI5Tnu6uxfpZp3mNeAbg7lxp4j7JxoU7A1
+YuUIKMz2VzjDo09L/yPofw4gDYODc4x+rleHaa/mnF7RZAGTDNf/Z9Y0cehaCjF
j5ejlefP/vXUdyAqbVdqSDw7+/TkQeu6RZpdI5XVrEGbFj5owne8oT5X+VbqZLEO
du2dWUL/cH628Kg8D38DNR+wET32fqjgrmiZ0cFuTPcWTOQCzkUkUOYRzF6cwBHv
PcXVAB2yMEV5iguM5Sr1N628lnnHcw5dwOuKMULpmSVangIVVUgTpsiWHf79p/vG
+vo8P6xXaieyG0e7InI2C1Mta7f4SbmW4IZzuxyoMSAYSf8Gi4LrqzAbCgrngxkL
cadSUm802WIDtBnfdJ0xOhgXvPHWZqJbDkjY9ZtVrf+TEN1Mh7xX+/Tl6kZxE/69
G/9S3jhO6KPvHkndqxUxgfTciGhc1GK2WLyAavZ5WOJla12eyLuLdrTrKp3ctXIU
BEMq1/atR7pWNApYc/SpI34dh4ei6PhuAkun1o+aBsre1N68flUHe3gArbZN0M1G
LdLbbG9ejVGlpFbnHqy3bU4jXAyFa4HieIRq2UPpKeI9bsr13zTpRFBP1tc6tIqG
OWncs/dbDFbqh7UdPHbrjT1Yqc3Ir0Ql0wqIqLkECq0xSB9YHXswLJf80JyiJjUb
B77i50h3Tj84ilN4hgMmvuckr4gjhcbiFGlDfG+3qJV65Bz0Bi3BkEi1e2Mo0tZ8
COxaGa/+LgcxZu2AKor7SkbceiC6b19MczAAMARPXN0iggOm3tsuV9ulsgpkO6rD
fodU1Gnne9sY4k61QpNBvDGXby/GWNNfRAvhKA10AHpnVSOItM1BYYXHfYsPcCCN
Rm7BKQHxKL7NKKySmSMGicFpTBZqG1+u/OCeMAzArdF+EH3l2jQc4opoSK5g2xrv
yqQYqD4Dn+5jF8rfyerpx1aQBJJr5u08EQ8teGoscP2ue0ENCzKmgjk4x++MWJwX
5xPPPVdXfFhAQWeDXExgKWwsIUnT9H0s9rcaf0WlUtM/b6JEXbukCnZXzcmBv6MS
UQt+a0WKvF4Qd7VRBsNufO3f7F6bMkbETviOQPdBdf2tukrim/azhhie+VRwsB0d
7XVSrBbRGUQI/p2CleaeyZBPun6WpURAYAlLPqr/qDWywfrEpuTiHDlutS+GzETp
NaVxBS+6WZRQunrwohEkvEzbQd8//sWE7Da7x/67M+ck4W0qvKn+eYLH6FmMdAA+
W63U/oinK1fizPoPFr1ewoKWuXBev2hIqyGhb0svnvUwxqPdGwRkfdbh+YYFsrxC
Q6rQvROpOSmHjDPU+KdEzunhwQ9hiXzS0wzrmaAcHmjzauzJbwhSpCl40JkSmDeX
fpGdc3/Izdb5H+lj5k0i4ebp75EWwIDPSodoiMLDcab8fkLg87v+F9BYasbCr0P3
Wxe04ZwSCewzvprxpq/PGCfJiPDbnDjZVCWBZaR90RUhJJDyY8H4SyBHIBUOgrGf
7u5r1yRCGIY/WBtEPBrc+LzXYC/RZF212UYPz/1eOUl6IxBqePj7EXayWXsSrHtn
3WunLddSuj0LBHlaU/AgcsH0tuCvi6xvb1/txLLq1rBdYELs225nz+hJqJbHJpqc
rDzn/iaadMR+Ds+eGxHWx1koOiKeNgfqKR5TRpeQTuZ2vz4WKbdHpd9YlYKXD+g4
CwDmJ65baNyLd5WxmiPDFK4UyvRq1WMBG6NzPnzfow1+C6rS79k5V9ZCrefWOi02
HCKhrEEpmbqrs01MwiEmb7qaUu8EpUdVebQailJD1V2QEsaKg1jh7S8w00F+He7q
JTeyOlrz7CBTIXhBFbRUWnSV3gD7yeIAuX+W+9z2EgbV9l2Oq36h2s3VmSpmIdzS
Vdpgs+x/GZP37sSuQZ7JTI+bbTn0gT74/mzdnzkqfNtDRwO8AzH8BWKsE//cCgbq
cyswt5w9IIHCakSzMMHqUHWyns7qLpKFdmYVlOJI22n/eLEvMd6HHamR0l5rrbTk
cF5NoAhGo2+UZSCB8Icyw4+LPgebnGP/INBMyQU2OH4h2PKyzP5u2UMy8cLegCif
rcznN5LWT0vvT530glUSX5QdaOfjAfiRXEgTQt3R/JSYTzaskhK3+3mDAgMHI/FJ
4+G3uKov2bFfvcJGZSwcxwd7rlzLW+zLdejRKJtTEzjVNysoXCSQJHIXX1xTwoL5
yExTco4vwXk5suPWHyewD1xZbQGuXHq1MnvZ4Zl7JZFWZTvRgcxPELjo0B2N54t8
44Dv0koP+oRgnTTwyDYHBFpfITwkj4PaGnbNvJqpgu16pjGP0Ej/BnHuB6SaXtCM
aRIh+EYqWRyfx4krKBflYsltfV0fwBHaG7aK0OIqT9Bjhk7bzoRSZTQ/K2uxUdnL
msH2UxilLgxDXBKW/NfpmsKwwcj8P5xEii+OGlPgjowJFhKzN4pQsezRabpjUSKO
5kj5csYzm29QwQB/2O1zesiA/jEjxirvCHzpMZuYrkFBmxO52gQG4mTlXOTEgLfs
rspaT2E3ZNeNi5NE31FRgund5my+zWkk+vMx7J/8RAb7nuYYNdUUuwuj2i774bSS
DEyb7vS8DWssSlq2GUaWN9SNPc6YlbiyOd6CwX09veKhiDtjh5WpAq3ulD+5mkk5
Y3zCzJ+UbK6f9hRyd3S56YcIWo4FPBEinFSIBEAASDfcr9crfs9J4qH+pTIiJ12V
UKMPXUWfxqnceaihP79k23EhGU8YGdxj5ZHzZ2SeLYqUEe1pE6QmSOssSJK59e3i
C+Le+9w1gnAjSJc4tmpm4Hm8AO55rYBKr6+M5k/E3X8USulTo1lXs76EeKTzaFq+
FPqp8ncCYYAsO0WYeILE9NtXXmkqWcJZm1ujyPyxEc72MZO6Zub/h3X5ZWWOonIY
S61sGZ5Gv8rzMtK4PCfQyk4Er7ONMsT5/su32W8KvIWnBQVKjb+FGsUXJ6KeX96U
H4K8HdjDmreLtvT8riNBu4sgYPEnCMUfewwtNeUCxlBmNI++otcCPFEXY9pLAbUa
DJzv1DjhNYXICspkxFlYbk0vTitRdDMfV2rKd8akjuWqOC3q20hrpKxA2fleQmJF
6bY+m4ZRuxUGUj6kbIFk3wfGy2dT7dBdebrAn/vGbVFVWOJNcl6yTa3iJ0EbvtEf
BGHZUCakeA4TSQuJ/Gv13Ve88tDo97JJt+dvS4rUs1daG75YyzxtmLyu94q/dj+a
wY6NGoOtCS51mxA6g6s0pCFmBKya2ggso58tQg5hlXp9lYaLKfmHbyV9NFjzsHVr
ZTpnk0jIpJnavbhnfSkOXww3hqk2oOm7VujG5n9726NL8ZbxfQviF58lT+jO3L7u
aNnuqJ/wCmglu85uyQOoKLFE6OrD6ZBgoQAS1tr/ZQaxDXx4kJKSoL7kkysDgR8q
L8sLFEDsYhQki/gGWLOXo2PsXNy0YE/ueaUPWFTwggA83DxsxmSZqyNvdl9kJB7z
1nuAcfBcuQ84ab2I8YI5YoOMXRKTx+/Go0oDWgtfhqHKhQnNVhjX9M63h76+k+bJ
ctr0sH0QGm5vr8w+zt5SC/LqI5MzmOas3uUVZz9CiSDoh56hJxUzY2j2wC8j0E7x
5XArK64YC8NcfcA2nHkSEX2gNH6SBXo2yEq7NvvPO+ZRDfySy3XfOpMVpNaxayGE
qG8uyjJiFTWUqqCBlKop/vYs31Pd0JlRdSIWJRBj9iUhSUsOl3rx4scAjdp71iKc
yo6vodAMDFe8FNzZOKEwani+Tz6NhZyh/0rD9WFL/jMlWAopwF1+EtPwxsz2VpOp
cLdruoS0vmvoY0tfbfybDaRl48MXrIcb2fr53ewiI53wPDukMZh6ohQvbkIbCapv
g971iihyOTLJWGYgR2N+eFmA2b56tgzPPeBJMjIKHsf4eNdve1gLT/hbCecPuKHJ
DZa1AG9H+gfSPYy1Qy0ueXZdHjnWHNa6Qb84K53GX75JWONI19Lg/xzjs1Bgte9c
ifRIPvDirnCXgEovVIFsx4kpgn/E7iKjMJmwm/ep0GyL/lfgeVgdJFD7cjGxA8jG
8V5oJMGGbNXkCa1/n151G97dZ/Vt833AUN28z+k0GHJzlF3Qf+NCf2Fv/uYVNx7H
PUp0XEeL3CM3IhlkHtnRvqyB3orZsFICNjF8SvohwGajmiPj5d7yD7S9muv2kP8o
2kP7vOZc7MtQe6FvA7+uRMbpwJ3qFdlK/KM2OQo15MceoYs0103grzSY/dWS2qy3
VAVPnQCi0VRGIFrg3fXjfQe47qqnJyzJBFVOM3EgSLoXeXddCZ2gsy5essxOsVVg
mwtugMJdB0VEGkIALPAgeA65gzLGRebRSlyKZpnwbt8u1ORyJgxNf46Z2FqnhWOO
zVP5owcqqmycrvBPMoL1y6sjnCzXSkiEJhlPOdYdOjyEWwP5IRFiZmSyStevhB4z
D24bPhP8Gt4gNLn/3r/34+Wq5L6QgyeyUgA1VcUbGDJlnxnrvHsdnlTcs73pHpV/
YtSGsi3EON2ltFmIL194RRPDBoYlYDWRF2WE7C5xfznab0k6wI/7p+UqXwbab7wT
hc5MWNnPoNp0mDakEhdMu+Nb9Fl448nZv71dFj/cRC9mPb9CYGN6d7EWh5lskbLE
hlGfqC4m/z9sfIscXaONog/U4xGAsAyoEHMvBfEK4H8JgQXfheQdDmp7MB/dXHhD
DMGUwRllhc15fn9jr2ZLUnHCALAZB/oRXkupIFvX0avTnK22DWBRJNmT+k5AzfWW
OndbrkgVm9u8spde4pkMG2+m16I7yoFMBB+9ZwoOq3XOAa+s/gcFaSguTiJs1eNy
3K6u97QOWhgS0mMq9024DHapdGsEnbHAeUJYhB5GwqgPIldPoApRs7Py+p05RnxW
bkr2DLYLDJRmerJ5UMA6W9zGTHjBhCAIv855xhLMQ40sVO+7l1tQ07KU0+8Sj+Id
DoOb7HulTe/Jdv9Uf2P15Qc5mbEHK3GQbAfbuwqh2r3nBs6PoggTYgCeOQUT45km
FoiR2LwKS4ohjy4fbRi1AqXbT0GZWubWcdlybXL4lOpRGZzvHSoAfArgTBqPu6gP
w/W9UyKmYGq+TqykM0aUZAlAm0ULAvfJotLeYwEBe4fmknkiqUxCVhAmsHireNOR
unqR8JhgWXMiwUculPL1gYiVO4Ooseebp3xkq5knjqbZcV//hBjXUFrnKTxeYIxQ
+WWlMxU70VvJt5tdpiOJLSnvDI1jJMVdB90/sxv5N5WpfDa8X3msRMZxza0FqKUB
5sVyoFMI6ZS7SskVKm9YhbgnDa5xwCyRn3vol/SgHt1diowCFAElENUn2nO+9JjT
Hx07WeaPJjkuAwOUM3nxuZeSLO6ZppvG5Ht1SjQaZhvdT39rU/iXbYcccUMVh9Ga
Jc9HcSKa73cemjFU5YsPtRcTFRIMzIKgrC9rgazOxqrgQZfVvE3co6768VY/CXBS
uWJ/ZnHe58KZJP+o+phY0mQgUSS218oWf9Ep2VknkYImVBlmvHveP5P5/7NeFge+
umyUyvEjiSE9AccyKOOHQ9ESUS/fauaQW+qbTRyAmwH1qArHgdSDJfO0yfv2Pgft
Nu+7mgQh+Z2bfb7jnCN0UraqMTbuswEamzwvDfgx4WVFI6CgdNmA9k+9yroPPmr9
bGOOEUFFsoMwVJHV9rHiwy+PhK8en1iuucBzVxT5YrC0GxP5kVglHdXfN+kzkpns
zhva7gLMN5GSe48XPp5qNaRjH4VmqeVrPjBth+TOL/7HogLCflzirq2rbyVy70Pg
mN/9PAM1G/p5dHFyyXo5LiHZXXBdGSvKV46PwpPqfF2adhzw4PBdQOzDRWqqGvIO
GI0PNVPrYepHJMyJFBcc4ZWs7pWaZiPH0uNLUgeQFU4AlNkx8pyw+E6P8PpDS5Nj
akI1Nc6ZePf+0Cuf1pNtBtXRMqPZMoK7/ep4PjhHkEN9aWKC9ZG5fodbnSaSNf1M
NYclFZDoRJIYDMztLeIZgBV7aiuMO7h2e88QXcXrZyRRZizPWRsvP+3c13vfc1Iz
4qR+F8S2RV4FWdCl5T4nOJ2k1jeyE2x77+S2qjSFHaWtAg9Tf9Wz2rLtkAcnAr8Z
jXVUnmImJh6dbrn8xb9bZd3o8oB4SrYMu0nOKsAXPCMALIZQ/hjTS3tCev8P8xUM
6Cj6Zi7/piSMpChzbNUEIR595tFG+0jJVaBzeynFdXeZRpPPdWCCmbXafBSLNAvZ
4XU9cZJKerouhS4XGMp09CBG5tZMTIeo1b5KKyns9hB/z0o4ENId0NYYY9qBq7/M
cieu6TMkmXHI7EqMMlcHSQMEosl80M8Nb2V/iJT3zz368wtun0kxIkksjW2em1ga
RjZQbBqgeXINTXQbR+G2howqA8NhwtXJfiEi01DSowid9ikxO10ad0u1j6zRBucX
k2wj/RPU04qLNuMZjwh+HVk1lIxaCks3ykr34DJexUQd7rnX7kheAduhg1nxMc/w
TDVC/toTu+RN2KwGMaKQQLva75MKYxpGAqHCzOLdlctXab0ieDKnxj7VCjfkZTfS
D8nD3rw7xf3gDIWxTo5Ev0rHIYayNE8SRfatHdnQS8WT3hzqAkeydTdgD0suz+sP
IfpFEjYBtLk5VzvZVxUqt4VCMrwTpe3PNMHFRKphEDEA62HvmWssFO+5IA75vqO4
4Mfdjmu2YLBWrljhy/SXNUCk173WkpLWXs0/jpF97oczrPygSMqucgpRzzLWy0Cf
zeFsMiIv7VJBG46oif46KAcgUVACRDVsNKgKcyP9pV6+OgVfPVY+V3+R7j8Tx3+7
dvQK7RJbh8Xa1Scup/hGgX8nZkEdS/+gToUT6YUz9z8G2kddbphB12ZNl0wKVFFo
GylvLwPe0PPtKyLHEltQrunLUw8q1GiVvpjlOnahPzIez0Q/DR6FP4DTGSur3Y0H
kHjGkKxc8Snvax6qlvKm5GPqqqbWaS1Yk3ecVf8ppPeOwufyrkq2nBd2nnem2Itv
tkdhMz8dn6jNR9T94BITwVTXWJCKr0Qb7extmquWknYsBx2rS++4fxQbTHvNxEZb
rJnxnQg8sbu6j7K7qJ3WWSMCMaLr5ve9XtVFJ3+T+sTeVD+zZ7vYMcANnJtf7qqZ
V3iDehdiq5NGIu3iBi2pM5FxhWfdFlGEajZaILjD0qXlVIKALg1qMwNlgd6mbQnJ
ziq7Gslgwyo3IuPFAVXBWFnuZgCQzktLEjlzMA1W2KHe8z6EL7bkvAitzSIXtDvy
7jJEzHD/t4E8zS5RqvC4ZTvQu9wugbdqw7en4fqqi1bEBYCjrxygcI2VSinR7ARF
z7CMm6B0Er9gO8TKljKB7FYapdpM1Nz5AtcPedqIxWBDcqnZOjvRwWFOL5i8k9L/
Tpt7MgBzOjfHkzO+Do+K2rwhVHmAAsC2iDY7zjn5b6YVsczYOhfR/pmaFMvxknUl
YbyLV67Pv9t//a5AtOCE7FYIbOdcSP+qJnV3jL4lsEEuD9TMjDhuhAYVUwv8K9PX
i+SWE51i3aA4NaBQCvMxm/iH2QH7f1apSwGg2Mwwnb5/wAwPLCPuUnWXGqP1BVqT
l2mc/PyB9ZduTlNMwElvRa45RTCmXELOqKWUmtXY1ItmZEbpKy0Xh6DH06Bm16uB
VjHQFHQhxuzSkJKrzBT6COtFOH+BsrRD5GBm7e/OZaboUcABvHVtxmwzxga127H0
mIhI2923sWn8HGoxl1UVHt99zKAS2dJsCg4yMluABCMMWnz1sv9baKEPceOMa77g
Fxl8f6xu/u41DZ9KdZCqgmreCMNDs8bIbOn6Xsz2T/r9X68wXP9CRYCd18QwdQAf
ngFWkyD4J7YIy4nUXHr7fjXCUUpTNagdPBvbwqhRzZ+OhHlcYSY0kpJz5HeHS61v
bvkdw+kiY+V2nVK22pPZADbcxjMd/YpW0IcE+XYwsHNRBjPrQe8VZbPd2ipX2LQz
JBsU9VzWwVfYHHub3rJA8zTPpfOU1PRWbZVgN2kY+JFOVgsPLBArFYOz5xaLaN45
wOVFNbPRd5R72P6e89d4Zkxajd0Pn7OB6wHcyJALT3fpQA+8d3iNikdW1e2nI/lF
m9iNrBuK2pjRTsvwTPtYArUdCJusE3MsAVqP3IWcolCLhrfMWQ9a7aZs9/ICFqoY
/rU2TrAPxLOrSleb7oszwHsO/d/4oWGLNIEXh7SZNScFCgSbcx3usR2OFW7+Plg9
L1LOpSUxIiBH23gII9xOULXrYVwS+/5b/jgPCHlSfwRB4AYzdY/yMcIM3Xf175ax
EsaBDTJu7zzd8dDhC/GNYPoLoc6GCe8z595PwtH6ncGpAl/NTNSeVTRxZOv9uULa
8eNuMJeioWDmeX8UW8Z0c5mSqau4D1HC9GsWItmNPwudOGnN3QxzTSx7jB3ApH+V
Gi1KrJvXjoDYfguT4eeDAkYL9DWNLYq22wT6ngeaPD1cPOLQWJ+WNp86RchAU2Yb
dsSuCGLIsvEGGSD15Ts47tIEDTmyKiOudbe5UKdW+pJXDPJd/xYQ08AFxhKK4Wq4
Mn0BLOG3jgsjNnwa6PO+K26AdkUvt/pZ2grgKxKsacHKjgnCDRDml/7GD3AfS1Hq
X7x64DULDDdOVYpw8gK6B9/3OvghMWx3nVTC5e6VYfDnnK5s6r1nqIHON1ZmhAoF
/XRqKisfzC9B1Cjrq4q7Olatjsmjy+hBSdO9b5hBwKxenngJsD6euysgST56Lvkx
aRdv6mfswnOn3LWYy4xDd2wV+BNnWiXw0sc6VZTqP2YLUQtyS5p0sUn1xMWWX++R
EpkcXbmIkK9FoUzjNZwjTSiUn6Rx+i+aQ69Lz6uOCylbZG2TF3vo40mUqOAgaHhQ
abewIFUfOHuhp4ueGx+/6dAYRAEnf1egebORtthNyXi6JXahBSGs8r6jRLACepCX
ELrVy540rG3+tD8+M3m2lbOAO6qlc9/CxugCJL8k8MAkWBZRJr7/K+o4m+MgLGWL
a++q8kgy3VPvusRrFuSqtNElDdZHs91oGj9z2T+P2iDCvWmI5WARo00U36MiD7/L
xdbfmUVjYHO+OVN6t3AhvDjRzoVoD7vhXf2LrWk1stJ8UMsloQj6v9T7RwCePaNV
wGWLOw4PaBTq++YmMYBpw+1gxMg5L6Lcf73mXff4NBIxKFoNBNZoDSIrizESqJsU
MUYB30DVKU0SqiuScTO9gXsEuRSbazl0g81IgIREeCfvJ+CZJ5a8/vhNCJJh7bKY
Vq9PeRwue/zzKKVYvAi61ozikm2sdC+7wNMEBEria/5h5tz+1n9BRdli0KOsNgsG
s80HfjYIDqWZ4+ydB2EOkgU0kOGFnQLe3jHMe4g4JtTPE+J4de4rSR0YbchjQsKT
gCCC5tYYqk2yhZS1mdUqEmmgKgrPyi6HloZYDeXF5dqM+V5XAQBZ6CQ9BiQPGUc8
Tbw0FpNBw5bw6x4jav/ZfoIQeZmLKbe/MXeiaqy1wkNf6czyYZo8gTffqbgYBGcC
+kqDi90JmlJSN69vdftzMJYfNfGdMoGhZMbjqrGzGYA50GGvEsgXJ3jseUFXmlvK
1xGFqH+B1CocRhBfje0jMEDjgeMfZVjYIaI5w4DSGS5pS22kZtd+93Eb/jRMPt2a
8D6iAdyXWCYzqicku+3ymQ5mG7gRreJaSy5n0eNa0crv8skwPZlecR6Ht4nkguxN
mvS/efLA0JXdoU1zDEO+hXJmNCG+KQI9G9DrQubQgx3ifMnMPH3voGM8no1Lr203
uvE3NvC6Eu7dWKlxrAG0haXZj1uhvgQ/HnxBnfd1ksAdmsZdUTIgLxd/QpDVJmgj
VYrlUbNGFDqWEYMnsR9ASX5BybC3RUyEXMmwBa17Dipre7ucB0kM0JslxIkCKzoV
DIn6AludMTRuA/SX10I3v6/HbXA8GEgiRu4WaBe5mSuY2G+TjO2DRv8JG2ngs1d7
krJAt0rHUfo+tUU5R1v6Fw21q1Fc1PB+AHGyLfy/JS36bfn68MhStBlE09qR9XPt
/GByGH+XIn8l8AK0KXDIBgfcisnvXnoBV8A65a+MsVsnVSAt7+Z9zWF1AjMmX7ll
4FC1tY7bdYnlcJjzykbVZfOH/6tDs7HrX92q+X3vQUtSBMHDr6D7FA156rR8gDma
9Ago/CjyFPHbbjqZvOyBkyupc+31EJDljnTnPqs6A8tyKWZDUdYjEPCtnmS3WUp8
NYpcleOAfCon7+jzpC9zx28+C9AijsgKOR2AQQ5y5iSEIlEJGIWHQXNgQ6IeZ5xW
AtC8fvjFTy/29RX+BoS7Ih25UzmpBQmpgQOSiSpY3vCX2xLCFlvq/+CkND33O0vg
o7Xql/vtTHxiUgwIHjxv1Y7H8aXTgxVVpwhNhnCH7uEW/4BY6y9XlsOG+j9RUW9w
tDFkQQSXCNl9/EL9rdos9okXs44oqmf4zPuXGF0aXbeLbNJ8SX1/Fst76+PH8tFc
sn/ilu+ajJtsAsbPlXRn3mFJlVPYbBDOU21W8w11wC9UicbQ/3j8QBolEFDo9fxA
R2g0yohNPL2HY+ZMT+0OIk3my4LZf/9pU2j6UXK/z2pzKy+A2pf6d0L0OMhSCp6N
64eE+5xuqtr43erq0JleHlMI7uPCMIENrjab82QXR3uH+9Wjm5nU+k3Ys3l3Jmoz
kA22oXJ1icjiNOosmR0K0phIKsS4qM4/f/yP54Z745HqBM+dJx2pVQNyDNactnBz
NfsPw78pqu1ljp/z6fREZs1khTSDBOTZBdzIFvW1gFdMmBeWM57YU81feTLL/JoB
sp3ZUUp2HOl1GrNTqxd6NkXit78XSJp7FbX5ErLrWH9zRc89xPZ7P9jyXhBcqUHj
3BeXhGwReFCeM/n12oieHrLX5dCLA8u0dxVur8S30MN1AI6G/mCmgkLhh5lLqNSH
1fiIG6FcNrEuHrWjDGOYah2uioXu83QDFSfAwIyNEQjIFbsKdllH0f9c1GjpO3Go
Tml2s4fL9C/d0UelEG7MS5XHbjKdg2wjykGhBhEZWdw9ZAItcGIcSPUIC4C6qHj4
c/2uh6mE/xrzPHWeD/AfgNo4y+yMqz71ev1vzSHM/DSZMUf0FszG4Pqus4hKLBLH
p3O+ITPFUGs8NnTLRx0DmpY7AHSb1AmOG0r8BLmo1JJiRYE9h/HE3iAy2H7nt5Fd
snGmaYZiDvd8ZaRbqqAADaNeILsZkxnLWjHKBKWAX1wYLNed9VLiv8TLvPg4bt9c
T4VxsV6cJ5Xkl9nmfJcLmVBmg5/1ZJhYRWVfywzrCts5Yhic343PnIEdwTGEH22R
Y51ZZgcxNyl1jYAeynPzcGk/WFNyb+GtT1A+Iiob9Fd1nMAJAdu+NYGzbqWT2XXJ
Mv456R59q8B0nkf1pXZ354uNJ4uJQm5ZDZq1NBy9zWD9XfeDClYA55xGsIZrbFzM
2YoqbdPAaX4kMoBlSsm67P6FHtdSLdWpozXAiJto60i4RlW4/aKPx5/3fubN4cz+
xLbWGU6yXyr9wNcCmeQ7Rz8Z6jYxLDLmA/Y8LTuCZXqiga9gb1smb88uLCAuUwgz
JpZmIiFtDyZmxW3SUPVZBFHzzCa31MLNju4ibD78bMi73CFEfoZ3j6VmobdnHXsK
GYryRpz3BXwJb7ipRfLiAFKEv2Hip+9l4LzZ0X2GyKlwx8ZCRiYV89p+48Xz3oYG
2AH3+LvxuI8PlQq92QBrxjZuHDVaA5OZVAm1OWdiHHJj58p96L+u9iZLtth4VR3k
H1Q/uDfs95RhLy1K5V7R+DJOu2SZ0kEnyVmnHjyFf57bG02nNfm55rIl4RrGExxG
5o656aGqNSmK1/bj9AKRcJkyfYq+cLFdIZrIMJLNcMgES+wrP94GSRvgNq0Lbiwa
qsJC1w0Brvmb9OYFs62Zavl+ofjP8z7G+/YQj+HmoWVIO1qeSxQm4OiRPgvobmX2
PrGg4ntJXx5mk7/UvXh6fLA2EqQsDM3fXqAgFj5rVG4upBWL8QF7YcuvXzY2f8/k
oolLT3hj6wLKLfi23cKn+/xqSIobJfIbfA59tYeiNWc6N9xkvMasqfhJLpv0SG61
ZVER+oDqPUUkz73A5nlZAD40SXkEmLxpizyK+MeSvKMRpgoNb93gq1+U1XtQ63+o
c3dYvUNDzIVq//+Fn/HN9ZvLrMiiaLn3Hmo1I3JSe+Pq3/ao6dw/xT/cpV3ERsY6
qWVirRqGXoVYHZmPOppQcLNo50JqhPWC40JxaKJbrE9k7BDiYS2uRWbMlhQaPwZN
BlWKTeZ0LGLs6QjhBxH7anfJxBL3FCkcWqQbfDXUwASq3ol2a8wIG0Hml1GS3tbi
Rmeu6MBG4a63WvpFvRt+TjRfLFAto+2xcN8PbdCm4hqO9DlzCABn8OUGiAUjvGMR
AM+zWAsX5yxxndvN16UcU0uIvxU4Lb+kd+ATXWv2HU9G1/S4T7/c7CPVB7gMol7+
M1uX4K/OPXuKKBkn6G943w6XXyseW3IlJtXttax6tB56BcAB83nz10dFsl0U2SW7
C8unuDdxvLgLLQlfKB2FWH+2VHF3vyYdJDwSD5RH9/eZWSV9B13IP8CGHoyxltBM
YvgtwlhwKgPEtPTt00dWXKuozrAQSuwuMfys/BdLKnDbAQCQjvchoHnOi6Ed7jC8
jg0HBrE56ZZQkishwhgvMF1+jrAZ2CXfUBxufkYxQeG3jaNxflpO0RJeV8VXwlYF
QejDfkwcdM3tKuMkQ2FI7gkvhipoKZJ6T96gWcVKRgM7Ck39YxZeFDuu5PE8aA6m
971twszGEq5aEODqbvAQc1lwoTGjHh/1K2MwOSC+TgJdcXzEqSFnpGlHbWMfiD3L
bL2GVp6sLAvX6eRpoNpH5OZjNzndcnjacjOpBAG17KbWVEmWrN3kyYUhB+RsTE3N
pHm0J3Wjva/uyU9RzL9/xuV741/0H09JaEZQ4HIpGFRF8atBt2fZympKP0oyKcNw
A66NCr++Qyj17UJQPhOLTAnb+99oujozyrZK8aLw4ZTfSPft3MfCXYerfAca8qgt
3Me7gS3z6qn0G5IEuhw1JjWz4b5SZGun1G9+6H+EvGcoOfNaIcAOdpDyDxIMidTu
+FqTC1oTXKfyDfoKIEg6d5cbBnZJhXx1Z/M0RulzBsaOGQDMcFSpr2YbjpgtXdTs
p2LmtHKEXVA45FyWXSMxVpUQSgYVaj5Mfbmf9XYD7nQKqGYLkcmg8jF/IsPDqquf
5mPcqUwzU3KQsiUjbVXN7H2pGUi2D+uulkFPmdEMIZ3t5l0TWXs6JQQE4jboHowi
taQWuH30i0wH+UHanepInc50hOlepdJazIujRD0g15Z1vrL3hEkh7mUQm2tvaWD1
JHbC2Di9XT6wguslkXtBPqxXzT9MYZuab/Q+b7xcMNYZ2G8UkNewjYilnAssGrX3
8UEvUz55mNgGLaMeGPwo4O2hbulj4PWymDj8LiZpRKNQOdvnH23WAt/hHs7uieYC
or8Pw6EPPzX4HPakHn1s9nXKuXfdWjv1j2Y73c2QHBBhpZMDbWLXz3Y7PgYXP31N
Qa+xwttYcdSyftF+36RO4xU6YrdyjwEFRuumwMIollx2sWjKDBc1/7m4qBIcIKlZ
5oKk3SlzFnZdNVD3MO9PQA5u1lVlk3oJLjYrEcqP/Jvj3CmRv1jQKN2UjFiGH8IK
gPllzTFS47H9arrq5O8zlqxVClU8u/qRIdj1LOs/81HC/vhyAaC2MYyCqypmQpjl
zmHeCkELln1sQV97FYln9UIzI4oOeIdybDfnUSgYY9vqNVKg5Z2U0oJ25n85ghX+
voR1g79Yg64VoGiJYqhBwDprppyrJy6pKRb3t4vV1C9F7Cs5COa9EmNto0IiU6cB
NG/0P1FlnCTGnixFVLAGC6p6U3RuaLxkJ6bl9+ik6qxFMmCEA6pgNS/YGxCTQ6nG
kwNJ/EZMMwNUdhiQa5/X4pQJyc1m06wE7p0n7HXNnT43V90BJ4f2GEnik/lnHkB+
Js4qcQMNkb9fvBJzQpbwLCdvuaEvb9T3xIRgmAqrtr3k73Z3/6VzmxF9pR2SIxEM
ov67Mx9rcP16J7ZAL2umlTxP4vPxGhVGDMIUCd5KB2ZlWLObBg4XQ50ajNrWmi6y
ycCpUsjw3r6rfDpc230Gz93Tu7QbwC8XCiK6WwDtKRuWnnpnFXOEOixWG/kQsOFA
yxmaq/FDO1g5enak+vvQHX0ixe+8oxH0uqvl5JcpNrFNleG4YjjatO0UZi8kz4cA
Rl/A8ywhlCeqn+XX3G423KnjNnykQk97FO69BtYqr9ZeVCXukCKS5lPckHfw2pOe
elqKWGIuda9KzL464g33D+IcoNtGdzXQWqTM7M4iy1VSeCJ4bluJ9Hft4O4cUqiM
4A39TKnaJMKQvWVzkqYnQ+pxYsNBVeZlGCY98jpgAv4O+2NmWoZgNe3t5ETwFLlI
6DcxbC7ocELpvNSbPmRpI38OQDva8JYQQzD1eoDjXE3GKsan5e/RpGRypaQz/qTJ
zRlq7eoRa1+89lDwNztE+pwYwYsFNDdoKAWg/mYjfwv9Bk4HP36BCl2XoxPa46yi
GxtmjJL+hdN7zTJaEJMtXEzUuEGOp7Awn87ttiOv1julSvhinWazhtliHvMbyMm7
Ah+6YEo9MX6rU50PGMeWGKo26W80zrfVQEuiHIb67wsbE/x/RVHqQqUp/butBcCF
dCFOa4xplQZFLMdBPhFR/EObCAA9o9ZxZaWWwIoGIxth17SQp0xdzfr9HvaUY98+
pDuSdLX33rqSQntwD8Ayjqw68CR2TrtqqMSMGAtKBk9Wir+i5PtU70BL4I9SjU4C
JU1CJwQLOPN56e/BMMHxA7TjM2wMabTiqhHkRljFnQQCYg0m1BDnC7DCSlBiP9Qu
5FYzVIAgoTAgUlYcxlL9bfl5qDu61pRdX2Jif0aOrlBXnvTfix9eNKNKa/fb4Oo/
/+yIrr3aRYZnNRBf+QeQb7No5SHZhDQu3nvsNyFoT4D9wCLL0r2iyEFEOyhqcvrn
cJ5vJz2CA3MvgRvNAHsfDG6QnxM8d2wj3JGvjyjsM6KbdnUbNBGvsTLtjYyOXa6I
mep5FimtP2WzkO1YTp97Wpx1bpPD07oCHOxshkSqssgQfUp14u/mvQ7u/v5sIeGX
fRhe6YgnEnLNQ9PqRSXuibXZPeU5RA6KYL/jD5lL0v7F4Oy/SYgavX+uyEt83qvI
xgboR5bMKHDOsFxrG/EBzUxrhLJ9bdCSJVAdNlInMZjgyWWKRDcGnmDH924FLPOO
quH4N23ZYsS5XbTcItjaDb+he351bZ3lKl7MmgH+h8mmzB4PeoDRjyKnbf2YHOqo
eJIaqGUMVl6t0CoSmKbTn+vd3lfK6P1iNjlMKDenSdgSTcS8Bpx1jt5L7H9Powk/
76E7XyHeHE3IboV4n2QI5704LTA7c0BP7BaeQXiipFQ/t+Mq81Srv0kl/CvL09qw
H8K7H4O8P8PcDzLe6BWZSi0LOu8lJAa20j7Srbrl7mDdTIjto2RecF3dvJwqyx/c
qoXuEJxcDEljgmTSZfXYzsKpT+vIWOuNk1rEEZ23JGu7AKvyNPKew0HIuTr8WeRS
BtLsOWGYb+ts0hAYI3lg4LYxOnpu3Z9GliX4ACYidKUnkBUIqE5PkqWkzZmOu3oB
39CsjmlcISiZFuRwgQHMJB0IoIRAe2x245jTf+xG65NoDwiNxXQxzDeW5QOPSXPD
kmhreMrfOd+GNiEYAr2xW4HZjw+Mz1gEOtiZpcfAJxcOTEqSovxupzXHq4cK6BrS
QM8an4CzOHQ7yi/8BBPAF2NLYA8YWmWcqPDJS2p+wC8ahkM9WlUiw+v8IiwV9Saa
hwcQ4/5mZpvc2ygQWAirwNFUjuWm1GSnGe4TzPX33Kkp14neyb+q62KkYAuOfzRC
gkqwhLt7JYbYAcG7rUwz62t4l3+YIi4mwEtB3OHfdVIQN9tYg0B4oLb2rWyTMQix
qYHE1m4dcngjHj2bPNgB67ahwkcg3fPazfxRJogiLU2JA/WbCPDjxlPjTCC4WJzK
8wvS/0+5jRCDhsrWMp3JaeMwhDCpxmdzGco1u7MJ3jiMaU3DEsSyXODCPKSKHuO5
DT1bX77qKpB+BqwHO89lVJZvFU1vxxwCUvr/xiILkp8WRmruvLzml4g12EUwtdC0
ud/+ixp4qUbs5/+QG3buJVqWBv2kRGTtUnpkgYDab4b78MJOTioqq6WJZVlbGpL9
1mUNlg3l36LH411HIoYtRtKHnpad8FrWBrKgt8HH9KAlhM2ViJbOh5ueOG/x4aMi
IJyyUbi4Wa02KfKMTosvxhmB91H+hX0jNNVS7aiXOuMuWmB3PgJuTVR8ERzKuOei
KLj1GHYqWJ4Bxi9UteH+tqr7Ov3d4GLc4+T+B0T6Uibhu5sZc1Igx7G6hv/voz3w
oMxDRhqqYiiPzczIkJrViRR3RIzRSJ/52hyzbzFvrm8MmHpk+OdcZAB1w0SmZkg/
A9ytrAyNT7gzk/kOthNmVqZLhLB2heRB308Jz5BQ7XIzSoW8yP9JC7FUat0mJTcY
cEbr9M6hHRLrn1t2s2RLSwPN3cxb0KMC84mHdFksYsBVhR1dIEOiXR5xumeFkHyj
AbS7cC1hCbqsIy3UQTf0TIUfSZT7Xj+dAags816AgEsWFu8H7Wx2gr6zx0nUAEok
3HMtyn6LkMRILuasn2hK8ea7c5SqhpRV0Y0ynsdLn5SktdmpHSu675qSo7YxWEc/
yrr09hNkNAcCCvg2TwUshVfVQjW3baE0oDs9k8TcoeartLK3ly/gmlzByR84Y+Ab
UUaqOrQeYDbtYmQj5v8OY+LsJCuzw0TgMcZkgEaYnGZu7qRk0BvUVSLR7WPS1Tb2
vlOknJrXtEDAXZMjcSMmfA75CnEcy+vxGL9u1BiNYjHzKiwbsSeoNcru4eFmNKdB
wl5dEm/WyWEBKJmFtWb7Hz1NZJBUb263MydeUEpOlwZXUmJfOJdo7QxM/Hlq9jIJ
YVlJkYfAwg/gTz/qjYPbgHwhW6tEGtt+gJjOy9llpHD9EDPnxQb1DmDz4fUzF5+O
GHLi7E7+OjpWrsgrBSDNGEuAvBjU6bcaSymswzTZXUUkfTsZS3ZJk1pMAVmOOZpk
hbIX1idZy2u525mD/kp4qzupWUmYP1ySl3SpHC1Ok8JXZp5IAvQwU2u3md3R6+SG
oi9DF6V3lVFtqHe4kA53RGBiIW1VFbW5sKvfqv1Gwp5bI1WWjXx0A/M/L69TbHS1
63k9V9g+gLSnqEMmh9HwOfbz8lMSDOtVE9LW3I2RkSoJgHXMbm+VLcMM+38OAKeB
Z6ZVkcTOtV2SfpR0vPZ6JPxyNHtiLcP0vBWsqKrkn9M4JzMYhJ42dVDLy2ZVFXf0
pFUFtYlekICZny7SU1qGX2JPVcPslZsHxH+wV066XMWcyIr+q+BXpDJxYSA7OkAV
D3DkrByd2R42iMawYPlDXFCQNHeIoH3vwlBnXXYGURAPL+Qd81nf3tdCbiNS5UjQ
l4+XDfugJR0yr/CzyjbdIilxcPbNfgy8Hw7l86guotJmY0CJgO/2Oi6ze6/8nujl
i17wAelpO9CbCoS6+a/vEkZe07OvADQryvhHN0kAFjhCDbiwx+XxORkuyzlyYC8X
PRyCscBz/NgDUbfQD0w1LHNTFFGTpCI54U8yA7wOfNPxmiJ4H75fmM+Czmarp5hQ
F0d0o4bDbfUvecVFFon3It7oIiFC/dGI4BJWv9XNue7zYYridSv1EJRs0QXcsu0W
19FTuI8orftokQIfTS+XfXAWU6F/WIhSg1ZQGeZB7HLy+CMKWOyHLiufS3pm2gKL
fmtVUHB14lfj5utDG/BbQ5H1Q0VH21zdFQ5yvJcVnmPy7HeYBe0V7h9Beeln1/dK
/T5b95ca6/Ti/MTqD4UzRNjCAcIalYaQ+jKSrsuBHIns0LKwXZuVkCwWryx/D5Ym
YUsHaWCCoHAlIXTLcecUOVYAhaJNI2F97agePLbAy9v9yYvbwDeclQAeJ9+xS1z0
A63wc3STwVHFGX91+V/NN0J/57jlNGnR7f46a9+wGCTY8Uqyqcwg0ICvDFg5NBUZ
yB9tJHCyQvPUTsxxg91EdlNwgr2E07K+Bqr8Wdg2LgOnzpmcF2rMBTqjJaDDSTtd
TtQd6NColx9BoloAqjp6KhvH0vdGLlcm0OnW3J0PUlJA4ZUjCUmiUG6WRCAs8Kgo
ct/XJvo3fDtFsEf+xNmnDdQtBeq1a+0qLBMwwMzQojwWATlUSwxtDWxU5EgqSxTm
NUHnpq/MmL6hEh46KjYNNDkQ8cTh6xXmmiKL87l2S0dzZLehiC1Nbv8uKhpikmos
tr8yOAQHlwXpnxEVmCIGvtkqiqA3wvXGnrGeEhIdsWD3a3jtQwtZSnCqd0WGooiA
8Wi29S4KxyXpBpXJcr1oNfXyZkhnVN/ZGOc+6wOFJZqNc7z/Lm8dthOqvzdBZ5RW
ZnzhuxZx5UZtyIidFBGOM999r/g6hXr3fLOo7kJLy4DwT8h7zP/6LXSrLgsQPa/Z
jNlu92F4IwUvbyOG4+9x0tEwOu8ajVlgMonX7cT1R6GA0hEDkNZ97YZiuKdf0+pN
AUv57UtCZWxPqsR2FP28/cmzBmAh4U/8IKrQ1Nw+45sQp7Blnv0ZavXylhNGGNxh
rCesyJyoz7UqTor9RrXxH1Kqe2GIZhe1r/TfiHK3+MRLxuZNNeBPbUbP/yEh9OxQ
gNUZlhSn0lkoTPZKKC7cHQqLd+UdWHUWq+CDgvUNnlWJdiBiU9nJczD56BQcN4Eq
vNXV9Gl/qe2oqctt1/NF2GU1uP4DnIxPuk0htxc8sybalb3BfiwDJrJyjSK7WV/P
ykEPXJxiE5MaEI5fR3ZAVWa1xNj/SpIUOki4fOwqaoMBYVEL+QgOPAmoiYid4rJX
UCTpulD1YhAPdUQAarpRSY9hRS7REzYlbEXBrFl6jOsvoGhhW90ydk+Ialbffj4C
rBkMt1/YnAyrbWDV9T95C6fCUj8ye7eVz7S5d9aAtS38P52YAw5U4HQSjKmbhwad
No9sHKCZUbdsx2AGUKBqgkmS/+sylLzjU3M7ExKEXO3J8a1mygXcE5ilZu8NoUk0
QsZudEX+MWKg5rDrn2Xmkx/5NF14Ser1jiallOA+/ALgASKFXBJ1JP9jqxXGZtEW
rg8cy15+puw5sEEf5Eql54anBipKH8iBZhoZJAn4ELvH/iWFnQyr7aeDXrooB/zG
HmCQ/H8geRJQGqN8z3YrGvb74XnaW7KH1sUpWJrJLW1cLUtj5MT5LSUGW1lT8fF2
h9XyOrcj1ZrpDhrxzVJrzp9nfO3a4eHYtLCtIYeu81sIMS0mwleMW0f6IyABIqTR
KLrLnirzE2Z/W68ELS78HxEnr80vQEJ616Aq6RI26F642qC8Dk6+jUGr4pVEIpXe
mjQzs/P4Zgvaz8bX69ZFLUacVED2bliuY7LpR97jPOBwTHFkaPp7wFTbl3rtV/u6
b0JmaLsBQ/5eL04JUZ5kFZA3KDRr7gbKhqcPavZT9I+pNs9HuTT4lQCQYW07kAiK
1gdpVYsJiQXMHshq1hRPehHEu0lRqXGlIfZHT7352toiq5NIu6giqjWGZNgsHBtJ
I2vtbpldl97vxA8f/D1Ch41QGIpmd2fPQXT2c1EXTDXtsl0la2oJapfTsW745NZN
HxSDydSqUrXb6xS/jwS5sR3LRjXJXRQvfxkdvXpL/9f+Y0YLIq0O2IbmAB3PWtt+
T7SJ6964LD8opIHwHIWVuTAKHGAiSVbHssAWoXELiY8pDTf1e42HMLpQnrQ9mcXA
+aFqkSfmflL+QK441Hh1IrE9IxifbDc+1s/gb3YSPxiT9y2xWvt80egGX1hMUmQl
GfAwSb6DJEDyHZGsyLuKxop2XuK81vxTGhT+Y6MWoTBSH7P6qDQ9IcvGQjVhMcEI
tbB+ClPZO2eg1lIEuPX8S/873GCzurrwfiGEzA6EUEON4RyKj4VT2NxWcrUanuOr
J0nJfZwmtpr3fSq8X83NWOUPaEubKusqWwnHSNgmO3xE4oP9D7K6LrPpUcAsne66
EH2byzhxUz/NtNNd3KJ3TME653JHffqYUuIRIgM3DPFItheSo6weIfkscvm5L1h3
6KXE+tMcOs9f9aCrYUTpxHUTe6oNpLuL1y6pYqOJU2sicPLkhyfQbCWezffuUfEb
kxrz/Z2qrvGIL6LsrvjA22x2K1J8dLDba2/Cu129vUfGdR0mcem7PeFyI0qhsDEQ
TKK7GAEcJrXvfdI/am2U1HuHOOnmZVAcHC6YXmwFvtsX6y5EBebPEVUlJekPsnYO
Mczmj6jA+wYcUEVIgU8m3N0wguSy7mMAE9+6jB6J5JCQgeTwhriaaCF1MhWDztFC
Igw+EZOyM+YtgZdtrZe0xT46Z0J4Ls0d2dlQ5WHaiWiRLUAao0TdptwVa2RTBGcf
lIE2AHRjkZ/FFi2N/0wv2P+mIukrYgzFxDVYZ7gZVOO8eDQ6vpvTl7T4eRAl9EzW
GXMxbiz3+H31bkMgDOciWhcryHb7KHCoJgN0c/HpTG7Asi9+xe9SQsiCwZGFE74w
kTOtdbV1yj8/0NHLbsC3ewmqUAziw8OeQRnCV+g5Fy2ovcjJqobDVSK42KY9ojvf
gOo/mHFv3Mh9GZ0ssmTnKyiwSS8MCcoLOBEWKKiHU4Z9qsa/I/brSO/VQyNm18xt
h2/sSmr+XdD7tBTfNh4txxaq/2CqgQH6FqogeDJHwhMm6pc5qNMLVAoKqXC5sceW
w3RcNd2t/oLomjXpVLiBgA77I5bBkrHtiWyeVj7CkvWCMWJ5vY8Oi++Ns0vvFqpe
0PGQcSB29cHc4PtHrHuTW2Lrzv5pVMHvoP3jd2cmn5XHAjjUc7lHUEfGrvwmUR6w
g90YXWJUzM09S7D2Rqof2ExH/GBCHK7ciYDHmj4HINUbXiBWNk+0SIxWcjRzPuuu
GeoF/tEbzlQCjmJ6r+lT+Y5z//I8G5R5vLZ7Thh+nxslkMatoiAcuZ1U6VTScR/g
MQUMykC2FSY7UX7mdpHWJ2ybMsactrPljG20HA4MpiiZSpStVTIOqBYf2bMc0qJK
e0uoCwGhpT95GcKVJfK4SRYUDuUby+tr/pIuGkv18nsmgizQplJLk7IdklkerdV1
2MiY7J2E0Mss++A1rsvzKutyMxZTfMLc0lrMR3efG8LSqwnjQXFHlrI0zOhr+jYZ
rHQ6BNhwCyMbQm3XwQDqWnusd1y/T+Mn8s7R+0tchXeMIug48qcVbXX1XhJXRi7X
29+IHS+xK7KAQ0uFmIACk9cC71RT1v6Mbozp9Y0lPC6yMuZuaWIbLUzfYq9mEwXq
V5cOqwZR/z1Li0cflffNX75AZ5IjXAorpzOzsAp7+q44DxPdyVjllgVt4+Ch8JM0
yvtBJPu3136JC767dOECvJjHLegsxmO+YfOjPsVynLgtRusBG2VbTQkUg73bBLTX
xdiXjnRhGFgews2lyx7pPkA0AIWZc7D41EKpECyTfBTo9d7A2viARQzRHErGX5AM
iWo2Eu0mitrhjEVx1xMMPxMIDta0J0kA9ScMYGkylu5tjIcMpxLipx/VebtvMt4O
99klZPbvETlp/s9fK26WTWEWLRzAKSsBcSsAwR6vHRKRcaxrQpnjBKR0OhxcxPNv
nmPUlM9vMuibcZZorIoNNlLUAATJgFr7nsDsOGAymSzTG+/eLJQ3TcyxWVrYzXYO
o38bsc25lu/urzEFW+oKu8mThVx8pbFULD7l0MZUyBkSandHxbjODAbHKrXJNZUX
Rg5Mn8KjxcSsRP+i2MJu/DgcFcPNxEQE1PkJdejM+d3BopBFUAmSBBme6tSY7Lcg
qy2PtiUUU+aLXIBNuW/Dj+r3XQRHFq1FZ1izrtlt1Uv+xKzrYE4XwwxqMClTQ6nO
WA+x+8J+LZRAsna633xo61eJy2YgkD5U2VnUfTyg6IkvHWVegxXMblbIVLFb5DPH
jwapqL0yAUuff8dvVLVP0U3H97Qlz+C//e8ypRZIEtsuxszOZnyt1tuhFamTLydd
af7dAElWLfaUyQ7tofMnETJWok8gKyxLFag1Pbdove+o/QiihXAJ1xH/Tc1q8Em1
Dt17UHSKsC5q4FSDDAg/KqA/Ml76iMOhzumEiQL1O/UGna2mfLOWHUPEDLRWtW0C
rFQsLUlPRT5jqcNJQvdm29zRV1DEkVRiIeW5eBW2mw+MaG9OiIeyeuqBB9q+Zq+W
yWGov5iK2+FZJcTtU8pMzSf3y06SJP/hx2uJ8AFnIJhUr17wuxYZHdjTP9Pnbj27
np1WasxhAAYZZfgzTXfxZaF92+xbX68YAPg7SLk1m+d5eogh8Zga6lLpCsWAnRak
bLhFiWDDkjbcmElBfTzPP010enq+WMMbmaW0P1NwkvgHmP+4oho6vw5fLws2PJqj
W0I2RRq3bG2yW1bqmJcxhZULxxLiK7QTS2SvEjMQN89lBGvnHnyG+XRVCdMX9ag+
N3+pJ+IX1/uGhWkS4eW1JgVCAeC6OlM91fSfKdyiNTWXyDyZQS/RW2SYwqgiQv79
Wh/im0F+wXnvUzHHzcXBOhwCr3ZuztYLOsL/jysyaG8MR4VBsuY+/vhN33PePuCf
z0sfin9CA7mjPS/xK/oobMy2d/y/vp7ZeR/4XOEKjWDvm+oLAVZL/XyAbit7HriP
Ki6ASRueHAK2lkxfTAaDU+ssaHDHjg+i2NnF6GKm9zW7hgq8nJZ5Qp0pFhdwSnqU
C0n2UKzcWNdq91miJxR/VozNZ0Dg9jFaV13n/5Xkud+OottdCz4CbLf0X6u+mvdA
lc9RgF34dTZCnm1QwGv9VEUAJtR/BZmjC227xEBzVb+dowmuRyG/Bpg4Q+56oKYE
a9EkngSJVXv4tAGQy20QCgjjXeV+NzU/radFzeYk9XgHwxRfGBndZxWQ4pL/MrFS
jwUrT///9sSrBdIP0GxXhg+VjWPUZ9PX4OGoh5OUjeh51+QtOP8IKDle7hyKL+6p
LjnUqNmB/pvTY6CPK2DcqYiGAS9hRZafjVqdmPqnK956yC5+/kdKWqh/QkDIO0O7
8A0nsdQavFqesF/Huf9CdEInw24J8IfFmgCHUN500nRBQD/k6G+xcOVFqNysZWPD
SbrHmSKM9P40tz81wnQk7nbM8utCKiKgEZa94kdKaA0cL3dI3XA0PODo2rz1YGcb
vTN8wYNsRiqisNW7l+Nbxe7y814pSVhDWDdAJmBql6XH+rrSNl9NMNv+rBXW0jLJ
Rz9aUg1J82koFXtEfw3ZJN6UOFvUrxkqC0O7dzUq4IjQ93fe6GLukKA04m0CYvWW
jhXrPWObEc/ui3TBgAMG2AgXhzyQn8tS90gl96oDVTiZpLQ++8JpBZbWiqMwMfPt
Bt+IUJyZANbh1QHdQ5uXDAYcYWJVRtmav2X2pkAfLBBPMauTZkVJTt111avZ+7x7
E254ZZY2OWXGFRW1HnuZs8SYQ4uc4eBBIuw7l2lnl0OmIoz9eQ1HizKZwen0t+Zw
nJVjjMXfmTJgy67z15d+dpZJ9DSijMEmt70oePp9plvFKtja85GU5XZkG5spZRX3
jiq6oa4OuCyxxdzi/rOqeeKhUJnxLxHk2nEOVFedh59s9x6OTd6jN7eojbCRwZOu
FCvTquVSLPeRJoetngX+TyUg4HOE3HoHYwMORvymcRI4tZa8+PrhfRYNXMnLdTGs
7D9pLV29CUvY+yUD1graNjikRjNL6BUg3dVrRPPpdOhpbVdnWVBKfb70bnQ/gZc+
wJOxNukpgEzC4A/3xpeJq2W/A7KzAMMpbhD/pu9XBZzCqXGjjtLQ+UnmPBsyv5kn
uVXGG0Ys0q3k/GFaL4Q1FC512/UBVhha+isDIYZTs+ejVHSDkjAEmziK5K47cUiD
P5s3XRVTuslKDfwjVBklnAAcOXqa9odkCj/kDcoSVPBIAMLJ63jXb6erzsB2F6AO
GsP6UftYpuB4XWGyi18mTTbfoSe1BN4uN+8JXdKDZKyvMEBYumj44KH/L0OXirj4
G7SRlT4rN4JIvkHPBr1B+O2zgjhKGbj2hiAyPk8oVSQw/0eKH6p6yK5EZxxUIpQT
e6eeERG6Siqwoi0z91KaIVpxAhIdDP2BGFORzmBtYTkOgQN2Iw+HHxfl6AvoH4uk
6bWhwEWlyWHS21tks+D6Y3pnxYPasrz4ONFg5hEblwl2/V0XsgFvdr4vGgaR6okQ
ZXmYNby5xqPmKIQxlipmrdQAOgQKs9JU9OQcJE/zyWkXplEgFN9YyL5Wz+3BTlCZ
ez8eUHnyG/c6RiHNkOo5EMTNj3Si6FGl44vTExN3wfDIKRkwJXKSXS9Agh1My5vx
H2jS1Cff2MofwYF9IufF+U9Lk6cDVn7gbKMZrVAbrlu2IUKr8YPGgBGPl/Z9gEM4
nnR9hAckPvIAT8VA6+JcLvaLruK3q5qaHChW/ArfR9IY0hTcof5GsV9FRtUB01mG
535PUzNJVoMVQUlHZ8u2I2aKyL/YC5g9myr5Doe52urHU2ASB7ibKOPRz0FC2Tnm
pBSNUG9Ye3D1cx21AmlIJic3lK7dv2UKxCvSvg9vcHz21C2Mlcoir+HmKZKxHp7D
brH4aVr82iXn8erw22cZQk/dXN1O2PaA3tVaCyx8u17Jnk+3hNkLKN8LKo1c128C
H5UbxDc8R3zAgcgcfOnXn1UiSyY4WfI6mgmX2HTyVwsnKL4tXzDCW9XKbth9hh7d
t/eoDrXmgAQqTwlBb3k6O8ZPY2bFJ9LuY+F0DYJPuEi8lkcNZRKbNhyCakXpn26d
lMvl+LkGGgJI1hjONSXTCNbJoBCVVn63nHFjwj4raxCy6Rk7RWw6CAQvstfsEX/U
MUw23Gb18iyKWOAV1OWKu15wL6K3caISptVUbj7IH7VlnWxHReM4aesND9MuA/FO
y1w9mukNx+mfGJvd5D1lPTdQh6WLQPx9HQRg9ugjBKrZmlVU0Kcbj7oDP97s24aN
EZV7H1U/wxBpiiQTWNAvcHCmitQeTYQoSoYnJC1ih5lhEX+tb5z6evveNTw2xbZ5
ZS3j3cNYglUH1LILiguLwsotsZjmE1wzqIjVnJ/ZvijE2qMFE4sQt4lLTuhuVsYh
8FDvZdBSDRmw/tIZ61JY7x6dmjZEo1S5z2BIVOaCjc9LJkJ71HedAyuDHCreqLFD
ixJF06COY7KT8yy3oQxXPIPOB96xjpycFQUfqMV9dOx8thxGIE2ewYW3H0UPWInM
tuxqHiFKoBjBslEYLExBNT9M84doePx4CB5B99S8qPJV1vm0VmYFgxqYjKf8jlj3
A1ETIcMFoN63bVs0XvSLlmU6cNisAzrzepanaOcF6OeYaky3J4jZtI2skA7kwmwC
Dnu4k+E3s+8MIzeAohXjp8PVi7OCQxPWDlResIEMNsWS1lRsGtRvh1fhoHLlFMsI
uIA9xvh1GYjmsOsAjVUAfVC0rdJg2V6VErba0OJPgrgm1xu2ePxx/Sz5hZQbykUc
M3VKT6Lo8RV9stlfymLUW+xfJb9LKYZnPsyAK79ZGSOpSzxff46e/rfOuCOQi9p7
6FzV/kO3CdY2DDWPqG20TTNyX1KFiZB7YwS2UPYyxgWl4nxeSmwGARyXsGon0FS5
u1wA8fadHfHT7C+oECpnPxccxxTETw5+3fIuUPw+qQi+Lq0+ydZks+hWJ8T3/8ah
/8LThHb7jzLnmOfGpATbiR6M5mH6rX4whdilcL27RJfwcvuN+TUUYbsfEYFww5C6
OiVwpSqZlKSrAePMEBPlNc1QT9NImcP6P6m/onSz854ET8ckgW2rCImJNq6UjpXv
uxU7ZyeDIzqaCV36D9YoNgctvcFINXyyZtYT85oVKKvJZnF0qqYbd3vHed8rYTMV
crQMFJxeC78qnP6y+zqCiyBjCqczUB3CFUzEFcvTAfePWXmCkOLRhOBCvQDxCc9s
uN9ozKqNB3phOv+REuhPkHrTKCniCOVVKZiTqPiGYkEUWXZETEerX6gcFGvJQ5Ed
HZGUpXhX94Bj67eyC36J6Z8q7ycAwtVwE5PVd3Ssjg0kKY6uu/9vWDZc/xAVIapY
8bsm1yHyqsGT8T+rAaa0in2ZDl+IQaUT6eCmUg2/HUzosf5bN7vhmn0/raoIKQgl
Nqly+QOY2vT9RGOehiRPgr5zKipZDZ7OVOVhzDKo3PG+kMxv3FyIpWuJGMRu28ZS
uiUoqWMp0qJaXlXYcvUqA/hyrk7r20Ttlvg7huGcf/aolBK2doYFLIZr18yRE1HG
9Og/J2N/U2QkF23FyfTa2pQ2BJer8BcW/TQNRjnSizDvic0D+Twq5HOlmvNBiP8u
+jVJdpoWrq7dnQYw2TPt4XLy1KqCcEium6QwyEScWZDKWfJHpAp+7QEd7Ig4VPPk
0P6iS1L+cEed8r05irIPnuIDXCz5V8Oudo8hynVGfvu/27lGU1NuQYYQroSaW1mz
HHMOK1wnL9nOm+emvtQfbASXBxnIKDzx1nvS7RcpLPxHd5K4I/k341GGQ0yB1hkV
K6ODX8rGLq0FOWpBBuMBj7WspU3ao2snisXAMcOyxaAf0Ss9MlVH6pcBFJKJXsNZ
+XDptXPbDDPCa+bvNUIKHZN7YOdg4pTNI96uyxEuSV7TEbtEYeqKomTMywCdPLtq
TVUubrfFYj9/pYuKv3fO4utbRLcptDD6fAKyHR2hVK3ENtFa761i4Bd+syBoy19k
H9oUZVdGfpusXq6U7/YkOj2Ini3CI8ClCoHrc0C6zg4f9WDNrVVdOFih83snqphv
RYmMImokmdOOWkhm2UbIOlPLZrNb2MN8hC+DWMjAD5UzydLTvfe40JBTi21uma+O
lvYfnhfuZVb/FRWFez7AwDYa1pMVUBOM+YSaKUihWDL279A12ZpzaHbTnciMx8wc
kfgXUJhte0whrf7sqjNXBvLvh0O3VBr1X2Ovh5bAT/gLrPduJsXCNBH2ILxHhoAo
euVvMiVgYNZQjvn7DKbkqeUF+iYKjDHjyKIJcY94VRyMTPTn48Alre0iJQtiJ2QG
yWpw95BFtWzV7mRFkdtIMZuBrBOUz2ccGJqMWviFDfgctA/YYfexM/KJm5xFt3ia
pK+/NAQc1aOQxYDy3RTkiXS6uTpCcVJVbetvhCbLdidJftMhp2LDS2AHiZZAK8h9
Iu/p8NKsxpoG3wd/3btz/ayD+RLAVTNCQmz5ViRWAZ9xz5PR4v3XLfmn4ZD9Slhv
gGFxu2VubeclUK1N1ir/HBryJ3tj3gXLqvTErQajYPk/B+RaG5J/Xoti+2CPRsBd
PFfbHhCq8CwaNmh3GR4yFgHEyYQ+Ajki4RZt7dfMuyHb+D5wcAeRjdCLgLIMYywt
pvhkc6RuG4wNm+V48j1ZUZfFIsDbq/+g79Lb5bCbajFryau41KIJfEnseAXzsOEF
8SHXAHQqR10QX0Jq2oOO1bADQp+wqhV53i5g98qpMRMlqEv8w2eMzgkrmc9NGuXz
g2jsG+lGpKIe7yfKWyO2L751DhH8OY1JMBtn8ByViAkfk5gF6fqHR+GDRJXBP2Hb
kmHtczp3+YYCbEvOesjMz4A2Qm/r2FzXNYXMwT7ps75+U3xCqRGZ3pvEJBkMBq7f
/V1yDniXohm40ZKwlpFBUr9+Xyuy8mlhER4mHDeZa5gvdykc8NwuA1saWV/COroJ
0Ow2PYBghgtyEHWk9kwBB4242YdQvJwStAATbHy8LJaNJhRtzJtTHaDC3x2sI64M
Pet0fvHrfQbsRthHshxm945bQTI0Gf4U1gYDJCPd0eSLLNX9XllkNZnAdOtyRFuU
0P37sjoy4TJfx9d2jxDA1vpx4N+AlK6ZzK5EcI6j8dPdUIvPTOPdP0Pj4gj/JUaA
wX6VRBs2nQ67RucssV5fOzqHJ0/MKfYy3lDyuGMJ55fbUPzBaUvauR6702eraVnK
cM83JWdmpSv8c0zyizEoNAIP6p2TAyx5K47qlT+Whyh0QPcK3jH2vNYPTztsRlAG
6HHEkGTp9Uw5hRDK6jJLlWsqhOUnMfj3lo/KuaPJ+BavcvR2fvTfC7vOmVmQVPKN
mpSwSKokKdxULokzWtgp2ibEG+cicElB2hI5NF0ShQIXbaEEnxMWA47pLzX0rh3O
+U2XlPT4Y4LM4YU4zAAh7trVsqLa6n5GZLFF6vRzogaiD7rA0kCN/AapenaXslJC
fX6tEJXunssOShJn0bRbY8OPRj84oSiwgO2KCwk/z/4MbpTptzwIfoXd/XZ9Dt1T
5v9FdY60A8Eq+u+XnIHFraB1+3pdfF68pgscP/nFrQOf42WI/rT3Df5fzawa8I3U
6lrLqBd2tThdYi63vB8qNY6GB0XMO5Bfns5i08+x+2EwIH6c2Y7/yzU+w/jCCWwb
g1N3wCM10tPZA8vubuOQM3FQgxg+swluEavHhEJ3MMahLp6k9bhuK06P6Imnal6d
Ng/r0GZYNAmi4SjpemXZAluKTEpERrhG9Dx7bdCDkFBYPohTdRQZLSc9q4VN63sE
Iao6ypWz7gJ8Ahq7YljfPEj3kKFsaQlX3LTMVjpQ4w/NOsRxSXPOlGn01li2uEr6
cnwvv25yn3q9K4ZkSWhzEU9w0eC0rpc75waWmbiMbyW9aL32GErn5UwFLxFQuSTb
bby/LOzNL52QJ8vrYikaPwRs4QHwXMjglmn9IwwI1Psza6dhOb5/FVK9ujVLgcvs
4fAiOncZ52s3IKHJyAWhS9qu4ZcCzp9tthdeE4YDzEs/ik+70mMFkHOt39aMjnBT
9dY1tIrLO/hgCYemVNMvjs36xbwVQF8O2ciWmxhZ/J1Yt86N8KnAqx8OzY6+noZY
5GW/0kSaTYSYRJlp0rrakq/DV0RCcksAfKyeHzV309SO1lImHA+2vUm3o/WMxXEW
Ef7f5zZ6dzRWYfrdWtkUhDS/PqitALNeCPBdv75QR0LXByNLUKvDSHaMmrC3qy7p
Pd+nDggFtIFs3b2FgXvFA/CKMNO18NXFheZVCKnalx9T6MAkHPHI7x490kaNqPu6
gbRXKfBO3A024aYN+3YsPtFCywnFZuWQbJul1ZbialowuSy+6nXflUUld22qlsjB
9uOvNMEaSt4WoKsnziRgJRsPV1Oq36o7kmxdyhHGTlw4diZLoF0rIDL80e5jJKng
GtoPxDH85iAyLaynhjByxOorxujlLwBE7aW/b8MOmGrYjJowlPK/Wi7BqqHfAvv5
T/31MiolkVX9IjqLZ9MjGBHJhU7jopxooZ+o4V/VZqttCgPlIo1XvrX6jvG4Mc2b
W/VLQF/FmdfwHXzjnQ1G4DILWHPVsNVHt7YeOgIUcpAFJb/i8j4CkPSObM6GPoto
Yh4EomRKD++MNaVB7P6RH4u+EJWgKUoCLRI73V8Xhz0OVRjFcI+/PrlFzKGMjwsl
N8Q6630tYO4G0+YmIx8urm1WdfRFsisKLXiOvV4CAH+LivfUpaBYu9w7bXeYhvGT
pn1rwjLp+DmrcqnTkUC4kIDZ/o5pX1/1egpFaNI11ijv/zoXfRd/ZaWh/c8m8do7
MhvZfPK+nbshQZH/kBp63yTj/54BwPUOmmB5W7Vc6Vq0DrxdLK4TFi+6dLcl+fCE
SOAN/b6wAaAZHxNyw4fwJ2Vy85rNseuJhvQlLBC/rf4oDce/1c+YkUj2qo/T7224
t0lm61KB2yq9LEg1ZVnlOGNw8fjgKfDeGl73XeIBUOERhz4pdh6e/ORKU8SMmqjo
c+q45t+DkNnyK9dANJoCJkrI1ijfxjhkDWtIrSYbdci/ctypEqjsXRDTmkJ9R5dh
pv4q/7o9bSJrzoDbvl8nNgUiaHhF15l1jgmxm6ZsF/uwzDFLsZnHz4bm0v9Wc/As
GQdyFzzEmZooUubR4CiwZUV56Ax2TmNcj0Ov9BmrErvclS3m/u3a/MR6yM3+sy9f
OKXkKs9FqiMtAHNQYVUrMYU9a801YNQ1uEs8cdxkI8m2luxUAzn6ujW33amxvFob
0K8hHkt0a9UmK0NOZstvojSzeRmm7A/i5ZqTOjXIia90GMt22jqiy6z6hBz4DHPH
ijm0hypMiz7VUIgWrdf7IFXSkBUmnMZ4KPJ6Yf04XrhL3+KbdMESf3yVij4aF29u
b24JFx92Q/zqP1Q5t9MuPtrm+iNKieEppl+O2C6aDGcy7aDjE0gP9XnGslXoWQX+
Z/4HYYsAgjthqyVFWVw1nT28nf95+ZG2oWP6LGo/BuZvONrT+0UuXnij1vxNiJQ5
uBTXTxKuTPBWFZexpzQS33Yky+5bI4EfQ4ktPf2lcRSc5DR7l4hk+SdFqYAg7o6q
jvulsfz+OJ9TcXdLIi42KNg4ZJA1hBXx5cYBL2QfrQCQyyx9WFzeg/TWi8TY0/CC
qu90q3IOYBZWG5SAgDpppCge9Gv2F5Fzp5rANZ/pub/VTh7xlY86kfyrfPto91G4
FbrNRP/o8eKCd0+rUhFdjvOeHJg6jxCS1HE/9hGp/osUhGLEv5zHRFCTaVkStja8
qNMJeRzo7na64Uq/WJtx2E5c8PbjA1DZalGf5+pbvKGILxEQtj9wGHR1UEt1Z3gK
3NYH7pk+neRGeJPNT05Uy8qn64y9+5KqZl1kCNrlfoMq9VFMd/fIEQ3H0I/xliC7
4FplhfG9IDlkx+Xvq0mgMJHZtIxnQ2fJgtBB6+ffFdkH3mM27Ilngzap3by0Euah
WJqgcl0K5orF+jdRAQumkrJQ1/2wXuV9x+48bSVJlvDhFE7kkLtDwTUNdwmwVr9m
ZFpF5vbT7ERjV1L1TeIsowaHhGuU3je0017ie8QegWYfRiUHVtclIVQbiRA1n4m3
Rrx98PiChYyoF/BXgxhF8pDt3HlfQurldHJx+bGG1L79HQBuoTYH4npaxrjdKhGk
9DLB0Q120Nk96DtOii8E716WPgEFvw+bkgKiT54KB9HEv9CqHEfqAqQtUfVTBKHb
OULEufx8HETi3A+5ouRH8u705MsMeeNxTLMeurW6IoLWpepa/iqPQiGL5CpmYv1N
RdDtH0EG09feGT0Re/jC0YK9oedIKX2/nFF6fIqfsDJ/qzNStjMah+T1iksJfP+N
9ANmG75rMmN6girW7FjXYP+AtGYrnsqmoS959oS9L6C89QwxOOHzSs+VtH+wHHlY
MOyAA50KiyEkR461aFhJ6t/fqhD5xWM+XNScRlF0kQdqGcGv6xxPTw9mI1adV/Tq
VAmqgIFkV9NG5AheUoqQNbf/zdG1O++7nvzmBHDZbqyEf7sqNFEK0g38M84+ljCU
YH1WrlQMaNIvJ1m9MecJ0McGdBS6qfcJTQWJ0MEWFn7wt40wZ+SUSM3q+uswQs8T
zPnujHgQ8l92eWlwyHE3FSZ76xxn+GcV6PJl9KIn4HNyVrqUmT41AULadrZnbX1D
RSaYu7kz95PwpuHvilgLEaKW4BS23d0tdyxSNh39NCQGkMTN3xUEekUqPQIzhEp1
zIpAVWSffeNo3+Ahh8gJ2pf/iNvQhhu0LVUqzS4T0GNFMaVJfCOyThcS8+IDGco9
MTeXZifrOvuEeYAgdrGqd3jCOivQ+nx2MQrY6BGzC9S+805Spun4Tucp4QZwOX8e
6eJi0hxOxpWwO34OAYhG2obKdQjtKgejspGCkvjNkiTEZFfVmS8kgXn/Yj8x/nhu
YA0lbYQctvXVXCyvu799LLTxxph9OJ1A3KnopRqwqKQfDbu/VcPjvAoWjrXn5z3F
tyICLnWfehm1SrmajWwXUXdHqXCZg5CXF1h3JARcFgV0L80S8XlfQwdP8Lc4yUOU
cl1IV5v48GRP5ihoTnKwO4Q6qMy+fTE38YGt9k4NW+IHSP0TGxVA/uMLfxMfV5Mu
W7F2jinfmzWUHCIQ/1/Y0EBIWDYsDbm5geML6U1hH0mhgUbdE73lPG0WDelV9UWR
v0c1JCts9aNwZeWpJDFbVb1N6sY8Webe83SrZXOeIP3c+KkXxvj0+jZ/qs7OMaV3
rJf41M5zNHoADqttLzLwhIUUX9l8S1tVB1AiSHc1nADeqRH+5LfraY6pqLz3dUZE
WlGhK/Bb8hfzbK2nip+d7arAR9XjLg6GXI40gKE4bV8U0ot6GUw/Yuwyi5KKtVln
x/indqlymkZkWI89KguDIU9xHRfgwpUjRNCzqqP7QQFBUqaAv1r6xZ9l9LDLLfHP
y+r53duMJPu4/hjNMZJbZ8wC8iPMtxSqm1EYwzo7r0jqqjTn/DK6Y0n0hUheU/A3
S78G66yr0//srZs96fd8CzQhw6tDTc1aKLUG2o8vf50RgoQEhA/dTx0NtyiKdkGe
vfrykXjeSMMkOxMCeyPpy4DxcMb9STsuGW9MS0c9T3GiF0qXmVtd1HpHV30B9Vaq
GyLJujwcXoxSvIwW8ru/ugY7m0ZMbDTTKK941QopJNXBLj7VgEtI69OLCyiQwluo
Dwx3aj8K3nTLcZKLOicoZqfYEEkJsLDT0lmWXgDRm0JQA/R2agY6a+jL38G3vR/O
lGFgfiYX9rDc4+VJvFpZemcglPiUtf3EU8AeDb6Xzm+33EMiu7i8+XVHAPal5ZHL
Ka5nw0udnJyuUFAL/jN3NOkhIlKqJ1OtXhJwptpvlkki6QpfnPu/5OrnZwqyDI3O
sKXjEXVTNEusQnVzci2YmOH2ihRc0hiURHs2c6Wd/O9eprCadkl1YWHdQ2rAha4G
ScvPO7wcAWHAurXnV62mnyowyoc1IWW60ViRE0Hi8wMaLKPNN1U9/FklYGK02xAP
7K0JjaKGJQa7FOJRfO1P0bUzVVE5qMcle4CdSTzfOdXx7AU/jJ8iKaY5KLldgF3V
vLpl6gERrwza8u4oUFnf4FvEmucyXkoK7KZVmElhHDmUD79Y0iDwuDjcXxbFvyr9
FjoyYBPffqhGkbJfnVd0rI0LDLvdSmI0QG0IpYQQk734zh6kZdWdMme6Bbz1KtAt
nqeUgotpz9NC4v0H2F+KaY6rjuSzibx7rccT/To0G7jGOQm6RwkY7Lbj1e2oJ8mM
eFAQS1MNqjCqs9/7O12LYQQRSAVNmWOAXteahFz187tKy+LSmaeIh4jnURvy71I6
px5O/CZwzeuEs6iUZgsUKxVsU3ayxZUi03yKKokWljS/f9aBKrQO8OOJfc3W94E6
ZEYC09ytlzVx3o4y0L/TwX44IzbV0MDNJ3+h2dGPqSD43hOKcJ78AKXU7EKzgwCV
J/5HAeWefLupzPc1mCqTbhl3acntmwnGfZFMIQDuPgRKMzyE3iw/05fiDipzgmjC
Iv4CyuOsf9Pbl8efvC42EU/pyJeoME28ArUGyhNLzLtrKuRXJwe0FAGMQRQTsqsj
/vTUtkASlT+QAiJzLCKJM6Ho7kQPxh/oZklIssFS21oehW1azivLbJv0ATidI1Du
z3QDp52URdv/hkzKfXPkIJjtplf2qW9j7UQ1e89y0ODSBiNA0czACbWavhmRyQiA
kdCW+Uu1+jkLkp55l2/4yleY0/hsr6uNOXdaROyYTLUxMqJR3kMGch0cFJxNMmQ0
yll/snq8JKfD+aod3GJxZMJkRb1LjiiGFqzuC5uDBXxb9UDQSx21LU/6jV9xK/L3
GucPDIXLZ+kh7C7jlnhRfn2s6sbLkmzpmNi/w2w2+6jjZpr0u8MMHrTFR1gh9u6Q
3zitGYCiU3Oe8rWsELEwyo4rReqle6bNkOSmidSQDQ/PpwJLm/ucIzPE+oVSZnk0
vw6EMbN2ek4CC6IYKAnQWcJLKk09I/tPvA8oCo8nrt/mlpPAJOyFyDvxi75wdxgb
8dbppF6yzQTHT/mjpO28dhOifB8CBCR/4zeuKRX30rwjRMUgTXNJx42oml3zFAyZ
+Hfv/wF+6o0RPR/ePhgo3MG7HaTLXNpWcox+PKJixtIuBB7FvdbF8CV7E1NIOOKo
BwecVCGWRgIIIMF3vewJ7XBX9l3AgI2+xCe+Atdu9WEW+IocPTHSz9YwkeMJf73d
FZwNvnuXzbdQCGbOIzh0x/rKDnIzZGlKhG/J9G6TStYTUJ651oupU6Dl9FN95N+T
O17eqEsY4X2XgMSY6/3Gt7MiuxG03ydxTg5ttZ/GEj1ugdKfjIlpU79Za6HbAQwF
5IGemkoUP9bhE5Klln2HXYd34lfCkr+MUki6ATD+1n6KQDnpd9AvOfE4W2e8nRMx
/QAJ7rdrbD/oOMgu3VCk/5Pvs3EN8W+NmJ0/ScrDXBkkzgZx3uBblPPHxE6qq2Wq
UhtM9a85864YVyR3oid0xwWCA959NnlqbX71T0Dqm4pO1+2iipoHaj4h7rsiFdGe
SVe3s2lJSTKXbzWlDAFTuu4+0D/azvCKiORsBq3O1dOcaxAMuK3z0nFH4Wx3/U1m
/lC89UK9eadnJDXEnsaOkAD9USJbw/eiFU925yebmWKTkBVAts84bfWNgjWnzYu4
p2dPQWmdlOs5nMQUMwn4STt2zYIWNZ8H2ni0K/lMdff1SzSPrvSwQqsErT4l5v9f
fF4oVRMXFvzbmWqLmpu5jK+Fe6qPhm3q9U/Ov/W9IroFscn+NG7W8sDJXt3az/NI
y9So+wSakt70gwtKgp2yyCYD//kzhlfHLC1SFFRuiwz+aS6TXYA1fBGLtA6QiBlc
206HObSdIwVhdgh33LRtrt3Ln++fEV/3BEcYICwTlee06yCxf88QOpmKc/GFBCxP
7DFHrg0iZ9totTcKyTQcshTnVcUFI0f1UmHpHeN7FqtiKd7Pkrs5Rj23eqM+600S
K9IV5ydsxp8W4DJr7RFx3kjV7gYHQI/xBaA+oI6R0qA+2q3XAdlKi/maFyg3ih84
I4fWXtvKM+7hJ/XQTinNT+l+bVLECtwnvicl8Cc7Js+m7W18ThaLHEGeb+aI/tBF
BaZtyqNOFtGEZn2o6/K+ARf9dBC/PbU8yhFjhLa4ZjTWT6Un+lbDsE1O8Y/3iJDL
icZ28zT3uzNaatdv+h3rI1JB1ac1srP0XPrSdY5TpTW8RVIVtTqmCC26lZEl9yPS
iP6QWsV3T3sQ8/ksyOOtdGWQzLhAzmBISoEQ54mXEhZkh1NL+emhsM5fg2zBqQle
BBB/HB71T9jNFKvcoomVZSjBxAWpMYzInW7AOyMepQ5UDp/lY5NA80Omt5KC+mRj
2l4r8p1oHHRDVhbNniT1T/LBIjwEswtLeYPWzU7xMx1pjwc+X1CP5achYOQuB+aU
uTmhXVjViY+Qc/5qsT56V69m/gF77Wi6AOoIXuPiKYHZ7BN4cwDevkQNMYS8D6Ei
8pmogZekvja5HEfRVrc6+ECBPV4hSEWjLUJZjUbARC7fCk5lh0rdzu0+yoy7Z/fV
vqi9ZUpLu0xLYgM7U6FGASHEzg00murL3qRip0SYK7HJpR+RxgcW85hUBeLZyGH8
g+Zmq6ajLnsdL9FIPrz7P+NJ9rimOtl/M5TLwaGKHd++s+d+Upp/JunnodxfAzi2
0/ou5u26OxS6j1W1a07Ku1SvjAFmj0ACuklDgzY1YXO7PSWPiXLiij7+FqSpaQ0Q
/BW0QmgIHCkmQ4ZCMlAgrjxUwfbRFPjWcabvXZ8sIhJafNsTXoOGlH/lC03OUIaQ
VgOFCP2VS5VpSnSG9S2hPRmKwk85A7sm6KhhVIc35mVO5Jl6s1wUuYR1y491PzPD
UzqtZNKa/eLPenRltwqgn6aGrwA4FWWBL3ZiI1If0Uh9zsydAk0Qv+CrwZp8e5tH
CR/iEpk+cTku8alZLp1+K/Hyqa6lU+/5NH1lS3zZ+7UHFTtl+ygGdZj64xzh6uTI
eHFZjjPt37rqsrJgtTZqXuDHpc3TMS3dgw+mrHmjvljTuf4LKW6YvtXZFAjODrE+
UBE2GosY3Iputs4JS+wYi9L0VCjIGcHgjx9KqCv+JWgceMM0xqnSFLVttg+M5bc1
j5pUgEEZZAXgtkAgyBHdbY8cW5HILhthidA0gEHfx/KHl7hMRShFxAdPnbHNlOh1
B4nI8UaZdcgE+WwHaKnKx1X2kd7G/+Z8pXeWKff0JfjyxjA3TFvpFnR/FyogIx0t
JmjDZGutVMvDNyq3yPblF9OT3rv55eGuXPVuaE4+lHEFy1Zp9Snhv0y0djIY67ME
djjdIq9zzuGRDm4g7SnxHiB8ytYiwcDFsj3J30dkiKOT8VdwBNI9iUNBj/UbR6VS
kzA15hfgFCSqahT3ZeDG/R/VClMgZ90psZd6WAROiNybznjB5f7OQNhNj/qIBCei
Nu/Uf6faeo28UojCKIdR0kd+b85cbRV3vdc31O0UmUyipXYwvAUdi4Bk5F/eojuY
/F6ebYGI6CTXvYlZfSrXtHKU5y99S+V4DBN3HhXmq3Wh/CHRuVvhcWQr0LaY9TMh
TRN3/m4iNMIQ0Nc8bLXRMDKEoiNzr8NEPIO9juxS8IUdcDNwmpm0tqTUHsQMpXrA
trD5gkAgBbPNQbAEuFdbwzqWxeo7LRrcbiV8A0pgYyLWWPcZgEpotbK7X1fZNbk6
HvDUw4FccyOOcvcJsXQM/bDEkWPwqVkEeU0fbn5qed5ARTZlGaLL3heiETpAoEMe
abVsaXYOosBPsuD3wiqTknMRRfO9HMfI9rYZgXlSFzPAaBypzI0fIJ5YoR5KI+FQ
ACo7lgqOOuSAhVi1sQGZ4n8QAO8XJdDGzQ8gwMh03xitMy+KfATnORiBbHJTa0qf
ZdRKrN/QW0jEnRGP2mJpuxCp80h3q3zKb993seczY84rmmMAFpOHTr1TE8k7AcOF
plcJfuCoGQlMH+s3VXhvSi5SQamLtu/s5ozwKTIvsQKsGXeDG7dxf3H0h+EUAnut
r8g0BkvtUXtUrAscP+nYmDHTlsAoEGxmBxR18NOvs1lzevyw3Advs5Xt23ACVWOx
+Xp/5eWJGBpuoD891A7NZlarP+MgX4AGl4bDERd/uHOhwC00wfinRVbFPNhSO2yo
LLVr+K4ZfCm9+8E4dKS11Fb56sDYRNtBHWZLVI8+XOOFUCobCHORfuEaaHUl+qbx
5oyzB7uaIq8f8o+sLpiGlFJQV4GFSnK7gouV8miJcaW8jyyE7P8kKrruovwqqWmr
06Dq6Skap7DWRZhjFlRgRpRNSs1nHwL6Lc1KwZt8XunME+vOHh+R90+TQxEsHaI2
NG1F4nBYOtTInVTNKuRdx9NirgcA2RRW/l/8M77M9jP130p3cYBECy7OMLcwyZml
0N6FBpcems8l23eMnrKUpbIVO75WrvrSILuV7ql0TzJm+8QJfMJ2yMr6eEoIVxSk
De3xf5DtsfGKKSUG8tCHZi+FCIpBG9o9/su7ZcqImdrORxol62mc8C9Y8yFYE62X
Zc/JPYHGnz8USUXpmMetG5hcrY8vYOn6rIMuz+w7jSkYsfj0dAtUUmVvBCV7WkiN
qy6T24/5qWr9gYG/vn3EvaOcWTUgXXgZj07X/+Z2LHgbjhb3iGRuSSpNn6vc4ee7
pOKtJVOyAZIs5vxuORy5V9yFl+AGUNBcKekS9gepjff6Jygg3EjSjtuwkj5ivluq
AsD9dsdBrEikinw7M4ShcJfDLS4RwWsDV32VPdgapnWWkttEgmXRLvsclDqYj29V
yKPCPrs/81ArF4qQ53iJL91L2YyFgOQe3I3yNF00i2oc3+nBy4Ipfe4sahDjZqpH
xiaZFTArB4MJap4L/hU3a/yTZf8C5s3Oh8uah1q1+IojQckRtkMDPL5cr65348Az
LQTqrfmmNrHhQtRoCF3STj99neDoZROK6RS/OjPDcU7qskybcQxnIzMwWnp+jgnI
GYQhme1hR9sUGzoM6mlNXYY/07zqEV63uczJlbwkqhFNLuqWC7nRsFmh8rMtDEA5
Rvn2Zg1cW1a05jU0Lug253n5Rn+SzDMnxX0Oy0oHf1P77mM8ULoIdnjXTYLpFXrE
ne2lVY6Gv4CrjXpWtXx6wQTKc5efHJVfsvty7ydYgV1LatQTmtSL2vwjqQpTZ+4S
+WLqTYEpzyHy43/jA6f8tP5QiIqjxpIonrv0ZAvYmWopDO7rhsyW8NB4bd5DyX6S
tQeGduWY2bgMpdzErwsPyWX4hTGYShwhZRDQNZtrydE++iES4vCl6mpC9BU9bZCW
MDkD6yZFe506sz7WoQfYLp0VgvsVSYlRAOGA4BoNv949iHPIy2toHFBRLI3KFEYx
yo01/wLtxGL1N3NcgL/0Ge3ldM+5JkV/MZ8/ZA46xbdmBVa7gKg7UGo2Jz7EcufL
5JkQqCG14347aUBqiUIXsVUaPomFmbpv2ZzUMDgxTrd1jlE2YFEWQtNBj0ZCrJIp
Hzh+QOZ0pLRHAcTwICjMODr/skM8TgKpSxlxC9e/jDQohkjTqTIHK+rNLosavPWW
zvj+vp2mXzJJW6OpZvgMvqMoCZP7nOS+eNCwWq/QHgs8FMbu+SrLn5xGkzf0xXC3
bfzLBpWwfG2wUu8jR4N+Haj9EqdAQ8/Z0L+sJIe+S6AoQE+5Y3Me0+xh+0M2lT3G
ZZvoojyUICnjJPOHq34toZBvyMXz8y9T/l3x9HwBJZF8NXqyOch3QkRgjAd71djc
vbHTVpYKj8Ou7RYP5Itpsw3A4fd+2CKj5LFk7EFJOdpGxY1VfDMBXlbfHzlQrATT
MZ7e35y+ublKvTo85ahNLNijZ28Uz/qEXbEjZ4C4F+HLlhi+OSmCiBGTLVvL7IH+
blnkGOdeLQrW+xAyGT7X8HDMAcaQBVm2gTNzNdoC1QhZ5r24QGqmiV0Z+qQcEzbJ
uF4i7oFxNsFUJwr17Z1KjJVoVNvWgQLzMifYESyFFu/htR2c3CMvllntptvYx7mL
UKc3a5hJfReJan65/yOvT3iPVQsDxpZIyLfXmy7pul5m3WejaY8yKhjDkLDpKmUw
NMxCd/M7+HK8Rv5+Q1t+GwsYUEZprhKSPWjmLOLqGkyABVEnv98Yl6G1aSxG+rTg
se2DRmRXjUxrhtUbWJ5uMpEPkkPYoLtrGajM1gMvKy+Jj/u7buOxWNV90q/zLyN+
xLrmzvdqNY9KyQhnavZ8XVue9McHbKEWJXGrjhn+PGe08u9/hAcAjS3/cRir1OVN
Zzr+bxErX/TFfAlJprVkdETfhbc3USAT10zKWK6I5/XL8mV2cmDKA2L0WLMAGDjb
n/N75F//nvS17ZmPBHIKN+fOnqh4ZirHQ555LWW1PXMtjgHP0XMGmhOtXYV11N8a
uUnTyS2ZBdmRmJzbx6ytZ2J3wDv1FMZGYGQvcXznMMbknF1V2mnH304VzPuFJaYJ
5wrQxAEtXABdeknVM2ZGAfwN5rrwxwNC1encXyAfSTed20t/+zaGJawOU1SLX8y3
6YXI8CeFF1LpvE80bkjP9AIKytxJSAozuima5DLRKPE9zMXDWHmXiLAvAMnP9ATh
YW0yM6/0OZIel8liDPs8pTRnGtc1r9AtaAho+I8bzmXNMMP6UuiPd72en/nuV0BM
u7zXNFQ5uJ5hrhTUCK/HNhWCB8dc4ZqNVCHcTBOSxMzK4uynuvd2XHDkkUKy3HQS
z0jTBLalLyAwZ5RQFWgtreZ5dgKWzdnBBzv8EbgEv1e2obExFTYVNjpt1rlMFAKl
BFELVXF48RsubrAXthum3BJHKjP+1HUWS3fpsmJWvcATSrsZUGtT13nNsgDC8RlB
cSt48t3/cRU8rroCH/P0Jiftv7chZpNXZhksfP+f8C/zZBTyJxH5uyp51TVuMp52
97dhgJLY9pAtXXDhhJFpc+UtPp2a15/0DfHlzNG1usMSH1+eAp5EURqFD/Y0L8U8
rNlPiib54SU8DtPTGMZaDhkY6lp7MQZjmds07xs5OwcZPxjlSPX2yVkeL4WE1DtN
XeBj0lQ9JUolCMXL/lnjiKXxPbHMTwwwKLwEF9X1QKtUPLtiE2dhP0IKHlgdMoL3
A9rwAvXRoxaZ4rFDEE2ty5eDHRllPs3dCWGBeKGWyTD8xD6x2E7AOR2Wxi/iKcTz
w8VJgHON3slwVYtLw0UIs5IesGE4uYgvEY+6Hteh5BaUA7+hl5AkEtB2oRVbJyTz
d+eThX3hJT8qr7+oMsjIX2bFnUidqWN3rxuu7RZEdJxLDE065BzdDk22jE6KDJ2X
ohaOjITIFwF3cU9yUSiKl3VqM2LYwQ46o9JFlOTl5/vigloC6M1oAxu0/MCTYtQD
60Ml3QnJz/B4KTv1xF6oLkcFZtF6IaumHqvzO/zNwsvG2Wus2Ah3hnGyhKVeG+rP
yk/YyphJcn90ZITxsspFleVmngIWvE2+OZzJuXi6bcgfKW8VFmkOOr0aRPrdhXEh
7ja89HKq8kmmfDa5aJPK5zgWUnSF7+5KcbCIwPmVp4YV8uCaO1GogcHKN8oTtxKY
48MiuXw/1xWITaTNW4Qv3GJtwVa8l6HJY0S0bKIVhbxVU9RLzJFBAAqb9UtsySPk
MKC+HljQRlshoidF5x7rztQKiw+gpMnNqIg8bpr2kWi6jbtbo59AgKkZFRbgUIh7
d9dIoYfjyAU7EYZz5+D98dnn3DpFg+BwrZ+0xDYQwDQY7spambpkO9GvsDSdSfdf
8MX98Lj12SGSGkPQUOsTQPENZVftPtYrBapbqiaoTlGp8zbcPR5L0dwx96yfmrb3
iUUs5tRZ83ki/txRjVy4sBljv5vLt6UsS88a3ufFGWkZgSNHNev/cwlc7ZjH10hk
idMx6v2Tn20wDNHlDxhYbr7s2153792NiKG+SePnIb23f4RGoVM48n8N2QBq+Fwc
5+iVl6/Cu+qZ9LVmVdAEIxRtcUakscF3+hBZ3WnpPSweA8Swdl9MT9EezS6qOOjE
LLC1fd5YCNCXnOHw3QiZB9XwAuFT3wqyGeu39Wzbbqil/HJYK7FDIt3hT2GUE+iX
lnDxu8cYy3km6GMEjHUNFrdM7D1rugsEQWUm+1iQXueiMJGMEafZt5tRCcYVFFoh
zS0njk05oWeiP81qWprjvfS2UdxFv1ca1DWU+6SqniitFdKWEHu1YoEEfa0e+2zj
jZQNTS2e8tvWAVHvTCUD5/2y4WdKuVSLw+boF5RruoSKHu562FIXJF5/bNbmBc0v
qZA0On9qSckUN1eyE1XYHFBYyjFVr19qL3NcFNoKNyT1ZCkNpJt4RQCDTEcDB26/
77j4k31a2pJQU6OkhCKzG4LZqaq28HzEU5w3TnNQtEx1ptr2HjkXQ0dQ8+ggCKix
kNA27Uj5wVG6QRkhSa1TR88rDXoB+ZNgpDxkc18dIoUgzHyevtwEcc1E8+RY3lqk
DxegNVGsUpPdtQJzZuM8s85g3W6eseNf82T+89RELSEt5VNLXb6QMK0d59azb0sS
8KZwiLCAaomLHigyafs9Wwq+DBgAHrWqEDz8D/ADrsA61W08tItUoF5ISty9LeQV
6Nt7pHdcAxxBf1hae6tcWaEjJJHlLTWreZQYGAbXOudTSvGp/FgqF3ESnTRT8uyJ
xNgpScH7WrKXBB6g5peuHwJYR5s/ki4LPv/Hgj4ty1wk2TEqb+2oDTulped17lL/
qPTPLh7qIgXuI156Lb+PUuqmsV16UGAGiBWAyXIzA+wPWRzQUp7nlBFMJ5Nmfs11
Z6mt3QNpa8MkVVdagzkk473obVjn3k+P+CjnqPYhYu70f616jym621w3dELNExiw
ju9H7X5v2tjgC/YaK2bGj2Bs64KuKyfWZksz7s0vJdD///g53VWM9W66QHCQP44+
eB/MBldXWE0yqq4q/l00fhDQx4Bur7yCQU3lWzBV5N/Ampj/3xDZ1SWMNDZoGU2Q
jThmzbrsOLdsBOyVFGspOV2ou25e+O3EpbXuPqQBkInf+JT6RKWTTGjoyklSsoEn
7Oxu9qCCggUnoOECRjrl4dwvDtq28mO4s6wcQGPmxmG0ybiPxh9IgPbsrpJE4daT
ALrbaAd8esQtXQSC49jmIjo+vRLMfsuOMY97Cd42QWwk005bYr3EA9tOl0VoRpzp
EZmORoPH8gp1nw6Km+gZHPOCt61DgV3XH5iXb2WdgWCDwYIM3TVcTHz3C8NRTIA2
e60rYq5t0vQk1/6SbXK/QimtFVWSLNWhkkl7/9adMAztn1L2C146i9DndZq/3ikL
rx1bE0xsMvZDD+uD3LEhtala+3Pw9++TEm9v4P3M19mZAKv0LoacBLWzkrcTKnYx
MZ/J6noU9LpblnvgXaArFCcx06QemkchC84gv+LQ5uY1YC/jUcL5gZ5rAlPkESTe
IckW41YusmqtE/c4mzmI+jwzquhVks6SY0DWf3DB5p0s4EQlgTC4saC1PqpS2voo
nKepu3N4rdJLDbNBYQdoDPGqtZohZygFa8MlEyJyqCw36WssEvDg9qXkrdjq8tDV
uAyP/TsSfK6PzzJOdTHAyjLf1MXP4bWQMGZXO5vFaFpjroSf6iAm6rjA2m5jV5bE
svXF8oChyyjuon+F3nM+faB2blk0YY169r6R77O0S8KWQ6PH3vIL7EPqkkmiWMhX
88Fp3SUTKd9lNil8+AvJKi+FxlTyDyzEgohNTbrrz05DDg/A40W5qoZWOgvlZ8sY
vH/I5Iq+qcwu1sTGAuaj/chUA0lPIUZoXiC8CEfYT+8+2+6r2lZcMCb1R34FpOIR
rNApKc5hPpTSagW/+LIvvkYGD7xjB5AjJHcS6MTdGbFtS2M50MiL9pfDmhlsQni4
qpepwbqESPK2M3MRrwaOJmvcUmujStgTAeE42oYAhVnJa3yGVp6lw1qNS+pRJwuV
1ltjHRJA7Y0BnKjYFWrNhcRo0svdLffRL61fHfLxeAV0kjwHl2Kwyf1rQbEtQZFP
fVYxnB8/9zmB5+yP10HOvzrPECc2vuqmaRMHmo8ZDapVz94xPY5qgKPHZCrgu/7H
BXjgSaZklLDZ9mQUfNlb1uiNOUJoHaHrw9PKY4crMjHNUMqs1gqBYsZOWLbKlHlK
GUvrDaI3Qou8sqEyDBYXx+Xaax8UnwAeFIf50GXd8QstBYr7yr7QYjZd/id49obg
LcBmfU7+wALswpM1tI3yHFJhyz+cKk//jk17eLrAs60lvBIMqSTJoYvH6GAuSajQ
SgJbLLf4vZRgpioHp+0dGtE+hXW8yeDCzyf+kC9LkdB/kXzrPcNUxi/xPi453LTR
HbdGMouYWtghn6KlYdrYXi4EdbGQf0qIqiKjPwHbMs1tIvljl61OqpSm4vGdtU5i
T/DvaqCSQmeFSj0YGq/1p1ZCuQXPa+/S/MLXmhdVeFztl8VM1c6udxJ+mg2OX0a7
P4k3ELa3yxpR3Y/Wo2lSgINAlHlk1MV4kbuNIaD8J+vo69S29eMj3eI0l4NMEOhV
72VS2VxzuF3XE/j0y8qoizWLut1BmnyWflYdAKLGmurxqfxsdby6K9+1Xg3Ki3sd
cv57Ntfz0OcSVQA1NqMAh0axJz9EHQznTOVWdXeC7TzFBmov5/6NAz0hkTBUrWX/
4YVrO6y1gAMAvX8lqb4YYPjHNeO4P/lo/eysMSVNyd7QcZjU3U+s9xTXcS+k7p7l
b8pZVfnNqwYZdIFxcqnl8350kNuq1quk0pXCgqEX4KPzABUhaA8M91rJEKWB2Wkn
LyEtBa5jdAUN3Lzir/IhsB8uIliB/Uts3zdjSTU1MFt6TW4excWE/0P/TfRSYFaf
9/Un/oTJy7Eib1N1dlYdRrrqIl2WfqlPj20ZQZddFkU1OP0Wcdj9w9F38A64UQHS
/oASt/Um+k2dz7OQulhrS2I+cwBiESnw8sYEScJlOcLsj7Fvqt370i3C91f9F/8f
X/6XZg12CdRtpTnMnwEizyzq61p4Xs3HMEtbwOCywMYKrXRzI2ah9DWewKGZ1t9e
H20uJG3R31GisoLYtCMGYiWdPg8vwVZFBoIhxcGsva4YFlcX6y6s/VBged7EmJB2
But5Z6sAbfUvlZKe2U5U5WTZZK74An+62jC5uuOabf/oWyLsYmvW+zBKiwe9K+Or
CoC7R1eAPs13kXNeavwvPdP3mqmURleMhRH8OzXG/yC6LZO5MLsF1GvD7tn8KBRq
oJg9jTDUODIbidJ/JZTtaZ8fiZ8oDsFSqtBFYHW7r18uh0m5iT/ggDjZAC5uzRHl
WbS8HBGDxnqcgf9RBBIyr9/v63qfsdOleGKMcXqIDmgnaMuf8u56hptdIegkUtx/
oKHn/JOpnlstREKWTmLkojdng14owPv+7L8oIEpZQsWYdFFqYCWuJpsFPAB1SJV3
KhlQS2R55vdr6QQtc0a7aOgz8xupq7VZRa7G3T3i966qDjCCO5WMMf9lUmuSBcbL
e7kytp0wL2qJKYYxzRhx/jCUWjf09D2KObli/XJ9qrFmOJ8mWoEBX1bfxqLPJC51
D0ss1BZPobwTWx9bH6UjJ+H3Rna27LNLB39VNj3eu65Winc7zx5OssAG0kPfEFRq
rw2F0jJYuOmxoWO3UAuvRhLcGC4T5At5vzoULMn3YOz4lWFSBV9/kibM/R7tslrR
wHIoMTif+LC9m4IwI8LpJNSSP/U/jWy/RFsfW5e/1HGRFfxVwsRK8UvatMSb4xFk
xxmZun+szUYnctJ/58+45vYS8bJGitZP7oHyvAt1k1qiZK9UQp/Pdf7QstiLi39/
4HW2cgu/YHbQECFfFI/nJvXDjqduT8ZdqzVCdCzGG8L3fqByraBBoBvHe0OLwbmr
womtEFE0gMPZuzJcq/hG+BYyL9baSfzZWAwXyycZ+fYQDYXFJISPsr4TueNTbq2v
ZNULgolw6EfXwWlF/zQ7lwGnVS7AmycWaho0LR9yS2wfSUWqr2WnRgouBJ5Q9bU2
46Tq2PIgcVS4v6TvNdACpcF7buuxQLEAmptd3nQCFPyR6KyH0ziDyywXpJ6K1eA4
KXEccrnOr9+aVJX44/f2GEgKO0RgnOH4YE9U6uSrzHQYg9+yt/R0wICarRBXCUi7
8a1PTZ+bQi2MY+fEYXVBbwJX8KAYsZY5kbTd/IPFN6pbZAf47giQ8qDjq6O2OBU6
u+dLkHtVEojbcSFv90oP2pA7EyxlRjzsI9hqCxwrzIFzBAiO5NyX/cKbWFYTUDWG
X9WLdCEJRitFJ4hIZkHzS2+YTiOxjKRUH+HlphcRDnSYHa9X563/lPUObvRHLLK/
LrIThzknYFu/KxFapFllmX4upJbtOk1bJZ5wxLonZJm7vaj1XvnK3ZXm9qSqCSnT
kiBYM9Epr4JXdm8zFenYLkekoKEc2IglJV2eKHCTeQ49cjY6rLOyY2BgYnGXKS0h
ndnn2Vc2fR6q269D/eehGaDPMflZp6IdurMTfVFwNRlVR4ukuUGj+IIDaAGsEmP5
vjJs9I7nJPDy4/7JOlfnBzj8IHY0lPQi6qCyTQ9wgzO6MyKy9f4nxnCg8mv7PmZt
c9VqxpY1JlafcfQgHmMn3tNZ6wiQD++RSlLJEj3BWmq4HijWbVnGPdgN+ywmeYTY
CLvk6FCOsng90sMxk3F7IA7iEyfB77PjyswT0Lagc7FX7suU8hOZ9os+ofAWL04B
sEIgmogWfWZGiwAPOPIeuIh9Xf/cq132KCI7eemqjjpCY5LuvMiY/2yu6uzIzwY4
K1azfS26kOvqZsqoHLasX0J+10AooFmmYF/SnTB0Q8sh8oW5ysfPM2LWJBRLSf7D
HqYuZnkEHoK9nBXYTeFTO3p7uCwSFGYR3NlWbbbai1PocDf2axSVwqr6LD+E29a2
ADS59LikI6y4CsuB44xOSl651KQ/ihD20tJSpZ3i24bD6YEGgPI1ioefpxJwU5aM
nmgvU58w+F3FkDE7Z1VmYKKoXZ5mdQn4xBdfoX7TNWoefjjekfGacCFOVVPs3ooQ
P1+dhvWYD/LFB06HFrbuOxWy67m7EyFbb5bOBXaVonL8wfQCWXBK2XWIB2Vj1Dr+
aXdR0ZpP7uBtKGR8be7FPfFnUJNRN+77wJ3tyIus0rtmIoIxnGoimyUsO8g17WRr
Gvsrkky82S9dgmSI8Xg3oF1EhcydpZyhKRhpQzDPpJBLW1uiSC1MARF8f/1Yao7E
bt7uk63YFiipn2atlD9t4ex1IekS/TGXqjdL4xNuILJu5gjbBWQdmLhwxE1X7c3+
zZbE3Jtn3whQydbBvn/E3zyMziR5dihWd3dbFggYVnH/bFswHkt4sSuiR4k2kTfQ
3X5VeC90mreknEq086grQBdS8HEnaL238EtCttryUMyyOvJBrSIy+Ba59HMPHv8o
UimpRETJVReC1vv+sjl/emECe7894xSKyIb6WM7CGLOR66BYRaUC7U9giM8KlRyW
ihFkaOlqn5eX1GfN1JnhiER1v6kg6kbWJQgWNFyj3TP8z1Wsho0FCZiR67aiMXj6
0dXEItluJxbQt2vqEoeyjRipYwLljSWK+x0WCzzz3jErQ0ZW33yK8GFU5QVSuOf0
IvD+qygQVbq/cFdlakf1zXrGT1UNh/yoxqaF70cIKw4cVsxwwGemS8zRDPhNSjp7
fDF1fRnvxRtk9uo99N3vE4824zMHyd7h212aZbFKNuq3l3RncOPbkUuUit+S1ajZ
dGCrkwNX/4tJ37lq7Mzr+BkmQjQb+NBHHkcHMLTaQW3o8GqIRRkDDBnKtl+psEZu
p/8nvr2vDcIL5jKFPOQ8mD8aMR6OXOyiUWjI0dqQnxnVcZSKka5WQTPlFD4l+vA4
nbwlMSedYts/nWpGa60Z/Cr4ZaPtQ/C7lTBlJ8mtt+CqGK7B6YY/hsB5MPT3RQTT
mDsjIcBMPkR3ycV3DtIM1kvA3C0ji33QB9rEt9igFq5NRrDSSAsoksDHBLwJWlxi
abnga+3GGTVxe/CtghRyPw90ltmbY/+OZk35SgiI38qVqmyQE5Q4EJ+aZVFH42n4
zTUOKvxOiEn968J+4aP2E9gHqGA1nRyjmtEeXgt47TmGPLM1zNs+ux1jWGbyYUlx
sADuaysvrTERxmeHcA5KgH+Jk/hF0ZUEEvwevQn8uB0pzmgC3iRqUQWiz1pCc7zz
TK13IdWRLCoRN3V4Mlouq+EjxN+vYjs6HYpqv4zKb/RZH8mEgPLLIW9rygl1jrMb
VHMLbZhFt37gnzK1/X8gNOtT4dPAmhVTffcsPXlnlt8KD2nZnCBVULECoV/ARl4j
xqufQLzxgcN9mPXr9LssMhyt76l9YNXIhuy5Gcg/EIbRoh1X1IYvSnbyg5VFy8tJ
AJ1zhLcpjU53UObocR7CRl43Fr6czyfZpe7ijGZMnY9iYJOoIIpKEmENbXvasnws
WaM77qr3n0MlGaNgPk0VU6r7ms+HtJSlX1k51/N/tOh8coa160JXW+HIYqCxlPjh
h2VDzCv0RmhxGvsh3Mz2BaVErqGPULQuygoCNZrQ/7skx/44ZtcnG5OhR40Zoiis
5vEbMjPSMFPm6T8HWubLnkr0Gd+pNilbvWaSAwZJTCIhpZTHSiJ+mtbltjYnHBbs
Rts/aMMl9NEceXXmjCTMxlkZSURvGOuyfOZzPYeYXHSBNaq6wCWzP8L2nzyk6oQL
WMZpzBEQpSTmIS5jLNFqGjFCflJsK2LoiOnWhjj29xLWCq3ADOMUCnYeRsDMkWEF
bdfyCs4jKwUo2JT9jzOtA8WtvDmtHr+xhB54JbvlxvSUg6Rs+HosvEuxTKDi6X5s
BAPoFB3422tLCJpq9olMK1kBWhdJPmOvY9z3r7VbGv4BIvfhjPBEe++3y0cazATx
r/LflkwoEI0wMt6iq/URMDBP7VhVG6QekB3W+9jImXu/iakhZZwtUH267e3wepeo
kaz0od8hJA1v0zz7gKaT1KzxQUZCgTyczehkZ4E6bcq7aMcf038370lEl4CjviA9
VAhnYuQ8KWN8a5fyovWItAw3YTiz/u7iGN1yHXRPKfMt0uJaQv538zMpXVjiGAPd
8w9vcKrjUbZTmiOBOPRtMMmwoLW8bJLvKtJLXedOpXz5JjvN09IwKNTdyp1dWtth
wr2558E0ucdvOAVW5LKnoQCSMPS3tolGNvpa5W/PT6Emp6lkOLlTBrV1hAovlrwb
GqBsq3jzuNbvtV9zsYyZ7UpSG40u7hHxff4fDbgYUkITBTukSk3K36Rm6FOjjkgz
VsSsQBIZFat2+cNnc9evAmzUC4/1LvdxNyReuwhKtbL21WIC5Y1nla5nvmcu8+uh
RYGJ7U9ZuCyDn++YHM+x+Yk9T7PjHnUJygWQOTY7HwEaQBQIxwThTJNPDiaGorZl
7Z9GypqVxd6zA3cmVenrxygLdxTHesrjm+SwsQrqT4uwio2mJyGAlvHvPDvI0HRO
MKBViYeh2/Yg3Pi0e4Iu62acERcMSTnH1NqnPez0OmNwE3CjE8khP8F6nzZl8wLU
i/OX5YlgYidHig0LoJurNbyIAojZpKfGQJnVCx5iAQGZRqGTv6Q403d+GWd5/3kv
QXc1phha6LmpgS8WU+cFR79Z6WgcNIlgYS9lpwU1iYxX7bDmZjNXBkznIt7+B7BY
Avwms6rs1wQQTVX50lF4Q6sUxnOsOb56/xCvpL8KR0nGlLdD4pExz1MMkdJCFEa2
VmMtzZMMq53jC9yh34kMe0IjX8nGBJ9t4cI/Hyu91s1hx+bIoRH7cJ0EmzKA4WVJ
WzDuySq4HeAfpYk1iFhA7LLldoV0wc5XYoz2AkYbDd0E1knCjI8Voa6OJndPzACD
O+6FH9rdhKNC7NX9WfGCMe1fFD5vA/S8HyzdtjQ5N4MOtvlLhQaUvVwUN2QQig9z
+N09pTY6XrGT/dteCRHHUMTX/ByUS7yF5tudfg7ABDX924OcCfY/esXEEhxTjI6F
HtwFoRxA/cUIkk2ibJy9GvdBbdcJB7fFmmsqpHfKqOznb7DC0NqIUm6ztiN3MYaY
lSPnPiw4b4PgkgHsbrWn4fRkClrdVvuv/6bkI+D8nXGI3X/ZeDA6xcHuRtpwaQN7
sceQsh5SwzmLjcghCFjC7i2ywr2cBQ6LG1GyRGPheZj0HVzjm5OweCpVUT69JbE7
jCk+AhzWKSRzh572SIDtO0ItktKmD7KhNzfwN/0PdrE5aazqoFqMW1hGUBH/eFxr
4fShgfunWhxuiiQFObY1HMCLBI1PmAXaRqDwU2u8DPC8F0b48HB+bAaCQ0q+kV6L
/0XFSyv0K4R7Xth9s3zWtw8L0V1DmFOlYDHovxxPxYsx7HRvNJ8/3GTYEtMHhqTY
IIFJdV6lNum3a4crqgJ1x5kcGrXWq+IyN0neLyBjZt956BvfVRIhSBDPssmNrysM
zaOeqQszeNqXRPrWEHJeJagJRck+D/Ob9aTk4hO1PJCe61VWc09OH0+1PUrz41oh
6/zSQYMrlOHCqS/THtDP2TEsz6nqAs/ByIBenmizVJKqZTdpWloA2mA6W+kZprN0
R6YkEJZrY/sS52WSbRR7FfJ1UnLBGw7qAjvCaJYZVkFwRP1L05PDrdcD3jHu6jNf
JCa3s3qaF9TkLrNQJZZPBcOF4GdZXCSy7TeLCIkwsA3NhQ5wC1mKDPeWEpN8/A19
TTwZh/eTECjqzIIWMdkMRCQxLmVlE/DVnRXHfhbFgLxwl/LHII5hhw1DjIyQWoTV
I26TZm2XQYTZSlQEDF9Tetl5tHv2B/pra/cp9jeZLgRrmxwPBnbxYTlTcFPTadi1
K88lbkMeDQQR+2T6b9v1vrGWqB9fx9r3V8Jr3jt2V1N1AWcCWK/FrR6e3wt4Q8yV
geOtpu7Amzz1z3URWnADnqzvCm+ebasdGOflD4QaSfopTV0nD2wyMLS29fHXI6d7
Ume4+O/VqmpAIrzhNm/8ut+C0IG8TOdvtQ17sgneMAu8kjSaEUN40lwjH1jD6Nqq
taLLrrwHU63TWg8/f8qMCojXpHg0ZjLLBaojfea26/NnvVDnzPddjcOMFgjoFBcW
4W1DbreF284N6TXcYmrfX/ALx6ifFGeCSVygHRJOt2LhnW1dd1n0rEm6eCo45d+R
moCo/GYsjH9f+Y4WTnzkPxwKFkbg7jvIYH3xAnKsjRHMjGuF+6NHPjT9LB56nX2k
5krgMn/njzWabO2OgXXWDaMN/vGACNEtU1ayo2dEMc1tyi2Xh2aX3RrViz65RXQT
ywOFkHL5hURQvYG/oRiYAmvKT9LNJ7s/vHOTokIDGSxqpzR7hR1wmRzUVvnbm0Tc
DoTJcud2Jli1Xa1al/p/Yd3nOp/OWnGg0V3J9mFefyUo7VRnHQvOxpCEfp8Dp4ks
l9yM6ENkzGVt+JdYBxSuSr0xQi1JrCoF4Hc3Vv6w327Rbzr85r/duIYxRkUnVPGO
qR42vg8y8euS91RxA8ZFH29UIXwNIfHtqXXsvwvphp/ra+EQEtIm2wfO9tMdNI62
GuU16Cgl2wvHwKup5ZS90gISbNEl3h+F3AT2GzSn6YdHNhyAG1u+aCIRdA83Y8Fo
aUi5zGNMFL6dXCM6IyTgEk53UCgRSKb/0RW0CW2wI6e+87jjfpsz43DM36BNybTK
YaN98Xnu+f5cbGO+PLg3UmfV5XT4G7R8uosCkCtu3XoEnrhVHYhOMilnaFr/yi3+
4ZOAsWshCJx7d9JDhUNScszTqjSfM435F6l5V/kCc1SJLf5X1u1w6hT8iSvGEAyh
j0Ol1nBN8XGfGisfkPnhPTOA4N2dzLbOuNhprPXKRPJgQ1tHaVUQdfPEZLE5Zi/S
ik/Cr1oeq0USvLtH9IkqAHvA/9pFPBE5HWK2W9Qo+XxAeISkORTHTM2/nhWcpLwR
8Y6wvKMK+HD1PqCfSlHm208ku1vJrMe/7+tpAtdQDMk+AkE/+YufcAQ0dPjGlVrs
CXABjvi0DbR+/VWi3cOVpeHne1Gm2BBlopJSu6i7ny4mUYhpAxLA1L/YIX3YNOHb
6ht7/ec9ZwQWLIb/2yf71oyB6RVZa2rHW1Uf70rcfoNwbBx9FzVbt19hZkUeD6Ev
lymS2qOqfAgf/vAiISGECir50OL1xszmfgyYWaV08OW8YAM5UzgRTQcrs+xp8K4V
T5mE6h6XZib9qbvPlhy9GvfO6vGAvey+mWL5+sE12RbI36c6Q8i7EmvyMxvpRw/+
Y5gdIMTzAIjwRn07BVL690v7V9ryh9vPJ0RN0GeQYEpr7DUlu0fj1DnOrrn/3thO
vIBC7GBRLSvI4m+BP20p6w7RNzbK4FQLt/5jccaXqptafPyMftUnwJrpwvR/AHoz
t04N4tqRcNejx5u9BLAiqc2myLayKF2ayB01WQ3tG7vpPRZXx/ndRNEI6sFbzr8w
8VCSubOYcarZH08SpxZiQQZaS8Gzfd0lfzGrIhZzcenFw3MkZ/JleADTpbPIJKmJ
oU11evjW6I11SCp30IinmK0B33Z7p8RVtiTgxg2CRs08qVzBd7P1k4m69sBDpqMh
bx6QA7VNdxrK7pKKPxAF62YJLFgZ6TMdnmC3eDqvdYzc3YY0ukyohbSwvuGJQPcc
bBNgiQe21pqY5c4SIIScCLY07v39stjrQ5vgjSaYkwDx9uf0khzNmzLjYBi/9wVm
Fi7YZg1OLIilB+I5d+jis5SPOqCrtmUwOu2C493JNi3ee4GvnaHU5RYuLS+mJUGX
mVc1nK8MWeME/MN0DxlarWsx3CVO76Yvpt+IinpXzaJ6r4615vHYTllWNtJ0zIrl
uTLBTy1/3Hj/igxm1DEbqEWY2vgav06sQPVkDLcln1RHlihVoUoCjYrlHq3xI0q0
B2j/lhadWxN+GGF/yF8He6JWgOC//kHPjRjh0Y5vPug1frC9v3fcdfYpQtFciCWE
yHgiVO2EZWrcz/jQ24ns/UoHxLucpQrXOIb9Z2mdmHUGIVJGNHDGkIczodnH7q0A
4QuR3tRI3vDe5OMmAxtfXuxEH19Ii19jDZ1hnG5mptbLc7dzg2V3EwxXsnJnmt2q
sqwzXikfFMYSnZ4riokmHIqLPlMJmKy2nET/DiEA5UebAyDbTkuoTLg6ihc5R2y5
u251Te6Q9n69u0qtitLxKlGMfb5lb0tyiFkAaTth6hX3bl/4cM1NkPwUeib1A0Wq
g/vOM4PQ5UI3cYxO6SIE93ewvGGFOhlRGgPeNU6uxCPLMQVdKnX9TqM1M5JIKHLV
RtifuME/pisPzY25OuIZbzrxrjUF/3vfENhZfYIthuSxQbXmTkh9B66OF4FD0L5W
yGRl9IqA4fojsXqY9LAiEpk2IvmsE/GGbzw6ZnW+sIBD1dkwqJRpANp3Lbee8v31
MnpXkI9dFS5ohgB3tCDtdlhx4jI1Q2MNqCIUFvGord9McmpXaMzlrLyhiP6BwDei
NZqtmpH/qM8s4Nl7l0jxCD1c5kmhbmbKvgakP6MEp2D12F+flWu15nKT1e98/7Ee
MijomOcE+V7oeDTQXPGOTWpnncDSeQoq0cw4uuOqronMHAzNarnd10D3anqAG0qN
8igdvaCwrdZbq9kxV8WV0kD2owsdLFDl2WLIixqaretFaogjumA20ASFkbSIZw/O
XvdtuFUmIrAAtCNPe1aVAXfVx6WR7XLhmADpFl/aKkfpRWSu0B60Isi7nPSe6p4P
pDPpytsIdNtjbWF+NZRQfd8i0zyDTo4SpJei+MkQUVVD2SlJFg5TnLe2EYOzeeLO
akuEpdNp4bMaVB2hGAO3QJvfkNwUwh9wZlaTJtAzya037XERndOkiXrPmp7pcHf4
k/U3pbVkBqW9UrzQrGO3kKwhEqP3cJ1SKBrbg/Sg9TZqt96caTziCJ7aQg6qfwEQ
Hcvu12zDsO84AG7FbS82ouzn7C4R3Tjgb/kjJ2EWbZQ+Lxdpm3KCgnWMPTlHLIoU
G9o4sI/sWlPXVrK/ZkFt2dXimZ4FMbIn55qKfiz1sihrC4LUKxQNV46GjNWAGLw3
qTjh676VS1/1c89cqxBa6uw02N/9MZKJmEejf8hF0gLnp3iDY9YvUhFOesQeIwDW
Ud65QRjQhFSrKlQQvLxDvgjFex1xgv079rGY+7g8wKGvCdAPx41/jS17Qn0GGQh6
SLTOoT7V5QoyQjmh2VAW2HqPrUSeFbrtSeW/Sjw11zuBsuzUqN9ilnM6ufAPz1VS
doqyFETahNIFS/cteLb4vYUaLc25s6UFTQQ2PJUa0tdkDE8bljcVBObEM5z/fV4Y
FtO5iSIwb/3VYJnRAVGXr6qTE7CfovsnwAmLLqteoSQbtZQ3xPOjGbeQC6pNGfYa
JiYIJGMmy6Yo6CdMXm/OmuwOpaA/WA2er7XGOFXlOoofHdkUbEFbEVhJUwhOEBOt
Br9LYmUJYBAMyMq8EmuCNcQXfd1CYC96Ds35uvmNsX8hLI7RBvh78401oB7va9QF
xqwoGoxwlvq7eC1o+9NXZPz5bWiUId1kXzhlgItND7oB0k5YCIPFNPlu/ykPuBxc
2DRI7qjIF7hYAI+xr73BssA7yf81VPJ+fmec3csfxMPpMr5gifdJ77iwCXq0BklR
PxzxGj5u9uSkvFexqT5idWLnWG4RPMa8MbEZRm2rYmWkh1AO3w4HLUDAXwctRqE7
cwoOWiWHpnJaqiKAdJ7rEVSts41kLQEKsHo8HuOQEK4THVNZWc8Zi2QpbDCfl9eO
R50s35Oa91EoqlgunHWzFuMTs2pTWth05iL2rhICsacHjb6Rm1+4PAW4CmR3SJGf
kv/R2BUVpPGt3uXKzfqlZQsnm+MDa0rPdxde7+064MMMUhh8/oz/aPU7FsnnouM/
x6tL+QCzYQxlKy4sr2KbPpS5ydcjCFZmfQlrqHDojpNL00EX1jJ1nm1lsAX1mxkG
4GL4h/g4n9CL6c9Wbp5TFBnN3WDL8SDxVeTs414TzI9+G1e523dVimCysP7sK6s4
yRC/sCwsQEmekp+FdLmVbbt0ZlV7fNMybcmNN3jWcXRoN9aL+i5OGpqCiPY3vLg3
mvl3icenut3D2yqykMSodJH5IrkruDFfoutGbzliC0gsil/2yuGGrxjc+5mV3DOC
pP0COy6EVRQlq0mKpJvLrTcWhA6p5ali3kZ34zaH4WTbMh9pkmsfB8CJBCBxk999
w1Dw4CSdOkIPW2U9R62mc+C7WZGWx8vsodUsPt6wQv49B6uDBUF1x9Nc/n59Ui2t
h81F8XJ/GOvk5wSuzIvSpUqNSdDoBOaoG6vjX99ZwrbZoD80futjsK2smkwNCe/1
WkwEHuzq2yfaYGqox+VL3QoEgkS2NMBXrYo1rv/86joopnmGSB85xWH1nVOu0Gd1
UIRcx0t8gtL3urztbIVk7rQspl02huqzm4AW1ZuxrEGDfyKHh+CTDsu+u9j35sNC
y9X65BZ38QFu+iR8z1udy1qghUIjAq1ZcidUMPLrkLxcWMl9YbuAgGdvXUA3m3T3
BvnwZHjIhHptw99KkQEXmsKypnYooIQ0IPB2E0MWpiRayPJ/Er4r5ynIj/kS7+uC
UdDcq2JcioxJ9AOdcQ/xTE8fSBOX1RqYoG6ooQSRpXV0e2BJvY4axhyr1aAoUbOu
6CyQZ8MgPsxAYiyL4xj04IQ+VWz+6QGJMF1gHF6mMY08wO3fr8SpFw3T1AE0w0v8
yf83C4NFfHpbdGeCNOEU/8+UG1cWvHLApBnb/+jU0bkSUE+4ZoUU3lOkEuvhY8p5
P7UeoxrtIvRKFPQ3Es/7MvzVfw3cIEVmDNrD/wUjTC4ng6U7JZ3lBVHNMWCBdUrp
sYD6fFpxfR2uZhUFxD1x9TY6JUXy462anZSAVlLILXH/c0JVWn/phUukUbxyNUTs
8SjwOkbqtU88r5XvuD5W9ecRbpPsvPTZ2WRJjHIlF7pRd2VPPNxrPI8DcecMB9sM
XuGDX53OUr2EGg7z8QslOh5cBZa0CR2VMZiXBvhAqpZHKOwQrZoX4wNWnMBzmZnc
m19eXTYivNruX17x7a+o38Co0AQqPiNCuDmEkt2gdeZJzRUYXzVDai++uIL88dC/
kuIhqLe2flJ4PPa/pX3B5pU1uhOnTbLJyjL3DkDW6GXpjO/X5qMOuqAGzXnHP9q7
vIAbJPeGJOhZI2l6tjk5Fk7XJll4tFDzI0xk7BCA5OsnB7YYoxfDa+zHAi4Xz+mY
el8iD5wIYKw0tsJZR71ZNy9ZX1QDnqrTvEWlPvvKpcuz/3WFyoAJ/IqVjKxpq1ik
/TS1MoDSo3iMU06loJ0XrA1oNXAbBAOdNIglHB1wj5RWvUCYD3QGeFGnO5hwKDi0
YyKKzjlyFGyr496SpbLCN8UcvwRabIpC/PZSXRw5qemj/NtgCGwLFHnefYDOJlZ+
wZ3Lmbc6x0ICAhkNu3L5PjFvoIXt0ssFIfgI48EBy3XlbohUXTc+xuHv+/SxQAmO
9rQyC7z1y6s55nYFTFT0rgadZkd8yjYn6Akw//zxJar7iOSxBQQRASCH69e+lTrA
cEctis9Um8MMJnpeCYJgi3az2tltAJrI5uuL7zijZdPDZhUstrge4NT3GyNZuJkN
L8bGRNaHrL9OvTjkdeKOqH5clS8Rs+zahZFP1hEKY33vxD5tjTtVQc0DGlX6Qygu
hG/+FOoCvh1555Obs8BbwgxPFkR9Apu8nh4jbAGs6XK2c1nckLrice81vZEesHhm
Qqq8XYIrCsoLV4kNEwiE3NwuWQuBY/nwPAI5PdRde9OoP55V/NuTvCXPHtrkqU+g
Ltc+p4y3V3OTdRZDVsesabiLBiihqgnhTm3khjzlJ9/rdbZHw/d2XaCV34MmvHVQ
GgpS5vbCs1w86gISdyRphNr/wSKzR9OV64tem0pyZTK83WjFIRZiBj/GsB8vFV3U
qdvB2skCtsxsUs2ouBR59wbwYyklOTORyu9nWZ5nxzc0EA2d/rZf7BRoX4SinmSJ
lPTfrHeQa8+1V6/JEYMFstQr4eFvKCrOpwkNqE9V6c2BIIqUjQI15Mmjq0nfRL64
0ZAhFS9JTA4jdTRQDMf21dM5BXuGxfsGMAvEi/aY+sbCOCCiZlpVSC6bE1RDJxmx
pHLbxNLYkDoiJrKTtClu5sTE9i4VsURLhXs61qG1OVCJkYQQoOpzv7BNpF72Clyz
X2L4tOff47yAsHjxFapCRU3V9yPGLm/JKbgIaKnB3xjMCBXCVjR5sJnYv5KMKD8x
e3tAmlkexe3QkpniiSmwnRx4JZMxZVFj3ccNyJcMgEIXLAaqvSmrO8ugSGOk2AcL
j52eFSyJjzuA0ZJj1pes9QUrgFY/qomHLrRUH6CWrVtpJatnuFfSJFRmIsiPzRuq
O2jefJLH1tYZER0eOD+UledVLzFfe+2o2M2balBrD95MEI35hF3cYJq4GQpCvJgg
QIJERPvyt/dPmXAidb0+UB7BV7kvNeV0MrxIokmKs9vzTQJnIA+p3/tn2bXXBaGB
kzo9T/36/XpPPPNvmm37iMOA61Wyd+NN5Kie7jtKC++jwa9K1agQT8IJWOq+kF02
O+LLuighjQnmsE5v7pjlQU54mkfS9ByPdMuzysKIuHwbiZm1+GbjsRe8HFmcovul
2LQXiH9om8uFjnPK65WD21VWLO7qCaQ6/LCJSyHqBYnbPl+UZjYgmXMWRoWEwFDY
7F9p3WcLQb90cqcm0zOSISYnRfSiodq+8i5m/Hz74lwSdXqBH0mLDs+WELeR9k1p
4/Ku8nhtkVxXtGWfA2kZunwidNShjry6fbIIgT7LEZOGdWIZftrK9Jr59Mp3Uzkm
l7JwQR8Vyko8rbkRwMkWM9F86waj54APU+Erg11KsEZl9dPEqHkGnqjCL+kBUJ99
tj7omsrMYfYB4U6pz6SWguT5b0opapxd4x4IcwqbdgNPCmEbA4lwMHIh1ZUasIQr
t0yR/A0ksl6QLZ1Y3zFS4opHQJoqzdVm0m2eDUnJzgsaBE6j07Zv3EexWFU82/ou
FEqkZXT2BC70yL78BJfGESMdvrdoHfoSPktq+EQ79P5dSSufnnAb50iX0W3+vh6K
NLpePtrVWolZu1iPry6Cx0JZ6Yx+lHVWlRZVSI4jHJvSkniEKH5WRC1Su/pJldM4
+muWJS0bR4KdTVc/NXYbYrfd/jGDvtt66IqKNW0RKWfLV0oH6hlUOOE1YFH/EF6N
NdEAseLLWj3YkU3ryCLW0oy89EbaA8WeLCpxM2rxiNCqTp/Xv91O5VcwetF0eCIi
iyDLHk5X34XZd3U8YgchXM0d8O8lZghjLWpAM2D5NxlF5J7lc+r5PL1SCRHpHvsQ
3f62fD+YjgPySzob5abMgIU/0yoTmJrJ4+Pi8EdC3XJUwIxmd7nBsQh0Zr9nzKvx
G480RqB0m48it1XVzWdfmpXff3Tr+7kGKs72C+X1CXKsvpQanxfOKJ63Jib0N7pI
2K2HHbw5PLTnzQwGWFEkilIxHglYX2bIGpUWih/WG0ZwIr/8z7lZAr+k1RpBFOJl
yCek78juxQISOuKofS8/85zuFm54gsNt3jaM77X2rIF5b0H+IXFk8U4pW0RXG4Tv
gIBJYDgyrFr8TCsimKULJTGkVjZKWobI8VQNVAuqK22htoPGUr1YjqFYB2CJKzbC
6bZYa7KIyho8ZtqxTgtLv8DmaCfnZxY/6QMIro/6R/Ju++bxMFLPkBa++OItHUx1
R6MgWVwuGsPqMdv5n1dHGWvl7X8jm+N7zJBTFHZ9u52edGaJWEV6gED098Tc4RQo
w+QpZ4MGTVQFz3Z12O0SoMN1nL2V/X03EaJHWQY18G57s4N7Nt3NbBejKqzZE3W0
5TqvoWpgX1d/U9YZh2n6xltr8utHQTyAPbRW3PCLw/Xn+WOl4frnpC/f9DSx6/SI
yVo15AB7/KXz1H/LOmlPxFWdcu3xj9p+Zv1Ksd4XlQYg4ecoajICsotGpak9BXA7
yJJjd9ySThJeSm4Ru/vAxUMb8OKJUPwcfhxVWq/z4nXzKEFpSwDsDhrVk96g4SyQ
6KsXvarCxp5rULMSPWYTOAQTY7CtguBIg2U5XIwEifG8Oy5K4MxIliyXW7HfuuXx
qmRe4KDy9owy0feNLTl3gYuAfaFRqTEzMYMS+D0Go0kFLRM8mpehVlMjhsFmKtrG
HDb88quENl+Q7TtdyK94p0cz/7Eh2M1VV2vxiLK03zQUOTqu2h9te17vc7UujRWi
OXcDi0FGIwyUuX3B6YdHQOVrwitZ0SXXFuLC+8v6YeCyFoiTWdTu8kwKamFgYBkt
paCR9wDPlE4aJ6vFT0QwmQ+c2oTyVdNO9MptnwtCP7ZXA3CrPeLGevKF4mJfcFzS
D7hQuWbKATzs4EqbG3UwnaHNuf5h4cv0LNw6i14BoN1+cW2jfJtLWjwtNer5fucp
f4ICyidyLqEoF3eXstU57VAvlJLKbqdvXuUXD09OBToWP9IlK6k+1CcOZd7jrXd/
lH55lw+rrY+948T1h7wxeUEPf/qCTjSlP36h0w+7lZx4gdVYNAAlJzf1/P6EHg5R
iB5riikzOKv2KB+5RONHhj6lochRVHJImmyZB3NZP41PbixIWc8Km7Q7SVhKPE4y
jwwaEnVlFSIgAKO6k3+MVbnGBUYRpKx/d6XAMdsujbPNljVhBLCGSj1VEcsxOX9V
D74GUAEia2NIGRAkW2Yp/LatfXFd1y8iPEBgV9CA7iUGSBMwTLBzjGwRWoYg3bSb
pcrL27coxVR1sJAqPZjGr15+9mNjToQP+Vebn+ICF+cswmAoSgDaf3SH32IlA4aT
un6yV8Ew8CPRtY7rZVF1+kaD9z2hzS+SoqsGyLDUFiJQBDfPh68qwcyJVXIyd6zv
XZpUd1kOuw0p2C4Eczy7HvM5dqANodk2hDGxT7EO0zJvBOTlOofcUCGd/3/rAMY4
v2o28UT4wQMomy3ejGdCPXI+TUaX+a4RYsjodnK6JzSCH6dFemsqwRHL4XU33b4O
odP1VDAGbsf7Ba+bP1xXjGEpigNNJN+QyqWdGAnLrLSVCPxEqNf1agNYins/K8to
Uz8+46hQFKAQ0zP7TuQMPWgVnPw4GgEqme64FtjgRDziDzaIbwVldiYTFHX9br9B
3xeeLZ/JJnYr2/oMO3EO9Hy7TpvxGSEmS9c6DF2ZlMDZRS3esGDksNTXkffhwH1v
yaNxlHnbH0sT7EDfc2Ljy1V/Iwfy6+XBNSBsx/jcTe7p6BaRUwqj2ytwlpbQIHH5
PSZ4qHhMBDMmAbQ/PokhXCt6w8EqS6btjd8GW1bhB4lSXMNvVxzYCfHFZFHflJBM
pafOhsszzRDSENRHXKTaHmGyA0Q9hSBemOJkqr5YgVW2vRU7fm0e3mvsbr2oBV4q
nA50Q8gjz+YEmzbjSaswQWiwrzGIu9B36rN4lL+RJMOK+T6uJ1p913+NOzGUynPI
HSBoYUw2iigL9qJ6NFKD4jrw/MgE4g65Jxvu1e5m80ITVsffKKJQmoY+izg7BtIo
9sEYzpQBX9Q8rJHwi2rw3ylH8gWFg/cOV8ehmiN+odgHaTYlu9owMuN4ZwTN4wjh
3Pcyhejnr1I+4ZBSz/sTDWXXHzj8WyUwRyuxUyaC2rImFRbDZ2sTRrD4MZx3tfDd
bbwz0ctBfAqUUTNOEW9yNvog/HyVEwQKNJ50p7XfSlp56A2Z3V1Clvt/k9fmnpi+
SsKfkfNqD/zVFqMHFANAh5lv1es5yD6TioWZic9d2W3m6FKo22yJCdzetNSN+gY4
jOlQX4+OpqGBC3inCA1tmLn6FYJ9L0/ax7pGxdojyaa8XuUSRkvrA1O7njNU2s3p
k/08u+7HV/Fymk0a8pBYfwyKuMjaH5Wf+J4X0IZ0iJ+z7cogMHeILPw8Wt9KouxW
U4sbGYCrClxQE/quD5khk1f2Z44ykunPE7/tISwww8tT3uNQF0QB3PiD3n9H25nR
UwNhtMNcrHAILzxUOnKInJ1WYywlqzzHEbGjwtyQxSUYnndnapCHDCgx9oFAFtyw
gp8MBtXlReUScynxTbPMSwzH91Sc8yEGWpi8gS70Fsq/mjuLDNLCvYBnJ1SrWJbx
FHXTVr+leIVjnO1IeWztiNKFe5QqehRsQryyNCU1uP9k6HFro2YPWlwL2aZ8mpPI
Opzm5Nn0kWPoVcY5py17H9ZNsT9RxsgVj3XuLLhEyE/wp/nopb0O1iXbgApTK2E7
AtEGO+DHqvSwo7Kz42f+EdeDAaLy3ZIOsmqsOqfk655qRtPZWWhTVPF1GCRbsx6U
cXqB6bgot3vkPoO2TUgx5OsseLay3shBHjXLLbBke6v0dnzp2B/3Kq1bKvdydFdK
6gqnH5XEhHaz61HMQzvWrt56Zv6oKbxYf0jvEAbG7NHO5Wkws8kFExrXgbfrYoNq
6AAJcO0oCOcO5ZvaohoGuI3RnpWfQC2WZ1CyeUGfgOM59ftc+8FQYampio4nqNoP
/8DUqCNWS5pYiXURuOEtcr6C9AAd5+upXQ0lUKDAqRP4iMwNNmwyVcSoncABZdKd
cVWCenAM0jEbz/dvd8s08dX+kRXhkzqH+Egx376FY6X0PPz8J7G3PxYzzbNLwaGS
L8oArnkK+Cyi1PZivrPsiLRtJAJ72IoqPDFhZva98ahsJJBsYw7JU0o2TLaK4xsM
aU73KwsHrRj3Ty0uclcJ5AKsbs3ls8T466xhCt832sishAC8rp7PWgmSL9Y/ZQAd
Y5pE3egF50pELWr1bK061HIPHUk7dxvVMMJuzxG8U/PlrwjwZOE5tciA53gxCOb/
2CBcLXIuo+Rus32+vlYuA4Ntq1FM5qqsIOft/dxbta5E85q8R1lU5DwHrD+p9Y4I
/vA/T1lnn7WEyNTE7keEYg0Flg7s7NuXTumFEzPiWPkLX83LMd88L/dMHGxGCFKm
hf9dNfy+ZDSQ7AGzDgQPt4kDXicOnkEUBs9ao9k9BFyVib+X4szFeel6yECGhhaB
Ybd4dAmVEHF6C1mMTYs/Y6opdFaE0YkbtS0xSSrBlJi7mMceNhnA6RMSqpXQxbbN
AYr2HOX3CBiGm1usNDCDqHKYej/7VSZVbXuBFqT9k1A5w/Ywyn79Sd9j+PwP0JNF
AuN+JnMKx5n3JD2EDkC/hjd/IhHf0WmHMmVHITH+4tYVIabKlhVKPCQJu/4mbZdz
UW+4Ss+RqXWvDa7JCwiTyFxUuqk5Eg0uQGPUI+usy7VWy+hagdM3uKNHeZvuldKu
kF+xFrh0F69XPuA1WR9Y3jgkjKFBy+4FHCOUxIhYyvyKKqnX+cceRkPfme4wzU92
NwN1eyFrZ1VAIB+J8N3yMqBtKN51R51uZk068qfxXuy7HUXDU6pLUV/iXIlZ3DxP
FvFX11H6fVhFESX/yvOp1i1mi8NaGpcfHtj+MzwXxKbG96bjqrlPhVzrC+Sm4tdT
Ly8M+B6dIhkWe9jYMpqzQ3e1wt9HNIILyN1+KdUX4f5oAJ51iJHb5Lg8RWIWuh41
eEgCUHGW1funwuJiCHvlX0/WcSV37Em5IZ84ByYOTwN71FltAkuT1h0u77KwTH3c
mvKqeFovxgt2VDA/U4L51ddgVN+P34wEKqALBScRRXVHI4dzsLzWt1Xe7gLfIiKA
F0FnCM2n49qOBq4WuJmqhw3pxRX1/SyPXyIfcNjixAfEgPfUNq5nBM+MsrQEHhu2
ICe6g+ETyt11pdI8+MukT6kN91PJ02C4efWW9Wspbn/Gshj65Fnoe6iYU41gbZuf
+fTNfWYVE8pks9bix/jivjSWzne5dAIrMq3UXIIsBHL83tD1j7qDQwK05eg5mxau
6W4KzT4aYkfe0eePzwF2RIJNlZ7AnmhRfTMzAUr9jbha8xsFfeJCbzEsYQrH+INg
Rsc/zvQHxOhja8OXm+x4tbjrw9X0MEHBJvtb1ZE80yFY9giqI3FCvaTZI3StiN+a
dG1auL6g2MTXBzXRH35ruMaoTa8A7F2iTYXi9nyO53sbnPiqJ0qIkCCPervvrWnR
zHsI2pNLA3DNhtUKHNguf8smPRNrcJ44aAAjXfC182dIr46fhIT6KxRs5zifFuky
RWkvalMcMupZoxpb2/IQx43U4JUKzc29YIkBzK974HsLmaZTvXeBFAb+I+Y99ax8
QXwr6pzvDb/Ynp7UlTupVliTHWHxxFrl8MBB11j0bH2Vm0ta18b5lCPhYj9v1R+d
qIwDjtXkMP672GrbDk/XbpxlBDfZLDMg5zzIcIr1HtEOhaAR8L+IJfk/M+QSYDnF
ZYLLv+EGHBynCj0gO7DmAD85ENvkgU9hRJqRItLfksa4XiFj2IobQznoS7QyxtrE
vFqggS+jy45vNWeJq2ubqaHze3u/FptxHyQPNOLtE+GZc8PuoKM1BmtU36uyRGOR
4mgdN/rAOZRcjHl3wkrkI8HW6phTJmc7n2mj843O8ZxrdtS+RLKs9lGsr0XgbtR+
KeTnanVMm6T9GsWlJRS6TipgAP4G0E8YaVe7Px6GK5SkLeWU/+teJt3jiHoVWdCy
N9jfw34I2cc5vhOCgTC+m3vpsAECp5cEEzWrCIp4LhC+NB3ORF7pOOitBKh5TwQc
`pragma protect end_protected
