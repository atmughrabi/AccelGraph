��/  ds��8�g�f��k��Fۃ�[��5ŭ�$ٙگ]p#j��b�zL��/�e�_��¶�v|�����R�UZj4�dQ[-�89)�Y�pF�P���y5w��q�E�%�,d�����c����M�|������gJn��~�B8;>����j����6�X����Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9��J�<����f,D�"(E�@�,&N�lſ��S��Ui�+w[Ê�Dm�1Y��)��tQ=�7P�@��>�4=�ڈ�3���%Z:�a�ǟJ�]�)�Ca�x��n��{�(���f�����\*v��bj��Cg�།Kh�l(��:�H�������_���X5>�1��N/m����\�P��WI��Q�yuC����J-�rɘ�z~�UOZ�2���Sv�_�e^\˃]��]���u�=E����u�����y5�lTXH�c���4�Y&yζ�bX�y�����qO�W�_�����g�dWA�e@�d��L*n��U���z�M
���Uq��+�p���	�⸏�1�Ϥ5:p���
�;F�و�Ϧ?[Xp5�=m�}"jH��x:�;#i1��}We0�l�&.U��\q@l�:�Ν����E�sk�rh�/�#��|A�PoH�i n|�����# v�Vx����4M�J'���?����'��0�q�-fؗ\��\���#[�҇�q�a+��W����"r#�a���SI�'%r�$����h=c���N3I��ߩ'� �A��F�{&�$�q�h�t�ϯ4c�Wx�4�v0�Iu�Ԃ�0��p_���v�2�X\UQB��ϲ~��I�p��a�|`�ə�-a���T;���64PSC��N�1�oy�į�#y�ǻj"���tƼ^W�1��a|����>i��jɅ5�4�m�ŎGm&��
M�\^�n�p���#�I	�z�f�Z����|{S����ٳ��lހ����r�A 6��I�'�#����qS��nڣ�"1�jlmY�u܉f��������q�������:�h��B|䨁��D�x���r7p��E$����dK�E*YgD�z�Y�-J��v�A�;wC�P}����:�_N���ƺ�����@�%^���1deɡ�hy�Х�Vzj�3�]��Xx��2�T�f�7�̃ Z���B�c#)HǦ/C����E��S�uz��v��vr�w3.�����0}D��F