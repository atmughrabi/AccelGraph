// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SZXFDRfG0+VnVHWpiVqlKZpqbtB7TcR+Rd7yGozgRVwP+y/G1NhlD7CiQ5lNtw29
2mnCeYiQMQZKaQIvE36G+dc3GGvgdwqa95UhnrpuOxm3c3iFLaRGfzRBdzxVJzQz
Im0uoOh5vJs7SJxXZBLJ+280nripBpXe+4kshWSzj5Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8080)
65UmKMCCPjdLs5GfYCkjCdwdzMukjXYKFJk9rtaN+RAbXQ8dHR3gp3nqKAc91ANM
RMoiZe4unXRP74MQ20jCqRM01zJ5BIUmkukkoTFHTgM4V2Am4zX3TyOXlmoM74NN
YXAbj6pG7ds3UGNfp84ocdxXnhLtToMu8F14QYPlCZ94AVI8Vv92MxY5jHBKbqVa
Vl7hyZyF3ZRCeGCL21Ww/rCkO5dKRNielU42vzBTQslBQIaW9RPn/MbGXKhFEoTp
igGu3D1ZddiK++v/hjCQczvoDbTCvUIL7fx36jgGbjg6qQd+TnbwT13kQjwxUEtd
3lUbKzlXC3e0lih3j7UiudbsglRswR4o01vrJJrWO3Yz85VmUMWg4hS4xtmvc3CL
0BrK+iOFmYvcSb1XslWAtkDqpsewrvrr/hk5NbvXlviX74G0LakTqQSn4GcyntWC
MdJXdVOIcHWS9shd8A1NC5m4oSeEXaOCpVu/aJdf49jbksUmSCZ3L3aYyrWwnTim
raWF2jELCL6yPcbNVrpFpvFGSbC6z2L4bREXQXQnnA2bRIh9eAItL6wRocg+PtsQ
7MoEgdx0zpZQ5OI1d586/Ud6G1UeHrJZ/wl9Qicn+smfM05ScV833SwwLQ7oSLCh
28exv2xyRjj5deoOflJ9O7QTznuYqNleYklAnBfMxpqnNHjLRoP+UAPfMmEPVpHR
BikYS/qEn4v/cYe+3790O0RrbHkPq5OEhzIoBsh8rurlCpKQPGD+gbJe/fKCIGbb
WBWzZD4s7CiVcYypSo4cd1d0xcQwaBx1PKzfwv5vQPKl/cTVD5u8Rq2K8f21YHHR
Xsxvqdb+HOQY+R/ZIZ9uBsqv/WgMitw1B9R4k4c50EI8GLMROFgX7anyO5W4AwdP
5MLV6aQV6z4ShjiI67uuYSMaxrThvEQCM0ukwXQ+nuqEgbtMEimEelc35vegTzyF
B3dDlAJBqJrrAnxixCQ/RMxbZ7TtsgVhZOthYrubvDLeboj3/l41Y1u0TjkN5SWU
wOl3sd9iZtRGsfOtV6hljX+LwbV9MzrtFrdXV4WwlQibAtcxIFCZS+w4y6+c5pL4
FE2h6mlaNv7FFB9ZHDM1ERWB0y5stt03bvtTQ684V7UebEdpq0e2omhRPk+9lksy
5sCANBrZ5E0CgUy4uD/iEPAoZtcbUqqxMzPFTJL1KL+gkiIA3TT0iDJTNKZ0oAPr
3csqlAtKqmQkLGhF9qJXTf9ffkMbbKCa0qjU4ObFkFahZ3B3B0N3WE3XQxmo4z2i
o1XXE6D1TRaejdcrzt8LniSvLhYhxf2yroAAfmCzZ7hrsYCRh2384jnEjG3jIa7T
YwzQaxNxd2LUg3NZy9HaSEhuRxULKz1lNkOisyc/YGJPpHHsX+DACF3w2grZpYN9
l2J3ARsB6I7bs2eXhkp2F2qDzDP3rYFICJ7BpEYJMhauPXj1Z1o/d/xWxKoVDxUg
aWno1GDSijADqSk1DUMLnFe52BGm/e1T1u7spktLusaz2xXosRQn0Wa6/wRcj3qf
OOOtHKENU7v3KnXbfj32u6RVuWr6+Zu/ialRi0qwLdUjkN+GpFYXRHSGHl9M/XmB
Oere8Oevzge8xjZ+cvqB8Pzf6/xYbPkh1XA9lgVchLmjOZ6p3bQHaPTecYZvqoNt
KUmt1Fc688h9ANI/RVvZLIxz7SOskdX5D47jBDqMhQAASu3ZaSeU6UbqHHSwSog1
q5RdT/IGVDnqW4FnalmeECWiJzwJvNIQfN1pIe0On0aUzvZMx87vm49qUNb1/MJr
PEiWjIaAKk1E/BsJHaNlRRwWtxnINBHupnSODg+W1s5+xclV0L8VNGUcygB6kWo4
Q6OGfHPAda35POLvHQasBQbyL5gMqBp3rmbFWvIuIX/LejMeNt2KytRsDcpguEBI
LHFN2M8n90tH68VABRfacMNvh0izdF2uAZz5wfy5K81BHn1ewKln3vi3vN+aKmuC
p71XrFtLLTs6gL4t6t50dVHzyvhACzwTSjOXy1GA9UoR1p40+gN25jQlkpfsxW4I
xx7xY12cIqSW4MlUTIxZt5KCfWhKSnFYSJAark/350BVYiBN+3spuQcv7mftmkwM
n8UkWBCHvHVAucVSuRxS4v/vH7MuwrifxyEEcXv/P0rzCUeIGtucNL/FY3Ed4/i6
060A2eSOw7kd9xC+fnYWoRtNu6X8zb0Qr36AIKTUHfyr2Zf9Ik2R2qSodJmIo8pz
WWbjtIJDsQ4YwUIF+0ndXWseXM5tSnCGTVTSWckVeRKBXkBsYcWz1l/QjV1clyOY
iFkw5X/OYk17QDjKiuV5Ll8Te7tTS1Bqq/C069+YDJw4D48hynjsRDYAgOF6ejWf
GiyZM0xRnVMwIO9Fr+yRcEi6pIdwgKEr2MgYtCMFQkegWls+QKkppc1VmMcBauss
11KnwOAzZh1h/0/I+kqhcNK9SXXGcF2lHsRCaD3JDhfhwhKFqBhgz5XsGd7qEAnK
2oFyjLf1DMP4qHu/mOGUJt9QC+r0BVaHchbCl6MplIdI3aBbOtdZlziwy/jBG2ap
cc8NPoAbyhQBsjRkVgnEjVM4hPWFkezHvHCONnDwwYl2pbi8tAKT9+uHUnjv1Qjf
/HQkoE+GSfyynQmTpFABam/7zkq3P8IF4YCEQwhERy0IXzuEIcqTjzLDGAKzDG6V
onxXwitY28WSkmJe6P+PvNrzJWhF/TuVkAkB6Es26+gENqm/uaZnq961bQ+LVKUf
sobzQHMz3jjl6bDnF535aKsiuDdekVu4Hl1cyuuDHRvJ1evwwRbaZVrwvYdqV9ET
E28V949vu+ad+IYbwuflCZSxWFQmLTL+ho3IGdchCyS4RaFez4ech2Tow45T10/3
jpxN3wO9QYAHImszU5URWTENSRi9Z8cYSHF4uix8adBcC9tAlDiwQHD3t5G22Z4r
+8VZPYEkKh4qsuMF+VGwJrrczbM5d+72R2jfOYKY6Ev8VmGlCLHtU/UpENwZAI5P
h/g+H/6GSK5N/d7Mn+Pl3QWTYDWNrrRVz4zLRib1XXdaWYv1PfjFV1x9PuUHQYr3
M8m2LomzcbR2L0RBl3v0nUWlc/56TFo4oVnnd7uaTTyg0lXjzPVOCJJXzeF/RSOX
oMKQTSQwKoRezTiGPjIklIczJmtx5Gaw+srSU6LPmx6/+rY0e+0dV4rr3nKfdrLE
FLqIv6tWil/em+iS6XxIrbxKOPTw7TDr8IBapftQEDM+DMYPhdGNSkEUwusXpvms
DiOYgvq2SDWgdL0OuhhHX2dUenAvzeUtk5T8TtZEDq/GYs99cIBVOvr4xtWPwcZR
9GIClQx7ZzTSca7dXok9VqHei1/YaAZl1KfuHHJ/NL1p1xIp59devEuck7s86iRr
STJLgWE1OHgSYiNH34Xlll/D8MopEMBLLGN4ZpesX/GycCjLvPaEbsxA/dGyrzIP
8A7ak7B7flmqMftjQzuP0r4ZVCidSzMXzTD87MIO4cvA7vg7TUo9q1ZUUC9/frds
l2VMW19RcKnp99qUwAbivX+dJ7b0dOHFiaeyn3WoVii8UigsKR7ihnQplWnF6mkW
OmZeD6Ov+DRreelOaFPYA9Vd2mUcmvEUy/RBlLf4HFVZgN/d19pMyUeChk+D+AIJ
uuHNeoSqFXV4HjvVJwrJPmbAHGCiDZYsDNFB1bbNR9DJTAIRn1KXYqdDCCRPxKjy
sZJI/6wi4W2XWD33l8FD6WUUai4MjfBVSdoWrweidx9Mi6J62CSeu5kXnAei5tzm
b+tD58NdNkk70itnraOMRckoOiOkyo+dSMzZYP+RdnsBaJsDZpnnvmce1HYIPQno
V7vECl6LXNemBPH3RrxclTGJOxsXuv6uW15mGFyLuHBYTNjgcciXrRA5Wg9OGDXs
1zq//n7fyypCUcwqea2+bRElkeBSFjpmZZLAQOrlEDE+1sqZ0WbcQpqE10ktIi+7
j1rTsW9cr60g9VoOIErzOvZuwHPcy/93GgGUhJurEj9sB7Ou9efgGPrDFh5HTgAy
aLpqRaNnIALIpkj712Rbm3KiwLLPpVyT+l/0ddeVMbLJPWUiy0PK91vswD8WLK3g
Ecdi/G0ICCHUHBdP6/WG/+Go+LFWKjCxJEH4kDDqBl9ZKyfC17kCZEdmab7x3Qri
4iOdi86NK3KYoo5h+qH/6kIzc7F1k26MZ1JbuB+puNJkZXNHKpOGLKg6UASPBBlD
lH+UYQtd5fpBVGbWWLvhCjtZt99TreHXqx4kaV2mqyr0bg9j5DjNRRMxnkX0kQed
TotsQs1DVx0Z2NV7m7YACQHX4efZjm8A7/s4gkXpM8MWQRUZ5X70GllAw2UU01bA
3SEZ18BzwN3klTvjZwpjNaFoOKUFXKnoMfmCUHdvNuOvqVz/GZsYvB57BrP/RJnx
PlP9EZYLwqPrE+IXZHQ2iBxdtp5/c+GdNzZx+Zem20AQvI/9QpRhjFlValiC7SMX
Vs1oUyoCp4CWNq4Jvx/Ls6UW91VyBimvA/KoGpGCbFNtG6F+QYIdyaoP5YB9ggZQ
tbw6kqfg4mAlBlYKspQI41clM6ybTZ7qsKOLjreuPND9LZvLpt4g3KUO9S6AXJwK
SuiYwQ7FEPtoai1b4bwR0zyogtSc+rB9fE9hVDhUsgzKUEqXwrTrglO+Q0GqDFZ5
a8pFzLc/dD1y3141TquZ+3YvwiXHbNt7rLp1RU4L8tgY41RVSPLpHGiXhi4vsu4c
efdJkK6meBW+IpqBvXj+0g5lyHqZuZG4PqX1ZYy9m1gMgEZKWdA0aOU1NlvaEFba
gdWWDJGZXOKdqZGFmIjLjl1kNyPsMJyhziJlZgL1V6yN0BsNxHjy25AW4lLdzNF7
4UTmr3ak8ZLrg+bJ8X7ueK7GF5otq/Ytt82c05TtcjMv2F71o2fcadEmBcLG0rCk
T7QrqHEWTHM9OVlg7Y6GNez6cCt8K5SsVTRsb92gcYxRL/DV6C2VHlkZcoBBMKM6
OhZtupHnHqR3PoX/AzmzaX9fGrYX1ivDluJIzN54QQSfIw6imXhJub0ce/wYdSvX
RKoVmlwqW19Sx7h5Fch9TiP08XiFNyLdLohx2lTTGQy6awul2DMztEQ6iCzdlXZw
0y0RlcM7tr45JNQ2uTYF2H9cR6TEThGxjJKt16YdClPQmDL6qA4sZBTYpFdSIa4U
yWB3MRsrmtK+YTb26LjScXp+PPMfXc9GfF6F+ZKoVgPchRy46OV0s7jGZb6ylQVF
Ya0n5ulTdu3bZQR82eRroS2ThKyN33r0tJunWRqKdtsKskUVfh+YYFiols3cvJHt
UQwSJ12Rhe5synNq/FtwOVYoMipf1z9okq3ZdGH1frgPpkIo68Vx4FqZ0ekuGvYI
VFmzigYzt1Zkqk4qsc09l5ptQDz4dfJ20z6jD2wkcmasHhsXAMArCp4j4U1wSSwr
PUnnFZ2QEY3VXRjwbCqLDQ0jWdyQMvapVH1MDivGxtgnUaegCcxlLIaL4txLXq6J
XQlkjvecJI7ehwy2pmb9pyWaKVkqT9siVjYjhEtAFhqMBxQNBDdMTE2v0OTX3H1b
btHx9vVPDMDdxRF/tcd22oYe1W+ptA959L7Hn5I3VWWB/5xFTCSfQSoG+/VBcfAP
U0EHmnB37JJW0fvEVXnZaTXhoOUr/IkktUmky1IEwNDJfE95hOACbH3yCTP8pV+W
EWJ9ibzItofQsq6zPxCH3aUpnKYACT+jdy7bODDPgNU4Tpyu3Pos6dqieImzezeK
IaQlB+RuHt4bMvVRyabjaQeE9vOsSo6MYhqGGPbXx0nrWQdVS4Iyb3jhON4UHoIf
8h8noYaQq49866PIWtrPFEDBzWytZU6ApRp/2QT/tmwpFjB0mFMCYyiComz8KTDl
BJfZpm0BVUmNRrFnpMz8NTLYiC552FjzvQBZvaxaW4Prkd7ywtWPqd+tSqUL0Tyq
cKPSRplV+YedhfHR7oDkbJpj35LzwoApSy4x7cf3Ra6wSeutu0IoyLlnbmBaksGc
T+LsCZ2pjveuC809y2x9C9C+/DsNwfNbeOO7lZ5c1Yoj2PthAmzhvdga4iFZ+VKU
ffsnR6rikxmr9CHdFJG1D4uLyNNmR0cEyzC6+RVCrs/YnG5iyGJkLKme/aq7PkMX
BKRFsoPrqeon87cTIuKPxZNKkBQH+dlPPtHELdTC68r7NsKCbLUdSjeG3nJzLwMG
WKf/UqFiQlcMBlPoAo3PFf7CvrpeBbMcOe1RYmXfpDNtEvs59ETGN9U76Hj++eWE
L//DBoYlTuPB0ob56w3PB+DfIE8kZ2d9TmrtgOKnC+30anVIsH6jjI4WIS49c8gN
CyYcdsr7Qa5EPZmWD2VuImwrHRteYcTv7StKwJ0kGQFU21xRP0xOdxvNitrknDAB
tdo86r7+rFvLdgpgEJDk2XgwnQ3F+2RghI5Li8tSLWwoyo9n+5dRQBMfCcTVQnCI
eMGpUtLLb9XFJ+oAXDXzZR/zMJ4x0FiKcdhPg9uXjvK0551tp4Fdc/l6KPrllyZu
P5wHM3rmZi1IyL4Z0jYmEtR5FxpzjmB9/8ekXvgvgiWaPu/LGvWFRBvovNzUo/n+
DNdGwAhiirvipi1rx5XeP0zidvQTyuZR3n5yL/TV5JbTY147o1aY6mW8AOw+J0d8
iZH4SC8DUhqsKpV7oMBFq2HvGbh90UepSX7s6NHkCuddTx2OyEvWwjAk4wSEUpQm
5Z1qycWqh++Qdl0iJ8Hpk/BEncI266HNY9iHEQvslpci5G4/L7rX4cB78lzVCEDc
/nTrLu4NSHcfvx395wG0DOBmvObSwnu5NfQHK6dsN7Wdoz98HYlSSDGw2yilfswN
aaW2JkC3nMY0FqRJu9RDJxwRbtuWXFkiAL/HG0L567j5BRQeaCQZr2nag0Ul99QZ
zxMyLlUZM1EELXOwzrtALSMqhmEeYFOjGL2Inr7T2pV/p/uezlplwP2nX42GI4Z0
fuhUt6KuBQ0LNmHR0rQuP8He9eR1M77KJiRQm/3yv9LYdYp14UwkYU/zm0B06eEF
eXmM7MaSCy9WnaAXkAQV3y4UmH4JW/fCFb0AXpp5cl4O2RtaUy7VqQA8DZIiqp31
RoQRZaeIr2bzDguSdg8TCJ/vuQtjHdaGkJ6grKCuSZNDb2eD19XwWJ3II3APmc4p
iDKx2Wz5Iz+ghuxEl1gMJVryF1r/Al+tu4SXw5KJSTKgyLCYVFpaeVT9vp8x6q2R
F0SeR7ifYJdzDjEP3iYzhHhj+oXb4oxICwqtclWyzLhfT20l9IX1mLwQBlgRrpDj
XgxcvRI0/mO2Ed+jMPYGYtKvPm9zPR2makVV3/iBQAo6a/uByLlOao81RtAxLbbe
ZNR7p1NvRSf653TiqXQsgtloxlSXSc5P26HdV2rJKcg9QOrJzdp3KGY/p3sXn7bH
IR/cDwXzqJC2RnkpqiYgoMMlolEr9S3Nrx6usAw0wX+pwNH9nONWo1iX5inrhOS6
xx5IAg099Yz4JVY1Mb0noHdiP5LqtszHxpH6zjLD/2cF+YNkXZW7D7y0O7pIIAWD
yN/Lxe7BgEg2VEQnP72kxjK3h/UyWBoxCJh0uuAekmEpgozFPBI+TvRE7vDcM7Ng
bMejnvN4HjXKm61hpDmITVxXm2U8Q0Pb7LkS36snvroic/RBNbShxbUfC0mFyxL7
fidtB87YT5EdHKTNT1TcTHhKC3h/SHPlruKxYB01atf0yiiwQcuTeatbx+30QuOJ
vZff0YRFcRA6yDlGbV7TGfoV2h1gbbIebtICgxFdiG9FQ2r9sCQYKH8O/wuhqHXy
nMd2QPggUHZDYAyI3KM+GyiWmlW3BTvsrsUjTKAnF2a7aH/2ZBLcMrsV07doMZVj
WO6ZDYkc5xrIn0KMyDso2gP/iF0Q+JaUVvIvcMDbRIIoB9HALLjRc6rC7VssJ5vg
pBDK4ESc9Xs29KiXmxaC2YsjLP3QpzsHDJwscYCRR4i8nhQ9GcqBUDZ/FO/nC5ep
z4kR0c31kkWuqB+MyaVmzMYAEhtDbF+zP6hiWLvkLSca6q9KhOjfRw0rj1K/LyqR
xvKEZUBupqQV2/jyUaP2rU9UcSvUye4sZI6hL8JyRbW5geptB0w54VeexAj5AQnJ
JmmshhsqYhcfGkF8lbn2uIv39thqfrvh5tBSsT58OplXluE8cDL/EdbYX09yiMWY
KZJ08xAKq9zuB2FDL8WQRN+OfoSujDMkEYiU0UC9/v0sUJWB8I7qyjOX6Kr+aFfF
eKnunpZAqh2Wx/6DGRLc0jOo5+e+D1cnix+EZ0K9M12tPCjW5ydj8XHfSD6nW9tf
bIulJRudx1wSnIXTvVbbJl3dIdBSkGBSymuEn66D3LcQNyHyF8fDle7nhXBSb7wv
UApJQ+hAwnfBV78zjUITUvXlxkTaT8q2dcEohgeEi8x0RzxGVFluy3m5o05U4rYc
RAoXxXhA7PYnArCJK2fL5FdtBIVSDrptMHFg8nxJ3KwX5PJKsB9hYBeT8LTP8OQK
vEVuDzecqOnf8L39M6hdaN3TcByZQtA0NvwzqncpTi0ZLeIw93BGymtbe0o4XfzK
yOrBakekjX+C35mrSjLrA3UPzbqaSrdb9uL1J9RHVf1yAXqld5clsCVZxeeumInu
U+iiebZfBtOSOGGltTXEcELh3BxbQhL1zJfaTlj02Tk+/nGQ2jvq8Lv+HIAiyD+O
WsVfAJIqNLJUenwEWiGtHACSPhTy35V6U8APzUCH565wesqGYobJBKNfub+KV32H
c/oNdy/7YwQKrzKiRwRKRA86oGSqloR/h7S1ogm1bNhfrkoyrIKkbHEDIDT032tZ
b+ZRjbXBUYgRNhACOoKxSKVzFcWILrs6c+a49f8O5/rLiEOz6mB7khwi+M6DIvgj
3Y3Fa2hbHiSRSD4rZEXPdHHf7fYei3F3ZYj3DizgKJLeeTokkcdo/FgfbqXwS5/M
NUGbf4zfsguyYzJnqSP8cNTBSJQwHSqTs+YQIVptFJtq3qYOHsYv6iOwPVScdqx/
bnU9FntN7sBuubBxrZ9qfz3E95rVZ0Z6hS1XoEZ+IIfU+m8D4Ndsr7Xz7sDXSien
99/PaIO8sKPWqz1AAhx5YCFYRuf6jUxCufaLwNHwEiaFQ137/nLm/3Q5h0320tqR
t3R1LsWlbRlwE90784rHe5HVlg743OugqKeg7233bnez2sUIwcBi7Kp3sMwpN278
lvJYKt4h4kELBW4O0Vu1N6niFHt3a9vaFIx3T9Ea3IIr7VHP1aSmX1V6eVoNLb9A
6M3a506ufgmddM30ClfMODXMDT7EgvqMeOxGzzRWwTXc2mXs4AGnKLA5a6dUr+ER
oVId4PRUgrY17lztgPZ+WTS6Jsa6odUHVyKdiRQ/vSX9um8v/wbj3yTGBSY0fEQ5
jPpKfvU5VsqgWQSAulECjp7j/PTRksbse53ePUpDdUNypXyOxO3Pv9Y9EQfbfu3k
BVbhxU/LOFzKYjeFYBzoDjlikqnSWXW3mA504SHVljMTelCC4P6apPsDOBGToyuY
ZG8L+QEUceaK8EeV/6HTi4ZCQuhPHhfBWBXoO9/kbC8MiBAOCVhebHkbWPl2iGTX
Bkx/umsyQ7zwR8C+PFkPuE2tdhz/EzDO6tCRyB98jW6v3Y3s8xwfrNK7vXJSlb8f
6tyVTRv9So49T9QDsVk4vEoBGE//o7tYlSD0XCz6ouKC2Kx9Dl4CVVvtimU5ca/T
bDnPpNunMBXn7YBCsSEkrgEU0Xi/IX/LczIMwx0d7ex/dgRXmVOe+0QRwEwB5hGs
ZlXJXT4OVVaXjDBM4St87QChyaDXwzxAQHSS+IZ1khHYdsvK6tjDPr6li7KCukAI
GOPmnqnvirEJ3sKb9a2Ozh0+BjTqWv4uHGmHg7nvEDsQgNjC0HGdhPjCZ9DfIFQm
eEVUySsulfcdKXJ+oOTnzYCG4Gvr2RqnMNv9fdyUAcJ5Fz43YwcW3+A7UZ+QnNkY
n4cDf0jKo7w/1rYoM70wja8LFDTNacNzlh+QFKn9Pa6aKMfCX0AQWHv1hX4JdAx7
rXTl3ZJ3/qCcVUarD8ThPa9zCmunk1DOSMqKhnqWSzFy3iV7ka76icfWOOk42vvR
Zf7S0cqQuxd4qt1ZxGPMFrp2pdYlER9O3k8TJd6TdG13NLUx8ZihKH2HkgRrEOFi
AKP5bEUqPjDQmtdTSDfj6sVQU3W5IM+xZzJb8SgTS91Hu/7QiTAfZ/i7JHZppkq3
7tQJjapoU1VWtyt+aCJxTYI7knTwXiFzCTfkUTkmL10aOs75RYYxA6/qcmPK4w5z
+JzwnawN3V8sgjfEi0Lx/JX1ZDltPUj7S8E+Qia+0hOhp53QMIsjH10vNZSQq7E0
37+Mp9wMy6u5AU6MDY1zyFOezTL5LTCbNktguAchZ5xJ/69Ug0q/ixTiSlydo/4e
TbqjA70ZTgYzwnl68HdvyLMVMov9uZOSYzMVwmd2fsQAHb7oOGLQUwlmrfgaNs8o
sA1DibLtIW2PVNjeh3YtYyq3TMUs6WtF82nHpK7n+ai5UEwKM6TgGdfJZfrrPqd4
fB6ZX7fZmskiv6xr66qLwBiZ/PoqiOW4/SrHtis9cfY5tXl9X3uEotfsQTJu6bX6
oP2o1ZcUB/6Jb5XCG2TSD8UHrEby9WTLgx9W1GV3VA0yvDvLwb+M/aGJuPxGgO8o
RxV4TKaCJKPKR9xc+5cN1XRAOYMtnjaGh2E+tzNmhQBC4vaITykFkuacbO6P1y4n
bfp+78TxHWjN79aCoyrr6g==
`pragma protect end_protected
