// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:45 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XlZa/rSdb/vgOuOFD1xtM6jx8m1EK3TMwSjYTKMmFmmQ90ocQD/8cWXMn5N3h3ng
RaMOFYL4VtT9XdOLt0RrkHJn/YkX3FKr2map03TNuEWXOVVqF/X0RMgCKnZL58w6
CIfKGQdB0qo57KLDJMTH3lhi1+sfcnl8eUFQsJGVt5g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21184)
EQE4C8bYxASvPZZEjo6F80Ll0zQ1BcGVUSyn+879pMUYPQQ4iStDA+avOtXm4zjW
Rufm57AvmaeUB8oXGtBp2mv/fJXfeOnEPFZ8Nn+w1Ldhar9rcyz54yFO1Sf3H8vD
bcdua1Wi1t9GObR20BjU+57yeB64Xyi+YYQufbqKbajbrnUUBaWTijQT7gHuJwfm
GANetz40cvzrxBeJ3Xoi5wNLxGBtR202DyH/Z5rvdcuASNTCFYmBM6nk0dvplUb/
pPCvN6fnO5k8N+kUS/k4xWv8PnRIYPF/5hBgR1+RtpD1RgoTHzDx1TyULRFTuONS
hXjMkeFqzW0sig8KXm7XYQ4rBAqKV0+BqV+kg/D+jzmbeddiUizmhxiJDm8T6yLF
BU6gZ4mIuCG8PGWgmIeK4G3tkNma7nZAKU5AGZdOJvWR9e47DwiocbofY1grOrrl
9CtuJ3+Arsu4pIgBHgKQI1bUx3kJXp+0NmoLG68MLJj+VHDrWY+8yFm992bIfsp7
ZuMssI7J9dg3/taxJGupAHG3KEiVHZqudolmQrwEqTuAoJcDb5YG1WWiYf/i5a6Z
Rh7n0qvn7WweKS7DK6bvBfj6ndRf7QDRzWTTysCRNuu6o4KbCegSdygnSE6fJG3F
vqAsXX8k1MQRJJvWD+u+SNOoVcrRV+ycm6YNFI9OKinVRXelcuQKUMCf4hiI4NK+
ZsyxztQxF8Frv4gY4Z+yOAKPXo6b5wQnzPariK/cdfYGTWWXhKKtAtZqqcB3YPrq
/54E4YnWd11DlU3rgz/fgLDkrALCs/4kTtea5xSEe703cxTs9hK8w0VqluWU4GGt
Jo/BP30J+uC5AYXsWaC621IQTva0HJYwtgOZCnlSFVFQMa9u9N8SEvhFx0xOP95r
7NkZVPkoXVEzHSAEPc2KUT51hLE4qZtTkd2+uGA1Klkj5LSwASY1Kyd4mUmnURbD
BUuyLYg5w3SNsQnizdBiB2UuGT8Ac3zbJEweghEo3AJL+vOGxSPOzVdqN1GjNkFp
w3om3dZ8ORBvkbHcVfxVaqOqQptRoRF6ipDoCi/u3BTMA2NY7x6e8ziRM22coawN
t3wPVL+CnZ+Q2njp9aQbMBre67uykKjtUZRfqpVZgAt20dSATXHXMJwr8icQ35w5
wcxEejKexzA/H8u+qM5wmIPri1EoN1+XakE7w2pPoKqaSzFtBt16pY/xleH9GP5z
NwukK/hRJKBQHTG5Q88QsFpZeOHWEuPJ/A6t0IZRCZTzu23RVOgGFGem3f1cG/6Y
W3vNc2QHmAga80zhJSdzbnA2kplsLjLEz/WFNDhty8fdB/Y/FB2HeX3wFuJP8N89
qG2OWHTSSp/8m3UCKr1OMmq+wtL0nWxrlWeKW3QxbUyUXuEVrFSw3q/GrFCa2xgb
CSqeoSpAvzUwZAv7DeNPL+1yLBE+XsyNGokGy1O8PoP0zO5jaFOe0WP4Hu1bOQ0Y
rnf20GDfU469qBY4VRKwpq2lnU5AttoPRXkIuMTjlH6Prcr56yAB8un7gZgnQysy
0QptofnF6v++3jVJGFlAPMXN0kAIg2rt+n9LxgO3r6YzxDXl+lwRumLQrBUy+s3P
MqGbjP/qVIddEq7vpWDLPnf3l+clA0PjdFyvGUXF4D/ghuBgMZ0h/erVDMerNSxg
YL46XHzcH3FCzXxSQYncR/Lcz1mE1BxP4vovQSu+A5GZBhBDcSTW/CEajJk2p81W
J4h8T4IeXJMDUo+Q+BmZNaXo15PsHvjuDR+3FClJBMpwbfvPmLIVWZUyFXVpzx10
3ThqxPJLmOsojDI6HGfUAJLB+gg28thbukspRrg1TP7b6Dt0O3bS5L3+4TuqgSUK
ZxX8HmY/tJHUD0uld6BTCRUyu0niB7ndrZ81OqNrlPlq5rsvB4o4Vx8oxg6pWBvk
JBzp0HrSKLX6g503NOYAZOSCpmp1skm8alp3EwstG/1+/3W0nEH5iyWxetATFBZW
4zI8owM2ZQ2uiay211j0pH5uxDucMIJG3Qsx4wUIakJ6DZr2InR/WH08NqL1AuQ8
+JpmD+v/HgmVvjGi8rRHCtyE8Ui5/G6Rmz0XCyQoeTPryOE78NOxoT8oFzUixmc4
1XA0bgcqk5rLqFz8ci3uqmkzl4Gjaw+HNLXgHYwUSsxCYPTxYD2VSu6lCHMXu3UI
mhTawvvR+JX54knfZfnKL5Q+TSymbUCn7tCLy53n01j5taX4E2fNxDSLlhfLWl/6
KkQXEhWAvbEYmw2R0MDd6k6Zb0UIr2ZrcbJhkof2IRZaoCyeyaeLhES7TGzHP+9a
UqulY9QChwfrQHWl0b1jF50W8woIJclqUUIIYZ4l51cg6T8W6PBlj7mBGgq+7Kg4
/+eqjGyDvdWOcIXGGr8A4ZHGmRjHIGR1VQvHolWlUBK/+JkEdlzCb5M+qXRX/RvX
QYKMjHetlS/4q7VljC2YCmYq3a0g88QSD4nsvPxhfN0iHDcHmNBKm9JA2//PAg84
PAR05sdL+DvmpJAMGhELn0A2v26V252Qp4K3qlVEcxsIzZLfRlukxY4Bbuka5vqF
MOz2qb7nA25KDnQbV5rnPjOAWBzMAVMJ5MQqbIPAG55NDvq0ukenO9ZZNguuJuHD
BaqcKa8nvbvHDU5cUqtrnaz9CvXh3R/rVKLVv4zcJxdMshcGm1HLkB78hz9x3s+E
m8QtAoy1exEuOal/GSoocSIfye8VCp9i7S+f8tmcpJvm60LzeJ+rBYW70u+oVLES
VkuQW3FnbPSt98/sHD0+oEiNAVP655fN90i+731+tjA6S93rq7s1QXH+XmCn+FdQ
1C45QTq77njbtEqIk6lzPG0N4vvwvKR0XHeO++NxMKGbGwed4a2UGbDRtwWJH8S/
BnQPCUGhMwg8G3oSJQwATn5FiNf44LzX5ikRuTUbuB3fsuE3s2yErXmVYKbP2UQ7
/xSmLGdX5Zuu4PQ2sCaVyrmiWqes7NI92ZRpQRzEigojQcrrMLM3AVRhwCUYMMgV
wFKYFWyoWUkFMr3OfAfdaeN70btDCW2+bEjwFm29SW1NfAAOrJsvuym4kdXbi+UB
8sj5KpwScq2aAufkdiU1Y67slC5/rAILTnwBtfKoqgsy2BY3+uzSRpglpbBbjRQA
5pjmfeZ7pm+W14pPLauDvnaRTFgwcONCmUZ0mo0IesiStJogT8+Sp9mFtjmDgdFd
wdND8gJv4vyUYSYG2glATfKcj0OA1sHC9HzQK7WF+0RWCdl5dNo4tFuVY18aIfZf
dba8LSShzCHxjDHW5iBT5r2AJd/ZNPmz06F5mqFNKtEThSDnbVabK7Ka0bblfbvW
31WCbbKA7+TGZf3K382rcfhoIBgjHdiFR1xM1O1G+sLXOy22YoewaRQRHWNBgoNI
y8RnAl4qDbsoaPfkvMM4eb32mnCeHr40M488eeK7unqoQglxcVMt/WdG7vDvmmdZ
jp++CeDcXgLeudQjYEBShVtAFsoHQyifJNdTJ4QrdSVW8mVOOkS1F3qKJqNFRmvP
9AnPKu8jj6CV4yXCPL9hF3JutGNDrRb3WFjD+oxz2tXzFl9ci/XsG2WumPIixFYR
awE8i8ackdGMBSinGlWFCGGcK7B5HFcZskbw12ttoFp8xTO4TlKqD+WmzOMOMokl
I8XTAx6e4ejx44HG6GhjBHhVTfVgY78Di43/ueTdJYsFRnP7y2pKvkZfb9p97WOc
PcAlHFaxRlua1YKln/TIytdnIZgI9QewZDk+Jadh63Md0tNGalhxyqG+UgGXzeuu
cHTjNcX1waZFf8I4uF3MrWICZUUibd+vZK/oOqNrXaqrys640yzXVV/54btqS5wq
LiVrT3ltdzgpFFiVWOXsRt244FZ7UQgkZithPZ7M+WZ0DLYB++HMhxalrA2RL16/
FviLShdEVMb88JpYAOXa0kbYZTtbFd63kcFbov5JA4ha1J1q9lmVuvuJIGsBkyDZ
A0LBrVssHwFxj1ctGXbT+mm/w3Q6ZWVNe0xGOYzsHsibUWvCXrbbykqQwnRS6NzK
IL+8+GZ8PSlZXRod1irok3xFNnkhQ8+Z5QLAC2A+LZuW0fD1/2wIchdnltUdx30c
tYhbhhcmvrbo/MoWLDupipGMu2Z/SrtoHiYuHTlZB8PV76kPavl5vL8Z+0418kYV
SOwK53uGBJqGW5R/QuLw+un6Tu1AXi6Y6TXsyFT/sLf0OYu0xHeA8p8JB/bfyiM/
+/iz2yks2iyPovuJzWd3AIg/bVMEvjjxDkzct9YgCeWhPNlEqRKkuRPnqyvbzC2E
G40SxD8Pk9W5sJAqPfrG06Q46t9H1zQPLG7Um2eIQVgeQ9lo3ruofi1E3BhREDYJ
QiV07Csuoa6HEI4OpzIDBsjqR5heD6zV8Bi4c2lIoYlvqik7OPtUBd72XqXxt7tH
sY0ONTJ9OCkeE+haV4xzFcTGTtAmIinvL4pl7zqS4sf1rlC+mZX8561BlX6vpl3U
Ql1fE3NdCGF0RgnLLh79RbWNg2RkqaUTOVoOhk3fHqV3dlbufIf2Jdkh0tmP7wiE
dui2CP/hsOWB6dd2hSA8Qw9Erkc2WdE7GmFsw3wfbabw1pVuPQ/InhwztdKybUDW
DzA7X4ZxeScwNiyckF1C8APKmNP7oZHkY73y6qJvw1eaEmVArwuPASBFBpnd2o8r
NGDt3YyTL3QSv93dzAAl9furGJuwA1N/K5+fd6Sydj0PPLR3/kaW5sfYhwpEV40W
G7pao5glXC9pgn7S18Qv2MukFhj/S9Ig1XEMpLFKKSbJSXYcwru0xL4Z6oUkWFuw
QiGUJipvq36wPKbSfXOX2AjIRN39lOc97RYTwWUFYRM+p5yQdtP2TgIV594bMRkQ
80WU3rn3SPGBR8QbGAxARZV1j8u6Dtcbddp5fcXMFmKfvz+pJcUnzUiffbAy+Zah
GutW+Hz8xSLrPrlg5vTWp1cU0CryN6eEsN65hoCAdHRigBSAFH1YjGfpnqaF/4It
ScEd59rmo4+DhpTDCRW3Y6wiQhAmmehXFKZOC50BGZDdXtpxSUrkaQ96OChDJxeU
MW3hj+AeOOssLDxCUaswUtWxMBsbXGjx6HysTZc/lRP7XV71VWqL1QpNQcsxvi2c
QXbN8qEicz5+G0Lj1Xvbjc4eVLpImA9+8xFo97FUEnwtjc/BDCH8IjBtAT2AwiMg
K4V8ywXQkOvc1o+TgWMYB0MZ4AKrWXQA3DsWGyPIuNk4thw1dLTOJuCJlgP878iP
j7RxPX4txQFrcK6iIVXqGNq8lNcxmy5Fzf6Wy4G2fzwNsZMqlghhsqVxgXAMjCqq
LRKKRPyQkRWRHsxr5G3BPRHB0haN3x2IVLAe91mt0UbU6q1wGuAb12iawtmI+S6n
ByDyDBicWZWrnDUWjjnGdJv1HeezNZAmFlH/WbYTdrPWpdbF0m1UTBhbV35mH/7q
/GRT1f1DIMy2Qo/sjBIEZ5nkyPcF73KoZ3pFP4Ss1l0/5tRFMnDvNaxP5616heA+
4xl2yp9D2Ph4E4aNrRj8wHOymXOE+tu04UXUk9iZ906AOyzzK7z820izC8NLmrCG
ih8EcEp8qJMzzZLp/LWbsc3R8xWl1LIM9fmQjw4Oz/BImWp8SU8CDUEpdfxwPvXO
3No9KNJEp7ypQ8/kmqTQPnBXUQfWEe5MTZYrYtmm4cLmEgbEV8ZcMC6z+hN9tyA2
cYRHE/KKIL3p+41jV+JgXh1G6Fe0e5hEbygR/ZpQ4++Mst0VjdY1yLb5ujL2ZuTk
SkL5dLN5bdSq42n95ivv11XEGADr4mD68ktp8QOi/UJNf3wfcFHEoHeAX/rgYKvw
leQcAaYGVLCJxYpm5WAGlZTggITfZEGx9D+mwWmYsBQGn6fMV6J90L5ou6TwZ5VU
1QsBbsVScFW8n2UURbbqRKU7Zk8FcpiPLN1kAnUNAL1Xawuxpi6M2l8lWUW9IL1h
MzV3f5AisFrNxhqW8sNifyl/Rilg4EIgN1rBg5LLdbP1hygqBkfC7GtvfFapO9gx
arCpJgn1AjhYW8G635lnk8FRoFVyE3U9QZj3SGGGyH+S41Hd2V+o5iEqfTbq5ast
PZKYE3hJz9zPGS5dkEdbt+32rsPBRMQ7bjPmLjA7vK+pbpU14vxOdDlLQBu0ndI8
xfCuLBGPaufbjKN4oCN+V5Zzq/9xrKLxDMiRSgPDnJEwhJaO1O5V4P48UtUMLjuO
TQQEzBRIb3OgKs1C14VVXlrCm+PraqMjt8TGN/S4XaNuF7Nc/rsQkxX/TfFsug32
+0MQy/tTWTqB/Wr/UqcHtB+FW//xvTYYIDqGsdMD1kCJNcp0H47gcLc1bmJWg2y2
uFfaMadnxZgxb7+F0p0Uv8akTQJEeRaBuhpaP/RWtwGcnWO218CblAG9WLh87U6G
yPfjJNBnzC3awBfkTEVRRvX3odBGaMJSYPLUogv7MlULKvi0fscVhTi9wW/bzS1b
QEvvz4cjqm7keRHz85JX+CDH674mA5NLdlaLev1cwy7+oZl16wpSUImhTETGrrvl
c/VxJi35e08ruUex5g+q+tItv9bEVhEepdRefXFq37IKIKVBFcXQOnfm32ZTqH4Q
klcvf4Lc6S6bZfWohSkmnr/1tc53EBNt79KOGynHGeYnb2O3U8U/J/DutIsjf6L4
8Pn1EppImxt6D2ZPRTyLetxTUBlzw3sA1bjpaR5MxsGllm4QZ8NCfJy/ZjHCBb1k
qmVMh5hQarcZ1ZZaeiE5eyi2MUaPELr6tbpmwRomTg68PNiH7x0MsCzzTvYQGglV
t9xXkZa1/CwhEeMN/VxvH0MlMoQFtTbeuvHYSyADW2Fb7tg6ovV79zLwSoOQX50R
woUsmIyR3aD5SDCcPNKk6b8N3f1zQWDlGOdcitraOK86amKSnda0sT14lYvMFzKy
5HsqBymOIK5S7DM1/IYeHBTLoetbS5dZRJCsnzCQlgyvLVmHA0qYdnPSP9WsHdFo
XgB0DmDqoOyRhdqTMNaU3SUR/iS1UVyN1+s4GTrJK6Ew8vWHN1EuppGpgz1ybGb+
h40QguwO82Z3JL/BLF23E9IN/Com888+phUWdVHeZmaR9oU7Xy4xWes+4pjF74Cw
rhdSojNS2/hgTz/qu1w3n3horTBnOG+y0j4un4Frvv2KPhMiOsMguo6PNiTYSLFe
4lfhFccdJHBurqvc8Guxo5l2rbJiy+pMuzg3giWyIwwB+GlWdyroIJMMaYo5poJQ
x/eIdH6weSt5qedFQORPUQQnPsOJM/cR6UUxMnrw70W+sJXEdjtYQEjVIJng66yG
FPmhOA+GTrPGYGs2GNPeBvAqCs+B6Yd3q6sCdhsJhM+6GJfCzZHPT7Vi21iN7cqL
jWkT3Vx7uXoFsnV+jan8pgb/Y+QLl34fQcgJ4AMM+fHwOma6S1zm3by4r2eUzNYf
hvTMA8sGs29CIqTpSzKg6GkafOGMLl1ZNgfIXZ6H44S5fQTtRnUev22Hi8kybk0Z
g8RmDI9Xev08IEq81NhPoOS3BZYytCqwtIbiJTOvaNlcqJ7kRBeYUdihgwW2cl2B
xWSbO926ifFUYb0GM1NDSeZYkM7L3HGZiQfE+JSPFYoru4pkTB9h6NWXRdOrvGok
D0qT5tjFmqcpQ8XDD488TIvQkOdJuGIP3+tlv6HhFxpAil7n3lJrAKeDyBlHRn08
HGMB4f59M/GcSP5QwYXXDAod+Ljv132+7bhR+QpEYzobqYrQ4e2KLc+KcKBeNhdG
gLUp4Bg0zTbnwnpmCZSGc1frc4shDI2ohonamyXGgnf2RiMspu7E7gYhwbGmIme3
MpaxxhaG/fZzK4262y0XAG7z4HDI2WHBD419dkg9887Kg3xlbeG0Yt5P22BpKa1B
LgUZFKPxHQXS3bxgegu+/zleCNpWmyvlsagJkMLRZ3Qrot7Nz0igCnt5t/5ZtKwz
eVdN09qWbn4ZShBrd52oraaszjYPzFeJqAv4Zi6Nrzn0jjhYaVTGfeGljjQKzmZR
/IXHvY6brUd5sdP/nblPRvvJUvdZ6jyrXDAkQtijYFR6YtYDvWktLpnCWyUWsypn
5AsG2N52ZNUJiV/k2jqJxHIZCGKEo46k/1dPQx8TZpMnHh5c5iuixlLOZ3p6Pwsl
1aqJTgmW7VqzQzXsrzLKdFL4BwH2cCl9yYIQR3Qo6sWbcI/sTttJwViLrpDaVxyj
xcfLn4LuDJjmwU/jx7RcnRuYcIlz8rqdX/YdSW03j6LPFmbyyvyo4+lH6NPTzE6E
3BoBs1oziLs1vwpvo2Bl064261+vxmDlSvge490gLJ70I/qDkb2S1xZPa8JJ4A+/
7UzDA6KnmIM1kWc2lUeqovqfDX1+KVfdQtKEsWreLkhLxP+knOyAF3UUtWgbY6e1
NMmCLpBzKMsC1K75j7Oj3swjISIyo4I80qQ2QZl5LQdezPeeHxg/zUEl5aK+suDO
JIq6/JnV5tHjW5c8amIEn8XVZf6TMSCq5fOWdKB+Br1j6/bDvEpF/PAwJsf3K824
Emfq0JtcwhHcY6abrx1fKVvAJHVjF01XLHaUpcmnY0iwDT4DA6G/lZ/VgHzxhFmG
5C92myTbrEiElMOKQKwolbIZPip9UQk0+5GFkDKeS6ZIBB/vAQ3ogN9lZ6nO0BJg
rWKOI8SvWxPKr5qcxBk1fHpN9Nq9SLl0rdfOL3+J+lS9r2WmylN4gxaQk8c8w9gB
0soKSNU68IRLaNX4YTQbAb4rxWd5zgoQAwoMvvlSnLI/s1Hw16p9TdDWdJdMpkzy
42Kd56uKg70hdlfB65T8sCx1kDOWaaxn9+QUTsaq4LHnu2+vuLl05jHcvtuz4vcr
iOzGITO0EptJs/ioU4z7PkHUAHEVeCyo77on1sZEP9OuOpE/91pUGE0uR/VWXUqJ
rKJbUditQrToAg7ij/kkFk+P9QBcGbV3u+YEel8pEO1CS1gM8llQjVfYLE0rjmQo
mfcbB61AdQ3LYJhuDDBh3WgwIGWGCt921AR5jDrNwDurPT1MfYiW0WSGTDgrXg8A
B4d2LLQxiF5m62QQXEMXdHgvcjdEhYaTjwuuq4M9zQpxsE+XuVEpi8senDkTm876
nRH7bz+yl62ZEO4ek1Qg375KHGdqTcmJ3RzMjWnoqJ8gEo2AxPZWr3TqZUST4s6J
7UjxxTiNh8W5JYrkHrFnR6PVpqeuTcBGThkcSUtX23NGoCZkfkgphk7quyi36dzn
bUKl9pZTrhJ4wTDFLujbSifwIkl2KIgu+iZ33q82pGIuvgZKmrRTVI7PEnH5nHmj
4/3Z7hxQWoJ33x8i1gmzazhDjEQIrgjmiz+SYHUKUk3uWbQsU2IDpaBOjbzlcwqb
9PidhVgtAUmAPJe/cnIThLses1ODfvOAeu4U4v8P8/tnkLKvlq397uOvDpK0Lq5D
bXi0FquLwZqcNDazTjELsvcvggS2N4tVL6WLnJFugsNnaEOUcU3sXSe/c2s/6Dyv
c9fRF32oVrbwcY6pLw168KfZtdaNxGwpWIX7l+Erjp04n2S+w9qL1Hxl1pbikeK2
4P3B+RKLgv+A17z1/m9/ilvJknpZ/KoyMqdO+zGr3o6WXa9zx96kp40Rr7rDaQ3o
IDo280i59tdQ+vNsJRzLBFHBhQSePuD9/2woLLEpO2IM8lLiyqFeMQ9s9AhSy1bc
a95Bz64x0ZKrm1bIofFMcbEjIIqwZ4yc6jOpJsXw+D+9izGKfljwY4o1HSGZJWM7
VnAyez6VZQLMPTNa+FqUZDhzrDAJ/xDyGEHy0fM3h9tRiXQd6nLBif6tks4g6EHM
eWU7Hp5kRL1rB68Z9SxMdoLdzDjFvpWDoZ+hx5gjAT1SSokD16X4EUhf4mumOL8d
vR6nVuCokVzzdRn5JbbSZccVd+RKnUpwTnX3PSJjdotI1OZPmvAUUS2IOOXnxSJY
3s7BGXw5XQNj+bW8LllAQu7/PUfOPOrCBRLL992KIqylKpoT5wIsxrDOeM3mv9yZ
HvAGcXs/Tm447YGZqwkGR0uSM10ifSkLgke5bYYrWit8FiqsyRpdXS/sMHeDNYt4
j43DvyvdcrpIW5AOPA9C0rtDl34g7fUTxmuroFuTPhcIeifYt9yL+mpsz6kI+eI9
z22xl+BoJGDkmXbeVI9obe14PnzoB19R2J7rtXI8VsfAKfqaHOn1dTOgZzU3ec+/
AQ4Bjw7/pMNJqEHM7Jp7Fexn9K7mF9YFNUAjtxJ/F10mD4cOVAojR9zrQ0wklyIW
b3VNbLi5OnfU7PCIeonu7pw2z/8psXvK71IrM1883HPdg3nEyrETQj40k0SFoyJ2
7zTOkhRXyc+Ml88MHz4ntYQIoTb+WG1aO0BlvNBMc0QaxAhD/iGvY5R6W6db3ucr
uPRn9j4g3GaBrAJBzjelqvQpYWY5B2QdNUFmp3qLG3Db/Y+nqPk1Mi3F3ERuN1rO
+ZwyhbzjWG4jzgyoRKkTetPUT5RQmrxZA5jB7sm3PYSgWKSwPEbv+QUigblKuX56
ENyVwVZL8r+wioKkjBP3/qzl7Xt7FEvCNxTqoXyAQOE4G9wCAi3vta4HoC5eJtI6
g6PS5W7H7N20dvW0hCyPtvLSqSQEmlElBHyjOA9mZey/dY3ywOe4CdMF8xCAcE83
YnFQDirODlGWc+b/KeLRKs2mz+SDb/CtQG15zVm5PcMsc48t0/RrITmpHb+/St+A
3LnAbPolb4NwE0se/ufkLdFuxGbszxSS3d28DHAcB3GBnp4utNx8v4xvt5c2mIPp
m8Bv9h7zBkMEaaLc0szD0cCE6jxTRVAVdOcgRlPS8MsGD+YGl3mg2w3wHCYJ4vTK
cHn+ewXnVEMiPZOuHZpH7j8xQagDLXIJ7zIJReZoUxu55tn3MTqk3bdMtltUk38w
mb2l9qFlncS2nXuT+wTHhqcMalI0sHlyklwtCXZIBQWqmlMFTp1VmqwTWCt71g36
eghdeXmOft4GJbA3zJBBafY5pZLwp7vdcA2yo7YiErzUd8iKLUj8zzns3PdmExma
O2YgCV+y1qpERDBmGV6+k4ipdfsAKvmPO+s0994zKZJdZOgAedQE12q5M10jnpSX
LvGfgz1ZsuGaT7KzXA5WlOIUBnWve1IbOcGwWFaoVX6hJfWVtRykGkOGqiEci3rM
iWidfxipkjWB+xN06siRriac3/C2OrnDCQ+gr/UI9Fy0vandh6m36PvjbNmfBs/5
qSLaykqk1tzn0yH/IIrGtgk1BfWvpe8pof6NQMubFqsrAtSLFglVtM1wuxOElo2x
5YKx2Kw9BM9fOjMHBhtomnu5hYCjrZZwwnJmuqw1H4omvVZjYtPf+FG+FRyj74sP
X4h6tiCm1JLioCXBRNiYfM9nL3OBOD+46unm6QkD+N1N7WYbvajxYqWfbH1KzZAU
mYHB9YPFT4ZVY/5aVXIZ8/Y0hy0vLTaxRhg1bEza+CVGQH9g/Rz30lq1dmXdMjWu
fUN1i9hNGctZQH6gyCiwEPJIrbWYnL01Mj99RWI80O8lPdI6bZQoTpSQB5CxmPLL
spSegSirTp4jUgnuKPmhIxncOCKPZnY97Jvh6cjzE2TiD1xnYrRCzQyZsDp4M2dv
U+sKgpmEgg57ZnPiCXxUXQMxzsLirVmoBFMGCisYZmXyh4WM5BAc+EotGHybA7Dg
xiFtvsvb790CVzNnyZZ9d/edMjQu781SKocM/tAUGen9PWmH7Ak/3bD8cxU2f9hX
/z6ppWMYcSwjgoWMxFHTBfBvdh7aOqBPUxN+oHd9yDJZZEeTQTuK1ZShu+h6tO4E
i5smvCe9414V7Ym2oAQvUiCzc/Wmwzk6UtlvfY7xeEz4Wd49U+8FPXGHmt9C5UGH
yKr9NavaJXULFj2CgLZerX3Rr9leUqq0XudZyx+NlLshCaBtGjctwA3VBppwE29q
JOlYm1enybvIdE59b1FkVszhvKRRiJmtTV3FGtBFVen3zAACHLrflAcBKwebZrHY
yvWC51KlDeCskMlFFLNFM6+AWhGe0Q829kdGmrxaorexuRdFlmECOP+kBpLMCRLB
IyOco77MewWW+u7ZzlywubKqGp2+kd35PrKizgw60gNk/EDSFBKxE5uNoqUsqWpz
ERyXuM4BwKlLa5p8NiQl+fY+jor/G97Ntr2KmUL3c/wWqYiVtRFsh+zfa5lVvqva
axmwodDHXbkcTXy6Bn2CEKQzuBJ7wPniMYiJQVvTQCNL1cYGlABCkKnMpSh6JkWL
mAZzalWzpLzs+oRSolxSBqeh75G8ddfptrzQ4sSI/DVXGwoqWT3vG1XD2tbRuYpO
maeO7igiTqnCwkKTT1dLJCF00GriGcCY06bGiaPoXZiOJdMB3DhkY+P4PpAETbsq
16lw4b7P71rJxGxBanxVpnod22AUoVaim5QEOLnd0zCf+1OIPPvSK2RRAEOaRrV1
ViZOZD1CG350yaKUuFuewExkc424lzLPG3zo/2isPhHaHp6LCUESsIXbkcYwfUIE
b8j5HwrSCzWpRzocdkBGd7xPxZC+4TSVA2gdf5QF00GaUgiqn78bs+Ii78+YcCD1
Y8Xff8tFJnhbiVop4lC19XVRVgKnwni+cq7iGzmQ7bXp3dvJZLkEDSRh0cygVrjY
CBdc+sQgBFSI9eXg96yJOxu6TXEs9oVHcIsh3IHlRqrKXofL2Pt5utRhuSDfLBCY
qsHdwULYsNpgb2K6vWnRYczVpXDS3RQdUW2BhcVtBP80Rs8kxiSExETrFlrP8jWO
2UxWfaiioOycf/27/bIHy00JirzBiupKJ7bQ/HpAxobIqfucPiolYXdCrM8RX96v
INaJXnfQHCL+Oji1ypcum/sOgsFJ25frr7P0qt0DxwjyjtdFr7DiabiY/w86bKLo
qzuAeiSMpaAPtLpRuLahJaFX8JiJuH0Rsn4Uilkv6nvnEWJ2nkn1+IS5UZ+Jk5M8
u9LjDUZUaUe/KiOB6QKTNqpDc47PM/XBfRUanFqPWRRgY2BnT7hABhYi5UkasNwF
4+t0oyS439JstjpW32y9vLIyeTAJZg66FHG2+BZRs5AzgVAMIIhlq3f/EZK5vgYp
NADfhdPX2WptZtSLnJZwEbcfrDoeB9MfD0eBoKkEViffB9uPiHm/sHzH0iM0pBXJ
zvrOGKJ/jrIAN6OzmcvNQxMbrJlP3reNlCUjUiYkDxSSMKFS3FUqgeMf+aKZ7INj
DBwfjaRriQJ5vTpQo2j6ELjvzjKARh8JAznUnhCeWHYkc1bu8FA7EbnrXhc749yZ
ucOySnxTFKOfVNNcPaKelQvphDm+ERbBBZU2Krn/dfJQpu/mDLRg0xXwro+JasT9
aOCjryo7zM9oJcwLCn3S8HRijNKmgvP8/xMmsBESATLBdVak7T4wPyeRJMeJN5hp
+8TAGhVBm9SMgN754Awl06xDzyT1WUyMTXSXudU8q8kyWhTbZ9CIKebn0kBCBHlT
dT2I621i4pb6VTvA8R4F8aPZ6rm+mx1y0s2tGGkVgaTJ+8uy6Y8RtfUIzxjlshif
0CwyHNqgfOqNG0U17sa6YatNccHd3Xw/JI3irMJNaHFg7K3BCm3GydklDkUj/X0J
RkjIKZvbuUd8mA9ZVVuI2UAeIbD0JvOR+om9jRPlhie1EeHU87HMAbH4OI7yFW0m
mLzR7yKiC1dMxNb697J9NqwmoPaPm9V0wDMpgRgsCmUHp7+FdZoclKSLOYt6p/Wf
Y3p5csqOanW1iSvjrhhGqgCSF7048xqKDODoVgRUAoOIK7DO8fxP1gjDrQ+l8oUz
meWtFbGFFSG42sD4e8PQoS1zqERV0KEGHDbAamZH3+jf/rgQKzsyq+ZRnqz6Finf
FlMgzrgxknKqKaldmkJNGmJJdIsm/8zVpgzS+JYPG8UWls7kuxGSi7sYZBBQSpg+
Pew+czVwCxYQCQshDo5nW1Ng5RSuuKsVaUwb3JJgzsb4sOmLbv46h6eHS39LKMzZ
DYyn7Kceg3MRDjyw9kC//cLp377wUwMztRT8aJJmYy28A1t4Gxu6IWWDttfGM/K8
55of9/2ZUOpxHVRek13LKRq3RyJSZMAf25AJRBp7X3pNf1cGKfzIzYS4NNWghiaF
2LvzSDGSa8FTKIJWdDlfuSKgvVz0mVltBmDKMC77OHjSJRftGLhdUAzOJAC6lZmC
GSugx2iZLt/zWL+djP46nKnGH+HegG5yf6XIcqXTWZ45UZ5aw6wp+/SVBxDyMHgw
jP7/GuvB2I+1rzrLUkRqXWzIb5skmPk6pTH8h2ZwJgC+YTK182vHHHZCRv7nMpJg
GCuTE0JSzQpBrdXyftJcGAdz2jTABpAyIf+djKdvzFVa+Q6NevxLfY0AxIVcvjDd
IqKJi2H2IoUPmalHKhNWM/6fMWJQK4fjBfPUoA/4AD/WtT3eQNMyCT0pCGvkMPKA
6J99RD/vAoywAff7kVLXhvsvDXfihPs/5d2vHd0sCoq+EdU3F+5GnGbQioNF7ZEQ
jnF8r9RPSPp+KRgARoaWFd/IH2X0D/GV55vFjmz457d5iMOmBLAGwRNpXujgr1RW
1cdhZXk/+v2sSb7o5iCWOetoPPX3nNjqE57mxmhQQ/eUlYuH3OyKKxq0YENuEe9V
78bdP8G6+f0FExyi9+pV8fbnoD36qgtbrLxVF+jJGPbqTQ5BQKJBO2vUX+I9WgC1
bpzN/LTYIkLU0CJPgQ9wGr2gW1sGOGShlfNASUgA9pwf4W/hvx4cOuzAGqwODJ/B
0bxCp/oWoc5iO6QQFgmdHihk6CV9kvTYRNT+GCfHMD1/ESe7+JRFt+N9EjygAud6
92kh3Z0Ij+w9IHds5F2jcg8/3xDgzQd75VWrQZmLlhp4+wF0RHm0HC4U7G3Gj+fv
ogAldwC0ki1UeTdRi1G8gelTnkEVFtbomxA0mICBfHKTgIO5TnPjQMzOElgyyngB
tFFKhDfxErsv2LH+QAhy/mEhFAnUd0nguB33Inghk+xvagduXB/nUgBg3N75FH6s
//tzicQ4qH+vhAIzKHrduQnGiN2ZUS72duQH8cFGZECSMlq/OK32SngveXAw5NFD
OjgDvLjNgz4jAIpOQZhMOiEXE2bL9+KUklygKTUvFnCzzvMIQdYpOwupgRq4ZxxJ
MB9gTRa734JI1mpBb2DYLJGUsjpoEuW4rkcj+VxD48QTfWjIEzYcvyMlPkv5z2C1
ErEJBPEf0CriDeKKp2W88yN1u/gXXYRyFm69vJqHLlOKXcJn21PWPUNkdQNlxzSl
/+oUuYIVH4YXlv4icK1gSIqPGzRUnrCLoYw49mbVo5kZlsU5pjzzc5RzmqL328BY
oghDwT24ab80odvalYVYCjlZASVy0M0/EO6zEc5/oZcaRLnNAJDrTrdQODMzJozk
s74lXnw/kVOr8pt3EtOFLuU2Yp9xLAhHQ5v+EIl66rnCUNIbT2jhcismb2LkOSmP
nWazcDb2fiL3ysEZtMn3GQ7APMaJRdEpTNEVkyudFvOTCDsDy8CqbmqwQ3C/1pG+
U6cLLsJU8/NCq4qbjLuNRpqKfdidncldzclvWwCUl5NI98A8O+NBJkS73PLm/m3Q
emxnZFWSLhaPgCxTFbQs98dG/yhiydHPdw+TwECEjBXDiF3TIhr3fb56lO5Db7lo
FtPc9wHK4u7Mhdisc16cSUHMjXTAvcIUbTYITUcLXb80B0mbDaQu7qW9u1kDsdPe
fFiFL+/s3BHO+SoXZwBv5YetT7Bj9ReEtoLWRfkOb27ufPJ9GnnsQMzEOKsQMC0g
9O6WEPh7ra64yLEv+t9p4/SXuCwC52wb5wS1hhWS4xDS2IJfIL4iKZ6aEEQ3eMkS
yIa/1XPfEmvML9d4T8qxQ2FVpTtwPb5yXx9ribrlT2oh8Fl1YrN+757dPeqhSh1i
kco2IK7NRed83YbrKH9aca1fF2DvOKAs3mDG0tLw+52VvGOg4knCKDT+zGvSGIut
3ghY1IAuhZo5iiyi6TQrNKDmSJWmQP360i4FJXR0Uw2OhInF7fMU7JfUbigR8wjv
sXcb42J1mIZIBTM12oNFAJ7+pIFlcBbdWrS8yq9MFY+5l0s4jUeXhzIsABsxBXaI
D8Mx39IVtvD8sN8wyDkQCWJl+l2cCXFE4yNXnTstQ1Aj3ey0pacajoREA3uOVUwJ
TgJEbikbAR6n/wyT60gGr2IP7ujKbcf30n+/TV9peae0nzJH2SgCEDQLpIIoMkMs
RRNjtbg8TrYiOYAGp2vSMSDfpLKcB848Op5+3NkjuwruqfpWGVqlX2jDSvUSFS85
AryG2o+kLLC516JyJ1UJTDvHri9M5n6HbD9jmNP3U209dSyN1GhPAd6iz8HjJF3r
gm98XALbAzM8PLAxfRArRfIZxZxlK9PcuJ4LIfROfAjf6i7yVAftEkAI2KUL5tr7
G6p8zjQncbuVo35mv9Pvjk3LJW8Zb62kVzkh7W9BOGvdVCEo4N+JCb1NtraOsWTF
Cni+QpJa9mrZ2FMpuvWPGGkWynVOjCvCGwHW4vPTjOr2r7WfMgs5sYvyNKUlXldZ
PTbvqTgf4QVAnC416b3YHnAkLWXrU7zPXQykfhgYiwEwgH0fFl0N7H8Ue7vuphDa
WE01/A7dbLlRs4ZRrSpb2Cj5Ln/eRkzcCkpEUGzwPXuPt+29xVkAes6HonKJx5W7
nMTBHIwsnAfAUwbjhDE8wvEHWPaqla3WNnKFxB2qrEB0LCPi0is3dVxvtG39z1oC
D2C7zpkYuy31NK67hTNMSx3ZOK1crC2uR4Wi6RAG/KNomquLx+LjXbo7rjJIkPSX
9NNly3/6jzYKr1F+ElH8kJZzKMfnHSQXgbNLLItrvBoEs7BjHRQCzOp904UNca5g
4J91edUt/nqYBsVly/++hGpTgZSIEKgry626+YLkzkjpea7JfZ45CKw8Y5mhUjKH
dTZG43YpxDAD8P6jFIB2VVbY9KKECEda/TCWvj46gh9tIX6aQfH39rS/QrtJboYV
5WrZoMndS6bmU56plrwD9/DWGjLGCBwO0lPbOTfx2Objl858Ed0NKGwARLCOwiif
519j1KMRElM2LSPRgM/YI0pulSoS1d2VZIau5NJLEuYMT0dyBOx1HO/QN+80hdgq
diu6HOBMHtspWyDMd5NA7brhhlimmXR/MuLxgw/1jqatilVyxsQxPat7/38GTmn0
nlXTeu+vsG5GZakTM1Rt06OXsp7sOpohca3Ad55VP8N7iWQsWxk1kGeORWDxfrwX
qWkWbpGC4XlmOclPar2KBaaVxa/roYkEM3N8vNYl1M6VXCWSc6AtsbExg8Af5K81
cQKf7XKMkPwE7l16MT1LqrJzsdXtLmEr1Vxit06kbopRHKCc8Tcm3H7YWLhPQlbj
F75DsD5A6dxYCkbs9iOpaCQ3BQZUuX3SeKV5yED5UbWBfbbwd2kV8IXd34GZ2Kd9
JBi37xpMAczGZRToLfpf5i154aox+dzFRvWcPDkvpBKxeYj+lGyTfHLXQ+XCXWFN
b0S2e8TqtIAzzQiRJy9hwOqfbtlY3Si5drRyv1/0+//luazKAi2yPpUu9g91KQOw
w2KKlctpEa0New3VdKNyODdO6hMqbReBDtwgVuT4Pl6vqdUPApmeU2ojAzIZYueh
1dT/wkhn+nbJLQcWl7Fsbk8cGAqKR2g/qH28Kswlad+O8rptsx0xjqN/Wrco/OZQ
xX5/1vL5M6oHfoLv0sbWHh76qQvoer8lspNYXiyVhOMjYZOc5Ti+roVp/IrwNr1H
hH4KLvUxn5ZApJcICsVnSTnR6nmojx6m6laVj2BBIcVGwGSOcEfT+trKj4CegWIj
U5h1XU5NdCRoRfUUHFGnkfVSxGPEG1J03M8Nkz0KkonKwF8OerIcFYZ//9MmdJiG
A25hdVnmV6zsoJq2GGE4QfwCTtZahnkeSNlbh/lWnIgsDWs4Jc/ABpyAAZabXc8+
TRYuj6l4vgQkJsl3+jZDwUUXUDt6Dri59OD8BG+jcX9ncWbxti4HDCs1JD2WoN2T
37oo8CvexFJXisvWjJ30roRYSiWaNFVXFBgZ6BSU+aWtsrOQk3K6GCzX6O4y6kmQ
Ka5ZoPvY/m7ow7OCzM/GqVGQSdEno23TvCo1+tQRzRm73TSRqv2BKKqjpFkZ+XKE
zW4kmNcjgVaqU8jyjsiAz8n4RYPDuyAM/ZO+IH4yYq3S677g0BPzQl5EmXgP8GH1
C1lkdfRtosh6KRwrZ3CFPxSREUDMUDOdpzGRP1sjv2ZsI6Vzy3wKtcZDdTvYNrtg
rkU6eyjHa5cf6iXEgf5GyVs1/NDWdOwlNgMfGPHKffdG1pNPgU+wQWtpaBJWrcvn
Q59Y4Dxqv2mOOdR8dnLcVXEFpI6xBTSApbHBPkQnt7Stb76vOZowdDSrn7j3V58h
xf+ENTQwBQK3UGDvwWm4I2YF7EV7sRwf6ZBvfYIuTQaoaE0a7WzxyB4WGepO9Qcw
EwsduDMa9vLt7yj7shIHlIoDPexIsFnC8wMmbgcPOM3fsYgV9WoLhYWWMcH2uAPK
00fk98X0ykrexW6+hYOpWUbhdE+q5xNIwFE9tvNMx1MZ8n5KW+QYOtjJSze+YktP
GW/VBUwTB0L9ehdkWg8I6yIr7dOGTKzMtgPkMTR/I4obEtwiCCbEfbF1TrsqBg5L
FLjS2XC1lajOFkZP7XEzK0f4kTsnbwADJntB3AkLQXM9CwUCJlczh+OlqdAeYk9M
/cmUQEtqd8Y1XZ+6J7o2hd+i3RGR0mMxlKUgOolyR/GnLDX66er7HlC05aeIr4SX
PkKxBooMMqAA8lu/2hD9PeZ4BbfNKIlQsyrGgnGXiEJQIClp2e1VtLak8lK0T95r
CbDUFhHih3JC1QSNXk5+4zV60XL3Hi+0w73X0Bguz6jnpRyBX0TeShxpzC701M5e
PaeYjJKgp/5ld/8r8v1TTEqld4LwznZQDhv5SJ41dSs+gbzfs1imDniHX9Eg/DMM
XKEs4HKEDyn5Qs96ughPDn5jshbul1D1EQIqilRUJMFQtEfskNG9KqgfbTYhHY2U
BPGQ7Mvual5gP19TMWp8J8UDjJ09GbGErXED6mlbTqwP5JJq5BVu0xK7IVcgmGzq
IGkSUZXrsMkVivSKv23/sacXaZxz29O1J116cMYwUXuvN/trnZ3Mncl46hW7nPNZ
J7HYj6mHV5HRqhPCyw0B6VPoex2xhv3wR+jWbZIDY1/4dymkkWhGYkMykYMbH97v
i0+yfla8mtlT7GsJt64Qxe44DR/M/XzFyPDMYBmah1niudCEkRAHObcO8xKMexxi
KvSzAdYN9N3zYXO9sIVy0l3I3IE8dG3ES5e4Zh6z7l+6cDVD9QUekQl7M1+D2xmB
ooYfspTYPqeHW57qE1tmAFRzoUiADcUWtwmJ2tweN3KX73bbRfLmIXd8JG8b6Xqp
26tEY8C4eoPiqEznLKlCzDFIQ7N6Kk6mI28sJ9DIDYyAPdx3kF5B4SyTyi5ttBOT
nzJ6+781KVEkiKU6vPufO57ppzvFyeuMrlqXjnYiRdrcjPxQEbtcAJKY4HUJ8GEt
9+Dv/YRtwLfxIBedS+zoDt9MjlI0L8zZc98UejZ2K+OjPk4hDfHrNogp7kBCXEj3
VPIF4A9ry7QSQ7nrNcBtAw3LCyLw8hWokh+82CGQEPiY8+BxkL91+K7knqONH3SF
yZJGew/1nv+jFzLbnKR0HIymn8Nc5flAvGWKifOhplfRPvp2LR+td5VRZ/MeYKLA
EUWLdfBDQiYygMb0NajMDaHH3tfum0HDaiha44qEbgdnKpMTtbc1gwWdNl7fm3VX
Rxv2c8tTiLG6QLGhtagj5DzKHDJHHTzpkapiSzGQVDCD94eBdezcwvsYcXl3xcOp
gCdgsFq1tfYR5wyChtjMyVawq+inmDO0CrgJWd8aIP7Yl8ty83TuOYnI9rqcprSK
UgTL9oeA9eh21VBFq2GvPqIY6rSCXHAohEXxhNtDuU/ohApd6lMPWdYhzR51F10c
rZy6WSQD8Od4BxmeDAK8reE8elskihNvicRxlYGdyAlA/mGKVzLndkaFiV54gWPA
s53GnR+9RkPZYrJ2z5G26cVq3siQG6pcd5Jwj3nuToZ3FYXohkDOYowLA0RcD5Sx
AnwoF3G3WLvq12b7KrMPjwZE+Lhr3ajVH406p6yiKzMLt8ij4ikBIZAOs4x5nc3L
iryYcNlnZ/vax8qYgqI31ZP48kRx00nKrsN8fJ3ASKXatvOnPxjixqL4H/iqGQnR
baVPYhp1N2sg6T7XolUzMWd1FCfDPPcl0aIZSEZ8gdcUT02WaoFky5+8OsyWWYZm
9Z4D9tp7+2a+iw82jxr27k2VaLuzLPYsRj6lC7rnfUdshTaT2vDrRNjfAcmbskSd
VtTVsvmOW1Ey1cfMMvF1k1iOw0vTpP2mcrLQDpnloryNguGZSz9BeGbw/Ei/4efK
lAxvuUqnzeOUsCsg6z6D1bUyfA8wRREjTubvA5jM50/zC3/SaT5DGtxWodRXvUpI
X/BL4Bb7schYo25uMrxJJ3wywOc0tdaEFthHNBlEXsHqZI9CKEfVb9+KCttBbXsZ
aw0OB9avSLtp61tq7zUySL+tr4iljnp6xF8pOCUvLWNtBvnEvCL3Vhn2WDk421MY
1+5jBhXmZrACre+xfhUhjRWNOO8Rnqdd0tWh2Hi3mv6LWEXYgImz7LxworVLYfK4
S+0Pukhdk+uOIXbYuzCbQXmQQxAaZLKPZWm7Gz27WwVXzSKZ/nYoNKHzDYdOppSw
lV5yD65T9m/KgNaR+D5Lbrwwd9yVDGX/D0BvR6yUQ5E8S8eJbDknLsC1MvIuASwx
IRsaG+jgMHHSIL3P7MXfuop0o6MaTrrBEEvzHWVzqNg0rZtsnVd6joYSe2KKDqg3
PbjcKxSpIIunIBprEO+Vk8zR2Nvdl0dC7WMuEbCA5G2zqn2AeVhXy62FTpg12QpS
K2hyscr6snsvSWDsw3oteUXi1iWiZZku+4u/R0ofbrLvb6RnomFW3+tRQm6niwgB
jN2SbPf4eydYkWwgcXlww+XRB8F0Oe8rafk7MUojMJaLnHMZbC0rP2n3RZeFm1dR
32tN0b4eZyGLcVKG87s8yBT3FXdB3Y6q2l5Ri6Z1ffiaYS1qTbV96F3DwPJu6pUX
OB5NfTHB8jANACT5Sku2K236dva2/TDjuLhJ/5VX/3DGpJWCpbyTwC+WQ0hvsh5a
4whzddX+jfG0Fvhgg4s6REaWp0rRxUxki5emTCWKQz9RHcL6RyZcbKDK8I3fmP+Y
72vPZB0LJT7WqxjeZ8XfiWkminjjp/QVSOtsIIjasCIgd7YhBGs+5XtZpNXEVlo+
4md1SpUT1kGozEYh70bD+8pot0Eo/e9wQ1czH3KBfCAxfs9dFZYusXfv4pmsbPVr
G1UrG+CAmy2Gtl/0hW8EuwS1Q+dVI7zXb7xnkdcQSrS/xxmn24G565jjMPegyX2Z
QrjfbOiNwDbvhsP6nmhZyvWTnV0VPgTfP5xcFOqxM99wzFnrveU8LbSYQEDSYYZd
3UtE43xDAcDQcaYwLe2AsmjAe96aLdhG/5aeT+xGQ+a4L9PdiA2C3D30MFbuvgqn
AySGDG8G4rrhll4J4TrfbiHUMQLOmyUKu1FYaKwI2Cx5/k3IWV9kRZceooW3nOFq
qiclq6Oi8r6eW7R0GlwGnpDLMbfkwzcc7DxhwEN7oWXo6Y2l0CILO3+y/AvJJtIw
R2ETvWvLPAPDc7jiWrPCrYm492kQcS1tifR43ol+0waVm48svj8KUMLFtxQ8xGLA
PILSspzGCZOmMvPnCvKZKpac4tkLGB4JpUoiLmI0wTjBRV3eBQw7qCOQZLfMx8FZ
O6B4N+ehGX6gZdrlnHtQCPiHM3D5csmNDpAfW0TsSTTeO04YEjHs9vzw+gwQSHrA
zPuhwyFi8o16CfsKiSsEMPaeyOl8/okXJFDjXtk73zvKGEZPISqXBCEG6phCgMg2
jvqimtd49M44VaUb+43eMKLqCTIYtPZlLrhAWL/Mfg/7LrP65IX2AoKxSch2WEGx
RA789wq3ypmyxxXmzREeWsEGihEyCbHPwd2uM/eYSVE1XVpOMI4Q4VURjGDK2fIF
cQU4PnPoHwJpX3l8crBxrM2fHe9+tX8D4gBBu3pQPutzOu/QTLgfIEUgTh1Pw78t
ocCdSOTRSZT6/GXlbcqbFs7BIEn/oAfnDdu2znZN2OR5ZqVSAm0S0knFrVztk5Ey
dSTVRZ6WiPE9d3N8+sXKu663N8Tazp1FsQC2QFg7p7ljtlJHLwkRbO3vvWU9MU4q
uHq3moJumeo4dl6MzG3n2q1LAUI2z7Amb3t3/gmB03t1IWUClX7pXUB4rRI5gDpy
If7twLxBUBSFK5ejr67QW49YFsCgBkl5DjHfMJ4X1Nf4mkCaJ+JAMQz16HyukFzQ
jZ8t5ZN266rfLSZPqkUhTxsJ+gH6gvOZ974f3jsH95GaIab2bvLmc0lnMq3OHxGb
5nt4MogugCYup+qtVBwSt2zXDN6Z8mwBhLlsMj6/e+qTEZ7yBWnuvRZ0DpnhZZa8
TBRX9eI5DpbRb8AqjLLOZvVFlvL9TUbYBGbl4Kynd70iyg+l38Bn04lxK5+H0k3n
YN0M26d7qxE+uT2cbjjSMv8oQGAT8KtjKf89rsBdC0/mo8k7eUOZ6uixBUX0IOMq
tZJWzEMixRoKFii830gKYlRMHeldaSvZtO6s+nue1WudkZKOUCDz5Z5dMn2TBFZa
ybgnGUfqufe0pknxOqgLy6wgjjjCcvSMA5tMQUnQ4/ChN9271D1NjzfIi0OFnDQl
OKf8d1OYgtg1scez7oOxrbex8hJxnfYIjCPBZrGywGK1OZnkNpt/hHjHNnmIF7cl
37AxN6QkCBg0IHRAjPFjy9RRIlBsaVmMhKL/dOux4sq/8UNYJQ4L4Y3pI4gn+WBL
V/Vf3tZRE7Owqyts/d608j1VZPfybqB31tg1Du4kYdxjtoEVbxpI66w3IdziUQLW
hL/hT0+w0ifKiz8f2GJTr1nj6yvqUchFM7EjAcwKdTvYehTOjSkjLw78NHSFHyDz
+z4XAjhA6qQDypD2tRMhpsMRzsqUvxMh1HqbRnfZR7BnsIh+5Qz/dFHOdBRti6xu
zsOpeEhi1JapgrSY57UBjdK2FL4MRnbs77aXeLOAFRqKEEuyoxA8Y/db4IR4rwUO
MSKr+7jJgDMeihzAzOfPFh66thY7YT2pQpunNstz2pKlVc0PAVDfmtYNpY163cCp
FZ2js6nZC0dopqGfZvACh2Y8CtaZfvciuSfSAMMUITCornH5qXgwtCrtJIXBbXhQ
/Vg1X5xjy2C1z9a3X9PsPIljCaKOFSkc2T9otX8c6/tO/JlKhzQcSZKdSqUfSZu8
d9915o8E0HKGUdwXljhux0XrDAX7i29o5RDWTFmm1RXq9aULBnPmowVLSRTcbnox
hSXlHppsNO91e2LGRonZAOxFZ5OmYA0B+XjbwUUsxPJMh31e4VBXG+c841AwRSFQ
mEH5qOE0QPuXelfIf2fCwNrd0CqDNCdKFmomaxsrsOXEAW9L12eaj+pRUt8wwmpv
Cbpr4SfZiEubUgJWIZJmyzzVid0gSGaUqPpcPF3Yz5tXuMJ4nPpg+CA7S+dLfqtZ
2bxmpb0HGV26RoDBOI0c838DHXhT/s64Ns6C5uLTpGnJRgtn51F5ucpSGgPqjoix
JcWU/ogvUcqQJHG6CLRHqpj5IItMu2HtCoPN7oKrKHAGtVYFZ85nEAZssylCc5Lf
MAfiUDrFvnsOBF84zLLHB9m6pW/1MmLQX4pd1G2k12uRbDqcZT4Cq/pj/M1d3yQp
cbk3H9phE7vlj/IqCXTZassf1NFn5iq6wYhj8s22IIAAKRqoKYwTcytOaSjqONFL
iz0uuZCZENptU6j0H8vgZnfmgGNwQyrx0UeACEQ9qxCGsl34+jr6ppIupzcWjseP
+Q8TlqZa1MVx38CjerPgoHUCiFwtQ1ihXql7FoRyj0ozCWqmm5jZeCaxddnnvjhQ
GJGUv4GOPMMA5a0pQ1t5sQDZjWN8CBopjKJy4QOxzzsfsbcy5fciJz52qxE5SOzT
FxkzsVZjJl+tiDWy5UOjkG9OZhILU5k4jlT6kNnkyeAw/7ysmonJkMbHMsCfu3zU
ofWa9nnHWFi4HtggrmTJp60m7y+UPt9KBMTYat/4SSo4d6YSDd/gnmtXPAYQQf2P
xNVVwJFK36A8IyiM68Y11ivhTa5eUc2Y1IJeAbf8ezQ2hBoeayh15xuoJiG4le57
to1LW3yPQ8D75GArem3Ttu7JZMB2ViONw6BNwe7YrxbLS7oW+Bri0ucZRxTdvV+t
ZHc3dD6p25vsvPq+oyhU11vk0qctZ2NdgZMTF5HetBlK4gyQSfnkoIRt7NK/COeO
ZTX5lRD9EZr2zI3jLqQzWybBAQtKFiL0E4JqSMXwLBy1uvB3plUfhk+3Unb9MB/5
YdT07hQOmk1UnYmuD5lz3BiyBQ2CcttLY0Jg2LDr89/rCsKHgm2Abk8y7pgExGrp
PqnuOxIB4JUU+Z7wrdhALTdMvjpgA8UH/NFMRyixH2TgGeSJshF4Mhx53JkwAXR6
u7gARlKCHwcFyrqBV8QNz8GHAG41nfBSar+kSmKXqlWFl49l/cciSgqo+G40VVpd
Enc9WOPwM661RWPJ7ZM9q+ac2LG8Py2aiJASDsos7VinPUoM0YnDsMtyAlcIwPv8
siWwH9nklcQjcPblRHtOSCE7bnLPJ6HVQAu70rqRzmW4crenFUdspQ72WcTubTzy
71+eJlXRDrA2onTkUvRftZHx0y6E+o/NGCzL2JVUA/TEuU+TY3UtAXcgyeSO4WdR
s/C3dA5ttYi4PDX0d+ufJffd9+Q0kA3CawZ0PX/TPFreliPwcg+Fjey4q5Y5y08p
i6V1YlXDR+jisONyk2V2i28F7v0exKyNZe7r1UXc3Bs3QfSO1NHV2Xx3TAF4skg1
78M0fJtCHK45okZb43Qc16MVf6+pIAxj4Td+ZFGqXKlhUpHWzIncsseQSUzAfPbe
tfxUJEG8EHMh8wSUtwwJprQ5KqIjZU2SQvKKoMkKzbLvzlv6RAUC4iRIOnQJpcpi
7om34Ng9uZh7EQwJo2E11CvyUU1OC/6U0dHG/aWX2z92alczy7PcG/r5ImtD/QFl
+oJB+TXZeiT1mQvjPjC127BeK1BscvCw/J+SKirRLLUu/h+PXbrrQ46zz/8lagCu
j98RPxYvjhudSP/007k4JkpKsuT4l8TI1i6EFhwa0m1ZQkgRelss9JdVCLBRMWnD
xtJOLKyjRTgvBuTweXYnFFpv0Wcc4+MfT1cDBHn1PjEVzrVYm3yRPc3E6piLkWQl
gNBXDt2QliiBuI+R7ESykZoVauUGngsS8d6PidwCcR0pdM1hFLymTcsMgr0i0l/+
hWOOs7tP4ND6OdBNH+cvc/hPjaXZO1PvVCUlzTtH5Ywgd6fkXqAEcp3vw2Sa+3Xp
ey0vaxsV8xNwDRomjRWzEYjTPYM1pu1anhYXiY/a/Hk4UjUcOayJAgpKMWR13E0H
SyupLimNZMqEo0e3HLzwf1uu4BYf1hRJG+UB8GA4nw1M7/bKlGE8a1Rnv78T6Uhp
F+Hf4F5Sheo/sDJjG2eORFPHWyMrIfzSvZ6ZoLGvQEraWr71lSUiDd1rcdPK7Uiv
m3hsWsNCVoxrCc2bhKOm6Nktzukh2WSG8hCphuFOz7YNblRV96hGBLiXu2xm3euI
OsMzoQCioyHod477F0a5+fthu13NXQDqa/pjJ3XD3b6wl+QRfXFOEljIWVObZfZH
DchUbvYKPAXF+r72KvFY8m0NsBQhWiNXrI1dOCtP28KnzEvLHgqNMZgcc2qHGqkT
6MC9/TKgJJ2+9qSzfGSGoGZ9bcGHEdhNMExG6+FmFcytdj5RgfJqhmRJOzw2pLgT
0S4zUEgQgpfKPjxNcc6Xaaqqd7dwooLRkXT9m4jbdGyzRk5ohfNeUY4qb36TBQ8u
rd4iHfLA9AjH5oHbHb/MY7YzrVsWusqmOZ5vWti7w/L3WrDcq3sKTAL9ovP3d8Al
gmUhDG+qekWEhNKldYcnaN++22tSbcJkPZFcRjNJWHp9POPfBrtJkkihK1d0RZ2m
6/a8c7Dzo8YiJbbUUfoVvfehkvkLdhiGvf6nQDKxk77pTvWFP2o+Jjg+VseHdmZv
OpU9udrJFV3Z/04R6A2ZQSAl22T5hx2zyE6PWWlN0NR0HPjlJ839XstzzGF2UKx8
3IK5Z6N/THAOkI/S0w6aE5uTI+PW74PLBYExxHrZhcFI/k/YkkI7LKulJFCE+bLJ
Cg4McCF4zXlVlAfMd4tB1FpNo1nBSqD/QPp+yS1NJeTApqzKgfX4CehwYAgypf2J
X81jdxQjkWyvtPyz+3VxhROKlkcWjh9VZ/jeKei6o5Di16gB3BK4K/hSTuchCcxT
lYMNPRCF50na+svsL6QcP8DMuWBtjxP7125oKbEtdK1RFM75p6KO8AjmkGe10a9z
tOILProF1At4WlODRbGfZif6RQLQZcR/dqGnr3zymRWrHXp3CnhM/Hw4uqH48teS
BNBD6kn3/HqxzhIwuMJJaq1qIpMjFbKroJQDHrJ9c7DhhejwJEC2eyLCCDi8qQGz
NicmZfIcyxw4YNMW5yuEtWUESWg/th4kXLhEaojxzyV3P4cjPW/uNZL6dkND8pFv
4mR6GtPY5jMuO2q07xCEDqLduIULbU5yd8te1npMpyD2kOBSl/rb4RictgUm3q/3
Af4VC8IYkKLoHARO/30qLK3d3cqLsLLsZ+QPLH9W6muAGIGNwSCQkhypbOeskYSo
mbejRffw2W/N9IXWc/I7o2pQHuChoxs7KBUsNe7/SjP3QuQv1s7yAoxQf8dLpNyQ
/4hqBiSb44cjDbzUlpvM6jvzM4u21v7YtLi9+tVwKBQBDGYaXTS9x+2w5LRcZbvy
cnQR3JUq/Tqz1SuysYVLgy5BtiCeJi2PEymlekTMG95AVT7rOc6GKzYfRiBDkbhR
NctlqpCFCXFlFA0sA63CoQrKKlVnVf+xMW7RIaYCxSa9fEEmNWDNnU/Z3wH1HIul
408NITEuBAjd3s3UshjbiCBZ71gaGgfz92TtRO95/Me2qbX4gbdj2LjhxHnKkR16
5hd0KL5DVpRda2JI2xKXhiPSGa/fs/rVulR5Fk+5ln1ucirYWP4xn4y9uCZkUlof
DAq+jlcFG5rqpOdPczaZm7DzrYyu1EHVk7dYNuKQlpMQxgH7qTv3qHSG4X9oQQRO
URoEdPqehVR7Di31ADemciHpZ76GmonCaGFTJLMEtX2lIWFUXg3ltm2ofLkmxS6W
y2mcbXcqbviw4ZUafSCUQz376zTEr/lA8V+0JVr7p8XwQKhV29blD61P6qbyjJTk
5dyo1vvGHZIg1YFjzZ9FuDqnj+6qSfYSLgtPnCc0N2HJxUsMq53p5z7JptLvn08b
6tnxIeCGUkFVmThHGeVjVtyE9EvZBod8Uw1OKukG/9gdMEl4ul9r42qG9AAJrYPR
y3vHn8HenzL/cM6behuJk1ww5czI+uyfawuskEaKeggGYL6R2451NHMnlQQb87ul
eardUzZnHyTpd9Bx6QpDviTRMzVp5n9F6LiSySdmhQk3N0gFS47VZ+qYXnQd9prU
aMvKr1MySzIC4klOw3k+V3xftWfBThZapa2ilKp9rw49lrSHGseIqZ79hksxiEOs
sbAEtR9RDWcRbI4Iqxbl7Datg4TbVgkdlJbmjXmddmOxGmLd/m7rzOvKUZD7IiVI
obk9gruO/TpDSYP5oVFYXlwCN1dV17ysNM/EyRh6JU2Gy6DDs+ezsp+Eim1huBvt
NBqZMj5hBxrr+GzRZiIQ6UqJPqIJayQa6McvwpJ7mLGRWCv3OI6fBfzwdfgQdFvn
lCz2s1p5vGvC7yqjVIy+foixNEYAWwbm+/t/AH3QqnPRd5LhHor1eZNFqKfSSVJz
iI+L7MpKTB9PKA+tvitjPP7YsKRyFd59+pjHbtJpDiDH5hze9M54I38FHGBdrbRQ
T/jFtkMn8IHFwdrgx9pY6eKz0FCggYDF/05NavL17irH2/EShI5qV3/bs8lbnhfj
zwmErcSws2rpWF1CttIUAgnYeLtyijyowBiKp0UV3qJbG90x4Q/DiHZdxdnAxygs
wvNz1QHpqFTUaCLULZ1x3kUOPlxv7b3eQWiiq5NoqEHiE3itKm9JFEB2maMLPYRe
aug1Rcbp51jYKvsg1coGHA==
`pragma protect end_protected
