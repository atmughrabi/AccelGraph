// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DuA20BoFqZ9b+RHQLCCq+79NkIKxTy47L8wgwJ/iw/7ulRElYRmL3+GXeWlDWQ2I
rlwdHXQCi+8qLy4h+4WImJmbP3FgzbL/YsI1+X5VSkbuVWbY3xybYu68MWfcKVzk
3BE7PK/BEghlnHn+8OYFhZF9J4NskOXfjy9iVHmldLc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3104)
n9M/QLONeZeGbdvDuREKc7N5R0PB/lNrqiELDqxh9a7vhZQCb/SuNUdpQDuZKkdx
CXLCyj8X/dS3qDGmEEXdFU82xPQOpVvbBi9g1mgnyfqdFTlvI8f5KFIEnho9Y24+
E3DkmbXiOY3YPCJctaNQ4r97Gz5kOnz6efcacbekcmVqjqHiibq2NBomNzwHcREq
zXvdk+CXsShjCCaBLSmI6731tv83mY/Pde2Za2XpokLkMvtyUBMO2J38gKnQwcZL
/yqQkgUPf5vGDINLuOtlO5aFuE19uMgh6MsSgKJS+5iQ+WThX0iSQ557ESI1KeI2
uS83Xx/c4Hdvq/KKyTLw/GblEDF8Q9dNx+7eCXRky35jBz8L+RnRFiFpd7qGgBUw
J4yXSMkNpUcI795z7rNIJNH8CU1fRx1NUBBHmnv0MMRHFNKIWqhkC6S/L3uwpIll
tit+XMDRJtBlgqxuyeICAykN/JYjt9vbZ9gDdsgdndLp+IAqXxUHXWKRcS1R56xN
LNMviTugq2mmwVK2iqBHg3pyPPB90CTkgt1Ykp4kPpKZeZMr2RB0mZaUp2ugknyI
UHM9PTTWnyzHY+C37da5/b6K+prbDLuKAhiQmbBmsIv+a6Sfswq6AOfAOQTwBCtN
p0CkytFjBnkj2whX16DCqM/OIYsAaMpttd8Yc3oXRqP3WF/h+8S+b23JCQKzdubD
HVIAWF2VMybCOlhU+ZVB+lIW6GkrqO2I8Wu7wEw+EBS5IhWuH8zVo/TYlzajnOCM
M4N0wN5sT88pRFdm7ZnRkJXHHngelFJiAWAwwOPASosK6DpYpK35Y6gLjo8yX+wD
13/YBy8fvTHnm6ucoVjN7+AJy/ORThCjpdMRu8ZCRd5uZBcJap0OKWI41UdYAlfo
mbWpOb0w1NVV7aoGAV2b+15ekBD5ZBb2rGcG3aTmoF4LQe9yZqqR0YT84v28CWuK
t2I2kKbOw4GuTP58dfuXIYCfnqWg/WkQJ1IZh1CNLH9/XuFpBgrJneYZSRUh6Ud+
wOJEhzNDUrPye8bFY937N4mTcBUD+/IAO3abRVPTQIVSUbU4bJWTmsPx+z5qkzyd
jXNdadqyWY/8LaIEJzokqPvvlLgaNpcaJmOGpkJz6R9J7VwS6WhkN1jcc2VwgLSf
2MUE825TyiMzBhxemQIMUfKL4HDqaQNPFiec2SKkFk3sBwIkd3iKmd9Ip6tB9sPy
vhLUvCwpLBdwQSqnC9O/+NTL+d5wZpz1Z8jpZpc8BMWSiFKGtK7Hnp2qZR6/PFrR
1GGPrvQ2PYXND2ft9GWpuPAZEx696NrQHOlsDPiTyDeGwtqh7NYcmkr+QI2ujftU
OvPNpzUHH3nyoR+MooKAQXPhwoTSWUAVMTsU+JRuCChB8yoNS3SNUGx3OQE4qZpg
lQCuy6jYCcPMW+Ap0Z81JmukjLLtck63p9HB22WHu9SEwIk6CodzF4ZjvCzgws7H
D1Lmiu5w0Zs/bX+wFW46m+pk3ZFVgw4rxJ9TBBOh2MUWfQuEqlg2dbS0DSzQNtXk
UxsHliddh2uy0WelkRCTMIMUeC/oG0sukyqvmeRU5sm5qe66e30VhujUtUe85EBJ
dWbqUGtm2HpRfEzLfmKfmdnHE9iaSe0VNQuoVQXfosBHwLG3/B+079kxW/gYODk9
5j1v0/yZnagGVtgK/uJBjqXgZ+91KC/IjYRGQmSE7IVZPgWF4Xra+xLCpSpFtaN1
z8GWgclVb13U5ksOCHXd7naUzoS4+mrrn5rNwca5gLFn0avQhWoMLqgyZL0ISPsV
FmhsWym1IBmDh273BtkWsvCSZvncKKZR23t/r5JYM2qfJkXBayk7Lgvw8VeOuMZE
gLnaIOeh7m8eBTqQ+R1KvxE9pxwmTEU1VJaYnCN6jC4gk49dfsQoBNXvQXivba6C
CCmqVXOgrRhnJGSJyvviAgugC3tI4ZHHYajrHILVcLYr9cwesRG2tlGMS4M0OkfK
qX58X2ixjbuolpKIp+kTFRMy5khKezLZY3BlQLJ42/gi57PxLWmIFB/xqOfvaV7R
fgLAsaulMH4MeHvdnghMRlqG2nkpQnC5mz4UtfpdYo/mCGRqfN3BwQuASOMyWttn
Ic40wSC8o5aWmgmKPD8dbGRBU20aBF46Aw9e3i20w3xuuYH0UZrZkqOH4cSx1EUz
tBT7n+XV64Uyzrf9C+ClQ8UgKGDet9qEy3gli1LaD7OnK/fi8ZE+yRWBNjuYROAW
+orPt1YuLXHw62j9IIczCf0Pgs4zoLhfOGUBz1xfyyoEktuMt5oj5MyO6TnMtKGa
4FECJ8W+CShxsP23juWX5MF1RFe7xw1ugxXKtqTCHTImiD+x3qG2n4YDv8PDGJJr
HnwcgNBrJRmzx3qLN6DOgNfPJTIhwGmRaMx9ozXvw1EcA07uF/uk9+nsF6xkStVl
WAqkDjucZsZx/S2uiPD+XQm3KpqQ4OehXKBT4XPVuSGrHJ8MZs0pKw8IL+tVmWFt
ooF577m/kddzQvrGHHpRdYmEmay8PENroGI+/rL5flLpEW8Bb+bzbw8JNDIXqa71
yVekU3a279mCHoRMeMZoo7xnR7ll4Fo3jf8UsiiTmNRWdrF2xWyaweXecq8/vdPB
gKobmSUkB1Fa34B+Uo+c8cJ1bEvNXlJI+xmRTUW62j5iEHyTMgHVmo2cNU7uIx+m
NwNPwVNDsDiFi4cn2RB9YC6XPnMCqf7IL9+WglLk/whCW/2HrlsivNcSyyw6fW6U
dB5xGCVXQqrI0Lehi4EVfMJ8GAMRwXAXfndsnSjL99JT7a3y5cHQNmnezDX2R27A
UmJGR07COBEBpGJw2rtvXrsen2FlMUf+ipjFK3YNdUkXvrb8hmdcLpEtXuOBOVTx
WLdXyZkC+klJOrGmTudQKgFen+u7k4tfTXyVF2c2ElIp/TmLbQ3esw8Yf8t7znJA
ESIAYJBzu532qLEMfxj7DFwdU1DQUyjFQWJiY1ABAakBNkL65Eu0XOSxmGiZUJZ5
cgZcGb/fNnM4uip1yKHSyzB09OIsQBtyGnOvoAN/vSc2A3FU8dNMZgHDJD2Dh5Mw
FZbaXA1kr2iSAwfe05roDpP4VnyR5Ni9VH0nkPohvmuw8bDlUm3Qa8oYpL8EO+hG
hdkGsj1+20NtwE6OHn4NmmAYXqwSE2jcGW9oEUrksrCrZY0Wkw1J6xO9fWF5U3TF
Np7foWmKMS8Lz63+fOd+PJyNzdhCGfdXePLFPw9azzM0CA1bwyub9+M/RnGiKf1R
ek96HDuu1Yzd6FhYZRc0dPJSDGINAmZS0zOijGb7NsqzrVsPawmK3OnvC5Gp1i3E
dKBIpuRGKwV6VWZyWL+Vl3QYrP4hVYkVgZfcxFl7JWx2/2YE9wcpJY9ciU850iUF
Q92rSIBPq5KUh/JwCKyYnAHHrXeVzp813+0RceGNCS6Oc6FHYiDa3aihAB/VlZpa
jM6VlcxycRiVNs5z8iNNyPquIDamxtLuIjJxP20Wmana9UBnXoLkCk2Vmr7SWad/
IsWiRz9dWBnDssZYTWO2bS0tZKvPwwv18tfJfxEnoBnbDXvoaI+T9hP14rMxTuNx
UVtzhkYOGPZfNjU8Si3KxKeD/+UQYcB+FVoK9lbrq3JCHaCBdN+N/EAbfdQ4Som9
949ZusGy7s5qJ9RW+LoT3yeaAsE2mISDdeSkt41P16R5CTYflT8IivjiophQM92i
qThZycQOsGBAccAUhRsapJt1+sYK6cXGT6LMnRWPO8jAVNT/E8xBMpgFLFlBWbqk
NbjcQVlqGS5dT/i18gsksWG70erCTN/bYA7eaJfhW9SA19iSArR5RcdhP44FPBCk
WUnaULhhY6MdRO/poFsADvrkX9E8o/W8xU3+GC1MfnvqR5vMoVl6yHZSAPQ1Fmzj
d9eMfJ7Vj2NIOzBjywRVZRi6JzV7G9rXHtRmoadQoijfJBJKPH1f0xmqTw+GMgEl
XP0wnBlro5xsFZFBIB0/smTn5PXmPYlFG7BwVgseyIKEPsJ3RgqIY3gMCh3ub9FD
fSSMXmcMmRfcPkIhXvu2PMxuUu9FzqkV5kI9WYW6blEhwcTSag0VfAr2ipCv5HA0
8yRbYRctiUCpdB/chDmNQssEs0KagJMDh5NoLgKe8ok=
`pragma protect end_protected
