psl_vgpo_inst : psl_vgpo PORT MAP (
		datain	 => datain_sig,
		oe	 => oe_sig,
		dataout	 => dataout_sig
	);
