// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
T9u2RLp07IOFh2MmVKEAx9BOaohNlCBPdzBDV3Ey/ipDGMpzFwp6vSi2fRn9YkZO
/76Rb8QdduRtrLiNQvYcVUkQhno3GkxzgJRtBwoQwA46rS4/rtsCm7wgJNdNQrix
PMloalMdrLMh2LaPT2sXN4uwwgyC0egeXJfquk1J4S4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13104)
7iD3IVNgOzr/kM5Z4vDI7b8ANHSy5is2Bbq7G5BxMG9khIazWVI/BuCn62hDG5G6
HwtUkdwqsBAbIfDCFtZwO4/bJR5DcJGhl8+4iR/vKTlazMXA6FIofI3T1yzzdCyM
nCygCrAQqkm5O7jFOMGh1XsGcW3+PEEJ6xT00grS4hWu1tr+fmaJE9nebjxOMT/B
F4MwBfSmMp3yQgtW7VT2qk571dT0+iEtjfDDKA697MspelSkv2TBYZ9giT2O4/0L
iPDJOMeSeBop4R5+YoBoaivAbdq6G9E0nHsLTTtOXWHkR4MB/TWe1Sn7WJgw8upk
GMIpL4lNuWClvZFt1JB9drRrb38Ty3NTEzGynbsnle2i1rjtEtlO8nMUco5eYrCE
0FcAMQqnzwVh/zZQ1/aA3tIB7e4EjsxtBrtvBkF1HAwrrws2Td0EVLBQh0SXWN9V
vy5myKSUKe+glGjkKfZ2lqJ4TS3zKQY4wU6hcJ0UTCRAiy2XAR8PySxJBCEdsr1o
aT9ZPMLjKxk9ZkwrREWVqibgE/LU8d3I1IymZcMtEaL0bzFQZa7GGmt6DiHxm0Ai
mzMbt53prQFrnyyjRkmuQJbqBm1OgYCC88232WlonGPVHurVWfT7GQlhA8qFohFJ
KLuqsHneKMizEboS1iF3S2QFXdkVB9U94YN61wMcWog2Y6G/i5g2U9ToDkXzJA8p
RKFs7qB1BzLSs6Jt6HSRogZzRruEJHzhwf5vkYcynG8DiE9EmfamXQMaNAk+/MIZ
Hn8ACAIk59tCPm4eTgh2CkmwT3lYxx+bZOfj7+N5r69NhR9/G3mEkD4B6LY7tl/s
MXCC99S6TOtfz5yerHHQMATa2ob5VedhmR12XTTzXXv7oFONFprs/ccPz8tG1jMK
yQ3CJidDtEgkPP31iAchqa86QkyZQ1hxE3Vfa1tuGwW/q+oXszpdKlwtVXYKF8qx
AV63kkK0OolA6NIySFbxVUHD5yv7umvq7v4C/dJ44iyXkGx0/k3IJ3KhMOGmtEQs
7TU8vhskTwR9ms6B786XVUUlyKvDGdQTgY3RuBJg+5UQ6WAwl/fFaOqdCJ348KJQ
kqIApO91UUe9HY8AsWamop/iSg/NKduH10molLd4V0jdt9o+wNy9XDR+GybN4TFY
Z9efj1kPrY4USzLG1S5GGowrdlhrXSytyAX3bFQslyVoPvWsk/86jFuxHjGz3uzl
yaj8VxjVSmX7j9Rm2eSaQQSNayHvz8UzNp14XJoKvWx56UOonSqquAa66p8/1exy
h+aBbk/9Bz1Nrgy583zHMp09SopfFAUpTlCCTrNvXXJmUj3L6l0ZyYyB0Y+WS06g
A10NFypk70RQeDKCteq4xyRm2dTCbBzUWhOtmz0HFJsCjmEqNCXybhhNTxvZJUpk
o5++9YoimlRxl8ktKpMBEgnsDASkbfdPb6tCEoIbTIgDtAzSnkby64Q5Ay5fFjWS
7lhl4AcMKS6bAaACXftqxdIQRTqAV85DOKSm4nT2LZjjltKhBvgw+S6va9Vp61Yw
00zlTAY8mEZEo7SPvNB88fUK9rIrONXMbnVVcncmt0tB2reGhKCvp2FJazXQ9Adf
qXj4qUkSjjZN2kf/ZNqFFLIA/XomySE6p+Hm/lMp3Q6btP+Lc934WolF3dTFhMed
jg9QcrirjWFW1KYKYeXXX9vJvqpwPSdQTJEfNay/xQOWDimm3T0ZGNkbowSJ+OBM
3fl4ARUQu45YnpymD39kT2KWrRNy6z4ohKgfnfDKiiHAz7znD4sf4Zx6K817+AaQ
6AKN7iFwW4JTzfQ0ledoUaKGqlMrnL7O+nPPYjJ35aYWuLGvS467krTslh+3muvA
Hz1scJRWKUNKW91o41vOZ3LyGb5u4JU/7+kBWzmYCp1wlYwRsl+h2KptYRZ5XUGJ
t8nOd89Kyjc2H81BK9eYco+KA3f2l6uCfIaZtRJg2hkLa4R/THKZr3hmRkfoz56C
gG1onpGq0guqmQw+hnXNC6WlhBjhtlbehDueRdflkXZU73MTGmF0XVHYx+/QhSel
IQR8yherYiNEu7zRDyxS1uzPAAueosJl+jS3UV1IUeSDsQwSndViKF7hantN4ke8
sFeaSAPhE8XAcnF4KldDIWdxertPBlSlUuXq9rnuKVh8u25UiEfPKVeaOZvxcZZx
W6uqYdIusM7d1MdtwZuo/RcWKzjFFUFPxkv2Q3uFoous/u7LuS7Y9HQjJp8BGKXE
1PspCnToI6/3/YV/fwY11ZcZdMYvzj1fEL09BHybLvRaQ+JHGjjprBTouFvF5K5V
CBK4624nZlDOp3vKZAOC8E4iJMUj5/K2ekHtATTOz1xoniu3Ycp6Z9RZ6yog5Ivf
boJPe0w+l55ExE6C5NeHeTjTDi75UK+jbQsDjSzp4I5RsfvSqUzCGDQ7sY1mP4m1
vlA+yQ/bdxjg4dbzhdKet0Lr5B0VQXC60sWT4+MXLt8NF36vVOsW1ecUSzpKO1jq
hmccNwS2mknBRDYaiKh/FvxLURgJ+G7HtHIJAyGeDo/fFMmP4EYwb/wsIx19r7e1
kS09cYy6auqIoWbUojP+jM8DEmIfUMHloNLxYJcAgrQQp/0fZon+cJM94MpGgc4e
Uwa9NiJIyK6hT4hy45l6gti7BGuDqp8jpv6ar0oIhBJ4TVMe7MXTqJSqrYfEhsaA
jYOt/BQg9tnH1MzlLysQJVcyvsbgYX3rsK0twizZzrRv3ebaaiPq7ShGoSGvoOeS
/2787EemOkyWu/razGZUc9PQoPY+CShsgRhRJA/TOt/Uu27b/g/wZw3MIh3bCILp
lG8ej+aCKNZIl6YNk9+pDKl6TZOxdNujB/r1sdC77/6pQNWR2r55UZxukyoQwGTR
k5tvWSR74oXVw5AON9itNdRa8DvaUVAJta9pdxrLyfWSWTIUXXLWv6eCFdVlA/IK
BgJjMzOECzgFlid8Cakk7S6vztt23XylR21015Kr1uStOASOyuAH3TDz6duZhPBt
PI5Z6kvFCIjY9kKV7EzunToPU5OzvyBFa/a0wqHz2jBYHATkQspCVnrb1yocse8n
Mn/AXjn+whxSDxNGvKFc/2vUV1UImEx/R+pB6H+HPXYSAwh/sUDhRgB31JKXfdnT
emizuXY0veaSK8TrZL7aPLMvZhGvmGOv8xQs27XfmMtOQN54viCsuOYDSjFWU8ro
Ix7fLYpXxRBauS90o4TYGS5O5HOBVwY/e9cWtTIYhBFju8oVqqWy45BxUWszF/+U
nip5Re+l0rVLW55FM+2NvcibhAckIs0OUIOIXnR46n8LbVvAPAvVHpNxdOmt1dKQ
YM3L9bM4tLpeqK4MqVar4QtmE0T9oW4Da5sR8b2IW3s57ffBDyBUHn0Equ4sNCif
b3Mk2D4R8nVuQFcW1C3gUfQAzMpLU5CUdH0V0rBIIDFrmuLl1x2xWhySoxTRCKSK
NJqB3Y+2puX/xPNwhbYuIgsf1FZBDr8Po+Jfu41a2b1vv7qQ4IJxRoVoUWfUl4Lr
a0Zkdoob5VCBAUOG0fpyMJ4fAJcwhtXr7Jq0fNPMgPRp0kNmAz6Jp+ItwME3UhA6
ZxZqVBRgz7G7a8XyXSe1JEhnH69EkVfPLU3FMEtYeMDTJp1A2BADn5qQLZR6xcA4
7QTAwygna0RAvvlAHgXzB7SjVdaE1DbM7WDDQijA+G2j0jqUUlvCHHCSieSL5iWi
vCLbix1EdnbVXFATCaeiH66ZbZSjz5ZZ+SzCZxTVBiAv7zu2X89fUOGi64GY1G/b
qQ9yZkvJQqcWqFvzvJTxEhFpmgHg99vI4DdERXkVX/Xp8JOuOdteLMyYUebchB1t
cqyZvRaKxi8rjnyC6zVfxMfXsEv3bGvx9SDJEH3MGBvTx3h6AMI5vsfddCzwBFpL
wzsESHHVwzsKw8GSOTUV2kAhNqsj3h7lk+7oS7BrWE2Qjyt2cdna8qddRVTqwyLj
PNAI5q4mZ15vjbGKjDkSEuYuvFgc19dwd+juZQHsYqN3cexwevDgl+SdQPrTWV+T
UEsI9d593Qx73zMmTOrcY7k9mIswqESmFP582SGty5LTrHjur/W4uVeeYXsCUDhe
cqzmq09eI2RDbnRgJJ3fQVtlQ28Utvgla9aQFhHHXHlnOXx9QC28ZDTDriZQpIK1
xUSPHkUUnRPXedZL+N0VDNHC2PjGutAEvtVA+7BhpNdNqgE5wjWlYjdk10qCvPR9
R0xf8hCkPiRvfBCBe74CWP30+bSDcsPGOnfYIKxoKOcAcOqw6zIo6WFA8Z2KrvpF
Ucx6rSUpSIvQyhKSRprh5ZYR8eDVx61oGcyniuTQvqK3cUt4KGJkpvxXC+OQzb4q
CmtHd5POrvQQ6UJLfPC9e5R8SCY3lrSOcV1Vco9QoZen245fRiW1K+NJXmfFLXXF
84dFwWzhM8qWs60XKFvpLopW0VT/aDWnhDYCgTX3GZ0YLYmlxjWyYU/3fuMenSy6
R2im1Cr689VsaF7c45AI/pxWCvcsbOwakHIk+RV1yRw0Zk2v4bZR9IsSHwehyl6l
99fveMdPu5+XOYDkqvMQMK+H2TguSskIqQAAHs4yvtFZd8xXjFhoX+/E62QVIidt
jdOY8pOVVc/9gGPT2s3DHlgGByFexjKgWupWFy96oCTXkvEyKxMA9QaNH8V0f2og
ZTuRGzjtKt3rIgBhYWToslU6MgQwmZ/CqLtXEUEcwPfvBeuYL/YI1DtS8A+VrJ34
ZJ+aYyW+jpZz0pQimBTympGE1SRPSVC9Fpcs+8jrscYvEYY9N5O1qeBnVmxuoBiU
w1/1h1uMgG1OOrU9Ekpa7qFFfXs+gD6uz79/DfwfIXIt9VLRtUOr+nn6OWpy31Fu
4+pA8Fs6eyMEgk1g1Gq5wNzotZJkUNXLi+/UpMxpPl/94/Vstaebmtykd+ilzGs+
Bts+CrOiQkHgbE4SsvP7W9y7na0B0USeqgW5h7Td6nQ4otHuNzT8jBWemLjhQGCe
cArrbZUc+WAuHcyX+6jZUaLv3eIho+zQ3DV6DeDzoX39/a2meb+9soJPH/yvpb9a
3uLDEmG+37qiuioeJLbTUdK75BOo6JvOiGVFe45fqirbGZgVpttlSgDCmEESMXk4
ArpdyBsTjC5wdQmNWzVtR/t4QQotZSXt/b3OHXTKN9/siL3TgXsxCd3e36WpKgfw
lOgXkxkAMwa9ChwaOvnLoQua46DVJbDazEcm7MN1RfIiCUS0Eyi3iY4Sk/N3oI7R
/ydCXTe8O0TD0meXd0ZjbrP1/X6bkzwbr8r0QGKqCDSOHHSYYAfagls48GEJywis
MGqEwC9v3CiMYRL5dN61C6e+LQ4CK0IAgA2lwDoehBAp/fEcgQTBWlliRs1HovbP
9oV4rX3Mu9Lm17mIoHX0cDXJoGJH/zgsP/6x3yU9k2/dMGEkL2nVplo1myO42SvS
pfLy8CVDlV1RkTxrXt5vRYu05qRyD70EKsU1KTXUwjr1Fed0ENk1NVayf+fxDn/X
Oy70sG0iUovjylqDzsjbRQhNDYRtPfaxP5Si2s7vcLqD21ntNNf14DNxaTj8XgfV
wt8rTgLV8tFts0gZUMQuDJPhZaF1sosYqACsecpPzsMQ/djs79XNXA7B6QLBCz2I
cTWjntIh/9KRavJomQjbcFV/YhwgO/WBFEYAGwgTv3U8Ex53soG4HhN2NvrG0X/n
kHIxNzmxIXekxdWdWWAd6jA5YUgc6vFgQ+cDde5woMj5YZQERHjLlb+2MCNDuFpW
z4atiqNEBnitTjg58QGC1Dm2Vips16D4Rz9315YbdgK5ZLPix2JTpCDl45IRmFlv
YhtU/X/5XHCDj9vZS60raXsVvBYIDqZ2nh1F1TLf9Y+8A5rKjaPJJFcpX4vBeoEw
YraZrhs05G4PFvz5c8S8i8I4mpb7TGyNepz93fFkH3g2y0Na8o7/No+kfvnnmxBQ
haJNr+oJwAEBIn1FPTGgQu8aoxaelrw6dBfn2Fpquxl23Q8ooHvtHzC2eSeLPwsU
wfgk0HPMB6v4EqVcD4Gz5BTLBdSh8kidCrc82LPiu5e/lvc1KSn3Q17zz+vEREzS
J7BN0yjAmQdkzi8woBrEjUuzROt02Qsgkh4+jJeVmXBMPUwO+0wFVC35md+0Pk/F
41N7y2LmaQWHAPfTp8AChdgR/AjIu1FTGYfceUUDCSRz3bB8NmyZXCc5QtLYwOKB
uZ9Sa3L+3nG9S8F4eByTcfJvh7UVJQV0SwEWhK/iwYFI/dvSzKVq7TzCWVXj6Z+A
KuLMTs5bJdJHUabnlSwK488YxtiGcxfl7xZUHt8NRfRCe9T1dCzi+UrGoSvqhJIT
zLAzBXmkUo0QmI9WdPcYtp8tK/5sVJ3qFn9NFx/2VEjwpU6V+1lTzZChWfgdwRJa
01zSdoZqkcKdcBAj123J2nza6ozRHbdw4XeTHPMgTlEVTK3B2CChOyjb9KOuATLL
8Wk6OnP990QaF0j6u6WSHfW0K0J5tU782AULbvHW/o229DJNCVte2jhp9PE/MHH2
XgiqYqHkZDniIeCUwN/TR3tMcSftoCWMMZc+Zv5ATAkRA1N+oyD9jWQ1rYKc3OKw
xWtMGUYcvmQXS0LHjFdeXkV34rGRFpyh/5odLg4uxmVdsstIUBvb7XGt+Yf/QK0c
VcH+t6TNPU4nXH0dQ87YRt5rT7mDn1FogjJ+LtNO9choJ1XpAWErzWR8H9Q9jF9C
qp4m0zDq0BNDutmg7Btpmt85C7AtdMQknZcSseMWHGGiGj+FgHYMqCoI6vo9y0UD
0va1G3uiQ42NM9dSIaPmHfyYVUy6RgbPCLUx7x8rAgc1zN1SJebSoaTzJhVIcHPg
8YDikAd4NskldcL+RwCyLLK5px/4VNNOxEkrtKb1B94X4Fz6/B041JNzY/oqxabk
zx1YOdJy/066fegd2nxnJQmYeexv30bROagH00lRuub+mCtkGeaDDT9QHNd81JA4
POpiM9mB2KawwbAraFERnPG/J0BaZACpMKnPCU7RjVRmuXZa1vprRSv1xMd95NLN
A349sEng1Dmb0oMnXDcv3MDCtX7mxGBq6DiLC2yADjcSS5xawDQB/J91c+finueR
rYu8NFCXV6VDzFOMxsHXbcwgvoRJ95d5VpNpsVFHB9j/3yd0weCA7NaN/gCmzCJK
/IOtGBekN6DEoU39r5DzgxD7XP5Lg6OX8BTclZslVcnpTFfxulSTFUyza4LWDXBt
lpnYbfxsYjTZVXS6oPU2hmXOCeOknDckZHpFg6FJzpl9vzoATj0D0aw/4qcB7Xgr
a2pfH1r6ne1qKUGf2tUmTD9MC7GSM5Orn8952kIUnHU0mzqQh0tdisBHsmk7cQNH
hWYUMxiI3YOckkKJRwV9rB1+h0XhYABm5vkydneMcvOxbRjiejEqTlJNTKlgLgVo
hSgZR6EVFsaphdC4zIiJmc/3YUYEZ9CQpjuHu00qzOluvEdobOADGM1b+gH1iL0Y
f7nW2A8+XQzwaUmvObNRHWa0vUkAJRkdizLT1aoDm1C9sZbkpfQqI8Klhd4Fpkbd
u/2lg6QAlTdByxyMdYXLc4G3WnY1n+ILqHipL+DsuXxpVdWo82ZqE4wlCRGsyN56
eTUWsgB/csCPog9WU7iicFJ3GOig2i4yfjSDG6V6ArK5JxueruziGm4vzJwKP2CG
HLpAb4GhGGpnOHVQyITbdQqAvV2vUeQ8dhNBpRZBaqJzMouxNEBZDRusOCGoF1QV
0U0KzCuAIU/8jgDKI8Ri8dv+hVIghh+ss2ApFfJ6zE39EnqBXUhHhgqTf970TZKv
8W0eOaR7zAwVdfMdEm776+Ty7pCEsmMYSYqTph8zogA2IWj00nDUJBXg1madyVAj
1tCOIXlee2beQt0TYxqM4ezMItP+abExLWyHNxv8rTBhNy67V9CW1Gtz3lM1zS1t
NGCNDmE0pJDnPt27b5tp2O+P8pjLifiQlgUfTZltuqFgQRuk2oZSiLXNbA2DXQM8
kVwlAHsHMnn43etJj+uKoKxVzH1kUI9EwHN2861yclTQBR612VvQw+/YcyuKo4xm
8xJNASfm41yqbqtEOYH+LimOzIY5Is7pMPf1PLuSC0hXH5oM84JmUzj1Srlwwz7h
H8INUi//rWQPxfg81QVBVbcN7kMHIfowdCrkKzNkc1ZVyaxUH002ptPosUOEbEjR
4ihFcWXd3hndKfiw9VIFHLxYGf6Zjzv5V2carrcCVHfo9n7955/pMErbi+J7A/hR
XJ8+POxYfsXN/tyzK9ReZL1Y7i4EdwBHLJd61Od76th1e7Pfy6oyEdeAI+CZN8+X
TzyqslLDZ21Jd45oSt870EfuENQY7zEh4CfnnCvqsrAyLopwx28GLCAu8cEDW1ol
U5pS2W06/idkFDhuW56lApOMYCRRrNDhMv6wHz9uMO/GLl5voTisQ3BCYDeNXw6C
KPjsktRsrlqCfiTyueFfhVcKSXOADFw97ddqvxGXF56itE9WXK9woE+kul2xI3DQ
0OEcFAe72epU4ZgCMsnCh/U1VdCOhJbumJUCBUWN2G3yvTmAohlenoKgaQipZaJs
K5QDtjqgSD+gBUFGoP6pTmuTaorkhDlgAIDdZEB9X36dHHRLArnTojb93DucnIJe
No7d8RyA43XqU8XmWwhAJqO2+28vRthQt9ItLj2kWhefgxxD239IERkmp8wAruCH
r7K75Wogu4KlVYFaXMdp7MRlR1bLyiot7UJUdeq7vN6zb8h8BsVa13+9smo97Vw6
LQ4EtWWw3qszrwN5O7hKHEAA7LyiyfjuLamts5j2RiYiwDiE7WNoIfztsx2H9Sby
B+Me8RntgxgBH/CkAcI0/dFrqu1Sq+F/kOCgvvFvmz+fbKbFHoH6GBviLh/xMS01
CO+5osC1InPeHIpbgI8ZjdIkLg9/3NhmtLhXKhsT60EmjW2AKZiqRa1uQPt1OxoI
wIJRZQPbq6DoItwEEhNvmoY8JBIUrMnnhfCF4vcOB3uzPbBp/39lZ8mgK4dfCzik
xS68+MXSL4+Xrh5oWBePgIXlCBRkKAa5/wgNkEMYlf+zoNiZEk2YK6iOdeA7Nm/Q
u0nOfqDUOeIutkM4lN3tOxK4UTQLi/3xNCPZBgTZ6GZYRALLebs1HOQnlFe9YAQP
5SCFZb1AxW2hPahRVJSnuS1ZrQD16bmykL6rf8KmmfigZ/GTnkdxNCMxlzW9NNwr
FA2b515r+m5NUUXm/AcR4qlzbGW9+9vOckhRVJO1SgPs6cQt7701mVccWjRrht5E
5yzbJogeXwEPt862UK1Q0rYg7UNEPPKJVpqyUh87P+OPQpCv1KbF8mV+C2C/HJTl
IzD/AYaFnhW1SKwXsSqMB1lprX0kOs0G4Sz+zZPTmuYDqEkbEv3Zxfb6Axb8oE0U
f6Jkbzf1ROYZw3LmrpeK1mZsgMT786s+i8mUl4TjIuNiVGp6hkneLTNWVdAEyCB6
kgUVELOV+k9YfLxSuR0ilgjX7rqeFNjBuREzOcjjiDjhaaBF7GzAFAhhlsb3B1kx
5WT9fk35mxDTG7U/bsEy1fT6xYE/Efvxgk555Y8x4LYYpzA5F6aU7l7fTulY0EdN
TJ0ywI4hSgo5ZZealU+vWcsCT0hW73YWgYxuQgY2qEHLZx3ZTOynWOGS2r64zOXo
njleXVZEoXJgS8wun7sqc46eDgSCiomDfhwLOiBkAwfYNYU90/8Xx5yzNIrX4nKr
9PRihEooBVenpYQfkE6LWWjZYdaQec91/aey2rZ5OHmdR9IjvLJjVrqUSckQot1X
MBKzJ4QHK7o0D6x6KLTCNnfwaRUV6Evf6YyCN4tBCxyvwk3KDzVLKspQuXO/5ce5
flfBd//m1QBx/28eMilhtKvHbMuN8twErlIONgStvlzri6XvVjJOfxbDc1Gi/PnY
MPe1dEuKjOEw7V58kheM69Rz+OkVS8JQkAxh3b5Ea59DorRGZ5QMqJnGZfasqrLl
jXBCuW4KhFX1VdCvHOW8FBRToQqfnewBxYLq93WJejGxqGH5GS26tSon3/WLqO8O
5gs6qHNTBroW7kkpIrs7W7KYH+HOfUZxvdsdc+n9NwQm0aJX3o7Hl0o/B4+Afdlh
gvWlskxRxA+h6cl7JV2CxddsDNsZObYPggSDCjxQpxmAALHdhuDe/B6D0pbFThdM
BBmK/f4gOcZqBhtkLJnjXCwynvfv5LhjyXfB7LT/fZLKlUmyPGLo1idY9LhHrP7k
ZTtnJ4RPNVzs+Q4g7SQznwb1BD3FkMrY/4DqU/pIe8WT7yScZx86PCfAhjEO2jqm
bt1vrp/R6UuV3ROgFPsiVmvsmBHaWoPuXdEdtgOttmw+5Qa9ohQ3iqMi4OsmocQe
3/xc9npsQWMdcqCHHFjIXfwWB44ZYe9Mw6naf1czaHvZKwHrT1qAIDEPLRXq1sO7
r4yhP6XFqAGOJbtIgMoZBJ3bcw9hwomZFemJyD3GWPmg+xUD3z8c08cyGZ+SIYC2
iWVQBySr8mKSFS4u0R5RkP5uWFt2F5Fm3DL10N2P11IPMylDPhpmO3YxBVrGKTsK
T+1GzAsrsMgnLBoq/fj0ZBSBi/nN9aMwwAGAUpyAhpKkADIN+8ms5pPyBWHMLYCu
17sq+V/EBoh2LQegxsILTbYIKA9c48JihEvcdpTuzm+6wDXIC8lEakGrYzOy1Nvm
BclPse4GpLjp7BlvkN01kpcyO8gIQfXLMDXGPuVrIrd1spSif1THWwtrJchowabd
NW1bffYvdd2lR6TRGmVAG+JtuDZqFOxmbtOGU5Dl+JQD8bbIhZf8gdxzjsCG+X8L
oTutvop8fLObRPyr/c1z/IIEoJiBzgy4jyvWYtQqi3r1Q2bjlwRAzqk3S9tU4WNM
L5/lYRoDGzRwxw3IGid80+3m7j+WaFS/HU60sbUpBzur/B/oQ2L7U1vNg+5rbheq
r4uwEeFv/Z9K25/ef5EdpLy6y5tXAnM8wqlZYeWg/GHVrvvOyyqONviKbL2yHD5U
+RT/QLCiuFborBDqJm4V+SquseJqL73f9Bvu659j1ymm+atBlhAyXpFWMTi5AzVI
WUlfqRv0/+UgqQYSMj5MNAXOUZQDPIUix8eNi6yera3qKaat7u4gXcnZJVDjL2GO
yC29/LGPlhbKK0PjXPiwBWwgWafqNKkAZ1WerjAj42CgDF++qLHV42cKtQ5Q16oO
wWjyqRBYw8g73AauZx33ctavTreod+ojYNf72MBIVh0sM9jPZbqK5rrGTgt+5QIZ
kyOZZA64caYrlBQhsfrN5lwwXs3OBhTMLO3VGy4ZKfPyT0lypIlmqSaT1zM/zl7w
FMGyq+30yxOqM66sHDGd+kIlNztH7Uj9E4e6jLabGPbj5Fj/zzjpGl5teeSzWZSV
ssWICjmjkfVjASscnJnFUtz6cdmHBB86SgQm4qT5h4ZiB3Ma908j8MY9cKxHar54
LOJABa1fLnd88iKAIAJ1mycGW5y29hlCn4S3fHmDPOcUk5jUsFnvB3MWW1iPooxo
XCYqEcMQNncpK9V9gIreyoLfKdKQwOOfjDDVTUCJr26gw2g6faJ1pM9CGc+dxJH1
5xJEuzyxwBHbbUY7KC2/1+rtCN9QvTesPPVsU7LIujjm95Sxes2Km3wZRtKj8L7a
HvlGmxs21yoz5b9CA520T/TluohkNX8v3ZFQZr0KQ3KsWcvgtmGwZz/VuMWl+NNL
4EdLOKNv6j3VPbHVAGX1EPrU/2lVnD6U9cN/n73AGNdtZg/fY02/7YVsJ6v5aNdG
XEfBQ1IeCpZqEO6cJ44xdh6C04MtZrOoevhNnz01CyWDJSFUzjnbczxBpmqkQxWk
+3oUG8FxZzo49kX6MTcaM9UM4zUP9Xc1xt90PD5UHxj8MOhQFXBE8iR5+6jzsSJQ
fls9fjFjrauQaQsI+Ss9+WO3aOJCJzROfKSxmugXO21Oz7jM6w22DeeNC1+Hl489
RUZvpBjrEfrMe6jABqHRwqAVmFlQRxmWBK6oY2f7AQUWjedkJ0FDTi5A1Np3yoWS
M3sZ3eH3WgBAo3U71+B7NSjmO/za03svXj69jRhGekXgqSHZQ/cM1SHs0GzqxBdq
vE61YifdMjy8wPy3LL6icB4BVXio1j+YBQT0J9ueFJ+RFkZVPIAxMqFt4IDbwb7u
d+jy2FMZ+2yMcI8+vZrwFs0WSWzdX1fqtOicK9rpCfyhUSh9qm9xCNw8/WdY5SAw
rbaq+CE7Zt/zUDx2uzFu5+aOFwUgEepe2cHLYIm72fQWSJ1cYiRRoutIeh9lDgfy
eRFULHYlz0nT9APfioG8l7S98mJ28lGQw2++wUebLdZLZYK/pa+oXcIlojbJkrRS
iU0u9GqVfviyB9SaI0iFIZvl78K5W04t6as4JNIZJsOg5nM++BIumFsGilDiMsNm
3GklDmgjrwAVGP5nqEP+vhs1feMTwxF2mkic6Y7qSGuRx6NQ4oUqMgHfBbiZ05cx
kgOVe8s/4prD1CXpSkKRN8zK85wyujA34W0KW9h87e3a/SsOFYoJj6q/HwbDvwXS
4U/m84XTKk2S31SSLsfganwHTGawil8moxpOZ3iaQkWxWWtEpuPoILreApGqAHMX
P3DOKshuFYFjt+ty5I7vnSSOf09dT/BKQAC2CYGegqtr7SYqzz9PO9nNNuO6M25X
BZ5S5++lHVTJCijdKBT2rqnf1+TOscyPOgAsqvpEw799MmzYX0qMSGyYdKg+tl4m
iM11g1Rog4Xy6mSasqgF4o/nSICB5MHGTpbwjOr/PgRVxg7tU7dq9GbUuhTUf2sw
8xbmDXgWbhoLhpbdWdsLbXaQHS2b+V78cJcatBHMyb+wOgS2HRsfj1piOj1wfFVB
ePEhJLpU7iTYGVMNj466HfA97Htn3zNr81Rf/rJ5pvsnFTyL2t0m7cier108XTfU
+NYKRrOpI6ewiZ6abcK5A6q//nn24m/iFAAwPJDcDoo5NiLs6oAXHNdkJa5p+f5l
9lsp8lqKRdyny5MNYcdmwBcjgaph5VP9NuBjTgcd7N5dHbH02P4axFAj463VLmGs
QwKFSZNA8abJUj7nCTrMrYMMJ4yvcR/sLRIOscdSHv4xD04N8OlrlBeyL2qaZvCJ
D+yL4I/HU67hpDp8wvUrz+dsqCkwb0oSDJjk4+/M5MoMZd5R0jm5W6GtADY/wDJA
c2SLWEsIIij11cbz86rit9iw7amEWjDKTZEr7rXrTJjzTFFcUMeyJOl0N2TmoB7M
2vqFkb+ZILMUtbWQVcStK+3A2isaxmTKyjFWtH3ybXIHafMiLu4GEh9aXsVrWCDT
H/Xfsyk+1z+wp9sJ4kAuQOymOeTTWed03t62xOWDyKHHIg7F4TXHqyUj3owiKwck
dLAVpeNS7lu4QnKSJZSNiRgFcRMGKJHxhtSBQNUDh8lYTS/0KAadAyX0XuvSDsMn
XWF+ewc1eBYawc8T2/0ZmYJP+ow/NFdK0Sg+gfno3dzhTLcIGFkRk8BUuuQy+Cnr
TiwzktB/8T8qeswm18mjKvRhIW3tbMjvQTOhLQChBSKCKvH90+csQtM/YKGtn/PR
Yy7STAOUJQ7jerzN8xM93Jgo78CKBr76u5iSaiJCQxj3NBtTpOFgEem0hsunY6F1
p0/yfGKr/maFeu66hHsnhrTbj+7h86ab3lKa240a5CNX//6rRVTe4G99E7aW/K3W
UuAW77DQLCV4zZpky8OaTweWP1wEcqoov5eb925goo1KdHN8lPmtZA9lQicAj1Ro
ve9ofAFuMgwKyyBhBLumeQrV0HGxVgmDVLTu3Qaeo2FL3jfQEPzU32atMQ15sNrU
TYczdMhkMkfP9FQZD6UYvwe7SKa8yFXYHAUIPwW0y3Lx0gQ8hrlPqAluJ5SNMSCY
DwRb/bE6xE9yyjNAXzrd/O6WiHIBp6+1eqcbsDgkWZphQkVUns3qZzJZJ4zXK8wK
svyX8Kot5GBazgH/mHnKSxav+3MSYHVT3YJxgVry9ug38KJFIInQZZviDk6U/yxe
K0K7hYBN11s66j7tADEx7WF/L2hfLOIVhr9jH/GoUOT5f/Dg6jrJU9fuXvNj5Qcq
BZvbISRg+rkmQRDW3zEw6EjFvs3K2LuW1s6vI0ilMzehv4hRidcxmJ6yfqAoxxpn
+MdXJXy+hQqlOl9l6IwYuwTEQxoyFeXuE4P3z7PH/Iz49FFdA9FJQqQopoV/bDSz
owPLwp6pEDPpgVMJSZKQT8m6cuVJwcDpwQwIAWSJiFjFR1H+s5HkFySySLXCX95o
5UzCHXudj7jgrlNzmsywJ/px0OSRLlTE8OSl+drT/Tsv5rtsFLUV6/Ij4ycrUB4g
GN37JYjxT/pqC2//BtKAjDlx3ipcBmaDjAC8yN/eVlPoPebn62w+nejGbhOLp/si
gwAaiWL8kfv+K5vlSA6zMHFXZV1aGzs9WFRYnhWfmAO3zJ/INJDOksQxHhgYutqm
EC0Pnzer/Fj1AayvIlCOS6DD7MTcNap2Xle9Csd7OGxAa4h+nvEXN1pDwnCejXxu
ZV6uwSBXJlexg+ptXWweshRbdXeU2HHKJ0pE9hemZ3HMiQ8nsn0iWPA9NxGKH03c
nn2hMVazvw8JXGpvMK6VXq0R+p8wt3QAzYqI1jGR5X/2+3mLnlab1Ts3sTBYQXhi
oaj5tJ49CfrsSnp99xmkrOTr8CaRiT/hDLLjL4bHmycpXUXAUSqEDtlmJ24zLTHq
HeldQERRT3VaDoeXjvd0LgsVOfiN0rTFq6gZ0l+tBB0qFA7jVaR1I5M17T2qfUEK
cbSxExxXC2kp8dOsFlqEsVZNUV31nGvdgcapgc+rv14cbIL3uRRPVVdtawOAdnTH
oSNqXSxPmYI1nCws91gE9EeAbais+mlq/H2qvaXzTPhLWaWA73sBaVEZVO6ykk6q
9Y8tA5lw0XKGtkvTDTXHKlAmdSzryHebT3ppCTqZ4pkpa9gnOCsIh4dzzlFm6qfQ
DO5XixDPiH8lMpcS8cHTM0MIU356j0/hP+KlJaVUuzQM3OVTRRI6HoZ7ulZqEuoy
QOLkt4ivplaVX3+k0xC74BoDBrzIZJ2yP/61IB8QjI5FaVAha/UyKOR8t4S8WaGW
XTSBS9hhy4YQRSsxJl+NRbma583qCPAn6SITtnPJAKJAuKOnbosWbTfXJo4x+Ulv
RghqVV+TPgq0NakuS4Ynpy3htYb2GU6R2gnHh990pVI5J4w3/+rNWP+Cy3sOHBt4
FaZhkSC3NacQb4UPeHIsoY5selTils55TVp278CgrMrpeVavXtoF6uRjXV3q/3qw
kxbZOrdXgUn+DcX7lFn6MPx0r6wzXbbUdMHk2tF/3FaZjO5dtpJRXjE7yNdTaZ66
g6RBjwNlouzn8Klmnxy9JLz/I7MiEQeCNP9NLG4sNzUSTNe1EYnZwPs1H04Gkbsh
HnHzEeLLHHCW2vINpUvKK4nIYibAz5DmY2l2iXoOGo/aW8P4IqdOXgwC81KAHmVE
gVw5BLHDaScMS0S1AUqXG/pXJTqgw/tepKXBguOQ56W6OSdGksNUIW1R5B3GvLd8
VhKcoai0GC3UdT1eTWadXFfcF3xWYnM8m73nJ4gVGsIb6Fj14z1L+Pu0FB6HP09i
JyhN+cqb7z9te5xVzR2olr3AlkmH0x1pGhG1ELnZK3VihbletFspLISleCuuZZp6
iaVa7Ku5INCQbnFQusD7yk/3cI4lSu2ve/XL7nPtFLK3wYLt3suWbB7PiAbZ5GKq
qUWaEHf9uhU5mBCYRtvCXG6fCGjkdPgW/iUGLdmfJghFpeQszGHwSw5fr2ig2zI3
Q4G2tkkDK6fk6ozntepddv1lIeUWDl4S1R5LJ9o0vDwSbZMPjpmvJM5/C5FZb5pw
FN46w01LvPM9H4bLku5polOV+oGjkIn9q41tA3p3XmRdQsXYT7Zzf+aFV9XP6xrR
IT29to8nLkEOK+akdvN3ovbA+fQ/FddrijIhxpEaWC97+ExTQhk4ZtXy1VuFD57V
EaO43Zl7XNapIdltQdXvaAwlvGYUJ5TfN9XFVuLBYZFm87IIlGz1dpvRB6gqMl0E
Es1I+j7nvAoZfGTjBJg45joMGPq0wVQevXoh70Wavf0RbqbRqh+mBfY703w9weG1
B2w1Ve6sOOPsttuOcEPmgvyaZORQegsmMlRwlhvuyL8vsT4VlXPzqzzrwzKxgD14
OQ81yJYPqzoP14MGFbj597FXwmAkQaVVkHS0W02nzwPhyrcbFu1SvdIiUX3ffAT6
ILT2d509OiE8ioxhOf5ZB9c2Kk/+q7SJW6TJjdzWcHc1fnrpWeMBawoJdDd07ZBL
cr3ZhBRspYgiSHNIWRiHiOXZB8/Z57VLIdmlRZ9f0KtlQ8zqdca38/kYrkhKnkpW
2q1SZBRfw1f5etFuA2WixkH8sWF0KoAbSMoDFFA+WYsqnFRYhPBHXhyjFZ6WsmEd
a6DhkSNH2cgCzU05U+UEeptzWGJPsv+a7uyr9VpIM8MTEr/4lcKwmmVLzCbokSI6
xgbZ7L+bStTGNeJgCxiO1oIW81cCxgMgzYva5cVRIIpmFsAmvfl1hFtzYQ7+etvy
IUmvnzO7+GrIT6JwUGAY7ZA3N+dEfBXDsGZ8eSQCeaWRrulP0EvXuM7KxozMbVoJ
XYNj7C6toK7/0fQs8sox+K8ZHntftUBhgRhYzIk7cE/AkuP9wrLVgUjRgRPxWuCZ
XkVObdmaf0r956NNgvRUg2zK8qlLm5g8G84mfz2rRrszt5Oh+M3/oE9FimnmgbFm
0p6ZjkcPkV2TN4gm6t1XpxPE8tUwKWMRLOAIIOCtBCC0MMf/mt4hoVWzbJC4P8Hu
Wtk9OBb/BA4NAhU3dQQGP96y5KSkpkZOIKnNPCiJity22zL3weOvf4PPCuNwXy6L
nHHHQGJgY5zX6fHIL27n5NQaDCLDYOQNy3N/8oG/PsEwCCRdB4YzAKqi4lYgF5TI
YX898/x4Mq2t98LAT/opQnlmdDzas7U6/FnZEoI19aMTwEVGHa1kg1bd+NGMfHSK
B/xErZefBZzwOfYWQFFMppmrZ5EFDc7fPELGRykCLdPChw1hu1ig8j7I/G2e7wkx
dNHLsBVjthbUUevq3pmpiC54CL+EGvib4XAvEXdwr6D56oirok+OXxwuILJkN4yI
v+5I5gcdE8DHxYRuejAUcqrVJ2ut/xsdUO7HIBgTXPEN62YUjCf886LdEaI2fEXs
KUfj8VMM0TmR5i6rL3fFGfOyuFPtebZyGjc9UdD03xlI3lCx7JWXJzPfP3bUzynF
k8xz2Uk4iu5Mok+lPM7CTOA0N2xTBcgkjfbYzBAxVQteVc58eTeQYU39dFmeJG6R
VhAqNgQFP4ea0oAbDxfyK2IJo4Vupn8KArJE50pkqMNpbPBCcI+K+9nCIZ9jA0xN
xiP8gIad7Gop8qAhtXqDm8KCaQfff0fu7m06M8xCgvyubNavoZP8lMV69n2L5Lam
`pragma protect end_protected
