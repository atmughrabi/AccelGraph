��/  ������0��l%�~j.��i��!g�CP6/�c�e��J���zF�Ƨ&"�!�*vaMd󰺨(ت��n3�Jk�ؚ�W����4��XY6�S6G��8�M��
X��7\t���:�Z"�9Έ���ӳ����?��[�z3T]��R����<��}���Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9��	/�%4 }z�9���eo��wl��%�-���k�L貹�jA�	�;K�EB3i;��ܠ��T{�TU�x�"(Q��d&q��Pq����K��x�נs���`m3:]b���Za�������tg��3��޻�����9���$�� t������f7T���~p4k�I]ӛ	�T�diB�8='�d�eG�2�6bO�	PQکwin]ܱ/s�����s�`p)#��
�c1�F���bNs��%u.���v�6�o.����F���{�?yJ��?�0������k�3��E�0�<nP�|�M�P���dU���N۶����Z�2|�C�b�'�K�Z�n2+�M$z�s�y̬7{Z	����՟VW��j<�&u�lSK_mK��FȒH�o��E��Ėb��~�E~�܉�j6o!�b;ǆ�]S��b�z[�/�[9�FϏ(���/�l`������{�^�"�����N�W�����z�~ �߮�]�̢����%�M��	�h��
myr���Z�i��Z'ײ��Ꮥ>z^�d<ҹ ��喼'�`>�FF]���H4#�������s�*MWZn'ZO�zv�g��C�'ۥ�|��qg�I��pQ���uy�h�N�f�i��AUh�u!�0u��{����9�G������AЖ�����ឱ�i�aGU�(ϗeE
ӽ,���ݗNt;;��v�㊺�!�44�U��T/�{<���i�:�u��{������^�8�>��솺����꛴�Oz>Ø��:RzU����<�m���+�3il!��Z���
�3���{�?<�]"�v� U�@��'��D=����P�2nzz����gp����,z{�gJ�g��'�(8�h�T@��`��$4H��H3���d7c�\df7�+x�Q�M�BЅ��F�~��Q{�8��9R<�����p��Ir��*�~&9❢��dO�J�fBa������