// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ecv+CoSGNQgNFknUsO+Yw4xJ1yuZYO2pNUbgJrIA2Cp/ovY/hOiiScRlrQQpXu03
p/QCRDI1advMZt0Kk3n+GitDJZGRx35imJ59RESNWacpw4DgMl0P6qC0qRpTbZix
yKMbkPuCfqG95eKWlqPFfgkwtBSU30Hjm9rbYgvmqkw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8448)
T5MH5EgUWOZpTRepcAQC3GVCyln/qZtBo/43j7e0I9cL56hRH1QCf3Bd8RBygVCJ
G4uY+5/mpMVW0TygTtomxtP2TW6e/K1PftuvALXRJxpAQ4y9yxqlUMF/wNIbvFTK
rvoIU0p9jmGVeooAyJ/Q0bl80bbS3Latso75J6+Al9sKdH1n18FsCB08DAWTofVK
EWluUqe2M/ekxKIDYU/oFPAqhBYiiXVBgCbvrMRwCCOjHxww73Y8eFt3xgGZlbR1
TG31Wiq58CCgcfxWCM3ZgEcpcqpj+ejattmG7PDvSVwGY42MseYfUbzKcVvbG2a9
QM3TUyug6Ge6cdV9kdeaIVRtme85QRMjrEkeUddXrhau0ufNfOcUVouKwjJ5brVi
A1RcSK0Sd6bsVq4ohkRxffzI9/TMIEn6NXlJCpEa89FL7cmEn3bAZhlCfGG6h4+F
hBScW/HvHTtW+8MxAq0DomiDJpO96fhN+485MGxxSulAYgfL7DYMtP2OVzQdikti
kdcECoqHZKWUFlCbe/Ytf9LM1WA7oM2FB6mTszlx5fufuycRgk7SoWbXpoTuMzaI
bme5eC8cnRqpP9VCQaYoLLaCIgoXpv72CeVWfWeFi7emI6Ec9mpgEF6AekyGS+Fm
BxU6TM1UVQI1WK0FZ1np21Pjr6IpFi6l1AFfcPcdr1GGt/zaTR4nPSH9z7QqDDhh
f8V6u10DNlxTxAuix7MNb7SpwE4L+/jCnJL94k/2YH0O1brQVwsrb6SRO9+skZoK
9oW2RS/WfoKtLAjU4m73ne/HLHihI6D57KqhB6dlU/sM7r/XyzVKK01gwj3ClDIm
sqi9/rq0S23ywIYVfeQWBNxhkAbjhCQ0JbFDI/5cYEzAmRe3ToT/nbi6BgrqBLUf
PzwEVfA7qtz6RDw6oOpOMVpuvkI9VWiPctZXt6JjnbUMu3wOcfUQDodN+FDkUx2T
HchgZII6XzbfeBdiIocnsQ6OcQSK8W9UhAfjC/g/1ROkmTOc/mwAx33aNmXsnG6Y
lGiCBkic1kM/DE+Owd/8Z8MP+y3BbCoyGF3dpkIapK1MA+dtPCkbmrebLzYH7HFb
v0hkgkRIlnFyEdZ8woYUZ89RG0XMbLxChOoY348K6S7j4nm2FSu/XuvWfYlmTzcR
Ox6rXISEmnx1vPQuncsE7wOS9i6AFGg6aT7+mcp329HaVB7xHNEdonGbH1oGdDpj
AEOIyV1tX6H6suiGbvOIyPk7dduXOiMZglrFAQsxGyl7s0KVfevWTbsYTAnWZMun
hPMTnzeidpJ1qofgkI9GpOm0ugHt+Aic/13Yrz153ahPRm9mzpekPoygNdSXyy5v
TeNCK90jWMQMoE6Tbq6kRTUct6/AQTtEO1he7SVv4ffq6bQO5PL4Of8Zwa1JHjU0
2tbt8ilP27MQuy9MH8xT92Y+cD+jd0+8mZlbEWwdZfL/Vv2gTJ/c25+SHNSc2Rq1
A5q05fGWl4GN5vfPYkKuAHRk+lIObX/WfGRZasg/ofGaemmtomZ9QfGBvzdcduye
LQ6fiPj3Oy8t/nym3T8axrF5lzJzM/XUrOjyL/cwd+wlcva7uUNuGvgXlxHujsRn
4dIqSvFvqySr7RcDYxx61Rh1fpBC+0MTUtcn82VBtJegRt4dl5iPyAn3oit2goCv
RHt4uO5g8fj2uJPUTEiJblfnj7/Z80z09FMBlMmXAl6BQylcjzXQTfsw7UIm9UkW
RHXDs0WY6OxhxvwAkTqVjf9VGYCkiVK0Cf6T+5CHSN5Xe6yIAjgMxldAYexkWOuv
szsWgMJSAj9M9rlgHjU151wvxkwvhjdPMdqbc41AtIqT4GWwcehA/E1Jnau7zL/z
eVjlqdA+yyUEu+f6FLd0k5ERZPTgjIWNWl+9+9KnmqRhFj5VM281G0KAMfH0oD3I
92cpgyngVjMJI+G/xZKKQFctWAAEJboKMhwiFNANdo6T1MPfAdbMsYlLlB8S79dZ
ENKbJDulLLhKoLHpl8QRN0mXlozx4Ir7HlgH1ztnq3a1FvFIPDgReMGAlwZMVD0a
Gp4D40l6ARMTNuxQch8aDmq/0GLSVYQPR7TTJPogbF8Vvy+xLL25AULAg6KduBJ+
KMm9dqIfdvwSQjgDJPqTn2mmbsD6i+cK7RvLCCNvtzJZAkH/3Gm+A33T3F4X7UbM
2gXHt3qgH+VyAVPw/cQJRtM/npIGLRUc7bzM5fwwkYieWvreKtYqHrATr42G6bE0
lHw9zxLcHmdcYaiEzzPL9WzQkU3++jSmhwhVA0XFKb1p9JZG+Rh9/tEjRH9jf/U6
dhG9nGRKgZod95OAHkvfgMobHBPhT+5LL04rcGKrTLXIkKlAsEYOXGTehJw3Q10z
arqGffTyZVA+qcNg82Ovc+kLrE4PH4OfmZdXRZHRChmWJ+8to16sM8A+CO2SdT6W
tSWMFRX7p+DgyLdiGnpqaJw4djfpneowNz0SSWp2gchpaetnR15oB37bwCwU36qX
0FONKmTwomVHMikkrwz+/Y0jymL7apRtbm/NLPti4UHQwV5VXl3rk3FEDHTjCwUf
kqIZ5En0WM05oXkoMyM6HRtRqH/j9h3xtlA71+V4clvnHYquNNBFw/oFNHJFjOvB
zxrBjdQToWd1fkhtdQ3gKOSE/5JlA60kOJPbDBgX8ZZykiZrf5QCaXc3vyyXaH01
VYKllz3eiRHGpZtlH/YoXXSgr9YxDbTAGLAsMPiz150rawWotto/Zal3FyMqmtoz
C4tx7Dx/WYONAFfVCbHtU8PBq+xqpfFiTvcCJ/sLDv4Q5x93/J+y7Ne5+dvzz7fc
1nP6bnL4h1oXpwDjcQOusK+9WyGayD9kzTTZeDj4+fCe6G90WbMU3yN9mPOEs+1/
zSnQWnzf1aBWB6nT8NZ7RJmfBnXg8wVN2+gNu7/tg5yknKkxVRSjk4ppMM9z0gd/
oPDVm4MBiclcCRC77+4XsmjxCpZFpXVZcTY7SqO3p7Ds747H9aiDC4nNmxGwa7CY
UpuAO8GkPAMWkJa+s8J4+/jpkaZBti/hZ2w9+WLGJOZ7m9u5v5D7K8Xy1/6gMUlV
wfqcGAclc7JIwqKLkkMDwXlMCq3tUPbiynlXDCNRZoWqNTGAQ8aeOvEIR5Dri2hu
ir8eE4NJ/0WnahkZ4gxHaWfiGa7ZCjxjbhvwXKPBO8ezhw4XiKl3HnAoJ5UiyeLx
Y79lkXJD4rTJ1+nCA5fCTVa8Ped7WB7K3JvCQvAoed78cNmcklToNXwJ7Le1pCHR
qz3bsP2JU1lQHmQbVHFTVFh4gwv6QozjMjgq6R0L7D9amej8hk3xSbMSw8ylvv1m
CHBlbmUuy1IcZMkKWqwusJSk9zrGGgy6DXkmadNKKiJJOZx5DMPak+Uz7PVzHTk5
Vf6CmTlYMlr3fqRNybjG+1KuCzO3J6l0d5QLrkPsu4vE2f1TqMVD3tpaOxzLt+t5
Mv+riRm59eGMKVSaWdholSiuyXs2BiiYSQp/j8YyQYLNAi/GPXj6AkfGQLr/GW94
1zS1J7IanxqiuKlpKvgOQfZ9Ox0u2I0I/K9IZd2K2sDCVq56lF1mW+oGO4YikUvo
TbNRkiU/cK8QAF6BDvPlAWCMXb7h6w0g/8NV9fjl6HwZ4t+N2OOb2wHEWDgTqBSZ
mzCQWGm4/D9Fl9jphpXiGsKNbkKuqi+PbY0UYOEH8/3nYtDInKJUfrmvNO4OuQnZ
7gUhV61KHijk0AQ8xmCL4cQ4LDSY3XCOO7+Mkqauw7BWwekHlPv8xGnuoSb7XPCW
ePh1rljBK6D4ak0G+l0qTp+RliIPbLME24+UGetpvdrryYjjxHYXV42Pcvr0amG4
zVsF61iOXcjXQtl2OWQdi84N6svGFjrYDv93bsJR77Z0pHyY/vA7m9zDbxCCRHV4
nfwrXQTWagTwwvcOjzFfJhrO4PwpSCPdzVuqioKBZDOyUUbwP8rWuq9TJmyOrCzh
bVQVTSDb7hueK1eLEVSPufGKy32wy0k+Qj/VVzW0KUC/GZvzMvkj0eZT2Im65Vve
fA1UN3RWgcI7uJos6xWXzBu7KuVDjqPX5PZE1tke8n3VZt/X70aslzTZjB3XPnSa
3hRbSPrzDcmVxEFKdC7tfsS5wo+7oig/01I4NZ3SukgthJfxyVQ8IRAKOpXOg20x
yFQRI4cg747/DlOX5ym7rh2WpVlLlxpKqZCeJr6Q54YFD59QXw3hQg6t8UGPsZQx
Aj9WwxAjwsdt2rwF0b7BmRowJKx6k/Z1Aezh+c8sgLMV7auTH/lp+6CeOE41kLTj
/fn/8AkH2mznr77ee99eUk4NvK3yCNc6uh3zHNLdiSF7ql0jwd3fQHzvRPm3hOkW
SiU748O9JUhittqvzEzPNL4j/AaIntqycUOTfSeTjLLk0iJ4KlOr8+xbsns0TR9p
GXkWRUhx++Ueg8B/KaGrfUjtAGmcyBV8cZLgK9xHj1boXF+jZ3ZtAWIjDCk51lMi
Oyg5H9DNAelM/2xG9hwdMreSLJcDQ8de/ayGdePtqThdh+zrjX8OtxZo6OW1Ounm
Vj4VZe3s3DrlbNzIqH1t/ne62E5KGXMbkrLqReJY2wEnOclTBvYue+Kkhp/jVtiB
aD+1z/Wgv5Fj6o9tdzywnw9ziJF/tQnCOwq4S25S0qz9lHBCDyhL1yxjrBo9dnGF
AirkKPAdKcAEYQFeb89OKAMT6tNbEOMcj7+NkvELsPspsELLvC7bf/LMIXw66mYO
AcoEfW30snb0nOTGXDDfNcMAPrQCWhhvThcoBy25OMYqc1UmfizviAb6GgoWKL+h
cxs0A6fHIUzoI4p4fwOp1eG9O0N8BJmGnA1b/sjpgAE0239VpN3sqAVIL7KfqtqF
ycXmviWszZsz7hjJ4y1lBkfqQcDaxCHeG/18V9GJwpj6FcVJeergg/fw4dThS48I
L2d3Oc3prPpSbJebitpb+qCebGbXj1LHHwZegJAuimmjta3ndvj4YlHWChRin0vz
OHdT8jYcUmdbMWi0QWg/7PCqkJMz601ieCaSqxD1aIVC9iYzf4X/3VkX7Yx3j/ka
937/nORdGygK6Ztwucvi9V0DcmvhquF3GXakaKxqQLu/5wT3Dgj0YhRz4/Wa7YVm
9nEIxYRfnJCqTpbTMleASigSbPGHKcwCVOAIhCGr2fWl0LW++sK7PR4X6ZSskRq8
9tWwQRp8sGi4BnSBGThIpZgUpl271ELU6zzft0ic20ZIX3JboTO2pF9DjHuMT09Q
sCDnfRBxR2t4nJdlnXcXiq18wo5EB7VgP8+ZVPMxoMHbp4+/99BfzMV0ak8jXaoe
J8b93pZfvu76EBL2VBC/66/PNir05cJ3spDQaTP3NmINTRGKk1EZI3NKSDJgxm6q
g579W+tnaCayNgDOZAWi0SR9Xs474tx06V74CjVYvibkE3+L0VLkTgl8xKK/O/th
Qxg6jTHO/nDz22A7vZtW6x3xRhcoXpdeLkuiixZOEqmSvaF8/J0c/HGZhUBxpZiY
CmXQ67t18IIaM2KbfjbG8r4WBHEycJEsD4oa8BPUi4Xhy3a2oQfLOp+9rPnT7UTB
R5B3xE0tcAPzl2hbG91LfjQUlNwBcD6fv15JlToTLSlnHaSx/wnsKbuzQbdJlJI7
L/PXOJxFAlXk78NS4Z7bfmGb9121u8qEvxwBFR5jFFI8GIW83jm48kVPfm4AWWX5
alfRXbnBqK2N/VLNVsK4LH/M1kFsTNoU/MAGFpI4YJeBdwuVzfb21BI3qPl5zrWL
DvhIAaWVEHBFPmIH+kslYEQYsbWfaOnYMhUWJRI/XJQVxMxLqMkKeCAtw46tO1gT
iy/C+01ZI3qvNtiM2Wl4I9T0Tiqr8BmezyTBEK0hZi4w0RUD+iIomMqFU2c+8ynm
Q0hx1ngbAAOKQz6LLpnUoaTTYv0bJdKHES4TIPwVMxzve/tshqoosyFmjf6K6N9V
IZgUuRoaEVm/20HV14oj1e6yC5HyA+cEoGG5LZoZuuXK07VEc+O1wFZtymvDVKu+
HH6da3IzqNi3IqvcisQdKuJS6tNFwPWpcej9gdgjOtdXYixjQwfIcYBTszAlKRm3
xA4mLEfgGAbn916McDdYMMvk5D0tHP/TsnNOV24CO4yTj+2NEjs8HGwX3O1mpkso
eqsO5QzNf3h/pxtfrnCRNa1tUHFWikgxdlKVWlFPVhXqv4UNDRoRBz73J32nlkMm
CP11T5QiA5/LGZhTcR9ISd8uTvJJe7++Sc+2Ii8MlZmTVdsxZkvoVHEqrSPrPEOJ
OPU4XQ/RhZ+RinKEYy/qudK2xmKftrKTUfI8KXDY6zwafTzmxr96d8aF/vMsGstW
LiZ6WZXsV9aNz2u02aKmXjSHRWfMVYFlpAFan9DhodvLnHhYl7pP+636cFfWJK9E
C4oXQiK00YAIwHuabsiKAq4HvUqm0cAoT4IkwRGWL9bLLj6EKmAoJdxZdEoaYNtk
jN1pkXXguaQTfjRntLV4OYc55r8vtOTy55XXoymiZupDcPgj6GGT0WOdT81hTzjW
BhFLm3m3STdjh00LNgObj3pX2OabiTojX7cA01zKaxV3UUHL0m5J2qGsstVsXcm6
3R6tJpaFg4YMSy5RTwoOxWLbtwM1Dqpn6pRsp5UEqrokc4Q0NFffQpIGy3C3yC7O
LSitdsvS5Z8z9v2ohDDn7xTPYshg5MNwOksEJtAS1LSpzqpxnJBJjiYRNQdljma0
sksnLifCQnoyPNc5qh4TXMdCQO6QVbbrLfSTXIgUOa7MGRRHkArXZd8gfjuydZ5P
yQF1eT0BX2gO45O3Ni+/7hvz6tLoNeqiBwmclA/oxnvqeMsRAmpNC0OxrobrxJLt
nZOiSTIwLb1kWciAb9ihdeb7ANByIQ08bZQeWtY3ph5G3nuT+MWM0eILq5pCwHEL
URhog/jX3m3j7L7p/ICSsSCJiuUTuSGafD6HzAbn6Q6i/pzJEjCBNW4M6C1+fOs0
vxJRlvoSg1LCECXeXuPGpLwsrGh6+Vp6jS+mcqbKtmWImeWrqemMREWgPW5fqaBl
Cwz/hSszBLJnrPI+EvCNTa3urbzkS3KBitiitqNjRXWnh4ig0ucdBJGZ9u2HF0PE
pMTZ/yoQqG1V6eTDoQvLU0Z4V58Ca6gVRVOxabq98yx+t4sxqdW8QRShQrOlAbwT
iv0pZyLcKaqr4JHJccjdI5wj39XphdGI6+oyx5tjlWvXLQhMjggAwYtxU4jNBfAA
rSO3PQDquRpmpr4opbEYWGmlwfhu/h/SYt+4l9hwiFHeCYprnHspV2KL7KfbOBX3
3lY3UjRQPJIMdoS6Qcoi3gv0kRJG+6DWzWNAeYZRHR6CGRizlapPDS3m18JpGk9O
Wkw8aJRBpjNZIxgvkFzkLDUJPz3rgO7/tx8w0v2rdpnCgEggstIAzWyU8g/6/VJ9
+HNKoaUvaPxmqwaCIqeMND1xQ7ALASW9+4L3XW3oCwiVPuV+sUQOSrsMUz8fhH4z
BD2wBNOCBbyqt+nx9ZvoaLHsT+L+Dr2mvsvrSH2G1DEH/xlEPL2pQQ4UDVd7AFAA
/2utcp3RBXk6wteehBHrO+xJMQBWotQDhkTsWArYS8uFJoX11lsqhXEKqkLbTTeN
VUpuZX2GrBknnv/LSDXTEskR8C6xNZxDbqzEOkUo5TAHRrPvlFyr4cBKeRN1DXmw
aBg8T/wLUdgIsGfiO2K1YpDkVrupuOVKGXGKpUSC9+HCWSavu1IVzfNz0dRD/Sik
diCkoH4iM33gNpMD7Miz/nbz8QMVNGQf+Zve7gevbNIwPL3Pczu7jqZXpWpYhkKC
9h8L9Jv61aG7O+NQPAVOChuBa0pslE3FLMPqK8wjThsGQTtSeTagBAYKsy6xPrsq
jU5KfXqs9iYUXij3EMHXrkCZNPn6RnH/6lYlhMTDKXTAHdswO/6fdQfuf222Fn8n
+HaGwjt2pKprowVq6gxNHovH22uPMrUebkZWzEC2aVdyhKdvkHlMXmrUdakuWVQT
+WtLnl+nNM+DdewaBAS9xDXAysqlh9V70dtMRLlZyGOb/KaPOJRthydNzzgyErcJ
U3MqJncf9vvMv7W/HPyNslzkZZFKnVTsr3oDo1yPaWTAFP7RVl8ogAtj/tiX2zb/
Tj1K2K0fDvr+FRMQxBdoYe6Y49AFlkBE9Q2DCj//iqhzJ2GpnIIpSL8QgTav7jzO
3PGj0gXqJs4r9XUgXvOagl68dZSfZ2czuPqrb53m2oBvnrAfeq0E9rDJF97SYXHG
GzZGM+aNJyqOw9ORryGHRUxKGTvhXJu30SZEaL1kN5vWuPLRt+Q7PONnon6UTMv6
Cq8CfVyAmxAIaFxgdVnWyyMyJfHyQv8xbu1iNqXFLT0reol0ysxQLRbz/0MtcWRU
0li2OjWc+C3Kq/YaBMU0MW/2fALm0doJNOdsqQ3AkBql9cUsOjS15c6colQZhMf+
yu7ZUsEb+oZNSyTUHP5KXMvhesFqW/fSyp7QqTj9AMKJnV6+xjG1Tlz64DNunHAG
7U0ZpDlPlpnPUTk6c6YX+dhwHd4sw0ncVkw3c23wAWT1i/S/K516UryVnAcz+qWN
aE2yeYW5Blsnhn8j+Vy+qoU7BCQAm1JFB5nF2LvFjbjU9UeVBY55i8xhqmlQqvzj
66r371LkjkShTL27N02te1HS27FmO921YCIiMsAD37n9CU6qa2gI/AuatV7lEoqT
sj+WCLkO8YGJVftI/cza3Ro6uTI2hbLQZvJXSz25Pl11im9Cd8eZcLr31IAHl+K2
AFJifviNe8i9ooaijxxLbZE6hGhYggEhwiuGuE7v/dIzyHPgkYhm7D/FirC41YTR
pDrhUs39Z8tdkev5F2YS8NFcHbbOZ0S7siern4jjS8OR/YNNAoIaa5kQ+rOEGuSe
fiibzl8Y8yOS//ESxZFqh7ntfOzff+HM7hTG9duq2maFjivTfBp2550NffouV8Yb
zhcCz6kbNbYM94chFpKVlv1Fz3DTCT+1Uz0BwbSDUN2ygDZmJsi5QWuTUuq/y1W1
EULiaR/4FGAbBuxYaTthY+7k70XInA/mBkUycYZWTQf2nZKJ3et/m9c7h/kTUfoN
4jiQ2sM8/gKs66r6KUXUPcGThEFHB3bqWYWjscaYIBODgMt/akjXVby4GGJb7Nhc
97uw4yXSCp0vUhf40VRy4K7ddwknCtUwi2d7SJPpKfNnaE5QTRdNUChabrcKa8Jj
axInMChoFXwf2zyuClVREpPLo9dtMxR0LLFUyq4J4iHvUAgcYzT39CO9YSiRFvJl
hJKRI+rhO5qnyfxhIHI9UO5VojlC99wYJtFlwZatHYc/cYofYTVIxgv7/NyHF5PS
AehvBIG+epxG/vZRT1facQlytBQzRefoBUN2Dc+TvqxyUsO+LH9UiK2WajJyMSKs
0k8OUckkfb9l0iRXZ8CFqGuTK/uTlfrekJwRJCzZszi7stihfHr3xPYPXjI4nVU/
cfTzB0RwYXcrMC/OIvsc58dolwN3rlLqcJBJ/e7cNWxx7kev2RiV7SqL1xEvu6xp
rizTcvEktt2h5HD5YHeorvcImJYwfWz/txJmmebriDXPtTDZct2iHPaEv24m05Ji
pUPHJT2X2g2psEYFwCHcFkKhNs6UbsUwsPDAqhCnvRitjnRKPcwhPseEDyJjWsik
ZNt4Zz/IFwMb3zgHX83NUB37S/2t1r0T20Sh0TgtwGq6R7Nik/givLR8KZsji9J/
sZ75Vtu13qgyzSMZV53tN7BNbhAJUhf4YWNxM/E+09c2VdMRtmyCFLDaTcfJfhEC
J5Z5m1v9DrUN9sTKvYZMeJeGmMblMC+TapLMM06EC/uqI/Knv0f4+Si0WLx9vPCt
cwSwYWmoRkM+9WU7TB1skmM9z4OWTxhsn8d+evU3bPd3MaahjEGEBrYI/P8BeXnt
xVhtO2P6ROPVMt08Zk91d/I1QDU3DhU/jgwIhcvp+CuLroWUIwOCfOQpp3C1/i04
zukcMUE4qtftxQRDX3UaDga5dDPXRZu2cdBkafNeusFSyWridxTFN7V4aid9sCya
iYRYZMEDNzhk9Gj+nvR3Xhhut8XYuPoDrzZhAJhPkKOCAZBPPhFNpQiIRoqZHmZz
ordHrBQS/u2WbjCIxBJpnsaQ/uN5I+tJ25qoCaXsyIAp7hRAH3P3OtamiiiJm8Dg
iHoAYGyxT1qnbCimOsr+rldxnkNlarma8zFxxNO7mMWq2ImvjpHbOsefcYPwhOaK
tfI3zrRjRXM9LlzPorRGoB3Q7YN8vxNk/HKbkEsqRvJBayYO37bGfYaQGMfTBdJD
/n0kYJdr5OPjy69eJ7KEY2YXG8Hgm3A39SCbRF0Q5aBsarS3eB5pApGZ4mDlrtXj
+xSvZkkeMdEWuGDMWFu4SKwPLzDPav+p36WtqR8KdVTMCjmZATOB/J4VPQMigbrX
Fv3eUofWCGZLqsK4RMl1Sf7e64b4ttxmKH1pCke7plKIXw4E7Ft+fxQFa18hCbFU
Ntx1im4EFfiYsbowQPFTThZBtOsQM+F9AyARKWFmYN1IVCpuU5iFxlZ/3KBouCTO
SjuiJ5NKU2zpNW28kQR1sWf2Tg2VVyvEWfbU+pwPwCCp8kODxtrQ4+jCw5J4WdoF
cEhTlrtaZ4uBrlgrBwGGbn8pDCN3YDFWMQVK28O0iSsMMS+/uMnH2cyH10Qbo6Ow
sRekZHWPkPJRozrCpzrHNY5jdkv88cRuotBZr8TrGoFE4eSulP30q+cIFodIsti1
gRTkPZjV6lrudBXkB8VYgojeKNKcJ84Qn8iWF0lZ7Kd7IPQelUcrPwy9UrLWbJh1
02McWox5UhUasoT2AirGOx6AuV7CLZ9oCAL/Co7JtJQf1ve/EZULV0oLEFEuaEjO
K+c4uANkdtq9Ylq+w4Ycoiuhh8q2p3AoVPUONI34HdFEo7xYnO8T9Z84qGEcEqZm
+Y+jBxA7Ec5EZ8eGmX10TlzLGTgsvJRgXpUI2EE4vr+uSyaHeRH3yOBbxNdCXwx2
hl8/L1zgWSB+acHCBw/Vv/P0AmCFQzivIi0uebi6V6R0HYCIA5M6h5D1r9aQmwgL
sIXG4ZaxQeiLDJoT3X6qMGCHm9KQC/U1+lHHq8Xh+mx2vILR7A6wxZHous86s8HA
1IivOouXoKDncuFRu52BnkpUfnjGByKx0erZS9B1V6lKAMiNmnOSaee1tBAKX+GP
qGzqs3yJRVmz0IMWnxYQdPBHP8VVJIfSXs7gsa3Fb0Un9pTlfeX38U9YviJ76BJL
`pragma protect end_protected
