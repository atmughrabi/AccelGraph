// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BFURFyCJcaGScm2pgkImne61omJ+Vh894abmHqdJ2qsmzbDGNeX05nN0pXnirA/6
vpTV/XkpeZ3aC8ho1CI+msorlwY8sqpDFqGWZZKASJhlllpWjvkoBdKvuoVDSstL
WAdsu/BpU+8ii8P2J1mqNT0zURqQDjiOZEHQa6G7xJg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6352)
13j2JbDuOixxLZLf7YaBtvUPrV43iT+Us2ECVse/KQa9FOSJfD6KRHqzW/obYptk
ie7L5f8IgRWRV54cPOK+0RWr4P/bbrYEiuckn8H/YR3WZwDY4acxV5cUehF4xGVw
lL98xDZW8sPt9wEr8CesSXz9KKyNaUio6wvWRQhZlL7syvyH1x1K/6ERj9QRbyAP
Q8vPwzIDnk1FqSZj5cxjcF8knQm2Oh467llTHADLazwOhnq62xg4WbcrpfFMfuYe
oLgIckZTz4e9Q9RPNLxyzaxMYNcgJUnJBIX96dFsDFezKkRUdXfWC0lsOqb8qeWS
cF5UsH+i7+3fskYjmJFUKrNrLBkG0pIwQRTq63Y/6lqIY1SBwX10aK7swZU5pdK8
bDkePUVhnvyw/OuNCJG7cnkdT/WZeH/q+9yVaa5u8KBNugBIFB2lCdNGBdxRng5O
XKBIwCpfYhLo5hmffgeENbRGYuKJgMJrceOf0cjLLfbNlMv0EFjmKQpfQQSggoAu
6ZP56XWEt1EJ32AHLFM6tolsR7RFJUo+wui6JdvO/w6rrgp6F/47BOJtP7Vc7xBe
x1PGjLm5KL+dl6fZ0jb5lcnC4JYS3Bx8qCNhVvvp09G2fAUjXy+tzGm6ZXm+L0ld
9yKGsGiv9cNsOYBggPtAYk8wnuV4+DSGT8g6TcI0YqQwT+XaROgE4pGaTl7qJgcX
Kzf8Nc+h3x24meKg3LDj26hZEtUlNtZ8eEc/rVZSFXHD4w7mQ+9C3x+JIhNaP7tm
sIOVNIIouQUivrIZFBQOVLA9TTYBJUIYGPoJnyYatYBi01kvwF8a6Clhaj5zAo8A
7Zgc0EgYLSHokPJzszrz9DXyhbh75kIZJB4ZJRV2MMeUdJ1dr8d7bLLVkJfWsO7X
7rQ0WCIB52HrhYvnWciF9ZnLoClZcnEbISHaEwqA/8WYkTIOq2HXoxPMwt8IUxtQ
wleraKh8eFZZIB3EPDC+cPCtt0f3WzHv2ZENKOrsahs+Yr5ctLdAlEcYODTIwMmE
+nLEaZW9emve3MTRzAcNWxNyi+Oe1lpcI8EMChoqh1wnTgU8LSlAGJ8Fz5WW33Go
RUKOXd1M7cwfcsZjOE3wbIGI/YxzRmYaAreN6HIuW70TKXYJHQfRuMFCGdfEk02U
a65G8h6LKv+11ItodR+dRuygNf7b8MLouZkjBeSvwak+L1iviwzUV8h0x6oMbg7Q
W0lEF9pdSTBA2ocUpTCuzVWvJlbMb13Nc+qIJHvTYEE43NXXNTLyV/TMJCHUr2FR
wagi17kc6OIteaBgyplnenhEj0jo21M451G6gntnBxxpGPgjwpSqaQ1wnVcPcB4o
I99PuAIyDdnedixfdLvFPFy2WwIlrFfHEXHS4bsBQnu5g+nCEzIoOL1j0TiygPyd
9HusVYhwgxyu4LAzyiNCg7w/lguFyrTzwo92WxLT39K/vNAPjz3X0H2mktkn0reV
a758YLPNaVvzsjUWF99qonQFOora4+26W0PPDeyl4xqVSCrsVoj26m7M8hKwfUxr
Gbv+Zx1ROOrBmrcRoml7XTw+LsHCuT2X6UHvAxY+p86RDPWjAbbWMKHSuzGDJBtP
l/ChVBnk/0d5FaURvXibFIztjzr8tjiqU/n4i4iwKpepRNqPUPG+kTOz5+80fp+A
4fqeF3EElEfsUm3HM25m9jxggya+5AbcnNw3lkkIInXrkOfdLP2Jfoaj+ywbORXD
pQCi6WrvnUunZbedx/ZQS2DtbltHs5sgie9SRfW/R2j2UVtjZs6+1ExThOW5EHia
FqDPIeSsSSIIDDxKbEMMXYnJWHFboHSMmCh0pOm87Ln0NyoasMfLNA4q88+q5rUu
ltVSJy1sN3ww1GtTeMr+4gduyOuk6dZVuapMdDECa3tNwvUMvuLs4kM6sCFn5JZv
4Y6Y2QdZh4D+mdEejCEqCXsqaStLXsVGXg0AxvI9QN8LhVagdQTSSLauOyux0ECd
68Kw7O/LBUbfLPRyuLzK9nfw8tseKSWwVv3FVOvysHdlyaC2kvcuyysrEwfiFpfS
1u40JqjQ9sI5llD+6n5QNjTgaKUO15RGnPzPg9WIB4+0+pwIQ8G1TRIZqokfujNo
b74uykXDNTWbAc0nk7xOqzVFENKeGn0FKk3nGDtH33irVotXbHbOS/LWpmzrulne
VXjmlWVCppObXNc5dqXaKlxUPWDAgTyscGMrEBUx7+wwXMkcJiQe60NMFx9G79Cm
o8jcQOepcEryyxzRYgU7AoAuMZ7lxeF7SlKpK+Tj7K59PFW9ez5Jc86X1fqbjPW7
6yibc7wYfgmEfOEJtoocBP6q+Y39qE5jr6vXNRA8Rz1sUhSQUaM4b7Z7zYpPvgBp
hUJ/WXnbng5mW0UMhyDA04779YJQG8DhcFubU7i7LRs7NxbGPpSOaDGf9y/AVzsw
wQtdXvCOccJD5UPiCurSokXPGIKLPbOv+Iapb3Z9RZK3SbNmD5unGBnphMcLIEkQ
f09ijfCp8R6uufSJPEDVbuTTIjmZmPx0IQ0Zawv0kJz1qQwFVGb9kyXLJyBiu2lr
RLU7XkN8CSDG950S0h3o9VHCv2X/2DJ2Szo0DYoLfbTNxkh5vHJJ91iWotqrq85p
UWRQk8cqcyKuSda3VfoeE4Nq9E+NYucnKUvclHLjCTDSbrXUYc7cL4WGu/4trGj8
2mVDgU3GhKr3oPztz78jL1IOSxSoVgIUEOd4DW7PztR1/FDM21aFBbL5SY7HDJOc
3ZQ59a4DijElae/JZx9ZfJv594mBah2BHpAkaRkrjrrq8xVVMQSduRZUMr37ssBd
p1q38x8eewYV//kaAbO8fqjDgCKGdGjKbES7Q/mlAtKRFagZRMEMiupqeKsHmU8+
/SG/2ggzLAU8WQeb4+abcaeuyjLl9JsTDu2nXuTpDJgRHnJY4wmuVHuTC1yQK+hH
iuNJu7wLsuwDRdFnPrXDfCgzxnE5l69nK+sxVCILQZZVWOwDoT9DQjbEIGgrgnKn
7qG79hOLCxwDfHYDi1JM/2Bw5A63MpJ1F/crgvXcpn5PbYYFypiSVO0wNyukoKiN
gqZIiDKDvOdo0PVme//lrKcyojImyfSfh27suobkFiWUr7d6ND0AYhYTNIaMXuWI
bamMPmwxkt9fbfmvjYwnJDPfKecPujOFKNt1EbTUavgckEJJlsflu/Se9rg7wPLO
wihTbaEz7Rh7+PLrf/oR8v6nqxWyspJn4bz3opmYHFPzjFi/8+7Z5ob+3yz2KzYs
Ur/Vda+JRlIoYq4tgeP9olForQEFRe1cZ35tZ/8mJzSo0QLenWkgUeXLJkMQX9Bt
LN4osu9FhEinUyoj3+iPLqpou1P8HkOsvByPjeF9jycIqooWXEagQcBkUBHzA63V
6BiLivB72TPYTYPJa+YgLIf1ESmzp7NxZYy/cH4c9KtVtBBqc3xoN/5fSNNueEYl
we/ukJVV9kJkry5iEzgwFop/g9u0ymXLo6sW1SEZhPslIEd0MeV84ETnjndSdCQb
9awoXvdgFSKYwU0BzxX5jIC+vDKYZpLjfKkt9zrS9mGY0H+CJnv03axT9LtCedBP
KQyHmb2TpaKjRe8d2E7YsSoUM7rvuBg8+4406Wy+XBRV96I10t0qkbWrcL4nW1y+
8RO/FrQVCMlIVbtoCY7LSbmZ0PE745XwXi9adf8R7yVueGdr240FSzPpw98NJD8Y
iVPoHy3hewIyYYXwwtq4QXGwmOr2qJpACjGx4b/9EuItgB06wOp+CBv0dQrQ2d2R
15fwH0w3rVmsMFNOHTyudSxyfY0nhz2K0FCCH2trSHS9RdfaX9ER008VcdDBu+3I
3LawOU2dUr1IE/2emw8hsJDGys1/vuqqQL4eDyaTL+crqofBqX0mGRNiDlOEaMh5
ChXcURBBooABx7tA+CnqWuEsFGel07qB7M1NfH1a2c4WFkjuJx8MzI+JHVGqRkQN
iwwLah8rPFhkATRaYobq8gi6k5DKi7F7S6PceE74pZrTzf319F/Z3r8JwkJpIKz3
aRM3wtRa8vu6D7MWcpMjfQaSmM/QIVQaZUMi8biGQq2PvyNPYCn8g3LmoRCyDhcl
ccfHIzm6d97Cr1f1xhoum7OIC7xnZCyI8U7ubyXt/6Es3eGjnjXPwmAQ83k0a94h
Way+jZfGQhB12MAiSGXX93DajTZ1jJM6DcxHCy0VuMoqqLxtxhryNC+AKxP4fE2b
QojCtyMcpR4YURIlhJ8yfR0ePwTrk1v0NR929L4R6JdVWBkrTKEMg9bXw9BMF4bx
8JxRuUixOFBzCudTetgTTwMZPXPnHMrUQEa/Jd7NbgLhhdYLkY+O8DT/j1Sa1LU7
xY9m7YtUUlcIm2Sz+O4oxR1t2Qs307uwCzm4q+W6njnyB+JuqT5p/SbECTXjmAWk
kxuSls35xNZ+lZAhFqyf1bqKfwGUbhbRYz29PkuXaYMT3rgSlX6ccECvVM7LU4Nq
4zj+T7RoE5SoT/CSAEgNX0uu+yhnFxWrL3pveCOZtOfh/1d1QoWWhIEGaxDatA7E
xawFb/vlNnWzVWm3J+ZJCgyUcwhbuxj6loL7Fq32INaMJ8C+j8ucOn3Gy6OsupKZ
AF915hueZgjsrBdoOHm+mgG27Rx6fWMMOGD0jgaV+38OgdWDpcfwRTR+/ZVMMuDC
XbkyVBb1MMcC9WgkPMMtBQB60wrZu3dnhk9Fcra/6AAmUNB9WTPXHHW9bquC7kaV
2XiQe5DC95lINTGX3pXmrx6v5SKcyKZZ6EWz3Pdmxe5u0D7dZSfov6Htq26V8uKz
XVc8iwXynMTLtE39vsflKTXaQxf5Dku2s5Xac/Flf7VuGi3HmX7gmVENnNkBHiRN
kFQATEzbupAOwhEGxOycDwOhOptsZmP+TyVT0KHW4QJQIYo90mvUqJHOl9zC6HOH
KbYObhLxLazxrahVnTvjHwmZDVKJH7Lnvq5WvQzcO3/BDAtNQxmWGDXKn/P8jF/j
12a6eb+vt1sUw5tWK/E3Ox+LF9X4izODqEtGqEKhH5lWl+YtPnHut0r1WS2w1bb+
0YL6c19kEZIkvcnEZpUO1hosnBVxDV7GxAXgycw30fOXr9QdfcHLIlVGbPgszNsq
PwPEN1r0bs1hUkkGKUmjbJWeBe4R7WSCa9nsFq9ecBkklqY3n0Q05BkNOyVu/IUN
lO0CUalznXdNmVy4BlW1CKZv7At7offlOPCAm3qc7Pg33Fliiqw+bnQaq5f0PdpK
nF9dzCjw8mMn7ijATtLxS0R08+MwduYL+4Yonl3SASxzF8n9eKFxdvSXkessJJdB
AbzO3dO6OAJTbx32JAjB0S1k2hzNOxZ4LiSe50eykiAKFHMN/OgOKxp02XtODCIY
llLwNTpNpDi5yvUUzLPNRi4dANsOgL8zrFx7OVLvr++85/f0A4K8EYAhc1maabkE
ZPgEOWJ/sE1GrFy7S4cIUwtqa7dZ8UEKI5NejOd6Q4K9pQQn25NAtes1LZouwqgC
9HCuqP9LXehX4YVdkOD0Wfu727v1JjAw0WDhXzu7tFcvDHoKmvhmS6BNx0tfRowL
WrEnv0WNFhUmBrTSj4ll/gX5RSQ+SofsWoum1kXgGhl4Dk2KZRtb9L9Mmls+rRaG
xgyMImVBoTQ/g6oGVRhagVm7XocgEoSGEia4vL1AJQIjRV6VbJSTedH+/i4EbBl4
j+1SteVhAShqW6ltDPy0Gc0hFeQr6n6OkvJvmioqo3V2rPDWH2lWCs29fNteZvaI
yV0O5rXW2BDLKBfuWsugTGEZwuegQHbPTYDnghROGJc/tgQ4ZyTk8PwtTt+kqW0v
mSMUONuQmyOh8AOu4miqaNS5k9mlryBHjp1O0Inw3650OPMhTuDZrNpK8KEubdXQ
tD3pj5j2llLAgCEZP9S0FsjE1Ibbr+URRM3ZsIP9+GD+hm0dbA8kBLFL6KLyIAhy
6JJ8ph33qGr12sj/tDhso+tQmHQnuYkD1mkeCBa4FBZsPxYz3FVX8rVS40wii5X2
NHC6EOr5LQlBy44xcs/QTnbKdukyg4h4FU0f8raT7MINiY3Fl+sb9QSB3ULcwkS/
lq6SQ80aiPqo5CbaG73MA+mOah1b1ztEvl6ftFvYRy+YUXPjNSxyWQ+R3FK7R9k/
C1pkm/NNDnMMpi+W8YE4YEh6fN5FM9gTod59gjK+GQVv02pCY+SworQByMoFS2MX
a/0TRPpmQ7cMvzeqHYq8IGIv3Dl8Ia1rQuDwBxu4UPmLkhizp9mFTlwjOSMK3rOA
l/xF/hKM9X/Pc8FX6tug/JNPjYV6kNRP5GW8oYB1DBf1e/kvL4Aq070MnWlFXw99
BWJM7DitSiBF/gCHvnAiDNKMiKiHZa7kBP30KR+KpNYqfBaqzgepxgRdtI1n6mrN
8WrfrHP5hHd3g30HvGe/9ADPozudqH2OLhfD+FRMxnFP+TUaiTpLnLDOXLyR7diD
e5FHEY/sUO35RH6VSkq44lcLoaAjSFEqpMlpO05lgH38rUHtbHk+u7eXQzAZp0yv
w2i7OTlPaRrQCAysWhsQTSr4k6EHmStsD4xHO2jadi1kgu2NqWaiX9cxCOAChUoM
q6b4PaBBzu0iK1ImpdwtHilHWCy9bUtGiROGKQ1dOvHXHP5sm1h+lZfLrdm6xA+I
cmzsEGFUsp5v2HqY7SCKezOW3XDjUKpPXQi8mZLN5ToER6vZ4z+7JzaCtL1S6E3c
CRcVngLxuKnLHek1SEvzdqat5EV9/XvDWkUW/5SRcBUyAEutmRn30daFocpWFeNO
MGTZijrZn0ysO/RKA6Sc2B4IerTcJLPHH1Bs5Kp9x93wvz2Fhu8NM4avK+nNQwuq
dSMMARo9mJApejLpd8QSEDvtOL+ys2bIPs7srpFbBhYrDtdaqBuEAe8vlf3D4wBe
Q1Pyn1vnKrkapHMosrFXwn4YrluRvHSsyffcl8k+lCXDFIXLk2CPiJvIiThExGtg
Vp6SenhnJ0jZk00sakBiBLEQcCBPDoIyrcpwZmNncqCwHGAhemJWqLp8jenG0sK3
Yr3dB7cSulv++KTe6PMCHbmhhb89rPV+ZFq2SqYbEiDarrl/hFOrRhzEFxxSlhmD
AS9rhzAItNEFj9zPVE954p9wEstH5e53WhO+NsZCUmeHUgYRYwiJ8UbTiERhehnM
LcH2aVyEJsmXyv3qjZkQJkaah2Nm/TTF1urntz20szxIdWCh7k9vLRuH6YK5LLym
p8b8z0qP3TfUDuYKWyxyPNaIfD8ElvCSb42TF5vWRFFiYvs205GVWbwWlSAirt41
5P/cfTMoNND8W+yUfs79TSbA1flazvw9xt9AhQg8o5ecmlz0RID5lBinwhm6LdAr
tlaH4sP3NXiVJGPh80ixVbXKC99xIjdAoumrmYU5u+59UnueMIO25bWmz4nlOzZ8
mtqCYJ22lx0eo03rh67UBlsONE0mIBHSZjjMMTaOGw4GEUL6VQqHOBLSN8wiOueG
rs4E/3YSws3+jTH8VFGnW5IF0SXtq5ceev4LD+3ogXE1f/KTtQRztfvS9IGLCH8h
78Gymuv1K6pZRFNdzs4qkZmfUhqkhnRRZSjxfHETP6XcjCmMvF6OiiRdCAL4pcxo
rxdbnhAlDDkHBOb4L7n6SkHXlk0D9mZKYPyRsqB4GJmaXfKFxcKUoRSR4HiC7qx0
PUn7NTWoK40U/3jyXV9lDDhYjdaFpkFyJ+R+aDZ8036d6IB0E4W2vCyFSP9IWfLU
kC/jY2V9WD6GnqbeS68WD/QldcnsYR6aqVTKhbAfr5iYwBATiBYdCgaHVRqvKz96
e/OXyAxh82p5itDquAfNSYMoHpxUY04ZrxENt4Ca+Ul+iaNIKmdK07Q1mA0wQrFH
zJpAqmU/0NZuB8uIcDL+LPcyMyeB12wDJGm1IWTNpnQ3YA0WK4lI41WjVhXaAtOh
VvDPPtxlNvWnkOy9ZX5MPy9sC6XhEdSDSSNJA4jnzaBQ6tYqfZFt+p8VaVdF5Dst
2XDGdv5uV+yrZnsgjN/eLPg7Wdipsyt8qWiHt74PPSye1Vs/jNQz6xlvi0tnw5s0
VdbcAxe5BWIW7CCGHZSCLU6qIILvPwGGEcwsugA7XjIyej1UDD/p22twunYfmhYs
sH95DuxYDusmAmVgCPSa/BZTFK7pgaaSb+KwID89HRqqG3eIP1emgzd61Boy7eT4
PuM4321lCSasKl12foxswdpTsaHpaOzkBXGttdewbBWcj7mjXeAbS1G/LIudsB6i
V1Gv8XKPFPdwMD0DJK+ud5X0OjM27ZXjXayRJabbSWb5lTw6uYQvW5/IcJmPQoGN
eqbEbD3bhCLYc6EP4aJFA8599HcwifnuCm075iz7pIAIoqmzj3DPeXgVny1AIH7Q
XIB3cb7CLnsNaqsIKthTn+ld7uBKsC5MzebYKpb72db8xXUoKYgQmsPLfaz0gXSg
B3I2OXFoXKceYmMzKLZiEQ==
`pragma protect end_protected
