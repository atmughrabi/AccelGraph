// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
s3h42SHXHG7NnxuDH69s/bPhyxB1Unz707E5MeoPyh06tIb7je4qGXyrXg1D+fTl
XVmwc7q8QzJbyeAnrOC9sniYQPfIXxHFt1WffLGbuA/KhLluH+YU1E0EdRnyaX7z
dGma+S+yp0OrWVSRpK6OCuaFj2w9l3jZ/wYMNebG9uI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29456)
a2QHYqynIyotez72t0ox4NKfSGC+aRc5tmsfAQwil6f/nZQQCPFTMN7XtaX83jH3
HBOQt0GbyT2Tgg3fguAw+rIkca+36IpZDQyqAE6IS50tm0c/vn/ZOpAIw4JYrTnB
VjEyntai3geC9wKXssPtubCcQy26Z8sh7sRQ7UMZk3gAf4b/dDhp/fj/60NnPP6f
7okmlrJhUqY6GpWN/IFutHoSEFrbT1VV4+36rzK01UZj6TK6ICRd6iKsYOP1rRSv
7gF44WTtFQEELhE2VQL2XlfDTgQb01FD53mpf2UxnQtOmbapHlzUOcJ9ceZu+fjA
c0SosHQTmMSMNoDhKms/jW3mymS498evbQghb873RUjLCje4bUCGjkN7cH9A8MMT
9xVeGcdCqZ0yraaXbI8goD8kAMh8xFMvAj2P0OSlhjDHJpV3W9uEP2U++ZfA2CEA
NMEUBuDE1VPDbUiruK6AAahlqIdLHMc8Ou0Gsk9h020VWzhVn472tI6e2OO7YkJn
r11OPbzSleT17pNjqpiX87tGl3wfSGQzVz0wH2Qjcdf1fIsJ7Mzc5as+vCV2V2Ou
KfF1AO5mlmfBS2z79x0RiVSTeuWxu3PcyfKxpqcsNFr4xgpsWW/2vks/m3tYX/Jq
svyoggMs8Cj8qKNDROtXVOzOb+SZ2WqAMw0NixJ8iDjUDsRNUp53DRChV+taxXLx
kjsNhzPjiSJTTGekwIXxiKLRcBFY5Qm0WEtwXZKFCrchiI7i7RVO8RQTdPPnqgZl
IZ6kMjZa3Ld7Q7BgCJE+srC+Z1iLgntSVQLosG/n9olmfRgT/9qSGeHRUBUaJEll
tSJjBmOHMSg/IXY4nAWbRWo6x/hSmNYoeZSL4nADna8wOJkACGRUGa4MS/meZQVU
5FF8M3NjrxxFL2vV0v52ue7uLadLqyGajQuMnBlBY7TIsjOysUwiVGAJNvjgCn5n
MWQTm8u6LvBV3zh/lit/mJ4oBV6WDUgLjNeAl6GuoxkSe4ukyyygFqNnT8BvvfsP
tpDgD61SrJEvNitJke94SPgZ8iplMfk3f1KE9Gb7OdqYXyIU1Nu7fvkIqiXMwzte
UWYpplXAPfahPvgm6aklWkHJJgmcYZn87c4AFv7PEWTieQQWUC2RmlDivWgmhqal
IdgpQT8BFbwKdOZcLpuBOn9d9cKjQAbdE0r87jwkvnIzPZQBOwnKFbOtGwhLEl36
mKEA9FBnHOd0w8zhuvHzFfCTfixZM9HRL/XhV4zKYieS7bpL0uJeapwjUY3s+pL7
EyfXrZoKkUGdmBKpzDuaLx0pYl4O2b/UVNXhC8g95Cib1nX9CqWnJF1wEMpAK5Vm
t1cdM5Z2hhEeuKrXhLy0RCN83av3gV4lRmpinaoUedwRAc7xovIkbBWlJMsJgnx9
S49xF8BcfPKMKuZ5gvrx3efZ9vSD6jysYZVSgPgE/14i/0Mg8VQmAJAp1bhzPVoW
8Qu8p9pBXoJyAg17yBRzNTtLQQvuMRDuc6UuM5CZAIFKWQTS//c06O/VgUgnHgVu
Pg7tce3SW17K1pCcEHB7728TOJj0wzsuXO6WcjNDrl8gZr+7MugQvtOoSq1MygEM
lEJnjgcGR8eIrUxkAB++ZTpQ9q5zd3ez0q7Ob/stLSaqZDc8Ol0Y3vV4QGdtHEom
lyyMKnMxWiB+LIw+UZPz6L9sSSAt4p0FVEJy/53TKFE+ZMQPmS9GrXalpDJmV4w3
4QkZIAGE0w6ge04Mxvz/BLvRvEaZhsMViblKARm+K/cj2yooQQji02is2/56dNnI
gGLkGHNln6wlvKGqqxqIjcWXb1Hp/61Dhj15vrFyj/GsMgMR2Z8Gn13ZcsXaNR+h
Pym2fJ7/0c4S7Dj6saHFXGh16kscMBoCwkpx3Q6ULM2t84eQm+kEsz5KXyEQH25A
dvV8CSaIuJDaJf1RoTfoYY5smrfR18FVGVpgtGs5SEOTH/xqLNKAxtQAsMtSNJvO
4q1BzLpYxPexabDN6/YuuBufd1PwhAo1ek+wjECtVVdPfFz6M4pin3p4niP+sqGm
8hA8EnJDgoVmuZc/hJKtpveXVvX9FjhctuvNr1BTF7G/REky1+Y93XjxxERhRqCq
Gq6+VoFs1ZdbnAHXvqDVPDQS3miYMpk6aeCqGcmNHL2a3rfUM79Fp3uDwBh86QuM
bUPXL+SASDRsrEkSNtzIIvwVIVl30a3oMxbPdnkAJKx0u3vBc17lRS5gYtghOcW4
bXOV3pkSgW5XQ4RFOdAMm1sVvFuCRMWSNqj5TgSQkrsPloSqkSjg1XhNAEXgjDUG
f0b9LJ7hWUfWeVS6d+0J5OIynVFwpWER60Mg65mXIVZV67H9MWdkNdDarWaafRlo
nFkcd6WuN/OILZVh7q2VApmBhbVcHF5d//L1zekFmjRQFpxLTWicm7H1Z3zAKZPl
PzX82t61OS1arlGL8sD96AIz9j0nRbHT4dgN4HlEgPr8ZB8vIWVv+qV7hI66KVKq
u/iMlwoMJsr/TUYAmjiqFbURoa931U1tpeWnlXBYiGpbJ3XNH4J4fevVGqB9YxpZ
3CZDI4bh774H505GZ/w5ZimLNyT8Y3iWPJny9bOT3P2iStI6nFl59UJhBHUdkRvn
fhQRksWuEK0lOcDu+/zG/nOgbXcAiQaa19dpiYOZlEYsR3+ciGT/iAkzs+d+IoYq
xdF3CV96eRgOpRF4X6DszsaufVKsDTFMlLvIaR7ZKhclzVyOlOPsmEfFOyTXTujy
pPISd1D9WKYjf0EI0jML8A2qWefAcF8SXIE/ef9w1FzTz0zqcm1VCJ8rH2bc8GbD
hmF0iuM9K3DcWmzzVmSyYcVMyzcSgXw37X3E0UTv2mWc1k28ufUMq6n4M+7QES4H
p9Tnt3gH518TEZYnBoS+ovkRjAxLOgd5Q+1ies1FfMQtSgiDW8hMqltPY/Uj2LPj
1czDjqfwv93IYiepA+qerfCNCPrHji8dXb1/MchBGzF0FgMu0C3Zi9q7x0Hstm/i
8tGiZEzCJiFNB9dwtO1fgyQYzHH0rLJbvK6xvyZmd3x8osiWTacDQWJNQoCcCRjD
/pvqlBuu91l6NuoWzF4aSQ2QdcoEwbqJD0+ez1sz/OwRxTb7G86X9oLJF1N89pWM
CXlPvZAIS2Yp7iIgaoCHgoGEwUDpaz8tc3xTTc3czkeyokinPRLtj0dX252piT0S
vZHheVGMg4E6dGvbHAiQ/8E7doL58kPxwm3Slh5yW+gQxHcvrOc/GAukN/a69Y6i
QtmAoHR3Un/Gi9anwNEAjEUjmadZwq+0CW12xdL6t175GNeZDTkeX881A7qqaZpP
7xpVtImhUbuWz1c/u88jzoumIjgruqso425L3NxGscmB4R0EuZtVqZlEHokuo4iU
Pv50ozotyHn/m64Ysur2gqsg9Hcx4qrgI0/dRucaPrRlDRKAe51GDvnSdzdd7k6v
a8xAsEozBQw5f1quIh+h3U/beniG74et602rMEnidg8cJJvI5ImWILbxxx9FJ035
TpJKTsliuC4gPMM/48J8y1nQU4hJH8DcKMO6V4o1D5beKn0a3eu6L8TV60yAFYRX
yi1f6fNVLHuhdS2KWLGmVHI5wHEgCQTuyvWDqkbKP5VTYMk1rH9HKcWDw4D2jwrh
32OLmu9vQMdKJOKXUnHcKG4boq9CIXvStmIlNXn7oL1r3TwMx520kCR+9WReJXTf
uldutZCTASL5JB19Ybmy2j3pLCmG4L3vFp0hNLJHeAXSE9vHM8ZBczhNfk1IID98
56xf+SNWuZEaupcLxREizbdVVBAsCDA8RK54CYIhlFVzBcF0a/w2NcVfRo/oseiY
B/Tg5cYzPyFA1uSOIsJZ7Kxv819keJXHrL8C/aQLFctwR/XOobXKVeMONBPejMfB
ohseOnaCm3a5zZmJ4+MELl4TF3ESr+Vsgysy44rVIdeqZRTTsTDqWDErs2nvSpoA
XBF7nWb6YlVHipjova8ilGKfltkCImCl38PNmGuEj97Y8sxcazQoSgJEm9pqZFNZ
cmrlmxOSUFQiZWrH+2/bJiJadu437IHJhWnlzjGSJo7+bRoLsNJGBsl5Luq/hrUJ
N3Ygxex5dCrl1xbqd0yEcwhM5WUe5q1S9szE9uFxwTEZNFms+cCKMeduAhoxTxtF
1eN/2HIaOhGUX7lXmVmFM4W+XPE0Yp3MtDO7k35iOQ3d3Pp9sL5T4E07tjbNkPIO
N05yvFANiBGTDofVrofArmZPsEI0rdjK/2lrubW+/VYrgatryte+Zbuo9BSAJ0+l
mgsIQsQzludPz6zH9E8DvL2YaIrE5zRU+Ykn8Wol5rmMqORAJKReTVPHio/DwYk6
gI/bMG9z7XW7ER+JDiDFzecBgXJHJm9njtmQpLXlZT/kez2aL+XeAH+RmxtM05PL
fE8vSBxdj8pBsI2OazqvlBVdf26lkt8XU9o8fFjWsVb0UjUocfqmkrW7KIJTAnlh
D3cRwzYGwraZX6JA8YxtwHslRLljE6Vn2kjDVOlkRRlVOLneCeiGIC7F7+94JS6F
YCTEAEblf9o1v9xJ4xlgzQyrezxOfSryS85gZCW6SsEiFy6fwYKItDD5n+8+/T32
JWfoyySpbUn5BijVnWzcghuKI+Ik+4kZ7wxAHcvvVKFc2e5wZeHso/PwFaWVFAcp
rz2/FYu1x4l87dIP2eShjUbv+wwV+Btq63lREa1ocTTDceQSJXg4V+Ct/VwR3mV9
0c3JeRsvlehAEGfjjQIK3HcR9t+dja4L7cFEHsdEJDV63vagdteJ4ZKm0KIVMz0u
T1BVcTXam5uBcu91hCLn/5UABOlbcEP8ecIirXMyFlI5drBOHDxOXkqf/k9xFUDR
lwKur6mHCEiZasCiVSkmx37gNWHHLInpf9UyxuAGczif9q7ANzXqWqBnm79BW1cv
gfir0BoXootvb46kS8xcwiq/QFe2j8aYTXyG7nGdzk/RdbEUPJd2UsNsPNuF4YhQ
FdwDkvo0MIl03wAGj6tpYzAbH8LUr0Bc8cA935DcLJCxeLbPk+hl1UpShbaAkevP
IL9wiPvSt2TM9uLnvvY5ZVEfLs60c7hMmysODU45MiNs9Ks6J7GuicCuznr/NUJ9
9lD2fBF0iL3BxkPJxcYBcBMKnNaYldiApn7whQpy39whlCDPhj3iWy9e2Jc76d44
T6R9Zs+rUnHmRW+Y88Ak5Ti/YoSddlEBW+U4wL5beqKVSqYSdOZlWAfnizSo+n0s
1Ve7Yiw6qwsCb+YQSPsS2B64jBdR4oWOHHIqJN2/pB+sRWvZA0yCtFrCee3nq1ld
R5DvmF1hKthDdWkfiJwoD4WylzPjkLvOpUuYvSDLql3mxxLlS+uca2DAMhqfs0I4
/OrxwY9Xqs2ljvzW15GE8We88K3+ezFFe86rS1rNHjlFcEEm8JUcdH/9CEpkC/Cs
oZAdYciWAjUS8Dp6PjCZFsO8Y1BVfLBfSR/4VJTCFNR0a7H4UqDD/ciJqxtnvvnC
/EcSZtjsHK/lpG0Xdjxy4JINaWid4e1XI0uhc4qUZ+hRvjdpZ+yP54tXsNb4TCOF
10kGUUuaUEAtcUGXn8mmSopVhidC0ruJ8SrzOCQJ/0tBrVezgNumEg8NK7+Pk3V0
1w8hxut0C5uxteKrbqF2DyMrRUrDvuZEe1KnGTRFjpAFOc8vblG2C3r6qRPGa98L
5e3eGiBKcUP4Rl7NkvvWip9kBVLcAx7oznUMP3Dbj45gI/b0zVYlgVwQacEqD8Ss
Eiwf50NU72RkiSngRG6ub+CbOvF8LALTBFxDjinhlpzRNFPPkmFo1eRkz0SrmDUd
MtX6esJ0hMYSLvQAxa/9LloI2dl29nQz2DyW9UBbXLy6rSk04TYg1owc6DToS23s
R2s/Icaq4zU/iI512wbdr9WB9Fj0ApxMKZBgd9HMtv5hQ3GzYNWWvQ4NdIxMW+pg
1ndSuwXGq0h3mnbmqqc16xYI0xvHi0z+IVbGR7Z7g7ILY/EPtwEcrMBaeifj7Dmo
vkJ3U4k80oowwQ/cydYP4gI/bxVda2Rh5A4GKN7bLWLbs6YWdVc1A48uZKaWf0QN
feiIlhB89SnMXeYpZ2rTziGrCb4QXeHWxKmb7xOwCV++A6yC1DGdjLMKnMSUJmGI
tJlEQYh24fls1s1Kl9mv/z+HhakY48q0at5HnkofjxSSNgWapQci6fxXcxeXhxZZ
UgJ2HbPPcVJn9vsMOdLcvojgmpUcQ4Ndp0Zf2uSZr1XECJ9c1xYFBtXQN/ExJ5j9
0M1j6x693uf6GldTJHD8cC68IseiZWEa/VZer48C5urXYIVmC9LwxrSqyE3CWWzL
wsFcMHVcUMyOoc0cZsOic6WE7elL4hOtDtexE+IuHcAgDVJnAIKguwcpUMXqsh3Q
JCaiujRd5DqFUKqpe0u+ESXp33FmelWuewqOJQFj9Tb5p+cS52aCVF8aIrwUlr1d
1HDzU4Ll87rhukUCsqAjNnqsRtuOCM61iz6uYjf/9WX+yWqr+LtzCb96c8pvuPrk
ncY3uSex6EW363uiNY0tpPoZ18ZwWu/NQTRB1ezkcX9IyCN1coJSJFmar2pw0dYQ
U+tDTHKU4lZBNs+JLAEx/tujrWJ3AsjYrUF6czsxHIKU3erqJxG3kvciRmEY/ekB
4qkghLoRszwBRZcJj1o0WOtv0ztb/FB2afYscX+khKf9CkO1t/PlELr+ALL55eyr
J6YhVhxQC1rAitkVKdldV3HVqCYFWxaAKOehI2TnO2UYeNJiRNWDojm0C+0DBgjo
u31lzPh0bBEBWtgQngAgo8YoEEAjWKvikU555QwzXAjD1pRNAXrrJUcY2yhPmObk
SH8Y9hdNWPMGkxD/OCaNy87OaK5qyBUQaJHCvp1rlviWztGbN1XdnmOycadUB3ip
kHN2SPOwRHA4A3DyqrkPZTaFWYw64uSNuI3r9JCM6bN0QsFqFVOPYb8nrVF8lQy/
zslSodl1CRAiwQbWblkiGUQMPeZy6sImmHKXK9wpHxbNRvyVgQPoYkxvddWB7aXW
+F2mHXxIXyPMcxfQanLjdX/ZfM+HsSTu0tnfoegDJMYVo7wWRb8fNJNcJ2tNRcLv
1iAgFizZUFN14UkJWsoSTBELiAD+VNPecMq/MhtuDL4Tz/8ttVV7KZv0WbSl1gNM
WVRhLxfoiktPR/WXKliNAPJzUP4ZMqLYOIE+2tGuQ9jOf4M9n+Oi1HG7JwddY2RP
M2EoNDSIC3WlgOOmd6/kHT4RmIssxE+zvff2htgA3oL188BUcyzwR4F2w1kxIB6p
Vg1DXBkGUS1P8NqFfrtyB3xDTASJq2K6VVDewWVTiiF18NNmwFji6IV1IV/kJSeF
DwBIhR6RN7zoMvf6yUv9di+Xhu0DoIqFsT2/s4oqYNTbjT0rZymrdUqReuqksIfa
zXRrCspV1dDcVtciMtzePZOPEwtIKmouxJtdqfFbURFELOq0wUNQSRGxrBg1sgu0
czOpygzu8TRL8s5FySQgP4GqOvnQcGgDzs5sLtoWK47lbQwFxpE0eYnKsWEZOa/8
AXyWU2TnALFu65aAwZ+bkFUfMeS/Goc1VMFgyD1IjzBqIALF8skZBXaWFzZcTIOG
v7t/osNupB6Us7IrnQIvMpcWYc0vgJQnM36q/FIAwuKDIUuRd4S1IEv7clvZcq9Z
9SxUmWV179GVUBFa76haxrScsOXzFVeFRv1F8NfpxrjveLMgVp7h3/q+44+CSwez
AGG+qO34tcmX0gL9OrLmn7DjkHjRfJuVwE9uuIeoAd2zyotD+7eyDaqvRL8t+9cB
e5aEkGqWvNw7uS2y+9oCuTKYpr2ozVHM1ZqGTf+mKWkMbxji9Oz52FJT09AYhmTL
wwmSCdmVYRpMCBW6DEk8eJUHpSjx9HNK09moLUhgNNJ2DRv1IfkyS5Cb8amlc85C
H4hyq0otK71orLr47aae5npt4Z/A2QlLMj+Ax34O3civ40Iebh3oCMsoCE8G6QLV
cmNZ2nx2TYbw6K07UHEx/w+Q6U45eLS7WkuBsVfakFds5HuAyQlAFIz1liKTLDad
xKo92EcVLy0WDEyEuNG/BH8gR/9iF3ZnXSZXv/amHS/7cJ17G2HrDGXGRLoQOBEc
/Tw9yLJHoG7p7MIkEZXmb+ADlI0z2PbIN4DTe77swbo/Zd6KbMZuKeVvJBxaj6Z9
U9Wff2TdFVChraPP4WvzqX/ZgpeouO34xfXbPPxMlBaIbNKsx2Uy8MQvcDVjGZ+a
3Nm0ic3xzk41fEAYihatas6o1KXeYqqtS0wYZQk14vAWGORC3tr0MByZdWSwLJZn
Tk0heRyiRgc3ElGnFNPz22iNf/Ba6hWw7sUStLh87vY+lCywEoj6eTIRCkqL3gjJ
wb+5UeL0fKmMzTJ5J71RlWHnUyuILgb7CIa8HSi1jw/EVBPwJweht1vq+hTRqp12
TVzR/9FaEfhpaFlpkOfxSx5fr/zBZxgez/LPPfoxx5HXDBe6MoXGc1se8bWwgA9y
hGzuRGmFAl0yZgnMhrLyzzCZ0lPjmr9HH6XH9paBzoiAJ8eNvDLFOgqSSAwazZHl
zknwfFjoOE5AE6aKtjw6Ccxlx1adZ7mYIPdbHcPGu9uuAh5QwoktkCRyh2QDdkEi
Bi6xClO+DO1SZOOY8uUMUrUt3hnaB1RJ/T973VlHDMExTPF+VWIi/A3YEbw/myAy
SeBIQ2Hq5NEOhQaZ4KLZPDDgLxYWTveI5SOjA+e9ngmQYjojHZ9eF5NHqEQ/OCrD
AeAGqyLLcx+yZb1va6zUP4tWsUb1ES8LneHSA7/9nLoNeiMPr3lCv8aWZ4DBg5PE
0kcUh9pY10B4/wvTOB0qypGNXZ4k2VwpVjGfDXEMEmbN4YZxuWoTscfFSkPLVQQF
sUhfM4HPyWl2xPu1wqGpGiId1PgiXQu31PdlkgvIsm9YOjXj88mnJ8pt0gaYVoyC
yPu+mlzWJ8+RZ26X+gLhwt127n9fzedVj+ZVGYekYgkT6VD8mEXaGRWAab0/QhXM
tcMWTNWNCqrRF+ctADG+Ou63wdz+MB5gGJSVYk9/RmPFHO/Ai+DWEs24jWDWutGs
dnQq4aJpONcigdbKkDEzgC6GYXv3dpn2JxvS28xjW2s5e2q6Sh06rNkgtUthgo3Q
lJCUFfvK/F7TzZrHgiG6SJQLtDoJh4J6RtNwZSnMG2yTEQZI1AMo+m6cJwSDMMyN
TvbQhaTt5PS88829sKzUD8Pfl/P7oGaibqUbvFurEeGT4uxvrbFuRAYu/ZqC+42m
zY1RV0gd3SKa7Ce05QzFrub469Ojc17jfVZLADhOj/mua9EjKIMrrWtLDAyIEMOd
9IRMcnw0KcezstbNi87qDmgPV+tIp0czsRXpBhAsD/Kza14xTxaLyiJb0wnXu3lj
24oaj4vfV2YJfnMAek0UGBAdiBWEGEnQuaiWytuNIuaVBo6OydpOzk2JID5ghHYu
zZiScezXw/QdCNBFOFlRh2Y/aiLaE4n5Rz5uoGYoIAtYAcJ3Z0sk4vkxsJfvwQnQ
b24ye+H/Vqwhh2+NmDz7l9osbO4HFlztwUZFrP0LP3nNWP98UQP2y4yLYwp4883w
Wl4ViopKz6AF8K/Fr1IkJKCzKka4a1ZzVFwG9fveL0Roig+KIMC9ZLh8pQMqisIO
lCOBAzmyiulbPwRmT0GL+23GjVTrkDzrdWsiC9vuBR7Y5/qqkcPMzX9NT2LBeeDY
zZiG6Rt0YLJ/pK5JEkt1Vkm9P7qFLOI7u3yGHUHsoGksXMq8wktViKKzqsOYjtfK
sMTh0pKPzK2tljhDQppiNaP++S38ktthXhy8cKUjGbj6CJq3W9IOLeqeQAZAAEkC
smHIM6COyso4Akn1SAhdjvGYPgPXTpDHkjuHG4s7tvYP8otPYxP/FqqOVgCIRpWL
wvAkIG+T2f0o//097HDnlDrU/VFnybXi96COkFpmckp1y9BY7zx9p5MUYXuyFWwG
YRpI1GHtzXm8RUdrosoJbk6Tzxa0V5BIAguonezWurpV1zkM9P6dzYq9FEwsvoS/
T3kPEUraUVlE943ZULDausJYl1BmQ357AH3UYrCS1l2jCbVljL4OsElBnJ7WjWn4
s78axB1wyP2nTsaoW+lsJENVmrRQ0Oq+C8u1aq0OR63z5vqR+w2LiHAS90EQDrUp
MM4BJ6SeU0eRsHsImP5C2SXMVCca4GvsZ64I16gvufpzpNNf1PY6Zx3G9Q665LCn
RinYVsACTj+HZyy/+7ty7ggY993j8Rg8hFib18z6iIAiYDiMvSWG7R0zAw9B/Cj3
Jv0TV91dfg8899VBlweXO7I1bX1WsAeR6FhLQdi8zplUiEHd2Gl6Hv0CHPBGGK4E
F8zM1z5OkjSF9nf7sPhmvdmg1tSpgJa/nL+1L7T52MohryRGUv01uT4hmwZ2lgYH
qTMWH8QXwqRU7gPhIFNfzHjfJkB3PR5sNIOy06nS4cRMqOQKUJ8EJSUg6LfXHspN
6Y0vqj7knSeFr62ipOzUZcxxeupAL31g0omdZIH5Vr6RIg8frSqNrx4yAd0rSPeo
M+VzZy6EIy8WqLjcti5cr+ckoEQMeVBTNgdpWeWeEUZTuAqrzKbshZ96Zn3cQ/kF
W/xNQpppyX6NRmKN+miaQjQXdQ5+0i1xF2Gwm4bQS5zYimz1GBoJ1d0TLuL1R6OT
j2s8QGdLEmwn8Dcf3IloDcCGF109oBrzkUyK6pPnv45PDmgXd/twNroFrdYdcSOn
PsqtNpDa5OHYwwvwfXBXSvqlLTD10ZaKVSR56hWxKmBr290SdtDzQbG1a0Zy4tew
XYDbi6Tuao/wwMO1rZ1OHKwlMJGIDTLoF6QTJMcgPxZLfPiabNqLX+C+lipGNwnj
fwBYmH83UCMjMcDRX6/gngYBFPeCh9g3XVugvwGcg98Nz018QajLP+3BEAUpmAD4
HJxgI5S516rLcn7V1+7kEOPB87gb5GA6l4ofNf1up1z+o6qTUJhJnotwMrP7NW4l
KuIoM4kCUaQ2Mlp9TgKMiLgVyUERNh79NHlX5geiDG+SigjRReky3BwcuVZIoCS8
r5yyWN0Uv3Q88PseDxovEIN+nzo28stgHRVmXrgYNCgyjChDkfGPhwXphrbiflnO
B9xbtPtRTwQJPOTrpBEjXGvibfIN7rcFGPEgQ2Eo1DFIM20OGtY+cz5Zjmcl/04v
6LE1LipD/hFm9OYxCN84WPDkmLG91QnJwWEk80OcAAEUi7N3h7cYtUPhb/q3CuG8
WB3A/motvxNiaVQe5oyg+GOdHB2liAqLOu3JN+nP6pmzk5aiT8+ghhjYxluqxVoj
pKqbNEc9y2inIbz4PC/oDsz+2VhqtQ+yuMUNfAYEuujkAOZ6X54Xz0Vz28vvk0kH
7CyEcwOExZVc6cZ61Cc1UOpYcJSF0yxyVIbTVqbKYLtRM5L2dXYpgPyDpfoVnrSk
xxxtU+prQ/OvXmjf66yPE1C24bEtifvhwbfoLLQ0wNjn3wR3LKW5s7si6/0/l5hV
BEtlS2E3/c98zEIS0kM5LAsqlJBdVckBf5TIgPkfbv0ld0rF+QrKlVlp1SHE1I7Y
FSxj0AsgzKhpn9H3S/LMqYxSw9v+g9WrZUCKk2Zh6X90dRinR/axAi+2nO4zlgnT
qDX2IyVku/eNdUwFviLJn+GGFQW/iwrYgHo2zXrNbcGOySNAr8D+DSR80d4xBzyT
IuwBsQECogIIJpTUPdX3tpQ58jSmLLZZXEFD0+t3C5geRzgkxHlgu+Apo03GsNe0
OKtliKQ/e9Kr6EPR0kvNW5LaHDvC9Sjmq1HHl1+gUoXAreBwRr05AGUEI3qLXXoC
BQSupq8WXLnfYaQ9yqGXG/Sw+CiWrp7HiHQmGOdcgZT+Jog4bemCkMg0GRaRyqpm
rl5GfsNqD7//AMwwkbC6AoumV9eOEFi+kw5aSItSXheJGs2HbvoK9C3qv9Dso1qy
Wp0hy0fvzwA6IMYJZ3NNCdfDzJ/ykk4Wj+HNDYv4HYuTz3Sr1ziTQll30l6qZyH+
4oDtoayjzU7BCSjcXNt+prxdFaF2IYxheBuZq9FysgZ4kZlGHz3ht4NwlcobHGBe
QsJ2ftx1RK32u2ji+N0DKLRMFKZprT8wal73QsWSkdbZo8LT2nkS5cX5nxfHkws7
yP1smjOVVUQguB2wj3QZfFHvRx8juqXIMcZDT9S3ip2WUHjo1jI//Knnqe2xUbrf
EFwNwwrFnLYA8Vy2jOe8GXigFXSuKnKmMaqgIWS3rY5zMQeggZ4WG6Q0r3GPSzRe
U/FtM5aF/QXeiBdWhjkCdL4OG3MeoxaBV3sFkG7dgy8GGjtih30EBQbnYkxvmlOe
HFB+7bA2GOpvHDrbcj8bnQj9k+zcv/y0QEiSd6IGH+F19aVGJqwFxve3kr4qkjyO
6dAxMl/aN/5R5SqOxKOAEEnp5qpTonKqJpX63EZFjQXAzNkXI/t3aYRDBqIX4lBn
NwrWW9XCqvAwXloBsLej0FBirVXY5c7u7COfDZnpba/pV39NC1zbDGZcdIyWlqt3
cLT5aECOpfAEtv6qWYHUiheU7IZA5+TbGjAld19dUYYIiqQdnWB8bWjV6XR+TJGt
49yIQA+Zlt5ZcTWDRJ58ULjVUiWhWRCtUD9Njb02SuJOBogDQJ4zM0Szgs6PdUj3
fQwCcORDo1ris/4Sk/oRC7LWFXEutKKVeYiWo7cgQZQykn1Zw9NwCcqfA+h0TKoj
aQPMPHooBen660ak9txqBAHA3bfkLqVJnPrLQWDq9nuO08DCFhgN2qQ5gxW0NZja
AMMZGWHWHg2DNMi+IP8tfIUOpD+/BURqO5iJtwMZkEo6l3+efW0V8P3bW8Im52NG
oRTGomUTNNv4PYscLlFl6Du++8ao0xLNno+hqWBYuUelGraReYktQoSDIeIDSoG1
49cgbqFTZimTiaaDdyl1oqraGbew8lerNYwi+KXpS4Gc4oRNFzqNHBZhIx8gKWwp
bd7/dPCe1SKSPZoOLaB5qrDINxa11cC1Nj41XNxRmvz1WF1O6LoUR+iw1JC5z1Lp
H3EbDoEhK0FHiaru/7cFnaDP4m1b33ydi+s/JrP+mBWlrbrs1bH3uFsB60zea10I
cyUq4B5SQzZx0z4rWKDyCUAXQNGpdZ5L4xNIcVODXZgqe1JHecmsHAXqLq7qs2Bs
FK+VtENzAeD1enSt9VaZ7qrfEZ+oqTJEBcc1o5BHoPzgGR3B2TAwYVpDfBr+elhK
SQBVCMGMO4dYqbjVWZzwA6iBCB4pGIlOomOzGDZjMROd1j8k4pRtNQLdUzWSkzrW
CrrbhZwJk2tv0aiXik9NBfbdKBBActH3wd34pDFsa21bX8w/rtAbhWK358+BE17r
FDM6k7XkVt9Y5YkntNHMKcWEovLLeLWEROztuXEGIvmhGhVOcWt12pvhpRFRSMnt
A9WyV6x7Gny6SONml35XiIqAuEwzXKOQMFhO6qOvEVrog8SdXjqxbOn6D03aCrkC
ifbsIm9MGAaGLBJ0/GivOHK8O3zPbPpZytO5fgpoDauQMFG3TF0xfzdBNuq2IWwO
3Lvf75cU/ILbbRVju7Md4B9YIQ53mnLFaUeSlTeIMbqP52kbMJdTBU4yNFUEzHmO
kPnRwHGlii1PJ9mXmp0iDLW3asjtic3QZKFuFEUyh+QDukBInvmT5qe5Hr69BRt4
BVrF0tmnSddapKLHOtqhvv8h2A7eHhg8ofQQrvQrz9ToUtOw/OzIHFk/KQNbp22t
eVyPQlU0UlpSoo779uHUCuGsY1l0xj5dPAxiFbJFjSFHLZzP4jxx4Gbo33yKItBQ
aSseKkwzJ1CnEf06u5g0fJ0OCWndMKaMxhMwbuQGSXNr6w1WcE2A8hyW2odBXzHY
IDaAYt34xGzHFneACn+ErbbMWaen0FZPKZ4Py14h5dmwkXAAhMQ7UEmDsQRLQJXt
Xsf2y7qGpudJKp6m7CZgFXUDNrPuiRZCxLwQDNxJ5Sl1Djus5mH2iZOJxI+4lx03
yPvd/bz0IOmpMPbhPHNx56cdpp7/gVN9vi6G+I7Im/OlTxuwzoa8IsNKWlCc2ijT
S8pdSw5jEMP0DkU/aHbyChLxnIzdBtJL5a+IWz6ijkgKIctUT39/7d9XWuOno0Xe
PCff0Pt6CKEdEAk1tYLwf//JWK4VzJQHO1Sk1RhFAej48E6GqEofqyQWi9vmMd2H
q+a//5pBl/Atgil7iuVdBr9/mQPO2cP/A4W93YXEVGs0++NBUt53zWhyE882JcHQ
62iHsgEOMhFK5vH4XVh26hbkEvAi8+LQIjkJXwLY3xdFkjde0QoE5oDHxMlcI1Lb
OdHw9b4O3cY1EQdhZu6tY8qw7bWpRgnhnvS9BqhtekU4ht4RJnafeKhuSpuRr5CB
fAxC7DAMLJ1kHmZvxT0UT19Gq010q2ALsMY6hTZORczAtLxynIdMzP1W0HqG6Xyl
Dm5AsDreYXAZg7LuMO9DNa7zJo73IHrSFXTE7cGR2FjALQxgpAVN90rrpLUsOLAp
7/Va8FOia6w9sdTurqHHa4DW7KVnwXNZ22mKAvOdsRgMH4Mzz/lFgENHkp7sN5jX
2g6FA7fgH69XZLySMkUXC8nMnsMqJdiPrid+Lpm4NQoGsgtpklY5aQj1WPKQ4upc
+RUM8pqF7DGvYJdgou2xpRbzEt/ltdLsiOrSacBHMxoZjfNQ3vfWcKPy8JoIhbWf
N40iPVeVpfxTJbTfkfmoQ2pzingk00LKI5Jt0AHIiZBsxqSjgNFWPQb94QIQ8iux
rKvWsx/ZadAZPieJYxOge2DhHS0XFE7p1ZApbmN9ZwcarLNHDZE5Ofb+Bj7RRw/x
rkaUU4BnoHcVSQ7biCOv1M/mhyVQkvOLi1ypFoE9wATftgeKjz1J4ygB8Ce7V8mL
mgCXNIYocLoxh398RTn7i07HcjgTlqbCPrDnduqTBZjrQoVi2bOivbMI+1DL9f9C
YBONlUa83nKYotHkeP8hCv4jKbScMAUQararTAOJ7QKASATAIU0K+o39IlkI/UC2
Ht4jLp/5az3ffZr25YVNpQTzVGxPZMzpmh+FlK/WQitNvedTliERo4XZsbN+ipDY
0WeOkeH9b9oTKg86ktuEbf1yHEhVgZUUNJ0TXHv+q5or5iWuZrIaZCgzX2Se2KGw
8UHzOxjazrGJ0X5rMnABt7e0PHhP/9j/O1F8GOSyNxKZKDeNeLszm/x+pE7l7aw5
hV/s3u4haYwbg2n7eZ1/PhqmeLh3LcLZj5UX3NeE5cHprEkNKKBtVoWEG+YBwG4p
5wNBjlvm8PDQ1/CghDo4vC5L6Esd8cVv9BC/lz3hmvduHCtTcbPVTl/lYuglCMAg
euoglh132IEC7noLrJ1eOh/U8FMxytf828wojeIFBRS/xvKkhsFkGsPpEl8iUxnk
n+FDLe/ihz74QeG417sUssfIn8q2qBh7Fo3LWFRwP+uqzg+4UQ22z30FMHHjQ8z7
M7AJsgtPtZsdqAOdcPwFdbqFVYgM6IsmRSq1r3L6QiVSpY3RLypxXzVL3PRKKBwG
+JgEJ7LRJ3H4UZMwkK+cLvqpY08Gum2kOT9om6vdfP1cQLNLCWl4E4UneeemipLw
cNRZmz+IRBgl+y2AyVma4KWDNk/DwCWmXecMZHA9q3N6kIRRaU5L+9y1lv7BVsV5
q17zlKmjvSdJMtXtPkuu1LWJ25BrkRrmgtnFyVKvPwnxGW4xmaEMO85P9+pzwZA0
HuHfIERWy09W9+J10Vx7A5qxcNi51Nr1ReKiIEsGJo2xO6bUxFNrbbBAnruCmSj7
7ClR9N9YBFOBP4I52NabOq/2DHR0nfjecvD6cx2/o1tSTegnCHUstFQX0zBahU8I
duSuhRUVbT+kCtIMH6uN+NsGiWLJP2YbZB/+XWPuReVmroDuYAhfcJZ0s7hSFFPV
VOIyMZRMP24j3CB4vXUNn3PGzvpKChAvC5MEwvfUMMPjf1/ybJQvVm2xxN0O9ECY
AMvouQQWOcrLe589mdMbQsUZQBLfbRq4cirdtmqmRyUhZucyFSUjiXldxACWYT20
sJLJliFftFPpqnFgo8l0Lbg68nyaOQbyeTEmi9VXdzm1Msd3uyT95dNRfrP18a0M
GQVTn6x2bY/PDB1Ia23KbdSMkS7nnR6amyq/46BdkoTORXxDEYSyLJYhtobdr6xu
jxTpcRtO1nKHUcwmlGCCzBVO7ZJobYrQd7RmNrMUqb7eUI+GKid0XmZgBRTnHzsW
MPwwj39pZpZWf/J3Uq6CKqlydw2y8q0ly+HTdBl8rA+jfQ/5pXSDHanYk2o6+0RK
LTNP1AecSf6PLPBF6fEDKlpwfjyjPAV8YLjMyXhpBqEEV8czBeNG1jhcBTCuXM81
5gszixnGEzSLENIa47NqMNObIzz/JevKl1z324k1JOhasn/PYk9tWwiTUoo5gG8W
kRrTSlMvCvRR0YWahgjXfoXh5FpSDN+gjwY/jfls0FvemducMebaNChxP02i4feV
3MzLwM04oMzMGPFAKs5xA6+EkzDN3mou8xShhPs86uc8y7q73Z6x/ayT4xT7bOwc
L0BrJsxX7MoNhy7DmjrAs0+0uvBLRyQtpuJ/Wa4iilEJLttBN+RnRDgqIzyHEi/0
asRoN+QqsaGomB6Se3ursGbEg+yfcv6QO2h+Ppx4xcQtXmAKOmYrXZc3W33Gt1FI
cWieXsyruEf+Ty0NyA3y1UY+gY49B2EvgjmcAUAUfea5opRHG6dxa4rt/7BcReTy
41Amo70fpi0hq7wbZvCCpgNT/6UJCb47H7ioS3ajR+zcUMc33huwKiNzPTb2qTB5
gxRL1UUIBqbG8xNAx/zBddSl8e7BAIhoiIK0r98qju3lHlUSBflE05MLoKgwu5DZ
cNMO8g9d7axlya6vqKxMaffLJxvvVswu/7TmWIV7tbSKBdFeb+MCdpjb17QjimxZ
+oL5M3vTQtbCZQwn1w8+ELWptHE0oo3aVVwuAbMGaAnBCt/spysJGp7vgWvvMNV8
gL7BJ2Aaf1UNH8BPdhjUbQ4SG/voWzfINRf+WU+dD/iWWNZcNe9N7v9jepgaIk/f
FluGrR/3VxxHdtCzwZeK37V8d1S5SvrYI+vLZb4Uidkn090Qirp0Aaf05bNc4n6G
4VIHSK2xq0MEAJFV8ihYbTXH6Qc3vhRxkkiXPXHtnZU4FMl1jOMo365DGQ0MCGeG
8q+YLTryzu38O5Ajn5yabikEx/fOfSbGk20C2cks0chyGUqLig08uWArI2zGeXyx
20Fpfvhq1qbtMpysDBw5R/Ujp/TGo6GiByD897NMb0XhVC+O0ynt/iORy8AVXXFw
f7fragUrrjT0ObMDVcmxBx0NwAo384ngDe9mkzfLtCWMUu+MvisWTXFv8zeTQM4n
Y+z02GiHrIV/V3YdU6fNM8kekTljmpNmNR70J55sOnkYMPm7H8rwVBi0ekPLoxG7
uHynw2HsdeoZDGsoG3pcgbTmRhHtBUIRonfIZAYGn3iWzViGwD2GCw5kSjrk6kb0
6F9gSWptLIfIb89JYaCN2rte9QMZtzfasceaAVDps0OWSyq5MXu0IRaa6zRR1/rc
GvNZqSESvui/0q2XdXCaoQQ2WAkAoJtfOfMBir9hG59eW+LxphZhzeC5d2pomRre
IuoFlmeM4GKfwyEhA1DwXGbD14OfZS2MiolDy7YGIB3HzvXrgECP4E1bF+wiYbb7
55B8LlrPdhjQjnP/ZKYZPh1FgVQoNniHPvJPgDQA6Gd7zbc6mR4wi7CBWi8HfGEW
V5AvPj7k59AE0wBNciOrQcLDiCO6nnwKDoTR34UWonN6TBzL/dc/yEemN36rJGyw
4c+DswrXEt6qr5kLBEsShI659ggvgFosL/cn5J7EpHKXa9faK+k6CKDtUj5Oo+Lw
8pykEm8N6QjUP5hIkS/Y4xY0lLs07f1YSnY8lZLi9LRS9JnOkj14m22+PKZxXgpd
zN47u+4n1D5UAJucuSHHKONlUxH/oWwLfHdxlOQGWT8BQIfsk5YEwJMa/olXlV/q
0I+e2vOTzjjaD7uLpxeB70fStDd3HvNnTXO322yrqmYfNSTEWBSekhiWTVUQ4Szi
3x3jUwOv7Su+3L6XZnt/CUAfldiUyvBqiLmVBn79foHGUcDXXflLn8/rIo4Bcine
a4qSmBm2VZiAPWL+eXhf4ne5XbyKERC/3MqKecSI4ePH5COON9zuO0uJafv8UIKO
eMYtbGIVjOvc3OCoA63fPspKcdNZBOeBVgfjPe3cZn60aeX0jHI16e6ntc5FBQyD
xLScu7eUamoJdtgiSVeaeW3f3f45xi6JgNYbPEz4u1Jvtlx9NXd053HkKhYuTuh4
GaQFiAH7rNcMrTjP5fEwTZQvtbnYN26mb1b9RsqRDJApx48z1QLNDpRrfLy9YVMn
/2r2sqktnO52v3kfGDkTOpxjuf4ELWNfRLUbQlI7BCZLo8QGQPCiFUSoYzBAoyS/
VmCUFaqoP7JcP6o/0PlFWLUKs/g6ctxid1K0+htTlcGH2QVsjhdaq8TotuyOvxfn
Icki/0HqWzzsWz4oQF3wuWO20cMPWFebmGPeYz9ymZmymVOLHLhPaGUsQDVrdicZ
rVUc4ZcpUFBv/DpA+y2g10bcErkqWn3lLU+RimoZgGRMpvkSJakutDEXF7RsydDf
5LLeHQQzb08iXz9+JEM3ZyQgSuYk+Kt2AOjawN0QbHTmv+bSVYrzlTTeFHmlFeDX
+06ODBfNmzkKikz3IbWUCYXZ4S92P7NL2/G8vs9ZeISTYHG5bomWV8Hhb0E5jkym
xyGJZllcJC6bDAFF4XrHazDqc4FfFfhWZl9rULxFtGPtUO/uiKmaA9veke6RrSiu
T8RO9QK0gnHK4gtjr5SBVWKHmyoc5ITMlsEVH9bQ/zc/yHYmPrYGNbtDyUw4LURt
egtxMkQ3RZK1dKeFQEzYTPqQLPl68ouPh6z3qvq8ircDrfPhHiKsRlwBt0WFU1DI
qW2ONsPFAa1Lz5E46KSGFoIWjvYKPoZvPwwATSfN0IDY0orwMjep61hMzD6LRVj8
YduDm90vCupdqqrdGn1oM0IVaAGQNvZru83nImNOpqmm+pjXpGzUyPw4ThcsU4kS
YECVp5sYSeVkh9XcU9S6CWLQfBGOtwRXhgP/3FKigU6hGZvPJriUhiYs5XfiU61J
VuXbEQMGarB4Th5ln1sL0k987BWlc0QOHTEZDkxVPotgSpeZ/S1UKoxf1vKIJHjY
t01hs4awGXjvzzrNfPlwvGo9tUzSyI/v1VSiOK+FrHrDIvGhORYfGQ/VQJqP30SJ
8OflNsJDgTLeuJfL7RkJ2vHCGmLiKHhBteiL0tnqdJzsrHzh8q7MYq9xj9iBKvh6
HYSElB86bCh2l0woeSZjqspPiy3d2AdBaiHcbZHkNjB4YZ/8wuXvBhn3P/XegFBg
GzrICVImO6AwtPl7kbCqyfxMiLPLvy2PWzEEHGaLE3H5SNOMrjKgmY+MkDsiVdCW
ZuUcyn9Gq5fZMJetc+HPBbuHf6ONJFadltKn7A1N0TgSsTVMjSSfa+QQ8+N8L1C1
1B5925RXnHUCgaOdyRSXjyQ+bD3FXdlHvjTaj+ko+i/iItevg/Z4jpWqrEeOAH/c
Jm1jk0D3vAcpalxvrTJ+28u5v23Oagsj79VPvAbRpdJUhPkmla4sN+bVcvEHyP26
dnr8zSYAFQIHrnMo5jgnZP+OEAtFlFM57xfwO8YHwLMaZHEinzUc2UXVvL5FDbl/
nEB+bUhHz+6bvutJuhOWxFelB7qGuVLffkJe8+gzu9GAkJWmX8ad+oUGv/VKzVCc
M/cOoW5kOMTuc9N8IhFVRKuBh1qsfExER9GrR9VETmeYFuQjdTwsJF9owOeUpRfC
uwaX30mpbDpdCozmcFIsISlp+fTmesP02Nc8OLuXefgwvFm40YSIQcIBFS5AYi8o
7BWgieVuIPdBRerZ7wNofThVLyEztB9TWXw4h5idXxZol3HpScDHPcQPWxR9BeQA
qo2yckdDdW2ywV9qzmVRioQX+yME4xyC7Yxh+s19wL/TqoD119Yw/3be/R+MhF/9
lgoL+VMnR7pYLDX3+Lv7apPd/bOPdxs4koGu1hoHahaw/SlA8NubfiOzfSOGZv9f
HFhW33fZEZOf+ipPJVJYbH23stY5FiAHWXHHrlLt1luWJ1Pv2acrecrb0lb8wSeJ
tI83tr/Z/voShDygALtwBgrtiizV6BrLkUD9rqJwKWTP8QHBZvbyiWGq8VOMUBvr
88EVphAiUu8T2ZGxR7myvGhrZztFbDdYeGvhM5NU5guw1Ef9n7VKWF/8TmiQgafM
O1jYFvsCjma2uIeTX002Bi9aNUgrr5raPxu0z71SbiCSYO768mcUvWYGGEaeHfWi
HP/v5/+EyimJk/YrwFi8T2MHZdefMDWSRGBODR2bNLa0PqsnalyqPVw/eU//ksYH
0e+HELTu7Ii5BjkT5UNOUhV0s18B0YCp6iTPeHrEGdB04IyycRdRKzNUQiBx6s3C
GSSnfnHTEN1Ca+WCbW/QRvjoOW3mA7cDvyvLq0ZxPQ4vu7ucsi90P7t5t+Auxfme
wPpOeSEEhBlPzyFgAFVXXH+kkcpYHCYZoE6nuA5kOTwFqVM9FwBOhk2i6/Q9Al60
3+Tq7LFdUw5IMBgPQhtLDezZO5rYhCIVfpfaXqyzTWVOENbdsGZqPVTfo28RhxsH
/0fC4s/NddxDJu17qs959F2uQPbyW8taG1FA+S2MOvwoWS3cvtcuqnuxizpJnYP+
AjrPKkPewkrnqTdjNEFBc28VZMa4mzDe2OJUz2UyPB5DvJ51RTZkDy50QnyGuktX
TZ+EeDIURcirruHiEXXSZYI1UzfiVZZv3Go8wTiw+SF6nzKoz4voI57Lq5SwiwFj
356LjMfZG9nMySjDwIVMMuRHT8rHrKY6UE/eTb04VglNfE1kPP6ZbTEYOY2ybqZ4
wyBMIJNrvsKvjHEkdXMwgpOQUUZiqZZc5gNWI/OAtKll4Zw5CFS6tTmdG3FcrZeO
jm7n1UJaSJa+SUHN6qkZO1JLTG+MKmgqFEY9LsWHzY/BeJEGvN+BRSQuNEuvmqKW
ax5uGS45L54mRNPmQ9M0pUxJL85Wi0B6BPWiADpDu3eMD9R/Sw/3alkH5HpOF47Y
ZlCa6dMPcZ62oxsE+aXzNGJSVTf8Jgu34QMDl03GrOIFQ7iUl0TebejGuzotT2Rd
C/bMQR1uNhxNzqcMJuzSr4TZ/LdFngxVJE6DdGR8zLe394a12YfqW4c/JUlWdMG8
0dWa/9NL7t8s7TlX4fokuMb0pzteKlxvWYwobiPD+lKlR9fT4gJD/eskJ8bF2p5Q
r1qum0kIlSd/lfZYfA4Gk+8wWiJJqnjvHXCQCpLD6M587pNH02nPIkZ9fgb3wdb+
wj40xlcUx7N4GgyYcwFf3gCo6Q8l6xUjnnRAHDICXavljeVIY7A/osbnlbk+NU/b
9QnPChBsCHXAZggzLaWm+j7qzBasHJvcmRoX2Ml1wUHm1lXjChBQj9bIMZmuMdR5
dEbMNAtCwXWXNDIsjYIwd6zmrEC37URlXJblZFpcu3zelq6M2K6OmpMzOJMTWryB
+DVyWU+MF+8LN2SNM94L2nPcsWIvhFxPBDNDqi+G5a+5tZ3NOcsoG8zp9GxQFowd
dSkCsrPhX9jYAtlstEAbG5V5C63IN7xtYl6TS87p2zEO+pKtb1CUSWjPzZtXJ3yF
CA+feGsQTpeNu6MQ6wt9gtkwWwPY2+1+bXRsYWLN4VYOGrNiNY43s6lWPQdr8QCj
l1I3oniBZnuoW9w8ZJ0aB9hfj27GpIVcXrcOpZXBI5hNim/kDs3otL8TmcMvwM2f
TYpvlvAEr26xI1SViPqicKnJJrdZQX4L3iP6zXMIdg9bAJELA2PfTci/rOhn7WmA
tkckhZx+CyFYqQmh/sjGah+FZ4ycBi0iwGijeSCni6bs69u0i20yttXEbz9Df9/m
4rIQxblsBm2hSfq5F+xUYj05BGmBbVAU8PydDsbQ7TEKgTOp3d6/T2HFNFTNwDkc
bRv+Ucska1xiY24K6hy65LLYb58uNGSQ/Qtk6dq7XFRMJ1RtOG+fZV93bFbqCDlM
e2MmFDnh3jkF3uHv12zU4gHgo8nJ3YpNztXzFS4rsBruUf+R3lZGAQgFy30P+RaE
wMMKfgV0ay841OlFMGPKwf0TjEKwCJQfQIa1IwcS0sr2VaeIPZNu47TeCmGCbKUE
JFJNFVvFXkN19fJW/KVJ22w9iLBIq3uUjCxT9e4aoq8QSRrHVx5n6IlKSlTQcQE3
eSP7Uwh8ZQxGwDPy+uhSZfY7Nzp3HPNCQCvi26QDaUt3btb+MxHIc6/4mhwiGABR
OT5sDlS3hulmOanYJAVzSwjqH8GfXb0lPbItcs+4oGjYRmBUQPUH1+stHEJE6mXO
TiR5xO6QWW/ORJJPou+94kclfqqKWDbbntFtj2FMA/oyRjxOaHITFB6Mlj+BU9yW
rJb0jZyTQYS/Q9oHk8c/jDAZEsNKW9Tmbq5zLFKFsAxg/rZUguiZXMUOcZk05eJj
FRAIiQ411yV9/cWvUnUzZ6KmSuPV1kpZ7ul6YgkeA17F9q6x9ZLhhfwDAKn8TTvq
pdLbiGj16L4tdwJkj+Y/e08mLYrwsuSOP2VWnGJUdQZTHv+O+uKJezBULSTAXhpb
x2fMI2i+ee+vAqpGXc9ytCRvHXjbPwgzcTnMnNW/3tHXN/yoBaVEY2CBytmtTu9E
4hR8kYJqgnBcfNgQyXaLfDH+t3nAB2cfLk+XXD9avUDI7Yvi/91/Yf/LqPIwfgcM
y4ZscfdgecdWjN4YQx6GRGXRmJrATUeHg+T2/es/Z9Ui8H/UDtvl1hL9kIoINJGP
mvdNlzR97vLE28WbW/q1seThT0cq2/ToX/pItmtbrOdpBik4bK58UAQFHvXn6ofG
WkioUNSRcUAfzOrvyVyhVQlewbLesqNCwHWzg4SFZD7POgSk/ANPKTmdYPNQhrwX
RratP7FD0eu3elD53rxH+aJuSn74sOZbxqr7KSGjAvMG6VYnSeuKAOMInWVeo3cK
cB/VBL1GoLO3uRX4oiVZ1GycdZNoy8Kf+34aGPBV0DjOGowFx+XtsjShm5A4um1R
QQKNxF+Zl+UOggSSkf8Fg8Cbf1nY4MZsu07S54cOj5+G7gD5G4ubaX9tAW0kPoHT
vHNb3LmcvNR+M7S6q+nEABVN8mzQvC4xYVMRwb0KDYmNWZyvxQJvEiAolW0EOZjN
kijASERRwLoS6iwA6iuTCIJkBiaQc+sHofXkyvcf1XItquHPQxX6Ax6qPfRO+Z18
qN6kQ5rUsShdm2JpQi27W+J7SDI1SVm6xqC4pfgQKaSRqB9/9kXaI3COqBYq1QMC
3XoRCNuH1y5+fXkspSnvtaq1AhQ7T8l7BXmql70b2E7zN2QS0UsVCtnCHlZuYiLM
xY9nqyfK3XC3xyLyZBR7PoaXvFU9AjLiISlOxQfq8SR0sq+n7f31023Tc9TK1p+O
XifOo7ZZu/0qu1HzsV+tMOQLQjh34A4wYi4oo63lIPyCDLUFgOq2Y7/07jJJ/Sa1
O8WnAqva7CVcpKxpAimAw5u8yq+TpRm6NTPm84VX0VrTnDZdJixitHEEYKB7bHLq
niu4GeEIWEHuG3XoNMr98cLjp6HuRZm4WBFxmR81zsKk42Pb0FlLJ3bq7+yORuWA
7CesS6ZtCzuD0AqZENo2ODunGfm4H2kCBPg5au40yj7CwfY2dNO0o+/hcIhPWGea
06r/Qo2aQAj95bAAww2R3yBspMDsRzSSR9lz7on62eGm20J0DMRiP+bc/K9jWPdN
cKiJ3Wk+e4knJ2cl7G/DgUXE3rmqZPaeh9KwsE3oAUjlq+UZESmkwakYM9UZKxaV
9P5slsILVCEp5o6/MYpidtL8ZyyvSbyi6MYjWEVeErzci8gGWrrm1q3X2tR84wQ0
a69R3yNr7s+sCVLrRXhKDZe0WBGGgON3yV/AblItBEEr7rMnZbInL3Awhxdhkb5c
Q+X01SjBBvhciVVPQ3eVKcLdcn4Bil8CEAXKbINdZOvGId/zFo2KzZXbGU5s+TsM
dNMny4DCFYVlg7nDKFOfjk4rSSiSxt5+oLTg0Y0sOpKL8IDtUnGmPAP/sgenDB0x
R/QZttlkcilQ1+2LjSZrKuDQHZQ1g7kiHb8Lyduw9WB9ASNmiYjILtubQtgKG3DL
NUclDWiuWRxoU/EkinanA+zZpeM9GoI7d0gwup1z/OTo3biNCpecIZY5baS+HzVV
+Qvtbha2WKHv02GegQ4/Gy5BBiKoJK+5hFuFSXYnOe6spHV7c4OFNF9eZHGoo78s
K6lTWPZ8yiV1cWyTzmZfHWvcdIQsYY6EtWZh6aommmP1FUbX+zweu52U8nUj8dl7
I6cEfMgbaeI8zseH22oRkDWmdTLyagh56IgGdbDMXfn3L9g6vS1BmF3qzvpQeypH
g1BxAGngBYeDpFbhFcQt28RB7JgwTwg3Q3zIcDlk4sbxsEl4Q+FNf7idIE1/N1b9
o0dVNWbpSyGKa3MwbMnmwHloHpNCxh31M69rLApC2r7Ka/GwiOFftq0UB08Nioro
Y6x6eMnivfqwk5RLrlL7Pe2YdxXhMRPvmKae38y44ox25cpafzLvAKibVhl2QtME
piaC3cisr8WPgys0lM51FukzF72+TaHLLpcLmJ838AGnhnw9bJG11ijb/14RHlfc
dOi9D5RdG2dMacl6x8BDLoxJ4y4j2nO6quVT7UC9cyGRep+BGo7mB/07KSAKDIoM
DavG8KS5YofgSfqZu+cV1rfOV1CiroGPxAHYKtO1UFZOn/2dxAbOx6tzKRWr+6bt
jtn/OpNqK9lr3ofilT4BdnuhrQD+S12CxwP55tQ3+gv/fMFEJC3+88BuQN8kcLgw
4N9bi3jwVyVeAo3MoV1yuTLIEyG+cILPEgfiUwv2MIWvpz2NC8VOS4QPcEspd1Xs
yZ0oIoCBoC9gGxeYnUDv1yZRKi8xwuSGu7hXruAEOJ6G+aGx1fg60iwcjzYR0LXk
gIlNaDv/rYm9RQKvcowLBsnsGBn0pwo3W/UX+/p7u45a5DP4aJQbSSwHzo4epND6
X1sIG0iu2Sqz3fdOwet5IvOCTGo3T9lsWbJkavoQ55d+y8s9Jk5ns4IMZlI3BmHJ
/90HKRfT4WXuHKCiQL/ir9FRpPucTIWUNKlqAk87AA5KxBnN3TiQ8M+4lFLtwx+s
36Zb7IZWpUhQfc61iuQ7zuaXRVozZjRY6O+HWFT3gz0Lo+R2vhLuJMFFNE5Ql8f0
IHobmJcpOcFccPLTv0B4WHvAS0dt1YJRmE9hhUigILq4NIuhlr7JqPjfk6eohXmr
tLSWDL2UFRnCY5wJAsjgC7h6V2nuwNQlebM3NvS35JIexCkOp4bAZD+oq8XSBZ6L
/eviyYXhzxFptOfeQCKFSG6iq+qR3jkaUhddgejOasjx9r0wxIVw2S8NT/e8DHF9
0QeuK4hidMUvMLLF8A1tpS1qsrHw7ZTs3MPtNBrkews3SrUwcU98A8qlOgA2At2h
/Enx5FKnELtnximDd1TnaHF6lJit9wtSpWBsOHwChaWP3QRYm80rQxc6Fdn/MALD
f7uEPvdE7brodxUlAe28l1htOINNsTesoK87xVSHBYc9mCOoqKeB7XtAQalG/rAO
V85ZAzUOj0TEcS0gDq+PA7L/4UzXh5DrW9mhdsb8qSnVcx19NKd/0avgSBXFlq/i
xg7J94kODZwC6Htbc+o2wvZOgRDwD5dQeTXtDQ9Oo6/H/TOFaTOnJEE9WhLc2iu0
Rybr/4a887IN/szokkEv5nfGlB7Dp15iNV/3+bxq89SgoGo4YUDsCxlyFziHK4SL
ZvrpUdg5hrh6vYORFnDe6W8fgvQbKC6XpdjlvTqui/UcdI529SI+ldRepcY3myyG
S+MTG7xleCuCDVOP1DGrA5FaEANVKIK9BKq/LSTqB7oDQ40T8qW0wB0r9F0XeZ99
iv2qdgJBGYOPecV4RT9mJFJCeGdIqeUnH+AcwOBo7q477+yWdb+QGitdO9QcUBUn
dWph9KcrHRLI46BbY9YjQpM0zugFEI0XFV7sM3Trq3SgJnr+MENd39kQ+8oPHwNK
WYum/RzZIRuq2jLjc4mikFY/k8ht7N7c+edu+l11pEyr4kZOA87yz0u2nYxNEvee
EOHZ3tbvh+FCVxO4gCeXLVKkiOmU16y8KvZQ0Qgadtlhl5Z2CZmLaxm3ezrb0Smg
jK/FXew2j9bKK5jPht3bnOrE/E9khdeD0t14qXND8v93k+6PKnW5pq8pAwGjRg31
yokOkxrEKZX0NOEbfjEmZzx1/rEGBz0RJcLZkMhQ12C8oUVg7/KPD16qvA4Tn0QS
pjjO2nlR3BPo5c3J+qCyDwNjDcoZhip/Y1pbVLUvKRKXhmnTws8ffbz6nxsXE8Bi
BCC2yM+43pWHPWuVHxdRb9cIsw2haEXsbzUYmVT62Jp9TFwwMHYK8A2h9PaGlppb
qky6QU4T99zHjyGFdUNg/Dxwq/rk8ekoRAn335qCcDXabnpSy8GaFUTWBo230pad
NsE6Ckd3G46dXPjsis0L4YBZBNrQiuzkF6zmEnGo/h5CKwDpDVSpK625digzlKtY
EW44ORRn0ydfLk2+dT5lMRcUK0eWo/gRWIyUGeRAydMlBFHGMDZtjZwoYUv1eVEw
cavkFBjNug6iGKHxnRU8PUKPnHGs6V0LPgszHBFmg1prm6QwYi8kY+FPNt/5Pruv
8oGVYdIK8dFAPnZg/KvDUoNlTSg1uVs7wfftSQE4M2bqNcGjrqNxscVEbnELtwYi
I0uoVgrFXgLUGu6VH26C2Ii3JWzf0R1/ty3nsDr06HNIjdEpL8MUuT2/ayQMyP2+
KOn3ZG+Uy2JYUg6N1CN2ef8yG1geH0H+gaP+u0jrL5rG6BZ1NmQPwabbjb8add/9
OxE8Y/Bl60sgy64rWQhAsZI01479iu6LcqlrOkKn36gqHMWrWCwsZyAhqdQx4mGs
pPGhAJ4JHF8r4G54DtBfUz0QQSnYPxQflgjAMCTAYQ1zDBMkbzVeP9kWZQWOrx2y
MH3EKSdwEdzgatX9giyJrgBdpP92F+Kr9XfZ/m8E9DUEWqkf5YjW1jBZ6MDzOJeu
IZ7Qt1M8khvf0vqV0+HK2/qhdKzUnRS5gVvthWfqOKRzuR0FX5ox11egqDgWME2I
h4P18w7lqH4m0uEF8Djiwop9qSmnF42Lg52uDdFdvcCynpsw/LAzc7pMOkyPx2x5
NstALBNhpsQFbI3OWhowh/6bgLoResN+fhrH8ALXXDmxHIzHZHZ/1ZfO4t9Zz88Y
MLdCOz8SYEmwrITUL9STpd9CrnJ7JHWG94w4fIrxc+HuSWju10ge3rLa/UQtvdGQ
ndKVDqYYUorU2JxnM5A6NuXq64Lil+H8hcCSxNto7zXPWuZEmFyerquRvonBs3Sr
PAgFOIBFYUJsxN/3i+jMeEZGCQCHh9Mb4IDm0kl3J50vv3BEQ3V7NO27V3VyRAWz
XJ499paah4+KBkpWe7D9Cnz1KvGOmlboiEa9Q7mjfOJyMVronvHe7M8P7gI+sNMH
UH9vwHXWExvXY32t/Tk316s4LsyzCHo78R92mhXe8LQWmLRTes575Dzs4J5sG7zo
uv+6+zbWLufmG0/ANky0cdyhDEA/YvdG9WBkloXeop3UHRoo2D6PzhyPdiKFWru/
uQ84NEPgHj3sMiPI6WVTT3+OUxqoJrUr6jTR/LfdFEjB+p4mLUN/P2DWjVcO5fsy
OoCqaKNeuwGy1nlXxYpQAnrmoa0kv/K4svVfbHcYEUpEXT/LqM6XgH5bFepMyyDT
t9EYsFhAsWP71qFQd3KRvp+KYEW1uNYDFyYX8/iYEc6BQI8YaA8LsYTJDOtSNBfc
VedNMn1aIjZyh0sAGlAjIADEzMg89yVvL71b1/4uAnPOHrxyj6wEY4j6OPsBxcam
9pFMeMLYWHABBODOweHKvazF2RAo3Z+8RW9Uo9h/DzTFUfaDUzCl4GotKqEC3v1m
FJjE/FhVIeuZYMFiVg9YmBy8USlsVa5YWZPf4XDp4ClcsERvl2lilTPdytLBNWvu
8kyQMWykGou1skELtNz20+KvPEUzV6eQw7apW51z3lPDG2jSUj18E14pTAUFfwcC
3PCc/f/N2xMPkOBAd/UxB1ZWzvZicNkoHzV13onDEbulFmJ+DDGTsvrbp/+V2JhT
HQhRUx/vvnkzXKZDaGOvwJvhkrWkRzwv+Nr5HxSKbHLYvRTYu9a0dofgaBXn5u4/
b7J7gw0RtbDVqq8FgyZakPJohAveXqqaXLeou/zZJfUfrykzENUkVvlxRqoA2K1u
+LdXKV0XgEJliJdbRhferUXV2fRuw5/5QXY9iLGVlDnsQ0PrzGZXKfP2vN63PIJc
mH5aLsc6Yg6yoOROMqkfwVZxo+Rk7f9ojxLgYH9tfIPLw/B/O8T5xFwz2mNh23ih
5f4X8d7sOTC3oNcclRPKnOUiALUvhBumuQ7gC4PW20X/FU4CBLPlhQztz2Rf/cVB
BHKY3TuBsuM7yWP4m5J3ZOCLRkVPlQmJtLXfxxxoUdmRseUzCh4UV6Vihp8Boc3k
17+W/drdSNR/XMAmWuJ/L0Brocf1JolqO9j/e1r37SEXMWS6zveObGTUIx+gUq+c
2NOTxBr+mu1O5SX4GmRM/G+UWg7qWOb2EvE1Nfc+9h21Uu5W9/OwaTcIU4ZZ8f6K
n5x5qOJcgMUeYMf1d+MJtmC72t3ydYXB/7WcvQfGg0pmsocKbkxkTIIUWRaeFib/
z2YDq5ER83p317C4wWjpHTm8mi4RXRKzgCNf9VJMcdGNO/KEdQ6Z9Tq1sl+y0BqI
arE7uDH+bOmHtz+0+Yj+J7aMwLPIP9xPW3+fsqZokt+MFqNNLm12vA5AEV5A+gki
NY1Mq5uKnZz+Cl6xP3kLBBcpHI/i7b9Imu7Q74vxTYKCyRBCunKTD/f/SaJBFo4t
ol64AMErwTNFTi0kDxJ87L1AM7ihW4rWifXBmL8DmDxWqrpXlt0s9cNFLRyoIXBE
7ZS1sBa7uIqqyxQ9csERBwlZUEy+hGrfky14atn3c+X4p5aQj2Pfr+xeb8V6TYZk
XUG+PWRsbXKt5dVYplZZ32Fwn+f4jXMUZ4NqORJN+6lVslnKecl7NCLU/V+zHRA6
gD/me5JlsAwQi8VA0uvZ5XHC/EBJ+z1AT7py3E9VL0d0wfOPxHnlHcJ33fMttI4+
mO/fbokPKY5bCo4Z19nMH7Uf49475Ez21h6IyFy53eZ8FZcIIQ16f31ujhj6OyaK
1gNq10/+IOIKYC3f2I37KiTsYoXT/lWksjTK/3MZPRduWXyCSlIPybR1OiNGdbXi
UdARp3x4DUNHYe8e3ADUJC04qqBIlFCoA7g4P8385/qPpMw+KLgA4dtPFdFSqiWz
GYeRta+IeKeUeBu2NC9/BGOmh7U8oomuZvSzUm9dZvW1P1sENssmvYCv04LrNNLT
M/+bM/BczNNLOjhVnRWR/Jsx0MpreZkIqdeUdArpVVBR8var/8qfjyXsbvRLO/21
m9tXKii/Bk08FnOODtiUYirLZaJKjkHBA77GKqZnr59H93rMEB85vCdx+/QTWAKG
spinYQP55hfwaIJrWWAd0giRyPRBKZp/+rdrHjmiBgmc9gvXJx4hh4mtDSkJuRsd
0fKSDeSh3HPI34NDXDJkT5nFyIN8xQpIIE+uHXjZy+4q/Re0CtKUILIwYvltTOPw
xzdrxvGYEGvIx7G9fKR+GekqMyAx4sMIG54nLVZyJExNZLBvmGz5nMwH6VFzvqU7
33MkRvWq3WwiK3adA8BGUzM1RzQEM19upJXUOY2Ejmz3YDj+8Cv4ijSZMlcUS8DN
nf6/SENhvnk2sFvIxiYsW1FKQZaPn4y3MEYVhJcbCyqCNNYYDeZ58cRk1eQIeQiE
reTVaKXR9DFzr5l5Bz5iyIIOdnb+V2q0f6Eath7KXCqXolUFWlx/wBgnm69Vf3m/
I+9zJsua4PhuCXzuDJ04Jn1BpmzkLZAmcZzfL5XmSPKiw8/233VovCRk59xsXq7u
iWuiC+Qc0VuAdddWms6c26frp2A4ihE/a4jZ8pVf6FDT4TAp5mcTzmGNvpG0eRNw
MQyYVVmvOsGbXONRs6Cfx8UsNkawbjUJt+ZvPXVZf1+yBl8aO/Vjy5CbtWtygLir
30rBdEWF/NTmxp3M1X96Be3/hwl7lvs0zg2O3UdA6LLmEf5CUH5zqp/eQE+mCeFr
k+VTEySq6CwGRR0W03W5iZmROU21W2aVHbtFPMQl69ASUy83iGKMk4PQdVrL4cP2
s9ZpuH6xx/4ECOB67Qz4b4nclV9E5Gg3MIwRrfH26WmMDdI0eGwgTf+V/eFuMyYu
uoYIveRC9QfAOAruA9EQcsWeThK/2F+DL5e4ANNNCejjpwPFD0N8kR6seJOJYvdl
l958hXdXD5sPixHvui6XUQiNkak557crweRrUeGUZBQyJbyTf6FWR0Aa7idiVm83
4iI/KUlzBhHqB2YMPnkeMwLzfK78oH81KvzjoqHsyXCS+9t5RZ1gleYlI97atUqV
JpXyn/USrX6hZYh1/yRVtB9LMpwrMz8glhUpTh2ElBd53gsfDTrUXzqwFQ9Dne20
FNUcoDVjphwoGpKpYauFZVNAPpWtJMSiZuHfSn1lSJ56jILBXxcP5+Kof2iuEYB6
eQbaY/8QKmUk8UheQEkLICl8Q9jr1fjWaEXFstzpMHuctEBEibyEzgSf5sCTPjX7
BfPwE9q1Mr0uKyTjFB4NT6AyLLGIm5wMvK9z1EH74FoQSUPqPZ1kKEsMIzDSRBQk
i6a7VD7PyKFIZqPejk67Hpjnvi5csZth1V7AsTrMEpeGR+bkmhBTZgwPzjEjJ+6R
xiP62hvQcS5KdGJlUAz3cfTSdPtR0ZAVXiB3CqrdXEKU2QhfVKhHx34FiIVb4fpM
ekvo9GUMm/jHX/DjQfnmVzFkSHlSMkrvw7QnzMmYQno1cavO+EPvcbySQEfmxr8z
NKSS22cwwKelt6Vss18eUJvnv+F0iV8JI/EHxuiRktAF/pjaibfOojhdCGT0P3/S
sDClxhxdYGD82o//4zxEn4sA09VTftNu2/2MKtEMYD9Es+2ANAybJAwGRkXH4WJx
RqFwzfboXqohgoYa8CbNQKgt3Hb5yBbGgWHYMmGqzmSKDOt8cbji8bt7Q+lAMLWa
/EInkc6cVZSaPXMoFbje8c9xThoXwQY0hbySbYppgi0VmXVTBZ/WPODkIcICmOyo
HdGdInf0ZPRaE9YMiOClkVzQROQ7TCp0NMMPRB3jKJBxkvNmjdt1taiNwGUjyeqJ
NkMt494QbImDaqZB2hqzWRtQWzhDaOLoXdwVzpxMto92mDVfizTL1jBm37H4RL4t
xXRRFw6LR9WlcrNxs218XOmYUoBuH9unSUQmr8O9lNuiywD7GQbzgaTzHwF30KCr
dKlB9F0TJb4wqOYY+I4jM4cXFX8xX50lpueSHx6JQNtlNQoiVXeMcRnRANL8sLFK
TU1pkLEIDGB7kBEqkGQgRue1Rck6ZeRzSPirg2orBnYkWfJLJXB1Qc5cTvccuNJ9
gSY8b37K/tjsNcpbYTlUvETT+EF5dF2KBS4w96p5XOhhVO4gSuVj7vf80Wk77jAj
yjceInj09WSO6wiChkNztdx3zGEJGqOgxSD7dksY6dfrNnzJ4YPTcfSnJLW+4VQX
Pd2FYSAHou9T0okgBD92zYHceOyb47U3tF+8eE8moWfPJdiW/T2U7vCIJcs3Tzik
FnYTClGAV9ow+1LdFM2tb0xo8wqeaESett+YUVdHtk6vJcR8Y4h0c/DDUCDum3Ai
YfQZWFNPqiBgXG/WsI5d6tLOzGXadbJ6Y+gejvkOqaOPPC9wVMMLCLDSdecg3242
NWNb7kTqqO460lU0WhAo6mpTWbQrLGcfkcp7SYl4h3aNwCE6U9VztzZFP8cUtuc+
95rsOLdd0dxG6vQSBYl81NgRW3dROo6uwnJt8VjfIecvp+qEx93xGdToaYyTXQs6
y/PkqV330GuCmLe1VjL/LBqUypt/G0pYH0l20KJZOTE9iAEttYWHfDFRZCOuXWDB
bNRS02kOaFEWbJHt0Jg7S9unLDWh0xQAUQ9QrJJyNfbqO18oyevD9qyo4vD3N6aO
MiG63L1OvVskqceabrNAqF8cIxNqtMR8lzXsARhjYfgeAiJhjul5kAX866DVgU1Z
bWhJmlY6XAqvv1P76HhQDlBSK05pcXgbWas+cVD6LLcSsFrEONwfTcj3RCzjUr8N
ONm4nQGfNGkeEWBY1yIooF5B0XFKsgbU2TcfO3kH6VcYGALltFi8oGdL0BKgRV8k
XmaNRwTJUzG1fpGFAPQ4JhjbnRY+4Wb+BpMxUBFZGttf0bmFJkTIdCNtkih1rsQ7
MKQb/3Dc7LN7PX+k/o5rcv3hWqt5YF2h3KKcqVHOP3QLcsSlG6pfgJ2vfeEUVkoa
C+TJ7FltpRd6uX8DEcMJa9sTf1pXmL0ybgzr2hFfyEpGCYk21utAkgYhKMODItUS
ceq1yB6X1zctfNVk3IajXmJNK7FDaEaGhI6/3nH0SPBGMHYt74XoMW+ePyE5VzCg
yQ8ar7HJUx9Y2iSnFYlM+uWEp5BnPuNH+EuDV+IRTEY2gu/NVs+1jLzGHahJT41b
cmThyGsNSwHBif7KDHBDFG5Hmeo6khajiWGWP7FLUpslc3qP4DJkIWsm0fwWlbzn
nAzXzmqsr4A1oIb3N0HlOXwPZrz6YFyhcOz4OZHVxt56TeXME4roh5UT9RV95t6j
EBBZy596II28IbIzcuUfBS+lLN/FpHwvxlSmfBml09lsWxr/IOzBuGu+7nBhDKLB
ZC22G5DnbEjhod8iPq6yO966vR3joAZAsq4BtD3lrXiRKNeegLUULvRmkS8t8kzR
ffcPFvVPBYYJWqhhcpG5DfJJRDpvqB530sQuigeonrsKeszhOw7ApMaSwo5mjCo9
azVhqEq5dMGwM1gwm76sJx4/h7hldCTtugvnLYDhGJCmL8NBbtcF+rtQMAjKF/rA
LSEGMyvuFF3GCcsvNHlmCKo0dfdi5tTdv375RUvwSM0iHLgqwPUYOBeZj91s93Xk
6RzYDiemyL+j3Ntjce3G6Wm5UfTRCeoCfFmOZzv3XPU9+Bakiz2/jrgCv4+pQZsh
0YV5pdYrtOz+gQldeGkBB/Zdrt+RN1Ux00qJDCB5ufxx0XjThFkRygBKTtJ2ENKx
b0/hwNTsCj1wSvYVZ84COccNg9pZPYWez1OfpZsaAjNgxPQAR7dCB3MzZlqdFdGR
ki6wSimL2kGmaEkD6nA7VCSYKv95eTJIojOEYE0lP+5WEZVM+uJ2jl30X+weNpoi
N/UWrUkdacTi8qZzpozloBSL69ZEVmyjP/DTWoIjQyLlT6tqpHLqDPDxDfRStUT7
1oTna69ijMyuefCgw+L6LcJ/pnAENzD5jR0fscfxCdiZRvIDIXb97OyQuSzFRkKl
Vv1Hwev5WA0xFfNiJJU3APQyHLJWGB7U+395aCMCiZUogER1101yMvNz7wlyZxMa
GISBXT6DFSJm3L+Aco347aaAo42EXR0/eeD/16u2qodNIdGESr6dOsLzN100RJvU
IHrOQBKmUPdW7Y1SZrxSX/eiSYJmtlCBAlkiflymSla6PLkkGYBv0mOAvxyRWNH/
UeapBaa/m/WNvAUuwRwIcahPDn1sQcuFVMwE9/YvHiTXm71cUTWx3kopjvT9lTiI
rDufN75Pg0NV0++uhatp5cR1GwA4glgMyGVva5RyPvZbYu1yZcGLCdcp89IGwm4b
cWB+A660TBib82WNaPtRSQaY1OAX45ETZx1FZdnEeA4GPcEwpBupavMuWZYLfNKN
GcWPskUBOzf+xx6vTb+ijuKGppzyIUqtn8W6mthj9lwXuPECRWktOupuV8/ao4+b
cpz82g/MVCT4s+BD3ulvTu80fpA+CTpat355MI/EvtxTwaQmpCjNmAM29TcZpp6C
L+RgNhpE91E3qJq35J3wiKLkj3fSvJzex+pXm0NOwocFY52UXsTuA5Zy/SqgVxxT
WS0GBUARLoaODQ/rdz4lFYIlfsFmWSMsqOxGIRlbmRDuyD6yjbv0FyeEgFiPTjPg
E5Wa6+V9LtWnIaNCemhGmTg4QhQyoGmLUpb5S6h0Jm4b0zDtAqfigXy88TxZQTB7
XYCoMcLSBXswRkXd7Q7WSuhf05cKt0mxoC0Syc6V4o8zMFmQXN4vAnoPDROwR8tc
ZiRXK4GRbHTgDlEHVPKzpsebJjhDwF7NbI+3UQvHjMk6dks/DFxSCUaJFpMFABTC
AlxqBDq6nAsKHtDsuxmODp1Wa9IDnb9RUPuAmMBn5lUOY+3bLxKCqMYOMyko9wm4
2Iol57EQHYTREtkKytGNOmoCC5o9AvIl2v82//+Uz2SU58wwDMb3mw2skw/xM2Hv
xnw59DD3S0OaxSSBnrKU5lG1XGvJShVhPPB4wTtXLUOdFs5Z3IbPJNEzHoKNl1RM
PypX/IWArVbNrvl/alx4LWCZHEUDNm08fqOY9NYEyJcb0kNmAYy9TQgz3QB/S2bu
KNwdI/v4gY+GK6FXILEJhWa+2oOfrZMCcahMtFowSZAgEWXmPuCc8WBUg6KsIaXJ
U8hiAFV2DJOW/eVLCRWeikKxz9pyBMcpxjKqxMZ2Ozj44Z5fSxUJNgZ1Z3NZiCc1
x1UrC94PkH6ooWvj0v8MZgYKgRs4xxWFVWQAkiuXwzh8x3UklEr8p/V89pEGORW0
Lmqa083RrBBcNjmr9TjmGNpqCsldtQPMS7CfjZ7jgv3LIffnBoq95LwvyOHTuxZa
fu680mP4aF9UvG72tF2p1jPxmRjOPZh72JdfPiVnSaE+PbWx61mPzFeKXuhcUStn
1wUKt5kVG6foYjd1EC3bn7W5bQRpZdNGJNXOrwoYtTtlqwIvOraRmTV8v7Pr4rES
sv1RR/shcsCog9p1Uu8bSIz9wBnYXh+fvMF70FSo6LU/wTTaRm5m7qgNJKAyv5uh
wNkX8uQPjUaIQJgKkjvmC/sbSlj9qORti0+5cE9LVchwSZqqgaRMFX6psHffurX2
bza464SdNX/GPJthjv2GCLmMKazyERWM+yRCAQSpEchcyxJb/7ziZAycRAxm5VVF
eO2vTVRR0mgnJVMDbixHME3uKZKmMNV4OqQAdwwQXfqzCcLv0li/HJXj3uYn6g3c
It9nZVd5959fTy2NrMq2wEQ0IupZ1KU9q2CPksc2Oylwjq7hMdOzgE8qF5pEVkr5
UR0ZE8vQJ6ixkEHSVowx/UnyFMKFDVzxhQP21Ldca8JNgi8Xz1WwwTkimrev2SgV
WUpMOBy7PgX8ur4cyE8Lu6lrSCF9U5FmYY+xxMGyG6QNLrfAxJsqyz+inAuLcTMd
7OGLhN6Y2BOaUyChbFNd3UxchTj/2rPCfmvflWGqBd7bwV5Ng/rGMAKtknxVcZzi
vV3/lYqr6PUI9oSMetXSHpQSpXU2IxZ1hXN48KXHYpBh1f49QNAlWXxJQtdDzSnu
7Ys04nliir0ub5s56c6LgI8B8WNxjbx/3Rrot1Uaajq5NJQnE1Qp0GU97nIn7gkC
yYU5KXV3VfResOnK1ORvXqGgfjkPgB57MtLGmcGfC3PRhA6rcB59awrWHkHkAg80
XA8O7GI+2V4DmOqzdyY+n1u38Jm5XJsOJXusdxbQJN13Publ1OIXgnLbjLQ7M5OQ
ja9Vyxv9/RmCgoDh3HrBlxTdoFCfwUW0R9Rmq1CkPLrk9Gafsp/AKosZwPBW92eC
XBOim649ZXMlNefSKx17hgrqdVw2gej/XVFUgXfQO1EKGXRIPaTENiKjvJDzEoc8
ZRcGaC+4Y3EVNyJcKvTs0g0GrGbpnNgupPswJ8OJjxlOPttZvCa84y3rrjL7v8zH
0shRaOw0LuVEYGOov4mE/ul4GJ8N7mBBkyOFEbiGmKBnMovZ75l89reiUk0u0YvW
KYWSZTOuNsI7gd/6yPadn6FhYM3LuAgoWgnibROJpHvF33d9cc/keqzgwfMfvrX+
lULcMq82ftofB9W2SbWGTYDur0DbqoU7tDiyIAsQ1082JIt/7ghSbvApP9yiK2xN
jVqAhFpwtz/4Z/yGDov3XYPZlj7B7iD/UQ1/nbdgEs6yvhN2Zhq5curyW9StW8tz
nJzGmu5YGYSIY3Lk1MXNeleNFYXWLRT8VZAIPCDP9rlEes0D6d4BPYR2SLw4F4t+
/TWSRoR+Gtp51Gb6gfO5WHX56YIggkwHZaimWcQy/3R4XX+bIf8coJe3ye8qe9Fj
0IJZkjef60p5qVMkBqpD+Xl48oPHuw+tw9eF0cBrmEFBL0raj6BBkHyNnaYFIN2h
m0BwECcTBKvsK4tl8CS+9AkY9VfDxqdVqIYQLQBQ3kc8xNoNZA97xjFzeIxFYx7K
MCfy0rMBbFIMcrTIYQSljMmL5VHWWKvvtM8tPl/Dw2hQuB2dNulX4ls3eNsPfslw
EN2cA8X4RWrz7sLH53uxfEtMWcuxfmbFi0mFxv7LnHSgRAgMfaNQJUsHk47kR0r+
cM8VRDMNOlHcBv1mhitxz6VtFzR5Sc05OrwLIMOdEouKdj22ZmAM9m2pqU9N605d
4G5IlrpGxofUkjSX4CA6I1/yq7G0b4RarxbEFiI+7nkENCNTlLR4P9YGaqRWI742
AeggZvpqQ4HzajFzZh1y1f8ohGxnsFGb5yR8ffVZll4yMN885OJy3z+6X8nnImPg
tVLflOtF1cXap3XSICDsjN17BD3u4YWVJWP26Kdw+QIrHWQrus3GkWqJniWol32Q
sQ56jXXheXAsJ7BvUC1+JLDiOokxg9kTkf81HvYtsbn04UNRFu+H7VVsn6hr69PE
TnrlKovHrNqHsjqpQk+IY6dqECLlE2Vyp/BMep7e4nGW270SosM5AApTwEiPsZWB
uYysa0uxFlj+H3aJdSFhmsmJPv5ubzGdB7fLBpCk31d7XCeD8lgagTokcdXPLmWM
kIhcY4WYPLO6ItVGJZ7blPwYm69FQxdmJyP2IQ8YWwIpjxGtNIvOQM5AGmGjMFDp
QBujFSjngXJwSZmWyyHL/QtEXPQXdUPwly7xPs0ICYVvMSnv/tTsTKtgwRi9Z4H3
/rDuYoori+KJlKorWdP+cu4FNeomFpQJPXIm2G3k/5VnBWJtg/DNX6zWxngSkMhq
REFRH/nAi0KReMzFHNSxexZgpgvjf/neuhk+pMMWOp1vKN0Dgk3PYSqKeyB15sFN
DUc84FbqDr/pQf53m3kdqTZzR67jYig6lkV1Rf4DqpuD/DhYKfxO2c6SNmO9T2QI
4v5BjYyBj+TncVG0i4vmSU53j2K/9wN2955734H+5W2jydVl/qxHHyyFLU56P6HI
j1drbIrbDwszy7AvYKus4BR8Xgu7TwRsArn5jPkZG4ig84c8kiEWM2v3KZ4gfKfe
I8J5Aup+WDZbN7ek/+uGwM3lgKAuroEmG5+mFeQuKN97mARmj7THMRoh+PQ3G9hu
A/u+g9J/L6CY5yLjSwXh0y9TmraD04Pkxea7Bor4pjlhGQyQ9QfXeovQKJ4N/pP2
2WXCY5C2fotGk3NFNpYUo+LphOH3wIvHILmDMe7+Olbs+TMQnlufzRzs6nJkhT6e
DwaR8DirYp8f+yh/43NcxToNXM5jQQc2dWLAPK8/ZscEE0bUDZMV5MitUP2B4y4l
7dlywEcz1BXwFx2UyBqdipMNbP+8gGDQ91UPZcS05Kqv9a57OJFSZkVgk9Ersvr5
f1XxqzbOIJ8ufvplF2RdFd47q1k1zJyeFUN4wE4e0tNYRqbFcRh2d/FecVurFeJY
TmblBWrbCS8C24JCyoz/ZHSEv1FbNewZ+TV9LQ3jBymbz35k3w5oVBB1EFSlGGQL
fcUzKeTb+vFwpAQbJowNQ1Kh+w/dzMrInlJl0LmmvYw22M5Xcj7XliMV3pvUKlen
mRKlNTgeRcRsWg4e7IXz2czbTwIJlCcyL9M1FVG7tLAbYufJJ4sK+dySBRKVBN12
Qg/1GKV852cHyrmLdinxuzNLlMxclY+kHjAriXnNXtrehtxlZ2X/+cRvI3ItVUUY
Iz1GKRS3nW4Z61UWMmltRORQEuGnjoeSCXHfqgZ6R68mmi0q3A3vFq42JmYyYJo7
HRaY79CoNmfC851v/Pa8PjbzQw/ijGnNJSuWliYmVOjc9cHth1gF2xLARWtIg1i9
Iie73vsXAlJ2OcQltw8ACYJezzIb5So3JRCr9UAGju3DKAJXEByM0y3+m9BcRG5J
ZCoeIEgjaPgbv0Pm4Kk1Br4uIXwQZis+pCXYsukJ5RH+PERFwc+EmpaP/MPJQiCB
IlJxCwYuFx9CLubG+1XXlRJgwQCH7Eal9Ww1WN+V3DhXGQuKdb7WWucFsijZaiGb
zIUh7o1bDgsjOZxQrZ8SAe6m0LjfNd+3gxIzOYpPU6cvYXh/OjRAL1RX76/4qIfx
akPqzKfgZkmlurwkAuzozDJnEcXhWHwZM6CsvN6qI8ZdWpCLlCbwPTzzfdDKrtih
ujs+DmgHQ01CzIdByRmyESeb7/JARt3nz+8rBD4N6aoKnhjBkf9BGFa3ojxeNYep
eTCu76wCdiHeaBGzkquohD2cs7oVpghOHWOZlu4l4NgVoPBjj/XGHxPeTOCKZlxt
2PDmiwmmg0WhwZw5O7Q2aHKZa74MGeVJbtHIRHyu4Rpg4WAvw4gvZ9biWHFJDQhT
DE+J8xpS2ccOb8V9fL59bU5K3fz1WRPGj958itlyrAcVCOs2JvisKtQwFnq1Q5fW
JvIqNx5f7o9Fnf7E/F3+yjGhtyV87i7go6ybNN0u9Jt7NSjaF4dOfw43+qKbL5H+
bEJpF3XI+Rz7UQDYDSseiEw0uNriyhRFd3+XxOtUYlpitHsLpiKoJpDDb2tkfpIq
23jZG/hT5Sub4rrkSK239wAhprJsFP/EoVueayFpbEjd4FgJKSkulw/hmvannAGG
Mrz6thZ09HBzEPy5YpK27gEujLSmQTRZ//qCcgTk5rj5n5w0K9Z7gaJDzQxbOuDq
rJUcBBcF222rZ9+i1q+BgrQgr6YFSR+6/JbPhHBgjO1m6+gZxgIP/z/KkVCUe317
cL270d2i1fRQUNOSSCcl9LVDsowUGs61kOBdK7zbPo8=
`pragma protect end_protected
