// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
s86PnTQ/O6E+YEBP3vacSap63HrAWkwllT6DIymjqRNUhxtn37iAC8biuwZuxgwn
MYYCtsypKMSllHkSqhk9cBfTlk3X888p95/oYgo2OfNyW8Ztxh9TL+RJAyqEL193
+hiAyERaAwVGPg/JypUSJm9oxrjDf1gIuMuFUtqs60w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 180896)
Fi5q8dtsnIwisAFxAySPdkhN3oXamopKVlXM0ToqpT2DJ/oQl+m1/g2HaX+b/jPs
xgH/0FHmpyHPYXk6RsMXeKKH79PvditiKNSLu6n0bFwbdwD/7clKU9KncW/nkHz7
WWV4+RaZO5z+IzbZ1jIjyq3SRLC9SLujnLk9mm0jcl4ZqNe63C9ifaBc1GV3uPbB
t5oozvCeHyS9xCdiBZF9Iydzfa3g3vnuYb5R1K27HkMvY7o6NneZfInfjZIIsKFe
2lg2XChVoQ3XiO67+UsUB8QWQdX4tSE6oHSmpbFo10yn7tzjTMoG6dMDcFlEZkXc
DIkScdS3sJ34fCD30r2KBvOoO+3SdomQS2hlC0Q7wu9KTEinvIj2rfH/GYUt5RZX
O4cdjZp4f4kKgMxzluaz3Kn9S/rcfUt6ES+GqGaT12oicryT6lhKEkUKep1mc1Iq
1InPikISKQo5YIGrymc/n3BMEwUeIdnix+w2iIT1lpBfWs+09ObIL5evvDMXhFKZ
pIwXOUXgPqZMAlUWOnP71qLe085rut/EDj7qiZKwsqsWnxH/l867Ldbx9+wsyFo3
g8HHJ7yLYyEQ7No1Ne4+JUxW8dC2B4sn60cEb5EkGHtCosm7NABzmdkXVGeRrCE4
k8oFdKTgCrXwm0IBcyDetfAHe5HeOG8w/Tvv1d6EpcR8hvlaoNPXp9xAStZEd5uU
C56wg1QAD8vn9dv+k3H4w8DEBhmd3sNx3LtdMPzyVIJa+rZpdEGxJAl/ONKy+4g4
eDOZ7wFQK5bpRdVKOER2WtO6HVAolOU2QEw28dqp6+okNEz5vWJqtimlA0fDTZ3c
/0I74D+OdP+qaWrHxOi4RHHRdXNwFqq6r5acXDl2mQrDa9CKMLkaQWyAwMWgXBKK
OtvTkc5YRHHUVO9LciHEJmvYSdbjRtAKDAwhYPIPS+cnaXYmJH225/Cp0G9/jsTv
rjrID3S3alggOOrNeK8d+STwCCkpnQAdRXfW/ox+6Ks+ddQ0bVFJjWM1paFI/ZBv
iI/lUaQ5pAvK3V6QNPfC3MsNEueN66dkB9FC+E1cHBmRDwN38NL22K8KZ9cIlCbu
cKwOuZEWuFn11XUKdSarqFwzSDZG8x+l7PcAh0qMErLHtBHQaKEv1JVTTtW/gutP
aqENYWgkGbPptYIqxcbBsQb+L0jJCNrw3Nkep2Zz6zBnsGKa1C6xXqYEcEMUZNRe
gPJgmjXxtAqYDjUjkpdjiQKGxHS/b2XNmxI7KFFodOjAXACa0476n2gtxcL9OhML
4YPivA+qlBQa8AqP2NEhRB22iDQDsMWdNrYRcial7WWslV/+wU+xihTi4/d4KJO+
irD1PT5WrlFPallIAB2wX6cSlSjrCQDxY7OCCHaSogrdxlca0J7Bq7j861ExZIC2
85wg9sRu3pm5E6pV3bd/FAatz2aiIeYr0RNgtwRbWu+UxJTaJvY0hk3JaEq+ZzsI
4MqMGIf/B8B9aYbJ6lX+yvTZQGzSUKwqPiB9AqW3ZUvtwUviJiLoWK4hCpnT9CFW
lKRJyWMMdwSWBaFqJ6BX7s1KuXHNqeId4wRj6DaMxW75/GzpgANHLw9tTnI2/o/R
pyB4WBiuCm7TY1nqWY5whZuDkovO0dddTkrQVsVghOEMY7jRMw2bq6bpVc0AWGCq
XF8WPROnnwxatH+jPQXLWo27R8YxxRjRpW68xwKjaapoUTgb9eqIBLorOf8N/ES1
pkZCc/z7O+BbWvMruXqzDtROt/1A24ZajhxGQEHSQ2x9nZKoy7HNZQInmIA00GQI
+cNOv17E2qfdmyAVqZTsK5rPihZRSwoe27IkrCz2IKmZrX6SCBDR+PogAj8t1au2
hAnh9CNdkSNMMZVMQFKtkVDmayPx0UPRCM4DAKcrVrk2rm2J9jtBoDiBsx0K4I6f
QX2qfcSbuTVJAxrrxBV+NaWCRZj+lDBNciWdGEAtF3CzIFac08UO+/ftgbeD7PUG
41IaKdmWWsAKirXRwNAwQAnHUkSGO4tWGoCnFOnISKxXpfHV58hHHvG2ORXSBk4U
kFExVwXSsLGlyoXBa7HWaG2ti4VkYCQpP6TXNycIyyllV1mZOp/E+GK6OfHKAqSS
LxW8Dgw+pt71ZagUNCaOlbWURdobByLAoj3hoVAFfxY5nlhMfpPPfUWyvAc7sTU+
eoJGmq/ZyVSCAK8gRfpb2GWokG/7UD3hMyvpvl0DgePUqsJ8OXH+PeyOwwAWjnTK
Z9YtdTDT5GBRTi4h0KHzxhBacKEWpnh9L6jsk4jalV3H5lRsaHyHrs11DVPQfBuI
VkbsE9cmPLu1KUQeVnX8c6ahUlSz9JHY+QsA55Zt09Ptto7lDL9hKBzrLcCD9qGm
XbfwCIyxGlcDoBcCkcQ1rVtJfz6yGuuSxMJkuPbDckPnzPcJWv9Q4wT+xMuC6NS7
8CKUW88axmXvRU7/cZJtPdCmNZ0V7pQAJKRB3tnrfvAikAPLIKF1QWIpZ006/sQr
xNIXIMXssa01xN2/quNuuR7kmgMHPaGM+nuniAHgsX4vwVuyrYcRk14y3S/JvO/F
lUXZrUO6DqclGAN3wxqOODEOG1HiMGwkNZBFDwNdpMlt+I1KOFBL/m2KXtk5VwUp
j43zcFht6tMRSOqY0munvAkaxaBzlnSHIV5rVZ8/Ft2BQqvuav+I6J8ExUqN0VSB
+SIqGFqTdvH0QqZIqLTq7PgUk/n1oDTfecs+BAgQDQ0WfDva6TwFcyXOcJFinWAb
9jinIQnUwSjM6R1fAI2KT2dcin6Ytj5WZdOezPm0fn95QMD+qTDGR9zKnnRMeyu+
AT4wHkfkQrz9MDH6WwtLWx49iWtNrlO9j//UHtrUp8evVND3sjxU0A+R4YTSaTKw
RSM+Xd1lOJj/Xu2VtueCznkk220N1UYoZaBKU974jhozMN2ckjgnZuj0AqiGBeHm
dJFejLuZlhz0h8GwVj9darDnJ1H8GDqDy+3FYic63iYac66ht16ppCA4AFpJao3G
1QnZMt2xeGHo6MAffD7ZyzTwTeN7YBoPK7FaghVcXitQt4juE+hEwSDEx6DoNE+9
qt77LYLs6lXJ9G4ClMI7q82J8EjufBgkQXNszcjqI+llG4r5ZlndE1gAUDr4Iq45
YalX0t4FVO+YAvKwfAFTUL//H2Aat9CByiiIDHUd6ieWRlMZcHDEJYgwM0TOrfuc
OpGzobvJCAn8R/vMSrbFb+IloRTwLtLAMe9oqLJ26Ex6EYOSW14txlYmSlnw5M0j
mKCXT8jZ2O9+K0P0hcgClUHU1PkrQnO/rcIDlesmWPB8L7GA76yN4m8HkN5WN/+h
cdb7PMlXCSQlGR39QfohveJUOFJN2hikmB1xwZGY94CzLUOIuLZdMKqWIlye2N1O
7PayODCMU5dDFjVWiIu63N/TgigEq9+UHL5bQBZASzAhL6LLDBiFYSocj0WKJN7B
5FYkMX9R++odBiveN9lrMAO3li/3FXN23JlW6wYAciFsGFHqnNWoJ1dbd/CY4hfi
U5jCisVlDFgM0cXzQd0j4b4Nq6IHMG0bQ8IbplaLkNXHI1T5wXxnpd8jYGizacp0
AC9XXXbSuxSpahS4iq2j2nNst/kleiaxYYsnIqX6jmKbadZ+l7phj3DV95tIPUPs
JSmIPRYOqM8x6SjrEGCzjN6b1gBX08/SWB8mp9Tk69ECRagqTkTAlJuez1OMa8kB
lTh3oDjkH+l+wT3a+pAe8P7JPan01nAy7AshBIj40oWjpOU9yrxr0h6YfchSPNqR
g4jiOA4koXdTixIHPZ9hHu7iuSV2Tu/HqUi/tVwzSRkNXg/JWHp1BwTnR7wBOVqA
LaUNv+1SPmodnm4ZDfRMvk0LkU+83uQxSkTCkYw+kZbWMxIlKpOtPMb5Q8ertxIa
0YD0NBLvVUl+wm9B02/1/pzYHsFmMPLsINR32Ua6fZyVTwPWpqzEFG9VUTZBljVG
5YtKrHmMPtrqF1fPqCynREDX+zQUAZu4q3NQw+oUEwEzvPVedTIYCyw7hn8VBrRY
LEwzq3sADkSE4nCHqoXqW2UzPZ+5kQcHnPpootBtRxeRVuTwaNtahcK0im/xACIn
Xl209c8QzNip6PCRW2d7kT+/XYBmGqMaC2BnLhwT8BqTvUv9Er1me/TKMfBOI2Im
X/Qz1J07TGPCzmghDXvlCmu0nxpX5U+g1q1k6C6MIHTM9T9hDWowjQPzbRtVAYJ5
u9h9gUgd+ijzQV5PBTuzi81thz0CC7EVgphFL0o4AoAp96sycAB84AFksiwezC0t
/b2/rFBL4/pr3TuHOOWmBojJM0f3fZii3VPwW4nMRrdqkP4i72ZVwohouPEx8pqU
dsrLUIHYP9xNrczMHxvK6c0rjBd5ByFiTv96OltXKcEDtAXIRxHzhloitH/GRsqI
Aq92Ug9Lcf5nRt7O5pksCJijD2S0qV2/Q4NSCGr3hUUroiVcaF0C7d+mj4kCXtJN
vqGrbgp6LTYkO7a8Jy4nNlmj2vnyEckrBuS0MJGonbedtphcUoTBX1xidJAeIhU0
os4czaivxizJkYRIFlzx8E7/5N3JUFwbstJP/qMv2Rw6W+maiwxzsg8W16At2IKK
jrsE2yjsFR3dJsLjFcZeXmIAonUQEdkRvhXSp0qvmUVnFgLOnkUkze+FYdbzVQ0g
Y+1UoXZqYOrGc+ejjdkJArYpZGEEcIEkk0EGw6hH2tk6Z3TfzlNnBc5KUinuZO/o
rFl4uSB9jxlhaN6MInarbFKaXSYvh9nnnEozQ4q4OdEiTXD+Ly8kaCVSeWWLlmvQ
uIz+B1vLvMPQrXeCD+/QCEXjX3Z5htMEGI6N/nXq1pSoCquV8s49TBCPwkSGvEZg
4Euq4qbQSB+DNaTWTB4fbf4MhGHzOyiTu4U0x+NGLqUrDQRG7KtpeXibQkzAMQoY
diEJ2WQ1H7H1PocI6TNdt34bT/Mw06uvcZPeqRrrDdwc0hv+ml6cB1R88FXrqX2P
9vfaA3kVieuiCNnBIvmeqmW2Qqfx0JXnHFreYwcR+hHZ+YY+mwsjwB2IOBUzJrtR
ippd/ZJCSNQdaJM67oGj/5g9t2BMpTftbdItmFcKDW2ecQ47A4I3/kQriNq5Xonq
44/PjGuhnj0oEzRhGgAe6yq45i84iHTS5490j7v8apkpMX0uyGy7TUdcJB0qd0sV
UL9/M0/xSEzDE2FGJMFUZuWFSzF1SSZV2s/3s2xinGIaUtf/htku/WfBwELqv8O0
LpqVWi+Ypyk6j8HTzAQrBpNYlN5jnVMQcrzjRY+C+DGXIitLsRQ19B00/tmYji9m
HOL7UgcsJxYczW9ybUl083X6Zr8/IU6iO6oxHxUtDeeFgU7zf9HabKM+oZ9W3MHq
BXQ19dVVSqynFVsuT+4GuMKndi5pz0slXdXsCI+CG+/AlEm3JPia5xM91g87b5aa
3nNbZEBbeoYYXHDtb8+xpVh2cQK6Nvw8HqlLCoarf9Bz3JH6IElRxU1Nqr87ppDg
wtw/PXMtDSP1Dz14FtoYrepT2Ct3VvzF+Qvx+unpR3QkW5MFG4Z9m22d98g+2oXR
aq586FqgWgct0nwkGAmBCHjyEiVjUZZgb0HfkWGn5hubP2WCL+uA2XF7LYcxhd+R
4SvWhPv4dBZuT8eQD+H1qH2Cfyi/yffrLcsypTJRYHxXpRWGH17eIS0o/UO1xuux
pXz+fzEIa9BX2v1rCbeBcTjIv0gWOTsjrynACD7RVWKcxIHHPJJWwyo7w/Jgsrck
2XaRUCRhr0jdONlNI8OVnga4rdUwX8xNaEV3W+WBy5JyNhutboTyp7TLdvqyhJz0
z7yX7OWtbHPoYVf4Gt5aIelEJs5AOJQ1zpyWHL41BmmGVdrso6Cd881lhMY4Kqrp
5HA1HzzGh3Y5L2c4f8+ttR7NBP5WkYOw2WadJRdtGzUKyFwLv1zAblvk8HNwee+c
4nmtVbkGerbwMWehHSH6NmU/tR193rPQITIgVfAZJLoxfy58UCXhNYtbB5J/aTVG
2zz5EYdfSNJTwdt8LJNdSOyNFQD6Hn4IZAxxD6Ey9ZJeaaELW45BvuZ9y/PIeY7a
NwyWWn8F4wNmAGGMq/zFtaNEYD1IO4iSOQmc/KtRQcq7AEAmMDrtB8Ed7jJpBEwD
2c6Tk3dGDn4Vipb6uqZvSaLDuOAfv+BmoeqjWG8IoKIdf1OnoZ3P3TXN8RaT8EKA
UaWu+aivwRZ/yDuq5qW2y0HDNmgETtpNnTMm0ObALJMDAHSWY2zI13QyibVkCxac
5yDDhOMIdnLth7387IkzXj0+I4px7DALQmFchS5OCNgmkMv3sriAe0FtdwHQEYum
JtkMcLVK2MJ38NUrHfVGIYpJXsioWmLJM7ggRUQJcItvQKm3/3PY/2BlYdGge2DP
5uw8CBsMnGL2FAqEKPCPeRXGAl48YWoS44uWMdPSfaoyB5171FryTptfKZKkLsvE
TI6iHShN+KP+LFS8CBk0/6yGYBmCWYHBxgm2RmdHGRYMmimjoYgz1aC2OAtHfLbv
YYsREW6Xe6M0QKwIjcYopWQQjN0/FvV8V6KHCQFH0xfNADLXuCD8sQkxFixY4tIX
7MGjl9RU7N9jLi87dChEyyN4F5PhrBowohVylI3vj73gJUhvXl5wZtES5DA7B9uV
pyQk4IPX7JkHTb7yKJseSjz1LfHe5zpo8J57YukwksfwK6YbTTPkvAp4XH9I/03L
FTogvtrZInwJ47lO9sKFWC7lelDsjQYHNp4jALZK7koQ7Jbn8YCcOWhZs7aKSWnQ
5Duli9EfhnoLKaq9uyXP1DZKQfTrDU8uo+r1W6+Pk1Y5HPdEcQmm9jO65C7APxq2
NE7g7c3YdoysuUzz14yh2LE1UmgObskIQlSY+noR6khbyXcXgXR++UqWqQv84CbP
txUi/3Jtg9C61JzpwDr6wqrZmVjhdfrLJumwWZQtHSKCL8yWBJPgbCsOuvRlvuac
yiLp/1oQHAWpr0CyXk05DdY4wak4j2TM7iT4aJIgxvl48f4N70QdmEm0ci/zpfBe
xSq6BLOQQhE0i2qjgag/PfSm28T3Y00+WWjjQHZcnIyWc6+HA9FFitGOnlRDAXkR
mqtY4rd9kClchY3FunKsfPna2//+QPPMsmVLqawJnnBVGsBqLNH56F0H/sarT4Y1
pbsbcyv4YPe6Nou6QBcaGEfThkw5WCjXEz/v8YkEjlfN6fPVOUJJmtCv2Hmo7a7N
djARlGZEi7wvf3g1Ohkit+R5Dcyd28mq7epu3qU5w/NWGtgoAr1/A6hnynvyig89
q9nhD8Vj5uQ3RsTpVk6vfwumuryKEh8+1tyh3JhGRXeEW966Qh1NjXBVVWST/DqU
0TvDtosZ1h9+LH9ZFn0mpHKhKeHuP0/4OsR1GpKzrnisAa/65hyC/p7GZ1tp4mSH
F726cma1NuS/8Cg/hnPypZEk9iJbFXM+n8FNRHe29rNCAp3yk4SN2L2YzbEvcGow
vb0ttC2Qt40iGkrsNmjoki9ivc0w0PBETgPQCf2pIURwnnf8xt4gpyHzAFLqkjhH
zrK6fnIjDa2TognS+VTK039sw4R8UOePMJoE+huSQlhOg3U5xv4YIogek+i/SdJA
6vuQ5/FTrRSB/WBbVaFiXgQazsTEEFF+g2ja680akMYTfUHDTH3bSuyluwdLeKXG
bavnpiOz14lZ7rz3rnbCzIJ6NCQxm/K3w/5dhDOARzXtWi9ie5wNZUqoVqbAMI1f
lfsCASAGncTmtAUqXyijkiIQ9OnIih9CM4UeqoQz1g9mK0J3a/P50F1OeEW+FjfL
YVDAuAwioSNbSFRqC0fv2BEuvszSKD5RypbOxoGveU+UaQzKPQtrEAoYPXZail1l
HeYuV15zPzmlqOIAsfGJEGutOQTO78kYWHRKA6RtrEgWch+ijSIT8af9JKLoi2rA
gRjh31vdmwg5Cp9y9DvgZe4frND5spw1U1BEUpuAN2DzH1zHHtH8+s51ePPKVGEM
WATajQjdbQW+zHHN8AOyWui4K9JOI9wog/RIuXMHghpSoYVAm9lV283z3B3Xyr2G
1gbZaaYxw5MPgt07xxiawfDnZRRGhDVMuF6QR+g1BZND3mLTO0j3vyZCB+V9xpOx
/e7kLVJtkbplEFvmhpR8hGx+5aXKaYfiWFdtuZDcgpl9mG6lZwfJByLzZdJSDHZA
3lGR5feFM3QqDnokE8EKuCP2E/PwFuOvjpQOQoWimRN57AhJf4rKnV0murJ2KiXu
6UqKFGVWcYoGqfEDI426E1MSRLYEEINQJkm8efYTkil362MV9a3jCbTmn0oXaPbV
lniqNTyA7cTxoDMBljeNW4amr5a7RZVHkuD6QOKMgzpVNnXajJA1ZZIvHAxuTAzG
muL479BDJU/fX1izD4GCsi6/MFVcwANONEkuAa736VgXWkcGSnTGYxMVcWUk1Z01
QBuvBOgkwtWZpXW1pAQQtRD1+uM5DxbRTTVwIrksZkg9S0/UnrkwrrwFgKLNibSw
RblfRzMSEsFTQSM6mrLPyRJOEg8oL+Fl4KJuK/BLT75Ak3pRmSNkJRdLHTAEEW0C
5NhXZooaTcqdIRLO9JenAt/4xAjh8hpa4XpL5CQXzAs37xM7e6tAFK7yh4/or52R
l5Y3b88Rd6KaetPCg6GRO9exxM0cNUsO3Cv5Ufk6nx3t4CLEyeS0a6PH9EIElZhm
5a8WsHERe7SufEC4rqTku6iBDNWvv5GupJRWP76TUZfhZtnboUki2MW4SsCwBN3W
snamZHZ4bUfVn9T8L8jRVBv05/FF2nMeSrs6gJa/9/OHaT+rIYC4S1vI06ub86Jd
0FOnSmAU21d5VRGooP/ITBn0heFng0+mVvQ5k/dnusiDLn/Y2oe75lmZtw4Gm22g
do8u8k0owcO2SR7k79qIdcaj4w0LX/9vKe5aEwOdz64qZGu8yQeFgG837fbmxRMl
0EMaI5+pwWoGnCWlerheG/ckkVWBQvICkLzMpHjYUwroOOCMol7t8pEYex4pZ7j2
G9/q3aEuB0uHLLMw0SSgZjjO+HHWh6vUQx9X3jHa+Yegb8IeT32/P8HXXYP1JrXt
X8svLOmFCosHCwFl/gEdgEmaecyifdf7kE91bvR9mU7jRXqJWllf9vNTZqg062bx
GjkWeZvC+kqr2ILNSRP4FFFpVl1h5KIlA+IUsgJsGnO8dDhdKLw3ykr5eRxGcrBZ
n0iI+3agKHLueT/VBVFf24g180ihfQpQ7bkKvfpc5WImKExe+VYLdWkRfG1PK9Wl
i/ZoboWB3IFp20J4D07FrVtYUI9yKS+M2gvWuiCzqzJSucfe8v3xGgRWTsXotyaH
32/+GyRl20KAorApT4xE2fq0WGnN3TifsrB7PULuOU0jlOGzVwH5R7xOev1Ik2m7
7kcapx52Rd4gJOG+YeEAuSfIstR/xTp8sEXTCkQ3RDI4Kwzi+rm+FrSGJqmT4Rtq
2rw9JlMcSZU9EXW+dw0Dds2JcWj7TNpV1YMMfnAbB85IosjsSfqTUdG6DLgS+O03
2ljrcdfKt0j4vtjtWITbPhaEAOW3M4+lCAztJIufoNQkFH09+pGwqgM/pRCEgm+1
8l8yth19AM5G2lk5ke59A8iLT99uDMil7vTqp4oVoe7z6hk/3seoPlHX1S+wZlwo
UtMEaY1t2SOXRY6kIdQDWjR+xiVX3wpcefJlo5CfK6mmQ4cHQhk8890Ci/jQa+zO
AqoJPqbUF7TyTzPMKdrE+NT3difiWDX+zTFsVau76bDyFg3BSQ1IvJSbn7EvCWze
js2zoUor3QF4ZMGNNOcHBH/DOuauvG7SBrl/ogTiBa5Rcfl/808Jhd2is1IxBf1y
mD35pl/LhJM0UB7lGwPGaS7FWtMJiYTERadKnvLXcXcaQFPttBtOfqA2ks/cjBKl
idtjihRMiCcsPX8sJDMPhjcUMWKCe0y6FV8YNmT6fPwSSCNZth7CyGQO3dKcV0ZD
hqGpGpshGxxZVKgxJ92EMGpj/snWP7GXd0jZiqdjgjKw3Y367dpyWl+S0Aw+MZUg
2hdIL4Geflwf4vJPtOdrX7yjEQVrgGBUf9FOMj1rfLZZfbvMyMbkGNLLcLeyw2Dt
DXbFFNHrPUJy3FZfy18+rMOIOTSL7IoaLgoL/5etPEwwOil23GdD+E2Ynl5l/EED
jW5pQKB22VdZRwg/qbHyOg+Uup5xc+lT1tVTztCg0gbApLgnrIQ1GAXDnEo0Bysy
6+Ng6KB9lkAmB+32B7QjTGykuaBV3yqokyKyOlgZxPa6/cEJ57KD54ZG9xGcFsHZ
ImPwb6/NCrRAg9EGHRmXSYlO71QV0yAHsKGhYb5jv3j98DQnmtY1K4BZo34JdQp4
YEM+rGDuI4xy+mlM4Xp2rh1hmsUNyazxEsWlQVXfbFNsMGr7auUnPTG/3bFR3k/H
6B2NZHwYlF4Bbrg3EmrxWLkDEWeAovSSDFR6jYlL06cVYGY4v8tK1YtU8eT3quJt
OZxH1V3drcLbFmh9CbjINc+8mym79saD0nP840Q70x381IygN9TWCK+JBy7nuSjC
OuQsMnVE11PqxqPBaZHjwedhdFCrawXFKTAepv4o8FbA3UFvEKNpiViSTHI3rqTW
SsGnNhn99m6mL4UOEHnzTFNJvyMZcD1NtTNxM4Av9hSCesrC6bMwpGFP3e0KFGfd
jNJuAnjXPc1iOPyW4dXg/JZ2+qlx5m1N7tbqoOXVD7zhEEVYfbSIptCuoZby/9ar
7uMfGBmyYaLRQ3CqOEeW9BlPhIfKyu3UWdhPJC3n1m8UZrz2gesaYI4bPa5gD9IF
RyQsm5GMYytebVjwNxy4Cu8ZjZV7YbdjDrC6scVkI83ft46iQHzPnctwIt9Ir6rh
sWSCvewzz9duh2EWGuvoIfkTBIz9o5C5ARg25hyeqbsLUnZM9BNNKeHBVd+AQFIs
TcjAfPqOpDqwslpr+iYku08max0ENqQ9B35YjLVq6J0T1hBuqHTEEs/5dawHZzyz
yw/snNCnE191hUn+vYaQ/xXgmJsgvkm1ltS9TEiWc6YbRHYhNOj2iLQAscjaB3W5
pMl1T4GrGiT+/+KZGjBe4wfGDSPzFK0+CvMMb/C5QParMLxCI2PfQg7kNAhmhGXt
/mgQgXYtDMXJStQKk7ZpzluBxwEYUKAIUexLMqPHs+BZwkO8H3AONSTY8inPCtva
F3KWgEMNI+9kroXADo0DVa4sOFxZXJvAPJiJe0WdYScQEgV2dJpanXHz5Pk2h3nw
pc/nkFGqVxCPmdp3JBFto8Gou3PCTj2Qrip3W1+rgul0ngPmYQy9NRrKcBmBMHVn
AZj6vNmowCcB1fklxi92Q9K71rkpy3asYXWnI+RNJWPBpmkMOHJP1tnj/wSPAMuf
fAV4LmQw3562REfBHCKK6wYNTSV58gcFw+ehsfJcahLkRtZhWvU4ZimqS2Pad6N0
Y/a0jz4HBSnwRPU9wUetW24k3ta5xCD6CNwWozfHtlcf2AKP7b64QGaQzuQ0j/Ol
O6wBJc9Bowfx9k2py7JxUmcSMjzjOevaJUJQ+uqJcHJ1f/MR79+D1CwuaPWfkrMW
vJHuZyf5zHI08d28epGtiE/BCcMRGlFzFKDdZCXP1cQ5IyyRWJJvCy8xx/mvDHZ4
lnNTdhBlDaMtyhV57N7dfRBIzBheP9VHplydO7mPGkv5+UHMdE+IoZk1kImQ8xIO
jiG3m08IIQ8PdXbWKCHkqBwx0z8BR2rN7PTOtLcabz1/3km29AQqGqJGaIr7sMeX
kvOlYtNmFyHf5gtswhGcHm4/3qbcxFhU3cidgFPMdVA91ofUDzJ5dKOzBKssnQ+t
+Wsz5fvX47qwxNhIyHBqs18jKnYU5viaPDZBILVVooO7vf2jJFfVRVq9IknhOqEG
/F9hBfEKddbDPvJioZFWbYiVKjEq/f/3YpyVnklcB2o+kTm7NdxkoKQyz6dY/1gC
Abk4WLRj6C53avGHjF3V2v7Ulf9+yMArh0/N+gx1p+LNlkydY97NHafuEL9pmAGM
lYdrbEAR3W5DvTxwkwRzBBP7NqlnFbfHvv/r6KO5apoooic/vpsJWI8cDSwyXuze
M0m0EIvt3MIUkUltPOkFmVwJEaigYWo/csAjwDLxtchfeSy/1QKMwDyxYgVAcyTR
xOE9INIFPVr7+JPu3tSZ/QGUai6+qejB8QgccTxuFlvcZ4WNY+WZeAk0EqzeDDUr
hBtepc5XaDfS2Ntwq1Zu11w7l5u4Wdu81kp3+YCJp9eIvXF5CZn/6x7CcauG+zfi
q+CVWcRe04PDzC727VHN4+633p+f+hCzLSiDgTip2X2+xqBUvtltqzN1ZW8HDw8g
HSvlgl+6P4F8iZ1R1M8ltQ7EvhNZz8WQRbNZc0gzFcZgIvzUMHvtPM6LChmbIrNQ
N9Sen686Ymho7TGMtPrpdmrHmNVnfzpYy8ti1xNFOUzr0J/bul34uRoYJXVxuTmo
9CzyKbtEw9TTRDfWmhdB3ZsXOUdAho0/I4rf29PcM1cQzyoiXBBrtcspvcr/K8EY
p3wbmsoDMP0ijfdZv9bFley8vK0Miv0uPpY5mbH/LK56QFCh00b4EQaLWQ1GGm9x
59gbmW30ZPUB8ZEy854hqLuwIm3+IUttGMYgYRY3N1GHoN/woUtRRQG2x8ab+gjC
rFEaqn/TtGtYjNcSW1LccI5cwwwiyIo1ZjyIVNpILN6cMsmZGr5EzdOuf2eelZhs
+NBv9xUmSLj226Z3qcBw1e1tXfVnS4A7UVC3PIRsupEaquXI0ALTWfZnNRPWzcOr
Q3gzlTGgb1pMKqfahzjqpYANnFM9ytacu88y02TiOranPzSdrodeVturDPef08yG
bHfwCowzGiDBrOdT0EY92NjtMH9+rZm13UH8YGoQau19VhEv7Ea5i1OL9WW/4q3x
YXbJcWjbYRmsKxwm9ElVsq0FzR8Qqytr41Lfw5dx8k1gSXDjRN9+pQl83OOIfrAE
P0fL/lEVtjjb6IkVO1Qdo618cbe6ToiQzApnVcW2zJsQXMjr2gIHu9/cQ70Rv8Iy
NwvJMk1b74L6rFm7JcZZ1/rKhca7xU9MUtv9xvqdbMr2K9gbdGmLrY0uoP9DJDgX
Uafhtft8V2AIEhES0hkH5xSDKmyEiTxRRfIP9Ak61EYnfNhqHL+tugBI/D8G4NbB
AaWTNgPiEtcaxdEmekkZRJ5tZpvC+g/yMvgKPv3nW6v1N3cSGByWv0mb1nileGTC
QssabBn4NgKZnvZ2CAGFl/d2td1wLtUOsdbz9EYVvV3TAp4wkG2adDFrMiX0UQzM
hpWpqhaavhQNRZ/DaXxH/jhbTLdheKeJuuHR63XmNkriyxWv954RH9EP4xJgBe83
bApFGZEEDmCK3d6a6i6qu4krgpSBLMxabylJwBmdiP2eoN7OJ2rBYHDl8CrE3Rwz
ht7bUAt4YaNDD6OEMr3VPKPmaJBX1uldFdGefqbBpXGZlP8oMjL5fTBR3E4Aqu3w
zxT7YbGibM+boIqGzthXl9jsUwzog4LErZYaDMZ3O/xJ+E1GspTVbnSB+C6vic7+
+mmYPtioA/FLkjjh7ad4Glx7CCna0iS0q2wG9biSwjXoPeYM1e9pFeUg8Mj+2ZhC
7QCqnyFgQwveHnFxf/qjLFuzVZ5dkWXPZYw2T1pGZE3Klrl6UhxmxdRdyCCvbTr1
uqz2a4yMklE8qxNBdqFocbPs0v0xt0RXfNY5uRgkKT+FJTQ185Ml4rj5mJ66nzY4
krsIwIaaN5gWWUb7EtopPw9mxIZyRAe9Wzk2muuVGGXv8q5iFWgzR4gLeB+2sRDW
SS1J3PWpzHbxZ6q2SqaejHhIV8oDIBo5m7WbIcrvWDlci4UuJC4ZRdIK8V2cTY7W
KA91wov0qKeMpEOG0SFAsfyIuTKVV+afSB4P4bs2Nb5yPka6tuG+h0T5cVAcC7OZ
QE8FPnVvWBuBtOgQZ+laYLGK9U5X+4CWwL6spByAjwUYesZWW2GSgIB9qU4ShrQJ
m8o3paBvybucHXqTjzy9AFaFKEtFMwjS+2Kqq7v1FIV3XCxZ8PIq5R5pMNl3kC/D
jybSsJFT7Axc9jraA/ZTGSdTgzRTHWlNJRpO7X0xSlDzbAVOkbvGVzW4QzGzjWB+
gm8FHSOoH8jtM+sZqZfeO2QlqIxcC+Qs2/vs6BuS2ICIWjZ+g/V+3suQaCjIFvPp
Z7bydkR3C6tXq486Atw9/1+XF/EuYTioYURjTa0DBpWXuAkU7TTAkCfJ48tjdlan
3Li7HWflGG7NO31J0/VYi1uDzpEf6jMBmhCBhVca4p0ECZahmgiaF/545cFRGJTc
WalMiCjKIMpNXHWP4oMoKod5xjbf9TAkYbUXRN2J4hbZKKHPGPNtIFx9fPSL/Lbe
HwOPgE5nd3deBV/UL011lfZgLmhNsZ37PO8S50e4CP7aC+nVeboFILBPIU7Dk7vF
cb1SHxr+tjo2jHR4/l9V/ViP1fMffVTbV+dsa4tpxEeDtKw8FbMA/dE2P3mcM0vL
r5J/xCd39YM75sP0TTNCM9+Ea5aUhFytqF/6gjP9mKuQDxR1Fm5ZPuISMc94EEZW
1IjZJDVJHViRod8H0pGeaeT0H1VPohug0JrRNJ5m7E0jzLGBgvAhb/Ph1u7Q4zj9
WrkOmpZXVnKpc2DGY19B9lLX2IivZxZAnPcGX0c/UKGh89BYFaomWPxjA9BZCbqP
7QK7k2zssXouHw4xIPE6deH+aEpw3ZRE/7LDItQL5bt+ZV0ymfo6wgQpcGx1/Nl7
nD7yxSJsYh1CM7ozvnBKUAaGrNo4J8rxlCjzto74KTr9QNoMgZwgGKBpBNqBJCrw
9dVYcfnoLWGpLkA0nF/PYpnIg4QUwvdPO3RMvoCF/d8pc2DDIwemsg3umfidH0jX
YGxs5oy7/PYTyXlauK3RZF0W+3l7SWo2OLQ1K9Pp8edpZAYqhBNuqSxS4rRbYPBS
6TcHeWvY6c3W9XKIOSvsC1yfxTxCGxGjsZ/FKpc5Ev94lhm7lthVrvwBQ6o8N4GP
G6Tz7i/4o6UyUxq2q/NyC0agkOe94VO+PwE7AWQFl7tAx2gZoAk3wZWe2c4iuzSo
q3M99QDc6d0u2qhKWuSQkXGqYCCDC6rpctx32l5tcEDPZ4a72vs+ZyxwAop9W+Ne
sfyZrurE3/HbqkC6S24Xy/3CDuPUyXZxiFrw4+Vd6A9HC3ANV0Mw1kCmKgQO+HML
jvrl7cwMEtIniCz/JqOdEhtzmZwBTNCD0zTK4n11ZeFMVngNAaaozib5Uyof5lIL
yyX9IOAtcwoaogwPqP/8VpdWydpNTXI5Rk2SwY4cMTW+OoWLvTPyWMkwlQHZ6+WU
skdosC0z5+YFON5/a9H3xlf/So9tfAC89ocOnfd+6hD4yOhCWUp4SJGvT0SS7Sdh
kWSGetMgAU9jsp2pOa/1lUyGpLF3JuXq5LVS1e6tMsNIceAaFn7eniytjHdm0n2L
SX//7dJjOpjPg+0hswjJxFQ2Z2KIiXLkp9PmQggmakjDIBecncYsII/TxSSe3E/I
Ijg3Ji7dE0bi1lukS0HMkfO+WidJoQBn4mc0ZDSYSLReJBHJPVkwIQpYaEfrCly/
haAd5VkT8pjD2fNWTp2ZT0DORS8JNEYukmvI2c7xaRUKWBmvSsds3iH4KPk0jKcY
ZY4+01E5+QF66/czG/5Ak8hadmDtWRTSese21jmLYB8Bdk0ZzrQlTya6Ip2LfJjx
s/cDcVWSXAzQOlkr3tgabRrXmneH0gdHhRkguuIg7hdghmUqItfXj5qXVz90s8CT
X+rq2mmbBdgV5RtUKAGu4/9hX1GD64ce/MKGelUzghsT1X1G9GXinYbwc+zk5O/Q
qi4toq5F0nseSOvLkWDNEgP+KEzXVRkxd14SrCo+nPDvme11shnQM3eBkID9yZwr
F867IW0mRMmzpaDXDU85rUJNHlv2KDs+CNviK/ImSU8yygtvgfvzsE7zeacrfiyZ
jYKUyxBpbOYTzDlGovE07jO50L1Pi2fP5BD0aqkpbTqhnHG9kc0OEwQet3K1HQaL
r97NiXo+WKyaAvkf6l/xDJAF4tgJBLQcKBpu1QPCXKXQ0VepNfxn3s1yaZWkwok+
24Lsvr2N+IeBvP8X9kEYbhX3vMu3CaZ3GcNLXs+0e2NNkwUgkTRgHUjuI+58Bs/W
SpZrJpxD4hbg4MU0Q4tTKPfbRgkwBAjG99ic6hwvLU+uXJQ81nzMKXVuwMIasGRT
amAj/2TgC2v3ZNho8P3fahsYa93kBqKfMbeF3IWjzSFMVpkj6e9w128kFOjcr8hj
4Jq3TZCID004qQlkZULSBKYwEZ0GOxJDnrTVgllZSYGI8tv9SM+W8f86+CSjJL83
rdmo15qmvXZjtQp6f6FVsHuIQlXZGZL7BxG+Pe5ASFkVWdl2Sh/SjaXmH97XGcWD
7d2yhKgh0AxYa5urimyz5O1rEehb4zTH2I1V3Oe1NFLO8XDGhfMok5lOrrSuI5dk
IO1S+1EWj+yLoGszbmAj5rAprLvYxIJW7mEkp/iFisAfvnZlzIxVJFZpocjz+ZB3
r+Cyqrs7toe00ThLO0SsMg3ifF/PjkWNLnwXL+oT2zd9i8cB+JFVVZTphLpmNFkw
UutBmOHqcVOe1GEAWy69tXqpxctxWzqv8jR12LHtvj7bPdogWOXe9PUDHct6YeXz
iWEgWuphzht41uOENK4iAhpl/PPPwxxpreu1ZozCAQ8an97J558bQjC+Fj7VBMUW
FnQUK4ESpHLiLiHEqrF5kJmTpejszhxzpkLLFrS+8X7RAEGjH0noWH98AX12TQ4X
zKSZVuxpG8qJkIBg/lT93JaDa3WKFBo07zlo4OM2FRQd4W43FTAYHwgd/W+waOEP
MaDEutHSjOUlXXCgLqn5hUUdznIEYri0sUTfa8u4LMKL23qD9XWZg+sZAUM0NZ+E
/BrAb6jL2D+K4+UvYa2rW00naUw/L3ozJWTtjQpGqmSlatHi5HhxLOkwDrxkWQhq
zrqI4b9I9F2rzOmlTUi78d6o/qSxXHZ5R8I762EsTnsDjfmCPnZ+3V/vL73x/r0f
R7/U+VkmBnGmnM9TKHh2P0t8DZRHBuJRTP7NI6Fbm0xqfKAwpl2KURSokzC41Ztt
EhZreUy7S1AfdHMM9rSsx6XpGv/K8PEJUDN/DWj+s/Bx0XQqp2LGehcOocTpVMKf
j1rH8axZZRZfF/o1i2nbaaQyL3LDIwkl5XfGiJMwtGCzWzSg5KK7TAlwyHsM282k
EhFKH0w6npZ1ZIRCbcgFS4gqyOlqptpuxUHjXHJeyX31YoiBzkOw+S05ivkVkEXr
daO04O70hnh4C+5bmwjoROtm2OGwRxixNQg8G6riFsxwVuHS/2dMpG0+Z8QYNrWo
4Ilm9R4rxpTmjWm+2CDoP4ibxncnDbcJTe90AOTphbmIj1Zgt6Q5NrKqruaImbDF
TOoShimn7T01MMqJ8Po0MgGLTz7FMGK9/IVZ/H4Mpl/35G5ABNo/dKRHt5yNAEoO
2ilor8f0aa8+cxF0lcm2WuICDClS9RWYhWuip2aS+Utdvk6eCjDBcya0b+tgybrj
lzOEN2VJV81HBlQtEvrCkVkWIhwbSvT2PJnwOG8ZJ3YJpPzfHkBwwvtUj3dQQQB5
EKBS3ZTjm/12Zy6wLygr1dzJCQOwMEfvCY4afgz5rDKghW0+Vatwz1TM6tyfwAo4
bMZPEBnLLzbiZ+0JtslQ/iaGaKsbPyzVKcbga5kSdu1xqdYkvWuMt+N4pRipLV6A
0pPZyQV8ElAkslBPtYgxUWloBEeT0HVWvP8d3lr4thIoZh2OZVZBnqh0JbFRh3pn
v6a5WbYgr5iLTT9IYaGi23AyUtd0DT4d5I/o7l2v48t+LECkvvpnkIs0yRGTikvl
gQfszKIrGfJfnxqHVmB6PmjWyjGGykkEc9kagYwv/ES1OhzBnqjc0QtLICikUP+s
7LQZb+L8gnNw2YQpUuy3HnGSs1kj7j8KqCGMzo0a83X9mUUeRVdC+62javkKK5P4
HShLwrQvspsv5KAQhGnqJqWc85M+rkEsjzod7xqfm4zFtfgs5UdOFksjGdMeeBCw
iOqcGekeZipByXMiywhrToijpaJts8AT+6YXrGP4Up99TDOomGn0QeHUZBgUKmh3
OrvKoFDO7S6Wx+YQoLr5WibJsB1zoWeZyszmZhTTwLL6rc4pi5u121T9XA/qNQzE
clXIXrVMJeMdYUDPueYfc5DQjZn7f1E2JETfRTZyAuI7TTI4R79Fgrz3zh3Huv2A
rPTBckIN+e3TsokGhDMJXt+2UgG7qXImyDrhnFfYUl6qjAvf4//hs7yYn5h7Ue4z
a9mUM2Ds2MNLN+VIgjNRpy1GXnrZOwkrCwF/TRSJiZjIfpNsj2QzSY3oNjcuoeoD
jFu7VpTijILG3KIsqoaVwa9J9mDKf227Xj1OjKTA5hGlZK62nC9yLyqajBrbfmKF
vkiRoA1Oo3zJHs7eHAwncSmtVwSMqU8kwO1M+iAbooatZidPmosIltNXQi0dGMrm
VHIUOrm5JvDF5SwNrBbJJvtf8jPd72E9apyYt/lVE36f5m+oDHmU9F6yr9RI7zLp
XI2xC1n9XrjsQMXJOkweHI2k5zUo7XNavK6rIUIg66Y4qsYQnlAFwmvpPH4CE/eg
UthGkiYuPEOEy0tVOzhI6HFSiPL/no84L8xjKjbSCeihY3+oApYm1kCOsbionmsi
ahzG/VH9rM7ArnPXwDVWuj5S3Uu06CFom+PeqLMqUSdHsI3VV1wlCd6tHhzDcXp7
W7umsH3tK6Al+q7EsvqajzHMZzIqnLmHDTS3rT+nXMe7FV1fWxNEhRQtyEJaDWPX
uLLq+SYwatoYlLkU5GP+gNFOZtz6a/ntuc5zOJUpkhOJUdkwZw/TD4MpwXx6fMZA
ALCjh0rNw5M1HuaoTuly8EeG2cbuLzptnihKT9lPSeuPUHm7MIbVCZz2UwJ90Kk1
C5Hxo1DbInS1C/wGsmdlpPs54TJJhYJvCWDEa//dEH93SgO9DE0NCJIhzBsvYL5T
8awuktG7ftYURBIrV5rV5vT+3GTvff5BpoHohJRJey2TE1WyzHPELqvRRr/pchTR
csaiEAlSTgMFNAk92Q/B20kGPvNLdrOu5LIRgW4hR1tmgsIO9dIOSxyZ2Ut4xRQD
XdhH05pIlByR62VoI6EPt+xdxmd6rbAv61PqKy5WT52Boi1rfX234W6qtZs3n0dZ
IM/sNT3yjHYwHNceMfbZI7Exd2QH5y67mXeZKF4KCRz3LjVj7jXHwsfbwnvLYW/j
ITlgBbY/TQ2YCw9BvxPsZxOEfmaW44VXLzjH4KaRCpsrVS7PTo/rGV9iFrl5Pf/C
73APxQd0MRl6QCxYHtscfeK+JsaPX4dx65c1lc+T8R9XQaul5g+ggMaz0aDS9fp0
pHf4LUKX0mxrz3215D9sjAYEpe8QY2ESByn69LnZbzaPDBg+ryo6RkZV0QcvC9vD
fqwSsvYrRuMVDv7f+kTjslv2FryiJe6J7ism+ZsIF0RiV4WjdwJflbIriEJegMX8
QR4d0ySWMIAPplbkkee3P4ibbG5EOiINxHySSIElnC1qGs15y/BPJ+qWKt3q+sWa
IEcJ9ph+02lSCdmeg8iBaoVEngnJqp0K/YnJrq9HXD3SNVztQWFWhQuVpVSJr2uH
yBOGd5NMzJn7MpVCygxTv5LSqUNfpK3c5F+jSbpJHKZGQKU4TJeH2wpUSwmT3X4a
P6SZyyGgDf4Y0DTcrCvFXmulKOHtyg7CKnkl2XNH77YGO18oKjxErGPIDl7Mo9ll
uTKurfSbNDGTOhrP7Z3NEyiwjRHXo15oPzu0GTK+CLZYT+zScuh424r7b/w/vG7H
TZiyF0jzJZVesuodRpNfaT3ju+p6ECBpjj4te62BKopeWRVBgrLWQ7qW6gt8ZfwK
noQEjwmNfOVdumUIUTcycPAs0oCYKcAXJyZT5WTM54hVg7skUcheOmXaEo/AxDnV
+zBUGn8+42lLH6LUNbojzJlFv/hhIb0p88ubibZHMbe6ZVFJJPsTqoxLQn5dhmlT
9DPEz8z+o2xI3g2t9G28KFQHsvOHVIlEMbPxjm3gsL4BmvAWADZhgeCKJ1xwc5fj
9xgrBHRs5DjN5gVNcM8r8r5l6YJtavNEOZt+F1KaDEkTuzGz+vU1v3q72NvEoMSY
rbSRb3WwDfGtI5HdfaV2Ux/dPx1QhJR4MCCdMB7PLoMBGvZjTzc/1kAksCE83v7m
eVu6jr98zJTASEdMDAZhQOC1rY42DfKo0FBrEy75iQapYcszryuO4szVmFx3c/Zm
e2k9uxdUJRzltro4KPnJrXjjI55fRZ4eLw79CeBD+ZKwRdJ2asfoxA7Riaof6hX5
C5WWd/FG6mqli0kUzOrQcWpM11OU0IdXlAgmZs2Di0SIkMGjoK5w8QykBGYj0V3+
kcQRTAubxe28yp4ZfzEeIXsOY+XhvH6/XlINdqoVak1hIDtDJl2nmNYXdZJa3hrZ
eSmaXRo41iaKmfKBpcBFWW8wP9OOPrHGrOh8VQiQTzH1isB9pTHfmgXNVezq1945
Ub50XzSz8aVymrpURVQegnS+4RIkdrwpX3G6T4ojp2/uD22g+463aXq8d4JbKMzN
Y3IZMLCDzH6D0UiHWqlGiL5jwfUU+5iX+Y/K2uu1d0HQg2nINcsTex+ECYiOj/bQ
gv7oI4k0Ni8jf3yuofTRvTg+fUE2/P/CHdQmR5qDYziH5KReW2GvUbcX7UWVWsoF
JVo3e/Hr+/6qkIhvRA1bZEi9hRek/MGwWx8Ph8RTkNqNy/UunNDhOt5JR71JUzNF
QNLQAsu7qObxOYWNrjuPD5gwJpG7KcYYKabU2aZxKQi8BR7rxuvjy3UY7kPD9XG+
OrO0uNwPQAfeYCKPIj/UO1aJN/gCffx50Agu9EP9sucNAZ7ciLPt17ETVY74qgI6
EjbL55TPCXnICkUh5b17qnaHWzp7i7z9dt/fQF1sb65BhmE6/6KeqCbKTy2dfm/6
2UKJO5bn9pXnRenUBHeDD1rMlQBVpK6eDnYyJPCRg6ATDLEXTZAubEcZBWnCMewL
55HU14c/wB3A6WZ8H/SUdntlFGVlW5ZplbZ2oVnPVUQS+mRGEpiLu08QjqeZlBBD
+K0aV2CiYTMHASjvFI6dY0jy4uDVBcZA5Xye/z/3xJJTKec9HE3MFBOB4Fq/LDSM
iME5ak4Ct55EbftPdVzedQNjK9ZPzOzxl1j3EVifuuk4VCUcmIvZ9EMvTdV7ogHc
DyYl4a7FGL5uea4y+IIyC/QQW3vSQ3IxQk7YhrXHBRd9Od/brKSqxsteYEWGeix7
ys7MNLrRQK2CgT5TVHCnpCFachyzFps7xKEFeylaTt/aIwbUaxXnEm2fLMflBzm6
Xz7rBo2xgC++V80hr/qtUd4PKeLp+ifmS3r9Xna9VZGOQEgDnRSZxf7XYj5DL8YU
T/U5cQELiwaXmDnSoCbr0hf/rBii7x8qgDQzokFcJMqdIlZkN2ypZ84rhNWnvfbH
x+j6i49VMx/jy9vcYPRyIXuPPI+eupIonvncQx76eJU5C9wR5j6E3UrzTkcJ68sA
6GaigNzXyLetRwSBnhukgD5Gqk+1oiNBAIJ29MNdAbOX6mV0NhC017j8EkGr6IRE
a1Ptb2tdvLAfH/dRyrhdaof3NwZzIUUcv41Y9K+SJTcNAoAEhpQeaabQBVlqH2wc
6Et3J8ZYtqZn+cM6fljPttSH12x16spZhNwwuOupEb5ms6fR1CcN4TA2eVsa4o9o
TB2jsg2WKCliJYLfa5QDvhCybqTqZJgIfYl9eg6mF1qCK5dxNaKjCffaQOL+eSO6
Ob+54XDta0LtaqSliRKYio1spijNt8B41PMGJOmpIcWIjJpbbqwlV5Cs8H7BWW9h
aNvI0dNPY2ntN6lGYY8gqWHFvInntNsL9dXCIJBwLVS99wsB3dZhT6kPBjarUtoW
qyZVTtBMjCE8o9pBNVhkavh0cFOOUh16jDZKR44Ss/EA3GTWfbNF+uFov9TAOkbC
NiSqUKcBToDntIxGLREfLzqP+mkivVtBN6ENnVc94CkOM4s/UdcOHTKovk6AZiqQ
kBWp6El713SYl0uT32Ig+WBz5sK94UyQhu/pIlZfdLQ+2jAqG2DJIUIN3uLt1R0E
C0XEz6+TEaNfCALAASYgE48m22QkETw5UpaQrqThU3lU7+eQor/w40HiEAzHHdTe
+1gFxs8SfPasbcpYQcVI1CZabTtr/3hFnq0A6lAkaulbwPJiJOBjsUnKU9A91y4U
r4wDL/pCpaCvPOjLkhADVrPwg8XqdkLgELXeRr3FVB83GwS6Jr5S/ctL/+2vVzvq
6+ZFaIzA9wSZG2/O5qxa2YdSvjs1bwNuF8SLLKirYbUVadHo6msIbWEQ97LSzXQo
MynJkr0tgZ7NNDhbYMIXo8kbv7CYF2ov2EXPGkglRDFmHizg7GEzVlqC+FM/+Pey
Cs124NOSrfLaBG8HbBL2qgUvzpay7z5iarslFwZ/kzsCgVs/hQjTvqzHzzGkTM4V
2hZy4eo9t9Zyk5WHpYY47thRqA5vOrGxh3pPXS7zfKl+IiWAqgSFk2Wge633O1KI
WXcyMGb/RL+qHmqqILFh1Z0+v47fcxwQef4uPj0xZm5Qrliz1hr3fB0QbOmtKETN
5/kbf5r7Aueub/vAcNGeAOnwAIBckmU/D0Ce1LhALxaF7rvuTJYijJAKPa/haMt3
V6Hn+sCyRht+HxoRJyr3gKfH+5Ifmqj3DFbILJodM9HnqQybwEttpSwY9lk/kdyx
V8faTwZI0NM5maKCI4GOWoWI6edoON7bYRf7yRrJDwxB9iEL9+SzMT08WINgFYHI
2fY7oe4bKE8yKwrPTkIuTWWvqaH9emwKqbjdYFyE1mlHJ5lBDt8EDa6sXnlLU4HY
UKVmHjC6cIUhtZ5zVBDS/5gPlv6PASMYfPVQy09u/7kXCOYAXnX2f4hXrVrd/1wy
PiYUzCqO19d5DcKX2rsP4FKb1CvjmX+dmUBDblPw01K9SBTelSbvH59BwYzEEJ7Y
A8ZyYRfl5sWFImeNr6YQHtBJH8oUbY9KHT1zkgPaBGtcsb7YEUFaBe4zu/pGDunn
GyfaJVdnJSzfMU1HzNBNP0w2A2gS06CCXhCCori5hLZQHjSVBwVQmj/GCMEgZzYo
9bN7IDMK9ujhpRWlP5YIez9AP5TGuerAUGNnz/4tNUhr0PEhtU25vArO2+yL7gWy
238ElMi+pd3S+sLck1i7RZ1t8q2uAIjONpWvgTpO7qgtmBTPpLeeHAIYehNVEj/Y
4LbpYKfX6i9eUo2jLir/PhWfemcO3LjPF6A9An1s44gIxUk8ErJyQ8t0yDVD3l62
n+ycJX5g8ZpUS90KgULxs0OmaClCuI5v6UNuQZIODZCUj0L+/kyyzKrpeXBZ+Ylb
f1VetAWWa0v18VCsV22lZJiOen5zE3WvP3sJ7uaSg0CjMpYE2CEeh2hpW9tuve5/
MKlU7FeaaEBQ//GcDIpJwQITFdBE9DN30u2sxD0wyK0o8C9yAMhtO9LtCxcFn2Gh
7zefV++Xwd6ezwSEy4z+KwGNFaIg9ynPCpbzcJ/VkeWov5CE26cYBaxT38KscJ2s
VfR6tTx0N4cHke5VQ197yBDkmKZFjpXqxTnfETyrM3gQAndM1ALkccoE3/JsbVza
mpViZvWcXRkItq21CdxfH6UBlWJtBbtF1fVPyN01SXdvBLInFuidpO9CBYG3Fx6K
rmYBGFnjxluyCMhA794TTGQj/gMvfIDGMwe5I2QyoPco71HIFPg36NIbVYsbF2lc
nDPuDU224SXcq+tFHGS2pcy9hoIIFfwncqvEC0+ldUTDZqsYtvLEKsinq25eN4kG
r8IBpmqBqr5BKgemfzWUx3K4arlqJzxyVmVC+m5SiJJ/fTVVkBq8OCHh/y+BgqTQ
0CWCHWtzzkQDEHfZruPigRbFzjj5aaiexEqryye/wSmNzTT1pp6KXNRtA78WkAI4
jZb/5Z3MQp/bVz2mKOFoOaMO2gpIDQJjfCD+Yw5G760cWB+W4MEH0AKr+bIHT13q
bVD278lQqPNNja5O3QccBVsEqYKU8PK2G2aCXvekAeGYJWd19zJhI4K5sH6ENl8f
fI5hJhuEEXQzOguT68rI/2pZtorpFFtnTIKY1I+3wfy+9JXGEcEdIrJuWJ/cBHj4
oB7pUk0rMCTNfMB692Nmt9LREVgJF0FTGrnLja7Cd1I0bOJqfV0dGiqgoymSrWHg
Gq9wh4r8WRK76mD/27hX7idQrClKSLhE5h2rVi+Us+cMGN4vQW77Tv7eaITvKauq
ihSDGtmKxMRWnDbgxaKww4uMhdz4bTx6uQyco1NyDq6eIyaWjxt6LDshgkGXKujV
rrjwL8RAaYM2kOH+5n+k1l5BaTdy05MTds/bk8t0xfeeuaBHwp+dgQueLdnIXzrB
oSi2H3YhXdXKNcgmSBGC/iHEmWM5/A3tcqimmev2oQsE0G2ufo2IUlrT9/OpAczt
67cv76JgwQgkVva0kVOfGjQbE2RgreOBoYvrSZyS3VUA1GPUIRc2IbPd9BC47+i6
xQ0AEk/n4EW8x5/dmrI9sZeNG878FYeJFwVqC3cOloeKdT5UgIo56XAmcCzUE5RV
XYkpDDP7L3mGef7ftDEEzv+BBjKEOkRWBvY9tiLiOo/DGU3LTJKaYJAoFXRCJh4W
Fdc/SiS5zVvbSHIsGzS86Vu1ltTHmCc5XV+jG4hRMhY8Gnn/Sz1vwqiTic1YzJ3n
acGAlujrrp8SPS/jmjGTgTXMQ3Zn4UdyWAH/zt7TlooYZURsDrOCxDY+FwE6o1Zt
oj0zq104087fgjrtPxzec3EWVCgLqfYY9WBkyoh7gNHxT78cqoxyU+4fGeL0NdUx
Ckf/AzICwHbbgvRGLTTDJBRRaMg7LXcGgHU2H/ZqfEbv8L5y42ZySaF/oZJfeHGJ
68yjEAVu2LsUZhj4miWuMi6aDHQwoAa+uAuPQF5o2IyZ6ekKy7KijXug5ZRYescL
JUGVLjXB3KoPLmOHODpXRgG7xxn7QAV3QI1m58tyXdBTHC1YcFl4g0bAWYuxAGzU
1D0jB/H+19O7HeYgrMs9lcS++z8IAEMumk5ltVq6dILZiBCgLjEBHHF/v7R4keFy
q23bZEFFjsEG88ud3nqT6TScZLCytVIwGkTQlFy3TNU5+BGg76pQunCZg9UiEYA5
z9JDl7ENa1Q1BN/sYN/6YJFS/pVSIJT44UNMaxprCLsocMbI/KbjmOIuJgAd0GmN
dN231hJvoS6/z0Hv5wLf7bExFtZKyzebbCK2+J7m3lxo8TwufGh2ii5XZ5jjAuFG
2eM8IaUd+X4+luxZAgu4IRH9gUvicrLLsUViW+UaLcgwpCbKVrzO3B2nZnsw/mPs
8nkbh8vBUfjDSlleVayHYuP9jdzDT5t8Tl6i2t9i8oOo8ltJQC0Xyg+x9erepkkf
7DAw/BxX6jvK2jUBpIW665s2IpGNAvYwiyngL5aFrn+Xabb4LKTvi4L2hIdZ8ea0
/Fj1y7vDFrB7t1XWTxaEMxAI8V+hQ2vH+kpZRhuEw7N0XvZh05R/mIfnotZZK5fg
HdhgBlB9Udagfncw3WhNYm0OtNhBIjnVn6OPUILSfh7sAG9mzWVrPtVufgj39v+a
lwEaKNn6V3Jjlpd/25oSs9G5q+s7UFX+lI2n/4ci11USMFYsuieKOOvp8Pl0iX9v
9e8ynklja8G8+4O3/PFvhXlcoEQ0Vd+cq1tZCgRaMoFGSsaZMP4KDR4uMnV9x0jX
5t1A7DIQGkANswiEnLKjSmc1UxO3pZBbAKhqBKbIMDk9SJQaWl3UIbkSoU4Ledmu
Y7g77ZCdW1RugrO02N2+fHJNfoOitcM9scAA1wdOBvGpx7wTZa2qUSuUjeEzK1NL
PRIDQUqBU7nWGsBzzFv5el4xmi2ROBCnooHcNPKayh9Xy9iSkYo+T3JVc0UT/Vgp
j5hCg3a9Asl/6C+5HWg1nxS2aY3hGNLw7rhzR7pgMb+6bC7TOoKCjgmR7lIXEdGI
tpcReXReR3ryolnAa3khjEy+hFYZEDIv+zdQQegEx0vXdJMOFwESHrqS9oJuE45d
pZ5Xrux97H1G98az8PlHDAp36Hr87XIZcgVl82taL/Bk1XRAT7nnEB4NARcpA6w4
22iE6+j3igMKRbbA6liSBlFRj6fee7TCOAfMnfxgAGy503+kxBfL2rZeTzWjBvhL
7tPK5eTwzkev02h4uzfkLYJtR5rcGqJpUkB/VHo5YY1LHXe+7yvSeW243WfdU+oQ
l9itmTZHUG/Ld9bkKj+nd5GqmIKNXwVMhnvHRLaOP8GwE+pdflu5yG77uYeFODhE
GAtBnCnr+smFGJG7CazqPTKEIr2Q9f2rWDCQeWd1pnN4b8VgOJOeckKGVLfOv+IH
zKBPc0OwwCWdVL1pJ3Lew9yd7v3W2k0hVi5PeEDyH6Jg+TwV0s1sVqImTeaImQqX
ZR15F6/RQWzfLpnvlBSzaOTYi8/xIwckHZp50GUWcwpdJTVo5JsaFY/qZ8BfwIGv
JB+UTVYzfWJqmEd3OTBY5fSyb7KlH3hSlw8lh29F1gGOJn4mWISoRz0SS35FEaps
UjQrqtCiYbX5r+y0i2lWmqsGsTARUWE7AwFmxHmFoLWHC4lroIWCezKJlDnRbWp7
0ck212GZDXOaANLRBDK6IUQBPRJlE4DN4v7AdD7xESf4TNUzwo9igDQ4ceu7kZY6
SRfrxuDlNxD7iR2JNMXwsDLrfpvmnUkNAVIEvvI/I8rX44CKMr3MUmy9IracKOLS
pXzRuVshNF2aWdOeweaTCAQYoYkb7fWTZZhn818JdNP2ZpQoUqbBMt1g+vXjNjVr
OuGvBpg/qZ6+B8CjbDTd26e9t7zdD6Mvna/2jLkGxStTivltq4Pw0AnEr431tELp
e2pXRuecrOwG7N+WwRwQ65aIyEWyp6KkpqTgEfJ6OaQeS4bZbzo2oqFQA2H6rZMY
p6mjCvQ2liiXZuNNnYR5wKE365rENd05uW/ZSsZC3NjxUKi5qT6Ulgdcp3/Bu+Iw
JINXPBuK9Hj1Q7NJ8uFeyR5Egni+PWocqJetkbpkRVspwc7hKW5hw9mgxLwxTbvo
zDTqBn0IHEEYQb7y09ZKEJkUHk33ArO5rAb2GQesKKOceh/HQI/FGFCRMY+B3isz
jutr1ATZPoT1uzo3f4h26C0mDIc8AXE6lS2GhqXcaI8AeKCYwjl5kLhHagu54o5K
f5D23UFDHst5ffHNNRPVyup6x3GjAvY5RgufLPguWMOPnBlSmG2afwKKkQbK0jve
epMka+NECS/6jIsoNtW72hpvI60Dfcyqtmw7XuGW+t24l1tikcffw1gUIpzM9aMO
uAGUOBWqhJLtj3Z7NQobB5xDkuMU6uA3if9GwX/ooXd48UgefkTgccew7DAj20DF
/fnPCwZEGZAMswJRl3c3djw3FqGcGYA/UkqLIQHn+g/g97Ozr5TLzeqyrHsVJlfp
TdIT9kIXlxVfO2dMODspbp8iYgn3RE4UQ3VIUjve/pHqcqY+hmACzgXIWqHEdsg+
HcQq1pLBcpPd3vlXsC4/AZcqgLwy8pmAu4foSV/W8/F8b6Byax7mHVcGTDZHS2Y0
iInqh84gMAjDHIFBOYig8Nk8RgxItz9o8uiuaPgWO3UZ0G4h1tNL+viwu7jfcD16
0RwXHbauHEnpWecf0KMaXdtCqN8UDXt7G6OhfIvwQufQs1B0MLyorQzLXzsqBP9G
9RGhYwNlxfG52AOaTZ+mdjd07rObgUN1ktc4B4rRzfMQNeDKsb35N/AsbFpMbEUi
KQzISmIhmjhw5u8RT7/97NACwNnbcAZGElxi3CfLaS/whqobd6VutmEMtqS4i1Qv
R0yj0VgNtSQKco7wo7VpX2DUprVBiuZnrnk6zB69pIEG3P/l7HhOKHQvEOtbpEF2
nd45WE+XpwgaLcScem3kDmSFeZzEe5poWMh/PpHR4EVraxaQMKTmaULCEQfVMsTb
2CmeXGzxAJ9CkXKCRcWlChlU0s8FPWkYU8BIa+JHVW8m4jEMmDJK1RYErBdmIPxN
nr+qMPOydBDSeEN8GmZ7uKtf0U44H9QoLTMLt9T9qm4RBTJaK/swGVta3Quc21ET
ulJzG7T4Sm7JV8f2cVcfFEobwf6z9QSdBcv4wYR+Vjn9CdL5kc4xFkcnVpwtxv4S
w0KofM84KEGVGMT3c3jmS1JbRLGGOKsbZCxgBTOVfXBbE+X42Qik1VIiMdTKTxmt
nFSxnCiSN3GaclVQWykS3L+jUwMpDcaOcVEig9+A1jMrGsuui7eGSsqQoIFMEIZp
cS9YYFITeOfIHT6B6Ip9eviM86oXnZrJWBR1oABDPsN3WofsdpabY6pEUl88Mvj6
7alzIaLC65ZpV2P+l/Xd8vXToMsK1neBdSnuafw9mGp+0Jl8j2iZ2RsIBSRRJuaQ
3G+HDAhzjTIwWPsqK2Bk+CeUTGp3U3tNFB/rP/kF8IR0jPG+zaDIL+tBBO0ul/EU
+tD4OFDdwGEIsFSeAj0uM6dbhhGMnmMGUGisAw4qLfEAqq29SyQcfvx72dlvxZiy
lL19zjwchunk2EJPhcXRdxYVrJo4xFS2jysmxWIvdotzVkelAvof6XDpvDj3Y4Ar
pse0r6CaLStuw5PXxbGZwMCm/pxiNmgFq2e994qcAf0STA63FIwungZEFC16aoxr
EJW8akQhFrE3A4ofHOFyQ9EWm4bnqGQVKlyLa4hxH1ehtUsGFhBHNf/Hp4xPZT8d
vGWXU1zAR6ETDjO/k4F4GgppWJoJqF4tb0YD/gGTgHBiyzn3IdTvg2LTn1xKdmIl
wd2+CoUwVCLu5PhW1g8YVXegt15HFWgkDR99+ucR2NGDFHdxHAlOk3/4SX0Jr3FQ
O2Ajki0MIxSsROjJ3P1ONmWqOC0G4x0P8HxXoGvWvmE1gKhJoFDyxAzO85FOvgQp
2nz+UJvRs5EzCGB8/1VdolFynuKELMtbvcaKC1GVSAaDt4tBTYbOkacOUG8KzXaZ
V45eOidfZEzzVb1oaBsBcgyxPkVHN2ZsTQROCFQ5mFwMuxnEEbuqgYVkPHyuPs89
SWQn0KYBkDUjiRdJBERLXLJeS8PcQeV1EZkKh6XS4aQ9OZX8xZJSFrDqvDbq0J/b
wqBV+dFwO1Qroi9pwqTjNsSbvn6n68IZdW5vexujVE0mI7Cx2wtV5ZezoZqHVDgL
D0A+cG0HS8y8VaQsMEuXMgLky+X/F3UYpBnATUPhwTflbNLKxSZqsqI+RGFtT/B5
ZTYVgHghXI5fg+L2Bkq+57J6oNYvVc62GJfuIRnyWsqeV/n9bBNmTq1dGbLKZoxr
4eVB64CROki/rcmbHfVxRkqWx0fDhVq0oOjn9Q78A1HQKlNv5LfBIDo67Kt6ymYW
kBNXvvo/Q/XXg9+zMDgDMKVbOb46sVV/4euNHZ3vPhc4cjOi0hjPaNeeRwAM3N6b
MCt6BFmmNQYsWKgketiTuDMcBui1dNlSrEvxjkFjl5XtxzkUEV+auW6TI70wB1S0
hiew6R29xjcDMctyZEP/kMlY9oevm4mgcHxB0UwJQ1EhjGHFD6SNiD4RcNzG7Hh9
+NAz1IcHvn4aV17IMRr1liP2DyubrISu77zPEsb3IcFPllq+PTDfzvzdiweFw5/R
vFH3Qwf9RUD3e/e3L66pWle4HFwt6BFJrKTh18OeZX7ftaoEfV/4B7NAPeEywnLo
IBeTss/yJrACfuqFq66KoZmtgD1zdGnQbI2YEu+PznQlQRPXGftFlI5vrRCc8Mk7
0rZcqR4u1YygrX+cGdPBZolq/nHzdUSXpCs+5TZekwXU4cvuPbhgGe3yzPW/JRn1
O/X1B1NZqL5dEkjrKM8ARUvEsA6kirHxvHJMtGJzjeoPuzcLQKN997ejPI4SuVan
3wxNQeVE4PixeGfgay02RJl5ckJifd/N4+/TltcpIHbkzq4ZORAE4+5b0N224o7O
jamCIRVn/NsSVt9udW4KwFThxcTp9NjpU6nnTGiFtMoMMxtlpJPhLx49wN/DdnOi
Mav5WuJ99WYdGEBimPnhUfuD+O2JmDCBCkS1kC/wgkgKYicZU9u5U+idgPtlXzK4
y0FAdQdjEKMDoWQDlJkpYKLt942DwXhgulPGwOgzSwPwQrvYRQHPqK3E+0B8j36A
BE9fzpNKsVB4n1Wmrtgkdlua79vU+ZnHrEWyOYx6iO2oPD6Ez97TZsdzIEfhobH6
WadItt3OtL6gkyqQNhwZUtrFHb5zsl7reB1exjBx3n0fsJkONk7Xbg7TFYZVsG3w
F5vws66Q0PWe61bRI2L9xGukMmoL+thwP9/M5ZwIzUZYfJEjFnZ6Wrm4Rk5xJqMa
A67MvVyO2gMTDLK8r9CYBDThtsIxG07Bra6ti4yP2KSysSENaeBGjWjjyaMj8+ct
zPuQLR6D9yg25F9GTj4K8xt08KwAcSDhmR9tD0X4GH7qtfxP7HGpbb35gtI8icxQ
wxBx57GEv2RLEJD1vETh300QsIaWaQF+6fwYrvw2urSzICj0d+4WzB6OsgRMjfy4
1dUFqdWibpCeDxIYA325X8bD9LRXrWfZIPSaen03JUj+Wq0FYVqxab+HAfqb4/W9
pXdQoEnTQt2g8+5LIJUy0sScxqqxbIEzlH3+petT3qVQdiNeO35t70rS0Ig2y4M3
oSKaZtIdduTKCLqJVhIvGB7Xb4tBX5l7lTxrgegk66l3nwzDctP9BgHx2tVcI4sM
OrnqqCGi4PPj8PMnHvaixSsAWlgT3DcdZ/8VY3atSTo7+odFYaNlRlaI3PLr62pd
fR1ffs+D6Ty/qVpwMXnc17LdwjgqoX7OqHdSqc7hbMnV5/1FNh4TrERqmzgTdTP4
4Y9zcBqBc+I+wRlx5xCWe+Tw1elan/hJiSlrYwPnX0ffKsLHhLmQpZGcIaR133WG
Sf7Z0yud9LVGq+TDB+LQJOgVJ7ZEI+U/mevrRfAzwyJ+7kn5mi7szKKfV8IZYD6l
iAqLRSRyviaez76TiW0qXuinV/msT31SKUDw74s01DUtYQgPUxPIzRmxQd7aCNYf
xMiFJ92NZ6C6J2oUfp7PzkjPYcFl4FGwyqQr7aG9BSBYxLhuS4nfeAxm0nkob/ls
xDIR6EZMiKonl7ecsiKD1uQThbEY159Z+AwQHPzuwuDFCMIQ/fITLMauxA/AZ7rW
9fALv8IaDz/o/DJvVmQ771gQLwrXkikuSC+BYBFWaq1p9k2SzvVmCyui4fIozblr
jgkUxZzfbve0njspFxd5xiJb3GGCPOICybDPyvCt+j6icNxFF5gjQeOCPCNZMLZH
O1ILo8TaXfwyevN3RimtEqwBrtJi57QUBSOuJ9LR4f68UL/xfE36rPIkMRt3pTEA
ptb0ftgaX64/haw2dlMPNsyYKgvZmFvCx6FRmKDJskIZh3e90eJF2Cty9AN2IsGo
HRdsgF9c7ANe8ZIUmro3CCkG2BxJZ7NyaJhp98xM/r12HVGHXgCfjBTpNdWV+KnG
3I9GdBxAcefau2fXPvnDZHOyB3yqGkdweD7VTqIHKv1kNqZAByMmU2vdo9df5tfQ
G/WvjS43fssR+M6DS3ggblRxJ7YxRImThyG7jNj2ichIABxXUmjGUQL0Fxs3Pl8U
90GKklOEEF/pcwZZH9SyA9jtugcdhPV+2HulwnylTO15Kp1Ms9vSrIvivBVnG2We
yNKywpzmqU1AxIBm8OWwePbrEyDO9nRbyJugZdPXn5x3VCsiOyer6M1yFanXaVJL
uxr1Kj3X+5aZjbEWUg7+Nzb0kUM+y7j4t+LhIp21qZBDYhDY32eVNbiKzk00dTRi
sEuG5VlXOhOjqxT3WsiLfHxSxpJ4KKOI6vAC2LxbdP22BudiLfZ5HzRbbJI+cvF1
ToWxhZ/LYVPPap3NJFg9kG7humOkm2N6oea/M/K0EoNrkPNIS9Ff6HxAen++hEH5
z+N9GozuUX2PqQ2gxvxjK7keJse9NpOQ0XKUfYnA/FB/lJEb6hzp+W10J8lz9Shg
rs8Gr3KfiiBlUfyTQ8nvkOWIni/lEGWltrQs8KUh287FD431c7t8vNj85PaEMLTu
mx18dPNAQh51sSx5gFKmBrEDrCh7uw1Hjl3LFJdBlVRbIiM086AvhMgEeG9nrfn1
kP2ZcQVvysm/Oul+GvqW23jY9o0Tu13gqYHXKiD4tud6KR0LMWmkMsXfZxuqndLf
6I92aIRs/FjIBjRCUYyyh236kKKyREYs5wihinXJNBfZwVQgnmrdnthmTEpvFmXa
DF7h8olQkvwwnDGbefreDrTW+fOS+q5EROEwuL7d5+t6Ly6IyRLKOhVc/ZhS9efn
xTN+p+CzHeb8UXTFs7DMxDEmMIU+mH9JPPFxCVFoqU8sZjhw4j11PN8bUh35vtPc
OJDwPHD6yiY5YOLde7ww42QDNAh54LjqNG41NSXKnAIdTKL0caNreJAwOvDktXdA
N7Tx84omjIurYWVLLAWMVH6lYFROXlJy0fdRxVHqj4Cwb3GpRZcnEkVMlW4rK6ET
cYnRFp3D395lCQCQx22k03fyy27jCARI0k/7KQ7HSQa9mDHYyhgDhZ0O1FzGcRYj
4LK/d8pD7QZ9O98gNA94txUgh/9M79uHyhjdTizJo5kJQR/ZuZ2JNgMUqUXOXEq/
VuOiQl6TROeo2TTB6G7dmG/C5wGMF8ktdwvAIUP/RRribKmNYIQPUwjxTFwlAlmM
2xTI5Ga5hgKNeUPh9MH42d0lUolXXc4MUnhOv8QPkQM+zqxE6NvgH3oIpmnzMLjF
IgZdNY/g/1vzN+bmxzw7xg3QcDpDVpVGG6n+EwFrR90KXCqLn1XSWl+5LgmhmyVq
VyZNAdbEcpMKgQzSeReXiQ3GQnyjH7PYbZti+YsDZS05Ydi8GB05cE6ddVpPM7r+
tJa6tsiCVyL0vhQxl7H5qBwYWdWPzbtRrtZ4076CCut/hzZE6pLBgZVW2g5NT8y9
OEwqkGvpUY3/Bt3ZBLPt2dHfq00j7g4Oaa9n6Wo75JBJrbHOgr7xQi/+G5TAt3Cn
tFHM8GxFwBQY/JPfQXwkSMzaN3EnJ1eU7re7rq1gjen4riE8ExkgvOZWbqav2epN
XO5g6KQPeqIgp4nimszdutaYPAEio1fisx5d8Y8vvP74//Ue3FR6SgZ4mSwbDUG1
dOaXZuUIqMYqhial/Yl+QchgcD6906/wUCIb46PFSvzsRHpHq3uSbdaqBG4jKzLH
ylTjRAmERQGzH9fftdcguHI5FSEA66KXdBjaKrf0zD3qsXEYVnJzDqcFLgHR4oIO
1YwbHhY0yAP3W95pMFkjTnpF8vaSrQA/YqckOv61Ubdki6bkjq8LxVnb1X34l2ax
EBS7D5QpV1nbOZ97GZnMOVnugNvJP0R1CCCPAsJYL9pas4Pb8MohC7UhzzYlDV0J
+GTHPjTKmtz1z2XNhFOxQy2sSSI1/Bn/Je80gdOiUjEpXjDZllsEnP84ypEmPwJu
c+1cQKpqXLcwJ86cAd+aFGTGgjueZrVmZ1V8qyD3ynUQoB3+D6sRhumRfHcZ+Llx
6RzeisHPQrV4bArhaVHRIxsPFYU3u+bdmLCBq6gnAeYWNdyVkY3yMaN58rPj8OyU
63XJg4EmWpG4UZ5IZ6ZfYGjCigXRPIdmTtDNF3EwLrEQOMuog5TyEe+W0+SR+cBY
WHjlZpKSRYtSjjuvtZS6F2lVCOUDGOpUDATEQyj3pj17pxz0MM1symV82cDRXtN4
JggEM9R/xmbTfcq0zqJUIrbp0rtVpt3jTUfm8Vewes5D9D+u0rmP3vwQTs92AiIp
Wrhx239WlIK/bzFqeXLoKfwESua0N1JV0mhzVN7/8qllqVYxMyRQQStuo/x08iSu
9Cvyx+ASX65z2uRC1vorNQBHvTzjZJN+dZsGKA2L9cojcwga2ZzAqhS1JGi1l+ol
Iyx/lCuXDG09XPOJmORjYqHJn9Jh4u70WLFNem8anKlg0L0T18xduKmnPXHP6kDD
SVtM+lcMZE8N9cKeZ8QZ44n0a/IEgmZUhoRsapBvoWLoSWIN5D/3P/XQ+kihJWit
Z3TssHFcZDtWc1ggIbVMp7mAMeFlOGcSqV8kfxm/o/nP8KFAYwctXxopowj7kPEA
0U+Y/7KihRaCIncQawdqH17iiPMcUiLvQ9MbTo/0Y6IJy6omXepLFawTHDehd7ga
hrfQhZUZGoZQni40aO+LPBusOEcnYs6zLFs4u6kpT7+2NoaoKErMioG5MJtvjx2T
lNjEPRvyIRyZsxffegNdryf2XceGkzWuEad3HAe8j5k97JAhqX/XtorTZlHfP7wO
TcLjMGCl6uuHmz12DFUGAWKyNekSTt7NCaFTz+tRCC5fMZ78svG4yft2KZWxrFdK
nPvfcJqPsGwrzguoyVibvnLwGlSkX7IgrMAW3oW1wleq633udop+eHfR7iv4KLpQ
U8QjUWeCtmk5GYfv89LffSoDRUf3ApAaxggNEGPI9yEPD+q2EQVq4JTr+ofTWJy8
+uqAj5uTc8NhLgFUIK+UbzM0UUA+gA3HSQHPSqfukehfR7h6meSoIIreNqr2trwG
SpN93tCyg+2VdPK2qA1ZGnrVcHgRU7E4cSV1v6bu7FTCrUOdX/2Szj/5VWQb8aeH
tC32ewwl5dNdFWiMitTute2PuEaiaZ/H/CxT/C6RJLM8SfV/ClGO8PNx2Sfp/G2z
kO0xaz9s4eLheiJCWNsz8mz870lDl9MpLIbzmmjJF4W8QjEtLSk+HyPFU5EoL2Vd
yfv5OdrZd2N7h0xBQ+LoC1c3ZwuhuLpvzQgKZN2/FhLrxmmb+tlcQ4rr/BqVbCUd
7MPtKzBmgwtOFuxcjUe4RsaZWilkZtlJfLpZES2CkyrvP0mBe+YbG7EwLhO+mKY7
7NEUnJ8NRzUbRrN5G49iZLn9Mv0Z0KmRs2Jloe9h2KC4alooo7iAjxw9gvRKY3ut
dPIQox8P/Sz3DKw695F55jg9x4INAiig3yGbv3ZpgwNYuEXRCf2TvJKjWLLiPS/3
bYLZMoRhKnyvlpja6N/g7IWwipK1F6JRMCXM1t8d+2/8QFBHfuCmfsmQCRM2bJLK
v/bm05BBYbMlB5N5oZOac1cjrWxfyvLsopTXxaPOPUBWnVUpMRjMcU0/2WwgihYC
uCqvpZE3VijQk83n7NvN7QW9aYF9lnbdy9qCgdX7/LlpMtVYHDmeVDFONTRsuhK8
E7tBaBj+kPyFd2NtfZzJsPb6S06pG5w6uMmh7qWokjz46kQeEHuLCEKt7z+qE1hS
PoEV1RppeCd8q6bLK+BNNPYYNaL0dikviDbf3jOGQU2BzBA2BoGKcM2pipjUtBg8
6vrF9MIvjIsDSd1d0XLGmtWLA6BB3zcuOW+zYDkv62LCT8AvQnBhZvh5Xkn/ODzM
6W5RzijwfvHO92SmLCVGFb/FckMDFzdVAARQt1dqQCEwpT1hacY6/nNectYX0bG+
WUenCj1w83fncxeds8r8ZX8A8ZgsLE/vE4XglCuyZKhDQjHUMSL19UQxxVclyy8S
1sg5KRtUWTegv48h506KZpP+kqxDYBzZydPasVJVprz8j8EtUGNWRmH1k5xmSS2a
vI2bmOGVa0fyn17w1W/X/MdiGrGX2/TCYpc5apZ01t3Etb8rlTZepvcTpGzVD7DN
kWfSDDWWe8X3VKEXfCEN8tmrAVJ8/C2nIpLfFcwkFHMsI4p1z8H7Dwn1G+196Z3U
oGHN2TNbceEMS3z15ECzmYbWoXP5xllIN8F3y+gsE8PVTaLar1SDaEn82aqmFD3w
YPvj1ZmWoTToZ1kc2gBqd0/Wa42gGhFTzHD6AU+Oocs6Z5dQrpUuQyuYpp7VFyvI
CdPSlDghWwSX9RsuBDO2OsxnparAErjwpF1c5bkskstJB5jzuJbR1T7nEU49TQMT
vReuZej/oO5eJogqoN/RpsE/wITkdnuy4Mvx3MATUsG10/Vi6LzpJ/f3WbsZCa6Z
KL4IeHKxa5GZPU+EQNbOPEaM6kF8tBZV0q1d0/mwy1uMSGrlk78YWYbwiHbvZWg+
VANgiXVYlCfwslu/5u3DJLSZgkLSh5JARGI9e+3snopcSMqD6oUL1VnLUDBxA7KU
89QBfCdKvdRCczQFK5fxhU0QB9MVv8Ll74kYEVVJFb0AyHo0gDhZWICXuyPohGBB
8jhpFk2mXnaL3P+bYz4CCYxE3ICLnd2P/y3Z5b+WW+T1oW8y9HUxwuVFyIoO8Qbo
hwnrpaisS9Bcv7a9MuihSxWayA39w4JFUsSHpb5F/egPiGMpZccD8a8xkoFAi7/4
2/bvJM7j0PzeyqU14g0K8oMwOiXhMmTLx86rIFKZu3APaT2BGN9L8hoESQwEago0
ZpaJhLHJTL+iU0ycQvtihijZNa84AaX9z/sF5k8dRpljNAYgBb1QRmtHUVEjyT4A
8c27hM3lbBvZ0IPki1OIVUqC+NRhwumoUsjb0vxKOdb+ATMu4lhrFQYAVzmEO9ME
kSGSpcLkV44Xwm0CAykayuECLK/Nnz8toekweSVgDjFdyO/OhoCuZjB8kQG+vrov
S6sMi5QAv1ndcv7f/p2L7Dst0dtZQi40++442BnCPngr1+xAG/cNpLrnGBEso5H8
T2mVz8hseqI9Dsr48QGw3SPHB10AZ5T0sw2Q0yxIctVKzwhoa9lVyW5rYKdX2wwZ
UhWxqBdzfY2zEktuI+CR839K9NT6FIi+47XqvrsrtwWr2zbdjx1n7XVd6PZtqXvQ
QGNI2Fp4UXCzejCGrYxp9tVtQ5c7CSSgimTSo7et84IG1UlyPG40Aq22GzNA4mIw
Dc3lXejG/B7Htd0x53Vg9HqTSB6sWl8Uiy8YF8pDhR/KCMwScMtn7yi8YeRJwItN
CIQaM9CfkCZV7WtdurWIH+kUe5sCXyZZAM6wtEQIX5xOqKNtI3/JrWnPd6kLL0D7
hi8tQpYHbAbanrZbg4/d0zgHclJag4Ag6VGe30+ofs0gbt2yGk8FrvzcCLaDc1z9
O7glPdsfQnUFbUPgQM18U1fGeARcrCJf8CprNWJ47H13dRS1UJSErzXSrcH1RrH/
Ly2RZtginUHGPhHBeO+1impp0GQyiDbJDnhj7M/GTy4Z9M2VyBI+6JcKGIni6dF5
61iibvJQDCJH7GkS2M7ydDU99AJVOyr0BmnGIm6F3NDoPQWg9lAvTwe4aFBOYD9p
Bcr5/ykkhF1IgeP1QzpcAP995X7Kle0XXcrmDg2FVGmCmQ2hnZmzsDpjpzGWg18p
llKtSe9Vi3/OZ5IypkNizi69Z0QEURGirhzNOhqvDLjfvFiAJeHGtqpHlzsoFOxf
T3+KOZZ18StYAlnCrKfZ9Kd4cmandUlJh9mNDhfTzkeCZpdFtbC8nyZosQ9kkoSa
bZDrYqlEa/GybTg5dNuJ0t0xusOJcKOnOrVV4MtDvMK9NXCYmsn5j+NwRvmcVZsr
lAzLl7vO82nbQKorDsEUgCRJXjMCzOccJyF4wSKAjLrJPvOXz9M5z0I4ksDY7kSi
dMFEV6pxU2KHQbTxr7vBPx4SBpmHNXD+AdWPi/WilvBLLrBxUZosEtB+Z9Nf2cib
Cpwc2zcDBosP0hUHQ7zojgJzUQ4E0i/qpq5l+OO+9nQXxjcOG7SOOIUqFSl2Syc8
Rut6qJLX71YR+4JPjv5qqpqrxMM1yUDWt8rJQ5N4kyNl5KryW7g5b4F7X2IUKXF2
29joeVt2hqJiOpVYzpjtL5t6osz2slN8LgQ/uonTDPpET2ARzlE+pdUsvqLBY8Wt
bsHoLOFeXBN1bTRYDUXbzAxLXcdp1uK2lrEouiqtIVFMoMFDsv1vftY6POJBDD/b
hAoJrOQthQnFHSdCu6rqXQOtfznp07ZELlgqv9Aih9O1accISPZ786uhsh8xv8fw
rSyuc/Rm6NEvK5yMO+R+AZsSjvStHMueB89QURlSC2pX5X4cyQhE2P1uVQDsw1s6
W0d5LUtUME4RwzZ4/ybf8IcP2Sd4qpEL1J6d7QCdOiEtKzLxkFa6O9kcuw+mpxm9
j2vfp0MwtSmmAx14MWpSqEPQ/TgaYaZtsG278ZgfBipJ1MxEBwBfwtT843hXVGeK
HEVhTWQW9xFrw3oR9cU17zEk6yARKO28Wucpgdb0wNu0lGODDRhkl3zRQlNSsyU9
BLnF4Rk85fYu+5h4MOm3TAHaW4iVYbWE1Nf90FhoMOeFFHoBYGqyqab5kOLSVa3L
//OTVAcu/hW10p7z+nnVoXoBJ4/5SMBSPH2Hov2vfusygDJ/0QRIdwhGxXtMXFiK
nHxhn1mNVb9NfhtW01+vzYqrA+3vBzf1xWb1ZYjMXO3vYmH1K5zaCJdqdeavzBd9
rtcazbv0rPdebxZnFEv4x3Yp3ebjzQ9D0EQI1dN1tQz/5C/CrzxRMgQM7KbwKDSI
ytK055XJGtXYnWwEdZ+t41gcjeHq43emsFZa9YFkVgnNYB3JowzPL+bX7Yjc3366
i1fF/IfA18AUvPK34B2Q2qW+BkfYHPDNRc8jxYi+FQ7mhU8/Mj7dW2DSXDtZmXo/
d8sbFjvIofea6frE49+8ea2wIFx4Axm3POn0sK5su01pzMkkna809ypieK0Ct+vj
Umpz8Y6g63x5zYmURrvv5VaoJM1P3/mPGX6h8mEF6qK8weoyYw3OK0Mj6w461SOL
HE3HpkJlHE8/UMfm3Dp+KmUgescf5onkiS06o867CmysFTtXamwoa2S6E0BLW88B
BXLGp5zFB5Sm8uHeiN186oSEz9eCVEuuUF1R8GzwtlQOi1zAWjBSlpFjgKo6FiRw
TlVCo9ZOs2O0BNytDOSaKdVDuVipSmJZUdoIHjAOdSAQRxe8TAc2d7ziIIyuRs3f
hqu9PLirC2YZCV00ktW0ag5yY/70xKQdTSUt0yCH9lH46aDWeZ8SeovX9E73ckwA
Ii5S7pybivPIA6bCN8eYtEPONnAaXVFu/oS/hMMhJbXakO7DuHd5ZqI0Z5kE+fJj
/fyCZA2tiRHTk7XdKP7AwCn0lfRjUXhIrwIueU25G2EA59W9/df+7Tz1xc4Y+KIX
P2g+IlydBPSs6GcqXGft9jGz0JtZnqYyU1US0vGUYX+RiwEeCebVuNeS++ORnK8F
coR+3iGEA6537dQ0CveCCHHoB903x/uANPRIy64J19jYP/JtPHxmbjJvEEqPTF3T
lTOaT8ekvDW7OzVaUs3ocaoh6iPqGC0wgj5uSHLUaQvdo3MWb3Gn135+li1YdLWs
OHD5bFF2wmWlQ6s0MVgaPkzaG0sroLqQP9tJiy5U6Es7S8XT+gj2ULdLyP6nsF/q
aweNLaqz+PAn0zWD3JMzxCng6dtftz89Y7AowNcPOZlOFZUdA0uxuNg+W+bgmvAK
VVEu1dXXx4ftEqVUStsAHGszgX4lma6O/RAPhIa+iFpkxY4j92PmM0+LVDx4eYqA
K15zAkdlL1FirSSDaknI+UVNKnuKqU+oGpvn+IIcaWCSEv26S18hp/w2X7CsU13a
Vc/TztCP0FshWKGqWN8ni2YKCPDRzsXoOZ1hpxyJExkvcxDKzhz6d+OlAnNQKAer
2Yw59AkCXCcVq++CloCshwFHsiLYweVx2oBhwcWDNun4pYErY+6IWXBeaNskcj/S
c3ddoY78X6qHeFQKL3cLw8AyDoNQPIolCssnvTIbmZ/3xssqaVK9LqlGdGo/Stpr
erZxIh3Tzv+zAIZ0M2qkkQk1k3paGYMgV1fQKgN63483o2Gk8e53hYofZkvo9PVI
0RWmE3kajjHx+rcfj0N8xFlxYAJT8aeB5unnLPhMp0lYYzpCr8L0RkeDQ9efzXoL
7yehphCQ6uk8Ypx8+9OfGpFUDIsHGK+s9GBH3iI0yFUNYJFsVpz1kVun4G8ZSUDd
12ou/bXtna8dNHRuhh9NW9ErZSY8FDWOlbV+0zZG94LBRj/qPY0n7T0w0/7OWnhB
RYiYLWS2KIYmp0JXyJj1JRRfQNwZNDF9JndKNUo50Yqzr+ethCPuJDobHGocisRa
zibWCsTilIZPFH1EgA+FLKgyvPBJydVrRWwZcPyImU6FunUyEldM+xNvYley/U7v
biLNv9zSQJBiYmCR/jD4W7/EtmU0zsWe7Q82DaSXqxJu93p426msQ7oIHXXUAT+F
OoPJpcUn2bXWxs4jNZTugNcn2vzqDMDLoucAUeRD7NMICydU7vwxkdjVjomGCmEW
xWeTLI2+eowIIEvtgwiR/1vgkbYjVJt6iSR0ATAEZZutz9OSi/5+V5iODf9yexH9
z+/9lFxtFat27+K1G1sGNEog5uZrIHG9ffeTdie2iYfSHB8yFozozZ1uph1GXnoL
zdw3M3FyxF817sY02YFXVtZJ4/lxTqxIiUT8QUPy/xGVCJzCvOeaKjRR68QFe9S9
bPw/npYFVeyaGXzNKSp5YUM2haxcbNL0s/EDnWgV1RJEVt0JT9xk/m7A4NEaIQFK
Sr++sA/byf7rwlq9qMhAwSpMs2Ny4C8mRUN2kxp6sNGrEfT03WQKkVHOL03H0o6s
vNnZxPOcWckVGKCSRcQDzOWKXN5M3Ft9WMDoFOIgwqucyNcp/V/XbDRlyZSCIYSr
0UJ49iKoiWgfAk85zdo6ZMcBkavo8uU8ww8vRXoUVbJRGkacT3eZk1nIzfnsOGEk
ICg/pORcHGv67L0yunEZ/aBZcfaikIu/6V/8o7JxRaMkg4Batqh83dywZwn47Atm
Czdv8bv+aTkb1bWpQUzu2IGTfJoy9V4gG7jy79fhwi84ZHDXgNh0WN+pPErzHvrs
69VqWQsvPjj+GPjydDe+H22ls5CJCwpo3ViS7503W1t9JNtg5/U0JdBg76Pz39aA
XYivN8Gca30cGu58L6G/AcTJW21IjG0EEOh4i23YXATgoVCK0+QjMZjBX5u4L/T7
xzA+SAchscmVDdxZVA1gTAQ8mkqLgh73gWiYtaUKaZ8aNBUzs7Q9YvJdk2/l5i2A
539J4QSDiRE3cgbCEeI9ubHxPb58GkqBqoMQZ3ZGaFn+ehW055//zUY/cvMhsTJn
xmMA2htBMKxpvQD8sNHPjUChLJAvi+mjYQenmANOik0TkvpDTcayDTwHVCWSBe0V
7MZwdTDMTUgY/QeJ+pHluM5/t7cxlQEpwMloT4/JYqKO1zxwdhysxzV3gQl9mTt7
B6D1SYunM40YwWEA+j0dxH+3FDHbb0QlcY2YVNhlm+U58uUa2S73ipEwoOj5jblj
XNNdEjDOSNFSOzGqMPKDqE28ICdPhUgYsFARtu0kNNBkq2N7/kiFHtJQPjxSgIxO
pVd9xH/H4iKXaX+JpV+LsWiTzMA/EljHh02na144BjoQcAqdqmXgRXy+Tz5NUZaY
PillBRJFnnSRp4IiRTbPgT/Ot2rRDTfCp+vO6vl110j2lkXVrukyoi0dwlS3dncB
pBpPQ+ges4vjT8Egb9tD3vUwXY7u478O+GFKPrjNwLg3ajGoCi/ldshoNZO7iBYr
SX8Z5Txgq2FQjIrT4zHs7FLLmpYpsWOyVhi2+G9wXkunoB6kPUOGXMSyAIprIJJF
D+q/RS4ahIn4LYTTR5En1VtNYpz+CL6ZVDeJix63ejB6+8LYqXKa3P32cfrHOF87
5NHGfPNKIYSvAOrYbbs0zr/kNSMxuhZttUuDuMxZ7FMAxN06Es73P1JZC1iqFTdY
vxtNA3HHS8tiURUq4LCKv7y2yV3/UeCA/IXukYFCQ7wPV59flXHpTot1/unt3CEq
V/OFc/vvCpM8EHW3O4EM2RnHhNkoYbWxvJIYBvVydn9mfSwInMW6zuF1+A3U6tUw
5tqc/s96GHalG5rxzXFdfPqjbMztm8cRVB8WPMJVPCBMeGVz1MQSkyQP+g/eT2Wr
V86VEBMqAWoIfLeiaEnhFoEOc29gsVlxyxBxCPn2HeGbJNWblzcfAjzLqKlnSEc0
4fHnpdmCfm8u4yJuysgNNGdhDcytZ61gz1E24LsHevuCMb9cT1/P10auIzK8miuL
g39PBpV6TrFJfp8515GiTSP49LSr6kztPEQ/cPZM1Dw2HdhvPqvEeeg78HA8D5r7
uKyfnpuzAQh+nIAR5jaTmHyZrh1bZX2OfqlYfL/pZm2bOJROZBVyUDR64lZuKDl1
f6YdZS5ZwX/o40RbVDd6vj3mSCV0S2c5eReZzK6rErZK301O1iXswEUPYbJcGugu
BfnRg6B696sbvClkggTiUc7Nse1qnk9USkdJNNnAYo7lalnnbZmRjwIyGHiBx9mv
Mp0eTl3CUBgCBOD5KZHvFRfnK0eg+SknejRd9grKS3gt0Xjykv60dVrBSt1Hc/mk
pAHT+Fsc+opQ8+1IzY44Gh3Xc+BC1hmP8HDA0vYdIV0ilUlZsvfCIjEYibpNlQJX
UXGoGYJvp3I1gRedu/FFlvuSKlIOf1ddgMEMl6PaaRpy1oqH5nyTSFY4c93zT0hK
+kuiCCMiO0lmi/PNNT9+Ro4OB4wzS391jyoxDYO9M3xk0NImoScCpYSi+7254bv/
8sBu3zsTxGMVJD1o11Dqo2RC2sniAkzkrrxBKCGTKwLDca/1UuXLLSwbIr6V60Ep
6joB+si1I7U/LkXeKKvmGV96p3oWR/zzqHZYz7JFJSZfSY3A9ffhbv8fdKnBhZDI
vNA6IKXie8oFXroCQgXHXYFGXA4Cp4cG8R3LHsIbVVTrQrbJiSWH6WoJODeeN5MR
if7d3AWdNhCaCES3bSfRehFE4DXTbjDcW0N1HsDASKecvT0EMiL4SinHjvDYgA2H
fjUvBjYYzVph4E68a/NR/Qqw3UMuYl+R37dOPr9ctptrVEUrUpY8ioVsy3a/w7n3
ZiJE2tUTt9Mw2T5Nui9/rS4urdcrQ3XXgaVh9h4ltCJwLsLDjPcg6mheZnOW1lRN
KqO6VPBNaIfu3u9RkCGBqDdOQYH8XkZpJYD+9B4+2y2NaaZmmRPRD+DuzWstcjoz
wCHQkHGYYBBY+Tx3V+Ge4V4nh9uU60v5NbRTIbKAzMs5e3P8zw1eiikyWDANZgId
qO85VS/Aa06LKmsAeJT1K55HIvGX1QTewPUlHuDiNPPECB+j2oIAe2fBgftwFAyA
p73sJT83DggBAVnGmManuQK3K6NWwYrwfi6aeUQOjaU6YOaKTEpKGkYgwd2bKpqh
/Pwz3GzjRe89VmD6zNTGCTEWOPGndFOD8s5Wrq+hSb8hagEbhdKgp/Q160F20kcl
0wn2rprqbmqyq0Osf42eCneRooi5QlKACqoAdnLozEgjTu7/EiKcPxeVgiYBOpnl
xwdB/n5zJbh/sZxcl7ahnlI60nRWGWLj/JJyrpfeVlrypT/ya5CNH4FXSF3x+RlB
tj6rSrhKCqNvh8MlAJiJGT8p03nG/WEdHSWwwmg44nYSzeAVNtE1YUzU7Io68jAQ
MOVIGjRAT78kqPPZ8pnRVsHMZyxsgPJv2Ekdf9tXzErH6sARMbqnuIMna3qZWVPi
062R56lzUaGklDbqbDQSkcN+lDSvt7zu2ZsOkmXwzKHtP8upwEPOM3FWm+rIBUt1
b7CrZVJkfQBJIrL3mAH6cKHXtPhcAu0RoSV8FoclPvAJTeadYoXmXJYZwitMEtGp
8BshGK7gKsKi3EVevfMkZnFg3xqlE1pLOoCvtkSvGe7rY+WjBdzv7j35ZbCCo6cP
4Vb+bKYVfXe6Z4Jlla4Ctox9UjOEXx9BSuCU4M6WinrEf9V7wepojpyOz/kz7vZu
Pq4yS55nVHUk5Tx7zriJ8x3FZipDT21cHG098f1iauBNmrgiOuJwuigWad3Yye2w
4JQT2BNNWu4sBZoGwl1K36DrqQ6WA4jk4s9U2DnKXMOry4hhF2OL+3gSlWDWiHKU
6RX69lPqXvqNo9tw+JltT4T33eQo086nBLpIjfOGFk1+vu2lLUiE9p8aRBgGT/nK
i7LvfPHFb+VcKmd+0VhcdHeAso0gFGgnF3zUpKsyQvbodVG8ozAVt90w7RTIWoB7
a5El2MBzQt7Q4dC1QNYaf41p7hhK0Wd2XpULLYDPHKCBHSJowB6X7Ji1tJeuxlWS
k8K+ylhIPjfVJSgjeTDjeT6082ZNXyoXlCWbqDkfR25k8jDslH/wqd3Dx+fP0ZMu
hQWHTnUefVFXJJnpzhADcLXtJ7XnogezjZMd3qJd5YZqiqNbWcZcWWtT6a/KFw52
dMfBBFdBa2tKRS5LjEpc6Ikz+MeA9v35wVD/k+UYpmAlIMlkdP2sAKRM1aGpoacb
SoSJbTG9wWdut5zmSURZ5ILOVBYCflItU5VLeYPUKKH0SvCqxnKaNqngQ+itOkaT
b5lrcCHmXIAiT7E+nXqong3PaVHH6DlrtFuL/cto8lKLq5ClEkRzLR3oVnG7JYCx
gYPsdNLiVtKBcVVTALHvhYRbJGwC0VEYx4LD5PCS0VLOUojNfG4XJiZqKQExzCnh
XUPZrgx0gGxy/fkz+5YWN8Mr9KrMcpXBkeMfhK/1CFennM+us1rUPTPzW0EzXlOB
zfX6rkESC1Xojjmi05KU42w/w1agxE9da4n+k15YqmoRcW5J8joEuqiKVBpedRzr
eZJEdu9jGL7HF3HdX5latqS09+vI+HLQcWftQ32c8mjZEwrNmPLF4vKyCMa7gDvT
+V+bYbb8OIEEWNq5mMHEqvy1kcID3IpsI/U7bDyIhyTKxzl4LtMakHKRlaJSNNb/
L9nYqAYRHdyduF6pEguQZd4aWsmRB+nwkhtlAumbsbjmOl8B07g+wSo8Q1p+dFes
LVr+bSn8r+TuBoz07Auacj7rQ33WKw2xl7wELIvJqz9zRTtMCDEo2+XEDF2xX+bD
XtdEIOpFx4QEGGQMZIFThr6QkdR2gWOff2RL0uFvWr44Wv1N0a/zutZBqs4ZQj5H
l5awiEuxnhU/5vNKPobQc+0YKe/TPS9lkcHl7LksrYByFzigeoi2+thW4aXQaean
OZIBqU1FpPL10HtkT2jXLIx8MroF6n1DzNQqxUFMU6XXDYdzNrAXcAhR6BnKOHVd
6Kt1widQ3lgGs8JQXvG3eYXw4VFicqQkJ8l8imlM6T/MJvOQOJQn1KOefnCQVBZo
82m5fqFe7JMPY+2A/8Mbt7JeTWPifKqFYoEp1gmadDDmXEGRXkboD+exO53ipAcY
6DvO8CZco9hPkACRVBJMBY+XFG8JOIG9QtqLTne91YF5PKiS+J69rik1Ey3somv9
y4MDvRaCXRY50tB9UmDsxQWfahAClh9ubxEx3ycuzB3jEsRcDvjM1V9/4NkW2vta
TVxgNWWNJY5wOay60I/4qa+imlrF+ObqmzT+VVGZ8NSjeISycXGhpipnH+YJTThM
vWUtJeDjCJTe8KH4wG6zfaex3wMtOFVrrN5ziapkKX92ym2TWVDa1OFU59HhrJoC
d/YMfJgYXwbokpvIQzhj19lk/UNCQlQQbznujHIJsD8vgvjIneXMnlzf4skV/mGD
7Im93YOQct+KnZOBKazg23cm9WNSfJ1gNfAT0pJf5cV61xZLhZd2Ed5jc18n8Lpt
ZSGs9Y2t2aXg0KzD+BtYM+a898EZPO4lKA3cFQrfVURVEa4xFRZj9NGNauKrtcEn
vQcSPddngjWutySpLGJs04ipNMg4GBeVIB0R4cRPqWkpA/0APnudu5QKoKkA7V5M
yfeKoI9YzCtA9ibCeoJKDnGFJHJ9FwrXDMpMozwir+NREZyROMrjWiQqZBEVPet2
2ZWmjTcfTTMwqjkacv2V1fBQV1BQkEleswrMIregmjkE4qtYZ63JSRTjz61glPHq
b+JV8plM2JqbAR5WZAFupX6tvmdw3twCyHbBuRVINND3CqYhgBmuBXvqtpI6I8gI
mh84CMyyt1PfQcSJMgKm0gj5MGYzqJp6rAlFN6UFxcyuAqKZo/8P9kPD3HvCWVJe
Y7Y26vS6mgYzcf5fhOP1jdFlMft6TWCTvoKzK6lKoVSI9fcE7HX9n1H10RsZ6alM
OAbT6HYELnL/WxdFULVrkMbibVXvM+q/Dhy//7mZg5XniS0HtQTT199XfWe1asOU
5Pc9/1SzIjDlP1uiFcmz5N99iWZpK49Bv/qUP3G26n4butQKoddLiwa0gmL8/ygQ
SigRV+77YyOmTWdN5qSrN89WrQyOpFjO/6yk0NvMXzGSHYW7VdO86FXZBGmTstcT
oH3+qldDKnyOsIoAhF6/8vAI6sFxqPjpHfJddfZR+2VviqrGEsMyLV+0oNAowXba
1WqWdranbHN5huAnw4290ktW6RG7nwbLvOkF6m6F4ZIG32rlCBQghcNTnDqChI2T
3bqs97DHMKl1ShKhK2T1gn+ATTNW/DqTSRD1/slq5aYXA80Ixo1dFKQ1aP7mPe7Y
QEzgzu4rTJ5zfbd0RdgNQ6OOprIO7/vV5csG7bfZKz/ljoJKrGpyVGOnFyMNMOL4
ZRTgUghIEZNpT3kY5uVRGhqek+EkIySdXcPAIFRv3UH3dSFZixfzWJSQMmKrbIY7
T6izuMadg1jfnC8RpEySQlGDJZ0Sek0DzaRNN1jInzsLLZlMwxJqWlWNg2o1RVp8
w3wWcF0/cLPOJO3OhVaLHZ9a/SpYubPRrN+8IQkbuKMUSLYeTSG1jTnvIMtmLMC2
w6egogm80Or13yN+jUw9pJ7tyegTZI0PWPhavuJPxGmUxWkMSxRyGSN/uCr7pKqu
R2kMDNA9GpGty7hjdThiHnjDRqcerbaRqHadY5M72vDbmNn27cWjoGAQFmf5sOxo
BLXyuoujQZqDIvmXHo8TYJCxI+b+w75h0NTqcTrHQRkgrs2E6YW+p5iuwkp/kNbS
kN6d9SGvQKI2Lm/r+k3VALlDlTaTA2xBsRv3kl/w5+CiUfELous+H6rdTMkHBJVv
KsSiCSoYdYCqTj8TbcqTFIUXPbpxyVKKcydCog1vq1bMRtH3lalEaNNtEd3AXxDV
ujbpikNxqQkV41AE20nTjQEr1w9B+miHDQuhNRba7otfZSIIWm3aJw7HgNhMr7b4
owoEBGyHMSJx2p7w1OoyQ0tpP44syHkCtNB+9BYPM7pWHl0PUw7wmoHzxXuB5uKd
XnvTGFqUG5BONR38Aj/LTz70FB12Y7U7mL5s8g9Js/1swAc/qZb5bL2T15NW9dhh
eCEoUDVNdRG9d/FwQdZYqKj336C2b+cB0lzmpfccTKB8JzzI+HScSTRNmn41bdLZ
fjBk0jGNepSuL9bWEmv9/rx2Pp6ub/s4KTa9k3Voa0y6Ppsq+B375mJV0Az7ID3w
MkN9gQaxbU2j1Nsp/otG/yq/JKNSOq2/iuslPCIRqIKTynSjkr2Q0eYP4BPd3Dbh
+6T/gto5LZbdH8XF2YuaTdC+KlIEL8ivaWiPZG+tK2Alhv8XLbfqNe/QPIf76Cfp
3+oT2DbqyvPJK375RFZ/tSqI9mP3heMSQqbOByX0/3Oj0OqyLP9rxnhgOS2HmRgc
0ZYRSYuG1aBq+K9yvnoJTGuFL++z1P/l/RinbT+TcP0Ns1ZeiJUTAD1yGt3nSV5M
ygG52+TIRyq61r3YefuC52Bnx8IxlmSvCkl9QRfxv/8d8TGU7vdVzWbx/7pKSH8F
Mh3AJfCZk/HkLJjUpiu00ru1kiNkoik3VnsYPvrVKRXTC77Lo1Hcw3OSb8VSW1WD
xwhXNa7oYNplLKNwQwxXE9ObD3FqIXYRa9LsCl5OrJS2lVNIgaw6PQsSGOAFvCj8
ytHbliKLtW+Jx6bibIaxe/NyPqYWoE1Bo/VP0DRUTBNHDrRkGLvImKS+QWXwUMi8
5ZUV5fGgN97TuomoAGJkooP57JOGKsZu5KH7Hu1V8Gr5gSyN6gPOpBVsqsQNsFCu
OaXQbmX1OdbXGOIXNXUlGrZcnMo+aEGIyV6c12EeuaDwypd7JQre0epbfuMCqgP5
MNrSuVRUz4YbURp6QjLvJEsChV5GtmZrspacMn1Yp9s1sfr1lFBEBVt0KtqOx/HU
zY4A54xBhCTbxjLNFp2ZQbJdWWQwkMXLQsO1KuQ94GfM/JYGxS4AX3cPtmI6ixrC
h/JjQky8Gb5pNxGQlRg1y540aPJ5f3wpwk8UmR9sx4/gDy9wOuBeRiD/tt9jAO4Z
/XPGPR/DnKP3crBVo0pZvPg51aR+wEidT5TEwyRp7zLpG5Y6dwyh9RHsRbnTmUqc
KBIjhZ+XLzYIrqgp4Q15jK8Fht1ZAwjVbAXpFFwYmV5R1HUy/cH2ihBXky4FqqzZ
zXfhj/oj36m+oBUsm60dvOy1HVIRuVDH40xDLSCj7ddArFVXExyeT/CCUneiVFBR
WN8BJu3D5zxFEGCB20TfIMk2A2W6t47uLBhLY4C8Biuou5NFY2LXz1sbSJhHk5bc
5NvphNS1wcv9lQ614DsRToXErrhy8mJvXkZ+s9Fn5WM17GF+zR3+mln0gO943jTV
EpY8ykWSJ2yhUsLATMYxg0k/CORHu85QL/cgJ8jZmCJVqB8uK2FdPWBUauhY+NZS
nXDaAGyfYpjh//DJR6gwymPcxUSQ+7Eq71A/LJamJKTFCzH3YbEd7klsnaRjQh2R
cTEFM+tEgznGnxJP9okXkmz/fpywHN7d211PfEgcc9hDD8R6Ud+jN2Zc83VelJVl
J9LSdCe4HBwtmDn1ELxNxMd4raHb95EdMbb3/it1AwWKE1JFpJV83fgN3z7BX8Qz
E6Nqzv1/iVlXznu6DyN7scJV4I1r1ySutfiNQr+0zNvXwJROLVL2+IXumJp6VIta
TS0Qcw4GSOUAjkSGgRaxWjA+E8nIs2g74I0pqFq9DfDx6avQdpxWgLa52F9o5dQ3
RTTClnY5hU43N+aPGZapeaB/Ez5MSORmeUA/aYO17iBLVd4Fr1fTDv1wj1XUgaWO
otJcz6Wf/bJ97KppEEGDNHt29Upu3NlzjEKGq/EOmaCunTI2p6OyDh028nLLHPFc
EstGCOYzWlo/n3Veue3YgSVnIR5XYHtYLUteotQK+WkwoP9JaKxZ7jug2Xe8/szq
s6qkoXq93XpY50gZzomG+5HVK4m8Q71WU3FEcKvma+Tkh6uSwPUzyEpFIkiJp4sq
cXqZ6+jdz2E+teRdImzdY8H5D+K9hzJCnVuPN55L6hWuJerReB3xJwcUDF/g4OiA
1cQrPvKpRsZcafK1ThHHECpueRA/ytD7VwKoPVDUAka2C5lKzRQg7URmbl/ZpdnL
U/aYTMSrcAoJEkM4lDbvUueIN6H1I95E9a3zcfGDBdYhbXS6jW4V/DDMafMhh0fA
kqaKZpAd7nbZm1rFZuktr2Ase3Zd9r948OuvUGCXgP/FTX3aB913VeHr5chqL4HU
vgPpyZjQ8TJbxipjZryI23qDpMJNX1Rbzbz1NSh9h0keJJY4BJtl/Ig1pVE+zPwb
fKNnAjpzUQVsKq4SVHA7bXQZBRou9Bgindpa8IRCH/xWIYVog2HfOOGs73J/oHr1
1g7WBVuZ+gBOssfyvXmBRvyclonkFUiuodLhb/nUwDfk9HRoclvBxQmCMfQZt9/Y
IW8NrBEGE6hKQ/B0wRLPkORSvj+SI4SZSb2r2dJV/Y4+x0GrvuWkCv9pHFfcUhps
5IAkatQrh0+DXCcKpyiDDCgVge/pIZkpL0T9Gw34Xnmpbv4QvAfWWgTwBgcT2hxe
sXFQ0kED1chGUICPLUukIKke378pKgov98o0vLT2I7JT+RJ3Eyshkr7aLrRqD8tu
RJKc9XxMWpJtv6z9uUP8E6MBprWv6zMtlwIVCNmiO7PXSbOxJFcxLWJ3ZVFukAlc
0kxJI8/tEGyXngMKrI/nNIQ/G2XzDJUgtLfAa8tMIaijx6wVwNkZTfGienzSg4RN
SXBB+uakqYJMWOYNU/oQusQRKurs5cYMc4PIsmDDdGCWF/+OC17UzNBCHDZoUX+F
bfayzBcJEGz5zJaBiHIZ/P4GJhzj2KraCIOMaksE6wxLBkRv+VRs3QEYSwWrdBu4
WWtdxU9Ag2L9dH0vvyjM8qXBW+EnYVXDa3Gq8mtAFCemv+BFUREhi3KIjz3uub2V
I6Qo/ksyIN0eNPouCfPwTza/eiZX4etIX33ekZcMvzDwu+QZb2GKmzy27aNdzgKM
5b+izP91klSlpU0+fyHFyH9nQIyNUr8ZsI/aLmHZRHp5jNIDfYaC4P9VStVw/Z+U
c1foV6fjhUf2ql1BspQTRURH3HFMHwOTcCpfq59ujryhbqeVu+r3Wnbg/z4ANu1L
JkcqSE2R0dQQ67lf6U8c5t4EhnGxyq55a3RzH0Pbjx5EXOPXa0JNlowUfr12zqj0
6X83Ts2jETqXnBpw75KYADXoAJern4I995kV3pQ8TsPiTfsE7SyUtPFF1URNv3sL
zAmuPKNg/0sM7c7O43OV1fJNGAA6qxlprwfwa//zAdsXVtBr+fzlaRG3DpNc4UGC
8bpEs4ZPO9DgSdyS7R68HndcPP+VJy+jeJu6AudVwafJkuYa1pekkDLB+o7XSwsb
prmZYTN1MsUmtceBodB1LSn+AF/pqQa+RtbwrxsUraYpn5OGX4bQQNX1W3UiKJaq
cyEDBGmOFzVgeIliYnqy8NpT45lB5OOCVpQD5q3vIUimkDynX6KiFFCvfNxy6Qez
dvPhH+yL7jMDAGYogfB8c3rHMM7YHcAwBcG/BJJVZVUjs2yeviHMBFDbNDHaL4+R
E52VWvP17+mEjhyO6q3IqoKF5mVG18udrRMaA8xbcUWjYuFffB5QomydA9D7b075
P58BagBFxBouOMQx45MhsKDzsVYM36p7pF6Uto38Y/FLSZiSDE6lk0JHNa6Z8e9E
Rza/hXwiyaD5NTvCpI3Nr6gtBSEzPw95sxhI3Mrj0iHF12hiAVfwcVQBg7OP1tNU
4LWdhXzZ7ghA8oRYSSipyYn3CoYa9Qu6CL/mOeUfz2Z3gW5Qu7WaFSxJiCj1RD7r
XVOL59GjLyij9Ekmu42uoQC6KRoZPbyy6MEJPsMZ7jJIkv+WmqPvfkpNGKNryVIE
yVtUPuQB+6FT0r23/kQwU5IbxZgHVDnJL/Vh9II/6UCsBVmrp/CR+VUxdc5Hb95W
Pq99qPjfu82kLXFO1vnRmync/N+YoHhyKaHtA9afeVRHNEM42ghxbhpAy9DPYC5W
LWAj9sx074TK1V75EWg5ixYYD22l/kJkZwra9BtRjzLJrPljndU6m6axKO9Yzhgj
wmZ7nzoSo/c2BDVwMaw1Mvj9jeWCvUJ0kHQyrUC3w1HmYe5v/hYxxn1Juh0J05M0
kENKNKSbvK9CeaWHzxKdbT2JoGZRNqnvvSRrNpJIhYezBrvAMv4U6DqUHpF7NECE
kX5x04y0X6JJgMl88y4X2ffw/DiTIqjWJCBqor2VwPeAo76kbsGE4Fs/tioB0oii
PCV78lcda9co3h49c4ojEBFd8IV1XEJfePqSeDMGo1xojoryXRO4iN6L1HODQT4v
zPb99DfyxJ22uVszNQiKwhXDaBuqmsysI/wxbx7n62kwuolwi/DgszDO/5TiBiHH
7M1jJeZY9ETEYqglm5g3rNb+VaN93T26DLLSkLowQ9BFNefqkh1JRN/3n5+Wrkqz
pVZlHbFidvZMYoG+qFLa7Fmrdq3lXpNvU+EgqJFDH67VwVozGXQv/w8MT69iCU6l
EWwxQXc7n7ff8kAPt3PIuEo+2Q7+q+w6R0kjWKeVOI/kiOJihXp0+0PCV9IZuwoU
f0WDK6wJiDGVo9WcD1RcBpbj8HnqzhyK4EddJL5fCpaA1Y6w5DYl45i6poKGMJkY
VPsnNdEhgaAhrPm9pc3MOFFueCZqQQDxbOOsqJjCtIvD229EdPN8UEwr0FfUjLG7
aWw1/3E55U3EP6UtDGVADDPtGnKxPbe08ze9ueS6dER3MZXg4g/T4udiI5q+h8/n
3AQjd6pLV3BHP0n6zdh+xbENzjMzS8k6ANLgOE/e1eUqojTglV8Op5ZC+IGIVtHk
CTOLuoBpxg7o74TPys3R25kZwDBF9qX3pTiAmD0pH8MpS9Cbbo5kkSANdlP2wtvm
zkfFH8SvK76CEC8sO/fav7ueY2pfu4ZnP88MqyFVbcbkhvVtKu3Rspt+lLYfHX8L
jlXrTQQbL8xbK+Un6qg7hzgiFYQ78HSamks4x9ZOqEI9DwU/+4sS+UtD5YJNy5x8
l/J423ZD5xR1NbmCCiDXcMZM0KgGycGGoZcd1ngRB6sysGLsGrdGBMetbY/RdtzJ
ZB0qWEqGsbut58nv8cxjyywDMkTVGhh49CgEefsMmt0K+idoWiOB/rgdsd+g2Ywe
2722v6/tzXZ2Cyoc7h5QqNXbh39XZyaZi2hCYsmPwUDP+0Ht/TgcRLOOWN0q2GBx
Iop8Jq5snZUFTRC2J9R4Pvs1M1K/mRsels93roRu7orOvDr+txXvM3g6FGwPIWEt
KY4/BNEmDlZ/VouckzYVxVt7ZpRm1+y7+SR0t1VcVFzL+CYmwP0b47I1iuGLU4eG
dZAV1/XsCQDKJOwG0KzZw/qD5miS+GM+tKb4rG+a8NbLuXCfMk5TsJ3XHrQWzM4k
8oY5Wuqw4q+SGmGkFAFWgdfDJTKzFrigmzuYEDWOgLEbdeEGGxndXcISILmz6KPP
8M64cZ0wpjmOER115zfvoqRlfkeCQ1txcrKDMM+HDzC+76pOce3cbCIiYtLWxJY8
EcGS/5biyruKWZcos4Ct6UnF9eFVsA1ZmQNzeuX2mZuNxV9k3rr7Dvcqt6k/rOeV
vA/UHmf+KE+UWx0LELtu2tLe5bOhbUCE08YCWGg7ZoOy3jYrbWXnfODiNCuGA6wR
OwcOJv3fDX78rfNU1qPCp1sWHZeBQesoeawR8x0Q5nkKNJF5A+i+2oGIXDH9xwKP
W/iubGcGCzC45ZySihkJnF52+0MIdkJ4flPlkMHh5UuvxMTLSS5/WyWR56D4+ms7
3xqnLDK2LO175NzF8o9mAdBa3Wc5UbV5ossbDsxZvH6MkMYA+XHHt5Vv0TCfwtD9
OAzvxVKtceM0nuqm+KJ9iLw9PF9q7yNl41g2Y7yhUIyCdkoofUZz2cZgX3iQvPL2
5RWy7RzJ2X+nYiR1Y+bzc8/596MtKEqcxlXC2LViDUExugw7xlaTw5pY6wU/MfFc
eAd265OzeIPMHRV68P3o9wC4UlF8hGudtv7XrL2e2mNumNtMIbvWGC4VYR4qn1c4
dJtGIw+u2hb5a9zk0j5wZcbn++gvCveYnT3x1ICuGe0TgxRANsAetnx+fCs4XZ6B
xL9hU0ltYpvOoLUJAqRQu2qp4TlSi5MrdUeLX+95Cc/RF47VrEujXie0W1bvcKxS
yR4ZqmaswL6X3wBlK7mVhPmnLRsErJuGfN03HvqownXuRytaFFLz4TvrywqEndB6
mVWFXMT9cYehWZ3e9koSQlSNkrr3rRn2T9K+gXFj1svDShogmORUVJrN7FIz8GFp
fTDi+Q+djFm4M/a+QK7j5SANWDkx1q6jfPlOpY0Y5yfet/Yr0lXJU/TDF4Q2z8dd
VyRcdEBeQJHrnrM7CBx74YSVmPSlnsdr7YvkxfDb3vcfZuhnFgX10JIAv3G+9W8R
zKjT9ILYJtk15kD6Bw6CaKilOTo48i3kHIEAqENPcx4FOOt0NTQJxV/SYCE+mk5x
ydxD9Eb8RPYrMQiT6xwQdPE9q9iU7w+SMbXgGJf6rbss+kKqCEEnZpUxoFlomjCa
R1w5iFys8Kq1SpL33CSV/s+o7tnxafHFPC53uxDaRK4q1kRNRz+G3zuToZufVQ9y
G8FVB35HCtPC/FYmIgIotZdnpyB5aybi6QXVAOWTh+xbBN+ufsq6m3obuhiLScAK
LbHssSXuN2XWaqI96cTAmBCvcorLJ4fAqo0KMkRK6opMB/jc3PQDyKYaDqGSTpqM
lp+Vo7KdOQImRMFmpQ2Uwo0kmk6sLWgHZRBpN9JktuEUpqSLaMhYGflQJTmCpPOG
peX46R9dA1Mm3r4GzUk3rSDOULSKnAt65XXFFIxmpFtdnbD93SwWqn3DQlJyTdzg
+iZEeqZ9yp3hlvkq6Pdx2SAbsataNxVay1xmspqTGpLhZ4iGIG7PpyWHtWEDI8m0
PaWDfId0dxNucqgqi8MRlH9X7D0m244S9KyOh0hSt/smL7dxnjPE6CinIIv2C9wo
6+o+mOdCX9nYSVEdemKV/0G2UGVP219iVJB/y93RV3JP7Qbh8JC3asUlo8CGuORb
bny0DD1kAW1KwJZzsyZXwuo53I8zhGm7lEENxPNY3VWPUVw2KFChsvH33Jr9Agoh
0rm7NaTHysdRPVg9TjWsDuc7vEVG9I17SOXEzSSrykI9lX5slIDpuHJUGrghxg4i
rlDfLOEFzbdswd5D2J+7Z21kn1kIcWL40JnP1Uf6xGNF3Tj2ELJ45WyornG/mqTZ
psAWcwr5x8cFj9bSiLIP5+cQuRNFelSl+PWPUOAWKggChsc/WEqTZeRl7Mq08Y1m
034dXtLU73fyzM8WU1J9EWtOJNvZniLDbe/kUew5djAohZXzCZed0792CM1rttPC
kFC/x8VYKJbLBOvRgcTm3o1KJy7KtELj6WH/FJ2jABda2ibsU6hVEuB23NZ6Mvt0
13vr7nibDs1Y9NMxUHjc9fJre2kMcoMemZwzlrvARMMcNHDE38p51HuhN+SvJH2t
SJFI+feaL3QHwoDFpSG4N8qXxYaVN6OzCyN8RFdg64OAG1ZasrJ0sJcXveGIaIJW
/dl1Q/ggcq8kLv4leMKEltOxB0vhcFKOq3defDibbcjS4QzitidRQO6EC4SwBpMT
tbeBznaU2nqeA1rJoJN0hKIPqBhf2LPPBqtMRuUPmsxd4usgeqN8uxi+3qWW9tev
RrhDLIp+o9SgUCwERdsu7fpp3Ju7P+iVHRrsGy8pypM4ToxYlNxjLKdQ0bBU8acp
hBq7hMWO/10BW7I3TzzdVNSzOggS5GkCZG0FsYiOpw9zLUf2IuK4y72XHZ4K8G0X
ScGP96JUBgKIUFPHsc8Cp13IEW3DqqdKAL3cbs2pqyRuSdITrRqNk4syfBkWZ6TJ
TPPQQ7XYeddvt0zFjFLLLlfBM3Ut8Q5is9sQTZBoVYLypp0bgKIWSzrFj3S7XeMs
DgOaP1zsVtDSdffiyJU/MqvY0U7oiHwk5zx0/yHoYnfXMPJGzZuOJvtznyb9iPI8
GoKXmBy6VwBWJqBZbxBCcuQ3DobVTwFl3cclRGlDn+rp/pTE1rFvbFzerEQjfzJN
85LZkpyjE5++qMj0IebFIZg8gjEDGTSp1AR29P+GhEUgvf8JjXo0WmMHkd9K1Gri
uDRxkGlTO267fewpR+HvSRqA13n4ymzuE8Ny0kKvGiPQBaWBgIAoo4FWHqBug3TC
MobfJ0nK0aPIdeYMG0s6cFkw7RZKqnd/ged282axPUauOvhA7BBOhxlMut+UjaYV
CEo2MOsvDlB/FESDHogFYL911NqMT+lJOvrd0e0R2ThDgF76QOtC+gtgs1Wp1u3Q
Q6VnfSrhPsEdnZbSRa/aBZbqLe0whPNZng68ahQ0dQO/WuB8iOaleKtl+H5tdtmL
S4zPtwOgap9xeI33OLNapeVat2a7dSgHy11EgZ7XZcH8zUHh26SyuUjrJjG0rchw
ZXIG+9XYy/bFZznGaleGU5DxdvCnro/6uhTSfCmERk/rb8m9VX1tE8nqB1WJgVL3
2HiTVV2B+Efs5zQx+zduWkR7SFmR7e2kevKaDeilXPjJXqdrIx2o2QUdmOdRybzQ
0WCVRaFBdKmUv6yp61XXjeZ289brH1nsVWpulMX8yjY/uDOI4FaNtaf/O3jUy/uB
qKbdv6gtXPTFp8jGwJhwRoJwOD7JJSmJ3RHBSPcaKU0x4Zt2ffx9ulubxvtAiEhU
90d0t4NdHwrMe6qIPnmh1ATNKZ4G5MocNcsDOyTT3LZjYbzEUfGaXygBXohvUYYs
g4PC+A8Lt/9IglMtTRHtDCw8O+Tint7jnCA54Q9mw1fpNl3ahIM30aceW26fBGWr
X5wsg3gYMLXy38jjCVP13ZTRZ/WNpT5ao3nYYZJ5TgIslQm79jzpw7xSh03a+zVn
VjiDw3MsyJbg7U5t9ShJSJWO3jJpfTQQNH2h7AWawOOwSVERJfa8u3rycBqtH8a1
AXZeIfc3Erkkkyo06Jez3DSV608i8Jl+AJangrsf6rV2ZZlI/7GJdFO7DnGhGf2W
Ho71s3qJblUHOA4Bwf9ly5BcwhGLS4lyxdmT+X6B5Zp3eKGyiw7locAiIjWv1Pb2
qXa5YPaRFQQnqO8G9NdSh+vZmJPAIs/JRnxTTRJT5XAb6AFvmu3zfpqneub8MACT
5FDwrQBXH04P/Sk5SZ1TE82dv+Eewt7Tr6yH2zjdNIRlpDDw2xePjT6mSRgFsJSc
jxPC3pm/YfpljjGRvKYopJiAx5TGIH+jvuV2pFOWLzSdyLJcMwTdNsnSVUU1uw4R
CibLO3jqBXCiiSvCl/6qDurDBC1q8/K9Fweagx+A1zD+l67Xj0Kr8X4r7ifc89e6
egVLVPZo0xpnkqNzIhrMGSyCu3+cwEdhmxDb7j9fArFVRTUbNcU/i92ySc0aFCKd
RFJXLGaClwoSa8lpW1WS7+0Schyo86pAgVry2MlOIbltgwBD7umG9o3MKoWTGfKR
675Jn2K7dkBzE8DOBkDN+iehCK3DY3E/1588h/2SO+c0fuUKYn+SGJqS3NWAtWHR
RsqgwVINXxhN85QXVOE3fkxaM+z5qdZtDJr7dIEeVHEHNKwILY7xC2NfwdebJJ/b
6d2yrhlcBPsg2qbD7y0h6aCd/CtQhw2RvgfkU8mcyAhvARXeXKFeefi/9/x8/sZ3
NQtzZD04ehVpJBOWAMKkv5DKinkjIAHCQEenkHDhJTeUZ+vbEB2xqeOj5YxQthP1
idin2hD0bx5WyF9C6p2ruK638Ty0OumyL4+8ueKqUXXkYjcEsoXNH5z4K3QKXR6C
th3KplMAksO4xeejWS+oQhdwCToE9i6djEJgKfENsl3H6S98eMf2xVoXtPZ9v3zs
2WG2hWEwpGEsEoL2gFRj8s9q5vaJjErWxB9XmCi2Zu6F52gp+1Cmue55153/y33v
DB+/RaDzSU+Ew9rk2Z2JeEdqcSBYbaEhBCIu18sH7oJ3NCeS6Vef9wwtvbLzjQp6
ZrnJQQlXkl9abAC8j76LzHqqQ481Ey6CJHhz5Fau+uNFx3+J1cf8kgtZlNlzObZq
uJpLZTi6kx/vmcYqTxBVP8+9ZDyrrd/ImSwNTF5/m80g2ZCycFVQiYcqCMepTHjD
Fl9A6zo9T7KYwOY9QOmGBzxRyqZgLLWOkZ5SEhmcQVUwRR56TyETrVFox07g8Pk+
n/NkuV+zK6M61jkcgStI/Uk8mrizx8TM13MQeaclGa/kaUnQpFUOszj7LRBHZOXg
ueWH7Gm685DXgkUaGSt5rDgIZbhE2kwI3Vz9vDg1kvwU+FOV3yoq7jF8SCBb4GXW
Lr6laTOKp0eBcHnXV2yDv0V5YQCGjRomFz2ZaO3rvw3A1o8xLn78OQONokAzxVe6
6bQbAbn+zv/aolx98IWOAeKRavKF9KOUw/7peQzcsjJvCBns27L56t8SrBd5skto
RyRYJg2GNA99wU8Ie6qONPy90kvCZLoxd9TmtD+/MORRJWvC6Qan2efocZQrxCCX
jumeN3QSeULXIpcWSvLUBaMUY4tcGot+3QLVkTFeSyvF1O6udpldLcsEv7Z4/xfG
hATMU5lWxCAG69AeQNRYavYuPuG0VklbfIrfjcrQLptrYCMuVlHUGCEKMsqGVeAN
BI7mJOBM8yaJutrCUlNVeZjpKKoxJJdxJXlsC6tNnB699j6XBmKCmLGqRVO217TR
xFtv/EX4BIJRVMIiHtPyQQ6RQXly1DM2lji72LviYupTj6dQTLNeoXV4sKRmRQBB
8jAQbxAwgWHkFDWnxNPmE0suxtDlqTPHkPY4bnoAmy/pefhQz+ikjHMYlZLe+yhS
PQCEd3LK92fDj2SIxcQdFsz7GSK11gP3DJGCb7XIeSFVjWMdX7CnvbGBL0ePvW56
dBWs/s3cFR3qqO/mfcizfbKWgfNVPn/vJbT4ab/gww4jM6eXyC9n0ChEvdx5Ir9S
FbeUFDzmLqAPXcqwCzEoxk08mC9OUKnrwsZtXaNOGfHjCOWjwc9FVwK9tQTHUp6J
IgWHF1mBth3rd298gUa7DR+wUSega1UCUhnLsUW/YW4wxd0yRwJ/4+afgDbg0lJt
DkEdSiURpiSTqwmbizhdgfaG3KZGr6Ci0DoF0LYjFr6muc6T8fjNot3yIGM8sOHx
sy7akfrIZDymJTCBWygh2gu+EY0PqSOEmK4xqRSGJ1ADVTUYsmRgwWVlN51F1r8N
EZRe04UzNNF7HyuDEUO9eeoLd2WVsmHwsNFU2PucuyiMM9EvD07STatWHG4Bwvo2
ozZERpb8F+Cp/pUnP9ZlNhQttv8JWA4OxDbs/SbrEVSu4Y9qhrivZIVw7DIf57b8
b4Y8ZGKPorcggYDOVIam8/yX6uE0T0Ving/fylKUgGDOjvO7vRSpSvj4P5B0AadM
vc+BUExx6eITIuCxxBBtG8lxC5LsthiMDssb6QI7f0I0AzpfBZ1AXmr1UBxk9sSP
TJDAX5hAbpdGC6UxqAVhDR+MT3wJGTeTwlVwWw9e/Iie2fk/PJhScqPNVK6d74Aj
9s9xjJNsOIKhiupJIbymU2AdHZCxSiIPinF9mqDpIG1vpQ3B9lbCINagpbVjKXd5
Mf+31FIIu0fwjE2F1BvfM7ZCYqaEnMQaKJuiD9BqvuY2I5Yu49FepkWuBTw3W6WF
Mu15fw3ie/08mAs+HSl3XMqHSUfvmRncBi7l1xiLplP6jnXVIWZYD3LrFbuptVK5
3NxCqMdP5ocDM4hWbRgnsIAjcP4sRDQvSfVNubgibvbG5wBbloEOAyixO+ra47dy
Oqgu+1nmud9JZjMtS0aXn29mpsfpR5v478TUv58mZ+itdO++fWHW7Mlb+BHuyeZ3
f7nhU9qxOegNTdJEOrSQHL3N5YuI6YsLcNjfD/qhXsw9gDEoykDKUXBtqLvs+zGM
zRz/DirAhiFYdddV7E9lpJf+QD5HZGk8N2j71QI0jCmU0L+vpl31txpDuJJ4pLv2
iFclQhXx0y2QUOgcoutQgRyHhiv82l5SV/yrwsOCn1o7XwcUed5FgXfJnO4dXVOG
AJcLqUnxyeTx8sSQ5w+CN8UeLZsE3aG9MGarCm18aQV5Xssfef0gTpq3+z1xVmBh
DKq6z7xN+fso5nZ/n1OkCWBjOhAc1XS54M5mgMuo49my3eMWKQ8aTimipqQCSTT0
SLv+CjzR4fucM1aOIiuGLWCCniLGwMbyF9Qrin2Y1YzBc68U9npTp4TPhw0u3Hk0
Jm+asF+bnw1MoboXTMoFMJLHBxlkH4QWBp8vxAwUyqzmZgOrfzDanv2xOdvxyVbY
RQSDO4EhonppJP9c6RnvSKfyKhSIanSQ7Dh1S+XSTOSkNZG+i3LFaBz2kRv/dAxm
pLirk9ljnHa7bP4Od1mM6Nb0HQSLxj7xytXRYD36HKqhgqPoLWUnlEaKIMT+V6MT
YS9dy+gIhsEVZpKWl8l3WPlSpmikzO61tZkueQ35zoSqNv5pDXOA1OLgY9H/XRc+
iPe4h/Uik0EM+pjAzn3yet1hcN+jA6ZDJvvkSq4EX/A4JD0cweg9AHcILKZZzF4R
h/88WgfIC5wQxd8g6m8SZpA/FwKj+FWuxsc5n3YUPzQ9CriC4WFt+1DR4NRvnfue
+OOQMi8GQDcDSnNQZjQTccyE+/GDyh9V/5J07ip46KGIZXaRdUJdPRAPODEhCRel
vbfuT3puzCcjHNVbeIoRjaahDooa6zkHC9Bm7JW4rntE58cChMJbhTtZNc2W2nBR
v5Zjl1aUGKgBgib2Rvwk9sfrqS2mESexT10RjpfSPXe9pk5oVryz3sMJ8DgAaKxz
V9q6VbyRU8Yc59FuZypx95g6fzCpF1CFOjL+fp6mnYqrDcLPOwAlXFT+HY9joEDi
b64DxJHbSrWVJwCKmCVuSzkUGD1BERMIyLJ8J1f4zMa0i5UpAnOz0rBxY7mv94zA
mdveY7wISovOv1Pr4/UxJimuP7y2Jrbj+HUBh5aS1dDQkfo8V1Jf45Lw7YabKxr8
E35og7RAoxlE0428e2fNIW1EQ+mBUtpes+48JtYilrr98xG3lGnp/ad+j/nJWlEJ
SpsbGrRPgFRgn04nfPvWr2QWRGN/7sreFELXBPyqfcrw/ROCEFpoh7nF9/zVOvc4
WefMWKC/8bPLbfR5rfC1xqCfl7RT9Jhq+7S6qnQDphaPb2Gz1Y7tbdSdtFbGHHsq
K/lER1+L4c+WGRr1/jyKkL+3kDBuIXaxnqLpsWtGc21uzIYSXypkGoTLDoSKyjxF
K6bifGDvpg+mf5Pj+uJi8wNzE5UgcPo8zH+STNKAN2vZxiqBcZjTE7qxUuVYqNNA
30SZUgSc+HtsIFWSY58IMeeTz8TrHIsWGp0vaFZ1tAFVQhlNfEvOU9TBUauToS4L
k6oz8t7B4wSd9IDyDyEHSLkypCR9njUZCPuCtFZxrXqr6a+2qHWC6hqoWhf5Ef64
RknePszSFuYep9wdg52V9Pp+39mmQm04b3j835b+h6NoMc6vqZgNZ16eQeXR6xM/
FTG018YGJ4ZGk/hO9E3d/KpT1/LMMUmmqHdtSGNRuYvbrlbLZjOg6oWUVTKu+d7l
8jBY5/OEM5S7RgYnqGEEyt4S6geFurE9h1U5k53nGvi6xWILbyqZnOWWQRh/hnOL
PaDexBIx7vt8ogO/qwsdCdimeTG39Xo7Fu3edfQNmMP93tq5Z71zTdsGRRtsnnju
KrU3RYwU6ET34ExJk+ZbUvWgLxWhLHca/gCtEz2FW4gageF2CS1lIQhwRcr/0d/O
piLYUgc1eJ9nfCAvn8bTli3mFz5Iqy7SBzo9WbMt2WsUNjXLndWasfl93OlgFOSN
JerRduKTdzeAdQc/xJ9nhDcGQoC9XUtxlZIdjZ3/81VpuuEI4GA0d5WOeIJi2Kxc
h7IC83mDUDP1psAf2TPBo8+kFmPrcq+mKNa1tmhWyhZZ5sssMfUH690C118mtf8r
AooJgX9GDp2SmBZk0UJGW0P7FfrgQUX0SvuZpJAeLEm+1EzbYzQWgIIGsASsNcyP
9cVxXdFEMGjW+PFQHJeY1aUUSVnQLAXCEwka5N+1/9iP2703kQqdv8kBAIw9rVX2
L+IyefhXwvyor9lJ+l1THuHBLaGXJHzy/EZUoIhYR9IMNUSAbEOnsDRdeiajM1Ew
n+ctJIP+YR3HejbBnKd/IbuW191ZY+B0McyorrrZxjVGJ29EyUosbLt4DDa7mSUi
GQVOaSUkjjCKT39T1g6xz2JUl6fI/plrYN9fsznrU2ROuW+yRcbsA7/W6WHZZcLO
1dg5cIB2/UUC4U9VRwFbI1UwAnv6FZN/aDB2XYSJOaGBDfeVEdx2FZ87nDQysUcJ
uLaOO8zshPUzRYjrdSqa5guM8Gc5TXJfmkC782BOgu88noGJf2eT3B5XeCDBl1Rx
zC7IFnMKVSYRBW2aklW5pKbJ7SucyjAY1DRh7KHhNDzghA1JOWr1EsA6HHiZ4mhI
v0g0dJo49NBdT1oLD4AoiSGufR4QkXbl3x65O2W8fEKJFcxhmTQROXMLo6+WjZEO
Kv0rOvJKNwPHOoBnCRvKl5yM+CXTw4zALiTXvdDV6eb2cBSgMQfHPUqEJNO7C+TK
Wt2ECWrjsEupuA1mwTjOTiaDSdunGwZX/l/PXv+2iCF8+5gm+CJ9DOL/KkrIMuK3
IuQj/Hl7Jrfe7QBlk8nVfvG7KzvJc4Iznes5+UIlMEJ9qfUMlcDiRz1bW1skI0Xy
E/zAU1Bj48ntILjVk4R6fas0Q72U01COZPsHU+uh/2bgQdShdrcd5I+X0B9u0qwR
lM3tVH8xiVN9eZygsOs8EDK0gwFmFPIdgtIaOKW3ocWkTMXxmOzJuQNXH3VHTvzB
xJbtecwkn3ZLl4oajsjPebUDfnKZ+7s09tZoJKyWPzZhJYSgao2jqHeEs3g+VAVs
h6mfaEqS2D6uqS2d66/F6Yj3QIsyijPd2J/FDiIj5hvpeg1nQaAomZT0TJtz0dRD
zkgr/mKtW6XHGroBn4/MGcgXv8vu1qLtoUhYaZeRu6KYxYxiwnWQQYQczZW+ygJX
+QeEIKJ+ERbyOgIs7RuF/8f4BVWwQV111POHZNbrX7d1kN90eOB0AgZIY1nPQzWo
tvKIIt9hutL/Ah4knWesmZ/oaZ2pz7oSqPXChqNVACgf1tGKi4Z0n7QaNQe2tcn0
k/Eb/PrDYE17PAeBHcAfQWkUxDebR36iZ3W6EM52+WaOLXRsrTbVYxPniHRwK+Lm
IWRZUPZBqK4kWHk6BjVV7cK4FRkdktCOTb9a7iWx41l05EhlL+M2C+TrwYkND+f3
zgSLVf9TOmoFTiquSHe+ElppQ2fs88ybaahOmfUhND2W330QBAR3FVPAM/7IfjzC
AFvQ28VxJ+M5/2xvY6V09EJZPttci9QlEKh+niVOLyGEZXZIYpEeIKr7mR+az1RW
xwC0aF/KbSapnfbOpKJQb11AyttyD/wbpWsLXcIw7uHtSHaJYXQCLeWv0RZYZE8l
DUjKZEgzXD1qkNnvj/MsixK4dVjiBxwxF+d9bvQGMslVWIDVQJbz7sldyP8jx/2e
RjB05oQ1rsaJU8cYlsOICqh4qEC6G9WTGTG6mPQOhR73p/0CPNPSAKAHJJk9IiCk
gvdhe5EyVKBVGhp2mdPRaHkD0Wxxb0pEkULOOOEmOJUDPgWsQxM+UEh8GGh7n3EL
Vlyy049gNeZiOdCiJsN5Mo47Llp+tEheImn2zQcUzMdzRgPsU/+2u9WRTWV83x8C
OxhnzT7zySy/OwEx9WZkQhkN15qKa32X1tXntWEkilY6J5qc8+SndYEqBgjKNWX7
Z/IqD/EJkKDzj5xz+7gI27VOfmLXI+yHZ+VsEyUMDfKFbgrYJx2XqJSIumm4PaXf
ZCq/5O816zqwxBmYMhkY2dj0A61Gz0r8MeEjlhlGT9wq4oiwpPrhJVRkBUVW7+Cg
GQqs/vrXAgUFnINesvhb23kmlZrbuWGi05MVVKuwNk9DVBjyA7K+SdVyrXLhp3vC
Rn6ODYGE1SvmHftfM+Gu9Q+qRtq/49JJSawlluXcy5o4AFRoDup1JJ33osikSTm+
gK3SYK1NtiPRM/oe1TuTmeELqpVVIzrsexiAWo2JY9sfvLr6ZLRRGkldov+tZzi/
PaMonWfGJ/U1S5PsliyHFLEPZyFQ4BOF/8kMzxMdEU1BHYzQs15sjFqaFhENgdeD
szhBPK/LOZMxX8ldrYl0a82/++0U1ncaFjyifQIBtUBW9POuhW8NMxUVNTg15nbj
/bq84g1Nt7KyuKzGOPY3i7fWQjCGwrm94yZP3UqMuavobTM9kAzNTAQwGYVEuFOA
WpeB4VnMW2189F0SWZwpRaBqtntvBGhBS+n4zRS7vOK5pEfDGJoc1fQUE/LSOkyM
j2rnE0NMp4AKq9L4m1h6v5E2r3LMCxCfvkSBkXJ9+/pmVI+uBCThv2VF/7NuwCK7
vY9j0WHd4rJ2uNmaApGI1xnYM49v/24yv8YMuivUpC0vSnQ8nHbluMiP/AREKzkA
CbpDRbj7yLY2kvAh9giTYK0A9dYiW/TLoBWJsMYLEgmC9xMMn0xovJ9i8nRQeiEN
IoOYFNSG/w5hi0GcTnE5GBGXCJcnUq54avvzETsav4FrloxF7KNwJRzNrxPVAmSl
oPCJ4IY0OvRfMNAJJag7ikZNiugCIx7E4S4zb+sgnndYLcCa6/qVQ8tXjA3MOG3c
7p0dACbB1UpiBxpsgGIcH0tzgidR4OmisD1BRo6A5SRXcm05Uaj6GgC9s7VjipSP
mWPeNui7PnvZgllm/cDGdYFLha4v/qW4s9xm6CK0x+/KJMTe4mElTHickYF1PrsG
FRPfcHZAFIkpA6JwICNvlTE2caOij4hi+ZXUxGgImyR2TaS0PvClJlo8/IPNuTjO
a30V78Ex1o1Uw8buqEZq88NfHPbXGGOUwJT/nhK3Oe9gov82XKvqsIJRFWgscvDl
ENH2znF/xcdg8HRdve3gZHMRngz/gg7oBwq91dcLd4tmmyHrF3cHRSi9MMxAt6y2
TtE6YBg57LfM3Pw5kR1RkZEXBukKvREl2L2nvkc5b/SlfB4joV5xXKLZcW5O2HFC
zVEswGXec1XbywDlKcpFz40ctdUPRJs+Nfvu8UuSGlI6COJRsghvCvIbzThx4t1K
VeaFy5+5OgtZqVVtukbFJAohdrzbO6UOA2UnQV/P5QAcBKVPYx9yXwaA3XFfp8HY
OxTATmOeTkMw+kaz+nUK4Qc1Fd+tG8bEf/Yp6hKBF9apBubttbG8loYQagAhYDhK
G9He3f9DTpPUY6RRHOx7jto/PRX77PGHJYoh4tW6AcilVY/GpY1ACUz8/du6EJF2
Nhx1A4HsIqaxjqsvGL6GBK06f9EBiWtWMl0Ju1CsYQ6ZhxqTn/anCEIxyOi3WFge
v1TMI2r0s9zRx/XpGYfjrly81GdEhX/xehKM6/z+lsHksi2XOim1Ix/fR3WIpqZa
aDqer06ocBMM9UYl3t0D8410hXj6N17PfqXqFSMqzNX76qR7D/M9jGKOD7kCWPCG
SqFUYjamXmz6I73nDDEatdq1VMz0JnISrIg+3gEvxENaRki4p08sinRiACRYELAG
mjimVfzrVkZUzieCRURzuGduCwT2wEF1S5KHQv1x1z/olrzQ5wN4rbrnddghDlAe
OGI0CDhjJFbafPtBNxvKQbrG5BfiKZh6J/LsgscyEB7lbmjY6CssjrLMU5AwH+6O
CIDDC89kU50VzBh9YH2ek7Pq/ShSwKdX8MYFew7ce7cf1KjGqDdmvCcGD70EEkCr
2R/IQnigGfa1CubgQgioeWbe8zWDjMYdo4jUSeSXT3Frd4LxetANgSjlicJg76eX
53kXAhJVb2OhzPnYf3pX6KHQ9vmCT+Ki3K9+nXD3W20mOhNQDfFLQ8AT0pS9XK2I
MkgbUtwLzcYuDvdrlJ01WIRE5RVQQLD3JeqEYQCAQAFQg9nEiR1BpkLVsvzHFKo6
JqGgBhiAebgfqK3YLT9t5fGS2nhcXhN8+Je8fQJwattAJHksuYXpjJnu2eQ3on4x
Nwj0lozQI1Z43UAmrQhy9Plr8Z6mzNTff8plaKVJAxBxvuH2ivGd7FhJ9ZCqRNXF
+PrvRB958eaXeI3BMUKPkSinzDZcqyZTDyQIwQGrm5tDc75mTIC9cHej7Z/ZFiy2
nvnFeVOyRhemh4hR8Navg6oFIg1PNiL6cwRBBw8ZZ7etXPOEC9rp+4kJmZASy751
ua96qLNgDUwDE5m5pTdH8LkSIuUOwiMjgk+YF/hamcryvwru39xLgW47DvoCnGKN
ZSliNpgoys2mH6+ni6WAKRGAqgBqW6Kh0QwB9rdjVFQ5yiTPzcrpxaXp4cODP9iA
CBm1Iejkl73Qq9/28o6XDgwDpYnTHBRBGYPRfF7sT0EaGMqjF0a1JBJ0f1tduQhU
cb0kanPzo4RO6T8somMFu3wMFcLDWdX0EQf1JecQMCDX/bSXC3dPS5gbwOhGBFN5
jhkqaXrhJRy11p3oOwGgYr36PS8gfcxwfgrTGAemHjxxk9LOEtPAjhrAZsEFuYkJ
bHE5C9qhU8BjevSPbQO9ATgFtcSRYPdbBjj0ceq3E8fYdGsyCoZ8t0OzY6/YHW9F
TP/XXPHJxHISrvmjJbejmYvHRBoiWwFavJmJDodDyX/f0vryndQr2h7rfRGwXtQO
iGjgma5Sc3BD8fTO0LrS0h+CP0F6yEMawtlz+5iP+C1G9RsLLp1Q7rPVM1jRe16W
Rl29+t3P91MSJnJ+JqyUEnoaV82r6EzZHIrzacWKZbG+3gn+RB05QbQ8Ud9ODt6a
3r9iZBXwv53z3e/aknIivu5nOeCoG6zvAIJJ89JW4JYl3o+d+tjz6CxIfJ813yCt
sPOOpB0360T2uDbFAafYQYh2l9zY3dwnSKQt3TVI8a05eob8Il84bntkDZE+srRE
UXAaiPxqmVO7By8gp40cvAv6/Pu5Xcl31e956r+NWl7m+IGifr1kXDYj/cmztPVv
VTZGvqSC74sdhqmUypLE94P/T03XVClrr5XNxtV3k7bQGe0tJ+PmurMMvYznYhSg
sdZvv+RrADyVUsWxGs55rTvS3R3yNv8CQg/Tv1tUn3N/1h0lOMU1A+0yuj+93L6X
ROAiI3AlWcfKXVqC8b0Mz4rEulqzP5CQ00ng+dSHKlwd2WzfTKvxt/ZVmKjs+7xY
KIKjgYFnMCR0WfhVqJC95VDivnWJoqmbe7xlkiFhMr68XQnRssdIA/pm1anDy9Xs
DNH05gpzARvKuZl1imZhcDCiwZZoQQRxcp+yv0aA+A4Ye5//+gpYR+bTwJFYrwJx
d+UWZ6Rm1p7sLJJVwfv7z3S2S/jX19Yqnw976ipkmYzisEKiKdYegZQW/8uZOCm8
AUk54kVZH+cPogVbh9azGL5s12oB3sku+XwovfTFzfv3rWh71sot8/ctNrHybpRv
fBJncbrKghrsa4PpvH/w14bpvEosvhQ/N29swarRgnvdp+7g4H3w5NvDKnotovl3
j4RrQ7CjpblmqqgQTSNFJ5uR9y82jy+WTvyG0EdzHYDKaNzKZUhGMvIknFN1758X
/ANIw3uw/AaOqyus/T1ojBkNzM0UxQoGpfOKUyE/yWGVFt/LFQl6Erh+EG31S1IW
/rygZr/Z3s/YGgulM/K1x7VJxuyeG4rKNDuOU2jdDtKq01kOzUCMBktNnj3VqCU2
KNtSwmWQqODHyp+WsCKikGOQ4N9yvb5F/wBqqusEiryWSgoRuUuvpP2OmrinOf1F
HxUz4KFZIFBar7xOHqhSDHAnIEuIvmneu+oAaD3lIXRAMl/auS7WYItl1aD236N+
ZRio7Fnv78SGjiXdqzA1T6KLAtUggEg/YkG2IWM0DUiOU1OT8AQjKljfQ+thEbPG
HGGinovCp8c5gRXmYl6kQke5Uq5u8JZyOH3dGfA7vT9uM491IwTWXeWEt4u4zxIx
avUsyyrux8zFd1vd1qbyHgAgTtf92PY7Hqm2hUCEBIPglTOawJy/fHr5cBgfmowh
ZiETo5Pbs03h9s3w46KxbMo8dhb+3/ho1g30By2C4pSawhwU6krYRYib3EBvehwc
1mhdk8vli93jflw3wYV6TZ6FuWw4aJ/Q/m/itLPn9cMMDcDiQT9UzxD6EagzGLZD
dH6buFQWvNc73VkXNkXlYDZqBBlaB/eXizKMw7tZecciEh5Pl+2uSN2nuq5YPBSr
mm7/zyqu08ClZE8oT+BeHSxAE6/2/nvFq6iwvOIW+NCj+N62YrHw5HN+Y/4TX8m5
67IdiUIRe5psHmfj2GXiGg+EZz3p/hTXED53tLCHFeV0nQOXdb+ysNaQ1gsk/gKf
8WFyMIcEzOnGrOXYHiSzxol6jzI0gYR5qR7q2Wxdm7O2DgRMziguBxGipQqEsGFo
j26MAqjs+NDDXtcNiasTCpPB1LEro1WjLsAlhG8d+sEBIqgREAhsU+o57S6Trifc
kfibJYlgBrlGrW1SKaBjJgrLo2vgOVWhDd9OpyR1BtfY8+ZBesET2BGmjSiEB2Px
OnkNb14l92JRjTxIXRydBgov98Tq7jfHfKBFZY7XgI3elzfKF8zZ7Y3wchJ74BIg
c5bpGrfyOUpguTg/7SBDoUWFwSmbybm1eAwKrFg3wREI8Kn5jUup/TpyQ8OC0dDl
6H4AVSZYSlPmnS7hGpj1COFon7owMTTK11qZvZdRreyd09lmgVwRJrp1pKRGAYrE
u40d+igXa487n7J8MPaVIodF9b3prWwDgbXrpxP/OsJ5RrdzP+3gaIrEd/NS7OUL
u93P7dBR2epqhrDgoNi3bHt+CD6xTrh1OHOXkdAd64vdscX/eHoSNZpV6VFoMXAk
Iy6prco7C3ncoHAq578BknP9p4Z7UQ7WJBt51cs8PfKAgfhZ7BeKxIqGGxiM5Nwy
Jd4jlCNdbR0ZwPsw8kNNUb5b1G91dCiRaIbsD72k7UGSGeD3unMpac82TBv1Cvm9
Og/nSYxhBYRyWFJtIqZCYQBLJttv6quVEZpyuJ/owjAT9rUm9ltCGvyAXMWWWkJs
cohLm84RPi75+zRtd0rB4uUueTJ9bweuj1WKKBWP4DzE/IKPOuH8XEZ3isc78l0j
ULoVb5DmwnVe47AWE0cVZV/9nG8trTsfRel06D2/KhPYQ3TuZuNJdFuImtQAnJKT
u+et5AErLsN+u4aIWY+r/50GKNor0FKTLyQoA3eK/nmGSa9H0rd0xS/P6lk0ccIB
48JRr00l1nUipTaiiNZlRRwEMkRnc9DNvikXw1L+JwNWXVuOlMd/26mA/MH4WhMI
mExmzKgqXE4UM6sXXoqJloiJMTvQowRGCXUyUZ71AfhrrnQkIbVhx1xoa8Mlzfj0
wEVg6+hCcmaIlGgS1LT9am3webHvAyV4fEymnNl8Z7PTkHmdzt85Rw0x9Hj3THj6
Gp6PDZJ3lKDTKBFiVPjjNa69IkF9G2n4fGfAAyhZ9GYWz7DBeVvF8bEUi3XzAwcQ
EjSmjrWBkL/wFbPpOsRLVpcPmGZStuJi3SnRKWOtpYoRPWGakxKMjNBj5hdrSzot
K4DBjJSCK8ovzEM1P8rqp0JQ0IzAmKToagJp0zzrtbGcwRUZM1XTEU649jiUFlel
UFwVGOUs8pCLyzlBh9PdFDTipLJvrEhl6TIEl/ui2itNYvIJJ1D6EhJtfe4tNUjt
xV0PmD2rYWYyizmlTOj2O9KbSBAiA5AleXjkmpQ+n4p4ocxJU9G6GvVDKwT9AOPv
bLzGEpTy6ItwzPKCYwWJd1I1wugvxaDiNwJR8KXe1mRMh0bzhlymCnKxqfDVTNDy
zUqmqxk2kdmb6Miazg4ClBg2lxL4bRuwz9sCkIRQkRNYcmuZnjjk8j0HOnJJ5Nsb
Q/+erh+bg/TGwLxeL/b+CBn9K/P8MR696In45TefF9UchOoWqhbO8ncJgg6Nf7cf
NME3rjO+fniwSi/bAHcgS+pPLyD2UfpCA4OerKDi+3REfaE2qWRR+qDzn+U7ixfE
87wRgaIB93NOzo0Dx9t4GUOigWZPehX5XytGoS54kHF0dLT1+V6NCK2OyfMIiKBN
WAn861AESpdAbms5E14S0EEjEb0R88DsEOJVGhJh1Jv9aJegydo5NTOQp8GsEs8r
HZaqkNvJmu+PXbBVa5Nu8+Sayselg9SjcLxHa3M9pt7Ci5kvu/F5jse+3AAXvoU2
imEroBU6j4swiA9vtKCh6W5FR+NQ6aP+sUxe/ZUXDWRqtRQHv4t5uEQzumTuHuby
8ByJmQuO8pdGW3yVvyBeO4kOGv7KSA4pcRZIg/1wye8zCmjBAG2VuCGkOqPxDAWs
UT7DaXYCxgpYmAZq4LGGVzLA9+kbfYZFpbuKxfHh3eSjZTz6lvo7JdNUeGCgic2e
aUkbT7Id9igZTdxoxHrtgd4x5Dk+pvE/2kHqECyAgVvVARz113guT0jARdeAjZMb
h4PDOVZYlGb1hXB5GDCs85hQKc/KGhN/84/Ybf+4IgjQ9plaXfY/JJpnTMhya5gx
Q2Kt0of6IPNwzr6I+qKiT7+mRfMw3DIS0BLCXL5Yknc3D6P2a072JONDpNw70M4/
ihdSEI0/E6bq3A8wpG9JADhjg2LbiOjzKs17RSsiNjA0zvL7KYLPTFaSvQZ74P5S
1oEHGTaQ2Mc/1AHzNAxIfS0aKwqB6MNFYvFGXj9pZEnbRh7xWp6/o+EyDcXfiBs8
peInHZSHGpWRHQkRC0xFczj8oUDIchPDSFdQcLn+DolqT5ZgjHtGkjN/SKB9jruz
ql8L6LcG5sjudU9ERyqpj5hrlTkj2R3fmfwlKxmCtrxiSJt/nL5TF22d9oSmXGoQ
Nb/ACHSUynSS2GOQCMsq+f+Ngn9gUnuiUML5+DENZ1hytEAw9KtmLU5uQCNrC7h0
XXfsaMOAlSXgX8z44ReSQ9fIIXScGuaZnzDXNLxlB/3ExJa/apfg5iEXkAUh7g5e
So7RGyhZcdW09ga/p9hh+vtpxn9xQR+mV9QmXvpE/dkIHbOg+5SI2EIuXdxjAkfy
foUDrfFilmudSzHoBEklrIMW5LNY6mdA/r3WYjpAyhBrZbWhYTBJzMNN1ljsLLkP
h73paGs5TmFDoxhYeGyZr871vnZeA7fSrV+lvEngZL4BVJFeqoBPbz2JYRV52qBP
VXBT7hMeAtrADnjck9swZBiTd/wcHBkM4nr5zhwrNRPkWF5qZ2Nj4YYz+l4CRvYu
rIJ+Xro+hNhph4PlZVxyOJb6JpQpODtL/VgTfRSlgA8qSVI+Rxt6pYZrjLE++wzO
lWFU4+o0UYgv46WI8rMPaypPpD6dDKmXX1QZtPxl1fNiiKB6zs9gXeAEjCLx3lF2
loiU5zCQco3DbzT4Y0eWJjb7UoxT7BDXwdaE32r7oZatJKEJi+sVQ7veH+9o6kWV
QvQNZzX+qfWfwt4JPGgeRe2+cvt7eGNK83EWGjkvubY5F5uBXQOaWUEuc0tgiDxi
KTHmpyPHn/XS/h+ixRxklQp701luU9EbGgelrEZqLQcDb1LbR4PXLJT1YmZiiGid
rCDgXd2pAhFeC04c/BbGRKLZg4fSdsDoOQ/0f6+EvQ2t+Uvk5rChG4cYrGRGP8rQ
+kKtEmw60aKwdPb3NbR48efD6tLwrlEoUPj/YqN9pnayTcQI6tczM4ryxsmpQEVb
7gfXn/rnrTEwK0mqRcWzZr1qoX9Fz+CJ71mF4gTgB4yuLMxJMTeTHlqbcaO5f33G
kVbI4ix/kUruN/P0k2qmWVLBEioUQPkJZli5pBecosWPo3gvTqCH+4xnzQNd4LKX
Vr6niqFA+TsKpfKjMScMlaLpKn81bPldy/K0dYzG75lfFUnH43RpRYHuBkyxN2ve
mjOzF4C8MamC1jxanmFKM1SR8hztDrn/780pHlyHqCcXp/7Tb7ko0yMEpO/aWwpY
ZDOplmGzWatfycHOktvENNPxYWwCF8jer2mjDsnHBK/ut7EXVUeT2cXg3z3MHBBh
sjqPT+7BS7eBWHzCDXxMDqeKoxlhCRGxK/+bFJOGmzZyNHbS6iRHD2WD1OKNmQ2l
jMv8WZdsxg7KEE6sykqNEhIcHbAmI2Ilz+DcgPloUYKS4f2IYYMJ5h73JTPKhBsd
2RTSs/oooOpTud1OLyYTe5YRF5I34jZtNrG67UaTBWEpR4GtwshI9YmB9C0/q6Sp
mK9QlJZsDUkKAHw8Cxut0IZ59ID1bUrx5TejTOvdK0H/c6UXSSdAvzIaZKNa9cNA
EN1Xx4wwkC/czFxLl5DNcnCzx4rekrMAw5uM+X+jojb4w6CTa/Xi30C9Sd1SuLnW
pHNDX8XfFRQRr/1nNLjubwOzCMg3z+k0jZ48VeJNjiuODP6B7UH31MFfOpJgz3y7
peIJ0rqBFZDCLX1in8UFwy5TV7du0rb1OQAWswcmKJ2RZasUIlWGu/Z5DJXl1AeP
3cXkESVjmUJ2TK9a0BeXvD/snIq9zLA30mrzvC7alsU688oGi7wmFf3PiWwq7Ef0
hm151W395VGX7HdfESRjLcaQK1jN9Pxkg5iyycSf83aVm9sMbyJcSoU/VablxM3w
NtyrZ3SmDFjG0IvyaynvUiGirn2cXGk2bDx4/8dEcZEeQUQborfYNaOUsYqKnGse
finZb9ObTfmGOBceR/Es1fjUKryx9ADY61JekFG5unOrQMzrJA6i0BNXEfVvfV3y
Tumm7IWd4kdXgZsDfF+VdODDLSaMko/bV2a3iu2kBgvHwfOS7SLQegRYNWGCFSc4
8k4CjKA/PY0vDThNOV87z1j4u3Fz7ghWm9OwRGJqJq8aVLAOjcjaX0Vje2DHygEJ
eBGq4qDU/BFTG5zwjer1h+RmWqfPxYay03ToSp7WBz4X9BPwxA4sv9zZ+eoAGgia
a+qRvljf40gZ+GwOsSp2EdaHkHpnKb1aR3K6wfe8SzRFWyICUFg6NwQAkEHf5BCD
WSvKo5GkRNfQgRge8EoExV5JDDkSijh3t2Fwb3H8NdD8Xe6XMFZPb0MJDB7VkxCJ
vkhaWGFas9G5snIa7IkfoD+/to5IzwxqkJIs1yHzRsfpXowU+dAypWJH6LTyVJnc
bZXC68QVUZ/51RnNh5hlvoOQt2sUMvvNezYUXIXJueV19Q/mfhIVTuqHdyEW4Cze
4cfez16SagyJ4HQHCWQf9q4uEn0UWjVOliTYluCCv8Jd2NpU89zBy8MDFUdqEUqa
NXr+9ua2u8dA4C+yPthUaQMbG7e133RkU+lbsy2tAjuhy5CvSxKALWGDrhbG8Km9
jhRtl7JNsOz2IPTkqmwTTK38yrbAwNEv0Nkw4xbQw5lV9bkoF9eq+lFa3SOpAA15
nV1eFBJI0RpVvW0fsms8Ya7SqpTQFrSy2xVq6gIiLns2ne7RXhFWS1V2oCGVFUma
RfowWUKTYNGnHzVv/U/yVDiJnD/QdrpaRKgjAZipT4hOAa5Wf/wt5UkkH9QWbHpk
GeU2ti7N1dn6EOV3P+FkDBh2UDd/kQIEhflm/K3cqZYFexZ+TlcQvurn1fQMGiWn
PoOpujnJ0xXZBf1ideflCrwYQeAITpq7evKLzJjQkT046iPGyTeMXKTSGANxxhEv
s0h3zaQgtA70RyBQw4Ehj2siHNsPNhXtMXTRXo3aSF9xjq5nkj2lp6JaewvK5Cab
Nx0mvPl4pBfcwT8CQTq8sHWI9gZunjFC7UFWnmeUBkFNEvZoyL2gG79sDpJPgTaA
lhpJ9dgXsifpJYi7SLnT48+qJfn0BzQkQjnG6dqtwYFhX5KDNbhSwzaWTxg/ssGO
AtxGhAZc/Tthnc+nxq/vy1XUxSJd1VnLmgzw7PTjdneqMXlJrlsP8NlPPUFmgK5u
oOYTRSdFPlEt2c7SEOz5p3s0lxuc178uXKFi2gsdt/bkpPBA8Wdul+UDSSO2cAB8
dZIKsiaalukxH0o7h0v3q4QyKUODw35VfAVthIFYZ0mcCLh4pAyyb0nbPoTzF9rf
Cpb+NZ+XS39fRxgXho2jDk4GpolyZ0YEKf5iVKUCGtaO5mryrZX8Oju+G4fYx+Pv
nLf9TVht+cDOwg/+Vu/VrgrQZQNRvyCghIeMyCUprdhQ9/MTsYqU1SVTiM82auvr
rUxF3pv0csVoYL/5+K71KfjDrz32XS3A+SL2ikc+NKy46PRnzmDttfjjpR1inQWA
RWyCjh13STJRgfhCv7tgqyeY8FyACCdciGvaYyVMbs5Lx4FZbBKmuvWtvhtPKBiV
88ggUYz2+F5Gtar/UEt4PMFPvLlRrvVrvBFQLCNRq9MemQro20xLedxmUNSyTUcf
2sfiGALY+lKd6YGElOvLrtNGXKRRfsYUEOW9EwdZbI0BtPoiOqHP5HigyQx8451X
Qgg05SSWE7kDJcEXnqaLLIe0Cf6OKUQv1kSYo/sblyPAtvn9rvt7aF7fTn0V7vKq
w2sTjP45Kp6lfJsgIYBNe6G5eMj+0UTfDWuKk1E5jyZr1+ovM+ZyOQUAbxv84J5H
lK42B1CAlXHqMj4eVuiKLfRkPVzkptsalObouTymgIt0Y0iu5j8jZnhD6IFVjPrG
I4sR2fHvPMcgQrtiqX8exsirSJAp2o1IF4b8Yef6dwV/1HafqBxw5qbwgCfl+/B9
OFIXtw+euXvE3xRCiIgfmFWlWXF+1WU7kZ1q9KtAZi2WTdB4IPs0FEzyzspCi0Ac
W3wAauLetR/CJS9aICkSb7KjX3WH9rFLgClZ6UbjvKHsBvj7uBx1trhZRine2UUy
ZzAfr108v9AaRl6hRj2MKouJBuDuQDqxYp0XD1nZgkwFsFXDdYvsNbKRflJjON3a
8OSXeheVK/SFLHLEL7px9Za26iYfgZIBVlk8/2i4z/UZ7r9kCyqMYswlxrZQbvtx
L79FIdIP3zYigRY0/VedF43+Fl0H3StGqSfKjkgMQgrSt4F2rEnzx+nESfncuHWe
cICX7QNlTDTODycMrXwLhlvECJDmv8uQiykXSSrA7niFY8AVj3g8ZsVDmWifzWvs
aIouZNSLDop49vZntbgL/AfvYpw78I3bFkhlaG0OtQ/u8L7qWsZMCL16SnQbLfZN
ax9GRr5sHzFqSBbZfXvO/BpNjVWgrCpNVr6hwn+xxQczQjadZxnLRDoGIQYhS4jG
eLs3qshPtcfBlz969WjJsBeiC5pQi8JisKHyVWgqncpdSp4bF544nVg1aeHyLS7A
g93BCmPeoiMTrR11EH3ZFwWeYFYKkbRrwqFHGvy/x/Oq2cwHGcrf1r/mNaGlQZJm
HktVKSHe2b42MQtJol6Rk6XhYvmvd/YGdE+ZPst+nPFm7FdUqO3PJSZ6FdFakJxq
Ndt8E7JduXrPdg3f/22XATWccUinpZbYvA+iw7Jf6DsCru04Bf2GKWJ4e+NS9ldh
ByCr+nPZOZsWjY89I6lW2dqimx8rljy3Xy5XkUPQGO8/VstruxDftMxUIXeBl4PA
+LUPToKegD9q3VdrrKeG1S4b2SuuEFLVmvh41/K1jlsYsDXw3f5J11LC5F7zmsAt
wKeswNNjE63E4u5PFtmatjZShbPDTvmUYeHpiACppsbSh5ukFtVXrZaciGWH5bK6
VOlZzf1TiJEUFRnNOiqRJB1846XBLTKhvc37AnpWIq+9HghWvXbx+htebbJK/q0J
xVBm/WMzywe8NfkUncbhZKZKj6T1QaPZubloLK0LdjF74NtUTOycf83UJPptdPIc
5nQo2nMkzl3NNrW3V1WRVt9fUZKSUMXjtvGeIvOv09ViLw8mSTFpEIwPFMyXKIan
Qmv4soJyKjeVNI54J4LrXWdvmYN7hGLouA3GMqeSVok9qQ9Y62+VCB04MfocQuUb
KESbFh41iW2BmXGmOkg4dPDh9t93L4sJ9qdMBAXqxhwGk9R1QvfyMXjeN65/BJAn
SCQC5Jd7D2ojus6QRgTCA2YXRD1Pg/8BjQ8rHMvPdl27nWDg6dgCei2+sy6JfXaj
R+TM+Ffi9hVAvFCaFx7rXE81CVqQo3bXspmw4kL9QPdvwD4xlyKIifjuKY9Mqd8S
GVMRuZtfI3xg5xfdxy8SBz7Hxrhy9FrLPGHJm8eQQheJek+vS/Vif+Ht2uV80TDr
naLAtdFFrZ36uDkgT3+2Na8Q0uwZ450OXRQ6/PfXb0nNXDWaWDcI2Eg6D0SUA1ub
jnaAn4HIOcMRO99zZy2BiPmCSVkGZE3HUcoE7fSR3NayBSOY6DL6xWiZ/XqDPoVS
pGbXHefF6rTCKGsopFJFypc/HtHbsjWnH4XxckOp6RvF6EibE90W5pF+2nXouyQ7
K/svk8pIro4SnHBAZAqpQwAOwyfj5sKohX12xVpY7hHsCbHkejlkeQVjEpc32IQd
fPttasJTnxQTCakzHjaMaRDF7FvLWPNmmzBNb/LQVlq03vYGtacms+QumEr2jaQB
eXuT6R/xFVSeDg2kJLr2J3NBs518pNKziqTuEScyENFcx7J7GGfZM9kcPpdTZFUE
z3FyBJ06+JBCCDB+bCC2EuP+E7AbgB/n4wcqtlhvXbi5wjwhxp80Yr6QJMIaCyF0
RuMtoN3XqLBBqVsbx8qJFiFQ1Rfb5W0K65LLKEGAGPR3WoO6NZoInUdjKPsWiFMU
S66u3A1/gWY7PQ4wPJIzdURYofg6Peax3CvPe9xI4UFeszUJAPtRGGj5QB7RQO5j
R81jCbIBLfFtAWBTvirPxWZPtFAuRwgRoIHCynbKmX8ZShnCF9sW8ckgW0R5XSn0
SvTe9U2qG5fW0uxJQVcYsUJS9MQ0FOIcmCFydi7Uysn6z7Kr4epJ2he9PxUtYxFQ
7/qjprfg8FVneJ6in88Ttjw0+7QM9XkxMxn4ohceziPhhOuin8x3cNRrleFD/hns
oFoNALJMuQfrpjwyns1K7S/jisX4C3FkLcOoFGV05URelEhmcfwElqeAeT+xp0QR
T+XnOpfn4mS4WGXD4De8mHB7ekYPNNZNqrCsULHlef8YaDpnAvACcPTS3dUp+d61
eib9SuQNoOs/KOxTmhFZO/C7FnAi0134Pf57lfbdvTRYCiizhddO/0M5RRRLjzOv
EIGvou1J6GcIodLgmpZtBryEMmno5H8Ib909ehVxJXxeg/HNH8LPpEeJHyRtOOrN
RGGcRQ0/TzhMycHKSsbIilvJAUUE/b8zsOSiQzn1rm/Hq5oPpck+tVusZxFpfKqZ
0QwLXBLu23PuSToplwetpCLSf7R+7s5VaQcdpq0jnnhIeKeb6RtfAN1c5yeACwGR
4llIs6MGbLNkX/LTvwa3aPyBT8uDCtR3mLVRFf5wYb134uJDSYHgSi81GrIxW1Tl
bwts9jwFzM7VfStIG/ylZYn/4DBe3serQZUeHZ6tPd+dzPRiFCJVWDHwr6N0Lv7j
6Vr67A87XMpxYFiK5syItW08WNwrW0jI6qhnD01Lo1tral0XC/WvAH+oWCkWOmsX
7X6+vuibIjdGfo65EB75PYBEHVpRvc4troeUHOKPJaVvBkSojGik6CyrxlgrkiOt
OvjHZK4o9Fzapg7GTXG891HzmFJv3kCymPPjtjGRsc/apMOOE8B1+1Dxh8EDRoy2
j1DVoWn+/DXElJh+Hs8ArkA93HO0U1U0sm5Wwry98//jajrgSwG3HXT3Ij5hdXZt
mtgMaqEEjVB4y3BGP/Tae7COtJx653Ive1tLikFUw51zPANNIx52jnjM2xsDEqqq
Eydnwl/9Tz4YX33FpLCVK+SFlQa96GvvsJCwVVwEjb0pvNVUFpGP7lg6FUpJE2Fe
2x6tqnlE1SOD2BZIOkAj1A2Qyx3Qk3Ju9FBLWKfDnDdTp3ud9tOb8Q9XXmK52mYJ
ORsCpBMICzGFOoqywPoZysfyO0j/Ldk/AmXjpITd+MSppa78YJH/1BmglI+2ZB/S
i7xci4GIlRCetGF6C9OHf5Da9nmbX7c2dfTy4wr9AdUGrBt6WQcSY7zEaMjCaH/f
Ocylke6EnHLZWa9pdNAnDMwD4y7Tvh8dHcuQM0PCJZayeqQatohGBmcBgHMIEHps
jNWw8hMvNJq4oB/UrS0BC/rAdo++fChM0OiyHJhzJEfQh9RfTuLj/kzndfMZnRyp
nCO+hw6dUiPo3lP57zBnlK63Hn7UnKhh6f5DeA4gMS2xVz/tDS4I/Q+rOn/ZKQQM
L+HdCWWdWAFZEJpCBpcgxUKDBMysKRC0winesrPdDk92Anvfpn0McAkAp6t6+kIw
7GK2BnOkjMyUDkwk2MEDjgF+sEZGViWYoV5xi9sC1cbgjXBKWIxvA2pK/C6h1fno
tIrJFv6qikAcleYTPqdmweHQ6EPXFj8LJCmAp0tzMC1o3Lh+oClVd8JxKng7spuK
VXpXSP28DzQ/hCzEq5C6TKHHgh/dWgs+LjAzVqj2fYBZfrz/+DJi0cQ9AcJCBkgi
uxKkoRncGkTyfAV/rUnod+PU2Tq8dG7Oy9SJ04F5VRMAwXwjxIsaCGTSdBI0DkFI
Z8SW7Q8DsUqckjA0cwV/uq34F+KRCjRF4GmAyyS7q9LHE0xqa+UfDJcJhV4wrz2p
VwM5SdBushq2gZJjPqV5OItyEGFYH7bYUF2z2qU1M4U0ke4Hx7GGmQZvYUcN59EV
URE92kZ3iCvQuX65XowlacfVKx7gq5cC1sqvkL/GKhe02YsnztZMsT6ulPX1zFaV
+Wo2CmA7IgkqQIiBD5mqPpYROkiIgWQrAyBYHcSm6unydrXFmOjimlQ/F0SK4p9K
QiLBFzg2/b1VGyCqk07zsn9US8NVVNxP9b68E55+h/F57/W544d9iNaeoW7Iozrx
LKsLf2d4wyJ2Oedr1g3dtNQMjRfuR9fZ0Vev1fm+Ccn7Gfok9nskuE3BUcdLh9Kw
RMq3/uKDDk5ph5ALFQdRRWvzli5BpNWUmO9lJ4G/lXerY8nBEgAAihEH0hW8vFhk
pUnRqhf5S8sYQJoSS774ef2YqakB7u2fsveFvg/wF6+7S7A0ub/QuyrecM/vKR8W
iz1ybfbCae7Sc6Ec2fOsRXsCC3/j0DdJB8P1aX+7H+7CJ6yebPEZkl9TA1QgqbuJ
V2ntKzxCAl+Q+aWN+vjMgJtBetlOfdnOYOnvWPncXPGogSYHxwzyHYUEgGaDoL2B
StI5bB3Ai+9UaTygxaaScMV0dVPm80KDenO1puWGdhq76KPjO0VIGZWgyo096Rha
kbmL8/eBnbOZxiUWJFcMP1iRefbE0UCj92VYvpJFbwiu12lHXw2Jdf+hU05iF9XE
/E+iMBvTzaGCPeTqc0oy5SJwjCIPYVpzi2Dp4jwYgiMoPEd8UjfiG6VytRsE4cCC
AQQNeOVdDyMCLVa/AqEdIYBIVOmDuSek0yE/GR4tO98x5hDUFtdyQEiZ7FGVD6DO
rD5okE+Yi6f9XRXVuCcD9r+j6OW2lUGpWMKAQrdUoraZ0FosM1W7WnRTmeL+/wZW
tZn/uA2bA3hmg4KnmbwQ6mqO6uoFhLNdjBof77W2KqEd6s5tvlPLPzLuo6bo20U+
eH4JhPBXmuHbkNuy5kLiagkQQoRJzldb/K+qug8zb5a0/zJlyNu84Gronuctr9FJ
joP+lgX8JyRwY+IrmgtjlNI0AMC5UKGvbh/lgCVm/PVXKnbTAZJ/tXu/BmrGM6c2
mEzKP8aZC0vurgrKu6bO51EPYXpwqymrh8kAJSGQ760ZyGQ5rMUIBhx6UeRF044y
VbJ0u1hwy+L2j14d8pXSI6dyj166gd4ofDNmnaMFsAReSZ4OPNTwLqFXK3hYLhhV
a7LmUMauvm1V7GLVTT9rJnPGe7o/sLaoAwdOHgAzNrR2ZzBNinw2OD9ICT2EYApF
qTQIufdNCXp6FRIlvtlzbmzejAp6QSxZff6Dnuq5ec01nBottLOEmrGourXp47Fa
EfudSMvu9bLbxI5GNySOyd+y3f5wK/ueB9XZzOJibCPEO34plnss4QO/UQdvo3aV
/fJswIvYw5YS0/0o9n1RE2cuSBdvVlY6RznqDOOzCnONo3ufZ7k0yCcbrWTZ4QSI
7M6UU5+Ycmg4FoMR+Vc+oDPJIDNxwM9dGjR/EPQFLyXcyNRYvbqO9C9Iilxl88cK
lBwMg5Ro2p7qy5yWeY5ipSDj4jD8753H79t+g1ieOE5HDi4f3iYQBQfy9Td4CCYs
gMNERO5g/A9hKv1Okdq6g7fRMu3DIelFPfZlcERET6GEp9DweJhKDVC+L/fYTLuW
UCYWnIt75CSUbUp6g/syAnjNU2bbhnVdZkbzU7iIULIcDLm9r6fPnCCeKoJ6svLo
/PcK92stAVThnaeIfcev6e2U9v0c8T/H/cRK2HJyu6I0IHcsOp9VPuCpo9WBvoDG
MwouGvDQogJq3EtnE1FJ7xJqZ/SYl/wY8FnkyPN+RF+0j51996i4GvGxQKHqbWGn
6U9UYyvadXrXn5k6SKFmr3R9Y0VWdGn4OidoF5yfhSx4IvozQWNWQOe1D47nidLd
IvU/LjcztpjpIsOu7P1iw6UWmnFk9cZ9yGZqZy/wXhe3EbaDmeJaFDBgNgW0v9je
LayaNqT5bocaO6W5VQpysyACMxsGs8E5DH0L5sIqCQhdu4m2TKQY4ncWj0RElqpg
B/gSV3JzbVzt/fchDw0PnXMSroTYnaj7FvqRfYs+EohaTpP0UPgTH2pDrDpUrrfg
UL4lydsY69p8sjpRb3PetBWlAeYLe9fsZdE5zg5Bn1dQ5TBZt4PrziZzlyJ3NOW2
70AC7+uD9b10qNz7gj5K85xq89GCCP2L9g7AWCRrFWKUN52qQiExNGDh3RQlni9i
7mK2K5hRkZOu2vXnJ2TcE1CNX+Cz2NlthVs2DCQvbOfiGDWag6T220gYuuHHmVWd
QBIOn89MOOWpRk7X2nYrQwkX1+aTA9sDbDuW0Smhihmy3Yq7ZPKQk2OCvAjYEF+y
lkAQFO7xg7JkxBXQYwUqjHf4pUqH4idwAwyWPKgQY4X9AAoTrhtT7VwoyziesUrN
k5KUHdxHrKVovPa4x3J0vViDiCEfTH74Zr6u+tawmZq5W54n67k88Fhw7KHg6xyW
57zfSGs8+lgnP79Uq6tCB3V3jb3B3T/dCfzaI1D3rcFxuZGCVx89DrFY0jH32WoB
QvrPj+A556vwjqZ1sqB8Ha06IGK9ZPtrqzXTRyXJM2LuhA3S2C8oHMB6LY0eBsQp
ZlNcvb0U0eX/n4lv5R3nVJav8KKLLa8xfpNgXEET2r8SvKk1zLq5Vq2d6RchP1xT
QlA7pmLi4X3p1vcfymQA3yaR7Pg8AzHHWFN2QGizLu8iFT5ySKNgWQl4hxVBxcyQ
bd7d5E8/5cdZXRcIR/Ve6cnNeaROS1waana2VPTuX1E8uvx1ky26JzTOImUXoEtj
iAB+qkNRAaP0H0vb9qQ3OwZy4waWz2HuQOxE6MvvLTi7ixIoHTvI3XKfdGeJ02E/
CqBGvvDkmk5WCYQrc9PPrHlRENDHzAkzXQ8ZPwpKCLS+Oc47kJi/g7LQbDPtpH1g
zyqVi6WjugWzRI8WyliwQhiOCsFa1fDbg5J2XSZ8BdmKGuJ9fckEXbDomqpBZBkQ
/IMzhYRVELLzjU8M/UwwppZmo+gSKaWsWoVPNCQQEm3B3W8iG3xuNpY6hVXHW1Tm
58Ilk+/IGWjcSNziUgCRPRq6tavlu/VvQtXO9xRjjdXmgd/EYFfmxj5tU7irz+bv
KX1KdsNUO3H+VR3wryNKa3Z1qVd60RFNtHy29DjkQYKT2SiJsfADdqtyHSzUf+VA
G/t9OQ64vZhswo3ornljaZ/RSUOUU8eFKZCJy+79QSnAF5ktDoKxipqyrUxXq4eH
58SFuxw+YjmP4B8j1NWCfMGO7iS/9VN8HcyZaCktBZ5xHeU5fANSHpktlNmk2gfl
IKiq+RBpCay+8dIQ7eVmRMe0Kbn9zEem/R/DiSkQZ5mUH6nQ8PyQIzv4fCWs0pMp
e2Mn7RukwK0Vc45umAoqYYamf0rYtcAskX8WKmkroBUBjHtMerTdcPKgo6l7AYDh
U4MrqbTk2oHKW23m0a0kfDuxhX5kkM7gOcofJD0xD0dvFQIgGtDUCXcnrOf4ONUX
BHbwC77UdQwbkZy4CpbSwdZ7utPG6g5bZP6042MR4neOWYkJD7qYIpcgBzrTMiSP
1iadOQR+PjQD8VJ9usANUYpKhYozAA/cbyGwkpl/G5PzSJ9GAW0yx99/tZkWHvYH
UdhDZl2ahnN9VlnMKjo5ZuBcRvKFBZAIMgJhg4Ty3J5U1Wve34+Kxf7Q++o0I5cO
E2jCLVJVOpjYeqcjLX4Ju2lKpmgxAmgL6LeTIj3afWqp/Bl4w+waJwJFxKD9Rd81
I5c3uWkEh/+NU2iG64jdrcyFkRnwcUloxat2yKgjjzaPQ1V5ryNeIsY3r7eXkSEp
//cFyTfd2oVRZXSlN0QYpQkxxrcQen+NWVTCtsJwMS06fAPiL6yvyyCmWOiVbVrU
0gn8jZSOUtoDaxvvN40gbnGB25ncEdMM8aOAFoF5MUgGfQ1biQ1dGgWBJIXVpXFG
XSZeWGBRgrt2KV7JmYhgDpHG9cRmofwvL3Xh2wxn054Mzj+nDXCoGcSx0MQwG7nn
NZQLVp/EBF4QrzMBz+Tpv2yPNMpzJnt2+cKRVHrEf2jBaEffCEzSNUnxW0Y4Lb57
okWgwNiU6yhaBKdy/3abYDt/cd6BQ98+L1ycUHxGDxmwVRhwGlMzCjrHXQeG8WJ5
Zf+MoF1JZ7KDtG+T/l9takPMo1MMZinfuToY5x/KGVKwg8ei3+qxmgG5FpMY7wug
v4LeMEMpNHX6N0NTFxUj83XbUOhoqyP8dsMFl9sVJIrga4Yuo7fxUKIJ/UztzD22
1Zhdm3VbFS1Qxd+lyP3sUvUIX6AXBxlcmW+RIrNaE/HoOYiVieEfuZ/LdFA+6HXk
ejvwdJDdTbWVIXy0nz+IqdEbanIBN9yYHEw8tN2R25cjho2dNamSX7ZLc7XUUBuK
JfLFhqW9XSBrHcIPDR77FZ3iQob8gQTBz/II1bsbYIDaE20OF4dpJsxnQFXsOK6S
mkWLBVnoZFXyMGIRfSYb+Ww5gdLmByPWx+IrdT7fKZb/VT+phcoMfQWwyBVYRa9U
td1DLWylU0QJxcD1olXzlvAet57fyJbfHb784/eM8DKbBpX3f+klTHnex9/KjuvO
GCOc7tLbgtP9z4r/AceBJY1+mJPQAcisEJmS1nVMPwOGxrEp6T2xZGOtjxIHanhs
zz48tjN6Hop51WXMiIlZ/VI8zU2BKvVNrH6wzsjzacCXY/Aq62b7HrjWrVbsUhZg
o4KJI/QAS2uXyIZ9PLeE+uueC5fiJJFIyBDYWZE8qhls72HDW7H02TMMyzF6ZnbA
59AIWW5NcvU8nUkIgB1FHdYssFUdVq7qPPocW67yj6odTPawosaoHwtgLkL521r7
NXvsOb/IhBGFDv7dYEdWsezFV0N6DgJBr0ShZ3jGO37MXxI9erzj5SiV8YaYRFAI
ASvwCeAu9anN4xY11zsgVl1NRVDWGhJiXJSxCU/7lZLtTSYvG6QmpiKj/pkMc7Mp
mNDa2Xo6z6yBDpQ01Mo13nD4IOwGYLDHYEXyWVWZE3uea0c4yNqSMeWSh6p8fwE2
dy1tlcmdSMtkmtmQsDyhJh336QibIADToC0aqC6AT3Y4XbrUek6p23qJuwvXureV
+IkPCDzIW/CMuGEh2vNfkT3Bw3vArldd4jlMyjGpNmrQxqGjTZZqAVHPRxnIoExu
tOlJsquR6DNLoDmBfQRAw5M/bqKGyfCN7KlhZPbRXeLC0xy5wCrs7MCDGfjPBAlD
K3/MWZLBCnmfAJnsRVSaFkji9IFFAm5hxvu2TZt67NbHr/As8OX9ZPdb6/WNte7l
z0YCh+ijdR9EEQIgv/E0wLqW6Lr/+TwB+u0FE4U1akEXrT/kPQy3qBVSQwEcEcru
F1AWyzxG8SV8sxaHjroMW6BZw/BHMHVjt7OXPNYw1WQUTKP3LCWSTFIkOIV75ZJc
ssUfRoBmQs1PdxK3siSDoESQpP1kXTyhLaZ4xv6QqtmZpt4pRz5vJQ8GWz53wYXg
/ltnunMM0VXNlO0gdF7VaxoiJlOfejEYouv2NFVZBVSGJn+XPSFjbsR2A/Na2wk+
evQgua+aPEj1qUaKeaHM8uDoQCUp72+1poKg44MWQhDDypQFDuyxs3XNg40KcOzV
CUGqVl0Hf0GkdSKMZ7IrKD87rpQ43JgeuWTlK51PV949hqF2/25UfOjrzQIBFbr0
RaenzfZVYmpaZ/IMOMcRxcLA8srPEm/7yVOX3Y1HxOcMKfgTNh8+hINQb8nVT5x1
obY7IWBYILH7VmNrjMXHR6qKk6rIrqZvz2lVUj5NwVilFd7SpWkoGYxhrINq3QUK
vWTROKOrcoF6Bhifsfjvqo/jmGvxI3HD8pDgvxeRpWMlDAKDGpX58gjbJSCJSAHD
2aXcE1Mjwp+1kNIg6DceKUY//R8egNWxp3o7ANp+2NObFPfkerDkcv9PHsijM82f
+pUVmMlBIXbg3nioZfNWoL4U+DdpE5ZN8nhaAcVYvjfdCvkTZfh2zIJ/RRkNg7SO
7ctwNWiAtxFMdkUVW49plyDQbptTzwb2S4KMxSR95KAKK7ewMZDZGVCUf1/AJg85
butpP1pUCub4ATTTHL2c5sqqAFriFlRHEBUyW9o8FGO1EPCabtcdYviuGRONdLk0
jQOqq87ACBUwkjfRwy1hnbT68bC4TmsvN509zZ6TzRpmOs6J1EJbnj0K0TR91ClI
3b4zZufDlbkju6Lqu28G/3Ul3bAQecJ6VHLiB+dArS3PP0oWD1gjzJ8RnZN6NV+9
aT6oxyL0BwNdX4wykP6E3msR2dByQbfAr0FPU1u7T9bhVMaFKh+Q3OuOjY+Z4kVB
7uvLbHN2JrTN4LYR0qs7qjIM3NmyY+rgeLHJ0Rc6HrS6lboRA2Uk4f/NxMp3z0sH
zvlkA3aj0KY/yMje18KoLKODEVUrwbQD7D18s+7JfG+bOVnEDTou3kQCxzoa2FeC
SiVTK48tbQFkssj/XuoC5uBwikFmrHE96JYiN7xE0th2gLFiVZtopkuuCHfUqhUx
CaOpDgLk8pJIt6q5o9ICjvugK66WBYlExHD6SQH0V/9WpYHRxX3AqCaUF9P44A1X
nrjXzzFqfVgwxLm65esVUhBXAgTjcw6Fgktb4id7anBIma+cH3WiZ0fSs+uPDuX8
+JlignoVA4QrWoUSKQuP/DjfrQMhs3GJbtVjA4ZeAI3sBCBGfrnjurSyksgroBCZ
vr9iFnO16U+KlkeAZii3Brd67h9l5m8L00QuQ7QoP/bCLhRZJcqkjcgWAEvoSFJ+
vki+tQzTxMAW2KxnbQRl1tV5gh2is8u8bedaMvMn3I+HzuWcC0sdokgxDPe7ExRO
mSQg+eHe38xbzCsYL3qImMZFBDs+BE6Zt5fD4WA0wWi1RPNxxCwUkvhz9LTt+N1S
flpTPxTX4+vt2dJZS6IEjapIycAhhJhQxLahaYePX8AMAFH4EESWR5No79S867hS
FzaW1EXSsqudYLSDtQhh0BrqFByRZCvQ651Io9AIxqFKcxyfU2IumD6aI13NiRUr
3LCdsvvO4d/y8YGDpXWjzJtUbWlOUZHcBpJwTndgiL2L/Ok1NEobm9fxW8sWWaRz
joT9iCZ6wshr1gxz+QzKWWwh8cTMOdfpbS1UNiqXjLoyVfrcaicm5wMBcWWVtw58
u/F5Lcwx9dD73+q5xAP0W8ZrnbLwtQxe8fhIxLvv0FmzTV8UXjl0TNRG8z6u0yES
sMiJI3uDlZdbevXVDr+zCtjVnaWPs9k0n9E/SANFblmHrvM7P3YLb4gPxYnI3nPv
9vJoJNzFtfYul0Zbu+FDm63e1QzYPLFRB7+Deb85ue60vOGNCHoUtRrAddSnWCbz
/AA0MG0mXC1YQuRtNq8/q9CXldG+lPRMQ63x/N8fnLAqJwWuwEMg/Jw0ws/kcn0h
59n3ESLJdGZQ0TcP0H5uEZ1D5gNaczMU8SXX5Qy8tjmSR9sTxnMUPkg9AcpKtX1H
o4X9NxJQb0z5xAqMr9hUj/4Flui0YS1M7FoMcAijp0YhguQUu9yEzHPeIKcn037j
0Iug+1pCEArkpb0Drsj24YbdQieUV76Jem0F7DQh3HLPYr/gkePqxB+tEwRCwDoi
eur6ZNNSXaEv0JShly8vOd+IG67lqv0CsRiVQljfcBTEONLvAQG/W7xahR/IkxH9
E/8uR3v0NvTYeErOl9wOJnHcDakHrCnehu5HkWPGBZE6D/W7i1ue3Kj2J2HZe1Iw
HSLa12AQcdwjU6M8p0q+O/C3r2OVL0SOyn2lumfc0Lq/b6smU+evPafDDKUOtVVk
Wmp9Rr1Gjg5yada0GmuMKZWXkK9N4Y+1WeEGokDW/s1azi7TqOXgYM32TtxJzgcd
aZTZi/vkcGdHvFgy/s20xA5lol0bhu6+kS/rY7BwFtDDnKCIIe6JJ9Yae3KfRN7N
6hCRqugdF2lLWKEfUBUlMCwfKIKszKxLB9qb9uUVj4gVhr1GpjdSmWdzOhBdsAzQ
NIF+9MGLGJABksueahdRUPDCwnUSNK/R5s7sczobn4GoBz1tCMd9V1e19lAfXMcw
+N/Fw/Aimb6gJTmT1SCaPFJ514r/34kHJUDy++H4xZhrmTBxCh0BhqAm2fEqswmM
tOMrHZz+SuHMKSt7tNALSbhpVZN4eVcDNsdB9dxkfscTDNEpRmb/aaIZPd6xgceQ
11e2B8z4nr0izh38DynaEQTHW2VpkXfhfdp105wEyJi/JKAV/cN+HQYrd6YSUakq
SPKj7Nm0mrnWMOLN4MYys1A3E91NRIcd7gL6kh1YeifgEvPGGKqYqjKLajhoSssA
bcQYD4n4EFlk/s2hDsx6mgYzDL9dSPXEnDBGvDXzua44u8jHlq6PGbOxEZ2Ph2lh
84MPHmTidr4x1Sk4ihjmEScqNhWndvKzXwM7eqoLLVDUupb6a2vvOyTEnsVPcKeq
WDvqPO7xHqWk006KHhhvyu/UbIxC8Tf3r/EMxFCurAFu/NVRtvgKB3Cw5innXfLb
dGmC3PVqEie/vdS2/+0ONVeJ0D4A8GD/HM9SNs9YBHi6RsRJl70Fi2Zumrs7SpO9
NQgywa+U88P75RpLDeCmrPUTafkI1P1EP8kp7BN7lVdB9i3a7Itkc+Vy5rYB++ul
I/y+VSJGfCcY7KndLrA83M91kcWLHfA/ocou0rG5Zj4DkGGc0lbI0vq6sRO6pK1C
Eolu6G/RFwZRDYcX23/uESakyyKzWBRCr520BM4JYKEAmOAH7Lg9WkSca0TfKqwL
UHlpYxKHIW9OYolR0aoP3a4vvpgWxyEgiLtgOyWF2AnHu7EFpFAix5QT+W9kGdme
cgTQQix5xeazHabcWta3fCV8vfzky/87KGeyIxF1gehiK+RecSkbcAhBuhMTGc8J
yIRwIeObaH+KY0bOAPZgULJFZjVFFAZlLLJdRgLf6J3nalyaIlhF5avBiCZ7Xgb2
ye4DUMsZHv4zCifrCfAm6fZM2HApKjbyfilkHOvk69mpZPeC4tiKaTJFnQ6PA4HJ
fUGJYdjqDUFU5FjRlLgoVq6K4M4pNqYIkM9s0QOOYWnUvgXZQzaemlqu3sK3td3J
f5zYejQcR6v9pllw9rchZ7gfxCCHsaiHM1MzilkVw9TrMWDSL1yCmTf5XXJQC42B
dPdl9x/08opmIYYMnEOYYT1B20HITcbep2wwuoeRTh7WDZBcjnZURGY25i7GRJR6
9+ABEqYkP0X+XqUAj/VCsSbd8QGhR3UlPAaUHW79HOlHmXY47+O0m/xzsuSWV6IU
0xQQAtfJygdNyJa5A6JgB4siJuX3kojJnUC6G7ae89ejzd9UMUVgZ7Kd2bX2Zchv
+2k1JJ0TYsEuJ2Pokq6B4ZdSFgHOTUqoD9+vrWvXLAK54KMLbHX/7FmJ3xLX4+98
oTkkYER/r1hbTvmYD7K3ofsi5UC9yAQ6u1s9JGZw/7Db0l+jKIHUwlGbdAChgYgW
6o4CCVbhJblDCxuY52T0DG8u6yA/kyQcrhWGStCdP6TTFUj481nryIXv3mhua//x
G8idTKTFyoXC25V1oq38QN/t0RoHAQD2BJ4mDEF8phLugQmP4es6xKD34gwl06xy
Fg0/ROoH8dfg+bmGqWtO91dU9150T9fMRUn6JyHeuOCy+/5I/2kLtMIHeN2j2RXq
hW67Q/TUJhwgHZ92HLOeY8e9x9SgSIR/CpIIcvC5/FRZcuO+7LLLc9d8x7wmL6q2
TlacD4f7Od/kBOUiteznFYlBopf5bRuFsc26MSxp7/8vdwHAq68K/rI0rI8Y364T
XUZ/CE8MEE90a8LZr4sOMHnOzl9r7r5B8w0qDYSHrzIVn+50YN8wCqeCJ2V8gkd1
DS+K2NjoYGrVNDJ2zVJHzHWSD5CErmzmAUGUYAdIiqaF5vUyzr9VZPQ4tRJ01wgl
Vc5IwY/KTfVFg2YP9H19il3XXkFvWQsuT4ud14h0b/lOyAXdzWwO+qmHMvxDG/2I
ZQUnGS2kxI80IDhmEuDSp9T5wjEeXQy6ztEGa+yYltMbjFogLKaBygrBocWPkXDU
BJ2guQRZWtcmFR4W7obFNTWCnEMQCQxxxzrxVnhC1dc05u2ZCJNN/ih02XLbAB5M
gIPIwARNKCREj0BbxmscCNHGX7cWDOrZZE9awyR4+tKEN7lhvO3TDVJw2444qPWq
6PGEodEyRcxz2ugn/wYg4s+MR5MY9WMdwLTBc8h9Qw++UblFP3g6PkQZvULB5shU
99UC0MKqM4RSCWfXUubR8WNdxPTfZDjb5uMOoIX3Be/q1iQJSCvH4JhEutdHFVl4
bScz0bSZQsKkoc/7pAKi10qEgTPkuvhTB+EWkMQBBiELnwzH3czIxHHFS9z2Mniw
JzzdBIuQk/8GklyAsfJA3mlMsBolnq420/q7mxGzWSNFMG+Nwrbnhd65ZaubJA6Q
M00A8S1oWKoZNHk/Eqsw36i9PC4jzGkzLMiHOq74f4nL3inF4p/7F5G42eOgy3xB
DSZ0wWRiqyVZqnJbpejTXtnF0ZaMjecOhr/EzHBZmzBrvj73gX1AYjzg5NZ3xm+z
ImcmCgm4kfbKLxLw0CLcMW4X0LsyfyhvQTBX3APuMWlqbPsGuNChdvY77qSYgEKX
8rfpxR0VoUMI0gz2Sz4myXB6Yaag8vLDYY+t5YZI8xv+ul9C4nLf+58jbVS0Dfvi
8qjfdY7fLaCr2d+mAxLkqNSpai+5PYedbp/MFwDBOXD/zXWjMiCepdGbBKcd9fub
wi/5Bvfd5wB/gjUTlBoBnB8KMXE9IqSKGhqWXdAVz7Tv59awS5NDN9/y4+vGcg1B
zz834uoAMeqdYEGuZuoSssewptbg2PWU+AIpqzBiibpHcK6DZL8keoziO/bKarlY
gue+RKzQndYmke+p3YZjV49RqDo1DZJoIJdeJ9qvTgb/254CwV5l0ms2GkY7ma2G
nh5Q+jXATNw5Jcjh3t/cykE8hNNqywBdvRoJ5Y/+w81p68004w6EUto+Pcyazmaj
hOzkYoJ3pHeXYurNlqsaVi3oXc7GWfvJlSn/9wsNtruiCDmNNTV8H5nE3auAkMwG
eiQC1tHTDZrDnGGqRWNrgvru/zNjTaaF0KZ6cuqhXxYfbetWbUc5zufmFbFxea24
RQsOzEz3Vuw/e2FNgF0jqQ7MViIwfn7RFjU98rr6/5buq/cpQCTOOeBkq/i23YvU
OkB0VSodYqaVK+SV0OCcgDLEnoQe7iaTvxxZaGX6z+vdTJSFGWX2HrrqM/9wVixu
qd2RneC80zWwH05PtpcbHSgMJs5dYtdWde0CLyJ597HY7QKSz3tL9aWbh1y7RM1s
CJKsGoIe1rLj/OLq+EdZsM9ZdC7BOuTClvAosUhAHm36Ty03zYQUS9g3LJUy/11e
Rki2xxV94DcVJqfh2XRHmrgVm8YQ4JAbC1NnWZH8KpfmSdHaltmNt2BZBeKef5zj
T3FlY5T3CH5bTSKOgRqjZxlSZ2NxvjHLszXAyj43XjsFKYAi65YZdbts3jwkUbQ9
mgVMFZwuRf1+OCFi05aDJEHYnph2aCNXPaVJxCeqiuzuzvQsMov4UOFFy3vVv9gV
R9TiXgW4xR8Coy2MW7+VyM29lrg3mFq5Ih9uU0m1cVpBQdwWnMglGkofkDT2X5MM
3dhNXDqrUQQbX/R0vJAUypvq/n+Su/Y7eeJm6qviOPFKuUG3/nUMFrqvg9s+mOwo
nhKJN5mhJltnFSgi9mm7Laje86XXxJ5c6r+V7a9sgtIxByltcVQEmwWv9kSRHiEX
Gvjn0Z3aOb9/4Ui0UqOw52EV7ZVE7YfrmM0uPVtbk977c7I5mXKNNJNGjL3JJVk1
fyT9ZfYzCyCUcRIh1sfvzuGBBoUoJiupkrniQ85kBwAncZePGnt/P9zWjZbjRe0x
edwnOMiNjBgQUwAuihQNn84GkVtxEpR52S/l15gnaFpScwhUpl9QFkXSvtZ0om59
Gk8Rvm/a0ZB1JStns5XmqSnN5Iz4vT29KVsrSwTC0aPJjoVB/2U+aM7cCh8IITko
jXnMSnvFGt0cr42WNnvTJ6e+CERgbvNrbx2xNp45XAP7PBSNSn9VxrxuyhaYCPbb
AjH7jJsJiG/uxszxTS4q/EvQGuVkasVL9SsD32G7YZ0r1ERK//0uxcjbtA9N5Wjd
13HiOipaHe4eWehvLPniOwf/MbNd5yvQoqTYPHIykyLMEtfYrbsdv+21x7/6IGw5
lp6cb56gy3lRVcQ4AFqcnHu0UsrrEH4TJ60mhpzzBtphlctqjSDrpbFcAg2mtVUC
uoa66uKpkBzPdACdl8IDtUuMa8XOSk9zpqBQJv2A8ttvpuhzsR8hwwI1SKLuCT1d
oD88yFFBuwtKcqLlt/fkmH9XopNUcmBXVMXru3r6866g+itHMMkOfszfVo9aGrg1
vmPs1mTADQcbitKe4+ZKflxFKT62CZgESmWoEMXTgSgk77gZ5ypFqBgvN0C4STSE
gjBbZdIpx2VfzKK2rrhTGgVoP3slzVp4mltyIfWXcYkBFiPTjQUSvHoKHSNSWYz2
ZEjN16FZYsY3DM8KlQFk5CQsDzXLiQMNDZ4bjWwco7/uc+kfJzbOfl079lJ6vFRp
uIwgq8yjEawuhT6OZPamXPljLIZR9eB8bXLKrJVN7LL4gKMtCWfzHRDSxEZyMEdw
1lV7hLYqgihgnA8RsHpVxNJOAUnDyPj4eI2p7T0Hweg1yP4nIe2iDWWKE3cTtWMo
B3U8eEfpXdTvP++G2nqFZ790S8QzNWSF5j7FmqeOqk3jdHOJnKM4OWKHio2XvQAe
WCCam3I+UBmIdkCStlJCdWiU+WMcjJfUMyfxb7XIznxZrpADryNj6ktd/btueBBL
rEWPWCi5mW7mpFXjGGBrjOWk6XuBP1UkJBqCKAwK0GaKKjbNqSLGREICUydKNVna
xGjIUD6juq8OB5QU8s/KVOqiuvutZSjg00ArtLqIxYXyS3zBR9a6Ub2sBsVG+GEB
50sHVzJpdfxhojDQM1mf950lLVOydUycZyWDQV0hYN7UKFctegTYATDo8lzQibHJ
zjlGklRrtEbvgKSsJu6nfDG9JZ/vQyMUwtzE4+kkC62uTmPa7Uzte5MW63ziAN/s
sys/PkOOkEVQJG/v6ZbSWKeF/4Fsirqt0PoQMAt4tdW9stcJZXqLrQ9VGaCURC+2
EFFkpNgPR+i8ckCXCOsASrRrJ508vLJWQHmLyQAfIgemDmcSWzZC7yUzyZlIX5nU
RcXiwJ8mJ76xjuayToSSW9tTs/V9IdpXroSbYfAoG/uGhf3r2sD3nlFg4VJTcguR
uDSDX1OvpuHIt62ZAbupWR8TzTl0ytFDjTnB6CdRrzg4vgKknQ0E4MYfxA+KoxlE
ezp1fXIHI8pTNU9IBWTGrOzsVgiagJYroocwM1anK3x2YThB3wcZ2i9Y6yED+MZt
hmYNIC2hTarVU1k897pWs0bF1RJWTgeN3IoVlTXefBhL/rf3Y5dbsEByl8z+mD8b
1KEL0ZXDJQZx9pktrAY7E2fxQkcnooWcAxCpihjBjbp9c1y9uFu7UO23Fp90RoUD
SCWBm7S9UTzuEtj6eEW9gMkzWqJozIjEU6mWEDVev4f+kGL8lHQBqcE5vH3ZEG+O
7e1P+lYHPRQNbTfMJlUpCULDr78iYTbi+r/fEIDEvpIz6Swf562ocVSaMO0hr83s
d5dORXKiSViqYUvamz99mA4gCfhmlB12LiK4ZaNv3hHtK5OEd8eeWNCZpYP+Y9xT
HkHsJSFoaPAgae8Dkas3KCxW602pDydu0E2s/RGW8Eb8zSWufl/A/x4CurmJsDUU
5MCVxAjzqXSdTOQXCb0hzj/Ur4lnmVFjXMy+L/aLP6OujB/hhf//gduh9pf2X2Jq
M+rHaU4l0rcc85DKqZx33nj8jmBhi82PnHb86PEkyUs/pydHvvZNx4MqqCM+qJdX
kMZ2HS4SBgcd0oCiS7nqEq2Y5gegxZwlzltrZra/lpZvuTPLjmJtkUxBW1UBbyI8
Oy1MvJazc0Ajs1OWrjpvZFiUnkspy/no6FCDKmxIFLjZL/pQf1QwYtX7u1+sofP+
YC9rClLHIfSYedEtxCaJimmebErXNKSguhXooiFf9N6UC+OhBX33uKfbG5lMOD4P
O3P0WpbVbF+kPAQj6WdPyfPCYVtj9EcvhmgsUvFbLdyS4eumiI5ef4Mz+BChxlm6
+MDJWN9xSRmClZTus8ORUzy/BK4CR9ZZvcs8aPbZiUSBUggRTPCVEVrgAStp2o6S
/RliPd6/2tpoqeWg/MOKjCUcH9IWWGBLYRVgPiDOL77Sj8OZuwfLoFp3zG0hEH3M
fsgJKfoluhYYaivvpyk6ArhiNXURacjB5vUl1604aTZXliCG2EGfTaEoB8T07wHu
9Txmn85kdUI4V3SoF6McFjBOuypr2bDZ2hPVEg5mWND44NQvn7RLM7Ld4dkpVatI
W3jtCHF5/LmPHbbuwbVqKnGUixVs2xUHPn2yqTkFDplrYsv3VqrJR0daQNq7xQXs
JkI1CilRmrV0lucazT4nJH2fcHHTa+mUXzzGwyF7QE0esguf7mzWxLMZaMT+x6Wj
v0/sUHZ9H4k93qURgdtlGa9Pbmvj+RvEkPcMSrzmKhMUGCB2CmtWrmdMD9GXZrYD
uafoSTPgoO4f/KcjJZmPQ82ovKuWUzyDYCJ/lMtU5hcObI83iQgqwnZ9nH+G1Jl2
ohZwM+3LVql13ifyAAz0s08e3L1WPV2VJC8f8D8JuAZT824lIivnqTiQplGXt/Z5
06+YAQCtxMamxkXgqWqUdluWGpJt3d5lxk/TKtM1OeBgj/+/E9Oyzk10S5YIfM6M
Ykyo44rDDOHyyJ0YJAN4XzMMOLubccjdGkUrgdieYoJkBY4emz1G/xL8c+PWsrSj
ty+ChaBFoeFTdZYJsd5kK4e4mWFZmdkV4XiQOM5l+GhcUA71071VvLXgOT3PsCYY
VJL/QTvL0bKzHklfZXznF38TvOZ/TR173l+xOAVNieeiIlbRerFEWz2nAPaTCFxA
ujuPAbWjprNRJS6EwxSWGRMnk6B+UcPF60AwtVdaED4nTMIoRcylncmmW9fuCeUU
S0Q3nUTVuETbSsijcGTb34cMEtFnogmFsg+dWnwet1a4xk5paRiptpG+sQqpyX6e
jGuHJywrKd2HwcEKBlI9E54xBYbSm3AJ9IfZ55PEZP3pHoG0mimEEn7CfbOtllnN
8E8pwB7RybwlApGCRiyrwH/uIGeXcN1mq09yoMCVM7hjyxOtgsdTCpyEj1/zjYpg
Ja6JMwnI5FpUhwhfBa9zcLv7biy86vQQjz9BfgNzP7XX9wMdC1sw0zg2tBk96Tjz
7038n4CymCL2nvraXH7f1kYB+S6vkMkSxBJSIT+lQA2m0cwpiRckUvU2h8wO8rUN
NRXXHOv+CmJuHfURQFfCQx1K+iqlcgSeuVGGr5mF1yhedG8A9XRLnnJFf8JMtOLT
nvD9fq4pKHuE24wACeAaI47qbToK909A8/WakVrWLg/w9Rjfev4xQLuZhqPDAkW0
9hlWAHQS5ng5zpYgofXrcrgqdz93dTESrnEAjaPfCAA+9X1SCRd4tzliSKzQF9ci
+w7v0dpibvP3UQqZfa3b0GSCKXR2J4fR5dKXID+mGz9zare+g4q6xp4Jkeqi88Ck
S2s2vpiYXC/YCMhrQsfMFLoXUMALZQ0OXpZUHg7N8RBzwNXM5wX8r6+1iQoasmZB
FF8vlafSIQrtnKyox/PyyOLTjRWkmaoLCOjqMNe0cJkDlk802wtcUnhQ0i3v8XBs
dNV+yQjA48Gha8WVFdH2JlsIGAMqOwBR8saFnwPUiH/6GFitEVlBUcUqKGsD4SrC
1rlH2Q9NYCZLA3E8GofzBfcWv8ma0r4Yst0pJ2N8XtPPIWmESxrw6OQmgNj9wxwl
BeAqQi4th4InwqxhbyTZ2DXInHmkGZga1VehxokpGpOLvVxR1skmjM/hq2M3sQrH
mb0WU/qrYcMhg9Jt/Zbtmm6orkzQvXRzq6aZsiVveUnls6qcu/VtFPhZ/6/2/igy
HZVjmyki/IDLI4DJYZfPlXFYLMf+h6lNDtD/2dIT+Dym4O2vp6BJUKUJR5RTrDTK
SfAlgTvTiWIL63iLhRVhDrm5F1SagTFSE0eSS4IyIAifwESdx7cDUo4ir/1PIg3C
56maa52SX/lElo96BQ3HbmeDpPdKeYz08px7MaehZjFTHG2M0l5s3DQfyGuk+1B6
5Sdni2D3cPO2z5CWGuqJAP1QWYjCeIMKIkrqrL8V62lx/u1WGNli5m668haLukjK
7+gbVnryIaydHawmuaSPhNklYQm2eFHsXjSqxZ/xThNGV7wqVHsZAsjkrVujMH2b
A8kirji3QeaeB7HzuB/2tvVAqAi0RVKzUlWsERKYEWEY310JR3sQXZUG6m8VGBe5
lyBDsXAPzSQ4rHEPNFCZr5FqqPiz+FsuRPpNpY/RlcV1JZCExR6lL15vFE8Rjvvu
UH1YZR9c45t+1jJ9/o34Hx4ckO4P0Pr+yqrplFCZMmYYVeh/SsKIVOOfkoAVZE8Z
ASzV31WJajTi+3KY7ORxEGgro9fD1ylmTIRWWN/VqFuLRsyLJUmxgoL6tVA88x09
+54KJY+iFJM3dMuH9ahob7rrGEw5RFqYCiSQ3ayM4/BLYReiR4NI+vLyWw1CNAZF
LFOfzFAUUeMMtjnxWkV9X1UcKIdIko66dPS//nsplwDakRHTWUNpJojMNtyxik3Q
8FaeoHONq8LjrGfkwxoOvV4j0ArBPCAQzmefdMj/WFqpRcLXR7DgzNAPqmHD/NMg
LuW0iwgFD8JDdVYxZAUpF+tff2hSRZAmglua660Vkb1hbd/KrgZlR3rDz+vmWS8R
3RjRc1yI4kieTUogfuzoPxQo7hdem3Y4dE68dhlcKAzL512yMozUy/sJ0NWltMCL
bnLNdZVNUB7fshcdNQOCM43C+QezUFUpL4q1yKvlCU88H3GnzpN3yFLour5g9uA+
MNctDOPRxQM2V9N5yqFIooXLt3lzsXmS63AIxodw6QciFcc7FjZ4lGM/jmZqFE3z
jthC+WqTL8GLHaQOGvwbCVwJmHtrGnhCKzImWjd6JPLQ41Jt9WZpnvOUZRjAYlaL
jB7ZaAzLZnMs/HqHlqRSxPqW/JKH8OUtHuLxyONRkVLFfaV/oBVJbRDUh/iBBaBY
oLxJT3mgU+0HMXSU1GdvXOzUt8kpWRkOGphsC4qmFHdYq7IVBI9Cdcsn3MAEpiOS
jPXvmKK2wO2DQc6mqZc3WISyKtlRq8RX7gpFye0TG5lEKOOQRTvNpAde61kJNi1Q
lZ3KE/RblCoyxfASVXSEyjr1ep3yEbwb6XvK1cEWPJ30SgdFafnpysdNNhbAsmMz
8kHjf3zzO0SNgQgDd2z+vjxtUYBfHVt9YCnZ9mUpx7vSpH/5hq2nNaO+cXpQPECH
1UvjasAdJAyXthk6P6XvjdbsU5DFW24A46mALfmEThgTGQjytGaDikA8EybaWBbC
sDgMbmdCj9M9hmthSso1Eq05a1Mdkr2NzGZcEhPMgTgHDMSucqH0q7qlKCOaLtxV
azqGtpZpcMV6hS5clgc3LdlXJShmZ6KY6PWtlDJW+HAaH0ed25WOqHZ9Rh9r+0Ut
OTWvrTGRxB01+C1baZBDhnK/KoX74dWoLem3FMweGsEhJwSPpgGNlkmUEIzRgrYI
oiCXJ8mmDeZ5F4Pc3maVBqNwIRxBuwQeoriUlfAz0dwJMxiLfCJKaJri+GY7jiuD
Lwg45N71WrO2m7lL6cqbBcRKcBNbm7L2JPXyR6n6+PtKj4K5S1ep24/3hMtm43UP
0jcFBnXIdGDTXqRimHbZ0p6v2bUvZaVuifePDOAe1LAfTMxM4UfiOONANKijrsnP
PMepknpJT3ov4i676r74KRTwmB+5+lF7quBJxreuXdXQ1s3NB2Ndop/tyrlMOuHX
RPigYuWDEia5neNm/duq0cAbDdmPhURHW0M+0ElfyaVAIj8+HqUecUdu7nXqApg1
sIORcPmKICuZUdjbFw1ULe0fotVAt12v+mo5NBPIDeUKm4BiLR05IGMfAfNY4MMw
uXaBWLxPeJhpoMmt6NQOKmhTYVYHJAm988uX5bDjgiBqnN6sX66WSipktuPFDVGx
40oTbTFRqSH/g3l9ezy+YQidJkO40KyBlGy9gxOYOEVwyZY9qoIvc1rcF+m0SuSe
iL38AprnxOIy3+1kPX3s06eMm+eR2U0MJ2t9L9fwd75gXz1nh8eGvrVL8SeLyZot
qyLeoSCDHyX01J6kvddI3JNYc/I1veZHNlzZltuAcDXIC/KXvNhevQMl5FrLnmJv
PHT5vuq7gHGlTMbqHQ2mAWNHJ2fS6MAAv5uEy1yNsB5LGEqzvM6f2JDyq5wnes5o
3uZvmYlUcwnXwFNDztteox9ASU1wLehHkWl/UziEjzxGtJbz9DFcDDXQFAR+CVjE
WHC1oHFZ5xPoPyoVwsbDwIxEcgb38EVqCHiR4ieMrfZOY6/oz5eNtNiQF8fs2f8R
OntxVqgZmJmkAsDoheTmzLwTiOsusQzysphTviBN1FYHtKYlXdcITXbqpBVZsTZd
HY9NEj18rpC4m2aXqnJUC644zm04S9krdVaREEWym1mX3+XJDVEIti8nONldh38B
QEWiVOAUVT7FolhxBDl0Zcrd2M6YRnV/fA3HqcB3QotM33JeEw1OqsfMfpLd6K/h
+GvDrmPCUdtNoU6OOiZMe6ohzJI88pW4zQtY0cpJ+8JLYIOo5ddqXJAneW7Gc85h
xIYZg3XgXADAZSVCgFyRKA+YEo47yfXkyzjRlAGl8I5ltCetWwSVLWjTydmrTsaQ
p+zymdrGI9tJQdT2RlYunxovbIG0UCFfj28NrFaooMY8i/tG65gxBIDKJdfYtiRS
G+LANSdmpqyTQeLkvGjxVnAWKgS+xe3AqaAydria/8faunGnKg5rGiW3lkK+CIVi
tSPNaVTzQhufjeTznM8b9Upkl3wCsThMw/AsPQJTxELghK3a46Ukm3HT9xM4Ozhj
abkNRV3NG7YLVXm6Ml2vX45ioaCGjRFI9tjCYuAy8TpCfe4P2SivMce/4wfaCgXj
mrhIameCIdmP+ryCy1P+Uo4tarVPBl1npl3WEIK2yRbryHUFmx1ZSVBOpl4g+VX4
wKggRDU0gLuwd2RE7DZXhn+HTamT2FP+kaeAynfSE5azSkv9fKJ9jPRGNbEpNL8U
SqAnhDthelfIb1lu6ZYzYKuVbITLafWsEgjwZPDOMo9QrXrt8gWZMISbV2qqMrMW
3AS6EhaXl+I+oHN6l6QowZij/3c2K3cItMbgW9EGYWLtmOU93hcX6XGaSwNLUisY
IkLBSe7r3ZoyBDWwMRgu9vj8mXadfCkjfhYgVazNs6hAAQe2NKVQjnhWFkULBPp0
aY1pcUH0ZyJl+gLkWruPu3ftLCbv6oxQjiMWLlgKQ/8OB3OLBiqq+1Lxy/6bneJ6
2KpvfCcuuIsYbD2iFdZTaGGUYsg0+OwGg+YhpD4KNN1hZzkXix0G20g1+JUSOtVS
uGi4Ka9TDf6QPPnNQrRb70pu1xII5W71LzCoO9cuV5cf36tlxwlrE1P9quBjuVoz
c/nR2ZCkLgnraKFU3gdlVDlH0rY+aU4ekr7ISdu0MLkrIGyfd+H+qT3GkfjjU1Un
QNsyHYAzahleiknggTB/DwCsGiCerebElifoqvPpTaLmWC7+Qhl+94PIkfzRUygi
5Ii+5qp8HC1o7YGuiTGHddwCNgm9x2p/ubmCioj0uPCSkuC4K9r5XFfqb08d/fY2
zqxyWPqfyPHGLSzBKW+qPDcZeNZv2YMJuPvcWLw0YlHBudpk/Zmuw5MywQt3EH5G
6AuAjp7rqemC1K1TfFnBA7XBD0YTuNYJ87KND5vrQQlBj/6AgR1UW7qJmFkUOgpo
bA9RYdMfzGT2y9seh/SVen6Mt1fGk67y4egPPWaj++N36pzdJVYp7nCs8txgQyz3
lPRvLU2DPmjD7fdzyhqA+N5iZ3HqxDWHEGT9AE8T+LvvFKeRaGh2iYFqrRPv41pM
6JNNAiwTnshVaOnsJTrgfFdVpPBSt2wh3F1hKmRMnuAxAWxKCl1HSa6wvYFiPEyk
ypPG82WLPxWlqtrz8mzP9XMw3+f1JFHtQnwDtVjTFrFRi6NUKMwBorZYhUAvv7dm
z0pWL200Urnpn5v91e7H4ADTvyotUOz/7HRTEXMyjwc0Iz6nF2qfd5h/AoeENq5e
Cz0MiIb4ZfteV3GZfigDHsTxMZ4GkYVVt2gGEUrlz9kwJ+oiDSCMs9ROCXHYoer9
kbsAS4VkUswc/3N/fviYIwKDuahXBpXxbABHEhTg37ePq39WmvzFmear4fx6DU32
W0qdVJmvAxGGkvBSH+GKxUKL9IRBI2gMeRneSu2ozh1zQjUKiXh/wZMdfc8YH/fR
1GIsQ9PvpqAnyXak0r6Fl0xj1ck+e1Uu3vjf/A5FWuB/7jqljF1f5hSR1R9MInU0
mYCWuGhKJO/HiLqzUNJzav8VaGi3nUKslIqMMuiZn1n4GnHA4fd2oxjdh5yYnAH7
nZ/sXtJ8WXULSwTXgHxsGvb5UvYy+Y69MdCB3nc8x7ja/phNorcG8yfbkAbhSdM0
mZYdZqEFlUuyroO/3A0y6FuUnz+nx/o4AonrZWDFmyEeaC8I1ciXGwdI00o1wbQl
WXOUrOCZ+PoVVahRNG9Hw+ubOke+StOtWR2Gg4bJR9PexfHsZ9dXxEkvFNuLvQ4O
tykgqrkEzBlH+qrhOKXBmntnZopGO/rtXlCcj1vht05bLyJTlnrKJvOB3Z/z/5q/
kIQ1knyePRKUXX2Hynd2xGktt0nkkvc4EN97btzgsFnT5VtovGa+F7aryEgDl3S+
spnxNFvKnU4r+WVfoKp9SpO/A5cJRjY8FiDu+IwbNTnzh5sV6EsLVYuoEzEckUQ4
JA6FfT0P5Bp7lOyqIKes9Jr4clHEZxXCmCpcKdvK3dR2XMBdLcBcrPKAgrjj4F0x
rQCro8Ch2GOnSKNxE4nNk1VZs7NqMaQujc3KAJiQAJlhRtbVM53LMuD46oLjqWLC
lSsINBoeHidda02zjMqQF8OzoTiYR7bQQyZezIGauCi9rWwvZRgL152AyJu3IXlP
JxOOEZjhPxgYoBaVP+cfnb5/qfQSNXyE8sPFUfyq3hekVmRJjlGXB30Kezzqy1QB
plIB//yncJ3iPkdRl6v7dmUb1kliCC6QhR4jv4QraYl6Z7ro3irI9xnyn+7lS8Z1
rtp5aETtBbXE/Z5sh443271nQ/nIgPAt18o7+lXsBrpNDtqHVyGs6cF3FO0tX8Vn
rK/Zl0P/cQ89QuAO1tUEVANEEsZHOQ6JwMAhKrZ7O403PoWjhlTR9FHHAqhAVH+Y
GkwrctkIQBU40HZyeATmm130zaAFnQY49J/LuDt7JewkDu3L78AWQA5TroOhAcdz
hdI30l/upLTNGZKDBV+PHdL8BjC7hPEbemwFLUEgbs6trSvXNPJn/tpqsSMkji7T
E0jqXqfClTe5OcaFcLdvVwbWvz0ZOQSq9UQckgA1stJpogujh4QcpN6aDNlYUdmA
oXOtwq0V+4JHeSLtXxRcMek784+kEQT6okHYD1lMDhWm18qwGRkD5SyAl4/00joV
aGhYnIuSaiWRWJpgdY3BTJHnfjTbGZqp2j7D/fugMuorrOMQ/3WP/T7WxxsMugWE
bEm/f9Ao3nIlAjCM6TY8W54CFK0Og2KMBhH6CpaQ/F+tCXf70uGw7BZBndYIiLmv
wto4g2uioyKIIFZEtG3AUvu9eqnsWAXmPJm8x32zrx9eJYvi+W5x+dpgQFfyvlK9
uLt/KHShS/cCtwDy7hIGWZadvTJ1Y2rTmLy9AJqcv3MP47ucjelq9YTYhElsLtGy
NqD7jVVY6t/DLojawdZMigDpQdBovnZ9dOK4PB5u+ZS2EGKfjf7W69RKBKMPXv7S
QbQTZbRznhuLrplmqAQxKlqlONGkROsgDAtU1OY1mCx1ZM+zp+GGekLMM6wgnoww
R7R3CbXberLOa0VSV2PAOHS8b9od8eNQiCZ3LWm3iu8sUumzlAxVQo0gr0PQA76Z
POahPsWIiBzrojYjLBACVNSwBfFJrEErfFnAd4vcKtaNNIDBecvfZ8j/WNgRMEB1
R4w4jjiLNgv/C3ExpLxdP+eArW97wsJMHUbId05KvmvNfb7CJMcIwLRVJSXFOiKX
ZIO5+IPsoycTzAh4lgE3eVglzFxak9QQwEfC8HVshcWu2KAzqYQQ+aQHiQefiHh9
4K2gLWyCnAhrLOMdmYPVfG7/bc5qTa+T7gsd6JCadsXhShM3UC5G0ipJRrwzIOY/
mouCgvftHfoxsKfo/CjAKBhkd7V7OE5bREiLSxOK2qIKaxD2UhQ4sMmdIVLPg5EN
gDQmZbIIYw2PPipM4aBAJ/SxQFyxL5cRh7CN/WJSGSwKXzPSGTTtR5+5hdS888UO
dSSAnE7lI+GP9VEgifgubwWHlU7ztosqNGgKiEuAE++RsT/HDMVWikcuzY6Y9nHr
J5iRe3SxMq+L+zmcpv3TZi+OFt/iRfQcsyaiprcsQ4aYDLd7UP1tsA2U70TjyOKy
fzl4NQ87Pod1sUpxdY77sQ64XprXk9wvPMIMaWLJJs2F4qiwJRolZRwzUh6ksS7m
gq6IKLzxsatcbnvsMmQwFnD/ia10ddDquwuQzDVEFT2cAXSuZ+hf5IJSQBZFd3cf
R0+K7w4RSU1077xcW0eMjIKSOjFGVgcxrRQjf/jWtuZliiE8biytFo6g8SToKnr3
bCvaePkbH4RuUbzmLfy5sfatrDkqpZR27KIcg9CSgSoglRJ2Cl0hUSUIVa0iuxJB
S4dR3vds2GprMUsJ+IhD/K6pY0wqmtmM6LJdXlBMqXTaFwWXSvjuqB3Vnpi4iSYf
h1EcYYxUP4Cnf7DwCex5wSI/5dIJD5FQi3p0RREw3OUmn1jODKnOQhtU8ufB8UZJ
FslvOX6nLanOjx0NgW1eFgzQBwY9z+UCFkRAnuvlBGLrzMzO0eDYHBk+4/qGdIN6
BdH/wGP5ISc4OngHr9QxMC451o2o/PiVWECyfbdPTsJODk4WTggshqwmu5KWn0Tg
o2vyuXu5qT6fN8Mq0Yt1fk4H8beD+8xg2CXUdzS3ggYBlBDSWR5Nw7PKk3HF7bTv
cmxTzmraOxMkmubTH511klLuj3K4TyS8KRkz/QZbycmuseBkMRkKZWU2lhw9qga5
oj4QwaIINztca1o+9+kDT7qojhu0PuIP1ggz2DUUFJUB6yAUgu5MbPQQbDDns7Na
0wf/0el3LhGP/3GTAt9TveUzLsKe/X1LJrLLfq6En+OC/mrZwp2bkCpY5OBSuOmN
KsZ4GTByxatbvoY+z0q7Ok6iE2JsAFIOzy6Aex0NLeEHCl1dQUp2wkjiwu1AQ8W/
zhWElnMve/MGjSgu4fjFtSofHG118+2Vd6+iGX/n63pzdvhHET2Lmg/ENPiYt94X
gtCwSZK9Pxdvko2RBeIolo3QWjscnLz6CKTJFMXK7MdzNByqg+A48lrIrypv9Qqj
3mN+VzLnon5wTS+HUGK5GpWgCQg7G8DjEAhJxih0+48ULCJ/Z9505BkpO6IlCuL3
ukS2qyN1MJHJ1fBYnpwcdtnK5q9dz8cBK4vv2xZGTRZiwo9XUU7J0QI5OV82IxeN
oxcai8ygViPD8GvPdpRBbNgS3I8Rps/wftYkxmBpVtuIqbKqG5lYSVz4RHwwG0AA
TULF49slQTKlmnFowduyAWtH3QPucmJfx3lURNrKT6mgXFiPiNnkJXHpagl8VkGg
3dkLmE82en5ZXrgM67+3OhX7+XYgySIQIi2Sp8DLZ77aZw+gNwj7GtO2OMsD7DSM
gKf9Colaq71tBkMsIYy5z2jZ8dJqRAX+XJZwPYqRRDVGrLCcVN05bZQ+uzBxA+v0
QbSCJH/YzWYyXxYo5789/udmH+3RO+jfTFACK9jUXajaww5XHH8ijdqFx0StxsWV
rJgWe3fJ29qZSLCyqFKX/6DkIsEBeK7zeDrswOuBMl8TD8kOhHWfHMZIrEMM4fZo
6/xSbcj5neKL3qNDVMAr80covNsXGbBO+AhaEUuq5b7Pa5e3+ay6am4KKKSwFrAx
6PYpMJHNuLvgpTT0rgbDuHL8FGbVGldcyyy+3R/6OYpv+NHL62xFTgGEfNhPigjr
npq0qioWKLagMEd5ZJyCtzn63bpOxwXFFhOlxhPhhUIYLYhVTgO2z8VQ7w0kHeuV
ntLC7j/oXkgttikUIsEilm4rmgfWt739xLJQ+kSKcfioq+/iL7OEmr7xAPSYcPEp
tw9OwY1m3LWcJxuvttNbkvGlxPIIiIxrTgOjhc5tN4KaZd6Liu+1Yn8m684IZ2so
dH5ERxTAXpQSrNED0T8RnkiJOMuAsV5cIUgKuFDsc0P/6ItPZwcdsgy9GcyL1uWu
fAEvHPRUyY2F7U4xEXcs4NJST+2WoUIr0ub2PVAakgngiOFuOwRzXOj+2oG6xXA5
BeLHWhuVsRpfg0AcaHVFPwZaa9TZlLLuBXcRD0Bgc+FfR5kQduocchQ9QZ6RAxKS
BKb4ypTD/x1QZJ38WuXWFxbI7q92BVMIvnHv3ZEjJEmtUSo0oZrJyHsAQ5B0X1mb
4P3HkgzZV3Lytx+P/CXWuVhXGAvu5el1+c6tTEYsAZtsS27zUdJXb38yCMKsSCZi
0ZXzpRFxrLrEj0XPXLdu+9Ef9NiB4VV5tRX4A/e2z6wLFH8ppkpHgfm5Vwmo9GgF
FDFMtlIOWpy5HdE88VLnpb1Dsb0Ihmy4vY/DON1zj6enDJNTWGJssjUdm2XL5P15
pW3v5gHJuHPI1Sc0WUyBDq1swjE1ZtdxwT1wdGBMbMjqkJGMGV5IOrx47rJLhfoH
6eEtNdpbGx80nlNMMdT6tNpayAX1T2H6FXlkIB/eRdbnm2awpX0UZXLYIuVWHgNJ
sJP2XEJVw38rTwqtff62/d8i1f2gPSKzDi8yxrOAG/nuyO291SV6/iPkdeRHPlMm
9DfM1jjdwlsV+/zDKqkrmS96QkweHzC6TRw8VInLNoJ/xraZNVd/vb4A3nF7hd30
M6gvJbO0bESR8HEpQnyB9Wh9zMuepLB4lCIVJzemRbPU9g4+uBRu8izLQ8YbQS+M
Uh6eOvgQ6tvRDIg/FneMxnwU59IG/nGNViL9Pr4IQc1fKaTGaEV0CyJR4kGyV/T9
0iVnZq7yWrkuzEHwK4w0GtsKNkc/5U/XlTD4pt7KMdDf7r0xMckvB8LkY9Y+KZ8y
pBvobeY1r+UaMmTjOMn/hgc+mEEE4azwpeyvw9OROD5mol8TOekDtk00umTZl9AK
g41+/UrYw/SWlIbu04App9+fPJwL/krgktHfpeCUcZqKWKiMk7sy/FcKv25qkrKE
P6xRGAyC0UYT6+ZTrNlyqYazqjnJtGNHg5FM3exy5IOqJLZqbnc6xawMZ+/lHUbk
tMSas5DEDwL/S9P/Qiyzff475cpMlnpYSNNZzAjnODqRUwUWd+NSq1VsXw2hulDW
myYTEFb8iX8bODIp+5xI0E3ZKkQrr3ePwxHC8i0U20pkI1Lxcz69ArA9wWifIK2a
YI3xngHS3WFlepmVDpDAYecskBp2JcTz0bN2/njA+Jqv4kkkWykhsCBJubDKCaAA
LWxtkjcfF7q97gE9J/Xa/YQkU9rNcgRtawge834pr69PPPcsYJBf12jn29tgMHEb
DtVIwk0qTWpwGaTlAljrJ9UMlU2gPW/bn26npTbXV/U+CX73qV7FmCCVwqFI4uu0
eQPYNqZdjSP4AWRbeBKKEOTMnXwzjFQffcCb5HcVbIhtknvU0i33kVMlFko2ZKRu
XDecXLcQuR6zsay8LDCp3KfYduyhnISbbqEA7rSSACgydDpPX/sgUy06onkBe/Up
4IuK1PdjgzPcfKOsBOJ9Hp1nX/nUcjQEzHvVib2vKD/x5mrBX3rXaZNgT0+46T5h
wjxBMkxHL7WWAuIqoz8Sbr4y7ilwxJrPgw66xkCWCip82iYwgnAIB181uGuzyUws
rhOjycIDJ3XjDPAgZ+v5xT2ea0Va4Y35lHY39Y8KA0HzBilMxWOAKMLiIlt6bghi
DMJLu9yItcnrcJehuLM+yaDuxbsy1xbZfNtsZaJtOY5VuYY83XFRMznYMDKVs6I+
81oRCwd/YMaB/dk6kZ1NPlaNpnGvt9Hx7fZR2nTHF1pBDs5tLEuKXIymfaVwFJeo
eE6tWsF3Thh5F1FgRS0rnkfEMUPkK5T1qehmB4vpnooRw5Kd3zirXG0niC+Vjzlo
a58AB1iasnOFNbIjdYdwTH3oucCkpQ+YD6r9KF2VveOOW1p9ZJ3FWw78aSZd1DjG
3eH1MbCJNs5LN5T8H+Ne2QlZGVPS+O3YzKeqaHMzKRp1SzoUNed5S709/5nGbQaG
wlRRdb8u6Rs8wK9DPboIeRD01WjUjEWiDHz+RHj0CaIlDVasznogCAgb1c7BolQB
AS3wN+T7I8GrkxIMBOuPGQHRenYW/uM3NiseD23AZCNNdLp9V06f1kf5zTUwwtQs
jcdVCZ2plbSf6B2FnLQHDFiteZrVGGWfT6EdHKCDaO2sJeuWQ/D8qjs6GLh+01UA
GFSBKv1TP1bHg4bilOEdTFXYM1M3R8f7RlYbAtrpYjDeW41ScVJJJvNM5Sc0kAqQ
siUPfCFbAMVt6pdqwcLQ8OJFyTwKlwYyHOYQbS3b0LjwaVGHGGyvUQGSclaC3hRJ
arew/heROAdmgHU+T8bLrymEu6SdZMAADyf4YvWXN15e+bMIAIkDhhC+Upnh5QfU
s15Ocd1NCQJBUga49XDy4o6WwB6DleisKCtILyhQVyH3n25/HNIz5id39lBpDSKy
QVs5J/uY1dCSj4PpVrkBzWlO/CYtpdXCG1uBnGDLwvREQ0gM1kivaGYaHgnFcTL3
HHXrQSdBIXRUJqZOdkMOt6RT10h4hm8olCuh4BjnWKQz4seJP8GlGKtMugqZZIpI
3g2eXrxu/leSwWnrWFVco1o2wjn9+yWH0LxlvgoKXvTZbWgcB0e5cVMavr84r3E7
B75EsN6no+djsqKFGxA9Kfe2DP6h4n52KREhOurRvAH9CycIwrhGdIq8+YeirjWt
3BGEcLRBkkD1217uo/J2s4QxrBpKhomPagG7Fviq/E0mvcHbo5a93Gi8IuaGjqyT
DDciTnUbDNad17NIj3w1JoEqDM3c8F2htSXhXcWNrNmrpmC8jJxcPmglsZ6uBC+6
vL90qlMeWjefl3RRi+LBRBReUoLn/EZxhZtYD9mUmxxWaFRCBSbJtL6kOQUzSXfM
gobETiqf1gwZwdWe+6gMHn9L0Io2tWZdmaes1vyWhqzCaIcar9PyAPY1Dpn1nRPT
HbSITzGspUC0JJYn34K1YL+qPcnKYH2JZTyVjz0K6x+lg6gcy2XWqK5agKns/wFC
Z0HiHZMh5WYmhSURxVEp2mb2R26cei0K7d8c11UL0+29HY7qlrpOHb7Je7WFATaY
XuSQwoi6h7cMa/MQG1TJLq3NvZ+rjpXvMxMA6kd3OAQh6yX42Pnu68/lsfRQsm/R
dFUrq1UDwYt2/+uElTaGG0pAuNlaPismby+IPaEUtV3h+cbrPpHkjVgB+qmKmxtZ
IsL9ORe+tJRKPvy8p02OA+qqidCJBdZcxugVrYoXhVNmO1/qPEA6H7DsYX6XSefo
dEyF2Qw+nH6RjdE9z2JWf5dfMMnCDGDIZCltkYSDzmtCsS0N5pAsx6Hoh69urQjC
aXvFO3Ibsf0hK3iDAPZaFcPtF2XA0nOAoqE6D3lTbE2rPeNI5gIZyNgQ8I1eBNM9
sMRfScN4d3fAX7ruBnIaDMXO7Z0Ibaz8sON9gaFoJorjHBpLpX/UHDV1DY+3v25r
sUO9YKW1HPsdg0Y8rEkCmTZN+fQMmiy7vSd+cVCMJub4gs6brDxciXy3iG+wX5s/
zvnxDlIvmNB5yJWF4r4X+QYIMrSgfpy93cCvA7QvpRDHdDW34yqSeSLHvEZ1+e2f
rZzIaB92J2qFAo/hbcAY6EKZOEF5T5nIRpxFbst4dgRv9S7urDLpMniDWRQ67WmG
GkrINDYYwoGW3Jl5/Phb2GgRNHPnr2mW8SH0x2eHrGBAc5xzulpHevC0L/ZJw7dl
RWlDg2mWaGGx6ZJeqnwE5/rV9/BrevkT8w47c1GEL96I/qrNHd90qWtqKdbU3q7y
5qsrJqkIYMh6cukGN1g1xD1d7JHCldMr/KghDC+yH5N0wH+TAZkq3nehxUl/USSD
zmXAeChSaiQ3bc+W//5QLPwoZQmB5dx71IS6EomPPt5HJtYj55dwGS9h9j+16mPP
7pzXeJ9DZuJ1aoRaJaBDzQzyaJjN4FOkIuCgwHpHuxBJBk9PyVP3+8Oh1fiQEG9G
kqcbzeGfFeJKhtN0Aewaf4FyL+sbevPNBpVPUXJkRV5K3VKXb5uf45xLjrP1xW9w
OmQHIWELQxEDSGUvZO9kC0mmLOA3Q9i6o+3qjInF2cO7Aq+hwkZGGHsub9FN1LOL
lg41+wCkrSmaSvsj5N/ARZxnpHrfopQysrJHNC/rpHYw/V0BgAASVbOJLu8oZOuk
9HFbrFgKUOnZTnO0OI2xO/rj80Yyi9x7a0tCHIaKQoK3Jm59M79Q8ydDro25N+Ql
Ehs2cQwXHkGAFA3WfJfTaHEFa7RLuq0pb56q52c23pIPq7oSpXAbNkgXGZHSOTfT
U69sQ/cPRX/X+qwH0IEA1BMIj72gWM1Yp6Sc31S28DdBhfk6eHSs7/0LDXQIMKRb
5SZLJVHFGtRaZhQysygS8Wdbiv23r95Ie1fV1CclcyfLFr52n0XYHV38fhrTgTRK
HWmS6n0phWaiCFjC13Bs14K64C86tVDO7o0AnvNsmPT3qg6jmOT49xu8ycTPO+yL
vwDaC0wsJtqjLPqJL4m3618ZOOco/liQjSH7QRAeBuKw57wbkvSACl1EVgx+NTZd
lxqeQeC7eHmAoPZdZ6jAOiUsF6I1PANYq3ZEp+e1VsrIVXH52QCmu457SQx7eH3z
oXzNPpwZ+WrcQjK/fs+zAKTUcoG2gTCLWaHaX8udAC3UJ1GkHrgK4O3SY4G9tbiM
msn8Xw1eGCaTcD53vy0hTt6FWcbY7GVoSTEBieR/1FdBZEsJdPfQ689XwTNkqqdH
AKEC2Hrmav7+4qBgTYmg57vahx1YKkYJGtFWyH5kRST2YiYVGyftnO7n4ZjrUBT4
5AQ5z+FB235wqn2LEv921sjDV/0iJHiR77RYyM6QcoljwoGvz3UrA7APJJlrgP0K
gbuMGqG2qEnkeFONcgkivh5DMz75Cgi0Kb2x2OA7qJTDFVDgWF9pu5VNbYluhegT
QWj+kN3EMQRhNAu/2nnswmqlfoGJ3b5aPyKI4/QKMfYLHesNRM+jdgBW8BK47BF6
pOAxJUph7Vb+2qLRqnhpyIPDsyJoW23KgRT2LFQy43/yp/WXWdq3eHVG3XPWOovj
mtmjsXn56fEvaSGDNP1wT3omBvQxhEfLEEPE3GO/XeApKvgov/hsrt72Zi1Z8ESi
VouDrOdRdBgWt8D9ctnRvt3UslqpvG6oVfnHCO3BFoh6DlIWeJ0AAGKbP/az+YQV
KxsVuOdrVo2NrbAF2ULyXmqGuo9f4lKOUULZ+J/77sq0RZa3yWXhcATwRJBgV7dW
K9My0kvPYN/0/H22uGaI5HIL6PurXUrhyhBCddhGWx2Fa2d6K587uhWr7K76WR2v
Vs43rChxeD+Mv5OuY8eyqqA8DEq/U8MxdboAm9tjwwILaK7xR9zgRIPIG9ajQXUg
lODU+2rjnDTJJIlIfGpPTf2bxrPkttQ2qbjuku40W66P8Q1kW132PIlvcAHVu4Na
hC49w4iAYoUJYhvxm7abpjHMdYaaRYirircy/K8c0p9pRKKBXlvls8xJmzT1J2kS
/ATeYOvZg4NVNEJ4eeFbn4dB1tQmHlX1cjciyJ6UuQ2dEoB+pFs/AGrBOeanPZDJ
Qbepf0uDtsuMzOWxe+ueX5g/jvZbl+NH1Yx3vCxCm3JT5m4mlqiFmbsCKZTRaJ6k
QKNyRM0Qak37qh11GDxh8xZi9Xq4W8f2RiPCPWqpm9Fcotw/wN78N/aoLbBLh6bJ
i+sZh4wY7lpiC/go3DRG8o7kAUlOK2CnS5GlbWUkUOWGGpOfGlmihmpMqw/wKNOa
1eBa38PgEeNlGwb/+IkfQ56Q7wgtXzeD85QpcuKprpwe9/kfKRBG965SfSABrRnc
KvLQYPjPQ6F3tcuVbi8SPM8onNxyauT2s0/NN+yQAG5mYUoUNgQKYwybscUuWmqQ
kdCdfGCVTrgKXz7Bkt40OKuTSvJqheU1omzCjkasKLRjbinNHJFgZ3323QV2rE+7
+ZX28UDSFeP6CaWmVyHnymwYwGzGV1ydQq7r51WE8/j98jjfdQEHUPFUvSqvbZk4
Q/34l6wWpLSc1S+eDfp0IR/wZMJqJvAg3Wy8Zs3Fzxk1NMThH9cxnwuJfCRhhXlf
1BNNszYb/BScKZN/UmCSrXbilnsZoRsMGaCLu1rrfomMHV50B0+bNjFPSVqpl4vk
coq27VwbrVabJIZ3iGqr0MfnOR3MBj1KYKeSb87FHaCxaExcdXo9Cm2D/sP2rwik
eNqR30wjez0e+DlYvDd2ReH+FNGS+JmK17kv3TD6SnJYcbrsjci7k5CnhxP+UCHB
QipK0pAWj3JJDMcvG2P3lvS8nbRg7dZGjEmGOkvJ9K5NyuSY83fQKxleaHVdoixA
q+d2Ifo2e6YOggS/qyUMbdDCbzuCWjtlYFB4jllfk8Sh2f0/s2MQKElSj4iYtiIJ
jckipS125aMVjTab7D5Hc08U907hDKnroEAFeqbLbyWuRHWmwTg5jc7yxH1yXPB9
tPeZ52EY6TZhpZn54Ff9DV5EoXHf+feDy61WR6aA37AbFutTPuquPsOZjXkFK2By
WycCfYAI6V+EC+5hCrtYn7QsXTAs2c2Yyqf8gGRBiMb0uc1W0RE2v4wiYqudKWW7
uf/cxdZdUvEsWk2W8hNridiIknF/FXzXbO6/pvowY2key2tyCmFhU+E9lmpN9MsK
4ikARFg+7nXeEi3mSucW/iNskS3LskLX1vFgn49SVqCpQB/UDFXox+qrtQsoWRdz
Kjy3nb8zXPok5c2YTvdbOEhL5jguHmuRzn8gMdT1zx9sPOmbZsjiWHh2itUZIkkm
gkqh7BFkTsFh7tvYznotv6T8m1OuPD8i0haZCFKFSU1zs7mYkbcVpBroO2MbyWXb
Kxi44ZB5FDVXlLCQXASSSNATQKDNF/eaCBg4iRIyToAm3VnhYv0bwCjhRA52hgvG
7YmErQumVchve+5I0qlAqEr1aAd/tsl7Q+EG+klqO8eYf/u5imA2xeOPy4IzvqKX
Tm1dfdL8wVUHulDJlakM/p8LSfmlBa1OrdJP1gFuCKZlM/V6iuLSYYEqFomTvY72
22aFOti+vaM5niyP3IdSBr37wzsQiPzvaGxKnOGRGS+4neYPINWTbq795PU25KL5
LgxSRZxcxPYLHSMkMLGqE9WsZ94g6D8Zge3vJmbjCebufpoLfsdGChmKth3i20jw
BDRqltzjvoaUDSGFMX2mVLfmEElJTL2HTkltJZLj03QY1gwRA3oZLRiVhIdbPgkI
C8Mx5LYze6IhW4QyGeZX+tIUxMvunTeCzcrWy/ldSUFpstEJ59yfIpwLGeHB2h7S
toTHJVP6uWpw6YnXd829Ubg+k/A98h/0tuZUojDLzpCSjWlgzDKnsP0FOHM/IrIP
f3YtCSh2u2umgFH+gcHIaAPSzeGQWBFfjFX1Yq3BEPFkKEVm8+OgaxJkiTlnj0QS
/eisWkJmRBYIrMPTRIGVRMUU0yJArm0gyFP6eeK/Af/bu0UzgoAgzWdkR5qLnLwZ
RP7KckO0FBTkj3Mld+HH8WvIrZVCDbH/afN7N3JW633lk997apR865IWz5y9eomm
ru8lE3eRnBzqq77qFgurhSybI4R+VWnDCGHc2DcdXfg9hjcrcq4z6PvhWAgbxRn8
0x7nJ0vIZ4YVGAC+JzGlmnSf8ei4mXbc3XIcrMhEt3jxQyQWpQJKJWM2lDjtNdWK
mn6/bQe9HR685dbvGkSY8il2GXtORjggG5ev4dZiYSk0S6ANGgZ3CfAJ6L/uqFgD
htKQ63e/RNQp1aHs0Jq0u5YZF/xvscHwtgj4rbwrZWU7V7KAF8CODLLpd3GL+ZLm
eAz5EYuYV6sthM99d3ni2XXudcZIPZpoa4aGspp9oIBWeiixedv54GuvicODPxXC
MFl7rbc0KAHaORPESU4DsBkc73LCLr2Mrwk2rzmN+PPi0tyqk7+beuSPhxffG83Z
jUMEZT4QcdI5yrx9FIxRiTTjohYCvWjtqpWHG4Cy6NbfaK5YPITXVVIIV4msdKJd
dW1I5Yxc+l13/R8ETCO0KmpJK+kp1t0erv5ggQcQkwOia4s1G06g7OFz5z9t+3kr
o45Y2piDm1WvMZ0/4kueI1LdfS+0I3G/M55orHTIMlAoN4Ssc1PzP8AbY6JzjbJN
IRxBDjX8Y50Ns+8kKHuomn9IepQVQuUPIpKaPrJjnnaTOoeExJVpvYDxNIDVv01t
SPWYZakyCiXHYl1ad9pxZDI+iU+r+xUIRAMHzsRCry2U2NKbx8qhJrlC9kh3YWCu
aML7SimCoPfbBP2mB8XYGonlnFupNpsuf67cAUn421Mq4upsuvD0UcQIrkIJMki5
5skWsPCY7NvyL6V4AEkp3WxOBxlBeLAeelPs3LhJLle4RWRyEuRWzRGBZ3mHfAN3
xbGxXOg61CCS33a//bYTTyLshZjl2L3zEU/TQVJJt6hxFYG1M4c+WEaXdO+aHMgf
qvYlFW0E2kmnNqBbcFYeIEPQ1cMcT6CLtf2j04qkkpmT7CK2kLgWPAwEtkLESnC0
3ObSrL+m6zBm9oZuo2qkES5dKIXZT9Eu24riInmvPJ/tjlW/6QLtuBHBe7bQZpZI
HSNY9/+oHdsI9qy4F5fe6TCzKLbQw42lEtD6KZFN9jPXc82e32Gc8Nq1dwL8nfrU
LyTP02DN0dbtrKosU1hWZ2AkNYzpQvGT6nc8wnfexz/qrWhs65Nff6NsAznX+LLO
sVzXipcwm94fJXfpepf4wf8Gtqq+T1MxMt09IxB7U95w9a++fnK9W8o/j7vgj5H0
u5gGp3bQ8kfcva/lEwx9JMZvxFvfe/EACLYR6FdF1Nm7YiXpy3jBaOGtyVby8q/s
8HOHuFQswhNNXXUF+fYBwTD8ej/FtYtNJskeZNRbtTu0wf/s29oiprjwxDwpU4n9
KTlvFGGPhstARGR6ZORHqR4exj3Jce5Uwpf6OfugmCTv1c7vG6jwd+EtTPY/O4J0
bTfelDhQwZa66fPMYtxsDA0TAtMje3DHQ3fDot5+z+r4mGSTxj6aUkPWhQWt3agw
JNoVgC2pMZCs7H+5tSx9WPKHrH5aPD93CmCYmtwg96RycAfuy7+ARGJgKek0Took
Jfdz4ZycJAn+ZBBP8a9yWtocOxFXLItOOGXSW67ZjE6FvLsdYNjr34k7jzVvev2q
ollGNvDsiuZ/ed0osYxfa2lFzhvHI82kQtG0nIADcLhHSpLuxrn+h+EEulNW4vmE
p+wRMfUZuCNz1S0MJRdHgrUMIYIkxJDkmc+yqQrb1yNwe6du4PRzh7byyu+ao6C6
VARmG94XtEqaEpBoVM0PjzkXQ5ie4tmSSk2hqCv3i+2+zmzRP1sPXjqkaECtgouh
hg3KdixU+ARTfZg9AcHxGmqts+z4RCG9BMSiRjfSfRO1PWY84uVkNGs7rSYqAHNk
aN5N1TEBeeLIrysGbAqE06OeNH3JtteHcfXJswssWMYLW5bPiepscU+dNn09yBny
LumKKyLivHrFED28yaIihgsYvNARWjW8GaQT1+BkXzK0l/BTMkq4JIRHMJI3UgCq
DvcIp10Rh2wPt6dTW8D2xKDoWpFxv32MjtO5dao/GqZ83fFC/SPcqmiOgwTmurD7
YqgILN9tD0Uocc16JcBBb1XkBgaH/CxOJT+cnSqTQPkb1aWWmzxFWCeObd0C697i
1lVLNKo8XfvMMjj/cLVIoPQAMlPLOz301Y+a5XF0+bQl9qtiK5rqKomB3JvE/a2m
CmTXFnSJ+Fi7D0d8WS6w/PiaWdAcgog7IQQUwadLQdGjhifp1kSizbx+6gABAPSQ
jcVYHWeGRxul01Kv7MZP1IWIxN4weH+She3k7YJf9UpCLcb/zbj4FL5dLAwGdFvW
4qkDx1yO5+Yv9FwfL1eSrHNeQn4jGqrqWG1nyiDkqT/vYeHqqd81uSxfSkN+vE9R
p48yhAgAjB/+XHnbshb4NMtiQTw/0uI1pnPwqIT3GC+eaoAtzwtDfdhgeH2GtcL4
7cgQ/dzC9puZ2UJb8VxpVlDgz06VA8G8YphWfy2kpOC83NBHdmOU6XLruNOCtaJF
4hvVFOt4P+g0c1m7TsbihDoGFAHyWqaOYgoBqVuyLFPn+DfbBhNckuh3aAnAc9Pz
rcoIjtl9gGRwpJjuau+OWdPgrAAf0+UQtkE85jdJ7WzZxxXNeRzQNwJEIIB8GFxn
A1iMTIdHZdToSwARtzj9qbjRxJ66ktkTr7Xme5zHGgBE86EYE+rJmfsJwql4DBer
rtuKOSNIyLw/BtWJ4NaOAca/O5cUFkqaDoZveJ6CZr4RDijfJeioNkk7TI8t3EAH
QvxiLVoAogaJ9HuogMAf8xJDNHcM+ehJWkN6Jfr2eQVlqlth3XT2zNMVXjFwFPYQ
BbKAT7nUqESHz3wHPfPN0RZ4SvGbX/2C0HMfZR/yKskkB8UvkaVAcTaqFjSvfyNj
z+b03LyHU9yPESt+LTYJ47ODNCQv0weIMZekC+1wpZ/8rJqQ048bTH+wrq16oDTo
OcLdO5cNBTcvUFBZNflW4OjO4KqN7O+tXkijb/GlOBRyUiYOJj6TO9i+I4P7yo38
wRKCv3iPP92EZzP5+vH/qTzrKah5ZY8UvCJk4o+WGF17UMlAulyvVhCl1zeUr+WL
qbEkmDkraFbcNSNBqKmzrcpyXZBlz3tQtbMsCSGJoIS3lZuZDpRxGNou2FMQYCW4
VwNKRjJXx+eqOTGrCaNZmPN4UdXfdajZKRlgHN5FvQNfUKFzYjxxeCbo81FmYOjT
DNb6Z4PHDZCXH7q0Sep7SzyUIVlCGjGKaLGMeLpSEqNEEMgaXaqKmHhxmmTUDWzJ
Ux4aUQWqbPX7O9ghdFJnOMaSuw+5FC6XqcpTi62qoV2vQb8rDcf1Muf+PvOd6V6G
e9ifAYGuIjHFSCbqZ22bhGepLOi1e8luQ6RDU84/wT9R22Ymvoqpwplu0SruT9ST
zK8qw76bM52PVDyjK5ZMuQzr3hoVfdGFxViGP0DX0EcsuvzilKkCEj3h5oRIfPQ7
BPtY+rH2hTpvJz2uhiKsd1damcI1bRHGm5Q8JU62pvkg0jqAZAgScutwicaTfD93
MoyWRRhHvjv/yThADx3Svj7s87ELLevHqybxBTDJBZKI6xcKOJB1JRcaTKG4108L
KpD+K5FHZT59IfNt7KNJRgh7D7tc1rJuIvfvZYyPy0dEMOLyIQ72cUpFzs84yxWS
W97ScmrIrwbu95Faah6hQ7LtgDeKNjpPSkW0CybOTmMNCsXGrE0M1fgOSqFT85uk
gf3t0rRg4DITxbZmO1bOauNn61h/R7SQizexbpZTG6/dHz0l56eBP/El2VyOGBIe
7/cgqQQJKpA9RExcdTOSs8e8k+z7MwKRCQnUVbbOUbvU5NPmxmqUzsC/yabOEo81
PnJ0tce4/AdrQyn8qYhF+f4BPKVwyjYNSY3uB+y5iPG3ETjqLN9p0Era498Ug3Dk
CjdX3dRaI2EkAwYfUzpUcoIjX5aTrlp1xyu3JK0m1r6IjBvvn0uesN+GNWK+gvOY
PEi2p9nW6UvfoI2DiVGeEtNodimWto9MZ/ZWNv0D01UOmHvlvqndOqFnHF/jB9dZ
aWV82LVzOws9NghNnE1PN23vq/34Rfi9FW80BjXjen19DhnGgu5UppKP7DlrsnSX
UcMm1nru2lezqpFX8/S6Ld6PMJx01/8no1d8fx12GBM3fpHPvdcB1El17LT/jRe4
rxHVGl6yWcNxC/7+mariTsD2Gm4AaBP3IZsK4LuZxbkDpJqUw0+PPJSYQl2ddUuf
HoZCYWwPFjaudQMaOJkUcKtaJ6/fXzoHp4nCQS84USqkexXmk61j90xWJ4iT0HS8
UFTvoA2RW/G3qS4oZGh0JRiMrZLwK9c32akNuMC8msgb3sxHC130OUxri9bvt11a
w9eA7OL9HS4zHUOKZPqfxqaNyRbZXEz9+p2kWOV0FXdCUbQwtlnZUtcPQ2JiR8t6
1PIugwHjpV/7iVpugXG/bNuLnLz2whAsEHk9ybMyTRmP7htcmA2CwlNs76Y8TpBE
u8pKiuc8V/HdzsPyvv6DGiW1nU3nLUVVIx28OmB9+lluHzvzz7nkBgF2NaBf0xJi
0ZlKBWf8VPqQEbGBt4zvV0GUpnGV5oMIs8adHz2840+UOsHMgA/t9Vuezx0c4vm+
pwzs+RG0G4xqoto8wyrR4ruoS2qO81NlcGdpPeCqyuS8fSE4xsjHyW+zsRyiRHyR
+Bs2YnQQOYM7GVGx8HXhUtFjCsbaSFWNLxrxZNWJs3Bqvf3CZ4ANXKjgQbN2K2Oq
odk3oo1u9Xh27obay/2U5fJbqkaxim/S5AAHie/lfIIeA8QyCKPIDQfXdnXWQJ5S
URTqXPDkWK/e0skyOoK+L55+BMe+5IqVxJfY6CEuod5vRr7aA5tTUh7MAmWjUC6o
eZdL4K0+y0fgsbhXZbQ44D2f5UrO2fZkUPP5zW6Oa048tXUErLvlZBcrG1LAz03S
Eg3jii7n8QVp/vCGTvCtTCbHSw36gq7X1rL35S3YJI4855vp7r6j5s1diQ7Vdlsi
UKsnapGQ20BTJHGhmVmixyr81nNek1mWrb8aXKNBURwem/2EdKo9SsqjvlbnPO/z
d20Ht06DQTTelS7BSdK/dfydMUom7JYoB8AzWug3YjVIogfZrTnr3rvayS+1tNQT
i5cMZzK+bORopnH5QUKUczaFPs80N6a6HmiFeMoiaiebh9xErQWYK011mH0sBi8g
COUQpFW+uSC5hqL6zxloZVGWQqbwpcdkd4cgz/2aBHMjG4EHTlVhYyX64qlsN8gc
8xGNne8kXAKbKdtZFNPyyGueskEZCErXBra2QA5nyB4v/VbLX8tAXmZhZpgc+Gxr
R1rOSV2SzKLHW48zm0CSHJ9mw93Ogd2FkIQcjH43uHlAvxWoTf7HkQt7P7NwWbK4
oMGN4cR4yd+dXmrSRmHuDpA7NfiE725DPZHvp/U1Bsw+rZUHhsevvHiTs4n08+0z
STeAMIVl5PgTX4UV3WrRMPI50SJzaFBWttGfoZsPe7OTml0uIbc1ums/3Cfr/stB
XJqIjc+WXXlWjTU5Bb+k4iAMkwUKKwDpLmZKssgJxLmUCbQBvRSppJsHkEqVmuuh
CJ8xrJEbsUH/IvOFFK1s3Gadaft3eVN1xuDWyuRw55yy4bI5nIYr0hsvdKjSs9jK
w1OptPt//1RJsJujptM21mW6i21LhJ75X+29uYXK7HlojPYGWyqL7AEPvFdAqWeU
M2bqX/Mih/ZhlNYGx9sSZvrbqsHYR40C9EAMu2ploVb6O0p8Lx4tTaS95avMbli2
NnfndEtOgomKAhscHuRCuE4G5oecFEQdrxAUEVxALYsJ1nl9/iUPZ1GTlA2AhHgi
6+fr2SbAIQwHWyVYOgbtp2j8b6uE5MP8E69Jfuj5xhZoJDvGT3jBmqok8PJaoZNu
97Pzcx0xKPF1BWl733LOv6FquFxGhzyWEoq7EIRqHWgxKhN0R5s4KdzG0eEl1JyF
nCIMru0vT89CjT1j6S8Z02EXDURru1R1CJPgeEygnKh3kOLTAEdRnDJpNb9+G1SV
n3PSlu1ulLlso4vyewCLmVaeYFbccAKJTGxGTAv/fYKek30Urzm6Qjsrk0fTS3Zw
MwOazhosXy6xden4TbiZJcM8nzjGx3ayXkA0y1x6R+QVEPZNEEQ7Qow7B1sevAO5
W03fgtTvaMrJVgs7qNGfAQlsLW8MgphLUP221TNcUehN1qeGZL4R/J4+I6kmvvEz
sZUsgMu9J7IoLZj5Rtx3grNPErTmU7WdWiBc3TNVsApNqYJc9WeQ4aY1w1DAOZQV
37SMHOdjDah6fmjz0ttqu4rfpO/bFTo4RV9rDNayntq8UofPVMUh+R8WSyPxeiUg
ihOmhWVQV364QzZ9OHqvCgZ5uExsZRi/GwbE8hm5Bt14cPnsYcrKKaTJW7R89EM+
Mqxwj+YcA+q1nmurCGu3Ve0nwVBDx+QWN27TjVx5OQA6RdxiV2EowqEiJg0VslFd
1+mJI298KInZ532RAn0IJMrB6ainN5NfNE+/v/6ANI+rwOrAJrAm72pK7qlH331G
J0SbF1D73oInF39bUd5dkBxbpgeR4cs6H+rvVxANqcXXu29VzS8i4AV3n1Ay16NE
Hc0R1LPG9wG235iWWg+E//vHPThA7aKOhSp8A9r8QWiNjh5lT8YslQr5lRyscvac
LCI6OOE9GJK4wH4Ps1UR5pT23g6t/UR0MNW3yTK5SHrcLWwHwH95gEBfDbh5NwLN
Q9a0u34Mm4DR3diO+LWzlefW7WQJLxeXjZlq0B0O/IXMD+iaO0ClL/yA9QAicV/A
EApAI7toXpdKcscdGwVbGnD5O9o97A8ukXpsne+Hcv9lWRT6P0azNLQgaELybdpA
yf1AiO/5fU5siGSxHBd/byZn/KTPtHISxm58VaIt7/sgn01aOrkc4bQ/q9U19yog
CpOPT0D5lesVe6/d2+ZhN58sUbH8ohskPgaSeVpLVH47/HWq1fJpY7vMb1KoqkwX
a2UfpticAJkpzInT51U9ZDCwfbtWN3juirBHBJ7k2sL/Id8lm7Pca6iKezoM76+E
XD+z+J0b/SJEN+cq7MZNhYsNWYyBD41pLUojDSRwfkWq+lAD3XW7Ar9iep3FDTUI
ngdTxG9b5+fX1e+JR9wjjl+n6mQ5hu4AZfove8G1SDCjODR9KEqiMrNhkFIsgREC
QHvIaBM8p/K7h3ypvGoqtsF/gs3inyWoWhlI4cLTDgGPKU9Xu+uOEw+MCRFSiX+I
ieivky0/1UbT4yikUcHAau0h3w6A9VNv5DZ+NArH33MwgUmCb+d+fbVqQ/It6umK
+AVTYRhPhCSktQc+kTT/Y3xg0nnvEEbEr93bqa+l7xlb207eWw4ORfvsF72BirU3
26OeQoMoKtCZPc4PBDyD65FjsFne835zLmgt6be8tlOf4l3D5eTCSwQvjNcHGWzj
thE5F3/0wLkjS99aAb2058m2AojzuRUOe+8Bbq239l0x6OYVq3DeOrUr6qVOBrJk
gfNYga7yh30TIWFa0rwqzp0tqwyAl6uty8LFtsmmgFuU/0FSM0iz5kn4y1FCrQNE
p5szTPL5rU0vnqx9mL2xaqz6rswO+YP/9jH+brvwgRJCHALZhGaLlqw/B9g5VeIR
/g0MtP/jaOrwQDskoQc3Iid0AMvdM3c4QTlzfjjXP/nyUdiUVUh6xf06hoZkhNlF
8KaC+ZG8+D61UxKaadfmMK6Dfio8g/Rm+SWbPynigBTeSwWXwIa2QxobVBmyZEHx
qYQ87GXqE35P8WihqiUY5Q1SFw6T4/bnORZefm3lA8s7sSX2pi8GoqHvzHajJkPH
eUqYLNEKggs0EvB1Z+tTlozxv7GDb35WuFFtd/66BslEb8UPIe7qLlGqQ20Cyfzt
Jx3wAlQY4Xbi/UryI3YxwWHwKKwjcQWwTdISwZoNz5SGnGmgmulBu9gb5XykEshh
agw6g0vesbVEbwaJW3eIcSVo5+aRX0tIvAJPsVNtgORR5hScy+xSlxuspg61K2Jb
eYnuusmp/n0qtf3y45tjhvHuV1pVl/fFxo6edqiBog2zK9RbpNtyEYE4GySjegdc
OfQqtmeyW9qJ3D1fI1QXk59j5817rdNfU7/eyhrGepcxLlkAJE2qTpXH4Qo//vpc
ZWQpBL1MkCfxQcfrgeFPQ3yOhqDOqv7c0rEWKZN0Gdr6mjQJihormVkDQWWh6FEh
TPabpIUHC5VZh/WA0tCYkBNESyxiaUiyQnJenaG1j49kancRqhJADcDbabgNq00X
0fCZzSaa8rT6itvxWqzP26cBmNsPLeUx+xL1HmbjyxTSfrmfYpNJzkVbK2pOl6e5
8FnY9riT40Lx1lBpfr7NR/fq1de2dWMDPdJCSiqUBbBG3sc77Ehb/77kAbsUMt/f
OJD6FLxJUmGkZS/nzdprtPWXSyNojsvUPLDD32OSxslniQrjx2yTCMkmPEESUsej
aOHt+mkdApnkRJWriCHe/6/IJycxz/x3zO8jXhFuCZkdCHcOQe8bsTeLW0cgHFBi
HQMIhxDd7TFRmlof2mySLyM+DZueUlVdnZBvkIQjf168l1YoZYF/Xp273fMwiD/V
zTai8ekMP03ZRwNMx3p55lRzAqQ0xFG+jt5YolS8DJM88F61NrWps9mlnRv/vUYn
Gjx2TjFLZCnVfapcnzUPpQ2PB2pvkhEM9x1wCmJR2KIVfGtSuvtX2D8q5iLouwxL
84UUeLSGBpTxInSeCs3Rm8xjwH0Z7mgycMRjzItxdqRwqE6i8YazvTIlfa+nVirI
eH6nyGOFZy8shCFaBm2h8UUveo4Z3ULMyhTlbtLlgK3x07pAhDjsdu+eUeik3PUl
pgPtzmDmr8pro0dYfDnhNUMKDYMc8Hi6epmm0iGaCeXwJTiWJogNWzwl6Wo2L2q0
zywLxK7rTM+v8jcj9tzXmVMH7equ2NEzYbXjrFRE0dDp55a1YSysqTaSQ0fMPC3w
5+atUo4H29cbqoOOGBt/+P3YePg7+E7BycnRHc1FUqfA+kDpQ1Hz6GojtM97EefZ
c91V0DxZt0Bu337H8zSXfWp9gg/6hEgUM6S182VPJlbcCPs1OTTgKuojIhOZAtau
l7uaYntLpGRRys1xs8+YMN66GDf5SOf5X8GKrW3ZofaUR/fqZ/tixqmDs38o5jBL
dXBUm/u29dNX3+9cJiat+YzOM91RcqRs+wtA4AebWYJ488LQzu7j5VpeD1Glniq6
0khwiR8hamruLuc9ofW84Qj2DkP7/Fhi94eYLk3oprNKKbzUQ/D/IdbNrG8eEauP
CJqGkCFPwFK1Wvl4xrp2uUnekpHi+v168gkfQLaNmpXkznM18s8RiJSpKPSJGzug
eIYM3Rg+g7FcNG39UQ7kuvDh3VW6anWsbdCBm5BzZTnEYYy4o0ttk/onqqpzg5a8
5j5eenyK/b0vXrBS3pIlEabmTceaKmB5NgW4jjalCIoeqUZ+I1bXpf7QQnVQCPfw
rA+mD3yLddCU7TYOpmLWDMX0AC06tDlvL5kc+PGQBxbMgEbSS2xWUPu6aaJS3l+M
OO32pZyr9wIABr3wX6sgvQaxfe7HFCuNhpmFcqZ/uc4K6QqFgfn/qeeuC2x2yaol
CvjTwIgrJCqMNOrz3hgxhN2zn4csR/n9kkL3xpFxKSZvkJOJOJ/pey2SG5rz1ipN
6AjmztORwgjMRlv9AcFn8MjqdfAlTXl91z379WBbA2uoipN2jGs7RSNJ0HctcduS
Ak1BiKgA8Sc9pQeZS5upIUbar/b9u69cAWZKeU1hL6NnB56CuWrPertsI0bTZuHM
whgp991GTXTLfWNDcW9WLKMUgIOOycL13+z0M7Gz5Ff1R4ArSTg33rfuH4GkAwey
SIwUJdKzgdihH5mPgXzDk+Hk9wzumTz0i0qy+/F255bk9psd7/vluaeA/un+TIGR
aTMdd3uiKv6At1lM9sjxFnLIJ1IbF8rWonEz+MueYRKlgmaLAw6HXhVVxyV6OPq0
K/F5gNjoinqO5dMPYyfed7BCBmRWCvduYpNwYuCVwfiEiP8xWghqV8zd2IWbkR5e
lJ4/h/A19O/ydDdmS4e2xlRepOKo8n27DQ6uO+Luo0GbN/rCERwrMjl4qI4Dsphu
Q5NStLqk7pGExmyA8jl9J7fOMy3ioC51RUwXndCjmQ9AwC63J0OtRAP6YkcRbhO/
WIGa6Lb5+o1GpjFWTc6K2aGlLvl298cTUqhrWsEg2nAOaW8fzVMNUzkEQENiQKNd
P1kcRnxpxvSW22P0XZ69lu5MU7QiTAf45h3pA9jsGfdAeAzIo79zToKnySIP+DNw
24wAdt/IVdMLLGGC6GNLjSyRHBthrgmUv6o9LopZrD0l4fqAyOB5k8EPd7RJU2/t
tDwxqQJZunhzI1VbGWkw9302jmtt8pUeJ1AeqdHNfQEDTXML/q9WaoN2GaRhXwp+
tO0vUgxHWH212XeU9UyvYqe4/JLUZIaV+kjXP6nmJQARPiIK71M+3gjoEdRVpFCO
bcxoof56UcU6Yeu9N3YajExFBLNcFoZlVUD15fKT6vkvHlDh7xxHWC3+VjOr0hm+
vs4ySTXfFKNJoRaGljvAfpdjm24kzID24NCUGA2g8O/IAnwGkKWfL0JAjAkE3x0U
Z4V9Ih0JAzIwH16fhrMwctVVGxbxYtvk03FyE1h9hDuyiL8X7IAb1/6yu0SbSitk
elhSNEjAPp9wcRUG3byLI9RROly004CXhdju1aRe+H6gg99BZKc3j5MtC12YVFH8
o5robkr4vbfCwSnJyjU5Ma63CNIWhnUcMWzt4Bv0TXBPAkvbNLKU4eHITG59gi5k
+WfUrMi9TPiAJk3Z7KtBZI5yCS2+D/ITjj0teCrAD+Vku1GCZijWEq5c3WDluXgG
t+CPmVmrNH35W6ohWQG19ebxJlB3TbmBlhvas7AUAVuDh9Ymx1laQ+j6BZJeFXTn
dg7xpLCeIhRr80O+1rsbjvGtkJRwwtwUqCKgCJ/5vka+64/fy9kTNPBb5IihZ3c0
HEhIJCZBiNJguCpERwdagilZps56PiEVvIFsC2dEQxTL5O7qlisN4pc913BiXV93
SBBqA+0Ve6vlXu4djjJHr0oCWttDQ+YiF9p5E5A7fG247GPBU1tbW5yFFVmpGhlT
JaauDjRsfMqPFB9yKLiMyatGbglNol1l4vbDroxVOITUTt8dJ3UkI3JD4HFKIecl
POKfpLOwHR924al0uP+hBsTcqW7p2ZgTRCfQobzuXxQL/csg+wXlhqYLgtiAxk8w
a03XmjQ6Go4nC/jlOYUTFrhJzO5mOBt5Bv2OlG+UQUrsynO3Y4/wFow8t7NSjiTH
FuhpR3UEZExcckfFttPMyzkLlLx+STrBqca3sNzjrcL1Kjjw94thsJSVBWXBiA3M
Fr3AA2ODC5lE4bsENXfciwnxdyQBavmFAxG+AhHhLl1xLEt4uFclA7gexIQj9NKq
Wpu0an0NTKEpPc932QMmmd3pnCW6EdxtLp5BdllwC01i46ywVrPec1bCrzK7Tw13
epX4QnyOCfa28TLT3raQCY/6p6Ln8sWPNjQDWEu9patQortjSg9GYXYJUWpoAUCk
ePu/MuTiePNr9e9jdIhK2nDUAP6aX2/fwnngXEFLC5jAel1SMuHrIS0GQ+rLbBh0
7UwSbaP75sA1s6aAHhI29s/ov9534KojyW/W+9oqpNuABRLdaCR7BpuqtMLiOT5W
9E1aIuFaADZV5eQjiXCTI10LFBI+4dO2WOHjfn/gHdaq51Vxto//MDgQMEenCX9B
mvFU8ICnJ3GX5ujkM+JVb0okvb36q7oGVZbv8WPCNcV+109taALfAaX/f2Yldjyd
Pt8hkBMS8qrcaM2oYCtadhmY0wYIHEtCwuAV762+h98+esJKxO4allJm5BZUpxGf
GwHWhNvDPNM64a2X++4QFzpr8gZHNNu/bfR7EDmk1jv8/BEPKHVxcA1fcR4aUf5p
wcTPdKwJfBXp7MJKhH1CvIhF6KVJJqVgtQSZNFnKrqRIPas14cisS1W4HkuE94KY
moMC/QrQJhKrXwzSysTynkvGZgNDDbrZYnyUreJlEpdo1kIOE1VID+ClNgBpQDKZ
Lr2OfQMo3noU0jdtQ8QwloCfxxwolHVIO6r+L7pW7oKzoyMs8uGOh9GW5zOlfgcU
4svX7nURxonPdKB0vapvP1n1pu0tojHiBd77cJZSnb5KFhHRwk3DpumT663cF0UJ
AIxLSKRh5LJVrUa8TWZqo58euXgFEAY4Rc8oI+nW2txS/i4hlMlS2XcX9BQYC7eA
ZpfuKL8dR2+IjdCWNznm01AENcwYI0+LqKqSBnOnxpnBaD85WNd+zeANEKQ6PP9z
Zyct3qlE3MQY3Wijo3vwVNrhSxwrkB6ECqQAHSGEnSxAMyP+Ckhy6cw57Z6XlX4+
vnXwkJAG8Pn0rG7rv849jSDVmJTTqT/bb159jC17iIKUy2dizQT93mLRUcDrgn/e
C9/0HcpMXXcbfZnaKhpnPUTvii9SFtIqD5uw03QXsGpmIaoQraWbZVrDZGPbUiRs
0dp5PRZySoRCA0fhE6PiBZnanyZwfH7hkpESVseNR+/jeTQNoww371ZCgyvQHyVk
JnN9qx8gsH7L2OLjy4HNOxB/P1U02i21649Ok+IoQak2PnXk/ISryUqadXf7op6U
HHY95izEmAsTkDtP0rpSBqHPPxUvEzNq9cFZRtuI/P7wkdXrFJlXlEFLhkyCyRM7
DDD+CSSck6kWacus0+9t6Xh0ON5rWfcvnDwFVrhH3FSuJVdRvWXc1JxHyfWBhL8D
5WTI98KNBlx7TSYKABPakLfZdhgPS+twrxQN4rjIcCmLq2eB43u4BnGmMGtwPq8s
QLoERgm8m9wQ5Ot+9yZgZHpiuy0jQD+3miJ2oXfSj7br3DZFVOzUnXcQ52eZzINT
kQdnl3pNmuoH2LcEjXJ4r+S1yncjGSd+8z2gf1UH3DcnVhs8dN7ioHLgD7F7ZARA
wtTkUJVgXHh0tYRAGaeCVbre4Q/YeN5hb6GRGJE0Wqj/RxbqeVAiGeywZ/nvJrZn
5FUf2YsWsbaZhUimRxDwcHmao2mWyjEi+9ZRqUioZz5eupe3aRTSxwPKeDeV4NTw
S7yoWLvw5IQlkSFQ6YuFybOgRMbkN2KcEkAvqIB0hUrAyr0H+0+fxzZfv2ENytHI
SLpH0WmPaTDIf2muLUwAnE/NRK5e/70e9fdTVk+bcHxs/5kYNUZ6C9hF7uOjSYc6
goT4FbYLfmDcKWmwPKe+z1xEmV7cJvyCyJjz3y00OxYkfOn4r4ZqQ0MyS2VvV77D
O8d+0iZcRoWzK4r4IiG6O2vUmFD2B1AphCPA2yyvpqAZbIqYcxKzZJP8X2nOC2ri
Hyr6IgIDMsh8BgUFoVZmeHOTs/4x/VtZtduwSwdEWizC9ucpoK/5wzJNwqeu9Og5
WPWcR8j6RoAIixj2mVwY/lUbZcMWs/UkjKnMbYcWtS5D8h/H3jesum8DLoLxnuPW
7P0e2VDeMCvmMCCTSSpeQm75DBoTO7D5z1SfEGwBIZsmWXtzl/UFLIceaQ8zmcAv
0Flh+U0qtsp2xv6krJMgIgnl2V+OxhdEAIgpocVN1ux0QEatj3UYVGAFJFXzhLK2
/C7VR2x7I+aC0hBqAa2xPm0qc4aN5/10XPe9FORILSfG1eohJNn1//siFrcRnf05
DPnDGL3tkBpNSocl91i8ZJ+dkfFWD7FdeF3U1+zyAU/J5my/sB00uMabw78TdOhb
B0IYLgCbvdm/qPOr7Awkf1/iRnEJD4We64rLSPFS04WrRn4HJjYjsQbDUbd1vqUB
lEyJMK6y8EywGOxw6zgQA5gBxgcEmrPlmVDh5Uriz1TkapKmTcQVbOpMMe/L6dXD
SrTZ/Beotu5q/EUOEYN/4KL1fJVQlph6W9ZGB9huVY7jXxvfumbIMpnsKZG6gBzn
Gw2zFqbgnDASu/wnD7+SRFmxyqvumvHYXY1wJmsNI3PFK+yhCxM7lSbfrscf0Utf
+0T93SVG1hhesSOwrjUenOukqgIECNgQ/9oZVgDys9cjUkuDk+3TeTdmvNIuAw+k
Bt6GeXE4teSKMc85mo708hRNbZJaqdkcvbyTpxNvYp+pzzbw2A8GJW0FwCV6wAXF
HU1MUxuIMIPlp6ZR5OwR4HCfK3YaeVRmLW/55IF+K3SOAQu1z5cnw8nhrjmBuSjw
N3gkRyvdfGq2IwdicqvAwVnmhxIs3qOSxmx3Mcpq+itRVJ6Wuo1rIOKSA88WxpDt
8EBaNpmsuwDb5+holTAiVSZTyeuZ3MnD5rYfLpKUKKcFiawtChUXKQnljPJxG7Oq
0Xev+aim0F4cNBmDzKS6xvd1nJ/SrRi5LB07kKbXjllQzn0zjRgm7cKpIjwawJbF
vscEUAtajBDYILc9J3Ps8MXlZ42FWOrkY9EOi2NGKbFW3jGldp2AQpCWkqtDq+tt
/sd1grG64npw41ES0Bs4ZpSqVA7ZGM/JFvIZ/9pXpmW/i2lzzWmO0tQ9lnSfyuSJ
wilwN/I+pBPYSrgZubrvCNCFzSzixoB8Bv3Y4jpUIpj6HSblKYvPTtHEjyZMJROw
pEF0dBHOttdZr7kdGlChwvNZxWmG+QuT7gV5bMMBr45hxHwe1LlrK4y0AKcnEiWE
pNUeLtcC7wRiJBv7xJM2g8pBTxszzFMuYd6i3UE6j1qvjLDqpoRP5ig/SFfifGns
zOFUKBm6IWaNgMZJSHFG70KV8LeC0WDdMUROfyJcL3fVTSbCsF+B1l/NtX5kYCmz
sLA7gHUsVKSRnIdV6bbk0G9zSuIszBoNfprmHay7lWC3M2TIPKFoAGCXDjV/O4Hx
Ys7YVxt6xNBzF0TyUKE94Z2iFsiEtlf5jqyqe9v26zY6nnCD3RTSEmHClYbWAKls
EcFXJwP5WlX4Z86ndUdGAVjOlVOCf+3Zn5NMdPp3NYjgzT9ut5tpXhE3hNoI2OPB
nQTEqaEHyUdl8mg9Z/nBh3yzTlHGB5GWgCogjiq8kHQvCZprRd25UtHHx7M3YYTn
wQwUbTwJnXNRGWg3dxM2aSMXllov/UZcWZd+IoY7g7DLaujaTIu4o6e7Fmsaog2V
Rt0ZVj4FIJZZbNboru31Sd7GvnLd/gD5WPRb4MAGioUcVtRfj3VONOmXPgIm3qWI
I9GNaw9W1HbxiTROxq3oYCIp5zyJ2fxnLoOAIOvvNW855TbtmM/Y2CYnWfP6pPlx
RfDOsyMPQ2XrwWLYbHkOCKqXEQ5Ba0ejfL6VZ2HUpCB4p5TmviBeITdj+6EnxPgT
fZuosrk3Vj235qG4uQkbjmmbbFBBJCwCktKYAT6DLpYtN5l26NGs/o5KTTZe2t0I
fj4HPxDOKOAP5vbqM2FOO0DI3YHLrc7CUpSZBPBcoNTFCQcCrzYRPl2ZbDXGtj3Q
tpg8cN2pUe12QO6bKpU2DjRJQcJyGaeLrblBe6K14ApGRNQbKpUlFPSZCZ/+lWRb
zyZiLqdARVmY6jRxajOeqFDAVSEd17Sl29SlsVALKpwibj6dWWRqEuNJieIQ0Ohn
LDoz6yL/2unsAImxEri7n0FWjT0Dszcpoln1hptoyGUUR2ZOdpWhY9rVoiNunrS+
FPU6kuZJt5nHevOiMv1/08ipNRyVBaG4xL5aJHjm73TQ2iObfDgc9zBEDZNYvh2G
HqN/JuYT7vTpXQkRkgYDzcebNhWv2ELnVZw99qjHGhv12R696DuACi+NjHrjYW9G
81Ycad0VsRiavb5SFKCIlUDesgQV/tPcuQwtw550df1+pwtr0meQtqZf122FISpl
+wGrkqdvpJYtoF4N2MLaLkzZh3pYDbnWduPdnJYeXlzC3OdqVNyLFWLq0oQ3D4P+
gZvqCoeWCVxP8IHPUQKPRsBYch736+L2Q7wt3vKIMVxqiMHBjxGsIBXGgaERA73W
YzDHEoQG3rn5B7ZijGO7xIGwDPTTxJrKzEHhl4mWnTBLZfEbgztUQLHptPtfqJsA
sj9aQsPg4cAJPNrxGq/yPtWI4grmvS82Z5JGrVF82qFQj+CjiAG2148yt2Pgp0Uz
FUwwb9CNBlcEP9mWUE7KTwZMACcbScwTtrH5qWWXgy/bWCpaGm3xHahXze+oEGGq
XYI7L5C8tEV75bNHy3yT//yRIH8StQnAQBsQDOi393aTxliJF3bsVc8WnE51GMpR
N47tMxlVLCIVSJuTb62hLkoDqfJ46aCHJEjjVLFDV8ysD/KIYeKSaS8xgjDiq9fP
0Y4LeGFiZZ46m7BgygEuO7CoJ5cGvtyS4G47VgKJA5H6GoLrj7rc2U3nJ3diWYme
ah+5xs171ZBVs37QH3oA20eQWSIlQHLLesK3cG9sW2tOaZ9qaj8wIqKsdj1qbN8T
zi6hMrynYuV9CdiIBhUu61YWp/H3pjHKnt2GwI+lBPEiEL6tppXueUSJau1Msuxo
omh/wO8k25RNUsWOAtQJZgZSvRoYRPPj5Fh4F05X+UXNR3VP14RTOdvE6K9K7yUg
XyL+0Ri/7jF5QWS4pUpgjCAGRDaeAUhmJLSLUHnBI7uYVSGtJq74MvNRRluKrVtG
MDmcFpZIry44+dyZP1zLueAf54x5BMMla4EPr0blbGRibRmN0ioMvDVE7n7XW7Jp
ySCqIqwGbBtZQ1AlME1KTNjyfi601FBxOEU4YNsIAKowGznRIcknj6Az9Dj8xYZv
vTzhIix95n+T/76d5ubvKUoya6tEX0H3ax+qizNyykfoL3x6SRo01SSjxWmhP5kj
9nUGxD/GOd58t8ZOA8V6jOEuA+CplvYTBpFkt4luu9O2flqmFw2ycI86VG7FEJMy
lLOrx1MMyMVhHL2G+jmimR9tw44c2P+fuByQDvdhB+MyIEt/gOPb3N7+9ik8Pp1p
D7E7pHDr1Az7L1DL24IABKN709tKRJHi/QBP+bn247MWZkTrWPy2djPkG7DGXHTe
QYTO2yWVU8dQLARbfu1hcB3uczvYM7tI3Hq+VXz023zfCLjh1Th2jmE/OL4aFS3P
YpV7s8GsK2kLRGx8+rg5rN9K0hHzLlu+B4fDzHnCkVf8aRhNjNsKmyzHOtdZ4g1y
Ah7bYWiiRGPCA59X2wYGBC6RkL5cdV4IezKZ1peZSzcy+0xx5VCxehLy7IMBihND
jBz5eKS4sBWFoVE6ON81gssDCURQyJ6Jc7LKz5HPRJ3QvG4JY2mupiUQMnvUHkZu
b24MoUIFN8C0c/Jm3oAX6hB9OT66BQ355EhHJSqhP71Gwp0BeuRPKrt2gGPSNLLQ
nOf9XbL6HE/Zuw0RuEXl8TTh3wi9Roqw8yyvGcmuONei2bXHh5LpzQ/GCpo+umeO
gh8PXdEQb0Lkc9f89mGqzWcVx6RMUiJxkKYyIC5WMxQYnddkW2IY7g5NaSu1afjY
8NF4mfeDkXc/3tfIURy8nn3nLMUpQVjSXLHmCZPpGyykMF56tPpvt7r9M3gi8rWo
fZzg6U2FlpJlDgUZndTuz2tnVY5P1vJjy0BEONxmf7xgIL2GjmBG3+RBfWWK8RQI
l8MCWjtFjyPD39ws5/conidx7wXPmUwAPEZP96zGDGE+YzbuYEmsYfSWgwTDTire
erBiqaxRWeDTtAZH5dygGl9trR7lDfUqz1NN/+UlacQXNDE6KBhfso7cKQK/C2WZ
eDdpVcUMWJnmadBEde3wCe0FRJu7lE/S+aHS+ja3ZnFi2JT0ZUh8cF2NHTj9iPiG
ZV+f/HdjZK7N0lsRisC/W8J1t6/4af3Aed/2EELGpP0QDH3EGaGIlIWKd2DVIkCr
DJ+WURM/z6myW6y9MMj7QpXhBgQnQ50bR/5eeAm3Rkf5kSxwFNg3imPGmUwKzODW
N670pJEzJGfmqgSZv3x2gINQ7Idr+6ms1EcIiK095fYJPzq5zUaeMST+K1vMjCPm
ocy3XCaqXup2P3exenKPaIp6W5xRdeDmQ5pxeJRWUBYUzxcWx5ui2zmSnl7h264J
CzcYpTD6fOusZ15LpafNAKGBtWC+yWHa+ehU20N2CRRMMVy0NYDfbq3Ta5/RrYXk
FM3H76wlfujK0SOZEnDgVhic0TT7JJxFy4n5U9MJ1Zpuy4af6CCEHLoiOhUNygPm
Qk46vmv3VoiMfpAa+jQedIiWWWYVAglyUD/hSHCXj3mEysKTODcLEd1zaEacVkjN
R4+bxWff98gBJEtH6uylVal5JuhEMK6TvUmPt2zGx0NxLhWhJdVgO+Kb2GdM/I18
mlw+GnepVoPlMARw/sCyVMVjgS9LYDdzHeYKpWp2X4hAQWHWYy1zSKSI28USuFqm
39KSpZIwtiwz63KBTO0BkNPVG2zDR8ER6kf4XJ+IEi9U6usPOLqidX3M3P/eUn0J
ophYGEqP9CIBK67sckuHFSh+UXdJxpWddjRQVWEAtuA2GLyUdQNM1/eFl582PeN+
hatp9c1hTCgzWENp6mQmimIO0GaGHXP/5gtmCQ6K1Z1g2WRULwnayLjkaLuCQ83B
q42x0SW2/hYauYIb5h5gcr/58Z0IsDq/A+7wu3iryHZJKwMxwnoelYDz+7zMbx81
+2yj+bCG1B32bYnsaYNjCMVGHq9GHzwheiMt+MIaD5lMU03ipVk37kgg+fJknq23
POhqP/OFnYILIVSALH85T5LxfGXdlTJYmeapA8RJg3d9ND2Nfs9rXCpX5nAJbTIT
74oltgrHTwZMi14bJXyr4F4g9RZ8hmEuW8QLwgNR3yOxWV90b++dr0gjpZzE5FUA
8pgOc6axPJ4sTO5gUgecNhhdlF6xXwB0ebrmwi8dsvJS0KBVBra17W0WKunDPwB4
n7IrPh4obUj8YWFW92X+aQWyABxMzjV3dK0OSIOMHdvwOGsLhlt5y9r0iAVv7IsT
R3FmcfySC/igNrmLWyYziWeT77YHH0NPka65pSUj16QOf5igwO5j52ABsaeoXzPs
z/T+tJdttaSSdSChd+55/vT/t2nwNBGtxQApWmmxdIn4laGpajR1iVmrVZJYbFaU
aMG3I04nYX/LHqGPkjvDLq5cMhBUbvmJOr9zFyGYeB6Kbo9tsLI/ywfuTWV4CT6E
cKK55PjrJLfGtGPrdFCbkaCt1Rz/KWlQDGHm0avWs8KJmdcwe8JBiXVDTRGqGhcG
x4dJGaJvn5AOedPGsb5mOUgDKZGXW0xX8+TdpCpcwhaYGDZPle9B4M70YW++Tyqu
2w6Wu/teDIf59kuUdJdDdU3PDPIne5rXwOQRPtCTURWuRNlBShvcI9JMLbp16TVk
falFh3pEZdXAafB4oHiFIC8o/ZxbqW2rf1ScvcZdpV/huJxYuq/pmebsDXTVaXiA
tMX5ZjghUQeiMotdAx4rtwv/xBGtv3Wjf74S7V8ztrzrkDyMEqgBlQqOojJNk5en
r4pHkqUEbfh++hM9Mq8thH0xof1ZL8ogfIrIaP4c3gF1W0/Pl1NRt3eJsYpD8ZjM
lhMSahABfZ1tbUJ2uu4Udhi41bOdUe9guHS8nu1wOROot73fhAOf8oyLEccgzQ0m
EjMZ2V/d6Vn1f8sgE1druOPDV3Zdf2y218gl8kYv7SyR2A1fdYYmACp6DHR4owUx
fszmDO4EfTV/PfphlG/ehHPjU9Wj6uDqtDo3jy6mN1LHdJ3MhcBo1JxJotpysnKU
Cb0XW3wOcZgZeaL/eVaMwcU89vvVAG2RHkH6Nqef+daE/bqfRcbLvVb+gLwfYdZx
s2ceenaE5D3bzAg52ocHxPg2M20mZ52SMXeDVKqQ7+gZim7I4caD1UyV3ma0xUF+
gUfEdGdZWd8zaHwbAcYmDHq4KlajX6dV/lOQdngud5Pd3RjaFF57U0SGfto12zZE
uS6BaCltXcr/cQdG0CtB/EpbtSvdS+TNStnRRsPV6BtLvqJHZI43/tqxbPyftcnI
qUCCVGwNJ2Co1J89pgTX8m2bpasOcNlMow6j7lsOzXadq+arsLr81cR59B/VnWrm
Hwy1iLIsGU9XDXJmHFI3bza2Petb7aYf+IB1xkAv/ztcSQncZFu1JFWOxCthKpnG
HKSdcn/wme9dXVmpK9ZVMJa4acZQy71WQJsQHkBhmi4/S4ZJivmi0qlgpKBCl0iB
Ywr5RWhS97apOCJAB9I+TtA4mEUArI9TEAjtYqjsG7bXNo1cfksTRhe5+BvHJ3Mw
J0LaZlg7+LM7Aoiq5kNvFigdCeFD9IdY/9O+3RAy13Q8yo4Nfe65C7IxnUmmGOBU
KibP5xugN0uxdwIntqc9UuU25FRXZ1m6Wt62fhmJsE/WGTFFf1vLDEMsQX2AMISm
Mux4vSFbD+OYgN66edtDgXwYsaCQjOH3O0tBC372PxB5Okg8fII1ur1OCT89SyfS
DQFZ6/BWcxj5w9fOPrskBvgLpJl2k5ibAVVY58P+KGF1DZo8SdCDMEz8aXBCjwKP
lDnK7X8unjT2F3lg0A+5GLNxx2UAR2Nnspym/UU7DGmEaXSeMra26FTBuUkydg84
sM6Mgx4Xc50vDHou0LIUG08AF9NGvJD85htT7sqxEeU/g01w+1Zok0dUKyZ+7MbX
wmihZ11GS6DDZwU3rtMooxZQl6agqgAjHbyZ8hYkkZP/n9D4jIxXc0k6SQf8KYgS
TDzkm+Cpl64rZDH9WaYe3XFC/2Ff6J8hFTAFHWVMypwZOZM+qT9PYezmLahB5/P+
q0uUiAW06kNp7E4gSkivAKDEqyOZRG7xPJsGM3Mr6ndzXctR13piEOIp9knDmyzi
6OuNOMYzXqmri6UJcrdyD80Td5/7SnSZ1Zt+xy9tp0YgKxZkRK9bgq9bIz4hDTlq
Kq2aklAna6kDIH4rXB/+dtPVnV5CHCVblVS9wCF6F19i9BpteepKG9HX+zDOGo+L
UMHacK/bXvqFSUa5mNP0dtDsVt0huRWsapPQTS0ZT0UA6Fj0D4hMo/7/u/ZFOzJX
ghcWO/JlvTDKPue9+WLXPDCfN7BO4438oZvnhKWI9lG2wqKBlTdV8Y6MwdOgNYlL
I+K1Jys0pCqLuYLePa4NZahxWNblSFLOyrlRkvEzcWvPRmrhf33JJ54u/IQJG3hj
zcc0ruJwx3EbSyvhui0KYM+a24788qgYZI5TBWvdToqZnZtljS1cydjZxIsWmTl6
wgjQnf/SsvlB1k2vVOoDGj7qBEJ8OgSVT7FzX4czKiG3SHMRXjjj8QlU7OgA4ClI
FeTs+EokdkxAnTxHJUHyVofRvNCGDoS3g/sIjueLVmDvPRSjEUI9WEIFP42YPKWE
IMac8lQYGFhaWzAkxbL2sc2MvTHcYgdshVEOTBg4IGLe0eqAN4W0iftcb2GZfhSA
+HKQRt+uWNOdG6ZON9iRzJX/u2cqEXXt6DJdHmP2Z5XrWtlsWHkJw8i/Z/PbC+zB
G7587tiu1gvTkmzgB/MJMPLFTBz0xsZUScU1Ph8f7AQlM6CDh/zsKVeZr9Clg3IQ
0vmr3bUF9wrlExVhM1EitfOlqbVa1l3Drdq2CNWO7YKlCgF/fueppCDYH2X2iMSr
FO+25PO3W3qCqOsKdmNrDfCrb3pr13C8Cs3oEsdOlVFS9IjnqyJ3GZB52mLyBS4i
4e4XlN1mkyNSSt3tWEhWlxLpRdyLtryI9WMlhafUGmYr0dpKoiRAzLbCUNV2/pZR
J+1AK7onZA/1dMX5UQnS+wUECwpJZ9ibmuH132SMML8yfGwE0xnDYYTnf1d5A5zM
7iQnclFHFZMkd/cTvadgNTKMvxZvxJDrQM/gwUSnpYXYHTqRmwA/iW5h760Tgekl
pfXkp95vbZTMmURDCb/6+SD6LKxljcmFD9fwRDiop12V3MfZAW7aWItG941ngXPy
ixaTURWLFZAs/fb4SJcjq9WkOCMPT+uv4R9Tu81vOuTA1FcCrhdIUAo4dFTwX+8v
0Pl77UNz+qQ48mQmdAND7KsCkg73D5ojBpZvzNFaIYcRwIgQhX2N79s47tkBWpLu
VVSoekun+9G2e8Sdiq7po3hByehMejEKCWkGR6R3eHAdd/RPgKx3sXuQCsOmGtP0
AVoTYFxnGO4aWQcc9v8qJYRQa6mmT751loKHIaNBn1ReIDtjWBRi2HMFQmxlwCED
RALBL7r6F/zl4Dxzha9FVS4gkNRBnrZyXu3z5p/CRppK7GjlHrdL6xHksyHGTA5U
rPZjypfC5LXWpNG+9v7m0LL7w5oM5QwMrh7t8UXXNBqI0Mk+jAz6gxr0BHUSrvlC
ydwflDUqj+jZoUhn61HRqdnLFfUDacmKiISozDBriaeYj7/3CIJzSjglVkVWbwJt
e52aKXNngxSHpuxbXTvg0CTJDMjqzwZsAYccgK3Z2P7v1KxeK4QYAwFAeVkgIBjq
3J94FnlTop+VxJ5XLp+ZA/cwjY27tfAD9+AT3G4I6ccd8fMxiAKKGXWpJi7tfXbx
I62vbltHGFb1AWQt6WiodeoAf5tfYYU4Vvjoy6jY51zSnmm+BzcAQvBKFHprJ1tb
n6TnBw8Mjjt+w0CKjb2akbdXO7KglZBcaeU9As8QwQm5RTrjwRsujwbqMd3HXmFU
PwOE9VhEPxe7FFIA/gEyldLyFqfGLHX7UAZgWc6OUJ4HmWx+qVbAW8qTOOEGfuNM
8DR/auP90qeotv/1ei+szhhicCR/Jr7GpIqTzSN0BgNLrVL/uNP7A8/FM8iBby7h
oPa4Zm6VPVwnQ+stYKw8NjfeFs7iCjX9qeCBnFA4e7Vb8WCnhPhF4uSjVLg6Xgyy
opfSWkQ1g2PPs5W3AaaH2D8tI2wkLPkxvjAHTLnh/t6CesMvohyDZWH9QqVJ3hgo
gKyIdeKblJ8H7JrDvmVkhdrpDTM/HzU25KvR/ghj51At4Es6sUDcDYP1dIPBGHkA
aGllk1vcUmZ8y3gzbi3eUJLRJAXQ2HRmo5PSAjzgzzdDZWvna9KWoqcBJaY8L4qg
J7876y+kLxC7gcf3Sx8MJ+fAgPWMZ0Qrrb/LG0bqueIetX881GRwIdjRtf2S3QSn
l78rPQ5goHBhzLUMVNWazl71p1G0u8w9UZ9VFI5XwCS+L9Q9dgaDkzkZ65aDQhai
IG1H+LCbP9+1F5Pqy9WPBMiPUUyy/P9LVNWhjG2ys6d24m1IIHaaAdWFbrTSPxh2
d5xaKogKaiZlYUt+5Z4TpM1LRMaswvkBD/uhxaGGucSsJUPmWR+hxpkoQ5I9KDHG
e0lTlDzmcZOwkNiWFj7+okftyCJW7dLTPPKtNoIXk5Qwdqwlwu2Bgcyg2JH5Wsdt
NJcGFeyeYdFI5QgpyA85H2sxsTy+IlyOMnr5Ig1qPeT1pT7kYqQ+M3KNjZiI4cLM
1WeECU/bJDWVFc+TzZJa26okSHWn/JD0rZ6e7To52u5uM23ymY7zMQh3GJBt/c7T
I2vEDT7scycHakxwNLbNOB91cvLzqgCo9SA/DloqCmHQbAKbFvDXFv4kJ8NVEtE0
CtVmifEBWAi6YXJHsYfjsGMXmhD2DJeZ+Vj97MufDLQsSiR2ANAfvNHCQ67eMnk1
J7Mekw86VATIgv5Y53Jgs905Y0R8bNHo452qTJFivNTidrr+etE84+ovMyijgpgx
WZe5sVJd/tE28DLadaYOS9TQ4Dp3sWgP4qDwuT8/xnhCY9ajtZD+kvRgXEqLEJE7
+Gl2qjLRFEqpomQr8yvlVno+kjCaz9Qlv//UcSHYMtZspAL0YOauI2EA1yvricfw
dfShtQ/FjXLzPe4krIK95V8l6bqA/A5alunAUJ3qNqVuDGb0S0OXjT7e5cOdHL0i
a1A42dAIAW2ihjzGQ/hPPBlz2PanqdFFxPWHEG/bj+IsQlcFhKKFpAw0WUiWc3gq
SkSWDSoSzrIuXHnA7cGdbOO2dfi+vrt1vkwFQfkeUUQYLOZcu6FZYOJKBZnbJlTT
fzF9SIOeur5pQWyxftFw2sMKk0MVTeRWwyb3uJNi2QMwO4OIrDiEuOHx4FqardIg
KOL4sciO2lzR3QD0P0Wy7HlA5czU4XdAAyknDQoZNK5PNbNYQzkBZF0+1uO8p2Ek
5hzWsR8WHx3AsM53YXMRUnCj2tCWAsfXR2jEcrqugT1w20czetyNgMRxvThZPG8O
ezAO3GwV+l6XYhKnL89E0J/fEEADr+S5XLXHmRGPuDVggSZn818+/gZw5a4Nasd4
ooZnnyxbiIzsknsPUtBi3FVAlnyp3UdsKtB5bUP5/YZO8zeqY8sb55KSHD87ZdJF
zCHmOv6A8V8dp2GXL9k/YC192k5h7qq1if1qZ0hBLtYdbLhKMpZB9vmeZcvd8Q2z
tWdT21U0/9H/p2QnT67oTNkSXvgtnsmzHmLTHKivVJAEWc8RwbYOGFmdUWC543Kz
ZBCW7FGzhCWCXXhFDqTuCaR6hQLN2wW7h1mayzuxxW4tiTIOz4xiV7M1YfuLGi7x
bT/p0dtlBH9eYHunpsS45+lYQxUBx7hIKnidQD6r7EDV4nJVmMzl5qcbuPJQM5Da
EgqwvuCqT70dxMb8u+LPaKqx42xrTxNiF7TtjB31FlJEGiwDoFLxSv3IbnNOog/a
lDk4FIEbl45R3HkzTgyzWeURgx8uMDez+8DOSsJOK9CgjLnlEo/R5Y8jULPfoyqn
q3qJE6fGIW0Kb+SzeL3WV5QB9NOHNqa9SYFJcMccwEY0BLeAhBpczmnNHhI5o7mJ
AFoQ3kCS1tVlWsm0A84To7TxYNrru972TWXzKaa0iUd7UNOgDRyaFqxY0PuBRCbB
bdSnfBQe/8sPdWX1mfAUZOjp95hkpnmKstH1kJ0QCYQ/bYMFqad/GD7B3H+a9DGy
kcOvCuAom0QdhIGuyYMRda0jLfzjPjXGHiqJ2vOqgvKi1r/FGMkgCkCtiaBat9MO
Ju49Rv6qlN35uGehgvt0MsanBOs8Q2AMriIS6LgKski/kGU/BKAYqymymMypeaXi
SVFMkX7CipNB4n7fP+BNKq+CzhENPl3Prs5dni5lZyLtdlMB95fun01HGAhT4kif
Py35+vrxuU4bi9S9n1n00QFyHCRJI5CZP+pY8uqZHC3UUtFXtHJL8E1kyK6dQnDM
eElk6VSpf5mfS/0QqBUJL85m8IEKnRO/Tww7SGaBfkwYbDuB4vS3QiXpKO4DcZHq
mRbbIq5JRiItUd9YWptHrnYCSW5FRpXreMHilVZcOfeMdBNu6L5GI8E8uZD8LQ4C
cFjWP3O7cZlI5dvEHSusKUk55eeVTen+SZuaE1Cdx7IXmwvpyKOoOVMrCUp1IgS/
C8fmccm11XoLbX9UOYrp0defv/ndFZ9iQqp0gxq6qn3u7OCLU0BL+GpggbSxQXCE
GWWjEENn9QGbs7MW/NLeE5qNkPTUwQ4KbWwN0VlrqJdyycsW13apwhMXmvvfoTKx
YlFX9FsS07aEEZtTpDXlvtnZxewDgIlsa0dyb9TU5FTx13YFyQLUv2x+tXySE1oE
b1pohuYrnA1XCZF2yDcY5jm/c5i1KCBeJM1qzlYZ3PrtPlDLfaE09ZBJWF/c0+Zo
eaJIzG0mrLWpzNp5KSiT+7zAfp8cBchLphVovtGgQKtDoK0MvWG2HNWe8eGlUqZN
gDAhoDX60mot6oZtwaeWKRM9OzB1Nmwuiq1lYZ85qzj7BynEyvIIbaL6vjxMiuwE
EAUsyGKlOTLr811kTb4gcwdWbpw24pVu5jR6iHoly2BlpIcpDSrNUApF4NZVJ0k5
HK8o1nDSlvqz9BLyx4sxDZu+q8hRu1HzfLlnetw+ULPi0bj52dE3T1WkXNt0gO68
AiGriOzqDpwyGY2siDmiwMWds7lPElhtnmvnCTVFIHNXcfo7TYbYek13L6PmviN0
u5+byUxNEH6dL7NmV2MvZ1iIZyIlhMcFMsEYIcFJULk3Sg6TroRjA0AsdF/MZI24
zJinfxR6vTXPg8iuX0hztyArKW5JyKFVIhkUs97Am2gRmDoKNhATp6cYR3O2WUcg
3vKU8gSdZyAEsAK+daipzHkbWc/918iyi65JfUIrIWZ3SXVLngmr4YMzNvTFPbrR
8mzziH6qem1m+wdVTbtwRn5m81A81ipXu/LaTj86seGZH+cEQiwrvWsA+odUsJu/
GyK3HkQJR7Ud2JDr3TYadqKS4vBhPn71cF6/HelE4l89GBttbmXxQmaxbArGsc/t
yJGeyHyjTVyULkzu/u4JGn94EYyoVCP8JGK7IhsiTVSUOQor0pnEYuZh51jpKl3S
zfkvkzIlx3Y8nUK/XVOaTnVyAeZx3sQVfdKbP0NiiYVT4vjIgchbsjlPL/XXewhO
8dcjpdoWelzYQpZIhxK1bMUN5CwPnKXQdafWe0LBSMkxIYWhP8HFwopoLIr3ivjc
KCFDuG17Fnvj/EYIGQWigDOZaEHMaKUflYmSJQhFp2AvHFftG+Tk889/h5msDXos
FhX7biiyDDoGRXf4DGAyhQZnwqZEXLMYszSrQdRzAZ2l5mZ7mLmXILLr6epMXqWL
V4adZZCJ0n0j9iNmMeEtjSfg1KMl3sGxwEf3iwU8DqitjM0OfnXGH7+fIKF6nCNN
nllunP/7YIqq6/JXiQgo+32ym1JHB2qRrkRC3RIfs1pVjZ0yZLEworf3gTiNMYhi
mCnTEefe54E1EAS2e6no7VNCrKjn9KQNSYjAWb9eGrEn0Dvs2MnnyZjOiL5nA9Ow
NaZ3l5eaPnrCyXHpXuLneVhpff3IA6GqxvERjqvPbO04lCeUsvR5twLuujhhOMDy
7kI/ng+xav6YPcbBGltT3R+/0DPsV6ye7bF9+iUaZBUKSGUw7Y/GWeqdgX8GfhOx
MmQYZmqZ8g3RjQOaLNNmVprK/ba1cFpCZRtLOxIZteumINAACsX1lguWuIPvMGHR
Hu7vnyL/jsjBgYLxJox4ZRkYvcvg8cG+QzFkFZin+1NKh4lD4dMUTQpX+dHsTj+o
2gpRWshBu+dLxOgJuWMbxiz2KzPf1ljmmBBWKOgFhCm/pn7z54oGDmM6v6d/odYY
LK3GYMjRkkDR65ZqJSeTS2rNgOiZmoWhJGpeTrYbF+E3EqrwvX+0B0vMj0/sxtoz
rPix7+k/P664EXRj0y1H7RuCo0aU4cqndWUVbx6eoJq5ywR4EAsrNzuDuGSdahJw
9IzQFivYG3LKwiY3Ngkry3MypGMltlWEg1UcYb1NrikfIkSInCjh6ilPzi2UlLWm
a5rIQ4M26stgmUSn1awrKjWlrT9j19XE0VaFCcvQCofLxg82Mox0FADOuvQqjanh
1pS/21FGTfswHmvob4a0EKRMt8YT6wSFL/hIT0xC9vVdxEnZrwDo13nbooNNqNAM
y72X/zJZ2+bfo4PrFiQgG+u64+lVbPFHF+/Xy5oGClV6AMd9CeJYa/iUNWcbkv4L
Q+5A2X8bS/2G1aPxEKzzUfOWzB8EI1ZpocAQ312bH+wcTxErM5sS3h5l6rvxMwIL
Wv5LXRSwipuYiHFX2uquBzAQ46Ht5miOmdBQtVHpeM3109PM6ydcQzcNFJszyxX6
vnjEBizhomZ0KucjpIvPU+nsgMwYAU+A7ujy3YRNJIUAaJwQDM4pDt9hbU6l/lTM
aNJUR7w6WchbeVgZ+hjtjXVyQtWukWRYUKehhrwoqMDU6E8FFp91f6L5kgHISkWV
ElfdatKKZUcVofauMK8LQfXvN3huOA4ILmRvSV3LsvePvXkmZ8PG/N4pwXPwC0VM
G5o2afJECUn5VeCn3FlfUexY8qMwDFa572vyc5OFw+gjgzs4o25U0pWFeT1Ej30S
YK7l3t/4ydEv7g69YdqpY7LcyoXjjOJ7nNFAvtm4gThwjeIaiEMgdycgs0on4QpO
fTkujz9zXaDZq4PYg3jFdN8wPc8tRLq+SCBok82L/O1WlZd5ZkB/mExu1iw9tYbE
jwd48c2ilCVTVTfm+ROnQfXl1MJ161UMwQ3rEPuZP+/myCcGezlT5uC/052e9CSs
Z9QsY6B1ThAR9dJ/mPeAh0wfA1lKf8QINhAHMfcvwhOi0rNobNTgGnfBIj0Fxhdw
Eeku/dEWUSFs7kjmU55qTyWLGdzU3BYv5o2PJdqIYis5yw/jCM2iTLrBsOCB5sV2
o16OIOUvBaGZhg4Z7YpvvnxFJLxd+YL5hVzStWOY7BgHLRImhgLhe5CJiKQ4hOQU
YFvXa2mpkvfPwlLDicHUVpi92IL30OlstdgbGyOLU1Nct7QkG1GPiCV/2EkHo2BU
mZB2luihyZ7CxYxJuS7iCXHSngyYAFt5hMtszi8EEf1/9zxXgM8S6FtaGjGfxu5g
BvfxCoQ8tV8X4VCxEHA6IvvarRkW1WSxNghIR8lj1aULZ1CSNQbosjVaPhstjx4i
hjnlipjqg/8agrgt9wZOhFtUqCQNhpoXayoxcGT7ArOSUgnAfM9DPtbm4L4Y67Kx
rWnLp+u1A8DX5LBazDH41/AgPaEa4cdEY0sE4oxvY/g+KrECVT3vejdcHQYZgcTW
vf0wEI+r2OBAV40GC7Z1vkrAIgJHSn8LCU28d+uiy0iv5ycXwgYoVp/PReGrdqJo
lpSO5D0gMl07qrg9FOArkytNSt5hxms3RxmjKegUzL+RACGL/zR9m5cHJdOfsM1X
QANjcLCAInoZeirsw+DAvPxVSQlalFVXYolaZOE/ON12UlxBGEq5q2S74bJb60a3
NNMT0UOfacQN6hTLtz3pNTuP6kHNrvs7qu6vn5i+6aNFf50Ggnf4VQEuIwncrxb6
3LjuArTZGcMfNTpu7nunG1l2rEVxtxfjsu+GZqHycGoCsk0IDlmC+KkmObPbQssx
YcDq5Zj/lV3hYGVyLOI9guja5TjaVIxYNjN/ZO3yqC1YnqBvTaQi1zF3HiTyAZKH
JDxR4LYcdYSHMN/aLArEe8GbmPXysYO7BHnzzSL/3sMMDB/7pV/nIrF7fcvkb68t
tcPtJ0SAkpBYdM8f3F3AavWbD49RYftbPlYdjd4tUQUT6/M5GD1qZZy3MpXbYH3/
43JOso6uGz8VhxHMsiZ5aX7ytiOEhan/Sf7TwZjtmXlsI37VW1RPdK13gStcqUGp
j9iC3vHWTvA1GZhe4CqdkKM3kW+pF9h3dfwiaQDbFFirmmriWZCX1HxirFbdeIsD
JzFoAHJzypHPXwX94d20pKOacWzDERXJZq3KJKkjcNl4K6Vy8dmgctTWWGBcf06M
MJY1r4iYeFwulI30d2AZhxFAcy3r/VsERIGeBFXDV/n4/6sZjRgPx76FLWjrbLIx
h9XGXm0eiNIkODgTDSgeeIhtwalZ6x4CfN1CRW7ug6+DOihJ6UZnDQ9Lvi/uo/7r
TbSxV3NJKAVx0jgRVY5YKgNCoWcJxQdYgTGbjc/SIA62supkQ+44CHHjvkTcw9RM
ChaCxAFlIckZq7RzzTdPKT45ZGo772Ka8Qa51/++GwMkGGyaAuRwwi8sw+kMbQwI
qrrKhX0NzDWkqP6biR2CtcYgVp82cT5Crr0DlJvcj7qA5Jh003FN0XJHPTKy5GLR
aKJBMbru7S9gdJUwKDjs9I9KD5yWxtmGhgy25uG85FSbziBDvXm8JFN3lYqf0nwL
cPkFk+4gh6aLkMHBcq+reGxHoTleB5hHXKJdvWlif2KKGMznKfDDQUDW6Hu64MmK
AVN8AoNdSIL8nyiYmSLISgK9mwelY7amsdgQqhBP136Y27ZOtogKei704jRMe/gS
Io45TOBkHYE24QD80JSZ6nIgbrguuMuFJTn+z97MODX4EosZdZJQvfSAVeBTqm2X
G4Itz5bO0BcOME/lhmg96d4dZaNCqRFfiV9VUzay5VQlrTdS5/CSB/iQVwi0d7Jb
QuGPoo3jxnxpvyBrUGAZ5vt2aYYzS/7zg3LnQmce+7Y+RfBpEi5fsSpWUcEZXEw6
/lYjy33+ie/l1X6loZ5HJAlzlkxI2a4WDaAecCoUt0eKGahWe7NYx0Fkz3CktQ1m
0DJHZodLNNudWYlen+sk3+gePjLB3Rb18SIsFZLy0X3n6rmqy7PX/yCXUmKM8gjx
JmliUVrqmkDC0yPZ+kpaw0bk7jW2i1YsjKR22au8pNKJwKo2jaSYTfyIv1ga88HV
vhlf3+GtuIJJA9qEeM4wfwOQJNIC74etERlXk2GeD2vxIeshA//TsTRuXkIwzK0j
wafi1bAhyfGy8bnl/xsQdJO321OLnEbYok6jz7qRqIx0HYccO0w1WCNz856I2jYx
oCGADxZ4oXiEqGlMQTFiNWksa4qAqP7rMgN+AN864dIWe74lphN8BvuV5ujJ3rtD
EgOLauDrH41P9QAmAsZGpARn/GeyDZ3p0HmAi4p/yURujImB88aQnGdKBCbTYNK1
F1oP/D8gcg5ZeXSVVqcsFxwA1IVKepLLgA0MEMEyOE9QXc2ad8/3lPAtmZfZ3Fl0
ABumIf3O7NKR6vWUuJE7upmlr0tO7I27fSw30v/jgCGLvOF6e55My8EwaePPHTO9
hjA7GOHcoTDOhgjgE0eisTYEkw/TiKnAjsPT2BSxPf0+YjT8HYYAQvuJsTuDkQue
J+5Fc1/x4VIAKVcL1/cWVI3huf+leltST/lZK0vvnnvISo4J7KfmV6Fsv2kWiGRj
uB16Wb7+EspG1Th2xIGJWFX5o1ufZVMEcJyMq6L3cfa7TikCDks65dDRyhGCz0nj
DtW1xvHbxj4LqQ2RbpdgJrFFcYIOh9YIZa4KvTzNWdhYW2IdFJ4PiQOBPiAoFHsm
bqF0ajIDaFklvsD9q7Q7ZYADgN0622xsvZg5MAiHiZd20OXO7O/FmSIiC804/VnM
ePTh0G4aUmDEBu2COU9iPcDMgPfzi58tN4Mi3k6B2wnY4NgmW5GgpB/Yc2jCzz6r
HwTncbJIakNiyrmkT4dSBMCs7qsTlMz5Ofumi9/1mjf/NcyHweUe84RKNaFWjW7O
dN120I6tIWRgCHK53wRJG2LPnMdqdYFO3tPPZ5D9goQPHVbuxaTRjSWXqUOWGLy/
HlbNaU0owtW1ERlAOvSr+6Ibi+AjAiyg0vdSPbslWUZ5wbCdm2bcEKivTMog27/J
I0ziLEDRcZ/Egi+MqY1jNYLvsg2pJoGfA7QWsT5qSMWebrKs+uQFkdvn1IKWglX+
44nHaMUazeHRAB9N4A+sZN3xLgDPDDa8UQYz7Rdswxs5TCfeVrIhpomVVigMoGf1
NyiCxAfe3LuJjMk41Vh8sxevNq1OMd2v67HALAZvYVsLnlL+MLPIor0o6oXzbOay
WUsHIbRHu6xE7m0LC1e+57MGo6H3gxZNe7WiU2kAmsVRXmtGKfEXabcchhHeChXa
mzsKAJaLCAewYBXQxvVcwmZSpkXSMj6XpbHK1/PwET0Am6Z20pxVrAvAyKCgdoR0
++973UveM1G5IAJ/7xgx6uUtOwHNOt2bv1DP5OgU4hH72q110FDk1DUXURV5/rYw
88nBz/gic2eGviGo9Av5sL+N2nPRQCuoi1EiMnLDMXJXpMC/Klmf6ulJQvwA0jns
ZnXTmWtZbAU2+aW/K5MYGRgPHPd6vV/FQ/O1Dm1sre040F/jToJqzZVj2PPUIlYE
rr5XIVcAMoE1LcW3fFjo8DI53Gvh4qyOioK38b2Iw8txKOUrcVWkXJEnmzt2Pi3b
7YbBRt6IErZ9k3sDRHzJ37O7vEy8OK61S9qbOMVxuXyE2xqfdTAECETjFTFEv1fp
wRLrmdC4ToVIwc7h781nFZQT+YaXzinMFFgtvDv65EjdxF2umq6RJHvIqt8I3v+T
C7r+QFU/3qNBgKPb8BvR8/JrXE7Nay39FeraNpiNrfpHm2U/Cr/xusvTGyQfyZt2
E/XKyugkU/JjShRAyajH2ZKjujuYmhzX5V7jj+iRAPt7LlEaFdv5OK+QU2A+1tI1
GhCt38FT/ErF//f3vu1uotANYcmhItGjrwqsjZZvXiVYqwVxx7zNC/1fqujDjFnF
Y7syW9T6qLObYukObzJZlx0Coi1Q122L/BH4PSWiDFkPijQRVq+GfPEE8TzQosR5
MrdnuEOpi4/Ibb0v+++udru92L30pp9wDkfR83cFdD+kj32BOLqOwxiRZ0p0bnVD
lBqZ3+IxVDdqDw88Xm9bJBuJTIPRMDgcyu4aJsdi4HBl3e4CnRWVTXm4PN6CfmSr
UkvI48rZBEuQwSl9sMav/C/hjgqRus9t0zS5C5OsxLw0INi7ASKnYan2blvBcRRA
uZ1lq763UOMVIBPVzbTtGaFKLSFSO7g4QfyVzfJfWMs+s0dvCetPdLE6FywgR1Q6
hAqtpuHV4t6mUmb/pDdPCJW4Czl7WyZvLJsZi5oyVylLnlQ3TafnntFSO0Gflj9L
yUuZQpCVQG7MtZ7U5whTcLARVC8tHca8kk+e4yg/H2Dfb9PPKu5mqxRLVynXaDN9
uIslPdYucYzFqSc3dSnuRc9DGsFoBIL7y9EBO7aEy2E+U2cmWZZFkTZkN1pjIli+
vfRYav+jO0R6i2db9uIJUi9kK39tkiH/DeT4o431RTnjABY8Z2tAZoej3zev7vLu
jVWIVKRP278nevfD4hL5ruCPeZII2iTiWMqg3D8eRfmVcL/WOLKbASIMky99arYC
ZfYFQ2LFYFmlHhtAoqcbYwM8UJ4/CL+H74VJB2/6jxbneCVihmxkz42xnaspvf3q
6TJUQLpW6cB/aRzdmmV1DuWnCdXy/b/KU6fs4oorP4HosJdUwzKTAWQyZvCQ/b4w
eg5sR4sJjd8Gn14Sfx5eJvmaMEgAq4tASljn819yoV15f23yt5uLiRY11lqdXGXV
4mVsw7hooW2s14B9C5hg7lPAWM6XtXMnQ82KgXJ6W8nN+OCP5Kc3fMi9oj/8LTjt
q602SIfI1+1rJOz9fHiv5Mz2zbWYGQ390SHUAZtKhja+IV7kgrHl8chPU3a9bIRL
HLZZVtJIgc4pRU3Xxu7yJ3IdYCNvYPBT47J+46QhraI3JHXpG7ZPOthIb3uaX81z
L3ZcaQaTM0dfa0bElxk+6reekvu5kiuUJwP6JWA3Y7Dwh0tnM6TEh3fr4RTmygy7
4rA619DPLs6R1ma6vMF7ceTfpD+qhDG6lX7LeSuGbBIVmyOEzXHE3+rAvg9+5M4q
NIEseAh7M3iGIDVSo2rtLPHSYMm8EnAmxFkZ5sxHR9Wg47aEdAbgK9PkfsIkdk67
0WMBDoKMxRIbxW8MMAWRCvhqiGkB08e+oCIrsD5whga9ZNBNaxB7dxj+rRU8mEZG
SVLdYVvLOxJCapN5O2LK4cC/JBD7QM4A4yAszb5a0Q3KbPjne7HxTaN/odjuOG8w
0sJdbkfFgK4jo2yyLmTtnQMUbUvE5YvSeSp+ETHva+TtDofjRWA16afiEezFGWVj
FC2Ap/vDvsZQcBmalgjVB+6z/UP99v0Po4BCjYar0T4N+VzWZGqdLRagFjyCGfJh
NRckB5cqj3g2s2v5J23ES7JpVmQcr7L9DAyEe9Hq0iOSZBlVgdruy9X/Dsxkx79V
XlGJuujMLrbmDeG4HQE3PDp1IPZGjevtRLW9wJ79vPdTGthpusam7obMzZdnqes6
Rp+NqaqSARJytZNgD/7ZdE0sXzBv1y9bZ8hsh6dzZV+GkiOz1cz5ryVMBnxzBQ/U
KBWPk0mDiMtDa356Z9eIQTDdJ7zG0bAsUKlADq7wyVvKSP3/YCjJvS643M4Dl5Ck
iwXQ5Aet/ueyXJJPGCrfxAECZC1izI0NzApvKKGBOWR7RmU6g/mBStvHfHYl7DyE
/+zmAR4Kk4vy6NarAsL+klvn+4/YuUegdXPqrz2zyANSyWbk5kYCYWwe0UpNtEnN
qp5M6uswxuua+ddSD2ngk0bNSMiPCyZEwMvwQqe37zmnZ2bFhP7Bm72Hc8v+P9S0
pud4dQKmCov1vEaLwCdA0ApINTU5ZoKJG9IfvddVUm+JGTJcFs+wojQ0VHjw/Blo
FaIncaxANMR2hjVm6nfAgmGLXP+5gjbfHB0z9gMZwiiZPAZlwRA5oH0DAqnxM3dy
nyD462uJRDnHUngHmuHitV3ibLU+v2SgvZvVhHnD2J3QHTnE3d9bLvD7GN5Eo9vE
wfAI9sd64jokfqmW9h985VcVJ8c0i0XeYvpYDun5eagiCnZ+Ho6c6m7lRBU6X8t+
M1xGnI9uUsyJYn9rkUQNPyuyfCU+Ppwoc8qXI3Joe1ON2DCgOt7qNTZnvatlX2mq
s5VDjZd5fCCBl4jZNoeSjRJqjETh4Fcs+bnLkf1kDkOmAE6hlZg0BwKG1oDlOe7r
CXXcgZX46+gsznY3Sx0psZr9mxwHFgOdDwcYO2qR7NLhPvfMYIPhrTECpBWv5P1Y
kBVq+Ets7TLjzhapShauwPR0YbO4j1PoiC4/WXsYsWJJFOIiPgPzm2o4Ii/HjKGC
1+DeExPuGHzviWBJt4lDX1mbtXOuXvTRW6JaH6jq2OLZF06AFGoS6RWX+NxEZGRD
lXyvj137BDNj9iwZ8pCopdmP3MxsyOGg5eO2BnJVNCfcXiq0NVgTvzVdJujmQD+Q
L+gFilK9o77+4Wif3i/fv3xaj+1iijzPQ5ue+G/5tfLNoHChpYRLHSQy0tycGjMW
1LT+3R11Lls2JGWj0Hlg8X7LFH2Butku31BbmQj5fN/xN6KMmmvg+P6shHIIpnZ1
Uh3j5PjWlCQGul5CCBeoog/TlNx3tPDwvy/rn08WdjRcYqpvWJID8+777p7EUrBu
IqlUcX6x8RTdebXvf+0M3oJPR6+mu3SRrvFh5OhEkz2LY6PK8U979uTBZKhgbFwC
NSQ0+SuwQ1oh6xjspx41t39WKz8+NtHNQ+0BzRahDAUWgsT8J9cRXVJQ0yidsKH4
BYaZ6AtC41VblYIbttwwkV3BHR04M7MLWwjmGC6BZlC1KbmerAM6lHPFRbRDiKXY
JOA/edSrCbgVcniGrX4siGyiHISGioFUQYRQkUKhUWm1SXyr73IZSx2bXWPFBriF
CsnZ5WvX/j6NhuZKAZcntHPw9H75if7E5ZpRfT6ZgY/GJkVYELE4DB9Ds120ar+H
7EvsIbbKMayb2Ni6a1k8RZFjk7658UZlrTf0iI22sgNOffC5wczhb4KxZbhKAqxd
35DK3MKEO9S4GcWFLSe9WS5UpzKLLRnHqbuOMDA6Jz0j7rxFFYmLMQz1Zo1BZwie
/CO+6HLIdmkII95T5ipW77q8hOhl7MbAM4kOVkqFzFcT8pGMtfbB3zz82dfII/9t
IydYtsgsw1aK3M4QpegkOrMvVoxU2XVQjOl1oSC0swoTs28MQpvpFKPVmDPk8fe8
Mf/S2iUvatb+rOPMnsMJ2z9Ogc/vp2XjjYINB6ZzZvCsEF2i6U3T+vtu5/7Wb59E
v1PYp75t2hLW3uRzbMcbcq4iMqQaBKLDz2YDOd3OYC2jVj18UVFNw99lcTk0vSGe
1RQvOpqkmauiotaAMk9pbvn77Eb3rM6YYOlw+y8jfoCeBpjhgG7kXrQ7m9My5wFr
Y+mKplSsh79hdP9ymPz7k0QWn+JtI06YX59PHQHn5S0UglCX5HedTLSCjHUJ4jLp
quHrCTVdKAyCmzne9msfdF7O9es4W6PUs/EFsrZii2BdW6kpGpkYzGiSX1gHzUTj
qiMIDLp7PMvAMstlg6g/xm93+HcxebFFLn5sfQHrGNaOeXdw2Ley/wSLJcvfUHlB
03x+fgG/CMFPJzY5V667zzvQXgPNABmoMXMZkKxlH51blGU26w3hvxMTjob1AAGF
wEFtdppAWwTHlLCA0lbhKJ0vRR19HcIubpyWaN5SEX+gL6ijJ0NFvVDNRFSuYlcS
gNW2YWb8+ekOjgoPIRuy2CjyFwnbOLwc4abAoKiuPhBDH5PKZvsxdl4zZAQVD6Gs
k27cePfrYrqvnKUORXk09it+YJSRzgvcNtm9fHAZmxxMkZ2BanSAVTC9tR5kQe6S
prh6QaTW82iORxZC0yhTxRPmtsEE2e6OioCChlhXeLHpzC5n7Byh0ORTF/6k0e02
tD2iTF4nouerw/fu9RqOULWl2GljoUF7yp4JwHMa5enUKc4GQfJJo0VI4ikygxYF
/wYHCZJM3olrU4JNIWFq3gLaG/e2m97STD07HTTtEAfkl/ioPQaLmL4S51WoZoE1
og9Pnoph7seBGc5Ea2Q7mmFe179xR8lX5VWH9sH7+C7FDUN8uU7jz3NhMNJ9PUDl
NV6NLdLjyNHFQdvgg8vWCTQLNYdRufhnNLti8CsazKhe95kKp2/miz7jyKTtjzy0
QFoJgrr4HZL6cjkw3os9skRD07R2eR9qtWBouJkvH5KEiwOaQafGPj+kayvmKcCa
PM2wSiIS1vrNGt0VjvEPNW1yT+m7wR+4hjqAR8R3t5Ci2qPKlZTh56thP90v1J2Y
maUQx63Bv2+iVpmggoW+Em/AJUh2QAaal1gK+8DPbtA7FGGcPNDB8s1qewm9wFIC
NRoJn1tmXo9ibpN6SE1bTPeSaxTbuRGa2xTGXwQ2Ya4y1OicbCCRX3c7sijMAdsu
+NY1NwmNTwXrkjaJq3AVq0wzhJLS64XmqC3+efCZvHQWY976Y+8Xr2K4XLYtm9SP
9eN1ijpljjjbWh2zopy1/BxPCiyiYpzT8+9x0+vJOeskoSAAqwDAndrr1q4Qrig3
vd4Pg8nO4OxYnFsMHOI/B8LwFD1NQjfMsA2zpkmfsZt7Rg9I3V3dIjU8Ds7BXHsh
gm02f0a06XDB36W0N6snmSGYWfI+mMnjXVvuQns35aZJnKvoVFAI/K+usl9vwLNx
kfINM6nXvEk5nByPihRWD63fZuAPtB+EUPag2CapqhevUQX/VZSFE+03lQN43jrR
VWFgND8ilBBhr8FN7xEnHVzwmwydXxNOtCyG86enc5G/5bWTU1fA3JttylzXdipV
OS+NQWe41q/JgfBJ7gXy3LNmd0j/oqQgZdC2HLnYhmKgAROO+gjLIVQIJvQ68Fq+
2jac7gRdXpXuHQk7yEQiatetiLJMaRAdL4D9qdeAlk2oJAWI9UOYtgnq2XhPklf7
vR8/8lcICB4o7+XQk/GiyaQf+yLoJaEkZdzXVPOpGLiXLL3czMeg2uzT1ZCcBMmL
1gIfLNhjf+CeDDVq7PVsyOVRo1AlgL+p7uXP4KARAh6iVm8JQAeBiUS6x2mS5rd+
1J1aX2N/YsxRPUOkG7hYN/qJideAr7VcUnRCPW7/BKnZ/ZhWmCoK4gpYtEW5MjBq
X9ebbQA3O7mYv4KgtwSHpdEE356CAAFVNM16Bw94UOifec8nAjxO4Dyc57QYpTKr
RMbn+EuJym/fkFV09xE4yZfNeg58OY0mThVzXXqlErONWxuHFiVGgk6yu6LRDOI+
7nqgDE6Ai/LK9ZfbNZrtbQqDxCbsbi71Dr81oV66b/fldVn7Hx/g81iz2nG3H5Zv
1/YTfU9D4DmjgfhLwfBpzKfyApwlsi5OTpqnz/Bs9nTv8rCzDvzkxdz/bdHh1olk
5GTU1z5tpS7ey2BUjy8VvHjsCg8PaR5WyuOTcvoFCgteuHZBOjdSlM7nrPBmiAmm
aV2GGqoIUVc4N84jsnJHh0+U9Lu/Ifd8h25mS7ZBIMOYqdBedbdbHKBr1d2Wc2jJ
HykAFhDs+73vXIOLyZXtrJ+xIDupkJaREhiVQXZpL33TfpKddCbn3vzoTgY5lRPW
QDZgQt4CtQmwOxwsENPwW0F7w7Jd6/t/kuDS26ZZKc7XRi7TkH3oKPDKprxQQy1M
SgFvwaoK2Vq1VcvxGjK6ZJjm2AF7gJOJUGmqf9bePSobwx814an6PyIKdAvFhYUT
FAwwvlO5ZAJxhTbp+AU1399Mm3sBQYx9PS0mBpjk0GHkG5xNJa/x4VPMc5hkmb32
GPo6vRUargtn5R2B5wiVuX2YFH3iIdAIb4eHSAKQVPW6uWlOTUWEPjKS22pjzjb0
dVcKLOUSOBMzS13+BQtC2BRuNfv7T62WGhZtfGz/U+kn2hbkdcRZBz2aBwSvEybM
eLp5VBGe3pw52w1Nw86nEuPJwpd6DQMqTEUL5rCMj5kSiS3OQrYwtkRmG72SuWwu
xTjUv8bbbc0rjSSiFzXyrP1RfBzIMoTpleetyrFq5uiqJ60VU9A03VFNzzEqXCoS
ptpsNm8XxJKTH8gHEz0xBrnHwbxLVEV+1I24qkAztOWR43erWd7gP3s0p3kkAaOG
Xcw8OkokOED7tp8bfiUW2Wpfvuzi21Sdp6fBKyxpAru+d7jNp5HsP2tpr9hnocK1
uGZEjwDQNoELn1c4wycFR6MgEZbvbCMHfVlT9dPhJvOmHy3KBqXskeBQVcS8O6sd
P0lTykIOgkjInmguZBK94V9DQGj19zn3XQxKb4jfSEJ2I0oJt183ApT1Yj8DQViN
quvOBTpKKrXqoMADtQKzaLEZXmToKKwRFwRiBtbVKyFw7EwhTblYEoIzppQuN68A
wr7u//JP0uO8AxQKfKcWIKFUgJdHAVkk3GJhcNS+oo3pu36BA1CV7x8/XoCNAVNR
36AQPdu1IAtCqU7UvoGW4XpEzZtWJ6WcpqROHhc5/GTjjtzFV1PGCCUIh/3XTkh4
tF9vafJTnPuUDhfTOJE+PJA3uz8zYiwl+S8A+nEp+nAXPkfB6gIqp/MX8Ke8D4zp
H+ZMjzIgkj0G4gXMPKzUM8sddvh+Vi8zRxA2cuEUii0ruayiIQabg/tzmGXzW94O
vLpigel807pTaucfvyGyf2aspfg2NmfezaXBeXPfOqfvxjrZJCjTe3/4mtw8IYUS
tjq3lFXyaEUdjneOPApgh7yrpORDWj2vrs3vPiNcWVz2YPV9RFUifrnmIG0i8UhN
giEqsVq8qzeY0vF2YAxbcDqPAydWKgJ74auF7MetruOleHQyIeea8JZ1sOaH3Bpo
ZHOCeVeMAXEQFc/FwdNIt6F/6BvT/Hw+OFt7KTSZx5NngKj7lFaeJwiZBiOgQ6cj
VWeY8T90wSu/Gx+Pi9/Ln3SUCuTn6hwuVULs4ZGr8Xd0gd4shFOPVuVTfsA729GJ
14koVtiiMHWrPeSUtA+BHEnQqe47tIFTiKx1pO4C52KXQGZvQcaqtfKbyHWPC7up
SHtWUcNCn5zJcdG0GFbCgdBAose0Yr2APtYquZyQNsrs+4yHcdnQRUbE38ieEfla
CyA5DI6JHbTTDC5/LIjFt9Ph4XBf0E0Qv3y4oxlAB9emNaB8Ij2/pyZbn4x3XPck
dWvkMYgf1S1igoaXeqM970VxsZ60kFcGtS06saJuLTufUFv8FjepEwpxuz4D0taw
kLbp3eCUeFoQiQuQv8HmhsEVACXbrV1b+ekU+vDAunflKOKyBxHg3Kdjjx+hPKKR
TzBoL5W+mDgAj+FNfw77pBwrNHTyk1NhsQBe7g8H8XWeMn35qQ7wa2/ivXOhz4YP
Gf3M/I5WZRQ5jX97U8kwXUNYLVQ7j/vhbaGzmWa00nEY5fjDp9Bt7UgUxxFHSoS8
3Mc5DR3iFEkEsTaieY4cU7svWbc7j2r9pyraToi0lsCcGVgyo2SDtnRseyQ94no+
sRt06M/xSzb6LSu60m/lq+9i1Sz+/4lLkSsMsW6SOcWkHtVX5VJyCeQ0Gemqkwk9
EaiR2LYrY83alqCqSzSIZtBJY00HcGrJD2ea9XeNWWvER7fgDirypzbAiYh+/POO
q0eCvmmoUhKnhuM1Z39oXs24UmsH1h9DSvaiHMbUS2oBZKdxiPgGO+KQ7dY+2832
qPA1Mq4pNC9u7452JpS5+/ZhnxWRaPQ+VzVaVnH6tCYTFurVgF/KsuP2QMTtYZsI
JZBitJjf7IgESfp+xLNxxdmC1tc1VaXlmi7EpJd5VCPpEqHDAbmwhSsJBtx1DjNd
xov+ID6ga/uN5x5qY2zZZJvZKgOG/9cgSg9M5fgRUqmp7W9joWI5jO+NZRI4x0D4
Hbd3G4pfDzlEUeVxXGrpNAvXrlbCFPnJDOiBNPioSMgCaO/bZISy4dR/UknDp67g
Vqi7rCwXdVhHcXNwGuhueuE5L4wwL+6HgkMuiiPVXs3vwZsi7y+fQU0TBJ+TEfk0
z2pRlSfOSqfNG+eBynZewW8ldyXgzMcmKeFxasEjhfvSOVA59RIPnEKgb4jq2avh
hLyEngZBdPKPVHeQqOKwJFbiKInfychKl0qDOe9nXo4yR4qJMz4MdiOjfON9b9In
4jbCV/Kt75WYuUaGpg6GE0VGWpiiQdck9CEUYLDA89I3PONem/6s87A1WOBxgTVh
I1cEgbDXcPX/WxKyYeptoGvwK0K8Iu8Pv4zQgaF+0sFiIjpNvTXB5ScESLqT4yeD
DaxHEjsBMGO+qkp7om6hhiet0ZgbNHZHOU8NBi4rHFpZ6pSnMJXjvrp/XynTlkcB
Ush6QYCNIGtwHrl2K+ZC9NSaw9qYGFWTco9oFS/OTC0LYEg9TonBaUr1J1M/Cci0
qbtFFFYtJRA5t4jvADiF3IBw0ZoxRQasr+IWMJE4lBSmMkazytLyIjOrbNI0eWzw
3mtDSwC3entoHMt/0jd+HukKplFBmkUwikdPA98VrhVkFkIbMpd/OUeg7kgZb2qM
ghazZn1+1M+KVy1ccQNQq3md4HOwxzIE/1qUNoTzIXCvvvtcNF/tmEVfkuVCgiw2
Ay04wh4vwa/5istr+/4cGHebzqjSqZF3jn1/EbdHqulhUUhuVkGH4SihIXd/GlxJ
FBhP/KuvBsCJX1PjxSIl5uIVNIY3EKEaYoXUShOIyzhn0rnTmccopD8i7+Z0I2ls
20oXPxkcIq5GiEKORBekf/vQ3HJaM2sf/uv6pjQDVcl6x8w3NVi9pCIFAwYm88GI
/hinqEkYlBErL7FDMjv8UacTp3TZWBDyfrQBEV6DIsUhvBx2cG8h5+9gdl52X6/R
tv+qUdrKdJ6j7PCcdo7PCGWYpIPxTDHvrlBvDWrXXOJ+VWW6klafwC3cqrFK71L9
4083Mhp4qbU2EdJxod7Qecg42L2iBb6kf8MIRJny08h1fbOwa0F3uNjzecGtLDtv
CfNB/Mk3TM/LSh8O1+p68hdOQii814Tx3nCzdayOL1KC0zZFO1QiZPB9aKaiX30p
1GeNLrBMovgQ2SoKHcBHurIGsMSZBIW4BwuzcIGsoy3qmSQ1/6Re7efJd0r+vAKV
WrgGxKm4/OYs51Pkjl8rtVUTgAwv/kD9ZSeLGBruIAijnIBQly26eBreBxNb4A1l
lHqZmJqx21kJeTh0fs3EMolpZ9PRSkk5zjR1DpkweFvbjPhBUb0Pd6jdt7mColMh
kzLafDaGHxiNH5h83anqJnj1JKsEvx4v5DF3Y81FdjFRXoU0GUS10UEdhNBfkqMW
bEaW4dvUicTRhLfZduX+B6Fd2kUfOx2NsvwD+Lhr2XBPCyLNCPhHvEVU0PDO22Jk
/x7JYs8hjErD5Tt28VhRc/eMfiIwCNriNRlaKUbgf1Zh3qWT/Taxl8y+5RIGyF+N
RWFWOEjdKE8aWYucqkv3ZZ+muzoKbjGa7jkC1WGZSaxJUDTqTBJTxatRtqTLIWkH
SnbFh/FGWgFcJxH3bIDyH9CEnFwb/PQFlJX4a6oM93B12JagWvF2zPzoP1JjvN1W
dbSp4QPC5rFumRsv9qAXWsEr+W1dBex78QpD6iOO26fTHi/LFhIeJ1huQBYs3Wsv
W6D9Tdlgpst/7vgYRZfb2NXAq6kENIpfLKNoce+K10vTAWqknIvETuSu/kuXTnz1
KCnRcJcn5CTrp25f2WSA/1SfapHspdTvbrAp+TlIAfBRsohVpDXSZjvn+LO4ENK7
6TsMkkkRWArDjKCpZRg0XgPTnBCqc+KmcaeayHaX5SbMfE47akJp9goksRB6DVvq
ZYbT1PQKWiqESwAlso2b0c7Rq5ZWhv6Uh5A8AkG5/NTQYCcg3o8YiIptsb0y3XUU
oPkDmNKGqwFAVAh/LiDqw7lkrrqjHUPFPT7p66K5cJS6LFdoN7fGo2xKw/cSTINd
KQ5dyiHrlm646kjqgCanffsT3+CQRsgG3BVl8c3bBbRdU9x8RJb1Sg0qZGrgqSjN
oCgJ5gVWF1n0FXFcR1oqru2Qa8SBskC4mMqw8/rAS3NYW4JdBFkorm0vzl7JWZrZ
un7lEPrcRyFKQaG2puU4fGX9WtNHxUXW7a2XwD4Il4t8uFj6c0bwvIMa/x4Rp3IS
GjH/AoSH+xqBQPGSNeb/7XBNkVJI9pNJkI4WZG3YSFiszRbiKsV06uuYvPJQx8m2
kq0wqxtinLuw9IOLtfxYYGBt/HLnfe14g2r6ywAO22qo5wzWMhKxvtBVOG1422zU
LJNQqYGkmsMDN3Vb2zXPXNCpoGezksfvlxa0vH6ueHRzs8mhzJaEwPmwcyLIMa2Z
RBJoEMe0obFXK3TyzLMJW46tRZVmGNXhoLo6npu4dWN3PutHJ64mS0U0bY/S2Gjh
mopZdTVXs6DCat1nkiL7nVH5H36TKH/8zUrMcXAo8TIDJccd+2RNvk8rJd+HD4l6
vCXG+EB7P17hUGitpoxLSNDJy8Sq9fIar4rGPxmhS8pf1uKqyqftI/lW2ilolsEQ
F6xmJzHzBrsMiMxMolpO1484uwD4WSCvy5kAc2DNYoqbJXjXscmz2IWdqhjvWYEc
DdSQWIRgyyAEh6UE/cKDSOjYauXi9tO/0yUzhomM8Ls1sgPl1SCBGVTmH8gF1RAl
0I0F/4COVjP5+TUh6t1Q7xnWLV5oq5pDd7l7U6GmNNDwL1QIwmk8sHq8KvKX9w/W
JdHzzpuvbA+69D9K6aOr+ecxZk4SNSeqDNW5m34BTWRyfdKwdD6Y4iMAJdTkmsJj
659g+TglZFCEA+Zf1gj1cbw1j5yKoe5B6KsuXonTsO0cUjKigdFRtlNsS1Y/qvl2
mCwgE1oER9xIAQrCMPDb0ShFY8hernLuk8Ms2JdEooQgHZQiB44AuYUScV2v4NIP
Xz0WMlTODM4A3RBIJieJwzrwvUDkPuP8dIH9q6QrGJWwsYtgV9+iafLXd9ijSRXf
oJsV8Hfp4lkwMhJlraZU8Y89AkIEw0EeDoHLBH1er+BvKY1bAT6FaMVB0YxD0lMC
13ZE2vGxVBqULcPfafuQz2G+GyOLZB0f0Tyyg2waGXVogOOusKHfQAuPjbMo5pWu
kyuv5pVFNX8YLFnOJ6JRMHFGobY5Jg3+KV3L2hAGQBXgKSVIcIQskNazBy3zhGPc
1HItCyzFPB9oC/VegLc68eiqHHZ5Gq+HaY8YOLf8D/Z20YXLNYfj62vy2hEvtSzn
BRIzXKzelBb/o3Atm+NIan/Z4qgqywyMevEIxd//k6hXEehHPNwpqSzvjY+KJvYA
73BJnpiqnydP0DtFnaGO8gGoedSVCtpEoj3EOxyqyzC3W7CpKpy2DxdfCkD9Jf8s
gqV8hiFRwcMV3+gAWLIaAEwQjS0+y7ityoq1nQ5hv6EwQON4/UMVs+d7htAGltrx
QAjQNrx40nX0dA8Z17ZKKt8Kt+7HCZxR5yhJX2BIbdqjVHZ2Yz6rczlsP3deQW+q
Ni02EqeI9d/LS5P2gh0XloQf0X1BXn588h2AF2GIV66S9Ti9jU2tkI/5PDrFVml4
cozqOErOHgUDABH36pNed6R32yygJ8I7/xayd19oq9hwldNrS+r2322IwDKBZSqF
5sG5hYlhzIOKwiuIqSjDJQylOJA2aaPYyqfdBVItLzPtVgNaL4HqViOrXtzFlcSe
/uCHX6IRWG7ziVuhF+c6vO0xj6WYNWLiFXoXxO1JRxACK5IGTMPhaH/p0dWpbYnZ
8Bt+yWDi9SUVx3tNDX7PP4XoyHaXBQnT9kvQtUEsu/qyeJLW1WH5/BnQdA9JkFoB
NR2raAsmAd9JmYrJEzJA45i69hDeO1SxDRBWildhQPJpif7jA+NkaRoCkihUBQ4S
S+6AQMrgBCxgVV66glhNc0vKbOAoudW3bQb6szznREkenH1uGRcabiWyq7cpuQA+
NOoWGNSs4/SUydXYM0G3l74YYNjdPChNY0Go1/sHbgoX17WVny+hCSbspi6ORhba
qGtLGehszTssZQD5qgH6urIiOv/rWIlf294NDMU2Eqa9YcMfFSV/N7NXMIh+Eeuk
YqvbspTsku3eaeuV8zxN/s6MD41FiPlkWUXQHgH6fjF8AVbVU87Tqch5nt5g2mTN
UMRvkz0tAW4itPOGbXjbkaD9EMTwfe/yRC+QwGp5rXZfMc3iJMVi0f27vnN8Xcbz
LLUtIaUGbP0a6kFZ3iEIo9QqwS3ve4HB3qjYuGF+H4h5n37Z2Kp30yiWwtCglP6Q
KddcUu/aVrIlApo0YkmIE5DirRg2hprd43PmVxNVajy4noq4MDAB+CZoA8h0QDP1
y3EmHPK0ekxd+D4YvQVyPiZSDxTHN+C9WIA3EwHPTxcGFG00ebbj21BgZOOMO4S4
8N9LjpySJ7LvBfgx71Pu3BpCbIEU0MEROBshUu+gPxErZqHArikKWLevo4dY/Gzk
VVVbCvPtIDjf4MlUBz+8OUroaJa9DXgUqcaW1fPWcfsaov3IzeYy4Flt/pnM5BeG
QuxOofBEBcxI/+4SHVq9nVYzh/Sc9iy/dtDyQNE+KRx+P3GRLSYHxDvYjxER7ovX
zYiI69du9QakeMU7dQ6gWOLJPlEiagZuPbGcfJ1fztZGv9qOnlA2RoEDh2X3enMZ
tY5CYHDAOkdtjdFunlfBlpi+DH3KdJb8u12xN4FApIbFWyAigTSqLK+/7S4qBBWX
p4nLg0JHCYbfcG9KAlSF8d1Z/YC+dRsY0mNjVtW565UajVZiYnr2B+EPm6cJ3WDE
7y9sEKgRKif9eclFIzWdGkbbUzDV0N+9B7L91dmfDccnsUD+cUGC/ooN2loTl4zk
vnX/ih6QOmnO0SKSy6PNQJysJo+ujVRgsJR8HQczy3E5UsNe/NW1iTbQoz2JXa7j
OVzHRxA/MSdi/106o1Kx4+CM1gLAyn58xOaAW/uyz8OHTtUTu7gjea7s1HKRphPG
Jln4H/HFQhajUZBa9kL1m63swzUXz1XyjSdkTQYugBzGfVVYcWwMjZ1INWcTW6E6
MKfBpGIpzgiZVUjHCvGSIDyStmViH4Nx12UZeLHuwuTVaSdf4Z+94Om/VirA0xhL
AcYsoDcfSi1Buns1OzRvYzKxWQoVLyJkYuRAJNqvM43Q6EziKrfoqJPlKv762nxD
3iUGzA/xi7KzpCv8bIvsGfnFUrcjKRR4ifQRBsImadG2wDsH9qOnEsPuUDqlpfEa
rtSqZscw0cKAlD7iY5joH7WnqqE4SjNtaa6zhMYL9fPXYkDR3xpRTdqX55OKon6g
1lLxbsitolHzKTwy0o5GOsi3ipKPPxoTWrgvT3P9ssHVaxf1MzwBvtM7N40HajZL
gaXuio4qkCySIGUVhpnmpVo3UUMq3ZA1Arsk1RbywDA3nX27/nRDQBEaRIwa7ICf
gEUsJud1caMrqlZpJtT4G3BXdlYpg7FV4EJDGvtsRxXkHGq4boK6T4O0yZLRsztD
xga/3OIvYVC2H67h78/xgaUKKi6JAGmkGtoQTJz4LCsHLdu9MHbP3zyx4prftO/s
wSb4vZbJeFyGcs/DtlQ21JlOYcHDacxBcCuq6hs9h5+RZwGDzGYGtDEiEN8bSqUO
bbqbXAK8EPiMKVyFjaTgzS7KwxPzTvG9lQQDAkyY/IiitGMubDrjokSBZllRNHq9
bPMjD8zKgHCzDwsZ+oS36UQW8NZhzYikskP92wudD6jd7gkZOn0s6qdBQVSdFcpM
dkzPMPpVs8+FzaX95ulL3qFUYS4VfFK32BZ2c15gc1ITcJnJEIOuIxrnHIs6xcRU
GOJ9RwEkqrVKL3ghMuHHJyiFADt49htBqaUdiucC9jRctcrvRW7DnmoeNTQbkcyM
VTAofGIw2VqH5oScislgPK5aXlH6UKUNxUyeRJZeAmdK0wm9RlaDarjcRuYgZ9YY
5I8/hn/w2RfE6XhwG2a6imag5zxGS0Lyi5tmrBoPR445F2AdMRFSIwBg6WCgsSHs
v73xN8ILwdx3JQHvo2s2mU94I2Hngj4O1Hno1/fd+iFMB7AB2GBll1nOqPtVFwJw
o+bZE0cXrYNBd/eGNz6Ky2cDh5sJGmXeCH7M8Oe0p/bTk6MRMLoq17yuc/Io5Kv6
qPQCsLE3j2BMUCNCsqqBSgbJtygW6uIPeULYDdPcvoLPf5wUn8a7RI/EOVdUgj7U
JnI23aITQAm7Le2LMn+pLS1IVlKI2id4f9GjyOsi8a2vumYHSGCFFD95E1MnESaB
X3UhSrmW/zxtJ3mNeJ6NDM3HHs+GEqjDTy7c6AXwEV9sCrqKYCJjCAyCOQrDpGAY
uuaqOaXNDUrciKv0VT/Yrdsu9Wuw//nrphQMx0eJqEb9Mvc8YTpo0eXYmop+4ObS
tf0zf/pTD8nNA9FJ7ZL74VTu4+aB7Hh2U+8pp6M37MXuIv4UtWHAXghvwWRDHNxu
bhl3tXokgkXRQhKu/WQTdOuKxKH3IgZAmwPrVXVauQdMXli5duM5DVpwqjSO13U5
4w2odSzkhy7Qc90R85wMXTdUYBLoJ/NJFUA7zr8k8hWdGv0856zReTjI3oK4TpLP
AYWUWsrMPwRkx1fLKFRJIocjm8CDJr2bg8X3qAaK/dd/YxIq2VvzYXExokLl1fCt
Mo5ybMolfAAg2Wejfdo+Gg+bBOYMAaiNQjDP187vGR66BbU9fvA8cAH3fxwMuwzS
aRp3EZZCKgYJDu9qCzDm/GBZR+DnT2aJp383BkfMul8mk/blhJIU9pESOr5fFtOE
EAkyv/+M2x8o0qi7q0VLTqhP6INR+R1ViffNk9GPJt2oSz06kviUvmTyRfs7Xw99
D9ahRmS4jIp7pzDxtcr8gUDr8bJAYSIbJJI5bDWak7a7/VbNliqPOgeScB70Qi72
dB5UZ71UjkXZh+MQoSV8gp/YkAkmM76jAWW8TMQxosf27I51Quv/Ytge79eIBtfS
HVRGLRKOHh4O3YMYAokYxFFmYuxddDDFEiRWS7nAftClbdjiiHcFTu1944DQgmaL
i4CMJ1P7R5bArEUnhoeDn6a++IN5CP0uZZzluExRs4ekOjcsiH74M/FCn7MEBj2S
uGCcoo3xZCsLttR06wStrvVXQLZkYGutV54Su07dGakSDqDcp3adPwmi7A84dvgV
7Y3+9vSm8wI4flHq5JuHaFjMqO0EV5XYdno7PevWo+uvUFR93Nok98PsYn2Gx8dD
wQcNHGe4cDKhJkKvdAmYO9/2qUizK7fI0D16zsvPbnja8L0dc+4cqs1AF/YAomQy
6nZiAHfhGtVji8/yeMDgEsnnJCtNk8sVUtBg+9IbROhwIDgO0HbRcvGDYRtS98Pn
K5vSTk31wKo7n/oB5zLQlBQZrTeJctnM4RAU0JJrQGN2YWVAdw1TqNMcpInpL4Mk
WL4096aF0BHKvVB1CsdfcjLs3QWuaRsQv/czf1uZpeGCBJINlO7z5SUkGSwgR3Cy
8ZZOtBOLiM4l2LYR1obYASHUSh8dfkdK0SLsMFy5IjZHUDqdO5BvaY7J8PeiVywi
x9vrOHv8e+JfUPzqnlRKqcHtxdk9/lFBeiJ89bL37Syfk9/nBwjIRRrIS7v2+fyU
aQGWdHfiqClKM/uvWAcFsxwU8LnXBPXuaDuP0mxUai0Iyf2Y26fMgTQdFdziKFWU
ZVj2JmSNMkJrPjL1XSMM4EaTE7+39QIDQ6GuSrv8+3WhAGIQXDSo9UQzQS2aJVeG
wVgk1vArYTU+YzQwj+8YDgDf2tzgOE+DtAw7LjSfrrPiw/R+kBnamiZTXmLljaq2
DoaqXHfD99eU39JdzilQBjkx+KPGJtFsqH1GATuw01rK6FFKWYAY+AlBZhsy6P24
R+upkQEXpzARINKkVi7haBNEmjjR6UjBt5nPBVO9VtuxLLhFyPE0EOLsc/9TJVc/
UPhfDb9T2UU7+mCqMPSmO0VTevGB2NxkU/072y3doY1udhxvmohPbNcxtIrdqSsd
zyLyN+bcVq+Nc93jApJTM8WCgdrVFxaT+jSFYwdbCX7fGUCNZTvBom5IXlY634CY
yJ3SGkzSdta6oo8I7plzcvQf5KZ9xVjHuyVT71NBGAihQdhi8fi9tU7r+Ft6Hv4y
B9PBYzF6+aOnwkmznqqnrmogiA7UsUQ4LKYwr15XQiSlfD3jUaKsa6IHq6LfIjc2
nQ811MgRH0bHsCSxExSytz+hz6iJoAWyXArc4aDiDC+0TlZgN+vxEV5AwKYdWnyC
cPHDu6yOaub2+eHILp41YsVGhH2g5U9yJUyxJd9zeolcteqMlJbodmSj71B1XySt
KXXQD4JTmKsgqepCmGeCju+Y7IzaljsrdQy2wMJHjr14edblbJL+hXV9U/rjGjiQ
GpFDmKcF6Ew9L8g3IL7/mmBozeFlDvjwSHnqiN8uhEYFzg3xTmQ0vI/dd8yPGnK6
whDnwhuiipvLJK7ugsfVJT0mA/KYQgVlw9lEsSCP9jaPGMM/jLqRqgiujdDeOwJz
ppht+2Z0wbyO8yTeR+LEfOqhheBwhGnySVhAFBo4X+INw3CZsh3JUEHGgpGsIca4
DSUFDOPRbfyvJ5CiCYUCaQhvmC7eXOYPq322phdkCWJdWVMfWYvFe4REbxrzYNgQ
X3hbhCsDWNsWCcU1FgfqozLXfDuokwJzTb/2McbEKfyLxd4dkButo+n+iaYdFlLu
Xjh3LHCewTMTk5/vC2sSgeuciyuSQRx2+TVPz4Ir9vCzXmfxuWNK/M9yQZ3n3isx
LOU22D7B+l4xACHph0oPeWEXkt/i4JCWfpSPrfvSgtjchyXzdnfVb6p+Mg+py0V6
0vXcQPoqSXNdkkT4rHmVKjGiIr+ziNkgOqfxN+5hZqjyPbGdWtofVhbKpBpTKXj/
yWYFz3lb+cHHOMzZ4cp+JItYZWauq4vT/DFeL3HuxZQSoCIi/Lk8rTesrIm6uB14
EjmprKstmn9Xq0XrsOgbFKRMPW2Ay5Y5nf+dpxhBvOFZ09lWmmVKwzI7pCQ0iHLT
9aU1mKh2BiaO8VlNjwrbx1Mai7aWuGnHcE92a/2NT4LxyFZKuPb0VGmOByN1ai3U
eJMG1eacsvf6PqotQJubF6mdZFylS1EqZurdEk3JCt94WlJIFBiH3c3gHE0UO9Ap
K3cr62yIgwTQnQoGwjXAKSKGqAWMBD/wYuOUaEKMWfw7Gmvkymvno5pfa1rJd7TT
3J77M5UcXdHW2WrYAPtK9D7R4LgbyX3ZoikOugD0E1jU7m4iuhLdMVMHY7UV8XZb
oYzMDHX4sukHSTYEs2clGbkfRhacElfxOput9l9Vqa5yAUQrOdpYB21kfkbYKjvQ
Uoxlu963lQvB06zHeTkk/gggb10spT9CmYZnGFlAhd+Tt3kUcUm5kT2gvGCBWcrO
zL/J5bv05+sWcnhG2yJtbUF8WXcIBKXm4quTjFI96ABy9O+tiCCsgyfmRuH45EMP
IzZ8Y/YJiKLObDNpP6DMY3infwst7+4D9eC8fw/DFk1+f/pK0GkauGy/fUKGBv7g
evVGlXx00rQkRHXc2ji0S3EKTqD3AYmlBy/CmUsGxE6Koj/8OQXTxfQ+xucriB+b
Fy3NCGDa+ewHDAGi44hb8Gv2dSak55X+yv7qHuWV9Tzsxp0KlFPFn+XoSyAB0G3P
A5ih4zz1yRPON4RN0OehxWRNE13oNhxPBh+fRo12i2imjNRECG5eflPqf6xqStgw
gOgUSfLjwp/QNSMmxGGxl7BNNExMd/dWPu/UOR7UAK2JWgNbRk3YNmYmQpFWmmyK
bpW+T6qSGOp2HAs4UZZif7JcTm+TNxRUGA8kO0V+XvFMntsyCR2IBYxqiH4J4Dcb
NaUohv5xFuxRS0a0uklteHrBe0v/ioOUDDOJSW/0YdmSKtlg8l43G2bIAFSXOBel
0qrEjblJfY5+Yls3ukebzMAZDBcFNJq6+bIQDIoGzJUNm2p0Njzprs0OoQ1eryEf
dvJABC4mQ5/l9JHuMJYIu4GhPtbO+vFfrbQTWsl7XR/PwAY1rO/POICy+Bb5Pkr7
0eyrD1iEMPl2UiU3iGMdVMze73Jo5CZ1lDf9nwa0Z3YIoTm2M9oxqqBV0F9b9Nis
KJCANoJqDs1gmaCG0H26yE7C2ChwcFk6DBzcjpcKsnsasbgTeniRWqGfOeS1veXP
9D4vO9ZCTjPeHcfgrY60om6lmYGJjaS3wHTDm2LEL5ojawF/Zs0lGkZ+IBamFOss
0pSRhRmsEL0OUTXhyvxbxmwUvRDEAq6zbKCWWCCCHr24rETZQIQTnFjklkKqHE4A
Irl5eJK3+dA/5fVcmhkpGIJIcuHZRXKWkA9UhwbpZIFaScaMjZjzKF4PA64CQMcu
S87Om3K6WdqHNtYdCdRctnNkqVjJ20LmWEdts9uI2t6IfcIB6JF/tdlvGCL9bo0j
YfRmwYs1k5vT72TtzjVLV9YN/E8VgcyXTb4ZEnSyAkizO+ByJ/vx8SLam9wY/PZi
JqoIvAHKfnMhRDDvsPX5LSCtL611fZv3oqOk+KS+cyKvezXO1rcXCHM8J6NwSALC
gUOcTXl7abEf7Rl+WTPcWqzMbTzsqiIIVli4in3+dS7Wf/o1NI/aFUTfdn9DrWuV
b82Jd/ditvCuzNc6vT7hnm5TPOm98Kx0tFPBj65bggxrLgsMlW5I114pNKLtMiKF
26Q/fDwGO+KXvrj0Ly75IARTu+0pFiWpcxpehQzcVn0IhnpwJCTjjJ/xnfK9yGiD
OD722GeSEmZ4rBPqNHM18kOlFZ+NR9UqPxycwsWE1QGokUURE2XuY9/F4leHqCbR
+E0Z3Gv6usi9sUXrAW+0T8IZHzG4V+pwDE/tpHkwr5X9P8CTKRLZ55u3uKoMl6ab
LkKGppLQNx6jKEIt4u6BC7ooGMC9woIJa3K7ZMuldLOJhbYb1XHWXY0WwB9rKK0W
6aunq3lH50Tj43oCbouVRQy+6Kz+YjeJ13VlerR3UuCEvl4oYm1eVlnl+4zP34Bo
em2yH+nV0JozkUQV80/o0DOI4cvIHDeUYL95Juh7B4rfqPQITSB+L8qI3pkqUpXZ
mUhZ8ugiYWix1ppJUQAJeolOTFaC+OD/5usgOb0aCQCmk3850+bu/qcQAhQxxZAi
LLhDwLm9Ke2oZhTHNUXsvM6lNMpxNI4qexP7UWyQrRMpdqfpUjPN19FwdPCEor0v
QMw8mb7hfXpteNy75b4AgETaMnKeNwb24w7QUwjrGv0nYDbjNX40lFLZworK+Q1z
NqBDN8l2KyC3Ta1/1nl9/FaC4s2Cg9IVhHPtmOyG8H8oMJRcHvJRFaRVqPYBkeva
+ZOILFV6QQS4d2Sahb6HG21OhGqdvJyZWifYKI186peeWEfxqRIu4mxGCF6Vvvka
fYmFIo3K3J2Q5N0IEW8TmECMmqABAT1scVABOjHs4WhrT8Rw4d8Y+pyCsaoE4uIT
z0J1yNXNJbna30hSPSJG0L+SRANy0vYBQFyT4oiH5t7CsPrh35YvdpfEBXW+j/37
U+reQblFcue0KRrw4m3FAJ0bRtZAFnqVSxo7q4fXYldmZPSqK0U6UBQG+cSpn+YI
Ak/15KjVAOGljwukcxVFmkVSvqvKIew0WcJfDVjIT7Pl8EWIit6D9zkfZcku6kCu
SnJcIWbQWjQhAcT28Zppc7WCXgw9jgCYW9T47xJS6FHBzGGDfmjeMbFnomT5AfNl
pGfHK3bQIpnjntRlQhjv+oF5jHJWBgXZbnENhzJ8pAVGcUuG6R2JOljeB5xLXeDm
PaJkqHKg0ITg+R7EWk9jb+9HXBI1n8qeKRlQSDkKUUbIWtQO3SBkZOE1pSlhFkOS
z13CxmaxOE1HVbW9RzmZqclxgGs19BTZn1tVh2fJI8v4QoaY97xBrejjki8dJMnu
9AbehDowfiN4Vk1z4HotRQsoZjHywu2dAYAIJ4fHtI6HaYMxLheySpgOFkgjc6v9
yrnR7HZLpKcuh3ygyRO1L5s9lmYPFTSbbzI5pQYEJ0Qzvld+DdfaTNDvdvlgHoIk
KSXa9WI40qdzLUs7RMk5OsGapeOrEYCiRy06f43Gy+lB21XqmIhiax/UTFfswMSm
M0yQR1FJ9422DcT2czPaH1X04RfGfTe5Jfi6nJArWCMNoF7InuKVK8P1IdiUMUGx
ijPJUoIBX3q+60juRjTlnBxwaB/OCpKeJA3goGOQETvXueRQB/Wtyqq5+IIrs17E
hikcwhC42PPnbARBP9wKP2CGJEunZZaAu8YmF4DM8KA3/F8JyE+b3pAiOAfJDzFo
CesS9Rsrpk6T1tD8eL2QjY6RBgZMNJBxUi/r2nh8p+GwkR2ea0j8ljTCcF8FvpCC
v7bdeanCXjgVwWnXaFb1zN+EUraqmOdmAulPv2Wl7P/ei4QH0RsP22d0gcsvZmGc
RZy8si8VYlur2988wYIV7PHQzJLeTnGR2OealTNLgnksx/BrDX80Y3RR+d4t2UuJ
yF9L1oPFPV47dvHCPAc+ZMTxKjQId9fltfrniQtpKyQGHJe9DdNEzzZ5QrivsAJi
0fFDUffL83iHnOszd2TVutAcXDv766QjHwhcfRCC8aLd278fNf6xnS1FuOI0MKv5
crwEnYj5tRlQr8ETuLlin7lNa9VuXBtkJQv15tV8lEhDP02a5jKHNNsEV6EW7ekP
ymcIIlgcjwxwvv/r5zLQ+mn5aS65MpuNfwbaUkU2hE0aVbBqV3ldHZRab8fQN+bK
ZbOZD+pFf0AcRW9ZI82g5NIr95wVf/HvrRwMPy78/xVMSM8SCL2VQe2eCTGyd4Gz
ZMHxwwWwUz9EasJunczlYGHh77VmpfJzviU8WhjujBlf/EdhVfRQIaGR725AjBtK
bjNCz+HnqIv1S6i8RYVqyZ8/RPeKkElY5trU5aUgbH2FVImqrm88etyQjNHVMr3e
HWrAK1uu61LVMtbUYTptZQF5zvej4mNg8pcVL7S8Pa09SsaUBi8lmU6YuUiLs7hv
YIOnrrZykjzZtqr/6p5pEQnEuJ3At1oPb3gUSf3+d5eKTbaysPZfPiuVhybwaUs/
uVu4XOCG17RiqWavt+Bh8N8DkzEPB5cIx3GC66XoTJtydFMReD3we11d/QvnXe91
hMpvYfIS4ejINkPrdOE20rsD78fjxEr12wfd3OUQ4dsxQYHp/vPE5k1relzP+8n2
bXDMwRpRBQfTF1wgo5XvjdRhW/HD8PWjakzNiDOUML4f3qLfC6qzKEknc1MaIKOB
d16M+/s0sozhN0cEMyUL7wvtCvOT8wz8GiBhA6alWJZxSshc0ZWx90JqU5bDQqIo
Skc8phIOdC8i/VUw+K5to/Ew3FwaqH5vbyCLEqdIsuOjXVOzJPqouMBcnwjJbgzq
tFkLjgQreBcQ/at+cEinN09274m3c6OipkKyJCcgPNMImxaySvyR7W6TWEZEvfcR
/Ei8HRg4bIv9AL8oxO/FkJktEeYGRmPiwfeF2WAnWI6idtZQaSOrilqKYjyRzOZU
VCPxKbC6JnGLFZStXBT5nNJxfzdtLjBZ2p5nVxSBbhQ59wQ1LiXvT+LaiVrDrgk2
54vvNbyNVswBR5haloQShBztnjYgqRYsvFK7QWcI89yetrffT1je4N2uyrYNYZwG
rIVEJnG4P91xmqR4n13D8vcaMtH4qLStA/htJSwtkp5BFvLd/shSNrXHmRFT6hjd
QzDpI7SkD32Z46BY6Vv/FzpeaKjz7sinbvrjVLKdk42TAOd8OG9yP6pwwJBjd1Sv
v+s/Vib6pNqt/OObm/p7eAAsrJYWzrybcxQc/L5AUsdiyafnavNswh2ezjBONtxj
E74Lh14C6f8FyUCN8q10DpvEhQCizxvor8HrQs8hIyIQB95FIOEqYHjupxNlJKMN
1f0JEm15ep//ZLSpGX+H6BhjWue/KCl1Ub50bgbSwlzgqabiVGVohlaIogQHWXOD
5vVrIXp3An1JErExziPArdEpr7uNgZLAc5EmYc3tSG7/GBNBLMTG4TK6nDfgLVDJ
5sFmbuPY6PXVothCX0jBzBTyAD+xHYSmtZ15BNNgU6vE8gEIRGxwDTddva9iJOwO
8TNBJ3iZ/iB0Xz9ZwueSkiEhKi0HOyTFlXjvcZMJa9F7/ie8nkx8z7dFzC31wGOx
9a3C8T+5UXr8qqcUKTrs/5q2rr1VgrdBKWrGT9gWgz0hwSv+mcJJMGPxAOShkPS9
xOGmLCH7WnrZDy+Ctp4Yqajds0S11myLgjH7v6dD6DO+jchZ6ufl/fZhLs14dPnk
0jNG3ylMcU/jJt44E6tb1415kGxBexxL//Ywbd0VXmjvCoGJtQL4q2QYMrD24OzR
A9zt3WKDnBxfahYHDz7UmC3HlOlYM91MKh+kQi78/KEcN0YCXbuq9a4QkFTUYLvD
AD9ztGgfFqShT4tDtec7kj6LkV+LIb6H7Q1XFGhGAaY16jEe0i6GmsVk5/9OOtb7
R4cNSJ02pCIuz8MVY5L5gWh0CkJgIf5zk2kbzwG+Qy5ACCsJ+UCThIeww6/xTUHa
ifH0Kmu+C6GActBQ3rWuAQRlotFeOL5XmlyEmY3f13qs5PqaKxVhy4XrRfdIiXZZ
B3D7i3esP7p8d9KPMo1QlDW0GTz+pbdvmNACfohPu67XJdSE51aOVLBNvIuIe6PL
O004TswuEVwb05i7J+OHylkMRaA11W7o97mxfmOmxDCOi2ZnQmDMsdIRTO54r78k
uIgaZ5gw2Z99YO6mNNzVJT1trulRanSNapFgOA12zHbL+LiuNHNkeVIVWpI2e2sx
Dffz+6GosF0mOD4QF0P/tPfvc28MBm7iI1/Er0H7SFAvfGMz+k1jWtR4bR/MtQRa
xKsjjpeT5mUUm8vivMuMP+tJ2XADvCH+DbUibGBeh2gQKGDpQrVDjARGR9MrIlra
P2sq01bCuekqug/oOwmEhsFQUqpB4MeGWs6Hy9blgo/3+pOY/bt0AtHlGZ65h3Xi
waA4/hv/mmkqai1X8DjLZKRJdobO0V1UKhCQvToVUzHYcHVJZYCuorxjSJsGraPN
cMro17NwSL/OZ6dQNUTmjd8T6ljk5jxRark0y6zu3NIbX0vBxW5wAVf82GDS+wmi
rciQtAjAyfVCUD4ZEh1YAcDxq8W8ME0CaWaPHqR2IMks3lrKgufAp2iXErmSGggO
ZVjmxNTQo82r378XM3FdURT8Wgs9A2ROrptA6ND7h2z3jlEco25Xjh8xywjNaqwz
dU73qhVA3eP9wWaLOIlZVDLbtJaMb+S5oOmNd4Oi11PTGK2u13IRyhgzq+Vl4tcI
5M6Ad7kD81nLgEYwncNLiwjJwl5oCmjs0MZ/1BC0zk22xMCgwZMIRQeJXaVjACB+
+/3i+GeBkAS5nzm/mOpNcgLgahCKW8wmmHsgXNKqvXjwBIpZcZM/tptQyDD+r3Rj
iPNQK7w7B6iq8XY+0+YCr25Ct4+ze7guH0vLuMkm5Bkh9nr3KJTfFiDuV/jHosLH
yYIAbqUH1Ml08yjKavIeHOWHzGzpGBHMFF8sxC16AY6VtfyglF7+gbr61/8fxs8e
4o1LHEI8zZrpBTNMNJMBoxQj7IZMeQM4Ya7urosZUnGbCI2nXS0gdbx5h9Ryv+rB
Kg2nh2fXseOByW0rFVe4+zlAuPYbS2iye219EzwjyDpSMtSb2TD8ILKX5S5HDkA2
VeYYd76KaRJ9pVXl2uw/O5EjhvclMnySopucH+qvbzfH3xJd4FvYUEtQ5Ofd3o9u
2MSPgTQ9sYn1rc5e1gI/iXN0fmqNnpETg0Rf/jc7Kd+WED9B4gXzu7PsWJNYF8Sr
o6Cge3kr+GZenOgePJ5tv6mq0svCaxaVRYa4e7dCYZMbFBN9RiQGv69GUaaqvf5W
Jc9fzpLWrgqaaGk0tCZ4ftx7Pj72YtTBwwRIBLF74cWK5YwTmayTloXuNufkbQIh
mDe8rL7Ug+lIn9lCfsQmltNP9NFq5acGsb35AI5JwfFu6gXF+x8HphYZemXWedD5
VBWIIOvXaT0s5UaYRT+FgKvpxJDPtDZHZ4qe9J5EzRqFdGTn1M1uXnWSdGSYVT32
5rmMugTDaMJo4Cb172ONV17ZFMwmbDwSYv8ygmT3Gj6MWZFvSGKWvtlkwGzluwFT
kn24YTMWIIlWJhiIu0LTl5WpYRK1DFVTvtlCxWtFGuVeMSCU5fBPMtKQXYi8Ipqr
wCyvTbSXTGMynekmViQf+OTwNJvTchdPc4Yo4dK4eAHG7bhmuPxyt66kcqqIPsy4
5dyMbblLqLG/xZLuvxtZStUTl8TrBYtikgEBnJbjOEzOwL1LfABxP231bKpQXHEi
17Q1uq7euB2yX9ZfN5KmaDL2KmJcT0015SZo0eMY4OkqAIzyQfscZAzTOluiQ7Ml
urmlP0frh+oQaxV7v+P11LoN/SgRgZBrBRrxd9bcfFjNmFpuSI9gqO9H+RsLir24
JzzOqm/61vH6IYWu089E5/Rdqm5dXJOsFk9TRv/VBCikpcX4RHgP4nrFyJy/t+qi
O8Hr//HP9DetND6oSrVtukYQ9QftriqDNyz/zOoBwWywl7fAxaFmRvv+Dl+hGCug
4P6NWLD+uPyIy/xN6oLwO6IDVjWmfLi3xM5wx4UO9qJ/ixRtJGcOGbRV+y7SSaO1
vZthKPcEdQfFgt6iiC8TziqWmh7Vu4GRq9BmYWcTypS0mtMNqtgejasaGCywzIPD
STkIN0lg107FwXB+2N0OItNqp70FxC6F/Ap2fGB6V9L66dOI6c3Kkm5HBFGGF8q7
qnfhHSVqO4o8NXqiryo4eKsTOwu/fllqgu/HUT1wdx7tiNlr/Egyj36uiYCdDo/a
fU2Nv+KRJsCWwgu66IpNmMWJ6n9ynQMycScfZypBczdfyDYLw3CvuHZEy8F6gJDH
1rAX/tbJxP3vvp5gbjvXQMxr2mw84xcvR6plH8sl3eIrWRKqVN50xf4ZgmmuNFE/
vemEdusDKJHGtyms0/Y9YpAeRDKGkyjljy7ArRUxlL90RIrXsMwhoKHXvm7EDm8R
mldtY1++Pcs3Y3+QG+9I76m88MerxqPYuB14BCsf+rVJbc15A1gQRnTQewEaULrf
WfiJRvyylvgrCetMi9wooMZLHSmk3Ea67E5Cm6aJCK1Vzhsf4HuiD9XsxwuwRpwb
rIsXhwyWaXs5mPPWaTlju/WpsTG2qSDP2QviNGNPUMhMDf9xEcIRbDvUzVOl1BdP
AzmNepaWtw6xgljPUr/vqcEIQmVhSAAT2+hI0Tfum/q+Hc9ZwMRe3iz3MsLQbjfW
ySuZWRMDOozqNRcCliYSpF2/iVBwBimgOj334tgPElerInrN0+n0lIE2zmN0rRc5
2aAU7AcfkdyQBKnHaYd1kEGjhIHM0lcae3F2thwQxuEXoadomYswQPGZ3tyN7ao+
cAqXy5RStFy34jzuQtcyX1OpBsorjAwsdKzP5OAAq5qQ+3xIZMhS2+E+MR4A2yHb
XfX/HMtez3rHzF6TpuVl62oGbzTLnp8NknLbWJ6gZCbpcEqrvDJ0TxGWrBonX4Qg
hEMsa12IwzAIoRhci0jC8TkSAI1LsoQiztNo4SSpt9KjulQmbJ+z8TEUL29VG0kz
eYU7som0CrCX3xqJ8wIoZj/cbeTKIjAJ80CXb01Wk2TCRa9xThZy18Na0WxAYORJ
2sbvP2DTJVYSk4PxUtDuCarJO3uPh3+hFX9dGPbfTDrmisUIxlouJM24iEVrjk2l
8CUMWqtLCsiFSgxVsm7u4ZSQ2uKB4j97XWZD7uSokjYZMjeVjt8vufnKSgtqQArt
PuaVI7iIDaGE53NglVlR+8vGiS+M3j/wFgJJ1UHkG3Gspg0X+WXWVvP8ZI8riWw3
f/kxgMUKAOG4bcYtdCYfTlMghppQYcr29szTpZIDJk7WdFTasKzMbu/bSqByPIY/
j4zTpsJO0pQOAoav5qxhN0Wp0oQieZFT+8vzwkleg/WdO4fcWwvRXxSnumjJoXKC
UdzuSUF1VFKdSTKkUSqXtjJTvXdIDjYFRUZdMIbnieCr4sAp0JLhkLBl1LsUdIPH
4n7vFBYgloYXg1qVcAdQoNBqamf51nFvtOXhwSYYdjewUSZ78rZ4tL+b4FV6u9jO
plN/pAhL3DutjnbNC2YmVE27hRY11Jiz18rp8kyyXDnCSx7KyDZfnzDgYu0OrGFv
dLSwtcQit2L4Y+92abMw21Wx90lKcxFNEITTPoK08ZzsFyH1HWLPeM808oaqQhLw
FgR4h0js8LuKTzL2367x7bIhJyPr3bX4aGJTmBEI7uQzOc1QK/bGg66rLMeKQM9T
TNUPRrKBpPNLq80lYgbhjwBi4OiuVcXkt3KqxUF2Ns0i57ILIcEUjEUx+qIghuSn
84zpvtXSNIbA2xXDyeflc/W3U4gAU4bi5GjXJmZWSc8tBKqk+JBEcvBKF7M0pT9Q
6DuRwbeJp7IMjPFTC+z9DxX+CS2J3v6lGmVHMoBrgDZGQysY9vwvpwRWnp/lAecS
wCMiupc9G7eGml/S8j0rSwZeDCcpIVNZbHuigmoZGU4rH1kKYGmCxX+3zl1tpRCo
2vZ+i8Y9DRsFy0sirr07Od9HlTRvyqN+wJ3EFoRtFUihOZUVr2oqoQ4Za36aEtc1
Fue9l6sbSpZTUYI6dItxlygrFVzQgmrWYUHMVlhpdyabBpKb1dVvx+c3InoNnEMr
0Qxd9dAib4/ifIQ7Uf0pKV1YnoU7dv5IPzTOvBnbWEJHL4XqUictpeTbpmTKWv6a
mCGb+hDkc/6ghr8W1ZdbiIXPiY1wpwXp/iOJxqTSq608ctpxJnHeNNog26hEHWSo
+QmHIH/GHyKf5jT6W7k7lPquiCP9Vn/xwanY86VQ4hqcgt6bPkndMQb+OzU6a0yr
NqMSA4RPuCmvui+LCRbgoCAWaGgDco4RiHCFfC0rED0BknsRXXT7P2U5fSH9NmKs
4EU1DhM2j6fszwUf+ErtYxFhgxcCEG3JW5nsRu+kmf0bwtApTf6vWOAv3Fj6YI3b
/i+tfB4T4NtXkIo/UEAZ11ZpHZ45+gSB9gsEADBqr/0kKHa13JjmExIn/KNvsloM
vuINOII7xII4HtljeK5FeSYftIOx5BL5z2SbAyAjDDtQZtlVItL50xBrqbT4e4h7
fNDV2UD5tZpQwPm/pz4wceBX1q4XkK42Bbf+o6KPTu9vAKnshizxovhCasjy9b32
ZeH/liJVk98xLg+0i7k4g96kEdoo6mG8uan56Otv8HxWoPavwEe8lych+OrJBCm/
BLzHloFGNqL+32GjAI3W/hy/BXi3HxUj1Gw8sQl/nEXAW0uMGhoHn0W4VVHbSH5C
8dK8daBkR+SRKffS4zC2W63Hwi58OQmJtMJIUqUNWhTOdjVQUKXel71bq/eSkMkd
zfQZmZdrniP8sW2OeZKFHE+2q5b2/PTd9ybw5QXxdGAYwvzB1vRpupjrtZMFL4SQ
98s5atgABKjcNbrOWy0k66U8XJg0FuuFut2HcTrgMkoDrwWKm0T27qc3GjhdVQub
ph+CXcEslQHT2n6NW/Lw5QN/M/s8obA1GJqCp7bW6pVog1J82yQvEttbopmNbYjc
IF3UdlmwHIlvpEdJUrnrxxdueHN8RjVaQYX4Zyc28/fKnXEH8d/LV5Rv7U84S9tB
G31LyF14S00sRgK4mS/SCoprmo7S0BrMBFsqdAuJyw3kPrU2dfYhhOp9PuNlzUoG
Ly1E4wFJxk1gxf9Ox71lmwfrJpHiI4e0sEjgRJ/JErUYM9RwXO8MwldEPSXV8vYo
mclbJ9I3PCGw/bvJ+c/C3tIua+444jvojEfwxxK3Jpz+u0BcRc5Mm8f4R/ntZl+a
HxhapNA4AdYg/F51Dnn4l1it8/3ff7HTqQQaOspN7MZEeov280Q8Ta/bXPUP241B
7Ym2r0QCmiaoOSvN8PZJC/5yK3IM9dpKmPrczfjBUlgFvTQ++U/cAqHSLdvN30pH
spYRnTHPPfn6LKPr7a4JZk2ab1ofnxgS1QK13z2UxEERmmu9thjq51v+2b5g5ZSd
CEMsV3D/OIzQUsIsGFo2sIWmxzKVUkY8sJ1iCeAW0gSUVRoF3sCEiZ7hCVoWmDJL
NNDOHyrNobRronCUKdkOCVhc4JdJXuYHBMiRlJmis01pvYHzPoU72xIABcd+q6f4
PiYXihzevQjKLMSHkqWFesxMn/LkrevdLBhULB/kH9qei+/uhTI+Tq8zCAOgD0DR
ML84TKl7SNWJc2GFSr+kRvD0JOLDCSb/+wAel6vp2dloKbRnyIYEu+yuvDh1cEWv
R4rOoF+II/jFFxnwQ573eDZT73okBic4nCBs+Rcwj8d7RJVHXvzLhLwUbbpqs7zM
9ySOKpYhm4vtZwIDaSrhgwvaKdlUsHu6whF02eUqPn7DwyTlQ488TNMTwKHuLMHO
uuaguaNJlpAMqMZ9+F8kUOWP9uCcvTtb12xK9t2O6cd1ASqhHBoem7f5x2/HaVLG
DcmvcmLCAX3JD4JJb/bnEj6GEckZ4MsAcikTDWGP8L2FsvbcLeZZE4bS5+Xr+A6I
FVRgYEs4R17fXpnrWfLCT2VxqiAkNfxOyXGeNdWrMXl6S5Ddr575N3+zFYFwbiJK
Q8JwdB6RypSCqiuCtYk30jvC0dSVm2HShuQPx90fl5EBPN87HA3uKrzijNnuJKJq
0AIbu9B8ZtyLGfjizQcmxRiBV3lXUmp0h7ZxiLdWsNEV+hL7Z+Fgru0EKH1lHw2y
3ZDpcnjW5Pqur4HxnptWqt6PXr6BxYu7+I+zznoVw9DIdwhbcGMqMW2DNMwTMisl
e6Pttu1SyoDvn2criJlhDey7eyknyEA63gTqapODJrzQKmx1e5jMOVILy/smcaYI
qnKixWEnyCO9qdaPQCjcKhJl5PIG5Uwl66PtTPJO2OHJ6boiO7i0f/f6n1ThK50j
jaVKueVKY8/ANHMYoZxTGIITp9ilH5d5jP5JiI4Nuqqn6qc54lQV2XBSJD1L/VVC
F8Yl6Qafn1JShrrP99ooLDDafkG2vT/nrxYAlk3Lv4iqgiD08LFUUDnRR5QZM/dR
pyGXIZEeFKDwRkV9XkzQDJQLbHOJCRKOE1LWGSOA/BXitE+DtQr4Nx2g6WcKZ/I8
/EfqxZUSckm+X2UKvofuaRtUrZhav6nJ2bB/U1oQBZ9lIlq0s7KR26XTAl+C27iL
/vJAIRL6nUo2W1zeW9qX8ykY59VpEkdY1iGR00hXGEXkc4OOECBfpDKcQYc8B5+l
edRcl6hfe3lJL6Rl9ijB5BdtkeU8GnnKhT+e6QKlQVFLm0zHISM5U0sW1X4Q6BG+
3GAyLrp2EwNC1qjyCnZ7bALbX2xGoxpDxfiAzpZEbm/7SuvKztf9pi5Iizy3GfF4
DV/AJ8XyTdkPQTBVXGrWgXSNFEwwbE6HiV1h4TXov9heMk15Sq+lJWVISJFd4UWp
vp98nvvq0oEZzsKzPMU2Onj7lSmwVjTyLmdqAHoMtuIwQugws0OX35/kT3n58VOZ
9eVHp4wBkHseycBDEG1t8Z86OPUzHuI/CTptt1y7E+v44bi+8O0hqMV66T+y1YhS
7Hxn8a0DFKdlW4w0eAjjCnJ9XRDAb5+3bbpCja+9EPxOzqRBq4KSyPhoWu4exsqf
lC4RllCkJMAEUHTKd5vNqUPW9Y8X9lcSqYaQZ5dtD9Ia42awgOmugaIH0yaMYLUU
bj0DrkDIDRN4Aqq4hiAIyfXWMIeTKOxw8T3vZ1I4Ot8w7vClBGIb7xvF9VGJgBmx
OHhHA2Sl2q+fjRl/rYCcZkWm+V1NpGSKE3x5q1H7Vu9jEMel3TZ25T2tI8viB6EJ
RAm20urcOjUYYmA5zrgdF37T+dOPepMN5XdfVv5QZLYypvvvnKOA7tJ9l9pZdodx
RqJ8C8MzG74fl+ov2yPmV11FSywE6g7JUkDLHyYBY+HYZ4pADY7iySFpzOC84HRd
WJw7DcnBidSfuN2sbDs9cY23qedUuRl7rrvy7r3YkYurG/bPEV0CRjyreEsxSXl7
gXEzt/vrD2Ryt19+N+dplzUXTYh9Gar2jJPqf6SVlMTJ0xo0oo0+faALgBK0MTgi
EkZOGwCndRUrLCvM7+spylU6wQRjTQf7gCgPQzBKMeTkfFcrNhs5+pI+0RXGdVH/
scZPQy11zPQZAf1hn666JZbYxvhBzriMrPZTMbfBe8NzbNaIkmIH6zgsadKRiyNX
jEt0wUCF/93TDljob8FlY1/gflzWFOpR/bCklIUAKGnFzYKDyHlrGxTvoGyC5lvx
uuwIBygxugaLJLf+MdJEN4ZnSZCmX7JcrsopI2bie3AIFhDFfLK7Nw5X40K4b1Wp
a3R+3wmGhsltpAVLyX0ImR6UyBy8StG2RBewB2/lWmvIjgbb8F8hgTLo4PYkbWuB
7SUmhtbS1nHj2TtMdKg98W171cYODTaxLgM+mTuefrnUFvp6XRF8mr2uroy+l0Yp
bjMdsi6brgMBPrZmirrzF8FI8CyPpIidHRTOyVwANqe4Yq9A2wMDQFJFYAIx+kNH
OvWy2nurkGLWEogBjgAJ+yUrXaWznFWPmwnHz0RQoIlLofS8Xt48RtpiGSWw2EWF
pVX51sYYfmxult9JXtyp4Iu6TKjm6oyhJOmKLYGUmdatHedCl5SRjE7agE+opxMr
0eJlx2w5aE8xTAHB7v9fWpUNJOmMeRAo5Um1hxiSLrHC5Yo9G6Dv9xbn8NaAmsUm
UtmSqPuuYV7xcEYlA27z6fuQRkiLsRVcoS5LltXOeb8TeqX2f9XskMIhO7Hvca9z
eeUXtmlQPbB/byrH8N6kw2jr/WgZ3BJo8r++BGPWLxtVvc3lp+ywHKPEkRGTIc0G
qx1zJ6jkjPEH+rNKMENzEW+/EllkSYWvjdTq6uydLPQFY5tUSS7zT6uhB+qEC8oi
G8Ne42EOl+W9DLDP1SxuVlKGV+ewmV2v70vH90XTvz81oT/5jdAraiOmV1nuBvEg
m5M/UoalJ/WehUiSddQEB/Vzz0Qtrm0S8DT7Ijp7c7PXUSGCh9mi+iMGj6cjcPEm
txamNUJ68P2Bl1jNYkQ+HwVZnSeKX5vuK8T6dTP7hHJZ5dWb5rehWDIWKqmKZMiB
DKP7yWb9uN0JKtnnSBHnbFNMm4cX3nWAi54/xzUZmWBCakMLELlY1DcIjGs2uMio
NyXX9pSsgbIxy24EqmVMCV8CiWpGrkl2RGmu8r5xlYD6GZ8q0zw9H34FENuxc9bh
UQE7dObJWLW2HrvFBak/2l9XPRCujQZm/JnVAT/QXrIKXPD9K/a9EMgFtfTbc9Ci
PAOTGB+UPWAJWway+i+rRzSOSd1oEzWnz14xDNBMgoRwwYLs9tkjcO5Xv3mK2B4P
x6JQW8+EH7M2VlK4OSovuHlM0WxD0evr90BwT2XYEFlIyQEfjbczWXQvc58EjfxT
55CSFlR+Phb9UGNeFr6n1K/l/QgMnEm6ESm3/k1Gf0rmOxgnZZVCyA4hFDJMH4St
7VXHdGQdMxTI6gUQ+zCb5LplMUwiJlzOv91Qz3HiQvqGOvmoqlwdw3Hm/nuhlSap
cY79/0hu/X6sWDW4Hamh3y58CYotujISFd/uyFIGWV9UILIZ4v8FYcMeJIWEryHm
6lOTRz+QRsoAZh0fYVCiktH/2Tm9E4HemRm4rt7NkT4ZT82Z/Zk/2RCZEzbZqVCV
hr9drL8mwr+kbvZOxjIDkP4fmIcYkoSbj+6iJFopXFIW3uCN5fitz5Wy9J3aWgwd
WqiQvyFJFyQyptc6TDU69levbXlwAPY/pCvwiQdXnkixdLhlD8k8rivDPunW68p6
4LJ2pvKUMhQdIEotMYRunQ8i4HHgoGQQx1KiZ4X0wX8bisKqUOfQDAo5VuucJrHC
uJ6z15mOtDuWSzOOdmZj6thbS4sc64Wc4CEZ3JReBSPiODtyRHbcK4qVCOHxLMom
qDszrPMTmnan3cWQjsBxFo09fry5U2O1vLSjuhcq2QSMVLwal1H+IfHA5+zwI6ks
J955QComPg31KgRjS/1h1fonunk4LnQHDI4TsQIaPubG+LH6da0WPp/OFD4BVPpW
BlgiKBp875tjrkqiMc3ldhan2IuTZVdd0O3ZBHOf3gf6RA2JQLB1a5HSruwFlAvD
7t8fjwe/e+a3jKpFBy17I8tyda9hpkSxOfJ+kGxsHVI3grT6txTSddqbo5ugmtxB
kRvFAqc5UWhx5ubCuBTZCEEJOSpl1JnCUJT5yAqSfhhOX707FRuzEtm1Y99Xm5qp
fOBB7/5Nx6SmO3c9xHrOSGRrTq3Lky63N/2ntFJlROivHn/tZIpNR5gika85u1AK
CqRkRJprO4Dp7yCBNrzAYLVFOqikL+XXexI5eYckyMN0ML7jX0Eba3rHRYgmFF7o
AkXoAZE9sWBOxsO31ivjgwVm2/ZWlSZAdKPvAopCgTuTAZ+8rd7jd5QszwlbWqzr
TH4cWg6loIPglqpg2ctE9891VuAe/RCCrEIljt4o0JFENWGT3NINA5e1+cY5eK1R
Y/NZzL9d+XFTsI0YcvQhCS7VkXKWX1cn8hd9xlGy3GmROjfCfSbTX5ns6CLv2UIy
XSyb/RrbF2rWOhr2DOuQpiV50uldY+IoUvtTS18CaqTcTK9IZKijvt6QksN+eNb4
NmIp+aFN+NapKT+yQ5qnvx0pyromSuVV7mChtwdKCTn0sThUkRu54guPwSBRl0m6
v+fgzl7CZP3po+B4OFqcb81Nc/WAbxfKtwwgAYz9jaIyhZjgxsOlDCaJqw6EGXgg
bSiy4vw4BO+ofbsIG2OTygBtflzy497plaZlAqJ+aDnhmb9I48Sq9d9sR4Rf3xI0
Rmg26CLRRhM4sPrfh///dpu2PGTL517LOvkEAYk4obrHJGe7B48IMLCIkMls58C5
kW8amsmmsaOLM//sAR/Si72qGG89GpZQl+XoHKjeuWzr932iSfMSonlIk5hjUvUD
f5BS0Q9XpcR+Xal12/fPoL6usE083BRdcSnIkzctqqtRTfHJnGM1CEtFe5Fot6JE
EpjufKZ3pMbZrqy/YZlGgLLSC3Dw5o/L/xbYeXloCpdr382yJxf5mLohq2r7IhoF
Hnn5oGFYEro/tMiqg/YQO1hsgwBMPg2TLUKx8+fXZMgQyZvuSMZBCXe0vXZapVjb
eWpcqKfQwzWF1n32r2qD01oXi3gDB8T0hr56AzN9R/xROT6vr5dBphhP3Ua7F1q9
eai9/kiDqySlcloBGmb+EdKu8gBw0U7dFMgFhOkVcAmnDleMjmuw/0kbIHdopem0
NPaPR3AUuXE+JQ0oY+nGf1n342JGKnNJCQP1XbTNCCDbL9i16f/OL8DhZImvwYjS
Vvcw8OpQ8vgIhIJWUiN544n0i6jW4K7YgFUh5bIepHG5f1ciHrZvDp6uPoB6x4gQ
R9aX/F2SkybsNz7zGyopwYv2RMh/3MAvN7ruNlcrFjvg4ojBDPuWSXTs1Odmka6n
97O7nM1XqxVHr6LznjXOYfAhWpZhrsdIKCvmYGbkehsdR3ynRwEmvQ4vc9MjjY4r
bwQYL5LUPEq51fMWrzIJLOVyWngoB7c38V9Qov8bhWDxnJH9Rg0I6rgogyeFlxod
4lmZ0RrAB89wvyUKn4nRkJkLzxb5Mq9yDl3UTWR//xWCZH7SFmZYod4cZMcVwSZL
556Rnvg1E1zpJ3GqNKHliksN0m7y84j6Fc5N66J6YNQGcLz7R9/iLN5xhrorXHPy
99qTU4xsEOyUCzLyMtT7UUjbh5I5tbDACskPJlIUZUIdQ8xSTltI/Rdwhck3HD5P
3zsiAmcTqIgAQ7aWh27e5K4l0w7r9Up5uNIsIB6jePcEYaLR7jkgBwwLz9/VFUbz
KgXkNnwZdNnww0KzLBB7jMJp3/uxjENUeVFzxuhPrcyv7VJ4ejRZK3r8AV4GLU/P
m85lylgKo6lNO8VNPYQFP6e+c4F+c/8okeqysX+aK8f9MFDWVbrPdXfO0pD4JicF
P2LvrF9eK7UPb4MA/7WeoWaRU5nhaty9IglohW3kptwbaczpN+iiZWeAaIHKysAs
zTWKvY6T5JmY2ATHy/wz5o854AX8m3WvjwXVcd2Fz72sa8IZm5TM7Izau6lViP56
wjUJHD6eAC+IXEnG6ahCBUCDZ9HSoI2dXvizg4h8FZ491lHlhb3JbbzbS9n4nGtr
rX9EhEys+SQYKNMHzWWDzBwFg4H1y1eDVwLNoeF7BHsX71NVVOX9yC2qjOGgukKM
u654Xqxk6ww3iSUQRy+pLHTQmpKBbK9IwlsfD94iO26hBX9bfu4L6gkjbdi3P4/Z
xZSCLyCKCAG/NR6xPVm3GP5/V1iP8wU12PNCdXSgKeO90cH4awjopYBDiRqpFZur
/u1EZPQJY0cK7p8wOyKdnl+h5gm0NBW63mCsRu9+zrnCKnz7qH1ja1PYhXsdMoDy
tsWfGIO0ixC4XrllQsfBuz5rHSfIKMq7s9L00XDmDM+lAdfbmbszJ7jPSqoOBiu3
gpyPBlJ7Hd21VXJ70JXYepYOoGKiPR9Pocj04oJ3AfLOkORAw2cC4OER5GZRxMN9
8DS25LxRItDw4IyxRUZ+1OzjPFCpVMp+7YHZbd3TUodwYN401AcQNHlYDs/nnl3x
6kt7dUmvaMcSZBIKy9McvcbFspfSwCvRXkWaAz4SoI3MhpJ2DWP8FG0APW/Pv5gp
U5D1tr/Vp477+f8xo5H+xrb/F3Mjv7z0OyrBLHYJ2IO2fcrXE4MEJdus1uW7gtJl
Dn6wUj+nLn1esgc9IWHN5BqFQ0I4xEtFGflt2v4hiT+KihjvME6CLKoxwT39kbE2
by8AHXg/PDq1eFO9V29eNZiNX1oBORgkaXCvfat+7oCHi6zpLTR0e0YKdf21VlD0
n8v9PoYdyAMSopyiH0S9uVZLAce+kZvj4lQQk1QPUAZLuL18HCzeX+j1ltpeuFe2
2tkrW9ccOD3AIZpRFSBRJ9Ok1Y80CRfJid0SgA/Lu1Y8GayNrnIMpFAA7CwEW11u
GDD5b1AlviovSBJad29YGckCZ/im3i7tOjbYUCLqmodYKf/ckAcUF08AMSbBX3gK
NT14d3iSYg5vVmQm8ArrwO/+bq79OQt/gdlKmHhvX+Hf3t4PYDqjgHPWWr0K6lu4
Ip2ZBGzA/kwvCSEg+EvrW7sk/x7TNSc+oxcsykZuXEFOklaTHBJXUGyxcygCwHMm
GrwQznD7gDQTMSB/hTvKn0/MkOR8FWA2ttuOS4HpV9hgdSG7kwv4grZ18l7NWiAi
McdNe9SOCoUWfeSxBBnJg4pi3LbgHJbeOBep8F7XI8PbYgpjKOJdS7WYY7rAnNbY
patjGuTDfh6y/Tny4WMD/EAB4BoYHCs9nHeMcahygZH6pJ2MXpwqbw4yUBMTr3b9
1k6SQCzmZ7zYsEdC2A9RwzltV3CcG66eupx5czA2v7FYdXp4Roidm4xEjFJ1yivR
eoB3LgCRXw6hWuE8BEvwaGlhSIQ0m2kGNEJGIRSDz3enijLwWof6Yg9QUbC5MkA5
IJZ5+8nTeDWqPYg8caTr/R7WlFVI39yCUcpJLiLdRqz2zVEInuNw1zHu20NoYvAT
T+0fFeVEzokhoP7Prqf84O7u6L8+3UqTpAKx66jwFduSvh41QWQMHWrXy+v06K9x
zoZFgKzoBhXobSknszBXq8kpbM2F5eD0GB+AwxuxSrigWD6FDNxZ0rdzIjfVvwxm
ImzX0bNs6fytHqhUxk25kvLBLzJbpZgaq8NgHMMKrjur82unw2l8RgXtqD5JHo9L
XZFHR6TVBYHfm3vTePSzq+K6/mW7CEXiguuF1TsDNr4PNGm67PFuJRMAgV02rUUB
9/jb0xSZi1DmO4GuRgrHKqAT9IR3cB37AsnC2XOdumapLBv3bezl6XCYz8AcYEQk
XyHAJP6K3BaNufczAIdXLKG76u7OqBPE4Dy/ruKet2iFEOUXE+NovEwhHoNm6MrJ
1N7WarIeneynr0/8BHkd4VdlVMSNSxnjbrdgzooExlw/QvNo26e+NpbzG+PMLnKe
2cM+uBIwbgPoaGa2z72ryURE1ljfMhehNI+60Iar3uq8d4FwvlHnsnSJmwP8aCig
lIHVSKOznTPkCgFy5yLfqdRj6EN/2aVTXf9fJZ6AuLq9Zxx8HV8oV6Uh3iW/ST02
QOMsWRNpmE/vGgkYYRsJKeB1CvKsGgwx82A0Ba2V282iq+R6m16+3saz56+9NKFD
s0ez+QpMfLIZm2p4C2hc00NSGp5vZidwi46x/3m4FuqKOX8MvAvYmy0T3/WiK3gq
UhjJLlRGHgb695HV8u0nq78hlQPEyJjYrhZkBDOX21dfwwF+XZ1t/pyxyszBBh7z
W5GNBghrX0icliP418L+b8+DPbOzUVTSqu2Wl96P+QxVpKxgUoCGONeZ+iJjsRw9
q/wjFsu1Q1KKP6OPSSaDcruF+3lPW0qH7NA1uSO4OMwVPlS7NVIQfw1yvoQaOF8S
PWTTTh/wM9Uh9HzbwNRVJSNPOxI+UlwsFHq+BMy2ep5cpWBrgE+1jtrw+SruyFVG
yLTIkoABXO9BxjKqUBG3nm5fdxrwPupWMpOlbV+9yMvg1TQta8y9vEpo7p96o1Jx
gLuDUqEjISvYQAhLmNZRTv7yHtHJQMIF8hbEDeccyEiUcQR6vTvj3Y7gVisOgO5U
WTSoVCDgvWeeAmz5uJfd0BNKUQxK6pBVhk63LmqNAVtiLj7qep0CIB2Yjf/BfWS7
U8hpQfXtIojQUKC5H6JhQQefzfNeovveNUDo4KaAScGfrULitC+QoPguXhmcPhme
rh6XiASYaAWdi29almCoKqMwMlaQCb/aU7aGzP2QWzNpqSuz+ovNcGnJXstYta3x
qMSk7HpJzeYp9kmSd43ftpft4R3xZ79abadJCVKDzjeJWQmzJSAp0n3wVFJZeMEJ
HME7jdShPp8G5Ry3dYpOMVm1FYCDSle4PL+cf/tO6BA+tZSJ1TWtR8FripvGjAIM
3GJUjjeLQGG1OhnK23Sn5DQEFDBL9p1yhY+nVKfNh7cU1jp1PZ6DoMeAkXxQhXVB
j40I1O/5hlvFXkTKgUHjM6PcrLr8TGOj3uvTUwLBS0C8lfjKCcqNzJ+0cZljcV1+
2H+8Of0Wzt5/8/FhR3j7/eC+63P1tY/KeeAkRCHOWpZ1YN7GzdwpJii6cM+Mjppw
8/pYhveDNDw0XprxRwU3y0AK9YQ7eNXf4mJVSaU8wivj3MjCt1yOaqUboy6gk5Vh
7XEjIXFoSjapbRYuD3jhK7APcfo0xeqWgN4nSg60ess+Yc8aom6GlfuFor1anK1F
5x8TrJ/3oMXwNPW2y5kNsaIcdajprIhnc30aq+Il9aAAz+ykbH/cHKc7/chuUfTF
8nzNk42nhni0By8s8tQubivRrGgcIWCCRVd/UO/6wbleqAERP8ugEvYqIiHakDHA
KaN90yV6kwDd6Woeyil+t1wVjCdC0jfTBnJNBAHtqidtVxT8vqY96mpF1tlDcVy/
VRHDSU8xBaHBihaFeGlrApO936QDI7YYNgKZKssxYMtQVJ9pbFgJ9clQYuu3nbxh
DbJhcsdRBOBavzD1we4asVhWHE6ydD1Cz0CGrPFnu0IyPO+RB/3aWoQBq2ooRELM
uedmlL3PvaDg4VGkBEsmODyd8ycR6NUgJwmgNZZtBUize8gIi6XnWRsy5lw/powP
RDnzbs5/HYOrsqDO43hpytmulVRI7msvl7GQqH1fl6rjFbUJG12uc8GQ6mc7bLe2
kJm7/NMwkeHGpa07W3Mr7VmU9M6ik7MCJOp9wvqYMIfwNw70BaVj6XI2hCHSarTV
M4JBj+NCMi0vK6H0uWTFGVTmihQQshklblgvVtZupTzhgRHf+OEig7i1j9BdRRTj
tqAippT6KesL4pAfLR/lI3nUY53tX81OxJUoMJgiLEk1trFQ7YetDdp6xYIbW5wG
1wabZDB/mKcc1h1hFS+5elQlNIe//xUnl8MzHlCw4Tu4Q2FHf2gDlgWlEp41NfaO
KQuWe8kV8q7ADVmpHmWw497OK/tL9EFoTWKL5tgu/IF+TSd/hTeZg7Ff4Xrp58+Y
qN36biglEJdOCPZQmD76mR/mW9MmG+4nkTDT9jxn7W6S/ZBXOfIlV/t/1QVb1bBM
5IWfGOGcJJtlWWQxltEOKxj7s1+yp2J33aefchQVa1drizO+ou/6TlsM9aK5alqv
IoxniVJp0oaPmFQbbmyos/0C4K1hR1icgN1UZgC6kIs76OPLFTTqDz8HxoYLD/bt
xYY5RrT43puGvI3CrRcwEB0u3HX3mDiE6KtdnivJJTi97WZrCIQew7/6yfOnM2Y9
sNIeiEDMmUcfakoV6jjMMBHpbYBi9NsVouakvCn25nmJU15huSj1X1kMuubPvE7K
6cEzAd/giVXgDTUmZkEpvskRCd7RAbhzN3BgKIfU7I7j0zBwo7K9chaR+obOd4Zw
1MSIPcrdvEukw1pP/VeF7favz77RPupxmFAcv2h6TZI4Vul0dwjUmChqVwGsVlGI
KOmvPUVgEnhGE4np72zYQbd1AHlekOvCUJbLVl+RXvU8j8yuSERWFHxtG/rXLFqV
yG7JTkXsiOgaLPchWcaUysz8KhANBQ9x7aGrBMjFQlufTQibCa0c46v82jSXWB7f
xXyQHM8ix+o8eT4aB6uUxyagqbyRReE9+eBJilivESq7IG/sRME+ZCnHPMo6M4Op
bhFmmeKNPuD0IVJfllqgEx4kv9DGTALyzsFyMRB0lVGfEUzYI5o1NhKwQ6okOE+Y
h5XShsWcuUJ9BWxHbuyB5vBKJkMRKrl8fajpXogZsY4lnKXKICNc4SwQsYY0h4LP
NrSleWLqIDeVk0dcWJZ9l1Fia5Fcc6O2lH5hs9+NLqFrU9M+iLzzgtIf6rzhckXL
DpfHhymqK4lqbgPBPWl6cqVWuSNE4bl3y2b6/kbkWlbqHd2nDUlXZPS5ZBwui023
DthKixNTwONIUigaeCPMS/SknLSAzSohPZ8Hmzb9kDbqDPrZB10GFDO8y3eTvzhM
z1JTjEhSV6bdq1w2oDLXIx96+D2G/6KmjgwhYBDwsV8KtLD9Idps2Xws166nXOrk
N8zr/GUiaMbFnxNKs5R/IJhMZ8HpdmzCboHAps+RyW8BzuEYZ5+o49Hut1shJN/y
H3XxY0wkr+Q0NnULGGfvdIDySBtU4ot5AY5QAJqzJxyiMne74pcbpJbCfpjq5Psu
gn/DnKgjJgezN6KaSzSaswWiOZiWc/rc4JS2Bi+0YTzjSNpoGHfH5I8c1R353Kc4
Jo1FySFBaWI7ojVzOpIt9IOqG1cjd2XtHJj/d5ZRFha4xXvEADsoZlmdWcCdt+at
QTbeP9lpdxzMvP2bnzsCCHhh1esU1hrZflnBctyi8nO5zQ4ZkD741z+F8hwNixkg
wZD44cT7yYwtl1g8jRXCbOiT4iL32GO2VTlJ40PTwb1vpPJZSO2QhE8QCbuz58VH
TzR2hCDyuKTbKFul3lS655e2xrjHMA57EZtYOtRFaJUqpD2CQGBDZdJK9eOBRhLU
lPbmVnOD54ohTo5PBs/u9aLVE0/OBQTcRe5gQxEEyoUrLQzMjRx6NbTrhkWCasGj
eKHWQlTCAN9r+exfikX1/APFORiwgHhPFOO97pPFVoPs1A4Foq3U3bCJhXxfVZFA
zudb+twf/5NjeO7BvVvmWe7TNLx/TpMMCByhrF8qJ2oUnxirDxoB7eA3ckxgrskM
Ku2VvCyTegPbtjmeBbU5BA2fOTAw8zt8+rWVo8d8YQ0WPqSlQgiRm0h7FqEXzp8D
+lvkNYpYP17m0WQHBAbiVKi9Z69MrhrT5zbiZpIDDzTJff2+CjXl/fDnGF4fthyL
WkBti/zKoa4w6eO1HfEyqGC9xKW6sqFep1aqn98vNQYoTpflIEumhQ7/wnVuswG5
EFHBRQ0cIaf4aV5TOuJg+FkBiWWhppppEeXpzk+fCVS3vZf76DtrHq1P3lBro8Xk
HZDo+mZOkR3q6+LF18m5/yh1WNvSKJzE/x4E9rt5aDc181HIJzzXONZYfKIyzJ2z
DnFc8vGA9dwx4yr40Xc2Fr38/KeLfMehZoLEptsdu1xo6/fBT8P1cFW95Ok2RPkK
bcSp37Ccipz62ov1dT5R1E92RSM9gZNG9z3KLCQtzWNKrDMSQtOP0exMZvUIoyfD
OVM2eO+/cQfkoXQP8iJD9pYuZxEW3dNvxsz91Df0vfsZ2zbeYL7tMe7EMZDKal0V
FP4o8DnAnQsKxQ2DeJTSS38yT8z2w7WNo8V7i0bpGkrfA7X2ObtuOm8j24KSC7fV
GaXATU8uUGEPX5t+xvg4udGiml3vsJ9fll5bPawDZkeBOG8BAmVrKxtvYmDhB7Qs
cz3/T7D5htiwpGT6Zg3wSjqF/cIZN1GubkH1+mcLmi/SGS2kWxeeeZOxvEoBeyP+
ur1GDIGz0yl3SiqfQs0RynkIlptZzMIaaAHQqCHcK8EbbAih6xnCvQBtgO9Jz0KR
uVCH9dY6osUL6RIIv7qWOArGlIVHv5mvbaGXyGa+r/+3pPVIew2RRnFLHXf+pR7c
tOslGgiw8IIHUCGU30Z+v2G5fNYTXMvgIYe3FCgpkzwgRroq30cmVoP1K7jhya+U
x02XzeWtc5F8VX1qeZs5WYXr1K5F69HRFg97IRDeFNRA6VpRTj2bIj5Js6/s/Vi/
D4WOz7hxZ2Qoa8LZKpgJnvVbcyXYAwvXWtOZzlxQPkzf0qOfhmanXuzOqaM/94J0
ngDEkTI8E81wU7/pnHOWtDIUhiUIhXZSAd8cfyjFrx2phJ/SKKxMOmZJ3OWmVlZd
Np6kmp203YUhsCHJ3b58faxCJ3zN1Q0MP/6yW/LgzTkiUIjqmZd/sBteDr9m/bk9
eITYmYzvlzbGsCkom07V03cLKFM8fgAYkfEHaaXRjS/9oAITgu3fyefiFdMIv6/I
WIbEtHp9mJDWQwYPyLAQZ3wiS9GItcMl25RLqSbTPBlBbyoaulLo7VvuwGIHeCS6
QAPaYpEgsuErSCw2u8vYrW2R0f36XMJNSenz4aZd4fe98msvZpLm+68XUw8KySWq
pN1fuAKkIo/4Pg8svCkY+dKLidhO0swn4gFjC9uGWW9eooy2mmW+b1mn9QKQSkNZ
tngh+jzbu30yE127nj+ana+GGne6NcXb3Rbw0wI65nghtK+SBc6lusQw5feU6zxD
gspVWX5uxaEjpe047JsKgVuqAvIyoP6AKn7NFIDnrJKVOUc0xKouj1rkWlghcq15
38rpupOWK2oOAZo0ICs/TIitjlEdMnqJH5TFdFAjQyHUoheJvfJxuQcL0z8vKYSd
qkYB9MDwSiiBs0pEf/n0vs+oNX2/HAKxmogOJZMRDchpG7hBObUbLKxg6gJgfGUX
kD4PSlfZY/Php6qj+s95wdjn9Wcbaoqi5wM14z94ikTNMklL6Ibk6rTzFKNhV5jG
5OgaBwo8H8/rleesxg42gbdOBdS69/JpapiB4v+JlFyYWjILnS91seZ2HHiSgZxT
N1uOPPeJzqvqa4pO+vGGBOMSQCSOMFd+NqkINFOIdLgN3KGZ6zDftLViZmA09DPH
u5oleEJtuzOFOfy3mZqzI+R6rBGH90Uiug3y92ESxM0DgxFIqzQwJAo54pZGmpIi
9HZ2VImH/HynVooYyi9MEoCNIE7VgcT6theiMWRhk76txHR8ukSWHU5oK/a4j8DP
THHdGyqMUolDKekSI4EoDII5+h9mhmfI8ARhnTPLmU3dq35Sk+gtTP5FhmfyVhAs
RbQ49Nn9c79XZOAE6AB04Wcxox/blUIyO5nEBxkr9J2tnDgf0v/wCkvQGDieLAw3
tGr6Bg+VUJ87+airlx/KnRxpV56yObq0GtDEOhyInmtQWPPbzUmC7JiumQvmuOF0
HdjIXkfy08C/GYIeeNpb/vFKNSIEzdV43/XmgGz9NZZ8bpc9SIv5ub/O4stoxRDI
G5Ei1zmQhj1tqyqLRe0f+VG6Rb/1xEmR9uPi+krik81uLDU/oz0Pe6Rfutnyb3Gv
sQ/HYqfjhuekfuhp/j0zBDYDBorVHpwo2s60i4mC4TTUZueM+mKKTQxUFT/HyHtl
lt9CHQQ7L9aoK7MgNV6YpRzlUp9FiScBP2xOkAD3F7dIduxP5tUigiKL5ygje9UC
3dx6Wxis27Dgk9ouZ6FDeCnwAOGL7P/wTyifh21gIEwjGluUmFfCneOBkVn5mM0j
7rdZI2hmQQf4xC2WoulAf+nsfMJbTPnzOlPCNRW85BSSqR87oyF9LNxx5XPF416u
u3lOvZrA3Mefq0WTL75lVkOMv4eST550wYgOcNqhgYuiEftBFG/BpvZU2MCA+SLd
92fAflX+kgEtyFt2OpKPkXfwhVkmr12bMnv9vaoPhmbDbm1a+eNcdJVf9xpunmGA
7cr1dp4yzq3sMvO5zd7a64vno9TCXDvAdF9NFeYL99hiCNluoES86g2tbxvlSIW4
VrGjLnhC+PRb8/gzLYQ2FD+Ck8RfcgelvHDRdbwa8P8DVN1eYVsNNQSATqh1nIF1
p4LUYQnqvGUNlKIF5C/Y5Ils/2YxGhYVfbgUlxMHL+oD/Iah7BiO7IK7gIXmQmJM
AYwIQrf51PTQKFtSg8pJeaZjmlZN7j2RF21L3RNSTHkVTkuF1xx7TO0HsRgvrVJ6
hSGistSiceN8e0uJP3Mo03x5uORZLT8q5OKfkA4dUtWrhRICj30fnkB8Ud1PtJSH
Iiyzmwy4F9cSWbt3Qex27So1jcNoOpu3zWP8yogV9mI9WVkiax9D8oc/QwPKeFva
5KR+RcaNoHm6ACi6EeMl4yey+FvSU9bgWOnPjwBzrvtdOxsY6Xeyjfd6EvUd3PPN
7Dz7zKI9IkDDBlYbRJTEhIx1SbrSsnudfRZo+0DmfD/k86lrVEm4nUIR+ZU5x3xp
26jHZSpquXrkq/PJ5UmAnONa8meMzfpB6yssSosSmMiEd3yYvo/K9HMsGWslOsAp
QMKqevfzz0VCIP7jPeCYbzYlcvvQqm78epkZQg8R64frmuJtKNdRujS5ZU5laYws
YuhG507wG0A+wsyl04+Lf10syq7uIvgfFE7CMyWK1Ane5hp508RcOUse9DLPF74K
NbtHI9rYLpTdGsd4C3YQbfX/oDo/COxZuMhT/gt7+NS0rTh3nh4B9trjq97EY604
vZZAv+q3h12ussWgZR/craz21Xjjs2Xfmrp/EpKaBpLROxTvT5Z+0Y4RIvvPQXr3
Sxzn+j7anR+gqPcNWN3IqbIL8gA69tLw0FWL4tZOkkLkOfnqtgPJZvBZMz7WqLCp
tWepeIPEmygKwLL+rSTdURC+j8lDKbjM+icr9Bso7ex9alOiSO2YIgyfaI0CwlMf
YQX8rlvZWmALna8mxegyWsJGGeJWoB31gHaf0OHCvUBu1LNG3QMhGivEYZRFRXHs
0SxFEZ9E6ky4fkk3n7zPVqZEIQ+iwHrTh4/cz1YWrhXINPQ2OGTGfKC9RHAkhJsh
Zy1b5g2NTGxCLiTRpIqT5/kOA6R3lGmatmVJy23iYCwyRiil9OvtQyoUiu0htg6k
+q+7w+APY0CEuepzJ3Swjd+DZPdENqZir2J1IZidV7LDBBDpSB+b9CFnNuSeGZlw
SeQ+j4VuyO/LAND+vPoKVvmKP6BllPYaL7KYtv7ccy+ezypAEEsza40FCDzrUvoz
OY55eygcM3lYXyrx+jdhZNtE1BQ1/chJnIy0eiYHLrVpX4tv7GoqIJ84tt7mKqvj
vbsLyGKDIiOSuCPt0s39K88OgfNZGibTw197GFRBUnQNUIGdlqlle0tV+eXKMlp5
9kVRQZqQyi/FdpUNUHqnABhaWGpsQ9PB/a1dX4df0D+GRD/xBV6s4MGenLoIDVwy
QnkS30ow96M5byBzg5jnxiqXXAkLB5QTEEWiab1sMVZyelK30EiBHF8HG9LSkoS1
FIx5LmK8rQtuc71Tv/7n1xU313zoi1zDFTAy6K32e9J4osuieqI44d7h4Elp2P+8
EGfAEUZKsFbSyP8IIgpeHe/KZ0ii1fwCffnyUcTM53zKZyk7AwF3rYc26AEAgBV5
9G30rI2JYx46/ZuJ0t8pLNVGsEzrSuyoOIDKe/1tPz6twdDSBAJkD9ltZAQXv7Jg
Lx29LlYMUUptfbihQuhk6kNMXuRNhvIoExfx270zgyKMvqY5P1qJDiaTh7DgUuhS
jbYwH/BUxepKAYOHdDztKvd8GT4IT3nmEfXLmfRTAVLNTWeNoQyID2/qfPSu1vSO
hSx25efCguwgiAsKcXtkmgeSzv9ObEdmTtbdlej/caxm0HUFcEHUxGcuI4HV0b9x
1Zj5pbZzqMIwb8XxZ7hidMxp/gD29HsGI28KvPHJ7LmH6J3VY6Pt+g0EMWVrk0hj
dj8FScTjijMQQ4baW54CqA62A4blkEI1lJVqzs6oL6imAWDwWl5Gge9VOUzm9L5m
dYwsgnLEpsh9iAp3aO9ScdVq2WcYmwIKLXAZ5Fuv00MBO9Qpc3poY0fkUs8/SRIG
peVMoCbvtxUS6zZQxHcSu6QuaDeJmc6/GYpWUjekloFffiwO1WVVaEj0Iyyqcttv
0pq5CyME497/lGooaInouaijhV8N1XGbbONTLHzVkf0Oaytll/0yD468ZCmWpNwU
u5a6XkOhZivJhZ3uU1WZ/KJfmcLwmlJLHj5ZWMWyqW3xWijHGKU5KRGmReLWNU4b
rXmvxFlwWyoZR/sPmr1WgkcnUwAj5yw/PPsk2Xc7ULhf2g8IOQjFDIkIQMjISfRP
chpTv3rFfEz2Nbua7thCnMSEAy0bW5AMW552bOokXYShP5rUItmAv6rzXHlSOkR+
bG6UxjIZp99iANPVRUbz6KMaD0xhySZDM7EqCoAoJuqOQ2olYTcWOlW060iXw6b0
f8RocNMDfjEhPLfoGrAsnGr6M00ldL+ZBn8IgK6aFarD+2UdgLidnscpbrw0AOQr
X1PozVRIO0lTM48wKfR4sFq4u1KqWIazkiYs+Bsh36TipBAfxdVjl2ux4oLd6R3Z
Tg/TIGDy21badwn66uojzeZ8Mb7wHw/bdCFK7IXI8LB4UJJAtgJlpD9R0cudkLHh
KFSHEUEaKMcfa7aXCo8siobaTIqEi2SzCm8G+NIvyvL/GnR5O6tPoCL2+UV84ysU
x2woZkzqfJCMWZbTl+ICsCB7ngVYQkh5w6re9+7wL85jrCB0l+hd3eTs+JqZizIZ
cxWCycrSDGRI5vziM5h8gC7ZdioPsgFwAI8nCg2uAoalSnyuaScH8YSeD6gub+TE
8XZ+/dEs4qfyTN5Vcd86hR9YrMkRnvDiowNNZX1xSgtGpt9baFolWAUVQgH7WwT7
xYj67dGRjSHqyZUB3jYexe77qgJ+KjIdTCRac5xy0u9nzsGvIraFHs1jPpPqL2Td
2Z4mL2HEFoOV0GhYG5HfpzRzctyj7jYj1mpa8mWg1qi3hBtSeqZ6DrKUer9trS6O
GQHWXqkDMlB9XFdofARLH7+zCLl9MqJHvFQSKIgJZSp8hsj0XtEHetLdvYBL4r6j
nLp4wtzKVyds+5E7mmmQVvpLqltydz+Od9dP/DH6yCph5L52n3dwgZhp6iYGSiQ0
z7QiFQOJmVU2fLVKKNIH4XGK06NWc1pjmGbaIaWgB+zncTleNpM3NGY1Brc2MejA
oHbt6+z5Oh8gsApr22nZxlY0Qqxnem8VsFjSNhZK35sBb4N/8TH8j24AO82ArBm2
dFFocrx1YW5t/H64AtkXmbZjaMiVfvrfHxbyz3NQQuZ37JQL+O9KLpyiJztGG8AB
FolOAnqQJ5k8+MMaD4hul38klE5jPC1vd1S6YkRotEayiakwi9QlPXHblHQTyfJv
Pc5lHRC0ha/oa68ywwO/4mFPYz7KZ8clDzeB4NfWUMzlEup30rTP8Vi4bwYQhRpo
TFd3fVUxgR8giV6+CZJWUCOJ4Fs6eLMsoMfVCRogqYDZ/1zW3fWvRZELyM3T0JFk
bgiaN5X67jD4Emf2BNdgClz8mcL7risqv4NappwFspe/S5kuQhXDmf91rW1cpTFJ
3/F+OHpjSPF8p/JGUouuHrmhYLlUDneC5cRlTHMrijHisqeFH6b0pdjn4GyAoiB4
vvSUHRT4A1sxvc2oOGmr5kbPliT4TL/0TqFvVkgE1tcnjL1QhiRFsODZRsDsYoCl
Sne0mTGgku0tjTwvCASfXasaSgpragrWECJRcF08N2lW4ICwg2NfWfgDVHrAjZB7
Iw2Qk+nQ1kA8xbJOEl5VljeHgH0NbEjh7KdIwKyHJObShoN7SPzMztlPaVdPXZXF
6qvD8/m3z6+PLO3JvBFtDPOvF1CFngS+MZ3QgLdnsTYGcd7Ryu0FmDjPFrwHfTSN
LiKCUIu6aUe5b6JbAOmsPdfvO5u8KLvrGUmzuWwbhqKXjNkdYLRh22tvBgshWB/7
Occqu84o+IH2Vw2IzANtlrt9N65Jm2Rd3M3YIDCcq9FvFYdVEKYW9gptzd0m/eIt
wHVdoy1+L4C0Em5Pjhy/aAIl4HzpqSHRMBdU/ZYeC4NFv5jOV39lR9prT2CC2BLz
VLLcybPGzu+nQuJRndfnEVK4fA/n+xzCgfyhbRBn6wnHokBmIT1Jm64PoecFIxlC
ZAhUOjnzsy1n+6ShUONHuN4LdctzPRLMVCwfPUiM+Dk8DB2Bzz8839hb7k2sSnc2
KQkF7EPCy9E4+9bQqPFqVpdX/XqWuRXW31sboIl/djFivjP6OjpIBi6auTAYNZrE
YVe4u+yfUy/JOZmPdI8OZvughLgfbIgHn565j97GgbEoMQFX4AqUccv7XRRUehlF
COZDDLSuq4s70rTbDBDjHY+PyYpUm5yauaPdpejarHx+xpVjBstGn/p6R0yAaYPO
H1qytZDXzUkWAFJhqPWvxhV74KDWxItuH3mp4OHWc6YG8yszPuZfkzI8YaSFfNVT
yrVswSml03Z+7Mn2vvhpcC1xinqmmU3bX38Lkjrhnepkrzj3A3dPaNqz55ut+LSS
GZhhnISmkEpor8TXQaArt71d6/rZGXoKGC0MT1GNIZ/4YJcRUI1SoVufZG4tZxM2
b0MUNysBA/fUAQrYRwenUdufoK+Nq3R4jovne6vYTAc5K1bMJQIifvCtPwiKpbRf
AwMtmLXfOnaqkE/7ttHm+E6HDKSvY02L6SEITPoJRoYKfJYxYsOmpCqC0A8KQr9/
DTFZI6N6grdygsh6fAwHc1kquPiqrJckxvzAE5TFjjv2jeqxOOXtIV4p2zxzOoa5
TH36Ti2jxwSHKfDoJNdHV+LSQibGas5LddGmOZPNZR6j4c1CMg60io118oXdFIxN
5jA9hBgAli4nQ6aTGQQeMtrkz1laJhiwOiwRdRjsmUBHkl3XOUG1+UZ/fTyfuL4g
pzhvPWYriEXoSyzFv0+0d4p8FG9+pqq9BsvbLefJB65zdohh5nwipwjA8M0G200F
h+lFX095eUSm2uuSTEeoG6RUQjQ9eI//uw+uuQ03CtPbTnW8WNQx/qsvSvJh3jiu
2c7ea00z18yLlIPTqcBiaBApBFic+IClGcQPy1/OHJeXsj1+7gZvDUwe9ekAsl8c
TkSYbfk5Cs9VKmJc8mIyWODUfD3NqHb66GWZqhgULvubI3/gUVjXn8emWMLgCAss
yTp+uB549DRNXke9exPKcHNLezPQLE0DBHHcUYI3s3Yqn3ve9PMh7MpGr5vMlMDf
+rkiR1zEJ+MDyX15dQXeY8/ma1QTHHahP/SbXK/hHFf8hQgxDES2JuLEO2UdpEIZ
ydOy83xOeVBzKwAn2LHYXlaTrgGOUzpscPTz1wyX4G9d8USdY0ztIJ1cmQrsokuA
A6L3LsZMnxcm6vSVXzt5A5Bm5j5igGV8WRGq17k5dfxWfaOAWGjeetI6IgdS15l9
LRCMJtMOCL2BzR+OPquVjSDDjn1EU8BIT9t064yNiHvX7brCQvKD++57TKBVjYjX
wuHrirTuGotLVIdyMVViaux9DE2oBMatDBUvwwmbeDZSZanZuIimJIzVrV8Zl4kW
iSHtVz+4/djiDdBvCLPvb2aGRibBVe0rY4RMcb6qhd9qjxzv7wJzg6T+SE1ZmueH
q6i/9Vt3t1YcALVVTJvim1G9ElKfpSsaP7rw63W21CArg1LXifDHzosexT5FU6P2
WbEDBX0qiRTL5h9zou2Sq3HjpswpjPQjJO2KH7CVNXLkNEAd8Rbw6vgkdXXudWEv
p2hQrMiSyud96thunQxUaCpaJdZcii1U00ajp0kU50gme2fsI6E1ZR9r++F77EqN
2PT1CwwwcIZuX9FAuL7blSTV+to3OjeqpnaDHJSJGCdknJMbVqU+zyU/JDDk4PSc
4N7cJhkRvLxS+v1uSzDrY2drtjEBPXZQj5KoEovGv0/FKnuY76+5bMIlTvf4qDTE
iDd/24o577TEWTDvO9H6B0Jk/O7aIEKXaMNVNqBI7/wNvK7pDxR1GU85sGPxy8hy
Dt2g8vV4uh9QtviZVLX150pzLGsMEUoEl0s0F6yvX1AoAuceCGC21LlO9BT+xb1j
NOXyjJgZ+AwkEBf8/2MynKFVzs1dBJQek+2ReTYPCmgS7sTem0CT3pZLYPcTO3F+
czFkZaj0fPAFJWiS2CT0u00gM10AHtSrz3UWe2BeUHEFu8yyK5srexRKm5ejhqXl
hsmWEVoQSrskaBTpKh9499FBgdd2xoXWZZWCoTSMAsKs8XE9Mdneaxwyx+qRUkxJ
Z5iy9gwFLocqFChoqqlialyWmORKYLviIa2gwZP52HJpdNFrm6Jb6k/gaB+na1tO
zDK43VPCWhRyezLkogjkQaRygvLZymtUgtwnqaB+2s3c/8Ytwor/6F+xR1BNYbO9
SS7PBwm3+w8bfC6r5vg5xtWVZFa6MkKSMsaM2Lwmn1ABeyDxMfXsoM7+65le9LtQ
/w4fvlUNrvxmanouJu9siDTtChWgpbU6UyDPNxGVoDvqIwflgv7447CHsSOjWEQ1
EqAUM/cusd8FFALDcBNlr3eDxXV1B/hdLEnpYTrbC/9i27tjEzHGxOYYQx/XTUON
8u3hDRBx6+ytl0CYh3IJbysoPRMmQL7+kpBNRqz9YDwpxIcHoWnsPu3kgWPqEpi0
lBrk434O8OhkYj1MzuXbIy47tq+PgfHT+Ixbq66Iit5kpo91UsyF6SyFb5EOS1V9
wwiCQ6ct0Fr/gMSxX7t1FH0dxIono6XK3rfzBN0kV7yAaDkB4s5fSx3LrIEMBBd9
QTGbMesTPgobqweah4HXXt/Xv8b/wSOwEH00MWbco7/iO05IaWZp8gT585Tk1uFx
/twONJYzTq8HGYLSqWBrg+X0raKq88D2jrUs0DbdxZodgcOMacLGzsOLnXZuml+U
qMortdvPwgW1IvJi1FPXr0HnxGcDCn96StKjnLYPqLIgSynsbm60GlvVyE2i8I3B
4HqiJgFCOB4yuU8UiH/IBQWmXtqjRAW8ap2GBS8AZkNVqF+DqT0gYuC9L4fB60Wa
jqD1cjXXqkPCV9jiyi0wwYaKyr3/fZk6gkR5b2TsPUOfz6KaV7+mQZOJUzJUqbeG
mD4/l3PRFUq1IlJFZfvh45mGee0/9u1NcMt3XVz+6tr5z0dnMrYrdzUfx6yl3cz6
G5IqVK66DmqZP1NP6qaLxCmxZ6liVmQf27cubVfVQezWnKK67N1BmlRqT8uKn8o0
iofZt8/AE4VmO4a8D1c9m3myQ+nrkKbMSPbON6Ey40OEoQsSfDbS+6iqWM/D9rz2
z5FWagJqTUgY0bnt+df+GVfKAKPdoerpEmjtZEofTa3XLwZLa/zC0fGcr+cNWUTq
LqFmIksQmjIrBYs79IGGMFQg/Z+1/1ocGp2gLUyZwynkBKD/Noq6aIgyiwpIvYIV
DC4QPjBujsUiqtZxZ6derd/3glvOyAnZkTp629BnEbY89WvNHTYC6r/4Aadiyxr3
pnwUvJWzzz0FmBs0nBS0k5jnkOaDYOaKdiO9xwWReoLVu+d7OQTUCRrXXmJtqnbf
VNGKpz79q8CsiWM7FHtq845ZxRd3aTE6Mj61aiKUGvGhwajx8VmgvnOMvSBv8lT8
fgcbiYAG8VoTAkkLkSqTav5l04UkAi4N8JxypMGuU1CDKc3aokKwq+iWK3ZMp9pu
g4losd9U8mH/Y23R2QpH4pxhf1HDJx6Qs8++NPZrR+z2r4XNus6qel7nnFMfiWOo
vec4Tib381Olaqm8PaTE2EmBDrm6oHNEapmJ5G1B3bJ1KDg2bhLfFs9kuwNbV3Bv
m+aEC5YlNJ/zC4ufsKPXiy7v1DispIPchccE/QXTMjjcvgJ19v7XzQh+MrWs8HPc
fqvccliPYnEcEPQ1+gDWCG2d3NawAYia++HDKiDMhe0uC1bIrdJkBFv74yAwTNSx
8BscY68Z+DsDdjG2XfuL30LkqrXGMbKjXS0JEXzo03io1GcoHggsdi6OcyQUClfn
vohY5/4Pr0t9wEuGdu80jOM1wkf/jLw8fKO0H31RvcTKUlgU/sdwUmPFJMtu4mXV
njhAcBb9RJnCz7EAQLmAmK8oWIinnjKVHRfypy9e1yOWFbiQftDMPfIUUF+GgQ82
APm340TGWH+B9Y723e+qULXa4UG9tWrJfM39UawPTOjAmu2wL27wK30Mz5T/rM/2
i+8NU4vx70h5QPpVgGpKXqZHFZZZqp2ndomDqXso7b0Is+5VUeG8ZQGP2TuUIWnV
WSMLcJHQIcFZBfgy1ZfocXN8eOrfVo9wULYMbkisAjhsPHVTPYX08/xuf+XmmOAk
MRVt71bO79nFmr4J4FZFttsjyjC5MEd9lFWUA2f8G/Y4Nal8yE5JmJDFNHjzoPQd
EM52fs7jBif2+3T0Y7z0QmY8Ki6SkbOUiYVIdhGuSEEkRJSri4AB5gWWNTgV7cig
TxnTZI/b+MK7iV0FPeXcU22EqeDhQ69+vhaOmfTl1eHfMR8SHYMT1y9OsNKb9UdC
uSQUNxTlFfMrhjt9Fhg7IYD6hVd0GI2lgZUU/N6d5ihdh0H17eEDJ11bXqCPR+w/
/aRX1MxESV/mHFh+NqtGFTChijLGhrxWBlWaEWF2SL+Loo/EnwckmT8p/h9zhK74
ng8ihH/vKlbc5SReSsHWkZYpX2d4OST2UkMRacaUQ90HCNRqJaZzan0/g+b2XrN7
WVm/RxsqznqO9BKyL1n1zFaGvm2WE3dm/jIvKr1zmXd5F+Badfxueft0LIUyjqxr
mxRt9M4nPhQGNLZRkWhVuC7Hh7GyB6aKNxgn29DWWTXZncapfRtsFJUJ6O1Qp+Cm
JUBH+SF9mdn8hurkw6RcW7PLekbt8+Lwrk7EPoo3TJAdywJqRUQ7L154RmD57ZC4
+uTENl6q2OViIcDugXcv9cgwWN2IvFphlRywk0fGi7fZbhMcZZ5lVzAbRoPBOFj5
8vIKVHzMkP5AS6kBn6SxGFQu+mODl5jKve1qQS5bBPpYaLzWXA1kFoOFarAnl0JC
xspEbSwx4bFJL9R8zrlDAuxOyfQCL4Ff3QDfzHur4IVQsCsNJfRZN3eon3YIc2VD
CP9R57yFAWXaBOlkTEzJEq0Vzm/RPL9Mnh4P2ebbnThUZ+jVfjawPYsmPR62oM6f
CNawtMls10i+X+ipf1cl2N8D09LR/+8ns5g1b0onYHSAghzhKk6nSthZdO37gi0y
CmDOYcMgznHJ4oAflZSiTntWFEZ/OCbezEV0LqgLh0HyeeZXW+2Ivs9/KeeLRFhL
WAh/Vj+2XX1wemRRlByEljYvaNn6JDVZCjswgkfUMcnmKDBes6UeWZr8nz95Edg+
mKHkx64crQROcO/1D199l+AlU34sd8mJfQ8gA8EoXN8HMcJ1Isb1fleIVYN+NQBe
dknZWukNyYYo2MXH3Hdx2YZoNkAI3KXIwS7wOAlsEedI/VnWpCIaSCTFw4iruDng
dJhArcfO5e6AVE/P3lhoaBi1785wFXp0EXufcU9Xr64ppyxxfbK9791zMwvQXiyt
Pmau+EY1USvt/FcJfhr+K3jyOOY3m+YnO+tN1rXTm9AGyt67pY2ahMKIZC+U0Emn
Pk4nKcu62IV2Gcx2iaq/5CZkM1faJN8Dd9e1y7pr3U3B3zlcIYfFwA03ewy/fSQi
dVzV/gugprPrwfeTeR+PBauTpqL9TR0G3ZG1CcRxOtijjHenyhl4uQVRkp1KomWd
WzTx8ec6BKKVcJ9rJytI6eqRFOUyPWHlaXZsKahdEO3ZpKE7ZkdluzxMwVpRdVJS
OZ9V6w2LlegS/Z/hU8XHliv7BgSSqmt1g26bQbRTX+kWu+PexBdApaJt/LdGVX6+
yHiEfb5BM3CGX58IkG1wXn3F0c603UDiVERBcbioahPmbxkb1hieVNqPEPj8jk3p
BKo6aXCwd5iqXp2S1EZElY7tuC4NCpfFhYOzh/RFlpkCEoxvISxlOcjvQVCSZuH3
Xzu+9B3Zdoa5AJe6GTiZxEe+vMr1HqTAmqMp4PVsnZCc+B+3jLw80E70sBX7kpYY
48AbJR9sQtXEcOPp9HMPuOabwozOSFtkGmm4AU36p719gFtCUnttXyBm+2+9qEQc
NoqMdBQBWvOxYJMMSZUqOwI77PZYm7aXdsFQm3YuonSV3bpf+GtVe0iXz+4KYhCz
UKv2UgQvMnfnpSG+4mGMgbfTFeaFq3GE7PzestIGl+S00+zBV+60irFChpyJ8+71
W7APiZysh3sYCjuXaiLpaCdThWmBM9F5+zs/swvMpaK9spn9zHklCwC+nzd5w534
VHgUInBwYNkyIiMn4cb3qlV1CEOerQZibpC7F4OqOt0LR/OgtPkKe0e0HPKFPnOS
KOsubkdd0V7dZCMsI7CUNDeYJDe1pYOhcYCd/P5QwmsoIaDK0Z4URsR6zS1N6iiN
rDv1KyJKJo+DOMA3YNJQEDmt6LvgIAHmXYuPC0K9YOpD6RHmBwW98xgUETv8cA25
nimbtxyhcob0/SP1tcnOQ3XRh1pDO8YZO1u8K+elYFh6KLDGaKP47G7eradCfzO7
9lvdZU2W/X8M8BxZxlB2qq+/NiVYhV1vo+DZLk48NNYMkRcRTBXGrRNbMHXBJciF
Lj4Yx39U82t1DAUg+vAmF3kgeWx3i+ePte+EsEtNAN1ioijfaHYy8nORYFYHX9zv
VdQ02FwT3CwsZysy1V0yah3TrEisVQXbFn0ks5SN3ly9HOgQuLamaFIpRNMREEc1
vJCD1HRD2xiMVm0aWbEMqne/UXe3CgZgpLNE4+3tsaX3Zo2FM8Kv65sr2ZiVfAH7
BjpGl1VhVAkBTV7Ib4vLxuPF0RLZ9ZzEXx9sSA4AzmcR3ZRs1/Fnt7cyj9fEoA1D
ijQan2cTnZlVvmOrRUoMwBHINaMnYulECwRG/TwEgcbgqetioN1A8MYENKT4vfZI
Nm18GFDOAdbBAPsK8D5kpk+Ci72XCeCzkTluFOoQEBDf1EfviEPhbwPuDk/zdLDo
6ACu5/ve3gM3O5N3x1GOv85ytpR2Z81reraFx3i/lpiJc/R2RyMsONR8v70hhZww
6/Q3AhX9fRl1DvkavQVD4INLI0jTp5Cn6507umXApP5MuN7BpgbNWuNVhWPGo/k8
tJh+2DgxwtcfQR519iY8Lyel+Br+6W2pxFwok311V1yYDcxBL7XggQEMVsGxZY5f
k05nZV5Art6JsEa8LttxbRIrqdJFPOL52mYrPQEP0ScPsnGDU42GPvsu5aa4XrOi
RBI/79/0AgMLpHhcuniJsKaeu35YMooERcWGq0etpTg/f7f4ewjfUZgQ2meBc/iQ
t/vWeQ1TbShZDi9MKOoTBXCDjmQjQgPd8PaydCakVEGK9Gtp56NE1gtBT+6Ap1Zn
r1OAPNM8TaDyJ5/gtOAAgQUMzJR9UYAFXEKdqUGuACJWMoPqqi48UgurmfF6a3WI
OePi7BO+gD6dxJXvDQWR8Zlyjr+sOMqPBKWDmVWeTDaaHfsyr+tgwq7CPw8gAD/z
osULGaDU/KmRDszctgEwKnJzrjnP7JZvCKqE4BE16I+iKhsAc5ZvsffBCXlskCRz
TcQ5A9lJUjpS5FkjFuivmKCx5pIIMPE/yJw88O2vg3ry/wpyv/Kgxz0n+viHB+AH
EbE9yKtbLrRLuFpt5rr1z/nvUdejvYhDy4uyMB+hiAzCViiEZKXrx76iDtiD4Rll
ReCsILDqcy4YSH+4JoKefiaGYBIkHu/kKt1/vrmW+rVUIgq/2/hSqVF9kNcwkMrs
etE42hs8lKvea5b5yz8rKrf2OokdAGE8L7hR0WuHnFfW3irAkNLYkutrvG3F+NPm
7yrmlwgvptG0+uzjQUI4f1KHy46oNe+ZHhaf3HQo01Y7Nc4ulWIjqGJQ3axvR+4K
8MlhhYI7QVEjj+7p/mVv1a7emo3I6V36rsO8+k88HqOQtkOdntk3m96/6NgYK/D8
L5u0FdTHL1g53plyu75wZN7QJarZ+RKxFLaYkwKFkkGn/BczrjfcfL4TMvt/9scS
UIwOcN/7DdOmpYEt1AY7erXonPXpYg3LVEtienI1n/9yo8QijtCa1eUDtGWWl9qK
sD8kgkABn4wUzY1Fx+kBYc/+rD5uxrlpFAXUTiTHWvLYHUgG76u12x2lwAxleL4D
5b3jGYD/hSWvN+ruUhW3AARkPYMbbn20VlXgqUGLA6SjaozDIm1LNwoVPMBk8KGe
p9L3aJ5vPzNzZN3Rx5ymFKF7GIy3ujXhrWc+vugVD240QuBjr8lI8gHr2aPOB147
gMCAOVIuaRZ5Ab4f3sXiS9HWkahxDR4PQstytpYwCmfJXEX2+7TXPM/SFSEcWzpQ
1RuE4YXdpIg2xr/auytd7IiXtGxB+3CjiD7fomvBdlUma4C79q4T7+nseoV+zrtn
w+oMUbo0yYDjcqfke0JVUUHV41uWZebj3J+NO3UYMhdBd3OH815lxtKrX1FDGMkq
fogb002CF2a6wSXKCcjnPhfy+ChA+rslMah9xqrqjW8hTdDBWiLVLtbcIWuQe+hR
4VkHPvJJnsDLDhaCKSn3vww/5QBYhIVNcrrt8SPOmCZ2JwrUvkhFM29MNxAxX+Au
FGgZusK29cClo1jfRJLPHh6X9Rrk7C+f4KioXoeEA+P1To7CDG+CFvNdc265csUK
XpUNsDtwaJEA5Im6gDtfDQW5PHwYXds5v1lQqd9J1OobMs8OZ4tZB2I9zseWtN/x
+YtPtM+7esGW94G3jjmSz5lCr4rLSM/0zRMXF7kuDiOJqLQA+C3HIcHrqjO4vwFG
HDnyK+FpmxR5a/fGZJAmis+6Uf4BSX/j3dI6GYXTLvcfK244ePTszzAKZtuvtA/R
homm6ZiwfSEZ+wqSdDsCJavYetzEmDkHASKyJTODZaP+qerREridqdrqkTDN2FrH
0nYDIdW+UHKQsxdjr7RVY3Ah657ixzLICcOwg9Ts54vjgAqvJ59rd0g8QvoTABl5
JPk9FOsulUPDB3wLLkSnsPnTM4mAC0DQljEvS1xeR+rjev03NQaGufAZtNVT7hIg
87mdYQ5pkMSOG8uV1p0b0saqmtghwHhuVGLOEgm8mtcjTkBDyULugXyknK0w6VEf
9v3P7RiAoShO9C50TeLIYFhILQyWymGdlGZPDsx2dxjRzCewWhdgU5jzguUuJjLv
VEDaSFMo+KCvZab1Ec/mr1MJS65yRIND9v3LJQGkP0LaYXJkt4E0YhxLUmeVRU9U
F9MdFqt1lYVD9Y+ebmyA5v+cJ65Ln5nGsWMSkYb1B3IitBvU9MaHQBD2feEzC/ba
xUcUbldV+wr7Pfa3oNWFz+++NGc48hEAwha04k9FN1GxVJZF0DVGC0R8gmQmEKzW
8elxQut3Rd9xq6T20NWpGUOszbENMB/LnOas5YlFzuQN0ubY+ruX81EZAD40mnuo
Ma+0fSd2aXVM6EDgIm8mbd91OBBFHLCw8jW3IHnmNhvWDB6HnynG3dQ6l/AspSbV
bZBoOBGa2bsJOz/tqS7Gw1zj73v4TeS0KHQ42o4r2ZYiiCXPKFcqhW1U/0pFTPln
Mh7WWx7thx8Xrgijwb+gtZBtzvv+W5qvxQ3xsMe+0sVxE3GAkTnVyIk/L0EvA4z7
e5eYa46eVHy/aKZIcf1hAl06SYTFVxDetmq1QrhcTp6tZSLfJ3ohr7CtuwNMowsN
967WpLyFsy1lClSTxh55BMSuIx7fKT6VGM7BZ70DNPfjyosLjCbWl0YGRI+hYgFb
aujA5xMPs9Pm2tN8itz5Sx/8hMNcKYnL6lU605jRgKvas31vOFlExMquvZGiaLgB
+E3ANNDFSpdsRjeMeWofsJk0SiizMb4cCfN0cdcdyq70TNQF5qZE0wFhWmjLLIgn
Ze2CicZ8gkd3DVl7ETcq6IgaGZhoUGCkNsedb6IUXLZQZnXe9sUlY4hfKoMb4Gk1
sI7AxPlcyzAWtIIu/bIvx3vHzMCpU/bfFflglEFv+KCbDbnNHaBN4b0coAXHtjlq
86Jj11j8C8OrwIAQH5A+4QOjVhLUYQqn3nEMemRnK94Y2SD+9/VAOK5rix2rbnYd
85ByBnsV1zSB7KCDHtDyHSU4XPITcvz1ZSJnuZxY1+N+GOIAbed+zu1jN/EOGyqJ
kASDS+7E7fSyU1m3eu67KaUkWWhQ5G6eW5+TnuQGw+fzpxFJhufCsSkKTkWW5ORf
pew++Kxr6Ftj899NwcnwHVNXKy6jaOCZLWDhaLYvhQzGsZ4uSdRhu8cZUd4kQGAf
Warj1pLRkZhLWPx7YSdibHuVHXUh0b3hYLzAO4OTGjjCirj7a4m4AgfEeeOcwS/2
2z8hQBy1JXwo7q+iZYRb0dTFLsrNSHXAHaiLrI0mHPBIj2RXUgGeZNBFMokauFBs
uCjq89xlEeQsZCHY4wolr8oVr4q+xRXsxD+mHMIZ9zpy7cXiGTUyl1sL6uvWYIpa
jphsI22njU5lD4sx3069jGBdu12s5C1QlYGx5McCUtYu5+7VlEFK9I3NxFBOWZHJ
X+2Xps4Dy/TCfxUPtJMqPRyrLNrzCP/zhL3mluGTCPlPrYWK+29qRKcX1QT+hGcH
JsE282uu0LZma2sD1aZS8KlvS7wfGXy3J+i0xTTHgZ1AhDUYYMdd4FLcUNWnbeOY
WfEHzFW/yIsN5YjZoieQXfSLqRbxD+lXJW4pocfe5H2sbFcC+f4znwxjXqTS0SWZ
FLT4Uls5Di6ouGgIPiaanwcedue+isN0NP9AFMSscB3A7s/nrOTZA19ctB55D25p
aQw3Uhn+7/sAyyi+wfM+iXQq1vDx2suw7q+KvWtXNmCN6Z2q9wAR6gtATXKMm9HW
S9A4l7Uui+srIUyZAHnkb7VB9pUt6e/DyuK9fsadXd0ziv8a4Wya5cnJpIn3eG9Y
f92sOrTXhMpNnBBKxgw6ADOiPDreqL3kzwHC/Es66w7XaO8wyQQHEnxd5LdvwJW8
91/r2IIqa2YsWIfEK5gOFtDbyO3Wop93zXdNXf2aiy9rVqwuiNV0Gf+cO8t3v6oI
hO9+ke9G09Y8ifiTaMXo5y7ORvt84taiSQ7ioLhdImmhtTthEfXkcgJL2cHSsZ/T
o8Kxs/gn5UpEWS6otC9QdRRLVMz/aa8CaSvLHLAWjoQbrBzIb4QCXt6dk/dIhwhr
rPQnAz8tSCLxnYaomLXbL1aluZEdBulgFj0bQfJLz1r9niL/5hk3egLDR1Aeoq7M
8BpPzYuWQrjHtdJymxLeg3TXDdY/hxcjg5M9k5xNxSKWJwxYaMIKWzPirHs9Q9X2
kt6saXzTnLge9FdPjbSrrfyJlxpatng8bQXDLLnoGTiYRgWxPXMo/FNPJcZ8D7Js
gA4MDljId+U8nxNqT3I7HVop5BoW+a4x+W+d3tZ17eF9RoAtfBpDf0U5LXV8pySl
rkTiwq2cD2VhdjIhcAG34FKFcu1j7ghsVc6J+QbLOa+UQZ4TcNl/Fn2mKHgjBQJX
obCNYQGakIUujvVV0bznXtLCzd+/rH8IAxrj5KmcG2qb8LN8h72ZLCgmUoG7/VbF
jrSQSc68SpD/S5lYMG8kW/mgSiDhs5iUf17tWXQw1q145vOdKR64G3yVS6MHePZh
qRunpo/hIGwadS1S/C4nTQ6NE+L3LZZ0lJADcoqjD6Mk02/jnS1GfN4H2yzkAlT2
6UoFuzGdzFoNh9M8/aPNzKyQGRuVCWNtnYEZMRa7ebPhIVjQFTA9GUODrS6hxMW8
7DtWk11K8uklqmF7+zPWGsb/7yNsPJWc8SXl1NNyucETGdsIWiTydFsSkAmiXjqZ
CUr6yDFFQS7htWIwAz4Eo/AEefJ5BLU3kHPtx9lA8HTEfJB9bzO2Krkt99U70jMC
xNbeGBttE2ltajjnD+TtQCAPDDbcpAfqFJxbbvs1rYUtG6L5OCxQ2GmIqu7kKmHk
qEY2puSRdL0Dhr2rAirtcDUDMBw7FxBcwouxNUqdIt/bHJgUmHhf9i3TZaiTWNx+
LH/+1limPfpyHudx4+AbkCDmtr2V0V8P/67/6YTehYqqVZYfjSUh8pYm87k4ujwl
h8qlRUZVbbAuNcwOVR2oyXRKlRGA+MAcEn2PvYoMayIKCEvnjZHxG3SBSr9TK6kE
1Pch8Y1MEzxA7x9zEeEKl3HjvkZIQ8GMmhoV3a9/U18XO6j+vD2b7RKYigblp+ox
gzX4MNYIrsnjRBu+4N2quGiqhJo6LRYdgB22h/3SrY9K1UtKr3D3pwO5KpXjDP6q
Q02fcfjy/tM6dng1ZFzUssOoTOerNl0nbPZmBK23qhsoJVs55+v6G7Ic2wxRfRQg
fk3d6XJw02MUz/9fsCKAtrTNUKyLYWYMKe3SASSWt0J3ygzam1QZYARM0jZ3ZeMl
Csejyr3ioUChcUw6Q71pBiE2oacA07G920Z3JBwZmGi676RCw3nnQ6TJRwRV23eH
9K2iWAqpZDvANqzxfE3wxFwRM5GFrofmLMOXpj3O0NPN/F2GVAmJ+1lSRI4j+aKJ
kOiYUT89OagYn+B9q1xHM4Yy+3lafakVdQX18YmTLDQSeHhj7JZtRz1jgb5yNmvU
8Jo0gtCxEVRCR8oAU5L/Jvm6pS7K638FXBONNAVbzKVCj5UDF15zgqh2iboh1s/f
B75z5xsFGBnllc9w849vgi1VS1RaFIhs1BWnkUmc5kXkUPjXDqqgK5h358gYNKuP
0mk0uJguJUXRZ+V02lpqZH3WzZHzLxvCb/U1gr0z1eigP28nYrpQ7pQr40wjD9Q6
pJM0HEtIbK09tlQoE74mUdQoe9efYPwQDPXsvcfW+MPBnZ4uffSzPmHfI5Alv9HC
Tybkss4in5kp5YogyHXa9WrrjaxRTvIioAnOQB4wHONjo5HuR7uL0GOfbC5Ap6iC
aDJ3+a/AtIKBy8wmz/VgaR5lRfTj7uklX/LnOqq5ZbQ+C1+uajrDRPkVmvloOtnV
lbkceffc1e9PrCUse7hqIEkTdG+qn1euwH4edwSN9xmGdkxTCnhksfCPjlJn2qwU
8rXHgYgK79+PGYkY+gAXtTJCw77cPDI6aB8OI85C5YwdDEWpk3px7kGvdVVI7pLO
LWKWp6Yi6wIwPyDXcXIBqt9RFu0EegySoVturofVv4f1cqFFjNFMidI02H/u9xeJ
VHRdI3Y7vtgeePsmp7DfkPvsbYACJdxXMSr2ecz85kFvReomD92VZ1iCF2bv6fgc
hy8PaO/FzwHE6vZ6pu+CYUfO+QuIEF+36SXscQZgrWhfc+B2FEhVVGBnSwVqiltX
41lxBbhLfnHdV5aluoauljLuxtBO2KYuB5hHKwCqteActiLabHDm6BPYcCIV/Rd0
m0+yV7Rwt0E+Fw2QXPYNK9qiTRWzqwizEDfNhghCq6LMzYJ5jbAedYKe1965Qp7T
GVgDacAaj6Z3wBp0zmkLec+CaVvyHcuS4B+adeC5ZXnQazdhRWjjkOCtBe7GdWUa
fy7tI3/OYTVQ1k1Ha2Y6lAw4gTEz990GBnJ3Q5W4dNOgdaLXGAhAx+H8kNRR60ai
gv1fycOcSBRTbFSAsODl82TEYJeCThnS/Cs9urJExLqhxqXdDOi6QKCfVoFNpCcx
ORgvVQwUJfYmFUHsO9GemRZIvd/7Aj2MItWBC+lcAZ1AQ7tRasK8AJljwp2zR+F0
htMPNRX0kuO5ebZHMpMxg7WNZCbz5q4iikVWfbRQdeF8+K/E4kKwJGmr5DFbfVLE
/eDZ1dN9nToYyLuyDXZZgW2TWB3/Hwb/htrvt5VzUQfnKYCz4NGMobZXFpFvhlwG
dO/4OUehJEVXwPiYsExg8oexL9oOYNkmV5cfGG5R0RLzFXA04qqYCDVHumwtn+gz
d1FIzCd5eDph1MH96mBqCAMGxknWpOZ80oGPPzZmfUEHCzW5lMvS07ghWU8m7FRA
wR2K7QRmApwAyOB7NxCShdy9TeIX4/I8oz7VO1iFfImMRaWQKRamSmC/VJKBumzG
eQQ8uEmDJPKA/q/YzVWG6BsurZ864RGGI9gUSlwmnT/NdbwgBvZp/oLIgzvdVRWj
rQoQfNN5M1S8DWD1pw+APKuUHka+AuOQIAhNWWGspaPCTrwgnC1XnDjRMHZFjCwD
G0n0HrmiRJWX6UU0l4vT2+xtXiftdMuKZj9vhIjb3FUJPYsDMXCow+sbIGNOs8CP
OpBGnt5fyn2qTKrmigh33TA9MWFfjy+ZGPU6yOkqfexHmi9MoVbTUZrAUkdN+BW+
EW5lkmNyuHeWDIO1ie0dIYuCRwg1r1vUqnzY314UQAAzm2yTYsz2bL4yzCgjk7Sc
lvkGD5sAZs/8W0zgoWTPxVKvHpLUqocRi+RBQlT70hCLF3X5WKfylLSZWl6Nu+vN
dSiluKf+MfKQOtveo9WNCZPZVJS3R/R9ej4hptAq+49amDnGiwnJ9bkn2qepKj0w
9Q4QMQMwa66RDqNMexhlDAI6tYhm4hSVsuX5hXUkRNweE9LOp1VJfvIS5Xq0NKAw
PfbH+ZR3/0J/xiAvaq16YVJQModv6s9Dw96CZe9NfwR7m7Vx70BUuYuiW2y/eal3
57GTCzAHXHk4/w02lFNtbF3pHuw1fVtreetX9j2fUOW+JhzyaC0v6JZyBFcuNqkh
rXvVvhbXibUSAPCCDjcDoWZFpkdZSU1bOpPLrRCj4jTBgUfWhE3AbgqV4D2i6mUJ
wTJonSiSu6VzN3Hz7AtMu6ry+pIui9xHNtpl4Iq1Aw95H80QyRrkwfmuBPyE+NdV
3US8Va0A8yIK1DB3D/OM6hoh5f0i/2yqQUSxmGMlc7RCZxApCgSHVwHAlYa9m4us
0LUKy7l8bbJEU+cnPWt4LRUxJJXZc677k+YQocl6wMzAql+DeCJ8NBDhJKjWm0Rb
jrQr9GVN0VgzT8AqxzbkymfqgWYaAyZpTPfwmyAY2RQAl78KZsxv57fmnNotx0rI
ZWCGx/vrflVheA1XD1ado4LVU2GHBjo/yr1dAUg/Hd37qDqjoa60oqKblQ2VaFj/
EE8WMvsQSKQl6HV5Mel3I/UmZPw7acowFSiiCd9uVyYa+/Go4elri+sW2mxOvDwp
/za+hWmhWv08WXZ5wO47AaMBwvQ4+X5ZSB0Mlkh8MeAkNtAe7s1IXZ2gBXkSOv0Z
i2NX/whvyEFyVsSX06f+Ka/Jm4uPdY5iYROVnSi6CaveeO1A3rSH11HPu6DrApij
1rfsIRLpDjunOUC6mGFa23U01Sfusqi30SGXLpyoZ4MsibwGrR6HBEVglaCYgkGD
EoWVs8LaoKyE/m6gdf631x+iY/phdHbgwhT7UHGGeC0UWNpKwJeHK9/S/KUkPFCO
hIZtzJT1r+VndpO9NmBJagnywe4S5+g0tT1ENcGdhyoHMXFY1O4MWH/kCJLlfKp2
HxOKDCCfkKOjirvQJhTeCe2Ajf9mJ/3ukTNovWSMDmy7c1p3P6SxqV23Eq4d7jew
o3MKhP4ZTjeUWB6uMQ4XmFaCbrEOuIiR8V5PkhwvVKlbDnWKSuFUFtRIypl8AuvY
UByWhJLQOsmXbiwtftwuS5T4t0QGD6L5aHYDMIHVoTi+0+CgX1ugrCs8QXJhF79P
3hJmNHllwUL/MkuyRGhCQFxIBkCpK1cZdf+XArPyQcbiLOFv1snnoE2Sh8dlKqTE
9MBdxvDGTMuBqz2yJrT53lqFIROafuR1IZ8DEyQ6IHzb/hGpgegMHBU/lDzkD8nJ
PMVre3+/HrUwtPAvC7j+eoH/erWWfUle1zE4YAg4t9KGcbcBMJjTqta6TUPbNrzQ
IsU4wLtW/TA+OhaRKd7myLL5HMiLO5GSCVd6Tl4VfkwNmclomkle14aMC55+z5aZ
SDgRHpAllcEJn93I1wanTC+nupt/rHUWSiayQ28DPtE54ShhUwlNFJEC7tdowIaH
a7XigYkoF+KBrx0QmiN4fWW81ws75/DlFWSxmbC5phFmGbjVMyA4oBZP+lyle6XN
+QT2g/1ZXePJVvaevkiXmliNSM3jxuN7339QmU9hOf0xdSSFsDBNbuq/r/zQW9/d
Wbp4fEUjes/OXekkPBiZ5xc1k6HHcqVjQZqVXlClBIKIwUKZYVlDBeo4pbQhNGRk
BcBh0uLfK4Vkx8DdJ5BmLCYxNIDTmixFWboH+HN0ok621/3zja51zRUuD4NMxA84
1rPJQ44D1DS/SAhUDe4XA2+FYrSN0qNDKpnIfMNg91fRNlqgpl56wwktuFA6EkzA
gJZqgzz+KAnkY7ZvDUPOdvZ7UvnMA3y9m+7Ss3NkpuqYS15sa4yGQ28cc5RMx2QC
PO0tRdamCC+qMrinmXoRq1pf7ClT7S43sXwxO3ZRMdOH5zwO7FPu/KLXXiv0sHE6
nIiPTdfRF1ArtEYt7pM99gWcXxQ3/82fjk+myZ6RA1/FiUL3Cb+EV9i3SYk5KVR+
DXdF9XGtUuVtDUcobp/tvDhbo9fJw+vft0IO+bqnIwR3TZOH07m9DZUzy25WC1Fo
PKsq6ttXs4NS0vmliQo5YQOSF+Lg/1tfVJt7zxMJ6oqAQm8wa7bL9IRaAI6d57sV
tJZAZ65WOxP1JSUbyfaxJq4+01g2+7TNiFc+iVn8Tt0p1VuMbLO9j8a8p//XyZPx
y8q8jq2IiOfOtTGGh9B9pOq+9maG+0PREgLXVaHe8QQKJKlDxQ0gZgpyo4uoo+mh
cUKqyQhd8ptmDMpJu9VN8iRdgOpWpGWAjyMbJJUrqA/w8rtz3oA0ymXNKfElltA6
oVBKsppqzf5zWYkauQ8tcR1WXhfD4sZ1WFHIjW4rK5KucOZbElIHyzQSqKFT9O+f
FKenYuFPmIBtlnCHEgI4pr9lUHWNKftcQ8nG1ozrLSnhXZJlA2+XK1Ut64P7kt43
daHDFF7yyQNDp/VozPO0FX6EwghOuoXDASX9uWQH3beRKppDa1Th8O/9hH+TvQuU
jfcujpbLsojaI3LF/BGPQkWzJpbZMETL1ZPQxBlw3lyzxuc9J3qqNRuTJT/P6Jkn
lIKhNkdUwhs0D60pLNF45yuspNtKnKEkH7g7ivFGDbQO1Ejt3v4Pih/7ff+l2CXm
d8bKK7RbKvkTLBPlnIgsv/CpMoyqEHSluu6hK5MqUjBYgJlcm/YC2ZS9mHKm4ksb
jLeoR1v46Y7eKzThlnDSTcl9z+q9krh1WVfJsEbl0QMrBwygTOrGWZEo1PliMrf9
SPR8Q4vcbGGIICYGmm/VdrAl4rOs+NnFctT3euvWJqd8YsNczge9Zat/vrmJ18Bl
jJdd36ZmfF9r+zqPoKjVaEmeajpyobNwSLv8rXObmgTLpRgYyroyCL3N2LGfGOUY
bh2OH5PD3oqxMPh6dqIPntcl4f1FFP+ryNrv+i1ebip0Z5fcAyReplWkRbIZCXu7
fr0OlvdAZCMX3UrRWmgLfNa7WB1cJUHj35Nt/udW1FK6cqJuEsQlRfmhhhp5K/CU
WfvtcAxqQpAX1raJhuQ4FbAx8nC95IXwJiVwuizQiUnkoSkpWw4n2AoySxPgkJmn
FfvluwfdxR/vdZw5344p7jXV1yw+v33rF2SQSBtVhjM8yE0cG3RpZNQpcCNrWfMQ
/i48CRDoIjYt3TqsWorfmyhPpEIXe1fd7HgJ4cMyImvke4JnVWRHkHU4bkhk3zCD
9orwU8Mc+fePv/iI3mBi15cDs1Oc0bU8DU64zqDPH18uasZ4o+hDiKZXDYWdLNRe
IHziix7TEh7Cdi7M7OdSfso8YqCzuS6mj0jnuFKyZN90lF9tuQFjwu2YlwC5a8IE
2wQrO/srohdGigzbCBI9hT0rC1O9pgN0IAkbBw6L2lQgMJQAPqQYNqO9IXaDAGQU
Ifqd6/DlhAUHonzmZm+tKCeUW+LkkcLQwK+au4h02Y7z2wYnvelhgcf/hf/0CZNS
quN5cKwQ9Vk/8lmbJsCgBsHsZzReJ9+Cr4/ftmSB5UxRsRQfs1vLGbEc4Hjj2oX9
odZQhHwW4P8hZfra7sgAaxGpqkhrImdM9+1neCwkXzMkv26QOncKYUsra01iMbQ2
UFZLbrL37ig2OJ5v0eBxBezJgVQYH8S8mtaQlsOsNcqL0QRrLLM7cmwEbC15dY+w
fp/rCTd6wIYx97diGRtMu6dzIlqCkfseAxD7HaxcA7QK8/QgqcxSc5+Mw2T0W08u
RA4ly+ZLuvUU3o7J89g9NMHtbfYBVmwd4H5MTbG+n7xGueZKSvUQUbeDs0MxiGrH
fxJ6jjb6S1hOTdK3NK9aWtslDaCCUNu9+tLuaYI7FLHiJTkRgCpOVCc+a1eFDBWc
bB1mmBrZocCy06QKqyNxrB183sUZuE8R7aUubndtwcWcfGV0w8eKjOq6J2OOAxrp
29neT8xaZCTvn2a/MGfqtOMg0A3LJ9EYxxAQ0oQ1IeFGMfaLiD+YFX5j1G1ZqN2E
iPwixb2MfcDEuRLb5nQu3EhpqTlK2FfaPadwC/7GTvyY8/FlcDie9HmzlVJfmuNG
fqJSOj2xmQaMKDuAkP3YKKRKsglRcjovDHrXVh5GINI7FvmypX+vUQv4IAbcVJWB
yYoQ6lqJ/ZTT+1edBk6XZIZhp4NfjIcP7n5HbkO45ng+CNxZRHCr/XP88LfKwwIs
qGWM3OhOuWmT09pIwCyt/kjKuRLjJCMXhYrbkK/sj0heRifFrkB5kK4mTCeSdB8f
2q/vfRUAoX25eleLWLY/ShRjnPqdpFeQOpRAU9t3FcAfJOw2cAiaWyHl7xw88Wub
ArmWFCnsepAY0lKchVnulFVD2VgMhwlUl0VHZj/3WXn589Oqjx0CMmCTLbArGedO
ZhJZ1rsv074XcTkdkoI0LsRTEpkyBmWh1HZjwVdn/gTdi58mL3x1cv+//dl7bA40
F0WJQXBJvNlB7yDjLizcyOmj1RyF9V2cw71arXJXqyqm39UofZHwYacs2YezHaJ4
U9f/hEbsg91T3PWcYQoremqaMdeIHt1BJZutnQKqm5e6MXm1iOLeu2T3lLM+WvuL
5yKTGO1DpAPT40SButL7cOTYX1O5rhan6+nDVBaMvwjm72I4sbpPMDcNSYFTahhH
dAcidiSOAdPCk+HK07E0lvuNfCCkAgtIXJbsKi4jkzawwSVG1xatw0b/2nGUIuaG
wrMQFbaXDnPBdmDw88kwurluqJ0pgdZiF4Jl+s4QyiFQGnzfB0MDqdCHw9+AJdDB
EbNdg5lNiz8IyrKZD5ATY2k9rZQPqco6k08Uy9poauahZgvPkGvcUDtY76EUNKsu
RmFevZ5luplJafS74bK7apKaVB6gxmIWXkv6nnNmtIQmbUD9ApIY4i2BXlQPZX45
bfJtK52ACSl0hKZwYIofhvScoj90Ij3RYEch35UDfL4xrwMQN5TWsgwCipAg2lIh
dfhdO4l1bmwivLenuwe2YMxDr92NGi0Y7hMAgpugDwoExfg5zjeIGXkE2+Reu7H9
ICEu6hFaJ2hpS+5adWzZ/J1JpZqzAHpn39It1/XY4GzzbK6Et4y9tgOuMvLwsyr5
frmwL2CBCO4oUc4sgtV+2DAivNSVL3zJY6+mkMWiueEZo5+EaRtHsA8PiC+GSzv0
toO/KyoM+Qs/2FuXETdzF/LI8/hGJwIoz5ElmZBG/o0Ht7B3b/yz8lFYZCT6o5sA
kyqg0w6FcTadl0qnNxsvspuV7fRwVVCysDpFHvGsZ4Gi4ZlTefKz/63KqM7f8cjb
tx0CH3rxvfyx+1zawgssiSmybI5GkIsC5Jhikb0+EwW/DnU+Nv3YimCiuHhJUwXx
JHU5h7ckA4dZcxNOQ+gijYE6PAf48nPiT5tY2e0uRlxcbqLVdXR3tBBYsUEa7n7o
LI9Hxo44VxsBA4HSPnihH2uoGnaaaM84looekAw9FymKmf2Lbz3PKY/4oqMpZoUD
/zrHBzpOfPZyNJjdabjg7gg9CuaFfzmUi3Hj58mFP6Rwt3vv4kpuBLtotFPpXWIv
tkv6zmccQ0boQArEaCZU7LcCIhX62LVs0EpHthrxIbsekfidLT65TIKPgQC6zsea
R567yETMgmDp4uyvCNcQrPwAPCRgYelMqg1KMF94Hy7ipIcohAgyRCxR6JtBYNeF
HD/ez/6VuaOxT9KMWhHohfcgdsK4cTzu5T8HdQdCwmeXgUttzxb52lTb4gLOpbFZ
7uLDtogH+6TQdpoJKQlSsR8NVfgeDnhrYuy+V6aET5R92VWW9ROVT9tsTDmXp7D2
Pcu0vgX9pQhJBBsDm/v7WWbeN6YuFh2tkr2435k28TPcYxATZ9HMSs/CbV2O7eGM
gy2+OiB9qS14JS5t7y8grOZALcTZC4dhjgmSYKjv5LzVz9yEjva8mOPfVlMetOzK
MpsKZoLP9csLhvPKT/hqzGq72LqO6gbS+B6BBwbrernsfgEf0itjzrn4RYHvZSUB
9ylBRxP04mRG8bS3imjxbMoNSohMWBtOPdc+rS/PxiQ0PhGLw4IoaziAjwzn4TFe
6X2zBvfc/z/9WiwMMJSToEPmiI6HeDsTrqIBtD/zvQSj7+Ik+FREEYZGGy5361Zr
NBiIF2K7jsBpeDmPbFoVgYX/lLu1+yNbxNa8wQ/LPOyRupRSOQ17wgYlnOnTJRjn
iwzr0T+pghDfrs0l8UNowtGGyYa1vkSdWJofhMRNCmMvzjsJiKO1wBLaSwkp8Xgf
7u8/VLx2n0Twk5Jty1kPc4NY8ereD0zZvYVeLSgPlMTuxJyE/hJFSyG0Zo46QKR6
pkIIUoY6ugoI3X9NmGsOW2A6ccBDLOEgdUZHQZiU1tzQ+rCbq9DzFNbND6bPcoJV
g/7T0rVVcdz2KDn5ZT4V7p570elwx0IybffvQZEgNCcrgYomTiQDpYpiA4NhvtDw
vKFXZ0UgM9GtOQnKB6ZA7haOHs+dOsEqmy4+VN5IyFhFtPrvSWe4F0kK8zxrxUCM
mWErTF3brHUIJZbjTiRi9EcnX8yGu/0SJh5G2vCcy6ZHyH3OVPit1gkVRrJ/Wjnl
bErxXlrlm1vqJ+FCghR8V1Bq02U96uSg5jhycLzUOyd6KxIN04Cn869jGoSgVjbC
Bm68mSRBHN3Tyw0ULKa96paueF64m7Om2kLqp9w927E6N8BGlnA4ObBPiRbzxs/H
3qWLDkyPk7Ie4IE6ICVeThQ8Pb+LqsVokpyJ2l+CL1V4NJk6O1dNQuYaDhrXAlkD
WOGfZ+Xk69uUzvespUIL4hz+CMm8Vw1gojpNJ037S+z2eI7aL2ZAZDDOybdfV/oV
KemwptQ4jZdyMauiT4Q9HCuVIUr8wiwv51pe8fKPvorm/PjQcxDNYbX+9e5Czd6l
CVce6GZiPEG6cuexe0Wp9aF7dhEktQ+3Ux+PWZzSbsh7/gowhKymLOiHgqrCoNoa
XPr+ma77FJyClHmdX1ZOw6CMcsqfOtTslcUf6TkuF8O8CIDv2yMIRhM8uRxKx/sg
pp+t2Qj+IgVw5sijsOiKPvqT1ZpnvxzLgGSecn9UOMw6BKr9wZsFxGoYjXPTr5q/
vB2bUjlilxn55QlxD6JZiBVrkkNw7toM1A3mjyX/fVVkzW1y/drErfheTkoy+bLv
FZc5zR91yil6WAR8szXN5/rirho6S8puriq+C3nltd+UVbwDRWq1t+b7JtUL1W+Y
bU7BIUvuY6wQjWMrg+Y18Uu3Kg5VvQGm3SYz7sctBz7CPFIO+/WQhLK5IKmVGfzO
m+tv3ioEkV8Bc3kfeSxbP6fceEP2F8jHxfhgTo9L/ZCxgwbHmO8V/EurszSGAFks
hgSww9fEu2kSGyJzluKYPzI1nfFlFLHXuqZuq9bv+T4r4ibU89aqkCSckimwnCil
f/npvGTLo44M5TH8m31aYsQyusWECJhMx98/N2TDL1GjQSCYaT7XVvH3A3lLarAC
V35SnOlkZTCxmlE+m0cKHdyIaJZWLs1NWbEa9ASpee9e8ZcfV6riyd7fpmX/7upi
Q0TUkc7VUL8HAX2wWLl4T9B3batAFvkD24MBwYLVhA3ZmUrouxnJjVn34sf27lAp
/32iQwCd9JZyFiEBYrGEjp0uxAMosTuXFklmYXeSQMY6uMw5zgL0sH1R6UCfUsFT
bunKi25hT0uMZpecbTXftiEINh24LCHCeuGoE7pvBHn38Bi3pMSF/RIMUipKsFB2
c7nHPryeNTRurZLA7WF48lN4yVhbR7eBjeFGtHf99SJFEfFOiV99oiFFhN5soLHb
DUQSoQqyqYHrfm6Egsfxu1TBG8pnjuLokWTnsRAoW6fPDjkwHgMNUmij7lr5eRZr
DKFQUFWEXzC3+ta+EASBMST4s7Dm8rFVakAGbsxT86oX0hjwMc6IVX7gSqcrg08Z
89wnk8goi7Y8dS3J0mTnEQgMTaPnuTvmXVQTDbFMXmBDJ11XnKQ4B5zXfqnFMA3v
tdeUg+PYtzIvk+VokzKeV6lOZ2/bE0r+SSPiEvlYJo493xKTjj/UJJnOH+hyqMC9
RvTY+FY18EFFpY9q87r18eKwivRdrAVqBDVOOTC5P5jZUnkZ4KLkcrTOk003sp6u
LbOJ33cV+MZklTS/TsMgRrNYEuVnDmAfC7P9RK3NA0iES0vN2x2j3qBQf+rVMFdi
+ot19BM2XwoMAaRaKKUBDTwSyiQk8RhzYn8EcBwyC65KUm9EP42osxJLVCFc8yUW
3ZaxbkvYpfRrobEhetJRq9ENA754xmJmvHRQ4DVv+e8PV8Kq1YDJfZI9pZzKCuhv
eUu93zucuKWBMYfhoh6ynoE0hT+ZIUNCAeY4pWkdMZewUe5tie3wHuzGRUXT8EBE
vfOtqPeI5GMIXrbXb7EzoSchA1tNKClS+zKmMCwe7Xhk3q2lNABX458bWSN/jqdP
CAeV8pS9iwpLqAMqWRgpx7lyLDPnCjflqzadd2E95gTdvd3YfJTkl+dqolTwVBRM
1NlZVv5C5+5mUdG9WhVtnFCgpxDVuV8vvn1C+eWEHSlY3RpZn5+QKrnEcgjYKA0W
NMMXxbQKSH80nri+Y6cBdaiEgEWpmY/ZAbldnqfdQ0bxXFPVXtT8cpRBaP4IJa90
xqamRhGCGQsKAuBS7FqltNlNb63QxsPHERsUWNH2VAI5RLlepZVAAuexZhdOBQvj
3BA/fH3niub6eEGYNfC6DC5q0dMUGV28Uy+fiCG/NLWGlZa4omTNYJ3hbD+PaPBu
2C+ANHluEW1PcQgncct07UeYd0LmQFcVb0TbPskSgO9mNZY11qF5uwm/LmclHVIh
pDQEILgiaQT9HiDWI6jm/tUtrgPNc/JwAw4qq0qb/MenscC0xOdlO8cqLL1Abebl
/wD9gJhRkb2SsjCBUHNKCXQNhxIFO0tEyj399fY8715sL96taUgdDVfpfLmr8TKL
aXlSm2YyicJjyTP3uJ+YbaYB+VUkZqts6NHmmJehO/GUJ08mhYf63433XJcS4qh+
BFsMxfNrVdDUo4ZDoPsuYVgZ4wKwkIL4kbwB9y6MJZJv8MfOlEYPTvw7XX4N4KTW
+2oi54sxvaQwNzAHymWewtnTvPy4H0nlcB8+wN9eMPAyCow65sHlUwCu+Hg3x7r6
2dZHR9KLbH3SYlvdrvYxw0TPdxa8uhpAzzIARKF1Aj5g16Y5xye4t7o1XeW1priE
G/Pst4P1fGa1nfrqAgFsueCiVGgel8a/Cu427DxY7hnN60XEV1+10ihx4+zUtpPU
jdn8ggKXhu1dKNCGut34MAnQwB2CVjn6F/QWjFDtSi4oRxp8m9rsRfBm136Uvh1c
B43DqHAPNIjMuYRGKQzU7zMwdsHzagk/fiuSFoBCYk/+6tlX3u/3Oi5NcMmacQ3E
PcVCh45SynXt9R1Iwxa4e/9+/3BqITr+0i3IIBsu535AkOdY3z6f+aUxgSiSzkRO
Kv3xWI2g6Ypn9e9TeHM1ObBELLdTQbHKQwbhYSnsgv3AiOoiR6erwMbnfVNBnSGM
AP4lAjCk8UE2SxZysrQSgHMhB1A7O9nKbG3y3fg7ryDg7C7MncLVuH8LdGrcpTDP
+j54IO1zMMRM4rnOxrD+ePngLKLroZ6MquXcAO088syYCps7lEa1hdgHVVp0EFT/
Ne+kETbucoQVMeLF96g8MyeAQy6hWliRr3uoNyg55nqjxCq/oi3qlYpuq4IOPjQT
TLVHj7oPL2LpIGllu/U1RwfwaGLKoS4VKYKsJl8o9LkiIuMiCpqtZCut7lDjKRIY
ktUNjI7RJtJ8VPl+yPxYnjRuzxaw7jgoWZC5ot7IAkR1e4+ldjc4HLLIvOZGSHr+
6C0wPuqAREYG5n2slika6RSpFbhD5wv5rJE0htW7VCXFGcgev3EWUTL0RnsL2D92
4leCxs6vo2qJfA8RqL9Khlbjh/qAMmLLNlgYzG/xCzrbdZ7U1defbniLbVeHcEzB
x4gnZ26A1Cnwi/Ta9FqdW4I/l/Z5ALkFEHuBlxe5xbpkcZDknOFR7v7+/HilF6D2
VQn+ofypX5GIBiC+Yea8eDbtfRaUTExK3WAYS3LqR0vwfqWE622NUwvCCvbahL9t
wwaBuc4Sc9sKTqcTNmVXvoiTAryuIR8cCLpwMd8JMZVVO8gNv7AFqIDrDJqBf3hZ
njxNXu1fFuwDrbT6qfbSzN0kky1NubQfagob3h1oJZeReWpuCuHt8JgBf9YvCTt/
NT63OFv8sVqLIZE+R41vx8Et2uUFUkjJrOY2Dnix4eN3KUwmF1S+x5FMAQrWGlh7
j+lnr1twP9C7vTQRG3Sf/yHy9lA1w1cPgGCaQFyduu84g2Zp7HcGqORTq54xMTPe
zCNLajYLo5kqrC+tdthU2GeALXYRfkMJELpa/orgcX3nJPEdQy3vg+Q4N9ZOB+22
1nD+1qmFNkWgtS1SDBheVonv4tJpHtVnK5vPmK1/tqXOHs2LHWFyY4ZBy9M22p/6
1OH7HgX2biTc+S/1F2xpCxnStF+WLXKzBEJvDy5dbxaD1rg2aWXjxghwVFn5fWye
eEdrL7Fzb1sFeAXJuy3dRkcWwR0NftZF5zV0lYm/d4uJZD1ukbhJ06FWGZ45qNrr
LVVOPvm0fE2Sw3bj+d6K+S/8dDKdgudakghNprMecDo4yj8f8A8auXfopiqX4tsA
tbSHw02Avy8EfMeyGFOJGHchqA0S02jNIuFmhgJhL1npe7L7wNLe2JVbyGyjBjSa
Q0cJOB83ig50zbbEIQTe7v9pGoOvnMXAm9BbwI1j0FZ0ZhNZHjxKolqGpWEqOmde
VuNarUn3TrIH/LVRYZ6bsOdrVzZVWZlEcivyxlgA8Fz8892+6YfXLORUVejD2xps
Xg4naxGkCHOX50onE4y3PZ5cMmx58bUt6vACXycgl2nay+Tvz19jeB5WFNcItotL
rXo3Pe6q0FGV38r9Mx4b56NX97P2AANe11GZX3Fh3Z3AKEzN8jLZTjKKL6ihdVS9
DYVDVZYLVfHxNzL8sFVde2puJY8G2CmJm0l/5223HziFaAmbUFR+mNFADvZHH7sh
Qdy7Q+RwhObzuqRJPuAJZvJRfaVjBgrLQt0VjvpTIrPHeWiIA4jdd/45rktt/k7X
tyse+Qd7c2ktYL4RJLt+aGSw7wH/YTxeIgMqqROtmsd7SKitaPqax1m+8EE0LBrF
iQUQggrqPxBFXlZXjWymcPMb5PICQKzphalTtC8eW2GoPg5MZJkUwCr9HjO+M8Ud
u2YBp80SoT+5InHnkWgsYPjZSAiyu/XpFl0sjsgnLlZ+BH5m4N5NNdX11fkWnS22
f993ssWHSdJ/ici9qOsb7CUmweEpMxBMe/9OmO2Xw3FhAgNebK4lcadV4ynLmwLP
dykZV3ikSe/YMgyPRUraS7/2iSc5xQAuTHdrYp0MbJh5NvcyTJg9EWTX4Nnevkzx
RxAdR0tQx+k3bEymgxJeNCO4dzxKRZKXCuI4W0VvbjJC2seu//X8Q/6vS9pOle1x
4a/vL4NR+cWraKYOlU/Gdapg8UMdXgkDjgqw81xh+sfophWK8ZIDFYX/TKGJxFMS
PHMqQ6xmZY8vJEYgYqEKVeKJAnMoIP1e/wfXdqrqOsjmHbTEXNEEzPItfVqWiKbH
6v+Z9Xu1DH0STkKU1VgZS6DF2NRiZkspNw+N/DyO/kfQUU+132x2W/1qkFvs4uRd
b9KfW6GjuU/ZskeZOsa5wcM5MftnQ7JtwBfqRYCXwikD2SLhaZMTJU7DdN4JrimH
YPwbS/I6MkXZhptmMbncNnprXtHfq5NA3jPLZQgoDkWs3hULRwJ0Jlysp+oBoR3j
D7CiTep7WlUvM7MpgNoxItUy4bcYjwEUM4Ae/7ACTtcv/9RP87VyV7bo40qVxtCL
+aNXX3ZF6s7VTMrjtcLHTAfWi0GpXmY3PNH/BBCduT3Pvk7osSdQL69wUFDIF3yu
FKUg7lN8usrNYHFj5OcF5wvUJIJISm0U4Stx79TeSc2lNnmwTtudiwz2DKUv6UI0
jRKtzsnCibR0Nf/mOsahwdRfqx4OKw0YmC8WwMIoASPfEdt9YJkGFQV9LE3nxHNR
cAjblwMpqIB6++O4ct1iH8zvP6OcVipHzjedOYnhj8if6gm0ZHiauS5+GiFSD6Mf
kL4NLnociZnLrzARwOPA49nn9uLn9a7UHZPnyp4pcaIV31avyUt9dTDCTHscj1Y+
A7wm3K8dWW+RvA0zhT8UciDgtvh4I38nFoir1ZkYvQq6izBVZxDCHv23KgrGvrNU
49c02WzVe4TKDwUhnmG1sb0cgVg2nTteTVAsNLGzjXBbKbbrt336a9Izbi3WbBC5
hATtRW832etJSWUvv0wiXni8XH/bKQvbvxHMp8hOqeX9n3ecvDGtQGipaskdOKov
+/ROLtV2/umadOoDX7VAHcftq0s2B/1isG/kIP9eH6IbpcHhFuDGYoG6D9vGl7en
oxnI/oyXyN0/NvaynjWlR13pWKqGxdk38Z6e9P1ZMIGuUTzD7BC7mUBH5YSs5x8s
5oIYbkQTQd1sKlolrjAlvz5lje2cmMaTr3tGpDS9pXhI0e6jvKG+B3YVtpzq0ASg
3PE0dOjniAmapZkEQIoMsMCnOWHB51tGopd5t5vQtwH/Plqj1X/b3Jd8pMWOFlKe
qT+y9PnSehlmujcYLfXinGikw41A/LZUDeqHsxpmkWnLtUzZYVDgZUH7rqApObMP
FpyWvb2DsKVVeRX/s74EEY/951Q6MkzElN5RRx4TATRA7rDb1lRFgRIdOXswGOhT
Y2vY5pLXVVBrv2mAy0a3wuZ0IgkLqIQSpeyEwpYHT+WDg/KfYyl4dlD9SeeYQwn6
icIh58gDjyFtr41Hzo465EA5m3f1cUJDD6Fe/SvuYO1ZGHDu69K76F8tA+4bfT3J
w0TZRgqI1cKPD9XNCUGaIWpWsc2ukkwwszySGdIQwn+J/k0eN7SrvDDH++MobWUV
rA2GaENzlrGCJic52rQbR/j7Ma+TVQanGNJoBjtjE2D5/3HlQr4hNyOnV0njVKOS
UEBVYjFFuTUJheXKhRSdw81QOJkSH9zvtpPqvqLgMphzbE4VHGPm1AXLWnm03ERn
zqUxM7+0bNUrNlIchEvaQa1Js52hyjEoyplWQLFBboO7cAxfJ2IVy13wHhXuOWBg
gqgxXrb6nZ1vqA/DOmiyqSwLGWtLCi20XvheF7CYCyCr41BolzEOXgqoik+V8N4w
UrbFBSh7Kjz86qOYFKMQsDw6vkJ8eCArDdcckpVks5JSz8ODzSev4CBHlQEWavGz
5j/J3BQo3O5va/k9Mfl8yGXNbfO2rJC8Yyse5FN0rRS4RAmLVFu7nYl8VT3cvVqk
HQDYnYb/VCwF6UtagNb5J4+8TwDZd6U6g1zbxQTU+pa2Kfu2Wu22yYBGJ3U17KCT
8n8Iq2Y6ndZnvkxTaS8YIAEsnGNj1/fW6CK4ExCfxbH6FB+g95YxVZA5mcUmZVqx
/4DdFGouTzI/O0zD2C2qtumDdEMW2FaqWtQzLKa4QnWijgWMsSVeg7OybgOijwsN
LrHjcrJX/VRb7n4Sa1zhCTyjEKjgbLD5F+ubQ4riFfTKdUtdezLKmMXd41qsbGzv
48ZiZLEQkZfpQWMl3dRC9iJWN8QzwcI60v1KpITvlEKh+uv505D36aWYTVH9XWKD
eHPI0I8EbujhyIGULMHKZc1MwQw9DQVzzeh+leTQhz13TG4UjEhSybDgcOXuXOdG
pe6HpIyShhqwiCs9qlhItLMO5qG8X1dwc9LRdnV/Y0Y39IL9NN5m/6ta87gSwoOx
nyDfX7Rsumsty0RxUTvxiewwMRezqfWescfCswY6OpDrC+0gDJw5jN2D+ATREnlW
CzGd/JD4iYKVzuM+q3/StSKSpPrUlWu7GEb+1BTOIB8cU/2PeTeG4CBc4CP4gq3n
yBvUXXj4NXWjMrw9ibZBN260P0O60KJIuSTT3ywobCETka+Irk5ZFzvNGyPUknGA
Xzn8YG6RQpV7Ga0bfRO0dwOGkDBNiN17/oDQ5GktWML+EDYGjEPjDXI03WB1k4f5
dLJyidwjAip6QloC0h5kcPenZi9cWGkk0T7ftSl6eRb276Ee4hpPyE3klI5MuYC/
P/8ZN6MQtnUC4q1oZXQgd1Io1jJv2i4qOJF+aeDcLtnxVHE0TOjJlcDgaIBfrdxf
OUOPKoZvnfNZOGnqt7uXqlSmFGEbcuFy6+4tzYIFb37fM0NBNyK8RkIWbQLt5u/Y
59s6PDMdEqzR2+PGSpHtvAYZbkX22Q7jk2/tusRwu+fqQCr7fkRhRDGJcR3H7EGq
8mR1PIRUc3AKNAOw1B5frhAl48B/73uy5IqaCRznbQzkpcYaK2UUose6LggZAAII
XRMqN70qqusUf4G3rawKLxZv+VwdmIwvrKBDfauKxSwvPk4InF2mtbVbEqdRA3Sw
+w3YQ9QiGL+QL6qTDWq/mIZZ4fpaDNW4fDq+Jpyjd5yHbwKXVbBN5spjSICLlhiD
wkE3n+sJG91dMlewFJ9g3Zz4o4v07+j/VgJeGn1BmQbQneRMMn66cTK1aPGIWFXo
JupudReqzhshGsO9D6cEuB9/5ikt7xvjrp9v0SQaNj26+QT39E4w/37tTMXjIu+B
91C5+KkTWDQrfIoJs2ySn/CuMQoe+43uHPfm32dA3iNkpUlZOKvv9zoQ/6KPvDmh
3Jl/BU3bdmov806KrQ/6PiqT63w1rILg6Zy58mqavNI+77TVRXo/N2Hprm+Q1S7t
Deq4nedqXHrtUKNet7lrVtSxukDUZqME8KFn+/r3nbG2i8Tk4AWJJbWC1HDrkw8F
uLWehzkAzeX0l9IbWSZeM8FBV49jAXq1OA0lNMuAv//cFWp5k4S3p1FvH5SrWswG
5ayMBZbKGQbSdIBBBjh8+Mo35dINm/XmeV3yw+dNlBKZkNsl5mH2s6+6V6J/tTN+
zAz2M/jgveQS74FnXSDAlADWDL0wouux/R/IBs5WEzHyYQj8TC7D5Nhnbde+OVzj
1hN4+2UcZHowrRuBvZZ3D5Wh9D6bUZgLRRzEYWrC17MZnepSr1jJ/qtdwXGa0X/c
LJyv01K0aasUwedronK0LF98EmOCYhSgv+xu1t+xeobzJcLKBbwxdKSJn/wq/cb3
UMiFpEkI8gR2V7spinA8NpHi1LFC/9FhnJNmo0XJ7ZjzdDqViI5DjtSu+jzNLVkD
gG1gOjNn/Fq6i+pZx/oJIxfBMPx/lKiLk4IcH56zJ0Qs9QfIm8VoVU67mJ10UbJF
M6mCPbVLzuNok+qxIRuQErlsgQqWJrpdL/jADE4liB/BsZNeGjpxbGkyp33E87hc
NWb0zYiYhohErZ6zD0oXJzg/d2GksUfV2nEdnOMorlcMQbAYsD0b7wQhy8nVPmgW
C6XnHfUwY2qlTuAAdcN1bv7JE1vyk0ekRWpWK36gVXi+ueUg7JYRGzgSjxUjH6Hy
KXTlLAGYZXYHQVfrI4MuyLiG+svzHGos5eFQTjAYKbh/t4AolZ+SzMUpjJrtayN0
QnNSYs58ysKoaAr5vbZP91RQALwWHznnZR+cE1hq+Cj5CXW4V+0TRXQtLqNIC003
Yzd6AQT9DMYlhrD56j/H+3e/qv3P2yRqd5wDxMZjVIVFqdvSnXyXKMVkn0hkGiJZ
2gEO1I882NTFg/HCLwiuN7CIVfyFl4AzDGRBd6a8qKsB0LRW9QRnZGUqsxNqA6mC
gume6rEjBuFjnMGy/RMJ/jESlhVwNj8xa+Mfaf1TXUwJ8kyJPNue6UtEOuNb7NUQ
5AHIGCz6x8Tw0Ssl4u2JNjtbytEZAAHc3ZCVGpgH+RqNp7SNRmiJBmvrANcCJFEc
InfaBHxCv/O5hhzT3yGoQzHSjFDP7Iw0GmSgnzDaqhXJg8VOOZVjC4I0Jk3qYD75
q4SVKa1Cp8DgLY4TnSAFYt5GMIFf5bc3yUanTDGRb4AK8ozJhkeDBIcoWBpz9icj
Jv+7IJI8Y4k/R5Kg2hZzcluQS5OX9/Rpu4cohzjlKNlOvfTIPNaCsud2upkTJX0a
gq9Mq70xHp0ocdU/zp9MtoFgAE12RjQm+7VXiXK5jdvV+WRqkvD+Qx/2Ett82Y4R
CFWQNHEzqvDAmNnVyFsC6vWAC2RRIQm2yzmzycW3S2W+10Dd9ojC0OVY41wh7ZAt
kF9a+8Unmvg9PNWw6ZFas9GRMD8JiZ72XuzhVsBZuznP96Onb6+rQaa6GKsk0wYn
b+kPqc2cJlivgxEFbMElRb2Qbf3re0ZIZD6zrtsLaM1FipA84VPh1jIzTFLi5/GX
gHnk7stLv/pOIpfFeqan7Nbnx6xNm778Vvo7URYGJCgE3MgRT4u7eUqgF4bXf6e6
nPTHusv8QrJwIN5C3m+K5v8dr8l3VKPqJ8VCKwJ24s375syLCXO3hE/jrhC5gB0Y
x3yvmmxAKPe5VKrNX2DuA0xaGT7/kZ3SNhS3ptjrkWMKu2AYGjL7caE0ELLLPMDr
j1I0BFWOtgcxuNOS9rFEUqcg+8JWY9LCtgEm/OipX8tEIdYEHUJ6O/VZkmlvCG+4
3vX3AqAxNUrHJ7IgO7ZpnF2ba0U8FIBNlPQZc+VMu4bMfj3LzEJafessPV4R6ysq
XHi8rGsZ7JmOZfkf9aEvmKogZS4hTePeHQkSHljZUzkx9WVObPX/dsSptSxOntVf
I34x0NuejMCHJH7MrA27e4R1cxHNQOo7jxpbIAlM+Wh4eGYCaxtBmeIXbm5ByV5M
8yGsaZBJ0LqQGe3w3s6W10LLiLpE3HZp+UWCxbDUA6KeUKtzhXqIpco6+tYWjITy
ufy/MyEle3Z+Z9tpwKDYAHgk3e1ktfbLNhisrX3uk8DpkcGY1fQaUQrTdoR9ZcsV
H/HtCVekmmE5tkXDn/fMbJKesgKTAk6npxfNlT866jOP3nRVwP5fmo92dMPv7vo2
aJhI955F6yLDAuEgsf48PHrGV5NAodmZvcQMeV0AUmq4dYNJPVIgm2hoTan7HSkx
u5ppOep+41YEkg2J25iEO8ptcdrpuP3Xta78mObRlCM9YRUMo8gLcN8opJQdEQOE
UL0egxHTLA6yq9iVVuDcV8mcLy9fro8hLydDBMyckofJJ+KkoyursSAN0gu6WnU+
VuaSzDszJj0quECiFusBqucH+fw8BjqAjlT0R4jLVVfqNB6z9lSz/6UVB9SLMgP3
uVkCBcfcFsNz8i+6jH7TI6dmHlxWh/4KUhH5vI5sxP6Go3hnPk7kMpXDJ1gtxlyO
f5fcTYyNEgSzVzc3dBWRE/VXmKtJTWYOMzoD4vyBGnFiUVIe6gLquFVT5FS8YzKX
0u4FKQRkZElnB8Fd4dUF03y4fkn1yL9pNBOvvSdvGRy9uh8oHB6JZE47Vt1huWAL
YbUEt9aMrGbwNqQbbacPRahxDyWr6AyhqI/jcwYwHvi1VB+nPkcHoPZPoce124Gn
NLCiKUOUs7YWXaHWTo0iGZfWeH21lH+LU61hIGsdGtf9F49WqWSKjukQNkeYXAX+
eEfxtsEoCzVJ5avauXCEate1B9Butz+/DmfNKWVUZOEf3V1MWV0XV/zlnPaVc9DE
QDkwWbmP/Teldamr4PxKCtNBeviBDWIK4m27l6Z5gYpdaHYV6sd0BCEQERtPLd6P
wYxzfbmENpcNjJLG90+okqG6Eq9RBphTViaAPtXglQdLLXS+4+RyaDwLEJyQi/rf
6ESVBMo5W6S8UWIcJuMUgWWRcR5ygGos5m09n61u1uF5Oc68fM9Ic7pJCpabaH1W
PjWSRkfvaeaRIySlhx5au90FW0JNmTPVWYp4grFPzn1mhWSitsxP2rPaA9vlT+0p
/bU9bWu2k3ieNIR/4mvkV0l6hvPSFAR88Z8lM8592MZkpGNf5Ft4JIz4QWpnk4wO
kcn6LMElha8jaq7G3vOVzDqKW8WRJowlEG+sGzfN+Epb7uIgpqCHb3nv7rqzXw5x
DBeEziltS9OZnxdw4FcRXQUdjv4VQnbHfe4UFbkdfvZV/abuViAMctD0maPiSrJy
uX8Cvl/xBFo+gHgmKglZqCgsQFRR553oqbkI5F4Zia9KvP9AxxjlFNyr7FqMSp54
HX84OG+zcytnaGNU3P7QA/goAGSgc8cMmCOMJ2I9v8iMsg6GeTNQnWRnvO+t3aqR
pvNCDGTW8qSmBOFIruHoiytQN9zin8IPC48MjokZdAujfLyEQLtKd9rh6gz4ArNy
qHb15RuV2LJ3sZ9LX0t6m9RJ0gs2XXIgNIHWKlfFC8xCtiso3pHm4htBn5lDMcwT
MInU5bms5OM6OuzUlZFGPh0yXhUJkCWjOjc3VCN44SQYhqo7HmppZKmveam74G5L
gq72bw7tHX7zJqHSaB7tiiG2tHvGJ3u3XaOYVHaDo7SDAgJSIUSzF3dqLqPfhmDC
eXwDzuFuneONQ/9ECrc0kxe4i+JgUYa9mFramqpaUBWh/NlfzxV+b+RkL819TNLC
32SrDqVknGiKfDGQUDJ1RBAODntm1F+iFxdocMPtX6Xr71wTftZ6Nc/1AeZ//7IU
e+71VmjQstPqjVGvPpYqp5RoVadKza9cKOP0ncItfw+z4sou3DzWkCR1+FSQ5KLt
fi0zp7Z90p3y+oYMzWeji4gYEswGBYbD6/2tB6unXIbhh0jx9yVDzpr06+Ojz4ao
IMSqM8DSh2t/L6pNUVBr1hXBKMwTx61XOt6uO2YX/5vsEoWcEibbODFVOXXsZd7L
KDlyvhOngNrpO47FjEj5cAoWOYg6ffXzAlGRVUKwVICG5Bt23KjE2uvhgUuPCM19
eImpOCV8TZgOnFSwHcmAvR9scPCGUkIzXgfMMAfrkZ9ETNdrxoXPpHfuDpYqNeb0
mnW6xHULzXR44cfgxEvELpZ+wCCaSMqN3OyM7W2mH0UVz/2okwEgutqh+cXJzz87
7gw5GLzLdiTdXQbRwCQy83Ivt68uudG9IwiL4eAWb4HLmcBKelz0aUDpfpj1mjua
2/js9OefvuK7vVd8fLaYcFN10p2z56zVPWf1ouBiNgsaOw3Up5PeDvdn2AotUNs4
K7oeJtWLAxVUQAYXcahwh+903N6BAATQzBPmZp5QAkOaJkNJiymLrH0I9DoURaG9
DqVf5CD2gMDFio+akGU2VuZgpzFcjxxFa59hfKef8ihDl3e8mG7QKQX1xrxujLBg
H5g8l6kjE2KobUfPn+orfEHdSHbDzSfsEqbjlI1S3nwgAlyBUdteqrgR7b51/Fxk
rlFOPtxhJ7aNWxFi3dO0N6S8myB0Kzu7gNRsJCiv+tsFBhTSSdJL19d9rzcM5S22
NILhyeC1lD2wAlBnexCEH+OVspuMI0NcXG3MTuU+LqP/cbj+antYywp3/r3IEaIL
YJpC2sNFJihpT8HAA1jmtoh23g6JRaP3+5ltcro7NUiHUk3vpfM5b8MXF8/S4c+g
uYwXLh4MXQc5SEURP21TtFxcd7hNt9iyAyXC7oCEAsvpNQ1S8hxWDu/ePxtdhw3x
pPwhlq28R8+YjtDJVtm6QBF2ySSa2bGsboyMx2mOvls/3gP0S/FT2j57KG3j2Fsc
P139UzLmpqkRRL8t08uHESoBHaFjFG/x7ao47fWCW0MxQYnGCu0vVSXsZcdIcJ7o
XdfjXKUc9thAMpEkpYOr+Gp0irCQpTEjWkoDH29FqM+u+ZtV6GCY+iyxGHYrcoAp
PlPiKJgDTEAMbc2LjwgaP/QReSy9PjbPK3b9UWbWiBmEWcuTcWMU6fX8l0Y7XOsA
UXXp3rGRhplw/e6rG179kdd48hn2bcyOmuOSqtAERhqiloO5K93Rn2yVE7UFqGB/
1pUcrj1DQQrg5DK4LXX1P7r7VKNMcBwQza4q6ry2RMEDUsGQAOI4Jy5dlGCjJsbF
FKi9gA6HnfYIuyAKgCXc67VIMBWjyFY65KOlIyXtRg7bB2MUg3+VauceXzaI4QSM
FEJ1mUGw8JTr/2ph8m7O9OgdDJjvfIfUamVXAhQBR9BJFdhoJzqQJ7lgXgosayDK
ZwXTMmPVcC7T4I9TRKFvLNdwEogjtgLtTopP7+sz/3FXsYks3bd/k8LgSDAXpiCC
yU4fB9jZqo71S2jmJJytbtpPx5RdlB1ljJgVpLsYcbWTRH0oZJVAUEHVziyj2woF
cgijUC30pp03r61Z19oMZFkHhq2sDAcTf1bYFYj++Cy1ttaAUaugHnAMrafd5Zd5
SPzjI4P7CbKJvDY/vGt0/llw8ceNqXep/ziqvahwPvP2mApYNQRQc76fJn+KqdpQ
np8E3NiAqTM5XHmYccfoURYyqvs8DR60zl/BZe3aJrpZfp2WM6MbNOARzGklR4f9
FH+W6j10i9paCl88+7I7bTzJap+Ii1IEJ4OgcKCFGsLnKTgKuwJMyF5ULlqvTTU2
YcWLaLVWJ2AhRlvhZmyL8E7lMN7kEQt9iV4rEpzZBLovpIGx+2l+zEMjyWDCTEO9
PvRLfZ25GGT40B0+A2Q506n2exca65wYPVbhnuz9yHJEUB45Um4zNb8JAmSxucxP
fG+5tAQag2Ck2qGkK9vCTsrrdyGjCXnZbE+ypCsj7dUZEW1uBn/DGD8Vux9O6UqZ
rZOn/NKVCaxQ3yURuN8tONbWYryiv9gLDeUFNdtv8xi1a46xe90WxVLvAoq92CSI
/YSlQrCUcZWe/XL01FyjO4ESAAP0N5wsR6GiKuG7F51nFU4EQo0+3CMDuhlZFPCx
+8TUsm1TLpYJ0PZduHeS8iIFRDv91kZjtV9I687fKo81242O8zRkSvzSDcFgchpV
LCGI4ndIOALSHxfX6J4h37WPQ3Lb5mOD8AabrxdM2wRw3+Sx9KZch3aqNH4HEDY0
kHGAvhC1ZFk0cowrE6ytGxAeYWY9GTrKTm+g5gxW/nPSS86ExI5zGyYJc2VaHRVz
6q0yr25BT/X9gYeuQJgsEjVRXw4g6SRA3bjxSDwEgeouuwzvCKuY7ST0u9YRXEZY
W7Rrh41mcEP8qO8jKXQgV6NvKNQcSwVpOFovi8pNOVrwsQJl6boiKYeoERo7aY26
qSBn1cpWKzgtIKHyoG1hp9rY7sEc6nUf2aJ0uMRsdPfySOY/US+WUnZhEjOk9/YC
0GWnXmHFIB7ECqu99N+h79Y7vvvXUlAkuY22lpXxJHrElXY736o4JRXPB6+rVcfg
2K4BxHlZonC3j9cerNuTSO4mPyv7DWZKzG3K5wN7CyG0iQ3TaKIuASTBKFE4TgOn
4QF/j+nRz9zUHrSkpCm5mo9naA6WHsZV7PoYNsRywSrejF2FTzAy/TwcRpcS59ZB
wxZnyEUh955y9fHhlV3SPsNawIc9v00zvBf2RuU0ojYeTByJIGUGUSY855Mg/teh
msS9vnim0hmHXYt7m/zm48eY/lD4ibmfMNCxbgPnkCwf6R1HJOuP2Xpvjey3TsS4
1jhZWWcKWYwWfdPF3zOFjUANns3uRmxzjc5uW8aiBQ63SKEN+uTp2tQNUwfmYkN+
SV35CGl5ccM/nV3Q2BfJC2w8KYa9bQ9nDm8aXZwO9wAGzTMYKIpywVjsxxzOc+nm
x+VGz20Xq7F0bslfeT/lXNqt9q4+zLr23wF/qHAALGJ78olsZ8q9sf18NWs57mnZ
OnZJy7h0bsuoMvDEFaYtB490xSni466fZcbzBlv/8QufHazC/V6nD0hyBRbnMDYR
nvkj6+fzNhzvJeSxq58dB3zEEnwzKRuH2QB1HyeqYuSamVKQtpfQM3xLFGN+kKmy
IPQn7Q8GS2jl4OYBf/RjRSl9UU1UhG5H9bTj9B5VCTZpDjeBx9VZYz8JHpv9vD/M
Lq8U32Du4y6dBDTaXUJmLNgAMT0fzd2FznGG2ybsmZpKJB/1kOJuZeU4vF4TNopA
Z9XvQR2V3xoBFvEHKXc81J4rH1Nbmp4yk3MLSkcH9nonq+v1jDws1V17RmISZev+
9qMrSJGOcYUZ4642Kiu5X58Q8y01fRnH0itEzfwAS/5FpN4DT64cpL6Tt+KC5Tqa
nbEJ0FjAmQog6D/4PjgKy39pNr/3E3MQBKzWpzgrkLrOiqmY9/ASVJj5PZwq1XKX
EW8jC9QjsRqboZbpHivz7vz0+8ObF2BiDc0tK4k0S0LKejm0YXKzsQF2rDyrZoI0
xyswAwgmtM+K1O0o3DYopfjV5BniemPP6EBDsBKALFIS2Ae7LwFy78JhO7VUBAPe
tf6JddXyMWixZf9tmKiYHUmJf+pAtR2T9i3FJQoqCVvjkbfFaZmhQ503mC5TsShQ
jNilHksH3z1aGSbIqMp/1jz6/fM8wpXVC5wlX++ekkYp+RXlKyKn10Q7dQjcpzJT
SkjIDQ8ExvdpEFGrzcZ+Smii6kE+Z3NagqAjUM84LleyDW9nXEBpq8fHKj15JhS1
i6io1wSVVaq8wJQpqae5xkcJUzS77BO/cGDtQBoxQJRK7ZUrvlR+zqDqFG5ki64r
7O+Ofz/F18rJcSaU0Fax271ENSOkzY/uzriA6s0ZTlmiTIR3Ssge7tLXcOwzsP0j
uQSGt9eyDFkNTPEWIm4gq0pABDmMvopoqB5yuUkwX9ivHZvo6QjNO4AZVSaFH7dp
23VO5Oso8UkeRPjgVA2fU60Qf8Jd9/CE7X9x4SCsVfnfdKt4L/7EFi8Je2NAc4nA
l9Q3SPeQEuAxv+hxuJRhGmbarnC4sAC23zgHQ0jkhdgashNvEWtuPzjgz2u6BPAL
G3ZPa+3O/KwdUYs8yrMMmGnGUJE0Is8or+J15z/GGaGuXSXx+7sEasC7WSiSfzXi
1LxcpEGHURIE1P/NE85I6H2fPhFWmamoj/VpY+VU7lqVF+PnqoFsmRLJnciJleJE
clOop+anFDeI+X3ywxnQQCpw9YDRQr7Mz09SRnaUCGTBQV4M2mH8AtX70XJ+/Nyt
sHu7mshThHPSlAYuktCt2B3zHuoGzoAW3YW0gJvvpI8cifLfz/1TqwUNzsTbBjy6
CTMZU+3V3+roW9n/xFdyf7LzNcg4AlEtE2ZjQKomJhniBumZiCuDJzxEQwiKS6Uh
S71W0W96vHJZZ0RootxXm3fdeo87EwcpwlUpNCdmcAHC7X/91du0BqqbFm9cI2oV
dJicRzkFGkCpYe7e+c3eQUDEkdSiZ4qsPi0+fyACYNRtoQj3gWld4RjbI+e02PdQ
agWsaexLLj8003ZwnK1n3WZ21uX0jvb44CC1X7m67yxBKGxNnllbJB4B1Dz98AgI
PFRCObkKJdyniLXFUZVjh20wnnZZos22qckt/c56WdhU0CCDmgWfeKq1Vc6XeH1O
RttqkqQ1fe5ZM2ssg05oN40obHpD2Y+EEHTp9DRko5d6k1Hq/JAHSJ8H+bOMgVe5
ou/x2rRGwpW1vKHYcVlcdrE/9laZu7xcxcqxE4QQf0yKjPvKky8pYBNVMV0fb0f1
s4LjQWiCUNm2qDDWXaHJXNEHQnYKE73PShsBcXWjNYMHLtIEAnpkakU+40KCwzhu
VXFDCtTnKbrG1XkFz+CzZbHdzqIgb2jGCFiwJedbNuGbXlsOfvZuezCbiZgP/P+V
IMdPezgXVjUYKxtZiwQVoWD8MO1yh75QjTMZiTejQgZFREjveZzsugLKoM3seiO8
2o1E+LruaCexq5kbFHlZx9TpZZSb/3oSO70bRJKPb6lcyHWPVT1oekhBQUyD6EJc
D3B2cth3zr3pYiL+qHMrMcNEZQUKAsb0XHQBTrXbvIrGJ8wh3B3aErcOZE2tEPi2
FBLy3CK1ojZmZsTdMxpuUL2bHxnOpSMpeCprxjqh6uK//1mZkmZN7rp7WYazirhH
uF04GCIpfpSWhWHXC7h4tk8auMv+LGCr85SMck9vHMeTTWZHYb/9mXCVUr4PDIWa
dlwldUGzPZhfkSbU8b3PuE410IIhJFPSEDSdX6R2ZNtXLzfzMaY08ZiFabiRU/A/
KIe9F1udXuJuIu6a8vPTJdeRggRnqDZGvmC3nX+pGoQdVH16toGLPDO3BqsjfEry
IsXwXrUAgdlfT1oETPPUmrs9oL1QewGyHSyQtmKXJ1oyEB/8yviJrP3IgAsoQvwf
c9sJOyf6Yyos7R2FsO7fplvw/hnGqLL0bTpVhPvtpp8esCm91wdIO+vyNPFr9pHW
VjzR7ByqBJL6xxDG0AAUWfwk63us9bKnCzEKjgpMK445zuuijB0Ngt99dYZSEv95
vGZvEy+xZ7uXPLX88aHl/nYcZ8ZV1ychG5sxqgDuCezBkLPGqt6vuyWIDsyqm/Rl
WQeqLJmIYRISljxJMCoZ3itvN6G9K70uB6hGU2nU2B2Y37fBMCY5tzQxWLheKAzA
KhJXAfX6eqqWpTAzbi4ZWmZhpT3GiKSBq6L6l3kEHeyiY1BlK2hUapcZ7aimz7B1
X2Tk4uNlZXBSuz84eO/62kd6sKWCei5ft6m315eryiW7GAJwTAmUl9ccjCdMHKV4
h7xNDLueqLI0H5GGFLu2hirmJl0HCx0v3o5zUCVHUT32ku89QdzO+DMvbRYnibVw
P0MXPzTkq4WN8u8QjaG6syf++k9lfgYn1mEAIRYRGrh2txpKfvzU8nO+pa4Ra4V3
tTon4plFqa797YP7e+Pv+dlhsQ5VXQ5od2Y+35Xo13UR71vd1gsaIrOMeQoGw/FC
7+iZbfhdtZNjA+9qOWgK3AaeDzM6YFK5rUPnp5akd/KRkcVfs7QEza7sT0C32OoI
3URAswVMUYO/rBsoyPwnODdOU2QgDtsZg7DVtfzPBCu5sRui8uppjtV4epJW52rj
YlGL8ti5lBFOcvp1NZkFdez22lLToXP8n6nXpmLmzmp67dSlUZQFEGjIxM4qwshN
et6YAfBOIFnwH9EjVygQaoAfV8kMAT6CCLAAkzNjBi8S0yYFmYVvHJLrZLEsSulc
L/i7Qi++/XTZ9zCiHU+jWE3tWGkYE9Ba4FR3P/280YWhuYtWM0gZsUe7p1+ZP8Zs
SZbgMKRkqJxOJzKUEsdH+Mc7XO4cJBUQd+VYBQ67CWRV7lgPXQ86aG+dEw0COyUs
wMtl6XL18fbwnM54WTGjAvXOuN3sJwQP2OeeLP/ilCNJJPthDgYdWtBqCrU1OKvl
VVezyCwB82x5GFde4/0SxcmGQJuI63GSWNpJ9+C+eKda4Ugp0qHI0cP98XMHLntY
bN6lfTSaDn8eOLTb0aaX+DjAZ73aXOA9UPTQab2Qdbt/7VqJSDzE8+jjXE8jsMMg
Lg7pua5Hvi2lRBpHYGkcv2nHXdYMPtwyEADzGfk8mkFfqjuUJDkQWLP4OP/My9r0
fFcvCBYIuXBm8FjM+cLeVpUh8iN6+8myIjSHlKJtmr1IwJoSd5keBMi6PoGJWB28
zS1+n/bcFLGMKtbm6epRlIWBtcOj5E94GPZ2L7scgoOj7cSVSx90kOatk4RkOFJZ
pcIyxbkCH50kdffvJVNpHbScd5Ekt5ST1+f4596THtl1eddZ1zuuTm6nywpjRlrC
gUAuFfEqd0qnC9O+J7NgysKEWr1BnPlOOxzmSGiS9ka1hcYB1rirZmgAefCZjRjC
FQqphdKeI4hEGNbn13HEwMTw+Ps9T0m7B43uqddxj4RE+IC1KRY+BLkdsHYs5QOB
wJcSah/ESmNltjEa04XPET8hzia6rKlh/x8+RL7OK/slSa0mVKJAA1VzMB2czcuo
sy0c69L4d28SYQ3NwTQDBI3fiY1wMpUOWfRt4Y5ExcTW5B4TI3w+ni5eIqNcfiwl
TJVP7qnJkpkA27bhnJybDo/rRuqsBDrt5eyyVol8FOJhIcPDFkexKHWfnVr5D4IN
jEhofRFDjBGr/kCJ1BRgFoXQH/J2cer1pRjb1CPDr1gCuCWcUtZfBSzitp0br0UA
09NETvAaLEvh819kYK4LA3iz5TgK2MFTM2fAZ3wjf2Sp8P2JEDZ+aCBUOxn/jOS/
Wtf3VhQkGxQI4ZMpTDclytNtJOyUfbInCM/BBL3cD3f2Qdn7L1V0n1dtgglKB7dL
hXXM3I+98uZnolDPIiRs6Nj78oPefTnrgclIztg02/zwZvuOo4tDvdPlHbyFsANy
kEqySl8m69to244kwfDaxIdEgp2Umc+k61r2jk3i0GbXt5acH8sn5kuM24fAtAo+
JwkUredwwDACdodDbgHLqdw6fqkmA2AuP7KudbwXJxJoZ07BAp0Rmv+sh4Ko2hdC
d6fyYUnW++JkkhfT/4jZGX+Hr2Hqt1SdF/63CBIElrbX+ajJDs9MC1bDaNKITx/w
aKKEHkihppk3r4VFIImIlZQKHfWu7tD0mhPq6E/v8EYUeh/nsbetEkZu0zUAGIsn
vYl+8EKwr1eDwnje68M/9S0GpsqicNqLDGqj85xaPCARaJz3lHJcQh1H0oGxu08w
cf9HD8SE85jnaK9Fusbnyjlf2Mdbb8O7A1fR438R48p6XX7ZylGHwxIvUP4MRl/P
oM6vbZSHRD/UdaUreZ08fkVzaIwT4SCL7ctZq8d0A5no+zOlebCy4nPFlUWgf+Tb
VMvqAteO+qU0IpMnICilJ0hdfuw587RIAaRatn8JkQMwmGYsK9GtXrjNfkLuP1I0
wK+NHkQtYV7I2AO2EhuQOQQ1uub6PTBEruRosfhKhNlM6jJpTLmNeTdso+UMSE8F
RO4RMA4DprYWgliaM95GbGtj/+9aXpy9FXMiRlH4p43U1OzIrcWfk08aiY4YxtjH
QaWAjJvkzlEwWzmIyDn+Tw26H8e7spGQZE1qjonULYLaGjvHWFGFahG+0p5Zh1vt
9GL2K/nvfSPaFXT2erZDfqWwQHvs28pHbJUTy+/jkFxX/de6v/rCWbZKWe+sRFWw
ZNrWQVIaxthPlzE88Dpv07hiR12HUeJjP/XTGkRz+yp9z4N9DcjhuMx+4zY5sb0K
tlDgEzcPRli4cECSiylIShldCx9RLTvJoV93jtuxvSHs/y2s5otfPA/SvaKD5DxR
fGniK60CmhxL07oM1G7rrr0aAMi4JUVRs+SLLloqaHPskPAqL9Vig0vuILKNrN8U
/HS4NsYgbhEPJS33DRYpE2YJ1Mb4OmSSd9LSioPbmFLUNbzTDf8PJeuo+Eiah/db
lL2kSe7U8o+iJm+she2Sn5rrkQ+dcN5RkYhEevCbAS3yTpuuaaXZjtXx4o1KX/FB
K6pr99hOIqn1qnMxRg7pLLhQotGaPOyJjghzpixXSXnptEOmMbopceF76jmQiut5
ntrKJYJtblgBU4ALwozcD2ERtF9VvLZkHfnzNmd+QT75LIdcqEGbYFAYMDWasmM4
jQX8Krf2WIoaD3N9hQHwLkePKfSo4SOiE91JU9ncn8NsxwIhScF6oEqsBFQpLsbl
CUo3fAp/0nzCsDW3smY6vQF7TrJ8CkUaPICOAIAf+nnnBAsP62eB6GQZnaFcZ//l
KDuQD8PSRv7vEx5yfKzSqtCaRxmn191+EF9L7wCRBRpU1iBb2wYnH/vbclXYAS0z
worOujNuGnSpgBZq0Mf/FS2p/FRi3Sr4e2mx+EnDPW0Pa7zFEpvWk4jXSEftE7eC
PrA9mF+0GyQVovINxXfQIXoOI8976TjcOhI6bl96X5Wd8ne0uZUZw5WFmJEti+qD
mC/kIcAHqpIJuRvkPH/WBOMNcdRBnKUwRUrWqaKZeX7Q8Hgvyy/NFn02yVGzA2c6
6LAGEcWT1d6+kCX1KVI4gPo/L3mahZJMDFnPFd9isLpPUbhv6yCsGSI1unMJaXX3
LDfLONKpZcF4jcb+MPfZ7BaBOI5kGiOGAsqe5O+zyt+oi/qlqEItJ8/I0vJuUEot
ppsiZuv591mfkC0MhJENYOFjGuhoV0xpRteRmQJxoJARrfOtG+o/jF6oXKeLhtUm
Y+1EiHzOIpUAWv3SpL/hX1l5+JbW2Be6ScWcjXtCb7U0/+Szbe/PA949abVXVk08
eMxP+0VXd3+Fa5a8V3XGvhONO/XpZ0yTLnqKWXYXKAtsKFmeBWJHXXEeSkR4VgBK
SfSp5J4nY7sGknq6r/RdhdGjrsgQSBtO5SGhP1xV6W3HW9ORwzRUc5VTV1oieBzq
wgdvt8rMGDD2Y+s+F20BANJy7s80C52zH0uMIoiZqWhGww5p5Tzx5IM/Mf5cp6CM
AeVVewzQm3PG7GY97YCU4B4KVD7xtajpovubuJ7a01S6cX+qFkkipTPjJ0BhKrH9
6yC6hYmN7mnX5P1YumsF65AyVaC6b6pTfimDC4AB+aOgA+bgoUbO50Cyc2LAG7NB
8ysCxEv5s5mk9rpGhtAiSY4kkT0/ABJei6l9fk3lKejLlyUoPAa11vP/0gJbzJD3
RvfRo+W/oqlJzBGKV5z7Wxn0MG1pjpI2OFYLg1XJIPFvjLOuFVa977AsWNBmKhiS
2nkQdkBIkv8ULaODZmFEn+wSmYg6ZPQrx/w4A4Ia+KlYiSIcEF0qXuyXAIhfF1tV
fjFgsgmd3LMEPo0qFN+yCKYTzgfjqn1Ex4EHB0tP0aARYMDs8DH6PX9QQXI6j62B
+hHNCc+wERN9O0YSg1aL7WvCXjvKbYe4F1OzPlusgngScpqcjZQZ0J2ZhHazue31
oT5W/h6xLREHerCM/pf0GXNNW+yeIncC5xs5n0vuOW3465S+hl5kPsRrrZaWyz5w
2UVOPBebkVVcD/kMI8oReUiIqyDgitjVp9HSdC7v5QsmwuwusJofB/iaRl3lpoWo
AsvQy5eiHULXDonT5UfRWofTkM08ZfICOsTJZhUjKoyA/OV2GnQdN5eU+ugupW0t
tZv2QCsd8em+xAYMD/VjHv/W2gM3yb8JcYEu8uttXpS9Zo30zdGjuxSrmKJ0VTVE
Q7ztOx7gZAbwGt5bMMogjzygJYRW+x1+fDrBReU8yfJu3t/ilqv+H5Mx9VCULMaX
bHqU4/fEBUNiZ+GAv2HqO5o/eHgw/eGdwwAWArJX34uE36JiJ6coelpR0e9lEnwC
+Z9GENN2vmpJAOAi9vhahaH6ZJc10LXs9wiHapBPWVW+esjmcaY06D+D2PIfELOE
74wl4pMwPKM8IMr/wP/LharPBt5hbvYqmDpAagPG1D1kh/hUqJJ2ECwZ9EbxgSUs
wPwqsNWy7BqDCX+fdxwLX8s2lxmHcBZ8/ms1ZyFBV6bDG8HywtfeblCHNYoPOie8
RRgkkYV6bYmRVqBMPgsAYHffNF7Bqvi81ShSOPNfJVbbmFmfPKylHVxpkSQoY3Yj
/cK2lWMQERfE+oBBT5uQNb6qxgbj14F2QojCvB1ATW8DzIeFQTcibAgdn2udn1cH
istTKm8UN7Z9++X07h+Pj/hJsjmT5qDCvNmAUNwnXMbAFxuSY4kUw3xsuemcvlMB
NSAC3COEhF+0Fo8FnnPhvkR93R7IBRpKfjfXJLG3S1J5HMXQmSeD1CHHegm5sHxB
pRQVJ1xIOonMatoHQhZ1wUE2D4jcnxyrUlBBOMeagdRmP2vZ4ykTDmtbMh8J3sHo
jmSrYJ2za5K2bkSaQU50IHh8Qe0xSdyMH35LUpPOGbIye1T9j+EI6ZRjwxv/yhSl
XVKi4aHOb3pa8KC38U6K5FAKAO+N8mvf8gRxegNjZN76KKw69FK/mlJudTOAi/xL
Dky681p9vE0nTeWzV6R0Dc44l7Vv0zfThJnYX1n7qanJrd7chJw004Ifu79Nwzuz
HzViIlaHcqAjjX1zscfBibR4ooQsur7V/cx6stI49Ml6FaR7SQ4K46fXBgHeEdqE
WJHCSbP7v/EkttigfYSTgQf8nTH5M8jwucfZlChGof1jyW0kB7eCXZZU6fNb61IN
AJq1zvjHwu2xUUqIx2M7WhUethaTCzuXctkAgk5Ev6BJYzc2oi06ueS2ZxIOqf5P
Cgso3Twkcuur2yytL96mHvFzmSCUeAM3+AmlkRAzC6IR+qG3vGn6U94rIaeOgLRh
bL1UBpH7Opi/21kdPjLDiW/VYau8Vu+k0PIWbNWX6K72kJb2mEiUBjJamIZivyWV
3R8s+us9ikD/wnCDNMBdmY205iEXG46QdVc/1Z03JGMzvA69IUwnPDPvBP614FHn
VDekoC+C8KQkvL5wW9qyOHI7R+xxwjceAtBnpTHNlpq42l6Bv9Id7szRqP7oQ7CJ
cfBPE09hvutjnCCHFaWN8sDfVoWE8UrwGjBjCm9dKNY/59NO5xTyppSnpDk5xlWS
cWKeitQ6uueG76OHArjN0YbjBK2GTCkU6g7JUelcm9vwQXtpYWnqjv9yTPw3Q+1t
OgC2n753rMCFH6d+0j/0E6NUSRDpmFTxWmvfKlyEzQYh9pioLGHCuTZH2kFanUjg
STPF0HY9bHfV0lkYL9bUedk6s8w1d/65Pgmrv/IjodxHWp8f358soL2ea+BEdWiU
Mm/7bX8ok9uxqI4k75Ad66vKNZdVth2zLXQ9gBG+Hyfcy+0ftSobLYlFGXhPwhv3
18z3kifbEiXrUceZzTe7W7dWUomhy+6U8t64bDPgMpEta5AL5rxiJ2GypRYvQhAO
GHLqEpsXlY/A7AwsDowf7YXkACv2aD2KHzB8RXU8mvbA+T0XwmbBRGqYlZfi9J2P
qUPLBH305cv2SFkBOMTY+5UA/co+gRnfFdKE54n60hzOtFFHt6lfRljt3zdUgQC7
YydNFIXt/dZXyOPQD8o+90o/BqPYnPx16G1Rb+xl9oYZhfx3Qat2jyoZfRwToNwc
qq0eCdJ1Ice7uSvJPUImj54zkLAEedKxA9zqd/KfuJ6O5SPTgMiUs6mp8P08FP7l
SB/mCRzw7DfNbLvKqz56UCNPomfvBjkaQVKeZ4xfpBM9YCsBYR1pIA6LgMvPsXG9
b3vCImCXFoSP3or8+/Zl1MvwPKWibpYQeXTJj7SfbFaRhTjsN84jWbev4w+Ly96d
bwoKT1lN0uVfBxf/QOSB8fnYX2CcQ1ZVL0nKlvhJp6DRLRAy699tAW9yCicfB+fh
1InSWXpHc7fAtp/O160nKFS6UFojJNEpWZ1owxot8etZ8R+KFXmDhR1qB79HZoju
cm1YKxA3u569EImHS0VCUGc3l0ipSW4us0qrikZcVaz1S6kNLNu4vGf6wl3kvJbV
/BKQmrsmftUPN4U5uRQ4V3JCS4pTiCfiCwp0bUN3bhyQxNFAc0JnLUmS+5vp/UF2
d808HFBuvckkAdb1pOb2Wp9zdy0vQ5bMnOS4F82dst+UtsHwjLKiTeNyb++dXHGl
t7WzWvc+Ua47JLL1x3hgZ4w6gxxh7OWepJpctm3YYjxW5s3tC9DcE2K51liZr/uX
fHSM1jUKwYw+0Z/COGYjAm1FvrLqEv1YTajYvEsXsmA1/6Ji9XwzFuhiWkHahxJd
lgbmRRGZnN4L4Qr0tYYJdfadyZ4TpuF6dyHdJ5g+bH4H5UkGTAYPaHU2HLcdjv2G
wGvHpoLeu9aYc4WTS4E57mwkPi4c2yX/3xPuOuerm6lfaNgs687VRTHy9+/bUBRl
tmQD7vtfE9Py6VfvOYCnDaviFJy7qKJYhnjW2PVOIaaousTqTKJocyCTT4xhAWKk
tiKmjMBCIj2Y0UFTSK4yjyhcBS8kM9sf1lELnDVpqTb85EtAnvylRWn0x/vsP8pn
MXSGQjJkkCqGCTDJWUXbBRFoH5HFmpA4ktdl9wdCEsNrq27kDCMrTl4rVQ1HL0EW
94dSMjibAiOv7sTP1BhZTMgLXSbrF0rr6YJ3PdLi+dulVF/5Ckdxx/VpCqrJiqw/
ipsCewWwZqk41PQutkHo8RJn/zEO4s7qeB5gFj+qb39T/9UE9fwyv2Lr6djtioHH
FPcindsLIzOyJrZQK0/KCC5JNzXPtsfn5/bj/7IRsxrcLFyIxVt7dt7L5l3Da8gN
b80L+dvyzh2b3X9imajR2xn8yKfxkBDl2qXqVjf1oCfQLgIub57FgfP0T6P76ApC
jQgNsYuqRa1tU/C9L5yyxbZkRWcbtwvT7tGFQ7LENSHkGJGp80R/TAcoT1+4xUQi
bNuLF26PIx5CvXs71DITkfCpEfJ025eUBV50Kc0vGF9x+lTod92eJy/yIBdLYWHN
YruiNxeGN9R+wuns9VYh47DfUkeFfVXm8Bq2PUXk3+CAl34or3L9UxCZQIvfMf7F
ChVlc2137CVBFfknCcLUomDpyXlfiGkzyTrLwmVqOLO2Vj7Zw24n4uuLWwSNHprF
U7LostjK+TzfOh+7GtZ3ImEGmqy/nvcmi6aHSdgbMa7EhZbejWaaMfJJY9l42FSG
Gn1orRz/4puAeQau9NRFFeBnnm1LiQtUjtet3fceWCTqiB8luaT4DkVz3vfqkV8G
ET64BKxcGW1fEkcI27Le5xBy2R3BNiKiPRc9gZxJ5Z8aQECC8BPAN2zkZFsPCjnb
hRol16iWCLtiXb8F2CyvPnZ+b03d/rOuvgdJ5uIZvYhcGM0V1N1iHYXp/q2OXK41
YFtzyRb/5NtRtErGmsury/uLoyt1AQI9ez2GDkDp7+K+fa9xdGVfdicL4/7AJPqI
lWOzWSw6nxkzFrytwttdmsF2/bwx2yogLjI5QaoBD5l7vw0aqPLBRjlB61NwVL78
wQM1uUPE9TRFr8xZbKyXnhY4z+CmDwuVIz45rcTfwD9I/I2cs8h57hqMDNZTff6N
GQjHaKLlZA12nV7PCoj/Z8om6NOGckd8nMRpYApEBE4gg+f+Kz9AQXMUqsOL7Bz7
hxYk8VuOnWcZ3JCIqWgeIsRxoiuD8frdgXquvyxeG//DwpA/3uAmddPZ7OyGfuYd
GkYOEWVMAOtUuA48armuiCAcfsU1Z6D2c/zwvnkGvcq5VU0qTCd1oIvfz9ft26EC
VlH3iGKekkLIf+a7wGKI6R+Bl+vR2LYWIQkvVi8i9+iP3Vli5ylczkzVgCaY/Dxk
XlWClUZb7q726pOZBlefI6LsX2fv5yQA2ThVMcBuVjffLm/suOtunGGzcgX+Ja1L
hFU480w2/wH78etLs9IPD0iH0LP0JxKA6zWPJfQspUcuGlBw71YmMbAZbXHVVxuP
ZqQatWmTS4jaopGUSlX+XIIhloK1PCI6yQDM0tfmyuh2TtU1hnVb+42WI9uIX16r
JBPnDafjJNPpUlv6Pvp0zce+PV6lBKg0dc9TxpCadr4Yxz5KWV1ofkIfjo5x6Wf5
pGvM/y23RAl1+dwUCGPmT6pDPcn5gpaeufzaZJMkMS0vGOpUhA+p8QN/HGdVaevn
++0pRqSAXXxpprG0LNDA4A7TMJ8HvL0UFHjQtuUX1QymFDNsNjP4LXtrrSLwKdLE
1iOLywhQhA00Dnvb0FLBg/HSXHzBfXVTHsErGF5SbLuqFz9IC4NIq9kpeAfp1toA
nf3P40KiYnc8Dz4GwjNWlgjL9k9aw2KdUlDgGfQqV30GFkl4EDo13ryzNWAIatQq
Ov7gmd2fBVOMtk9tte6YMC7+F0gQEnZTXYdLl7WTG7u9Olws/W5YdUMLSbDerUwX
MO44I1pQzz7KfE+qo7hLIwrorS5wAJFSTLD2bJwB7M8+t2zmdJI/VrCPAQJDehFP
Jti5zpsfwbu1B+pd0nrnRUsFRW1dhL2RbBViEds3qOCaRcfsk8mtBi6Ls9ZXFV1x
N3jBlfjTsEoJIF2TJ3FFhxG2i73hjN2VzcKt0CqvVp6QtzKI13iSL1uA1uB4tIUg
Fr0P5GQ6RzQ+oOLXrVMzG+zkw/VyPiJSBzPuonP5XCXktnPaTQXM5FUOItAeqYvA
fHEBre5AqddLdHvp5iGKh/SiGCE3z5HTs6NUApsGZZD5uKHqH7wnVP7VyX7ARGbk
eCvP7/eswUdNFzsELpcCpOb9RXX//2UGcv6NCwpJGdEJU2QBQWJJwGKmxCEM4nub
LkCbVpPDlXPMwnP+ph04sPBJSgR5wdnbb35P26MfCku9fKVV9Ai7WXEdBSEX6/1b
pqFCkxFxazYifkIMmssxA6Nc4BI8ChSYQVy/BGJW/gNHHhCu2Oyfi7rPMxJiTkUG
qZQYyn30oV3uJrF/SAqT8iYvWBg3W/1yV8zOjNWLcBhXOh8P6BSgGWaJp7traj75
7sLqC1L7yjIpEg6c7CMaTFL+fDe73MCJaoh/QUeINzcCxpkZRtxEZqeNLN5/G1mA
Tu7Q2UA/q9Lhnl2NdfrXxbjL6lEKjtbxOe4ilJBhEBXPZ/aeiQNZEXOnPLXo47VM
FO0nz4GsLlRJrWvUOowsA8uFSH7eev/Z2YAUstzdMe3kvhBuq0nseLRcVANOxrzo
tdCzF3shrum90l864/L1OMWVze0+qejaTEpMgcT6ZWHmQ8C6/QJDvUeGZcktiQVz
vgN0Qyy77Te/J3NvEVry0d0JhiaOA3LFZoq8ph5vjVZ8W4p9m6QYe4Ek+5M87LHW
jHG4dt7hPa637mz44xIlUy85o6HQTvQK+sK7keXaMfbQZg1lf6nx/L1fxJOamXUX
b2TPKI8HTLTPOQ3HZ5XgsjcSLdKUrwauKoXKl4acN5y35lqyNHJZ1z4YAkiSkXZl
llDhazWZODc3fKzgK22+C2Mb4T1QWhhcIhGMli9K/aCvuDic+DmDVUN3uRHmxjMS
mxqeOOFoKY2pudf0Rtf6DZJgaZZTFHhQ3RgP45mNTrpc4MBYmYcgEBQ409O1FW3x
T2G5JueZMSKYerl8I+I4Xy/zjAeEF9hOSf939wMLBTwICGXSgQvI4EONr2HeMpQx
kkGxaydqN3gqKjTZNmek9vkoMEw/0IvJ9i2OkvhbY/LPVk47uicDEPga3SQFO7/2
+KLzmHdVS7FCz5u6xUAnMEK/Vqb9PF0UBMlj8wM7PDl4025TApUtcv60KUwrqunP
/4ykCCadMOZNXv7jdrw/GcCbJHJTJyMzEbe9fTFIsrY0+j++8/k8/KcVe1HMMkCK
lB5IY+RpgJe00nJn8qzAtpeW/vRMx3HdCG1MXfnPdF6c2ZEhZExls6LPAECHrQWI
VwddA1FOlq/EfirpDk5kZ8y+RgQ5oz6WlMkrc6vt7ltfl/oVKaCfhU70Wnn0Dkr2
1pHPYSN0SWuLcP+7mG2ppCsv2/KYS6LhE+oL9jfso8lqifaZxdnOWfPp3WSucEYK
VCNndwrPzZktnVvyX7x8+Z6rSyDRYeK1jNL5dbIiaeKRNMKlxsU9vbEiZpV6QxQ1
5Esx6pVX8h3YLdeFWVk4d/2mUmDCKYqoo3OC+SH/dInkH9B9YWPRnIw2rbYYZaQP
56tWvuNSE7ukuDtYNKeaxAtdlp3GwVYnAUq1N4XWv4DmdnBfQA0WN8D/MI91M7Y/
OhtqVYtU3+jNT+/5DRcbNkaiJDT2dk0xW1YeTDV2aB/oke2ysVUcV1WJhKrb+FMA
2wayiD9LcnzwGpLtkofixvDxh4dDte1PM2C3O3JoahRZyTCZptXvdYTDEaE6tSgr
/dVy5hXusiqGOYOjPg/rOnvduAscBW55RzcvhJZymQ94twI0c/8yoouADtZuvNnu
NagslKsyZMgeSl+55svnXTUiOJseHtmB+l0ENOLOfOtW12xDqpv5k0ErR3S4HkSf
hOFPm0AKjEtmqGX5/IB3XcO+bNuxgyx0DThVzEdoHFFpusHIFHaVw1AhhZIiGV1F
k43ZvKhTOt+oaZi0M0ULwtKHCh6yw0EyEz+gheIfGjnrrJn231ZeUF81VylReYvs
KFPPvE+ZWolhMSHsJcYG/NUP8qtSkhs45wBwosHaNWX6Adl8oDg71d4S4bp6N8Wn
V1O1Tv5fHrcRg97Tb+p0OMbnclL2odxyZRAW0hv3FGSITNkHlV5eh7iIQ8D5G4SF
dFGSJuge9YSaRPV+uFB69BmQ2mFssDTDXuY97JeCDMB33I+dKwu/UsTm+ZxFxC6a
K950xcGlVoZYQWBzoYU7yus1rqyhBbSAudWPHN2O2hdnxdFQGzDyDDVVdSSVGB67
3WJYUqChYJNHKJ1m835wz3xFxIGN9JhmdcMZNQFMOaDX6Mduym+eU5OeF8LXe77K
8yj7mXKZ3j/iCpp23u2cIb1l0Yxla+ehnldhrForLfD+II7Xgjkh7RDrte4sLiLM
XoNs6OfBYW0xk+IUORpm9X5rZW3FzMJdoOqwv0Jsmhq8wP2adbEBot37OnIxlG/k
WYcaE5KGqUafQtCCsxPnT6cMg6c3SdX4z3O9DZ3ufDAsI3i3GJsEZUyffob8TGd2
sFIrort0s3o5RRDZpbjVomuO7d6bvfMfW8LN8H2toQqMxr3rodfL14tKBBAqQ3pe
thBHoQlnH5NmM3OTJZR58+szPfHrJ/d+hUHLj4snNCcJ4oO69Sp2HbmtKYkj26V4
ylW5x7/17X9D9NFqH1zfffd26qT96U0wtjFfKsmPPSPKOI3u9CAeF/lr0gZsrE1F
yoeIlCw3kItNBeG9ukmEbabutRi4c9Um1yMrCXiADUWZC8J51R1+8vWTHRengUFp
w7GztucXlSPFSSpIxEQNKi/xelr6frpz7qSQZedQkANuw60m9cpnu3dNlnC2zTrR
OmsHhHEccqd1RKwRJzqzJe32O7d3eP53tK5rexe4g88bUZnnAX9GlgNEtgUcjTYQ
BxEFTlIfDHD+ql5/6YRft8ixqGq41OM4XWYbSOgDzEHMIf36Jky9uyB4CKLeiVcj
GXUKEIYPSsPkIVaknRDKJDwBltdxpbuPYvScAUW5iwwjNwJChvswM4kq5VORbVZL
+fV+rw1QH7xQXphKyGygANzg9HYMXlTE9vVGj28DTo4fpg8M4eev0kUi9qX1+maH
Zv8TqgSCWOgyDkcsdmnVySvh47N3WngRaK2iHMhc5IcZC9fdUoQssMZYF0zkbnyB
s3yODdZm0/n5cY7BlwXN1FLx13R0hQaxXs+jOZKkG9/yXW8eS8AXUJ/lBodSTXxo
zETrhMoS5EUDCSEkpCPLSivshAZ7L+n/+6AABjiLvssVTgbL6XCNXXfXM5VMgJgI
JzqQBE5F9C4wJMwGtPLVpnW5hyQ5sq2+q62857jsMHfKrbarTKbNt8Lj14QfZX/w
wjVFIXBukgLWugsLS7JfVKeuRvDzoZn+kVE1F8bNuYn6sZE30JQTORCbcB/T1quv
9o/EyTWIl4RUiLX1KY/3nw59EFAuzemDNrw3qxWcnidbaBqVxiTVKKBKhoobmFLO
fR10vMOYOgN2YS0XtkzHpW5IhOeD0rTTAmM67TnaAUASrr9sdLIpscJzgmc70tvw
MEOXvqI+WiNmuhd4wmgpEMT0ckQaYDX97Gg/IkI07iOrUe/h9vw7lYuh57S3gW3R
1e4wvSIfkYDPDhUAluxLYfpbPOuwk9LAfmlRZ5HHXkhYxQnBPg1spik/Yqumerwx
EkAnTLtJkfUw3eDDdvRtqVYDCKUU/zxGEomhweQt4ME6JTEbqDJh6duusdSaJWOv
OFTaH8L91y0MxEHAxbUlw02TkuATvlSAVa0SBsvgWCegVwD/I2B8Te0IV6LSjwAx
2uEBIpjr/wBNTXKVYyG2UXdZKx+9aKNabVoaaVEV4DionFiXl02Xb1iaxUsYBu0d
Erzk1SeUzLQeP/s9UhTkwQZRYSXhXn0JSQe0lYsQgxIIMNtmbLDdr/B6fKUaPLvB
zR40hU2tD852EWuLeOtO/NKRv4x3p9EDPlwgV+EiRChtu0ew5Vxww/EuKSQF4+3k
luI8G9u/b//xK4ZziHRtjUl/gXOhDKOz6MwSOtJdvuD9T4awr591A13IGr5lZPom
gb6bX+krkJVQBipD8vAbPVxIg/82umAJVR24XK4MzOcOT5no3t5nVXjwmXsxy2QB
KrJfGZiZO5ptQp2CwHh2I0fgPBWLZBqAZ7W6Xr5VXOsodD8u5h0po4o4gd53d2EB
OZMpTRGhBxmT3ZrDTOWsoh2PZ9WvTaF3/hT0ie0TPy7+qjm7/fp3M95++HcO69PZ
RNZgeccxk7vRBr0q6B9kr1MWHQvTswJJezwkV593KgQ3E8WzB8S7qqOvTc4sVDER
rJlx5awQYl2sbKhWk5R04AgqOfGOGE5+h3dWwdGc6O9GWK/bGDoD9xnRSRK2SW/k
epL4TVS5jafDvGIH/mFdBF8FvNRl6NMQSjQdAYzX/3b/wLIpKDOUY5nAAoh2nqVp
aTRnPvHnr/j7cqCDXofOfGW5aQqld25DZ2YqUezRIelVsVe8EG6S0hGQp7eSICkJ
LiAw8MLSPBqRU0qsOf5D2DhjehN2msmEZwzACi/AN64NpBNDQ8uMrHUx1PEyJaI2
h0PiTn1K5nqhxzmxsR5jpIE21BR+Y1V5ULB6y+tV3vZqRlI/L9JoK/qiQw6vquFg
GnfU/qo2d8UJh95W4LIkotYhJk8OHSUtl80VfTnD6KAFn/qMUHNHBRczpBbf/CZL
mhH1q3f76bwnEYIQjm2ITvhDylQ2YIqnAY9bx8k8ScYtqqBnVdO8vDGpksZPESKS
uWY7iVevncGpnnt/NUAVoBMheIaQhME1Y9HpRiHs6OVn5FWMhNPOytb/iGliJS7P
cINRZcYT9dBEDPV9WRoANFya8DM4kAW6TgCEVCIsP1ol+sG18Q8rYUT1Agm+7XWW
oI7QKJCNPrtjKNuyPielX9uV5nVIbcyzdmwLX1rv3HRgkIYTYOLRBF4UMNKHzz/i
A5g02rvtavtI2fG9pCd3R97UWOZzLz+9S52q4KeQ1QIb2938lSoLhDvWq8fK6ni4
6c41fVi7h/aZXtsJSv/8QBWpYzpoAukrIdZ4voy3Wpk=
`pragma protect end_protected
