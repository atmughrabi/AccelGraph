// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HV=2TWLH[J%&T,*@=?C="O[+31,OH4:Q)((_"%G$1>O!@+S6F4J-#G@  
HJ\_ =+\35@(>7K]:BVK@.5?['=&97)U[SDK8NJ-)<KGB@52!?='AA   
HA'X,GCJ)\_-#8\Q57K.V6']/H%OGU]3"$][PRP2JV9\/I_^G4B.E%   
H7Y(P0_**H)=U0*Z)4[<-6EM.+C;Y5[M<Z,,&Z!K]7A #D@O,QJ3IY@  
H;HB3>.@-EE<=+%43-<H.K:GKRJ8$"Q%W24\=6J2&FX !$HMD6]-7]P  
`pragma protect encoding=(enctype="uuencode",bytes=9680        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@B_C:^X-'V( TE@V3#)0O.:Q%I!=8J0OPO(^>1J^#0#$ 
@D6(;"B&(8%TW**\$\:3 /O=\F6/;9C8*\C'Q-U\#C-\ 
@<SYT$IYGH3)YBA@-F/@@]DF(.DM6%&.<X397&QSS3C\ 
@_35/T'[*M(6,*F@^<PL=B'<N@\..1$+JB&;.:],WG3L 
@\%%:[A))8Z)YCCPQ784$E UI??:%/"Y6,IGTSS@78#L 
@O4;C!*2]/GC'>V0E="4^N!/0\QQRR'Q8$>5:"*L,M)@ 
@S>']-1FV??[RA'30JF;JA7= P4[J]IDK:-."2)-X7W\ 
@_A_VQC)\)Z_J*5V4^D(XPTH7R;Z+6'!HFBZK,21*<CT 
@7'>4-OS1?A9__U27:Y. 5W*H&;++ N\?U!&G2=>.GA@ 
@BF6 9?/KE^-8@:MYA0IE"@W;LL8>FHJ)QKR^O:O5DCH 
@NXW29W66D\'"T0-*CV;RZNB.LYQC,"I0JC6G!5\)?KD 
@_<(94@P"EU9*\]8,.##D2E6]]YNQ0%+Z]ET)OM].97@ 
@G/*L'=0^8[2'?0=E0ZO1MW=9+O4R=6!V.W.(!2 /F$@ 
@RF_Y7O7@;<4<U->^FD5F[B9]#91@ZJ' JE!&""G\VH$ 
@J(;CZ=[$CINC1^3, #&@HI]>.Q6M=S."@)KWSP"@/M\ 
@$R=*HP9/!)&+OE:VW\BIC%Q724_!9!??1CN"=+SMW:4 
@T"+SJ]BEVC/H@WS)@HT^O SBI;D(&8*5V^(/UR404O\ 
@53'M[6VRQ_K+(_E#1Z[_4KG48+ZX#'['LST-2IV&RC  
@;G?.=MB[[M2YP(^SY<>K__FDE1D5<O>RS4U\!]8?9<L 
@C?5S6\?<I3G,IO*-79N_X>W\[WT"#$-8&(DN;L3XJ@0 
@,Q)Q_P0R1VL=&&X =(W-3R-"6/O.'6W3%YB'A]BYYM0 
@63^5FW].48('D5]O%!SB,YW-8\'2Z.-X?;X<!>X^KWP 
@3(JEY<UV^:VZ,0M40<I29<G+57F91D+!R4K,TR>%6'L 
@5C/ Y-.A_PN MR*;@#>8$\G0U+E!(Q*/@$S)@ /[+)L 
@*T0+G:(9SVA""VG>&UVP?!$/,E0)&GH2>%7$&^-C=[0 
@;&UFI:S3&F:=9=YYJ&?DF,=+-NB5I,1FR_Z7:,MDG$0 
@!I1'H?Q58AU&[%QYI.$;PL1>9WWQ.%O\C8>V(,E,N#H 
@.'Z1X[QUMH_BL$W$4@VBC;W@SII@8 RY:SO'@S!8*%D 
@U.NZS--!$;C_!$P,OW8(YWLT! #-1 C%,-\*,OJS1[  
@L9*CKR%8D-AG*ZQ]#AC)([Y;<#K%%!(GE4BSVPO\ [P 
@:WDI':SZ7,UW=A POJ10F"@^9Y@-V0D*651[A2[8'/< 
@LH#7OCQ CZN%^]LO><^PVXN! R%&B=&YDI3HP6I%SRH 
@_I#?!0;XJ9(^*L1QQIX0RL>M27F:P5!PC:X+%3-*3I$ 
@R)J$_0@_E>@%R^'46.3VH +'H7/I8!/C4T2,] "U%'X 
@A:LB@R^.@4Q%64.YL@0BEG>?=].V\:5&)WL0*1W7YC@ 
@EOT'2$:N1L< B"@SZ/R++ZG6+DE#+^TM]3:)B(L3644 
@EU:G_\V%)B;&3[#]SG.[19?<#DA\;:0L7=4M2WW\NB@ 
@Z)[).V]$*KC"!&T?;_^LAKJ[:C"6>\ELE'WBM>0J_(4 
@<Q^Q*#"?W"A]L\^,1CNHK'2*IL[='\G%WC,7K[KY,SP 
@3:<.EP=C&N(0(QO9C2QAG4[E^XK<0Z)-L &;MZ8"!9T 
@0WJWC-Y0S]TIK,/.';N ]YD+R0/F<]H#3Q3Z#QY^VK< 
@29F%,DS4< T7JXAO&V3VH/EP]H@BQD_^3+Z6<XTC'1< 
@.D@3'MT=]\#DY F?H=9PY.2%8,]IV_IN>SM3:8#.7$X 
@R,=;3OF,)4XQ;9RLR[P%1JW;3##W AOO+ON\S#5^!78 
@-(SU+I>'+<:*:>ZOJ)RHA"$&K5,TOM64A:YRV^S1 "P 
@=Y/NO80)AKBNHS34<T7'.*OH,VT-V!J#RD] X.K500, 
@@UDP?&E%IZ=1>L;.BMF)EVW#+.UU;'KJFZ^1Z-.*RO, 
@\E78U$6W"OG.=$&BX9\IB6=;[[@NNP]9?.3VAIZML;( 
@Y9RF< S%2L5=!AMLOHM1;U]@205/_!_VXH5Q7$K-*@D 
@;2QJ./N%ODD>!)J5M6\6*#%^^ZI93T2*Z<8KLE-HOIL 
@E@TE$%\Q&0XFJ ^VN!NI)J_VV$9DCC )I@AMRJ[@OCX 
@=D#P8Y#^B6_.S/P9!@9_77^)A603'_6@*0EM]$$_;0< 
@,]BOM=?U2&5"9!,\?(:$$86,&-3/YU['>02&H2L#NG0 
@X/N+INUH@MRX%(BE'3]-R6)+%EZI%HO4IO\GO<#JV:\ 
@)>@HSW-E=SQ[!P!@(8_V!09]B_FKZXM'= +2.T);<'\ 
@[G 4&#HSDB*@>?WY0A &97ON>Z.BW<$6M,F<+G>J7Z4 
@"(ILY!\0[ZM]<,=2:H>-C3+$L[-G\OOMSIMNAF*2&68 
@/C+%*IRA'SNDXG(\T5+<8)H4)TAM).EYPW#\;%?,B/\ 
@NZ"S$(U1V*<=UDY?;-K!*0+G-\T[I^517YXRO1K0(>  
@$^E]88H&GAW"&]=_<-UUSE"V&KI%!S#_M#*Y9H$J39X 
@KJXSW Q6F4>@,2>@!+1(<\8SZ#'4@6J@M'^W'/U1\3( 
@-MZKE+$4DDHQ/VBM?<X*M"E<E.!Q99)JN_13J*;LS:\ 
@5KR-U0P)O3Y:LTDQNR]YON5"1K* A[=B]7CC<RTOE.L 
@>?+LO1&.6![&*^BIR<:,,$QM]UN8-@%5BI+1$T5GPR8 
@#M[@:(FR)#O=(>;8]GA\$%E'>PO[?XC =8/M=4ZO7H  
@?U!;UQ=W_( 'F+4:L<0%IY*?/YE#YL3??!RJ!#J!1SH 
@%IN^K=F+[!J11&%+=83]FY;','/*[QIX 0+"<6X/6+L 
@+"5'7=(W!ECBB,B_E+RO(YLI]'Y>"NRU3&*#F1[/0($ 
@A(>.QGY\HS07(DSD@+-F#-3#[#8&5<61<E"E#])(X_T 
@OK!<GY?M^-/)(H-;&<+36YD[ND//Y)XN^CLV4#IGASH 
@!%RL>Z"GH*\.B[8S!?ET4-\A#)8Q!%_\/)-:5;DS/IL 
@'CN#PY'.<)^IV>$=#F]6X4!WT>XF53T+G:':&=Q4BB  
@$\N$B#@BIQ:8[?WHR6!SCV3)]4[&S]B80^9^]LI17.X 
@B33X8C(CHQA)]1G*[+Y*G$('RG)PD<E< U5'>]@&RM  
@'@U134>N+PE&04(P<F8DU.@,H'N#0=H@$M])<PZ_=38 
@LEC 8O;2]SW3B?EL#S^NHNFU8GZ'Y5N4:/KLISZ6W+8 
@&/A*(9.!&WKW C$1X V'YUC(NO1 OZ:S"%50Z<$1 QD 
@@8I$OTU\ 7$>VKECYS8<2*02&JIDDWO<&C4KX4H+:(0 
@&I&HP"\C\%E6S0Y] V?.8@5.?+KG^8=2;\X+N:54IH@ 
@XKS?S<+E(U]WZ[*9X:"YO? ^B&5X'0E4H9RZD7G'8Y< 
@ -FSA"X(X"F?V?GL[T^;D4V&*U-@C=2H3*W)5;;FO-X 
@YA[]QN<J7Y!?[V:@EC$JD@_H=>BW7*HDGI.8L'$#O0X 
@LUK9.R71F@AMYJFPW*1RCX$\4B\'/+E1?$8L)OQ1'CL 
@W,M[T7;'S 2-%A!HUD1?A1%PY)8KWDB-^W_@"WT HCP 
@Y"1V,CO7R%L2R/8ZY4ZDL1PGB%S8B.A//75KU$?B0!D 
@L<AN"<%F,5BM*O$/(B+J#78"\WM7AC:>A^C]I:I3L%8 
@A6RT.OCL!.-^)5R&%V+8J!M-B^WF9_//H]H_<GAQ&W< 
@H1;O=QED B,L.0%112HKR/UB26.V&6/O^?G/@6O)%C$ 
@I3XQ&[(U+/%UP- CC:89*(H@#HAK4OW U_L%MD;+K/P 
@[X'^.(;[/$QC<!=&FV=V.;4 D5RI*+SI V7[U?,G:[8 
@4 3N/I/O$2R+P2-0!5'2W'QCRUS);S<)?V:N#]S('2D 
@IN2:TWJVGIC3"QZB3[==XW=QE=?M?%U;%3$]9),]BJP 
@3TZ/^]/?M]@1 F0D2&J'.B0X/'H7"\C_D,U1>OB"M\< 
@EIXN9;>2Z4W./\B(+^/$0Q_*= "U6+!W3!T1OVW176H 
@!EK^M\X4UO5K>KS$\HM[;)A-;8FH"Z1A-MT^C-Y5'Z0 
@\P\[(JCL,)]R_*3O2MWW_7EYUKNI(XBJUBOT@<>(1U< 
@?ZA7'K8YCPD3Y+E301",%CG[X.86S_@4X0\3X?C;PKX 
@'YB7$H\D\"R_TOT,Z]I6>!!OL=<G,2WL8>"!2;U%;TL 
@!?,C9@G=,B&;R79L9-#G2H9T!3E2+Q%N/S.N7(?')1$ 
@,A9G&[9@U41+"(JDQH**)^/\Z)MH]$0LIM:2&!0]8-0 
@4<B+PG125P$GW89#)X&@)+J>>D-2XP6"7%SW_U !A0P 
@^.&#Z=+]5X;\3+EM7@U$V(/AOESRB"I9)BF?R($;9$4 
@0*UP_EPD>,YZG]FMS>T92_R%+L<N "+B(*!*4*.O:M  
@L<M(]NDRR'*(3HYNU#5](+"O1_:8NP^K)N"&?.BIW[@ 
@B,.C-U';K.CD<C.F$9?<A4A",X?D1A<2[.^7=I3DP-8 
@,G#-W)<H.91B[;.'HB")274.--4[B8LK0C%>?'UXO @ 
@,>9FV=Q*=:6^Q2Z*Y8F!!#P#.[^A0,!ZZS;(J#82S8H 
@KFK,\0 183Y?$%P0([#KXIN]KV[^RQ*7H$X[N$IT]G, 
@XM))@Y$KY,(6>'_QS?>TQ)Z+4IZ46R[*>>N,&@^,(B( 
@-SG>#;4NSZU=!]JMR>)_28IM%]@]? ASVOHXFQ_\J , 
@AD]05V\EJ6B.03Y&B<H;)XEI(*HCL1=6_*Z%H"DI,CH 
@BHBZZT,ACZ8X0GNMU[@,++L>HB/7J4U5GP3(I^AP1L( 
@S>S93C3/ZE*J<8X"$BC --U/[L12WOY95#FHFH@?]*4 
@")_9M;_DZ"M?'T[RR7ER'O28\S<'6SU'8/IRTNZS GT 
@'6>5J)'+0U\I4KA$#'@\LP#!+97)XJ)L+@9$=C]*#\X 
@J>W4>'E^DP9ADF%+PWNH$!09K;N8OSSL>BJ.-"6=4F\ 
@S?:&!DV_?SC^(Q4%/:+[$O;AQ1RX'*$;U.::"W+A;A  
@G.UT!_W4"4*R?]/]C>-K*\//\M15L!N7T[BC4FHNU7L 
@<J:+$K1#M*4 O3875\2MFK< /W^D3BM#$EE4^LRKYBL 
@'9KX=(PLFC#6MC9=*U.%W,!<\1.%W'^_&.J2Z6\GRTT 
@<-IF,<@0]SK@+N,P@]!!2"_B2U"4UD/: 3[^J/HVW3H 
@WW0N^/F&-&TJTDBM?ED7U=$:M_:Y/V N+CG7+K=?5G  
@HRE$O\'$[%/H?MQ3#@A08ZYZ1;EOH]Q[$L/3&,=33K< 
@#J(H0NP1UE1U>W:JNX5Y84 Z3T=19-;FQC64+1K[^F, 
@BYH7S=)1 T7%R5PN24F_(?BLK<HJ>:'[9C,3FO9-L2\ 
@RQ?. )<)TFGWM!ZC9 -VUX</EHN,)1,T>-O]C8B)\!4 
@*A:5%,F4#=^/Z*X !XQYQ[:TF5Q,]!S?XI/KVP,_[U0 
@G7Q7K7-=<='+8Q)?Z"K#(1=@DT6EIBDG6UY#$5%_)&8 
@JB.X?@>R8>1$:3G<ZU5V7CU:-Q)?N=#1Y/KFZHOU1$H 
@*[(*1109<VE%^Y3Y[)WF=%7NT:K47JX!><DK%,YAZ10 
@Z* ^',:$YQ/H!K&[:,A+2C8 .519L#/VYRC0BM)D&?4 
@I*M;."6P<T<*):JLH*;=+'80AV]XY<T,3#AS,;_RAM< 
@+LW+FI>@0FL^3PM*<%C;9)10F NRMVP5VSN5GDP)M]  
@=P21HJZ-PP1/_V$P&;G+'S4?, XW& ?Q0)<:I1*RT0( 
@KL[J-@TF)O[4<:3(J++&3C/7T@U1L1RL^D]7^%,['0\ 
@_X,O&<M^U ^[4QH82$3=T^9:1339FGN$2Y3 '<-;;M0 
@E*CW9<@%&(9 ['4-G@B:@!B2/Q47246 AM%@X,*<!G, 
@ 2G:^V"*Q:D]+I]RUJ.TG*Z%#,-J)"9+&C5  )3RE,H 
@9WI:[\JP?]W%2'3WB<-W2\VZ9W5D8RX $/=)*"?]U94 
@:\0PG^<#\N-Q%#P?[TQ@X+>DJ=;0^9>XO-Y"Y&+TW18 
@GXE)[DWZV CUUV8E".J&R))/'6KLZD7/CSM/@IXO)8T 
@7 ]GG:5P&A-%AS'R8NG: T\DNP,'7\[C1TQ+'P*PRS( 
@$D).M YY[YJV:GY2(,3$"N_&JEDS+2+P<H"X"'^8&J( 
@RSU=T,X:LPUXI]K.M&#6N]$*;J1,SF8=I.=[EW6\MO@ 
@9+CO.RS[IE<.^H).%?5EM3^"6.R@ ";TPCF"<^B'W1< 
@.[)[]>0@%(7;^TYAP\:W)YRMPN+[[=B*:^9S5^EO4RX 
@_%FK]2>'0W)NS&8>_#(&CJ-1OH1#T810NML-*_Y$<Y@ 
@EL0/Z[H0D%$"D"A RM(EOE)CO+]")< UQY19E+TLF&4 
@?6:*+4XR%9[_/$/GHWF3D9V91A'21P00>\VB:;RGX:4 
@PC_5A1:<T6F;U(<!E!]=Q-V6'Q:1Z.DJ)DN@CNMB3"T 
@D=-#&Z:9J(FVXM-75N3S";V7919 Z3=N'WSU3<I+K7X 
@G$J+70UO).O:4O'*33R;2(8]\@V9!TGZ[4(=_EYV-%H 
@QIP*Y]'![?8>JE]2.LH&4Y96^7X]60(KK$<M8ROH]YH 
@>&N@2AJ/2 B<N507RI/G]BQK'\I;ZZGQATX'R-.S1J, 
@XXP)J61SC@V-[1E.ZS[TNX.XC8V[KR<P.2'$90IG9\X 
@",YHEK7(P=OI 5ID<_NY!'TY_AO44]@8$&!(/>(?F=8 
@M 6>+'1#@D].3Z$PV:<MQ+.%29CR5FR%+;SL=F8_V&, 
@6GNL1R_J=(3=I7[FT>*EU('A".K)>/L!!E"*,GRF0"< 
@6_/KCHT)L(MNCCG\CK*RL;KPN2WVYL?9&6$#S[R/?I( 
@L_K]L(<RF0P2>NXF'C5\79Y0 @A/E1\^I;#8QE>>=@D 
@L6\%LBU*W=F73G6%6(B%@B$F5US..+^MDV3@1P8P7%< 
@S4207$CZ &/63Q?)IRPQ\AYGR.Z9>&$ !,SB:R/SK%4 
@;J#'5*:XGA=:ECRE3K^<,M@C\)$IM6EE27/<UQX2:J\ 
@2,QO-B8A+]HBP*-U&Q8A^)5DBF:8&68HT(&B[8V_I$H 
@;%4C_AMGGS9;4!0@7+#^U"I,J*$A>)JV"R;2]/2]1Y8 
@).'@ERU*VV 0) B;7.20!R.FZ"3 6VM_&N/J/2-@WQL 
@#9?=EJ>L=M1Y?VCS(*V2R01IGB>I7RHZSJ;?CODM@N< 
@QQU4%_-/= PQ @Z!$L>M*==PFH%-X5S$76WVO@$Z!'H 
@<0=0HW9?OFV!><][9UT+]KLSHV!5WQ$59)Q4)R6VNJ8 
@B$MM8PX+G3DGEI>N[9*0B$LL7+V]C3>N4)6YH&F-%@( 
@- 8&:F:4]D(UJ9EL&1OUG@NP%6*KD]TV"?%-_;'%#K$ 
@S!YKE0"AU,5G';?NKN$AK;4;H[2U.YRL);S<FKEN:DD 
@K5,4@U4.@NIII9+=D65<&^C2<3L5_'M!;2&I;.<*)7, 
@W.#]%[J#FM4TGT&]#9]>SG\V24YT]SNBB@@G$IDY(;0 
@/I/$N]8K;(S/T>&F7V2!'IHHGB'OP:@@OZ6']P6I 84 
@+QF&'36N"LP,+M=-EYC(,C4#PF<99:K=_CAIY8+_( X 
@)K?H2V+<:L%@SCM:8<5.VP;<%*H=XF@WKDQDSK]<[/H 
@5]&_<=[C=  8%A+(N,5SUEOD#A"N=D2_R]'?$'6<!KX 
@L[Z<$1F;>HC*@.1<LWW6S*Z/KX%3 AU:(WK@#0/I.6( 
@J$4V$OJ%?'3"O),E!7-R5@9DBTT95@#69PW[T^M$C.P 
@QZIFX<DUFBWZEEXOAM!S3C8H0X+42R<HD:Q.=V[!>RL 
@A.,URMXK%LS=S?]8!=Z_A,BGDE1378A9G)GGX01&B"H 
@RH$0ZYU40PNK9],&'_,R;!%P*R$T<MG'K;B[F217_V4 
@X87OK L"T-?'O@S/_-[FHY[GN79$4W4]6X'.B+.!$DP 
@JO<<3 ?ZOP(8'QA)_1'.L-J-:I00G:1/3M"0U+!";2P 
@[\HK+(5G2<:]"=<V4Z/@5/?:MX+^Y0,.\!IZ/EQYG!( 
@E("2=[OC>KHT53U!@(>+E$Z.,LZ!P?;XF8&R(2;[YDH 
@7*6EDV3&8:E\:A,D(".+DJLUW8.UW2!28]ZEL;$YBCX 
@FL3)H1F$71=O_X$INR^'U4I+KZ,=TK8.>Q'27H#@#(< 
@??^MYE8;F3&A.10M;[21^:#B2;H%!JV_*M*Y[%/N"^T 
@T4P*Y8K1/+H'T6\;@"CLZ,4?].E=BD9NEMZ )"913DP 
@CNR\'6B%-&T]A)6>7DL6_GO,))W5<$EN!-52$57E'SD 
@Y%D3@DRF66(M*\IIU%FUZ#A6.,EZ/V&B<[+*L24N17T 
@]R^_U;M9]N4-4-8V9LR*7\*2.M/$-6,\@0J%-,?]'@@ 
@W'T?G[M*0+R*=O+5@H&[ICG^:(OS.7,6WS,76=2-_&, 
@ ^X=X1&UCB.*(30N?+*D$*H8EP!?Y<#[*X+^0+6?KB$ 
@/[?Q0$H@$U22,A[,<IT;[KY5"<56"ZP$OXL%?WZ*-<( 
@*#3.2(W UY$$DR2[K,^KCVL%JFP?[5$NP:>CHW$SV&T 
@MILNM@F_1:J2"#QO53&<T8@O T_Z@;&PX&6H4S'C!:L 
@,]VK0'MC<H1M;U^_S4#< =.-M9MOE9G)2=.I2*YKP!P 
@$>"7:6GHG80Z9R@*Y 65-T[]#,,X-(ORZ?<B5RR)NW  
@']\0RWX=QL P2SI[\#AYYD*#_=^S118=4!HP=J,0HW\ 
@AP7C2Z<F\0@;PE<(OM'A%89$!E5_R,%=FKG)10. 'N@ 
@L[KJ5Z][*S>RN4E$]O<O?"RE+AJ/-0SV))AF2>3^QF( 
@V>I-@:X.X5<4P[<>8Z=!"0A.3)W&91AKBCX%UW[V'Y8 
@4WKHL-A/6]'1),K>6HNJFJ8.EOG4)^-6>4,PG1(5*"X 
@9 S2$G'JF568>(<W]864&V98',J?$G6U)L-UV+Q3PBP 
@N\F7B(+D4R5J'*D#:F]-4-@2^RB"#3P^^[4X)E\A;]T 
@VI]@4C6'M$2"@.6$%+4GX=>L1SJ<W789"&4(A^<BA/D 
@ZO9RK]"34"-(_XM;/F5W($UU5M/B$VY1V-JFBRL]O,0 
@K8;(R2;B335]5XKF%G-C"$^C7_0Y4*\PM6#S;YVD6K8 
@P--UGQ%E2_!@[0[KZ*$")#W0G:W=TY0SP]764(F0BE< 
@7\IBZ \_S'9Q:<H&1@X]JE+6/DD:W7<%XGWRY5)-I5X 
@D%[U/V$E&4LW:?<_WDVF'CG.QN;P$!3?6T-$$[1OQ$D 
@ DK7HFL0$I OK9<X9/]%]-[2$Y+@5!A[\[Q-A<\N$)L 
@3.-BOA81LQ#EQTGC\T)8@^.YOL\\2:YQ;;53\72!BA  
@5#O+>28M,"I"L+ 8&*68ZOH"Y/:_4Q$O*9BY& U"LC  
@G)%J(E1JMS] J #6V[+4._=8_?4UUBWS4FDN6WK. 14 
@9;-[V?IAU.Y*IT^=Q2"<4=,A(0MG6[H-L!0Z\#KG9PX 
@!;9&7@$.TD)!A( Q%*HW[),>[$P./YO+8T/#9)"?X2  
@'@$R,VI/C[;K&#8;QFX3+]XXT=D.'O.!'*]:TARSDDL 
@MPGI#)P,Z@1T_5"6)7X5WK@>]975'^IU;$=U7\5?;P( 
@:JH&J-B7+A6M*Z"R_C=JO\I>5\BR+53Q,C/4%Z>)W0( 
@T ?N%V!-0.FU8T'H(Q\(7]3W%+[-<QWS<P[]P&BJRT4 
@3O6J";BU>O90KE+BVBK='2?=Y_<H\)[JMFDUHO7\MV@ 
@S\J+E5\M(-%51X.Z.6J$^\T.E*^B!SKW6X9"\E K'R\ 
@4NSANO]091L(HX??IV\1OYX1!EE=Y)\"<>)W)ZP[CD, 
@,4.I0>K;P9)K>QYOD =_OY9BA#7^&!E_3S.P-X^SXN, 
@U%D/8GDW)= A^;H/5AFE@B(F4%2<K/(,/]2T,_$OVJT 
@#XI->J]ND8I+1"3R=U +CE<(BT!DN3B#Q&K)DN?HU ( 
@HDD"%(?KQF5?Q[VB4B/$&HDGI^03+\55T6EZ) M3,K< 
@>/+T;R=[=^<:Z[A24\"-\3'=*OXIYCL"+B/);U"X=1L 
@VZ\O#7$>LZ\,;43"K$_7VEU.3F!@'9^#"(:D="*H@1$ 
@GGGKQ<B691KW*O9(N2[E:!(/W\/&D*M"VBSM7_=H:2H 
@DSW+IL,5]QY[![(LB!M2Z+J_MNX#AC2!XG^-G[B'DP8 
@^71+ O$N.]=4<LA ].?BR)U2R2)C#(Q@J ':"CZV,K, 
@:%]417'13A&7N++"*IX<^<BTG+./'!X0XBQQ+B4<>:X 
@A=R.]J-UKR0TJ^$;<(.'_>-TQWP$JW8Q*<3R,>CSV,H 
@$3NE<O2@=)A?^3X:ACLW00ENEXBIB? ./O6_BF;2J!P 
@:8@R5*S&V"]9+KSSYC&4=94#\(OK)EKZU1FA=3XQI&X 
@@FL8\>9M,9PM;U=DX94I\,J%$KI.T<D)E''9*ZH[1W@ 
@0@H8K>;R)%EP6AT>OBG>&0.W=NOE&E-NB6?6[[#?YU4 
@$H6?4PVX5?X_(1YO' 4."[!4>WYR\#S,%8NS3(5P>4  
@P*@!<F2T%MH7A)M?=[>!WPD:#SKYL0.ZE&,:+!6_IXH 
@4\%&U<=#H,I<6PG2G6IBQ!@9[80<"/KA&8VM5X4#<.\ 
@+TP/2AT%LT=+!C$2BRKH0D49U'U>0(.:,$02-93XJ P 
@_Y/ ;D9UD# ]W3,^I/GBPHIH1W6#%(1KJ+"DA+4V8?< 
@77LX$SD79.2#C:O?L2NFA )JHF>"G+NCR[E*-9\^[XD 
@E\ECX9?I^F/0O0JU.#X$[]9NP*.C@F<4RW_D(9D-?N0 
@Z3:TA^T7H;.VWFP1A!E<XD"%E'XLGP-WJ_O3^E8&I[$ 
@,8&MRB0@/^#P:TN/'XMG_X-#F$>B&B8)O<(:[6N,]P( 
@(#*-W)J_]'D%N_V* QUMD,B_->]7;RLN CA^6$KIXE, 
@C%4TRYOCC<-W_1QV%5:-!(DGZF1\;G?;ZE*;7TV;E   
@_SR<%SYF;CT(1^.,BJ=X,.ONHA9*_<@D1S0N<D+R]48 
@U.)A&SM\4 "+ ILQ[Z1^X/O]TP[/Z04$97:D]@BU>>T 
@8]%Q'0&JZPCQ?((5DC#;=5U)!+<&JT!7!A/X/LHFG:D 
@,D_](LO33F*)#3-@23<1H\UIR R<2.'0&?886"\:9C  
@X2*VLAAD\&QL!+(Z6? B2$Q%P>]_9;8>V +,6U&HO/L 
@V[G+Y@,328AH-.>E]U!A&^=U)MX9V@C4P16%!WX(Y@\ 
@2 3X-@L[$=+KX$JA#U<YC(J%3&E'-97/=R[^#85:JYH 
@Y%]%-H5SBQ<N]N=DTV@T]G"S%_VQ2$"*L$E9N]8-V $ 
@(U9K1]GNV$4A[1@^W&SV?O_CK$UH#<8JK&3$"/\%$,T 
@3URFFKO4&6ZL%WZ&(6&R*/OR=+&ES,[D8\$]W#Y+TY8 
@N93F6O<J%(;H:=)/C'4D#L?#5@!Z#E=9!BX\;QHM7#< 
@HG+9;"Y-VH:6Z$Q.^UE8YR  WNYPQF-(@^1!:DMJ%S, 
@IP_4DL Z%K*4U;6DQ'!IV*$*P4\EB1D4?],R+S4N?:0 
@<F!7$W46E_';4,L_F 3\33J;#]%F/C,+7;#P[NQH/ P 
@Z!Y>/]BIN)/G:H)6#9RJ1UT(FF%-3GE-N._L8,6@):P 
@Z--I_8#3+Y,/$>31[>B-TI#Q@'E;.2?5N"Z0$1G%0(4 
@AU'<LOCN"@R@3<RV'GI-!*D9UF,R\:RA3+0IN<6Q?H\ 
@AYU\"6= 4.1X',9X+AFW9A10@W;A58 5P5X[$$6NB&( 
@XU(%I4C5$%!VE5:I-(L&,>>:T06,O3=R B'_&WZD5&L 
@Q!7TG+-N_H 1-2 H*Q$-LWJS'.I;OYFAZAI6)(F8EWL 
@"7$8QVD$IT;PT.5Y=FJH,JQ@\P.1ZVT]3LY;Q=QHXV@ 
@]C77H7E<"7[Q,3>#J2GEDV=CQ6(_9SZZ@2C*QGK1?!D 
@ QIR"KMC<DOHC66YCW'D&OUXK&B[]RD>;<#-[QCI\EP 
@CT$F%Y1J=?9N'Y:>0<T*%,696_9=O)Z.,B9O-?%Z:5, 
@BWT*AZ1)%^VE\PLRTS#MMMY^!SAB,-AA0X6<Z9&&/O4 
@TMC,)'0O0[QJ#@*MB^J\"+DECH3$GKE>J+4==9#^4'0 
@\6>!DYP;+4'?:^VU^DT_%#Q#"BJ(C=,<Q4 /W]0Z5T\ 
@CEAB@X:GL*-< 'VIE).Y6EV+,3:)%"7A'@F'.Z-K_YH 
@._B8$?UAP>^=O;:R= ETL#34T3WEUZ:>Y9]Q!BLE<XH 
@NS.]*CVCSPC3#7="[9G1627XUD2J?[#C(>27&>I@)Y$ 
@2;=S<V<:O; #(LZV(%O6*Y1QHW9V#SMU+Z,DN7K);D( 
@9$3<GH%S"=VED8OZN$"LT%2%])EUU!-37%)IEP<IQ(T 
@^F4.0PDNM<JCP\4T@OT]B%,ZGD6(%(H4_-78LLU YE( 
@O3+@I7[V_O&NAI&)_E Y@\9X ^C\@)7("97@7N63U@D 
@XZ=Q6?2/!7YPF?$I-B)*Q0U'/F8OUEX?PK*94+]\Q(  
@?MS2[)"YZ1<![^_D3LT;#XNR1E AY]C#$:9UB65+@J( 
@R],Q?"&(;?OK]#]ET_E[NFA?6VK?DXV@9\IZ*V6,,(P 
@3S>89%UCW5.ZGV&(TU'Z$CG^B]4G5=_+V7V%:!*'# 4 
@^H/[<5#-6!J#@,[R[ONKHNT**HI!=IC\'_EE0!]I?(T 
@W_OD-V]R#]"M9=K^9 ?]4Z[*H&CX,LIB(5_HC<8HDX@ 
@\B_@.0N@_WL/LE$:3:U7,NULW$'^SNX6&J?ZRO7@^YD 
@N%B$%@M98J\Y&:#-R3H&Z@X9=M5=V9?L@.-1)EM11@X 
@.:OAE^I>N]&[4@.^0?3_L#<*9<:=XXR9&\ICF]CZL_, 
@39^KL\3;,@Y7U6F1KTNT!&OS$W2?DT(=D"(TO[N2=S< 
@JQ,J3%Y1"Q I0ILQTN9A"'R9!H:/1V-0]&OTMX-K<(X 
@)<1\4RL=B*'@)L VX82(3*S4#U+>([BRLY0P& !+S?< 
@Y'N._I2B?YBD"!-_]R=CEU09TN3T@U-ASTIR<QN#YV, 
@WP8\0Q=47YGWVM^O,WQ@R4TJI2":Q,]^#IH>IL^:!.  
@HNE;+7@X3EKHL)Z[%^P&PYAI]OX! 5.V-P6I?#R^. ( 
0VP82[&+X&]+KH,DKO'TUH   
`pragma protect end_protected
