// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k1ckbU3gr+iOEzrks1RLwlBU2q/rG4GHGyZ997Ky5Yc406B0tUhcy2fQBgcS64Rs
1HOYR5FRECAwAX8ohlsRgWh0Szb8m3xmvGB8yGerzzU9lEWkBSNawznq12BMAvW5
ByUuVeLZYX4DLxr9w2DmiWdm8Po0LkScbT7rSVtfPz8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23264)
LyX+3ICyEdUp9RhIWMmxGFw7fA+SUxTs4DIcLN2KJ8gv03fI5hbk8BI+37js0Yz7
CKTqSPf4JRckxTgJe0V4eDCI1JEL+fBtDRmeEV/JIxToiCwoN02faaV5qfjjvwvK
vTrihInOLg+AR3Maweb9/3zGH9t5HYt9QM2PNdWnynB4e6lzhv6z/NC4mOzmHXDm
qCyDXqKVspAMlltNoyY3Y9yirT2yjYe2ZmWGRT+A2JeTiqBGmlhZgCdXNpJN8nfx
46oOUGXJQesNXANSx7HLcwGK0wxDe7Vb1Ucq7BJzNgStyWO98VF99NeJ2E8JHySn
qMZBn8mFsx9Ss+gY2wuvGZe/H6nzWXyRkKDBIU7SrRzVLwYY+DmGwf0N97PcyM9g
RIn+gwBw5AMbHKeK1Cnlm024cnYDDCvM1AuXQgfR0U/ZIvYZEu519t3wJStHDDmd
E14PbcY1nB7QabTES0ZJkdDzjKb46ljl1hdNEFe35OjHM4AEeNfG8z48YYr1eegp
5PgU+zwLBvuFqiXf/V1a82mWuXKr+TuBm1XGg5YkSSz+oiPP0Joz27HSuqiYxDO4
XMRf0//08UzC8Hv7ntCV6D9dnabnGggi+qYC/HVThROu1uF2kPRbmjbvUAiDdQFs
8H27W2xrTtYboa92a8KP44tK798dRQ538SWGfzRvVi+di/3AP25z63lGKQEivzk8
FHj76QleKG90DGomL7ccddotwLmK/79/IWeWMDA9u3ToKXEPyn6GYYG8D98tIcoy
CIhzQOrDfcSxY2va7a7IrScOU9Ojf86XrVUarA2m7vX1FT1N2XvQStIe4GzfyDDu
8cHwSXDK9+0Pr1Gg+nGfuoSuZem+skMlQwTAvizUl9oLGizmkPzY7s7W45ozXfQ1
6wM5cfLMh+cs3aKl5wk748fGx0FkxJnuUoe9/iPeQHo8Vo/KmsNMcnbyxBqNyvZU
Xr2+9qqxCBuh7vUHUF8mlhwfPeB5J3yVumUKCFgpFs4GJXRuTRKSxQunYP0nP/Nq
QAyyVXKgLR24Qo5cPbTyr01Jq2BPziFxkMsZCzlg5gZy75ZBAIh6/TG15BdWnd1K
e/1RdW5bxXaX4I3ZcTZEf++Acba9vYBo7nq3iKR7ChacVacPRq2nPuVYBgH0Yaa4
5MHOvSOrQqHFdVEaOAi6MalPJ/b78eR21VxoYjddSJXJR6zZNd0LflFMnMAFV4Hr
LxXpevfRgbLRhCZM16mYJVOZTdqt8C1EdALjFTMPaF4IAHP7izET+UQ6OCxMBhGd
L/aSfQ63XDY62GFGJPK0F7yVRd8MWwUrDTRlCQAwGmrlj/3esIIpU22j4t1dcguO
dVxvbEoPHEOLNxKnhNqr4GuroZFFk9nViWF5x6AL6mk1l+vjkdjFgdOPgsjmILe1
oo3Ofoquvpv1FMHwpoRohXJZlpICfseu2hGsNdVK7o9YN3bXLln0kDPb5ccvyrBw
zjbdR5xfESusKmzH8NseU8DwZCEeVBtQC66HBCwIne2hszfP/O+XwfRI74lTXIKb
rLoIxvtoESjlQjTohFV8eIufgWoks7lkZi9k3hsK+bKVwlvBVCNL5FbrZjn0Dc01
819XH8e7tHPDogWYqKVvS24vngLcYep5w2QC467r70JDKmHCPayOuiqOlCwemgcr
8g6xBrQ6AIot19o+7Sr4FZbe5oyExL+qze4LFUeo9tqnP1cr0mMmrT0hcLdBfMbf
4RS5rK3cdNuez9d3uCubolLaworW/E7TXkOwRedV3+E+kMPBw6RK4WBFuVi5YP+E
CQaZjsQXWbwSM3KXuPc4IW63+3QgQdn1tlXQLKkiZ1pQYaTB94G0joPDzrI8jY8m
MjFTuJlt0RGvahak9z+UzI/QzEj03/XW+lvmho51E6MAl3vzvbtpSjuMF32bL5KP
EJSNO3qqBVY295CLOw4RAgACo4bqxoZn51AVj8N5laUSKcibI5cwue4vfEapp8RM
Ap2FkBChyd6OEUVIILHgzZftXi+tcdPYRgtGp6Q5FRYjvzA8p0iGKRZR+796uQ0f
PH6ILUz5a32w6/UhrErci+h1eVSVUW8ZQqkE6AO2oiKpoNO6pvpAdpFTvOa17pO7
u/MzlKU4Eonvs589UYIPfSN9I2NTxozlhZ93AABcVmQ7CcIFXHSA8cL/O1Riy0LU
WWW5dsAcFLAq11UCYBnO5FWJ+zqmP09F3DCztOcDQ1fAbxTHGKywj9u8JJ+DaETK
dK5oQVNqrJe2+94N6XYhq/JjfhVs/8oVkSyUWqNHiWw+qHwh1FKvWZurYR/VjOFt
Ales6UKjOXFVT03WwN7tuF+BKbyzkhIm9X9zgycH4M1/Ax59eWlbsGGF5RAE8bOx
+z1yKyJAwnvea3zykAVOOJ/M4KwhMqas024Qw8GpHOc9vJ8VxnXucZmyj+eoKLPA
Kf69FzsTdk47AJ+bV4UTDuT/7vESoFwxCaBh3+7DVEEsIAXeDBZXo3PjkjSGYUzS
9viVWBAsy5yQcwB9fliNR+RcWYyyxTz++WMqul51TmxQx5N5CVz4fk3dygNiciRI
HCIVWitRNJhsjbw//p1I56mmSzQGsOYtkzoIn70XKFnfo/9nYDpqzzlcbDAyiyof
h1xGGfsDEXvHNSJ/9QCv2WQVc7LQaPlsdev9GrKilb7i9nuhYzuDPL+aCM/S5PiV
qx02G0QR0KaunaKCFhuTUVgXrNwC9KCuECWvfuV2TeuNDNw2oSoP1uEXO17djE2E
puLUnwvPyyRCm8E86kzlcIsGvdE9iUnBHkg0ckIcjVVNqqLoiKJ9suN9Y8djI12X
cvVlAuKrwoV4NLrjA6DQEjNY81sFWHiZxsHlpdjGx2ESndgZkaoLB8cgWW80gP5i
IgwcHV7zq9PAtLivxu7CAvTGAFByGgPA1i4oPjZfsn02xcYM0+6DB0tY7dnsosLo
3hoqODSrnmXTz3aktv0Rkuuuh5zqEcs5teBPVU1Kw4pf6hbmQqJLTYOnYMCcfEnw
73gaVUW4reGtFkDSXNOMop2cGGvP5263H8b3hTT0GcMZ+v1Z1psUrw4B4MlA0/OM
nvZWgcA3QKxazHY4aRcLqsWq8HC8L6YkWp4viNRJyOAng4x7u1rYrbZSY+p3g92C
8hyQJ8l9EveVDfbbjQFFOe3Tqb09Tj6N0ISidVcmdAPM/4RleUcGUjpSjyEZLLIY
oXqB0gR9oxBIHSCvL28cjiNvMbp2b/uUKWQ0al6TZR8ntm3XHSI2HO9UeirkHetw
ksh3lNHrv3YqBPE4+pmBVxHT/LZub+Batacwso0lOIZ1Th36m8OpFzf1bi8ZcjIv
BAbvQaaFf2Rdg0cxlBu2i8sS3qvOAHcReJizejhCxVzs9Bsj3/oLhs5h3nPOUh9i
0zni5W4rZPKv22cQGdMeyaqMhGNrTiYV5weerKN/pn3XkqkCGE+bMmF2i1nd0lqq
z5decUSqb9NpntF6V+DbnqBhDSXAV02iP66oh5WwCxIc+csOJRBAVE9b5QodTZiv
Jsa674Sn2oqPBW/q8+V2dgo4PCD+y5o/iO0NmjXMfaraIz5IxX1aOLMtiNtkra/W
ou7LvHT0Fi40MRGq8gproOveBJhD7V22J7wvagM2/X04dX8rJY5XF2dT6o11ZK2J
qzqV5/P7l7g1Io1AOuibkkTUvHGWp24NZZUZkWE5rw7IYRSKAAr8JSxqS+5+tY3b
EwOyxfAEjhdvXdEuYl4N+O7v4K5dvhM0Pxfm3DmU4M/GmoBfuLLzrWAp6h2w1RgC
Uk8uT2hJKaZZHw9sp8/k++i/zChcXX2IJncRDnyP3utoTk6W5qs7AUIqKL1w8722
dL/vfv7kxP7Uezi6YG4zkwO3aHb/gCXPiQePAcqwwTLLaAc7kQDQeLpfPqXtjp6w
ycy2sQJS/7QqpE4l2NDQzM/hoKXryGoiS9B0UUo0It0d2JyXSkTbUI1sFkUOBVet
z0pvxoDf0Gs1f+K/AYFl5th8gYU9InZfx5rVtIMInyvRQJ+eK0HrfmaXCVs7Rc4o
yhWaxDbGOXsNVMpKBsPcwT9ftfzaErxYQEgHqRuCnrvCTSGOtp3oJE8nYu68MmI5
IZ1VgXyE2ZXVpuA1Xkrlkk5sRIFnpHNxQBDOU3Z7FVLlYvvduqGvgv49+Mhf0CTc
Xv+Fb73uJJxn0CdZAz3utJfWM8oABpCN1hqgJ1UNXkWv4rpGEFOlcI6eEftxEP8I
fX8z0FY1s6CcDmumIUbGgLBV2CIjiCWjPSsV2dR6yILl0TahdMCDTMAmugBowZHA
trVEMNybRqVMabOTJI+W0RVv0FKauPl1hLN35zg1GbKf9Ls1Esi9x+KDMnDyHlLE
dNCp9PE4N04wwLirYeGX8fUzWVuchw6RuPsyZ0D/6Ec7z1usSIpsccBrtCFxcLPp
RhjR1jTGuuVit/r0fwUTizpc8n05Dymkmij/hDqV+eIKeZx8TTNarlSJUfRsETxs
ygAIDkrrvfeUZj/FFXvYFcGxwFCbSIQ3gdesmvsdoH8IjUtrhwciiJWujXM1SLIr
GDILv6t+D9nD2YpF7XEsR+epapGowsNwkGRXQcv3LbcAca69zVuA7uQi6+PLDpUW
/7i1gDiGWht2oGqXk0ZJKYtND+gnA8plEc4bVgPQO+drK8o9dgZ2gn49ayfqzDT2
Vpm9oFWPH2jffhlxu4rwU6nSonOJ+dXpXQESzA9jf8NojjTZGPir2PR5O6fznrB6
1HE83zFinJ2EtKlfDoo8HiHkjAwwmrwZcdkFutQk6ucVym5Yma4yW07fnybPwCVZ
mVBJbR3N0WXLwFId3Dof39oK9ifLNLzeACsrxOaB8oIiDqAi9DQkV80sUEFtSZeq
lIsmRElTQqYaLhfgRwQB5jJQ/KPkYWlC7oTyUD1F0qddgaUwU/s+zALL3leJuS/e
9QlzGTCKEgx1SOeJK0hAUZ5YNDbMCTEMy5YdFgMGr8QSAhIrdjYaG8NKCe/DKPfS
wvbB7g6QxYk3D+0/10p/iKsq9Wh3f3dytwM9NEtPQXkAcSy1DIGZUksPBPzar7w/
DWkA9lxR7G1MyjeCbzFNm4HrEQpfahj7IkGK2vo9svzWGmaWXaZsbK3Vd+aUVPlB
TBiScAAci4i0FiYn9+8KY+/Te1WqjSzOe6YhcUxSz3mhTA/5br6s+nMIpcxTshvr
zWs3w65n5KDyIot/UTzdw4unNEKGyNHxWqKACkzCaviCOtITxawHeBtppFRv9qof
9A1Q4cSrX9QQtQhjXxh4qkSNLSzcEriYt99DMM7dMVeXmZD+jvWsx1mX//a+rm+f
CFSlSFGovVK7v8pGZC54iVtzibnB9aljUiNdYAVSNvEtDgvVBLzdm6Sg11aBhto4
G2sY2rvJuJJQslf/7/SxOuaE2wdbKmYYOj49T2DtNpZk/PlgVDN2FyatwmFcMZrm
whQb6mDMI4LJJYePMwJIRjx6YKSZw+flxBInadCeg5DZJatdZmNIKZ8GlY6DbR5a
xG5fh83b4K2GgN7ho0LlabaBxKzlmbzBq3Zf3PIpDROY2PeElAs49KYcxWn8Jf/B
lTJRDfC0qw8r/98f0VO/qKuvYlf6STaeue7szZyp9fxTerCa1G3fCkBoExzV+2AJ
LBfBJ++j84Web01iP5xgsd5clJ7G2s51sQUfPqtlYaUAOT4BUHAJsm0nZ1SI5Kqi
yLE/eZ1qkiG7UIZbXR92OWKdhYw8QEljq6800zKUBTt5zN4ge7v7Vjw1dE766pEe
BMNVKXofYlFKS5c3e1BD8evKr7E+VW/1lgjE2f6G34OxQ3hTXaybroXZ6G0++v6p
k/IQai8VSzHFp1SrOKKpmUPiZ5c3+3xo/mHbWvmdkUkDFGvIYL/rdGpTxfIczpJn
r1wPP+nEeh3yPTqf5lPsGLGOiMHjUF5ZIZYknmizHayzx1veXK4KpgbkBTsZ63Rf
s/bfhTIlC5QExKEpGdxwYwy3dSLbETiuQezRO6vP0/DAOsh8G6329t8qVjLm5kas
Hfk9CHNpP+VKbuKWtlpjfy9B8KNNYnuct0j+tI1JmBoRawFR0pjefVMW/vQ9I+JW
XPQzZEOFSqSSEa5yB5Np3H5+JwwKwIlXR5qWAKohsfK5vhRcXnr+dH2aR78cGy3J
OfkVwSZxezprTgvJKWv93wWFBE61cdNpsrO5V8hArej8Aljks9vdI0mMZrT9M0IE
l3H6MfWhOie35ChZe+eP+Yq7EjsvnhmvWWONwz7gif/iHO81yp9Nfq2OyhSD0XVL
ZpodzNyapq7s1DM91i2Y8JTKQMeD5O6R4QMtQLjnDL6cutt91PwSk98s/+D1HOnq
Qs4vUvZboYUa5/0mAGxT0+YF7t5b7Mm1e7Lg6Gg3EruAZKK3rn+mw9NuCJdspprU
LIb+ObaTxbku5ZdGtommwh246asN0B28Mlvr2mJYKdrtcHX/xPawKy3PgDBuIS0E
GpRWayxrjto0XwUsW/vBTOLbBYq1kXzPTHZSQ8TLfz/J0KS5O3Q30S1+57brgerO
0Q44xVwxyFXCJxY4uLjUXzbt+UzEL6KRrH4N370jgM7haSu9OUkvKLTzOgCsZjPH
wIL4rZgM7ozf7Puz10wn4NEontwgZlJwk3jmlmgL+Jz9OXD1TjfB3KncDxgPxM98
8b3SJPN0OgiqKcU8eMY4fQOMmRu+83gPWoLdcmBNg7bQXK/2+SjpWSsfBxxISK5+
CqE7B/AqDt8wnQNexsdDIOswQ6/1JTZ3xwnI0VbqQdKgTlnRwlHD/ZUmxa8aXwHk
YmNXzbLepRZSzrCmucNBFdVYy63VmqEIeLB+fGVq6DS+QtpOkZEFFA+0OhlJopdr
rs+ORWzxuwLNIacZZkVpbO8hfHpEIONYSdmMEzrUJDwv6JLnRbgwSjG5NVAv626R
+1MH4AErZOQhUPNn4cA6x/NJLOhtrLZhmB/bQjn1RvSph0hcrC+6ilMiTgnbE8VQ
4tQdZ2paZ2i0xNJfacQJAMskSm5zisLcyJMoyYlDkf3lNEcniSkpFlWXvEDEoUz1
sQt9yJ6F6jgRLfbk1sU06S/HgMqz1ftvOQa5JsO0OWvdJo7zZ8d6jV56gEzGFsB5
im2nV3BAodAaVRztEzLYsz84wxBy4h5TitCbl+wdYVGUEqZrKZHud1aoNZ449rXP
ehNY/H1KeplrJ0kvaU30JRnjYP+0rG/Y9uSpBE2Ms0JCRKMbS/LTKsyDRXBbF90N
iyvecrI6ii0h+sNZr7KgYlTHQYAZ6fHVXnn3wazDslrsFuuVeB3E23pLC1WJl8p3
E44ychCNclmsIx80inDKeOvXhGfClsv8p9k6JjtX/o51T3vajbleCV+X9C8ScLNR
hp4/L4uajMuCgoQDGhZfLRusHIQ5HTBkHz3tF/S9V+2zabZSfgUTL79FXYEAwXHX
nPnrtxAYWDwfzeDflgKNKE33D5OHM1+Xae7hcg3bv8vr27kXCi6Rg5qS9AsvmTG9
u2ZFvlmxkPJTSv0Z3NB2DqxBeVhjDXFdy/1WNwnCCzJ4D2oblhbI2teNijhfi2es
Ay2kWQteL9lKzz+1kP/zerAqa0q435HHHzm8q4nk1P4apm7XssUk9bwYPvooy2nk
P+lXu/pAl/VhtxAiXeLW1+WJsGkNN56ChaJqF+AzX4Y78Hd4y7MCSojBE099XrLy
JRNc2SvzERhuZsFTnNxlDgguW/MgLA99g5ozMGrfoQ1Cg+m+K3r9PSuKrYup7kZ0
hBUoOnEf7/6HzQozsIkAETmY8QkjGOFeMFhZtu1zDDztXL5ZhUG6KwUWRZ2qO0EM
aYl9S7LLHigsN670YP9LY7+Hcdt21jshT6ij/O10qnOBQj7EZ1aKu/xLbMR9Vgg0
8ZVYM2+UnRXHfncO9niFUI/1xaJsMAQPVL8Fd7FPCOKuFwXuGupV7CYkYjnybxoW
bQD2FMaoBAOdwc2uaxgMWlBqOh6wdJ0E4b9gX7Ogn7amQboLt1mvcjlpHxAUrhRa
EhGxFysL2D6AE+utBOK6Wpcxe5AV/hwI/KmDhEStrLTTg8sRFwRA7jn/nkBstPZ3
9EXEfID9LRNi2Oj+pkF0sW8ME6/USZ7Hxzsgvt7jNJkytlibD5e6B453EqEPBD5K
hEqF3RI7PtHSBV5T519NMpRfJfSAQxYtFrUzE0gut8HsstDhFmL+q94gonrcdQbV
O0j8Awv2suhlazvyenLETFrKI0ti12u2sSGnG6Z5aQl7ObWtctj8zWaVa+f6WW6W
QhcKxTxBy+1oi52XxJi9kBjh7Gpv0INRkyICHf7K3/gbkecQzPXYq3kVNt2PMeCk
zZebVlOH44/cbAqNMdMG0I7dXzvUY2ENzhce8M0cljFxbPnLBvjexB90OYPf++9J
rOSYpvBA6lZCg4mWTrXjh3mCZZEyngwck7FIummP7SejOzyuu9N+8RkvTiRVhXio
qQe6zrRg2zO1TP60r/TZ2cIrMLnmx0PQHK3TikuROoxYxBeKsfLmgHfsL9BPE2EM
g4dtrSq11ghRs0R2V0dRrLQIVvatQJ1BvaKvmGf9PAwTT1/TacPWujWJzC+I38JD
Iu6eky8XINJsnTbK89OjZM3o60QR8zP52houe5mnWSD8C/0u9c3zfp3pssEVEDkw
NTmYNse2GggegReLLgI5lkAGgs0Pl5Qs/fV2TCx+JI95XOriTAl6oQ2EvVyoCfNH
qt9DT0lJk3uq0R0mD/rKmc7cGTUnzokXpXeQZVj7PSdFYgyPTAuMcy/ktxWmw5Fa
4kpxppcHe/aTFXHSVLV17It4U7/LdQwKt9YpifgkYr0+Qj3WPgavQzW8vZf12ND/
0wwUtKQkDvI9RXwXUHxU8psSS7Zd6RKLIvOJ8cR3y/JQskl/Dhg2DRR6Zhaqlobs
/vVkCUVaE8zmMVhkyfh0NJYukqXQhfbyYkWASjJO82Ofv9ax4kfs108EwgsSbHlm
jqMoS95hz3FGajkxlzpQZ011QDFqCbnSMYtQH0w2EcCUOPJDdYlMYigphEcOn91u
zvV48UBzU6aOHoOJ9GUZOtS1I6xHmaUNBof+WwY5XrHMK9Ds8QRTGPsln/XBjgAd
hy+GyxZ+oW2QnJZN6BhmD4f3lDIFuKItMhzHao4SL3xmYhUfT+dllI64defP/wta
JwX9VAR0/zBb8u2E1Ul0SsKp5MbD8sh2zA2+bMaLlitq5lHrgt8f78YmsxflPvCQ
vy19AIDSskYe1c47IAu8HoTrdg3JyjBb8/IvLLY5h5hk/VocLLp68yBSyOFplc9k
yRYspOu/1SKIDZzYCp3B89jwT97MXasIldeYMKAQCuZ7MsWV2162CWmv4y0ei7ld
6XFuyw2QfDrZ99nrxmrPcR1eQModybZKWrOelg+74ehf4oktqx0ISccfReKETvtw
l3J5Ws8SBNSlMaSXJGi30Zm8wj6RPcw/UB/XwvHT6wpUbXevjCCK6TQCW7bqCB9x
elXOXsKz8B27MSHWCFIITXp3c6pdKkmD1XX11Gb0RyVE4diJQZPdwiJV2njw/gbN
VoTLqiR65hl8aCNb4fxbMHBfKsnUtrOl5ZhMQ5iXOV3EKKAOdlnoaiEyKl8mWSKx
1KPzEVoKRdn5x+cUKdn9JsYG/P3Kf7ICrHRwTs++7IHOShPYtmIH4+CtRVs/EfMm
pGX5SorftfUarHkCGUbV2QoZ+AnvPeLn1PaZ4UMqcIsqCZuKkwUUAK0XORnTRLb5
Wrms2e69Z186KejUfZREhKO3l83Zu6+rj9xfNZb9+4RQG05QP7WMCeTNKMk+8EZU
WLZekYtrjkUIddFei6cemX8wJ0JoTAjIjH9dTwqigmhRAYxbCXYdHVVTCHS6FpM9
y/7FPcxjEf21j7C4qGQXg6c72V9YtAwtAzPYv8qNzxkbYLCmZvmIDwzJ7ehpmatn
0YR991eeddF3pyrJZh2re5ZHLnjPdMmas8/lAsKbqyW1u1WGnm0t2wYuvegnqJ0k
sNts7h2q4j1izomojBYcXUaOXW2XMqfFsPwlZaNuJrvXRaJ4VmmxOYRiKhxE4cl5
FPfja5IFoI1XiAoqiQbLPSskUrRnUTYl0McrcXU7h1++nJz6WOLcwmZzCWszb1UH
d/ik3bcxYYU0PFux8jJNc8FcZsfxGQ+1IsuOeAXSpirDcvkEvo1vvy9hI26YPl+0
VIE2x5m8WK5WgpCQW70fpgNLdUCNxAQc7+RWgfbVmBENwRw5l5xkiBC6Q+0J5SSU
FqP8oKh+2G+JJnRyFWVLcniohkSKee1BNsrv3k90vDoSVbPI38iI2GYL8b8hIqeD
PCtvexpTy2n5wytyPVGAmDc5i7gG95VrGGch4eCem896rizjst1cjj+uGSzApwjh
iM52SJ6BRlaB3vtSYwsPrJ5hv0V7u332FrszQ7LkanX773Fka+0t0I0B7nuXtQPU
b3WkV+wrUExjP7WyzgWngtWfN3dfymp7mEH0MbvGrNl8uvjplgsHpt0P78iS2gtZ
eblypIa2tbd5LopmRjlymBcYYHHzYr9paSivPQXKmOuHmDNIz5XQ79Vs6kjJcQM+
gxyj8GrQvRvwUHwjyx33lfoOm+k4o66/5y2SmNGrqvpHpaNetMEAvZErQqxsp8wS
5z1+84hCsmWLWOufAOpcWwY1sR5bgg5S2hq5E9DFixWelO5Qr4KZPL3NyJlvf6aO
RKFYXJ2uP4bs4FnoYoAGAVG2i64JPNx/WG7J1yq4eW7C6vGIjijrT1OJjetDQaTx
OFmkPt+Lugw5+1bGHWV8aoYq9/WwZp8XyphASN8s4rVkoMqgiJjDgGXTkxvn1Hpw
gZUf59jcEGlHadhKhmpYBPQUy28LtXMBNYfwCOKxwhy4g/onm3O6gjogxoC8HOr9
YazQLRz8wUjQr97PDWZ5MZiQEwTO3qbBNWPurmTLr9vVQE9JZltPctr2PpXbcrTx
xB8+nhoqlKF8l17LarOcOKdzd1wvoABFXYwdPApAcmGgH0NnsEZ6Vfu7p7Wmmz8d
gXid3An2oLpWyHbQIkC+MJ82ToM0+RsKvszz+/5tKqDV1rOFWewPmK0oMBQfurwl
hkxTNZ4GbvLzDhNSkkXHTU5sDdDE7WX1ImxHUybP7haJDv/vOK5Jl/zEBaCq47ir
XeXbar0ZGvGWFatAW2rvCn+vxfFxeM6g3CBp9erBANLMnfOzWQm6u9Eu1FvL2/Et
xKusNdXbxRNEDZ87ZPpz0xjuroqAzyWLY1+HUSSaG8OKicLL+g2xbo8HCoz8CIdH
LU7zZGYwtMCQxY+sQHP9ipR7dNGnlOtRTROFo1FLBFRqKQ8XtY9r7D7gCGNDZVIv
6D7R5wfmPZgO0/qhvOBrsCaBBk6eZ5tpSaQDdh+JAl478LG+9XRkgcqBWmAc+23w
z2mU4gJveKV5uGyolwQv8aujh3UzTYVxs7FLvJanNIE1fKYAQa7Aj5Y2EK67VuCy
idOd/8vb6dZ50eS1aCw/vNcF46eQxc9Q5PbF5b/ER1BTEnzcFDc6yUmE9Tj4DKzp
/WcyRy1lxK7NE+0VlHplcjMgyH7tWfRIXFWItpXPJDhEatkkP0VBhKClUzsEiOqP
c3GvaQAFsr3Qcl+BtWzlJLU0Koh510FzU7gWTvxIDJBy5HYLhgoLFR2mFbFrJvl7
fNgnVCnxCmKh7oaoddJYgV/KzVvT8dLl7kTHhRWaF4GMRZzsBzwHheXepbJguEAD
mxB1eTF+ZMgKH8As5yZm7qcn6nxZlcajznlMKZ6PXEhh378HpgmdRbY7hms+OVyu
GqSWt/Uo/wYRb4A+Bg6gPoSusgxt5Ju5l+PZGkYVxwR0tlemDt4ZQhbPzUOLMyzJ
9wp9+SR4G7edujQIk/Y5/9F3HfTy64/uubXzFA7TFi4a8vFMOw2pnFNRmK7NJgZc
d6yQy0HC7OKlg/oKTsIMi/a0PUnqCq3r/NE8ZS8dKUchWyZiW+BSsh7wSNB2hS0y
ksU0eXld8SsUSjwO4VDkA00K2civ8QX0raePuYkigzyt/saKZSSLtQAg3YvneOtd
xs6WsynnSB8e/0QlTq7MNdip4TT60iXtimYPOCE2/Hf/BhAC7IrXLHGiZ43hjYo2
FTDYBCOPmEYJZlMBWV2LbpTO+qg4z/p3t/n1IRisPKqQpyv3yeWNukwpT8a0xIkw
Q4nXzdXUu48/hwk5AFG4IxE2b6UyJLDZTIRF7p23kh9WzBVTjvJbip9m+47bDtXL
OSkC2kio1uUPXz8wiAlJuZlWeCku9087+SyX0SaMa1BazAeuyQU0lim5r6NDFUf2
JNAaTPwpxu5bFBVTNrgrPzs48taP11mJJlzewBxpVF6PqXgxsX2JqYT2Ue2xbExd
8dx16CraBelUM7Xgk988pQSsyhgU5OlcIib76G7ckKW1zYdq7FbN51z5c2sKLeRq
esi7nZI5n/DeITWSIT89POmr1aCNxBsPj8DJ/rC0dvTSDbsSxM+OFt7JgAvLd+bd
CCCwXAA3OFOGDKcymq+OKZStsoh0T10OJikW+ZnRO3Li9D3xNVI1ORXJfnbmUKdM
BDCQh88Me5tBTPRaDIy/8ZfLssBU3ORuGK+UghT639RW7YHwb3hYeuKma7G4HzAz
PIN9tuCsNf/Sijj54VG70DeoMdvruSUyUEyBP503u4r/pflA1GYcMYwLEn0V5Avy
ibb3Tgm68s48fiR5kLqVlrocu/BweYdteaBvYUDm2o1VyBc792KOyRRPxewC3Ii7
u+2OV7dCS4zZhgKmgSChcVASkgNqOX1KrX9BQRA9pIplromDAhwpTpvQRBcY8zft
fZJayLJjq9W0pi4MlnCz0tjabqToeyhiiSnxdT2zgqxMsDvlVYV01H5phDcuZ0Jr
M/uADtjO+e3tWaMNtvpmKj5ExLwRBOuzDs496EMU7G2QNpeXsp4Gz6PvIBkSlW8P
dOSE1Jfz/pvYCWwTTTrv6IxihLlWT7gMhDACnarpe9iB/Kc2FhgYIA8tSdhRmiz+
S3fivyjdcFw4eZogWu5RUu63YnlOw5Ins2X5p3ZK67tGPU0AT/RYrxxYMDOoC7Er
YpQTB4OGAqlyFiiDVygdOWa41fE/YUncVLsXmChFlF+2SHeV7GW6cS3s4Os1vBVu
QT+YBui8bAq/bYPEpQaaUwyBwN5n0uZPIkAkao50+s78vPFZbIkHsAmjXIYQlbF1
tINBp/g/3648sbvPpRk6OtSKhj7yH16/FPVJZEpmnq4S+fAcjLB4KjXD+TdbUIxV
5WBKMxrD767qMy3+bUbklX//nWWQ57CgrWxveLod8wJHH9q4BNgcC5/fhhhipv1t
oVnWyECh0IIqqSkUWd4tpIp3GphIAKyaATEbd1ApiUDPAUtUC/fwnULhjUbdx1kH
aCLlFBQErixUAjVP3ZcRBvg1EdNkFstzhaGQzkOcqkQ7D1qNH1ehFBZ+q+6Mrph2
ztuLV5x20oHNo6ZLgB/8E5mTzDG0vPAwAE3D26bfjd+J90Wiy/ngXfmlLRcxZ0cR
l6W29qFrfzxYoT5DvxL8X29VVZ7yWpAjQrA8Vm+gHrAYntbBx52jFECAY24woMjh
2LSHrVPZiiPu9ZT4hofjwDAcpAbh07YXUnq452gdGUP/B4Q0qIgc7gu+ecSqpk1q
SmkmfJ549aeP2b0RsGQFWuf66i4Mkosbm5Vf8D+wv8Ja59hJ3dxlUbOiWssQnGiQ
WY6v+fMH73+My4A+PaFOUleu8J6VT0kfml7xUuh+hj9Lgsl//5729/UzB9j2c5Ka
Ws5YPXeE4xhyYWt6x3ELpjRLGuDac+z6x0voM+QQJMG/G91+Fe8ws901GfpcdF0f
NstQu3Jy7sP4B/16uFP2F5sFM3Y3zpdgns6ledjfBrhLhyPcadXJw9DG+TOl+3hy
aJb/gVAio3d82mg9WGLnuB0QzZ6/et1aXiRYwN9Bg/UkBkpEUBZTAgTNLDrRAy8d
xUpMOrZITyct4OQvJ+hL4Lmjo/oVPetnXz8mVJhDyUfpYzVdXOBtkb8whoqSiG2i
FRARybdKNBUUf6aLrE6cWUeh6XvU4PXUpzhrrehuBK0758ng+19eyg6N8xFcyhqc
mpCI4kNVP0g7q+fWT300fZg1X2ujhmYSaNuyNL23Noh5xSQP+z1zvYlvVNeiKvKx
p1QmNM7C4Fy3YPbLvguqJlFGBMsJy8LZOQCeRyV4C0TQ8gZpqxfsOmBLfjfAnEws
7KwB/p8GiHZLW4JUgvGPowUW9uhFtepSz5WCUNnFGUPkz4UOKbrxXs8cbcoINICM
hzZyyG9nj/2FMPo7jsywxsm0ce3EqH3oqdrS1pLKXjrLpLHhxlKJObgRdOyme44C
DpMyxO/ryxrsuKW8/kW7lIkce5sEBjkuFq7MrerBORpapadXn9JhvSGfUU38Xr//
hz74amyQxQ8SSKtfBED+3TWnBq8fLKhOlkMuIccLSzXLv1U8QiE2lrWjLxSTTL1Z
MS16MSidtG/mCsbXGUMz37dQZOjS2MrnPWCCstOHZZYVCEkT9nYE65QYlWkvmxop
nQzo6a8rPrynppDMQTSl6ToLqc379dZqkv4UX0rw03dPDg9uwW/2ngQM5RWS/vKi
BQ+NE0gxp+G6Ysgb3I4mr98P7UHCVDYTnUijrU2dGNCcobMROrjFJrpBdZCVmhH9
ExBPTVgd2q7Y/AjPFmBhXbRX/bztshH48NzKvqgIoplqKfHFc4myU8bzhfmSTiSU
i29AYDYpcJsMu1lF9PUaP46d0wyrJQHqfwQlYVsM6/UdiJot9wK7yjd41Sg4/l7G
655Plc//us8Zpj+x+Es10gO1evG1Qqh2hZXTFxa61KvZPCscG/bRqVF1SK6w+5wH
0aLH++e8jMFWuDRaKH8LfIXErgsCcYegaJ5K9EHFrgQcvC7Vk29MyNqXSDZhwfN7
RlciTb+x90WOtQ4Dl/w/VNaBNPveoBbtAwYdh76Fd69gKgfL41tosHiXu8ztwspj
yNHtgkt9C8H+YxHXS6ZulDRmjxBWvZRpReitllaAAs9E2p6VqOXQokq3bFJGp8nY
jrn7fbBJ+mKPYwGtHgyclEOp7ZB/ZajumBtb9OYd2J7MQyTYrZZDpMRhi5y7+HfP
25jGwWTgXkd/KiGAklfUieHGhW4/xPQGLe98qu8BJVI2nb0as1RacE62ki2IRxM2
pvz+7C8++pCi3xi2KlJv4kv0ivvjp+J5BjtE452qO55jZviz08ObtUD66eAUTJUp
6gYyIqaPlSh0ZUbDzRQQqugVn1E4nquXsui+XfTass/+KfNF020qiaNdGszSvuzE
WQ6Usvsi5pAucC1gGz6JMsgyvD+bd2sMtAfoTMGS34slVjyQo4020pW4nxf1O5N6
Op/S5uIbjDItPtymBsiP/WUtT5N2EXH4O90i2aFZK4iLHivJw4dKHzrNMDRYsTab
vgUOC5VnA4zpzdlF6vh5iZlNUDjdgdDU4vuBWqzphLughP124lHFmrkYLXXX8bM2
JbeT9b89NNnmPW6pgIAaifoM57e8pg0NCWaosaThcZoKSqyVmIHc7nkU3malH+s6
FVyasAn2f3mzKdz3d4bO/Ih20g8muJImcBisFdroVDk6kuoIx8pnuZRWDBqCbfHk
zZgNkARtj70deHOtr+DgtnXo++rVBHyYNIBlWcNRdcQlwcUCSMp7iR5CknEpSFaV
E5SJrMYmbn6t2Frsa/NCsGGIc+uAkfdchmREOJ5mn/uaNEwMMbASCGKE/8OdWk0c
3N5QEHxIdtufV90rdTlTo4Ujpjy3pMrCs74TeiSjtt1mn3M/AkeuhvR0ETD//5lB
6DQ01xvQoyXfatPu3Pymp2tIv6UzfQs/GZJdLt7cqKtzp6bJzZant4AcntzVjXE3
9mN1Dx2UmyQ6oe6WSJBUtexBOo6GnMRn7jM9u44O2bkdfq9pe1cxHeJo7D8HGMrN
r9AjCA9r7urJ9ic57kskOFr0e0LiL5764yBK8qPqZtBWcYYCwvRXk2Ba1ZKRiXmR
35rzUWoj9FI/tE54MuFFo6422v30hVvVo7r/qi7urpk4JW7c0KoeCqpkqJwXgjES
xRckE2hiICBXQP5LlXF8V9wDPhBF9Rgf2/oGR+N9kyGOIN5jUFsoyNRcT6pGgd2T
aKanJ2XyWmn+4nbPQo5ibtvQfoW0KpoB6oIcio7CwkbyYl+riXRTLEP/1KlMM5GN
eJS4cmqMMjSQEOY/Y/8tGTwD8jW46aBmOKXMzmfoo7CJZdXjKSRX5YgF9A6UCt3J
l0twg4dAXMl5xVX+4wcB8+y5JHQFQ9NKlCm114oSu7ECk4kdVRT6Pp3bRVV6Ta5B
h/kbDsYtNFD4hHM+ZvgGBli2x2jA5viPOYd/ZiSl+fzkPJOwrzu1hUSLSw+kJ1jE
ffcPw2ooebBrxY1nd+QUm+NwkJVHe2W5qA1xLvP9X2ZavLgfC+w/ItyKuTYiupv1
ULMrtVbJt3Xeg4TKhbTX/44mdGJB7CQuRG9o3Kps7wPUKQ2Z2pXGqHCKmG3zXJpq
Af4/Muycf4vF80+oA7/i3f778tDiy6IC4RNZWdnZyxXmYFPcOBWPxY0dKmPpgJBw
l+LqCDGdEROrn/bIYdUJrL/OMWLzSpbX+4/tl0wSaTqCT7cU2GGvQ3ezNORFUOAR
lWlvy2gGdLrRnkCCAVGfUdOUKJ3HlRwuHCBfkD3RWy6zOYAOT/jYguoVRnfVkZzM
kI3nElMBkYocSeWKpdTCTaxN/nYvBvoJhG5YCLxLYSWmSQ1TcZagO5PiNkAbHBgC
iDJQV11+NWKnMMCT6JkNArjmK91ij8amCFCsWOoQbNYRx3sx0DisOezs+15KpECw
TBEnGL6rfkpV3WLnEOnj5M7qpLRMAJtABehzXk68Rh/erOdwpbXZ6MrVqnHQZAUk
FSW/fAt3cJGdOxD4JnukjrvFa7ELJMeGQyTlt+RSU7UQSfmXeJ8mPijnH6TEBnLG
Zf8ETw5EQbYpfULQnydhrBpGewcaAah2YDi5Rz7c1+gYMzRvbPuj30ZO1AVX+Sin
1N6y5zqFqaOL5TM2S4rR4yGcuojpxgSgKjXSoC4IZRt3tipGY8ZE+Opywz9cnN/G
GCKAMN9Uwsbg3xCxIjhWZn6f41m88Dw3Z0KHa94PRrObo2G3SiLEBwoDxufkv6ZH
3uHfVujEksjSgonzLxkt084uClZxaLTDzJn9mbKMLrUUcjMwEezNXZvn0wYDioO6
B8J+Uaws9/RznbVNHO05RpEt4WIWftL+wgwFUnh3EhxNRY3fF8F7Ffg1G87mnFa0
SdEv7Rr4dYnpChEZ2wCogRU5h2sP++ecK6Fyub/bcFbmn5A39LkxMht191jIoGmd
WnWfkLYjd72SxUbmpNHDDPbjmKh5mfDEG/cL1B+vdYlpQ/bHL5uVbHIYLZ6RILon
uc9yErWpER/FbX3Q4eqEClXA203qziJqPyeimT/6yxnsr584Ccy/Sq8Zh5e8JyFV
6FXnivqejQyRA+YEaRSismwK2E9QAIW9eh1kwQrHTC5DnfFNuvRQ29aifPO7n6Yc
Gtl89dnC1AkC7z6gX75aYMFW49HzE+k3PRFF7ijBnU0gCZ4K2PznlnObPZ533kAG
AbABPQK9yo5zzHT3g2Jdxt6U33KAnttrlW0w89ZMjPRcs6ZbGYe6yJJMGqLgx0EI
ng2pdD1v1b5goL99I70WrCP39JlZrWwOzQqCJoZepegtSHPfHkLfHwLORDYorqGW
QtfdYBLLagVocHxk4oWBFr4pSzDYyf3xNyR98tIF43teW3Lva4aj5JtUAWjkemEQ
KuoF1hCLlIkDR7bgKTZD2V77LKZEv1UVfMvp9ktPl25oSaseV9/N2++IL+2eoNQX
WSVp8QqinWFNXmgV/HHykoVST7Zw9Bs03iTqi9KNFmSqtJ8+unzFO6DIkPLTjm+N
LioC60Qj63K7/lycCptMItJMwpv21Zt2z+ogRT1q34GBYvZNZIosUw1jpHmTO6hJ
JbS2pZ5V7IhpvKbctbrw0ilPsiJZ64QrAVIJ4TlMfIDZu/qpjBiscEKbrc29lQbT
CU5Bwp6arVezjBLRF+ljftHgIs4cssiUlkwE+P6djnVP9Ab0rn7mbAEgiF/p16xU
cK2aAZu/BrXn9XTOaKdaO0HM14+2gd5W2/YGB1xG8viMjcmsobxiKa0NkRuasRc3
LFEMGAsPU3u5AdRpJTFtlreaQvghfkPu1OwDLMUERrA3C2+ypTAjh2HSDfO09B0y
hPk+ntdqsFVSbZsU95fYF8nu6GXS7LT9GU+H1EOEb4VxFB86U+vCI39PZyRuZuhU
wG3ZxfV5x4VX5YFHaYwIqXQHspqRcFN+cW2tGriibESJaFvBNTBkLlXCEHNfHvsr
ypfT5VEpBIkMxWjih6FZudLihGkJuGkdiuehOP+PsGx8dp1sMssbrqH8QshrmqPO
OQ+dcHwsiLD3E6vcGbeFHp1ap0bakNeBy6S4EE++ux6CHNmrMR7OOGSHeSPnWKeB
0WcltjNooHperR9TjETpBlVYVKzwUMOJnB+m/loG9ARsEoYCiet8SKwm9iskmM+Z
zBxEk3y6VoK1LcD5TtGr1JlrtFWfPsY6BWqIqrC1fju0fygA7bwVy2RoGIefMVkU
W3MYjZZzNMUhNgyyx1HWv0imlGhxkTUtTRrjN1jNIst6DhsVZRyrA6JMzE7K6Lht
Rnqiaf5aJ18N73fExlBnIp77ZyTQwVslNpSaL5VMs87qPthJKMz8JJt7NX1jj7fi
1TXoElfmK1U7TsLDKzhedm9tej94iSSOMBdiDKBn9TyX8IfcDZ23XkvLzz69aKZh
Yl+H47Pibl+EZSqaYwSajny3iH+CsQviYMQ62WtIO9tjdMDMvlfmDwZB+fiY16GW
ruRm6DUkL9rkZwf8ZNeYXBMBUmsXNp6t5pRDTjyO2SydfIttyyr7EwV1ygsG5v0j
H5rU9h7kLA+JFA5TLdzFf/dH1buQQfTrw9UZ/8ecA8eb52oLBYKlE5H3UHpRGzoX
cHTx0YhylvetSR39EYwHSkMlibCDaZghYCdShhBvxeB2zyD2XP5RzOeKl1cNhv/k
rcLXQNFUVZZ53NH55j9izwBwoR9RRS3AW/WGRFbIbeI6JOHqRLHywh3j908TgP51
aM7FnvEFaSc9RVzKohKAvuTo+SNEGNHBF5THwalmqcB2sxnuyljMVypaYEnI4Uj2
Uym0+r9HYlCAcLDTGvxe2h/LT5Jf7XJc/m7TZgHcA7FImagWT1lGf7eZVIfbxgbV
Dl4sZac9VvWfjcXdg1M49rMX6MgKtUYT10xI6OOC+mevY+fGQKk6+exFH7QGUfVA
hXRYMbTadtK48WQU4/lNYtRd235jb84O6VKaomujuiLIfOOx5q80ypCFEN0lEFrQ
k0qeZfK5G9BqiIx4XndxDZs28q2CI2qJegrxFOveTKuIxI68d5rgpLOf90WgVRnZ
ktEnMmHacT8muv0Z7xwE+ry1Q5m8kqt0NtQfLNu02KqFXRqYQMbmAXkvJ0GY1zT5
2TOHjroUFlMSNF0PG+Prifo6DkLWS99XJVNSGnSgTm7O5hwGehCy67plnhtn/cVY
pkFI4dHjKWlFVRtdCm6EAj5JcwHWrNC8gStFb08g3Y8Y9MTPB6ZokKSd951q35ND
t2Tg6GzBuJfrmpPEed+KZnzDa1XsjUOV+CQ0iJbb6dxjZcguO2U9M0Q7PtkisshI
yNvWfPHtBXRAZJ+KKC+ta5m/ThMoNOMBhEVRySfiS/FMjLTNULkTGA5AF3uyXbHl
Ke1bAz61yZ5IwCIM86UzOGKg7GgBCEGSDoFzWGVKwBg7rQS/XZTqZLyqYq/gTgOd
erD8CDwZ8/wKgwjbBkg3Epwp/cv3H9jjiinzs82HZbdMrDSmiSIs92htj4XXGdJ5
MXFrc79LXnH4Fc9+ylhm5CNhQt0oI1q0sRA/OyGEA9jD2zJ+HwDWrvdDnqqwf5JQ
SjHjLWnJNMSXBJhCuNAkE9Jpn338vgOAG/knuelMSIeWm7+EL9HUtatun5vhNFNO
80BCelu1g7Xp4W9mYtvQKqxt2Cuz0lH4M5vGgVBpDboMaEwGCiJ/GHgondN17wKq
aKkX52ZmT3w0ujiUykxLD4kkEGsGHL9d7O5jATfnLSVZATVHar5iyMGAUtD2cvW4
al98BdUP5unmSmoqcfjzwz3ri18OnnR1TdsScE4vzBTv7NYJBuSn877Z8CyBfmYA
VN/ORqlEnznP7oV/EHFEvLkEEKfehk5YNQKSLsHjebKaf4aUSLAlDEVj4dL/srDL
Q4/wooMwmC9CW9/3RgoFDWwlVwApUtLzS8PGbAxioV61MdDh//GzF5FvV+1Z6V9X
RZ+caLTG/maNcT+hWkh0X2xfvbG9o/4HJVWATtQEMAj4qZiTFBM0LRETiXbFwK3l
ci7ZA3C5xUakmgO+k/68UDecr83rKgGZvFW/A2M111YVbjaewKcMDRRagsuruuWl
4aYp8IWLCxB5FJmAiiAKy59JcGevUsX1YX9dDB9fTwaPIRSSnyHwPgi43vs+HIlq
J9WCXVGynpfwx/05ybraU/A4G0EgfxC8e1vQ+WnYxklPVibJGe9ifmP1C15VwVd9
eThTGmQBzS+iw/pTUbl7adS3wkJUfaK/Hg6QU1DhhGmP2TS4nfHEGIrpG4MEusdK
3pwd8uFvtaoCccZNa6hRZ7Tt2bG9Xwi+Ww9/3eTHNQvgIHT36bDAyky1BvpoCiRJ
To5UpraWqn/57Ls+ECDfypkVKZV0SHoREx0KlyYWKnZHBwQdAi8AEcqAB8+yoQTq
cz6I2KS0x/D93X+VJkZRsT4ELSXh/DKy1Y3oUqrbNfFwr7pJ0oCna+aCF04dbDGr
fQG9BIvsKfVwyx+W1aGnx5VCXdtassy7PnV69Lvwy60um6BIqoV+Hurl7mtJJTGC
Ww7DKXdq7inIjeb1j4QUbSMfgJvf1n1a+JOWNkSm2Gzp+WcJNM7+oggs1Lh0zZmZ
czZYeAleRpmZVaMhwX7cwEn70RufJZ3WRJKNnFc/GBR/o5N6Zu4LlCfh9Aw4vv1n
jBaw8h767HtJGphWAnH1H2nMhPnfrLrlOhXHlKLy6MFWQSgQ3RyhhLQz5XLU1SpD
dHrekT7XUJ8dNxpOnx+6dtDPSVmVFSUq6As4WZGP+Y/6eZSJHgCCna6s9bdBjjmy
ISMT8syRBOSiqp3LcFu8yYqpK1MHrGZxnC65K2d7jqpdtTMSiF/c3p65ir3fbPDr
JdKuEhNTwbjvrafxxI8Q7RAG0cMjYCs3yFS9MHRmk0lgvQX4h/zYCbZezNtIAuAf
dZEC+hz4c8BS6g5+GaQzk6xjdA6SoB43lUXEIs76x5EmHYuPM6zt/TB1OrpRpjK8
TR10vidyl195+KiLSLNHqxRzBpGwTnluLaDyKWWxSqFBcgCtr8NEy7yVHNhbW6a7
8FDCFpGO6DzOmH01KbhuCNm8O5XIYb7gngxUfQJn5tYLNklVB84sS/axgNZZai1V
rK+Ytxj42kcbOwY/LBDCGs6BEdz8vmyZks4S0PppShO9IRxPji4kuNfEjX/8an1e
tutlpT1LaxWAeEci8RQZwzRUuEpKuLpXTSmqfy/pd9ukLSoiVwNKxaMky5vm6zki
oksfIrf11eiOBMNKOx9eCnpmowEHwf3H9kf/5an+755mytgLF9Q3oiicPJju6CMS
4sGF9N73E/eLuauirqF6Ounlz4mu3Qry5e3rhYX9YugKxwVywLujCyw4iP2tD+G+
9zqCunn7cRFP1TNcbvS807/GS/LoOsIRbaJp2QwtDi1XKGN14GJAAm603i98llt1
Aw51oNVlQWCP0n2wSCNY6Xqhfuix4UtxWSQxRDMVJBxPdvvCBXKA/y7LQkGIZa8+
ymF2j4TFKYMk63hS2P1GVmxfg7nLB+THoQAFfvmPns9q1FOqgvkAOH0dOrO/2Fxh
6vf3b8Lje1uMdYURRJienR5hj1BJeJg3GSKiAfLNkB+yRYPXnBO01yvThPS+AozJ
G3ohfaAJ1eY/uOPgye3Jq+FPp9QSKON3p5X3DAbCYmqbEGEw5GAMo2YK9A2mMhWm
rqj2/5Fd5ty5pkLzrhCCi3b5R9dT4hoH7Ugln4IzPpwNB3JnLNTg/WnAspBnntTj
9V0pAKJWXPrBP1JtKHnb+bmUrttwBmWzT3xqR6M2a7eMNYlL9TNwqFoHZGT4yELH
1cyN0M9SuKOgR9jHFppTjkdyHXe73Gbyj+0r3X+/CJyGcs2LiOeV+9iv7t2ip4ms
a5zA5cgRn7AcD6FGNyo4yuRjOHj1uf2ESLLAHmumRMKF9MG6RRVWv390e3v7ucs9
W68Wu6D3qUcLlJ+LKLZdKUskJ55nszWPtWQq5PXt/pRyBdCcPCMayaW0b3I1hEII
EXiN4h2+4Pge1dPCrmFgdfY9Z77JVyboSKPl2OkdiIywR+vMCBRxYe+Z6Mf9AehK
qaddr2ztHySiNrS3XOFqKbaXgKZ8GNfS7Y6fV1UqXNf2DuRVS0ZVwDumtCPOeSNg
+pT8iBja0HqiCxq1vmfZsEQh+DfGNCryHnR7Ha2swg5uarVY83bzJalBpzyxCBC9
r4qqnfU5i+E4h3vThDb6GPaCIduZXhj/W+I7VY/Rj5BYufw6Vr2HyDzKLGeR/iAe
TARsuN2aj5aMz++L5ye1dihqKxVvQbXj5SJ2ViKPTexnIWbdHg4A/n+Cvx1HyS88
if865V6R1DzgkbOcwZsSC45wwqhBLhw+XIJr1n11HN6WlCyVAz+BTESD+byR8Tg2
kumKhDNF1tvTIm1Eywl6SvQvVi7faeh7L09y65+SMw02rns0BlNev3NX604YjHIa
gjdfJj6dvGpdtKHsVROCxZj2B1VjHq7VjspGb+LAHxrkJnlbdYVDZeEF8S6Cs/ft
WO1WpeXP/IES/ZpKvfJqWHeDDe1Rz9Xlvc1RqkZY5BmWiVxst056q/XzGlmTWwnX
qMK/GhDGMM0+ASdZZAIsnLSvvE5Inh/W1l0p/2yx16PxWVyoIX2WCeY/MfQB95iO
+eo+QWQdoiRBiS9DeVFbAdvYU6irebUBt5DFm4pF4RfyPiHVVBcF1IMQ7E9nifvl
MSrSFqnU1eQY7mmCbjXxljbbwBzC09fOqW1AMYtni7YTD6U2+Jx7Y/jWRukVrqHi
6T8mP1Gmi5iJqAsDAQvkxgqUcBcZFwC99Dk4VNxSUr0NNq23P88vNKlwl0guIeTQ
nsH5PJMjhIKoQzN6k6daCAFEzL8tSQ0U6qG62kQUQgXH6g2w2NgDppGPrsOvNKRL
uDE9+MfylwlagxuhMOUQdwafleAg3IWTA+JpZS96V+C053AdGZclKirp/dI34HoM
9ZU+p/OBoIQn8kTqqAMdB1pcUTuWIBSgYZgjxzVehgK6oJN5bGTv6JBgEP8C+Rro
uu19NDqlaxK+91zu4LgUOdEvd4GUmQwsVWeRaf6SXnHnfPVpLcyVZFtnTZihVQqw
IB3hIy1fasIh3MYzUMzy5yafqXHWAHsV2Z5GaKNQZCPfgzcCstRT2RTqzJdAvY1u
XfddbeiV9NhNVRAys7jC0l68LADrBkLkH6gAkXkw1kgatzW6gwtcbYdm3DoRHKv4
Bhs3tB1aPZrpuE+nfQ9O2KXG04zQlU2u77Gto3PLfgZo2H2JY0StVJIzNhzveA1t
Bpe5QvS3jlcSzPKS1GHoszJOr2zExo8NR6jDW8zlxdi1r/NE3JOlHwN4/1/6sUKg
2jLH+AyurIKoTD0Wu/D4LvODvxkArkhAkBasZADLUAmNsj51FIXvuNdczQEABSYy
X6DXs5ZI0pbEpwVExVPMkG0O9zH9yk4w7wprqHOWEmTR2V8Pz4tEMG2pxKJcWpQI
3Ewp4UGCvx5Fi9Sd8IxtMLyjamdqZdh07t+aJ3EINiMzXl/fxoP1HeARfpjzAKZx
ZTpVwkzMESSIiZ5QHtLnXha+/KfgZxtEWayt6pRF9vfrJWTPTROGKRkzWO7a8Q+r
Q3eGQvrXL3whvLyerbI4CvO90GfoNc0ewW2lbPKmgvAe9/fqNdai246k/MfSvogK
7GssQl96WO4yvphbYeEW4O/qQ87nWhzhc3ppl43m26A8sQNuOjuXjduYFm88Jl4P
ZtcvgQj8DRWfPxEMB4TjCL4zllvIcvRp7u95ptByyN1qHTl5F2BhYAfWkIgLHNg9
qi3ja78sz/yFd9VNEyyqhuwBGRkkbkDppb9w2QjoaANfhVj82qw/C1yKAd6rp4zs
GAiVFEHVSu9KuC1gakmSdcOTy8sIaIwS+/VcNs7pJ4MV0VWx8q/39cce7eyjZC2P
4iAVv7MKKPIuVATl56OQxsK8ppJ3p+LL0ZfaLraAchcMnvoO+dbRh08/p01Rmbqv
+IgrlZJYt1p1+I5HBZo8reSOQM3Nxs4xBG4HUj5pyvhz8DzHp4YSsoALibajIrGz
R0nn3fvEgZsVMIzKStC43mmY0iKlLScTv3s5rZzP8eNZeS+SMRlLbZXOmdhrxuWo
PfIgQyvc1ExoIpv/5Ag1Pnr72gzwS+wnEsKNPwuZoXogH+aI9HGbWElSgESLgJhh
NYuSXIq0FSm5c54sbz1sAc5X088BhvBkqL2fjM4foVuHjXEBKIJmnmBZtguGE05P
saBkzjiMc5admtrcKNemvh+9VSPBppSjT1Admh3+e4kC8SjTl9Q5uvVOuycrko1V
5eD+8SqQZQVjp9pgV6vj5mFl2mKuDRpsVShtYuRIa/GIsa4MGbFP2ybuRB4ZF+D+
C51Qo7u/DkAoWNm5gNVZq51xeJl02dbpGRpyE1p18wZgPTkv8InFsFoyG3xLlLrK
sgVXn6bR6lKT57sw63V6aX54pt809asZNBUhjBACTLajR8QJGhmxiQR1+6p4oTYX
242kPxZpzHiVOfNC/it6Hcra/msOnxI8r8BhE9Rio7nYCHo8DUflD5vCQXhz+UPc
oke8lC/pbdX7LCml6vntgD8TvEV1nzh9zW4uLGtK5dKFvTE4hwBFkqSEpZwhyDnV
W2PjEPMZ4tC6HuugrJVLRBD1fQL1a35wxAW0ZV5fpJMP+8FwOCkDnb1FYA3aPcDs
ql8ZOL8Ck//s8LnqmAb52u/GvgGdW8b/qPn8wUaCnioaDOgLqzdu0ewDSL/4PTm7
ePANoGH33ZR07wKA6N1jltKrNS9X75HuaxIuuqsiGr/zI/Yv7arHyUb48FXVF13J
Yk6FRjrWfBlYH1F2+N980DjSAmIyiJsBpOypjrYlEGAUZiF8KSQ0FAkqRaOQbjML
oIwGy74BioUWIL4UbEGJWeFN27xf5z7qMxYUvlLlvnEwlJE0i9ESpbCuqLfKnXc8
DiizpTM4tvJwDNLJOOqpUtNngRVrVTwQIrVfmZUuxbmCQd+NfIRcEu5NVJBqFynn
bYuveBfNeTdk9eJuUtUM1DI47Rjr4fVooX3X9RKT03ieaoBVyN2ieUScSPoeL59F
W2IubWEnTNvj+gFrR8ezwbGeU1mdtrMDkZObyiucUNa8qlyZhd1bRNTVYnpxzYt+
F+T4YDbOESpgssnutj7mrp4y9FBOcUc7CP7jhnA7wpQLyTegiqw7ElqVfolR+Ag/
gZI2FdMkfHMex6FM9nSPdZwbNMcrARgoqMXl7QpZp9oQqiwQv9+OWzqU0xtLtMBN
REsNJCnLkwnrsnb3lV/2/4vZ2rH+Xq7w6DqASTI2M+1NL981BV9xT55E60elWuf1
4+IiGJgg2JVHt5BLHAbdjeoY852ske8hbaLn+LFFvzdDCGH1YqAymGM3+M7CZdOK
5i8/DYFrkMcDgDQ11jekkok/K3EsJg0E+UTEH/KxhSakQxoxLAdok8Fvx+jHzv9U
si9sVnndEPpRcg6zX09hFRbNuCsgWp4IvqQT8Qv/0poswV40LJGbBL9VOjGR/vrG
x4ZX8K+FJ/HkHNeUoE73bzs+VDaU6/Z8LCAzmHqlbtgTeUF/b6tLFYTg6vpjcx7Y
J9/g7CgnjHP4dhGwOEeDFtT1Gujqsxh2VCEd1QeMCEUBylJBpgCZIxK5PuD4dosj
arilECXljIKZqsKIYSMBdVSlGwLcj0uTRm2pWzyMK9y0KoDFaxZgFE7+HEeCCaE/
l9UYQwg+qDDj9Ul/PyrihbDPDPKXxu0kdKUeAGP2v0M+8CqJSb40itjTVXpI3yQk
7LflEFl6Gf8o8gOTpGRy8yk6LE1AUBeBonZpaR6FdqNNaobGPJtYRjtCKQ5TORBk
xueJTygGqJza6O9NHgYh0EXv0h8pj2Amm5K/1yxGKjnPRhwdj+cGLeqrhNU/rvIr
RED39rcGrN3/BKdWcoc56gYpyG2jfkSxU5O5OdC7WPgHkCnDnFlCMS4ao2E33gWp
llKEGBBYtOeuY+04pw7K11SAgC6i95WC58kEl08K5XdXgBfRt6mxeULCsQCmqoqF
B1nh+l7EcSxs3nEYdQUHIizSGm9Fm4TujUvGlv2QknVLiFwb1kNxJ8x4GbvCKkHz
Wm2mBiRci+q5iJcpdPKWy+1HdzRvxGsccpQhh3dcPZA5QSAtemKalnSgcbZDjXqJ
0ACHLPm69UIITajP6jYZksJKnTS4cM9SAelomjWkhAPAekC+s5AJhGbZ/g05TXmI
b+hlsoww9pNyNEYQLFVgEx8mzE7Vn7M8eNOzOOClNoTMjpcEMxhCIuv+PUsqHl0q
dY38HeS2mdTZEmIzbS2xU/bSi5SoNGjz2wSqxX6pS/cR3Ba+y5ff0S5l/4RGqZCB
DvbBh+O3dkb3lOTJklfVLm9UzkcsJOu/aMqTAhY/c2ejm0ZM77YwJMLJ43R5Pt/i
S+uS6kLz47YUrvGljb2kGB2E0/9OCGSHZYxdNpLzffU9c92mMGigpF4B1rfG1jm3
bD+UDNKqxTDIGGeFuDfJe9M1QExpgaXEjNgXInSPlv5qXy/FaK5oIk7aIGrWGSar
5tInE0zCsTJPam6zOIiUutfO4tyMiDOwKovAvQb/v6N+1r095iHNrKcS8+NdTUfx
QkXyhkMplM9kMBVZ0gpcvKgc9aptR7vps61ptId+PMR3RQ4s5J+19PnU+MAwlKjY
/zDgyzg32D6RvHVb0KtR1tvR0rgXoj4PT+Jid+a71x8hK05hrHzE+Af/nJlqH6Uf
clPwqbrthoIzzn75adxOtiNTJ70Uqa90/wnOvFv0KsB8XnlkjaVX0XJOH4ap9MJy
ojiv9FSrafLkMbxJN+blzpvWKyzEPMwYrBwkAcHe3v9+KGlcwQVyIuyTyHsMOkSB
6ijs5JbFRSX3O/MuxUC8MYLI0h0CwKDT59KJoVmMmuQgSyu5noMEzPWJdYQhMMHm
pfEWc6M3yIA3xvMHLIjz0LkrbK9hD2zEeD5No3zPxCxy7GJE36S4RU0L+k7wWr0B
WhPIqdwBRMFwiGS3eSNIORpYfGOsd8z166F/VWSEzMjpjcc6mFBsvZWqN5OcN00d
0348EgwYeYgiock0RIUvpSGgvKMW0lecsI+MvVdsRdzL2i2Z8rCWpJTakGsihaTo
BVYexI+1kKTt0Vg1M/hPFngnvukTK28njW8TAyyqpHtxqmUaOjDfyj/i2aRpLZZt
6gAqv3DBn7VfzeJU3BuJnnyh6pbZVx3XLtfKQEOEbj9f0nkMrwX0h62H3IT+KJeo
QU1cPYyJkiewCxfkeBty9HTbVhK3q6ZtTxWrFHvOssigS4BdsZbhETxADP9MX66H
OqTldir2exlGLoD/WRAyNV0su0UJbw8ZrsyDcVED9vRxvQbi2g2lCvu+hVt3XP8j
edm3c+Y4Qh8oRE9F7iD4EZT9/yPzZUmrXF5cE7bGqNrru7o2k2SeIeSjFxl7VuUF
wAFV1LKO9PghYhPZpodTGLoNoC1qVN1bXL9scVVCWqebv9WBzxcDbuuunhxgbf92
F4lNh4vrD69kp3NU1zdoX1CJB5eYv7gpnLwxXR9EPBSz3LArhlLr1rrw21B0xZn4
dg/72svlDIikvV0WuFr2k4BgTykrYh6dcq6Tk0HB/Uxh6W81iGw/CseE+soD5HKD
mmB8EhkhuBMKFmBF41YKDV9v2AlpZDzdgYm1svM8Bxr1ZBYglQSPagP+PNUvNIcl
uA2jCY3AFDZLkSKawpunGc5mP1tIemG78u0A9gKpEUgIy/+vq/tRlnRd8ppDFl0V
rRd5ctNSPNdBwq8i3fF07hg/RI0cdoHgzTxboxNHIsNh9fLjG8OVt5Mm133dy8d4
aXNJgKbkpUGE9R3g+UhObv6mY5ug7KDkllUfcuq3c1MmHJRbQXTzs8/Pn06fZVJg
c/A+zLmP95U/sskThDS5G+C45w8G1PRXWna0e1EOfgxssGmu11myao2bKPRzPWe1
/FcE5VQYBJLj0lYB1ogA+pPkQAJ6O0rNigxvFVyeHWovgHtT6qbvHK1W7oZdOxIH
dpgal04mN2n5iQAO93sje5YCqNPjUMYWTGp4eUwkvYg7Z+VsEDsie9Ma02aYi/iF
mUkEgEC80+pKWJccr1n7EHN10JdwQpJQB7LWgma/UOSQPsLifJNG3waHj7Qlhh/M
a5zJe/q3yOj5FPK4fK75JzACNikk6KCBsmJNmWEslUX+/1YELG2Q0WbGZ4Z+IZvQ
xNE0xFQQGqvoky0i2Hm5DWuGo/m1aZg0New6y/JHj8wSoeDJE6P8CbZiiUlj8Lhs
RQonAt7729LQoxVW814wbb67nVUPimoSHvJYQQgy/B1woQ/o+3f9HAhGbKvKUijI
Bq+MfRm2hAFbvDhYV+Hksl6yQVXQTxUN1GTSqjpxAOCoNYdzOsmylARRxpTbXVTD
UJMmqu7UZl6dYteoh5mP/xQlWFe/5CeDoTylyDUEU3ApCjLSAjWKqyUSs3ONPQRz
Og8QlKhZscwrZJaeLrwsGeOMqc9qA++tl6A8d1GhmPWaJKZMOtieV4DCbqbcwx7c
zgiiMacJ4FDnM2h/z4oeUf1e86u/0DQwCvbe73CXUe/jRm3Oz1rnRbb3Wv+fGNwg
b9Mc0+bB5nl4Jdf73o3vb6cjlhPF0kFURkpu2Dp5MiLnSORABAeUQkTGfttXIltY
C50G0zUsz0WHqblaqADo0Xcc558GHGSNdZHnKxO+d0ok3mb7Em8dBYmBy85+bzPY
gvXWyywQCiOoXGY4fe+fpqqCHRJdxa5LljWvHjP+8pVf6wTHjxh7TRMoowzE4cWz
9efG4gxhVf2Q1LNiIQQXN0Unr3nMUj4QbGRvGO58Nvu38TSYZcHHAn43kro0GUWS
tlkor9dkxkMeZ0+8fBP0jWukGRAEuJ+jiB9UBfuixCv/qmHnCMxmSzcHnzEWq5GG
OAlV11hzAEn3Z4ISAX93JuOyUlTY4dCgXR6FKCjTyGhJSey1b0lgYeRVDrLVyQaM
oYVC/Y43Ikozpp7R5sZXjh9WQaTCvuS1huPrndvdNFmfoNp3HGwgvF275a7WNZir
pTbxBnocqnzrEd9tG7L07fCQIfcMD0IEcEpV9veheO8MC4DyR6A+sW/Bw5UN4/g8
1Q8fSco5dgBRu6y70fnJiutL/bvK85kC6acd1n+WuLiO7sxehnS7ws8vb/pGaL9A
SQisnIrd0sNwlmj+Kjiyz3Heo4wpQU121Q1OG+BsvpxswmSZz5TVbWYSVBNkIJ1b
5u8rH27jD4Gp3qzeM0IgqYDAAILPflctKEvofdv53hSOXp+2k0Q9G+/Hqo5yU+hl
T0kwHwtAImSzYqxpK7oUuceSoTqL3MQDGJNDbsk00yXdAM+ypPL49XQDmvAdR43z
QVBLWDA4yP3boo8ni/oaemUYtuq1KeC3nGSnya4vYKj7Y8QwonxR7yZ+nDlNb2Jh
PdUmLlJ4ZuP9m3VYh/735db3tvMMrNnqU5QC06301JhNPubT3IyowiBy2EDGenSQ
Fyv7uEWyLVir/Q39BI+uG1ZXE3AzuZxs9kA/p5Resn2Q2sMwT971w38nrtwr0n4H
fODaGCcG9GqlCfYEP6n00vIuCas6fcq8sSjuDIK61PQTHIIgmYt6NVALQcEWgeUX
RA9zHGaQegtuCJHSyJ76Z5KspQQODoZsd31fgn8suUBlMl+7yjAUss7J7b/ZfPBd
HG73z+fYYl0hNk6d9jma23v2GJSwYFuT1BRaQ113Kp/Z57A4lDEc/n4bbO2sdKUG
HWFxsb4Hkq3A/DS9ZGjLUciT12NGfVvGBtFxFqxIi3WrgMUNJc8Gl02eGBgoQwVe
RkT/+p4SsXuExE6vsdtsOCBLC6+AapE9Llre6lnbNnh05I5eYpDV8/FSGlXReCVt
Ytiv9sI7JDjBsewSyYqVRv/EhO17IrCXhagl+FbsbxBAreX1cqqY8VOlU2huM5Z7
f1FO3f0CuQ4Y8XjQ8MuIi4VwZ+s37pERKjh3uec53r115JZ+uiiPiRW6POZkDb++
weqI89QFv+77VoSl7XdnT5HulI158ufB6lY52P6vc6dnUPSI3oT2KC9mkFOxsF2i
VK6gBF376wIOFOyEwmqbmL7CNnAeBW0lPX9GsQ1HXwr6kbkqNuO8OCh/Z1zOQjcP
FhSA0og3/0iK2n3vpkBi65HD0MP82Cpxkd2O8mcoQOVk+wzsYZMrXr0Fmevhpc+l
S5C+EiMg47xk8kgs+SsD70OZY+ZFzAfkK576dikPo/1J2+8TmEwWv/MFK2J0vW9W
ETMR981BUbxrgmPu9xjoPn3vhueVkhtGXIIz/hvjIj0ALck8B4h+Mwms3VKZQ8Rq
GjsC8Waf1nWiWdpYgch+CDtQNBT3oPpQdIkWY65xRMdtfUZJRsiiMqINzw52DbXC
asCxCfci9nFYP92a9GuiM3m0GSTsCV9o1CkNGg6SZa9gpZaN1tmHsDiLOYB3XbUF
Oz121i6fNkF9urCe8e/bLpOHt6ET+IxId3Tz5MtgWUhne97LfduTK8jS1d2TFnDP
Mds5a6cL1T0N78nItZ1LBeaXfxlmJyKKDTCtRXx8kK1FFekenxbbskb9iMmRKKpd
qpxFgB9ho9u2Vu/Z5lNa7fwlqqc8ByCL4YXvdTx3Nck=
`pragma protect end_protected
