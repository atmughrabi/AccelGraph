// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YqMCVXrmt4tqKH0JAT18DcTDw/GXbjrpVQlGmpb6GwzIfw2QLGW9bY9zFH5LYCEl
7gYTgGbnexm29vuBmU4OKWtHNx2AWAFC2NK2oms2oa8WO7YfMEUo+Txx+BwbRG29
a1eOr+2dMEeU8K+aIxRjw4DDhYqCNwbf7Bc6oe7eyBM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34480)
oYX+7Wh92FPOFKUqredXsJzC8em6UWpmAvIbbSzhidyPLNzjiMMphEc8p2z0JBJJ
zPkdICcL9RzRSyz7vrKo1hWxjRlabFB2nfINHGbKbZikSXxhghleN2ObhgwQWIgv
UYWV33SPgE+uXYTWi/kRT0di+Mum8RWFw8EYMFsO5+6SBq+kX1mNHioBexhNvAx7
oiMXcmvXcXiBg93PsCuLZSvxl7isI4nLWydIKkmCASSJw7wH8la5svDBzLEfrAJ0
liNaKusyA5JMp+PeJg2nxMYBEJeCAeB+0gHANIhatHWK7B+9UZPO+BWPEjQq/QAC
gRjYCokFQGlV6nC7aCTNq5WDn2+gnqqtNACGSA2M8rrie9nrvg/A8ulrWaVLM0pL
DG6AJ70OcNJ+JlajKfU/K2rJWW9lvJyTtD47+IID4ZgDLTdifTKKqnIjEoPiPggb
ZSMdPtmknAZ7ewZHg9GzLtgFfcBT+Cmyw8rv6q5ReX0eR0Aa5S5ziQZCeCuxc+SN
rUEUFzufP6Q/4wJwtFJ8kMW99tFrlEPFF7AnwIGWL+pqvBp5+vpQLwx7UcMhRmXN
Ljy0CVOCoaBkfQxrUJhd6vJ7HhiP5wNAp0L3bxaYy7cWcsJOm6GBhSP/sUhhxP2z
ru6zydZ/imTcvr0Pstz1dovTNd7dDTrerwqhCvGM+7UL6mPXAnW7sTHQfu4drw4m
my0GKTI10pfYljwE7J/DIEoULETHOBF1WYA6wQf19oyQzjYYpUetkH7bmMMNZmLo
QaerlqPqrYE/Kq2bBigbP6yUt2HYD2DwMEIoBsXT/aMyyixY4Rn38iAL615CnB91
jnY1LSFmDwJTDSwBXLpMYWRgV4iaEptcaUIMHwO7k2YpfBdwwN05ODlyC45KkO4c
6CwATgWKKxR2W4/N6sywbF5DZxDNVuEaP7If2xjayXduFM7KbMhgkbHRq9uybxik
bjkPQvk9jL+eLP5bPHKN/AVZyLybhoKEwvX3lVKduch/hgV9FcPUdI8T7VaIIxi0
BdjzK4pYuYIlwyXmf6ZMfjYPvbkOmNwi/8TqlbIbbbYeWHEEM+VEZZpPT0GhCn79
+Ky7I/Qs0/SJafvdw7Z00j3WnDIigiQ81JeoCRlfBm/rF2x8u2yD9HV3WMjgxs8R
E5GO5tnO5dBreJ1dJb/cKc7HspMoQXV19vJkyD9DlpV0jxwvI58xsiOp9NhSXAEL
3VsCVWA0CR5QudG3rdcO55oqfE0nUHAxw0/w4gNHI5h92QXePVlVR9tG574w21tm
oO7yLGSz9/QHO0y/4XyGB/a7Sns8nJFTi1tLORiojSmnXLu+fbs76w5uYYiQ4Bi+
jqfHjkRPLe8O+c2JU55CfxHbxplZEhb0nBHF17CmG+dGay9PVtF9UAaLUXA+nhmi
fe+1mufDxDKcrkVuN+yd02oXMM6hu8FmE2tMLwWnfnZDgOONYormJYTI9JEbcn7/
nnMXlYPpxJ5XmlBD8C5oBdSwRfM4e79jvUUtGp6p/uNYJzuaTNUFuKIAMU0oWYGp
ibmCizCCq53nAO3NYK6x1RCG5gobYkvzIMmMAwfvExfZq4yNvrYxD+P5LX0WfGyF
hhlTo3k497Rt9vuHA/1lggypDOHTS/KexbRjPWwosqqp6dwi6WccFCd9GRHiKGHs
Rx0QvJdjgwJFFN3zeZ2T4rCF9sBjRKq9VsZ2zI9+AY2SZpzLpF8BrFD8J2iI1i2/
45jtA8m7MMgS5vHwWU8B6/bP2It9BRJU7+SRgo3rmTQFD3MPC1NZOHWyiNnqJaBF
YDMUZY+cVlORkohoFM5t14skTlQFGpcYwJMUot8VxaVa2trOfWn1NkGhw7oFjs7q
D7WRxwTCEQqGCIrHPoPsydRY+NkV9+o2OIXs1S/s/iIQzA0kMpbFp02Is42MxnSR
bKR47P+/4lLLvT3ZnaxfOqgPSal5vbWgkQw1iGGp8lYqkzwdyiONYoVu6IvNnk8X
t7oJ9+nghoH8uA01vFGF9kkcMbSx3RUF0B2lW588wTVY8RJurjunD64DAAUHUFlH
3JSLTZG/E9OStTtMkxN0OCPSmgnmLVtBlo9rMEQDp4jeQUEMHMb3/v44y/qChHeC
JsEGl6dej9ZRgkAMmgBfNb7qRr3tjFUTSEDAPqg6cQmQFw2JoamteRI5FXIFDPTT
2hUW1eVe9tKxpWI0PjBO60LATu0QtiP9VkoHp9OJuXVOIlJFT4HTkTmdWo8HwDKd
VMaSqYCl6vz6TGJgF+iXQzJWxWG/vbbA2yalLB6+8NyOJSoddLyK+e4u7gKcZ1XG
urEk7FITaBvqLOB1El6I9oKE89ZMiJn0HLrTqovzGG9ymUkm/UsoGDZzTw1FLI8h
MEcoOWGTWVmGwyFSGvALxZo/VAJfQptIXoT3AGVUeboXSdGckctOiW2b6k47I6f5
OaakxpKqnd4wE21LbPbB0JvPui6Ox0Ze7G0yfrVXrotqlE6sAZMM9U9frck0qdqi
xJgYpXdxDAgpqBRTEAPX2gc0ctmf6XhyS7yRaMeAAJ51eNMlhf21KwA+XS64C08X
tKZTW/q99FbvyORIuRS2KysUgK7IAiQ9FsEC7snRp1QePBLfCV2osmH2qdFtbTa8
Ww+Ya+unsrSDMZDN+ufdxGpJQE0nRJ6DhiZOvAs0M39v9cZA2M3GLFrXTIYMrk9L
akdQCqd2q2Q2zgldA9ugjwl4rF54GOMDWLI+9Jp8QwYgWJTdCI28ytJAa2mvLeSs
Ky7/Dmm3XH66JPEoAYj30BPWDWHOyhAtCP3R7S3JxFvvi2E0hKrYoxXGIrPHPr6C
H9msfwb6ADaZcq1Ajmks6OzGa+KiTzFDeBIi/c1GmCP5czEJi3L8JdJ/DxKCM00z
FYUSOuKnp30Osm0iaI3RAvD/09yMrgP2/xwTdYWq69evkRAk4bMhKIx6nqbeKFuL
MNptYhKs+Je4d0XomHbfGS0eQcFZUBhXVEpg4PaTzhSB/9U5m7gmS1JjCkkJqx6r
q8iSvU8AGdellMSLKe+thBRsqe+M/2tm2iBsMfM+UGjJtT7vE0x/WhXHHD92649m
/jXP/C4RpC6Z/DHnXAfO30bHRRx/SO49VT8JrsnONc7SClKGUPXmb10YS3fnyOLZ
uaVzFhRe3ASuHJ/aWsK7HJEacYlGaI5CTgBL4A/1Gr7wAmUbe5Tf4j3SATv++v7c
FhYX5/2cpbg0qo7bYZXEUSFElMxSzRHKED21mSnu2cqFJ80gRlFNElFP8q9dcvKW
Yos+KqnQ/y8ZWWG1S0ZAx8PKJcCllSAcQAQn83tDpCEFiFecRR875raZdXTTG1yS
8r6BH6K8isdF0iodr21z3GOadGpR1UM4JZHg4qlQVgZEOreGSIWuEvBnr5x40Ou0
nGHJCmGgMHLMFA//ZipRese4NHkNSXTl6pi7daVXfPIFqlF1N0CjJj1NRVkOsp+P
hl/lbDhlPAk/CEtrrzvuhKTWtgcbruVz4zNmFGW4sgpF7LfNg2CpD2/2lw1mr5fD
mO2t0fi/PPT2DqphnqY+2HZrlenyLT4Y1HxB1dYeXF4cAHlzFk/jNc3gSN4gOTeE
p9R4njy3eUulYjYLBftWcKwes/9L2JpjNJlhToL/DcLG/5xAm9d043lt1Fgyt6eA
/rnEzZyU6FRxqZUIzwUX6HAK6Wn8QZD8aRrc5bcrxyDDV78VtFOWV043NoZoux9l
fwAeMESbkceM+FTpEv3lvIzSUjt4t2UnOW+YfOAvpWeo4AsWZjTK9kuYAM4dDqHL
r40djCoau5pVwApEeXMpXm05P0mqqkUgj5JjNamNb6kgEBJDXH6aAzuylDi+XJ6t
74/go5MTatQIkQIFWAisoHKuCaERkYNB1dSexoqKGQLM2I0m3LYro6u90uf6pzbe
x1od2zrLjrTaW55cBF25oeIHnODxmWoEoXWtFNzDpAGpzGcZPL7dJmoKpIFk4n/v
MfLkFyL72094tOsi7K30JratEuaMmLeCDCd2JU7JTWh5J9HrdhCmbQ1Reh1vxAVN
X45wLQlFt/FU1OAXmlLdmXMwrIytqM6fXmGjhepN/7mZZ3EDkMPM10CRRT3HrG6k
LoyvONT+5ii7ynE6/l5XpdUXyp16TjkcUNaG8txRA5sHKJmdfRJ8+N3IMRlI7JMy
asZpoarzz2nMNrF+w3C2ZhKVtE4GVKJvlHLsqbln7qPsLynzWFnG1F7ig4C3CDXz
dEg3b5gOYVatw/D1cV5E5HRyOChitYws66+lqD3zqlg1r9YQmrWmT5BWvWbGfOC8
uvLQPodkFx6DkxR02heW68gWiwgid6/lO7xdQ+1owlhmfSp/sSAW4oLwGXr1xLMj
0SN/sMQGIdpMmUDeGrk1XcsQojsPC9mPaSjs6uxY5Ig3qv5XXF6B4FUfEsjxIP4u
CE8PH0uSIPAtZdmG6aupdZwXFGpos52Pd1CXNU429qRSLJ65L8pkSmtevik1UGot
roo+UcNEkpospyqklLLu8CGHuYFz8Yc2cVKc1a0EFeXpfPExBWRN5OTuB9XjezYX
ql0EXc1bzPZf96xNPctfOvOwV8dOCQ4NTG7Vt4S1+gNbho1gjrM4gzCyHdi3hYTS
fsCfqA8noMa0FZyeNWD09/xidMAAqwDpd1nEwv1IIAK23hFd7O18TF2l+20wKW8Q
BqXfU+jGb3VQMHdfhl/M0qVhY9I0xiGID7yWcaGypvXaxOP4ZKK6iEAO048UD3M2
ulVJOgR90hrX11g//M3r3+dVVom/SXg/d10wLUd7BbvGzrOKlItIHPLsSmhlsTAb
t2UT6z2JjGSB9wVY1n8My5yZSMN25f/yAri3htaTT5oj752nOo60MD3Fr80eWqWn
Nf5fxS8dVJ0/yth4gXEqH3iWk1ZonSq3GfzXbd32w5SU8YMJLvR44j7NClhv+Y4z
1GCC4gJPuF90WAZE8QvGM9a6FhFFGr3cH+Xjp7mXGhNihlhtslIAJO7T2qv9QGMC
uArpghhuiTaKIlBBgUrO5wAnM4ISk0u/9l0jS0vxDTfDkRTLq0eSm2HSJdsrKnuW
HKew3FMRKrn7VzK05jFBC9QpzOvl8km4pKSzDoedppf4AAG0rp2HfOd+V6EDq7wI
UcjOzy6VhTLimQ3QZuejPFWLZeDmqVEhEAKbkTcIp4DbfuX0SpaMgQ6V48/+9GMe
4ZUXohpKIMtMGqu//NHiawUGorGZfYJ3IM44KMwgKWqZhGVXNJK6hGCZKxzl2+oN
C6Ol0IMLtnGRXUAzmAEPeB1GfD/DEilhIOYppDJTFXO52YNhfsWJ9qpTUwslUV1L
QdrPOax7oQNih9WfSQ+SIM9TXcYQYNzWAqkkw/F8AeUp3PRHWH7nWLCVfBmkTtll
nQBbjd/FA6THquMffseGTVO84s4fsPGwiIPNkTiraa8bXeVtwBi+IanE7ao/lI8w
BGdpkil7/aGhQR+Ougc3i3nvlNyzSQVWXxcoHF+nUuCYVVbtq2uhO0rhUkvXSrre
zIf+Hdk0eP3mxWc39lPeOb3I9vh+RXV1EUqw28D3olWoVN3CbDVBUTjyvTGBR77j
0+b5/SoCdYajFyTfFFzLzposl1E9SP5mjvLRfQAdSZqHvrbDida7cGmb8m07r4Bf
wl2ZhJO019QspaJhfZVQqHa13Wse70oaf/WG+csbGouhiybxNe/UbWyvaHzzqxO6
yuvYl/+9OrduiY43UE/dJd4Iio1sa+g3hikcUJ+//EeFFvkXYdHS8ds4GoPppDzD
3okKMZwrXmqaHlK8VD4n86hORZb+jFfcHiCk3xydt3aQZP6pHwo4HoG4wYoGe1JN
+OY8gn6Snyo4uC/syfvdt8LI/NBEhO/LJ5XzWNijNWLiglmGLQiK2ndOTiYTIJNY
ufyez3ChcbdwUYRJAG4VQS/s0Qy80Q2X/Jb7bgjh/rVHjfH5Fe8FrjVWRoYDBjxG
xPLGSPBL2gjM9rY7MGnLmbbxhKl7KB+SrmW/GMd4haSvhDMebs8b8NZ1/+e2ppc6
Jfl/V/ujyog5lI+M6ci2espxuI2qV1MdPx3cCLYTNr8u9xKvxlJQpK7OipKWMOoC
GClMwBz+KA+wToeiccMrp1O1FtXTDq7yxRDIBeuj8BzuyyEFjbx/HNi9Kdcbljws
Akek53CXaMiyuN98Kb22NKwxT1uvPW4C1iN3Nt5hWwzmD5tqrij11EFjfXf5s1/Y
7Wv+cA5aHAI3VhnWE0C1rHBpOgssDFPFaR6/h6f4zex6MNco/tXSzW7h49wTYtPj
+E63b/ABCtCpbWxCnhdx+f7XZQ5v9Ce/842rttV0DnlLcVdVcSwwY3kDLUhxAXgr
D6RDkXpoTxQllflLOQEG8v3lMK6OZey96MlyWHHmfg5lCGbqcXEZUpYvokdEGlbV
7MW5MoP520n6lm7/mvTHwQQ1BIgOYTXMs0VuTWqvYmM/a2IP7kqMHV5a9cG3Xbqn
DMKzig0ykbHBDjL9a+q8dzOIDytMq32aaVFIZ9C4zOQi0zKjSP6g5ewxp6fCX5b+
KpVqUsNWOWrT7XQoXOrOrAZx4qrMpUtN47Kudh4ktpVU6W0kpIEkcoBSiWG6C3vT
wfiVh3LlxdqyuCUTH69/sg1ZoKK49hjHmqOrkBpob8FrXzZ7FwQ3ei7X6CzHv1Tu
LhG06sUGOh2IZmlrkrJ+Gt/cZYRrWhxJM1t9+ozUoS8Ajp0eDO/D/SXnWXD+953B
n9rNOEs8ROcveXe4DLoIPb49MWfA/GDItrx8/6vIzhZcEvnDoPJ+ht9dsPHm+r+Y
FVWdMOVqkyu1GsEKLLuBC+xy/aNcAJbsqzcGxwNgNPXpPKnOKJjZoToUyP7VBCeT
gXT1U/YICAMhoV/wnFjlqa5TmLWE43YuNjgJ0CFzvughjvAE32O57ETdWqQ3JDfE
Cj/5R9RoqaGD3WnVTM5OZibGbtPzN4884sUuc8Zk4rlXSyFa4Pp98Lewl7uVdQQO
oiPkT4XOenI7TySo3YmisRohMjwDqrOJZNrPz5vchb4C6/hC2Z0kCsUHobaigsFE
/LTixGz40/Y11LnGJl4SMis9VN6YD6LB7533bTaIR0Y/KdLrZdNX230d6Dw/nMcN
rhcmUcfz5eW6oQ6n4bVsinGhnZwI5jxp3VRTkvVINgFfZ0IucXQTDXuzpRNJXokT
ktVeVtGyagAAf4DBPRfaHMUuFEOFiJszf+u9QvkvotK40FavhzpBf4UgXEq2mcnk
F0xCSqeSFFOZlldj6pIQLS9bePo5zxv1dhWPqWjsJH5eDomx0ClDahFCqnfU6imo
GG06ZJoy5ymp4gD4u7AZ325+sNTxH9oXmrvn71/yY+sCO0ca0wOlqRELjuhczUbG
kAZGwraoxIa4teu//8+LfhneZ9kO9AULQX6PyOyvwdvKOlcR0sF0HMeGIf0vhNuB
KSqQDTg8/IuraAsQ9+Dk0cVS7weTZAvj2WSeTP68r/6eQbzOvq2pMWUPrUNvob3Z
u0IOKsRY6PCdbl86KddvxehfFval3OFIcjW4HMHYfxKpoTDIyD5lf+mngPRyTGLq
v7d+2wsCoT9OjC+SFIcupXiwlZ/aAUrm7aNAgWAMuONhXcTgLJKZylcrdXoCuiFB
7FDfzfER3IgFO96OE2ahckuumkg3cvAYFDHNRZfW2TWDyB5J7QSfY3YF9UGm6Cp+
wE2tBRjyAkfkaRg4Nu3EBzVkNk5HI20RZ1gl35+UZlV/3zuLdWHgJIr2VRnCmZsy
UTIj1mzbTLXHdnFPaNvubuVWEdgLwhhGSB0CU5fIm2CrkYOYfRhedyt+79V1jHkk
PfLKn7XI5ZB26BUohUkEIWkjf3O8oA+3yQlAdvM3CYhwyVeybEevstVEHMq+eTFZ
1YR8ejz5KowjSCnO4/wjvdEevKnQ978aPcaY4sxAcpgOwpElXOoxp7aZ15jws3cr
+VuEEL1nYQgz/md7U0/H0jWo7SWu0XxRAbnCY/mKrZPbzhrGFfnsNlne2DqWH9UO
Pv/yT0114CfyTK3+mfruANi7SLWx2eypBhwKcaAbKivfGcIZMLyA9vIakNvy+YPG
TgfR8C9Ipy3+RYip7Klp1t2ctHQHV0A/fjQnFpRd3Ns44zeog8NukbUysKnM49aO
d+qdRjnJRhYj7gpG1qc9A+iW7diFimBAe05hM643a9hyj2MZhvaEpXgUcKNB+Poh
mYq5+pUvD3fICSi96YixCAEOi4IeuKCFwfIV2nfNq/o8F+3ZABLWQcJzBlKaDNqB
QNJbss2IWX1uMhTtv6WaNVvz2AtQuuc/ZSExwvzM9kZzfT7TS6Vhwtl9wRf9HHHK
1EmHuIX9Ok+SxIJk5i2F4+Po4VIuudMg2cdoUSaCW5x7XbGwp9/Zy+bs0Rj4ESMN
RMQRScOzbq0LgSau8NzjfhG+e/vyEB3bPVV6CdD4TWRu6Z0PF2HgwfATZhCzktZS
tLqOWZNlB//RDyQo0XIES/F3ZYOAeBzD1ckU938opwZkf6jARM3lQqXAPICanDpZ
80dPNLTkMhSQYiDp7rGsqfwDek8ClLgTYJ0A6cQGz+xGt3Aw6Hfk5qJg2/VWFsk0
AB3EbjyfZI8x0q5twpousYKiUobt8Lp8qL2puzeotj1YOkMTfUpPQEi7pluqvDgR
fjFPaGvSendMeX7gq+bWmjIzAerPZqcJ5iojbD75ucZacHvp9QT4p37r32aPXv2a
9bEbkdzlSMjGdC7WOOLHBBp+BEyE233vE4i/Xjbm8WC/hXNfZYQEjl3P077nWEhC
DY1iq2Uxz5ppIRozkAa0/UpDDA8n9qcgG9VU8TcB1gYgclBKGSJC8bE76DeM8jhK
pmh9WXzXJbBOkjdXEh1i4om5DjAqYHUbWYN7UgVBgB0sm7b6/7a4ytaTvUHNVVR9
0ykTr6VA+rtpnVJx6nJGMIHAVP5RF1J34NFDcq2g3f2FCImKYbiYahxCtHgoTIbZ
w2+r30XsubBWz4Wq9YN2mnkdaZvT875MyyUqoTzWkAOqdjpVw0adO6fydckG9nRC
93+BSghrJe3OUu1HZU+pj8YXCRVHmpXaKRXvI969rmA6Bb4peUZ25QkBaVlryC6R
aZmsYbdXScSPgdTvtVmtveDqPcpj7bp3c4mUQrs9Ec4tPdxHMoC2oBmg35wx7zYc
9jORS5eANB0Vi8Lu3kxs8Sd0z0OMRO73AGJ4pMz2yKSn+5Tb5lDof3AD7idxp3+4
k/tSJCEgnSdWq2+AWKOdbSaQoOViVdVzjQkCMRwyfDlqc4gWQIwXivuGQkPpOD3X
g60w9t0M2YLq6h5Raoa5hv4fzdk8QiualPza4NqT3lAqWrLpj/lgo/Iu/e8GSnJp
fXQFNxKg1dTddGvo01l9e02JS3bwihJry9FBW+7OqIcfftx0yxehEzN5hW+MULKd
rAYuyGQ5B8rBcighFkJ7PpEUY42CFE/GEp/BFteWIDzmQZmIOJhNseNH/PbU14Pm
3pJmNbgP1AkhVxAMll27P5gjt1OF2jUr9bPKdtMdtygivv7kE31gxiFtHngVVcd9
4h2Up9E8WLTzoy2nohbakaVrnYl6b3QFjuIUn+/1/NSa9/+XKbioyWn9BfUGeAqP
73rsBLRLpsf/iJauDTw33ECHQ/be4J4C8GL5BVk6GKd3JVyas8Q5tfdVpvxqwhmP
9qc9ufMPSn+rva+TyqHVBdAw5cq+dVZ5LgPhWUf/uJcnA3etXRqj4wOgGhP5A7MT
K2rHbRBPCU5m9ymG6Sfz2BpAePXdyHD8iESMUw3QozSbsqZ7g0v9gNk9TkZ4xS1V
KUqItfiJ7Wski3m5ilF+mISVE8KhBbm8mMvx8i1WQG9beFtwJu5g4dAclFK5U3WC
tKWJQrvON3x5ZBQakk9pZDNS8rxr46t7Z8byC8sDJ8UwcssTWifKTPc3gNu0Otmb
M4IzKtidem+72nlggTwtL6iLrheyonOzikjM1QQ1vpwQEJWa3ZPKSqJai0gGE7Pu
QE+HTPptuew6U5/hO7xW67oatPzBQMFbvIO3cSnU1IVpF0FTqWzaK4MHFWOc4pAl
0FdFNqMAz7kuSUR4e6+lM7b8smXbK/eynian9lz+NMFHujETDmyXHVisPWUT/EyD
Sx40w/IbU7BvCvHIqWlJsK9wdwD2UkvBVHbkiAC7YcpDxE5yRFPBhtqsaQv0Vq1b
kpBoILgBMDyiJS91nEFhUdOSMgp47//kHnmDd5c0XRRxCor2l0Ym7X23JN0rsFF2
bvbtECry/T/5j1V4zSqiKzAvVR2KYqll5ardLGUyC4dTbjHtuyNxDg3Fycbp/djK
x54cgYIJvPnqeHG2qaxIKV1BsKJM+erRPtApslL9GplOD3Xn00L0BLO/5ZEKxN2O
5fFh0xEOQYMNhHl5CA8PG8/KsOzBSvhROHCwd5gp1iyOeE9S7xGGc1eZ82Cc2vAC
kFs0Jl9E9h0wJAR+6aU+Ox03/BYBmvr6dKzhdD0ptdmakxWFw8wqQvrcEv1sqSgZ
EJYEH6smJXvi+3eDKUYJqrVPQJsJuaON98fegbtXnTJ4CXRYVmhFZF6EKZEOv3om
v3cDm9zRia0rjq4JKTHMoVWoHQGz0pSx4i6IhRZe/Q0uWFjD7nBnVfSjtAhCOTnP
PajdFs6eh2KHDm2HlDgdO9L4eX5vZGm0tjVpBzSVOCc6c2VVR7dVgQbJz28wcs8A
aJMV96OokawO3DPGlWOo15MW6oIpLv2VUiIUC0baY9y/x6q5zvNKnrcVoTdfrZuz
mfiVzavHraks80L/f8D/GUS75T3FQfRcgXwUIJ+muikO8nC8LgkBkPvBVjRPWxbW
G/d+JyIyWGANvJzILUnPEAHrp4OR3VmzF8+8Hf0N17HVsmkn6Kbrb4jZRzKDOpfG
vu9va90qaORBLuubdOvpkkwIxSojYuPQIuEN/4MlBxmAbxDBTLEZGhPJfJ57lPIm
E6HQ/ylz0uogQp1CLF1Uze1N0A/DvGoc5etAn55pr2AKi2GnPNxZrrZe8kaZp6ox
qbFFvlI3TRRlk5ftQW5R/11gYlQcID7g7P6B+bA/90maMmKMsOnZwxbsWiwA3DHq
/BDUoIfTtuN5+d6yBDD7oxaX6k0PHCNqB8695sUNy3EckSa0G7OxF4UrFVVNabtp
NcVSNPTk6pLC6Ie6BzWo1d8UCE5yIklzAHgh8gicHtGrQ2QUhTHciFFxcSFcrjVB
ZQdxH80wv2/FL9TnmoBuIIYkmh+HgvxXzoHCAnkjdev6RGrmMmbIf0EHTuOqP2tK
4S2uw36ZCiaoInZ3JE6h/emBwwZKquZY3U3c0K7DstGukE98cjfvwoUQZDrUXgUP
0Pfj4X5k2lypenPfgyQz4Voxv/NgbMqy+At+jZFR5s3fXrmf504O4gfBNvJCjPj8
msQChaIF+tPnH50hDFKu+tddX1SL2BNiSnMga+wKPZiODSm8/8NkPBdwN3ymJrMK
M4Np9FPk2GmgXKBXD0G6Cf6PcM4UYEALV9Sbi/rJuq5HzHfvOnUh7XUMB2vouHVR
fuKBwt8+esDWIf4HHdDnDOEkOP16hy0lXwBKNTjLdHfp2xXSrd/r6qtrjf+ktTf4
dpUoRIzHGV/l5raGM8NBzBAQEnqz97vgTQ0bslkhmFZWZXBOaAzeoPKrS0Iul/Qy
qL+gX4F1rIwSKQBkKxjC8SwZCx3364Ej/+1RiU3eL63/6ZGYt+DhxEgguK74DrVN
4dp6HMn10YCCbK9WVbW0QOp6PZuu8mcSkcOHIQjzyS7g572Md4JW951Qa4CPTo/L
3OHScgLCWRYpO9c7uJF309WZ0B30QLZyANpqr01c1ontha3CRiovNZ+/TdONxFFD
h1n1z6GuV3l0ojvScWkZr2M8fsRimwxtptTW7+kd82g4ZLO9Ck2isDFX6Ct8U2gc
IgT67AFhkIvF2HZa0EsebJ8P+F/9Z04iBG20rimwnk04yFdgdQJ0ele7u7SvnwqA
jbIqLBjs9YMA6ZkS1I/Ko3kTc/qmjHCj5Bz+RR/akqDYG3aG8Cn//J4jEGEib4Vw
qTDx2k8UFg1DgrLAmIRTMQvdqaciMeK818JZFgToDLPtYsq1uySTyUkRfpHSH2N2
YQiPxj24uub4EqHqeN68DezoY85qXtXRCqyt1sQOGu67lK6d+Rxa6aRkxle67K87
XADorY9W9ZtMYSJ8+YOxz4I8ZSkkY/3zIkByOvLF4KnaYR0XchEw1qLx1qPGz1yK
GeSiREpnsatGtDW70C8WlSFrK8yBeKVSpspUPJDKFd6AJdDoPesKhvmu6BGkt93h
pNaeL4gzXPeTyJbxoRLFp6F1Lu+FbIKIlYyZKgQzfy2DE30Ffo8qr8CLV0oweqmv
nC8MxIBWjjDdu2MSD5D+U5bS/qP7KzZINV4uHy6xzxjjgDRva1pcw57/D1o5bDtA
fKePBQ8L5SetFBJuo/HKqUpT57nV9GEt+zGC/6WjVUOt1wWpRD3sAzoDd+DGgQdx
BCm0YYHrnGfDfaI5Dszhb7OgWR57EHXDvr3GVPi1WM/1mTK43+0HQmQYDUyqCQef
0UuOvgI/OsD9KgvC7Crb7ASFAN2mBRaFR2CivIGVS9hegPxf0gVS8izNLEiwihzh
ew2iSF7+hcVJ8sTf91zZIm007E3BJWrGbuX28/fOCAIx3vVlUbpbQnIfKZn16DDZ
8uxQ+FlDGT1tgSMkLKSYE6ZzkUonrjy02MJ2wiCiASRlIBER7IiWUT8uQBfliUoI
zqj7HtsqG851yzfjrSyOH80xt0qcBIerY9627lpEwU69rmZ1I+zB4wg1TLoaq0Sa
fVE75YzSRI4fMRnpBgXoHAN/Tdq8yWGlpFHLfSklF0WXAQ464L4jNhazcOX+sWBE
FFh40Fy9dorgPl31ZXpEHJruF9G+e6kIP/W8P7mnmMu/ZIBdsYOSnnF+iLg4Fs0L
zUUMJZ+4akmZn5s2ATiFw0Ue02Y4cWVjbAJwZMD7hbBhCoJQn303Oza7FZE6LSEk
G5EWSLR4pMDFGrT7n8XrfGCEpk+Xxwzff2lmzUAb4mc56tG+0bWhSMGBW6tx2kBX
T83+OH3TFS4u9uz59+uRYGIzG1QvNckYCcAOYdf5Usr4yOOjnKTVQnt3HjxaTQzx
z507b76e+7Z5H2ultoyRLJi4dsPJn4XRFXMuWzKqU2pQ3HUPf2hbNjhOHoTXpXjz
eN1QxXzkL1N5YnCpXoltK0fT4WpklJqw2YaA8vTkQvpCluYWn6l9p0r1Fm5gwoFk
6bGKF2I+3jAPjCku0YI+ePWzyCxJum7LdOuFx6HVaZEXEw7C/UF8S1dPcUM0e+pu
9s4rr0z+5osQ7aPUENdU5+AEAQO1QmtWkOOaducnruLfnAwN2ATWpFp17H12IZIS
MQFfc3iUBWsNc/Gs21WLjoDXII8CDXhqjDGe5jsoYTEgsiwb+HEUqyrkVgHC8P4d
IPK14nBOeSBr5LWr6gWArplkq8aMjBDJ1y0OuXVcMw2uJCRl+9qBNQdVmcPM5bPz
cOmb9rpUqShLfqxA2L5WnCir6Sb16cxx7I571rIek9j9AC/meqPkdtDP0lkNhH4k
bSkaxROYXUz6j7xvOd+uMbsvVgojwhQKYiElQO7Avq7cxVEVxvvaalNhC2f4hOA4
uWAzesHAqME3HyqfBGEmqnHExOtXTXtikHIJcAeiQGN9gWn+dgU0vdeo0pf80WaT
2Qez3moYCdfNdbW3GEJTsoaUC9vGmLeOF0q884/kFMrbg2tTNZfFSOfnW3k3IINy
BpkdM8kyKelgYect/5BnRDnlZBAl1NNGTUHF+CiGbGJqaMfG60c6QHlACJC7T3hh
0A8dj91UJCNvwUQ6RuDHizkZTq5sVua9TlH73EgxqBzsK6/aCfb664z2YD8jpRB8
EEO6i+j7NGqDsvSIUIpex/OugcGs0/mpRsK8nFFAA3a0Vfo1lpP2XL4NvxROqZuV
KVS49U3H3PqzHaowohJ1fC7wngLPhE4auk7awjZGbsPYZ44+7YOk2O0u5m09P/hI
vclKK3gqs61athRry378xAUGJiVKE+ZTpC9QK/1XtBkQQ37wpar3seN1XmAb7ojA
1ANVanT3ymHYG+uz/wvyVk9hCRruxcWVLswg8SGYAm2kcD058aTFtEUEPXDysJxg
hjjor0wrRo4CnxILT46BJDtzsrs2Kl4ZjZwYR/n59ayEtTc7kHYkAz8LqseMN7kt
np3OWDXd2oX2SH7P9h362bj8o7tHEPooqIGTBuoxuduFb9iKRa9zQcZuWThtyWhz
Mj7nGED5rasZkZs15vnoFRqwsaCh0Mc1qCjVp0nL+tJ6VU1FJ8Ao6IP7XxvChEXv
Eof5sbTX5uehZYFNid9klfepkFysdawRIv8DCvhELHKkz/1YR4b5xoAtb8LMTfOH
pgeUREjyNB02wZbCajZmH7X9t2Z4LKYwmbn3j7cRDuqgExHI6HlpUNk14vTxhJYy
fZjwToJ9njsVksr4oda+NGEZG2M/MhxmeC9qQFpDYEqWKzdz+PjCZqjuza7KJEuk
LGHSwvCQE7WvllzXngKvPY7Ne+RjmSzm6CziA3ia4OfhZmzLs5ip9G9PXai93PjR
GHZfckYlZpINo6VNN/SHCcI5OGz6F3IB5ooW9NvouJmNpMfkpTz8LuBwK+zG1pYm
SHGbb/vkpTpRm7ui2+lGiuhdNvIt+WT9u3jQjeYiEnw73CfSBSXAA2Yt1+478HvK
qVdLesDITnS0orFGNktun7gxWXKsin/i2eLRXfOfykEm8NUl7pmPYVKGKtz60mZE
TMGOVaeKU2ZB7vTTOD8oG2uCvzYltcuV9hRuZRcKmUvT8kZdHhB3gygW9EfcLp/F
3t/a0kOrDCbZYimCEA2dcy866eU2Y+55f59ncfh9pDsP1q9dchK5+O0g/t+vfION
u8tdDN5Vj4FUmB1xDi+fcXg5l7D/vh5y+r3io3Kxa8oSpmxPUzu+eWk6GRE9dhoK
K+0Rgp/pAH5L1wNRISt6SyK5OPRDyyswtP+/H7KTdHZPSxj1ZRzMklxyw/ul6RBV
TxC/wn2WL4lUPHr9IguO9OiKgXiC/D0XIbcLEq8oLEr9b5ivW2ybzPdiMc6k+sFy
1muX162iX7dWlY8LtxHuN9nYMlJTnjhrQ5Uy0HREcaA6xzWN6rPA3jxK395ZpRRU
1J3uiJ+vH4idIhVxvJd96c5uk2x7XGrai5Zei/AORL6z0KNnwA/cN7sbyI8OK1eZ
fh+JoecjU+9unEoXFUl3JeYZDmDXLCmNctpLmve/3vQVWOo+94MRnzzrkHq8uJ1Y
4HCqQ+omeupnvhnRJgOcjTVRs9OxnbJ0G0N/r/+HjhUfMBgwV+0eXvpcWxtRP2jx
6vaq/yd1zgU8ZcJFjDuCpXUJ1QodMlOP/Q75NtwEoewGeaI3dwfY0urk1GCYx17O
xC4+f/30lnPEHOXD0f8p1fRpnY6vuM/98XZ/vUOyawP2ro/9AXseepXJNHq3BWZx
+nAFALpi4rnZI6pSNDasc2nxm9lYXH8Ddh1c4iJJCuJhKpQeNjTATxc1Z8S7c3VV
N69sK+61DRMSAdsvn7/lMgHV1pzdgDaKthi0RKjijmw4eM+aULDEo9OEHDJsdkyL
y9Ma7yTkvty09/7DC8cXTCw0VRanmQ5veepcyrIFwoUGcjkx+XKb5fBm/edl8/r6
6KEYm/YqxeG8cYMmEktz4MhsIiIQrbWrlBHtnHyJPOxzrfQnIs45SaZNpteTJGTQ
WdyKWR1mGkAnPFGGo4+k732oGve2b6l2SozF7jJmscMChAk0sXLLCFBrVT40O0pN
NM9wETaxCeeCvK6hhH2G+KzQftsiHXxVlndJQOTLjAK7QJxDMAq6Yd3Sit601WGf
/16nGGjDHhDdtE8+lP2AJx/LXAgW5fmV5v35rgHYoIOiwQV57PCj6GCHymTZOmYN
KN1yRBCylFaNUVPOZ8KeEf+ed7pgUOYExLrW0y3ej5W4v6GRBkyON+lZ8jYcYP2M
u5mtKtBXt4w4OULS16G+oUCy0Mg/Xesgo3QSjYOnxdsCBPNAupI86ARq8zt5RQ+A
IApRsapRE0I6CUGIH37+XxOqs7ITirTal2+QRhdo5l/5ZXC6LMKtdcMX3yyaBukt
jHmIvt1kRFZa6CHLtfHPWpswwxAKNMy9Ks7vKFFva/pM+xRskWj6BGlZtIOmtej5
b0DzOt9tZQ4WRdel96F4IzakyBxMJdcfD/RQBp4QcbUExfbyL//ZHAs8vPce2V5G
Krbv0nl6V4pNjZ5SDwb4moKPnOygFXl5lLrMpaR7+A43FmUV4QhkeiwJDnmb2crd
23P9sMG8cAWNXu7lR3/vg2ardR1Mq03J+qkqvi8CgrD65lOFNE89E12FwHvATPB7
aimyOmOtsPEST5hkYlA43sUNmEJzPfhqYYsdzwZEyJlLy+Zy0Zd+C/VVGjKg/I1M
4PeCGV2vZQa/3F9Ln8fkarqY7+D8JhuoxthN6egdwtfW/2g0T5fB7cMEv/ngdywf
+V1HYkYU6Z4d9oI6B0Ix5vpXubzxGwbFcym2EjC4+yJPpc4289aDUFC9k5qFRJDL
I4q+hZm7OXnJf56+GTcQ/g8HGDNqm9Oq7SdjxobrJwrAvy2zoxdHeQ5Tvr8+Tklt
SEzF7p20oVVNtNxTLEwANP0J4XPnHncwwcUaW75NJLIqInLlpH1pExZmkZWtttLn
MHOWPQmzOYOvqwg7/bjiCe8zGejJyx4fK8pbc+WdiSH0w3gO9Cyw55GBLsAwnfDA
pIR5EnKCi8vZ3bp+77IQb/7TT6zkGZ5HIqaYkGA+zf04Rm9Q4L7bLyj+002SO0co
cOQZSyuHuR/ZHGO4xDFifhmP782gL1mdALn6QmBSSpvgJphZDBTG60buFKlMTb3Q
sFcMko79Hvb166TnzzaUHGvamATdY1ix1sGG1dEow1TeweG0wnSp2I1WY0dhF5a2
kgZe600eyc2N7aiY9C6PcwMZ88w/Fq2x+O3jduu9IIxYLgW4VZ/g2+xFAJNA9hqY
ZpS10PgHG4CBWiuJLlpFAJZs+hIL95r5FXFHQjkkM+2voWbnLC0IKZtMSf2awzYA
ZGNrTzegea0EOFZbPVjjhgyFluw60qDRUACFpRHv56w71MpqJPJE+LZgQ2OUmz8W
kfSGIME3ykL1xmmXsag9X2D2Ei8eFAPfPw7srvj0xaP/u2cQn0SfxOdjugzPpq4A
Y01TkjGsHzxCf2HadQGFv9Lhn0ph5kfiZQUWYkucdNHIlMFmhV88KN73eH++Cv9p
Aq6zfn7U2Ec6VqT7XJZynO9eFSnmFHjzdT9AGNFfqsJX7s+fHLfKC+OzQXkFesaf
HQM+jxw0ZOZE+f+T3RvfevJ4KAzFzRh7iFTGZ6pLR906X/YiyLUQdRI39xXP1tXp
1R+YILDXYezgfo49P8qAqt+4aZxLpV4ZtXfXPFlW2AzoIhRQoz66e2c+g3F4Nwum
ai7E7bWlx5kZGR2DBUGjOXEokhwiqxon3pyAn6mTnOsxzz2yrXx2qq0hOimX44kv
T6aOw6Mro95SwRnZBCx30kUesJTMUbcdgoP1SUavIAlerXIRg4FrIkrIEqZwiH9T
DWJcUQWqYaNjsn1YPYxpCwvpYqGMId/Bt1QaWTkgW6I47BZCP4f7ca+9K1HkVZnT
6CfT2fufNMjfJvBQDZ0EluuEwkB0wqohyexiLU0E28DAzDRCr+tYH1vJPZyjxU6s
XVMXUG//pVImCQ53ZWi/KCQDbyHYprzgYKKUllRhN5M0W14Jw+rOZBVzJuatWMyx
/wiP4AoqpqYfNydC/T7Kv8BqeKTgUTzrQbv6zmyVc84WYDHXQ1uzSjkq01uANqex
eK2W/ocJGzEjXI4Hr2hzlS0UJXSq4zUlmObezUJckDPDW/cYRHvXwjgtiQIhOnym
LOkEyFMReST5kkemtTg+RBF1a6zGpgAAKPf4Bk7PB3RMEoRvq9s35fsdOUEm3aIC
kwlYseAQ2364nraCS5S55hdVvmISlkukmT4N57HV/pg8a15lLMPpKNq+ri+OLMJr
JPT4YDGiE3i64wEWK57v1s5CG8xecLlRMS50hHLYLwpSTSwTU1EZvxdzpDRogb+U
svLCyHpgtMWeEy5AHRuAtpNpL3Q3o98ZNMWF5FHWcH6KkXZL6XpqtDjIJ3uA86dg
NUstcSBNX48gc9Pa6Lns4VLwC6qQjNiBWbGyaC6sTWlLJ2PgLASkpzvKh5JrhVK7
thccmP6m6CwshHPSJbjFOwIT8dvGmemVYKowctTheKnKTVTyemtXpjUIFEysIaqY
P7QA1KQkSs2jcY3ePJ05Fo7+WrJRUH6YPj4QaYia0BapbDvC2MuRdZ3r8b9UbLDY
3YN6h14ZSDl8Ci29Ku8r6s2GiqhbySHqqENdrJLi8wgHZEHzHJ0oCMR9FW8gyW1O
jxlXLU0xIbfbaa5S1NbHMYCrVtKUGqnYb8zf0K+FYaCg09vIgRvgb/g/FfqsKzeL
Tw/ItGJNNd43W2dZq7FIgcrM9Znlribg3++d/72TDIGqmwfFiXYG3O99klcUqDlE
cqMBQMPI5sN+ofhEDm6E9KYGM5veF3jTw6irUiOK6vt0qBmIIAoy4egyqV2pjMqK
kLlhtHQrhku+7rTQUduCU7d/oUYCn1usr+PzxuJ+7U/BtO+T1QoS3MohtZRRzh20
4Fnot34hthUuDTcnEOSytvobCW3Sfpa/Wb15r83eFJhGdB8Wzji1L2E/o+WtYHmq
IrP9Ll0A/pOr1xuKAPflWoCj0VyhDg9icDx0WC8eIJ536B1P9GsPbHaqqq5Mi5yD
7dLzxutJdDSDOOJvmzIsyaf0AWM5UmU1tk/jS3Z/b2igWtmeBiX4BZC7RFhYsEhq
iB/mZaArfZ3mq1qLvwkmRkN2M+Q7aqMqsUpVqnpC44T9FxjxvPIbNl/V9cpDsM6x
k3rp+PPNiGRkTbjI7jtsC8F7cWJlGlx6spuO1/8ZamrAJiX6OFJAUc/yC/Pf2b7i
TTDQrDwcgGU71vPU9I90U5pfCIi7lbVrTOeivFPwlZIfTEIj7dbogy0yl14EMpCu
hScZ6QFolsL01FHlI+yvBZcEyJNmEJBtByQbiv5pECmSAip1xV+UfqyV0S7Ma8BO
LaPIAQ5rOIgFA4rcOx7NgBph9OYLVGIKmkvdPZwN436IxBcvxxJ25eLYwqB+oxW7
E7vYEIO6gQMmv4GQQIimoDOdIv/qhI30xWMuwC1LGFOPwMTsPLu+UFl7Vuao9nw4
pOlP7othIkQrfm1aADksVkzY5OlYZe26rvoMT4gV+daUipw2IfTDKEuW/7vHXgTq
sDpSYgt7VmWoBdJhgHgl3D1/zhZ1ifs6TPOkbEvx5gt0QXM1Uu5XAnUl+ziWadHY
LOSzIhPCuTGCuyI3yJk7NFhSzCkGf2bsiCt3oC8k3QhMpZbkZQEq3DkCYvTyTLqw
EGZmTqNssvVLYcq12PCrEC3CIExqsMghOziYNXMmigmr+Uyl30R8xZNv78r12E+7
8i2w3BHBl5jqOTt+NGR2LJfpvlz5RkWXason0btnyU16VZMiaZPSRFobi7bLuazm
2uD43jDospAL6vW9c+1lkzX9lXIEZeqgsDXQKWQMFsIneHRXodXeNCGS0Jeoo0k7
MDd6UdBkYguG5E5Z9MpopXhmsp9l+OmXgO8Pb0bsTzo9iAApc0zUTb1+x7MHxtFW
A0PKs7X2iV3RcfCH85dqwuYHvhAuSMx4VbDE6kUBuQuc9Kk6kKll3ZiRXXXjxT2S
qnTHWYWIUShW7E5+cXu0jI4YwwCNVzT7OJcXeDBOK/swp6otx8mzV2bSADpPi1Zb
eUXD/2sVDuuvM4lgzxnfBa9Lx70j/VSgA11TH69RRgfm6aoam9VAB2xyrpgg3kw+
QvdKgUaMTS+5HZrKzyQCwhCmFjkVHeToOiz5tvQKFReOH5x2uBYijhXHZiDi0EDq
5VOW4dQTqUCecD7HLa9sFzacZnBrxJxc21+4NMT5psnPtQowkk0Qw2Tt35MbFnXq
Wz36D9YO/A/LBopSldeszMV13LmeLzRnstgzPvONA/KtWqLQ+uPC9aTHl85L2v6C
zSpD3VFmLL8n2TpeKzXgoxnfqOmYfx/Je93LO8jvC4D39QkKiGFg+m9HOHs4biiE
toWbAdQ3g94dKmmr8Epl9jsA+DgsEbiFFtTJ5AKKr5KhTEjPbOaZGh60moRlZ5eQ
F29jUvP0ydMdsi0jco30GJz4cWS/EZx1cBHFhUhU6Xs7q0FPGed/Svy4lL4qc/G+
NBz2/VsMRTsy2kSYj9XmJeL0lgpcMOQkW0mVZQeXrWId8qmh3jsTQ7/aIT4mPHV9
z1TRzPsYhqo+T8NIkun8szKSO0SQA8Em+tP8TIq5pyB/dnC4JD1kU29GFJz0FbLu
lKyhs0Q1kI81ZDJ5gGAlGRzlozU1QLXDnme4ig/5C7XDRwllXm/dqUgWqFygLNJe
D+cwfSXxu/PGuHxWfTNp8FwEX1V6Ghf5dB6NX2ro4UjP0CsdNcFqm5sIJ5OJ9c8Q
OJ/g/IAgB9DfMIckspqYNO6dDPZz2Fd2YePIZJGzYup0pgB69N7vmeCcTsKDAvBX
i68r+y/RPvwDUUnnPpiv2WpJO84Ku2BX8i/IwFbZDkf+0SVDCTIL/LYVe/goinhI
ukEAQICIeo31U/+1uf7QuItXg9z6dFQ+b0gkYEoIZzyOlPfu9hX5kKBFvmf48UEn
zMV0mjiYenO0Nf/CfmgToRhir/4woeLZGdJ6VdNoPPPvFBIT+/s5Hj+D0jbNeR8F
4tEoptwnmfYOLV30ZUVzVuctShJMM0Ti5JP33N7JDBB3V756Y2vq2p3OBPBho9RV
kS+OuhJUhNZEgzC5iI3sPavy8sgwkzRMEqGh4gAp1VpHbotD2brX2bnAlBFtRUIn
+oRcDwDyTLJzZ1Ti6LIPPs00fR1kCLBZs5fogXZ5UnQpPSnR21CneIDlNQecrhvi
I+pY5i64B89T32VYUp/tQ8e+wV0/wVVI1ubOyHk2SkV+J1Msm5QE7CoFxHFuxKlE
WWvFgkCoMUrByH5SFyPlMV/NDiGuINDGzuvTshODrQwqouA7i2MFPk5MfjeiV+XB
cvUNPLpn15bJYJXLaEssW0UhhYBKFRnLkZzHAh0aUJiwjRtmF5Lc7L68WnscUZvi
9cyzlmlfGLvw4wYUkbDEV+l3U7Pgx8cERWiNTC5GodufHdBFHw/w/FdAc7C+8+2M
qOgct748u5Cg/aee7eZnVo9Q6MdG8Bk8yeCRjwUnPZ9q3ul17vbDcT6iTNyvzJro
kbCbuHr00Zp0Z7YxdGz75sN4cG/QuLxaL21tUcKIIylYXPnPAQlHr6h+SnFtDNL8
5zbmsbtxO7po3Qk7XUoUZFGgD/K6CptJq2057i5EoK4gWTGiIh749ULheknoe0J2
N77sA+7AT0Uf3OVFxi/BeZp8f8qcXNTRBVkFZI8fOL90u4UwN010Ne181Kz6G+WA
wpj9Wci/LO6rNUoYIYREUN3rWlKUD0iegnedrttOZRv4Zu/ZtAbwkscHQeHKrwhj
99+qIw5fl6mZOj/BCxhM6d1VcJ6W0Glu2Z+xJrOjKVfqrVw8ebWOdftbh1oXJtcD
3qb0WtlGI4c58y0BSANEKvUfUisVFsGQneTsusDYpU3H7Fhn2A7fTHxEoxilmPzQ
ylM6u65+NY6KYIG+iOkIkXVwCJ/wGCn8ivBdI2W881+D9S1pQTs2pL4QRgFe0+e6
gd9QMV4m44wAw+djgYiqOu1YVb1SRrKvVFJWRceLZUwzecsTtS4QVzr1m2PQRqyn
C9Wqi+EEOCA3G++z42JJqabgE7Sk8pLEQQ7p5qd5rr9fNy82LS3tYpfpeUjrb6ls
4v10fJn6Xhb/SANKxsz82Epk1gfB6+uYh+9OGV3mLyPYYI3s//tnDPR30cr83ZEd
MCaglKug8S/o7y0BbQxnPc81byAnGf5W9x4QspHQSaodL2QoqCWKM5hnerVGPh8S
e7UvKlGzjb0em/TlzJkZPb8YVdYF+tZGKZG1QnmKThq1SLaxaI51JfSUFin95ul4
zXfo3mziidtcnK04Tnh8dapmXIvJWkI6C1UZER3BnYW2gR3FMYlJSV7veRqr8WTe
ndGNWA+DsWLhTOKiuiXKhtLkmMqcC6PBzEh+TAIBbU9C6EOEOxO2A5AFAUEQ+rIA
wxv+NKOhEn/zHHv6OMV7Z22Oa8Wdp7HrbJZF0muhrAP4efI1/3NT86FoxUvTYncJ
Cl+zHqsXy2NxUU19sVyi+8TbYGM4iIy3tB4J4wCMXrfdvZNxHRCXMppFUHYm4ANK
qaffdwFhPCZaNUKMhrH49G9v3wcWKO18Nxe+pOPTUEwk7qr9G+226gvz2Rv8YfLm
B27gc+w7bEpINRGyWrKqelEQiuWfUoVHZB85lyBfscORmIPrRm83F/56ezCkU0G4
Mgzs9tgoqBAuQbpbRW7NX5aNAYMy4i+fYC+m8m38i3HBKd6wuyKGTAQ3d0tEV9cC
olhqEcZKZNeSg9gZAq4Ulefd2aH6dmXFh8FM4Ls4KCB0Gzy84rF7poJdpcj/CPLf
CXaXrZtcJyYCV5Qfh2PHzdK9oQHVCdMA9uBta5mFwHfbQdJ0Drhj06cKqse4R7jF
Y34OMspEwfkoTLKs819xBsmii4XUZV5tiqs/gY8CA0Ye+Al8GvlpihjQJnDV8krQ
sfMlZoMf3RnZdDDyuf8OlCs8ycL6YhEYSQHEyz6T1jc9yKLH63l+4PSGhQbvdxpb
CIdZPb+A0GelmT1Nkgi6AneuC+oiS+fBDbqdlxd89AEKLKn+lTGaj4Mb3wWNOGJ9
udi0w09sASuXeHZCTwt6UMyCKTqvGmOkmDrJlSE/49mqFELVTRS3BaZgjMniI1vl
4SRO7AnQcbVY5AC/AqHihbo0Url+jAcs5kniq+WPus8pCzpeCpXFQczztEGsSkpR
VnKmVnuUCKjvptUQZcZ6+k9Yld7hFyMJqz0qAge5yvtH2C+i/IL+kd7qhRL19llg
phsp2XKgeQkcdax3f7guVXTHJ9sVCBz/cd/KGvKgCkkrGSXMDbUmCXFK8T3mC5YM
ZQgCpmSYkd4KgtTYFozjNC99qSdrwBPr5rZeqsulYmdO3x8MT7iv3OiuD1Rexvyq
vKMyk5CnTgfpQKIA9DY+klihY82oWXbPsHaFJObh5wIfEmelV53ho1s5FFW+0tZ5
BieGxVHmBw0V2MSO8W9jLyIPi0cZkUUmaCFdUXNN6oiWEAqDTi9SWPn0Y76D4lgM
dWGMHTJYA66alkjWWQTuugWCcM5ZUCq8vGUX0e7ppwRqAHyW3zDlPxQWhCDpG7AU
MMRU/hpQ7VkxbT4q7xNT5HyqFBPE+vbPnQVTjVoPrkktbtGS3vxV1T9HdiWas8NR
1HlNuVKCsxAwbrglzPqYl8HI/8M3YFhi71soJ6XlDA6vg5N6cZ/CUlE1HgwiZucE
byCw29fiQsXTFNC2Sbpl2iA4T7lNn6UKqHLCCHZSsNA2DNfBk5Mav02iazozjAOu
8a4UapQ6wSO4/pVybPkrbRICNgtrClymyvBZt7qtO+Al9oHhLShdn76MMK/TIwdW
YTYeZmBHLMIVllh8hwb47IJFfJKYIgupKPowuQylemmkZ7giOH7QglCp80EzgBa0
u6c2ULdhw0CQnfpeE5PhNtIysnFL3jqiAhl1O0lhKwR+/1qwbTONVHTtgwakIAE9
alIcjE7jU59TUdyRjhB0mqFK7gal2ArL18CFc+9JlfHI31z3KUvISpROwev/KHkM
K15kPWGV+d3KcrqlOOAIYTQR/gfa5mCuyI6K4FLXbBhrED80TKqXfP6AdReyehVJ
vIumsyHcTaPSioDZFQ3BIGyeySbGz5axsLjMxhBzK9oNCK5t7jeVHt8nMqAJYkT7
WlBvzXMcIiQBNg4xiE48w6zEKgDo+cnHTeuh8S2V/Os2ZqO0qjXhiqOXXb2oIB9C
Ec2oDwGvBBNUm4phgu2Ak0SjG+6BnuR7yZOWmu3usKF/WrooNPxhDyn2CmdfXtzY
pAcGYs4jleRov+Q90EyDjA2dmb/HEKHm39hEwNEE45v8kNYrHzUcZfixPZXlgrlb
keP2Z2DQZG8v6WhXRFLglQdM+jhF+94U3U4wXvof+MugToTtnlLF07EbVKm5vfXU
jtD0fsJu7U/LUl5GFUb1UhMBYKXTS71xACrlPP6GoX3JJvKvuoQVxz2gfkIvh+28
OmYF1z5rajAr7ZAKtr6UAqYyK+1ezekXGLYcpDM5XTEY1O2Vi45TrXaMjN06rdhs
iPkWXjF0OVB7QkgZi/CWtZ/ze/nv3RUojx9gCy2K83O6zYcmarygULO0uYoOsoj4
JDD+nbi5re+EwvV9hfhYJXxB7EBDnluBQy49MClshKmYx0Als6jkiDaAwfJnUAKy
Qj1kACxEFmbU9r417RO1CwkM3W8v2JaAWUhZlI/Kf97JMwDWAo6mhYXDJXBjUSTc
c4nX1ruzrFNmtk0AgapNonOnbqMnxHxchx16iIfFnn2ukRAmDVn1UI1mEwGzColP
d+jgCxfusqBrHH9mrJNCauMu9EUYMMUO2En0yUmRWIwR7HGREQIvqgdsSMqsyS7q
xnUXtJpvZT0QOX/nvgOjgnySF0xO87zNaqzL/PTCnHVQR6pdxhE3kZmBevPOVCv7
cYsmcipmyzA/pgcS7IbeVu4LaSSU1aO53849yVmDq9t4VBfx37jPEDWdAdeWLXYI
7ZLy1wmZSltJFoZqOUC6xRve4zDD9eicZOjZ9Xoqv+xAjdxgnHI7SILqSgKsXo8B
sSClVcSGkzhW6c7BMSoaekT+tFYv2v1SDe8lsU+IaMoy/uNiHyWgFARXM7PyoK1C
Ldur7g6Zvo5b7qtcyhTsK0DxV5sgOr0rwKva650CpsqzIMmQr/bXEuTh3O07YCDd
Q3eFZOHUilwvqyLUtxEn8K1E7vH5km9RXyPLrpdnKxEFsNr5fa1I9lARTlw0L7nr
57mwnblUoheg51wsJ4vCIzC4R38azp6f8u4mw6F984fmh9JGa7jwkK5FfjQmPhHI
CTE3iJ2KIlNROW+/ykp5OKtCOH+JNr5IIjSMkyZPbcinjQdm7egiMcmeobgqGpOL
1zhlRJjPl7fyYQz6LKiEyJ6xyBUBSAXlCJM6D81dftwlvZoJyB2hW4/l2+4lga3m
/q7JG1tZAtxNfYFXPI0EkURd9voVARLuIewsKRsnFitA/70vliXiaRz7SigyfzT2
jTfdI9V5lBjTetI0mvMoJuvdmFsF1HP1Jers2JUmxkfuzdpxc+ZeHhnQOxMXMjiI
6yZGiqVHm5jQjpkhGIH4RedJVBhXah1nXEgS1DvZlU0zMfpRTBk+ckcSPu0deJ4R
nIMtC2NboxK5JmJkIW0meEsBG2+19jy+QjhB1oxXNJRGEWHO+XO3l7Z5IhIL4foA
sYnJSOrPw7fMUcke343oWqoDXc8MUqGX/OyN51i5cD3PVv7R/rtNBICNA7ujMIGS
kZiJ1FSyR9Mw4KcE7Bc/9PTs+V2Abvo7bMJWhJTcRFoI+XpeBlzctmgA7ZkYnotz
ifCo6rT+M6zuqyumaN3tEIItDl9mj9JGUKzmIFXFEqQihyx8E6+dz5WNDW1JKlbR
uZ4lUEgHmtq6OZVzOyX2GFyt19K1oJ15K1Z3JJEVQ73SbmlT/e5z/5fwv3JXIOUa
wqbCd6ClPfXc0mn5Ke07Ft18gMBOBoWSpg8fpNjl6YW+BN8WRnCxOrKk5IXorOAO
GnI1XhlASvOCMEg/UJwGmzl4q8wAdx7mqAb2AuiF9/tY0Ju9t6ERYRLW+ijEidb1
kbkTf+qjIXekfT2muFPpLC13g5pXrFk77/2+bi2N7qqH+As2vHL7/J2+quEdipb1
kCZlwcBr70Mylr3A3B3yzLtLqmcFCKjKK2t32NKtsdE6ibcEWuQn6Gozhkc99S/4
/5lTa18S8oJu82WXyQ+PBNEk6ktg9iUH2OiBJVOPFYpwssnm2VoQmWD9uELi+6lq
++cVbpdolhHnaenXAioBkxKeF5+VaMRAV2PUXP3kipvW2KfkucpbyefDmIK6lZhK
L413IPCTxaRGfCnzjM4ycOsOSRJFa39EzO0uyYHNDjtwBM8SgXVL228X/VEJ1Iy6
zpIqi/O+bAPa75/F1AptswELoHxQTXZXMTDCwm7L0/ndwQJjz+g3/MEbXpMN11jZ
YaKhvWbutVopQLdlRAckrZsL+C78P0ftT0BgDu9febKzUlKgjJG5d0DKquUMmPKB
xeHC4wUv6EjUJmYsFvwi3qbC0vY231zOqVt8/ZtoPx7OrMpVGjWCz/Vf7c5tpcAE
PjayCMxpU74oNyr0flb+7pNPNpf3A6b1gqeUF8GsMeMz1kvG0tJ3TzdLjNkp6dbp
efrAQ3z43FPklL8KFFHNnlOCz/J8uO8hEo/gHZzaqICNAAt650IWzTdSKf2ze9QF
2phyh2YpXC5p57XIq+VHh3UY8qcSCTDpQVUAh2pjdiMiKrQ+WEkkehG9eUxd3FB1
OT4KKYxlatWe7B0cd1hD00p+K7upWywgwFOvVJt80dktFLx5bvzaCA9jEzVPHVEU
8Bu2rsz4LTcTnQOVqPFepcEYr4NyRWUUkxdSc5/y9gSMRxNQC/uwiJJjbVaUujYN
PU9F9e9UJxDe/r6TMZ1kq7SXaIVGTqUYCqicDkkYOHwbDBPj3YpB00UxvQx9eb13
Jxjg+FUu9TF3r7NdCVwpmTPD/azIVhfJiXoXSSJDgAsigA/OsFs1R4PYKfNkyIlB
DeOrgjGGKB91FZYyPaaxWogFhsPrG9dBpHFWEnfJOtzfOViF+1HbpO5/Qjt2cM9c
4IT82txuS2FaU2ZOFh/FnZCEzf5D9odCq0VYhP9ItQF/uqGU5vr0zK06cRPdenTZ
MjIOH4feDdYMvZTLmJtXDRDBoRr4IpGG9sb2tj9gX4CUc4ZvoXw1vBjQKlQ3sY/A
e0O7/iIL95uWtmZXhRrzMa9Dji91qjCpVigc7KYPEy0NG4CtYV8tmKdBeIk2yman
1nnnaj7ZR3UaEkImZp6nHM2kBcLCz20OCm+4ZYnlbX3yqgKlGzy1TYbTR7i0pxA2
Cla+UWW+N/SBQKn4A1p9hSj+rYcbNJNbvAUGYBbOmGuW81sn+A9TgiAJx2shrpNS
4bOgHWz4qXPXF4cQhnuI/tv9YK74rcZOM3wxQQSSPuOKz0t9BZIauK1PBDivbIfl
6egzG2N6QXkiIt2G3oSVtPRsvTedmJHJ2cGBqUz8eNqnAm4eeH56uDWD+RfZmlGp
Nc8mjODLKBxNG7qBz9N7WTLSSXq7rI/uP1s/CS/7CYRtgQMrilmhCIBIbEoNWZ8T
iWscvVqNCopR8ET6/DSZ6upi9y3Juh3rZS5d3K1c0dlJBX+W3vZj1GVuqrnoZBQN
iMqFcTnRkiJz8nSpE9t4tgbeuEsZ8CXWVaXqOf6w3PjSNb3UKfch+jTRKhAfwwm9
hv3R08C2HJ3hwXGQX9EkeYgfFiOGqhJoqJ0QhXU2diPESBtKgQFYpEBjjO+SR54B
i5Vw4PyplX9kAh22g+1bi+CaddyHR0Ub9xkPefrMboYDfpGPPC1HtBsMYbTCtxRx
GOGdhoO+NXxeauhZrvFShtBg+rfcrs3klnkPSsq0wsZNLyfpNYkXOoV8cfFFtJYf
IvjyM5jYkcw6J/1Lsnj57aw9++LM44nnWEvYDTPkfa+tLUu4SamZuhP5KrnC/n6V
DpxanaSGY2h9RZhUSQnYc4WIqwv/fQN0LTcc/daZSBakHf1dXBWnUxCXl+xrjfSp
cThafuZSTdzRgGdjEDPl6oKAjCuL88UntP1tHm9WC6f3VWHBWKgZiMmXsT3wl9yy
qz4Uz0jn5lVkaheZDy4WxjbnelkV70QBJsYm614SZ2L6NcLoJy1SCfygUHJbTz6J
nLjiAQRFWXA7pszmwXMZkc1CMugipDmi2EoqZ7kvtGl0LwdJHUPrAIZOvinFYJH0
6e8PsbRwdeItGhJc7n2XTqCWK6GBNomcH+ZtpUbxomxCT6aKbntFmfVbUsMWM8FM
6ZVv2tnaDSORUGvKwU4FZ7XcA6LXFqAtaePCBS6NnOJlnuIWKq31XkfAVQDIK9K6
ECuRXpMKXAst0QpVUZeIUd16nxqmDnRSJ9KOIQvEHqqfT7WkOPYNDB9HrhuN1lSf
HqdbEtDzvVJgd+0ySbEYxtwkiS0WP4rm2hoT5/xh7QboMEAT59A6wrbH2BdyTeNg
eXqLqfpya1G/MZmAxuebLhiDr15l42PuNIXdVUXBotLtXND4LJEwJ/TyLybxcJsx
Gx0Plkz7G4zXsT3IZx7n5QLTHcQS80uXnSuKPrycKTUnmRAdj88ZY30WvlQtmC8r
EDWXwQpfQcIpXn6MgEv19uXIMNVOaRK9/wwjk+nS4Thzjv/KO6hI6vWbzxzp0URB
wgPevuA+c1A6CJNivplAznAyHSrSfbOh5KY3BZ6obohMUoLUFyrM6g0J9kiaN/ky
FXExP5AGvYSZUej1HfI5Go9smgRaxdIOXA6GUxwqNlYqzEr1Q27ujkG+orw9uXyx
lABjTYsvcmrcz066a2LC4Pi1IZn26MkyheFi6zQ6LCRBhAUeP5zzk97Y7vI2IVbZ
/6D8+Wb4+RTA8+btm/VPE/pOP5TYcIphWfYo0GoiHWuhe3FjganoG0sZcS9FtoGq
f7ObsyD6mvziv3+EIC+LNTsRUt9ECM0cWFxYytZWKHDxdlxY3/Hzfg2XymQ/md8D
GUEGKlZKgBrPiXRgd85qpv3kkKYc8tbwRLKB56EL6ZHpt10swIICXhf1NrQXdKJu
gctZ/bT4vxTbdlcn9kJ/iHBjH1MfCwPfIVq6obDV0501g0i/csNAsZ0UrnxOgxaM
Xo3BpcSl+1mUI1bXEPvmwpX88XtfeTAcebBkFIieDERwfvlqui5ObCvC7lsRVvog
UxohWouAX3198TcJ3kwJ6Lg7j7ZunPGwN2b//ElByv9nRcmnKucVJ6MCS1J81qZt
65pOBxAqPAcIb3PGTReoI1cxlP5rRWdeb72LB/g0a2jwYQB1a0vte63y0xnoAy0J
/zitjJmfLGBWdOQDIFWlJsQQ86pBPAROoxEtP+kVdvr2YWXHmcKy0x3FDgw9kFIM
o6rNbDP1vCG619sUdHOjYacggSSInTh1E0l5ihIfjADhdb0U5yqDn1t4a/dkQ1Yc
gZtNGVODL6RqGO+c2kF2rQygn+76KWSCRK3+fca5noxyca6ywzIQKU+RITpe3pB+
jGPthoYJCoFxH5IgeQtBquDOhINgbXcv7yM6ukgR3tf/Ng9yTjUcs/N6xNVNF77L
4trTlMfctPna+13cYMXNTwq5yIofCeXgIOyFNxXTBIsOIbn+hZYj0yHaE0+ITJrd
/rVGJAux33QjRLm8kC+Tsccf1l7SHJnFYvcxCK4VhNxRjsfz8UUITxPDDTXv7j3h
WYl2biwYf9pR8JSAPLPH8JaM5c3ph3wOLakSRkcHhLFR83Y6x27UbQ1RaSBmJH4M
TDE2YGZXKN4GI6nbTjYXdxG/kOEOoKrzctjXhACs3iGkpKkOTwENUHK958ZLo6Sj
meTe3dPDicE2Xggv1TP0zkSUHY9LIUECYwpxBdhzoPRY4VrFngKmRgSQwcqroq6/
DXe6k7OEuslpF3Soom8TGjWcuvD+xdSGTYY/Z6oQQl7fc1ghGHG/GWEA3GvCUt+o
yW+PlQ7rwubklR/ycRD/YfzQf+nb/bcrlF2c8vw/L3n2YrWG7FnUX3yn6Pyg1hwB
PSPJLVdxwz1OkLxljuuQPcshu5koaIWuPSplWF6hKanUyuDlGv7eSAGWD6aT8WN/
ccd2DHLkjQqmMfeZycmJys01ihrq4HipGVVtIqLRmoDYkFUKsqNL90dtC3WmxnwF
5euVsaupQQP6JVtskfo+bGks02VJ16l7O4BkKcsVuwXu9I2XyAjww50S8YdVFR2g
wfUG8pfiIAgqmZO6sXRuRDNsUCuyat9FaztsBu5L+Ew9t0MW9orDGy4jKqMlAd6x
CGqkaA4CcR5TdtfJ+6zu1sCMhVTUACkFACD7ymNq8fHIXYf3knq/9yw0McxxE9nQ
tthq/m+UvxWYjBpiJO71lU2WgK5qVuJbgdjLmfsLYF3u1BPlJWLu2cDqpqddos4e
zxU7rs8nmk7Yiba0a50Gb49Sde//NoRvZTpTT2JwauEGHUdYG3XgAfdl//HW74yW
j67Y/rGbSaMUYmoLeV8+Jj77OYgne4ihkMKblBQNPaYL+LVKc5dXzOXVF7A/DN4m
bHq8hlc24yy8H5RbWXn4Iie/eUQZVzQXuAeHhFpYKEBzP6UjoNvY/h6mhk43iisY
MRzoUf5Cqr82HJeiSYgfROtBifcKvgv1b4GLozU5+6AS8agDnIzS5668fp2GB/Vf
2wct9/iS8l9RD5p9jS4wOxUE4bG6ewhrCcJnjojgdrUH4/9dgOITFo7K55U6mAA3
x/E6rezGrGKHeCXof4t+qUEfaYH2/PmzEELd0C25voW/l0EPficX+BQaoXMmEMoJ
LXiWdhH1hLHnj2QDkjB+DKNew1y37NFNP/PGB4m5b7EUmNBVIqWhBPpGa06tEjp7
J4B6wboqguzpTc6UdxT54ggx4UDfXSlZpHnn1FSdoIwUWW6UlEZ3KCc5MPaYoY3j
F1bdlKBxoxTf9Xb+lBUXXRWRDN72+gF7uvRWLf6l/Lxs8mG/cA4dszTahRfnVFQW
7q/q/mUZn33Oz5txRiSdVb/KopfXjRc94jfAd7xLQjlfoYcfLXQZfbIeza/VHrI8
qm/fTtUIS3MM8JjtBlPfFshxRCCKQZ8r/7Df9hAOKySGuWrSt0B5507ka7bx0pr1
JZvXs2llm0pe/BZ5YOcF0prX+xyZ/Zzo6YIBGdgYxGe8foWAoLkBxJ3fwXJV01Ao
L3hSkv3JD7IBhP1AVZdHjZSqZEIVKPISypP9hsRo0K2dbVYzSP0ioAbY5sCY5WM0
vcETq9i6cwiaI581gP5JibDICRI6vMSUyT68E/otNt3k0RE0Xr3q9sWCCBTETMl7
BoJ7ysMjllacYD1pxpFowaVstwC6UsYK4u2sZag26wFYJuGU4o4gdj+rWw8cE6L+
xBKTXJYtILfNPXqGW5RBzPJjiZHsYrs+9tTYdbPW/4IqUX6LBySF4di172KQXlXd
IAtMCURuSPjSwGsEWd7xI5c3UgD55aZDlbuUmxSzpBmBVsKzQCS6AW4qyaRVFc0P
pPyUsPmZ3u7WPtmWvFEPJXrPja9S8RNGyjtVULEHhhoYMwk0ceRKQaobNhnaHK7/
XpMvPLsClHvnm1/Kbyc9BCahnC3439Jyrby0vavzca/y67iJcoEcw7onBNi/o/fR
XOOmK/2wiQl1bqxCkfjL5E6m4TrSqZGOUnqgHmIGh9jbfKYVeEBzzLXYNp/e1kbP
96PRH4+6zoTDWjuMmVL7Wxset1Hggt+nORIwmuIVa9WzSXEsJyqcbEU4jNyAhZq1
a8Jj4I/kP7k2CIDpypFO26qXUChz9eXlKfz/nt/RTbaRs4+fkA05bTfNd/ZH+dS6
xEugWX2JMrnMZ07HX9Qr/mk+1OA6O6D+GrlF7q9xwAh6nCtFsfG/OD9at4C+5dCo
6OHJgvnaRVJyO1cd9LUcGMvGt/kEY6NDHWR5E/KZD9AU7KxHxCgy5D4eY5eTee6h
GaU3ODERATXFW4rrzZ9Gg3i8qXCjVOHKX/el0soqkDOkBAPvfekiCW6gj5JrSbIa
a01Qf3HDzSS29ZnRRvEaTEjHcQS+HN67Ul1Otum46dKQnDHxa1tgG7XwHonIPe9s
zJXzGCsp0xDHCLtomVskQe6CssW3tRQ1kT1II8Ng4dQXWpPDocaNRz/xGu/PQ/El
dKyB9gHpX/TYuaAcrwf51hyMjYuxMqiSCmJvqQejp+1A2bdk2nXzmz3JLwJFKLu+
UjwC9Oo1Sn2cB3abIxOVfXJcN55dIJlRdLFlXERScD9Y9IgjzDRcG6fU3X70xcto
AtFZ+VdRcojcMwcvHkTRBywOy4b6dm0eG0cPm2E7L6tvsvDUIOxag68Ig76q0pNO
RDKHWq5ZkLQGge6TRS4ZyF0tjAx7jWwwFZ+9n5q0sqj7CjYocb28Zqp34WJalcfn
pRPBoEyMhqvIiStxQQ2527edFgXjw98JBm2h6SGR8zqFTxNbbDDIRZ7zSPRb/iy5
uebHtkGkxQK4ilDZ2g3k2FajNsHGh17Gz9+gBAePl9EfAx76G/aPGkvJa182rrYU
DQ8u3DxTiYFyPMeTQd7+ddpgVsMNQAh5tQV4W2V1T0Z1EGMazSsRmCD3Z62f44ls
wji6fwI1FwgynnZgsA9asHeyG9MPOt42hLJi36pbWJAPX+kE9rjQeOcXO6SgiL/I
kkEbMnqudgq1tzR/LI5MabvKRJWA10lilWToL2Dw4gNB5Owu9KHJz9YzC+wwhlU3
I0KfQZdAQJzCEyfiJ2mTRWDnwnXoTg0rMqOJrIDy7SvMftR9wQxULSKMC41mVNYK
dpL4N7FH478PPc4mwY9/J4sx+WtdZOeZ/WLLQVO2FBwVLOGXLrSyrtZZH/6veOPg
ECZTtTIK8ytHotT0wmV3azYQ8hrV4yHHR1L20vQRzftRgaW7fKHe53LdSgWu2Ixs
92RKlAfUEaTns2D3lYL3pH5LodIfwVfH+bt3rm97OfhmuAmgTlY5yJQASdDiNKMY
BgGBpHPSdQpIVbLdQhz3Julw/EWj9SKcXZgTHoFROSmsmFX7Hu7ZVu5PveDx0eSy
/rKEoo+gQ2nqb+cePJyc8tAF+rQddCmuZWJF2Iyv/qA1Za9F+O49k2lqZQsl0iG9
peiox2ctQUeI+jApq6gSOigl/eOEO7z+sAkllTNVQwqNO5R5fMOJeog1cDjQ3WRm
egpr8x60yfg6ybVS9m8hqW9T9bs42URqN8HPB7sHCjo5wyv+KBEmVn7gCA+WmK+J
8YDkEVCpg/D8E+DBL5ivtM2kLFIJNadgzaCw7yhq0gDG3kTAwF8TozY0aM7hbjfj
+Gtj7U0S75aWAyBE53m0E/JikzLVKf8JZjdZcXCMFNS3pIS1grGD0dtGLMCC8nem
Km/xeHgHDTnbw578b9WheY9VOjUB0Q7u/qgVQtLMjoglBAB4g87go1LJFvOh8LON
i0ARQaQEQDit4Vewf9BucZcQ1W/9oMgqVULIHrJTT4aJ2td5xK2G/MJPhfknYuta
SptBNa1pUFeDVy+LJJzgxXY2986pvsfGDKgp7L+9HpM4Xpzj4uTqJXo5F390sDRX
zxhd7FtFfXvLEP7kldyNq36Zsx2bdgiKFkGuWNkyVu5/rG8lhQnT8R4gczN6qhhH
KO1nyUW0tTR35Dy7f8G26WlFI5rP/y7j981QnLlY9B6qbnYwyFhLwzOxZdNy63wN
WJvR3fpgBAPnvYDKc1IGfsrlq3GmqLwuj3HBfxTi7nm0vYfSBrOMu9JbYJUwfhJf
rkdV7Ka5FhxXTpE8m8FlgM+9hqRi3jdgkvioERT6os5BBeUBc8Ux+fPTQiZ2RAS6
45bk6hT+QHpmC+fr+DfanusXmhQlNwDco9tOy6Of9VTmDdw/E5mg8owU9SK120jN
U1jFjayxz9esVIrwPzqzcbMmSWyQ/I8pz8KVSRRvpJGiDsY5jjxmdnVcpqBSyXS8
aPaeGxjA+CNRydNv8/6quqCAabakD6qCNQESnoOtGCEz/axUPUl2LZMSg4xX2VLe
CjyzDwyPs2kmeguFDR14cypxisdpGDgeX/0h+5X1x42uEhJWC5Kt8tjGreTu5r5o
oswzl2CzgBeF3N7sZF/pObsubuPTO6n0wBX0tGT8NKrGSiFHLxVMwnEDUilFv2oE
336KmOq9PYHr1C98SGlAAqmvZWYCvPOFcH8BjAaS4iIL9yKU3jC0pu/hclbPdMap
1ccfmeC55ZxFuWCNzBrTlLqhQZVoksH2Pd3VuDGz0Fz9HzdcYXAqdhUJA+DifRJJ
rPpthuMmHNahGzW2RuUe3BGckGtZUfmUjwg3w6PE05DwDBS8gZTrsVhbbOVXVZhh
JjhvDI+4QMsimcqRNlgmdWnBbFF3XXbRrC47HJZsPTAtPBDXU9d7xRDawVwTzv28
coKNKkdk4EXO4RixVd/Fu4qZMCzncbrdPUfzWl0wicpnCK5gW4HgtnzFeG0zcMLh
Jh68dHyj41XUdT8zBg68kMMBBVfRZ4SwDVfr7MYS8RKsfoo49at4/a1ypcOdsUFx
qx1Huy1Oa1KmMSIudQbQ1U83gpEpsKEymQaPE25inCbP03DddhWfxZnhTa7CWTBJ
uVzA6/2FqfOvpN8RSZfMYo5b49IwMxTuu4NsSfCQqYD1FvcCXdJOndF+GsUeGknP
ajNO4zJSCfMm9k1AdDfAE6Ggs0fPq+lirXnNYcOQTeRvs48BxNan/l7ZRfE4MA/Y
gUS7DaR/DYTrugJuiqWB/o878BFCVB3jtcRbt8eLhmGD6fRW2wydEt9ZQfLhttwH
bfWppYGecYs1qtLt572QUwAipbtHD95K66d7jwdFWTSo0flE8n5YTCKPz8D5ULxT
SoYJhiS3jzV0p/QbyFaePG5LIQPECL5jNcr2FhKi8qCG3sgK6phWZ/ht9ljhZrtj
cMf94wIscbHngWFjwUoa1RbKRvmTxEIxwVyfHMYOp1l2Bx3Y2rnynhAKrIEFqnpw
wBbWCiR4WZzyEzZvPsILaKbJfwDokgQCnqmjgy9GuSku07Z+JL3XVGMijYN2F/+X
0cnDXK8AFO1XnzAz03tua9ZWPOYpHyGlt4Kgl7ojAxkcd6+nbUxFGXGGIoNZ1/Cy
Upbm3hDaNkFKJMcMEX6QZd51aqR+itVFELHqtrtfhgh3kVZ2SJE8TMXEOr8DA4qO
yIPej8aVKNQEifJEUahmsjCECYWcrDCvVyBpMlZbRJIAIKo2AXbpvYkIkciDkvEh
6Vqga3rMKu7eMwAH9uuVv0EuBZW8ZxC4Z3LNMCuxkX+bUet/WeZrSCft4/K6Wakn
Hn3KuPcRow+85t9djs9a4YSlz8ES/N7boPT9PS/z1ojx8/gBdgTjCsdeF1vOtrm0
BuItRBpDeCb0Q7TLBglUkxpoHqU9NEJR45YVtG0U7AdMetn3cLVsL6vpMqlFCF/4
gDR0Ycax6yLBOKQhtDqFNgFpFA7+dXRyXl4mNa9vD678DKWo0lrcqUmyRPlOYPKk
lkCKspd4jHmsXxhI1hiBLuaBP/x7fnUDsZoUk0bzpwkcVn3FM2C4lF5k5YNd1RDm
HtDH2SwZjIW602EpAG08z2v8CvFq/54aBNlCSvasytJhfB9v7EdErupTdI4sJjO9
ZQPZnJfmpnTK8ANChurSn3TpRENndROp6PzpNhjRV/LOCACljw70nT+98pLSaKSK
1RSP2H81tZRWW8uhi6gV6IC2n828mASDb9QD6072cTr7iteww1EIASU8ilbWh68N
F48q9cq3fzzAjncD9etAlRtDciq4rvGfNf1JIFXLpaf8Hgp6pl20HgWIa+dAqmMe
wMdZYPbJsmbwV+oAK8WLOx2WSbbYOUht15+PDSrGxgXyyUFDJlVUO1VyljZeZOhQ
ygCwyqV93TO849IN+jxHtlylON7IK4mHr6ZDD8LCE0TBPoPAE+DNjWzRyKJZZ53q
sRrAB6TRYN2FJ6uvhvuAnlVN+vWV+8ADntiSpLgIpeJFRACvbH1X9e56dD6QgGpY
hroMk9avPgCAwfMg4X5Vhvv/HZJN3Li4F6Bak6rWbsd59BnS1FyFodg9AQTt/ogx
ywO//McysCgPpOE54ixz0v/sgvvN9UNAwElDTPRfh3YmUPMaCKiWyvp9ko1t072n
PaxfIx8lKIEBO6Z2PEXrXIWGLI4yuH2Ea//MdtREDr8iAZbzCoL4q0iHXC+tumBa
fzPfo9cyEWSkG5Q7ueb1ws1KxSSEcWDH1Q9asv2eRq809dRSF0YG83p/4nLjeHql
C+3qWtAu1taRfvbH+aP1hJEfRsveduE004I6xXUbDXGEgzbu1QuRwgOMMK47CwwM
WrQtm6ArHV5tVlJ2deWq1dtNiVvIzU6y9O1WlMbbuyy+m5rknbYen7ku2HbLJbAV
cg65oJOup2ondPRIuMocUktSFqa/hN3IRkuU2TNL7hChJB7puI4DqJC0ad2rd8EB
jFbrzUsmz9NVJumLyp1bclQDUP6naqXahl1H0zGyR8mkS4TYRJp2kyg4UOjYPr8o
rNeat68O3Eay8vfitOom/g4ZKMb+EuL/1xzs+oQw45OzpSTOlk0ZcfzHLY3ckAaC
2YlbOAa9GeOb9WzWU2ipsdYySlVajbJi16Nb2tQ3qPHvYgLQ5DhHCH96Us+Vfpgx
DfX+svjpV1xM/HpeG2JMsFGWqgFtN2w8GKQmAl2qQ+z5Y7lPRboANsewOQODzqfd
NrLDT9lk50SGSLf5QiROYHFFIrOUMxrTxerPalj6eXsepmTN4WrwKS+N03gb0CaJ
OFuCO1dzmUMBaOQmvMLsdnOyObp8k82wRE3Ej7g+wwotbzIAey8NT8hlt0ue2EjM
nDgnalSa7W3PRv4z5hsp69d/Ajmt1PVgA985dxIEMv1rur1KaAkfeiqC0AIgqcos
n/FAWarhtorgQoMZkPEW47wB62lC4bFzqu7BlXzio7lusXIzpGrG2bWx8/dASHAF
NSwDjyL2yUi1mpJhQ+VuNf9g/nf8oBPdp+0/Ru9nza+cgeqwJvMza3IBqsnm+cDe
hZ5sYPguKkGSQlR8SaATouy+h7zMKXXCsGBxTocp4nMBxaTv2fIjAOidjoX/kJIv
/YTCcXYGCUVQFDEZvhMqJ6iMJZ/XfgS+bne0tG+e7FrQxwu9QtSa06ITWGvUvYHr
pIx/wfTQ4e+UV+gJRBQmtuMSphqsTdOQP6vI6qi9P5hN38GLobPtqMDCQlRAsTL0
MDaC8Hx3j7xEuHGfO7Gfh3uaEwdKnaWxuNUs+VGSuvMQLDpl6HYR/H3UuJFfPo5E
MhdEjnUK8mIuzVVYBZfydxw/K7YcPG0JBD0PSiCuxpNnEH0/n96MV1/rbql0fYbF
EIjmtOK68vRgy+0VbGZ7sOjHKW0MESVzJVFYt0AFQEFqI6oqJiQntsCGiwtQ8K9O
5DwPJWVxWuonQe8YLFEQqzQ81uIn7KMt63DSxaTAdJH7vzTGW7KPejK333RmIde2
NgGhME5GAnl4Pex+CeZSY0FwKowkvtdj92FTPAw/cKSYEpDI+3DCPyKO57tz5WbL
grJQacQrA3phdXLPUIwrXwUhXQ95HVw1EpL7uRyG7dvIxrOfLbLt5rHyBTzJkwka
kmzNpIa7ADed83JV0KJ8Nd7YFmX9UvePSSv7YWwnlLefnQni34+1ZFQeXNW4dumb
snAJzQf8tvsHJG408B7j3M801/sIpKQ+/izyv8gDt6KDQthB1oARFlrukar7CRvq
gr5B7xQWp2yMU7BtMd7iOS9jRrBxfMK5lFXqLbhcOT1flSTj/y2G8w7cERJcAhKR
fZRl2/ftxOzq8ixiLO5G/PQRbaVRrDm0jd/EcFD+HJ/DulzeURY5nvP/KRc4cdQn
Q47TeFOno4t/7NBHcRFAhoMAzRMaQgCVM01s9gL/ouI12z3w7BLeXjT5FNroehfo
eaRuTT6dvSKM4MTY2dNOzTaSzl03sv/HHarwvJ9okwKljDaxvsdk1JEdQRjMz4yl
RglMSx4sHr05YK8xC0eCTc51j2JJtx8PtCZMQpGi9yDKtspDbFxpJpq4ofP08grW
KL4bU8mxn793Oqq2McA4TW8/KjveltnvGxRpZTr4Xnr1N8MbPLDlsGpER/a22y09
UWsh0TmFJkSs6IG+dtrEKlM+Wt/PfPRRwwmYd/oy6yQafbe4e6FPhhaf2kW0Ka6O
9dGtKAHadsDdsIGJl8BqWa1cTpXnDakGiNgf/61lfYoenKpec4JXeHcq0vs+mFuA
fPJj43ywnZzELgNr/jCcdgcmEBHHdPMlOlAzE6TcAxLJSEMax32uskrCtnP9bPRl
gC+/9fTA1goOYc8lZjzuA8vaiNg3BrSrMoH/B4HHl9RvuovttugpPZsJccspES+g
AjN5G7fk/zzb8G4+gDpZvFfaQoaWUUiQECLfGpRFtpwd1iRJgH9HwLICD7ys/z5A
NM382fekHzKGL5Cd9t2/fBBSNyAXuUGhg3sON1DWQwkCmxVEoWgWoaOaia9DJTpm
0hAZkIdyKLhBrgnuuL3Zf4QwMRv6cPUmE7qd2CVbjbg7sb5EuMRgzFjCI9xY49qD
CIrXh39Eex3n9jgG7e4sZA+nLwIs23FP6xSWjTE60Yft18//Nu8ZHqZe6xJxebU3
+ZvxYcXFg9TyPSIQGiChiin/rRYm8SZch3tU3GsY4ctsUP1atF7N0RNDOtFGMGCy
kp6CsKZLDsx1BWtpJ9itLRP9ri37i6wVSXJWJL6GUg6Tsen/AxbCzOdf1w7iV6tq
OMnxWc9cDOoqRsgXXGrQB3bXlVNWxz6BYzVAd1nonNJQPGh89SpFp+zWlT6RXgrl
Je/M/6KJMjZ3OY/sCC+bxpOFxM3srpgVKNOVVyZ0c8gqG5IznogNftdEKFDstIDW
kTDboyq6703gVy3NZ0e5FiqQ2ITGvngb+ysX/QfEm3pYhNQXF+mf/53w3gLS+C6u
OTLJ1xvqJ6mC1NioG2YtckpEaaVFmKuhFqnSAU4ixPkjc0N0jrxsAItiMR05kqtX
A8WYHuijnf4Qr90CrleSilV8IBdANv6zdYI46HtvW1Ly+sO8nUYSbAh+JxxtB4nD
VDN3kHXKZHYCrkLYCKWlThdQxAWHkGidUm/dKlzinAWxZHB6/Vayl1vLVX+6BC7n
nnsnRs+Q3ICt2rxHO3ERVBzVuya8j4kPZOaWwe9Fq7tQaqPwC1hFEyuNeygZXx6r
AefrA/K3zJwycNiBvcJRUQVHis6s5nM2zd8AUFxcATk7BGxw0Lz6Qt/JEuyqYud2
XHPF+kPVfTiNS1WrlgAJlpj9yxb11juqvSVWtISnql1h305C0HkKjlfZE/JNngPn
rR4EsI70KuOIw1hHbSVs7B520T3tyQQtrrrMiGi4cZoHZ0TxKCHoZKToF3ljVL2s
NTYr5/vjamFjhghgsnvCg5QfL8QisekTJ7U1XmAhvSEy7ce43Je3ity7hPB6qf36
u53AqgrjMxY9dGhHrP0d0dr7WhVwvvQIQx9RxC4AhOsJH+pON3hNGBojzdyiybOL
AeE+qkw8HgDxuMH/nWFw0BbwKuOss+zEKaEUQ7WqeWlq47C7N/azCipCjf9kR2FH
MsJZJNWwo7l28wMUEKunPXC3QykfVNRqaXcKO0yzGg2YVDTja5sE2e40fyaXgqkz
8+PH7YW5szOF8EdG9BFz7ah9npEk2dB1WQ/TTl1VnRuGw56NX62hy2gm8RlZa0lU
qiGtrqhMKhsbdKuaQczXFwKtMssexMXdlSVzrzwfjIV0b3GSuvAyg7mqKumjXG6L
cLL+1YGnRE3KXMqnnxJpCW9zZlB80idUw4q238u3OXSI23R/pl2lg0/uC7G9iiCd
4uie/a/N2Knl1s0QgKqjVjacw882OT/EWYGzB8d4T4L0sdgTu407jDUK9MOzp73l
0WxbuhbYZ5TitP3AmRG0LbVPgcELivf3Y+gPTteVjsE3+jZHNkYDXIEC0Rydl69k
NTj/y/ugi5UYiDFPWvkFUQTqlFwjdo5mURL/+Lk2XKQ+gpYFSQS1fjYCKrMaxrXb
4FNdxjZRC7+qV2mf/twNz2Z2o1tuT9fbIp2mfuuyjjaPLgBrC4fGL1BD1tekhAvH
diVPhpLY/r3Pm+jODIMFidH8bmwEeF5e+7s0jG0MQOpGSqlM6Jfik4mS9dt95iPu
8PFXVef0Myc5wt8LbRr3jJJetoe/Fylern/bw5UD/bRzz2TQJlC4TPUw3bBmHP+e
oRyc4Z665CKp9sH5TWdh0uLAyFD7OUOEVQ9NeY9xzkb6fxat1gS/lsljj079tS0R
O17CXM/ZoPlDvafreARAE4nDsJNOnzlor+OXxKeNQflRO1YMWqIQ3pv7VX+XbL8w
EX77Gc/VafZIcIBMr3Cb7GKL7qggLtzW1rI5+Vu2K5pmfWrEydhsmxOrw3PghQRm
z++rdoObxSsd7L8TX+VrncVHzmXr2ipmeLMhtPaxJfYu529Z3DeX7XbLsotGgh16
WXZk3+N5BslJtQDpTVP9cvX5NTZU64Pgzw73cIrFjjjrtqCcZQL72x7pQxRfpg+9
MUljU+dlRDRotXboVymQSnIthVztEnq8+llNC8WfXj2RxjZj1Yn5gFaHjB8yv0bT
4EzYNQC7rkA6kllKa3rFlQA8nf2KN3bHNPp52qau5+CsPuO/BOzTqMtse2SvWeCq
LZA01xjgGqKqZ5AHCPQ/6dajYOeQhsgMpMG39VlH20Rn26FAxHXjQfHd/GkBDvCG
l2kn5uKRxlV2JuUCiGrjwZCjzy/sLUd5IsbUJjKojmUo62olhlXNXqrUTBHsPHOI
+yhXpEeVQ6Te5saD1edZeLClsGWqhXbUV2S+RnhGbqnmQtnPFUrRdkgApHqgfc5u
E8NDJu42vsL5W7UPx+Hha7yBdaOKInmdCu5SbaPaKD5QNjPxjnH9zudSGakqp56j
OZZjDk+TTpicj8/gSF+NDwvsxtkHk3AhiNZy9XFi0RWJG30SUK8nzbFBVhBoCMDs
WeIlGMNyaRo1lGI0p9oXWCFLlSqFKg+ZDoExrY7LyXyNyhkVIwgvWD517P1QhQoE
j43ZGsVU+hjtzeOuy7RnCwH/PeFTJqjbYEgA+vuL5+LhllBjz3+AIHouzNfgT3el
iVPMWhIaUQyaJORuto0NG/f0ya4pFzW8ofSf3CEQu2WkxpBAUdA4+CObtZtrHT3B
ZLn3x51ALw7/0HdUOFvr0v1msVqJS7my6v3TMnn1L8gWRjfIl59CgONWmemqN5/a
lEQQ95pMBJa23Z17RvGn/JV2v2hmFmlW8w/iW52zkzpSkKZND84Cbcd6dS2L6oWk
z0KeOMx97J8gC/1FiPmNpTk5LKq2HOZ9x2fwuJrsnuS5Zm1g+LU/Fs/t4KPyWJim
AYBHz0YyCZPskupEaaFHHWrnhA0ubcei64BJ95P7YmK22ifFPSdkxNEmw1EP4AUX
RnEIJ5+Jp7S3N7HKSHkcVsFtVAJdqeghULyF5RRGMNR0GRyX838Ebs1Nw7ueKbXr
JKxgvKl5969DD1nJcy+fRwjf/8U8pfO/LXRFUFuF/2HeZUJTMK7dKCd0NXfWoZ1u
itTY2F6Elwbufci8nAHngLEYo0WErAKzfvKJn77D8/rk8jKXVJYQgIegfYiJBQCT
DfYpAwlOAUJl3IzVWXznxtiwbUaz5bfxG0fIaDR+hMXG9AK2GKdMBvjna1pHIQlr
XA4iYcBCNJiSLwwGmZId3bg3rY5CeWBh9cJP+bqMxD/VjzYeoUU29O3Gl4I7nJVT
N4r0lbuV0dwH5LWXcoIYOgMbKRuu29liFFbRxLGhjako42RT7bS9IUZJBI9QWwr3
Kw/bzsz4BGhodepTeBc9b/YN1qsNwztelPBw9kflf8dQ8oSadidaF+aCCWZFXSbw
Jl0JFvG8uHUseT4u+Xb41Uy2+q4q6vs3PP+nYAtowgGpR3IMMunLlfP2LmZ80pYM
ed8cOJVFSY4Ksswd2DkmGGzjzNoQvG3JqFu1Zly3Mz3OqddhaBZK2onBhclgfhHM
/lDwS6D38ZjEGX6PmpgOCLyRczfSRDR4gWlT3nFJJGavKT7PvjFMUoSRaJxEvxDi
69YS6WyYB7YbY3n5E7al5Vsacjw2oRcbAHGNCu34rg9SXE8uMpstAVEfNv1MXA56
wRgv+EttYxmlY6Glfh2h0zbsDAOwm1Ghb/k6JjcTOZg5tovvV0dxP57i4PSWSZHI
5XABfPNXm19dIoXAjdyL1N6xnTT54RquI/YqJ5+t2O62W8cbFCh+bn2OhcKAtwIm
AJPLX0vRPLUlVMqM9/8yPN5ioa2cVZl6UvDO3Y3DbLR/u0NA0PaXktBGzinh1Mca
+OrhjNNtT/Zh8nBh8scsub9jSmgoRV5bIIJVIpsovmC47afHzraLZFCVkmPacZWH
CeXddJDH86XWRqxmOpRXFxTSx5b0og31IGyqQvtREnIcw7vg4LM2Kt2WF6rPLJ1+
3BHw7MwzbeHkLLweStTlugGGQ7t+XyhYVmfmK/YEi79kIaNfhWHZGb7pCHTtAB4m
hTgmyTCDG6/ibJ4WwaWkBWrhQkBkm8IXpkyanklH/RG4bRfriieEf/DPEAfnf31h
wWWU6S1mao+rEdDFGqgMBBSRdZGL9mXsr5830qlFZ2h8mkF12BECeSovrEkswL5T
NfQdUJb+SZ3jMPxTkPQ81FRqEv1a1U4VVORI4+Sd7twwsfGiz91vIttrd9h5CHKr
+4bVn2+4R4YkJmX52UEy/MAs1Fx2HXfBtlXwPfF8V/UQ6c4kxDKzNp++iIerTeSp
K73UZQ4t0xomt2+t66o606qSPaEWLc/7ejgc89/oBxXTlPxDa3kLje1F6d9cTlch
cPiuPlLR6FbD9LmXqsd2AAIR7w4h0oaL+M0y8jKHfElSFqG9WjiPWguPwfDc4Kzx
2NUHS3Dz1JJIWoW+YbYYMXCNQNaxW/dcGWhna+ZFB7JQBNgNut4kINxfqFTmg/ej
gZ9PVd7YKlZ+T/YP1BxsvkNUom2xLJBivIx35+wXj9HrUppZmWS9p3aNpGTcCzuz
lN213kKoPsZVgyPlbJNGRiq1TQf4RRgRanQLnSl3CbY1TiovkR3cj2TR7PRm8K9t
2ON3RMv6XaipTLqcXVeu2X1PiMmIXa/NHrpvH/0YK0TiS3pwgEWKQQWciqnN0wMA
CNw+rtH83oEi+RZNklGA8NQMnrXH93hhG5T/o9MeGTaURiHTsj9gt4qtVVgAiNto
ddJYF2MlrRqBPFGcnkRrBtHsK7nf30Eqz/pxrIjEqiegA3woEO4xN4sjHNFOSTsT
WM7sSEEQYHdOyr6Mjfv29ErmzKQCDc9h9wW9G6Pg6/XqJBTVGfudEo1sx0Qsavfd
ivsrPt3Daw2xggXv/s9f/HfOWH5mdIUF26afP/cWSW30vOHCvp5rgIDEcz+8SlL2
qGt602DE2Ju4m2TJUR2AQgqyoWD5Y0lsOOcXRA/0oVfMkYZiIKHrcET6LJwpELY2
EcEYeIEI5FzRVJbceVeREH6EBLS8U9fF2iXBaNY0i1uPJJIp666CIVGIB8sk46WI
7XIIRoiSWMixsNakkCTJSHp0timmaWmNNCpAkfKrbjgEyyKsW3HLz75bm8uGyx5u
UxNZ0/DRPFs1dUdgFEmOOKH45z+0gZGVUmsP1dWQz35a6vxYLrBBqxdWBc/MlsZN
HvelUXfVoAIH33vr8T8574uO2/W26j+b1Wrl8GqRKbXEmJrhAEFeosN0RLxNuDXq
69u6+E0gfNCOhzoV0jKTwuGijyscdO3QiKRlTLRPqo7en0LDdLyTmoJmNDxXzt8O
BG+ZECzLS0l9o9WrMqFVg4nl6lBZDgf/tEs34caylB8I0hDL7vAuOcIU6Yoe8uun
x5jrIh2lep90PFGcpfpcRnJsHd7KtTGAU+4W/SGWHkuQ6e9bEUtK+MB9nH2Cbn62
83dunW0ugu3ZmcbRZ8DGDenRM2Q5cm8YuYcNfzt4Rq2YNtMzGEdISjIaOWIDt/lD
YICV+jTEq5NqHMqjMqKKR4CULQRAFHG6f8lBh9DzDt60gCBXLhaLaF8lHK02nvVD
1MJhZcd+VDIBIAp7YYb7pB5p5taXI4X1mVKsR59ShkwZK90nLRbD3UeAikUijNUC
2ECI6/fuWgaLxxiBu2PZV71ShV7aje8RCTqQ6cNsGFU/uLS//jCAoWxRfoCgN2vn
dwD89nraRbaHCy+F3YzJUuNKopuNj0ns/C9D49FvVKTktZEistLlmKgPZbkG//y5
U0Y8UuyaA/k3TLqqbM0x09DXHiwhtMPXWAcDT4bfoqtXBk5HmsFYZpZlZTEqNUBs
USpjx7/1U1eDs7SgKXjMvW9YhUcruVWVk/TTo0GB4KjgG2pCzYmedAoGcZoxTszO
fLY6iLOSqbL9IvaCbmGmqI2va074V05SrzbCpEsxBkGPvgjzRGUHro3oyEq7476g
2YkMEoM8CiyXmTlPhERghHEJa//eALRHWULJBKpQ9HNYrW42U0zlWnJuARva1xWT
RYuqM3v/T2c0fRTpPXcSSS+XufBBbv9FtbaHwpVLqtZNGYXK5aiEyulO2c6KNc+K
K3sE1jEM1jUZ1sZrivbCjRJKIDGGkio7RHBDINrM8ZPJNOpvG8TFEBywAALCsJeT
hSyhiekPZMzTJ6w5YcTTJbxyWYYE91QHy8tZKG4AcgKY4A8VR67Crr7gZDkQGlJm
g+3hE40C0fwzQpDp2NDvQwyhuF+GhrPWAKYyybLIqutrlnfs4rEVAfo9HX7BPBpP
3blRAENat90c2MPkddj+6R1VQBUKnuSGk28PP+NomcXV8l2q4rAb2PuyLlEc/MnQ
4i1LQaQu6fKyANz1GW7p7tCCiV1QhSnrZyhq7ht4em29d4pc78nAERiMY4OaWBjw
9PrC4nCyEPurP5LPxfS4NNBU7gg0e9LvIbe9AxjRNbTIDwPop7sGfk2pafWrQyYq
7unFnUBjgqu/m5zd6H+4M7hSRk8s002GE/dmbzucOG0z+lIHnqhZuyWL1i+yISi5
z2naoPiURF6gAK+R6kD2OwkjBcruNp9wjCeGlNsInBTKP72Zq0bLL89ndeh9c9jJ
tcmkKCmxkk79Oal334kkzppGmTa4MZ7PDje7Kh3tPI/WFF1K5nPV8LbGMGGYrilb
aHmCB1zGbrkz4U2vdwrFxWiz+6e/VifnyD145DnN+8JOa0q3q22+8DvrgUwcQm94
RKztgLznO9/X7gLLzKDzZE7h78Q1OkpZs9Ldo6vWozQb9YwD73KW9MBqGEyFNc2H
9G0qE/1ApC01zuN3hZO0vX1NOpbCoLWwXttHpym/O+AsK9WLeimEae/AxV+VLEk6
1NHfYfm49xabhAPr1M6eVEWSAkOfKvJ2auwhWY0fZB+HShfVNdstYUQ8//oayOsy
QbRuIkcioks9UJJUD64AMiVN1ZB8hCc+jWTeuaynRRutDXpXwr1Onrg3SESTpxCr
Z21/89fSUqDoxE8bWD37XbbwVEYY3wiMs9YEv8osilqdsuuXVnkFF/mkbb1k+d19
AElgNLcMYZ6IJ+7a7agaLznQWp35WSea2T1buC7L7nmfVeWEgm+RoaipriOQ6kNr
JY5H6uU+dtHnQ+VaqTYLclFiB/+WNsE1E9666vcSZJhQQmWVlzvxUDtsY2J2+SY/
If71FYlW8J8HF89nXL3po3HPyRADCFS1zeSI51jyIp8gdIGkQYACLQZmK6iQGj7P
5HantmNxumgxRJF5Ah9ZzV2xXIYNhp0r7qBSfZ1RQkjSD9oCCh2dc10jlOzuEGcO
1Z170Vm9Cr5HtJuwzYggTFnN0T2sdVzmpaNxdsWavPiq3skCtTqbpZy0xyGX7XhK
/2oosaJATSzOO/zzR6TzWlBqjQS4W/vG64eN5ZDXf4NUGU0GuZs+cn1E/ZljrA/E
qP2y32bVWeDJAzlGSciG6QnGBezbHRWYq+JPWkvIioAMbgVqVoHpjiAzm+rgbemz
9saUwlf9UehOItO/8w87BjhxTbJbb86xoRGPkINUEt1gciMTOM69okBhGHy3v/ce
KWX0RyjZm7nR6hz4TZLKlKxZMX+WLOXbZffl8r8d5E1CZtmAlfEeyXwJfO8F0vDG
559Uaz/3hcMaNvG0dWS/fWPmyYjmp6jYYW+j4Ah2VhTovpRxYvpnQsHmuPusRWv9
Ix24zDlxQbbKLTfB4jtQqA==
`pragma protect end_protected
