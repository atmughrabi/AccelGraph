// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
s0FFplQHaGv4iHKWO+J96e/qtjEKzwo68P+PNabisXXwwyDey8778YStswRi1lrt
zfb2ib4Y7InTTIh3sqKXjFBoMvC9DTlAhnXzxdBwtyFBuc+8pskdorln5qqNVLzN
E2tVp8oQNeXI3vzEtl0879bPx+bBJL4SQk2z3x0+7WI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28176)
Np5UU0Fus3eg3nFPBrAHOLJvF5b7dFzMvaO+E3rGlMlD+QsjTwGMOYpvXFjj+djK
7pkzUaFfBTSOaTetz0QPOgpEv/Y+Lkx6XCIwizQI7cZ41n2+z+WjUHDCR5TRpVZe
2quJ2WaOoBwhNknA4Q+D1lNxB24E9zXZ8ZKwIs8FqwdYYgt8bvBOZbSlYEZJOUlD
bHvRL1XnFO16gOyaKzh+Cg6fz7bhrKbc9G9F9Ya24Ex7lc1hwkatL3JIs5upheA3
Hj/w0Ry08rz+yL/wFz98AtBM3Ssnwrp04/1SN9xwqzT9w0Xpn2ax0fzDCj6JgVIc
TddhmJ8xqexfi75Vk3yOvG13rvnPzwrhdpcaTfw+ZtKCjmG3OZLFuyQrS1yY2m2I
JHw5SNFM2G3zrM+007RLRG9SM9SFsAekknX0ItmW1KVoi85yo9c7DhkQBrY+EulL
a4h8SifDZZUk1Vn+C8U6R/LWZYoauv23LPfm8sjdb8G1bZ3V3VrdzHmTbopuFWPX
Hew1OWVQP0lFwKo55Saaw3QwRSPUk4YhLRAlQI/lrguwEI402AdFKCisL2ad8ysx
kFN0tNOuAFmAO5E4jTsrJ+2Ry8akzIPLJaMXca2hl+8iWmT04MGzh/77VsGkLbFV
fBsX2SYXbwJ8eFSwOrp2hg/4AqV4HVZf08iV6oXZXc3kg0KyWw8DcEMrpTQ6bKXD
/nD+iOI4PxunFjw1pHh8KdJ6u5EZTrnAhWOoJH4CcI+6+hvVgzEFC4uqT7EJyht4
tyQEYNXjUUEx4ceIGjSDh0WE/Z6+HOYbafVHn12qfDSLlfY5fmBes6pX8cNx8MFF
+mTqhqGALe8is7wNJ9y3JdL08XrbWA62uvCQnB5Bx9gjYvtUzCn3GeyR9RWBTCrz
F2f7zwRML0t3HUq9k4QHjww9izJZ3V30L6RxF4DsedLsOS2oVF5ae6xLCGDguFAU
Vnevr2ZNmtSh3Fghu1rVdKIymW54Oh7DAR/idY26J14+v9uz8dClxx+v9Ps+fLMJ
21I44sOwg/G9o5qCje8IP9GvgYvufkFcj1kmuyZwOwjs2UzkvyC2L/948m6k7XgP
MNLO32x0Vc4mqV0jZCo+ZOH9JnrIQrCc79nxS5MBOHX7r31eZgbV2eNpAJoGM7eK
m1zRXn6oN6O0QmMdnLumhtytHXtJkf5RRLp5Qa8gBPwyQ+LvgN0i6/ObAW6rdP8d
IigYSxBfaN7Z4IaV65lgM+CA1MywyKAemJhWLSNr//2t3hN4vJ2QXGbBeyvr25rz
ckB1JC3+Z+vyqTiyOd6E+moKcmAT2vpg9uIMOqcIfObjbYzizElQyxYtoLliFugj
ps/2ed0shV1ErDKnFxyX1+Ea5qd9X/uVhdIXaEyCtatMxVzIbnJswrJ7p/HnXNke
n5zGg8E2EXDkLV3QRbmmXFGpae8/p2fAwiWv1qm6fhUpc6U+bC52olFITNb1T/i/
OGhmTBCD4e2pbK7L80tLW1zECr2uaCuAlCGnulw0Kw/K62M0xSS2rr8WRKFN/9C9
aojsIhOFprV/xa6mDPlkSu428Mw89PQQuMC0DiX5cwxZprXWi+NznP4GOWyLsJoR
Pt2vKz/zTcbnTgBm3fsXVsnYd/iyKGf0/377y/J8DNI0FhPbYJOhhyEqz4gA23KA
EaPmmH+ZOadik67VbIWicE0xLjIliz/GzjOyhFTbCHBidf0s5NbdXyVAGrJEcEBS
ua2tkTxT5ElIFDigo4ctg5NW+LbHF2LhCpvznB49OBXtuez4wndM5ie0yffSgqkQ
pL98tTPsXQV0MC556nWE4Axn9SrPaXTEo6UroLb55SU8nvl+88LXFnMR8sJkrTq2
j9GWUYdzOy9xKrTvVFC3c+kc1s0kkQ7vuNFJRABwL1QRF9f8d4LOqh2Yli1K0cjK
SJGcRI+h71TTaLcChAo+6pGr6zEOk6N8q/VOXLE3LQBh5GA6LEK5+UFjycxeA4hL
7LwqwBr9sT5+pUpkSKUW8WTjOUvAfgzOa1UY3tqgOQn4btEyKPoyIntar9zQmZAj
AxaHUGi5rY9i0c+NmTeV16A/BA2jfzAy5kl85BHe1FymfCzwWHjpiZT2SSOG7oB8
OpEhbZPJ4PwFn8DMZhmijUN5qyXmOXOBACLCSOMy34dXQ4vvGKCUL1UQ2QY1p37t
fof32aEJLHr267q3qsxehx901JtuBB0SnI7evRgicKfsRlQ4r/jr0QDGYcPruPeJ
yKHTAEJgkCgXK8bIdUgj3ZqA52jBAzXPkEkdYU2JeZHd7n7kxp8W2oYU0Nht3Fg2
QZ/JPsvOMSgFexfLMTQsN835Grrjm4/VY7gDZfi5JNJGT2U/SjEjdn34LT+uDYHd
rzGCTYe86wnIqJwqDS4g6wG7g/rWo6FPAmAbNTKhIC0lnkiq0/KzEDs1zbe/Pec0
jzfigspw19dkYPkzTA181y/LCJcDQOuQ7ASHiiNPd3E7+tJQDkXXI5ExEy9ixjHe
lT0Db18EHnSdxMJRHGhyS9clw0EKnlVmn3ZfRnwAaUhedpNsOASW1m1TwfOdRbsL
+rBAc9RSFjOD+8dUU3kphFT+G/H8556LF5+tcZWz8kzYb0lU1NwOY/rW3g8tY6U4
42iD0Aho5jXDoZQ86DUMJHqU7oYbJY4jAeTDTV2vfTXwOieb9aIl4KRLY639e6fl
sknMb73EcD132S93GHEHTCnAM7iRrus3D0f1MzA/MLeAa09yzta0wATGiUTNXQAh
kx2HtRegiZc2FaY4vVPFe/xMjwGMvvOW+UXJitGi0zJ/VFnnO6hfbNXotnduH7zN
YfMoH1QB66QKSQcouM2703p2a6J5dOg2uXOTSakEuLbDuSPpYSkLSLhj7vZLzPc8
7YJd49qiYMGegaio7/9uzQoa4hc4kt1jEus/jKXkWGWmy9paVbgEAwiqKOANLidB
nhXyy54KoQM65qm1Kg9E1W8gHa9KOCjhsePRyL3MpYysIq/bvLz/fMJEuW780Es1
HHCNR1tIF+g3RjYLN9tgJ5TL7gtqwRd5/aAYjuGc46tt+CVVsUXLrJETvzWTef3z
farrl5Gjt0CdiOfwa8dGdPdzDn8hXNmg1XxioHy+QVy3R4S6XAfnPVZIYSMNqg83
QBlovVJG7JplIjrIZF5HTUyZpPhXiBf4VMY2foSsUEh2od9ljcOFmU0XzhI4X6tF
dW7JtX5HmbdWmiiVA7b3PQqTIFCUxeXy8GQRcm2FWWWLR4i13k7/785n9XHCelK2
pP5qOVLOJf5gIg44EPKi0w+2/zJ366ZdZRqaZa35H3XpLd/k7qJ8CVfSwSK/FQEN
bxlDRFBCe9CuhLkxeNNlJ6UZtNVTS64/baGaVuVBgupiF4sg3IznsQWUaemt55qG
Fy1HZpsNZxoUt7kazZOrX/gUGRP/93zyVQnsx+tpZtJyz/TmtndukUVr1ohtKBoG
g0Rj1c2uKBg1p0mkDGRoSoOM62532OhitLlM0prpfnpOubOr8dV5zYjMgNwmEUvk
QSLEyo9O/zaRzL8kJE3FzQ6HWStrshAOgxffJ8j0nltCHNHDwCa+9dFE/MZc5hqf
W64YKq6eLlHBCITKXomVqyG0cXyZFES8uiH8fyk3x88yWuc9dlCbB7EPi7W+sVVf
swJR+z9Z/roH7FG1ftjr9Edxnrpv7YU/5XVTUAHHuLHBDo8z3k2tCp64+YS7floV
hIu19QqLrlMaVDHD7Vhqpucs3GZru1q/xeR1rhT0a8kGRdckz8X6FbIHyc4Q7G1K
a90KcUm6VhDfCVwM2zpTycjojG7hp2/x+5MkMMoclFsV+AcreRjocKAq83mptcyz
UqSYyK3DGRpfDJkzallQDCROKX20WIPxsnxVr/xiP4CQH2OHNbK6mZIKi0f5Ro4E
d92tmG331o0C3zRgxlEP2MkWdKztyPVPPwJXE9Tc9zIq6fhekfPWH1gDBtpmt2t5
3x82gmLg524N7ToFR4/RmpMCFgOLn3DPinjkMB7oGQpZkludDTEKaatv1TdBzmkU
2ed1EWytl29QGCh+q20EStdt/wF7mMJuncJRePdnECPTkI5GcVLGPR1QYwuMjRbG
G3z1G/SRzpCm6zO9Mm8TUHXotSHzyjqLyREe+IN1OJ4r3jziW6RZUkr7o8moqqKj
AIvX4ZG81Il+he1lyv13WS9nBbEnS7CozYdQQ/bcrmYmTX6dihDk7yyD/ROQfkTI
JWCmThrNNiNHP5GDB4aBWNlgsfsSJvw8LbrrHN8WA54MiOQasa16S3tuwpF7sKg6
7LvUQNsftwwpBfEUqCGb/vk2b6N/1KuWr/JRsMTqz6vu5PU1qSNhNryf80Q4Nr63
JMzGoDFEu034wCO67Xo+Lp+TC/7jOQrqOBg4UrkKYV16ixItfrsRLE7hCQzf2X/7
/3nm45vmMMCaJxMYCkPBHtPflFG3snGRxNZ95HmIC3Yj9lXPjJ2PdqBF3Vg4lCVq
PJgbkhBVTWcPEq2gdnCVqDXq3F2mGgRUwWcsrB8YMh0dN1L1tZqMRhPLhyESER4y
5rtLoQ/n9mchIGim1T+hvPypAuR/NEmc/TewWXCnAhguJNQp7dEEjNJpy7BruvMc
TVTSce5qDnYPfqwFnJRJOOngLF5qgoKCFr1OyZMhS3SzMCLooq9gm9O/Uo3kk3hd
MWLTshiqxAPAMmC3rqdsUBvRIXVK/mPZLfSEeCrTXZA1hgya3YPe1xe3/gfrf1m1
ZuVyHDFwdxnqd0oVEJvAetdL1q0HmZmcrBWlcRWe8M+2hrwSPIZB/ExDG8mZdSfz
FAF6mOowbkwb23hwRnrq4SDq9IxZ9JAVgzmwWPo96h0sK2wcUpEjJzdF0tamFcb+
2iy6w8qkvopPd/gWmGPoVnwQ+BnmrWnLWB7hQl18W44CS5mHR5gHzG4U4G/Pky5+
4WprPbR+87hcMc2O3oBaSDhWwzChxHVQB4r7kgZHJbEJfYv7CGF1GDXc5DVEHHjD
YWJZB2zUiDEj8iv6P5bnThucn85d79ME3HzrjdgVsuyC8YcIayD5okIbkdGQupH7
CtsJyv280PFblDAPmiDuaHmn4pEkmHq6vjQG8Mk7BWEPTIN8BokKLKWQqjEr0lDn
XzekkedQRVCzfgv+H3aWSafaYwaMYE0JTYkwfoudpqMNcf6QZb43GUy3AzADLh0w
xaJaWwxcuqoPA4a59miARR8Qma5TlMIdPVVccHFj0KX3NlHQCAtBm3EqyHocI1gJ
286GQGHUFJtuYExwLU/9FjM0kBVcPToy3ov0FyK9AFXR12lrOQsj96WgXpjdVj0j
0eHP8A+jnq2Xb2cqXAizEYNfMspzWA3DLszgelCpGypJT3vROZw9wXkEe0bJ07xh
flFUQUOVkXsCLG7v9aEuYo/w9fSQYxRYg8Nl1EjnTbBevbPPFW4Vv/nFhXdnvnjY
qSIe+tsXl1zELmMfA2PIonbFhVVL975abvDpwP2+Fzzrb86JeHAiB7nhXwGycja5
rAT9Kl7hB1UXcxM87PaA7Tp25owyEeN6TvQayPpaZZH+XJWDO4YWAHaE2nsB1ctJ
iz0w6wghk7OF1yyotazEObvdJacQmWDXHkYL1xOSCWLsEsT67TEkeXZLRnsByxse
QjDM62wg/ojcfT3KLea+1UlZGDCJpH0uCZdeIN8k0/eRU95/8NmuqI5+V8GXzlR+
zfV/lJsGQVfsZ2f33BXdvWIXr8esJpDgzSfI+j/ccGfSgo9i9TCPiuvDo0Ddsyby
NtJOM0SyFLp4pZco+J4DErF8wclE/YriW7Vopz/gOyD1atd9HlOeC5nIRrq4f2Uq
e+SuEUv0JeS0hTScWFGJ/BjsnvJdRMBqKxk946cZrgCdDfvD+f8sPSLnAGSg2Ei6
mnS4/qOccNSAVbrrqNfSKjCFHJOq44djM7epz6JJ3YGfwdkKCfQCSjzVHl4A+p8g
5BQD60uWZnaHf2oCs7FJosifCH5b7CGD9sIP68+pjCKzJ7vh/c/gJ3QtLfIdap2v
vOQENj2xATTXteugiWMVPA+92BjDHLLu3YXBIT5FSVGCdUnpem23+ASBJIJJGTyG
GapIO4SUDta0eSsBW77CW2XYqs2bUkgZV22vXQizYJ+n4pgAxn6/lsTD0HsXYK7H
q3AHIl1BIZE23mg4GDSObPLLsqTOY6FkrWoiC+a3RqMNnF4s1vo5mci8xzdXAgOp
DNCv8BwIxhmMFTPhXS/Q1qxIqBwCu2Sp6h2fMIoD9SADxncxvS7uT4A1DsmVoOkp
GinODU//DV1A0xnE2tr/DFx9lW4sIb10VW8sWbpxDIFZKTV+0Oty5+nA1OXwNCu5
MYIYI8fUFWGp4eYG+aqEimV72lj+XWyAMHzvVyvyW7nyA6+61ZVf6XvxhlyXOzWt
C6/KUc/i1Q/cyJgeByFrGBD6xr5n5kPDK8D0m99MIJ/BlFrsUuK8euWm4Oqmw4bP
aJHEw9zw8VeZBNwE2Zn68TwIGpHo3Sl+/7abXZKGefb+xxwkh2E0ambExX7b4xoV
4KluMgFNvKaSXeb3/hrFF+ehNFf2fCSkNmSdLTMEx49qe9GPEiTmrsdIsAGUPjU3
DyCCSC6wGUnMpgW5zmoVvGxzpiv3kvEUNxuVWvMu2eaDuSl3cNClL59e1zbdh8qj
BX9DLq/OE3vpmhBI+x8aABQ0I8oEtX+iHc4It1pwzrtdzzkPQdWFkBo6av/juGZn
VrO5ug3/j0NqB/CTKjfqffyutFj+ma7ytCxzVFlEgq/VLrUhMdXbmLK5jCjfRXV9
yJa05UAgh+WINU6USoJAIOrHHaaJ5CyMM6yqWf25dNV5M3zdoO63teCNE2zQ7jeY
ooxLbCgRXk9121JSMOvw7WblhO0a9PY1yaOthc1EKkgk6y+j4QjA/aeiFbzB5XQj
WMt6BPGYzm0YNAeVMi/u38C+2Vgg0NcLwBSAVvlToiiCVshJF+/m2z95hs+mwppg
9Rl5YMawUm4G34ul3uimQwHQWJuGBtILZourFjqkaBXIgQXh1c9roptO5d0jj87y
koeamNL+vaLSAL8Bi9Jv8qQVEfbpx81yDn5it+ZTAOwk1oqhnuHuENsWYWJQLHS6
GMQAu1YRtyfsHHb/sWwvZqFjPIOPxRKk/nhXerGujm6RgECKgbpyBv0h7CGacAIK
N1/G4vt+63idO6WcuJgmZi197vVh/9Msa28WBCZqAEBDjd+rHFDvP1gAeHiHJ9iT
acOG1TGK+ssyRzwfz3EHX0grLNDeMx0ruHZwAwdODhMYy7sE/W4alpMcSRF1z6CK
ru+OsDGIGZzugOfuVyHZYsd8Nu4nucb20uwRwBnbYSuvw542I0Dr4tn4DoWLgYjD
rFQRZR59lA226ead8Zf56+6ltbA+yUC5k3RpZtEIM0PCJ1FT3IPCH9euHkjATHmm
QpriGIky+PpGHBbcQdcC6DBL/DOaKQTLuSXUn34GZvfx2obWwZh61GWng34TiefQ
C/nhZE5EcXAFwQo4gOasLnns9gTBXTfPZTvR2UGaiIRoGxZEwMIo1C5DE0SBOGat
dl/wnvclnV2U9jbw1NGGhoezCIhFNl2K5HB2PD0vrfHfDaV2XCOZVWRy873n1+2d
vraWEf08Qs/p1yi/derKFKfAwJJcSF9r4GHOYJGHYXdZVj7arjdj7P3TMntY9lGP
XdoST/psOpHrVf+1NP/+s7JbPMlNuy5jnl4sYn8/IotDJKJpmq/CNEzu9uoumPW8
Ty4HDeOMIOvsYzXaAXhqfKcGV1xkprWh+GIAab0MLCiy2hgT2HnoDH4HVHEQn/+K
ISUq4Lf2hVAb7bSnvfKxk9x/BWXmzV2aYWlz5D4QysSQeUwhZfKisM2VnNyDqnl3
plNUc0KYGeZx2Tocp03viiRqIW6w+RSTHEmdU8UI5dfaLBOBqypY6MeKUIQ4/WwV
wxNFyNduF6Wpg3ll1T9VA63URraLD195hN1WRAl48Cg1NQ+Kdvf5qUpXO66Mr31Q
Yz4Jbi7Kv3TAkyA0c7bBi7U9XHbKFpaW69czDKDdi8Q0wbogt81xvc66PVED2IvL
neZXOYUdutTidMJKnZbzWQH8mR06sm7oZNxJQGWXXnd9Zl7pGaBnBBKXnm3/ZsnV
fuS1s/Bc+G6D4Jjn2WhkQ98VnVFf7inNciKTDJIdk/8ehHIKOvuYH9W2JYXvpjog
cEbL1+TYAadcnwjSthebXNrFWWFBmzP7nCCX++Omq+FabzqSBPVpfBcciq/qyXrq
M4OoE80fOn8EfGjMkKcKcgOU9fwlPBEKNNxHHEYlIzYQ7ZFJ2XX/tS0f63Caobc0
qJH5490S4EJtuJU15q86cN33UlxOQ6kVsdpQXY9e11g34vdsL3JCCJLmHDa55yJT
qJ/JRoKlNkSRjU/MNfuluYEOQTOGNVAYDnK/8yM8MdNc97xVKEszfPimw/+Wzp5s
ENRy6OT+g61e1GhazOq9fWQXY4Ao0qtwfXKxl57BvYdbZ3LwVyI5KotSeekTAO+b
fo0f9FgmWdBCKOk/+VsCK0x3PUZr/6wkIWywzvZTCuc70ACDLBalKYUsH4fw7Sm7
y7vXlt9UKERz57aHucEIv93GTScXdF56Wb+bDNP9HyVu4XxP0NQyni5ncjJgS4s2
lVxVaZ9a12mu7+Th5l2Ew2ttBcahTlVG61cS2lGIQ/vEVDF0Wzwy9+ADbS09YIhj
trXf1dazk05ovqll+Kow0Cu7R3F8bmn6r8+L4RIZYOSPRhsCpcnLeElkXLxX016e
DpcUKZGR3wfisViIugARb56WuCRx1YrgEsUaWSmleetXex1+AoVt52urlF5/vAp+
ASC6JJhWaFEFMXtDnUd1wKLKKXcRnHd6Lq8+OyAfGEtuU2Vf3ooqHyuSje3C096v
DuHOWEj0JpQ7owbz2dH14wsxMe17jtuIgtgF85K7f7Ies5gV4mUq1rjxlNH8Qx/R
QHE1unvIgBw78IjdZ2/LZ+Fra0T7yK8xwwtsrSe++KdYhKQYsi8gPlYVf8zLroJz
REq+9HS1KP65zl8K4Zxh9W39G4nyScNqTHJ/1TbVSHj9y9c0MtQcFkl2spttvlBK
upSjVzobd2R62a5gxFMYIjAOtlMrnS69HTujmgCtNLYjJDCAg18/kHiwZb0X47Ie
h0fXnj/eNIB3Y9ZLmYpaevZzMtTn51YM3I+L+yQS1/6WWjnBArTWcl/IL/PV04wy
VA+zPWN7lSJEdyFM3qBf2c8T7xiH6y7xkTyl79gPr6SJzZ/pDT6S0gZ8kFRwG6jv
7BM/MnZR/MSpiDnPScSn6mOFADoDIZE5v51mJRUs9wJW2PCzKSBG1GAERg2k3pPp
FuC7Bmblo80X06wBJ86xu+fUogVEXpnVB11S3L/Qhbo/79IGwpV8La7oGg1Vv/Et
c0Cn7oWDOx6nYF3MBarw3ewFupnj4HfAtjPbOixuOG8JS/MekHUDFlLsiULyJd8V
OMhWtQgAP/Q3dF2A8DsIv1jrK5SjfVXVxYGZi64FatjyAk74vj3XMHALTAHGA7sH
qWpvad/bTIobDt7VUJWc/qlkam4MEQ+JOqX0YU3eklfzAX3RfwYThiCUaaCi008o
JWRxhw0uFjg7U/nL0OdCD4xk9413z6RyBfVMGyMw6N8XCsQjik7+xrXW/SuLYvmL
/xRYrlDY0fD/0hPB96EY50zB+Jb3OP6U+8qVIn3cYPfsEn4szgUoZLpuHxNiu+9X
9KFk5Sq3iNRsNaObLbcdn4O/kiMDghW8iB/S6NrShzVxAMJm0hjjeDGJz0NEdKX7
rLrJJxC6MRjnRy/21RAW0JTMsweg8KvrVU6XstHXROPfSFqd9B2kLhjdkqlYyOrN
h//8avDbdHng+jwOJ4cSTTOST0J54DYuYYXh21ybqICPCRXOJ5wUfGMQ6S/DB2Rj
IuN6mIto/A98B5QSDwU3do6yDjfmIv6urGTdDCT24TyEJBugQEzOUXZauqTTaWQT
mWC5gWahPO7VPKGzJZj0BGRyAvfBy5GMMcWyRbGZzHZ2un05nHGdXrLtAtTDmMk+
1ybkREAHE9pI6DMZPJkBwg1846Pq4X89xe9nN54uXb2O/HXlYsG6kwPvfm5X5B8I
q5vqXFo8Wk4nsXs7iBPgiUSbaRhHZd8oKgvEKNMRooK82jPT343uQYr+lwlFILHK
wqd4FO1HSHz2Ui4/o5dfXuUQ9xIV6J/ZCHbNTVV7PBRIpI1MopRc9jSJv5DKLaIh
7EZRTLVO9dZrnTY5/CI+HPktsddBt9TjQU0+XH5n0pnXidv2RAQJPQuRqnIrLVzg
dC7o3r5W5wpGlol76dlAjYRLsPgFjbiKStrcTSnoIQdwiahychpO82ziHUR0QxLd
prVo+mJRZI9yx8F25X6Qs1JxMZvxd/D+IxFklHa83MVxPVxZzHxw4wllIkQXVV8M
Vp78FSaGXlbRc2Rdc94hXCxzqxcNjBKOYOiouyKXc4Js2V8V/DXXUJw8LVZTuQBB
5z0j75J0Hy3yjnV3CNZQ1Zrk4JX9/7jSjmjk/6es9F6453BBaI6QKPDhsdLYLnio
SwCTWw92NG4/3V2diWrrpwZfXcb2ejisvP/EZLXBVP3LXJy4ii0+7/kJVVq4bDw2
oqOLkp3z8rr2xAw1xLQlZnT25cp2rSr4Ck/6i7hNzz3k7UjmHT0xeu8ppuHoV1rL
Iqhg1/pA9hwi+LaeWwh2PmzfzmB4tjP4oz3yc1S4moZnSE3WBXobew/buQ8SZ943
e+iLz546Le84auSNMH8fqUvCJJeZpfI8LI5C+XvPoUT8Aj5PNMZEudPF9vSjFoX4
bqg2ABqnqGH7hGs2ZICUuWA55xJinoBwSs6ZWp4c77mA5d9rJARPQ81lmAfEq7Jr
F+F9uuxGg2W6/h7SNQIW7lKjf8+fdFyeLksQ62tdwvve3W1wcEYesDMl3PHQlULV
pAyQua3SIcrLTurDceNHNexqJ8WlO0gAHN3W9Vt4HBfh2ii4/gStfngd9vg7m635
CgGS36W7cND9GDrOKnOScv4fMSjB0IoJ0zjOydjuLaVwMrvI8HIkStjMkwhuhA6b
Ng7TsXONK+RRGn/v+YkDF7ge5YxeZcuew3iK5dlQ0nKkcx4CFnmqFUctvMahm0Cs
2BjKFLeMaak0WCMc/QlkWZG5RWC18neON5d/Lh0t1kovVmiWdtwXIco7Ibkq0wba
Zi61wLhtGxW0XZFiG2Kjsvhql6sCtgVPh9yjtv+ZANPr+z+7b2EaRJfvuetugQng
MG0gqsdt9QclkcFw9w7gzBb7OAOn7NO9izpitbBY/JKbVvKAB7s8PwxXg8zeUqjQ
+vVn86Fp/zoj5v6R+7fHb5px2XGHdf8JxXqVYZnB6ZO5rKWmq6sXeCfepIxLZt6k
Xif1Fbuernn6gbirN1meUucpY4Di/kl37PAyWs+yQAbdQTr7SqRwl49pS1pi7duT
ikPH0aGXBxQvJK6Arh+huW3T5ty8M0ZX8cn69msXZ8FmuXf6OhtJ90Cl461QwI1s
+WVapMHVPlvJN1cuc7BJU7gg+zM3NYdRl1jhUbmmWK0aMpMHQwOxhQQbkQsszRse
Bw8wJhgEHs6xDp94/ymkaTWQzAjFP6BlZIZz9o4zOMKo4xEGRnOzLWHnmWGbogee
gHwzRSFtQgFVv71d68dmda69xNxs5d8P7AinZBDFqvaxDrmZ6YgwjgQy5JxBpRpu
JxXF3AJ2XVGl+MKi6pyIneGQMStkr23Wy0C4oW1H+/V07USxD0Z83bncz9o4jqSk
v8XA8icm7NRZwVo7oiCGwGMSrWHoi0kdBaeswjz5tbIaC8Fh4744PCPpS0kgropB
ryUuE19BUsbUf04i+a+K6VNTTB8beelrhvojy1vlAb+NHzfQn7ctMJQr8al5R5OY
Pv/jwxiTZXccIa/adBkHgAc1mljWPsAzGR4dpx1hpJDsC+dP6siJpgCeifO/7212
s8Ez9MNp84+Kh1sQAQT5ItJmghwSRENl2PbWQDhSMVEriM+fNCT9sMDxeEo1Zxnh
7pCcbWG8gGiyeuhzhfv+hWwbVKIaGePkJAHHKYKkMiC2AOlLaSZ5ztScH0ofH/fG
8WOR30S9DrJHLK8P3wuwacIZi3AgOIDq5VLJEHcq0/npneU5++yBIeZx4Bgf+/5U
PDs/cuqHHnb6sh2ld+5WQGzIcSVHL44W5rAjYyiTb+yDcLU3OONoQ7cdUs+FCXZ0
aL/DIF81qoDrOqLBtH7Y+t2N7MG9rIGlqcpI3g62UtiR/xMPeuAGRyLYH+tM4t0B
d03j+trmmKY3RS0xNa1YSTeULGVsq5WqvyHWi+IGHnKHWJj+Sudy6e+U5osVAAEP
j6UplYtVNrCiPhQmrQ2oGlVI1r7Nyd16r0+VIvMzCIzk44IXedr3/JFRRTEIlYUZ
s8Wb+jXdExhNHEkgeWikEG/1d5C9OLnbHurANRpq1+cH7OqjXsRnUzlGZsgGKY+L
ylgLSP+P0AoR3qGvgLdKLrTC93x6d2hECkbpdeL1wvJtiCgGg0OdpVQPcNa7pML1
lvlUgbhh7kXf0A1+y5tmoYhYVSZtn7WINHXzerQduLXMnxJoEZbd+HHMhENckNrO
y3Cmz8Z6XRBcFUGk6e6tO1UhG05Vp0ec1Gq3RVORbQpIloMHJj5YUW/Q67l9emqi
ODTHvxMmqvsu9Y++rIvUKTIEWx8aK6f0gNxHW9D8m9VhcYpetIbV8QGgagQWF4NQ
9HojlHn3XiFRJ9a2ifzNZ05cOHSmhPMOWHD7XI/OGV3lhql3bIxcenyMUWJaPf+f
fQ742Gg9dwXffYpdld8ikwgVqyKPGYwDbhiBMzYL5ScfLaHiwjraCfKnsxlPwL2P
oZR5DDG8PtICV2fvrYUKhc8tUUil3QQcv4pr4J1b1R0Mu+bdewpCYRlPIZrl01ka
71cl0qmFqrTL+64/qJTCSrkihfo+Ja7V+ovZe7JCE+/CeztVjIxSoI2nw6d5Lfc3
nw9kHTQnBVyKneM2pS8dzTxwY58bsElK31ZXtv8c4Nkt1bJK4MYSC3URv4vciJEA
mp6vSRDv9hc29HToMAO+WBBOuTHAYowAW2bObW15NiIkVkxjbCbsRvTaP7oNhsjD
wIHecw4lIg7/hZcPMP4o+EX3V7qG7OGRpG3ET+eVXoYpiL/U0eymM3qROU6t1cMJ
aKBKca3MT+lUMPnd0SLpFD/+05yn3EPdMzT2Uxl6DfupjP/q5CxpVncQPKimpQ7W
k8BXdVpzlyavQwjAu5p4gqCsgvq7YGzenn6FRuEPCE5y8nupjy7egnIiY14Fdbdr
0AYPiAXIwZ2+QlSL7GyBFtzXjnW+39nS41eTUwv10vzauWZy71RU7zsJSXT4/0rA
OP4ZVwJg9sNtNJDufGKh7YDIbvroj+d8QOjPivOLnnGKxkc4YTzG1emhzVvapU+P
J5T2iTOcuuOX67irRSj0mqa8i0xBE+4dL6Qk/9LUjEzZ0AyrVHFDrzkz7OBL5TMZ
VKJG4NcQbIJaRnyZ9SAyOLHfhMixcJHfCAneouZLnZPv+s1mRnRew0KqSOmBpchQ
uLE/Ac1RLV3yDI8mL+rJMRuf2iLjls0e6SzbhbiODsYF5ggFmqwoYXgPzylPqI4Z
zGPXIxNKjNDsUCX6X+4B+WsMPAg/ujq+yTELbanB+lSOoehvBCbEAT14374oU8lH
i5k6YY9FrC2OZ18Ej4RsIH+TGwZ+h2vje1Lyx80lBsd4OBKr188ehLSiuTMlQSyb
ytIDPD/uKFzWQsyDMUOKxd7Xa8nBGtKTUxOizHCwKyDdIleVHiPl2kW2/PtJoee5
krlncBADcj0zTPXCNxet20S9cqXN47vKJO5ocz38m0y/Asahm+El0J5XUvt+iF10
4YOnXkMuJLTry74G105oY2enL/jST4LyInkwMgsUPE6gHjcKLb8ln1FIycaxQjxl
wcjGl51463aqptJeD49V1HWD/wkfUzqe1liL460QJ6T8LGHPtmyZDKYayUx/sDok
Rv+D7KRAP2ivBa9JmFPmxEB/MJNtSfWxI3A16hFzu4iiAV4mIbQ9EAFli3EHeIFT
PqxYa8dXjVTeIHkkaD/AetuwV4HmA1KOw6BBUkei3JgwRbrkJdQRhS/5CKjscU0j
Q1ql/SH1aUkUMPmEJ7YhJ1APSg3P8DFbiR5JUckr2UWTzD8fAv22qWBq3K+9YNQV
4wMAWawM+U7JxdMuF4ia2w38sZgFh3RRR3dDUsS4R2Jzo3x/O3VoCPfM5RaUlrKV
y+Eh2V99lQKIWrldbx1JmCH8ScVachFuq3tcPqprDD6Do7ablHPK9/6NNuteEDcI
X0KmHsRANEjLP737K1dOOxIFDSXKE+P4T8p46plgDdkDYaAEOjvp38BCx3swJHUn
DMz6HrCM85rJYGII7YA3FovBPlXP6A2ieY5GMaocxrG76Ed6EXdRd7kd6nzL7TC7
V9YbofNBxLD/xPMaBaJkdwC6vae4zy5L1X9QzKu9kJic4/HRXZb34HfPFGmQgHvd
wZjyXrE9kqRjc22b2Il3cZ75gQyVDMCwDdPOlp0GdfFXoIziU0O0KsHiTgi6dPfE
Reo8k/0F0eLFalhW4KAB2IrAhD5dTd6x5NZWbfMvMpupNYmNm1uQk6WfPkBVU6D5
ym2vCyIsUrRPE2m889OhqbACjHuTEu2JzE/qDCSXsi5jutj1rvrnseygbWJ+ocBZ
LwSZq/glXWq5ncpie9kvgYW7fXQb+RqLFjZBOeqdpB9of5zgv92qCyLkQheyEt9x
raQbsDxaUQzlwFLF6K26G9zK8LTGkSgdg0G9jpT128ZglgMaoUkTunY2N3b9nTdT
sG4bqJ5f6+b6Ji+sGzn8nCksAFlqQSkuXnfLNfHM6Wax3mPfNYVk3ui2YLgswFWH
VchUiY5cZ4UcQa2pyPb76xw3DXqHPK1CFBGHk4ZRYg0fYVvsHkWH446vbYmfHgNE
zhVlGfoS88HiG+rmyntupTWti+WuOAj0FS1ZefAoOZFJgskkHt+lj/lMW5nwDae6
MNJKxxge7cwpHo37nBtrsTI9HayQzJE3Wj2z2wRgVUdqgwAjyQa+7Y8zSwVJsvK1
JGvk9rkOJJBPBipNkmi8bnbrrQrGBuD60QJyTu/qp8owNUIMEd/tyW/V3Tsd4FCT
sjMuQUEXPBiq1vMpx2W40o6tZPjFlMke/tSQqbVydFlsvbl9QZ4aIrXPREie+DOH
eGunB9WZ0ALCx8OYQkJ7q4i290OXNvbNDcDDBvHLwPI8L1e1N00i9DqsZAwgf3cd
qAEesg8a1cT8p4NzQHklqydifsqUdSXeoT2SHMn5JeS6EzTuoxwY0TLcEAVvIkDe
B611/xXCz1Z8tLeL4I/TrHx2D0bGrMjmFKZobNvGAsH2iUv+J5QWBSip4rdv6YEf
X/sOub51Oi9fL8FFeIDEd/xzZYJn6Z0LLv3eB/5n4Y4j1sMIUXLZXABT4AwYDCk6
QYtrH30ZGog35//z7FE1Fn9Lt6g5Z27h/dGlywhpzTa1r4CqoKPMeolWIowWUVO9
sGLLBp9HqODUeDvZ8sWI0cEaDR8in1tmi12Ebpwx/vPg2zbhVO74uxmLFbR8d6OS
gbxFJRXHoTttlXoGLVQgHxm/rIRxgqY5k9fYZJny+yifX7qjVtaYmeXB/NtzAjV9
y4VlSqMYts7xyoHb0Sid5bO1TC4fczpA67VuUImzRHM7fC5fPSaH+bbm2kBCAZIi
Hq1GT9Tn7Z4vz73jYPt8gbMOXTzFW0Wl3RSs6sJV5bUZraKL59+qf3hZSo/8nsPn
gLmeEtr7g2URLPgEOOupP+Rri/4/hWkBSrTnFxd/qeCVSYuEEQQEHAr1Fx2kH48c
h8ypzKeoiDWRHJhyJ/U3BvNBLOl0r8//ejkE6nmaHp7t+Ghd/aggdl6wSj+sw7BT
8aFzw3y53zEV1ErshWM8i7G0Orp5JFuiI0iv9XuE5EJbnrOh8ZSL02h8vKUvZi46
QSq1Ir3dj66vsZNA5jrKKMIkhHWu6IL5WHRr4uDn1GAceD7qkcdnMazqCw0PMzoT
dzqVdBAKNiE3ewPrd4UCHq3cztsAPGvZTyF2YmYB1SMqUrQFPmHEIqsYTgLf1yCw
psvYxdo6qa6f+c0z/7IuuJFXHsl6msewWuXEXBTwwv40R3/wL0TmlWNLeg5aIe/T
jR+l22sYgmzKq8Jdc5OwljrKdehOrXY6YQnfw60KmraJZ1BsvXNzTrM4jvGc6Xj+
EFnjNww4chMNj8K4U1mB38GvmMOk1SCVx4kvw5e0r8EEVtSUMqq8g2b68SiO6Z6U
tGUHvg/ogyDZ/juQAifQvyXZurgBljqbl93MWUgS01llnt3zXcO9iLMx0QyuEODT
6EimuDjHArBFOcvQAD546Fxu9K79fzZqUO8D0+2Lss+yoCJHxR7yAe3oGpht3B/g
TpE42YVtVCQyRfjJzRN9h689KwwmdjFmmJThkYbkoGaWFJAT8z3ErYBp+mMv1DzL
kHlbh9VJZ0hd+w+UDO3Js2A234Y4tJNXURaL9JSKh0dDQEtHkt1+DBG9Ib7DK8OE
39h1xqiFYzSMM/a3sSvFs3kPVpXwlNwMvHXHlgmWSoByJQXriS6f4CA7Xghsl66A
k3noZIa9PQoc5jl1u3Oa+ird2Gwl8v7TTPL+PE6CvngzjsAugKziFIxKnxabD2oN
OzqgbQQnZFGPMbhm6D2rwJ+LpKV4y0U3T96O46xAL4MJfk8zRTAqkIodjWm7J7JY
Sewa6mYkUTTE4tIh7VJhwGE/MScoWU11n4J1JnDLBd+6Ku+RObZ7c8Cjsbusq3s8
tor3KqTpyLTlnOqoibQF55jaDlaOrfjQIKrmgUELiAEkCm5qFHaqV2xLa2gd7KYq
bpSQP6qPLby72ki+JJ3bdmByN3yTf41h6e3T0GnDenW8C8w4npa0WlbKSgAOxgWW
l7vkIptqwuEO+OnDXK+Vge4lsAYhvv5H1mUg84OsZvZHoS/s0ghX7AcDHJG/75Mt
toCIGKW/TvxzrYpjPQ2DXR75K4HQT20OoWY8NSVHnOsuQbqtn5WshZ+aU2uY8imB
4HSPW/nP/wlaOO9fC5uDFs5u83PIFANuMnynDWFIIY5/TV19I60L2h1Vzw4JJb1m
IubepbTnNKd5eN0f92wxOjVc2TIeOeMvDbMZzylDDEefqGfz5Jlo91CXSmbYb4pD
KsX4TK3b+o7g+X8fNslieiY5IgmHGLzh4RTx9LfnabVsmzZYoXUGH2YjD+AXjtsS
DD/gkhYhr0lSlhhH3JZU5dXF3OPh1V91oXdSjXStSBehvDnQoM/vEK1NQLv/Xiul
eHlc8FTENbVYdpGa1fZx0cP2L9rDigE8F0SkoivUhEHtXAfQHxNWKbespAMqZEkC
LTMmKf+11RIRG2UvAmhvuTNzoETiMo238FSh77+qU4dXXxcc9CMq8iYP8mpJcV6M
+0DNT3J7V0OOr4xQYFl2iZkysLtucTxBFV1yY7ahN3L1bWNjasMBs7kdPnnmFnb1
Tan+UGZJdYJ87lT3gIwHbCfQhScsqOkQJxbX57hDfWcVZ2O0wDSbQwJt2omF9HGk
tpJgsflV2p3pjP11n1ek1C5yw63DdjLM1oc5zklM8qtSVCyRsL9xEQwcr9OnjPDD
5HxXot5Ot2is7H6G+Vw2rnKZKy3G5VVpmPvHcGVk3X3dbHpSiud0vDVt4dp/vl2Z
0zCwW+9cXkaOeiXoEwjZWqbJYWOs2YV++JShsX/VMlq3ENncgPIa4qKjI3ZYNERa
s3C/KzWsJ9e1AbwgtcWiexah6AsCnE5bZ1bAbB09rRQQCYSxcNHdUYdSaXtPrQi7
/0pI6xm450IPwbioTljdUyRgQ4KfLacIZMySG5XwjAbAq8FRZZ4oRB+ZKV0F5bew
7j/us+bGCQAY3V11F8s5nzrDAGL8r3BrtK04fNt4xMNm50jHMi2ddRpXzm13AqUl
aK/VY3g4sqOZiplwONrRG3q8r4DlmO0ZiBD7bv4DCavOoqvfwpD6KHKTpppVySyZ
2WaflugEpN3niexqBz9svqyJlN5eB2E1u/DXQk6rJE3xcKbZ3oCw6qjN9C81H7BJ
TzQABRieCG0bYT3zMoGPSTa0/dCfZ1785OcyOKMIndkRDBvvlq7Q+SdmCW1HZI0v
MOUUj8pMW9ZYq/1o5kB4ygW/u4ojMPCuOoZUSMTUT//kvcQcSEYA9n/xGQP21Wql
VccsQhM/F8ay8I/Mjy+5weBwuDgSG2YyBbZ45tZflWvQ4snWYfLEmFu2TRh4ge2F
ofuht08PbPPnANPaxst3ldB4GFfS6CP0dRlIGq0wTPlgHRplhcERSkQrmwq9Qfqh
/rz3thGdKQMNkZWTiBjCQyT0YqqWlaRbaJ2yy6KVOSMz2j7KjtvzCpjdr7fSyZqU
Hrz4H9Jka6AS7yfJFegselV9ejJClaDZgzkmIJRZmQNXDpE6dudkQgMXX2bZPmft
FwefOr/t5wK7lIYzD5MO3jtsgGUK0KimWoM9sdDJjC7FSVftRaK4+fNmIDiaGixK
zZA8kh8XytECIOkjvNAyqQNiNRVKqZ+Otu4WuiRAyYMVQaC7S4gbOHuCBLOcaA6P
vYuuq621bLY/UeEjbJffO732j+Jh4+8/j5svZNOP+PglW/oTFIK+4LgS/mthUjQ5
rXkthqE1jraGHhABli4fsyBdqSEGO9XR56AvSXFfXyvOZwbULs4dZGnsPMzPDIhi
jnB8WhnyvqJciQZuWsqloIGOf9Myk+VU3ZssrTZN0EGmkfYOaSmyyCadHEsCBsh3
LXwL7HQkz9cbqYEbaKMdJgBaMpoCWZHzP6zA1pmVV3n9geQ/viuX43rz5mh9Item
khBJcpYYH8ccSM91I5tDaKVM+Uvsp323JS41UL4V4wVQshIOpSXPUIZ/Vd8/Ef8S
SZxE6+bIwH1jL34fXqXpM5aYJAW0CjkpErp59oCmfcHYKMhhCn+6KtMa9DA7mdlq
2TiQMeOoW1KcOKpZwayLTv+GX1KiFhPiEfsXMIWRKnQknkapDuFa1ytwrnHsEeZb
6/GI8U+yIhI2R9Wdpjll4Rt9iQum2pI4YdwWIMwyy87+R7pFy0cucazJzdPwjyaq
8dsWLWBO5mkvkpfSSqHQM0xInp96a9mbrchxSPtwhY/wF7aGg/26LNdJpUxR1M68
PcPqQBa2V5Zr/fRbZiZJHytoFyK9h98fuYcfReQf5YP5N/n/91xeDF/MgAFFkVhH
29e5EWsdsAOK8CpmT5gfVwH+OgO0C+76gqhBQWNuXMr0cC4juTam+4aNAGIHfzsR
LUHpl+bR3xhu4/ISAoi14YgRYNj9rn4DmvFfj7PNA69nu508cH6e2eyztOirur0z
Oj9RY7zdkWPIPd9+C9zc/BOtcaqwJka4acl9q4cg+AJuPr7w/vOxU+uRFhgGJ6JB
7EkY1HTFY1/r+5jAPdRopipMtCtsMKBO0QMuEerbaE0tjQDiJ6ym9Fp7nbXKgYZg
lJ39V/BQHIL6Q5WAbpxTydIO+bOfkL8jHqQEJOM+jzK2ttFpCISiKcPECnJjPqHY
JOvry6pS7p9jzLvfkf16dCrsbPBcvjdKXR6BaYQxN19/9QmI6tyYbStoVbJJFsNf
/wIrq7Kr2Ieep8AHGkT31gNzSzab1HXjZ3GB50Vhl1SIWY5g7Z0S8B9kMmmwFLvu
UVghk2Sf+u5lHFFHTfW14dGx1O8TAdO7QlpAQXhWz0m2gPVUmTfB4xrGcSqLuvQe
SaPthS68w9nqjp2EydmUl0vZQQ2LYrCPE8fWESZyOBdjEsbcjxZcdKmo+pbQ5Xri
3cCGIqpcvlyNcT5qR0OhRsGjv63BF7wTZk74vIemIvWjM6kspRmQQP3EOwc4TMUa
9/NENS/1mEl+SCU3FhJGjK0j/PSfiwf++9NHceFp3GgMGRJGdsyiyqHsDWd1zsgP
3VArWJ42xnAF/PgVNc6zxfY+eMj6wOCPjAOg+fkYjKDD+ZvV+0Prg9PObs1iaMea
aE4F5X0i7XAiLVOjwxUec0ZiqwJsF92is/fwbM/aiWSZcptpq2gsHcu2b25mWwtV
9NOHo4C/utJHDBThXTkeBDazsC1ltsxZWCbCqN0KZPRz0FPedWLY7nwHgzwoqnPQ
u+430R6L66BOM0xWhWMJP3F97/4a8TUpZtIITeQiG0Dg06hfrbMTET7psCGR0ee5
OGtZAOKihbymrHVovHodmgwx9GfdzsmDtk5I6RPtblK9ltmX1HqvGDSHCrEKljrW
bxcTpDw0tVWy3UCA9xuCboRQ+gek8wGrRJMRQp14uXKrpg8p+hKceijXqRsntVAN
kxA0CDTkloi13Se6G2ABnwqHgPCtKt4O4VgEqozkRnHwGDyU0NsEjpeh4uq2fJa2
LhDiJ8iJyesraauZnIpniir16lGM6hjzrYHeFavQYkjaG7/YKZLtZoE3R3sM+Zue
zhwohaUjy9pKz+XThdDwGKn+ZIpF6RbJsTqnQXG+v8Ka8tjVX8DXWxeoJdX3YSJy
thIgSYFJdpghUmTvdT2TxXt/FtYXM94clUqT2DeasdyJsSFMJxVCFtIseaJw706P
oKxwLG2TH85HNLuFxPSXVPB1sRQ8/V5FdovN6dm5Cd1RW1GkC2CRVLWtf3TYoHkt
KKKDsYXqhp78W+CpEho7CnA/K1ztW5AqUuH7XXcv+OBfDzV/aYB84Ik0UACir8eE
6mQ7RP64UCkzzQSCkWHpU+7e55VgCZoGYp8L1AYouvmHYDJ8N3ZAOtnVi9ZF5Vu3
7E/CQ52aFeBVhKscN9ATq31iKojK7snYDeeLr25Ap5dwIXKzgDTnKSkLihFWh0zP
O0eZY24x1hXs15+amdm+fZ/2n5XdeoVZVfGAqoELRbMbivbO7B1Dw7rVO6tgAsMQ
u64zxcQl+W3umeLD3G4gG1PJSlrWW8uIgDhEt79FTMY6LfPpKifIrFbGcZLLZTt2
WQf8GjJBOhdjng7MlKU7vgCY5uM1hPFN3YA6f02JaV2U4niPXWrHFJT/RWXUdNqZ
Z2pAuQxvS7D0S97e43RFPgAXVFGFOkuDyHse4nxbZTz5XaU3IK4LmTyM2ZhOZIub
vq7gllyWoeljxVJxjo3RXsAEEQa2Gr2cgi/ep4aVLb+ZL1Ney8kq762fRoK5SWp+
0yGDPndajbMvD/xa13WlLDYeeTrtZ/8aIVyA8ch73cFO1kdCuKOUUWKCML2Gq+El
wGOuMO5xBIIT+zH1+NnISA1qO/Ooy3tEvsuAKW7jzcSMexQ7Wm9CJrWrBGLqkb1t
GbeZwiFWJH3tVN0Ujx2OUwtsSBw9fiBDWoyroEqSIIie8VnCymiObeBasjUYGUDW
T2yocK9b/RDBa07bVoiv65kYLHEhVqJzWq0Rz1Qty5PJgcVGsOjsp5b+h2LHlBk3
x8J7EqzclZ/VAycbr2eGj82rKwmMNZb5i4p7C4SDTq3Bhj60S9AXH8cYv4fW1XHG
hP1Xy2SA2E+7sHlqcfaWFFbZTAn/sXNNCSFH7wNPFvo/RGxTu5Mjd34jvfo09MfY
1x8KEl6XO8ktBBBzZwvWFWiuD6fT46FJEhPipQPasrW2JHxCOfmNrSakpCZgKQlV
2sIRh0S4YOic24pAPbu06eYoKH/yJhXaqzctlOR3HfHGikNqCHC2rrpQqtqpFJVs
ZGwodnmRm/Zn7zgrhARtfU2BxdY113XSh7ZrKMOfgoHaj+0uXvhYGHPI1wMDWb3Y
BLC7XaFYth+o58MC+Ew7kjyz+YIbEzi7NwW9Qi1BzArszgQ6ShHwD0A/pbTcFXgG
fFy9ozDzFjTgCz8UFvcEISje4g4HYRZxxjd6B+pKPueypHhfqCQg4XPlxjYs3DfW
zAeP/kV+2r3A7p2Uus8PTjYfRIUUlXmsIXtmu1gdTUcqUVA6FLwyz8Nc5ZSmFJrD
RmLWvguxW6yrc7ZZGnI62saz3GHKlXPpWwasGwK1PHxxPd0dQlfaTJB1I4BOA6ts
2svhEicFN5nheTATq1elqkF1QW2/LTJ2HsXySFPrc0bmTzYtZGbB8nY9wBm9FECZ
O0ceen4iK0LQjRNjFCcNVqEQadBlaCxmZ6uqAU4L6Bzpl02Pd/SO6CwBhByBLszH
0Tje4bjzSEf7gP2PBMJdSrRnKDtdD6YAu0qrq41srPPXul48rIjyFelITAQ8Q+OD
y3OLt0orVA7duMy9PcE1UBXAPPIJNnQwxIywp5Yl/jo4CU0+G3XzMasYbobxwSXa
dP9NXzniViBjvdrxQLlwSuZLDB+bCJoEybOEBzqO4oVryElWRDdPblreK67300k3
HaNnKpKouqGrF7ZS6gRa0nOoQM9BPTNB3lUK96IsOxABTk/K6wO8+ei8xEHElagS
uGp14/PQpjGS2cFEBqWsNQj93XDwts1+cp59atIIgKQEJ7yOlaJIiIzgwKDjBfv6
YAQo0uWffo3RBlzmOlhC7o+QpDLukw7o1CVcH7M/1kwojKYcfUn6AYg7J8/IQrxw
3u2daY+m+m+fRSfVc3t50Li6IkLsj4lIHOHMu6wcKhKpArCe17jO7Njm0OK3EssQ
UyZi3GrSl5CYsL6HGyNQf4JMX7frwye30hi4RQEE+qixkcYRxYbit/QLvIKS61su
dxQ/dtl+Ujf0T/1XKNf/xZhzgtEvLXfnvxWqXZntMA18nIvE1ju7opjAN0ZuSWmw
1Ns03/9yTBTZboh0lmrLGF0EVCfQHu6pp7TrPmYY64TK14OhXlemmW5CJj9UdNt8
knpBx5vDM+cAG/C2uYGSWs5W0L9aCfpGWwkBCN3kdTlaBOJXougsZctw/g8dhrSN
JdaA/Ri0yPk7jP00k/3otoWbU8nvgFULeoGpVZkwtSKNM4jhpFfVB3jj4TgsMvJH
qF6z18cFyZ3hQldCkJMgNYwwndDBKanebnD8k3Td69Y0+exO2XjsC2gP/JL2eM4S
VZ6GMOU2fFQvgwHbiUStk0v1Vd9UyD0b6pyk2QYy/5ZyhKjGwm5tZ54V7iHVc7CY
7FiEJj/Be+HFlVfcEOaFBRg5+/4IttipKos7ReWOkmEF421XsRDqtV8qF+DZVDWu
AG7ODq1AKrZG01g/ulphQtwCl70ZDOm99sZMDQ/8IFG3Uzpzb7F5BrVj3/9WreeH
IOBKUCeLbpnUET9u5wtuSkUuIeRQgZeSW4rYX2AxnBU1/TlJdH1W889XuRK5L50s
mTmwIuiSM5OACARJUfeyo+oHUL/CO+EPuSSazTXbTOD6INRH5nIhOwOeSCNHnCci
Xol1RYE+gCCHeCRORYdaJB2MTWTmZ3kwE/wEp+8/MABmDoPjpCiTjGC1H/1Aw0gt
KJT1Tvz8y0zU9i+0oW/KD5BIaP1o08bInJAtj39Zw5Ly7qZ27/ye8WQJpYhk1ucr
DqvCExee/eCFoPSy9B4vSJqzodf7e7NK5Zw73hijfrsmVEkLlbZgCdI5xAL9bCif
ANIxe9KR+rhFouilJKLjngjLXSkcJu9tIGyI6Ay2hQqgf2iicUT0xPNrKIrU55u3
U3biWUCjQDLDnQdQNoNruyFJWtokOX7P2Wz+y4oAbc/lOYxJEzWeNUj7vEUFOAHo
KyF8C4tC0p2IjJN5l4gE/NOnKPuVzupQkHP9w3ly6kn2Ze6MQ+2PG7ADazLHibrK
mPBoLzCESHWeSblIBl2gy6oUcIp0xoYbjux4KQf1niTDopCUcAHH4+FrywOXxPlO
Le3egqFrpkY7zH07IttU91nZ9X5A60bNO5cARYQL5Tl20/VpD/IhbB6nvKNwnnsQ
9wI3gctBHIVTCeWinH/kzaA4vt+cnuQRuVk/Lz35oQSC31LpgxkvKSiXiwaqSa2n
OyjBsDy629XTZmRStrIleONqVULIaSygNLd+71cgsg5LR5sbNu3vsYJQYB0+cSb+
L56HtyGQx/9an1OkTEIZ49KHfik1Rjnrph1XfLZJ8DBhiQxfBeDqVhN5+3GC7E6u
Lg1E7J54eLUQ3P6q7K1rjoI8X51yBt/tmwYNegXSDC3yC32FjWCzNj0BKJVCXhOu
bClM/9XSFcZNQ/o/8LqNguo9x/SR3ff0PMF6s7NP+WUpo+ptesFEzzIKLprSDXT5
PGQjauLuC+8TlQvk44OJ7xCKppCKH3sr2Lj7oinuH2OnZzdK8OGIdxxvmgSswDji
14GDFB7KoJRxli+VxA0Dpwtu5yDCxv1BOdblKv630cgfigVt0YAIycn96Giew17+
t6q3Z0a/o5o6j4vncdUsWZ2pXvBRuJVBJS9RPXfVfvBjisT3Xr+sEaKoseNFNCM9
3HCzxme2LY5HJMXKYwWWdAm0p3LfpjiwL8K8E9CjnK0l7o3CGRkyI700rlxPGl3G
/CLQOBThm7VDVeGhQJLc6NKenK1OMpG8JJ3eLoPHzuI/bcpkq5OvRyjkPatSQUiP
3TYUzPzdUPTz+WlUwTPWgaSKUZQgwAPvKGQ6O3RG/LIMlK2hbjoWyYNL464Fhal1
SLbUmeikcZymQqweKijAxZWbrKGtENFh507QdnUu27TcRZckMrTncEcJ+Q5U41KI
OGtYb8IDC4Pk0b3Hg1AfoNoCJSimTAPEo8u/Ooawu8RmjOLuAoO1VI3c2et13VLr
mqoZe+eV/95KE/wCQdS5wCYkzsuTnF6gSZwIjIFXHdztOGY/0rbrY8SI5LBjuxfG
pqNhiWFm4egzbfcZ67W2gtwzhjSPf5/q74t3kncfe9hW+RxWS8V6cXYW+hL34ens
yPqS8Bjgb2ZQfgIqamtfrQIcHXH8kGh9KWM0sHNug3lDbwIE03+RlGx/vtBoDHcH
llkg7qnzNl/CuxFeBlNq/1ZU+mvpoUTpqXmAR7sigCGgVx2g2BEKjvaO80ZCa0BW
H+B6QPRy2OEKeyaL6OzgMHdNwF/+rbYWDXhDjfia1HeVYbsD1TVZEu2qeFu5p88c
zeDpUYtZoiffcmK1f30x8+uPffB2i5WF4ihdfbE+Wz/i1OcAAQYAnz8OlSQ4o0PT
75409QW2/udypF4sgHc3N5OwoQfOryFeb8kUWWVU/Ksu9/nDIBTqYO1+1J9ysE27
dfK7D8eXWvY5nH7abqfaBEqcHFQatxOK/fQhgDxk7IrTrkkcvxXBhM8Au9BxhTke
kpX7NsprHHHWjcoYh7Ky4iZ13tygkgWjxmQvDJTvYpaUgBV0mWjRZMMqI4mgUm1u
1ZXhNUpCCtGZa1kkI1DaqK3yhN/XndUtFHG0TOOUEDy8LWCKiT+6YkF9LwfE6ZZe
umGZqKshLLzKz66SGpvEb5NtGBxr7Qt1VfMyI31FIGQe/5HeY7lmMN3j784iur3M
nTCjQtfX6pFdSloEcRCl0S0CTQ6DJ6S5kbFaBKME5tk4bJd4GlnzNchPV1pocVdQ
BTvgfUEIIwLw+2hcM1NeOk89RagmtRnphElLJfudxHVcjd8B0USinZl59q5kghhz
7JU5as1C4jDue4NVpVtrk9mLDqVlI/2csQ35Uapa5bfwWHYfEvXK9O6QvQhTorB9
iG8hMVfYSp4Zyy5imHLJqc7iAM7tgdQlupB3yjEiSHDGe/LUH7yBEQtdloMo7O5u
asmnuUYz7cmllRgfFjSO+52fnGUj+M/hAF9W3aoEss/2K2/L6EZHMfT8cGV2vmfs
7mkUHqpGEfX1WcGheaKKq1JW3FF8ByMFg0xWP6u51TEN2h0L6FcIQf68582RPwSI
6DW/38PwpFBS4+5PzgNOptbw7bTnEvF9CupWXVFjNJMEjgy85U2F8XHhc1JwZNXm
i/cWPpN28LZnsDCET64RIRsSlCDD41NlM5SisH0QalYYkFUlG16Ov6Mz/7iCIeBa
7PVQfcQimvZgZapBPNB2AwoFv+XZO9m6V/RItQkXrOXQPZBc9NfmvXgSoazKLeo+
Kd5XOATYRYRWEE/geLkS33CrwZjPqLLDag6C9JxrC6Zr5vE3BfEyWsZyBA5eR7Zy
Fh/BTxiP+TKezrDKmpye5BPhmKcSmCYatDZZAjtxxtRcSSRN1yQDgRJjkdqrPNZ4
VGfve4R8j/QQmspRxoYH0HlaK+Kl82BSfTL2q3qdA15BUeyKNu18b8EUnj+8WbeQ
/ASvzKMfFGA/UMMwQ9eEXjkx74MbCa2b6nwMFwjQKB2PNQpj5qkY5SfSBJx5YaWw
zxg+xdavwgSBlPLplXZl4K0xQqfMxfjsxy1jZJxEo10dCcVrJM4eio0tTlcfeROD
iUbJuGr//zJrq89Vf02mUc453kYmP53Au7xhLcdBI2wSMc2yVzJzuuxepA8YgVVw
kNYSAaEhTmLiB7tDwAHIMtrd13eNsIT8iMtLEyZ2Ee7D8P0SkbVALNYG63bNRANA
0z/6O14LzzIR0icSZq5XNmHcLgwBWrCVszOmj8Ngr0priuPMn6o+kNOHwEqiqEmU
LY5vGngBeO6/g0uWZInDhIswhciYpEBUC5YD2dqX03QTj4E7ySHxAPudhoUXKbL1
XRJCtniQ5VXjGY5DbAmfI5hD9SacdNpQB997CqMeXhzE6m7mpqTlwZiXULcrTJrY
LiE4YXX4IiQ7cqd0DAv9VFZA40OGahwEjiL/+xNuX6XHtaSYW8WFK1VWJTF0FVZv
laJ6cMagV3PJG7x6XsGDQHRS0yA1RL1bfM6uu5cwF+P9vYwP8CmPrnxpREBvIIr0
mFl2RpEVLazxsfmH9owEMZ8cSdOv9gsxgGkvMVKKaM/sreKjezjjd+SGKtHFxRGO
bilOUIhtEkskuBPZNSkLaxKlzPhqXwlRMLDhb69Mcgr4zErE/8UJqMlBmm3THx8f
L66WiPu5BuVFj6zQ8LrRIFCBdRCBsOg+zyYhRs8McOIQJh5CdqrZ8RR7mBlgMtAR
eww8V0/EwcHJexGJYMC7x00Rm1b0eHGZU2anIvPr3TDTmAP+WUhJ+Jqvjey1HBCR
IvhksMw6EfKhpWiuNhyT9XRgeABd8QxgaI4Wcp18/uoN0NF4mOzKtxDUh0vJpLYc
qZZYIJOwKHH1BRnKPz5gN3WWmFKPCDIjrFvZ47rCvhaNxYh6qhTQ1mKdWOqhnwNd
5Dq2g55DDOBNUH8r5dvgUAZIhitpe3K2oK12Xorjwi4GGVVXLACoxkwZB5VVz70H
JfnAhiH47If3BAKtjG7AcP0o1ujFqluwtEOemL9km+jzy2RG473sBFzdf67HH9sI
ceeAW9Tq6a/zaYG4MRkRt9TLlstprFNFEHVA+WNF8+N6FgpwpuatMfo4TDReqU/5
3j205CTWpK9UWxNy5bKCkZZmFJdD3Rl+PNLedN1p5jWb7c4hBOc54gPF51lsvJHf
zh9b02KaJuxnrEWmN9EI+//mriQUx3v3XxkYzhZV4vCLk1voE5bObsUe/gQnDP5n
dE76rqgQ5zEhWT4fxMTblWiSeQLurLcNrLOb0B78xmKAVZwu6Lal8CXmtg3x5D1I
KbxZnJHfFBdhZvIXQo7hlQ+dn2xZdOnyuHBORui0DDde/+XTBX5VCEWjSaQogQnK
njZFulhlT41CoT1xPWgJrBuPNi+2j7OuHY12GzNvNwmlubWi0M3ZXchjoBqH0AHx
ChgIkcsKTPRmHITIVm0mWKYS7uK2/iHpwHTgDpSU8aThfugmDKpgumlT6b+mkFJC
2obvgGPrPdAQ+hMeG4IxAHGmi3rpR2pk8tOH9pg8SZRIWKTd2D53yfaMCxFz9Kbt
GsoI7kM2kjZe0LDMXzQtWjwsnAvKIVAX/0TSE2GdEKNVgCaaogItSZ00x8dwArNL
UM41+dBV2Ci+kpTb6/hK5OsHBASoGkWHFSQa8C+B2jw94Wh/YnK8sI7qnLN2A/nC
NLlxnFqF6qNseQ3pUdBiKLJK+hy611fk941MseU1puN6zZgFD+kjbtBz1p88JCUQ
N8TXdf6aqCW/xLpS8CBQ4Njf3JluzhBuenPur749rHqss70pkbE+IUzZsBHpmtEv
wKTDHGnQFwXo7ooPJRkBHy5cb6D/aNnJpWSmskRzpHO0LYJZLkU9RBRTV/2WQ4KX
efrDLGfBnV2QiCLE/BfGZ+5DVPJiXIBWUdDXqCwFhA6I+GndJzj2ppYcyNcENpOB
FwX7lozkX7MIUdIeXfz+CH9c204xwVyE1g/zVRjjuWctBEmFHxPdt8JObuB+SHFL
YkwJSBQhbwhRoWuty9LjPexRoE7E4Nsp9OtSDDssPdb74cfjPXT7LGHUGIufg7bY
Bm940M8jMNGlHfVbO6aRuF2M9dBxCerLiIHNCouU1UMVSKeQsXH98RQAf3Vvdmhy
upmkDBAzp08n1m4CzLnmZo9iBuwyagXGjS55eglqFEhDFGiNGPlxr5OQ9pvwap27
ip96ojfagHQ1ccOlktT5TBrAnb+sw61xI6tjWgVhnPXfSklLKbZ9GV/w1h3fplNx
Cl+iKjp4UrtLlIq6hdFlgQD8ox5sUHXV+iZkPDiQOQ/Fes/N31nKian+obTDg/wl
4I46E2lX7OVyXJ82QU8Scp6KD31QRbqpBFR6MXw+rgcrg+d0AQ4ArEIBbQny8rmW
NPokVdZie5t5wcDIg7TwkRCmvOrd0wcgC6oFbgN2sZZqvE71DfrFtarnNd/bXNfn
qUlThn20tJU3ggf34I1xws8OaYcFo5S85bhGB+B+z0LioXkI6XLWt1yzfXRgMjf6
uP185QrSlIEEWYt6mf93kO3Kl//PhEPE47I2R2+Dt9U0ULx3C2c8Ccs9W7j5jQB2
x183RQJPjSkZRW6jgV1KU/ih39dk48QBM4PZFZvbS9yzFcih3SsjvdfS5VIHNSH/
6pWUyLHkwfRxlwZ9HzZpaaQclJpQ8pmROeuocVaF4PN9te4vVrRp+YiIfoc0pjbu
r4tCnWuyeDnLBa/onxoJyCdl4buVmYaO15+upAOh7L6/L1TU5De7zWYx/b7gjAdo
nzt387mWnPg9rRVD/BikbeZfK/AYd62CxybOQxHqA4d1jy4jeLa5TllVqGIzA7G8
lb4R4YVBIP+RYt/ul+d3xuOJPZjFQF6uH1+CYBL6/qYS10yZuWNeVwfofMLzuJDO
32osgxp+/jK8/ZQNCakvsDSldYsDIdHwbvUTWXY0HdA+EnpG8zcoNfDeW0BMDK75
08oR9LsL2HoCxJ+B5v6GCEI2RG0qGthgbXnjCHkpROW+4OAPBVPhuDiwsFeQwdnF
cipJbME1Ru2m7uqvJGCocY/Z3eUOrKKuwalGx7P2EIdXrLtTLphxvT8Jo6u5D2p9
OUFRbOAmYCMAlCL93G9ByaVlaR/fAB+FNhewn/JWeIjHdy1IGsTDTzCg6jy+bceG
ciAsaaOxE+VpvHXtIyYT0foT+fdvzvfyP2xmW/j3YYwpulVyJC4jOjqxAiQF+MPn
8EZv85/DKeBOF6o99ywOwkOxIhagMapi/T4XZGkGWiVUMhEXZX4aig6CTlCy5BTY
wnpA+E1MctfmmLn4yJATaHlVQJkQHP36nc+fd3kCuSPEVgUszpHbRsnJLNEjX6ke
34Ad8yywvD9Mk/Ck7xjyzAw3N7QelShL4/Z2ZIF/Tr6wci543k7dXnx396m1S9mQ
JqVu7gfTz0hYsmG7AQqi9KQampFtKgxByQAVshy0NElngElLql5tMGbd7jua3uaj
yEZA8EZwntRSg7o9lYo9xWVo5TgNFrokPCwkj5Vp/wzo8L4Aa2Q41LcyAimD2gK+
if5/dbZ8xPE0zielEum31tv1tBtlLMYvUbjdnoOChJI7iJ07/4VW0b4Kli/l4Nlh
Yk6yv6o8YBV0exY43Mt3ILQZQ+xnqotpDOsc1WEn/jVuN4pPG8yzbcFvl/aW1FRM
2093fMDYQd3fVcfchQ5XJud+bN0DXBrXhxr2CKctlTFQulBOlTdSP3rN1Mx/7Q02
cCGWn130oRyIN9acCUqwyZbV6HGIkSrRpXcknc3liw/zIIcxTreaYzjmKaiaIkel
hOydC8pQAfH6lrKTZlbw63v5PNpcAvzdJkq/cqzNkJ5ZwTXRN9JnWImJqntYDTsC
2X1vhEZ9r7Zvpn+dSgCeAShjTrTquWP6GmwmLRx2Jl6pRQb70mh6QtW/Al2px6XN
YQAx6/wnwKZQmB8ucr9Bctc7YemviBGiPOIrt20pZPWAvpm4G/7c/zSVFM9iD4Kh
ibVhRRy9KNy0LaKvpPBoFjmRlBfIdO/y3a995U7n8bqAzt45ZywoJdY07yLchEmD
OjcVdxHYCx7aD4BRIH4a5rNWlI5M+lTI4ZOAd0RNPGKnEoWmL8bjCQAFPJ5mqoF2
6EQm7LLzmeyq/yyfIvA4bFstk219l4X+XkfB8MMP1ysmH8BXT3bV4uGY71LolgBn
m8vglgc4N7hSBIkTu8I3xKoq2FVv0rqUdmcJR92SsJy8Na+iOiz3O/dXGWRYcGZh
s4pmwIpp5HO3u+5wziI8ZLfVxeU0jKQ9tXhaV7qoIYe94teXLbnEYZCUDxuIY4pn
ndjZlQfbOBxZoxUgGaj0nuCjltacXYknWRIt/MRhPXKJzIj3nsAzr0UPeeQj3i/A
pEoNDHFscPrJ/txNz4vfCJn0rBPTtUkorZRmB+NJ2u6kffSw9JOtczuku4S5hoWl
soDv+Zmi+5Ztjo3KMcsHLFn15r1ordO3X3GCKaOUoec7bIZGK6dxK+1MUXwnQ8lI
H+z4bsGcYagfpjrVyUUs9D8/dDBdXrAr0xT8Ay8658YlJDQPExqpD91uMRgItJOe
2soTS+45Njfdawm4iDx1VC6dcbm13qfgMIP6pb7k5EZCSrykPRFp5SpYYKDACTDO
foaXlO0Nl/SxORD6d6Rf4kP0mdlWAne00rm9RLZyGPC5ohlZtHsP6g0l7WalhXh/
SB66ZXEFelU9rNNiirAIA8VJE5siB4QFXFGgWqKVwtKwEMFTjrWHSkYhVrA/vV3C
XEweqIkrG/ifdgh6BxBGH0eJN0vJgspvDJtNALUjkOrSaJIeYi6fwe5ZY/GBwek7
of+C0W4mg4Rx9NJfRu/xh3W1AALzhuY8eCh5iA/Nk80IOh/FRy+b3+SaFmXd54XA
e1MrKNUGA3NVaCsRkm+yin3CyK+ZvX5+AYNgHrdVvZ0J6P2ZIbF/WqJD8d+XM0Ne
sNCgOrqBE4hucBS10gZxCgpa9Nk7ZPFOu1UHUlbPJx+X99fodOtHVGQia72v4SzH
mjvzFDObSMrkvE2VSQx0Qo544/wHyR21NcqU0inLZUq0wZBu66VX1sbrBu1gG4CF
qM+3VoAd4quwb3oTLQjeMrgYIr3d7G2L3ArDsZRfvxuq2JxSIU24F5WH8FUEdJ7K
i/0ZUFj01asqmNMH8s2bYdqOO4FaAk5WmdMHkPkA7DznThDQE+mNGFOdlZfSMe43
AepfRXoSAhDg40oQu8CTOw1yVcXxYFU+0mGQ1pK0mrRxNg5hpADDYRwRerUpXVbu
JhOoao7MQc97hQ2dzqpdbIZ5cE9P/x/NBCDV89EngPaRkL7mx5KGaaOKh1gjmYY2
QwSBgsOnieBkSwNkt7IPsREWXOjhHeaNxAEDD7k7yhc0ngGDK+HRjGiJ+4ALIgHl
Mj4pXP3+xhg1X8A09X77+8F0vwnk/42W0WMY+6r0La1SmrrJ0f/ZHS9t1dA9GaHy
dpWGN5ii8jdXMdAQcpsQjddbM+3kIyjn71oQE8kQzy87znPyfDsumZtlI32fgtN6
j9j36bT/f94brzHNQv1iwJyvxfLQ9sqjbQa417CLZxz8KtI5DOOHw1PLGeeSf6Gt
WqElkPGHTZCt2MVXedr5ngSCK/IJKnr08ZcipmxulYTTl6rdsC85Uz/rkGIuJc9g
rByGOpF0jc+TCaYTpCk4sDY7q0hR1KscnqbvgKa8s4o8pHh2/nZB7U/8ZYRmoJdL
AC4hDNhNtzRzPVLI2x0IdL7pX82HAQjtsAN+Eo2AgsZgMAPHVZHKwnaPPkbMelwh
EbhvYaknWUq7YTMKFh6ClnpFHchcR9rhquSDGoiv23X5cIA0DdbZ+Ipn5Y4mL5yj
xMab8Gx1Q+uMtQ0lhsUaKxjygdlQW7qPIopMcFF7IND2/vLr6FcMMGiVRglbP9Ek
PoPTUpTnzk8hJLXVSQsVz6JqTmxVIMXCTSCo5kgTmmesOvSEF2iPGoLd813gXWBE
VbErjsp00pcSkc8na7WTOdrC52q9Jo8h/fvFhd3rh77TISzxRys8jKoopzrml4Lp
hrxZeNDzh/9QqNNbnF92sqV1vOHz8g8++C6Mphq+CYZC/3mV3qKOSNbh+MnyfaOc
OwCw0HgtXH4EHB3YNLt6S4fYr3B3KFcKu+wcdWx4JNJKEUs4+swtbnY/rJuIbkl/
KOEjScJ4Ad+EmlX/Omgd8Ps5wbnc40FsqEVZHCtZLHNL3hywbhSaM45b0rx/vAvd
tjkL2b2mEA+2zIb60ipXxkyQDHdPl+vnRrasnUJDHknWW7BhzSLqnI/okDHRomG0
toIjWO2v8RVEi2gdYDdMGIhoRAyIs9TljBJ4Q5K8xkctrmaTFWpawoUDHRAKTlQD
pR/uPZ8R22QOdqlFxm7F7muknVRJWFqxSEBmmzw1ZCNpvGGk2REN6Y2iwhS5k/I0
jBZHwFZv8YJn18l3oDBZfGk3fgYgpk4DvbB7IFZU7Z8Xjkzf3EZQTNVjrtPewxx0
zvyGGYzR5/iEziSp7ZybfA3E3KR9pc3RjXlWx2La4Dx50BXZf4jAsuApM09ZPQTs
hr3JPb19KyKCu5zGTBXO2Pn7FDQdIqBlJCOULhSTNmfWE+lSkzu/ZxF8z5rU/+Ej
IeZZYwTPCQJD0ByPCE5sI/kAKimDCWUig1H0TAS8qXAYSQGxfPdb0dg6EdzWJYgV
15UZIDVejF+uuzmJhusUa3F8foR0z+8yZli/1TVRIBPf0pyK4MFhw2JPhyUnCnoy
XkFfUBBF4tsfuqZmLvxWfxqphxcfZfVd7x5VbXjzzH3JaJ7mxqPZG+3t8C+ZJILz
f4RLny66v+hSPKC5fKUekzgEj+H/laazHqQ71aHQcOLqDKdCRunSG2qhdAJLz1lX
F1LfR/E4Ks1REOXlgGRJaJLqI/0ybkZi10BdLrf1kHrKw2oPfPHT73p+wf1hdDoe
yeizvb4Ol24AyWHAw+c5JR+v2BuQwifNXdC629BxZgn6XsW40bSGUo42dsSYLG6k
MuoLw83Hvd1DIf6BZ0H+qlJ+aSQ2l50hiQovzsYouonFs6zzc6Zsw3dT7V/E6ApX
2SC/mG9vFV+BHt4ECX9hrDx2Ju9jtw1rouK3myNQUEPTEduhq/a0utuwm/jGMXoB
7h+DOrNyrPSFfSVLcLOjctCWuN2CguocmMMKfTygcHvedoL8ILvKSJMe9YktBZ5u
WRdWkCyLFDmHfVHaGSPt/JBMoXC7hDWOpaRsYYpeHejkSApb0KRzBHQWSa/LJOrI
HdNoVC80bA6WxwbTu3wbDOyZQU+OQEolezkJBMZ27ND++DssRddJZojQ5YRJ+Vw2
5csjTvk+6ibgbXs2QQsoBsyETb2rCtTboopck6RtxFDduizm9pALpk7Fqv0/aydj
5rpetG2Sq9epLSeHxuK0n/1SVuVWgXrThQUsxfRCl0kDjP+EvnZ4XcixJvNGQqzA
rfj9V+Uv9zKT2B5KfZ1oCOf3IjDEqDA9RbBWAd6uU6eVqetPTE9Lxa9muHERBc9w
RUEfZkdCcu29vGITDaseAcrsVuidcFX3APjRKT91dd261IF82YG6TzzGnUnPzDGw
OgnI5kdE3ICuc1jmjiei7Ln+0gOcyp0NanFdOu9Z8UuRuryyWt9WkPQHwNcRUhqO
Zj4sM7ZM14bttpOvkf2O9gbd/gZR6rADOHcJduYznN2fGeEiFOrd7JCD/Ca7F7/+
NhuCx4Z2CCegg+cFM64iDD/lA9rDhILq+Limy8AVG2WPTeS18ga9pwjYO6KyPz5H
J1jcIlSqC2mTatMMc5ekfpcTjqdUCaXt03+MEN2mQSf4UDr8BlrJD9jUsIrMLdZy
aK+xGUtG+6kySx1G1NOtNMXkBmCFS0ZreQVIxP98q9iADAX4W7dsKMUjK13sHw1W
KTt72AtV9gdEfz3JVO4qksuaLeUeAIVkfqVViu8jwvM668uVAum7dfpBDa6HXZaz
NYHx3rsHFoAv/4FI4qHjKdNLGIeprfM5Q+GVxCe1bdRZbCmS2XzVUV3PPZ8XjHFC
KlVQawPZzNt6wyHjb/cEOIysaVxvBJXvrF46ZQgYKqk2XXOhLf3HQMM3vpbxN84S
mhUh76mCoLqHATWBqtuVbZCnWnfUuFATIIsdWB/4S68ayyedk3tZtnFK3nPZyswh
8mzV00ER14FigkGcfoygXbjjsHzuwogThJe2MtBieEUU37p908MiyFMA1W/B37fQ
2aIB+C9CDfQyOUSC61nQ7R8OUL+hZCCl+fCN3SXyAJ6ebtc99etH9P4f7CnV5jkn
RSOTY07hnNGUxC67N9/IhL9tHNuVyyZ860yFJv9r+VtK4HaWLE9iH8xdwTdMUjCx
mlRVNshgVwaSimjzOy+Tonkr7irFdrACoO8pBEfBCTpOc/djSk7llWbWqoveeWvs
ZBIW2BA2ChgbPwm38bGF/CjBPkSWIwDTlOIE/Q3BpjwZ6uHcrIw/3Wg+UEsvHNpp
/DtrfniL8Eta4ptLA3fjVgD2RKgtvZc4+PdcO4Dyru8pcR1rGLVPT5wFw7I/rWEa
22eIcDI4g8I817l+kkMmoLuQo8VzWeAjE9hF3yqv7CAi62HUrRPilwpqG2ltzoTO
jBrgWhYeW+soUEiRO5iQQ5kCQvmzWom8Eu0CVVsIUJ4OUnY2ANW5o32Rpw53lj65
zG0pGTyho7j/jPhWf1Rdvk4nroH+6sFBSw/cwJa7JW55VNTOIFd3Z81a9eiUpFIO
7+9kagnlyUGuexFjtmdBRbMx/COpiLZzW5BlfKTR+JZTp9dQqUnaNMSzV3PVnVK6
WUIl0mDcK7c/9O/m4PXfTDJTsl7mnUBwe+xPNq4UWvR63McIeVQHEoamVob1Xq+e
IudLMh3/atAh8blq3T4YsyByCO139YSxbLhBHVIWrr3wOMNqAbaXGCrux8Osvdty
4UGKnUSCbHLDfmjnQtwQ9gCMC1oSndDA2GveNVGecmRA9jfFPsR6eTBpvTLfjkFZ
5TIJe70QxLbWCdZZID3vUhzboSoLKpTNdFKwMCFDPAjcw6APz7+ZLZm+g0V/1tlF
1pp6BCtnwN5jhkNMiAz8Ixo9VljJkZ/Q4cYnVSWjEk12pWrsAjv/A7Sf/K0IEyVI
Kcrnm8MdS0YdAQGupifnWX7Va4WR7jvZUcSVRiy3qoCuuH5uydI+orBKRg1hsaX4
xiLgCYIaU8RRHSIRXuo+j3tqjOmk0qSZlq/h90EFJ7D8DlPLWKxKckdfbiqY18vP
k2+V/htglUCe5ZjaWD9AkcrbexOwC9ZMUkKEUJ/bHq2fMt2u/JHSzAUE4XRth+Ni
u25mIVIaxiYIQMxF8cIMoUCIXzL0PaO3RBfHfxjdB4SQYx0Iu/lYeyhhnm6CSbRm
NRM3M3g8alSzpjvYuT2Xx8IXnwLk+Xxf0RjwcHeQSAH3glz0+NcJDq+FtBkljEAA
8YfX5O2iqPEgqF3jr/fUpe4dKxtZ1M2HCc/9Mtfal0aJkGzzDuuV8gDVjFousb5N
HOCUEBVTzFBL1bOlM+x/zQlxJz6/R8d8qbJFEGZimL0qwnBe8vOC/3i6YsMf83RH
AszWpMvzZ/eXH5IVRk+stSMVz1tN9Kr5YICGKw1yF13MF3TjOqugJbb9fM5sxsFD
dy9i5M8LSzxIA7So+SOnfM/egOhLbTa4f1Nd1upFZzoHuQUAdSc64IewMbfb9ahp
f3n/NMvfVhPFBgafKhLlGBLCgFLqscclS3GzFK5E67qhornskHh5YbHJD8j7zdaa
8fF4H209ub12csAX1BAoiuVLVZAzwdQtjUgRv/beNb5Ejik2cuheLoLuysQvF1/F
JypywGsubnB83+k7M8q2lyDEkE1EkRNDOBueD3kbkDpN/Ea+xOTDqv6wx3/tvu4T
xkHFJiLlzj/QOpaWKsmPivR0mxbK9En4dGQaQgXkZLadOorRC9nLS5TP9dORs9Ry
vVGa4el1WsnU8CnOMu7gi2HT2drIfGILMNPkknhzJ1ujrTTxO9TBgcBvu3X9yh8v
n+i6Hn6cREp7LWZsxczc6yy3ba4Z5NOsIIPXgeSjfs/xXGt3LEy0Ure3Xyp2DgwW
CMn/8NnTShN05KYv5+BhLgQWkmxAT16iZKH/9t6dykt9G2jVQcIvXszMSi3LUdy+
J8m3azG8F0psNVT7zowkFy7+ikA5Q1VhBqKMyLvuXkIzm8EH9u/t1PHa5VRFB3ri
qmj2wjUezilnNWj6AqVbyVrqC6AQvDWb/hkQ58HadPGCPnoiFTVTSVKFXt+r5wqX
PoOxH5RnZl+mOhKwQoeqiftDfD14V20oqAYpzRCkBfzGjejmCI0NH7DGDvlAisH0
lEda10eb0m7P442hvECWfKB9mDpri/BeSIkm4VgOJXpiPdjLU80VCQkVKPKc0kcA
l/tdqyHNPpkiHaePeWA9fSk1drPUFhF7NT+9iEiK57e/7hxY0hG1J839pvtpiRDT
Ubo2KzIy2xBrgGWEyQekkIZblo1Jrj6QqN7uSAjDj6aAx3lejxcNaXPKfFkpE8RC
xVjnwgErM55TloifNW0rlsiH1aw6t9n98qQOIhi0gn084dRxbV2c2uY0eoT0CIit
J4aMcvGrMi/rQ5zxGpxLAtOA4qtf60DyOI5YsCWa3+C0UIkzKV13nRORsWgxCVsS
kbAGO5k+HcJ/1R6kNHWN605lDl/QD01fcXCjGAWtCF0ggWlJTuaP1yFZERGtg8HH
RqfBWBqllNrwT33wwPc2/6aKz2ynF5mcSbOm+lOQK/Ft19h5ZhKTZw18wxzRGN8W
DDECv6Nydf2YQc8xoo3O5/GoisXr9e4VNYFoQj5RJdZw/vuxNNaJ5YsbMguuKBgy
Che89AfQAk71eQEvPKpF2dadZZcWYYMoRKTE+X+yCP+Q7ypzl90et//VUE0zASpa
MxPryvK+vw6gmI1T8BmYwhoUh4WFXIsr6EeRI8cMpXCi2i7jEeuUKSI+V7HlKJel
9gyKJBWIl9Vd2ullBDIFcSKR3Y3yvgGOg0r0aQzSNsCYhX+UGeitUFJqETLlwr9+
+5u/TNeDHRhc+FMmqnU/rGBIlt5sZUEsJDurhgemZaj5aUhzwjhU6h/lTX96M+f+
ka0IWT0b2aCCALql79sdiIAG4bJ+bLoC5IOj6+BnXb9uv5jA1vt4IVO1v4dH69ZA
hrHad+VTFQslcStm8hMiKI5jg3YcAtYHBHpgFbfki4vGFr+ppC/jq+LpXWJmndmJ
DWCyDpM6XtxMrASUHkVtSrnksCEUpmhmmctrcn1oJ++YOTisg9mMtFXICASiawIl
glgCviUwD/n1Y6u8O++quGM4EjGTEG9AbUCicMdRYsLo7iyiYmMy/Yt8lLcg6VMC
MyATBWI5XisEDLjmh7nOsqfmUSX9teyLhnCw8qZB2HZ70gfZorpjuMrl7B2RG8Nt
`pragma protect end_protected
