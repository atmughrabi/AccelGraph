// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KCb6GGfmR+jTzObLZiokNbDzAnsCqV6Vu/WgJZYWMEegX403tPbbIgkojbISkR4q
u1iufDLCbeOVu9JrXikP3Zexsvf9UsePeqkXeMWAxjfzxRF+sjHLLnMYvGRsckZ5
W6EEcuAT9mYrZ5fAZg2vve2gLu8GhlcXK+6DSFu1bCw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 126704)
GiOc10/I5v/IiFyHP4bg9Um+NTk7hVwWXQ3Gc1wgGi02vJNeki2+Y+ZfuEvD6X7e
XHlyNdzgnyz/LlMQT5pMxq4mMNTxkQKftKcHbP5Dbfchpl+sgJCXxuIVbkTxsEpu
Pj3LJcncYsurlwlaLX7pO7wYj5RpLVcVQmsIGRueQydHlTCiHlq2Mo2iRKYz23Fo
SYlpAp6Wp3udVSGSAx8joNmkt/v8nZAcwsKit2fD/jSfcudDlgriK5T66HTksLX2
THsrBuhGwWH2r0YWVsUjRqXIerjtBxWxy5v6Cy3YCnFH5aderfh1gCGXgHxPgcsR
K0cQttAxhC9fClW/ZqakqLFPuAOIwBEbVeet6LmnPsPX8Dj8k446ojkFcOsUOUxR
mtZkKI0KWvJn+Eqyal+kXshyEM/dHA/njLBSq3usJ2SIwwy28S9DrA6yqEa/pB87
E6SJK/WJT5DHCV5+Z3fFG6Y8JTzhvW3eqcz1B172gYTVOYe3jkIZDVcFkvTsG4g5
BZdgBRdLcTOWQW8G2Cs4yy9yZ836zTmfoCdzRDAU7EdMLDkpX8V2NjjSxeN7SxTW
eQhibWbSSqYFZYHW1qKVu2Z4I2yiM3sAUr3Vuora62lKGu4dn0GFhfGjsRGRBdfV
WTADtiPKmzzvdfZ4i/pHbZCtmgVxjcaj9qUni+UfNzWDxCgzEL6OEgNK+NmWPZHC
IKfJQ/L2dg1FWlT7/+9FWrwFTp0YQ9WE5q5IjUBYl4VOMj6C+lAAZe3XsOIkXBez
/gksol/r3W/mc+oR+WmQbe+dpZ5/jnVN//AyO+aGM/3h3v+2isiyE7hTsbo5KnX8
Qay2h8rMDuvHX9048IYA9J4Gw7uzG7tmLFent90UvS6QALPj2DPopDi2+xMPuBNG
UBdapOGmTwsoTMfcDsXhme4qEJQerVjRorCjuQtpQnPxWgavyzc5KjME7enMu34O
cDtOknfvGOueTffJYkwxaor71G0GBGeJlgCJ7ZbCzlnCWq/JL03Hyn3hanWfnFpB
NsE0evs3mVjMHG7pc9e/3OWllbi4p5a5m/EMk2QqWQoLZ1mP5XU7bpz0rh7xsejX
4vYoD5ypDckQCTRQQJ0MsnjDBMoNVxZXcJX5wlviJxuPFkX6tg5iZU/HFeSoQX0K
RvGqjtmLTMHNYl4sbsYPd5wnpHsTn9yTQvYJbKBKWR1ncsfEucInwexLkw8AVKos
1sNMzY3ycisjPBB0syeRZa+txMMzOfQfQPVJqsDtCFqFtmnXsZDyUFf3M+jnTZ1Q
k1Iw6QVoV2efc7xk2dIYJKR9pdby5al2SmWBNNjQU6IfnzIiYDnbXpAadd6ZNtjr
0cuuyvgOa7lo+PPMJ1bLij2y4wjOrA64qLRzeY7+Yo1qppP+5fN4rD0skX0O+kWc
PqgarrFYm6MmjiSyR4IHI7H6FRTVWsoEe36SiGmv0Np0R6J0KruSDT6CMA9NwXy7
0Gvh5eW+pJaxOb0EmYtPD1FVpubFUjbV6vh60zq99GubFJdTqXBbE1Yz+cp1ZB4p
XrkbkTL+rUfxNTlqB0an/VSJQwjQYr1qfUgwWhLWYVUqyp//4SDjLLC4W8sTX3hB
5H9dQMfKHYa1IaZaRLz9FC5biYBc0AwATKABXx5oNn79JuTj1110YoCJwIklxXyd
XFr1h5eIbRz41YlsBBbXUDwHuK8UrHeZN8v6uXdLRKQfO7jAumwmgo+v0fRXiYs6
3iuMpc5YHyLvAHQDAxWyDCbFIGS1jUgaBkapuHf51a+VsAcnMvKNbBzTXdkWapUF
IvuenxwLw2if8Fb1gHQmpmytZ0GgScdZ0jTBvh3WSOK7W34rCGLEfEfNhTFArEER
GyrfTDZ/XapvUwE3JG3dU6nrv7ZXa2XWXo49+wm80yKp/JVCmJ0C7xQYhY+df23b
EJn0rZuR0qpQT4P7C+Oe3mI/pf56rl+XX5Je2GGSuRo3TAV0qDlUziIVew97gJPH
3y1V5ylYugPpTx/dkdkvYtGfaFb7h59fD5AvDy1eWJoHR0TlENp4ha0oeM2Qc56I
o3iNR3JI93W7aCr3YakbX5jgDxhwzz1gBBAMUyjXOpYgPdXC1Gb0/zwqFNv7cvfK
K0MLkgxrYhiuxBeDrVUDZMnmpfuJhiyBoURjmFhBIQPRhH3T91c0nUTlvkqCVWe9
TEqmWQuGovSf+dOR/ZA4gXb3uO9fh+K5cgLty9w485WGkBTZ/Ey2JqJiGZYa8vWD
7U9PzmN3yrF0vbrA0+HGAoJPnY6f7ikQ6CaCSV/TK3SoZydbCdH50bTisyMFLAec
MlPqplPhvI84Y0D48Pjp2S+aYyU1H/dXblsAR/1upXisq3Ag641IxWiGIufs14+P
bw5Ve9oETOPq3FejAJDKFVQfdsGnOwWJkVIkuF1m7hfadnyyJZyunvDXTUZIUzzi
M1zEgkl8lO4AEwX7FZwnBqMD6iiJsi2e8NRBVlxjHqn3rNlzh8doi/BisOcAo6XN
FAOOPWKckkrK9brOGhY49jbEXZTpuhhvGyUjKN02O5SPIne5es2w/yEA/6vc0zAO
cyz6zDKD11IWok2x6H75bVKiZIvQ16/tq2Ati7rF422fSj5DlF82Dgwz7CxEqLuS
YU5rbrTOP3YN4/QuvNZeTvgOT2y3ocRiIsmk/lbCVvOwc7P8AjLStHa8atxdcktv
hofIUJs1kSskOe1oyZsuS8B3LTs2eQW9f8Bkn8kXe6MWh/w5SXwourPNH3+nnpKs
i4SAne3t2b6gHEEBDcR+K5ntoqpuZlBKIleP/00r5+sSBKMNcHARRuD5GyxNrBal
HJO3ZDgSqQkjN5BvnK5VPoShulqjAyU9niuv7iTMxUr3hCyfFBMl0sknIJXcGdJq
eXD3hxC7kim4SrC5OsearzLk6y3vDFDVe9VHZoG4t+HDXa0TavR7PkCQGU5dopb6
M3NhOP/RyREMUg92peEuXwxhRYSk5lrOM3HbHn11jhaXVgs4QtypIoli1M+PS586
jJnaBpToHJvgJPaaIvEtJjteGe6PgQGelqW4SqVgGCpgji79y2+quzU2hd8Ab1gQ
qXzwLC+T61na4IQJLvrjirWagLq5N+o9yUJFJB8xeyZooMWeovBZcBol3GHHkYmf
Zvv2Z1wfFCXBsjDVy0ti1AOnpccpObzKRpQIwpEVNQYw3b2vo5ouNyJJAdIH6upG
mGPJKsPF+f7U4dSF8pSydmocx8WPZjggM1zQFf2LrwTX9mfGjBBSjUsIg3E0YrWz
+4tk5gyna7CCZJO7X9S83ko7O9wqHbCc3SsFNgNqBaiiMK097Tb8U4om3PwI0mas
rklGv3H33eF6fQR9tkoshz3totXrpt+L7M5x6Vz0tvpgcf7UamsvGNU+MaY2ZhbO
CNvFDkAsiSvd5k0qu+GLFdI9AUinzNfH8M4DcSPBM/4tCwagRx0GZpkBSxTpuizF
qZ/NERTZhagMRYWA9AkW6PmPs84FlXVHEVQF2tMUmqXclOyprW5O0WMkuSsyUPdn
zBIYoYjdwngq1LEu7IaiCHUkLm8cef0rKdKPKsg7FX2YcFbbByQADT6P/fbDyNd5
QD4q2/svN3fOeGrB1TfrEMxRl+2HowclUK3YdUp04q1uWtCu3OnWiQAQ+vsUnI0Y
Vu1KCnD3uVuoh6KJeX/Bgnp98aVRspZegknOG3gErQ8yP++LFTuihdP7kf5mHu7D
6BaLPXGfCG7/44gxbN07UTmEXzuvi2PIXKMmZ4CWq5b8Iy3rAMS1iy5xI2cFp3h7
0alb61pZp7/AEgzYKTR2xivC72vwyaoO8+gW1QMUMwz+yR935s2M6SWWgq3W1FUg
UUbtaoeCiM7SjzJkoPTok7ZA0AGfa2VolrK0TKlAgv0O2eX3BArjeXaJjkCNXXei
plTyX1Vx6QA3h0j2COAQu27kVFwBhqp3MEewMiFTxz/ufORKrKSmZObadF8SN1ua
ZXiiA5ZRO1i0e7lOIv7rDCcuxE52vYqH68gZ782mym+5dEpPY67z3hOtIdPaSbe4
CpFQ3AwmQ4IPBUXBK6HR45ujjxTIZ0jqWFI9S4y1Ayj5WizM2hZRaICF1EOxjMox
gLrqSujLIK++jPme+zwBzMSH7i4WlO/WlKdl1bsNA2rJ4LnJwY0Er4mtS7JtBfGb
JfRiDSu9hEw/H7ZNHHiEZtrrrQO28FlZtZQO22ig7f0pDgDXK72cG/HTUydjVqbJ
s1mynx/7alE4uaLfAyeSlYBrjPkTWQs5brTzgNRhyRb0oZBXhKQqPVl7Ezw2FTQd
1Vdo0aeKGWprCEdRhBt3GHNZP13n/o6M3RUjVKMg6XmpyivNCConsvkbR5YzeEot
J6zaDatuyN9fxU1d5u2E+w6MjnKBBZWnMXUhSQn4dSfRP65yWODv03fB8pv9ZPYT
uc8qPwNG/i5/Jz7DlyjsAHT1NQ09gxH9tEz74Q3Qcak9l2vnNpo2AnNImDDNZ9OA
mBweCtoNEndpQ130eI25r7qC3mgFZ0m89asVBhKyqjNWTIWCKXtdxqdA47Imiou2
7kH2lrzkbViY/Si6IwzOhrm+x72pTXZlwIYyeZBa3YqT+FZvnBsXiibM58K9rB2q
SUlvMIqMra2nM1yOnqqJLMLjYVRbocWKvAB3vrGdMfrFlU+hjyHdPnKW49eB0ank
yIvjwJyq1kDaKqc9Z/s6igmAmMjGvVHS+3HJSQmLUM4yMxMbzLf/vCpX5DSy61WS
Mg3V6QkV3EKFntyIoKlshyQgK2hQJCBXhJ4Z6UugtKICkaV9f3lm1Jhs7PWLagmK
d0PFzbVAZ0N4iAnlmIRyaE22kgtv76CVMa6CWlGL/lWYhnNQVDUMWLtKhYHPSR+K
mFcRVc6Me1MbTYDIXzc2lGqCUD8rg7IzsgFwZ8lM4qNpA3e0WlNlOWdpntIRG2QS
aSL4JNbd5y8Zfp73VXyz7SPhPHfMa2VFJKI/cxWV+gLBBn2okOyKXmQEq8jKzkVc
mFtvPP8T5x+rZa5/sbS+HkN2UchUY5ggvfNoKMckKxIZk+DgQd8Q3RrIWClFVHLQ
ewgDBoNdHy5GGIpJjvwAGP+P7GIchNDOZU4wUWRgb6Eee9H2OlIUz9h/egZL1zI+
TidR9fjIlBLKaRIm55yc5IEJqJ4zpLU6hkfN6hXM+avVaImYgFEFSWpywCel4PkJ
+zFQEr9L0zff9Xf+Mw21uZawsA4geVBNNf+CtH+ProetN+K7rWEo8RTbd5XOepc0
yBLSpWSZeo20u+lLtiz+p9mntPEXcCnFPINw8aP8njzrMb0oMgtLqk8pzphVnIRN
gvaoC6fBkwOy6EgBK/iuGEXi0nEbJKVTphR2mxZrR4T6eDJT+wD7T0zfvVKMdOn8
TDeaZx1WfKkt7n7AgmrpWQAcsPloXgGzE0SK8uLrmyK2/v+ojMP+AWW6mwWY/YnQ
VVxGOWLdbPnzb1yLoc1j8vG5ZTVx5O9uKga6P4CR+09rvuWWi6Rkv6s3l5r7rBJL
on7yH+C1sdJAMTdnUR0WNH3WC8uPCR9o6fGURGwuVWLLx2gbgnJi/9Au3hbCBAWi
cVoDIfIvnt3fh7veaXcdqU9vJ5H72+qRiSfruAUqteWgrckfr1gJKKg1iH5/lXNw
am0c2u+kndm9iugu4OfU4ECEr8FX9tvKQmtB2w46grS/hab5T0egCrYD72Kdekd+
ODj/DBJg86ZzXwucNOAz0oFH8P9hSRv7M3WHRm2Fptf7CvtDornhbhJg2o24twpP
+8LjY4zxAsrW3smDZU7YViO+0kH8cTdQmnlXbO8apE0ACFmFvo3Sby6ak5Jr8DWX
nQ0jTcorT2ZGaPbUf4zS0GQu7schC5dRiFJOTxkaCkLPu3xgAiC2daLf0QAgqUmw
jjLRLd3tEC1X6g3fpldyoYlS0uzBqXHk+0/BZIOqT4eMX1M1KI4ZuLXuov/mDxJm
kHcPzO/950fbMUb0JLcHMVPqnj6CFpCrL4xkPZFRDNhrErw2u/RLtzzVpa8CMzhy
ERh8Kt3G1NI6KIHUGauqYLNO8figZtqGkJUd/ZyGF0nIRGGST1pYcpfo78xgjvAk
1eHx/Md1zwuzF+so4zG55EZBoH0C+hHBE+nj2no+uIVspHLgH8zMP9UyiNiLqnx1
Taxcpd2fHpV7uMjk+7Qacfma56x1cVQSwNwPm2x9Dn4fH6A1s9gHv/myagP2pPM0
9sewf78DjO/+7RNqomSrNXmQrIZY5MCwChCPNqq5qWJEjwNRY6orHoLx4fFRfCix
G+LIuA/F2evl4a5bsfRsltIlK6puQZRM/odomDjK3Di4Z1Z7VECoyBqbZkXicB4f
3Nx2dS8tGdwgwIfhtVtru3+QpVr/ve9ty9q9NjoF3GOYchl3bafvtrFToeypRvWN
DzEhkTB4P5zoM/HL+cWR3sAT6JdoTLbaki5LOwEiS5N5e25iVrsb9hBerFnZYuhN
1sH7BVShxAJzC52NYPehIx8Qtw/S+Ewe9K4WfjXvW9MkrQuwOyMTitwBgrn85i70
wDX5v0JoL296OiyXKZ5n8Do4xcoizwXQ67pUP7zj1+jvPkdCxLVcSaZmKxE1UwBw
uvrx+uqdUqzxl7TECQNeBMXXwUVjbghNDrVzY3EYSJC6w2Boc37YuI0+cY5/bYZc
OLNo7cB8TrhvIkCVMK6vWeZ1D2oWhJthOWvYdVwdqefaAGu+3f/TO0ffAQR2CxZx
PBBjS//cyIKpMIIcMzQlJ5UdjlXTlVEj18DraNWl1Ax9y24wSfWTK9trwuKBbOsN
MOmLqEYGK2oU8jextDVv4pCNBU+W/IWrQuw7qX1hHjyNnrltCZO4DiRw0b8oTFZB
4Ix57D2QXcfOLemGpSfnjk+dxkk9ZuyN0vRC/dSqaciDRO9NUfS/yFDvmi2ep5A1
pQUeY1MCyXpRcSg/5uPxFW6LbFIZeV1v5ok2pDO3EJwXCaTmFvGYBp00F7ftFhUX
Y/liR1yJSx/msrUzWo5FkdPmKhETaNrtI8XFi9sWb1RSmDu2NkJSUiixJ/n2MAEV
Ljf8vYYZgX26bIKn1DxVP1XFcLYeyXMImuZhmxjdL/MblC9yZN0lMDuevZ3uA22c
f24VdtvPoHoUET+/uEtIk4Lb91zZJbPC3lzYn1vbSbJlwmDrM65wG4KtYYaKSWjy
/M7PrDF+8xj76hdwE01Ugnos3TlEN1DjXQbbmao7pBcGB/RiNZutkOYqqnnupFW0
XNj7mSS8VrVwUR1w7qoh6+8TGDuShIBGNyhOUNXGGeiaTXGNu6lk4lvPmGytI9JZ
OV8VAKMfVZDT4arbGE8cxTrmq537/MOUk+X3LWLWsGoeJvlN5p1P4Bbn9TtMQiNz
3SbQVjpX3TAitCfOghYohb6FKtKX964e++7JDdP7WAD21OiMXb6BvIuHley4tLL0
esODkL2Cze6iQB1FJBz6m15Rn2pg/1AxTpGW28CEFKEKKRzZuHFdv37ACTQBUD7p
vVUz36zWcmyEcw/zjCjW9WstpfQ9cyf2N5/4G68ab6IvK1tc6vMkq/EA4d0AIXLL
aW/CuLzOV7oNp2dcUh08y7O0EjX0yhjH+RONqYqSs0w7gAalvSfhkw4vOCBRifcf
jn4mq/EhGnHm9v8rcZ7j3ziUipvbtSu4r6B+XOAXW2dShVXg+Dz2IF4myRWBviPi
ej3Qe/p7DVE0DBla6RjqUVFF6yTIQxMEEHffoqN2fWgyOVSCRvNtHehlxAhtlnY8
czi646YFSxpQmDNoVi2yTxf6IHEsG/oMTmbX0va/go0J8znzKZxYuvBV7PvkIuuo
dfI29/38pbWgn+LMo5sRGZHhmTWV3a7oUgTysTH7ZkqOPBAPlTyV3oMWEMx/cwwB
2hLPQkIaHKlPoBLzTy9pkfbxF0OPxEWgopWJfjuBietl9cWnNA8KmpgoCeaoGHX1
2TlyZpzTdYEL/vk3mYi9ek1mqmPbvSQX7vSPdwy19BpCTsFhnQddcrxe3F3nSXvR
3hjcpgwDTLDhqcGO7TVIjUFsP0bGNRwGz6jN0AeCQEJpVU/NVRcmFPDa7Y0bNA7Q
Y2RPzBB3DSKGM52rj5DIp3yAyQkoKPSm3DwnUrZSFfjEvroHnFjNJHVDFPzunD7t
d16vZw6DZKubwH8bcMwxH9aSYr3+keNbtaEJ5pFkQ17rBk8ZBknwRXuKbAYrtM9o
V1f4GibHkErXYlU/j1mxwSWN/l9NKdEC6YSuYTWVtPMtIah4ixZ5VdI3YPVkEsip
J4SmMfkA3Y40sTm8Msm5qn2ZFiSY4vOT1/2BWHISOy5tuMv1k7p2nMeKWxOph1R5
b+PenlrBKd8DqIs8IyZ7dxURXIGe1OsFSVUBLPb/RfkOW1hyYPYPsu6sjvNpRv1Q
5a+o8VH0qfzVFO2k0sv6XeWzepODMLCd8+X1d4gBJQ+E+t9VFFwkfmdwr0RJMyvz
r+NssV/0+mvixZ2XFl5FE2I4f3NOZRqJTxAOrAvAd/ruOeyCaPGzCo2DyF/AZjea
XE+RlLjgPvbNdP46YAjdSFGYgyiepZ5FzrnTdzXrVFHIL8fWMQcJSHg0LKvRh0QZ
1cWBUE3G6T64JmgO1g4PcRgDh1FbRxyw3Zuh0cL/MFH3RLQP/21DxuOdJYS/wngw
GiwLcttLZrINgwCl9pdgXV/NSbhlXj6aK+zi1D+Xc9zs/PUWjr2NuqYYYcohVP5b
8sCQgf5jYVGx0MskDOt5kwQ1UBNNQrqgXrdFyHq842YUutro9WDPqUGA/GoaF+fV
d7coZXhWa2oB/78Kta7gzMXc+qIO3YTFNznChh03h4Kon6w6A5IG62gR0FY0Rfj6
PuClgnstTBmSqUlTSnpMRcAAuPtKNLy/QB3Jbv6gsaCp0DTmKtmufIa+9zK9hK2s
zmxUesVgdvJz/uP2AUqxLts7zTClQe6nvvN346ZS7NzXJZABjpJ5RPAv6wwfdRLN
zpcqzSzpyYtdFjlbKyppwbMzKUNDumP4ya+YbeiSHOFYT8IGSC09lrYXLgB6IAWj
h5O1Pr3ivEeLYRbntqk7kNTAGVk9b12L4Tzu5HgT/bpgf/737Q5AgHMrD/xASa4i
o9uSeZqhEqgGC+crzkDqJsi7ENXMqI/oE7kYAC7xy0XVqmZz/50B0mYpEZZ+l+oG
9fPz6V5pFr/+pDWYJ9ym9IkCNwNclMPpXTLxx99wjIDCqN7LQKwjDkMNDlPz0WAG
M/GG/6ea5GtGotueZ982C6Rs8nfQKFyxTEUU8cfbkG0gjL7U4Jy8048zDsKMT0AN
kx/Kj4DnriOghbcRVO23piMKY2StZgaNRIbb7Zxt5/gb1uzomvyWRnmR+Ov2kX39
Wm7ajTguLX7E7j9CCCGYrNoZxUKhD+f3SXx9qg7HQpxqJlU69ZB+naK0BlDd9Gur
sTnzBLqKvWG7VVLg/hekpZ+mtrtMflzUDPJ+eg63Dsg8I2SZCEBypkCEuEN8Lj7e
zYF6p7k7hwYPkUTH1CIpAxBPfLWbK3otjIBiEQD9gX8vuJlDPzcyvB9CXMC6eZqq
xs1aomj/PnwNxLVknum2StYrnvr4fycL9bssB7P5SXo/p6ys+l6tzgJ4+hau2h7s
jkyWu3m7YrQ4Sdw6cctwwLRYBeC03eFCBzDjIRoENR6HZKbdgvhymxL/iV4ctyEH
2XZs4UjrJEc+vZgZ+K4I/TWzy/kadY/KA3aMQ628NkKPwAtpOT1d1t9sCUU0j+/Y
shd/Sf7g8/xAF0UJ28W5EvOkmYypUfUgYRa/M2qqsxJQI7FaGxegsbJUMWJMbKIz
wYOiNiktV4zQmJUea4LGWwEZ0mQ2PzH0hGg+Dm4Ax9VXXyWqwjViPrA8zSyyhpJS
OxBgV+OS/ELysKkfE1P6gGeFaNAaZNbQGlY/1LmxNYgywlguGC71DBOvmc+3gf9k
8aEEGI5COaJhI/cMiVqsWU1oQ/ldWINbyJVgE39zmanXvbONdWTj5NAGYEYpQrlQ
FCN0Nr20/vuH4KgKNE20Cnx3TctxHjitzRXp8tkNxxT7dBbWOmxilESmtr6100c2
BWy0B5ENa6GrlYDCiRTJphGROLKbDxQl3cHNnffkiOOANH31NKmf0p4BZ6qh5+b9
Qy72ubbCT9n57Y50W4Bo5DIhkeUFWQzxlS56qV0p+kvfZaz2cq9eaqkczodoMdze
QM5whXnlRErGerS/3La5i0vhTkFSIRi3wwr8uiwMdyr10L+zbO98+0umuMJbkn/1
xFByVVmYkWUYGADR19/XyJuG0v8+Ojlasin9Z1iLiQVSSty3GwBe8SW88Esg7hk5
zB2LSx3azvlB/OO2mSzR3Zpm9tfx2XxPglQ4R0C2kK/NPErKmhGpzDdUyFQmVegF
4ysN4rdkqD99TCyhXe55uwHhp4WAtmRKT8eS2eU4elPLcAUDeoG1Rlf6WZNn7EKZ
FaAX48GHRRkZiVOrFIu0pZHV7E6jcPfjmny1vO0br35fgPTF71ZejP3zZxl5vYBc
r5KbwPZYFGKT+yFGHunTkSk/MxDkMuXu+HmZN7/V3So7WnWmJRuLU+HLVbvVkA3/
jUlZ1CDaIlGs9GnhFNCX9psIp2m9E1rZNU4+BGYVfHlkOb4vnwH70grt7oaJGutp
wBAKB/d3MZ0YziNfQtXAE+RY7qC1p/KrIja2dy8cp1kv5mezwYv6+avpRTU7eYbE
P3cHm78vLsi1Lp6eDqaBBNwF1Xs04GzdBziG/uSFESToHTzwjFyJ9lSOMFcntP2o
rWnxZ/l5lcO43SOnBucNshjftBiD++nSKKr2NBH/NJNRxUz5r8HV5ydECtJf1bT4
RnKnnDa5YfIWCsaz7pE9kKKaLw/jHjELprgr+MGnOEBv5r16xEZ6QDx+Cuch1OVk
qaob6NVseX5aoKjETdmllhiGyVhIMrLqzn6YTqke5BzieLT85UfFORnzyeY0t05+
4f2qEL/1zrAJOUOXMD4urYZxOiT0J8A2iB2uJNNXfzK2JgyUmQrt5CZND47rOEOG
zgdqgzXSWHaBF/jZZRWoy+YeP0kEY8qQ3y2oZ1GHYKEqy3QMK8W5pf9l1aWYleGM
ymRbN6jKdeX0B+jNlzaRdP86O0FCyM2tW1zhwdaFx3Knzov/9LbF0sJk6XvnnDyi
TjRZEQQ/n/0NFdDAb/eza6V7ROOAu+7EC7Ff9I1SsmeiFbDNQdkVt+0kYLxcuf4v
45U+o/Yv0J2N56+4NHd2Hc947+2lrT/xIOHvNFKDh9uVe94kL80opsqH5+l0reSD
2TFqvJO4gvxgowUMr3t26NvEBHWt7f/9h0FhJ8DdhufYvTwa0OWtzyHd64lEU4OV
iYMLfUTA9+I4jvd4JiAkSZRmXe8CQH3PMl/EpBy7rFjXHDGns0n3sLOHnu8jqToi
81omaNXJIUYmcn2zZRJSyhC6CyY6zBSZOTrjfB484XBFGVowD1IjxFUOzpdF0QnE
cSMB04Qn3gjngWUJvGm8qq/yEjlzOWzuV220LyruObCT3Vb8fBxMX677IbHYClpA
u7NI37gPrCm/KZtC6gwaxDO+19YpPe6VqtPocxUWtRG8cWXuTIJHcKeAGNzy+DNF
hkzDRbFfn/c5ndKhoVf1Tkd74nTXMLWI3T73snM4B3tUUtxVMlE0flQkAr4xylbu
iN0AVjFQVINxwIoDRrINmnmgNbluXIqM7yUMSLJJKy+LtLiBcZMtHdlw828fkd9x
2Wb4Z0S4JWOxuWcQ/s72HGj/mu1HHnClRsvXfKdY6jAg0H5n5S/RGEpVPD3UU1FH
8i2Yp8HEMpC/bar8pvI12DtJbxqsZ0ZejTVoKNGwuu5NW6svnjlU0nfqMU+0ryZE
1zV2OAEZpi17SJBmR/ylzQc3Us6ddVdFByUo2AcJvS0xfJOvs8j3xs1O+nbbeDq8
agBxjMYUHAqJMIW0E9IEtZRaqBP3SMSS11EJ6yGhRs4NaiUPE5OYsN6igtq5J02v
+gKM1XdOeAP/5V0vIxNXbQ/slkWjkh9g/W9WYrFJCPln3YGoVSqtgGyG9HPLp41F
S8zc78fEXJ4mWRfn4qSgm++Yzq6dqv8za6xE1c3lU37238ukzSb/nMmaSDn4TLeV
Ao7gQuyxXYGM21HpzpzsfQ2YOdsYVV+Z6fmbBgNr2zY/9djHvg/srCQ0nKLI5zxz
DbicjgPq7TlH6V3kLLkyZ+P88z5APJhI4Z+FrgT5Awr5QohDJfGO2eEfRbihhxQy
VETxmgzN3Vmfh4mJKDyW+m2HEdEkYVmTqevYepgU9ehmyaU9ODcPqw4EXJbKTJCl
r+f/s0YGsM9SU60lI1tmLIbLcaixg5dgorSdAohpVvOhRV5COL/aZn2KijlUOh1V
jOXyI87HUHwrSAhwSFBCn+TWFdzFLvBndLqzffQhbnJdcb1C7W1cCinTU5Dcs6qW
i7wQyL17Zg/t8gpkwOLFV+2PIiy1VyOWWhcZWry7qbXK4h08aN/VDgkhkBevANlg
2lwxvU042cM4IvpsL3GjWbKiSh8AfDT3QpA2oSNiPz1IafcjP+nt6Kh95gzSEfao
5fKqarrH8Gm8Qyuo/CzUDEulouskFY/6SCCqVXZgBulOcFqhYC1cNs0wzWFMqDWg
AN/HPZosMaKbL9Im+JZUiCM9ZcurNMNNJx6MbvU4Bt23b3RlxvVFOCvZWV4cfcdP
JPBGO4zXidvKx/dgyh0L1VlquJKCzDfQFIDca+Eteva0Phbqv2iYHc0iyKQTfgvt
8OdH8PixClDVLNUSJhK20+XS9hrfkC3kXFvkTJ0vHtLYmI4dGQnWa1z5Wj7I/L3z
9jRGmUJVjsXtB42yjpopIYcIfzu6/eeqzwwUIPDgNrvwQ7soaP5/lZ1dpBwWPGR2
OU3HKUBu755rHIgo3AOk82Wd74jNn5cDp5m+APTNi4B9rMhCKrquE+n1atnhoc/+
XqIVQF4sIWlgtG+yfaf0nOQZYGv2bM2VUvJR/GVDJoxqfiyydrFMurcAIAg9RjhR
TMJkdgT6kYaof7c7jEqX32ogywY4AUji8YP22/+a5s8QQFzXBRQWsFPB9fse/uqs
DLiC0S+0YjzHKtecODg3puxtUHgnkaMV7A1DGFQBRq0deqq8mx+Lafb34kS1eNi6
c9q7eeNVAq10sjcO27dl0B0Pv2pJlyvTPq7vmeKiMxj6ufzvVQHuWPo0/sh4FUwQ
3xx6Pzj8pAkLo5KmZZ1BSDLVtsDaxmWN53EEfTX6flZIB2umhfuR9Qztc6FXD+vy
P3Q3kR4N8IDeuXYITxltgotHvo3idXbMa9xoj76p1AO+p6rHQ+yRq1X0i2//U3KV
lmOP/OKGkhSs5w//vQiq4MpesFob7X/lcTcr5IWkBcGiM5/aGa24Fpq/G2LuVfOH
YKXoi1XRg5WU9GUBYiOrRf2ly7hGSmpQNsrd5NN/AkQQ0ZGmg1Ewde3PE5oszPum
SnuMDXCU37rDd/yFgC5ZYw84f1TzH6CphExscWZeTqAMY00bmVuZ1djg68v/7K23
dRB7Z0MYY9PRcUAj9U2j/I5kDh2s/0POxsEV3nRxCnRoAM+GeQ57zU3wDwsEsQgb
4rDJ7rYeAIV+Bv1PnHWNXpIOsdSr72rhU23F0C2CHZe6HJTBpU7+6DxhaDB4C6f8
/J7k9W+KZNnD1BdUPrhpBwKGQEgf72ZYcySKcb3BsOpYbBn49AkX7v4bzS1oFHkN
HV+QuliB3aWDE4HvcJJiSJFCDrlVAScrx5g5zPoQMt8Eu4w6+ePjhazkKfYfJV60
itVk3+Y5ceOorLl56oQ64t1XzlG0xhshH8sE1McsjCOsPzvEVGXYlFHF/176Djpu
kX3JnaUD8nQWHXQYbk/ilKqHJbjpMIRWAvkntLRMgDRXR4ScIYGUu1foi5BFeHhr
qVR3eDabVFLrQPfFh5zvxFcVe2BZVpGd0YIGPRhRJz0Mmo1EPTslL1a2iolRmDkg
yoIuBAN8EwqyOomKq77I1yPU+XvqMHRwkw3SKbsXIJIT+9lLB2EqBtkTY56MnFUb
1ARN74UThEsKwpp4/+BLXhMgWNMqPkcn9JjF2oHoLiHTXGZal3tTB3IKLS/Fnq7g
NrY+8oJBqJO7FN7iZmyyFhZOskoXSep98rHKM2eM8SMreZ9/JrQGDfDADyL8gSoU
OZ7rzov+PUV/WA8DsewCO94FrJpq0u/R8Y9q9pBAVWXWV6PiCNnx8jD2kdogtoUb
W+GCDIvzcCWyLhpXA6qzK0bvZDKKMcBJbpbFNAXh6fL3KP5dKi1LnM/02tVJ3+HU
HVNfpSZMH9P/axIQuHnsw+amhocjt+oQwn2bPTd+orciJu/cUxNQNzns2mEr8Q9H
wo/11sNo1/Ooft5HXmnuU368RjwbY9Gf25/HEC19hWmMUNAZAVq0scK42gYqpoxl
kqzif7q0DMhuaeN/La0XxqfNrPvpEss602Lu9tSBDrGOxuClmlKDYokgVLbWAqF3
C4G136zCTFwUxkX5gLY/gb3rF39BL6d11+MPncviFMzXWvSFGM40KzyTqL0Q1aLV
Ln4iQ0mJcfrLpz2D8KnMNCmHGoLj5Vh1w8SA0s4zMNHf29pK/fsNMQ3jOP7k4AKX
6GQ2eIhj3tW31DNu884LYxf1t++8FpC7GqXJP+tyWGd28PTZ2QQTjxpLAnvwpyFx
kz3eIaumwqRn3DV7OMjh73hg5O3iYakuzdF8ZaW+/WN4kHigSmE2T4hGcGbolUzv
5jBDUJedM8STQtfKvurFbfCsczZ34f8BvXx1mKK3ZJIyscZ3R0AkBCNMnYcq+Mqi
rg4G0yBnPvxG6rdohA308YVrMwTyxVdUR0w4OCfjC77iGdWbzGB6nr9OQRjML2SH
8j3+XcYAi8O4CUpGYKGp6NwN+epzj2Wp6Ygu66JhcOpyi1VyxlVybebNkeJ2bfiA
rdfN8yxmiLe61xlsWhX2OCCoAohfG42fQ7soSn8Z+uI9Va82mMD5VIbRo143TWbY
G8PEQI58EVCRGCTLDJjFbWkcu4GV/NYg9Wfwstyx4l1C3fWT8OT9Txl+sYvhSh6c
ZrEPnNo/J71RVSvcfBTyWFAfrD65ZQ+MAVzSOqG9HrMv+M1FxHDXf90SKP7jdEAQ
voDAnGSXbmcRUzIvYF09884wROcVY7rLEitvMPwdQs2y4KQsMOiNiNERT8K3tU5Z
0uCiLTW5P8x96kdPZJrGrdj1naqcHZqjtjb7GzBMDnhQSHGXue4yvmlfmMRTp8rL
OqVjstUi4dHMVLeRCMbXAjTlaGPyiifQMmmk8Ldv/qs4Q/2Y5W21a9dEJ6MR0t67
QXbjIIPdx5pbPP323tNlN36r40EvU3ZfqUfrFNomxZsWLyHlcoBcE3lGigd6bCo5
pwTdlN4yDYFYbekCP+yMJ041ZGZyUpIm+tKoU/qFrNsx2zwmQp/x2pYlvc5RQDUP
olGr9KyBZwMfyws/IOaJUvfAFQ+rUkgNeyeQJ6f+dCwja9cR7+U7gq7HQj3zYxdP
GVS+YZVMFsr9qAXHQF4TOEb9K03hk5Isc4qTNTUo/uMXhP3tsbRBj7gFoP0nQLon
dv/xzsuqw+y8RYoO+zDRbjtNAx8fCFK0tJ79tMgPpJKLc7LP9ZpH8xpzJRJz+vgp
0HipUPT3Opdk2o5+reaWnWBZ9+T5MQugpldCPK42l2uG5RIQrt3tVr79I97X59Vx
S9jIJP1JBHmK0N4Wk5DcCay2Yf8fNiWLpvhSNWFDEcickYsURBKVOiI+TWPD9Pr1
jvuyTVDBsRXg9XFkPXBckizPOGbDu3udn9lRmxh2vkpsqB5TnYXxVCwJZsbKhay2
zGIp60/6vm4t/gYwQefuIY46YyzeJV5KByiWj8EsU1NCRwzAFUtsJ8gbTLLmU7eT
1yJ6Zj7s7a71FBUry5svmrudO0xoCB1RX9Q1i7dlGSB0rs47/SCy1NdqeYyC8r+K
yHo9hJcTB/UZ6kZ+QWXU9mgHUqS5N1e3gUj268fS7W45vjOvvDwCxZ/P8l4sSUO7
TE+LnAVgVg4BmnouEPOrSc5dSebuBvI1Zr3S/LwqQl4L/3kLPFc8uiS1PXnhylbu
0O8PVz9zvXR2M1mng08O4d/b1PT5uty0xaHsOjOVHre/0WijPNtMJzDHpMiIQ2J0
3NEGkNfqozdPyA67scgQ+ye/9eFkHk/5JHgioNgvW+7vFmt8hMz9VOTMSssWvw/H
6HKlq7OpyEB1WPaGvy+sSZlKAd7Kz+B0EKCK2oltpigNz01mbz55MsLicy8FXeRE
IhMDWFaakAwn2EKd+NWslPxM0QBiMrvONVdYehjxFGiMx3OJLSbj0vuloq6kjE3K
rpVjpJeSyjR3s1Rj1ItFaRTONLLUPjax0vOIoqENgRr1PoMrZI0CE1wAbLTineu9
RSbuP+mioLK/zoG58RayBf8HZeplQ6bAkGnLw/ZpYYxxGtwY4gGxZ+ssglQwgveD
JQeLNvDiRCU9HEdkSU9iHJ/nTC3+x7+lGbjrTPezYYpDXSeJy2Y8YO+h2B88cC9x
jVktNk35lHUEWCKtA4EbByzzvphBth/2PZFMLUaAZiyD5n+iiFauHTb+UfW1dN0B
0Dwgvfh6S84kEeyU1rsZiFyqQ/qFwLfEX3tAZUOT7rmQ9bmKGB9pX93toWL0zlcU
fy6KQC+JiufidLE7vb04997urBzpts7Z8PElpglXTaoNhHA7FbQRKUahbVZJLYxA
3OaNs2nbMkEuYNedKxyYorvIKv7xUVE+5DR7jqvyQmYeWZP5GySh0pr/G7Q3VBJf
SZRHXG7quZgTyPnqs3B4fjui0mlTfDTjp4siraPxHjfRd+lBqObklz5W8abV7kN1
QGXvPsrJU2EJnXmQo5FUPfgL8tObZCF0GdfFKxRqaSHjvyEZbtZHCLabgqHepiCx
OH061xAMaTFZ3Mxr/3mzrSQVYIv1+rAOVTloZncgJlK4fa30IwXssbvilI6Eu8uD
l8z6z5iToE5wMnPMz5u1oWxIhu8rKUmI5IrGU1kFEeCH4LEh2SPbJFiKfpQzFfya
pXrrtjuxOd2ldQsItWmps8PXE75YoPeVOJzXlMR7StQvs7A0gBTkun6jqdV9jdWI
z/9zaN2c/v20vSYiMr/2Lzlq71JHTHAfgH7ISfGPOw+3NApOlbxlwh5OB6X8V5jl
qTevSZ45ehkubNY41guEEqbjEYc79ei4ZF74e30hB9ngzUEGTFXJMybYMbn1Zq4u
8JZDS9Fwe9ZLmqBDZ5xkow022bZuVh6mh3OUijh7UKn8MCC/FQSm26wOxsH+kC4l
S7XFoW3dHM38aRQlN3JlXi6ajYt7Fd0L1ouoW7q9yLssj0EEfMTnD7Sh3693UE6B
nDT7I6NUWi6jC1gBDTiJTt+vrxWCrriesGlzT8M7Uo6Oxu+AvxTFlmyvWgtZrjCz
yURoQ7vuCUZR3vXaAg2crtrhYZyWq3520JypcYhksMV1uI1W2W20ow1dQa/+M9G0
7ure8VhJ8B+BgLDg9sOL1/9ia64hSnNeFlTaRapnEH9pyCt/uHGB9FNeGvqEVT3N
jTf0wR+d5G0FuVNfSuTIpYADxZa+Nmudg9Y0De/9rV3jOTY0ufjLwOv8st3ND6qy
AQd6Dyr5D+kXo/1BApZERn1JiIZWPWLEWwXZdgzlxXBeMh1WKEeWIXYD3c7FAChC
t35Aou5SZ2kzXKuw/xhQdtanXYt8Dji2Npwhm2m4MFpvZFSEy853ru7fx2jVJF83
Oqzuwun2vegLzEObPr3Qr1/jV9G48xzaFjjtkM5bO3iDa9NBHmNhoua5Y41bVqT6
pF4nhINB4ilFJhOLY2v5CPyIktF4mADMNlnZ56fgeohJms7iHu+q52TbmOooXFyc
4dbVEoNx1uVEyODCQlW7SuuNBMvtr59QeYYIPXcO46phSOg60gDRfUlZEZxWAWyV
EVvvSUUKMyyjKhP8SHbubB7xw3P0jDORIb/zqjkM9A82Lfi+vq95W/bKqdbaCuu8
3NX/MFlhEu953OF28vHR/5nOTIIzdugdn6iHkOL/wcoxEIkIj+UtDOOQtJQWSUyK
xO1LHe8774d01idMUtB7WiPfB687BA1pf7j8D4gsej4lvE0dM29PdWpvOO877sQO
sBG4eMjPqiXfiVC4ziIr1Ff2LwOm8aSQnTuUAFkgirPtJW5Q6d5RX6JAKEFt3yFR
N6wcZsiQsUiOuld0sGYl5lBQfaJ7S+ylB7QPSl/Mv0FAmSb9ARQl8JoihD0yLaRQ
cZ+/5OFMw9PA5+jkg3dU5eaebDFjQO3QZOCKtDz9x8qp+v+VZlk1PlY4QYWUVgsG
vC+v+32bH+gQVexmoAgLhZKXOWSCT7BGHNb6biB0kewqfk/GWlkowu9Qv6uaP4Xg
mPEgpjck430d09nA6WWcaYIMsBAcWg6Myw1Zi7nChIVrBbr8SSk593nsZpxI8b+h
qkLDYCKY+VkxMlN+XyshOx1mil7C6Gk0jAG/Z9ZDvAIhPgqSMJmAzWIGAAXU3Ye0
tg6OfM8MOIPiGmYWeNMMetndPSB8UEXzx+mpnO0X1+xxREAn6dBE6CeYnTLtdMCQ
cP8WpGSc5G1fjSBTlgqjhGkIWeh0893ojigFxQeN8LxKLADP2DAdrj8R9Dz1jjrK
knqwoEK4wiwTR/uxyA0Jwza8LoaZaSvHJ4cpbTjajp30v1uaMJeLlrf2UL9V3eIM
AjkP4rkoHqwD7gpEDxzur8fbYpkTTyIFgmvrRVZls4diNUUAGu9/dGK98qyJdS0c
/DQIB/KZDeLHfghLHvQSGJf5XM/7jQNvaF2Zae7Ut1orB3KbhFXMwDS2h6w8/Skq
u6aGxtHF9UvRRkqGp1ThMRn8CbmKKtogG/eYgO10B1yNyWgIT/+2yrRtOHqGDqdX
mMKsV1n4GWlDZ5suLuID+8C3PHBrXDb+aYwXM1pKgItc2TImIWVtDEWjsCM000fJ
y9SqxvLhEany64MEv1S2jN11GJFkYeIgeBIrno/ztWZA9Tqex0rIbbZAgJa/Tcce
8dgUd8D5nvkIYd52XhT4SyiGH/uBQ0UC0muzDgWFoORxnZxjRVqXJ+vmKIiXnxWr
3qNNQQRKmEWE/BKJ3v+B745ed9lWGpmpfQGy+sofNmf+V6lzwvUrSDza92Ub8WDz
sy657Cv/w9trB6fJcLaKm/RKU0a2AwTrS0bLbD9kdS8cwLPiOtjvMdF/HROD7GNN
3CQaL66usI90sSVKD8FlxGIW+R+i0qqlbr7iifpJ7/UuaPMoK/0GWoWawB5104Cm
YTq0zuWgdcs3WSlpmMch3YDMe+STz2bLxuXnzBpLPiw0EuZJoV/lStrM8mr1O3T9
Ay6ewX+fiwdJLuvahuz/ioX9w9a/e1xD/1W2JN+cD+uO7UQI5VnPyAGkFYgLn8ou
2DCpXZmu/J0LXukzaEEfaOCjouTsI+0Gb/iJiutiyUjhmSynsWBqKMhD0CiMwyKi
ZWfFNI5fVxkaQuFxubdTVDkWgyDl2+sx5k34Uy2cNG0lMmzJnu0rpAOU8L1HHIRC
urLzL5nFvyesQTVe+gSKeWD7nYC64Msq2pV8FtYZSOKfhXwB4XqFET4K2GvFYhd4
JDj+uBoHxD8cY9viliSCEHyKyHHj7dfKsCf06KADkR+5e6Yt1cLwaMisypwJi6Bf
RjUqStKa/x5EJuBJM9GruJBMQORrT14J6037h9Am1dhhG7lbrftgTZQyLAZbsb6l
nqYa1s8tYaojHeU8QkJ1OEqvNQTY1WCB5ipp1mnn7iCCcF1i6q939PjuPiRbXZUx
DDAOhNXZaamHzSjcoLjNc1aHvRkH8mJwM4Hv9HTTtmwGaPj5MluDyvbuQvjFWw+g
OMII+jWYM8JwJpaqGMB4QL5iGzAMuYFP93Q6ZGZuAiP6hw2SZz66hxuMKc/01jM4
LVHOZBoszoIci3myqXhxOdhh7arE2TNSkjgDbR7idCc4eI/nUVvSjqtTNw5+A8bo
r9JtsAyG32/Msl506uTDpRlOMHEzHzoxj/CUWZ32QPy9v0rS4WWgoE3Dup3hUcxO
HLqWsUA8rXGwgtWWrBIdLd28cfyBKxQvk1aR7j+exU8pG9iiULF5chjvzihjza1J
25S8pERyARob010n294aoFK2b1TLKw+ZiBBTs5K+UfEgIQ7Y+uzgHRclZCtlYqyQ
IDrDKoqJJ3LGcNntVs1YiXJ1my+bwvaA1S77fffFbnQNdCzliilNk5+Fu9zNP+MV
WXWpMc6bLx2tKqon/cOD4CECplE8Wkfd9saUTr6RIlZPQDvWFRFoj2g5LyaHJ5of
1sBYfovtXjt2tXwkZPWeUKHq4R01aF1eTuQrQr+Kgjt536tJeSzVYqaKc4xSmx10
de0iSsPaOQ1hNby8T3Xri8K49yGi+m62qiAMkWPfJokxriN8pIUJN6Shmg0fX2y8
C3QLzLiwp70ETdNBCBZOhBzjtqiYCz2tWxaRSY/Z+nwbhBy5NML7lQe1GCAfs4E2
ehQDHF7cyJukaFReNUw5TAPjS9z6n9gAigq7xbBnLC6aMPzwULwl84GxA7XA0hwx
DziKyzGoOP4PXXFfXYGgnL3TNQUiXD80Rml0+BhBTMhssrFaMDxo7BgWWZE1tmwT
dDaQ65T1IJqGJSVrAw5+b5K0pG8aTE4YY8faYZXR3YKpGVf1BfWnh+G1pFMNXSyc
KgQ/SOPUi82bYfpl4soI4rxOlQhRukO3U3Sh+7sDk/PGKpnpa6/XOtOURU16LlzC
axGPTjd67yivrU6ZP980MEryy7jPzWKMjRX8eGCtEJw80qfAj/f+PSjSYRWKjKPE
j2qtVrC1Mxr6UvZcZFJMiPF2dq7nQOszOpcqtth3bV+lDQK6b1/Wb8wwoLSRicG7
mxkQMhafFmbZFZN9wMPIrs/TuSbe1O06k1BSGBOSRERknjKGBXuttUgDKZk+1kXi
ebj4p9rhqPYuwkpz8xf2G2ZN7tX/a8+utsIwjjOJ6LOrE2JFGq2aZGu416esGKH+
G8cZaFU1pCx0LmZEdVzAklVJ6UzbmMuH8P7Muge3K/3p/72GjCjkn0w8dSNEf+yJ
uDAoxgjPhywQSR1OKaqc1UmhqnYE6yWsJCbYViiNLzM6N2tq+kXx3cW+0M4qIdZQ
RsNw0D4716m7kbh59ha1oyeytG0F3DsJ/OyuvwWYfTiDYwyW1dgCIioQgXttIAlh
hHScDfwwa/C30zfuPjzj6eWuVWZQz19nAop5SHk9KLwh6hvtE417u8VucwZrKZcF
m1M7cMrRHnVKqHXvj96b9pCzJtV9DMpGC6d0UfPwIGRmrn+mGEENbZiGMabV6IOL
RrM4yRR3dM21+eLGkfLfnOuZkOGHB4AluSkJxMowQ1HFNqkteeDq2eVszKXNbjIC
vFOJsynrH/RNFYERqd40EJetMGJhJ632TDpEmEOA5zevHDgPgTyvcK5gaJJdNCoC
w0mkLkM0mQCBKugGwnUMu+dpYPgW1FcqXd4tzSef9y1SlRtum+XyIUqHOjaLhnQk
7Jt7xwYYJSa7MqiEdAtut3GG1cLFjuGjmeFNfd57ONlNSuhjoENIp1dDA6rvI+cp
E/qcitL+OBmtW+FoaO/kov0+FF9D1kYM3U4CtqSwpnPe1cJIYGzxz9xoEQWXHSLH
XegeVsyaX+Kg0Dhl+qes2M9si5wEGc6J3kImLclIjKyMVmeykC9fmPXJedW8obYU
n9nGohp9LPS/nqC0y4KUlqvSrUvHo74stFkV/tXC0SeRNYaI71fcHbuZ/3e1zAL9
JPMO99QpEhPTvLMElmNIbLeEXiwCDdVX5uqeDUF+kBa6gFO36Xkhi7nI6JLaF932
oTv8aZ1Wfz9IWHnpBZPvJoMGD8jkg3bXcQtIAxgfQLtRpAiCcvLpI2qYoCY5QNSE
POLwkbP4Q0TJXYyaKls5tTJZ3iPzgN2ymDC1Bw9MyU6R8CsmH0vUxVzr1jTsqbWY
O5FoJQ9tMqZhmDPuxgUZQG4KycyLPtMJmwQnsLZewWFThNml72FAlr9x62bXuRXF
U0cAwStW4sgK9rIJdf3qVew11KEAA11MHLlAzXHxUi7HL4UFGMdj+g8hNb+tNCgn
R6VrWN3qA+JBGOHl2ioUqMPQw4m5omOzrdiTer2Pk2asM119cEOUrJQvCgi4YGLS
x4qhyMn27Kg9G8Gyor/F7WRGKgRC+03b6pyiZt6QW2tOkTqmK2AaqAeThSl9ms4Y
SJnPyzYU+oDBp87Z/URrt78LG3fmjLzk2fZ5C8pZn9U20WOR/RJOsNmkIHEkuCJN
Hz7UFMFbjOibxV847E/kJc5OVD5tf/RbbTGXxa6wbTjery40a3jB6l27wP7VyPrw
1mXOgkSwRd4HFtszkWWZWNE3/Sd1CXZEFMCRll2Kc6GU9+jkOXuRsxZq9SzE3ELi
nal54Z0FVPeIo2H7qYRoxQVyzBwB2SS06XekyQ7XorEtcf73ZDOewTFSDmm24dUD
dVEsuVFPnsQ7qARnm/yOVDmLaIHwFX+mllzxabSW5rovmJzh36wII7ZMk8K/gwUh
XJX2uKS+BdxYSH0C5vBefQEQKHt0FaXm77rcpFKR6NuGF/iM5pccZrMQ0EQHJXvr
upbOiIocNSIWmmSkBQ9keI6+rwbYva+LskMzP08GLxZXO8n3rnpP3QiIOGtaHdh5
tnaYIpDUHgR57RyOIFc/6jFL7ZmlnoJknudrnKelVTMEOCzskNHTtoyTi0LhXK9m
l3rXgz2QMtsCuLixoaLt0vqU2NaHRNrJD/+uDC6DnHoYZz0wf6VATRxi+lkmmp44
2wa9NbpvPjEuh1CW2y8ftTLFxyn0CKpUTj2//x2bvbkrtRR1928KdMtGkOCMlH2O
VtS5yXy9IDomYoQ//52Ur4skft4mkZji4Cfxebo5YNKAOqcPTpy5cReCgb7Y52Fz
mc6y/HFsEGTAfVRLydFsZ/Ya3plBKJ0KITx+foNrcGo9eJ9sZVrWp8FrVyYfrFXC
lEHWJiD87gXJIqX7/NOq9rF9WKV1Os/MKHFd3od19iG3c82eKOftAws5bcgYWOCf
S0xnPZofQVhlLLZWwZqr2SuaamGRhIA3KR8FabfIFFqAx0mhC4EmPFSg33/ioUmv
Et4bUQ1ZelTB1A/au01tGEjh7lBqk+VKtciDwQJopEQ7khApH1kY1fHbL9IactHo
Tphl3r0MtMO5DFlh5O0pQJerFarxquTcOhboBuIV7882y8ycPWlPVg60BVto/Q9J
NR7cWTqtrii8bDNiKvtXsei/x0WM9LdXtcsCdel9wcEAcz+u5iM3OkmUnf8A0m4Q
2U++plKKhtFbgKrUhUszWuLXJDN56ERjlIfvzVoAP+iQ2YEjFYsMBhobFzI9/C+N
I/BvnQfWEut8+bxI9PJm1dpRmVWmpxDQjTbylx3lM9coWmnMUvnVer3ZivvNruLL
oINB+/dnG/BjCjBR9ukPoDbvGlMWO4ViXylXWMCwPj6w1j8HdtJ8BHVCfTMuuTvq
KMe0QJhw7rcq463wpuqBwJnBM8cxq6uqZ6ctBSmG9VJy/dWz1uq7NU4+kbmozcHw
WM+zVtN2rC49mpA6ZDbj+tOeAiJRxV+F6B8/69SD5La9kGkNhpIC19LLoopF7qp5
oD/JLzJom1rMsSk4W3Wq45PvNM59Q/RWgbhpgvr1BC6oHQRK8qpkXUxWAXDSnYkl
pPTOffuYGG+60cssyyF8e59b2WFtFhr5at0fJA3B74vDx2fok1tP8Fu0rHcZl1jh
V1+mXwozBDCYJxcyMHneT6zfMPACxQpYNTDInTKyBu7FG6MWm5JMzJNNdwi+eOFi
JdEGjFnbcwN6T29NOVrBax67l9F9o1P2h5GDb8kSGg+D4ZadY6gXMqC2CQYkOBo1
8opfW1QigsAfbVXfTmp3Zx3qhlSnoTAIaMOkhDITXDA6kXKq21XJa/ii4AFNBuZG
/pp8jWuTH5vcoiArtTVJAT/NOCfIzlFoO5EI4gFBl919y2bQEopiCh+ePjfqccQy
coJg8ZtSIzw2yg3O8UaziMECa6wNRSLGCzN0Hc4TTKjxsiNwVrurd9IfC5ZGpWK+
9lb2rpSMTl01eo7tdt8rbAowYN/y3UI0cDaKe8mEHWXwWhW9b+qfj7wZBJH3qWu1
QQQSzGxuDpgizx/d9M52DPot42sL1kXe2oHcfNJ1RbPsEQqWLrGSAVRpGTbbYWAR
57hRU0X3cozYPirwp26JuLpnc7LFzczhPtx3jZx/aowoavm0oqLtF5LYwHevppvm
Ep+YiMp8eP+1MU2iUOCGmXoXCjNG8Uq70st1K0rTZZLTSMpNVukeYIGjBAGEbGyV
kypdjtznq+n08KtVf3YEjrXu3mH/f4bzB6ERd/Oca041867q93YlcqDnLlDu+1/J
i+oCFTQmAssKXGMYjy7nLgGvlWphty0l/zzhZAIxNEdfKOhop/DFLwBO2jEkVdBK
L1MqJUKgXr1y8NDLrznxTd/PWFPIa1UT9dyLRIXVX46z4tjYrhFO0/EOlB6TCBbS
AzhoI2xDdOt7lK2L/Pzq/j5oklUN/4YD4nhK6uBQ2+WU8JWzi2pp6mEIFvFLd0hJ
aI5d+mZSP/wd7MHDXw4HVRZ3EHI9ii5r/fQ0yBMgZ96IDFBVbPD73c5TIT2amDfO
v9h2UDcXH4wl8UfZjCA3OwCqxwLPXDmjcs+s8mlb/5GN+jyL6Ct+hIHH56RyYxYQ
8s/Idjb1svBQvnfemt8Ln96vcVQ3g4q1WMSqc2z0iVBXtNEs0MZNZpVQAwIvNiS0
kAELj3vvW4rayzh2gu29yYfZ/hZOucD9UchBwvj1ajlZxwn62sFsdTkcAhERUWam
g/xjo98AIQyKvPJEngOdpKPsJLvcr+zZZ1/AJuKi2k1FxPj9FTs8cR+rveZS6krO
qTNHcwmE1niaodi7bSvb33ebsf0aQ36RcNeH/dcBNB8Mbvw6GfY+ueqqz1Zi6lUi
YF8/+MwnVHwFkzW09vNaV8nhBAW2LDIxpdWePni3endEdP2gscf7ohm8/M3jn19i
awUvnayPfhgQCw+OzRMhGbQyTXB39i5WeHJD+oj4dq6Q/6EQqyY+EJQjHPtX4CUo
qhrTAa3f9KPb53sYHORpe16OMhlq5onobkspF9rasSEjE6Nw3SyqJ1NE+arOVhff
5n1etrsZLmScI/CZnt9FL+3dKt1Xdz9cTCD7fi5RJKO3EiP/by8M+FxfF8nKaMjJ
NLyS7e2dbToIO7owi4ahUViQTyZpHVwXrwa/GSQzlZa+S5w2IdJ0ANuhWCBjuRrM
m8Sz7G/AGcX6mTL1ak0HxDXc5dpUHt8VMRst4DgkQBgRRbZNXGEQrgNluRxYdfMt
Tsfj1dWT6Xd8eZQYhi0ow9uSHdOepdlXSX96qKjx7oNuQKPzgq8p7EKRU6QOdfP9
IIBr/6y4/RkusEyHMuN7m0+AXnhdLVpyTfAtMZR2l44inuioMfEoSa4z32dO0yh6
pTEHUK1cS3rKmKCEx1i32HIIA+ZW0+gGGBFlSmb20ki315ATFL4tu/+FuXwe3tDD
2sJATzZUhqAThS1h5pqrwKncnNbzIEZjh3oB3GUcMy7PifxHSneGRpaNqxsDNczR
8JBdTGGmbGbsJA0ctkVsX/3rcgYrZO5yMkE4JJsNzaYQXSJkz4bh+gHUAojiEgOB
jVHgVnHYCI1Y2ZfVddhIDdZC6m4MJ6GgeRwcAuuZrE6ofpyn4dKNz9y6Sw0jQ1cQ
iv9ukL7AqJKaNkkl7BZVDwnNqK9Dw908pGDCqQO4F5e17taDiRzspeFtYHN6vgEX
6ATIJQuStO2DfNJZoKGxIdZNW1+pTuZ79wZwVGBBviV1QKcwfxEik/CPB/7pGsmP
amBnXvZlrUSHJW+urXYyVlWE/KHEHRyOaDGurqi7GQ5vQ/W43gPlN2WM+0TNW503
fHAyYmMEUoLxPm3AkLg5CFuQQSip8kmP6fUQOqvWqnIjKQ2r4etaD7oTUY7qub2P
b6+PyfEEvX9mrgc1CmxhfY96lmhfyMh8VP2fvxanGPnnAdLjUQ93+WoMU6qR5V+O
4eCdX0SoIII6Tze00HMljC7ei1TH3JsSetKnjg2Pvv08+3+2zHYMlu+DwXCWOUkI
DaJXOUh5hAP3oJcnczNu/ycduzqB/90EuTxIAHf9NHNdyTKDegxHRjHM7osDVi/b
ixC/gEZgPcDNEkFa2NXZAo2mHPaa5fHtJ824atNpFfZbQCLV+9J2sHmYzottIipo
vDxu6582G9XDrGFLJYJ8Rf3G4ggQHItN0tVmIJDXFmlkQpQXFRfIryApmjxNqT2o
DY0SAMQvvFub2wQCW/uQn2nWiaWRA+u0ownQlC9I082MXwmfDhxB4I1Tm8UjnGGX
GInz2UJEs6JTRnsbS/OGCyHbSUBLZErGG/fJZbpjYqdS035Ry16Zp3eccyq9ZNfP
EgCh2/S9ooKupWs0tKuK6+couKtbQSESqfC3uW+1/LkMlmxwTSoAefpdhvX31IXy
E5RUy3z0n6wN2dERn6ATxpeMMuCpp8VlqILsH9na+Wq0RX3p+08kMdR6z8n3wLhG
j0x4TvX6tOVlZhInTMs5eaWKi7KRCLAVfLcIcMEB+2tXYSCdngh4/epW2bmiN/W2
lvaXs/jysjy+XidaG5/hU3KdrB7NjTcGdIa+NrWzbI02NoWBbSwukL+UECcME6TV
HYC0j/lZUDhmVEiN5iGyW7fJTzqFamkTAVyXPnM/KIKgWPYhUONNLKuRa83YqMg/
rSRDI9XXdXv0B3uPXT2kPPa2jvt/XvdOtZSIqjF2DayW9Ix2fVpK1eGEcqH9dHCp
fxQEd9fx/dE43nPTVXSrsKEqZ7VcffRH83vv9kahSdjnbVcB9n+YOHmO3RqqRl9H
nH3wDhYqwkR8vRmqtb5YVQ3V91NLNFC6FDdH4+WG8GGuMjObq+UdbF6kqol2OqRX
b42NRPqy+pbVQarbg/eGMt03DgOaBm7LjQyBCbVns4OQckDUXc5mJfNk9yNIKm/y
kE7zGgTMguJIJEDjzFuyna1vi3ZQC8m64MevJ/SeEdm9gVMnaDa5IOFvyUo7/23U
TMs6nHNhS3Y1IVTFO0lCPQGJxsz1TP56KVGc6+PTUUburpIRdWt39Cp+ZBho/0P6
9y5LisuTFYn20EPHwxq3MPpnpsieOLLxIjkfxA5AEXX0PuSnEMd6/D+1zl9hrHtL
FO2kpbbsRM4cUY9LH3P2aDqwh3Oavhxfh4TFecYNIqzyoUglCk8bg27DM349S/qu
GQrw8RdPgpwM2RCKwMKXOjAzLzLsrpl/a4pcY6VQvlZHlI9WaG9x2AuMQ5G5YcI9
k4INmZ8Z9S89npR4O94BWlV/UXgMKehEltTlT/WvXvRxZLh11uvqTzE9qaw2U0/O
f2yj11SsDde0+/b/wBVQz3MtAEq2v9ZnDYTi66Ap0V0VPfC5+4qHIftZQRxrr+3d
7pb4dMJFhMYpgaGobxiOSa/J0Fty1lv/AwuBgNFFIvZcuNlnKh5dDdxJek+N3030
1D8fCXU2uxuNV0BkNYOSTkGHnbSFieMSKiNOSxeMGGyxwT5llsQEIiI6kIr6q2j6
BeXMHHtAlPTXYlgP0ljf0Xsu8NNx+nHkZbalKqSUzSy5gudC4VUxnQi85TsXXFqD
tAdp+NAZrQamOsXOZaqCTUKHj2i9C6yngCRHym5dQFqZvgpwdCqDLvyGT4A/i/Sx
LVDqdb3xCs3FWvswj9HeT/dQwAqwlMDHRUAzTH91TzJX/LHvvFEuyFllkpWuN7gB
doxHxUvj3DUXbS9fUrh7SfC2MPgs89QiyHJcsOZqxv9AM2EUgjvfyiFR0QA21YW6
Y844G/dSzNlcszlqk9yWwUlzQ9J6rB5hweDbyWvDXa13bweB7wvoqjcBnPW+TM/F
mE0JeUgZjelbzMXul3v8LF3OOYqjIG3zlZJ0SrKLkdQXsTwOlR/NKFf1S8RQODIl
ydHDb9QgW02w75lgm3TX4JfkCJ2Plyc60jeME6M/b3eiAKOBc9bUYRw6DX/ICLz3
lIvbnyome4LB9V4bbh0xNFFgTapN8MjAIWKBS9x3WbbjN+AsbH/GmgyKLATZOLRA
cOCduDj4iQl3+24LLhGie4Si4WL8jA0fSQbV9bDbFEc/3nAq8r8CDcWO3aqxAWpc
ayk0Js8OgGZU8fJ0nHSkZ7oh6E+npAqRM/2hkvLBubtw9YFWoh+FBRpdP+dPFlKX
NPqZSFc6y4gC0TXgay2MzOaWRO2AgKJnvnNkvo/c/QiL+CTP9nvOfchxqk+pakRk
vRUZnsvrlcrU0TDvaflmdC8nGgd2DhllncPvcmOh7Lpuu9xbKIVGffQd59iJahVI
2p4fM6sJr6UOf/cxXPO039RUK/7PTvVs3hyNbqNLnwdKsjj20FVt5udldWeRf45M
Cu3oR9SlQNNMfY8zHl3nktK/xGSYOzYt/EVx6NlNsf5m44UttAl8pYSOQyYbr7WG
GolJRVEsYreQbcNCTZCnaWuSalhIo0c6Z3Q4dLVrLsJ1PaFG6BfX180Iakurul1O
zR2aWKFC6Ps6ODGzxdL2v2FqOvlPweQOaQym5xpZBbSTYg5pAVGPstwSLZEkAWLL
pKpzcz57fQbutmr7vp8e6ryXb38ejfwqCgZcIghS2z11KaXQqg2vx2QUA6GaZsXi
E0Nxis555TjmyaNI9sv7cvgOp+lOSQZQ+WJ2gVmHiMDYmQkbtYP12e7jk2DzUoYB
pBlUtCY5AVLNfa+gnakQZ4bl4qzWinlnWxAOJ7LkMAOmP3ZAwXuEUFK8LP8Vm2Lu
bAnjqWzvOCzVTkg9QU+3woqypYkx7XdGW33mqRNUeFVPuw/qJibsSBm8N83FGW9J
fXpvya5IAdRRLJIJCiPqNIDBnCf/0tg35s0hi1gpirDSxhuoXCoqdzQC/iARalBK
jOkscNrGsIy52iOIpTUPxG0AFHm8GvNNHTtZ894onco3fLFvcbWMUGLctQZkOu1b
SF4UPhytP4rJS+FX16B+/T66ZIRcoRXpfc8zkQHJ8kAX8UQNRj9KMhajC/GFJk6i
5RCwNBSO1/ayz6fVLPqH50WvT+Oou0/7klmWomq7Ckgh2n76AS3gc+2Gei+LCPwh
qUN6mTMffmaBpdc3HpYHWL1JMayKxeXd4khE6Rq1eeFHeKMuOVwd75HKYzyOKL14
AiPz0/jeHBlWFRe7wNlmUHEUMjQtGKfJzjBMzANp5eanaxEhMk9bZMGxmr+4tHGs
a13p9t+cT4JcmVQbXXESNh79cjr8rxvd+rtLr14bCk8Fhvb2dOoIsYnCo7sii6JU
YEfcJDaiV2DKDnNofSta9M6lKvxPct1rMqjSnaJo5lIsP4ESxezvzi9CL0+A0vAF
AtmN9PXDHXdzJQ5/l5xSlFdg9Awf54K7gCW2FCDXU81Z7hjWhndK8HUEZ7/fHlsm
xoK+HKac2vKOrtinbzUWPKTGgqcEiKgcLPwlOpr/pS1DGYsMcpfynkh78JMt+pYQ
r+clx5XClA+a6wpM2b3S6w1vLAfxnDbMF81xbRykxc7Kp07HaA6LMeExxhxz/ZVc
3biAbaQQlJGTvEsZ89zk8xn9IUNdnRfNKCcFQe9aDwkPurLPsbHs4vJvfLIHH9MY
ZnbdKCg3xQESysokEueASyE7pMsB23R39DsOQ8ubc5k4GkDWoUc+Y4Vf56XdWArB
TXkzX9BaA95onA9FwHtR5cRL6tPTX5n1Kbbs4JI2xtZAUDqXNY7JM7sk24PbSsdS
gM8aDs5RfiWZjo7SREz3lnmFY3EwrTy5U6drWw1rbPJCD3fqwZG9O9r7T2Q5lytV
lVjj++0+/AecOchJMx8MLXGI+la8A6yhPvNXH4WPL1yF9vgDfg5V5gZTPrl1j1Bd
OjLvjR1wgVXxLy7BzVEl7HeQUXWB9Bpxg9r5zYcJYcbH+Hoccm0t8HKoJPwzFMbY
rO7GWBNnvn6icgZnnSjABYYG7+BJSfe29Ox037OqRvumd7mfAijyPwl/gXQuACwi
Ol6/xzu+QamSsL9CkSuK106RmnfJHXOk6UmmqFB6HSVWSbNRCqeTjzwsYaYNTIn3
SK5oNwx9pFOUTDQVquYrGNGAAgZIDz0swaYb+JlQVZGrDR0a1/Affo8jSwziGuRe
wCvMAKWOSIvW9HY0/FIDPud9SORbSTkKENfe8/SS6BQjhKlrigJgIlZvewaWQgoi
YmCmNz+z4Cqh7lq17VSPvUoi9gypTXlBxgXA+nG1cLS2j5ugqwoBzNfDRMtFj0qz
HyC/wxIB8aHPSVkgvs+8JtkuYNjJLmUVgA/SdC6XTj9vneT9uLNLyS9vdfcdGcAE
TwhmdVqBIP3KQFM2hX6eMHS0vWPHGkDLDjzb5m7TCO5TU6Fxo6rkH4HPMzZKsDie
SXRBZXcHOXzwZLPX+vpOJ2858nkupRhj8EbBKy2BaKmtr7qj33W7fAtk0ojfOyyZ
KQMzYyMjVUEENxpHVvgKPi1rOyjkLY9kIV+0P+ocot7qQEluQ11wSrGHJrzFD//V
NY7FWHWOEyfNqxHK9HW7qzCablWdrNbsplEdOdm9QmwGn9GBZ2EjrcRqF+bsWKc5
Hf+pBLYa3baSbJZiffeMTsduK7l8Ozk9fOFZtt+fN4ba/YrX/j58jURhE6pPoN64
rapo5SeCAbff3WuZmWt0n9+1xm2iIyMoTgyvDr4tWZov+Ue1aK/Td49Fb47yfrOc
Mirt9BOm9p8H2CNc7dgtFbfq1zMZ7KXp9xRbTmwoqqBLFD2oVgg7SIR/6mIGd2th
fZBO1DtxqjSJsk7aRG+JXdN6pUWj2su2u74KkFQ4dWIC1/xYbhlo+dYvKvABvNx2
C4ZGuF8kBuEkOmy4d82e9GjlEuS3i/kAVbP50nlz5xVbNum0zqk1oJ7bvaErgvK6
CL9AG6wV6mnm8dtWixHKwpUGtpAaE/Si9aSGH8+4b01in2o6ssNipM5LKCVyM3ln
6nFMR/ezFWSWJLzBxVoPBKXHFBn24EAQDAc9yQO2dOTfwIrTumyqFleSliNOSrNs
jApvxWAUT6Drvm/+7YGsmxs+o7+/UropjypMsosO3IZjbRaWRIh3luw/sPI1+mHn
IScAxjC65TBObOWulFbLKNABH5vJ2iBJdgh1F7A/Y3h+QqPVEeC7JqU3XxOXbzbt
qFLwwESygx0etp2pLvMPBm8qjpJGWNc8kHH4FFZhhZnzqUzHZ58EYFYt0fMLwaQK
TGG+kZ6xTGgAYUabfT0Y2+so33UeIlaj6iyCMNqnQjgMSatuhmhqM69JU4XLcTqF
H/jRcFvM4fB/wISyt1HFcivfpCXVfhz/BXSW54cXqUPIc68Ni1Bs5ZOA8WCIVyGy
Y+cXeAZFHJF26gAb33i7Kws0mjpWwF5N0w1RC3V+jipSXqakeNIzYHIsfg0TiTLq
0sM8Vwdl6mK6YcPG0Q+ZXAoLtARSvri4nQC+Se20aOkmyZzFvg77J1Q2VsqYiZmx
uMvC/Cb+RigAhX+mpyg9q+XoRRduio1jR6h4j0kfMYF3rmrrms0dLpmuLMAxNSAU
9P8kUSq/h1pF5ZZtuxbWb9DVYd6RLMm5U+eI/+80g7gFI64ASs6Rq/+pgupD2ZqH
OghdJMgFZ+C7CYMPA/QpLlRxHZz+flenAiLKz7VYBxetGdkSrWniHptcAkZnXWNi
lOG9PBmmS2gaOZvG6fhIn+scsDUO8DjJ7He4OCeieCfczE8f2YwfEGa7czqsOD17
kyEgH1x5q7HPpBLyU3EpnVzGjZTilrrCMDl+waQa4q76P36NPWDdJmcdCc/bpWvy
ZXMO4fh9cHb2VLp9wKsv2XgtwR7/u0pSmzrE67y3Xe4sJfxIE2xh52zrhJr55n4J
62uPz2wPdXqcU4FSGi1phLjmWeggQgIlIzwEZ8H/75uyfEQVq8P908SrET1Mi5jm
/GafJ+lFVDr5oC0BBYJl55aFoTboKWVZ/tXKDYYtnDv+4pS4rTTvruO/MY/n1yF9
17MdcrjRDIf6RUJJ9W2jJH4SzZ2UklZmRXeDUMPbV0eEhCE/TvfljONuG9IQlwec
AHEw2g4Rz9+ddt+oEb5+tQzT5ihnpOHAvzHi0zBvHl19pyUfme4HjQrMrYETZqn4
VzwtkKFCEbt0r0LD8chP4mU7FIwtu6tgaNueoTXXJqC61ToUByigpule++uQ/q9r
ZNCz0DCFK+THwT7yjpqAGXy2WIiFVd7x9f8Kou/1snCFWDQUEwuyUbP3VCLrJX2V
TQ+j42kU/PPGbC9tvfTSA7jlAbHPdDyRQ2/kEeHm3J+GVf/KV4hRJcL9pAET2cio
/fJjVVlRxOd543W4bylcRNPfRuDBjld3TVL1c6mPNAhYpwRuC+7SXYVrUBDelgHS
bPaMJUduRBiTAGrGrrFJctzK3e9WS8oEdGIVZLKPlFOehJT7JdxobDJvAh4X1Eep
qN4Us1/KqLT3vIeaTWvHvb9rhaBjCoYV8hfAdGkXEe783qypj0Pyg6YzRu1Tu7+l
S3yiFm75iHPCxD6elOb0E98k7uOKET/y6TBjMUub7dA60MLq7mzVfGqAv9uC9Wvj
aQ4oRwVReotToBImLM5gAWErSxhrty1Z4N9gETt6k3MCICK9yoMjR9LtXcQdI4yE
RvqPTMhaIdhou29Uku5A+MUD8oBS9GVAohu3RJSYC4mWfgfF/rgfoxPxeiuOf847
7qOTPSFbAP7CIYOSctBcvRrzojn87vo8gqVIdPPwAIw04GAFlgQWWN8KeIYIyYAV
kopJp5t/4r10ubp9eTBAu4TA3ss8dNzNFamE06QHwrbeRLOsvQQny7eohvkyel2N
GTjt40jnfs8qmRjHojd4O6ftgwwP8PMQcrGXrKIRGR2qKBR/qD2GvxcTMprzrmU8
kzKeWBvwExINzVVCDspFlOaRh+DqPmZ4jRGubUufzSrzmjKHSh7xEWxBGQUwpk+V
r2waue+VPTPb2hpZavsaXfeQoZqfr/KSc7CZrVikT7qCQNhSIQQljJQjonHO0G9J
kjdzvraNbqIi74CXZpT4e9OQ29v4jU4cQ+qg+HLaEMdhO/gIhOg1p3m37SIq51Sc
aiq5Hl8QUgH9GCJXRnQZoya6QFObuBhbVUoYFoUmZNzZLe1FVZIbcnkuPkQE44hp
W3MCIamp5J5JsvyEQAUS6HS8Ghocw/Cvg5mtN1W1CIaVLtiaTv/e2gLKejdddape
jREi8Zc0GgmM4VThIhzv0zjK17p4IMmgiCjm0hVZcz4pMQLm0VMRnjg6S7E3ZFPM
YkLWgHrkKUna9ZFesm6MYnxBFlfHOTTtE7CCDRoN6FZ7z4bGR/WtOarxpLy3YupI
bTCILWp4VRj77dptqVwQlu4eElUDWOXR/cJVGB+TjOm6NSiy9rf/ZLqyKXamsMR/
AOcEl5mcju6t0Bpf4opZKe0gyubpcZNtq1PErdeds6Dj5Lyv4ItwOXiwz4ApRSxm
P9yF7bt+Al2vgdZ1RDKswbeHkwmBNDMBmNKHWuNOe2HmfUYeoAXL5un9HTB78/3F
F8a/gqRWc2ahsMqQmdBk69v291JMTxqyPp1uBDBUTU5erF8LdpD/Hk81fUsDc8U/
5aCtPuXKTCyRtLfVfD6KdhIeBIGRvmRgAz32ZHJzg05zmxe3J9PacvzuCu9y+5cc
O7WBy1fDLnErpCa3MOhuDdeX5uHtLZnMFpmP64Nf17GG7/IEmcgX/PkYDR0W177Z
u3qc5lA4gmbu8UP/YPyRzDO7/bOjc0Gl3kf1psDhmCbuOMGNenHJjX+6iGMOHzKn
CrEWvgNZqG2c63dUI4XCAjh8cIKPCvCkzGhbe2oEz784+uCE9EyzIHGPnNkvH3Dt
QKArHnGMeUYB5E5ij3RxQonvhjZWATIru/RLat/6JXdmapNTSB2XKYQoXiwj4Ist
EWfg+1onp2GLUItBZLsGkKJ2+zG0WKgSiNOnNCh4F73tvEyOqR/maVVr6xANr+ag
O72enolJwERz19UzUBsEV6iqD0SmnX3FdJ9SRUSPBAyMnYnKygIGKdr2uhQvmSU/
n3tyQIYXLuG/qnwtzcVgZR8K/Vlz5n4HOCE/gelwltk+VE3uKZCxgs9HUkQWEUkk
Xni1jMmUmNszSnWM6BPZphqdV5DTCEkois5Ohl8nylPFFD6ObWWEhMsoJxqaq2ci
qGOBZQDJ8Q5Zr/ToT9PsUNh/ljCvl5s0Q3UhnJazcovLFOZC0lIDzZhAQLlIvxl0
4Syd28t0AoF8ySR18DnDESseMMPdDMWsBCxzEMl2DB31fhFM9/Uth3c1KqnyyvhV
TmVyz4lVo9sZdw7U5Oi76kCYW6jcVYQovGH56VJBP9pp26VgIAsb3t7d8avGz98r
mV1Jk1W5rD+wWNOwKEeb6z3UiwRkUWB4NjMrbhJqfX1SvZmT4uixkrAYgdxIyCqp
Oy6sbVsyBUAEFdf+SlCMF2IBFDkEwSDecSjpyjgG2gqSzQBLE7TwsEQiWw6mMMAP
TzgP/0zVNT3b0wOKO8RsD04r8OvBNqod/O3DNZxGzYXDKSqC5MxcnAaui1ObsnKq
UtAfcocZ5EZsKXEvQXi55UyPDExNrLBkBbeB6x+YQ0RZ/j03qsV+wNhpAfy7d6aB
iBWgFS5xaGwQUd+qj2j55CWclVpR577XkGcsV0qf3dCvDOGO1byfJzrHlXHFz6Tx
b/rYwfEHiWmvkC1vYqRwhkUwDDuHbEna7x+MPZAtMgbSSaRdvPhPOhKycQqPBQuV
/kXYhuPk9JvBatobjH0wQsIeoFEBhSq8rZ0ae5sZueXt73yJi13UqJCm55vC/kRM
F30Mjc9COZZDeaInIcw2IUgKnu0XRm2HoeQp9Dh8RzzAN70PuHsZtgv7B49+RO5u
j4LZQQILt9YQLGqY8XbVUYSSsyuoWwc7neCzPlrSs7Zb54OLDpeFOVHDB5qQ3On3
keNUr8Hw4+xtHGy9W8XOSXu9ITzu94VVcbW2TxbDyWAcjq9o0T69joaoreTyL4hh
jBG5ItH5umHVI+q9n27Ir5ZmKOkHdWHWtRG21UafmK8SK00ARHqbbmLt01FF3JSH
h3nqnuy3eO2vPriob75ebECXiI4Phy7V0C5gtkz2V3+J37zBdq0rDpfTg77cdN5F
WzLp9H2OTObsbEJQ7C4Kw3a8syPnc+O/e0EDASrZXcv4A/KvULmJsJW+QkYbAWh4
nWKQ3wStQHBu/oS8N+4k35gxY5WgutfH/tM59hJpNwMyPWPxxWYfqyGdvjdlkqY3
MByL2fEmbU50VuDoQQtIfXagh8BjM9ecdfQr6363DXxaONKCPypJO54vTezWq00x
RPMMjSJYw27xYH2j4/B0AlpY+XKND1K4ycOnNnRnpE8ghW52QKIyd/S58Zo1vvLa
qS/kyfFBeTkN0QdKWMso/I8Rvb/ZMMifgdhzOTW4PasrmoCBB2ERX3Tx4eymjsJz
AKy5V0Bud/iFsmKSAmD9uoN1SJgx7h6zXXA5zP6HdrZvCwyLmP5f3TqomHnt3KWH
zkWVCA685qohpZzQFkbMUvujj5+O5JkMEPu/McfNd8XcyTvKTL2xLSdHATJ2KsZF
4agpxDNTYzCl4adnYbGGAKvXlfV+Uz9soBFGYqI/aFyPLPxBtghHF59l9IAIGKDx
uf39YQg7hT6tyNsTJhqOLp69U073hFrgGOVf+fI1KE+cfn/TylQtBfj9uHrRRpNw
kGVqO4T4SjxokPqTOhtSJFLOc2ghhg/bcl22Tp1B458LS+jRwi4Y51+LOGICC7gq
RUU4kdEetFlvE0nbQvtvsZ9G9sFJuaAW7vqQ6P6a8yNozcXxhKsLOWGoHqBR7Efb
tQTxKs7ltpM/osFrn7vWMOmg2Y9MAH4j4u3utgGoiyA9Y1cMFn4s4md5l+3ZwcPu
+hZaoa+Ya8FZHldET18u8JUt7MYA6K5W5ovYD+q6Kx1/171jXzDeihNEiygT7fD8
IoRm+s83j7TKx6fYfaQ0DrWEmybeLgwRryHnagcF3nqZ5wyCh/h7vfJFCkbdECUF
5e4tPZBe0DRiN1PiOZMoXXhIHthpY5WBt00oGkolBNwXi5ne5ixYxLovmYI9eeDF
4mdhcYI1vi0THJ1wQeHU1FJf5q7RS4mlcslv/YmJg9NB0Qa1+FyibXN/8Dqc/8o0
ZA8zCCfTMuyARH+RGMrn6m7+JI5U6UrWkgdzDoI8hXkwQSGlrFa6s05NfnLL0txS
zhb/1enoVElCnO69nz/PG6gbrj5YQt7ZA9FmmVPsmN5NUreWNfiYCWFtXQCO+DUy
eyb8dW2Ulhcs8JGt3POGHCuUpp4X2NhtupG5D/d5OXCQMJwIivYLbtdwWMRUq/pR
tK3R1BVsZlHI62BNarPRQx9TDOWGRlbIxM9zFXEE2W7GEGBlxPLgnMzQrM0CfO+0
5JN40ZNCuBAn17lD8/fTyCZde0upAICwmAfEGCaSYXWS8v2KhyJZ663uqIDMeG5Y
CmKp2l+4HUO+eAr5mJ+QuMwzHAkbuR8ikgc0QUr+Na29Y/EKiN6cVvld6W46Svy9
7kTK/SMyMbsoLnqcL02eohFutKpCr7P06EheapLpZN4QzS9v27f/qNa1R3s60EY6
cHYE2e623u4wU/+w6itH5NunO5ecltIDZ3FMp+eOaMW9b9TPnxuoAMwZW7Ku33Jm
XxvenAT/9l9+Mqte2MeA2TCWRhwZn6tMR16QlTcIMqtUtPcbEd4pIGIY55WOdS73
BcLYnN/LofBf9sBoeM2rDGjxOJ74xqICLrOn04V+flAA2x+7cjUuABkd1p6v63uJ
z5lWRDDYx8jaabO5G/0F9ZLVncikFY8BkYST+LnwREHHGmKZL8SPYBcAbf0Hhou4
ZrhSxlQ3h/kDR5H9XQZbwH5/PhJBPEAd8+Q1R/Ov8yeP/FgaloiC+TFccwnmvaGs
WusOp8j6sFJxJozrH3CJKHd4q6Rb6wkhgOvj4+/fpY0WdeG7mpuG0pXVPnikNyF4
w5tCicY66AUksTT/8xK+s2aQ5z1l4TbdOOJ6aT1ZoJPuNiyGSV371lUQLorDVIIU
RP0VEmm/s69X5FJjdHjVyT27Tap1CiAW0aZObqRn4b7QHqIlJ4evd0xz+x/ektFs
EjC9NxvJoUHmlDWClRN2w7EXwuz1/LOecaj7KSwqQj1LaCwnTcAzUDD37zsZZuKo
EgqnglRCz13FohD0QXe/9k1ZiuuQQyUOCyVM9pZDlvooLO8rpLayVRm+v7EgTJRB
NFx4QaSeH/ccG3N9a1kDKj+gF+bRyPrB4Rfp7yp4RJgrDCL79j6GtbNEAvGcH5LI
2yM+zAsufRxQtuAMyPBagMIk8RJBqAPsqMriuLcukVwpofvjEVAKRDBPcAmzJC8e
GNenXkK2xCKeuH4jo7AaxTl3LHtlmo3pWm4t20X9xuY0fJsSQn9+M4yCBhZlIzx4
w+xV6r7AOQKL2aA6d07cIsvteCbXmpz70Nvu5j+V9WT7Q0TACW7eiHGTVd1kViFV
6qV1YYrp+LJ7oCXsIRyB6EGI6d3+6KS4PeVYjUZBbmrbAxqLlkv+A2J4p62a6/kf
FcZN/pqz2gdVxfdsxAuVZjSefps2QuOkVlvX4ogmkZecAZ6RIj4IiDSPSnzsUe0a
01gfMCKrlXpqybcVIvvB6RMHKVEUc1JYu801jsZN08VnXD41X4vffbg+E66/Ci5I
BQcINe1Hrn90hF2WRlaxP8D52rtdnHGaOmTslKeIK9CmS9B6Jc+PeNgMNcjLYqKX
X4PmvgeBVmZqUKhlGpddoSHYfr0IPr7cGaQvfIgQnji5yTol9Rc+2JGEIEymqEH/
L5gnlXvly4EVMt9A93h750pnxurimOLdE8cNW7kiTCLCqIOQMs3bBWrPR8xq79oZ
nPg6xivA6s/r2flzrnnWc8ND/GvGDHxv1HnL02zsJQqtiRyuDj+whke0kL08kc0I
/6PqNND1WQ+T1odWiqhjcoIZDZrTR5jCMHMFoCOUiOfSUOgT+ZqRfnYRVl5Y00tf
6yefIsTWa+Kp7FkEAVEhnZekoITqcsYEMPKsvp1bw0FIIRTDeRE+UY2+Qgfue2Ab
t+5BX02uv8yWbscr37+fodWQZqiPkPnIkv0t0FLUdJeQC5EOyAevI28c6t66oCto
/ctAPwEjrJJvW0c2n2USLcOCGS1iiLQjg6uczs27AeeSXJj1jsHubzhncQypllkM
NxkcOybAcbmmhziLVrSYV/gVITWUBF7Nb5cHujgA2iD0CgLu7APNbzboIgWK3yG+
mCoTvE9/dVLbIXc80dYoD+oiiMcJMCZVNcrWNW2eY+l67qJImRDQoGsz6oVwoaKH
GDmlqy8ek8D0UngMgNte7mw5hbJUK6XIlNLYd/cxHISydviQ3QI+nfo0TEeu5S4x
KYInQ8y+F6OGlaDT5cUCqpKsaljiKoVIlexwn+iDJylI55p25JX5ndab+JM37TtA
519ouFMf0c1xqc3k05bZCjmunzg3B1ZcKzlt0X3EG6Rlt3AetoOSWgrzh6oloMep
CEuOxg/2yCjHtBnvuU6PKtZlmyb/RIB3G+6HaMPuOpCpkNAVG06aJO//89c8+AWi
92qMVQBRT+xK/6A3lVipb2QzSDv3KVwLCKiGezpv3E2iNs1JeU8MXb943EYVr+8Q
ii/Oo2flVpjwyjXVXkane1YtuAibvjBkG6lBX6/qbi5Kol9KSEwsXvdnx6WJ9l/p
yrgRDyekcGV7rwVV04Gzn+jfg2G6H3IjHIWbyXa64kh1frz3VdUZz3t1wvUVArsQ
v/fW3BXUj7Md12RorxWl+yfXxBDWtihvvO6VIo7EufBZK+/n8+gJGZD0Wq0YV3kU
fLfHC9olPmT7ISgSbSDF2Uswn4WKCoMmyDO5cstPu6G38MRoyYY5wSaxj16+6iUK
3TttUS3wbvWBFwBNteeUP2ZMfFoPi8BS8UcS/WsV7x9iRWMrZRQJR6eyuTyMnuPZ
tIwVLS30916fjbs61XOD9oACZNDfJmxrvXBijntq4kqBUwQdwijNNirdXI+sbZae
3Gfd5CB3L/BdUsXh2uPg+mU/yeRuKExbDWZ8KQBFMHaGJ8PE+mQ79XiDY6/3/U9Q
goJDKz8ghQKzogGKKLEfesQ5Iyfk94QH4QiTd4k5oYBM3WAkFzBV99uHlXbZ83Lf
uY3t5MIOec/NnmrCEtesudaypN12eawsHBWXPVjNeGS025dsfc3nieOAqLkCZ01o
T5nTBUnw7ZskneGh5pxUt9KfG7wF3pyZKcHqo63uNKRzxcbt9z6YcrKHUU/NSgOB
/tCBDblSHgkzAjxLWsxg5Hh2xZFSHQqMpEtmpSYCvLfgVDKci5U7kcts2RHwC+Jg
KfIkeXRX+QuRwmDaWt33AafMvIOpq5xsDZHPEI6k4YKH6uKvgAwaXzj4tRfqJUtZ
w+WM7YvUaT0zefKaFR6kqUgYNjonihIESlgHFy0CBlcZt3qQIzv5CDc6bKr7ZABV
V/LEVQrnylFInyy+U7d+SF1cyGKXqkFU4fiOcZ3V/wUX9PKaiUFZ2hRm8D5gou84
VvEkjXjKWaqJi54XhTRxB3kUOrLu7+7k1SKk7wu820+Jbombet0Exzcpb4F49NAZ
KUqsu8RGcvL27IskUoxRSc+aQFfJE3lkD/pUWHTDUj6WGx1VdUQIsuR/HbSNgfio
UpjzPy14yPDiwuKVkx6dbu4qMS6XFSnrGrQfncV4xAQPik9Bk5dt0yYF5HBocPL4
tuMDZP3QSW7pHxvP36KhPB7/POmYiPpsqnDoy4Pt4oq2PJJnUPmuCR2y+czmeoP/
hI0sLQ4n9kP08Rmzm29Jxjccoz5bAdW2DtY0V7g8hax8SUFEBEejUnN9NZq0Nou4
cV5JsO/9NDTyzWf9mU9gyhRDYmQV0EY1QoqWAD2fSQyrUWsFYlYN9jax3XaD7oxP
/m8MmYjKYq983w3VLNS5jzysD74dnRQ9mcYhV+wVFeLlJt+FTU7DiSH/2Zcpx0Qw
Lv5fwWSHWX9ZG6TYqBxj71U7Ci2Gh4GHoDV3exluI5bLRBurP/qic2b2KWDvFZmS
N8uvCYAGhGC6U7gKQzBaKTfFMKN0leSTnTO66slWMWGcTmkZ4JdfcsmX6ljcV9jK
weIGR6xj/y0xtehjaYZA1OXM1a49aZc1KmoUaHciGy7gRHB8227lJ0NnJsTxjCx/
7hWlO/PhaPXNkiDrkUfI3TnpnvZnYWJ+GDcj9HrZ/+s+NGGsfho1f3SUZsrP4exv
nXtmnCXoIdMm+kXqPQ68NLfNCjkRpIoMQ8iqju6xmuDehytxnrUMQGpnB5f+5orz
gpLJNua2dP5mdapx1FB2TN4BXtoXnGwKwGVfxuejscpgZtv4mHYTIpHX51mNxlGv
j8wXnMMLhnVtwTlKdTo+o+FoC1dYZTZERWE0ZY/VGEbGSiFquQrRlj22jj49yf84
+hYgYb3MmQQJGjcxKsgs/ir8r6vbudYmZhsp8SEIripcUEF5q0plTVR/6d25yOjF
D0kt6YtSGqM+bNUPmoTGMrhoroqO7nFveu36pBGHlqjEUl+FvTcfaJuv5nngOig8
2PqkbgiwoHkkQuBsxCoPy8F2lJG5202XDSHEeckMwqwBpHtBBlj5m1yLyJU2CwNq
Dqtc9amsOs2PE3kRiNoo/t8+PwLWH69Pu+J1SS1qz0qbYASFezBhxbRQ3q06FC65
dNjXfEqh8wfrzk/uHLQMqAKMB3rA+CjUNGz4R9NdfPU35cOB64xA64JM27mWzjYA
HG3jZy0SAqAz2+jQXN7WMTihkISJAApQ/3kXLNoiidb3s/gRSnAXjDyI4uYV/iEK
e5hT82wYdfmX4Ome7NLBF0fvYxl55tv/v7CIO8iCd3L2Zu9VVrWvPKxjmvxQanQs
7K3xdRHn5qkT1KY1bE07OOKHvUJNhK7fmNEjlFEZvorzE5PFcF8w6DoA8VOgOcbm
XH7KdLmf/NeA6VnDZAbHdhLghg8JtB8bZpzagmqAVS4ksHMKAkTaY9bqppQ3Tsti
96fBV0DAe+hT/zp2uQyHzB7mZxoXSx3Hqrme/zrPUUc2XrGqhPlv01qiP9ByzPnK
bJuPuDGzaaXTy69CYmlj3FLtcbqPxqT4cbzHfbS0iGC1/xDTUIjptqrvgwU05yr/
wlGRdF5w6O1OUyelj6X9L2o7P1iB1bg3Ehp2Iuc4yy9Tm3Zm5LEeyK5jWUTy1W0E
LKpGiJGLhGS2Mi0SBuP3cneOBWNlQ1pESDS7fLvClVYhW5uQA31/J/nY5WZM/LVq
xmKRzeAtk71aX0EvspHejMWz1aBTSxdaO1Vv3bebZdUQKbzM1P/P+3URpbKD2EOu
m/G7VYNj1WfqAgSWjNEjLBUeK0S6snBs96cgptwD0xYM/PZarehzv8T36II/2AxJ
gp71hckA4yLFp6BBXT7bMcp0SCeIGAn3zYDzOETqOSktD3MFRhPOMhD2wqFUPNBX
ODPY4BNEjdGf1AWgi0oCzrLOSk5jZPN/uUpxRmQ3Qc9LX8XWfq+5EV68R8pwmG2V
j3MTp3ZuByRKxW3rDkvH5Uz6qQRjXFpAIyOLFJFsnbdxhmVtsupuzxGS0nDzq3Im
dbdHVdwwwfJ28nqxsYNQNg/+r/sdVnfiXI5a5w/TBbPz/8wiBgnpSfjQffkR5BaV
F4ZW2H0io3seLzZOnl6VR849DOzZ4IIG12lzseHvla8Jj4jszJXf0qUZLxzZcGMf
SxC749Eoot4+XKcOo4VN7dPEzrN6Cj8oA2UuAKhYdKN5fMWwc6ZijCjEZ80+oVYH
E0xvTPWRlk4CCE7wKgnv/wCFx4Vl/80ywz19Lll+ZAHmHqhQHwgo0hG1gP4oko/u
jjAxzFcM1lx3315OfpvKxHI1yizkgQKgCHrTMUSU9S2SwYgHZSj8LXEJ2Km7rzxS
PZrL3bcJ8rZCai2kaHTrKGksAVRufhcnzNaIOl35yRbwjBlPBjQ9nviK/BtGyIWd
gUavq/FINIV2u1OF8w9F6ZXR01Rsc78fHYgMD6vdaSmu/U3XXMiO6eFwwvXm1EKg
NK9l8PlwrDWsHSa+Iju3aJQThY/wRfIqMRr5TdPTBF8dlBCYaMKr8hs2UbvsTt/5
e7PbTDu9KZJcwLALjpAvFeCuu4r9H8oYSMEiVC6quKVYS6J7NKdXI1FO9oYIX6Zd
sIGNGQvpAkbb6vmWS5VZKQkPp4C2xAVCCMkDSNtne9Hm0gdBrKMeMPnZgvHVUBQM
IZGqTZy7H6PhGNpgEZzTZBGTS8pWcv6unSucPv/JEQq6rsovVw7rpNq4Z+LrDr1G
Keil54YcTb6ugPt83C20BJJSedyZ2GDhBJJbJvy4gsuw4Fmu9m85uPFw1yzZLIsc
Xqm7THlV1jCHj8K4Wo4nrvSxalF1by1KiFO8b8XEYYmN93ONOzJ18J2YCjpPbAu6
z9buwBL5KzE4YSk7aP87NzGtoNuYBQHftO0RQv3A43S/ozkjPcDbpe17Rx2MWERv
OVVjeLee2YYf5+qPPS1KkFiHtIi4w7hbgO01WPpLxYkafsYd/3i6JgiNvvZs0RTG
cQJxkxQsFcOk3q2AX5gBdLvEp7rGOzs/bKhj003ClIjjtUW67eE1j97p7EJLB1gu
9rEFxXez4lxl/mRSaY4mTygwxfoMMqAzZuY0ugq4JMZl3hV8IJEkXtI16zd/iwTs
Ewa7AXnTgb7GC5WU1wyauR43GLxbU33JLBMyl9cU9ffUDN8qb0f3KPpSbDsnmMby
jjy3cwVRJ4aqhvCrSahopNIe6RgIHlMcMCcBeP3IK30wm8K0qlTBQ6Mp/mmnYdJE
3Vg9mxgY4Y1vtCbGV0m7GFab4mGu59w0C+ouIKOSGkv0OeFxbM6lMEGFWozDpJ/J
i2NEWUdblry+gAQBUdFdfHl3B7vnUkj77Pb3VLIiwPVcamKWCmB1vGDcOrUBMOfS
j1ikKFPyU5zRythg+9A8VmEYtvTXlqv1IDfI3qEP5FtiHhlpsDQetsw8NFqxXF+v
qKSMrEQsxom6Z2ZmZCuUFx6Y4qDLATEoFGXl1hLElWxG3TYOPKE4JCfk/acSdPKB
ulpqv4rnyOLyyyxBgqsUFMbLZ7UzrYqv6ibdIfMKch7lRhRA2YxXdwfy/Y176phC
VCiiHRwR1WRJAweObE0YUf2xKSGkyWFgxuyv+IL7qrY3VH/8Gd1GlJ4JBL8YRkIC
yCihPfyjbz1sgt9C3ffDBOgUvWPQ5eEhVJPIiY2wdhKI8caLfhtfU4rzdqbaPCAk
JyaeqeJiPMpW64E7COLMXEHq4KnTbCRAKcWmbuf2CaJLYBWYycRAP96Cke+Tz9lu
N6JnaYz+5SoEBKkMxnC1kvrwpzZtshjcW+Vw5RBt0mZZnqiL4bf8+AEXgqcL1oVB
RXaWGo25v3tVvyc1NnKxTK9JaGE9hZdrE3aSg359j584t3B+0tM8Rp9MVGrzI6Ut
qUxKH3mVqhP2G+sc+3YvGoaSfmlmxZ5npNTF1Jouyl6tBlauVr4XhTGQvE4elLjP
fBADBLPRVG6q2Ru+9/D9h8fVFWp79aQMLixXVidLnBY6fqjpYY3wRpEfZV1JLhYw
+p8R55ddsMz6q1NbLhSQNicLXetpsnDm/laOSyfCnnoOnNAro8RfneypJDIhZ3bR
Z4tWWJB/0ZPbBR5GmxdY0d4ftOCHo/dSOudhPFprOdVt4MuBUlIJt6lmn/0Dgjvt
Ye1Ayp2SsPFLTRatNVkDq33Cb6sMxRE+Tl515yJBcLhcQXEygkGXFP5AY/4tVXPX
TIjuODMybu9d+tLMtv1JZ7WY+brRhbIh6Gzol7ElJCZOkKDZtCutcBGpU6JeRE5e
IduUv/CJqMQT7tdMqxBBtd/iNgZpyJyzm74N4eWceSY1P9pSLxAZtNb5LCSMk3px
JSYEUDzIJ6b9/dKByU+eJp9M77GiRrGyPyMNfgzvIObj4DMr8mTbKevtL9zw3u8x
0cBAe5og3A/8oSIDaheKId321JpsdyjLVXDvH1JP0/Qj4AxtOI0J5wWLcSNqeu6S
0IpUPmhAdqHuJFhovKPXocOHxpPfFuKDLsXH4YjrNfzu+LQwCj9lFSrBaJ4sry2w
ky3EYauRe6v3xg3DsYz3FMPjGRWI2+dZ3ldTfRfJCUWCHb7snJVOFUodsSoKkYHL
ovnPyvnhdJgA4tcWWT+WcpRGlb2DcY9yQ4/uwk2KqGbAqKeWjiI6iKUtO9rdmaQo
t/+OQ2xBkiCpXq1ERIHAFE/ZN1DY55PuMGg0RZgF4uqajoy+cMECXa0WEW+5Vs2j
I8B10b+v0BGGhtAB3TEJaFadu9Cmb0L5OFXHakw23jRqF0fU3X8aqmo/ryymCxUF
bh1BlR6aCFNHwxYnmjRFXalsV8qwdoV02UHO9dZcjpwD4+7hIoFHlJLXtQ57JChQ
UtkFAQySoUhX7Bq5Lb3agaR1IPtrdCZRlAQlgDGpl6k4e8MY/5EhCB/rLcdGu0/Z
9o2luf7JTMv+I34P+BztDffzhAacof6btL2xQTkTd5bJn2oYgZTivKI6+JeXAc4v
/mUb3hE0k0Ym+2jNsKg9jTc4R/DDW1Hx/LigPbALb3WL98m6iV0cImmeDfviLRH4
Hc7xFIsJUfr1AHnNRmad4HT2GIaks+l1xrpo8q5W8mtZ7DREMgP2IdBzZ3bNb1BP
sTzBLRX9OcR6K0hO96udnAHZazJugxNLBRHVsOxCvPuBMGK4lKKxnI59S/Od5eC6
IMv8NC7o1YAgshHN8RumlloHsHlNLkcqTRO6OHwCtVN51lLMpPLrh/Y98tmKHdQZ
vF7QE7QKc1I4nRxf+LJlmgeNaxXSYCxoa9qzUhlX6t2XCssKx+O5B0aP94F8Y+2L
AHMACmfcOS5b3LKWcnTw3xksZn80OHncD/ODI5MqES3NZIrlLbsv5xz4moRmJ1iT
SLUu+q8ss/GIXezMUDiXKFGR53QfXNkj5IXVuiMxsNF385W/c3/oMf2KaLMka6nd
a+Qg4wH5w65frDkbvSjG9t/hjb6aowaOUZWrsfVbOnjBzoW/4VHXVMvn3BIZe2/P
2pkly24uQIRS7A9+W5k1DzSdHV/01WbssGCxbwZjoF6yzvAC057ePlWarHjuwFkX
xhNnc+G5zu8BaMxaHTzLL3rq1rfdCB9C/9twu+9NHhdr0e/Byu+e5wBYjmKiWXO7
rUwpRw4HRfv4YeXCMqe1aHyBmg8W7zHl0wkPK4q2mUFWJvHozhuthAl97j49p1tN
dlDoQibY3Cjg/x/TDpBVb6wt0/0Y022ghqnrkt5zWpNZYVV6cSBMbSSPQz2fUloU
X30O6raaAP3CwAbFcfuSoqOJ0xKmf6x7/kKWlezxdi/cRYUr3YQ5WjE+JHRrdpmz
jfee/5eiewhIMbr51CA+Tnq2rlNSr+sH/GpmI06JSidaXeSXSy5pHsAjFNM5rpPO
94b829MBwvkXjNY2J5wdIepqCIEvTsLJFKc8JhAYI3M9EqQ9ZgjXa+QnkJdto/LX
qvR499xIDyDJbgS0sY+DCyOuT3g+vr8oCSjwvjRZqEKOLDSeGdrCG1IsecIqrdAi
qv/afbHZgn4iUg7gBCU+7zOdpPEy19GedcvuL418Y7ExxYOfAxux5z2fOLQ8FNon
aU3S2FHNLb9SE6Q3gHSNV0XYp0TfVJ2xwjdLEiyUnZHviyiVLXDKCcUYuCrwVVKM
0N5FCcAB7/JN64wBZm3DeYT5Eay+Dlr3XYH4WPaznbb6i+x8EL8DSvklLM59ELKD
xFaXRyzqbinOX98bwSAUenA4BBtf1Ti67DkS9AV7mxXgahzLT+unDz4ZsNcIY0MI
4gX7lvfs7fcR/HQVyN4nTjE9S3F7NNdUV1PmHEJwfDENQQJyoV4FOQ3o9SmHN+Uw
+2uMVRf2zSS+KzDsyHQ+Rmk8m5RJHcl+w8iBv27V6dkqFETMMhzQfe0C+VDmxyG9
cDgaFQfznQjwP0GjQlluU7MQrSWg44vMHrPxOVfgIBALXdp/hd2FtbiJDC2/OuYM
5FhQ2VWTaTwdH+Wtg/ifMj9oKL4Kkw2N1lcs05Qp5GxqA9XSCBGCkl9Ghrn/ZBBr
d6uYZkcVvWK26M+QyuY4vtQT9Y/g+NBf8N82YK7uHdtaA3QFwY5K02o4jaMv8+Oo
Hma4iagPNu3aDH8Jfp1bRBvxDX6VX/pLYihwscacgvHKt04rLelgpyM9VcErNiM5
t6bRAVbIIpBeCJZGaI1RRhLZ22/NDi5XAoLO/5wpz8aommyuvejSLQHBn2PSjcIr
S3fxP/ijeSJhWCdOOfya0hlTOcVvCaBKicqgCGD5s18zTcdrfEF9kUbE3D0qXf6G
AKBgSv3raJ/gI6Wym4VueX0NKHB6V2PdHCHqOdyAsMk8PE8G0rSpQzk4u471JLLl
ZNkj6FeAwNtkBLIZECSrFKIZMkJUfHCZWCEtjr0iIiGFOz80RoNb86Ai1H3YvuXY
kL7VrQK+1peQ1ZRMtw9P5PzQVpBBlojQ0GUdPKrMjdhFtUbxtaCY+3Btg62thMUN
VgBEFzizZsKN3SyrvstVfYQIlWy7s1pPJZwZEEPETlFDhHZm2TLUnSHFAbqucETp
QGnYWTl/acStYjn4uhzBkuqxh2Zv7J5hxVDbn2P0yKswmDrpN0QCO8DHZbXFo6LY
JH/hpjWI8qF9mztd4DYqqntrfIEj8amDNpqzw95UmlhfGoC3Fywyr7H2+HiZCFnP
ceJJ/c0Bz/vQ/TCrihdMWTFp6wOZeHzTGWN0I7OSazvG7NHNkDvkHtw9fLgxvbSN
gmwND54Zn4XmYGVjFyNPdMUlJOUdXL4nzDCAnNhkuyCbpyZnruQLE8D4l7H6xuWb
OT55QmAmOy603Y8r2KUVj8+GgykxfnUD8n4yXpmWg9xkByZ9B7FCIRymHIwia7R7
OB+lpsWUMtAbE0mSXhWGyru0l4dLDgiAUp0irGam6wx5CsfiT4Rthvx9PArb6OMP
22mAToSXt4l7YTNbaXn0+WFtxTJhcvlqMMSt1lPl29EX3yD2gWdRwTwtBczl56FV
jAqogP3qoAHmgRr6qopm0plPohhYGZsEy3yTDTdTA7N2SInyO3MrdLKwtoXH0aK9
4nKnvmwBwiRYZy2pbXvmi4Y0l65d/eaQ9jwuTHCEl4vEIM6Nn0mtYLqIhJL/zdk/
KyqxDd6IAiTDEmayxSgY8YTMAHzZ8vTFzKPZ9Ba+UZtaKPadaOKuCzv2K5UWy+FH
1TvIURuyg/xnrgPidYdt+COA/eWT63SZ+k3n5v13Tq79YSF6J8S/bRIftbz0diyf
iD6fc88WADIAu4S9vPl/0WvKfNZY3G7GjBUXW6MivH9MgMgpu4J8Bwwwp7/ZCS1C
8Ld/nfLUEncJdW04RfbJQtQGjlX5eHOMhOMcpQlSiBWk1o+cY6DlpkD10QiBxtw9
IsxU4lk2vbVurN3zOHyhiu75bLD9wlvL8y5mHjNdpERkjjG16nK5s++RMq8G+Guv
cEDv9/C2pm2ztWBk2LPnPaOuiQry8KDNhMGOKmlPnyXWObXb8Gke2/s60pMd8dlt
/G9dOZQTpdjzYiWFtI7QZOxx7v8xitqTDw57D35s4qZthS9rKHbiI/hgLiGaskm4
Gi7AHjBmtyojvNR6+RyKotytRgBsdTOt3dx75CxeNsOGQlCTG94O2H04nERO+u7F
7EnezTKjTXL8VWskYKBDEkeQXKC1zVfFeHHu37RjZgDAvwHIX7k4CNjV9IW71e3M
/+RXDOs+tro7O1Do0KQmHpBW57nxD0sUf4Ixs0x74HOqC3+Grc/zuMjdFf0dgwFU
PeapEtAZutdo1vmMphPumlpEB2RydMGoIyffAcbB0hBSlsg06ldnbseARmB31zjy
qzIGlpfuBPtUSb/Dc6rQdduxlJBLsZqDbuPa/DYGgNg45A9yldmPl7cp2WaoBLJZ
gJKU5Oly7zeSWZG2Gqyh3e/IT5mZtcuSuA6so5lKbaSMZq1ksWMZAR3s+NmKEjQF
lz3dXxK6RyAke1RsdFhcRRaina7o3liFTQJzhoIpT5hhAfSfaTLQiQOw1+AaqsY0
DeHaozhEF/LvcXlMFdeyH2tRJr+idhPHTX/NeQkqWvPQQld/qFQVIynBcxh/Ezq0
IIv8yoRIA7wINaGwagLlTiBiw/JP5bZZT5qSMU0k+EOE9HYNTHmvSiBwa/CR0g2W
vAsyRwLsChXci45HSHkwhwG2NrkAC0MWyzlxSPjNCJ2igUiQlpV7/MMonnFyGi8w
pgOAgVtVgn1fug4oZDpQ0cMncSKcQN51cAmAZEKrQDYk5tr/lQXnhS8xqpNn+9Pc
raqeImPIiv4IZhtc05gD5o/rObN65UvFHAmctblKI+PiWIiNzAuWeLDhha7IjjWM
U5/qXSulFzC+Fp/nsUZvxKnAUXYUpl/cbKcX+W+LanhZxqvjajwKP+sJ0Ydsidvn
E5e5gRm1uuv3O+Ik9JMyyVtIBp34LHGjt1Sm5FfEM8BWBAUkCK12lBBDWLMW3arQ
gNxEgD37Z/XxcHgxB/2v2oQLKlPsEt8XuedtkqmdqwJlvOVr9ICyBY5ibb7wfwR/
nRLoRqhWuuEWqBrQXrVzlK5yBWN4IdH+s9HSGR+U01wDM4OkePfbh6gjR9eZanpZ
9PaQfpJOnAAVR2pRWjIlED7w03c3bB69jqeKbn98o8l3JV1kt9Dn1VCiZfd8tbbA
Zqpo2YvJX6k4yCP5JhUoWqCR9HYFbeUQ/kDwcVB5PtuRKPH8dGhGf808m8FYEmP1
2/Txl+USxP2vFnjFQYPhcBw7pQPsv9/rJ9q9C/69g2zi34eJYEwc4rroR8Ay9OEs
ywsNY2TUSBfK3Vdm/bRudBtt5+Itv83zcymbxPPdj+pyCxeFQUFoeqavmkGBhnFJ
eM9IKR12uk2cBpgAKDEIzgXTfp0jPHmupEwCFUEPiUvcLdpasj1+jQM2e3U3cDdp
Zah0KwN9gShV02grJKhvkQyM7VcjNwa6PHelsc7OO2pzKtgD2z7H4iqiJIdNyd3g
NEcoFvHAPHoNiEl5yi+lsHjHvH6ikJ6D0NgR3Nh0h7Rrcm1WD9gcRLA3pNTiimEx
bnLKHsV7VwMwpdXKgjHmZIC7Pd9GovGm9LoG5mdAhx1BHGH4kaQAIg/vFgFlCcAM
kEscIwQ8q4fCqGUR0TGqWAIRq9FlwqNDUoPbfTJZOYcbMnhdL9WTlVf2rBEbJZfX
cFhhSeeoy5FQX5FbGpGCtjR79azSQTuo5o6mIWtohXh5htzt62QddpOCbQz3i536
Y43OzVLwAjqGfgcQG9aN70sHJUmTjXGShEE3ZFLEQoipL6jNZKQfyoN1B/ejTszO
HLsLyrOfTsZX6yurjOHkDmbGWSljjYpovAYbbMfHoDb8TOTPcNq2caDYtjyiTabX
HbxutRzh6iOg/GLNua63nPWCgTvLgqoR4G15zjSkCq3wwNX3r+KRus7xsiXjDVjY
vwTwShTmegnrrzfkrgsFDMHZBKjqWRiknjxRwAzu1GU4DKAdvbjW91UzkIU1fwVo
ANuyB1EP0zIkIPH5QcYZyO6PUl5xrR1IvKaTNZJu2XyTLnrH0GNEJf56DlK3EpPJ
ekTc749ozUsJSJa8G2Ex609LzzuwR7nHdUWA4MoWKWVT/kTa8EYzZe/nq85XmVdK
A4dVF/mf1pedADY9V5jjsLkOJd2L327bdlPMo14eqjiEn4cFRQnbHyANvACTaMOT
clbINfKUqwBNwuyf8A3uRjkpWG8ten674TszcrznD9taDp/4c3jg8D5BHKhgif2n
MSmnHCMyOPKa5+gEaUZr23YzbHUlfhA0sCdgxnUFnsNDf+GdXl5OkjT04yiFtwfb
mMw1dPGdz99gyTpDZYHrn12e08W+YpUgg2lBJfAqshLMbPrNheYmVqLsVWbMy8lx
iY6DnqMeMZeLCp2JYoSgHq/kxb2F0b3Ibj0KxfrZywULlqvR6YOPN51aveomqh7Z
iwVZR7uYDSrWBkR5VlPsbeb3bll/5pje6ntO0zI6VmgpQMyrsTXtVo295o1v/R5v
wJb2mDQMERdZV1G5BQ5u0NFguT2m9w9+6UOTEmvIBNUHF6/sCxDFCQjbCHV5vYqX
J/4If8g2fSOK1hWxGC+CC7/2uR+iXPH4ppGswe/lh4QXU7UQFJL0xrXI6eTsXwZi
/ef6fB+QpuoRmOHf7mosvTLzQE4nxFtS8vKC2qbidhnLoBxPTglnwa0UtbTYHT97
qgYlQ3R2ON3qHzWMC9jkmrUUU6KIUXpt3xp6AIvI1KvVcvQAIKTZtkFysvznJQ3V
kq+KGRUHdOrWf3Bo8QcHDRa4MSFK/fZTRbEjHGZsMqkXXzGGOI6z1Ushh3/7+TCh
SVSkTGx1Fi0m3IBlrU6bTXTfNjy6WZl0RGCoTXc02jwioBk5/Vm4td7edMenfEcl
Gev9zz19Tx/aDbdRUZPr18MRQB7DL+FBK/AnOZ5YEgvneZMIo1d8VwQBCpFz9cal
2WKh1wj1x1jjZnbXrMZjoh4pxR6ggdRKedrhMMIamD0OBOu6KEz8rf0OU4H00HlP
2EslOak7c5k8UoNS5eeC5pBn7iOSCSVumtZedpnsGlfhFUPKdqByDXsj7Zw/b+CY
7YJCawossYja5gYyIJxJnUDMN0WmAzT0o0Me2ug7Lm1w9FulMoSIOqyB6Byq13WC
jDdl9T3jUqrO8dymu+kxLTq5TInUT0ID7CRU/kyVI04aDdzbIwINIKi4X/j/39W6
WpNjMPnOD6fn3Og5T97IDdo1OZDlFCOBIQOIV9/6S3gaUfCnRBtr9TmHeo5n4gzg
KVPeP913m897AQTT9W2Zhtlkx1U67aFsHnsrZoFDJLDWwHUM/+fVXlx7bcx2/YSm
tHJEh6IgyJ6Q5fZdXxSeXrUc7PwLBTfKSAjac6w+Z2rA/4P83f8nCT7qRrxs80Mc
ZqdzldqjbWGIXCVjfK/FnI8etVBEKD69sKSC0N80TUtXWHpoS89dCuDnslBtu6Nu
5VaRPGJQBDs0uKZ5MhQul9Yi4Vmzaghl0OnjWvxAdGYry1Rf+WU4N+/PQBjHwtEm
FvdJf7uQ1sLM6yEfod3yhiLV3sM1SVEzgI+d6/ph9AmGHf7TCSSsXEzbM3kCbujz
uP+2oCgP+V118tYYW9AeAEf9QGy4Sdkg4DwD+9rWj+HczUFJPDVIgLfHLZWDBwYu
4wZunkC740F4w0lvYeOsf2AgJcJCBcC88R9ehC8S+aAxF8GARvTs+LhfMwkLRV+G
xB3wCjE+z5ms30Cn5O9fYiWDreIKNFLNDMQCPn2lDBxrR42suJc3lI4lAaDc/mbS
j5YvQ3km/sR9tQxKMCmeHgoZOTxEQtD6f12AVVCv+lj3ejYXdtCKIdFnvAWMrbPf
i9BdvbInnLA66PXF7W74H0x2S5n5npP0EvfhjoxsRUmqojwoeSwr84HguYJkOL26
Kf4+pipnT0AYmxzCLx59+JwQAhrZo9M5tqQtQzGkFrNPaKPCTlxv+5HPgNLqWcRi
v399ml+Iz/yR1uap2PNml/VJzWUu0nIMQgvIyz/EarhTFOQ5Xue7bjBIhctabsse
gIgmcx/tUNzSwM9Ct7kLVeU9J7SUJWSu1jp79G4K1FQzNKy9scfdMfMnEaA00qjK
16Vk/7WLFMtkCN6m2Mr+5GzSjMQ0vsR59YcqDAPD9/Fs5m8d+f81SuV0AEAdZu6/
sx/S+fhsHXrE4TJRFk5I8pw2xcZhROoE4ztuLXrPJZyPHFos3x9X4U3xuc7P0VUJ
JBnzNjO5uSvyZVikFypkqb/fDFTGUxUTnrNwRe3B3z58E3Rf/gBfmrStYMtnrvc8
TPJRJAlzrvNZl8ll/HPwoQnwMOT0wmga7ZVpQcWiRYH0d+UPkOkzX1FijWES8sQD
Hp71kNYpw0bi0TFosprRw0dOZu2bMPqJRAQamT8a+IYRntkC5Wdi/MLp3lWqjIfT
rL+mnhoFltxNVEUTvKt8lEhwAdt13whK/sQVS3NAlJGW8Mb8NaYmgKnRcabojXSU
xOvr+UHMrV5Ouq1SAo0soLoHMU5Ft6j4H71oGlNaakCLIIZt+LD78jVfdVN6szgZ
wysTuEp0eaMQKO5suntziDM7tSobRUJ1d356PmNgIzbNTegBpi8jabj6nOh58kJM
WlDZBP1MVMZp2q1B7UJtPITxUbizPmPtGspjB8MQBsoD36YZ7DFu9OTJgydif+tC
Ear/kpOjbwj6gkEX6hvD9D6WYZkSYJ65Zxdtz9UONjD4zTJkYE1xncZiFmVrBEqJ
5FAIoafCvDGzHkSKuq4UQaHR06nkUxTNvicT7TXNHhqUkp09mOVOYpIyguZ5H+mt
u9uRmcmpyRCDEMkYGK1neyA1pye9uBJxP4tbkzn4PrhJh0WLQZtY946EnwjaMn/m
yzy8RjSd+SDjxk993yNcP39oFti+h2/9mPWI0nX7GsQwWBgnJVZEIA9NkyjaDEvo
PjB8IW/ELzwSLJxevK0O+KMJ8Sasa3T/F/fXoWVKU3+HikxZfI86VVGxdqFciANA
nyPMoue7tpn18BioxDhxQgWr/9IIr7K1NzuIAot0Rd4bs5+iYk5X6RE2k9gcRe8e
vw+xhSHxYR4uhm72ME2Fxh11j0uVSXEm8kHBuaDmFcwfCi4SkTFKF4FK4+Q3VoVx
OVL/wYTUu+H3ubLXQMMsj9mHfypc7XhOV5iInKJWBI5x98dpIb/On2XcZ69D6F2M
VECGEOehEBoD6o1wd3RGAA0v4kybxFFUnkb29SKzQzF6vsbMAGG/4ombRxGQoo6M
OzVd+KaBDA1br5Zqjf4imHP61KXnKu9o7jzF5XjJZsRDruAKqQjt01Sy3KWnlBhD
ZA9kbxcp66KratYQ8FwXa0yAKFFF8xx3nl3IMxUhyWGQJwJMJAWL4gXbvv1J3NqF
FHVAtouiDmSxlncZfu4d1ZRFaBqAhTgV605dQDTZMyVn166rP3EHLRukk91oijTb
akuDMrosJZag6Y86BK5bFboIlA6S/dz3gZY1Xhq296qGkvExUBFYGbkr0MR9uLr+
1bJF6QvILrJ/iNin9Nm1Uq1vSlfa0cVz9uGvNlm+z7pg0gjyR33QIx8z4RgOf87o
2RredMkwIp5Er8i9m3U/S9BVG9rzDtTa+1xsXGQr0PVeXnQs4oS6Tp9ifisxnkVe
50/3CXKNo5iMGaX9YrqMSrNw56wF4LckjlfcPwen7pWXce9+ahF5scDSmP+DNeKq
hnbRhsx27VM/Y1tGOJvXatWktr6assFWDE/NLS1J1g0LfIZ0SJaY/3yJzLUE6VvO
PgYqTn4Jh1xl8zOnd6b0mvml753M/n5vUJ8chvgnPvT9NztcVTM/ESZ8r5/nc24Y
JmiWMXlh/4maYAgQuZ5QhEAQABKip+BU1MQJp47G050wm14QiYXyFr/zrEURIWx/
al3wEpjlT61Hcysfs7htSBNJLtfE/zMy4dW/DwGHe5fqsfNc06rGhVlmITs/AtWx
3UTP1oVhGr6M+0bKY/SdOv9HsFAjNQQ1UdT/u6hdBcwojpS241yzfnj+l5TgCNVv
AJ4AJc3mQymhMOolfqzxIK2wno4KetpoS/U23En2lbxBUsqjdhpJcpepaOK4FAwO
EoErgnG6j7W1A4B5Ci2r/vxgMlbim9ZmT/20nuNX4WGlVtX4nk0TjN074i5rHRPP
Eeh4my6Uoa1BPKu6CkDhPy0NmIOMkTs3/dCBqceWkJCuzr65hZMWz04mgCzyNgxb
UOU+C/DgQZBbMZ86Gfdk3elqx8PTFn+MDemgVgtM0EbAKVa+59BQ/r2V0s5KKV3/
KRTZnDZYIulUyJNSwjvdp7HoKwxZ41repZIEWrVfxnCr7imGDDqA7Iv9Gd1KEDhl
0k2zhXqqdoXAVGiG7Nnol6ACyQ2j6J4n3Dy3GUK+Mr7spJmEbNLi0kV8krGaqnUr
/SPdxmIO/TTLCPGaQpt/WK8dXrH+lGZ4uyw82/M6qZVd3B0/w2qq3JmEq/cBy2Dr
gzCSOMpOmhsxlBGk9qK0v8185nRWYSb9AwliKly/rFyI6j82xo9XmsS1VAWcRkZH
dVZ73iEBS0J9UiwPkUA+6oh4dOAVq2z5oSx0KXFVjtmCgShWT2tta2WURH7FE8TK
MDyyr8CUdHtYPivXEc3MsIe38mPfhvu3W7xkve4pwmcfiPDs33GXTdXz3mMHMHpq
agqf4D8gATTwg2Eufd5bquKZjwJEXIj5Qv/0IEW7p6p1iIw9FovHfQ6jd8QBQ/g7
hV4tMLDFJ1c1oJHFadeZW07dpJkePIyp7MYx9DdoQsOhCh6ut5ttGI0n6iA7agkb
yJuOP/lTfpTpyaupiWu0eOhgorR9lT9W/MrLzgsze6dtvagj3YNprIcxS3D7RKKf
U6hPEkshHAtfvESzht/lH3kOrnoAVPo4cXWykcO9JNCe0aq/5VTGL8Kw2B/VjBh9
AtBkcWtHuPkQggmMvR2IBYYdFDXZCSERPUgsOnqzZfMyMU9COTt1ix8Z4iSkIbqX
VDu8waXCl6sLZ+tnHnfrelzp6azADH3zlkBuvNbTxA/3oKmJl7jIHtsgIWoQ2iG4
fldd8IxKqZaXhir+8tFyevMnGoJBWm1t45L33DeszFGxsCof75iIlzpJgvc9HEoc
3U1cb1q3yp++6TLlTZ2wTbIT3c9qnl9dE/FA2w4/tostJor7oDye5M50sK+jKhgh
4FtkUgOcWLNsuMnr2TpSMroU9j8a5jgjDfA69iendloSsZgvbvWNSEVrsok0yoUM
zC/9GFpINOidz8zp0Yqm3bKcB6DIcO7v9oZUgqjY1qBu6UwCZnZN1HbK2So0EkXU
ufloYwwV5WBSYVNG8ThHCeUHEDBBE45HeYQ5JdRQKr9NLf3FZYLl+uHLATys/7IF
DZidsfYB/l2XPBcyYurHkdT/XBiEnOVPZBH6Y9VZhRUjD+6R/yZDxxtmr9Edt4Uh
MA3ePyrNaVJHnAlVJtMaQ1e/yrGJAyL2cFmpzcUR1Ki24FiKkrPNmVepsSc5L5o2
kxPbmW61F4gwYcinCg1Bi8hdXzifl43ZYRogoBRULzGVmRfFdQeNKyQwu42KM3XC
5qQkriMukGooNJHdK3Vel4QvM8ZFsIqQhXUHiLKxr2BfZDyu0Yq8DhhpYM9f4GnF
yk3BShGu/p07OEcC9CRuD2BwWTkM1Q9xRZ20L8ZGrWMizS7UomQM+OuRE58X/09Y
qWp0dkjcjqa91odmkMk5DHpIZ6NwhtGIOueR+lKWip4GP1s88+oYR2RLEHoruirU
AwYtgGJLxvAiM45ccuwrJeEKqOa/sVyDqRKb/8YVbsC+UQ2eKAbAbVCyIkWHrHJu
0gZ4L8i18HZGS7sPVtc43WDltnsgtuyFepCn7JaYtDR8MGz2zkuN9XtF06lybHrG
tjNK/9r8OtwjF2qXYo1al3QWpZKYJW7VbosdTHhaMX4fKplLZWuxH2CEnvz7pq91
nmTbQIovpvE7+6u65Zm45m0d5EetE2xtP8l4tQ3SDsY0q4CS6/dKbVkVCJMcbeEU
YUf5LhEfJRQY5Y6W7eFzD13Oj++SOTWuC60MB6W7novqz2QzIcf1eCe6nwj1UlJM
1h7k+lX2QvFOHHfIfYePzWOFee3M+aDcwd3MprXGmUV0krRnBf92+GVtyVHHtB+D
2AU+zVnHj26fJiSVdlYP7ZnYE3mMzWEx0ZJBI/0cXTRSSZl8Ws+RSJHexjNZQqb6
+3lDb4uoaFGy7AZTc9DYhdDQ2ihunpoYkEFxbzlOyXIxaC+GDUedMY/kR0ewp9SZ
acvTL4EMJ+qFuILFLK1NT4/Fh52StTR+EST1djkweliVFF9NAeEUHxrUYvWUp/G7
4T1wBQZbIlt3YO/FGOc5sXQxpCo92k4IFEBWh3M7xDZw7LZW4E/StPIARhq/wsxm
TZ5IUMBnZD8QAFn2ekIbtLe4TVG53RTz6NhABxfF+wV3TnwGsxxhDZjdcx8kYqzW
nqhsHxQHARdhWItXPeb6dFa4lULJepjOTS/T+LtUxQYTz4nsL8OKdGg0IGEBbC8c
0KcK/djPrr8NvGB39aHl5Q/UYD1dWHAWmOjxi0hW5gCwseLeQMGG4fMZI9MLpDHu
UsJMB8veHjUBlK4WZTtiHJcFsPrtppuJB1XA3H9nkV5AOAnMwZc5PULBp/w8939A
i0yD7402bif7pnY/ObY1Rw6fs8uihZaTV3s1AxsDRyC7tvippPkFX2m1o34+MlnH
uRrorc0M2es7I9WFIk7gJ4rdp9k0zSNOoY5FOjqEieE6o6FdScUA2DPKqdXZ8+UE
7qRCI4m5gxt4iXkiW0yN3Umu5ftbMiJR2EsMYUGjnDxgeSdqpqqIAITK6mRcwKcj
HGFWd+fmsZEWDtMZl4GGBGUG147FF6mu+4wwzgjSrwmSGq06Om+X+lCAJjwADmDZ
L+SU4CYlCGpS3C3Wcn4Pa7lw1WwIxJyrqWFZDe9ZAiW9eT4ruhNHa2d8PAZutK52
RoRlPD7lLQSTlHkxQ2iuqNHR4JaFNK8+J2xvmxt9PqO2cLaPmwJjCgEIbp0VzJe4
XylqaTvhH0YFK9hXSQmDIT6pIa1frtInpy1y56an/FEOvktLQKdBTCzBSwO8D60u
ccJBvl4Za9RXO9Vc7i7eFRF12XiKbCuELaSf9Ljdh9z0IMWz4fHk+PKYmvE405Vv
RnlGvUmtUVQqDAdGd1cz7w+RD06gcYx78W/6v9q2e3GryM7xtdt5LzBYC2j5VOYW
Pu/37QNjRqr8xD4Qb5yVdcQ3wGtjUW/c1SJcKrLXAG696Yg9T1KsCfTdl7iomN7x
TGwzG+BAoVOJP1QTR04vLGfiqeoxXZh6YZCoUQTidGM20oygjWa7E0cmaJXh8XYp
DB7qZBKLIMmTXMMfPGvH99gUvUAQqu7PCcgW3YSfWuu4XDA/uLvCm7b7xIP7/Wvf
9/TzSYCrBYon4NwgcDb1t2W9NBa0GAh1nLSznOKFYstcHy9FgQ2sm5EcQNiRe4m3
cpgPogwdU5CNxqi8wdZulHHpfdGIKaepNd//pTOZ9PK0gS7K0Fk30XFXuMBvnHzA
thb/NlRI5VbTghm4+6/mGXaQiDEElg9gpqjxBJkO/mizmpDW76KhT4Dqocba+uIA
eaI3eP8eeEZttNtj8n/ebb54hKkcK4tU29o1EXJSd+GC9SOMWmwHjWgVfUzrW0hw
yepIKzuSqkTc0D4EFPb+dvb9KUAqdQ/+J01JOEem85+olwAFZdP62KjHAyEFc8fZ
2QTEMZshD8UG2bAkPb2OiDwZPQyfFCuCemcmsgvloKMiKg7VtPdqRGx3JqKLZN/4
DInXOAdnCPthN06nGpYVSptKXuWpwU1U8fs1vWuTj2O1krRIVY/ITMxX4CybTVnI
N5k+dW9us5WVfVqyUAdB8y+lH9MXzMFguNZuJHtb/b1kWLiPvTFQGKrxeFpgjdMY
gb/UEEu4dlx5KnsYWKX2OP9yPF4vTE166FabiH0eJUIbYTP0f+bPi5J7t09ZtKqk
e7tDHBsgFpP9PFCEjzkbUmM8/sopc/RDm0FaFqEDW9YkgC1MGT3qEQzrFp4mgRQA
1KKlFaBh2+vJUrS1bRhkv3F9ZB5h6GFB7izwyST2Ellnh01XSke39PC4Lr9v28Ho
I1anSwBXwgqYZr678bP7Us6Is+u3vXicoJisKE6tpZrN5e2gAioJ4oBBDwDQCFro
9hYIJrWZuG1OkTtlzTSA2bxErx9CKUoABm+Y48FsjDFi7dpTN57lUPeEmKlXzdrx
rmL+EYVX6aXTs8Y6FvYzt3moNZaU5O+JCwPEmmPPETC1SPQOldIU8rRn0yyBBchG
jai8wpRcnf7WZ9Q0/OByXFBYv8mreTVk/eQeksswhWA/Sk2cB+OFunbMYKXRGR4M
HkZykSQ8hB9I8z2FKqwpuAPNLFF8xFEk/if4Nju8MKAH1Lg4SzKfYrWo+UO+Kilu
i9WadDNeYPDB88r8OBz3ReOxgzSoPkbdBZ4OpWQrJQBf6dZcjZRHOOy2ogKaYwxG
jmp3mSiCZN+ykT4Aj6i+gS+xrSvNgEuGpJXDNK3Sf+cXRWiSs/KkgZcFcIlykX4Q
adaAMSdk3CT5tSuVt4uyiUocrafeI/7Nyk0bVunndAw5wXfMk+nnfvVmEQ1gutv9
IbQ0iBm9lcAsZ8lEDJ6NijuIGmcenT3RgqiqumQ7xdpG0fvSxng8kbdKkYZNxJnZ
4N/9S77rN9muKQ4TinAp6q+xbtRO+CyE7YAzlVYMT5TKzUy2wTWWGz4D6yQ9pF0H
cRrHtg9iGijzu2QlEbS+I8pJf0tnLOx+bxmvxREGdjUGFmg5Aib52phSHHcNBkUh
3ndDmfwQbRDhCm5SaQnhp43walpQKPwV03DTxmNzKhd09l74NvpbubJDV3YQ/f7q
cy4UaqWxS7qg5hGoS7bFerQ7d7v6k4ENcSQiYrpgZahxO9kbeJEVZsQ8Zry8x9gy
BwIyuMAhuRtCzbmiLnDF3QBAnRSh6vCsQwD2A5iD7afJvL0XsvAB3T/5Zk33MdPB
ryqJPFNsxBuUkFDxQk0ORpnTxnF1BdC+8+Aq7DGavEVB5p5MxFVY5jXMBDORXWU6
x2ppPhm6lEYBUrShyioiFW0hibmluKadShF7PJjfRvaCMa963tg3MgNeSTaI6kb1
Wj7zQSq6leuBD/hQHYtwlSvye36eWXGfJj9ahMLlLgWGNLHHty1RDgsNYhwQ/w1Z
rps4MU28VsYwWfoZ4euR4i7s1s2uDwm12KdiQfgWlUD3fvhK+YwzqOsEz1EA9S8r
tN0qolngDtPppdO+RXB+1hUtvPFXXe/g8OMDPPxxQjddY9Za+LqB+5OvaRZjeiyA
E2TaxikkFhTuj96ehboLM8uGX9Aa+wAax/1DyipqTR13skLP44Q9QHV+IRjAZqKb
XiRQcS9OomROpCBBy8+F/Nuw90GgR6u9pE9HYLxzytynyWM/lVPAI74hL2nDey/C
vo6Yonwk+laXYYTShjTQvwdUdyxgl3p/6zK+IbORdBvsw1GcxIV4ICHXN/meqL19
m6+KxjpQ9tw7cQ/jCiCopgo0gIr05As+hAR14WDrt++xtuJoIgCsDGDirSXs9o+3
wRfgdPkc2O+99mrbVD8nT3eM3A/KfM7l9aX++C2MDNNWIiW+lMNnRW4ynRrPRu/G
3fqpvNJPKk06tfA6BULabluUcV0qGLh8Wr29hDB7UDZQnEZ7aoKfRwlL5R6cN2gY
tujqIJ/owhEtg4Wc7QlHQNNqvihRVVCpld0Kfj1wgDSStYwntVKnwHOp6iv6RJ6R
mJxJ+O/Z4IjKIFrYC/pZhW3EBI/ZCK9Xh3x2HNK0hyxiuZtgVr5TUb5mqJWsa8ib
11eCnfrH25ZzVRflo/bx5HpwVTAmbuOC8BqXRySgbew4cwCjd5cZVU2uG0ei99m7
uKXMmhub4BMQEyM5fzGq2NzWBQ+GpekTuyT4Ev5U2B1VAll/pSWjTqz6fjrQJ8oA
KT08KJVO8fx74iR6y+WaSC38EUHnkZjlHrDj66CYBDQ8jElvpDQZPxU9OvR9KEkW
QobSQlJeK16vDnsWOgosyd/IQe2ySg38pZwj7GFzCYh3HgG1M75QYdYHtLF6MtxY
/k4Y5o1MBAbSEyRsO7RUx3njoYRIi+F2KaY2Yp16SX233rf8Bi6zW1UFgbImsINP
axLnx7EEcjY/ZTU/XJ+nObcnDJhQkNn2Da+6gKX640CQ+NYQXkMZdNZ4Z81b2IBW
9d+yNDP9Duzsm4mM0aqiJybYChlENWAQ0tPWdkqBMSiS5l+OG7u7TmYkgdcv9Tfq
5C7hf/6p8qWGv8rlLosCg2A6w/tqJY5qvGJ3tl6VUwbHSwCfCINMHr2vOfq9MHZ0
ZZqeXSiN8PLuGY+qk8cHjCqISIHS3I6G94lLLQ0PybUm5XFybGrPMzzIhGPStM96
RD4OSYTV/db1sSZi13aNEsyXL9c3vuS+sbbXCkeknxq7/arukWoOuUNT3zjDYea1
yDvu3KT4Co4e6DXjhpoSU94TrG8l+KbbjDHibPeWg2//OEav/TfedDqDfQ9gB+3I
ZPfFtpK9re6I07Stxr2umbTcOO5maaI+YRht3Hw8jUprF8QG4H96f3edyM+rBup8
YdGEXjfy8DUT+JwSpMhK0yJWUFw40JFmul03nqPwjEEBwEEw+/UNfL+m8MfTsVLg
UDMTDZWX573U6a6VU2dCioZ3ShnO+n8oRAPoQlOT5O9n78dbrfVZBB3CET5EBWIg
knW+IpN1RjbNqhV2diKJ9socv3l79+ZOoZhBl4UeMe4l9Zz1426O3Ss+Ysmge+H6
uxsfGzau3K8nV7OlB3rn4vyaGdrZ8RMWltLjRBr/99SFqrkwKJgVZY704G8YrPfy
RvjYsriT6fvg8wK+lrCduxvtnwstQbJiQcrb/Sj41VmHiyqGzV8CwndZYavwLaxE
nhI6lpeV1su+15VTdiopnCmjs6jHTfFRInUwm7Qsn+YSGQ/PU2d3IwPdh2Ch//m5
fHUaz5w7Zj+zfkgwdIck9n4y1lCHkGNwpp3TRY5J6XHdGbON0yIXLlCVjf3v4ROW
c7+gbmNtlb8PQnphsNXKqYN57Y+fb3WK+VC0xViwvgoLRDitbfEmO8LHXhA/F2j/
RGm1fwpCWzwFHyKRL/dPnb6ytKBiV+GuGcYnJjD8Dn0WQRODTvmTjcfMRbmk2LKq
pef+Wdv3+UG4yJ8dYH3OSmNTpnIqgqcTUVTz47r4U2jfP3Q0oYhsGSqTEQ8axqIX
o2wHxP834Lcr1Jn1NLFiZSz+K+9ODhw0EnKynOmX+O1iy6ftGwtPG53k1cVdDo+g
a6a5HNjaZXi+isaMi1tR5TeH1gJeqVgey5wa+rU/tADWbij7/qaM621UceHyNmxK
1p4BFyLeJ8k8vgPgxyKkoYSBYFcVx+3sOvMbwvKiYAOcBheF3hdhkvbXII03BB+B
K8AVBGQd5zQL8ykLXv4o1BlwbbThObctkTV0EctqQIVR5rnNpJIaZYVK2wpzk1gs
vF2W7IzyuBNtOpf/AVCSzapdigQ7C60Oegi5PRX/UZBPzUkC2n+Du16yzzmTSvdt
MWBB1In6ys6ca+Co+E3VNqXAXR2eeEZxXvNFfsRwiJvBergDK2kN9koCuAuy/ArT
eCHN8v6bJ2eiz+zXMyZMeRUGmwKnna0na5RqCL7M0SyyOyGA54KMjYy04qamrWM4
jF0B6q0FuyAU4U0XIC8m6ySQw01HNGSvzXhMgjqG+WJZ7FeNvaynkN20pB04T9vW
4LSiP/m/CbcmDdkiO5vbTwkrzXl6hKxEZXZR/hoX12yUMwXwoh08wu0GO5Ll4lyl
EdvzbFubby8pwlKF3gNJcUcZBsjmE5AVVrZ82q+UbDV095YTCG5OFfPdxvinqbtV
hoQIingKO9WV3F6KHim23Y6VJ6r03B0BIxePJjazJ2Dl3I1ZLQwplCqvN6/EOJz4
xE81YwC0CBO8lAqfA4RuRTqqzvoEC/umKKv+BbZqzzB8Ug8UFoiLLhTQTGU8jKkw
/p89oEnPMg95jTXzTILF+bvSe2Oa8ptaGa+fiXA380UwVZ6HTlYW+sFfSdrLQXYw
jxxkRiIOLdPbNczQKRiH+Uvkw1ZgvzvzC7ePq6bI9LhdU4+YmbRavaw82EbBT+3H
Ff9pq8Ld02Y2t6Ae7z64MFr9Bwu/Rev6G6nehoqhFKgAkqXfwSqAy485SlvEq0lm
WaMVZvThwCB9MRYay3tsq/xzWj//iIU10aNonPf6k8iuExhM17BGHQCFnUn3uvD4
BJKE9AQQgnTSIjYxNj8XpTXmK5NLclNeAsHPMbLmXOSFhe4tVedL7UdXI6xXahAD
Kr4qtYFsPMNsTEAKlbybYwm8igXoKY4b0l+y7v/J+EsOsfXWxIjPYX5FAFRb58wB
JZBeAo5Rf9yZlkqbOHItTaTngzddRsED4d0uNQrEiJkKW3Mas8SWPAXEIbLbajwq
r4rcMHdRVEx0Tz/vgrZXzMLaNnMXgb0mpPSKHmcank/LXTS5bKOjaXkBZu25mkZg
Qzd5Ta0qHg8DkupfHF/LuyBnGgX6A3qzaCbd999X1I/yySposjamBy9BHRcood+F
/qXqdskTZSpZLDCBC2REpaMKPaB4UuxSgNHfpKYWTx1zrOSDJ2izVpFqBfeUNZ0N
q3AEOUOooO4jFOrJrlpc1BZryWbSqyTMiukqIaqNaLBOqljB60i938cdOAaT74l7
QWbMa43HduzKdk+YHO++reiGe6kv3bRjs6bfU6xTVSFPNMEzHSdebTrN280GaOtW
ShDB8KATHtNH/gS1MkwC5eBxovy/3CK4FLbFojsPlEBaukoI+JzIc/8wRKtinRo5
hEI6+PF/BDMXrECTpSfwS5G3avYs5N8TDYsdJnH2qB8WvV2LevqTbIvaBLHYvRqP
Aco4MIx0tuk3MNIT5d5ni9d/U2MnjdEJojPR2dFhziQ8YwtBgK5KYzgM8B8pi23t
AnyzKXOiEl08QKoEU7S8h71i61mWkDHP2WaA+ksi0zVdxNEsOg2uakB2Qp/QPUNJ
9GsqSQ72YMijAPTvcaqDG+8JUZd4ILgarzqluWHm4tIeGiXFiWpABx8GGBxW1ykJ
VJjXnOcFUZpFTyg+zbL3htJ/m0NqSjOO9OdCeO3V1/I56rNYJw+eQSrrAGeqOpIM
1ZNZKRNP20y4XYrsylxUxeLSb4sYAmQTTPRUkstMYQq75SglZUHTpqiMPI/DuOeH
aBxbpvkqH5iO4fnyBVu07WoNoB+YoBq6TSJy4TQMWqEiO9F4TC7U00mL0bxrATDo
QgeOA5waQoMCJe9fiFh0zeCXR0/IB0Zrxkx1I8JFMqlRjGlvr737xlc171E5rUlL
DMI/7T+J2BGIfJGRoq3g4q/0MgXCR8HnzYl4oxxhc05LRRmKodsnTdh6F3LLGnYG
wdaZ1FVHSawfdeZ+s7ZrTKH/5lZAi6dyqXGSVvuAq14jqtLI3N/P2h6OP7xZs69K
hYG5uSKQfFSZgtIfPaJJYRXQBLstSe4GQG15F9xhDRMte70fng9fWK2Ku95A0Uvx
dHwx9Bwme3UFRpwWw4V3K8kFsWhYFEc5R0tDSVWK/KWB98GuX0EnN7y/YZXUXdSB
ahqAdOmh0NbTVGXqE9/cO6wq4qYqI2p7zii8BQidUG/Kk7Vg/EGfyVbRtlTARpol
VymwND7acXsWoapuyukufrFK56zU8NCdn/whPqtC4+hbw7GH4DN8xfwNX8Z3qhtY
kvDrN8/CRbBFS2lIOrim0k8ypXScDM8phTfBuYI714g0VFkp6Hl5ESfWM5KH6mJj
vSqW1YuvpPPuoB4255DFI8H3g19RhPVAqPpxcS4i9VclpO53bAqr/IjrloemTSIs
RZnIANzmDvIX/xmoB+fxOdLAoD/TSgvCN/PskD7GjUzf80CAdyCD0I8P6j0dw1B2
ntSxqscwWvRc+4dI5PYYVTUis+VB3BsMR9jL5dSPdELBW1OUuJjkrLV991IwUTqv
SOUkpyYzqHr0IcwhnaL0agwsIbLbmcjU8pcBRtJ65wJ/VOPKz6sLhJzlhE0g0cME
E3BudbuT5PuXBT0Xzn3EOFz2Nz9Z2dI9Ou9UD3DuIX23P41wPS+jR9iBpnb1AeqC
W2o8BdR4EYilFf1qrXsZ/n/TnGIK6nyHyX4Dl2OzP4BJVARNaNofKt4ml3cZXq9W
26GAiW6XjQxYIxnbbs26Kh0OtV/hoT+WcYn9+G3vcUM/hvni8MIpQVqA2Jj09SAW
+TAghcx5mJ5lH4D4nmHpYdpPWFoi5Si+7QyjLYSAnK3ygNiMH6KeSTsGUk8SBO5H
OQTm7xZkmEpxpxa7WuxYOlmNPGNpxEPu87tdpcdhlQuvzKNOyyFUPInNyNedgsxf
qTO36uZV73wDZ1MupSbQO0jsX8XxTRMl6KrOmEf9qk+XwNl0mBfD62tC9o40ABWQ
8fuZw7fVyDYDOdzYNwAZuB53mOXFGNqf1fSGfbg95sDcPsOs7gi97xGtz1IyTfZZ
bBswbdoVQ9sfJAlk6IfmzAkFsBJ983QABkEjp8iu4isxXpdLYe6UpF3xQTToLrML
TdGbC0jvLvMwPh13vq0I0j3zzeon+5f3/9jXGZrRZfUbFTDL0DeqTgXrwxYfuoJx
wK0GreDteIDNYjyeWhb5i6FS4NkUi9JxxpAFyCNjdxpyC6ZCP5jkNQ8Ktoi21nmI
aJv4xAxGp3C2m4UtUrYmddC6acHVjJde8juSBbmPYVzma0Yv6cpHixoUKUhGn5xi
oMZ2ouNjyb9bepNBigzAnrGkGUWwq66KDG2yORk8rx/1x9IIeMITLFBc7D6x1f7e
eDCOs4p8HFpjcBQ006cvh8xpl9hmN16/6Jg73HbAehOgWjzFLd41KkTI/atdSCyU
rdM4rBA6LQEEdcNLtzVJV5D4HFRvVzEwGISxcKY3fCLZwYsAHd2ldKwrKlrMhX9J
/yaSoq6+0kK029BCnSsY+4LmmISrED90FSWJ5j5LiSJFuAC1dyDqpFBH5CPJtxme
NOl4hor3jpAIxqj/KOVBkMGr+Io3gju/9zPk20a/tRpE/d/BVZGNl0pABh0erxM5
P+fVM6LhJ31qVgblZ67kfUiLJSxE99kdW4ZxA3Jn4sVm3OuXpQpCMfpjFyxSkLfr
a/HWqnbEoT5ppqMEOzqcIdV6mV/6alwvhPTuMdOkSjYCO+DZC+lOKmXY/w0iaFnh
Xvl+4OIb4SYfA9Pt0YCGNUTVL9qMjlYD1ejnu400YBKfqJEb0cJPvdy7zOsS+fm0
MdpHEGceG4PFBxpivisPHSb6xGSmBi+D6lUARjTooARWJehIktsiy3iBkTOVL9L8
yDobnJcRIF4WX7zofXShQM3TnmYCqvfo9LNm4W121SaaO+k0+PtwuxpghsRxoM/T
C6K995XDyvvAE/gC3V6SV4Y3y3q6clHcZbJPZnYo08Hhqk3jEZ2fkJN2WPykzTmi
CFb5WyRaCyHroF/8/uQwbnEuNRyaiY14tiCD/4ORG4qKOFhGm3807nj6Y4pTbnOR
F2rpZsekUpZMZwdzxvois26ps8jCqt2+AY/lvLNuiPHH7xecQUuJnDil2J2gO7U8
fbZU89CPspM4kTPEXOphCntvCeNhf5/XBu4xe67zWT4DM7d2XurWWG3szdH8F9zZ
vW1RawmwJTmBIyJ4cc/ld9AJyWlFd1Jms62jG0dbbXTYUA9w4Ty/TZATNTexlf7N
CFjjG+nkQmn/FFjxX0Z/gENWn7+C11XzbX7UANvBHW1mNce7uy5hSz68hxxpBpq8
bf9+TCm7S4ymIdx+i09ms4DHjZiu71HwPB2aG5Ulol0VtcCwkvO6d30ry0eZh9d9
QuDtdDZ1n2KxFwT02HAqu2TNd6rHOHR9EkLt9K9F84yxJTP5ZMCZbmuhixWJH6pO
y5A5xMEgkWXMO0uwzk87rpgGwwURuiUQaiBfnyL4HbSSFCt2pylSMkywUxHutaJ/
lCDZNUW+qdw/e5vfSMCISHuDXeRHbivgjpYvUWdzLehP/OFfqK+3dKp0dftD7Pu+
OlgfchEDq8ydg9J1vzHynqUa4wnyR6wQftb3OEtNJ6AGaHVox56yBFReQKCRAPLS
V5Gu11q2ym2Xg2xB9OPmNi4qT58cK+mjSQ+mSDJJJgixANsL0PtAx23LZ4bnq0HT
bE1sQKjQin3xYQdbtR0w8nzYxgaP30VFo4yj3Lm4qtYWQWJ7B+xUVKgo335xJcXm
IVAB5MTXmnnjXaReQ67oRCqwmkH/U8zslTNjdb07FlUoRi7KXyge4Q7aVhBBFRLZ
AvDOTLt1bbzQP/gTOsLQ9G6xjtM+p5lcXp73U1qVKkRMyKpUxqhJxm+3FQrjy2bO
Dk5OoMVbxr7C3xrIDXQGSzobxusKRdUO26Z33A9MhNf/8fbHfttm9jd5twOOtzVQ
+wTOezfLaTp+u8x50OSzXT6jpzvmq3rzyphmefq/g782hHcxoGVKnJFS+ZJSg8HZ
k5RJAYXZuMjIwpZVhwXiaVy9oBxCXcU3ZKYE4iYWoKEhFQqIk+pSZsCuCAzVBrgZ
Tt9By9RgkstDthUFuKiuMyLmtHeCfkFmEGFC6or94Y46Pr4dsqPP8evhb90AyaDB
7/dXmW1dFEBkq9u1I1KpEWBOjMgwaFOyMJog0Wxi1wSn2xAIC5geah6OzArQJ9fz
w8JktpaQ/G34RoDKamJU244ixrwIet79WC2NrzpmaIGkLHWqmlAAqvUnLWp7XyzP
7UKWIagVDRmzO0AhcFidzLPlUjV3/CTfAu2mTlTAlDoxyfBaA+yufgIH4FWf8VBe
YDGyy6vL7U38sSpw/Y0pk4Eh85X3xhiI+QNyXuiMeAluV8yRUXAAdKZRBAwd8Ouc
iq1Kd4hc3ORWRPDgbtNNeVDklYd1sdVfgAKiBU7BQuEi3147prPhiFZnl14t1adX
IY934YBVyzXL0Y3GQUUDUmngD//jgY6fmLhCUDDi730MSWF4MakmWPMDYW/MAk9a
zSZnH5S7uX8ZeqPJXxOaYu0+fW0M4PAcxHWbqhyQPJNhao+ihL6MN/tUixkA+6A2
W0Crt69oP/Vo8/h4W9RXUTXGaGddij0peYkfhG8M5syhO2XUHPOPQ1DlG73ZOMiZ
+X0C7zBwwTlCE0WLkJgJy5CuRQsuEst/vzR4dkHN1rNmoKhfXC5d4YoIdnWAwJnV
uFqaCnhAFstMmaCo/TFQUQN0KguMRg/B19SCsbZUK1eAzXfekOM8rcqLIBMcPvym
y18am4IY/ZHa6iGcock/qFKDE0zs5t9uhoPTGtmXIT2DfH0gPVbUZtbcAls31vz9
Q2JHWgU4z0fBEuFUHkllGhS0T7p71yFCQRMXy/lSgPXUYdZWTRes3ENoT4Lm/qQV
5oEb/JStmZ1idrtZGQvvGpuPTecHJBpRwyGXhRaQPfTqH2wyto/596NU3zQ0YRJY
+WLYb3VrOnHVmpyaGZZQ2ae3CjziDhITGA0dEkMoY27jYZMcz284gOtLDvQhG64g
v7g1e8R2UHbHaLHB8f8+o+4zx720HlOWiuAbMo9DZzB2Ftb5yx/v8z86KWYi/51h
+BYcu/7RkUSMssBP+S8cLjN2FYc4sx3/VR2xo/ACGH1Maxq6dplZmwcgjWabZSH+
CNpX5Auzlodh6UWcDgCoBpblh3T9R6SLzmBiZq+7egdL/IfQR5BpNl2EEBXESnFW
qnQh7BPXvpPHvQtpCoOrlCG9V4u3/GCsySYWd0nTDXlYnW6C6+bEBPAErwJEIaFQ
GGa7UaFL7LuGmoPfCa4wn4HHLPKhEXIqCx7RL3yHfL4qS15xlt1i+RryQmLnriaG
c9h/VW4+gHIk/LKM5Vt4FOvUJ08N9kNsmBLcFyIx6oJIcZ5rCNHcDH37V4r/m2GI
541ow7tM2hl/2ToqVvDwqSeE+oVvC15LCYRMYnM/dPGGuHe3KOQp9daZBGpiu1AT
r1Aoc84UupABhLeFO3GMRO0nJQ/UuzNLPQlaLmjNj+fFwIBCpspBIsaF/pyozRxs
5LcqfOma3ojA22HP+LojAHshQsLsT4CmjKvl/djC+UjPzcAmTryKN9aD6OG22izn
wMgOQKBszBXGgOr+Dwqo1Pd0zhkeSAxxfm/kr5I81YI7bQa1Wpe4t/cc6QAVSJNQ
3gJVTzMYkAU18qC/ks7PjccFAY8/X7uGbwyxU6osJTUIzoSIFv4P2RAIy7x8PSWn
nplb9FZtp+7Ev3F8e4pOyO1kjV8SOdq8PpsoDRlcqyMpXhIaYE6vEvKLNis82RBq
DtGrP+24BOEaVMWFLhg2FebUSUcN190OdloTV0zxETBRK0WE3bBabEIo7zDiiANf
MB5DvuWJxOlAPmM2DijbA/olTr5uo1b5VYfJ641HAdESKoj4TZvFqfgB5HXNLVkm
m9dQnL/XBSR/Uc4OucqB6FSiPZEdxbmA4LAhtKVBLfbhYvgeT/Dnh730oPDt+UDp
55kz0LnA/8CCm7PoidKUyHbU/wM0Lvg91MB0QQDuqlMNeugD4ZIwJnle6mPYrsXK
o0ZgaCsRU6cUvCGpS8ywe6Ulc0rSNPEkIt5uWEyR12uL/ot+dN0R/ByIkDzYIYto
Yf8FF/E3aJor2cMAAnH/gWo8p4G9KWDEQ3y89rmFo0xI9EMUYDQJYdUgG00pwSfi
AFqdUf0gGEaKKpygP+UzMG1SYG5GCTaG4NS87fH1R59WBQuLCzMDTJoHArQd4QMR
MemfARQoQM1IFfzLbaqKn0A/pCX1CxFENOl0natK9F3fdBbwn5TTsHprywWUPYeC
rWykxQoazGp13ykPQf3+jaWiNiVGfkENHLWYDUPof0ik7WH9jiit7NytlFH3+ZEP
H+LLIU/MMkHyj93AFFVw1/xxyxuZGcg6eW6jxSj4hTnhaMiZmrZy9L3cN/0g9V/z
s5QCQj7pY5e5Bi7epxplTUWyewSFApImQxFuAu/MYdCJ1+9BV0cwv+s+zQKRstzn
5J9ZY27BP1m1hQQM7pBDn9W4AlNiWdJbOaNYupnQbBvFqxYpx3tl3ogTJfabPKWr
PuFfa4BungakNBxZDFAybIX7gKO2kTG9i/sPmRT7sKE1XPJ6ZCcOXvqO5Kyq1Mqv
oBXlHIBgRMQ3Jb9bpysk9wHYvv+N4o+9xNLK/JNRKnlPMEv80DklwDOKxrYjv3Dj
NHyXLo/bSm2gurmP9Iew+40H7pvhIiBDW4kXdLuuD3lG9K0xTTPQvhMrhaXvaiFc
HbdV+IGzL1XhBvzYdHQJ4466j/pZpwOyhwxQY4riqRU+EA8F8jdPU9CS+w4BE9vI
NIPrQoyc9vpFfq3Av5TKMPnnKJgQGC3+ehLb8owc/SUSpeLaZfrRkwU4f/RGEzS0
4vChwN1129+lWfTfan6LXmMdiryGDPyj59uhnvQqMo+eY/0C2vOxi9JnLHoK8fYB
wsqEWoTYheid3AaWTmaKK8J9Mutxx464/Ozr+4EnpaI6q27CbI6lPhT8Q7ncAs2M
A8Eo40A8MCdRETo+JJ14CrUWqwjNt7WPLTBhczpheZccZ9CId3peqn49bWosMfFG
B+5ozoRp2R8WsNB752kRVnWnedXlrx5IfdP5O8C2eJCWLPJdK7crMvxRTqS7kvSN
eadHuGb4Mx3wsqHdktOGW+HEBqQ7GjneHDCcUdWP39XCM5A+dvVZKaea/fUeg26u
j9niWUWhm2Nu++DptyULS3PAfHNAfRUJuG2gb229gVAYU8LfE6SckaX72RlEgMPz
X+e1Geme6FGC43SxK7eUh+19AWyf6cMvqtWDzP+f1N8msdQNN7PNgtT5gmqRV3FQ
O40wN6V27yoNFroBkx6NCmSD8SN23C9QAA+noxCfRBzvBq0eq8RQA2Vqf1LLlryX
qe5RKgYIRE16ekClyaR/jfAXjmXeECRf2YnQ/AnMB8NcQRQWmPmgJqHRc9f2dCwh
5Z1ljDXjxaHgQXULw2qaG19VA5VLHXpNb1okG//G1UVPFroqnuIWYMB06IcYFyOE
zAdEAt7GgvUx6E1qnbvq0ZpaOE1S7GQgDEl/70GhlxfdKiPGHiGKvQ9UMIbWcFWl
vMjn8d1dn2wwyBTnCRGadiUliomxzLny9b1EwB14LbXgBely3aXXGCDRTRHyZ719
7gL81z10IHcDFfHsf1ZhYP243pZ99zSd/0dAgQe0kZGuSK92CgAaDWFrGpTl/UoE
xoMV63aZE+Z4E13MdUe6672EcOWCoN3Eq1x0oMRysFf9qLp+PeTWbfwZGJDB1+nu
1Eu+yUCdEHCqvVaoSDDq2JZTje7glnKjCysRg6yf4GW/OGn4YyOpcC4ItXR8ug9j
mG2bSYIdz4GQwqw0OcuLU0RetBddxPPwSsvhlv5/HAA0bnSe0Q2BEaouidNqQiQc
W9zQ8kSiHJVel+eaZDAEehbUeBE3SKaKDIZf04R3oY0HeI1avH0jNZkKfHQRqAoX
qphtrA+T33cKyBozWNB0tZ1BuBC6AH16AS67ODYqNs1NV2apv4wKuo23rNEZ346V
WUbELvoiymgheOjM1xpdjN9mfGprlq6vu9wNn+xKKUJx55tkgZute4CLR998sN8B
oMq3qNn9u+0Deh4fpYVOUFMtE25xhKoFSDqgNKStpX0lIt/DsKeer4+BRPB0dV1K
JdZGgSuFTDv+sOkIqsPt9eO99Hsm8uhKh5mbNRgC7TJ2s7Oz1UJ9NLfgjLmn8V+w
PD8abghxnd6Sfetl2EP/piVm+CdSPbuljCUANDQSR9qBn1oIQhjdD3XquYtPwylf
Cc5eG1WP4wm9GvkN8AXBMIPFeyI5nCzKHHI3wK1arp2iN7zBAmHzUnZSThbaTSVP
79Uayh4RkiU6rjx9pyE5zqBTI/cStMXurGMun+quL0kDVaUWutkHsDL4q4EYwdjs
73QYqUj7WRZ7JNMJcs5rK9rdn331tEy5fOOwQC5TBlfx6LJetOVRo2X8dMU0AOPc
rSnU/Gceweab4isFCv2NtaiUaqcKTQiLiU3FGimFci7cixUWm9A0JEk6xt+6V64o
1lxCaPn53j2n2OZeuG75iHxV16j4tm+YOPS5I3PlI6ldODm2fVCoFC79p1smJSYs
Tf1hvDF6PoPc7fEvHB3494xMMIMKMqA4qAup9CizJqVH94b9rfps/5sxrLK58g9k
C8N9jQH4eZCT1gD1Fk+YgmBWtZi7stOR/W9stjK1Zt/S9NKS0Po3NT27fzol5rX6
vVEWk/gN9hyVgREExTpgNHqESFXxKsShk5WUr4gMzsgJBYxXGN/Op/sIzGDhtMgV
7Zj4ngP8E7H36ycbukPkbB8zhUuPPnL3GfbIK1nyTliyVtYsXF30D21Xpa3eQlx4
pYf9qe6o3qDzHL/VH/bakWMEQeV1x55xCKZBgN0hFSagrKphkgquDos9pLmWNmul
JUkZeYh9/zFeGsJ24ltOFyXAro7p/8/y7QJQnlcdkCDNK/s1AS6hc5hGmy+Sv6ws
P/Mei1s4K+ytsOlx79sOmqimsC4+LnONb9TP1RFnz4Qsxnb7O6lGUiAUVRSwILia
mh/R6jx8g4Vrsq6rOdvpvDIdIFwoVuZ9BwDq+uJzwJeRUmCQX1PIxHGoaetDNTPU
vsOAjfk4QyAb0A97eAB83tahin8sVi9KPZh/DXzsSNe3kMp56iWucFKO6/T98z5c
QRQ2Zzb4LiAOjIbtAmFhQdzO6I5Ofz9E4a9EKoXJvxMqhPj0NC5b3c4FVTZKlvrI
Gm4i7Sspfva7c6ddIYceICh1Qn4hGMrLgrSHZZLGhpAXxtkyzEgF69NvzgqC5OFA
Y8Q0DY308wPBkDChN0tMK2HNoEzOJYcKEefCL4TQns1zxMwQCtBJ0+xPrAb1VUcB
FfUfEOFbgoEITz2Detd7/oLKAy8uz21KjQ9GYaPY0GZTmWu8m8Ow6q9o0e0yKyh4
MG9AoZMo8djNOLQ/iFeT4mAb9rpZsxIaF4C9F1DHtBwFZaMRj2XklWRc1hS21TES
1If5SqwETH9M4eHBuB1x2eWqnxgqnxaChBSoPc/8ckzxxPtFZ/7iMDF0IGofBXEg
C6oAhOgyosIx3XvUp37ulfBDfga2OYij5CpAkVUjLjWlumsd7JGM7YB6b9faInuS
bWXbcTdB7SDcLvQFB6bzi+4g7Oa8fPJt+wA4nk6vqy/kTPtF/id95lgMEZ+NoGUk
0N62z2PlYJHHABfit5Nv9Amv0fhzri+/KngpO2ri/VWvpPngeuVZd4zoDdB9RlCl
WbaPQTSC2kpj/aE0BrndG4Az35rzSemPKn/Y86GYO1GfT1Jv+wXBBK6V6BdWEUtV
4VzoD3uuRjhoU3KOX3Wj0nyQbHvdqtf4kwrtcwkCp7FTUc71/puSvcUfGzOwx1Oz
nf1AiG+1w0v3i7TbPDXItZTsJheC8F4ahXWLXHLYoUcQDOsJUjNPiMkkO+Sw8uVI
pV/AiNLYr6RuB3YjGmoQM8DYxSaGHcuAaPxh8vFyvTdgp+gCuWCms4AEvVfN/rXb
LbCaevdqqUV1EV/GR9dW1pQL9q5dp0LvCbUm1yd6C/fxBFr2V4oj9oMUjK5hin64
28pyIC+GHSHzM0TqUGwbmEOTl4Dowrdr8czzIIRfccRSnwOqph0rOy8gbFMQis9j
ucuMpfl+Z9gXZjkhOAeUpx4DijKkZbmlQLaz/OzUNe4Hle29M8rzS0u2a62wyCCI
xUrZj5WBjp3bDlkd+OTRDfnsmH5iJSgfyEn27W8POvN0RRgeM+fT0yGaMmCVGTrb
QN/iFljFnKQgtSWqIyJkLEh3ywamk3LjM0z7mBrwjkm1K8M/nPVeu/++N8zYCHTn
MGqVA4S/FPZNL1q9yp2HDbmA/vxzDYr7Fu/WnjbhOVKkH0/kB2W0pdL2xG0UCTvb
EM7AZ8Xv3GdrONM6UkttK6ZpvDPk43vo2KfMQx6lgqYpWUPt4tWgUmpxPMp7I1IA
PFQT6EAy03W3COtJNgO0fvQKvq7XcqRbZT3IcB/u+PIWSQJxXc4Xiof6z2bKqyYm
X6XaRWDQvgmwjFllwv1aKOtCXqajuflb6UWuE/J0NTk2UrxuHxPUHeEPRTUtq/q8
FpIGQPadkVIOsFNsdITsbSwvv+XY3QGUOk8wrD66bxrhcNTQqtUE7PL9Hz6+ezpg
6VGnA3yVJRowwRpzc+4cbpigZB8J71rknNfvgwf0t3TXZeVZzXxi1WSRw8+8o0xd
mV24YroqqeBzLZUbd83PNDgCmA2BFkMWfqrEgL91ERllNTAmiNqGWNyfjtBHR4mP
H5u+Wbt/vgJcrTuEnkaG1yFxLd7KqQSz5HFoeasvz6JHPbs2GjZwB5u3VUFFE/46
SJT+QqAFWsLW8rtDnuHh2Aajo6gZyQETzhZH0D6LD9h3Jtwob4NrnTLiwYtDwAGD
bO92gdSbbxIDadZ44ZYvQepr+4m6Kt8CP5/Ra8g+aCRBtDqMJauJcLg+BJLF1bgW
3vv5Cg3iMw+dVgUUjBHt5D/ngImPwBB+i7CUzQFtG5h1U6umnA6C/Svnkon6b9V8
/KwjiEF3Fgj7A6/TxKLQiZoQMKrwMkGTfTB7im4V1iADsG3iNNKYLJRC7LrxruZI
Fc9xaCqGFYEs8qKu3FzVwRI38YHPU7GOC2rTYN9bYBojyHo7AtogfJtYON3BPWGk
uWw7U540cuQsTzX0aY5Kk880HlaKqBGJNMO69QU71STA55huzAL0s79rnbfPko7Z
DWjgZl8Nsy8C2Bp0PAHouf10DLXpSP3FDtjEzwNDWrDuD0O0UOAtz4X5S5XzNUsm
4zbQN0NlwQ3HPhRlSvGEw9IakmT7ok909kUtzQloNKnpljzEGht6fGTBRVx2Rhx5
MSmwe2plAE2Gle2uTpS8AvjSNb5W3CnG4tBOmDfVoR2TxSb/QZuPchv9KmS2yTWk
zSAjGbHEBp3JZf0qdOSjH5Upf4GJhoYA2c6qpcIrBhq8jS9kLE6Ts9nuWCP+XU4y
u6HDOV3VSZr8njH8/1PPdc37UJeCUqCwVI1e2ZmPB4PslWezws8FwY9+iD6bMPoA
YkHQhNKAUx7lKkUTQ5t36/7CVWx1myTd4Q0nDTc4msV4UWubAqdyKM55fuqxevbD
/AkWPwj7JtuCre9e61759G/zIITrSR74iOhCC8MhfnR6+NtnbBRR4WccyjJ3KT4a
H/+ZRyIgh1ISuYWxw8IUlvITKwtvckrJGeGdd+u2lRu09Yhk4Ow317MEvRT/Xj2I
SJTFqUX1TMMg+M0WbYi75PtkwcuRmS+q8S5vQiGliUJB8hOKud7tgWnx7XlAhv21
bL3YDGEvOp76oR58PRZ+qc6Z/1a0Q6HJTBBS/DfQy0dXUNiZTyl5F+fw5Ch0BDcf
as+L7uH9Fq59hAQsFfs4m+8ahDzNxhTnJHyS1Qb/oHXx49JwgscWKIcm9lSY37tj
7GOJGnUe9XGT8jMgrhZlS0gMDEoEoqe9pVYFshmA7FW7tifykM1ttEjuH604FAOr
s8DYBes6t0CNhrdTjQz9AD62d6fyKLK2PyUaPb06xYskoub54HxHcOu5xG3QksE4
TTiEYdd9o3GW2oNDMGgaz7oLO4A5VQd3RKS5QdPz1/N1mVJ6ErNWGD7OYVL13b1d
sUo14CPG+ipAqTGp25dZBghVz0evTYHyc0bBknm0XlOXxBLCntsyBYbm71v0gc85
Mhm1nAuHWKX9nPmZ8vaowBgx34AL2G99PQKCqrbBY82/bywJljM0nuJaxRsP5lee
TGa9gse2B16PaYGM1bOzh8IoE+E4GPS1CZdFHHabuhuoOeI3ZqAAbwsjO0dOLLyq
OyBAmR8Z+0lkgmJOh01IVPiazm238jCmvK1lQSRIt3mPQuBIX6F6dRkE3QCNXjJk
7UmXMSXKaWUDIEeOehu5kj63oXkyYwENzZhKhkQKMhj7ug0hIV7cTYXTeEJu2S3c
lRSLT7wt6y0jlRZypd9rjX12gylWcxDdcXIIjIil4VA//XaumNPEGnrx093hNqfv
JUSlU7Q86nEQEveicAVYV6RE1v97ksWCICKdn1DlUFPx9DqbPTPQk48B3BhkCf9Z
Q7iY07VmNtAC4prvwELnmxwAsvI23mR0Ua16Z1JsNv3BZhhOMeCDUzRgJqaMHk0D
DLOIjXdRHIGmdFRwVRz/y0INI7u3U7q/FtQg1S6XwiTDQ/hi5MbEJp28dymRL3qx
3o5umQfd43Tgz48ePy9AE3gB4EDI3KDUoAa9zo1bEDHF2/qAgMpCZjlLr1VMBul5
Z9gRiSde77O5N+BtfumQCt3Rf4UbcpeTWwBfhn4LbWvSYoVzknJEUKzlvd7PKZWF
3+l8SV2tckD9cjjh3fISUY2VKnSifnQ4MxsmD4+n9o6J0H5odTdouKcT+R8+IUA7
wkrHQ2BCm6Ke0X3BKlAFCm3l9ruoTTN7oN8n15skz7Lv6/YD2sSWPqCUbE1gwfCP
isddT5z+m8Er1ALpz8AVI5Sy5FaF+WTsxCw1XfSzvg54Kdl7eWNtTWHCbOH35bBY
nNhbWGS4Xj1msrs6ZCrpp55k+Cl+HHf/6eJbWBMc/qURv5J5UdKWxqBHMxo34pmN
nuVbwvI72WBpoccOMYL043t+xwkq4sXQeBRdFgrWjstsriMMYW+q38aoqKdtlP13
VCHINVAHbzhTMsMBtsXW2X7fAMX+3rt0D60tLO5Xeskdeo4kNLtLqWJh2aIDrCOU
7DRQozkD2OAacjROkUzv0BKWK0wbwDlUX793jInrG1u9H/33QSp/T10Xbnwk8BiV
7Lz/hUUo4bDfi0ML3v/ud7bHtzxCnUwwDyXpk/n5J8iVuh67u94hcX2kz6TRK8du
LhhZinvpKY0Jrr7eKK5n3dNYvjFWPzSUIUo8Zr0XTsAFsmDlvgCCH31PNBygPZjG
0erLdi98XZUwC5Vedgr6yhWSdTU+2yMtDctaLlTduMmwMZbbAw/ioReD7mYlssGj
FmxoD841rSard3X5DHu6kiLtn3viCATuYKQfmJa2pfEDrij55VvGBp9IrLPPgRrO
HBF6bcWcQg/GxgiPfnjjQ8tNUPtgPjrOwMvEf0m+vyi5JdLyS/KSnFgJsyp8bNu7
yx8GomuAHJdXjBFwVSO0nmwYyEM9a5leyoBqp6l8YQssd06CSfQgq5pAm6DtG5P8
0zodqqzSUjA2oL2R0sBmUSAdeJeSoKzNo9JvmD+ABShk2X7m4lia9muTG81NKdba
k9CtNvLqDksRFPOurmyUv1xa8vcJg6iuy2iUI+akdggS+VDV9JipFnEtao8tV4KC
kmwKxMOzVMogX2chx/s/pA7DAFq3aEYCRdHld7MJ1S8phK32bu5Mu3vzqB9dBoQR
0erjUIrQGTnrCLR7f9k4BRMRQxBHOh45xmFZRvI9+dxJBUNco6JGrDbQSiC/U2KM
NsaPgRWJCL7wxE3zWnKnBqmMsHMxsS5xxveUdPV9nR++bJLclONYvs7xTbFJZUk+
W2DRVsiDlSvoye5wIAbWRRgR8XiMIWFSWM7QxLo91wlPTtmSd67u52XjtDQ6eSaH
SGAj7R4OnUs3oCou/gUwlDlSDW8CvBdRgX0WXZ62xAZY8JwdpM9U8h+vuY8Gpv7c
yHpEqPtHUNB+ZqV/4oFAFOxfmOCZVg1DmqsNAMAWTL0Tf38mBAr5ofrPYbtf/LJO
G9bdTRsU3s2N4yo+qFhiA065QpHnP7fkcX5ETvudQMdYGgI0GNDDFlQjqdZTn+DS
n8SYTypXEfF6s2oxTNzpCfo32utmfNqP2zYR+JLo7BRft8YIOCo+QQ/Zcat3Avpk
lR4fXnaIEUvo9OOn8VsmAHQquKBx5xdxqaBpnTjAHHrBLWxgeiZb93Bm6vvWdJCy
Rx7npwrvB9GbpOnav19aTaGfZEYmGC+JZR4JUwLmLQ+rC5h7QUf1NBIp/ZVf9FlQ
lVTOCIhYs/XFeJ35hILPcGJPZB+VpTRJjIvZ7qmC6JJ3BzRQXZBdgWJWNt0rdzD0
BnMzJMs47oA5gcKxYgzrpkogNY6sQxPJmZLVXTDDrOZ80mDh0+JQGohHqdyqwLnI
RKHorKWxqQQnPiWNmo+0GtbRCj5jgstt/68DgiPy5CwcG5JdZ92kr8rX2Rar/i/5
1JrmXiCpl6FT8QJLI2kqxs3l1kaB+o3hhI1PWZkseNwmNnIRpV8SnsM1r7O0pf4/
VGmS8gK5QZ4yGZQ9LAXIg4/uUm+fw4Na1gpwMTmGYUvq/aoCTLzVhplYxf1FjzaS
mh8hWjV+hWd0gYBpGvipUXjKagl3pTY2gVXHq/5Huh1+V6Zd+14rj/m6uqs/8lHX
QImoQd8iMWUzOm58TSC4W8Uysdi7eYG6c5uem/GzRJnlQRw8XIgPM/Ovk3JJxDvi
pmGZLGAinoP6GayVEHQnNGZ4zglGWcD30oQ+1LdRxlI9nlkmtptL1K6iZ3H8jX1d
wgVZXD9gquUpO2Q2kdOKOxcnbUmFPCFPELJVYT1TqtDZ7bHMWFRP1dCcME182uCM
BevjEA6LrOQt3H6MuWPZTQ8jooVDAMi1FYNBG6allbCOSucyMR+GObZuHuav6Ufg
Y44kjiQcM5gIdZ8E8AnWrHcUyWzllPfnixJJ/fvGDM7bmh+Tcq2TPoaZ3zYOdlJ6
ybTkAahU0iIasOVrXUDj0znEWY2d/EJ0j1ZPdx5KuBSFEJ+eLsxkd1rkBqHq0UhL
+Uo449F8GczrcnuogPaP88yYM7yNCyQNefZuvv/SUTSopyQBs/0D9q4324CuQCpk
39tYrn9vrsTWfAb60GFkvqHUgwHnxQCsZmQ3qmGfY5R+k0Xf9ty2zToykjXLF2Eu
AfG10lbxyCa6TD4ckxuMxoOKEhJru8lSDi/d2ov6Qht4OvHEUU2AJQuCRjZmpkIX
+bsKgS/HpVd2SiWzHFF36iagpB+rFI1XxPjoRiIc0woJ0MXANnzWa/sgOVNk+Ssa
QQ4zyGm3HyBUHQr68hKCVXnjFTtFtnziWCy1wLLnjvqxvvJ6mLwR0BWBK5uRbkoq
wiyqpvC2YGriQ28hQZucygBWUaVXZ1VUE7+9DGoRF4InG1L3z5OwDOP+A/bKbQ6x
oZzHmrLMWztLs2fW01JXdMz4I81A5Spuvbs0m3DeiHyt5rcUVN/Sl92BYcQG9BPv
TkI8rdbpaKZqbAtFPFyGycnuwuY0BFNkARvaFZDEnsq4TyHFqW59hW0wFZMrrad9
xCPqKbtdOG3pGPTjUyzTZSnI/7g3APbs6hQfeKhYWiG6K4QjjgVISlgttRyoG7Yj
kar2wvYVT78yUNM1yziVXQTnkyFUq+L6frMS+EqnnejV6ibO33k6+nr5NSewCG/W
Bqznubd76xe2C6BPE7cNmJ3UuxzVtcU5HWPFAZ8jXWnetQrP+TE8dle/jTEu4o3+
b9bd84E3TAi/u88xfIxZ4plHRT4n0nMTaA5p2VagE5oBgcKgii5Z4SzTS1e/Pn03
jX8RpYc52MqfuCtUjBzUrppyE0eZ4fNhY4WmAujdgt+mTZDAtoJMR33zTCMAIUGy
2J/JdmyIn9XJnHd9x2pB6ayxxaU07bjCXKBj/le3xp95BJL/C9C4RAdehQbsiJ5z
jwsn3VKjwPonTqyjo3ifM/fSjvuWTue2Dmrg9U8ZY6Bt7jpUbEGrBpl3m/1ohsDA
9EscVSlPosmIeOmWsH3uy8QP+7VYsbF7GHTBOTB+xXTI8mNn6dIDLf0/55j8hZQE
K1jLnZlwaf0QD8va3u0T4WO+oHHlnEY1Vn3ZjgrNnUXW25k85+4md/u8s2Hh9kMt
dxiDQBTs6axG8oq6ewhASYiGATrbW+qiCHBVzfqX/X5urQBjfcf3DaTldyp7/fSw
k3p3Ssrb9m/5v+IyjoFUcjnXI3O7WVu/icFw8hr1J5i8TOuBrOCPKBXwxfaErose
2ZUmIVu9IEq/dp42pk2l3sgidAGTV9eafQ0t3p9CeuEIhqd2BtCdJWaT+wNaBVTr
5qKoX1WAzyJVIut5ozbaTSO7FjK//cN07cdkw2aLUwar+ITh2oME7U1gFOsmp6vx
OEHbJDnIzbJezHBt1NGh5aCKVteo0KjWpIGn90ea3nlgBg18Bx2NSBzlF2KMJ4j2
aCDSDuSf/0S3oR0Y0BE5KHMs6jbt1URZI+bxlWAk7pZBrdl6324pZKMbPV+ECqND
F6isQPDpBtCWHFjF+ZJXcIsPEkKZIQPhwAFrgFGHbhIQdBmqH+w7pAM/gpOVF85V
DICR2C0b9Ib9GP3XO0k1I9vk3eiwAyaL6sGN7Hc4wH47emankaHSUyOVkYTxpmQr
OBWXjJVykyb5758hjQjkT42myYdtt0+WLLL7HzxFKrlHh7yPV31z2npRPLtfyCTG
iiT7OABidk+pzn6S09hbZToxNIsoqEHixY2ktl0kqTwDyUjA3TWA8bCUoG4UI2Tm
pMd9Em7/5teZsdjEkr8MzQvD4m0ZcXQubJAQJYmF6Ld+syOb3K89FTFpcRwHYH5M
HKLMpdWfoWPYDk4UIhNJ8Ct8HZIp1oOscuNNxxxkq3Bi0bNCO+fZt2aEaHhKpXpH
3zO31vdML9qd/mE5N07LwLIjwi/2D1OoO2oXpX7iGV6LTidi7FqQhJffjdkkyJkb
QTIlUvslLmMCzNzFGsh2m99iRjC2kz21siM7QFgeWJsU/2emfaDI799VWFeoO3vJ
qea5afPrZ+G9DUTzVWNW0x65u99coVd+kPeLjdgiOcXGmG2yQJgZGPXGyiaDD6ss
alwTN/kPVbRn4DEuYupdHiLOAUD3yIcjFWjfChIQioYYoQCU6InZyLkLNJJ3g/eX
8ep0HEQcL1/PWKUCQwpBXZlsx7NliHNCZX1u6LsgeuDF87ijUYi7KTQ6joqCnLzN
5dCBO6CHk7GymrqYIliZ0XEaRAfwcDZnK4VcB2x7tUZwTZFOxSLpAXSFgqftDOaj
FnBdgVRwrKD2B48kOIG7yjSaUAMWTibIxpiuItx5UA6G8N0T6vqq2dlHy5iFA0Bk
CadHhJ+Ou677Zb0bTa7hFj5NWrlLNsecdkQR4Nx4KPwkonWE4f799kEG20WEauLG
pARam88tb7s02WINPQ/dhE7yw6GnBN+2E/l1CAzTdpP09cnsYW9LZfxo94ciQGI1
d6+Awfw4+HUd6Yfd5uroEuFJ6bIBCr58R0JgkqayT97PYKYBCmfFyHgqOr+nCKe2
OjGhYSxuypMdVlFp4gHoAxfSbbI0xCreh2cW9D3wpusgThnCKpdfud3a6mzcV3Ul
FY9rz2A4oO8VfPRIhFSKKDWhBGZLroh1oRB8NAh1Gxeygx6DmW9DcJy0vD8Uk5XJ
uupA42M94ABMBT0IDFPGiKeQJ77pKoA4yDRmQaac3JXGbYrOHSRJ/dhknP4UFHlR
uW5EDes59UNudFswQFC0n/t0imUDG4QtssmXY70iZbGEj56rpen9rOy7IPYhUtCr
3Y5ayyvbAZ7MU80t/N4RfJ49+rSebcOXVPfFCbIWunTQv5WzV45kLrNTi6Y/i4Qx
HpfVinX79XuJPiGqwEevKw6N8OS1ioMEwy1484GUd9dIP5Oq+pCPhEuZn2Twa70I
RntNZsr9dF86gCCUivfCF7zVR7wM4FcFHyAY9vMeLrfflSJ7xBXs6LIpCEFpO7O+
yrLnC7zX6XYEAnWL7qccionNZi/TdyXdFT0oukWIQdIAWypN3EIFQBtNkW1rgu8W
jQhUhkdFEQVeSLNZrN2cDjiKb5lQB9r7i9oesl2t1FSuL1Kjbp963aCNIzqfkN6u
vVuldTzB+u2tbqxLHatHUk5L02wCBw2gucVY3lDh8abbto0MMuTXY8UC1hvt41R9
8U5kaSdHkAeJ+ThzpdJCMvAfu3CvkCzj1jaJEz2RTq4EAl9khl2jZHEsZsxCozM0
7HAMsDrozrO00leB74tBGpRNOU2GZ7k5VnjinGE9DBekq5my59xlgfDz62TeYSeo
kYa8T3b5TUZlTInBwlSeLMPUjGtzW1l6aHMFhgm/UVXdMbXQmVyHA2gjo3r3S09f
6ZxVBmsV0oIeQNXRaLLmQ1/4dGwu2t+vpXz2sBrgVEdU6UcPh/qAEE/+brTIy1vL
Nhkm/mQ2FduE5vdLpxIE0g0ejinklg8yVIdjTYiIRip8w4TlZ3FhjL6PYKuXdMD6
GQPVtTR6uFHPWEJ8EOt5jBlA687O9lvfKykc1Bn5pmO22tJY5NsvIifKomp3F2kp
JDmb+TqzoPXbt9ZsXooIP94XeTUX2dVk8Ze+HGaE+tlwYeKWeOaDvrnFE/2lrxK+
9PC7bJVe2ZcQK7J31nb032EAMhD22nXzP/nD8U+tlaxw34+4dr8YdxMXDcrWBMBb
xuZ7BGP7jOMPbszkR/65/3gLKxEoWSWcP89+kMCZzf0Mxmu7n7065+WrDQs4OpMv
HCYzFg6jvV1/ophfm6EOYU6LSY3hvSPIw+tkzf5d3F1tVQQYDiW4QkW7nENYCzhF
PR3Gj+YU3F0eauWJFu/Q+9LJZfh76B08AyfEzaLyK+rEwPqqPV4Wt+FKX6jq7yxS
MM/0CvUdTr7HUx0nMyd8+ZplFbw0O81OmqqZABG4QpQgwBFOfnXhysolv9qHv/U3
vtcr7MlyHNGJQ5EEtCWN4cb0F3qwJS4A337VgYE8lfHEmLJaUwvvxtqYISUTm7jK
iL3nCB43icNbJE2dWYyvKs1yekcw3wn2unLghBDQqrywNclcfoUe++wbKXSvkIvG
YggWra+1I1cEGsguUSb0jVpDB/+4tnYEkYIseAn+zk1/2QwKnjECsbQWPhViVtGR
lliZMEK2cwl8u1rRkliUdWhD1qDqNOQ0yWAlcliw4CjDQEuURHDj13BGBl5i+xag
Q0ws4djYK6ox/E6/ymw6gjuDNb4AOB2Q+xzvMMHzcXsLdh3RRrYqgjy0OnVguNM3
sbNqZNv2/TGmLEdPriKm9SnURQiZEixNyPhGheYOFPGZ/m1Th5MOVxSdJh2lpHtV
u2hgRDc1HVzNx+36UlS1gfErhkvJH3CyXLfgtl34odI+vnFBUMIL77wj5OER4Dbr
9F7wB9ouopfFF5UmNaSFczNBfURx/GET5VTYSlUwGZtkCzM7y6VjbPdbBbenqdon
pCYw44TLwWTw76RVU9SRJXYwK2/kCOjN1MxbRFcJXPifR2GRPqz+1tUHJgOhEJJa
UKBnwKAZqyjTGw7c6y9VCUaqMXhwmwDKa6bOsRKQO4W09dSzPu6MZ+kQO3R/IQz4
nlRBbirvB3NX5VndpcgwMGQQLtzQ2CudVuPfvFsyfGK92jbGj0uJKri8h4JopHg9
EEdLj9wV7zFRBf1MlvHzO2OF+IDZnA4EK3G20+RWuQ+UwCps7ECndcvotCUJuRZf
BpDTFb5QVGjfGG3ChjbD806PNO647opMCcGY4KIMlYQgS8oGhAGdmJltlzvFfAUQ
9WYaoUK1/hvF291FMi+NsWIc5bN6+EQ7pqFEDjqOCeIt15y5I+zl4bYyQ837OIAd
/CsnKDFZ6/MgmADkzp9pxExhm5v5hD7zXaOGazayR6TfLrQopjIe2tqu3+Mq3ItT
FxMMgB8Ay6k7q1/tGSF06TIW4cFq0N/c8zFd3S8lHvnDTCAilr6OF3aCLYYBnca5
R0f9ad7ZA5ttxDsCnT3pCDEl+P6FEBydLrolf/1XDr2AYF1bofdALh5j1wr56FEw
zOVU9IdVwxHDiDEcgsnzu2yvzWvpabLDGjRg6d+M7ZDU5sVs519RZ7J2cjazhcAp
fwZNXGi1kAD4BcYaGwoazdeGf99L/SwLjff2JnxP2TEeo2rSB3YETxFdL/pPlMDk
OiDtMPZGgFK04KjP7vglrZrLbKfNQWVfGdo54VJ3iJFilGiSnrx3SmXF/BRCn3mC
pXngN88C46Vohsvnzxtw1s0lWYRboOhLAyoQaR4moEqFMePvMTsGJXtuegjrXLU6
xrQXAeEet6YSA42WDJ7A4gV8eZ0Qh+q7J/68eh8vc9XZiB8HMVZ/crRL2nuCPc1y
xwSVKZo0ZsvRZ1FW8AcME1XacSPlXX4IS8BOpu/OP7rwxAKHb/EaEt4DkjhPgkXq
yd40YBYtFNpkOdywPv9iC4twUeZNXa2IqNXvIj1tUrGzTJPxNMFZsNgYcfmf/2Ba
C6aUgtA2v5fpHpRgW3BpzpNHwg+bwXm+xxGmzm4WqRCuaUil2+Db71mCrSc2JUyT
VwXomtShcQW+4nfDT6+ZB3WK0Y/wY57Xn5C9X7+z+LK8/nA1Z2hQXesiyyAd1Rg7
QTKOna5Yv3wAZNOCS0Zu3roOjbTt0aJ+gW4DWEqEfyDtFXag81UNDKBLSl+hTWLQ
YuBnwfFC6qzpKw2yq8wOUyQun9NFnN7722FhYPejwhy38ELF+K4Rct/MKWPxUovH
BY80DwcFPLOV6zGskGSr9PW08rcikv+bk+M9F6yT8z+ww2Hs1SJJ4R66jFkEVfId
cqvylXgRwPk0Q63XnR4kJqfVIQITVVSMwr9DYGUBhBGF+u/ADeUtxbgMc1ukkVXR
yAP9d36ciONldnfUYojC+xyLODnAxNJ0YmYdZjlqebM2C57+Lb880kYIRnFaiBFO
HKscz+RXmTQzGAbdgPgRFi0kIAk0c67kka9fFIy2IbhzLH7IPJPcmsxLnQTuNgH5
6dXwry6n8Q1rQcvsSGFYocAUJE015KefXRVIMAsJEgkeuD4c28vASEnKrPfM+t1I
52FaM64BSyKwXBWjhfxJu1DjUxbu/ODD05m7wvFs7LnwZjqGhdDxYmZQebpVCt3u
rcgk+4ZeigXbs/vx1fsI3+yl/4V/wAmlJmUa6YC3pOVPU9fSC/WyU9EutFFeQ3of
Qx88920vdCXrMxToC662j5vJt5sZvGmKgI/g6wpAm+h94Za6ViDBW3vROXT8ySK6
b90jdJ6YwB99PNrx86x9dD3rhl6pjo1qmprB6tLRLxa91nNhkq/viF9HYieJK0E3
zoXeKL1ZAwl81FXw4XSE1UZzLiRgY/dCOgwY+rqba0LRBMK4yedwRBBm7s5lo/DM
bfP7I/aB56dyXtfQAweSF7L8QACEMXMG378nHskRSFcXFtxoB8vckQ8XvBMUzHPx
4D+MfUqEY8SB3OBeV9mdHP4zWENv1pEHEBP2nNwFj84I9qD3yeLcyZTUArR7bs3/
PFVR+2ECCZcu1IalFBB7mJC9lvC057FSmCvNaph6DPqHfXY2UkKbuNIxm10pnM3a
3yIOVukOiAWBprp2Zz/X/NPmeEKrCcUX1P85EDJITP+ng6/tNiVfdOrCA9JvyJmx
mM9x/vY6XktdFU9BQsQLK5jlUkvtyTSLAA85+GYC8deJ44OQg5Frpp8pz93Q7JF7
q0PuJFlvWTTdjb6iEKVE8gMAzJdWgE/B2uwwKLg75/tmdOW7Us6QWCs7hEEgMgmQ
GEvDkr4npy/9DLgI8jueHOr4JJ8MOYHHtF5xHnF2T4miE2N1OV3SNBqB4XBWOhBO
/Zpf0Nh8x4qDW/8FLjgFLdsZeYf7+qyTNaBim7LGUNrUmgOzaVxRAtoSw3BwcvXz
Wu6KF1L+jhp2mJuXXfuy6d63KwUHS8tUeNSM+NOEil0kHblFCKHFBDsTaCehAucp
EiU45AWJ5Bo15KAdgywM3PzbbjnZRsJ7aCB/hLrVMBDQETHCGVULMyUVyMkzjkKy
9g53RfQo2dFKxPgxbRsVPgTAhL2KwtBVTI0Y3TmO843ixvaB/no2s1oVZdONZRzo
sSzF8QrB40PuH+ngG/QBm1lbQcdvneqFfdoxOerBpyqQuj5cT0uMhmL0bAKW/GPm
y375zo8g8GNxZcwP8B4Xw4aG7KWxtNLbpPx7HSl8/tWI/55o7DT/Cncgsll9oB+9
dcoepyatncDCFKNeJmtj52mHfsqi0MYVisCrx6CKYp7ob3j+JtFDGMUFSUVJcs8J
WtxpCs7Jk/1CvyhoO1j6jVUrjKMB+rYFPSAur/H/g6WuFy+dFV5LMrLz5beXjewv
/qUQrMQmGeP9/CE2nanj8HdugIeJclcd1YTiFiqR6rdwf+4lN9gZEVNCwt9/BeqW
7kHJ9W+Wl1fGuZAaOAtNFIiAsdZ8LLvZhn9xu2PPr7AgpGaKbBvjyKZdLg/CYfkD
RM5jBCYQcpOOkISQjLdCjjrEaVyxdNPfafF/9BTwKPl60936clUOIAMmrVrH1JWt
kt+N2lRjC78HBs94dPRMxst+cc5HELaekqELz6hHoNp6KyLkPsYWOTcEkod9UDgH
wuW7WiBTJeHWeihC0scLAp/rTr6get05GCCYS/v2wfQnItqsibVGoSyKC9Xw+SZd
RcwjKGSSK8agUrKDChnw9uWN1LGrUiRCrfE7mUaejg/jUBtx5vcQ70g+qTasVdzh
l4J0bxkwH/tjenD25NAgpovhVuKFOd4W40rkedlX0Uyl5h65DwDHW7vv4RP6MqaP
K2z0rtlQwHILxcrM1LDPNsM2GRr6lILlkCFH3MwgzZLfSna80LUQBt59ugRAfFHb
Uhjrspe7xJMBRxUJ6WLJ+7+03rKorumLaNZQtxIknwzFlXbYiKI9WDS/8/NgRev1
zYYnaQl5VWtsKExUEujm/zRb0LJpuwqg31uwydQZDB4PuEUa3oXw4V2OzsnRIeYc
VvnF4xbQufkRFIt9uchWxeGJ49/FlqzyoYXFSpEzp1pvURfNij3pLRdke//TPOHx
rhq382emDZhY4fkaSfkdDVB1Aku4OKbHnstHKs5ynNQzM4p/+cUuXSmz6mv869u0
SqWuY3GpVs1WC92uJMJ9DMPQ8+Z2OEsJSEjTJ5eslSA02gdWAiP2r8e3EdwC1G0o
nZNBl6MGlN0toXmbYK3TzmPKrfcy5iFv+iSRR3YS3izjVlmCuyfaG/RmqWj647nJ
pOUkHzAZQ7GBKxJIMh1e7Ea4B96j8MPeWhtecHoQtb2a3CtmCnwlwqx45vsM3ssY
IAHFMqj9+8ykJt8SZ6VGcUHKGkbJK3LZTLDTpoBAArI+2vcDSnYfSG350fTm7hPo
wmXNx/s/5qhmrLWNYtPGQRrPmmDmg4hylRoZfq+o0WiVA/glrdk3bUruoODuI0Jq
leVFVWG9hioUh1GzRvkGxWETZjBK55/0gpoB4VUW5ko1w1s3glE/nyQpKHog/wn3
VQxNIohDmA6/I2MNMgBapEziNPLKbaZI069qnR3Ys44oHWWqO3Nfs7FKmd8Prf1H
oHENhWAtSjsWz0/7cQO/Lxo9DvUf1/AHIaE7lem2YiqcY/S7PH75qG5Fiz3IlPhW
PE61pqsNCJ+CKj8ua8SAEWwmlWdWUoT/adqF+qNcCFtlQJHsftDsYqOJFNfB1mrq
zJ3f1dibGHdh4rbsHQ6ZOQLlie8/rsY2B5cSROo+4QGi5JhE7VEMuGaZnC6JWpjc
nN5JjLod+tdnxMIIHGL5APrXKU3lQk8Kd5pCYrrym288vjkTtLC1Zs8t+JiyYyfV
4boe9Gsz3I0uXuiOdkThEIhk4Tu8qwcaqoJCcsz45zwWkVPfoozzgmxg/PhZa9AT
WkKEB0bRPaRY1yjS8mqMr3VcfvRjUSjfGR8Xl+BWQh3MUrN6wVY8dbPuv3ImXzbB
86JjFstbF/jmj3+6IfkZYCbc5m9FPb2NFc7q0imLq0FxWngVB1ukqKK8wyBKBcjw
KccMyMfzuiK+icpBzGejTyu1wLovSQsowtAiHU0N/fAG9HbD5f3TdCVfJ5eTA2Iu
QcjOOPwOsvq++6oDFn+tp0TvC71eKQYcbNqqTr9ZGCIEmDmGlX5jqFtNmU4nSEeA
kKl3NlNzxQ7LmepJL65BMxzA3ggcqVrx7nDGpoPMcqhvGMFJCtn5g7XVgkc0YGZp
qyNFwdetrgB1Ai+Cw6b1gbounmgjmqGmAdHqZ85FGo4QoPMkfU9h8XmJigCWP8IB
yqc3vSEkgIa1ZCWxz7uYtlijElKLfPoaIQWb4El1Ky3K8n7KkOtDU6g1TxWhdeg2
EUPauZzXY+pOdyxr/itRrZiEAgeCbr+AcRPn6/hqLbBxyClIaCwKVHi/tFCqHdqq
WfBBBvWkmHrKzm1VM81oZcdbpPgx3Vv8e6ZF7kMpqDGc7Hs/WsO4B/A6MIPrTsA+
yBYmgpnhe7TkR5x4qPAGExC/zhNeF9nr3Pz+hsS1F9R7KfEkzHFZFVJ219I/o3Mr
62JGGs6aRmvk+edrloyiqMYOqEZ9B4ArjdhXSB6bTmK9W+FuKtJ/t6+R3gSZU+xC
sI4yheHYRVgz8JR0jHTo9V/pZWCp5HYEY0z/8NpZnYDCEwSxGAUYkWxZ3LYIHfms
rx7EKM46N1wVufOHZxUrUH5f5fgSQ+QLDsa7QVbDSGI8D8S+eb2Ln89jEVZaIw0f
A+EsiLvIBR7WLnJcGJF97bMzUmRpEIn8X5JGaeTOuAZnRD79uqLrKUDnPz7Q4pnL
SvucKflvH4xVIoy2N2o94YOmsu1ivxH/epG/EfyC8ouBKnYFgTH5gxn0E7DSzAEX
MfGUUADK3yB8D3LjoDDJovjZWX26/TIt95mSedZm22HLVkS6+HzSzrA4O5oIcOCi
PPwgDJljto8/aEyQEMdg3FgHU6PoQ5lIZsvnJhdah43yh7Sd11Kp7n7X0iSnAiIl
+mlBl5GJPIZuZgND8F0p3inioFEez4mOcAxCKYUbLUJkI3TzPC9AVzwiAzPIGTjp
vN7To1CvYfl4MCviACfoTZSLvRojHFtGhDcWomLZ3M7SzFq5kEONaBce/KgShbJA
nmMTFWttKZpyJDhZbH6ZvvOHX1WXPgwAa6H97PFBu5BU4a7vs5zs/DkGsQe5IYWS
CtEaBKmKTh8MhASMT+9jc0oy+tj0z8pmvxftE6RwJztIG8cL902HF7+7wibnKhJD
9P7pq9dygZ31E41nNS9YhN15HT+Rx/O94L2XbhnvuJg6iajC/Mlweup7Uw3Eh0Lp
qiKRAq+i5Vz4XxJFsG/x3uHzyCfG3Yd4YWkI6QwtJ9Y5QmAWjoJzOfdrBj+6rrEx
sLSrBcuc/07VXRAvA9ZrjiKlkkTPAqTvE/7ND/LnpjX7CUtsB4312rWyJHA8uMsi
llC+IBy9+DXjt6b+FLx1dgq8+G1bOar92uoji+Fcxd+X2Omm8BB77IGc1M4Flloo
7IxPq1JuIS7Ghp06ahPcoHR4xBNM5jEJdEFRFUR3UTIkdPGmnPft5HeuqCDTbeo1
HR0k1RChtnGEz06qWYujmgq8c7o71C2XpKEwAmUm8+cooDZtvhtIozojWFON/GkJ
GKXWHOlEtpbOem/epBP1xe0E6xgo7OuDfFm73nsX7OxQstpxAXmgzlzsMiUY+C0w
q24L0FtFxseCgS9vwFh4B0ns3QWYQXvbGxodeUxqNCw2ZUGG1YTLllAtJmtppy70
3RtmD/aEnuacx4n9qOrxIpXXss+0lX77FHGhATMYAEKoUX3DvlqeWTWFNK+5AC9t
O8HmTVoHXxISUxwMb5XWJBHt7mxo7YYiQ0y80pl4umItn3D9AOU4H+JQNoFbEdPK
f4pPpmS1atKV2WwaSYoQTuGpgUwh9AIN6dON+yOtGBXhLuOWJsfeHlpeGTLdjxkO
uuT7LnrvJKKCee9nly5XQkhOcq3mZ6xI74rtgC3SP6PC04VNaYpyWdBALEhR5556
R8lyiSjHN9rn368oxfx/rysTsTL5ilfLa0bWCSpHj27bvasT0MgOj/ZanIt+Nf4U
IVGksH20PQxkklo2SKTEBO7a4skx7RIK1Dpgyd6UNLtbXo0v/UxfNjkEdVxV4pSO
Tt9yHMzHRFXg3xDBuRUheG9Z34CRUXWFk021GJ0/XWZ72MxluoaXSvpWXiye4h7o
l7LnFoCly4SfkqFCQxVTa6qPgZ0XnFZw+2SDi0CVV4v7Xl4+DvaDX1wuAc2RcbKE
Yt8h43FDejSllSoSDtKjIUyQH+YZGf2YKzur2Ua7ySLAdrW4OjmtB77F+MHwpaIf
yvRwcVniuzhcYId/dJnN9Kz3w4NAzUIo3JRoUxWTOs6WxBrL99W8jCw4IexVffgj
snY34//3qwZkj4FcEbK8FXmgCn7zGJq/r0gKwSpsPVCoTBS5+cOtFpnfC6Kag5zE
R/wxEgoLX4+I4Q8nuvE+6+TkowQLvIAunHdjJ69wAvCnvXsVZWUL6ZLB1ZBktlrC
d9HAt7+m/8aMyeK89cI9mSuiN+BmSvzarq+niqfP/kp8A7ORg5Rz11xOakslpp6C
57/94jhiMaPN9aZMJMmLgxt6neCN8MeRo0Qy5N2V3731LM7jgCI0i4LhxU5FI64C
jGE9XVmsvT/9AohciHCHGYEU4OLipDpvfbGdwxbwp46wuxTiivqmpXgWp6KdchXb
oWDOKcyq5tfbJT5TYdl2F8tZZmbYrWz2aNkMqKr5G2rh20EundiXdaOlNYtbXtTL
/3pBt0kOBruPQVoN2wPn7CQVfK7M9Dbnx/nKcLyZduPnrkt5KCRuTVy/RrYoZ6PM
dnTWr9RDMS88ox6uJSLT69JAMHi9s5KhnPpDo8C6U5VG7R7zBJf1dbWcIg0G/fBH
aPy9DdUmUXvNX+HiV9JtZp99k7/9wU4HVyEevllpsQ1S7uZKJXbA0vvlxSoFAs8m
CDFbxmkCdlx36q4ZIi7vdK8NoJqOU7O2I+PSK7+xFQLVd7SVzwMj6uXFJt43HHWC
W0qyMp+w4AHx7Xe1pYrkMYsOr0DsXCgAgyXacc/v0xP+ADGzYlMcjN0hzzzoBYYs
pK6vvoL5FAJt9OTe2fai4O+9JETymr40msdBmQCxvx+Rrlz9QvSva2yTt90aytTG
2WKXMcAgyDTJkn1vY2J/d7V282N4FthEVEiUyVANlDNXV0WuYNaKwInLlJ7AnmiB
Z7zAgwBiaiwFGqGCUYfCC5moWF1/uVWeY0P32Em1sCYSZ3gL9GxgdFKs2P/RdqjE
3Ndu9AFjiBlqsAIH2hMEAnwsiQt98EDD4pAU0cFU/gqj0JIZB0oMuks7ON1i2RMo
X0lhkLyvQaX3LXRfN0d8qUAXpn/Be5Yf8LOJop8oZxCN+TnscwD3dVIUpvB67LQJ
MMnD9i+bXRhch9wMdX+p2Hw4B5ZLdv6YjIP0k0NiNQqjE6a5nzZgOzVCndv9/Iz0
pDa0TXN8SgGfFK6Map9PItn7eJAIcZZYIhSkneOuKhAEbuclifrERIW8RJdDuOoD
5edY14R3kfZo3PYWLygOSN4Ih0k+mLoB6Zss36VqTdInE2fzKcbilWe2Z7fCu78c
ybkijnNZEM8Pd7I/ypbjEmnDetaVGBU3VikqD8vkH3OznE4jtDy7vY3nfRiLlweB
ERzc2FKI6486QoddMQGS7Pld32LicdhGBr1WKM/KPpLU+ZeGfNQgtmCr/jvoAjgm
QZiXDCsJgaQgb6rxTRM7CmhGmOPdGAEC1FurKY9Vu7nPKfvjRdkbmJ4aqqvb1Y3t
rvBOECePyENdUXnrqYHQy+B32K2jvXn9kfEn4IMuXHejSWK53p4EaXH6dKPvf/Lb
ptpPtckCo7J9pTOwfUu+W+yidC5aFDEWUgQ+J32jsoPwEtGu9Me2o2Mg6TDoG7bd
cG75wQiFzm44C9HOFtNeb+QySW+MpE1QBLQRuEpI5WuVQSICOxyubAdciEnflbZm
e7TF3iXc1qeM64VfaYfwH6AxF8pW3VKxEnups3GoQcN7ZV8s+8B2DCvzAmAmhlrx
emtw61JSR9s+CsEHyV12w20C6sIdV81OIw06bq/uTwPNrhmc5K7XdtkcdviNayFu
VAzw4dqd4cTywZxAkv85qGCxX+FvLgFApeUE6PTlFENRknVIGcrhby8pK2ebEoDw
IVCIJX2eI7gNCUiyHxttbs4XZ0fkmWOVv95rqvrLrvnao/a6nG4sLUEKlsvT+J7t
rFdyRuirCMlmlRxt/eSk1YOX55pptsQvuUq/2kh+7LnRIE9Fo+cvxWtSbMqUm0LG
G/2fYTJI6Yxp1799kxIVyGEaY7m76XmpexU6DacNk2Xc5EwNJvx2G20L8uyCUYxm
+ESqvGrNYk8zecuTTBaw0wPZOQ05XA1E8reswy2PEGnQjOWltP0rp2jKtH4OF6mx
V4MrqD1Dec2y6d7b/pwchidvo6Jz5kfmtmcn9EMsqAtII425ZktrFsz8272oC8Cd
qYAHJu+lfm1/95Yr9vS3w39lNFZiAfzRNha23Al6FqDifIf8jIUOwAsQTcZRUJGD
y+JD1MwEdrcd0iKkuaytFVa0aThGcsTV9w3THNtGsUEQuukFqDBXZBzo8iXNvIlI
LHdj+pL4D7/ZgnVQcbBZhv699nhzy2fsWewoLoA01aAVwMk6RVirBNUAI1YjoO0B
13C3AWdLFBdkEi71bD3ZbFe4zw55gevw5WIJi9G5yUYI7moywzhJKAcpDvCmZ0m3
ldmiL5n88ej60nsb/c2rfiIRNGbHBXrf8whDuKK5LVGHE8iv4oByjSna0slV3ud1
yeDGWqgh6/FZ7DGL1AMtfF6rR9mKvbYZbjsIQrPwcASdd+Yu3OB29BGnYGUZ/MMz
oyoV4TQbRBc8mQEQfTpVrwkCIr35w/puoOAAHdiquRdq/MBCh4fai3eSbEj7L5pM
CGAkD02gdn65JI9QcocLtp94Om7j0dgXnNypr9+9hrRfdvKRLdSHRWE638QKKZZ7
dggCC1s5rpuWT4XYIhXUClDDgCdWvb/o+mV6ak+7KIWkV4b7V5zV98I1mmD1KyWD
UDKrf+QPw3niaFbR5I58IvrR+Pg+AIk3KEw3HVUnIgSM3m8xZiJ5AnQiz7tnYjGR
/lkbbpIRcDe35vmOtD3pVAAa34wVmDo1inHGbJFAOUBiy5plKwzhjuzRrwQISuDR
4mQa393h5AMIdAHbewvgX9/Gwm4n7B4+pHyKnz+UXKxlcXC+ddJvXswlRSr+ZBDb
mMU4rCGt7tkOTmD13TBMf2Pj/g3WtSb2ABFurmfFtatzp9+p8gBKFEYqOwg6wKSh
UlqMMH38Xxwjh2HUwWVUpgN4Mpk1cWUmVhk8KQa/9DAeZbH3BsZai9cfH/QkyhQa
x+BJRsISMquv+DaVTMNbWdhpSw7CsXIh85Q+ZDroeEZBab2WWTuXY3icJ9wt9Dt/
aAxv3G2siY0SCWqmOsjXwgy8Xi6mUt2H0CPZ8KemK1pLMuvUQELTGqAmlpEQGqf6
CLksjQvFJ6Ygszf7D5q7hJnLRx9LNcUhURlhc6vI6E8C8MSDs1H8IGCU+/yvVELL
fWhNGpuRYcUuXf0VvvfkAQ9Z5M2EmNMArChGdDzljGCNRkmABiDBWVkqg+dO6amb
nVFiRN7nXbex6OaQotxJ4BtX78bZGIWIb4tISfch8TPOLZONriOazeXqhoXdxwrF
YjIXVdHC9nZywhDjEEq4BICcFbreoPK6DZl7GCKabFTFy9gKk/2B0RHEwHU+Kr4T
uXkQIoSMpSu5K3luRCoM6RHi4cp4p8PlLZaTQrooVlDdARwvAtI7obUGTu6Vrmv0
JJn1w/ISM2cQ36HTjdqrrpMVrZUwyFlJYrZyU1HJih9PC2YIif+GFpZM07OJCnhO
/y3w71eN10mUf4UdZglWrl8LcbqHPlieB5P1nu8x2ukqg2UGc3NTGU03+5ABa1Nf
GI+plLTFS9sa/uU5tkz3XGiH9RBsC4GJIGZSPbOhHcYx+5FLWvnsaHXmpeHazKZb
oe5Cr1DF8dkkqay+D25C5GtcXu43haK0Cl/gFN/HDCvaFznec2nU0HpKPOr3WoL6
enw6QmqEUvg0dod1H5xWqMaBM/1g4qvNjP0TP63YxLwFa9I2SIzBB2jKxFiTpzOq
dGZNSAO5TqN1qYoY9yXOfVGVS1Qd6T9WKqrv03BLpOMdyZDHk3iKyWpxCxvhMhmL
LSRe567i2Z0BTYYEIkjZf+lDER9q1xJBQbpenR/SHuIwYM+whHE+0mxzRvjLi+vP
DURBSdZRViCIT9VSeAXjU0zx8OKH+A/mU5Ekdkokk3ZSQxBXFDsEI5x+OVvJ1CJn
5KL3P6AyaDPelWnphDf6Y5NuRBKJh5fgZnKKBLYY61AZnA19epRMBp+xLT+gHXlP
pMUeEZdNBK92mm7lgD3ZL0GRTXfihtn5U/8gfykAgF6WWyMvQznjK2DoM2117aZH
HcqWE1tHkUEB33Qp2K7W907C4fapvJmqZMYx1PHT1vxhl61Wz+XIS+zan7qVfl/9
rHaunbJEGAsmMfIurrHArBX0pQDmAaWzIUzclNeEZu5Hbwc26pnxt1ZtYPt2ca3v
SNP1K1AkQNuNZeX2K6awvcO8N5k89xJFCex2EgxtelNp1tAvmdH7guUIqUFB/3Eu
KyIX8Kozd8gVIWInZ5eU1Josb/ESCMot7KcWK+bqD/rUv+YmbjdB7GBTDWG+a6bh
lSvEICPcn1LMcLSnrTQ1PQ7KTdRUn9Rkaq9/9WRVvMXK4eLpbzQKWTlvH7Gjo1/L
XxO18irGajCRtOyJ9vEwRlQpGZcb8lEEGOTC1mYaQY+PfU+9QBfYGuW7dhTn3qmr
cjv7pFIKLKIq3kHY8ib6JJDOxLElyd4+INMXeoBvsVxeGFREh+K9HchzyvrupEB/
pitwRvRJfuu9bxSxAv/LUsNoKS6DRYV0Amqjl/PwYd3rLb/A8SdnQCEVs8XEDEDR
pTOq7EOPcxuo7nrvaLCxMDBhfgNGeUt9OgE3ieT/yrEFU0h9ukcMEBwoyzZPUtsW
SWezjGL80EcBpIT5qIqlW47pvZ2urI8xFJgPVnVSWj7Z47XKfmyhUagTLmpf9nFy
yvBsIaCHtnG5QzH41MwvVLK7wbRQNwwTn2PICryV89Blhm8rT9EcUot1uYXALFYZ
syeZSiJ0U8DdIhOYluccauD88DWs93cY+wN8sm2hXYFhk46l5wcCfmMzE2/qu7gE
bby/xeInqgLLtwlP0DO7P92AwLDjj6k3kHsoWjN1HUzrPof+EMssMroDCvqfSLVN
xeZ7IyliMMPQBa7sYdPKFN//RPOvBDIBOWfNQzpcqZ+PJ0fwJwRoeqV9I+zEw9Us
T5zIBtEGND6pHX+KriA8tZeJ0xWO007WTgZL2fikHH8D/meYVgF3uFwxlu8CkVv+
GxHsdmkc4oa+DAeetGAko1x8zwWPDuTSEszigLIsIreTtsk6fQ8slrJmkCdV6epE
1gvEHBj639GKGbJMRctHJDL39yXt0SF3gQqRu/MHeivuogabHWOXT7noQc5M/HS+
+5NdAUd8mxFLiGEqKaTa4C2BLceC1kfn6PqPGjMSMpJ7BK//LVJPU9UWsP3L+bfe
9UgzZeELRY9Ji6uMOon6q9mmNKGZD3TC9s3VxBX1IlNFGvrPcYCcooRxpXOOTdN7
g0Up+DtAC6vqJaGxKBZwO1PgAAI/e8uWovKHK7kruO+uiRh+/rD9piJl28JtF0RI
8LmbRQFtyoiinJYn1S55qS3a//ny87EVvZJ/3AZ+o4nThGABEis3xSVTmobrien8
LBonhmNC+ZS9qdjXDjeFVinTEAR2lTF0t2Ae5z3GcCzlwL/0yAqEmeA87qTrLKc7
zgxMB3hehlxhp6NMrHjRn61tdxeJh9GPbtmlTBOzaVqG31Em9+ZiNWAcnGPMbX03
qRZvC5DxrtWK+pmShC2m/MVvfXy4wqsVu7uzZE16cxkt52PqYqOPutIkWE0cJVHE
QcLmpa3BUuozpf1j4nnHm2GEkD4mx/SwmdxXUyBPSBXX9OkiWhwZaqZs2KtobKN3
b7oO4FvxU59JcL+Y6SvmfxshUdY/+rcqboToARdEHpsawyxcpG1N35F/Pyb+szth
DLBzWL82rY5zWwmC3PEZVayGxD4k+kulWt8xNwgSh8zuBnQsxBZ30e9A7FhJi9uW
aLWiXzN5qTURg8mzRuO24WgwaaNTSgFevS65V5ltLwnWnsZ51qwP4Yy8+DXAug7t
9E7y50gSG9vecQGZP5korGUnadvExjpoBi9x4HDWqwyH02TCMkjkuNjJfdGFWc7P
VI1XIRCJUSXQuwTsylPVdaKZ09juB25w7obee/OIzCqJiQNhuufoXyGGjRw/H8kT
ypPSEWJQ8qesJYyOOlTbAfAaUfcSsHcWQ5nsP3gz30RmHSF7bAUiXvi1hQCiy+UO
op5WikHf3Qz+ws4+DBiOM6LrgEzPYRedX8WnKh/FAaQuSj/+s/RGJoqoIOOXEkNT
E4cjYPApUyJrnSed2GAf/1w5NUbTuC+1q8yd3KJhskNAbveKtqw79RuM6GocydCT
q2BviT+/lmK9Kc/IjtZP9AwOdfpacHIiHfyEicb3FdMleUz84eT1ByeJqSMd5OFT
ylTvewANX6D6qYq3ElcVZQs2jacimZKmDbG+C4yOPi9B5Svz1JuMMVV54jNHKTD9
Vs7fHMLNgrWChqAu2KRoXKTVZD5adY1MmbuZ+lZ33F1DRvrIqVBpUnPCwhhCJ4e8
obiNuNd0+fekGooH1uA2ISHxmyWwWhh6JvCTys6x7qivYcIVvjWt9Z0B3Gcz8Em7
K8uVBsBa6+F/eCGYQzr8gpZ0/4mRodHcv03G8YrX8m77n5RwDO7hV503fvn97zpf
oN5PgqN58bloeJ5+I4GFHsTdQ8U4Kkynnlhs1w5ZrmK5YuPPTW0B0IP8MfnaMD8n
xK31xzhS0j65zXWPZgHiCDPUz3gkFmu+EoEmqX+pVFWg18tWDZ/kDC8pyyvBMt7n
r2/+5h6afk80ZpwWdEslw9SU+qOqpiaSL8pYemCzm3SYhcqtDLoaKaeO8O1/GqIf
oSaOfRYScvEge+45fFu3/IgmRTUxfcLWv8C1+F1nbKpxnLx/9d//m1qlV/IwNkHb
y8MvLNP+592cbB+lO3hwPz0sQ9+VfjrHzAdBu4fq3qyS+hTE5tIwvBLl6o5cMjBu
c+fO/f/w2+NwULP13J4pS4hznnrtkZy/TS8IE3YeCY33C/V+fzjxkfb4br6PyevP
mgYtYsNCl2Lq8kRMjHPK9Z8rGSDXf72qEqzWgbSuWG+WLX7hrWUFAMpoGQw2mDLD
FawNbmTYxm1GLH+1HKflg8PAIRtqheWD1XBuL93M2RA0s9waqGWG+Xdx3gglXNZX
VvpFhRoZjWlBRsZ4jJ8T20FYar5CPw7hSlhE3zGv1P50hmopn+KLSl4z9GuIPUIV
WZEIKZ27VZayPcOOBwJdjTY6yI6fdnXZMVSrX8IdzxZ6qcF6Gsct9CGmf0O8/Fru
CehGqGvbybjDDPlZTto8ftVjM8a/iqmnWHoVoeI6hHfoS/mhkKur0FPYoDK0IbEt
bZiyFsiY4Qzv4LszAZbZSFCDKq+BTBJtEQiiivQgxoL1rDc9pUBNORgr6mEJHeX9
z5WVzCfKUFCWonOJPzjm03EbydcdliU6LsqhgFT6F6khnD0Y2sZAskdvCfJIW0IH
yYaNQZWscAGkUSp++o0Foehx/W1yoPsVWaFObNxX7wwSzGOG1bFjeYGrjGGgr50b
qxB9M7s+/V6dQ6X5/D+RVaMu90kV4YURaV/YHLRIW+SGvhlOYY4acL1iFopAqWvs
UqS4YFogS5D39lORBDZ3MIBA8NtEf77y2FvTRJbBU5z/gWPNEnlOYLkSOii59vz3
ax/nNk0uA3mqivi4JybRJbBtsXHNhWOv6wD3h/Q5c6XZtNxE4W3nXbwEPnW8royS
C9abSrXRlTD5Um22MLIzE0ojaC4qwT9lZxnz94U5LzjhYKxn3Uks9IxPDmzhBjgS
qlKOoO5TMAz0jt9wgR6tZFHgv0Ffxk28+C+MTQSeu6vs8WvXzKekwGicg9diHg+i
B8xRZVfKoyV8WUWsR1fJyhGMc3GuXKLWpP86O43prWDE0KwOHi4FmGC//9tDGiZC
eCz+Nw7673OLrt2geRJ+6qYU49kRPsxixY3tAXRYhGM9XWiz90daVa0WFYwgd3DU
MUqNFmNVwLsXDssqUAfPlkdEdyaTlRwXGNt+KJPyiTGdK6mqG+pAdxvrvtNAGUB/
SZyKCu/xdAcSI9WRbEZ840QK00WXS49R/o3bsR7VwId7TjWus6Ln6em9n50Qp+5+
HH/QKKicBCfaESoIpIlC7hWH8kz7octwma8TpnVad5aEYQXCSDH72Rp8vus1V39Y
Bu9XED4v0X1/jS+PogrBV9vRZZhu/r/SeoHUcdiTnhfGkEpLna4rjozuyo4IsnGR
umzO1xqvit2O1piV6pZr5gkRqGJVfJtXmd9eQ8QMFOV4wbP4iSyXBvKN/JX8GtLh
R8+0KPI8nDVFt/7T45o6NsZotpJKk0I5mRRcoxpG0W3VXiwoc5FGWacmzTDb6zsh
926FlV3vTjKMApVTslffFYCWE66C1lmtrRBWolQQGN6edja7k/KwmrwsCwJBvElG
wwtxHH+VzfhCR1kGTH4hIVWcjzSFWqs8l7/gvin4kqxhTXkiq62CCHALVcX8wbgi
+Ac4mqfQhO34fAXG46ml2z9bFOcCsIERP85n42m1uV2NPkkAjev23rMFzTlsbCOK
H5qkkPV9pGHf9vdKsOiZdMUQptxOx1EhK0ELVPjt4JQlr8BlpSddfCREvMU9SBc0
OOVtaeX/Hc5sFedNNex4yxgX5geg3qDrE5Lw7ZkZR4J8IJxl0LVIKInVKBqyTRYU
UPPaiGlmSif8Dk2NmRl2nIgpwEsrJfomR4dU/tNiOX2gTat6quALKSsmMyovwDZ+
7t6U216gDpp2pJuz+FDEwfQ/WJ6Exh7mPpTgGgT48QVSVRgEADNYvX+GT3jqXKRX
Mv4mVviIhR/gcoS3R3+bqvgwT5umYVrF9ERtdns0gdXSLDwSPBHhLpShzgo0L6yS
caNaCBOo6FXEuSGIp0BSeYC6Ag1ncn69mAK2hNeu30SAMOzUR/ifNJNlAmCs367c
MJo2mCDIDkvAUr5dsvWyhHUwQ3LanYPvuoTtKLo1HuTQEDrw0WbSetxe5WCuhGTE
QshWRCGpMI5VPsko37pr2LCHzuoZGi4SwXHqSUez3s0E47idNJzkcy9+CDzQlxEr
BjLHemhIdPIuM/TmiUY4fDMEOFzGg8FLpchqe/7OZqmgQcx1aYdkDJT4IJgubyrF
nhN40RtXtyTJt+mjS9zYfZun9TFjn+dzjxOTITvLu8MGUlUSKOT3mK+NOSwd718p
ciJVPkerH4f+D4FU5QyYPFUkl6DdxLOI25aXpS1QZMADrwVcjMh14M3n7zR8YYtg
8WGHFZGmAdhNgcLGmYLNwVHoHQPFCbdcbVUe6BP1N9Lf5eMBZ6H6Bdw6cNsOEKWn
9Sck6gHWUMoByYyTZC3bFIiaYCq/4NaEFT0mQNY1DRV46z8g1WqHJ5ClswchJv9c
uJGBJhqVAhjUNCIeLZJ/WLqAD374g3HoOdrs7aSy0VKNcF+7YLmD4OkEQrcJ2Eyf
fpXL5NtykfQU6BigiBEk+VeL0YWVPd9lYO1H3PxK5Osgg2U52F0gV4iNYnEcskW7
D8r604djr8qCtFjamoiM9lm7SnVpNIvyqeNa4bln7QWXt0zWhXuzrJ/IpJyHwprP
g6hLZIX3L/3f7eG9Bufev0jAJkCpeTtbgi2kTNrga3vgoZalyKWIadZ16U8r+AmH
89sB9OP8Sx6YP/GioNWgcNq3m90zxxb97/rP53Y6iOiZBS0YT18hGLu3LIueI+MX
KGrnM/W5Wk4I+ZzPIzqQRvYzXNsrdlzPVw/LMpN46LTPOB6yVaZjJ1b7OpNLwLYc
TGGR06tSuB94c/9fwdFwNk2dudunZpknzzuUH9fspddGcjlmKG9t56W/uEenWkFP
Ve4UAadyNoGleOp3PgSsr7MEhtKz8g4pSZl0Iu8KpS3MBojHzy8JnfRJ2PuhkuEO
IrbnTet4KIjNGjYivWqenZWCv36TzzVzUgL3fHDgXrz3lgf/ecKB54sYb8nVkfhn
G0aHaL+tdB7fzBsRpWP6rO9gVKR72TFv8u7Rtnt97F2SHDONXWrOtkMz9zbocqg+
7wv+tjhFzTiWLH10hC1BNYSqyub0pIURyVIEO7HJ+JrBoVIfracXMpVNGkzucCQm
Cl7CDDHN6CqTK89Gg5AP2NqOMHzNv/yeDO1sMjMMN+6OUHHnOy4RL+NgOHhvbrNr
cf3NE1FjKTSplVUS2Jkla+CrWfXu6s7PlhmXxKwQ/YEW0tLWxtKstNBitCvL67Ik
ao4WEH4jNLY83v0yFHwBumoWCqzoM9ZOvVtMo/CTZcuXqoRPW3XDNGeW44q7NXdr
uClcFZGHixrBnL5HZAgwMq1xYjN2o9g+jQ69KFV8ZSIjY0U2xOoVsYDyweN8YhEG
4UaWCpAfTfVmJ4j8Ra6nbA2bHKwoUIC5Cdiu8Ey9mB09NDEPcNZ79+DtF3KevMwk
ZJLUr21MHgmb+Yr1tPlQfgy+voPxFn/fI4zxeCu3W/jhNUGFRV9c+Zytq6teQVfG
rVkzd8Z05mN/DIO27Hpz9jtfIMa7ngfgPiDhmQ/tbJ8XibCJ32wGFeh54crKAjAe
IDrkXobh7XaG+nNgGlV4QpOihTMLD3UO0jARRCJ+AewVx7eVMiERldLQB922+uk0
R2VeRmZNNsfatNV3H//C7Op98GvF3qotyH/vwVQRSqkOlPcy0s82B/+gSvvMFMAt
S7lTJ1WmYqyuz/34TWjbgGrEDdaXv78oO0kCORYNuzZPbDqOv+XMay4bmNewXvAG
to+nYOzABTPk3m30WjMJXAsp8nCdHBHs/xL7H7DVkMwLRAKESEtlF5QbWoNP+I/f
CzAejDUYxx6cyVUewjRO/MGgAegZSdbVzBH0F78xVOQMJkdwBbNpbl6I31qUxT9u
f7kSz1lQ31qRZmoHN27/Sv9+hALVSbjPb71MA0QxS5vPCqhC0Nr5TuguOiHRdTQE
8vwRTeAnJ++xCmdE7M04AMoWiSs1YsgMajNyKqF8WNsduGZAQxBou0kdHxkKKhTv
sYCCmJ09OWn4k/QYg2cJHSpI4UpfxegJNjPNeg8NmuEqb4mFg52iGeB5LXEJFfyk
5d+4qHuw6/zH853TGnXY/auiaumoyjw0VUlFI2NH6tIA79swS8DC9u6ZN7p8QxF/
HS2dk5IpV9E7Du3aXGXiGbWTz08NFbL8+FtCxF8g956Opy+R5JLOoWCzy2khYxeM
GGviWPm/FsnVQJemM9wB81ZlFAEZ+pdFKEPRjn1E+NT9pRDrfGLYH8O5NNRmGfWZ
VRm1fzKKTHuSSasEmQj7UGzAS8vYvdPpV7B+UVOGshRJ0Jahhm4DVJNlcci6Gcu8
cHk/yGx26EZBnvkeGZcN1/i+iLfQoCOaDhdgCSmDGMb4VWWYEeKw4aMgTRB9p9OX
Gn2QvNZKRi+AOyPDcL0jivCDEXKMU29AbJgEmOGgfvRsx7yiLJWFaXu3g37CzmUZ
4HcvhojLjzU1K2fAcfG/QX0t0ldsH52q9uKhbH6mUVHPz370j2yHh+N1/DToz5iH
138wL/Doowa0iAVMKDIKwaJVPVWBln1aIvrls50C+8u4JudjJSNXkOM+4coz/5t/
sFBRoNjrQa0PfBzQClWe0idNDDp/YTfx3tP0Qxhoyq400FQsBoNgasFe0XBPI+IW
kr+Y+0alI73Wsrl9pTShGVl5N6X6QdSmngpZEg8SXOZJobd86U55YAa5rKf0O5zU
fcm/2Fj0smyF1Go1VTIjqebMjcsQisgPD7EwTE2Cjpz6euwA7RAlnuz7bqcFjj2b
lZNL6KskU7+0AzcRXmJBulncYjfEJjQ3Zpgb9xYYTOf1TnnQCLFr75S5raQ5yB3s
MEmBhxr3kU3oGnAqv7Gxjgvhz+J5DmvvHzBLwqzeT5wzNmpHoynCxi+Q09f5LFt0
Mve0wzz6HZkRYWeX0bY4zB6zg80X2zMfqqqhVTyEdtuGlDqNg/Ns1BW5PT0VDMlm
lOjzmt6QaPmKp/BuAxwWDqUxrH4YoCxatPq5qoIiOVhp4L/bG/0fhmfcP7mQcsEn
JRs9ucGK/GLrGjQX3zwlthzdnp0MbAvvqcuk2IuWEk0dYNaACNgrNWnEl/vUejXQ
CyfyDcRyocK2uGFVsCz6JYP4tUGVz6L0JBW2uQbkdbs/eTiHGiEBw7sPGPazYtAB
k00rjHMg22tcG3Gfe/5ppxYydnIjk5MBhu18Nl2kOt/cEbHBxGZMwiMxaQ8x/4zt
CcZjdyW657/J3w3wKXtpPdSQZ3FYvYDYM2He5ChLvLWT4SCbWoNZ+kLUOSjOYhzP
5UJsJ3Xf8BLlFvdNq3EBIV6VEtWh0UCpiTUMw//OKoGQOv/4Pxax7ETiCB13VvH0
CEU0/QsEMPpCv73LmrIJoLTiGYjYbTMPos/NLuTMFf7ySYsU024UjTnz4+PjrgLD
oBK8Qc4ZkjCzBwAWIzrfXCVordtO2LD1AcRHO0KRMPqOsI/OCEwUkr+8A3Oa1r2h
xAL552BqcGdyuTz9Qx7YSOgmtnb53TgpilLLFnD4pocqGJn86YsI8/2OAGQGgu8u
Vhxhr2GEU1F5XRNHeGbHLZhe5wLkMkskkJi9KKAXZ97s6nCUOE85xdHb3PuOuGSt
w2J25d4qYgM3nI/1y0BHV6VSIS2Dcl9+vJSPP5oUqD/2+HvrsIFBivDj1d/rQ/nn
FpmDJ6Ilbnl90Fa9b0rREDjSYoJQf46SSGzakGntY9g/5Fr/S6PHqhcBfzO0sEj3
C1PnuZCjoNhF6t1L8hvv6uSSK03ZjmAmBZlvOvwta7N94UrQV8yipksdJUj71qNN
ci8WM75HG86iO0qNDwF1G95ei+stbU0bxjqZ+PhHI6WT7OkaXFieEwhQ/Nnr/ewX
G0wZSxm2SXN1EOIJBODiZOdbajE8TKkQoZMVL2VZzhi6ZPzqTX3lb0CrkKXnrELg
WGE8E8r6K7bR6pJakLyeVw1UfNoKWIJZR4jwOJLVp0QwcpqaWn4/KVq72J9lhs7c
h6yNJi7YKC8i6rQ7R6Em+ur9gtSel4zSKpj8nYbQtBXooF8AF4EM8uMYPpNYdFyg
Eq3JTkIdmkZhfPN95Idd4CMr0Axa+fKI7YoP9i7hnlAzrw8bQB2F0rXcl1kto8JF
TZixejPmm+2FHLEQ6d1WosCwrmWarh13xkqkHCkJQeVkoon9UTO66t9gbdfXfir4
xgFWGc80zeEd77Rn01ouWwBI8XGu4LOFBSwCGqMSyqJYOuG2IRfUOvXKgOmA6dwO
8efLq083Q9ALsJtfa0fOapPq20VYjoaMg7xRldKtJUDqub1QEd6hAyRBYsujz9MN
wnhqX13NGPxyW++kv+rbH8eESKS9Z2Pm8DgQgLGvnDYevLfJen25fwhWC90EHRvp
RF5teEc+5+Mvohu/RPB5Vu/LveZqBeleb94SgrM3gL0TrZCM9v2mfuPEiGvzwVtE
JbFyZD5sMNWp2DS2wdjbAgzjy0XySextf2FwYOv6lP/Jx+wAmQ6l9k3cMJzZBxiw
GoKCF/uLdsWa4XI4TLD1MBdJpjPQvi1wp86yo/rMNTHjxxibb5rq9d5XmGCZiuXp
BtnzSWIWxrAABn56zglsWuPMEgxYzj5JF7Bqb19cjmrnIr/jgPSWlgAws5RLL2nP
3SCTdqnIh2TYUNUVUwPLxwzV6P5avtHccaZwYUdRl3yGLLXKbcWocYNqGPH9SeM/
Rpp4Ndb9WixdoSfDCf43myAldhszklm4fkRC8OTqq2GDmeB7+teqyWIN49XPsu70
Dms4vaohLXoSgdyYmPOJJqhdIOD/L/6sSKpMzrHB5JwhgFbg4hxmMAY0zBDLH3Lj
q8hYD3B37L3JxQtPnHdgf1yINo4hP+iSCTUr+nW4WHC8cHWfu60KmgKlwkwhws6F
bBD/F92iAr7pr30ZHRYFzRqaFMoLQgfLxWDWlNkPZas9K65bppvnWgM/wQ1R1MQW
qFooeeoqY4Plbwg3eqT7olSthwir8DLqRcs/VqXgDH9NPtmWE8WnBo6mJws/lGHt
m1gmzggDJk/TzVIz0caMAQ1/bUr5XSNjofTFewe+pst0QoIDr3m1jq5TeqDax1c3
WgzNZUTwksz81su6+vDPEtJQilZEemPagIjEP2yIJtAM/JV/M3owd4FvFUCmfSiZ
aOOXa57xOJYbS9cevNDCrDQb+tUMtb8tV5U/s3xzOlyGtA/R7yg3vkNGE8sqD3FD
zgxEwFT97vClYc0IrDSeifLpDEcNb8tUMc+fEoUd3i6vfaBpXOXF0/OVoX/Zy7mg
iWcB8mKnmLNWLj4FJ+gFZhJ9vukkNoKXsuUfEQiIMotYG4qM9to4Vr1gCPRdyOAA
WI0ZvXeCQtf3hCzey+Cp6/sPFYVf8AmNkUHQCYFmL5mw9Wdx8JE4w3l8hk+9QV0R
5w8ipJdQn/XuIBSKAhBq/nRadwvF4V2RDpsoLDvZWl6VdlnbQiL2XF47TOvaFf2i
GwV/EBoD2ptTp1/Fu3Iznd7E0worXquD5q3qtXPzEsokjRFs8Ck4k/AO+p265IkZ
Jf++DPxPcjhYU0QE7hgQX8m2UcZMXmqbN0tSZUhI8uZPUIsHAZQn1U4Bsp46prS1
YWlhFBrp30/REzqZn20yJx8oiPJQPvkpBaWvmVgS3EwW4c9D2YBZ2jw3rG1nF6lg
VkLfI5Z07x1M1xdXqPWqDJl/F1FNE3lZcfpwCZIwyfqRBjDlkJRptHpacIysJd41
pb86QECq9bYHVkvB2KG/op2Xu6VcIc/GG0lAMLQ/OX9n8ftZrN4RTZQfeI71NDz1
2dUewTV4+ozG/iZ+ZkadQw7Hl+mUJN0qgNasv4CHbJima503MaE2lEdAJjye9LMk
ad+UaBwpzWV6ggbTd3dBJ44RLcoMNxRk1AavXQM+EOBiYDnyDxVbhVhckZbMjoQv
hTCJyXofgbbAo8vWEHVr6LAhbR7hBzsTOUeZpaXTy2938nCEmpQmOrRksUxdOsqS
W8hSUfqOb8pEplsIFTNE49fh/STinF4dp4YJVTMjDe/XtZm0J+O2Hs/M3e4R1SSI
qlhiXPDF0dEdTTfO0DVhzN/0FQk+tM/8tDjakroV17vfYtPtVQ+wvaa4GtBnNg6n
/DE/2LGJN9K7M3ecC0pkQNXVkeu+zehTxwqRvAp6BXD/jUzUsi/X2IPfLF08ktfN
8jf98bcEvE942jw1z5/+dnXNf7IcS8+/qvIaw4mFautKIkXyyKIE4W0sdQHKWMVK
K+mK5K6g+fuxdeIdPlCWr8cpfsZxNsqTfeU4kf1ogqjdLP+KL4kpXd8d4u/ErZYT
XkMcfk2oyNk5CZuLp8bRluVMILXl6Tiu+m9dxjyUhS6S6Ic1dWgzjBaADDaXHqpO
fGALSJgdJD3LspeKQI3i5NsJut2SHX5Z1f/YnC/6dEZ83Ox/9UvbOis4x2w/Xaj4
7azKggV5KTtX2gcLv0dGY2Alpi6nKXb0RLXUusstswzx6vODvtEgZ/qIj/0ZqT+J
TJoXxypOM/EY+qIaOZmyihOP9cm3PnosptET5NEx25ehH79QxmkH+scInMJwV0VS
VVOtPuCm0qrSQsBIa00pSHGwncLoby75gFKcqEMYYBqbNVdGe+HcdW5YxicJitSB
BzxRMRBzLLgyMFBdO2KDSA/6NZN4TEKsqx9tRp+VXLgn+ABrHkk/FKBGCFXGrkjR
ZXGgCZqQ2Yi5mrvthSMWXi+LeWxtd0Tn9N63rksycS4K7dTfvVRiNRAZRgsTHRZP
Ch90BQjz60SI/is3mq21hJIsI65Lx26i7CA/7eGJKVJMyKzhY3u/6l4rl5oB+d6M
jNSGbRaGO94qdFCiTJBGrgm5fJuVSVY0C3K3mxa/7tgkqAkAZ91nzga198ZYAIJd
LylXqDYemPnry6aKiiZXCGV8zKe1bYh9aeH4f3sCfa0idudUAcUxpMCvKXRyXfmM
CEA72igr+5xBFgJZbvf0bJtFiFlVJsOwkfbD10q35l5KZbFQUsY/f8C96+Baa1PZ
i5Xl5+Sf/VFEpeLu4Wp7RXCgOTIQh8S6jdZJq0Sh7qwukJ95I10Fsu+mWP69vbxO
fu6pvfJRhe+izTt4SBhn9keCbc2XR0rl+7oe2Tx9AzFBccgYXYIAZz5UrfM0FbLk
tYtmlwRx78f+n2C8fw97ATZekS7quvn/cbloFTr3IL+GmepEo3BbxpRnGpm9422+
uj/FnnsJWlKr/LSR90s5+Mia5LuIaLa9Kc5wNfy1zavkg4wEc/AzqR49P0S4bYyr
dHcVy2qGCS+BLXoI0fmr10XXPXLjYaFFQZJPDW1P3FME27Ud5jYqSZqan+oUiYpQ
cy64h07sjJ42k5dFkWsNEGvhUbMuK2mqGpO1AI0oqQCpoeusa2ZimmegUhtkT95Q
WhbZVo0XLLqCAA+6SzQ0NJ84hyl4pp8RhorHpCNvydNnzponZ7ZcyD6zW+ycrQW6
Taokqf/j0L7RpZO8XrLOqGvJoPcvm1ODSaoo2a3ZSAquLQD5biMICb+GT87X8ksY
DEDhBVHcu2S2/hyzjm25F9rVIuFH4kzWN0hBhQ5SYVZUTc3F1my9V5YIHk/+Ko2D
f76MWpEYN2BzyyfHogqvnGzc/6SGut0LaA6MdoGTaUu8EBVX5SjaSJnkcev2Owdu
n9Qi47c5c3xwxHw6GIwuOgpTgcwOxlvNus6gwtxha1QSABj408zVCgXbJ7hGgdfO
3TCZjI+7Hy//vxzw4m9PprIK5rhT2yU9kOD8h0AiA6E1MX15W853puTcxzyfepLU
eIDIAMLQRwZ5zvStHEuFJNRHdAQ0x9U98PoUMkuyM+9F9/YRVBPOIy6LJ+UsanbA
0Dd/o1Cuw01obnTw8leRGNfpnNU6a0IAPd09swpYfShqSGNdGNXJb1gkPkPQHix5
i/UFh6X/Lh3LCmp6lP9BUGiKHK4WpluAor7OSgd3iWa/XyODSQ0fcwc3MTNKBYUB
wI/EFfk6PMvyuuVKrbhzUp59oMktIsk8HYjSHwp2RoOrPFVEzOU5++1kkdc1YpnH
51w3HSTPnd4z7Iie3jgCwTaMUPqXv89B8XZ2E3nVuR6nKiOu9h9yeT7fHhrTOxQ4
JebyT1y8nFsw5Ffm9oZb2rd4N5/gqaQCsOg/8o3TKGWpolvzzoCm3CMrQ5ykkrCn
63ncXTiS8kVl2gljpXjkxTNzfIvbmpjMGk6zFRcBxaLpSo8bCEV/LkuuDhACPYmj
XNIEk/lGvrnUVU1LIyi/pobAuMVGIGlkq7VSwfIktvyeAoFZdamO6do7JF14Bi5/
yd63+v5sMKb1l1vIXToXtmdnlNgSSr0QiRBAaHdmBGrOd5mlhw7VbKjXOrY/KbL5
yc8bl49tGx85QGdzbDbvvNRvrlNuhIn8GHgjzR0TKiWyKc46+FF2pLF4JVivCEjv
0JEUiOoEXMAVse9BTtq+UuLhf8oOeOJ0wcTo9IfXPnDGUtcVuJjovyiEnZB3+UbP
p238IDECjf1dPwvGtaXCJbuCgVbRp2/lTwDZzFlSbAuQdXVQphVI4VCPZfEKezUE
u3SzqKW6D9KcdbFQ4kndpE2QAcFAol8Tupv2dKFiSINYtils5DRPmkbmMUuipUY7
KKUWW/8BnKbDfoLP7CVGeE9U95lP+8NtwXKnc9Gh5m/WdQ6FdnfxvTYBV9314CpM
4RowmnzF9zQSYtTpqAUf6mIORcdTcZ//mGUvzCyHzGXJNsL/S+ibwYIxf70xMmCT
Yah48kK8ZEI6O+ndI9OYVwOlFtLCmf+R1HSDW+W6ZycUZPuZTZsfjjeHHWBUcp+c
wskDUCvHQp23bMuAWcm+Wstrrq6uguJB2M8RNCYL2YYG/D8QxzI19E8E6thmTeYA
eTRlbPbh28Dh+BlNd+/tP3pa9ZAy7EOP42c9psaBZDW9J/O20PxQUrft5EYSYLqf
5un1H6qGcTdcNbNNWlsxIWk8NVw+cdCLWRBJsCYp4famO9ZALFOUpyU4xiGZ4Y70
g5+nCgVG1k3uirhh4cWxLuy3qN02aGy5/2NjUpVoXfAp1+AuYrmnzBvsnuaf4RpX
m+NDqoHyrC21vkLX7b2SWxx5TQDU3zs9os6WqR9CIc1wvJsy9wkMxxF4K1TJ2EzD
gk6XFQDUfhXWRka3grKQqK+xa/G0IIgGKCu+mU/muo478QhpXvvVFZJ2NkXiW9rM
Jb+0m4WZQlxyrVz5nQdPwGf0DgkkuH7kczy1Qg0NatrbnEqtwQ/YjmHpvJXQ2mXJ
ZIIZsaWVqHKeT32MYz95hHoj8FBKJqZF05/WqUZxCDmHI8LztMgzVJ+4UzZfjfqW
GGP6k7Ph4Jp3u986M1ka1NxooYn5xjnydsL9td3+w/fBkyD+EnyZQA/ATjmgj0ZA
+nEDplGMghF4wnHQLhVhKn6DY5PXiOHtsAG5l6zZ4ge3DTbI8C/edya/Vb5SVNEd
X6LWBu94gqQTat1/EW/LHEsdPu2STjbjJWAC+lG3bmhFH6KsxUG3RtVYmo2+YiPW
fnQbHu9lpOob7xGTPGh3ptzM0VVnGgG7LduhmRnwQG6wS53AYh0qs5KObHdLra/t
z5ra/DG/5SaJZ3hbrNw24TGOXGtHzOTgT5PoVZJczIGanGW4XgQQeqkLRWau9Ggd
Doz/WgEzQNHx5fNLN956YaYTWatW9li8VUIhPMP2hZac/31dCDIVq5dk3mZ7HtYl
Bhb35bRVSYlPyZUAXb2pRnUODdgmBP/SGhhwdNLj7XWlvKZy9sCP94S25ytzegjK
e6M50gUVhQqH107YVL1i2sy7BiMDydLcJ404gYntmuFn8NSJe3PlkphVvlaxVmzI
h1MwIc1IOXzs9W9wEayF/CpD083UlrMMy3Bm3MYRDmbO8ubXQBB5UxfMDsviUugV
N8BWILEv6Fsi95pZCREcEuCGz6PEbp8uasIzXuCTRztNzoAlkm7rHCDThvdVRxaH
uryFXHaySxrEOgysotzrEyf9iuT5E8PyiYDu1JQ7JVGt4IO6dv6QkhepDfxxayd/
2sZvip4qsgkISD5Zb/cI+w+W0c5T10VfFDFDg0OOq4VsdgbjfZO+jqecZohfBF0t
/X4kaHlvgLA6EBXkNMOpAQbn6EF5XkIZ9CGuHDUEZqVblg3HKHFZ8r9SAPe30Jq8
ht8lz7IvE+qd9qAxFAN0mJUtB4o75XC0kdniDHiaGRGKuZznQYE9o5cvzMzX929B
vOgBX/bpO4nFjRAGKQATUCJ/kQJ6Im9eSdYbSLzDQZyHgBw83z9tVtcZhG8pYva8
4gQN9xBS6Y2ZdFprAk8I4HIMZKNH628As+YLb3LBWiJJ3bXwsrnlf5zL0x1MVSSq
PZ9lXfEmtDF96z7mg5qQEKwPjJvHvvU/B1NJG3zaqVLRGkyx6Qkh5krdNPUUGRxV
lh4lIcFiI+Y4IYTjkzSGlxVQIpj5COrw+eJp3FM3m2zPsw+tvL/+5RMq1OyG9ZYj
ZwOQgyttYs5yUIV31XY6fT+kqOJn0H4q1dnwkCExZZ+GbcfQCWykhSevDfBTS3AY
3npsuZx1ZhsrxPy9zCdWL3y5PQdrsIOhEbGYg7klimPTllbNvIn5MCOAmEs/lVxk
FwMm9YMd/1TgCZurZRysvyeCKTcNQr6Ozx/fjP2dxepsofUyxVNInfQLLapQw6Ni
Du9YEo2nkU5Ezv6we9Ccb4Z1Ut18IyhDnkBYkdnzjhqLb+VFemHsSOSVdjP4ZyBj
0Kocpz1VIjiVxdDHr5oG7G6YcPnhy+JRUZgeCofFmzVXIcHtxsrsojKf+nn9uIOA
aNAlf1W51fXYi6GmtPTCUOSW7QDwDv/jzBXzMkXi2LYTlb0l2CCy4OkopO5KF7ZO
IQqBYaB12bXq1K2DhyEN03qOLGMDJX2wPhSk3ZTmZ4gZsBVnLjB6yWeXlSCYqFYS
Rud5DX/gSDYIdS+3kyW7y9wPleiFE8oWuaaEwCzg5tP5UGOt+veLIdQQ9ljZmvoR
QNyNkOY+rUDYTQivqQg6Qdd/9pplhK7rNVv2MkkMtWXc5IUyl6UoPKTNPlKQp5CQ
zzQF30ZGQw4kH7wlASOkeiRBD4s2hn1nfYa7xgW8+tbepPvYaDwQkv5Fci2arvB0
SsC2Y//koLb1dAz0NZ1E6yRajKRxzYbHFfcePc9ALVfky7IGBPIYtwj1AAUxgzI2
2lJUmyBRS4lsp+lOCqP/ulNE1BKp7P7+7Oiy1jX+iHIp9uWGQBtbxp+C4m+Ou81b
KNr59zNw5iSgEfEY2vNkjlQp26quCEYSb4uA9LpkVvXvZ3ojNPN/3LvlZD5MNtCE
KTcsqLS3bGTssWd4DFN5XwEPSDyQSdIwi6BhsqOabw7FxwNiUak80HMrawitj1Uf
uWG6B/l1ZkGHv+7cAwDeY/IYUbha001SVKViIP0Jh93qtCAGT9AN/kZ/m88ltsKI
E9TlUU5r2LTh92pogxNA6Y+yEoC8ji6ONQaKZtmPG0/pBo5SuK5dQ2gckdHBTJ7S
PViYsxajPI7ytd7Hobqh2EZ7la9sQylbAM6upbFKeZ6AX3U8Uxe6OildF7Pgtqzp
9R/L5bOoeM0rmQgu4f5Zug9+EnrMkB5YTsfT/fmcFwUlvAV9kEG87nbhbSGgcNyP
Ohthwker7vkPpRHGXFyBDhmmBeaqfo5UOV9XhVuVdDOCqedFZF/5aoa1jnpuZlOa
zLebvON1vqzOGnNZ1SrG0pSKAdrLcCZuyd4xdSN9rZ5X6XW9K1+ur8oDY2mxFGai
9s5ll2Qm3fMYLxUeF4eQXtfxK/6hxDfj9cHB76lxTgb4WbWBv/ca0zIK/Y/hKVhe
DJ0EM9tRTXE4KwmIM2nkV5VAYoMLooXAHGZFquYETvidUZx+ha5Kwifp/zDrCzkx
O20KkN2q6yNWBxqHNGy/Xp0vyibkuONXT1mrvqE/U6ytCBEXcJuu52vUPF0WByrA
UiJLUYG3Nbk8GSyi6MSu0xAuEfvVf5OfsGlAL25/tY6YZDV9mSTNzRzHi06E0AYj
cP9ia8KSJrojFF4svUJ8rMEy2Do8oimDhG77E7hgp+a0c+aSWd7TQgahG7kkKkuA
Z8DPHyskoH82GofUrMbsz3dqpO556GCuWClu+eGvuWkBvHnBxG18Hcp3r/uNnMb/
xY/56VQ60aeOqcV5ZBiHGW/hXWI5zJZbDfjYjhrkk/dswIRFthe3aLC2E3dEhfJH
ohf9PXpWiCOrtJIfyRsvlTP9EQ9cU+5QDp2mMsazgMRBFVaTE/lQGVR8Efl95JZl
wRkoC+7IdGkK6cCkjtmHiRzDHqB7yJXIp77SlsBWrVysUAQe8J6jY7styUCNvb5o
otqglImjJ3tEASU/aIyVFnBEc/P0UMzW4wkGk04QwXfAaD2sjtdtbPkedIH28Vet
aZoLgMA9+v4Y/306wK608DQTGPv6jE5visi8JBl+Jf1fnjyoqmaujmZNXO4TfRIa
mJN8/wIrgtVXmramH6/p0IScDdvxz/SGCOY8lu1RDkpX9xQo3oUCjtFBHRVYDH1k
KOGFHrGj+AVxH5ZEtA0gNhPXcZYNkEXaOxHWvG8gTPcmeMXD6TJMKZEIqTpXrcEv
u45NiOj+wKxrFPsaKjqHj/a5XVblUsMRKbeeksWsQwbkzx4GEfin/LCQHr8aGnpz
SqvJXLMFIKhTPWenHFRWj6OKhh1cuMFmINCWEpupytIuVFYOj92g7DohgFy0rAPt
9JFlGhj72b56EEN94tVeGPL4zHrkQlnhsJ0FHui1AEpsCBI30he+oiQCDTzbKs2f
wXaYDBwRLbhSCSo9tN31vL7/oVVxUuRkH9KmzShPZJfyAy+StZe92fRKDZonAGlF
yHZK9UyKm95/yMgdh2eiERQlN/lF2+l/IeV1Be/5vIdhzbZTbFWS0nQYWibzDdIf
wnouuVs91sS15dux6yfI498cx7BOoNWmEc2Utg2Jc3N4CdhBScPKwLQbbFuCxqPi
tCQ3aFuyk7HE5N7LVfvcLiErMYJ9ZpgWucgJjgeFr5AUxM3R6UHJbOpELArUX74o
l1mBwLRvENEYT6ttxsUJqjaVmj7T/EkeLNbzG8yzoNaHbatWZKDiMHNDP4SI/iO+
9jr+Qnk3YObo/I3oQShrEpRc7zZx4KBQ5prFUTw741r7I4dcSy0/ARvsYe05nC1M
+RH6FCNYHLiCiXUYao3waAQ0bf8TZjExdWrEJyLUPpXGasqUDPDzOAHYNPkG4Q/8
RjWiRusJaNWtLKMtPRmRs1jCfbBGXS44qTNshC2f00UVDfYj0R6KU7KPeY4sk8Ux
rioY/SdJDp0SJMKRg83pixZCcY3OBQA9JSH7FBstbdbFKg5JWfqaj6auwCqy0sTE
mXCTRlB1bUvPcRsoJRW5HdEpI7KveKVxB+xzZHh+UacPLHODPjBzeSWJi9dJ5ine
IGggTm9Agxfz8RSHYszj/vY7POXpsBntIUFKcEBDLVgYEkifWgA/iId9g/R5b09u
yxDSw/wIbk3+YRpqhUo4kzbiLtsRZJaRMWOnGVmoau7ABMYTLX+ellR5AWJm0wVk
kVWPaXPfJ89iFVxYhMZOQWaE4IuHZ2szmliLxoDT+PmNzpAi5q6FjIQRxFvqfXKe
fQee944REsXzPO6urkJPNtHvbktpVuV4Zn4aQD+rYctwcgPEWbmDOHcfkIMCSX1k
UJBg2VjrtJtTj1qREJbtSwrtWJm07wTYc/IwDb1XkN0IcVvfm7GZnObQpZElIjQC
s3qJf7s5DO6O40F2CFzuAJvgYCMrtUag2kPDc+oXgNp7VkZSZAAxWR5AO8A5/ghw
rlHX6dEaulEMeA+f6j63bCgDrByZ7x7N7PYHq5s8K88PL7e3GJ8It/DPPnImZMM5
0K4gESZv/teJJqQtC6IdPxx4X073oSZnPL7wrF2wcoS/NZ5uP0NNWCd4wnvLgDe/
wxfjAMyE+ra4KX5eBkqR6/PCBsH4eb3ErTFL1AHH/hb4DtqUYstXdRMNXTphRvIZ
g8cl1VAiaw9TZqUnx455lr8kuCpnCutPkeJcsieYuhhdXDKyeZSLP4iMh+3e1EEs
/nhLi3qyNHMqxgX5W7u1V/TZ2ufNi54RmzbykRD8pr4GG4bwHKzoZ1favlfeeXd/
6ghORRVnvFqUzvYYKN1fZXwmzEcVPBh1slqhTMRjHrGV8Rizj1hJzEGkW0NWT0al
qvM3ZQIiumOM0b/o7e9VSU9K0DPVJANp6LrO8eMnPYRnW8QLk9lYzhAoHkacaVz3
oABaDK0RqIacBeKyL91CRaF1Mmhgyvztllp2SSDtE2AcmRoil6A+0CzBEBGiZLuN
iuW8vKwa7TuzxIylj0Sxj6TUcaZjRMzZujhHsaL8hqCeX6BWFP4ov7E8I0bmr6WH
7DPH0j4vlt4UDocPNHSkUHQEJ7ETU5k6K1hHNsGzc9b5oeKYTkFtrRGNiUqo71ie
iJTG3cZx1apimGt8dDUg3a5KHcbHLzqKEj6ve1hWZ1skdq9pch2AvYHHLWJwRtOU
LrYh27TQRNe3N/eFTdsTKbmCplkDhepkL8o2sQRYZLHH+lK8UG/q8XL+GqenjwTE
fVlaoXUnPhMybipmoxxS+Xq7UkQIzuY2a1vWjTAtjSMjBdiRsFMCREM/24eXcPbP
UzSm4rYwzCvnYLTOfz5rRquje0hl8XPzM1xdPYLWFQTSH1TDsDLUCjLvyNAGinee
+jw/mLywMvo3+M4uPreEOS5hnwDCkxfwpJDeBFOBjtJecjC7ZzaQgaN3ebzgWda4
HTFJ2X5y+8FrB+rmLaX+zG+5/vMqLZueP4py3LwDEJxkSu8Nr0u9eBiI549cExlt
WJBcfGuMYGEL9EOxdkxlAJSv30bnWUb2+8hTrIPyZMgybQ5RzmPzEgq2An36o+dG
Pt8jrG4JrXGUg4YdrpicQjpYpwWszn5UqYZWhYuUU0Dy9YbOUdsFn+gIIf+CJvJQ
CXCFX8gYJCPhWpfO2uIKx/igVgbib79XSEHu+vMdJjiQjO3Xc8+pL3bx1yRzfsGg
AHbqCzJaua/NakCe/tgugi2TLuDVtJlr1E7L6ys4s3W9ENJ7ZL+KrkaQEl//RgHb
8w0LLLmEJSWvtQfK83zAcmhFbKYGxjkJXM1tjoA6cSpTBaO0640y6Dy2bxsa2U4d
KDRmsa0jWjCYE7QabQRbDi/2gdyNh5XJt2EaODZtFPi9ke41JM7dIDa2JGXo/iVa
vTU53a/HxNkxF9H3Nog/kAspB84oqNT+AeOg3LgVvhjDoWi+e0vaAKSVfhBK9dpX
WTpMCiHxNls9FnGfRXKbdVGJ2LnD6HYNS3T61QpSt+YAFwgRj8D6QWXZa9YqQ4Pb
8Lj0na7c9I4Z1/90p6+8x1c6SfnsszXIONxwJj09Etd1YYKFRYMExMU5rleu7y5A
QgiBEJn0mWSNEdft1smnglYy9cwKpR4U9On6LYVyKw/V/BQCaxD/lLEb4kdZtFqh
hIT5MhxZl7yMhWMdmuEovVkdENx6Y9fRK1yL7Z6N5N82aTm2JbBVwU6cTziMfMiq
ok/F+hPjlazYz0LaDDZ8xvbV9+bo6H/MPTumxkMXkCjgRsyrStm/i3n9bv1fsp6x
Auet0+Jh1IYyVeooaRrq5o4QRDJNdCy9szt72GVRc3Yw4jzrmLt8JImCBG++7haC
7k1uLP/yP5NeqGszHiB1WdHXr73oRA7Uc3J7J6qurCLUQM3OtDy7oRaxIFbsL9IL
r8ikFyRzCG8z/MBjuJZgumK7O3JzIg3DWjwLQuZ+H6j/LZy4SaBiWSkdNpljnwrV
6lz9Elo5GNoC4Sdu4xDiF8myFIACL/88qfyyRafV2sMKdgzNXwxeFv3diadleBed
cy1LYa2Tt1AG5cmag8dCxgwIVH34eBBjjMS1H07B6R0ES4qOT8PjyTGF3FRkRq7Q
TNPuBsj8oooO+WHFHFpETFLH3/eyy4OzTXIURQFS/sfK1Fzl17QOJzyrPC/aeor9
4C4t5S+9xLou8tg2fnlYn8rRUht+5L0cfwuyo2cLMpK2vhMu1/1QrodLy2/nPQpo
93OF+TBm1JwzTOuFfqXwhQWkHHoDERzgFLbTn5pfC7+Ygl8SW0eMdUuc5AOsdxMA
7JVjFT2/MOVFJ4L0/8z7V7L2lJnoL82OhvUXiVfxO0YPAZfjQFr8MadiKz6Dna94
xj44qc66ROyKwZP5kiBWWjH5bD4js3M0lQPL/XW6YIi79e6erQcqdBu+UnycAgG4
JG2rEeYt1Wg7WQVaAnkZ0VLOIDzorOJ0zpwE+/L/hZ4bu3UqZhCouh5RYccm9x7X
byr+vivRAprKYOPgTjXLT5LYA1UltDwM0Ykteqd3gHAx5ipGW1gcoFFM3ebSve3j
YT8K42X9HVd56WcS1QC5jeYKovSFYJfSrbrl01purzw9wqfcV8JYqgbq0UpqKSup
384zLdIeQeg9UJP59xj6UFHHbBoddxMNFn2azhyN0R+ywMKx/o34YocnngIkslXc
n0sxZ1sJ+BEeR8/sb7qWX1bFB2g2Wr0X43VU+SR6W7DW8Tu4h2YabwTfUqDaP68v
rsYUsY4SsMuG5U+iEF5pfgw2ovm2wE+nPda124pWKLW09hN92pzbj+JunI8tOL+y
75Yxq2s01w83TOAHAtnTsvmkMrJn4AaqyHCWcimxt02truR+gfn5lbdLnnJ+Cxsh
AbBZKcIc56XDY5nqniBv839oQk76B4ysmcDDSm471+9hbupIkO60h39mgUxLt3GO
AnFxboSKPdjM7T/96U/eDdhXQ27+wdELcf7SDuh2Q0NyApa2qvPgJeSdw6EvL12L
fq2MPqODpBz5wyUIrZkCpNd+/4JF1lS7sBZB8h3IvGx4WgOLf3ZL+iH6MZPwrIgH
f/g0vFY5VVfRF+pr2kLorokxHunlJBDgsMid4UpTRSWCDcfOua8R48xMnZTTqIqU
gc820uicsxBZN2i+2JVs62WlbVTQfBlSpqpIr8+jLX8mRXSuvraoFVvSjzGuEXKq
rKihJdOsLnc0JKfb/V+dnww/n8l77bEKG1revv/RDUOkT4G4z9JcLq0kJgKt40C/
ZugU/u7OyN7vhJ5CEEzL1lwTwuO5k1N4UC/s6kSLbM+utfF+xGbbe4g+5ssd1kau
gjsRMiu9JhEy8zirWwcd8yxI9yYGPtAtgFhYkbleOiHNiZajOm6Z1pl/UXAMkagP
3w2Lqvw8c6LTJPEjJO/s8JvyS8Hf/9I4bOzcFVZh3jbTXKXnOrywQeo/VxysC1i/
lKGs7/EY2/TXEnSiINIa1e44b8+gK3CWF4AEmgT3Rfnht01ji3StYcrWYrb0EDbo
8wgkuV2oVrUVAuosaDyZ8cctZR17xBUOhd7lrncDDgiJS1pfAWWol09DpyOS2SZs
cbt05aYERgKtjXFMJjt1t2yq9U3MujwwOLC57eRwyva4XPDmpiND+mTZox1Djjyn
2hdj65fELF7BIgqpN9r9hmiRfXHcndiR/dFYQTpvKml0YfdUJmt9TCqE7p4bqroD
byfZFkcvjiX55SSkPU9VLLu0aambuwYNOtvoqE7WyeCEvvgaNKmRXxENi2Mi9EbW
O4lVNPZUmt+uSi1/PtpbzW8sMT+OgJfkIdSEQGmM1bTB/yUZ0y182oY3w3QC2rum
cnJr2qWDRgC950hMFiIln0hbm6Egy28nbGozM5ZrVgXBsaeb7HmYwJ32apHGe7NV
Vjago5jQgCt31nJ5Hx20SASFADhvoIrLK1xc4hrZKxjzulu8POiKSjuq0fh8xUrm
SsFDCJlyhTff+btjH1PQB/pSrA93xhB8OiEzuOLcMsUwTYOxGJyBMbh0bJLYH7/h
D4LiQiFPidIbGYSADvDOAOcIMdA6e5P/kiXpbFXHsv+SClzpreGlSYU/Kog1FKoh
psQkOAcMy7pNTj+Niq66BdoNq3Mql3y+anm3QR3ml/LgSi+Dp75Ii/88iYPsoEHY
ooaC9eh24RR/A7UPyEDR3OKW7kTGQX3liuSSBw2ZOkfJ9sEPmdqqGWdf63gB6lXP
ZPVCqdecxJQr9IlKBj92B1L6JuGa3iuC1L9PGYcnEnWZabjy66kF8aqhhUCEb6w/
RU+tuH7jOsauMg1mUIRtD/mD4xTDikDvSXo1iDGuhY3M1QbFIy3BzQFoGkT4N+zU
WdPxwNZJCXyver/KPV7xkehNiDS1hq8zl3U0MP0502Q2R3LBdkC9KMXSXqxNxSwG
gqUc4s1ypCQbUVQJDSIqYjIJfbe8Ga6xoj+6dnG6uoMjdNfc/EgQMjfpm5evrURe
BvPl6QagH5l/JD5GGOmh3cFDQKOSLJtvCNr5XKGuSA096GkUXkkcQx9FY7gMRUMT
Cd+5I+DhwfuywMxRzSINFdYjB2B80Dag8Chv1EZKp8VVty4gSbjw4ZILvaaEG4c2
GqQcab5Rhq1y43dJg7rser9hHnktUfmv3IwEw8l1C4+2s9l5uSr3hlej1jVF6KO/
j+fcwxSOjg/Zgv0W46AK913i4Jj8b283vcE9uI+npuPmGq7AFFbTgNcpwSQNSVVk
cXxD0VkmGm00iCs1WSjLTBMWrf0Kyf2xbQ56iw3Y13VEdxQeXoWWzH2l6szPxAO1
N+SvoIvMD7bkJJHjXdSb6K/MpN+Q8i84rB+iR5KFeJEdZjduN4GzfxJUHTQshCiD
5XrRsfW/sfr17D5VS9/kyUrNKK7EG9pMTosRArn9cf5ltJ5RfaW8HOZvARLeE7+b
L8VwxqW8FDnhzSPwaR+FYemHUsx7Xrm/aZhmtaVmra265x6Sx040uZZyU45pTFGc
7m52Lw/gAFPdj11yCqufxQvTM6rhQR8UsaaGgR03HFDjdWrymS6QXGh7D+84dqtK
8nar+b1Ml0V84Cju7UJCywlXPgR2Nz88u1D3bDBOybi0I+kkBN8e8zXta1HcsQDF
RintfLD1ww/GX/xZgWHT8k1ixi+nQPE4LGhFifmJSVXFfpbhLJDDCkR+iRXz+TR+
yNqyVwc7tp7Q3KazlYTbG8fliL5dI2ycj5d6J6xhybhBkN0iOu04Rrp/y3KJvd6P
JLLKWnyZWcTF7wNxsfDe6tZeKHYhP8Cx/MYtIME9TXrI68d6Q5zTLjWIZZTxFXxt
9jShv4Xyt+1qQ0iGO0XWYRWm4HtBBcfwQp4Sj0Oo1eEzRYKGsX5/xjFlWhPrjdmA
pdRbIOCFFdYtSJzQ5z8wDpdJcMydqSHUqefzVJjo76GngeOKOUu1gLxdDWiSVgGp
WZtknwowm72njk+3pwNG5VOsrlutJ2ezDEarK69ZgvPx4HtTylyA1Y5hU7SDe+KM
uDdQ45ULfC4qfao4N01ZoCDRbbxNnqBYA4zvhPvAGeYQnB1B1A0w8y8iC3EqTEBP
0aKkdKG3I1ohsFVtQn9UrbtvZsDG/HpJK5EXgVczrfbS4i9dJhATeusLfo7w7cJh
5GpvYxesqR9d+L5bgYxXQEZ9krNlOmqSZyCbllMl/F7mP2QFXYw7eKUocsOrzkv+
w6pZ6wPzirp17JWU7notjQHKb9NoAPPLreDul7fYTfmBhAA+76kYMpwUeO28OXtq
iaYjL1HOc1if/9FiVwERtnhgcCyp2nhlVm7+7R1WTcAKzyriReUoDFQPtD37YZLQ
PO6U0D/Zhxpo004iZUUHVlQ3/IGijh1VF0ZqCPETQPK1+IR6wRy2XfXwABnh5HMf
L65wp541jWNeAdyPtKLk0cZleCg/rRGAioqA+SvzeguqueSgGkXRwTvnTHik0QpL
MG/CNIvavvIeSVL5/ef4nsdsILTt3UEkFTgtgTsJkZ+c35xh71k7J6oV6w+kMiwb
lWapC0+ynq3y8rKRaeunnfIS0H/w7n8Xq4IJQNKbyyykxKOQ1X4H/mZ+w1dbst3h
yAR2OdC3WktJhBtyMgVz7gYFTTohO3u5znisLSBaUZOV4PTbncku+uZV9cFMCROu
jMbdySxtdQ3ci7pAU53pVNzWU5ZBA4lxi66w+9bDHhJVM1hvgCDtvk6+wr5hZ6gV
QsAdZcr1NWW28HBFKzbGn93uii6EhjiK2Lnnm5ZDX2spJ9omnwTaA9f5iS3b0UZN
rrJlXmkCNLYLnwHfhPT52FI83jGvCoIWDsHZyXAu+h/4tAiUeAnXcgGzR8V578fp
m7bOkTXkQfubZqFpePr61CFxMrh1aJdb9RNGgqP2z7Lzepze0dIjDj99Q8JxuAY+
WH1syIdy8/F2RIFs4HE8CFBYqEwInf7elOYGopTrWphI2oJYirM/pGqPAZM4jlph
Ct7YmN6B0KRhvNwREbZmI6T47fbzsCSWRVgL2mqx4KaLIZDmt2ADxB8xvmpP4lxl
sXXu7psp9xmABW6DhA5pXztg8LgUFW9H7T3WCKUoZmutAV3+gHoF+GWzWy5WiWuK
3ncPWmjK0PcRYNk2DBGMhpvauRoDz6aD+vTWztG+GcEVtnS7SjQiMg/2kcgc9aIn
uNgfuncuxARm8Inv5tlJvilj8lr8M6i5pBzA1z/50MER3kH3gWkExVsls1kNSO89
26vFf+jTLtYEZt74los7yJJlORv+Vy9Rie0sWA145wcjxQYyKAS6dOqvBANDg4L8
CIrISGwEo519r3XaWi4Bs8MewKV+b5s0KQXo+eDyGO0IjQukOmDLwhAajn57YgZL
VTahRIOENrmanlRr8EnQbCeGNMY+fY6t3gt5P7LvKIE85PgQ/7nJ0nmh/SuwTud/
dw+MIIWWmgOFyoNbRC1V6xBXYHF0N56IDoNwTWLTjkivaJ4rbkkfGybXjVTB+rvQ
NOb3//qKPjT/Y/2g94Bpw9XzKSj7B4fuVEkbtNucHacwnVIkqBdn0fWWONRAk4+5
lSpIL8anKYsiXxJA8N1B+I//8h7YamViJIRn667VrbH0g886l2FE82dTgLFfyXZA
FbAVggIXhK2XwnpNEqFEcNjrgvpjG1CtlxFYAqKLNJ+J3880iJsuzDPhOfaMKNYi
uPJPStgnRzaj/s/ybXxRr1WnqnHfq2C2idHyouB14YT8lvTmanorjvhNUOGc/Jw/
iGfKkmcq9+n9m8E/tfQNp8gSaCFBI/hfVWzADrLYqb/hOCKU0gpNk8X6HnoQseZw
77rn+adBY0+RPvSahBEChwywlZ8fBi/RPeG09L1i8FBpZpkF0R3K/RHJ38iTS0ls
z8I+R4BnMQp3oOiUOL+7zRlDfCLG/HCqNIwxaozmMv7FLkeZdfn3isLIyEHjcz1z
nUOjb8T65jpWxTXEJnSMpk6ITqtRCKG/HBUiQCK6c6PWaRA+LUPg/DOjXOSfY7AE
rRgpDSSceh55WUnViKMi6pJaP9MUwwEMEk1dykd/M+GS8J/D7Z9/Lle/nopXOJMV
ncQmBmVkz1pzMNAjyojIrj/74RhjLggRt7qjTXjLpsnUyCY66HF2Xe3RleUVxCpn
G56JsDUZwdViHIgSkhF/Karl8W87tSeDhOghhXzv5B7WM+eb8tDQoz+FevJEEUNV
qYx/boSmIaFXVe8zhjP0Oc9kH/qy18qb4noPw7qpz9aSKYBwBpdRQpH9GF53Jvmc
DgACWSDjMBaC9ZfsMnFwmWQIl217+XQsQ7Cc1w9bZmHncU4P1RXwNKYovSgkEPAZ
aOAhD/cM7zN3ZkHQTrpaMWiAD2rO3wlHFN4IfJ/sW8b/rCDM+DS6DBoyW9HJIfwo
Nb36l0S+o/Qcdg7pr097uXrhMaCDIdV7I1aTf0zRsmkFI4BBkst46OOqnBU/oKKZ
rH3fOWt14azFQ9CAuoS8LnaJ/pZ8B3XAkVizCWXLFAHeTkEsT5S1Atb3YJMPBYni
mpg1KHRCOKgi7G9t3HG8q9sMntOskd0h8St5PcV5rwbRxvdBGNRuMtZiLWJhpeOs
DPsu1BFwqKsfUsA80PsbK+hGeO5TLzNkLXqS0UUFv0EQaS0qltFAxiMrNMx8wsaT
xxMU6oJf/a/KJquJpG4+H9DIaICryN9pgsy+hUhoqDsFFSzv0pTjTmOEt9vqcjK7
dL3SZulLdPQ4zEKO38p9rqgn628hRFqtwLtDHzIxxf9Ny++h8kgLGg/Ssv2KaYge
1m42/pPOr7sxoBQ+1NobtWzXLY5wT8eW0Inw6G4yrqliPQMPqxBQVd6awiHe+qHK
+rcdNrFqAdQhiHN5DVdwphQl0uaBCasYL81eBNBWtdjhNYq2tn0+Yf63RSD2+B0J
MOCbYBM5Too3IARSbw/GB06TmT5N7geBQZaKZ/4CA1Cic9gMuCIghBmB44dVr6LX
Jw2pbra73SuStVOsVMQv0QyKcUjUgV4Q7WWZh0aGcU6UfgFpp+XwdGvL/77U1jz/
p46TLW/phJplsC4oZMuw8wmfl+j+KIzPeHVffi3BFuiU6JszA1MGwj4VZLdXUCXT
KJJROgjOrNqiO4RqHNF9nA6WkrUli3KrsorkyW5MPPnZGASwk9JywMuH9U4cvf8a
HrI0UVnEMNS25TqZtsyz8apDpwJZE2CZCWiHG0RpZJpTMKbJji9Nd5NGPszTFGbk
H+2wIXAXLJTcW564b3YhFUXxrYTnMDqctK2i4KoO+Xeth4K4mNWn4VMCF7UDA4ub
XvuolnPS0wuSrfOaWoY3CKkYpAGx32oMCjpLapuN6LA5lHbsZMWss5Njeb9bP5DC
eyiW/5ZHcrJadys7LeL7rSthFVmvWHePdvUVU7IoP5Vc9FI6nLaBctmlgHuhRaEP
oN2rLjwI7MJPtXRP9HOH1bndIHMAxYhU+UH2MRwnHfBmLqoI5d7FDKdWbxQtkcGh
/Cl7LEXzS0xCiHs/R/GyNDbbtk64c3ik+mAFriSYEwnukVgYsaz55UHSnymBjpdl
Rfkjqjo7V5QKCOIIrWcSMEOFjvksgXdkwVctDXmtzi5qYmRLREL7X8y8ZlDrm3W2
XExnPIYhRhGymWiQ8tMpHkMwlUv+F7Gc12h1bF3hagMUBByQFnjnJdp0iiRVsxju
tlKB+M0a3QJm5iwoT4rsi2ojmBW25w/D2vllhRfu13LAc74+4VZkZw5oAMeB4fie
DuZ8Dwf96IdIcGLXGTFNp5+4f9a1vGy5RROSJmYRYups3j2nOdQTxCec9U1snpto
LXKv58BLapK+ogbR3wp/SQbcNhDKdO7WnVz1ZWAOREFQ6Pdl+MYyLJbTudBfknQm
2NRyasirDmOaW7yEZfS+zLNbDUlnAQ8pJghVY8ihT9DmPQo4hVvQb2TDGPTvc07b
5ShBkzJnoMmiTmtY2OUZP7rh8uSGON5KmmieifeWy6pXclKYB2xHAMf34XWy6h2i
zAwBD7fL0Ybix20qCNctclSZxtHptpDMHR6DmQB53KPPcH871tI1B49rsBueR5C2
1t8kNFqL7EfGVUY8w0tggPkKrkxRuK3O62KqDCHGrEVE1eHwI3IrmtS6KSnd3amG
9lwjVkzzR49r9FxLdfw4Dmfad2E45JHsS7vFTK+njOB1CfiCZSZ18MeEYJgAcZ2v
jG8lDev/Q8fzLDonwXjibYw93qXUQIjXcObSFviy7pGHsgmjRsgnMCTruNucL6jS
7RD/BaUgdSO/fRznYHZP/kZ5zwJpIFnm7stHY/jlY3KyBO/D19P9AgyP8Rhfsg7H
E+jrEtpqWBj/cWo6JhR2ivOW3E/Pu5ldx35kY9TBGgYVnKxldGPzvgPLNreEOWlM
9PeWf7IYsikpm7H4jaUWZrx1o+JvvKQMVorrtuvGn7WAarUn7eK1Jsi7xCoeNf2I
e8AIx4hHGzN7KR6fO/y+0zVFCrba7JyzVvhu4MWNuyCcAeS2NBSPd94W0Uqz21lz
lP5f8PZbVZT7t9bQYDvtqF2SKq+4ODlrw3zFa4GOf8GpN14PU8LxyrJ4kYQdfdQY
3NEKMXfxC1Yuj+YwAWIKFj+H3+I1hv9mMgWWVirVPIxSELLtKEI30AZ9FePoq8B+
8mqESKxiomujNYKUxvzfq09ifsgheiZG0CM4A/ALk5lerN5feFG7RVzSXKkbVqQl
vXh2iBWEAV4vXz+u9e8ZCR/doiGJDzy86/NxmRJpL5Wjn96ipkdRE04AItKmYrEu
pFejgZnioda7Vy1UVAqmwrsAGDdgoHGVdTC6qI9iIRt8Q5QHRN1O8nbeejiS1qOB
PpQqiZclWfHWMe1tGnYgNuA4Gh84Ewl+fxYXMuxQUNZOMhpsbd5jJXHOYcD5f18m
AD1gT5yqfyjWM7LEeKIfg/QaCeLRNi7odexQk5Nt87AyHD01xjCK49LsO6lkaXGR
tsL81IUlXVblRtLs2JURSMPiGC7pS4YcT/9ne3WNJRykf+ccL4GSInpOxj7v0j3o
UIBZA7+Ov9uETzDXhEFKLgOx0Vy3mUog62459hk0gd10islujqO+XgE9LwlAu7nW
5aOADkdqB3BqlPW9r79hrfD01BhxOuSy/NhALOUSBHFprrlJ4xK8lAlEtL26XGtz
qVG0/q2s13RhXUC85htkLYT6KnCZAA8TlACTVM4ZoGyqQfHoSW786VAELwLYNXSD
pguULyXRnBm9BcU/dqDz6OSdb1XILDUD3tULBLO6mwg7wmElNbUpWOIJQIOLwu5s
NJ+9z2yg5uHU28KaXVQ2uCnqnbhSJePnszCvT/AGbaVLq43pjhac6WvihYzG+QBx
deApUVJOSrkTISgbgA8YGleSGIKoUsWdL+5qKA6W/V9eyJS+lG6kpkeZoFRheEqO
MEWe2ajO58JpgZS4nYEFyTFxuI2TkNx3opczlJm3fZPLhlOG7TJOUkF8Oq7CvH3/
W8TcMQlSY54P1eepa5oAqh1RSiUNOmPHJLwtapKI9GxiC9QRX4NUzBNJD8V/Aa/7
5OS/+eOFp//UsDV6D2OQJI7rL7Ep70O5sdnUyryF3vTPD+iizI4KArtOetJ1kVtr
QeaUuLvd0LyyUULNwNLgfmHdhathXToju50X2UXOXMrtwybD2ZOQyPnR2NLc4hfq
MSU8qlK9DBqQwxRv4eRi/1Ws1mpudj7eOgQ7vfwdciREKdx/HMkuoQDeJGP5oK3r
oMNb4syhxMYbmu7kFc4ePdDWkv2CFDMsi4LEAyEavrUvgtVCDAsDA1pt1XwTkHXj
6rjbhK63AZRWHs1Tjo5N1gYF/QXokoyjbVJPEYJnp8PQ5SJvarLp3LaukWtL0YEV
ZSveY7ShcBXisxjPbkH5Mhvlf7wtwtZHCdmgiBArI6GpIkNKYxKsUPJ9Z0VbUsGn
2FRn/6B2tESmzG76F8qrPy/dL2g46+UPRR41JS4qcT0B9bMZYXuoGmy+/CB91zly
NcSFEwMQvHwzFBLS+rIAM/SGBOGH7i2tezg7sokWHlI8hErKNZNo2UpDSGL7Cbcq
L4+iOjZS4ZWbGXOxRkquGFde00t9kJE0jJORU7fgx2Jamhy9P5M3/RuqyKTipyv7
yZGQa+aXTiljpsZx/bU3is17W6cOpktvW6LYLotqxUIe3y6lkIeZFYvdzAy6aOdg
8dXwwUmNvMa7OkAXMO+b5Izp9y/Nmcs15AI0InDSN88HZJTGFRHPBkhNTdCsoD6M
w5tLkirzjU5lQBaSUcChKwSWwAS2FFSlk9u1tQxiWlSriPud1ctRnd1dFxdKmc2o
5V5c6jxu1JyPxPq73FqWjzB8vkiPPbpdGimxWrK9DRSlja/W2EMcxZyOQKgIg0+e
ityGPAofQu2h542mEqv1iaT/GsCpjznFT+t6WLHUAPcAyLV7VQXERozr4oiceV8u
DovEFF3r3zelfncSxAilwCCY1eMydIvnG7O5Y4oJhiIbcIJVFgJ5xrXSecw7BF7l
m/UySL4yBIuhkNS8DbWjnz3wcgkA+Tdtmi/6mVMXa40loyqK5mnVpRP0p8mPYS+G
EdgXxB1nnkFVHngjIXRlIWLFyDFKsjAOdzKnO+tELvPSSkiNReaoNZeidMtPvMYJ
NLYzs3EJi863mmqIGAFhO05lSjB3rNoMoQnXCnMBWuvWvL5Gb7jAlfnUHLfxTCEP
0jHHcitJgROOpCJzq9ghcxNRavgD16SQXXVfo+HpyYdI942y6GK488B0asHaVsAq
v+bbRkwYnBgrHsUPnGUX+y46xefg+tWqazRDi6UBGygoGHJKB2ETbL4eGFkrsYp/
acW+ArzeZ0lcxa3eV7QQntzrnZo8NqzoHOXgL3ziLpA6413jfV5YPjeD+gqFeRgp
QzCpGHMG+kRW739doKVzswe3+YhtK+ukYBGcTA9/JucvGKZVUQa1yHBJYTV1q3me
0sD57a5Rgo3YxhR6iwOEM2Y3t5Bm8nksrLtiSqIsW8Bf4TMNk6lgPWpGW+QM2Muy
RlgSvBNrYZ8mmMGs4OtxNJADM9j/d562tbcg+2Oqy1nFyFmYGldbgTp0tTV61P8f
YyherXkDcHVsq95EvOtsahQvIfWuaUSoqC2K9K4ZjH1boJMb4ykrA8FsAjthAcug
czitP81gj+mIkLY7dQsFDziHchJFIQos+VO3W81UKH+2/s6Od44DU8lVXIe0Lkm2
NJqvlImGdgBMvQT17C/Bd8wK+lIhD30Tp8IhVWHTO2meLIKzUDbuWPEe4vrUouAb
S1K6r8VyfUetwwiSxqc7F+2RkjuLz3v2pliETJ4gQAEAVGQvB+6nt1DHd9jd6Q6k
RHm18WddJP9eI1i3W3zkQNvGMm2xe4XzhY81TRo6jsClNkbOBcAdxQWeovzjDK5t
ShF9dTR5HgDM86uCi9bDB/mOUkZEK7kDZnsI/DsNiC2PeWR7VYBHEuwdIvaRMQVl
oNcVXkOUzN2Lf1ISNjBKd/EbXupC6xjgHGx6+v6DItIpP/Gbu+P/B95i8i5LkcQN
Ss62Q1WxIdNtygM897mP6OOG7vOEZXhqvt9ZYikx13ZAOpmeBFK1s1UI6JcP5LXd
y6h61OQjtMfpVOKCk9qQ774c2uyVafz0c+nvAabtC2zeEbBy+gSaREJiWrBecWA4
YIc4KkcGIt7zmch/j2Intj0DQ8hjylHHAj+9Xo6xJSFQT+wuMUKQSxyp087CqJzM
hbC7oCnVwVFRHRXuIKh9aBtkEzl8WftOTffvDTeh3/MvpvWjY+qRqCKVTi1BtIph
UoCuFugMVxqGCuGIdTp44QT0nHpfnANon0Kz/bjfj+x1hwdmkgd02bX/ZPTHBSc3
wmLBulSsDsP2xxsg2uLMbJgyHa25Ku35/qmvqVzLRZIdhiicwXxSCu8rO8Q1nmbQ
YUmm96cB3ViZJihKie48XN/sNkB68UWPePEH2QNS2xbtNrIAcmX3reZ5xRTWdPeg
Om1e4T6K2qBY9Up1N3ZjHKbS4IX975I3hFeOKyjbFXXVitm49r077HFAoX1V6o51
cU4V2iiFqXTMvgQgYXOYtTAT79uGPwMdqijQqIA1a4in/9XtNQB3RKWjG2+W/Fc5
BcNbBfWQyK9l/nZIQzR1zhYPgCbqY8DkPkznHSY4f02cRNrRAJEHD6lyNRhwdS5d
jbEMbz9oXDlhhW4Tq+OhWhd399g590HvsVXj6DEKi4hLMOr5zvDOIap1L6+QttBC
8R/0Wc0agkDo4ILs8tSLBvCCEQ0G0kayW1gB5luX364Nl9pMuUMGtqF0Vp2oyJXu
GZmF78bMRbImFbmRXo22aGcD6lpdPN7ObqCyfqBsyA2aB1uv4//JWwVjnIeKnJ8L
qEUNm1avu8p8AYvaG2xMqppEuDBfF/SNYF4TwJzJih07tQN2cj2UQn/+pRWtoZh1
70FsPEKX2Z4ovgf5mVWeQk9sB3DiI7a8HwmOYPUHVuR49r1KN65UGR6mfrCnV7a8
DKbhko0Wzs3ddyoOCggo2GW/yYuTt4NjCnqjKoJDIdKqxFKyPS+HDErv4GlYIkYU
a0JwvA1JWXGOytvj0llvvJGymGDHhSjcL063hRy8x6Qha0xgBE9xl+lZCHEVU6rm
kFbqkKfFnUeqKkQdHxLwQdLRjuVg+LqsWeoh1l2/R8pZPR5UnO+I1juYGBiOp0a7
LkynT9dahAW1H9YdfeZ/EX8Lwpml79jT154f8/7by8idfldMiC8S0orAsTSwtPCe
DrSxYK9xPnmSFCqXeGg+QkKQk1WCgGjBwpnuc9ylJubSEGswaXNZTPgyC8G3phKo
dU1AP2E1PcyFslNX2CM6CgQcPqLT7fZ6F8QXQRaZ3V5YzWe9uSifUk5kgeZGmwu1
p6EPJh3c16ZRQog6H8dICeDmYCJaVptIaDupBOWCCRN+9JEGE+4cTrWiymWSwgc5
lx14/19+sXZAyLUB7xQ5/Qav03ga+W5CdZVzduWaX976BjQq+YmwKEfCRe/xBUhs
9bY0dKO5pxLxwi/uSd2rg8L42HiZ1/squN/ewGTNMeqdjPuTIQX50/fKmD3jg0yI
Dm5vkLoUkbRCFrwawMMaLlFciRxk4DZryBWJYE6bGOGeKmYzMLO+3OOsbmmxTpnG
igSc/SXa4TxWL3zsO11008Tfe+goQYLfndv4n3fnzVK9LR0L1GDyHnRTckKL1o+E
HkUKnUkCWj/bTzzj+B7HLY/5NzuE/sVT+QJN0Fs9hC2t6b8lkI5Ou51olRFy/oDu
ntWBR1gc6NcOvCv02G5T2g7oeZreUBuJfA4Q8HtuHbH3dpjxotxHxAckN/Xyhlug
N5sUGQR/8jkmKDruZz/u5H9DjknIvL2nmaDAsH3XEmdt0y7Cl5qe+9jCNcnqqU+F
jg8Ao6mwZTara9vySs8BhuTNuTFEVAuBGF7Bu/0Oj7fVuQE+1Dsw5N4tph2IgeX2
8O1E5mumRAwqu7a3ItDktsqVrraHBnEfYZu5DpXGA2lE6sQVcStDEoWlAgOucgEn
+435H4FAxKb4Umm16uCVfQX3S4ShrqcuGIw/hgWwsrxe6Yz8PRvBgOVOKSTb0l7K
rbKFCAHwvwOzEXR5EnlhWagkuxHV0PAFkNhnSKrbZN/WvcnQ1144Ei9JEalsILDh
tmpSVhSNGX7ScbRVbUVk3766m0KhhKD10F8BQe2Yze1Xsbx6iOhOzmhSgJ0R9EwA
diiSFkGm8iBwvzGTsXOi98UacIQ4ZxAPGbJhsF+963rsmjIj4p4bYmuO8tToJfgb
FlZT9tSihuAWsCw4VJh5r7obTwSyBYMr7l+/hfSS/nDPaLAaASk4rc3WefnYxYuG
4/FQ1/oVkO8PK3dDW+Mhyfh0x/9qXIEMI95uCt1gcT08gktJMcA+78oJDR6/+tai
Y2AXyf5M+LImlHszyoporQD7Bcqg7HsUehZ/oDEa7QbS7BhcEajLi3Swm7C4sEWM
zwjIssSyYqr1KTmsF1u8nR9P6u7gKYIhCnEawtfhw8mv+FcIwmU1EibJwvtT0Ln8
G1tCzBys6h9BAGSEY6L7vIK61bAvahepMJduXElF4mmAzQZfTbNiESck7S59NyzT
ajvUKZasgpyBdUfOTwSFp7uDCBPD3rJ1fpIWqN9ki/9eFXUS0toACWSku9Ak51th
qCc+TJGACvdATzuQLbtv+jYyJdjz02dfFCIxcTqgQjsypFG+ow/Vx73uP4sqtob7
NAU0YRn+CP2zOJqze/Hw76nDFTMrtzBKHFNSazX/eaM3f3xNIPDdFQsBpMdmMUg3
OrHNiXfcUq7dty/F8vqTZ8bi1ZdvYTcZEBweCk0Kzf49dBVmjszLUJvtrG29RFCS
2ed/E7hsT2e6utGqNsoS8IokpmIlFRfQiqJbotYG5qH7L1FwdXd3QZvOFbPA0G2n
6WGEAEEEWxwlaiOccmnRpq28hj44ny59A6kBg+pKzQDhTXOWpZnsvA9sfh6kzPSL
e+byEYSPSRhS9anEY56MJtvWsv12mgM0AZuHrB0pfqLYfIX4CvEycpDPpq1dyFi8
3p5jso9+INN1IaOPquYFvzlerOkx6J77I63HuLE5+5v4CKx4PtSjq4UFvrcyFruO
tZv/pMJRVMRWSLn/VlcvnaGhIWEcyo00k7o4tbJR8bYpSlH/SBfBZr6i40l+WZ4x
jllA005EYeaNUMjfckXfWB+foXpzaTNmZlZ45Ekp0ew6CPORjAjxo5B0TcyoY38T
1PtFGmAmTptzv/tg4R6TT7YoT0KCoylHgduaFUd8n87qa29MGbi21Uj9qZ8PTrwe
WL0c95O7WepGnNyYMJG81FCwL8IWUT1GZkJyB5a6ptXLynTIDlvPjBVXuXnWzzd+
bFOHS0Q99WM8gzcm1zXPLKmLm5+ArQ7gzJenH/rtiblI1lJVpD4Ym95gf70sD6dN
z729YwxhuhkBLhp4LveohNt2ZgfAOaDxzhOCU5ywCuDqe5B2KuljGkylfg96fqa0
7NSECQMz0o2P+Dp7b02iODdpxurYeWbQMR4UUNivLsmlGuoP5AlgWNECbT183Lwp
I6Xz92KL3ZrjMCvXsiLTUrvPdltuzF974IoL+oly9WrXnYwfo6fx2Rk+r34TCgEp
fy0Z69wllnmfAjMbLpvQAdu+NyP6mOikC+cHFKGICiurb4hZ7TmJd21c9a0qSgZk
8FMFsp6pIsS5I3tfp9HFsvqmwsxHuj6TMjnbgo4+kmuqAYjaebFC+tju+FT0Rj95
aAzgAtK0S2209KmUeuTc+zRnP5cQomd6A+t6Dt3e+WamyuCBeG5iJ5j8fnZ1mu9S
xfOtVwDMFUhtfkoGLJ7WVg0hWcBNGfd+/djQqQYHictoWlAnf1+LNT4t9kE1Rvdr
35BLiq4cEnJ0BRM1NzavjiysZYsFWAUpVcfswBsrRaZEQCpA+NuGsQyQHSKZQC6j
1rr0oBs2gXBfs1PH84cQdaYzTYDwiEgfpd+4TM/O2B8ONc2biAmxaczUB6SNa6T1
eq+zPXTLJT4MUJNXTO0DaLlANHcEtsiFGy2hcYNpJORYv9dENjG/WDs/z8C6RFHN
EPykMLtR0PgPA8Em/Ce2ca0x6+sDGSJxCsxvh933zCI3lva3Fc6F4JuHKbgqCAXl
FD054g3m+NnBFNI940AadnUEYE6Kpdiliikrt5P09NL/N5nEb/zru2JtFpLDUgWX
BHtZ2XVZ2F0T8zNGFnB0/+RpiJumFhPGqVznDp+FWxwAEILVD5aELfCQxmvV+V2Y
OG34UA/U6euIUCzWVHfrciUtEdie8vcai6AZzoede9qWkAUdz12+m+O5EhbtZXcd
B2iEst6XvwjjUgKFtuk2eyUkKQdstwYFWwjZxPzLAwG5WCRK2cyMuPC9HhSPIeuo
S75moTFQMvNFGdc4RYn8hKOkYo594Roj6OpVF+CpobqgGDrr9OKfHXJaSy473XSS
O0KYyBl+IeQAOQXNxxXDZY072tsR4f1CDF0pVXnl/ViERKM6m4TxUbDF5korq8Pw
rit3GxOIqPs50bQxp30w2HDNzd+T0yIdrTG9xbokvj8q0/N8NsLeOC+jrGhugW06
ddzJ02r44tm3+lSn2BMnUmq+r5gSklaFZI8XvAjsiHZUIs0bhsLkuC1WacD1GwDx
l0vI8FMMK9rtSkAM8k2gDlH+Hb0UEGSQmUDc4aWFIR6FlAhLpxNUOmwCrHGi5NC2
1TbVGNRPlfn8EPOCmoEj3/Hj8SI3iIqLt4FTvBFlLBf8rxjEQaJBkMcQ1gMiEzeJ
uBK82EdZwEV5i1/Z54UQhKIt3sszhLfrdyIPJ5hbAQtuAvbeCnJgld3sx5wx31SY
wlR2Uoy3hT6qjbgymRipjUPyuf4EDxaYgrotpHKHR1Piqt8z/YtYLOKZLcBilDh+
ugTkXV9J4e1FOUM5BY4cSeziz5xJbb5MJKEN4JOrMk9wfabR73SBAyn0pwYxhOPj
R6aAY1K9hpK5QRwiM93o3xmVwsPq1H+UE7R0Uf5VpVzaRCckJpQKVHZ9xmobxVUB
Z17C6tPZajo52PenTnyBXlOp9H8h8Qac7BXaaufUBNjid2NpMpz7mfrP7pA/HzJJ
smncSIMsxWlHXjHLMfACM4+WGFZSv2AbB4YXWILJLwEYdw8cI2nnBzgn14lowEuC
DElhrGlvLyKR5mxQI4t6fHoVAlgoA6cpV42MHwu8j0lovZgXZy9e10LTMnikiuaM
YlYrgUx2NrZlALRLhSNGikyZEi0Sk1A4ZJqNLApYv8uuJcED6IpzHURLkMr2cAlM
NlCJ9A6As50GvBq5A9sC42tK9nPVIrDY8mO17v07ZPT0EnIC+XBDQ1g9j+1l5IUy
61HL7q8ctWhJrhN2zikoGugQHXYronpgxIVuHbSHYhzWWkdJkAYGMueh5qu3gJcY
/+MgJiHrUJJwXHz/2QQeMBC3zT8F87a1ZrqGNuk3GMo2VsSpVB5ofH7K0BvhpZGV
qIYjoLfoWvLcJwQ9lJG+EeQt8a++qhBJhkDjzFfogQuHUfuCpN9z/BWbp9Wai9Q0
guI8mR4ZN5YVBqiVdwOQYzb31Go26rkOlG48JdCHOfTs8v032VJnhu86rOrJd0C3
rZk4u17x9jZ/tVqLjvuIEKoNPzSJYiY7K5BRbBZ6IYYFkeyyETWskHtj+pXcvlWb
MrVQeOb9Wd/bx+IwuYDcvjevry38N3S0UlBCRRPgxxyarejOrKosWCRDQ8i9Q9us
bv3W/YXiTz1YQk+jG0tdnTDJEpoQFOl99pU02jzCh9241lyTI9A0EO4M0xw2ILl2
F/Hvnqru6AJha2vVR7QwUvc/45DZnvAzoxgtARmCNGK9hSKY5DXkUaXuE5BcA799
RTeb68npaa6tk8lzCyNdIwU/U31kGnjn9RlHG7t3zxaxtGyl/GRD6JJ0TRBs2QRd
e4BMfuLYwvVk6KZWrl4gf63wzQe8d4nGepFkEHRu1O2YJ6EXpsZ2Vaz+x3/klcuI
sh9k1ubE8rsSsXQLCGUbluV4ZGOOyx2yTMe9hv6p8qxVjiSbGGcfym4Yye2VuZhT
euP6CkDoWH9CtmLsEQjXx8HHhXODTIdiOgHmphT9pQc803OYGXMDto2d4N+DbHRl
V5/XFs1D8GOxRs7XDUelpsrXwoncnTdmCd9V2Sy/X3aNNjg1E2n+k85WbzOwtNHz
aHfbQ/qYPsQZoftpsrd2bYROmm0BiT+bugGnwlN0BlOWOvXtJJvYGI+0kXVjxFDY
uyy/FdDb1PoDE4KBZmr2Kjn4pRFh0W8opmkEEhijPsFIQWv+nKUY3Eudtsfzo6QO
kphJkEMh018Yo3xuKqRO/VoowCZz5yBLADG6D/82NPYQ2xerSXIygwV0tXZNqOt3
KWr+HqFKXUUVGWn+sVU1XDtlar6F1JP/GdSGEq7hcS5xekHiARP4ygIi+qMQGWGL
ym1YNA5XY16PLIWErijszn77Uj+MtMJ4Os0s41UsLW1UhEM3Eiz9G23EZLQvG4gn
7CHYv+yU0YcJg38UgQvaOrdAwIkN0ckCL7ksQeQe0kwTkyfos1zRGuicL3Lcq8X/
QLWPcnoPcNZ5owIRX3oF9npaQWgyQk9XUZmbHZz84GFyp8YCrW+I/8b/gh5hRAea
DbQxPH18LdVTKJbXa0Q6xso5o8mHxepurWdz3FRuSaV10CUSaMdpu0q7LIgQ8460
FGG4U0+7qxd7DN4kbcMDs3LxMNAytctGGgbGGwDyKVBzW+IqTIvjkPdYzQ0Uh3RA
RBuEwAUfea9h+kHEYnnK0sxMPOxI//p5Q3O9fwxdzL2B3ZzVVwKMh8nWYbtS7dQA
BJT4UI3CNSdZX0Ow90K4+ll6K2B6aaK/OIf/VnscGA2XBQs1NSzJIasYF1hkW8mc
07mRMdiWN+ODdA/A4g2hkgYUCqEk2XH6tyhXbhue7MQqFbse7hQEEsSeC4MXZCwt
AVpf3pgloRGDkBlu2KcFeXuUm53YuVz6WbMPiFwpXOtlD+3z/ewyqY8raMGcv9lr
1u7prlGVbQnK+xruLq8EWv+BOAkuTZlYyBUkowKJ+rSNXKHoQosCfgyniSx8RQ44
42HBZV4eEaBmKJR1xHkDPAfU06CFaGDuyT9JAcq5xzTwlsDPOcjrBL9zO6QtQbZ+
gp/tjr4wPSB8NdWjgzwnHpSPg96EjeC1bsRPF2+wo15a6DA9BaKeTYChGrMSzwfs
DlK1+6pHyTyRQvwq0fCVZqoOJzc6iFtczasj1KrtgFjhWqQg63yTCFpY+f3hRt/8
z8ToSiIdEi1cbWqvZu84NSClLp54U2ir54VmgrgXgLvA0ZJENZp+nVGAzemhT3KW
7t3jHU5KFhnDru6DYDPJf/LCdwuCKjEdE4heRve5p95NXEfWk71zS2IfTS5pK3Xb
aoEGVoJLvyrIZKXILyMpv8m4M+X5BOPe414aKrGhwGbXvPGR95chvHAphI+oWK4t
exIWc+CWWVVTeHj3YpKq99W4iJ1MkMJwqv9hdBuKu/nL1DJ3pvBMmfqMJwAUv+mv
8CsVo5sEZV0YquSScxvGwjy0YsO1+68rnEXFKcB7BNo2LzrC2lU11FLa0k9eZWtY
Oe3zqNNN3JRvgUt4IAn2uO1N74985ckK3FBt3MiyPBVv260gB3pFse4EX2nOdQU6
M7KA0sAdK+aUpt3eHW2m0ie4vnSJB+9Pu2lxbHAbdyLyIjIFJ67gCSVUgtNDNSPy
iXah/x3BWMc5toFzztdZq7bXn+kg5oobQXvqS48tea23xVV6CPMtkXuqr0+Yqdel
XTd0xOyzmirMhmLSNjOhNuKi1HNcOWCoy7TEkrYbFxZov1OYp0LunKpYqJp27/QW
xgPhGWUjpeDvbb/DHGxMNk1fsLwM68wuf9Ipa5EYcKgwz5NuzIc7o9QSalqrgDDh
3RRsj0O1YqsUDfgz7MEYo6AXgEGgx/Phdk+d49Gx5wepZqDtzz1st7QqqkrrQxnK
aO/2XQwxIdm8l44S7TE50X4qPLfg08uCx6qre4keKIBluv1pUYgolXIiHR0xtOAb
67rQneIUCXSBiPY9IvWRk4hEdNNThDrt3ryzpMYHELl3h28+41VqMB5RrVGyNC4j
RhSg4PFl3WEVn0PQ6nrMx5RviGj533KuwcbDvmChhXsiS01gmCjDmTroWa6lC8tg
ZjD0E8YuX+6y1B8Nchxne95s+H3aEpety/aDotOUTKWEcI0MapqAv1vhXaE/WdCc
JddtrkVV+7UtMdg7G9rHxO2sYr7VzPnYu9p8hgDxjj4CqTl4UWuqVC9G/CmhmDhd
DfsSjM+MNAS2DteRzQs0Y9YCj2ItAL+IKjwgD8BocGNncaXElmIyLXdoJfXm4pSE
0Z/YnJSxueC21KgherSnN/cCzrDOCCJOqRQpIpwOSRK7t0YUmh2qcasNbKYJ+dGS
EnR4OWkqLt7gsP/zbislzlKmWiSKxrXSzjl6rBIv9arJE4W1gF1pmBa/024gvOzV
vEl+PQ/788IAh2HZ/9gasdLgOP9ULDEqyVEsCOSf1Voe7QtoceFkMKmchDG7L5hU
gy3QvVObs9+WTBQ4egBJC2waLAFyOgL/85PEzWzY67fWKw9RtDjGVezQSqSNiDTp
PGpel8P7ZBG+pw0bebGpahA+BZiEKPPj40FBnSwrk+m+AkfjEJnlsC58Fgw7U7iV
+IAEeMzG+bsqdkMyDiqu1zED/2Ag2dGR7JkL2UeSZeNKCyETVBCX2El0PnrUb9+1
S1VsXAZR14OivmMaEC+n0qJBXZADIIf2fb1k5TC7dv3Q07FiAjqs8zqdPBs9N+az
Vu4U+YasqI+E343Ty53yReSY8QdJQHiYrg2bDkdrYomTUL25SLXbv6iJAB5ioNXi
UkzoG/VtkdwBmRqPtdfZAiJmUXUkz0a0+u2+RQshxhQRpCOtoouwp+iW7q+3ohEY
ojMeY1Ah2l4kXw2OdNgEnM+X4looQSi27re70VmR2YxF5Pa8yTB7TflwA1g5IQLs
0mQSwcWmj2tuKhBSxBV31888oufv4e5wrzICzLQruVqgMFVvitOF/7efCppF2kiU
KKkGOEbjk44SUkasQbWCX+kcQfEct5DU7gGuhny8sIz9Uqn8hWnA27g2N4JT22l4
MpHw/fwtbkCBtqhC3PMM4n/wSI5v4JjfMd7NTkans7sJ07Q0gjYoeIIQSEMVQ5wN
H3yEU+HUvE2fcOkn5FeKxqHsF8ambNdlWozSs/ooBooSpjf2pbw/M/OCcgO2vDjq
rnDbBuV1ZWGVqPG8hKozZTLCyX6jRLXTab4LT+Z5tW12tlA4W95ivsxuQ9FKSejr
wDSnZLTjfzJBsOcjIsv1y3b785ntFxLCAyuL4SLmrYO8h4YAID5i2SJgnks6ZKQE
G0WHuxAfxkp9nPHwRjkV5S+Wt9jJqGsa5k4u0jhCalEdnhuMw+vWKYFWDPYZb5Ck
RoyNomAAaiDEJRvO4wby5/IbNNZBPEfbqyfbNmtmvaob5QTqccu84y5+L38HU3xH
1ZyflHUNSk459N2nFFF6S+Whgj4ZnJE6kgvGUV8/Il1MpCD6MakcpKsBpON0z2Ia
tb3dS4XhzPM1KpytNnaiYEhx0+mww/aLN+nh+JtERZBwOrYjMlOQ/cugmgNDMTeI
tI9/Qg8JySs2oLNuRi8fV4vbD5lh12vxNgxofQYKuUtUTLLN4fy3D3MITpLQwkth
kyPPUtyObuJp0xVfV46EbfevrAv3nNaU17d6sQoAivurI4cq7/4udJ8MA4MePXOt
e0mZ1QWwQ8H2/6H0m8TIUskgS/pkX1n1PIJ/LY2Z4BbvRLrZIX8h1yW/nuEIqL9n
JWpb86cQgiFNf2thnf4PpNpc35VnLbqnsoJugpvpibpCKre/p4Hnl0thOFpk+Hzt
NbORz98MX/su+ZGmT+3ukxI7ye3KKIaDMPU1FTfAcqY8izy49jog4k2/JQBkmTP8
lio4b+xpiYjLkHaF73w9xoOQz8hphMQk/0pvUEDZB4q6A9kqo8/Bk0TYvA+q+Rqq
1Ws7KFiT37NtWCB5I7EGN8iy3OT+mpbcdDtkMdd3UesBWitRAwDoCAQsl4zZAsR7
SiWAwGy/tKPD96haIyJco8y7VRWU+WUWs4C0IXVkKnkWp0iRX+CEQlWAHf6uWikB
6RaIqQ7bzH7sII4BvjgvgCCtS9yUPT+QQafNSdUOZsPFihj9FdwOOKoBjzS+CeUT
8dQQ2+uBJ6z8vg1XdXK8NmgZU8IUzPs4ST3MJgIH/Ru2M/LIdE8UqszwglskJCbo
WF26SLGQHcBQq1hUVXyxITAUDfhaB/GgmSe5HQ2ADkPlH9IYW6TBY6xbXDCBsNF1
hqeLeVAngr5nMnjgQXHhXfkfZBof0cbNVVpaciyCBSfFwFpRM6wKNy4iBvxMF33z
GJiuxKu/H4fRrqVL1RPMdTO/A9RYF5LuzZtTYExykJozQ+yEkl4FXdUYLQrgtEPF
+t/DWU/6FpguEEiCC+GNE1zeRuqewAb7kJu43vXRac81uyA/XtateGuUcFj6I+/u
gJgvlJJH7FrwFreZBSg3Pa07rOQJJjWkoR7wr+AGaERqatydIOkwyipF7DTTpasf
rskboPOvIliR8KPKP75XtkUGApTHA2xKd/sZ7z2KJ6YFoRPCzUL0m+UMw/bCJoNG
RUCi40cX5py+rwPkRBwXAI6tDdugwXjPS6Ui6GQ7O+gipXAEHuHtv3OsNAbbKxeW
vzm9K0wBYjQ/CfdvTBMP7/nBC2cyg4/YsbASgJvyTtXLkIO/2YBQXXYv/+6TmLLu
EIZKG9rk9cZbhhbjS5EjJZyB8M1kql8qyc4umNC33lyC13tkbMhsSpRGpQRxDy/C
xyEAz2p3pI72jggC77e2bsPxDKYdSnoQOCKLA1AGiXgciyTD1hLaxb/CpZKzJuyE
tM18GM3nFl60Drtjkdz1FO9Ph+a7gS5LkFHpJqGg7Od7SmQgKz1bSQpHnis4nMSm
YoSMx4MqjMCZ5qULyiQ5e2FECCTKLTVeMn2umzpezKYvTsv7TQwmXLE/NTIflZaI
DJKhu4UCUKGTDbbk3id7hDw2CyNVgw68nsfkcNHoedAfUM0iupREt0Vb0lZpzcGY
3aK/FngEf6tkadJVQGilOOdk1UnOE6D0kWo31jjVqWrKKL5k263TNFJ4vWzlN9Gf
585kq9rhASmKY+IpLxjhZ2dpK/+mHZMLh/62cebz+7nyNtXqzlCHOOrvTbol716O
ebE2CDLJjoBKEWkv+REkukN5IEIeGzJ2Y5YfgaWYLZvTCD+8R26MG6be++87q7gE
8+rO9RRcnn83rIZJZVmAxFzQeFFqb4RguJGBtVnojXLquZJN4PyrQO0k3oac8KxM
XCRFEsOHsLhCAEKXKJhibip2lEiLes1BmQWZfYCadn0v8MPkWmUAG17IbbdLEzvM
GDlxVfhK+Zs7PkKdtC8O5tH2ePesV7hDxfdMB0vYqiKFm6J9lyafEkTpaxUiHqgI
sPEqBHN0xKMBaBopMxonli2r0iYLXbZow6y7941gm7Wu6Aar0yrX0fMjzv3Ej71q
x/wPURDfYAJBv3EujsCiUqyZCidb4pgjZuqmVktl2njKAX9PitC//LMid9PRWwta
Fm0k2itDNkWOtvy89LDYGGRB2qzJkg/HZungCToK4LAdN8QaqZmqT7EXprqBGfM5
2X6/GSAOfUs4jWPWCkgV8A0wkpzuWRhAhzUnQyLVrlUvrCCucLqD3HaHVW1H02fo
dItgIpreFwDcaTvyimU8uIdrGa/Lj2CijGxjEakl4xbyT0pi3JqEJj6bUWGbXoum
bDKvJ4Y+Tr+/vDNKAEpjxNHz0lRIA731blWElP0G1+UU0BWaYVEr9J39Qy/ZJqdF
DRrvdwHqRJleDCexrwJ7hpgYlG1oKCD5KtUbMJ5teYfY2phKDeg8hQ82DS1LNaM5
JhMs25WmiYmTTI8+etRiaa7xlRKgfTWNui8UOk9qSk6wFkv+0lzVlgNw34K/fn7o
ePj0kKHgLMUxxQC3QDCed8nxThDH8o/wQUw/cDTFCbgnQCt04NhUr/KKRWllnSku
FGOsJ/AITGyLxw4iqMe2H0gAH8fZUrvJrFN1VQfCuH0fSgK4eKNJdAM9idZRgTnb
qia6T0LZvcvsI1WTLapjAQIr2ZSCE4KQkV3+unr8p3XpOw2MWnYfbQ/wkius8sKu
VncayQa6CATYKwPAn3NH71mR3lp/2BL62Gam9/dCzhqMBHD17Xbv3pKF8uPpZXXV
yegNgzeIjFLP9kDnty+RUNbgHENTiIzjQxcrOqrAe6E1w0VSY3JvXjBWPOewRSe2
KKfRbQn4JMrpChnIeBg/Jdsg1Ml5O4ZCl3TzscgF/UCi7FiC3Jyea5CV9v2K4NXn
J4SqPfrlS81/5lkCcLtI6YjONdbSL5nLI1qDt2b709HRY4vGvi7aiLoPHNFDtxyo
gesAZl7/qVdO/3Sfi99Pu6+QdZoYxlYD9pNrtMdLNaqH9Rz+t9hY7yV/QObAw9KX
fgGEYhF1/hFRLEiy8AGyrG+sJCAVktSdGMb30tluiQYKlgBV9phe5MgTyymjE2Zg
YtB2wHSzHtA+JuYkNKgQ2ddq456AqkaQCO/PCbg7c9RcWBqGNRXGq/BrK0FtJrIX
LzJO+OT3mlXnkES6VceIuRNukfQJDVU0NSc0eSSjUwnY+oILZqg6ydjSzwezvl5L
Vzx+w+Y8O6X3DlXhOAqoe34+6hgjrgdaAPqXp5yJvKwLDBH0Y2aQaTSFRSimnqGX
/NDNdkmkWxd7Q+9r+RuiRIWRaB4KoBByx/4b8UY3PhLcwf8RCYAO2LZRM1C/7V0l
oJ6ufTPeD84BIDqlxO5kYnvmZc2k+ek7zr0MqzC3CJmjLIMNh5Bcbe3rhRjifOxg
BKWC+cg7y+Jxf9qzxHnIRRiDGCRnTualOQQm1SnEVKi5iQriRph1k2nS6oS6/pab
uJc73y5hqHj+7x6T+jqUJa0/uEFEantyL6Vci5c2il7AiJCxI3gdzryVIKlXeOEp
rG8g3Hq6nJO8qgb0kkg0zpLR3uFz1ScYknFCVhL3O0YxOhXAtu1hLGKgmn9TncJh
qkCcLx7el09usPuqdQPr/zTHOXuBWiEvK8ASfrsBbS+1gC5VYHC7ogzt+Uhd/o3J
Ou2v8BVSe98Kcbsm/3XAgyX+MTKJ07uc5atG5A7ofwGaQijv/OK921d3wtHiDNDi
Pgo94kRTav9oBCPGU8CdkRhkKCdatHcS4gSFgo6Y1DiXLHYGKuyRqtAGKLjxXbEL
coKZBF/Sp74k4+HjfcLn3ClGFsktr9pWUv8ExQP2plZBduLl5LoOkFUTJB8S2Fx9
OIEguE1ZyfArQHRtZ68Dmx2TvWHT7T5/uzYlZD3hSnrdj+98U2ApDd1Mbua5Y2Nf
Gw9GHaT7td/gVi2R1nW3zJRSlSa0fc7Axji2T06UFhE9H6E0j440Xhk+M2+Gl2uQ
UZ7c2j+W8lIKb6Q2tiQv1+oMPp1cQfPYdEh6CH4zd699anPvpGcZzRRznEX3zIJj
yVQ3Ww6L+NF3Qx8q0Mdo3tCnj3J/H9GuzZ42FI2gAQjPe7cQtzyAN8DNkL52a5Yg
Q75jn+Pbu7fUP/dTzgwRTuwCW+72FPbGOScYjkGUWWbF4TTx93MjuFd/blWmD+iJ
SmRz7WeVlDAuJUJ3M7dnpKw3YjJ5FsFxSD/OOhobuMYN/ATje2t30M4imRlLwxzE
dokgxx6qS+p8fZUL95Sc5Mi1bkxKmBbA4PKtyKAyci//QSrpU2Qhbyp96AFHrIHp
lATXebkGQXUuwPe9y9iTr/V5l1Vmhscs8qzz4HjcTEa6D0XtH3Idh5LWT/tEsNaO
bAM9fm6TARA4w5x1e+PtJiTMZFRZlqVfuWBnr78Tn99mVeFmQMRpM7UyePqG+2/u
dWmDPZ07tr6ORn3xCNvULhz9GQjr7AULSJimVG/mzp1ecm+C1RnqbNSNU6UXCwuD
CbWvMhjhR4kyi7BuCsvJOKxuotdx9snx1L6tNj7JzSTWAK24H9Scg/82wLakrXFj
TYNA1t8jCJEWi9ZDqA9eVygl8m2XxQrXuOF2MaQ0d1bQVwM/73HdyP013Fzuw3TB
nuZSDLHKDjaX4CHVt0jy39t830qPf5z5inCo8MDJrfqY73q9flLvOsRRYgjbsjVy
9jZyBMU0ukfKjS9Y9745/E4vSL7ejMZiUDQIPjbpxAyN5QKKWQ2/kIcVLt4vTZoW
wUiTefXHLjRJK9VfshaevP5rtoq9YQo4clWKSmk8z8k4KwaUKA27AJChsalynIJ6
aam+gaPF2qzcjbfvh7XjBjNj95w9i+kqSq1FiyyuGqWU8s1Pi7wFaMciE84wT06/
naAA+J0LFb8xYfxq9Ig4LYPnTUrXxfMuD5Ma/zQ32Xy63T6/eRzMvX55QfJOdMuM
U9tLXEMo05CBJD7/niyWtnllLzovdC4RG468/AiHEitOToGhcSIIFvL1YX7DhXFH
tW0nAdJ+0apsS7Vjo80BjgAy0wUdA5311H4KiekVGba58I33MSpdraYw8KR8Isn7
aaixXpTBHN53vugRxMt1ie5qD5yghHolUkvk5kbls4RS8t4DUaROzgQCiD9hA+cd
cmO+QiF37hUQR+Urim54+QZ+CT8gD93sNC/FjTb+1SsYUiCQo+HeIDMBlGqurRC8
2PqCXjB3r+bPa2TiG4yD4sHu8txQgalnmIrBOASQaGIqmEZaPTGUkmvFlFxnvPLv
36h9HmOZwCGTtRv4st3wMWfcWNQSYLG1V+RgOpu/cygd92aa1RFJJ3WLM8qIpGyc
MZewWSJnOuuuUnKx6g2gXFKXH78cadZPo0I5+FKZiyESgbwqGS9svEaHyEomhZzE
jb6R1jWvoRrI/zsO4rk/q4iOod9Y+C2ugUwIB34Lt0T39SojcAlqe6P9//aaM8TH
V+JlCGJ2cKQJ5xI5mR4UfCXeJtz7cw16KMbvnbxZtE2RHLeEqpLI6NSJrU9+PVYY
pqMEVCnMIFbYrqikkVnO4GYu4BDmxfmfH2lR9VOJdlz10BN0xxgEwcjrq7wjXvDM
aanPjfd9fZZdYAnNhnuyb9cPloNPM/Ap3b/9qRhT8BfUU2QZz2YKTBhZ49hKgmcW
vCN+jR3e+hqjsqKAOMWZx6/9zUezt0CfamYJ4dYsRWt0VXGQo4RiFIdWo5r1Nr7h
fjorZDIh/rJV7JtWrnxMlfx1ABTytaaByc7Gel3B8XBZ4AvqUrJzq2LUC6zWq6jl
zNIrOtStbtN7EDPF8XblsD2Ma6Mbzb2wY8LJqmNK2XUvcfxL2LaZvv/4TU+XjMSj
wX06XglN3ybfgBThV25663eQt4YHzgC83Rd8XATMhAnKQ6kMwKYMEnMJLlZrePTU
GXb/SYrQ6/IklRFkvX6RZzify1tCmNA+4ZA+gUWKbSRT7rGaRqorMFcPUWHiXpuy
1RVrnGtleErzMhpi04hV5ZVHHkp9ELC4oxSfXU54Ap8rMQ79GQV+u2xN034p8ZHU
ykbA8IEG3l6MGMWmyb9vVzCw+G4QImN0bbU/G7MvJrelZfr9L9kQDSGWF8VZF6/R
U2TleeGbPPAam3C2KSEvtzf38R5FvVzpfGUV23M/GnFvxds602aBudEYHqwLolzK
X8rZBzEkPMpGUPTSeEY/89ZgXr/AB5FBc4VwplQ4N+lKFc/K2EEqRYRtn64v4L2b
J43GItN3pL/LnQm5NVml0YUdXZKQ3F7SttGK6d9Co8SfVI9+g+U9fPSEPP7fUL/P
6F9VN5a8pkzrfM1i2zu1a0oQLo0DCyrpzs5o4PaR6nnY0Q1rFC3lEGfLwJclhqXb
nsZM96VzWoKS8/++JLEMmeDXkWpPAsmUjuduwTh05bIP85qbPLZU9inhqdjzUcHJ
43JReMQd9mxvwchcVi48d1uqIcKXeVLKX+pM/AZHid2Bqi/3tm9iLzn2X38ZCKWn
aIitZgSnRJyjDi/U+EB4H9oqwlrKiIiiVjyptcV1NgqhBRUJUtLMYrf4nTVMk5uI
tsOVp1CmzxOGiFuriUCJ2PaIh/IVpVfIUhofwUDWClg1IyBkWkuNoxu2Yc2mw7wh
/Of888YuT/e2R4uUojfG2MurKPd/ABm04jFI25ka2hWuUmdE2geAznyP4QyPtdgx
32KHG8z4ChyapWZ8WVXKGLZjC3R79GapVbE65RWf4iErw9GflGZIyROWkl+6d0X2
Rre+Apj3cVFdVh0VxdbV63aCgFq7evWCor3EzZxOpbLeZWW98HDz8TmiD0fBt7bg
feZIkSpZ9RJJTgEHi2l06t+WY2c/n06rbFUo9eJK4AG0UVKaE0tyJHabybRuof+L
jDC147i+HgYJxQDmqwZBKx+2PGIk0/FewMiOEgVfXrseJUJm2WWJKfXNm/FK51Yy
8pr8FEYNZ4wxsCSkH93NGz4h7RDqqLc+2US32fcc/AfXKyzsOhSLtZoa7WBl2g5F
UiESVmAD/y1ygdK719xMxDGN+OEk7R6baMor6QCRVj6UVoJ2BBP/0FzKiLhbfA4Z
sRo6o/gqpTbMFv3+zj1Gwn+pRAjcdugGoxhqtnJd9MO6IY3V/UZgGtxql/mOnMKq
1RYD67TfSlMQeGdefhaFkqunFc5LF5Dn8KI9chPKkmWovt/qzvDVAw2cXbNKTdzN
BEt6p+FOaMMHS+FxhIBZ34IKek15uha3roien53u453soubnwAdHjD9b990SO8fY
MI7pAJtQ9FI6vr9UsIIr3M8HNI8QJde+Bo65m7AUVeqWU9dZWEVlCuFZ3VXqL0h1
KddeYJS3e94QPewMCfzqFADehps/JA/O2bV2x2/thDYCfNqmaRfLXkLAX1mSYQLj
BfAuLalEeQzDlXZHrOvpF8vN2yhHltlZUPA0hsd5azSLygUWA6pLbWAfY7ZAIHtI
bB6xvdvqEAA4Aeqq5LO1evKiZDKGmam8UZQnk/cLBYpDS2X3m2eem9PMuEjuZ+Ff
a4GvXB4GUwJqTpSyStVL0W0xBx/wNzhsfoybgoC0+lNDeTStAU6L8T6d/3Ib6mHW
qS8tmgk4MnclhglchS3sroF26WVHZdcQkz7NNgMYf2N3Ln7VwHX089EC9ITOx77S
rdUd/I58pTZ0CabsHHXXvxTPYLBOJ7iQOjg4rAg+DhjiwwoXteZj7Z3smeXv6chi
+AIkFJCfBIxaw5MbQkGOuMkdKcsHkpS4EptUzOLG4L5L1GpQCV31LHIXa7erLBCK
4I9fYoQ/4KL4q//JEIA0X+YUybQILwcs++30V6KcoW/7KYxlT/WNR0rctVwS4PQT
VwHfuQbHZYy4JmpOp9zxNR+81hKGSJVS2RZGp0a8Ztezh3agxnY5moU8783soq8o
APfxTjVL3E+AxsOWrIC7U82Ld/3fupUXeWP6t7UNtWz7KWzObiSOWy2TmaqcjqPA
9BltZ3zt1xNmhIS5DoK8gxl0peqYPL0ZVePrPZxEFp66GvBYC7EYS1OhY1Jpt68L
iVwzUsoRJ2Iq1ytRwBEOQyqzRoPFYqdF+1XWSXHtFyKuKExQ7tMy64VfMx3bXhhV
lTOQ9IJg0+Nop7n6idt+QYBPaSWy97Y9z5gfLevunmQranJxn9Zn97dBgRZLJV4+
2R2U5Nlki+OelwVmHQXb1LpKGpUaHFiUnRmakDdFwJmWDrQeA3VOOZiVye7CqeKx
6IxKExt/pU64c91V5mtaffMrqiNvvkHYmfFCyJUn9XBUjBH+LCWrIq8kkdADHUoh
p+nxcaCUmXEpnqaurb6GXE7aFAaKezUkConMX2CodrMU1IU1nN7dD9VXHnEChaNA
iDr2Fc/4Js6/9p2mrizYcXw/dXSbDlzoP/ChihABHz7XoJtUos6bAFzO5/tNMtBU
tsEARA2vmrqwk+0uyN1WeZoU1d0cr0nwLYzKGl9P4dghuk69mo4y0P4lz+H7Xh9S
reU1ZtMUbGKmDFuku/LSBUgLGz8ffRCxq3Av2RwHFovZnqvOjhMLcTpxOsUliwle
l9A4sGKxyjVHqXa0l2SwgeKcjBd6Q/Lz9g9j0I7TR38s0QPwd7P+BO/uhwjIiIVj
G6YLLprFu53hq+OSCfkZ312JoMTRogsDR/PTwUTO9r2i5IXNqjpLR45lRL9NEuXD
rTqBRdwToQx+r4AqbbDtI3JG7yhrKh7lsdmSxKYwbmsWSQA+qpDPzFqI7Z7ByjRk
5+ZcvUL8iyNWQsq6lLCudksluPE1ifRjsmcD3oPIFRlwCR3N+it423JNWdamYP6e
lTFCzDE1tw2X3fR324AL/c9KZ2XEE3nlUupxrSmSgYoArTv3wqc9pJs+QjtMIcdX
ynu0eChL6UahduJHZ63kWZpJORi5Cx9yBoiAoXdISZFeqtOtxkWSxlFB8zgjKcaw
ssJbQcpRmGC3TTMl3+USTV1dZabmu29hQdV6ZGGmkFNamuMTkYuqVWsy1IP0pK73
n4seSUQ6r8/uT7are87Fqw/W6mtTjVvJl1R4r+ahZjnyl0hchr6Ul7E7dm+TDlcm
h0GVqHWhxi1TPOpnGYqQ7EPa26HDY1hCiQZrrvei1E4GUGECIkhUHUJOZNGQ8g98
caEH0JMk26tyOur2eXmFNZA0UX079M9QdTGwRohL0cOHB+J3AxVx10mQbbXRrRkg
0GAxhVuXQ/q1XnweYbslvUjksugZ/Xt3z5xmRfufG78CV2Lc2AHcfVwrv8p0nflL
8espaXxajLKYvgzqC7o5p1eS9DIUZT9c/+vRs01m6VpiZXwDPugyqGtHAHfMK9M3
2m7rHufOrsBu6Ap/mYUD2hfMtK4eJ5v7K/cFUtY/7eKRpsdpqbve8gZarr9ZVgvJ
f3ty4H8+RSA9VHR/Su2eX9fLe3Y+sXDbQc4P7yoXGrtSp4D1s0xB9C7nAuyXYi6z
QUTfPEzHCojaEcJihg8HueBri8IMm905O4lZaMPhyS50vBbXrh2b9j00d/PHqDov
JX9bc1rCUbX5n+CgpZrJphYQDZlcCxrBCpfUZHiTogGknOx+8Xoxy3UIg4Lw+HdG
3cKQ/+IHVGdpxJi+oHHThhSOE5KfIGKPV+Ng2I2Q9zOTbx8rw9jTgA9SptqCFLhR
5/ja3f6/gbhbKLlce3sZTlH1kqnZrelD83w9BKyTUjqUwV0/M48zks6lQvtq44lo
4jrPOdSLsq0NfE/VfT+8B2tFuSv6IvHFH8b+azAowse94QtFTdV5k7L6/DkTZdmU
j+4FNL5IIzbBXr/HptGokVRwiUNAYqXXUKAxLEN/szlWip8Pwb8kfn3q7lB5tBgp
Bg3YiAi6RKC12MmZ993bfvFFY+3CFTOJ0oPQH/YSyYOYAbToGFF9iu7P+ROUbQXT
8oscMVNaK0wqcva9fzK4FhSggIZ/X5bIo4VkihSAcQuIg3Djy9niuZAgJA6mYhhA
GY6zy2aftu2Gtc62ueoa5eETpafZ7hP5d0wApIOFjluqwxu0eZND5OoAUznr8Oh3
CAuZpnjcL7rYjM2vg+qXmAyLU6RhTbZFYvd7DDN5Lt4RyPA+FbSlNnCdb5WZ5fIl
S8Lj3TiFS9PfaTNM/DvoU7iSpZW+x8i9LN/5+j1eiIjGVn8/Yu/5YriLWJ65NrDq
gJPB49IxSGRrcdb3wwEVlkuLcQeCK3tOH6DCRdZLbvMSQMOw34dJHS+FxyQT6MPC
OO7CgSTyUzHEwi+nKiEdg1CwrDPvhsli2Sej0Ch5M97W7DtB5fypTQtJ6h2CINRb
NE6nmj7RzFEDRfwKP8Dt6TxWqgDnsQsSne3B/Y1mhMuHGqhfmIczBcnf4ZwR+gSK
dZKkHY2dpkC/KQdY30fM8ELKgrSIruV6MZT/Xx4Lq9Ks80A1ZtuWnHHlHC5YTJLq
udRapSyrWcKf77W4kEZBNSIwVBmolyXeugjltkR/1ZSexmfvuR1xU8sR3CmNRtOL
Z23KmLb8cxsY6jEH4JmR0n/c/pBxYKmnQMSxHN8iofeX7QL11BpuRAlZxGNob+PY
rcgUQMozthcAPTFqJ6lo2p06PvyvnGIsL4Ii0QJS7NDCZpAnc2Q37YXMPxfJGoim
aU+L/FVYR7wlMYAmN+ndybBsmmwI0Tdm9PJP/A2YzmaJqPlpPlWkXrrEe9ZII0RL
mQFLvDZpkjxG+iYGTSuQfAPQ+21QSC4gCKvDw12gB4VFjtSH/SgyKEDrPnft01re
B7G9tn4M/MI4j1ZLHiQ/hFzh94N20K7dxHCEUfxpfnvdHZxKoHKCycnY4f5Dv1Uu
hcdRNq7EW8/ObDns4qZ3fRc0UIv0H/eyeAaR9+xYKFl0QPpoeQo3Cw10lJM+Gr8C
Z/pEs5jIPkicFfCGeK+MrR7AfiohaLFbt48EAogzvYY5kYj7sHe6QJcdP/Nf5YL+
ftjdBA7ob4jtPQiMhhWStNSqAaPhdGPPy7HqIopt5FyQ0fpiwgEKBYG5+v44dRH4
4BKFCIyHGofwa5KmqjbRwdEWT7x6GnG8+h4dwy/v/fmbXU5WFD5qlVBE/WGYnzyv
SGZaXChwP55o331sCfsPdb0R201mnemhrmm4j2uX503LDpjF4WMvGjdF/MuLPayr
mo5knQ1C+4h+iDiQxTe3GRrrYnzyEo1ov7GYEcPA4hB0zWifxniOD2E3qNXGaYJS
D1/hHfV00TB9nhWV36TFkPIB5Q8x+2yqHU2mb5fJm38efTRjmU3sfIRr/DhaMNnR
qr+yUCNbM9z1tWbeyUW4HsNFbjZIp8wGXJwjjZi/UoMTGoMUELUVwZrnzZsaWJYi
eyjqCkhShgXKNLD95Lh+2N/xAZPfgbpkO1UjXnILY2177rHVkJ/vro4JpymrNq+1
9+BWU3OJF5EHHlKhJdIIDpxdcmg65AxKGYT8ERjpyRHDZJz6veN8IetIUCPP2mKd
+/yW9xHd1Kk0EWKfl/6UIS877NLQ2mAQRotB2BKpAIIIGodaWZ2BOlHLwMKBvCss
+a3JivhMrPFNd0bo37w1AiuOui9ImCOTlXD7LTpFJVZXJi3hVm7YaWMNgUKylQi/
Pr96tLUaiPH6pDmd1M+YaewW7AGnIe1Vl8Z92CJHlJZM4xi0at7udJ2GuxT9kK19
AduhDfRW6V1mNRu5FbbrO05N/wGzcU29yj/Yiwv5BL/q9T/5EJQA9mTOi3Vchs6j
XhS+kHoEMqxbaoMynqO3DiQMbTcQmkOsRGNsoquaJHCTuddBKhZ6YQcW+O5AUXid
mD6ctINY6QFtNR7juSvx+lN8WZ7v7xcwyoAjWOXniQMeIVcYaDxFpZPj8OQbY45v
q9HH3bn5d6OMoU8q03AtcmY4k6TWnTVYL1yWYh+6IvWLDGGhUL3A0GW6Qkdt2KZM
synocSl/QfGfOrWsqR1WrxJlcrR41vCGHeXqD5WuTsJpmm3WL2/QiEUNphsIgomp
uo660oKxhhTFdvkfOm/SoogbfIMpUnbydxS/oe7SlRNCWDQM0KU2hs9n2bN0lSwd
NqgvDbNO/rD0rHSYVeVlYsZVsu7SkFPTcdJM1rVTrMlpnw1KQTnGK/VsS4WAhiQV
RJzbwR9XUH1SxykcKJTAx93Q3uw1spKipwEtNzlCAEeSU7QWP2Maiq+X9deZEPNY
smKdTapGWahOe1YwPgOwx4n9A+Q2QixSTzZBQXlXhEeoSwltSsTfoL3WMlVTRibh
aK5tr9TVM4aVrRqDOejziYltwsnEL60HdQvxeqZTRw0nEwCm3NT0ubEkaOa0Vghg
UsoR1mx1UjuOOPeKed2S0Ca09saLNZ09z9kpTAjNYqAxybqgQCCyr2fUSoXBKoj9
s4qbZTn34NwE0ZHgqHZPS2ZVYAjz/E1TKBGRdYrpraK/KhDnPFlzdb0iegXzr12F
2a1iAIcQwc8zVbn6+bWnPlVnWsfsyvOBNjqL9TS64oP+mNql6VJdyWC6lL1GXXAc
JvcCY85TyaDh9fKFokQaU0AuD94jNfedf/De1WCSLA3bCEElJ9TlecAqqYZhYoCL
yNy34H2MJNp3ySNwDWW1eizoGsr0IL1reELYg6mAAkTiYk02Z8zdN24/EU0zujxX
65E5MkSAaV1jKCX+lKUWfevKJ6k8Asp6Cg/TvsAhofGNoa4eAhEy4qbZaUzhoiBp
8OiiNAYw4MgHeCn4Y2tnOUhqlCc1YeZyKsY2+/ee8GrCJKUH4qSS/VmEOOPkPxFM
9/c8U3aM2UMy/BJY71aqit8fI8yiygktS4IxRn/CS7jT+3ffRIdvYMoLALbjK3Om
FM19bawGrAi5Xqs/87H70subsL1wyUIynklsTj7SAW5mim5j4ppGne0VIER6xKNU
d6F1g2iLOGoOpCse6h2JOt55aqiQ1TqlYByxNwxo+PH9EmtYjLpjfoqm4UNpx7on
zIDrlCAF2on4hBfOKKwyPN84u+4ntfDGLpVZyy8AvxKqa2R3Arvh5RGrPT7a+Vlt
IDfae6dtRthL679nFbvecRI8fBT2iT2ixnWY03Q98My0tT39J5DRq2yscqFBRhbj
00c5/tI3ujQeCnONDegYVk9uNE4IEMIH/3r7yD435kP7Tb1W1Fu5Y3ZqZoMlBvS2
dOhn20ifIpXBAirRsF7V+T4+RQy+NIyMQfZ9fCyz2Sb+2fllaaWArlA8U4vWQAjI
0B7qaCJtQkIdIDEPB3tNZzft25Ow6BjyyZj/lmHKrpREanqPBK5sOzhs5Pz/SU3v
yOrZbH6t7+3Z5QTa2atYs1uhTFNoXN2H8X9llljV5zi9wRsT46QH7ov7hZ9aOqZn
tty5zw/RyDUM6RGZJaYydTV5odkCXyQYR/TZME2MC1KAkqco4okO6AxldpVQKmph
LecEMGxifGactsxdf5sU2LiGDv9JexOtU0A6JgKepduEyp7ahsFCxQjYrRix68M0
Y537GQ4u6Oq0ytndG86WmIlZi840LTGuWVcKxQbjGzcRUstN1EJ6CHfqtTglSO2L
FAevEZXnJttAKX0n6BurIXs7k69yDwB4grSMiDqOmA8CY7LEcMf+m+Fu/pR8RYkK
mn4spmvsTBvyVFMg9iPbXHhxrSglANI0BmUcA5Q7qx4TW53rW2UazUbyY9U2hRX2
rO0AC69Uho0uti0+Xm0YD/Hv6sIaMqvAZStU7oNbTND5a6eZpFOJjyYhUf+JXp+j
rcbjG5Upp4pzpjTWcezEaDg1tPW7zvdrJvcIzmAECKur4VcLX/jnpUh3z0tuO1E9
2JhaKTX7Kgi6O6Nf1sFHT7rajkbnfKm776gndxk3dw3xvYHT7u8H3A8nl+ma8m9v
0Kj6J69Mo1n2NllkhYjMSAauxtnLODQmcKTaS09aDJvBKhFMWRUWtwXZZB+krEEL
iopqJ6l4YVsCjZub2ItAR9PyKrcAmWCQ5nf54iePkJ4kughbRz2Ap2xOUQ+/8EOa
ES++pas53nyYscF2SmKNah2t5r9Mf2mN4FpA9ykgW+OLWA/ExTgp4hRdb20DrIa5
TWvaCvV+ejiRaVXRecr6nYtaAmWzMlBD9BgnOcnDAmW0uf28swnuMb4XnM9AfNBL
YzgkY7i9k0i6NGuGlF/B1LxtweeNQXQJek6aJJqisw/G1oI/PHItIj6iXgNiMB4n
R1+DpK+4tw3fs6sEGqNgUV4wdqz8kPUi/i0AA+4aw9z1HuI5SOVQm2R7WSVZejHw
7C9ClDclkADyMbpR8VtQ7SKIWJIc23S4SC2+ucpqAEb6G5Vk9zLxKBlf+7wEm9iN
mgJELtLvD7YrcIrb4N7LEo3p52KeVD2tXB5l9nGwAaPgEOhtKRNR6VCora5SM+aK
t10g6TgABLxut36lXQ2ee/17dWOHwQc+TSQIaRCseQWYAMCvkkXNzdHWw6i0Zllw
F8sG2+PHM3nNegtLBr3dXTP45hOOzDAJIdCKj1Azn1WTCVaBEj4NPmg41duiASys
H9OKnstFAGIXn3GwjO7DNPC/Rk3M966Gyf5bbj2SW3aHHGbOmnjWONcalsctqDcH
X2OI/vbqFZP/D9aeIkMo5e4+v2rLAcqeZ7knds2t0Mj4NIzgb0wTK4PYX3TXrswy
70fCk05lw3M27Dpx7sP9Up04fq/0hspaQCwMfCPq5YVVMvlWYUhYilNCONBoaK/P
1S1qIqPidiJ0w0LGpkbgswoHZoHq+/7Tvzu30XTui3364XTmzumrn/z8cTjPFxkN
tguzO841+uPGB7/HJcbPuFF24Yd5lQtMRu+5KIVTlUX9GPt1QbuFbgopgYOewm1p
IimZRH8n/1LDVuhfM1/w6lalQNyc10WyLNP7mq7dlZWZitxK0125yQD4ovRNmPIm
V0a4Ig9GSlj8DAd+i/rH0d7jn7Fbs1jXRiPSCHi1FelSXEAMvy97+v7zp2826CRE
vA89ZPwJJmIESyuX9CP95BX+UsGM0KSxmfg06yj3pjH6olKiFqzlln+94da5pxbE
lH6fpCslcEdfKPVx6TD3X0wMjSWla5TyzMDaWH+Nds3lqeYQOP+68LsstyI8U9om
owmeBMnlaIYvxllANUt3id7UQ/n07iY603kQosvinFWAKc7sr8pX/sglrKYywXji
xwQLI/P1o5t5KnBR9bE4wYYA62d5UiXTtIv2GYPXmsxPhLn70qFQKYi4mHvHS2Wd
dlcI+0NJFGu+lqUZdaiR5jtag/bb315HLKOGndjpwmCMDzN2LEBJYMuYSxTa9qq1
+bawgKeMMkem2pH3QBU2Ov05j3kqOlL10btXZ3PmzcJn5kxf4UzOPPCqElVi7AUF
mkekHUvqyyV6pkNKsU7n7mDhyUA3Pv3j/AFwyQ7ynP6YRcFPb7+zoNbHw7M21ECs
XQY36xo4TTfHiBIoO0yS50ERvctQsJsF+aaWRa5cE1FsuEpypVAM/thA6voV5m8R
nUuL/tjy10Z6sZ+i75i/JCht8XemKV/mc7s4fpHBALNkAJ1LcDtRKhnbsjI/5Cc0
sFiWnA1YFPoTolYq6+4RusvCaPem6ZY7YDDItayDiZ1S9s5Q84h4Pa8TZdXn95z+
bWbWubbmc4cO7D67WS2GBX/2QOTYv7d62nWW/4N2roF80X09RjNAYmo5oNdBqBXL
lHx0oASxMEkWMMSCAbHYOEWtNKqwvsx1PMm1/K/xIMKd32iFjlAIPM4OY+ZarRAv
KRHnAzc/bhZFuYcAl2c+21QLgERb2zGAbeNnzA55TvRwFXxAkkr2sEvPpkG09XjB
1+cvJcYkU4maNkQtyMMplZQQEEDoYjW5l4e0hJtwosiADAISy68N7y1SRB44AILz
qhW1RcwXmSe/4E4CsyjbVq4+k0wd+WzgjWqo0hQNduamuluXcyAy2Xuy9CjhquAT
HWBJXzqPOr9ruR9RiLUL1dm40ZERqwaDqR8uHTSZdVmYaTDFdJZR/cN5G6d5/+U6
dCkBKYSPpED48J3xm3DWFOVaxwgNOgvnVeNEa/Vcz6lcSUsG5JM7dy9CAYfhvE4q
tQgf1OQDidr4rz/ajeNeD2iOZW84LJR23MaruFCR2IWIIya6wJvWJhqTl+KNF0Xj
t4vvyNf29WPscgWqF/HrtDzqXsU5tJg15LiTw7NLvdKBcR+S3DEvtAXdn5mLdu96
Nqk3VLW2r2S9FsvqcEaXoilbhlvibScojT2vb9+4lWfF4VJNuJo0A+Wj+hih7Niz
brEWFaUg0XzsKZPODzWzg7CSZ98gUuYrxhOzh/rAfJ3JpvIoq9eWT+WCnwDtQTIK
hPFZ3Eu3shd7y9h5oy9IYWL7mHwGtv4IzapW1DyjCQdz4Uzrx9ZmytPGxqDJUBBw
QR0tfOXHfUaDgstgyvbKNXl+IcwEJb6PI4U/lPUCWBXUFXcMXoG3aNrn+blXS24b
6cQBqYD4Ty0HeFQe2HAfaWPJX57NXeDPBftC4vxDltWknOlw4O6+NpvIvJGreBaz
wkJRei06vD45kjveW8jheYDYK5kZ00NaAdUZK3K9B/5wq/R9gcXlVzwtAW9vST3v
UeQMO8ucsNmnP/nor2gZZ2CxQM1Syp04o44CETFuHxq1vkKtXZLQ4gWRYi8f5f+n
kr86798cZPsat7kcUTX8FJbRZ3PFOipAHdHQ1+oNGhlMvXFOa27s+cV4FR+aWgWj
imO4hAacCF9IV/axeHNdU/ZffRty8Wja61HLxmOXEGF+Jvya+fZtE0ErH4GUWgFR
KjPbHozL8uBvwBwcploIEK6Amt0DaRGT8rSu/mvb57DdKq9D7mpdjBfrytC4TlN6
wdWzVysY/K9KTgvah//Z5t64e1ZWh515MBnkorR70WttXxv58CMeH6PaLlhT/bZI
zwI3Fi20CsfxKcSiqC9rPzq/cwBdPqGjYMggeIj8zfH4CsB3yuoKvHbuv24LCQRw
KiE3ExXmqi6yGoYkCVeb+yzAXGU3/b4upPqq9OQ7BI1ufMJdQH60LHC4ZVoKLWAR
q0WyGoZFsc4aGTv684eemrtUOYvzE9+hK/wWDEq7i4qzlRspmBNN+cZ9W80/4RNz
WEV4DlB+xC87AA+Rttk52MnpTQImxzM4vSs/Wv1xVBPsG9OrYcZAg3NXv/+CyJSK
OQPdLCRMoz+EqxfbvdLDqQe0JGPD4lsVjQdwKUcrATbgw5Kz6zt0oliMmXnp1OIK
2dwBVMSMXTbaknm5QMt2xtxklFmxXXPZkUoJvBs5Cw3rq2SgdEs9+l6iDaNg7II7
oUTyBEfBHX2afwHh0se2xWQ4hM8K6W+d1W9fUXucMm1yFiOIRY4W80eRxxoohnQi
JwWa37kV49RRn04TyqeKP8zJItqMW0rnxRvm1WNQfl2y/BGKabL0SaLg+lBwHwQ3
t4nJnZGwer9uwB5rTK7H5Rd7eGRmXvodbAEk7xE1qsaM2KEriMoCR6Zq0ouOxuvF
xsu+iELkv+FD3Tl4rXPxkiY+V8+6g9PSLzXlBDWYblqaGdu3S0atWWi+ws3uKPzQ
E+UAcSqRi3cqla/eCPXy+ru0890OLBM+uhWOZhVDYRlsAnlht9AI0xW+hC/1pc7N
s7A6IjgdRsxyN4rqIroqtGHnIipyWme28ZKXLLpYeDJdGYu8wRw60SBLFteWUAy1
UhzmLCN00TZ08Zdwmbqcf8RKAwZ3DWqMuBUqyS4vw/k/keiXiu/6/YFIHbUg8hjb
KNXQaNlE87kn/uu6PPF5mlOVH1ZDDaaU1ZlzJnFtdqp7nn689HXoOjijKm9FIjj4
j7HdByOeAJCyoDxagFsolsGqepNYQwxc/ZtCnA32PS00qMo6C0ecgLOTIVZrwg+7
rwz3oJdwkR98MTk137yyf3hFhRq0N1V6E00W13ZLIVrOdgHMlxMJ7TAGo05FBZFM
dVNKfJVnWBX0ijrBaaf3ipZv3JPNiDxZ/oWVbQWpFcHBIDwoeIY2q6/2qBMklLyX
wXNHQmqDE72P6vyiYdjBu2laIKOEJ5QDtLVE57BQKIqjDPQyQN0C/rpWM8tykxk8
rg8J/mZr3/BSWSCXj9GuEK5tceC13UgOkDqQBhJCbQKme3NVnI197IYwh4P+sZLn
NcDflN17ZIMRXY4R4N2ZrR42O7UjkfOi1Rk194cb66ylkoPLp5QdTdS2z9HluXhe
T28AA+ZEqrE22TxOxrRlxo02j8x3hY2L57v3FQf+5OLvX7sLjlNNZnkiGHCgePOK
CMuISB/SIBJ02IVV05AmYKfqBUqXnLyx3Gj3lH0p6q0H9i8pmyE68GHmFvRnuhij
nbWXAPPvSugEvt0ymnGThK3/zWGLaXoyy/BHmerOLIHr4FuJCUh1VtH69+/BYpir
6XgpfqBo2Oj+RclRu0GpnfozlQNx4sxrwvFYuhZ0SuA4wGsWFySTeTzQRCrr6jJv
abk9lw/SDsqdpt9l5+frwRmorkLuLLTjCX1gEzs84hdGb6qExNGNElPU6FGCz9Jx
EeeDGr3gjwmIx4oM9iY5rDCK5yQObakLHPwWLF5XYKTaYZiJgBfo7gu0DPmhDFI2
USOOc8E6DtnxtfUq+lmbUHhA+xzahFnLqRzlTikCV0q4lJ1w8loQEIv/ncK3JuBC
REKi/k8kSbLk/jelagsB7q/QCXm+A0D1nLf38WnT8CskjfBIQ8CfoO1cHzt9iQpK
dqDgJisVTa6LniXQ7YbD4BXXkdi2vn1QgMS9xpR79bf6gNPj61y89gSm7ksQXSZU
4Y1q+En+uoRPruky93Dr8EWpqloNGhJeYdUsI5a35Frd9uhPilA5BmJGyoi1YJtE
TvoTF25HBnO1nB6HnsQ/EFR/r3CclbLZT2p9OGX3bMIMsjUKyP9TJ9gW/nUTDwt2
HvpQDh8RyA/2KScYHpK7mKKRvCUeZr8Z9uqEu/zR+Vbu2Qd0wYho+ukkuRJEOi+X
nQrFPVFmh6KPk7P/RR4MDVKhH/VBINKFHquq1NWcjOL+zNfTqs9SkPEBLGGA4fAy
TKuopQcmW/IVL6A/4Rzafig++tQ5o/P8PKDUeTJbFOJnCFiKw4ORQdqCTfAAbN0e
IuJwUIZwy9eK7pCFROeYbhh+LsPtNPxunU4YHnbrJUkACzz26TUUCBdXRmcLsZRN
EJ4pMe12SFHicKAqx4ZgebpOoYXBqqrG3ij73qsW90zrjUKCh5vIF8yNxpjdC6FN
cwADs9tJcQVfQYPig1Y8PxbvmxOniqcNSgg7ELrq0pMcXON3/dMf1US5NTcXVW42
zftY0THv5oYLGCPHxkFMMy4e3e3VOAI1Gnm0AR5QWuMlq/D7x5swsBFoc5sZT5Ah
n1VlU67k32oasn0l8znwNJN3SHCzChO7OdJA/ZojWzzxGlYh9mA5fVLGFL9nfHRC
0rf3T5+VYXLQqaSvndMoVFXueHJurfR1ewWDQdNar91iJsSwZJqPH/RWOxP+EXbf
JM3RNFML+xfM3i3LAlbL82lapHwRQtzJfUsNeJIBMDupuL0ilJi2i6u8leyHaUWN
5bTF9VMDMr+CvLuVNiaydW82NPUiCD/yDpu/4/0VFxErd0n0m/YX8ypstCu9pcGt
+g3ueBFxNfxtQMfcrMDqfHmEQuidZ3SYwSXHpQWNjZDwkbEK7Cs8WXSXZg6h39A9
AWQy3UmQpl+a2k2Rrus0DiUb/mULSxxcBOkJgPixLUeu3rNOkBwppB8bmpyygtOU
m3iY456zyYkkN7HFeBdwQ7ZvJF2DLRY0F142zGvOkeUrIpDDVhibfglDk6PIJ0TX
eSJrWxXuOh8DjcRm292ttlotXj+IIZbEDPXMGhp1eoZC1yBzvd6MOYrVIQIHZ+ix
HzhMaMs52PhsuiLxXqQu5mbUS5wRetLK21En7KC6lY2uIw9FWWaU4R+RzDx8j8i7
HLXU/v1PISHwmK9uvEyq6GgL9ve3z+PhUVugZp9fwaP5FpBZebZADUX3w+usgRjD
VYi2qLa+9/iw+PNttYH/+7py0s6heGAnRuJKEIV3xMtF0bERod6TMG9YXtWRiw8R
9MZ9yGfmNNb59nJNWfq9KdbchVNEhwKK3J1VPZhyKbRDVQPVTskYaBnOBzgkuV8A
tyi3qmzgxi/ooR/5BPJfdS22mNTd9RApWskXWYLnbYBmyZtli7XAY0BCSiY11KdB
pi+A5AfS4vNdcYqkLiPPupjoqZSf4aEWdE/5fcQ4xgV7UQPXg5c/8fE8oTV0Gcne
F6VSg264hOAPtjTfYhwZvsnZidINi9qA355iYEOF9kGNIzrIWmhifllj6UEweEnb
dg4Kn8qUnVGNCtHQ8U5HozK5idpHVBBVYkqZJzLUkWPlPn9qDBID1Fov/nxR9iOy
EcyBb7B3FId3/kScfNlXNmsuBi1/M004KwzUgMSEO14mmoOb5wVb5bqUYTO3Pjl7
BCWv4Ka81yfFn0/FnBAqHMdBrBNM9hErFLqH+3RoBkNKP5XHpeZKzSAZOQov5Cyq
pOu4K4yVu8fD9PVEkX8yKWDprqQCpgHwx+gYd/l/CG28aUKNPjY3aEkAdYndIC4t
HQ/zmjeZfrU7tzl94sRcFfsRMSZhea+09SCpr5ZXWFM3cHa59fzx5bs6VGPEpsHC
/n5Jl11L5sY4nCMx2I0ZGePICgMOgkKOTmyZbnA24cBj6M5l3UnMSX+6axgcr2xq
U2Z9ubP5TbZ8Jb8/MQ6Ar2RiPXwqri7D96f3+TCEqXDjWdVvZ0PjwRARLKrhNJOE
atnZnX06rytkyC+umgtL7btz+mB4krgm64K8dJV/qf/ENyNaGUKROX2VXDqplMHU
kD/CLwAoUYRFHJZomShGgkV1Gsl2itS6/tdNGDTZqrpl8STzDLdBwnxZ2NLBAcmf
6j1s6IcfcziRTIg6rVpr/X1nY4dvWlEGlLBSstGx2cCzeUcRAq5Lkw37D4U8y6aW
SWXseaGvVE6VdlEKf5pTlxjDwBLkam++NLAhxIwAuKfS3WyD8bfO01d16qfqUD6N
kbDFUXHJOg6S5pVAI7YSTlrN0APiE6lKh8hQzorZllw65B1bBr2EtshYVqx7Mexf
xXm8BAPGouUql6OQyXbYisqpmmwEXpD1xPcLuowLfymkWNeWdQsKHP6zYlqGUYwf
0tWcLrVo4Y1S+/FFN7+cP7+OCNsRSzc8LoFK1CSu2qoJE3lf3lMH5AAbfjdDHof1
60N/40vXDoC3fEDz08BMDrJFiPKnX4KcWj6jCMNINWP5tF2kcMECg5kwEEV1YtnJ
PfsAODVTNRGthZIzARwrAxLunajw1EGigN+SW1hUSzUcX+VaNU6cvaZ7FA62C6Dh
i7vqbAWO8S7TNk/ZS0WtBQi3AxC1TOrpZzxYSUMK9Xf3TGnw7ZSa1OqnYvygyEZ5
mYkJWXf2kfemaXyZPiBBQP2oUgAx0vBZfvYV/WbwyRvexjpV3zfEeXK2II+kyEO6
IB7VQlDfQLmO2AujwN8ppmuQ6RW0jd/CdzkQJg8qUv2SzdhUQKPicX42OnY51fRI
o6mEoHA0fluv8wjgaQJ4GqbzM74y+1vmWYunaHo31g89Ei6StcLO7dNebaiSQ0PL
5DX6voSxvXpwwMb8u/md0n2QD3z7ZI/A6/O0k4nD9LUApvrdgldXah6TMABMGT7i
UghSUCRaszEwvj65Wy3R2QnSzlV5qyg2Taw+fDyUzV3rKxaKUTYyoDXRKz6DeQQs
6J2aF7gpTGGD9DFljpcAsJ+yLjB4P7tp20S6bPGnxWUdSKfJ5IJBgYHegumSSguw
Yr2gdjeU7DfOnj8WscC0WETlbZKigdeSaoz3Bkoim0VItgHfzLeaYx5YWthrEtX9
u06w7YFn6MiJ6Hl4wL1ymyp9rTsohVE0rWJp3nsiEtJX/xqQwhlFVrjdURSnRTOf
aWMY1XPucodcL+yhzgtme3pW+4l0AayO+FQTBkAt+Hjryb47z8TlQg1HPTfG0QB9
ZnzuFIDvDjJ0f3bnCMRM81yaXRCdEhl296Hlv2phZ300iPSQLCrv2WsuTkKD/tMM
PqcKcpwj2dECiaRjRiNXTCC01Cs281NZ8T9qSd6gDciR+KizvmFnPbekJG3nAaKg
lXnqZ04GukENYIeqvKaunw0xTZvR8/J/LZA4OrkdOX6O5JAzQ9an9hIR4OmoKq3c
AptzsOXEY5h8BtKcKRKJeKw+iww55t+QuVtrYqfXorausuNQ0z7hpCqDu0YpelNo
PeF9HCPF+52XYdlIQyMyVvAcoSWJd4+fkVRURpcy6WrW1ae/IwHvFuJn+zvlucEa
TAoE2jFXsyJLBuJRiuUWHNiN10QQ9Oa8vAfBbtd6GPvWYIFKVzQbNxr7NWK+1G1p
qbgna8aQ0BCpron7ZUq+UBBYX+4nr73MoNtpxa2b2kxltNGVi1ycI73CVRWpJe3A
g0bo2Ves3v6Jn1FFqctY93l2aASlZQADOSeQ/aBCuaePAPNGwWAc1Hr1u4ogMcq3
nC1wru0gI6ypc30cPrqd9X8/WTdDmCbO4oqfybAyM6doOw9qoqqO+zvuKHM69+t9
DJXQAxhrot4MFDAcqnHs4Bvk0c73LfHiTeECQtoNoXtdGGAgh91sIuSh7m5qckFz
lHiDaSlCD+n3hpN/IHtR5Cwk+Kwp/E1gcXHUYmSTtbqQreF66uRKDjo6FiTOFpGH
7ySVUhwekuLOJrQgrwRNx5hVmVvqAwLsiZS/GGSpn1ZsAxSsp2S0y0pTnBkDrtuS
JgnAdDxhRAmYnmQJXKli3PHJsjQ0sBgm0zSRl5EzdsMCTALyZhXytRFhkSA3uJI7
v3wBhlXA7vlUWDwwOjuEVYhcHh2xOdcYQThdktSMAgHdkM78KVPK1kNawgtBtoh1
CP9K6xyGjcOdHP8au24yzpG6NdzJdULD8mnDzBxmyfLoLO0JW4YACht4ISIiK8XR
n26p++2UQpXb1NbMHAh+XRSlPqBrrziaabZehJ9EzBnjmolPv/R6jnOF6T+Z8Gp5
PF/MCY9++HXX/F5k0OuHZqQ+FmED8dI+4Yd9HVV0A+7W5T9mWI+XxSgMnInf43oe
HKTZg7oHb0W5bdnJXs3XLlBw3gfFDy08kIOcLyKXs0CKmMxTy+h2bRard6pItmBb
wRyKiIE0j7oa6LCUfwDRpYCWYXPTLN5aNlITfiWMXNXNO/RoPZX8srst+xq76xxF
s2vjdHwFHuQzpb1kkXH8nkJP/rNqpzXlpkoHYvbT1kD4NhkMvgVBcZr9/bhlODPq
nm3IeYGCrqJWWZP+Rn+2kCKodRVbmBJcW9w+5sqYMw3M5OJxp6N1KzVDsuKK+x8G
bmWajpsgyNhkEJXQu3B7esWE5ifvEMjB4DwRArQMNIjfCIo1EobBFZSPjqIPzavh
6i/PNcro0hiZLlLl4TJheUy3U3o9R5mXjliEtHikRrH0DEK3RO0EFPoly90JwBHa
W7/iryr6h4qEOMrZiCtT+bxRqkVZ+VEnoMfzdccOWFtri5oGwmHeforxIP6yhfdP
97VIWgKNT9TRc8qAmj68AvRT3xs2ciMNUaUvTocCrcI0fpftvvadLdXlvcFJjd+d
0QPgP/dOBtq2UGD2YytsSPdyhT3hIBHzrQwCfNug3QAcx6Us5cDmDO6/LXC6lmI5
c/jRPUvrdW9E9bDPBH6Q+3pXeEbU8+59rFxrNhz7M/HeWfJ6m0W/rNlc6R428tJE
rH+9UFsv7+mqFFA2cxXzg9aAChTXGAFk1++fDfvc0pl4hFHQ6r73wgQj12V9h5A+
4wCZd9kb5y2e3T7fGQmlIN77BlZC1Xnzehb9YBbLoVfs/6/T+/3nF7LWYPKnIWTO
+JXg4fAY9A5y1R4fagm9P2KtQs/aBW25+LmZA9jN6QYKb49FMVY574YJKhhsqa+Y
ztWWqlhyAVVCkYdeYGXVXMVZySkVHU3Kjo2OKibkgrvmZ3weqMzNGV4dZ+O8CYxy
c10FaDlLcC4prYX5AfXgYcdyo+eqIORaesEkVb6JAISYtAT6i/xO7UqtDSJukdNa
plohSw1lvRcgzs3JVH01qLZssrtKw/RVQ6TGJoVoEDFFzZMhX2s9xH9gBydYyE+K
DJKIkxfP/qgv09t2KS6AO80AW/6q+loi4/Ku7hpoWKwErVPFMVlRQwxk7ZZu0Bpe
7BASnS351a1pAlv07CoMqywhhfZhdYpBz54qKRD4RtanaAIAtWd4azj9sMIw+yti
LIBibUJQIh9yz/LdXPN1v5sSi2x/s1A+Q+goN82Tygi3G4iF0KbL28YvxTgi5RtH
W5J950/QcLYKROIvDaTSZrlqmthzptasChr+07WZZFP6Onu7rmxjv6+v8Pc7w0y0
z2kjoS4QoQUba2xRM/EJmTlDXC0ZHB+l6s9eEq2Wj8K5NpxPuRE9AdXuNscKAhFe
7P2WdXCuPqDBdLaeyi9vUmyIvwyu8OyxyA6r76KkrWZYvkKMdClEgYegGToImzv6
G0FFtD3v/ronIyavfLNxWbZ7kbgvje8Uro9xcw2pS81v7J2chRPirDPtQ+s50Je5
FSwVVcmxNdK8ici/0o/g3WceyoG1Pj1DWswxOGwOfrUlf+Q6KCXMuvtEVABVe3Oj
d2fP0YZ0uwb+3A2L7z4+wFfa89ArKQDL1SSBJIKWWPwFwe+VjvAMkdshq2CUZDtg
of5+EJEOI6pRA2RPO8NCAWVkPLAPw7bbW5ucc2BcXrItHu+t1ejD2PpNJ4Mc00jK
IRe9YCqyIT3uPbUMJv/qx7q82MgVq++HqM/LcvzcZ8WdyMtB/JA+tqIUzk6Dt3WC
kR48FcFoEb9mCqfm18rUAM4R2ccMOhyUa8XHLFrSVAa+2dOoeXIYRuB7NBGvvnos
p16iZwGYpNInJzpfHXqMH/f/7RTW2wBjz+T92j/KMQbw9R9Zz4yAPZMlcSA24Lxx
UXLHsu+sjZ5liMsqhENg53C9bE6zuRFJqvaKRrygGhnIMsCFyDBbeiaiJLsb9kOQ
jIqh8qfr4VR++XvBI4KSCPa9ryMt1Zf8nZq41CQOdU6jRERnBkOW6qrL5G5H8vSb
qKVH6ij9izSxHhEfEz8MeiQwXD/iz665yGBhy6A9hUqLrV1BfL8DuqRMKlG8uNPv
Wtc3CP5tXoCQK7TEnKxYakreDKEMhppP6JFzz9OOMCAkcEDMCJy+3LT+VdzkfhmI
u+YdLmAaj8uXRhGS+JXoIZ9Xtn5ChR8dHBe4X/vIhuZdMl9sevB8qfHjqo+iaR3x
VN9G1b8mvWf//kgyYApWAxuPIZXGuJ1sBWhjU6GQS5Y50K5lzx5Xa4igOvd0On5/
SG7QxgEsfa9fQZ3cLOpZyX4F8bSlbclZkdVubZb8Q5qpcC09B9Sos4MsG/7Bw9Ok
KFLdHkrZ9O1jdvoxH4F1i1/IBHrDCty9t5m337Pn+pEp62a+K7idrPwvaT6MiNzR
9euAgW59676E9FZN6mNTLXeBSPpbYccGbnTvVCpBVfBv/41OdlSQsX/dp8gmzPRS
mbacgWRADgtgs+8IBr8TwzIR1qZzhpIHoA6pYQ7Vnvox7LhyJr6WrlyRinR8xwvz
WjRWxWbezRMiJryiyhSY9m61YvwzzxWkMwWy0eOhDtBhgFq/X5VyA9QNxhAScVZy
6jGSkJKhGThOyFmcTmoIkhqHMWJ6q5Tr+cLBMFth04L6Qpb95KLUhmUC+6O5aEG6
AqUNi9j3IRqvijEq+zMw69fdI5R+zttulfc7G6R9ygSAbsDNhOj7keSm6BvoMJGe
5vHa/EMZo+tNayOPH1Ar/TgA9XnX5X108EFSTJj7WPiza9mD+FX+dhMwPkpN7t2J
s+4cGVWP7UdOmMW9LXwnM0K57jkY2u455Hk2iuWTzX2FaAgEHHtt9hOE5tVE9oaZ
asJnV9JKpfEcsdPvBcM9rxjmPHMenwxUe9fJxQDEt8gBMLJD0ozMC3Qy7u9Xw6uN
i2VrE+e/Rv1tGbpLoehYddpl5nITgrpcaB9TUHmsyRUqhJn7TPF/CGA771wYbSTn
+cIXcR7jPPa+VRBdVL/zg47Tc/MPmC5WdhQ2g+hTKeKG28fQc0NFxhEkrNk7PqKs
680hNh53i26MJSWucrxMKo01gppTC1t2iJBVEXx3d16SnGrV/RZwKJ5HSXg9oZp4
VM7KBjBfSOhMm7eEx37mDPgsCIDMlMganfW42di55EelBDjI26QUOxFvWJpFxT2O
Z5qOQ84x8Q5ghsGjpiM/g+78B6EmInvLiBhVI2eW+qBkkmz57OjcmlVl4bFs3KLS
a7dq2gLZB6BLdnUtLgUamTo/0wnnEatXRczt42itc8dqut4H8eaG3s7PePHxZAgW
IvvtoL3hQvbigxS4dt9WN+G359aVy38Wi/fsomOYsWYOzyC7q55qifaXNXqzGLho
+5XEhqAGEfviob9bLJg85l/7b7VQbZZzHyrafmafDsIzL8ZIynjbn1iBUneKgbqK
8awN2uBz2/fcsMuRlbZF3H0R+p8L5s3PUvmmTP8hYctxQyYCMln68gT7H8iG93tr
7vJbgE3m26iuQ3vBRuaDPmhLp60yCAf7ha7VFxwmXOY9vx6unehPqjBIw5ZwblMo
IJ0E/1lD/EFYjlDowedg1+WqSFhEGZ5b/yAUMAob1du+DVZVdQDJUNw/1D6j+QRb
ZrzLIARYpfBe88LoInXIX1IG9vdWVjYicE+m5XXNv8K0ygKkdo0wUIqrsHLJfCUx
8z3LLUppbL6YsrAt7qn4IxGkfpCRDbWYWb+gs0M5R4d9q1fDqXRDUUOX5RHMd23n
5LYFeaH8cLCgofWgdhuSXBVs+Ti1TGmbny7vnvnnZS2gk4FdJnejGbHDIQH+cO/A
xvwOtSq1thyf9CG0SNoGwRO6pVGLB0QWnQo90HF7qSsgPW1OHvM9qd9jSq0tmXtM
Z2ANBxShNDTXI6ahFQFJ+x8kfL+4VXUddqD5lokjL7pX1bfY/FUfNLqkW6UOziuO
T4rHfr1wuIeCTjOgB2L5L4yLehe2xn8ozqFFfv/CP5KRy8DfaEatVu8SH3QD/zpo
2PITd8wXNpXfayIV7ikXJxBATSVYcUFoGfV1FPBP/G7BaQz2grDCoWSVyUVgn2zC
SWSTY+nWNjUfHD1y1VCpX8f+Qc/HCqZ2NaTs/xMQ+Gpf+L+P7eua37/jvV3QuxsR
mrPjKJFaA22uRznfi3oim3QrYqhiKiI7IMR0ADcB2A99A6lMqyZhTvfEeApVUzC4
TYLCAiR1+Vcb5cKfiRwuVQAzx+DB2MLt2kfBiVPQQLPwTn4SLcB7fF4ZI1oGtYGu
0qiZy4UyEyMkLfEvFeWNMgHn74qOKZsm8aoaJhGTAXNfOHlHcpYxVKLzG20ze2uM
AvlODvL+LdJCWHCivypme/9z/36mVaoLbVyzBNLS3oYKNeskRHI51iDElFj8etPu
redJTfyp0hEEFpq1jjFFw1sjISU6t2ALkZrLaV0SQvCQfWJn4jFNMoU3L1ctpHQM
qS/hgWpKl4opBkKbR9H/hkH0FUiv5wiYCXuvantDW/+yN74DNZu+qSj8aZX+GeTy
gawMD7Hj0Ya3PLJ5uI9VgZ2h7oOjHkLzwm8IxnAHHCVTnI9S3KAhy3BiljYegvfY
YI0b3r7+42wfBgeG5KqCfeqCd4PiYUdIekcCNvfm8mO5v8rQcRJVFM8IXH6ZNawA
z3dHh4AQH1sIAdH46bAKZmKxMYOswrbd4P9c7yVncd4RMQRz10jiaQu+uPVUJ9jX
YSYiVN+qMw3pmoNDKM99V0XAVvNmDZjkfZsh77Ov1pMq1R5emwvUNF2vII2y9l20
lkkbM7D4whYLbUUeUiwduyvI+0F2ZKdQuQOo93dIMSN32+CP1b4bcq69Uy7KvFBG
5yxVjNk9vsIT6ecW4creu4NoB2hA6hE0ctuwHsqZdzDgoD8tK9tmGfv3g78KhEbM
k90NIRgqiq0kA+lDVWRY8YubnrVnODFCYkEILTUzcyDgw/DidR6zsrUUry2zNhmv
5OJj9qx2CXXsBnoSTi4FZjy2K4v3eXDx0y8UVCRarewh38PlI9yysIbjAxuiz+6R
Aqasqup785YotZ4DceUiuEUEqD3U/NcCCsnaLuYaQh7GR4pPc58isOfv5/PSrC63
S1SgyBZDIixIpdaw7A1LS5g4q1IpDlANMrLvYCKOou1HYjSR5X1IMFNjvB8GyQXr
2k5muoUPjCER0l7R1lU3KHaoXj9qReKe1Ny83QATQrk+tblOliz+8FQ4UlLZoO1P
PWVxc4dH9AzSEWoO7KtUX95rSQPo9PRDpayltrMrXIRUdiq43CfNMMVFqdeGuPjK
pNKJ4/uLp/jE8ygKbFSCFFcc1j5ur1yD7Feh8+9sAT+9ui0HJvcFJcXcIqiSl6mc
lSWQXj9yJuEREwIxdviGYo7nST1ZfOsuAs6R0jxC7WTQk7IAu5/6CHfHeI7x3+YD
gDwsbNI/glrzp0dNLAULMTRjHAOGMIXZhKpLjyUtSdJ0RKcatmoP2UtO5Ca4Y1R4
qq8d0PC5s6HBN1CXulLAk0L/R7fCZjcdjUa4xJngDLb7oj0XDKuKIBSbNGIo6DY4
/BS09zc35+R0tsYJfUxaohq3nUC5B+CA+I89lKGhxlof/M70ymagIAa8smdb0+Ry
f1tcmCGI4bXzdaFV/GPO+M0o1akWRIuktZm5UEihQYtUA5BjcbLDg7tY4SLw8k1r
FCYqdUqc9dFndzVkBkYTdNfuErBuJ7RHXJB5koKCfdcpoShtlJaAaxtM+UOUSRXR
KrJxT5gtBmJq7BDZxSqlVtU7c5aPtRhLjWn1ucS79ZZqSJe+PKTHdqsjQ/cr47AP
dDJQ4kb2xtB8y7MWgm6BbO3oeb6qHgX3FOoeceG0ALzeMILjLiX2o+61qetAKjsB
cVj7YEwi6nnsyq5C+JOpSq7Cvt5ALEH6WQJf1NN0/e09hLfutLiDP8lOL8pjmfr3
9uoi/FQt2dxNsJAx9KifMRY++j8X6Bc/2Q4U/DKREk++Y8yRROCvuwCjLRVZ2cW0
38TwIVgXk+mS0Bs380JoDEih9Ju9cbAnFRv6FrDYG2L3XYmTl4twVa4fmZfW3seV
8keSb2WQP+MNSLx3S2pROQUytFaJcNQQeFDRgt5h0h+/aeAAz728G1JiQKDIqos4
N6wlXCd8Ba8PkbjIMPZFIpCXELHDTfLbxqOpN5iTNZXgxOhBIGjcmHVLupgm0/jp
RFwUTEI9u5dKUUcRVeaXeFxjo+EHFs+A0UihZ4pCx7Zyao5Y7Z0VWxEkBuA+6rfa
VfT3Ccj7bz9QNdpDUfJjNQwU1r4pwq0r+PhK6/bBrP/zg4llGXq1qmLfLgVerE26
/eZng2qaJKn0FbHXQudf5GKtRlAA7OyBEXtpgAF4gYh1GO61YH/wdWlXEoJFQaYw
dzRua4jPFpKZFFMeSjhpAY6EFIist5qnwbaBV/ZZvjXqh4tV/jM9JZiRcqzaVlna
WNh0ZDiNcQ6Y1G0pQ/vt5Xsckr5ULv5GJ9xEWEvwHvxslx7q1EXYmXiUsBEz3zCN
6+05PBluwOnptZlxINyzm1GCw4H3OOoKY81M9vkpl2B873vR8sMpihGue8g6dXOb
zP4Egki88xqsFcKykFT8s73dv/wud8nE3+I0/8di0orQZcAQ6jRH7ZtBwhUVKRWA
hjW+/jZGNvroUK9WvC8JbBiQjjTxMpmZKxQjH/IQychcLiXXmsJVT9LjmTIA+Hxd
VQRzkE0qn2qLCMvrXylwnZigC7e5x1N8fAGVdiO3MZcrX8jYPD56b+S5dmwXTTLr
BsWfOaH9sTz5I6wAOjiYNljPlBMk7ilhI+ZhpcWPHNJmbjEW3fytryegGT4xQ1PA
pgEa9/6q/rmfKad4gFGYg1iyVg7pPtKT9uklbIxcNWOduTbf1gLB2ykqrRyP6ALS
k5nbsiky6HSwqMO/6cKSad0O1uCGdshzXwgtAUAljm8PUekIbvMF67mAA7kpzeG+
Pbxhuqk1NK3Qa7PdxkaYvnAtiCyFeCbBQ6Dwjlj4dOOO6lnehTA2Xa9Oosly7Gzy
B2dKW88bWqcEA8FjC0fyXpDHlpaBqGUlb1DmF8/4A549PNsp5rK98zkIPwscuJA7
LskjkjO5LCSuvHwKLX3hlT8IT3I2AMbaHo32fXzTIrpq/ceVh9uvUH6XwTFLowkq
2u1jBTLOZ7HlRfvxm1olixHxY6QCdYDqCN8WLdWJoNTW0OunUkqKSVY2MaeXSB6r
G4OHiL0m+LuVbw2WVZX2gysr617GWeVNZdCTzLKzaR+3yFZjPhRUrh0rfHMhIWB5
BsBUFM3hOWdMTIcpJgzeGLCsgsSoq2PGmiiLO8VJsR21o8/PsKla0iCxjekfRvV4
7hm4JlGv+2Re8Qt/4+y9ufXdkNFJKYF/HzxeYgiMlBlVINlUpzjIWu8bIuhT3jde
sgycyQE0S/03X6UiPAOkaNXagJ0ECPMHZT6apWdlE+XaIGN3K84RpMQ/i4dbOnh0
9moA9Dk9bC4++dk4nivRv62buTR1fasb3u1HIqtd3TfALWAThR7rbBPJuOKYIwdv
Fjskxq4laPLHzN3K/aw8E2HS3SsdYUcj5b1Elwl19PLB++J/LpddY1gLedThM9Yg
0gyso9E5bQRm/DKiSFjDLVx7wfaFnDJJb3U/0FLBPZvbSqlmBwkFXPMyDFvKDncS
0I22QulUcAj+9b0ZIVxuWhenQ8HiTFn0oQOI/7KLPTrHJDvEWfm9b32tkl633QVq
uHyxt9Oy09ZPn89RbOjy7OR0orNTCTNAU01O/3JBHsYHe4yq+45EAULAiI/cNsdg
dwsvkbga3Z72Gn1tD5uReH82ZC4ZFPAdjPdcXR3StFJbiIA4f66KLOaf++VSwddi
uN5iZXRJyTEkH6TtCve2IO9OBe/43vOSj+RhC3X3le9mF/8AlVIQrj+OiUIvslCl
mcmC/yPfwT6tXeo77XWCxaIzpsGm+kmXNGoc9ZW0clMllnHH159JKYAIFxQ+jK6B
N7Oj0HU/bLcVJVF+UT9kL4moXvQSk3GILMwoKwxSSwpTwbb+J4xXaGxF3qIxZ+3e
AUPYOp8aq2ntAB9eGZefxYbngYoSAPVKpWYlEpFD8mq87zlXnXvO0CJd7YxL6oDu
9fK35EAhkRZa78yV64gWao2HH0s4g20brkkfqTwYSCRQ4X7eUUT6ZgQZeKjraTO5
MqH5zBS0AkP4md3hfyb/VR9vspuSPyhAV3YVge2dSazAa3KS/WiM/MdeNRTsLOBg
Io4dxN8yVLOdo/li/UjiPZh4EHGqkR9Z4uVn25q0f7Bsg9j15f128gzXTp2NAbLl
J29qmgI2GnD7wZxp7mrS6uXnI2poXmklaA6572SyEZ/xARKScEUyu41XtzmS0vTZ
9d9PKkDcsROJyLD548FYAKaX+vQqaQjacc5wFHNQ3XQw8QTSiW9fzIHWQ2qdSPPS
ekWtmpFHg3bQ3zF61NWl9E5BLYlEWaZCyu6CZBMcKMYsjoqsrGtlBK0PUcJJaQq8
lxuvlmFQXdQ/Z+SwzHD0re/DSWFuspywFnw7zX/z70Y5MZm8nuGo0jBhNaQTFc+B
7WGQIayJIboYryuq/CK1Vq/PvKxUA9TsZdoKMovnd0x90rURZjh9FaHLh3cEw3ro
BCByw/Lle6X2bZSXLwCzq4CeiQffWrt8plNn5bhzOjMpf+6vrWkutJgz4udjS6c0
CbhZUVuCzl22+RiH8MdHmCg+s96vsB7xTcv/+WFBitWFaTI6DXj6vnO77riWWZgf
2qF0QlZVeodzPc4KooQ27sVfAYFAsQeWQqSqxY4BWxfkV60CNY27mM+Oi8JBKX/g
fWIb2RRqtIuiqGNhqLkfHXy9lTLAuhdZnRcXg3DIEzl2Plu1860E1bUaSVD/4LDG
2nQiZYqH+s8PCI7rmDESOhFmC1yu9eARm3aWHwUwApunP5IUK4WR9TgWu+896wvl
1J3W1dxAgqddNA9ASdd2qpQ6ssHTQQAkrFsKXtdJXHEOa2RZ/TJm6Ir75YbauXLQ
UO955BrI7eQgojTVOWMlB78JfbWpaJK4lU7HKjHfK/nZFHXg+/sI6M+eubbYxFex
uc0NrNNNqDV2eQPy21VEtMj1vToPXNayLaVUxwCiw6V0PVkoLF0uGsQRo1PIKYhA
Cc0X9481psc5EAV485cAs8Vtwp6GD478/vFwQmdDwJrxniMukBnqQKmZIJyu1EUW
XIXoh26Uljw7wLCjGHTUKm66DZpZYvUz/MJjDFbLhbHNo40EmpcSrJBsOMHrQrY1
9oQEw7PjLLtVdDtosFYXiUesMgWevI8t7e/NPtbn1uD7Z4flbXVVdnu9hhMoO09P
xv1Vdb41NjO3TOf89KoDgMxFylchxow0jvvetwiR/bf8dmKoLrSEckU0pbjxDDnq
bM/q0XPtQ0AboIR+lzjL203RDWlUwPkUiF4TSr3iQACVcsNLhZmn8lNO5MQn+jOC
aJ6zXrxrkDTG5I+86+VasedNsM9uDfYEjw/y8SdT7eGwxnIRl3oupzXf2EGir5rM
q4bf5/GjZVIQFxhLpcrFA2tZ3Q2cjIHhpHshNfM4FVZ9I/OsWwywv7r+455Tvfw5
5Is7zDVGvgEH/D1RxIwKJO2UswUZU0QGcVRpHkC2yU23QW80V5EhXT+buWuTjr6i
uG71UkAJthEBiaERNlBQMb/ArQT+ctYrU2LQnFdxNiwHp33foI/eza9Y4iFV5mL9
PFeZDE1SqMK+wF5OwVf3Os/HxABxy6sLmSA75wq7+6fKkfd7nAMFcDVSl1FeOWN3
hzDrq7Vp4Z+okxD/CfcH+TWF7b5QPNT8X+cq9Pzl2bpj4GSOs/JQNVBqkHcvAKFD
/ZTgtYfNFjq8HfQjzaVVgAG3ZPn7JzDXM1sM0uOlH2gXo7paQU5bEPeEaM5ebLor
p45d/NBzgcfytQ5sn2GxmuR7jU5uBYt/HaXtGHWStQU1fKwOezHLTekx64zX6yL9
PCj3U8WtJj4EGld74V0GN8FORV75pKd7k421LnyKW8kMQq1TW3uVFIdyrZmecFpf
jPee5j+SGNe/6EFVvLOUQTk/zzCQKdaVGmvlk1YYemXSEQVDt7+6yKf4RGc3zzxw
+rbmstjw6o0z65Q0KmaP59aKR8AIzHQ+o1Q094v0GnVdrzGcwDHdE39djbprMI7Y
Mk0Qo06FzI/1Tast6HJ5jizZN8rrMYhArZK0igj7m3A0ArAjayBBgcueD9CfFy/L
D3Ma2IYUZtWHRBc5m/cRmUXHWJdnPcn/QVJ6cE8AjhlOCmXCt6ieOpG63/3+Y5gq
E87EhobSsruZ1KdiJEnVkZ/oWMTBahsOLxJwBElNlNMUnJZBpTYY9NwS5/HRmNEW
I3OSs73vZCXMo1L149uKTq36lllUUhdZeWR+pwfJ3VbLFQHcgD3xxGby6qzTOcgQ
9jVmymEPr0rpBiaIKTwrMYR1Dh/DSzHVHhXpwPsOeYyHvZMeM/K1+g84aM/mqAUL
7LFdCG1/pXCT3TvKx+sBkoV2JZg8PtAirQ7M493cYslPHdAxEixim/iT10t+tqvg
CSIf0dFpt+4DZDKyA3ISOqzIHYjkNzsC7VfpnAhHfcymudx0JnC/dBXECBBfOjeG
gWv6KW5/gqxh1pgPAnrY4kh188Sjbz3YpMLWhVOzkUE64ec4fD1KPYmHn60DZ2/y
VxmExdfjerTk2Vdr+XE1zMJE9IEjFIwqTTvcmxcQC/d3gCNxS20DbcElUMm3P4Kp
dXUuP6R0iqotwQFYf12mxeXsKWeKmM8hJ0+4o90S3LOqpdapJ0YHEBs1rhII8sHX
4iSkm0qL9UGGeJchHeL023+aA3ptvzgcV1ljamJJaVG3bQUzLca0PZ0+FxJYoUO9
lmBCBPhpSHvk8TXEKUxUwUChF+1+bWVKiT/El9emou6lkhJlsffKONhuYz/Roe/i
rkSvOlvfbWn72eKNDu/1ziRzIuGokwz36rneR0i8W8h+kzuvU2dGL3WfXgNjOaIq
zgFo8MMuDGk7sYOVhFbR3eRElOmcolWkBreaxX4WQCjs2WWH7GkRWrg9Nf7wSI/Z
uKERuEcygLcei2mDURk5LdrsUhCfUHdnj5kXdYSWH/CoRSmST6ts0RtGIcw4cJ6o
mM2qQ8jIu8lzjJb9tsaVGkWMkpUrnPjj7rdDCit/ZhQv+Ds85o03vXLa2RDDlHga
/pyb/3c51zFwAUXcjtAKR7+FkNMZSDzIAZiYw+qrew1I/WQY2Bbl8optoAwe38Oa
YX5mLFcRhApjQRZuIuJF8AhGURh9YlgdtgLDc/9vGEEnXa04tJ4tiL8Uz+hdwoJv
+qkZaSaww7oiWvyE17WOEczpho1gC1y2EOZ5LAm4rVmEhesKpqThUNi+f8yPyhvx
hfr8FHVy6kMmS/kEiXvFRYLXGT47QD/kWqxx+BLTeO33TXAYKGW71UYMVnPDaID7
EI6f90/MwSFBPTn3jh+lTS+21rA5tJn2yQ8qk7t4URBzkaMiKu63KtP2SkCF00ZP
JG81mJg1lqPwaOgxyecVGiI7XFS1lBSL5O1uWZvV+V1XcxxXeGBPQV8qXmMm1NZX
xPrJscUJviyRbiJqouS7UB9AjbBzCt/dSnxvJa8Nb1Qj2kA2AKF+anZCkicP3Q/Q
AUua7O+EB7mXPrTG1uUhZ+rwBaN4Sj3Ces/ax4mKweRvrMcvhp3T1mhusGGrEZf5
CDosPzvByjsfRDXJ6k6eUYqJLKLdsqzMgOq19uo1QZakNphIdfRM8a8K0DIqlvSc
38a5SL/EXBYP8IsirTNrXdG02ljP+F7yXXePVAwEnRYF32gCCG6a9Z81B1IVMBWW
O4xmTtq2ExSsNzQWRsChurWq3Z55CUAPzGYtWB/ykb3oDp5a3Gyws8SVdcu9UdMk
h7KfyBS4qla1qNIEXqgGvUqIRi8k+GxvwjCmPJMQ4j4r8dQBZBPdkohERHWK5Uve
S9AngE1YcxNhUx5fCBepczNRngRUi+lNbwM3ApWu//GWkx3fInBER3ecTrbDM/zR
7W69UTBPfAIINyWajPdsiTB93pzuGjVN2IETKbKGqP3doK4uzDAmevF29mdGUfMT
PvyYHRiB05hHwuhKVOShk7DYRw0WVJFKQyocJFeNijUSdTsb5yn8+wMLdKQJTLho
BKHWlucxhispUQWyLXG2Y6CJV/5ezyceu7iaJ4I3BrIWe3BnWUVkOgx66n/Q2XsR
OGYpGOeIaiRfvY7NVcITvD3IKqDpUQ7gCV3IGh9ZJk0gRaqMUQmPe1bIlageiPVD
7Ok9S+Zx+2YWuBB5oQyZMxmJVPt1cZGd83/z2zadQ37ssRf1BdijQtgbPY5d0EUa
fWLJC06pHiM6tdbb6ZDEWfTuJhUsywxRAEw6zicJnpY=
`pragma protect end_protected
