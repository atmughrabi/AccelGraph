// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
iycw8+eA5kkAO04fLiuDYCL39RLYDbbX5c0FKECbNc9LZgbn79AbVHNot4/XysPN
qWPh+fv16DZ0s2t2ROdypnoFTYXm0LHdWNo3TNwUtCF5O1OyYZe93Lw5Mzeo6Z4u
EuZLUsC1yBLKMenFabjaGYomtYK8BfS7NmjSv3ii/7mqq3PC3i3G8w==
//pragma protect end_key_block
//pragma protect digest_block
nFu7rNzKHNyILLMzKhVPXZKQRVk=
//pragma protect end_digest_block
//pragma protect data_block
UWPrUZ3xNJpH9KQ+yM5Vzv/Er9giQCdMfv+38EMp0B1Kp317K8JhGaZMIiv+wPnS
5KRg4uXn//zjbGAfKieTZPUDlSAkzPW7BBZRNtXqwueOE6nSFBc3P93NU9rQgVP2
TNp/GW45FbzlUNb/zvaHMx3joj2BDVp6CyC+NZs3MrOn0VVob3xgi0nehPwp6qPo
V1i6MuISubqF4lTvTagaQy9/YGEAnBA0Hy1ZwkuTZJ1XTViKNjmacPRT3CogCsai
fOWbR4gqfCjtJG6fsjAIp+sDg678k1YOFTlGWCneogT10HKqACq8S6ULk0i9gv+6
VSLteM+HK92/3JqDEQ8A/1G0YsrSlWEjgU4OYtyFMF1b1fzD7yDZmzAijY2jYm7G
/DLi+LqJAWvD/IklTHrVD4PKMimYeZOXRLLHXlIDt1H9uRJGfB2I1yB7pI53DrpI
ghUora8UMnUusmzLft5OPDonyYBeQtFJ7EOxDkBQQqtl8iX2KRObMjB+ovjAwlpV
//dbLatkJtaMJ5QLtZFieM+JMKRDfzzgmcDi/URSHI2DcEhPSEBzu2T3cr/GsxjF
hpZC56r1WDYHisLjPam8YwXOuKnSlc6M0X6y2K9w2Bbt5kSSgVlzp9cQQIkfdIqn
UxJtH9+5I5AZHLVp3MEiglszJtveLml8ZanR9fD00Vt9Tk4fkQlXhiml6LcHmy1m
Yx4Fl01Zz+qIZogswnMz4fUIXsi3CVzugH+XBlcPIXjhvGIBLATiiCbt6yZpXYt2
2YdsjJ0jftSSqdjvOuZI6wP5ks4MUHarvJbOXGjNR90Ww/gyvmzD6vlnzJ6j7HaN
v20UwXRCI8PN8/j95qm2ZPYWFIWTMlZjZATMyD1lJr/jNcfn6KNYc18IaEP6W34S
w2Xu7QDUhYqhEaGNxEV9NEu0TN6xFKVMpFEqR1RuGsWsXbv9sSy00pQAApxoS2+5
lB1ovlx61Zr1Gl8Y3t/N77c72rWMcSNRi4JT0y/hTgWzwq0EfFRneVqWp8ocMzkG
aNrpEDtMHQLKZxriRDu+wVl0urGetiWxfNDeaMx6dSBTxxoaoFShJsijt9H0vmOO
JXh47hOcu3aQsTllaLpJSuehXcd3qMu8bfWh7ixMvYrK8uCULba2JEgqnGvMPhRk
+7Q92a0C8EQaN90lYg103DLrZ+EHBAt3pIWdioKjkxd4br7VRh1yBh8Zp67CFCr2
pi8Ye2tDknPokKgI4FTsMtYROfBhQOTVnbCR1J94XJTqqCQ+SL297X/EC3tmODLZ
u88r+yQzNB1TcepCnC6+CG/MitWjogZYCA3xxGUfV1RN/FdpzTrO5MhIJGJMUNoF
5xVb3knuucdghmnRQrDGN2dRsxA9KYryEMo3d1WHKfQ5VUZKEUKFZzXT6ZCGD+bY
zAj3AbFXu7zra1Wk9BaT+OSk/+9iwpE2xIl/CVbQsuLwekFG3qc9ICKAxUTerHko
mp+a3QsswXoMLLkrYMvwYtFWHndwd0/6ddSLB2OFs+F9nZJ7pw3Ag5TaU9J78Ncy
tOB4fk4UxDRloWF9IuaP0Z7KRcg2gFRODdlS8N6c2w9qX/8DmVIw6W+ECW8ry2Zf
XO0Q9mHv27RgpcKmOWFf5rehPi9yhWXW10v35OEGxv3gjTWuhOiVdeqGV0D4yc6f
Nqcl0MNjl+xIS7de6gScwCpm035s6enHi+H3FBjLRtSfzgAnHzaW7YBaajDMxarE
YqMLqvboygeY9spf/uiDhNAnKHCMdQgScKUGM+8Zhk3Tu6rP00ny9QfWKxzoykl4
zNoQpHrmtVITiaUeegbuHfj7+zgXjzUYHb9C9aVm4wF4VaTWzWX3YO3r/M5+jAV+
NX3V28MZ/ZH3nrrUs530WBlkqSmvNnSfQPTV+0ai8/SgGx4ne3eT7mGR1fd+x5EI
CFtANJOkVQMPtXjPdcvdlUyrsQ1Sggf9dTb4V+vwHH1RK3Dtl92YaBWOxNZ5iXVA
yOM8MxS/xqJj6WJ1q3flE0x7YJ076jt77NRfhJ+iZt7QX2EihGREoCj6W4kLW9D2
c7Jwm0tkpq7FB/A+2n82F4RNVtmc9aH8wJ1iFbgqcG6765ss8WKZ6YhWWT1RbgvT
BdhwKWA7DCAa3n59yWTYdP+oAh06vql0maSAydivg9MdhclBhaT6OPJS3F/5pZxe
w6Ov4LuM5rNaxuQTFN1CIs7kvZDplzaScQl8jXf1VIv21E3gypvyDyFpyDjzNDgV
h1KbX8Jtk8pvXzUmOs+d7OD85xfbdyCnG7F/DQGPIpssAXilXp3Y78JFJfyA/Z7z
lemw7AGKFDpbubgNXFWXx7sv1jgGb4TZjX8NYLA0yyaHgGsVTw1WbitFyXMKmIVK
YnzdRZYKumB+nv/vLLsbP4t7qf/RrjdBFnRMocGsK+pumpwe9JfyNMx588h6/7vA
fxrXQtpwckiiobuBIOMv8WFD2yWZDU6WMY5EIDWNalHdQ85YjLGU67vZwm4MQdeG
HdVa+GvsZbgedN+5xNWY/asFEfcy25mzxVGwZHz7DS+vfHiqYhoJRty5vDHmTAEm
QF32991WS9r6QG7Nd9AmRYLwFFvKeGU0Wca/ddJYq4SrfS2ZXSd+46leLYilRcO6
qGVLmXaH2Ykuk/FiX6pIxfSQ4hK9yZLEH6anbt/hJ8mZ+kINZPvfY4PK6HRDHOgO
q/hVIgPDzBGqR/v7/ubyUe85lW6Ee2ohhYViv6uaNUUJS4Vj77V84zr5kvAcmzl1
dpiyntFMK4ASzE9Rdc3JjxRAbCG8IAzDpfi1bCL61n2bCA2aXOQYdo4d84QvNFNO
ybx4B12NdPElR9S91QBhHLbx46wRoaU+yDGvcUDddVW62X/+Ok4/jDfSDSEa1JVP
bE8QQKTRpgy9pf1Fn8NW4+p3Q8WSz6M+DzaLQYj7fgrNNYG7AVT0mXy/aMYB2Gzj
qB4RPY3qNOq1pBsCYiKGOj8GSyxJbCvADWbGtG881SVvfD3KgUADpB6HPNYJ+pJe
AgxRFb7l0Ph+9GqQ+bps/9wvO1/W4YL0D/BHb+79MTNeGJCjTkLESMxhEDiMuXeN
Rol/w/lQEESbyE7slRn7RY6y5gU5ZXpNzMKMSL8eRD1Z9ayZ4DeHmpoGvW0WfF2D
9mSQ0ljpi2jPTrQ5GqjbAeHADHgRovMaw7lrbm/J6l2O3ECaO3+XOvF2Sq2HxE5O
3dIZS1BUYQQIF5JDuewl7JRvYlgFoABe8t5uMqHAO2krkkTVvMmUoBPk1Uj1LJk1
boZTtJ0m7cuNFTOZ2dARcKLWb5ZaMV7nBoosarxYKDghM9PDHRO0HAN2O2T47sVP
8AbEAx2Q6b9jl9KmWL/mHLb0n7guIM7OjlPlVz4BMTq5I7n1LOxAG2W62D0p2g6D
i52ElCcxZv0E5cLZXE5SKvA/T4N8BAvI3gQzXOQ2xQpl8qz0Y+MsInC0oPctKEfK
ynt25Hr/3OVbDA9U2fOWv82KkBS1UgWrMHAbvburQgGl2NeKcRpuEBkV7uSCgfMy
01LwcPdxmqROHqvNJO7pgZBGoxm96rDuEUxm7ufYziGGM3K63fBRzd2BF8Tzd2bt
x8hnv7SXtCL8y5zo33cOQbb5qgvlk1Zna240ms+G1x2i++HDJKmdd5e3jyBSXD9M
PUGfoWS+QUAfUfVVJfFYC72tipnuw0+HCVy4Mj0sh8roLvLFiOt6ParSReizK6xw
UOJD4DIu9Xxaho+zNEbs+/ZIc9b8lm5rTN1BHQg3MQVXPTHRZ+QgVPPlpMLPCIst
Wjw7Kd+UmzE2PeOV4nes5+nc5W02RMuiAPa9OpEpDbEVgN6/SbJ7HJUBRZSvr1zD
Sjb4D9/kDthg0LatWn2b3Qt466oU/gC9BIuiPTGYjZAUBpSVaGPSBuyzzmnAXBwA
gbWXcqnnY4CHZEYWCPbnD5QMjeLKFRXlBmh3npMJ1k+OECkU/Ny8KWBfO9FfxHeh
vklDfyQdmwpJWPr6oPx/ouwvGJdXvXktTJqyIZihySIa7XpLmtRTd5MJRuwHZu+u
plG2tBCz5Gu5jePtVPxER/WLxgI7BJkVXGLtjn11LdoJe82lqiCtJavijwYbTlex
wRuyEutUWGMsvO1i9zjSdwU1O5U32qkOkav7vGIdi4u5x9Ew5iJUFfPdNvND+j/S
JPZFVxm+NK+MouS+64IiIXgXqw9yulQBhxVT+jf3Di8m12T4rgB8QmFibe22s4jK
/pYxa+9QYWKaJkOw/KbehmWQgEqN6ozovb372STlXPDbb0rJQ965kGEYSe/Jsxu4
G7CWxsqMkniOANywKGy9gto9rR8o0FltFNuDolg0MiYa0+KgAVQ/xJzHq636lFgs
zqT7gCU1QrhOsMvCaUdjAFHrjiq/E0GRI3yPBfiEz3+AC6RXEf6CWmcM17a3l7sp
VPl0GvAZELyAMzdcGtjEYh9I5YheCgR/s4D7PMlY8cd6PCduZ93LUqx6rsvqCDxR
yb2u912x58MsDQhiFlu0BstOf/ymJ8125gEtpAGA0/jiVpKaEjjtF51AXzgZ+aM6
nOCrznhaIsjPaXwBdOhyp+kuWoeMHL/3Ps3hur3Nhl9B8L9hXSw1wibL+gTqgw8V
YnifTR2G8rR8RXHlL42OEsaC6WwcCQf3fi4+o8pEKFokGWmnfWC2S5FtggmJ6E6C
vzKyFYTNteQd+pKhL1yNdySGaoUWQ6+YqpPzNONJYeIlFtM+q935wPteUz3PJsuO
NJrmZXVi5OmmbNpBNnQ+HtkyVNck4Kdqef/fn0ArD8lDGD81456I1ZHmsCp28SO6
wgwDfPU9VqQR3ObOp2bgnjIWpb0ouC/frtB8povRyEIFvoQOVZxO5IQ0rU2KKjWD
oPZv0iC18DfyqI+Li0hKAos1kNdotFVKEzADas5DWDyPv9srub5gf3H9vNipD4cD
lfpZRyhHyCrfQI4m6NV/g8Kzz8e+5TRwaEcpJPj0FkKfuL0KRxZiADMUgJuUmF66
ShVrl1q5lYoBMXf2VSjBIZm6aD6fK5/i1B6AmlxTLKpa84eKT3eEd11wr6XgtXTW
1nxjhzHO9o+i+ZU6UMKQNpVElTeYvXOkBwGDfIHwqIy4TNfk5to0VEQAM72qILrZ
8GGMgNkIW8+Za7+FbUXUk9nBqAtiIHEKh/tB8c6LortGiOUN2y0crqimxQmYXmtD
cDZ/og/TzQiN5d1wyhMyXENxCOvUbs8SaEdKReYYbkwPFF41Tt/tGu12iEAPQhq8
xTdbgQ5muepfe1U5cxBxRYr49q2f7uajWZPVw9IsRWbp+MOz4LqJRJn8IiBWJmL9
F8lxKtrk5Y7haXUH/RON5gYdT9QORYTMYLcCDD10fogY+5pZEkhoG0/P4TkaKhl7
iHivM9J6KZFXjusXOJmYPmSattC6T0nK9BUNFo/Q6KwnrCpONLnmdQ7kmxIcQsc5
aqEawjCuD7uc4vIQ/c1CYsyDUoz/w2cBYfJB4prgpDQEF+3PwsYc4zF9BImqi8VX
vyMlQWTExjJSR0ROoeJexMXnwZ5aNYTM/xNXZmJzpZmaBumPyn2OKsPNvySj7/Fo
RFsvKRMj5k/F/6Di9hOtuyh9MjIqzpDwnDIxlpjl/OLYfDiT10hLxdaWf+rz+Mnn
HZa1sOLMsg3u03ZC+5aOmsi7YZU0BY0zPnLKYrz94rLww+xI66ZuY0RzrVW86juB
nTy6RdUW7MG47GD0ahfTCeCD/PAmnFphn1OjqpIrcl6CMfP79wr+4lfB7gBUgDIG
fwFICs0wXW3sPdeKnEVnuXUS7IJUgvIbNWbRC0FA13IaSg7l2p1ipUBeraziX4L8
tVCwcfj8qPgdnJl1LCM4DBt75C+6M7LXRzj4y+z7PLseKTcuLwii651gKj7RiHyU
tap+bHt4/GzjYBcm0wGNXOM8j+NbJUACLHMwqiLssPq7ku3ki1jFRuWVbvFezNxM
Q3ETjF6FIBPYjLt1QL18pX92lKeeUEO7DN974tpbujz4ewPkenpV3bWUoSGyifBZ
sHIH8L15NtMLm2oA2ISkwmw+h1wqwO+kr/a0RdMSC/i/gVB34Twr2RLKh654x89+
WkEix5RkjchCWxztzOhspQaPPRejuOplSjtrOBbPu8AtI6ZK1L3uQFf7oyZoRk4X
yhF5nqDt5yxSfi4Xl45b84u1rSu3SrFLm1m03fvaFp6DFsL9EbsUDmL8NHVxmPYZ
P/apExzrhPj+KIg+8sozRMD+RJvLwZd8DfP+rArUh+Q5HiwYwdjQTnT3+1MWOAhS
rQ891uLlyeKsfY4/9tyE0Nw1XISy56OfAlvgmnU456tLl0irLIOO6jUt8LhrTTpN
fix0ziJ9S3A93bKv/p5Rl3SCKpN6MeP43ZVZcw06ckOW2k63HUqXvUEACMk/dSTA
6G8O0RMadYlp3ncA1TpHRVVEq4f0XjHRVOxBp0im1jwwTq/YPu7zD0mq8Wlbbw/c
f7Gz4l/Y1HXuWMsVX8Ba+B2LBBb+MrprlQ85Flmzox1i1HvMM/Bmz2PDe/slRMQt
LPz8rLZHxkFDngffH9Re73azIhgejSA+kDh8VEzYJryUXfjN3T3G2eAwvC4mfQKE
RAD+lUFtKJ4BwDtd4BZjbdLILDQOGuWPrVj0oW3w33W0EKxSG+c4Q5o06CCGK0xO
cXinLi6KJoUhLmL/EHKDbnX9G+za1QwXRh2+wXlkJ966Ke1+u11IstqlRnfBugFW
wU1E/lip9H1eZYXq9OGM63S+UNSagewEAD2Uzs2OHMwJwcoS1ZYC0F3ZsglgeQf3
RsbQeKEKaXEKIoEIGeBMXM7wnKsjcXKkTEW8pNzBi88kZc20quPtMWA76voIQXHW
YL+m6RYVmd7lLNzHbpz+6R4OfnaofSIxBkAGeJF+vd/FNXI/YpOtl5S8dvIrkaBo
j2yAa115CWnj+F2iPYDwXhXAsBxAjD32Nx4mEDYUg4T0kyhOOAPal7A42PxZWNoJ
RkwchREHZ4kf+zSVYQykR9Pw3SCntrwHHo4PlJ/THsAkOfpyKORtZ9MTx7z7yRww
B2Svs2f9pJ/Udb94kUImxUAlpJiN/WTOUeuTb3fADkVJp5Hhos70SLdRPRtHrGJ7
mmAVrUUE2dgF7kqnIBA+9v2gb6Q5mTL1Bjnknud4gWIZ4W9JB9kmZqYsaMBtgjmB
i5Y9jeSvMsrg7XskBN0mjHh/qPVtJXK1c65Ti0W3XDxpve0E3kdD24CIEa2KZdSF
gucfbvodikq40tBMetV2SgI+Kv/cAZiUJjnE9FLrWbaCLPTOzVELaekdUvewo125
2Ry7nC7sEpkgKiLIymDYyCjnvwKGwDFMSU61NbIOlA+dDrMLBwO3s2y9ux5wK5s0
y9k52nLBjAf6gGRRKi6I5tghdaquLeq+n/KHEh+8o3qtSLql4UuPlN0O1IVVCMnA
firK8BoQNrTtYJiRNtMWy8bpQ1i7GCIbrDGGFwDmtDw6VoSIIuBaUS8FHmvcnTFE
ZrjrNmODitUTw6pJI1illO3zPfpxKIoO0/YPt9pIblXW1xIjhsNL4YswmfIblEQI
rBjhzHhhW1OCR6TtFgtCOD9lfPDUfMZp0fkWCCnJyCN1e8Z/hEaErX5q8yUZ7ACO
qfb9EZYjjBfAGO93lLAsHqtgSyAl29BQExAFX6ZxpVj0F02U0gwNtHKvUpaC/P6c
xW1Y935JdRC3UuKPEADRDRJjJkXEhyVLEVVcfZhZtjWf8oXwowuYU6EFkGCIEvFa
00FNRL92FuWnjskUnYWOq6dzzu4fPOYYJgpLL/PpZoeukMo5tnFV1e6xfZGjSI+k
fZLiR05i00yLYQndiO1H5pWYT5153RzPaWU1+GdXHToDkqhUWvMnByi5kh79kTv2
E27QDMriGSd4aV2o4DYzOHoVh68XoBzdSJIFhWaF2sWjrgxwDQoKAnGprFGTMXCB
+FK7LXsDLovA5aOFWl24BypafQfQd/BqSLrBf0fNI1ctdgvjv3mVC5GXIV839qJf
oI/RNBTgT5PGIPX7/OXssnnAyt8au5AyoYiFFpuNUnhl5VDIUAxp9teh6ppW2gTB
/sH8B2R3jEa3z4FriaPnG3D5O4mvBl7bEvfCSuvilkDPNonn9OuG1amriYppjfV+
YdG+jehXV0hG7gK3rAmEpahDqCMHC7Z1W0K11oV6Rb6r2zf9HnHCY74EeyNUO/C4
pUF/ZyyVTPEmof2w91FZAEo4KaRa6p/z5veeSWyxVb5x1YedG/CUtUEYG4jAwsdX
qJxzsgumKBSPCHn53v3dA7uJ1eAmvY639EzWyNyr8yrUSBm8fnD78yC5ijjN/VSW
XRkBBU7O2Kx3tWeAodx2aN6Mf1IFtWxAa4/3gVw+UacbWBFjVzfu9KKQR4X6DKj0
FciYhXuQqBsI6f6cnkRs4jqOid5ykNFc5Xm7JkifVFKR9YZyiZYOJjz72/YKuv7K
yd8hjHW3300/njbP5VasCCB34W8HvsbbchG0T057ofF30W5trfvzGXo7s+SYEuiu
ErjWkCpCLfTjwnhDyMkVJ3nPO9b9uU/qcDq7azwXWrvyJEBgIEpo5hIxwR6vACva
XkNeuf4ZLJFOzBRiJHSuppQf31ZpQllxdzpdyY+mdCEryNoVuZEcNkHA/9qG1rTV
Quaq0yENSbQNhljDcANtk8ftwTijeQIsDNwckqbqmHjej7To+cbCGG3rVw1+Wrb4
wwenLeVoFcvg8FxUgF6SiaLmhQskYjJBr9XWGPPuFvRXw2s1C8s3hmrWSm+LZy2l
3ftlC5bnfSlu6Yk1pRDeGJvzDL6FftgDagmNWqrNzsoTu+4r2ODDZMNCQ0uJwpmZ
zN/fPmSr69HQf0rGLh1nUoxoTyJQ+5GpLaoLL2DJYz6mdCUxXdHdq6A2HHyIeYBA
C8ma3OVHXtp/O7pv5yY0SU6NRXbqiZa9SaZ8KhJimZxaB52rpmRW+Fp0YsshWmSr
D/MhlUI3b5P1SxVkhgX3rmjnkK6iUPY1W5nWOQsUIasEHGCZDu8bt8kO+jIsYl3d
YHR9wSLRv/hI0Kb2ApNUpnaiADIhVaJ6IQLmio/uMVjfiCd1ai+MBlTMw34bfD79
Gx9msvloViKXmwLIFoo9oAWpqKtrIqvk6pxEETh6p9UxHhLGO9YGdxdQagKGAo4R
vNJvTpuq0K6yc25xcPuujHSf/RZ3BYnpozzw1/FJMWOcFQOjbvUxrHlHE3Opw6Yd
viXhOGRahD7VF+SiPIRfDvnUNTUCOudAkeJ4x3TSoUe262OLtror6ra5XPczCCB5
iWNsFSvEQFUsdEGGTTHCT6ak2xwhrXHOMIirBTy435ntYDbsywdXU9dEniCHlL7w
mgE2373x+p7Drr2wtUoJPFgZlSjzs6hDwaqQLiP1VHBLvXIlRydx9sLd8IOe2Q6e
WXnk6btCsWwYb6YdIximfyyYeQMJWgIpCChL/xy6LBYLc2Mr1i9Gy8rbwlvX6FUO
Ww/Gb5T+SyTm/DQToSeWqTIrJxBJ7fV8fs/aFJymWa3a1c/tkRUKuWUQK0zvLMIv
XJLdwRUt3Qcc3TrQDF4vNiocKUWPgtLGO9VlH1TBXlCu94/nBQEVni5kba+jZDfQ
sAjvPDBvO755vSQa7TJtms4GE6EkMQZ2hiG3D+pNitfJ/dJXT5QKkOLeKkeITH4A
EnxtDoElbzXM+bnbbdD1kFZXEZwhlBIlaO5xoMlDAiwUu1678Us6priynCAgp3g2
jzg2MUMlAiN4kGMEghqIKcxP+yiQnXkd31pZT3z/sgXVUgW0Nw7vR+2x0o1wX6M/
72iOIE5t6KaaroAxGfW62eJ1C989LDG04LcwFXWkb8YKChpYlf5ycq9x+EIlPPev
6PO2RbXvhoyt4u20XZoLFlQJxRXBtFFS7ibTB3lFK3FMkfDUUNrFH7ldtXNGCE5h
IKT1svKKNqUxY7R6hKoYwpQ34J2v19SksAaQugrkAOgDcdt49NPu8M2g9HRBRVq8
5Gnbdt4ZcQ7y4HF9itN2UAXChf3fFInXTASQZOhVoefw95Wwgm8yCDsE9aUYXZdG
XJo+B07AB33yHg+ep5iJW7kB9v2OchxWe/6ZEtTovejD6Wp8Imf2U3AIsQIMoY+v
gIXIEiznHtV+3r8GZJG+C21tZ1aK/hyGG+BGjy1tLDBWviOPZp1KimwOxrP7VzPm
xvSnTOgTHhdV40AQUpvPRc73RlmWJ7M2tMIRqA/DA6QJijP9N9o/bFCBFmmo4lUt
JB73y3pW8KM23LQ4GST55n+8cfF2EYJW19AtIFJb9p6dy2mtbB2BDEUDg2N/FsFW
Ar01ScDy3nCMngUGFO5RuvKWaQ95oQHfXfDeBDeUOVkErnhnOVeEcalYFgO1u7a0
8xLEeNr974/eQiyLz+cV+BYOEUJ3jnxxtUs/YGp9Edh29Rpsxvtw9XxRCFZu7CBb
NG5Mkw9Vk+r12s/jqSKaewr7C2MA5QV2a1H8P0vQ8oErDFLQw1TEiVARsIq9kNno
H+6mCgSggqCjZB9vz8qT33UtqJrbvJBCaqGfsWKBOvWwXwVp3wOF5T/8uYuvTHpZ
NZmoFwMSC+Vi+eBl9WOj6m8HA6XaxLZfmqBy9+ir1YhE/pLL39TZ3nFSIBPCJBkT
goeGrnE4mEL+6chXFfmbkK+9mvXJnP9T2yusfST7RN9Tpq3vik9dAVkZ8KCDZlB2
fr44InXWqThsu/CsLt7/yiz49b55TzyBn9GFZxEHdm/LIu3lqXV5o+d3bofms/m1
aQGySRGG98qPceyd1gSwKmw/YPfmxYyWEyEEQk/AU5eJB0RT5q+cZrFufK/k3fSS
8qz6p9BdTrlJdz/lbs2GHrDvGzuOA72eNry27b1AJKBdyfvwwsbn9M5QFWGIXmoM
/Cej+LeYBTjkIdQkzt9HmlYzsz9S6ggVyT5aAaHYKJg1ExUNPtqjyiPEDXmnerU7
JxCNcOvQDadD7R0/qDiOIXzlFJ4m/OcsNeZf+HmoxfL+sZ8KueWsdK/NYMTCIFWv
Q25gELHlmb5exxYk7q8ijqlxbk6+VaD4jbA5g0RvAmtGiSRt2pygDU2rId3DSCun
Q74hLGl+oeuwC1WEaym6u+0WuY5nYLzcJ9OqGEi7tz3XInrTpY/d8H0HwQAolYCz
/oEBgHMOVKvsvKoCR9JJwrI2Mi11tUP9M3HQKZG8/Dz2nhQQrlQ9wxLzlgT6zYfs
1fNN9OjVVlGOaxqylnDlm6Phq5+F7uYa+QUei+uAyzJy+JtzVI3axnJwNIdbAAry
oueyh7jp1xEKSNP5IGc7A7MDZPmK4ps6G9VA+CrxldXh7Qj0xqs29k8o5+qErnOl
vSLtyFfpocHXVD3pZ5muuLaPz6YLaUythqPucx6byH1YU0vdtPSyQiVsqhY48lHP
2c/F86vvJSD2bBd+HuTjlTQz7hWNfFbwl7zkhe4T00Kb4TiaFq1eoBlXxRFg/HEJ
Z20q1C45uM+OVuYc2y7k2Yct8zKpQYACZtZhziZy5DIqVUh6TwEv7GfXgtWl/qo8
lAxRCrVgVs12sfPPhvyYiCxPVOGW9DGgrzHgGHVsa5k1h5K/Ir98q9foIeXyJISU
pMw9VNEdTNz3rzJTdn2y2lXq2XWm8BuHR3JG74dGQx4SHXxGgKfTFB/hHgPT/nVm
jl0E3yUmhe46AMeA7FtfY8ULLuSEaPAuOKHLFJfMY3aSBdB0MVCmew64oCoulhJE
jaRGcP+guX5O05/86E0bHYV7PgkFYBiaHs5+hxhvo3cGff6V2gz+7JnvIJnsVyXr
I7kNJCVpNiBJVpY4Tfb3AcdrCYleA9/yID7ByRBdNGmNXtdrMaYvrJsgYVta4OTj
shO4Zwdu04i93igi8uYPCU5hidyDP2ntf/Bto18tzTDrV498+b23WFQA3QnNjNzE
6feHaW9MyxIaKCxBDpGOmuYUNQl7vosGQ5UKECTR1fvHphtqY9OBfwXYTR5PRjfZ
4bkcMEUSOD8fEEz6TNk/NH1xbpkHoRNVbw5kzFeoH2OGVdKG8so4qrOQp1dbSLqa
2ILKfGTDKH7FUkRs/dHm0TJ1l6AK8uJULBITUgP+I52HfRtSSXitJ1qZnmIYgg2y
T0rt5iv3r9o+BTdU63uHYMb7rjpjWKW1Yt0kLZtKpjUCtBzyYTfKM/roNi6YAy9E
+c3KgeWZ4yjG3eq7v8VgHXow08usW4djrDOfsyqwwbAPd/srIvthhFGd3UzfKnUD
rVWQE5M3ISwvOUQ5eZA/DrBNPaNgMKUPD5ELbA0iUS9rbtSG1MZpd+QcLywksBPW
upzHZnvm3xfL631JNXCkIOShpuKFt0xsJNQT8DCxc/thq99Cmr9EMK6KZqYEoCYT
z0uxBa97N7Hkow/EuIqpT2MTMPGbhTAMKeLWpT+D8wDwNu1uY5vKKJSF3Irvn87b
hZoVgTGhuXCwFd3o/eLGI9kQim9CD7cZcI1zJTn1i1smaU0hKFSdFDF25fpXrdfQ
6VlgRGmfVWosB+oVZ4FdJzKy6C40x5ppW4H+87az1777Z/z+B0F6G3p2lXPq1WV8
f/6s0JZ2rF2M4XQgxraPKRRa1qZl/r/Zwjw3M05SJ7LWugo6SgRj89+hA0SqQ/Zs
VcP/aTi6R9bhAcLNxYscxrBmkZANsivC1hwAQz2gNH59K6xXjvCKcjbfy948ADqH
WrqJxvpdkUwFmQ9qf48ONYBMaKkvK7lAgc38fB8ILJjb3WOJDxlpuzw8vx6x+626
xn5MoCQIx9C1GF+Hh4KthUIYwzTgus2XxxL7MrPE1KO1QKecStlNWmJTLZetdxDY
RNDTMyBM1o6b9J7Ol5DMbnZBGw6U65CtPrYI0NpKnWXzkBi90/W+ttYEKtm117L4
mS9WOXhTFUpX9IOq/bGiiCSryAA0PapTha5JcVSDicQ+Ju8g/ODozVtfcqwZIusG
PKcUIXXdLSbrBHQfYb1r3Gdn3v1zHVKpr2fYFAdOkSHTbKd5JlQCb1oPV6W3riba
V8yDBZPjuBzKC69QFUY5ApX8+Np47Ae4C0MQykoITFrBRX3Lv1BaqHD5OWExyJJG
noK0UOR4kKJSPyRVlltqZDLt2jBwOK853Yd3DtNjFZwG/UOooPsG1NR1JQshuAqd
TmtFZ+nrcTniiL1aHSMae+jSbKeWaF4z65xk1b9YOYeSPOj8rWJjrdsuWhbswPbw
5X8HFhTHkdg16LpLURWKRRPEegwVe87SV9v/e48jdS2R9nv7Ftf0eZB5hkkMK88I
90rTyCzK1ltxGYjyt8nMOLfowqTvELZ3wesFuJ2b3t32UvwaFeD/VvMTYBvv+6ZK
7y7upv9gHqLWPWCzUK7FtW33xpsEbKx9AJ+83jnPxCFn/iSIowwp+yKjHuCKmkKF
h26XS/a8CeTMjEm0aimVBddKER8qSuVQARhV/6/uJOCDqf49lXas84CPFfShb8Kx
uQhNa8qLKMoRCXMqjWOIS3TmouhlxkS9BYAIFDcwXuy1e0Ogjvju2ognoTpJoimd
D32FSN5eebSqXN0ZxgtAIpXq5RdoAQhPyzAoHJjvk6WlFDh26twY+lIq3lGU3Adv
r0X9qyLwTsctB1keTk7tu4SfBZlKe85FiwqforkXdSaglH3/+Ur6+9EGs3SWKG+c
AzcCQw1yu9qa3F0qHPxnhxUabY6hw4urtJ2E4NYtZZ2SR3bj7gyDfknAva9/Qb1k
kndTuto0YRx5LqnrJ9HK6kzPO9F7fvmoR/1JxjwcnQ/p92X3qcYjox6Tc01l3wnO
69azPxXMwakwkUdmRCnQvbQ16PNWGmbfcPVYB1GXwBix1HAxT/7qVJ6p7iKCqhd4
rqIyMSJRRySOldX95Zg00se78OU5dTTz6umwDccHPJuQ62UaQ7GXUY/g1oys9P5C
TfxPlvs3lSpYZ0YP8tGN5/u60C6BHow4450G35OltHlmidW3d1vKffHR1upBpOMv
WgpQ3YYdb+pABhs60ZGAEGHr3SrjOhKiWz6sJK2h/1drNdkFYzBh+NcvxAACMBeG
nLcwEnNFB7wydSXf3DVES5LECAHd5Xxbv1XATch+DH4aiaIBZDcArs9AodzYPKND
Zmw+0kCgfopProRJnrxRgmCr8KIj/E/DLmf/qaaOhaZh6zZ6sEjW9Jsa9htI2Xbj
fY1EzIOmPHXa7MS2q2nzZzhZ72wotHjtIJo9ELnrknb4IA3NQBks0KTldYiqw2dr
9oxaSswWWq0K+KfRZ+XgAOC5z0ReIcStYO600MWyQFJCNi4Th6wNK/CWS7YEUwOo
n2bWDPtoMBJ0RjF50F+cynp9eC6JulLZBK3iq8MBNmviTQI3JJzARPFmsJRHvR6W
/7T6+LP/t9LHVXvOq9EDDwirIkJVnkqbNnpgOHHuG9xruyhOfvvCjzaZIVFAB/5n
FcCL9WD0IcWVsnCtFmmQ65fA5ce+Xma4hjU9TMDyepSpfXOGlk8ZUU/9N1bm3EQm
tdQqf6y62cFIMK3jTPJ17M0YZmHwxEjA3JtgR6h3lxn/BmXYG1nqk/FFjBleguum
rfhYr7UiFyGnpW4Asg3QKIJwbh3gR4luSQoJQczqXOY8lVGXN7y22fk9RYefUGOu
5B+lNZKXLqnxxfGwXSG0E/bfUYnTJnZ4i7SjKdUemcymDjMzkLY4NWZmnpi0s8Kq
C0D/uxMt80M1YeiWsJ4rM77IUoLD7pbVo7s8ge+LfbK+ASgfaLLiPTg8CbV4FWyZ
Qet3wq+2+J6TwLyn3vP8uZcGMNVLkw1t5cc2KKAQEWp3OrFc1PSiURMT8iRcl2Y4
6/XYe6DMEnAUv6xpUpscBvSfYbLDdjfU5dRuQYN14lxpUxfolCd6JZeTG8kI7iyf
I8GVvxrB22hr9uSqE4Z2jzCdi8JyhnojuKznOG3OU90y3S+Y1Jihf+RjJesGYZ3O
hURUx7DYO+08PGhHgFA0VT9/q0e+lg+X8+/ippsn9BNH1CZchkLsADvwTMORsa39
TA4TVcdcvSkjIUoFTwwWSf3oaPQ13k7mLWcnl1SA8NbgKeJQq/3tMU3hff3wGqMN
1naK8J/wufeBJG4rhz/pG15kLmo0RKL6dlo06EE0CsiltM1/UHpj0qHcMpGOqgiJ
c4r6Gq9H8ohXHowV4aEJa3nsTvxOwhsGb0F/ShLzzeNs3C0QODPbPQ2uQcJkQEtj
8MQdgHi7mDeLloSOOghD6cTxNJIdVLb0RmUoM5fduBRsS5IezjeNoF1r6kT80i0U
bOgBS1MsxCxgQ0PIPXy+po31Nfv84pDd1r2c/iSEbdIxqNybZ8ncDjBVicRuSiwv
/XZI1X9cyabTE4wLa4X10KVULLl70IEuX4dv00yF7WEK7ALvgMfm9Gt8l7pDiZIU
4YydJtmCSYdvjrUdm703dNKd/KwDnm/hD16tqrmiCR/DUjqDnZ4USEyw7Tfa3yYP
/HVrR/lF2BjBag5ufpPZHOmLcbtkdII7yPzUJtCFX9oBUKTLGW2OyG+hIwGI3IO9
I6geEx/Sy3Yy/FTx0hYfHn9ugAZGLwvAm/NFf8UFY8HXloEHY41v8jt0umkepGyQ
hnoNZ63exYrUTDVd/bJMdrdjACs8mgpAMrH7t2KlVg77xYJFkSKW7bRavt842crx
o+PDpFwh9McOB/6ZAsRpNQ8XGdgSptbLQjxcWVsmDKUeEPJPR7uCW08gRx6RCTpx
1BuQJbM6GPqzxP6x9eHSgDrSF8ViS5m+w1316KMm/234fbXYAi5uFazx7kIorjjn
gLLquYBI6iuatT76woMzXsba9f/R6pD0jG07wMyTFxCvW1O8FJhvz+J/nbdfY0sc
FIkpzXQ7U2kV3fp6OLCZkFNp05ryRUQn9+pLqg0SsYpcKgbUmD9U8wXnoowvL7C3
ZaEI1n3W3BwlvdgBjvq/2lt8fjUUpq0BALq3P1Xj8W9/Rltu7b8/peeTdxcOI01w
+pZF5VJ3dXsNYJqY7jFJLjaHDLFgjvsMh6DiCtSI7/DD4akh02X3vpr2b/n9C6mv
KUdhSiBYzQMWzrO8nT8AS7J17poXkabdr6K1uY+XbgynwAhse07nBtIvUjv0w+kH
r1m0tLtvNn4dOFY8tcXfXglJa3MYxFd70DMpabvTcudmXAZPEXyt0gj1HxcX2VGc
DUQ6+S9nSzgAiOk5MbjO9foMl9PxU5B/oupRiO9INHBhhsubgq4KvDWdYLcGjzDc
xmR24nbbcKgOWANJ4PZXyNHcwpThNyXsqYFPZGuF8NVbfjvZ6DAR4EWdQf1JVm8I
bNvOX1onCnhdAVIFLM+DORN4khuLYTI7wp6GvtuQ3sjUyvkVdGbcUr0vwgh/hYif
n1U5P3xJd8o6/wDE6IBpqPJ8uDzRWIPerSVFAutdL4O04cDMvD4ajbLDP/Xhsc+h
jRRECogjssgooepmGRiJaYuJP9Nqgf8eQlJSWAoSD2CFrAUcQfZSyRSo746Hq8Yo
424+5+YR4X2aMNlZ5uGpAreV5CW9elAqCqWlR8xDojCi1kTPzB6NU7aOMKFWNsWZ
ezuv46ij+QP0t7wbQZchxcoGkVl4XHAoM3LhwWIXwU1LyD304NartDH9RNQDNy6H
HizzKD4ngnuP8dV616CwXQLfw9/rFDz4eRlsP6tNpIJnU2HV/mB2fFIvyg8dFxrF
zDjOB9lwoVURXttdCgc7m6J2ggJedvYUlDis5eHzzafOwwJy9JlDSdA5cXObqN23
fgCTrGwuYWjCwQ8x+v92ROQxGDOuZqgNHB6mHRDDmCCyX+0MQjvyuSwqTMPctrPR
Ewmffbs9J2I0tbjbp4SG0WbQvAd1BFMOp3cj2L8gF+iwPe/nZ2UxY/Od09lNVnDV
70elwkwzq9+h58X+8I+kclJ13cmu57q41YrnoM4NrSMCGJXTL0r/u/W8WjRXZb4u
dcHb29QWQ/ZXbKWRqpZWOfuj8jJgo1sEswss4YDvqKgv4j8h5e9FJUgSMkF2kLa6
/A+aZqyHUXf2BMkv/Rmd2hbNTEmlXyM2gVv+W9TqyKSj3cWoew9TxjdV3D7e9uv6
aqwPVfoGV8BEGdSIp3z4c1PfZv4NP/0jlpkiqvM+YWR23CPD/1ytzczq6rQ5IgOJ
m1R8/AwDBGhiC0z2bijnXW2QAb5BrjAiL2xjMLnbpVgnbZyeKIyN45xxTHSC5bQ1
+xZzUHwa5iko3kPQEAsJni4Py34VrcomdQRbXcZMdZMFc6GMuEq4O6pelhD6qH8O
DSEkji8N+TiBCgOUkepfntu4LSd9LS+SalrYQhRmmyBdRVkN0KZ44B5PT4EW14vD
d3mtyPpAun8DadrSSrNKi1qOm9xtm6v+nCMgU8eNJ5dHhGtXUqb9LXGMe/6vKinF
+5ZwIvFSeX6r73DbUneM//d1YQ2svN3BiRs04GhEtPA3XtqtC2Z1+uf+yEdj5HFf
MJFTXeR5glIl7uvCvgVvU+psQrG3KJaZL5Vyx+sXMlLDJS+QdCqqDt5o7k8OD0A6
Zns896h0eSP+dkDSCeqFnnxUOJeXIklpOkLKCEzOLwzqClnbzEj6xevPLU3maSWW
qJDMU2LjGj/YCDvDNFTCjK0UpysyI0pzHVhiv6TKrEWf3fPdSQY9hZ9dWHm4u5nb
2WTjVGwHxKbXY5Xc0e225oHn729OaoDZKO1r4SjkAmcTgD/fYeDdi2dB92QJO5k7
acAQWUyftDfvbtQP5x+WGiPCIb8T/Ho73NJoielE02Mj7Y5lMROBm+RE60LAgE9+
ifHn7F71xN4nDf408lglQoT91TrG7fL4xyrXRhVFEvPr7R6X1gMgn8JlmYSC/v6k
LqHcJXSBJn/aB2SZaq0rM6jyXcrriQ9r0OJrLK7dFWqSGom+VcBDVsCXyxekI1VD
LgoNY7sBDfvU4Bq5ipcbNUJ5yxHGmRwnShtUeMLO7SkvBkPIae5eGXO5wM3c4ZK6
v1kimxxS6sciDqiJp5ZRAcBh7qYpMvrapFl8AVZu1ObY7pEjRQcnHQE8iuODU7fF
5xuoPvcEtQK/IReN4g9GLbgr4gDcVipkR9eQbATGlBEkkUTqTmcpo5pc+HORQ97G
qKRffVTEKQuj0hlOtiNd0Cpc+CtnCZ2jKCdPeZ/mCkK74HRzehz5WqZDbxpSitY+
14MltsohhxshpxCdXIh24Nt2hgw0HguFhpw6zsV5WkIo77HJD6z2Vdstqqs3ckvt
FOGWt2LnHfvSqEZ6DJDwwvzxi+p9/peew7KCryL4FR8PniLg37SXRv630Yx6MzQg
jRu26DCdxehVAqFVDdAxJNaVZAhYru7xVpGBTlOmrPcJnKwfcdtt/qsYUXjkww/I
V12xs1KSI1Bi7/GMHnolzXbazuzoZ37gg76a61zP1gRK7C175bbP3oIWve9mhAKN
AvWwiKaXiRXp2/9XHAw2J7J0i0h/M1Wx0toGXc/+sSGexIJPGHzX1mD4VYK3hOQt
mFLJgiIPa9VmNtpUj63akkJbAUDvouTyikk7VDFYRNDADVt27wAdTsn5BEIuI9oa
TjTnU27wqtIzMxM03S3z1q51rDmTJrFSlcyPzY+rDeNrj871VW2fHETsgn/d5N4g
x54csTffuRozWCo94jMg9qf6+PauH/jrhAuzNWKiyWOzCKWZ8eNMQK1lwvQTL1uI
3g3Y66xEYQiFAYwriLN4MuYRmfByCitK/AkFhvL0XsPCqrdAToP9p+KrA427tIdE
wiPXGIHd/6ctjQUmYTJpLxf1esy3HQ2IVBAOo9DbuoPPSWOZpbpWqevTOsfe5Svi
YmRq7BvuswiNZFujNlkKnIq9TC7uwS60ypL/aaRfd3etIOvEW0qJi/ihmE4VCOXx
dzCrrPtxobVX3jpppSq5RrLFjx3DkFQ3zBgXZ52aAzkzagPHdE6+W6px2d5WpGaq
3Jokbo8GYO3lDYY2K7kj7PpGnvIoA4cpkP/D6PcSvqh/Rtia5Jg/+EPfoJ3PDLaa
SnbIDV3s6OXSZcviXwBBarSw5DOE3sedSGIu0bS247u5WLhxK0ONnMT1x/hDs9Pk
VgVx7gmM2HdZYnNilEECprWTc/6rpNAeNNDUb7slhSQuVfvX+xKSlYx8mytEge5v
Jv8X+lQpjuGNIf6mWFvaYV3UnUy/NtTO++atcBMpapBGjoKnXpqjc6EtJW2cTQao
SCuE/KNrDukqAp2zyrhfNeZH5QJzBeswclElVeUVNQIHugFqKn56R7yK2tKXYaWf
pbpBiqc5F4UEm0ssDZY3oMyIqXtjHQ0TcXcWi5Hnea5hEezSVQObCvvA31XVfaVw
WFhEjogN8R/8IWARes+Bl/H3awH1/ILAPbSvcKETHe2xHNMy1oG8GE03hXPYVZs7
pR3i2CtISS9Bo1zbgddvS3G6sQwXU8BXWHXFYfBeMEQzyBmfTb6VBsWR/cEgOoyk
nu9rHQIclQEAfJ33F6CSO7ceQ+g5xzddk0wXMzSQGj9GMOYL7bf4ruRAwKuCA/I3
2frnxSfBQ6jW/yoF0ZHvnucW/PmODrdVtkJJOz4zsXQw41fZ6I1sh1v4QONj1Yrs
dQyS5rwT8reVDr2T4qsuGdurreI/BT3IaHDrgWd+yxBo3BkqevE+Nwngvq7VJrdv
fIT25JXgAm9PLhxfRFOUgXWcFIHFMQbAqJq6j76MDo72h+4w6OUDH4dTH70WK0OB
3m1X80KAO//Eyr/KDOahaXP+o0ZZuAqS0ewWGdOSf9bLiwraFAgn6qL1NSkhgMv2
KOUq3NPCMZw5s8WGW4RP8Ib/2CeCOE2gY36YGFULmc7sf9Lx9BnFKO/EZ1m92C8F
QQRSVmAwJXtG9ZDY8bs9QlxVJ/D3DRIwlASzvZRWJmKhGommPnWedxMnAl0LO43a
Nm5tnUiWMRo7sRt0QqOGbznx1dPs2jEKVap5ay/GEZ1mfPk83GOC9C9q304WQIW+
D0CY1gYsEFmBrnUnkbpeoHA1U8Qd+3PE9G/mMMzmupeJbdvBRq8lPqMQGsXrSCls
Gn1mfbe0nHyzMxZfcEM2ualnrV0Apszh7QhqQmV2WevuUBAWJCu+wbHOjCmT6cHc
HLXeF/xNB+RzlK84iFUWCcEdRAk3DCZeKloZL/72V2jwtCkGZQxjqmeS1o4ajsmH
b9fICDZvTsXoa6oghr/GyKyruZ74S55pgAldO+7A22SO/KfJ6gQRuX3nbCu4DDip
HfSDcLLMICzMHh4InfXsO4A2S2n3aasBlPKjD7HN5lw9481RmjjbEufpJKNnllXI
VmvrqrOziv2TDpPGdF4fQGAUnFLFoKbOt7N6LG+XA29tuFM0PhrKUIUiGJ1harWl
qKUEM2HxPjmv4g0/SfTs9qk8Ze9PFMP9XHTYK1NM40iUae2+YGbEbrqP3R2NeGpf
9r1xg3aBrlZ/cZfLrtNu6/DTNeSUt8HkqyrY96JzzKTeYc8YQRfKfkFB8zLnEo/T
ymEnA9sFxCIsn1UjWWC8/AJrJNmNDoC97QgfR85wti8nPTC8L7h4jDpMt9zo9Opf
ZFXyy47EIexn4YElMQxqVnyDJtcTroVXB6AtzsfiiiI14DB0rj+ve+wykKI/s5Vo
aPm+tFHSI95DCZ9VzuEa7XybeTZUQkEoRJIVQBZoETHNI95YP4gS3ethUvA7bdVN
2dcpIeMBgWSB2yGFn4tdVlo2DSmo6Q5FCP0ZR7Z4jzMbZcWnAsA6p3CAH9IHvcZx
dLCat98eJAW1f29SnkOg7A9pzB18ViJY3W3DyMgsaTp/K7gFM4BnUo2CEe0hrw8Z
8qdpPVbUb4dH+gp9/00zqdzvTDZH1ELBmZ3V6V1DQj88Nhux8THEycQmofKr8XQv
CrOuoaBvMiUBSNsapfVmjtaxViTpVBhMHRxOjB3V2nv0D8MtWyOZHqwWhwhTVdUv
TsOxM+iEU5QqVtQIMnRmHlDLuMGnU4VeompwWHbGx7JnYVrBivAr93dtBJXbnE7h
nFcJaAoj8DWqfCm/hK6rvGe+R06gif7wFu82RzDnTmcSDW0PU7wwTYcAsy+8Wv5z
lTC12mloe9WwmUrfxlemHTX1HtbAQ3lb/weCHbLUfz0qT2h/5zUtRRAlfCFe3QTh
s25yRfdIQRT8MQTL965brbw5QyqkbOaIUnpR+h6UGxoAO6tZ6sG1IhlxQNadGQOF
BjujXBi10+0IQGYJAyzDwA5Lv59pFTAWNdVMG+QwRMAaOcFh0xo5HgGTucSqee8h
nnsCgxQfwP6ptio3vf+CmiDnXl+EyT/9/jBy0fNPVTCiJ6LwmeD/Elb1RQfWGZp+
Xi/vaTpKGqO2SpcwNqf7SQj7tUX2LRLS5IVcH30w56iPuC72jbqoTi2jaX2RVd3h
4/iggPbk4G6XocLLKNci1X/tcI5Zh51/9w+eKL/JNdedb5o8WgxL6MaflyJofTof
gT7Pf0wp+yATGDh4V332tWwZTIHAgdc9gccFKwyPJNLZFCP/z2NdU8/kQRAb2Q1G
H7qPkWk0DuNpHMb5NYiJ/8eNfwQdwsfjZMG7YDduk4x3OoCQF33zvQG/z+NznuZ0
ph4PNRInyKr54o53QJZp1RpmJ/sq6/2ngxPyTqA/MYYFbNzI2eQyejAUjwQK2bmp
er06FAAdrUgzaKO5tKnS5IFUpPYkZpKoYey0DKEwal3oK9IqjK2xTp0xwQv5gxhR
2xdw5jTVTI/mMZi4w4bIMQU/hq6xHXcn99B2GgDRaWY62SnqpRKwUwb9R6G0bhoh
aDhokEf83EC/1JTolItbn2i2oGDSdecRs6I+QKhX5QY+3UtYE+A6HUQFvaRcB0Jh
OX6Zdp60O9oZCAb5Ky0/7vvDrjLy/8vgoIRi1PUkEgZ1xQdPhD8Qe8/a6toQVxBo
3j6lkc62jlaax8DEdImmfN/isJUojqiSKnT6xuddwpY00co68VPg8JzQ4+MEtYYa
DCaE5KHfde/lrtwMgkhJwJtUV0D1xpczyeIxJw/bjDvNIcBitcCvQ8/K45lJGDpx
7Wpbnb9gqpYcQVgkdLLtbnu8UtC3B1Q5eEEdC68jxuNyiGndm7uZAjYWaVvHlHwP
oBMQZunCUcG8R3ODF6OuiezD0Z+fNSmRhAB82B3Bv5wg0BodlAs0ddvCayK6WRPd
1SvZfL3gAjEOAgvKjaF+ZFM/KyqXpsENO5SgfuY73TThNtL8rSwiz08T67poan5m
tCYw2m36+S4y3658bcLsDfrur5SueCT6eif43xO4Ut/Zo/sOXxmgLRK/5erHzwwR
zpEbx9T7uzq16mxx1Mj57+ttjfz+7UrgJnZOmzqf0OBckauxjFrLBd5Pjl82Y+Ex
tba2n3968s5+jvCOOObJHre+0CtKIFOVm69/zd+NPIR9E2QyrtJYbuuKCWAK1iqO
ScGIa5Y9Ds9JTMW1JXuKG4uPjzgttpEcSTb3inw4RHLFuaz1pO0tSjhxjm8Cxa6A
741gavfcLCve1LfC+k5s23QDby8kk4JSKqc26K/vcDYTTKeQMG1iLo2m3EcXbas5
wG/E3dDVhIE/NwUjxN7JvkOVcDr1JMsHD1PQDGFx99LEEpNDDfe+v8Evwx4biJ2C
yLJ+Q3jXYtlVxmde5//d0Wjz8o2Q5yoGHUPHkjqHEK4Icz5P4RDuvtDoxcYP09bx
RYUC149XPi2tpeBwC9sxe+47DLZxh5ZwLSf9A4IEVJS+gdLkzMaaKFXKotor5y7i
ulilyqOEP2lupQrylbkaQcyuxPBTxXRgTteA+wVXDntTaU864BNYSJqWhjNLExHE
wMEO6YDpt98+x+onQVrRWGnkZS6j7YLYZsxppcvxLCRDrNRlXj+H2nUAAGn4opy+
46uZDSqhh68ZPPATZEmM6sW7MvInig6mIDxs1K9ai2o=
//pragma protect end_data_block
//pragma protect digest_block
11PVCoUEORuuifyXUV4tmuJ/smw=
//pragma protect end_digest_block
//pragma protect end_protected
