��/  ds��8�g�."O�[�ܳQ��4��j����1 �v��c/�$J¢�\_����y�E�Ծ�����riiFr&<B4l��[5U��f�E�51�3��M33�5���FeC��!@�U�@+u��+�I��!��ֵ�t�5I��?d�th,��b�de�PQ�Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9��J�<����fS$��W���_���_U��L
��|+�Y0�~���97t�|�����Ay�,�
)����ߕ�+E�U�U���f�����.]o������Y�}t]�<x����<H2��9*!Z�o��W��L�3�h�tN4o&�?�����h��%9�Ԍ����7�w������Td�N������^G/�����կ�	�fP�xY���"����)���ԭ�2��X�_�[��5�R4��5��o\I��H�}$ 3Jj���i�ޏ�<�'s�B�҈9Sʳ���0�O��8�
�D[��Dܢ~����+ow�pc�`�����&�9;!�Ϧ�s6%jS��jFEu�vaM'�"�؈��X-�/τB��h��ʗ��M��Ώ��u�#[G�z�,]�G"3�Q��3neU�(8�"kF��eo����:��#�h3��$_a��oh.���C��ކ�/�K+���5'��3�\[/�Gp����\���	�����(IL���L8^q�mF�n-(D����T�E�9��/
G��6k*n�";b���3��*�AD����ʪ"�_-A�s*=�U������$���vnwd��J�qO��#"?nJ:��T<_���G�^�e��� �G�eG�0��$���Bi�&��;�M�T�S��?IS�Ꮹ��c_E���Fy�����:�|;�k���s1�ė��İ��8܀��44&�Fn8L��Q1����~���0�n�;�[��R��bK�D=�OD��y�9Q+{x|�ct����Q&��������"P�<P0�J��&�3b=W��{s���r��Y�mC(�OOu��p��� �@�Dˊ�Vlr��*��itL���^�R��������n��,�9X�T�:��L�����B��)eU� �CDSȳ|z �4S1��x]Bi�(�bms���>�]�8m0�>����a/ t'�]#�� ��Q