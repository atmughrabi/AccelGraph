// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iBWs+U56C3FRg/9oKsHd5Q/sJFXDKhGFlnfCd5W7q1jPavaPhb+zLoqEQ4FPIDlk
EhS/3L+IZevQTO3uni4mDXNIuf1FXE9OG3KcligMu0jZLF0GXD5TiNOTmGyaFY98
TPXVD/IoNwKACZX0CmmHk3WZ0uhrmrhcn17JSe/dGRQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 132976)
FbXyq0eJ5YyNdS/5zUjEudvZ0DwVefa+7VheI3IqI5QwlF8U2pwIfHOdI4l0pj6D
hA9couUDCMeS7aLp+kx/zN59qCe9ktT45OUkXzB9AB3eyz/prvO3gRP+E/bE3y10
3oeZ18zE6j5jWR6y2zlVoB+7JWiB0+X126hO/c1JwDLGE0g+09ijeQdqBUV4dcxJ
tsUtz/XP74E64sdGzZVSe/BGtvhpb60FtJxIK9z0Qy+r6VahBto8uJJC+HQPgPlR
lesMerv9lUpr6aZBjBo0ujjbjm8csiWz6vwU37rfh4aqmxFFsUf0863D+6Q+69ok
hLlLs+H5N9I328DfmyY6J+Ov8sPDWgM4BXAD23kxqZV+5IdHAMUpAcvNEi9BurLC
3Cb171FethBAtqd52LuRUzzeO4YYxVHb7yojbGFOodhesko1Zm/30FXohIwzqS92
bZ953ZNx0y5RqVGWp/QmHkhd5Gq9/4YPU0ZjEjDs2KSxHwsl3d6RD0cbHNLNi26U
ZeWX9fxE/kgI08GZorx5i1YenFB+wpnhfpfXRn1W3HQ0SXyQRI45E3m8Yu2O+aOD
SvYmMr75pAsb0GTsbLZuqEYWPD/P1gCSV405tmKuZeZPwBL+2W7dSllfmjoxU5RA
/zya+anAMPXu+LMfElNH82YV45zd2h3Ii9hn6VKLr2JXFr+V7L0CR+L+IDJ8+/Yt
b9xMe9XiYfNmSXE+Pm4LijL4NQ7xd84hIk4jjvWYWgSPz1/8yze6lsVS0lgZ0crj
8x+LkGxBqlG9moZJyZJnrILxx7ky+SYce3+SQ8QuOFiZllsCzyoWZtzbRoioSaRq
FA3n7YOvB0qQqZomUOQo+Hl0cye0x/knMbfFetYB5go/ZN9Hq5stPyXY5Lf/d4a1
crgg3/37eQsgQxSwluJSghdGtjJrSB7bq+u0SKcbGbPwpcA21hPA/49sgQgvoeqW
N384U/UojmmCooorxe9flNQT15qBLChqqSMMxu2N/r62iYCaVcvh1vMB9QjBRp9w
08imOpBVlfkgjH5FezvGL1O7G+Ma9o6f9CFxE14ybnpWsfZTfFqFjpKIWWh4dx+a
fkkw3czcYPyRDfZ5zZCb/wNgT1RAKgWa9RjTSrzKUiYJXga6d83yfm7OVGLy20tl
JwpyTC4Na8Oi3FiO/TIBuXp5MigzJz291bpmO97UcOjsYuow31RphrI3t7wkxe0/
g4Goc1aF8o3c8bfUTBQttLMZGRW98SETbqmNK1rcMyXq7uyiYl+dAnSnH4JaThIS
ZLwZ7t6rZJjxaGQMp5ah0VRgGeZfIo/dNS9OLyOSd706CVqHl8YgwF0JjPiUpydD
NkSBDIAkk3qt3XS3AzwvmBLOe1KzkHSZkp5COyMBzjH9YD/VLxalsssiR+SLlP6K
V3LSISFN0wqFoXk80SxIsK6KpuJIHV9CAeQS8RVF0bTEbsB3qYlUhugHTjI8yy41
/NG8vRHCYJ83cT4EA3Za1Fu0J+gw8V3avk9b25FpOwsg3/QrDeRzetY+bn6EyM79
LTsZddMFuDhkKDbhikigRgFXDSQ2KXiZWYuEtlyTmo4aTcqQqbvJ6Bx98P4R+xsJ
OGZ/l2ppgu6eSWCbarA/+Rh1rux41Wi3u2HybkedHa9i+Tlr4dlHG5VBz0uwcMDx
exvNkIZ+R6Vrqi8CoS8ZnBoSjp2zi3myX1uLnVDadXl1v82Yy3L5d6JALQvRE7gr
PS2EEtRa3KqnEnQX1HzHXK7lhH5Bdse+YUS7pCy0jP9XEcoWO4GQpSIVEXbcOnr1
SfVyxmAaeatK30sPd3Ri5rLaxukhpZFG4j+zoqMKdiuQQdNgkkLLK7X6DGELnMZD
aqeeVM8gfiVTD298/VA1B+P1E0gTeqvmPg2DmhCBlLmWz65HD4Fmd/C2LLayeNk4
b2moT80Kn5oWSmkWGpCPvJ1IbaJmyLQp/315Cy6aHmTbT4foRgeYz8GBJlq47Gb/
4WJKwOzlvrmItSZplhSOprx95MPF4m0856AU+X/rOUR6ZEy/y8f2yRTK/46oPgwg
e9yY+2zY8fXjmuBsnTjCX/K0diO+nIAg3p3PuykshL++RFS+ywB97Kkb9brkiaeD
hZhtXD2LYAQUHO0F1AFzITqcF0V3i4cPAzWq7xYl0k98J+qTLTrAX8/Og59d74R0
of8+A5kJd8wpYYudAq/cHTpUDk0j1Y0K+NoE6vcQVtmazLQS7AHmezYvGcZfcXI1
khsRQ0QBFCis4ib8RE3dH1g4o+XTu8GnCLwcoaCWPLKYQO+ER3QZwj6j9iJmBCFy
wrfinmFmrkao9wIimNDoyGPDHJdTD5ooldbirkZ/2IHY3DsWWaAv5jO7FR0JCr9r
/2wRT5NhV3o0MVqE/p6IMbFxjwUHK3+EIevVaCYW0IRavh/4o4kNsPv4aN2Z85pu
8nD+VPlj1ljcO4TJu4mlW3aPzKVE+x/GVO9SS2RMpd350w4SpRyjFJV/UvDhPDGc
vH6rdPcHgupOqw0TDkUkCUJaFb4Y5jNnFbEc87AM1pMtAiBC5AzieNhGXVZKaeIh
tkc0A14TJMWNpIGWb5o+8lPzY/YgjzPdWQvNNQnqKOAJNOwnznHP86eyRyFIwYFv
GRbs4QYrzTiwbyNnrTA6KhqK1iWSg3xoNH6RUrzRyoWYQfqO4u9IgFgn4pitNqgg
ZZNgt9td8Ft/ctRsIJwfMaiyz685U4idxWobwWN81QJVn4ch8iGqtqtnOr6uY5C5
nWqdQMzMQg2HEWlekfvRCeYTuPmZYudxGwty3ECdQ/3CacO7/26yhDRHPT3vHnaz
XWPhA1TvH8aaWXbt6i/MBpc65V6enBZH8jfXEth9JbnLJGCo9Sw1sOhgQjeKOB0S
XIKcTPCFQFJITMvPoUIr7t83mnuAS42zUznEOWeMzwdUMOc5TgHju3GMf5oF6Osi
OpZlgmsCZBmTlegx3/5cu5pSos8Gy/ir+9Gnb9GgXzg740JmjUcZVntUp2CP0jlk
wW3EMtBBxdZg4ID/blvSTtQw2uQHCozywaWsE2k1/7kIMtK6OQIrfP2NpdL2Ms+x
rcEUWFIkCuhqM6egaNulXVC/ZevJE5qv7so5VjfVT4sfmLUvHrz+3jzHPnMN7vaj
GRtTZmZ7ScPpHIp+VU2AKwYgXOJCAWZYSV+Xxov2p/y6VCKs93gn0DcEaS0cezO1
CAEWGlfPodjUCvG7VAA2wYl2Rfh7qg4kF9jdvDntbgAZXnU+CA8vpGZkr/To53iB
XF3ukQSNVC+H2DkUnboFwG1hjw/9zKEuVZs+8jZfY0sncODQlMK2X9O+EpcGIxBQ
GRyLrMLpM50i/IA9pnKKqmraa+D3XggeN4IVv87NjbMCBIhQ077nh8lRwZFLYuoc
8UZcF9HhlNSJC/voF2kefNxUIAM7T31dIfTpmkv5g7G75JtxrpNX6Yl6wr6jYWYF
GUIGTHVnMxBIGp6G2BqtMdFnqnn8/ZWNJGBFx88bLQPULNWS0TpZgGOeyR0H58am
pPLyp4WwKJwZLgb+YAHlF/SFv/Mtq4eSzbT7cmYLA3aduJAsm6dwAunyxzvghcSH
w0vYtg5WHnQgrLvExhjW4ZW/BJ0k9pG4dIq+WzH8N2eY6qoTUX4vo1ok9Tqrr+aB
iuGXGmej0v3pW3OXA4JK+0HyEgHA9H2aT/IWqY19Ro+RhFwuEya4LORkVhdDOmGF
8ZH9L/7ibB7j2K+S7/PJNPAFgf/2rv2GyaGtBP9OtORISY2Gv2xN5YN5bjFvBKrG
K8cNDnzsjF/ICRErMN9QUOP7rTIo2l5EyT6nevajfHEiMwuAPjS/QqL4MVjBLB6d
oelB2ZaRDGESdkrigAbIbxsO31Wb3hILGdmMNRnRMT1fBv803OpvQyE4oxcfcUtl
981aUsjg+ZpitKhtGNHU3Jqc5qsSkuJEgk3arLFOWnOa4qFex+ersXwxSaJJJmKM
arUa1dq1pgBBXrpbbjOp4asCwU4DEA9di/WRIJ/ibaT7/69s9D/6ZNB2Gb6Rzxea
qTtJ4jnBM3lch01RYJAxYEzLsXmwHtgesbEAcOdr/8tX+hr7joHHJbKBB1C7SiU9
5Zbg84yh1m7piosp/HrRVUMsD4GzWNNHXZBZEs0yU1/NveQVsjhLzu3EXL/tyPfC
UE9gN0rqFrcZ1ceAIpZ8kIsOb+a2OzoyW2D4IxrasaIXwuOpR7y8l7bPKOMQkigp
c6op8vl/5rJfTH8o6qMtMyKTrtNcZZHoYZI1A++eJm5GG7s019Rio5h0aOuCp4d+
QZCUDfAxNP8EklLl05bu5BEAddmxMYtHmFH/Ag2liyoojnxWD9USIKFcYRgLYhYU
cVjmNik1gHI8d4C/iMW+mpPHtLZ/CRoKsbvuwEp+5HKxGXbIy/TzgGYjkrfSuMrR
W7SZepjQM+jQFQ5eaB5bGCaQpXD8w+4kZiOURKw02XluLnCRP/7s1pam1zMZLlnW
cXKpdcxpBPoUd7SbQntTe5vtrgBD6lN3L/M+NEpWNyNHTcNU6sdGjNt9pAfEZAtx
I4kBagBrSzf41TE5o3dEWmoLtp364PkW7Cok1CUgaNmKVRV8OLOOMWEDq9R/Sk4o
eRijo8vyrz7LM6umvCzPcD4VfnH3jbYN5KexM+YgVSGLITGbqUQL2wVvFQP2u1rW
w3mFUO9O7VSjhwN2pdRW9LN1IldBCmmkLy+jbnHP0jvDUCIH0HvAFTrjAMk4AjkK
1cBog7KYPxAWEkLq/YnmEumxmse62cKP5gAj70T4MIcSQl0bo0A0Ew+42VEXrDti
xqkkBIU4e1oHoJKiT2EgSv/rZfRl7wO2f2EMmtJgjdq0tEYggQJdypgcoudhnk9o
oRzaiiVWobey+k4dIGZKuPR6O8zsCEhL7A2Qi99MID/2HnsL88VOFEVnGl+nxYMb
f+VPmPFzQAZoHfN1eWO+fbkjT9nd7vrzWDKSMvO7/Dsdeaw/oi0jWy9n5EbhSqM5
JGweHRpZJ8zQIPRKRTT3K5L26k166RraWuTD7MtyEVANw9n1oK8eIouMz/AUGea7
HfYn4fUtOsiPQW2fBCDsy++ByjRBgFb78pXLxfwC2EHn2AiJzIzkYm7hgYPHguup
FrKluZ8iC00piLju/H+muIXoTxPBNSiThgYx0dprg3Ico24LLcbfxlQlkOkrgOCQ
UAfPZaXGh2Bx2E40UV29DTPdvna3vrQsoF+YlTp6tQfAwiHfRIqKHXgIKUQAaaT0
Z0eB1lgdMJZTIPFJ13HjJSn4gTLkhrolgdo1NNOLrJzlj1Bw+kZVyynGhlPvalnN
+EzWNGQFm6Fig79mpXaCReESVDQpZ9vfoAdHflOIQBldnuw3m2xknzDzbXZm9/cT
8YxNerbeJ7hYWNm15UnCMPJkGGwgqLcxD9XZslapStCzEI7kN8IeMCjfWPX0LjaL
c/sGWo5BqYTJwTJu0HrKixWcWhWeff29sREpu+XBatMf82byKFp5ym0noY3KJNwX
KF3zOkVhV4KCRmdvpQiU9dyXUmZhoT766pZ+2rnr9+xS8gFjyyvSTdrKDQ39PoIs
qRiFS9kHuQzSwtl6j5K70YwJFblMvYUSOoS2D+5lq1dZMIbcoEaP4D75Iv/X0Ltm
UDjHywCTQ9YuAqpNX4FioBXCrFHoyPmGVn7Z1QgMzkoTyOnx6gpyLOMnYMQNPVjC
LYbiWLiz20ztZhPDo76j0vtj7dFNG7bWzM2pWPfv8SkKWvwkEozQcuRa7+NdDtLY
SGeZvPSS8L2yybjITKdWbWcdGBB3/ighfXZF2qmKVyGtYrtr+2LxGyd7S/3HrwYA
AsxCIin2MuWBu/SkJVpqeM+cmgV5SLVYSsJQvYXQJR3r124PmNBmGYltjCkP7eZz
ps+f1m4jSepw1wiZATWauphclPSeIJ6UHlU2eQjhfRpAGG4InPkhbzQTVkfhnPvo
EpZg6lybmNBY9RqyVNegtBZUDSpt2TwJfJK4ZNDIVfcpIBnmsPsdfr8ExqD3FVLp
2CxiInami2qzRSawQxvPjJsCbDAdGx47o7GHWdqjL6nBPFPxpCkbrNyFCYRm62ON
fEgbF2tfFEXMXcI8e2gVb7dnrhffFQQJQJdjSZZyP8B/4sYD8Qm15+dtI20nO42b
40i/NSm379RKYTAK/k8X6dDLTVp4xRsypo4m3LdBzY7PKeS8f17f22U9/bQzWG2c
JW+iFLZKlnaojskC0A26WKMmi5sXnuBNwWFQ09ydmUzs83rEmP1kfvoSLUoiPbF1
DkyQZpcqmpoDSzRnZTTMBWgvWqT55L+bkQiRCFJwzZG996gP9lEmcTq2tGPeNUOj
S7mu2dEz50hzLa2lLKe3F+AufLUYzOQp1V1xvKMeBcA1QktzDXSG+6rG1AfDGZ+d
BxXVcIDDvC88gRqXQ9dVlLWVn5i+m6Pgs+Cy5FQ8BKxBsiG1hwqrhXO7QuE4686C
yxagX7y1UdKiO73Qi6l5wGoJn7Pkbi3abVV0ZkXo3v4AWhOe/Z6pxn59+6MeTor/
W8nugYZ5d62SAhbuK2FjpPYwyF9oaiQVd9TlVxxVlcZlko3Bf9eTKaoigSJdAQKK
1hrsGbMEq+1ya7bBMjrZ2d80xI0fLXUNtVfx9bZ1z+NUwyte0EmHgbXzqdlV35iA
eNKPneJiBRM6k2NjjRxBJhJtJYC0v5wvAmH2NghtflwVqooeu6uFYgDwoO2fmkVO
OHybrD5U+9iz5dCXec7sss51KmBVvJX+X1dX64r3YRbLxDWO6UdaIImsd0LuzU6Q
DUET999cVn6jYYltZrg6lAA6H/12/6j8FDSdUu8kOtavRaf/XCZjKZfw9gYvtqKZ
VIrGOlKDZIMdcBY+AlyHEdzNHIZiAghKLCcefgXAsSWaRJXFR7d0nSIpEHa69eDL
huY80w9yVyCrhT+GgSB+zrhWKbcwSfO04Of9AQWe5JYH6w7a8ciy8EuF8kWeB8Ia
ipvHM3NFQA2GreaZWvVyHX4/f5PWbj70ZKJDJ8+gnERFG0mzas7/CPVUQKN4BZsy
c4vLCjvLWHnA34veWUiZ50BO74+lPPeRz3W6y9TRCswaxR5rI1EGeD0LSJm8xoL2
qQtmDSJSWFasjUodtp/zN3sgfwf6NL+mVQE2s1A/uo0dRlVaJh8beEYlwRc0WHZd
kat7xezpCcbh9FziJYEdty4pKtsYFREJyr62qjVNyYek5WARlbvHD9Up9c9GI71B
NA5ArnXisVq+C7ek7PusrwHJTRK72dp0YNe2PS9DA8zRj42zPXYCQu3Mge0aiJ0P
oSwbP8rnhBLohD+aSKDMzOsyjlLcLJd0aFJtSQBAk3t9Ct+CFEjBhcYD0G2HfNra
DHcER0yyuyArpU9T/x8ctIDEuOnzOAc092SUt9koKTIWF/Zxg/jAtSjzsFFhFJmJ
WZEXiPMyJPQyH25gNSQ1pPKxQtYZwYYxobMCrKTAVArjyR1EVUv8Z90L5pxumoT9
H7oisNFZbam73VWfnR0bJLYKx7VlSFsZ0JmaY/Av7ngqdsKu1oY2lNBhA1tnpEv+
efKoYPLhONGnMo0b1tkffZNAPLc3OCgD23EpMempbdCRq+vRHwbSoWiSiJg5fTvS
QmByN2YdVmaLc9oDjyqsWloit+njXZdClBVI/Al55IjVLC9VzQ/juAJFI23zLUC6
tf2NXXPCY0HfVjUsXViUzLblKUHSwZpvPBPQihd5+galRMUFIfx4ZVbBbtM8Hr10
H3XkqsRD4urGNUOUGzOJWasxIr7xUFvdFIg//fGgAvsRhm/0WMt48I9nQMFJv1dq
n902T3V8Xl6h5p//MJ5kbbfo/lPOPaaadMUAAi3DQ3hL3gDhFjE6eXbEHnqdDwSI
VfO2sqpWR9fB3dDMT/+eVlRzp4zHSYtg6+UGAbihCnwhyCeGIw6r3MT6xZH+JJV6
d9vFHwAULijPuEomft8TGzsWoymMYDdlj3XDcceG3bMWvIRQ8nLatLG7xwqmtAcC
OygeLfkPjwrwPnInvYv/9OobKgmxwkhnDsvWUexchO1fuVq/jdlElUtR/JCdVu2Z
cHa2DJItISFZw3pJfwJ4mKrH+AW8C2dPGNYxHjhOd21Paeekiw8AEY3hqMglRgYy
JsaN3YkpnshinfFHzF51LA6wHbuyr41NmdZXM52vqWNM8jLm3Ge4XnQAHzV4Sri6
NfaQM3mm5f6zc+NYla+0D6jXoAfWYgaco5dmG1affU8T+opqoE598RNv8FOoevZg
NHZbD4ZiD6DRvWbMce0eSUa/cFvow5x3Oxi53d4B8kP20JuJihXRXDCBIEUrg24H
DPap0sgqXKqv9Ku0f8CkGDC3ZOhCHb+9ktOluBK8KXQc46ro4ZRIEcSsodNcRX5S
NyLxmymAGcXta+qlON/9fb8dv+yMgwM2QOOgCOtLscmlLEjJ4soN0yZNFbEn+t1E
L7Q4RMgQnYEndNmKXz9pexn5sid8kXV5IVPwforJNwR3qjv85j8Ks9LMZWFOwL+A
ULqCaMGiMQzB9WsTcyQwVUyO7OTNBiS+tC4Ou9+1j32mdmwt5sNTB+h6kJBod29V
w3EwNP+WkIil81q596KuHTJ9pjl8vyyjHaJqCyfpqiFbEUOUKpBral8K3T+2nH/R
hixWeUqlGHge/xNAw6UjDCXd9G+RqmU91Ed0eFeOYDSM2gdFGhOOfLMccsqRVGla
HWGD0qoLU0VcQWHpm/wKOB2teklxgrbkD4Xz/2HtLOkej7BqBi8rxjKDunRvFF8P
dtAlEmsL9zhQODmUDN49V0JMMBIVMKFdfJ6SOMiuVL9fpPem64S8tTQrCcDjz7iw
hwp+CKHIxW3z+n6cRZRnYxMTqqRaqdPj7tqRu4zbTkIqTpF+lTql31KjBopUeI4F
i+SYH1W5JmkCwstVnCh54JPC9Gd5V65LnyLJVXeOx2arY3JUpYaMpImtaYTZic67
dR9P0xSjy6HuHN/ShSyIcQ6qJJFaRp0/Hc9SNvet5UsiuMZrdNxJdqmarJ5hHSyo
a0YisarJhOYkDIksD3as1fbGnSbXAEHJw+kfNJxbbiwoGW5e0fujqme0ThKP5y56
lrXyVhlSUWf99RbbRDfpJri79o9tQwbfyNYsfCpE/GjBKPpDlNSeFrgrTVp4hQrp
k17nr9FDTi/4owdqQZnfWdGfO4wEJ+tjblyseMBx75MBV/sv4+VYNL9twSQURHNA
/eZpJepGa2yUoSv6N/U+cZvaxedBWIkY/ioNcaKUd7SPf9NmnSekT+gl/FQxOPne
qIfh9KkEXJxS4Zgx0fziMGGdJyb5j2XKzn82Sf2qgCVgbapTF2uvDI6SsAyfhxvN
BOS92Le4mIWi7KmifGBBAbqIPF8czV1eHSnPfUjrN2Pb5vl0t5aMJTBClywi7bp4
nwxo4h4h/pjw5OnCKspExyVLA0mgvnLY2k1WzvZPEUu8nZPATOWH6Ba2f7GtiKgc
+ZROdCRytf7BxGMbwiurc++mpVFWjFACjFYCAXY4/9f3WdYrvrKi8yuHnPDAFN4a
jJRXeRH0KOYrMsELswmKB2sMDGJZ/RY0uzllJqCN6WPFwZVM8vexmr9eYZtYMado
pPONh7Duub1mWdrsM4cuHeypdRX8CMd0Vl/RI/8crQo8PGVNln8NuHYTK3hqmotV
YDeEdNYDZVd6eL8/GQ0Z28SKsYXAQqBuUhFJX8Jrzy2tETTA9gfXI4b0kdNbKmJz
P6iGNZRQoo2bHmfiWPrVJ1TG9jyokHGTiAwojfjrHgimbnT4rxB2s2gXfL57EYX9
8cXLWL9EibsfekWkdLjbFj+/uUGvwztWK5YF9zehDmIhezA+ECHOG8wies3qADLV
S5vJIlj1Tu7hyuubXwMFKFEI0zxVpcC4DWUI/Ba8HE3i6Fxb7yq6VB9crw9eTpQA
hN3kNuhKDRsKA2gllhfVe5FlKS/cDF9/MH+YTDMR6kAqwL9m3Wp8vY5L5kDb9xX3
LGDSXvx+Xb5dUmM0tjGFh8vipVI0BO1jD4NuH1ghxgk4hhtBznaCa15Pqr9aajk/
7lQzgQ/SUw/4cjIm3xPCfUVSh0YWgvhE/8EafcdfpZhPNeyNlKtJ6ZUQ/zB14kd3
HU5Akzw5asWKKCCLOgFVmZBjDUOVj4mJnEdG0Vz5yZyyGyiDNoTh+HETevnc8alY
FiDK5TqHLtAYtv0BuAAtMuv5QyHjzTMvTeKYswpT8ZhbiBkAOdu6fVdGlTTLpnPD
FHy9TsEsH9/SEF166h/bNM31/qw9PUafVZ3zzUohzpgmz2Ea3yLo6XwVplyHUiQl
AOIR9hobqDOrEJMzH1MNkkKHJjYYCzc9FAUYHmn9o0J9j8HoPufn+6eV8qrKE4Te
+MjYxTn0rDy4bRTwImkOD4tGfO9f4OrMVInUPNcPdVPumgjbH/+qjcuGpBaOUEJb
NwIZNE4lEXyERXs0Df+9ImNDlcTL5VBpBXpeMArUwagNPmwyvW6XDJkTIbxyzR/K
i2jLPhlOWNU1V7Uc2NYMeRPx9N6G1p2xRPD7iXvS05HRqhFz32itPOszSUygQfUo
d3T05GjbLgWSk5gepHRGrVBVCln+u10vCwcUf1iyvcTsa7FewvGLtNpIQZ19GCZP
ajIHwUlrX6a1A7uJM0j2E0E62uzzHIBUJPdo9RRQ+pdRuR7hZx2QmKV1XKdkBrQB
j/fBUHfx1as79R+XEL2iY7NjUoiUu5G3t9pU7b6ArzJjhlUdS2DyJI6tHKcUbe8A
+1VDt0zFQtwcX/IM+0jJb75bldt91V5lQY9B1icOS+GV8pYDKnmqqZBLwssuZWrO
wippt7SEsW63q8iVYcvk8pZ338yOZm9MxajwN9ud4stjXwayF804g+oxJO0EhhIV
WZkK0lth3BoiBa6XJi0qnjGsOR9Nm6U4EigjTvC4n4LLCeWCZjWkhTToNy0mzddj
a3k+8yNqLATcMAMTsBijArY3Y9orRH+KNfQ3eE/36NAW4ZHDmupuXLwoatniMFmN
DLhaDURwGqfIaUpAEjj4SSBlPsMBfCQg8s4QFDslqHOo6STy7S44Cv2iESZrMTD2
klvQD3RDsTQdF1cdhg8BlKTLPlqJ7Easf7u5GSC7/GleCYO7LPPTuh0rcRxkKN5n
MIRSQcoZ27CzjIerOsRI/EtZQorm7CDdcBuPVKD9uIZh8C4FpeCF2L05jMBKPn0p
QYrGb/zMwfE1KL4LTdMbqpWphNq/PVbIb+4DumiPMeYGeA6R0ECHaBir9LP8jKYt
6zgmxx1JB/6yd2NI6LIjV//1ZNesLKiq0MzUeyv+8BUMIbv3dCN2EjkewjilIbsx
k+M6pyBoYCw+dK32gpMAgykcht2sxdnZgszhumJAON/D7m24s9p2tNATyEdmENoq
9gH9g1HoKT+QPu4FK56bqKKq3a/5r0bwR4cdmpkGq3HYsYg/awxeseDd2OMLcA9X
YgY5RVGGVG3sd3x4m2Lee7XllJU7Kz3tGnPBJbiwQsGjIJqDAba/31FfvOsn8Dmu
YWoFmNHxf3nTiO9hu6T0QMT1pHZFoi70Bs2CIiVNvbmPlNSuXQUkJbh0oeHKNMF3
lRdygbo0+4MzDOu1FLCtghYwURr98lfbwrTEsIF9wqY+zmF6fQQxAuglSkUgY2s4
VBVDZY+QqJo1PmSYOYvLzTzHO5wlXIVhvC0uM0SHOK2aIpezAay6qJiLM3PzZuBF
yj76aI0e5btotrzunESgeyKeWvwtf8PxNvXz4nnim/P0FnPWbuuVhJh96+35CFKU
3LrFPx9qZ6hmo1qGiCpwjYKy32Ory5K2wZULy37Xi3ebxXC76yOIMWExJF/UGIRz
ZkyLufkwVdZaLm5jLeCR7F4uDF9X9QZz5480HLm6UUEaoidTBeHl4nlAk9tG+zzU
fqAFYJzyGuc2awLhbVufQd1l6wFKzlY1sMVMGSyCIJMhIQ+n/hmaNPGWCwar1Tia
Tk8T1zV8nTyrsCu+FzqoRbRzJTgHbvBf+xnGJYGW5UkOFTPMDIWVMGV+fAQ499QI
lPKz3R5wMFqi7Zqt9Pl+f0taiqL9oF3r7ETgCzsGaNaWPqbW+/wdNJBzBj6HRbUa
pVhYAc9sRJCnqg4c9U1qw1N1AGy9JMtNtHffCC/EorXNWdC84kR5WULeAa0Vrqrd
axU4m3rtA7wAe7UJa+xmGmMYfPXu/mIXdp3U7ErnP1qtQP7ovDiiI1X9X64j+maA
mZKfGwMQODzMIKihe56RcnauEmP6fMNPDo3XBxCN98oi2ZAq2Obofq+aYqxU7KkX
5hlymAeBheJ+k8qLtJd8lWsI9ESxrac+D65BbvNrVO//gB0UdFBhPqw9Ph7iLVNv
gfHk8eF9FJ/Wm76KVQ4EDE183aKDa370Yywtzx/D8SYkoli0Tws5zCDeofHHPf//
teMLUL1BFWDdLApRz+PD2GTJ3BuSuR+ACZnhISEpnWuD8T0BUtfx/c61fW66Ejyg
msrxmMEe9+xaExPP2Vy+7NB3BlCuRJDzUPZP2AglbvP0MmDHCUCBb55kGrVJxXnv
A9oPiF2mOuKZPIsXyiYLZC9beRN1yH2IIZNg9dj7Y9fz64CaHqp/tkRUev6bMZzb
LuOdASawS/XUr/U1fZC7+/t+Dc5+fBLEilAif+Hf0jLPticlv/0eJKyrFF5X8ZEo
K6Z2o9HG6WYbWy8c3Y+NHSHBp4WyuD92qTg4dQ0029uFMklAiUkSWUBj23AHhRS+
V0yV/enweeNwrk7LPLxbbBLxeIsVq+ekypYl20K1YJ0PPWYvhpRdz9c7NRPcIACh
cgOSaGbQjrYhcYltDU2ylb/SrkSGQ8UZgefgNnH2aUv+Pd/Ta2K0H/XyeUVXuDLo
lt8wWzyOso86NbjDyqtjPv/wV31Cc1bcLFJSXRmRmXQ/I5S2MzTKn6nT7CbY8rd7
PRolZ3z75xv84aICeNklofyhNXoA8/mGvvcHWyv9Zsx1lMT/P63txQVWV4awYE3Y
xPWkl64H3Ckhl1H64z5DoQpo2T7PdqlktTbwQmg7oJAW8zh3xLnpWh+DG8J/aZL3
l3NTB7G2slffQZNwUannoPncNkFmb29DtMlTUkFXLGLnLnfG0VTQ5YF30Cqm6QoF
FACcVI8MUioB02lUrWHrN1BZozDCH0vrWORDyRWGqsPNZ2O9bVotE3ZpQp0VMWUv
BBbahFeUeO9UvfCRJ7LezZbi37ah4HXC+hD3hPHyef4az/587udvs3EOMKTBJQH3
lTxWXmtRUCIpUhvKNvt0XmCG0jP2SwtYLPFlOm7vrRdU6Lux0cfrhV+26wea4QlZ
2RglKI7e9fENrAUdcfyhOicUj215lIA4Vyw6gCZ2+umlSMPuhOZyswoogbppKlrj
oK2pi/xar2/I8RX7zTSL70a35Z+bUZM19msKFCiKYsOr1vfpdXcHPaRBTujv/Hys
3hc9a+yqqFQxo6aU1XH1Z4HLdyN2Wc8kGm1UaqBU8zhjgMJFMx71/RfW9RJSbitm
YXyV4TrPenv606juMCXlj05KPmEROCTqCF4GnTZKUHVY++7WE9wgTXh1ShePlYXf
rlgTFNKA0Lsy1DXW2mEOwQO5smQxfEheIkTf9Uq4ZHz6p7CLg1fH2+XQWbY1OuVh
yszMHflCarWykaKZgVDqYwGkCgA9LROQAqMdws8GWnWKikv9MUjOEW0MAEZFgO7I
rnbBThnPUF9FknfpHlhxfepV+WXNj6D+i44aD2qDa5RyJSCiQF0/s9He8pOKZgGy
B3gTCv/SbyEx+F0/5dxc3M/WOmPK0/K4++VBGL7W71k8l1OjKL1clSiD/FXhmDla
1EiWT7xWGsepmxl3dEp4y1HqWskTKHPplSvkpdjF6Bg1CCmdyXG+euIX/0Ug3A2K
q2XrbN2gnM+evqd2zwaKnnIFmBshmtsTjGZF0xXUvzTMbqIQ15gWtcXOTZeaNY8B
cwe22oljbVhaRHpHJz4yszk6Zoj5g1xtzAqFSgKePyV9VH9uV6uGdB3rFyXGcwme
i0BEKPhmUEW64MfChbgfsl9D0vH9wm/5YuEzShjwJkdod1+EHgHLG7dWVccOeIgk
znKrT593ANuFqnBoImGjSMtBfNK4JSYn7o39KYeGpVGl+CIidIM6QbIMyp4tpmmQ
dFmFKPpVCUry84HN5PPs0JfkmohmEUnz+hIYrdSZN8Lc27M1c3Xpwd1G+AqRVzNT
3UiOK4B30VK1dKG18h9gCzId0msyvruXc1CWiawUt3GCht8TbqTDBYYHI2tZfZYQ
3ZhOZnO+KoIC/cNtf+gQ6NEiw2SmM3R0rzD0Q25g8r7NtcQPz7r0eG4864IQbOZH
LKP0ESeMhwEq6XeIYK8hb4phpbfSjP9VcCF3uodG/Sdn27+28hz8swnzcE+3DgDo
knQHe1M4KvlLuUvBJAa5dQQhiCtE18qjk0TGM/ss9xdMPmS0wgxgl7x7tWdf3fN7
Rlxta6VCQS6u6PfiEeWi+hXrNdwAWEQKDQJrtvCpNJ31/32BvNvQYtOEXQtKlZs3
3zUc3jqLL84wQ0Z2mdgftCP8x+4gzpzb9rxRebwKnUpqlYxE63uG93mkfoOuhdvx
dtmmOUjBjKxoeLB97WMC+G9028/mpgqNvtCqhJ2mplbc77BzXNCH6NoQ96W8FK+D
GOyNZrXh6iCyuXXC44/lSnUqPSvy8YCxAO4MlQoVtq2Z7dQY4re4B7r9iVIIYgSh
Q7Apev0wKyAoSi7g914LtarABAF/bubSA9WRGBkJ7Nygfq3SLrAbKxeJgwVFDT2S
kaFB29JgHuleCNZBwuvdAtYOc/lTT1txTXMcDndoYreaOvdpWNoX3d8y5T+lBrpn
Dll21lABH7u+RRl3uJTpQu8aP3GnaaCgMI6qX/U4rYNtYEz7dy2+kPAQvwyMJDpe
bmFFccZ+cU8t7S8LB6A22knFI9FDkEQ+QZ7hb49OC2GLETpEAjoc6JqLtz9r+FCP
b2w/B9J0nhey9b+uJw3QfbnDxuo9W0nlkZ6fEosxy2CXYz398YJnL9oM/GUCNWqf
Rn/lBlkpcOp0fj/s0C1WvTKpSUZyzMTpqaf2xCqivtuYe9lVQzKcOkwJaLVG5JO4
D9IO0Bwuxq5t6jSjB1QrtHOjy7p1to/oTJysWEuAo5lqyBPCvnFZX3Or03hF66W1
9VvGheOPEAmNVpc4qDki0Qk2eGZEqjv8JzbAxLz+dPgCohYaZJwrZl5MlB/FT8iF
NumI1V7zPs+xzlsyQHkxlRRzo4xDBD8Ro9eSNuS6HB3YNgsuMarBmI/Tpt7oAx0y
lx4/JZ/pFl/xGNLUkrc+3/xtensOS5OVShvREOxhy8PTjqcQrqVlHXFtGg1N455e
IH2oVclt+j88PSJ0l4/VGxlUq99X9qrgjnJ7ry17vCay5PM88nTO1zdtD7ibf3Wz
jYhuvMQiPnh+kuJilhcB8ofVTpDcL1QIAkyBevtF4kg+2UQfs368zAWIQ6CG7Os0
K9O0yYtjGIsIL3uh4VPuon9ed0ZBWd4bos7w4NfRmzn/SvU6r/34gaUFTNG5zjyQ
duoMJ7CVAOArdUFfUO9OrXqMWyrGiO9e9LJ83WFeDJqYGIERSxa4Pi/kMCG0Dlgg
+QZlEMybUANEqMSsD9soTnKCl8CQxsQyGvJ7KbGdcfTIOExDpeGpWSZk12DJIB/X
NMhAOFQJ3N2vVzJ1Ttc86pYWU+3PJYW87yyj3tGIarwJc12IqcPrSmqq+YU4CSgP
X7Z1FxHxQe04c7XAv+lsSG2LhS43N88lfDho2jrBCBz2qAMl/fS2YaPYvFWnSdSH
kNuVMwJpTynMK/zNygx7amkJiSexWEZKxMb1z8yuPkBRLfJZwUw43Ah4wyGoyTnX
cyDx87SCVY7mp/gYqWv2iuwxEqPBeKM6tml5ahMVYHxqlVzfJbNuKL8O6e8WwbTd
KWTqmMLncRBgiB/LAaY4HBMHCkcq3wzc6cjpjl6cU9DFK34fq2S/441SBW3KfZm0
9cS8Imyiie+rDd6BszO3HCGqWBt6/4jGJjkIhyAuilTyQ2PiCVgUFNMTvz2Mth7P
Wm2mWmMQ/7pw9MaOx2MPCGbgxdV7bZlzbz8TxP/2aSHTHj/0qZ3ya4Cm0p4tjUzk
dF0vEauIIJzj6qINa16D1DmhxrGqEA6dhMjTpEV998rrJoGgWBgPdXHqB8ovNhT0
xJpyo0nYTX83nnEdQVnIo4nd7UyEKcYR0ASzICWaj9NrSdR8l0xbL0WggnXGE9QX
2nBPPxRedhXVzcS1D88AyvV2zWCwwBSMINYmYCxrJWGAHSgWv02hOW2nf7q+lVF/
i9eknYrIWeL+VlQk0MAglFCpfrSonFz/g2kGMgitABfIRMSEI6U4uHWphuP3SfmP
4G9zJH/jyDqY6KLpBDDna/xocPnwk3r8ftE/qVypdiBYUayjB0nQ4bHofUYSkrGW
yzWdOb726CNewbq4PtOt/Mm/mCoAyD3gc5mryRGuMwYiDlVQCBokl/pKfM0nAQ+1
lBnffNb68l04PzLHfb8M/PLuqKXt7EQrigvPStJWBx1UHZ/K2RtfPjBMyB02V7Bl
GhmebX95YMXaNk4MVh5l1b2TIMJZB9NO9NCBM/7V7OEN/8ZNpqJteE5c8RYrgZ5c
D0qLl07eZwwwmb+XmaEFa+3WbYzwmL46/X/Y+PlTFJtZemaGTgUq+DK4HiCqSKXc
XMHjdrqowcmaEE8PfWNjCuxF4tkJKv6CSpTDjlgI6JY5UL7k8zHMSCQE8Taud4IJ
3c7E+IKJ7lThMa1gxSDo3eHHg0wPZbOy2pxZ0djoSr2NDGS0i20TXIcz2/bJNEQ4
XvD0Ca4PAqhrAwW1n41d3omqMpzxmmuAIiHj/HpK8x4TZW3as4XFq7brMjEvBZHI
euO5g7WaiyFeiB+xzFDNAH2/ZNz6JvjCESb8EcNIyDbELLkjUuXEwWw4kCU8dcnO
6qWBun8LnDx1U3JXO9sq95lRXrPUPvi9iZxn6sMGAbhF/nA243x2lOnLwjjhzOGA
DO9HaDkjj9O2/xVozUvVciQ5SwEaUk2tGNU+JhKScr2luhrUPvsycaEwWvqD0nzM
RByGzxYhmzMKjFg4S8TgPw8i8SRuBO9SM01fvuTfwGtPUsjJzVLBe/OGkgwHeomm
ToMJq/gKsuz4B1lnS77ZuaBp3PrNkHgFFD5PWT0vAZVKrkdgqJeUF4XlMSZ3fx3B
YsXiwVfFkf4j9Omq6smtCbjuuSYJ82866y3xIdiJDrVG4WJTSiaYV2LeqircmGHk
HZLPp3vaXpP3FDLnfpG4enUrG0KfTkCJyxXaPWc8ZzCvHe3miJtu7f33/bJTNdOI
LxULHkibWq56qHuh0Zm/DzwrodM7S8D3557XiCyoIk/GpP7lYsmAOMjsCh+y8uIl
110HGAESerLbcdok5BYWNmz9J748FuyHX9tRV2hFm3TjiNHtNM8aRUtTrcIqjWTd
ObpdqdAGTZmxQqRgj10maRlXiuheRTBW6fIwS6r3Se914OS/PNRlA8Bal8dye74a
3K2QhyKqfjTEvqU4/9tSMdvj4kVzx2OomrTe2VHIaecfFlgMNQr3WZGUMz6qxRzj
h7sQMFzJ2EqnjYUEgjowM+vImd+5VvwQKClY7/k86EltR457uQeJkxj6dcE0o4i9
n11To7lahUuE/sGsk5dovEHK0TNeQuHGhmMT7N8o2HwwMFMJqSyoycjQpSlSax49
yDiTErRWEfp+dn06rjPNYODLbcxR8lvEm4YVmA/ok2FLPUfrwYYevc7Sq8DNcuWA
wkTLkgNwJXC8X20MptGHBfb5DfZ1tOtd+IWWZK3dDLe3xulNHSn7dfwmgpSxW/gn
7rVX9Skj97jskV82SVRT3wqQ8gy7XuL1W2Alv+P7YnczwvTvDYKsfx70jQOo+3Ua
8YEM7Tyk/gibnoQyWeJjV/7hw/+YHdNUgw9fMnaUyO+cKIfeS3/CdqNakBA2/q9X
H5o7WMOrNfwPpEhIk1A6zKEZU7vyOhCpPDG1HZcafk0eRRM59yFJWfAXvJfXLSrt
lsHy3xs1cY3fa3+b+kWlP34u2x2lCTOx2nWL+oNu1qPFSnZFxSq+uw6svt+G1oTG
zub7A0BQUEC3FhAJb8+8VUiaWhQoj0WPSrQ8HANV82KQrmwNExEWLf0lWGB9GyH1
kdrdLWQ4nzPNla3s3qYOKPkkkXKvRsbE0h/2aAVYblRTT2kqyhw4CJZhnXsxKJ9K
HofcOT8i3jNyAehAi5xTLVO4UcWu2Rztxj5AV6cuBwRGN/IB3abOMl25BgP0AqMG
vao0LIa6EAzjqFS2C8/OhGF7a42jyVEzSrJpoRDZsNS9lIGOEVxlV2xEbJ+Tbdj7
V18GiCtV3M4E8edAP7a1IAiiYyGScsYRkCR3ns1uHyLp1d6dBeCskoQ9aK1HDZ8u
ucIwDGL42zHWKHkmNqmpkX5Ba+sQd8WmWtL8fRALGHNCnZfBm2aPDxqgd3Zr2OM9
8qlEpUXlugYbMSxc6T+5m0FOTXrkAgMhWyrqnQiMhcuuI/FZBqnKq0yWaCIeSNgZ
W+4KyvGva/PodJr/fveeofQmEw3u4z2tT891bKRhwvhMU9Phuyeff7g5YPo4WxiT
kOr/OMdVJuWME6EC1rXdPWO5aIUwonV2dWMwoCPyeTKWkECc2jBW3+HedPjXTI79
rXOQ0wNG6JhXCIwIeHdDqoQEthCAtcbKYdyalZ2w0IBOau5oyUjby6XoZSn8IiCx
9kBmbfNEmK86hQVrq/pu1VBOqYBGkO/DUOM/nnBvh0JC81GJqnSql6HUASkiRHZ9
5alY3U3PnLpimKzbxvLClVgWx8n/aC+DkfS488uIX5z4D5mLANmVld6C0bIZm66K
5OVOsAiBwJXEx7JBu2H4D9Sbi+lY5jIGQy/AIBt3mCnN3wHbuKuZzrakiXbbGI30
xZu6hsqYhDU74ptoiGespYTApKl7vKfzsRwkYTeQN1UxqUhX5lDeiniwU7FYn8zv
nJPX8RE+VxiViyns2KukIvpWnL402sPuy4GqSo+Pnrr9P0JK/G3FQYEom4Yw3c3l
TOlUO3tpKn4IiZzd/IJa2hGUfPSOHoybVU2uSYeM2wHsG0Xt+QK5LjNv8Fx69mWm
FZsXTHR7QVuvW1oHMl44SfeFJV08P7KyhjxUCpZ0KFwN2MxBLOjVSCLA8eBx3Ijb
n9q2R6YwQEGsWxGcYwj2GYIel63Av7zAdtzBXWNI40tew0oNktiBOVc5xEYLyXUS
kqUxMgw/YHZ6T61ZCloefre5T9ros83+jvtxY/vY4NeGCZdY8sbLan6S07uq85QI
0vgDA+BrLMO1ymdn/QIXRefGj2uq3Fz4Kz8j05Rwisjs8alm1eT4VpAl5PP4+Jor
HtCUS8IEKIXw0Q+FCFJdSXe43F39HX3xJHOts3Wu+i5RbdC9sf4lY48Oa+7vZYas
U999lXSe8N2orRADc2g3C6qXkPSVdkUdv7czxoW/IcbPj/NSIcwe0EWjFFEYFJF3
60AfTm8Zi99iGUOKCzO80SMcPbtIWgREDiqWCnnzt8sg/ZPBXr9Cjyi0MeTSRg8D
XRuun2ju/spIJH2tNIsbez/YQPodlMrnDW62FbTtgtQWeQyDnqFlaN+aAaLR/Qa7
ZLYY8FIZzQC5VUu61VY71V+GvBzZZ/IPUReceSIFBIOufSfTfEuJBRje26m9s2wi
o+Zcs0WHTUwFYLUvyERopuhtZ6luLl4vCKwwml4u4+Bb912XFQETUAPDj7safSzv
C7MfG6R0cuh48qEuHzB+biqmNosPMJEMHgOaAiqxtVHQ9c1yYPkBgqg955jXRaJ4
7UbP+7PMxrvl/zdkmAxjfltVYcKAMo2rcREgJt2WFmSiKm49JCzovqmK5WnZjceu
bpaWlpu3Keb5K/PMw7MrHy89drOfhMbj4KhB/5qY8QTI2w+o3DMeNwMzHI31yjbC
TUmf1BFIP7S6W2mqVbTx2DVNWi5z74dXRGrswCOGaA1lmSOgtL6XBgT9AB7tH5XT
XCwkWTI+rhPJW8FnMhryqQNwavMrbhR2j/WjeFEMDTqnO+xuqhqfflv8jg8fcYJB
E0J931fmNFQ7KxjqvcnuQ9RUYCM6qKIhWnFVCuK1POrpu1vfscwEAYI6yE7QFFco
CyKejygfS/WLRcvcfZQBKq0QdSn0fkPJW+CLrCcXYxXbCdF7ebdkEcMdnobUSc8X
uuE61sjBKK8Ahwl+U5quqICz2c6keEw5RBSejZMsidCa/p88fjv/itRql4RSdo5U
1WWgH+ZbKB3m9Iobi7RXYeyksjD2hRab0+okgGHVLkzgMFu6zPR7+ouANPO2evhS
y2nk7AkIUVhKfqOwo2qojR1rzQza4x1Woxs+lNXAwX9M910LBlc5FZcOz9nVDQaN
fIRa7sIKJc+qVpLjU3vH71m6BrJYguDAHOUsgnV6YeOhcbEwkUa5zjvLKfkjjjHT
myyHNuG1/vj5MGO3NuyO0IM8wYRG6oz6Wayb7bB76mx4y/tozr4oZdcmP+qB5YR+
4z5xYgsVcqmoVg+bLXpjLdFQ+8w77YVdf5syN4aUjYX9inNs8TrIG232hN9eM3Qo
RC5ZgwamDZlHy2DDQFmV7vIWO1oRT0Qky8msv41D8m3n8G75tlfES2zChP/rhvEG
10S/URapCdA6RLlSczzTOK9LZfcj6hup/PyM/2NMfVQ2IqQVxu99GhCLBny/5k77
ZqTTCT5sbaPk439FllybOgdDH64pX8A6KMrUwylHpzWEjcDaniaOwdPKJspAK4IE
hXx1UcNknsRSaz9k3ziVbdMtLqWfCtItMfSLXeV5LSd0SJBkmLPujXPAl4UCqH/Y
65tWSBBcmRKXshgmhGtprsXpt3/bjFxTvikNYOmRMK0mC1KmbC6VMaMWrpJG33Ii
XjfQjnuQ63V2UXKUblDzWO9BP029mlsjq+VnVVyMFc8/QXpPEVaxnodY62K+zKZg
/mFGM7Bw5h07p/WT5s1EIr1kGffhZQvmR95eHTRocE09fxGzmgtjmXqm/tAKhDRl
2rw4rLsoHa4PIr712gFmXkCa8JG6Jes634hniNYpXJypVEb+YHq6e1nxTeXfh0pE
GrL1LsGkuutB2DcgXvbnJsntbKO4nDIR3Bi8H4FhzKXmJzIfMC7rynZwciYpDZop
wc03KEFn7RTvd+ScAJE/vD/fnTz7tpFlZytlk8RzD+DfL2ECN+lwrUB3SX8E2XMU
YR2GDuuFCOCmdzaEQj7nzOmiQ57RdFLT02JQFIh3Du3xuLSNRuLxAXLDXczUJLze
ylZQfPFUwNVCxFuCksRUNbjzwNNHYEnupecgMDJIf2xWCCAKE/FUx2VzG60qJAQ3
3m3CAaEeTHrqjYp93WrF52lDg6xiZHoKKYfJzdS5G0w1OxbHg4FB3H1HzmZEDIkv
MUW8xnrMJesc++UOoHzoPVw9fsgplzGiedHRan5Dnx3vw0BLISRKgJmc8fCJrdDb
gW5pvYpWfhZZsWAZXcmPwTK8tuf7kBHmOtOdqJopVZUmJFD3pd88/rH6Bm6yD3cc
nW4NuhfoJcax6LhLSD5Go/cjxJK5KeRx+/iSgxlXA9OLqDho6dphiWu5J6BvzBak
oQObeIZ/R71WueXxOEBgzQW/utBRIIC/ErOxGYxDZkP1lJgotqp1PPGsF4yuorOj
FasOxKfoe+dUOaz7o9wn/GpFHE5/s9yItE8OQ7IL0y8DUhByFTBrEVfvYZ9Eq1ob
w7KGJGDHvsiooGKl7i1yfK7f/VvkqWlAU9hRnz3u719rcAjNQwShAq1PPY5d4G/5
qX56sffvzk/3oRnwo6cRSPiXeOaYJaDws4Jc/PgtyPYl6cSGFcoeUFMYzjmulbW2
sHJQn74BK/mdUQT5f4OFM9qo0pEj6TV2reFMKpjkgGe9mCzi1Xyx9k7oG8pofY1t
2JuB1mZof8axcKtlIg2FGaBmBqCoXR0pbNV797hpLK2hlfTxJ21etplTRGUE8T5Q
G9KBCZx5XK8RxmYUq4bPJS5/PyHLmoTcVzNNgYrsPfQJPrt0ya1J3Lv2ac4i5zkQ
9TVAFLjOa0nDGwTitM63VYWOgJX+mwdoFeGCMpg8EjBvNhuMfFQ73l5UgmXtyzMK
RVzWOy0GEuv+v5zygJAmGBvqDf+zakgWyMBVzctoO6ZChi8kG/EJz48gvB+8nAUh
/CSjY69HazQvz0WaMral50nLSNL+59OFhAOb9QZLqyBnsw+oRJSG33zBMkMUpzlP
uj0W/EKwcn3v5U3c4DaqfJqS1q/PFaStwXhms5ruK/8GjnNnaiXoN33leV+nxHOE
/scpV4/tK8C/7h+OqthECPCMZF9mAfYPwiYdTv+DvfXwyQMwJLHRmLJfyDVn3WJi
OvEXvqcGGgeTEZNAygWMpxNsgFigG9cUQoV0Z89jXLLXV5sQ+Pjr9PCeEMeuIrci
uhivKUw99jp3nmT8fQPngj3l41NI2gDMjphdW3DJYMLR3XpaYaFQoy2Cs0MvOsXA
Id2zFmX23uGwhZFMWe+M+/+JjReZpezPfpB8GHkvCyfeELETaJELSZAOjKscFiUf
+dJPwUF7QfbFXKvT2BvAD+TF8Rl9TKFuiJuJ+bY0n/TPkWrZ6pFOMP2qlhbXtQyo
woqiT7s1C6AQojRzWY3FUSOdEjiwTUGNc1v8PB2yxrJh4EvGZAMR1kQ9VvjAOB12
FPJi7rKPKDQPPzYv5SeGOx/gtMibYHJhGwL8tvmJJ28WSV5cHlD0PEo0hzJnyNdN
EGNCw06SUh4oLjbWLnIcMPnObz2YYzdrjd9b1fPz1uqK8LL20/iXfLUSRZkTskTg
IcrsghKhZe2LyCXRXhNbagr63CaTF8SUhukJ7L4CEq7IoWbvAkBXywhj2EbT0poE
x/MGx2uOrlFKoXIswu59LLv0ZW+oBfB0IVy+EK5fRGrEJ2cSOKo/IDybwmem3yf3
31+VZO5D1p7GIatWhAy/ZEUHoujAm/k8PEw03bQf+v1KThYnFu2aoWJcm5B8avCN
5uZWcRl3TRVlCsv1HjFGEDu2vdePKIqJI/4Up9XipnSXYAFDVo2AqT42t9/mj7zc
4sc/Kucc3FoTtp6pa15OfdKPDhaSK36WKBjfJGULDa5sDwDYKlkFKH4gaZN+0IYP
coe5RrXjQKWdacKOr2IJL1aNjN1zLUoohAWFsv2Ae+lV/xTBo9NrTszDjXzyBiCZ
+4q91oYsuta6tD2rl94+tzqrIX0bLTCnoHjcbcod4CJHPr/C/XGyegkbVdiiBpku
FzYPSsAgTDsqMZdMHtz7yIkZMK2i3wqa+PVkUF7EiuzCilUQA7gRa0O63mbNbYkm
uI2nWZioH4vbJnRtB8HSbMoBUcwsS6mZG8v2ofz/Xsm4YM5oDoi2TYZQMUzRUio9
ARsDvell6It9dJcziixnlRVGEU5naWvw4kOopbERpSCpFaxUrBfjzZwGZvGAZO/X
YfBVfvmVsW05gR5S/oX0D+zWhogNqcwDdhipdYWEee2vDDg9lDBaUn1t/zj77eC2
9od3szankdEOLVwMujqaIh3z0IUqn94GcWVgWoyqeoZxLMWgkqicSHYjNKT6x/iW
NqiZj+rTtrEW4RNGM7FPIA8rpnqoFmbR2pDT2rTJ/+RGWL66nWjUQF4FtSUTJp2U
a4uxJ6rtyA6QCzcJ6whF/o9/cjNF0ZNqBD0XR19IdMLvKcMwPa1uzfOlIYzbjtbA
uqna3hLSg/SO2wlQbBDjdDIR48QG9wtpdnzLFvS6O/+GyShfLGAsUURy2bDBZY8v
X0lMsSmKHxuc1YwElpUjTKVYpzVZzramrIwvr2jH71e7+Cs+FnVpudQRYWimD+4Y
e2vcG6bE8zf7aQf1oPhUr3PlzAHDybTLPo7Ds1uj0MuZCe5KHW8WMIzM3o2eW8fR
M0di64dZoKf9ZsGfQ5T18gUsNWbjfbmZAn9edAF0qjsbIjZ7cpe3iW6UQ9LNLAWr
F6CWnM6CCN0lUaPN9niJfvRW11Zv8oLnYgAXcUxHqY+vs+zGNbULCrLbjJwFnUz9
BLVd50u95TeVQo7uVmgPgm3RlHpdhZRiintl8YGwUq/k84VzWhWTxzCJcljZ/V8q
gObAjE/046tUvcM9IzkSga8QUP2YBQzKcOSpDO0zFet3/SNJnPwuSXIyurRcNweI
CgLdE/6UuYxBcLvHdlFaEdp8XMj3fYQOS25WGgMi+PCpId8+nNutPyzsWY6Ej61N
/Lw606YmFnNPIaXxToPo/Zdq4+PXgH3r4sUcgDxALN30SqAOGFncdPugzKzyS0O+
zyqXtXbfxRcOdCBg0aza4YjPt341MNrtw09x45O2lh9ZFRSmO3bZgdN8wQ90o3uF
stQ0sWzTcC3iv+PVdyoaAlUse/mItyy3w9Xse5rWtwjTGg2+eFah/kUf2cFkGIad
Xdl8xAvDM8JWz/yk0WijaqcBVQCaLeAUe9xPrUSkZPjHPhZw1lzDEJfFcvYXe1CA
QauuYcYWZHQIAad8x7q6VPv47iXlJym6zyoRqHKAXF0ILgd+S1q4cPFEKIfdqRC8
4y5eGR7mXOJw6UdkKlfPZo8VuYYBPpL5r+tfy8RXiE8Yaotjl2B9oEdoGYPwJ7FJ
s7ylLy9+cNuMW2f8rPm87h7WYnUH+uokiKYnTAFB5FWTV4pK4Wypfo9ip+iWoVtk
G77oWgqVPTIjOxsc/46SO322iLc7Sh2XtYecIh9BZGZMPhZjqeYoyF6qGWRTvl+q
YhoYdrLjJCTJJ4VCSQmHUg54Hz0Nxr5RukUbF3lRL4DpeAh8X3nZsMLpZfS62oYG
55nYkv+lxVUHz/6Hm0bEOzRbJlAP3ShKZssiJNifm8fqdfBk16pgai0bAub+CgPb
FMw6GHycwaiNRjmumbtHUzthGjKayHof4/gBspqNtw8SdGpUikonhclPsXap0sNR
Qai3VoEpr3E1iQXHstvLBLOhs1zmuVbbQBlxphAuu4ByNemgYil4fnCfgkxnLLS9
CSwZoODWIh9gcwKP4P8SlEeI6iGdEfc8ibR3T927I44MAIczzH0oeuqxn/arzKgn
hjg1b0en+i+0ejTK5N4zjtruiDgEzOpMCfXrfypVTJOS5eyhuuFIdCOL4CNEHB8z
gzpEB/pLqeqFEoqhFtrOH33yHWQnAsMKZZjOYVVymqZlRNB6YxWM/7kGNAZvmChT
1L6EgN3siWyh8akfP/9z4nJIKV8WCkqaAvK4pM7IBOsPiwv9H6Y6RKLSRBeNWlIs
1mtnMbXOVyVdSmHhpyf0XGtChtLC7tlZDYxsQL2xMOGzW3n6MW/HKp8u3jWXgFB7
mzh+rEmKyDYVQEmCOtAOioDrrJfxKF21sfkgkCavGFXd2qhALcElRDbZnPFTsQXv
Zcjlp9Na7+xUGRRBFS6EDQX+Kv0LFVzCHbs6hj86CP8FHv2gtBg8GstkHwrSeG7f
f40fio9h91QezfPtLEoL8SN6xYf9xr9FfQtL7lv8Qv5AT4Zq4q0Lv1pckxQo+ISa
/Kn1IV8afvkdqaynLzSRto2/sP1BAKsO9stWaRyMHsIHowFnY2OoCxduofEbh3Du
ZjZg9MJO/pvLOqnatjdv8FaTvY8odYatMdXr17sACXbsMISi3UuJNW4K3dHDySFn
XsF83BYcdHuw2BrvDCttG/vs4Paizf7zwOHEHNWPRBmVZSC1QBxOeW8wblpk14T7
9Z+nKBKto+yKCmsDY6rDUzv7Ii90OzaSnS7oSbUzVltKUwiPkYfEMk8+E58s0flM
Gz3Qkvn/qRGqAhm7kA7KopUUBZpPXcSVaCOs/EQ66Pg/RJ1RtnCKKyAT3hLQRQth
gTkXwwHfjk4FkUOFVbQWOI03URE/BrM0mzBPkMSgl8daHEGF7Az5+a3fe72xUSqU
56b6sRBgrjKzSloUDGWbM4Y+1VDxgyvyKh1t8K6kQIWp8cZGUto/JA0QVMBQKTHL
OCnlQbqHaVB71DZR284wTFXeGPe/Yj0A4cc/KLuE6k9sqR/unvN5XrlY2Fpa1CqO
ZODyuc313te46qWFx0TZ0lRpfxsZb2jNNHHC0g5gi5wFqdrNQDK1BZ+M1ZT2SdNK
A5Hcvc9whaokX4Zrbo/g5CCoEKxFPQadveTWNSP00+fDs0g8knPQsniOJR17zlBO
QIoY5lBm9LkYwX0pSRDVkT3Fya/D/IsgMcPlETE+116ujGCNjNdnyY4M0IFldq41
qRUhSyWfVi6WcMsGujXz3ATQxQxxxY2mt5TjTkfzi8OddWerYb106xJPNIKqqjKP
JUq56wWj3uzSx+81P3YBDLlOV6yV3FewueM+velQx9uLbL6hG+RG1SdfEf74TW0W
PV+Q8Yb3B/5Z4BjhFecYNPesUJ/rPsiyxxm6BlZtEqsLJ9hYJ8nPNflQZsY3Sxg5
5M6sIC9mbAjIgyCF5LgREwu2Qjk5BM+/yrQMfEo/+Xnz/8UTdErduME5nVlXD4KR
rcd+1vUxcQBhC59tx2O0aKW0fj8tUwV3G7N3lGGuvIdTU9TTRc9r8P2t1VMcutCB
KxLLA91Osk4OXcy401SPsFxxM+/g5Pk5cLr5qWAS8Y0HLexOsiSjfBAPU20bBTRd
R1gJAFSA/tyrJwQofAyvbWIwlmAe85dSenA12Ug32CXt1stjzzeIybVFF/lPPnfY
fPaYJ9LNFt4wx/i5SLGzbPdDPln+BuZD0uXGJ47n/tf3B0YP0FtvWUbLRp9beRZt
CGx+CiRxbP5OjeNt2qEAlz2xYJSXpwYgrCEzNX5mTK92bNjoK6wn1Gq3kdDtVPxi
t+hBnsK7A6ytyKho2RG88xDm4OnpnuiInmdoFXJ8bS0hiwrMtuooR4PVFEpvDKKL
bbCp0ni69i/+T9EpQIXo6wbhqGOslbROxffNNtTRgx7sYlwT+vpaPJF6a/Lhhw/m
l6AOP40t7M8Bh/tYTBMlK/pFlFVwQYpvzQy9ftK/6aAzcAQQtDZFTszARb9dTdqn
D5Zsb7q8d4IUHQBn3xnYqq1JYtcu+pepz2hljaua/fJBfewEGwQrDcf3GJV48rO6
9gbh4v9DRVA+cPavsBh/BLsvxtKmrHSkzV03TZ4it95KjRpt280ooocUOUfFQwJr
KyQBHiGDO6PIiYVXRu+iTzwvMA0YFqNkZZyg9nUydZlIbiGofIRt+oxgYRizwk+u
XKcrVILWbOaSX0nmDGQ5pjBpBdTJON7kdHhDeAuJwuKpGD+XapWtopQ2ymbNOWW6
6QYCAbyntfSBjgDBWbml4QeVPYryj1DBY0o+sPwD//3y0jB+WhgYPWkuiV2RrlzO
TmFnXDSCKJnAbF9uwEcuLNgRod3f4o0O/s2T/pKjhtjEgqD3FdnGJmQqr2xt0Teg
Ez+o/Bn8gIe9XFX8q9eWx4R8IcRCWZLbnboqhX2tTgI6fX314YloQulpnurK5nWq
iPkQ7Y8FLLUyQq2xFNeyZ7uJrRPenyZgOfadqqtsJuIH/VtPWRqNSY2M4mCwpmr2
VYjkbjERk274dzfdQy/MFZnRmS0iBXeAS/iIRVEQxgU9LF202dGyvbuQEBjKA1w3
Z7JdZ72xrYwFU6OL34HpOzrujwr6Qqqv+UNNBy1FLi0Xu1/lB+ceWk8yr+o/lpEl
9am3YjJI3ZCkp/iPURdT7a7D0cxG10RadamPew6uvKmyFwm79RSF3h5xy4CqFQGI
roMuyGLTVlvmAHQ8onraanuONI9/FxGxc2rL+M+tAtA+/WCdxEK7ZAkR+AFcKHYj
XSnt/nucbGpTo64afDjtoMrpr+CMX0CmmQdwRnnPp0pVeF8pQS5YV/bf6pG5ksTT
ZqozL0SW9Z+wKZSWjlC0lIQOr9pHONEr+A4mTr4D3EM2PHGPNcH/s86+Lo3fIbpo
WNHG/nN5KDmd4JRUK0gk0xPZgACLOf7sxg7Od4OSgMRvKVtNIOPAAjb0oiaRj3JD
uWFOvIU96uBwgQbvMduP1qGjRhG6+yOViBfNvRWXJJ6lPDtjIQk13E0wRlrOUucO
iLZdCaPwfImkx5VNsvRmWoLV0ZS1Q6W30gzp33DgGRNsjxNOpqGOIaFD11ljP2UU
NQAAPG/KKhGyavMM3/oZ7/lxWISWdQr9b1N5P/ouN+iTRhzMnx/qShIynx/3GuRa
eqsVYf2atE9Kh6xOwGlWypWKVJAM99zCI59SToBjrOczRqYg7qz3EyG/pbYg8LKF
8puiw7OM5jBtxK2OC42z2zqSAW9WgekfzjZx6eGuJvL9ffkspyxhzYseTUAhA/tw
4y740+r5S/no2rW8x5G4evfphPHhOxmUOXdH2JZVwo4RGSApbIqpWXeOvB/jbmBg
lxx7ABQSPi+4CKmcQydZABV7EVj7WNaavH++qfwz6Uak4+eI7WlvH/UjDZCw7qeA
jKrqmnagMu8bwsvdINT7yuhwiZo3jhOZ1KpDS5iVQo6mB/ot6QSMd0PbVUO/MGZO
MMdIj4OELkVYMi4Xf1WSsRYCw3lnWGnXKhneEo7NsO0D/EumlFbJANloUVt0kY5Y
VMxsYb652thKWtF8ZRpBAR77eGf2Y3Pcr/UpuAQRn74gQcAnfZ6cxSLRfLj3G44f
Czp4aZ0QCcSKaKDfbvd+chWAhEn2eIMjh9J5Psl87Q65iY4/Rn8aCEDu3VrGeEZi
cvmXAkFL9n/RjDuHI9HDHzaFyt51B5wHw5bfpgGdi2nQUkBhotVvn2PTO8NDxb2Y
vmkcuCnXhTxTG0UsaiQeNhM2tWiS2NeNY/W3gjvYlcUHdVccpkjKUcjl4QLg/dR0
HsYalEin9zuO1luTOs75L1LTsctwQpibNRgBosFA7q6r7mG5BQ733rymAIeGI0wF
GApXjdiIlepQFjVBfVWDzHqi2E+E2YMvHRg5U4PWEjwGtNB9QsrmlJay/qmU1/1R
6HlV4IokKutq/RkJOoiH4GtYTrZqIZqExFWtEv2vMJG/K9/koO8sIkIRUuPLKUJd
R3sdcFHAJyD2dw7+xmyLTschMfWed9fD7qk8gbD/oPAd6FIWYx8m6iFZW08nYCdE
dpq35IeB1z/2rQkKp6ButpQ29APURSf5oRFP36fMojnAn2dJzPq7cIqfnvoF6Y8p
3w7/gz5A/4y9BjaG3565zaVJXZzE6jCPCrkPb3IiRy9wDopWHaKQYoJXgl6SlJSC
h2QjkjpJvauUvQG+Or9fIx1GL5U6dLrXyH3eRLv0IX8AEw2epdamGlM0FDZtsNxv
7hJfTGW6ECw5ej1bih4cdjNhzrRQ5jbwy47CYeQ3PesfzqJbBWAaaTBjBJBGrIbr
27o0vnQFqHeJLQa+Mh3t0sADmv7K7mTAQ7UVwui1KLBVCpoAH4IVknSYI/WdWyrJ
v1MSZOFk1wsJ2yZUaGQdAR+4m8IZV/thLa3nQiSAbWQo0CaFpoHX+P8D/pGwPhxO
R5ZWQgOQxoubiUreGqNlk9Ip+DMXWMz6ujZgjZMYc0ifAFDTk97K9iU08IN5uR4R
n0rRm0WJF0zps0VrPnkhKpbmITxc//8mx+fEIUSvByHk9DQ2feQTjn7/irtTGqVU
K6BRy7VJwOkPRc3xPZXhsbxuS/TVS3WUYJRTMZscNrqCnKCHJ2eq9qMOXV3Y5BGr
3yO9ZeQ8+iQnjbsVgYPiGRNfV/3V49pxBpF/efYT3MNJRiaZjnwd2HWWGL0zkttQ
HCz4Hvw1ihj/IlS+lx/dcXRM1P7HLLUF35yZebc97oOP6MAU8Wf4qG1knKVH7GIT
8PwzFrth0dgR8UFXWeeKOB7F/ABRit0rQqcqIQVe1W9QcQTw68pnFQfT/F5b4Ehb
ybtv/JH1WPlPVMgYWCOmHqJktnvS236pHh8GgfG5J+wu4LNlzqg1/vwGNwiv0J2Q
kcF6r/3p6JJhN73SSkZsI23IfJvjjjgIZsz0LdmWeoIHhQyzuhZapmfhOweWDzWp
m3QplWVKQdZikwHR5bKzjPSGpedBqvjNPtDvxnAIvB+OnBkW2pjWVYPFT5ug4stD
fMUu+E8XW2iAB85m3+1wcR0HZrpyOexDaXywpJrP/isa8pFxdlMR6Uo2lKR9866L
B39SOr2EI6EXoz9Rowq6iP+i/d+swmnIh3FzKVs/hfgKAIauMPopmBLV2V5Pb6TQ
OKTIDpZjP3bmfAQN0Spysp0AWdBvE/i4+5OCqTA62CSQdf2GW6E5LZCSylyhasj/
XV2QHr8dt+DoDnSgqBVSKYxaBe6vANQaW8hbdo7I5QCTEWNklzMRY/FXEkEvCkGE
Q2e/QjoRo8vtNIsI06iFyD+8jioJTBgBqSqw42N7jRBW61ILQCn9GB+GkH+8akAG
s3AsosoZ5+EksrYY2KABw7kR1kRNn0ftA7TH6OQS6xmfNUsINLD6bLRa0wOFmJ/J
zFeGfruWeH/PRnvy+pjY0LFklxeJzKvFE5oEDByhR18MFWQNpo0sALnkdYB05ic+
GDrkF77AngyTqae6KSl9wBsO4Ai9IDghnoky8/m5Wmlgm0c1U/DBfmu6RX+VMS5J
N8mnr40kAbG44eaYj65Lw64f90TEL2o+jKIy/1h29miujTtLubpMpSSL/e9OH9x1
bc+3hjwmCBkRtotj2TZSw2DoJc1ZJxonbWwjJUxP5SRH4XX64jI9/yvFRE0GvqVB
ejJX/nBSCTr2wKJPafX5VehXItD+rbm58qqGTtk4EHCCsL8wv6EW3TaKbG24IAFJ
rR/wWvdRAy9BVQivM4ndfC32/NY003kZfbVvw72y4cToMt/vBPKX9RFB9Bk+v1TD
DNfwmaDVyg/V8QWaTuiObU/cGDN4nmFbzd7AEXms6P8M646kTzlpAUMBpDu+C+yj
kbmOi4I1z9KWatftf/p/oa5eiFhmV8wGWFdR/cTgDXKP+/aKk/xEPqInSocRA//X
6OiPX7IeyVAU6r5GdNRspkgJHp6+gfq7SHSYOKE4wWiE7fNoWQYynGVeYfoqA1Xu
yjRGHvcDSg5BxgNJdXiD0F87k1lWSH/G56cZXW+n7a72YqHKr5Y7Y20rHSGaHH8s
UyjSxk+3Gkro1IyOsF2o9FEJEOPausFOCrj7TnApJzI5kw5do2CPvImtWY2uwGGy
7luQi3Ownhl5Nt07EjIdt960vJFcStbKQHeDzxaFCXapucVlr4ssPRZda9WU8AU4
EKwMFnx+zXAIjlWLYcYI0kFQvG1mh6daiPQmoT4LxqlJ5QRTx9kwx+VG8V1/nHm5
8HvoiPpp12SICwPgoykvEryYmTuWwoHW7j2i3hLSBvqdXacfKUcnTcbl9dSPolRK
QB1CJupxPq22NxsuAMjI0TC7lPbeAdIM7q40OS8xdgzJAH2y/2yHtw+XVTftL752
cXobtYyWVYswT6QN8gXUC5Azr/q4vzNjyl0YXkWUL3CBk2tC/eAlnfAulbGl/jlk
oOm+oXx3xmzXo56cGBM7uIMUqIOGIDgSvHj034f0VdQ2M8xF7wAFl+msCZ1tE1/B
DNVmYVInJ5AanAzl1BpR7DHESb5ZiAKjOBXznVRlLKiTv74yDohoqVpmRlHPTmvU
exKPj52VU+KvzHDU4zUINcXPmc4D7b2kIqXqBB+e3uYMgFuxn/XMiwUlk0nghega
XjiRXrHfk0Qb3xeWPYvSfqL0zSIvtFbOkIeeVWRdt0hlHzT9J/Wz9dJmJ30WRLRC
R4bVDsU+fV6UT4DHx4tnfiLpL5PM5f4RE5uIooK8jqLh5tf/kFGPL0XqS8bMzrpR
Y7lDkIFcqcMTy+oA1MeDZdQWmqku1RRiR/3h57U5vFI57nmZOWwoVCHF1GFPs90c
8jwWIeurCRZuQxlPUeKyqhrXejC78AB6v+g2S2dkHi8qZM7dEyh5m3bT5aQjHzbh
vqbD9cQn5BuiFDv0xucnDJs7wk4FWWLfEzV+sidOnB6VhXBtonvKi0FRP9lmA5L7
tZpHwFZIJb84ygn4HvPQ505z/iH8OepRGi8ApN3nnUO9UA8qKkQ5KiuJpJTSctKT
KXtQp/6q1+m+nqwieZp2lVwaguwsdBB7QojH8mEG2xDTj9XPMckMyvqaU7C5t+T2
lyJW3deQaiOGD0mPeoIDZqnn9t3A8qM1OpH6yqpm+jqO7+KMf4CFE1y39Iwgp2c/
vnUM4o4dIgnS1FUKOd2RSMEus5u97qXBvkKs0RH8GAKLwEfYGQnesqJYUjKLmr8u
/NPf95kAKpv/5QHRyT/VxMb8p0Nw1aPYcoR+1BFHOZiJJM0WSMiIRtCowQrppuIk
v9R0o8KoMyLwbjCReNkRpBJZxyW4F18MUHHbkbXMQbUKu2yPs7/BCY+jDBjR2VoT
AUvejNm0IntcdjetAupMO5E1wzw3yOTPO9KcxQNPkw36b5VCQTrfUe1KMPRhat/S
gUT49w2BHwAj5LcA7wyvPalBJbx2nRccJkdHEEWeBf34AhTAReXgHeFigL+emjQD
xL09rYoe/Fb+ZJ063vmfOs9kwpd6/qSEHk5PPuLmuzoAMIj5CLD4717m8LG03Cq9
CeLjkx9myzGAqXje/AhjORPtfeDD9TR85kWEzFs+htBid8wIZfOkWx9LgDIkuhUk
d20Esni3/VLS+6lHcglN5BIMDXpoUn6KGxEsIpSwbR5KHhsYeiWOvkPPV/06Cc9/
7lbUqB3L2meu05QgVC06koE7esa5sLQRT+dI5jUNzdnosqNlo4vIlhe9gu996kKq
DsgL5YpyZABJULRQOiqEaC4tcq76xHls7yFT8kgz2eMQ6DSzVqbDSv16gUyDtfwt
fQsB5AL+79GURE+TLn/YwI+R50uHDFG+dFN0qkjIIdt8C4Wc9XyU0p7l81Ww5WuK
E6SR8Wx5GB7jMvMhKFIhD/z2ar6vvJlvSFdhAkccEaRInweRS/bXqEbwWv9c5EtR
KH9kYb9xxqAk5Tva2XKIjuXqQ9nauvur+GpEg+LfxO4q9ZYLXoF3dUYt0+ZAlJy/
Ob+wDv2KjeMoNQ2TsAFhHy1A3z3C9RJXHPUegEEwCiBVLMcw2OtzTJSN4w0ZhIrY
xKjarcxH1BLm/O55nKgxJ0nlyuzSY3cIYG7PJS1kkWS6BhC764Wr0u62pk/5wFFi
zFDFkD4j0gyGUloZLidVdtGNRVjWfD+kHcSIxICEq7bKAQ6D9Q3TTtRnw9LZgPho
T4O/msUmCl63pjalHfRC+RuRKiSFxNXY0ejmeqNBJuvqtDJGWtrjImRS5zaSk4g9
BTrUVK00zquKRXYVyZvSmhzfTTlF87pUTEo38tRBCDIZMR2L3Ks95wg8uqgamIZY
lH84Ypeq98zFFfaySn94GmxEq2R5wGAjDL9DDUgwN6ModFx6MChbmDk2QsPWkW1K
r1qNmrtnb7Jgl4eiV93yzqgfH9kYxH1P/QueyKixR7E5ndIOPcvDdTCoixYkCvl4
4p3UnnGNkaA5MYwFx5UnB3kw5zepRvWLVpVD8k6n3qugFw/iArat4/36h6ttahYq
83HvsMVFge4671taqiUlv/bVfnbdJe5WXQYqQi+rVZ0G3tnOizOc0oPQnzhDh+L7
k0moHtwDbmB2eogCbBqfyFXahRt4my8mF+HUlYAIb1zMlyNkyVsrLkGId/RBUtL9
NZoOpMIscHCFCNWL8oIrIia61I+SYhBg2ssi6fWaXfdze17H8caPf3xw94SMHSEl
utCtqBbLW8jXCJE9QH8Xlzl7vq2ZrXtPWJp3cLr0sywLfKzp9CwbOowDfvLGDiDF
0c8CN1D0z8qEmS0r7RCu65+UH7shUTCtLLGtMikTfl/LnmXhu2CtMl89hC6Cthxf
wd+3PnQiPv2UFNAU8VJ+K6cvGkzdg/zuHn0YQ6Df0SMTWkJGghHa9PAIZ4EpJ73C
Nh46mXAA6d9nFqErGgxxPCVylXwakUbX8GGPvg06AiB2f3885JgH7hXHPjPQNl+V
YHD5lYp8kKlqwPwLHvvOGzdLizwVeEPIY5xNEN2Twt7nKcOjWRIKLSkcPfdBtgYe
s4pkGbR/ulR/cnG/XZ1X73rdBwZ7s0iTS9e//DelLYNukLmfLxApk9kTxaXHLoH+
j8nplaXVh4wKl9mW4CPB4Bm9Ya4bVXFSKwhVeokN+EBTyqtDkraqI/ahZVFDgnlY
7WcZ/iCoKXke9zgv38ozB2b5sNUKBXB2V1VhLjlhaORkVxof1aRWm0VRbrnBFf+m
/de578fLzzpxf1WaBChc990oomgLhy0vHTqmrMDY+b7McneG3IPr966IjkL5XKzY
HntUiZ+Uvgdiq8OvxlftvYzo2nes+0IQBNfUuoOOibjdzTv+Qh6jdgXX/UZQ1oQH
FSqbQcjiaeqrR6XeC9ZlltSxEcSyzwoeXMe74cXOPTHmSih5mk6Y216ixG7I6J6m
SRYpTnLYeyWi8MRGMDxuB9qkAnTkULyzd/SRN66YqTiCCCWoG/KcOphknYPvUHPI
9VyYVpGnQi9haAkq38cPdkU2faL529IMwEzEJfaF2L8Ha74aisamUiCzJT+Fu0tf
TqTqpEKi9rYUXNl9cRuAOTKFfbP3JJlqPmnrLjTIoy7dwS5Um4nitUkAkVOAtHAj
HDrcH/530LMMIjWLc0MQapNkmEyEI+rbkedXJdO5eF1Ao5lkzYS55zz2MyUY10dk
EobSB0wnMUToI6OWXHkffitJEdsNyPJWZ+9z8skVZBbah46jvo9a5WvNRNCz5aOs
8Li6tmBSQmIjL4NxQGllmfbMURBBlrWyLfnXg1DJEg80jceH+cDbS7R6b716CxjL
Q91BugTNmUaMPzbeb5oRk7GJ4hG9InW6L4gdXCIFp1cIhf00z5nL7O5g3duo5LM4
zcOYM5kRT9Eqc4eq++otujWhvj6dXSNVE/ezujxW83dO5NQHoIeojBi6ITm5DPQf
eOXpJPkSCFtDgnujSaQNJ2EJiBC5U9QuUUyi2pZDI2wjsr0MJwfBDVk4N7HgSIRY
5BSpPHRz4N9Ekg8P0KiDd+ZgO4XyjJL+HDvv+SolbDszY7eP2YnYBbmjvhYVxXfU
QggMO+//KM6vL8hjMCJdul9l5U/S8hTOddyHFeOkh9Ae89GzNu8QpTEBd9BJrqYr
cbKJIFvE5s/ejRltBIED+x/y5RJ/MvetUJ14qpMxUB44hAGd1CSftq/TYPbfK3ZY
Gqic9wG8BSSDVuOkKyj0a3yOcg3Qh4XxNitu//ZhWBPY619Yzqbm/Ao5rOXrKF7w
rtbpTx7WwXgi0nLKX1W/gQyXYqisQz9szkKMUm09MSMzHLx+8wL8KToOtl6qltqj
jqpT7c9PoQEspspmFoOQ7tjkyWWagaC8Hfwo7A7r1V291E0xKEx0o6unGnZ9E/8o
z6u2yq85cer5IICYSUE/lm/Vc7puvGsJCfPeN/YC1Vx0ie24NnMCh3DI/OKS01bW
HKZrzjpKFidjqmaa2nQCW7BOaMM+UkFJG8acJAxTsKwFzFgT1yzkDaJdgBH9RGF7
F/fCpcJ4jTNpepRTXsjqZQXFstlH5BIlcqDQQQHYOVRwbKVTar4Y6dD20+E0X67V
fcLVM4s6AXwZOaKDekqxuE4IdxNBUE7lwB+ikH+Tps9EcwwL8ZLUjkIIWzFsi89x
hqyVRE4AGDwuGIW7wV9FAYJYSfHJfhG/VH/o0PuwfbfL3pN3mYbNTT+wWvIcr8z6
oYtjj9mA7mtVCwOWtbz+POGIOJs+XeO/ksWdalvGCNo6X88o24J/LN1hKAEBMh05
aMaQgH1bFSTJ7vmHttDq92DAQC7WDcYatX7V5h5PnaEwTrkXFUjvW/p4YN5FB4qK
xVRRbMiSVwOvYPsl5LS17x7Vb8Cjt0KTRmUgKMfE0Q27cgdKHBL8KdTKmGLtw/OF
tj/W9MG1CQbwPKy0glbsiyHeC76o00hWxVT6Zc3ucLl5FK//ZTheK/GoDTWBeJbt
b4e96IdzONuhxTqHJt2AigNGyWsjiZ+ivuTUc8pCrLv61s1N5p6FVmuBUPcd6/MP
uLptVlGNhcT5TYgs1oMZeEc0Y6De6+hDczeBHfg4+IunzPcw0xOvs9RI+/lTvWVD
LyN77ceOxLZ7/0oEQwmaEM0B6T2rfxo5Y96JAk6rEZ9wyc6WlA7J/T+QF64Jz5MX
FWXw2VGtqPqKi2rag3Kn/DyeggL0DozdZlNbdviHV9pGeQ9NHtNyl+bmysQkWyl9
Wi4LuuByGOMovDGUMO4d7Pu8jGtKInhDd3m3MzW1hXDcNqnKT9Cnmuf/3MrfO3JA
gfYuE2VtSR55CgTAXdE0HocdXURt13h6Hu9LwOFexJl42EHnCpNLCiEGd8XcEypy
ADu1b+zLYQXT7m0SFmsF4Km5dX4VF6zIeHUvLjvHOXMSz+dfImJ27Y1netF6luqq
k8SB21Ulgv4orWC+zdcjc/jFt2wrhF5eWrYr9T1NUPf2y17v3Xe61tDTQf8HDfXv
FV2Sh5Pnh0Z35dcGSf/ECnnIoOYnnBZO1N6cGYHkIHMiDFS0amZa3p5BIVs16MrQ
3nY4RwOX1bdmkQ4RxQK/OQebmPOgcwVqOGK3dyQpD+JaBJYCm9NbJxwEnsdwtw1W
7ZjGTm+TzqlCa7MVlUTd36H4IjbUzsKeEze7DaIrH+KHd3ry2FpqUMxFq/X8liMr
e201/1EMA+WhvO9G0NDyQNQKLReYmHcYj33GIr8DbtHbc0W5cs6aXJuS6CvtIAmU
Ob+MpFfEEr7U0P9Dvi8r3fCxv/o2tIawUfPZNaRdsymYF5+f+kKHagfIqdZvf6Ux
oQZv9d5HKelrkk4KHpHBivRU0Y91kDLvFZh8HPEG9cJdWv2DbBDrJwifWyzdx3mz
ipWguMfZfjtrvjrqMnlHitPQEv2WhCvxCNzbHqvE7JakjbTnLuMKC6F/3gVykGae
VbtOoMXwpTw77l6hkHeGFKcB/tL8Cg+PBlNeZ+NAnSN6rpvzWvS7Bi7iVx2uGgrB
ZA90XghEPQMTakd+VlRI6gQbxKENKmq70RvUS9e51tK3eTLUjDq53GLckLcr8Gn0
QA5UpGPLc09Z/dZe/8u1V4WRSIU00l/Ih+jyEJRxEsJ51e6KqwNdkC1Vq9Uq3v11
ejd70jHnYZ5mhG+Y6EkpiryZcSA9jYdu69SRyLMvMXK1TqAPadV2CAQsvkr7Na/+
q4tro+blkuKqZMRCVlhS8mGxDeOB7/IJtCkRLqyMGMNBbUFEhfNxeFMf/d+ItfXw
tibhZC5HhnrOX0v9kvlQgIMlURaY+wjRs0CJyrlFYARixRtZXMP6okoGceM1RFiM
CdhAVG3Jt3HsqO/cpxnDn9dyyOeOhWu+VB/DreRwrQCpLQxSGY0kl3daWrvfodLC
W2eKPHEaPZKAKMVtvGFZGuxxJoln/7y0WCC5/bD8VamVxeas/JUVmVRa8vob85gy
DCo41l9han5Bm46pEp8AMS/v+vcAdSKWclq5udC7sAPPe5Dyodk7mIbL144z4spZ
LS0XIHLo5nLB5df9gnM8MuuqtVyn4gkfLhc/d24ocGGt+/vIVdtcThu55hgEMC3o
sWo+tuoxDvE9MMg6uZcOeRSjXEKtm347CSxzCO9Pq0lK9HmIdJoJqOTuuavSbFht
Ot8TXaM5gen834Yv/jGIY/4lS0XANloyM+1RLASciD47Datd4eYsS/PEwhZfKEmG
EXoYqHnoHQQfC45S1S4CZP6H/YqpsZuOQn5obw7zjDBHzuTAVfIa6iCL8YYg72YC
A9eUAB1JXhwzAusnPmDbLJkBnvSvVIEkZR3RC1OY17uZRJbUMFKbL/IBLbdLeDaj
eHTp0uI6AGonLJkFDXozHcJvqppGQAV1FfmF+zhq03kwWkPAI0/NeL+aMvienR65
uhZ8GrB9uLXjOYL5VH+yqKDJjTf/IFuA2RLguAl8u/rrw+DadRyj+eY05ReBWWWU
PEmRtQraH8fvmGu5mUM+29PhweSR+dDkdYVxvU5nre7AqftMPwxeosgklOY1serF
0FRHkvJda3izj7jeq1rW1r8OsDEKORnpgDkhHiRZE++qppmx5xBxjUA1pd9n5peY
52xtSlXTvrVOOUpS642AgS3UVqHf13srkF1+YqCYIhaXUdHrwf7Qgw+GjQ2AIOpf
7KuW9URYy+XGkJxBKL4FGwi22XCwunD4zpgtru086aNpavy/JEYWnSOIsuk3gRp2
hU5sqIYgpw5AtgJ2PzjSYisJvgzxVTRWQP5ppFavEgk3JxKnRVoidfkOenIFzmDb
YdT9M9qLxlXZ7hF/4XyTB9ktkBb4hM6QXNN+ikci9A0jkeqrUZ+us6OqIAwq7ucc
P6e6WiDSAYeruW28L46j90+rj0FLREPvgija7Zaeu6jxUqJYLL0EjxvkoKsHJEt2
x6vjfzgnYWWYy6kqxIGoui7m7rFym+doe6nef48228wCqm1iGn1nLJJU0WzFk+3L
ABOS0P0FB8dAd52jBodjm2nXxHKwtX+RPV/llM05FmVNWvm1s598OBatJpJhn2CG
e3AinqqAFbSPDpa3DhQN4ViXfCiRxYfxWhsJh96xLcE8R1CB1GEVsLRlM/91APQQ
FRkWIm/GN7/GzuDh4aK0CgzVlMjOJiDFPTar/+z1jrUYUGFyQXc4VoYGrYWd/R3m
4nfnDwFPcc27l1FgWy9dG3ZIhUZQvdEA4aMXB+QUpSoAP+PHQxsX3OtM84RzHNLF
UhOm88n7y37ATeY3hUpTxHdHf0MGyOFh4yBMv+AV5Fb0wR3xLHcTljk+lxz3tIX1
AgrKHvu+vqn9KZIXjmlycVg2UTun488s5rMUQADS+QJtzWFG26C0bedxzaT0cku0
IbzgwyGDUiWllTgv1dFyJmjMLfQ990CyvJVPUoWjkm/BE4AnlXZKSs65JTw/v2pA
KEtUdiR+dQKPap31+K+p3iY0LlSp1FETfYonkEFdVh7/bOlYqMt8XIlEzNRukFWe
wUhJB1f5u7K3+xkxSW2zQA5xh9SISQsApGPcqfrvf/q+g70cIXjrLAD1MiOVhh5F
vCb9ugp7Xnj+nWbN5xvp5Sts1HtTjWsdKQRkf+L79bX9VyICGcsQm7Guklo51Qis
FXGjNSKoIn6FEgeSZ5ghRixbxZWmhsfbO+7T5/rxd3AokYh18UYqTdVRAyRVKnZQ
akfPgOeRDNF+0EWpKfRa4ZPM6LWfo/bgQK67gL4bcGQaGw9mFH4VU9a0jdKwkegp
6mQiL4CEecjB0wx+2srNxiXKYse8Pgasq/MfaUoW4OWccddqZwP1e7HXW3FQLNJk
TsEBjuBRdYnMIoRSaLA0un1jNjOpP7wiIyVafiZKVNPJ9zBBwwqqrSoMkR0XB2LN
SulehwWOQiOJ25Mlomje0RiSAMe87mp6LrAYmXCNkF2DAC39VaOQD648WSOPmX+v
bLcC+YZr6ttDNrEC3yJRc67dnmf1Q5OUFUzhYCohmqJc4bOfv2MgY9Utsm2rqW3C
kLt3F5rChRHDlIahLlqhyG6ApoE3m/Hy07nRrPo42x/bhTS9S4dDROd7y/PAlhX5
guP5gBg+5DXnVR/DDJLz23/kniAUkDAcVO5dQ42TZUlEKaXKTBI1ASIg8cwiEoCC
u+x/u2aUWV7w/I7KfCcNaO1/nFWTCk14Kp6hKs05r3ZOKBQcACqe317cowCJ8q6Z
mTU8azsvqbEC0JPdmTd7kDMhIi0Yptt4poAs1obLD2tWOqYh+lmHSnhPMLE7FTxZ
z8UrzRS7511T2vABjtMllKXJAGsoaykc29budm+8TWCkhTxdCbwCxY6r83YWX2L2
AlXhRjVoOqSC0IJQub8W6/bRcWbaYKsccsaq0JrMErQNJGaqeiphGj76dyb/JaZp
nLbWQolJWmOnqTkqI+fU8HspTYFvC0dA529rHD2OsCHWhmqa5HRJHHF1jIUqOa40
dJRHnlyhxOp7ejQsbDHKiojBtdHwiO0rbnYH+PhPPT71GC2a2BuRtB+9ZIa+2p7o
EQdJLZbF55TPtNK6xn0E9ZqapMt1Bxm67OF+/2hQSeaKL7+sxz62/HnYT1iNfa66
UDU4nfd3+K4usgDFBrAbWf1lrZEu9QwTtTUkg+i/H9/YOTeTw4byUKNq8CS8e0zj
bCPB2eYjTqB0v5EUEn+4IDtesgbXkEyLX9m+2QvtXZGIxxErw5Lhq3DNRmDsxqVO
lEmT07MJz9wDXG5KYCr0dGL2ve8h9T8BFunsm36kh7hYauRQRtT6lTv7DQLH5rus
3siCd7qxItYOZBv/O7yHqXk9GnXZwQMKrvBYTqcy0BVtVI45iGnubFLMBVYf80mU
no0MkLnOru0kqyYCDd99xKAg7jd2O0qXl9OWESH/wgaLDEdlYIFP9L/gv16jdZ1p
20K1aF6Diaqw33PyevHdzUHf9/BpNDlqW6tybu4OEAehlA+LbCGt6ifaUut5Ofao
qlCjBj4Pi2tz7L3Va12rnJb18A6ttOjBD5yrZ5HYMQcnm3R4wXHWlWo6xnnevN64
lhfEa9eX4OvHdCYnQ8fjqvHAi4F0Jehm+WYw2hGpJl6Hf2UaRxSCDil36cSjyWMa
cHXhrG3ME8Gyit9GIlPyZ9jPbdsMcofiSTz+NX+wYLInUfHlnBPtJNVwsJvR5HW2
Rej44TiGPNkFtZNJcqi/1QMDy6Wr9xT3K0nHmpso4fNxOQP1UkWJaUsnb9/ehDoF
Q9otu6WpnyaRYNY6Z3PrnZ4G5iRXnSd3xLZKRb1GP26NYmSixIwltpQRv32s/wb/
7vBK4mH/X2MOtaF/BqylgkLSUleqf8L55YlgnUbjY3L/MVofe8qCxaFEpysTmg7+
fz7yIXqcPP2a3x3HdAomYEfIvcDarkuqJnsLdEF4qAIfJ0YFI/IEL+R1rEAwpAie
My9vQemm2eosbeNHAVmepB1PtQzA65axN3UXw8/9COwC+UODftUMyzV7iRhEC2Eg
8b6cXGOSKJCUlWeHT5OuiX1uzff7a02xi4P9tJF3IBPEkho5uBAQafIkfWxjv8zo
RYFrV4a5fOLEwVEnd87CQQ0GOMxwUrMliFzyKqyNh4WSniYuIYC12zx40N7vEK4r
oP6V1qbSq4W7TCegNcBzbyZVKrOCViVJADLj5aC0DSQQ8c0AAtbvoWEuMnV98NyX
kNHCYdoeRHxel3gGtGzdHzzTZuqhotuKBzDbekYTlMYyYvjfkx4h7jfNNts4aeAc
dYP3RwqrZlKj/OfR838+Nk24B6CjDH/PVnJIhuVIA1hLoG1D6XsbUCTyx2WIN4y2
PIKqhe7Uz9Gwri7ibGUS0t7Ezmwhgk5m4/PppRujt49vJZ1c6ay4O9phPU/jbTZq
gEe68Ic298d5W+Xqp5wAlJJ6UecYGq3HAKSkvC7dIuPyGhUIIO9SewobXG3GrEai
qo6RaTZNv4r1sEX7CpJ8eNJUlvQYW2y0o/GArtxWd5m+Md2ewLb34hbMuKkxdf6T
pP2LN6CubYL5QZOZ3Mmso8oQx5nrwH0Sm3wiyJg9svViwjogr9pxgMvEY+i3X3ip
P+L0Fso1OhoHfM//HbNm86xL1ivaojTbMNGuGrkeqj5hhB+w6iCJsHrCq21uFepf
DsfL8lIM+FaZNJ1+4WPKFE4t1cGMC00U8h1VVJwLDYBqbb1m8ehzry7urVGRdexV
5V+M/AN9fyfLeNVgdbMCJtMeUl4+B+UdkcMsB3UsBaVhOk6AZ/MSkbpHz+WdE8Hn
weUrvOqFTbkSOpZBtCOspj+yFD0L7QxfANsBLpuBfj4MtNS2Hx9v0VE1SNcNPewo
PzSE6npSk4z7C93M2DevLs2r1zrNxCAQGo9WtI+c4Du3m/hTLPcWWWvMP0bTDLRV
EE1vV47m/HCkQk/nB8sMIiyE6aIVJVqLg+gKQKbV/OUs/f0g0IbsQvf3RA4DKCAG
3BMu0I0Z6A/W08boAGm3GDtcK9BaKDzy10h9MqLo8DgbRVT27zuDNvOtWjV3nHiQ
hWtBKNkGPfnIGp2pnXXgMRoKSs2UmRnnkUE95QLr8EvOtXM7mlKM05a45693B064
fy7O4eom95qjgkI9h+PJ0BPJMpKj1dqaJlUCOO4C7UFPg2JNdOeW/S5h7TPQNqPZ
fsHERUDU1qYFvwxacE4uRQD7GbxB0jRCZmDjo2bASV4S+mXJ00caWjbEshUOInK2
8XI55Anwu+OhYpLUp4u5MAzrqqdYSZwhC6E4qFiAJkf8+klsudD4JyUDSgXwfwDw
taE/KTc+SguR10XELIP7JyJsSdewy/HOAZj4n24VM0BHbjmxjdjsi7tnp/VShaOz
pP8ODP7SerRO93ex/HZz0OaVxG2IytPm6fa3FiSHhMoJjAGmM5wUVP9SfCCzPUfp
abcPs/pjGBL01T5KtIZxaYDgELc65JxzoiYU4mUnNaeC9LwsJ0xWaOe+NRx8dnPL
f52xrV7dQX7H/3sOFJyo5sUjpuI5vzDb7akaDQgftkwP52V5obtywkn+SWQ0XxS/
TEYoqRF746qfui4zLonATBZdtRQdU8HLfADlwGeKJI8cd48hnyOkNGGj4+zYKbI0
15mCw3PeU4aAARGX+CPo22xa2AlM4Xu03wS0ir9EVnRPQYM7vGK3HYAG9943lS4D
5dPkXaAXYoBNm04kTpv0P4fnG7ivWF/VKOEQyOKHLft5UQt2ZwOQshewUKk4nni5
PZ7GRcucfJCOi5daOTYBBsGp1eFBy3suKEUMDauDzDl0c8e9tT+zXmbI7v7fHSfA
AI8EOTSPIJrd7LR8qzRfxUdhjr6cXq4qXlkk/qy8d4iYnjdafy20Jtr0v9ZnXnTE
8u+O+P7kscnUv6RpLmLEC8xL34L3iQtel+jc5lvABlsvwfx0iIRdyZnZZSxmHIZW
ZR7lwAwJnX9l2T9Rj6fgTnwGRowSmtKG6cBqshmIsjRJnNcOSvxFhrW57JYIUMgX
SemEnxZChSEah6OOsyJi7RB3HIwHB5QbDIqPKZWEV+lOpYhPzz7Qbtxmrh+IORw4
I2Wri/AZtjtF1pCrQOH9vPugoydLBoYynrGBSoJ+2ow/ico6u70aKF8Sw4YLaNfA
DcR7aS70I3K6QQ9AtWrfi6W9jmUQ8/2xeoQGdd73Wk4ZGpNzv3u5Qy1zMQkMz9uB
srXQRsUgIDrMmDDCUE62WWOgp2qkdiDAmn+Z+lsgUKXSe2P9vbkw3tIBA/E0j1fO
0z5xGI9/t23E5DIBsp2ghPS7eGFAKVXxacYUmFibJTaGKqwQPFcyQE7Ddo2uJOI4
VoB9vX55oldzBIaHkCOvcEW9Zn+P/WwbAMNicWzig1yTpREHOi6cVNYs5PBZ+lYZ
51btLecKeMnuVUVcGAp0ZRWeaQQ5bYoey58JQ2IzOk7ZAvADKlXZSHSfjBXqo8fi
YSxlJquIPmY6LQjtjyj+Wlfg9TPOEVIMwZRDe8XFhXq+Yiq9mhSzSPRLoY5M9/Xp
UuBjzjs9ggg88U32DRRYcWarL+Q51rRraxd6zz2UQyFDHQ3m6fXeJex4G+CPhkjM
OrcxuwesM+dvM/nrzUYA1Gi9eq8C66vTa9RgwoolA93zX8dfSCLIF49XcG3yUfb/
i/fI9lsjeYrTBI+NvbWwuiCDhqViBObrP3kVaNyUH07V49QzgSONK2zqRbFmphbV
44Z7pv75OrZTB+LJWqrM57CJwI7d9d+RwDu5p06l91yz3VnvlwqYVeQq/7jzQPCp
KRmBfcztwcazF9T8B12c5yxxtRwllrC0V2IOAw13o9Y7DdggEWX0qn0LBcq8DA55
HR7YAHqgrjjq5YHLJ7F/ZoVuBzlTyAlCfI36KXcAahoOjwNXhCqZA4rALJodHKb+
IlskvVovrPjvgyM82QyF8AOfmqL5DHMQfAIlfRXpfv9JyrNzDSpFiVzc09TzeDPh
xlbd/N8Hz5Z+ucHqNB3sp611RaxTQunchudI6KyKYUBdPZ9T8HEDt2BvkhohKOsM
n9e7hz/sU66v4CYXcEDoiX/X9L4HV9t+xbzZGuB1cerDx6vWgOiSq8jL+Q+vZarA
IgOIr3aLvWZxRGaktIvkTAlDcjKwOGMBu/CUuuEoTJL/cPIKL++k50gkwz5y1ElL
9ffNquJjcs3MQCxSnq4VJZ4F08v6niiReFrdftCVDBAYRz9YPFzLRjwrgeafVM8Z
GLc/G6u5pEljd568EM7uJX96twHFNLdDsNXIvfASsbw63k1tYBKTL2+aM/wgZyPh
Z8WtBN6a/gKpuYi7kqy1+BRVhWuOvvvRFaLI5/x30Bn22G4jOSgWP6MmH2L4Lvnh
Wn1ll25hXbK7spOFaPLf1b6a2wd3bETEcFUpMwvhQ5h6tsM5nLy8b9KhlON1Jz0V
tEZ7hyVW69qUX41QZs0z0HPHpfhcKLdlszStIwP+CwXDEpgm8kxO/MqE7rxP6h5Q
IMpMPsXj9bs7hbe1yoxR1+4q0+nt8Wp+MBaO6PdD2WcskeVYoG2+y2/gTniuP86L
+lKVbaNRquonYQ+6qRyjIvPe0My9z7ea9nlGq+AaI3rQvd1iAmZzu4GqBGvIVM7S
cL5MniLmzUZ/Rhx5m7tejTLuhVs+DGv3Xs4b/3R/DC9MDTzeVvQpuzYQ4wxvkCbI
QJaJijGbAZAUeU/4T6qzc9rJm2FmoopYokDP2s7EhTLSYLVq+HBM/mycADGex6Rr
VDV5BiftveTg3i4gC1jkYtKlKSh0+BxyKmwOdeAEfbWWUU9yk/aK19xFV8tLAWWl
0SLbf3O/Ziji78/gdrLsFWE1eYUNjJY3VgbIRTt0W8XpV266KKEOU8GS0XKallJa
Bpd+IRI98XCkbGSlAXErZUHalLXOyUQrlg7jaoTbb0bMXKBF9s3Hj+8HSr/x48TE
FhcjQ16Hg+mCwPK5o4SpZs1Sd+WJXUTOfhGX7ekSCGPbJZHTLrEsVE6vVqyBaVvT
eet8hZMDnqxPfhUJZNomn4rPdbku9Z9q5Eitcu65exC5AurnXANQ3VBgfgHMKfjh
PgDadS8fWySbqkrhaCU6bMWFAC0r/MymmlX+vOJK0+9gx0QtPjOEdJ/ayvsTK9jc
SwT2RzCPGidicSmg8+OOAItfYWAzAF47qbjtxo2weZR6JnVvYjaiIFfXXCBb1XqC
OA9RK3BSUzW0YYUy7z6tBUkAxSOyMw4YKr6l0dA4wSx9rO/xcqaFm6m3mmMD4SMN
5swJEnx0gIcJnzKoNO8h4XYGo8tzaiOtqAlT4tUkE1N3QX263pzbpBpBGnPbAr2t
B4eNIvu5FAfPfSgYwLAm/hrq1IIDu6/0gBRDYvReo2o9pqvWY3/GoJ3PMx7xZzRp
3l5B0+Xa77CM26s1e7XktyJB7e79GQfa3rrsmcQ7+1ukKxhjC7HCGwphvvfqXhD4
/F8g/2uzqPWIXJ/1jQcmpQmBAWeOa7FnRWgF3RWkfcItpqpo7jD0PFIewkCTtjQW
13gWiUuTWVbFd6Ap4qTW3/U9TXr1vkyplRPRsDc/dc1+43wfD+UnCXGAtQBfrIjh
ntwlne3NvVgZgBzCKlr6VlJcnwnWpkKp/5WrwCr9WUzqYHDrPCkzEFpTbuFereCB
D0FUsPey7bJP3aXvh70gCsDEfJcPFbpVh0dYXS6bRcD7ZrgaxjaMYJHHCOaOXT+b
qtIx6ToidRWmkYUcJtJSjzN4b01+wcgzAvdRQqcWLxTAKs0TUl8Dn/QSBEZEtGir
lMYuYfSWJeRJLgL6OPM30NWITgUkFCTMEdjc4DPAlFTSMfI7ndRkRbt1/owuyHqg
SbSwhzsuyM80J1wc3tdkddTUAS0dhPXaDYE17AnBLYpaXAQayTlRtL0ep65MKh7K
R0BHo6DraHLEX9P+1Bg6DJjKXxjh2Vla1HI6DxTpnJm5FwAkDdUcI/lVPPWa4OCu
Ydux/+uO5+F03SLLBlcb3Weucypd1ubCtL9bKi0GW4mjjBsJ04isP+Mt1N/vd+ih
hDTHFi8yMyb/XDKAiyFxAbCPRCFrSdvrl/Z6bWTYMiPIMNvtyBDezzUosaypFCAD
UaSGL/LvgYhVQnY/0Vd6FiUYxAOEvBowXEK6psBVQ4/ewtSCN8PjO8Kc0krUalox
RkOtVvNv7P92s9pzl06g70P9A2N0LA+xCuz8TxA2WbrhmqTr6sFNqpBbB6XEtXSL
mPOOR9u9nVv60OQ1jXZhU5VHvog+fmJZP48BPwcy9IoQosFbaVgokRxucH3m0x1y
47033KqYgSO+g+ZG5P6+YqwhUcPxuT7hpi0A4sGoyAiwO9gQBLDIF0eh135RfQQP
potxcpVD4T4y001VVx8ZrzBE7bDQvl1zm6D1GMohqAVXHVHuQOpj7eaZVwQDWRIx
H7cPs0tSFMx/uUY+iDnh3LEUVwGxmvtDE6jfIJe1JYP3objIvAO6FBQmim+eE/LD
brp9ayjDw3ApCzKChIGNAG2SmpMgG4kg7oSrN706J8bkfFPLY4/BCOWjrpdUKbVQ
6jQXqXZElyYdXKbzJP0nw036qxOG80Us/6UJSgwQQevxylI8Uk5gsovGpWzDS2Iv
jAw9xhtS/KAWZsJCQvvooFzvwIY0KVfn5mqF4s3OyBm9LLkJgNw7JX1VR4vxsmwT
kdf2yUrR4Pq4n/abxR+PjEEherrJI0X0cp0ZOcYt/kl/lfntzKFsPV2npSBkTRpJ
KBlIQYdYbRw4lylIaDjxDar8hL8qTX3UWJMHq/lm+YoMnIWLMiVXrnkREIparDrH
E4J01tNXG6FPrEASLfRAbGedlVam5id74xHuHe2bv0WQKCVTUU4nxCskR81IdxT2
Ry0AkCj2mw/UwlJHSraJ9kGNlv3gSs6faZzgfiLVXoID94t8SVeDcycg1qOSOi4l
y052wQG7+Q16WYZPIEqxqlrVRk1rD/hdSuTO7fZzm1jh5O37hl/5fMM9OD4VFbyX
qnNK3D+ndc2TI4WAWOqWfVb/kePG6s5PWrjO6efaqo6lFae1WHOe9dRpR7zeo5UP
rRgsFV4ftRATpbmUxgWQN7iATkdPxZZ3UjRp+pgrUB5GAeW87L3pVF7hFy5J2MZT
3x/M/GPBaX95gJCWJiXFWFlt3NinY4ZHqHQm4tHBF6T4kfT8jF+s8IAB7xGL26Ts
xunt9RUv3gT6pieZCz4liPyL0FDZ3TJBO0qWTPmySiVhOb6R87ZY+7/rB7aotdF6
NNjZFOsyBY0qGphMZQvYVYk4pF3RneunZGIHRVZ2RJrYpNr0lGtgQhQdxmsdPHyl
1d8Nn3QrJmD/t9MX/a43QONzaJYsriMXkK0pS7tHjKkENBMKmhN4cas+1xr1DWFv
hG0cVwbit3nOUmxoCIYIuBArybYeRfvW7alk1auasIhoMXJdn5pvu2Y/M/MJheIt
a6TmcDdvss303uCsI9HoyeChFJJpSieUvM/EeQRQu2yO4xc5H3YGyFbJmGKHKjhd
5LrWZOyTd1xmWLQqaqAlY+8isyy03qkWn92NVGUbjlGmuOL6fx4G+TlJsDRMABNM
sbYZelCxCEdGmI2138Yv/tnJGSokKqgMgysJqZRx2006GcqE57galu1XbFET7dWw
jR+++JpR5Bz0/rFl1WOXUSLq41T/LNSSUJCEmbcLEax+TSPQJt5FJ7lDGovdmYPI
DUhlk4CMOnenDbGwtEmCTrRv47hTkF5B7stHBchOc46raaCLHZlhd/nTCJe+LnpS
Xj4sQIQ213ZjVgljShu+cYaVNs4Tb5MEFMq2Z830fPFanw/MLT612ot1fJUg777j
DfkGszwwG0NUuPEQI0m3jv/uQr3Mlu9vXwfVcNeCz4ggDN566LJLTPKLFSWZ1HNy
6cfXDxvU1sdOoJmKLTuAgNb94tzz1YGYIi7N85XITgqQJ4S4NFDdswDMDvu2wIq/
t7pG8hfUPZN6wZy0Vev7bwCFUbJjzTDD3smJ/7vgoSNqTLtWltcVdgBDru9zWGIF
eE391NK3f9Wzw31M1M6ovmc1pPDhjsnKNDGVl5lVF4rjf7Q+o3Q2xnB6L9dHxhyQ
26K4OvQRLJOjfvHSGt6jgXjb9SRw42sqQAbUJTgBjytiMXTTVe9yjc3TNi9sczBY
4UrW+1YTncyVEWM3SiKkE65+U8emvbiLzEo8MZ2V3sXsRGHgbHk5R2WzjMIpW4DD
LuXY4xPTRtB33/+G1o9HfNuHAb9c2HwgclX7qxxDiEX+zM3jtJe1xCw2Q48a8tYf
YHwZ+tUsfry2vtnovmipeujdMAMci7oXVYFbzAAfNMs2e99zgc4oWkyqrKi2+Xvl
8+JQWoKWtsQS2R833meVHpbntWpEptoRIdtK3vbgd/2Z33yDMR/AXxp9/p0+i4d3
+zXM02evz+nCNaQUYJ7jy4Ef8anzVX54PvEtPIMoDT8k3Xstj24KSXYXO2qPGeDX
j0B1jqh9cw1MV+KvDM8JjEmTuPiRaPMpr1JjpzA7hruwZhzxiM07D7BhbQi2IEmx
YUqFlrV9s60AUIq1d7nFvnnIxWvwnLXSxyApkKcixOyd3QK4P17g5gSIGAAfUaDH
Qdb2IFrb2YUJiGFZPPqqzG6DSZE9on5O/VDD+oou/FapgGuVPdcV38f3bVHUgabO
szAWXEKzJgAIYFTmRyzzMZJfQmlL//hkchV5ZPOlzPv9sLI9MIC/gzR3KzHhLi7r
8Qxed21jzYpv08ZdRkz5iMEoLLrn2ordOx7e5t94p+TSg14e56BosVLcUNJkxHLX
VzJxAcGm6LwttrUkbl9AbhzR7KZ0nO0pJzFVkbNIR3Rii+cgjpZJOmiBx6G2aYQS
IzCj5WX1Q7lU4wt4C4YF9UjWDr4PvR9UAOagkN+QGrOWvwgNITGQMmzHiOychw4D
bVCa0hF/QqyEkzhI64hLPGuTcfihwDXgZXotzw6rbMZBDdrQl8L/KzkkakgyFnUo
4ZcZ1sK8ORGcY5y4ppugBmyxjplDyNEvzk/OWuZyOpm0cDf+Wk1y5/QcxGl0h75U
X2m8uxHEZMw2/yoQPtF0Ugm+4K82n/TmWJJkahn7lGYrKzO7tnokfigDq4+jEFnJ
EmROrexYZHuDJPi3QQ94RwC871lvYR38CAWj1+moi+VGFCXXwOR600Km8s55y6z7
uXbBchdjSwbwMJfJcouxESbhHXhyCm0jDZexC0w5IokecF6QTHEOkj1qi0XgTfax
qXN22jvvzEuQGArNWtbf1SdvFKu42g4ET4/WSHRCEUuxu3w7e1HBY5u6ZSwtOGlr
5hnApC5F27fwbx7dwAWoEqyyLbgczpu97bcYr8Z/QyieYstlrXkIs3qUDcT7M9k5
9BZIHxHld7672RtFMFcZYKH95zpkG8nW0WntAvZUd/o7EF3W9CNqli7m+OduinvF
s317Daq6f33HPnLSWLQcA2eQiEnyJrPRwHf5JrJ0S5bughsPx6NjdcfB8Bap1rY+
w22Wsi+H4DZ6K+OWM3qYRsgilu2KykKcL7qc4c1RAYr50Zfomxuv4KrbW1oqjANV
3kY+9mZkYKtDS+2+8bWgvZ6ynIUMhGzoHpzFMShTJx/9swjhN1OdChkXXcMDD1GN
Fvu4pP13ZIOX/nY83WaTDMQVOcz011GwQ6e61QmvX9ibceiEjcVOre7rIe8IG8bX
+NuNjlzIL91ob+qSTVJ6C8BJcN4KNUmSvA22F+VPtT4DK5m0wl1xrI5SYY4m3bS5
7e82BWkWaueFRze+YLJroKRc82cHRy9UfaGXXUflu5IoJ45g1v53zUctzzu4lzw3
hGsGfdWUxxHMv08dweY4WV4pOBky3nmzpKzx9WZhcBNvQkNvJ1APeUVQmlVbN0d3
+ZK6N1DKrKqxu70hWgO9u0rwOsfqbIjLUpBYRhCR65EFKgeaOOuWSH93vBFyCKde
XHXpjmSDrzraS2JsAwkrrd19vU0trE+R9kOoVbgWNV6dCenV9mJ22m7fV4Evt8jg
J3VYvGfV2rZ0Vb9tOdN+y8SLjXh/RDKRewy4A7Qlft6Cdkl6YWlyUZH9+VyXY0Db
W7e6fEzc4G9fIm/EuRC0ngtDGeCTNOTyh5qFugERkd2ho/8yUJrNTGDdz1vLI+Fa
DSkvbvGswr5dpCP6f7XvuOWKh2NCGrzkHI0Nhp0UCpNRBcIuKj0UXxACN/jYi6oK
NktKpZPam4VAHsZpLZ8Z4LcJUGoCbyYlKFEuW8V514usZyoNMjP/W2X1fAkH2REe
f4aRchw2XUy82LRxumulUyUk8ZOUg/MqTIk8wR+dlrhaeZmjAROpJsC3PeyNGhtz
KSz08wotA+Hm3l+jjMopxu+jwr8DWYdE0zEbs4q7MViF0H5ECV3MrnhAWf3dEN0M
i/1NI3aHRPVHY/49SQLcCPqPasU8g0EhRlXNOmxX4RU+RAXmIyAQbChHAbyRC1Si
QKkD+sq8WVrzx0smLsRJpwUq5R1RgPM83Znx5lx/gxBpPs1GO3LCyFGNkgeo94LV
L65GWg9jrYqkIrNLwN8jLh3OtjoTCgwEGO5REvjvuTov/SWWwszpZlpzGFFvXT3T
UwdXt5LFHChaNQLhG4P6JAA2KRP514egZewiUiwDxI141rBimTy+XLzxWNVEaQs6
H2hc0UkOLrAe0TufCgODXtTIcoNHmjRh2Xx5O95gZyadX+z6Dh/n2ZzKqFzKa3GF
9ReEsdD4nSkELta6yf+GMJiUQAXWRuBNr9jkIqERNTmRx2KBw4sM+VKAvCyKLtB2
BzAP0paw9POB1WtdgcSNEzqs3UCJtQ6QSEsCWQxJxIpdHuNFgTIscr7vmTt8Y31C
yDBZZqEVAXkly1pBJmkuzYTfBjZVVNb9NAxMpwfEorHTMIVU+Pw0VUNu9FabbbYA
2N4vKcpyxmAQZBveUS6MUsAkIlevb/9YnF4Gsng9ylgbfIFeQEth2Rl2dSPBtIJn
IEPdQfE8I2xugEHj6E8+jNWKj0bZ+6ruYui6wUYHbiykdXDfHmJLUJL/1pOTytUQ
Coj4lTrEnOt1RXQqR+Hiv/JvEc+bD0O9iFQR+KDkkFQ1cp+cr6N1rY1CATHON1s3
MzDsgDTXBdZWJuxA7jBQ0tAQm5Q9M/spdhm6G1WnxFlgkb335CqDEl5JZjaN4VNl
mTGHhtHoa3ofQVl9HsEym2jGIqmMEhhoVr4A6l9GA8fKKJPMA2MwPxGhsZLfLGUG
F/HqltcJevZu91xzEl/ILt/DZatTnnEmWE9c0PKzCV5UUJtinq6UERk46fBJFwfq
c/RaQuYfMGZiTKGOZaMrqR5/A7EXM/SauMSvgIh1z7QeHwcByhQCEeitol12UtXD
SZZsRurQM/FTn/t4yiSdj5JFKNBUQ8Iqzyy6ihi6b/aERGeRpjxAWYMgBOB+zGWo
yv0jja9ecuSbyanlsoga5cW+Zc7+ddTLyl0G46/qKgE+ndKOn0JWYZnj5+zvAfF2
5e/NARPT7IPajJks6fOw+Eof4yFJV0edwi8gnFfNU93yVRRq0tyzt6wTyZCRRMiT
RsJjoNb/Vuc1jDoOWA2bE6ahqyQNu0lwb+70909rO5FSAKghAHFo0YW88OM54ls9
CiYsNTA0dumNAPusvsGGar/miUWzvotulffqidYMzaOc0Ri2Yz23WBANTYMM7xDD
VymSDZtCMjiAknFk4Sj14dtub/ciMr1zk91j8hg27Sf1Wpkci6ZBGiOQQ4kh/ic+
Pztyt/tNrj9nb5DCnva0axKaIgeEDDyJHBHZ4SLWtGFYSeFdvMaKevfTDIBNhhpx
giBHZ0H+h8D4YcWK37Eu6TNS9gAzQMXtc6LE0vMPa9eh/49/5Qd4r4s907wRfx8u
Fesk2AWmt1DRtOUDwWMqqQih6xuVhE4J0a7l988fk0aR+1nq8teJIeCmgXP8kUqV
epdQsWEaIKzaaE63lVKjf9BHIGtjrTcSWw+lLRW9RVnqNxL+OdllOiaE9o5ch3mW
VKD93VHg6QsZJp9GqITX3lpk79JPjyBpZGf8lfyagpiRBuFEsM7aQstqr/uPvSeF
5CZrMXzWdvm+PBHbsWVBIuY/0PTW+bQX+t7dFkl4p6thMueBfcebvEglF5FC/dRt
cVyan323BEljQ82mzZ7xT3FBJEMATeznQ+j13JrxhLl39E+YW6IIxNKSd4utaxtC
KxwSrsrPTWRt6oZdrE85npjyPE5OH8glkn79SZhPIW1UxHc4RuCeTFA6KK8LdowQ
JxrkiHeg6MUAxBu/Jxrwef+ezuR3Pd2bQ8/nstQ5PblrNAT8O65Ot1F1O0ZTgsbY
O41r9OraP4gJWr8QskRd70CNOp/VZqdjh7ym/CBWSL1PASXUeLQQDYmvgSXvr7Tt
iHlhpRgaR6YP4JdM/XmqRdKUIswH4EvSMYNkRet9hD9tGK7433nSoJRaj/mQWNKa
dDpq4z+cx2OdquoistZ0xLR/qYHw5HNxRdbxIKdYECilqqSAjCLSuJ2m9ZyEUVh/
vemPKILKDSWROxl2PPOD/YdfmAFEDu1af5I+lRxgnA9DMKhgGsw2gXLpWaJd4hit
TXBw6434OWtPdqeQ9WQLctknK4ivduPnKU5bzQmzrdz9nxKVXlq/WeY/7EQO6TL7
eZsxD27bvt/nvDx1cK9Qx1pSO66mzaemvAEAvQ2Mgxm8zFgfnPuKv20k4vQnqbtz
fczSuCV5nJsyjo+q9vUY5f5YRqAsWjhUc/F6gyLblJnkrjhWDUzT5Iv+N86jvDWc
9hmlZfSuszWXUsV5tB7qEjbxx/Zr8K9XODP+l2hh6PSwXjbxFbQ07+ZTnMBOvGc/
4E+n+eWrVEVROT/gRnqdK7mXbAeuNozF6s98L9TsJWDZrgUW7DmTUyyDUjDG3VjQ
X6iC3/q8o8NDLdgbqQtW9W8+OERYKUK9CRMtwC3TqJSUQMr6tI4414nFMy4qIoZ6
Dfb/hvbp3tbuyycD/ErF55845QwgnAU83Y0QTXNw3IrkzZkTzUzyo/BuW49XiMdH
WT9klALu4VmxHvWyRNG/zhbiBxxuqrlu0bTF/Z2Ipkg/izH/nYjS5BoP0NgBYHjy
yZJIMZ4WoGnpuyPK30ltKwHLdrHdes/OeFrosXvOOZNPUwmLJ08jMD7EbKa7PoRe
LxKpGfMEuBQbyPTvri+Ho6Ni3Ki2ygzOL8d+336zSOFlVNx0i8klI/sdXuz4tQT3
1rRo3CVi2uv3Nq3IVwQfj8qHlOz4n1wra1cQJd1Ygxhmw9YHhHiz1z42Jv5qbvqo
a9+Hr+wb/vZQTsAQw0W0NYGd2eRQmFPjAz8UcNhYmAyggZaeLsfWOmC4EjeQLeVH
73Kgov8YAb06BAJ8A5qSFlXxhYKddfz56fxrdu6SHKc6HNdrPtyMH8pAJPdquyJ8
Z3jmDOq0OslTSGeq9/M2/Bfsk2+/W1fBsjEELn+GfK+s7GAUyu0BS9VNxRj/57Qd
+6fpEPjqc1gepH6C8rPR7z78MZy9EhvvQoitu3p3eI/zOrMRR3Bn7i1X37AVt2o2
rV7kBkq1otZpF3du0xlHn/VQ6ugDRrwPb32vA9otZuEbvXgPF7Bv7tNTNASqqlfD
GVaJ6Tq+zUf+DbJuc/aF1N2CYZC7Qv8NmCdHw/873qLB5/mRAydwVw2lagw23djw
I2XFKCGOzSAQwQWF/p5R1jI/FNADSqKvWgrF+ERVjsMsmrOZ3NMzQ1XblMC70DtR
NflxnVE17AWpDV8p6+S9IcGtE8WCWaOrd9p3fDGXYe+HMf4azbfypVQCGaoJ5DBH
+O8bKfjo+fUlBsJxvUGpiMQLPWKkalT+ZOjHxOnqHkHfrAKiudxjmaLZxKrBGPfA
17xP5tm/xk2BSkFb2YDlUPN7JodixaVSkasRQsF2sNb6+8/2T0znQaFNZIpZ0O+n
8+5FGPAH/zr3C+Jp8q7pqwo77grUBBtHqo4QWeKX+iLG8Fwb4F+h+j1jApLLK+rt
ywlK7DwvOaRId5b17M63Z+DDD8J3Zpm+KAAPltyGsJZmErHhOeTHN0+3w1N0plI7
ed7oEij7A0HvABpKoqEoNyXa4CLx6Qg4AuH0UuhuHcMnhYLpl3+wJu8xpWKFhj3V
TEv2yKNptTnGfKccOIoliPu4yaBe5pywTaDzzRhnJTuEI1gQ0ciCEUW3YdzC4h/L
dTo6GIi3pVckVMkAvdAeWOCi/bs3uj4kQX+avj7qOA2etq5ExgvkpvWbyVaoy6A1
c9Cjiah8RINspZv9I4Ffqsqi1cPE5leDOFQWaiKl5Mmd1sTIuy5ylp1KcDJCFZ22
/g/nuLEfZTHgFAiTqDatVu36+cC0AKxAK1NbSYoVdnAzYfCDJPSRb1n/UQtm6oCa
zt1oJ2H5XXT11Aie+BRAbZ+dEOVlWl/9KkoOFsbK8seMVqPa6cIPu5NYqTLR2fNA
GQO88KGiI/Rq621+i+/Fv91Z+xtuRXWFt554z/FeFugrfskI50GJeKYl+a0HAR/M
A3p1RntvBcXTEbFx0QJ3/GvjhZL8hSw27sze6mPDmshm41fZo6Vv2s/D5xVLl3im
vqAT7anwj2rT431ldIdUxGc6Vw0iyGkQDAOxWKO06Gv+Ss33asP/I5aozfHhSps8
0430zRdxFXrYwdGsTdUd3nD7nehrC1gCTFhtRwPqnGflTqK+h/NOoCJ3TaQK7i+M
EoyOBBXzkwvojJPHx57XsQvQ1v9pHzDon+54kFTFHIdM5Cyf6/IUIyABlJlYOKPu
FRihd6VU97F9G6wPLJVfea8HoF53ECRVehsZ48KZXkX0l5q1W5lej4/ml0PBMz+T
j+LDvKKCjhPWf8p9BuZy7P3kumdQ2/BfdMtwgkBXzThdS6JoqtM9Mg12P4wLR57A
nTn+7QIDik388zYvlTKEcXLtndS+vRY4chn0fLZkFiA/AJM2aEezy7pIKefNazPF
H85bpCAztzVmthK0OAyCg58dbV/qxKzwgQc4vA1BB1GUMgp7NvXrzR+356JugPK8
XG7vWiPGtGCvLg/0waRAXWeL+6UUig9z9M8gxWegMHiqrujw6gN0UclMDuDBkFLk
sKmYF3ylwf4u44n6Wtj+Y872lfB9vGMT4dIHLDaNC+YuxYyIoSGTT4ozQX8EQzix
ajTQzr+a+LED8sr5L+TU/AaC1FHMAXj/ZdjOMEfHpmRkHSUMAqNNkHB/pvI9GCkB
UNoJTWThB7dPMi2+SxVZZWWdy88qC9rLEeJoAQpJHkBTW5vSoicTJ+qWR4ylmnT5
U0lbTMFjA47ms3eIiU7YHIzPYALHiLUjVRdi8mRu+a02FJKXysGC3yvzjSLV/Iog
kUgDyH++pUFDEwWiLypVvM3zPiCd5NeYUguqLISBjBwHM07U10dUD1gD9XpENhgz
FnrK7YoAEhQDG0NRna0Tey7EnG6qvMTGk24uhQTWsA/0t3C+GkZgMLmL4ePXw3tf
johsB3sMIpW7GULNUpZMPz2kY+X63zc/TufLs2f0p9MVNQNape8zNZAj6TGsfp2Z
iiqT0hvVLgB/FxrUVzuhaZuQXuolCKNd99e3O5UOLWqPlPcfakRxXDjF0R8h0Ac9
teye7D8eHWke/UqD5iYGVaGikYPMXnFNDGwWAhEvPrJeQTTGStXJK5zPGFr/UMVD
GaR6DgK7teo4vLYx3AsblgC6K7lPYhDc33BF3xAurzdV5MalCZwrtJ9oJqIYkdO1
RO6PgvmDpDvbfxBWpD7SHUIxM7VZSeCr0a3vZ8LVYwfE5mKGUeo0hDFSWX+xOMow
GdEVcbDoJ2DC7q5hkGIZ6YGpYXt168WiUbBG36UQcRVVovGFrTShEPKuNwx0tRED
DJ0UpfKeGn0IzReOrl5BXFkCqg9VNN6SjKhwDw8mmtAZcExm8APhTHZPlw3AyahV
d3ADvw9wDaLB3kXxEX7u4nSX5w11Pj1W3BGucUxS76PGR1BCCFSk+fa47tDcfEr/
gvpj4NGFnynq8jgcIfJbCgJajsKd6zLXMhLQwhHnJW4BnH5rVy70Wy1UfSP7v8YR
4rqMI7O9XL6s/rfDyjZFjIo2+dtN4F2t9q9PQUr4Xoez2/elYq/Uez7jcSpMo5Wn
0I3h6gE/PtyMnRfoUs252YSzy8zmCfylAWxVJq76e3ZT632s6jDymMXTymqFu8vm
3c7Jm72Ohnxgg3zLfHeAYYJnSKMwaG0xxEcPo9QIvR4jaXi9k6+n/lqEh7fK39Ki
33olwkhoDb+qUtiGiMoK3Pqnl1bBzgJPe1szT842xEPgwl//zlVLUzHmvv3B1eve
g+1sSgU27iKTi6VMwEUERlyJGpXC7a2O3rDD4NsU1LtdHobR2hM6URbMPVYwvPQL
IuJJ7rols76yn7JP+AQcIarF4XCnnXFO/4FO/66kdcpGPHmR5R1lK8Vrdyy4/bnw
cpXRFB35/ANNipp+Zj5i8JPHZgfA6SmDoabbCWS2NhrwA/KqlVHgdObvxgJQ42pi
blS4uZ/1omOCi5R13vCcJ09e9cdlmodRYYonRLuqtLDnyc1/LL/a8omzcBc5Jzlm
F8nvCUF4kp1rURoxHOMs9nUVtabg2qnvNDpCubrTxC3gSkLDDDUBbVWrmEWXPt/9
8AMMJfnyhf+rAXAOPRWU6l665KQj7aw0XIE8P7QVHt5dAB0bYD0iUX2LIITrTLiY
HEL2+5cqwIIScLaEQM18jHX7JSfEp5szhVn1urvAHlYzJDdEif8Sm1uGW9CPnNnJ
l6fuezy/rA0qolxqs5uIcT1LsGSZSRjXjqqXV/QzGkO9wJt4C7Rqh2mgIEeMqgZd
G1LP0lOL4KqttEXo7IAsW13C/aS0D2QMRRg5yuaopG9cLIpSrW+c1O7SBC9sTOls
P73WhWjJTPl3xFQy3LvUAWA5sryY0BBM+8njY2Gp2fsRd+4go9+1YDTPoSIJSUHg
YyeDku01vjQhJK0Oc9o8suqvDP4Gc7+pf/421CUcps8R6k1khxH3bZXZWxqFTJZf
KR1NXyKJPHSr57K3AdLQzkt6S1zQj03MFBdc3W8w9wWet3ZvnvrtJzMu6I6N66Bm
HAb9a65ACIkr8iPdrAsryv8318LZ0194mG43gHLpow5dNZ70FBaZ6huCwjQyYNB9
+KOFxsQF2iEh/z9P9pJ1bTYGMsgFkqu8/c+ROB7a76zSlH84ZjlxNKjR7+kof7+x
UAWTtARlInhipVco+Qc9QM9bY9Ustd3LScfQJDapJmg7+bWEGxC/n4ILJY2t7T54
u4LmblYFNb35NeuC7Vd+6S2ffaf9Jetr2X/HQgW818SiBeK4dV+4XpCmjzuNr+lz
6ddChYCynmQ/x5T53D/ZNQIYOfxfrwUhM9jD7ophBrdCCbEZ/jlnUqVWigNN7Sgd
vJpnYuvS22iGFpPQyNcS8Z8ldhPdTISp0thukEDktKwYGcOrFRo28DOPcYXtnL+a
MD+dHyt6mZ6BKzP3Gq3HehRLYk0MGjnYtFg9CjJmsD11e2T8kj608CQJGBlDjqzr
jkTNsVYdAQvvUL4zOq+PDSbKScJAn0wq9uNYU5sUcWw3IzFWDuB5mAYLKGMsJbrg
IoVCuJK2u0VnWiXCBLsMsSkL52JdfSjP8mqJ6oPj+d3lOklrWoMl4w7BCIcpUL5t
M2qN1F0qxSOboWuIjA9VyuUF/3fUIY9JBEjHwKxIsiDZaiC90j15dhuPX4fs5z+y
KbHgVcodJjXl/vOknAIQw3HNZ+39le8YY1+K0Zr9qZ990bop1X42sc4GDN3vnDD2
ycuGw2DZsbLwOLHBK1drhdliDLenQAxQUIbCmCVeEJC/77TjCRVw6GQPgbrTu46o
R0NgIGE4NBDdaDrrp4/H34HNODGSh/BQnOmgvsMxFPOEm4iROE08tHwriiEVKe77
/9eiGPL+6g7OxsV7epOtaHX7bsGh9uUKbyiXUV6d0jpGpxkYW7Axxb5rVIuE10m7
6PItG9ws4IgNsKys4TNn7MvVbwb4fL1fzDG3MHtdNoCJ7p5Kupuo7+DprV6y6JgQ
vK7AVsSf1kYjxiGDTIRjsqwRM15ZnzUqpAi9NP2jqsogQPpDrCyeYAHYc/wQQ6iE
Nt6BXmfXuDG3syiP41lebjCkeAsXZrZeud9mmPCmAqm4Zeod6BpDkxSZ4fTXvGAX
ReVq3z1lnc6uyVY2So7XbhJyqUkBjmrWLuCS1zeGumt2BBWPd/45H8plhvqOaxYR
JeLiXgb6G3ocRfHggcHo1tjrBN5FW5rG3e4SFVHTC3EMLCmkKQvxTiWoZICnP1ar
zoo7gWYqRPlDZ+d0jL+PIQMCjuqBswxMQHtUZtcvSEbAWrM5uqErX24aihIDpBsV
yhdjgmruCtRrzjvthnhDUDQA6XmR5RBeppMFv88teNWmjrC0HHBwLFxDSVMRQm0S
awNEFX5GcZ09Fn7oyTRgCMLZUo7Fd/tdv22aCepV6GVCOHleN05ds8Ua4Byh5ICE
yq4rO8D1eI0AwwI0iLfObS+mrRm8UHYNJLca0VYy1SZfaEvfAvB7XleTVHcTIRcz
K6NBcTUZ47STDTtR68iVkJ9vHU4eUA5DlfJh/D1Y0gAaznh5RitII6hvw8VEDSqH
JjI3abNghj3elsUF3A8TybmwmWB6RP1BiF/dJKnLppIHJ/9O9291pNbetKS5UysU
lW83aecALKSoIk49OH1TmUg4/N/QAlkUnJVdPiuD9pkBb2n+lC5V5+5YEUD1jQXF
PgpVt62sGr5hH0RO7Q5rkup1/mCrubklGU4Hlp64Zs3tsM1/rwK1tmP5n4hVoEeG
insuboKPyqi/1cJqm32fCvg2hyLb64CI0VFHLTIrDil28Qif1f+1QwmZPFVOddgo
RyNWOL7rlVUE7Nek+Jf2xp5rDjciLSm/imfjstKqKmAlFnO9c9xzLdi8xyFXA55v
OqrUPYOrYbAIn9enGav/SWUHcgzFgktlkpfq+RgdIOzozC1y4y7tMi9jTeYgxgGx
N3RnhGXp8ASoXUD8KQhUAiSGCKSvI43MAp4CmaXxUsVzxA4jdjLePuuyp2i3HCVM
4/rOPj7vm5R+nWhciStMjPG3n7n4WPAyxdxekGECCO92xsb/vNJsWJqOhFfK+5N8
f1aQJFjRPQ/YbVEJYgexsDtdL4U5JEDbqtB/VBQJUCmhFy8pTqkqoD8h6jvioY+5
TjFlzs31kJPUnYPxfB8NSSF0o6IEWFq2Pn8KJTGQL+oC27sf2zwbu5dMctJGbqtX
QiDuPs9EhEFHqXqQXdLXi/4IfYS6FIKwlOtJHyALh/2fspYmCQ6dzgLR1L+KSX81
dqZHhsN9hDoSPsWPDS3rcdIa4vvI4Flz6akK9dvD1SPfQI/QiCyrymvAji+hEmV7
7XMAMHmxFjF3FTr+MeEGMO79OdDStYAnVmrxSLwqXVrOrCwSuRzZS9zW7Yxtd9Ag
ABM7XKe0t11eR4jRaQf3uYpSv/5hwRQG0KqPLbxakx5P59FsqTK/ykVtH93snSDg
IyQX2f++PHtce96AlCi94kio7CabEcnlkmkMX7Z7NyHXzNE4hJ+gjEBKxvhUCUlj
WpCRdLeHD/I1NGAIbzZq43GL+7vSx1qLgVktx2GGbdqm/u+13XOKjsNKb6igVzsY
p0alKd76uLkpCOTnQ//52ZH3+/7HSlqIRzp32RaXNwmdFYZ4yaNkfKnKOhwDs/Kr
0+i1eUrBmyvNjaeHTuy/WowQ8ct2ULWqFm58tXAN88KqL7T+/vZM6FOKoQKlC5w/
A5ojvpyU69MFXZWNJhxvaDgZV+9iqtP2yOQ2AKE1h066KTzdde9dfl2MgrlQgwCl
kZKi5ROUs8iVr6dn6x2VpOAkdQeRZ31hd2aU6GG1MByyqvBI8SRmWDSPuxiBgslU
+MVvqZmXyz1LURmF84+zch/EiR3fHAk2wxFoGyQAr/zhZfKW+Wt2NB9/Wmc+mTmu
IK3V2LfI1kdfS17JqfgH2bn7xbgfw5ZFSsZdwU11Fyt7T7jENJTgwyQRuudP4vm+
08b63TyuhUuVcN8lmV3raSOwp3YJc+dWkumLuyeQQOxMVBtfXkwxJq8aT2zHOo25
Q8q0E6m4GPGdKGks9jBVGvZ59bUS9oWS2zyKY8Y2FeJpcskI3u6zHGjZ+jP/zQud
nQ7uBwaXlxz1IildO/GIMx0dWSwthoJZjLqaKxOqmBg3wgQJ4OTb4BbqeYO+42C2
ZDycI8Q2tjrRDqfoZPey5JgKdh/GwBAs208wAgHuaxPp1Ay2zddfaj0elvDq/z1E
ybYqbfaCtWPdUmf9gI7aA7eF1JxO4Pqfgn4g6ETYc/pJXYcdcZGcOLpIR8+92T5O
xNYAYbFKm1PyQpo0SsADcXAUW20wCVApC9dJC3e5MZp+Y1CDAdJom4rxGv6AD/vb
wo9oQzhjrsUe8yvas5qfzPABxcC0weRtvbsi1cf5lr9IUyhZy5rA5GlA/oIMWsc8
vIJlxcd8LgyBYIra8kSO4bfMORQYTHP8k5Gj13ywcbGpvm5Y2ggwl266INwDvWGk
Y1Be5crOiSmrvUcsHJEQ7/nYnt1lowzljsX3TuQqM2jOaZJV0E1sau+dv4h9MIO5
zzzsYr6jGDbuy/3SihPCi1sMNncc/uTFDr5CKfz0x702G6QiWv5ElS1FNS3/jPuo
+KWp2vtUdVplNaSH97mUKOG/l+Jiui2TlgAOkkjkMadgIVQ5lVOcczP6d+SJ2Mkh
YHUU77ycbhxGTNU+EXFIVpEJVSXVpcdnYhk6sDbjhWxWqEdz7n7bQxuYAmauq8RQ
w4hqXQQswc1Jgn6pI0nsXwKtaZ5ZAx6goMWdwC6vbIaFE5VfwuT/5febu8JXpr4Y
gk1CeyzcCYozfnMmHT1uuty0oF6sYFDJFxKIVF0mGXPebCMzr7ZrbWCS/bNvcrFJ
KEFJTAbc/pSA/XL1Pth0HlMGm8k4yHnOIHDOfNuIep2cnf8aCJw90PnTX2CcWDIt
IsajpQOrgvCYSTWY2rLrs38y3M6OaDGhyFjND2+hKUNQONWMFmskf3O76yudxLaG
s8mq5mFaCJKY0RqfguZdXXAmgYzwrmJRXJka1Aub3Baj66NSv9y5tu6Us8hpY2iO
9yD6o4KzfFt5eiAlGD2j6aL8eNJxwVJUveiLgQoPFcAbUV/vE0Ea2n4TjvwYBF9n
W3QH3le3RXdWnIjRcKsvUUTtpSxhKNBiEuJN2jtMuhE0UlVZJ/P9szl0GNuvKVkK
SrSsXIzEOoRvYjv9FmeXKV78CstlkZi+4tY/7bGx2B3QtltIsmk0W2BDXx3F4Xsg
WYZtzkIBZv+w8znFEwUzPrVxQjwFZOJgBrwFtfB2pGKQ9pbmcVlIG7XmqCpYLwZt
E+XvM7QIyV0EodXjLvI1Ahop/Jwy3CH5ZpDSwA0+Xpbq0xv4n6jNP+sqaX6gRog7
L/jtl865/VouGbNfpBLs3w0LBoueTwYNhtSfnywDCRFPWQ9LP+v/k5BUNSbo7Ffa
7pM/kg3TqTs6/a9Dkm3rwHfz/3hC9xciXFgyEFLksRNbUt3vdruiOdwmujVEs0zB
aAKt+7P52TDBV7AkmrSgY6esW5Ti80YM0moSbk6HVN9tTCqclhTYSQSqNfJikFXh
qOJMqjmHwTzYuaA2SxmSC4TM6Q7SM/unKYMkH7mmehYMJlN+PVrON0Ot/300dojp
6BsEl2dyF4MPKEbrOd5CngQSSpiTTPt9RAAtMADN0bvtYR13CnOTwXeHo+lcWQrS
8V1PvihGpBsoOSfTfujVyaUuQiQK+iulNskOf2oKSK/kpeWQ95DyMQrWZQY1rgpI
EykzsG4xzTx1EbTodD+4jpDOxIce4Ozls9GfYJM1WaDoVLJEyNNS85sVCfVqVUaN
iOgw1cq0LddBD/FzgLO+WllenX0Y/6VHMMFvMKE4855LdFxe2ogAqE+RXVTcG8uO
t94VdAe0mvqaK0NLwgt4lVAHe7MP25sSIyoowSusdoZ+5bESU+5jP80TLlRSqGdc
cUOnoNwVby/g/qDZkulzqxXVR58eShfLGLMSW0dplfpmbqyd9/TgWIWxyg0SzCNd
wmRaWZ2hfh6wPljK5/dwM+QGCRAmGh8CplIJnWmAwhFSYtjeuX5KnaGzgJLL0UqY
qg8zCKPg11A6NEp/2uZn84aIDFmVA7nGgn4p+9q8CHcKWrj2RQ0KgdLHq+8gWFym
Y25dZZg2mcTYG7H35o8UPwrZPJwzuWiE+8c80eIIDGArsmKtts1kJiRLR+hgGn6o
4Y2a4dQ9LDNtXm0Q3IhRMzlkMtjzr1acbWY5D85bSn0EkXaYN8PcPO+EB7YOYW0m
wDbEBCr4irlRrwHnCRWIVwQeAdLr+Gk6iMGGkEepWdUq6iRjM/rSwbXblNpSosyB
U1L1YAgu5ECK/JWjskD9mMrjgl2KEspQJJ34tK3b0BRxV8EYsJQIE+J06KJ3T/GU
lUjnEV8o576eM217D865Q0/TLMZ0UPknh2lqjSCiRmizFt1nSeNufT82KrftaL/J
ZDUG3OUHI1r3TskxQjLCEfOELLdshV/YMWrpgljDP41J3vLhNBZfBnpMwN2/FeRH
rSK0EwTa/kt/sAk1efFDsGeVr/+1IE1nkZA1mtx6FXG64NG0j4dha5cngG7Z3dQF
IfDjecQSLRg6Qiw+3ESY4Bk5XduQlbOdIcxbBQy25Mky5ovOh3lRftuB7x3XcDn3
Fzp5Qz2DV1eh0I4v7gSKrngsybhJ26OpwQPHl21kiPqZEEBVAEJoO4Qm38EQ2x6/
sS6gTRhuEPw7JG7bLepX7QDOCQVGGZRb6U+t9d1XPVuxEjhg2RqDAQfOaBoIUiFl
5DfkywMqV5NYNRyPQI64ZDfqkV5EfNKfEB4R6YCaM3Ni0JCRA2WZpqcM1G8oahY4
UeicAy8Xg2mzk5vMPMPLxiSoJ7ahvFuKoz+IjF3HJEos8l73iPumwZt9ju9zJSba
cjrhkvyUdAvLhy0Ui7gECs5c+rb8O5cU/iyvJsfKxMXTUppRTTlNaVFS2CABg1RG
hbvyIhbe2ac9wwaT9r+ktZu85tNF0gnpwbmreTXk3YZPZyZGl5P6HmJyJVYqJOzg
3kA3agOneqUYA1jeP+B95WSJTwrX8tQsTELUuNQNngEl+nLAtcuvCOcHU8x872BR
ad7fzMnWUlzo25TR6g/VCmIsXpzPJBBMx/dm6vKR5YP5V5szFDAXjoG8TpGvLXVK
63xFAeJk+GvNGD2uD7s7naRQZJ/yzUByvJQee//IPoGZIaNcVEkJob1t0q5TKPp1
+nRsO3TfQIEk6qV1FbB7l9vplphFNdJ+ba0ISowrP13H2mIMZtSz8SRElChRn6PZ
9MN4CRbk0H3EDtW6Rrz/sg23Jb7GPr9hbZL/l93sYvrmhaBkPGaCSSVzPFQSRQW4
sGknGAMAb1udT9x70/c+lVSzLcbQaUngPsZH0c6faCqoOlTnd8YmUv0vir7isl2H
aT7LyWKECne9TrepOiv8wUc4csjo3dm0AO/pHJNSCb4KmW0hu+WsIy4D2peC1abc
Ojt2MEFimziHPZlvKIk+Np8xzTt+5Cz+nkTQ4XvT1lRNj49LCh8tlytRdRZflW8V
EG5vBmJ28vlaKesAjbN7E3Vz+MWQaE9qdOcoakY9cP9NVwx4chuTxpzSnmrNkx7/
spJZZPuZ6NqWDtPN2Qkk9n3VELdM/fYvqIZrKTrzTcydlyo1Z2VM4Nux9FB4ulO2
GUI5G01QpSAUwRU1XLFUjc42ihiXNXow03LW7VKD/KNCXuPcBMzARALTfweutz5N
GZ6/4D5pT8+sNjFisfX1AMYbtXYGVqBWB4woiHjCAx2SR1IM5jT51kMHomD2YDMh
0Q3NnaQ/ZVTfrS5e1XqOZgJfeU5r0CgXbLVDVjg0COXcgkVo9heP2sE3sZFLBUyI
bu/uDc562vetWv9IumRUMV3HSpCAQRsdvNAYhLOsLVGm7cUy3Hv3csOUwp3K4Hbp
IFOm31tJS5j3Z8ntlbBuu4sKGGB5iq4voyMs6naUSR1LnN+TBVQkTmiEwWwn5Jl2
ebvCeNkjRukSe0k5inRYN3RJ9c5tH+HRZalZIDvhUVlMp8VQUWZTHr9zMOcG9iZ5
Dtop/U1SqMgi9MSS5+Pl+boxBwchUqo6cEf5waRKWaIn9FENAu0yxc99gRzMAh9Q
TQ4fPdfbsk4vU8akWp7/HwJUgnGBXptf2bqYzRoBm6rcGrfNu5kFdLaL17c/5tEZ
F9EJT66UblzJUimLZu/VUhrQmpt4m84/yKNV/wZSUGKlC+IUpioa9vS1V2BrdGnW
nJofsuuATBr90loSZd6udIo4mKOY8f9eGJFq4s1GXH2s/C9jP1UKuNDmpClFeB5G
JwheJJKi41WhI+LIxhzOUd1k9gGG6xyzsR9gSDECHL7Ue8y8+AD77glWRHa4Vfc8
PzjpAJmqLdh6bm+tVf5BnBuL4p5HUeyRJ83zWm867Xkpfn4hOSRy8hR0g0tEiMaT
QjhxpPl4CkOaU7pXKUAo3zh82KQ7GyNrXUxEyDBb1UDqI9oDdnL8LSrILfkfL/+j
vJhYWeQxiI8qFYIzlbPOoHIWCfR4dMsPtt4tDFemKV/1JNIJub3+oyHPv8ZxjaVW
ixr5QaVqb0pgjfsL25a+qqcYGomPrlFUDtNAhuZX6kBvaQ22bblMUmbApmgYIldu
Sy5bfusvs3wd8dYPk39EVYmSiWPbLusoPMO8D9JcnzL7teQYDAQ9wGH3tNL9CtTs
XOKG5RcOXBQbJzrZbmcqxWVGkofkqlgF0462ZefJIG57rTBTiV+Yd1irgYMNbdU8
JalE7ZOLPCvUGq4teZrj1glenS3qVT3fCP+c0VWowEpmFZx/pG6tAdCqXmALMBYw
UlBc7x8XzmDceBFf1CZ+k8ldmMPSIZmIlnlx0ABjE9iRxncVPyKzYz0954EeUASb
kAh9jo7we5gqwspH7HhU77SIaXX2DKSTvdC8kXwpxj6oVwRvaLVzqzMj6sQF6W8+
OSrebhdEK7p985FtYbvEZ59AOwwy5oUtRNnHnXGwoJa1PxD4SHt7MGbvSvTKt7fB
Ad+y80CH/wzrzMqNkGCYPXvpRHgj3TOvNGIhrnYmLkHiSC49BB95I4IU1wCd/xL0
rSyejKblUikx4lqkxNot5Tuz6Ertmn9XAZl1/WvaAKGR0CtbOQkjk+G9Nrld2Qh3
rSBnK9quhV8bisZssnO8l3MYxrc3cxJTWpWP7p1PtiFVRGyx3cOkp7zPZL0OHM7X
3QDpDMMB2cLmCcDxoVSw0mo/ruGKBvn7t+wdUTi2aa0k7OSMwXjAII3npdAEvfiJ
EIWg99qQ6oRjWZVd0ctUQ0IXGcdSfN9FFiVCaJqHTU+Biey4YveCkfpsKIRn5pKj
BVTtnHd9PEHngLViuo7dziwrkjnOUCgQIKSSWMrGKeicY8zeEE+C9VJLKhSUei8t
nb+aogaQ5Qyh5S1jo/lP5NzfxYaU3HlyJqjcqpxa/LAkVRgoGEfkg62Yn89fQ/2V
5nMHZ9tPsg9MlaSNmWbGwud8EHONVYDvgkrdcEx8iIEXC/AleA5IOMb81OJUJ2hZ
KdGTGF/HIfqdD7jNdRrch78hz6okFsXhfXp2iuM5D3hTHfAXmt/72yC34RlYDKrr
Q40mnj6QoWn/hXSSyj0BgK3mf3YDN+OtpI1/+wqN7JmweiL3B0lWOBjIcsVGideJ
HWE7pfyTkMzAMTf30cmNmfdjx57MXW6bO0CPC5o/pKYgA2Olitu5sY3GCq+mHrfb
eyWWU01XbjYzsVrxrcSFwD1NEEunW0VVtsSJP9pwV+kbzn/i820EmRP2RitAjLAf
tPCB9Vpp/55Ihtdfnqg1Ujv9GYA3uxUm/ROrhA68eaCQ30IJMjjuWS0AmxRXH4uL
Z5tBx6gCwC6+Lx0Jvz3tQ7OS9KOZBBXVw17wpPuOxapnAQYiT69eSxOPoZEMWXxy
VeJdl3/KJPR4nFONcVms1pLcipxap1Fdpy09odHL0qq6eVkng4jjKs+5tQVHj8xZ
IGFsukW6y0SGMYFh3trWQy1mp/CrEOE11oz3QndK74axqq5GNKSdKq/ZXgMavb8i
Vflg+RxzZQ7TqZnk+omvUvHA8bfbfWIyrJc4xvMoQl3C371LSHlAlIj14Xd4sM6N
jcmrbL0MGRa9OLsoWqgioQisccPLGysqHKbwa7qBe9SJ25fYWpAijBmoTV+2T69M
GNAZZ2GI2rhamihEad9b7SSMDn5yT+1l6Q503WUV6Uuw7xOljpp3Nns3ggsSjUCl
Ko55zZsbvGpgFVt3E2RTXIm64lgFz304rfq6cwEQr4KU/mmACn1dJYQRvUqZ0OXD
28Vnp+p06rbWSa//ACch4NvZ9R58PWCqApxYXnbT8c9RltH2S/Fm60jvuHk40B0G
yk3sWt8M/VnagNx+hb5XMTZWygx+Q1WDOO82+0v9ByJJy9xzFUtsCNXgYhFnXEot
jVCVtca7rF5ulHsgdRe2MuvQnhQX79fRwp1V5FUSGUBjDT0bjDHNZ8zFNQ38EFHl
4JmzWnmN3oaibY1Xi0RhTDyFAdFxJc2ki4UCHB9h4v6Vg8fEOqx015FL0aWPlBoF
V9PiVRTSh4hSiJbxFEhzDOZhGn18Mpj0Lgnvt9Q73lSVMiJ6wmsO44QoJD35FBgC
li+4ktV3fKr5YEYGd0kCoC2ghOvJXrXicYfMrM/FaYVL8cudKt/1FQri+IMU7QLZ
823dHHwIQaKFiSnMQgrcKOKVn9MYH6jEVle8NbJfo5JM9EAprE6WTr1BuKTNRqgl
mNy8WKSQz2pE46SslUd43U8VnS0/J9ZGv+KeP/vBHtE6TR9elG7+M2FT2GuSQ54R
f797TzmFnmSLV146EYFQCM0SUF4ODqcCEFxB24/st3jlpsvg1boxhJzJjWLLIvIL
x/zeiP/+AWzUouzzTGn2N2DZgOQZLnZwzaGtjvxtYb4Wcs3H+aaBNeRUWs4j7lFs
oG8chrKl8UEnUqmckZokNHU7grJ/4RxREDEM533YWa5klVnzxPSAI8YZAHV0sQKM
hqdEFBx6oWaB7vVrxMep/krj+Oy+GAW1cIDjdLmOHOkBanzEBK5EVw/og+ayu42+
Lvopur3YW+dFwJatjXBMJAg2eIUafpPXXpwl090tVS64QOhHzkEh9nhmDYpJqGfh
Uc8rCcwfzzj9vELP0OyAQsto2B/1zZOkdTU3NeDXUt7CB5xmnSbkCxzbVutvWE4u
8oUDAOXJPFimtaXjCOsTYTeQJGIXDWgyoLy54Va+U7mkH9twxm1W1xAuEX3rMLbi
384M5gnYpTFEp5EbDvjpJrVU0JIORCPXFYffTu1SpqiFCEKHbOBdYkvnMEyd0FaP
sUw462au/1ow6f4crquYD9tC8BSKhrDSJa3LN32tABFk7vE5v2hnYksm9asb9pD1
LiNknsNWq/Z8brad+DePKYrJbi1z2ur02jwrkAbavQJJ3dJf8VQN93TZxGIX9KwT
6O6Q6buk7LzlPXRjiDTon34Az3LFDY4BDimmN9wlhT6myKctHM1m0hwumfagZM9z
9d94XQ4TtwWltngYR1JtN48msEshSRyeAZR4pdlQByMRPk6dqZv0DMo8aIKQFoNq
GrYh/6+BjLXA4zDOkAzTPcDpfdVmMtRmqNpGt1w5t9kxZeOwNtKOYY6rjwMbUd+M
hMn5VRf+Pxwf9aKKNUoOW1ixlWSZ2HK53mChInr4PFBUqs9IIUXwAfLKGC3q7eqV
bbm9R3cvLmbAZubMTodAfDDcoFbwUej1W1RPCg+3GHgbjpg6v1DR8eYdd0t+WFzV
C35zslGbLRwQCO3GzdCJQ8QnHD52hfTzUGhRnO3O3jey3j9U1u/EO4cmkQf92E7N
4yxSfvuxTKJT7z3RSSuZcTQIDjkgYpXjD3ac25bEvh4maLorXkAeZlXQmcWzCjfp
U603d+GWBoYmTRxPN3an81cjNOhTYJasOaOMdudemqoGtkI9Kk/XRAgTxZdsIlvB
p8dGUh722o51DpcoRJyvNmxs2TGaUaFS/UCbkm5HY3VvA1zJ09YvlWhbI8w0odu3
JfQgI+yem7sgXePXQA/UhbR0/e00KtYegTWS1Mra4VZRSPvpmuoQlPQsZmpIz7Q4
Wrk0lzeyu2vpa2mDBLTe42k0JSXsKnUG+hsarHWKWDUFkRiuceM8b6yuxcPyVeiR
3hn6ib/YBhgALmxdzF+u5RRass5GHvSzco/t8DRD+OskralLTnB1q8MRoGuEK3za
syMURWTY1Cbt3azv+ylTorbWgCrUbh8HZ7ZlvX9OOvXMMAuwxi7DhcisS/J+4U/Y
CEJej5GSa6ZOoXH6h3xvvco+gFUzB3t0LcofSjjHSvDMnF8PTxxzmrvluliq56G/
V64KKPJJwG59gKF2xamJ2yp/bcCQk1Gy1BM9Gowc4ri08wofL0ahOH9ooAs0NGMy
gcxrbLf/3Ej+myodEUIDdDtmj+RdWWOtpsBE91MBVbzZx18q9t8QRAeRDTmxZGCT
Y5uLBLYb4KfdA+YujUSbYr/Dp6GsOtwBSpqPKYb/OQ+7BQLZwS6R2GGoQAg+5+gZ
dHWftwB2ALMo2KuYPJaceSfpHycmDfSM3KdoCQiYS69YppKw7f4N1Eu+kPoPUoUi
5YlenynDR2POo377W03p+ExkpMwfuX8A45f74CuO00xfnrr+IAQBHZBUEPlyk/We
Tx0ISfz/Y52Xsiwg+CTao7g37mNPLQV+m5MAaLn7jOxWm0MkA0xE+3zc7EQB2NZA
tUzBJgRGNpHhpllNFwONXlah10L0kLH8JJTg1xQUATWdmtGQ7DsHF6wMxW6zl/hb
NtsMaxdMOiJXNnywknT1Aqzhlqyh4/FsGiMurEM17vIhUOhFskABnL7qLIWBNfp2
V+Hw3jS8Jz467lZtS1qy61QV1vgqBnVjoihWDKrNNVo+LJYay86N5tVeFCj0j+mS
WcwwYuKyY3O4CaD+n6cltD3B1zExPgZp1cHr/NEKpAt+MP3+RMHeWsEqMXPbZ58/
k6qX8Eh8vyH2Prb2H3lWzXRVIQciEtTdeKEz5cMsqrmOk3tPw2BXr0lvgZbkiEtg
knI248wMz2Hy68U04KyGfwVdCe2uIXfoDDj5/iYhrGyOaZ0JBaPGo2YGnkomIxki
Hv1tHOGkklre0J3jxaTxsuryNIvxjOu2AVset28DvqJC0Y1V3r1lcgvS5T4Mjgvt
5aK2A5OiVrsqrdEOmhtJDnrX/Yh4xWc/y3e0LZtffXLWSMnAUvDU/8K4hA4oDkSv
RLAK11xoG+rRDT4nm4RGBwdAF8QCzEMdMceZpvEEAcaj8rqBXSlbRBjYOm8C0/nC
5Hw3yf4xNVvWMlaE+5A3jiks95Kj6DPWSs0QpeeYLfudFw27hP0gCyHqQbtybZoP
rycaSO3Vo/36cQv0JfOGB/+xPak3f/5rWAFCAbd5j1/K1FKtC17FLwt7biKIMv0g
/tatG0hVp0TEmSxtBxkerzpLXvK/EosHfKqvXCmDUdE4S8GKU7bWBlfo9E6KZlD4
Ej0FMZHpJH0t08OVig3Pknftx9c3e7GLyq9YLp6//NB0wVSoKfAwZvCSC4moflx5
Y5Qd4Y9q/G+XpMlId4LoiETfjAl7Vw+8I15wmH2OgVaH0lMnYZYOUA3POXYqMWAH
uXm1EC3yZBt/5HNR7jl2lyKcmpTXJfeLrCkY5UM98jG/14F/etlGrG4GvQLx2Ovx
NOgyv7FtmEsxg1kERElLAB3UUlr1ry7dCTQORnqMzL3pIraj9qtoAZ4WTu63cryS
81KiwQF+Zpp2bn+yrGlaqXmX5VYRwY/s48dD8AxrrA3GlSEjm0+PFHbj2bc7sugz
I/3yH/+5dgy42ru24YfQQBVXP2zIM8Y+H6TM/DtM26Ffpxl/i7h6gbC6ALBQAHe3
GXVpdMsQhhVZDImuD0ZBE4HLdcJNZqf9DJ9WSHyTg1RJfGtfowDBeVtyUO3p+5pw
hKqF0OVEPXIaPvMPeGKCBuFLz3N2V0cU0hcMiIa+fx1cie41a9g6r+do0Iq8zcf9
x6OZEQdgds1zgxgaHqU4xAHZq+N2i+dgnGEATOg9nK1TsMzMyozuErztfjjAf4zx
mlRfNOFW0sSC/mrpoAs8kbIY3ahLldXpig/9XB72MdQbnCcw7yY0RzMW8Z6Gqz1r
rnsk1FmlSBfvzLGAJsQbBSF0dqaICQtQNimjkVcAgsixYBs9BeoXuscYFqZVDKST
JRvpeGu0TSzgmKyHFNkqFKvjc7CO/2qRDAZpMh7rn7F2UUR57ztX3ki7DyssCDP9
RgX9OynxlcQV6HSgMubT2tAc64JzQVe8nb6JqCJXX0x+M2PrtfulV1S1ar3zlK75
SZ65LCVC/yxW0UPQg3dEV4iijgNhXDovqPdLt7IQF1PrH1Pylx8jgg8MeBFyn4yN
H3gEammR61fuaGfKiggc+T+sIQG35KFmbu9qkmBlcZ7NMY8K2Kg0IHn0OB0J4LXM
IkBJDFFCNKJLiQA3j7Gh6jJctDD0Gv7nDyygmpGdlusZauv2xI1EXeeVaaGGgvv2
SXz8FkLXf3PgJGHuTvHXHmytrCjjXUdoB5HeLh5TWEils9xxfnadNWO+6bFsFiKn
nfy/Y9U8Q7NbZKlk43bfmchDTGgMrOSESXnG9HQT0AwCoJEcxBU2RNHhYbuEFkFF
ALtW9XW0q54wqdGMEqy6Nw/L6BhaWjBdtOq853w8ZomYMqMa8B3BJpgE+gS8Cdcz
szn6ESN3zXUjUIj/JvdMq7mSvsZBzeqc+lM7vRU7Ehw5UuRnRil8IwMKc//SSAZt
08AEG/OmoCotrPpBhRH21+8IijRsfSJXvTaTbzhNmk9Kk0sKn6O5RnQaRbyZem3p
gADrg1xG8kmaJdPWgy1AyFqz5cYU7Sn6SQ+ILYShMc7hOUFzWppc6Rej74DJkuaC
QBPBqe8d74jyioYhLIa17gH5WL5VCTDXx0fXbHPze5NCrxrHAgp5E/QhP512UAl7
xIA5KO48OGqXVtt19U4Cj6BqLHqCEnvCuWfJ0MI05lP7RNvdwBccJhsc/XRXLkqJ
ZaUPUIXzNQ9QOTkBfqAZLJLg4ImHbX5wYnljutiVyQWqMKWgXUZbB4P/RAhzFYiF
XXu9puU3edmJnK19DXvO02PKAO2TssJMQQpuc4/L4d6PHr631hF3mStWtX+M8oth
Ci5fq0NZyvl4wGytRmQL+XN5ZzoFkOeA+sH8QOSDalbiJrESTeWpL4iVfJBcsyuU
S3ZabPPCUhBOHbUQFLUlQP7n9hpN33ihnFeAFYx1j5Eu/Q8F/189ynRd1WI9CnC0
6r3JGHz0Tgcl8LS4Mr5MZUU4oZlqc+it9e/rOl8g4oQNEAkB2L/vBhpj/bGRP880
ZW8gCrlTleRaxZJPHXP7P7AbnHUULIxJ0F6nR2qQfjMd1/yF7K2O7pmRw3yP511y
LLIXxWcoamF38GAOCBgcr4H2BgOnnnQTa5XZ1GEhQxQZ51hM0dN940Prd8Nubi6p
Yemo9iS204laY2yyyWQhW3oUgaW/FlxCTibtHi2UtBnxzlXN/qw4HaBp7/9bIAGE
ptDoGf8W4TnqGPexpielPM0V0D5cL2Ps6VIlqmcBPfgbvOAL5J4lOaeaUvi6occh
3pDUGAgn0lehWkRCYzvaiH61iWXxkW7xvUfQmg88WYt8ZLyY5xS9GnU84/hyDatG
g4nMD6TCT/LiTu7LXrG5gm455CajrUDW+4QpmKhWChh0yOdtr7WCGyve3DIvo7bM
0VDbA1aTDhtgpToWEgp53T9s8cM7Vvz1RqUk5m5FgDdaSOPDleQYJ2SCx+nPctoj
/3sRQkaxwKYzvFS+gGLP+70MgJHgrrN/gLvKxPihBfpLUaiVOG/BdCxCxXIDjK3B
ddmPouyp7olYzNsU6b/+7KbjB4aL0+dBN3UMn5xtlV3CpzF+H9+Az8YfxCs24Mv0
7WOa5HvED+FhSztqJ2BL5Vxb1ZMml9kYmDyxxBegUa4JQw3FcNdB5hIyi7mPj5EA
l/nT3tLI9QlpCLjsJJu/0pt6sNwiH9Zc18wtYGNSyTtjoya+WkpLcxpeWMCvrJBM
rcfE6Ln+2uejke4PI8W86qyocmhEEZmcyOqeYpTBqx1IbW5E4dyVCF4Hh5Gt6xbq
jnhE0zlfbA0v8sLKYkXCvIBnMKZ+4VRy9H7gt62hdhJlRx6y1S0hxXOLZf7z7W+Q
10xK/M5+cFGwyR7zRLCFFEnFt+oJNXOD8tbQAB8pYgO6GpCD41r8ob9Ksxp+Ml00
rSc2p9ZxfeUVdrefCrEDKw54qvSxRMSA27tAF7aaaRHnySLavURWeQnP0V2bnDMR
U5ZjOzKY/Zjrpf8kSGBXSUo8CV2ksx2RKQcF/OVtbOOt7LB0Z/ceqBt9U1xU8IJB
yxW/ZEfvW5EAZd5lKuloNvwkffNzV7X+EhpRi1ProG3B0vz37FATXh7eNIUOyvLC
GFwuf0textLL6W2JWgc2AfpUvsLVuHDjB+THtKL1rDWE/v9Kfo5lMwPEhekkaXTN
fnMSNj16JwlpwQtGPSV//urbC68B65lR9uJkYhjJZfiwoZsWr+jz/FrRmvxOH8Yy
jEIbe3oEv1PZ3MMyz0KptCklZdvImixSwpUl4ByVcQDT0jFY0yUc5y4WHwCWimIE
zjNWqVXSq/aH5UOFnZ/mj8yHfTppCO9geaX0jNsCLL5ssjSPRt0NaOJI8PaWSg2S
vziLItOpdT4vRm8aNubaCFs8dZxJy20YoTY8/MIvPfpB4f3iXlqz+3EzPemoqd0x
+xqurrOXrjQBlHTGKQ1Q5QTcF/bJnYn1IgWUqfNN6n+VsJRS5sdS3jorfFierN0G
C9/Hlo+MBC4kHKuMlqDHGhzGSAuvMFv0aY4MAO6PTsqfGspny6pX/PaQF3QskVfs
ZlrMng9mnew38mG5ZXeiwTqG4UjbNaTbN0R+UAIaAxVg3hMAT5kKwpnpcU8eVGU8
TH/XNMCHfaiNjogBvP7SznS4xi+Dbl20/8A2MiawunN5aWfUw3D4Ej5BuzgIO238
AOneAAMCm6k76Kq0sznSzVaGZ+AQFW6IkXaVxd4St8/rbe9dV7UtsGuunjITXSQK
Jq80w2Te0UpbGhzlDu80bPg5p6YhPJH5kiBwG2v90sOMb+rur4phQj3A4GYa/6Y5
0fwkR3yCc+vRAJdDYVrfUoqcE28IlOBrY56jwO63pBIfrDXSuh4nIRo1QDaLy4cJ
N0+gTwcTlpbAFX1k8vJTMLBeSPGEMGftLocAnEBnnwfzAFottmrUNmoMMT9XedHB
ztb2IeBu9NqjcPOKMCa04/AEeLuTTssxUL2PFNmqynUz3VclYD52t7Aia3A1MEXj
UvnUV3X5REKLp3E65c7XkWnk+CFQA7PKAyVlOBzvxnQvv0bIgC0SlJghm62Zurkm
hOBf/8n9ANDGxMFwri+P7F2vs9Stf6/gPREg/ofjWFJ7vsI6hlzMIsKGrYsXC37r
OYHhxwSA++sdN9BcbX712hW6ildygvFZqqJAeOPEI+CTwAKMapcYtkTcxuxDLre9
uzpNCxVsPgMffbl+4KHI6hk35II7phxTX5eX6pVtewayzl735Cf2MjLP2xo4m2rs
+JhdzeKdkd++v/Na/uZLWuxaElIo3tPNh2DVoCixzVglPQ1HanCngcPWrQRo0ggX
jdM8cn55sOCD9OarxaVRYYE1OGwTwjBLMOah+4yLw9N2bpncYytlsIDY22WCNHQW
VyYR7pHgKD4scKl4GPfrDsqcjZ6GST9AxpDWDHc/ekRrLaFattolPIzErKBRd1lu
70dlIRw+z6wj5Ij2POlPNpFJ3BAj5E/p/ihfd0jkOBrnEXql56H+L3vbS5g26i/+
IDLYH+cmhhhAGQ4RPJzzLJUlHTziS6Clom1FBQ79N4kDK4fiT8RHqzbmRzxzwpn7
qCs7GDjDeCUFC94KbdDH8LchpY+EBNlNxhGLLG/QRDKmIxYNWlt/Ymn4Dul/yM1e
DrODlhVSVOvnz2qvKCW3WlvjbFXPRA3wfdrWIO8h7546dMM76r3U06SkVxUzm2k2
ydLz+M6EGFRJh0g0NaBo/U7FUdtzWp0VkDBZdlL/QS7E32mBkv1KCtnCaYOQ23/g
nna6fIDqIzOqJtkczrIX+2PefzDm3/kTZBXTqdJ3ifl84Hk/xJSnx6/WJDnw9VgB
+aL5JM8smzRJ9XdoV7zgQyhZ4Ks/8ObaTBaVewr05iSiA4vM/Q06t5zBLxdUC4Zu
McdaxmlFtxzPM2uYXM7zB4TW1c+4ZLaMuva6vsdc+Zzb5IzvOxXdr8WvF/Acz04P
cyfTXd9dzF7ImrYZ9Nm+11eWfhhfsgkcTEngjOYbbe+gAjIQUl9cxlu4JU+X+7Qe
lgD8WziDDqsrfT+igNJUIfkg5ByAzbwd8K/WJcAecajWlFv8tg7NjYyJ9Gw3UxFO
XyMXrBJKcyd+xR9IbUwZcRsZPR1OJp+ryIEs8m2ojqcjWeeMS7Tp8H9MOX7P4g/f
uCzsphK7180WW2ZrF71lTEM5x4jPfcA7SmNEAha0NhM4Yr+vuPUB7h8okJeEoEq/
6UXQPy9OR8h5G4lQTYWoo4rLy3Zdy1pj+bS6Z16pEYNnS/R5Ia/NVpsviymT1QgA
kTxwGH24gXX1Cn+OnPXFN80Di5u0ddhLlaD2x7EacZ5+vUL6dCXU96KHHrsN84LJ
s5Ml6GvFkYv1xjhhTdf47Z+w3Js4SePGzJBEg31jZahXr7Tm+sHyAy+XoeNZ46aS
BFfv80MMuwIXFKeOAEObK6sMP6Gr/XaAC/c+CdJeXjTmqucVzUTrG1merw92Yi47
Yjnozqxbos57zUGVnpPCZWjhJCeHHx6g7cLIdeXGPI/9d6ewjMokPPlce6qudFSy
TLZIVnCs+yTlxe38c83egrktFC/Y4ufQpH19tnbY44Ctw0y8Xj9j6UYKJb3Cv2Dq
KSWX1zR7A1W3dYc8ATHVjiB4USdEMzVjMC/bUd2N7f5ohTayf6EN6LQW7RIGUaeT
fAO0bybsaS8qPiel1saWgd05QZI02i8ytc0H8qhIkkMjLB0Debbo/xaSh2S6Lq2X
Q1c05fpQ341BxAvYE1qI+fVdexRq2XG9iUC8ItAru1GC2J4DCxurYxEEAET1Og3P
Ev2CXekdjQjAlnYKCSWrdF2lLMaSVl/nqRwR7GUThTKCsBmKc6A8Q7BBoWayehJx
/uMWCXfUFb2aA75o0NsFjI4enAG0HDj1noCtKR1TW1mHMiXiZhGIBUkss1e5sH95
wgjpM4GOw6bg9mmI2PU5uwaq8r8d2V15MzMGveNOslJnZJDoSDZYUz78PvcDr8uq
7LVwetKR8U0PvCIuUeHK3YS4UIJMfZ4mDFOr9qCAoiRvhMFRVoh7Qg/FPHL0XsKY
H95YOLEagvpTcE98lajj+ceRKjJb6KFxaHHTcF+/R5rzdVCh78Qsa9msvIBdzi0y
Iz9+mQxMTALRFEkrV2GZkkn/wH5TUywjhnQkaEDWB1EhKmIJVcdH47Pth9eU16nE
dB6bEyNTmbJBDh/ed+l99XqtA0s+IPBbRs3ohpMRfVNiGpSZIioTJQ6OUsF6BSrp
zrZpoSjU7cYPbXDqwR0Yo0virhfV3z4U162/df1PgB7lNixbbK/EHPc+ZBrhXe79
3H4/ayTF/SP2HfLH/pt9lPT8O2xrSHnMaiwx8CGgYgPFy92eNMN7n+M3CS/PT7IM
TIuQi97aXJOOA5yaUXBqCCyp6aanlmqhAkUmxVcGBmK3Poe3QCwUTAwSQlBch1CS
5/OpGDOehQJwOOoVMNE46RWpSqMkorQuAHW0B+qaDXQ/P6o+LPVYFPZH7+vCCWDN
vOQNJKnxftgBeRBHOgovNX2gedFxaZpwcWii+a7EUB9ymabmFt5LJuJNzlWzq1nn
9tp9Sm8GJ2nGwENYlexzofXXEjGQZktXvxazZPUCiT/a8x1bcSUCv1HVzuWd5TiA
VUEfRQVWFUPBcEK3zTytXjRbt5QE3QVa1kfhMO3q3hN8NFFpgpqzJul9EU98D/j+
/grHRmwh+bILl8NG5jNccsThtxvlA1pbI47+h/wS0LrA3E+oE5tl/IS7JS0+tUp+
oxj7DKJZHl8mWR0ub7Bql5z7KbIf2LvrEp/wl2M+UiNIOTMD9dfvBjAdgXgRxdEc
vQ0nNInRoSsW7ly44oucgjE7QlsYfZahlkxhbyEZS01pEJLyQzkiP9lFiHF9Jx1U
/enjx6/B89AVHD6waY1iTNsAru/SooKGHfxlMHKqOF5bifMCHk6okqjd1YC7vk7z
aegMFNdZTqIQovz8EPsp2ukaVOxbGWInbL8Yy20j0TsC72i0PKsHruWntND9T/Dr
81OLYX+yjOaKdvb6k3HiWnEc35PxrgU0qnXo47BRYTXq+w492EwMuS4dpd6ZH4jv
BU6rYKFpwwTfzJK9ybFdCqOCs00TsbF4RjZT2lr59R+KF04hnC2aQjEfnxsagFUO
/NkgvjgYw4/P9y2iErDvy2wNF5ZAsViBiQ8+z+MEtV5axTcRupGt9QJEs1W10Owi
jWQEjoB3owaFc9KiHPwaKQrj23+tmhA90iN3Mv+MABfo7WytYy4+x9lPnT9l72iF
rkUJVvg2bMWxEZPL89Gde2U102AHfAvYfwUwh92Ix2YzCs/EdMEij0wKQy5+vv1D
cSMzR1BNbp+DpgSMMl1TfplO4nDgtlY7nn0KV4TO7bwbXVskM7F7HOoa7N8FXPsv
wJI9ahYpnpdw/X8Ba8Ih8Wy+xotpyLat7qABchcjnaqqW4bs10Ix8FtHNM3YJTcB
THLZGm2dptgU5zZTB0kwFqUtCUhI1w78GqaOaGh3NmRPCt4n8mFwLUjYQ3e9L43q
6OeDfocHeCG/zQLLPdjUObx/z7AxbtQBdX3oRwkGQQ9e+s1oT8Q4E+xE2EO8btpD
POybAo8oBuam3I7WwX58AKX03jto2YEht9Tugjiuky6HG1NxbCV+6Ktb+4DG9Uqd
U+/ouxxBjdnEGG99ABiGQbN4MO4Gi4Ik9IaCSKRaPDvvZsfr4v26PF3nKF395Tt6
ggK4EvcrVyCjG9S0tMQ90sCCGp8CfbmEzLfdPct/liVqovzhtLpPbn/TpRQqrlrk
DKBntDfBY5OHbzZu/4BDAnn5b0wJ9Ro1q/qr6uKwUy8bkmoQTklZ77pYi2AHM02H
dyd33TvfJl7e8VbvA7fUKnmcYB+XhdfL8jqnYKrHuSpOZ+JxVFsReo+RHrecKBcr
vJMrU6MlZIJAnLQQAREQ46ofCbqAY2LbwDsHpHF5qO/uoWsweh6/LUTbHmYhkNSN
rpe5uyZa0zcjNRKuAuNKLUoxM3UlCoKUHYaO+5WJpeiuhpFdp/3snjDPSCY5/wAQ
IA2B4X7ckNNTiW8r5pSQRNDegLqqWNU/VjKnSiJxayAPtAem/IJd+gr7YhHZ0Mop
VaHsZxuAn9LdHEBmR9/2xa4DAUECUtU5sjCjf07uX3yGhpbJrThOYBOlEO8B6vKc
XFRjkGw++huTU/ky4nMkLX8z9A0C6B+2tYX/PCJ7SzSOkhHASwhAdGuyNM5usNUQ
QTNEJDtqD8LrIngceckPQfaa0DRQLbp5zSadx1bvLYnwq3DNPweEhLUypMJ8313H
Fv/1uSWY/GSplSvzivo7Vw8I3Q9DVNTTVuxze1ndg+s7ASaZmihOVabbtA83c36o
3mq5JiDCoZuosCXeI4/CbqLZwAKmiu7XvREMmDNCdPi1AN+DzvCV1+qoaVCRHiJy
CzDPqgH/aSDXhtj3F9sGtrdMCrX0LAMxHAT20720isa47/JqhcvWA0qLVesCCd0R
nqpGmob9v/iPUSQhfKVTF9LRTeU8xg9K6v3sbCIttpKphDxHqmScVeawLO1yqg5g
dhLQ7tIGD0K6h3K/zLkEAMn54ePy/SMNQiQbpn9h/p7wY7EZAeuOQmrnzY/VWGj4
JzaUzOzymh7zFTCD8m4m1QKKzZE2cejBKoo8UN0605o9UfrOGfupC1PHiAz72hva
Kna/okPPjYfldagcjdou8kitFmXjQfjFQG70ujKDLk3KBrmeGSG9rTekWbftKmgT
ZhFGiUf2PyzRnYp4Sh8kiMrlNC5zkrPcC+tgX5GFKnyrCEc+dENFbNfPBLuN4LM+
u2tMqGa0pOouGA4JgVrYZzhjYacxMBBZzD+jVxYpP+rYzKgU5M5/UQdVcxv4tVgA
zpz3zlV/epUxLD+UinOpfJ/KfMYQ12o5pTZrAor9zDMb42eFwsSsXpiP6j1rlfRd
OuTaQufclyJSyyfQlgVuSKkQbJ0CiBL59p9O1VCYfQdH7B3mv9fgxJ4+GBUxIYfI
kdao0wGjpbbbb/oSCsoWY6VnGuj4kueFg/kDzNyTQ8uPRm2guFz50eqnYDDl9TeE
4gH2mI24HahYRff8/wkGbCM6ChWhx4jmRB/RBR4Dhd4T1jt/iZMjTZktpSYkg+zo
dxNiMM7PHt2PhPhEKOpl9nVpRC134HZEuL8LLpYD5ujMUNdDCvNmo2MtOolD2gbg
hwjWvz0dT/dKuoyut+YBCVZyYpjGATr7M8VyRwBYKExMEx79qpqb8PYl8CYWrxbR
cRlCZsG+NT7/FBnN9oAfnrGzeDKFik4Cvi52IjBZ6ru3Ocnl6vdOUpXAY+xvfQvz
XIvZiRUF4D1e6Cawpbqyd1UbasRJV3b8whN3V7EIxBXgShYCF7Wg42mOtQwWGP7x
wLOLtO2lRytcO6kO9bmTWbSCYmT+hcrmNKNURrCwNkJpc8YSJBBvUvMPQ/e1H+Rv
scfAcyZUXhWd0GbK1mD59YuIhCZvH7PXDOVu5pZ+AMo5Ui1XAm8Yn24RSAlxX6i6
v9pXAMntRTittdttIwGeYk9rEPs71XFBU0fCtrY9iKzHlqXYb2IaLS3oJMzxgmwK
cyIMoFfJwg5Xh5vSjYhQOYGemkivuW0W/PAB7SvKF5PCFakw+i5XOrpzJ0M5XU+k
Q8cy++9iyL4yV63DuTKm5MhTrd93J0YC08HfdMZuYvPvjjqiiIY3BUffdh2FgdS4
2M5aAtFbwMaQFDzzdR/xkGf9GC5cvPN5hMVkamZ5BPVWW2Cgl2a54YnQgyJWFcml
Fk9mHFQbpkoWkHCHVuWNLKLJ0dJrascPktoK0DqQly0hl28xOhma53XNX0ofhMch
KXQ30tV8J9uvq/bG4T+ZNRHzfJ8Ep4oiHfagVonsCQKmJWzqDDWr1cyGjqB4HT3U
MUuukmtTTB2oMscTTon3slEPj/apuEZQX8vb6jUNg3Atisakog8Tw5FO4tiBDT8w
ZEW527WvLTqnmI0wMQqGmDcFs7SXjoCaaSDrXGSvlYGoKFLSk9ACdc76IstXt8Oc
JnirtVe9k55fX+f7cFsORmt6KmRWNNy6H4xG6ZdLbiEqTKTwvAuawYajTeBWWl/I
hrK6Bjwxo5CWkV23GyDYefGWDSUndwo+xIdFX5AEC0Q3tRrI7k3yaSbgyAt2rb5S
xThNh+1fhR1VH0L+zaqYSRHRGgGe+QzAIzKFUEBID8WUt5ABaFKFFxv59ovmSH/z
a6LGz3HyA33e8bLrwOhY7kYs8F4qpZoVZc0bmXrmiNm8mZmvepKyPkgtMPg+x/3W
ixTinEbmgxpE5lJ+SKbhPEL3G9+Vq8/h35SKryNDYKEc9UkdIWEts/5fpg8MPnl0
/6mqntvafs4Z0r4/deb1Aq76JNn9eg3y5e4d8UUVavPVwVMvvV6N2NwpdstiJ9+G
wfjPyV+Mo3mxNZH6sraGmhnmXWfTHbhGX1A3Yfx7z5tYj3kAzTpC4EuRmSuwEWjj
U3gmvrUz7AEqezNw47uuSp2TaLtM58Imr3MkZKkP6lrLE2R5RdFdm75Kcw/XCO4u
Ce2meo9ANGcA5C9s0biynytNX4lCmNvcXipceBu/cQi8SdecrH2VSHC0sTlJpkJc
w9Ajr42GpzH4Glom340tlbWsxxk74OgRlfG/yTc+3u1MBrsiVqOfbVw8KmXvqqWB
Li2DPhwu8yBRIlBzqI6Cui3lUjyuKaPKhY5gbWw7QWL3CwF1W7V4aBj50+w+JzjP
0wsPxIb0Y/I9yevkC/UWMoZO3+o1ljGrhKTvu78bVAgJzH5SgcItrC8OEDE8pZdV
htPWlGY/jd8Fgogv4XD0jsKccLf4RvvHif0Ble2CogSUISxZOvW7g/jUVbv/qrfg
b/N/Ydk626FDI8uXj2pVnSk9RhFqg4MOv03zp2i7Z/y6kHBzjrJLVwyjmC8P+3M8
npXKRqB/QllyfPVzaRTrLWQRjAkBytJ9vT9x4vTDwAGdvgE+AJyNQWtpps7zE0dM
iY8bSuyHefC6obShNy1hkWPi76/ixMRugp1/7QvRaUgl1bPk1HIwvYJpcnx3nzZi
PgnRXxz8H8pSsIXxrtfyj7K2PPPKKGqgVlgV0kJnRMMIjSus+hu8DUHmF622P8sA
KK4dDO8HYaCQi/n1dY5Zam0nugSjC223mFJI83DOJmkvN+rTsz4amkjgwWo7afRC
ubCd+7acIVxt8qNfp7jkDlNuSWYLABquFmHSFHEqqz3Nen38ld2WjHXYOxuDU8CE
5qoK6Zy55+2slhDYiZjCRPHGovXaUuRiSltbBNLBVonputuOGEKroecH3lPXw/8z
0Tz34AacMTb9dODPbTAQnAadibP5zi5rhv+WfEGGAQ+Y7d0+NPc1kR0eerZBxTXI
DstZeme7BJHmSOt+KCfYf+aDqn28zoIpLA7vOPi4y93BqwvcMHi2JMR32091Y4dH
bae68BL0/bvoMnlwbrYAPUYtVgidppT7Co74I2NXJQrEnam3+beRHkYEcdQAbnyi
uHz7K16ZXkNwNgR4miqVKWFTUWHCivB7WVxelKpsUXn5dKEQ8O9q/wd6F8+NXaPA
15gMpA5nBY4DohhbLXRu6SCuc1bT53Jjb1oJlXDfnoIFk+COaBXjupf3p3SaDShW
n92G/frJOFBlCQx7+TBw4Q5sxR5GPjez7fBz/yntSgX9dG5cDInoTzUbUCm+fPWj
AznFuZiAeZX29tIipu4REn9R6BCfUyfe6gz+7fKYXWnqdE1KljQeJ0MRjEyq/YzX
SGPxKcNtvY+DSDB1Gokzo3jSCIl8bIE9YxZRMX876Gnxvq0ceRjEQ1SWUAWBF3a/
PNw1h7xG4+dzJh+co+6IwwZrnDMPlC14+neHORZGpp2MrpXDmLJAlD2rkTeHUsIk
B1Ck9nuoxnS+Vr9drO/47HfFuMViPi2IVVfKkubkiLReTrzPPlHe09t0mBrLbfF4
+wYUfH8L2XBs1SfgVKMLKo+F/RBgxQCIuOzFLHHO0Lpa+lT6/s0Mai4A0Kki8SiS
Du7e1J47U1tRv9zLMSuwEbXtZ+iUpoqZG00EZrY0rmJvLXi4NzPmbBzEhrDP74i/
0JCKozuVloPfjFFZ/wqJUQQ5VKapWi9qKToCFRp04dhzXih7C6J0XM3xp2ajsTPh
kH3ATf0/K5zrfGbghEJ71IwFo1TfXbCnCs8MCA6piH53hAMo3R2vN1UeJhAE0EPi
A6cJpwQ20Du+xlqUCL0tLAvd7uGMPtQx9AXQ9TNePa/YBMTrsa8YhxO82Meq7mZe
XMm/mjd3FKInzYiLn4Y/EnxsCZ7KNbYWT1+k7f7ZT74Zp6XPbY6BDUiKPKNt7IC2
eRcPB+UrEDXrJSx/SucucJr/xU7EtwQAF+WkZhpuap52qOHtp5WCR5toCXy5IHYQ
rtfHgjDnqZq/qlbDzqcBCWmW3En8BbSf6uK8cM3PFDb/g3c97UY+Y+awdiMbBunF
2inECPBIZHVUo8OL2gexr7N5ZPvaseY2P9TwhH0MaMMrLRN7i5nSJNqhpD9WalfR
wz2h4vXZzg5V5D1XYKDr++qGxR5b1DCvWdV9rQGR61q13tOvygJNt5PphaoBgBhF
NvkU2cZMZWIKo1o1YLHkhvr/5Rj2tR2D66If6WDnvWdVpwnLnEMAUZP6zB/2tRNl
WchUcDdCoRcyF2zaqrOgZSFLnCIvTNInhndysXnQFgNTI3XtOeDxyGVdttSUr1a9
TI9YY8Ki2T0FTW8rcHiK8gG71sU8JaoJ4vk0YJbg0mdOy6ztaEunsxkipZ4BYpao
5LhAWKjuigMr12TJO4bGheEgMySwRplYR7GhTN5QMJM7MNJht0ANuQgmGofKQ9XH
knqHw/Uaa2WLgs6bH0EH7STPoeDWL1x3xDp+v3r3fR+dLnaIjucvnVw2PMntTt3j
OcicZ85C7cpHJbFFHyTpvtspcz1+u6onP3x6J+n6yG7XDMO4Vj8xDnV9LKKlxznC
Vk7+jD1onhN9PwClf1YlKRzAAt6Gf3yszvrFwFNWzSVuvtAqMJ6TlQ0FRU++29jN
qOyQUAfVUqdAsYJ/k4cPeF+ocoRChfA6kkbb47lP0wL4K72sNI9VoHhDvSekbClA
SRTGCGGQzFiX1O4bCvDGR1L7nnRCr4U8R0vJsa3fcKRrIfqs08CJlvSROCtKRckI
VqLEYO1JTv0LQZerxnfHHVD8CyFt1HRIDNv9LuuMJmx59t8JGl8lta8Zmp9Tg7of
FssnSE0RamjnPNh5aqbgqAITzcsDyZT+wMKoyzRJ64x3zHbW8geug+mDbmbroWNk
cx5cLPuLz40HloC2hifsya9cEtT+lrereVHTaGBAbF3nFpxS8z6CPWC0Zg2sDDKX
Jw25ghLRWLGYROZxbYcXUJSrmu2vAn2iUkx7wDdaVLmHNBkNB1EL0hEjinPwI2V8
twkOF62TbHNVHIkHaN5XvMAZmPTlbZiDKt2Ge8bcSlymwZSWqtNbAUfmIo2LjLXH
sf72wnhVV0Wo787t9t6eQX2gR6vfMagaqo25rSU3qynaShe/wz3yLtq/j1IcjU4I
87valGwd0AFt2mL4B2m+WW3sFxZxTDizlxAooqmojlANETXOpzjR5QSeq5YqDlyv
O8ds1aEGYfVDrgt8xIZGb2Yik37qT48B2DQ+0yBXQ0QYKlkEMWha4YVF0958bH7/
eoIkwujW0eVbR9LxEt/IhYJpGB05oeccH/v+2+ldjWSUCUal66KoqzWthvuVZFIN
F5UYbtlmxVfBeKWVD49+JHIUsiVfuxjyOtK5KWzVqQZnonuNPx7Myb1H2ofHd654
9ItNEcdxo/ZU0nc+WVWNmfrHPfamR3gQZJ0esF85A9irLE4RjKCSMrSos9iB81tF
kBSwmyTBLOK5UfdTQS5btJw2xGjcv+EKqOGxXg0JwRiiv4Q1Iy7hjVN4GyS8XBcJ
vBYH5Tcxff9I5N0Jk9Y/BRPJmQ0oRbvkaJB+6pZGacmYCu63OjwnhAZ05RmP8u5m
7DEmkYHoYcAePwIjY187sbYpF8LUPpgNOeFSrgjJ+2Azg4lQK7MmHAuHSOO3xnpP
RRN6L1g15QdeW1s0axkiYqIgzkNdcUKv0WFEN2JkOGhguFGWn9V2joFN1oDsTFfV
1HcMA+OEVRe4sEoMXQb3wvfCUoomROOIbpjAxIiLsvXT19yr1UXU4i8ear/H9nZH
RGes2UGsWDNO38dzWQU4j4YwdANuyYm3YQbhIGijEb4ALyvKCv+V4CLgHHYIqkpQ
F/KXdRMRRyC3Uey1hb/T2Zd1wH0aSAzM7Oe5OhRpoVv9rg5H99NgXYxlat1BeWTV
FqfqXL6NQQdZXxes+/I865Fcs7YU8Jr6wlHikzhvuWsj98qtZaiq3GOys2AropTI
jlhtTFyslG3NmlWBvzEL9MBzVwPhJSlVQzJ03ur7ZGX94jHp3GczEbbou5fch3ps
mGbZdFoZq45dGmGaQKxmlvVwQiCOYRZdZY4vqygOLWo0VvF97eiA7uPavxxwRRJi
biwiFqbpDqszp8+aQW07IiH81PJYEeWyTDcJuEjCOPtgsSnRZttIAS6tWUPp5X8T
LU92tX4yOqJQ9BpaMnpKfmM1ZVlLUNGGJYRXcmwbd9Ddy6IogiEFvIC8PrlTxHXZ
+7VMnZx5v9H1CY6YtpcTIcmNrSflE0LNhgKaPQWFqQk0IHme0l3BYMgDIa/AoXnj
8pkmN25EuYGLOj6xhaDfkSRvuLyLtClgHn2XHW/ckdUysZRa4wFcB0MfvR2kBmeE
MobwbP6u/hc+B5lblymMZRaHuFvIIOOFjilcJQV1jE+kIxjzoDBNyumzn87Wnc+A
JTMlEDO+hl+gMDLCsTzQxr4s2iDQmWKm2LYHqMFumltY3XytNINuyxe5ThPKvMYm
hsMA194yalFuZkkQws3mvXezRoJno+6k7+yM8d8o32F2zk03iXXpE8pCQbpFAKLt
hgCn2BIR6hFjQ6awVm5KZ4Tkgcvye3UfgcCmOJR5TkoV9HoYQPe6WyKql31p76GA
lp6cpIv8PkNn8Ct58pcm7wRAkzN1FbO88xKPrA2TDJy5CWlFlbIhSyo08EqKwpVy
fPGOt6RY6PQwS4gG38YFvAOcyD1e7T4CnYjsoy8xgIOyzF0A2w8YtEBx5BkEGxzo
sYkosgO4VsTVGnZk0CLYEPhT+5X2jtyW5/BIPglS6Gpi22iX2aWcOLJVWag63axS
EV2v8FFTsVaz8X1rR/qXLIGYvJGibTYx3LTfpIYVT3NCi2zvT8EOtWOL/ohnNFoB
EOTV+7ixyV/LNIRQUIrdd6t3bA10Azn1pZHZvzE8kMHkGUJNAjjr/MymfhA+Fsjp
0T97n527Vt7xnS51ZFBQZzUfY3XJNOKcoXH9hVzGiPdJkwvS+6024+95JLXIQBtg
Emv3BR3oFVpFMRiAZ1COY7qZUbdoBup8XYgS5LQSUe6U4OZFsAVCL7q2nJH247w3
al6Ug4QQJQLb5Ew5yEfztFbHCPBbCBSWmevHK6SJCtWMRN6AhN8E9YQ3LoRQTBDy
Erm6uXtYOrSOPu+JD4sESJ+/3zcPxPUqqxUrgGJX2SqQMdCt4b/RZSdsx1v38knI
dgK2JWBDWHv45rvDvmn5Iyn2tehF33sq9THPaWqHOCLPt64qD1qMC46I3wAXs6aE
6wHkj02WflGNdg/KbkFY0wf+YrFDJrFtb+AfOnn/B607mIkmwlltbtbCzZJLlZP1
/3QcwS99m/2eXgs1Vu5qytc2+oiS6bt/p0ysfcsBlz3QRtov7bLlqqLVQxPJl0/E
0NPIlG90+HtVtkDiRm1D36zLXlAhe6MVri+36MEd5rPnIpJRl22cDnjwJ5iMIHMu
8+B97VRZvQMdCuk/K1I0SToUU5/gO4DbdEi04KuYL8ZuRJeGJGVZd6kGrkZGnnBs
eRBzbuLVW79VYQUj5H+k2j68lBnZU7UcR49wvIQUsKcVL24bAKbIy1TtilMPclyG
4bzjPvcpcrg47xBpZ++T43PYkyNmTJl7os6GBBnvC1sWDcwcFVLl2IXnqjYSeWNJ
myl/nYqvxybGsh6XbNFWWNLL5q6ewlar8BOC3WH/IWjNy9fg7qagj7iARizR4/g3
mCDAyNky8oLlii7jBUVmsTKibcVXmp7UC34xYzj7H6zDl14DlYUbDVtslIZM8Hqw
X6q58ubfLw/XlRVkbo3Y4dEgdggJg/j9g7RDNxv+KIFhcjTN1mz+a3Netc9yRCme
nXCksUJJSK2ai5MC7te8llVfyOiQF0OrgmgTeaGaQ3VfxXXgPkc3VsTo0D3d6nX5
g4ELksclzLfeWthR1hLo9Qth6goxSowdfgxhqDHCw+l55pGU8f8gOJHwNW6rLT8K
hqsWT3CFXfdCdq4GkpMLussWtIsazBBn51ZPzU5B69+h+tpMzBw4zlVkYJUZSeff
Gj4QIWBIp8MeT0limhe1gDDeqdDDGvZ/cmFacnUvFViZCkq/qZfvKfRP422dYgjS
+p4yoqXmJxUG+b0NJk4n5YbYJ2LxOexC76McjDWxlNblv5u84bcjFk/xAV87bAcL
4ZG8eU6pwCZlxXMVvKX6EInNL9x4k6w3xze9GUWK/ePaQKW0UH3/vqhYy2hMn+fb
7WMFINRAmJr9iP+IB/pGkVRG9wuVdlrWXRz65zjFrFmEy0ZPMXe/ShU8ceFZTs08
EMrYucJWRMRAjJuwsCZ9DAwK95oDVT7cGYL7letFuqvktDD+v2LzAqznZ+Rk5+B8
AFGAtl2W813Nyhth7tVCW+A5/XZnfWbemyfq1uUsWpABSUunvBWjYZyi73RPWMzx
rgf0N3gcab1ZSRko6JxKyOjabpqj66nvnLQcikQ15SbcDRK+6t3R2R3T3wdNEp/h
J9gVl2xkvorIGERTp2fgCl3HxLCGylyHPEebZnIt/dKBsQFRp/hg0spqe8tNXyOP
DW9D7WQarOMPGD0Tsmly6tsWEKeDU6CbJn2K2NAReTXwVgp2vkoHRMT1wBMxLaKu
jycOn3jLEsNytINT5Vt96AuhDgROki0veIKaXsUzx1VU/K4rnWCxm9kIkE/U4OFZ
2yb2/o0Uh2JE+BfG9T/s8YtFx4LOwfycW8/xbOXcY/c2zKX7bLJ9sEwc6mSCmUhu
gezxlywzJZ/0iiKpd5AIHksHjkTjS4JktqZUOmCPzK3wRecWqScHMKeF39VdOAjN
JhpALme48Ey9LOx5JFOG/VJzgFf0KGq/AWyMPlnza5DuciToOoikqfVThccSjRnR
SrChPDAXPUsNphjtVEJ97NLfynK5gzo20E31h+aAjTtJZDxluFz9Si4vjNp1HD0x
2VmrC8Fl4ZrPqjk8+P3wdTSPReF5oHWfnjP8+un2sFFOPXp9GT5KamJpvl1XLL+e
fIZJViinsQktxFRynMShHfZ2rmYLuL4TLlK9PqgzW/IHShC0WVCL54eXPKVDAvEF
4v7jMyaFjsbaygRIOoF5COLEcLcnto7PWxnoI48rf+dD99U0WRi1+BK0lVMfvwJF
tq/wtM0vAreSDZT3xHDmBUb8LA13pgciSfuk4SwuzzxERzOK65PX1brjakYnzX33
grFGEoS4qMu2zIlP4xIcSskX532joWILQFKiXTwlWEcY6DD51EvDpj8FNhI1I7wC
CxIaNNUcquJX7gTMo0Dmqp+iTji6V29LxmZ7+Om7MW3Wu9EmEUQR/5Aeip2p9YU7
egRkADrK307KdMxK631vu36vQ6r0PGwqGGIVeDeIciq0Ae8n0bEHKsGmpLHkPf+T
SxHCKeuJ03pFVDNZ0jK3VgwJ+2P9DS3cKtv8+l9McH8vgUPfczwNLKCMvVmLx78S
71AHyFnRIjehVI0sNATIc+uan3lrEzVYcQfW88oLvyskE9tuTyBeMW8gOdciJGiu
XNypL6KFSYPzTIbxjkzZhtuI0TvNAg3fI+9COb2HFRbabnH3CEKBRAjBuwB5plPt
awFpQGfp9kvQfm7owmOL7AGp97hAUFFNVa/E2T+x3o3t+OpFB/g9OIMzMpZ5TSKZ
YQXXbi1eKd3bTklDqQQZLWxsRxAxogVkjw+vuHpJ6IAKBH+2q6VL9qVsY6+CRFEL
KrUI71oMN2WIJbNV4FZig8yho1+Td/GqizHjZvpd6d3mqDY+0yTUmhA4BJe23jgY
JZuxu4u2y5dheuTh7QreFLdP2km7OQkIb3s7xB+8dDWiLCwiGTlXG8aUyWfqbuMr
Q7zYFd9nvEZJVj5Oevu0ihRTbgozwsTv/dBAJ2X8cGW7/Kl69BV79BaaQ7Hb0UYq
LzLPivjXqno/UeNOSex3vP+b8cCJEcdABiBbAvVYUWUnwyGLIDI2CaNDGRL/x1kZ
tx6iqDSYFKUde0OoGsTbYaBAWZWe1Dk4WP4trrFN3cM4JkspPiTY9w8JTkCDnlx3
XSaEwas63XhyUSX6t/xBbGf9+rTS84Xiu2GKw/kyXR76wXuwIVK4Ms/zMG3Ty1AK
7EO+y1pdk4nvgHTKjG145pkf+wUNFJjs8ZNtvMjP8l5cAKzdX2jmQxpqP5QzZ+Tv
rCVJNBWNGtbazxTx3G2okNc+ay3CzbWM6/RG0oyGGCnXFtagBFHafT/8zyEVQeWy
k6Brrz7OrGqC9RGcWOH86hHKyNw2GAyeNpviEBTFptYcJ8aWkeBFun/0Zyn6zgKN
D9Hpx0zPQ0uhMqBv+SRHf9B+zOUhJHggx+XOv+qgRBOnpVY5h5mwI1ugO6BFfCAi
FZOr1smW7FnYpGKZTMQMMYycrM/QJNNzcPVQnZLyfVTnfgSovAJKuRU5v8MGP5E7
4ZYrmJbaBVo6lGD+CODDSTVedK2rAZx3QGJf59fCE3Kj5d+U2gm75KGIwK5RdIyk
A5WY5mU9l1Q4+kAGqHjcfnGJsCcrL+XrZcnCdPB4eVzwl3p5WY6tciKKuWEvxkQc
pFEPM41wz+svC6BjPbpzrd/BBLJX5cQSjd53VXe6YaAQHtYKLIYUSwRiY1SMyE/j
T+xd+WWX0MESAfvEsjfd2klDVqvSEZw8bVuuPqXu8g5V6E4XtmLvJg1waZYrI68j
fOncElZ8DgI/zTND9LLwnzOyL3xYyj7WmlLvqBQtU0XHNeCYcrKD4GvC4+YKAMu3
H5KZLuLKHHnSA67FySV/uzw2Tats1Orwn+yVu/VOHQuA+Z4nl5gBd59NP7/YIo9E
/LoSSOgc0zq7ZacT6PVTP+z9AF72E5LOYX8GVM1MiIANq29ih41nZKWLJ1zHNX5t
/YmxVI4QnFq5eTZ0EekLg8fW2HlY6VMVB6DGK41mcUswml/kvBpwGPhBXOe5OQ4v
9lTviBy6xjSq/8l89l/kqroK4ppOAqsRWE0NIT8r4z2ZD6KwXq1lzgP4BOlHvfpr
ngPSBIR8JT2kiFhbkWZX1GpeIAcjLOGKPnPgnRfP3PdEF2v9zCa+qKcqsIeo4tvU
bxJRWjpbcIUu4RBS2kxHbFWFUHKZVBBbbeIY2oarPZMonUiW8c2JIrtR7A3I9z5A
eDB0c4mIsDWabacxEpSGFaJtLOLMk75PaQWTD7CzOQ3pyV3Oy74kieIyumfJsjTY
dfJ7dpeYCQdk7yMfykD+8nREHsNHmXgKYTrXIPHmnn9JZgKm6Wu4sJR4abhnIzIb
pW+IUVXH/g21Hx7jPcIeQVFK8VJr7ibyH0CRgC6D0LS9MrhFcXgwNy7S01ZDfxvQ
1RhSry5fOajgsFRigj4ehlHYMn75dZR1p3HVYlJLXEMeYIRzJzsQw4e5ZXq1cfLC
Sz+ZPL31sXwZdKNvRjvcxe3ENbHKCKKXvZw3Qhy/7XTW97WUpz/G2slpWHIjSdSH
N7xkvGdNI6zORra7z+mSJ8b1Pnnksn++dh3QWH3hLtNiX9XJHZIEgjeakalYqiCa
BC9nKZE8TZck4bbCNrIGku89IpVwu8P5xRIAe8R58pDOBOby5rnfYpjcG9tfWDeD
FZNWzVDp4GyIx1n0AF5DfD6CvFfkhFq5L2a0+7xRiHK+Jz2MxJQAFVZPVMRJkBBH
NakkbgRQhcsMzpEq2rwn+VK+d7w3FPlz/XgG28e0N2etXAkvFWJ4I48x3rrtj1GA
XO9+FFEzHyliQjhp8x2jFCH9UTOc+bUa+uulgvMXEcknACixMbzTVxUP/XDMqW+O
QluLzXDL9lwdkWImCEudhBacaKzBXVnBsh7SttL716qTXzg7hItlevOKHxPylLjX
E+EpyPt+/eMJcEr0+b1/eXQO0tZ2UbhIw3kf4pHTr2miKnSen1d5rtEe9FuCTx9K
+wReqAanBtDO+L47ijK9GiRvIEt7SZQawL+s3C4CUEZHGH13F36iowomH6BLm1uV
FdFlKt3a1bYq7ZhKrOww6RWSkplrOhjOlbBKQHbYmRKbBPdPpzqGFBotIZDwI6Bw
OlpYV3+tkhQlN+ZeOkud+0r3ErYsInlApg9Lx68ZamRNhnv4xG4nGZQTFmJ4P1vN
OY7EWs9RBEUhyDSuFy6gYPZvwyeUYU/JpKR/Bh0otporiKrwjVUAg2rca/5Oc7M+
Y5fp2z1xWZ66McsPM9gjyIdAgChLis1IV8kNIZ2RQltTv2YXuWov5plJtZlINk9P
Ggjwa9oAY6MkdQ2Lqr+mzrq16S7w5vjYpsXt9u597ZXcW2E5yBXvdb//O2G3Srq/
Qia6I5zZJibiaGM4ZqSAARo3uueQ5Ve8lbfyOxa1Xwig3nK4/a7wwkisBZB3Omxu
8dWKAltivr8ye8LNJfhYJmcL8ztxFO9tMJl5v6Uu91gvQA6cVU2uRYN/9W488l1g
hER0zTjeC3tKo0uyav69GZsOo7rr8lIrwG+8i6a4Z6GYjHjbpoXgt3BvrDYR9cYu
1UZ2Q8Yfu80mpaAeZz9+9I57lU9prgBwL4g9X6A6WLswybLuEsJbbopLMIbUr8sG
Hw2BA0p5sLIhGoq33f4lt+XIgmrESnPqYxl0hQrw0bKPCslet3KIUi5ShF6Oayw5
SEt1JyCcKsr7mUklUAv7bh1R2EtdVb2ibjAtzljf5NpRq+xoBIYj6Uih1RDReOvk
AeEDqC3tsmMGKGkFq+6zdPuRRoyARa/6OXEPebtHIfQczWljoza89ssWyLgIlInH
qexZBSqRRHpwKQGyfoioAsA+NU0PkdTaJXi8DkQ3IZzYBZ2xF2uouDuBFNtcx2gs
A3ZHByA7hl9KwU95TgBqkTgJgdT5YDxa2r2SojIKs8ocFHLeifqx/4lpbd2IGj6i
JyWwbgcHeLKBXYoJNqZ/n4IdHZCoqFizi0nN3fvAiEkc11JuhnW/67caQ7hS25Pk
j9L/AFIFp9/oHpe3B5NKsHUf9dW/oysYdFkCIXMOhymgC3Fd7DEGddYZ7Puqn2yZ
+RIb+eUA+KO7RtSV8QhlD2otA9BWPyaCZYLMH4Lv66HuSoYJOxwQgSZ8pKRQAEqf
kbUZZ/VVAkuj0mLOHtPVnVPFPs4RzfYtytuiVhh56FOuiIqovtGvhNx5p9QtOh6b
DUiwiSDh/xumCJyLNc1DramE6A1EfdgjKHB2HS3H67FsyqPFtjQ9SBBkvWkRUaEM
w3/+pPFeQ0hFClAGYKY50/NE1+EpEO+6oDsf11qddktKoLlgumrr3xBeJX5Xrzmk
NNR+9lhzV1jpFbc1MK92tMjhfsKqiFR/nNGlxwM26Z6dVm3K9wqMP1DsBc8A5hxm
/hRSmrJS0+EdCn3YO3Dz8fViJJRvvbLNHEm3FYwKljRxlfSX6RTl0sojuQeEvR/h
pQrR1XgQRGejaEpw7jzkeNQBhFqyKeAlnp91h0dkmu+5B0noxq0qJMyDrhv9XPPn
b0RTjfKoONW34WKlUwWOYEI/vhR6tGd5Zni+2T+vn8m+y/hf+bC9n0lM7/3zuIKx
RES4l+6q2aZ+P7tUWwRCiJTlnAgt+uythe1vsaqBqRbmqD+cdMncW2EniEYPkaWa
ZiLRcadQOyUjwcz4Ul0qRYBP91DdoRYu8fmyx2psBuaEYh1is6fGnps4pqsd8rG+
MQqz3BWSp4P/rayUZoKemw3Fom+45jLcEsF3oTzlI2UwvAeF+clabIMnWozvZzfZ
Zl1arMytyFO2YOqZZdqzSdyomwCFRa97l/M8VKEGZPr5oWBMYODls9us8JoCeVBk
NIEY0JM+QkOrCsR5W0r4yLQ+oirJdTOxy+lNF04Hxn2zN/Ixf83S+TJiZVH2WlUh
bwU6I+gqz/XHRincPlC1nJ0HCkeiYO9z5gcGGDVxWZV2R7j5jtGb66UAht3Lva69
FaEEAHxWcqAA9RNhRCkauQOGnLS02bhGtFEAPYBfwk3faSE1Sd6639K6VtPACI7b
znNoz4jm4BY2kzl/BsLo+BvN1QCImRC6hKr9wMzTfiG9KmsU3MKaUK/P04MTQZsO
jOha+/Qr0uy2sA6MR8eltefJrfpyNDEuCsy9gPCEgM/j0ACwYHl2je+KJfLujSBW
7UfYNNFCSkWGMZeuAA1GuQjjvveCFRVkeon2xwgaV39DGhrqfJdvl0ioseX/Y1v5
4TzkcdCPxS92+BRkhPG8BVcgQEAsJ/Mf7CYaVY6EQmZD4slqGBbJZtS8+sozTFxt
e7QPKrSLWFY0asnLrsC8aZgctmOFLoE5zHnUHc6n/remCM3T2FHHXwMhPm//desO
FfJdMWw/LcdqT8RZd89oHR1gInG5qBYzbbySM3tIBTW78FTT7IGHhMvzRjgGnpQo
t6WQKI5AXLSpbzuGReESviGywy8shhwg64DjWh7n8uNZTG66rQhP6uxNUrQ85zWL
lGwrDGH0w9mPOS+MmxUEgmHvt74XxGo5Kc9Z0IsVyLk/oLINJpi34coV4vSvYD8o
Q/2O9tvgYGpHKE6NPPaGTjgZKWUhgKJpRTdTBkxPng+Z7idmgaXPPLbJidhnAyOo
vlzK+aArVAYCpDOy2BqRH/9YgUnbQs6U9tpyHin8CeQeRum0PEXpNjOVuJUCfEQk
pnkNp+zIHwMpUcl35FlvoUuEqgchZF1AjSZcrCjWFt5eFH+MQIK3T4dfxq4rF22I
bAJ/8a3K/jx9bPlO0WDYybdNd7WaFQwvuy3qXhe75y7MeaaMfqaecsOOILgfE+IX
awiSpu0co0U50BSiA/ZH/dF2DEoDIC7EtfJDgKn+RCmmVqKkTKhWpph7a+M5StQC
WlbS1WEAyN21eCW0fUXYsonG2J2hZl64OUIodw71xuzorl+8aHqMSjF+2kchgGLJ
NNCrVzBv1iU9UoRuzKm/GauYIRSyU12vQp914sahkkr7vZ5U7m0iWvt2JUtF/Ahp
0OxwQoDx5eLeBOjFk2Cu1MnYDP1W4Yuw4jv05N8NRKcQVjrBtXrlRjc1Q976uLL1
k+LjDLb5CecREcSNL55EKzm/xXrDRiqM5vBNhNCcTDvPVJ+TWJxIRCG33xwMbtbQ
yzymKudIMwjP7dRcd2KOGVRhhMtfRgk4PNOAPcIpVGVfFpmYR91lXuYiizIW8eri
wDN44DNyAbpj/9rev6efWDLFhXr33KlJZuaN0GBVASCXfya9vHR+4RLVSfxcIofK
fL2UkENyaVn2DYjJ9RZK9KGVIei2+6bQe6uzMZwta0EuRsXfjN08lcg0d0uFjTb9
n4GUlXbjaNeexDEF1f81t2+OxjOCpJS8fRpdfpAJVR2mvLyPQ1YfNQJtLDNtRyik
WxRZk536TGobsIc9LfXobOFI9XcKhFVLV1CYwLH/8hh7pjaxOItPtwHSKI6EgaME
gR3xyW/aFs/3uUTE156NsLmN8vFkICjDnxBhSrx7kB+yeVSQJfDOLPAgGGqOaXS6
yLIRZqlBrvnNsaDbmLXRDLlzqbRdkX4n1CV9vLiNWfD5cer3ef8+bGL0VO/FpXqu
PByVBBR0IxqiJ4NdtmmAyV8RyE4sXth1DfeG/MX/TvijCcFfGw9rQFB2kdst1xuH
ryIepI05ooEPvXXBxzLbJN8I37RTEwXUdCZaOu7ZZh+2dXT8a+8/HcxDWopakFjb
NvTRowjzc81uybpTaGjxcpAczELJd3SPVlUianub4imPdGS2kPPLiOJKSBOJKrzB
Gk1v4F0v9+2RlfwZmWxdLpYooqRT/GpPjAaEDSUDqTfUhVJ1QVrcp/gyjDn41gTI
5ZGAqZif8SF0VR2RvyP7gc6joPZgYDJ8DpAwXSsTK8BAlREVY/3laQV9IENZe91e
1GFt/4S0ul6N1s15T1vuwhecgQgDwneKNKNu80U+y6Ls6Qm88SIHSAsEBLhgEEWk
9M5KopAMV9zdJuhpdUbdRFR7UC+9b4DSR1SeXtTTY9Ea7R0/NScpZUmfN+zGFRzq
ItSSUzZsqPYn3pmHUXMHnm/5zHXE8AH+HYR62g/bT+U54bLxgLkYJ2bhvcFlgche
BfJXY+aB0cXzaDwp0/tG6/7Kb1mV3KFdclPsEgw3HW7lOMpJYW7AbC2uLrdPbwAF
gVAJann/SH2x+a+QuBq0qf2DD4csH5OUVBHVJc7u3nJzhhuYnVWeRpFyohs2t/kl
PSJmL81zzmbmdJnj8clt6CxQ1VBmI4dwQVOOWHuMCpgGHVvpTUxrzya1AaQzXnPF
BeYf4nYkzaLLCF8RrAGXhqojUMfjDCzDdDp2kC9Se4rCrHs2uzmaujVvSdxGMCCE
DQymkyChQPrBTJ3wl5xTpY+GmmUwTeTUdOrkRvy3/d/K0Oh9PTOwK1OWEp9fTBN3
Nl+DkcKzy0eu1eiXgGmKsLOfNdLgZ63u86nCZE4VfuxcVLCTEUc3IaYEWYYI3Cy+
/01pJ4rNZJOyZvZb4bWIwBT73GRsm++PLtB4ZaVWdQgywe//CBU7vLF6M/xAjDsI
rCOyA65Knwf2/e7KjQLZKbd1xSZoTmVkJYWoEnkucY8BsfKAQBpIezqG+4YDoHci
QTmqcbniR84hfeDZv/U/Zronz7D/j957h3jByODA60YiIClYP/LKcXKiJAsUXTLE
iThTrB9kVzjOPtJ1FnFcjEvxQB+fka5zTHsHNBwKkP0B6TEi+ebsvTazpNpkhfUo
MFCzmchHpca/9ts4k3F736NKX6H/8m5BABJOja1qVIB8yVG07JgGVk4Gkbgx22X9
Gfdx8Yd+X5xtbr+BsEcCcxlCDHMzO8oUQfPUF4m5cUT4/XRjjWH/rqa+7APXroPp
4s1vUScJqm03hHqkCHUUW3RgTNPVaQgDZDJExiD6ddlaCHULoN8thEL/U0V0u0Lp
DsbcraP6wpWCunjD0cdajPp7zP8jnMYLowK5+JTzkwgRVRA6jSa0XQ5Uj5G3ocQG
M6w0MT3NAcKV+fjfqS81d8E+NPaixO5Vsrbh9FryYoTt/xrzZCc7GXHC2IKx9rWR
WP5X0DQ2QihKng8kvaCaiwzR+aNH5iJpbGW8KMO4EtbyfCut7q3KeFyOFTBH942c
1wovjZrjydQ77tASVUOpBXG85AVtMgT/gONBwLqXSMCRPBV71PBz+AbA8aGTBt+2
AEbfJYB+LJpnn0scshg3WKmMbykskLlARYCL1nkB9N+LLaPkdqNIhajL9HuJfHng
Izx6FR5/Nb9nKjp0u4PPFsJlfeUce8R9BfTgAKImY0uwCuzwkiA5FXnG4DhZw4xE
dvlYQsBEIXJ74E4qeTOlFu90+pIjO+Ut2p/ThLz3bIK6rVZ7xuUZIsoYgw/Efm2b
qhgPPvTGr9x3jfwTWVPRmQIyKK5EbCHl3wpUHez9eJLudHK77NZzBxxcDs9fn34K
wRGjjRbubgrwKFihfC7+FqDWnb01U0Dde/uQkiq9LCPxkPdpCb9bcHJjtahq5FYp
Mdux9D1gpvXc9c+OQIomST80h+tPA5HmJ+ih9vY83RsBgQ1Ah/YORzm4gCcJozeE
wPwp2DsNXgymmGeQvVbTL3l8G4mbZIJ8RtzBDKGU1TDNie8HhuXuiwdL4vgL21dy
cc+VRY0N0Uyx7woJvCxH5QPVBW9+imrcL86y+7J0hMMm/ijDMwW50BSnzOn3H1EZ
3DGNNHB0ZPSC5XgV7Mf86MT72xqs6ZqY9pCQcw+6RPBD44ACZxGK93NBhBzOTNLT
zDYefGMEEtRDlP2GBg9ztmXR3bz3Od5rknakb1HNgx3zLx4BGdLPXlgmtWUSkBx9
sdLUExsmOGVX8ef2c74rs1Tq+0w6G/Aim/CjIu7NzWAA0uFVm/4sKpnJTQIxUBPR
HnAv5byCjhjPwivccc5jy4j04hqIjWQ8Gs64CTtmDF08pmMxPHp5fc5cMdGLhXEx
K7lC+ACCDmuLrDJJA9Bpy5LmtUojHp2RmRhGtqPwFR5f5yto01N2avAkRpvSU0jr
kulk9ctkKniHpimBg3x+sAsOhstW/jiQP3IKCSEHpza5f2ymmAJTZ8KNeUKgYynj
wxTM1WFWExDzVd5V+ze3SQburf0w9SaRknfbNFwSSo3G3Sg9+Fcy8Af0HABJtH+A
ScBtPdBnW6xK3V/os9yF6yis4ItHQyFXH+RZiyL7W9CtBrvQsep4Ss2aawEVlKnb
He3hJ0SS8R9kWWoYpgyqhEakyw3QltnRo28NzxB/GcQJfn8h2WJgttLaA5DXsQ6j
wpmmU5JuwtcyWbPm83t+4vbyjHeDvBPk/rfg+Bb7Q0EmzZD8giLuL/EMk6kV9Yyb
yzerFNMou9WH7ACPhVhVeV7Pf7Hex0LEugQhXXq/GuijShMzDkUe05n7Qz5EEUzt
vouqLecbVu8Vtd0Fg65yocV8eOwvXbRv9wBBtZoDiT2JVl7cU6AsZGKaPKtD7H/w
pO2BYYVQaEVbu+d7EX1xjNMGVrUYs3zv5cIZLmpxrfoJ0Cb0uttjtUGiVgdtZqz5
DajExsWkRsK5acuv/H9udbzYYot1lozwLfnqugS2RPBimMMbe2cMQ99Yto7Cfvxz
x7dM6WeeyC92ySUh356SD4mR9F922VvmPZSHSI45OeMpVJ+EFzmC4qqYl3j04ijR
ECMiT7gQhdBUxmox07Ys3P2Pypxu1b1DnoAoFZYoefUW1j/6LeLDjJA6MkbiIiec
pgQo548R96h4E/pIrwr88IYD1G0jSQordREmDXBgxxeO6GR5ObdRkNdI/CA5o3xu
iDOTFk2n1lXvRPOXI0A3Gua0t7k+o+apuhWzyUYST5sMhc6Z554IlYayW0DrREEb
+KIuEFLKPRJPyYaqa2K1+dkTtcPA/aXjy9xn9HBcOcyTkPoYo+v2cpgR2dj0J88o
aBCamTqtu79LSYSYkXaZ245E+4l4deZVDeKwhSIiUzJjLi/0FAOyPkOxFZth/jti
Ziu1yCp/6e/FQ3UxcecQNIahcfFJPdJrXYkVADiuRoAlZpF5C5uRs3N4iWd2tB8k
1O7S245o75J/XaVObWKTrOsz/a9YcNYAjq50x4RxdcMa46Z8WYebSkNuqI29Pp5l
cAxkCaY3CyFOMpFG5PQH/+aqoS+IdWljqFTqBcmTbi0YOSQXTPPkuIfuXDDKP42e
C+JsbHd5PvlTwk+uB0tY2OklOy5vNQscG6ahMXDf5FlVNCvkwxey8UrZn9hlRa4h
SfjHrjt4GdnLd1TNRM7TS5wCEKYIIsCIZH4jh7T1Q3K1psd/qWaw3YubwsJ9GEeF
91YfFsLvEuPHuGBqiOBujZEh72lDknxLashOOqWYykWA5AZskoeSSz51+NHnZS1N
BD7VpoDbey4F2XksUVjHcdyEP0w2jnD9q14x4UrQAzr5K1KbXpbgrrc19sG/uJ6f
cjITJg5mWO8LEIkzhcvjoGmuBMO7wTZtRiMqMqWkTP4QbLBn0nAxJhHOWGDu8kwu
txeYz+Mycof7tZg3nM7zaRKv6VYvDteTrsfoGg+Io2uuQ8mDBppFHoiWYFbUhj++
9x935MjIQvSfDCLnK9IA+ilwWmq8ukxizQ49BMVfWA/hwHf61DhuPL+llqKAYt3w
otIFN4X5xbg7YwhXE/i6vegvj9j5+I1LLH1WeXYgHScnADI6iCIaim99ugnsDG0V
YNTZF4HKtyk3Ldc695wIwuZBRAzpGC3wrQyOs6mF6tY42iUh90XmQXHQSF/jd87e
auOmmEBrqqO7MwOKuVHvFESYZidrCtlvw13Eoktc5v6+dvmX02hquBnaM3yRAXeF
BmWLrG8K44HNcMdKBAagI/lcN0qUCoBjuo2Ww3S3uCXxXHr8Wt1cFoLaOdRzkKVf
LoEJ6z8K0vhRSqCfFIzVWeYGpGBMfwm4i3g0cLhH9sNv68xTtUmDPsGbMUQpw0WK
n+Xt3hTdig4nP2AFcYkT0qXHCoHITodxEPdcHzWVAypWZgcTyCfk7JZgvBYihfV3
daox6feDhQN+Wzmneei1QWt/3thgdY0WK0vSk8Mw4Dws5CrBhlWqvvo3bwZZsgdX
+fOiuhhDM2Xnh/xaUVDMSAn9Xut05k5EPSIB91YOfHrE4oqvamlH1bY5mKsEgmuc
EsiPGLeFAioPhuucLXATfqR8bYs7SAMP77ghE2grun0nyEDRBxrhmPfIGsEk5oe+
NYHa+0/bAYQTIiJdYL1d8mP1LT2vOcIjSVyo75/RA2CrkjlveWqoua9t969+wZ9h
PO8FB5bnbXatlIJnEmRyqbGwKEIl8PuLwNLddzCA6h5x9I9wgD3wYTLLYDyPRL1m
nIbEUQ+Yx2i2WNA+hBD1Fo5cGRfi9xBDBpiCUnhqPqYmlWCN/+tpgwmgHbG4c4H2
qo8YfEXnW54uns1XoUufW1n6XaW18UNbwtnq73d+CmVviIOlp1N5PvqmS7xkNxaQ
dY/aI3llE4OAxi+S0ho8ifPRF50JyqQQ/1rEjN+ZYouipJZ08t+i50yyxEyNcvJ9
QjsHhJXMcAUv/6wOKUp/Vn0zhSi+rN8Ju4dHWoDGzgISXSqNy7FiGNC6BDTRbZXy
RyRmjVm6eIQF5iNkcSt4BgRjvpEDj3o4IK0b3mwgC1oUhzF9Cmp7gnaQuQCwYVqm
GRvvXCyQ3P2tzQ7P6NTY1B+VgzBHgrskKDOGGCIJRpk+WlTpPaw3W1VsTSPh92Zf
xNNCPkn9n9tXgXmkYtcg3hmPetMJWjY3wMVfs0YJbpk0zLKkpKuPK79xWFr0o0tj
IkQbakpBWI8jhcmrlYlP2bf2Oy/FoLSiENY11sGz7h7azsF7HBvm44CZJwC40sh3
u/bW6PYfAoEiYvlG3YOc9QihHDLUViOdpnze2BTS+QQPC3N93tKwXdXE9Ud7q1z9
e0HcPEzcoCRHrw0edQA4V1j8Dn8tVxVRhQ/95XoUwrsZr0nshRBCMYjaAzVO4qc1
2c3lotJdneuMqIxBmpiB5rAuBqgSfci7Sm3YosTvHonHQBD7wZdQs8UMQBRbpkxa
eOGVOHNXLvlBaNcRqRReXdLLmqxy8gG+duSYsQYQrUdBeYHBfdrIw9eoew2Dz4LX
eJp2PtlJeAg769/ilGTwC9klBpPI6u+4de0g7XqKjfNZjGy5nhw45WwLj/+LtPoo
UNyX7UrxnotWQy2M9AjaEwPltpkDtFHdf/Oi3k8urFpXcuF/jicTyU1fkR9Nw+hY
Yc9GgKCoxUa8gmBYoV7U+uaru2pIUtALFvFplgLOLXzQn6CQdmZZpEN17l4qHFv6
rEkCK6NpwSkNYKmasY8RwCoCu/OVqTy5ibjUyUFqlM354+t4JGy5DZsCdo9qdVe+
yf9OH1dT710j8D0quzrvsvb6Yv92RXGDnhstzHZkEegKyV8fdrJ3IqqHNQoP3pcP
kX5lvIAUuBBqVaafmxPj3kaEkELLsrW8vLOG/3A5ysW20ha//F9mwVmIz4GlZwtS
Oix8Hn2PTqNGVraoESeWUlFMnJyvTDUhnQrWFyGygwFA3MoCkBkqNzTJ2+7actHX
zaUjEq9fkjGIMz2heU6lyo2WFkIMUb8J9x7Q7m9ZyNfnzHi/4qwIBN2+6aOuCJLM
kbcu0tOej6oK3CRPBnoFjpiu0ETfLTJgvjgJ0sEjjIVcl3Kblightik5N+SGM5UD
RqlMFYzpr7iUFANy1MXMUAH4QtVNN4FXdulDse5BpXpXobAF654bSBbn7JGOwIFq
sjYHX4OTcX3NnsSkNijcXT5bHvTnlQGGsLMVPJqbxys2LDorUOIBh0mHXPoyHeOe
pJElwW9U41kQRmNSv8p8vM0m178xArMC0Blx3NZoImsiPm1qr6cSwrkSCCUWiVYR
mEKBesSrhBMnsepRihGg4DnfWMh5xwFV3pj5sAWkC+IUzsVrZIBAhfvi2DbrZJHi
aRueA6snsfz3cj/lvwPp8AOnZK8KEtEbq5PaFFFQ1kQMub3bQHWPqEqyiVJlUBNH
KBOJ9CsP6jdWH3gVi+l1gHeig6WBHzXprx3EWwdxkF3l2oL6VK8IyTUxUVovHNEe
MEZlZF5JPsGezmkorppufp+JTyURG4o77kIcZbeZgEcRO5C4x9+gt6+A+Y7kM10t
R5a647OOLh/My0mLTRUzV7Qsvg3pbmvVJPYen6jGbP8snGFE2XEBp/SsDw3t/Gcn
UIo0oVh+xlLI+4Ht3QIPvgrrps7WzVZBhGSM1/Sua01Flrb9bWDPilFc1VhSaG3N
qQ5YIAZ3TKKrUD7crdecu3pYSh6+GLy7UuPcEHaOg8kavv7xTnXWSPMYunpsYhmS
r9M6yH+31SEjlz7mpM3LW1gO67i8bnsH7SHt93/ptBRo6AHluTUsqbEQkXofgLQJ
C4WDUiQt+rftU+B77N8E0KkekDzmlFd9aRfwjmCtqlbqBdjtf/RWdWCSdOvjOPje
fKSx2WyfeMLkTpC5RpyzWSR4aGRP5num7AJ5fD85SXBo/L6sPekYuQogPj6f+CyZ
Nuy9+WPrboPvFvWWTX6Z050INqerRPTX3cjnBVsgk6N4OgjHkKPyah9pGXXcvLfq
l9yHm2IhjCN4Pz68uGtiXysC6M9yCzAYwq6xT8BnlPtOIcRRm575lR/fdKo6jPD4
D3gb0oqkhPk4cTnIbOBbcXlQN5qtWcbmedeI0BMaqdUMoszQzQFSZ5qb7pPVolQh
SNcxhMb+Y2mWCaxKddaHliq4lAk8KuNkw8R9x5ETgzyo7WGN1jgrW8vdqAgIKOeI
66iK8mcFa7AKC8WrtteCi6nftPPsSqblnZOMJ+0kxUsXV7H9MqnTZSQyuQNIYk9X
MFvcmmDylLd8BNZofbWfQWmhZPH57yFmItr9JYDqFz84N2m/KLqklGZEQDDrNluf
kP1n7aqLP2L16YKnfUkyPk231XXtnx6AouUjC5Gi06miS6ndldDZB8xBcXWxjCkP
pOUMsFToeguTZXKQbxU82YplAIPO7rfNTy3oOANXVcFZXfvU9whfa93Je+l8wd+q
hTgchdvW7h8oTrmigkSVrp4tMNJ+hsnq4owPY6HoT9fPOJ5dRkF+lW7mIY6x9Ppk
D+QXahBOag5PZDeSMQmNiZq542g39rnzH2EiC9RJw5p/pmcfrKbtdREMMOR2bxH6
U0LzrFMPIT5C3If5E2z9J+eAuNGvlu+7re+2StfBuub6Tks9qEROkf0ZPBXqcmyr
Sv6V5n5B9Pj9dElcfUxUUddkK6OhcOr2ETEQZY3exvLzUXbmz/u6ZJYyC7Q432bQ
fPELLAbF1OJkXsC2/6Bt3kMCKTBRrN17+LgiQfaQAMxDDVBSxa8JG8HVEvMJOJ2s
OcFgVF4q77nGIFudPkgEJUno5Xv+DtG/BZ+YUqoj0G97r1/pH5UxIs5VWUlMPvp7
ac6bnK3+t4BNoFjj0u/vMP2VdooHvUuciHZW/5UOA50UhJHy45YzYN0MlFiwaFAT
J/cG/JcisJ9GC/0iZcFA/0OZj8Yhh2fW7g8V/Y7PPYFmoPQ9yhekqociVRdcTuBl
Ek+h2V1RyvIl6gTl/yvqKTxF0d3zRX5Q9VjpA53HNiQFH+XU0H2r5eRXpUUNOtT2
SvMSO9tR1Y7J43Vd/1/wdP8tbSrYOzrV7y97KA44IBqow6VPqZwACA04X13+FN1T
1IZYW1LcY+pAxkhHwu+O+4uRUL/gM49bVUnaRCXxvzyO1t6vM0ul5zOjyWm+oSvf
cnzHYEIYpHJoh+L/RqTlxXq1YccnNDxxdl5/Q2sh0Yr6wzOVSIcXKqOUVeffClmX
aeK/AqE7dRm3Rmohgvfuohh2M1uAlhaafO5OQHuUI1S6oDpv8MlauqLfMQPXu+Pt
+xroh63z/XtaBcxvM8mcm9o9GPkNSsCrZoHFK1a+qTXsT5jnq0UTZHjrRLgCs4hG
vR5plaQhaZIfPC4LGx0/DnFvRvuPR90vw7IiOmQpeVCjAglYdNCnWkWv7mowlAir
sYVI74www0EtaZxbUahExXuXQ42NvPGQwcZl0s4VmGPagVIv6DfJu+GRyKgWl+Qt
atVGkmfw9HG7GHuUNS+2bS+hqtMwlneSGoaQhNv5cKPA1uwPUJQF4JnCJ7B2qGEN
QAeaYfY1mNufN/5dpW9azvkeQsP1zJLrw3qor7vtCQ4FoDhnPjw2w52x853PpIsx
Z4xaJaTJVWc6DPA2pUVmWwF1Vh3zIaLJ/8DnwsbFkfYGUowoLnVSymD4ZdZns6il
h/ollwCA5mIyF+8k1DFO4U1jX2OqLurwt58tMPH3Z8cxg+kNmJ/ifie5BtQW/6sX
BtoICJsrzNWB8kxNa6ZP6DR0IpPH5r4JLsgu14EBFu/Mi05z1Jg8bO6IoZl6NcRB
sugRtnVcEaqeO5IOms7ZkYeKPCELfqcSbPmHs9Frj3+rwigOu2BuGppJLSqtqn0U
b5pOSwEsXFXguY1BB4itD/eMcCmjTr6LlorU6f18kaRANDIDQtBTULDcUAuDBRUy
YJEQuWjhMKFclVGgeXvcbrnUekLHr0ZhPKmV0Ey+DaukKUSKgAlgfRJAI3COOGJ1
ck6ipcOMAh1dN13doym1QUWs380CMfNk4IB0H0q9cDLRMNLvhR+AqvrHtRcOBqpU
jccgJ9XzfyTMdk69ws8Hw6OvwHe4k6WMF1MXb1RP+SQdkPkQMiY/FNMdURpWxKU2
slmmGYKEH9ux9a42t2nxwCQLeesCVXsSVlKPRzAXA2DL4PV7xbsyYG1T9BT9QQqC
1jBKDU495Wq5aRLLn0IY0PpYsyaL9qPjrtQBeIQvzxHHqyV55uazyqeGfIQJADUS
tH5zyQ4uFVCwGIliGyJE/DCuxZXucVGYNc711le2cLX+V7vll6/kSBRiT7t1rRHz
tm6XujZlbM+yH1oJ07xkpy/6C0oTr64XcAtyrdxuO+lIf2Dj16BOKZDLFWu0KIsE
GtVHkHToQLUoHVfSMEVLVmWleHQqRzdvLAQmg/AzKGvCcGQV9kCaVNFYtZXMTG1d
fYXZ+Mo/3MlC0/BambJByYxGxzxmwwyMeXOv9gdYfeqnVyVzTje1Mtt/13WuzIpg
MfyMcJkE3kl6DLRC2d5UMHbjGVEnMpV8M3P0F7PQ3N4AbamJhx1sXnaVmlV19B/X
Al6JMmDYJoMv8TniVgZjISgJUMWDHizHUF/4HhhtswZZ5ojmN6czSGGvd/jplzXV
XIzKbjWzqh4rYB5vw5seIS97R00vJ8uIZLnb6s3iZ5RXfSnLPZLdKx7DV+7fogn4
THAmakBDjXuu2nvniNzhuy1MXMGhJulRbo24rt0gfoPlKEULWDoeorLJ6r6tPSwP
1SXHvBCr5IY4Aoj9xbrqyvl4ezyNmJ1zc/uS8BF//mmddkg2sowM5dnX1utoHp/r
2rIvDRXqNMFJXe6REWMOluZgT9DSWAC7rblgh8+8KnaOlxQOhZHz8FMfkc8pWb1w
U+fgaIo7Ykeek1v0VDS/3+HCd1iMiKAcqRKEksZM5upHQXCmHzV8dH65Z4ksPSo9
zmNHVd1kHm2Lm4H22Be7kMFPmJwfUd+e+2A4IBUsDssBObZRuY+HTrJZAs31DMQA
STcbrNTEVqbEud7cZJDqSVDkJWKlAU1Xpe1C9UBLtkjs+TGUo5+6NbJ7/8iTtvC2
lQM/6WaYY2O3rx2Q4wVW6pTGYiGkyxQuAmbHYCbqS5te/pCZMtKNsnBl2HPLlPOv
HUVbJ/o/BYeisljX4K70Gn+v6aIuGl3SG81ceUuvqX0yuZWEGz0w6yiRJJdD/OOY
3ck4H2sTFcwGR4IgpKVKxWicuZ05EI6E0+jJv0C8vIP1HqpHp6D9UkSVgJ4gov4e
eFowFMtJguyP+cthey9+7EImpIFpSrUssJm4AjtdeFxa/imw2B9Zi7bMKd7o9Bq+
pd/zM7+F6rkSXvEa1sVwh4MKvB2k3bR980dyiaB3pw6joABuWckPA5B//SHRV0g6
owdB5WhyirqZ+4+NL2rU6hv9IaDOwfdFj6MXz/brHACQ6FjC6CAOkAbT/KBBgQkB
NZJyzDiOEUglB8jp481m+eGkDhTDKTLU2/nKy2R/UW7mPL2f8QDiR6iUWQB8AJCo
a1dMpbYuCnSCduc8ZroigUlWlZT8y6H5jcygybHoT1H2zvdOngfJfLAq9HpRitW+
TWQvjA93PdUVmsucQuD6LR/UrCpCfbacTwhcXN6+I8kRRn7ZuUKqMGDzFnuD0zRT
7feXlDgocMJWe2SSFi9XAsTbON8un8MEVGfRuxXknt/vYAfyZz5PYTfu4EZpFMM0
J70t56BdvgrqIoF8kNlauhYqA9UNUF1Pwd6WiMw+8nBROP2EhsHjGb98UzhrB6iS
3nZ+NgjNk5PCayI711ItuVqr1lej8FCsEvYtrYfb42dbnWYqc9Wor+1T/Dg1XURr
LsTuxIEq4ndXZwIVUgPHycblBiTP8wqS7sLj8jf/TgZ5uqe6+4IjzaLuTt9zqlLH
D0w8iy/5jo/wuf6yQNmBUOvo3AqMHhF8e3gEvaoeE3YJao1/97d02g6xAKTh6Moj
eu0a65E5A4ymj1mhpNzfFPr7c1bEAWRrwH5JF62U8VW65mR+dCaMnNpyybXs21SU
7cOginTjCF5ft15PQg5T5zhD+cLa9Qk4JKf/8RX7/lAvW2hQfbYl1BOE8Bie58Sd
Ry+g7gabjXtZ6AavDTlZ4odxpMikoiruLuMIV7t2uhAKyVCPyXzcno+7Oy71ZyHQ
IxRulRwyBjvp8Ge/R3QgqDUElsnEmsOIGOO9gS/7ugQnTFY4XN/bZLw5Eh7q4UBF
JIdO9LB+WlMI+aZeqz+yJ86QNM79sDiMC7jum3dbqQsQI5ClK5zQUWClo/QKxfx7
TbkZcSreJ0tlzjgZetCykA79/Vdo8UlIRaPqtsQxWF32fuincYHlPdwpXcCeq/38
EI3Dy75MGG7G52JktRj3qGD0lNvnDaEMpqDCwKBsAnrI5C47DZCAubvErbpsq1+e
sqUUD4aiVdL95+n+9GC39fZvYVkEL7b2RFSamk0Tudi9R87U2oKvasHAoPnSU5Dl
Gy0Irxuyv5x05RNNEAfBSwwr/xu3LrNe/5b4PF3IwdVur3u7o/ieHDTCZqHKGphN
B53ZMeDzJfP3pN8gkILKWVakhQb6bclGZfF6GFQ5RIuEQqp+GwZGduoAABwlbFbq
0eFTcA5vPQOCG0Z31qLukk7ByBnDWd5OlsTuj2RX3YRTCniu8FHsg7Mu7Krb/oTh
xECuTLohz6IYrJcVwNTRnpTBY7Xoh1zPiEja7P0M8z529oXgfwZEfINs8jknNAoF
217Dra3ncOM1JleP3k2lpIhah0ykVTV5inPSWHi2WXkqwNgQ9TzlzmwWYfV/BIyc
ugDKlxs+a/nQWOvDszIqfdNsXvAAuTrvHF7C9JcXv0QJaGwyYUutdt7trhYadEcG
qg0Bb0lExlnLHG8K7ClO2r0pkV6G63SG1kJ41WxCH5Q4Q1lu1IRF44WJyYUPhBXF
lKAD/djP0+YL5Vb0STMmCYLZXHtF0Meo1vS+mR2gpw2J8vffVEDXXKUipxpA0hRQ
bprLtaPZjflL6m/7Xqn2jgQ+nXcAFAzDIYSUFwCWB/Aq8JhpOhJhDHRfDmt6Pp2B
x+7rcf1DDu4lzJXCNZK5q9ooC/UW5yWWMk+s0Y7cKciZkTJm+gRz9yubke6TtBnN
8GiVzxcZsltQIiJydL2re7x8uiSm0B4AMst3aLkq8DVnkbv9Bh4We7G4iqZSr/7d
lQXaOwVqoykrZPkkCP0UmdWEshV7Q0+KlOs9qbFsSK3jgukIIk4jWfLDegjQ8S3t
6G4nL+qojy5CrnZKeVCpIBaZY6omprAsFqBMKizYAqiRF0cgL2R9oYalSPolJFD4
kzRnOMYjZZHUdLrh0xnzvdeGIkqNwy/uIszRvazBuSdV7LHTzSiL9zXIU0N4WPH7
gNfa9aApnfZMWXf/GLwedQH6dqZYw8eeA7ZZP0QfTHPwJN1tMZUrqV/hFc84s0TG
/39fpoRXCHP0Yn7+782mG69BDH18IEQVyk8RLbMzJ0STs1XH6uwjXcMtsBOOp1Qc
WpiHAoXnsxu+lKXnlvVTCiM074SqaJ3+WGNPJDWWm9l6evn7GiAvH5VwcQCAz5Fd
YxUwmZPEcgtZrb8/jZpJ7+V7LWFB7s/CbV1ml+A0Tva3q3LWey0H9trDAfb/mrG1
sRlm09l5vhd39YmAixxc3j0NjefoHWB+f6ucFOdzI9zF3T/JXIlYVJzUtZxQnXYo
ln8dcI6fDx+j6GAnj60YxiCWor+Uwnt/Qu0DM/7baLQU2jJ1FSBcoDFoQRLRdNIb
v5lyevHhMoKRFk1/BCgZ38/s7MSdxDBPNopZsNWCmiGNOxuhdqt3CVYQsZkvqIIk
XOaMx4snn1MKBC6sabTBlJPUWA/0srAEA3QYoh8aj7P1rsflvamrDavyFlB4gtU9
4VW7ttjYfinc+hEERTjiWEWHeMdY/WVe/5S3IOzw8goNi0vxgPhbF8h8v35D6Qc8
G180+j94iU5HUn819e7nKc9GYVjZb4dG5T0ehG4S8QjJZo+lkwyMK0Vd7+qO7tUy
3F40Ob/xukuiT8Q5tPQEd7bbbxwDkFOSPzFAzGLlOgOew4/8hgj+QqyJ4yptzcs0
fr2RpmLZDeCq1/FyNG6fmOP2r3HFspaaCB25R970dvufxSn/Q7OdbKf00FqhMGFT
ek/CFncC/S7ASYmrKGNb4bUADYfftBOEwyrO0u0XGpvQY+H5fSOVzfUltqzPLbyu
edwDI3gAJ+0I4I43msz/W0RcHQHKQyZ2S4crW3nJL3mo2kqnI7Vd5xGWqiWGkjRd
qwlrVNfTf9czZGvvKek5u6Q5TDw0R6I/MtuI8WOROHioduCcL8EdpEMWUZwXFo92
D5G+cFYAm7Mo1Afa+Xi5Us5oxjWelEjVpfvtlvrCqeDlBHbKGXXMxTlD8NADxfc1
TZWCfNXjnQdsrNVYOPycpDfeBDc2oRjRWUzIbsaaffUi5ldH66Nrtou+7Cnf4LmM
cBAzY2rSfwfcyMOMT2CWE5UQF68NOnH+nmZpLNnGBR4lJ9WSBSUNZ5vD/brHqlA2
hUGcFJ2/1bu7ICFUBk33w/YwLuWn6aXNzWdsxz7Lr5lHw4PTIctdknx+pqVuNT48
Fl0QqHoUIhaplm/J0ON1jPsCpYxf98JXGnvDuxHfufPy2FYZA970K3o3lVyOfKok
B6ZU7JymTdyMtxepjDpLeIpx3xLc9N5m+NKdKcmHwcfqBHSLCVdPIyANt1XD7IH0
99IET3t/GxNcsziV7SmVdru4s+O46HA5lwzIl6BEn6NOzAyFHC/Qadow9z4MpRTr
8O7v5W5SrIDrgntf9zAts/c4UIAxL8nU3ncVqZuv6pZCK5YepgJ4A86bno6Byn3r
bLK1iQcbyIw7ewmNPcbIE0S9dPQaERdntTZKjHOO2A4wzalZuXxI8EJTXCF9FEM0
bRhp+rsbBKFa4Ib6gPhcdnwDuCU9w0mf1vJhceFSpvDmay6QyiA0oKU5iHTzT5YW
wjNJrcibxPhO2Nfrt3oF53oKzPvNehXC5tqqqlaPMUixSxAMW8iV6yqAPkUvsq26
IMElhXs2qKVaB0CBw8I8ipvaBklkqKA6B93Z2PVHag7bCuuhKy/3AS60PwIUwVGY
fY/RkdSOKJkZcyPT8z3NuHZk82iE9sy5hWRDl5hCxPwzX2yhm9CZggGIGlHn/ETE
Erkxu5o/fi12cX7f4f3vUevv9QTRwzC6XRF5xGNIQRsOiXTt7FUfJxvKraK1g8h4
8RyWNpdC2/xksEGcLPippGeGA9pt4AkzGNINww1Gb3F+HPXg5Se8hRCmeZKyFVX3
JpMAwTQbZikypP2j532cAMqbidJDwuuLCXms4gmAvgX6b8MBgBGx8M2JnkGBDYPE
OPAUnFBsfH1uZw7V1ON6pSyMvXk3srIUv9QVF3I+e2wRgRNsw+0XYIzwnThTqBJZ
OKBPGKmCRe/fC7HLeH/2RwzCJjqI7ATKflY55+H62mEaw4qh/Zz+aWV6k8u7DF67
V4e8fiBTI82kU2XgAXQny3JmilgEFzolh2aWwaC5GO/Pdp2y/K2DWauKWei7f9kX
SRpNDucK4ygsY3x/d20IU5IbmSSbAQxU825V85ku+60/lnmAKgrOdXqRw4KyHhk0
aWc4PwvKuTfvy5AIBfVM/RojBsPZi1+9t8AJiZkQJ9K3PdVWEtxXUqDkvoyykKZ5
yN5TDBLHCYQEZEbujBMpYz8/f9IHJ1Fy1Bf+x0y32F9jKzITReINNsbciN04HdLl
sStUcPT1tCQbG/9hb3qHVMBg54EavJkAdZCi/nq88M4+jfSXr5pKnxzhYqhDbzwb
zlGvbBp6KC4Hso+9a+c28g9kTTgpwqG8ht8NX+pXz90bK0xuCCLqDioMVuPr5QnH
zRUd1vKSYfbCbMo/8shhOCw6kLtJLaUxTXkW04ZpVsdEg3aCSMKxFuf8+2k+Iswv
eLDYj1v/Tp47PYdphXu7F9z4QxpGUAK0438qQQX11gqUUzyCgiOnwpablHLohpty
RJXSpOMy++IodGB6BttTLE9YDMOUk7LZSwjppAFMcm/9EBxjuZDFMiwTI1uaCOe9
Mp/OtrTY1l1zdhWDdHu7DAvK2/OR5fjaNP6wdKiFy8Tij8RtiifKTPMjQX3UdxpI
eC0ImTg2Wi6yA90N09QL8a9JC7ujrE1zbPtRnVjH4U99TFFbt/x1UWsU2B5VhALB
pRWTfyUNP255Z+gtDifzsGlQ0qqMWY7VhCx8hvVoMXiH/uKetJUd35MWfFKIUwOR
GNlN98G/nzwWshgPwhU6iy49QRo+8QGn312t8lE0kqFUHVfZkYvdUs7A9h/CwYWZ
b5298Pi6Mgs6TQGwg1vDCty43CkRAxetQIwKKd9lRS8HAXoDXJhB8W5V7+JjO+Mw
zpm86x6hO9UDSoeKuO/ngp8SKnOPuytIybyaV5LWBhSQkUECTRCQW/aHKVCHvqRg
HtRGlv5Taskrzabjy4di8Si8xkGwZapo/xS/Lo/Njz4CGUpamlV/uXTu4OtTONH6
0w2DlDXoTZ74B0YsAqHn2EfZKvgfEZnh5VByxNiMbQCam1gSzha04INZFCUOrkiA
uqeiUjzxuXu7VgZ0U9LrTKXu1leaH/2MjodGz6M+JO7rvOX17R3eOsAk5kP1mu2Q
6hYhiwhM/bhCnOsH/LLwpMjaqTwZ5TWY/hkQeONUyzom/S2PwKxf5h/RHNzJOzPC
FY+NRyCYm8DpJIMNA1/WrvqqHlWMiLm9gZEgw4p1h0jAHdOqnlUqYRaifPJkMyYl
UiVFPk5atbOEn/dXO+lLG50XQSW3eA1XoMsMXH0tsdPRO6RbZRZe8G0nvO/EqiSr
BVkhpiK7xck87VCD4rAKWYZrB3XXWVOqJd2Wvxdx/V30puUIP5ITcKLMLwxi5Fm7
6+Ee9QDU4aI6S7NB87+zpI8xgdrZSKzmvEcQhZ8K5DabCXOVzJAbufUl9CxaF8J5
TVnYak/DQZ0cUbd51tP2tjxNtzCWiZE/DNIkpNx87mgBehw/PrsdejCG/WkqYzYt
x+FskZAIWmnQkMN0+u206iKN7ZNtbzHsVK9/+DvCaOzz04aST2oyJHq6s1cHJcSs
uDR4BeF4B6T5jm1BRgJpaOLrBFwwrpqyr/o+vFjz0UzB9JYVBy7645s38eZxPSUv
bernFG5iVmyzXoUCdF7tVc/iZiG9VvdDED0aSTE+8raMQN+vCDj+uatNitRy3Otr
b7PuaA1d/9q9zSYFLM77mXq+kTMut2ei6Xw3UFm5/qYjNF2wZTiZnWyN/9++gNa6
+XBKMdMicjTEbfzVTmwirZ2a3n8gKcHShM2QhSleeXRz10JryVWH9/9ciZwC6tyn
U9nOICXolZbVvge7sf1JlQpOxgRHFKmkA0/TVWg2DH23ideMyB/T6D4bvdKD+3VM
iRRdB7qJ95AjZAsiHtrWr9TwplGBbKkPT8/8U2vUCnokaJNC/N4Z34fD+SuFXcsi
XEIDlmRhHO2vvOFi+rtpf4MEon6KkQUY2oapZyBgow/Lrxbfd9PQJrIIHam5FUKv
1uEf5ZSXzRiqRFWVZd7RcaW+9TAusb2hqsaFEfkPNnf2B5IuhGQqncjbaBtmGRcY
KLRnlXSitDMNro4PtPjkHkBOKwR9BbuE5SmGHPX+YGo9kB2CIbdefwBMFqEjeSDu
V221pX4TczPknAJxYg+eERn60BaywKJlXwgnBBTrzYE8u8YJBXbQ7Rm5UyXAtAJB
SPe7Orz3NoABtMeEjEPT/51C7p8ohq3iee8fGsFlGm+Vh2ZWKkbBcs/hT8mrCsyv
yeAIVp+JhiT5V7zIibYulLPBiruXAn37dPz9ssg5/G+3sF+a6kib+rWon0sSkgj+
TBcV9JgdHTK/na0POg881HubmeJH04hgjZFAT75f2i9LTU9CXq/cvoqBBSjzRB4a
iELtYVTlxKB5SYi14HCXIZfqyjCtlriAxI5nNSYpAioDgINMk0kKRgRJSFWq5pFz
cyIlmpZsnEJX4wP/PTQHjZh2goQuly3sqpR1/7G6XWq24/0xyD6wUND6iU6+KSIj
bCY2Og5JYCEwzMdkUZzDvRRpc+gdUjvkT2mwlw2tiz6iLtX2WeX3JkjyFmzKoFEO
8C9o/wIKRw3DIq8TwkUb9DS+2pNlslapzFOG+NhNacPTid6Vw6HQ/CQRD1S+hztM
n7nzvveqfVCYt7ZeZGJUvXpCd5ordbxhOjPr1Bn2QgPYa0OivycXDenyTrYjABjd
A6IVNmAfxEwQBKpd1CycLkchv7zzw5dIf25Eu1vxV/tg+76ck/KIQv7H7Jk4Zd1t
DKOjdOYAf+ESqK8l9kZ2iMuK+Tlx38HXbO4cilZpWV8jLoZq8AyEd8JL9B7abtAY
a3kvkekrOw8Y7NVymIAzH7+qxJ//5gKvXf1ZfuSI9Z+6KduhATM3vq7CdeT34v+s
a4TXJk0vrD57k8LXIPB9ouwXEm2UOUUuzqz2TxhTNAU/asuMXP4NE2aX2R9F1DSq
zMez7leNq3aqGd/kUB0JdRvx4knpnTUAxxTiY20Bk9EO3DbFjLpUH66fNiIxQb6q
5+YAW9p9NlRfThJWZoemUyD7I9h7WHO3YDqbMXzpFj8iCnZRcVrDi0dMkFGZFXdZ
7oslYWT0PesSpI4ZlTqcOE1AW0vLHGUiJwErFLN+pcnw0K9i/u2/FtvjpHkXk4u1
wyHw083uwkcXDy30pK50aILxF3k4RLwmy/4XR+AL3fS7WQEKNWKDlxBfVBvaoF9e
kRzS5rqEsg1OrHdoewJuj5/viHkxuHfVjjIxu3GeWbzpbUZv9fO9WuPqoRNYjYMB
aNeClUdnYndsg+4nGB2SJ6F4dA+0Wu/Gsf54aqZ642+1+HdFazZXInqXDh1LfwOv
QqXTu3s5Lo0R7yWPPoNBkhjyVroLfuhXJQWOIO6GP4E1xcWYhUbt4oeQsZVYWFiq
MrdXzjS+ka1pu7nvKDmyzMA8ypNrxz6TnbVT/7BD6mIrGOXKgN35U8ecE6AgXP+h
Mk/9O+JAxRBRsXz39mJ8SgKnrTPf2gXGf4Q554P6RidGIICXvI/s8IDKHLkIYgfY
OQjJMyZ5n4jHn4FGZX1V3Fn38m1nvSOaMrcN3iH0VVxeW+GpHd9Rt0e66ti8a8DZ
TxLexiPchVKr2qhnPm/YlfRxZQcTOYHFBfehbrDAP0rg1T/tFPnxlFBdgNerXIj1
ucFENUT2ReHgUYedtk2D2vgf2xYCNK5rHyVyuPRKGqDdJtjL0HvgeDDYvyuielY+
ZdN6PF2bK6pS5hmheC14epNmJNvp4xZ/o3HJ/iH3xvlnElmBw4winEU46kHD0jH+
FYJaeP5FOMC0EYHlbWK8I/XM/7GnqCeLSUhpqsiRh5CKrR5KsPIKDQGjcbLlcdhY
4cX1YGDYOq1GAbJHsWjTKds2vLttdFo7IOO3As7CmHbF/JcnMQJ0gNTlAUQcOcEx
mWsOQC8J3cBFUZTTHz2WxabFSHCj6X+x1BvjcBd8id1JsWSsFdK+SHB3NPAmAyzS
AbAwYLdGOzAj1Gny+PRsxK1ZWHl1bB9ngCD51a0omqnDEcZa+XUF/GGjz9KYlx1s
KWKudtveUJqOb4KJTcy5ClGKB+AhNlF0DD3m4Ai07+ujYgANDtpWq9hnSaddYpgn
qZbiCzaV36ETEX7OcE23zt2Ku60ihP70UHcEluvtQgxw9wO8Q0PFib2HfICz+qxv
EDWhoKdyrhZl7iKoT2OtMKhtTim+bpTd28TBHeVj9tFWCH3OliZuFNWc7qmubniu
JOQnfp11A3pUwwV1g76+9bHoIsPs4idBnn22UieUlCwSAbwifkfqBfYjopWNo04W
+Ma63ZslzRxPvjxEdDjJUgv6yIUEa4yyMSrAiqQQMweTRlx6lZ48hWCNZj/erIU/
Vzc3d9eghrTv3pTdJgfIcDRsOtoO1GfvCB8vkS45SIeNtDoDLp7fY0CA0Q1bC1da
L6BjvhdBbp42KmteIqtt4D0vlVNtWcT6SFTQB/mdPrKqyYtJYhgobwB679RVmM29
hTFa09rGYIh9SAYdIGjK4lzJTd1VDaE8IxEPrJoKIw2fUMb4nRmt3JXo6Tv80JsT
Bbaj3YmtkVDVo3kWy16558iRnJZ2dpbnLS5rND0F3hf5u3Ej7LXrabPwDQZ0XDM7
XeosvjzNEr/js4FGdzgqrvezgTZ/RAE0VGFEolWCLPadsxqUink3v2wUAE9ReMTa
JEw4wP2Qm4bj7tRdky0w/75w8hcD2NELULYsid5HnjQTbewmmRxe5KUczA67Q0hM
QG2npxyX0+2AlUiPAwav88Jt046zux4yoGVg7rcoY6D4aw0yNlb9J5BgHVxce410
znuVeEWqjgi5Pf9yIWhklH+A66M7Yr8NJjDcr0Sm+YvWKw2cb8svZ/1RIfmkAzcp
lDxTWMQi7kQhTZAMswncZUSQ34xuDmgRBV684eJTy9BoMY+Q6aBpcBczIiOoTSJQ
eOI6NbRGL7HXWTke68p1fxt8uXNYeg3VaToaBp8AaSirO2a17XBOgjGooScMdmA7
9evqMAWsxZb8hEG49MeddoJ+QhPRnZCD/LtXBmZp6G6OnTmsG1ste5Skm5zzMFMg
oOMKh3qtbyFikw/V7UmpfTB6uAFDu5IRvaqemPgTzbLu+lREpO42Nx5uVVW7IPfo
GpLUMN4AH9wNrZlxxvWeSjmroFL2v3irQPY3vwfd36TaVJSCKhR28fCD17Ie47L7
BDzvyRkMFxiRKPqpTi0z8okhd/xgpLBpMZHE5RpIO4xWUXZig0fKT6K0FqvJ0evR
sltJZm/lLE/wyM2wMmdsEbEG/9JTxjaFfiCG9IC+4OszMxYC4QcYq9N7mJqTWaZL
sL13F3ewLlCsr2Ej3HvrYMKRwZOFqSRWuOoO+qXG/jOKXwMDyU5/omOCE4nXRl+V
gwlPpzQHAU57zj16d6yD0oCNTXColLQOApC3QQIG9Y+aWrb7aVJv6qQexBZUqCQe
yhIx8xpOCiZgwXQ7pSOuY0J2JVaKclwgfCOKRMzqIlIRMY/Ck3it7VkKwKEcqW19
3b7F6cbAEzJT3MlkWSJ7Ln/0GhFgrpLyDpDDQ4vDmwTSsSjlME4Osfmj3fJ9yAzZ
FQkDHFhuEHPHsg3wgYTWWi6f9Zy1Z7BF73C6EIjdF/LHbGxcGMPAT6v3t07dXjJM
pxN8ESGpo8JKirYWdMk2TG2p2vFUaBcyDG7BMyopK8aKKTc7sGyQWHg0PFh5s94b
lMZl7R0zFOSt8mRGNQlXLK6gVM/ek+tIdL3cnnEYTupZCkz97aUY5VIgUxiXonfV
AMw7EB6t0hubW4cT5O15hgme43+48Dg3qD0aCey7IDXEjQRrkcg3NBIN1AJjChz/
q0c6EekqPSCgkl8ihMLmE15auouL+6ffbggvtOHQ0JxzU/o7x1t3Kp3WUfcf0h+n
SYxF+2UhZf0G/UfORofLvXJQbw0upciK+Lk0SkzRN7c3cntkaBn/n1hs6q6EoM5f
UQ7Obn6hXP/iAQA4VbzbS6Ny6vbY/FLvv+tOuIkSPzQHlkfgYTup7QqXQZP3S1FS
+FI9+VXpuPLl5hQauDhO1xbwJXGozo2gNN1azKPdNyxsR54ubuRwhOeRqW5bY43L
1Ptzj7LWEIFMv+SlaVs7H1SFK1B1uhENaHxiFN+mvA1DIPj495vTVavEdoB3ahTO
uiaUKtoFFKRK7P/gwFrBfAc0myZMhEkDkhfuDONmpPLXs13uWMpxOVgEzzI9tgji
i7EHyfCSifYpNUKidh2H5s7dscOnRCgPpD/sLmfSPL0ZZBbDlJBp46TCQXj2if9f
mxKsrJdniiuMqmylkikySxfCT7TSDtxNxZDwHqVCdes2IfjO+4esmtV/7X/fGvLD
3ElaTrpdAiVV0LLNvT8gd5g5MLQRH8xKW5EU/klFPt9e4VCQqS7ihIBO0AcSWN2y
DdfffJEBGVN4ujvzKAxp8iht4kbTB7RauaMGjhBSrvn0IvQT+ip+OXfblfoLwCyu
qXXJM12iGIAiMT2E6yholP0MgNRw2n/918TdhMLN15RqW7pE0rJgich5bTEaAOjw
f3lLRq3iDaRl8lO+3vYrycfyku+UPFBWtcvkzGBCfwcttDxN/dT6MtmpTKPhLT0X
38wo/Fj2T8CsSVYQn4GQOOpkoIK9fx66pjgfgHl6NDuM8vEV9j9fCdUN51VO5Kv0
l/yDZOczRiHL4TLkNBt39cnazyYz9DnzDo3vLDSvC8v7wU5v22QRt1BeepdxUCUO
DGS0AfBH3PHOMODbC4j+MYo19yNR2zoStGUt9VxVEn5dzDuXWtzmf/KvogEYmSKP
RwYzSyQIUDUBfSFutzCZ1knfk8joQgzez05jXqU4JP+vUbDqrYCNlQj2nm5rx2XO
FiiRkv+vjqD/4KV9VTnEOrz+hp+7C/nWV0E0MXHfDPLbi5fdshp0gslrxAoCnsPc
vZ3YwEiZXToeyPwqUIfGWW4w9f1DB+tNmPBJToGp3mw6OmI3hzyKdYX4TLtbyZCM
9ZjpH/CVID5TmBTkN2sYow/GWH0vgUvUcp0K46Fbr+o1TsfUTew2tEHeHQ3RYj/N
QrZ6YjRDzNIWYmeGKf/K5AmMQWBKOs6+MuF9E93y9/OyBtSLitNIcWUSxHTVn1J2
OeTNdlH5SBKKHVAr13WEV+CuY0NyGp+ZfVIc1SkCzAEzP+YrkJ4Kb7bHxCKh8lO7
gvBriJ22XLbW7UTaJnmqHqXy90zI5wH+BD2q9tqgLtZ9A1D3sPavy4dnDjUi6P1R
SPoC21H4oPcwAxDDTW+74Qq7/aRGgYmNCeOMQ3n74rzyOe8MaHLHNr4rE+3FrtzM
SkvNnEYWA9JuLGn1n+Fvk66Dy7M84pB/Dp38V0F+nsqz37yk0k15LNaoCB/r7OkP
d//VmbfxTJt6L7Z6wUYHV43qD/T6PqfgQrmDPxOlqTxslk5CVA/6mnECP1yZRFJn
fIobbuI0/Fl9x0fq8ux0gBD9QJQXdEc/UquNm6JDiUIuI8HAqsne5cPzA18M2Cbr
TP8Rd3XJRVMh7b1Zzvg609OHNpcW2jkBjzX8T7Mhd1aYsTdpOA3zFFbPeh5alAuy
TsPcfrZXfVqF1pid19+GkVtWByUw4S3zAQG9RqS4Wpyay/MxnEcjbLz7i9wuSVW1
tVJ7AOrRiotel/oKy4TBGn92SNmJvoFaONxKOlvj0IgrZf2UcVXgrXyr4ef5U5BS
Dcsjer/uA42qQ11auHCsZ/DNF0bq410W8umrJz60vk6H4cN5v351CXy0CXLVDU2h
WUIc8zyOI/Q2ZixAXoUW85xhReoh6QBfD+2Zv/pfYEt3kfmYDbvoNzXDrfOe7tze
MKDxiWkuJB8b0ceT/sdXCIC2/HunA5nqGkO4Ccq3u4n0GMSJeEybAuFpdPMNt3VZ
Bd02o8WIqOw0sShhSAYVDFfMQ1n+lFObmbGiTLgc8BsC5XiEIf3IkPSzx8eLEFvP
yyXsVLRNiRKbeJ8bV5jZUChxNP++ANM1EEbQ/fau7t0SXOO7yQUHaQO9toT+p2cd
4EIdXsBxlF+uk7u6fmYe4uS7Dlc5qXnBv6SQlHz+uLFpNr4t0yD/EBU45JZutuJy
MKcfdOe63FcjDFh+uQrj5w1ZCwqBy12uPouGmdgY7/AnpKrngMWUgYTR1Mvf9G3Y
kSLIs/+tkDQ6drlP9v+wn9Wg4sx+AopXCQhe+/bFkDZuE33b6l7Vpgzl7ov6ilU+
cbLGut7KkWnDnr4XeQ0j2O4NsfEY8TBhp0E4xy857EX5vIEMWkSQk9WwsckEJdW9
oxsin3voz86CVw1sqUKECnfU2/FwBqYnk3RS1jFYAyk68ahE4par8ZX8UtGZVudP
8sOtvhhHPeiJJ+9Cfnd3sTlavrV8ZE7J2+fJfDuC4pyPBeL6AiSjfuqTy7KZTtRm
vC8+5L5dbx21jk+/jgaCWewjIqhs+cppwFGpcIl6rrRXtzQWGmzatpdHPwMkLabY
F20e5LewJrygPMN5DEYrTLrgu/MUSa6a9wSGVmEXlUpJsmIfmdP0ZtF+yjCu2GMS
RGZnnUsTHNZtW8Kp9OLJ0QhsFhSvQx8yCN2s05S1TMszjABjoB7cd+wsuIw7IHjb
+dYHC8J+ByJNE6mvo2PNfsNrClllyk0+QzWimCnKx0c7llv2kWnQNQwgrfii/TNp
DSVLOugk1Y8H1Bdoh1+rpC0bJ1Hj83ssOSgrqu9KT7O0gSIwoOL2g5e+lsCXP8S1
mKDmYghJoo4UkLbEq5+FE1c8dZPkrSxm3ggBLkgJzlqpa3Z+Pt9gIezPscZaypqf
VCbplD3QocKTEq34Uau7SR/wM922PY9lx7rdrYdzWRc5p1gxk/f4aCU1Tq5OQygy
oTt0Hbyc8fbKKrv98B1YmzxcN5G4UHtqGV5p24xgilVKXJNDrQpD0hnpehVb6bhG
q2359YXjTmWpzW+1RASrOenIBlKyrblcBqgH9IiC04l4fgDJfYeREwWg9CvSxRls
B5/ssLKLUljNJGRcr3+H354TZRzRBqK7k2fIhmWe5+qS+aQYijWlFlHmmVmNvVWj
IBPt6hs+m6xHYGMgbuEC9kZ0BOkjzk81y6V9cgJleY/ry4hOv3Lt44GH7ywQ2YE/
Vfba7NpPtFu2S0dh6a7kwmVIiDUDXHS9LK8WP26mhS8FkvI9Pz7/Fem78nWdEyuK
Ni80VrzsGpKr79zrmW8XrygwA913ZaT3A3mlTTaBEgbOEcsXNEqqwgdp/2itNnYN
tBKsUXCExMUtN9ldJlnP0tJwo80MnFhMWIdXHpgYQd6DmGw9lsKSOoV9H5rY+opQ
JM1Pu6xq9e2Biws/qFYy2IMwo09DmLoyqYuHQ3DzdoiLi/lifIFliL58clGyK8js
9a1LnjArB87HZ+IxSU00Gwrr0bs0W1DnN+9Si5Kpz3jD9hir/l2M6b8UTBzN+2wL
Fbh56zuMd+CnaRI0vtYC3E0MRiIFvxH4OwBUB9h9SeMips6q9ffQZrKIXUExLIeq
rfpNbZXQnW2i7WWOFIO2VwgE1cGawUejx+uhPMP1mfCrZdaoPJsLwNN+lq5EIYoW
Jf+P7gwgCYeMXTyBZYtmn02lc6FSp/drQF3DXY5mIhbu5s5anIkxqeAoh6Wl2bSG
7G//UOzz9MTttCJ/BNYzWcLX9UjSUjFJ46gfvol3HnMyc2hzrirnjpMH8190uSkO
8jtffRIXAjjVt/FyuiKtCKugpv0u2RgKqkn4SxsfjFowRNXycVlcBhOvAry9NUvq
TTgSkBtX6A0OxRL396mzCKMqYu6NQLOXbM9TFCSflkSOejxs8S+kFbLIRJSY47jT
dHLsOArhUF2Yes0gOXcoRQafh4TQghoyow2OLayZLQEpOt9T5Qx5uCFJMO2Ai1hg
/cwSCI1aXp5024IA8NU9+VDKT5nseZnlIO5BrLoqrvKLN43zPfuQBhAlrUJUMFBK
uvOruQPeDathBAZl0O9sRAL6L3M0dt/JGpAmpmEwViw08v6Jy6A3Qdx5n/kCDX2P
r5qAaYeE+838I64PzoxIOQVqhwGwGLZMQsUCdVO8pqij7lvSBGbqlZuXLbeI3QUx
xoUaTvbgPx+v/iB6SwVsRYJmmeirvZjjgAc/KLxGwBMPlZJtEtek0F7pURmg0dZn
BBMh5c/EiEh1tNwTlYd7nsw/ASUYN1qztTaN6vM5+AETOUAP1P+E6hieBgOmPPSb
lpfs5jEGc1fyBlmxAmXWKp4+ET5NryyUnSUnUEUD0NqnuBcfsBib0iUkHTH5J2O3
cxt7fmVN7XJqby6TfJcqtgt9nloaje+Piai/uK2Sq5vG0I/CjjjU5Newt1Wrt/Tq
OTjyOKpi+VCfSQwWeISrmvf6f8pXxLftaiT8moEK/e/S5W1kDm2qeFqwhl9XHU1Y
+DgpG0zor7baaabYgifCtRriTyXmVztT9LVtCgI8ChT8arqNewEiAAJjzQzszuIX
BwnLF1UbCI/GWt9pmk0P+a7NLOLyCf/PIWv+Cpsy/B+0n7fSSHhmt9uITHijDOH/
GIagxVkd4Zj28o7hShZuvPYsLVybZ7quE9gMg9V0dgFS+SxRuisAr4hdQom4eLYj
d7kYh5WpowZZKAdLBq9fQ/nX83H49bE8fXHu0HQ4QRZRVe6FyEnZlixDTzrw7Wxd
2Ce6Zgdk2pSK0W9wwXTzwOXb3zCJlILF19ZpsLK1hRj5oiWbIO3b6eXA3AC1IyT0
pxotqQIyLjK43HH1IT3gHtMJ45XIdThYAD6F3/0APVUPxzWh8P9Eyf0o6jy1lnAL
8viuMhMSV9jOBA28QrfUCqC4rmpYl7S3ALrgeWRoxnvsd6DCvBhaS5UlcwvesE7g
APmB/x6SFoXubPQw7KyR64oXbsq5W0TTHlteIO+xpyxbhUjNOUGuDGQPLRfVUx/s
+l6BF4BKdUk2yKCB3DdVDvd/3JTJolChk8by9+piIUnQvUwRfzWKTpOKuhA4cW03
6oXnJb7qRp2Ls1mLIC/GOhsyY85HLujsAKqe+ZCIi8Fs/IAk6QOnz7hFvKjrfCfr
PoLcW1KHbNF2lxIVWapsNphJE6Db9wMw3JkHCPxcr7S2k6UNf23QGcswSxh3dIs1
CxC28U7bMbOIKB5oG7rVN9aNIBaVyV2XvWvzcxaCRkAYrkU/oJK5/BaF6Pjpwytw
VAWajbx29FiVIjJV1sr0gUHUalUduCa44RygsNUmld4JeKypsBDgMr3wkEvzdO/O
U4Bs0hVam57iMvUBJMPUxMHRGWuFKvewWVvpdFx2gzEewUveWYUZY96/W3Dm9XDy
ekigXr+7mJBeox7YHqDH0xb27cX5mW7TXC+ylG4wpmNxkxG81DHpDLOWw3gn+RD/
jweyyyza/vJUlzL2/u7r9gPFX2aGORXFHFu5YaIsFQ/UbWgVrrkF6Ckvb3FFwbSN
ZN14cOPPHEPqztrs7rlfSMLiBkLjQWsNCfP0yzZqc6FGL+gVeI5U45peUb76h+HH
YHGGYakbLqLXkcOZPIYi8gT+aORWwRJUGahuhzaZBFCkqv4I5eWe7eCjmt9P1FmD
+ame0MxOpdWKismM9EQURhvs4tnLKkHzmbIG1jcuUTmFX0innoSH82hn/u2VAToi
d6eLkKcNxhNGeYnMqnkqOU52zDZY8esGblq1t3msl0av5lc0zLxE+xMW5cKJBsc5
BzrTPBIkqddisq/bcvly/MQ/fQJxmWCw7epkjZEeTx0OvHYYsDr3HR4VzHEBBSI/
ediwNlx8p51w/Oz3SqIPDcCunpoy4I1SMxvELj9WsAlxLPrujnC/xWbSQaPxb5jh
mPtlGJcQJK83JAeJSbikkTiCbSs3RLSfFhl1iLnp8JjYF0+1EqwRaW1f6mavTdFP
KOoaqSUw8OASuBBYjDbBicDI2pZUKaYc68one/NxlSxl6Vx6PPEqfY0wMjgumh9g
Vk5D+pA4OEzkp/Fcpr3AZo3/EUXoymK95SmkSHlZw+kL/ZaHF4slL1og5XdThAvn
h/SN797bQQmkJE3pGRZaAfPxEecQstUo6VsNqiyQU9LnVMPo8sd0a0mEOYml9oah
EoGh2OSI+MLJNzIymjavYLyhB/T41aW0Xc+QowsY/AX9iw/DVKKZZKMkUYIIH+pB
r5UO6t2WhOs3cd7cmp8VfnDd76lhpzStgALDaJwTRqacsPLbD6AL1UJpRDO8oEqz
XIjLMnlS9LkGNhsf0B+3TCF10ppZge4OARxWRHdtoCdVTUgk8MfVmfYFXbdnY5OT
9pHa4+zTexf71bNYu3AemlrkGzIqbANYq3m0jwcF/IvKbUADaXsYjAlAGPFKmiA3
6A1ue0/O+G732i8sv7Ci3ECiBqTU66HS2K0aysxmKixk0ODEGhW25cd6aT1PqiQG
OF60L2/LsyRsC5nqknavgTfh/fO8tZ4iov8OAmMJ0a7Q9b4/eadoIZlJXyVhQxwe
QQQxmNtx3cAXUnzKg5XdjBxYHSoumSDdflaIJ29GXEDTeN4uUJLtFYHb+nEJYwo/
gB6Adu4Tgn4DrKPbh5wvPRA29b5KDbcCy1PsQCVXm0Koddci7nuNJGM0SB6XaJAK
o0e0DlYZ7ePMzTkOoa9diKzCOMX00L/7ecEYGC2uKdTjSRi9CHrSKlCuLFFGtFxt
QtqQESrQW5Q505Bfp8QIkcbFPwpIuO+Q5hJiwYxJEZ46Oyn1jR0KZbn+crsin/hz
1nTMjbmak3SwU7gPp8WLcczxiGHBmbuzrl0Ui1VBS7yWMnKjahk1q1aTkeIBn80c
FGGngGZJzPnSu/J3v8KN/Qtf4uA7bAjWZRZolTwmhTFjqs6lr+VqpQh+OHkccWyz
/6sObi+xerE5gSWmhrPWfsFZ5OhuYAW5+3Dz39bxyik9SEom8Q7NOksyHudxQmyR
C/ekdLDtQ2Z+bYEg0vDVNjBQjlKXEmnF/s7WT0RMKzs1XIZcF8G8KGmVaI2uqhBg
oJl4O+D6IQ6g+T1Lu4wkRBZ2+1IC+LbhLWmVM7ufCo/W/9Hjau0kQSUiMwta3BVs
hIOA0n2/KBgDwymUmaihcfhfVUxjKrCXhYOCYcy5LqjDxubwMz8qqJBF2Ic94P7I
q++HGKL2FcDxbsIRqlx4f7abTEHeHWlmw4FOi9uY4B/bmy5uaDFGjRHMGLubnts/
IwGmHmRHYIY2wJW3DdfWhrRAHWVleATHe6ZlFgUUR23bhqIjzQGKHuCYfdgPoyJT
lhouS0vROjuuUh7fdsBlk0lGTreptZ2a4Xxz5gL6XsJ1EuOMZpKHaivwNo1BNghm
cGdumbSgCrR0w3VPZy/0kCCZwkiOHv25mBIG3OwSZiyQX7DIUzAC0O0gMv3DEq50
YBCdwHDSkMwM4yTiickawGb7eOQ33bg+9JQKpznSUd7TaXEJo2K0DuGxyLqtaSKs
oDp6iFowAV1vdzKaK65QvhFLdzcPOJ9acnMnVxsXKS+dHbN3Q9fgGgEiPP0AAyHA
UKhzuvFv74tSbk+6j1REXoRxAXH81Ryp98jBtjbCUFsywUl7Rb3vX8Kbg18CcEOC
Lx3YRs8hcqhcEm5zCIKkWiWspQKhXeNL84fxUgwBUGL+1eO5qXJ9s9ra4YCOVyyQ
+8BJeIRHuNmP8x1pw1pxHyzbGtJxj4mjw0eMiyBDXHVEICZWp9DrZMk1w6l/4ZKl
fQfBD3xR0edLl/b8hbZGabuNJSkBDwkFI2ARWUWtwYm6ToH/GbRceCmoFYmeGirl
Kj+/DqvLl9HwhUhwaQMLo5MBs1T/JC05U0moi+au7Ecoxy0AmX6wEnqdrkeYwHiy
bOPaYVqpZ/YglXcRJrcRHsqWiFwloJpUQcnvrsz8rsVv0sZ0TI0mB8fAyuJELAyq
00EH0Ss3H0K8fbhQ6xtzRuyh0NgzTpsecGtRVA7z61OxKhXYa0IK36LrsynyZdG6
bdQhueitpkpXdi0gkyv7XNUJkbjVi2VoU2RcaP1J/NLLtXAoIlgmVQfDPuLfBpBc
QNi4kxvHRansZqUFK6zkVUopWyOzryqz8mEAj/BWzCFY3FMUzZvufUyJuPvZ2lht
SW2v7ufQ/p1dtXftiqWatbFgJjVjLXiG54vUDDLOvc3jd5DwNlnTsR+gbvViv2L+
uq9CWFMZoL7LGTxxF37iQP72ACNgsnGUZIrvQeJ0g6DPbzVS+03/JQEdr4TUR9q6
WeEyvpX4N/Dmp7+HWD1m7j3VMb8X4zIAdrENRipw6PT8g/4Qu4RcbqBKkCLefhyo
ePcX6Dw7FOkeoXQZ58dbch6VOGiE1B1ZhpB0Br0yzuPFxFHvnKb0Hk2J4lNGkkXu
PSjvJrycuo75Fobc9xSu1UDwXNq26jUbqrdmTvB89pdMiPNvqqqOzw5VV8xTsf1T
MVWzso0hQ+RVDIAvpl9MBBuo0s6a6xIHuCYOSP5lbweGcajt2qcb3w679FIgejkF
uVCSTzdwUeQG96wRc82zo9F8QHOim/FkZyEFhFxVIrlEUNpgi0Xx0SEHyNDN+Zb/
rN4QGTlc7NX9jlUISNVd6qBJR5edK8GwJkq539w3/BrucXg+MKDVWcqbDf1dGxKu
Rw+m0dLp2a77zA4JV3JhZJg7rBPay5hW3KCIBcuOlMBy4QblBUsKStZPQXvPguaC
YEyxIJF28yoiRrnH3LnUemyqaI57c2EzfYBL83MPFoARoKA9xoDkDuL3i9I0zgRr
BMLUYBiMrler4V5j0nT2tF/jSXFf0Ys/NgGXjIWdU59A2HlH2gwDPY+5/NbLwKHy
O8wuH9AqdXNWrGX+bEEyOstuOmNZGlCk6osPis6PgH7SeL/R0Ci7noeDweQb708W
1bPPBebaU90eX3Pt+PPBbpszWSfp1fnP79mkup80flIT0U7oBxoiH+5JdOwPCCM+
8GUBNwmFAxH51zCOB+rbIRHk+R7jXpfx4pvJ7iphXylC5abG5cspiDbqGTrstrTp
8h0a3UKO0FMy7LE5QV6kecp4w2eVIlf4KqPyt21e6ADcfduEFf+vnY37L39VvtXU
5YWkqmyDWL1RRlSIkdf9K6GplKl7+ZvEQReuPVFIoZ7M4t7lrDXUZv7wo8VVASNy
vjMlrNvqSnPwWrcrXVXUTjSITaSt3DB8MzjNcaHUsJywJS3ZS8Fbv+ja5JGmhEy4
JL6d9azpHAqvRi/XGCpzgMDsuehn3zZenELYaTlkmbfrORBkknHTzjEDnPdKPnXL
6BRPDpnuDUXszqWwI3/6XMNPMOASc9HGrzeDLqT2mwvjljSu6lKC82pUQC0reIHJ
p7yCp4o4xy15jRjHyblh5tgDmKkNRmAqDHHTyZgNO6ElD2Yi/mhTfW/Zvh1aFdrP
bHfe8nB+RHvtGe+A0rlsrLfBEEc955jK4Sr8Nh2SyWtEcww7EpVIcjdfXGevwd6/
8zXVNHXK+LAilGfjGO8Q/FzA1jC5XJa4uq4CkxjSWzLQdqTMOEGTaCzbSFQOaGzL
VlqT+uTw33U3JzyO6+GIzwP6w7x70JuZ8W2NJijruM66VaBp5QtXrDX+4I67YBDN
MRMDm2JoipxBCIjNUMgiE/XvM2ZAXcPCHpM+NuR6bGR/93dlUmXUzh6qDiVmJrCV
8hOF/G9lEP0PO81LCHuK6By3iwSwyKVgk057weMVWerrh9WSv4znUFrp6KagZwtG
x+HwHivB7ser8A0OESdp23JlEmantErhHYb8B88YVWSSwfxAj3ofxfcJbynLlVwx
2X6pouYW40ZXa6uleip3ySrJUVfS+yca7ArLex+cId3YGa7OQJ95l502nI4spr59
YF6vqWsJMaWoJ3jDOuTBJQtIMzJxj5Tv7s3RZLyRpWr5HVA1NZ3JkyEvKkbqVDcs
V5/McQHZP2vcugRPBditVGg/OC+YgHIiaoCBuakIa+9s2P2csaHBZBRWjsYwH+5f
1BXSqVB/fJqvObjtxbrVk7GBWBaxU5jMKjtBJpn4Hx2WpKv2SeEgznay0Vw3ELhk
+SEPsGlY+IppyUfSJQemY1sNhH0TTalrrpGAL/gKZFU4Bb0iH0eSBZjljKODCil+
eSt+8Ul8BIHl07PdULVWx9Lfc5snHsX/D6ZFkpKZAsu1Mu0H5q3UxvoESOME5EBF
beu7RpQZ0+OtfWyQLvzy8EnN1205ZkX5Z4X4Qbz6Mz+zt+m11tetcv25Jag/d7oA
gNLCSg1wqIONyXf/BKtwllyrd4fsm2vF7LaW33fRZ4h+U63TalzIh9WhXyuiQeLK
znNrTQl39L6qkR3lzL0JX5xVulupmyFE0LHgB0zDrluCRIRZt31joepAs+BTLqGr
H5La4mbID4xGuGcqJ3QbFZEXrbvYDPvOOa3rnWO9ZPtCT//vwBvaYBVcajZQSspr
Le++ND3T8c8ICxYIhoHo5Oo0dWIlJS1ycjqgpOZ4XTGkxM5a3X5tfuh23TC7mrFf
/7zBiMYYuD/LZwZtUF2Nh9+7ezTLmqsvLRO45amkWPwyc7emkJC3XFQ8wah+wZ8S
oBvjpjun6WOX61x51t7PVFxWRnwHeLXP1vXTer07lcXlErJInKU9jhvNXfiE0xoX
5MnzpF/bJQMTccY4S3Z7jsHpwdmud/ig5I94lzBTz0klNCb+3BuJP+l/WNvI7reS
wwJPxhcTWzv2OrAwdfeUP/WHqxa7I80XVfNM5yytstCH0E7qZ+n0RWldEDK+7aIa
zPXmYmHTzQ5m8wY22H9ZwAyAgLr1aA3Q62uyMq+T3qUqaq2rkFZOtjJEJwjuxy5m
UM18hTUWSoIaKwpQYj874ZaLYfuYIjTM3Zdjv2qwl75EWRtribAOvFQhyelTOHlz
TOCLO7KKukDZcD4mmlXta2CBV2+eDWq1d8i6RtaXjTDtt9Z7Oyvoe89xjdsHUryW
ne93k1cZ3ywnrR6Hm6Q56N2buF5s6sFKR8LQq3XfVRLtak8MeYEkbXgHhy7Cq00X
wk7fKl1M8627BW163Ra8Fj+zWFBgHX7dkloQyUhKXPIMg8hgYdC7qED+JTokK10o
zTbr77mzX4gzQVGBYcWJdy540tz6Uqtd45k3UZDRRksPSjGNE1YIENz4W1fvZODR
NbV/EgbDhJ974sFkZqpr3OdVskzp3Ks1RXywqyTdG+KlqT+3ifAlvtvIhmfIrlmA
tdlLqyZfQE4dg9nYxtZxt8uWvSHSECUDy0GnKZySXGsdyGWZkY+0maJZNwnQKgOq
45Q4rWBcNgYNE7p4qajYoI4gc2Y75xLc0whsclpgav2Ry0qbQlmjpTmE/ohKqRWU
17Tw8/QZeiDXEpcRR2EPiEmrpIRvvtJTMuDzmhuQROkQu5OWem/miXN1hdpPwAfG
+agLqsZ3BiVTSRM+6Je04Q9XAqfN524PbgNGakhom1/z7L7W0EXs0ox26WJI5yoB
/l9uf/AD8Qaa8/VxYXauI4L2+Ia91/+eCUHWPG2xooUPV+HeZiOklQulzsdjKhG9
fML0c3xnQYuf/s/8sxxgfEc5jZeCcgg1uEtU4uA+mKIkrKiswws0Y2NK8m5BjGrB
pnGIXKUdKX5fJt4zAf9L6PQ1W1s/9o2c9w5TAH0fQ54nBU02tM8ZOULbGWKRIYWG
fwdyxn+UyjQ+Iv1nCNLqX0ri3by5rXxve//4GzRzHcnkbbkP/4yOtI0eeUsG9wBn
mhenmZOvUpK02huDVdL8dhBLgRJaRkzWVujZgFnTdEoYUvhI4Y/A5BxURAJrSZKg
u7Rpaue+9sljvmFm9BiQzw0mj04Ery1Uq+aIUU3YeTkknzdRw/EZLAqfb1boj7D0
avMQ0q+2Nl4OtoF6uTKN5cCRgnnHp3Dh7uHmhhWYSu4yrRxCJab2132tSW1VecQj
N/OFRy36pFMpUZ9Mn9z6DnI+2DCKLp6lM5W9PqIkqUYEgOxlIiQPTf46aS0L6EeU
Tm8cTQXZWLa+80q62v5Ndg1azQLhT6TAAfnYs9KTTZBRFEqQLAJuM1byA3w+4eJK
8SkfKpdEe9QsV5ttD2vykewvf04tVvVztzotSIqafarpTB5N4iJayFG3E4tEkmCN
qzh81RocKcHmVO3UkiZFQEsZKW0S0u1aLOWvemCKHv1P2Rdo9AQXZ5mR9l0L0EPS
fvXV4qjLLpEQ/pfZKfKwVIseUWDNMCAAnhUjKiVydMMNg0HwOgXteetgsyU/e+Zz
3NJ0mHfEFaoCuryTg5QutC97ISqjtWPX3GqCa3uHVeXAtBBtk1vu0z1Ezn8W7wpI
ThN0I8gsA0HwXbLULVM79ZlSIvval2XzjMZVoFjbJG1P7KK/q84Gu8IPoxeOQb0M
e0mg/RkngvcSP8CI/UucMkkS6w0PzfOGUpWfDTodrhc0HUqz/TKla2cgXyzNu9zH
GaYWB6JPh8beYWEfWYSFSH5HZVzroOokWxQrOvJKp3sQy1qakipdHDLtxemF47f2
UMkuI43RBn/FYBRrxCMVeq1Mt4gVJU/3wF/orjy79GPEMQ30cFtcgxso6r2dJqA+
xjQyEiNAzH134n+eSSI6rl8afySOFe7+rLyFWGaWsZxmgu+QzaxlteTmTqSp0jxM
19RPjmuFpD+Q6Fb9Dy2Y+1L6Iz28woMNXuBOPksSGTYGm96PlNoIUpaEMouB54CU
BADT72n+eaVsfcL72WWEt2t5ME2ELG8neUgiRP/VggZ9pR2QJcmpWylTXJJFVrXL
pH4wAqpLittsCPpXHDxirHBdJtDR4IdfD+2Hukqwc143U6P1ptLNgFrOasdPmW9Q
IlPM60qKOO3E3gNkr78g+tNrRC3jwwr5vHgZDycAGGP+GZJvtbXp/eUPHAfd6aue
BpocWTfcXl3fqgxowMvrodYz6raepnnbrDxkFA+5R4VlwJoeTTHT4Tys1dEtJW/P
2poBl7Ntz2ooZ07JI7d+ptnnh2k/J4ihrIcWu8mm+sAsanSLu/zt1XSHxbF000Gc
pf8L/gIicZia3bvs4l6wsqmIe0eMCP84MOznIZlT3kAe3LWsd2ulphPOmLOsJnkF
PXzOVdSVU+2Z7IO4VF0qeTMQvFzs6oI6O5s95Ju8FiWZjgibe+uPQYWSRvcjqFjf
nF/bKHw2fXVp2q+HWZBkCqhJAUI91/F896llY861HeDPBb7kqdr8fVUPdQcFXtGJ
09/7QHPVbyKUr68v/k5ZpRRj/VWQVsMet7FDfKur/lc+q3J4GKJ1RIBZhPRy9R91
9FNbdYzvFZYRgIjxatGAgIHWvfLnWylVksbUOiIYaijVnFNgHKTLaD9pYcATvhvX
0DgQ7SvDr0WQw228QzWcuKh5FoLDt7fSWb4vSgLZqo00myyMnvIKARTkGveICM5K
5rlzNV+2pZDiX+tPDfKjl7+TQGRdzNrS5MFU3zZyac9HV4BhuXBvgBXPIffva4Dn
8tmlhVmyoYT2XgLz5r9R68A0ZSyu8L1QmFyH95wTvguiw6WLDK5DTg54EoOtrFuR
Nfc2VUHrWN0PH7OVlv/hmdn2qmUrz5QO2P53DBn+uiElkeTFVmkxcgei1GPstN9e
UWyhXPFJjApBXXKGcb0I/YqmOl7ECGlVi0M9+u4IoOhawVxltOCaX97Xet9sRgf9
LtU3Zsty7e3wueyGqKDS1TgTZl7+VBBI9zqlvP494v++M5WuPIdOk1NvQwjYPl1R
AzdoCX3KvMTPygIvSKQmkoWkFUGYEgXXNX0X/QSZ9/DQN87W9EWtjkquuHeECGJP
YoTHf9G1gnXGx9V+YtvaSTFYT1bhKqHQNRD7079fl2Q+nr/cUzMtjzVAmXUYntws
eY+lzDOkNSfxQgC28BzWjgcgSi/7nFaj/ZZedKV+ljfSo6NedHZxdDUzlo/t41D/
PsEqH8ySzovuPL5LGwzBKOAmyLj/PhOFl26LlRPFu/Jn7ru7Zwck3xWP24P7YRBU
VqzfPV/pEVzG/wSIApBemG6W9O9ygCmEO/9Kalei0RCSqKVF+cmAfoojxuco9C3w
NihnmkdcG20KejlNK2mgiheTHiLUyxUDIhlMFFaPPRSCUsCCu7N0KU2wqYxH8Xdg
MzaTwL4U/bWm/MtrpwDljmnMJTC5UrkHiq6nIIfVFUsrQqgqYavlV2rm8RL/7faW
fXdkE/OMTzbVa20j85CCShd+FK6D24FxlznOJd/DYLqCr7yy/YlPjmZD9n/+kLo7
/mipbg0f7MCgPNALtWs2NOWqY8E5oT8cBdBN47i7q0lyzQJmjFkpWOmjIIzI2tSQ
OwJWuIh2zTsgDyyPnhMVvTlmIZk3vjbm+LzJ1Jt7kSVR1Hlvk9Mua99AFpiBP6NP
hROVsNGMYaaNPQSK7FwP4lWQLCTBErSF5kTt5SIgHeX9vtXDDrbBXKtCxMDlWhxp
MaD8lNzFWRsQrxuhW64GHgsdUOcXTnGWkmi4Cg8lf6AlEeH9gETfqGyYf7Z1Thev
Ujk7+ejwe7hAkcYq68gnpm25r5/6x9OCN/xVO2QksdSPRLAG/+GggbCvDZiuWp1a
g4w5b10ZsQv+eAa3CY60VdT5INHagFWhzP3dWh7X7v2RrhaMCVwhCVAcP3esuGe0
tICsjAw15HS/5GIGPTLeMFIDact4VCvTx8tUnzmwn/Yr0SX6NtZ8VwAs4g2o4qGd
jgrc+c1kz4oDe2j2EvIQIHp1ghyl6mWmIJpA7gNFbz5Zd1jRZ0O57WYYXBbqj7Nb
Saw1eTzFNw6CX6hZ4/PialBMsBo/GBKn4/l7nxf8krTBQkzZKcf6z7sZ2uLp8fZO
h32nsFijyhcmbdRD4AU9JKHGptJ407GAeWV++aJMSafqPwIdaQcXLX5rS+zpgjbt
a8ijsI0p1BjKKRJjM8eHIeLc2Az1Gozck6gTAdfs0qxFqKhKaTEtGun1GKd76Wuz
ASCP2BlwP3cbVWLS5Q7lJJqZY7d401OpcZZm0I3nnYQjFh4+pnSXB/B4LpGRcp0k
u+lJA2JYmkiMC0OeFFK+9mDKoZBdZZozjJ2O/mG0WQbVGG7DpGA0qNc+vVWtkVZA
8mMH9l3rt/4lnrfDq0xdMIwCMB8Q1zyvtoupGVd2CXfTzYNNNfs+6D3OsIRQ0n/R
3NLSSBvlwdbyRYMRl+dA1CKUmvKW9CGXW65lvsnw9+o7upsuLcaCHzTRXXoSlX4q
3YKUcWx5kt/xM5CeCKXVPtC2qBkRo+1cbDd5fLEeOQs3R/05hYHUMQ2hUKZf//Lr
5VgGX/ozoF87gk9NQs75J+j4zjjRGnAkEHqZNpWg52gCOKrd1PFJPKDxJOVjGk5L
lnn59xzgDpUj+LEXxjPdbEw1qQ/iKoL4nnubMEESWasNpdVhHmE6J06LhI20n9EE
aTW1OmK6OeRshw80ZEK/aJLDDfFimNvT4gQ+BDQLcC3tiCKG9AhOdSYDepmbUNDY
W1ube/SPrOYRErbS23IGJEv971mhd+O4ufPB0x2ZxISlyGLWzFXpxz3eL49Adovm
XZT5CNKeCNySI4wxbPptF/nJsytqxS4gUMNrYLpkXlDjbgi6rQ44Cn8FsYE7bqn8
HkNqvxpdPglDrR/2GbTdpZLjQudsEgn5SKPeExddYOwtnk0/G1k8BG8hkBBBUwdh
X+Khwd/I5FkQks/Dq5d0G69ytyRD3hrgCDwUZlZ30hNlBhUwVtkyzQCwFRe7GKPc
U+QRRhocClbL4xOwSJcB5ap0aw/5IRDpXomtrHg9EcIHeVN7uMhNkdZssDWcwv1j
TM+KY0iSCylW1glwhDxOD+GdrJaSjkVrEZ/SuXtbOp/WB2WSwZj2pBnq7AV1ueDf
JmW0gEajHZIlwCYt84NgakuY+a+tW/SS9/CNupc2ZjcIRW8SdViGtZijFoUbXcpa
7j/vcy+5/tT3hHQIaroI5XtkTTUiczhZ2PpVW5LOpterbmuEy8KGhEnnEoJBO21C
UZZPllIm6XFTac2JB2jzWieipp1iVLuJ1zOCv3fveAjvzhtTBw/S4g/a9g+/xDH3
qWRklLprMbmmaK330zBTdq4bUYQg8b0nrrvBHMb6OVRKcCI8BZhtoIWiqBhMkzl1
PoClUIM1DnM5EnavxhXKGodFLZ+4Qk8mYp46sIiraSrBH+jmucqChKlwXNJlewCD
FccENdgA/L+6Ftx5ZGJyRjyea4yahcjO39R00ke5pRqot3BRWKPJgXa2GQubuHSW
ejb11WbLLjdJTUfvueBVLMlUNNI+t9iGzUbhI/Bu24fvOT6ExKJKG3KQ+riLG/al
TyDhJnNBj7sMLxFeQ2dfB/3ymautrb7bB3GXyarGYYcyz+kIyu7LJ6QMXYPsQcvD
byZVLNWej9/VH7xSK64naGCGMfEuzKNF6Tui1sSwzkziIj6vkHUKLv/FbaNEQUCg
Wc7rEnprpqlEiU+6oucspz+xljjsvPl841pKS0LCWTRPOT3Ld2K35fdSAHEsmiVX
e+RAKa36UJJ1YDUSx0qVBYh7H4wOuU9WpGAmvbCNYqS9ZL/iUvFzqhPfr6GTWRzq
hsWse3/FoQCEDcdMXAyFpOUhEG6ct3b8ziEadmLb63PjJPXLneElzKtpsZ1c1kdk
E7KPU2lUaLkkk2A48ggLI49gOooj9xMEvQvXkoxzKNMLl4dUejgshIvvPFXDKU6P
9zemnsuHRYgSYIUbhhaXfJdijK5AZClcdq/9RDAraeL/Az5+zz+bs32RX7WFhHKA
vFrLVGoSxCHkM5+QKm/33k97YSQ35l3tce2VLquRK+9o/IihwOHq/Lzi/L6qFTRv
xF0v/STRX6N+gDHfZk5ytDcBdEopgHKJc7NfiyOLX1Qy+DCGXbnmtf6fvWtMpnNU
u6MKTtmxzzGxrX1LmxtseloQWo3TinAraGQDJwF0UEnxUz5yhYzmk0l0qkpcSt/N
j9Yz8RLL9p6JNmNx+IPExTsJZw80F528WkNMruElFWipdrygzdL9CNeG1TBRMR0+
+FbIatGEW+avYwI4DrkSMWMHAezPdzUqzzzYOYfN7YgbD4UiQ7I4xDO/qP8lmlRK
Lj6ca0zlAN3aEIAqpZHB8Vp5ZCweeU3146ESn76+L9qXR5k7ISgdVCpClSF8McWi
pYq8iZz1NXNC1N+TTdhb8u6Pi1VwQkBATVxsZYDQodmcorrz8wGLLpvmaQ+FVtMa
0GdoL5L+wR1jXT2P9kjpgpXsASjVE5ehDieG4W048t9cbGSpuVdcHHodR3PcWAID
jQovQ5bsJOyYRA8U7p19P8YTXw3qO3gKCUKMIlh2Tla2LH9E46XG+JTUUQ2Z53E/
vmZUStfWCjjthBLq9tusPMm5eBLzy7vClS7yDZxWIzSNtl5AGO+UugR1MjT4wQ47
MzxlqcagTGECLrAvB/a3tgpKUdSPeCBh2k17uzKHRPHztdk99cNUP+RRmnV7QcA9
UHlFZZGlQJDZvq2YZ7mo3M9LxKSk3YDyS1tDK3O1Q/grKBpq7y1SN2GQdhcFnJai
AY+rkd7lp4Ojsu++x6YgMXk08MaUNs8nlTCIfQ2Y0BzRJ+bqktAsdr9L/7f40LHd
evS+dNgIMSlcHCFzObBfDLgYajs/QxuxMYdRGbF7Z7Fs2zWsyQUuTz/BZ8O69kFO
vUfqNlEh7yuIoa/U7BP1obFHsharP6ggCKvvoLGcmc1fubGKm3JcXWRBG9yL+dN9
o2hn9/abxVEOlqpyFhMSpzVMbEB2HPAsxnWSo47sNGxHoDjNYNjeX37DEVGoCvCL
+9yornTqCqnYQIZ/HPlYWlQyzVUNqEmlFYA6lUYRJZjVFR5e6YV61K9DhhYaMVc1
2wWkr3RMSuiqaXz2JqQOpJ/qFkVE/cepr72FgKd7Vw7hTqSWhagGdy9NVZK38aIT
hxUtI7ase7MQg3sS0QFebMVsxQqNsSUxmu0GkDcBTn014L0iCwOMTiplfVoAaouQ
tWS0O56FnmRq3VN9/XuTXGq9e+B7aEC/VS0WhJTOrN/hJZcTF+LDJt5DDstKWXs6
k/uvhYX4pDT+ZbglPmaAEyP75iE+IYWgJKKxW4hCg8OuZPW/rSVzJ5G9KjaU+emJ
JliFyEEe9O4dGClX+N3M+LEI4d+iZi9EARBMJtYDkFa9Chzs3mnW868yF3dFO1Ml
QFjHKgXfzM2QWteaduF0TV/V7FrSAbd7q7U9El0ebaG+dmtteeXZJCYIn35igf9M
C6Jvpmtn/OOvkDM0aGsG88VvA7VSTu0x3Vwru5OPCjyn5ffQCbAfOrFl8x5WxeSe
pP/0WJTKmRAgj7vixnVRNNoo8DvtdQ+jZrIt0AbQSDk45w5DyomF5bJ8ppDi0xI+
b9eErtcg4wJ/8fICGv6QdaZ9ilv3jEuBjn1YUccMLA+urF8bxCPZbtIk1eDNcIMo
Zechk4rNQOmQdJprDaZSdpnkXTk1EHwLxLfWk9j32BbiJpKkLe3JBC/yBFFYEgaV
juywxK2G5FJWcFPXXHUEfcvMjEP8QYczuQxJPkd6vRlN+kPp89URBYmS8CQrzJVO
d9/Rsp5Ge8L3ik86GvN6Ta+woHPNGpa354AJOyFyfNXFXuh8JIv5LnnYomjpzm8t
WBXVfOipAOzoYAkofS2CBFch9H2xnItKkR7ampuW5UUbFukAA8h2i1sPXLv8xwZQ
DdLvpN8ENqkNtPgJ1EV4wCwQE1OUmBkSLPUZfbD1FruS1djqc2SGV1ZYcQIEzOPU
HzTmwcHVggAceW/mUbRpVq9xoRhjUcDa2drfJXr6+b2tfn3V3Vy8gi8Aud1N0VGA
lNhNVfB74kfCLiK1F39oYH0Tixpenn//S5nFVvwAmRWo8PpyZdmHzb8ogMiiDu6+
zeMEhmOdxOt6fzoJb/1q0l2ShYh5yA7DXXdfmoxdplDVhQpnKq7aEiGSyJTnRmgY
F6nlQCQF6SE5YBWCA1y9i24FkJ14z+PFnap4YHE+LdTwGQlocoRUzwtcYF/8hKEI
9D90TopmKbXhFiK/ZPYVImhAniXjuw7MnI0jgRfYuBf0C3riScpZKLdPAzFWa4BQ
rl8RLzO8te8SasxP6j19FJ1Dy+uDVhOe1nCJra2O32PYqEOvCpvshcVXgPVMPTYy
1MaAz5S0NKvoz6Rqme5Lxb90nUNEflXbDvlH+YVhQFweIM0SQ/j8qe49uy0T81S2
XRZjui+nmxC5jkdQaZRHyfwHfxsmUFr8JX0TZBqBT/j6UEFeI0Q+vwbQd/wL7TFC
awZ9yugoYEAMFLpbrkPA/c2H2bMR8mHI8X9Pg/quyGZivZpXkmrFLNfAZzjp4f3u
qxPal6302Bkefqz/qMtdULAq6v7ySzZ/BA5ETnszi+kog9QRWuz/7M+UHnQDxahY
qooLNfvQqLDmgLunr/GDXR61o79JT75gEvP9jigRM6PrHmYGsXkNh9J+29jFKrZc
svvrRnKq8T4fkbbRYhY/uYiu6vjBSJOWxIeOiJm8rQssCXLAW7ZhQegMwX6UyYEb
8B6sWN9Vmuy7e0Pdz1ShKNiC19dgG/u+SXRmc7Lywwl+/1Sqi56Euy6R5n5YfmAR
9yG7j5G5Xfymz7KZG5KP3p2QWkT9u7xEHEsPS9aOJgCEWIdZfZ677N0uDO28cNrY
TVIEGUnqf9hOtgPeO3/yScMYVRUkkaVrB8iYcZysw0TiQHcP56XRt6PuX+HVjnMv
CqCwOVYxsCkh/wTyMLwyfjBJlNTsq56nWAchUNVfPb7VfYywHliJLTuqcnMYQLx2
n/deSA2872jElKJs20JYdWVEltd8/lh1FQrB5mrxsVkYS/YUYYtzAkn/XDkv6yBm
jAvXcTPBoCqwBRgOCqIDeO272T71VniFDb45OG3T4genLEdHYhWhNFQbt6ARFCVr
uHXkgc/4QVTiIe2sVfdKTAO0lSdO+rSyVNoMhyrSQ8xl+XV1kRfZifg4Px+U3s9g
5pEBQeRkOWef5hf7tIt1eBHEfmzKRXV9gDAi/kAlfF3SeSQNPtkV95kmJxxxhkgn
g30oudW4/RqQA4rBhIjeDCfz04Tk+XSiVz443J+gTiWPnXQKF7UGaEpxWOu2o0iL
/yzWLJEpPFBzK5tbvFnOaijyrkF0m3rNac6R+jO8QWNzn/NVIUROLjw7t+f8kQGz
rWgzBjKqL4OyxLfJxTwQDmcL2Q49hQks/XJrONHTCOzo5D5r7x+Vr75hDQh/Qued
SoXMiAd9w7YGcplFKx/vCHEQ883NHibEEjbzE3uBTgxK/AvazIG+5ooU39SGJ76s
QrtIS4TE9K7kRVUTFBn/2mzl6lDXdl+b2+ZooU4Ey04NQgBva2n4gt4EMbS0+85M
rFB4e9iggdBqtRUzFoDBEWU1yIjGkqwXucCDSUlnaVhoYhBo9U4rSWuXYavmvLKv
UEmoFMzYK43XTxb6plYvvihqw9ICL4MUrgOh6TSkXVkdQ1nVSstMJmXgd0NSN7WU
nr+RRFU5sRls59301hPLKYCMGn3eW66m3X5qafKlxVebwyagZjTvMS9nAv/ybWuZ
09Hf3+dG8AU37T5ceANaL7XYkMs5WzMctta4hTY+PB3+QrPpq0VNgNUdJzzYUc6l
XTAzYoEQEn2ITrtYOnUInrw78tDbmWyB8v4l19t5PpbGnKVmH3Yvd60+chpxCuqJ
6rA7Hnc/6fjuKIrLw4PmIiZY2Ip0HNCuFH28yYXZDgVxrgqMQzkDj5wrgyo+rOja
sxa2OzrB2Pk4Vo/83e74Lo8IWmHXnnxGFb/mwDVHpt/St6LsVmJMKrLMHmpHZ0Kn
TmkAfIVqxXLwsIUTva4qvXj80HKXgXEHVnfDjDhJ+VYF+UgL32zqdfRbeDvqN7Zc
uR0hmTEeckCF38Ez3qGqr3LATsvyMMSpO4xoLjtf2kJ0B8uqmoFXG4T3OufApKDe
8RBG2oAlu1E4TP3bFmt/HV23R3L5tn1WxLzuJLe0JDhdTBB6v+bTkrry4k32I+MA
gZxcTXL5HJ8DhiVH28/6BVVYyt6NEah1qxpHHSsxktl5CQYuCYQ9ueRBK/VaVZ/I
TB/NxChLiK7NrS7WwjERhXRs0LOEcvOBSXpR7Qo/rpiOM/ZiMbg+S2fd2/9Wz86P
g7n0tJPR5Bu/gfzJi07S6TRaEN/GaRKn5Xy1v4SvjjMMWntDWGu+GBWpKK5U2wmU
XKeRSnK850iViZuW6gx/fHvbdVzPI1ZBXjqIQ7mJZ4vVOR66K1FSFXX/mzqvAaii
IEiXBxyGXHZXHdaT02rS26G56W/PGSqH3YFbzBKYkDrCx8SZ2xsbS89QVjR1X/xt
KHuq57EkNHWmzbO3G7kUEff1XmFq0Xtqal8E2KEp6vB80zd+RR7ddHYpBFCyf/Gk
BoCKRTZi+UERTIYsDXshXhdMypB8iDHKNQ24WIhSlOyFMFdpEUxtzq2MKIOtTe/T
tD0fJerMCPPlgikUPfmFom3gBlH4oiSYTKe4EGBaGvRBE6/jaV11vs1coRJYihV4
rZAn/oglOgFElJ4jUFAheWqbtHdp5tgGqooL6SxrYForjijp8xgheG9/Uy4lzXo+
cXvalXjWdLgXfzisClfTqIG0FKeu6FDaT6wXw4CC82VbQUkT2P8Llr8OWgMqB+fm
GxSGSa0G0O+Qxmr21jJEOVNo4q8+RlcT0m+1VvCwmc25ivtpxVFLrO2vGlaCGhmk
OPSenNWAtengYCpR1WXVAf5c7Av0inHwMFdHhHpZhay/XEEC7jVmOnwcNaM/ZLgm
AbURuz+0+RPYVx66vE2F0gkdxryde+KDzOT6iD7NZwhjSMHXAtwPu4GrjJe9YbZg
9OAyiGygNIXVKtrc3vgfDaAaWrKWja5wIbHnKuv2WlUg193ICibpj7m4RGkvtNZ7
JMrvQq976ZbRUC/85sWZU+Ao66eHXCqQTuID7/G1GidBZQ75uR69oVP0JpQzs4ch
LJTyatYfUn6M4vuML/SPJvTrrH/8eisoAxZMQazCaezIuiI+eRjMjXKglBIg0ete
97+o/G2zi0eOF68zUlwoOFDoZKeTrlr4CwcaUrLuwzlZaPyTQ+66SN8Tg+bU0XyP
6zXHbjGfzL+kaO4/w7SbCMLU7rgXBYSd6rEeLEUEip3jB3FGFkTAvatNLI1+/YNs
u6EpyjwsQ8fJvbVb/+Exjb3vLyB9g9JDit/sbSLcwvN4NHWi2RiWvX6R4wHvyveq
0Tm8k9EkfeLSBhEM2iwXdFHQ9PvVIULLUvpWdkq6xPeMEqjw6AFEWUnxVNUWyoB9
MvIYKTt8XNHQjhORF1eQRcAaR79zWZhvukM43UHlEcpGPJjICKalSoCj8eLYC/yC
LO1oqcMO8SyEJWC0cNxo8qPl4PbFM4IagsKoK6c91QezluWIi10QzDg7/+J95z/R
VNEgiiyWWt4Nb5m5oc+DOTRso31JBjxXZMNTMYa80y6nxdNCwUM6zWtBdyUinQJu
vnSYu3VIvjae+AbRdDKp8MVh3BqxjbJfsu4taqeKuZUwLLJOaRzRMnOjTYdnD/wx
HutPnSd+qn5EY6YODc8cEwhOkB19qcvUdzvom8M37llaWDQko4L7ZJyE2tWyC/Ub
gJfT86Nmk4MPo3JsjRGtN28Gvgz1WOAxwHzRojOKfbVFETNxtV3zbjPwvLWncxVD
+AURYDt0QVg815jJ2Zappo4MGU+NeE1biA6CcKB7ZjDSWKhGQAl1HnXTP2zPVepf
24p22XPkzuHRqc3141vIMgwjK3PmVKtIxULt1KkxNrdcKqWanfvZ4F7djxmCBZVo
JBBoh+8FG648uIU641LFDrj9gm3wszotzeQFynIGbPlcJ+e+MxO78aqjH3vgvQ56
O3fPo95MUdL0MCPANQj3CwmnFmdNRkKrv9fJB36hcOrNLIlXKwRumU5g/t6tvtOn
FJicsVIxlqHojV7ZouRblNd037xFQoWxlrKwBK/ppaeSWYRgvp/OuokkFbC1V8Js
eqO1OSGErqMc/ITB6W3yrsxxzjLEjehdcMLjLcBfhm1JxeBdEYMEJHIeEs5KBnpG
QjPRcPt6Aw4RJpgmFcwnIXk/KI0EZu0uwIT3Yo2guI7tyNwGlipGLdjj2xTRYdmA
sUfjAzdFsuOuYDjW8SRmLimfua/UDoSWGi82YremhxXhX/vnnnXUYkzwRRnbUM6b
lklHivOtQT5BGY9lW0Lh14JW7mZCTQemFFvvtP2R676LQ3UbbsRIei97hY0s0Cvf
prsG1LtvTpOQXoCag9I8pHvLqGkdYKeiDYg9IqFt1d9Hp0JZaInh8bGs0eATcPFw
OEAU68f+XHIDfzDi45eTsxU+nGCi+rr+2qXe7/SOyZS5gwo++94Yw81N7SNze8k7
GVVV5whdURe/qa9MLOzX4EbO4KqWGSHKsFKz18uzLSCl3GRWGY03Ltwa/vTRrqLi
t5b9KtN7eZEwkBDbhvHHOc80jhflEcTIYgmA4nutF5xTFhrplNqv4F8hJCLbXdes
vv4wHdds8+irz8d3dnnCGYFJx0DnMIZW660qTIO5D0WG2HIUCg/FFvfAteiD7Bd8
jnwmWdJOdQSEhEzg0f/7VMe5XHvaed6A5o7W+ElK+9RdGUrsfrVS33XIvsDizfUx
hePgfEhMr3uG++moivWd3Hb2RbCYyh9gDRm0dovbgtXaFZmjGZ7OtTZJOcVG+x00
PnUGDXSlhyZ7oliJYHqGR54qWpogU1L+bt43qBvrk5ImtzN5lGbTEBBnKWpPTlvU
3eWmUctsPCyTiENkzywxtYRSQHXumNwD1EBtbdzArKkuYA06wYsT9fB/Jbx1RZgB
HPoJ1MgQs09UCZ8r1IXS8YdXUV5hVNNNuTpeq2xJB3QFB1uo9Elg6h0EF01SLpgD
9Ljqkr4pYzl5YD/bCXt/+ubqgQ6yqa/tvnXBnmAHwlN1HSX35+30h20kVodPIS3b
6QSsd1aO6uU8qy0t1kXOdw1bBHJkiYbdvHIUR5c1qHMVJWi81/9DlAyErng1DexM
6uqexadFgWf6jWkLbRxHsWqutCdwV7DT6EacUPlX2J5bwjQkvdnMKMg7sbBGiM5y
yOL5RmpDXyWJUB5NB01sM0diX4/Iaujl5wuJu0rBlq5l9WQhr6iPYt83eRkInHc6
QJfLrxKCxXQ+nBKyGtjg8VwCDgAGBOyFqO0LdyQMy6Vu2nZ1WkNILyJFZgia/CVp
XfR9rKTnsSQKml0Igr10zkMj2y70UUwl89x/UmKMVHgIN86RYiPmdUm2b9FrYL1J
+D++Uza4jBEh1q7e8EtPx0bpy1xJ33oXebnCOggw4YZnaBKGx1iLpKKKdjuov5Xy
jbjcg9LT0WDGO5mXWwYZDoi0DuoiPKYFangmwMQLitItqzueHElOtPAnvfC/nHkY
Y0k3Uj8B3mnGSq323L7VFE/jQDZcQZB95KPxRjUQZluuhfUQVytd0EAMFDZA2N7I
RMM4poBWZsA1fojR9SRods9ugxNPP/Iao70vrrOgmcxGS8IXqTAXBIpfAt2u2KTU
7xoIW3CoVIMJMTxzVHDMtzpNWCRBq43phxulCIPTVH/GibDCF15lygYnPJlw9nV0
uX/NgBsSJx3xD/80AI+c0zOSFYQszv1p4614faJjJz++4QIrIIzrOToIFkXvdTMD
nj76ReFE9wptYisiukbBW40G7cw+djSMdGTUj7S3xMdCUs41DSdYnMbjbKTDCmna
F9iW/e+6foh0H43L4Dd4aAWY7f/6NBgYSoIQVEI+cRO1WQBZVMYypWJ2fhVFS7pf
FYg8D/vG74mH7WgsnJ8pdvC6dz4M5k4Bfw+0nHKiOy5nDWLAPX45f408QYSLNdfI
nLwThelLKDh0+NrILJLg3F6yTrJLZVZNnOjdQG2Nu30JWHo8ypP2OpsdCE7oA0Fo
uGE1OGFB/M+rieyBSgpXal754j2RSc7w/oHT3+LyBbTAemPVX10cRvqvQ3mPqHHq
vrS1kyJ8v7PO2VzZSAN0Klg5YWZh4Ld8kfEIBk/ozpbFBGTrjyLATLc3exQPePc8
r8vIDwOQmj7+OSLzseNqA6jBMQp1MMiOU8MUiEte8ic0oAvgyDB+zkGBUQ5R9Ilo
tNtHLrESrhkO9HpFCfJUOy5OOHr+TXMEq8vcJFvBL9l62SoWQaecs7/7hYVQQy1h
5iAUW59Bxff9uCE3qrxqeXnbF7XfFZ2g+dmCXSdGvRu+RaQUF16bjyOFCdDzXQhV
IvQ3u6NtpDUufKbBnKxDyqUq6lOKjXogds14coflyEykeJ2hn/fh2JJc0Zq/YLuk
LGpyyrT/EC2T6RTPoNxIOSrK+IIaBK+GS1ZKeRfH9pmRx7Gs06mV7+nzZ3AazNnx
9m4bL61VIVnOrTEa8GBbxMK5ZGGQ6z+Wc944oZVR3lZBrarRL+o05VDbUK5tIKBL
MVx1D+3v/Fici4V9dAjOblr8h0LI0vNwZ0ksN7TEsNvFDySaa9DKnZ1eRNcn1MiP
esHpwezSLNmpcz9QTNwWxolJoM5M5Z5r0JPv4/ImiVxFsLklNriAZsPTqKfSbKQP
BENuUL24rJ4jAtEPXNbuBVEnoxYSEiMiFmUNlM//mqFm8fYucBN69W6RSjPUoOLI
4rq31bMXXVAUCoku2/YKqcFjlNfBBSBw/lyA6OitADyPYmEofuiO6XlwXfRKw9MH
8iSIL2ZQY6l8Bg30m5TqlhATw6Klptm6j+EP6D5PQOZETKxgoT6MffJXTkjQqKlj
uvvOS22VIh+OpaK4N1AMeFz1J+rslrOvlN9vVxSByXW7jEI1g5PyZfc+OH76jq73
anxSYPC8ivbhioH3DFdE00Wc6/oCty5JWHgLWQsoX74rNklg1CFUuOJ5FYUxmlOh
yogTNDzknCeBa6uTQwdNmYUMWNF+ySLkk0DBFqzysn1VFY04twHQ6Nu834FxMG37
PU2Xr+cjh0QmnQfkPB1doOGJtpPkrsX8ygvi8b1bz53hozgU1XFwVjJnhNwT9X9a
jgEuLLK1YLxw1sGJD3GSQMSf5a+SDyAoG4jIrhVWZlCQXWOuxlHSoVkbOBWkOhE3
0dhVnvcRWwMbwCC6AepRDZL9z5YEAbtz5drwSfUShlWQdvF+lksrvn0O8JUnMOok
4cf6LtQs74MH6OXL/0jhVs7oOLsIqwhj7utXBt4QVHdvTKHr+9U0+og/GjUVUF2b
yMU92TjbSROVQPGznMYCSgXgGjJcZgHUR3RDAacaF9uL2GwAaVUNGagsVffHfb+4
kyneT6f7yDIH8IQUZZxNFI6NSR67ZqMFde4jl0QYNmDlDVLLjyJi3H3p4ZuPoy1p
P+c9esAoBtGSgvHE7wGq5+g8HSVgeLQkj5yotO5PbHQs8H7ZgUKeA3X5W2aytGeH
jt0lw+SQz9JPQpvAxaRJZcTjLK8sGDIvzBv0pFDYN1zyk97Xr2z8l9UYDqiuqqT2
1k9d7myPx+Ca8DcVppe3lN0T5vSo75j+NoCEFJKayp9jsFc22KtGBHPMsasu9uYa
Oo+YEu1xUBt4pZXv73Rujd6/ErsT3RwRuolIU2AnCg6zoxmfH8/pF3rEf9wvXlFN
I0/xcuaERo550U8BzXwAzrtZiC/u+yONEPpCUdgWcd9Ix10BvVytGOAgr9NvKOJ0
QhVo8mIrRiJNA7EwKaZcEzgIhGrh/90vO1mOqzLvbuFg9xDBDhZDuz96i1v9bygg
6mysZVmTkH428D3n0GgYmYD104yq1bGWa98KDktNOc/MGNpuuOuzFZ/2EgO/ssRU
TwpgPYuOg0qaeLRQCcEjVnkFVR0mIuWrVUb/GaDaiFR+2JU1kxR47yaGbZVpMquR
8NlNf5OU0RX5YC95bHo/7Ingt61zP+BLSrObsiNw/rElFnm2VbytjNiyLwUXmYtI
AZL08Tk26YflzkxAIcJRFXvbyerfZ4yBox5n2WvI7C36EoAvRK9zx8TlDkgJEjff
+9cWMFN+pKesodou2wcHqN7xR9RrDqRTtqDiCKvY0Lg5lxH1/rGq5BxfzXUBj2H9
VQakNkwv2iIxqR0s93HpatkmH/ZbaVxLrRm2FyZbTPIgeivu2KFCfldWqqApFFgP
EUyclGOoxJTnRKhRwqetpo/hJCtmyFUtt8sixL8AURbz7ElpVch3F5plGoKfAn8c
a807IRdY5c0oIH+l6JlO33Mys76TyWhPho6Mc3Ja4XrrfmiA+5Qz97ItdySR4zYJ
iSPD/IAt2DmDscW66b4UG3XvhCAxnanoH1gwgRn9YrbJDiCu81Fixp8Zw+l3R4Bx
OcOwmnBGsIfrME0qyLQ7udN8mHFLcyztzntc5aOSTykAGK8MbwsxP6CmkmHYZ3FP
59Fu5vkfJJUoZUNiPIgmUYRllBuR/MvwksP1ucEktrZ1024zubQGrDOgA98AF8Nd
l8hXrhM9dmYvxF+PC9KaaKAifRp3cw6yzZUaRswv317QjU91cYdLNQdbMuVWGJ6y
/i18DPlbGeB5OZATMyjYRFYGUM00KRz98rjusLhu1XE9z0e4xQHJnTjZcbEsOtuh
TTIJwPzPPNEFSH+lOZ9gIPXn3hhpASTdfgUyjzdhVmehSE9CbeqTu+tZW34LhL38
XlmxPtOZWifP8C6Rz9XCnY4hiQhLy96E1ZaxnPgH0F4iw04Vzc9J2/DqN0HpDN9b
XcEc4+m2sAnFFfEoN8j3B/yhJrPDFqvNx96E2s260P/omsGnV/DsRaVwDwH7SetC
KkNtfDs6oHDN4EgEDvvniQYVuP73YMqgLwWa1aKXVsSYq6LYY3E+5Yjl1aoy6bqz
sO3RMmdY85zVD3T6TZKwB4KazEaw7KvbdqOayK/eBsI23y6cIuPMNoUZx181B2W5
l/Vw0cMcSahRZitCQytb+NFTq9z8hXcU8l9cFfoyZhTopRLYTJ0LrStrqwHWtUej
MhuPCiwuZP0dTtPR9k2Vs/Pr74TAyHPu6I/GElLaeY22F7JBJHGzTXWdpRYKEnlp
40SpdPSxesqbikimbHP6SavolDBQy7aHuR4SmrTpuZQ+xBFcoxLaizyAwulmbGuc
4jfJ1dgxL/3HewsiV9RVslCozKwgF/pkPUjsE3IU5b8GEo2NAyNt6EZr0ePXKc2/
e2Nxq4WjztcNRpOqOjXmkeexBKf9QRuNxa2Yj2FS0K7NbzD3FdDNPTDs9qOrUcKP
CmWkRHqPf8B0DHJLmU1mzTOgmMruDtfqq7D9o8rAvH+FoMduv+TsW2b0YLkLhygn
4qUSrTJqJffc/vp/fEJ0spoiR/aHvnx8YyotivvhbS+P/ksi0aUGr7Pd+oOg1q5z
1dR0DKr9x2NG6SMIJzlvvI3cwPmuj/9NEYcwru7ZjzNzeJWIahL2e+JDvmo0x6YD
UGvM6Ok7AV4HRq9HM1y2Dzt5gPX4XkhwoiiDO404OanQK2aBf2f8X16Iz1tiH9nH
4ImhnBfBXY44oHq7heT+VFokzzwhz3tXhL4tSNrfaJESCVKQ1KQvdgiUcIIVCDv7
i0pphkRlBgOBj6EhkQQs7UWhDegJke9q+no66dBDkIkPm9pm+aurKIxvDv1cwi5V
EQO5/LCgNDXQ1oMvewOJC/rv9PwiDO2BEXeQJLtqFRIxbzy40dEkxqccNFQedSbQ
klUoj1+Dza3gd6XXYyATGYQbGh8mMU5t3RYY27QmFovCvhXfCfJsG96LOryBGmWx
lghoDzq5hE2/qBoarpn8Tfns1OsV4byDWW96UcuykOZLUTybJXGDHyMUhMZsPZiM
WnzoGiXbUg0KiIya0xSUj8naXJTl+rS3msm7cuZ9pINaCiZ3oNWDwEhmlGB888A5
VsSJZSEU7DuxjHcLC5VroOoClTKoCP3nHoMP+T6GaNcL1xF2c5Ye7NcnM8+0d+z1
cZTkOlpP6kpeHcZlZqpppbLtP4HOc98fNlcQi56x9FmMDRuK6wLQBsf9PF/stfcs
P91KsWPwLFiLkxTzdW2DkL4MTU+O2Q0c7SSG274t6wRXb2TALyCUx/VqG9pSbuHb
Vzg9ue2iU8JxXdAN3ZtGC6oF0VFtGel0oiiFjugj8zdGleHn4Cld/TengOxR/k/1
/fn2graArRGltENwE7UaRVioTNuzv6xHI3D7YpskXjK7lqOHPW3uz9yLF/3Mqi69
Rxtw/OBqmL7Cyvwt2hLtmENa+7HfGNHki2qhASumddenYsFbT8D0Tsg4CC4JllC2
k+99vnqNTgbYD6lv3tqIdczmGHFloI7UKiNBJ+5whEWnjx+804+iB7DovvuKKR7p
tJyaExXmYmVdlqoa2D/KGtM0ITDzq9l+FGuMN1f0xtMHRcQTOTiBJokW4Pc2AF/u
8jU12S9411l10itNxEvAHG+0cZmGa6ZfLrFL6mBfQfBFT4wbdZtwMf9sB+WzvvIz
CgHtYJM2Z+n8uRseAQLO+N83gsz4kx0OC/wDzdTaGAhUXBq4a9BevemKIQF/lmlZ
LniDk/1NuBR4jRMKdj1Vss557oxWz+CJPNGoHgzttjzDua77sQHmrMmmOLaXgx41
KNQiqgQwaqoBz+NUigJfOvMzVGkzCM5GVZBGtqLXv3wNfZA7Eb5DTJpGE4dZ/obB
dI0hZ7mujGG5XFZFT2BU4oAggXq2t4wCepYNl4kSawg0dpjTqGE8g0HTipvI1hwJ
zCmKIgh/HFi8fFjEh+hNinXQ4DqmJK584r4z6HpXt9XyPOcz70DQOTxWNMek7VvC
gtW+G+5KE4NF1KWUm9yyoqQo/7SceSUoIgRSEtBuWZ6wpdLju7AuLdth1YLaXGnY
fZl0NC2YdPH5wUFxAJHgb6tw2fBocRTAhL1kzVbgavdBgumwK2HcFHSRFoNR1QN4
z/Al51pu0/jxtgr+VoNG51gYVysuLUyeHm9HIMxs2cY9Nv37tGF3fwt7+xA6t3/T
zURa80niPGtSmKmsjtLMC8T0WpDPCTo8//yUXGpTJ8ZJh+iw+JECbdh6mciUKbN7
fetZ/1RRCMvug+PEd2K5b/um1qr7i/kxDWPe6yhXoSQt4Np6Mgy+wS0cSzVz6/PS
nA50z/GFJMRLhh6WMMo/ZgUnwiYFQSy1GHH/ByN2207EgfCdWWPM/OzoSSGIcDYO
yCoYakUg6qo9KUPFRwum6e01Jx5fM9qVyDe1wwHYpQeX5B2TwdC6pEv1YY7DB3pn
7hKw/TNEcmTwmN++i5zT2jrlAM+xEsr7fsRiUaMd2EE8+qyydHdt+GjGLIMhys+y
kTXFOC4Td3X4ADIFIVmJX/UR2bbUrjUJvN+xkiFqT+VQftDcyM2m+qFwexKIB5Nc
Q/KdoPtOe9WHpFNCebBsSXOgSonnKV8I5+CmQS4UX6usg7XPOGvUp6pc6jwIisvF
Q6n7Ukozu3X8iYd7+R98QblsBH9YuWiLwAwygKu/1gjwuj623+4X0uWPJAXxZTz3
QhoMF1gfOXmUBraQDApljDBSC9c1yoCaOHTFwqOiQkkohtFYtjRarLbL27HphJPU
2Ofku7xxiNwmyU+91I7vEBqFSn+Vk4JQ7i7XZT3UeaHzqoxvMyQEuEEaDPWww0fu
1HVcKAItwM9mCuEWwhUorimZWoj8N/0/LhGsdW2OCCE+aM+nCoza1Nb9zKUGRKfm
z44sFs4RhhDAf2JijF+jYOO14BzeXIvZWM5Bno236kmFSSmvgU7+c8MDhGPx8fGg
SQ/M2oCH7tDeVyjPoiQCCru0oQVJNkRkgoLS7wrWIJCqo/Q8x2gR5zORgkrjH8cB
umAolPx62lysPh8CRj0cqojbPpZ6Sg2KFP/z3a3YakJDNlAY9JQRd/s52LAaXIqT
Hz+J9gdcNuk3Q24GcizSZMnZwd1fxdH3kRYv7l+I9qK1hYLcL2NTLNo/d6+PqbnI
ClSPyCVxSnVjMlYxMRstgozG8RYafgQaDPJDJAyNPtoSD5a0NAfaWtBkrE6pl3KF
0M83mGYRATRDbvxVNC3yxV3o+uZ/2p4HLAJWL33ErCHoAI1r/MAtNixDKFMqW6bK
alyKJUvt9GSrubSqnCKjBpDW89+KQzI/uam1uWhiVaUtCafmTZ96M7nFJEHLmjVt
ME2aZA/AOD07+Seis+jjtC/zW2qchIX3hQ1fOzw21Yzc7FMpWb3rjCcncJawqgAd
yZ6cVNuDdNvXVjeBTaSTqKqbXZPyPnVjB2RLN5zJl1XzE2NKFa5tK9sazsRnE1uB
Uke1iFz3cYbeDwXmgmpj9OG6N/u0CsjFtV/6L6HNeTxieHsYsCS+K0fA++TU3X3R
UaFRpJ1fIvnQ4ScaqnpBTJw6OY4rgtS1MfVO6asu+bW3cNP6BOd/xbERfTvJnqvf
5vAkBZAdC9nISeer4lTDa+AQ5gu3l69v7vVRa9qfUBQNscbp57SkWXAX3CW+betK
udvayetcmqfuuw8hnpBNlzDS2LcrPRWBQJoL2NVSdth3V2FUoHOFS0EXv8MHrkct
wKW4Y1fgF0yRNLillslYFL7PIgbhT+qBFHviQsotpVeiYRQmvtez0m0feprxD0HK
CF7E6VxcFeUSzUS98p3GGqVJbSLU9kLYjLVmEugpo/jfSSQyFy0t3ILuhi3CtIW7
y8fVS9d1VKLyYf2pom7OYfFyMpJe9ecgBhtruSThk0+7Uv2NK41Qx56CpXMR1o3x
qIIo8oA50aX66AX7/9XX0ibPdJcGfUOL+CA8fT7wC0Tflqp8ufjtQnqmEQ5HoyKT
LhNo5k8TAXpeNd+unmp/PvN5CGZkRKBlHeTTVkBPocygBzVPMzEPlEeGVdag89LL
58z7dNM8aGWXtRxGc3lc7P69fAWCJ0zDfZyhGUNp4dp7E4aIwCPF1LyX8O014des
Ajr3m0yU0XW9hqwbbAR8QDF0RPggFJjWKLvJk+jttg9hyT/wxXmU8cIUcBpQxuvb
ux36BBq9Oh5waMFaEBqrrPVereCfCvKdFats3QaBJ5mgraI5dnZKPZA31NibbqGJ
Bn4Uj1LpeTs/g5rFSQpLT2mDLjmGNwJQpFTFFRKMqTp+OiV2LYTpTsCPu4okvxpu
Mdi0Y9pAjxjUNlrgbKZej4TkLXRWxbeTX3JCpk4vr+ylsr3n/T1eyZTqPqpwzckN
v0PoqrZY+K2hImJb1qqgRWZzJEhjc/iGINaWG/nqRKLl+5/HqRxON9wPGIOoc7Gx
1ZopMIEXCLAL495cllFe7gD3VvWXotm98PbFFyUGPzkHO4bNtdtmP6q7WFXS2uB4
2SP+ALqkmJIT1Wa2vqi5IENsRMFt/ptf2fvUIq4mo3d72Ac+IvDzlmQT2iZ7udAF
ZCJGqHjklmUUAhno5LgPLGYO5qJNnRMjv4cB/d5j6hc6eeV+NEAWONVnThJ4KiVE
1sZSzHvIqsnM/WNqGi1Baa+Ds2EPLpIu657iDl0YQJ+4MM36+kO8mYg6rVuN/unW
AF3DrqQYGU4CNaLI7zRErXHwpoMaFNybdluMHQmnrMoodI37k1Nf+elpI48vVox5
uwpvYVKJnCFf9W9kAlU8/KaIxk4jhF+WBPZ82dOfqSZeSywgs5LI9rGsv895xH87
92ErJuRc5TSr0N7duT7p/VqD/DC/RvUg3x0aiTFZOshWP9WlX7m2Cy1S2lUOEs8/
9VhnZT+sdiFKumlu0fTbd4IIMp5NdEFo2k+IbaXqX8f4b2hUu8gPmQN9KrN8hoVj
A8tKj78x2Dcx45czjpemtGeYOANPFLyMTZ9kfjD+sT+oLiVu5oYQNgqyqzc1Jknr
fXowdt60UYkM/GQaA/bdl3LK+w2pTXKw05Gwvvw1YX0J+g+78ZN+TQYiPDSAXQub
VYI1DZ2un4GWeX80R+A0MtpQM4QzmkVxmM2P2q0s8TFeRcZr0/pei8b0wfsibLBH
/OKY4XHu9yXlJj6bc6MV6ItdtJdKvjiyz2hxQpg2WzxNy20Hqivw8xL5e6/+CnYE
1yrjBvDBslYZ4n8jwVYsMalEHNhzoWpuPkLXkUtDPCH6JZAD3iUPC4JwXQPFNcDn
492Pwucc95izNy2kBU9Rf0SDGc8EeolLIDrSHLEGmhTMp0DtiV6vPsBfqlUTz198
nYdiO0UeFTgmViyZbcLsyaZiKUdFzN3xU1Qw1e+Pn6iPA/R1hWSSbW2/cZIHzh4w
JBZD306dymPbTx5D9Fbtk7twT13DuGLYAMa0QmlU8oLYik36rLe8ztMC5+nH01OB
49p//zxBX1v/HUoG/5OoplT8n+Bb05N1Z99SSl09hrYGOuP3a4xJxeNajOEIiR9O
Zl1e78v2agICeaVYFAm/mGd9Ae51pOnoBvWj864qyaHT2N9ShQElB/PyT8ZpFC5j
55fjdyL6Fj6PNOoJFeRAOo+LYns9QxtysPgz1zH0hTUH6VuVRW8mdyXcCYMpdrIC
fVy6HA0RQCnGzeNoXhgY3ogn2VtCU+hc+16ESci1yWyMxTAdPgsJZ5h+icFil9JR
CXZQ9oHh3dz6Mjso3bU7xhTX+X/Ufbyr/UzCcbH+nnY50d07A+xwz1LMV63NSABZ
3LTetdzD3oSCYLYNgeGTZahUL3yvJWRZsBG9MPlunpLwDkOeh9ka0WL+OtQUzpYt
66Qcj9snzPJBgJW2dw9Y33uTAQvF4SOmbT3GYyHN4UEwa8nPysTpiL2j0PqhjJx3
JWMjnnKA9el0HFAVoBvuwu4jatj5Yi1NaTFtzE49wJ5GLvUJHEVfirxs4Dyc2fOG
0dVT/dYhO3tb1X0HCwF85nzzedQtv2qDF1Un+V+QxXyaRTafFAMUte1dOAFgdOgf
42v9Brfdv9Skm9HzwOMT4m7xpy+9Ek9LkjTqJzgkJ1lPWKoghk9yCH/OkCrDvzXF
504mtk+of7SYTO+5Mtjmu03VjbOPXCV4gumD3IhWQbLpqySFDzzd3rQtAhtEUPgJ
77EK8a3KxW/8QAHwQSr2SbCyIMtEodN/XtDYC9p1Xc8dttkLW/x4HZ7HHtMkqZHa
mpH7p65tSqd7Mfxi2C9Xmhp4sU1u0kF7GHp7TnfJgBe8SeubrPPHiIIoOvEPkdBx
954FnprmadxKMNI+ptDq6cbdOTj05DiHocLzFQAKy5VrtScgDkbsBMNwyIdhFPjc
F7CMrVy8Enh9k3EjF97+WI0bM0nr7cGi/7O5GqHnI6KRD235Y+GBXaMYceFfmhm5
5nn+iQbgh5MUy3Zze2RpZmT5j2U/SBE+CVFCl/JtImJVHZh+Rf+VQChGjiKxjk3a
2Do5sN84hMbpd61AWayTf7j1R6ENlXFMboKlbJf8fG9Ka/WSJ+Amrqj6GBqLm8vb
F8h9yB8kfaDfXL1k2uIQHtq+BgD6PZHX+lpC4QtGy/h+k0Wo460PekjA6+Od9WTF
woRJ/du2mlMLcyrjToNWf342uH8rHf4LoddZcwfFIVnPIEn0Kl9KpKEA/Z8W3o/D
2AXKVq6JfjXNJjS5aiha5LZy7fcycsUM6+5ihuJu7LGhniS6dPtEYh1GwupSpLTG
o02o268stKPueoHhobFrddNxsWH98aThjtak6NRzSi7d8++sRF8byqonWreQf2Di
pfrIzX0LOGBe3T4Ie9YcCDtCvBB/s7FMmzNxHvKhqUp3Sk2uVSjuZCy/moxERac4
RqOoX7l0j+U4AVZ9ffz1Qmfr/ab6AehWlu1W0fieg73zrvKmlPZA7+6FTWqcgfnv
2QfUbbqnfAhFdvj3c1NPlSrQPzHyUEo92KZozrOPEojlalcGaK4nbkq/+t0hqDgX
CyC8Ym5j6mGmBV2WgjnpfzAPMn7yaIel3kJEzMpcyM9NVCX7NCgnAuRU4y7pnCUu
Koag4plKkDkf40mBZ5PveS+Y60vx0JuJotYwio5I5Q3pYsruT+shHo962rVpDGwx
a6Rr96Rc4zby0W9jL0bwdrtS7w7Qy1oOsJFmhNF2ZEIF6ofnJ7WoVSAOw7Ptt+cR
lu3/qsKQbWTi6RmjfMqQq1+R2zoPgZ+XyjsI5uP3rGmWQwStfQOAICPx3X0oss5+
Rh6KfZuoxaozUqFEKxFSnqjYYdYEnfLHyWHW/WlYN6nXkgm5pfgxG5tFD88HxktJ
PB0QMoimUv89xdWrQHqaV3m3Z4oxwgJX+Bok159x+5yggwvvaNAMKECSD+s/gQAG
9o9KMz1GMcE7ekjf0KphqxHdA0CM1oONlqtMvnxywA2BdLoktKIe44AfRf0cuYKl
FnZAelm6CXuWN2Cw+Eps00tu/rS+jpF/I5K91dkYsnzKiAMMCsmLVurVrihMSkM8
PqboYquHcDXLg74QYQIXdSaMRVb6DQqLm/PKpuuDEwjZaFoCYt5WDwAyIBmfVczn
9yb65EIZJqB6AgLIiEZMfND/C9aRC0yQd0XFGKBCTQan/xWH3GEXy22Tz06qpAT3
qUkCaPx521ETHVJYWVK7okpy/YynImtywXxidyAn/6s3zM7Amdokxakeb4nPu76z
Yvk3hmKMkw8qw9EORLOB8ZqbNX2qvuXXjFMLiIkF1gIat/AUDVc7PKhPxiT5oqwI
O6IfEMkVZFGMKREIaU+agva+4WB5YSY7FeitvqGGA2qhx1c4oDTm7YjKxFB2kiEY
39wxwaYU+mBTlVFt+Lg1uC0zpJF5IDnTJceXBHrSYlHUqH+LSW/05ZH0QSI0RUOQ
/xgFsjOlqoo7yg6lD7X+TsYOCnqBr6j3SgJY5M9khm7Bvfk4CKmpUgee9cSoxBHP
a0BRLE1Lcat2SrQQu3ddhKYqjgTWYzVXsDd+wZ4x32kUnRbCLSxGpYWn9ybvbewh
tPQPjzySUIkk4IhoE69KJnklGx96GC8GtSOqZyTGCvxQQH+PG/ka4LY5zivYE29L
V0NNl+y/+qi8FbmsNQkxIqVYTe1ZcjT2/M2J6vS+jIaauH9xSrZdn11XswPGsH2U
+Hl1x2IU7Ti2S+F3LAsmo/xMe8xLigu25xFdLBY3PVzWitrp8eVYRVqEK0AH1DGt
m+6FtyXoE5cd9LDLk3M8w3oafLW8YZvBZhSmYjk3l8XjWAF7ki6SOWJmNB0/Vc6p
trFED00Braq8kmqsnc1ucTs/96vA68JlckvP9Uca4CUTWCeZ9bwhqDX0LTA/WbYU
Fqt3X6zq4YwnArXiIrajmONjbZiSu3mCkqL1xt/e2JqyNuuF/p2qvCW2t2FJOz4A
WdTzt0bl2ThOwVb2XbkXuI4VL78MOdqpCBqKUsyaS8/8WEDFhj/rVqxSxWmO8kUn
aUwiVGO2nL928Pfn9Bgcwg1Ri2HEjSNVmw5pk95b4yK+/IzDMUdq1+SD3TMVXc13
ZAR6DPx+wa1pJLHtpIfdbLvddQWdK5QMvAJRChcmTAKbCYWxiPhI1pn0r3fbRnXN
Lhr1Y4a/uIRs0AaCsljzbuhp/qQRzLNDz7hEWyupWQxC8oPoBGoINUpP06va53YM
gApn0owjp+FUcaFryiOqVzFq03peVdJ2otZx90FW2gvWuv99CRoeSw5M7+ChtHFV
V26SVQIxJcVIiKJ+azP/s7Mqo+SVrwg8Mm2PWKi+2jrigxBdeWV2haoB44EtkDmB
3uh87CvnMrRC6Frv41/1ewQhZU0orNKXlna9l90v15/ChWNMdgx6gwP/Z3AwZDAy
3HjtlAkf/3jwjvfEQYx74LRVBMFEJIjjwqlF0xMqj3kHTURNRghAnzfgYnB469zn
ZXj277IcNBm9wj0l2ifvkuRps23EgqUXGYmWQuzXwIR5jzdyBxL1v6WAFkPt/W1g
o/I2IuzOTWFtVwTA7B1ge72NZGNtJIqx8Rv3bwKdIkhj6yR3xtqfN6R6Fp2QZYNg
ShuvXJVnoA35oxih6EqDNLI286C4L2KSCIfrUqHUn5j00+NUDHui5p2D/sPrg95C
Od4W5P/f1uBkyuo7zSvsM8Y1TwoWJFNDQG/Jd7ujPjiwQXl3VnaQI5eDIEPlltPf
WgM6p5h9e56tLU0eRO6E9rAwo+97R90Tuwh12D/+pGmG0g1JMhXUs/D4ie5wL/+Z
Y7oOcOk0onvoi0KMgtqgjHVjIa839QA6qED8HkmN/JxFS3YA5USmatWBH0LPG3rv
+2n8M51hLPA6DJWKYMaIgo0BjASjKYNd3+qhpYboV0yxM+MxTYDYs19Vj0TxHgfi
ihh8J+/Raq/vxLao3ENxfWPJcYZ1cHeIq9jgAVHceFXVmhTKpDfzp1MKdGfhoG8V
ODSWhiP/pXlTGL3ismYcjy3cPx302HQGHp5/NJvQT8QVM6rOZTSqzinvsS+D/z52
KTgD31OKV1vLs1IOLAMoavVFq52syHb5lo6A5pL1dH04ZVx9wZRx5mOG0g7NAqsT
7yUvj6TXPnZWIbQ43XePrPRs0EApeQAjEc9x29ItSU7O0pS3jnOTxnySrvpCBJg0
sZYXHzfPHR7OhSYgtku6ZEuqwGcWtQYJ2B4+P6KpOdCCkFBCjHPtnn97CkY9jdy/
/n6wQawyrA3z3Xd2KyyXcWuQZScS0skwcif3Y7bpSEs1nDr5mqkubUTwJkKNy1UW
lMRfp/ssmV4xHoGlgOdH+8S7FzrqZyDMfCgj+X2cp7x9jWjVX1VwnV51UwzNOq64
rWYqVlhNN/1W1AxFcCtEYAHolFhw2T/P6PSm/zFuKj5gQ/vINg39V4O3sXSh7kXJ
Ae3e256xWoZnOiPf4a88zR0O8L1UuBU3jHESoZftmG3bLOphOWbRckDrIds4Ql6O
S+kP51BQJ9W8N06bsNYRE2KUk/LbF0Wt/DLCVqgoIv+dXuxfckvj8yXvBVICmq0c
oZ0VzagO6cDkbmD7DjW6CIFn+/4TuhE0R5vbhJaCxQO/RuPgydxACu8fcV08TuAF
K/t4KLtqWmkqJml2o/M68TBKd+XANYSU+KwrtR1OHNfj15oX8IVw1UCeOuXzkEvQ
QRdgF39xaH+sYZKLA0Wk0wPe7SM+GmHxLxDEqB5B1MgSZpuWJgLw+HxCDa3CaNDb
RPAlOUUWrRXMPOVgJFiy38WUW3Lx6KeQsprZlx9f3vFSFvcIh1CSv78v7BbFb2u0
RNwLjHVXY9+y+vX1m3ubekSCY1d0WNVkUivEfXgaTD0wKFL5VIjHQH+oKa0XHFL6
m0zCEycLG9x1811iPrMxdrwcYyV+WSYL8tUcxY9NqjaXuEpix28ZngU9KLojHndi
JX+1ErJIwGInkhV064CNVoC+5LhScrdTpDBEfVDttX7SYxCZH36/vqjZMCKJLNA7
+3kLC5dUQHK7WLfWQftCje7ihDyy1igcttEB5oFF9VsOGZYD0rEIKQMqAsuNlCrj
26ZYWTglADRIDyHYca7Z2wS1gXj8n7ebTVdByLmg0+KzAS4deR6LAS+hMT09r0Ns
W1MT4Y7Ep6pPWM4/t7cbHOoaM7wyjqfe5gFUJ18N7A9iFc3vLbWk0q7K/ptuMqmO
9qHF2YF7PAhRbTb80ljavYf9IY3qId79Lv7m9+dyb+5XacSJ5GQIWe4beKVE1DdF
JCG4TCYdPxufegdYasefZ3TE/F+s/ZH37gh1B2MtNw/lzsBQgvwzlPVv4qA9hfWI
AOMVGXKx/fYKCGJyaAs32VPmjbAu4HtLlQ35cPPgj+TMwT4eMXlFTFqQKRievi1H
58PtrF7AIRvdT6BIQffLXO9KBQ2DBAapy0wxrZQGfP+Y8t/8uc11fhkwlMf8761i
TZL3aje5ze6d+HcNx6ZiQZLyuAwLAIXj2I/YqZ7PN0lzNFuRmvYaOFWi1jCBnyU0
nFm5Oau+dfGTBAi13VRFKBff/ubXiVEc5oA7CJRJNliNX/Xzpwj6jzJqHtRpxoj9
dKSk2n0QbTDt/NHhW7PrXvGpYvDQXQVRczHsDnJw76Z86Fpe8Ag8C7KP9QC3TPLE
wf+EZ0u1rf7LrAoGoCtX+MGGnsJpoB9+oBk33IIVJgEjkzVvKMaUbxZwYm8IzaHQ
6YFeSRqk9K6+DXobjCv5rpjjuXsZ4i4xBfDCEhIc52+mORotz06os+m7GWp+8cIq
7r2p2Rs7p4b8HJv5RwQnEDndt0F4FoyzkeXMtKmujYArR4dzpUkcoJi542B3JzwQ
mgE6XxKNxl5oKkCjqf6hnyU5Nfi1aFMbQoed+5GGs8k0Jn7iK/gupFn3bBhHa34s
5lI6nFD2VW9bG6C6fJn1lqFNZps/JPVJo/w8slN3q2X//yo6tmcJxBwvvePJTR2s
R/ekuLQdnn8Cq6bzFbKRox5NtMuNmZqXXEVs67ejRZtv8eJizy6zihAcUFQm1/4M
dDD4ZMr03ANl2s1Eh65rIuCk8HZqHU6ZmZwSo78spyQHOMSLDCSQEs2sCgfPakdw
oGMZzk//2Hyt0kKN95xhmxmId/TR7QJkga/d1SkXWVhwR1YCOT01t187CnMsXVo0
3jqAHGzuI3oupdpM49jlchsU6qoC7ugQMCfg1lhTiMCeL3lKDW7ueR36NEf/LuVj
IyUY/ypuQDxyLzqn2BKe/VhZzXgWreEYp0S0j7XftsLYcYUblh/WpZNaztqIbTa6
CExUF6PzyqianIvo8D2YS/jq65wfikzE9Z731sxOwR8xDF2wMdFXNMyrPVjxv1vZ
Bids6F7GG8D9iaQQzQ5s51l7mUunIvpSeFKtnaQcLzujcahD358H1RACLM+MpJdh
VuMiWUR6umW7GDRSAvYvwY2jzyn2A1NjbCYMcvyrksACa/U98xH6n+/iRXNuqtJ/
kqd4Iyr+Nc/MZs8z7tk8i1bt/Q/+pgKeJoXqjNHpIo8LYrjdLDSY5PxD0TIHPpXs
0fbLcsJnNy4P4uc0pbpyMYR/yjMcPQxuMLtSiF1AlCxSfQxHvczYHAsbgHtEEq6k
pVU6GGnPyc7kalI5fLuVLxjw2g+josBJ/hj9mSykarJWlzorI0A1xebaSL0JVin/
kZywTEo/Fjche+OHhDn60SLcGjda8gqx/gDoU51G0tqMDZrdZcMskDb9ntDnm/P6
4Nbq5i/tmC/5YHpGh96ACMpZxeaUSGD+hwX87KTePmqtKgro/Fq205r0G93U+O9u
0UTDFnFxutYGJAZc4/lngc3LxoAv3W/Ib+cslguaELbuZwHvGvX5guC2fhA1SNZe
PtBlUYZ99kaFPpKA/oB9FUotow7JdFuLsLc/YA3ONfPh6joRtNN0HIu7bcFC/n6L
G9Bkl1fgEDKOaMVCdNkELcTwS+wLd7rhcuF+IvYpDwV2WeCPmSdM5Ln/y4/BGCDo
E+5VzBYqNZP5yU4MAMQZ+XnEPWZUWZpyt+tHqxzV6TBmGKVkjeJUYEz4qVlhS62O
h1SFIiExf1U72DFzlYq1obnj1B+Fq8Ap9xhyjV4IeL2KgDqrvCX2g9kocEPFQZ7n
khPnqHq9jednGAbOytYDF53bwOX/aWD+kotvoxNX3xHnF3mxAYwX7b5uOXxTw8Ky
4Ld6kv92AQPdXbE1JQ3cQXQltMifd0/VG6gtOi5Ye3yJBuNJYo8DY1lTS1t6T8vO
Omo39JBkrBStEB9DVPkjY5ciYsAWe6Tfs2cGSQ26mRKINM8bxbT1R2A1AkIaLyky
Hq46xg2W1NOS1pChOT6XaD4ZH1k1kleBttDnqckeOlxF8iLlygapg8TkLQI7vr9A
q8k9sS1cNlpdwAaZXrkO5j/4cKaJkjIUN8voy++xzqJfAlPtERmli4RrY9ylYgyb
EtqDAsIgEYyHb1ajkwkJDLt80EYKFvgCY7KilAhFsQtASvmbrRz0r8UL4qiGWcEc
ANeLQtF3r1tbjNpSf0TXPjjaDwjowpmVx+UKTCpdDr5TCRc1ieidSQhHkXcsloaP
YeNn/+qy2JmLWkJnlTnIR/D7LR7yB8+w33AOyoFdT8+wUz4GewRyoXpC9ZQS2Ika
ay6QASXDsZzgSzNn83GN/OVqZRurGAAXTjuFEOLT0hJ03PYPIq0zwmVfWODrl3fa
nyFxnaLZzYnHrlS2vWnZfkmgOjJqwqk8ri2pkqoGPUvDNiycY11PWgaaSVL8aQTz
+Yxe9W4KKdHl6yh93mnTo4P8jPJUONIkdLkjxH54YaG6ffGDxDuhe+a33IsMcnWu
dfHEc0tzhRsvDTfyAfyJPQZ+0EPbpV43tCF5Xe2Wq/dmkFCJhfLJm0qwRuJ+2jvH
SogXinex3hyaOEvArQQ6dnLjQfSrb5OI2W0vJg3LsMPb8BzOywsUEnbkqC55kgDo
4+CyvX4eNQjqgN0tv0DiUVrn6ojMo7WeNAV7HJqiq5hSHC1wxtINjoRPutBZDUeR
yLaMKRCqLEuSeTmfppbKJlA4IXuEuJG5Xms/mMvzGCg81ClolnJjBLx0pXcoiSFs
H7bL7K0UpqDIFHlxWn3M+a3Vh5R+XHHw4P+cHmcxa4ZHUkQpvapyFV+VRslhnAsW
h85Ht51JcqA55ak4eJVsf8nS10FAoTmZig6X9FdTDAKoOA1RPQUVgiOf4s85uxMx
avcD19+UJ4Kjd1c4v0u/n47jY6+w8L/9OfOsFuf0wK9FTA60G8B9mzomAJkeQJkk
4QBIKeRHmYR2W/hpFT6oU8+g370vEZypMwwGAXfQQ2wFpnWgW8P6asyzKXcq1k4Q
SJHfh9Arwi+9W0BhfKkltn+SQLi59OhtolEGQBtpxQmrmpMgLELUtpLmRnKM/R7m
2qa765sht/EaKbqOpR/G9OFZgyNEBqNH5869D3aDrihUHyJSp8zvBKMgtKQvNEjR
4jR0ROUOR4mnCSDCktelLdQSrCUHY8iK5Dg53hrDVCW1hjoModocyfhVUXiWe2cF
vT61svz9D/0JfIfp3pejWFOO+a40wYpCQ9ovnqb/bSCdOdL0ZjirHHDkzItQEX4s
4wckTd2KhI9Ohs8q7LRVf7JlQcTuxe4zNK11P2SGNa1hEk8CjANVAeTaSfcy7o40
IOPnADyuC5kJ1+n/3pdVo/xaFQUp8WJZ9gun+7qCgbfFRGLMw535S7tjMLJGvefh
lP6HS6RJ318Q8RTLj9HeVvrh8sRlksIPLqsia7KdfuJmQdQFXM+DyiRAZeRwQ52I
HeNqJLvED1EW29mA66sGFDmBD6iFN6EpCmt17R5dY9pnGD1rgYRy4GY51r4pc08R
IiWrLRhzpJLcjH6cG00qhgqkz2M3RFXpdQB8K0YZDPY+b0Y6kOUyIFj/bmnIGwOL
hHDcTQSRCa+lz38Z5qJm+0482OH3pbmU6HF9RPHTvMKgctNyOIznqizfLiRkjtEI
LkihOk48pLU8F/u+Icw/oDurbFYUT3A7vLaiXujtAUOCsi951yOfgDCBDDCguPdH
Xhf2uThHhSPTt7UFR25DTnHqTfO7M66hSvqYna/N9L+66Kt96dhI1cMOXvsz8zwa
MqHdNQzViy9UOs2CS/O/exe+tigRhCSeArKbStSkxJHT3kA4o2SFrOMCiX6Xkk6N
nNPy6uN+hknAULr0xtEqmkd4E0KA2puaD2Z0lhce/rhiUA8aQc1HLX0NrwTpmZ0j
Se2LPSv/XCOn/h0HGKo/0838auy0H6G4jJuJKIatYMSKk/eWvUOwgMtcQh/AaHdW
y5rrD3dA87Rhv5mL+0rAWTpNAvmM0OFcJGg6YaKG/ttJjv4RCZ5UPwtz3mGv1Sjn
Rv+hP6z0d2vRU8Xw6LAiijY5AfXxMviynUn8t84mNKTSWOy3emofp+cjo4+TYjhd
VptE1jBEfSwrU2TyAmkHCqvdCKmWrN7zZR2ft9rjlzyt5w2hx6tJRKO+O/DhX3Ll
vFXmCC0mtSydTWpiwhOkewBh6XQQlJBNjweBmlvEOj0WlBkAtdvukqOxavGP4/vH
R4qUYPacl7DrGXVSs7fMsVhi+YBiglTojcjhLMdnWT8EwYuI4c8k9pVUyAjgD20e
bRuNfAEFEFFCHYGcS5VtCkcm3BsPZWQrqfXkLEHh12r1f9tMAIt3P/MRH5xFaAVK
M6VACO4ilZ2uS7iSjQ5wxw6xhlIbpyX9VoBhzZRdDSIeXw7Pe2ti957n8Fxc3ql0
4xSVT7yua0SgIfvZ4yLm1RiLcXnNfwT1VagEWQ2bM/M6dIlg2mHFRXjfEw6oWuUZ
WEZKhVUbD9cJFlsjCpP6Wc9gRuU0E1QRAj3qp2bl/VS7RvI1xrDptFoxDlNgQ/5E
5GMvo65fEAA1Zxiuy8mmxkvWshxu6XsGGToWU7JnozSeDWQUDQ3MjVVSAgm4qgJn
1NRtZqXZJuIzuy/peeRTidL1XQIjzlC7hU9LYaS+QQ+XDbKwZvdA947agYavj0YM
qJ8hhUklW/qFGUjpsh/+G7CJdk0eYhKIs+VfKjEjwfyAXcRed/oYMEPCPliVAWDH
rARX1Sz+2qbvqBBxpjKGWMtTbF24F+b7X6MbOjcY60XX9bsyuhlh+RJNibwgCNvN
qWx5Rn0zY2XcJ9SSBpu+C52YIfBrK0uf7rUTM+8wIW1P7dvRqbWnpOfAP5eNsTiC
CuMQNA3twrzGRNFYCHlO+390xdRFVpvneM5EzCKx1uExWNq2R6GVPjhGzxF+Cl4R
04zgQoSgm/2dopg/3tLsXTMqSjmclkvg0+I7ekVLcJ8QLPredo9jdjVfzW22psXF
Mq+DOt6MxdlLQOB3BSW6ka8L9K5RVfvt1/78TL/Uj2a8Kn24UC7mHkc0D5X3oWs0
kvvkKzWkaeZExpPgcnTEeQVhYUyDaVyloyhQKCjKC7xVJcIk/Wiua/5DQSWi6L36
T4ylLF74dHI+3n8T++m1IehQ1bjn7wY4cw37doiPaunA85FFbvQ754+0n6KuGjFz
XD7AU3EnVgluvz7e+SRl8j5KRELo/nA1QI+p+eaTS1PG8efykf6RJvymV209709n
GY6bb51N3hb0bEZp7QRTnQq7AlFTjUMLvloBUUYtkFSF99dHEDQH47QKQ5mwjeJ+
N6yIJfm0uyVM8N18qLlxpVtAPPJ5tINVuE0W6bKcEJtyWXRZvDgxiI/YWC8dxB0S
qZG36aTJkH76IhsduJNtfnrDjPuDER/ioaTH7Tt7Hcdh4B9pHqvCtbQG2xEa5km3
bKaL+zVfNeJqTlv+kYvqOo8Ukxijb8qnJ6IqKUuIR0kvOjbFt4p8GBtTE+mx7w/x
zi3Xgj9iSNXU3o69uc7+CAwaMzLbdrORX47/f7yQtxowkC9aZ74EnKEiKZ6nNnun
AsNPGbnK8fhODlk3r+nGb8FVhG66iCQSvCs18pWW9Z8KXe0JNe1SXHAaXUmFkJSH
eB0Ikrd9h+P37yWGJPJFCfdCtsPxqAE+WDYn0XVal7U9F7GMdSUz4QIzTQSXGlkX
lvfXZ5JzEszkk0VK2fiU4Uda/mWGAAcXS/34KcZSJOikUw74WRQ3g2mfqelsqlpl
Ya3N4/2vQ5fiF/ZN2Cyw2+lizxsWjAzgB81flnLZK7lTPZvaTUJ850SWKUnf4rGT
sEf/j5DO2QYyrkqwnM7zxJM03M3ey8wPi5WdOTBGLzsJRNyOye+7RTHwn1c84scg
IxM6TiI3pPoRQ+0IawARe2NXBmDt5cgSQZd4jXZIWq8lLcCeSzEyxyonOxbV27wh
6WPIh6iN/2JyG1153OJt7TzxsOMXizUCIKpjJCHJ3cEJh+iPAMTalY/r9F0vn2LP
y5iCbTQ3tQDRWB4nrDL1spfnZPzlRPC0WEEot8MAab6RvUenOLatV7HBBreN8Pd0
BjIBCPKpEIno48npf7z2TRPr+J7KhJW3uev2+S2dSQWzuZUvYY+2i04BsUHNPbDG
6B66gwR9+r7nsyUaOz1z1Lu+tzfz0RtSwMpGO6CfuRwTsnR6F3tMWOcAWKa+qmAH
W6yLBErLR/8HtlMCe1Ze8j90UcttEMMFzHxz7FSq6fRCeuJ3EOQQ/Vbe02L0jsp8
OSzcxiw61kKKpvAy8M59gLUX047sYihAoneKYgV6ayLHe43H3Gp67KM723Hv9wLv
/SOXfsRDr5jFS5geMju+MTDmLUqeiJZczjeCdWxLBtzgG36NW2CkymyyGYu+Xndr
aNDeH0VNQyoTNHB7rXukZxj6D3d0hMPIoDNTMNieV1FJ8lW3r6BIV/WdzUpPlikM
ydCVZAqeRaUxZgyRavUkYCRCYA2N1gS/cNSnkRpzBwmcVi9hq29r0EgPWeSlHSLu
KAmjygH9d1JKFKNDz4sFAN61n+Fz01KcSNdZpXfp0ylSk68uEmxm6HQ65ZeB/uAc
Vdoa/YWiYBAhMzG5q/MDGRrgDCUgNI+Xg9qp4LyAqUoOanN0s0z9vMNv7UPTvpMj
zo/HIMcF6YyN3emElx2UdDnVLPJ8wKScMgiN9n0AVpRfN6cHFz/vBPLX+dB0g5IH
ObWLGk8Xu+lvuVxu4jTVUtBvN9DKRlxd8xCYG5//4Y5C0lP5H623uBP2jnSJVM/L
oQFjUDrNj1Wi1tfICyk81BOfIpHMLfhQRqiVLDBOL+1wmZv0+nShox9tIHB4l/1+
RQTJjF6mEDK3XFWrgkGOhy1oLBHeJUcrosdCSCE7hd+PL+9fpSkxOF5j9aFiRkZl
uef8Dl9cdIsoXHpHCcx9sA3gh/SwLKmbfXJ7jfpAfyOIMR8m3a+TUgpQb5EdMy7s
FQPFtZ2J5seRBL7L+V82liQYDwDgcZMPU3uEF7tZw/67YCuGovtMx6A12Qg/P/Lp
159rd4xpcC9RPKkWK3b5nj51wClIuWvdrkkPtBO7A5a385BV0sE5iCPAJ2UjRzpp
bLvmmakA2K2SwG4pjFAD0Jz/OxCKFktM1gr0P67auYbhtDFCiJ+PwU+LzG6vB9f/
/pigAVLNTrNgquXJLPxU3znbDBRNae3FpMCGxwwl7JjLfyKfJB0Z7y7zahaOzbOJ
bjAWvzHwG5Lfbtu663q7fnyu9zrN7fwgf8EopXsUsK8H1kynLmmSI7CPnrGeZfkN
1PKKPOzMd6NTVOCMyXg/AjJTnmY/kkWEk9xCflfV/47GjmCK30p3MfJBeZfoBAsA
FgKXDZl1BNQQR1+D5vBrPpwndhJXsk1CDZMeGisomfDfVQYftVbV/NQCPOUYdx8f
jdeP+4OR8shGZPwk74wS15RKg25W2mH+TxXbx2zvu5JM8sFcV6t9C6JKhdV6K3Ii
BVG0dkVGGSEdJNOlUbeP4lftvjWBNGQwQ+bhS2brCzNY6wTJBd6Kof7w4J2lpB4q
U0b2egwKl5Oj2iXmWHWxiOMG2XmMhOvaAs5+0iNWb8dwDUW7yO/nrULOHpA/vH1G
OH0v9FpvGuuDxrziyHNPEPibMZrpn8L04pjr5mPKfXh0iikupgfEagxZwe1WsuKD
2g4oxPFnPGM84l7cBwZZdIBqtS/u4l9Y7PQiWXYtlzHASm2uqJzDUAyb5Jk5o+Gf
DUbMVbf7MEVYtut2hclCy5xlbq51bNwZNvQ+9pPcKPAx1CvsJpbaDkzksf/YH//0
q3tVn2QtoO5R6L1/hxkLSlaEA7F89xviRUFBnFfSEgP8cL3+RxX2FY2eXP2OKnIZ
0M5lH8Iif+z7cgZHu2935qExndgAcYgooyMLEAp1WEkios+DNdCYlrT+K8+hKNrm
oA/uooz75vKNEEZxAGtL6wYh3udzPwVkUFq1H8I8417nUz7KQcqaobcHwWGSWdgQ
7RdEo/KBoU1d+a3cliES6Vffy93fNmEmVBSDW1vzE19T387yixsqQlIE5fgI4/0K
bSys78g4C+UqurRAvO5YDdp2vEzXMJo0z3P/EgBDZZXasgtzDjzD2TV1mhqPqQiV
loZbECQILTq5iE61ssqVJzfsaLIM7+Z4LIveXVuFKA47VWNT2wBislXljT1CNZ7F
PamNC0m9gcc+cfRsWaKixxtNsxrNLibD3zTzdpLukDawyAU8i/S3ld7JS/iG3I+O
dCgzSKs3zRaX8CjatHfS8hd2FUxlUxuAJ3fDJGGFq+DV7bnfArpYZJCsqiREcDoI
NunPzt9GqUfRV31+skCLtIvDhMByLBFvxxs2OvggE3JZScGyySnR0BxG5ruJLoss
pw854tk1lJHPz0tlxAof11vmdOv+gMVQIb+cJfXQRbybJVPWjpEQodzawiHxl5hS
U681whAgh49o/poixFOSWbqUfoswBTfHT1Me+DpyfwADgkn/CYd3LPA3ZnfBPLta
rUlNEIm7rrBCWVrZlnrvvGlqU/tqXmJk5nCoQn7yCggWej5CWaMgHzEv1rJpSBea
6i2JLbh80r/6rZxAzG+EkDMGifR8qJKA/DGkHW5mZc/9aWfmySIG6BtmiXR4ECRL
4ecFQr8MIpnUtMjTKSGErhtLjs1axiwxeHwVX6d5fVlzZC0EWZf8GLgh81upemVM
/RwG/tzlUsv5J2pI5skX6UtFQT5oCC34JpDPb/8qro7p8EjlFyghi9JdOtsFBMIi
2p7Sweb5gfUaA5V0PfvaL1BDKiimq+iZ6PUJvYWwiouKaEl9Q7dNtMzJH1MIDXw4
c6elKF50OnSJOIDvD7wVHlXsB5dOlXBh+5+gNPg2ytM+n/pt1VLUuuVW3t9hRs1z
yysw7OOc+qkyMP4eSMCB9E2dgcHx1qMNokM+mrS38oL9o8l5FWqNEiqhVfR4T4mt
CMBA3TH/mpFIAYoNGBJhSN9g67yMnOHfpZtNLoGt5bKA/HWAJkdXEFEcQ+0yRv9k
65+qh+dYpZaNjYxNAuvSc7Yj/AINd/numzYxcgNwbz42MmiwBNsC3U2St7zenH9I
n3zXM9CKdHzYY9gtj5nh7e4HQ+mKZxYEx8DmdKxcYgoO8STlpMyXwgQ/dtNHZjzN
KU8pMnKBAtt808GTIHYBbcqPFqw+IdT8MU3CgsGtAuRmaA5n9KsdQRMDdMUh+p25
s00TuyJNPZmOXFcu5r0M3ImxS2jUB7EyiAJ6JQGBc+quMoVqVdN3w5XStbbVcn0y
IsWYjufuXdE/Q5worW9DCPMP1hSVPKh7/5oHdARrJ5adrJRzMN1Q7MZkoFSHjWyD
mu5keUgrFPDl3cRlacNicoSzrr1x7nyKHT5UdCy4IdvGysFF81j0vBnUPF2dMRJY
D9oEs9EUy8778dsr3bcQT6acTJXcPZ2WGdOhoUjiHEfnnQEAGRIKGnwLqLVkCPnn
DappqvIx93MUgV7uzsNoZOJMBiVBHTMwThp9epd+GXHSNo+csw5lWgLLgy0HAe6d
790/D6wt/f9UgJ8xP+m9x80aoTd3R/aqlAhYJUaoh0AobhKmMEl7fpOOVCns6bhU
alOvLh/WZ2fnGGs0rO6crHS7mfDoKE2XeKDnwfGtdTkZIBlyHgB9CUUY2QkN0N6a
unnyYZVTYPx/K8fRFRrqKOqf7wi7CYXUxOKlpZZHAy92xOswLOPWND6HB9GkQadG
8JJ/F/uvI9BRtcr7VgJdVWKyKWcp8L/ewMCchevxaBX/1kpJhsTypUat/EhonfiS
BpiUuTuTLhp/zHe0tajTjVx3nz7XZi3mJ8YsKAe2nTjGOe0XuzXMz7qk4EGYLakT
SQguUHlKyTortsz95/2RvNKgwTVc4dAxagxrKhn32zReAuzl2q/WwY+j0sI//Bcf
HseWaDoFgpdfM/et3pcWsnOsbfxeOoL3zdalY9nYHjRVNoxB5OGonMCwTB3TBan5
s31nmPHLhttxBjqQBdPF9ac2TLLAlaM1Sx6ceGEDj9nIIxeEK+nuo1wcIsyDgCMV
A0dO4/R5iQICZITxUXbKKp0XK6lQAi2bvM9RHkbS3srqUjVjwlp3Bkv+Li0av4Db
Nzp5Yx0UEyiKqkmFv5ImLH7bac9FvVtiK9LMSh5pl6Gnb95ree5gB3ykWoVTjF3D
ffUqANlyMsfA6XGJyo43h8NEjH+bM6DgO10sR0myYjGDts18io6EKeOp/q2L1g5u
dddW4BKvPdPUYc30A/vau+dP3TWFkpr6Ya4z2zG5ri2oLjQ31QAC53wtoX28DcJr
JeKee1GMhtbJ/3ndFNxTexhmJq0RCLm8P92zU9YKEDaS9gc6ltPyJaTKv8oBiOlH
XCEyEaLlR4bZcci0UBxkdF8/0yLZiTpMdkdjuAv68sDCUszxQL/0S3Pi4gk7lpDJ
M+qyYr33qAm09TOd7Utbk+Kn3ndF8Yho+R4b+d/eqtbenHEZCeUB/Ri7LHEDKGfa
XGnQQ7knNjM9t7j3iVms6xtIOknRvRGqo2RP6rVqhFNxY6VhgBmVtiqoLugXqGM6
JY99DUXszP5uLkwfVSLISeoHO9ZjMjA39V4Hcs5lYuRpRBrWDFXEuzYgEeaoNCpb
JUyYgWk4UdvK8KR7nzjopEnqyzkTrhxUM4L40joUotb75PH8Kq7MX/x5oyj3NEJ4
JSPd12PeV0yX9dNhRPRlwFcibgg7TMzOyGvn+ouGndg8BXhgs7DjcQIrAiOKZ/ty
tdGVMSMOI3wF0U962icul26RLC2y8kbFGbcSnCbjERNcNqc/aRxT6qNY0H13+AjK
a+nXYpclOYl9rZWbOuNbLBAaI4ZFluxtOq0VD+6wdUx74fKaS0D6QghdSZwcS0yH
+nSUJGVwPWoqp8g5L/G0rQlMQctxQfrVULmW1i4Ui/f1sTRr6iwkSdnHdaS2dcKl
h+BOU+qJZ70ZfJRIx7DZyfb54Ll3hWNfdLYWR0X9RMA3LRMXBe+8qPpVaLTzg6eg
YWKdzMRL5mkYw9KLp0d/aK8GAE2ke5YsEr9MPQ+zYKK3fOvqSTeQA01VOILyZhaC
bjEJBK3eyCkNcxKJkgacnxeQCSKHQhDSj/HwAHtvbSUMe6oBEDO+J+SFcNBW5lAw
xEW1oe8SO0V6B+UfkxYH9DF009uUzJlEE/X/zHmXR3WxsPsT9WTcf1jjxMrL0j/f
paUdAbhsczvKyYVmN3u7FAIRJVddwdLWWaiw9FaYeyfoUP4qCetxZITvYC0AcTJn
J+Kq6hTlJpIb48BHArKzCJwYAFG5LIZJsfiVaX+v10rkozxsnb1PTVh5+5+ks8rD
8Nbhi6P5Bbnc9a1bbBFOgcpvOLofUpBsGKVivq4O39IWhqbpC/6M7DVjfiHMSpx3
Nyy7ywyZ4voJC6FJLjdGasZuiW43NinWR7Y/UwoC+DNoKULcJOaT5WtplvIklLyN
19u+6E8qzRpIjoKULxkv6eeSx8c3k2RHwA/yp3NSIyzuBziytEUNukpU29acsu9d
ohjk0v9lQQA9/Y5W5xSw52NJhJ4w2CvnYlQIvAHbVXO8IMWFX85h1OdNlVvdQM4n
m6p2ZX61J6rP+blLMW4vnu5xj726NfGrOd6Fjb0O2Y9jiefYlXV9edKzywr9I8WW
MDf3xI045XmV6l2/mKwHhOB6xkLY7kmCuDTAd+uSResnk5SZ7wVLB54a/87qLNcZ
BcLN57i1/5eu5lMdzZMdelVzo+gM23sQAOYx9GS4n5KCucWw+T5CE9I8zBKcQpME
3KSAxcISQ+mz3xkiODbeyicHldnRhu0jkTs4EbyvYl2qftUTkw/tRcsPdeGSCdmM
YJ1PJ+VbXgP7iW4QByNLKw7T48g6Hdgm3RozpLXVAI6oYPs7dtsEXunEjsXlat7z
jDNb8n6JAVdwmn5mybd3urwiIV/KH/RSe61hRlYYbUJxxtNF0cBBhoDShE3meC9s
1OS3K5n9GdX8+18H5bfiomdrZcavaD5MkDyBd5/HoeDt03N6Ne7aepWeYpUCTYer
rsGNVIK2vrlfgZYtIKvkdQvSEVrTrssm4YiusJEy8ezHUNuCqJISiVjfVjq8hhxA
6FSlumA/DZm1MgmMTDctYAfGJ9zIL4+hSYfzQqMDGEndhgjOWyJl4jTlmzFG8cWM
bZIn3CS16I6sa1ru806XeoGw0VsOikC6Z3zm5b+eL+pgXN0l2ffHNgASG/Kf6yMd
7gBMOepjrAE+z72JNtRqJ1TP4+6gXJ13K5hqOgd89Bn501dgfFe89bkm2zkMpG1B
zIsL6hajONasdOie0R6wVLirTFNNZ6D01tcckFg1PdVkwYq31O5DEhfhOupZ7S8u
X6pihx9qyG+gnQ8e4x3GlmXb0zlj34qQrRcRI+GYPmTUXv9nltnWSuK+bRvNwI00
2jwRfzjvtOIr3GYgHOWuVAFHeKIn514qKh8XxcN8EqSWKw+w9wRXDTXRlARYYh4y
j3dJM+hKDHDIOSvI8UDVj6paCnaBCt7+ZPtmYOxA1YOKbRNLcz18GdDYHRy85IK0
vGjzIbvqUpA2iidJw9F1RgbcEmEk6OTp1vrP9V8gT/lHTqxvxiRb+iCmjrY8cOlf
sAb8rcu87K5+ZsxfTGhkFu+Si7adVFXtYuyMdJyGdtrm5pH3lWuo5btyd2LCAxg0
5yf5Rr67J9uzh0ajTXvHrV9645ys+0xYJXmpfl6NyHT4ulQKT5rDJB4CPLIrycR2
tjm/XWlhfdxYKfnxwbyDWacWZHVMmEDA8t1Wii/j0uk1k/yZ24rlVN//0a9IrzoH
bF3V9tKKtDnPIjXp2AW67ZMIaKIevLKcePD9QpQB0FyLOXpD9b9afP5J6+k2jTyY
RCY1a9Q7WObs5Sj3JWrHxhyLWguWLIst6b8fOQJyD5DDg6I/K+0Fk+d/W7OWDpfR
Mz7jmJi4/Alth2X6lBmRVecKqnF2KbiBD1zldu3X2BMvle9lRfFvDRwCA/+Og1dy
ivlNZfVnq6MX7fRPc+cki7bM4cfkHSBYETkhbE7Qac3JQiUMRH+mdw0kToOX4lUw
hClguT96d3+wdZb8O3N2bzq+jpNg2DKAagHrt5gu3q326c1eN4Toaxw03EQbjGUV
z1aOERfsNrEwzKFQ6DofdBFHPYZ7w7old9FF7leHhsudEpcSfKaVZeHrq5/NF1HZ
ja8i2/kX844DAn1GCWkdD+fA5cd2PtSJPg0qnoteKFgV/Cb/eKOzQOsLwWbzNvPF
oO2Oy9eCKFQLTEPx1vp/XBHxJ4nG5izH9mWsX+Zb4jmW/yzDv7Z5TioxY2hIy0yA
c+n+7DHCVz6yragAWfrM0ka9TLbxVEMKZvWYyGRyDLfv7nV/gDTu9UJlmVc+OL0x
7AOSE7jZY2t5/sBUdRFVOq1azI49QzZ0WTUZ7cSQRrfMZ4c7JM9yA9tqoaeFiOwh
GnmaZxLxDkLDJC/K3TkMJWdDL3ev91cf0A3TG8EqtR2fc6W5dMeFUa2E97Atm7Ex
T2zd2C4wqQaRbF5/QuGG4cJ9Lu+5O2XrpB5DckE/JweHJY2iRxQN9fHlnP8m8w12
7KdczeqBn4dG6vd6r2je1nWg+w1DbGZjTeDBW+nWHaStyP56nD0/893ZMESTPRkg
VujhipuuNspO5dtIDVEVVPyOIV3Lm+jZYrClXD5Zgx1SXaiMeia9xA4Yl9idxu4i
+cltXcMcUxU+UpfEYdC7gp2cGmhSQ6HduQvgyQ9AiB4DJdieeI1GE5BB9YPY9xbu
SeOjxVw5qkxkp7dUMm215A5Xm9VYz/ZCLUWtxHZUEQ5JOSlDv10OkrnBMzp0MAHg
rB4yMcXczOkZ5qAfR/URWGWCT3lq3w84WFNx1I5wtQNW+MsmJTABgeAOTnNAKB57
ZCLqNVLWmo6X3dfBlkUdGSTrZFe3NVR+KiULUeBCtZpJexqWDTdk/80aSwq+sHC/
b52ev8v2Qh3aqyN6vnx5jzzxd4Q6T52yWcjPlPtjjT7CoZIAWnl0NNKE8liQqRiW
R43CiasvrHx9zXcL++m6eUylE0S14NnO7t5+jwK/WTQa7KdYzW6cs5fm5sXs/nko
SySLkH0DmDI5+O1I9j5X+7W2kUQgSpzSQ0LtB/85X+A1MmdH3iUuziN4hNhSMA40
Gtd6tUWT1D2SWmlY1PqKG7YrGo868R6637rU2o/WzZJ5D44FAeeS766K+Ugcdr4z
JdL+CtFWhU40IivqM/J8MSXiwnFUYuU5BMCWxrzA6xk++M42rF1/9IQeGfEKLAe4
JbJPHwIQ/yLws9CmuJx4lbdN+8/fAMUe62f2x+vu86umBiwk2p0moTpwBDAcJI6Y
1QN64lRe2T4Fd8KLien6lPLfLIjDJl9BRfcW3zwcxHXQ0qulxfKAkvQgU+yjIp+j
4S/tqjC+CYekUBCm9f/3JgHNaufb9vYVA3naQiJPFUF50PAW5nn1oYpMEfEEgoaX
akHGbaj1g1EKI0kDKshrg/N4cWSNMGln0YPwLbM+gFoSUGlvBxsjjbbvrIyHV3L4
9ZUb66gniTmeN+umfN6/LpaBDzyn0cbePexbWLSYSmtP3UBn0Z3/3gswSc2uWdYM
SYDtBr/ILaIZlpKPL49hHMhGGh6+tSpkmmTZK4s3v0elDF6B87MRchH+rhvOp6cR
fRWqw07/eqKZwV7DQoGfvqxyjRAk6h550r3LlquB5CZIlRhffwThioGcfDwQn43j
uC7jt+FTSnpwIquM89Z0RDbwTcTgmC6kYVQBjK+wwCyD2Nl8pNiSSw+YKD7ILw22
m5ADnOeDgEP28e0DJbsdRztoBryHSVDPUBe6rzuA9g5iq/RrsUg2g9Gcli+GhfSU
n4CRW3ldYLdr/3Fa8ZXpOYlgD0V7w/2HLGPLy0cFeNztj9g8FDJkRm+vttmbbMuu
ig6CcFEMOYFNW9lD8wpc93R2dHPfl4t8Vy+mIdl8FbqzcQnrSWaP0tZDrSjVp8ce
81N00hZb81X6YirbY6H3ShuAm94zoFj0V93HtZCdzFkyZDfq7hcy0sDCOnIpQFwm
Kx6KOCpdhfuLFJ9icmZZC+B0tmWpusJJfq4q5We2YHkxOj4/BhyNyNOvM1bb5+Oa
Is4YQawdBza1qdWNEukIcLWLkza4xPnzfzOyYokBCwXDrC5vlzjaZLA4f95sA/3N
HxHdYIamT7o4MILpIKueqW9CuCWfjqOIAf5EWM+FiN3AiOmEGCFHt6Fvwpz+pz15
VHxCMMb3GFHrJLRQDbhQZA3MixLFwyARxJrpenDkWaE4vS6Vk8CLi7V6wTi6iM3C
wckutyngOzLkUIV231NNRTy1pMP+7BrexnTwBOfATIsPxtHaxKbgJ4kxhFIy/T4d
8nUnrtJsQIZTt17V7ZJGemx5cxs7TT2K3c+kAdxWLqtJcoAJLOnV1RXqK3pBVLcN
N3RfnB10oTs9N7fKQarYHH5a86f3Gh/JfWoyTx7ipqNi50WqO2fg9pn+zcWtJXlw
dRANp8/XtCs0hkeHaZyKcyRY4gTGhH7stYyzkLML8VvY4ptgyfYNAPBXKHeOYlSR
203taL5Xq/LUmOddyVizHtJUcyXcQBXxvCTYkjTBtDPmf4TMgP78Xoa7PcN72A+L
3U80IVLauQAbBWx0jsLNytY0PMBJUUcZp/u0nTuI+EaczEPzCfVm6MlNPxOvyDz3
IqmiOleCNtYA5DvNPt3vvMzTF9W0ALIzVPily6HbHQcG4TD05XdN1G0jnJqcHe2T
6k8GJHGl7gVY3BxGyPiENJJbPI/uF+YpWSqoZb+l3aZCWuOAyPXySt/nF3kdwJXO
OCWgKhzI4oRFGvIYdZZ1jw8PyouRRhKAJNHxsXyRW8n1FJOUb+SJ4BiByB/EbB5/
N9uXvQsvbeDczHYFeIJSCmWphcW+g0esGXdAOeoCYF83B1U5BkPg1sT01DlOZlHh
zcusD+PUVfhOmnyfe4J/WEc/me60AMDbUga4Q5C/IU84PftPiSpgJFIac0Fvxis4
LwWSAk1BYY9Z3bfrTcdAm+inKN0OPuSHv+mKH0yD6JnPSReqD5Tu68FjaoQjiyQv
a6HyupsDwRHWpq14g/4BKucv9Ic8HWJpU1n7SqSFuzH9Bs+QpjoDLxa5FZQdky7R
Jl+manId35BsNAKaDc50KWEOtv4WCpfhVzDEO3uxMABPaO1otleJTy6zuxHL7TZL
+fPfOVg9uvmhOTYSN2GR/1SrRRnz3CGC57CLbvuEwhLEngKsbR0Vhj7MUzDRL0l2
TQctRiZbjLQpJmGhxiQXCu0oXA7wgIon9VpnhKrCePCVA4/vFY3I2IupGB/DZ/pD
A6eqsfRsqikjm2rVH8xVf1DhGtPV3dtvk1uS3YBwmCMW8VwjlTgOC1vSvJNX8Etk
Q0VqJDnWOj2e4lXrFLgIe/crHm+qrgjOyKkmdWPJrV19IyJzLQapbddGB6Y87Vca
XuX9+zy2qTfhl5fR4KbIgRbIy5guFHDO+FFax2LgDlZ/zjL7cmtZN8PnXnw0HgvN
mP0f/YIVd7wnJ1kaABIcWlGAa+lWPuyfsofDE0Dr+euN7dCoY9haDzg+7RKugQhe
O/qbwptPnzMo5zsf4t4TPeVqo0XvivLlKVUu+1uKxFWGZsTnlvUrXKzJskq+15LJ
lf0MjGtzxr4Q+enmehXr/BAVqYhZbwv0qQDr0pS+hImeM3BfDwNk9LmqgeJZA/uP
kPGLY6oXjseDKt3vAQO4+Y4s+sOK2MItFYVlus+m6cP3OsxXEB6oVxKxOM8dMCRQ
/ruEYhnBMjS3RgBc39mi+USk/poQzX6nKmoUMHPPLxH/YH0dQGzDOzi6JIQywO8B
ytr8rYRjVaKI7J8aL4Ulmy8wzrnymt9cpxT6b2vVkqV77IIzUIK0iKmwm0fOAXZ5
I54CuDmxHoNw29cDulXflnRicg+x2IzJd66z8Dk/W2M/yrRyvZqzT2fXPMrhugFX
YDn4lpNUNYcv3Llm4SRHh7iRLJaGVualRPUPLRGgM2Oj1k0d54zIbweK3ysbWJHH
OyVD4CG7KV0g4gNAbp6IJHJC0Vs+cb4TSEj4+WLWMcQ0pCqt3rCMsAgPukXv2dKR
oh0srjQj2psdKQ3ow8urvLZQt+6R4cvEtMWNI2HPSSQiUT3JmAlB4oRM7wBmgdnN
ODY64JQCgYzr8QNGiz9OZoKhy58qYpOTPNesmcQi5t2h9B7y7K1FBkFg+OA+oGqG
I1TDTVIDnnZiIsKXwqhtvvoVnIeiL3dRVLS6Eq4KCk3HvswzmqiLKn6jaT3WkprB
G5mmdPkkA7MfYdw+frQfuip1iFGEdiDFISJq6OVkBpKBE23/WrQIcT+ZsScKMcJm
oyYapcH//JOTSBenPQyCaovijwo3A3Y2VY7PUH1zeaFtiUITz/UKCSoUM68m5GZP
Kl+/enRNlpgLV1CVis4j9cVVGMm0LLPviHkWkOIBbExcbbQ+3P4S8L5WQ0lwbB/v
Pq7V8WKfpPDJFGVzuR8T/2X92EZWURUzqmRBwqDczYQlC22jRB1zROpt0GwrVSXQ
SiXNryX7BpcHuTjFcDFVB051Rwg8wUygkXbzuEoSsSUjivfc7aqh0GU0xH8LdMzM
O7JHgGHO1ZFNxHzHOozqAbyZ3FYo4xvV737n9IFrzwtSTwZjkysyQa8c2jZz9q5/
TGbdCcOLvsigUyUmoQHPeiZdGtIAi9NVceTN75Aw1GZ6epYsmUwIxsYcyYnIgDLZ
4jADme/pPshW22FxT7LUCUS6RyoTrHhterF3hdkg7epnJKEXoJZt+D7bBsWTdt9P
09XwQOFMxTj4CAs3VU0Bo8JaQ0sGQO6CWfoXPTZRinZz6EF5YjbvqzZFgjLGk5PN
hJW4SVkdxp6kyaSCIFW4qU33aP8rpGlE+voj0Jtsw6qHOWs9UonYt0bxRXw0uFCY
RM6FtXp0o2naOAAb0jm5mf7Kvlj2Ra+A3lMpWY2dVLUTyWP7kqyKnh2M5AonFY4m
9NcJolZvCN632/g8XIszKCIMmhHBotOi2xgc3SXr3V9174/tK/vGdhkEX++MDVSW
NypGcU0vW7d8PYe+zykqjsSOMKrw/p9HH7etL11aPnVpcVm69hrc92jxSvVzgJKH
fdLaP1/zxAcaWcbnEjIWvzTKVzA1PK9qAgtOGTtTgI8VrooQXTk7s12+bpjKSlXG
L/XUp4d0Z3qMLzIdyme43/yt6xCSoWwVB0+yKFfJFZvstPfGA3lB9fVbeUzodMZt
bXfB5XlpCNHb1yoqdZkUISD2SCpkSdbEU+vOoVOvCTXpSDEXBIrvvQDKkBh8JILn
8wzLFBtZXa7C34yTNt9XV//ntso81XpF+cX92A9MEwAAj6IZMN1WNJdTfW+++Z1j
OZMtGyD6uHrOIDKJlXmn4uzV/mI1l16qoT0TpAMGQGQ+LaNAEUCN8dEhXtcgN1Dh
/Hwe9OgdTBP/ITD848IUhMj5R/0LnEcILPcCAFTvktsVOfwzXNu+MvIQj1z+LAY7
Oje6MRwobbTNdZ1MAjykeMLDbUE/eHABd2dSEf06FK1L2cbRCotdLrZFdfo6zJk0
9JY+DNHdtMsYRXhly7e859M+1BHx/zEdOeCBbjEX1pyr4sa8oAkGHoqr7NC8Rjde
kjgLHRUfoYnTcLMghzGg88IyfquSJXWbZ46aVcqGudXASp3S+fnaR31O2nuPwyG8
Ik3za6ymVma1dtRT70C/7PFUmJ8PhM5GpK0UlXeiTsRyBFDrbtrLb6nDyZMxDvxS
SCaPpfsQcpuNeKI4A2TTr4V5oB8CpJME1PUaPE1Gl0oJ2/wan8jS35YqkcFUvx0D
b8vBxqJMPk8fJZgfbGvIxO+xmpywy8iPOtf1kNuSfCuXL/1oLasR3ucPu/hH98TU
jBxfCrwWkfBZvERTEn9/d0u1Q0asyrCzX+hn7ig0RJAT6JVi7uSjUMumViMydmaa
6FBlUGPuDpd+nxI9Z+3Mvvx0Se9QYllWy1njD3oY6Y9ZwpikA7IQuHEIU8B4pXYk
ZuGoDe3Fl37ivKh8VeQH9prEfPyhgHIqJCxDCbbnuwqQGrpgWRxOUlKmed7KQKwy
kyNoc1upV/f2bSwhzGNiRBrAkzwElxbZvzVd6Z+Vuv8HUuu/IG73LmSPlZ2TVRNm
zgNPG8CpLDQM522yM53yYudcNxQtj/EJ2JbYNeRckUkfn8qhAiepXqQXePFvbH1E
lgLULZ1pszqgA+r4RQ/Zii8FQVjSbsy1WpblGcjC65ea0V4WECwUsKGnS9ZD33y3
VZ10qB321V5+PfC8PSZi9trTl9sgsMohKD0FZPxqZCVTFTxLpC9RRZpWXernjvv0
LoXH604M5HEJ0Ij02xPoaN27/fe1FfvtFa4tr/8wxrEEY5//62xMAnOqPM4smFVX
ycxXVsWRgBagBqoDJoD0GFrVHm2SOdkjalQvC/HIGEGc0IxilUd3wvccKX7Uw4vg
Cd1YvlifaMiQ8/cYpzfj/EXs9G0NSbbyFauWbmyDsuPkvWncvSZgKm/G2SPDCHBh
5xav5wfhc5bgFtwY43uDklTi0P8yAz59i7mI70NNWIYndmLO+rFnZwWBuA1BUKyx
kYf3WOTUqGnTQecgg4v+K79DdIEny8fNz+fnkADwoUpVUQ0xXtL0mzMv//CA43aG
hVtxlFBTVZ4Thz9Ja1m+12p3ptBTd//soiiFHw0BcaiK/VyaeQujr95AwaUC1ANX
C3lX3FDEMPjoA0Yf6TtRpov8REVjztIPbAigfrC2V0xEiwu8A433CswMV3d/jjpM
mLPBNSwsHiUkmBR+4iwQGyASawAvDhTwNJgmEDvKj37MM5eQ3bJ35KZPCAHt5qkm
uT6+5eNVmQF33Xc1nivnW6Rmy3tauMV6ct7zy42/+NS8BwzTl9GUAAuJYHtT+1c2
qXiOfG4I8BBYkcHo5nGxba9uuYfNasPXPKbqU6Hiv89gqIvvesvYUxI5BNL154Gq
y0D6wZfZScQCpIgVvN8oslY66E/G8BYMC5FdAE9VXVkk66ENUa1zjzW3ARAxFEP1
V5Ig7K0we6MMrjZM0aMDFRBidCz+fQ3Tp3oBFgkb5I/kbHOdJ68tkN9/XLRo6AWZ
KZj106OV/Q1YwHc2Jndj4gMyc2JS8PP871dUSi19ntkxodYR/Bo9wT5pyqYfYlB3
SZgH3XKJet4oAzVvDcXWN2XnsHxzYm+DKeCQ3/DRpjszyIhJxbQYH4hdB4Z4sy9R
KmS0OsIQqfdvBKo7VannjLyH44yR2WCmXDSkXttWLZRlMvsID2Nwvv+6SpSctttz
B/3cwguppndXjOtQ5wtcN2a4tQgKZmUcb9wt3YgKTUxlrXW2B4ZlVtr+7hLm+VFh
WnStoRamUecmsh/czcmNj5A27C1PFRrlxVGtjxZh7SD0mddNirC28hMaGxtMYLKU
eJXVaVd5Wy95mnymXP6o3zTKzKqThZQBEhKXIdX5G2U16YH+0qiGTYb/AQdrnAc7
A74fRP+Y8xPFrItgat1SA5un73OAGEWxpWrX6frBxHOTa/k3kYI8pPCfelZY/E0N
c8YxPfifkBiak9tBEkHA2ib6uXDpEdg22qenvcu8D9AOtLUQ4pNC6ux7NvTu4znc
yHo4WKWc/eSqgWVK6/TA5aClewH8d+aJO1EtFwsv2qNbOSvac2JoSLz16uko8Ylh
5YkfoWufmFjTfrSV++/E0iK4Gbt76ly5kom0IOuC0rJwfIKywDEdvDF5dpSfrZUg
WAKF1DylCijkrxw9mDUS4VerWruP6KbgWPGUPiTxgZseStKEzu1Cv6ybMs9qKrIQ
F/8Ncg8k7tifs9fan66k+UpY3zxgoYkpf8suJVEDr1+O6x5MIoBHbu+/hsUqH+tK
ozk0vaMRG7rkchO+6E1BCALj+9hak2+0I94IdBxP6lcUdHVm2YT6zSV5p82pxePh
GCQAmiW3TumnJcrqtxTyyCD4SJrnsu+zPN7I03VirYdQoly7xvhdT6tuYR5NotA8
kcAouft0vAkS9OZw1taZEMRG0JG2nGLi5/tjEP9tdQ1tSiR1aELy3dh2xoGpH9x9
clrOj83cZrcEvXxuzw7H4jlpb9WV/OXYFAgy2LPKnJTH9yAxyWOnXcPdsBwwBJez
JjjjUZj5BdYB+YAeWiuzHASBSC1e1/ijxMssXb3zaoPUrewf3v/ILfnoapN++dsB
Eob+q0hzQMvflyg7rNivX/Fc0NgKbdf28bDGirv/09qP3m3QgnPX+9pYI+HcR5g/
AvZOxmds4jY7ORINWR2wjWriiwrxzTjrz79NVZlK8sT1csuk26Q9fEuvobcpZa1+
daL4qoSoOzl2T5fERVpo2WizhF93X3NX6p9TzgURsQlZA3I0WJYG7n6apoyxrcc7
mw7QLn8sdwwt6KKueBDfCCy9VLD57hyYTT2/PXL3y4b5J8RpS5Vz8rjYSHkMmj6j
7u1wgM6pMcRK46AdCqrWI8g4zNbO8EIaBz+xUEfCosob86Etwcwo8sXY/WIrEYeB
NKkzPgY3AXfs6OswEaXMGQhXT4OiIyfgmSA6Mq3ONpRrpmc6ig9eAaFoqrbM09zO
h++QAGmrP6tlyi7Id9bzLm8ac1+JQLH5j/MRVGNc67Up3349eKYtIA5R4+J/PKzd
ZsMJCCAefwfUJcF2BjZ5Jb269pYB7plOyNyO2Fwn8sTjuG17u2pOK8TkzbOeDK0C
zJnhrmB1uaVV5/kB7amdisRaJS97McHkJ5r/RIfOnFM46Cwvt7fw2zHfTjSbG4iV
eDq6ZsZKCnA9FBPT3DY7UzBNO8ZmOvZon2z3yS/rpLJb9CRgeU28YRwi8VN5ngDJ
Z7J6DprszwWzEky6qQZt5V/cSGX7QkkqdUCQUF7B6+Jr7gx8jsweZG6qNR/so3aB
Np7paR7YdUOLV4kjNwHc8sQHm7qjPNpCewSt7AWOxG57TmYBsNCWPwzf62522Pgg
Fvgfyd6foObL2PDjYwLtCWE6IUYjJSevg8yff5jtEet2hgZJJ7A2xdP9pAHtAZ0k
RckvE7noTbjhXyaBEvlwcVMVzBAkSkcOX/9b76iGfziCCJ//gf0YY2oNWBlexnZV
jRVXRQxwVvgYmFxNO6SqYu1hNJ6ZzDal5JP7XT4wV7Tpc9wkj8jrzTHj8WZCJ/dt
3tvpj5FoMEEiNAzmH1cwApD2OtaZ2kWiSCJoaY/mYhxLOeUWaK1mhLpH/AUZnGyq
AV390g3OrihQDUXkuHfqqSuDGFXZF9qnZ1EeQBK+fPujcF4+GBqvEj5rPYqptDIp
qQHGec7AFqV6dL5cw1HCByPzhEcA4lE+RTlRnflTd3vXgku5o67lhjEeVnBJQtAP
VtLDU85uLCGgxo3GsmKHuwfrxz3urxSL4yYv2vlXws9ejl8ovfb21EGlREyRAQzj
0QpEsPd/ZNzQ4sDriwo2XW1cwsp+UItUsQgmMA+2EGXBrWZ5UyngTHZfeOZEJUr2
JnkO2SqeGBBTiyZzQ9KEXRyMY62uUBpzceQdH1PI7c4D+7Tk4iz5V3ygf909KW4L
vbCf4XWC5/bw1myFuxmr+h0EevZTXOxypFeJNK3k7bDH8Q5yDuzdjh1LIkeLSps4
/FCGNpA6eFcj5+gQMQYww+MmzL/7Dwfis30bmu/BVombBndsJI+ad1pcwc9kHAl5
1+bl7A33GCvnexpt3C32XAQVfTgy1Yvt5jyh4kw27agsWOxHNTckQwAZWb02H3Yg
yCzbXFHF8dgwNKq4L7UeUEblcYM1MqXbbeis04BTBujWEULU89wSYS7627yu55WC
Isa2XAQBRyPm6FZIjpf+52sO3/vMq5GwDhfat6tEN8BZP5S4zspo7nhESyqIpZ3Q
051aTCqNgz8vCT4l3X8yVBIMTNHbfHXOXeGdVw4t1N/IHFSElusTK+/zF6Mlu2YN
PrsyHSer3nxdLPLv7zzrG7uBIwT+k0nFkGSs8nv5URhINMlqatES8nzPjCxdICPK
7nMlg1QsqH5Ag34NF3etUZPc2cjg5epvm+YpjFJffHbQUFOnHSv7t/uPGpJiQrgT
0euI/QIxZcwlwUD2pmXypN1ZpZ13mklkMicxOt9SZKI/plEp+fHpSqQN3WPkGiT2
I809k/orWXjVMCfj8DTqGtQmgD20pfXJ0qacEQ4l4iEE3A1DtVNju0GaaVHPBoWn
4pbsUXXfpefvoT2S34xlqQhUYG1yw9GiLa/TAKnVCMfHBxaiJ6N4eWnikLMM606s
Q5+VXwrTVA1KVdA4J3OvUWsPuPdGbkpi3dVUYGGKgVV/fHqMOs/5h0eXzwhVb5lo
qpHNXR+/Rb6Gn2OxBJEvk1XzNDJQnlBVZguFBgat+GEC13/ovFfP6ngkSRAN0JCb
rI8xzri3iPdrNfGosm2O9b9bQT/2H+iEUdn38Ze0WuHcFPFrsmrORhlOYG2W+Wxl
FMcTwaAJMC12Dzwz2VJqFib/tJsIaY/XibLw+ruTSQGhN+B2gdjDkIKs9MU8xB0b
3MzZHMU9GGc+8Dd77P5VMF1Tdp0/53Czo62xe42N0WtNaA3uii9rIivMwYNrW2nb
gjzADI3p2+BdP1yvuNSUbiBbn96sRNUmzmMWgKOagE70E+OU0n/ivEIhgrSNjuMA
GjfhkPiCG+dtypGcFG1KgBJIEbs+B0uVBCBEIJPy6BQQMnZ6ciF4BhVzzpv57Pb8
R2etxdpoLQhtw1g/wOG1p/XBiKEyQWj6dEk31khauPg7n2ulI4zXri/7CY2YO9+I
sX+XLQO3BwwjGAkpQFwuL42OV1n5x8ykEJr2ARQbjIGDjJozTGh2ahKztJeu4UdD
mdn5bKswuBNx9n72vjVh5rd/R8jiBPULsZQZu9wWQpALMusynLaJl2ZgU0c4+Chr
C6ebj0JI++orAP2z064rihST1VxqEFkIdMKCavx/jZR585UIyDurUXUkKDq1GP3g
mCrfBFKI0wTGmhyjjS1KOVSIDXwwief9wpajx5TP8virsZooCXJk/xCy7QZ2OSEZ
lzwNN1ki2+5LrU5csZed0cL7yyPRH6L5DVc94K+o1JJ/Okl2uEUhdqiNxA6aV8xx
L9jjYp4sdFMJ/TthfybnzDa+qBqmCKmy6q2JVXAEB34CQHDBe1il1f/d+xEyREWM
zVd+DNZ4+kADtlE1QVuMgnHCwnw5scUP2w84kH/TjxRIfCQy76Ab00AKWCFBO/ZN
5txN7Xzhg0oFRmCXiUmtKiXmrKEkk+kT6nnpgepnwuEY9nyU7ZSSXSbLvjrVDcpi
6pcfzMo+x5cS1/ynMP97zClLCmeTSJduWPaYCxivBufluuN4QvbU3e3s8fh9PFFb
AgH/AhOsiZ0+hlSqHT2cQ1fU11WiE5FMMU8YaHCSHLoTBn+FgdKZ/s64ZMF7CMWH
vaNDGztToU0zc3CP1ZPkrTqgroJfn+DUaweoNSE9oMo6Iu7fI6DJ76DBKPYjBUan
h1QYsQsOKFxB3ohrEkOrJRVTAOJEdEbfw2rkBSMZcTI4qkAsPvAshtWAbE7tZCYU
zkRg9X67KE8PvpXx0yyIytSEeaVLyuGHT4cXJHpDLZvjNWcs7RCzy0xS2xTFUFVG
zGrsWZXELhmcrw/3CNTbCY45GkQoHbAaZ1JR+yaI5YguHn8jvVVzMOusfo9YytsO
LAYaW0+MU/QQFq7w0E+eUib8JUmTiG4m5Lk1NPiqGq332YeEgWMX0d/nihYqmI2i
Btb7b86Q1FM72bvqOOiqCG4GHEsWTET69gSR6uUNhV8ejVfeSa0u9FxxVpWiNv2/
Yxdhib2/L5uU/D0ONXSQxBO1YxVy+4nyn0Z+u4fjSjE9845VTO3HTGGALWWZqNWq
HIiuCGocpqz/iGBOmCOtd5A/6+1Aqzo+VICGXEEhk17mwYnIJeXP143RQCwokwKy
4oruLp0FIim0dlaD9CuKILFrCH3BAjub/AnE/rwMELu2NaxSA2x1cJ5+iPzKDwsI
9Iqqn6bY32+bUVq6oO4fzzdCWgUhRZdPti6+vFiG9eZNnDtTh1p5NYdxMRVSQCWH
eVX+A0c8GD5Hg8+ecZzLcaFQ+5zlferhq7Xr/SPihi2rVHYzE/67dfo+QB4sb20D
Yn6M0anxvjAFgToOfG5X8XufGIFOT2R18/BhF0eDzO6pI184bRTNzQDtjbfk1zsW
wuHpnk+Z+96nU0l3+O9/Qpwz+TDQj9oQ1Ci+Q+dKxlcgUmi+PZuXgEQumyITToB5
VvB7eQtigDMKl/60Z9GeoEQPlRUcuwS1yYHS3Hg92oERvJi8C9pAQLVCHhnvPhx+
iGuTfzkhtzwHw/dZz2hkOfV+zo/djFB9W8yLpOcWPE0OJzFL1lagHrFyeSmmG4r+
FCOTECr6Q0qn7XCWUT28tsOCJ0NRkIxGgbL8RwizcxQ/rlmHlJ18lBV6FSjDt9l5
rOLZFLQD1RtXYTF75bpnhQ==
`pragma protect end_protected
