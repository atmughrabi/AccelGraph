// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:36 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iYyo5JMGxpGe1e+F8HGKMmsXsBqdEuHBwWLaeJcDb9ynoPG7QD8dXj+HfHZ7rlis
ntCx+DqyzAq0424Jnm8UonCdc/dkkyqe69Iue2bskk9LJw4PPXgGB03cCBT2DfOz
kS+x4qcx+Mc93I1579aj3p3YXuFdOZaizy+Wm+kvYcU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28320)
L71yvcvHnAGRXIxzHdlwx0ahHmsr2i4RBtWPib17cHH80QOyjkl3QjqWRig2T9qX
nFs+5okLDsMk+0qbqeQLgb3Xg01kzQgeUaQNLxmz5mzaVAHmv6aXwYsryj5X6Mkc
rDolP3ogmZlWA2D7ISb6PqFplCeJJx46UbvD+qp43SL+rY88rBVzw29v+oZbnDsR
PbL8xZXzEPhMzn30tNVYWLlHzlTJJt9eMeDNaB5oMnSAQIxhhvgx/eQIaTQHQ9Rj
L4RMCXF/SYJG1oF2sUWLQNZ7S1/hQX3/nRuferlf35Elq86trnHGNHfw7R63fDYY
3aSgZMuorqs+dJgBhhMlCeqbFMieu0Cx6d3IpwtV+uYLJO6MVHu7Ww0Iw1HhTidX
M5+XsK+igLTYS01qOTDjEqtd+QY4ffBkPI4ZdSa3E7OZhWSBNQEdIDftiWBL9FQa
uFOF5ukd7XJrXhXe0mbt1lfrq0uZrGDweo9U/Yx3o2zX6ZoasHIxxZUb8G3UCza+
fAlkvct3LO6wemma2HN91U1cEEtYsOM3iFOO8OtTaHRDgzNMq4iUdNAK64VicUPz
6/v1mxOzP8pZmXzHCVpfzt5cYWc30ZzJ9yMq9hQL2LWI5+343sQ8VZjC6Db/m6FP
81TW/0BtyXrncYVTlgLb2dvlkBFQS3Vi7xUJ+rmk9p/yMKeSc5zhGhzarg7JHoce
WWtrzr8d9KLX/O/4KnsOgZJDdw0K7pd3Uvk9wkfF0M/dKcjjYFaqE80Y/DlwKDui
vLO47KSG+m2biIB/0cVrsZbwIPgasr63n/Kj10JJ26+/ikYIrW4kYAUHiwZ4Mepc
ec3cO9b8wIR7Z0yj7MCob3xBKZWgwM9R3iuvIxeod0MgjrnA4tLwuWfZ1dzfOO4N
w/mn5K2Kmv/J5P/oqmc+/MqTldZP+A32/cvnye7w6DAGGkIVu/2UCmxziofsT+eP
/m23qiKqy42h8IMfS9/GDuGsH5G5I/LA0bmI5i7CqVPR8MZtS9QO3boVaNeZAfWv
vVQfZ2k8Mh0z/7drMCDS1Qtdh2ZFmgiVxJNNTbqpJQbXlf+gMaIS8PK+vsDxzmhc
t28vqCiVf1s1lpzMV+/mV+cEdvBeawZo3YB8LkExjgs7yBRo1Acx6MeBSozqfxle
jUrQepeDL61NFsAybN6SQ0y61ruAW3atgh2DoZcid7OkI4I3DJxjADBKn7XNjeVr
VLtVUt1p6YZjrUbrKpF6+Krrm/6e2POecjt32F0TwChMOJiTMn+gl/fNA6vbphzK
RlOU915EJMrs3y63MGInEkQkC6XWRRDuPh7F46h8jka5PidU1wpiJ8ORGLAFlABJ
pmQJ9Ygs8KlCRRgSZQ47p8q2pfaR5nhrXA0Y3E/xk3CnySXsuTAUk0HdbaLVJMPA
iQ7rZHyGXLyslRYFjXrNI/GXcX+JHencirSc3BLw7QHcOhghI7EwtCrWVlL0lT0h
Qh2STTJHP0CquJjtrNx5DciBwS9mEI5LQ7lWdO3zbq4KEEspoRMV1eP8fFUsiS6c
3MeIW924UNFj196XNywH2AATtPJT/T5ZXVMpxWQO0WSDPnef3hVfW9jyEZkfJ75g
HgOpWkCjNjVB4kTaPZiH0k8tLrDMQxGbO82/9dr6GeMsfef7J8MKDOThE+RXCFC9
dITNlYeKgBNReVoiF6R09BmLZBmNnUo3OqA92V1313oeISNpyU83Kwjyb17wErt9
PMfzJa7vYt7B3oxe3VTFJNb2WnZvdUb2MUkyesp6n0Q5nK7z0mg7nr5jMKvDHP8O
F+mskABu+lHR8CSxuqGI63yygKrrsbYElnKUSCoXBy5idr16k8r5adtYPovhLFZU
m/Fr/hG+2gE2gu8ucrYzEvSfnvBf0lgiU2g1nz5utRq3Nd40OG9GvKZkd0b0B5zd
QYNxWhIFHKp/9dQrKRUp7igzYNPcrzJid64Tz5YtmScE5oYtyyfIgt7tBJK60NhZ
tbcbAU3MhOgEt1f+3vaoFx0KJ3tQAGV+q3hOyecNaA8ayQwbZ3i+C3wkU0kR9VSn
WPcV2FShhy9TxPiKL/niX9Gx/OkM+UbFmpF/kjpzElEHeMutHYFAA97DIxJGi/Xd
4FNaQV9IpVH3AbxXRmqBGywMjRYaxO/rJ1NXSxZ+6dHYVNYRvCavYAQ16siPxv68
qKv/3nRbZ2Bct9b2Zo8dd0tYMVU1VUiRS5pYAfKXPbbUB2qiShYtwJdgvpDFrNgU
QD3Z/kTh7hHwzOpD1HEdgK8lts1qF8BG/WAwuu6HpC5C9qH34qC+veoeUzOvOD7D
mhvn59JK1w15FywoQctqUPBcy0T4nOJBD6U7Ag26fUgS4U64O1wY1kmo3dLTHYOn
7muwAlw0ow1LQf62edt2uVyb3hxHpFLrceIW+JVNIg9IS95pvNNuFOWB/XGOl8ms
BsJ+LBYUPt1MZyWbe91haMzpB6AJ8jPbMXyQE+bAmS/fHLJXYAxD93uqU97uzzve
Ej1tp+15zDsBfC4PVGbOi8z7gStuxVjtH+P6//O4rKBSxtqoom2mn/0jAteOow1y
tDMawGRMrlEmBVYBGJ1pLVVPWFdg+OQeBetcREfucFNJ1uklvD8Kl4ASvfckWDF1
3+SjXfBMEeQE4WhzKKgPw4Kyx1l0o0zZmWZcvoBzAP/ne1bS1gXRZLfqTFkDp9e+
Pv9v4Rr1M4e5lMX23eCyms/JRKdGUmEyEPFi0AxBOTKQvIE3ppwOFOcTFx5T1hc/
1ziENKmk2ZBKg9P2WNdkdYc/z7TiNmS7gO/d1zxqXtMPanLhNgbviy4FytFC66xj
jQnPzNyf92yr3QS7CIVN7eEDASyDBiy8DiVv/6mLQJxV5QVj/w8uNms0ORs/LFQv
guivhmeSnUyeSD612nh5+PLSWSWfLgNPcW7+Pg2jjbQhoFmCaIjYiDE5GHcNdAWh
IRfnVI3QQIp67/cWQ00dsaLviJgjwrGBDzVoQ3PBuAymVhBjGDLx6eR83zYYHzks
4J7Gq5uwNbWkt/lCOScf2ioggGP1WrlYNajWu6Cl0XJMwXOyyMHg5m9MohTdwram
rIosvn59zfOzPkug77dwqjZmUFBQwasgyVfwIiQ/U0xMKr2Qbtb4ZEnsfCuUbN7o
5+qwoFCyOjlIV+5ZSq3q3hb4wlxkWR3gh+qTBlPL0zeAVEK1WFGubtZo6HMLJi/s
0eS8mPrTbiQvBiTV+hW58koNsRTl0KWS6UKuc1J8dV1UQAfCVCG12BimCKAm5HdL
B/SSUNyYYrPTYEvLASGAWsMkFLjY2FXgbcTqL9FvFt1xs3BShxOfAD2RZ7G5cX0r
Lyu5ymJEGaLiGhfNM+diGsRgu8veM7v1YrzP+YtGilAbY6gL40i2EZO7C1W4CRkp
gBSAnqoAdEUW1769yiy2DWYEsfz3ICAy444pLo9RoGqY1tm0rpHl53/1HqhR/YeK
ZvnUbi0AcKUnPqVag2Kux2LolOerBgUkXuhDvplWDN8KLmwBVSRNxf8XITbx3iQJ
iPOWsv/U4G2ApNllmqYz3pzq2sE5uM1iwPAonfwEx1y4zzl+xMbEZYQE08vmO8fj
lWt8eQZIS8H1B/X1L9JLBlSgbJ5Ygab95JYhAhy2410Oz6UvFqmU6LoDOkMAXB5Z
QcHmLwLDCL5Pb20so/Fi3RC71Sr9dDjixYS8Ihv76NrtqiKuqrDRUhJC6fBtw3+9
pcHtUprhVmXdbMG0L8q5mJEWdmNdPlEoUB083HGWf2Fuo8da91C6htys8uKIRwOf
7wXCt0UxNm6Q6i1tm+p43j1mXvZSdrcmyIQND4UsYN6wkNR0jUm3Chi7cwH3SqRE
UskX6x22E7Ypan8b6/sOI6ckZj4PNowLB5QteoGUwCmqqjM7elf2XlmKdiyF2vd/
g45TBEAVcx4t13tRo0C4rJu675XP9PPuMDZ8aAjPs03N/43PG6prwE/HVlzrmvap
ngi+i6gcQCM09/bipdItaWL8o0eT05M89LjJ7+Qd5vXBm/AzhdRH+eXuaLveQQqs
V+gkPzndovuz2eKwHgJL/uDQM6yxFx0PGos2BK8+uTwQ+azatpQLoC009GwVu/Pb
DnbAfTEzwxi0YaVz+Sx33guMIf2DwskOzZr/dha7zjy/Ogs2aQSMESMmGF09L8iA
0SxXhpVaa/JhQ1yOugQmxcYvJ8GZtYKxdVGGdp3oZXVWM3RfcgFICKCpeCtfDSmK
MaJ22vijC+azGpInc6dlj9omJCwx9ZouyvffoVa5+Ws5vxkF/JDMZao9rKcPuyB8
6qj6s3KBeNM1xoR+PoHLG+Yf2CK7SVRIVTG/o8bCuxlJC8gVn4iYblzOKRh7BONq
eUHsP+/1WhZfD5D3Uv2f7NxEhk4/ygqWI/qnYudVxCr75HWE94L1oEJ8JCNXix1y
BbMaHUD0tVj1KyxPVSgtyRmbagVso3eWdIYYZ74kwkFDTJVFD8B0wQb89bImZGEj
v55P74F0632GZbJgDEgTjH13wVwvArpZnlnNAq1LlW1OjqD1F0G6uIoWWf5Vopnc
ir8tQkmfH2s3GhTc90ZwQ13Vmf5EFtTGuRLstJ+8qS9NNs96zD4SelSnJtk5YrcK
J2zDXXTMmL9jgzf9FtsJCQEv1SEqzIJjYotM/eh4LNnAvLRwJOi67iT+oNUXPnMb
p/vH9YCHcKBokT/6VEYYWs9BmOto9UxDau1Zj9ccln8nAluwZNafNBBaVQbaRhv0
u531vGFvBn13Xu3EKNvcS5NkAofphu4lw0T/U7ZpHkegyG68ENwajc5XxWK1X85Y
D3G+zStb+gOTzWkeS9+HVTZ7rVTEFkb+tqIJR8z6c6NKtkR7B9EC718xcyN7jHp5
53tSOgbCYL8C/qSAcjLbWQwpHk6p66TqAFcgUYvOpk7ueRexylFQ20DquoGVrKQu
+ComrtXKMN7VvaweM0yb5WnXCnfweccH/HW1+h6D+OC5aq7lXb2dGPXWuInSqT9n
Su5Ap9MRgI8Jwxiki4+YzYodC+G4fyvFvlPNCqvquokrKTs1FTB13/WkqD9rnUzB
szVttUrp7cNKAr7csJBYsSD9+vLSAucsn7VwUWuDpjGJMfNPZu31TJxEpR5I/Aoi
Q76bKUjn1szUEbUAX+DwuIB3mnv4d1WoglpGxDg1nyB+l1fTWhY9INIrgzHrpCYD
AVtJuSRsEmpqzZcxLC5GhA7LYJSFGLfzgyv/9NkQC0Wsfmgn1KjQXhbsWyh66hT5
0h7TeFwM0EVng4ZBrZevvLqu224EbopGMLoR9UkVOKoFbIEMFe4/Mragvme91EcK
zg+pE89MVk5iQvuA0cL0XdG3Goy0McKGBDWvFzbGqARUJvrlucmWXdjmX50hF3RY
oEXtBDmF9mfplzZZ8TjY7PUJUtnHE2Hsy+nY084J3t4vght8BtzjjuMTfMHwQeAH
ycBjPJYAwMnGh+fvVhzMd/Opz7oeIh7iLQaLmHYYWbc4eqX9cRiDZLJ+I4JrpQB0
5IiUI/hP0ufPDB2Cvzv993W0XuIZLcI0mx4pi/UavVUINIO8bZYGITrtaaB+FpTA
YL3SrIcUto0a4+OForQdgG1hQh/+DyngYfFvgUr082S+QGDfLO9to+MucFArPoCM
hkTLBsPcIFHqh0ZsztP+lcyjrY8J8geGzXbvL55kgV5MEdFSH7/CPmJGVkDBrbrJ
y9bTz/qO7XxG/BrDNIl5hiKDd0rhwufNQKIYoAOSBDZqLF83kF1amc/xQ0PegX1l
kY461opS2t99BR/lNYxgKxJQ1785DgO/jo3Sxd/tNF37N0hNfj1cw88Hq05nOJVg
MIC77m89Hlo96i5bvsQzSuhpigJuHwwHjsyuYZB57lO1xp4BuSJa4+AqGNrI6wFi
RoaiMOSMwLSYip6LD1nTzI8A7UXOKlUD7ctSJcmojg+23DqB8Q9lBmrJBN2Tfged
c0SsmD0GvGS+wyz7OtEP+CroSFMYtfV4RNr/mlnluh82tDrVeG8Sw2kMfmk9ywM3
8GqDNXFv+bOshkfl+qovYif+/bjqPLEMgPo06/eBdY9zZWpkCGE/DwQrG6Z6SFZV
Mxep8vgsZG0WqRv4iDo3FfbxOa+tMQlh97LHqyeD+S4lJ9WBUlHY60pVjcaayATW
rPthhDLSx1w0Gj7swMvwewk3C/lIzBoVpbyOrgipNaBrTwpFqdSZLi3G7hWNZPTZ
lxneoTvjyUaVmODjGONFC1YY2de2I5uDgAEJ36MLQBUbdk2D1p10yVOmEed8pHvj
Vcxfc5EBdtX24rpYwCvK7AEc8jx/hEVA/Ce2Epla3GwFG7cJT0qczMlWvvjIRX87
Z5C08dDCGw9iRjh0l6DjKdJPtXJVPhOoO4yAEPTSsGs0L9c8LNicH3y3bEnVHQZ9
aHjwBisK1Dt+8fc5oEA/4/JvexNWt0bY3Q+LPCbRLLzz2wFjNA0kRyO4l/EdpIgo
ZucIPsSxaigjvGC1whckAjkHO9DA07LyIDtcGm22jBtd2DNqXaJXeJHiMga5gzWY
KOucASOANioEBa59A7OXYLhq4RCfDaYuSaRx4uT96o/flz7xXtcfX0kLmXLCURbc
WHJFRbWODeVjSrXtX4pVPsmq6EdZBFLQP0Y4ABFozUGxxV+dRPK3xC0JUPNoDh0a
cwAi2uZsEYpIinKL6n3KS96TUKKQucnYvr0DaBJVq7MzL/MKVax1Aq4kSuxryYp0
c+/Ov5aoGCKD8aanW5rsbw9sl8Hz6Amsxe4z47pCrv/uF26xqG3VoByDfXwluIdQ
39ukyepacob42lxO/7XDL2Ck4xM4SqwUy7qxfECC+vhP3nZ5NUdHOjFAYahkbicH
Wp4CsVzoQG+kZtH28qWPfbX6WWYY3CUpIwJUyNhXci70AjXf/yaAE++feiHEYrL9
QlauP8LEBIrpVjt7SxlpCpFBJDKLp6Z5TrVzwY5G7mWyxPxRp/ZTtlMSDE481nFU
C9mncI+O1b6qOzgx23QKvHc0dB+sjzAymguG/twr+juvmU6KyCrfpohywbqBBWae
S4DEnvzhDa8veLp9navB8wBbaDS/81nIrHg2StrmUBeG66YW6O9B8h5cJXengSQW
Zw+KrbOFmUmcaXQn+95NP6xFj/RPXYKHV30v2uPdABHzGf/IU0PsmRC6nFaAq99p
v00oZTKbDLVKSTOPqOO8U+N+Y/KHgDuhm+QjgvsmGqwAqzJx3F+yeE+JZ7oZv2EM
veVRPI6ZQ5PFs6KoDWUJ7hP7A1mgZPY67WgNnq1bwuoGVEMYTa2JI+bNaZA+R4Xx
qpVwdpzakHrtFwlPbAR+Z5q0Y8JHvzB4m3y/8UFw4DjtiidPFQN6LJtMVd3EG1ek
mNcGA/y5QosPXeXt/GkwP+ubR8YF6ENYHCkGq7HqZXEdnNBl/1/0Jzkw0YBKmPsa
OEqR1kmDH/0OHQFImuByjsN2P/LUFNab8hPKlhShzc41Z71igc+9ExN84uxNiffK
0ef+tZGIlVvnKyjjpehD2CBXH4dTXL1LwQVG7JHOJvReg/m8Gpocuvc/m1Sv3nNt
cX8Pz/Or2BUr6XYe5zputYlNdlfOsjlehh/gEvH60UO59Tr6CjkH2sFjxmsDZXPt
3hMHI6Kh+aCkx//Qp7w4dBAMeaQHOajbkfA862qbDgpPsUzuZ8iVNY+rhBRuc3pg
RlpARQVFbNIKjUOtdx7HAk/gt+xgritFDB7tQR99h+OAiKI70ZXLMb9skkLdbHwN
XHXFiUMof5FBv34D+2fG5smHnuKK+u9ksH5XLVHYgwhJm1UjtGV8MbkQnoKJq4XR
qMvop6LhB9lZcvTx7aN/rsF2XrLPvVdW6q6n8XtBiB1DLO9vazjNCvIsuopTXpsX
o78+ZvtEXYQ42ki/6etQm8xyYSkbH9yhrNYnlUqaapmEojJy06wbUXHa+2Z626/p
5JCWhHL402Fog3jg/KmoJW46PeXn4Aad0eABjvtHC7RVYsp/0TrjpVL3nMkwPpwW
MGT6AyBKUtVqR+rSfr3YkfuSomBrLnFV7UsmtTdSp28xbhx9363MS44hqkgNW6Ke
sv/9yyhY/AhGJ5Cx0yoDjvVUiJW+RI8lqJ4HbUYx/cNItTDT4vN+1ctI+DIhjRQ2
M9VA+zmEiGp4d3eu7/eiejohE/p8ax50WX+sJ7aBvk6yftaNZ+OrpK718FIqEGT0
ks7QeoeGSghBLn5++Xr2/luAMltqxoThhwacywDCMe7UxMTao8CFvcU9gCKr3eqe
9uO0h9z7jFYJFir/mUP8cXMRIPYdNptSLIGeUn6no1Tx840dvIB9dnbGQSGBfiVO
x2S1gz/qVdT0RNTYvHVVVcUWlof7FhX/rYHdXGSBxiEmSypzB9YzuikPe7PtteLA
/BTOrTwUXmOoirIZDoEJdaqRyO1KP8Le/mh9Imnhplpiu/AfW0aAH5thje/APK3e
01kBypuyEI8RyKa73vUdmnlwmO9Ua1XOWgZdhV1+pcdzOaBIpXnGER6qrdnhvSNg
FFxkWNmC6VT1FCc6iCF/GZ+vqdwEeGnOamaiJKVbUa2ny0sa5clj2bsXYxxxvOuh
gMHAqzv8oqMSOxOnGyM/HKhUfvJhHy7jLlgN5oArlMtjbPb4DptNN0zeVtdE9x6L
PowlWSZXWgGfPs3GB+cP1f48+g3OSsTtiQIlUU0hPU1o89TtmiVgqQmf9HBQlw4K
zXNxvQyfrhT823wcEM414ZurU/+FVvuoQLV8zJ1JUuY8YovmJ9Hj9+HM5QFIN3FG
PY7PZhI6+OTcfsNTRsICgfvupW2OI/rg7PMcO80nu5WPTxc7gpTv4KEZ6gTQ2pUm
e6VWQzNjHs7DaEl1lJF5EuEEz2nI0w+A7IWXMRqCNSyZUEqRVruX5IfcbWUu1GtW
vS4UAwhCRbxkjbOHP7iwHlAiIUaqBfkOVn2HLeoK+aogbr53JKsvmnC4VaUDBm0g
JQ12LcJ15c5W0dAau2XwLXqazJAypHgPEduVNyHTXW9+g5dUUwsHtqDORHg+oHQh
L3kEYI8YlAuwRBUay9LsbCtW96JvdN1mckU03YWjWVJiCDY4aexhMjGQhNnhUKcM
pc2NHrlow6YkaSLgB8N9yOGiFo4MFbLSyRRdj8kyOLMFCwg6R9n+qlubLo+RtZgu
4ZzQ2BZ4ndX6qwnBJdIsE8Phl4yBmYZjaN8pD6NEN5TZzD2N5cQpXP0BzSM0NnXp
Gr3dUaP7go+nmffgse7T04VNjmkVifOqZsqfkvePW3ORQsmz2wxvOwUsjAexy6V+
RHiZEjraa1dV+iS4243Y28AkqbJzJT0DDgdC0c6vml8X/pBBnh4/tq75TuIRUQnM
paCcGWRD87QFbEJbBMpduWTEyHpZ404dkGd0UfmnU0A1DcUQY3pD7ijSzrf+3Jh9
4f7XI10IY4psoLuTJ8SEbwGDxAOOkZL4SbnOMBzGYdltIruK8ypKYe65Lj20LicZ
drPVQubm2k+II0rh2GW8WNlnyTYWAQs+FSnHLcvwKbt8qqf9KHLHdxZrLbk9ZvJX
ZIqNt0TRuSVLuYgMZQZbzzQrn0N22Klp0Ag8c+rN5KXb9MOAPOnDx7SdC2dw/fzp
/tMXwHyXKK+CjcFR7NL8DlFf7fVfXYYy9JZa5r2yrT4h6pWwL0tbBsESUMvqTEwM
Th9C5T3ZfjcQOrixbmDpy7AerLTvXzDtEmTpBY1BLHa+DlENY04Npd3e6Y3QEVsQ
mXe6Morp/3X3y54LLO8/fNJvi8ClAI+skQDKdam+Z4UQCAHqEKHsQmYqu6ym6w59
Xd43yulEvxz1iJkK4MEjuXeMkeDigHBqsxM5ZkzWd++wvSM0ZcDPnscWB9jZ34dy
WpaSSz7JzguIhpMGgOzMWivx3AYevhgXYAdXO68EHDj5Gc3TZe6tE4E5lCN3v4U0
JqkvDh42JyvTAk36+bq6xiiGgEe4KTv8xhs6bQ3TcM35gAH/6hWDJQxwZ/dafhzW
mufABXYzl2hTKIFATdH76SBOE2DZa+LK+cX9fd4D5IF4G9IX7NhG78R9uU3ZtrTx
JfIAHESINdd22WBVdTIXZWDVH8Gj4Qip91HQ39IGGNQsE8mAB/PKujPN6UcS1wlp
4Sw37C6lMGhzywoVE7UMQdWSld7JN/RaDLQ8Zn+BE2Bt/tkyos0qL6Dzud7h7CQU
v9wLysTdaWtK0UBiu9w6hBd8+bMZlSu81E5/Z+xp7xfqdZ6g1WbXKepC3eeBF8w4
2vHz++zmM8nDnjnDYNKCc6hwgJCpOzRUo0DaIzIF37CCiqM6SSJjkjcdYG1Fr26q
eYwKMtvKynb3X2ydrp0OOHUCTHQyTDfOWtMdTXyt0Ouj5jj5xL0gIZDPM4UrdA34
TbwCcAOXv+GPhP/wFd+QjsAV4zetEOpf/fOBSUl7sCq1UyPdm4UwGt5ZXijdOqcR
ItfHuhAynPbpSJDQW+fn/hDV4HC0Crs4j7zIJ4CYeuxqCQ4qkZUgNbnhUW6vh1zU
9Mo4pZ/wH3BR/gwRsiV9Cyoevecv2sDGwZzsOUaR27PPnjBteNyaMw+wyzRVbtEG
aqisteZ7W2jxDp1A+VwwNowEbvWf53MzJrLSztHtxLtBuzr794OO+zMncbzbg3iu
C9hsFYyWbme1TeIIcWA0/Z2bBQxzU1MMK4EgVz3DmZBsTXBpbwg6Yh34hHREoWyu
0FPA/9Z/s/oOnAgt01HImduo2mY93aw/RL1IEbkmq4m9umjXqRm8p/ajoHh6EeWA
pJINeg4vGfcZsO71CB5E9U2tCS6RaM9vhzT2P61uFuKi7dSis/YOlsmYkvkxIewJ
i4T1aUnPILN04Wcotcy41qU9Pr6pzXA4Cj6ZiBsbU8V87x/2Lt7u5St6lYIEHpom
Alehoh0mtayCvUjaZ0LIpI6WI9UxFHbbkzIjdKdkSIkLjbv12wbGQoBAFd9IAydW
gSrSiKxuQDsEkZ7/3Er2OBdMQLyPOFFKazFB2eedVRJ9GjESe/RD6a+3cQ+sFlHL
qtEREGvVYTOCZlbI4Az5IGy5OP44nJVDvBwuvPBPe9L3XwBr57OXP4zbYPJYTh3V
tYGTi8e1a5eQ/lsczUgTORvnB+S2zykbUaNKmDzd2N5zybhQo/tAklBZcwonf+os
+loaXdy5EK4Y7ThggrlbC50dRjRUE4jAzZl3br/E+9Mi5AbatiASeNIamEo+QDpa
4rd+5H6aqCrXOzmpVIZJa4FW6lIsWh07CX2Vs4FOQdigagabuLWNyMYjfs/Kz8mM
Ls9WfBx3XLAAWw/VZfFw/Q46roxXh/pczmGJQE9cTtq4/lqCosUArEYf+deDNzBN
jvaCA4qtVfSUHDZqqPWQxJfjnNhC9xbHLP6YRHASmWyNZ4t5upsKrzD4dA5ctGBo
mhU699B2ONPOtovhwRUbAEni7vf1ZPDPLGghBpO8lgrEkopM+dIS11XXYZWQuncu
doNCv+J/wRiA92bpPOaSHGFEuyEQ66pp5hxwooUochKrLYjrqn/iSiE+aMBkTuJi
3Aidtum+WCTJRGtPbPTuEe7GKMWrxPQZudXstGeHhZ8GynLOoRRX3HC3LhYVwzqz
+nzypxqy+9zEmNV2fvOVwp8Gr3M7WK+h0xayBZR1Ky5mMRHQ69gNpBgKjqRrXekE
C+XcG/jBkGrYgVMSpiGkbc1pEfuzS6E49gGmVdwrJ4nC2Fw4LBuiW7xzX4nYKtMd
ZotdWdL64kYLmzJyKYKwZ/y/+n+8Y7mztynOkeLetZA/WTYih+zoi1l1U8Yh3bQU
BMY+xpl/OikQjEiXOfh5HqyaQdAcRROufnrvLMr+xMa6xFAq9k2YdGDh09dScxlY
S9N22lhwNlGT/I0ZHGfnPaZ12I8sV9G+OIowNbP+Y/o9O8RxJ3IMfnSG2t9VG0vY
kRdGdBbM9z60DPkuaIrGKA5yOZZaRFb/jd7lY753zyaCHm4LWZ1NIiLmm0LiWR1P
hxzGwuPJL7f6P3QaiOxDt+Udkhchni8GiOkwR4umXWHk3pvYU9XYqu6a9SlnpmRi
O4jEk3gg3eYsB8HYFpQOMnLE+NlSKZ/aNutLV655Gk1jDM4U05jqL79yiNOaQIAl
7wbHnEb4trwUo8uupFt8OHF3BfKG97KOGcQO/Ba0k7FSWhNpjXsqswPQESc0hMvC
qfMDNLQp8Enn3Zn4f8+wFP48stiDsIdESg4/XMRfLu7lw32PkWSUl/Jr7MortG78
uN4Mk1MHJKMfpxbDM6ttJwbUmhUwCXFeA/QCK2TRLaR5q4gX61DyLMz7naxmGA8D
kpUBYbyaQti887QCsqR4kboR8wTg3Mvc4rE0UnMDljPHJIDDZ/ptc0FgDv3uGvPO
F58KDKecA9GCajbpEsHZmn3JJ420q7oIthl3u8FoHKDjIN2Fup5EeFrf4mJoqsJ+
2tJ/I0LUKseYHeUFoe9Re9bTLKTqT5t82ANQvIvuQtqviTjHAqf3yQPDcTVlVtbd
d+MmvBvt4PK9xkSS39zR0Nhe8o64tbT3LMRv/Ijsz9k2wYkfopdKieF4gbm9T1KP
StJLE28Djl6OEXP3ienjDnuGkxmCcidPbMzGKYueIwJ/zKG+SwxPG6tD9soq3OwQ
bgu9v91CwiyfTnvmyYSPUp3XGeBXwC7U8dz6ner7BYzMuN3tBdXIlcvk8P0cqL63
7G3OsPHMUvAN+qUrA73WKiwsyow3qU15uwS6na7eTsmhUuSn7pLPESSDiJaI8vS9
+dn/7K18caVzNZUhSH0WvNpI/U58WmM83D0QDWT4uqqFKtuEJrFkgJH9Ztz7C4ly
wck4Eot+in4VwlXZ50Nkvfl/VQJfoAuvdEuuAOKyFg/g2Af2yN8Pvpe3SiG/B3OP
ZLqGD+ye6xONCel0FVswIOVFys0CUyDkAkjDdvBRqu3I/sInd7FJOjVn0GH6tKaK
sVPwC3wkUqmxQvXAXipnoHKrqE/qFF6mvZC00FrFB87u3fm9FC4dtNJlscn5DlSz
uMW9Sev6r8x+2MRg6i4FG96sjR6elYuNqFHaEr9KwrsxRWtFSixTfs73cxpYCSTX
rxbP91cMuRvBJo7QsJy7NiB6M8cFa6jEyVCY5a9HYvW9U3s5I0zkgGsqbNwkSMBE
UXY7SUsFpF5Xxjo/jmcKPiy5Sl2T19+IlVtADtcLYpz6/6sZsvLk0kWfAWUwZ37t
sZSe0vxCDvLXoRzsjfXp5lJR4JMR9zM92Rc+5/TWlQBvhm2zZwrEBSJ1ZQhhh+Oy
m1yY45+lbKWsroldCqY/Ba1uhuTUixUKqVGMZOEatCRUTguFUFzmOVAZijbRjjSv
0jaY0PkMRbFhnUZnJRc5qVFRvvdq+dyQBAbaE2zhu0miIO5SoRcSVbbr7eLqxDxm
/3+5ltawNVvo2zHzqVgdYl0fHYlH7f3q1sr1WDxxO/vbZdja1PMyTa/MH/8oy1Ph
HzoQphF1Xqj3cc865PDIFy3z3fOQofBz7n2YedjTSbzm+Blyh5DTaGWmGsnqpdpQ
KvThx87vkgusiuLkfARCUaMKRmKjQ8Wuiq2AIQLq02GO9NAdObV8c8dcSQBOvPCx
cx/Gj+S6/yIe6EFbGh2uiL2VDFbvX5Up+x5daCMCFZiHEUY1Y/k+6KJNw6OAFj5/
Qh7PKA+Jh41EftWStJdFcJMLz2Cy9KWXcdFST51iAi0gS3BQZSQVx7QTp+08lshz
TekqCwwZZ92IfqARB5JKCsLN5AROqJ0x6ZxBhqdsJoXJ4Id07avHUw/cQtashg4F
FNNAxgpIn2KvZNQA+Gb3zV5lg68/+yK6316OadlLYKJBwQ072GVTzb7tNHgB/Bge
XK74cGPqx3ddpp1kGNqwG+x+9HEEOq8GDSkAfrKWpTcr0YfLeVoh1W0bbQ7KhtMg
L1gNKOYcpCSqSki9ZG0yucMABsYgOhdP6m2YRtHGQRkR+Qd02JzMcgeVnnKcpQ/p
nDs4P6xaOO/R50naFsBjR5MHwWy4j8ROv3oz05igx0E1jODK2ESWjNcMGshUJ5d3
iLap88L1x3OJxO0ZqI1gYPEJaF0n8QGGlgyHfSz6kYwGzdgDN8kGs5/ybjBLZnuh
5fMaeK4ySlqJIqEsLMjNP8e3eWS4QiazKV/ZePe/6gGbs+vAP1lJ15rJK9JgZn5S
tZWAaZx2K5IAEpyopdfZDvte565mkLX7iZGBv5txg27mjEAbM1a+imZ3Wx+rem1g
c+ySXohH5yC8mQB5sOuHUzl8mHL2gbDCFekj4qy91kKD5WGJFJUyQy06UPlxkrg9
Gj8b3vVaBtIUkH2OBD4p9VibxTW1b6bZxaJTTeRpYYGdLT7llYuFCirHL0mV+Cyw
GwakMUCTsv9y5rToBZrButg/inSFCVi27yNRKCFlpxscmbEnjnoTGjf4494KmUqt
9IvJYVt5vW7ZN1/awa3mX+Ufgo1kMQ3EvQpvuhUtJ6Z98VMgECSkID/+3trjm5tG
te1aczBBpp6v8daGArB6AV6sTJymG64ayrA4IU8av2d56MBiqRMIP27QG8SqAUex
TaqNc1MXMGmIkmhIw7nkIWzOQcmln/LLAVydUyGVvCyonxjs8pZoNRBxK3Xl5Don
08GOF5Z7gUcMZzfsMDUqAfoyKlS90n5ruceUhEMajju7edtOTQRMKfOyhht4ut0H
7TO6GNqtVLImojFCLI+oRkrD/GIBMzs3dLmNrAde8ich5YiuvCB4AEg2E7e13xQM
OkJ2cUd/JWbsufQAVuuRIy+4WDy3w0rN+4sVZUatzpOuyIdNllAINWhfpdjifSvA
+4jS3B/+sXXZeoOLnffYFhQXsCM3hDG6s+/3mMx2pW/4VGDsr/UHQaWEx/2dKUd+
C1L8/Ei4SJ4cflWxMvBMVpweqC7V8H9delbQGv3x4WbaRbrLLiSRwlAXe+BJWc9A
VrmS3f5VcUdR8Er/bWaHkfgjYkMIHcobPWWB0AunpwHCcDNmLn63+/kT1xpTUo6s
9bLWjVlm+0/I4gq8s9eSnzW8NQw7NLD2PZmDxbHbY6qVFWkg2/x4/D8JfnUcq1c5
GAeSgE3YRjj8FxaT9J+I/IixHq4hBjR5DsBJfzIIgXs/RnDdj7gdYMnOcuZL6Cg+
FON8QODPdO9Y04nro9rEla9ptFKM7vftufvqdi1enK2F8M//oKn4eu7yKp5OGdZ3
UzPCn7xkfsLLkxRFII/eawTq3VryZkf+zTkscN2gMwIfbp5j5W7yqGxn5uB3vXer
62qhSOUfbiRJXuVfhfSkn7HOnWMtQxHkgzH0NT88iWPrnBj9ds3UTBuqbXPlvU8S
U6SlwY0n+MVcjrKI0QPxRCMS/JulvkGQzRhT6Ryekcl5S+JX/M6xSocdr824LbwL
dU9etlgM2e5Mavg6IbXVENkB9Tzx0okPlm0RRoQM6MJj9MZOes5MU7p4VtlXddZa
Yn7CvjieIRL8Ayo5vdstv3pUoOZvvUBtcICo2FaI8i4PjjbOLaajA6H3xxyw/YB6
yTzNAJhirwNJT/5/78HF64Q542I/SMfdYi3ItHTI/foVIsgct69ZQXfLeEFXiNsZ
F+iyQ2NFbovtZc6+XT8YC+I6hj7yTbWmSXlzrl5mmGGMHCKlGSQArMt6oKqzJjCX
hoPaeXggijyeQ4UsjxaCo8uDY0kBj+bqtfIICLUwSTvm7C5P2wgnHiO8ZwxAjUCr
6KYsYqUlKUMpN3V8y4WOXk0NKIowh4fVQZMgfHUgLO+ui3qlMBQLygm/xH6KJNYy
vD7QlhpXP9wS5tblXdwWVSc2QIQrSCQY+gTJyLdrWljCayV+P90t4NoyU2u4KH/h
qhEW1Zl4pZrHURbM8UIO8MHMU0kP885zuDJQm/A6yNjidwvC/DyLx0RJyXVPwe2c
Cc6InEtn3DsEU0JF/Xcn9wRHOPcku9+qVyE0eKELNkvypJiq50kUJNxTpcb1JBaT
h4VaGnvVOCkLd3Cilf2F64ysqBCDKtw6zXz0pqhLsOrkW+7yzE9hLSj5dvgEsTKs
lU0DtopnnQjrP0AkV6GOsKZoQRDfQ97CkxfduNv9faIU36s0rAG0mYwm4fyYvM6w
isUajSfeAp8FjVbe2f3hTY75hZrWjVZTMNA1cZj+OelVzXty5KBurXHswq45bQdj
wGytii/FDoEo/QLTOkQ5Row4aCluyYE6B/DU8kOgFLobRKNy6aCLWbB3dVZ1wE+w
1fCmaRBOB7Sz3x+7t2T+0roFvRruglZ4xw29HFDLgoJxv+9e5otMQwGy96rzWBpr
IwKpKa2osJyQX4DucaWVWSXMg5QbA7hlwKAiLv79iM8f0AKPRThpmTHuPxELJ+mw
LlXF7opdTMx548ECEwOmQCsOIAAhWmvm5BTGPgwQTECDlqjadBuEE4O5wEjz1zrZ
zNxV/vWxpmQ4TcPdBxPryQrDxd6h3SavS3O3AaKUIW/FCAul2dJZEIgscGR9Rf8T
6UH4zTolprlDi2W+XRx4OJ4A0Alt76xQDVy526GspPYUvxuXPKv7yMQFpuaSOCgZ
AQ1V96HMCEaEIwz9CpWMjPdEUtvXPfMcDCfw2xstGFQaoCbHrTyIZG45oL1YSJD9
8XJwkwE1qkqrwb13SUN9ix0AmZeEzYNN5+psFZ+n/VoNSCQ18dcyOj1RM0TaEP/J
1P2jnahUiU8ejNM7DhzUS79bJKCjp7D0ZmoTJUSgh/0zJ5ZnUmHigG+xzPyzRQ+o
gGhygtHMKSRaXGNgSw5sDa3BU1Rv38IetG3rBdLuE3OCydKguNToG5SB7Wp51Lqs
ibrekHbv+5xgS5+REO8sKgLVmb4Uoima14FRAsWyieZe01L8oMiYjH1U0H+3p9el
kE2I5YBYikGi87wqO6TJ6knH8IJqBAW0kvm5syy9AzTt3g36Fs3lF12mdPGRSThp
FPiH+L/nEqUm/XgjQ7plYP+1QkwqB7wWuDpGqI6b8YIXziRtqfm0JbtwJfYeHF4W
eYqnpYyKpwezuD+1Fpt8EjYqJnuGOKGOqm6FxtkuGGkpX40Th9lxjxA51scACm9g
1ucNfJiBbVbJVi08+4uECFwH9SySVN4cQLB3+a9FdS9nlpB15ssZCE9AbFSFKYHm
AgwkVk9wR5E1qFnk0ZQFW/WUTEHWNDVTOZomulANni/qCBIO/B/ts0SOH9FmV2O+
9MTwW6+0QQKQzVMChQ3mI1MDqppVZYrLzwPoZHrZJUbT7LIWcGdznSY8ad3iE0nc
LHdVDdwtN53lOSVO7asLKf3d4WdI9itQq6dvRXzkFw/1Xb8WVVrCzhIqvGW+BLMR
++kB53t5pn5xAkRND6iB+Pa6i+9eHNO5ceFmiw7yXO4AmUMLUfML21lheGhJS7vp
ZOGt/ELkE2P4P8hgAHa2GzP/9EwEB/vKsuZxKZvT2vkOTnFdTzcGa0RREXYLzzdi
yYduEVQo88lJnyPjAonc+CRgiyKZSefzAGfhRmhLHuR05svHEvnbXGUPx6xKLnx6
zmhIqvWGCgNcqyC5HmqejKc59ttudML+IVy9tYvyxuslU8rML1f8bofNS+n7TpN3
xvBJKUiDX5Nmh8Ouf9GXn2ndqYXOf2s26VihDBEJWN3wvRrZ+0OpL0bgmSNxgQMD
PbatzCQ7mVF+CJflupJGtPp8T5gASTlNKwloCMHfDV5qBfH6824mJeHl44XlVWh/
l93cax0DZT6ulnz3kzJh0aP9lcFW9chX+xLQrgiYpFudM1x2yF+JIvKLOVRHBj6v
yDQcudr0J4qz4HVq8FJObtyJ0RIKgxoaoWvoUGV02KhaNabpfyy8bJz8WVpu3AbH
rwWSN2g6k0uD/Zcfr/Hv38N61hlsrHJUsB08Yhn6tEPlSlgfJT9WSMMueI7sUbeR
j3KLENf0JK+TEuJAcpScYK4A3Fk8ZOBquo17dfcBxm/qOnuXChDHTEnK/0iC1280
tL+qywUBWAwEgtSN4XzeWNmzJU1rptYExFlPp4x1tdEhTQp+vYwLWkNZctutDfNb
KvcpAUIbenKD6lqsrUkCyzAVnX2skvIY3D/IMtEviFezct0UBK6jpAvq5bosIyEH
TPtJ1aXaqff9kflHr9DY97lmKdz8SkJx5wWoL0SDo71QnKDFFsr+3M1w1NQdx32h
Eq+du+GPpPW5xztE98nUKdiA16VNZQTTKlgTnGou8CIwM0HSK4J+MpZvxbpMS2J7
c/B+cdQtbfrNUZTxVg5/1MTuhI5jrj22YZQh6Vd8GReWQFVvBsgdyylP6D6T7gws
k2xsWBh2zB2dPKA4qGeuCkqN1lMnRNeDn50rbkjFybgpPNJy1gUpQ2kebiIxT8aM
TQrDKC9+5jzI5rXwajXdXzaC8VZNmIua5pYlyvQXHDrwobs5UkRqMdCURmB1OUnY
zGDcNzWrI5KowXG67FvUUNRAlZPmcN1dIkTnQxwRSinVVQbuuxzL8QH9LEw+2/Eh
0G9ip5C4YU5qG/jZCVfmySuY32cJpst1JG2LX7OObQ5TSR8CQidSQ0eXQ+ezqvzX
WfAVhyM2kCbhPyvyBdDE/LkN1rdwgjMBjCK7cAVfvor3ebuWpujj/1DnIMv03qV6
WAOARQYYDA5uSHzDgdHbPafMZQJh6sdji/Vfzt3Z1p7DCUnyRO4NWDGzsLEGSLZ8
47lOSDFz7Nptn/ERBqnWink7kAc8/1+7Ca7dJsyQFXBURKWV9Dw10SyMXysp/P+/
fT3GWugjwtTAzwg2Wp7D3uRiZG/XGAeSyCSHeqfQeJiM7SKXGBmopX29YAjTe914
7yK0fF8Uc21x9p+1na7iX/F6bhPrz5T4uhblGbLeD4EtkFlnPbCahcoZfHIg6zc9
yf9w/enYQJfxX8zeBWfygN42iqHh1O4LR7za/xxrodfP1j4hPNtF7/tFuxw7Wobi
cCq3QtqB+U3lkBxDAHHQhvrpVJYt/MV0hWKQ8F0idmJ11zJy3WO5egPiRG3ZpWMk
Ub+lqDDY5CtrJmA8PY5cEi3WIUz5d4PmirRIwE+Mr18FFIxCg0kuyieKlLnL4y0Z
G00Xvw7u2Ze7uFhdLSRVirRdnjko4bhDYQxNattwCgXHuxMO0sKm4UJ/M31OReEk
tL70EzG2O4IqfuETSa43k1EVe5mL0M1FeOWFzHQu1VE8ijm2uzTrVQb83iI0DSEi
sZMpVNR1DJoeUash0O9Cy8WeW7fa0Qrz5V0CX1sVydieDoxXzUtOWmXVftD2CAJ2
SUZnGDphOOwjO0zVJK+JJHJ10Izw4YsI36/vccXdnSFju7XrXcbGE26IEMduOtyJ
r/lUMgOPFIo+pW3bdMuFCg97Yr5r/Cobb8sxT50uKULU+DfjwKQmNMaGVupEGTpC
ssKRnoVyUzDz4qRHGvLhcwSxb5dTzoYQ+NRoUKPDGS+IksTCytNsmw76AfrhPT1M
clWqKx+EUkvkTUGBAiLq5AbwmzoZEBF5k7sxqQRPfDa84QILUzoYMrgOezYm65N0
aat/0eajuvSO4HeD31Ij/bE6LU6Ml6t5mh4lH1OesfaQIGxcXoFYgiXrMvUyJDX/
vX1yBOCOHIwspPaB0Kj2VAYFRqC0ggUr23Kpuc/50aGrrDw0FWpOJMUVoQLkfEW7
AgMxhdiYRR/Pj/vx8W+zceHvdWupQDd+oRhe0VskObMHUohZ1EVnuMb8julu4lR3
NoA7bIKlSRViUiHs5oOGzcSnG3uCayhdW1kD4bzyQD8by7rai60j+2i5x8LEwGtF
t3HrEgm5qM0yOdkBZxSEpvDzKf1tqQLVSx+x44Q3r1EIKpAoQtGUlDlw44PJWlPg
kNF9ojjzB90IgGlSDZcO7XaQ3kV8kEHba+uid5BfQ07cm1Nplni3eOJe4j34jxUq
FpZBb1dqIMnz71uXE9QaiKiMtbSb1p7YlzNklI2SFrV9x5q2qBiKwgA8O1sA2ugL
X4sZfqgChYyj/q6ioRbLizlo9/XOq6DXTDpdhCgZZR27/o+LjuHn2r3rqrHnnJp9
n7HCsQHGOJ4uBmUNFvz8cw8RvjCtKxGd+k5zT/6jwRIZwcERe7eExV3P8q/jO4Wc
u05egz5RODhCIYtunTpJFUhHh1J6UKAm0sxPTg3g7z5teTqgBt6JVd9ZfNmP0bCn
iamyHyVteI40jS6K3dyKT7fdJuDHincrCjhz4j/WWpFuUVBqdvSNGPahNJHjxvv+
fMUfQxeLlB9eyVK069RIS0pE19bmQe8+N+L8lHAP7n4liwfxEkKczEzVb1CkgZq1
JiMoFIg+xN5apJdt7obw9fP2uUra/wTp+/H9rqjp9NG81AYLIT2/jkb6wiwXhOqA
TgYEGKTkjozGK+vUMpg2xFHDOaPf1FGRHhFSXo2M2b27EpLaCm16xBRL9XpmeH8o
tEyTM0iieivqzW+kOljDcMPyvv9Gc4uvDvh+ZG0dYc2lIW4srsLjryKSpHGOMvlw
S5E7b5Ag5RO8t5BgMga3Cm6vh3IqqEe/ut1cI0ZFwZZKUdC3XDskMrPpTYp/aG/R
vnaqs8WzvThThRIBofe2aXA5RsvNB2Lktx/B9TeioSLDOZv/Ta+VCGLoD/RAvxel
r1dv4LBVsoIalrvJhs6+oTHhJtn6DhWiT+AvHqX19Mct8p4dkwCnY9EYjUguq4U4
AB9arh7G5fS9vhyKyZOmzoFG4YK6BibW//qZfbS26ohihf2olD/C7pMszvaBPbVh
H1X/Dm5PdOk7EBplJi3yBekVCtV5EXLbc8DVcg0AKY5ie2+ewMNcFckgHpZoxGni
hpoAOy+Uhz/Y/H8MJFa5Y/A7G7JBZbibxYBZBDHFVrKMlgpI3drLDXzXuyvJ9Ovb
7r+yDtJ4/1sX6dEz74zKj0KESf6y6MHEsMxFIw25mM9BOnZUirQ7TeBZPI28dS/M
s2j2gSe2wv8faNSI7BImFXoPL/9pnHeOiYRtVK/2Y1BXM1Vbcx/dr9gvvSwOjrfe
ggT3bpgIZKAiibLn9LbKJCrP1WXJoeIZrJdX3pBx1V3uNY7wuR40ZSIlphY+yUQu
VJyZy3nbP9v/M5MFpW2bW8PlH7CF3xIzF159ekydwhnU2NJsrPsk/k0kGmpZ5bv+
yO0XcNEfX4oxwOith7nTXmybWCBgnksZVaM65ySoABlSbBlD0l/SGilhEbDAbU/e
mwUDOrdELmFLNb9mcjuXhnH9uT8H3lT2V3+84eWtbP2oHLbRIwOCOFulbUgcWz8S
zd8Pmcur1j0hFwg+zd+o/jTiB1pFMTwDOzAxTpqgXCcsMAB6MqhV5HubYiZ04VMa
Kv+1UkG7mSIbJHiZPxBqHtzUGD1XDOFSsd54fZl42DtcZ9DZ1zMzcyfZjxjgaMxF
R/GwyOAopTncJKdwvH64QwFlQ8OOEvfNXhX03WX0+T248ZlwDehUiKvXqtXH+0lQ
R7Ym0a6HoAqi/m14/C9ZNjSollNWvj/QhxB9P12Z+KHFhqQVtmwP7UfjnCmd0j/e
15tC7xNNs9AipCMK6XJxHULX1S7owasi8b7F1H85nOp0HW1zQu6UXPqO98T/46Ub
yj0F6uAdIznWFF0/yEoc1Hd5WGJ72ySqqJqtyOnaWdwWZXP3jgxaq+P0M3oz3hzT
9eDT5A1y5E77J0SfEooHu2EpJHgSiWTgumVb42PZVOh6bv58p+KdoD7aUDOJyHbQ
V4iXEH+GSLr9HZKrgw7eYS1PTMmX0Ty4d3cwI5KTyQ+eauXtTjB3gLSsuiE3eJ75
7Hj7O5rfjgOtb618PBAB0eXikZeXSyEASky2krybWHw7JDR38JYoSeJKglJ+c9BK
Ryu6FdUVsjzvyotJgbHPYoyLJbG2/Bpx9H63BpoWPzYbWtJBryxubqLqrgt2jwCL
/q33D1dmIsJjG9ivKUk8z6GWlLQc2JhjbAuQxQkAMNSbvpblkRgSupMD0HfoL1lx
anRCjar5a5ZxQfNEyve5r2Fkep0GXZhLY4cIydUuRDGxbh6i0u7IKD+oZt6cxI94
GDAZXfZ1eV+7yVBkrzaE0zbxpdNd6QL/1+pMTVcHoQKbxYkJoXAZisP9BP7uEKpq
jer4Vs1KBQIGKdoJI5LC8/IWqw84NZvtRtYuSYX7PTsmhqI2vB8hvJSxN6KRas+4
VU0uvspCK+TpCsdJ6R0ugdwUgubkDdFho7ChlbuQuOJlXVBrcZQePlPltdc8eNhg
BaQ6iN9jYTQg2SbfBUO7eEhbBqZGUUqN2Kzj0h7NF3X0W7WQBSey8yMkdN9RRsMY
grvLHnQnPChmg0WHlwddAigx4zfJiLNbTPT4mTmko6VwBBY7YBG4Mi4jjmQlrm3w
QmxcOO1+7cpToxOrvGQvYg0ka/9ZZ4O5T5KkNv2dw6A0EjGxeXDk5p2w9AEMFpSt
ygH4ltPRfEv8CyKzzjF/KellyjIzWi9tZMzKIrHko0l2h20pyktxdw9UhCglaZQG
rnctxEK4n2egtiXTLg3/ieXNwFjpYcF//wPuJSO07+JoGdbL4cW2cgEeCac3LFNg
kvor0QjKY/4xjMvRhzSOj4knXefkRHoYMgDwpRis3QeeeA++jVe4MneoZ3vpajOO
jDVL4Ani3d2CAoiY0FH5djVpucZn23eahZe98WGE+FYaf2SwXGmMVUMcMBcIwCL6
q94bqHFyjMKj6qUip+J94q2iA6wY1M210Rngf8Ou5qSn5A/lpip/ZtM0DsjgtifC
GUiSKFfjSGVj0dSps8+RJ7f7pI5h4zlpt8oTv5KdSBUx41rNnkQ7PLl00MaQ40rj
jc5+/KBzmBLI5+5+D84KQv0Y10/ouzA4KX9zEFpovtgNRDdBZZETfCqAbZ3bxsIf
TWe9WyOzrvD0hF+vUYz+NQ/hwUI7AeIy9XwBCF7mWsIHwnlp87jTh1wze6mFKci7
1PbhH9onY5oo5amV/Of9PP+QclHUUu6HEaJLjQfx0eTFt2/42Keb7B91HCDvuR/G
7UJFFRo8MVAlcMjxOKvJx5t4pv+Bg/4V5sDJA5mSiOj9oIAvIdRZ/oiwn6483umZ
aDIq2hY7JPlllrhRF+uh805E1EWqwMRS4DgSNwDo8/NR/e/ufQ12db/h3KhWKW23
ZH5FtUmJwymVfouAYr6lo1nqY+Z9Qqk1EJhlNTDaHj2CUNC+0kEUdE0kfKyjkcwb
gcnPBp+UH5gyRVFcJ6w9CvzM9I0HmTSVkqvr6b/vCdKzMdpt3EBatGyx38KwJ9uN
EzT9bjEaQCLaHUQBF7oX1V5rpNiQF43KKLFU+gYPei1rO0eJkNGvidgsAR7CsWpJ
abnjNt93Y8+dD39IfnJTtfZ5QZOIeCavLQ437aJh+raMT79Mihb/iGslpmQ8vaD/
5y8MZA2OiBuz9mMtRAidAnFKOmJDSMsiDMp6cMOHRz+AzR5ulYdl1iYDJSdzuvBt
U9h3yjAadiTCL9iS4xYphKWq+VQU5MchOmgQhpYx3S77a/aGk0K4L9Aq5wD5gyeI
VecDDNHHdV53+Ps0L8fLq3GKVvDm6u7bt8tDrUY46TMGcdRFcdXXGwNZ2Q3aXdaO
3Y7ig/bffgUpbLpef+9Q1+R20FR3XJzOIcWY+yN5rBfQCdBxfSMTmvq+mqscFs5Z
Ht9+khml9lIO8vvRMcHfzhR+ufUTOcU2HIoQBIu5Lp6lOWfJud0pMSXm8LdkFoIZ
cD5DBwdSTBnZiYmbsWxQ1aOYZhcrO5EM0FbQUbX9A/aBAk8dbmIA8bO8FZ1qywNJ
F4J7Qk1JQuFMZDEC6x+n0QbXhy5iX5ZdGXGSNw3/+AxKP6Bzih6Jh90XmAbswQzj
9qslQfXCf1QbDy2ITE8jBWlFO9mjS1Jde4vraub4KmFpY9C6RVFMMPP8h7l+dcqT
CHRIR4VpQ4pROHp+QV94rkKxrL0VEl52HuVSmeLWrFx3dkCXHYdJs5oyOXdxkUl9
2y+x56EAjXG6ElY4bu9nwvGLD/HKjsTdoHXyI0yBWMEiVcnR5pqK1YlVWm5qI7+e
SJeAFQaNkW1cVObDMfzHaprIm9qaWWqJdvDz806qDXSeJNNuFUhw0Y26vcwl7c8b
iuqM2YsUEI4OJMZylIm5X8zGpEv56YByCejy86O9K0tEoIkXhQdLH475DW9nSki9
qusoapvKLJOVUwiqB+cGnRR0XIhrJA7xHeUY+1VMK7bbli3MBlKjl3RocyEYdoX7
lNuSwajzBA9An4AaogT/Ibtqmhd5gar8l9zNFrbuqkw6kuJi0M3NiOYgdrt984IH
409cnKvEgrCM0+5RbKJnZYoqOIbOeIUitgSv7hA5gBp9Wy0JLV732r+TmvtK3NA/
dywPbj00JVqgBDBQhDgnRcBM3gVmTr4bWd7KuA3C/2gKM6ISln8k9IbMgJCkzNtE
gG1oJaP2loB4BkhycjWk0lDTfYruwQ3Wo/IkOlARa5f3u9hmjSdQByV04oA3ApCR
6mHndxc6zRYiyU5KJswyas+QSG0OPTjK3PAf4SLOXyuq8UvkzoRKuW5y/V4zZ7Dz
9w+NjYwDOMdkW0+M80btVbxIHBJCerwk0QRBVpmpZYriaqnEYuN97BOfPa2jjHv1
4AfF1hKgmnE8KIxOpb59GRJFCJIsK6M0JRGebFu26hMP0WIQu31uOaOGauSfYZk/
C6yoaVyFFmh8uO7u7ur5xJ4eRLVspvRHTYwJtgfwk7v8kCJ7Z6eTVsLd1kwYLoaP
QtG6uipnreJxCX69edG+0eX876+XBhSWhTQSbB3q7usWQK3meun1VHj7N2P/+BLQ
9p+VvXJVoBR3lYZoEyED1C+lAdtKsYMtH7LquAvgMaUTZINPZOrkkI+cQj4gSFU8
vvRUXxZX5ew8HsmlV5v4MiOa/1+CcaD5qb7nVnqFRSeisfGUtc+mwgidKLgPQE7x
HuijGBFVw7T/tWb6J9Mueflu4I1+qQiKgCUAfGXbRJxoTAw6PrJa0wJHYi7mdfI9
QcqTr5k7nQ6t7avuxY2roCWs/9UPgTR3hbXqNQmrJGI9TpWHI88hORfkR4ALgIEE
810FgY8ywvxldntwEVp7i+ee+u/g1kHRFtt29ef3fwXdzzvshIzcqlCJ4GL6LD5k
nkyrxG/075VR5VZ2FtPxnJ6mrjEaep1eumiXSRs1cRX4v9rywkmpY8O8sh9qBDpI
nDVpW+6EA5lRw5kNEnrsaDu1c8jDF7qXFPm94AFMCEVw5fcwOakIoRmsQHkc1ZrO
hSy6kxQIDYQszuRovz3XvaR6ofqlTSWNEmJktmcqWGd6X4pbVaRkw9AaeAteVrBZ
z40u0VRdTbIjKuZQBEeBE4Mh5yOevVEVmYrjUAIJDGYNg1Lj1hKM1CYMTNBwzBVZ
GMx9c0YJXDh/NGC9SW+0hxPyNLFdov4qS8XDe8MXL/CH4VN87ea5Ml6qMqsB9YX2
zgZUYtFm6+1HWk1HKx9FaJ3jKtNv7ytMU6LGv+BHXL7a4WCbLGcib66TsDysnb6A
zXEIJ6ITo32BnPhtjAERZrnrzBE8LsJLLoFKr0M9uAn/vJ4ysXYnGKOjyvdc98rP
DgmLplod2mcgQukOaWYqyzl/77E/g0t6MPKPuaGpoiShU8UA55Op4CKpKXpaUHn8
2r637cbyE3gF/SvZbN2zwHL3plTiI2FjzxuyUaUIAcpKpzdNTfMmstZpDx0I0WYa
BwzNPL/6MlYP58/9MuGVNLKXigdLcKZLJVP5zzUz7vG9/Da0AY0tIQrVhy8ek4bF
QgQWMom7BUBQQ0SC/ADPvl2i0qXBi/U3fqh0fL8H4GazXsS3z8dTIFhVlbDjG0TI
sbDvplKzYWaDpLJ36/yZdYJPhZDLRIBa8JJrSbGR23cFdphKLEW/HB4PDWvyPtQX
i2mTUDAEji8E4mU+vv0KGg0XOWAs2cy/c9bl4opBKfP8g+OYMYygReLrl976h1CY
1GOSaOWQcBEAo6JaUb0K/dEA3lplocELAk7/kLUs51pIih0QgCa/HN19zTIp01T7
gnnQvXnb3GCsj0EE6NUDxkASzNBMLgCl4nyCAwHo/oC9ciCFS9ACNHaANRn0fwgh
TGM+Aipy7AwpHzulKT3AekdVLj0tCQcGDK3MyK8+p3MgEQsCY+3iZzPVUlm5KSXh
gLsvvJRnmD+rmu1BU0jhAL44/QeVmgQIjwvty6F9gafZMTzNmwC6uv9/pCiepIAx
zmf6yD37q3uj7IDRXtoVn5fPjpQim6oi37afmV9yOweGMknV61nXMsjyj0CbXzNH
qKUgxM9nNsAKERYGffWt3OMZ3BzLLgASW5lre4lc4lDgFPx6kJm2nmy4CCAackQv
DXgEwmFLsGHn2zxlU8jyXFI5pndbIBXNKTpLrtekFAiNJayCvRD+izA4MMLKpR9a
FB5tnMlsN+AvbSBc7KTZ+XsE3+C65Sk+KcpB2obnzVN8KLwu/H/QVmJxlBqnK7/u
zoRxcgg78NS46aOf6qDfaLstbHWOtdlYlhXOR3wANNImf1xHnxIM3lKseY4I3CBj
2Z1+L8G6AvD6goN0lVHP6CbnaasP7CivvBej99A/Cf7/899LJv1/izdrFq3M/QFI
dOKmggcjvAAEoqnyyVoeXfT7+awjOo9plO0XW94zrW8qeCky4y3NyOiq+Dm0MJW7
BBg24MVS89pH1OEbVjfTkCdMwG6n96xPkb79+8hZxNFtYZ0W9GEAzn8w+YYjDRS8
oQAhKAK7jbJZiD6EjzPqlbPLoFF7mkGp+NPi0P9MT2g3AbyIsZBLWkwt/PlJ8mrz
sascwtp6BPIB1R6STR5y+Me6lW0NuiNFmki6n2axO2SZM2zhag1wmPYgM93DK5j2
zGRep4IlQIF962rNLwewowJqcEg2VPDxwYyPDPpQY9+U8xrvljCuOmDu/WRNCmWD
XqtS6Sb0mEoajH2izm0HXFnQGxDEH2vsQ8MJpSyDcymfQ0ad3E6N6SvfDqnaWd8/
nSKZsWfkj5qNMjnxB43rYHNDjtPzr9QIsXuukSTgbvwHgVdJo+UEwIYiWY3/WCz9
VjiEksfjr6Q8WghhOLpatyLkXsM4Cmp/GOiHz+QanS92jtOdTSJ4fMP29RU8ahe5
dEpnwcvZPBWDAHhezOguDS7HTurQ959HcpTYb+C+kHNmwApg4fJ/yWZhhxySuxhu
bJ8xrwoYmwrPQAHmARDaYAfSUD37iXK8UDyJvCWewXvJGzIy+Pl3maqAip5nMmBi
ORYbSs26ZZ7hE2HcRSgF9Cy98gxewa1e2stkNy1eXC81SN1nUbMLhA8Yc25cvWhI
JqHw+y87dVKy6LOXX5kKvrZgjumigHsKjUixtlwB63QOtWKOF2nzYYGj8jbvIR1m
B6tdMhk4thJ6DV2hXFep9R5Qfl5ONEtjWH+TUdKsyDh4TSYL6wrZt7e5Dij5ivaN
/13kEwxmoQh/l5bhO+vXQfV2f6L/IhxiJBNuSvvzxmlLJff+2C3ssVcJUQefwIiM
Qju/NyYOZY4V+wd8YeaI3CbiJiOzCVDy3h32sOJGNkPOwhpsRiSqLlzhQSChLNTS
eMh3op1yG1uZNxnpxk4Ll8WhgKp8XxGUKejXeWwmYBaXS8RqI2xGRS1I5z//TOgr
X8K2KDMw7iAWLyE3w5wO2DPElq1DgTLsS711X7Jhw2LArT75T/qSxpUn6LSjPN/f
RKlIJ3mRhUhcjte7yKsvNwLLnEjaukwj4ZY/hmhc+o8dzDX6iHwPl1v7cdBs9+Uv
eShdGF42ofojgEvjuIAN9WCPOnNVqdFOxnJlT5TVulfbfW00V1oQXZQnEj6jflOs
ill3vgX3NB13r7deuOoIgYzqzcwXEnHzdHfkZHnp/SyRl0meBQRD7CGzZi2FheM2
5deUARFdK32EnLs/Uvbj1073RxFETzGdYUT+mEuf6kW3MysHQkkq9uE2U256veiK
O9wswi+i+MSvu7T+E1jXLCzYk8AQR6h2U1SfI01LvMcQouVtfXXfSli+Br7vI2AS
tBuMVau5SGpD9TjwvPAaX2dTq2mTf5ntSW+hYF3+GYcMWf6ux8qTKe5aX5JDZkWz
ktN7QxIf8hwz+dttK4Md4Nz1p/ZsbVFD1tTKRxzKYXdqdiNx/Kske//QXL/dPGWp
gIR7YmgM1cjd3yVvjbvJd2UzuupMsNAh58kRVJqJX1/LGTDaa+g68CJ6gzOetRDt
PN8BH3mwZpDGjHBPTHbKPYpQd2APQm/kBihqSAPI4BHwtOe2wKMWr12l4O+ELFFS
a3/YIObGW58K8vmzcnSfL3oynrs2WkPCuQlUcwHtEKq5X1sNiEoMkCC+hVwZ8Aum
mVzMCT9JBjHFbC9B58DyjT2gG7v3FI50E/ISG8e+rx02ZNWMxgbuGTk7d20CevVC
TQyhRAv6/kuQ30vIoEu7kjXAAA9OMOY5jhM4ybz9AF8Wnz0VwKOvd0x0J6ZPNCtD
RjEvGoiOgGSmm/ko0hhnPMTVHyktYBfKFyOGUhL+yKBKaC3rFarvzfMqHwny0PTU
9Y7MvNQLmVLD/7r6hl81zoeFU4Io2TIx/LcLss/G2XAC8/v8S9NC95REwXyKi3rU
jOZ/uiI3CozlG2DvVTb2Dy2D6Gg0ymShsseIS7rfS2ERe3PnhPAQOrXHfNOJ1IVJ
1yoRs/W/MpNvfbZAHlRWWvKPv/PUhByzv9NUZl/9unVEXTm3CpUynjXoIIROJLmk
mfL6uHXvP+4WQNdH+9mDDJamh3XshST/bhr1vmswzr8Y5eWWh8f3yB3MIxGwWzn/
jW0qFafFR8+i9gW58Xk7rKyDRNI73Go2PnBaxmKgX0EBzos2XkYmtljLMAY7PnEO
I7S8f8T1gDVNQFAgRmu947kX5Ko6IpYJqAaQdc3t9Wv7TI//epBhACwQNjGTnged
Ah8DR7fIMbymvA6CFOkb66r15KU4e+8YuX8un/E0SZVo7Kf90yRsZsL4EvsIDK/t
q1+knpbHBntLRlsajmd1Ga4w4oTkVFGauHMkQwU5spoZgiIk12/InL5Z0yfMov3E
uu5hUhat9ydtC+K1Vy9pmva6hDaLsRle9aBufOPpcygiJZhoLf8vLe8qIpWau+7t
hLkmq52qEzB0l3H418kDmyK8y5hVVkvSOCDw7paBgsl1zpqJHtkyGZCc5W50icyo
E5noxB9f436h0HeWnJd1OkcRrxhyNDH4W0V/3ZpkOFqFoR8v5m264vROWnC1IIhy
MkmCapxXQalxQq1+5DMT2b1rzCUL50sc40EcWsX4Ktx+EPaJrYBd4FfqMwFSTYD6
mJzC4RJQdA+N4Ax/j9I9N4VX2QiqC4jkuaGLXot4+Lo9l119p9O8nbHPSSe0VhF4
rguE9dd+hbAsPa8b9uwwGru4Mk5dYK7sjcvs5GX/3hrhgaYhtSISUCJpflzsCtri
lOteMPhOmBuzPNDEt+eVtRgGosEs1DGGZlThKtqiIxVjr7liTRkUu/G9cJfa3kTa
PY5OeBusnH2PmKoD8wzq2Nvv+INuX5skqg+Wo5yGuuhVCQM5FbwXpqXjqVhUrfaB
ygdnED/HzMLPNUURCDBSPpqXCWfHbw+I3bRKd/qgmEcJGiqQEA6jPfVIBEN1YFC3
RfqJZzr2Rw37MP+U3G8pfctnU01E/hGtAL9X9AA2eGypH/njQP+Xr8qRsPBxVTH4
G4HK0Y27jQeuAMpJniG4Uih0nh7Pd+5afVoc6FC7FOsrbKnlkZHrVYCl3wvjF8pG
k4tCGj6J5Bcv4nbhTS+HT3sc3ILrW4o47PZ4p+2334Kf6vtR0ofp8tFqGQ13AkzO
QBsISGUf/PWoevXm/fbECGBb3dMY15KpdehRsPjSXukasLFoCM9b0p+/e8ummOYW
4R0HSZuBEMuO05+H1g5tGv1HH2kFoJZD6AKxia4Bxj4RMUmqKTxWRieRzH/+KKW6
kUSGAaMt1S1TWPw9s5abLDH1fb6wOuFHJg17uH3wGslztgjLw4ShLtVQ3X3E6xoz
yJRyMrfgr56LLDIjMhZpVXf1dOTNZWZkowd9jwxjhnoqX8QRO5qrKAySdyCY1VbP
cjqCwo/9g6hWt0uLN4lYroSjwxS4OGz20E7GhcA5o147W7FioacEg0A++hptwwF/
CktOVufxy1QoDx1rAYxj5gDJQCtgs8tdDUZXa88KJ9SlkjdGnft/JCxEHTSTYXjB
vO7e4ThE0FLr0y8JMxImFD1ZSI1shmAmZhVruVp8HrtZVYz/bACWSg4ZThflvp5T
7lDRBwaw6sCIRBgzmDBYwNc3dY+sbOgmmZQK5usOzzSDlqyHVmg3V4udtuxL0nV7
a7VpotpegDEv94n4pLCyKU9Vj1i5AkL0zivhrXjFKswQNymxJdz8LKPd4AoKiWBP
ROlieDYfS/holUjXzr1GgMDAZeRggxgiQcvyya3S52hNC/bDgwumLhDMXbx13ftI
5fEMpKM7Cpi9wyJKpk4PSpbufEDaNZrEX1//KmpDy4tGW1y4qUFRnASvuidjkP8B
KtfQa8yEjYBAQvDYrxEn1cWNVJkv4qbVe2n49jproi1lRqy73wKoKDn2fRXYlpTS
EamZIBMEAbSfj3u6JlDU8quHlIW7uMO1QFbWqly76vU0Q/chhljdQFo9VnAXNv69
XfTlFyXr8Cskim7e4RbqXBFr6MyIggyP1HiMGlWFcl4fTzX4l42ncwPHZpIapUKq
kunI+hTXBTzc4C8eoPsd6JDbGvM1pPj6ypkk/zWT9XHN+q5+LfrFPuYYMPrHHMX8
aD/0nNb/zNLPXhbUfKhM/9PyrtrhESDKQ2G+lqvslRElWp67w0jyc08kCdI4V3aI
W8W+OoqeFEgRp1hBUUUuWUt8lN0MN3Wsy9i5jUyE9wn/Vtrc5722apCGydje1ohK
Q7x8eFjMlcHQ/M3QRMStqW21IxOiM9t8GGj+7ddQXuQ9949by4ROjTQdiKKECy1s
rwibWXEsHlUXJd+huEXcVnMXmV85qogv/573UB/tvgcz40gbELXjYtWhTHvajvNR
j2MJyVi7uvSJ4y6TYzCDVmpUyxTKzeqHgvCUb91UaXTLAsXrP1w4M+xocz72H5Zm
U8S8JPuc0ffJ6BcFTp0H4Sfi/IQCNJDckSVOiBCqLLSmaUWnenWnTzXWBhDGl8qf
v6PVf4faCq6pADxWzUgY7aeqMjQH2xPgh+PPC/P/rMr087MHFnV/DzpnQz6GvPLF
nHlQmNwpJZPF41QlgU7WpauAno+7aP2N8Fb9Qq/DBioY1J+FeDDqKyNIUi2y3X9F
K7grSegqekOuh7cI0SEe1OGMWOGA9vQM+IotRZFPPoVgkiP5s5fcSYrpaku/aNSQ
ifdn6ayJFFQZoWbP/yj7DINMMS5BJYp6MXk9R7moY0yYNcIZ7zDofvXQa/N1eK8v
faXDQmLpkmOEetbLRuzB6jfp2o8+s5al8l5bIbbkw8sk2sXmmP2sv9vwz/899tVD
m35Om1ZmtsUxdYoy1rqvCciIgcq8EK9Hgj8Fv9dDOECxgTrAZGDLIwDoTiW3V5WY
Xkb67U2EjxCz5x3b2+tuitw38cQLN0qqCMvEm2FNM1fn3zsE3Qqs4X1/F+16fbND
xIY89nDEZdaWECT1jrovzvkbW+8RFyQVUYN0dowhrQfe6Fv55PjVuDAFMtzDlW/l
7MVHLXInehVk0mHuA64nnrrSN7ttvp/s7dsScK/fkcD/6I6EuXz5h+UMdWd9Q2eC
e755Jw9NrVlVC5Rdx9xmwiLBrKHGKWBi/+Hk8jQBuhsY0WQfhrlTVtkFVoQ44OeJ
ngXvLqPlS3OiCvbYH2zXEzwHgsBFT2yyUR5G1j22Nay8EKz9kRX6jdgpLU8Pbg/J
hZA5rPOABA5K+QZi0h/WkLAhdAUIEPrqLqRS+3jZeNuBQJv9r04tZEjB7XMeKrXp
e1neF+JbCYyjJ53Y4DLN+bsU8FumZGKbRKHcC2VHG3+MvwA0LJx6iXbqFvjSAExm
zqy6l/06YN9wrqHCvsfK56AeEy7F8KoaQt+z0Ldbxc19V6jNBM5PNF2s0EzjdxU4
T6IpCS+t+r6NCxTe0COd0GW25FwKDvRKqWtjwLhonLjPd0xHJ6XD7yzKTY6IfHK8
SJm4IGfpJ88k2SNh96Rz6hzFM5HGek3szS/iEucAImks8Z5p1Rj0m4cbMyMvkTkB
kkDvZKqWPMg8664uAaKKvo9c0dInRVpqlkdv/M0hm5po1YOs5MFF01xV96aL1EBa
uaYBLVxLslAJdbXEbwd4eQ5snp27a/wOi758WeHkCYB5TYa6GA35X88SWOcSz+5A
X7m5PFsDhlsNs3sAQTnl+8/ZCIFhjxZhIPEJjMjbudJC1tq6fp1pekdf9y2FqWZF
1G6n/AKJq74qTvCVHcmsiBKQBAnmxHXsq+tWagmBnDhGVYxfmzZJA6ZGKo6D/Zmv
rWOto5XjxYMwhUiSFvWw8P2s8f0KiSBWuk0dNIL6W7gOPrHWGEXNipSbCGm+4Jmp
jV5MAex9XZJHpEYsXci4VXlT2o0r14nbC+V98Ii0A0+poQrHIwdfF0WIPN3Zn3mQ
SN2S/5GJLXxwiVhVZEmTPKFjovDj4R7hN/mWT66WhvXqLWOXRkjXma3XN2rpLJPK
2E8PuTm5m1cji0/NGo3z0zEyktdZbrRIMSG5MoIPNquArK4mNMp6U/ASnBflfGUy
V7IpNAm09DBsYelSBTGg2lCVWtFZ8xsVw/YiYMJhZK0+FYta+qwGgGw87tUhUC5M
sFElZ+GEbO+GeoWd/TfUaBF0GrVS4VRz7H2YO6xAK1CQhb7X6m6GWiQwn2zsid94
PVKROC6u83QS+ShiZDgvl9SoK541+bcJJoMircKSmWC4bA2X3KMb5P42z7r8GqA0
ioTXY3TyIo28JuTdTbZJybpglWei5QtidMV1uDUVUzAWCMtuZZia+Au22QNgO36+
bsuwz2dGPR8t8h8yDjcxKGl2DHgtrXEdDJM/p11e5sWwGjzlh/c+YAhze7QRvZ5q
WIenM7+TMF4nIFXU1yD/Ig6EtQCFT4XrHT0+oYTwEVrn/66RPYK4tG5//BVNNe5n
PagKCSolNCYOjzOwqGL+X8zfWuvE254cdZg3vJxjSUenRFyL6rkxFt7DyeWUeXEp
pPRbdAfY/KuphPasQdls7NwE4lmjCpMo0u+0b6rwKlcbCb1Lml5nVPgw1JHTZMM8
1DG+CE8bmhhhMRp2tLHTQSraZyHS+j1fAHPC75FWI1yasjzyvsYaKN1DgqCG5ZYe
vpgz8AsV2GAG6H7IKRHP/wv0xYT5v7NjWk3RoLGkyh4BTBOlXjHrrKQa4Qfz+mkc
D9VKeb2fu71NzbWs0lILkFz9U0nalCKAk7xIZSmHefljTNbHqgnX8fEO6LV6dfKs
ajD/vX3NMZ66yx50a2fb9WtgV+lDJeH34+OuAAnDWNeb4Vn4pGgt0Ftnyq/7TGHd
Q6erB1rTEtvNGfKjmRjg/d6XPhpk3Yfp/lwjF+NcooHFYbvw3COzRm9Q5kuqHMDq
YmR/PUvuqr94AxQm4Be9ebe+NJxRvuusYzevCtt4/ds7OTyZCUaDAv2lt0c1i+64
Dfq/5RPbjHlNrkGs1BaQBgazNcHR5Sd0AAF6186t0CtPEiwID1f/eeqSsW89ollj
7u1nlLzEE/tmH0xrSLTc5z857GmV7w3Eyk+Exjqy+WmWk7vPCwy16+T23zWiKiZL
yef1zXN1Fxb3pcHMkw3R6hFworsDJ37AuCdCWl8RuWDu3pPYMk5T0JW/NjC3zFvS
SjXiqO2wORlcQdtsPZZKfwizXQsd8Rav5x7y4j5ILcLm4IsBzwEZp+OlzW504ZBl
bfbIFJcguqiXM11fEih1zcFPZuj1S0jk0DNZ7oOJxvsQQcO9PVxXeQ7eUcAk8f0k
q6h+9AumB9Safpt6voZYHERU7Bfwoor4ubynaKi9jdY8oztO42xs1cQk5tR5LjF7
v2Oy0/lqF8PcIciJIvDpasdvHzrrapufjcXw9Wmy+Ehf/fPdl4bZlj+E2Q+yde9H
GPwyBYUF//hLhWZm9ZQW92qBGrxu5elVRgDZQAX/EiO7JP6cdEQVjx5ci0U+URbi
i1Ebd4pkS/FPcSRPQwx+qk+gehv6ck63HIf+7IRq50n5QciRw1YYnLYO4eyBl26a
ijqulLDANjUnwVhHsOJ+jGfCZ79Fm6g3momqinYCZqr9Vc1HIGdLTy8N3C8Z4Hvn
cnJ6BMoqlSTN9JKgw5Cx+EXyf0bJFoMwSXuTieFBZMTY5AYiTmafSLHVERdYkWuL
yUmll9D10PEKpK3MbAIcAbiwY9piMzbnpJDMobAgmS9Oe1r4hWnrHVVSP+MtgTTE
2/6sCN1+t46tzOPZSZknOSmk0p/AiDLWq5Ua8hexfbDxzUmh1Y2XEmTBQt2OQ9IK
BY8IbnoW6R44m1yQXTmheMICl7c6ISGidpCe3a8nn0xHQC3k9p7BPLUnXIsqXPyd
ks8LW6IznGX001FUPrlhZJnaeC871gtmZ8/gCuuLcPvUDUOnqu6X3AcJzqgGJG5E
x5UCox/VbpLcHq6crwc0p8w++yvks66DlKWQSc+EnSSfHQtRaMvNxkSEkGI7l0Dp
0YPQucoGL7oFrIyeBFU7mKAsRZozgaOW9p20aFbTBzKJPgj7PWJkH2Y9+VwspTsH
xTIV5MrRpFNgcIuxhBhU5D5CsTTJR95eNc9sp14RzM0IqwSeexI23Ip7SnmSrHhp
dWjWJcSZGWf7G6L/HtcnJY1BtP14yXpHvrb8rcBpLN5CII4ogGr/2IBLh61/w9ed
+jiFJi5V911CsaQq11lYyJN1mQhdHZ43lgrDVlVCBN/L0OgjfnQh5AXYTu0vRlim
RdWa66mNf/r5WDSbPpDfbax9NjUdw+P9N+6xZqIQlQncJa1670TBEzDNhXtBJgZm
Ps2/zjbZUe2kUa46t6D8eWi2ojWvet7TLpIJvzTE9xtM5Qr1Ma1HmKZkCeyT2CIs
JEO5JAKYkp7tQSenTFrHkUYmZxZcJXVgMaNR4L1p9AOpXxwLKX13260rvsz97E0q
o08Gp7E3LYYhvNwXzgoTztGpYIJw2FIoFPQNFjPBSqw+rSkRNiDlYrfsy3bX0pzB
rqAW6vSBTYgFCyJPtc+qHOnE5c8ZUlF1sz8AGNLOj7AdBbQxv3eZnkcPtvQvVWdZ
hyr0FoYLrGXHw+ky/3dy6CIk8nnUlMhNl1lM58IjZbYC8obAQkGGhnpL+DHuv0c3
BIBFvgtD751Z9Kph/l6OYjHxw3ft9hch3SEt4p6itpoW2VkeLTD+MTCsZtr6g/iU
1+ReFVmpOY4rRIUOwM3hdw0/z49xnePvpCEzi/a2xrOYxvi2stvlyAzk9gBWK76q
he7gKApHPB5B6+zLEKyBAdGgmgP9fKiTycbdzEy9hcyj+mLwChjzymdAaStpHkhP
ag/cl9BbZc9RFRyPyeQZ+wiviXy9O6G4Acz4IkHuKWsvb9sIiSwjNDp8ol0BH7Jw
uc5PUxfASKmOYcHCFfFGcpH/EYrO5PqdN1udcwpWh9hPwxXHAsbFzkMdBg1Gblpk
DhtjVuT0UoPDBO4STVGhYmed2l6b7KMF9TN4bPxwO/Uy4nkUEG+ljLzNth8IrmAk
+51DQabXIkw4jQBCe0rAvFGZURcdNVJuoIu+om58V+el18kRS0zf1vu69GBLnvxp
9bl8WNLlJcU6NiwMAC1bnwiQ3SEcObM3Gc/eQEf2LQqXzFBvhRBk5vJtCEqeYFb+
I2Htq8H0xo7yZMoxM2CDms3CMeErA6Ew7innXJUnMVsOZ3XUojF3h54rG1eDJsYa
nt2XqsAd41SELdqV3u3vETc267LcZ6yXS1Eg1j6KdjICnRxUSnvtTDRW7Qz3UuxU
PftbkUOoQMFSMhlt3LOiIFrreRrPei4P8bAqieSOnaFEeKK6XMgDVPOzB3p3Vqg3
lCTfRBG8hFtqAHBgY/CZ0q4GkYnBDY3MWFip4HWvkjCYtdS4NysEiaITJKw8TMIR
e6ml35EWFmr0PlSNNmlo3V55N6iwIgOGJbn8FIRecRyIjuLv/C/XNEDcn4IGPulU
lDXdv3WdnMfhh+VfNJEI0mdhutO3fsIPgERQNycgCV9WTCyuNlaJpVRSELcmGoAK
Uf0JLQ/thH+ecPXKCpIr2nqLKcdV4Wc3/znRWWBvu+lWmVT8brYsjg0lRj/2TnvC
rZrH+BCbLfCHjjNwXd2okHBVQQxh8vxkfHENzM0nos24WvPeTDK1fWxGR8rQO9Ps
jUO9T+hsmsd8LXhRYVxEMSSTLIi9BDfZ8T3IcWvbFfgBO50m2LlZ2Bk2WIlAPpBl
Tk39Hiv2xdIf7qzY0btesuZU7RYiIwBTFe8bz9Rq0A9h7B/mv/6SNjvoZ4X3Thpe
U2unIoiN+1YEcSmm/Uo5GWvU8gyQ00qJ2R2EPFQWDiZ7qrrQpWEG+KVnov/uRAIU
wFxrS2RXj66kTJHF+imrL86O1ll2KYzHy+Icgl7snFgupa/ndW7dQen3W9XUUPvv
BER9DuKclHADM2CMeKsgDCPSvZfzlf2E6hTEQccuB0vmYfFWH+nIOglUBEseHlUZ
woiIHllf0fp4gHRR4YmrnBhyaotrARH3pnlvIieVkDcKRJa5i3oE2D9iNTGJOn2y
vNyKSIl2biZ9Q+PAAECDfuWZAFFZamjUIJD4MCqW41KxTuQ3e3nJK8mBnZ7kgDhD
Rf+DHaam6qPSAs7hvnz89YisQDRwiiPhL3E5O4zqNvVMaZhMfYW7bA94N3dOW050
IIbBROhCwZhvNOyOQsfLmoWmYcN0Sn0OUZHwSBWtHRpQ9w19KmX04iulCUA/PBHN
NfwTXkGPv1vbYSpBiXjnRwbx1DhVQPta+F5UMT4U24V14q0sBOfKutuHBqxRYdU3
4OyL+IZ6frnQ5tDnUQftJ9seNkeonllN5wo3QVLpaEFRSDIjQEbss7HfTAI4cBye
BpvZaF7fK2YKxBH4avaXRD5L1IYFlhHbNEkIFUPqc6S4dNyoZQ0UdLr2u2GaBEN2
6vntYO4J0v7ZPZBZy1RUDUseDt2+IAj/iLs/0zF5CWch7Vpg6SLSmOQPs12U5szJ
tr65HLwuDoKpORyHmY7kdSYYSqtYj2Y0aXkwaVq/yI5YDmGUmCPKDJCF9l6BPcHx
X+auywSmcaGp5NuAIB/xXhYWP0JU5F2uj9tba8yGo8dDulhKd/V8FPGBfQUhiFUc
L01haL4pzl6QSDDiv2362rBUHBQ3aImLryY+W8SXmvNOUUAn51XsxnHNvf0V6H4M
+k5qOXUlguCJOB38FpaCk3oewnRL5U3O3jTeJ684jlJIKKbWn4k6WJwuDGqos0N2
TUnH1AxK+qtSqxlvIkMwHp7RS3ji6LrjKiBCgA7A4c5MV9MYW2r+lwQVA5+p6ZX6
gb8ftK5qkXkmG4ba9tRS0GzP/hqCGppNG5qxLUF+HR5lLDzn2Wxel5QJH6+xJIKm
JcDxEwlAxU61fiUujALKbMGHW6zIIU7V1hKVj6m2xfNtmc98LTUAlTX/VmJCX4kA
LRs/jwN5TNyB1a/e4N0CBxLurzhCJRKvDdHPGmDCkYHJAmVnZw8PNqLZFnRw007k
E29OviQklPIY0Zgn7CYs1mtqp+aB+ve7oRZu5CklxHzuSWZ20AvfckpXqzYh86Uf
mwnZqaCaYF0yyDUL9ndVZ78HED03Krc8CcHfLW6jRdXhIcrZzIeMd5PMRf7uh6Rn
KxGGDqrZKzhtBBf+XQBzZvZQSo4YAsImc92XE0Cuo4lCNZLJ/AsrBoEfay/e7ASs
t1lzEY7asB5JQk14KSiKHWjb/rVEYB2TNkZXLmg31nd97XLv61NU93FZIEVbLXr2
`pragma protect end_protected
