// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H80-5JA5R73[Y.\W7Z6Z>WWWQ02'99_<7OFU0Y@4QG$\R:"S/203K?0  
H!RO 82(,Q/F0!#_36&HUPWF\]NFWNJ+&:,NW8R_-+'@,C=5">%IFS@  
HSQZ:'Z0DEQ"22&BJ)OHF8M[<8@QE9&P0SX:-0,,4 Y<&FYK>!Z!EF0  
H,J+0L(*P 16=^53.R8?U?4O5_&210CV(',!DE]=H$S D>:Q1^U^'P0  
H!Q%/40J_-G.Y">YM*^R)EZXRR]9)(\,QJEC,S*;LD#I/N2?V7/)]%0  
`pragma protect encoding=(enctype="uuencode",bytes=13744       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@E"R/IN_F=\IWH2#8 &F(/G5U&>M6?;62Y_IHE&E^F\( 
@5>?S@9"UX6![ZKD6A2/1W4/=:NJL?5))(/@7<."[WZH 
@K [A[?")"+&G<T/L4J^![.R5R: 3])F+ )MFZ[^EVC4 
@A_UH[--R1E7[LX\UZ\T[D#%QI@8)W">Q'2-/[(2I,FL 
@$83=;B8%)*S_D+I^J)D-TNH!CS$@>;V/LQ[3&!5\X2( 
@ KD8U*0 <CW)MYC0@C%A6&E?_[YM\HI*/6DHV9TF\MP 
@*JZ//_;"T];PY63$!F@'7L&GZ-07>%F@5(\:>]1'C^4 
@T/1_O[4B&<ZR1(*/6 'ZA1F1= _%J$U5DCGX?6;B2V8 
@ANB$G&^+[$GOXDD.6PR]L)4:?5>7TB7DND$T)='0?[$ 
@WYF^?#>.'1-)\%OCV<9.9GWB"WVU_@$Q)OJTJG#?I1$ 
@.D\:))S@P8*@6OMJ2A2SL>?DK,);3#D]_":<2C%$.>( 
@=E?#M+#4=I6N)RM0>+)#'3*O0?*OI()"E?'.AY]V^K0 
@7G70.,=%5KT'R=$IORV=R=@J:4?+O +,U(^MD[8;[:H 
@P%(U2D@Q);B\5(YZQNO_G#]SS3GU!_ UJT5.!6ED(B, 
@Z9Q+91?.$;5I@1*&GLZR<G/_O=T"FMA7))]*:#4&-ML 
@O/HY@FP%X*U[9&/(SX^[2J FRBCW*+#+*9 O?:S5)]0 
@7@\<0(Z%K-NZ62"HJCB"(:;5JB/\PQ_H6GAZU39FI0P 
@E>E6/2_;E6SBMNYVXBBO=R^'"IA1/,:]_RE6<P.)\?< 
@$T*,*3S-Y,<K(A;ZTYGZ?5-^[ 9_X_SNH9L6H@\(.WL 
@X9?[22V1!)RW5O>=TO.824P'W9%ZDSOPNV>RD_:3N*X 
@B(.*4AI>$21QFZX ,I^K52)0-%!/Z%S8 _W-\%/U<6  
@764<5FZ+ ;#ZU=K@RFD74]?E/QD,)V3T,I8L\73Y;2T 
@>:6>E(#DY8LY.T,^YR\2LK;2KIR7S<<8KM1F[[UG\3< 
@2?LROI"H.W@ ;W*G=><%HU!IA0-!8^\IXJA*E:QT'+@ 
@7TY^Z3Z[W(0:^A)FMCVE;>JPC]=7^CS(H(;(4VSW,,  
@T$IXR[<1%NO2US@C6"4GH4!+0:HT;I,PG)]+\[=KWLL 
@*"R^CN8> 9A#\1?EN?R.K!!0#5.;?MQ1!@)FF3#@_&, 
@*<+)^HD06Q>TSWVZLVZ[7"51:>2&KR"$V 'U4>8+2/0 
@A KJ6)LCHNH>Q@"<K9=^ZVD5MW?2[$57Z$0)Y@.Z_/\ 
@N9,?Z\K#W-M=278JWFT&->R.K369^NT#):)FMO@K4_P 
@G$C:I%-7S<>3:W^PJ34 5D!V7'J]LN5X?P:NQL>G1.< 
@<-I,M-/(H]6XSJH(!3?>]R_RH+8FU@8A0&3-+HSR]#  
@G@S9S6C&+A66D+Z#\I94CQAK2,(CN')&;.+'M)^J-[  
@ )N_N]24BG::,LAS2RN)'[<GN4\>@^NX275'7NO\7IT 
@'\:A,=UHT:VN!0J%5X;K%L'%F3IQS \DFHJQ!Q^JESH 
@5M3#+$"#(@1R&"E<QH)!M#QND *@;SZ3E(]39&/;!OP 
@/.@Y$"/8C*_#A0A&JD7:M&PQ3*PUY0PU3=9[_NR-:8@ 
@&8N(E$AG]LFX-P&'TG(TUK]ZHU#/JJ Y&B3!^FUZ3UD 
@X6ZE8ZCWU5W],0\Q275,Q!8XCD99L)!51&V*!(?%BP( 
@=@<;SBVY!GB2U-0]Q],/Q!;Q),&;8>:K5#S6(8D3Y#0 
@W=834L*P_4X!BJ>RJ'Q 5Z7S[REXEU]60UO(*ES7L9, 
@2A/0S\^JP2L4W\34#)8U[N!I0O4SHB; 2W[&8V?8U\8 
@3F3A^/E?(+X<//706)>S*64V=T&N)1I(F05.H6>N"J$ 
@!!PZDJO>_9WO)!1M&_7.%8+DF0>>0=PCY2B]5(V3N0H 
@^18>KLJ%".J3I=,Y[LY+ WKW$*T'BB8CM&K.7:%_8 8 
@WIR8#M[1)>/*I5/^)M[8:&0^>CHD9\R<WW(H]<5?F+\ 
@RVL,>TEIJC5H$+8,M0M;$7SE&)1I/LC2.%Z)[M+!U&( 
@"5^[IG]WF^BO-T'\\I&?-N-4H]+JD$5FN[F.CP5I4S0 
@M*^>^<N)^.7R7TAZ.8WP2640%#<W+T/G>.)^/UWP'/4 
@@H@B$<26YV\^D_P>!O^7UU*4.(+V95&UX,<_ @K>0CP 
@!BRX5D:,6^_#DY3WX./8>5X$,]R\ZX0 :!?/6X*HDQ( 
@%N]@#74Y!0ZM#P";X;MKA4+0"A8OZ2*=8#&1I^QTNW@ 
@ N W+SY",>H,WRF*<B;5=XXN2UME9,'D67YQ?F4<>+@ 
@Y"V;4-:]^*4R7"2.IWI#V*S&D.EJ93M-5\#&\F4&DHX 
@[N[TKVM3C,+X$,KYPW>.6@2N;(V"#^C,^NN$[RZ/M L 
@-YP)JW,NS,/[*>[WJL2RTF$"?>'LIP$^7<F_I3%X]/( 
@3+8OG<NQ&0RY:G'LZ\'P#C4 0_T<126-B6(7U7<OVPL 
@G7D!A$^G J] H%7FYP6T2BJ1/6O4^8/.:_AJ(EYDI74 
@%8$3GI>M))K@%FR]\=ER')2\/73=@9H= 1,(\HX*+JL 
@VL>0AV7KL\]C*$Z^E@! 3/;0]ZG$Z-5_),DZ!\5U08  
@)6E0.I;[NDUO+U#SSH@0,N<*'\N0": +MJPDS@;J4P  
@BPU*,6Q8EC[<>G'T2]EIHON)%8Y OQ,4\@H(Q -&S@0 
@T<98C#V<3J!.IZ3]=F/LYQ_0\XWP-/IB:UO?^!F^.28 
@4I;%^D.8EOTDH;!!"5_5#")-1#?:.<"JK+M:^E0W9C  
@\IAQD=[[[PQT.QY)/7>,9?F_J1)PZ;(IP>AQ/(.S]HD 
@*]?N01F+DZ^8W*HB%R(#UL0?P1<XJ]9WW=5^YTRM;KX 
@7%C =K^WNH$"MBJR&;)] HE&S:>MI!'T*ZZ:(' 1O'( 
@PAP^L*&H<B60"#":[6YZ65#/T9\.1_%[/2+J)-=2W\T 
@4R^!?Y1E?J&/()"K\P/B?:!>$#['WX01[UO*19%ZS0\ 
@$"U)<_@OQ[7_#3E?A,#&YJUIGN#O610KR7FR%7/^ WX 
@S[UB'>9L2<[ZP+\;J*Y96FXLYQV@N8[J.GD;%LT%D$@ 
@):J&?/9-6VG5"!SURS.R(W\]:/ I*T8I ;?7=JNLM7  
@=R)H+<*- F7^['HPGBB"".:461>T-Y((P68_E(9JP!8 
@%.P&HESUX%"%P3-5=JXT%ZE,%/3V0"R6'=4F"1( 4T$ 
@LJ><.=3R. $\:5 MN(=R3&&?@1HLDHZ:O__N3:.ST)( 
@X)?]A+6\L>EPVN[#L4TQ'V#B"4LQ*$( G(]GMH8[*8H 
@G (Y\1J[ZX,[<.U=!6;@@I]_\^7L7S*+'(D3PS?QUX0 
@3MT05&T*YE-TQD<NFXB5C8W\<FJ8K#:^AKUFMT]23(< 
@4WC%PM+U%+2CMIRFI?_*20@_"(NDTBZEF9_Q5LYT</8 
@\+-@A88-^F@L3'VI8 )T68PAM/9K+%_5824WL.CJ%1, 
@3 8R5>"27I+NMX*O[<Z_<+36TUC/",>=V^[]S+5?>Q4 
@ZX:S0?,'K8N*Z.WUDOMMON@'QLD;*#W"^!@D45>0VZD 
@[DV[ O7JD=GPE+?/2!8CWX3'&!80HL_Z)FIV=0L2#W< 
@"FS[,D96NWNDJ6X/"8:4\BS]^RGA9?DXBB[8R1LD<38 
@N(KK-E'R8P\57X5NN_4O?&:(H@'[Y#II(8"$7T[A@GX 
@CBB50^N_:[/%&=S6/F>4O^-ND'/58<K)#JO!U(?JH0P 
@9_:T#DCU.?K+],CK-<I"$<JVP!;!-9A$F>3:^9;+$LL 
@M=S<H#O'F=_[E_7MRU'S)203H[D:>=^GK$AI_ ^%ROL 
@/(U],T8O=HJ7ET1,H_!;X% @I3^_[7K5]V8[.!P7I'D 
@,B2B?=_C"$B$L5U9J:U)AL9ZE+![)M[T-EZ".WG2474 
@WY5AEXV2RP_^D^NL)2#"CI8SIO<&4EJ0T+^="="$L9P 
@F(KDSKI_Q*2)V=V#7[3>T+NY9<L; 4BIR7V$IG.^0YL 
@>=L>'[T/6_.O,C&$*RU%^C7AJ:)B(0[_K):_.9^DGLH 
@[H5/F0XW !8N>;/S+R*=:-1A%AC)PM:J<&,)0JE%:7$ 
@1<V]HT<-M1M;0&U?P(0:0%&0&FTUNKMZC/EUKEA$61, 
@/I 4%I]T7@;9BEH354?2B(G4B=O6 QW8H+^!9NHIF8\ 
@";6^0G+&132;F[V'&E8RB0QCYWN-1[<[ $C"O$09[5T 
@;X^U4]!Y&4(Y@E(D@$S4>C.Z"H?J46?9?=NBL0%66/$ 
@NL@G(84Z!79(ODAI7"+MDQ,ZW/?.HM&O/4SB(](91V8 
@>7]MF3\[)VRQ/Q498?]#,SW4S3UNW;/UDJY4B;RT<Z< 
@0>L/'IP5R9V%=>M*,TD/BUIL;^GXG+7O:E\JH\]#JT  
@!DQB )WNXKI?WU!4NO?,I]+XCZ+_SF**T!OVM1>Z?.< 
@[YX, F7.R<U1#K9J[)V( CYY/H[V=!VRI@(OR0JWE=D 
@9_PL-193V![H727E^R$>@4%"57'6G)J4\21;=18Q'[@ 
@KU(Q6Q*AT.\P8'57$3J\VML;Z"2Y>QP]6ZAOSJ%A,B< 
@<:(V'!38R#<8<UIE7Y-W?Q(0.P2B*5<*]TV"+GFOYW  
@WUSV_;_U6X;;CBS%)**C5WNHP%GC4/P66(AV"D%W0%P 
@+$L%M\N:AL"A@>X_1<@]>1WPA<:=!Z/6Z^H%0!J<FF< 
@ICHQF^GL<=J[GQ#OTB#$+Y.!N9E4T_-SFE.SQA#.5@L 
@C[NP,&66$-XLZ$BU-(&1W5-U]&+ZK^7'3@MG,HNL:(P 
@Q$1KB!4+O-#O<N6L*=V##EVW#42-N&?G&-)T<[,3A:@ 
@*?5B%TUI2)#3JII]IOYA4JX!18NN^0<U)A(-J4)(Q2D 
@1RIJ2+CZT\D4X@9[E#<L3:(N,[5\1_W^7H:U$3Y]1>L 
@?D$!J1\]\3G8.8UFXP(2'?I$#RU"G-4;OW*Z%:DV3IL 
@\%"M]*!T2YM7/WQ)P^ONOR0ZIE#0.B.=+,U2A'ECVM, 
@NZ_R\NMVC] 9Q'!<LLIU[1G5G..?-F,8V7JF)=:*+NL 
@O\'AN[\P!.',8"(\L#L-"T( =P"?Z@I4#73DUS(3/2T 
@?W\Z+EE_>9VS+*O1"%N6;S#1FA^0X,_X&9([JJZJ_6@ 
@3!G>R-5X9-#<OCW#[$*;Q=PIIW4A8UZ+VXXXODQ%40T 
@L&5=[Z>84."3(:)9#O>OVAY.^P\5X-735 $Q =75)Q\ 
@K(Z]3T%^=&RM0/=$U[7:RAH(]^QGO1[\%Q5O-;%'D@H 
@R%U&A')'N)HT+ALMY!@$I*<K;(^5'-V+&Q54K>!V_L0 
@+@+Q@ZE6!XP KJ@;K1Q(_Z4A0H9E_D\:/@NQ4B6!%_< 
@D(S7NW%A:6$ CIQOPNB8.E@SBU2G,B3X2UNB2)'9N., 
@WMJNPP#2.N.U<Y_'X8MS,9M!MOWK=>'3,US+R4,8?M0 
@G!K"<5HRJKC/Y=NPU*X^WP49U.W/^A$W(E*XQF9^-]  
@AE- @%O-!N[D':Q4WM,Y\PT7K8$1+Q<PFH8-Z3_2T), 
@_>ZU>SJ6R,P@LB-F5N:#0UTWKI/5Z"9\=^SRI01@BM8 
@K !QGJ9)/&]7+&<F+WG1U55IS$:4S&B^H33&V_?FYY< 
@0O%S+3R*!]/H?8)#TW0[T)BM,L)'V Z5LRU6G.H $'\ 
@NA([MU3]OKF5[#8X4@,^(1.YR!+]TS(7'Q_"1(>S7Z8 
@3/%A&]\,TGSS+51<3( ;2I2Y5Z>?B2:YVY*7IA_E/C( 
@BVS<%8CA&%Z>8!OEA+%0F/F0!P&PC*^R"6WI9MHV2@8 
@V:9R5SORS@][\_W,0H,,HK.#YW"G=B1?LFB=/BR2;<X 
@L60\.)>S$@N8>CHF%Z>,5@"W.<UI8BC$_?3Z=Q<DG'< 
@QMNG5D>FB$@F04&LK2CB]2>5'9&S\!6AV2H9J4SMK6T 
@2/ZC-XR<6'&DDN8<9P?\Y#S.<J96#3FQN]IJXM!IR!4 
@;2.J G#E>&A\XQ\+)B&+VGG3RKR;FDL_D5A>"A<*U'@ 
@)SVXSV$,P8WD/V+WHD(8=5^&\&C<N7D/]0' S$CF^F0 
@@>\8UO3T'$JR]8"[*P,)LR)KD!,M[/]FL6N<5,Y9L4L 
@;6L13@LP#72\*%)T4 3FIQ:PU\/,O?JK\,/X3<IVMA  
@8BUBJ<MF&4DYN(O]J[_Y"[SZA(&==9= ?#8 %T0-X*8 
@4]ZL?J(!_0T_:";+$]<#(4&*  G,P4^EEY-7>]:19N8 
@_[?XEE9L[[":BH> C[,WYNOIQ697UPPOQ;D"M\,7WQ, 
@PP'MA9Q7JY3)CE8WS#';#(!X7JGAYW+$<9IDVBL-5,< 
@@6<A[$3= 5X(^Y77IAQ[$A;6;3Y4EMK8A2 J[(F.^E@ 
@H5$MOYC!XC1V4Q;8L2M'>9Y=&8-0C_6398*H>&3V![P 
@7IJZ.9B/Z-;U=]@?,Y:N"\<R]*9.HR7ULSIUQ.+_?F, 
@SA"I048'#.(,P$HB;)K?LRZ0*;.<L(FI'+7MK<ZA5^  
@_>-F[]^PJ28#*A(P5W,9IEY-!K"E+%!X"0IO[QS?BK< 
@6[O9%8%AJM(3-FKG@\3  '+-^D4QLS!:>E>(UKYS,.( 
@K+I.,_2JJ>1VZ?7WE; S9 #>E2[1K9<8HDF0-[P9^3< 
@]#6?^@'/.3Z/9(A3OCH94?N5$@3G+$-@Q_=K$JCFZ=T 
@H#B:A:,!6ZSZ U<NG8P/HHUJV'MZ%#CEX[2/2_PI<8, 
@%7>8-;']]4R^E:9.E97 N]UM^UND$$13X_UBT@8,;[D 
@FXX9'B3*)X=+N7.]VD)<O9G*.^92_[QR&03J_;Z9?.< 
@6RG:1K6*[22;KL[W"C\%_FL07\0WJCJ/4G58()7.'<@ 
@J4PE@TADI:QE?O?B>H/PSHO(Z,(HOTI;_AQ4P\TKMGL 
@J_$+ $G9QZ&;^6H6O1JFH)ER[R*(@!'AAQ6#AAJVA6@ 
@CF5I ]<CG2/2]L0 I7F%C0EA/WC<;E@6E)[B3(QC.?( 
@YGE_HJ6FYOZ@G /NB:WX3)VMC!I#FW;Z.(*62I*C+G0 
@5O9X!4"M'QR*\,DY]ZV5K^F*'>VCV@>F>FXQ3"\:0I$ 
@>_%/13PQK_J*[&_:; P&:V#Y]OM2Z;I0CO2U\/#D29@ 
@,N"@N\!%>X P2Z@N38RH70^2X^U0A]I*!-;V[YU"Y08 
@(J:98R!')G]0TU=OF_STJF!<;S\S S0LMEW B6R?[%D 
@9HRAFNM%"XM_J#&7H&-W!5.(^ZC9QV_?X=U!N3>4^&X 
@JH4CIY)SOJ#8%P:0;M9#<8EI5-7 +0HT2S,%AH,R:'( 
@!<BPP9.[O<T+\U]PJ7GL:)1YAU)!%%7F%)_A;[,7@:@ 
@$Y+#6UZU2^[XG64(@S/RTF9[E?U+!&F7'QZR*N=VTW< 
@)+S<./?AN+TSU*9^5ZU:9?0J+&Y/^S.$X"Y#@1@)<&\ 
@-954">NLF GR^K%&Q0"OZ(1>/SBRE#=.)3V36F0R27T 
@/X8Q<#J4IH T?9 X$#08BFK:>8C@[WQ")DB:AR_>@XD 
@8R#!AV?[S:2*X8_*N83>CP\20A#,.C>C*=PI>',*-5$ 
@Q*L[6-_,!DL-S$LD^T.3#=0H[Y&K-2>T*DXU1S":2-$ 
@XM)RH#G 94#@<J>K"760Q%'RRMVN4Q44R-?$@+/'48$ 
@J3"7Y.)DR*FNY)_Z9DT_Y-&2]A'W)7CE]#6^,X&89.D 
@B JS7[7RJ78\3\MH[:1W5VJB4USZG8KU8(E@U*"G8*0 
@0'\9,-W!@R+R!\N-_]+*R_@L(Z)J$ NDSD#69:W7KP< 
@/?/A7:?*F3624CN5I,@1$]/I"_P0NCG/ZGPA,+*+PYT 
@^U=ACN^0 ?$/+5/$:# 6LK*>/ O5ORY0 W>F.ETDI*D 
@\1#TB4W9:T(X#)/FI\G :;U,X$6L,>.")!F6D)\/'L$ 
@9=BA/G^S6YS19F%H3_(S)?-:9P:669 EJ6V2;BE36E( 
@G^^%K;'9V32_NN&5:Z<Q.9ZP85Y\GS 3"+]-CI391QH 
@=:T1!:F]'"8-(!6![?;B"+OA7MU)C(#/]R\O3%ENN<L 
@L-/>49G4)0B8#'GZ,F5X,_Z^Q$4CZ(!W1)=M49%_5C@ 
@['[4IG=KR2L1:=KZW1R"[C@T:5VV.WNA-*M1/H=4>BX 
@V15 &JN^W-"ZO.<9L_GJBN8G1 9W2B&0J^,BA<I<8T, 
@CY4OF;:3LG@]IMN<]EQF5P,B.#?D] 9S!MD>R.-B$IX 
@?N5E14UDX_+D)':4 CH2@+K0LQ0^!*E)HXBO0N/ED[8 
@SXQ@BPY]K,/5C_:%.3VLDE/*V/&8)9[&_H_]&\H-AC, 
@6/>??,?\04L\:+H<[4E%1X$_,QU7:<%D*7B:G"RS9]4 
@: 4G>@$6TC>E81^%4*YK*A])D?FFP2U$(!BSCL0DQ^0 
@43XC#+UF@])2D5\4B>;2D@VS!ZJ='XR(_02PX)67TF  
@9F<7LE\7)<<-=)+?%DU#X$!. 6FB8BD9A=$Q,4CF X< 
@X"$D8=A=?!4G7*$M0/.2V=Y8ZQE(+)/BU"?Z4$7("<$ 
@Y _0C-%&G:,Y(<T/"/"VTR;]1_43XOI%,;>T77W[.4H 
@)G@%(MWNAV_'"\Q[W6AJ&JD;_S$CBTR[#Y=,\F#ZNW@ 
@9N>QF"6+8F_-JI_$7'3## 9BSEIV>1H,^5CQSDC00$\ 
@4.G-X\EC#B%6*>TY2V)!JU@>K5OK(7=$CWH2ORGFKL\ 
@Z:#@YKR3&E887%=6 ,^'4U!&'M0]HXB'C'?WBB@[O7X 
@3[?Q79P?A$K"&B50VQS?O/*RL'1(#YN*).*1!R*->2( 
@-B_>SP*RJ*]-[XK15OR5X7<,UZ9_DM%@3?DK:;]WB;D 
@U;3O/N05C\L))H0RDI]& IN7H5&&B67[38^[$06.%+L 
@C&1"W]_2\AI^$&)3]XF,-C%1,%'VCS0H_X@K#,B,^?( 
@.!MA3+C.05%!=^^TF%R;XT \A#U*#6 5^J6 F\XMWD8 
@2H^8JB&7A^U;DU>:$%;).BA^QOP'5FXDP]W:G?U::2< 
@Z5Y3&(Y"V87%#>7><?:FGJ_W;H]#E^-0N$A)/5#] ?8 
@^]95^_K.HC9O^BXS^*I0UM[2E-68 C?8J9+6]1MQ5J4 
@^?!6VI\%BD/3QD3VL@U!A8R!2VZ<P8'Q!>DWBADT?(H 
@>E(L0HP#6P'2E&J39)KF' Y4F(P8(/0PNVT$^=Z_U_T 
@6\J\.ZZ 7F!=LNJCZT2XJ.N>]V\[^H=B@]?= BKODZT 
@HN'W1]=!^S:O@@J^T20-<2N< H9@Y)H,GY5W+V@62N0 
@Z+Z-<-9IOES*/*Y@V'#E<?^6<^:G FW&7-EGE>42%5D 
@@R<OD&QF"$%-6Y($S^TY^YXU\MD^;=B4X/4HV9,'V.@ 
@[4!K88^<<T9'^1Y(YY0TB')<:F>^&FSJ(>C[BYZ5&3X 
@)0@@RX%PK9Z+OP"TN_?4+?>_F/,L020"Y0AX"L[S.K4 
@-YY$]#_)\-.!<>D<!&)!W'4QK.=[1*%?7%WV$3^<76$ 
@X5V<N9UG)WC#YE56E(<.M$LD_I-YD+$#S _\Y]/!;VL 
@_\H75XCS+=PEQZ;O-G?QB$SL$:]"4MR91;!A?N+4:7T 
@:X MR0J9L>"F@YL*]U6\*(4893U 4M8.8J".B)M_UPL 
@(5^>?S,+81)1=#%5W4'3N=G5^%-JZS 4/G!:0@_HPO< 
@%$1$K5($Q?QDJ?=:<22]O39,5MD)%9>!J#; -.<;5J  
@W['V8W@]]A;8+03SF.I&RX<X7S>U2*UQQQ4PHR6!-P  
@@^3 @(Q(7"!4$\45,36"F$S+63$PO]4!!0OV,0.C,EX 
@^G1#UYK6C+TWS/ _)>Q"L(TLLHI&Y/@1G6X=GAN>?$H 
@L@I@7T#7"Z$^7E) #^&6O!"R[3#)_-S/^?13*B&OFNL 
@%#51"5MWC#:#K<21([I'-V",%A>D<=VH.PX!1->ZN L 
@8>ET7VG[)']Z.!].J7!BMHU [-DH?%55)QWSU:#6;F\ 
@PT0W)MFW-&5"() #<X$F.M0L?HKA$O81UNYF!O([ZFD 
@]?B3)37VHM!Y+:]AVDN2,F+^WAZAYPGWC>G"SE:24+@ 
@S9D2/4>HDXY_N)/BI\X&M;'\J&<-%6Y?.=$R,P;JPQ, 
@O&276$'FQVE ^<24_!)A9O-U=;(+W9F?;]NC_"- $D  
@)PU9@$=#I/MF9?\MBF9(95'(@%TBUA/S[F76:5B2GI( 
@N=-T\FA-0>P#[]KCXDV?F*E9+#1%3#$0AW6^RHD$28X 
@92OWUF-MYX;A^M]K?#0;M@"MQ,0@G6N?8=-F;S/_J$T 
@@*T;%/F@44O:_'(?W)J!G7VF"-_-F986FFR[MC[-I$4 
@'%"W"IL#ES(D"Y.;9&)6RME9G)F;("OL&.O\5@?%'[  
@%CZZF2<^& (%0+"Y9!/7H43QE.B;;,TI$01L&%"4)+, 
@)9$/P\]M.]CF-Z\Z"\JNE*^T?Y@P_FHV,]/QA\4K7&\ 
@"LFQG5_1>^+ON.=YVO0E4=\0N))<9R>/+%(![R/+9UP 
@&:*OT4Y*_:HYB81&^D(1>F0>NX1/V;F0?"O>UXZO&AP 
@4'./E+WHL'=YIV[BR!*\<#VCZIT+Z\.[[?^@G;BG,#( 
@YMLZGKTJ X:9[B-I*YL7W()"VQNZ2CU$ AMQG^55>R( 
@#2YJ72*]G2EA*^MK]U&+JM(<A_WD%>_(V='XL0J RM@ 
@]#ND!4WS,*V$XU?F3^/3C\&#YX\59TW* O(V+%@R:R, 
@8ZU"-"-?>Z&JAI:=+>Z$5ZJ>$[FJI!!)%@T[9+-L$CT 
@G_7D^;@FD!UF;7%=;@GCN(CG[V4WJ51%[W07WO?N__0 
@(G+; S6GF"Z#Y%T#XS"/A#5_FI'T6FQ"VE0;%][;^5$ 
@<'<U,_VACT=K*42R!3]S;8QF< @0^*9]N 6E/U3!+NT 
@$05:G /A>N\R.G9D9-0@/FYJYL\N\[':X$@NS0/71@  
@5PX1.7V=Z+F69%V<WQ83BSR+2\GSSQG>FG186B;E[2\ 
@PO+4D3:'_X+?MDA9/U"33$Z.OD#2N8X5/HNNSX]7^,D 
@3G:G]_*F",8237GJD#Z*OPH?K7[.<D"1ZSOZ2Z"I(&( 
@Z3/=P6H!W M_?.-;F+Y=TM+4P])GJ.4Y+M:FI[Q D=  
@;"8#/GSOG!P)$[(8@MC$HZI?B7AS18@1R/3AZ_MB+Z< 
@%M0XM$9X"<:U*C:$1N.:366(>\YW:,$P?S=V==@JG<( 
@G,KZ9:JNA)?0G<SK,O7PH;]6/'@1;V2D"AU$)]96=FL 
@Q]3^ZO1?T][LWHPXY\58"#G>ZG;:)BH&)FUG'=D2:Y0 
@=3D9*+]6YQC/*$+\/>].6#><(.8!.6N$IN-A,;TU[U@ 
@;CUHX3Y;%-$V-@V'W5]]_(!7)XQE0O%E=^B:D'6FX1< 
@O6!U*HV#)!Q0&[%D>=5Z NT1]K;DV+8R_G1&HZ?UQZ8 
@6.4X@*/Q8&''X7M!X8Z=NY+.LE&\X#U2$"[14Z*?+WX 
@^%$RO>J.2O^E;XNQ72WSK,)KL7[JGKK!OBKT:0/Q!/\ 
@EI*LY,&Z+*6+<41OTSRXGP/V_:X'Z27QDWE])J+2*>  
@]Q(F@F96I(3W+<LG;<4$M!-&)"U*&TK*IY+56/4#2,H 
@QUN!0.I\91$):;*JD<&"W:IFQ]P>KI7TV!2*J+NF_WX 
@CR4U],P=^O /I7R"O'<#Y^.E%ZGJ'EU26\+BU0U/YD8 
@6PI7(C^=J":8[:<$$,EV2O#8QI(Z\.ZAAZ*]A$?G5PT 
@*BG!9^4C&)*K#KE$ #E7]T[9?HH&X'7/\>W)4+BKE/< 
@@%UI^,_CL)M3D4F*)3D?!+JECK*51EDME#[Q'9)[^>H 
@0_^5B@KH<,G7*@GAMHYV@WR5/Q7B4.;.?LV: 0G^+2X 
@K)>X&RYR\#AV*'-F<RIP7EW*KQ!*5:S"QGO9>N366M0 
@6:)_22$BX,- O.)16#N%G!,.^-]8VD4?IM_5%5RM6"P 
@/=DJ8H#)* '**D#3<X4E=B%%+-7!>"\O\;(*8+E705  
@'=JRN )WHUR(D,^5W8:5>J7M3PK^]X^#RL1SDMPD+A8 
@T#2AH+W=_[3(6HR-AMUKN&^B#CP >I:WGW1#+1EJ*80 
@HZV&M*BI_I)N0B)KDY/A^2O3V#W-IG9W(%9,9Q?C[V@ 
@C6G2^#*> RCOM]?1SMP8S9N)4W*N<\SHK.ONM</FF!( 
@,2CG"9D29H+B]LV*-C?%X+P:"LA);;!SL:*:0VLCG+( 
@4UM"NWHV*KCK_M&.($ 8)]/]?6:"5K0"#/Z,Y@&9Q6@ 
@E+UP3Q9EV\@MM42<ZBV936%2OR,<%4DH=/,,.PIQ"#L 
@<7\#X;LMC_G.?YU=65T8@M*P+ZN"4-+H(=3JF==@XWT 
@]2"3%3\QW4]$DH0AXENA^:[2 NJ?L]J0@-,7?:U6H@8 
@%5Q$SQ,^T)E),^_L@$L==L_K<\/QL@!&.*4G/?3K-RH 
@8TYD9\'+1AN1+?C!S;'Y/$Y=4$0YS>@^,U#TMAQPF8\ 
@X 'S1KA7*>[=2721-<^MU_B <E69 >_(<<G3<F_DGP\ 
@%'.W//91C9:"Q^1&%&,M T]UV\.(4>.IUS \0$<G:8@ 
@=*Y"QYB),?7D=V1/QM9 W])<+F-3T\;GE7,(;QIQ7U, 
@K4/T=W+MU!]\+%LAI):,:]?W#NT@7&_-?!K:#T0B4&L 
@*0B B2X7 -WENYI;+0;BEYD68@$=!/"TM%!U5,?4C9\ 
@/.LP:>"!8X;FJ!O)]@)LVY3>JJ2>CQ21C'),?*U.U[P 
@PK9=&'4/M"+A29@N[W)T$?[7QMHWF!5\1EC!U+W5*]L 
@1<E3592&V=KF0]!7 +X><?[EJ<=(3IH*7Z;7=TH,/>P 
@I^/,ATOJ(N5)/ZE_*0#+WS#554#0#6GVDB+QL;[:Y=, 
@$K#?NM'\EB6=7 2I0@/(MX13:KIIB2@(:F#V>C30?P\ 
@UE+/=%D"O\ '\Z$T[&S_F$=2>Y_>B3%"^(3X9B4U6$8 
@?HZP Y$Y!D!3E',/'<V2(B!9:8?S4.<I2<R[ V6JU_H 
@&+5LC,>+A87P9J[)[NW)@ @N@2K50Y()-5<E?6+"47L 
@C,E2_LFAC%QLO,:';,9X85?UI#\S;(J/4CUR32Z$3'X 
@T-<XJT:['SOB%]BLTJK"KRKJK$>E^Q;68F3@F9Q=RP\ 
@W3F[@U7\OI7]'3VE,FYQ_,OYG'ZS_>")4/5&\][P@@< 
@U).WT5!E["$&Y/5,_Q/Q1AXRS6E.2W$OF3'L!3%@:0P 
@'SV]:K_?YFF:R"V:\=69A/#"R6@[D#6S59>HN]&QD1T 
@(',$,=H0EEH2BJUL4EGJ7*AY<^C+*V*Q8@@H#3N#7N4 
@PDB!M0NMU5=PKHI0>1 '3FR6_LM,W1YAD",4-I03G'$ 
@?# UF,]>#^T*8#H7-/7]DE]&A7E)KJBPP]JRRDN(>[8 
@-IO?=Z,6-;<\Q&M!E(V?L.K@/11E.36@"BI<23;.*H< 
@=G28+\>G$UM0W<C,V&"M"GO]F/_UD=;KI+3IFL=2E$D 
@;67-Q< S8!=L1%*:R943YRG(^1FT'9N\#B7_J%.9V0< 
@[ L>LYROSRP\_\B^MI@E>M?4-*[]SZ[-V&9[)Z>U)VD 
@.*S5#:+Z="*H_XT89;J+ __G/YRQSYSO3)/ID(3LG-( 
@0S@L]H5=]2L6ZT=U<"A$^]B[BE-PJR/?MW6%AB#*1R0 
@+"8;I[;GCD,&13V2=KNA&1'42O&% 'IZ?JB@Q4IMIZ8 
@(#O$#?A'I>0)7 C+ZRQV@V$F,=RI#;5^%F++?K_Y7.P 
@=3X:^/=P8P\$5JQ#WXAW<*.<8D(BC(8044]?,?LM^MH 
@3DF/THF0W2I,!A"P!8H'H??4_J*OUX#=_75KY!6S3]X 
@V>:E($8@!76VM5T6CVR@J1<BKV0(FIR[74"I\.]K+?0 
@B$B6<3S#P*%AS]._RF"I83F>[L,Y'K] &^IT5X<.H>D 
@==7',HN:C2T8GN_>NJ]7:MW[V%-)(;CGKU!QA\+;6T  
@4_LZ8GP?DNKGV/7:8^;1P:XLRN)+1+;:IAWM^)>0EA8 
@SMDQQ$5AMEGB4 F\0MQS3C)M13+Q[4@Y:<.C0\"NBHP 
@V*YV)/XW&CMQZ7.WJ;K".9:MLQ9#)Z^70I2L-I@S2*\ 
@BT9QB&R8NMNHHQ C0B2ET/ :BW113KM>]76@"NR_8HD 
@7 HGA;(*GJ([PQQIAT).U1]-T+":O7>O!_\,"9;AYMH 
@KER_PXL=3S.^%1F5 M :LI82XY(-A5AXQHUS%_BMA!T 
@=S-AXLNMKKTR(4A.!O"R5-#A6RN92LLBW673J(#,8 H 
@"*0(*I$5NJN6=+&+\&0HC"9*.'FMKJ/YN%NHLVYYLJH 
@+"??M?Z1.?Y)#^3DQBI!V&O%^-&/I,P\#+<[<;'3[&$ 
@53X1A\TRF:93J]O^H4=-E7P_7^M[CP"+ST!)DS*//I( 
@=PSG[-G^35)",EV$E+&6MRRTV#+^IRDYYC5OOV .<Z0 
@,*0#0VV0?ZR?TZ=<TBL35*YXG!SX'(#'(M@N4;R0BRX 
@Z1BV77I\?9*A%8KA]M$%C#QLGID0.>ML$V/;!(/FYE  
@/A@OVB91;<C?*,3]2!GC!.64CN); Y1S"I\R=TC02I< 
@&7:^[3'&PGWZE_.)2G$MK]*OM;]$*V9V[0V)P'.RCD8 
@@H_HY)(P.>L/#TJ7$I2]%@S*1\%GH!_;V\B$S%@"?0$ 
@EVGM8E^W);-6R0NSY_XA)"M5E=TQ-%(S5%11GV<)XZ< 
@8-B\.("P)Q C#H_LDAP2=*V+(H0-[+E!FTQ>QDC_;MH 
@$$</M?-OPEA>4?PZNVU6ECX29#:@X3U2K5@DDT5XJ8, 
@=LO]N/2&&986IG^-G&!U\7?S5?"788QR9#GUYR8-5HX 
@$I#%.@FDM(O^[M.743OI>O!J/IF;H9>I2$+-45O!%9T 
@KE)5SYHC@F-"2[K]P5LRN6-$_[^,K!0,[$7*IIQ#,=@ 
@4%M0_Y"LH<89%^1"A_^IWBQ0X*J:3/:E1*FT-;&+"<0 
@G6D+T++MK,\Z9$;D]")%9\DDE#&=,[_(#0#C-U,9!=, 
@LT'<#.J(+4;8&\TJ]C_+M+4/6705/,;1X>K'RVD^#?( 
@,%E(0C>C_HC<G!C@-KI\5I J28CBE)#UV\_7\]@=R'4 
@S72$*:#2N_X6=[F<##QMN#KL"X8? M"=2-M5#N#5O#$ 
@62B/\F?HR ,RMZ#A9 IO]WY_ 1>NU1IC[ ?GTR%)<!X 
@ZXXVF(R0,:&B/19GBNW?\.)>@6UPXFVYH4PU%"2_KE0 
@N1.QT#B.H*/^\>Y9%3J]WG'#IC61I"S?N^3JQ(>LW78 
@7#IMW6.*!6X9,Q>V-6ML-@\IA5HXNTV>^6[$C7L*!A8 
@E6"M/E]*9DMH8:T%B/*=B_<K#3\H737\%[+O#[%*86( 
@(:#]$DK0N&*S"D+QA[A^/3(S4)OYHD([!%0@LZZQ:?H 
@UONAAK42M3F!)B*C,;QRA>[E0VDE!I7"^U^;CA8N^1@ 
@/KHLW$\48VG;':A\UB/ WS%0'/+3-6CUL7YVGUI/"1H 
@P/UT.?)4D/$?ZZS"2]+_PKP^.9>4HV G(5<_WCX2!K8 
@PJ*%9V.UY?'\@M NVPWSKN D)9!*KJ-5OW):C <!G<( 
@AOUC!H*<='I+&=%IO("2<1FN:.H$T)3'H>G#RMU7U!H 
@_2S;? \LH:- @>$<E$';V4?\$,RG,R[TI5PZS&VI@_8 
@;MZI_S4H;X4<LL_4JH3_"#@*0[CJ8J<,0=E?KV70& 0 
@5\YD'-HBNX9PLGWU40#389J6HXBAOMS3J'"ZCOL,!=( 
@>OE1S_^-#U%)34^F[-2"0T[JH"VZJD,D0J2=*%-CH H 
@GIRQ0#XUQM$ML.L1CVKK)5.U7JS$&RI,J1'X+P98Q<$ 
@KKF(P5. QF[,NI%M.Z>B!%_-SWR0.E@C!ID\"P-\:*@ 
@E!O&TCYH/Z>*S4IY-BS:6N[$%OZ2F78T\'X,.@#L*?D 
@6+A;>%V\F6<LH\TI74Z9JH<O33O$4M2/SX6MOYT9YT@ 
@X"LM;P2U[I#BG&F??EH&GKDL.SLVKZ6\M)6L6Y5T.?$ 
@!]\>EP3>.,/@314$KI]KT]$H>Z4,EK4C7C)$-0^QU-D 
@5W@[M8(33(T>_+)L"H%K8@)"<SK<5'4429@%X*D:NNX 
@"#EW648'6_).=-B2_/8Z.86/?#J)J=6&]-*VG#M$84  
@H2SA8A]$@R\B;WN"L?\Y3LO\+SSIW)GZ[[5'N07BI;T 
@($]H)AS#HT&TGK7(L;F=1!(;B>HIC%5Y)(V:#R76H:0 
@7<668EZH965#?^U;J"[J:TMWP\_%U\+FEK1PAYD0J!\ 
@8\0-78B&C=30FR%M]X0ZPKI"22+_O85YI2>-E_E2#_< 
@KSJ/]]]QSW=!$Q$6H/+"RR<-_"@CM>150R$"9HYNGO( 
@[Y-R%6KG?^\TFO'+-)ZRIE&<7J25[ZXO>:Y[M/$V<B8 
@)'@L$;@:RZ;<W1PI'F2H<@G$(K9:WK]#MVD&&PP<Y!X 
@SA%IR*[19TS&2POQX!<OXT[8SZ2Z3PS!;7)^W&KUC^( 
@"4W91H?T L1-K./+KUK> !AN6&WGLE&B\/;AFFI'=4\ 
@Q=FT@4)3SL!H.F'E'.T[5T='IF_Y>ZD=Y(BM-!0PJV$ 
@[@76X%@\SQGOI<_V1?Y$HNPZA+A\VOG5?."76.J+K1$ 
@%8'Z?755ZO7 \+.6_Y?@3</5QPPNY5@+-I%0 ^@+S8T 
@G3 I.%P>9\B7\9Y^R2U?[QIWJ_(].KC?O-=SM7!H?0L 
@&F M;_*\<98M?5 "P. ?4%C_Q MHUKB*YS9>Y%I2OC, 
@%-88=:@94F+:W$'L9/H)GTCV<@EEG9T#3ZF(@T NEA< 
@[YWES&[N, LGS;##(X[.';)0Q#<JL?67M=P5<WY7FQ, 
@35#KM111&,N@LSAPD3Q(O[ ,]S)&1=MWST  77$HP0H 
@/TB D9 ZROE+,YLFFZPH6]RPNWV-+QOY:"DS Z]Y*_H 
@F[07CQ!S5/9SONERZNE<S\'YU3;7?ZSY^9G8EIB7L#< 
@L7Y5:SV PV*O[IIEUT6B@))^O-2<D@*+AG^O0U30T@X 
@XI0KT'?B<!ZTJE#608@5CS<BKAHZA_I$P B(*T;X4>\ 
@V42WX4)G0'L"E[4ZQ-0(^OF;#EM!":+*_'"$6?<C[ , 
@:Z[[[QA1!^^06L?&;A U=@CJQ8]=HZM/?QO5%YC@-^@ 
@C%,7BG.&^W#5/'XXT")&E))$+I7-]P]3_L76[(L184  
@A(U;?7;R]0G2\0;@^_"$!:@O>:$/I?O+8T"IC=$7AHD 
@BW(F-"U+!&"+2I,:[&]+=TP"6>:Z%&XWS2D::<=Q&;P 
@:DC0J369ASC@6, ,L?#SVQ!6RPEW;$<V>F//&45QI4@ 
@]K9Z5KF)W: JJ02?Q&._*E):SPK-G#8-@I5^L>P'C%< 
@@WH]MN:6;'E7,>)8B6->RY:BJTJKW9C+P^),@/*FS54 
@<^\>+PU;<Q,N9O=DZB]4C16:3Y![.GE"B']Y4'@TV_H 
@.W,*&.HA6BSE0-Y&4%F  D9D1<%HUCG6AI3M2%#_A4X 
@$Z[,BPS$ UHH,+]W=!;J=AB-AFN['\%%-LV1"H>TZDH 
@OE+$=A:22R3A3J*3ZX3E0)"W)3W26%*"QYK>.<ZNB>L 
@.V>'D8P2#MY^,I9/2KG;-(.C+!2.?R3^TN/EQYBY3!  
@?P1=T<<R2IAN*K&U]X:"B1J1_IY@!*- )201LSCQ8OT 
@"\]%KKK:R["^$/NL(4>E+8RJB@M&0K)=-1W&&:GF?&H 
@N3H# ?PT>]!:)5P>8=7:[&Y]  ]MVZJW 'G=%U-SIT, 
@10!>R5(9X'JB8IP+-,%'RF"1L?Z3D'NASF9#+/*14AP 
@961OE/$RBXT1^Y&)%>]F-S-&O*(<\1*TG$%OYPEM_U\ 
@DQK>[:>P&GW4&P8+<52)P@;CD\R*D-GS4>$>IKY;V?T 
@?_.=X_E14XF5D4:CJ0R0"9() X_N?18-S-*2KQ@B[Y< 
@')_7LA6+1-\TT%9TQ9L]C^\)P;DKDG4F(0F;""'0QDX 
@C;IDPGW]>;[-D"Q3>_L.]X@* F9UH4$RH/192]Q$',4 
@=A^^#J("<TG:Y5?\4[E\IZ#L>BI)$_%1%)]NWAOL*<@ 
@LC>PYLVYL$*XN'@\XP@M.*YI]MGEW$;,BCNJ_'NA#ZL 
@9;5/G[[(RXK/;GR%(MGGJZ&)&<](MKFE@=[N)#*!4 D 
@+=P+-*:T '=!_[RX/-A-D7%W4J]Z*5&(C;.;%AB+:%\ 
@+\!!3)"E&T9X^%P:%PF>OE/FC"1.WH_1.FTJ$MSU&,  
@P5S(7!!"V4W"+CCIBA<[:,]J%S_($:G"\%P.2UL+X^  
@A6,X0[YI-SDS5%1H[*#R5,C<9MJ6C$+CNC74N!2A3E0 
@H34T F:;1:_5@1#"ZUV>R;69,]R&K'%@H4DNO[!&^K$ 
@(^"SN"([0LL>!!B0T;0=*_0DX_3O$O\X5'>[1P:*4'< 
@T[#-R'KHNV$6EB[0 =]HDOX'!A']OSZG:OA<.EV%TTH 
@G]Y$I(3V6G*<EZ>H%S57 )YOOV@FMV8#_7&5'#7R/   
@8DK14R!3TX/QDD]GR^Q0.0F10\/!K E%3>/S.PJIL@\ 
@?!X[ZV#X"$%HH\'1G*B-:<O@:P%2FT8ZZ8K\:8!"WR$ 
@BZN"6]K\:]6\NVTZO,^\XW<Q=$P6/LH1;X\@3#.I!.  
@4WV$!Q>O6Q IY#.&8"2ID\<UTIX*? E0'GRCYLI57DL 
@SA<OZ[5J"%"JMAM#7<)/#WB X)W&7_S0=T<LUEHQGL8 
@EGW@ H82I=64;?4$G%1'^5K/BTD$Z<F8?ILJ.54.$\0 
0&6O*-_ZN;LE-@5@(?YJST   
`pragma protect end_protected
