// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WHp1VLCdFgBbszOBL4ZUJ3YjqM7h3YRdFIQj2FS7qJgs3tqzoVuJ3uhKRQzb8Fw5
R1Vc/cn03K2DG35t3pveGMIbDhZiRYg0K+DVvgRwFsvhbQ3Ku5wMfndjH4Uy37E5
dtEWFlZuzgURsQRw07iwCxbjNay5FTIKUgadvD4/1tg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 91264)
sKFJVN1yb26Ma7VblXXum4wUVvF8FniKmYZ6SR1bpg0ZVNkmrTxkQczVqXrajeE2
acf5jk2OT/U7ZtgUZFspaAZuqwhEoCUIngRgAu1jLjgzqmTIHIq8ZhuIRkQfjxMx
fSMjXLwwTgtLt7YY6+/PCWLETAuBtPMOP+nqtdYyFrp2NvzMxkOZexIz36g1CkpK
AzjLWmOBPMoX1vUQ3twhGWztWXRHo9xQ9rW1P6cajWkX/DXKSZwoFuKF89AvYUIr
LpBsXyhIMx5CO6z5l1TZ7XCpyHRjnXVxyq1JyDOJJCx7+ABnSv9LS6R/9z4PAaL5
CMMhbrlaRv0+egsGq2ME/R/kgCCETPra6gMDg5pHPXuH+aYV4yckbP5thUnsCVfA
8lnig+5A+J5inNnRWlJIRK7r4FJqourmkNkKTYzvxojGCFc8HcwDv2RFsVkFY4Eq
PO+OBB7GMbFiJmyhE9l3xxN6XtXN8wlB6FQRd/C+4WiTvkPH34Ww14c6VOhood2k
ngxPMJviGJkSg+X84Sash+hoVa1ESS91rl1oJ0RwZ6qAB7byfHjMI22gkh4iqgAm
v0r0238A2t6D9vIk0idZyYcdlDlvvzpjyXFnk+ChXuZrzrubrUgIoLIXEiNEYqyR
9HQ6g7BQZpuYpR5Srw7z4prHqOTDF1qUBAC93PxPvBmlXLbnPJRiPdF6lQzbh4uM
azz0unZWmSJXJ/fKagusydiBIrIPSA20RRGawVxEelyiYoTAbrIymo+K0kAZO5Ai
trTsFmh0z2NC7xav65jC6NiwmU5jpSHQ65wKhwh+gtlN6+QW1U56VfieIJQVCkmB
7VrWGyQyL0XCIrh4ayeHFn1ZXOpfJdNWGK/gj9rjMQdJPUAxkHCF/bycTyTwmULm
btd7MrgdCFS8zgzEEnGlGUfrNb5Yl79nsYD5OU65QoTgDlcT2ZTtpQdUk9n2P9I6
BfuneRhoY/rQLJoMb++RO1raat9avxQDA7qfoniYlm9XDoM/X+kL8VxkzX0tJK4g
a2o5n1veIVgcMz+eM/CjkmE0pXtxwCsjKtYVuOymK7PWrOEBrkUIQkAf2enar7+G
rKdh0Xctl0DYmWo05yN6hed1OZr+TJB4oKwAjwezRDgIIVUDKeLrc3xIwbaMBFKK
Z9/jwj8QLyEmKdkKnUgYPONSbUqco4PLS6RSBFYjbx2RKzjcuHufemDtKhXx2wZa
LDS6sgQ4kneezOdnHdNluQ5fUAZWAU/rGthNvLADNUbmRLD8abmP6S9nFCmAXIu1
5Fi1LRxDPEs1Tf4+0A9YuUJgdPKn7atR/iaVpsIWytdcrfvFB61lYCjzW+uD2D1H
gRFrNjUVuyIS8Lqbsy0NECXCJak5Ftocf4v1HaJBtb6NCmLEU14ftEUmUTmpsR3k
hJmAexSCkYSLYh6lcyK9fUqFLS1EuB/eKsLcS7GGMDL/kaQf/X0vGuYoFNQ8J9Eo
lqpNJuZTcgRIYxGXWndoTwohH+5fypunbzrIvBHt5cSpt3xt59uvHt2PJkqhT7xp
K6rpyIv/bSf0eJLv2p1/QdBrmaw1iMziW+IjSayKiykxBYPkUTVuq3n5cDaRJ/K7
I6VYbvBL90VursWhtQiGyXB/4XYJCt3rzVoqJJ65vX9wXgxJaK1CxFGENzk+OsyM
47niq0jBuHlKgY0qcKaX0c9qIrAoUGCM7WW5afamfRDwS9CQjGmN2Ct+91AXub1I
NRKhV/AdPXd/nJEkl/mq1sHmJy8My59pH8XzqJPvZ2iS/s2JB+mEbbTjObQeXW12
2CzlcW807sipVQdOrRKkHwAQvrMYOXIG5/2Go+XRp3ARnuVed0VuCqB9INAbwzTu
1mqLXxEhW1F2lFMMefqWe15MVuf3mpxgGtPa1vSRduSPemvzku5ysfBWLJKoL97Z
oWlHlXQgK4NxDUpNO+XtSdxSgp9IbLUDAxYRPG6q+46sQLkbHYQWyNVdzpJM2TU3
fsIpP0SUfDissqYOBnQxAFJ/gRNrF0Qqlpld2lzOZ6ePkR5J3Bu65Uuz2t83yEAm
RNxAOedjdUNFA+PYyczDIyMI6yPsvnMMlOt2VRrHw8L2k9tV8AUwIqpWu/vKMVoL
pTxLSAEyPXfPeTVlR3YXdjUbUTFjHtb1CrYsuwdztwuE/iBO9qPqlgM6USLqTTjQ
E82uR2KkR2ZR0a6w8+3xLEj8IThoqLH+kxsbDs9w1H+svPXIXtknxql4RlGXX+5E
wftvyX3oted/95aAztvmaz9bbzZMmaAQBM4fs3+tRmb5kv8gqBTJNVMOwFk9RkQw
LF0qhD+LOX/ga8JvDQvTljsqvA2uxrd1RQXKkfItqd48l3S2LNt39Os/hJaYux8n
KF+4bzGKt66QjebmiFi3xp60ffJRbXbN/Qu9stDLwbmiN31jJcRXs+j9AAvWu0hy
GEET6qQAu8uahLxqj+32NpjA6Ikbv6yKMKMEu11JX1rXO2PUP9qo5WkvjYVch+Bz
KsYTDiymmeTwiwoSYzsrISp6dHVkMQNV8GyEhwT8VowjOK9WwhdOTQxHGQn5ScbI
edYI83DVaSfewfZu2cqbnnKmAVmH+j/Fn3ZNS0S8eEdazQP1bcuop7P711Cean2x
pr0D4/FouFJ19QeSbKq606MhoZpF48oLO5+tBo48ITASkENW69+7/JoAGT/2A3hB
ZFGoQ/0+F23cjG73eyynFNFL1QTQvd+yA+ua87sb5e4M/K0sK8jaj3yimHIK4CHz
cfCQ3RZmwNSWgFJ9ZVZQ+6tKaccV9NPKb2cX64HQd6fLjA9mn+m3u/3TB2P5G9S8
C8qfddW7IUDFuBZ9z2NqbpObVGka0zmfiFFcEE25oJUbNfegj6BBeaB9a5/gHDJf
e2oPpneRRCkY17goEFSExfGePZkl/0yT7ANdnjNHbcIt84NxLUjyZbiDDPOlmOX3
bP3Szv7LQfSc3wlRrxwllBV7hFZPvO1m1BPq0tNeNfgs48NPEci2bxJlmEuyv74+
OCefEPFolrFYtczmLfYd8yI94I6b/v41CJHxh4pEvm3ycuOFT+07BaczYsKTIS8y
bXyzHWYOosogDpOXlrxqCBhcnuGEaIwnX87R7Bdr8PRrk8ppCRY62ryF6VQg3Tqh
Tr3GT+NRW8rontsEhGwIOeKKC9WQmh4ETKb2H/Lx0Q5p/m1+uZ+Gv3T6RmL81jHk
mHrvBpvdIWwkKd5pzRwR250ukKNa22g3NzaXUZlOMcqo/T152lgmg8bGoPEYPotv
WF67o3/sTgBEGsa9XcSnQs8IqboH8oVWzE0PEDcqmea43RssSIuWMwwOZfY4tLo7
cTutmRsC9RHnNjaWI+K7YJxuYMQmqWbWeCWQeDr5I4jivEsuDgDudvOspaFRXZMb
/+Vt/uY19t2BQ2Yqmb9/PBSOYO49I5Re8lHsJrS1aLX3i0IGW9GDd4gglhXVIlMj
ziM64ccoaehElQ7Ta/ENnnyik7zhnTEk9B4P+N09Cj7JTkZhLQQ9phjFY7wXSQvN
+vfSZMzn2jgdKk/YhYUlB12AXxbro1tqGAm29Wz2DsZbcDW9aN7qD0uly122DfEa
ICA9Li7547Dwdl+W8Vb1cY7dObA0osspfeNADBCSPw6tklyf2fOIJSUluq5p87T8
kZbgSHrAaA7O4cqxtLDhUfzpk45zA4dHqAKLUvbWhb6xQcItM8XKBz+dd9sEui1V
yt8WfWCbT6Qp9o9Rz9tHpEqHmz5Cklx7rNvDp5KtqDK+yU1vWSHvvG8BPd2opTYS
O9bK1Y1Eclae4m6+1NURz3dBswpRJ1HMH1hrOEhJ1o7SoNPHJQylbM4rb6Te3l9W
ZqPX9cNqK/deTPsfbaaqn5LDfio8jtCNA+eIwg1JXoABl+KVwXfsFUERmC4s7KAZ
Hwc9E51eXI3jSYCyQCoMlH+OyDxXVzfeoYniSFfsZZZDuULvjc6p+Haw5Wf+WCCH
PXeDTinlSuWzDW3fBFZLyrdp4ZpPebsD612V/9Nh3IwWnrXCfaQ5Lyc8AjFKVmU9
nWZwJSnzZ7pQMunKEgX93EKiS4nsbXtIOIoWohQ9FW16GDxHZ8vgeeOtVTs7PnY0
JOxiNT+LTPpJn+GCMu7VNrU7pj/wfnAIgN198AWySsMBdLSnVnbhf6o486AFtE9Y
sqGFu6rQYCFGFvR04LCAugznNAhJsdb31zciziR2kcHu00JaBNs+iRJDgS/NhSIE
xV5Ud5GN/fv7VLgW6OZzOmY5Dn2zcmuvGeXZymdDfbPRFreWpWBbuViMbt0+UIgE
9+YF3SDluO7fZmvXl7/g/V9Zt2LjBYIYwuDhr32Phm7/usUlFwd66k1gzSY9iRlF
uJOrg5n7+UH/xHUS7qVixlzpVzlv1E9HC9b4FKN9eNjQEcj6UcB2frDmHM59vz83
n4RGh/PWfiiQpmaPuGedMhv8Yyin5fqj8Gg4eTgDVrUXEQKqweupD7QI/yFKllkU
rPHgw8LDN369mUCjXH2Riui0wNWUxf1eORRUOe6pj5vryD1J0RfA80/Sc764gThf
AVpcSk1dfZl0CKmxRO1VlLtaS9ea2nMEFMQGbA97rTz5nMEQ5K65+CNP0gvSRO4p
lrEIsOA3nD9LP2rG8Ni90e/dW6K3fDuFkmGCSPeddalfp4/6XbyhZ+6D4LJuadsb
ilinVo+d6Hqoi3sih8bxb683tVhRArkxteK57HRAa5nNJIj9E7x2biyO1/IVvVZU
XtngVc+b5FwdfWqJwSBQK+r2TEI51Xvgn4QHn2OjZfGNV5ira9MdHsdw9Y6ayxvA
n9B2QmIWNftdhLF2YNWUKf4IStp8+7H0yhYrDX0xOTPRwzQEjkMuVKVD2CnXhHzi
DeVP7DIMm6+iR3c32glR3k7t+skY+4PebUxriTY5iaJifbLxCocBvQTZqcIjdGBx
JGaTUby/hxfc8jUy2BRzQG7PSrpvj/uNHX+BQ6XOvmOZg7ngTj15fNjTTc1mCSwC
QP5JOOCj3+Zl6n6DL2ul19qEthNxB7B0RKlsZs8qByKUcNvtaDg5hmVygPOC+O1G
iD17Gv1esJeIarqz9Ur+H0RzGiyJQ49aaj7FY1/Ed45C7faawpoUoe3WrVelPMg6
H5j5GfoSalTN68S5RlcLkIJw9ETzpexjxUu7iXU/cO5/SXwXfN157MgMs1k44PpV
lCrC6VLpfm1q1hqc7aSCf0UaNIBaCbD2uNhcG2tuGFzZrvcXWdARr8t8YrE2btBY
66l7N/f72zgoKmt0pBaeEZ0hcI7w0qcdUaUJ8wDViBoxDqh1f8G1Dvkgqk6PAOtj
bErvHTGDmWcc+B1IvVtu0SZRy/0WG98h94PeUwHadXkXXu5wNi8++t+vUSkUMj7v
6DwwHGrKmYsraCOHWxSFyaG/SRiSxSSJCQTeUVqE9tkiv40bI2USHGtfdEVTq6Pm
SdF/0Tx4P0niZKKKWw/0Ycbjpq7AwJqT0CuQF9EadeKJOVxLqtsnrgMmkGGmyls7
X7RT/repNoZbXqPu9jDiBWRCCuB8g94Noc5FyuvPgaJDmg0VbGHzuwTUPylrwX0P
r0fcd3Ph46oGNfoNo9kDP4Pf1wOyY8z3maZl8+U9FABeLeTMHiQ6akBY3DW+Nac/
crITPVgMixijx+4UsA56FRVPAX+q0cW215k+x5lA4WtDfX8137aSAXR2iEpxGKYM
hnYkFO7acnl2kEoAa1VSeNvyE+/j24o0Qljc7GiQDmE9ldaXxDwJsuYjeX8KrVJj
i6FbNomWUaggQ9t7DVVU3lLwPUZsnWH7h8Pe//xGgyIqkqlR1VSRRtuOgcOD1Ox7
xQSrLyldle4bPEVix+KTsZe3XjUBbcUqW8SC9P2FDypLmi0Lqm40heoxBjPqfPMk
2KECbLA6n/oGGJ1xDXqGVCfDy8N4nukCZJyJIQpSGcgyrFZ5O8YFL1+8U85zj6Jn
ErXnA19gPFc34FMjRsb89XHRF9+h1eLarwRE1/bDZ0zN/ZTFxR1TrjmaxB8MJnlz
YPaqR8sBd1aTIerTGup0cNUVcLB3SASQWhjColHVEcsdr0X59oOvVHWY1X8wADNW
I4OWFB6sXk1dmW5WVzsM2N7xmkNf9nJWCR4BOxksu09ZJJ4qKnwCyQKNUHfZWH9B
YgC6YEtRZpKTfAh0yrSrZlyk6G88Sx2AkQBwxHR4CX4Eb8PVhNsWzhd3P2kOMXFL
dHkeBXqw+Mc8Hjb94LyhwcR9xh+TiVwa4pgoUfNPfh4jfkrNf+2FasbDmjeg8S52
jdzvif5p82OBGY4f301sMuSNoehM1W94bm+1K9FEu2wNEdSw+5JgmRIyJwCMHs5o
gtATw5/I1Fyi22UnNVxjrvV+bv8qsUfrouMDxjjxEaqJ7QX26J7eZhOiGipQO0af
1pBvKH4wkauDzAhPIxJhdETgPIFgWlJshowBSWzwIlnWtNbES2fRyZkoWCXf8jR1
3SG8vSdSfRbURS535U6LU3U76x7Nqic97Ge1+uSEEmvRsszO1//ceBa64VvTZ1Z7
mZd0bKnbfmRsiYIEO/uPXjzkLcLoTeWgZ+IYwJKI/y32QhCvIVhSJW2Mncb0LFl2
zjQyBS2UfKmJbZbBEHzBYCUKYWaUDps5ukV+5dR+Ep/CsvuzOgkNQsZfvZKIH0TJ
Nj3dc4ZnMEm9Z8eMI7SdqxlA6XqVe2DpLJzCzb2l0FVoyH0LqEFv2k5dCbXcd3lJ
PGjsgWR4VMip69qtAlJT3zhzhu87uBQjlYHyU0whAV/oT5p0vS6w+1uXy4TzuTIQ
3HkhpVj0VoKquXRmnzzOExKUEzpTJmxF+bKahK0YLwns2B+yi5ujZiSq9gsu5f9J
FMI40rVJJUk5sOOGxHhYqaWCkkr/m7HCkh62ng7jzhuxhwuz1aUJscnKi3mGER00
bhUVo3wqWUwuxsgSXobJxBl7YayD+FpVt9n/acmMmbq+kuX4vpBR4IrUF3ku2TH0
MRugJ88zHjP1Dh3BoURWfhrE/uFj2jM6lXnmJME5ei/Mbkw2KuCwXviTIjPE5fZQ
zSIoxPKAmWuKC7i1Xsnpgx61/JFJbnL1bi9Yne/2VwWlRMXRkt9woO/Z7ux5VxiQ
GcNhyR/YkRNlOWW6uBupK21ecajdqaoJMimbGEXsXuwD+/PJ1hHJwTbx60/08KzH
lKo/wofaJjbJU6R9en+p6O9oupbQ7Ltd9Nd3mR0ZhVV6VNQblT58c7HgHZ3YmzKq
hpJ2ANEvg2w3DcW3VFcRspu2JSWrUuDCdUJY4X2tJxPhJOU4f47KzZKzbSyzWKxM
H3XlH1GOA66Evjk5mwD9gBlptThQPZueNxSDbuQh64q1PCKOq/q0zscem+lZczUq
ppmcUtiC4vhxkdtjOOQPyzRTHi6UK/bCtKQ1YtAr0MZ3mnwjPjAvk4OUXLh4k9mv
2uEjYoXu42C5SUBD39s55fQ0KV8iWDUSCm8njYk6eNMR53BvqHp01j6cdoDktIU6
ex/7JkhmhvUvGNVAwQcPepYn3jkAoR+6fUHgPrjRdwiCna+5lE//UFhvrPEt85HY
7AfYurpZEc9p8HJci1L5Ux20XiFy1FZQHREAA/f7GEVjUeL03yo72gCWnNUt+llq
rR9fjfVMDQCvZukHcFp5O/6aVa6ETkpDuXcXRNQtxYqAQx8Rk2R2ptYJs1SurFoL
0JSL0QALN7LYlr0CF8REKQJOVtoNFWiqEnmXffWTnO+9YX1XcY0p7gl+Sc87rIlh
kEPs6/OjVbu2D5h6uQr2gmThvUc/IBELN+hFTt4RHW65TpA79HnriRvfBdRBHs7n
8F9nZ9LPqXY7HSb0o+qe5XASB1KXrGcGRNelb/1dUbENmODuu7yhkOixMZI18Rlv
4kaDtrKBPPhiHqgkHkwDTNofwxnu0lSfnuG4Hdt/BdDdhlyW6ci23RihpcnfIBwR
PT2/W5uA3TQsxgloAISvCgO5ZUcP0mp46kcCFHtR/nSOsnV3OgBYw4if+kl71o3N
yVdcenSLsOgIbFq+XtjhEU4f5TsI5BX+6THPL06IQi3RJ5O70UQFB8X2JlWjyLXl
FdCBv2r3+w8LPUm7vi4mUPo3gwy25TTNbPxOtZ9+IqtP6btuVApN3fklaobrIjnL
0fzcPfAc8SECxbUhasORzw9zlxfOinuFaloMYVV32OaUkSDVRkYLLWtnhIABeliB
0j3nBT2PZyuZ4KuDqmm4ROLgisg6wXFaGM8GtC3C2pFLIA+KbuqG+M5s7uACCSmS
7WlA166Mzbb1H4wx1ujMpVmtvVdpYm7X87duNeDxHCshBhDHGxfCwmL2ERUzIaUQ
WESj40E6fnM3/hcNR6F09g+tTBT7iK1s3syc0cn8IW30Do9wVpuwdsDsNLnNIEdd
Tzgh9cvE1X8UJKqkw0scO1Oy2XdxwkW8ViJ956Wy5AcAyDcvzz42Y2aSGRh+erNb
zRXwFxtdgHa/hcAcMzUls52MD2owwePxLDEwhogLWarZ6nTiP7tNI4qaVZ/AqoFE
sUbiGb0+vdFdF5JmMhNU/kv+a3dTzNTWPKMI/XcjSWay2xL2q41/s6F/rKEuoJBD
y0ZGVgQ/RWo74Fj0WINzl7Dk8yq454LUY8M+jKiMp5jBAJriP3QwCoonRMwwUh+6
C96LlCUuUnh948s1SYXhj3Koad63JNJklSj728wGuPdrmxGvfJq6YMwVrn59gM1d
mKQd6wZConv3AtXg6OQibI+FAEWJmTD2X2iOgY0qEKQOYKjNDhWcSfozAr8HOLFX
rJqz8OAqwS2KYkiIRUG+mMuVInv3koy+Qxm+MWaMnEUML4SV05WI8QLLWCI9MgSt
8t8zP2xhPiaV4JBLv4A8c4l3SPa16p/a5+o+nsyT/AguRvNkFsB4f0QsshrvLKDv
wgGchGbQxHYj6v+SyCM8w5QtC3DnR/tBt3u2TI0F+RmD29GdvQ+LMFGGzsqnQSZW
IGbsVbcgPpFB/FWFR8NjQC5uQrgiPXy6oX/rRYxS0JhVehW/Zohuk09bjpj0Xri8
jqPyp6pW15N4VvUnKvmdUvt791Wll9RkgEk6YInTQYJbkuXo/J4/sV7GQhnn06YN
t/0Q8RGWrRhGhtl18mJdJcXck2ThNm01Hsd7gRPvd9QlvwcGyRZb6JHBU0DBrZ9r
ym8PF7B/rZSIAfWgWXP0y1J5ji9SSurge2KA2lZrXv/3fXkvqLqoRR6yT+sERioL
eljXB64Mmj3CyA0PhQPQTDA7KRQzz8xPLxKRAN63FvnCBZ9PuSALc6ACbj/vl+zA
Rh0XnzqevFTxlynixUTw1JdENiMARNq1fYEwt/VM3YBdgyShfVuLlKGNUCqJOZbP
/YwLILMWZIO4HTugmgPwpjoGRSDRiTFAPj/t9LPP1A/Yk8jvyG2QGZZr3LBs1M5C
MO4u0+OzkzJvM4QG7WtWM5fFRSFgnCz1cMC9d7VdiPIJY6QMg+M2POMZuhGxI6sx
Um44pt7c4N7cWtR53U2m3o2EN0TCvjuxPD9qpZkR9qyNNkAXCAnVXcrqZMaM575d
eJtBgGgDn7aVoTdTZ2iBXEqmTu3ckk8uLPPCArd3HWrvZg1dv8XW9U0b55Pk3bAf
oblzRgFzmO0O4KV9b0UVpZkjQ6bq4US+wIvGl9vHCGZVSUmryZZWGoXpWHqb+2/Q
Op6VIeEyO8jr4qKBaWAK3Phl2llPyAxRzJlsKJTXY1C3o/QBGB1FA9D5XzxUdaP2
GeIxmhllyB0TTccVCKpcvPA5giaNm5C4Ixk1TnbWDDLK0iu9VCWDt3P+02yxHqwd
3+0bKWLkthfsxLfAtDa8nAsoQGiY0jzMLSyxhUD2bgn6slVpfAS1qfTmRUdZ68+g
YkorpbzHiPzKeGrxbaa8/LQxddIPhE4r9KCzhl71koIvwMKpJRFqLz4gweBGi4vy
EV/0DeDnsv3fymQSPydZ4aKs7D9YkPsn57nYrozI6lOrc3K74aiw5G1IYk++LWMO
N23rXSp4pSm8QTQP4oHIgRkunC5BfQsqmW914sJlzulsbZbAv7oyKXCLmFA4AqnE
JvP0nenBpIYYI9DDq3ivL+FIl9Xq7RjOTfpa9UvSs7d3eF+g5xYAtiXaDKmSbRfN
3N4cXcvGkc96h7zArcr6lFNY07zFEEN0TmGq4WIDZsP6HyqpEuOq3sJMVQjZI7tJ
/Ou/avLKEDQ1DMYmvEZcISL9L5Xy7vc0b4VTOt1rdH3mrlSG8xs3wsRmBzFmPlt5
inB6AOR2UawoiZAvUSdgb2c7MkjZqUmkZeyZ/ohr42NKk4t1PpYmqvA7g0PYiwks
idyX8116INM8NLEuEUB3oPeWbBZju7txdbVCARxQx86Pi3q7pHe7jsMI5Gd51+f0
B2OnpzVP5jdAKR6ErtxIO+SB8dTuWWhUcGTNNs6bR6SAV1pXSUbql3N2VYvT23u8
JRZWgNHt1EwkElBaiYdDliTrzPtIMTfbVk/dKTAt4s/n6LlZDbu5ZqsEFvWbymxW
O4kFS/QQwjYaCFortnC2mBFM61n+HSRhhC4UaSevm4n45QhvFENTMcJ41EpDZk+8
NOjh27MploARbF6FPNYJvTiVPsySuy3RKl8356sPa7glCEOylb1eR7e6HaHIsQbd
FOzsqS2UQR/JoFdaj27s9Q18A8NG5BfwrooBPiKTT+bOliJDgRxO0p3fyKVDt5iG
IPkgMq8GuQZxbqrFUQL+xKZCdksMX0eR+O72piDMdh9iFrXFj4JTLE/Y20pMBkEJ
XB8aYKSfr6pZfxol/DTFtXli8JibNizRGTV/nIMIB0x97/8GP/R/+UEs1htaPAdT
SVzAt5qGEHZWHzLhkvkz3IyvVVq6i1VLCsUWBMUXM0S4/85m2GpKaI1yJ4RI+vB+
MOKkKt+yRlQnWso2kGQfb0JZplizA/W5TqaDSY9vO+hE0tTLnoGme1oVmgeVYxop
jRpmvdKEmPoi6nIoAoUwcc9YQJLdK+XdXYKxFbQLDnmBjGp4q4pMOyvbPiR2+cZa
+t0oxc9hhPvCyjYNHUSrOi/mAWElmlUQL2VLZsFI9nHJ0ZhFdqOsUcUiLYwwJd6S
lv8tO+b3zXJ3n/IXUyxHP86788qkZ6/d5YS4Fl8U4euMDoQOYxpS5UH11d59g2Ry
hK8+0n3pV4FC5ha3TQMZ3wp9ZrrX6xp663b2fQFr0Io2smPnHc0v/m5DhUDNYTIm
l6/3sQxbKPqWzK9mCwk4BrrvtWq/z2fVwfuMb+tpQO3jr4w9J6OY605pFBnJQD6l
lTL5sedN2JkObGkj6jMogD21Pb0YZ4XNdjN4oIYSH8iGTsy4XWEFI4O0xPtQfRj4
/RvEadZ2ud8ac4xHVoGK1aD/GZvm5KsFSfBPzuKFzauubw9LrF4reYGfbXwymQGQ
w1aIAFBkq2kC3FS1eWxhulkaMf29PRmL2vaFnoxZHvX/QSI//ZS43ESBNpBb/L0t
WudM8sDVRRwu3OfqEi2q3XDnv7LW5o2mtPCEa0dfrgeYehWIq4eDZOxA+oTbyqRB
EcNYv750c4/O9PSMJOPgl+O5TautXaML61h1f31M6NnEuJc52jY0mruF7aszd0PF
UyQMhrBAcT1Bhz72/kGUVOY2PkeoixirwOoz3M84UJFYRGRsJi5lx7dln5yWoq1W
mpB88JHAr4orUvirles7co32pVDn9nhIXfU82CvsbOIUlrRIPusLwFzqi1FXaoyf
h31E2qFtAQR5m1aYwWJw6ZKnCZtc1xfNji9UIclcfGTr0E8nXhxt6kABElv9MQzL
Mc8XdFf0MA9K248hOM8AmgNo2RbAyv2bXJnKWj1mW9hYrS9B2w53WIQ+Hms+HU1J
rj0/Bq32kW1Wxc4USoBGzBesdmplA4TrecaggEf8HkuV98x1gAtuS6n+IwNRmNWN
1AY815qzOl468PfZzTEaEoujdcFeEc+8oErYhjHu1pTf7qpAL8wT9AuSUOozxfw8
5RkR7ukdMBZLTuXDxp2Fuf+m9i3nD8/qGw5xvEV5SP8S5Bk/Z0vjLbf8q0+ztpTC
H6IPNi9J+zhYtlPRqahtez+CFxcIWjs/tMZ0mmKllZaMRxM6vX/k5WQdNLJm0A/K
dHXLGNJsvE9zfjpkOhhKC8ryOUy673sg0zl4h8NKlB2Rjd43vX4aNjntmqCqUrVJ
qRbwKJSTEnO5/9UXoXi7XlmIWGPFpZPXZ7oTOrkalp2UDq5YLVbjTBXgOqJVHIRW
IXO/Ez9baIWAWeZKSJJmAgClewLIOfsSO0YNLKwiw0s9Io5YIc69swc0x5EV7zsr
HJAY12XzUnkjjgnfBK1mnlLw1nxR7x5GDD4rUR0vztavUpfHv8XF58osTmSH3ej4
ThED5RAF5leNvdiJV1nFccPCqUSVgIUShTv3nt11Gy7WrhUzhdQMt9YR2HM52uKa
TDrD30Xzo93AmYHp/KVlOLSaC07uyvxErBNrL3i7ysB58wMKAOYJRJhJIEMbb1rY
NvFp5WQmFFeFkjcy4moVPykgxjk/i4rhbKl7U8Ve1tRk4OQ/TbDmpPfv3MLipNoy
rXunbu8/98PY96qFq/8K4jD/vovBgm7kGTjV3ZFU09LiFYgBhcIZert4lbCuYD2A
8ChS5uKxhT5y2fVg7MyU7s/RG7PRdSCyP+zK3vko4kvLnQbUVy29tF5ExU8ozVBX
/8qF6P3p9gijp3EIo3bxPLMs2ECgQaCsxPsEBL0QvAeg7DsIZ2wVDLhRxgYxeNKl
vYITTVgLL/cVfNR4HSImW7GB7s6wjTTfDwPQLNpsm84jOoCKikfQtlGqC8cBhcui
+xwPaCop+j+Tt7FQA226xUwNenEhunORvWNgEiyHblLk3GfPwnRrXdvBkWs7SZDh
dqatjckPZvsnT/2WVNHaO9Z47qj9CxL8a2+0BDLdIR8PwhGPn9fac31NYEzZPFTd
bFWS0782a8Xau27K0Psq+6IaXUlTEmIHTdy5E2UAeGGHTuZxY1wvOW1JC+mpqsgZ
tVNsN5q3XAtelwCyxYgE1ND4T57k/WRylHTFB+Q16w00OyJeiz3LIdvD19U1R6x2
Z2F1izc9wQmHkddODUNflbHhd10SF6eWZz51Re6kS2AGyxHAxLxZtd2xL4biazf1
qGgZlZ7VxFXY6TTeUKCm5Av0ZoUUBHrV3vL46PWlxZGQWq5MiS7nXMLPIoSr+JYl
VfVEzpQXUHTzfBlfN7mE/Xnqi/ZQuWzhTa4ylz4IB2VzrS1A7D1W/6XtXhpwXr3o
xk+1bSF9rYQP50I0sV80iZhhgp9H4PE3GF5Adq3vuqlr0EI9pVxKMgwHoFHUCEA2
9X0VRg0zzy6ti2gO24B+pQd+LCmjmrspabM9a92eKYKHDCiLOQDGyCmHblny6gq4
/4Otug1voV7SEa3BR4lEzS9Qxc8qHm5LnjZIFROmBD7VHhbrODP2Z7GraLAiCV2x
KUrl5nnXbOxBgkBNWDhY6AI7AaKP7i1XNyOMunuWOBjobLWktWGk0dnR4WVsac7L
c8+ECb7sBqET8KXIu/dmbEGW8pzpj/Xj+c3K+M2wMQJ1WZxeeytOXbhHhSBZwxjw
z6wPm8gIcNUFJ9462LFXklnIJXbH1dmWgIzUvT32KY4WNp5HektXg8w0ndv2yyT+
WOgRMkh6di+Jl88+O536kSyVmHA7ieuQbrec8Q+O2bT6lI8cOxdJu6uL+yDzJ/UW
xwqZbT1G9sj2ExssDfJ0qZ35Uz7N8ZvaDYj7FMoWpE/xl+SotqmqCGGpiXMooNlf
qtVrx196GF6uCTlBLDxs8Gg1PSWLKVrUWIOqB5HpE7uW5oXj55pZPH/m+uvqIzgE
coMlGm6HULPKUezUSgTmbphLqZuKdsuQxyw3g3P+Mtv7g6dIjOMM+x2fHCFaPCOS
5doEApce57+iQejGhLvF4aXELCbsqFH+AiAwiA4pyFbfBOHGe6RQkwDZXz8eyxay
ACSRvmk2MQe3dUdvstt8yq9m0XxSTCBnVKyich0Tgi9qgrGZ/iPLZmx+rEnwwUJ6
pTm7BOwl7n9Y+roKCJj8VWJUkVP4MV9czC09Xpw+M/BPTpqDQPJmUe3R1TIT4k8A
f0WNU1cxhjkmhj9aI8/Ey6dnq1BUR4Gbsr91I/N0v6EuFzNmYT25PaIvKCntQm44
49UPgXx2i1ib2ikexy8geZ+aAKe2/CaXbidV2+8VMPHA02spmTWNvh9TFXH+rsmW
5MGe46CJ5FvvgTj//Sv/f9UnhHnufrdZKK2Lniw8DNXVLwl7WCk8os74EPw9xrgU
imWIdYEos1TR6ZFC4OcFpz/qvwBr1tPSU396lwgHiZ+rzUTGZ8ZMeiBOHwQnKE2T
EtFMVZZ9AS/3GFdSh84Forp6s/+vm3JARQpg2b7E331pF+h7xB7vIAM8uy3/wGv+
jqk1j2UpofBXqMftTm7zyzI2T3kyihEM3lFef/Tf/nQglPIXH1xZxeHJl6+c0v6R
G2kcmr6vqERTxA2ufdFRQfCXkgWTMftHoSSWqlLb4VrNsTwTra9CougTy+wTtbJd
kF05DxmZvrIEakSGwHPzqStTIKNYZ3bfJHYUJY9EutXvKBDOZz6gLgnokTJaMOeY
yUETd2sOoICQDI+AOyFkW9/ffU1OcbqaW5VbFNPT5uB5EzXeTFK8m34NrMK1CErf
D0llpJUWigwwD0c1B9OisTaTdww+vjkDr605HA058E98Re1TlvlZkXHiEC7SwuCd
0yy2qwTmr9LNZIvGFUCzp9W/WyiNSE03+9hx2F24eQoyZjMh489k0sWc4vpBr3/D
l6U98qecFwzP4sZ9nWDlGPF4+BPocsPGm+mw3LOepIYMPioX3rByBr4C4mrYE8UY
Q/xgO4BbnzkcpTNW4oPqBCTJ4pmxsBck9VZ9oHKxy9Yl58ZGDm7SpAUH1DmfDGnm
DLjMsxFBj9ulYqg4KJ4Q8aCz2kF96s3Hft9erGoKXQfQGVLOkBDTpSW0jBOLTuha
YurgAoCCuMIVUPJRkR2XZ/2edgMUgQocxItL67eCUv98ANmMlp/6qOzj5Y9+FPns
DCO1HY4p09hibe2o2WWTDwSnamZXKm2VV0A9/hGFV5pV2fhEI6BoJA41Sm04TjMA
xvfWHJVFfGCw0IVRLVViXoSEa6SWRZxquI3M6X7ZTC7BewzcxA6zodskTaIiLwCn
fICixgRdOjviICIM2643KWd+Lr0a4e4/AfB2Rw2TBYu+pcc1Gj92f/GnOfgk7lOC
cK9Xn1KIGiqVfBb3WdNbZRyHKipLbvow0IXZLIc6xd4l7kEaZqSFeLM4AAQtVu8r
phaJa4E1HDis6LY8tKRPqorEhob7xzFrvvJAX09a5Z4cTOQ2oDoEVucpU+KvCWTS
1eW7WhoamBcNdnMWDFU+Az7n71ypDLDWwbjvWzpla772L1CXLoX6B3UmjakfAzyh
OZv5BNk3eSLgZkmqesw4lXvcfjw/pLTCWxM0Dced0dAC+jXI+lLi1xYrGHmVyIu8
53m7ogf1b/eV4h63S+6R6znOZXAdQ1lilH+w45FpTma9sCEntdwdpOcH7shdHLvo
qJo+qYC6fALXLh8wrZ7hQhge4yV/k5JlLxmyjlf81/vh438yPmQtCY3fSifRkl1G
Gig3Ser9jXX2kDwee18pv1UuY3bfNeF2+UM4Cv2ZXswNM4yqoOPm28LNXSeDAkwK
DpKwTv7mIscQaMOu9bzYLeOlq6msKXcQLtav6KPNqTbHhaqLM4lA9HfykHRZ8uhe
8IIhE6ys16t+CI1yZmNv54Wcwv9MgiX2y3Kv6JWqATkrhZ+x99lwAf+dJ4EGD9P8
EVYTuo0rO2Hxs5Rl6DOsz90Dz/OB2W/5L8eGl1bMazI8KVZgeXsG1//3Smhm6AzD
pQP+3PNnJwroTi2Aszhg/AOtn4mYUWiYBg+uPDwgqWtwTB+9wIAEv93SKz/GB26B
h0w8f9+hkaKwX5AUn7s4lPQH3gC0nhTGLmQtXyAstP0ezIkwl4IvuUALqGtGqboy
qtd7KzDJdQpbHT+BMyshPdbx8NNVimzJh4rit62YTxTilWCHInYQ3k3a4/wSBRFk
ShFxP5V6gO0hVGYIAft2pToX7w3nT4UR+V66QNPRUl6xi9UfWpfAMbC7ZswQDFQY
DSO+37zg4HZQxN74mSYae6r7cVoeS5ztcimmZTGktZ4oXR9oy4dXgrpAWMGLLDni
s5JnAsN44JCwMUP9cJN+o8mZs8AsaTXAT49jm6XZy3mWGJYjdZum/HipP2944VFc
qsMv2feGMjIKUBRhNqyqZzcKRQXxngVncc8eKik15VVNLgtzGa64MnTYRdtF99r8
mKEqu45gntwGd1N3g8fgD6jIsgXb5TyFMSQHVUCb+TUJaW/rNVNj/wQdKnIWormq
mPx2ClC/a3kA87EnIxpy1lTi/0yM6Te9ddF3LpfN/oJChWf3NX8aXpfq76CPhGnw
06xCBZLuHz+A/uDHHeDa6PGZ8Pp9+g1KUJq5JvPIb0sp6MBywqZ+oPOFxzy7GKGM
zn3gmoglMyrh9GJiB8Z4dSHNB4RmBuLWCjcSrv+mVAn9J+lHp04wuKXT2R5i+ta/
e3h4iTPkEQPx4Qif04m36EO+8lYfrzGnwLCSXbiaUxbtOj2/24zjXuyIcExp6LnS
P17e5ieS1L+sVLc99u7ln1jJ5NHiqw+DniUhTquab7IAyaOb/ibrbtjqyfsWuzkZ
OOHJXzcOL4TIqzFxJNN4n9ecfoCZ9b5U5gqP9Q7EaVcBfS7ihkf+y/9GcddCeUwZ
vm5ZHBSo22DEeytYeBIw+1234gQqsB40mr0V5Vq3FMJWUzgBgPHbhHv8o2cTg0I2
gCYPffVQ8O1kfUlj93g+O4xYH1sxpBrFDlLM3FtCaO1t55tLR3yoQGx19a7fUlKo
2MyV9z4kYxxsO66fcgqC+h6Kis9aIad7w5XsRkjed0bdBDi4xHQUQtNVt8Um0l5v
H4mjkpftCbPrIc5n8v2X8oSPGKFe+HoG6kcIUvpRoFriLT73QuVFRzTbZF7V3RNg
hAmzADExOb5tZGipMHE2qP0N9SIp8j1FKIANX2C55wS3LZwUmXK6T9TT6K9efvAJ
qDXyfrwE7Z3HOZ4W2Y3ERqCyBbufsL4yLZfsueXRkDXCiVLMtwZ8Uub70PLckm42
A1rOohAIish5cPlLOmje1bpt+rxDb1wjPAxzhC68lKvVUOmQ5qTLLb3BDzObhlvW
WRsyOShR8WbeOdohsP1HM2iHkMASECvaVJDm2JRMGZHu7v92gZKJxvBnpBH/hks0
6Q9dj3egJbFyrcXFdoV/MMnB50m7LP5xl6bBUp3q1j7jBAUAGbjuDcZVPSexcAue
1jq57T6AyuTTO25Krrglu0o6DQccpurjtFCyRiv5W7s0HnZbtGiMDhYniCXJBZcJ
LMVwzhBH4zXLFhJOR8Y6k6a22sBz57kcMvbjn7zoVk4PghYciUbJCrZvuOcs7XhX
xCf8A++w+NzPYnFoAioa3eYopFefxTfTvflr9d5GQ122h3ddm9vrZHObtBMM59Kj
nul46l18YwFlCNKtkg6z1UQGND1oldRnEeBVwLsSTeCAh7FMI69HD1HP6g1HoBC8
aeBmEt9rskmTGu9mCciLKRSxRW653DAWPu7w4i+ypAkfF5t5TSrB1b9s/8xetseM
78tEo6Qk26wmwJsgxuiUi9ByMLK2WL+L+MxZv6BdPc4ZDC/2PqIJIDyE2zQrWtOz
83JTcD/RirLZHSvXG/lkmdTzexBTPdxtCDucYVX+IA8AG/pLHY5gp4KaTyG2vV8y
HoqiVkmnsqauvMJl9lyjRqBu007OctVjsW2zr/+HgBPb1kgRRQOQmCydwlx7T6Cy
ZS1k8ztkDQTyB6JlX60NOcLTR+EPnQKijcCcxIWkyYj61GPlSqc5OPXz7EKTtwz4
AKXSP1+OSm61LPMFLTh6rfHRb430NtNdOlDljFEGb8QXQrNxKawBChB5hI3fF/8V
ZqnttUC0gqV9Et+Lesqd5HVslb22XpeIooQ4AyperhyFLgwm8u3xJQBm+ZNZSuEH
VHS61vsU5tGedx685KJpc7P4gViIe7gY7YcRKTpmGyzDo2VacB/K0Tm/M6Ov8u3v
DCeLqpLOndwbRMVSJsc1lsNVxFmLwJaBdF9/rM2wlb8ZGPqYT5syw5azmynwPmh0
FRw77snv7hXe9nf84rOgE8LGE/xS+9O/B8jHNqYBFkCYQJ0926Y/TpfCkc0UL/IW
jZCH4AdnBxj2Ft9BRqiz3k2wGrsvZjk5ureMcGbiQt84sSQBVM8MPyGi71zZBD7N
Yjiq06DUqXhkdH4Nwy6j1+y4lVjrU05Dz6dT+AL39qXbmOvQAin4byZrdBUv8NrG
/LePq8tmU35HYNxCHaGak7+kBy/2cr4r2f5A5nicMGJ/795VfoW1v5O4rsjqj9rr
KhJnjPpK8Ctm+uQfuERVTSF5HxEzQ3FF36j9UsAaenF6F2l7p0XqcgvJCd4JI0V3
2R1ee8OkNpU+MRZCxj7AppkWYyUFQXE8c+7vtpWzi50tDsbD8fEGZczRMSArpejh
Bsdjlfvtk3uNSB98DONoyBC856VgwXzUUFXf1ipq60hLDn8Idzdq8bioPY7SkTlc
etke967OJ1iYIWkaMZpBtMSOVR/nW7dkMwIh2+O0SUhT5Dpw0suDdvgJhx0J7luo
mDt9q/Xt736kfalEY5BchPqW2x9WrEQYfsfTZuTVtQK+qW++80hUciWkfNCQfDcc
bt2rX7fCSXjiDE7kBGrgNBZe/3BeJtDADdED/57y1Gfw5NP8x3CR0AEBNxLpcL/y
5WVz6blPNluBlONGfhyZBtT+Nz+jRmoxLoahS+tqrz3/a57lCorqm7WnCsarpo4z
ai1a6cD1Uyb8F8v0Or2f7zv/VKi25iNTIu1r2TEXP2xCE/ISrogOXAEKTj4NmjXr
zpyEaIXwhTlqrz2QKaZK/7NpOx+x/QTov3jgTAyDk3t1OP/peTbzq9jEQbYM3q9y
BIQ5ut5E7ikPmm5SAzoZ4jo2YBvI0B7EFhqNzXr1vQ9xLXKqU9R6Be/JZSvw0xW7
N0ZlWEfmjtfJvIgqLzw+ahbJ0QgfQ1SMsb1tqNU1B1PKhlbTJ+udxJaMTwzMkPDg
9U6RHa8UoE/UgEqFb0vZiPcQJrKfMCeBcvU9EASH/tEvux8aEtNLKRDlnM8NYwEO
IjAmaI+gUJ7pBb510ciuFbJOhrBsb/A5R3dLea4Msb1g7ckPSC0ZSRr+x9kTTh+8
pL3t3tkWEkxgp+uQkFHPdP5nI+8gyXL0ugDP0vPxj+i8AAlwkoPDZmxHnaS37sSU
AHa2VJf8+Ejt8y7teoDAsGxU9JXz54GR80f9z3uxFH6sMlpsjsQEMs8HWSMORyF0
hCeL08SyXGfdbs++bUlBYZxMKg9m0CG/9+/3eAz1d+CZT5KfAx2dD5MNiy5wInHO
eU+UvTFNxemI0yBjPgcxBzN3zV85toe/uZsq2VfGU6v0Tr8LKZqRNXcy//AexEq7
+7KiNHOpXxQSIUHoowI80cazjZ3/bDhoUJCPunPabd/qVcNiOAOJjoiSOWjYA8kF
+Xw9rgdIfOqJ6IoL7zsAcS9j5uQAi4uGOhON8XjTNn/dLc3phUfrGtdDxIeQUkhA
9t56Ukmh943rzsfCW3RLaHEgik6LCMFGJGNEd0ddy1DNF+EFw0PDB+r2xmsZSOzD
g8c2zlR2YpjhBGOglt2WWje68HeY6lMmtBw10IzPgRA6dQRBQSoQdU1PIP080STU
9rEERkFKnqndClFU3B2D8irDFa/dHAaZMAjsR5bdjNcKSvGuIMmRNe8AGTR7A3A/
dqMgst0rBAGB0gsn7rowRdYKcFQcWqaf19eiJhIZeI7v9Mx2o+44llRMYsydIh0Z
q8xW+YGQz44jklvfydM+HHwMCrMpYDeA7mDdyCZHkBO6qW5G9Fa+5q+HNJ9rXmvY
F1dmFG/2fpffaUHbSWslosZnICS02an0oyNiJt5990i2j3ObCXVAy7+5gguEiqiH
R2v4MdcIHG7CIbHF0fFgEArKAPaczGafrmDT3pmVdzA4JtqwEHUEZwFhvuuQKNmq
8p+JDCBJOKhWqyxk06eSVfoLKuK/OIEP944JJGgAyONNbBaw/n3r63nsU0hGJvOD
lPL3xlMnzjcJrequzDv9apHHKkn4hzv18gzyD3yIv6+QumZQ9MM0kfag0+eiuzyA
9NoTMkQ/ZinKZ19zYnr8WOUQFweLkETMgjEN2XfrP15j07RC7fTKE905BXX2NlNy
/T9swppjQor8ekmaw+lHuRXhaO00IIu1B24uOKg+1cdnIBJhrNqCfZGc5tFHQcQh
EUXTPfuBEV3d82dsAjMPhUE8D2DAC3HJP3iQbIA3O7tUEginG4xeBbUNM2lO1z0A
C7JTxvNzxHuMbnMKNz5o1Id+HgD+7PBGN3nrb9sxBHrOJu3MxtA3YD1kWXbSYK7X
+LPP+ZNzEDekBFPn1tSGPBRaaw0RQJbltGqV0GuS7LRxAKzEez0Y25fN+rjxoYwN
MVjJ3P+pgTVfpjXXv7KGWHkK0sp2TWRXHabKuReU14IQKHoFCg0ku4jzlISvPg6K
33q2xOJx80Bp0rN01T1x+tLRR+o9PIVaW8QbUxP4BS2lMT8zIxBtvwq3Ixw3eXNO
SCai77HsqdruORyYHciVHn/us7G2Sa0cv4fKZ1ly6iKDfn7rQ5XdjGe2qep58Q1q
NtkeBDbixVE/WiG0gxEmLc0yknOnqR/QVGv+oMILoSwwrmrNWI7jA7/hwFe1YcJi
ZIirKPnVMdeeYDI7Kmw4mMGg/m1MoJFEDSfnZQmkG4cCmjyjejVSEJHNWzcUlOp3
e7i2o4sZKR4ZWG6vRv/GkduQmPn93VN6GNIDZfvYUHt7dC3LmvkaslSJeHkyM1OL
3+FMGZW86jCBPtu4yKDwGy4adYv39yp9erBhhldc94rwdBcqtWV0lGQKUVr8v18R
nvxuauwWsyBSflC+NeCgra2zNsb5BXebXWc9P/X70NypZjK7fLNynLbgA8au9Jg3
8/g6vhjEXLZl5/nV38Jil8d7s0VluRCklsYhqJnZaCcSGz+xwag8zqVyP4ZRUlEc
ueHsKV+nGcW+zf3BUJpdX5rf9i6ZRjtaFSK0+BxcP2xk7OHrW0mD2ZDt0vrc90Wf
BdE7UyV3PRTf0Xo9XzBnDDL7fqv9keqEuknwc01D4ny/uLM5CzekAhg1EjS44YKl
j3DHJPS4ch8DABtg0yQk505kYY0l2geJuYrFiUcZCWU2OV0hYFZ1V2SFpFT/r2kp
78hexsRKwGlhHh30guGBKD8y61keE45NGqP9raUxnUAgy+Umfad2X9ct2Dlpqa2C
gRG082WM4kXWcTxWom/WqapmvVp/jIzhItD0aloEpUubk5PCVUczbwgw3dbPIGfL
yPzikw4zjB54WmgLGk8+nY/B6YYFiFWwhfiphgqOU4MzrZOe9nxHkDMTQXn0O70w
AVtuk47UfPDpSWqyjOBoVGkkYouHd5DEDjg1+yKbeqMD8ig03zn1iQt79lh+nsCM
ypLvslYxeUk48h1VnVxKHNWrzt1ZYsjs9C22tMeRhdE4eZt/LbCplSwfx8LCXfNq
7N85uUfS1xUJEjsRJvzsoIiMINHlmWduvkFsaHkyr8oJIDeBEKz4NzWSyEYuTjSo
PE/tdFBL8UjFtYSKVkV1k7U8uYgl3TZyYENeEyXEC5B/B0qvdPTYeLKNGwnkkzTE
WTDEL02JL1DGdYA6gecaLLbn9bpPsBCIc8J3Gg2oaWOMD8AMmd/ZLf55Y0fEYrDm
ZSV1Ah5TY09v2L/bx4Fo+Y+ztMoLCqSlKCw/kBEuj1A0vUU4Mv3kWzhCFJyF45yZ
6qckfG3mmHO4UhYnSSPJL2yQDq0PCI4zVLKiAbUfvsxXiVPOe5EkCIf0lg7N5Gze
eQG8MCAw41qqA/gZdG+drS2R1GF6H8mgLA899NQ3brK+TY4DdjwdvWcz1OtFdXP8
Y5RCt2i8TgJ/4AYkSVFK8c0uOYx5SvdzVy+xBuXQ3BK0SvwasxLHsxz9W2+t6zkl
sO58Lc2fiJUuOMUH/g5Cy6Czsp3ejIUWUDFY7L9xMV9ACArs6dGdmodd77d0bm3m
hEweKkgfv9YG+wvIR5vJv2Mw2vfUsQ2aYPjqvjiUGpsfsX7brLgpxVFHnsivuaek
rDOuHT15iboE6XQz+iST4w8sf4Pxx1xP4pp8nLZkKa47h0pxpluXRYQ/cSKYnDR8
ySzwkXgqmEgIB7OU2EYEyeE9rvW+UBMy9LX8IdK0IdJQMQvrjgZZVvFTcMKLMcfl
tvQGBB8NE79iHD3Otbur7sN86cLPBx4uKgv5h+DGdVAI8RmLuglt/ybwdKdTk4ah
9CN9ooheGlIpjeR2xpvf6GQJ5egCeMS+WrXOEgFffeAilEIkez7bakpGUjEX0rvm
B+RaHn2d134d2T2J+uSVpnPNU/w1p/+YKQhdswcZ+9Ma8CTjvwWr7C1kIFA3TfE8
Wj/6FxaI2otXc6UdFMChLEZTfyYx+lwp5s1uzBRxxAE1t4y8F6Jo1QmY0VtwQs7S
JloprAjfIs8ddcaOAiiOwx+lzKgN6wx8MvQCRxhr3mVrwUIqyePTmBcFJ6Cpv2Bu
RQBjSTY41h8NyRC4y2YxJEAWDkpZxyzLatOqvl6lNKLjUDn6wpBpVEj7wGvuzGCL
rWAfg/zbOIYJTZroKKO8ipX4Ubvb6I52kziQIUq7r+1VF2eED184zbzGXAURg07W
lPdUBZoBa6vlOlLT47OB9deYjvxjLsTuU9883GAIkGsfaDbsrd2ZWvGPEpModw1b
URgFAdbq5lL6/jtpRVDfcnwCPSBrwl3zc47HlnaZ4vcKZ7si1PnoExa1AhjsZoTG
Cxv2PPyj5TSbm/+RZQDoxoN7rTRNE75N2rACMLqXKJ79P38NDlCLRP4hHdIP5qwT
QNiGA+/yf7yKbbe+brYRRY8e4H9Y2WGDwZlZpC+PothWtwYcGY5veRbAC2VEGptS
6tYbcvxSKNC/TE098sLR5XglNVqYcg+DNeCPT3NOqWAupe8uIlbfmipV8cwC82qN
oPpjk2xYVSaUAXwpKp1Lg0RPlQsRqArrbStNG+A/40SAQG957DwKf/AH7BouIkwn
euZztZh838060mJe9/62XQvswvGedAQ57Ss0BvNci0m5e5yKWVjd0IVdmo9IMJ/Q
AyDUD7/TvaYKgjNqzvvw41Nr/rEpacICExEeyrimZ164sLLsbONt/RRrcZufPlGj
JDtX5qJwm/8EZj++/bQrKdGI7HM8V+A1PHGlHmhs/+k02oWbqn8BAhPph9nCZbiX
DwyFLXv6ZezAc8X6r8ybbwWZEETYSU/bfKzPBDa3vMV9xX9MwMVIrFaAF/crvGwt
uCq5K6L0sWve4Mvs9oJYEJOxqulHhLYjQiaVVvfVpk0Kaj2ARVvY2TycZcNjhFSQ
9/jxtVtftY/7PbF5P3xonmJJfFU2SPv0q1VDBsg2cZ1CbXlPaisRDO03xqoKJY/z
qvhwaX64ndkZMFescSZAsnF1b+gMiEe9cTjcIeMSfw20tylUyvg0wLAE8xVc/WT1
j1T3CaK6faaQk5RuSTZ9/JFDfjlUsvzJWxGuFyJLLQOwLgmRmIsPcuMudK3ygVCt
sffHOi7EI6/4SfNdgx/gYg08rv5wAnv1BfbwFYtIFvAuPavy1s3dCe9X2DNaLdit
gqHfOgnntz01uXra/Mr8g/hB2xM6fyXwuh9gVngIe7jJVKBO6A0SagtklyY1JKK8
rz2TIU+opgobg+6Mia5ufp1RG9NsLxrXO9/7ovxYTzxUuDpqBBv/VbLnBRls1LFA
6WXuHLTUA8yJvxHV4LBJaeN4e6Ps1nzEWUB4fINR7BoqFZLTfWQVVTVfQMnXkUPb
Lns4EuaXZlzj2zbyUSmm4D7DMe08fGFsYMMzSx+9vBhN2r9ye+iixwxPcfB3s3kE
0ziVZVJr6phyUBBKsH4/c3FOn4Ca2JJJf959LRw/wnNSEwOlR4Sig3oLfNW6BjLP
Enl/40DsW25kLAS2urz4OzWmf9OAyULeqSvW89uosqWzqhc6aCyncI7y+8ufO1qA
NB7X8z3HBB3lR9J5BLqWJFeUQwboKOkv72cKVc02lfEinnEYzTSGSRlUrMzYz/6g
YBB5daT1cxTiDq9KvzFuE+LpTOpJtjb/5gOIczM/Fx2rb3dmqS0R2vCHJUhciPLj
J1jM9ufhw3E/lDF4jaGdDYEmu+tJgl01hGBDa/Nb0v9jPeEtYFrKVBUOOFfdIonu
4ZlRTwMLgr1MlO3ohHNe9fxbeliYYMm8jyvcGAwE5gQ2j7QTGSXk3saxnJZ7uAbs
h3dNTCrDQG7ZCg4CpAUTdexi/91daR4Ute/pewWe5lG9b7M2PGOJG9JvoIPw5s38
iguMvTZlXhertUmR+PM0PHy28CncGmlubAWXd9jFkxCPUhgy4DJAGdAR7mzU0gGz
tZdJ8b3Wuid98y2lcMNlCBhWWeYWlj9lx9yy7E+K+F23TbQ8Getw3NlQCEexNu9p
yzz1pqPtGbCjEFIE4IUG94la6RtQ9uBG7t2WUpHTpWMWEsPNjejSpSPaT3VWfjIV
XeK6A8K3m0iMlzmnMKKWOcMDke0H7UgKbc8CXrt66Er2bSeH5yHz/0qf+hefEQUS
HhlSdC7SFo2laJADhDkVAV3NjR3TDF04tStFsrmkR6nc/Gc3M8zNWFT3QazYnrMl
NtSCoy+W966baKcbrqljc6FF1H9K9DnZWNG5qvDqgiga4YD6gOsrw929nKOrE6Al
c7IDyDCnLl9c8HJffwyI1Mw9onQ+cVZ0T3QK4Vj3Ss8l+ck4Jo+utiJ7WKJJ+US6
3aCr6PQL1zPMnf7ETM/m9ao1k22R2Z+LUYPEkgjvTeQkmB/V22j+ZzYH/6iREdP5
DHHWrixrzgYrdh9ti1MpqR19tC4ILGfDXrwZo4QFrKDCQRTRzaSrKCcFqVWrJxAs
hn+5kjREJT6tqtj0FgnyL/7fV0SxsZ8jtf6oF1/wzUNOXWID4UEIpUbIEyytxHNa
3FwCcxba7q2NXerFd+UVGkFgLqoJL26xj089jcN7RAknXfeNOwydwa7v5zT40HFX
nqGdHGAPYDQadvtbTo0P20/t9TiP+Wcfa06ezdmsA17PdO/DiAIqDQ3ttz3cgcp+
jzwMqBlOitlOxa4QLgxyzgB4h9fXu98Rqv191cZhKdB+AvPyORM5wY7fzqkropbv
9jLUs/1YX9eV1n1lJuHLqq+lmn6zaz/la34SiiDOsqxW/38nKoxGESS5s8NPTjWj
I55oj+4N3+1qEnLxglKC+aalOp+deLOoBda6TvPs1kkXwFxulVvwH7EplJzvRTPM
v4PLcBD06uw+X0mhS1NmB/fAFs4EP26riFsgxmMdak8mSrYVxSMZKDBn7ziMxNdX
3l6eOQeSiRa2FwPH7PnM6GZz3ztFPBWWfxCZh9GKNiNi4J1yFN1rT2UAnXThCrc7
Rfn7k2oxU7eywhCxlJA57Vlrd599jAY7NuV67DGLGyq5oto95FkEMLyh9wDOhVux
FAN30cDhaIp//mZbk1sujOp3DvgQIY5lDYLvMsnPqR/klXLMGOIVQFsXknHDS3ym
pA4tw7Vptvskr9ntsfCzborHxKftofvLgGJXTxNiaqvEzI4iurQW0p3xfGIAevud
2WH1slCV6TvU/+aymnJTWIVbkUbaoXc8+C1BvbkywU/rbpVtdFXuuXI+Ykp2QiTL
aOB6nrMn17dl+gnsQ01yJfQqQastIdJZvny4WzJaU9vDDBwFGT8ARdnwyZpfEsMR
19PnzCjOG/k1nUbQtWTvcwsAz1YrUdTpgPMinoVbDDRzI7h+b/+YZsVwMkA0r5A0
OWwsPru7zEIbYYwNLnTKSJrMuOU5IaDXV8gPhWNXvnnjRkcIDD+DdXOnd5WMNmeI
ndarHQMyKbIvCwt9x9VAxC+Jz6kasqH8cGyRWOg58m2uB8FCRNJGR/oCcFA7TYF1
X5kreS/xaCH4zC2wztGuRDyLAaBszacPDz0OPeKCVjTH1nW7YpXbcXM2ow2g6xVc
xA7hryDTEhYmbOADqwEZJBaJgODeot7s9EXJf+5h/lXqy95h8WsZBdtvpMhGws2U
2gd86zKmpNb+5eCihKxvuBmajZ95kgHwKlaqqZJA8Yc3LmWGzXHcqCy/smUFqqU5
MTuaA7HubUB/0AYNC/0kL7bAvXgT/AqHR2tS98AoMmFBFLE4bFGU9ytK06kFjTzQ
gcTn6IpIj0WwgC4P3kxM9+n/6zGudGyxpqBXDir/GYn9v3vZwh9UdGKXjLycDwEG
aQ9/GNqBGA1pOKmyIZkbPXLIcYMUZYQirtNU1++QpgpQCbWnhu3GwB70BMyByyXV
fxGH99hPv+lxG9t97oJlhxRU15HahJiMXLTRox87HPrW5eLQRWljrD1IVk3ft6d4
PmgoNL3VunNas4Iq3/quMBRRsLAlPkzcY+S6eoTYMxJZDQERHxV5hxoBgCpHRBhS
XGpKpIVee49jF246ZcorYxOsosL1TRmnbZFZ6UZt704xEYnY8A3UBqqg7J4tRYbX
6KykzgXKkPLgxY1nvrZuh03wjpCcJliyupOCf+nCX3mbjSNd7g728DpqvDFuAELi
JPBaVOyYPcf317VLmB1vg/yKtJoRIZjxJ7OaznnDvD0B7pwcfVv6Vm6avH3Nh7z2
zCaARqZzudwQ732RXRJjWi/GF2ND8F3Wb8FVctx1vsODV2fGD7CsEJKm0ZmEEQLq
5p+2Gi8VzBckAhymY2q1uDQkHmgcFX/M0qmjeovlRMkyOmuKSNnuFAd11Fe62GeX
7ZUm2AzvazuYkZk+iPonVzcLcSq8YBKBac9gNqyP8gmjCSIwYUNdTSTAPl/8AUiu
NSqMSUg2/JYGWbHoOifmH/CwI/gBp1EKTjp1zAmsKrLSHGgy6NNdJLKzW67AAES5
ApvCEmKDv4d/wLlIKl7pJ77L8fRTmkiM7ygSjRIvzeqcHYnqGtaPxNVm5IKWTDXv
khvJGUBfjtTz6mR6rGxGTy+CH1aWmlW4z92JxLT9aotce/93afWfqo5AuY88Dn6b
95ijKaVGJ0wA8dOVng5ZWpAs/4oD5eXqhJbeMntQ9EsSEwc3NPyWZbicXnFQjflQ
fV8dFThH4kw/ZAQ/A5Hb0zP0uhbhW30WR8XAlYgr6eN4B6m4b5e+OlQBwnkFT6Yj
zxGwt0rVKr/AgttyFaEsD4JY1NDCGdsuqFr9aTLseTeTdP1F2vsHNlDYEX4DwfG9
hqc+v3d665TB+Iz/Ah35CKbRk8ME8stiivAbPWOgVBtTcpLeZf0YzmN1piN0wS4V
7blR/J41q+VAeFRFLy+wFmmEVwRm2aCnL3LyCJd437IuTcMCgiZfH0gSBUvISIWE
9GZ2yWcXoArGBIvaVEm2w+ILMNopFBGDCmSdgI9Pvf+IHFvqpJEhZ3urr4SX/5JB
ulaP6HUq/oRTNI0oWV4oF6/3ueTPEnXU8YFQlv/hVC2THrcZaEjXVgxBicEKdxBO
8y9dhR5djFlY+QEIrzs361iy07UzDD+btAkSaIo1+ruhSl0xU+uqkyiq/dENX1Uw
v5IjYizxP3Bg6lhr969SoOq4Al1PpQGyz2WC7Y+TT3FW7mTzecJuAI+eNG+8cjDC
iXHk0Ykpl+rWSkVkYQ73plZa0itehW7z0KB5R/9UU07Q4pvdkndNZdwpROnqyscM
kSXSw6W3gAIxq4DlL+zm0qsmIz/Vs+nM3baH5kwtSNhPEUVLGfNiIcKgeErOxERG
eMq1stIVIiLU04B3JBH2dVI0rtG8eN95y4cNkmhEYkt77imC1lTvDGWcjAK7zpxN
1+UW0vJC1p2VLjf8VDfo1EmAIXuZvbQ93tZaaJmseegrNVWpsL6yG4obMtGqpzSA
2rHpqPJ0EIwcpbm5OiR/3PP5XefuIyAA7eCBFdxtEgZWAIgumaA7J9pINoUnPlMH
KdAZQ+JfHViNGrgqVXAZX6E1DZEvmHAO/pA3gf8SQcQiZ8GfEy380MC5vYmwgmkz
LbrYPSGZG3jsJ4ste25kptF1nP8zu9NDOFMiPKrJBtJW/mpMJc+YAObfMIGjXhrl
/8oEPmHorqMtJ0OMMP0MTdi2EAquenTyFK6781h/iPmWmrWH+A32l1+RvKZfy+K7
CsU9pjCTgHiynzUYIOVQBvhYgTiBeqayPTCBJBT6RhAB1sscg37upOF8NGRdwuz1
ZL366OBm6V7hzJiAng1WP1Z7XJ8g2BD51u14qYAVpTl3MkNaU2bZGjgkiMRclYTy
72FYumQkxRpxWBm86EGCB0UaZ5rT8h0uNumcTw8nM9pAudQW46aZCJBBUuIy5gib
T1jn0A83oG48/ghZreEAGPuq77BpweGw+0RHbPwn7IJJt0oC0oNaxC5DyXABrcS/
BEsTcOur8CXASOXvpYmOpKJEML89+qqOEb8ntOeRKWN3/UYGTI+0P/shfpSva4Eb
kcPxWV1Mnk83O4BbyJllYOgIiXdn19SMwmducti3AFWBrNl1ICTn+c2ypevI4Sn5
eRST1IX+WD59BFAvEEzF1EUvG+8BRsSingAM2q6B2L4i6n46Cqs3t20yFUMC5No+
04q3JxJrzIAWBXKjq5z7p2fXJErtB93nsaSRGiiZ6NDIpqhnSzQ/RogpmE6CTVFa
Bl7/HvBjPF76iUWO5lz2DVcTv4csOwPbMree+4FUnaOIB0v1FX95eRMLmq0txjl2
JLp4+5GMFHd2Gq++qvNgAmU1f0q5bwlT+yMj8p0lfQ/t4wLvrTh2EdRvhcohYGul
VSbbUdgv3zdxt9+u3+hSNF5tM3u5RojRVgKnLEkuy54XMrcjc9SL66jx8V/rl8Py
iepdJa9NzfEqVP/R33339XzJg8xHU/C1ckZc/hhHgim8BpLLweYkY1lcixMCGhit
oj9odNYrE/ucoHgVQd6zoygEDjlsiAOwdWmFh09kYx1t4d8Vyn1bC4vb1YRpkAwQ
p/4tfkMbHSn22SgO9+WnspIYO5yAfI27o7d/xF9leFj1OYFtzTn/eiIBxksJdq6z
Ox9HAhhugap40je1/brVd1qxddMk47/QPl55mWv+7ycnW9VSPvwIY8x16lfTOzBl
sUbg9mhx09XgYWcjGpxsHsPlQS8o6OrZW3IIqgi8KtnpKqacObVukEVYp5hQdcQU
0qzUwgyY9odNq7nCeJH4Bb4qw6JfNTNbCZgyN6FuBLO2iTxeXH4+WbOV2sDbJRDN
0XFx6omE0KMjSJS41BuN03f4yBX1f6ZulLJxZrO7aVLTlx6fscLp/lE5VFR4b/v/
Dm73yUZNru16GNWo1LPhf3ku/GzdH6dM0E4CgTcvKZ1bSm4FyuGu8kIkSZTzY3Qx
+hGcecDEbbDL+jkLkWVbjaVgOkeDmwM3oj+hFCf7SKrTx1nOWjT6Vkf3faZ2dr4R
Kwz7yyuA9xGLHKzBAJ2iofvqGaiZ1B3f5r1oDLFFjuGcEJkGfbjp9wcE+3Il1rPr
IyYjXYu40iSLwxTKQkGUIocvEWGskyQxnw5fLCfMMFpak07p1LUumBAPrYL4JQH/
3AwSaNAsSCrqA5KFUanSK3S8e8w6c+uUU8jcvjljX6SZVS831TMafjAsM1gxe88B
zR+QRRxnXHKuPsYQdvdKcp4wAmrWl/GBLJCgtlV63CtdHMpH+p0X9BMvFW92sJFy
PSSZQz/p5Tq4Gx2d67IGDQdPFzIdwFW5fJ2CgLIEZZO2zv7VsfbgjFUJO5PXzHjd
MPBQ67n9S9CMgRB6feQfKXFaMzaM6wXdFct0cpTaSkYk7YRR8JuyCv/hXF2IHa/m
0W5blNY/i6fk/Zx7vdo3oTo86NGSoNMFQ5nSJHOKaKflQzvmRSmpkhW8U1aWdmPk
FZ2pGieeFshkX8EfKO4uEdkXoxHwPjfC0ho/HzYUobGAht7m9c7TBRQI6rP5BxXG
3WYbfx1F+1BTuBJrAo5iHSgNlH8viwFLJUVDDWpuFgmCYjfA+v6ekFGBUyeq7re+
gvmyVAV4yQ5o8O94oSbUKPlm0o9Es+rJvs7yGrkrqbwdNGupvTeQUlu30EeYnYzf
qA8ORQkmNWiEwzWdCRLQ0YIZeWm1C6e7dafTOKj7D/K9ajo0hQwE7B4y4JzY6pcO
vN+YOa4a+s39bwbVdjlRGGC/TNemen3GzFVmKU8c7zn2Kt5k9G26l5qg33B6+w3/
H9s0dDV2eqqpSDrpniMj0px77sXgKczmw5qUCqJtf29kBhgky/sbagbCK/KD5R7v
0YUN1VdXqD3NsFdjyPJMfDjEGB9fR9pOAFB9sIxVP8MebRicXCmlBHWK3TvURTP/
lM4OvUZ3Ho/Ixm2+s1A/v9HAZU21Kbezwcqh2NCZpN0TJCx2BagoXKUI43wRzyeX
hXoybKjDJ4bTpMBKV4HVyag2eKPuJKDbR1BSkyXGCe3tlG/qn1PTsmV1z+BOK8Od
x8CXT750iOJ2tsL74m6xaHrB+8pHtuwN4fTIcwxxCJpXQ0yRCRJNAUYbmYT7A/I/
1aynCb0VyW/cuDyWcbjKGxueMmbYjBT1HBWfGVwKalwuMX0Y8imO6SZNgbL3qQfg
YZfImBVNyM8gqx/p9IbnEJmpE4DVCiVIt2nMYsP8oaoUUP/X+g4ZIFfx36Y9Ln9e
biURaycMxOxx4e5TH90tkIoongCxfEzBypD3vCIbfTT0QaBqZ4fnt1UXG9KFSVn5
OuuPo2hMXj8mYDinXXIB3UNnRuQx+zw7oCGSifdpqdcaMri8JzV+RYtZj+bi40qQ
K+BY0gOH+bHMpNEURczkSQHvPo3SodYp6YcA4UlDPuNf0gRwyMLIvvJUJ4fYcVsD
hHY7cGgWLKpUFghfDJMiFUIw0HaxEyLzIm1oUjlvvcx1VkoP9cLUSwJlU3n7+Tx6
2dRKm0QhQMo2lri96Peyd2G0+Y23ZhymXwtDrl9A+i5E5nZ+O32GPmLAk2k3N1qW
Zmp+/GJWrBTDgb3iRnPEj2u3sCt12FmjhryTG0Cx9NZNvekeftii/3QY2fSm7spN
iUjNeDO+CJIvzZZg+m2y1cJB0SnqRAWiAACnH5Ap6a6ctgoSNjWUs9F2/V+j/Nxc
8L7Jv/ECrCQUK4G4JUKRvMnC4f1nw3/TILjYKVt84eUIbWbMNmV/sIMjrDS8VgpN
Vkh+QkSulHR2h2b8gDm5RDMZ783WINHCaidKLKaRrIGOKQi5Vln2t3ikep3X1d5V
TrcyBPnlztnA+z8mSUR7LT3sCM/ROJDjZ70189JXRwOuprvb9fAx0BB5lGdFB95q
A5qx8aFjM2rKwBTl1Leq++QyPyhW2wefjn2NbXJsQYzeNnI5UT4mi3k/wtsUT0Mh
I/JrkCNMOHhp30yLsQ634nTri6BNbqwnN9JFT1ZNpi0AZUso0+HkozMmtm03fOgp
ryfTKEqN6Qsws9ARAH1XPhAOL1NTV+bYUHEC3fGRdEHOanV33M+D0xnXcZxpz8/R
UbNlrT7WiaJ4r4/4auJyxdOOvZp6ABFn4I6+47uDs/0grtAp2wLkoCR/W6gBWu7v
rKTWF0P8dHQZEObdhpnq71YF0wYmtbGJ3WNBtZlCRF25z0PM+G71CxxLTNEmkXA1
jyNjiERXaMdaxtNwSKR1OHvxCCQELCwQwvp7ZA2OoWBCGwxnGPyQmJlyiyNoKHGX
mufXfYpCowkFB8N28+j5aRxiN7fSz1RJiuPU8WjgUwz/NEY4HDHWyj5ULAtK9HOR
oKnc5Glvj6LbZBxMivLAEBhGPRyLkz5oU3KfEbbURyYh7LiT9GwnsocUJvj18jVQ
cV38RUDVF8vgS+EP7pY5SF10/MK8dzpsNrBb8GzdyIY9pjsGa0DjYh5Rh9cvLWol
led0pnGs02VeEXu5rrxWv36e/Eq0t7JmzrbzMESxaNWVdieV9HVl0593LJy/ErKn
RCrIC7OuWTdxRGsx8wV06GJ2Mp2rNO9FBMxgIM8BLy0I37teDHnQ1717QmtKz460
HLug7GPjy3hJ6Na48V936D0E11h23AgR2DcQA0nHojzrrFsgPHWfmcC1MoMQaGRv
6zDcYMoJsMyI+XpLezKioQ9IfwO14Y1t//pMG+WJUgK7E6YkqTGIjGk4MNlgOVX2
B5+OClUfFoNnKAD20tAo8FvgRZq1oBruWUwiiAeohDAH7gWfw4/oqkVEx0sAirB5
tt6j1ngXBz/a9Eq+LPNGwQ//WYxGynjEmfzmjg62HIi7uBfEKRAYKzIFrtLp6E4Z
uDHrNF+MjxvX/Ou3o5ZvMytExlYJjQEqHeejZl1bVeFfeeoc5Q+qvMsgTlnxRZ8H
yRUi7JjnZEko2M1KyZmh/vpCbbxIVpdrnnxKPwCgUdqS2EWBSrD8cr/Zf7zAp1CU
SXt+WlHElf/ghnnH+SG2beEbeVKlKrtbSE6LUlg2b8r4uaXVLJon/NsmvHfFq1t9
BEgJNBZKPYC9Q4T4L9uk83U6N9YvERGs86icx79GGsX+gaksJ0RROcCAp70DQb/v
ixHS7B1AWAn3gy5lZIL5oUvPuVG6Bld37ZGj83oKR5hZh7nEzmfMOKB9WRtVaRmW
hvftEsA+jakS0OiXZrBmCYMybENp2iajG2AOs2hyL/v4y/z/cxWNiej9I8zdAYkz
vgL8YVtjL/A09iWEnTuAzQwKOSzfA5OIL1IlUjKyYUGQKH8jyixUeNrFsvjIRYCx
5azK5ai9tZ29nFj2mVQl1/HCAhCIwxybEVt+axofF2aA69ewyLDlL/sT138K2dk0
HsbezMdJSUPxAA1mCXjYioBwBcaIaxrNjjpkVA0B1Nn2hD1AR93CeAVQ5c8D1r7y
7hDMnNL3vmCzGOMqBRCcYLrZasZuHTsOi+/gwz2cMLBBoGQLcx9/v5LrJDoGTJC5
xa4kz4afA+g7/4Ia5F2UhFzE9zeT99ECZfAaT2C2b3LCgfXjbaDISxVbffwtF8rQ
IdPFenZz6ytjFXs4bhggt8ar6Z6cwp0F98lAECi0JPl/PNOwk1VSn+j7Y5dBT5DK
yGWcOCfOLUQ13yheQ6T+V1kcDrGci+Um01XMjBXmh6v6IWZxNSONZjPQa5LDv+w0
Y9RQgxE65/+FTgHgRTXIvEdl2VS6U78dP5cNrCwD/QEfrNbFB0620ipu0kA413gB
s8CsB6izettk86VNYYpiayZZ0fPF1QXSh7TtYRto/W38FqLFGs8wCr//5pcX0JR0
ulpqaCy5IDZolkpQljI7zMKhsUb4jkVBan0If3owqRXzy1loJ9xMaqDA07OShHfC
LPSauXhflK1Z+lp39cUt08mklp2bkjmxOhkl6DdqRGDMilz01Ik88NjgYg29Ycdr
5kYeUksAgTT2g77LUUvW5z39P0LPErJDNGGYPvTtWPWbLGFUSSyE5689Fck2G9wt
cROqNpnnaadaZkw0d2bITkOp4PMXnwZkCsEpkZzGXTEH5joxPqb5CRvwWFMzKvEG
9BPr6voLCEEcTOnOtTbW/nIWXO3mSrckW+Xmo/P8ctXXqKQkACCKdA/fVheqC8Ln
YNKlhq++97KJgzbfNdol/FZuUrPdpzArqoq5NF1PFkZ9IzvowMt815SSM5uxjZ2t
Kf5eaGqwzEp7uEuBIKOkycbhUqSUiNTT1lhFAItnxdA7QamccCG1Ntyn8LArRx9X
yBNarbySZ+UtgMoUVVV8gLkLB+axPFxm7UgaoAfn3ckjllAs2fh2OYsbApbYJ8y7
kaNnIXAb3vuj8XYabSptrhaTkX4ycYU/aEse03uLILSFRZbaw76xbA1AN5kLq7UV
UWplr4VjnBvq9LZZ21YAjC2pMzeqreki1g1QZSQRnXS2bv+6jvqV688otBMrsiKt
uBAK71pJR3ioXgETuT9JePIfOSJbvX7HEXurHuTQWXuKG6H3HhBc1W8SdLBydym5
yFLtpgBckdeI6ztb4Wh4hSxZ3gUnZFODOk9mP1P5l6/ClPhggNo3an+DBlw+pbhc
9s82wP5645dAusEbaSB12u5caS8dGiPdyljMbhBgK2nKtR7cASPZtthkEjNd66ER
xQqleLaT0qZ0VVq2ciXZZZ7rGedaebJyokJEi1pohSt1qIu4jakY6imQqETfWleH
cPb9x/em7t0UFru4mZyy8KJgk0YIx4FaHnwodzzFbiOP3INd5J1+e1gtdSCCMyf1
QtdAZbWAcMYKgSabj3fhUfDt4NQiK9KTZCoyj0k4SYB5vier7ImtsL6gu0njk/yi
n1cufwfpTXACBKeJHDiQBBzCnBJcimqKeoWiTHXEoCypNDyMoJxHJpuvuAmSReSa
aiUgSpRvL6GkufMv7ad9Ip8+idUlxtThP9jhAX4RQtAPqCvlpI896qCk78TZ2CmP
kYx3h8ZbRKcQKIMpQT1YKryZ5/K86zddWXBlJgWhposSrYJKlZOxqpnTPvni5K/m
gmMavMQeKD4lVnHvWAg6oo/VLsQjfbwExGy5+GsNxwfXyKrRwT160UO/dQ2EsZJo
pubxzvgu9anx9DNURuWsfYAovEZwKnnqa+4h/S+mdd1P7sr1/AINUmBdpbHwCmxd
1zLHPAxABwVnc+rA1gNIpvlJsIJRq/JwKv9xhDgx6HYMg0rp39OBjG81bwdlPN27
9jO1GdoJBA9MQMMTHrUd/nU3ShPXiNE+x8NDMsEMOisqBzM+2gg4DO1BHtY31tM2
Y7ctyhcLAsXPVGKGHOsj8INkMIzJtZ6STj9xVs/HpsoMErZmXgGzYItF5LrjRmLJ
qJQsKn7i5cSxh7hKBtLSDYGm4NNa5gPNIxAtI4XkjjHc7Sy/bxzCGTtSRuiKmWBc
QQJyVnJ9Ukt9L+eiBTFleGxHz0nhfaR1Kz6+iK/VX9oOtPXBVrnYVxQYXQ+/vtrT
lIW9Nk5q8pVdGoy3wWDcdUNzZfHQEiqJMC5x0LdtI+jKwEZ0X16FlIirEjERNDwW
nDMkiiIjCWupJiGNIvLLum2durePl1c+I+CbbupB1orJpLBAUAV6rBt3qoG9jJNa
tRCSvOCUSu8qR1RKX+301xmvgwTizD8cjyp4bqCB0GbZ4b+a+ewhLFHfdwjhIOGt
llctDz6x17G0IoACcWsE8YCy1KuaSj+7Abwyd4vibH5gPDoB7Xn2F1Mxw1c0iQMR
guVpK9/jSc2EVE3aSqB0N+OYUe3RtouEuWJ8SlkfTFgNd+1WDYQeF222Xi8RHnXz
m8Yod8FqMuaxH05lynYsQn+rOJJkFJT/NiJ3WNRUqg8MYKWVryRuCp6lgYFJl10h
QQxiLz64O269uCXgBq0G3n3360Bp6rZPwLVgxTCbcqOY9t72KqhHv6xSc4/Uw7Z5
mV1LfqatpCEmXqrXN4dd0sx/KBmdZJVO57dUxrcxNuzicajXR/mmopZ0TY2V1t+e
LIT85gXg7fvo8L01TL/CZOcwO4V8+qEABkDGkl/YyW+/GLLzhqfw5FE/mH/RIs48
xugB0xWtiTMX/80oIF284Ks2ZcdHeu6UvOSAn6BvuxlJsXRC0IycfF9t0MjIvwhB
eIjB6audQgG3oRCtlTsrKIPsUGiVV2C5yiKjkuV0yYSPeSpPxDrDROE0meqYGeIa
9BO5uiVcTa9vQLJJFx20OTgVWo99XRlV+Mzm81D7+OF5sp2ZtpYn/MmJKBq2ZQha
GmEc1AK5ejQh9ZTBwYXZS3qowW3ZAf4zAk8CgMXSUw/el6NV5anO0RBT0qKBgO2W
PsWcR81Vq0FLaOu6HriANaulluj5e5+iamMyQ4ayTyEUHr/docbaNs1IO5uojMHO
yPYT7sy/+JcC/FgYSVykKQVE32lFdrf3Fi9QrfE3jYyOXxI/nbnlBqGvB20zOrI7
UR2AHQGbINApxbwKoEdSFnNo2zW5OMzMjj2ZGRH983gjm+q9DM3zU7j5cS1EmzMZ
iKAhmaPudtZjyMElsb3e8dZYLySQ4gK8Gz9bMUlrm9H4qv4mD1j6eaJHPr3A9HzP
MKdt8M8iUISIp8LoucxK1u9cKMlm/BlaEwvnaYeqEaqR/lsTnLLOHfN6VmIZRUg+
p11gwhsy/XIW227mpsDr8ZFGXzNCYA1u+mAv6vEh1QjxtOvBbKzICkTGcmhnuJ3y
5vOvG/vaXSTqVbDnqmTIb5GeG53eeEdL9UEJwxeef+TPngz/wYQCuJlLPY5760JS
0Q3fnwHDJI/8ZknzVzlNgdaLxSzvOGZqaCwU6Ie4nxMJ16NJCYIIK8RUHGLWY1nX
s+V7D+4fpcRc8XqvaxHHFgp3HiRfu812L5M0I/JGjoJ2fUEnq3Qrc7gApkf20R72
vOvZrll//YNxO6PEzwgaDyvbKQHGj9k1s2DhTSWdbmS/2pMZnST3W938lgbDOJts
DPVvAB4hn74hjtGO0BUzENoWhr6dyk2vHeF/66exY4ynwYSyfnmQY+ag3I2DVCy1
O2pcEZN+y5v4+OjcARO98YmfGJxhMpqntQXtRcsVDlb0NLrDeTHnBFPnp/IGOPdk
e74C07tHU9GI0XEzMcaaX/ezKm2l2h+mFxkbXDypGHT/kheAc5jj47Tcxr8CAkm5
ZzVoiqPcKditdyRfcyfYre0rpDqghxbDBUZ6eRdwHZvbsw6A8Bh992iV1QyHw2AW
CsN2Dm623JDrnL+PP0WvmmqpnLbdbndxp5oFHI2p1IuNQUn/Gm4p+DvctTiNulN7
rsOu9E16tWX25uqBFfcBGFW4DQ2KGgwPjCUPOnie60OudIEE93mOHEuWqK/WbiCm
Qli3eJtsEeb8Ljzstkn5j+LreW/0ieiK7+n0gdWSaeWltH12PhU6CQ0+9GUXwUvB
oFoSQDqVJv4I2OD6El2sGnnJGH7salzXcoqsmMiE+NndlF4kQvm+E5vPS1Mfapj7
EsEklgEGJOJSb6it+wJfkmWXXIW9ppciqynzklEE4/HgN5BBOwYwz2xRo2go7gER
NozOmJpdnrKE+0h7pvdl2vkLu9jQlOg0WsHMub3BDXtxvhqFGpTiN0ZpoBBkJnsg
kk3Smhx/8cFTwoaqmZarxhmHBbXBa7B8xctmnmNGhY4RbynzdNfL15DQ3XCxOmXv
tLq4jwqk8XFALZBndijBxNlW34rZxEr77Mk2O1XteGmPPYGWSGyHtCNfuirkeHAh
XS7ssM6yxRHjkwEOmpOABXSz49rmayDpa6At0JRlTJTKqjfJrOKc9Em6kTe3k2ui
cRItvh8FDXthpa/v4BwEQxGaFCjcoqw3nqFlWGTNtRJm0p/7Lj3xQsCJeX0m/CRo
MIq6lEOvjnd7lZFoRKQpaH6tPOQMN4EnMwj1AvfCKsqMmUCtogkgRVobbnv0OCfp
bIi9WYm8IcE9Qpsi9voj43sHZpBph3p2d178ZtXtnhLggoezxZshWAkUOHeINorS
NMhJzb3e24s/G5p8meE9Agga3ymMzxL1iTnjPmi4FIaykDHt8PhGDyj9PVph8/N6
kJ2SSLE+8SPJfgZBQuKunynD4l96RVsADDKa8JAVn5qGHr4wacHb+rtxwaMXm93s
bLjFw3DNgn0RXYrUaohiDaeO7l7Osu3fFd5/CXQHW+djrpn/+TQ+PPxIPvm5rE4M
kmv8AFXsD0z2y/LOlLbpnffXH0mbrUb7oDkNrkLNPcX+e57YoIa3059iX88Y/0KG
qOUi4GXdE+SV+DTqX8GsnH62SubRFH4JL3raAGpSGto9oQQcreAUp02AwH6kwSY+
wDWf+NbF7ACfftHVcxGoCZvE6yWlH1CVKOrePX8UX9Ga++5jRRjyCr0M+BPrZoRD
Q4PcGw01vlE1oNqzMK0m5Y659NEzKOQgpUhq0mLYV8xtl8x7hyWQDBdhQ59FCDSM
7eKSHxx0LYof0RJl9Xf6cQzV4Ax7Cj/mJV9G9AX0w/YAl3B3uTMRe0lh6f8J0ak5
wDWv+5Z60w8Uhr+kVNnR57VcDKX2tnjV1sqoyqR3DNXle3wucSYzgKJDfaC/TCh4
e2iftqA0oO5L2qiwzTX066zVdivG1LSVFBAu/16I7PnCarrupt+wYAJar7YWBZZc
AM1ZSiUu0yUSm3xRd9QNR794qibGeoXjMfeR68d3G5MNwnf2fuB/S1J3biHO8U8o
fMdqdpjA5JwtZH0+marj9FljIDjzQJ0tsbGx9egfs0yCHBQkYxbGxxKG9CNEo7s3
OVeb7/5Mt3TEC/wOxkWsLI0p6Y0lZ2OWgncJs2vo0NvrNs7s55gD6CVVEoUIpDDu
zv85jBUQRxPo/XsAVIhgJYZIJgeu8yam51LJ8gTvEWz/1Z4KRI4JLEOCn/QIksj0
vmG6+d9iLyu2bktIQ3M5DonHbmuMMigxIqqWEecW/QJZ0AETNEeIp6SAkMRFM/kZ
pP9K6SQGqOtI4LbGwph0EA5SODvf0yMh1nPOMeJqRtn6MLuNYD+DmYIsR0+0P4Ni
16U7ohiafzKFz/0lwBgagyaLrXoxS3dPrDPpl5gXBlk0E4mEyydGYAW4IvR9ebXl
d2y4DRxFG6y8WOF6tOssrOKBO3N2xqBo7bWCJiKh05IoaU45Urk73wK1Ea5ckXyg
eO22wUHaJCMAZL2Z2AlKqDmkzS03mNtxh5751UIuuoxTVBr2XhLlnAcaixHOnv9A
mIXJwjxyp3JTdOaHrZymx1rAycxu4M3zYgzeshJ24HQJSDhI8XLYN5FjI2w//pie
RoU/GwGUUahRAo9cdoMnP2Y4yaTjkL/msw/MikrHOEMLrHwEfZhFZUlZq8ACsfnH
eynsjbbnneM0jXfK7cRN/0KNd2sQi71DrF94p+gU3HkQ6ExkTezEyKmVIcNfAod/
THy0+VtinB4mD9nZA9EzrjlFm5jyohrJIPv2TGwElXEAHd09rGnKnl8ODaVlfenJ
iXHwED4EuxJCfCSesUi3XDNs9+DVl+dV353nRueZTMVLze/pmYg9+yLkmh2JKc+2
yQsJKXpszMF7pQiqNukyIpiRq57qCeMAtgoFJnuuY3cDNvyt1/I3KI8FSS5QKEpA
6hEbb2ICniTfkqb+2p3GWf98xWNlTw55boLM7ec188uwmwNyVn2j5AWTOyo34Ipa
4aikEwsgJDFWoqVdfYMXDUZiZbYY0Z/swmW4QVW5nYGt10SpWIsL1vSM5lnU01Vc
ORIQaNqXj2blrbiPh3bePeSbHN3VK/0GQL+A26q3QM3cXUax/mn9U77/sUg8Uq/v
+vD9GQqrmXZpX7t6r0IuUwK4kqXWzCD0gbAcicYqxQhgpRNgGQpQA7GzLwh+jJPl
VWZZIyybrKT0a2zdZldfSOBTzIUvF56TRiq9o0Xib5NWgGgQ/JUECpn2fKjW9qt9
1xbqYX+5bE8dEg64PJBeIKxLc+jF5j6YOf6+gOhoPyAmmT8Vf6ZyzafXynC/NrVx
Ux4YptadVBjjV7UYwdHZ86vvu6M3mchfXY/AIQ+N3ADqG7KVnVZwsaaO9uiABd6w
SQ9EJei9f9KHJIbYNWrb//h5HtPsia0BpFB7x6GKqcIoPod13tcZuxiO5u3UJW67
H2OUX8MmT4meymohqS7VdsxfaYxGzvEsK3mKC0bDLZtr+CyWG6kw1RuMgXB+kZ6h
m5hsNrU9LwI3tgncZHgp9ePFi0RYsfSu1pJ9Cty4N6/GHSoc+6VubVfPEYbRH86V
I3nPpWEap135vYj44Cv7bkKk0bmKkXXI3jMEM+EEAvDWGxgTrkxoVLaRVkb45cZv
49V6FDWnYo4sZgVIpyHZ55MIsb5c4q7kVOzgPb2rQkKJseXhGS4JEy2TMsWIp8QR
17kT4rDauSeDgIzV6o+tI95VoQCR3NSQOuR3lJT1+oZLszN68GkU4yRVDF20TQfr
EhtG2V4q+Xpr9T60jWuMX3JUOhfTm4BwErxGrrQ4eS0TkG06/ev7a92SIoelv/e/
m4I9BoFx0FnXAt1TwKsSptkKFi49Cx5qW7I7q8tHrJEOuw872aspYDSoTb3ayq/O
ahQw76iZRjxbBw3pBDOOXaaGCSgts1kyfh5wsCGaX86c0CyXqlGcqBdQupVi4Xof
38IiI2KcGt6aJt9iS7jt62lldQTC9+Ybs+h55A+tlw9zRBHbNxIFL0W4BCBg7xgt
S+cqPgs/ICKJf9rTv/qmW7sWf+Wg88HX7aM+UStKovZ2eH20ZsrILH9H9qlY7n5z
MR/HFTTcV+yd9mY13CR39ADiMbppexsyoSQ6gY+Vyt/nemz7LOynccg9ISYv5cr3
E9mKw3DfQV7DxMXWgnsEoLxesifUp6pxdA1sdHwuw8iBQigJSVH3px+02wZUc0Nr
BY6DnY0SaUKk/bx0FTgWASxs6Ev7y+hj/N9FTfkTrPsH2WDPFkRIHUwPXML3kXR4
z2pZfj7eaMY0S+sfTyHXaspSyeX18RirIVCGflG+YsGUSjnWMuurcTgwgMbOlels
4OhKko+6XTJ2hDWfeMDtyaHkqIJSH21otZPW0Qn/SJkn9Z2fI2W43fKPwbX0K7vO
zKbYWmWntC+magUtaTbcyRT7Kj+IA6gl2hyh2wtOBJsJFZmQtmlKd2REsq+HwtwP
XhwuGP61fBoLXa20yIYWT1u/ca9gN9d6YfFnZc/tUeuaG7hrh2k+P+h1A3PlWgV8
zWDzXssQzrlD0Cros5x9D8rHQSJ2txuk9LDQ+GL3WPWlQyQyw/BiYy/arjKcfYhR
Pfld+ktedVOFkiKIbttXKV7xRItmcePSIIO6zzEZLvto3SCz13Cshs0R1g+K+I4Z
v5y//tX4KK7atLqZ1u6pqLLmP1aK3KGVELm+J1QXsueewHbMQu6JOi8hlbnpKtcA
vmhCwqBhO3ll8anoBFmZOZ1xZQC+EN8BacAIhGav7ndHtf0GyFhNJe/upWJgClfW
uksrfG8QxWrLrfdumNeXEjhjoa7806zfR3DSThJn5PUkf8cDem4QdazcNay/RzhU
hcVtr+TpSu/OSwgg2mkOOTh/mwkvMQcdMLdx1BQ8Oj9ussgtIGq+JJd0Z6ZgPTgD
kExn092Y8T6NVXRxNgded/oS6QPBy1qISQ23bKAFchQgfXo1w4IUAcb239UMFBn/
rLqxPOON7hiQ0kXb4K1H7CBuJRnCX2m3LwwXPi2cFxcj04huvadfiZNM4vPEPnMp
lQuh5JsQ27b6Y/efmm2CvyUdCbPwpHrsJeZmk0wk6M5PDhh0GQ4fgyokWG3HxNhT
LDiyej93nGwCO3CQOygou8IN+BXIHyNE1TkqpsWRf61y85Ha4VxKd6uYTOlZdw7y
1kbcPjSUlhETDa0+ntUocXwuyyYr7l7dAX9ddyVAba/AQJ5QwprnsDIwJpb8j/dz
BPc9xx2Ziu40bQ3GfrqKKApSJzQ4wrGkwMSmW1XnEuKS/sdwiTUD9wB/2diK+Mbk
nYkmxZu7Q97KoqOTGG2K3Kt6HNxsaGKMrZbR26lNPm048wm55fhBEcZdSxKmuttk
APmHhfk7YHRI4FvzsLAG770YNxLKNRaPvsIEAkFdUAOCTvJUkADys1nvxfQk//6E
LG4YzuEFXFDWdZZVwZS9uRf4AyJBLQYpA2r0i82Fwi+nlmXBPvNepbL6s9tefjYc
y8iVSPFSAc4FN/ZZhc0nsgXr8qPvi3WGe5Z61TW5lhHXiblvdT3UZwd9LJQ0ljl4
aDLYt491xN2Dag4kYNlM6dw5u8NaAtAON9GJXwoGwQiNDtkCEdUonxhVWRuCf0aY
05JYxmC6cymWqzLl/OGD9rgiYGlmT9neG3/eAsOtg1czfLcSmu94QmOyHUv/Opv6
eHV5HPX17I871vfwMs5VOrw/ho8YntJN+El1i3mBs5OmGP6ffsYLjAB10kXy3R/q
8cmA2dYTlLlrxrMdtG2HFsca2yFbSU03rmlrgRItLnLgkwXbrONlHGfMS9LI8jCU
ucxjrepydsLE+IwJenKHF29Uo9cewnZ/C+uKHCbOJ4LPBuwvsG9yHEeOyynjAWtq
CxG8CZ2bCZJP7EhyHJ1X1DUelsHGYhdBNIlQ6W+JwZX9sQHMENTgcTTAhVmXkNpU
C4ODaVl+NBWxOBIZqy9ra/zFBHaQKmF1gWyecFxhhksdpW2WPSFfVYEQFMVVff4G
Bv5gTerWRjjZt9fy81nPr2QCBEMeBlGa6mV7qzmTnvZX45RO5zVJQrx8+Dnw8uov
fU+A2LYfNaFiqRcPOF4q2FZXg/+HH029yIi64uukgUbTE+aKo5pti8yAOftmUC5f
fiT69fUqZ5eO5Jh5t1VGt2bdaPvikQRGdyg3/b3BH1Dqk/5avnwaMKlPflKX96U/
Y1esagAUIOfQYLXGuA+a3AaOlfWSL7ks3Pj8+JBlTE0+gNoe8l3z5xPpf6gGUHdS
uv7OURO6Skqj5uj0yoYhfA0/RYZH6GIdJiDTVyG9k3WOt1q0d9ajxxbTZ2IzAnTc
hta6faqzQLRF5YI/jcyf6kpkG34+vQM8J25R89fNUWiVkL0EBDu1KJAcnCplbNuO
B5CRhwgeFFRLPthDiGUr+93M4cZOTiu1JTNT9Cyhkjq/m8QZK8dqTTbw/08YKSo7
HEl62NAhlsDRxeSrig8Zhu3JmpxV7TUJm6IHyQc5lLYHGI50prsYEPbZxAMWCYoT
4QzXqLhf2yPVCH82UQHSP3AV0BoIq04+FZOsmlI4bg9vq0svo+fmg4m5qqmn6GSG
Zs9FMtm6O8WbdSsgFZKatomhZxTrToxOlTNr17ygfKxDF4PLG4+hzgNTSzEJuY3I
9wyCLKrzwdPqd/ZzB3HHp1zJL1JEpc+Zbg+P6uiZm+xqQk2XOJUY1Xk7vScKTe7d
Vou5JJhvB4bR4ATOlT0RNn3FgwpadLkL/GfuxxLBsRFK5/iuPMEnVyqvUygvaWdm
YdTpgfmRay+c8RPeL/LEul9M8MLIYzIClOcvsAKakNaO3A5Fuun4XItahf20rCZ6
beRapoUy/KgE0B2afOup0McBUxnYchZqrIAU+egpyu9GyXiOWEAjnIffs/ukOUcL
P7RZy483RzCb777zvlmcxqKvxbd5obrC7d2N6f6JpVVp79c5ycAaD7EfzTQmDOrJ
rVxNi8MtLL8y3lvz9ZJi5UH0+dV31hAqBJHIcs5w8HEJETIg75dECNw7/ndtU7ZX
MS09h0z7MorIv+dMuQnUacSLsElSWGTSbvS5CgO5BFMMIKTi4cw0UBzMZcrPTXSB
Q8RYkgU2ZXGFjOiGnh9LJ+pxR0C2N9KD+46q01MfqKkp+iqpnggwtJmUINmoDvZ2
hXFDmMMgO2Ve5PcGNyFhMVS/xMfMcnas7plunMtTc/wZRHiJT9PHt8+6l5nNbiCQ
KEKDe9OshavLza6O29nsBOmpQ0rgLYgPcsK0NE/MJCzfC04kMwSchkL+YXZy1ZEu
18nnARIIyT3wugPEvk6QRhqd0JE1ZD6ORsiBjSDRIQHhoa4cF5J3YqPWJ43zZaJB
J4PUJzOE/TA57nCeiuchXW/3eWXMVoN2DpOgTAvxyhLn6DIoolqD+k557FBLW21i
KvLt9SeZ58irTenvmoP5n9zM76i8gLstT+6WWAEmwtzHO1C7wgyA3q3fiVxTYWuf
SLEPwrorVrazpS83IquCF/IgAU7/2CNeeF6n6CcLOHtFnoCAxCyrvk0ppF6LeBpa
iB7sXeO+mQU31/gEcULSAAiHgfpdoPofQC/SARDz6L0MA+UiMYTP7Cgz3KbQIvHt
WIAANasZWlWUyuGnxIK+MyamvdLi+EmnsYHkMl6Kcm4ZgpCwjX54Iaod4UeQrB54
fsmySJU0AgOVhCrtTNCDHegeDfVpqErEh36ImIpA7GJ8c7/oNmtusQmC18/Q4v0u
NIucthAtIblPoO3mHG+3wNYkNcpKsr+xR6N7h8pTZBfDqH+jsyreeYu6AEZPk7zh
U/VJDQz7K69/auPynrasp125tSzxTE4C9e3RBLJjEEmenifbhnM8G9bnVIlLHlm7
9VwwdePGCW9MbhJp1ykZiC1PKRilLRieKSowTsvJFkmsVpIoXi6UwOmZNMVV9S94
RsU4Pn8k9q7Ksem6uRTCEJKJLlDq8OleZmi1GotXMQJhPwxkZKuqZ24REcm1/8Q0
+9ocSdiTOAFcV1f661VXQD1RqvnKpVSq5g96iImXMiQFWoFd1GLvrcKK5xT/fcJI
nOWTUbBqXh45/YqHTVFR3jJ/HOG/tNvYO1Btd0uvyOP28cVBZRhGu9fC+XlrEmup
77f4C2bldNT3r9W7t6fQ21nNBe3aUGAb1vw77TKRRQZ0D5fVMWnYxcvV1f3ATHu3
MNpJEKjfg4Xu5k8RlrgE1C58JOviG8Bbltl1DN5z0JErF/QY8g2CAy+Fa3cHRwX8
SyncENTTXNWBJqcW76cMOHUS+RmXWP4wPQLtFlmP44n+qAnu1BdMF23cDN0Oxi8V
EbFvrGpO4IoohPEuOvkbm1X0g3HJohStUjAG00GwxeqS0mSEmh5tq3hUtfueQ/Ja
MGTDnUpkVSaSR3NZ91EinZwAB6g2T2bQxMfS2fpf5CL9Vn38UgJXdDc5k7TITyrc
mhlszWM4v3hSvo3VfCIFwppJaIpI1d/Txh4IHGMDrT67a16xMto/oujSP6ft95vC
7cGBNC2xrtMXbdQ9xE83+s9yNJIY/T6W5t4ic/FUKBNbeMSqRt2AaDaXSpbrcJeg
hk7qZgBanWmYbQJU32BmneAKNag1pFpE/7dBoOhqOHJee7q2LooQDAude/ubDGfY
h0e2d/BPZ3zIS++MSNKmc+dt8avaTlg+Rl3qn3NWtQ/bpUWUZNHhzt3g2+O62lIe
NigCbcOi1mb8KtrueAH1NsLtPFQ0HMwXDoG9nT7LUetI0A4TM2cFL26uRr9PuIvU
ePHVpeVRyUP+NSyKN9BIsGJPLYcHlbcC77DsjVd9D1BK4Wx615d1FRO0uoRmXtE4
mCsbR90Uu4zVIuCBJ8uc+Rzj6bJ5mIBa6n47tV+rJ7iwiJK8VAXjKNIxXllJt+xp
hjifKfhZK66usq8Ux08J4hPKCnA9ilq8q3FvAIlh/UPko9VF+d914Q7Dv/OlW0B2
2oitqn2WdwOt6evDlNsTV3YoCmdnofNSb5qMQc2rCG8r+pZ0OF9/9uKklFPx6yBD
dPnaRi2XABPjEkkCAOY67FUTNYa6IUfunDxSfmuQo+2JgIZHwqvcmPdMILNHWsG5
rzFlmQxVrPXghoYmyiudve9T6iAOxbQkC1M4bG8OBgxjdJfa1J4EM/JxUNqRAzv8
dI+MFjk6A8SJNq0D4RYQPnfq5ixM1Noa/ZP1n3qVFN3P83ue1LOIAgsFVrKV6f6n
vZ1pe1+KKMco065JCETCbl5DaQP+W4XeFCIHLfHRDwSvREM283pIDK1GJ2NWW4UJ
Vc2tkPGBTtlqc5O2tMTf1qxL6muN3UrE3/0IYppJubP7nFW3YwnQy5BFOlCOaxfp
K25wito0T/WAO55I2hqmT6c7CFnjBMFAXWAKxTAg9iZY3jgm6uJYObEjakSN6XCG
SSSSQtaE/rsq18meyZgAD7mVfzBpRgnS845GVFYtQk2vJAo+SAQ5dklrrrDM2s3T
JH1FNNTjot33nMHVrxlY9ox7JuOdK5nR1fvTEJRLQaPLtTvk2OgVJAR0If/LuDdx
7qXHN1dV9YYggskDS3ZUN6OgcKZ7qI02rsxV+tNGF902DrMCyaI5+WebIGaRtvq1
GIaxjSi7rCpimaUrbaleDw4ij8ED26jgPXMG7oeZsjVWDauuBd75vsw0Pch3Mokn
ffMkohNu1zOpo7M+/vs3EzYZYJeRBDaC1rRTlRmugL8FYeixUkQOwscffgrAT++E
cjvEvbX5GBqtufwRxIOtqULIEWBJDTSzGSlXS8DTzbdV2orDOUnjliUS6auX1ZJX
mK/1S+/6BFb78jM4faSuC3bZNtOxQFatTY2mmBFgLQROrRdbD6NoBD1KshgTporO
TpHSATYLW18qZRdGCaG1zTxnVvV8NX+ggeImerHzv0CyQxizDOQ/dlyds+hknZgL
4/0Oz2UkvFk1SR+ehvmzVVh4nCq6MyJH0TD5VKJT29zmQD3cbwaQFRRqFc9bprc1
ZyvTmRnK3kGZtWXiRCHTloFalTyzASkyts5uBVZn85x6XAuL82p/tbvl1s2Zy6wb
yySDhnOWf0KuNj92cBFUNrkQFtvD8ELIgF1st/DBaOFaiYG6Or52STXCrDbVqKLb
x6aoPheGUNFZojsmALrhX0sdGdljAw4ZtV9gEU/izjh5TCGdi7VYs9pzMX84cqcI
awo794puhZ4VuGewcBRtvQmI3WLAZKMUO+/hZE+jIeNjLduN9QQJKju2ZD6oVSTl
IbLdafDs/mgoj2XObG1QJptTDZhvk2KMasErvSVC+0FUtHY/8gb+drK+CUjWNvkR
E6fB7rVt+sp5iKsZmZChlnqoHQnjsll2CEu/2VHVR24R9+wzjDyQp89VsY4DEiOk
xBwzCiYNgcVb0U93MPNFv7b76tKMk6pTmJFsjBLQdG/kze7/X+8/STF12CYLHt4C
cCw6tlkVNqAH5GitULDqkwLHaklHc0KXHnCiw1kkvQb10z6o0Apjc3QoMGaa3mgl
MEVqwAAyb9Qhlk9tT8GaiNLg6DyjcTerk6/kncQERvvrdpNdFdJZx5yvP0zEEkeh
fPkoeHYnZ+bL1krket3fpwS8dyMmWZco2ouEMCgqv9RhF2SCnjMJ4nFIVD1QIlo7
sO3TICCRZcgyajfXGtrmqlnI6KF25Y+MSAb2ez4dXVi3IHUGaraHZKIwxneSmUaH
jQSDwDj7/dIQ9cqAg+EVhwlIBsIXhwBUR3TgFkIy7VjvjvbaM8UPqz6J/xsFLvnD
GO4bF7gAVjdK9C9LFbk4tUMY/NtmNdkZ3v9nGuoETftFVC1HxI/78u0rnizxGUpO
bKqSXsGCoE3xrubHRlQRzttN69P3B/Pcu6axPdCGycY6KCPiYdLsUql9UQIEt7UO
GJgwTaikPrG6uHSOaaDahxhr4LvTPh1PRzfGHzKOKzf/OqL5E3XWyfu4yS6hlVjm
UHWSnssofi+QsP3b6+R+SQ+YuKIn4DPq3V6+MP23AuKtQQEQAjnBMIPD6wL2HnI6
Z3SUFTyGLfxByV93sm1kOonOWR8xqJt418tLyVLamdVa8QKLsLOLsowDOIRZlKUe
YPmr6P2dV//aZ3YojDB1UDU4GNBUYCnLA5JXU/TWhJ/uIMqDfS87L75VPNzJs4/B
LDWW4CuALxzZsUtXlMVE6LuBP7TxDWFkTdsocfqoh3CdSqpumov8xyzn9es/agqc
6ly/77cyGESeIKt3iOBKfDeoahduT893/dxSd7zN2Odjd7AeJqYPhAZD9dINtFcO
Iq9da7kN5VWox2lSpFRSTt3IvqEZV4DHTCbwVzwt0GXvePUABbWsoMBc+tBRx39l
AWFzy45GKA3mcfEbPeOU3sKCsDmEqpqKbm+N9xHBKWJB4HW5JPW9zqCGYvRT+8Dg
85rV+diAHnUO+wvfiS4HuyPgKFwtfC8EfOrurDGAvm1qlTYhufUxx0FqN/z4K6Hu
zyVUUb/y/v+RFXf2SWDoT6yd48wvykuvMN7uX469H8mJOU4z8jVtaliLawFO+LrJ
RiYuFDdVnRS2A2VPDVjKX+eXxO1xBwOGORpiqpsqJLmQse182KtFxkdrXQQXoTzT
P2jeH4L5frVJKOSeeBpT/I/I8AkFnU3VDS5NxUMT9lEyI+axuEA+K+TbclJHFbYM
GZSuTTGuPWFTU9tFKyPKkQDsHo2UB5QQ5+CIzMgvXP16Q3yqIFpz8X9ct9CS8JvO
Q9js7nd82Mpf8fI67YVZWRijHFJjH4iX7zzkG93it062EpODdRMuuvmuryPKJPy4
0zOX5K1e2BWNYP9Vgj3D6wzNZNxgo81Xj/UAvNVjY8EhunuAXPgbgqo8tIkfrUE1
Ln3yzyEnUrftn/C42e/yNs/67l1r6Bn6skGDjFI9ocDg4GUCoev2e0NyVkCMSboE
yVlQiQ3DEhdVW9txcT06jo3Hc31uQJn4DJQtbQ+QUxT1vt4ldiSV2dcXN8Q8ly9W
poyjWBmoRI8Ylz4sVlhCXynQGowSu+89uWIKN2iY3yoMy3TctmNkP4yOr5dMEhQ4
UbBFSDO6+U08qDEFi+k/+c8JPCdEbHmAzu/usO3p5c5UdTp1/ZQvb87+Ih6Md3xe
qqkBiscJRDqPm2EwqLHST05bXOWCg9nJIZxTOCJhdIivI0f5OqboJU2wTwVhw46l
0C+QPz/j0AZ7WI/dygIeCp7cHwzRzA+JqgQ8UG6mwoBt6vfWYtDu/HPkWbhC0Vuz
ZM6vF/CUdqWSSXPcLu9oJUoGF6jaLqi6DOozR6V3U854mBG8xGbOrtbQyMnzBDEn
w6BfUrCFIsFmCznf/AkkOGv39h6EVnzfsamZsNXOQ9zvamuBUeGSJVGwleDYiEuJ
zlaqp9155cSzQqf74LuOfMGQm2/rYpVVLyZkrK7BdG7PfAU+3KKwWxE2BNId149x
D8BjDxS199Em7ezMxzexbOf2ZHkb7CDNL/NkZkyCLItDf/csY4zT0RtFTM32pm2F
nTYE/+tLruwTiUi/kRoxbVi4QEFtwJvao6sbWz6EZTo7uVaLNpse4Nx0+lAmT+Vj
oKXXamk2QmkOzs2u/om0UyLZ9CDUrEY+NLoWWVRyjVg8ccJZ3JUHBBONakbZF0j2
XMPmoF67cDMRO4OmecfeqTvaECG46kRd+B3xmBfYe/l7zK+D12ZHM1yfehe28FVi
PtiHcUH5MT1ItGqgYlolETnBbvGX+6NqCHypHEQXsM6xMtX8f0DBp/WSwBG2rROA
SUKQzZef4iFbre09nzPUYIbcjNtziXA0xLP+IeEP5Cd67LKQZJTjehTs45KeWiUu
j05Zo+ZO/3UJvFrZB/5d+UBaGoekwF1tWnDdopMkBoO/n08qZn2rJfR1gGhiAEQr
CerMq9I59PuOf+/m/O5koZhTQh9rW6K8gd4Bd7Lsbz5A/Aw3wEEH4v29E4ie8jbG
+UHk987A9Z7hmfmhvF2HE1wI2ryKTHy0tK/K4BFHRuci+/LyK4biKrzVnA7H+Ru+
KJH0JwpASz7OcoQbAEsqEhHNY5mvfXHHbgxB246d74B32KFzof/kUsSVYSQWOh5X
qDyiBeWwmkSm4txCz+udDJrrCWXTMr7f219nJ7HNtZA6U6O4v+nDLFhzalYyICvc
lIe649+11uXueArWrvUwAWwgpXcRXyUhRLKfaMbCBxadmd/DOCaZ9i24iaImZ+0o
+6UFzWpKXX47p+U/p+pLaP2CHoEdUzHDmbTlQ7AtXClMGEUVJYIs05COTApo1haC
XAzQhsBnPdb3olIzM6W+c0HLU4YZm3YGhFqZjNcDHzKOSyBhxcMfqfpF9bQex4hJ
eVWQ1GeXqzLSDCmZvp3d43lStP7MVAywvT+ePXJfOoZ/YRxooS4ILZ3biivbM4hu
+2Hdp+KcNW3rWsVRHrVs4kxTmd6UNICAbQF5WAcjcSN2d7MSaGDx5yjw9qPGZuJO
ejad6uX+L286MiIBO7XgptX2G65UpvL1XCMhdYYg/BvxLjfoRS/zsBqXq+gwGWfJ
cbqTBkvw16yNOKHkFh7HtpvVPMR9KGgz+D2r+OSkTbTZJyKB6mKgK4oqVbMcNZIt
1HV8gZ8z2B8moiMYq0eoDPi++8sIAaTzTi8SATpiVOpBs5crBw+YBU9C3g4fTxWw
A8o/k2kYDHoPXYLDzMJBUs6Dp36D9J7GcfUHaJj4c1ER1kDuTDUhleC5EfNxDr7t
ZjZMOo78TNwO1T3y94cRdE/uC8DUPp34rOyf4kfzMY9BkMyrhNeKHrJGhCpVIFxb
ogQ1XJlMRfaHINVvwPww/wzyBwYJj/j0qpkdwibXQbAUZSAN38NrLdYR7W7J0d2a
E8JnIs9gwC+EKAw4vvpjVdr5Fk8Q7NGRRMo1VCd4ObnM3odOR16UgrpZXrzuAa4J
LZi8Dvww6eHSakqPoLgh5eeYCJINlPIo63mZl0kDhTNHJQ/JYhkorA/IhAH3gqsJ
RCnGdlnQmKYmkBnJIGZGieTMb4TXuj21hz6C9Fm5rTnwvzYVGjepEUADake7kml9
SQEuJfRcYD/sRYmua027H0AWp6ukbsjavnwBPY2BJ2rezt/KH/I8Zk/4WOOqawkG
rn8fckAepvlEYxNFDtYGONIzWYF2jQoH7cuYXHpNmhnU9YIRbDTEESpuodgtro5n
xsus3X6DOe8GWT3k0fPxScmnwWaZH38thZF7+bPkIoqJYDP8jhutDFjElCriBOke
eSVTGrGJ8AWr2miHMRyrHsaIIQWvMs+yO1vh96IjDnMzOQ3b2nuUvo/74vMtpZjO
XcDUZfZ5JW2+Yibnf6sGcM32/BrewHDnOqRJA64eHofUttwT0HJZmDSCz8K5U0ie
yVV5MBE45lxsJOG2A1UVRGhxBfcvL56pW1gT9Dzj+B4xVuvFyWbMEHsdFstAVZ6R
SzGgfeX9bghxr7Hk4iR97eZX7jNQV6Uz24Wtd+DCziyf6Glvpgz1B87cJGielane
vyAMRWNmwKWgKwqKl61iFUtf+nR9+LYJiQRcpobf59K0qgQUAib9F6EDmfqr1Ul4
cb2KDUDkYM6uE3y5JLaooyaCmEZ+4vng88Ih4+4biDad2z6SCeof1E12/FRusPCM
Bt8AGwYhVCHc3bT2B3VzXlTc60g7IDsokS1MA5WSf+XKd38mWJvm7r3zf/aH0z0r
ORcFb64ifVRW69TLMZqqIhTnJybC4lpSh5g4CS2YHcPFGI2nRiS5xPNSR7eulr4E
EGxIQcLOc9jX1UCUAaCwEjVE+MjjGsyKj+RNAOi8XISLNIuTrSmmqjeKSKj5vPtq
+n3jbb8VXcX1rcvU6om98p36nIA34flpZPEQ8zf9iiOb+6CfIpKxmlm4y5aDQDOx
OFiPRCiynoUO2jPudvO0slopOzvdjq4mKFyXKpp5AHjnDfFzxx1Ua/o8maz2KJwW
+0a6wwc8NW7HxH2Y275r5KjFCBHdU6As4gmXg68PJc9V5NqF6DYwm89K4ku4jYfv
oYlAmZrz29aN3pjKX+eWFiEHGy0PMIzeaSFldDpdW1dSIWjnF1/rHlk9JrjvFpX/
cjggoaRwccWZV9Y2zE3QZ+MYVOHSZvGA9dmfjZCmw083kpxpH8/J4g1uGfoIF2eL
+HqXwWJDm6SH+tYKqqDl+Fi4zW+uatyorCv5Verm+ZpAqfUyJjHSqGOCAa6IoYGT
95GnjHZu7bz5g+JUmy+/8aLUQMbGtaUvMcS1m/NK7YmmhGlmyfFaGdA50B6zHgBv
9tgVqc9oeKfPLfLpRsCN0LycD/ObHo52InAsARKQu4YXIaIFPIDnzZ1rtYzGE6Tm
vjSgo+rTRoNpRsf4ERKfxtt8g0KWNsZS3T2X4Te0/gXJE6ijw0IAZmOEb+Fd+2Hk
YmNyjy4ruZ3oLFX34QdPvww2liNcHxWIK8eCyUTfRuAygCUTytQpWCXiNA9/Lr2x
lXwQf2kemeTF4nVwlPpQTqwlKypOCkMUdqG/yrRu0grBUa9KTdjvpqjXbYMOsShy
OHAWcSWfUV8KhZX3QDBCxo/7lCjC1nnD9UEgy5SNTUpg5MAY/EaDMApNQJIEpeBR
2zZ802NNn1HXodbD7ldYIfwsg9n5/RZ/w07V0kXfJ/uH9fLjF2tvlEFBcfn2QIkP
WLqrvkIEXYgS07afinJUnZT/sUOKXWPC8BOjEJZHcWwDvUP6hGNtgrhTSkYud1Zf
0Ea63xEOqXLEVnauHF8gzjuehyf4hzJYiJ2KMk7nQsXB4PBVP2bsxBHzb05FM8OP
NQuqYkVTeSotHk9xz/YeEDsdRPHKZJQ/N3QdmUugbpadDThmaPC6CVVvyMp42k9M
VEsID6FVCbsNqstZAY8KRFvSVlS1+6yQmi4HKrHLBsb2H3ypTPtU/07Ay7jlFqb6
TPBaM0pT6TwUpZl0e/y1rDl+C5VqZ2YjfiHeznph3MNkTw7iLEGoDhA73vzEpSQG
zqReUr8b6rLYoejQXSz9ocp0tYHVQJN4eaKn2M42rRUm+bEH+y/IfDA9aDG0ShI+
ODnb5KpSmzN8K2oqi1HkEvbcnZMfB2GvWCu1kgbOFemROIUFGB2FeUGOrtNGH/JN
AMjSx2MrRQ2LoI4qY8Gxnxue80L/LuCoQRHlzJRFYtMmqw7xGMs/U5ie8iBajmc0
r+Z8leGKpd6Z5WvB+qYHufuTs4CCq9Il5YvgbxW7wvefeRLargXTblUwGCZbFkuE
bpg0MNG0PkgbmbyTH3Yup5ndqgxGd53pxKw0K+k3uv4eQ3e9RUqcjXyQCDLuNLo9
kY5B2PcCCz+KoEyyY6Ucau6+3SWk/eHnKBNTz3dgvs4zF53044P5jb+iB3ilfo3q
UuOk6n/wyqTQUyFYzdtN+j4Vnrr4gfDTONPv5I4PQ2soP7+Q8aC4EERREdOmGj1z
CajZdWSdeQtGNqWy5BGrlupt1nGaf/YLD7sAf6SFRI5H894bWnZZvcwJIk4MGzFB
ebtdF1MQwynN+rX4IJtT37CJNyVnpx0+K6uKVlOTMlro+URQC3DCTH+jQcJH+PiA
J9T+uPoO50RzzLA50/oWofU9t2fnLQFPFHO69fpfYOsRfAmX0nr+FbYPf7tAvw5L
hC3Qw0aM52UhTcnadKiDK48oroaA1+M4H3iOKAmfNwa5FqSM9chMqIKvrxhTQKFC
NtDhwRzYRXXNgVwtR92x6sN2swWLn7NWhkA3bU2HHPSaB93sLZHwOochMVEAcTGv
svHO1RnqyAluX331nmJmyy2y+E5wEJGFP8CcvBI5MM0Vcre83PRGnM0BzA+1aUDk
XZw/1O+EOHkrO4o7EzUEpfkW82zd+MpGrQMPb+rN5AHHGpI3g9i3WiU3qS84dvhj
oSoE4HrE4sFau/6MTdviYhMAqKz86/wNstV43bVgAQMxyPfT/Les9GCCvzuHItFv
jjgp57OdMtK2xHUiW0jRJikDTJjOeynVg4RSj2oEgxcBOxudLqVPT3GjFyE3bNiz
O4WTfpmikMXCloLNxo02Tr9vIJKBizIDlndJ+m4xIMl4ULA4/KoWavKV+eZDHeIi
buNKCVcnvVgCDG4U7Y5QtucFBT61xDGL8AGfmWWzs+1C9Imy1Q3wtC5uxxBSby9J
++EVh+FNpwzqnyuhlePb5jGPACWuuLnnfZaXmoX5Vo1r9QxM2B0ezXy9waysOTf3
ihYnB1FgUY84uzolK9nWRcrF/Bjz5j0WFjLJPJaTOvQVxAx8jx/kVQsrjcSCyJE3
sKwc4h8p51KMTMYjRQ5EhZfKZN3Esbw8DL5dGsTqjaJQZKMVAJAC4A7nreeV8BjT
1vkadF+aqK0oIFNT2Z0agLNts+2PIoY4zD/DCDJTvR+mS2XjezSKeo2fNin4FcPx
+38oWWhkxDj3e7OoC+Hh+lk+aVSTwE86C66qxSrfPSeT3jwX3G03ZtlwiI8EhPgO
+P1QGk7Jq+uACkQR0912xuiT7suxJWTXJbxP+iPVcpjdvbd9S3qyjxqT7vXTNVo2
3o5ZeZz54iXSmYmB9hmYB5ByGANPmL1caWhFC8L+HbyFgCvKYgtbsoCehqEJqTqV
fjosojYTf1CNFTO4pA/fIXWv+/iGGSLP/We1FLK1k5FK4SMmcBobShFBCuH/mY15
rkHGTuiK/nV/tq7rhptd/+U+/A5JTOB48tmxTD4wX47tpW3/KBG+GRxgRSdIjghE
IubtlbdB7nr/EIlzX1ImIkbgU3ze6qA0bzvE5OvHHO+E6DrHty/Et4p2DpOsmbO0
KRYAN3E/7Y3l408lzp23uSuwguxiyMEVtxYSqlwQD4EDFFNz52u3ILAz4pWsvklZ
PQU1k+7q5Yjm4ZLqih163et1l6b9R6i5he8KI54ZGooUbJmAijQSL04wcEmZW3HQ
nELUSznXujC0c3NDaR+nakP0axu631hGLE3O/+MEqvHxua2XN06Ltw+c4Y4E5+lq
HXO9RhIVBWgSOElIoyQQNy4JqhCtR08eWDwGI3KvSRyq4KyDbfHEKhzATPUVbHJq
m2ot6PgSDAc50j2ecX6UxV3B2baJiBhan19iS479PQdjGwgQXyT8tQmhr/mumLcS
SzirgPwLSnO+PrDMrgshct/KVisQg2aOEsrwhE9ytOU5GIm3y6UJ5iKs7UDvGBEE
vwCguazQUL9zPbJvbVJqEAQCwjfN2FTc+g7s1uGzKNm6uauatag6pm/Qtv0FSQn4
Aw+2bfu8cquACJNrzisOah4VML/SCb2hv7CEXDT9w21C6w3nCREa4S2D2mUyPpfy
QEnEyUMlWvjQMqAApzx4uewl3Y3FsnGj9lsWPgtpxWrl6CM7yB8cuSdNSuiew6BY
laMKgiMGhKmxKLkTzwWgYtLjlgiDCj099cb0L+XQxPecdi9pEJduxzLEcz8hIdEn
Uo28jpUrKk25PBuoR0zDqW2vRVMkSk5/fR29dunq5pfWNNRd/mzvyBEn53U3dS3V
2Czgylgz0YJnrkfSZO33TD+yswqvThE4a8hDyLxa5Zr1+/mWBiZ7kxp/ZjgltvEF
v1rocCKA1fJ9eH9wL3vNPTXVIWmb+8mtKIxz6wZJzECJG2colgqBDiwJynk9Iskg
3aoHAD1HS7cqsfuZrL1ozwKvEl6WOx0k+FrWs3hkihLDzECWf0ocvdwt+c1sLPYU
FGiQv/YLW0muLBN+/dkQifaI47P9hBikYqSvsAOTRyeQ99UAk4XxriVz8OvsplvY
JsWOrusmC/F/LTYYRf2vKgW1HceRcOGHge/g5MFM3xBqNASVAqqombkNdvQvZJb4
vOp3LMpe9H0QKxHFquPU7vKeyvWlUI0BwvCcpyQwhblFe/23rBDwWqFe65s2raZ4
YiP7XgOxVYGtfXe/8nkNrQM+q3IuF0bsOq8x5LEW3ELN5ucTd/w5DBNmfX8BdaPa
vBiwVaWvwObvhrItPxOmhUJYVFO2jOwfKwPNA8TkqhkCmAoWfaX7GeIlMQpNSCic
6G/6xEIqusIRpo9b2kjrVt0NxdxhvfIytIJoX8BzHmbHAUP5xCBj5cUszRGujQ4U
CwvrZ0XQIBXWTQqLsxOYXbrDojp+e5m0LamPj0bDXQ1Ll2JxopnJ5wLW4ZzhhnRe
nAQ96dytvu+TEOS/rcsYsK/XggxMw1/0Ds5qgQjD5eBKjKpLZKwuFexfIa1oQaC4
YfTGYcSEvj/g9qEH8nnlAT2AMbVNeabxOORCyB2rNMwB5T1bhm3hOcq1KZvAKM8V
26Tn1xvHDtVj67CfqwmSupjgaUybckjlPJOCrJViXwG5ny9hkA2RFvbliEug+Yqt
XDecljuKc7kQ7l86tEpFuW+y+Ipcl8M7+/K4SocR9cz9yYWLxT2MqlEFArrovxrY
46MP9yPdBY9EuWp7VLSYY1Xsv4iTszJlHu8A2413Bq8Yfzkec91JRWRVgmcrnAs3
+OHIjWF4pUPI6is5piRNQGrpyhyNvUWc7jiw1+PAhFPgmb/qBqw45lSAFYNLAM8/
jN1SELJjEzpBd8OYpVcwKNvsYOJQM83r2o7BPwvscImHdYKH+RkLAETC0jshVyAv
hdwEqlMFlPqVh2bokC+PG0PKGEpBfAzX7knRQAVZXpXaD1It1xhL/JWzuokOrqw3
X9B78Wv1BwuLAT/Xz/E81AKTz39fC9MF4FM3fIweBuE38x0mqSIkare9AbhsvqIP
zD2rmUy/cliCz1NVu33O2H+UrqMkyUaNvJU7r/pzu21h+mUkjpdKkartoLYPE+/P
LOd5LlVON1TiReIyU1tffJNtc9AsXUWL7xCCDc8WSDxrg5LYST5z6IhOCEHNPg1n
bpeil7kOOwBFOntC20X3mWgTJF5gB/5Ms6NLZ8teyvu7eWuoiNTR8poHKbcs9dNM
iEfyu9UdLF65WTfIPGiIKHEB46DdK2+1DORjpm+L2AmzBbQtcqAlXyTkYCcT87ml
OPZe3Z5dKPaq1nR8R04hxJOOz8mqHKlAMvRVzCl7B0I1AMKMPdzNddoSyU3CySrC
pAjlrpatylP0X+g3sndvJ5HnfJxeFnyRQOAeDkD4pd65DueEK3IUUHFXS/dArGqU
t5lC7C2KLjsQYKTBq9RT42ImMfLmz5i9UZgFCdWvfP7olPNVVRpoXcF44K8BEKva
UiGUGlcoS9FUXVWyFNbCA5lBeksbs83Kwcxkf5MXZ2Kr98O0lWzNFkcou2+ex8Qd
qJC73bCQEICQNQGjNQgtMujhGYensS+vBTNaAwYKg+rj+kwXimYRqnt1GZ30tB9a
HkeXeoO0H1DdjEHiUwQNxuW2UgUH3rpV6iVhpv2Z2zvnCbGj6k2wCsh28F8uBH7k
7WPCwZercDHJIoR0llNspdvibPY3y4Yjv1NQ8FUJjqTP8vm1gf8fKgzUqeyGu42b
AL0p2YzNlbIkk1WFJi5ClXEl36D6YCkdVj8wKMEkEJPclg+6Tbk/1n7LjJM2chWV
OaETUjG6Y4C/iWbYS2bR3VmdyvAjEvW4BJxfuv9fVT1gH9zG7OHf5CS0eCv1YwR/
FkYQz/7C+2WMJyz3SK8StYSNgBXO+xTKuPi6/KLIBKQRbedhHYEDIygFPpPswtSU
kZAOBhlPqnV8Jx8cJqzOzhvzECg6fyJQAnt1GCEdJ4UaxdqQRvlsMsKfETwjd0py
b+ZVygz2XJpYg6vOsYMswAzrEbyEYaN6Tvc+jz0ulrKMzKTceRKwYHkqFpbJrshb
xFNgT5h8MIPtkWuiILt3QkZLTrJvsy5GJd4w2UEFz3lHg6gIV2IC1ePKPDmx2iYx
k/CQbTxUL6qiH/2c2V1dcOoX/707FGEAQ0EEyHiB8bOvvacq4dP0VK2EfQ1Rn6ib
KW7n9UkVTPE8DojLDoWflk+0XVJ8x0WpqUn8GyUogOlCuvZzYfLANLoil8J4TWtR
pO0LGGxVKPayoe+wkPiZiSsCBFeKERn/uuQr4mF8wbG6MnE3PEcPSwWKoAW1wYW3
qndsMz4zbfRldErVNqS9aUI10dDg/TPJXIJrngUZr4cHrrzCBWK3PuTkt8HLU/pn
pdK5XUVO7+ZV+Q2TGwfe9hMPN58vKnbSdFx85/ar1433C6zttRxV1XlDUOfyiOLx
XI5SWHlxw5BDk5uzC3M+YVWOtdP9OpN56+44lm6A8Um7gLAMLdW84EsPrK11J2bU
ZEK3b7/koX0qSsIVMJKXI3Kmgye3xzIV869nZvDMnDIJr5coc8NDKQrKlhI8CeHa
bbESP0RPhFJLdkx73SmWBTdHVNsUH0mr1Ip9Ra4Cj4fCBJ87hhcRRgD/9QUk5v/L
i+mRva8ZGCI9js6J6mmK5yg09mgesdIoCoUZA/JoU0CFv9kwgwLMoZEOL3MNuGHH
7tHcAUekATOfw+Q75gV9xkOs6KlQ6FvyC4JsauY8kMlRmvEGDfv+2rrhXp/i2+DI
2TeQsn3KgPoAaOGzUXns75V/r8UOIxsrkHwuXxurJLfdMnFhYcYbGfnilQUd0Pp+
BXUbbN7NhBta1y+OCV8AKetGhVkY+x4NXy1XfXXi9ShepLZpNZUT38MPF0qOi9Mu
NzQfRcxra6Lex2FiP6vFzk4UU2V4gNMkpvJl+2gzf2fDYqOsonkJqq9V2Ndq5115
San0HjYBisVGnTx8EZ7IgiLPi/BG8KWgxVN6A7uFC4eVbK7XsPpHs8sEkQY0dyJ+
oY7OyOMOdlVWs4xMxMQqCDmCYoRsY3wAUF2FyqtUjFbK1r77dtvOuB7TZaOYEubV
0szXy1vP6HKqlyWzdtUwQRZNX17thNnbaHf8KB9YMjz68xV3hbC9QHF/a0NVaC6Y
GV+D8Fs1qdTqkLK0tLSHaFh5KCM3hwxeK++/naU7uGx4wT4DilJq+TqwmTV6eUWv
xwYnBexShlZAnJGO07V0a8leM7ZOCBaxqQB6a9y0dcW+WdXUi5kQKwloviifVZyx
618aL3MNgeRZldaLoJ2IS2e20NNYnizCqPGfFtYEyaZA2wwpuDQ8gPxqy/AyUOwB
cWRs7oRP5YSAyHPLv4YA0OHY8mRashsFj/b1fOORxfWuIOFMWVbKctK5G8/mNrwv
l4dXFYB3inoHKqqxEu/88yuytp9ctECytkAOHCghRxwn0HcpHP1pYBxz2AecLIQX
Y4+wJQCUbuzTfKsCz+ssKnwFaog0OYXVn1hlLx5pneGXbk55ODKQESvRzodpp60S
dQK2ngTG0XAYV45Jsl0UEiM1pLLMoxpGrlEAjLtdMjgZ0uNKl7G5XvDF7lhkcKjv
e7gVik2o9p7N3rsXH2UbOhPSB+TawCbfEnbaCpxF9I1ml/pLOgCZNRW/n1oCUhlC
60VCvOlwnI+QSqbFkW4DQOcEn4QxSQyh3OqNMYfknQPTOWXXEnD79PceLj2+gh+2
mzrWdfvE3aGHeRPU91u7KKAEqxTMvfueMLcDWpdLcjQmCWHyNjFCyjqvloNyhwBL
seDHrVnESuTfelp0lboBla9dt49TO69MfoWRB7XCORw1Q9x+xC0hkjTVAt1FJiUc
q/gY+9A8a6vMiuLRLVBvqwupeW2i1vQ2sFc1UM3WC3JaO2rd2uvTrVgp3HR84DcI
k17bB9O7Zo+Wh+ondw2xAVkM7gM56qFPUq4/kCluipbMVt3WHLmIokTUqKnEUF38
HeT/PjnszcHz9SWxQSqeJBVxNEI2zylm0MiGeR4B+Vb0qMesAPatHIrhbKVGYwC/
CQX0KN4AVZdxDJfG7gwK/9eRsfbPYb4vBFEvZ1uMmhSP0pYSU7ED8wy8hjPr39vY
PFBdst1oH2sPvNQOBAt57dGs1UxcY/+Nmz8rYeP6kpPo9yjwUX/D8HQUjYphZKan
fRBDnZUgcZJlAuofbbNm9+K2MhpNyVCn6cWJ3h2Kp5whjxH9fHGhXHpPt6fKOyva
w6WdCMuNvHzQYvA7lR3ILv4dXZ0ozRKEk34nxuvHPnf/gL5X4bshbU2ybQWPu5Kk
81DdNY0J92VgGr6IUAyuzul8CGk+PqJbxjBFXpNMN8d6QK7B6MHnt5nwFyLqw16v
fcehRPsRmloQpucgHzmMoAeRv3WcZC00VyUfkjrvY7xHhj9dwpfKkPIUGNTi/kLM
C9+2wU4fLYNfUdB659wBNEeERRumqGCrRNuFblGUJQAVH5bRQsVP/x2xvMkQt8IT
f1iTFq4bwVDsS2KVrR+e1em2on0jgaTpzfkg1Cy3HjwY1CuCma0d+Cd0zQVbogtx
7S0ufyTgYLOohYxUv0S66XAFZQJt61o9YhlldoLtoHUlluGGpY8EWmT4lVt53Ssx
ztInQj6/aQvUMx0xzSMvhs8MoVttAf5m1SMX/yNJCfRbMe9aYslXojLpkG+zfdJB
t5CuXxiLLWOLr4B/s+lROnl5IcAveuxZyadzHJNCnBn1ISrh0qkm7KHclGQIVi3f
qR6jnWkzTFvRsejiaFnY4GGsh9aerGEoAtuyesR0p1xr4pRQ+ZZ6eLGr9FwzxeP/
BMJP1ziiXubcCwGtDdr6wHmWQWoR8G8hpfeEoE/csOqDwo7gtwjA0sQJaynz0dPk
Sxo2UoIQI8uHX84LRyuZm2E5RfL7zpSXm0EUoOPB0SxptZXRrmWcufDMNUnDpRH3
KIFhilK2hPFP7gVD+QvRtzXIwV/NqK7RWH3CydP/ZzgqojurijJ+E9HnyE5qSILS
gHLjRbajYIWnyRiA8dj2s/ssnEPVGV4zESQMnj6SVbG1GAhoBRuXl4C1HdOeeokp
gQ6iLwlsFQ9Ax+/JEJJygfmnf01SN9uZgHLEW2Ub7TQb+NoL3UFWZe/RpsRbxZRo
OncCluJoCaGwsbWOGL2dokP2kbFlQiZU2qfUvPHq2Te7XK+MyOLZpf9djuAiKWXv
sNwhXlB3paOnQVjfdf0RgFcPIIum7lU1hSUc1+ZUQsfrT0qHXpHeFSY44q8e+/0L
rcT0b2MxzDTVP/QMgx+cZs9hMT6oU55ywZbGqblGutHHlhS6Ad2sEmWZ9fjl4HHX
a1cUuU5WosCnmhi17Ppi8Z8S84q9I4QEpjn293AWJ21E49rY5Bo+zQaLtAPQagWt
gkpsNrowzFDQII8J6Q1inH78X7Jdd1ss06fnn/yWhc/OXfSDe4Gm+AqUjy42qXdU
oAbH4+xUYyQdKfX2KVfngcn2YNoo/MRdRy3t8J5St29wgbBUgLLDFJU7tkEFrrqY
1hlHi8+602XU1A+rQor4AT4TV+kzuU61FaETUUXXLyJvE7xlwmd12c7zYUzuPjca
0yExkY0N6NBReL963LSeQtzIiEW5cchbVD7CqTIAszscdI2R4t40XfhV0Er0zj1H
EbI5qx65SJNgV4LAp8X2HGZu4W3/aneM49Qtb9r+EMIqklb/GIjyHSjXhchVJwDz
E97mow6ci6geDBciztb8hDXopXauYKNinYPQH0vvdGKpywzrYOvyDVcYSiZKSa39
f1TQ3IIVX14kRGeIKuqdiMLpPVOfCwlJr8nm8gsetBgYcM3mrO8r15CHo/UeHmkk
Ptm3jaLSKks0XuK6j0CacPQ35DCZCsccRkKrGtKWqPMH1fnr/s9UgBtVYUFlL2/I
jMyFBlAgqvFPmMNwGZkO2rqOT5nucdN4jODk3wjyyCL50GKnkJS4q+bQEY7HvZv5
TA1q9Ikl+3ZGF1hzYFf4BCOSqc0FvYhwkioa++NfT6WiGkmHZFLL+qlMX5MWJ7CF
4C6D8PvR5XJXBsDkrMefzMeSL3VxAduXcYIArC7Z7tN/9bpYM2xzhXi2CbZ5eyZ2
1hk2TVGb0i17c1eUTJjMNCaXfM5DRTWNmGHUNwYuyypmkpPwd3rjo4BaiNO3F6rt
URGnAjhXtRnZ2zKiX4rh7QD86jf6qN86XE75H6IrZ6iuRCTAxeKLb1KuHazkreSP
eTjyOLdSHYpx90YClJ0DFk7KwWS/P/xCboQtaq1DO0F1akP6/sa90GlEAFAFpZJE
F6qgJv6Xgv2wJRcKLrbfARZa863EH/MXoA5PYJ0uQzaNTq5W+AEr/9w46ZsqNjlf
lLIlA9muIdxSPinfkiTA4x+Tg+TE8SDj3ucwkehXrwK5zZro36XHX3AYINnl/Y6f
gOUGB2ctbCjEc2VdPMACQM2nzrv+4KPsPOR0q8i9M1ADihYHVuhEXHzjb/6HG8mT
bC742q7JPvoWHRoNFem0vPNse/T4X/ZHF8MO2pUhpiK5+V0NqrR/D7cMTksWKLS1
q02LgKBHkrYwuSRtKal4rnE8WxUy0gD4oAiIJw0prwmkLdYP8nqnwagOyXh++xve
iO7R4DDQGSIkPLnMtbJs2Yc1M25/EM+H9Lpe62Qdmo+QZTAqJyoo76l3EwTQJVdR
gwmvxxm1PaIw2PCL+2G4TySYJvRJ3ibomPwZIcZQpuuvjwnn80a/4q5SQTf+3dxU
pEF9EzAk5xSVH/g/IZvNx9KWshJrek50J6uzQ/Au+Wg2NBqtF7wMKeofUZEf7MyQ
nw+xmeKlvgrLs5+HsxjzddQTBDIC5RT2qsRDVxqCjXu9ygnHTV05hj3kAL7jt8zx
BttTGDHByFIYzkAB1fJ27Q7al7fdDGSqUDrnXdiL5z9jRNkdFZSNuxOyeG8kk9ni
IWgBF9RgtjJ1w0H/E4Asto3xBcQcO/Y0yjisuNYd8K6P8WDgcTHUFHeQwuK7FNoY
wPhg0KiUwrI3JGoMlgCQzm6rj8Wg+UgH1Cnxo34jdOkYBhyKhJl+VhaB3ARZNmue
oj9sO9PoN1tWrJCvd2VYiLdZ0IuCBKznogczQdrcbjLtOz+rqSgA2/+L4AAPKCv2
uupFW/RNMcQbW9sz4KVhpACnjjx1e4Z9pjKkREXSPP8qEzgVjpvl7gdjIwWyOzRT
qtMmT1eX7bTZt1QIr+eAoDLwiQBDacIsH5jUoc0lue/WOvlE/COgA9NOJ4X6e+3O
BI85qpE6/Ls9w5w/pzXS421QLAF/IyANwdwHgFltatnV8gtr8v+jwrfj+6wxWuIR
ayy+5CYPwWORxKvt1PITcdrBaVplJqJOslFmTwt3V96hLBru6jJJ3PxZs+70kunE
nJf9kxZbupcd92RZuk5l0NLSW6a4Cl+ztU2ywp35XIFH6EGAwkzcWNZ3y9Xsv5gy
TGv04ATSDyjF52mvTU1DDV8t84QcPWN0/wcf8XpguadPaJ4/4kTbhm81XyiCcZnr
kusGBWIOgdGjaLdGZgIg/COFbiqIUGa3VvtWKjcRlh5jYJtdASSgw6JVV93wyJfk
uYKZNQNYxUtimjZAg20Ogba4WzzrqeV5due7LoI28U642R/yvWLdUAbyKR67Ed5c
JJjtZ5VM43/RutnxWzj4+7348oYHcKQ0QbtNpHhybxvIr5PoHaKSH9fqJ0RmXFUp
q8uJKyLgSIR9mmq7JshwERk0yWdbMjf/0ULaZU7BwfRvkkUlNxz49UdnBhaE0U5r
DfM7OnIh3Dj87GUvg+ez7KoXUJNFPrfnJKEXX4kEOrJCRmk8YEAAm3Tl2iZmpE4+
ze8MhrqjShWPcyRgY9xXYTGQdZ/XsCASwJi5OmFgBmWe4pP9XKSQCTFBmMdVej8z
KkySIQ5GxNZon7sr5CdJq/7KjUBF8/6IgIFhzh8s2S6ittAY1uuYRhrQnqVEZKes
0hzQo9Z0U8kS8qIV9qASYOttifKmyjkDO5qX4Jf8GdH4rBGWjbzd7mcoo68u/Aee
OrDh4nQ1U9reRiqwpeDChXlp9OLixIpjUDm6JtgL4AGWO+PeFs4U8wyPhFTtMRUi
O/tEAnno7eY71qX2AGjGaj4CF9ufekeFnRldNw8nptPOmEH6oQEPxfrc6Dp1dn36
Sl3ou2KSobIeQbGpjIApgqytJq1yPKI8y0hOw1rBjK+CSucYxJSiB+iIf8GcpVdW
dr8OHOLa2r41TYtWlNaI4lv0cgpbiRvA6d5jqR/gCHXMnS/IbknJrDvH3LQWXJhy
qNH+FvluxpChKFMShsvWhl1atc7rdsix3Me1VTJljDHN3ZM6S0NC22puqmVXEc3U
IQ3pb+g9q8vhT9o+w8N8Bt+lMCKUjqyYId5loaFKh+jBxYm96D38SYWZ2aRUSxCR
O/5MceQEQ7FxM+Fkr6u7eSeK5NIBT84xfA7Df8AL8rpVwtzDL9Qs41ukYImSFSmr
YCSQNGv34MLfF3i3V0l2/jIwslLW0DaKllNiptezT7lFCVbIylHzWUAaW05jq1Nb
cowrdjvDCI9sdZtb2dRbZe3b3cXjVxzRA9HY95M/Z4wyRgorDiZT72bupQiE29wA
I47igMpLsW2657lki/LuT4h4LGbvkFW7jt3kPrLk5RbxA2lU3hJEnKtI8VfkVnfQ
2teqLynXyDT28+FVY5sA90iqF5tJjFCBLt8xUxwr9xIiYmNMLbaP/KOlkEZqsrkR
vcME9r6YzHTkyP9aEcMREAkiTlLW3/WuXqqXshJAJ0hX7OpCgJavmhbLRFUiSpYE
8vSa4APnojSg1tsNf47lKUMjVrUSmH0yoB8sSQq3iEEDQLqKh8NkioeLzru3PNLJ
yFqByNQcg9gUYYCfKJ9G3Pjil8CBHM65di2vsrbK2/NMuEmP5xHwHUVBMu+ftvBU
gdedMGXJ/ncRk7qxOq3N3BbgsgyxicY/C8tZ7xYKm9D69ekZ2YXG9zLg0iYKW2J3
cOlKAGgSiuX7T8GAiWMOYrf6cYh6wRiexleGbf4d+L/n3eand4ws65ZhJFZFCDeM
MADxX15ZOxZy66hng7VG9uCnorofTifvCbdLzxzHNRouuo2tJ57T+L6Es2o8Ppbz
4CezLl7S4GSDzo292B1F69OGcwyhl2FHkTlvffx/WKdNWmB5IZwcU6CWjvdR1ARL
FZeUAB8/Giz6dOqlsDzUIwqITpSzWwQ3Rye5KOyITD8t0iLxcO+5SkjIXF3O2r9H
MmEkkMKpaZc9IYhrv00p2WdKSzhHN8/OnEOcOrwCQmaqKWf0CqQCbkuAiDMgi9Tw
88cQuCQlDrqeZpqdk0Ke9tp/2UopgW+Dkz7mdq6urMi4r5soeGL1Iu6K7k6qcbSc
r8d7qt/Dw1t7emHFrL7uqs/IGtfjUsqlmPdergz6bsEBqNK2QqL2K67fJNYkIVdW
HwXwvcpU2jLUDw32UXXlOg7zpoywSyENRu/nWtj+3QKxOugg1I9wikBAwkn29KIU
W3LQRXcK6muVvrb2w3pIN8T1ev0vyQ4HD9/tU8vxz1MIHVMvhW4kRlyH5HAHPuAE
eal9QfkaP/+2yaPHSxriCPaV5WuRON1JxXyadrowyF3U5iqMmIDkMZjThpaGtLM3
HN+kDGCNWxmzZltWGPPTTWEV3roMog7WNdMwhCc0HTtVLMrTOGcT7QeOZsR61AT2
yqJ4wKvQMCbigkDSB/yXOmcaBWL/up9pvmYO5OYJHq5wt1BKbs4fKLd1KXBYSRAP
OQtyDAprG8Ff7yA53S+YIx0C10C9i5YzIVQihHR4msD0S63e7It42hwWfza7o97r
bBW+JKDyCUmJQDrSh2ZuFJS0wu/dieI2OiyUCrztIb8hmvrA0nth/h8EM8s1iD0H
ogCr1dXW/QDjuK/I4fk7nqE2I3a8R9D/0Fus8/Tev+82xuUY6FCjK8DSZKKbFatM
g0QhA1vdXRgY3cEnUzNyTJ99C4WCD8Mpm13zjzV42YQgmrGrmpFNd4V/p7PQLa2a
iBnP9gkM0RMHr517yV+3GPFGcGVzUoQGxtF3aiCSz6YsZ+OXpYyU+u34TBVhjy0X
QIVE1ysCOvYhaizepBelGiMwVaET2+hsksFtji8avO4S7zMQPCgOqBzYqSsSB2ES
EoW3OCBYmA1tFAj8L/v0V2zWxIosarqDW4K5/1AAwcl2dN8//IYRjgvuid7MFh47
H/gWO0sTaS6HtR3EnvD2FPFKozDcwVzQ9FPyQSiPuAfctY3wbrIjw77vHVQ5WfuR
+QrxXVqLSBYIpdRbbgKkKIcl4kGUdjcU2xd4uHGleE+LSoZ1Ra67zr90JqjamN2o
67DZG+De5sXdwLcpzmTYWZncERILpp2H9vNosHwDh7+NHmDI29MQ5wUXRc7Fd7D/
H6kSJInHQnIuAbaSpp2LrMp/+CMLQUIogNsgCX1miQFuVDe9YWr4NwkVZF6CSERS
nUOm6SkYbAiXdGVE5TZkC7cYE5IVA56w291EX3PW4d/Xgzm4mDl//TSlDuVaL/YH
oMLjuHvZihJ+/hJY+ohhSFNgVl5YSj9SVc0DUQ6FtO2+3nhQCF8s7DVN4FCGQ5c5
a3Ro8UC9rPwQMUsVAbVynIGyO45L/dsxd5ibpM3FXvaK1qfiWF3fvv8BvwZch2rK
odCWTsDEA+WwjApxwddsFjWtPVeMi6xAOA2qiYjJs85qwcKoX9+BLGog5F6xSg3e
9Pe0IMs9ce3CydvcvTfl7Vx7XbbXzpSX55KXL/YsO0vg6dRQbtxIMxy3HFgD/Ive
2t9Hx1H5hM1TNor2vQpGCg+whpJlpsuibK8U1UWPyiwW/At72d7pCxGSWmDgyHyM
KF0idf9Em7w2ebwjdeHGmLvE13SJSgrvU140nuLqAObfOTyP4fR4oT3EDL8KGrzX
PUesgp1kMnTO+oh9UdyUOxCLni8VXprAN320BwW1NRBflLA06M0pGFaQZ0sah0Bb
ARYV5eNAulGx/tal4wHf2CIxvIDIieFe9e+0ifBVboORGHnRXZv4uwWe5YDRmtLQ
uzOcBJfy2MgtPFGcpEVeNRZHHoK4Bkki4MrbGD8rpJDHHorogfWJbancb/97pyJE
AurKau3OZ+iYfHDQBENh/zT7mVU2sPxfQqDQU5NT/OgHtlVCXMgh/uOqBcC3D64l
HDji8xjeWaGaCQOjmBB921prziE46wMpOXoZFMqR+h+W8sSsz9eRHneA6bV66qsP
zkDBkaqjH45KSrs4C0eiKfJf1TJbjeB5fBmAUihCWjnUR1QMPkOFcvXFKEb1VT21
zvwWb/yPsE7wWkBLR5hRItHQ25m4ieao0k0POLAIvSJLq86+4h9I1tG4fy592UOU
sN2SoEfEzjbsorDUmNLmULkDALTQzlauzRoUFKkJ1/QLYcCZRrrjQJeuRNfhD9gB
dbd1RyUpMFQvdvDjIOn7FaWg7ufJbWEweUpzbrxPArqYXzKlnvYo+tIyMD9/HdUc
vSnEIxaN6Y0olftSpDGfHkotjjOcZAOLraYTynC6nyqbuFrMrpHmgFHMPoGYdRpd
6eNYFA7D09dCTyw58oXesj81JHx4x7aMJm1EIA7OqDTe/YnvQbtHNVmn/mZUfU4l
w5j9UjQYl/tRZMWlIJ3OTyrWUjYGr4KFj0dxGF3NH37yJAvhrNj450gIoblIQ5fk
1JakuDRbhAov+AE8mGwc3ZH8y1ctLTCk+WrOh67h2GRBQNzNDVNDAHVsp7O+VGWo
KcVg2DvDJW1M5o5zqL07xeOv8tIc+0wEiyy3zceFmeLQpY7O4I/EA9gQKFV+smvT
vNIyEMhU30dxmS0lJhoiCJINbELINTOwR6ktM76th3NATMqOXb6rkncol3UxXPDO
wyNCBhiFWyZXx/1CV6J/4ke3UvPPD4W9PBfjQnVMZBB9XyTQvaDDusBzrfe9SdGn
TrXyL1hBDAt1mkak8NXowUCG2J0B/Dw/KZbJNf21mCFe724hwtwfMECVoRrlPwqh
FrzisF/rYUM+Y98qlXCY9v54az1SzjiXIdTEWRQ1dJx7JKmUnGbkmBfDeh1WywNe
zuT9vxu0//16x3KcTuZOJn7LPHbLI/LrQMTXCJEd8r8RDZOP8ElCNYcZ8leaONUO
arIIkKIr8cnCOwcC6EVwBxVHgZXXUcz0et1WYseYeLgcrBJrg71k2n3RQTwtJ5T9
Uw3cb7ENNtfszGes1YW2JfvjTCglgh/p0hVibnCyJW3sQIBJ1BaihU9J1/M9mmdV
OPV44XbHkNaGwp8mfjwNTA3FiJrJUXYN+oJQyZQynMu2VopYijizB44ooU1JeASP
nVcrTz1rZB5f3y+iAh81m75jVlO3lwGgD84Vw07TKgrJSNA5DvarIKBAFRPggjDl
bD+TzQhlNGYS+c6I+QX0TESP63EoF+kwuJP7krsZ5d9n5H4dBaij6Nmxi+pPj2xB
sb9pZSzWiqQ4e3xVQ2wfEJfpisQfSFsd5a9D3mPrNlJjJGznXj9mYeEFFDTKLrrG
RUW3+4QJjb37TL8bfBPUcjMWDjCbaBceaDho8p9mhi1u3HAqI6wSp79KhCN/INMV
WS0Aop3yHOeAHDkr3IOBFzxNbe5Q9J6Q2yMWMdNehMZS96jGoyf5dxkWRZeWyuUa
g/qfjRzEtDOegRRL2Y9U9RVwR4R+t0YN7E37/+h6Ck61tzIfZRpOsrfr0sViWUj/
ZiNtqckc3L7zk6IEcohxmfNrLj/0H6EtOWVl7zUGdYtnyCSavBH/JyezC2Aa93+K
FUasoaeDgvvBhyp/00Ix90r/N1RrTDksE/c5gGaTxNB3zyfhV3OL//RJaUE+usEb
9WnVTMhY2nqGn/4g7NBnIJZh0PIJYQhiIrNyXyJUkVBYBZuuU7b2FaDDRj002YEx
a0rIRFs9cgXWdCuvmpwW1CPVOPBYkiNSI3yA229KXWjvGvQWIhrc+KDCZ+kzrCfY
CS7EF/ADPyXDNImdMRdPSwG00o+Mq7c4DVHM5t8fsV9ni4f+Y3ILSnQ/VjVkEYux
51ikfAGyvvdtiBd0j3wQtRgBrQ7RZxgQkCO7f2laBV6sYAgH/jkU9ZMTHXtgTnBe
Xa3HDiW8ESnu/GYQl9L+Fqs7Wdlgts4dxAarHtACfIgB1ZzUGMtnSFIKyxrQnLke
1r9mUjkbTTfAd03hTBbZUAxBuInAD8jdkIjOLq1MbdCEz2NikgRR3iR9ovDCS0/b
SGEYSBBuqxx0fEPEemXSCT7Gp6vk/NdBvckTxmRahTdptnATg13j5Rt/+CTpCGwr
WrDXkMv9tmZodrxAEhVxZYXWIyi2FmXivaBnyvBxRCXFoXTAXixUc48Kaha5j7fA
poo/pWvFo1z3tSO1bU9rGj/tmdXTEl0bm7OsMizgss135S6GcVcWZQFmGCv7+avB
XldSbpSuvMjeO4Z9VCca8tD4+9WWuhpz6Ir0qxMfpvUeVvepsDNUnrmgXqb9DLXy
p4mJeYORnWQSqKvms4TyCrSMpPQZZElloTXva9sbLEdt7oGsNgAuKfwNQ3CaEUQH
w8TdOrUrSj2VekdCpNuurAQz6e+2xvfhTbbjc43jPWPr1OW9QTnez/fNFiO2IMBe
qfwgjcmO1+zr6BCD+M/e5bRgE3ILBYao6SR2NFQUNtNbXpIN6oD3EilLgF0tg3Gr
sWgDD0Reexcw9iuZf1FBQj4W/iCRQ1CsloQeGUNTF3xdDEGe++WXN1Y6KmuMifNj
mB65U+1d+B0x0kVO1Ln++etF9AONQgvKh5dQeHajLnsXYHYBWjT5U2PsAbLcH8qi
OQAc+pVx4YvPF7gFRh8WX2i179+s6G5W+PgfZePFiGiABkLbqLul6hr849jnYNzO
IaHEEL+zHRgGootnz8Zuv3XlstfIKM1ubkigIRh6rIsaxlXOfnKM+1h2DwgdgnLr
fKbqVfJKuBnZnnQiqbnoOrohDidtkr74mgVF5nGHIs0Ds4swy5YOXL7buQcNP6xT
jmOEbMWpHaV6RIBinqlqEFAvpWJirzihSzpUle5NSBYGkr7+prm9wvOkFsfbx0jq
iRDoufiveaIkxoBeEQdef3H2fmDG4FXWbfHVirX+AQYqHFsVmwOqc0xkPeMX0Nzm
tXEXwgL2Rk00Vb/AWdYi1PhEgIaX4DW/y81sz+0ixUvnqySKAUeTmHxIEFeMUkaW
kWD0NNgU0PtAEn7HgFU7eR815uMXzuwUcmgxqsRKZB/SnBaYqEUfDLGr5yyAi/Nq
8UHzDrIfjK+/eglQym4HOTM+ZsK/rWa4jTpseLP3qhD1hpT2IJfvhZ7jPajM56x8
wiVUIpBjLEFyYBrwIKlxOSz/7FZ1MNIkDPVcAS+YwU07dXnPztfrBpfOfJAQl+xN
6kWQLFJ3YHB2zmkT2klnSG2339FIVLh+v4r/KrM99h9NpSJTXRxvzqqHgu4kSKQX
e/acDHAFyrTWCt9Bm1i8lZmwjpLJc3Q6d3P9+lIQ3eC/48sKdLFteJz7BsPQgodx
nIz6e8+wuSr8e7IIFdEi+z66IIRG19azuX5F5hrFz2tkj1gu+rXFJ7RJAMPEWKbm
PNfu7nclg6+ZmOwonWdGzys6Ppyu6EG1EdUQKIqAPc0LBgl46xjvTG7tqmVjOHdt
W3YOSVE7Sd2PB2GNL/z9cTbrJBru5PUdNZPm4SzwX9UOjyvkoRI7iKc8BjNNE8ZH
G6snCENnPK4G5Xv8J+8uhmINbbjljO9+eW85XXdgGM7pHjUpfjPU93veB3XdyVDW
bpm9Pv88ZGupYRhwFQXQ7CRJeDQAdPpb2J24Bw3ZNZmU5iSefTyx+vLb4+VgZj43
Sg7lhW0JuAyFz/ZyF5yGzFuChKdqflngeCSDUTN9edqkKW8517I50ppR1wK4NIqn
dfGUFx0LAwfBx7k5J0IFbrJRLspNcm99Fxczyh6qLcT9jBvliDAsf4NiJ0hIE5Zu
7r3gJ7uX1aTzN8ntBykItaQ13MmYyx0W164JeloiFAYjKm6qTMPewvzo5r3XHZIV
GXFKhCzsIpHASvzpxxaJYux1LTB3tKemd5zO/lQz8WpuI5OKfO7VENCkoO0F4Jvs
IvqmXhnDei0jaIlJkFeEQ97ST6NaRmitwsEM1KOqPanycwbkMEhO4stDyrPExeTs
ka35Vxl0o55zzYwgcvG6MkdHR28JZkJRj9CwWP9bSoSyQVhboHB4CmqcQtVDNazm
FEkOGTky/ktKw/2KXmDZq9v2tZlK7aRg+B/ao+Oo4nh4sGl4rmIvj2LhL14D9C3q
XPuEmpPEF/RCNlmC3wfC8loD6j00GL6fQQM7Mm1ky6ee64rlmKj/29pK2uILmt7z
VHKDO1laVpYRApm/LiT4Wg+pBO4cYlBYzGn3MVRVvGAQaBqB86dLj39Ht0CmPqve
muUiJScAB5RoX7x/It1DExgfN+ILP0ipsOElGP07UntUVo4jvoTsTBWf0eDgFLJq
BbLejbIAwjqXrlO7s+KpTdG9FdDCa20XzYF8BlhmtXT61JfiD8UAvKJprKXProv+
UrRQ1EPl60Eff9vB36WAAInqBkqHHyLg5hRZ4LIMDfqwsMbaKIhSB63IV8e5dZrt
bhDZvFJxuSHdbguJMWH5swromIfpZ81s/i7f5fTalaw2pYz45vX7ctWZILgVj6Q+
l4ShXWuLd5hwtAAk5rabnF0AZDa6BUUIlKyaQrwREOlVIAL6XgAK4Ec5T4XD4YlN
00bx8trWGtF0MVty5TPqOq3dcyTQt1jfX6JuDT6Ctli8gF46ORBM0TDWpteBKWt3
Og/50aOr0y95mnHetZyVPPWS3LQAQvOFG/4cp/Aqv8+4sUtF7ZQbpEx2V8vYCG9R
/DwyHe7jkGg9P4sAT21KAjnCVou+zmsiiVBhi13Kn7wF3xffTBw3Mq70tC8k5Lhp
MF1RmLho3PuxnWr50WdRvoqWeAsVSrwZhQVpAJJHzpyy0bs054MAs6XS8Blz8w/8
18f4yKjpFvWITtNZBaL3fnJgBkaAaIQE5QA4YRfoGIklWxkIK7x8nrdzeiyeE/wJ
ATPv6QclZRsr0GouUnV5Ok9G/fTNhm5Dy7Y6YVfbaSgmqCU43Vbb5uQ8EzzZByTV
nc+NbpqMZ8M0cUGEkzf0YQB98cJV6EDKf04IrnDPSMgMoXrit9QxJBuypEl0WbzJ
JQ0RKp1qswk7ZPWHQ/0fQYHez7UBX3EPZICYnbp6HPWqoV6rV1wV6hQJ2tjulp/j
mhzgmSF1da8AAZTj5fEcYDQXWjlxHm82CSOHp+3a1++4j4CCx0iOryTvks8b0Q4N
l4EpB+1iVKGldZN1F6Jr5RT5UIvgxjbyOAN5XtMA7XoUlOnFXatsPsn6vTbaO94k
dyifmBhdhQdHdZIDoTRceTqzoFDYJS+KDVQvF17nyzcbGSx/Bq6RYx1cWY9E3QbN
32wogUld5s6qRb9JG/9StpmKx5o3uZLPr3SGXLhh3xkxKUz456Ik/AUO0iVGQkgT
4vHCMv8Qgo7vUmBtniEXu4JlaKEERukoZKzWPeWcZ6pxKoJJZhvDqv1qWGytwC+b
RRiDngBpQnoqeT7dhAXYhVH+qdxbN1flRRzHAeu4i5syzmpM6CWRSpV6adtBYaPB
lEOWSpqlI/42na+DQBdn+7HBp5cz+uje3Ql/3eC4SrgBYEinht2ZCozwxdpwg/YB
2O09k1K9fhTdwJvkVl3rd5mn5l3TBHLiUaO+jAHtHux+OjY01qwMza9kV31KuwdH
VQjg2m8zJRymgU3pMKaI4OkcQ4SJ562MypTbjficfX6siuGAl6VjE68140wDjHla
z7S03usGELyRNfckODu9fIMsbrS/D1/uBI40LM8lO3UPNeEErYG7QSfQrV0BGs2q
hQLGYUNRTgtlniJOEZNvVn5dSc76Kdwtfm5miST2Nt/4Pj1pfw7MprhIeA5fdxNC
PsJELpOa0q13mhY42h6pFTA2mDGwyUwAtBDR314pUgeh5TbydSTSLJK13biPjU0H
EEj3DqnXCQcK/wuWdtt9gf1onpDi5Ff26pZA1erbDspBFcgZkA6uZtM7xypQZURO
gLLtUSrfVDNVvW4LHTNF98u3EoIPnVVIFpOcxWcF/eIa6qtke40Nuh7vWvUAy3wk
KCHMl3o+9R4gj7koTkhEejEaQf2Sz683ntoMhQsw8xf4cwnHJCKxn0ozmWG6fPkQ
afaIV+hA0rhmwGprVmNc/HqpHn8e2J8YdXYwgdF1XPBVeYIltPQu1WLsVbT+JY61
tvrqSBC2raK2/f8kqblVMdAajli2GnzfNOwvCNRheawW1TGrH7JNY3W0AcMYH92I
Lp4CUmu8a2YTEFsQz5CKVF0fT0xZ7a8VEXP3bvBrYnJWeahUCfAkbBH4Lqhixs5b
n5RtJ73CPSsn0WdegD3X9Ufj2NblpyyshdswFQtT9zvnkRfiUVuCg/Xyf6F3/c1i
4vJVc5Ud6oo4RjX9vJhDspSULKA3ETtM0ENqrDoCfOt2cmeqArktwDAt2nQPElCQ
99C5PxLz98zOoCnXYsen+J6e692kDKyCWLyPPPB7+ZA0KxkQhzf8wo6RrHROgLdz
lo9SFQrKRbbKyXFl/emVB8PhGws2VfSwtv2DDKM6nGej0ycPLslJVoDNL+zst3Ev
kTYG+0SZ6SSyOwdEYbuDEh2drvdjEQuzlY9aFsI9rtEBDkUYOUvclFzQY4mCj6zr
ddWtcnrRf3RS/zcHSxDSBB8bN/0aLCk1Vz682jBB0urUxqgVMPjuF9YI1AAJjEpj
Brt9zOX6mFhZ9/VVilSveoDmuxdgAUnLVxK0zVvN+j+XOYLjno6ClPxn3YxsM9g3
y4af8oWpVzyTr4LlKIpLTmFN+dOrPV22ipBnN9PTit/d68jwhYrBG7RW+gHKZndO
WV5CFrTOQoHbX4VGB0kBUWN5f5dO2KkP0SbEYfHlgUmAYT+jDHRpMq7mFQ2ljbPb
oqAOy4yKThBdrQENgI3TEw1qQ9Bd4uyhH5hFYfMRtmDM+v2wV9E0Rx/Va5RHnZ11
XplCnpa+nUM9dd0eMWLqSg26dxG3GzeybruxfVEJclVxowEzs4OVoQOxze4OwcaZ
ejiaiXoVpnuIRR3ngbsQyxSER986wWZZHmUOx7MVXOHc+9anhy8tulz+KCtZm0iD
ZiI8NNyr8ZkrGiYoyCMdvSGstEva6Zc/A4GkJINDQ/37htBPz05J+7jnEm7p0DKr
eci7V6jwFFpm0C9mTfWrmZeKcZ0ehSLhZeKAMKd9rmpyHccl8Kp9lna4FGCsJCEQ
G70JIxdok2lXR7hscU1n0+MKEBEdZaWXO2Mei498Bbjt/azqViVzWoSBWtTs0P2j
PNYtDk92dlLEIPsejqI5Sdgx/TbdnGxZOVnasav4HeMJ7+HtTwD62XsZZj89X2Ch
Q9KdNqczQviwFLWiNICFCYAemU/rChcUxyPvQLlGBUd9WhM8vCjPuT9pRWpaG8YJ
0hNxaROWlkjH3Ig5EmLVVcg1n97JaNWQxoG4+8IrpTyi1CsCoOpGNievkz3vZbEk
vYMRBmrKkA3IvyU8lq6l1SIwvZQrYfo7Ia+Knl3ZuDHC/79i/aYVxKblOaE+iuB0
oe0glzLUuDCcbRaeXy4U123bFKvC0PELpPpvb31RLpuzjJ35qVFPBohH6hbbRIkQ
awEfp8L6pluFZVnjFbi2FlzgiyJq9nn7WU2G7SWAJN+9mnmAFgOmghA+blflaW78
0/wq69qcRqQNaLb0RIC0UX9Gn5CLpO2srC1hJUU4fDuSI7SH161dx+S6pCzlMNpb
ArJwQY+hudLFTm0Ox427qZvBpx0w7O6Ysd9/t0AeljbVCyVo0+nLypNob0OLQY2S
EcC46Hc40Z+PMdumE3uR7pJGg7LdoEZzSmiAglhawWzVxtn+Pc6Cf30PWC4vSUH+
2a+HcSPsY7jL9oo//E3zh+xeGUF5bEGMP7N512J9JK2+0p9Y7NV+dm69cV9UmFnY
a4+YsXdTnakqU4Ya5apomg/17e9TLnmPB53Crhnpuomse4a/x2+TtQJ1mGjbkfKt
UgsXkOXYsnp8aPLPHZD7cgt2mcaPlHwDbiCGzDaJTCZYIYFySysRK1AqegGCK4pW
R8KzVm6sHSdim+lbN1txQ6X5Dfpd0X7K/4I3LIyFXqU3uDwwlpAlPdOa8yHIcx1y
agtHPEdXduw9pWKq5z3479HxM4YgqNpul05J9nEHIcptxMcYSiWbqz2YPRLTltfD
pGmwemHH2vP8cbd+R0CDFy5jVpn169umy//bkhMpFfoLiki3QHqptGeRYOyZJiL0
0ASCK48kwvpYKgRxFooki7ooiG+L/l8tYL400AOZlgC1qsxdG5g+FQ5sglthsbPs
ooTLw/F7zEQgHvd/LsRVFhNfMT1X41GgYXhMCAlYR4V/y+xCMo5Kcr+akmCpXkI5
kVLN8fPATMyyILnBztxRQulyf5fVkv8oQupZq+X7+AweN0eB77rU3Y1Q3T+mASaO
NGqB0kakyvea2m528OzHs9Z8vrCCvMTUJoGWNF9+XVVWOwjvu46dTbAZzL7tdu8e
eE07l/HUshltNqyj/mNJbmWVmJYRb58owrK/179Byb0dlYmpBZo8BWTfT2H+gIVR
ubE76gwk0raE7FK7Y7q8D+8FcZSt8g2xnbbGpqznzMvSo4dYlf20RyONbyCEMeKG
G0TFvD9Q/5nE+dY4ATQTYoOSQIbIVMKEF9rfRh7/+Rex1jnumSR5Z52ofqhyz9Co
MQ4oGCe2udUbpHbUIi7wRQERkh2E91eaxmf0INmuKkD6OBv+FExRE2gZp7teSbMw
50VBVjKIKom/Ha6rQ0QULMs7oDF+qvt2XQd7Qh2V7AsnpfvLtbNEAjsi6zvWJu6E
l/zdGz4j5B4yoPh7jK1IvgNrO1V1JLVFGMrizp2DWQa2XsWv4igFuPSbDzrT4ux3
cFVFE6pYQUaQI9AycErrM2SJ6lQRr/uIsPSwlYno7LayHidghEAnReOW/ajXc+Ml
1omA6nCupSH9j+X7iYKJmZIiaxADBkzva90A7UD+ab7bjVclqiJW0XcJkivMTKDi
3dBwr6KgT0K83hegFPlEaLgfpM1bWTkz0jXlsYjVp3w3Xk18yucs6CAODqG0kk9Q
1bkKxhoxQKNKaRTA0VqJgI4jet7G2QFL4hR3Hx3RE6AhJefpWh8vJz8Kx2xAg41V
Jpd6UNTr0ERjHiUqOsXPxI8b1kXvjbmYCIIAxlle09ARTnzHDwqFDy9dmHSrLmAX
ea0sTkMVuboI4aYjXduumHECwOww4yA7nabyTmz//Abxq7yzkuqdX9rkVQlueJrO
0Rysxh6YYKaUsWERL2Bwpk4gQTUt5cgs2T/uRD3TzRKfvE7bBH6zDHGqpCVaYpmK
oVz9leGgN3IsL+vvGKo0wYWVUNDYJhVYdvJVGtS/uJRaC+LFNaxRP0xMPTsBCgRN
PF91mtej3KmQE+KG3CNGQHTZFiUwa/nXfh9us6OP31g/jPZeQCX9MeWY1sX8GJMT
+133bluQrQs/z4BT6SNHR0rdEML70nol6+MrqCD7GtpmFIv62lll4vtE8Ji1/snT
ZAW31agXH7IX2wJbf3erzN1uPpAmVan92ARF3WLXugIM2+LEKd2KMcdz1Gjp9ylK
/hDmrGCVUDnU1ztPDUZtGz682icYxs8izZcy+7liuOJ0OBBMmVSxBVnDa4gD22uK
s+fLcYmK5ZAVyE+oqg9+kUeZD1LEp5Ltr9GNVVf9zkvf7gIAY4Ab71ea/cjJfu97
m5iSUAK6vGQShrRqYSan9PZ8PCkcjY8bhkp9B1oR5UmB5NLAie1DB6BXIioPn/on
MiAGpt6lXVRZ6nlZWHQA/7egzo3bEzAQlg5mfYeRtuHfY51Z1tcpp0z+uX2R3Si6
zB7M45Wg2nU53BhRT4CrczwGi5M3cE7NSbDJAC1vo3YoRPp7LgRMwTHZ6ibIpxCj
O0+PktBFbMq90UGJmrJ9aA9y2V6JYEDPOKcdqGDkJLrKzsDiLXkKnhf5PbyzbvE0
QMgHB8tbuK4Ma3lqYfp16gC25k1F/HmY2udZqS43Db07EywVF00N9hW5mrAjIiZ5
zhKiwVbeoxzYGqvp+3jr4d+O3vR4WBj9UXxtVwrhewOtyRtetK95pq3Mqo5oD6Yu
h0WZQLLuP5ySBtbEX7c2aicDpCgaUalUANACPmWA+AMmuI49DiYgMJNhxRXsOL6q
biSZ90NvESLb+SIKvPa650bUnCWP+PO7SpASYQ2rm7ni09oPUMNyblwhd1NDB1Lj
9Y8IvOfJJpAgYYWl05ZPEIe1Zoi2EC53X0x3v6UHChqg21thbKrU/jHTM5mgKAtu
AS4wdF8JfoWxPzxw3cpbdzdwNGSboD30Us+F0y9YQX7lqi9zi19D4yPJOiUYRiNj
lcegfq+oVY6OKV+gusZ2ZOsVAdA36vOLjEapzrXuiTAUeIFS8Xkw2r6yMPRGBYPn
JmqgGiLS5PfpYRJvvePUnzMMQo2ye1IFTGp7vqNG/nKwD4hs9mQXT3zueSw8MMm0
L4HtqQp3Y/1ZARnj6uPDRFJr4H2wPwXvrPKb2axjo9DEJoHwlK4KWW/amVtZTHeP
BYXDjUkmPJyA0CJVv7V4uM01zbh7ewhKYRJjuSkwrnz0hUjXyAII1udQ8KbjKNeP
aGUPbKwi6ETe9YikO5ZcIQKU0V2K/LZSnaxy/1JtRZw5SAPOhNOTEILQ4vIv3AJh
xeZvBZxfyC8/CYmCDEjGbG9Kr6eSHrkVahYjDgQhRhNyWxr4S/9Uugin6mxlNxKI
Iq1jjnyGmfEAVhEEVxPFrmIPdD/U/tLdc59jDHSdE6S+Xto4Jp7bwFsqnRarV9pI
PjOIf1jw4NGp2PAq7BpDAHfNs+cFrGFSXBQsiKOb5jXhHUHHqTRUorQV289gRbke
1+ltnEXb9d/zvCuj6TKvvUeQlujHfJNSrVmvYoRIwwifEs8FCWx99dt/jJAetRAR
4Mqq4cKUalv3waYf9s4+lqiQf9qYpK6M7wSs0ymgML0xQmfEdu6mneDhgGy5n5ii
ZTWgY0dhdVB16MBzQzsBpLhWUGl7b7JXCGmrU2RySlZsFpgzsLME/IoZWvMnmkd+
EyBtpfs7F+5e8ZJG0/fRqVU8/epppzRjh3pkHc9qe5o2mwn9k0/UzdJhY4Oil4KI
JYtsCcqHsrkHFBD73LTfeNuaEjuIxh+kAFKKpGcRzoYN4mkmCswRFASc5H0VGhD0
DedDNUT2gCyWCcgCmxQBCBa4O07CgS+72ASGLp3vBsdvp/7+sxlmV15sGEHyVYAh
Ms9yxDLEaQIFVi3MaFYAA+d9oR6qqloadrMFm899Izf6/J8dAbLxQlOrTNozAEvZ
Xwp/DQJUzXn1oAbqjnonuZuqz2/j+GSMwFJ1msVbd4ENpHLCQ46GgJO8oEomt/X9
hal4V7gX0JKf4RFqXukNKZkcs7Eg6H7USF62gcZLn08NI50F/q3LggruVX/XXeir
5r0WhdhbNeCia8UowquprLGSNrJefN8hAh2UqLwV1NFkXtOuMLqPvN4w8Q/9HC3i
15Xu/jGn9sM1vDUEeWB+4o201nVes2CzGipX8hHfPOiSKVzMWIUKDlcEid5LKARa
tCCBysYlkgNoLGoPU7uEy8Kq6UyZExvE54uzdthYrITNUpPAU6/WHKO0QD/KIXPJ
D32QONKfgC1oxy1hyyOq/nChnZpMG5NJNjGoptNwyDT9XlTszbicP8/In0789O9d
fWm08xjGMnRj4a4rZn4DPauH0AV24pv6+/JAb0RQBYN31yCjTzW9QTfJgllrNoki
qFoPYxabTdSvr+/QV4RTV4V0vD8esJ+Gzi77hAyqz2e1YT1HO7nvjD3CwD1ylcUf
aA4hbo+Wk0kVAcQwDP2Nm+CJIzNW5GPNR/BSP8mqgLSo0EPZwBax2eXUWTdUgcUg
OUCPRAjH8/RqOYQ0K5Oy+I2hh31VX1Jvt9oIbd6es5T0OGukrLpVJtZZLvbJOtGN
frio864iOxD2HDhoW+eDGk28zGahKJVSSEj7f4aBWc9MvlhM2k6nfK7jctO5sfna
/6kinCXP0v2avP8xcR3PaaABHq+8SuaEuTwyyhJZ6VPuY5NROiiuJLvPE6UrBTAc
0B4dtpTYZ9lKrLaprZhN/vNGeZSZ6ynUQ7y1X4CIuwKpEkWdrH+B44RZ2hlfYEmn
Kl7bZDf3Brh4LwAfg3KVeaBJ5U5T72wKhXirpcniSdoXC7zKy7/Aq4VmmB2zqvSQ
0xMJpT78BPfoJmnB0oMhxud/C2elfRxJREMmnWb8RmIflbECENboSiSVG1yuLEu+
n4gXNFCMOkmBPU3DT3OGSYB1+eQ5jVuy9G4tUOYREwhiTeDdj/yFdVyoi9nR81pu
XVtNfmi5XxZxW4ETAjEbbDshcPAnyY+yZOmEsQiFq847aTA72cdSc4vUkugiW3UI
Is27rp1gqauEysjN8Jl6b4Nz8pyURteBaQQcm83Spoh6VYCbJBvQk1yiRTZ8GZzr
8ecPuziuOoUCtAaG9CpNi/6gGYRSwjDzFbwibJVu+8n8p8B4PVPBXgz5x03jK4p2
NsK4QGp8Ii39asB3FViTbu363LQyvvrbjVPc9Lu0M0B872UM7fLLAOlIJvyfi1Zb
mGdSmrWbh2pKgALvEmL1Vd+//kNCXAtGB1BN1TXMw69DXiYI2MxXS/6R/4IqEwqd
ehIwqe5oU9LYJw2JzKPyrlg8HWi0Cv31TwnpBLFX1PMIL2NPji/79JJt8KUv1KeR
UtchJ5IySeESqIIaOUo9c+c6+SVeFnxSru/XerENI+W/9b2xmTbvI+wJHsVl8o26
OKCHIB++NbBWei8LA/a3tUCfFGsD0pPr2wwVfIThtjyqVIwFfNfrvCQL8RdstQlR
IEK8p8kxuIsu7jXl8hFBB7kkZ4IO/+gXNwsw9nsC/zr1/itmDJs6ClronSlBEpAx
SEIMoKy/4/EGZw1RAT2wKl7i/IwmCNsNvQwUYVAIoyZVD6TeksM1MV61P55U9mWV
vg/qWGQZH2aP/UdEQ2fViVtWS9aQpT07ym5x6Ihd5oojkckJi0sTQtWDlc72wcxv
nZ5iGSX9H416FNQoDZWyeT4bPMXoTRjAOGDLCpquIiiYs0XFPDw2CC2CUI5MNVSB
33YNYwBQERA2WstvrWY3/Fz0Aq33/2t+EoiWI15h/paRRqXHUmRbQcHN0ENQCBLu
PyE92oQluI5yKpDLY88Zc7l46RfvaiWPnmXqza2sMlxRKtD3wbeUJpxp/N7n9ubK
NPDAtZhpQKVrQSyk98D/KKmHKKHOoiw9a81pharWdaNIjByObG5azBWTq8kQCDbI
qpFiu+VDvQe7ZKWTyip4Uhgj5Q/sdH3yWzPDNSJsIKEQ+t3wfoNO1AjZRwm/D4NT
PNdA6g6phqIMj2jIVPTjRKwkN/D+tw579f04ojF0MhrOe7sqpSvgSSOKJ0YYCgwO
O8tbOhl0U/+r49UR1fbEvhQiFNFO5VTRT6SaqLfkC+uMrlLvJdYnUJntt4oB4pUa
sQP/rNdat5muPm9TTraxjV3aGg3AOXd96PjJdvmYvE7HpswKF/A/OyeCYq5b0o8d
RbvjlKIJzpB4/cYFPCMvgWidipMLcR1v69rcfEnIjC4uPGOx/vhS894oUejWEsVz
7bPvQqJCUlHSTDvRX+7M3XXCfMUHkjsHDfsKYYhPCUDEddlwogP1SlWQZjDVedFA
2P7aQq8iaapfnhZ8hR3DIQJ+PSq//+97feU8eCQYBBbmnG6AYeqLjXCeeDvF4G3e
0qTnCFll4y+EaUYifZGxqCnQj0Mewme20dNOXWWv5rNdQRlZuG+GPZdNqxpwhkhQ
AmXebAaS1BVAYwUV1G3dCnCUKP3UarDhNF3qg129DTfv9vaLCaW1NwNeT8mOow0X
yRlRRZKMeiFWXDTaTDS9h/sENvlSSagxKamnOmUrpp1XZGsmcHhbxWeKYfXcVjQt
ztel+NyN7zySUaPo7bVK/ekNWkJtWIsSdIwIANc1xr7dKGgNZ2d5xId2kWv6AONj
KEGxVCoHbN9lXgPw3TMJfLnqi6mihGZBBPF+oPh6kJoh5eSHVpJiKfyWdqpFx9eP
3miCRqlc22PNSYzrdrgj4PVeA2q1WGQvLnAnQNjASmPRVcdCmMWP7E2yO4b9LApp
3kDk9NNCY3lbV+FN8/LyeYP9bKi4ma1fJp56g5A77O8RbrYo9yolKCSCmNWgf+gb
bF1Fo/Yd5ej18A1z0OPMbYyC4qH7F0ldf4uevkTa2RUgqLcJYyCR/p5RMHeoQ4gb
h4PaLVv4glOt59Z/QHvpfcTTlA1YJR74ndgZ2Pq8zoOcbbH4CEY7b5RUHmmoIAZw
XcldL1ZfIh3uzPpGp+xOtwqi2c1IG0v9DoTmq4i1k59CVN+mHCOVCIGfgmlSFz3t
dm3FM/1McCg9OhiQret9Uh4VwVFWhH8pL9rnH9QM1ey1c6oJz993IljAY3aVv85v
znReedaqU87THlVYCjqiWiv5iiJJMYBOgdrIYu5n4V0zRWxke7sdWUHYtC2D9bXc
3LzTlDn9CKZfiLCh5epx+ovOh/rN4EaI0+ezFhuTeuaFScNWhuH4HCFNaXoLFJFt
rFhJJscmsY4NocBN/TyEKwgvFDVZfYTnyonl6vfsdDIev5XUldkXDe8l4hsbCTwx
bpNPOGFajhXE+nTe93bufOPNMUKutiKTumhC0TAuVgIgCsrJ7jWOfwztm4751jdt
muCe+wu3o12C5PbF1+gRHKNaXhcIXDztHf1exUBqf3BY29hozD6LujD9EaGGrUlL
pOX4XVHiM74pZWU3YnjWfEegFUAW9csqNhkNCeXF7j9ypIED5Hh7lM6tzRMYprFM
Ys1MMkkcTg1Ro3au6KYSPJ8C2JskghrkpdLI6OUb91hZZZAW86F2J1pc0Pvqel+K
tPjuvvsLtiajamMmaXXwtJE34SIf4YU8ZtRsIU0Evm2xQN3+kxjiIAM+X+xl9iYb
nOTz5liI8BHYJkCVZ7hX09VB5CV0SZH1DkTd1vYDBZrzfnwhUqC1Bw5MpfggBtbp
PkSPa74hpg/lkyMFArYl58UuHJQ+Wn5BLed3YgNWXiLPeoVgGMedbNiY9SR0TcgN
8zhKjPodWTMMGMCmfgv8Ryf8qJNlM2ATTGxMb4vlb9KQHNDTMEXAQSxd9zR7tv99
rJvevM5ECOAXebbc9+uVMMEKh5vIda+9gorFKseH+3EXe5OfXqhm/ubnexiLs6fE
PhrJnbrZEFSbIl8Njpczs5wTYL+bdQ0/qHKpDhx1q2AS4L0v9KWZOeWmfFMosEDw
p7UwZFaA7mbcIS4+KzL/11KLHIUonFHFdlGqJWR6AZFy8Bb04iqxZG6SmYrsi0cY
fuoXsfViuOkzvraG2DVxU36r80Q4KnOa8cMzCBYmmjdfiDgwGJ2Wtdil17dAdhI+
9sOCaC9rs6UdUbtG0S8KXCZ101NkvrKj4xYUamnLDPvRDDWr6lRuNt1+AJbQzxLj
91hhADBqSR+73Aj26T9xEJwR6rQw01TCGJGG+xOgRGejtAolrwrhzx8K9wGBSswp
3M899T0fVrERVuKwtY3U5noSTRAMS8uNhB8Tei5JrD1FiN4YFpaa6AlcQ2+ujkUn
fIxt/veqRh/jSis8kzhFGPbezUbavpA4FLDvhJr/b5Qiahv3X1Bk7PD7xdWt9FpL
fwlfuE/rhUkOervYRJZaeEbZ6FIYIuhSRp8bTRtPQwjH0Z6yd+ySwOh+Xi4cHKud
en/2Uk+bJxNW6oD/1Rze/YoPpJV+7JQucFkf0WsBL9+tuhO1A+5YT3CshpnjTxiZ
YNq9P+3KAp8QAuhMFWCntxgIkCoTdVGNzWye9SRvEQq9sTArVhTlUTZKHuf/0/cg
/Gz5QsyPRsBkIDrIOJOl7G6poBJOd8xRVwmGq2cBfyN6j7Fdu/REnmGiYjQk72rk
pMW39DtVkC7SF1IVNBoxxWlMIwZzziLboP1GUoHsRo5NMZfiJHTM+pv6GuqzjpWK
rDJBgYpLQMapuzxCwCQd/Mutf2+KSjRdvNTHcX1a7q8hr/4VcYRQsGknHEpUKNnq
RWLEcODKsQ76Q/ZTY3YqWqhkU4N939xDJSAFoqqmTVosRC6TEn2/Czd9yikTmhVn
rk1QWUHFQEUHObvo+vBt38mqIou1m++hh1T8x1LBDJraMrPvZ1nSpwe4KCvGzW/O
ajAoFDYBij1yE8cUK6MyWP4wjmPvdwZNhFz2fjty3XsI3oKfo7HDytQuB6PYqtVB
48tb8tfLBF159Zf6lMluts4b0qJ/pnfduHdn+EzR4Q1wJcIT0Uya7bUP3nQj3XEZ
KqwSx8YMXNTHwzDU5Lv4x6o+COhMizAV+4uOlpL3s5TsrYk+4oXrZ5E8Zd/W0xeT
wewJH9Dypd/2Kkc65Ya3N6jCyjDQf8yFgJ447KxBmac3yZ/5kQO5LuDDnaCWfBeA
7oBLXu1Gmsn8RW7IwP6zoxh4e3z6C+ZPe5NfGIE6jqHY9wicvPIV17LxtboHnixr
ee5YIMyeCJgaHqiFYBv5gumLdUKcD1Ig5nzoJdMxqKkoIbAle/4y+/gZlyNcevxs
JKnCWN0zDKibrBlBAEVGJtJR3fZCjfr4lm/hLlS+5sAhpXUjhDYfSoCK/sHyFd45
EYCSPcI4IkOonzB+TqYxdCzCyge9mFcVOrJaMn35xuLDt+xkHkj/RsIErrZxDqa3
ebNFYamnAVWZ8gcsIycvQV+5cczZF3IwDRjRVK2zMhLcznIOwYrPZR+gslRn9aBy
b/rjBfoXEk9UtriE7c+T3wxqTS4KdUI2xEzd7mqGd5Tmnqd+3m08Mnvcthmnsf7g
PzGon5842gQGvOyOb+pz2stJ3xt7JrROv/Mm2vuHBff8fCl3oH8YJ9cJfDYF7FK/
/oNmrDRdRGdUtprIm84YGM9bPfUTYZCrspkOWR+xeiG4b6cxh35kIAHne2Xj9QMp
p2O9xQOq1vv0YXXOibP95Y7rtSyqFjIc4zBL7s6T4Stc0u4glatc6Ar/1lD+I/f3
uhd8C/SP/g3NSnYUJ7NT7Mzid5SrZ5i6iV0pAps9CXVP5FRKCZfVoTMQbKSTRgd2
OGb2Aj52+9nNZGWrmkQnHKWm5tk34KCZyTnNRPnQ92T9gxah51bz9dGAMiX5uqEd
Ern7vqyMIalnS3kPD/X+65kUE7XjU64c8TwqRZJhBFb4xL8uYo9PGggHA2v1g7rK
nNciXOHLaP8RyNjivw/fjm7ndpbIdhVVWodJaaHgOYlaR42poGQJirkqn1tkBO8f
F9So6X88DquqinBm1UCS2fx7SSZEeIXp1i5NWhOyEfuq6gYljtiLJwXxtfuUl1Ej
Y5KGUAU9MkYCvWkq+vbiVzwluQDe+8ZDHHoUsH5UV8VSJv/cIy05ljaer4k9ic4q
NSwpYTepJS/08PbL7vNNqr2qJFGQO8xpxeuqn82u/OqX/sjy1aDdDtJ/5riqSgYG
kx7qnIE0lSpqesse89LlI6KsudzOZFkc2VbIaQFkW3vBbe+O8rhiGYoUY+qjqefU
bSfojS0oVwN7nv1JR6AfwE51+5c04MaDfLoI/rKCuEWbj/vwfPS+JBmS2vtTYtzO
gd9lDEOmzQadwlwPwuw1NN5I+e+UXMkUrZJSWda3wu54eMi2q+3cD8CUIVGmVBMC
KfrqNIbxzqBPpScTCIzO/bhxml43U7DuEvH1SAC6HbNquuXWDBBxRf+kH6KxMSG3
g3qkXQaDxTukqzz9Qs9UD4yBwWH4kOBV6QOIyTSmEhRN39wfTKcpJhYYDRn+iLdI
wRz3GoQ8p1tQ3U+zOfRo9GmxySKY5CNfFB71973RHx8Mf/LFCxLg+47Zsq3/7v30
E5FvcJlojhJe80l+zJvfXPH+oZ57LcpMMEI9l0aBiOM3Gu5myFhNJZNsWRfEFqvp
NcMwT3/3f1ItufwQ5Sfpf0tXMP+tNz8L3Ubw8fMY4bdvcQbckyn1L6bmbEQRKDIo
yUUjbrME9WrXkbTeGi/LRcVUeeOLPRipCDNqwtMQpE2OKgXckOybIiF9vFif8T/P
yExl0167Q7V/ZRFNFGjJ8trEppUHgZDOX11l7DQp3LzDLECZ9HntvnY2nchK+u/I
Uy01mxAMnLY5H9KqWa9mQqadsYUjyTvExpw7gQatY2B64oBSC+XLX/gNjEzFgjoa
wan5qA8O7Fo57EWMKgclGdNZwkUmzbT0CF0Da/xdi1eWSY62oV297h8DVwzkuVWY
tMOktP9AKNVY6NxucLZe+8O/hnhpxldly41V738AnjcG9mUumNxUD4ABZOF9ffPr
eMPs0JTxZejvoUKfBpF0GwktPmfoFhym6rVqyf+WnnAynpfDMbImLLGL1JWReA4a
cmmEx9Mxxab3hfWuoRcjl1xZK1sa8CMsC7O9WCWGH3un91olUXfaG27EhKH46Boc
1enWJyiEd1W7ZmXuyQehRD59kgdL8bn+WmTubpjpoKU1Jza5oM6KLxfptykqI+cO
XqDTJTfJPT8V44X4XWh6sKbqFkoLQDivpK5Y+s8jZG1cdhcgMb9N/hAAQ+t+8GlE
x+g5h9zDbmqRNu920yygp3WGsw9XavMK8gkSS004SHFRpSFTs+eTlz9JW2V0WyUl
M0YDZalUokRo61DLBxXfsmnhCwoZXjAUOe37oiI9z2u8yfGsnz4A5RJo5m5jBGJd
ntHdBNgBLBOekEN8HpYUMNs2VEQDRxnCcLNFasuBa2Il+OZAU8/NUdZcVq335OYL
13nK2dDmkPQp5E7ct/4nSVemQjPmMNBEP69IydGDA4G7ayyMAxs9xv1FaHPS/0Nx
9Kd8UEZs+RsaoOY8EKJyBhFkvnyz+WW4VXGnJ+zXr2S/vEcBA7xyEUwaFsL+lqui
jAwuOKnOnqXPN4UaKgSYPKyRLddxwsuDUrG4HHxpnFk4EyLBuwRo1+yPPsbWYHvN
6xsK0ghritnmVcfXca828ZCF4WwG9qftfdvyLObKLS9WXQxvTGDNk9rh1dLFOLrA
0aIq17OugVCpfAdArheHykeZx6pYHE+7+vek9kYh8nZYjeQo26O7Q0HlN5WwWvRR
6gT7qVrNo1IWrhXBTSuPx7ZzYPHIlM79cZOPxfXWyl0FJLOJzHSTraF1MYGesBGK
iXLXG90E8CEgaS6YjzHAmLhEEAhRV16RhqQz0aeABcFoWESZOR2ogTJ+HlJ8ogQ/
5nJMZFHZ2y8wvMkjc0Q19aR/tCeUqT6S+MXPAqJzaiReC+IoWue3OHX7axYx4JmI
X40wWiaHlKSbSIl68UO7hqpgweGzmV6Gv/WawOIpv91uH4uLjqxH5mZxDcL6Nq1C
9Pdd3VGF5mSb1Picpz89DRbU2ApOiCSZDNfuTFEacvLQG/rOlmPGSbVqaKKNyP22
hVqZhgT7+7i9AtHaIWDcEnyXuL1jmVc0LktKUoHxK6mqZ2UK4TiNO7fiz+3Ni7ck
ToGPRmi9D1Fhvq0nsAP/eWdjCee9A1vcr25a62EnjXuhkmCtmgNlJPZakQ/PbuDT
f2VRmd9UskAwbfHcdoLujX6FqE7lENg5AS93iKASKaT2QsCwNie+O1/Y4a2RzLOm
Zw3aEjulfmIv8rHKr3fxvuVUnCz2WU3aiELB4zvV7nPbmDldIb7SEps77lk9k8ML
Lf8QP71zex6e2ok1tJ1Syn1vrLcAe9BxIutlvFaWSs/AKl/Tu7JDBhbwM46EtJ7j
O4MJr5NwrGlHfNHx0fgGIegR1/zYb90/KTqO3LYbEvQuFr9tKwwq+0v00UdmHgyk
SsCYHdMeYjlRE3osIjGTTMYBwpZXXLQg5uWuZGNKEHQNk9X7yUjREn5IRjNx8v2J
szcLtb1ITwTGEXkG2gWRSrZC6nvOfCGEYxpv3Re2E6lODttKM2fGybrXQ39doMyr
Qx7fLYMYd//wdzjBH+WGR4qaRZLdW8hAjgFi3Pxb6AY19YfxQg5szoATMn0deptE
o1Xf0wqwYDQxrbbn5RII89HqnZkd6x0DQtAWrkTYJqCWeUE7BgZ45qzBJ1oHxrHG
ohX0eIv5YM0M0+I93c0FqmA3YR8A4YxtaiRWR4HKdtcBGpWDm2i9l0420NRhAOJX
Jr9y7a7dMyFJfGRnu+mdfJTRDVHNuZXFOjW5JYTTIJFoxdJEO9OOR0CY0nU0a7rJ
jltI2sy+ezBuItWNzxli/oGqs59WYY+x/+s7Q0nG7C9W3/84xYN1qc1H9qLQx7sC
R7awgJPY6c/t7DJQg4S14m1j9xss7PojICqbv1m69J2bvdj4f0w0VUyR/zE1Yttf
BKAPDq2Sgl9dxgike+fyK5DNxmnJfYDWdBPmS/3jacZ6deUSIWXn+kK8llPUhd03
sey0BdPp/gDTyK0UoM9MgX2eDwI8BTpd2iODsR68msLQ1bBdBbhPe6dgP0+msoxJ
/7UL3yhfWcswZFyuDoamaJ2iIpnvuktRFdtUEylqJZEn2kXjvcC9na3SeT9wLwhH
4D1szVRTFs//m+1pYcuL4258VX8ExgN5+bJIq21HBq8fVHihn7J86BcP/V6BcEL2
P6gHS3hgPYdSai9kgUD6BLMbCuernXV1obNUMcA0DqewSZUShYgY1fApqbvUSY9F
aGvka9HWZn+jO6Jryu8PXwAeg3JH1XsKIaZQVBsZ+O8UoEONXJzGiwCXtY5k5HHf
Bzi1EJgzhHBcUYjP3/hx/6huHlM/Fszm2kzR4+mJkXhqV8xcUX1axT1aJ/lcjJca
7zIoPaBJqVtDWuXaDlJr8Hkrl0KBZr22iZS+jlPOBxsFHAwpNqKelRL95MMTiH/x
MQGVp1rbHB88eoXWVBMrbGVx2XWhrkS9i/6tWG3YrWONTtNKPBeOg4hGdmbjCDtt
rpFt7240USz2mfYfu2AnzkIoVvM0BcssJvXKfMofdqwXX3veu1pNBhpKXXwQnwW7
hqnPOwFR1xtBXlwDZtkmB2Le3qY1hLUmLbLGKXDNQjb+PdgDvsBNVaTGTTgiBQla
emkHijerO3qNmxGiVckHaO5A9swFkhecxYLsGEWLeFLCeK05rZvRregK7m6FAwB5
zFIb+YFPM2X6DEwuQkUFb05eQ7WclKLMD8X8SGIUNbn+hyV1GxLd716duKY/+a4i
9AbBZlm1KM468ruDM23esDbiV5tO7RDiPv++hSD0N15TXlQXQzPPHOA8M2tArtV6
MCW/7OfBi1rYmUQsmxkA6A7iFH48KbtB0z3JPokAQ7vrofoEz//6kOPwOioHyTf0
WKQMJ0H/BCr8++VWZ8de3oAPcSYbR/Mkce1vI4LzVTL6Pk4FYa36yZIgVsSRh+Rv
Bxpw+WRdsG0OnWvTD5Yg3y5RjrXd8iDSJf9/vvbn5ioHBc3o8Ax5HVk17VGNToKX
HhZTBZZ8hTtPbNIePfqEqaNFTm0jcPk+UGocp5lZpCyiybVo2e8hSC+ZOX39zQf1
vSF3ySo5JVEZ0kKnKahVV4dXoMm7rA7k+vqdEllhaiEz9WQGCdp8kj+bqKW3jaNV
ny8maH+BSHSoaOqI/h8GUOEdlIE/WbT994QbDKOJIPeQObu4ElGovXDfXrwPBMm9
k1QhEqrth14EMWz4ZaLGgny9JsqYlTh8bfJMew7SKiBeDxK7307s/QYLFMilfucr
HwLbesD0sPkWJ2TaOyQZXz4hSF7W6CnbwBuD5aIZaJ7dCfuJ/VtsP9LFehdDAIWk
TstD3oQ1VqC/GHWLsPUSaBfmB9X1EHygcBfIuU/kOyUU63LUjvzHD6a0DRIoCZYY
V4jn7/V2xzSHfc2wm21xnNp6887MHtIoJAYPWwzhILryXIqq7VRwFtSmVSJQRyY9
rTk3uwFSOdtbRfrjyYlYyLHlhrKo/lxidhtK/o61pr4xnzGp2AllbYkJ9M73Vv4P
a/9hrisQ78K+e6JH5rPPGwC6fpzBH1laGeFXPUGzMc5lyJlsyIocy8GdBMxcGVDd
Qo1r7pYnOrUcN32WflmEUxmdjeJws7l5JoHyyUWo2avUHgom2306LF/KoKCJT2JP
U1FkcvqxbrzgG0gFuUVZPkc864TnfsbMMF8rQtSmyocNLvKzmDXLG+uBZNF0N341
kJpaOw+zvIoUUNiQfeQnOUbMdRcAPvyJtxFQC3UW+6kaPA5PXp6ko5YdkWXyOplA
800VldatfMDhFO1iC269c8BnHpjJb8AgdvFeC1GfaBEGWzHseszTFdFmo3iGRj0k
jqkL79+vZ3NAy2ToI57+Or431AqNvry1euB+QFJRMz0ckxZL9bS11+9So69kr8Lj
43zCArLnrCq7LgMbFHNeod1c91lasYe1JzL5WjUhLRuWKpUP5GDTGAruqWQvmVgh
OhWdhZlVOBzUn3D08+BeX9c/jx336xa6SZ0DcvaSFUXwM18j8SvPP5RqTJgiYZFc
HwlEdIP/S1jL6H1xLbs22uopgb1TPVRLKPNc5UB3AfB06uAnOQU173FFZOAhA82f
/qEpaH+FlsVx9naloYvm7FmVh6dAiAfxpbN2cIDR+zRjzy4Leuc/+opXRyk9qx5Y
vbuw1rVQTwmOudjh6RZ2ReSdyJFHcq2YawjTHUBFHaUO8vm/xq6cBHY9moiOKvl/
+ayZ5K55VMLn567bAkdD/2EIqgLOlADWAXtD2gpu/muzL44lKk/O/73UK/cC9gzP
6xqk72zbTJUYE7iAHY1jehlVxFZ9XRlh3ou20c+UuVgD4lgAl3V0pqdfhtTdyRCR
FIz4mbRx0mURiI6XKDLqil8xpnKTZZgi34Zulwf7EUtcRrIUxiYVvWK7wxq3Cbse
teiT24/zsSSIzojOC6yz/IWTREIu31tcho0Q5j4SdHgtuzDh9hKd/ZIq68dfAp99
4IvD1W7T8QEUsb2Udi5CU5j/bm1RxTDDEqRy+UcLQUnDErjIWI4zouOL6iMZ61EX
VPIJQsnIuCOFYJSdnw/khC0DQK5hDvEucp+rnfQtzkyAdGboFDaWAWmTtbHpB+ie
MvQyWzxEwo/2OuRT9ut5bkVIQ6BhdsYptAElAEOwb8SxTZlJQ5RL44uFXK0LjzfP
Yfz35wHThXcDBLvA4eYd6zNtjRIBhX3uP1p7D7/oj1bpYj9zSvubJr4c3iiln3Nw
sbI6jexjBK+WNyY18dX5M2vDHiJSSmA3gfJCAlg7WCsUbVV+nhZTA3jxygAzFTCL
SR4AaJ49UYkgPKAiDy70aXM/tEiq1Ddu28WEUidTD0eUOktQrgPHhr5tlXRrke0w
iH5lmrYUed54techyC8X4Ytia7SYmUecEKXtao00adkzA0COMMuIvF8qnOebrhgO
HRuoH2aOYPzihmahwQ/rbPIAUgBYCbXHx1qAvwFTA3E25ipIEI9eKFSUhxPLe8bS
mEjM5D64h83teDdXNYLwgCm9mQXafPVEGhQJ/qu10bcLP1uYAumq8BJCRFS9gnVB
2AzNPrJEAd3AkSnpahvsXMCWuEO5lJITPOsSh4/QKGeKQrpYdRX4fU5/9pv52R/Q
1F20NQwXspy/d8vYaknq6d7BFCQLESextJRKXTaCXlMXUpzB4K1avgSai5xyXGKt
r0ahaShquOXiPEcKKo8U7OSmiZnXT3j4+fO5FCwhDb7YhT48qpajwWauaA1vkdb+
CCLaRXmwU3ODIfEQDu+YFEw1Xg9RbKa9/7EEeB94mGFxGMLnVXQl98xdPH32FFvy
4Ijx9wmiwRgp9SVchrpQFQGi5J5ibG/hLCUZG1xjt5ruz7KomHfnM2oqNCtksXKC
VkuLj+W2ufbNJfmnB4k5z9TITtrpRLY1cbpqrbC/FISGoLfWXlnQmz+UC9JGDHd9
/AuCZ0Ay2LnXsqpJ4c0TGs5jIl1mVLQTvG56SsGzBZb1eF96XWcvC1ln306T7sPJ
Pcu2gG9gRmOAml/ZWivkn1CRNnDq1zMtM16njYkyC+h8e/4URGM4kAG8bHj+u/2Z
foBPg3DbCk44OEVUKDPm+adAN5sLjIBeloRqmKAjSfzKLX65k085pupwNHOWQFjz
vurPCjR08tFR13Ec6V+5Z1TfhUsqI5Ok9j1OCTtWVr9K0/WmtpbmvZOUMrsh0urA
VZ5YRF+ZNFwC9lihjtVhF+jz6De1LMItazjt4+oa5twG0HSeqMYmidUrs2YzI6i/
rnJxTLx8AkFORGB0u8BMkdbcCasuZ5mruuHrp4Q4XEdDkw+kSTPaUpicGYQLo9Jf
BExAw9p+/Ax9gXFlF69r0VNMVPr0Hm0ZWpja4t3vs6Hvc36C+PKY0gIVL87b5SDG
AhNvwsLzodQk1pg3S14UvcCjg6fQh0Tu149iJtcTRlrRBU51hLw5eQ8LXRYlXU/v
8FAmpWPoBpn/p+Oe25ZJ4Pv0K4v686KdQDzgWuo48qCwzY+6NdY3CX4oqEF+DqxW
jniYYFNyLk1BEtXTigyjuDIRX1SjUq9AVUD1RJWU23QcXslJfWKmFY7UjVh6Rwki
bylaH/GxKe2Zar5bQZmldZ46aiteoojqmIc+Bo1UysD8eazoBBei4/3dxlnF04xP
MMYZcNy6l7p+S8gni0XslRrF4owULFNM0o6D7XbLUU0oMQFUZ9t4GbZWPxwu0kpv
ZMGD6RvyCYuJq/Wmb2Eqqcuqebl/PmhA12D07FvODSxajQZRB2PCTKKjXr+e0o0y
w1XECZi2cl0vFRi5gSvSI2/QIspkvgUlbNP9znv/LUglfbowjtsdY+nD8VOAEa9i
jyeioawOH///HW3Xa4CllxNmO7Lp3CwNCWcxyeZeBwLe017tuZbW/KpoXVahj1Ww
fTuNxQ9hbZAEpdXLxQP1IeRxTOgDtiON+sQ55AHaRpjFyoL/7qKUwORT0fQZ49QQ
mUEHPwwwiSw2dvdiEPGTIfS9LB5v37teBSYaLxxKTy7OTSK99hFxqsGaSR7Ut2IV
K5qcSrUhQ7yQyinUiatelZu3CB4T2MrD/BAZr5/7bQk0YBiuZT1SEjEDxFBDtRwe
aoMipgLS0gMyVhzrZxuOZprZjl3hF+Jwu1seTnS0CuJet4NsnG5dP+y3EjL4T0QV
UjP+UTTcIUMrY8Qo3EkI+/Nd0FDyfG7J6P5IH2Z17ZiA4/6RSniuMbWqrSsU3cFg
dMav110aESt0fVNEUbbuDJp3CIjUHsWScYqPtYPjKxAt0/HDGiEUtKeE/Ru55pBd
bNRkP1TQmYDqQ0HpY3M+PxeMvZuUjDmU5s33f+PuJ5gtL+TU/h6vFGC/Oj0wtJVf
X/a+NingRlVa+mNmczwI4hekV8iCFG8XL05+agJrinGlnvOa0yaZvIbROYtce+Gu
eZsnbAex7Ij8VbYPp8g6tciaweKKGVIm59C5EXazyRbmFt2NV5GP+s1JLdmVMvo/
X8pYUUcC1Oi3KWpGBbtnTZdayYjuMmKwvDCK4kG/uxC5VpwerALZDdTyCgxIvg1i
mxEir/HfrY2LqgpF6/vxWECImOQQf3dqLtm9ZEp1DnwtKVX86M2AKAkj694b+zuC
lu13u1s//O3vPkUZ2ewni8qBB1zIf8qcKygFjQifHmntX6GP3iJG3pbN6Fvu7CAD
oNBnKvla9/+kqACaz92L9hIh4uwdTJV5gGU8RYc/DCDKeRtC11CixPnC/eG9CJXH
/xkpi7BcOVJFf9ysDPSOHpNMc1+TOPpRmyn2xNMb0KN41NHMSX6uXtO0oaNvVLF7
Eea7xH+qLyd88mbNPU0rxZVDgy0fWQKdheozWv8tYxRk4N76gj/A2q8EPBVHVXMD
FqSkmD1Wy9nKs2jn8UA947SRP4XdwjkuOq7TJqTGLE8MDJza4GmjH4BfrudcQEKe
HIcDBygu4lDjbc0RKqvs7O5xNC+GcdVquOJNXCvoBDvBWK/Ze0Ihu68r+4Hloeuc
sEvM+YjZZpfspRkVENQRdQTnzEZgB6cTg4R+QCPHUSy8rZX6bhXMdSinThAXppXH
7bsook96+U/K+N9sDomDogbLic9JSYSa0ZSdgdEw9bq9u6/qJLduKuKmQy/JO28c
+CRBcgVLZc/C8K6fJGcN5ZKxhvS2UqFSGLlSxU5/+banXrsytLPsYDwaRLLOw25l
oG9DGkt35EXnjWyxpoVeXTHzUjU7iQ8OSJZ9GeHdIRUadSnER+Cg9c2Lig3O2Uxj
LCd1vFXdYSdCyfWbFUnYtgOo9wREeMZ0XsGttiUgVHRiRkOu5FWNtIJpZtxXqgP1
K5tnlGeN3J/1K7iomLnnfv6FUo+GkIq0GmJR7O3kuMgnrSkpD7gykvIZL6C3bUrn
EG1QDcIjuoF2SytFUhZCKQOkey+7qoUhEWl460OYHLIiMqv0yK+r+61jdXgT1XSV
Xxai7f015LRre0wMcJKEw/ZV9A+ziBV0giuqO5c6RhrjJTssCbr4ohSeXIc3M5FZ
+WL9DitF0KlKs3n35JbR7fAiD+46S6BC5DZY9e/QlqkQp2Y/n2bD5Nkodwi9BXwo
u7w0MIJmYCfITY5rBhlkJWm7Cc/ZS/fMfx8WIwNqkLQ0iwcCQDOdeHOrQjDwMyuE
Wihgs/KskuLJYxVFAHbUOJzBUMmZnpuMcYMXWR5IzEUlLCI2Z1MCf1uACefp+cKD
WilV0vf08fBiqNHBI9N6iEa5E79CUNmde3xWmJC3R5qwTkUBlDpay0wjqGM0Ody1
JpagBtT/YT8vlJWJojWqlsG8pM3lnfgoeeidWZm6KzY7bMRwICXZ2g04/EnAqnt1
4IVTIvnXapC7da1GY5Qwt8JJZGU0OpsF8o2E3ymS56QtjRXKIa38FjkPSmphiWSe
kVfc6LFIfyohIQEKag8sQaa8fjFjQkFYR6eXSDy3nBbalKQU3MPdvkqwqhpxcw2t
ErizSN2Z+Kd7jVpKOK49uaRhA3uvQ2S8F7f5AxqLoyAyxHx3f2btKq8U0vpfrc96
Ds75ze2By0LZuxTdYbRnt0TmTyu387RlfF8yBhMtOots3fQ5Sl/ruLK3gSDroNdI
yp+2Xve2n9OhCpNKhNtF5o5FNGzNKcN/Y5R736KHRmahqktF/uU/OWWhmoCdt6fj
43F7KmwIebd+Tqo4Gj/80er/aUaaHu7PIrjressQnagMTHdVo9T7nMqBArfJeEqZ
/zVY8ZmyRu9iCYf131sdYZ6cu7L2rMt3eANvMUsfaeL6ntMVHogrX94I53tvonWN
dpKlSDYhdu/G1I1Vm9wJdlh0IE7Pqqa8xHpoUiGIk7jcIpSCp2Za8mleOmOcAWnK
yjnnXh+x5e4c1gyVMxyL7EYCQbQ9k36y+oasToJzlbos+UJl7O/D0iK3K3m7HXLq
/TMBqIODYf8nFuT46Obr87nWw28TiDXTS4NSBO6BgtwJ+QKVIYSSPlw5SE2aS/jY
Qfu2OGUQcwndoQQbJdnZyUOIh5SfiwyKQkeOwybJ2o4y66ky1PSCIB3GffyZnml6
Um0GYxOk1QSfYG0aX1SWck1ZQwYXdPe1cZ83Njcumex2hzNAT06873U/2nutLxMj
KYVjjlJJpbLMTZg/jm7SGZ0TzZ441F66rkK9pxDexADYmyAB/VB272KoMcBPTh9P
CCduvacPadGxIaHZAv4XXB1O4o9KhKR0yMzdz8RM3eY6Qt6wOoQk+w3rfJtm7PnL
HOi6SM1nMNCPjYdKboPhxNZXkDtEfC4YRmz+KFICkDMHD9S1n4lxBP/VEKuJ9JTZ
J9EfjSJ9OO/QbRnYYGfbtzgr1HhoTsvdGxCRYeJ2vB4TttO88x3oLnyj7SR0nF7h
PNcCMIRtiZq+kTCJivkPaErI+cBS2gIP/xJfKNYM3Sdbuak9Kw3USecMSUoOy3uU
cJxX+yl6BHZIBh3EZbTlLGxvSNNk2WKVAT3TjWYf/ooqpZuj4EVci+Dh2KRXXkpf
49zV/sgHjLVvR8rP68rgB27u5h6ii3nvio7Hr/wam01o091oBtA3RMouUXfGMDLY
HxYe4tmfl/JclIIkerp9Ib/s3Yvhx6hBki5sBRWY9a/aH/aYOqbRznBcdwh0U2RO
h0yYh/w0lHIAjqx0iacClr9URNE+VlNfbwILv4Oq5S7JxnpPl/INNsAu9onQnzGo
DoZxZVsjUL+FZI3S0SUwQcvreLEjoF25HpAIYvRlnGfNMZPkGApchVRSeU48W3AA
shSriwk6Gon1rWGKrY7mmAM272kcNhLo9RJo2jGs8BhnQep/PM+U7x0ASnoryUG/
2b6CHENPmbiq9qY1VydY/NDKCFvG/PtfQIfYdQH2wFv8dGiR0HdTbrGIIQb0HiOs
4ClXuD2tYqEQcTtMg86PgZY1BYHeHxJRMaiNOP36Rcuchmj9IObA3QZB3Cl57BWV
HI9byWPa4l4hseFSVcwLCp6DuckIX/Djl27EzvDuyqeOXTSvx8pndHOlawIrNA2d
/FRpZX8LNKWQQprA84XvE5coQG9yi7V3NKcO1na0xc3SSA3rer75EfkY5zu56bWt
QFK5xPSK0jwR/AN6WpLuUB6iNtZytv5LK+XT+Dhogd79eh4CZl7yac9cFsa4x1K3
pTSasMpt9h5RtsHSiwRLsWTSXHkwtaQA4k9Vy23mXuWiZE5G+7c1AdJW0W7DkFOU
XdJZPOQ765o3jgoh2d7cB76jxwn70y0pQYrcKNCY7EVHz+seH3Lirs38VDzZhw98
l4hDZ7r6N+EK2UhnUI4L6Amk6KNR5YibQDgOeWSibVKqY1qaGe2vTToZlqVYtqHG
MF+QuOPdNYDYeUq3flcQKOTue+vQMKvMjfmDU19D97shGfXXYRamMmOY6kLXs/ge
gHthoe0VSJMLq4iO+aG4F/9YIYCrgIK++3TBmagJEI0uVI3NE1ZAMy9HYBBsX/iX
1JyByPfSA3nt7ra5tdddvYih1tvWYwfgXMI0lDLnjwpX02mAKJ4xNv2bvjrnSfMh
Lxp5eRH62LnAyzfWm8Gbv8WD/TuYRznVDYdT8y/nccZDDlWKWZemJCSr0cTh4q21
TXQpP7X4C9cupA7Kmj3lrNgBnzClcs6XE37jBokl6SYOkK1Qsl0NiC1E8R3y9uYb
G1EVr8IveXNP5wGD3Rt9l3FhkbMZYUNPHEf795717dGMw+F/3iGxrynPRHgwh4nn
m+Ibv9mrSSqwoEr8oSjdmWsdm8XMGUirCJvtbYNMuKfo4o6WA4hb6BrZH4aT5Z1X
3ekCECaceMhnuGJVW527kROUR3zyY6/PoEWjDVP+dmSsB4J+PgicBrkLFvxLYYS/
sVs7DDPJ6iCieIQZHLxeRCkENCgHqc27nbwWtbg41oej4RxSvIXheFauoynxNX+6
/nOMFs6cdG8AUQVbgLUvhSPPGuoNfCA5CjZUn6R5LILoBpLfIB94e5kdfhyit9kg
hQ21sfmy4yfMMNfXzT2987uhNQZQjjIg7u5Kz6HCDG4aZV6y/7Kvr7SBcn5kxmeX
A/YRbHq+5iFLRvSBtom752YCanRJNJ/ETbInDAffbVEuqM1Nx/IsIFkJGFp1yvK2
t5WpdmWdejnSty68owKEujjkqqJknOBf4afOlWirPmhXv4KDtfJoLlZQtE3wx35p
lEBAJ5rG70lmZTd+xniMSZxiES7eNAKcL7lMue/VKrFtc+BeZz+P5TzWPW0rnWFe
ojEW1Aq5MiHMfuzWkgdSW2iS550PHnc5eujQeH0xgF8tjd5kzsOlz0YXD4BfSFuZ
7DrNS2bXHIoySVYYDTo9pTnTmfhsJFYjH8tZXTQsHHP2mQZYHRxP+igG1tTV5LuN
U43PR8PDVEzjzPVZL1FUSyRF8JQDjX7k9NcvcBo3u9OY60xxtmwLtrCPMdA1jJVB
jzPZnvsDXwOIAfzHXkWlxZoDL2cmV2t1tjG3W+HWOCGZ02wm3MFUuvLdNQmmfvqx
ApwRavOfEckBOXwaT1qF29j2PpLBt410Z/a5kdc+iuHuONfoAsvQ+/Iyhv5LY8gC
yU9PKHn35m55jZNExWzWfY0CyUWB1CAKFiC42l7RGJ4OH2RXHlcDNyJylWTbbWJn
rG6FVhA2kJfRohIzZpENl2RGNzpM2hCxa86+CzGq+NF9/cGpYfYv1jzDTGt63Rsr
SIswISIY3G7nJ538G5tdiX3WMl3QlSvDBFh8Afwgu4Rrwv/yP4ivntbE0H5A5fPB
ylR0eEptlgEc5QWHqfdV5uYXrb81dXovUOz/yZdATBEUT4Lz4PhBF6rNIxMUFSz+
mq/3MjUAw8hEn2sPhY04TeT06I9z0cRlzNW0WVLYO91Pt0plhDCcYU7ubsJJfIvO
xVU02yJcFXyN5PwlpvMq4B2/+dvWxD6YGWxZUeGjC9M6uNRjpTW2OIK0bDjbUJDo
1OB8fONd/RaivRrikPBBuiJ5aLnpXq6FgQPba3cPzNZ3AT0yTrF3JvDx9f3agv4p
Xh/dpM1ABQjoiCi9uCGrVa0/qUCZVPe6CvVJruGRboa+rOyhMwOd4AlU9vnt3tKK
kevmFWI9zowCmrGYh7ddOs7SxRpPJLT/UGur6vtNImTrZI8WwZRFCAt+I/CDl5b3
h9Lzc7yGmqRO09Gcoz9pt5o7n0fRFXd2RCBH0zK9Slo8muRDYmC0S/VtSGwTeK2Q
oUs0ixhksOHrQV5AI87/rdyLE3SnYheBdKADXfzN/QaCHxK652IqHEfA3FaRUNEM
sTGxh6VEtHRUV6wgeeQI92kBqSb6B/cFQVPs+SBMgYPyWPJGb/B0HfpJTMLpeeYH
StwlFo5TjsO1WAWq+CSOJfgGvsmmv7xsuldFWzJNNkRQQ9kJrhdL0ob/rWhZgQxP
bfrY3GGsapv1mCptFJIf7601SP9dfc1vSK/Gfi5quEuSg2KN4Lgoo1xBD7wUQHNv
3/KErbrKtH/PlRlVDv15gTwxe+otgNw3By69eKfGnYO/LPoZIFU+jAKokMh0VTr1
195BY3iV7l0hGVlGRpIANP9fMCZIGFNn3/JYou09L0G4wWP5yTYdr1KBCWi+tvsF
EQjN7nvGYN/ujI93T6/PMjB3E4WiJzaabZRQopipOIiprnFi/ByYnfkiHmWHW9/y
hLWJd8PLmwOSBsjpcNcJ287Lzmz0nwnO8RD6PxjRTSdVS5K3jaVm8ehtgMy+ajYE
2c6P1zylKYmWoQuTBH/1WphDK/lvjfYJO0A+pJW9g7dKBFCDWJiaJqEdsnRIghoi
VtIv4Jggx12Vtg6gkm1HD0dmPMNl2Em6y9m/8z5YkgZQdnB3ya5swwsQ1TAovVXu
qlB2emS6zbl/5o6msrAetLIeI9kAi8uGCp+hB6RlZPQDWFqOGz//ViIgMb/olpMs
S6mLpEcXCutARjTR55pAsbcEkZQgoPGzHtHY08+JjvC1cZQpOuoqC7317ZtNWnnY
82/y5uHsarnOkOvtXl6B5e2qfI8aZ3VunTxXh8PgQ4avxLHZDM8Q6beJmK73GTcL
+KRbs/YhF+KodfJGE7HvKUzymyFwgIZDvSGIuGszBdWOBhZNXzHvLHJs9YLTdYbi
5KZK6xy/PjM9LYo0wSLti6PixG8ZDD9s51yMA9DrAG1sGGm3gTdkXAKH5dpxGups
oxtJcGLNHd4SadCf+feTJm+oJzuLuxRy+vOgjtFMY9C+SvIGYqHx96J/nEfbg7A/
3Ip7P2ODkDA8y/A6Tj0i9LVPXWlznDeLRCkvAenLhapGKOwDJdPcy0QKGOqiL/xB
lJyZ1D6NVPRUfrTNodG7QubiehnR8XXGt9HN4csOVBQHSv+hm5WWOhtp/GHmAnb6
3E4Pyrn3s16ohxaR/Ia8cefhEYY/5Yy6zBA8QN4M4QGVtuEzddfc8gVRS/7RR3yD
H7kNZtjS0yF+C8mEQNG1fpGwBJwAqDrXeEizq9rH9xt6BWZ+3xbKRxTHpMoNHUK0
mVxlXQJhRF6ccIaG4TgPtMko6mmx7D4BulQU3vFEPQS2dGarxdht/+45xeQGV15h
H69TQhMEZfI5u9JXkyN4p3RWt2Vbo9s7xf+Q7276o8f3IR0yg+XFdd3wX+D6CtLO
hEJUEswVe9TL+BPwpNZ6OYd0NEeziN++AHBa6e0N/ea4ryxLrBoJAue+nnYr+29F
Ahc0xIoQIc5qz0J6wrHt+qXLwScluwWH3tajhLuVNt9vdhJNVWyjg37BgYScL2J6
QuOFeUKuIUzSqA0lnxsx2DrkGtXJt9AU9hzQ7CnM7DD1WsC53sAMPH16sGewza4O
JJTUhVpPN75KZGRwHbhXR7+o2OArptTFZRxAOXiRSCngNn0CZObvlvMfjzZkpNX/
hej6UjyeRjJAMJRMp2uX8EOaM90JzZRuHVLQlX03sy0Z/4m2x2hooDnBwB0QSSmS
KdlpC5C8vBPvqm17BTwllSArFFMuQMs6fF/5QCv/taEG06xYEfTX5AVq2HqNwWEi
8eSZ5VmieBhWT+ujWXDDJdhMwo5TZAEILcHPtMmXVHxJE1kznWWc2rUFAnSREBXc
97oEjgIjmYH4lIky7hkr/EjD2lKGVqLKoG7tEVaFj/ZRcAa81wpJGzABuSz0jemp
gNe7ShjhFoxEsMA8MwR/TJ1lB1FJT/5YOWSlXpelzRtmuZoPlv30UwdcU+OHO9dO
DBy46IemRZ0QY9WuMphHeqhwwzPsH/fdaaVL9FQ+yvFhJw1q6WmuWzlU7IV6taNq
FSBVmtaFexcWeFVABAYFFpEYhwUi00IOYLJom447PHfQtSx/HgYCLvCWKJdUWup9
WFsXu8DF1yfJOBx2xz0fmtw858rYH1i06wogsKTgT9lBpi5yT96y50lCQH+ma0oo
HzlMhgMsJ4lJJcODsDbLYbYWZ7afjVKxMa0y0vCCSSq1kZHiKmGRgWdzYC93Pb/4
mmgx0E1zBCqe9pzVF2qeFYh3nERkjNy1RS/Qw4xmlzcjJ9lffdXXAIE5ezIAD67E
kCZ4HPAKh8BS5roSE8JTBWDRL2h2kVKiV2sAntUGAVYlnNx08RbztFV9eWUJdSGI
IKFe+zHqSwZnUH0RbVcHoFpoZm3VHxrYaSz01kN1oEvzF3TeyMWXeQEqc0L11ENn
0nVGAn2Z04tPp20siKJiFOkx0ejed6PQ8xQFxMtKzU4Qptb5MA5gDdGZCVwx7x0g
QrZQ+fcnYDy8jDxlJRga6E57OHePbSoP64H1Dy1sk/3sUBobk+WArfa+ww0mkr6f
UHbUWCReoTZqtl0pkd8QY2F+xgJNxSwqCLk/Mz+5PzOk/6wQhB2UwBVdtZR1ye0L
RTBb3ttLVTORljLROM4RZTMo5ISMgOeP8oOEnkgFqjPlQKgZ7BhD3NvWlueuc2jS
DJRf9zliDts9UPzNv61w/vRM4poWKUdEvYAs0fraBEJZ5D2SV7D2GonRd2XiT8Lj
MAC4L3Ik6EtCRnsTtcpuQQZkQChIu9+gC4t7dYIQqGgpRV3/ci8FQg8tTxcqPm23
mtwazsvHwe7ypqccyQ/U0WJzTjcbiHB+g1LmTYfdDtb9amu3Sn+73G8cAFVPS0f2
DMLbKFQTYvQpoBu/D7z05TR9ZhsR9AVXD1SKrFsU5E0fr/vhhDXJ4IWv4RBeaLAG
aGT7AaxKbf+0Z1B7WbTNl5U6DspY4tV8AN7MmFeYpJ22vl/KlloueZYonn1zzXv9
yUTBA0/Ct7h385pc0kIU7DtpyWLqDR2+md/lwo7Hi/hN6qX3/nAnbmMltRom5Ao3
gTGbVDCTx7Na6c/09wIRXWGd3ogsf0MbQ3EC0lY7uhSqjkrrHk3EyjD2OR8oRANl
gKrgKff8a14MxZZjDitaSyGVD72F9znhuvda6LF7TvZS5H/rXscwUdUeOI0cOJeZ
1k41quuibdHDpRp6bretatFlxmezXi4UdED3/riLPxab09jbdtwfxeDIRm9SEl1h
PDnVAe4maFjy9Vd/PdP5OjLQKRUxg2ktCK2T8uALVfaZk7vhzwpLYyrsjYfh+5iT
rAr0hNzeCYhaISltSztqkUKj7DACvfMM3KM0tTLg6cE6pgq9wpJEvjIUkrpuE8ie
1vi0vuo522y34ZzhXito/cIDMwzV6RxNoOQNT4DAAWkpC5OkmeP1m8s0DzI+E89w
N+BEnvkWrFCks/DFHqpuT1fqA2DomQ0dgqVDeB52VKmGptYwuevnB2m7PUKv6lGL
YBCvECHnn2BJ3B4yR/nSoKS8uGUn95C4nLjDM6tFDte1R3r5uAntkpwgL/mtWmFl
oNgi5txEgV0O3LsldEnbL7Y1UlqwiPO5AkW9h2P2x1qxyu0nEeJ8w9mSAniUD/w6
qVTP7LfKXUr44ygF35xOUZG1vvS+t6UrgwLI6P4HGjts7NtQjLGZFqgwp3sZpNNv
4Hjmtahz8tHC9rm8WS1eKgsZPKCT9pQXj8nCirGpHvhmY1FpA8ZsgqsU7XAkiTVB
xL7ZTVXQWVNtfRdFCtgD8yVT5DrcOl1q6dUcVKrE7AHpmY/zWw3lr9mPDEju7Zzi
0sst1OM4kH0njnz2JOBb6/qicwkOZJqm3PvZ5EgL6yXlLUoL0XQhjgmxPRxH5HCv
4pvJUrlB0RREQ4Qy2oZjRoAmzV4IDOqog0W0lgrAvO/yJ552Eva0dn45qhtGNpxj
x8tmyqYr0MCN7/SDtunWS8PCr8CLkFlkqxEmR2FQbSfA/pf8sTh9xeuw2b1zAgSY
VdqaWPp3HHd+L94R2VHnkGme0MefSs58n8wPduucs7ITgRGrIfo5c2KyBhq4qYJ6
CEvbhB1Yvn4wzC2wTA29MQBj6VHANiQnKloni8bC8PDxvnuKNtenjICg9Hd+hCjp
UEHl8PaUQKWOfMvos+2WDRN8FJt+iiWPUr9959ALDjzt2Tkd7CbuiIo2NpCSs4iz
HdfUXlmNUrpUcf54EJr4F9YIhJdLSqwo2U7iTophcBJrilLaeb06qi6ue2rEhn+5
78Tws8p7q+zAaA18l5KsNkyw5+kwqXzyiFMN7c7WhOMUSy1+k1Xertp9zUr90rhW
SpWcU5gmN7o0ytNCk5a0VDb6QUAnlTTSdgj/7bpQCHkY9b7uyYm2xpmIso/WIJd4
MkjF06//n11ncWIYCs5qbOLGB285hPUPpZ16D/l+utSokKQxm6PRPXj0mTknBMHP
wuCFbExY090Kq8KBePrXETMWIMPEUWlAAe9fK47ARLUbppN3rSzBG1kQgnjT23U2
vYb146B7utag3/N0GQjzJ5y36LQe8mCAst0QeuPY8D5LyH606fp2z7Naf7SBI7st
a7fEexhIXt5vErSoVX++L45VINrRJFcHCu/iM+mqLXoV+ZY+On+Z/PPeu/YUiUbL
z7pYEQOLhXUd0kQpDpQKT4wuUTVX4AlFJEmqlD1IcYpY0fW4vOqfHp7Wbr+Q0CLK
OuSKo6Q3eRRYCnvvCs+gdyLYe3mNQQR4P3LRT1Wd3gSsZnNh4CMoeOyL+EGXh3Ak
viJOZXWmM99tXw4RrO14wQAzkBYrD36vLIOVJuhZep69PAICcyPt21fh2zcMOUkT
1+slKQw4xxmoAGr5p6FbACKn8nf6DqLOT/V0pBjFKQHnfa7VRM0SxcXFzGUdujv8
VtCwlVDBJyv1PNycWhqSH/bZ0DE+aYA78QdFdf5CKndg7sAcKAisp3bOrFb7q7lj
0q7fo6qVpk0XDAKY2x3SUSEYY6xThELJvb2uUnbdL5PsTZAMGTnpV4TvG2ASqohe
ATCy1pZ/JwPRitaQ9TfMDjMrdwZeUbZzlGAPiDnn6DT54mWPO/aJIqgeHuTHUpb2
/tyKo/3Dqqi59/z4UQIM2QEbsC+mdQKM4dIYyaHziOUmJEI9WdywJ0nu118lDlnW
AVYjjATxSpGr9xWXCQSPe9kDtntAYCQm8CiTMbij/+H+O0ejscdNjawzyrQRTMWW
FMuL8QQQYL6YB0xe+Pqm5lBcE8edsPFNQZ6Kpzet5qonWGf2CbILMqqaZCuGwAnZ
i1kNlpCFAhMjd4lHuaz3o/WhsRfXonIx5qUEb4kZeNl4Kz5hgfVfIJ9PrSrJ7+Tw
hzZdv1e6JoCsDwPNthSbywUi5Jn5C406BKSULh7Lz0c4Avm4/B9MQYhTq6nBwYc7
NphXznJlB2MyskPj3bx2u+hfU6o5JT1vHrOMpXT5k9ikMhJaGwCveJ0jDRs70HH2
ZHwo3rSWjzPzXrL5K/CwyQvypxmIdcuOd/0djMA+IKrN0QiWscY0yG88qbZw9oFc
wNdt3rWQ9WtG8UN5WeOLDwYx/S129KAtapG3RA5N9g9Nq4/soAeUgNF48rBX+q8K
EirRD6fl06WQnNfiT6bRxgQAHkttu1HhnOD+2rFl0OVK6V7rblTB8LML0g68j9HZ
haqS0WaiAPQz1Keaor3AV39PQf8ZLrHw6xpA2yrczO42BT9w8tn/5duX+vZSp6Ho
3Iykc1Q2r0kIj+ukOnFoA0uEbQghL5iTmmeDfaFUKZYFV6ZG7WTBxToPVHLDm0gO
/4uqNaBSMAvPxq5BMdhRnSK7XzhLaYYWxIAqFpUOToWDW+EnUKCnd4N7cBD+uOWy
TqFXlOgqJgWYIYo+3j+vSYAo3k2efPBmfhJRa9ZUN5XdQkSrW62RxDQHZKGMo35O
q4Rgw7ro3TKQFwbx3hqQCWLqbzTIz433LNtDP+LdNjjMMKHgBbSR1umQozfybHDy
XutqORMA7fgT4PbcIdUHeD8MMYSN1j4/4UjaVOjlPJmB4kyTXHBRIG5G91Vduo/z
3+eORdcwgN8tjnTa2beMDspJR16znASMAE7eSfkCvf/nPEN+/6QXVSu6lzQGxzn+
9H80JYQ7uLiCEWmkS+P5EVSb6OckMDpbxmCm3jM2O1ea8vWmzDw+6tqbD4S+b8s8
WhKJFgqwEOvyCbRHUcS/OLP78nMavqOFGt/66GUnyFtiwSZplOmXF/rptDHcqui5
zhOPIjfwNwvRLQIGyy+a32pB3QhD6ytiZ+v9SStLL6ZIlijeP+qafS5LRIHyIno4
/2gZ4kltdPdUwmi/paYeyjTPzmvSluq2swf1bx5HdntHdhpu17tLWkUpEsEJR/P5
jJ4nO1Ss4O12N61JrrT9OC0Ty8LCjzp1bMsEmwTE875/zqstCThIF0M8c6iSXZs/
oOYGiJ4cUBaE3tnAbHihjNq8oZ4DE24Fei4BnvUd2IJ/tytfTiy6CqbAVHKqpltb
kKhZ2cXj0oN3/3+Yzfg8gqx7BA1x4xT97gKm60MkR6oRrxjrIC0UwzyOTtMOAf5w
brnSUUusHJ/wvHjHTYd6MgxQRTq6FbSUywY2jSRz8499B0Yh0xuHQpRxyHzLsMpW
ArnOk76ojPCkIlml1ohwQo7dRtcf26HZSkqQjPrAgaHq4xFF3Tbh7ssJu2xTBfjj
M+IyZAYgBS3rXiOku4xUeE8v5eOs860J1UMix0gBog4tJQELDBH7C8rJ7BsM4nhk
VMWnjRtgia5shBE+Ky0v2x+Rgg1eF7E9arcFEhnfjkdXaXLzg5wQJGoE6xWB7/hT
UY973oXCMRDzODU7Bod07tuuk8IiSblIqtJeDyLBNU8Ro2X+GwEt/gENBLM4NOcR
Zh5e/Lp3d+XQ5FowkkNWQP7ILPuOBpScViCBH/U+S/5Uuc15Oh8ihX0BaEBpkLEW
sLJ26pVVOgc2gKpI85ublWxMrz0oQTaiPt2khT66yZsKskkeCBcnGmEjDh6HfV0n
gtwjT6j3kdnzrTwAEuav69LGTqvyTIrE21Y1uEXZgiGdHqulFdIF0Q9PAqJIZFgD
PFc2iDEhFWCD65d++MEWPKK4FP8PvO6aC/V6IIH4jZFF1bAyMdTBggl0rggz7VAc
NnuKLRWYc4YNFqX/I5gLRGKkRDXLbXgW7tCIVv4+jQ3s+/R0NLmQmhOV/Lx6iHIC
vspGENmbtJeyCS7RshTiPmUjrZ8joN4X3p9Q6HMP2F69jthgrHa6dOaM+tLJJd1u
KfeKLo4gaHCGYZLnZBNLxuOUP56haQUaOzYKsl0lyEcgwqnG0R7EAiZ/Gkelypv9
VKX/6Uwg7FiRe5zaGsJUVaRWXgqus2xGHhC8oZsrwK5+yrEOIOkxm2cu1yNKkTXb
kydV/AZyTBjTVKaAcmUHArjy0EpmNIZIeiVe2KEqLAa9vnNOcbc9U75fe/hFHEgA
3PIXlkv4up6bmh0/Jsyg/kI9rlJhfUECjJAB455JT1PJnotleuhO4rIkFhiz80a5
ZuNkRwDcCjW3uuhWfJFULifhbViolFbQ90Cef/8fpgd5sHNsy5d9W1WnzVuO08/7
Wti5tNey0mQtDJ0Na/HF/IRKUg2u2LeLYDMOtxEiUAP8wR6kSUk8aDzdqBpN4FYC
SBJDmBMe4n4n7rLHjw7saxCQGEUKjPVfTM7xtVsZpuB7v0vYtLfOx1xKzcPSPXtg
9pU4qRjxolckJlTnB1wb+4XOVwprc5Htye9qm5pkcu75qNcHEqBrDf26bxTTEEzU
fti/YeHaP55+LaVKQjqq5UwRt5uApuvxETFqaYdV4x2mRTvY/aaWa1CCo4g6/6ud
TMiYeYlrVvCfC7s8Iay5WgBcrXvFY/iplXgAeH2uvpXer4CTSWC/Atm1aSjShbKV
Y/s8wBoyxBK+64sVF/ppMZLCyemDedxDCrWOaa+U/P03zy+isqp2yQfjC+btcJQS
oUJ9lq6WbbTVvzMUloBE8wb1vDphXx2G/zhRS3BEVyap90DKacKQocDuiJPNHDbr
te5mNJtZby8e53NsAnwEKETw7Gd/DD8IdnSP5MlrT3fZVHVkSM1/GfrDur8owQ4f
iaqScAB13Xacese3fen6kW1NWKOkGyLWkvyNPw6NDdwIoIa8m5DIcJr1ZcRayjBW
Z2lQb9RpwKiAalqTZzYi11JiSTdpu3FgORmnvHsKXS9E6YTNjYT+I96UwYzhbYQG
Q+Y92o6ixw8cWj1dNm0zCCVWh9vZ+6lSpNgjxCaMRu2AZmCZPGJRv4A0STRybKEO
X26gnF2tUhqQmkODCnq5he/2C+gmVffJ5lMWmBru4QR6VE43e0hnAdWQZsN9/HXf
6S7lt88d2U2gPQwXcPWGtki14kuzqbEqDidShgbpTkMGIyD4o0bpGqMak2UtUKRS
f/JZ6e6l4PRHHXbqvB6khS1DhQ/JlVHTWd3JkL7BQWTBcUP8AnOHfdPU7KP6NCEq
k5ACLLjbko2lOZMDFqr5WuB6hYTjhdiG60zRU1H0osHdjrtIqAkjysTmilpLTfRR
oLvov3zsQ7YyvG5eV6Fmzixl/9OuJz9TNg126mSfGoHNHcZijMYcfB+CBBO9zn0o
AHFWO9nRd6F6vh76E9NdLYGMyrR/QTGe24cbMN1uIuLIs6hPSRK5f6Koi+VDvU/7
WeftIGKDJACQm3FGpx7U29oJ8KIZjSmPsG26QTvKwS7mEGJcFzjJhsy2YeFaMgYd
+Je7viNBmKcaj7DsS6Zxqes4Yx418WihAdhdnxNL1PhzKLIvD85zM3bp9iI+LYTG
1Z5CgXdW7kZ/YWJk3S9hidze7CDloYcoVVeVZygxdbzEUNTwvoXQ/nGiFQzR1YLZ
dycBuFsjCfnfKIDRYztgIa59mOam+JgmcYGt2rAKDPRrUvUpbsIBbFqhzd++Bh+B
BY6A0IFnNOVsl7gRukaG0IR9tUWEm3vVOlB/413EyUsuD3jRlhZpkIHW7AoI2lqb
x9RLN9MWUr0aQECYp0VupI4opXb2lZHqtRdHjMT86UhVzK3pgNn1mnXDvXQa4GpY
z7Yt0BY0162zPg5iOidcYVXk7xKpXpJUUjDWiAjXfAQV6Cp0qAxaXdYy5Kb2RJ7s
/dkQFvv6B/L+na9fItjQqOG6ztBuD0FFqnaqf/4qyxuVAfw+WSzowr8mxFfqp7vG
W3OrGQZthlwrbV9QDFdiPiFTztCEm7zTl0SQwa/Waaj0yz33P6y9bnWocmejeFfu
uybMFgOik3U9ZPWTHacgjM5I0A1cRE37M9wTCyhnBYPE+gnZTWfg+fOJO+cpedIc
cCHH41HPoGCbwc/2KP//b2D6g940j5cisFTremf2MCnDHcxwOxfE6Xl63DYiEED9
8TBVPa2EByq8CoM4jc8VjPGXr+1OFaDyhXOxcoisBDL81rjnZnvqHx3oqUj4T9o5
DgIuYi/CGByYm259+32urTKszy2bJbqhg1hm28h2tC2aezL/YeymvSyXQ1uKrfhe
ax83Y8P3hCzYBD52rrkuT2z7aYOvVjmPT5T3/sdSb3WPSr53GbZxdFFqktnRNfWh
pwyyIw2su6cULqsv/Pn7ZAMC1Xa2SnI+xSqtgcCreirdA4VkYg+MZRXRF8hGZLfl
I298k6LfMSyuckqT6rORwsQAAoeeunFev0CR9nVant42Ics68tOtTO91adCtYhCf
edcBAo/SKHWWt4FENxzrwuCQSiISunJdbxtgLuw+GxGG18Okd7LvmaFLRhCc8XbT
+red8vBPZPGpVsK6SWa2ldXL0hBIi06bgDbRNKwzjACciYNlJ/lstfggElX86i7/
jhDh0dwv6pVPQZ/kQ1Ekw4n+4cJVyn+G34LgyweVkmpI18EHDhxmrAcMTKDr8337
/4iXcQTWgxuzPGrUPE1i8iNdQnZtafXvlRK8HLKMb31XHC+mpuSmVoZwIQCS5OGb
XqqrNiE7gXq3x9/m3xCX/pGvTz+w2mpV7Z4MKLSM0wtFKSoshrf72EUR3jGFStAQ
i8rDDHze3dIUjq7YJX/6yYI+u3kOfT7nk7SCWksw2TTU4K1ecP960fvpYQ6QdCGC
7EJc1pxV2+SFvr8s2JAtOYCaG4OEKO6bNtio4guKHVIPyj6tmprh7be1v9zuoqk3
hgIn3Gd3R4jvGHOdT2p9v1GJQm+CWhqsxBK/QKxIqsgFGYmd7KIbalWTn92wntJj
NqyNhV31KTvWMsTJch5NO5XPMiv7rGxWl0TQfLg45Kb6ntuc1QeReDSUjJh+R7DU
grVuwbxnPBKIErrXwjvS/Fg+yQznEkxqx4uYAgcJl1/2ZCQk8WRiFv7AYN0Dug1Z
lBvWgvLjjlcvHpHjpl/5b7yzzRfq6r2c0Vj2sKL62CJXukkfQUqaNd6X0O1P8vdO
IZ//6UW6Pg1IC6htdCApiy/fL3yL8k5vW5qPsTeTp6lwMIzl574gVT6kbnwH7ZVj
3TPqWi6MM9nE/Q3Phk4dUi4/qOxZYziqQ+WHFJkM2bgND6wkGJIc3tWggZHTe07N
vQXkG4+yDrbKsut3maBIXF/+QPKPwtm55v3ErUe4mnaOpwhPF3jo92UOILaa0yPN
uJH1P1HAdA1obx7ZJ5KlPT4a4nQlxa9EgkOG5ALvdcd0o5eiznEsgnc7KCe4ddBe
1ShjCJ6ayYF5Xxb32qb+Ichoeje5C/i5Td0DOUR/CRBVZMA3lEtRSwwyVjLOgA91
Uf5JrC2K8MNkh47Gww9PpBrZnmSaJi0UyPA8xtBCgoUqbG5EPZH6M4Pk9eYER/Ch
OBnqW8QIkpKy8rGP9x4PhlD/c/tNGeiRVFNUWcI/mG8yMTJTudlq9HIUfiTZI85r
M8sQtXUt7XSh53kAK1y9hZ7ywddf8yU5tBviZKVixJda3qG3DlKvtPAYcbZQLrFt
DaUJLd/qC5iBtgN2ksguOleL6SKY5lqBqb8hZjNJ5E0KzHvMK9yIxDszmAgd5dXp
CrUX2m8ieTTIazS7m8jNrQdcSExi2shC8ti9CZQantUdfui+dLlfoXA9OCMZisl1
w/8gujr8bVFNp3Dkjt+9GSag8IksAWfAE6EIpObvNX0NxMivshbnKX6f9Cg0aBP3
BzKMRMwfc/LpD/REn6FTb6s1EU93ssORysPHOI5UHmc3GAIRgLY2HZ0GozW3tnZG
t0RHSCTwnsvhRJqaLxJEIEV4vmC2GLyO88ZNJHpQL3MJriVfhjhszFP0WD6CAvgk
6rIkAz5299kv3VFK38Cij9KNR83JFbTYWPSm6n3mCDJN9Y/bySzD1m57aJ2XywGx
oa8dAHFvhJ0R1vT+IDzCaR1zCOuTZs1nb5B34u5E+hRNhyRKELo+iD0UgDf5crdf
Sq/ge3qrsZUlh7DQcHcjo4WnRz+E5rKU+Amvlfh3K7r4hel2AeKfgwrs1H5w++6u
8lu0MI+GqePymxIMa6Nl6/r11Xp8J2e0aNFUxS9V50vb25nsuuOzG1eg3SBzYHdP
qRSwDLOz7Md4bRI7wmRvUM0Q/BrEe2DW5LYqAD+4eMtZn5dafInqxGUKgF5DrAKb
buov3v/q14OHzdXxeAZPAkvbAsPlIbBa8mZlNS+hbPWG+UftZlBTtFbWI+i2FKMh
KXY19wKB+M6FmCkikc0Jk9Awht33eXoPmNhfWBjWh4WVSX5gwW71dXBfy1BJil5n
JralXE7dDfXOqzr/UDUcg9ZK8UvDQ8YTnmUVaVavdxVP+wzWlA6Wwv/tLbhK4/q1
L2c7Szp56VoYHyWcCWz2cepg4O2K4s5wluTn4HSrPWCMnFcElR4CPaU1RuQ1nC5s
BYwGWJyMgRutFx9MZNxtBdD4foJ6gGHaPeL7M/PWTLqKP3FxWPzPwX/LFa0ZgjDO
7LcS+fua5Tukq276+Vezj5+NzOnKEY/KEUJ1RDY9hP17BzPAPkFUXyW8dMiK3My3
QylhC7HDwpHhP6SrD59w00wSrf9HGxtfF1NU+/k7PDOFUPyC8nF5rEtgnp3HXbI5
QBcfZLWXcQqItWlGWkZ407AQCokgDwbWptILHFnKBDzftT0mQ940ycfft1QHoGPt
vavvAfgj8BZt7AUwlBjw8F7N4SJKSLP+L2RRNej4ocP4k7sobnetJQqOH+TEiEfF
W90BF04njKpQ5+89ces1kK4a/Th7/Lf+73KQjCJZLE1fk7p2pEtsLXKPr/GsdSs9
v+tnips6ceY+NwUAgxUUuH0mP/Z/yXAoU0rgq7ru2tWADDXBfHyggjsTxREXPbsZ
tM5oJDuyqClC8WlTXHvrksBrBvznFvpAFEI+dx0rinBt1cdXteGznfK2eAR2krqj
lI2YqoTTSNBxYVwU0o8db7RI3P9vr6H07tvYTG8VvvO+uHpIzxXXIQZqUmrXitxS
vb1AhUjDi6C8v5m5HgJXnXJo+DU7J+7PaTO/2ih4Vx+nqyzVDQz39xKCPZ+UHknI
ntnvrBqymF+7aL7ShCxU1NecfFJT1LfgHpSY026CbzNk9iDQfhJVWf4AxdlIzwEm
4KEE6fUP9VKIKAemi/GyEVZLyxkEuPJbc2N2wOw+8CgngtA3NfoCu+xYnNWQE3gs
QlRE/CRtlUzREyC2sOd0BpW777NFTChUtgHiOWWtpsUwLZDYl8XhGOKgEBJIgpic
UWIdWfthufYG23bZVhx6yudS0QgndUA7ENu6eF7vUUJLSyj6DxGLFyjmdD7JKlZf
H0+1I3aRaeBbLiijU5txIKxFvUPov9HgylxV/+BY2m13OCg0v9j9tCGE/I8LbdaW
IPZwqBHPCbk0Iqn8FJ0Ms+NJ5GArezRGPdpPsJMSllqyKz1kwdQ/0mjVQOpjVxkH
nCJh086ySQE3amUDFp1VAKmaOoA9u9UigOEYnJmkAr3ksx45WP4KZ5QGYSJe0bq3
hTHoOEYJ9HqJkVjToKkGtARnQrhFM09Mw07R+Nq4u/qCD0ggM1z2ZbcxYZy1l+IR
83N9a++kMCCA4zPiDEa5NKdzrpuARgUQi9FkY16l6oSMaC3zEc4aFDRtDFyEJ6/b
2fuKRktXuaKxELElmUDVovGvuHEOz6mbIcDMWuigP1gfPVZ5mmmrQtS7stulMqP5
7+yF28d8csg7UJqQNrX9Cj28e1bcwZm0lVqIEUQ3DdWh0RSWVnajSx9r3nv3qqd4
NDDT1tGoOCGwSuQcJDv1IFiE/FAc2HOPF6fDom/izihvw//TwykqZFZYBnnXmc9h
HfHeAr0xlgyXNErUKohG0NaFHW2GBfcnDJDelY60L3i1OgDilGelCrDVrEz05p1Y
F5aUB6R3yZ2HVngER3QloOtFMzvVLz/alCuey1V9uPH4A6EBx9GRvrFV57Kiu3Ap
cppQhr/d7K2iFdc9saUhUvRBhHYn4Z6CCqry1OHoEvmIYazirqaKPe6oVtkr55rH
DUTsoz5ycqW3XCjTQgL05GCOThUSLVIadx4layTBdZX6T3UP5ilmZjlmKh5mJK8k
sMKL5IVIkALEJywBK2QBQpRdqBslqlFKJUKYM49isKyPOdfqmAKMibyNVZGtsUfk
MQLbOJ05jKR4RHM86ZoVaWZffLfDsitY8hDa6kRLXEZX8TYOrIv8CcW8AwIojhac
wtr5l3ROoEhzeUiNL8qmhT42zjis/FSI8wc85qWn0JZp8DAXdG4onNfp99VQSRr5
VLYPrG5wNSTLbcdXRcNDASQ50QzLAXd6oqxnyx5c7hc+wanD00EqUrbLbdqOHYFw
VOYOZsoDI/34C7zY4IFru5G0TVn/uVeNVCxLPLeYpBdXMz+LRw4erA5XkAfHdN8D
61f9trBrvGGB4Q0GXyhKVImCOpVDuqgafG0LPww1YviKjLHvTXKKyEHVb9gF10Uv
++yIkLXkcxgluPOhVeTkqNBKPiCFqVXqfrfYPz36w7ooFEiWz8fAHoxzVhX6i2TL
NAkYBU89LdnkFp3GXEZn8cGIn2RzPWztbZy52TgiGYIhBD7wHsbnk4jFf7W/0wFk
9Sv+Bd3Eo1Ke3pbW7jFC1nGuzfcfaE3o0IjFJ55uUmC+MAUySHdjalHy3aXBqDkW
9lwyjJXY/gQlOeNohFbSJgEW5U9qYh5YFk/FHbkx0O0C6b/YNsHghpIRm5b115z2
khWKrwIzp9w+WNYQAPtalvlvpVs7AKSkK9ossQaTKxEA4n+Z1urvYrzBMGu3g+LR
VIfTUkJSFuNu2x6C1E6gHkf+z34ixeseF1YsvZIvrsCU9zflEBdSe2EfnafKqELB
Q+y6kSNbU+pi5XSfa9XKArpWW2DM0O+mi+Llg2USgFcav+xmhPbfiEvnDPz8ABxQ
Y+ubUUyLjZ0RjXOuB/9f4sHlMc/7FLPCSmhDcMRcu0oeIjr+2aXVQ/HGDA70BngJ
4xsp11ZF1zAhBB+HdMd4Y+r06iUpNbLfX0YSyVGuyy9GROtKOvmH+nZzkXiBg6fu
aiPGb09c6q6rwB7WqUGik3NsH3d2qt6uJz/c4WYobxTEkGiydRPy+PsEEk3sFrUs
HvnkdQubKzJxApEY7kJu6oBqn+qSz7mla19fHVr0vc61CwsQjBUKnXPov035afHK
LCr0Kf7J3TAEHSVO4phZ0nteY9AWZ1Z4hMH50tr4iv+TxfCdN/SxD0GJgv8xyHYw
N8s5Ce6nALq7fVIvn2nrludhpC27Q4+p66XVEvpjkbCyVXGzhSWW3vzqilveoAA3
tIiGgqw/hlQFGbBDyCZlHLZZIeSUpM76Mqpn4yKO5D8Zo8PrnBNSSMbgxtQbWA+q
cq6saM1bjRdTmeAxueyBr0aP2dKj4kmEiUloszDySgjDpb47uqz3dcfzQAkEbZX+
GV8tHLJJ1DXWKh2AQGTjfKOwbuS1mHH0Jez9qf3wl8wrxj8EZHbHuSdP9ogHTVn9
ZQ/sJB3qDNBSyVHfeqfSDCXxfKDxdf5Z0XiUlVlQwCmR2mbsh3JfbUbKRrntoWE6
qlKTf3IySkTlo6CcytON1G5wLsrz5E/+GoPa82YggmsMHRYCfb87f2FovGZYp4AJ
wl6YWOcSP+H3uXvd3/DSQGeQP3ieLXASMxzhbSsFY4YhW+aU+G3424ES1zkAWL1J
qQXyr3VL2p9ZheLmIvnSBWKVif/wN8TI5ptmdq/27e740JNSurXV1Y/LWnuYw44w
N+MZnOQCh563LXwDgbgup0H69P7Jqw2Vj4VvymL+Fo9wWlxIFk2zcjBE3Hk3cqD0
G26vcpFpni8RHNKlUT8hDNmK2KMNvhjO21mCIF4JhSvU1WrX79ITNAB3ePbGL71U
/nf+03wRTXz7ino9DGJSahPfI++odcY1i6QnrT8G7IXM8QO5M6DEPoEiqKQ7V78l
/s2T80asTgGlH/kB/TQTbbTdir8xAe2LKL5mLeQOlx9MrLO4DTndpVFB9malJO2M
aYfprQ8G/SRFcKkC80CW6Qzqat4Ukjv01eGyuBWcHkTpsQHN6oMLIyNg6FhMvAkl
aBMLW6SIb+nSLVU5L9iHXkLoX5e8JpUBVaOby/VK/kujd/3Co7Vz4SKG/oQA2taq
SMefAu+642wirKixvMYMBQVMOw8Rx1okdMXignzhao38XLg+gsqdCRHa9t/f+kHW
vJqsN/Ih5x7yR40XNSZSNwlFgjhUv14AI0/g4m5uv8n9KsG/v9KtZEzZhnTVYvXn
3SPy+RI2zuzFAO5s0TG4gvWo5DdDg6di6cawmBzkntQqMebgGX9e2cg9LrYZ2AQZ
lgKh3fBt1cMbAd5jR7q98mg43QHeGYMSpj3qsLkLjVQtkjCUWLj3wijBJRNbQzNO
Z4ThfHUkP/jl1BKkzc6d3kXWeX47Y/Su8190DjfrGBSMh22dt0w/BU+FG7Pu4+S7
KOMj26jIvAJpMgSvS6r/AqubdIHiG1H6Uq8abCGYiHCZiRL/18aO8iEJmNRFU8lm
qk/6qpC5MTFXCdZKnBp7gvQEA7jfmbpL/aJI+WbGevS0mcxMeUvpmeaY0Hz2q8Vv
/XjvieGIw1PzTLR76XNLIPAyOfJ4Hlis1waaP9a+iknRSr36abZPQGkZoG26yThD
I7JtfHIQMmzW53ViYPCNt2OqK4bJbXeoqwFw70JLoCYkIX5PkyWehQ+9h2dUhb+E
5nkaXRjV0Yq0QElL2fyQy2O0xy/ysAxYWvN3qMVMhTDjiUwJ02FOeedf2K1sF8D9
PlLRl7M6w5H25dr7TSB2be7R5mBHy2Ojy5Nm4N32AOEL7TGG1FWHJ+Fxzk0GknKE
vcvWrLQIn0ii0BPvugwb8pNfrXQiRf3V5EgMgbLXZERAfvKbu8ol1hf9jKch+MMd
BfD+oqGS4I98tedguUOQcYesG3xiKJA+EhFU4JhvVGU2qhidvKZTQmIJRBS8y2yF
iOGamR7bKE+G4jg30AfBkvXe1SQHRz7byYRF9ll/uADpJ3Cdrdfm3av5ifFQxAnY
HmLnlF7VEyxXLhXzJu0pTvT22dz7/fdjvg/gzsghomo2BLjjyuE20/+l7gNgD9/s
1S4Lkcws2s5F66jK7U6h4HP4nQyRAjQNIhJR0q7FboFTQKsITEYswqrJ8hJZ2hQw
yZJD826iyPKK/0NKxVK5jy3OITmnWPCjRlg8qGLbLa0J84cgOGxKupTjUCIgMqMO
c4TSNeFIe0cV4hRCG+O3t7SjhrxZPCJsvWTjRjzMYMqmCwxr9KG5NYBFdsWtlokg
VWpALQxdioMLgbKy1zPdJBoQEnH+5xsThabXzAyvv2MqWVgVwPypFM+U022Bopeh
bMWlrSI5CIDZoGb3ifithU06RWKrbw0r2MMqT555r/3xhQoTLdDcKM/4uDEoZtzf
ra3BfvftfeD8PMHJoFxPZ7gzyYqr4nIHRgnqud783gx5UCq+0Ap/rpxLtD0uZHzD
weWoZC7Qzd4a6eCrBDBt4MWu0ni/CbDDD4zT7SiN53dzuo/r3HlpFc6J2lLKy7ea
iECafFPKPQs81EW2ZyhpYr6jTRlEUOn8YOsoWiXY1f6vXOIe7ZgR8wZOojgrXrb/
e+wRXSDZwNULgrAYJKrKfUKmHXdJ9KHNlcEHcohb/rqP+8fKFKco7Q4x27A+8q4Y
GaAVyLe/BA8I5sjxXQsBgQ1zPEkz+ULSYftLF+nLA0fgiaPHnXQbsyoFvi1x4UCv
44rZgiF7q7xdqKgra/5DyKWlNoiUe/YU5IkGZMPV9EYdXV5NtLfLiLVbyXyda7KU
EWqHt8RuJ+H7tBOvi95a6w8vyh2RC61IeyAdd/uyplYq3RJ8orYHIrXIk/0rkaPI
FbMAPyWTbjHbwBC8KxvM/wAJr0dvJAkrYGjrSoOXRp00PnXYfo23SrmPn31y2C4i
ragLHlw6EHfqvNXUpOKDGoYy6I7NnWgDxnZ3zZHNYOd5Ugyv7S1Po+U/mV/1VDKc
o+ssKJtGZKTgXQZ+n7FVFEi0oKNMc1LwQQ+URh/3LzdqwRG0TtZnAjx8+8/PMXjY
+jU6cSwnAG4xz8/H8t28HVvbt0V5Kt6MrSfXSTK/m5qvPBNggmrERBGWpNDBjSx0
9ynDJHhirThSuJzyjZ+tIPAiTUsgYz6di3vetnpT/b7pNhMqU4SATcmhdiGVPU9g
hkYtEQqkdOpYJnBxOz3mqV6uP4mRdMC/nXhn2pGNP0IRKhNaBYmmKqDRIv0iS7lR
5GnsEdK18XQoZCkUPZvL54r3HznX6NgZcRGhngS+ae8URHB/WubMjmTSrYElbo2s
efrLza4Y9sDciKAT0yPz+ZNMgpz3Sun/p0TpdMZPlQ9UGOZXwsEadB+ecGPV6PVt
SWlQ0c2PUYUxsIE9YP/2im7HCX8nqDlgt6bmmBGFG8wunoCKO86brGD8/du5LnIn
3MDSP5oS/ilKyNbV7lrK+65f+NHM0bAAle8uZf0DkbNvdtqGSno7343CPUIiuuJV
H4mYMbe61LzHPfERlYOZ34hQH8RYz337UuswGK1MK3mpucvtFrN5faFUEQUIdiIt
fapLrjfCS/xHqlEzvJvUSLjtfxWjTpflW2x7ctJyPfCyJb8THtrr0xDSAzhPajq0
GbJAefHjMWwS7Qy2+o3ayrrv6rExuuxB5Y78uvW7kz1TsIDsj9q5R9p5nuUzZWa/
ZB0L6k92oYd2Ec4aaLPMGp+GcSSiw88sZy/2XdrcmUZlSlJXatj4NCs4rMXEOPNM
+kx/QqfYYVgFw9ZyTcliBqlMNHFyPKyiV2WIogbG49cQ2tnxUXOwzhbSsbHP08+I
hwz9nOuzJaeo8TwcmPN3r2yZ6gfGrzq9CaTZ14vNX8THyqB2ye0j5rVZ6ddF0DGy
+VB0qHBqkr/XnWcYcGs3k5/jCJl5oKRiDkiOTZegXrRHCVd3MmGOCuQcZySvqcux
PKkNqmujPSGV5r65Z5RMatuJ9cI5nxZMmpl11pNjsX1q+PhnrNMOzJGFyFn43sHF
EnMgjQQ9es21R2ui4YCvmvAa/i7GHM4PSBGj1Ua9uNCU2AmWrpYxW8ws+DlLPkJF
v10pZ51sahvaz3Tfo5N25Q+tfw0V3OQ3giD+kX93gXV4MkchES8pnOjmhAhpFYin
CB3hLBl5jZ1NslNGnwiNCY24tKAFyTAaKGBMhiQ3xmTixWyimnt7T1LAYNiTYBAK
d7aTGpEWQBwmR9z+4Qp91Q0MmvzK80j2amqprnGAdHhtHVA0APU+Cw4IZIYwC3Mc
a6f8vODZBkfO2C3SB0pPsatP6QrBW60B0hc4yyiT39efj694qek0ts1JTVp+QK3T
Z1vaMfwZN6d1OrzNu86ft7C0eXn4LT1KBZOJjfa1c1ersH+alicC8UIQ+Gs5M37N
vcILlxHVe5d4Fe+OkaHsM4g7FsZB6mVAdSbTVQpY/MmhWRnm6frWNS8IhRxqXUKQ
5nu82hQ44YL9isXRIS3hPC8Z60BkcLScQ2BsVbNS5K79Fp1Zy9d3N6qvRiaJoPwJ
TQ2fwrSNOfxCtRVFR5F06AHGOzOSOZdmqD6wgh5GpEXuLkIeVGJxaS7EGwRxfnsp
k59a70hTm4Snb2HDgfbV7AwNzpfnZrEJTkVwnst30onVKX1P1qDDYvjOO5eI17f/
CxwT/8/fMkq5YBkfPZ0y5K/Q/TaDVjmq1s7BN05/7Z9JwlZHokogbcoTcF4hNnJy
uU61eybT8dCKWzbwOhhwaduz6CEWKzGlf0NGwLbAW+Tg/vhyDpD59keHf7a5/lfu
N1Ut77L8suBX7m7PE6I8I6GsufBDjLH7GBUXht4u4WAIE3DuGU0Fx5aGUXETqR5J
kzCD8lhb8kU+BmxhB9RKGghQSpnTpRPfleKKXfKhNKPHetZaO+nUu8prnYC+J96p
Stk0g8m5I6E+ptM77x+UZrhbYsgD6ilPDHI9SgJgDWxTdB0ZPaWl5QLUDTGg7vtC
YeMOsiQokMzKW7hWuxiq39LXRD4zmNPhxREghnksMi6SEu0rGHEJ1iNN6MiIO3Hp
0gAa8M3kJx/Kfc35fpcr2VswFkr5LwZkAF/qLCOHlnzJLK+jc3ELSTRIew0/6Gq7
V8hL8NYTwhcu8pYo1p+VFW7Efvm7rsei6zQABNowRZpl1PRaNEOjYOLfj5BlxPrb
WTbmfdrJFek/WvTOGM9vCewQrFENXmyeB5urSvQuDHoNhExEteweDd91Y8xUk17D
57vr1wTGYDNBxQIwtWm1YpnGpm/nssauf+oKHepr8qrkiFFMaaeiqUtAmtMyXqrF
jx6HjBHtV2Q1Pv6pjIYjmr4O3yrod5ljVUXWr2oBVE+w9Gd919CdnM2eR34psrmv
sB2PZMf+nDGSpiER3Hs4D2hqIkmWvFOFPmM3B6+X1gpV/7dh8PdgwODjpjgZkxf2
Kds2rwezy5vnI1YLt7Kt7uvO0ViE8Khs5tLvJqA4naiJ5jTK9OGBBwtaqzqvDTDB
PFddb6MBqWr27DOMNpON4KKWL+YQ74oIAgA+PFTuCkgV5YfDgSeeOLCNrEKlCNn+
RMAC4UtNZoY6fiv5fmxh2W3/tD+WCNgFn2yAVFHxeuJ4tepxddPIKpXN2EtbrJac
4H5gf9XYNsKU2SENSljx4xCP8OLDqmbaar80NnigkszpxCUqAIlFZSUq+tG2DjZu
LdcY3vUi6TbmiVzx7e2i7SGJFcKdeKRbd0SaIvTFKWkxSSmPJD520WW/HpPyHrTX
OP9saqhguZY83odPo0ch7NIHHgr45esVryHdBoVnX4vI3ZpjUgAq3Oxn1hM75ybw
q3c/aO/Gd7cK4yA/LOl6Qrftj7l7ejT6fIImF8cUfNapPe4Ps5JeFas9aqLgo23L
3QHBFvHrh1mduiUE97ZDM8+ZTzioV4DRn7n4MKXVJL1YSAqdiqLJMl7ofMZTgz3V
86d9DzsgOueQEDr3HjwUi6PqJFpQCryYA0FeP9kTrN9bKQBi/qJAIkGy/mYtkmp2
oBcaT3D6x/wfFwDh8JMTMTPVO7y9slPzF39UI+jRNvWYpxbuBuMzjyHYqfEuAE31
ZZEtqicYjkxII+eo08xPd94+TEfnXAV6b6+b24idqQOCyg7+jR4FO6z7MELeAH9H
3vdQLNmc9wAXA/cTVKbIKIOEgZSi3CnKW5duYXnX9kOCATybWyGWiMbdszsfqbMV
QuDITsP1lsgJQYCKc+c2T+9JHIiTejfuYwuyzZB12rZ8TK/RInjHy4xRkUxxcE/j
ah9ptlbwsdPcBDQGHJ3U/ysD7rAczu+sNWElnR/9lDYgvF41iPQB18vpVrh1ivA/
SEmiqH5iaeCupRRlzzR4eFzqgtC1sV/1u4Rtc6sToDZ5CqXRcZr4Sof94RtqPFZV
xJN3zL5O4OwK1xMCFcjUQt+jRrI0k3lLO+rvwOx0I4ydT8s8g3aZAj7z0VFJfEgr
TVFONoTxtFcSSV4GneT5adZsQdm5qMMOsOnuo3JsdaNzrIWJc2OuRoUpxr3ZuJKl
didOX3Ovhyl/uH30U7CHy9moacwTOjsgvh5YqW6evf3jIRj6SromZ9ddwOct6BPe
GVACZy820FOajSZ8a1TUCOSYNosqUJikg8HCOdUuOW5mpO9gmv2+F07vp87mhK9O
SGoMAnmCQn7o2DrouJu0e5pMz4mEoxthQQL1C/jhKVJTTmeRfvVcMWHaSbKqg1at
eU/9yMbSzKtLkn1PPAn+ieNEvUl52f2LwAqPnhzCN0qlXV0VZwe670/ekJ5P28FY
QwSkdx4AjHo9+2FITQkysahb3lx4ZxFJuEmoZTmVeJFfuYEIF9itb1UEwxteZjRG
qDBmXUEPil0I75x8mBBRaKt6xW2lYXxV0l4gUrkvaiHtq5YMnMd1ykzWprHRdZzt
V3LKSj1eX77KMa4iPQVjiDEwBeqvUeo8Ffhtpl5Y6qzUTynrfNra2LnG6SD1bylD
P3TRTtqZiqrXzwkBH6wLfpt15A32qCGHogIPtN/N1ON2Xlw1L6Vq8sYUi6gDvTYl
/FeiC8fg5NX4vCfXMMbvTAW4rG2SrFkm1ks6Lcvx1Xcgv5H7hmRv9meHdqbkxINa
cFXospkRhOcJp/IPFSA1Y/qx8vvkDnmDY0trw/9+gIxH75WHEqBl/eQVgxZxrZe1
ZnZgG+dlWJbYqtIBFRdlhJCqWtjChEyn4WH2W6MyvNKv7h+0u3cSH3Cu5t+weP2I
4jgncNcZQ3Z3ZPh3vFQ4vnDAEtZ5Kso1InMnrZ6iN33/SndOaerAca7EEfkXnDZj
0IqtyZ4H2TlZ7eu/wn/1cEZataVVa+tfLoo2oW0dIN+C8HLIlqty93OgfD4/NuRD
Of+QGtJUA2X0t90unU5p+IUrygS9iOobtbqKg6uCqKtAnqGEy1zDEGzQq9WVDTD2
HWt0oasXFmqn1IC7o+BW9Lz7XBBLHMIIBdHWq5irzTZsuJzmaROU2NW+mrsTLlOm
ritbo8FaL/er6HoqqOTl9oFV3HYS6RAjJK0LwWQhLuJfcgqLInBer1YWKZODsYEg
gaBRxW0YVpoNybcedlGDHRTyHTlVCtxT+TX7PFTl0XxzfTg8V/vYTYpaRJ42io+t
4j7aIa3aXJJWQpiE8uQ3NwzvSxF3WIsnYvneadny/bfCz0bc2Vo8urM0yd0s2cZe
dVz5ECxJM45G3ZU4OPV4KOwTKrCTxJevkGUSSwaF4/Mqro0EA/eubtvJ0uYES+cy
/oy4caPMIf4o4PWR4vC4wOknXGUOoktHWZj39ENZD6Ap9ZG0020D+nwNVJlkT5TG
mWhZbth5w4MFyl2axT8Qu83jMmz1nN8WNrY6VdAzXpjxFg6CFu+975jBt8t0epza
GAXGLLYhi+hW9FDtMs4gqRAmscYjttugKeAZiDQ7rOUZlhOFBVMvzIWuLweXK10b
Z6QTNeZpkT+ioAaSWPM25DTdyP+1HGUkLZ8id7KtjvuuAjGf1eTYq1SbOuBbgXYB
/R8RKJTyfA/8QUZBfatxcLNOTThn4P2gH6MN1NK11GbKv55l5jnYfxsQewUgeqAR
N/sZ86QnCGCJvlGrY5mVZtQM/ghrtXemfZn2Je9Yn861wlckwVdrwVC92/+35g/g
HtI1FV1ZyGJBU8ejoJJUxvBG4J9zOO3NuCIth8CmFojcd/DUCXlK23hKztmTTd2C
Ze5/IIq3sUHKd05BXcncRWQJ4Vlinr5d8mfLNRVX/8tbkncLPl7D7EbJGgXCHRQA
cKoWUh7bLbAFV88uT9g+ydsHSZw42dXo9M0b6DGaaf1QvVDAFdkg+bepC8+Ron5C
JTdyBCQBtbsKa4C6ULrqwILhZ7gmo37/be1MN1g+1swwrulOcOUqUAiAVhj0rAoY
KXr4gdRsj4ws3hkOyOxuWTpiF7lFcS5PvbHJowIbjiArSN8PBAjch6mlxPn3slhQ
QFdVYkRcIxWdwh1zqCDoAgsU3YlaVdDGEvSv+TpRkcdIMDO+NH5UzYn6srCoDA7G
TL2HMVYWXnCo+wQu+r6O0MUyLukK2yrLTcRGMkuy7sLuhJSmwuKKuDt8Vvzdr7Hx
FLsYytmdV4NetgYEU0ne2edeFrAu+GYhWaE+JgpK0TqbrpAQqkTKRi3vfPfR/so0
38NNFfcESvvd0A1LDyNKAvpIDWpm/7SM+/f4HswTEwLltrl48Plk8fTRE7dZ8hGz
gyUWg/aZHfpmfNsoZoWnjJxVhF0bozK7O94/wUIoDk6+23MzASPzrjKMX1kkxpfR
qV3Jlmtgj0z3N8C5c9w4hvtOUPQtmsFLbO4bV12/vE/3JkMZaUE73Wbh1V+IdVBk
HcXmcPYySyHUlbjbaji6Oy8IBo3bNsBdURe0MvqNgLGsSM3uLJ9+wsJQnkvZ+9HB
j1Ar560EzQS3FDoVvPT8q9DpZ1G7GkWwXiq4qyr74oV+Dwbk+J2uU5/Vzh+aepPj
vkF63W9oL5FbJq9stSsXLr62gxEYYoMZz+qKS63U/fNN1JC4TpPu2XGtEfdMMeKZ
D8pZcbHB2woCx8iK1A2HDbxaY6WuBdx52OtJcJDwsiclrsNWjD8p/dXc8iLkA9Fd
OjtkAiZ9bSv1EsUEjczVZUB3B4ls15sU5zXWDbiUh3Yhr2zWf7jr1j4CDJF2TClc
bWaDeRYWJRO9+Ld+sKg582T+tgxwBgPATMjzgXFqjabbBCMLHh2nBN5GpjG/T252
wzv3LClbqEVAx+iAGPjOM9tZBuXjZBg8usI/cCi75C3yx2GtIFis+fqslXB7hgSa
aULqCbNdluUuu3lasX3CoxVAKnTbcr7WrJXng5ufnDvOypaDtGOqO7harSmGzzsP
/Sqpjq2ALUER+a8EvjDRkTP+haugyM20SFMBdnR5Gr+WBnY8wmtpFm51XIUE7TFI
R25Bi4b0MIAJt0slleAd9iZmQ4sn3yBnSQEe765NFEah2n9UtejTo1tkUZf+a4qX
6lNbjy85Lzm/omIf+bMrvWSmbkkYLTNvXdOQIVGD7XU/ylN1n6ULOPJ0pkfbEJXN
qwA++7V6zJaFr3kYOWdVZljvD7CZgSV2Pktw5GqagbRkQc1t7ReWl9ss9HKZhNst
dI1zXlW9S7NSm/LdZXzdEaURfdTmgwy38sWVXXL1btBjbtZp4QxWgpsVCnfINvKa
yLvQuQSRNdk/3GY4NeK3vPS5ex8vCzlKLc3rzuSNjBo8XUTRrqbDXaaqMoiKQEGT
I6UZwtZHF98tgrkaVgwKsDHBilOB0nMVCd3zL5c6O8OQBT4NETQhHhZ8zZLrjugj
a1dM7w0skCYJrDfcMD6bgXt1G5oUUyJk8tBUvYsnfJZu5xlr86LcEo6Tnf+l819q
+FTU4qp5Y8eAEXyizLQD18uFRRq1dI0FVHXZJcFvYBXJom1qtoisLvE591GTZvUy
iEEK6NP9JkkEYGhfIPDikuAkgMv+R/8iiHcfCmC3D7g7AMYA7aJT+pxgTKNYfgL8
G7qF0OrXDm+15FXGNhTX9yRq7Yr0YTY5tQI4JcYJe2qr4FZS90BRJPli6u/Bv2Bl
rv3IZcZ8u2Ti1u1F6NQGGYq0kPuYHqXQ7gXeZ02sM5YGM6tN4pqVd+lrRih4dPPD
XgPmNBeY284UnVY+k6jJ33Br28f8TRbAONylOn6Dzc96csfrmHyOnQXNeQRHkIxI
iWFCbCvg1p+7EX9PYVHKMqsrIXcOJMnC7PFCa9o9znhHGvHPt9EMPDtyKBt+GIhU
YqUoN65TO4YnS4Le23ee2x3voAFfH3co8EItYKu0UmIVfNSV6UmJmZkFng8VTkY4
F5w2LwERie3ZWT07WUnR9GkgYAf7nTEGgHsJT3JEBojl7ca6VZI/pTSauHyMOGPC
JxQL7f4zON/JsU4rtH9iXV+kc3YRRZtVeHAPa32DfhCvKrY1PJewbqdSm/CxSNt2
1wAjUiFki6kO9xX+5H2IHM/jEa0eEYC8KvoX48fCPYtBkV3JnKganLDDxRdkkjoq
GUNDBqdz+Mb7bvWXeg6ew1Bri5X/wNcmUMHWbYKCytnDsFXLtbL73WRpcfSpJTAR
ECiZIhEl3XnYRY8x58yU8CBRIF1d0ye8jBGTOVWg5ngKm2Pk4CB8rigmcetDjFRK
00tHzaWMSZh/6qlqMSmkEU2lsteyzcfmh5lrvVV4SRdkEWu0sglYqG+UhB1At4JG
3biLq+ZMsnta5smStSnUL5vhzXC6873MurMRNkV2HXXHcmnNO1k9J9AQg661Y51u
N8EXGuWzUVPPt3VIymPeBLmRn4B6P8fi7WKfqpVgETKMtNE59mC5PlWeoNZpDIH9
5iZZXpbqgBZWna/BZ6TshXFz5ELa8SHVl4Q+UlLTMCfngsItA/EImzg0slsJM1U4
Oa1QoD4u6zBaWY1FwGTdWgRXsmp3XA9geK1xE5MMFo8jP/enjdWmyB3WR6xh64ju
5bkYbJIC/saU/IyKA6V7BsyPnp+D5sBgCPV/pM3QTB54R7J/CyXFfE2l+JQBteU4
s5xSH/YAjOM03CU9rsjZBA==
`pragma protect end_protected
