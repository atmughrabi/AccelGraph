// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:35 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Lzo+bT5asYAbSwflqaOUWYnRzn4/lY8a9EAlcNgxb/YycLkF10D7v6cr1PbULoHx
MGsqx2k2W8wSUb1t6MN6k6j+wrquxFa2qXMHg4VIguz3SI4I8UCQGwu4NDaTpRZg
QedX75fv+eVZCiZdZx9vo4v56FhmkU4SlPxC5lqVdbE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16976)
WBFvFJ2SVLnKYjSCpZFBMuOanfVs2vjYnaRQWuN+6cp8JHNrLr1MLy5/Oaaa3trC
0GtYC48jnl4y4KDsTut35zVVMiDPwNVvi2dOrmk6Ol+EV19i/HW6ZyKxPYk5jzdO
aDThRjQHz4Dvr1tLT1P9kYr30yuWdjs5OOMmgJOLbDlVu841hNhZwBgJQY6C6zwD
W+ZMTMy7tSCB+2DwSSp0Hmpbt90D2FEA/FoOUl8w8A4uucWOwFD5QxTVxd1O65yF
MR+gWN0+B4tQ/D4p2Ry4LHEPXlXDHfJ/Gh1XDWTFMtdmPdb1j9LG+2TJfDQuIluI
cd+rgf1BeZGOGHcVht9qb+LZlJhSOUVcFjtkGSt/+DO+qjXfPtmDR9R6lE3z5Gu6
fSEL+nZ5AVUhbB36y5adP7HFGy7XjeJMRzGYppSOfvFLPznEZqbI86k3/AkhYTQ3
7dZSdijKtoCcoHnCmmmhsDKFzrJwEN0TieiExf7l+nZWHKZ23/XnMSdPHay93g0t
WbvHbsO2YKwk0Fb3Gv4reHoVo24Dx/HzorJ9JHud0+zJoq2t4XmwzDrnN4jcIyre
gQjSw+apVaIKLPAFn3pfptFOtfn7QvWIO9VS3q8MsBaZ7ImqJPThSFAAe+H9WW1p
Bk3dB11JOZ3vtZM1D4eXqxvUPa7zi80nS9B4hAraJRGDz+aTcr7YuOCNji+0m2NN
GOLvuVp2jf4dqVzHreeWjecX3P0JsssTHLdkoLxAZN5vnvEWxxRu+witsh3G6SAa
JgSb+6XNG/laCKbl62A7uV9DwS/bgjP97GcJ0+zC19KpULSGcnKlcsMD8nlwvIrD
4jDcO5hsntyh01iZcwKbHQRzpK997rz5HTMXCaOn1k+eLBZFqUtyBkfmfpIZ58SY
nw1Ek1WvHgD612JU/x/j2/auHlZNKYqdjSq4A8ufz1PTVsrS3rnc6P+hBtNBCyVm
RrrcCqOARlT+cthsvU9Y/peAesRJjOroRChojWR1DtDz7sqKnJ6w+utJb1gYbKF8
UEePe5es2RgKFQFjNXdQwzCd2CIQapFXyvDgwTwWsXaCNIzc0nPjkl7qzr+/9nMG
OCeZc0Ru7zBp2kw4L9kvC8LtEJkIHKD9hrzIuYnTLOxn+NQaEL+udgx0DpckAp6+
cjj5ssHbhXTlQYk/hoKQN7sHTaZVkunQEguO2cmou5kYfx0uTVz/GehueK1+J8Ic
cHTET9/FyP/MELvP/nTRhVWGg95Ux59jzWkanZ19W1NzgXRU4uXET2hWPvciFzqv
xHRe1HKYCnRvuG/abuu4V3OA8OwwPvsQu3RaGXWloyVAxePuv3mIWX46dgzk80D0
5ksLubsMcSy4+QErF6eorkws6XZBlIiigvnn+D/ZKsUpXYgAPgHYEUawScNIRbJg
R+IEOdOSMOdFov8zDh6G9MJGRIdRCZmeTvkUiGTuNv8eiIs0PIMgwaY3/aYag3nl
+kw+4SYUp7pvHNr3f3KXjIs02dRRJ7rBZUvmq/55HAtm1dJqJ87L+7Cegr+4sBDX
pErtcEdQhF3B6h7FClJQDmkhx2gGvKh3A8V++UY1AtycF6MhwsiIvwe5DA8kGtkB
51PmOipTVCjAEYDEZgA7CNeHgo92MnugBiUAuIonswhntxfnkzAgAO+fS7XBPJFm
+9U9r1QXXp8Sib7WkZMrICsGgbzMj3FBySOfvqoztWu57w3DsQV1/Qh+sdtsM0ZB
tLRDiqtWwZ9isdzrDlAhJ/WRp7TF+VGRb2joQzbysCOC6EQQkaQ93n+Ux6WqUhdI
Q+bcr7XQtTM6ph/vnE1uhW0HXAJjGOdysYVd1UOnOY4WvycRQAcLHwyVM7ii+WHY
dNlImkjkts7gGTR+q1iXvZWgUCaB+fTIIiuz0TD5yOuyh97gm661w5ceQom4B7Rl
LMpP+DlFTw0UmitR7kgHH5+uigylapXwhfCNGvHzWC7ONwxEZx2w1PdJ0DPhNG2d
KxyZZq+nQYNJBM08dBgzjqefQh1Ne7bCL5Cd8nLm2co9j9nr8cdxGl42BV+AdHOz
Fs4bKsL0K9l/36M2zo5hD138aTmaB4VhB70B+6NniHB7+pxQrr/KMwFpH3+2fkBI
nV/2BItrNxu/nJ8fauwKLYQ0355wPPwowqESrDggtXy3J5n/tlS77xNqH2cu2X0n
Gr2lMxAImQtwMvHgQw2kSd3sNhqTMFBXgnL1Z2UNgYknt6snX7fVkaOcYTaoFnWY
xF4ZP8Jm6eJISzT/oJrhW5dOrPvScT9h3vdvRVWLmTpJUGo8n+VoONsnVILltK2l
4Cb4RLZG1d+Ka+fZrXcsC0wTnJlZKYC7lBjtAqgZKwakoXjaB2cTfjo6F7vbKq3h
P8eH1BWxngTOuQis784Xd410i/3l7DsjpKLYg0vMXLivX1FaM1wMbmh25MVxcOkD
5QgGLSa8AVjVp+PChnapWprsBjNEuZXXY86uMMgX+eNjFF+6RZMF7v+8SzF47W8r
CCucjIr/25x/8x0RIU/u0FAE20WDU4YTGI38zU/6DVB5tp6DDa05fSFIib75o8Bn
lO9aAip/BLX7q6NwBwrf63rC7wxi+DljNWqy7xzVLUK0AHZbvlQFctJ2J8+n72Dr
5fQpw+/VCOAldzPrX+0hTh70GXRAhzByChhv928Ps992i6ZOya4T2eFTdZQCiBSf
CRVpfZvzdM9USp5qD6LL5KUeu9yZ7pLC4TgTPjzDHWTzpLvLRiTqjZR90waSnpRh
6xWbGWepohyF/nsUJIrtXiYFeILx+oUPAL+/DLcqbKFWq/vLlTV6+qSleBFHm3ek
TSJrkJoHhrSypjFz3h2W54LmeNpxSehYluu5ZRTIRIa4JrN2Lv08suNIBb52c7M3
ZyTMpWBTymVGRwDaAm8UNYiyeZBSgW96nWNlKTbhRUGLHfGLNsxraAi2MhG0oPGX
ByJvvM8JUt/RS60uuKo41rd/RGoiunrWx5nDYHtiHKanRQFFxupBsuILRKgPLuRH
uxucWmCzECbvQr6lnvZZgkIC6T5bkNlQsBDzyDxmIIsdkwR4uVNhPcWpO+nJm0oC
0kivazAQpj8zkbAlHzjc2b68hSLJ1koC6sB/Ru/1gNS0kxG9WGS93O/EBgnzjwGn
3nTEQrN8YEAD89lp2yw489dn7WIdDKuGu1+Kgpy9CUN7YPSkoTbqeGfDhsotbBuK
O3eDqBZvQB2ZanN9KyxeOwJoy2hLlEWSrQGANDarsyTtQC7LxSDwfUJt+UJ7ZLgP
UevMh+68fBpOsNUGkxepPclvP8EqItiLjzKs8uY/OpmHnp4pMVeN5nixgDlJQT+s
9Ij0SqdUuSEIWY0ggs0lxRXMfGvTkhyiQHC4nJn7OTOydKeO1tRdzSKMzOvkfg4u
sfNUCrPkHX/b6M4MAGeTolWHvSBr91xTBIyYxrjuMGpVZ86tqhXu0gv1tF99KiFe
TrePR0EGdxS0AdVTIyIuL284Y3M0hEwWoPAZiNhXdTHDDNvgPSuxMEX2S7+fvLMF
P1GCscL0gsFHsMfIi98j6nRWYD84mdILaCQ8EX7/Uq48k8dhcOOXmGr3z5vq9IkI
hdJcYalBmpS+6MLbT71yDdSmQdxVWDH1BpIThtkle5HKntB9LjrBA5yIo1ea4DA/
ueSvhkaeejr+VOVc/TL8q4RUXTJDA3u/62TZC1NfBdfWo1SUX6eCL4GZzMczMCbG
Q3sbfweUjWvzp9vq3wS+cGV8xmyDqq3CCkZ73sF30/lCaj/EeTcxnnkkFkmHLwHf
rz/Dqf/sKiVXPqL2HqLkDOKrD1Bi0LpXszi8yaW8+0lzKD3aoRCiFM3E4VqzHvca
5sKs1i4TaPZ8cRBsRtsbtAq31Rrug1Sq7f/UJayDnJozIxEpR0dXEdeU4SZ6PN9P
1wezqXqLw4p2yNekVGBJzk10uhtrElVi6Ii6/KvVbBkn8ketJgw9IgKixCsgG77b
GKy03x8PqNqE/s7TSj8/xMPZzoPN9hUipm/zLqd+49rab+BXo8BAh6k/3f5/Wdai
ZQMY2YEaBZBkhdjeSyFEDkh8ltN22eAwnRNJODvPY0fAgiTIXjl3N7BaNkfon1Bq
cNyP2Mz+NkWMDH/nzxr7FTp5iv8TucYFQRSMLDx3QOZQrDurUa9TrRQz9tLsz27u
EVgvJaecBltxT7vGyzNAh/nGUu9DkLuaa4bgI+Gk06UhkaVi9LxG1PnumQKrA61K
xn6VDhqvLm0srcun0evb6pNdu3DIlCtJqYjmt3w74qA2V9yWn+4XKdnvDIxYhB7h
kJme2rJVJtsazC6nrcHrblS8tMZvnmgcwxm2LOEI1kr5W4I07S/F8EZISPLuf0pg
ceEUEYUBrqgnKZQuD1K8XUBvmgS5OBuvx5aF7kgwL+rpMsOU8+w4foCJz2ueVY7/
Mmy7eaqCrrMgo4qbZ4VMqhmZcAxRVMxKf+vwGaBuwQitUr2blBeCkaD1PwrFF7HM
XHWy5qTH1Fo0dHszIICrcaMAx3PvZeY+RPgfNLMtGUNNI5m9/ATSZM8vuoIHWJFE
fUdfIMia6qKZyW24ne2+DrqUh0xKGnH0sO6CVpde+xsDykw0n8yqMDOP+W8HLkXc
ag1SoUcMchaOOqySbByrdwYRqOmyldHY5j0F/Elptff5NKeaWgI5akRY1voTkH/M
LPCi1iW3qeAFEN0CQUetzaA8fP+LOzMuskuUR6Y1Qf+z1fImqZFc4KRARle+HwaY
KSwlfr57UvMtoZQEThOQbAGFlXhMPQgHiM98caLYxyO0mu34kVPC9ok/vPFmRQK8
YKwoXzGITUeYAcxzzK7Lkw6I0JEoA5WXFUu0p+udExr3vSdNjKWkiWIBsNB/9Vm0
BUfysUUZfNoRJBhwYQCMmQI4zj2HdXVLbqPbRT4LA+U1zZoG3saJKGX5RU2dUfLk
HE5KQ2PmBRLcY4DqbgeDX6hUKpxWswzPI4gcJ8AW+pKfrQzE7+J1yDjbmsdGUsX+
tMAEQSUPLCgPmK2RjqLphe1iPVDv+e8EYGXoqeaodcU/NBD1hH59AHDtqg157Y4Z
MvJj1+ysfboXOMu6QwjXr5XIjEZrbC5gzGOkL4DYPcYWvqJBI7GOkmLPGr2QJRFA
uz6IZrGapXGM7Afxjo83TDW0pkjCcHybrFqER/fi8+kwaCzWq4b2ZQO+Gdk063MH
i1sIo0EAVyU7Ut4KJEELZI+EMAPkc4SD+RYHS02BupvyZTulJ4xCS6egQLY//iH+
yEyO1tTc06+x1H59TKYIG1MNzFeuR075C+EcEs27Nc4YkyTAVrZ5K3E53HO7Y/Iw
Js/pyqMT98IQDOLxUES7NrjxP00U06gyW4XGtFWxJQK1HW4vcobHZbWeodcln7kn
NSHeSnFTNkH9eXLSW9riqbd8NnPMOEJDdGHD3V2il7D/8dvERrTiWJtoPjM7fWpE
EeDVGyJoHHQ86O2HDzav7jbvu/IZxuu/zDk4kOTh15I82jGiL6IvOlPdJLrU35rh
k0cWjEcKc/v36T7nvKocZCiqWgMNkjr9twcsfD1x1HVEIDA+vWUpxglqLAwx2rqx
91Wxu/oGKe44kk/T+2qG0wrMh0f0GIDTcGd82A9Na59QxFNyd5M0vzVFle9ytA0H
MrbYtQRvnTrbWBQI/jzDDMX4CORZ5dL7tJy7gAgw90mTYZuXaxNAQcdu8VLWBkbS
IuB1ayoixb/t9ps9PtDAHMAWdmM5zIvD3hgGT9cjnyjWmP4dMJ/VxUyDCWnCzivH
pR94bKjupoVG+lkpr2ApXuAlOaTN5RIfZvByYfKxPSyHd8radOb0nYxDgi9LfMI3
YlxSDdVpimq/6xMyzfxubqiGNy1DKoAoC07MiKkXPNR4XLjWBD1fFdBWxSlFoo8Z
rogZKazgeFJCL1bqlMfelNwcDwZ0bRx2ieEnzYdPMKPPD79sHzB7jxRhSrOSEq3C
HmPtZCA8cyRQRe6HkmTBNLIjheGuBAFTBsRlXQR5AQ5JQwL4kjADNZFroTjxyHUZ
aEqHfbVHnLjtLOxqlMH/iEXZUpjD+EvCX9UKjWh1QR0pLuzaz7MfF+iQSSbcRj9e
PlB0tr8QZn1jHV2m49Pb5URq+1U3iTV1jjowcyPs90vaScEMq0bkfRwoSu+B59ar
oDGKrUtMWq22mebuWCQds3F8BAiptLCl+Sur5a4roBJGAzHtFJt2405dRfrzaC5O
X53lNpnh21APt5m/ERY7/0w0B/WnfbXYcLw/gr5Kwjri2vnM2XHY0CRKL/CowYXi
lvBF+Qd0I43BLHuPPN0kLFHYUcOa4r2sPLYGEwjDbirH77ziumPYHyxSgLk47tzv
HcIl9UiOCh9mWyHGNrkBDMpHeBlbcHb6Hl8692e55zO9HxYqxMu/GnRkBNAlHQ7+
VwHxikr1v5kBfRNP/YwrlSgqTfmyP+QampYEFfjRW2kJAgmwkPIkjuZ3Qm0rUxGx
YP1CbU7cux8S/puXyxXFQ3H8W9TsRNcQyIG8BnVVhnZyREF6fbWgrgutP7QeQUVH
vBN0YyaYAXFV24oZSoBgTNfDLqhQi+xdHAO5kcqQQF0QhkebOtgJQI1Z281wUOiy
SDR3h68UQ+49BjED29eqgpwC1M25qxg5DmEIeGm0UAYdmgSPxQc6NTBEMR+t51d2
V5kjbK87PNd1dOiKafa1RLx3C7RGEb4c+4PKjgvGkINs7D2TyAXiSNOWbHtrRAfd
s3riwyw6Rp5qaoxzQYoNTUPJ5oCm9T46P+704CmwCNV8chihbyXSwKpCUMm8I/qj
Bt/POIp+MhXU5/JKySluqqoX00krQtKGGM9eyLoDYXCkG40bvkXfDI0y5OVpTwU2
w7kRsKOl1azOX5Gvx5Neu4vMoE6aGTOtyZrdL7LS66QouOdNefP466hoP8C7DwMA
6SsxUNDnW+luRIra74TflxK4ppIYDnNbDGwFiLLPbdFk2BLHe46W11xDaQ0YEbfj
ODzGtoJ0/VdZ/zuEj+0FRaLlNi0gWICEPJhH/JuwcT8PWM7J4mIuQIl9xKL8eOCP
z5dZ5pWGv3bE2opPGfYtMSw9qgJuThcKAeGzjdx/aQSDV8Q5cmU1Bnpa7NhyPjyc
lrrghGRPrYSpaQAXE9Wx9cA68cseTj5s5qrm7TPcGGENnEJSi9h8Kt79XMhV09tU
4eii8ZnRVZUvNq5wHeF3s9QHpLjDd2RCcz/Pmw3fOAennq7TxvO02xtwW4Bh272a
4KBRwIDBlCYSupvY8JP9qVwaql/zL+PoMBpeZ7IYxuM51Y0/3VnPPL/KZ6GqKv7L
nW7t9NkZQwQ4qpypOHX98PN6eXYOuOxHb3Q9gDVU7EtD+oQYlv1z7L0oyjIxmZAA
UiIh7T2fgz1gsg1E2npc2kgBNl19is+9Re5CzOQTxEw6FlJDSGBcp7woXdNoPl0s
Zy+89SM9SemsEpdjz0G/7XTh+R1tHaogyrPHdvSfsv6NwvY2MMQwY8pg6znSdoMF
/LWY5eDpdxB9KpOybIiTL2DoUj1EkvssB6Eyr+t6ZOBkmOHpQnJQwHn1keWxLn9C
nWmvW7XIGw9G4AAZr8jIp9ZYAJSMNT9MHNciOkEZDPbeDpVuZZHfG2WC1beEqZ4N
2TiMJfbrBc3Hv5Qn/V2QGQSzEAtx7NoVtoSOQVxSH0OgM6z8Rby+Z7WaWEyxrOfI
AV4x9SN7teqxTrbdg4ADuzjhPVeeKJt8H4uK5Esj83Vl1DxIHR9W5yEtppCbfRkg
o8g2uyEdgtrg92G0BPTsAUdZN6H1EJqOzLGrwuKc25reCtfpwVzdJGZD06SCBJXi
ENq6m7tejETtMEost1lfD8JDmXmMPAkvMBl4NmhxxzOCqrgNFQgMZ6FSH5VZGadr
Y2to9GvwgLErHEAgNLjFu7OpFOAg55gIZZQSkEh7OHpV5S9uLWlhVszAUWw26WlD
2YAJAueKKs/cPyp6aD6OBqY4TOMLsN0YMZWUMsFwht+mvf3N4BxhtRgMP+pEfjjX
LuSMp2KS2h/yxKborJP3mfu9pnNyohaQ9vd0ginOREaC7PcVpJAzCTgvrjj6+yvL
ws8Qh+zvssX22RrPZTvHFNKUDw37sAblmp7xogO6qydb9A76IYf65RhmNeejfAvb
sbHNWz0SAZDrbqaIJsHeauM1UkmOlnK4NEVp0zdg6T4KGNe3Ws1JnBq+Fk/Pg6Pw
Oa0IhRv6THCHnKsjV2OJRyYTsizKhxmLIFCwpYXWVzJ55XINh7MQh5DE2m187wuZ
If82Dr9DDPqmcuoi6QV5uiVm2fQjwArtHgZBYht3EZnuSNVnkq9X7k9YdWZ1DzQx
+MQgHeXhuAn87hCUJr3hlPHIuSvgQeod2lnOHNO2bTguyHmVSXDQuxS/Ty9rGGkR
yhtRQiJxzuzJR+GyLUd8KWNbo9/lZT0tC1UfuHqb2ZwOAafH1OTaKOP5jVtqkIsj
3T4icJ2+8GGuTNEP/KVsn8M4VAjlAJo21vLAsGVGk9wDIpOKy2y/G/ac9t7MObm4
c9o31BrBAWycN0W8c+CgjlkWqrWm9q0PAzZXiy+u2rrPniZ42hMBYCxH/rzcqrRZ
JXE852tScOqkbwZ2mEbyRyoN0FQfR6fURAzISVDXVJuEfOav4uwqTU1I31sryesS
WSzXJ5dBZNeJ8owNOCJ2X1F92AoKKltP/obeZK73AkE675q+sb4PIjp5x+5UTTuW
jrwQA1uANkBwhdNuMxnZo3QTbO6WGqyZGAa/+lSlIwtreu/dt0jsjE7CWr+NXwD1
Hh5IIup7WWgWS96NCgcIhpWXXidxhJqhu0PGCn4MixqZgVawWjUtKebMHdqi5uJz
uD5HXJJ/kTbRtt2qw+O0xV6bjWWPkNhf3iCkFy7Nn0qrRbdG/bqaAgtjtdB5JkCw
mm7MR014faL97panLEBlFLIcKy/5RaLKYAJVNLeT+b/q9m8ySYZZNh7gXRuur8F8
mkObpDL6ludzXXGcrI5awx7ZmiEI08KwW9yFFxPdMKSQ1P2hw8DeBIj2yOwva0nA
st+tvSWwrvuKaefyCL/RlR88CDZ/BH9Q2hjzm9taDmnBQgLVJvMk0BhlHayd+p2n
UGW76tEGHQWzbaLwcTA4Y52qnpZ3WXQNByus/sh5zBmRAAz4KlihB/hZQDTbbowP
U8N+01psshnINL7oNFvwrVMdOxrNyPHhkQaD1J/mmAsAVBpEW053DiQ2mboZSbpf
OEVJ+nDfGJpxuabdtRdDH+pY4lcyddeV1Przul0MxyhtlTxclcRywfaSbPmtJ0LW
kXvh3bqI9ZW/tSPgBZKgpt13EpUYUHW34fRU3smoTsyyUaB4tZtaLrU5yu1l39ex
W6pxonk6nIIl9o4dNhbtpRODG7UA3Ycad8IWANamldr/OKbWmq75SuZ351BMb54Q
j1S7yEPWxpVALgR3TgjYcxdKW7Hd/RA3ETWmAEe5qtQcbVKLoTMQJi9VCPyHFGPA
LKbxjztQAm1h2Gb1ljEFUzYUwpbvdiO0/cnAfCd3ghXTIoelKrRW/DpMezKF5IDy
Q9PvKlyC3/D51/uYEJbTgyeab3fFVhKwuOfAu8jype0RaeRNAqnVXRgcAvsJQs6w
tY+FbDVEB9RQT/nbPL7ZWK4Du90AKbvnpbO97MTMvD3hjF/1a/LlWKxc+kdrKt5A
+ztfiUkQBTiuoyGi1PA9zaPLsd1GjSZHj7cHZUQyBF9LeLS4EgUoF/BxGkCXD5R9
HdilVaiGn+o6cA9rs2APNIEXOYogU3Y2Uvc8jf4fE4EfUytTQe2/LEHDtxNJRz/B
qGrDU2I2kchmUJjCMQJVAWdjZmbjJFLzirrUW8KRZCGsUdxGIYgXAlFNfaiKHIiK
4I3V5gtpHu41Gwtvnm2YV5xqzBgbNE63iztm/iR9gow4gEpm+pbK08Nh6wgr/GSY
XNzHTN2j0g7kF1Suk7ZDDHDpEBkC7Ggqc4Ht4UxB83udOpT2Pk3iM8/wxukuhy9X
mbqZThhMSRLdmWkpV7bUpyy9JO7kYd6DLDLN9pkRoHCCRqGFSH4Lp0zKgDq9J488
D8bM609+nWXI8nO8OesnF+Ntt5BhqN1zlNL/Bep6gbVHzRILKvoJ2TMDOdWMJeMo
dz7fNMOcx0tRNFWoldH7O6uvg65ZE4MotsDFKsiKT9jWqMli6xP+w8SN0LNC1e6+
F4uq8q1tHlUIxXgkdbN41MN24FoEbmSABmm2Ic9JncPnuAudUTM8fYXSdkjw5F26
Q8Y8T2RIczd7/b12rXmQ5kXYqv5eVc8Ce6p0YQXYUD6Ldn3AEX6rPQZtLYiEkT0d
pQROGVtyh5ZOzAOdKcgGS1rgbT8O4kPRUcP1p/LNJvSLIIoXYqH5SdqQjdGMVG+3
VU6/4BNGiK2saAtU5uQuamEjdlBdgPX91uiPkUQEOFYyXtex+rzvGg9S6QSWrLpz
tXYRvCKzwe9OUvN303Qv9iVYcGSw0cuqjkcqvMvbDKkOWg53j4P6H1KuRAd5ctox
VjlK3GRVI6zbQLxS8imOV7+nKqxeYEQRHYMVm2k2PIyt7t9AyH3rjXLmz9YRviWc
8MjgbZ/KiNh7VELfH4Uuj7qIWvIErELwPhI6xIfazL0E0oX2v342+SOkIauSIzkB
zw9W5ZfQMBcOxzyQmpxWNtcP6WlJ0aWq0/Ws4hhrryfAhvK8y4UPuoznnvo7+j7T
Rv2hUn+DJ0NkgBosULwl9Uy6hNg/2N6bELh+IMkICuqnNG/bZ433S/EzqyQ5Tcha
8dQtx8PliWDfLF8raFrdjqeQJZ1Z5vScEm9xFLnJLTdKJNg9pT+vSeaaXSKvNood
B9ZPO+XhIUAO63hh11RbpN3DwtjIGh8d42ArCdkXaq3MoCzGsu2A9rIdWqM3gWH6
tJf7WukqI1YPf07NdBJrnFJpPjyCay8QGgAcFi77ofwkOSQqzPGx4bgnq7el6wWi
Fs0tT/BzrwnG1gGXrdRPzLvaE6XJtpOUe+sdDpdyC4UV6rFSu27EX2p1esivu7rN
Q3qlFRlZSHcMIe3c9wTZyqEhPji5s4hToY2CPaXnAZeA4L2f5LRomEI4T3OyYbXx
P95/KPerXkYKiTu6zh59I79Hb8v6c4O0/s6jNDEc0bavQiTRYZ8aw81iSMciFsdU
6nDzKc6IPUontUMRN4i5kEbirqWLgYUX01HmWKReLp5xMhwjB5mujvKYUgLEvWFq
T6WgeSEskDS/nA6cBXZm4uGZvSPf5Z+DFrvlflM9Zzw0N/RsJObJ+H2gEnGaiYWd
JD7JCH9Sj/b5I0osA4iip1F4paGE0EVCN4bOjbf7zCOCiU007esFB50dKN3HN+uT
RHQo6l+PopORgz+CqIHBrgQ3WcAwergc79nrMvGUD3yyw9dceVjbAVpk7xpHjsMT
EHFTJ1NDJDMl6Pj3OjzaxAkBIN/ggfZtzv5NIR8e/3I2NFgTTKFseIvRZlNCsWZJ
RDrLAFri+5GGpb/S139cTkkk1L19dtZLEFacEBmv52siF7Nzanf5tDwoQ63gw/4o
zalpqFzo/rRAhhLw1vZfSJDAI52yDbx0wpJ9y2QTPw+gMVtCDa4eUn5ue0PS66Zk
GqCUch0G4L4KKw4KqKyDRaU0zcP8DGbVRDcuH60tPhfF0M4x0zyeATkjlMt+1Xoy
GhlzY1A6OQ0OuCC4JZ7+9sIJKL3GDHPh+ihDejzkTznDzTWl/wewdpkuZUwOOzWd
W9+C1hOw/xJH3UFp5l3G14nVzmjgivDBSgWp/XYs4Ruym1rvet9ymVTSPw4gAY5x
pt2tuEmWFRkCYhVVDDyHgB1RVI5qxtOIo9Hbn9BikLPmg9JcuBWTZlalg69g+hiA
vBw4Msv7ALWWS7J4/XFpoB9Sg1i9LyvR4igpyhsg/6SUalPua7zRbc4dfcMkte6G
Itn7wSCvXK9/uwHEY3uAOC9RiZ1P+uR2ssbaNBewszbMnZAJX84lBwk1U+nBiQDn
5CTWlY40T32PkjsLKdqLzpddsr4TVQ0USkO+8v1S+HQKSTplsZySiR0cWsfHomSj
DHI1+odrN7A0rkRMrJMh0uKWPa630BxCjFbONo+MG86NOI0Z3SUGpa32PMyf79WN
gOPsfiiYlH9TJV6Z27sxIo73B8TY5y8apX5taIiEZ1sAFVmvrJ/E2L3qzk5VmoIB
wcMHqAygKOid7ctb9pKlqKGMWMQ5KQfG8d8UY8DJJ/0nPgnBOv3B3U5uHNsvaGp8
6QwTy+hP3QaKmX22b2WEDYyMxwrzwkRdZWq9sm+DU6XXXFWaHyGuYg4+uGTW1wgb
c5WcT7BPl131SAlXtJqQ9lDq3tkSggoF+YwIDQS5mEB40Gu/RRPgi61zoWxEEgWt
ceBYnRIfXGw7wzTTmcCw/wznhIVvlvI/BcAtVRuOCFxH5QqHKV0dBulqa7yZJ5tA
A8WJVD2JE6ljoXP4K1fALTxj28Gk8K5n33Iu7f/cN5ze64++KXpVhbqunjbhTnzl
Jegeo032uvIc9Xzy8J96WbT/QcOaqMmA5HCQbcsaOVChO9GyAYpTXT5iQ5cYWC9h
2RdgRx1oRH9xAn98TZpzvpd/jQaSzXP4RydRwO5ihGYxh6lA+OIho6R6exXUdOab
ARkOw68sYp5L0jXyANbOQAnAGSEdAIQblQr+trjvm8wXKwrLj7itX4ic8jCTZSQp
it95X44EGlbECkfUPJCfnEDOW024jQ6Y+q5Om8Dv4CP1hWqaByRth3kBIrMkmt+N
WhSvQy5K5I85993hmx4PxgvI0xLgYaxkSgfXUkkTthHnZv29aVCqYHU2EZkWz6aQ
q080L90OyNSCORahhGjvPlme4OmiqfZhKn5PHWtFVu5AMnQ1Mwrb21vwbw2Fo93K
sE7evubUN3pCg69V/4KoKWRlvhzcm10EsInjBEiKCbU/9DTVZtBVJgjzxE8YPyf/
g+Vl0l5Qf88CuTAxEHZ26f7+Tg43vozjePjqs51XOL14k61qX+5xozfnV1jY1J5W
uXkseuqxmd1CKFX4244QGypmwqlQCM4wuep/NmtnqET5ZrgoQUpgyrsuIRcvvPAC
bCNkHTjo1+Do6Y/L+fLGZqHTuhlctiBGNO7aNRggKrVfQFOCBa6TGMOCHW3cv2nO
5753y1HHXZTPdBnkIDH/f/8bQeVwL9sYFIUaGZFq8SAv6sGPs02ZMc6Yu72qH9yx
/QBHrzd96RPRtoBdZK/j+cHiDE9w4kfWksvBG3MOCDmmmCQ9Z56I9YZy8/2QMIYK
qwNyCFoccGpOVxHmkcQcBTc59xAZkZiqSHIjsu4RgbPbYfHrPB4v0SPNLIeLAYfH
WzSBEpI/pZfM3TEeAMRcRmGrZEnA2DWWZXcaMIPLL9kP3WMWr87mDqeTSC8Ip5YT
l4Of4ik4zMQ6/3V9tFyM5IglEG0l3DerRG733arW18DaIMg5UQKV/RZib4UbOvKc
/jHpv4NeGi+HY43k2n8Mvqxy8IK97ZMi5J25xgJvbMBKYTPDeCb9TTJKKZ/Uwamf
dyvhH+rw1HCOsVNKuyY89YtE2I4RrhHMv3Taid9XuVkGAe4C69H6vfGYGgbCjRFi
eMvbpRk2YQuysF7fSvS3zpxBgtgDO59EogN1ysLnUUbGDeS6Lo5fr+GFCFg4nCfd
MeeMfsoi5+7wrVY1XLOvqLaQ6j8ZbHotfTVU3k4MCrblCIQf04uZ4ZosQPiPdvah
f6GLXC2jDrAmW0yJ6DsAKt1psISpopVIKolS+kr1m+Wufb8VWiXLOWBqcZEuMu1E
GRRI3iUaR8wWleynkhBk4GHNu3Cu4Z807Ptai8rm00gJtoXzR7DqUXCpxTiwdn2R
ki/L5uNOKSxWpmj0sPhyD3REGmAoQuxVYiodbF371e5VV+pY/VUqWjSUit0oqIxR
qCWaSe6CLjdHNqzOS9CYY4nz7lOe5q/6Qr7vNB8X7zoHEI5dNrYnQa/IgZq7Z/9m
eLhI2kuv6S7CP60irpKISi2IwpN8WW/bxeZBlcPgYamZNcNReuZV7PUyTASn94+j
wtg1BaH+8Ah33FnjlJ3F8rHCMaUPnnxAMmI3u7DpAOawFvTYTWtd0xNYj+eiOQTZ
PpOf261WkNo7Vvz/hzEjOU+oXjtszzfgb+aJjjSB+z0n5bg5zgapdJEYmX5bAhuC
hTZ4AFt4NE3z6vBIJhNuLHoVj+Q8jau/uYQBJIHNk09Xs8Tg9pWwiLGg5eWcRT6r
v5YWefRmsYOLOI5U/l8mNq/OQkuihimmD/mFhnvzFZLK0MwtKnnjIrQUaJJOvKNc
bhiQDI0APKrZuU1TZ4LGANMZilJoXHyzM9iXtsp/TOAMm/57ht2HWEWRMm5NqMHK
xIpZT094XDUt3fes9ZK85RzxMc7Kv7jxjpgnOox3mx+Xq9rlEaR7RwY62pbvJDDz
xqhF1BWvtVEbW2ewZxQ5OXrsvklpTE+Xc+aDmOrLIuu1xKJMjRyRaTGs/IohwFhY
8xSxh6mv1KELjW/fCpDORH1D7iNL/wgfU8RJKW5X8xRDo0FjoIRySNI16v3/K3Tw
85DZj8Iverwbtzru1LTQ9XJBWKd2kpO7hK7vnwc0c+lEIJCZvXVuIhrTYnZXRaa+
thEnzvbiNyp+HtMPi35GjwVQ1aqzvH3OHxpiwB6NJqMafyn9Dv+g1jJLSMmDWnTj
0oyj8DzkEM+BE3iomJlc87+IKHcn81z8exX/q1fYMtLfu4kAyJrHxuM2E47yo6Jh
KjpZFKIQ3eSZ6WL0t4SS8xNi1/qX1PcMEp3VPSiocBbW4CAuxv2vrgbdtxJ5O+XG
19nxkyuhJzTz2IUx2nsoo+IMV2NS94itR4piyZLvn6U7FUsOY/WaYUV6jriMo9yA
m0objMRPL0ZGK4eRiE4wu4mC9mUKA/ryyNx6GdBGJnNZQ/jxPX11n2CMn9FBf3Pm
az14cAZykL8AAmNqvz3aVByVtf+0i8+LymF+s+9vcrOxoTWXUdsRbAewzioX9ymL
GOAJUUADz8IO0QrZtBjjnl9ONaZC02YeZEwjlZcVJuV3ZYrTjpyAgF/viqKUbvKV
jYQvAFacKsgLHIDer8AsiteecsX7e0ciaCkc44zDPKnLfuDFcBlOVr6+5D6szdem
uvR6suv3ROo10yOqPaoxqeG7/9qkMvfvMSO6e1FsyCktJGVAu6VtBkbaeoe9hUFU
JIZbCCnpbKnPHfVTPOjNJZek3WG3nl5rYVJi4tZFlm+gVrcNEJdmeDW8dhZ+oJWe
X6xsy4PUtpldLXlztX/tcZHyT4d/cVwlqHePFK6EGd6u7PaMQA5S54emwkqTmyPa
HqbDATIza5sBV6lAN9lMTvNpFnyP/CkcJj9hLPiYOIoX1PiQ94A8FM5/4Dp9VBhg
NKnaqVDi8DmS6d+CY01NCiuf4ZmV/YoGvsop+593HPiwJUeteugvcx1lDUh7AyD4
xg4a+mCP5pg9+HaZOG7qV9gaY6h5hl9xOIsjh30hRm8+gwypSaA+D8uYhl+1wfIf
0ELFxw9CEOUqfLmEzc9Q/tbiNr94/MYt+7Z3kroLgCa3HxEheQ5TOLBt08oPIMxQ
rTRLsYmVDqqUNUPZJ4krmGXx1+9Fzxcpnt9PQPYn90Ta0Mb990O1MLwb3WZu7q95
ZSjPapMSOALQxOnn5o5SP49UJ1nq9IVlBwXMJhJmqW6gaCL9LvFyeoCd0zrgS+nA
hNCpkdNE77XIVsKbMum2jcWHvJIGHP5rbVUP7C3ylY7RBYU6y4xnhD3RpkbjSFnP
B75s4tH1PorKKobptG1P6pXBqecwPldlWC43rOPtX9RlNGec7akD9vZqSl5TCnZ1
6cqN2R2r+1c/pPlrx+YsSFB8A+jOmkFmUPjHQBfRZPTyvjgUwHC4sJeaw34LYMAr
VnIaxgiUcifQ82C7jPldm3ihT3mskZV/ZwsALJZVUVGuVh5NN81d2ftfTuzjbH5Q
7WU7dqjS6FKmvqrAGVtttS4LUsGgMtFznnGILhx4UBziwYXiBXXALygqTpb1GilE
uQ55Mg6vlHACkJVjnHYZaHEOObYM2ow0V0p4+i4XiHn46r0CCX28IUpkkA/zfAXM
yq59Hc3gTqc2LEanySPREIzk0MZ5csXqhPtHUNkaRJWOpJplFq3CBMcXx0EAPAjq
4DR+n9qUYr5KsSajyGzjA7jNIl2pTYDiwzzqK9mL34UK9y5nTEc7rxl7fcJlP5NM
a4CPu9TPsNaguCALo4Og/21Nhxtn1krHLO+Bkt/OkhjxLJJPvaEllv9NTQ8DJ7u+
mzb08I8hSOyCi5nyYh+iOyUXJ66SD0oMYushfffqVx+SGrqOgdEIX0KLv77XX/Um
mk7cKQ1Vw0labhac3nCw1aXQvBAyGs5C886O/hbew/dVc9hE+JqgLzOb26H0ZXdj
YAfizTh9h8RF43SDWIB8/5p9KxVi6FzvUBw+da+SXtcNC6itKdCWG7TqnmET61JA
hpnCvwNV3I/LzLOMIvrxWSr24xwI9bW7/R99Y+meUuGZq7VAqRDGHBkQkuW4ck3a
s15FiONKOvT7kloX8Z9b2Cqb1I7m1NWP9lOQxwgY8WPr5+mcsqfKxiTkFssyCLes
CSiG/zxIA20ZOgqFGIjA3B58FWgwhzf+/G+2TvueNxphzEOebXAmll0YgqnXaviu
wxZMZI3qZL0IOHuTVGTWmOCK4J34kT/etSyK+l8ccHJFR9E2kXUNjXwQyEtY13Fo
2vIbZ1EqiFlXdNN7aGxK+xDoj6pv5WSxo0I7NdHjMZcIaXc12K5ft4PNMaJaTdlf
z0sjDFBX+WiNE0zu+EEQPBTkcZVtO15AsK2qtcwY31B8PqxvTHjKzPAmwQ/ceSXF
MrS2plmBLoEj+FRdpM+lPBZc4lrIvYKsruNCWgsCWKsnHzYpIKZiy5X15y6y+pdw
9h8k/nw6YhjjzYzrlDaNT46IiNX3T+He6EsMz1dDuGEd82JksNDmk52zLcjz84m9
u1FpfW3qzuDRRo1+Kln8bn++iP1uZOH2Qp7PCIFOmVNpr2trCqlouwvLBKiDBa75
QbL43opDP73U4AvqIHxZ7qE/js3YKYxKhm7F8QeK0NQy+/2WQTyOzXd7vABC6TkP
mAHYJX3Y6vLOuXw1knUKw4gTCDuk0NzCAQ9eg2/SlaU+rEBS3vDNpjtD+G3eDEZX
zk3shS8XjBFnUHfu8Vk6fH6G54aNKe9+hh8Z2yx3GfffxT0V2VtnDDVRL8Ktjd5z
d4U2DHQb2YRPYnPLXSN8bb0Q2j787vxyuSq4RBX1zUC8J29evy5kEOxK+aGnnywR
PoBrOoNcF7sXCAOV+fxaW1WewhYEDNfImyjvcZfCf3nJjVI21QkvNxlhw2Rc3rxi
Msp+qWIKVRdn9gnGf6BGNYFbt0RVCIOp8shZcUqdnfe4rNB93fLucyigQxT9rgMU
ultbHT7jzsOoQDAJYTo6T8zzzen6W1TKDzV2PYExWijuyLYvQs5hTNuKKSW/ytWW
TOIW4ikaOASk2BO0YsZN1Z4PSb4oMAjUYO2D+De6kSePSBJDJiN/98Z4F3+qdrdX
kqKGF4IXtfK1pvxNM8DxYPaOOEiIivHAJBx0wW80ujXroKmMxzMAeL8fwGFR1OIx
8bMS4Ux9nTXtfoyKBJnDTXhP5x0Cu4R0rWwFKFNVQxt7wWKnkKvxP3wXwYtHudPF
CkVYxcRM/Y+visFiglTECjPPBAWH4LqEwM8ROlHu2buKwqfrL9gwUSB7aH4krcKZ
R9dkaDs4UPFH78XBsOW+eW1THqrDSyRqnANhwugwpoOg39lMhF7UX4fgVaoix0L/
WR923K3Kw6CohhSILnI1RR45+YnAZJkctaDJY1E5oy7sFWMEU4VMNHKd9SKHd1Tg
r9c4JaLEQu1XRBKOS/BYi2H8zmcEv81Xd4DZgGPbvbZTIZ6Y22OZfOj3x07ItN0W
hpqRaVag9w3ErY5U697t9LLbhU64sPwvcb6nCnClxCazb//jjqtF3Ft4kGfGW+XN
vD0t1tEWRM0ZaFA+FJ06b6QLLJHBOlsRdrXepx5DjKBmIQE6GxUaiuNB2ivNGigk
v9S0ty5E4RDqIfykS0XtxpMMeWpE1aCnfflU+jDERuv1dwYjjKVJ85sgvLoAgU8e
RFFbfdgc8DQ64uq7ZVTBam+mhFDsQhh/3FsJQxTfpN+4UVV1OU2rr4KKNQ6DUuwj
uIE63kcyf7y+/z2CDPhyGAfTUO6+fpCiwBP+OpRWBNPZMubjnzoqpdNMbDA2rdmC
DrIWkny3phgLwldw2BxKXbtSOXsMM191zGlZ38f+6xvzBi5zc0dh6KfSTnFFTF+f
Xx9OTALCGhv1tpLrMj22bGDsNaWmK1KhIaFIccG/g0Tyr1WFPHgvqkM0dknkdCK8
zwWM0odrKWThTaL2Qb94kEXQ/eFNbTBRJp+hnXGV9SlURd7+7iZRNfm/hcRADh2a
i/dAevgBizzJKKrecJmKLivuOgdp8wy5qVRpOuYGQLYgpA856Bg9xVGkR2pSYGo+
4JkvbdS7Gu4oFFZ5oFSmSZ/ZHoAF1uOUpmj3D6boS+6RZPcpdLrZwmDLnyqwuTSu
Ks4V2I9Bq9O+cd7ZiKwrehxp8iIVnFwSrMp8lgIgQqgSdlo7gTryV+AfBJADRlcb
THRXwZMrkA92O/6BqBFM/cjykk5tdpltCIMn7Uj16yS6PYGv6NLhVZCEYb6hyIQ1
ZmekaoHU9weiaOvnTrsdfDYg5532wqi6broGT9aSSb0lWtqdXwEzNtqaTN9Scl+i
UZFChY/BZZqQkZMolynPl2Duu5r04BauXtyEkiplZC+AcwxHGiH0BfgaF78y6l+i
aH3hj/U31oDSUnP3xWXuyVNW6uuSWQL65Xz8/j9CMryknh1TjZZfM5rB6UdA/iwo
ZUOzbDddbLIofiKdApyj6jBEJX1mKylbZn+hs0xwMAcMxkq94DX3FOzMDED9Mnqg
nUWMKWeQj54bEo+MtImrgoJAC4kvqBusADJop2PCAHN0+zU/z28tlPdmtOwSZNAp
8Wzf4Ee5X1DQp3FbeKnowYrJRWGfR8nFL/dh9dW553/5yLXmFzwTfmMUHyTI+mSc
zdAQwy4q8Ur07moZlx3/77EvQnxJdi2oBbmltvSAbShgmPJn8j2wlIbtxiJuIDaH
arKeYlgT33PHcvbpX1rcbEpytHFr7rrE3Nb3RTPyveCseTDlqU7uatKubj5jP3i4
rhfeRcjEFI3BA67a2fFJ1d+g4/J4IjB2NHh8VfaZjL1ShSrqnKuXRI8+Q2SKrtWP
SM/flbeTiZFQ4/cVaMFGycN+R+BDiFoSMIGMkWNN0L5nMKBOMGr8YV+l26ok4Xbs
PFFFuSOdATGaG0Kf31GPCQbC+zlNj4T16i23/cb9otu8vnZBS8ATUkfX/sqokP6O
YJNpFG3qprebzUITkdPtN0CZWxXNe1VszKJMggqaL6ATe6EY1CDs7r6ilLQ12x1l
MyZbPV40R1tmQ4ogpwl4kLQLRExdWIVPCIWFKRkfBl32kfA+ljmMYzwcVnLDJaXm
3bJ+c/3njqu+z8Pjp8zKSdg8wc3X5XmoDjLNw5wcSVMFXmqmEKgUn6prtYni6t3o
CFE6+IO4lZrK5/QNUg2wrE5J+GOAnQLcNMayKtQdqahYUP/OcsuYbWnedBSCX8eb
ilGtAV0wxJY+T2NMw4GUxLZbNuE5ZQpiJr/g9S3eNCWEMNTdmby74Htx8uAwNRRM
/zuYUkGLc3ddNsrFAYyYJG0segd4mvyF9adTns1IT71sL741HOav/WmHWKaz4TBi
9W2F+z4Oknv/Poiqc8AW1jxJNlUszWioIBN0HsOLIPL2yUeHxZe4nOflvmrvrWhQ
1aOaYkE2VnaPtCwVlqDL0+va0P4vMxfUxloiQ9C3L7Kfgq81aFLqkK+TYD3ovP3I
6CQviem30RK6qmT2I7lpTOm/8wfK9Hmbr2Gec8SHJI2SLA3kX6d8KEr+CHwJ75Mg
Q0nFTe3ps+f0X+7Th+Nznnw7NLDqfhA7E6OGCPG2UCh2qMc7a11yBCmDq2yFEffY
6SeLYEkjqSLW7bff2pZdeEFNfDYy/mlSTAZtA5U0C9ZFVmYUKkTMQI8WWvZ2Karz
6UdflU821oVtjIALZE3hIJ+lkpJ6xRJqxGgVAE1pyRE0DPzS6767hfeOPNxTZNBZ
bn1c0M+1MFmGwgr3U176T0TSY8zJNSc3H9ovtLAiNXXa68iUFxkZ4ojZdG5bsn8s
dwmP1ihtiB5mIyRu+/p80MCt2XQT4DBwabUqUA8n+asQjkWIUDd9xkwMnJG8DNoc
KzjjOeyLT5tpV6fss7Pr7SfVUkbPabLL+szWTwIswClh/ZgEgQFkZw4/UEklw3XL
gFnJWzOTb2M2tqhnXQq3OMt2C0RpA3axEMMkxt2mqUsOFlIc2x23pCXHMs2nHQj9
RaERW5/KaCbl53nv+WfEu9ZNGvw8ysohA6uR6/ksX4dl0j/+4/dq/Agox01xWpim
4P5zBUqcuHUWoDmU+rMSuxdsAzOSON0YPcLlRNV1FCYB6gZ+HvuP1Or6G02Bpw0v
jF9o77QRkw0hk4mB5hCR0pDW9awpjQEjKhGjh1YWviXa741mlLPyj3OH6f88kezK
C4hYSly6r0RqY3v768+kejz0q/CW+Cn7hGPzfoQsxWfQW1PrWLMsvWRaJiacoTEY
W0K00P2N5oPeRsB7qIYAssWl/29vnTSAa6G4X7efiLRgHs/4NEWHsuiTsYJGMXCz
rNEJgFp6X0dkv0MrgRmla53OJwtVTT/PdP28EHMB6aZg4P3occ4RgcywZvuzdtoo
mxKpjNHkvg4u/iRMHMTAtS+ifcDcM/06bkh4FHbEmRlETamnDRYzbi+yI/A+YJzo
j8kmzBpW+Dl1b2yAf3/wnOQ18j5ZYE6zlD+CGEnGmLzweCU62xRsY0NaoGtuDYvm
Bs7WFE0JjuWMMs0NsfeJbS5liB687f6XE5jpD3AVcvdwRLqabIzpoQL54/OV94L0
Rv7P/oeMTWSDBWu9TGcRH2zMDTR/qdZBS1J4kBks5goLyNXQvKnWK28npnc9oYqu
chC8Msi3KMAok3Pljw277SP30QkHcIH3bdBY6L5N8cGNzPVBuWCoGM45TiFeWyGN
xp9Qj9tdiOH3H4zgIteeaCY1yONcKk0NB0NduUsExeNa6YYeBsuyC9ohw255o2t5
zKNxbRN4CnMBfSCb5L6wknhHgm+iVg8kQ1Yrq4vsL2SLQ8wwybpCHshYYi6S42Ym
Nw1mimC3mxzFeJ+Dur+0652p3g7nA7DkaeS4DY99XvQHKnLZPsG95UBC39bUzoza
w7woOOld5YAbyCz2fHUKV2z0vMjpE2CQFkSkrc+Is4urZ1W3uUtbz/ujjUMsVyeC
mrQJXtbilxTqq017M0VCnVtbG0h6HkfnAv6qEV39amAa9Nkqm6Xmdjgs6+JfaP8p
aLB/BUCzM4vVFga06djRkY3PKIm3eL51K3Bbq7LaeJIowwDRax7qRnt7Z0GP0u/o
IPeusv5fXeiWwYXchrmL0jXUD0tcDDnxdrhEaIZARYy51OTXmn5ZGsQ9Z+f7ZabC
I8DMG5kU5w8mwHi1/crOG38tRD65lAQWoypLVDAXxZEDHxUIiEwIW6d8p2NlkjbZ
EUodZ427UuIg504Zs6rUPgT3SAz/NP3XIwB5YZE9bLsS//taoTSo1CJ7mfqFRHyU
lHrp+4SwzuCu1/goARPn9D+/Ki53ku6JcJMW9Up8qv/vGbfoIA8noMdi/LNFqIs9
yOG2cylmQ8rz/49oiMnXIu7XAe+N7eNCsrL/tuOzG6DQGkMiaROuO+60Mzz434JQ
RedKWMwBq6AQBn+NvgHbufh2p2Lhyu4qHm+KH8FrfKDLGpgiOfkfZXcfc1Jb2/oB
7vZ7wqEdbKyO4rQXFcfs1FmWpEv4O3QHZyxxt/02HBakzqcCY1DSREf2Zg4s0iII
PkLi7mM7iiWIEc0vhwGtQwVKI9dV00c8n25WWw19szbQRg4QwBPJkSzHPSwqz9M5
vjgCOpIglfHfVZvONCwJbk9Pev+b9/GisaGhmRKn6xLWWPqWEtBpWkjHPYL3XWPF
v/jMLhrW2xAdntAmyPmUf3xwbFDuHUWJmiUSd26OFvJCicL2tzLj8XjLN0OuqGCb
6V2RAZ6HxG4mlODTeC2cuuVFHjd/WOAD0IvE0gSFRySWg/LvrxEC+NVABUNTUuT7
mfjKbZGoec5HzQkothorIU2UkDQqkmh/0H8ZM60GjwpeRm6NFuGN9oopMZ61HbZZ
LTiF9JcQr8j7DZeL3ou/tNyZVmy5EwCWnG/kuI5dv+/k5HhvCyE84SL5O2vj2uaF
Kr2H2Nk0kgm+oQIF/lsge4HoJWxlYbu4mlM1FmrjzG67QKpPLNddRIdc2P21CagE
fkvMjSEbmccfGRgCEH7zwGuGChbzSQzKh5xOjS72dlFkoiCecaNNCmhgk7q+M3w1
zeD2hKvIvbRoWw7XZPpTrBVfmHv4O1L5dD2pXfETowDfb/vh7CC0phpmgabdRN7Y
ZRSB4zanwNxvdRkcoApEyPffXHf9de4FdFCzmDTFDKDwsQnRSy3ptA8yL0z26KHm
v3ZK3NEdEfILRhOsRXp/HCzwZgxJbQ91/V3uVe3HR6I=
`pragma protect end_protected
