// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OBcxoV+3ZiZZYnO4xTOBsBXnf+Taon63EijvOY/Dl9hzgZqHvmTGz4vtYKtoWd0t
tDNMrKv6QG43r1Vd16mL9pbjZr0WihoBZfCQTyBqiGulFeNhMS5wOVnIFgbN8iYE
oXPuvV2VAIP4GdsSJ9+8txJBN+1BjLPYNr+EDQkPRcI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31024)
BwNasXbTEpMmMIdfBCIOyF7EsrY8oWJMfLULPbHH5ogUKif1syK0pIut9LPuYjT5
HvQyi376VGiAoge7q41LZcDD95fn9rv73Hh//bVnltSHvBkXH97iiSGJkKU6BkwV
QO4ogpX4HH0QymPpyEUCtzXo4Mfxz1agSdoIUlvreXZ4DULTRv7KtWq3ylcdGQaP
JeDUOKlIg2Sxh5xXf5T9szTw/iUnObwMwSjdtkGNDmjFLKT9/SPDLEBS2M/8XPX5
xZaVD+SOLnifxxzi9tUfLASJ7MC3+jU+vUj2+mHFjGWqoM67NY9zqOZUS+k9ee45
0zVCEDwl7+U99+XI00U8DLVYpmCa01CG8lsZoq385/sgRkBhvFSMwDv2PL0/n71I
Sm4b2Ku/RDHftfCGpICYRK4FaHPEQ0l15jvq6OAjahKHBFdxJKhZHMMYOgjWriGL
EGy8KD48Hm8jWnTxUtMbH3719j/FGSKu+ozOc82TyaN+mCt5nxsrLvqxOEjWYbO+
7H3ZDyE1GV78b0KYJeDcwKrRxTZIqf86cFRxn1/pKhV6XQUpvFOJWvq1VhegombC
3E9Hy0k6VdSOXYDBLUWHUxYr2SrPEIxmL8F5sDtEcm7TCO1rGTkiyMd3pmyLa4pO
T6ZKM9pdKcD8d1xkd9CACjAF3mSRerTivdfpc4iiC4zJ3Z7zeXw6E5RWfiz6NY4a
IAbFN1QHrnBvvT1IwSjlkLFMSdkH9xd0SFHQ2F6pQdCP2t57k9wNftYSf4TwhyIi
33NCSMX4J+BCfrBREfXLrgjIbgxeDflf98eS5BK2nkjg6npwsqM56UBAWvgskXlq
4PfhVZSPNSRwDndBqSePBs7gDTspBZ1w2ZPadyOmEJz3t4yNJZIHh7yX6eRlSpEE
EK9L/57HAHkZk35sP4Hw8IKo8FWoYvMAc64lv9VKW54Q54WPKXIxSKJlVJNrv71x
FXz7rbZujHePJRJrmwHeuISQPQiFQICEyHiBydAnkYH9bzNGnbH6Jp3ub3FwgEIR
XWRCiOu0IDZgjDZbsC15zZ5aIFTO7+LS6mOkoMrOZ5wLiu6TNZhxgnwjSQM70n3O
6xuZ4IDL1k39TCz/EWDiijGP1u4bASTnN3fMlP24WD93maZUrUPt38F0vd7KnOoj
lUKl6BQ926Q4B8L+cx1P7S6P+yi6TzMduiM6xuL6fxpO6vCCLaOVzCOmRtGz/UbG
S9P6H3/xc8iPQHJ9K0FMduPKYPQm08HJUst+OcH8Q0SF1Uj2c0Fj+5aP0OewS5X8
RZEc994wtfhwvpr/9U94ZMGi13zwEEzLjEkCBE2liNKQStA6Ze06lJxwzATYYm/g
trmmFtHB00r1j5JkUJ9YWXHjEPDIvySo63YvZLST6TG43F2Fq/dKwaNOcnxBmLrf
YXHelslBlSfQwLaqr2zANf/EXcKx/5zGdHVt7nrvMMVjUeJH4oi6qOgRRM1JExxI
zQ37pH/kzRdP2J2hnoQsmDcBobOLYHp4geONRKomVYLdOnhxqXYKzLpGaKEZxY8J
eij1Hlub1tDjl9p/0MfRa35cEwavlPZCXqbJSw7TqeeqZ+SueX+nMSC2u1a096r3
AeWckhk8x7UrBPvEIWwf9NM8EdTlNlxtQI1J0z0+0nN6OtsBQ28eQSLeO9Kn1wpN
dwGcLYPdiAkB/Cvb2/pMx9CSViNNXxoPaHD4kpBaxFhUY8/VbtIvIz+9IyKtUi8N
yYamCKx0aetxi9uSzqMaXaoxr3wa2M3+ZY6qjej8JyWWobpq9XM9b70LLo9P6F3/
RGgdHUVn39mKNfueGiscmDDaI5dA3wnDFDYKTgIFglk/wKEUYkPiBfyk4ecHx+K4
CyjIgUbP7U22UxwJc5n4Nf66lpcqlAV1EUFVJKLEYLkttlm1rRT9L0OLtVzb7gsN
/BIN9BnH4B4Mi72eGBEQq+s1K0+iX9NWAD7nhYC2Ybn8at+gmIT6nd6t7XpPdcRf
q32vcr1HPaZ40whuY4vJxeCAGpZMS2NHfI0ft1BJ5NfheDd36VvR9hSTrip8pmI3
agf2hBjTT/BVG5Fx5DY1ntVr7JzYWe7zlQ/9sTuaCGRX9ukt+5/leiLrvmhgp8do
ouNiCkV8gn/2c/NF2tMGQkfRBWFt/9VYOkh5+NNLT8X8tz7jDgHWmGp2rIt9sZEw
29y/s/SmhYL0tWs4wUNXhPIzOdW8m1vnSyxUD6sZ29bM/mNzLVEaB0FiM1ThiCP1
wXDGyfgmAq0QoNPhDb4UttQyjtEldoj81JupzR/OoSrXy4pe9WICyxDzUhQ+B2UN
MHYEnAmh6hRiOKaHusmHPWLoG7kPoad8iwCTJe8y771fTl6xeM8Npj1LagcU/zxl
ZC54AUVP9bJyczPHMskWe9UjcPNn/iZWlJeJ7uSuytU1AaQ/puMdNvV6GoRoI/0P
skszp1RMoTzEMCippJ5ZwOsGLt87jNbnh3xZt5d2h4QRX9FGVCHPJLuNwUzMbOG7
g7sY2qJwpkGObDiVVZDd9a3OOQqH50eGR7s45jsggLHosE0eQr4ezLDhcysFJ770
U59aYg8WAVFi75vS9lTAvp6+YX3KtwRoUo8t/xQhYwG8zDi6eQDVcyx13nvS9tgj
q8C26aSQxWTIE3147E4nyQWzK+4GQCkC3KhN/toi8qT7TAnhSyyFDy19eTBaAu6C
mZukK9Gbr3qVZIm/eg0Auaq/zcKnTf1jZPPf5rS3gfcgezYqfsBLJUqe2ETMZqaR
fQkiGpKULPKFzb/F8DCelbP1NVoHWxO8kU5cEitLa/302IrqsaBZVr1JllSqM+Wq
JHL08j+EI86uFO/AeHaGnlwogblehcli8H8t7Bt9Ph8etJY0YOtKbnoPlXilwJDt
2mUJfK1abt8e8QiER5vEFpA6N0aTd/KqzTZD2mBqsV5hg+2VfjdbUTKvU585atWQ
BA+Xv8FwArPhNut1ykHsdAQeZrrTHEy0dFY7tfIVMsGQhVc8QFav/b/zj31kPxqy
V8IFkApqS/acLJugYr3qDqURovqcFE5QFNrnUCQI4R50V7/K7nYOFX+9tlRwKzDu
L3jsfCqwTzieCy7adR9DaGn2WLe5UCfqxuB+Pj4SHpBYYQe6sIzUuB2TNF4O2fcq
VdL5PrTy8rHWL3bWmu1/2yzFogjl7yrHs/If2UrG2aMUf9vV93zkMrwBIS4YSVc2
Kj6mydgobZteDDl/Vo8IkQKAz/c06HZPXFIk83JZRY2ZzRbRy+B/eo3QIwR5JM+K
VFBdUn+RMVfm/q2CDdthyKjHeV4EzJvsxlwKdi0kNr68zDP3jK8iIlukBrzlkt+v
tyiDfCAC8/JlpaLnrsKThwc3NYzNX0PmsNlbLI4aXZ8Mb2kPLQJh/P2Fe6oKeVDD
xdTM18Cp5maCkqO2I6zlAjEGoFvN+xtUp3aJX5PdGpQRJs95878me30LKrox2fr0
XMU35bEVHCJemJF/lJacI5EFUhDkt9W/360yCMc0tXb3QcwbXGqoFg+HqHseiWTl
rI1OoYMBKLV6uUlFukJcp8rtN4oeu9uGbv9qNXrcFNJGZo1vvds2KqRx0ke+wvYA
KLjDFTywL1CE4AUHYH7xJ0hg+OTONmc/yxzs4EXQpmMo31uGl2BR9N7xSYpgMZq8
nIFUsa5s0D8lQ4EH9cTS0WZd7XePcpnfMfCQg4rTs4QozeFHvMi3HbTK7Z0TJBgf
NqNafMpoJ9Iw2GlqAYBveOR3tHM2orhcZVqFwYqpSS96ftTKNAHpzJ+2y8Sen2+X
ku6qV+Vpyc2rHZLinkPpu7Wdyx67E1rFVpow5cAvRsaLdmMbtBYYBmd0+sfQlj8b
v5pquHW7TCaNnzRscVdXqJuqV0kRO5slEmQ6e3q7vPzNlNm8oe5efoO7b6ZcNqsX
r1aXMgtmbPJ3zOAjZnPDQr7r2PEy7UQNb8rhEuVUQECdzcFX0ssfx1wBCKfFWl5a
g0SjEnG3EcZ5U1TY7yG/EiTfjxNNYT0nL1L89l3LtD08iGUijIBSpcmeyZObYML7
aiKomDIaqxZtVxBx0svNhqCVOi1e4Ab8Qf06oMsHD85+amwGYZzq3vL1rUI9Bxnf
jHXeqgdYQO87JpSnA7qQu5yqIvH44a3tpX86bhMa6+Aj+NjaCwEXgPVFJiGljWXp
SOIdViXFRiIzHz1N+XRl2DkKyMhhZb4DxZivfRPDf+ipsjNhIOLd8t+BVjPGhcex
h8o3Cro65v0cBFBY7yIxFSmidTy7v2Y48NnbqQywK/nvOz5OsTsaAxpavWUETzUn
dGjWdknX+xpdpb1P2i2pW3CCnAJ869Zvqtipcwm/KAPp5483eBaabclL4P/3keUI
evSmDx+TbsnYvKpczHBOQKK4DMXKkF83rhQ65s2yodFdmu1Xv5Ex3mt+sVb1up3j
SQoVIL+BUQMt+ErvHAV8P7zrvx35yX4LF6Bn1rpH5/TQJdS9/EV2LDsvH6vCe/wE
qsimr6bEPjIZBV+7OZpf0lTWPuPsfRG3ks+pOkETxCyUkZgXzmoHLSWfQfeq90fE
Aztt9aSFuBD5h2wUWGhnUgbsDbDnkX/6NJBacU+yc1pfCxQzRY+JkEv58BWrhPxu
dPvWVdogyPV8ZQgDv/wLzH7F/zNRmkUBixX94uoE67wv8jJ/+DppjaS4jlnxTto4
f46cRfKdK6nLExzvD6lOVnlrxyTMcfPEUV0yZqMwC73SFp/c2uXZSUPiGlux+Yfx
k+7xyeKu6vrGw8HrqMHCpy5qQQlGnK8z12FG/R6ymiy51e7hIRQgYD2rLgImi0Fb
qL139Qor70DyDkZ5aiYOrpwDkhf+ilwHvZfCJVCGnAqd98oK3JiOtTTZr2Ged/L2
+q0DyuGkWM0gsnO4JFg7Kd+ccDR08hdqXlfHNBWweBi7r7PLbK1zV5aozGuJq7zN
GAYFha6dnGdYYH/Wj52VLOqJlnFck2iDbgr84/5tavEx7XeobYM/NT4SKyQaPtMO
tnYe7uLV5ndKmHl+ofbxamEksIGm7gV1VVprxbGjCptT5xxdl7m9P6+cVMzGu+EG
BeE5Sg3deaAs65kQi25REyYdl+OPJLxIzupvy/ME1DrK6deHnFTMr7Ndn9sS1TAG
FGXOy6/3YNrSEv6A8SMcib1J1IjxjhluT+X13dDqjn8c89f4K/GalJVgxz0QFODm
3BcmmaXvi2LiTBJ4DU4SIicFYkt/p9nTxic9HsclPoHnCm62QVpL3hNEIf+0RQCo
y6BoOhRTXgAD48+ql50dvOfkOAuJTYcSgr9JMrOIX2edqiK/VEozAVPIBh2INKDN
vKiF89jgMxeX6kFsN85nVLiUrg3Jj+6Lm/TeT8IRaFc9e/6pYxOcft1zY+GcYFt/
NIzATzuKB7BxEgFRGiW15GUKcoUqcIzsBWenyhEO38Xx0tEfG9zyaY+z9BuN1tZ+
epipuP+jAh/UWFcGB30VPYdTJoH2t6/6Xkj1zrhqDNZU/TL9VDw8MfbsdDhN4+yG
tjZezz6kvFNJdrYI8Barh0h15tuUXoCgfvagGHn2zFpxfArftTIooy7Fxg3Q2vjB
6bw+2VJr2O5LCWgP7Y1GODQyZ6pbhiPu8ewTIQ4V4K6keAPPDxFwcVet0k+OiNCW
AXlLlgSiieKclDs+rb8pVWI0gd5JM3PSCE5mwxH235SctR3UtoP8SB6XpZ5MEoXU
inc242AG6i054XINQkOVr//g/f+Gq9/ZGreT48rqqA6vm3EPd8dkohaGMVqJZ7b6
kyXiAUve162powHwT2VjU04ffjqqRxTOWToXgcj9bu5NSvXWG15ii/9gYW8QE7vR
5q540C2WY6mI+WqdP8OkFUKG6vhNV7HGsI0tWWnBH1AEjq+/7Dx5qc5WKCqvZVEY
UaaVbB/HfFb2rzrKytGhnq59htdihKZXLbGDdktFMcJqyBYAVW+E10YwfZCum1xG
pIg338u/rPisTpGXi536f7S8tGWGqzj1JjfrKAVQkZlMffArtCBusPBONRQYZm56
LxjPL8AcFX342t2zS/ldRQqLobjWrxST8hj9dj1VXZCrAgOwMHKh6AZjr9dKx6hR
G2OoFyfoPdzAtJL7acefO1NV5kYwzcygQu70a6+oqDksL0qy18tkojA3NXFMXHM2
E5pJkKN5VE9vbTgiq4rC5yKCaK0ADeG6GwY3YlCchrP3mtf1CaiLdHSUQOmazb+z
NQmXX87CWU6owgDfJrwzYdpCAHNGRO5NETf8cgZ2KZfpwAjvj4QVcODF0Vx0fUlg
lPUOoWYqillgJmPIHt05XoVu+92QfjPMM+kwyq8ppoze20Y7vSmXlfxBMRS/Tkmw
jFgHOW/O+LJqfC4O/m3tVIv08Vkm3gqzIj0FSSJOuYHeuKplQYdzydhXFSb+bENb
INsxIN/beYEgZFgesWIFy6t2xlrgAnDpTjKm458AyRgsoPL+hKX4SHVTHhRJste0
ESNaEhCZukLvWXM37OB9iRzcqLdz3cOkT5JL38Iv4l0X9jN/jpsN8FaeonxXFaBa
VXPGu4nTC9spnSZiO/JOXSUW9WnluJ/cUbRy8UcvkVtlJGGRXt0HAiHMKXNDKFPy
NgZxYsi8GuSGcxGcU+RwXutDbuEcj70w4yEVeqW/d9Tq9gN7R3MxRYvK9OW7AoXm
nxdVL2mMUH+jyySuIwz1ql7NYjXFSXsnM4kPkp83dpmqCxCsZlVhrp9eAEtBY9ka
gc/RXd1ziyWzfviQVO2lGJo/gDoi+/6iexIi3LdJ86tpTRvJ5Ld/gApJcQQhuxYL
6YcM6y4Atg34A9DprTq161dWzxkMLghxkDVApevHyX/soAjejuWO+0yXhiaSpDw1
fBYmsMY92kYfMNjdIWcc/+qYKvAdObZifDHUwK1Zm8SCPMToFKp9HqViRedfQJyq
AYC5JO3WGExBltqwhu6UMOwupvCe+8/3itaPq+Qb/8WooXFhGZ0Eqk9z8+44dQRz
bf6f3Z9CCveb+sVexpArl/eTyl2M1nygkHc3JMADZKcWqIHsI62fmcIGjadnxPu+
woicWSirTV++Ov0gQwP5G1N+mNifVaHWcjt31oO4F+ckUMQIDLdA2aVHdalQaRa6
TbS80vK3PLJ4lMFtbcD/7gMkkWg/YVR8KIrzMyABtvA1N4WRjRwudW6OXckLU5Pf
Q24Uu01L3yx7dtyREwfYNaLKLkcrAJUUNs1L+AccCGCeKxrwlZ3QWBpU7wzQ638I
Me/hoeaC7xi9GJBYoDjCpxbyCj9lgf4xASvc9RyjRysi2IZdOurQRUuluOiqY6We
ovPb4rfMnMlr0kMW0GYQdcpbix6cXf8P1AMh6cVi3T5owhm/z06cMzOwmf2qF5Bt
HxhSV0GumXq4ctAuJknp+kHbXt5lO9a9w2tQ7j7HqHRqeORaZdE7br0AFycJDY6O
PwHdXHbA7N0LggpCQPL97wZ5s+BVMDk5I9SoxLrWQC/pw2slYj0sasPsScEM1YbJ
GRraIqC0BFwAkVO40AA+y/vo4FNYrlwKxuMFvoqsx9kdbrPmA6MYPsHJUW0EL6zP
3J89DEuAAmAuv47Wwjmw7jq6ST6xWRgTBEz33VTKnsj551umdrFlGdG2ujBWfaBv
TcOvc8MugebMPkdNalWvq+wQ/ZHibjKsDI9Q3sVHCZSilcyreXlT9470D87Gs6qy
vufe7KFSARIdcRrfUb75PuJt2nM166bofOVQYxmv/bDMfZ89aR324zE4x486Wihb
AgNpb5+Xyk8LSeAAIrOgoTC7By59wO1qJV0lLBBILzwGOtJE6BS2nD90tOIpI46K
ixWu/ro1kI+uP8QnA80TusG0n+CV638pLdpwGxjyf8lfLl5aVHDYuJxFhw0LYfJ2
Kxd6BllxTKDxPX2PVi+My1SNeeYvnaJX1lgZlENakXy2yjz6Dtd8lYEWymBpqnVH
rmVXfNlQjaIyIrj5yTe+gPBNuWDM9VOa7aHOEPDXPxPuH1SMlOb1X5mQakm0HlvK
hy4UE6rRKN8OwQXjqglpdAXJHoMogO+q4/Fk609s+cE3nRZAGTGj6CTOI2VB6Orw
GK+2yi39zwtkau8IhGF4066ZiykzSO8Y50I1Yim7VQ1UqsyV0oEt+8fMZmfP+1gi
ohulJlXOs/KgZdAYa23WTQ/camaIm/cSTYJFasab/j5ZXnTPUL8Dcg2O9VbPreK2
C06GuGnMm1aplpUkq//ezMLpks0WD3EecLltaO7TIjiQt9kd50HrTNvaxvFJJHm4
gU+os7QcSirYRUL6QCJBnQy0lS3lzpGzmoa3YNTYo7OcDYcE5+M9XG8cgibmbgCy
NBkGbl0XFAO6MdvsWLbWNE9GVv3f9yoSqAq3xtTb4/8VE+3Yln18EtjZwXqS86vX
LIitgNG1iHMvcC1pPjzt7DI8DCql8XAB0dzFTpWl5DaVabxvduFxyZRpNfzmST64
4aHTDG+DMAyseZi861HlZj5QgUmu2K8QHnqrFd7n2dO68UeZOeLArH+LmeMS22A2
VTy/D2Q/ZhL/JKALEJJSA6YTOXutDWKZemzlW/m2MlDeLNWPPoq70v1zQr1XJvj+
9ND0fW3Re9wgOV/jmvCpheHi7Z+N+f+SVForFDVyohB5BeGfEgLWuj7mndV+Y9Bc
pH9SefZI7MDeCl7ZQX0rvQOGLjtJO9Ak6k2UgYiawLmp1AiUhZe9I5fZEasptjHX
vkhMO2AJ5s2S382mupDRHWd6YniuSL/U8De3A4ROxtK9SXWIwt5msCH3wksaK2JP
CSW//k1x2Wpz9SqcyqBIuoQOagmiYj6mnXiiWS5c4kNqi6vvIfwHKFOVSIglfZ0A
pAHzqbcbPPb/DQkSP2M5e4K9+xhUJ3QRaCIAClQgkFZLG5UMKtfvxOrknYiNFy4z
ZsaAIPJSt4EHTGAL3FFZlVQiq64S60qruqdpgeqkoWSZYtk8yNADMjcgLi65EhKp
GACpde/Es6gIuwoouBGYlRh++DXg3WVusOGAA8Nui23seF/vn1twxg0qn1DbA0p5
QcwkecbeZgJsrgJ0QCHWFVJyQYQH6cJLTiSGRyKeyMomoFxhRK0WzIUlsl5acpiE
86OikYF05VidOsIY2doPfE/8rxsXoNp734v1iEIQoZCWRhxV4HlGnjQHF1FK7LPi
3MtcmmkQ8QHgclGlhxzqLfCa84L7ksR2G+sdi4PsvJCu7X+wSZ+xAsS4epIhSlBM
y6OO7Yb3nCuhezmdTE8XvVH4kJRVBiWon58W+uhEXy3jJsa0/07IprVvsxz/zMcI
vVkm6VKKEftxreeM23NshuEzuxBl0ZNnTFeWD1+iM9iWrOFvYT6sq1edwFYjzQ+x
17hod33HQh0Vyed6u7YhC9lw5yOi6whTtZpKh6Dq9/vTLOdYWeW2JvltiFXKT8RS
QHVPClKqCmLDJzqvPSCmqza+B3m6rdsCq0L2sWa/5S52ouY1bJe6XCko/cjZzXwV
d8lxQVu7HXR0eXRwzXJCI2OJfydxbHCmmK3kPO5ZryuAaEvkIPxAWsWg8jMFLRrm
7KuTkFxNmRxuE7/Vc3rrE1ST1Z0PM4aflG204zFEkYaXCmIzjzA4V5Q9NanW0jcp
ABQ4GDRNJrgch2PGTfFtsdjc3QiMbPKMyrHdnXkmhcjU+5vxNz0Nqs2FJfvf0q6E
y2PMbM1LGMCfHmCPyYRYnpf007KvtyANT2ZPt2yU4ZKRICJ7qZxfW9DjcDY3MlvN
y2KQ/FJE5hjYqrld/pAlAjUYMWV4pr3QTWxiRq9I5+PMool7gYoHwoKFXdrCyNoR
uaXp/JwNtRLeqjZ+u6j8ZI0CFt9JUWuGjXW+oUe6PGcOzzqGQ3tkFN7rWL0xt3DK
1IiN/io/X8HTQm/histzW2UQEZByOChEjE4zQpNbr6rOlWWaJXuhjklTwl7pk1ga
E5VQtw7NvxTqMGdEJt4abjU7OFR+bUYG0TJII1YpvIE8dYXA/zH3SF0xCdFVYHmV
JeQ84y/Z34qtvVlyQLMixTLU6XhSyV8K9dN8ufg6rLHZY8G+w7JbqmscYX4wbv+X
e6x/YFraI7nWPkFr+qlQusQbx0bXMO+j7w2W8ZILCWaPTVPbBjI8HIFeGd2hLmEN
KR6829bV9Ym6ELTIjOyVhqD5BDvbKqLQoi4fPwFluzt9dL/df445+RDGoSuVpNiL
/Za8jP6m3dXVBRRahx6fPMfFaM8gTFx9+IXGocw9824PCFGgjhHzQkmi+54O5syX
V2EnXwZhXnUP8qx0qVcAbJzWYqsp7X8l/FhCmZ7d8wJUvlnadwUzZo918mVBwIp1
19zszS9C1RH39/W76J4dlGKovvNs3jEueZgI4+AG/G1JH+pRMvRqYHVDDnWznq9U
I6i2XVLr2x0OCJnY5JSSomdnnd6+0b+6EWUDkwDNyTaJGM5Dqfbfc9poDCa2rzcW
SgjVSbs3oNlN/4+D2GiHgY4TNBhfEjvnRVjgBo/VXJRxYgIxFsdSf26Z7KB+aIs1
FlbqzmYcpx7+1ysECwdC4riDGumYFIJTbFKaXvp+BI2kxquUMGtj/DP7Pqa+xI3g
LLstgKs5v44wnS7F0q30X1LAmWqXTuzJWaGzhdcO91YY+XRbYUFsMu4/qmBwLxay
MA72LxI4R1End9Q2GPscM9w+mUAPjhD+vMY7+haSHDAECmzWtCUTVO3NL8xj/UMO
LN6BvPSSpIlnQl0I01g8MnzqKOb2JbaLPwfYoHSqgM91BW+Pvp/roFioiraxE1dY
F6ouAmCfbob07Zzszb9Sx9Ab1EqaqZ+2cJpQ6O6xxHYZqxwpXt7FJ3+iEaaC0UN9
VxSzDQA5cOlIcBianyTvaRDX8/2UF+YIbW1+M1s62ILfr9VpavMtvORd6NlH9HT/
0sh54zotQuP/5q80B096dbsmIZkJ4HX9vDRsW7bwUgiTd0qPdWqJg1Y5ZkInYRVv
Yb5xPJqgtdxRaZ1yTnG2D+/cGM+m+uL7KxVYgmwjcx+jbkU8ROPzKPVZM3FlLyyO
ZciYTRGKI6llposlDVAZOWGP71nYqW/tvZFNBaRbC8Dqu5ksV6xlXbNebcRUU63K
/VH0EAYGlOxcOHOt/EZFrYLeMb+FgefrQvy/K696chGk07Fvab6tQQX/+ZD6UXsf
iNeLrxzGqVE5fhSgYaDikr46p3P5nZzCdJ13nfrTCMcQ3MLgIIvm54jwVPaBp9Z8
Ubdwip5dgTAc2LiDVEQBHcAlA+JUyYc+3zS9YZZ817aBeRGHdedLg9UznTurqOXf
mK47lDNcU3cUR9eZeguZrdDaYYrPVKJbaJsJOHNBiYSbngV2xH8Hrke8y6MmEdfd
1tKZul4INzCAlMCsZ3sG5YrzyWwWcqc3lMvJpNhloFGL1uWU+M1FRWe5OKKbBTml
abMO+i8Jn+Eh/7C9u6DC9zfTV4Ck4qOV3V0B7lItRYBoywvn3vh03NMdTvHSo0lB
OJJY4byszaRAhBZVWxYUrwdH4K+5Tk4xbAco6tlFPPxwyhIk03R3mnXeC+fuQnC8
w/3DHVV+qZlj5fvFzVGAVfSp3CpMDGy4Fcvc/rpBa8XPrLbijinTk/+P3/wwZOmr
S6IZlwRPMJs8Mcb7ChSQ/DlTgr4mdmBFjp6bjwuWmOcHbMkjdnSGunvNgeWPthTu
40CZeaEaMhjV9GA6FiJZOiies7hWQEcjZ0OEZQPHwrNdUEzyrgYx6W/LQCn5pwmr
WLHYIL4ylLkiRqgzJ3ZPzbN9m2lTN8RmMzvzlCDzeqVZW+RQCSH2HtrXoxBAUk3N
J9Fc1qrwkr6qL1oYDR7LCximnpJ754/TmfYNxBI4e2pixBdrV1P84UXwLQfZa6pD
IVSL3WLtpnzLzftFnhxsTj7kVL1PT2mDOVgZifLhXxLb4JLmQVGEu8mFS4NIsG9w
0P7qSfpuROjsdAJineuA6MIloi70LGLhjFRvWikqVKmtk8y6YAY89MilI/D1VqzW
54KPfdZGDre44ZQIjYZW0gxWKhI3MYkCLCTEfWFmjSrz0uIZzMcFF4cht8qHKfyN
VqFlQOkS8NmJACG1OxfHoGVkGnwzbC0APg9UcfBjaaaiOQRznKeJKg8k5o1l9DD5
NrmV4+BFgzMc4ujITszvC1RHGDg44iCO9mm00GrMAAK0hrAtPyY0GdRXxhaTyxEV
YxXvCAOXtsvJvND1DDKl7HJ7oqayLuPSDd+8bwI+JD6zU12BUCdQuolYT2+ACbjI
8wWL/WGGUf619i0I8Cvub5UxX72gbSy8t/lXFJDNXStDEo5dCeLSjY4MIsWpfwZe
IEZRMKmVJtTyRdOOjSJcPBn/QalRdavg9KC51U2ifT9vKEGQfcVLw9zTzA5AbyvL
OewsPIUFrGc7J7yOjI2TOgzLvLH3/tevb2VUu9pOEFZI3VKf4vb2+XuNY6+b7XRf
LwUpvEtVI3LgCn/OBdzhmup0toLgKVLg+St6ALLqnVpizHjZ5S1xkyCp91AHzUd/
G3CLSm+q8GUlZwqjKNYL67qUTIwNsc9p4S4yI+hwXSt9igYu/tnc+M75gbqUE/kk
h69CDYW/yoSeEmj1sObxlCpLLpvB9azqGqPeWyR0W1b55kQdnZFgYYO7KcREnGO7
g5bC0qAsFWa96JTmU3KyCvl4LEdb8gmhcgVmPV4IDuQQG2sB+A58AzJHPkPZQVN7
Z/MYl2C0XSbt2UE7gKlGQv4WO4A0+TyIYndU1kQn+fcJahvCfoueBMGCh4lgYusB
wv7jkIEFzrFBVYPRxqh1Wz0rgzU8UJq2fVf1qiZTOZni/1ycQ7MqPiwejMdEGXI4
IPfnin0er1viRp01zTEbNslhERdvabrq/0Dq+x5S9jlZGsOjbVP8qC5dDKq7kQGb
P7ZGOVDDN8OJdZIsh8841GnguBVGgrTYCoOpDO5L518UUSEhtjPCGuu09fKrNzS/
58cn4lcvOM5VRfZhtLfIWw6uDSmcout6HvpTr5pQB1UiotnELQmxgpLJxVaPmOle
GLVJJTtnl8LHjLcpw7EgSPS2VGedG09A1+XWJw75Dq+xQGq+f50tgCnIj7/X+3+D
9rl3ARDz0Qdg9i2bLDziJCrs61zYfkQk9p9XgGa3EQH4KZyZm6nz5KGJTNwYEbju
xqR6LQ/FRmXzXgUPMYdoTtBrjnuaOZeYswHfN9xHg5ij7Yo+C/MdyhYiNCDGqRmS
P061Aa3U1QwZqoLT11VGREsE1F3SMNiO5b5ekDiXj2uDgBbtmSmwrgL3AstekFEd
tJkuI3FAh2GQ5bavyK1Zyayxifle0UtKBCtYzE7U/Te3F2h43YOwqljAfRfMy2If
S0ewffUoF9dVU5tYrsxDQ/v9/MNafA+aJW5lssqax0pNH7vpufecb7ElC93o6yYE
tHz+Gv/fW2uUH3fVGu+N0rluwhQLM3qSXwu459cr6HLFRFIVfkvKMJWjlmZPxnSG
NfzBUZ1h5eKH6Y3Jl+HcaT1OHUuEnd2meTSWDP3jPjBlLDoQVu9ssPIGRFTEONbt
DY2/0/nvJmS5jZGskhiyKCZOr6FPqeCe+Nz1TeGdk0CQrRob3+YaWM4jce8No7bq
gSiXviEUu1TMUJRGfaBR0AjMP4fM3QVI67EUNJDxanOuDfUnSD3EShfpmB++zYCu
AmnUm/iHX1RrpNsHNhAjF6EYskya7UicM8oOIcLLW9BPiSK5JAyrOrXdGCigGcij
tvXbEsc2ul/hjCejQUT4nvANXxJ69OLOLycecP3SUG/NtmPtz1V2WWsYgrCZkPzX
RNLBSxhi7UptWyegGlEM6/xN3GUvGDFaJL5ggTxiyOjqhBIDh0bXZ14pR8M/51/k
I2BbIxE6V90Z8eLqA3uEJsKc2DuYjYtjite9+nljSUhXUJyyjVF1pIU5prUGvOaJ
PMKUy6WUkyLg3hk4icrtcpQQRDNDFwXXOGyh1ll5khUflAPrLKeGT6VAgpJqLL2Z
YkuanXcK+qDpUvCXxKHM+MG589cQ1FXWhWZjBquXWD9MVFWD8DSAwZ+1pTaBagLk
+g+GWJ8Xj0k/StrZQmy2ZqK0Hd02bKy4OZm9e5otaQAtVuEmU0WquZEC807Vhsbv
6JPUpGrOC2vehJ/k7y+L7IHolpcePH0sFnLbaB/1n6fcKnQgMfBPCdVPn4bgP4bZ
4peM2oioEee9STUEcBJhcYMcRTVadmXo0nB2TIwK/y8/PUKCXMZquRO8PTQyD87h
4Cmdc+a54DBj6EvdSA3ANSnjl39zE4gbHP6g19mUt0T9W9N7r3wuRl6sIX/fQZDO
2FbkGQ9cZGyRG9Zt3hhxvTN4Am2HdIT2b3Z9k3u1+YTo4H032QsIT0t1PgT4PwyH
nK1ho1wzkKd/4Et8VLkFM4jtVt8kl7hCorZQt6Le5LUvNpB/uUNQdnUhNakIJ+YD
7HO1mJ8w1P2p1koR2kDtOvAaY3Pvjs+zDZF37u2Z1QB5PomvSX3fWVOUWORUUUeU
qmyD7JsA12on7EkNZF4OJ25Y5SNB86pU1fknr2BEQywfI3gqe7DXYvb4X2KtScEn
jUlXTGTATmMaEMfZ4dxrss1bORSFmyBLipAYUtW+LFXlnG1oaWPjipObW9uvgBQ3
inZ9ADruqmL9mUAVyQUnPdh+Ab4HuIbVM+k5SmlnU3QNjnmC/wriAcsvEDdcez5Y
xDYj4axNo/aKsZ/cAqWsm3nkxIfGN1GIwl8eHgyw5t+GP804lg3WcYISGzfDwXo4
CD1FqHCiwgRC2Flx318D+TDPrYCRFI2QGEvw8uLTkvIHEF6L6Ddb8lxSHMmvvJk/
aKYnxm7yOKT53mJbY3ferFlRcXgecHsS6rAM0AiNCqX+5F5IU0u8KsImqZ8PzOD/
ESxF5Qp0nAbR3PidIlresUxIjnto6bT29YMo8d4yTqJoLfiyU3N+mBibohObghpy
R8Z2jZwscx2qqTDOBzQAzcdzfmbbj8vEfWEk+oyMvb8jGQhMU+bpCAVgJiUOTdtX
33acRCiVZUkrPAS+ShbZOGvSc390q83GqjQy5HCz7uXXnpP5EKUZJnyR0Jco2Mki
gQc2sWfFAWgleLyhsj/KIslnAUWap+yKXYAAljM87/whz2y37FNAJ7wzJG3MHJ6l
wa7jx+k0OC7QRFZfbSuzEw6AVCWJaJ27vUBtvGM7NLhcepeuD1M4/mG00XManopZ
iQrrWyCvYVhp+B707JalzBjJnZ1Yl2C0rYBYLnmPEYPETrGioqeyf4ESSzxqo4v7
E+eXoa8jzSu9Ar0vQ5Eu7rhEuKTt04nUIqtL0sZjlGC034xhjXYdXOHei2S7t0kh
OfQjYXu1IJGayefjEpbTzXy1BwbYxv+WQxuoeOzCbNC3FsUU/fTsfN+O9B8SSCJE
/68e+SCcW3Ox/CHK/vUJNHGo4vsVdqlvSPB+WXqL3TEtWTB2F1pIRNRhSsHkO6KA
yoK1WQc73cuRe0CesogDydNhYLFfBKaOMF9KGT1CN2AKDygFMn1zZNUrBqOr8Pud
+E8rtYbYmVRbmppZIXiwJYVY8BNWRid0eASfmow8uMwSyajxdMVBd0bAncndSe1B
11kB5vK15Pb6nuJI831v99Zo2/KHrMXu8SxIHHkH7a06AQ6q20ym1E7n40LH7scy
o/weRrsOJOiQsXlHLplsMs/n+o1Nl1s9GJO4r2ch68LIN238nZZ9oFxreMSZs9R6
LMopEAaJDHeH9un+GgC4r58GgzfzRJMgA4huwW5KS46w/uFCb56bduyTiKnhIDL9
pYD7BQ5cOzJKzGHYbgLJZTz6U2+LjGWVI5++r/nRZ4ZgU7zFH/1PNeF9YGUnk2CJ
7W49ealcoqwg8jxAp5tgDee4BPLGDoyB43gfrY4/l+gHmGVOybUCU+XvdC1b36nJ
PgUfH+T9Fz89r5xBieMuvuHqkiTDFrgyWZvtBxLoJCbcXYjnUe7hPQvpQ0IagTZ9
9IUIjpaI1YPO0Hpp3NcDwDvBxqYoylVYL5DgQr/Q5EtQt498MXZYc1kRUBx1l7dV
rtsAnYoMZurCcXvyXeaBHjuRaWfrC9NBQY7hSopuVxuKx5c5aKFpb8A2ofkXKfmU
lJmJw/e/DUj7cKI2Hkh+fqApJrMWjid1jdj3wRVrBMufnZmK9KaASAezCUDpQ8PN
/HzIrsRAFVkhiYEzA3pLMBvWHNUirsNB00RQ+FUTThBaJNXzSvPYNieBkEXeSd1P
LmOgsokiQ0ebQmZFWKQXy0YFVKgqYaEH8OAwd2qh6smOFSd6kokfLeDUZ5Njxrgb
3HyarQWtqFi9k5JA+VhdqczkF5lNGYmsCy6bcm9k+yCtyGZflglVKhMOBpk42AJw
6JNiDA3jw9c/ew1x7xXE+nhJSQksv4ouc9EzPq6ZigvE4PjYBCRyXJj9YBg4RfY5
RffoCkLTRax58z9jUGkqu9y6fSMouc4EcS9dMTSS7DD3Ws+Z93HuOW0x67CpyKf0
fYzCa8eSIPu3FROwWM4dRn83h76s0+RkrRo8GfeSqbu29DqoJcYd2A9m+rsVtLTT
EgKztGukg/CuMOnd6bnPwfUphKoQ8Y3LoOOFfnRofYb585OPZY334nnxAa7zFTSf
8cch762F/Huk6PiMNc69aEp7YyU/RLbgny/cmKJRomkGBv09vtTxMBBx8WsMmJ/B
4pLpY1mqNMtgGjIUXUHrXt3snnH0a4d/CCy1nGD5lGkYGAee0GKhqoD64JzepRv2
N1eEWtsyYi926EPp73dMTH0CrY0tA67mo9lFtgah6yHgnoXlbDYUGt/sVLusjyuo
IB0Wi+pYqekLJNlTwT5y9Ce8iPo1hGb4PlYPUMTZ/0eZvPG1Nt8IgwuL1ynYyg8W
oKSI0nHFhrGEpoBKkKMfSxGOtgp4xk8yIjiXm9gys17y2lgGkXOURqDjGnNDYeOm
FyuoDkDQ/tokildhtM7vmyjzrrJ81vQI2/9lhUJbP3cmMJXnbPHA7nli2VGr/0P0
AOBl1FQz+Gos5cI6aOjVE8+oBjvYKVtB3KHy7ZCSyT16Q0xWSrPS/brn9D8PihwS
CwQ6GhC2TwEyb3x+v7NHV4wylnJKQxWDqIXtKNs66icsA+snE6tZX3r137nILKuY
AO7OPaQAF6Jg1Wo4D639HrUlUYKO63J036zJRbKw2DUX9FZ0zNYGVKc8V3PIr1q8
RitbTa/XiJxSc5gKB/usjMoayhIX8jdFc8+tdkWBvephLyUKAo2Zk9yEcH1fUcUM
okkqW5jrUCJRGJrqBdyVibDteP6sIJ/cnzAerWeGQ3IRYy0d4CqZ3M8L9rihqcZk
HcoTjpIs/C4sHvlXRKUnzCZHi/k1649A/Hwxmbyxi05K6bLc/iPPmCxGpEPBX4Rv
Xrde0A1vIAxhuFH4Hq4AmhuAekIEIJR8pJBEOGWcGWBtjEMXvSNmGrn0lA+peMQh
Vo5KP3ZxkMPsbDqN27DKtEGgRGSTQF3j59QMt2Aoe3eXPiUgDMtPIdLMZw5v0POU
6CiAkGaU3kGulIz74JNQSRmhMwnKXMfn9rQmxFclejYm/ce3Go448XAbX1u3iDib
YYLNtfkM2/sRoyR24dP9b7JSPjXXjM6uvRJTXX8xCPouE+MKNLGBgQIQREYhhfdS
ttk9TtlSrh4aZmfmUnZ8FNPZIwswi4rUIPCBFce9+T9ZgCY1iznFr3YyNbGwnHh8
zRGfBObJu0odNBxuFxkH1aCjJDON7bseFRAJ9FtTGdFNzmsHqH7SjwuiH96VCNwY
altp87j6cDIL8Zu9fuVD8Gj6yBnYiNpHlZIF/Ckj0tjJe+MKy7aViA8Nd+Aoqdny
oP0ksLIP2W0fO8ylcrx/VNgXq5Aa7iYLnXkvQCxrz78NSpnvYu4jjLAN3Pk2az1F
tGkcY/z7coTPm/kZTV0ySzfNLUIhwNHrYM0FeNZO5+RTBDoElkkEPPz6qh6GKqwh
4Jd4wM2zln5fXEhf2dyCz0tOEShC3sR7RUuIxt4+UYug4Rh4WUysb0mqWmrEOxXr
6O9JCXnkj77QKdY/mFaP5UC9fniE+BqyxonIKqjIJR923BAYyi9dkN1gjef/zp/J
KZgqcLSgfvpF+uabdNdDjkl54NETn2iXPiSrJqkmOGzm5UjKmVHpkF8DN9e+fE/W
fMOCPx3j/c/NP0p2hV/XIKuhcgbnjTeQisIImRAyx+qBICphyeZNfpz2bklyxHWc
ClI2PfguaOgDQLR+GdGW6fTRC0jQ0iLtol2/AVfJFEyTrKnYDgb9lHS7KnEhFqH7
iX8vsVL9+A3jdTEGhLelBvCZ65oo210uKSJQroDhuik4j0E8CMFjCTKv82rjBBoZ
FG4tcuamsNI1kzQzDDuXak9OJX5NQ8Ax2Wni/cRtSAzhGB5nza7G7v9x2PagQdL+
8tD55zveuLmwMbGGvV1qAK4Eh/JF2g3O0FCtzqs0+DkvasbjAo+DetJZA11ZLrBG
lNNGDyKM1cBopGX/wXDIk02d2u/i2fJeI3XhSfI/fh2/Yo+eeRMA3E1dMXDJEeNU
MVYzBiJcu5o26dKySbinQjvK94szssrM7VyJAa2fYXnA2dwouniHh56jWp5OQRq6
6X7t9VPIPRSTZy3sE2sEGHQCvKTZUKh4pwEGBFD72AERvUG5vQ+EU5XpzILU0lwF
C7+5RX1dMO/6XH2f0mtuFmuLmTkiS6V+3B39D6pp9yf/javffpVry2PBtWNCeUM1
spXUFWufJY3m3/J0f59H484yvbnwvIhdE9w8JU/5X+8VUH2qu+YKwuZwT618DyV6
xNqGTycpKbfy7/p5wUz3MJh964BG60acIu7T6aPZWoQt1Ujn32trgeUsyKZjUk/W
40aHSeAe9+jglFp1TPzffVVxb722cFWXUOEGDcWCAI5oR4GAAY1P4yDid47Xcib2
Xhv1TpgPtEhrWH8vtkv+htlMLoQ7rD7/5jqNYr0UTw5fMzVKEpTE21T7IZVL8/DW
RKlp24u5N/m//HwqznL2vTzfc00GEbzc6+Ia4zpJLEnv+u9r3J5GBrmKyBD9Z+fl
klYEL5jKWgASwGE/dv4gAYor99LMGUoJdkn0bqnbWuLBcuN6s/Y8mmieJu0nN/rV
enMMIhGBdScFLLuEohgGmLA1bl2CRgJts3ZkdITUBQnD9XRcbBUagzSodz1If/XO
CMISQMnoDHPveCRuqaBSFp5xZfxqVlu1XtatJLxMkBXtGjFSxfZvkqBAPUvHgKMv
eHLVc/gnuQmDDhRux6GRBgnAcsFG9Iu1ThSH/bCMNIbWsoWrdrXY4bMFRS8gZp3D
H7CweoACDYMHvc4dzXnfFws5WrvvmdxnexFm4eSE50o/hr6cudA+3lzkjW53XwBE
SM9ZjfJCZDuErI1g5UrcMpcqvY+wYvE5G8M5nYtyhW28DcpemdMJg+BzNtD69wQo
sFAqXIOwWMVQzxceR0jbtWf3yyIsSEK+k9CqOgoB+/0TvWhWKjzJExLhpGNBqOOE
+EONqqW+3heWUNcIrFcTDF157+LeSUR8195jXfWk8Lj5qigPYxurrXGTnPqsIpcS
cSHcWqX1fTiX7MZIwJeflRMh16w7Dsg0Rzdd6OAkwFuaZTlHCQwbIJElfw2qHigm
0c+vbVPZnzM56Wtkd0nQVWw6zGO9ZfAw4pzynWP7VsV+GYzf9DIsouExLoCsu18M
YL5eNYSazp4dnKuC+Mqx/UBWz4o31skwNMUEmUbHH7f4RuceCSMuC843q2jtSLpk
zlixkCbPAkWs5IxygehxULvDOu2vWL5w8skIWn8YBaslPVp+TvIEu5QQo0OyKvsN
kkoGgQFmGGg6sSwNHu9rnDYr+HYGkWdxZwSg/gm/CjkFV9RNacI0XTRmzc0kpSci
jMjKQX5D0TVhv3UmdAKBBL8w0XmjzKKBuRHFSmRDXfNf8ekhntjVOR5/tOqXTay4
ou9V2G3Sdfp+0MOS752QEoQFMmgwrnlRxbTbZMMvGSWUma7tb2B+z45yucpx/ci4
Tbi2qj1lKQedOR0e0JnVScC1+R4E8QW3fKv6HwTkwQSvoO8nw5ml0t5dToCrQgw3
Secb1wbGI+q1teAI40wzbM9jspaGsTugX+fsVe+SWDEDnEtCJY0pCebo77W12V0A
Riw+JIPPL44AUeBIfRhCrLtf3RiAC/iaftU3y8vspHs1VTFFvC9PzjHuxbVVq1sE
mX22Ud+RTvpiTFUvngnG+gHGb8GTVmCsbl9Y/sHEh6J+Vhx43awIHv0qkPtcQGJE
7QGSkCTfdImTFv93Whm44Eu0Qq0V2Dw+EJEggUWmotYJ74tnkcTc7O6RqtQm4CO1
4C9AYiJ3NrEYPYjoPdpzvXCiCaHGxz1v1nSp5LEJqO8DyoccUZvThgM8lh+0WGbp
1HVZZZ/VdpBdnUMgos6W6iHmjWloY2OGwj3zbXdzJ7gmXf1g6GtodokspcWjcOF9
azagnfIE4u/JZPJJoheWagUsNPoy0JpCGkpvbYpj/IJIYyp6Af8Q8PyxabYxzkqd
9bi3nKGS75T8ve5BJpLCaKJ/dTA13ruwqJbTIYvM4SHOYK1DAI/zEY+0I2hEnsbc
K8YpaZkC7z1cm+fVrnPGaYakuMZdX3B2nxBLQVSn86vkl1hEdr8OREtzr4CvPBwE
q7YlAlfc/vVHyrPIWzElDymB2QeJ7KRx0Bg3ZN5X+CJUoW9ZhGEQnhu/Vjbahiv+
wmJK0De2HQKeRO0kJkUksGf0rxLCZbpUlWRYAt36XFMM9X6J21g3iq7wfhhtC3+n
gKlBiQbM+MmDALaMRhUDXlvM542WGnjooqHTNLaQeQ+t/CG48WcK9JhUyr+6bEKT
BMBBgQu4ZrCg2zsE6Qze5RA3sczFOLOqlvra5XlwRMWH/wT/FqMinSsr0id5K5B2
o51e+tPRr67otQRsz+/guWFhQIgckmmhuZA/TSIzgJ3F0QhgKE1Ik/kBkd4QMWl1
yw2Mwz6gGBRdekhissKH32r7hQ9oEOcdXFW8AXZUKVFj+aNWLKCmIyMg1rBPOcUm
oS6ZPqaJV0mi09lrYfw5rE7fxdP0MXTqZSr3+DMk+XLUx/vfMOMmUoBCbl2YXoDl
K54aEF2kMssgBJGKW2KMIlhbrgRvUjDyrG/RfpFhqwO08EwS1M8RdJ9CPxmRCtjB
Oac7rktT22+v5DTGfsV+n0m/KUKQJ0DyNaFqfrTFKbDGhBnO1nVsxhTxsJ1uEYLm
aO29ufRZ1VnxLIAO+IPigAzhG12L0iVwZXoQlbZJ2JxxDm5viPFD1B8Ic5mA8I8q
7FYIWA6qCjZJZSykYBi7cXjCE/vX4nJYgRvSiw6lWS22KIhzB7lSgkBCCKNj+/0O
nJhPf6B3HgVE29D7b4fTXZDI6zYugfDHHqZZniJ4+cKJiT9Tz3AIVcdvg6KUtWCr
paF5flYkhmqZZS6y4Um9nZT38nkUairagM+XRsBdPwOpAd8MaFuRMhkcJAUnsQPU
ZqzZW4VgA4OkeeEmPvf71bBxQe96/XLq1SYspXpP9t5AG+5qf8b6M8aOIYjkMVfk
bVh2H1MDwQq3Sh6gSR8uvCwGAHDnldSfESB1OV8TPyLfJ0fHReWqR03eJwnmcfzy
XuY5DuRT7ogJXLO//Y+Y/OK6Z3loZjQPvwyhcCqZGkhEYuJYlmjQRDuXGnVRC/0X
sQxT7j3aJwXPROLVenxP12A2xLJapf2jHIvYPi8f2pfg3n49DMVcTvX0OJd0sWYe
GG957382xwyV/m/xbFtnCymLXGJMCW3DX7RR2OD/rQyML9iY8ELEA8QRf6mviWgq
oxPM/kJJmTrGq2s1XRw345TnJC83+I+omo1XEw9YNoL/hKexnNOxX/gFE0fUTk2c
rDQtWNZofCDF0h1PcO1xGeUiSDJ1Pkkj8U7QeLOSIZm+5xAO3kToqFggXjpMfvTU
LsuftOGAodemT6cV4gWLFVFxXbXRbp9gGTlJML6dDbx7cXO0qAf7rR4Bk+zwayfu
N5wrsQVVAuSCM/UyYGz3+4tz7gXQ6nzVk0aPKB5qInMuGLx4Hmf4M89Hkzc8unxV
x45d6tk6RO158W1y7u1/0GitTQNWcNmuEIs4kidZQmbGIwgXMQwqaPJM5+R+0GwM
RaeyEVNYG+vAwn2YPHoYFvOHe92SOpr+qGr2cawB6cr5/wwK+toztmb7WjpwUZvF
g9pPaaaXKoUSiLlJsVNtIqkhlHjdnb2SjfXi791kZLVUvqdjRo/PJ2GggcxAbAuX
/p+Hzxtm7K3wxF52ZdYEQO7/sBtg/JIJQvr5UsaDb7OWPwVs3SZNs+Ox9X4c/J+q
FYApcv9k/8ldJ1kjLPGrqmLAbtUz1myCLpuWzN0eBRb4IDRwkmiDGf85tV2Mg0Q2
kOEnZZj91ZpBGldYHh61OfZLR2anvrzMcjbRQL7cpzaBVw+8kwSkIhMfdNJMlMYW
S+bWzFJw4NoGNWP7R/d5aBMf0nIHPXF6e9UIyO0u2YJ6TMYixX8mA/7N8Xv9FL4P
pRwoXxm0wUD16VY/S9S7rCgnkS8d+u4mvCX56vrBScuYsH4Q6NpkXSNKkD/GozId
Y4C1I2dm/odfKuSGwCTAqwJXkZtrQWTF25O4u4G7QW/TWvdbm9aompXtJsukUunT
m6+F5isd0oYtO+637y7oKfvLe0ImynovUadiHVLQykfF8/Bpx/9NxnSgznZ+eBcH
oguailLl+7O+OKUes2bAHkj9fq6As8DARNIQlnakkfkaQkcqwxB5Lmo8l7pxvw8O
XXFqB6s9ZcQwPasGWUQEDE+VA/i2Js8nr+LOoeUp/bEOG+CqcZ2aayc+JIziY+b1
7MfdN/UTwauF0OWhWyrPpf5W/oMZtWEjLqKOyl+xShMA1a+ar3D43CwtcccJdb+o
6eFcXZgUtdCJcfCuXK5evdoeMCi7xQaeiDPLxZcsiiTs2lJh/IZDwYikjmlVjYLO
K6ttqbO5YUU9PG3k3boYxF53+UoBKEtD8hGrmfwdG3NrIP6SpMaeq/Y/km4hObvY
P3W8ZFij9jhfeI9AcZCIl0glTCXF+LqkpV1HlfV/Bca6Wo+K5jXtIuuik9gziY5J
HCaICBq1RHZktPEhxO3gAou7S9rpiMTGnzYmN0yNKxO8sUz34Kfrg2Ko4nzLeE+p
hzquZdoMkuJjwEoAfIQkojFxrdU+Zn0M9WtzQWFX1ts2+DW5USiUh/jUl9hXulKN
j24kf6LqAuhBl6WH5qZPzoSGGL/h08yzuDdzujYMM84EX0HQ4uMGXXecQbDYLeNt
bvV4szevK6HzUnAJYKL6b/DAOLuaZeHQSHLm6L8QMIQBJW9FXT7iTShsNySiiQCU
TsNUTQJ4E4NlPyAG6TouGZJ5Bh2ODiDIsKi0CQP33D6pnG6gfKJYuqzhvdtQPuvB
hQK6USpfDq+cSYvf9xsqZRxiT2aHR1uRsl220jv5t85VgudqIeOMiZm5w/ohfQUF
ejG9VkIvLlCVMp8VdBKXWJHRkPZx1EEOuvFOV1otnfDjJ71VO2sXLzt6k1VLubaC
iRbIXKA0uVG5b3g3qF6zydz4FtNLj1oPrhH/0Nk9Lsu3ULNd1b2/tXLrj5nnGvO5
G7Y5ZjYel72y+MdgAfD1ruwZuYJgM7/+LJBP6/zp1pXxJ6KJPCsR5kdzRWE9106K
egVCYKohUpTDQCBvKBqq/zMC7N3l8AlK81L0200sBKBRO52afSHZtGuQnCcRB9s0
NRHe4KjvED6VokxcK6GeqgcuZRo6qmAa6m119L4SEasBEbcJskF9SYHwPuCzGIp7
uQgGn37SaHdbVAJqV2orLyeuyo9wP1/bMUPKhEa2YkvxX2pZl02PcY9U5eo2qCAG
eldCLI+F02m/dCnvmP2PnALZx2DJsJh7PQVdLagrIgAHGuSKUNAXiHB+dogDho4/
4dMKiJKmon8I5FBcHgFvzsdDsihYT4lKNN26+lGrddlDH9lrCHSg5Iv2kjcWVAqP
yjDgEV7Y0B7CTL2egm+VIHJ4bmuEbhR668i6WouvpSHKMuA2c52qnHI5hZ9jWS+a
BbqhN59yhKNgmjy0WIWLFIYLaTYeuUGE5ok2Y+S0eTHi3x0+hWHT1PddSE9lbH9H
qmTmg3r8VryGaVedyYTnuTZok8y6HmOX5f+pgbkViu6t1USEMeJauFRr3fnsTwGV
c8lMOS3LzZ9Nf4xYbd+/RgxGROsuwWynr98flrWjwy4TgMU5i15tTK8kAC/z8Fl3
LBMJImgxXhyuS6SMBE1Kf6yr3WIpttIO735SfahzhZ8HemVj9f53r1c+GSBCg4JG
nvzgguCYpKd2VpBE+AugG6w+EnRYKee1JC83+bDIAIFdRWwkoHe/z0tTNNU6Lw7I
XBN0G4mmxyABHPewqW/K344KsbUFQGkvGYh4l/g81iZHVy3BYp4K3IG+Y3bs91A1
uJfpmg4T6ulmob1WXF4gu1QGcv5cH0LPt6B1FwKJn4+RWDFuEu7qQacQ7klKBEaM
JRWPcFotiPkmoJB5gIcQIGIRrDGYjJjPB2ZmIfhsjBwLYUm2PzGhZmS6tzG4tPhC
phoeJgkb3KjK281YoOF5qvdmXsWVRycR/tKK9+h7dOvEWfteAENwcNHxMU5Io2qP
HKmcSOnNjnqhEQSNNvrmM8gJ4rBRGYR21xSWhTT3iBtglC+hDaiRPwRRl3h6Eoli
DhluISxEmjtW4YvSqqj86BRjX9Y7b80RExyOEhtSvGpmr2otV+Nm191H+nAAozLj
Qbn5j4roIHRkdKR0Xvm0vAS/6ncAt32wBTV5qZOVSKTRvKwvuCFbJRLt0x+0tIw9
r7MEeE3gLMVaY9d6HD6hSa98Gg6a/KpDu+GApxXha5rWy/wgbsJnd9v1hBzYmgOn
oobDlmqqqHqHixoXRPbgniHpmR+KhPL4Meupw1QPxTZBqHhAx/dSGIdWP+U47MRa
x2cEpaRhtO2oiyDzjuofQotXc51EPw5CnCcJbmgF+J2Cv7Wqzpm+oJqPiXBQMgjy
R0F5xxfNrtzHsgs1rxS/V8t9O854bBJ4l2qp3DreVLlTOZLI5lNu0BM/S4orA+ww
QQuQeHjRohbF2Nd5kAyDtSDepIkVzeei5k1bPEWDv12RWT6NCadU73khiZ4pU3Tp
r38uWnTbfRJAVTnOLpqeNmJ03EjStISf7fnokrgEqa6nk8+WNqdFtNVMRsT9f95F
8db5vyMLPThocA6UBLpB1rrfjNxWESMK84neIs1iqXzM/Y1WvpFkTiQ8NXtWX+jI
n4o/EmWW9fuR6a2fUU/0SnMToNVSXx3qFZyfOULlhtlREE8d7ZkJyl2Z9maHsq+C
HxqxJSfnrvot4oPUUGMB2rPcMVcJlag2zkOiCtUn3qxzTCJDCJRa0F1uBCTx/8tf
auj2BSUWOjNWWE8nQw7U2jTK9SUzj69otYwCBQwRUDGSjZcROhfBCcmSj7zJLX9d
xWG2QiKZlWfauMTTTjXt7bLOBkSc0Y/pyBg030wNGy5sZ3yiAiUIbybARITsMY1q
uCQrU3yirDC9uWfuBqHQ5q6d36ozDXBbFIare6ffLRKRXSmTQNkT1HjXntajOWBH
V1FVwAOkOMBRyTF9Mw7dPSvHeD0SgR5OE9DTq0wXpu17O0PjnQAlp8oMlMknZntV
a806ZDKCWGdwo/Gqq5TkqT4l/ERh7YXvsrl1dU94jh291OAG8VkQxBPf6olcWWah
uMGltVwHc8Fd8eBqsHkUEycki5MagyGIIoWrvXNK+YWFO33eeK6ihSaHgzmH5/Sd
SKOGe3yYqLQ7Prkd0g/M2X3Ya/LV0cs9n339CXYder7uND/vu0g7fGxebN+Kjmun
gzF6CLItjeY7dZ0OWd0eCs/omforDu0WlyIwWnEr4FNjEuaZCgQ51F297nfg5Kc6
HLQxc0a4/9FaCyZcq4Pv+iXa/Ve5tRqQFPIj/O8AeA0H0BzElThfd6dX62W4h08F
8r8UgPyd8uu1eiQPv9o3C6iv7pFgTVKe41NxQTA/81768cdRoCFZlWlife8aOBkz
pHM+cxO/1TN10Cdm0kiWtkxAvRBuW5bQ9nanYyn1VRx6vMc5TaCxFH5GtWvcdH0E
3HjL73LpfznPkkvdEvxYV5tjKQ+dMJDBBcdRrO5Bf0kwgoiXqPvA6k6g50ep2gxF
nibAEGW7ASLAU8q/qo2HT9dKH/SP2Iiw/PhqqDmpB616gAOOnpMSLiZPO9nB54V7
0QmfXpNuxKfj14JSfBlu2XF+YVffheD50WhUQB0+nhlPiOZgohcFR/Vk07eePokS
Looq3EAFV2ipjnQpo1lyCpkiUQTpxt6JBL4hfLiqdJQx6mbGrSH6uaT56wxCAX31
VDmrTGbh7SGh9W9QCXiODJSl1xcUMOJItBTP84HRjBg24DL4DQM2JGox5u6T+n0a
IzrOpDTI3/hk3gOHiYJKneMs/qOeIGvJW/entvBWr8dIvXP190jIOexZyWzeQH7N
9FcVFUfzlWbpL8KL1v5IqXbEAiiBSY+PAp0ByQ8Nf099Pwd/YLYSgjhYvzsDBQBB
YCiLjhkkm2g/9tdcIGxxfbvJB2p8YOcJSPx4YObMr/CYKIOrkC4NLEKH/ClPagPK
6+G7pYU4xp99eycUGIn3yphn74oa6ABScoZL4z2SvJJx23uL6WwAVxdiX2DoQj7l
JZSx7r6/0lti5zfpSEE3k7eEZP8XP7D3NyIVl/Zekp8fkREPl7G8aOc9G4hpSIWD
O1v8Pwi2HtfDvcKBcGP2XrNt/pcUl4w42FcrrYhE7o0Pybw5tWTlcGsDiqdxbsgM
UfmAlvuIS3ekj6juzgdnC2r4kHuvEolbzJO+lj607LXbaod3Cgzo3zS1TyyYLI4P
+M3xrY9XR1A4p9JU9WHURYrniK3E6SpEf5MPBGYtyOHgOXOf1DHLyfgbjki9w1Ww
YCB+E/OMqKTNo6IbpZqmiCkm5eekw/C+I+e/OvlxVUFymGNNEOKbtyyklQm1xeMn
Ru0OJYJQm+pfYpi3fouzaEvKXQGiODLcotQs+WMFyQlGRyN/sUjQEyD8yudQCjiV
WH21l4iItZ52Wn68xZp/FZcQS+1xRYxeXOzij+gG2/wpOPNQWglDglJVA75G28n/
fUiJMd1NQYtYe9ml0c39YjPQZeI4jAn6JbUccOjkAbSBUtyZeMsySvI685JC/78o
DaXNQIHtR8MTsBbXRXEYU+aP/aPDJ+7SHuVxsWRHfIudJ+j4T7zCbKXfwkA7wzMP
KqwqNCA8RQ9eiPyRo8ibmony9Xy+RP3Ch39EYxM0ATxh/1dS45ljT9wHbzXfHqOl
k+sIhdyHst4wN7pYxCqZMyV8wsfYZgduDLzOQiokX0UCusDp1xResdjPuSrrHima
v/KV9R2gl+66F5cG8FqJ/zWN+kkGMWiUtCFlWDYRXZpBwXvx90ZpDuSCCPiF8a95
1mJ+6OyrfYPoMe4RfdFsjs7LelgXxnXiCZ7A1WRah+vZBhezl4LtPHae2RtPFaRn
eVk2nK+qBNl2t7L03YAMvtCWJ5HLVmfC56KYLm0PIqJFog7jOYvSropPE3hK44ib
xe2+eKafE7U1DHOQ+15Kzpdf7sslA8iF3+AZgH3xKiVuyY/hEX7ZjkyTZrvuLZ2f
AKL01yTt1nU1ddoInwkEwpwp0PC9X4SVtMLRNVyfjQHGv+LnPl5UADkefJDSQ8rV
auFd9UPGU72lYw2fVKyivH4n40O2+PWLgusbo6CIfa5kkbT6esxCQPOBTS4OZEDh
6XDTWbh3JW4WvezzZGClfb1Hz9WcWP0HeXs7ed7NC1gmsqOmIqAav2yiU4VM/DMJ
UnumFoW4PZEutrOsB8CERGmlZAfyxfaTUroVRDUuIEPGXSGZjDwAA4t+RgcaIUAK
GZdIlq30n3q30GDWMp425L++N9ch/H01mrjliyhJhp1TXlwRsXS8V8N+qZTZNa4N
ocufMrLzgkApsF+ThdidB/rSxolTupoYndkWf5ZaXqyPWHHEoNrWxqLxsCfKQDKH
GQN2HproczzbnhVBM4KfKBfasWNtkhFyTFuzttN8PtkrDdr6RlPcBkUtJxysTDYm
FR5UneAeNXt6goUOEJCj84heMNjU3z6UiROXoPwJv9vsedDjikm0upKdejK4CbMg
25mVC7Qxvg+z7sIz8ur/n7oYsDQy1pIHdQ5xptrdAcNwuW+p/1/MSqmoel5dOCPG
d2ByO6nkvoQn6Cui1Z1nVrf14uQEJ4yAnrDxz71raQStvAPjeT4/isKuSHjYcUeP
Bs4iMlj3hgp4L7+S1FIFPWZc7WTv93X4joGP9uKap2j+ZzNxBUhw0gEBtWf7pe7n
ZfxkvOKEJ6Wo7kM3zIOw4g9ygz9P37FRQPwIsCcviOLEQcFH4fI0i/jSVC1wFB3c
+Rw64UTROsiXpk5ojcGkPqj/yUJyC74TTc9Oe5dgtMBImZgr3f/mNgkFu3vpWklj
9pIo8zp9PGpn2pV+svszdkSpuUMR/7/YRLwcEJ3wMN3okwraWO6BMYohX8KDBQb0
yxq5l1AUt6WLYSvobpJXaLGbslXpXtR8NNSCujHZs4S18RaT3Iqqozd4HhoVygiz
ylVC754+/AoFy3JNf96F7rEwlb5D5tdHHcI7ZM/XkOqtPs0qerBVYJI9SPFxlfRi
b//yH2IPCHrBrxOtcI+tiRCtfHsCJ+u4E+/i01SreWFl3tbMqP8ulVtxNZLBYqMs
cF5U8HrCAUAQ5f6Ff87MTVCsudlQTndVSr5BuEE7od9CnSrbHnwO1dWTaYwn0HTS
RfwAGQitp4ctHzG2b9Ju+LTtgmrpEDcbDZGdFk4LpKR4Gkt2SXvPV6DEXWj2vXfQ
1oKHbZ8N54tGK4eJAlWaKWc/iwKw3psz6OByvXyMcjcT2CMirW9xwFP4Jmoj8CKS
kx1eS+pXBLwanhFVuOaKby6COm2kBClgWZBmTY5UhiYEku1yY7G3vVgw2yDKEj4c
OCV4zH3rPfl1LCPEp8F5DjdZm1wBsb8AnhVsRGUhiwEZHgU8Qw7ZsGLTPmpz9VS4
0Lfxca4cEiR1KiNacHVfGwgqJKlPfsbDNjbzbpuP5Kr7CNEjvtc5AA3HCnkFeVLA
DPIJ7vmNqL9uepcA1a4EfURRvlRz42azrzivkjtjETyi4kjU/A4Vz8WM7ZCbMOVn
lZNZW5uZqnSCDo1ZGHXyTYRppdY8xl6OmXfqpPPAKvr0uyhvNXc/g9Y/1909kwEe
kDaJ5iGqdf/vDvfGbxzGHFdeRuBNM4G2KA36W0Un+scp/1GWXJHvSMYGSr3Yz6Sv
k1x6SRlbywNbw785ZKd0phdW0KaTmZpgBbLZ6vSNUeI0O7fv8mPkoiUykkerBtky
EOYgKhbliT53sj+GYpHP47AyEVxUA0f05yMBhJDcVSItioJYxnt6qR2QlHP3dgBc
UfjDjncxSnKQo2+TaadwXt87Kjd4ASUJ77fY7FRwUGDWC//Wfv17TbA47bCQzWUu
zyks0YNU7VT74hZLtjcdfPtQCf8w3Af1qZ8WIlZnZpDWn/qVpXOmCqeg2T8QaPLc
MNiLQzVwiwmQ+adZpHIce+GuHhuQtR5c8oWgB8bSa5/44rukAIhG1Jng8mgwol5J
/yhhQcRwl+S/Zk0xRubzBHxSp2+cF4f/XKm+Kh1BT7//A51Qyt0UOz7sXokjkNfA
vZAsLYNkNJBuepaGeNbM49dyLj+TduFGc7yh6hC928AkCg8DUUMo9TB9DSXsTWJw
WZ40QnSoOFyy+9iHK7vdc1WsYDloYEk+tCK3JTsjjfvuXlhgKvz0fzAyvwEB3PD9
qs1oSrlhAy0t2/+3dUp/ZR3DKWkq+5tXn48BBfOgLhFWqQPHZPGW3Y6N09qOcFQv
wV4cSsOs5m1WQTW63VQ39m/dAbn2veggBxdVLRw5KTvbEQHlZspYV5upyohMLh6I
c3FgSTmoxl9cO2kglH7cGJdWEWx7tfG1x5NjotO+fA5ZbmGXmx9j9cW1KFBdxq20
pMmaGGejQ6Os+iCXlipQ2wNyOLFlZAxj3BpVLiY/nPXAtcA9NS6y8P04vBO98Gxp
E/Gr+gDlYnAxfrZQyOuJus5INQ6S+8A0O/qQ1Q8cMxuL+W0T3mdLVJjNm2mS1DVE
Tx64jbKcoKYHP2QIU2IAqLLb26d1VNmSYv1wTmvKw3GW6RBiB+DpE64DQd2fJ99V
kNqW3lG7PMp8dl7DlliYGHEo8ziQNSYHMx5RbqyiRxwpkCFMVR3O/k7Qf4FHCI4l
SK1SuDAO1tmCnmDcfS7luK1a50xAtbSVBPTE+9zqYMXf/XXPjBmjuyJdhUcW+XA+
iD87vT+aoIE1nk+OMZv1O2SoNu50LOv8zvSu9V1KPzsZkoGuvrEvVT9Ofz7g8uzT
ROJOxr/s9623ICne3+AeudqB0E5tPP3XoyhS087EU01q7skszw8sUA+wumbHARA2
Gr+D7+Kj/JCoA/DkK2oXsue/MjsvQra5YWhdO/hb5xHMOVKn1d5/3m6rkJM1iYAu
v8AhkkXDYU6Y2dOrgJltISNxNnmvhYTdlKedIgmicsZQGVFK0d89xL3Zg8K5CCCH
8ra6cO07WdtmTzfU4JA77AyYNfSohP7nbugBSwWw1Wv1+8r0jg/9NuYr68eLtFQE
kBy6T+VbgLy1NUlMs4dwNLZaZLTXqiYdqV+KIenOEMpImapNYJvFrBwJoip/mmCG
XlI7lRaPa4sv7lt44crVUWT5I9CDoZ8j1gzomXhBzZcpqZp6ZRn4rbH+dyYmjBQH
l+ThC7hipRemw5UjcPv9wMW1R0hJqBttq39QvOlpKNRjcVZ5puFoE5MRNL9QJqlg
ku/G79BgEEpTP3xPoxxpinkIKVCZrcrwPAVMX3lbKxkbR/bEy6mMecW1nGPi5Uy6
ozzkgoyWKZypq7lZLjbzT81PSAk0OJ54IWnpDpRg4TY0dC4ujO4yyzXguhUeQxHe
LdTkG1I/NsmfLAQ7e/sFIoq7dBk66cwVCBwwfqBwG/xuF4QlAn/UFPj4E8UefqIH
D9FDDUCVraz0o1cachK0TF51eGrwG/iHaZb/6Qes182LzEiQUj35hR4s2nXnAcEM
sqDutAD/G0g+jwfVCC3OduS1iQZTwuMoipBlkYPYONqJ5Dt6pBOctGUj1u92s5ZK
BTr+fIFtETtSwVjlT6mEsVOZeesUEvP4o4Gy93raowWq3c0aWN9UliIWeok0h0x7
vTtpG/z5hgtCaLlvCBR+BeyJ/s22zXtQT2/TziWh1/MeK+5LK7JKQtIXp1IK+FcH
oJePEJzEm5gY7NQx5F41wvcH4LUlXHTujBHjxEptCSIGAPP7soXm2OkGWRR/gTka
QbstdMKe0Pa44umMLF4FJCizxIB03Xkk5eQ162fDtwemsI0PgGmf3wtkb8fn2Jy1
3l294NPv46T2o8jHe4mOoN+plL1UDs9arCfgMMkv0T5clRsRlaksM8fl6+PPzmWZ
0+c6+IrpTzZjoU720O5iEbQzyX34gCwE9yf/jL7U418ltRVmR73Vl35H6IhF5Ic7
hzsHs+2pG2Tm004IVPE+R8JjeNemHYynbPQCKBw231eg3/ub0LnUi4iqYyHAbykG
q5YBITUG2JSmh8ymz4urGOky8nJnsq+8im1Nd4QkYAI/a9a89f6yvwhZIUJRe1DF
1fe3s7Maz3xI9IjfHK5inggYp1/wu209E1XSLWzQZwA09dPY7B0ng+dpcnEC7nSS
Dsj/v59vTZdnr+98uuWAvj3bfMSXgr2yjVljCOvsS0/4SuFh/hOuR6W+xUclh9PZ
V+kZlKJWiNK4NhrVDeLLBskqpJLejDTNxOzo4OFUaY4dEnv+BnFReT1z1oSr7P7i
EEXJqFEBPEFOM88yyYg2TesUwYVVV4DxhlWdNB36cTm/p10n8A/lYv50T6jXLJ+t
JkSW1cE24gE7gWkiGGmbUeM7WOVZDKmEQ1MLjP665cDWel4m6RcUrAJA+0TZQWad
+bvpSyu1e5aL6dT4fWfEeGKnaERxHBvMctpf842yw7hXOwFYB4xuiYibBRBTEw7J
8LRynzQF3ME/4O74E4klQZ0M9MyHqzTRHR5vzYYAuSm5TMC7K/O6+DWMr3/wENN9
MejD0MlsHoVXk1z7GvezAJ4fUBo2IhCG7sFm4K36gSJl7UzapXJb8Yrr42zGr+LL
83i+GYypF+UU2mkb3TNHSyuJH+oem5nGA3IgvcluSWQ9P/BvbjMpV7SwTJyh+32k
RDjPa/M4GJn+hotsMsu3fhGQPdbXxNU/BzOqYynU5wwhKOgrw49o13YU7zct2+om
saDaKZHrLdIMa0CtBvEI7FvbRI07LM9H/tnil1/0EIRY5KPi7CU4L6InxcBnOUey
UOEThOXRtc1kaLjDphs1Wswa3Xwk8dK3Ls5Ps5A828w2yKyxntuVjfJwyoITvynq
dAQJNPJwxonbSt7JhVD1DKVJBuGrjMRJfcmerkkmSHoxgC9eiaU7l5qjs19xTR6n
dXs6tSTPXVZf+VG1eqR1V0n5jwvpiAdA8a7qfiV5TCpYBaQYRhjkcnSZQrrKkBpa
rWtzcq1Zt2HXDq4/IEOol98qbHmyXR1nNz8/ey4RK5z5UVW0+UKGivSHtsVs5857
CVuaQIPYHP/DsBCU6mR5OMDZ9ZKKyNxYw6h1Dbe8EW/0eIIQ9bzZfthI3DQFk+9/
EPfG/5qMfBL0vYwyw5e/kr5BmD8djNXFCvx22b0NP+wTU/W8PtJ1QEMQ8mIhbVR8
gDCUSqvVHRNrOrA97hHunvZH6aQI6YqJqzAhX7HFosm6y9jL3nKUQ0Zl00/JPwDJ
hQoKoFaBM5J+w0l2+uzS9cp7t8dkFBTiLruPjLMCkP2ndRFzeHfujz4ZKPW0M5v/
bPfX3wBdG/rbrU2njzE0Sp6+dMSDhn6YXM+G42K4Rz8+mvJfJFheGthrS2FoLIFb
RaJTwgPRpyJPgjJcsLnOqOibMrEOeOb97zCQ6tjNAPr1R4OpdSd4oeiCGD/tEQke
iXDOa10u2TdQwPjKW1c9zaOOpYGby+omRgcRpLtYU3zMOGE+cEhJkmk4K0RUeaCJ
m8AiKpiv4FEOv0hWH8yAqMBfa64JH26SUZvsDwYnzPc5ZlMAlAxZT6tnRNOls2Az
/MiKbahnyrkiTOn7/tQjg/dNuGuOXtxnUWDcCFT0u0wS+k1MKAyS5IKdSvcCAifi
PFFGBi0SCyceeo9iI04c1IMiVSCkKUy3yE31JdqRuHn4hfMF9/kmiefw96H1eB0J
YYUv2LMSFf4nNBWg44iqitd2uKo26yvnbwG8nXoXLdHHSFk3nyDXUKYphXmGwRWf
ACTN1h1nLc98mjYI/krPQUzP17QrKJn1BvEZ3dMrpPT71irhOGXwmtM7fd7H5Vor
6bszmK/Ay/GppU1TmnTo02P76PNrWBj1PyfT4L9B4pJX8I+DDqTKLvEeq2W9dWRB
WnGD+Gkv09kIWGs6Hase7ktKlnI5e1CO06GASX0ZMINlH5JiJOXbZmfHSW4hIaak
8U+3Ijooa7WBZ/4I8eYmwyxDB2ENux1blIQYIwkM+bjyvoLGRl0eQnlItXm5E5ye
bD1zFThBJyMxJDNTk85svuSeBhl9rsx9BFuaHUT6NZGOw2kRMj7hTMHzAzXvEDXu
D5Qi6d789yrenzy5MTO18yt3AlHNkMxR46FZ4lyMHAOi8JZCJ/0AhvpmzIzALIOE
3uNOeLcGNS/6COoX2zoesXw0lIoVjYCp7a96n5pEA44gfScA30qHJO+hO14afwOA
LPBu3gxzDrqcOyupYFfW2KwNhxgmiXWt79Ku/aHaG88KezQqUR3jfXHVz7YpWlaN
Qj1bJcW9RaAbqJ5AYVcJQjziczKLEscd1c1TUyqrptPHVY7WXmVHs85BmLf0wmje
PXHrx32P8gbzX45wFrte5yLL5kAmNSCP1XeBYQRYgg1Pmv+QCFvDarwS44h9iPSD
JeuRYcdomoZUhoEs6ZmNYSaFbk7ktFFTwF8YOexXTh1F7mbL8cmeKNsNFo79x21E
bJ82+pkZqK+muzFXZEjpzZ+qLGeKURTJRi9lVK6B3U1q569lY/Sg8ME3DYuaVz+l
UtpAw8JFbKG/36aBgQlkU1QRMLt5wjz5hgqCodlVOp8zvpCKVt1ZNocq3NMo4P8L
VW7g3pmbvQ++0eA5Vuf1F8631fMgL+oKYALqOaHuvGFhe0IvUrPD6M0vdyMQDVTa
Pf7jiZ7UT1QmOv5f1lTXt/gp+rn4hByiAkNnlHR7Lzj1RhMk1hz4H+cM7kArYPGR
sMiIg9KHx4CWzJIeN7tk5pDmdZNcmIL8FXnTc4mBXN7AdeZKpSBALI13L4ESSa+x
jXiYp5Tp0WrogpX3G/X4r0c27/YMJMiTU+OMMdAnyX+XUkwT97L1+OuSoHQBLa7n
t9Adh6bHmNVKzAfCk3yrxPHIc6p8vG6qRy8D30HpHwC9X8gG1GUKT701NTkKckKd
97/ycOJWKnEe4yjuuilx60pRtOgRVYd/XBje/XsI/TMbndhmroV91xnWe/PCq2v/
eQUow3Z1CzNP0ixEzC4yhWmlgTRK1Q7O2y+wajqCH0IwJXeLP0Q1Zn/Nftr9sv4N
Nnpomgv+G4GGL2b9R6K2Z6JNG5XEAKhApLH4OMjYY3xYkI63Gk3ZPvsYuEzWwikk
TJCEKr121ieGbShEo7Mcv6uKxcPnN/pTF/llwfpDZe83EhO2bBeUGpiraZUs6KF6
/MnL2qjaFlz7SQcstUTTjChlkTi2VTf2rQA47rpSLjxuvFR26JlR/PkbZZ8KwPxI
8GQUrw2+1+teeNCI+/gpx6cf4Vxpjup8dqSQnY3YVEygdgBbSBMzQiZFnHaJZpVV
my+g0EdLn2Xk3lBlAOTD4llZe3MWlu8uHeHREX1Q3xIc723G/wMUc3Sdlvlsv2uD
meMKxqFfuHj78yZ9kii5mgkF8g8hPbfWoF8EV7pMGTfgSBOe7a+L07KmA0Tth0nn
wOeKf9ou55RmJ0DXNM85Z61+Qb8wx6sQv2sWlLCJrfeEuDhSMkaEytA74QMqDOyq
/hVbrCMal2b2Vm+AgeQkTbUFmfTI6aNgmjNBf4XFWv5jNUc1sIduWiaK+JIFk8lQ
ofDaoeb8MTIBgUYMwKmMABsMJeMksTXHVPGkKp4I32tEb0fd1eKx1xqDKX6b7cTE
hLbrfJW8PUxuAlH7GlYiigT6hy1FDD9OXkKTwx3Dj9A6330yJwq0sd9C1zZhIRXn
Mww57IFo8+YpKQsd3vV/r8uNTFkpuN3+MiSpWigaAS6fHiOHyD++xSxE95vw5uq1
0VVD5I0GX8zpn/Ue7/nxSZgDOALCc7ANqBsvn0aJhzp95cB3OYR+eMYs6LIReWT+
jjuF/FmwVVDFXIPabhGoBwUjQ+FyKEPU6QTvax6sOl4TbWaj+4y2nG40Sv9cQNVc
83hOZm3uKaAIdZwAhZrrFNg9HdcpN1GCGkC+N0S8UUOkM7sykWgu7mR2eSb6KB0Y
bxatdkudIdHSlb88RlnorzzInm5Uts6615ZsZMowC6O/qAvZGAtws4DDARIjVMQ7
BrKjvtLCRWYAwBsMwnyBPaCMY3e2RkGfSBxg2n6cSVk4jmlP69tjJlbQdcZKHLc3
mrnqM+fxx86/wRfPMiKajZcvccMWSv3rB9jQAPSdYJRrml5nYUwqT4z6dLcMum3j
si/uP7gSZh56q7gxSlM4MdL6cIgHlUjdEjXz4XACsQjp6H8Ya87fy+WncgKIEgZ8
lqhurytStNIJTNazbj9DKwtlKbmXQQtIUd6oPxDjjugEe1K0PCDhq8/z7bqe+MaA
TjXWv0Ngv6CwNanNevuTEEc8LSmzAV4C0pJcFl4pgW3FbrWrRIzatAMfVopdyf8x
QYC6AqxxkeIUNMkA1onG5P4/cnwbvwXGi4nN7lEVLgLf3vEP/YzrNKkUP0N9r32f
1LinCiZEhNgDazZmNrEY583wnE5ZnCo7e2i08CSwE88NDMT1naiDAlaeQ5/q5JIA
Q/Fl0ejGjePr59qydTBDKOzNsb/PUJwMGdH19HK3mfV0NxS53BnVcumQuApSnncS
Ltkpe/0b0d+EZbTFwNoAkdOB+tlC2wVl/J8tZSK1O5P6TaAHhmklxNpS+o0kMQDf
V1yv/ry+kMrIfAMvvTRhjTlwEHDXNLoXkp7V88E6HuCyiHfGbB6natOkxGUaioUN
dRvHte3Qcb3EFyOac8grvd/S6OeD+qZ9tKiD0uyewrnJq4hhfKKUfky059P1S/CW
5eb7rF/kHufslQJC9JeY47tJbDAq+qBemzVIPkjG6WkqhM+uTCPIH0ALCLhafjrt
kJKQTU1qJwhpOOjnZpDPFHGSgds+fl8aasLl28S6QGpbuaBTmnf78uCCKcTzVS3L
r2xvrgSfiBTZuBPFBp9xvNOXPM6C5XjFOzQZD/LndAz5KsiP99wV0iERbZns+3Zr
V5xW4gP61Ryb+8M6okqS7jqg0BTT1K9nJB7AU/tk36Wkx9iXc0swoxN0QXjuu/aG
+VUMVQmKUl6noqNEAmRyERhZRy3BCVvagMqtAbFuF7I3s2v9RlpWO9qJKxLC0n0f
GFLVWH4/8lCGuaSedqSXSsNMwp2J4CUL/5bubG/6q3c2Kg9cdOSPTcFbtJOlpeo7
HkkE2yimoDebvyhW+oZb5lIfYPlV8EYGmohe1Ngp77q9aU3fi4gNqrnGyNUOq2e8
sRJSZ+cihnnAqYTzPzkORJirQsMlJlzQLcW2xNgyOGstw+FrSYWuAhFUDVnB7ewS
1sX2Vp9nYN8b8aK8PhTNsKkqwRjSNZmqeA64jLdQaoqyqIuu/bxPXrw1DrnaOKcX
NWJIArErb4bD+CEMBet4qu7O5NFdYTsOZWLTMV3knBF5pDroiN6RxAcpwOeFKVMp
LzHKdwl57PJWwgHjbL5SNHvgMauyRfeguwIQgwo1GEQ2sDUnPnO7Ap7zkmSayfsO
opA7HXRMVEPncqmismZoR5yADtBN7lnHXCZ522UjKxMzOPSKuLjbknLm1T/NLG6S
UbzAAlA1nO2o1eypzjLxbyVQ0g/Buzjup52gb8aV03hFh2WuqPs63Jyk/aaOpAzG
lXJ5rz2Vpp1oYlicLbHmG/eBlqpVwFoViF2b96SOsf2/xpBuGfcluFqOqpUyXzOd
lNJN92KOSzhsl42KFR80rcL6Rn6J9EdfSejOb+5X1537m9UwCoRNwVUU8XRtxQWZ
ktJ6rTZMbqP42lwD5I9zj6hgJgrC5eS9hxbY2kxD+S2oJrFv3JNdjHORqOt2Imfo
lTXNTrGXwlu23ivrSm7/O4VTePiH6lZlVC1OCNPUXrFPSuLLqtdWUPpQcYGez+Zk
f8vEEHzbyKqbsv29j0SxCmG5GE5lAoUvicTXAaAXW7s3uSDuJlpaZDfatkGLClq+
pAF9J1/fRHqvqtxvfghAhVocyi/+BN1NSItJxrcMWql62fgkTGU3C+HNIv9/ynWO
elfW8j6BbpqXhwLMX9NFJfkZQRnH7OKzQ39WiVXXjy5pTLrQQNjvmKKcOQg+XBxX
lOZ/Aam/XV2DB5Y8wgPqbe6WVF8aJn64fw7GrdmrDpPHsGoXwTCXHERB7OKH6iXL
CPjXUzqevsUmmlsRPllCKNV1LS6vdWSO0iWkoMVKzZgKQSRbbxpQ7j1m2uktL+zV
vAKu3cktBCfK1n5XQ3pcCbhvcE6JYsdUy8H+S4ZfPqGWFj8pRoW6ab1t1iq096a9
8TAh5wo8hvUo5LVluJBLi6Mqoad9BsrcGEU2JvEnXpWUZ8YLZsVA/smNXiyw6Mm2
BroYt6kteaqHAvDL7chEEuu0qi63k4EXI0bIAE2x6Wo2kHLGE0VtX9AV1kIV4WIi
VKOjHz0EnNcqvsXejiBJcHAEdJwaUrwXmZQB7ze7xmAPQ5Gs4q6VoNavqL/r7N1Q
m0RCETmUxIZe0l1AC/Ua/Osu9FmKfk/DW3KtCDh/BKObOVIS4F1THydmDLdddIxU
FjJgtSxUf/CVM4WsTRuADtADCDNZCxvHZ6CUTy/yobf5sKFREIkpQxHajNsmO5th
g0GfRSzcoyWWCd2L1zCRyAsZdu5BpGS2/OwarDFlFd7MWpqabkEsA6ijG6ncp8/J
FuRHxqH2ySVBXY7l/SAuhY8/Y2I1Fcw+lsAdkmftBy2wwzkEwYhF+FoZuxRPebpo
HLeqjOjyTwH2s+SKgFg+yi+M2MrlnUuSIQL45eIwhtzenb4FzUBj5QhPniZpd5ez
KKsyrWsE498eWzpBCOVXcdjI+4uvlkR7X5KAkSe1qLom4lhAWTtOHmUHNrSP5G0x
z0+MsP7AipprnviuU6ScKkFmR37IwbXBNu9VYD6hlPoVnEf9HIr4ezMgJmuDxBGZ
a/rUgCmoJ96nG0LDDT2NkkN0ulzXHyrq6fMpZQJcExR3sb35qTfJDGRCfkuy/FAo
dcpyEfBtGhY0bguW7sMYHDjjHeAql5OUPgANlkpFo+KDxY9jdm7Q614thPTuAJHE
2T5nOINYazfF2G9KOltJQYRfDidshdnYpuEp/NAuiuWgpPjrtNF7OEWWHJCI4euU
aSwM8AiKoK590HjQT2By+SFRtoeBbu51wnPWGS9nElG/TwTyOmU+6ELH8YThF9ox
p4gT9on/Z/hQEg5teoZwWL1Gcx4drUKsXqeuJvZv8DJpeHFrOWLAT1ITdRTSBTuc
LIAeAfnOEZKDu2E6Z41pGr5nOdPY3ZgthLIBOSFD5WAEcFUI8ZbP/3ioUW7+jwKE
+s/eU0RwP5XsVaJBc2/2ebZMUkoOo1cSDfPpjZb18+m69GfmXnv5ygKNFrgh+jo/
gC0nhd4qdGViBuupKINwATv5b7cr+5Z2Z/8gVdoyaCR/VfH0RCIbO8dVynOthxS8
oqB/eagDAhVusx/7bTPCsZForhLzjvhoFgM53Wr95pVSruq6fGkZoh9mxVP5wNI2
HqmEM1KniRtz/NbuuZPYykhvZI+uyvPN7Jn6IMWFj+Td8NPp6GOQpMi1HuCvIG41
WZPles2ofuHeOZB81RJPlWt41AKkn21/M06xeLikcevO76q0wHeGCRsc4u272r4e
pFMgldxHtNa80K+co/sK11fRbzpNUW5Dq+NlhmrGMOiZcsdo6ZIfRApwgWzZcjvl
PXo2muB1LRlbEuU47yLjTA5k0/xDK4R6MvWUVgcXDxdQ5X2ezCV/iX3PbEL5g8Xk
IJdfNjC31q/xJNDF5070aHoLPggyr1hq73XHi7duArp8/ki2B7Z1NIrPWYpXx7b8
QWoUR57QHyYwNsfW40MmOm6+qpX20XOVmnZMNVlS8yuOWl9QFgRakKHXn5Mw94Qd
6EPu6m/cv84l7CyfCsi0ZdtYrH4I1bgKRre8QjW7GOTvTs8mB8m+NXO+TxixHwgO
Wqmtu9L3KlmL2O3+4AxWwLi9xnuzse+0fT1w5l1PRHQ/wj3BFJ3RlWZ+lQlnNQEG
Dp9VB345j7evivNlv2Ss8iDpXIHIAnT/VVewfLsIqd6SnlR4hIGIdfcRLe0uzDAl
JGvU15u76i3jIkcw6lNfU/+epA0kHnHNBA4BBhn8qmP9y8UXFVlJbNdEBMl8OOfY
ZYKizrJl9LDq1hleLPJt5D6Ix087paeMbJrBwa+G5B1w4WWVr/DzzU1xuR6mbab9
tExw9Eg7GPaz+SsP1bOoN9VzbmjRCWFcBUPUFLpiOXl9ABRGqwv8OmOD40ZHGo9t
9xmohCPbQf1/2W72GwXOJh7MVrlH31h6pH4hiqM9EvwyorxSincafCpJp8VtJJhB
c3NgbGy7L08l5gKsTOLjyfUmSAz8FICujqKnAFMm777romaUfoQMR96rgID3PSRM
qcetky1zVD4pzdz8gI89XJy5MBJk44iQSn3/l3rYQP9ZiQHRw2Tkg1SoI8K/wdzx
x85KRbOEt6GJjEcJdePrxo+UH6Ci1zJhx423f6mWnHwxdhz8SdOg1sF7I3TvtXW9
Ep7En6P2fg3/hdj85SyS8eoh9qP/lMamB2j98upthFERTBm3Kzw7kAKo6iaCtMV6
UoHiqmbtjwHpvir0UY3h0CoR0CDeZCvev7yZPc/NKIN2PaqqbF0fMWkO/VySHS2u
xmw4uQtShXL7ejKd3g1QwoXCK+APOGLPa8cvvNBMtBX9ozrby2xyhWSevyAETUvw
I0lx26mSO9uMthcIOEh2Rh7hZA27S7UlpoBtXkw0ZqmrpFyjNrQI0I8ICX+yXXug
4yq+UApHzQ4t+h+Gcbc93w4EnicOXk2mKqEsVtmB7jXj3APqvrUIt3auUM4r4T2A
Hwd6vjzYLNCBPOoG+aYLg0q3lANZxkinSGgAW6SymVv+mLreL3yfREqikctu3ZEN
H/xTf+iQMJlCntG01Lil6E6KX1rwewMIl8NLZPtTqXGDxKcTn/G44iKQKx4+a7p0
11wZUKEpn/BrUUns0xsfYjYN77kv/w6YxQNNTEfWMIAkpNSrdRmlmUrJtlHE1vIg
oqoYGcIBVOJ18CLbq2yIzDVwy8GaCgZr2b5thWNTBpkzY5MoqHxS3jsm2JtPAxgp
e167LgDVHVf1S4upDlrt0gspx/Cbl+pnqtFNRJzrFLLX8DRi32HF0pmqBGlZ0fzD
NFa+aOfNilSb9ZmTAdTCPBs62OEkOymphmbZHfiOLPvf3WxTHPFEsHrVfLDSz0tz
RNVbQdEr/lPWZf72xw+92uIlk53XGC9U/A1uItYNVO8Fo+shLeF1qgJUFdIsIuJ4
jUgp4ELJPvrn6TjgSTLqcJQx7XICJ4OGx8Y9Sp6QM76E2hoXkjX+66Rl/yzSjdRD
dRZLee247l7ODy2EOzXOUSMOP8dGY+GBuDgp18g2xVj282mPhu6tqsS1bY05x0Iv
DHYa5TSClzalkyAtsUaQh2jROCbB5uwz49KAFLADDeFU/t/iO/94fVHC2NCdfDq0
mN5OXIa8N6BIwtfJMpIP6K+eJnQFzjCTo6TGRyYMLmME42D8n8BfKLOd2Hem/4LB
x7Mu/ATEpOPbSWjFMqs4jBoesAS2VDTRKv7gvmRRSs3SXHtxGpmiBxzXkK1ytttD
myysKbIpjC1P6CNB11f6yUNWPeF2yDAv251TrQWbWx+LH42n5tNxecP9v+V/Ucnr
zaQ8skNL42Kio1q897ouGL+zbnmAF19u1FN6qqYIDGfFWhKGhjpV33oqL2+lpmQM
ZE0uxnkZQvvKZEZkiMsuqBozcjsehePhFcbHByLD9B2HSi9QSJfz+9HViIeqcLIP
K8khhzpayUsfExKji/XY5SgY+erj96Kc9PNkNMQc+qNYagbevH7XIjMwpRzky5kx
DMpUMdme6u9N0laXkB/Xmx3TVTXfrfmAX1nv2ngnqihdgBuDGNnstcm3Z55ERZqw
ClYdmxQ5t/kM5TnQN/s4Bw==
`pragma protect end_protected
