-- pcie_wrap0.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pcie_wrap0 is
	port (
		hip_config_tl_hpg_ctrler         : in  std_logic_vector(4 downto 0)   := (others => '0'); --      hip_config_tl.hpg_ctrler
		hip_config_tl_tl_cfg_add         : out std_logic_vector(3 downto 0);                      --                   .tl_cfg_add
		hip_config_tl_tl_cfg_ctl         : out std_logic_vector(31 downto 0);                     --                   .tl_cfg_ctl
		hip_config_tl_tl_cfg_sts         : out std_logic_vector(52 downto 0);                     --                   .tl_cfg_sts
		hip_config_tl_cpl_err            : in  std_logic_vector(6 downto 0)   := (others => '0'); --                   .cpl_err
		hip_config_tl_cpl_pending        : in  std_logic                      := '0';             --                   .cpl_pending
		hip_coreclkout_hip_clk           : out std_logic;                                         -- hip_coreclkout_hip.clk
		hip_cseb_cseb_rddata             : in  std_logic_vector(31 downto 0)  := (others => '0'); --           hip_cseb.cseb_rddata
		hip_cseb_cseb_rdresponse         : in  std_logic_vector(4 downto 0)   := (others => '0'); --                   .cseb_rdresponse
		hip_cseb_cseb_waitrequest        : in  std_logic                      := '0';             --                   .cseb_waitrequest
		hip_cseb_cseb_wrresponse         : in  std_logic_vector(4 downto 0)   := (others => '0'); --                   .cseb_wrresponse
		hip_cseb_cseb_wrresp_valid       : in  std_logic                      := '0';             --                   .cseb_wrresp_valid
		hip_cseb_cseb_addr               : out std_logic_vector(32 downto 0);                     --                   .cseb_addr
		hip_cseb_cseb_be                 : out std_logic_vector(3 downto 0);                      --                   .cseb_be
		hip_cseb_cseb_rden               : out std_logic;                                         --                   .cseb_rden
		hip_cseb_cseb_wrdata             : out std_logic_vector(31 downto 0);                     --                   .cseb_wrdata
		hip_cseb_cseb_wren               : out std_logic;                                         --                   .cseb_wren
		hip_cseb_cseb_wrresp_req         : out std_logic;                                         --                   .cseb_wrresp_req
		hip_cseb_cseb_rddata_parity      : in  std_logic_vector(3 downto 0)   := (others => '0'); --                   .cseb_rddata_parity
		hip_cseb_cseb_addr_parity        : out std_logic_vector(4 downto 0);                      --                   .cseb_addr_parity
		hip_cseb_cseb_wrdata_parity      : out std_logic_vector(3 downto 0);                      --                   .cseb_wrdata_parity
		hip_ctrl_test_in                 : in  std_logic_vector(31 downto 0)  := (others => '0'); --           hip_ctrl.test_in
		hip_ctrl_simu_mode_pipe          : in  std_logic                      := '0';             --                   .simu_mode_pipe
		hip_hip_status_derr_cor_ext_rcv  : out std_logic;                                         --     hip_hip_status.derr_cor_ext_rcv
		hip_hip_status_derr_cor_ext_rpl  : out std_logic;                                         --                   .derr_cor_ext_rpl
		hip_hip_status_derr_rpl          : out std_logic;                                         --                   .derr_rpl
		hip_hip_status_dlup              : out std_logic;                                         --                   .dlup
		hip_hip_status_dlup_exit         : out std_logic;                                         --                   .dlup_exit
		hip_hip_status_ev128ns           : out std_logic;                                         --                   .ev128ns
		hip_hip_status_ev1us             : out std_logic;                                         --                   .ev1us
		hip_hip_status_hotrst_exit       : out std_logic;                                         --                   .hotrst_exit
		hip_hip_status_int_status        : out std_logic_vector(3 downto 0);                      --                   .int_status
		hip_hip_status_l2_exit           : out std_logic;                                         --                   .l2_exit
		hip_hip_status_lane_act          : out std_logic_vector(3 downto 0);                      --                   .lane_act
		hip_hip_status_ltssmstate        : out std_logic_vector(4 downto 0);                      --                   .ltssmstate
		hip_hip_status_rx_par_err        : out std_logic;                                         --                   .rx_par_err
		hip_hip_status_tx_par_err        : out std_logic_vector(1 downto 0);                      --                   .tx_par_err
		hip_hip_status_cfg_par_err       : out std_logic;                                         --                   .cfg_par_err
		hip_hip_status_ko_cpl_spc_header : out std_logic_vector(7 downto 0);                      --                   .ko_cpl_spc_header
		hip_hip_status_ko_cpl_spc_data   : out std_logic_vector(11 downto 0);                     --                   .ko_cpl_spc_data
		hip_int_msi_app_int_sts          : in  std_logic                      := '0';             --        hip_int_msi.app_int_sts
		hip_int_msi_app_msi_num          : in  std_logic_vector(4 downto 0)   := (others => '0'); --                   .app_msi_num
		hip_int_msi_app_msi_req          : in  std_logic                      := '0';             --                   .app_msi_req
		hip_int_msi_app_msi_tc           : in  std_logic_vector(2 downto 0)   := (others => '0'); --                   .app_msi_tc
		hip_int_msi_app_int_ack          : out std_logic;                                         --                   .app_int_ack
		hip_int_msi_app_msi_ack          : out std_logic;                                         --                   .app_msi_ack
		hip_lmi_lmi_addr                 : in  std_logic_vector(11 downto 0)  := (others => '0'); --            hip_lmi.lmi_addr
		hip_lmi_lmi_din                  : in  std_logic_vector(31 downto 0)  := (others => '0'); --                   .lmi_din
		hip_lmi_lmi_rden                 : in  std_logic                      := '0';             --                   .lmi_rden
		hip_lmi_lmi_wren                 : in  std_logic                      := '0';             --                   .lmi_wren
		hip_lmi_lmi_ack                  : out std_logic;                                         --                   .lmi_ack
		hip_lmi_lmi_dout                 : out std_logic_vector(31 downto 0);                     --                   .lmi_dout
		hip_power_mngt_pm_auxpwr         : in  std_logic                      := '0';             --     hip_power_mngt.pm_auxpwr
		hip_power_mngt_pm_data           : in  std_logic_vector(9 downto 0)   := (others => '0'); --                   .pm_data
		hip_power_mngt_pme_to_cr         : in  std_logic                      := '0';             --                   .pme_to_cr
		hip_power_mngt_pm_event          : in  std_logic                      := '0';             --                   .pm_event
		hip_power_mngt_pme_to_sr         : out std_logic;                                         --                   .pme_to_sr
		hip_rst_reset_status             : out std_logic;                                         --            hip_rst.reset_status
		hip_rst_serdes_pll_locked        : out std_logic;                                         --                   .serdes_pll_locked
		hip_rst_pld_clk_inuse            : out std_logic;                                         --                   .pld_clk_inuse
		hip_rst_pld_core_ready           : in  std_logic                      := '0';             --                   .pld_core_ready
		hip_rst_testin_zero              : out std_logic;                                         --                   .testin_zero
		hip_rx_bar_be_rx_st_bar          : out std_logic_vector(7 downto 0);                      --      hip_rx_bar_be.rx_st_bar
		hip_rx_bar_be_rx_st_mask         : in  std_logic                      := '0';             --                   .rx_st_mask
		hip_rx_st_startofpacket          : out std_logic_vector(0 downto 0);                      --          hip_rx_st.startofpacket
		hip_rx_st_endofpacket            : out std_logic_vector(0 downto 0);                      --                   .endofpacket
		hip_rx_st_error                  : out std_logic_vector(0 downto 0);                      --                   .error
		hip_rx_st_valid                  : out std_logic_vector(0 downto 0);                      --                   .valid
		hip_rx_st_empty                  : out std_logic_vector(1 downto 0);                      --                   .empty
		hip_rx_st_ready                  : in  std_logic                      := '0';             --                   .ready
		hip_rx_st_data                   : out std_logic_vector(255 downto 0);                    --                   .data
		hip_rx_st_parity                 : out std_logic_vector(31 downto 0);                     --                   .parity
		hip_serial_rx_in0                : in  std_logic                      := '0';             --         hip_serial.rx_in0
		hip_serial_rx_in1                : in  std_logic                      := '0';             --                   .rx_in1
		hip_serial_rx_in2                : in  std_logic                      := '0';             --                   .rx_in2
		hip_serial_rx_in3                : in  std_logic                      := '0';             --                   .rx_in3
		hip_serial_rx_in4                : in  std_logic                      := '0';             --                   .rx_in4
		hip_serial_rx_in5                : in  std_logic                      := '0';             --                   .rx_in5
		hip_serial_rx_in6                : in  std_logic                      := '0';             --                   .rx_in6
		hip_serial_rx_in7                : in  std_logic                      := '0';             --                   .rx_in7
		hip_serial_tx_out0               : out std_logic;                                         --                   .tx_out0
		hip_serial_tx_out1               : out std_logic;                                         --                   .tx_out1
		hip_serial_tx_out2               : out std_logic;                                         --                   .tx_out2
		hip_serial_tx_out3               : out std_logic;                                         --                   .tx_out3
		hip_serial_tx_out4               : out std_logic;                                         --                   .tx_out4
		hip_serial_tx_out5               : out std_logic;                                         --                   .tx_out5
		hip_serial_tx_out6               : out std_logic;                                         --                   .tx_out6
		hip_serial_tx_out7               : out std_logic;                                         --                   .tx_out7
		hip_tx_cred_tx_cred_datafccp     : out std_logic_vector(11 downto 0);                     --        hip_tx_cred.tx_cred_datafccp
		hip_tx_cred_tx_cred_datafcnp     : out std_logic_vector(11 downto 0);                     --                   .tx_cred_datafcnp
		hip_tx_cred_tx_cred_datafcp      : out std_logic_vector(11 downto 0);                     --                   .tx_cred_datafcp
		hip_tx_cred_tx_cred_fchipcons    : out std_logic_vector(5 downto 0);                      --                   .tx_cred_fchipcons
		hip_tx_cred_tx_cred_fcinfinite   : out std_logic_vector(5 downto 0);                      --                   .tx_cred_fcinfinite
		hip_tx_cred_tx_cred_hdrfccp      : out std_logic_vector(7 downto 0);                      --                   .tx_cred_hdrfccp
		hip_tx_cred_tx_cred_hdrfcnp      : out std_logic_vector(7 downto 0);                      --                   .tx_cred_hdrfcnp
		hip_tx_cred_tx_cred_hdrfcp       : out std_logic_vector(7 downto 0);                      --                   .tx_cred_hdrfcp
		hip_tx_st_startofpacket          : in  std_logic_vector(0 downto 0)   := (others => '0'); --          hip_tx_st.startofpacket
		hip_tx_st_endofpacket            : in  std_logic_vector(0 downto 0)   := (others => '0'); --                   .endofpacket
		hip_tx_st_error                  : in  std_logic_vector(0 downto 0)   := (others => '0'); --                   .error
		hip_tx_st_valid                  : in  std_logic_vector(0 downto 0)   := (others => '0'); --                   .valid
		hip_tx_st_empty                  : in  std_logic_vector(1 downto 0)   := (others => '0'); --                   .empty
		hip_tx_st_ready                  : out std_logic;                                         --                   .ready
		hip_tx_st_data                   : in  std_logic_vector(255 downto 0) := (others => '0'); --                   .data
		hip_tx_st_parity                 : in  std_logic_vector(31 downto 0)  := (others => '0'); --                   .parity
		local_pcie_perstn_reset_n        : in  std_logic                      := '0';             --  local_pcie_perstn.reset_n
		nc_reset_reset_n                 : in  std_logic                      := '0';             --           nc_reset.reset_n
		pcie_ref_clk_clk                 : in  std_logic                      := '0';             --       pcie_ref_clk.clk
		pcie_rstn_npor                   : in  std_logic                      := '0';             --          pcie_rstn.npor
		pcie_rstn_pin_perst              : in  std_logic                      := '0';             --                   .pin_perst
		pld_clk_clk                      : in  std_logic                      := '0';             --            pld_clk.clk
		rcd_hip_status_derr_cor_ext_rcv  : in  std_logic                      := '0';             --     rcd_hip_status.derr_cor_ext_rcv
		rcd_hip_status_derr_cor_ext_rpl  : in  std_logic                      := '0';             --                   .derr_cor_ext_rpl
		rcd_hip_status_derr_rpl          : in  std_logic                      := '0';             --                   .derr_rpl
		rcd_hip_status_dlup_exit         : in  std_logic                      := '0';             --                   .dlup_exit
		rcd_hip_status_ev128ns           : in  std_logic                      := '0';             --                   .ev128ns
		rcd_hip_status_ev1us             : in  std_logic                      := '0';             --                   .ev1us
		rcd_hip_status_hotrst_exit       : in  std_logic                      := '0';             --                   .hotrst_exit
		rcd_hip_status_int_status        : in  std_logic_vector(3 downto 0)   := (others => '0'); --                   .int_status
		rcd_hip_status_l2_exit           : in  std_logic                      := '0';             --                   .l2_exit
		rcd_hip_status_lane_act          : in  std_logic_vector(3 downto 0)   := (others => '0'); --                   .lane_act
		rcd_hip_status_ltssmstate        : in  std_logic_vector(4 downto 0)   := (others => '0'); --                   .ltssmstate
		rcd_hip_status_dlup              : in  std_logic                      := '0';             --                   .dlup
		rcd_hip_status_rx_par_err        : in  std_logic                      := '0';             --                   .rx_par_err
		rcd_hip_status_tx_par_err        : in  std_logic_vector(1 downto 0)   := (others => '0'); --                   .tx_par_err
		rcd_hip_status_cfg_par_err       : in  std_logic                      := '0';             --                   .cfg_par_err
		rcd_hip_status_ko_cpl_spc_header : in  std_logic_vector(7 downto 0)   := (others => '0'); --                   .ko_cpl_spc_header
		rcd_hip_status_ko_cpl_spc_data   : in  std_logic_vector(11 downto 0)  := (others => '0')  --                   .ko_cpl_spc_data
	);
end entity pcie_wrap0;

architecture rtl of pcie_wrap0 is
	component alt_xcvr_reconfig is
		generic (
			device_family                 : string  := "Stratix V";
			number_of_reconfig_interfaces : integer := 2;
			enable_offset                 : integer := 1;
			enable_lc                     : integer := 1;
			enable_dcd                    : integer := 0;
			enable_dcd_power_up           : integer := 1;
			enable_analog                 : integer := 1;
			enable_eyemon                 : integer := 0;
			enable_ber                    : integer := 0;
			enable_dfe                    : integer := 0;
			enable_adce                   : integer := 0;
			enable_mif                    : integer := 0;
			enable_pll                    : integer := 0
		);
		port (
			reconfig_busy             : out std_logic;                                         -- reconfig_busy
			mgmt_clk_clk              : in  std_logic                      := 'X';             -- clk
			mgmt_rst_reset            : in  std_logic                      := 'X';             -- reset
			reconfig_mgmt_address     : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- address
			reconfig_mgmt_read        : in  std_logic                      := 'X';             -- read
			reconfig_mgmt_readdata    : out std_logic_vector(31 downto 0);                     -- readdata
			reconfig_mgmt_waitrequest : out std_logic;                                         -- waitrequest
			reconfig_mgmt_write       : in  std_logic                      := 'X';             -- write
			reconfig_mgmt_writedata   : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			reconfig_to_xcvr          : out std_logic_vector(769 downto 0);                    -- reconfig_to_xcvr
			reconfig_from_xcvr        : in  std_logic_vector(505 downto 0) := (others => 'X'); -- reconfig_from_xcvr
			tx_cal_busy               : out std_logic;                                         -- tx_cal_busy
			rx_cal_busy               : out std_logic;                                         -- tx_cal_busy
			cal_busy_in               : in  std_logic                      := 'X';             -- cal_busy_in
			reconfig_mif_address      : out std_logic_vector(31 downto 0);                     -- address
			reconfig_mif_read         : out std_logic;                                         -- read
			reconfig_mif_readdata     : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- readdata
			reconfig_mif_waitrequest  : in  std_logic                      := 'X'              -- waitrequest
		);
	end component alt_xcvr_reconfig;

	component altpcie_sv_hip_ast_hwtcl is
		generic (
			ACDS_VERSION_HWTCL                       : string  := "15.1";
			lane_mask_hwtcl                          : string  := "x4";
			gen123_lane_rate_mode_hwtcl              : string  := "Gen1 (2.5 Gbps)";
			port_type_hwtcl                          : string  := "Native endpoint";
			pcie_spec_version_hwtcl                  : string  := "2.1";
			ast_width_hwtcl                          : string  := "Avalon-ST 64-bit";
			pll_refclk_freq_hwtcl                    : string  := "100 MHz";
			set_pld_clk_x1_625MHz_hwtcl              : integer := 0;
			use_ast_parity                           : integer := 0;
			multiple_packets_per_cycle_hwtcl         : integer := 0;
			in_cvp_mode_hwtcl                        : integer := 0;
			use_pci_ext_hwtcl                        : integer := 0;
			use_pcie_ext_hwtcl                       : integer := 0;
			use_config_bypass_hwtcl                  : integer := 0;
			enable_tl_only_sim_hwtcl                 : integer := 0;
			hip_reconfig_hwtcl                       : integer := 0;
			hip_tag_checking_hwtcl                   : integer := 1;
			enable_power_on_rst_pulse_hwtcl          : integer := 0;
			enable_pcisigtest_hwtcl                  : integer := 0;
			bar0_size_mask_hwtcl                     : integer := 28;
			bar0_io_space_hwtcl                      : string  := "Disabled";
			bar0_64bit_mem_space_hwtcl               : string  := "Enabled";
			bar0_prefetchable_hwtcl                  : string  := "Enabled";
			bar1_size_mask_hwtcl                     : integer := 0;
			bar1_io_space_hwtcl                      : string  := "Disabled";
			bar1_prefetchable_hwtcl                  : string  := "Disabled";
			bar2_size_mask_hwtcl                     : integer := 0;
			bar2_io_space_hwtcl                      : string  := "Disabled";
			bar2_64bit_mem_space_hwtcl               : string  := "Disabled";
			bar2_prefetchable_hwtcl                  : string  := "Disabled";
			bar3_size_mask_hwtcl                     : integer := 0;
			bar3_io_space_hwtcl                      : string  := "Disabled";
			bar3_prefetchable_hwtcl                  : string  := "Disabled";
			bar4_size_mask_hwtcl                     : integer := 0;
			bar4_io_space_hwtcl                      : string  := "Disabled";
			bar4_64bit_mem_space_hwtcl               : string  := "Disabled";
			bar4_prefetchable_hwtcl                  : string  := "Disabled";
			bar5_size_mask_hwtcl                     : integer := 0;
			bar5_io_space_hwtcl                      : string  := "Disabled";
			bar5_prefetchable_hwtcl                  : string  := "Disabled";
			expansion_base_address_register_hwtcl    : integer := 0;
			io_window_addr_width_hwtcl               : integer := 0;
			prefetchable_mem_window_addr_width_hwtcl : integer := 0;
			vendor_id_hwtcl                          : integer := 0;
			device_id_hwtcl                          : integer := 1;
			revision_id_hwtcl                        : integer := 1;
			class_code_hwtcl                         : integer := 0;
			subsystem_vendor_id_hwtcl                : integer := 0;
			subsystem_device_id_hwtcl                : integer := 0;
			max_payload_size_hwtcl                   : integer := 128;
			extend_tag_field_hwtcl                   : string  := "32";
			completion_timeout_hwtcl                 : string  := "ABCD";
			enable_completion_timeout_disable_hwtcl  : integer := 1;
			use_aer_hwtcl                            : integer := 0;
			ecrc_check_capable_hwtcl                 : integer := 0;
			ecrc_gen_capable_hwtcl                   : integer := 0;
			use_crc_forwarding_hwtcl                 : integer := 0;
			port_link_number_hwtcl                   : integer := 1;
			dll_active_report_support_hwtcl          : integer := 0;
			surprise_down_error_support_hwtcl        : integer := 0;
			slotclkcfg_hwtcl                         : integer := 1;
			msi_multi_message_capable_hwtcl          : string  := "4";
			msi_64bit_addressing_capable_hwtcl       : string  := "true";
			msi_masking_capable_hwtcl                : string  := "false";
			msi_support_hwtcl                        : string  := "true";
			enable_function_msix_support_hwtcl       : integer := 0;
			msix_table_size_hwtcl                    : integer := 0;
			msix_table_offset_hwtcl                  : string  := "0";
			msix_table_bir_hwtcl                     : integer := 0;
			msix_pba_offset_hwtcl                    : string  := "0";
			msix_pba_bir_hwtcl                       : integer := 0;
			enable_slot_register_hwtcl               : integer := 0;
			slot_power_scale_hwtcl                   : integer := 0;
			slot_power_limit_hwtcl                   : integer := 0;
			slot_number_hwtcl                        : integer := 0;
			endpoint_l0_latency_hwtcl                : integer := 0;
			endpoint_l1_latency_hwtcl                : integer := 0;
			vsec_id_hwtcl                            : integer := 40960;
			user_id_hwtcl                            : integer := 0;
			vsec_rev_hwtcl                           : integer := 0;
			millisecond_cycle_count_hwtcl            : integer := 124250;
			port_width_be_hwtcl                      : integer := 8;
			port_width_data_hwtcl                    : integer := 64;
			gen3_dcbal_en_hwtcl                      : integer := 1;
			enable_pipe32_sim_hwtcl                  : integer := 0;
			fixed_preset_on                          : integer := 0;
			bypass_cdc_hwtcl                         : string  := "false";
			enable_rx_buffer_checking_hwtcl          : string  := "false";
			disable_link_x2_support_hwtcl            : string  := "false";
			wrong_device_id_hwtcl                    : string  := "disable";
			data_pack_rx_hwtcl                       : string  := "disable";
			ltssm_1ms_timeout_hwtcl                  : string  := "disable";
			ltssm_freqlocked_check_hwtcl             : string  := "disable";
			deskew_comma_hwtcl                       : string  := "skp_eieos_deskw";
			device_number_hwtcl                      : integer := 0;
			pipex1_debug_sel_hwtcl                   : string  := "disable";
			pclk_out_sel_hwtcl                       : string  := "pclk";
			no_soft_reset_hwtcl                      : string  := "false";
			maximum_current_hwtcl                    : integer := 0;
			d1_support_hwtcl                         : string  := "false";
			d2_support_hwtcl                         : string  := "false";
			d0_pme_hwtcl                             : string  := "false";
			d1_pme_hwtcl                             : string  := "false";
			d2_pme_hwtcl                             : string  := "false";
			d3_hot_pme_hwtcl                         : string  := "false";
			d3_cold_pme_hwtcl                        : string  := "false";
			low_priority_vc_hwtcl                    : string  := "single_vc";
			disable_snoop_packet_hwtcl               : string  := "false";
			enable_l1_aspm_hwtcl                     : string  := "false";
			rx_ei_l0s_hwtcl                          : integer := 0;
			enable_l0s_aspm_hwtcl                    : string  := "false";
			aspm_config_management_hwtcl             : string  := "false";
			l1_exit_latency_sameclock_hwtcl          : integer := 0;
			l1_exit_latency_diffclock_hwtcl          : integer := 0;
			hot_plug_support_hwtcl                   : integer := 0;
			extended_tag_reset_hwtcl                 : string  := "false";
			no_command_completed_hwtcl               : string  := "false";
			interrupt_pin_hwtcl                      : string  := "inta";
			bridge_port_vga_enable_hwtcl             : string  := "false";
			bridge_port_ssid_support_hwtcl           : string  := "false";
			ssvid_hwtcl                              : integer := 0;
			ssid_hwtcl                               : integer := 0;
			eie_before_nfts_count_hwtcl              : integer := 4;
			gen2_diffclock_nfts_count_hwtcl          : integer := 255;
			gen2_sameclock_nfts_count_hwtcl          : integer := 255;
			l0_exit_latency_sameclock_hwtcl          : integer := 6;
			l0_exit_latency_diffclock_hwtcl          : integer := 6;
			atomic_op_routing_hwtcl                  : string  := "false";
			atomic_op_completer_32bit_hwtcl          : string  := "false";
			atomic_op_completer_64bit_hwtcl          : string  := "false";
			cas_completer_128bit_hwtcl               : string  := "false";
			ltr_mechanism_hwtcl                      : string  := "false";
			tph_completer_hwtcl                      : string  := "false";
			extended_format_field_hwtcl              : string  := "false";
			atomic_malformed_hwtcl                   : string  := "true";
			flr_capability_hwtcl                     : string  := "false";
			enable_adapter_half_rate_mode_hwtcl      : string  := "false";
			vc0_clk_enable_hwtcl                     : string  := "true";
			register_pipe_signals_hwtcl              : string  := "false";
			skp_os_gen3_count_hwtcl                  : integer := 0;
			tx_cdc_almost_empty_hwtcl                : integer := 5;
			rx_l0s_count_idl_hwtcl                   : integer := 0;
			cdc_dummy_insert_limit_hwtcl             : integer := 11;
			ei_delay_powerdown_count_hwtcl           : integer := 10;
			skp_os_schedule_count_hwtcl              : integer := 0;
			fc_init_timer_hwtcl                      : integer := 1024;
			l01_entry_latency_hwtcl                  : integer := 31;
			flow_control_update_count_hwtcl          : integer := 30;
			flow_control_timeout_count_hwtcl         : integer := 200;
			retry_buffer_last_active_address_hwtcl   : integer := 2047;
			reserved_debug_hwtcl                     : integer := 0;
			bypass_clk_switch_hwtcl                  : string  := "true";
			l2_async_logic_hwtcl                     : string  := "disable";
			indicator_hwtcl                          : integer := 0;
			diffclock_nfts_count_hwtcl               : integer := 128;
			sameclock_nfts_count_hwtcl               : integer := 128;
			rx_cdc_almost_full_hwtcl                 : integer := 12;
			tx_cdc_almost_full_hwtcl                 : integer := 11;
			credit_buffer_allocation_aux_hwtcl       : string  := "balanced";
			vc0_rx_flow_ctrl_posted_header_hwtcl     : integer := 50;
			vc0_rx_flow_ctrl_posted_data_hwtcl       : integer := 358;
			vc0_rx_flow_ctrl_nonposted_header_hwtcl  : integer := 56;
			vc0_rx_flow_ctrl_nonposted_data_hwtcl    : integer := 0;
			vc0_rx_flow_ctrl_compl_header_hwtcl      : integer := 0;
			vc0_rx_flow_ctrl_compl_data_hwtcl        : integer := 0;
			cpl_spc_header_hwtcl                     : integer := 112;
			cpl_spc_data_hwtcl                       : integer := 448;
			gen3_rxfreqlock_counter_hwtcl            : integer := 0;
			gen3_skip_ph2_ph3_hwtcl                  : integer := 0;
			g3_bypass_equlz_hwtcl                    : integer := 0;
			cvp_data_compressed_hwtcl                : string  := "false";
			cvp_data_encrypted_hwtcl                 : string  := "false";
			cvp_mode_reset_hwtcl                     : string  := "false";
			cvp_clk_reset_hwtcl                      : string  := "false";
			cseb_cpl_status_during_cvp_hwtcl         : string  := "config_retry_status";
			core_clk_sel_hwtcl                       : string  := "pld_clk";
			cvp_rate_sel_hwtcl                       : string  := "full_rate";
			g3_dis_rx_use_prst_hwtcl                 : string  := "true";
			g3_dis_rx_use_prst_ep_hwtcl              : string  := "true";
			deemphasis_enable_hwtcl                  : string  := "false";
			reconfig_to_xcvr_width                   : integer := 10;
			reconfig_from_xcvr_width                 : integer := 10;
			single_rx_detect_hwtcl                   : integer := 0;
			hip_hard_reset_hwtcl                     : integer := 0;
			use_cvp_update_core_pof_hwtcl            : integer := 0;
			pcie_inspector_hwtcl                     : integer := 0;
			tlp_inspector_hwtcl                      : integer := 0;
			tlp_inspector_use_signal_probe_hwtcl     : integer := 0;
			tlp_insp_trg_dw0_hwtcl                   : integer := 2049;
			tlp_insp_trg_dw1_hwtcl                   : integer := 0;
			tlp_insp_trg_dw2_hwtcl                   : integer := 0;
			tlp_insp_trg_dw3_hwtcl                   : integer := 0;
			hwtcl_override_g2_txvod                  : integer := 1;
			rpre_emph_a_val_hwtcl                    : integer := 9;
			rpre_emph_b_val_hwtcl                    : integer := 0;
			rpre_emph_c_val_hwtcl                    : integer := 16;
			rpre_emph_d_val_hwtcl                    : integer := 13;
			rpre_emph_e_val_hwtcl                    : integer := 5;
			rvod_sel_a_val_hwtcl                     : integer := 42;
			rvod_sel_b_val_hwtcl                     : integer := 38;
			rvod_sel_c_val_hwtcl                     : integer := 38;
			rvod_sel_d_val_hwtcl                     : integer := 43;
			rvod_sel_e_val_hwtcl                     : integer := 15;
			hwtcl_override_g3rxcoef                  : integer := 0;
			gen3_coeff_1_hwtcl                       : integer := 7;
			gen3_coeff_1_sel_hwtcl                   : string  := "preset_1";
			gen3_coeff_1_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_1_nxtber_more_ptr_hwtcl       : integer := 1;
			gen3_coeff_1_nxtber_more_hwtcl           : string  := "g3_coeff_1_nxtber_more";
			gen3_coeff_1_nxtber_less_ptr_hwtcl       : integer := 1;
			gen3_coeff_1_nxtber_less_hwtcl           : string  := "g3_coeff_1_nxtber_less";
			gen3_coeff_1_reqber_hwtcl                : integer := 0;
			gen3_coeff_1_ber_meas_hwtcl              : integer := 2;
			gen3_coeff_2_hwtcl                       : integer := 0;
			gen3_coeff_2_sel_hwtcl                   : string  := "preset_2";
			gen3_coeff_2_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_2_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_2_nxtber_more_hwtcl           : string  := "g3_coeff_2_nxtber_more";
			gen3_coeff_2_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_2_nxtber_less_hwtcl           : string  := "g3_coeff_2_nxtber_less";
			gen3_coeff_2_reqber_hwtcl                : integer := 0;
			gen3_coeff_2_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_3_hwtcl                       : integer := 0;
			gen3_coeff_3_sel_hwtcl                   : string  := "preset_3";
			gen3_coeff_3_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_3_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_3_nxtber_more_hwtcl           : string  := "g3_coeff_3_nxtber_more";
			gen3_coeff_3_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_3_nxtber_less_hwtcl           : string  := "g3_coeff_3_nxtber_less";
			gen3_coeff_3_reqber_hwtcl                : integer := 0;
			gen3_coeff_3_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_4_hwtcl                       : integer := 0;
			gen3_coeff_4_sel_hwtcl                   : string  := "preset_4";
			gen3_coeff_4_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_4_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_4_nxtber_more_hwtcl           : string  := "g3_coeff_4_nxtber_more";
			gen3_coeff_4_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_4_nxtber_less_hwtcl           : string  := "g3_coeff_4_nxtber_less";
			gen3_coeff_4_reqber_hwtcl                : integer := 0;
			gen3_coeff_4_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_5_hwtcl                       : integer := 0;
			gen3_coeff_5_sel_hwtcl                   : string  := "preset_5";
			gen3_coeff_5_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_5_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_5_nxtber_more_hwtcl           : string  := "g3_coeff_5_nxtber_more";
			gen3_coeff_5_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_5_nxtber_less_hwtcl           : string  := "g3_coeff_5_nxtber_less";
			gen3_coeff_5_reqber_hwtcl                : integer := 0;
			gen3_coeff_5_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_6_hwtcl                       : integer := 0;
			gen3_coeff_6_sel_hwtcl                   : string  := "preset_6";
			gen3_coeff_6_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_6_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_6_nxtber_more_hwtcl           : string  := "g3_coeff_6_nxtber_more";
			gen3_coeff_6_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_6_nxtber_less_hwtcl           : string  := "g3_coeff_6_nxtber_less";
			gen3_coeff_6_reqber_hwtcl                : integer := 0;
			gen3_coeff_6_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_7_hwtcl                       : integer := 0;
			gen3_coeff_7_sel_hwtcl                   : string  := "preset_7";
			gen3_coeff_7_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_7_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_7_nxtber_more_hwtcl           : string  := "g3_coeff_7_nxtber_more";
			gen3_coeff_7_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_7_nxtber_less_hwtcl           : string  := "g3_coeff_7_nxtber_less";
			gen3_coeff_7_reqber_hwtcl                : integer := 0;
			gen3_coeff_7_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_8_hwtcl                       : integer := 0;
			gen3_coeff_8_sel_hwtcl                   : string  := "preset_8";
			gen3_coeff_8_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_8_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_8_nxtber_more_hwtcl           : string  := "g3_coeff_8_nxtber_more";
			gen3_coeff_8_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_8_nxtber_less_hwtcl           : string  := "g3_coeff_8_nxtber_less";
			gen3_coeff_8_reqber_hwtcl                : integer := 0;
			gen3_coeff_8_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_9_hwtcl                       : integer := 0;
			gen3_coeff_9_sel_hwtcl                   : string  := "preset_9";
			gen3_coeff_9_preset_hint_hwtcl           : integer := 0;
			gen3_coeff_9_nxtber_more_ptr_hwtcl       : integer := 0;
			gen3_coeff_9_nxtber_more_hwtcl           : string  := "g3_coeff_9_nxtber_more";
			gen3_coeff_9_nxtber_less_ptr_hwtcl       : integer := 0;
			gen3_coeff_9_nxtber_less_hwtcl           : string  := "g3_coeff_9_nxtber_less";
			gen3_coeff_9_reqber_hwtcl                : integer := 0;
			gen3_coeff_9_ber_meas_hwtcl              : integer := 0;
			gen3_coeff_10_hwtcl                      : integer := 0;
			gen3_coeff_10_sel_hwtcl                  : string  := "preset_10";
			gen3_coeff_10_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_10_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_10_nxtber_more_hwtcl          : string  := "g3_coeff_10_nxtber_more";
			gen3_coeff_10_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_10_nxtber_less_hwtcl          : string  := "g3_coeff_10_nxtber_less";
			gen3_coeff_10_reqber_hwtcl               : integer := 0;
			gen3_coeff_10_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_11_hwtcl                      : integer := 0;
			gen3_coeff_11_sel_hwtcl                  : string  := "preset_11";
			gen3_coeff_11_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_11_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_11_nxtber_more_hwtcl          : string  := "g3_coeff_11_nxtber_more";
			gen3_coeff_11_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_11_nxtber_less_hwtcl          : string  := "g3_coeff_11_nxtber_less";
			gen3_coeff_11_reqber_hwtcl               : integer := 0;
			gen3_coeff_11_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_12_hwtcl                      : integer := 0;
			gen3_coeff_12_sel_hwtcl                  : string  := "preset_12";
			gen3_coeff_12_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_12_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_12_nxtber_more_hwtcl          : string  := "g3_coeff_12_nxtber_more";
			gen3_coeff_12_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_12_nxtber_less_hwtcl          : string  := "g3_coeff_12_nxtber_less";
			gen3_coeff_12_reqber_hwtcl               : integer := 0;
			gen3_coeff_12_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_13_hwtcl                      : integer := 0;
			gen3_coeff_13_sel_hwtcl                  : string  := "preset_13";
			gen3_coeff_13_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_13_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_13_nxtber_more_hwtcl          : string  := "g3_coeff_13_nxtber_more";
			gen3_coeff_13_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_13_nxtber_less_hwtcl          : string  := "g3_coeff_13_nxtber_less";
			gen3_coeff_13_reqber_hwtcl               : integer := 0;
			gen3_coeff_13_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_14_hwtcl                      : integer := 0;
			gen3_coeff_14_sel_hwtcl                  : string  := "preset_14";
			gen3_coeff_14_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_14_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_14_nxtber_more_hwtcl          : string  := "g3_coeff_14_nxtber_more";
			gen3_coeff_14_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_14_nxtber_less_hwtcl          : string  := "g3_coeff_14_nxtber_less";
			gen3_coeff_14_reqber_hwtcl               : integer := 0;
			gen3_coeff_14_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_15_hwtcl                      : integer := 0;
			gen3_coeff_15_sel_hwtcl                  : string  := "preset_15";
			gen3_coeff_15_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_15_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_15_nxtber_more_hwtcl          : string  := "g3_coeff_15_nxtber_more";
			gen3_coeff_15_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_15_nxtber_less_hwtcl          : string  := "g3_coeff_15_nxtber_less";
			gen3_coeff_15_reqber_hwtcl               : integer := 0;
			gen3_coeff_15_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_16_hwtcl                      : integer := 0;
			gen3_coeff_16_sel_hwtcl                  : string  := "preset_16";
			gen3_coeff_16_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_16_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_16_nxtber_more_hwtcl          : string  := "g3_coeff_16_nxtber_more";
			gen3_coeff_16_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_16_nxtber_less_hwtcl          : string  := "g3_coeff_16_nxtber_less";
			gen3_coeff_16_reqber_hwtcl               : integer := 0;
			gen3_coeff_16_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_17_hwtcl                      : integer := 0;
			gen3_coeff_17_sel_hwtcl                  : string  := "preset_17";
			gen3_coeff_17_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_17_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_17_nxtber_more_hwtcl          : string  := "g3_coeff_17_nxtber_more";
			gen3_coeff_17_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_17_nxtber_less_hwtcl          : string  := "g3_coeff_17_nxtber_less";
			gen3_coeff_17_reqber_hwtcl               : integer := 0;
			gen3_coeff_17_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_18_hwtcl                      : integer := 0;
			gen3_coeff_18_sel_hwtcl                  : string  := "preset_18";
			gen3_coeff_18_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_18_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_18_nxtber_more_hwtcl          : string  := "g3_coeff_18_nxtber_more";
			gen3_coeff_18_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_18_nxtber_less_hwtcl          : string  := "g3_coeff_18_nxtber_less";
			gen3_coeff_18_reqber_hwtcl               : integer := 0;
			gen3_coeff_18_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_19_hwtcl                      : integer := 0;
			gen3_coeff_19_sel_hwtcl                  : string  := "preset_19";
			gen3_coeff_19_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_19_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_19_nxtber_more_hwtcl          : string  := "g3_coeff_19_nxtber_more";
			gen3_coeff_19_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_19_nxtber_less_hwtcl          : string  := "g3_coeff_19_nxtber_less";
			gen3_coeff_19_reqber_hwtcl               : integer := 0;
			gen3_coeff_19_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_20_hwtcl                      : integer := 0;
			gen3_coeff_20_sel_hwtcl                  : string  := "preset_20";
			gen3_coeff_20_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_20_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_20_nxtber_more_hwtcl          : string  := "g3_coeff_20_nxtber_more";
			gen3_coeff_20_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_20_nxtber_less_hwtcl          : string  := "g3_coeff_20_nxtber_less";
			gen3_coeff_20_reqber_hwtcl               : integer := 0;
			gen3_coeff_20_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_21_hwtcl                      : integer := 0;
			gen3_coeff_21_sel_hwtcl                  : string  := "preset_21";
			gen3_coeff_21_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_21_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_21_nxtber_more_hwtcl          : string  := "g3_coeff_21_nxtber_more";
			gen3_coeff_21_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_21_nxtber_less_hwtcl          : string  := "g3_coeff_21_nxtber_less";
			gen3_coeff_21_reqber_hwtcl               : integer := 0;
			gen3_coeff_21_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_22_hwtcl                      : integer := 0;
			gen3_coeff_22_sel_hwtcl                  : string  := "preset_22";
			gen3_coeff_22_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_22_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_22_nxtber_more_hwtcl          : string  := "g3_coeff_22_nxtber_more";
			gen3_coeff_22_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_22_nxtber_less_hwtcl          : string  := "g3_coeff_22_nxtber_less";
			gen3_coeff_22_reqber_hwtcl               : integer := 0;
			gen3_coeff_22_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_23_hwtcl                      : integer := 0;
			gen3_coeff_23_sel_hwtcl                  : string  := "preset_23";
			gen3_coeff_23_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_23_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_23_nxtber_more_hwtcl          : string  := "g3_coeff_23_nxtber_more";
			gen3_coeff_23_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_23_nxtber_less_hwtcl          : string  := "g3_coeff_23_nxtber_less";
			gen3_coeff_23_reqber_hwtcl               : integer := 0;
			gen3_coeff_23_ber_meas_hwtcl             : integer := 0;
			gen3_coeff_24_hwtcl                      : integer := 0;
			gen3_coeff_24_sel_hwtcl                  : string  := "preset_24";
			gen3_coeff_24_preset_hint_hwtcl          : integer := 0;
			gen3_coeff_24_nxtber_more_ptr_hwtcl      : integer := 0;
			gen3_coeff_24_nxtber_more_hwtcl          : string  := "g3_coeff_24_nxtber_more";
			gen3_coeff_24_nxtber_less_ptr_hwtcl      : integer := 0;
			gen3_coeff_24_nxtber_less_hwtcl          : string  := "g3_coeff_24_nxtber_less";
			gen3_coeff_24_reqber_hwtcl               : integer := 0;
			gen3_coeff_24_ber_meas_hwtcl             : integer := 0;
			hwtcl_override_g3txcoef                  : integer := 0;
			gen3_preset_coeff_1_hwtcl                : integer := 0;
			gen3_preset_coeff_2_hwtcl                : integer := 0;
			gen3_preset_coeff_3_hwtcl                : integer := 0;
			gen3_preset_coeff_4_hwtcl                : integer := 0;
			gen3_preset_coeff_5_hwtcl                : integer := 0;
			gen3_preset_coeff_6_hwtcl                : integer := 0;
			gen3_preset_coeff_7_hwtcl                : integer := 0;
			gen3_preset_coeff_8_hwtcl                : integer := 0;
			gen3_preset_coeff_9_hwtcl                : integer := 0;
			gen3_preset_coeff_10_hwtcl               : integer := 0;
			gen3_preset_coeff_11_hwtcl               : integer := 0;
			gen3_low_freq_hwtcl                      : integer := 0;
			full_swing_hwtcl                         : integer := 35;
			gen3_full_swing_hwtcl                    : integer := 35;
			use_atx_pll_hwtcl                        : integer := 0;
			low_latency_mode_hwtcl                   : integer := 0
		);
		port (
			npor                   : in  std_logic                       := 'X';             -- npor
			pin_perst              : in  std_logic                       := 'X';             -- pin_perst
			lmi_addr               : in  std_logic_vector(11 downto 0)   := (others => 'X'); -- lmi_addr
			lmi_din                : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- lmi_din
			lmi_rden               : in  std_logic                       := 'X';             -- lmi_rden
			lmi_wren               : in  std_logic                       := 'X';             -- lmi_wren
			lmi_ack                : out std_logic;                                          -- lmi_ack
			lmi_dout               : out std_logic_vector(31 downto 0);                      -- lmi_dout
			hpg_ctrler             : in  std_logic_vector(4 downto 0)    := (others => 'X'); -- hpg_ctrler
			tl_cfg_add             : out std_logic_vector(3 downto 0);                       -- tl_cfg_add
			tl_cfg_ctl             : out std_logic_vector(31 downto 0);                      -- tl_cfg_ctl
			tl_cfg_sts             : out std_logic_vector(52 downto 0);                      -- tl_cfg_sts
			cpl_err                : in  std_logic_vector(6 downto 0)    := (others => 'X'); -- cpl_err
			cpl_pending            : in  std_logic                       := 'X';             -- cpl_pending
			pm_auxpwr              : in  std_logic                       := 'X';             -- pm_auxpwr
			pm_data                : in  std_logic_vector(9 downto 0)    := (others => 'X'); -- pm_data
			pme_to_cr              : in  std_logic                       := 'X';             -- pme_to_cr
			pm_event               : in  std_logic                       := 'X';             -- pm_event
			pme_to_sr              : out std_logic;                                          -- pme_to_sr
			rx_st_sop              : out std_logic_vector(0 downto 0);                       -- startofpacket
			rx_st_eop              : out std_logic_vector(0 downto 0);                       -- endofpacket
			rx_st_err              : out std_logic_vector(0 downto 0);                       -- error
			rx_st_valid            : out std_logic_vector(0 downto 0);                       -- valid
			rx_st_empty            : out std_logic_vector(1 downto 0);                       -- empty
			rx_st_ready            : in  std_logic                       := 'X';             -- ready
			rx_st_data             : out std_logic_vector(255 downto 0);                     -- data
			rx_st_parity           : out std_logic_vector(31 downto 0);                      -- parity
			rx_st_bar              : out std_logic_vector(7 downto 0);                       -- rx_st_bar
			rx_st_mask             : in  std_logic                       := 'X';             -- rx_st_mask
			tx_st_sop              : in  std_logic_vector(0 downto 0)    := (others => 'X'); -- startofpacket
			tx_st_eop              : in  std_logic_vector(0 downto 0)    := (others => 'X'); -- endofpacket
			tx_st_err              : in  std_logic_vector(0 downto 0)    := (others => 'X'); -- error
			tx_st_valid            : in  std_logic_vector(0 downto 0)    := (others => 'X'); -- valid
			tx_st_empty            : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- empty
			tx_st_ready            : out std_logic;                                          -- ready
			tx_st_data             : in  std_logic_vector(255 downto 0)  := (others => 'X'); -- data
			tx_st_parity           : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- parity
			tx_cred_datafccp       : out std_logic_vector(11 downto 0);                      -- tx_cred_datafccp
			tx_cred_datafcnp       : out std_logic_vector(11 downto 0);                      -- tx_cred_datafcnp
			tx_cred_datafcp        : out std_logic_vector(11 downto 0);                      -- tx_cred_datafcp
			tx_cred_fchipcons      : out std_logic_vector(5 downto 0);                       -- tx_cred_fchipcons
			tx_cred_fcinfinite     : out std_logic_vector(5 downto 0);                       -- tx_cred_fcinfinite
			tx_cred_hdrfccp        : out std_logic_vector(7 downto 0);                       -- tx_cred_hdrfccp
			tx_cred_hdrfcnp        : out std_logic_vector(7 downto 0);                       -- tx_cred_hdrfcnp
			tx_cred_hdrfcp         : out std_logic_vector(7 downto 0);                       -- tx_cred_hdrfcp
			pld_clk                : in  std_logic                       := 'X';             -- clk
			coreclkout_hip         : out std_logic;                                          -- clk
			refclk                 : in  std_logic                       := 'X';             -- clk
			reset_status           : out std_logic;                                          -- reset_status
			serdes_pll_locked      : out std_logic;                                          -- serdes_pll_locked
			pld_clk_inuse          : out std_logic;                                          -- pld_clk_inuse
			pld_core_ready         : in  std_logic                       := 'X';             -- pld_core_ready
			testin_zero            : out std_logic;                                          -- testin_zero
			reconfig_to_xcvr       : in  std_logic_vector(769 downto 0)  := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr     : out std_logic_vector(505 downto 0);                     -- reconfig_from_xcvr
			rx_in0                 : in  std_logic                       := 'X';             -- rx_in0
			rx_in1                 : in  std_logic                       := 'X';             -- rx_in1
			rx_in2                 : in  std_logic                       := 'X';             -- rx_in2
			rx_in3                 : in  std_logic                       := 'X';             -- rx_in3
			rx_in4                 : in  std_logic                       := 'X';             -- rx_in4
			rx_in5                 : in  std_logic                       := 'X';             -- rx_in5
			rx_in6                 : in  std_logic                       := 'X';             -- rx_in6
			rx_in7                 : in  std_logic                       := 'X';             -- rx_in7
			tx_out0                : out std_logic;                                          -- tx_out0
			tx_out1                : out std_logic;                                          -- tx_out1
			tx_out2                : out std_logic;                                          -- tx_out2
			tx_out3                : out std_logic;                                          -- tx_out3
			tx_out4                : out std_logic;                                          -- tx_out4
			tx_out5                : out std_logic;                                          -- tx_out5
			tx_out6                : out std_logic;                                          -- tx_out6
			tx_out7                : out std_logic;                                          -- tx_out7
			sim_pipe_pclk_in       : in  std_logic                       := 'X';             -- sim_pipe_pclk_in
			sim_pipe_rate          : out std_logic_vector(1 downto 0);                       -- sim_pipe_rate
			sim_ltssmstate         : out std_logic_vector(4 downto 0);                       -- sim_ltssmstate
			eidleinfersel0         : out std_logic_vector(2 downto 0);                       -- eidleinfersel0
			eidleinfersel1         : out std_logic_vector(2 downto 0);                       -- eidleinfersel1
			eidleinfersel2         : out std_logic_vector(2 downto 0);                       -- eidleinfersel2
			eidleinfersel3         : out std_logic_vector(2 downto 0);                       -- eidleinfersel3
			eidleinfersel4         : out std_logic_vector(2 downto 0);                       -- eidleinfersel4
			eidleinfersel5         : out std_logic_vector(2 downto 0);                       -- eidleinfersel5
			eidleinfersel6         : out std_logic_vector(2 downto 0);                       -- eidleinfersel6
			eidleinfersel7         : out std_logic_vector(2 downto 0);                       -- eidleinfersel7
			powerdown0             : out std_logic_vector(1 downto 0);                       -- powerdown0
			powerdown1             : out std_logic_vector(1 downto 0);                       -- powerdown1
			powerdown2             : out std_logic_vector(1 downto 0);                       -- powerdown2
			powerdown3             : out std_logic_vector(1 downto 0);                       -- powerdown3
			powerdown4             : out std_logic_vector(1 downto 0);                       -- powerdown4
			powerdown5             : out std_logic_vector(1 downto 0);                       -- powerdown5
			powerdown6             : out std_logic_vector(1 downto 0);                       -- powerdown6
			powerdown7             : out std_logic_vector(1 downto 0);                       -- powerdown7
			rxpolarity0            : out std_logic;                                          -- rxpolarity0
			rxpolarity1            : out std_logic;                                          -- rxpolarity1
			rxpolarity2            : out std_logic;                                          -- rxpolarity2
			rxpolarity3            : out std_logic;                                          -- rxpolarity3
			rxpolarity4            : out std_logic;                                          -- rxpolarity4
			rxpolarity5            : out std_logic;                                          -- rxpolarity5
			rxpolarity6            : out std_logic;                                          -- rxpolarity6
			rxpolarity7            : out std_logic;                                          -- rxpolarity7
			txcompl0               : out std_logic;                                          -- txcompl0
			txcompl1               : out std_logic;                                          -- txcompl1
			txcompl2               : out std_logic;                                          -- txcompl2
			txcompl3               : out std_logic;                                          -- txcompl3
			txcompl4               : out std_logic;                                          -- txcompl4
			txcompl5               : out std_logic;                                          -- txcompl5
			txcompl6               : out std_logic;                                          -- txcompl6
			txcompl7               : out std_logic;                                          -- txcompl7
			txdata0                : out std_logic_vector(7 downto 0);                       -- txdata0
			txdata1                : out std_logic_vector(7 downto 0);                       -- txdata1
			txdata2                : out std_logic_vector(7 downto 0);                       -- txdata2
			txdata3                : out std_logic_vector(7 downto 0);                       -- txdata3
			txdata4                : out std_logic_vector(7 downto 0);                       -- txdata4
			txdata5                : out std_logic_vector(7 downto 0);                       -- txdata5
			txdata6                : out std_logic_vector(7 downto 0);                       -- txdata6
			txdata7                : out std_logic_vector(7 downto 0);                       -- txdata7
			txdatak0               : out std_logic;                                          -- txdatak0
			txdatak1               : out std_logic;                                          -- txdatak1
			txdatak2               : out std_logic;                                          -- txdatak2
			txdatak3               : out std_logic;                                          -- txdatak3
			txdatak4               : out std_logic;                                          -- txdatak4
			txdatak5               : out std_logic;                                          -- txdatak5
			txdatak6               : out std_logic;                                          -- txdatak6
			txdatak7               : out std_logic;                                          -- txdatak7
			txdetectrx0            : out std_logic;                                          -- txdetectrx0
			txdetectrx1            : out std_logic;                                          -- txdetectrx1
			txdetectrx2            : out std_logic;                                          -- txdetectrx2
			txdetectrx3            : out std_logic;                                          -- txdetectrx3
			txdetectrx4            : out std_logic;                                          -- txdetectrx4
			txdetectrx5            : out std_logic;                                          -- txdetectrx5
			txdetectrx6            : out std_logic;                                          -- txdetectrx6
			txdetectrx7            : out std_logic;                                          -- txdetectrx7
			txelecidle0            : out std_logic;                                          -- txelecidle0
			txelecidle1            : out std_logic;                                          -- txelecidle1
			txelecidle2            : out std_logic;                                          -- txelecidle2
			txelecidle3            : out std_logic;                                          -- txelecidle3
			txelecidle4            : out std_logic;                                          -- txelecidle4
			txelecidle5            : out std_logic;                                          -- txelecidle5
			txelecidle6            : out std_logic;                                          -- txelecidle6
			txelecidle7            : out std_logic;                                          -- txelecidle7
			txdeemph0              : out std_logic;                                          -- txdeemph0
			txdeemph1              : out std_logic;                                          -- txdeemph1
			txdeemph2              : out std_logic;                                          -- txdeemph2
			txdeemph3              : out std_logic;                                          -- txdeemph3
			txdeemph4              : out std_logic;                                          -- txdeemph4
			txdeemph5              : out std_logic;                                          -- txdeemph5
			txdeemph6              : out std_logic;                                          -- txdeemph6
			txdeemph7              : out std_logic;                                          -- txdeemph7
			txmargin0              : out std_logic_vector(2 downto 0);                       -- txmargin0
			txmargin1              : out std_logic_vector(2 downto 0);                       -- txmargin1
			txmargin2              : out std_logic_vector(2 downto 0);                       -- txmargin2
			txmargin3              : out std_logic_vector(2 downto 0);                       -- txmargin3
			txmargin4              : out std_logic_vector(2 downto 0);                       -- txmargin4
			txmargin5              : out std_logic_vector(2 downto 0);                       -- txmargin5
			txmargin6              : out std_logic_vector(2 downto 0);                       -- txmargin6
			txmargin7              : out std_logic_vector(2 downto 0);                       -- txmargin7
			txswing0               : out std_logic;                                          -- txswing0
			txswing1               : out std_logic;                                          -- txswing1
			txswing2               : out std_logic;                                          -- txswing2
			txswing3               : out std_logic;                                          -- txswing3
			txswing4               : out std_logic;                                          -- txswing4
			txswing5               : out std_logic;                                          -- txswing5
			txswing6               : out std_logic;                                          -- txswing6
			txswing7               : out std_logic;                                          -- txswing7
			phystatus0             : in  std_logic                       := 'X';             -- phystatus0
			phystatus1             : in  std_logic                       := 'X';             -- phystatus1
			phystatus2             : in  std_logic                       := 'X';             -- phystatus2
			phystatus3             : in  std_logic                       := 'X';             -- phystatus3
			phystatus4             : in  std_logic                       := 'X';             -- phystatus4
			phystatus5             : in  std_logic                       := 'X';             -- phystatus5
			phystatus6             : in  std_logic                       := 'X';             -- phystatus6
			phystatus7             : in  std_logic                       := 'X';             -- phystatus7
			rxdata0                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata0
			rxdata1                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata1
			rxdata2                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata2
			rxdata3                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata3
			rxdata4                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata4
			rxdata5                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata5
			rxdata6                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata6
			rxdata7                : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- rxdata7
			rxdatak0               : in  std_logic                       := 'X';             -- rxdatak0
			rxdatak1               : in  std_logic                       := 'X';             -- rxdatak1
			rxdatak2               : in  std_logic                       := 'X';             -- rxdatak2
			rxdatak3               : in  std_logic                       := 'X';             -- rxdatak3
			rxdatak4               : in  std_logic                       := 'X';             -- rxdatak4
			rxdatak5               : in  std_logic                       := 'X';             -- rxdatak5
			rxdatak6               : in  std_logic                       := 'X';             -- rxdatak6
			rxdatak7               : in  std_logic                       := 'X';             -- rxdatak7
			rxelecidle0            : in  std_logic                       := 'X';             -- rxelecidle0
			rxelecidle1            : in  std_logic                       := 'X';             -- rxelecidle1
			rxelecidle2            : in  std_logic                       := 'X';             -- rxelecidle2
			rxelecidle3            : in  std_logic                       := 'X';             -- rxelecidle3
			rxelecidle4            : in  std_logic                       := 'X';             -- rxelecidle4
			rxelecidle5            : in  std_logic                       := 'X';             -- rxelecidle5
			rxelecidle6            : in  std_logic                       := 'X';             -- rxelecidle6
			rxelecidle7            : in  std_logic                       := 'X';             -- rxelecidle7
			rxstatus0              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus0
			rxstatus1              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus1
			rxstatus2              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus2
			rxstatus3              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus3
			rxstatus4              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus4
			rxstatus5              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus5
			rxstatus6              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus6
			rxstatus7              : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- rxstatus7
			rxvalid0               : in  std_logic                       := 'X';             -- rxvalid0
			rxvalid1               : in  std_logic                       := 'X';             -- rxvalid1
			rxvalid2               : in  std_logic                       := 'X';             -- rxvalid2
			rxvalid3               : in  std_logic                       := 'X';             -- rxvalid3
			rxvalid4               : in  std_logic                       := 'X';             -- rxvalid4
			rxvalid5               : in  std_logic                       := 'X';             -- rxvalid5
			rxvalid6               : in  std_logic                       := 'X';             -- rxvalid6
			rxvalid7               : in  std_logic                       := 'X';             -- rxvalid7
			app_int_sts            : in  std_logic                       := 'X';             -- app_int_sts
			app_msi_num            : in  std_logic_vector(4 downto 0)    := (others => 'X'); -- app_msi_num
			app_msi_req            : in  std_logic                       := 'X';             -- app_msi_req
			app_msi_tc             : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- app_msi_tc
			app_int_ack            : out std_logic;                                          -- app_int_ack
			app_msi_ack            : out std_logic;                                          -- app_msi_ack
			cseb_rddata            : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- cseb_rddata
			cseb_rdresponse        : in  std_logic_vector(4 downto 0)    := (others => 'X'); -- cseb_rdresponse
			cseb_waitrequest       : in  std_logic                       := 'X';             -- cseb_waitrequest
			cseb_wrresponse        : in  std_logic_vector(4 downto 0)    := (others => 'X'); -- cseb_wrresponse
			cseb_wrresp_valid      : in  std_logic                       := 'X';             -- cseb_wrresp_valid
			cseb_addr              : out std_logic_vector(32 downto 0);                      -- cseb_addr
			cseb_be                : out std_logic_vector(3 downto 0);                       -- cseb_be
			cseb_rden              : out std_logic;                                          -- cseb_rden
			cseb_wrdata            : out std_logic_vector(31 downto 0);                      -- cseb_wrdata
			cseb_wren              : out std_logic;                                          -- cseb_wren
			cseb_wrresp_req        : out std_logic;                                          -- cseb_wrresp_req
			cseb_rddata_parity     : in  std_logic_vector(3 downto 0)    := (others => 'X'); -- cseb_rddata_parity
			cseb_addr_parity       : out std_logic_vector(4 downto 0);                       -- cseb_addr_parity
			cseb_wrdata_parity     : out std_logic_vector(3 downto 0);                       -- cseb_wrdata_parity
			test_in                : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- test_in
			simu_mode_pipe         : in  std_logic                       := 'X';             -- simu_mode_pipe
			derr_cor_ext_rcv       : out std_logic;                                          -- derr_cor_ext_rcv
			derr_cor_ext_rpl       : out std_logic;                                          -- derr_cor_ext_rpl
			derr_rpl               : out std_logic;                                          -- derr_rpl
			dlup                   : out std_logic;                                          -- dlup
			dlup_exit              : out std_logic;                                          -- dlup_exit
			ev128ns                : out std_logic;                                          -- ev128ns
			ev1us                  : out std_logic;                                          -- ev1us
			hotrst_exit            : out std_logic;                                          -- hotrst_exit
			int_status             : out std_logic_vector(3 downto 0);                       -- int_status
			l2_exit                : out std_logic;                                          -- l2_exit
			lane_act               : out std_logic_vector(3 downto 0);                       -- lane_act
			ltssmstate             : out std_logic_vector(4 downto 0);                       -- ltssmstate
			rx_par_err             : out std_logic;                                          -- rx_par_err
			tx_par_err             : out std_logic_vector(1 downto 0);                       -- tx_par_err
			cfg_par_err            : out std_logic;                                          -- cfg_par_err
			ko_cpl_spc_header      : out std_logic_vector(7 downto 0);                       -- ko_cpl_spc_header
			ko_cpl_spc_data        : out std_logic_vector(11 downto 0);                      -- ko_cpl_spc_data
			currentspeed           : out std_logic_vector(1 downto 0);                       -- currentspeed
			rx_st_be               : out std_logic_vector(31 downto 0);                      -- rx_st_be
			tx_cons_cred_sel       : in  std_logic                       := 'X';             -- tx_cons_cred_sel
			sim_pipe_pclk_out      : out std_logic;                                          -- sim_pipe_pclk_out
			rxdataskip0            : in  std_logic                       := 'X';             -- rxdataskip0
			rxdataskip1            : in  std_logic                       := 'X';             -- rxdataskip1
			rxdataskip2            : in  std_logic                       := 'X';             -- rxdataskip2
			rxdataskip3            : in  std_logic                       := 'X';             -- rxdataskip3
			rxdataskip4            : in  std_logic                       := 'X';             -- rxdataskip4
			rxdataskip5            : in  std_logic                       := 'X';             -- rxdataskip5
			rxdataskip6            : in  std_logic                       := 'X';             -- rxdataskip6
			rxdataskip7            : in  std_logic                       := 'X';             -- rxdataskip7
			rxblkst0               : in  std_logic                       := 'X';             -- rxblkst0
			rxblkst1               : in  std_logic                       := 'X';             -- rxblkst1
			rxblkst2               : in  std_logic                       := 'X';             -- rxblkst2
			rxblkst3               : in  std_logic                       := 'X';             -- rxblkst3
			rxblkst4               : in  std_logic                       := 'X';             -- rxblkst4
			rxblkst5               : in  std_logic                       := 'X';             -- rxblkst5
			rxblkst6               : in  std_logic                       := 'X';             -- rxblkst6
			rxblkst7               : in  std_logic                       := 'X';             -- rxblkst7
			rxsynchd0              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd0
			rxsynchd1              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd1
			rxsynchd2              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd2
			rxsynchd3              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd3
			rxsynchd4              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd4
			rxsynchd5              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd5
			rxsynchd6              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd6
			rxsynchd7              : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- rxsynchd7
			rxfreqlocked0          : in  std_logic                       := 'X';             -- rxfreqlocked0
			rxfreqlocked1          : in  std_logic                       := 'X';             -- rxfreqlocked1
			rxfreqlocked2          : in  std_logic                       := 'X';             -- rxfreqlocked2
			rxfreqlocked3          : in  std_logic                       := 'X';             -- rxfreqlocked3
			rxfreqlocked4          : in  std_logic                       := 'X';             -- rxfreqlocked4
			rxfreqlocked5          : in  std_logic                       := 'X';             -- rxfreqlocked5
			rxfreqlocked6          : in  std_logic                       := 'X';             -- rxfreqlocked6
			rxfreqlocked7          : in  std_logic                       := 'X';             -- rxfreqlocked7
			currentcoeff0          : out std_logic_vector(17 downto 0);                      -- currentcoeff0
			currentcoeff1          : out std_logic_vector(17 downto 0);                      -- currentcoeff1
			currentcoeff2          : out std_logic_vector(17 downto 0);                      -- currentcoeff2
			currentcoeff3          : out std_logic_vector(17 downto 0);                      -- currentcoeff3
			currentcoeff4          : out std_logic_vector(17 downto 0);                      -- currentcoeff4
			currentcoeff5          : out std_logic_vector(17 downto 0);                      -- currentcoeff5
			currentcoeff6          : out std_logic_vector(17 downto 0);                      -- currentcoeff6
			currentcoeff7          : out std_logic_vector(17 downto 0);                      -- currentcoeff7
			currentrxpreset0       : out std_logic_vector(2 downto 0);                       -- currentrxpreset0
			currentrxpreset1       : out std_logic_vector(2 downto 0);                       -- currentrxpreset1
			currentrxpreset2       : out std_logic_vector(2 downto 0);                       -- currentrxpreset2
			currentrxpreset3       : out std_logic_vector(2 downto 0);                       -- currentrxpreset3
			currentrxpreset4       : out std_logic_vector(2 downto 0);                       -- currentrxpreset4
			currentrxpreset5       : out std_logic_vector(2 downto 0);                       -- currentrxpreset5
			currentrxpreset6       : out std_logic_vector(2 downto 0);                       -- currentrxpreset6
			currentrxpreset7       : out std_logic_vector(2 downto 0);                       -- currentrxpreset7
			txsynchd0              : out std_logic_vector(1 downto 0);                       -- txsynchd0
			txsynchd1              : out std_logic_vector(1 downto 0);                       -- txsynchd1
			txsynchd2              : out std_logic_vector(1 downto 0);                       -- txsynchd2
			txsynchd3              : out std_logic_vector(1 downto 0);                       -- txsynchd3
			txsynchd4              : out std_logic_vector(1 downto 0);                       -- txsynchd4
			txsynchd5              : out std_logic_vector(1 downto 0);                       -- txsynchd5
			txsynchd6              : out std_logic_vector(1 downto 0);                       -- txsynchd6
			txsynchd7              : out std_logic_vector(1 downto 0);                       -- txsynchd7
			txblkst0               : out std_logic;                                          -- txblkst0
			txblkst1               : out std_logic;                                          -- txblkst1
			txblkst2               : out std_logic;                                          -- txblkst2
			txblkst3               : out std_logic;                                          -- txblkst3
			txblkst4               : out std_logic;                                          -- txblkst4
			txblkst5               : out std_logic;                                          -- txblkst5
			txblkst6               : out std_logic;                                          -- txblkst6
			txblkst7               : out std_logic;                                          -- txblkst7
			aer_msi_num            : in  std_logic_vector(4 downto 0)    := (others => 'X'); -- aer_msi_num
			pex_msi_num            : in  std_logic_vector(4 downto 0)    := (others => 'X'); -- pex_msi_num
			serr_out               : out std_logic;                                          -- serr_out
			hip_reconfig_clk       : in  std_logic                       := 'X';             -- hip_reconfig_clk
			hip_reconfig_rst_n     : in  std_logic                       := 'X';             -- hip_reconfig_rst_n
			hip_reconfig_address   : in  std_logic_vector(9 downto 0)    := (others => 'X'); -- hip_reconfig_address
			hip_reconfig_read      : in  std_logic                       := 'X';             -- hip_reconfig_read
			hip_reconfig_write     : in  std_logic                       := 'X';             -- hip_reconfig_write
			hip_reconfig_writedata : in  std_logic_vector(15 downto 0)   := (others => 'X'); -- hip_reconfig_writedata
			hip_reconfig_byte_en   : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- hip_reconfig_byte_en
			ser_shift_load         : in  std_logic                       := 'X';             -- ser_shift_load
			interface_sel          : in  std_logic                       := 'X';             -- interface_sel
			cfgbp_link2csr         : in  std_logic_vector(12 downto 0)   := (others => 'X'); -- cfgbp_link2csr
			cfgbp_comclk_reg       : in  std_logic                       := 'X';             -- cfgbp_comclk_reg
			cfgbp_extsy_reg        : in  std_logic                       := 'X';             -- cfgbp_extsy_reg
			cfgbp_max_pload        : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- cfgbp_max_pload
			cfgbp_tx_ecrcgen       : in  std_logic                       := 'X';             -- cfgbp_tx_ecrcgen
			cfgbp_rx_ecrchk        : in  std_logic                       := 'X';             -- cfgbp_rx_ecrchk
			cfgbp_secbus           : in  std_logic_vector(7 downto 0)    := (others => 'X'); -- cfgbp_secbus
			cfgbp_linkcsr_bit0     : in  std_logic                       := 'X';             -- cfgbp_linkcsr_bit0
			cfgbp_tx_req_pm        : in  std_logic                       := 'X';             -- cfgbp_tx_req_pm
			cfgbp_tx_typ_pm        : in  std_logic_vector(2 downto 0)    := (others => 'X'); -- cfgbp_tx_typ_pm
			cfgbp_req_phypm        : in  std_logic_vector(3 downto 0)    := (others => 'X'); -- cfgbp_req_phypm
			cfgbp_req_phycfg       : in  std_logic_vector(3 downto 0)    := (others => 'X'); -- cfgbp_req_phycfg
			cfgbp_vc0_tcmap_pld    : in  std_logic_vector(6 downto 0)    := (others => 'X'); -- cfgbp_vc0_tcmap_pld
			cfgbp_inh_dllp         : in  std_logic                       := 'X';             -- cfgbp_inh_dllp
			cfgbp_inh_tx_tlp       : in  std_logic                       := 'X';             -- cfgbp_inh_tx_tlp
			cfgbp_req_wake         : in  std_logic                       := 'X';             -- cfgbp_req_wake
			cfgbp_link3_ctl        : in  std_logic_vector(1 downto 0)    := (others => 'X'); -- cfgbp_link3_ctl
			reservedin             : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- reservedin
			tlbfm_in               : out std_logic_vector(1000 downto 0);                    -- tlbfm_in
			tlbfm_out              : in  std_logic_vector(1000 downto 0) := (others => 'X'); -- tlbfm_out
			rxfc_cplbuf_ovf        : out std_logic                                           -- rxfc_cplbuf_ovf
		);
	end component altpcie_sv_hip_ast_hwtcl;

	component altpcie_reconfig_driver is
		generic (
			INTENDED_DEVICE_FAMILY        : string  := "Stratix V";
			gen123_lane_rate_mode_hwtcl   : string  := "Gen1 (2.5 Gbps)";
			number_of_reconfig_interfaces : integer := 2
		);
		port (
			reconfig_xcvr_clk         : in  std_logic                     := 'X';             -- clk
			reconfig_xcvr_rst         : in  std_logic                     := 'X';             -- reset
			reconfig_mgmt_address     : out std_logic_vector(6 downto 0);                     -- address
			reconfig_mgmt_read        : out std_logic;                                        -- read
			reconfig_mgmt_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			reconfig_mgmt_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			reconfig_mgmt_write       : out std_logic;                                        -- write
			reconfig_mgmt_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			currentspeed              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- currentspeed
			reconfig_busy             : in  std_logic                     := 'X';             -- reconfig_busy
			pld_clk                   : in  std_logic                     := 'X';             -- clk
			derr_cor_ext_rcv_drv      : in  std_logic                     := 'X';             -- derr_cor_ext_rcv
			derr_cor_ext_rpl_drv      : in  std_logic                     := 'X';             -- derr_cor_ext_rpl
			derr_rpl_drv              : in  std_logic                     := 'X';             -- derr_rpl
			dlup_exit_drv             : in  std_logic                     := 'X';             -- dlup_exit
			ev128ns_drv               : in  std_logic                     := 'X';             -- ev128ns
			ev1us_drv                 : in  std_logic                     := 'X';             -- ev1us
			hotrst_exit_drv           : in  std_logic                     := 'X';             -- hotrst_exit
			int_status_drv            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- int_status
			l2_exit_drv               : in  std_logic                     := 'X';             -- l2_exit
			lane_act_drv              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- lane_act
			ltssmstate_drv            : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- ltssmstate
			dlup_drv                  : in  std_logic                     := 'X';             -- dlup
			rx_par_err_drv            : in  std_logic                     := 'X';             -- rx_par_err
			tx_par_err_drv            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- tx_par_err
			cfg_par_err_drv           : in  std_logic                     := 'X';             -- cfg_par_err
			ko_cpl_spc_header_drv     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- ko_cpl_spc_header
			ko_cpl_spc_data_drv       : in  std_logic_vector(11 downto 0) := (others => 'X'); -- ko_cpl_spc_data
			cal_busy_in               : out std_logic                                         -- cal_busy_in
		);
	end component altpcie_reconfig_driver;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal pcie_reconfig_driver_0_reconfig_mgmt_readdata         : std_logic_vector(31 downto 0);  -- alt_xcvr_reconfig_0:reconfig_mgmt_readdata -> pcie_reconfig_driver_0:reconfig_mgmt_readdata
	signal pcie_reconfig_driver_0_reconfig_mgmt_waitrequest      : std_logic;                      -- alt_xcvr_reconfig_0:reconfig_mgmt_waitrequest -> pcie_reconfig_driver_0:reconfig_mgmt_waitrequest
	signal pcie_reconfig_driver_0_reconfig_mgmt_address          : std_logic_vector(6 downto 0);   -- pcie_reconfig_driver_0:reconfig_mgmt_address -> alt_xcvr_reconfig_0:reconfig_mgmt_address
	signal pcie_reconfig_driver_0_reconfig_mgmt_read             : std_logic;                      -- pcie_reconfig_driver_0:reconfig_mgmt_read -> alt_xcvr_reconfig_0:reconfig_mgmt_read
	signal pcie_reconfig_driver_0_reconfig_mgmt_write            : std_logic;                      -- pcie_reconfig_driver_0:reconfig_mgmt_write -> alt_xcvr_reconfig_0:reconfig_mgmt_write
	signal pcie_reconfig_driver_0_reconfig_mgmt_writedata        : std_logic_vector(31 downto 0);  -- pcie_reconfig_driver_0:reconfig_mgmt_writedata -> alt_xcvr_reconfig_0:reconfig_mgmt_writedata
	signal hip_hip_currentspeed_currentspeed                     : std_logic_vector(1 downto 0);   -- hip:currentspeed -> pcie_reconfig_driver_0:currentspeed
	signal alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy       : std_logic;                      -- alt_xcvr_reconfig_0:reconfig_busy -> pcie_reconfig_driver_0:reconfig_busy
	signal hip_reconfig_from_xcvr_reconfig_from_xcvr             : std_logic_vector(505 downto 0); -- hip:reconfig_from_xcvr -> alt_xcvr_reconfig_0:reconfig_from_xcvr
	signal alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr : std_logic_vector(769 downto 0); -- alt_xcvr_reconfig_0:reconfig_to_xcvr -> hip:reconfig_to_xcvr
	signal rst_controller_reset_out_reset                        : std_logic;                      -- rst_controller:reset_out -> [alt_xcvr_reconfig_0:mgmt_rst_reset, pcie_reconfig_driver_0:reconfig_xcvr_rst]
	signal local_pcie_perstn_reset_n_ports_inv                   : std_logic;                      -- local_pcie_perstn_reset_n:inv -> rst_controller:reset_in0

begin

	alt_xcvr_reconfig_0 : component alt_xcvr_reconfig
		generic map (
			device_family                 => "Stratix V",
			number_of_reconfig_interfaces => 11,
			enable_offset                 => 1,
			enable_lc                     => 1,
			enable_dcd                    => 0,
			enable_dcd_power_up           => 1,
			enable_analog                 => 0,
			enable_eyemon                 => 0,
			enable_ber                    => 0,
			enable_dfe                    => 0,
			enable_adce                   => 1,
			enable_mif                    => 0,
			enable_pll                    => 0
		)
		port map (
			reconfig_busy             => alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy,       --      reconfig_busy.reconfig_busy
			mgmt_clk_clk              => pcie_ref_clk_clk,                                      --       mgmt_clk_clk.clk
			mgmt_rst_reset            => rst_controller_reset_out_reset,                        --     mgmt_rst_reset.reset
			reconfig_mgmt_address     => pcie_reconfig_driver_0_reconfig_mgmt_address,          --      reconfig_mgmt.address
			reconfig_mgmt_read        => pcie_reconfig_driver_0_reconfig_mgmt_read,             --                   .read
			reconfig_mgmt_readdata    => pcie_reconfig_driver_0_reconfig_mgmt_readdata,         --                   .readdata
			reconfig_mgmt_waitrequest => pcie_reconfig_driver_0_reconfig_mgmt_waitrequest,      --                   .waitrequest
			reconfig_mgmt_write       => pcie_reconfig_driver_0_reconfig_mgmt_write,            --                   .write
			reconfig_mgmt_writedata   => pcie_reconfig_driver_0_reconfig_mgmt_writedata,        --                   .writedata
			reconfig_to_xcvr          => alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr, --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr        => hip_reconfig_from_xcvr_reconfig_from_xcvr,             -- reconfig_from_xcvr.reconfig_from_xcvr
			tx_cal_busy               => open,                                                  --        (terminated)
			rx_cal_busy               => open,                                                  --        (terminated)
			cal_busy_in               => '0',                                                   --        (terminated)
			reconfig_mif_address      => open,                                                  --        (terminated)
			reconfig_mif_read         => open,                                                  --        (terminated)
			reconfig_mif_readdata     => "0000000000000000",                                    --        (terminated)
			reconfig_mif_waitrequest  => '0'                                                    --        (terminated)
		);

	hip : component altpcie_sv_hip_ast_hwtcl
		generic map (
			ACDS_VERSION_HWTCL                       => "15.1",
			lane_mask_hwtcl                          => "x8",
			gen123_lane_rate_mode_hwtcl              => "Gen3 (8.0 Gbps)",
			port_type_hwtcl                          => "Native endpoint",
			pcie_spec_version_hwtcl                  => "3.0",
			ast_width_hwtcl                          => "Avalon-ST 256-bit",
			pll_refclk_freq_hwtcl                    => "100 MHz",
			set_pld_clk_x1_625MHz_hwtcl              => 0,
			use_ast_parity                           => 1,
			multiple_packets_per_cycle_hwtcl         => 0,
			in_cvp_mode_hwtcl                        => 0,
			use_pci_ext_hwtcl                        => 1,
			use_pcie_ext_hwtcl                       => 1,
			use_config_bypass_hwtcl                  => 0,
			enable_tl_only_sim_hwtcl                 => 0,
			hip_reconfig_hwtcl                       => 0,
			hip_tag_checking_hwtcl                   => 1,
			enable_power_on_rst_pulse_hwtcl          => 0,
			enable_pcisigtest_hwtcl                  => 0,
			bar0_size_mask_hwtcl                     => 28,
			bar0_io_space_hwtcl                      => "Disabled",
			bar0_64bit_mem_space_hwtcl               => "Enabled",
			bar0_prefetchable_hwtcl                  => "Enabled",
			bar1_size_mask_hwtcl                     => 0,
			bar1_io_space_hwtcl                      => "Disabled",
			bar1_prefetchable_hwtcl                  => "Disabled",
			bar2_size_mask_hwtcl                     => 17,
			bar2_io_space_hwtcl                      => "Disabled",
			bar2_64bit_mem_space_hwtcl               => "Enabled",
			bar2_prefetchable_hwtcl                  => "Enabled",
			bar3_size_mask_hwtcl                     => 0,
			bar3_io_space_hwtcl                      => "Disabled",
			bar3_prefetchable_hwtcl                  => "Disabled",
			bar4_size_mask_hwtcl                     => 48,
			bar4_io_space_hwtcl                      => "Disabled",
			bar4_64bit_mem_space_hwtcl               => "Enabled",
			bar4_prefetchable_hwtcl                  => "Enabled",
			bar5_size_mask_hwtcl                     => 0,
			bar5_io_space_hwtcl                      => "Disabled",
			bar5_prefetchable_hwtcl                  => "Disabled",
			expansion_base_address_register_hwtcl    => 0,
			io_window_addr_width_hwtcl               => 0,
			prefetchable_mem_window_addr_width_hwtcl => 0,
			vendor_id_hwtcl                          => 4116,
			device_id_hwtcl                          => 1143,
			revision_id_hwtcl                        => 1,
			class_code_hwtcl                         => 1179648,
			subsystem_vendor_id_hwtcl                => 4116,
			subsystem_device_id_hwtcl                => 1199,
			max_payload_size_hwtcl                   => 256,
			extend_tag_field_hwtcl                   => "32",
			completion_timeout_hwtcl                 => "ABCD",
			enable_completion_timeout_disable_hwtcl  => 1,
			use_aer_hwtcl                            => 1,
			ecrc_check_capable_hwtcl                 => 0,
			ecrc_gen_capable_hwtcl                   => 0,
			use_crc_forwarding_hwtcl                 => 0,
			port_link_number_hwtcl                   => 1,
			dll_active_report_support_hwtcl          => 0,
			surprise_down_error_support_hwtcl        => 0,
			slotclkcfg_hwtcl                         => 1,
			msi_multi_message_capable_hwtcl          => "4",
			msi_64bit_addressing_capable_hwtcl       => "true",
			msi_masking_capable_hwtcl                => "false",
			msi_support_hwtcl                        => "true",
			enable_function_msix_support_hwtcl       => 0,
			msix_table_size_hwtcl                    => 0,
			msix_table_offset_hwtcl                  => "0",
			msix_table_bir_hwtcl                     => 0,
			msix_pba_offset_hwtcl                    => "0",
			msix_pba_bir_hwtcl                       => 0,
			enable_slot_register_hwtcl               => 0,
			slot_power_scale_hwtcl                   => 0,
			slot_power_limit_hwtcl                   => 0,
			slot_number_hwtcl                        => 0,
			endpoint_l0_latency_hwtcl                => 0,
			endpoint_l1_latency_hwtcl                => 0,
			vsec_id_hwtcl                            => 0,
			user_id_hwtcl                            => 0,
			vsec_rev_hwtcl                           => 0,
			millisecond_cycle_count_hwtcl            => 248500,
			port_width_be_hwtcl                      => 32,
			port_width_data_hwtcl                    => 256,
			gen3_dcbal_en_hwtcl                      => 1,
			enable_pipe32_sim_hwtcl                  => 0,
			fixed_preset_on                          => 0,
			bypass_cdc_hwtcl                         => "false",
			enable_rx_buffer_checking_hwtcl          => "false",
			disable_link_x2_support_hwtcl            => "false",
			wrong_device_id_hwtcl                    => "disable",
			data_pack_rx_hwtcl                       => "disable",
			ltssm_1ms_timeout_hwtcl                  => "disable",
			ltssm_freqlocked_check_hwtcl             => "disable",
			deskew_comma_hwtcl                       => "skp_eieos_deskw",
			device_number_hwtcl                      => 0,
			pipex1_debug_sel_hwtcl                   => "disable",
			pclk_out_sel_hwtcl                       => "pclk",
			no_soft_reset_hwtcl                      => "false",
			maximum_current_hwtcl                    => 0,
			d1_support_hwtcl                         => "false",
			d2_support_hwtcl                         => "false",
			d0_pme_hwtcl                             => "false",
			d1_pme_hwtcl                             => "false",
			d2_pme_hwtcl                             => "false",
			d3_hot_pme_hwtcl                         => "false",
			d3_cold_pme_hwtcl                        => "false",
			low_priority_vc_hwtcl                    => "single_vc",
			disable_snoop_packet_hwtcl               => "false",
			enable_l1_aspm_hwtcl                     => "false",
			rx_ei_l0s_hwtcl                          => 0,
			enable_l0s_aspm_hwtcl                    => "false",
			aspm_config_management_hwtcl             => "true",
			l1_exit_latency_sameclock_hwtcl          => 0,
			l1_exit_latency_diffclock_hwtcl          => 0,
			hot_plug_support_hwtcl                   => 0,
			extended_tag_reset_hwtcl                 => "false",
			no_command_completed_hwtcl               => "false",
			interrupt_pin_hwtcl                      => "inta",
			bridge_port_vga_enable_hwtcl             => "false",
			bridge_port_ssid_support_hwtcl           => "false",
			ssvid_hwtcl                              => 0,
			ssid_hwtcl                               => 0,
			eie_before_nfts_count_hwtcl              => 4,
			gen2_diffclock_nfts_count_hwtcl          => 255,
			gen2_sameclock_nfts_count_hwtcl          => 255,
			l0_exit_latency_sameclock_hwtcl          => 6,
			l0_exit_latency_diffclock_hwtcl          => 6,
			atomic_op_routing_hwtcl                  => "false",
			atomic_op_completer_32bit_hwtcl          => "false",
			atomic_op_completer_64bit_hwtcl          => "false",
			cas_completer_128bit_hwtcl               => "false",
			ltr_mechanism_hwtcl                      => "false",
			tph_completer_hwtcl                      => "false",
			extended_format_field_hwtcl              => "false",
			atomic_malformed_hwtcl                   => "true",
			flr_capability_hwtcl                     => "false",
			enable_adapter_half_rate_mode_hwtcl      => "false",
			vc0_clk_enable_hwtcl                     => "true",
			register_pipe_signals_hwtcl              => "false",
			skp_os_gen3_count_hwtcl                  => 0,
			tx_cdc_almost_empty_hwtcl                => 5,
			rx_l0s_count_idl_hwtcl                   => 0,
			cdc_dummy_insert_limit_hwtcl             => 11,
			ei_delay_powerdown_count_hwtcl           => 10,
			skp_os_schedule_count_hwtcl              => 0,
			fc_init_timer_hwtcl                      => 1024,
			l01_entry_latency_hwtcl                  => 31,
			flow_control_update_count_hwtcl          => 30,
			flow_control_timeout_count_hwtcl         => 200,
			retry_buffer_last_active_address_hwtcl   => 2047,
			reserved_debug_hwtcl                     => 0,
			bypass_clk_switch_hwtcl                  => "true",
			l2_async_logic_hwtcl                     => "disable",
			indicator_hwtcl                          => 0,
			diffclock_nfts_count_hwtcl               => 128,
			sameclock_nfts_count_hwtcl               => 128,
			rx_cdc_almost_full_hwtcl                 => 12,
			tx_cdc_almost_full_hwtcl                 => 11,
			credit_buffer_allocation_aux_hwtcl       => "absolute",
			vc0_rx_flow_ctrl_posted_header_hwtcl     => 58,
			vc0_rx_flow_ctrl_posted_data_hwtcl       => 882,
			vc0_rx_flow_ctrl_nonposted_header_hwtcl  => 52,
			vc0_rx_flow_ctrl_nonposted_data_hwtcl    => 0,
			vc0_rx_flow_ctrl_compl_header_hwtcl      => 0,
			vc0_rx_flow_ctrl_compl_data_hwtcl        => 0,
			cpl_spc_header_hwtcl                     => 16,
			cpl_spc_data_hwtcl                       => 16,
			gen3_rxfreqlock_counter_hwtcl            => 0,
			gen3_skip_ph2_ph3_hwtcl                  => 0,
			g3_bypass_equlz_hwtcl                    => 0,
			cvp_data_compressed_hwtcl                => "false",
			cvp_data_encrypted_hwtcl                 => "false",
			cvp_mode_reset_hwtcl                     => "false",
			cvp_clk_reset_hwtcl                      => "false",
			cseb_cpl_status_during_cvp_hwtcl         => "config_retry_status",
			core_clk_sel_hwtcl                       => "pld_clk",
			cvp_rate_sel_hwtcl                       => "full_rate",
			g3_dis_rx_use_prst_hwtcl                 => "true",
			g3_dis_rx_use_prst_ep_hwtcl              => "true",
			deemphasis_enable_hwtcl                  => "false",
			reconfig_to_xcvr_width                   => 770,
			reconfig_from_xcvr_width                 => 506,
			single_rx_detect_hwtcl                   => 0,
			hip_hard_reset_hwtcl                     => 0,
			use_cvp_update_core_pof_hwtcl            => 0,
			pcie_inspector_hwtcl                     => 0,
			tlp_inspector_hwtcl                      => 0,
			tlp_inspector_use_signal_probe_hwtcl     => 0,
			tlp_insp_trg_dw0_hwtcl                   => 2049,
			tlp_insp_trg_dw1_hwtcl                   => 0,
			tlp_insp_trg_dw2_hwtcl                   => 0,
			tlp_insp_trg_dw3_hwtcl                   => 0,
			hwtcl_override_g2_txvod                  => 0,
			rpre_emph_a_val_hwtcl                    => 9,
			rpre_emph_b_val_hwtcl                    => 0,
			rpre_emph_c_val_hwtcl                    => 16,
			rpre_emph_d_val_hwtcl                    => 11,
			rpre_emph_e_val_hwtcl                    => 5,
			rvod_sel_a_val_hwtcl                     => 42,
			rvod_sel_b_val_hwtcl                     => 38,
			rvod_sel_c_val_hwtcl                     => 38,
			rvod_sel_d_val_hwtcl                     => 38,
			rvod_sel_e_val_hwtcl                     => 15,
			hwtcl_override_g3rxcoef                  => 0,
			gen3_coeff_1_hwtcl                       => 7,
			gen3_coeff_1_sel_hwtcl                   => "preset_1",
			gen3_coeff_1_preset_hint_hwtcl           => 0,
			gen3_coeff_1_nxtber_more_ptr_hwtcl       => 1,
			gen3_coeff_1_nxtber_more_hwtcl           => "g3_coeff_1_nxtber_more",
			gen3_coeff_1_nxtber_less_ptr_hwtcl       => 1,
			gen3_coeff_1_nxtber_less_hwtcl           => "g3_coeff_1_nxtber_less",
			gen3_coeff_1_reqber_hwtcl                => 0,
			gen3_coeff_1_ber_meas_hwtcl              => 2,
			gen3_coeff_2_hwtcl                       => 0,
			gen3_coeff_2_sel_hwtcl                   => "preset_2",
			gen3_coeff_2_preset_hint_hwtcl           => 0,
			gen3_coeff_2_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_2_nxtber_more_hwtcl           => "g3_coeff_2_nxtber_more",
			gen3_coeff_2_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_2_nxtber_less_hwtcl           => "g3_coeff_2_nxtber_less",
			gen3_coeff_2_reqber_hwtcl                => 0,
			gen3_coeff_2_ber_meas_hwtcl              => 0,
			gen3_coeff_3_hwtcl                       => 0,
			gen3_coeff_3_sel_hwtcl                   => "preset_3",
			gen3_coeff_3_preset_hint_hwtcl           => 0,
			gen3_coeff_3_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_3_nxtber_more_hwtcl           => "g3_coeff_3_nxtber_more",
			gen3_coeff_3_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_3_nxtber_less_hwtcl           => "g3_coeff_3_nxtber_less",
			gen3_coeff_3_reqber_hwtcl                => 0,
			gen3_coeff_3_ber_meas_hwtcl              => 0,
			gen3_coeff_4_hwtcl                       => 0,
			gen3_coeff_4_sel_hwtcl                   => "preset_4",
			gen3_coeff_4_preset_hint_hwtcl           => 0,
			gen3_coeff_4_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_4_nxtber_more_hwtcl           => "g3_coeff_4_nxtber_more",
			gen3_coeff_4_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_4_nxtber_less_hwtcl           => "g3_coeff_4_nxtber_less",
			gen3_coeff_4_reqber_hwtcl                => 0,
			gen3_coeff_4_ber_meas_hwtcl              => 0,
			gen3_coeff_5_hwtcl                       => 0,
			gen3_coeff_5_sel_hwtcl                   => "preset_5",
			gen3_coeff_5_preset_hint_hwtcl           => 0,
			gen3_coeff_5_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_5_nxtber_more_hwtcl           => "g3_coeff_5_nxtber_more",
			gen3_coeff_5_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_5_nxtber_less_hwtcl           => "g3_coeff_5_nxtber_less",
			gen3_coeff_5_reqber_hwtcl                => 0,
			gen3_coeff_5_ber_meas_hwtcl              => 0,
			gen3_coeff_6_hwtcl                       => 0,
			gen3_coeff_6_sel_hwtcl                   => "preset_6",
			gen3_coeff_6_preset_hint_hwtcl           => 0,
			gen3_coeff_6_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_6_nxtber_more_hwtcl           => "g3_coeff_6_nxtber_more",
			gen3_coeff_6_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_6_nxtber_less_hwtcl           => "g3_coeff_6_nxtber_less",
			gen3_coeff_6_reqber_hwtcl                => 0,
			gen3_coeff_6_ber_meas_hwtcl              => 0,
			gen3_coeff_7_hwtcl                       => 0,
			gen3_coeff_7_sel_hwtcl                   => "preset_7",
			gen3_coeff_7_preset_hint_hwtcl           => 0,
			gen3_coeff_7_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_7_nxtber_more_hwtcl           => "g3_coeff_7_nxtber_more",
			gen3_coeff_7_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_7_nxtber_less_hwtcl           => "g3_coeff_7_nxtber_less",
			gen3_coeff_7_reqber_hwtcl                => 0,
			gen3_coeff_7_ber_meas_hwtcl              => 0,
			gen3_coeff_8_hwtcl                       => 0,
			gen3_coeff_8_sel_hwtcl                   => "preset_8",
			gen3_coeff_8_preset_hint_hwtcl           => 0,
			gen3_coeff_8_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_8_nxtber_more_hwtcl           => "g3_coeff_8_nxtber_more",
			gen3_coeff_8_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_8_nxtber_less_hwtcl           => "g3_coeff_8_nxtber_less",
			gen3_coeff_8_reqber_hwtcl                => 0,
			gen3_coeff_8_ber_meas_hwtcl              => 0,
			gen3_coeff_9_hwtcl                       => 0,
			gen3_coeff_9_sel_hwtcl                   => "preset_9",
			gen3_coeff_9_preset_hint_hwtcl           => 0,
			gen3_coeff_9_nxtber_more_ptr_hwtcl       => 0,
			gen3_coeff_9_nxtber_more_hwtcl           => "g3_coeff_9_nxtber_more",
			gen3_coeff_9_nxtber_less_ptr_hwtcl       => 0,
			gen3_coeff_9_nxtber_less_hwtcl           => "g3_coeff_9_nxtber_less",
			gen3_coeff_9_reqber_hwtcl                => 0,
			gen3_coeff_9_ber_meas_hwtcl              => 0,
			gen3_coeff_10_hwtcl                      => 0,
			gen3_coeff_10_sel_hwtcl                  => "preset_10",
			gen3_coeff_10_preset_hint_hwtcl          => 0,
			gen3_coeff_10_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_10_nxtber_more_hwtcl          => "g3_coeff_10_nxtber_more",
			gen3_coeff_10_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_10_nxtber_less_hwtcl          => "g3_coeff_10_nxtber_less",
			gen3_coeff_10_reqber_hwtcl               => 0,
			gen3_coeff_10_ber_meas_hwtcl             => 0,
			gen3_coeff_11_hwtcl                      => 0,
			gen3_coeff_11_sel_hwtcl                  => "preset_11",
			gen3_coeff_11_preset_hint_hwtcl          => 0,
			gen3_coeff_11_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_11_nxtber_more_hwtcl          => "g3_coeff_11_nxtber_more",
			gen3_coeff_11_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_11_nxtber_less_hwtcl          => "g3_coeff_11_nxtber_less",
			gen3_coeff_11_reqber_hwtcl               => 0,
			gen3_coeff_11_ber_meas_hwtcl             => 0,
			gen3_coeff_12_hwtcl                      => 0,
			gen3_coeff_12_sel_hwtcl                  => "preset_12",
			gen3_coeff_12_preset_hint_hwtcl          => 0,
			gen3_coeff_12_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_12_nxtber_more_hwtcl          => "g3_coeff_12_nxtber_more",
			gen3_coeff_12_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_12_nxtber_less_hwtcl          => "g3_coeff_12_nxtber_less",
			gen3_coeff_12_reqber_hwtcl               => 0,
			gen3_coeff_12_ber_meas_hwtcl             => 0,
			gen3_coeff_13_hwtcl                      => 0,
			gen3_coeff_13_sel_hwtcl                  => "preset_13",
			gen3_coeff_13_preset_hint_hwtcl          => 0,
			gen3_coeff_13_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_13_nxtber_more_hwtcl          => "g3_coeff_13_nxtber_more",
			gen3_coeff_13_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_13_nxtber_less_hwtcl          => "g3_coeff_13_nxtber_less",
			gen3_coeff_13_reqber_hwtcl               => 0,
			gen3_coeff_13_ber_meas_hwtcl             => 0,
			gen3_coeff_14_hwtcl                      => 0,
			gen3_coeff_14_sel_hwtcl                  => "preset_14",
			gen3_coeff_14_preset_hint_hwtcl          => 0,
			gen3_coeff_14_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_14_nxtber_more_hwtcl          => "g3_coeff_14_nxtber_more",
			gen3_coeff_14_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_14_nxtber_less_hwtcl          => "g3_coeff_14_nxtber_less",
			gen3_coeff_14_reqber_hwtcl               => 0,
			gen3_coeff_14_ber_meas_hwtcl             => 0,
			gen3_coeff_15_hwtcl                      => 0,
			gen3_coeff_15_sel_hwtcl                  => "preset_15",
			gen3_coeff_15_preset_hint_hwtcl          => 0,
			gen3_coeff_15_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_15_nxtber_more_hwtcl          => "g3_coeff_15_nxtber_more",
			gen3_coeff_15_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_15_nxtber_less_hwtcl          => "g3_coeff_15_nxtber_less",
			gen3_coeff_15_reqber_hwtcl               => 0,
			gen3_coeff_15_ber_meas_hwtcl             => 0,
			gen3_coeff_16_hwtcl                      => 0,
			gen3_coeff_16_sel_hwtcl                  => "preset_16",
			gen3_coeff_16_preset_hint_hwtcl          => 0,
			gen3_coeff_16_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_16_nxtber_more_hwtcl          => "g3_coeff_16_nxtber_more",
			gen3_coeff_16_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_16_nxtber_less_hwtcl          => "g3_coeff_16_nxtber_less",
			gen3_coeff_16_reqber_hwtcl               => 0,
			gen3_coeff_16_ber_meas_hwtcl             => 0,
			gen3_coeff_17_hwtcl                      => 0,
			gen3_coeff_17_sel_hwtcl                  => "preset_17",
			gen3_coeff_17_preset_hint_hwtcl          => 0,
			gen3_coeff_17_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_17_nxtber_more_hwtcl          => "g3_coeff_17_nxtber_more",
			gen3_coeff_17_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_17_nxtber_less_hwtcl          => "g3_coeff_17_nxtber_less",
			gen3_coeff_17_reqber_hwtcl               => 0,
			gen3_coeff_17_ber_meas_hwtcl             => 0,
			gen3_coeff_18_hwtcl                      => 0,
			gen3_coeff_18_sel_hwtcl                  => "preset_18",
			gen3_coeff_18_preset_hint_hwtcl          => 0,
			gen3_coeff_18_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_18_nxtber_more_hwtcl          => "g3_coeff_18_nxtber_more",
			gen3_coeff_18_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_18_nxtber_less_hwtcl          => "g3_coeff_18_nxtber_less",
			gen3_coeff_18_reqber_hwtcl               => 0,
			gen3_coeff_18_ber_meas_hwtcl             => 0,
			gen3_coeff_19_hwtcl                      => 0,
			gen3_coeff_19_sel_hwtcl                  => "preset_19",
			gen3_coeff_19_preset_hint_hwtcl          => 0,
			gen3_coeff_19_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_19_nxtber_more_hwtcl          => "g3_coeff_19_nxtber_more",
			gen3_coeff_19_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_19_nxtber_less_hwtcl          => "g3_coeff_19_nxtber_less",
			gen3_coeff_19_reqber_hwtcl               => 0,
			gen3_coeff_19_ber_meas_hwtcl             => 0,
			gen3_coeff_20_hwtcl                      => 0,
			gen3_coeff_20_sel_hwtcl                  => "preset_20",
			gen3_coeff_20_preset_hint_hwtcl          => 0,
			gen3_coeff_20_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_20_nxtber_more_hwtcl          => "g3_coeff_20_nxtber_more",
			gen3_coeff_20_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_20_nxtber_less_hwtcl          => "g3_coeff_20_nxtber_less",
			gen3_coeff_20_reqber_hwtcl               => 0,
			gen3_coeff_20_ber_meas_hwtcl             => 0,
			gen3_coeff_21_hwtcl                      => 0,
			gen3_coeff_21_sel_hwtcl                  => "preset_21",
			gen3_coeff_21_preset_hint_hwtcl          => 0,
			gen3_coeff_21_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_21_nxtber_more_hwtcl          => "g3_coeff_21_nxtber_more",
			gen3_coeff_21_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_21_nxtber_less_hwtcl          => "g3_coeff_21_nxtber_less",
			gen3_coeff_21_reqber_hwtcl               => 0,
			gen3_coeff_21_ber_meas_hwtcl             => 0,
			gen3_coeff_22_hwtcl                      => 0,
			gen3_coeff_22_sel_hwtcl                  => "preset_22",
			gen3_coeff_22_preset_hint_hwtcl          => 0,
			gen3_coeff_22_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_22_nxtber_more_hwtcl          => "g3_coeff_22_nxtber_more",
			gen3_coeff_22_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_22_nxtber_less_hwtcl          => "g3_coeff_22_nxtber_less",
			gen3_coeff_22_reqber_hwtcl               => 0,
			gen3_coeff_22_ber_meas_hwtcl             => 0,
			gen3_coeff_23_hwtcl                      => 0,
			gen3_coeff_23_sel_hwtcl                  => "preset_23",
			gen3_coeff_23_preset_hint_hwtcl          => 0,
			gen3_coeff_23_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_23_nxtber_more_hwtcl          => "g3_coeff_23_nxtber_more",
			gen3_coeff_23_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_23_nxtber_less_hwtcl          => "g3_coeff_23_nxtber_less",
			gen3_coeff_23_reqber_hwtcl               => 0,
			gen3_coeff_23_ber_meas_hwtcl             => 0,
			gen3_coeff_24_hwtcl                      => 0,
			gen3_coeff_24_sel_hwtcl                  => "preset_24",
			gen3_coeff_24_preset_hint_hwtcl          => 0,
			gen3_coeff_24_nxtber_more_ptr_hwtcl      => 0,
			gen3_coeff_24_nxtber_more_hwtcl          => "g3_coeff_24_nxtber_more",
			gen3_coeff_24_nxtber_less_ptr_hwtcl      => 0,
			gen3_coeff_24_nxtber_less_hwtcl          => "g3_coeff_24_nxtber_less",
			gen3_coeff_24_reqber_hwtcl               => 0,
			gen3_coeff_24_ber_meas_hwtcl             => 0,
			hwtcl_override_g3txcoef                  => 0,
			gen3_preset_coeff_1_hwtcl                => 0,
			gen3_preset_coeff_2_hwtcl                => 0,
			gen3_preset_coeff_3_hwtcl                => 0,
			gen3_preset_coeff_4_hwtcl                => 0,
			gen3_preset_coeff_5_hwtcl                => 0,
			gen3_preset_coeff_6_hwtcl                => 0,
			gen3_preset_coeff_7_hwtcl                => 0,
			gen3_preset_coeff_8_hwtcl                => 0,
			gen3_preset_coeff_9_hwtcl                => 0,
			gen3_preset_coeff_10_hwtcl               => 0,
			gen3_preset_coeff_11_hwtcl               => 0,
			gen3_low_freq_hwtcl                      => 0,
			full_swing_hwtcl                         => 35,
			gen3_full_swing_hwtcl                    => 35,
			use_atx_pll_hwtcl                        => 0,
			low_latency_mode_hwtcl                   => 1
		)
		port map (
			npor                   => pcie_rstn_npor,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --               npor.npor
			pin_perst              => pcie_rstn_pin_perst,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --                   .pin_perst
			lmi_addr               => hip_lmi_lmi_addr,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                lmi.lmi_addr
			lmi_din                => hip_lmi_lmi_din,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --                   .lmi_din
			lmi_rden               => hip_lmi_lmi_rden,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .lmi_rden
			lmi_wren               => hip_lmi_lmi_wren,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .lmi_wren
			lmi_ack                => hip_lmi_lmi_ack,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --                   .lmi_ack
			lmi_dout               => hip_lmi_lmi_dout,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .lmi_dout
			hpg_ctrler             => hip_config_tl_hpg_ctrler,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --          config_tl.hpg_ctrler
			tl_cfg_add             => hip_config_tl_tl_cfg_add,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .tl_cfg_add
			tl_cfg_ctl             => hip_config_tl_tl_cfg_ctl,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .tl_cfg_ctl
			tl_cfg_sts             => hip_config_tl_tl_cfg_sts,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .tl_cfg_sts
			cpl_err                => hip_config_tl_cpl_err,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       --                   .cpl_err
			cpl_pending            => hip_config_tl_cpl_pending,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .cpl_pending
			pm_auxpwr              => hip_power_mngt_pm_auxpwr,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --         power_mngt.pm_auxpwr
			pm_data                => hip_power_mngt_pm_data,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --                   .pm_data
			pme_to_cr              => hip_power_mngt_pme_to_cr,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .pme_to_cr
			pm_event               => hip_power_mngt_pm_event,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .pm_event
			pme_to_sr              => hip_power_mngt_pme_to_sr,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .pme_to_sr
			rx_st_sop              => hip_rx_st_startofpacket,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --              rx_st.startofpacket
			rx_st_eop              => hip_rx_st_endofpacket,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       --                   .endofpacket
			rx_st_err              => hip_rx_st_error,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --                   .error
			rx_st_valid            => hip_rx_st_valid,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --                   .valid
			rx_st_empty            => hip_rx_st_empty,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --                   .empty
			rx_st_ready            => hip_rx_st_ready,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --                   .ready
			rx_st_data             => hip_rx_st_data,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .data
			rx_st_parity           => hip_rx_st_parity,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .parity
			rx_st_bar              => hip_rx_bar_be_rx_st_bar,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --          rx_bar_be.rx_st_bar
			rx_st_mask             => hip_rx_bar_be_rx_st_mask,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .rx_st_mask
			tx_st_sop              => hip_tx_st_startofpacket,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --              tx_st.startofpacket
			tx_st_eop              => hip_tx_st_endofpacket,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       --                   .endofpacket
			tx_st_err              => hip_tx_st_error,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --                   .error
			tx_st_valid            => hip_tx_st_valid,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --                   .valid
			tx_st_empty            => hip_tx_st_empty,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --                   .empty
			tx_st_ready            => hip_tx_st_ready,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --                   .ready
			tx_st_data             => hip_tx_st_data,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .data
			tx_st_parity           => hip_tx_st_parity,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .parity
			tx_cred_datafccp       => hip_tx_cred_tx_cred_datafccp,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                --            tx_cred.tx_cred_datafccp
			tx_cred_datafcnp       => hip_tx_cred_tx_cred_datafcnp,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                --                   .tx_cred_datafcnp
			tx_cred_datafcp        => hip_tx_cred_tx_cred_datafcp,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .tx_cred_datafcp
			tx_cred_fchipcons      => hip_tx_cred_tx_cred_fchipcons,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --                   .tx_cred_fchipcons
			tx_cred_fcinfinite     => hip_tx_cred_tx_cred_fcinfinite,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .tx_cred_fcinfinite
			tx_cred_hdrfccp        => hip_tx_cred_tx_cred_hdrfccp,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .tx_cred_hdrfccp
			tx_cred_hdrfcnp        => hip_tx_cred_tx_cred_hdrfcnp,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .tx_cred_hdrfcnp
			tx_cred_hdrfcp         => hip_tx_cred_tx_cred_hdrfcp,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .tx_cred_hdrfcp
			pld_clk                => pld_clk_clk,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --            pld_clk.clk
			coreclkout_hip         => hip_coreclkout_hip_clk,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --     coreclkout_hip.clk
			refclk                 => pcie_ref_clk_clk,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --             refclk.clk
			reset_status           => hip_rst_reset_status,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --            hip_rst.reset_status
			serdes_pll_locked      => hip_rst_serdes_pll_locked,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .serdes_pll_locked
			pld_clk_inuse          => hip_rst_pld_clk_inuse,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       --                   .pld_clk_inuse
			pld_core_ready         => hip_rst_pld_core_ready,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --                   .pld_core_ready
			testin_zero            => hip_rst_testin_zero,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --                   .testin_zero
			reconfig_to_xcvr       => alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr     => hip_reconfig_from_xcvr_reconfig_from_xcvr,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   -- reconfig_from_xcvr.reconfig_from_xcvr
			rx_in0                 => hip_serial_rx_in0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --         hip_serial.rx_in0
			rx_in1                 => hip_serial_rx_in1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_in1
			rx_in2                 => hip_serial_rx_in2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_in2
			rx_in3                 => hip_serial_rx_in3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_in3
			rx_in4                 => hip_serial_rx_in4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_in4
			rx_in5                 => hip_serial_rx_in5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_in5
			rx_in6                 => hip_serial_rx_in6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_in6
			rx_in7                 => hip_serial_rx_in7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_in7
			tx_out0                => hip_serial_tx_out0,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .tx_out0
			tx_out1                => hip_serial_tx_out1,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .tx_out1
			tx_out2                => hip_serial_tx_out2,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .tx_out2
			tx_out3                => hip_serial_tx_out3,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .tx_out3
			tx_out4                => hip_serial_tx_out4,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .tx_out4
			tx_out5                => hip_serial_tx_out5,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .tx_out5
			tx_out6                => hip_serial_tx_out6,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .tx_out6
			tx_out7                => hip_serial_tx_out7,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .tx_out7
			sim_pipe_pclk_in       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --           hip_pipe.sim_pipe_pclk_in
			sim_pipe_rate          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .sim_pipe_rate
			sim_ltssmstate         => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .sim_ltssmstate
			eidleinfersel0         => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .eidleinfersel0
			eidleinfersel1         => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .eidleinfersel1
			eidleinfersel2         => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .eidleinfersel2
			eidleinfersel3         => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .eidleinfersel3
			eidleinfersel4         => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .eidleinfersel4
			eidleinfersel5         => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .eidleinfersel5
			eidleinfersel6         => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .eidleinfersel6
			eidleinfersel7         => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .eidleinfersel7
			powerdown0             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .powerdown0
			powerdown1             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .powerdown1
			powerdown2             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .powerdown2
			powerdown3             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .powerdown3
			powerdown4             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .powerdown4
			powerdown5             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .powerdown5
			powerdown6             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .powerdown6
			powerdown7             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .powerdown7
			rxpolarity0            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxpolarity0
			rxpolarity1            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxpolarity1
			rxpolarity2            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxpolarity2
			rxpolarity3            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxpolarity3
			rxpolarity4            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxpolarity4
			rxpolarity5            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxpolarity5
			rxpolarity6            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxpolarity6
			rxpolarity7            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxpolarity7
			txcompl0               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txcompl0
			txcompl1               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txcompl1
			txcompl2               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txcompl2
			txcompl3               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txcompl3
			txcompl4               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txcompl4
			txcompl5               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txcompl5
			txcompl6               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txcompl6
			txcompl7               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txcompl7
			txdata0                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdata0
			txdata1                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdata1
			txdata2                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdata2
			txdata3                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdata3
			txdata4                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdata4
			txdata5                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdata5
			txdata6                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdata6
			txdata7                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdata7
			txdatak0               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdatak0
			txdatak1               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdatak1
			txdatak2               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdatak2
			txdatak3               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdatak3
			txdatak4               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdatak4
			txdatak5               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdatak5
			txdatak6               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdatak6
			txdatak7               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdatak7
			txdetectrx0            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdetectrx0
			txdetectrx1            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdetectrx1
			txdetectrx2            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdetectrx2
			txdetectrx3            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdetectrx3
			txdetectrx4            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdetectrx4
			txdetectrx5            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdetectrx5
			txdetectrx6            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdetectrx6
			txdetectrx7            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdetectrx7
			txelecidle0            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txelecidle0
			txelecidle1            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txelecidle1
			txelecidle2            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txelecidle2
			txelecidle3            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txelecidle3
			txelecidle4            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txelecidle4
			txelecidle5            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txelecidle5
			txelecidle6            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txelecidle6
			txelecidle7            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txelecidle7
			txdeemph0              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdeemph0
			txdeemph1              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdeemph1
			txdeemph2              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdeemph2
			txdeemph3              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdeemph3
			txdeemph4              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdeemph4
			txdeemph5              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdeemph5
			txdeemph6              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdeemph6
			txdeemph7              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txdeemph7
			txmargin0              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txmargin0
			txmargin1              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txmargin1
			txmargin2              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txmargin2
			txmargin3              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txmargin3
			txmargin4              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txmargin4
			txmargin5              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txmargin5
			txmargin6              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txmargin6
			txmargin7              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txmargin7
			txswing0               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txswing0
			txswing1               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txswing1
			txswing2               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txswing2
			txswing3               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txswing3
			txswing4               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txswing4
			txswing5               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txswing5
			txswing6               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txswing6
			txswing7               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .txswing7
			phystatus0             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .phystatus0
			phystatus1             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .phystatus1
			phystatus2             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .phystatus2
			phystatus3             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .phystatus3
			phystatus4             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .phystatus4
			phystatus5             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .phystatus5
			phystatus6             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .phystatus6
			phystatus7             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .phystatus7
			rxdata0                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdata0
			rxdata1                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdata1
			rxdata2                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdata2
			rxdata3                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdata3
			rxdata4                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdata4
			rxdata5                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdata5
			rxdata6                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdata6
			rxdata7                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdata7
			rxdatak0               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdatak0
			rxdatak1               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdatak1
			rxdatak2               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdatak2
			rxdatak3               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdatak3
			rxdatak4               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdatak4
			rxdatak5               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdatak5
			rxdatak6               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdatak6
			rxdatak7               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxdatak7
			rxelecidle0            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxelecidle0
			rxelecidle1            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxelecidle1
			rxelecidle2            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxelecidle2
			rxelecidle3            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxelecidle3
			rxelecidle4            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxelecidle4
			rxelecidle5            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxelecidle5
			rxelecidle6            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxelecidle6
			rxelecidle7            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxelecidle7
			rxstatus0              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxstatus0
			rxstatus1              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxstatus1
			rxstatus2              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxstatus2
			rxstatus3              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxstatus3
			rxstatus4              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxstatus4
			rxstatus5              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxstatus5
			rxstatus6              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxstatus6
			rxstatus7              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxstatus7
			rxvalid0               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxvalid0
			rxvalid1               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxvalid1
			rxvalid2               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxvalid2
			rxvalid3               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxvalid3
			rxvalid4               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxvalid4
			rxvalid5               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxvalid5
			rxvalid6               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxvalid6
			rxvalid7               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .rxvalid7
			app_int_sts            => hip_int_msi_app_int_sts,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --            int_msi.app_int_sts
			app_msi_num            => hip_int_msi_app_msi_num,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .app_msi_num
			app_msi_req            => hip_int_msi_app_msi_req,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .app_msi_req
			app_msi_tc             => hip_int_msi_app_msi_tc,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --                   .app_msi_tc
			app_int_ack            => hip_int_msi_app_int_ack,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .app_int_ack
			app_msi_ack            => hip_int_msi_app_msi_ack,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .app_msi_ack
			cseb_rddata            => hip_cseb_cseb_rddata,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --               cseb.cseb_rddata
			cseb_rdresponse        => hip_cseb_cseb_rdresponse,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .cseb_rdresponse
			cseb_waitrequest       => hip_cseb_cseb_waitrequest,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .cseb_waitrequest
			cseb_wrresponse        => hip_cseb_cseb_wrresponse,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .cseb_wrresponse
			cseb_wrresp_valid      => hip_cseb_cseb_wrresp_valid,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .cseb_wrresp_valid
			cseb_addr              => hip_cseb_cseb_addr,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .cseb_addr
			cseb_be                => hip_cseb_cseb_be,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .cseb_be
			cseb_rden              => hip_cseb_cseb_rden,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .cseb_rden
			cseb_wrdata            => hip_cseb_cseb_wrdata,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .cseb_wrdata
			cseb_wren              => hip_cseb_cseb_wren,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .cseb_wren
			cseb_wrresp_req        => hip_cseb_cseb_wrresp_req,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .cseb_wrresp_req
			cseb_rddata_parity     => hip_cseb_cseb_rddata_parity,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .cseb_rddata_parity
			cseb_addr_parity       => hip_cseb_cseb_addr_parity,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .cseb_addr_parity
			cseb_wrdata_parity     => hip_cseb_cseb_wrdata_parity,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 --                   .cseb_wrdata_parity
			test_in                => hip_ctrl_test_in,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --           hip_ctrl.test_in
			simu_mode_pipe         => hip_ctrl_simu_mode_pipe,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .simu_mode_pipe
			derr_cor_ext_rcv       => hip_hip_status_derr_cor_ext_rcv,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --         hip_status.derr_cor_ext_rcv
			derr_cor_ext_rpl       => hip_hip_status_derr_cor_ext_rpl,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --                   .derr_cor_ext_rpl
			derr_rpl               => hip_hip_status_derr_rpl,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .derr_rpl
			dlup                   => hip_hip_status_dlup,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --                   .dlup
			dlup_exit              => hip_hip_status_dlup_exit,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --                   .dlup_exit
			ev128ns                => hip_hip_status_ev128ns,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --                   .ev128ns
			ev1us                  => hip_hip_status_ev1us,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --                   .ev1us
			hotrst_exit            => hip_hip_status_hotrst_exit,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .hotrst_exit
			int_status             => hip_hip_status_int_status,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .int_status
			l2_exit                => hip_hip_status_l2_exit,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --                   .l2_exit
			lane_act               => hip_hip_status_lane_act,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --                   .lane_act
			ltssmstate             => hip_hip_status_ltssmstate,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .ltssmstate
			rx_par_err             => hip_hip_status_rx_par_err,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .rx_par_err
			tx_par_err             => hip_hip_status_tx_par_err,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --                   .tx_par_err
			cfg_par_err            => hip_hip_status_cfg_par_err,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --                   .cfg_par_err
			ko_cpl_spc_header      => hip_hip_status_ko_cpl_spc_header,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .ko_cpl_spc_header
			ko_cpl_spc_data        => hip_hip_status_ko_cpl_spc_data,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              --                   .ko_cpl_spc_data
			currentspeed           => hip_hip_currentspeed_currentspeed,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --   hip_currentspeed.currentspeed
			rx_st_be               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			tx_cons_cred_sel       => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			sim_pipe_pclk_out      => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxdataskip0            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxdataskip1            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxdataskip2            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxdataskip3            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxdataskip4            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxdataskip5            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxdataskip6            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxdataskip7            => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst0               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst1               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst2               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst3               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst4               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst5               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst6               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxblkst7               => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxsynchd0              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxsynchd1              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxsynchd2              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxsynchd3              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxsynchd4              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxsynchd5              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxsynchd6              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxsynchd7              => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			rxfreqlocked0          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxfreqlocked1          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxfreqlocked2          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxfreqlocked3          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxfreqlocked4          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxfreqlocked5          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxfreqlocked6          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rxfreqlocked7          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			currentcoeff0          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentcoeff1          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentcoeff2          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentcoeff3          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentcoeff4          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentcoeff5          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentcoeff6          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentcoeff7          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset0       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset1       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset2       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset3       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset4       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset5       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset6       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			currentrxpreset7       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd0              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd1              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd2              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd3              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd4              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd5              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd6              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txsynchd7              => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst0               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst1               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst2               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst3               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst4               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst5               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst6               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			txblkst7               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			aer_msi_num            => "00000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --        (terminated)
			pex_msi_num            => "00000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --        (terminated)
			serr_out               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			hip_reconfig_clk       => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			hip_reconfig_rst_n     => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			hip_reconfig_address   => "0000000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                --        (terminated)
			hip_reconfig_read      => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			hip_reconfig_write     => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			hip_reconfig_writedata => "0000000000000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --        (terminated)
			hip_reconfig_byte_en   => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			ser_shift_load         => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			interface_sel          => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_link2csr         => "0000000000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             --        (terminated)
			cfgbp_comclk_reg       => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_extsy_reg        => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_max_pload        => "000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       --        (terminated)
			cfgbp_tx_ecrcgen       => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_rx_ecrchk        => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_secbus           => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --        (terminated)
			cfgbp_linkcsr_bit0     => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_tx_req_pm        => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_tx_typ_pm        => "000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       --        (terminated)
			cfgbp_req_phypm        => "0000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --        (terminated)
			cfgbp_req_phycfg       => "0000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --        (terminated)
			cfgbp_vc0_tcmap_pld    => "0000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --        (terminated)
			cfgbp_inh_dllp         => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_inh_tx_tlp       => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_req_wake         => '0',                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			cfgbp_link3_ctl        => "00",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			reservedin             => "00000000000000000000000000000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --        (terminated)
			tlbfm_in               => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        (terminated)
			tlbfm_out              => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --        (terminated)
			rxfc_cplbuf_ovf        => open                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
		);

	pcie_reconfig_driver_0 : component altpcie_reconfig_driver
		generic map (
			INTENDED_DEVICE_FAMILY        => "Stratix V",
			gen123_lane_rate_mode_hwtcl   => "Gen3 (8.0 Gbps)",
			number_of_reconfig_interfaces => 11
		)
		port map (
			reconfig_xcvr_clk         => pcie_ref_clk_clk,                                 -- reconfig_xcvr_clk.clk
			reconfig_xcvr_rst         => rst_controller_reset_out_reset,                   -- reconfig_xcvr_rst.reset
			reconfig_mgmt_address     => pcie_reconfig_driver_0_reconfig_mgmt_address,     --     reconfig_mgmt.address
			reconfig_mgmt_read        => pcie_reconfig_driver_0_reconfig_mgmt_read,        --                  .read
			reconfig_mgmt_readdata    => pcie_reconfig_driver_0_reconfig_mgmt_readdata,    --                  .readdata
			reconfig_mgmt_waitrequest => pcie_reconfig_driver_0_reconfig_mgmt_waitrequest, --                  .waitrequest
			reconfig_mgmt_write       => pcie_reconfig_driver_0_reconfig_mgmt_write,       --                  .write
			reconfig_mgmt_writedata   => pcie_reconfig_driver_0_reconfig_mgmt_writedata,   --                  .writedata
			currentspeed              => hip_hip_currentspeed_currentspeed,                --  hip_currentspeed.currentspeed
			reconfig_busy             => alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy,  --     reconfig_busy.reconfig_busy
			pld_clk                   => pld_clk_clk,                                      --           pld_clk.clk
			derr_cor_ext_rcv_drv      => rcd_hip_status_derr_cor_ext_rcv,                  --    hip_status_drv.derr_cor_ext_rcv
			derr_cor_ext_rpl_drv      => rcd_hip_status_derr_cor_ext_rpl,                  --                  .derr_cor_ext_rpl
			derr_rpl_drv              => rcd_hip_status_derr_rpl,                          --                  .derr_rpl
			dlup_exit_drv             => rcd_hip_status_dlup_exit,                         --                  .dlup_exit
			ev128ns_drv               => rcd_hip_status_ev128ns,                           --                  .ev128ns
			ev1us_drv                 => rcd_hip_status_ev1us,                             --                  .ev1us
			hotrst_exit_drv           => rcd_hip_status_hotrst_exit,                       --                  .hotrst_exit
			int_status_drv            => rcd_hip_status_int_status,                        --                  .int_status
			l2_exit_drv               => rcd_hip_status_l2_exit,                           --                  .l2_exit
			lane_act_drv              => rcd_hip_status_lane_act,                          --                  .lane_act
			ltssmstate_drv            => rcd_hip_status_ltssmstate,                        --                  .ltssmstate
			dlup_drv                  => rcd_hip_status_dlup,                              --                  .dlup
			rx_par_err_drv            => rcd_hip_status_rx_par_err,                        --                  .rx_par_err
			tx_par_err_drv            => rcd_hip_status_tx_par_err,                        --                  .tx_par_err
			cfg_par_err_drv           => rcd_hip_status_cfg_par_err,                       --                  .cfg_par_err
			ko_cpl_spc_header_drv     => rcd_hip_status_ko_cpl_spc_header,                 --                  .ko_cpl_spc_header
			ko_cpl_spc_data_drv       => rcd_hip_status_ko_cpl_spc_data,                   --                  .ko_cpl_spc_data
			cal_busy_in               => open                                              --       (terminated)
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => local_pcie_perstn_reset_n_ports_inv, -- reset_in0.reset
			clk            => pcie_ref_clk_clk,                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset,      -- reset_out.reset
			reset_req      => open,                                -- (terminated)
			reset_req_in0  => '0',                                 -- (terminated)
			reset_in1      => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_in2      => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	local_pcie_perstn_reset_n_ports_inv <= not local_pcie_perstn_reset_n;

end architecture rtl; -- of pcie_wrap0
