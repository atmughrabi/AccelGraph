// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BnspwXBwrdaKZ7kTG8IgnyZ5/BRqzcLgeBegFzpIEItNKCd5hgkVUyH6JAUM5wuC
dtX795jH93EB/UkiCbb5+wbvBfzF0W9OSk+dglVQOh2AsUTf596aEmZE3/r+UTyv
DZ/PoDN8gvULu+rzWz76ZwVkUgSko0wDuOtskwritec=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12912)
tr5uzeq/bD22O38RkLuXZqYWytTVvzTVMzjaet10H2TJwyW0nLVTP0GbjsElmBh1
VYoqhlE02pH7trk+RqE9LQbOIaA6S5Agah8Li7WxwtVQMSv3BWJHfukoGuB2FzOu
CFcv+76V+kNX4hrx5aynR7fTjDVoGRksfwPfv2JMJnia+pjVlQLgEhIBZlOF2r98
9pnGxYyMYgIba3J+7Uf77Nr+9knlEOAHpdon4CBnKy7zluvFTLHtiEG1Sw4viE5y
QAjKIXz9okhupW0jFpCSnHsYUADYGQ+NkX6Ws5ewf2ek4u1zxIx0X1EYisGUZFKE
eFkpu15rtgSIScZ42DCR3cb6tXzyASVsCowxhsdhoB+iJ7Iq4uWbydksAUq3jbsu
iG3v9OIBQ4NCETEOog1wFJk3rWrVQaG+5kr3E6ddUKVBsy0ErXd2lXdCsjrcNKlj
H2ZfX2vt1v4QXlObtpfLGDQMBbvOx4TEPFWVAPeFSU12U3mXkd9ZcYxf+YKC+K/V
zjPNfDg/n4CTRFo/wr/GJ6ViEDfeUe+NWa2upThcbqYkKLGSs+UWFUVdmDN1ejQg
fQy+7/UhohJXUeprGeHYJct+rY/aszQ9NByiV6AmXnQr52D+BhLy31z9sb2X+tJr
ZVq9wgpZdyOruIY9Eri3TDF7vCt1hRTcmklSwCdWKEBH4Ltx372dxc37Br/Y6j1/
y0O4zbtVL1LzvqemlEhYd4lNEroqQ/mdWm5WdUh+J5zMS+8dZmYZrHW9bGVsle2Z
eYDGtrxVHFbASPHzOLF94Xw6aaltFxPLEm6iU8XgT0XstF+Eq+mTxyhCEApn71jR
2nD+BVDz20iYDtQcMwZ5l2tjgg63QRlvZVMvsr4bYnEmHXHl9jdm68JntwELfCqH
mh6OthY0R1MbmidihuqvNlrTdMze5SHsgVs6S3yFbQzuBvs4pzv6MjfAxd9eUBQU
YTzeKtnGOYLE9PSSGLIknx191gcGdmVoWnsOuHk32hIviLUEFbCgXKvfPn9b/acF
Sn0y7TnE+hhOaJ72paG5IfxPEBtBO7Q6UAiL3rVAjx/4GJMHYtsxC41VrgjOFlhZ
RD5+Z9VWk8boPOm6LETEn4sDKzWecF/mlhwJdY4jjaJgnxrd5edGvcgLw4fiOcJF
yCCniPDEWs+k8eOfYeZ7ReR9uJc4sW6b3b6Iam7ckEqnzyPJx6jE5WhxZ9krXoay
qqS5V0TZ6/m+q7RyrF9zwFEWR/txzJrfa89A1bFtb6y8W7jH5EbqvfWyrDDoX+Vf
uPx1vPxX9xQ/QyvizV6WvLaB1+W9e1WS5aIqcdPEsSi6RwiOGO03gm1MAZGp9kE6
u2qQQeATlRLgrKqRthomoKP87WO8cP3Xzv79usDhxMvhGz66c4RQsjJcaWDrMTuU
1N/WnOUtjTXB5SFqF2qdtNVUqFu1f7ePLsw2DV9TaP+c0S5ojKlzVVyIh4ApmVrs
OfpGPHNJKFP2FLjtIYHdLhylQ/Z5YTKykaHvkSeRgF19y3McaW3nK7FBFd8aZbW+
7kHK6lNpY6BopvBhWM+aXhHGPSenbtexyMadwofSj4M1zyqopE8Q/NG/2l5ymb7r
xmvAfH1AJmial0XxNSlqQ7h4PSZfxlEGu8vE53qphuK+fjaQFXGnIM9OJBtNKohh
taQGIDI9UrCSl3i87rscvr/fl1OyRdLrZQ1TCuGAnqbd+E3rLM7p0sckGjdjukTT
I4YY8xaYEWXkajoyQW9aMe55UabinSKk6mEwSNdAEU1b/9FJvJtSJt2PNsgnevNu
HFwp7SiU2EYnWwzLHrPTD4dzbdaem3BNuKPq43J4+A3lTBOyo3CDQDPgBaOuGTV8
2M3kaCnMrw+N4k6koe6+UsOOQgb9inTCc6j6TC3WA7Kzip4x7vAGauW90p6jdAl+
Mx6ozKqPl1VfHojtVMR186s3e8eRsuMW6KKR6Q1U9isAJhju2sSsaUK+RohSvd/6
l683bgZyTR+VCWsjO+I11D0TXKNLPfUJ9iKAqMN69fHf1FE5LkM3cvX0EQQQTFv8
Kj7wjZMY52U/dV7Ofgj81EkQNLwvHNztpTSyRLnYJe8declUDjSAWWny6QtRsqfX
ckQp+2ORyC3HUWR/5Unj6ZTjH6OXdUer6RKojY7isPCi2WPFlP13jRbogm6aQ/A/
IoC2Z9DoZJzbCnOJmxNNXn69aZWAeLOFJgFGE17pSVOATroaK55ylXI3rbAi1HnD
QeajPa5wyj4Xeev1KEae8rdS+wc+QfYMwEod6Fd/vzqxVgDKO/uTasrX2Tqm4LPy
jwD2bh25JUftW6JTwPpHPwz2NOIbg7j7W7kqPCMeCTmrMh1NegU3XVKeBbbIS/2Q
DgBZXwfkvGJ2fQzt9wgWrvZqBJ2VMPbOd7q73HznWMeJ3lMvEOi5liTPihNmkr75
fPytjtcXWMRbPsqkhfDz0aQBzp/pEfWm6rUatjv2APwMj9Je+4KGCbDpWqMnJsd6
rm3nL7ruqCEo60rzZ73XNznLKXvSfgVuIiZ2jiGScBr8eQUYTyIBvPGkiQFSkJB5
x8qGtnFclGlccWowG8PYj3Y9TupyvjeMtemkm6MUaa4cXeZ6V/QwLt8TNUciI8bX
NUSJnquSIxWWygCmY0gjO76qLLMrPmJMzIldi+AdfEYuhYf3BlwnonWAxA/rHPOR
gYcBsxvpHBNxsdofj19UudFgzmIjdrtUl5Ou54JSoUg4TL5q1IedXyoP6ZopzTPE
uWSSAIEjAgjl/HPVisM01kWyt7tY4IVLcWxug9ITb6jfOA1L5mi5YWQdRTqoQVXa
SWhJzSiqql9kKqMhNaRlVYaxv8duQvZIRy6oSA/LNSdTti96V/E3RY/wQ5yA2nBl
cIrbxXaCZhBSdK63bpiXJRl8JRw+uglBfHkNXVAHSJ0Xx81JYNIvGvThv7jD1vqp
kVa6jBhNdMf0ooq0NGy49dLWHkCFySqbjw2mKounlMe0DQCGjOEJAIrLXGLJFbR0
Pe6PHxaXlczJ17bGee6ekDuRfa8TWshvW167q3CSE7/wemfxFivgO4MRLjOEUWaQ
IdgifkWTWqPtZ8oZrVBlQIDTI9U1B50rxEwbSSG3OUXPNb9rzrgx9ExP26hd8vNU
2DTH/aeyqFQvFFGHPMuf7iUu81VRLdh3XPIHxE9On0DIfQJNJrV+vUol15Gf65Ae
R1EYcMT6706+hd66SKAiOkNNMm3y3+VXvij3agQIPc3bX1J/BuILyxFK7WNZvbVj
mKKQPEyeyr+GjcgEyptNTyWYNTgEPT5hxH6NFLqC4Ku9tDlSGchEfbt5S/elGWJa
3i1/2yScISh3E5Y0AbDSqtMJPXvJdBBJ7nwyENfwzuZ1KJ47U1W5O+xokeuLvDdM
Ej+N/amYcR0ICHH1ZHOlNCNqGTso6JFIAZg0BukDw89eb24G+dw709UFUzmbZsEJ
HP2CFKsYJvtt/PgRccvCn/QI/hHSrN0ebiJjjB9xCIptKAQ8FjcFNEN4yEOaRwgu
YzyPRzfQrz3kNnk227FUFjgHZ9OYNWJ9L8l+E/wQ7WfGqW832mJupiFhQP/5FaBh
SOW2PJfaX/2+veS5lv0kratmhLWAak/bHIty2X4rJRyA7tI59u8dROfVoJed+3EE
Z2NQ2BaWk0xHLjmuk1pU/0pNuUTUFtGdzhzmZmdX3aOtMFV+dIUONaCHQuvCFjKW
9rZAa4IwhfmdAQ6rkY8vb6g3UbOBdmneT5d/NpsBr904OuCiDfi1esvKLGOaSZNx
+R4G8wLezvxP0J+cO5QjTOAlDMqlULr9+ANb3YJSCzC1xTrzZeMIUm5uNvhVFcoc
pOe5v/Me/deMC9gklKzmojLHzGtV7Q8yfIYEmHLAsgluB8UjW7iMu/2LLopKBkHz
HgXsRFOjIUZamPyWZCcylp/HJ1dOZR+XkdXIjM01vaPsbc1A9v5KuFBKFBaVC+9I
uLlInOQNP9ubYdLcuXo/yQ6x2p4y3x7ScsPEImyiXuYFLLUaVhlkPZkHrkr+asBg
6ytEDtUZspNByysHNzjVRYl3QwkXAQC8OGyZPprg6jwz8L+3xSWVZNlsLHZSYrnA
n7y9+YKfqb76xRfYH4U88M8xdatgwYFMGkuJKYkYU57baeHKevCJJxAwwbB6lUxk
hfoi3aY7XtS0FdMDkLkb1eOPXz3Xeqf6bexy+omhOQbj4fBTaxruchAqssxNM07j
AC4kD/I1qLBRA/9qHM7K7GSm7uryyt7Ann00dLUfnNOQm+3dqqStKdmpbyytqwuQ
e6BohCERQcPb4uueYFFwiFzCBTf0S4cFBmucs4P/qS2UNDY7RIuj6MaOlYba+W5M
dQjui16YTD9Bqb/eD0dwpZrnwz9Esex92ymbaVzq655GoxkqFqCiUjmR6NE6U+fN
ktXN9Ih7Wh+9HyTXGF6EnsIejgqHC8n+/wz10rU4DkeXm6hleC/Z/RsjlwlK+2kc
0AKeonDCUPWQMaQxW4gFz7Ydi+Bo0w7wzd98a4dDRrDSrcQksLDh5J6DSa12Izdw
r4kJnescDDB4hrVHpyaA2qkkhepNp5t6tAez/0PaMJfPhehjaFw78YVSmq+Ak1WO
Cw3Csf8n73jgOAgISp4W9wFJoT5i9mQaBZMpR5+6Sf6en34Y3afkgNItIV56UVgB
TCXD0ByoQ4i3EbQAdY/4Klk9xu8IwDaplvK2qz2dApyA6ugxdjpzYirQNVxYSsYR
l276dX71g4yYWcjehn/iwTRG+g/PanWAoQzft38GOn9e6jloTLQ3n29a3d3Pf5zW
+RLLSaaN4NMBPmcrE5bXaPOoIhDOL8x9AIxWIyzDGstR5I7MQflorq5WL/jbZh7s
NYCH1oRMosh4eJZL5BWFEWsVr2XQp5jkbmMRWSvFr/Lagrp9Wt+3lKtAJ+NJN452
qh0q6wyGLOoyCHZLkZbXI40ESIGzsPYMX3O5hiTLBE0Fsbj9tp6gs62rSjkM8MM/
EEUID4fXSm9bLn/SFZfgV7FYVOxZXUqpCfD5xP8J/Z+zdE+Euj2lK5pS/wn3I7Am
iAmhASH6YEsTaoj1lqLv493hFlUfHaHnJ/OAzwP0haTbfr4L+fjuuhorKgmkWX0B
50v2L3BJthwFlUPiQ0zrmOFIwF0ZOWtP3qFVE8Wjqb7wae0InOVzbg3IkTyMG96y
NKZ81EoEJeWfgYuSX87/OJPtZ3sGv0+EfAvZossNNX3oswF4BTBq51gD569UXdCm
enpxr90Q4nY43/+Zo5BnUCvOJg+wiADiOGRX2zXzyp0SJigEQQCOSNyWAkk5XkK0
A6u3o2Dg3z4Z89hVIhHOn5ef+cfCJZv1kHJ6G35TfSRq3DEPOb1Gz8lwnj7RSVBV
CwXk9RtJsnI93Yyyb3NWiHVYX148PpTOf/wtq8iAlZJvcUVilsIEG0rHg3n0ZqO1
+GW2ZDiImW6/Tw+Dy+EneypzKQMH9PDLcdpXZ4MV/LK3fa/zD2f4WkF4XXF8bquY
IoLw2s5vYuzwZVMOUlD6TvmNqLp3BTLq5EbuxquDE8CHnaNwPoEzl1oiG6kdbOOu
gUTFt+zM6QipNfyBSN3idMCY9aXnHE34oB1rNCFXmxHckYzB0So1TlKo7hWXsj39
x5cy1RAgFe0VDYvKtNdA4eBoHzzXh3kdhii560fZVXBbaUVSWrpAv2rYHaOiVsBx
iDd7Fy6QMFgIGlw0Hp75EZhHKsq7Q5eIR9TqdYyUb0IMEbK3+ZYQO5GOerVB79Wp
lvXaZ0SaRM+Rmen6fl63j3GBs+0nobOo1g7ZEv91vaPqBd1IuSXna0CXXeVSgqQd
2CUP2SirtWyF4IVFycmLeLDiDdR9/wvGDWZX6hLfExANpnbAW/7pWApkp9brkqV/
kKMQEsYEghlB1hnwLKVjenwM53eU7HDXKrAncGhy7om4xr3fHDyGJqSXIqjekpYQ
nRF8gh3n3Fwe3CAw6vd7+WXn2/mxj+EdvOodNwnj1ZgwJ37iSU3bCdiARFu//pKb
Rn3Tbmk1PXj6EFBJCRMMOruxyLiht3rGS+xh6PcBQEVvV4M1tNZEGbBBeEJdaCug
5R7LHI6NQuKEIGJ2mgJpt5CjGj0ERzdTGjm5iJ4+r80K6gokqrwRFYVmRdb7XobG
pe28XU3/VQroVDNciUPFi/bZKO6GLpCg+N1HcBcPkMxZJ0NyQSkLFtvIt/uWP/Ad
z0EtXuZZiYGqpkz7QBtSi6Qzn5iW+9tNyxHk/bqevzS3oo4fZeYP1vaxiImHMEev
bHkGlRkCcvleeRH7oQZox8vrkCENuYSKxx7Zn76Ew0oQapAu7LjGfYg2+InrFQvI
Qdoa0wTg9+756n5TaBUhrEUcgbBMZJzwrzB0v4hl3uWGV56SS2ienNqz39jMAs0G
W5TyNWXf9nRvkR2moFtEbB2WJ8HKFFhZVLV5vKVzgL2P0BR1ekOHQOueg2Lo/BN2
mjPX5WbNTZh5nrc3tnZcXlozTne1H2nRosj30qarMvLo163pIVyI69PRfPf0bVF3
AmojmtYdO6DFKFieJm+vR56IqdpzUmdKuo62uHsCY9dxheXgkkj3ZNH7HloSTbX+
k711xk98GnLIvn0/SLGzxekP52WbiQbr0AK7nCVyP2yLQQE//ewQkFxHHj0cGrqZ
0o2ftoULY2Wg+0/bBoQJc4oyYywROAxos37H9br1XlFYHLUJRKr6iO2yzl9sDESI
xrKSwZWsONZyYsdFrV/e4Xi8gcVrPcJffvIP73DxXhib1GbCZ4GtcIhTHUt/iwjN
aSemBk754sHjpDuRjSxwwP33ozNhDYTTaaWZrfOwkKBY1SXeMgbPULRnpJzsKG0j
wtnuJQ30GAOndhNn2kyPBlSsj+Vb8kXhTP2VHeoYBHdC0tJJM5n54AA8i3u25/W/
ZsxZUv81v2+rOskTaVXDHF7hXfpRurqETc9ThYXuLzMdPpmF6ck1vy4r61WJzJ1+
HIHNkFkbVOxd5PXTpxkKgZaoz5ehiQ0NlYSmSKM7dvmXx7zt1ZR92CoeoMHid49u
7lqjR+Gt3zd+UZCjglBDTQ9MlzTCDDKRhlmFN6pHt5/kqcZuIOrF90bQUSe+qj93
RGDWs0YavrCCue66WI9ZYLi/6+WEAixto6hJ9k4gAw4whfhauzJFtHokSeyRNnKc
0KWwBAQkPeg1ygWFtxWAiapPZjw7O+19FF5evU4+sFSEcH2E/brW+bYky01L81go
8tKAYFwYsAOYqIuhF8QPTJF3lSy7tsUnqvdLpJDTkJ/70d99IJ1Xq4dnyKsfR9SA
KOs9qxsxrL6F/yp1rHc9p2bQQ6sSlHmralu7VpmvYSsF3ed4ijLf2zAcl+15eYP6
Q9kuRPAHE2ThyYf46govMmQbqWtBnAYJauSAAFzFQikLTdz6pfSUFYdz8cWmfykD
+XYSjtIZgYn1nHBdiOyCcH4al0JmfU+orPWeaan61U8O7wMnS6U/YOtNj8170MwF
88+ZVKZ9orovsUtrYW5KjXfJOVCoaNJim07sB5XwDSgndL6nISt3esuIqvnvDPd5
6T4WbUpyAhygfWH74hlGtN7iUWWLW6fgIPxX7k+u68SYxi7dFVrPleGrzq+tgjDf
eLih2DyVaMxa1ZtTfTzegiArbE818fg99uEoN1II9yWQ/dHmE4Wa209IHymemw8+
ueX0VZ2NFH37bLiUBZL+fAdmpcI8JNsE72nPYvGoVIQwNLDjqpNbhz6olwrV16ow
YIR+sHhxCvQoHOETEBGFixC4Cz0cSCPHl4xFSOXyTjr5EaiCgqfEJWLS0DqlcA9J
ZDhcuxgyuDeb18gX9bEzg8ENX5fTEjVCscK5z//pLxt7Cend+vk1W+/tjktMThNT
zSqAfK7Mg5MimhFuv9v285on51KdioEyyg39UHi8Ozreia6UwkmKvG2xIBYZS5xy
P3Uv5vnrksz8fGNy7YWKrP7gG59nDe39qz8ZqNrFHQhbszQT8+SVDmV/yDcvzqlP
3awoB6M++4CN9kYFNe4PmLzXULMjS6qdbU9TDofTmBtMzFRJVvpv26psthG+5oSn
85KN3SSNyn32JC2dRs8Bvls4dDk+2Ow/1f5nmvBPGJLWzUuqkpfwWqpZurKvuuEJ
bscliVV1tZojERM+4JlxEFwKx3kI7P7+GK6ZqGz2KAnw+vYETRT1pwAJU56EChFW
wookk6v+xXRbppyO6whCPQ2dunNyl0nHwCo07x/LDa5sgBsQW6KtCsCDr8dZNDe8
MxPVe/JsJRbgfhkBTWobaNHdZ84/DeZjd+ghIRbA3IBScR52DwXu9J+Cu7oKmdS+
35AMr7rC0qzSVck0jNWfaLvyR46m63vikaB3Bjl5US/KB+UEgO06XhrDhSm6GTxn
W8Jw62NmuFHBSWSPegtpaY5glfFOSvIt9W6eFVDNjGv58yAmw/sCjmePXwfQtsqp
gJCMVSmlGhTd9GcArp3Wg9oeF+J/zVpblGrrOiy2N3UwdnjrUExpbTRpSTvhqRwI
YhhSvrzAWjMQIyigbx0aKEZV6WcjQMiUq0EFPtqtqIwgrLCNs1YHbrmt7juBUqkI
q5XkbYyIBjnyJLBE64Yhr/GdrNyPq1eb/R4UzcIhRakGbz4rrsP0EyUzOFhkeLen
Ndb0nMF5eoajhpb4020/vJbQEsCWPtvvBjisM+sNEB6/UyZOGI1vOGnPipZWupPZ
GksXbwVJDjpYHbCzO0qFP5ydVZee930eQ70gHRoxt+862815AXbfokYM7C6CZU8s
lYVpbo2xYbc7mVIR10RPm9mS5awcxQa20IxWfYU3ZLBCrz83ZnLDsZrUtEfTj+6u
H9MMg+MS/zElvhRP0WtGttnBo1ISmDtc8URkKV/NHWMK1eVtdRq82U0IQKve5KA9
qg0xqZ75R4PJ3crT38qaE4KXNFeScukgWnav7dkiKYNgwByqJb0pzVAwQCY0HvU7
+DWzKyqdME26a9TyF8BSKK6369tcQckCW0OeAjZKRpq25Cwlrb412dABBTQBG2f8
ark8Ly/ztJdFLacSdezwKO5976nHUyfIvOSh19ZIiMCXh++DNo6L/0AU4hu7BbZk
tMtvwa5RMAXYPyKz4yd3CR1rsk2fPf4+3BkqyRNcHLkE9jsS4IvGGFWYYZvVIdEE
3Op5zXyfxbKbH4AP8FC181zzH88/M9LZ1j1JmNOZjt6y3GCrgOgDFnMIm8iZlDPe
pdnAqZn3n2MqjBpIDwqJ9csD+8W3TBk4G3FyS+5nSrZp3suopnaV/LT2hOF2nRFm
0bl9KTt7gL9h/FUsja2yWNkvijqvtkm2GZWDFgTtNh+h8oZ9BW4abGuBnSehA6Al
bcv47KBKwXD50WkBpJsRyu878tiTjqouQSCxToiaQxtup01QE/widfjoZaPWXgh5
p3dsLOdmgMmJWs2RpZVdQuyJAsi1P+ab5xpiO83w4tG0R81Hu4eAu/ep5BaoJ6dJ
V30XfRyku/IrcyIdMCJaQBhNd/bv7i0SjBftLYnR44x9gX9N4wlDJV7Mi25xLum5
nBMhRavdoVL81Rl4+rguxzIULTNozQKhrv9mDAj6+5WPlrjjnP8sMjkAgDyCBCEp
ABZ3bUMPRmsSFx3e1cn6wg0+l/siG3ITEOPl+qK1J89Dq2gg1UhdD+khUvdtlrhy
NpKTugwGpvTwoCfsoQYUjP7tWpO9B+WuDxsVTCPw7KYEgCX+9Ya0yrWK1dgYjua+
ajhiOQtHQVzBD9CPfWJEl4xc2j+JiaV2k9lFxnR441HNkqvRW5n1Itng+iOcJSgK
EOZbp0my7MOfua3ftZgAmh/D0t7dDNLSr9yen00YgD2GZFyTSti2ZOQ2R+hjjfKB
VTzoKCi/n9ddYb5mZYFyuYdIiHTQ02WNnWKBsS3TVZpBCk8vduUi81BP9ggVN6s9
bNTnePLki2HvEyVTziubNQSx8Yk09f8Fu2sdz+I5tOhTs2eBOguQUvq699qifXVL
Rq9cUu56/0BOMnlePOwzrC4sK1Ek2CIAZKH+7lEL05uzoSUBiVVO1gy+GakPJEub
NwoP8KpH/Ct+iXto0ulwjyBV3A7n2ddw4mG6muYsmqudwfVgvYATz4mqQj+7FO6R
j+aNlOr0bPuk9/YiwG+DZN14vKkhOU0Mse8iTpSjTU433GDaw/XgrJK7PD8zprVc
RXPHrejGfKCJ4VBbHMG3cTJvY6G9VD9Sh8Mx6T2Krr7FnJEBhd7N8e7ag0MDs5NP
hYgfJD8iCbO6rMRLudCEPK+tDHP21Skdrbn8Fvbq8AgWMasndALua8PHLR1DvHg2
Obhtw5rYb/XfnnBJQv06XzT7/Zze7icuKa2knzQrGyPr18rDIyk5THpiZYC6nEbd
ku1EM4/KTsEKFqrOYKn9Cf5bKQeX7jabrWHZTs6FSYdjB1ahvAo9/rmAM2ZMbIvU
sR85usq6pQsH3JtYRlMw5Lmeo+n4n7Fka0di0UuyPWu9AaCu0BXF3nqAYaQbTN9z
mRKwtHGdUFIssspHbHtHthv/jbTFgGx/f0UjbPkX4NX6xTuLyQLCJgcaHLra4PoQ
34RUme+cbZEPrAGqIkzrh+36Npxt3OY+yOXS+PD2hJGgiKADBwqhYNMWPfC7Apqn
Oq3N4EiVae0qIcpNHK9fp+/gqLIDFlkBE4zTPg7w4ybUfJ6Rw3imxcn/GYXz25Pc
RFKQnvwI8/kTiD5s1/zKv5443FnOCtESAL3gJM2y06y5xzIp+ncDODlKK4AV7bQy
OkMQOgmsP+8cXABjlniLIbnNu2kobNDkoZmx41oze2UaM9bgDywohc6kURxXaV9U
4UvCpmnNqpzFnA0EuDzYpo5o7S1dZeFx8ua7rDypEHdqHt2waJNsWtgJaq5tLDBb
h7ID5Sp0/yoUziO5L7lE6etcqWEtp8ZDTqaAhk44JvWOb8abFX8XaJt473wgl3hA
eKvfm9yZwhEibKxCxFIKFayVt17UNOHj2clP86EqGGngF7zG83J5NVprTjBKPORi
2Ju57MmvstkpovG+nzKiV0WxAxhU8dJAes2j8U2mTPNFPPuNsTDgr+n4b4KudZ8M
OR85K6SlkSz2e5UBvcKrycLcquFaTH1qb5kjH/UtyqWx+IZAXc9GbCQQGvcyZfYO
Yc7oU+v7y/3wtlV6tnhPvEd/OoQlBHfJdAoKYdZ8WtPjRaUQHMCtaMJIdGu8a50L
jX8StMFIWE+Hrqw1hsZoj0xWNBwjz9pLwp/h0HyXDjRLTCnnmoUTx0XEwQFOINNV
0V9UpyhcYBlp0T/Ve2v50hwU1mi6yEK0E5HSEw4M5jdRm2FwudhTuLemWInKIqJl
PMoJyItSpcOX2PkUCYyeVriyhF+GmoVS2uvELO8ldd1XIosJLNID7A2KRG5OlmQq
0xc3BR/NyJ0c0rMQ9HmVkxKZeGmWorxV0pCgkNtnId7Lp0+3MGPD6tD/CcNulcBP
YG6isu4d5w/bLO599DOEaupYw1ZWNcOLhevmmDZznJzD/yqcGD0v1gOl75lF6pAt
yoV15AptRzcfpMI1F74+BNAlHR8ag8Z5+2W7dz/2Q/1tFDzmgRwMYVIGcUsIDQXg
H7atktKi0MNBjRUXZ7zOS4tC6c27uc5eYsL9Cuv+VhMiTAmsg0skk0qAWTItV7lQ
NcIV4SDmGDbhUs0hk1TztVEyS9/PPnv60/l3Udb/B7lDlJgfVj2u8iy4A6Vv/UIe
E/cNelhNsOTs5VlWKLQKn+8PqaNCBhzKYquvcNPUuxpGbz+lfXskIcDwyYcYxtCP
6zAl8HWAxdGjJ13ML2LsOUr5dzKH36Jfh0DKeKBQL2nSfFA/qT/udcUiNTu6GOrr
OMtw2mS1aSvFdFjbiTG7y8XLiFecMkFibnkwvA9TuJQ7j4Px7ntQsBgzp1WRwGEl
qtV8RyHn0yS5V7W9ll8oBvS3i21ka2QCKMu/m7W+MJ3009mbsspzSr0SjI79WbyL
2h4tAJ6c3LfublSpGjcj/acRHLse/RhUqDt/iwjNiBD7Ido52MSbup2i6poWikg8
snuH4CnP1TRWvPVT4+BPSrUNNYD49OY9pgkM4ugJcBRMZ5Wk9GIoLPQUItiXCWjh
idoSE9H5ewTjPP4dAyyeXzLBV6xEaoukQIkYaKyNKa3wOa3DLu/wJaoyvtpe/RJ3
BgTjUSAsNIezK+9Rw+AETfDBYrpJ80bgy3d4L1tcI+3pRYHDbfESyXzN47BZE24y
x6AHDDwjMHgARBe3yqUU6m2u1DLYk4e87ceLkEqjmWW+HTj+8+t5Oe7PQRo+KY+8
LYLULdryyrY9KfOJVtFMT1oEikmyEanT+cBf8yDaAXqGqa7/9ZTTVn/Xl4C/R0bV
04ZmY5JvBcvANhHyUL8mWs6DsKxMsXlsF47/t1U5cQ1r74lSdnKDaTVHBj8zM0Y1
jWcMzgab73PKesrD231xFELflrf5uHQ2HKQqI6EvR96rX0FlK4CpJACA/Vu3AHET
NZtcs3JZUb+o3ogGDTo8CYUcjdT3hqL6Fr30GhlZuoVaP/D5sSggiBodNm+1exp0
nNyro2tDQQJE/OpB+I6iY5j2gTo0pmHOhx+jB9zxgYCWd3DEGG71hdzBA8KdcOtT
HatykPdkHgUA1wBuPeeLMEf6Ygvr/QELuHUfwpeI0R0HH3Ri+a4CNHyG34igdgtu
cThx7LABIKL+cU41SkXqLHyS6JNsp2weQhJ1HH39VwGNWVytUk57SFTXzR0QGukv
jeoAVZYa//pY6gh40ucnpAO4QgNYiX/VKbPtjSjse+5DlFY4ogt7YK00T2+wW9Sc
4Nb9khWTlYb+91xfILh0UzYQU40rFgP8535SOUhWBDuOBiXkLTYfNHVwdZNBfdNR
RpE+I8Y5ixN1LmECQn3foy53WVq0nf38L/O+vEFT7gdUrRfnPUTu1Yq1mkjHFzWW
JGaTfHbCW4SXOJZfsL56Hu0hUV2gOuNVYmEqDn32SrUJ814NNzFS9J2V4WkWsA0W
qbU+2+4UVHEC9pwkUvzqjFMxNki4cbt0VtjhonmU3QQHNS0ZFftLId9e44Qf3lo3
safk3gpnKTNgHnCrJHGC/KCqPmZBGb2cnUYbltrAybLX/Cw5HkQFajq4BGNpXbWW
8i9OCdfCj3iw0vskrzmBsne9UJnnBH1y3KQSPPaatAiP8Vo9i2WenC3RFRK26D8u
gwByQcp8wNpA0CMFM0eix27OYPNxNTWUHDhMjxVDNGBboaudgEgP8O9I4MZfh9LJ
uKKsU29GmAoBgeh7yQOgTGXNTwfe4hXTyOrRsV0n1fx2Agbih7RUB/Z2W8tBz7Aw
vJtugurBzEz9+R178bLpBG1YohYGrKD4xINcUtAWitk0xRJlNKx5XELE2xeWvFl+
08N8oTcL6rV+QwZzHMgmhf76Ux9+vNGFqtrVvsmrXeuMZo1YoaxHV24Qxvqui72Y
tBm8rBsYdeccB8fsQDYFdA31eTVW165ez87BWyLqL5ZowZqkaDpP/wT15wRyQLxO
+Ts5vkuGZsMHDJtwWBnJOwaBRsiVTHbLZoOPXrrhbdymueLk2HRVDwYzFXnaCBHI
InhnR2ow4u2/Z4UTP7MUgaXHqEVBYFKce2L5IbizTxvy4UKVzIrPlCAZvy/bHixQ
A+I2kFCetooRPH6DcGairwnimGTupEJUbZeLMnrcCKr3eKojsRMHjUnqmaSCv4RQ
6AWaG4crirzN6VG7rW44iHPpFK8vK6tsTUKVzRGhmJEp9M3u6rin5S2SQh+rpquD
4Xz8s4av1H6jXcKOmbvgWceOIWTLXOer5vjLLMIVX4Ypdi08h58+ByhCXfQhLVy7
vZGsPiQkJ5wWdobs3lHLiR+KRM06C8FiDbz3d7ONE2iDNB+b+TxSnCosPjZxZ/Px
f0+nAO5HLL0vV8ey1Bj0Otgf8lCigrNradkbMtAnmI7ixzYGPEvmUQ5qfnb6S0EM
LQHDnx3ie4Z+c5EJBtMA9Ju4vh9fUXSUIUGgJojXsgF1Qoc0nXw5OVyQpnMY575t
LZBjrBcXuk1u0iI27Jvt39juLyPbSel4i7VJ0mZGtPCbRvJ3fMCjLbdLLKEA5YMi
S7sird4ot5YWxvcZ/+sqiNdkc+qIFRbAdmU2AmyFhPq77lGJeEY4YrVJGX1OFPe+
pkTP+w64g5lmn2fmEDe56yhEP7vM3g50vm8fpMcESwUZJ13lLPe52WF6562mNdpZ
q71NyClmsZgzBbSLaPCZ5nwHE7N6iDPB1+i16b1Wxg1IY0/ONTgx2XCQJ5Jybqfe
EhAfNq5nvCXM3EDj8mI6TTCVwu74svlov9dVEIRMhrwRgezeby8eKsMuH2bz/1u/
F1u/Km+UbHaGxw4DhODAWLjNdPCw1xEgKUeQXoOTPR5M4P8btbls56Imvgy2FpOa
6n44A1IElDrALwI9rtgHl/ECaDKvmmwfIZ/CFPMrlYrKYZGWPR/ixwSGHH8fpg/Q
R2OYfWQPJn+CnUihvnIePhJ1zDgjmAMFaifiNnfYbTQYoe/mfE2KBpvrbQHjgbKT
BKSnYaKG0BXxbfqYZS0IHFG7JDOzobiwvm+JZrqonxwtBGTBIVCVQ6PKr4qcurJa
f7WJ4iLnhj0EeGsBpZuhcmUN0m4OrtkK60WFMKSEj+FBY80h7IVE8u9MVudTboVI
oUbnDCC0pA2jwf691mvouHqV04J+vnqM9zRtYNG9PJmsi+KJNeAx4Xvk2nd9ntH9
h3uajiufcYyJGflkkROU4Cgm25BeJKhQP8DH9HKDWulP8RPkR6hJN/AO6pEnLxd+
NVuGuz/KUnb6ABLQgNfQwzkXHPlpbmI9Oc+W72BEZCQ7TU1wmRiT/gYOrgRGfOp3
6YWGc9DPrA27wzzUk5NDhjLaJcArqWXOkHtWiTb3Bi3jEhQk5T0eYf7cqsZMCcif
8YdCdGz5AErhHsVKRndjD8yp9PyQcVAN1Ch2s2qLg32YTc/xBY+LweZatRe7sqOt
NhaASLKJH9xVY76LFAml9wWJVS1gxQjToIicdm+3jQT2AL7VHBVKx5TCHL6PlymP
/9g6BRG//cdQlrqUWtTFIOh4Pu55yz6JOuxGi++7UIurn6goRc+bgTzsnYtSxTj7
SjTpSJ88mLG7O83J27/kObsh64WqKf2MwL+PlFiGozYS5kCV94Sodsry/5ZEdweP
XqbPzwWmDfVXrUvPPh04PVwBlvHJcOEiKtH/khYIrLcBCBJGk5hnQPObXgTUL5s0
z+mMPzpJef7ioJjYO7L6T4jYh9qBrJg5RlnGzPi4F6xPFZcf2Kqh9QA4JByVWwHC
6G9Nl0tcuv8uPtfDvCr9a5jhuNS+8U6R6HMsNu1IVjk6lgLmHXVUuBJfRF8yxkKj
gM4XhpNnZNUlbz38AOoJFePMRaPhWAzAdEnV6MuwfrXVq+D+a8B5LNn4JVVMrN9a
y4wcQzBcC4NbMPKCbn9KUpRWOq1YZHmGnfJG5iaBL4uXJgjREB/diruoE/Mdy7Eq
9G11fruLlgDU9jTmtJ5XjhYVYE4sn/ws95iaqPgSkbmQQb+5Qesn1viROaGErdbj
BXlHn0Qkr0ghFs2IMgLi2lZbnS+gmtL3FsiD6CMQ0Uin13QH0OeGvYxRg36Iaimi
vRWTdF7OvURM7Uraan64ojzbxqWE/9t0HE16xGpf0uLJMo3rqW/vY/4t3qNwmznm
/e/dwdJkYbbcWkaX8bCjcGAdjvNYehZnErR117/lpn+2l94YSsHut4jzYWF17Ffh
7DueexA5gVFlI/PUQxYOqOymP0J63qtFsKqs/gWSqC10r4UAsqCJ79fwqzREbPai
gGR4bnXSBkOIbFFBeghaTrcECsPeDOeIlmmeOjaEEi0oQt3Zmh7BiAx9opZK51zz
oAt2SwqD1/vOvKXp43oqj0CGDYiGpqhi2ohgruMoWoX7qCn1O0WaCBObtjstdYeE
tQl0IAu0JiWi/itlCeZppB+hj75eFSx9GxfcWIQ5ETs8ssHPVjD9+HxjcW2lvUcA
XrQ0WYMiaXnApipLqp/Hj9vVBsvKkq+yABlYvZctPbERl94ux61TjaxfPR0LwMaL
0afiwcu3woS2OlHr8B4+uVYu79ZSsTU03bHGnbg1k7oBBnzpId4rUG5UvVLz6gRm
N1m4rCfbJEU1faydHz0GAIvbzYBxY2BAzzla+MWXBaenQizHHDJXweaXa5Zomf4h
57OZ5H4gTWDEdJTnxx7fE8q5+8k/B94W19vHF2OZrTFW2DKnmb0oA/hP2+xbW0QP
+z5e6oWt1pavjywF5oFR7bHVxPtZNm3cSXP9926muY1AQyEAi8xsibOTV3AlmZWS
KpCLy8mdt421ePEMtE5mejodZzYi/31n/ojK3VrKbMewx7+VyEHMPSwzvrEXtJQ0
LFr27KcyNXs6aPYWJ6wOEDpD3fXDor6cKHKwMcZF6t66fNppSs3P81/Tae+gQ2ZE
tjsB+NKubs7PwgmW/ibgLqD/W1YYoBOfyfndqG3juTOXYKHXQ3jZIrgSw0GVaXxg
N3U1+/UFf2pfV0vmOyJM3Qo2WDQo2VQm5ZxzJUymQ+mGT+iVmqWN++edQyXqZlFX
MARMB/Hev0EVatocrb33koCTUNRLaiuwkTsouogSLZaE+pczCHLuGxZwdrXFTN3m
1b/ul7GQQrTgR3IY1cHxC8G6zosP44DLH/wGdAICCDu92eKuvXzMmybF7DMLiE4J
1dEpCLRrw8r9KkIEamsBAYytTtD2+7XztBqe0bxlcATBPVZPDL8ra2lQ0DdSHROY
iA0H4a+5tq6mlSG2TsxVSm2OHq0gpuwIyLB7ylZFVv6pC9h1p2mpBWv+T25bHYPl
ATHyVjdaExXpwKG6qyWVHUp+V/Lix6XdMivj7/2F4EICrJaQ+Ae2ZK0gySGZb+0P
pPSoUZPn55PGfCspx8vKnBzFcXaa2bEjUAXkWdDQmdFTlC+hefBaYvnbx0lEO9CD
1jpOfwRLBMoMe3+9n/wtt5Waer7JS7Pb3dAQWUQ4rCUhQcFRlrxLs9b1yfFPNACU
E17b6r+e3Y2kD408HypnsYnQ+HuflfBXQ4MnX7vrVsTCGgOICPT3y/d652oAntx1
KWJm8nJe/Kc/1gzi7zD04/UgxI4WdeNtlyVFR1CUvT3nHE9cmiURDfUisHjY8Zlw
sNC0LEId9GPrzlGPjmqut9UOKGNLvq1b70/RkRTxEhcET0wgd0rOWlU1Jjlc0/E7
`pragma protect end_protected
