// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CO2WsXWMMYVQIZGtDdD8txRVwhGfz/R8U9as60WcmGamEIG2fiCxbH+UJcu4MRry
wtP1/0zYrSdVkBujaeaU199LgyTf66WViyEWZFVrUfjHQhWxMCPoFvmQAWvdw2PP
/izkbwEoHHsipww+jjdT+kMPFzKa1zMOxYY/6UDsXGI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1408)
GYKnBSZAXfThzMZ+0uHbzM+hK06SxesSsENq/TFpJN5Mm22o5q60+5pVh8MwwZIK
ipD+CinQP9+xQstweSiFdNBaZORYmohkCk0vZgz3G6bGNR4uVuFNp8mmy99tRNaZ
UYiOUGz6yN2jXQyKxUa7/3qmDR9CrKLQZXxkemlniZR0JSC7zfqG5L4e6nTrUFw9
PHZ+1nVH5aWxSooIbWBI46TipwRSn+8sKBEQ4Ws0CMfRM4Fch88UyVfRH/Ntzqxa
Yg/mitIfU+C2HfiBsDmGG+b/sRoR5QZo03DdQIHAV9XtspWDRYA6tK6pBSKPsc1D
Jv0p7ys021coUntQwYKErzoGdDvNZ/DXf4WV8sk739/Kh2tkQ92EwzQ7I+yNeutF
mB2whRG+hIhrfJM1w2LlppQzxGHW0hfff2J1falQZarP2dTY4I6SvMtYZh23plAq
Vfx0i1KaV79e09qGtlyAz3MNSyhD879rPvjQtuSCq0mqeSKfE3dd07fmJRQXXeiw
vKLiEX8mnvYNEvCB2L/eYhS0vPifSiQnlSYD1xqFk0STB0MahTHdTGMAxcoN0j1L
ekyjP2jHiiNuYI+8W86Cak00SsA1CH+cnsMEye29YBXaWuWITimqHLbuD1OSczpv
obuTdQ7WBdVD4FpRpU8GiMfA9NqbktKtSxQMpJGH5UVAkyiDngpyVbt1MfP36ai4
j9YzG/3wLcYD4s9K0ppYHrwdSe7c9PU0YVtTwt69yrtY52NGdtom6awAKgpGwXa0
qNrP213fmKjKmcEgygXkcik2JITeKCGEk4eEtQ5/Q6r2itW0oTTSz4dqeqE6jlK0
fodviDPham2zFHvfCYXZYR/1BNL2TpG219oX5pHV1Po30v4PBJ9zrfkUqx0oUurA
Z1xUceoZqZPIRf25uvpP0mJwESRYbbyeG+wkf73Rk3lhycnE2e8baZGmltoGw/eS
3yJEvzWxsCL5XzqjUS7wJu7wsFl1c3I5NqbF2xAMzi0ml/vc5WtP5sTIF8liMePC
9f6VvLJJKhG6jZdezBuF77PhZNdu7j3IrPl6L1LEuO/CLFNTa75vDr1HQnLLqKny
l9bfjZLJPIA4zFFfLJNZWVxGLxW0QwhlvZNYSRoMz0v/KBXd5DeJ3cbjPT2gSOI+
l3CuvqTCg1BeNmjF3w2iyZY4N7yVn6JzQDPbfj/35sX5UQQFH0LLbd5pxiDTHX4c
gOhQyOjmB7ux22PALwObw6WMM30G2DU7Yi8cPMzgxZ5Ebx+i6jkuN0z973qQBb5n
StZbiY7ph2+C3sRDGOUfACdB4vigndv871GaWgN7R7GDcp9wR1haDSeyQrfmMSl9
wOVo6DPlVOmsEtRVNx4gBkTOOyJMzGSOVZPBjV9PZdznwmzfdxRci/BjSAiyo+ey
hWx6Mbh08UpneO+NrvWHtnaXVQBub8/TNqa6/uIhzrfVplvdRfiUR/iXtQSFQkWU
m9Vb0aHMEps+k9HmRekOf7GfIdLZk4xPIG9LpAzjlHgF2Xp/8y8VWX7SrtjOy3l5
Jjv1bqMH++3GZqeIqUbrSVhWsotDlQqwggQurYF/0Sy8yPPkK1Jnzi/G8FUkPF5j
nLHr/+gyfV54FEvwOl31hnar/kbmGImy9C3Huxde7os7iM0sD/ZXTcTGstfC6rYm
h8K7TIjU+7BUunsN4Qm0jWBFdPwNa4B5qqU1nptLo2xe0pnKBQFuZ0YBNQk+ik3N
42NreS/W0m3zscOVc/GArDI0mpjgJQQ+6ovRLi/u48BfjjFHxvDrruexyjDoozwl
J9LgUev6X6lpkNnnCYnhs/+iPjtCUT8k6hN9G8/owhmUhdxdHWSYuyc+uqsvlw6F
V72z8ILm9bC46kT/2jRW+w==
`pragma protect end_protected
