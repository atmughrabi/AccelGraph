// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oMbrk3eHLJ8xFmVRTyESvdI7L4zMmxtIn6qGWdyl4FNlA5JeHJnz/CBYsCKYalRH
C5gVu4vswZG/TSIbIiqESH55M8Lkwdfg4IX4tNkVvPxIvQ738cZyUOrBotcgKvsJ
9VptSc5NvSr0RhVLOfU7fkTz+lo/uMyZr2Hj0KgF66E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 45680)
qhkvUrAzYnnzhClA1aQvmcO26vZRQ37Kw6tMCbGFo4wMkZbp1MQuLKxLZ6roEIkZ
zuOetfG6EmP4f8M4ZJ7FetSfGTjloHWBEbcoMevELyoY3E8UUd0l5fY3WnEXhgom
5Zs6ZOVvXrwildcVahzmVDmRWTh5F0N3f4Lsl3Ij4LXG/aOvUrKrEc0du2m5nwlA
LA5Us/gR5p20XTryVS04UcOmztsGNrX04S8OGCQJhGRrqcdfKKvWzO8LCLko9K8N
hkMN5oMWFCIoR4d+grDkW65bQ7EiYNUOGmSzkEZgaaoOlBk9VGT3Tge8OvwX7rae
yaaY800zBNu08cDf0IhquWbCtPVjLaV2UT0sK6oS22BLBULyOhWVvsedDkw9I9O3
4J+QwgGVxUHZNHKefGYE1f5SMkgKUwgVBeFR4dAX/sA12QVQ4smotkZUyFyp7bX5
6ThEIxCvmPOr4P1PqudlXvOU2+Sm47+edSC9ifUQpZ9zLtI+h4IsiIpIHodXbQ9w
wdI7MiYF7dbGelwIa9nmkCvjp1OImLioBBJdvo9n34oX3IwzoXDu0Cpqj+MZWjyq
6zahjc5Hm/LQ4LNFXrX9zGj0fh9kixxVw+dTs93DhjUgaqKEzy7rjPVmBa1c6Nfn
5jnMh+flm/S02VV3soxvSQ9ZGqGGRvSzT69QxlObdV54Xbxy59dlUS8GDC4hEQb6
IwVshLQtOMgiLqSaOC+8hgVT8gQiJlhaOpgO+Y9+0NUdq15FKg33jaqrMYypMSFJ
J1L6o/1IZQu6VqHTUhfsnUQNHPyR9b+K3+40EBVQMkIt4z19iUDyutX0dmqkOWP+
uzI+Q6Lq10kXGwRoZu+UMIzirVr2r8fhsBxVBpG+hOvMkZH39WU7VL5xcxo+E3EJ
I+geh6MCFN3oiZ9w3v+UuJPWRIyK5gkdUx7Q/0IE4GNKA/kY43q2EyAazL2OsQHL
O/7E1kNFVCv+VwaA/a8tUcZyyjS8x7SInC9nnSOmcjhs2IlfFJQhT5MhyN4demtH
OtoKDiKn5I7w7Kpfk8uP08gyNEQ3fsKP1dnossWjVrWJDlRu+1QloVAb1HUU7tO/
LqjAmUSvhBiR8MYlamnL5Ws/r1gpFqhc6WoonpGYynVvq5uTIFr0a3ZfCCzbnpkJ
Dg1zN6t8iyOqM5XcFk+tEB7wowbooFh7gOYOLjVSdFrS8Fj6eB6IHqUWu1iRBbRZ
5PUQSC4x9lqtvFk1d0//VaWD8EblNCufSs50a3WM9Lhj6IlGw8Jx3V0H+hj1K9OB
yAQTxsxHEqESPocMl7Gb5TA67COtIq7J/aaALm32P34i2+l6G7XZ1+8LlddI1Myk
WqSnCO6T70EeduDwePjs58DEbCs3L8M7rMxIFDaB+yFxPnH06pw0fcV9IOfxA0HI
OdVCXksSC69FsjKBT/IaBu7rJ7V3ZUexVDbnHE7JYVPyKzMwscipGvRwTmzaIwRY
v1KRG95FlBnk+X09wJOwof7ndZTd2zmJcGbHUIyzSujAtvtp6lI0it/6szzGgn7e
reXYNI9BdhKrdCjto1ouK1UzgcpCzlTxgv+WaSXRCdcGBtmGjVnIJkv2oK0taY1X
nm+cC8F8l2SMU+p7NW69brxWj9nsR1B+/O0yPMzryjJL9MNQ2EiSYRxwwYJ1Fb9v
i82JFFvHtJCmO0WRyUp3/OzRpbYih6+eXIZBHuBFSBcr7t0O2SIoC6VEgF8Trexr
lEd6DDLVW8HB0sE6aROYwpQorwLI2p5Dpit7iFzg5D8ARQJ4txMlTnVP+870ezzS
agYa3B6fvcTR3vMomGM5aFQQjDYCnVmOgzAYy2Vw96+4jnrbMF+4A8F1lKkD9Wz8
P5PNezncIGoWsnVJz5JGXeWn5O+fdS78zCxj/4SrQdS8B9Ff/y9OGwzAJD2VQuF1
/Qo8fWAATVwY3hLPo4tvo1FcLMgfFX4VmqdINF3tuhLAkOkahJMVa3YSGJgeGrcf
Y3dkjjGTlwOa8X1fD4PVHrr524rioOXkEkdCA8ccr3WKZT+kkl19OpLVp01Mkcob
wCczvfKCF5GvE9ajQm0r0oGglF29GN9fYcV9dPASr9dzqhjQkKCyQyOKkyb+JbSi
2DWajvWub6SYRkcsA4XjpHemyfhnu6AyvOIuKK5scZMBzUrNCDzOcrVvz2oVbvyU
jGELNBcQvsYlJq5oJJy9rA4pX1gLVxR0Sb3O2xAxWauWu5je1LDv44pU+v0VEv7a
ODRZes5rNOoWpOK77nBPK2KpKbEPaXhW74d0bfINut1Ioi35VJv3sHrzEBSPSPa7
gzjOVMLG7MRC97Yq3ZX3o/mBxsh1pCQc2t0fuWT88s/TOp/b/IrUMbeW83yI9RQm
EVihNNfWZy6cBBJzh3k6ni/dpsw+1Q2jUTmqjgmUG+0NFnYsApFhSgP1Cp17ZFGh
x+PlPU+noz0BVODUocquXoTBlHadHAPBE0W3FCLHVy97s82xeOM2jXtHko06rT/S
d4jNcKluD3OWfAETc3uPoUhLbzexfokY6CH8O7N/w/UuJ7xrkNsFvOV/49dELzWj
ZtcyvTS15pyDOP6HSh3TccUDJNCBtvFu+QFEC36C5+pOwOE6LB/lcXpBOPCPaAti
dUH92v3g/3okpGm6THIAc+wD2Eeg5VFPCdDYAXr41Ex6+8Q4dPhcD0p6SVb4pf87
czUXmQOK65+KNAjtstniP5o49zMNE/R4USbcoNtwbS7eohtJ3kMJuqxzNxA+9fJC
7iR+i1vY8U+3VuPnbegoeA+BRkZ708BxvLijOg856aG39m54ol+ispiPS//ROZKw
NAvAOAavof0kic1D2w/NHjuJLiSlsJ/qQy1VqnVEKqz+NX6iUOjPkoDmbTolt/fM
DLMS79mOGYaiDQoURaznTu+Y6G51u76SnCwWnWvA5ny9UkIMZnPLrOXloPrtnpm9
wSC0szDYp2H8kknSqoo6WyQ1dAqGbawlruI442RQz0ZADbYKuo/kbDkXTJM1ltHY
hYRlaoKrkt0NwJMABWJDChnD5NsDnmCu/JTwANM4oTusw07T7s2PlY4zOozF8eOp
aXoNh2f7PTwWvbvi13KZf/nZREdabkpszOgne0Xds9JXYOTlJ4+T6j9JVGfMHdbi
dXnA4fXa2FYx4e+QjXVb8FpfZGubEye4BD/VT+eLMeOMIYCul7FCZHZ8qUcKjKLE
Tl/gPP7MD1MUBE007xkJX4IxcaCD5L7aGFm7IFADtiwvBurPdY2WzQh61ysCFM2r
TDkfOGbrmyQquQdypaXfJunnH5NZM09GJ2Ea9kiG3GrGNoUYywn/mHOZuShmwL9+
QU65pd6WP02hOG/B67D0sCkPLm76DyowHw/D3sD0Ra26e4qZSvx/ycsHThVH97hC
HrBjSWwkeix5Rngeli0wpC1St89YBzv396EWV32yYURUieCg4by5ierLEi2heAth
/+3uy2G5o7DyZnqJeyKItqQJ44u7ERvu1l7lWxSRJ6XNuNXaqZ8oro7YmAWhMjZK
Y/A/yp/DIBwj02WOSDOZKiP3KRropYXcPHZWx4TjmrkNzDyy7/TRPtyw5rlatoPH
BJUt3MCtsl3g72nBRdnxXbd2FNFh1mMPbNFJYDFrHxBM3svHtwbUvHqFYQvFVUHu
IiT7aWh/rL6p+zbaKF4Jik3unwyuGQSXgNdnS40sU5Q74mLnT0jqpeglzI/DW4Cd
HWGkbxlJLhvvkV5yqvPL3sCWb72n0BdX01PKGxjavSHB/PxhC59gq3eOfQdvUl+p
iTpu3u2JutM9+lR6GlPsuiVAmjxz2oJ2gQnOX8CBHCpCmUp8G+Hsp5KUpB8FXWNL
KfKoy+TWsJJffeZuo32i+dnGa1RekwGjDYFUiskkZrXCV4KqQTfpJSrBsnGA74uA
JvjpfFtkQllbhO3s4Pr71Bc4HTfpw2atKSaSN1oXEDq8PayIpukak+fr7pXvYgVC
xfsx6pNAnwlIZikkr4auX7KU3TLLzsHl8GmyIErx7QORrWeWiqnY8bIXgCZTz/Hb
dnig8GBj2tkXxM0jmJCiE9X9DJk7nBtxNPyVICaDXvKYhovSqPoGU6Cp7amChIRI
Xo2Qx2i/dnjpEbeTQaNhqypFS4/EtRkLyZfyUQFGTo2DXYGqkdICHI4yS8sJSfAa
Xx1CICCa8TU3k0alY5Cnq47LioCVqDA+fKIpOSd+djbPpTVFhX0jzhgqiF6RKPqu
A5l7X3e3Zw9U+kEQ9Wghb+6pq0cQ5JlkodkZGhZgsaUUubn7VUpzlxyRXz1sw8sC
bZIPN8sBOqkjU7gcKNbNipeZD2xzNxibDW8e3uIFyaOICHycmFynqyQWEqAp9yzf
5sNVLKq8NMxJoAFah70kNar7FMHu4bneXIH8LZNuyV9KEvg9dKMjjoe/c73HOhg0
xeX272SnCbMeuw6x339reJVjqWh/cT3AgFKgG0tPvo73MJRx72vQn7gtUfbytyHi
sHrZguiVzC1eUlsDEtwf8htxBPyFR4cJnLpb0jH4haqKMk4Ii5XWNZL8+LFizW5r
Hwb8h+33ztu31Q180Ze3z7rdMAWV3SorZuEcgPlEN8OSPQGGINSUgOIoH4VhzV7z
etMrUpW3NHORyO/HpbKLHAELVzafEK/TKpLD+LqN0IUUMxYwQBmbME3RqWOYipwl
tQgPwmX6pQe5Nl1pfFA8ucCPq8jqEz77dlrhrR88pD8cjuFHD/MKwuOoH8VDjabD
HEzxwf8TkDgWRYQDp+3qJs/kdT2HabYqLgi/5JHmEbs9mA/IdbmO8JczQbU6Gzmw
1lcRqQ1GlXzBJTQIEYNowe4VdDpUVcJDoIDFolsWDGnVOgK5H66MVGXBJfB1ETJl
gXffCLLqwv67CRtoeuS8oqTzl1sUjLk5UJBotrrmWycMICa3shZGYXf/3T01ID7K
/PnqGqQDsYyeNAjDaGK1sQazVl0W9vsnOsDBQYiacj9LDiwskxjz3cGVw7YrpLnh
FiF0v8BHR2iGXvU3JThRJlHyy3QCa6BSg7LOmhBMtPMCO7JtE9TWzRXyIHNZDK6L
F8GtM23LiOT+6A3W1K7hQL1oCiJ4VHl+vEIu9k/Sn69QFoOXXnwd4IrFegO2y+Je
97UrUaEeJWZtzZM0dUvjSGfD7jTpEAktcbctMCt1vZTmNoS+gq2iXGe0y/KWz1tw
mXgIe8CtQlpjk8lurN6bAOD5XNRRvQEcXSgmbZLa9b9otoYXtr+wWnbUfN9tTcOZ
RAelJnGuYy8BsoWfz4EUvRxdyhFjS3UHjciIs8y9+IjdbNvj6pUO5km/DpN/71fT
FvCiWpcYjZUGczCOZkYfV2IYOFO1UIAlYO80V26GiGrTgGr41Kxbbs/dNKu90mNc
B0dTQMV0uTi4L8abAOccLJ9QMrvBETm9uCDoBbIYt21PJba3tdnxKvo4kJ5rE9M5
yDOOQ/3Fzw/uFMarsBayT+i9888zQhUtetW4GsEx+NuDDUkY9e/9YYWS4qVbf3rZ
0EwICPER0vTNPG+m7EFpHjcoXg/5+nLbvm29uSUcE1D40/Ow2hOaWv/s6n9nhHLz
vgsdlRchRJ6hzl+ldfJrWEniLus91KwaILnSVUd8dUlKXjl9N7aGfFFUVNyDbhj5
NpFQkTCDUSAiZgyqwnvNVOHQp+v7h18XZKAWmOssEh4xmNFxMS3txuxwmCYnSo0r
gkoWiFQhUgBDiICi6DTUsHWX8VM8fvbelRP2wVIqyNazvnJnz+a7NWtP1cXSa1rH
suAAcDzvLjyR0ZZOwefIk7TIqANtLkZP8/NrhB9Iol82tNWLC60Djq98Y95J90T2
E8DFOp1fr7suQ1dob9f2NlMAkN08KcOJioMGRAuVlrXV2/x/IodhC8v5c/OAJulx
Gw7vHhAi3H2vp5+ESrw04qKmnwbTfdCmkELMFFxotSH1tK3S9TWE9Au1CYH++b06
OJSz5Bn5Z87jqDVlZPHBk2r/y+PCH2MnIf54N81iEeUI3/J42CGwomvw1wHL7mHm
F9zfuT+MvpTwakhYDSPoB/l/ub/6ipyzjYeeM9d6OHjZEGTrYHPSBYh4gD5ZsV8l
ss9wJODOC7hBg3FUSjG+h4/tSYdnLefjre9WEbazUO/XDD4JNS16nh2wpmedeAj3
r4W15FAXinVGlKRQw5QX3lHo+h24lSpdTI+Suy2PFh4UxU4MJiI83TyacwjiPJJt
jav1OjDQzxYagKE1l2K9pVNwr62zMATLfH0qwGaT+VrB77EDzTTfMgp07rsfvFau
VjBdlaIldQXFmaRMRxpU5eSSh1IEbhGyRJurS6v+AhtR1c9NIDo1uHdUgBSOyeEl
nPVU5iBRDjgvbh6ZI400Y/dmZ/+O7gvD5BsPv2H50P0/yjRg7CtaWgyWdVdM7leB
QeaaJkBfJvzC3EFurqQvdfFjIcNTdxUyN+sUPR/VsNG1nWRJMqjBXtKuP/621NYV
2gr0nhBA7FCUePlW+CMrNk2EZkHA794g31Aj+coTNGaPcJmsRbiy9m7aE4BOKbnB
Atb5xxH1fkW5D74u1KLdOmsyIuTagT7MQKWfB/vMMIfYQE83glbHLqNsv0jU4Y0w
bbNoNnyYntIVgOFeq9akjOACTLj4dL1IKKjOzH0N5nbxkXLvz84BfBw3KxRU7Cge
vI6dacBzBgNNjhms56/KC8HOZz2Q/3MIYrSp+9+YoxPAR92JRArpVxDaOsIeK6uY
Rgcpc8pfyYLkEwFlEhQhBvwVNd9xVxF3a68oofPYmzIA3RTDJNTuYxMVDRsCQY/0
JWqvXwkL30gAJmfNBfqvAMXfxboj/ERxfAP6N3oaxo9qGgV2E58OYx8aN02JtAI2
J3g2qP6CQtjUmk9E2PE7jS8BELddFTyqJh4dt0EKZ4JbafhZsMdt9VuEtoUzhikr
pByXK21DWN1BRrXCatfZDMhZVYLc4rXkfv5eYXLrDjqV+jFXHZsQJyH3XXhU/9vG
dz+d5vmcR7yqdg0icuurNx6ck4H1lNHWKhrWj7uIyKVh7OP6pz1HzOp/cTuKSr8+
vnhfKeEaIDHyLhbReZczNv0AsWVyN+zRAyuJyo+whd7u4OcmtuWlWJ19ZNGZidpe
SNmX1qWiKy7AdIv+bMgW2F08zw0dxPJn1RlybiWA7GN5adYlyqm3LJhbccEuy1Qp
sgKOcM+XdjXHaBoqycYoLL8kIUKhbi3iXI9Nq6gC5VcCi7RaCcn1TKquQikoHZq9
oNb1RdQFNILJOsA/DhaNwl5m2HTBLWfUYCVIdCIjHhZBTlZ30PRkpS8SnirHpY8z
d+Z5KmpSIjKeGHTygNUo2t2e8F9X9kPqOH7HVuTjmB9qTEI/1RRFzv8yS1KRiAP7
y5JsGgn1Uj+XwukEaNX7jZg9QWbw52QfwcJws3hgxD7RKCbsbyBqF0+ARtSYXjtq
OTmEEE5QPPj+zc3JtWZWXxcnlDMIgIjkVhvjvIJ+EBrw0u9lDKcOdGuXQK3prwsC
/RyLQVQ5zUMNcZzVAeohnfLC6YtAfObfKTzJqKJ7AkOHFYWVagDZAl272IWaDkbL
Z7xtd2l4/hYSEsnUgSYiTJdy4dLbbOioT1socigKG73MXjEKfqLbwxF5/Q/zYDno
80jz842I7HaxoVGoYNI8SScZjULM4w4fp+4b+++GhyyPrdxED3eZ4fxJVNhfToAf
uwURpjtb5aVgPH2mhNmndrFGMC9meqx8OZ3K34y9kdrAisYWX6JvyrRn2h4fBLgW
muYTtOLgcAKCJ96Wx2QoRUHZprlcEo9qB+4XVe4IMu5qXrIjqbDW5W8aBM0d8zTi
QkkELf5B4z6RWuFmJNH33R5NW493F+wx0dLxlDd7g+nW9LP+vnLSTk8/a0v/bjO+
Oeqhpsj35g5ZSIKnyGaOs/92jwiq/fSwdvkGQQSTiSzXb6TOTev/xKmjH71rAuQh
M/Dl0HYpoh1CrJlPeV4G8PEdfDwXLqD2U550SQfYcEtqdzM/y3zC/HizIp9t1LP4
nBUPlJuXGLq9NS5fKwCVpf9zGRDriPwSwZv/yhlp2D86q8Np6ZLDopGjLUM+/mTL
GUEBEEYhc3zUpFOsnCJc91Q7KrRhk6Gp28qsLhB+RWsVng+OWCT/ZSKY4FFNdgKM
B4y2DW5/4lnQAMNNidSGbxMnG0hlZa/Wh3BZPVydFblRNKLnwy8hPZ8AOC9V2pJ+
9hqZS+T99g0kYsiXiGbININbXA8g2uS04/n/WjOWG7EAcYWVQtY9uBIgucDLr3n+
bSeDkZdy4Ze/2utnjSzUEMIaAA+6idqHK1L1nu1QKT9fOEhRsa4YXNFqO/it710W
e8pOl3Kg/jB3l/BJB5jgcYG2B2JlTnrdI8D8MaZY0GWWvTev9CoDE1fhlpPUE2tj
GkZxe6VJqEQwUZPypnzKc/KoFFFzW5Hc6L9PIEzzN3ceXumj1wiJsoOZTbSCigtt
e/n+R1vWFRWiwsquelBtdcHuzs/nehdWJadwR/za+ajSrwiJYUi7kgwE50R0yRfe
pUvYbAxdwODDMXRNfwl43fD5uF9qoE8Ug4SOhM7RoOblZ+fa4P++Q9weXxasf1XQ
ZxaP1+NaTSAcvdIQ8L1zhKmkLd8izpnL1QDXZPoNSw3nYQ/qS0E1zcWad6gZ/9Xk
x2OJxOApPQyv1FEdEJfRUshaMY6QXC9G8JqA0Q8dt8zd+GQbuWuAYmI4y+qFj8S/
h9FKSBF5mkB90il6sfocI9Xx8pNzr1clwJ6oIJUdvonUtkcj5Az4L5BVqbHL+0dH
Ay42l0isUnRzrQo+8K69vIMQsgEa0V8CU/j5Ag79N67Br74Np0s7LVdQqEPyNdTf
4FsF0dBvhZFcXxXQGT+DG3Yf+cw1Pa72AgGhOY/q0LIAW5kwiYj2TzFPIVzbztth
HGx1slMc5TshJQ2gJWprzjUakRDc+FqDC8E0ox753ZgNdLiTmSHMVClTuWZ8kpIC
1NLRnY+CaSDwe+W5A3kwxurObiIxT2rnakHmRKQTyzErqlawHCyLwNzudQecci2C
cqpq+Swgb0WMydhVMIMyQy+3CWPEX0UZj64fpufCtQFSA0zBtfTwPYHxsuADjpQq
hxIPUWRemGRGtOfbIfmEzgjEwciPTwQXdaT+DE7D/YZhV1AyGECoxLFfu593YTlC
WgVdf8FjclSaZPQG1ZAvDU+qUwphoObp0i/vAIBTE1daXQ7/fLL5EN9lMhhRtmNO
20zwWL+a1Vl74lRIY/+IQaBfKKhDUfI4OUDPKiYdpwZMeWkxXXMjqLD/tPd+ip49
KgB+v+hcC8Ua/pQsNUJ4XEXyD9TsRRaZOJyb8jHsidHQzXwBi+R4gqhUGewy7cMV
q7nVIJzhW92l0wf+Uw6HtYoN4n8YXOzD5Vx/KHPKQPsuWqJC/5H1DVi68Z/bThVk
MWQNFaBDypRWKmm1XkAGwWdSqa+diAgYptl+TBG0BtQXjBDo9dMGxU9g2nJara5e
6tFaXH3YhVU5ADT73ciz9Dy5DQn6romNE0V11LkC3+5cT6sJXdoJSHBY8CnZ3m17
PVx90kUV0KVyFIJQfbxYIHojxckrUUegv62fwb1sLDGgiJJmo0srirRCQtg0q206
wx9lTPshS4mSi22cZbsmBeg+RUXWsQJT+fwfBB69wdjC2drbr6zxCNza+fBcH0sU
cijRmCiyzqlO6FSv15oGiiywRNRhO3qYwz5NajbI6IGdTqGsYEwqzPzhccbMc0/J
QSPLC1XeobSBjuJttvog/B7mH7PIOA23GuAaIe8Akix5doz8vp6tchIFrXO7lP5u
kyRgVugW2YJZ9DmnCubhiUpJAl56PooWhWeGgudry3wqgw+nYpRmVXLF3ONyTUZk
7VX/Uv1fIAA2y01Eu8UlYBtEAoTGjc77z+UByyG/uKcjX1HbyHdV3/ZsKb0AvqmW
If6nMq5tyvj6PDou9tVQ4v9QCVnLB9ta7SAIqj2VEcwRpwrWoqIs9LFIkV03eqYm
HWZ1AVdRU912UPShb/drSPGMdgdtU3QPLcwKkgrrzAbRD7C0lwNHD83lI91/C7E3
gum8tBk36J6XX6FjjSwMkpgfM44kTMBWoRmOyklcxBe19gEcLNMRH+3NcFdn4hCl
aw8Bcz7dl+zdusC0GSsxzHqWLY3sQodslgHa2P4bZn9fRZAP4ozuNEGfyHsHeZP4
E+aOEeYHwY0jVgkfXUHR/QGcTT+D5Rz5lH/S5nqrlWuRt9PO3hTbQFyHOytPlXOB
79KK/GJn+RhKu1qNTlfwmXMJAksQuHJAtu0gco2reVJAzv7DOdRUygs9t88/D4yL
XAAnK4c0dYR0aSkY0NsleNhVcZPq9G0AkEgJT+ZMY/2/ySCeUczRihrfrlghO4zh
HX8pxXMe9FvjQtu/P5UGGBIWu4B6DuABLiTla898pgi0UVKEeU/nITDsPwCo/1dO
jyymm6f0wZg99eD4BdLwr9eA+aFpvOJNcbWjc86V1WZDSAwH/9HDQ4g1Z1JWCzfs
ds0M4yZInLhbVQI4kq9wUhrmAUQoTxtYFg/Jbou2ZRviY+Ds14viyAVi/ZlnLfkk
7w0bc1UDpvQT8TCARxKU/aM7GisbXO5dWT887+UBgCC+YMERGhUofqhrjIlBJxoZ
ky4wiaaxYMN2wWqnquuz5+uFpHIyIclGfMHQSniulDCFYvRaOzd+/9SgbJ5Q/tZV
LjS5eayOAzjmKbaQsEVKHyxxsgneK3RBNh5KENEgC1XTiPPR1Uvnu3XW3T3uzEqF
gaq58WYykdsj+X9XceFt5jVklNw02iUWR/hfVxXb1X0S+XVPbAHdUKrWbofFtGV9
TIGWVQPJJCvV4Ka05uPwMdpmjUHybc2+z1sqW7nzIJ+yTn7QElm9UJgj8+tzcqyy
+8IkNx+3N7RlBo1P2cPoRav8Z98omc1bkcX9CwXqamI8IsqTOm7GjS/eRBIjuRET
UzrT6FW46vqpqDIypWM4Ft8wbcBriLWTPlO7cg/LkEfE3JzVT2dBJrR/guSB9n/X
X+fRXl+hldm9JX6RhqfuBniy/tXX9WkPcoibS8eQN+XTz3NUp2wvQG/NXM+uWVLR
wd5Y02owAcZPzOid/8tgELh2d9XWn4H/9pN7Yxc6Z1EMJbNME+v6HOuieznZjCv6
7Ra3Xk2reAIgTjPtrdjB1DAbCt4Jgtl+Jsf40fJAYTJNclSuQ1U1JDDDJYUqxLPW
JEC257MZZMsHBi/VylEpaTswg8VaAqwv47XQIcu0ZaAXXvcKrOlVa3ZbDEYYxju/
/Y91VUgTtinOGZWiYXgIFrkD+3bf2PYSJX7fscWjl6AnTlAjzTKEDzoG21gMIoX9
G71rGxs1gWnYtPSpAuSdfMn+XKkJLwc860TwmqzA4gkYlhyKIDDUw7ETeF6lRqEp
/kL2Topoi2hNA1YApscatUz7Uvj0z9hcleuYP6t67UxH1825iAerJjZKtFyW+XFN
yg53BCZSNoaf1MBeN+m3+2yybSOeZXwOYbimLERMvN0uIgHcxBVNTZeaNpYe9Sd5
+XKHyt/Gnyag0Q3RenX1U8mn+xvvABxm1kAZ7SM66qldWCgpWTwXHtocWDyuUF6p
llqjRsymC9TwGua/sxTHig7ZZpWklBnPu1c0bc5tsa+8IQk79+3Iq53Fbu6T7WNr
vC4YmX5LJG8umAoE50dGP2TlxvwQ7H0JUuC6ipkE5+8ITXg8I7EW8M7kPux1S6hP
kM/jYB0yJHvAKfJ3Hj9UcKx4dkjblFXQ1+xS6E7cX5juqGQHTwC6axlE0N8yasvY
IsSncdILBjGpmimFr0V/kqP21tKpiYKhtAre2eIdPHDqh1b5JLubCnZSHBsWYZXa
P7Nn2hrJQ49GjByfKtBzsQ9BSRVCxgBjayPs0cuoISiWJ0XrrT2JPzB+yRvtyq50
1BsJC/PzO5RpeXjNqXj5/yzw8U4BgrH7uxePUsGfshDPndgJzrIdw5kjQMpaxr4Z
QG8oWvEs8/pKFsrU/UcXFmwTdZ5ppZYo+4VD0GtpFd+02HofO/vfNKo4vcEfTiEd
VrJPX6PwF9l1PQKBlXGIiRlyK+KqBz5vv64zhfUHTK2Xt+WlXUjnI7UMXTAjp5Uf
GDZ+x43z6z1V1KsM7nFusQKhrRt1NXg2tLV6X2vWdGTHAmdpDoouBMUh2XvZDYi2
pcPRiMVM8O9k7ObfeEafakkAjRIU13xuWQm5wr0Wz5DSEPYa+jInknxGfyebXQwm
vsakw2dDWLuizCRYdslKLWfmD1ldajUP5IU1MjK0MUhkZmNmPYeSE2MrxgOPD6nk
A1EY1K+tQ2HzocKtsQ6BMm5ByZ5l3m5DTIQi144mDV61NaDsO5gLq690gF+q7T3L
tbEJg0c8h/nr03BpvbudXzsnIYZizWLkrLtKh/waw5twOaw3ayI+wy9tiYfdiC1p
xqqg5QzLMIupOFmLaVbuFcYfzcKGPK05QkRkH9htz8bMeoQtUAby9CVnQq2Xshc4
NRnnbBYDzUjs6ULfcNPzjFmcbY/VdxH+Sz8ivTC4Svqc4ci4RKtf9994D5I8kHqc
Dp9GIWIrwlQwIN1Cu2r6Q4dZNV60YpEOpCUUN8FglEF7rzEFpVpgAIAdIT3czxzb
WsPGgSvAz+z4cPkuFnwsAdj9m1CJ3OS+0PoE7wFaCvrUXU57QykMn2pBWUst5eyf
OxBW91Cuon6yLJqGDdRwBGSU/UYdPK5zjifQW/XAnx3aN1Yred4v7YiD312cilJe
mZjYqnJ1tjKDB+gLOH1AK4AdqMUYhiX3axK02k8KW1U38neu0s3UXVT/yarJ+XMW
ZRuiorXCeBXfFsfAinKhEdf9uI91Wn7ehbzuPXEITo+8s+Rcwngro/WC8c+jBwB5
rqHrUzc54kKrHbXpdV/fLKAn2vS+3nB+g9/VFlGjzGC7MsSqN+47q8gR5J/wQOuB
vLUrg0oErZeNaYHImcbDRCeEVODBpnvi37dj6m40p2UOcu+3o67lEkmjSxvnhF5h
2/u4lgoE6NYusN1cwIt0BoNNT2VorGlQZnrLydd5Angx2tdl3TU7fKqSGwuWCofv
RqtfkV/tULh9O6JEl0nFuFf8L4jCC6OgWBkHj7DmV/d6vkxv/pQ68tBlPOAvuU/Y
Y2Hj6fUipBb5+OCfMt4nsUASplN54pB1KgmWUPRIdFOiw7kMtQcSQe6tgNhoguRq
HO+Q15vFgxqo4P4eO8riwTXH1Au4++bi2nocXNEjxna2V7d5uHUWyYxjeSczrQMU
jehsQKIv3a3g8YipN+TAYc3Diz6XvYNPGIqUdXQZfP2M52hw/63DjtLnBBjnDrnZ
lAC81tjD4X+Z+OJ44UGazDzDBKqfrJZwtw5LucSZDEaRT1ly+49B/o+jd2GjNQUf
D9l0ZPLTHrn3/jZLzzLvfquOB1X04b1u9xaHKl13xNxYjKqmnZp6tO/Dt29vViP+
hMzcV0cwb/louyKr8o8fDL+6p+EF+CyXaB6d6QjCeJy+iqn2wp2RScXAPdRs2h5a
DwRZnQsrk6UAlf2lNF+hVA637I2xJe5etrEhMDW4F8jr0fPpoEELZk7kJR0qJgfL
lXETXvoWSww+y2k//SRp/2yh1aXZDNSNgME5PXgqreEKT6R4ox3UBRnFEaX7JWxR
XWToMzk87Tvk8vO5MrAXfMS35WGeELy/Hh5ghnvhfz4gMVa5JGF7mvYlcYz3lyzH
50DaN/bmPiSQN78JT33nGff2gr28Gi86bwXSW6P20RsFjK5kOJ0xvclH2DJVd8li
2Zc8pKg6rPK7ntEVO0GEW4vIqGjisS4tR6wTXBy4mmuwRrjfARzwfJsdTg6/Rg/W
lxxqfVCBJK4QzVIGJJpf3Krk0KIkmGnMLq2zAMtVRiyl4QTZgzDZuGN91adqOYCO
A4nCmM32rGPbcvgRxqlgEXcnwy5W6cRcDTfMFfwyeze/Espm7dcXeLlR2Ky8x36n
jW0gCq43AOa2Tu2mjLU/YbUIiBJoqNXJ4O9YoVyqpIgC/4xcauxmTweAOlPVJ63X
y+ZLmXAgtsHT/yabLxygS0HTBnk8rI+AYQALGYEsN1lW6CG/EvAUJzT6fxXaZw27
xglMt4Or6N4Vb+H+fE+mYWLKobvChlhGoT4QD+v6GvjJrazoa7q89dPLLqqkaiIJ
m1yRloJ5F8ToEPqfLgTAO2XLS2+rkk7eJNIb7L5MuCYqmcvp3HWbdV2UEDj52Ns0
KDxr7aekSUWgLI2/eH8nnwb4YQN9zZtt5m0aJbHIGoe29iIqOPg11l1V61PZe5fL
cnfcxEIamARERkkWEO9cmONPysSBFRZPwBDvNVq4Dpbm3iKoqsctJCypi5OO0OmQ
TYkfkZdb5qmFbYKViAOirEztBhPdNcUtWa00Xkkp8y/JWoxd5PQ5H+hI6/seyc6Z
KpDhBQ1HT71sAmpFJtaJ99pky2B6wuoqoGn6uVGPtDLxY6g6bMwbqovopSx1jGW0
U1c1x9IbbT0DBikl4QTeSJzIsLeRQeGu4Mc/9g7FO+0NFj/kCwhxyElc2xK587PD
VAMPSBmMo52BtaCQEO4vcTaP2T3/ybUYogxHJRq2okpLseANDtHQ3GegS8GEmY7e
+9FN4YxjPv74l5Wq+aX9zEvSKqjq0X/7oznYSacez/J78xTAUeE2IOpitl2Y8o6P
LEFJqbDxmox+WRPvDi28HZsan/BlZSfiwa7iiRWyNrLqspMYolaEl57o3NeNJMYl
5hEaPnnM1vlR1NcHQCC5StdF8UUteLCkngdAihr7an0ingPCbL0IeTytowsTXcA2
ySN27Gy9wp6WRg35D0wR9V8spFK6fk1cYebIxO3IBq4sBA+CEFXmoxxpP6AvyuLw
1WUFT2CQ0FEYEm/I9y4DzFKpg8W7tLJN1Ka0gD/1RjUX35e71VUwyZw6k7dO9HSM
bZwD510LmiyVvs9wXrnVysrB8dTsA4TyBfs6nFHKBj8CKvt4V81gWvAy1iF5yEVI
XSCC+nt4zA050rBROtKTYhtNYrEoTrIqGp87mOneveElMNAcmWIG/EqFaVTipgCL
21eLiAAjJZhAccxolz1Rdfew2kZ9IILgBIfM/z7CgGVogQzd1srQ9nG/lWPHS1qP
5gxPJW+WOBazeLhWCeOVi6iutWO0QzHrzwan56DfVjtsdKos9oEub4eaCkCnKIcl
1hK3mNpR27WQZXlvtsd1As/v/nF7/fOEHfpa+d83paJio0N7mDffRoDb/xGSnp/d
zWmKi5FwlYgtTNKswKPIpysI5n3M7YCIYDstlm/ndZy1n3EActEGNJxX2VNvBAAq
ZbqLjbmaQKqGtho1fQV4oF3JxiROFR0c4Iif5mgcTRkXIGC0gR3c9uFiRSLsQlrZ
CuRQMecQP/2KXSiiqrHz54J1zbRurjsLQL5sft6nGi+gKTAn5rcDchnZeZPy2Yfo
xNaijP77WJPxWm81FM+uCw39cGteBhho0xNhk7H6OJX12WUI9YYtuw4dWJv1hRNF
2E6QEKz0qNwrUkbol5IANUQEGs18t49v5u56lM74hoKPwp+V1PVzw+K6g0iC3JHZ
VHhaoK2oBY+c/r8ODm5NPiRrWMBI83ERFY5bR0uCX2tdy1cLYD1pSqTFH1751/pk
9ktSI0kcOu7lHvcEgQW/5Nhs2w5jywPYUInZ/lrKxz6eH9Kr1P2SkqR2sFrSznlZ
uihOOvAjEPk0Uy3zN7GIuw5g1/THIyQlEBHHw+c2q9A++B1liKBn2flcPYJRJOEC
Fy8q3hKThvRHEr6xeRl1geWlpdoM/RKWZoj0vH61o0L8Mknh4hEX4K2xfn1MuBjq
2uA3ycHgUt84e6i4NatO7A4Q8jG6CRXyCkfWIIBov9X0QtJ4bYgfCES+ULRm/aDu
5BQlhlKw11ciNfEBwV69m+cf0wdaDH6YjYnwQZ51XSsmfH8fPpdNsyiNT/k1I10E
oOsZNy54/8b4S70fkc/MCv4eO1D2RSIe0HUJacFTGQA1PvDWwh2DBh3deAfws0As
cZm6HmOqII7mJIRDKbLpcd2R0cBKs+1MGT9Jm56FAb9I+21l0Lz4mZs8tT+mk2HW
4XY6rRDF1ye17h548Vg5oRxfcv8RtkG9Li6humCAJypu7Dvw2vdtmbo/27qRMvIw
HwADtRTlBbOL5kJyNixMILWLgVqjj1b4Oa/CkPdzlYPJ0GYbvSEj7NIdFfnByauB
UI0SgSBU+WxeJspXqCIYVSkob2axp9wPzCSci268Z0KLuLe3cve1y7bgTGzGPkVN
vXQnX8F5YhiS+U/bW1oLcJ98sblTTsfr5RSDH3hwL5B/yjmywGskk/7R1GeG2JsI
BYztjZgRH433eN9AWZUOsgNM1QxlDrevQcuzKo1s/khoMsGCZt0CE8jM/whn/KvW
U2zAJoXNUBLlytgpob3KsSbswWgS/kAVgaLKoG3XYfoNw736/k82RxMHk/deqCYy
o4fsF/iQm2x8nb8JqRzO/Xv+FW1jYoUKv5L35/zGJPs47WP0l7j4fTy0XKMBVErI
fHsuerjlzY7qY1bHw2Fvg7aaaxyHyM41/4c21+bdDmJO7yBwTUoCk9uVHTwaohlK
0acXHqYz/ZX0xAtmeDcDM4Z6LCWsywDClc0HwV2fj/REV/xRCt4eoI7FntuRk3w8
qANmx8uxOeV4fUo14FfXtlYdLC6kcl/9PSEwDAMBnSrxp9vQ1R4chJmcJVVB6l9c
nyaYbdQfB9BdgISzMAejDl4+qgcYOjBRj8K+Np1SBVu89M6s2XTIZUGFGf578EpD
t/hMsQD8tYYJN9fc+JZOuz0/ebJA+VgzF3x29V3ssldvCBKsob73hlKhZQHy5EXt
EwlAK2z3uggxTOaRELxKplt9m6SHoP7R6/PPe6OD2ubjkc9Lhg884pHrDBl829V4
pfgJaXBs3ou2aBLphV7t1qpKZ0VM5LwYnGzgKoUr9Wh3+dh7hicnpV23zzeY2eNO
LHAQXndRI+/TcIW6Yv1PsGImZqBCgJm8McFhOEmJHL3Ik6evCpCG6jyPagWIemh+
lMF/qGRdNM2SRCTI4sqwEFMRAy2/LDWIBV7E8IRM62mIIHNxb/EPU7mPsWNpOxkR
FGFJW7tYUhobr8nGG4HXp1fCZwGlgy2+P0rx1dZY4TaaFzU1i9gFVA65+Ff4i59A
1NXkm8UsToN5hgH/dlYnbHXPTvZD/yS/WskhcKE27KtYnXhzquzomG/V2EmfdZ8Q
ld3NYISRdS+b33FvLYM/oWvPPnIelzZe9o502nD3t7qvs2+QKXs4uVz9RYyMEch/
e2RyJAroyX43bYxhR9rXy7mtox536qsV+dD5Y2pzn3tkdAWQGTQSghWlwf8Cxzbx
8BtCG305huTETAQDFoPbpPTXPKJYVu/xbL1xCeAK7a/fgPzi2io5H8Bp7jZGe60a
f6q1UUGj7AvidQAer2XTLQtrhMERUygr/2vkqo8Eibpmw9Sx+pH/3yODnas1ZVCL
nSr0hHvBDffmkyAsh37jyknh/41Qsg63TO5otzq4C1N3plNnDUsbVmCCkHNU6xt6
q0/zc0X+r7VM3YTluvD1nEeQN4n6q5gQGNQPXGFha5ZpTkUw+HZ1LVxk0TIPNR7i
lDDFnTX3GBZ557ejm2T8hFymdJmA5zDmXbT0fr5PA8lvb5HyC84ikOJ8vHQFBdNQ
VHvFrEsYlEfen1TDuuI8cmdkfvRO527/j+TPHw7odBpxHUv4+lLfW2o9v1DoJ9cB
NlkGj7ozjv4zyZ+CacyJXcENsnY4JL3y58LoRuSGKi7EIIATeheJlkhuOGvcWEVx
QcpviJIiMxJ3bMpDTbtxj1iWVv+/p4ux6kMIdo7eQmTFIDLmPHGEkPzqJtFb2bL4
AHOljVYQdy23I81ypSPh21qMCBwh1lABlWLqZHSqx5QO/t5G9omobGgJcnupZq8i
4Atn5DnZXTXr23W5n14Tr7WmNqWiT+tmtx3X6uajQGmcFp2KMkbYyhxKZlH+Jz/E
uOiQhRS5n8GYiZx8yba5noDm5iRmxsvAJcX7BMMP1qqxAbR340NQsK1oa1P1ua75
YF1LXR/iN8vMdreYO9CRNxWaESp0X8cej9++3qgH0btyz89yeTDxqjlqeq/Q02Qp
O8bPko4UJf4OPKW7UzxEWR46Y/CYHUgCLr8Zwba319ENmoDfntym89KCcly/V0CA
JbFZK0ocd3dMNJyLCrAvgPfn3i7I/1n1tUKQyPQsU6qXryoIgltT7fuQb1oS4In7
QjZvww3RO+QhuxprbEUm46REXLFhNfeMgFKiuIQcrdMKgdJfZqtyd58yTL4DUWBb
wjp2UnTGWaKuXhDBBIVmBRZNejptS8lQZZlzkzqPsGOsus0HfXB2ZA4vNJ6/xjks
L7ogbHEMdfPuIBI+RWnH7KQgp5trGD8Ac8S8GPfDo9LGtR26BYJ3KcBmh2ycGYHh
ma/8GGlxm2pABORuoLpLVREbyHJoryQ+s2h/TtAw4d1g1Ab9CIu/FTikk0sa12Ii
+6NquOe99uX8ex2m2j57lcI097JvGqojzW/IMVSWttaQxDmt25NTpBT0Gr3wvS/N
hmqdBJp/WIBII++6GvQoLToo3QoaDA4ulUaCUbj5LSVNbWMR/eabKXl6f41B6pyk
AthRb54i4XWJW9hX7m2T9TixlNDkhYxRH3aTxpks3Lk8cqwSKQ9J5IeM1vTMJwjs
ysvkTiTQ2SWcfbQfd+PjCIZBLbzvXoY+puTH8NTzYGIba1T94g8YWxAeGe+xTlru
+kLM64l0muUO5A7QZx0TNNIQVZTSrdwrRKvNn3Q/Gd0c0vSFtc4HC0ltBEZuBuGB
k03Ba207crnIdLxtL1feC229G+VDmT7HhlE96Nvdt34tfu7pWTlG0722gumhuKs7
/GVi5SGOqDbTHGrt+et/D0JOD+QyE4ujpj1R6lWD2MiVLNkrweE+3Kz4R0TDyen8
1ubEf9qy2xAhBvp0w3WCIYSzevyyJ8MWREoHEsnneGNwV3tbrJoBjeMnvUFRb6hW
DKq2u0yUHaoELLOeQ/TZ4kdSdl0iqQcEiDr++u+yuy53nrrh8M74AC05Oz2ccZTt
d72lK9MIRdQaCRDDENI/p0SFhIqdEKwPubTSaa1sovt+XPi1cCFN4rWyRTAMFMRt
7PLj9ph7MKbV4oArR7qu3/sZqIbw/pSkCWrymyKTBHPQqYEEeDpIwIYiJspiccW7
imy16CHvA+iTRMFJ/rIiXkvFUAer4VnVLmDnucHdqZ1axQU6kaPvQQkPwKBm8ihY
xEv4F/NR/KLBaZ2/EH0FEzW+8lN3yIndBIJu4oQFap/pnLFcAaYLcBR9N1AAV5IC
oC0k0tWJJ5MwngQg30XOGwzXqwAbaSJda+IWxN2NYmTvuIh8OKO7NrQLI/VgIrbR
QpolI5LzoCbTz4iONqo2cd905f6KmXzLQVtk2NRersN4xH/tKaBA6/647vIbgtqt
QaGfUlhavEl3/7Rs6yYN183TGcIyFeoWW55TwMB2b5G8hOcUvt7h12pn0lU7538t
J7ITTd6f3vIo/DWaiq2pDhy+f/n/pMbkhg+UXefDSHYhsZVMOI7up+jnSGKrFZz7
Y+AbMoZqNzBY4+Fsh5qED9OzlXhr+y5ecwdgBpKI0/pgXnaALapgdBnbDIm9LQgI
dveM9AIumPQPyr8cUdB4Ca4N6urV6Ud8QYSHFlDEb6u2RdiwNgIwvfpbcE9cHH/e
f+WScqnTk2bdVvSX/MlcXsxsSfApuDFmD3ji7XJ+rnZPeZJR6VkRpOgWgHxxvCSg
wdSOiT+nmtFBnbU0n4Xq1zgU6U2ptRt96ydlU2oAx6GJRqLpRIYNCFiy64OLgvWy
4UPNAKT+5I2ZelrCpA62iF2KRK8E0yHH0mQTCArwwWpg/mlLv0SbM2yIBkCJqCkl
4/RIkGIitvb5rKoYcPn3gBl69zFiBO+H1ox+FlRzGZSDGTZaYp56X+V23zdMghZz
PYmXMqyDrrIZuvPN38aIP3BSUyyECa4cn4L6HFT0L09yJHTCP0thIBTt/U33bCTF
zuVD6AqkRhXgSgHBVY/PaVo47qFsm9b+z1p1E844vb345PtR+LQ4yWrFXPyE5h2b
pdCBnNH4QWdWC3S1aYuYjerLz40Pxyffex3+rORCnFxv2GWpKA8jbaENtlLMQEHi
9LDUnIAem+bJXXmgqhEtWH95FbI6wVGgDQ+Q5kaZjBbcBt/3zaqPxdMuDEDCpUV6
QEALaFN6iol/vHIEazkdma2nzsGrBSifEFGg2ACaSoLA5WzYNShBLZz/RcGmgWMY
V1+K1+t0k68dk7zJCQYvd6e3ufimTcqLEf3M/m3bxpmFcT5eQTvxZN8oAekizm64
tSuJZ0WKB1QajqsPn4peGA4zttF3VK6wsKxa2OrG4bx4eU3htkEUREiW6Uqbtt63
3BbYfjn4MVHtTAEdpKAAsLLFCpxHfjax3xC0Z6AjX3sKmx6wz5LmtevdUBuv3arn
OxPNVla2thx8CjuA3qIRZMBX2XyOJUOoMBXH7eU9rQ9E89by0PLDlKwJqktUIbtQ
H8/k2mzWGxZhY/i7jsEWqwCIlCuBd26M2i4KB2+LV543zxEbJgV8PJptdf3dlGap
43OxdiJmDMh9JZ73FUxxF5MlR4K5Tj+XNypmOAKyFUAp6da2f1GEMbwmMU8RyDK0
4IjY1x9PeNpGmmcLMwnId/OE2fKpKU9e29A8T3xIkHrFES+vnOZzk4crQFSPxqka
1SEdyV++rdnujtcIzC5JXQjYf0ZGF8EZGvxBXkKVVM7UVWnc90HuCKckg/Zd/NyZ
sm4C4397yov9mSvKlt7BbDVTwKhvhP+dzA+xf5A/7AJuJW6VFexsbqbRRUzD4c4G
SqpyluNBpEZQFZaLoZvDPO130nNzmxAkXACnC+hVdJ4VL4evhNmCEnbz43Quihqx
sqqI7muftf/FCjZxBUxUohnQyMOQFoFcgjTGU50Ei+0+D0dWPYgH6mdAzcay2WCA
YzpdqorR0hGBZQzZIy+lnM/9bgOctvraOSMbNicbbYX5mMJ+clT4A57PzhvozPxz
BjxWIQv6x1GFTeDIZLkfc2uubZauJA1L0szwm6uoIP4pR682ynQaNXkIm8mWyWA1
KHO7iR5/9tcWEDrZThOOPa3BPpltkAHzPOoWsNAQBRosZFb9IRTCKreN4aoJv3n0
vqEPW3itW0jjd1aVDz5ynXylmf5IsF3MXdoN+x2y7buU2s8n8OJdX8Z8AzZaWhgX
D9RpNlwU3QOOgzlLCTm8R2Q6dSBfPLtnI8pzGQTdLJUeTilPyLAl+VmYpj3YNr5K
rXXDOVBdgHiw/soTIjqKE3uX8bQyYtpKJaZ5tgAPmimwvqU7fCzG+doabCES8rmW
2RRtIKFwOc3Aubet1NFmbCLn0VTIEUfUaOhR+2V4u9We+LWB89I47AuaiOS/76Kp
7TOu10c+7HHhtCIEVOkh1GKYKVMAFaZt0zSgHO78xpnfX1c8GsC2gHGcLDt3zgNq
qjfUyhYpHC+TuRrJ7R4FUMg1Oohq8d2N9CD7488e3XJmk/aGGNbEWrdSClK8EZe3
PoPQSGKdaf+SUVON/QOZV/7/hX/jRVLPkLCDXf3ji3kPWirmh4dj/8Y/Y6K6tlGG
bbqVwg+jlKwC2uB7CGiLtpqAe54uOHzDwj0jgGa0IfjdyyIHtxPy8IbEWSXRADTU
VanPtVaNJZ+eTV6SlPTkcnvMEteHjubYuCIMAZm0R0DsxY1SeY0tx7UQQlqD7vyw
mVUp9fTNWyik1yNAh97NpKV+E+RHrCmYZ6dmsbTebqwHRmxlcw9bEUYvisTF1YXd
I08NwjTEUHC0QrGxzHB9XDPbCfLUzn8ZAPHvfT2BMPI4YeTLJxOuh8SsE5MZJKZg
s19jwLTjtOTa8+wEemc07BwTWy+vCCVITqXa1A+p8kOtuSNMwRUC6yuo1X/bA+G5
NnsUbRhCr46PHdnw7qYKUN5xZsP1tKG1R9IlPt0f7KE2VT9EjijqQMrYouzQlFuA
qFRaou0MssQmUFs5Nhx+gKapjvi7gux6PuZItrgKqW0VAoAi7mLfJ7NUMcV1mn4F
Jvxu6MTah2jUEntnKw3NUpPPp+1AFZ6NhYCNifQGHXfBlFyc3lWeoTgsbEi2sA14
8woVhx0FVMyTXFJt8E9Jq7UgmsdO6MphdhzGYyu8zne2vxYKlTRhns1JdHybioj4
RO1/rQJ/d5ZuGQZpC17zMN76TFFNv3t96nBtA7EYVpiMoY2mR91OQbplqzXpBbxY
nZ9MGgEamgXEMQtjwoVskwxAtXVb/mnfGNuazMVFb2byd2+8auxg9B/zwEoLh6ys
dfXGZM0wTxFh61GpV9KBcoI4WALhvUZBXc5GUl5u/ohITIPQBkjpzDVYuaXtI+SZ
6edyxVux8attya8ncYbdC9nbyiKEUQJG60YBEbt3sinji/nnwV1tyMZ1KGPMKtu2
TYhIoTzFhvS+o0RUkYuI83qfABcfBNuDaC4FpFWyeSxjOrott7SE0y9N3xqBCGGc
/aVC06EusskalWDl6zj82dJizIbCfyKeGkrnFOu9/lZf7R7dIslX8LK0XPkF7b80
9tRDtnzK4D/0oihrGZu0GI6NPZQFG+l76pXf7rjrFZHOnAZg1O32YSPvnwTPHCwL
N1jVgols4ZyYki0G94hX8pOfNECg0h1gZqtZnX912f2Suq+KMOYUKlOiuuyLP0oV
nSH+2B9UWChzzBZJXhk94/aAJSNAus4R4zcLfF2VsbQAbmisDM4f3La1zgKs73jt
UN+zUnQRNyXot4Sz3ddTF7b/8wPNA2j8xVCCC6F0PBVPViEZ36lcNwqSQgmhXv/S
KI5THZncuHkMJZDbkzkTymhDZt7gDuhstUaWBz7r/YZFWCxudmEDEBDlh8N+8cro
q+g4lza1LzVtJiXEikscYSnlWj1V5kWVn9kCyZVOCTmVBBd69d6w9H/uDcqaVcWw
+4pPH2tExgMzLZPRnh3OTV26KiotQejFcf3lmdJ81lU/QmRF3CtmntZtN9OYD+e4
Gu1JXztSYxtV0B9RF+oNfYwC0InNv1XoP1cJfDOtMFI8Fo12ZtXEAHy9IPi5nh2b
4rccRiv1Hk01ZkdW+zpVfjIi4r43AKb6jW00GKRWsX81NO9sQqDW4xL2+Wf44SBD
YaQMJ4L5eqrCRzHMTrKh6iA0AFzzPIHv6JK2LcS7ENLDxysMLWr17TJNHyxb5PMX
kRxIqretoyGqJi513eILKCD803KyDbe1Q/RNjQ0S5TLXLxRwCHLiKx3fMgN1GVJ/
ebm6XXXwShQHs8smEXhtxA4b57qevnYt42VnfeAejp4P+/WWAnHE6Ae9AiYA2tUu
nVWvmHw1fgierWFtbgkLFgcE1gsm0OaD+MXmuFxddmNOHM8M1MmdusU9PUYd2Fzc
BDjDZzkSNwIZM30rPXtMclHxva3cxwL/4dBNy5dZcd7VZwDNkL8ePD0swWSccHfd
ZVgO8k29bP/tB4n6if913EpE1efcWOifD5k9p0U30uaE1GhHqC26lTnSdbI8Xx9o
c40omMSJ36s/6bV/6Gvy6UyRmcYKPuJSJOGEoF+fc4Vdju8AuEIgjHt3UwLEJtYw
SB0jH0M86AFZkFOgi0shp/JAo1miQkkdInvczDK7FZxfwOVlXIDQ3/ApLXPvqMKz
eqBo6TKghpGBHgudZ3ceBmi45ygIeBx1nQ4Reto+Rs1BFz2uWXonJxZww23Fa4a/
OBn+oH668npPYsiDcaYI41CLnEIigLz0TpVlnclNLjb2z+y32Xj3/D0QcDnAZDyJ
8kN2F3btcv53GMAtpcF/Rali1FvepF9sb/cgP7FQXz6RQI7tYinh8/YiTFCLau8V
O+AbrAqxeMOhfsadu4MVF5GPtjHhWOaUeZqdHJe3SwEnnQSY4MlQJH5F1c4MkAlb
D55y+egsZCLi0jnQDkzxobpXRl38u8QUQ+ht9t7MIXNjHQc8ggiqL4dq7P6oheBh
+t1+o4+TYrTqk1geoG3rHHHWLQ3dHsyFgVsHFw2/Z80uAshMZg3eaX1hAOpJsdhS
ejuJ5rDqWCI0PAcLF+uY7oTgFgmuikjeRaCgCDcJUZk8hRmOovwzavRobqVJULm9
6pmBx2/h6tHRJN68upXoM3NJ5nMe3F1a+KuLcvgBmcx3PAwLih4jOmZEjQvP0TWq
ZXoaP6hjDIB7geW5Sn7520kbwRjd0kTNWFQOTabdSuA10zRVLhEeRW1AkzrLuQTz
E+PZNaFZ1p8Amf19v8rjUQoBIad0pTFLswzoXxXiprxkOVP1GwOCznyCpg++43WJ
Kg5V9wbBX1FP6Tk04meLLlNTkl1oh6UaS3exKZObsu0V+6Kl2PgW7imuJ4YiAOdT
PO7MkyXHNBY1IKESd48uZffiYw+5p+GKATMjmIRNwKCBtWXOB+5OkgTZiOm57O3T
fKdo9rx13hKDDSVANB9QK6r8O6IiW84U+c6Ieo1V/V+XeLyBZIcI44imMMDjyL3m
lYk0w0qDpe3Qx35EAi/vb0BLWj0DWtMfU6eauVschglE6C6kfVakC4FBy9npATBH
VRpHk6LjgsjIDHk6eFa4CmL2Zrh1mhVe0k0wAyr7AjQgw5NOUMSAy/4WB6z60kkc
XZNO3SsMYayQWLUf55ZVTIbzuDQXvxjF8Np5BvL7HqI6T182/WL0Md1HbCeo5csq
etQ+Zlq814aFnahofeqwW8J3zE/4AsVBycni+nvVAQXUUBK5otlBqlE3fQElljuB
/EsNQ3zLaDL2bxsXupBwqgulQLloFaTCInH2oVHCKkIFyCQgKcB+eLfW7DMrmnvQ
TN3sNAB+bWzYV1gUSo61FjWG6pJu7hjFn4xvjJMVNtFg/ftCa7E86m5n0jEwcshE
aZPnVKYepY5o/UHdUUBjfpkX9Z9j3HC5rebpS1LshCC5p/4u36cTJMpF0ORcSGLO
OIbJgyQGX26BTAryqFOErwnXXFR0OLtpbOUm1dGsRZjOy/aZCjBOrwBQhxIlQ4Md
q8qC/BG33SpieDxq5dlrGqrvL16hIO0nBNL4HcxgsQcgj7Fpg7wdmVhN6GudR/4k
ohFOeZYcsl1uMaG9co1/IV8JqyrHWyCj373ZYr07HFVm/qeRNJ17lKs26wKIALRz
90lTczXN41QOZQAc+Hk0QGOZiw2OH+PkaLNaPUrjds/n/ZTtJ2U/wJ7hIxVJ1UVd
KRjvJByXnkZuKvgeBwFrfDGJ7vpwPrrzVKHngKNK8BlpCUHtkGdD0InAzIVzBk6r
KsiZ4aqVnPzOefIwLbAGOgJrHZtpfJccaKUc+0E++ueN3KXUEvWt66kajRQ7hTry
MUYas7sHNiRuX/rLmNgp6YwQjfWAhCMJCN5TbsdT0bUPBL6BkzZMZq4p9n8OXGJM
tQGdKZx/v6KHFqnzOhIfejA/jCvSY1P551VBmGwxVElQcJG5Yk7OwcOVIrZ9UH43
J5zIMSXT3LmJKdexAmOwSgVH1Qmdv1fUnbcHAJxfnCpsNBjSRz0AOgANAhbQ0O8k
u+LhyR6mdUmBUHSLlk2nFaWpw5QYIhCKqfTr1jsvVb0u8EB3nw7o8T/6A1UOGfyK
9k0AOuTvFGLVfNoHuLuuaCf2GbJF1RHBlp4+bBW+c4lNlXHJqLkEL5XauN/BzqjQ
GA7A9i4K5aqVhj4AdzZ71R1BWg0A/9EJ1DpNlWH/5uguXTqqcq6vT+ZHAB1WkynW
DDWQ4SzVhqipoLZrvgK+9kVsXvePuBHYV0N918+FMoTb3RfBYHWcBdrutgTedluG
L+kBun/IGd1DXfTZtz+lboH5GA688UMWA/7axq2oeHUB9CuRLj/HDogV6iQ5cxu7
+IQk4Eib1u3O5e4POEo24g/4l0okrtTELmQ4FOzyJzONbnLrFpQ69vUU/R31wBjE
kxAAaFi1mvRaTnXAUqiH0wv1j7DsvzuQpixX8UkuacuuSbF5P3WJC3/xG79ywUv0
bfIBYjz7QxJSL6TKXAoQIyH6GfzGYUvyLCnSnMdyKh1ENkY/Jw5UlhBmtQe07I98
6/cjuA8USSIJJt/V2EXCb+1izVje1Um9HW6IH8iCh/kfWjrPhjCsnBU+dxuzXVwM
Ak05uTX7o6N9FWPle7PpZQxNyumWsCLgQfCz2k1c10HOefZi5qDJ9hPFZ7LwKDh4
kcDG19htKy/rk/8HXvSxejZ7elJQLmGVExPhNyP2kvUgxHjEwnwPU7jYMuDd22rj
wAqrljnJ8Ns+srHTKNcPojAdwRW+jYv7OwcwWRoHa+DDJB3QRITTsxn+AJhY21Dl
4XQ81LtwPdSyUHiqxr/mgR6mgRtoTVFFPA5iagUsEJiLWATsHTWM7qDcYc1npX2G
mCRyFMGrG7ErBp/ODVcSTDc2SFL/SbDOd9xgAvHECdK47LLLqg6FOU7oLPbhMGAL
Pxs2U2/AojJWeqTyjQZMxHWg3uMtP7PwsMNUTwUvFLL9zumZr3uLtutIOEJ56Gxq
vsg8AfDCREoZC+hxny2efUT2hTDC9UpkQhhJeNciyCsxGPXhLsf+S5IPmT1ydbpf
T1uI4lpi9G2Xavsc1P8Yg5LaeCPbMRrXc/jGJL3RxrMGQvRw8SFyWMGM1hjBsIcp
3CPlHdMqJOF6l0nMfsbTjgn3u0kP6jxWT1gWxfQoe+R/By10S/B9jKDNniPpHHei
6vkdzzOnF0cvW0zUVVmQh9jTCd6PfbA2mjHQWoCpkZea/u8oHh0obHPF2TdfkZZq
hbWqnyKbhzrW7at7P6Fwm9fctK/JOjt8OYbsnQiWkmxnmq8eQbbfeMlRWmotxx3t
qUh6u1QHNrx9KDoPgx7PkFbpRLoXg7jlNlz49S9ADP5LTC/4e8oXbJX4CC+oGoue
hThjSEuoRHspEhh6Pd5SlrUHnWYBj58JmL3R/U3HsKbPpBvP4LTDT0GRSMAQVl3G
AlZtxFa4/dGp05FDYk/tuPakEcanJH0KXVa/SiwwEnom98h5q1tteYCjjpBlfPMV
GQpIv4m+yWuREZRH69Vg7TaX9gyjL+5kWslM2P0SP2oreeAIMe1v2kSe+ShaSZ9T
+vOWl0ZtevYxZRiajB9ebTTKV9a3Tk+1tApKC2bN7Qq51+nq0eebME0Tbh7Wi1VW
uCxDla8LztE4eC3W8xTdmp1kbqfBI+vtgoYo9cFTVhOdAGzAHEHK7Go9lCPRvDtZ
uJe/dJHqIawJ/ohjIhBVTYYrm1zEtqT3dHfQZFZRoWl0H1ceT0vse01xmB005Ny/
5JkjciKilIEDHeGsvpqMkOC9YFDua7MSYlSILFnmz8TB3F4XQ2lyQ0rZ78aDmLtn
ygQg8Hmrs5ndFdfQPiIp9CXkLyIDL9ZTBgIeGdUKX+XiSttzZiK7BJu4iN3t/1Cw
wIwknM6yULEjuhm+x+ifIeKY/o5LElDeqvX0yGKXI/qSoa9PII9ejmy8l5Z8NdXm
VOlHGtrFIRWiMn3m1tm02junY+ktPymE1qu7feqMdhKt8xax9/gLDBXCVsN6t744
G3455XK8P+qZqYv3JaLfLXCOmvYCKxVcbLQPdbPl/eeE5BRkqJiiUtfNguwjxpZB
g8fGhwx9QicD7X7MVytUy0ofrGnEOWz4KKkbqeXnVZO4rq5lYytqbnbXm4n2LM+u
B2QwXRVnyrtGAqCTw+k5JQu5iGfupSyS09oWEU+BNMjwnnL7EffCqbO8R0NILUrU
z75Jl/ITElf8jbdr48NolgOW8dw3iUMMP/BFalryPAG+IuN246Mgs/IBlqKdmxW/
7vNYZ6+/sfrXT28Lhh/Mgz+3ibb8L1bDQQrCqo2DTBvsKt1MKFDzKt1fDWovSIuK
57evrTNLbWwDq96yibWKDwT0Wi4ifYEXzxOjVQMtGYnkCRmHe8YaPDIFawKMYc4u
fvkpHTwF0rZ9eycUF1SzOJg9VWv77TP9om6+F2KZtks7LETKxQbSGoZ/x/uXK3nm
fd76ODEEZKtvliTBYNW22G3HaV/2TaLX6LqI70v2vKpLsnTCGErJlgCAIsyVkZ26
ekLZcCQYFXgVuTxocmbNLpgccNxLpaZciGaJweruRUAKmnw58856TRyD5BYGKyme
Zjj+y2M8vz/2jhsOcxezcj5RV+QapFu52z7ZULzlVJLy1IJC7EuldNF/RJjMBBAi
2LSquWmSWVdFiOzvD+v5v4DlIBCxbGPQoQXifucIw5DYqQBV1ZaxjjtzZZV2KAGo
QhPxPxOrQ9fk9MPtX3GM51Eygi6COdllYXdRgn6dK9hfijaa7zqmT4TEITNXoC/L
auHrmYhFHMAhNaFoLtCGscXwcPSNcye1p5pv5BxJHwuWmEL3hIImf3tUS56OGG4M
9lr8IKlYGNQcRJ3RsFqPD98KabADnrvEdNadpuEcXYZtSr/jkiAvtIPm8a2D7ojs
7fBleHDDJhNxvassvdmd02lAX9bdZNiwkO7gANm99LQ4CGubJ8H7qDV9XON0sULh
irCl9PKMKDG6CmYgaNuRGEgVZ1QXse184YQ5SMTJVCNbxzVIKUYfgBtsbqejcLM4
ADcQ7XzAv/SfDJfUOQgTdXsg8w84gmCOkdfxSzKjCuVJys7yJdjtWh2EF1riZx0T
m8cv2U1ilv9LqQLYlMiTiLIItNA8ZU0ioD/XOEJCvRGMJVK52jEhI7S5wLijA/0l
3INEFk6Zt1lFlJVgnXiBLNTnX0v9IvqoRmvIJQPSBQ9Z+jqJF6beDiQC+3GptOGU
3Sa/CULVkpVtb3ZTpfjWTk9C5FSf0NGxancV7c+LcpTf03spNEIlMVa3X+vAJWVI
DrbRxbafHi/OgkX57MbO9TiJIOlI7GuKqTuzxoS4qpPFGiivr1kv/cE38vYaAP7E
616MLjCt9BevQIaW7w+UsWv3LJUp7WfcnIGKEuq+kOXh4vfNz+DHBYmpGxrx8pgU
ojM//zAKoNIguFR9WKLe22UGKB8AUGSD6CjU8jkrbyFavu6vD9zx1MjwkOPcDlyP
WWBpccTIzNFsxr8CaJCL+HQ4fdDxJSfEa/cv4Pc/+mQ7xr5QTIcFa5IC8ddaxWIJ
LjbrVLsLzOds1kxL4Q3B8w/UHSSXg0iHU+JzqSLa1cvTc4no4jzKdySF0ZHc4EP9
w4SfDG/P1+o8ltHyJMrWdETdr2cUEQEAGOyFps9PJog328HkwMMnjb6Ay+pASIe9
h1H3f31S/kzZIl6SLprMT9+N0nkUaUiYx9jWrYMoGPtg73r5i/qSpxhnsQ6Y5llr
3+4oGtuaXLpxIcGVrqste38JlYF1RsL9n00vjl1eIN8Wj94mNpVEDeCYm58vZ8A+
XvPHQDDYLB7NJA8fmlbh5dqSKDU2cdlSGTs7+o5bjXcyXjiYLqzZa7BV2gLkUCy8
hzf5xrUacunxe15RYB1xrWStH3/80EF2xdGrc7e21MuWO6k2DUVjEsJXZfS+QT6I
SNetTWnkqKKcpJsfpAk8eiIr79ziGP6lb0ffrj/W/slKYMSZry6OxGP0GL8nfKHa
G3m2fv7xWr9JcilGTjJ9l1p7L/VnWBbUbjK9Lub+F3CqLOZCrmM9Vfx8WuMlGkd9
+BCNds0raoxRzQwNtZAe6Ipf//KlKDvoL4GPmPc2rNXAZ4W5zy2V6tSto2dgCCcW
GzrJi+zilmnarXkt0ivQ5qODVttKazfsWqYQhoSlzuoEggBdFqqwb1ISNPeCtrxk
yXCB/Yb9gR8+cTS4uKMi1q3B3RO063q5LdV6tHQn4hQTzp+AdlnCea+zxnIYqG3N
IiEaRIT0TtKlMPh5pChx+YTmhcFXxjDtay7qT2zOg2xxl0ombxKzG2ZN38cymzXr
TOnKt+yD48YHBM5g46qiduqBdx3y3fxEnYLz6vdyHNXM/OZmpdlReAGXlCqC2GIY
1qOHwa043/x1XuU4JHZKRAvUz5kDtrcJc+FlqI67sNQJesZV9tGtsWuL1Zh2JIay
xm3x2WnwT3IGsAnCnvWZXgPpzg/ifcT6eDi5WXGv/xTsQkTD1sVuJQF0ZIm/mff4
fyloClTY/V326epR0zFVo71P8O1J7GhB0UMhLiQEdceKAUosBW9JXSQu76EGuEIP
PmXKYYe0V3fizolyRuzoQ9Qr6C/pmIRSwWH1P+JAABsO8ZRnhcDrcvKIjnywN+vO
BbZ3QHc/aoEwOeqcqtgI3Szj7/CnZhnJioxpHyHlngULm3QxAeO1x4Z0/Uhdw13o
POc9KJ5l36vxa57bpwyx5QgCnnmo8M+mPd1AeXWgCBDvoTq4P4SCDI2B8/Ws64WY
Ff668FNxC/1a2B1WYlSEsjsv0CByck+9BsYaGYOWbXr146WAniLyokiICujusdkV
lCiIAXwNHUUqZO4p8k25kN//oO1A290XDi6xzqXkKQXC10ylWr8QSymIzbvy7Zwd
yKdsVFahYnHs3Tyqa7HJvXLVgR6X0bdpP3YoSv+bXt7759JtGikkDHTELs2cicUK
P77ZDDpkn2bW8O+/7gAL4C6Oz77UawgSj5HoIAd+bAU+QkcbvY8yARvG1be/cKEs
8lbVmSqj+1c0TCqvd9dfcz3BAxER1+C8m4IeGA27jUqsAfPRMJSkDsX1iMq6XXnY
fKQux5/xzXYRKuhgxnsYkzOu6ODpMnWe3wOAS+xLi2W7BDsaj84vs7VCvEXZroOr
S7cwif1oVcibeCvh+gzlVInOe1OK6eVdYBhqLRIkCr0D/XaykhHIvgoMooAKM5BF
fUtYNuuDj2O48JBl9Z0VdPBCtM9EUMXe3tE3+MH8aUxz1LA+6hPhEXFyWelUuceW
v07PgalVlr2yPC9cwpZ9RnyTscPWP7p3+j8LSpg/SEMTgVWcuU0MKLY3PG4S9//2
umg54SgAzO4N+FA6MxtmuEXiA5JV7SwcAMNV6IBXQLHdkZcGPW7XaGXdxPZbBGiM
DjGjoqLGZSpeGPkQXpEjMay6sYp1SzJTlSP0Bc5DwBTj+gC1vYp+gFJARQPz2vF/
uOSkWJ/O5neGh3Myt/suo762UjIdl6fYkO/lkNVpy7odk0CO/V6vIB3+IEo6zoPb
rDZtO1CELNLOFvDOQ1z1bORONISjXxmBivvWKvyaoveM0T/zUZb+mpnfPsWiZIbR
aQJ+Vw24RO7Jd4iPy5gyO9d6mNxMpUdiedrPgy1KXWr105f9jEmAh3SsRsAqPJsG
c2J4oUSaeoKpMr9t/CADNxFSbnLP1NhWwLxeigvCLLVDE5C4ic0kalWr1ecULgr2
cPePMg3SXWoC+cozrkz4sshYIFvuuqZ/zIKNO5oeFLkyZRHzONZ79Jevn425zak4
hrcgXXA2DG4hKZOeYVy777iVe/JNR+eZBLaEjE2RF1rk+tybtO9FKZmwYXdXPRgf
xA+drf57xjJPE9Mc0M6+EkaLnEOHhqow2xaKu5xeG980XUsDvF1HDHOjOEAXMltK
z+NOEz3DErOSIjGpoZ5epZyOhrFxSwv0IC6pBUFnwRS9FjsPhdBQLGR0ivsm8XES
r4JxUN82tU5R8qia+M1q4jIdehrERfDRyV6k6JB8Qxe3HuhA6ViNyeXCR++CqfDA
lOA2JpCVTeP9WwA3Wc+DVHRlhqwwEvZYXc4WvG/WLp1oE4UDp2ViJXh/4+ruyl70
r8cjZBhyw7L/4NpkTmbU3PfK/+WXF77cYoVFuQWkXXMhosLxtuGaEWU6Uqh7kR7U
U3RHK/viGrzwaLHiyEkFnpeSqJ3Pqr0/qxk049WGTJVqDXZQLXWuI7gxGrfiINcB
Qmd4kJNmILJZehBBYc9k4/6Mg1gGdbVcMcXRZxzZ4hO70QkeuE5I0uOJiiGVRhOm
1q8ZdA4fitRxOEfkPxt8nz6qnbm6XxkHge1zB4ueuwNVBiiUaLTIM7VY8NzO7QM7
KoHLbuGTTCYrnTGd5bqgF7pwuv8CMOBlsHvUivdFB61mpAzvAuXuLw8lFdpfJzgD
lgdWOyfBfTGnmpeCF5FTQ9C3CkBq/UZfbIsG4cORO2sqPhhQixelXuibwCCKCDYz
5bmdIZXQxeNrNcCJK/1tQWoF9mRa7uZy6MMz9S0rOiX5gmmJHkbHG+VqEEZaNnul
GOk245/ioLJ6lzyx31u4N5yPp3mcHygjYKcGTCoTE26c+Gw54bTyGyh299F2tFl8
1GJczAQQs52K/vKzHL0HZt9/uqqZgUyJi8t4h32KkjOANz8FKantwvoZ5EfldIui
Upw9MpHruGMvuZP/oanMi4iSMkfXcoNs9JeNQ5JzRtzv22YsEAeerOnzczL6LA57
B+1bVxn5Xlp4r92haw+0TTPOsb8YUe1UhbBpIPFS96N6fJ1lr6VzlcSkVnposObw
ZFtmxjz4KhioJiNKsVYooeP1cpXolctI+/WfC3/n0TJnCUMd7gGvvXMRF8LuSJB1
2OkAhK5yRsZTRsR/DIwVVYzwkTNo9hC88h41DTw4ii712WK5YzuECakZIOP/CccO
hTh1r6QKuESZPt6tkv7TbPUZiHdJjehBJdOjpmmzlXbpo0NJfbIpAhyl1aD+B+ds
sbPrNFCDBqyIIcTI4t6KeiOtTqyuQgBKUl1ppHv7LPuAd7qrqIghNDgG6qQLeJ9q
TRlcOU3QVRTQU1JAnGUU9Rrn5dvyjp0VzPMBdkcwkXAGV+BbITlMqmOOfwrl+Fdo
BRo07Tc2sCO+VA+phZE5hSzb5h8DjvWZlxzw938vPzThyBVKu1vj/8R5E1VPjJSQ
7oc437xsKdsMTj6GsNJMNKdTfI23klskPfs31hBRWaHclTJ5/Xt/EKA9VHfM6r/O
kjAWEssVjlQwWCiUQ8m1P3OavFwO6533tuadNY6MiftdywjVfTT1GKqI5iicrWYI
kkWIx9cTHI7M+yEqYEuc3sHEFzVWch732DpnRDx8snu9XQJRFQkUd6TIkZI0TWc9
luhjswWo5Pb3ZmBCQrnUHz7ebBAGuQMn/Ean0mDRprMGQRcAqMG79RDwWSaJqhl7
dOS6zDp952TDzOj0GHBBQritieUAnMHWIjAow9jACe2xKEagjJ0CA2ThF7JJAzHH
OBqYCG8i9MgcurRH9WbrNR7qyzkgl33HXcc7VW8isGxIOyBQb4T/GSGd6LtlqMaD
2/7LBDamd/fcvvPrFWQ8e1j+FibE/E2GuaacwmKIFHJzyEJi995oEWcOINu1TXlU
hUWnh27JDJnIJNgBpUCjkleNALKJBGgkn9vVHVuig9hIQ6rF7CMPWFUJ7zhkvG+H
TpdHUugIgt8UZY8oT4RgH1M8tSUbv7byy+eukRsrB/QeJsaIexMfwHwZnehfE78e
puSf+D+Cs184LmoKKYK6I4YzqLcfcRKeQ6dpvSTpGXf9CHstK/cNLmde+LUUG+e8
xqho88fFnrX8ps3shOPsOSYq1E2cqOGlP4CZ8okrAYKcSICy61/1bI4nI2GgFC3c
w3f/JaaPxy7kMkfTjzwpWA1/UHHL30ede2EWeKRW5a4BWBimwY3WvmotESGbZFcL
1YswGb1JX4nDV4+30YfffZ1h6GSXy9BvFOHpnscCWFnaJV9QzxiPaNInM5EL7YRX
mzE0+PRjNsp9/OfL6T4vXHHWOUxIc8a8r+5LU9ByiSy9Vs+yq80puWiETakbx4g8
gkKibITmXfJiZWuciPhJB6AuZIZaHP4UtJfjJNy+OAerx1baqi9EykfhjScliAK5
YbBkSaV6GAkYCQGcgJfiySv8igmjipHNaSAb81Exga/mqsySUbHseI5g0oG2s4Hn
25tzPAn73xDenmYrwdQWwCYb/im8TxK+KDnG9G5PxuxXIDUpWhfm+hpR3ZWDi5cG
60bgP/hp4k16FtoqpVmLNizjEb0GJZ1/T6ouLLgyQr1zEUXGDa8/clotqqW9Ft7E
+QvPEF5AasbqwlJP2+D4DP8ZOBt4TozeLev5yz8FZRV5ylYturI0r2eVR5064bJ6
KC5+xvT7XMPBOcdhOlqgZNxWIE+Ck8sEoE17wRUZHQ7u3N+OXIMsP6mDAzCOZlBf
K5deue6FnUfdCPoaW/dC7qOjxanga8AfmcDxs5xxnTLd2k2w3xaErbF0r0o4r40v
gV6cRISQXQPc05aX1ICAZZBLb2EB21RzTRDVELKhjs2j8oxGjUTHVWPyyS3x/Jx5
696oubRd/4PL3jIWt8III9z6NuFn7x7ZmzBpKT7ggcNFFHpLQht1GHVZ2w7TM8Hq
p8ivgzjvUfxGo6kIkso8MDdYjcBNXifk5+PDzACXqXpbc8YlCip1YF6hGtq9HGAW
CQMTFM4ODvnZP8GC+RAqyRr6YocaJQBqECSLd0upPJUoygn1fmVkOXE1/UDXfSlX
aQ+uv0PiQWMc02PfB5ycSccrHQmfRG9QIzTDPnb+VPr3aQKpTIbqYrC+9Jbdr7w6
DVlQaNtT9L1KEnz8DIQOJlk7vdfC9aYo15CozIC6kKWcARASF+ytA4zCEjEs+fs8
Sr1bCmJ9m4csFG/Rs/8/v7BCKFiNmu6nc0bAjudEmgx7OU0T85Ahv6TOluHZvdaa
4FQISFS4ibNzqNk04Zd2aCz19LrfXkBo86TrlatVx7JAzXisMsVqzE9wP1odGL+M
a+dMJAlDp7+FVOBNXNe4Zs3a4YvaZVQx55VkETDq66C0EKE62UfPdzXpgA9XFHEH
y0vvOeKFnjeeQqEn/akpa35IdAVvwe7yq7HZa7g892xZSeNv1Gk2A2zxCOkaQ8sr
xVskq3crWwwSa6I/EvKGDaREEd6WNt1ylx6n8oTtfal04ZvsAjx//b+i1JajS27U
zMdhPAofPwjGssgklvPAXFvGjGSwW57W1LdupYtrU+Vsqxm80ZcOJiWbKYNvha3K
bB/zxeqeasNOh2uWGpLStgrkjsVKURXZOhp6UCscInS1cDm4mr4Em4HFq+ZNMazm
iTaeqhudGkg5h4Ol4EewhQE5EXS1oGFlnnnSlHPat1z92IuHlRNiCexqZ+Ba5KIm
f6sxaLDeDpm3EYfJj2oQfEfiXyZFp5PH5mO+V2ubLNN9Rtaxy86dXCn9mZsnd4ue
gYxwutKUW7Zl7tXWGVihTfb62/D9reyVd09laIXXIQ6lrM2V0dBnTzLWCaf8SIyA
egEpLrHOv/62nFI3SnkgZl+Iro2OXxto6xIegCjmJoE19zYe9v01LpjNbCFE3BMR
D4oJa6gcoM78G6OUoUhMQVRqU7PSNdQI9e89PtO/99wxTeTCg1NGx4kCH1gwkE2F
yi2SxUpUZro6YmBjIA4f9TqBRdOs3M/D4cQjAG3JcMQ2ymtvmfdL+VzYJvoRiTsV
ivQtvp8C6UC+YQ0YfQA/Lt2jHgYA/eevhBawvXTK1l5nVjM++YM88JAecX8h5Qhc
jdYzdbXod6nRIWnFIxqC8/E+CJW/I7O3COEcDR7vJYx9OiGd8l/2wnpUZq0fgGtX
bUt6toNrZvC8TBJAcdtNiEBNrxQ3aH+p8eq0Xsb9AEyyMLVOi8JpqYvPw4hICQLP
IB/9Yo98nVyTj0fienMe4GBSGftBIjqCiJ7rai2izqBmZ4zJKKeoZ2U3SyO3Z7uQ
QVz0qOts4OyFa1AZLSE7KUTw0ngtfEABG/k1mdEtjdZ/uBR3/sHdmD8YZXm4QwDl
mi2+h8fxKgZKiciy5PsRm20KVgv+yfnl2ywxYv2O8O/bHUgDrgVFKYupnZtKwUIM
8TYqrLYC9GuQ1f35FH5JtLe8dNpmpltWX+mdX+opQa4C647vgDaeIjrKtcnOkHT/
qVP51IWtr21AakmNM2gjAGq32st5NEVb7KeNFNzx9ENeFyK1YdzmaWifAIHJc4sE
n9aiK6Vxld3YEyg9bam9ti4BYjewUL6V3r+/0J2BPEYbuzPlLFBKD4jqm4q00F3e
Whjc2foCQ+28NMYubwGHaouKSYFW2BvKbYEZkWOJi10BSBL3FGksxxrG/tQs0Flb
F+IblL4DC5rm+RfecGNthy9vBm/M8CggXIibNJ9c5Isc/lCunhdKdripQJzoz+g6
+qhqIlIAIGOruHJCKYZt6qcBf3nnR7PmoF7/U6rGnBBMcDP+yJg1FQK1MIu1OGly
Vk1ZuE0PZms4OGyHpDU72pvd9LIIpSusbq+5fzSMzG23hyHa7GD3ZCouQYiqPwHW
tf9UuvjGs3JRoFPxspBb8Scddh+RL3OJD+tiEbtyBgBn7L1uV33YgDPDCPZvprCv
dwnvSleA7OwUemP/rDys666X1W979jBuXF7xrEpAEtOSOo972S/sH3XowY/TqH0x
p4jw6RZ7V7+1nDHFU+ynYYXkn4VudaGAjENpAb4Vsqm3E2bHPCAqyCgU2HSU+vYw
5jK84Xs3lg9Ew7TT1SlJr2iSX0+TGLGVjuyVzDE/BNRbwlPKtSQQVUPXaKdP4r9k
rvPDh0ztzuHYUPifAfGH4/3UCM2PBA4F3y+IBBWmBu2cHCwUJuHElLCATcs5Lokz
aNL/vfzDzuJTnMg15OxoAIAZuNLjTV/FGTx9DaYRtduoB+9anGET8TZB4QpGCqNf
sTXL4aIHaGoEMjlVB+53htNv4+nCm/nG7Znkgw/jjWqfQuCbBrCWSzcCWsa5UgaO
RzSRWUK45moml7JFQDik/+B/ftPKlZAZtqDtejtQJXlpREBBC0G+kTLybtje6Ns9
6nF3DfFcIymqrWLqvcATbxtEx+m6KTHZHb7jGol6TI1hVoCHg7UW3T68G13AR5pl
f4FFR7nrEgMBF38YHStWaLQesUVlZQHdszjcMUmT19hQ+ZqogBrg2pueHkHOCJIP
NhmioJwymqncMfKd0KsZBLiI8Mh6bsAW53Uy362lElNlad1CGmBksU1TfdjRthqX
hLzMtIIE0EYxxxLjVyqryjsr+m9knE5u7RLTQuM/HsAel74Kvfd84/p4pnA77Gjr
IrUE1tl4sS3TGGN8jQDPpf5PeEAu1iDBKARSNZWQF7yq5VnmwLTjDFJ8dKOXEZXg
V3C0ZjW1WI/7h26AFeYxtCrLG5POWoQzuCKAILPIZGPyHzvhLHJLJD6+QEULRPzI
yHDXKdIqUcFIfnm082Ui/zHSxnyTtQf02sp5mc6uTiAaWyDCVHtpEbGJHmwR3D8D
sxO9tKqvDp+9yUi5EyhzbB93P00AhkbtCG/N0cUHCDJM+V1nxsdWJNuHLPubrzZX
3tpUgqKeznwpAEeYTZT8qgt7n3WgmGHS9mlGUw2rd/FHLMfJfg4I+Et+vXiXQuaP
bPnzMtvzsrNdboyKEiQGDjT1cypY6MGWjBTdUb8gJyMBtZzRJJW7tU9rzlqwtr3C
D+a4mFHkdeACOxw3zTQ0lRnzoZUl9jTzfy9KY9xqJlKPTYcmel/HG1X5uCq1aQqN
a5Izt1wx9kquo20tcjP7SED57RsvSC3ACkZL9etZUQ9f8KaE8tVdTv/WF0AbTazU
Qp8Bjd3zKiauU1rRliMexb1Fg2h3RFvZnFnCEWPjwNk4X6jTW5IfvCVa9XRk9J9E
Aidz0ue1CVyiUB2SSmoi6xIkCZ2BiRF0bTxsVpOXHRx3qD7zjpaXeTNo1JGCeehc
GeIBVyg2Goe2gdthyt0+AcFpaV0t7BLnFEv0Sq/dQVu8Ml/ZjNggvx2QHgLC9vvG
9PEavZUKfPlGsG8byqQLoz13jHdRoeaLMQHm5aXjPmIXE1ku5zphDjbm5/c7vbn0
vcJXcGAalmhA9d22kDe+E212QXw4nWKgju00Ct9lRsqoFLsKqsPIl143ML6zscsh
XdFydC+p7o+I13yzsfR47tTWB3xSPKD1V0k2M0xm6lLTrNX8i5k84H5TOdZx9q1m
hPkI2996+anuQn238iz7PZU9ziR0qVU6Sgf/ezMb55jjpv12VFpvcz7QS+op6SMc
nFBPx4MMSWtj8GReOHiozawoS7JTvzvPQHKx9SRW+MBfStFcT43Ktf56Krrdvg6o
0C++apSNzikwvglFILkgsQLjeGPbqfZJTXddjSqMqjJ/SWCxwRO+7wQBbrqt46PL
Meyq5P3ufZ57boyNwomPs/h9c5Js7c+zhOD+XwWX/XmI9xcPE2IybPQk+MyZ/1xU
yQiOX6QBH0R5//frwalVGkFcBm7kwrOJwK/qr6mjPQvSeFA5OCn7zTDAq8WPcWpW
IUiccL1i80sJ5CvEkj3yFRgYQHklukxqUM7lBOadWSZ6KHSSzyHzVwi6UfNCNcZO
VMRgDprzpJPSOdVOjirbNi+gGW6QuBMwnDIfoStrjtftSBpwOcFisyKVoLBKwZl6
fgtvu3tnSvMhGqKgW3PxJ06FSKFq+5kvSAdwqve+GT5byc8RhSqz8Hx2LRlQimTB
Tzv9FTkq+snD64PSmX72V4PSJMkCN2l1XwZbqs+D3jEoVaXzVRGj32rA9DEHwH6p
efDw59LCB+alR8O4alSSi1tAC3MXNvSz322KIZK1DDrr0GNT0LfH7jDfsQvhzoZE
i5mYQ2z3VegQW53jSP7tQGl0siZQWTWM28xj9waJBij7/FQrigO6FBXaRSZRC11N
kpUrFhzG+kuzgvyIxE/1Iek5BsWPM1uU6t4MALgAw8Smdj7R62kt4EZAhW7vSk+x
HYku5nAwgGBKZsteRpi5l11Navt1gMK4TNwzx14V0Y3o4Lg1XpINMdt/He071YdW
Iw9vQXFekqXtspj9zk7d3fAShJEmi6ycB3Nis1quvYnOf8qAK7WI8THXelzihlUI
lXe2Gm0/t3nPFQfz7N4VOCfFaCfHvwow3NdGK5bv7o2roWg9c6ZX41cETGcdUQ3+
r/cr9CxL3YTTtIOP6itnnX4SoB30Q6kZcUVjgYDADIE4T0nMmNKgi28WQfi2eMr8
IlHXHh3mfONW8VaA/u/+qVTGimvuHu/GCul2m+qSuMpl5377FiRIbHmpPxZV+KAH
Cl5wEy/WFueOxq9ktuL5JcaS1QD9+Af12/3kMw+cmws7PXcax9ii3UtysmLoKp9U
y7gJqlqWJ6987Qf9AsZe5dEMHv+15u61vkOP5fy43fn9/JdpimxOF+0pFuFjx6Z0
BVpQqqjG32/tF6plU7sL2K8jiocYa6IDlQBI9WcCwHImseM7c/3sube1jBr7ObpB
+s+R17xbOJOruN6yglGVdvbRhNTocgSueXE9BwgXH8h635LAyW4QkhTCkD3rwfhh
wtFeidQQH3Gcf/tE7YVAppRkkUTTESPrPXOpgbKvP5InMR6556iB8OyWcOedKrrX
xqlaUEb0sqqlJM+a5306J6SVpexbA6faajf02T6g7LcRy8AYCcuDH92CD5xN05aY
hOPa+9vcdWkGUdZKvcjmFrv9aQGqsKkrhewynMgl1kmwJmQFyp6eN3IKhD02YIiZ
9S6b4ytek3CT25kDj6e1MNaL6S04P3eaUGJxlnSKKn0uJ5VyFgh07dCWxLCZA3Ox
1KfUBucb42z/rjo9sHyBdg/+0+6MSEvODCWKDFH2v8U81r1V6MwoJxGyMEXwbg9B
1NdIRIQTkPFSFcB2vpeLDxUenFqxyE86DnH0IlFDccjcg9PXRT6UF+JTs0CazZAZ
8VVGgxoj9KVfXsy9tNu5dlOvMmczHBkakfz1gAkiQ13IeV6G3CrFly/r3rd8g65G
xNMc/iHPiqYPKAjocYyU1NxR8++lztDMLDVTxvTlZ/nRKDtwY30fGXLzpZ9ipaDC
KjbvopWaWiNIg1DNH46tFRn5dnsyZKlM3pz85FnrhrZiEHSofbF0YDoave5D5QGP
zmpuF+tirihJqp8fvsr/k2ib3A59yM0domQdYO7J27KoynzoRvS82kQEWG9zSkv/
QlLfPI1pMaauT5wQfQV44UP+WMNyjbvyoNJx6URg70BTTip8186JdOVAl3RvBWQD
bqS1nuoTJ6znU30DB25ooXzpiQqy2jIEtUAOeYKxAkKFI4Rle9xQwix/sQTqOWm8
6CnBKh5OpM44aBH1Nsfh12QpI5g3EnQgVdF2h65ZilCSuHD9/aRITjsnzMLpisMa
eF4QXZMz1GRtjhtjkFw+Wakf7JSM/tPC+LdKNKUpe9ontf/6Xs3QkzL4O7ohYhrO
AfwkFWm89jVp0HuoR4xP17mV3ITYEfMEEIJsunViOZA39f/Ohy+I2MEmyFJkqIjb
8kafh9heOtp12X0ycQcItYgxlYssHS+rpQsDpe2vtjilK6KB17gK371+oOm3CAVA
fsQzTh5Ob5SOwCHPg+nrLsncEZzYyydxoGKnjb1vAiciewV9CpDnp1HjEqjl8UYZ
mt94SW4ULzm8ZD3F5bujiWAKy3XiNVqV74q1cB00ShVwFMDdAG2jq8zubTqxZk9+
K+fzL/pAhEsD4XLJDknBUo5qS7ETEuP0FlZOWIItXJlAYt+3OWheiUqgkrF3c+4I
ljETbAD7yNepVDFGqtJsc/10MaQkBZBw/fFdfQrZH/0FOawHgW1hDTKNUcukuT3g
y89KIS40+UZAMDZLAG0EK2ySpZ7Gxzz0BgeIDRGP5IKiGRVW/2vhOgH6Yh3C6hxx
qbq5q4INYbmLgVonpdlbGG51B9ckOmtQhILJJGTQyA3a46i9UdJ9DP7xoY/HsUK+
Tt19VJbjp76ciCwbsKRAiB055gxIdjPLlMQLH5vh/phEZubFD/klyBYU5GZpfLH/
r8jMnqQMR2K1lE8BLmd6LNJnSplTwYsdRywP06CXvkGC1bI+5iqHR1eekpnwYCC+
fwOXOOhoX2kpi49rH9ZyM1rlFtPhrFblNsffDeIpPCu0ezX1aLbOUrtIYT8tfUhM
Cp8iWNhwqQRGDwuSAlVQfOlHLkrgE/7H0sLf+AsOaNfzLFyicRAuSCzfanf+dPoq
CKpN0r09pPCLKRgQQv1MqmnFmImrmxruvZ0WK7A3cY/ij3UI+ONkdwBSIIjV+eZX
GpfR3WgY06hYw4OMEtX0R5I3i8BKrpXu1erR9AJhFOH6huxQEP7b0aAMvNiptP4Y
DVaAN8NyF/0IYpfiP1U9DFBnZ2Fpp+Cmz62wdh2JaWOHYeXKzTCO5eaVjE1aTfYi
vYajejq8iY98wbp/C4j+yc0GQROgDHARbomYh90EPhiZzTluTUGET8JhjA+dXkrD
NDANT3eyRzJE4zesDeAhQw5jZD5hJz7I4rz+/QUAS9iv5IPAtEVN/A0T088wMz6U
MlvxH/GqV/Cj9+zuYwaORiYAUrq1s0EL8IOAHCWfq0pGDDazXoyyRmSnGHkXjGQM
bONmNsxxblKq/LELuqQWH7qd3VdHta2EA9Shnrk/AXzyNFZJxS6SSNRtT/cjNjy+
Pi+V+pNrslfSzgn39SS2fb7XIIlqDh5RNfS35Cr8l4vYEQlNeDpOS//K+sVyW0li
jlLz296N33PmQ7XBjptzgNNvocAmYKijmRmGeTSy9HiwT7/jN3uRJdXqWrc+KRxS
5X4v2TVT/CA8jcytqRR0EUpjac0tzlCvLtzdTOTmKiSJ8vZyoOKFWKKT2BTjOiIv
qKgJUlyp5RxJZxG7TSRXQirVzOrEEFa4++PucfvPJEmg49qp8ZrjdYV8tP+uHy33
W8S+cVtZA3Pjj9KEpFmR7P5petBXBDYQfLG4DUtFqsNKrDttiW4Uy4RJ9XyLJwrj
Hq1H50RM5doIRH2mdmnjM4GFJye0uwiMpLSxxUwxfjTAn0b4Rm0S5QnE6ohWlqIF
wqbnUdo6fLaFbVOJbvkbsHKPSSi345RvNR2of9m5y8r6chsoycjTPn4nQGdqULpq
8Fb+0AZpRlrzSQSTOlEhTmgm4DmFWQ+6IWYBZPPe8wBc8htoHZT11pmpCInlTdbn
pVXPFQZJHPvlKIYbd56oH7zGyjN1RYl4Hb1KrAK5aHnuGn8APjOJ8xD310bJPRP3
pebf4XaQ8wmR17dc+Kjq0/3JbFJXJyFRzXlFVc6+pUuuFh04WzHBqtMs+xKVvQQy
AG2z+SgyTSq0ZDTijgxWktTaKxBBlR/Y3xMlIcRO1TRXXmRUrSx5WoQFIobkfrRA
+m6Usxx5poCFug0jiyGo0CWUg/K7u8b1HDdjMDvK3zB3LJ2Coi4FJVrgifJxtmEi
0TAunFvQj96MOd4jnsIo9Hz5uDdh3d3xl9v54MCaBvGt6HkSWxatWyo8et2fsbn7
I/2zpv4gdwtUQhz7jDo17fK52nfX2ZRGR20V5TF5ygfQ+TQe/vDPjwnZMv7NbbO+
sIvLTnUk0OcU4KqTNuHQ5C4aeKJx2a6FElWDaEo4MbNG60y4+Tma846nvirOZrKJ
QbN2s018w2engXdCyshrFxITlbOKM26RmxTQgT8h1szgzOy1MNiJZ7Bww2Wckulp
Wfr2fKDjjzOMkk+edydvSeQ8tN5QEF/yCOORBMSAXgD61CwKvvSz/ryvBaprypiJ
7lWwN0YalrnQ1IETpTuVbwdaZpTIYxJ09hFr37CMIUpf3rOpWJnrWPkplWtixjRw
QXOZ8hnQBZqjx51a5VbNBInvJej3jzRoOw3qMDEIk1JGuytVur+rSAfBNauxo0+4
t7d4/K502HRAHEA9bsqBOn0pj2npH9mav9Fl7vU99GEb7l+qq62iyLSUZJuga2Nl
U/IUKAGRPidsJ3XRq9ViC9lz4xTvZYvBD31dcEzd4Rq6vl6U0jiFbHiGWvKXWxrd
In0lj5VzEb2/+BSvFpoy4+DYNU1k6dB3xIyVvzoF5otfvLuH8mbj9SKMGh0mOPjm
YggNs33r/jXtmk7fiBA8i5gu0/qDR7c//2gm8sPptm70/qCtXMvIatvOe1Nw0uua
hnHOMAruey7GwkPhEsd+dK8Hh8ln9WsWjwBGrrGuNayXx+jbiY8+D1Ruq74m6KnD
hgoyWAMxBAtMSZ+02nR/oA5MZ/UMlHMNxSGMzWenoUYHoXaT/asfJdELRqhIiCSG
qDWIOB/T0TlKAY/sQEPktFo4DfseOxKIPWjgLUkhRMULcQE4rdmTTAHbD+BoQGNI
zE+y1U2v2RripDJGLRqpybPuPx02JjWsUXAL3bUfLtzlnsm7z4an0DBzQtdi7iyQ
pX+ekU3dSmLVcyPEFspTzIcxL5WUG4cyasteXr1TG5SExYERt2Ylqora7mn13rEW
JRpVHIYNV/9nxlkgRdeTIZv3NULeCiMBNEE1P/3oM9GNJt77RE6dEtQ7xALn2A2v
c0dQubPmpSlzPDcN8AJ3wATbV3oH6YeZOdxzaz6SuYxJTg/NbsTwcCS2vMESivvr
FhiY2HnBqr/UoPLvkdSmWgNMcySvKRcMdxMOdfZFkX1iCtmrYNISatwxARk5T5le
rvl8r3mvrlA1scd7UKpz9a/GmGnTTMk6qwMKM49WAp7KQEdBiDcEMGaFcx3a7i9R
yhH9MPsTNMi7lpBD+5yLm9J0kcupTvh6brgI40BNCRSfP1f6xISwfkzninh9nqF/
seC5R3r+nOdSUAEajZDaVfor3AQi+BBDZGiBDhROgx9J2Y2ydGVsRlXgiy2rNMcm
FzWQLo983Uz8p4298s2Aa7438lhRwbzppq+xRiEV0iu3ubVT9hAHjtx148eqco1Z
KYeRmQu4gDkRrpbDlqZyQe4jLrE/W0nluu6afYjhFSsQiwzzxb3jq6U06jcq0Qyd
8EYbSkj0aD53mrlIOsfQrc0F2ggwrUVVW+IhxglnhPegnHxU50EbxqBAbZ26Uypq
DBXKZHkABf95edvRGpNxSY0a0TsU90gxjmczY9sTONkUcIXq9m0IikWPam0vVN0b
M4IXNS6nGX6SlgIJqA55qmQiY5G0PEihzRGGT5/+AV7T6vnXK40J+DkrsX7bmBkN
Q4BBOhpnOEpTb4XTzoO4ckILlFYKJG87HhA0chiE1jcj97P6JOk93gNq4a+9IhVK
oLgh+rZXtYP7dVT5YXvZINjzH1lo1Ynw0wynkdUlf+IRtMWgDza8nM0OLnUAIvn6
AySA+UP7SGgWpfikgZqdhJFMGKDbD2ICRJckx5g6100q+YsAVTrMfv7mPoEudT8Q
mdvZ+rY0IPqFfKR0hlWm6VvTEWa+Gh6ZMyxAGASVNLHEED/FIA2Qt26NvtLWE5h2
EL7u1Tbg81TGhvbq+LK84eR4hnySfkwiR34pHDbrw3QKYgIrawS4qWe62qQ64RmF
wLAQyRvXl2XD8zXniYaW9FGE/CCIHySkGM8T2cH+Rp1HMMCdecP8U06xzwvZaHwg
aRXZ7UpxPeA8xlfeFpJJPvKpmsF2a4rDm7EH7u0FDcJgK9SPQnioet29oYQwxgDV
p31lOb+6iIvGYbZc/ask+qHp0iPfUV4wA/+7YUw+E38bTc2xGnB90G3cTuZc5jSS
hSZDA+3K+m2yp/5Kr4w5JUUs3on12j+zLVvLmPeJG6XIlact9Gk5HjDJiZEUtTTT
lZFgtnnAawkyhfwiywGPMMagb3IujA4mkpZdgBu2OfmtnXgSMiEyb1pSA1h2EiLr
TgJ0aAr0oc1r0pnZzW+dUKXIGBHHfLjoafYpotfXpFywPqq1YzbAljp1qankvO/3
HpALfRIJFI8sWeg7Wlwqe3fHnxiLWgNEPX+JkU8Shgq9yKR8l6bjLXrLnnxqikdO
2l7ZzkXaoHU6Z9ZBho4hCiGOTELMb3ijCseY84A5OEfdee+Jn3QTr6fH88zF4GiV
Vv6Um4UqwJGxl6AHv3lm8DEj+Ye0QYqrOMwLDgpcSJ3r43ATkqMBWlH993y8yToQ
RRgflGj6GU5YuvgRXRfEcgKsJe5ot60obllpH3avGSu1fZM39T/yt+wgxEh9c/MI
Hrx12jvIALyrez2F3q8qXQ82QwkcEQlbNpUNZnfmO7HJC6aa/ssiYK1j9Skbj0Ae
dpmEycxs3U8lCkO347wtC6nCZ0aQqNawBIxC+R3muQe8N+NPWXjLHTYvU4h/yV0L
yJ8XIsHzxvH2V1P3/jjjZkXyFoIQ0gqhgVGrraXuhEXREDafhr8/JP5c3D4isk3R
aFbBe0Nri+5v9Tt5ywWIngGHqlJFCLWot/0HaltFwN5N8tg8lhAqEIVjShUYPCwi
cEzriT4tW0jwAzmQEOhTXYNCZaAjC7qzAnU32NxMsnUQlbzZuRscK6BC0CZjgjjR
r2vtAJr3/+iG5h8iy+gUvcPM94o2LgvR/ZPaG/uNgiypZ/33CDeTr4IIqp94sh2Z
m1009zIgsrEWBAK2w6XVGnClkD/UGiMCe0ICZE1tErijpjpbcGmM69VJ7W5/CCZh
bHRyKXog7BsteQG77D1Kf/fmdvYpcEiGMCLybVkGw0ULp/Zzx5qUzzuh1wbt4rSG
fxG84Sl7Zfx9w8/RH8JLsDBHHlP3248Gz1/dncVWJYIHGf4UWwgk/zVi/Ebn30KO
kFKoxwgN5HmSLH2cla9Rfhil6sky2YiF1S8zh46gHWLh05wtZXs0F5kBqSBppuBp
mzYiDgBXEBuDc5/G1iveYinFjC201GeKAcUiKwnp+sCfMjdP/LwEPZoE9bsXdTC7
x6iNoGEujkKjua4jHHb7ssRVIppAqbzeCiqrrVOtYBzDweeQHMG4WigtWYHGcmQx
kdShEslMjUGKYTloEivjdmvnkdXGutGPyz6S2/PL5Mguz8/aKAR7vT8JJm8k0VtA
gZM3Zq5MHnNYw/hRTnmWWdQ+uzciyxlrnDmw3zUuGPJZKL73hne9KutySTH9jjcj
X6JAMv9TR3xAz2XZdjtC3kWN3UjO3mM8u6UW2b0Gz+wI+++i1J8apoLBuvyn04Tw
pcii6hqTOzTjfQPKFT9D9WwXOuP4BIix6vf+i6lMTEikP1I/xaLVWGtDPs4+FYXk
LF7s16VJm77uQDSJdF6HuFB4Xz2ykPyemVLexm1bqlAD7jetaP6F2RT9RgihZMy3
SoAIu7SYZI3TWucpBspQuB4G9EEuVtjvCFyRBuH4n3wT41TFxrUXkAgQciVxhP8t
cpVIMlAA+eqHNiIeUz5qXuHQ0yzF7hKgbTwD/OuIRIZQh70eu+gTulNBfUpK1bHO
ANUxQYFjKU9lQzysAHS+3KNYtbL/Y3d+Cu1oXL2OysjQspF5DsX/9S+mzIvTGzeQ
P6MNLc/+UwxDs94B/PQ6FNjbwAnRNyTOKLwdBQKHZzvyLgqFhFbigCDE5R9ffBhm
rc9YdXyXsX11KPK0Ek4nGkde9D1FNliHao1pGcMbBtebBBx52SLgmu5KZl0doLJr
Qv7DCfyKtHidPIyDaIcylb332nq2JYRh6bHJx6IN0mogdCwLosQDs+bwy6uPI/Ns
ZpG68/NpFq4qq59unj338v4XDlyKko6ISmKukTZvP483h08FiLL7+O2haSipAyqE
FASv8qv5yPl4jiQzUz5hFLMcpVIvhaH2NUPMdvoCMZEs7zk3dmKl8z2nhKmU+jZA
Osgw23coyevx8HAp/le8w/3cgniVjHUnUFsLwlfOP10ZqF6q18HcogERDCr7NArV
Iazi2MfLyYBqlrAQFaOsNJlSyxsA12u6aO3Wttkt1RaFHIDhqpnc9o+iQMBsK/rN
bNCbXQvDuvtACsx3a+tHqWeRrxTou2/I4lb7GXbrICDw9MEoqSxBv5eEshs0y1Uo
N+Ltb/zMHez7hkWkWeW7VBBaKDFnyICTET1XyFFP3iKlCzBR5XtBchae2NujSDPC
roee71wiXU6FAIJiswfYgfTRxnn7h7Umh6ekJDVvzl43qPiKJhhA9XdT8Ys5qZjj
JNP8Jbzuj6GpA0dlfVMfbIj2+MQeOTkLpe2/2wxGLZaAfEOtXHQe30nHPFw/QZcN
bIu6wYb1FMm5rcbvwjPPCwSRFIcexSMgxmILKPG0HJAGQqGW9/ayJGvjRCHQkO4+
d21Kqxm6b6HvOH/n45ME89FjC0EMEiZ+Pg/eQMbTXwzwuM3GxNjlVMg4t7tufzdN
J94K5+3d0gCFC7bNMvueEfB2lqQuzkykeEiNs62VnjPDveoTlsn9Zumosk32KkbT
miS8O+u37eQVBXdnqy73nFP2gm4etZc5AtXd4yiLxNTVdGJmIfqzQs9mDkYpV/9x
mU/8eQmxdO8sSynidHGp0KS9ubFFyHTDS+7zLkVtEjeIhOZPppSdYgoqGkAFY5u0
sPGGNwngpv+ZC4u1Ts/uZc2m881qF4TMr3lDoqp4M4RK+zpFWKz/I4f2Z674AZPJ
9/ZfVVcSoQVrjJdnhuNVG3OLanNjhwUw99gBOGwZ/hvoABa8NEzQe2IbrBJUIoWy
6osKhjuHY+wdyKh0Pfbw/Yo95lRFPiMb+35/sGOZNptWBM6FdXTMLKFYKzkLn2Gy
t7m1PQrGV8dw/pQU63ppvcyPhw2mBElsiRAdfnC661Rd6SY6gwyw100ct0Gfvu+6
OvmvIXK1bEHfmrL95Z5T5Q/0GtNIGs/P4Ge9Fqzke+utL7AY4IB8/yt8yqP2wZO7
sTC55AB/o0q+Ef/UA0urKJAJvV642GvedZCfRxVqlkzXDN9xmZfJUfmlLqa4vnf3
BPlk/7e6T90U+ILEJfX/8EV8+p+LR7efC0+M2m3BCTsCbr/P61c1/k7eF2xLNlle
9/kGihDL6x7OYGjQooOABVORVxzQczjmw65+sYzu1XKc5SwljhHxcp/WxnbkUVcJ
p95gqAi8OQvRkrzfjnWlLcBwNI+yq1AewEnETUTRU+LjdIZgCUdgJYr7zNd7sFHM
zn3mtE1IGt+zbWgrBgjt2EbJy+P1wGexH3v0ydnXYeS8a2dJNi6BIFxoI4ZI8RsU
TiYMx7iKWfqfS2XBlenM/nSLFcw6mvEiZGF+ANGcJiyGQXmwhPJ0AAq1+9EdyRT7
UutMxEF+O+XpLlraKNnkOmBuXwZrDi5UbKJkPYB1Znh4ifFM6CDvm5JW0g0tY0nD
hlOojdABk5EcgiI5gpanHkNZ/XVWwouH0qzcv4EQUTZMrcFF9DaX/F+NGrZIJwDo
EfLMfli1d22rSbMitHf/9BFUiNtSCATCplG3yQ/AADojlk+tVljSZ2x9uPEuNa9m
ln0OFQIkyBa4kYH67/FtOwHYdLuxfsL30V1ryf+7ujN/5gFaj/3oRF/S/VAvh/XT
KuzT/E7zjc/hLHtc9PsKTekU+uEjwhWptXEnuvu5q0/uIaeb+XNMZQMmk1DKHa3+
GneVexjhW6RDcr4THeeLsy3E9MET94Ujdd7M0IevTda1X44pzjvT+7VNickj8ZaJ
HXMWiGoQdbTQedOsjpgnZ0+2BXhFtflkaI3setwcxe3R5VtKvnDZgGylzEdWFHTg
RKguY37jiLSkrOUO19MiM10io4mgaJ63vRkRrSrzXIfE/8FVgWuWDO7Y4apnxP+0
BNALjtSOi5RApdRMoIZWu3/9+1j6ktnavg+fgtOxyWq2jEtTf2EgWtyONlA33rKH
lyxPOEHGLFEKoei8RbQXUJzkYU4X7Ucv0IgJu1BgS/YBa80f+GGrcualUHNZpJLo
kBY+Zs4Q4/mJTtN/7SdXJsZlWo6K7ltTdlksb9evXLs8hRIuVndRsfdj2TGnaw0F
kR8+eg0Y4lSOgC0WehGvNq+SE2Q24bxhncBlIV1i2ngayFlQ0bKhYOroybmBlLIw
E2CQrC0hoaBDi7dXq9KWS9zsqYbbJ99Tj4eXtaq06vShBUMKFmOZsC8IxBVADhzv
DH7FL+TjNBJ4kJox1UwojNLv21TOFgLIKOTZz8f67Qs7cS/KtzcFmdz//IaBsUHd
vRuPh8FTiPwpnUoaiFpOgzqMPmdqw3/0liapejd4c4bISauZ/kjxxYi2GOAtKhrh
q6QWrE4Irpu22m2awUm5XqHJSTCMHk89rRMlgvyK+gAvh963EHkKtAfYVMt4O5NO
c+wKGQ3zQTduXMc4zqbdmAQbKR2LbUi1qKZVcJ6xPjXlhWm8wE4lD6kKrXgp8KRE
O8V2VUTVgx+d6RcRbfcAQ6PDMmNxGP/q9NBe3ii4J7i8hOqumjYsHSF3zLvU4VzF
+z03UrPhPJJJiocnLU2UZ9i/e8ccZQLRSk5jskuBJjNLjyM7jG2+f45xDQ8/cb+Z
k8a3x0Kc9ZwYaAFA3tuzF8Vk363WS3SJ51RBHZLOSf/gwYlNzEgYb9jcgD8zYZ7y
b/xYXrcBZj90dAINCbthULqhgW84yXEp5at77wF3klEnKLlxgbzi+4y6MFdzxT+n
udmQ294MDQ0PPiYUungD5tkwoM7mDKpjDDOFD2cuxIpNleKGo3WDU+gzlloTa3fY
c0n3hUmHemyv3HMrFxKH2ag8gi7Mckc1YNHLttzj9xMMu1QEgTiOEb8Owpzg5RjT
i28tPRsS6ixzLOMZzK94fJMwV/5yjp4G5MdDlx7HP2iajMBR0wu1IP1MYt/426ua
JRjgl8Mf4UH2VnkORf5az/O0dRYnAxmn3Wq91+CacsU7WOkEnSOmsAgncVEEgHT/
+Z3mvSSJQ9agqpl76M2YAVv9T5DJDGIiCRmphrcGEkKR+Bq3UpQAgsPc6kYSxzL3
kA/qjNR+Rsr9I9+JlbWYkYm9Zypt+ewG8umCWJ6abVFK4XfWw7ZfE1ZXI99dBI2E
Icpj411CPbj3OknuJACWl3iTtMznaT0IPuGNdICd8gms/mvdRdwPSKBjtCEVo0js
k+7fOumBRCMaPPEbPFC/mGxuMYti0vzaZxFJbbv1XJT3j/OwojjXUOEPFlFMjdhX
Sa224HLkgHOgGLrOweFE7pq//5GdHTGhBrjGBPIxuQvn5NzUeeaT/GuVsqxqhm5D
YFvJECJHXvq1EeJla+fKkwCVnmQG9UtYYPEYharzrJQ8AkfYpLRsIlU3ut/1To5f
/ccwkyFsZkNrXlvKlS2vXAq2K5CzfiinUkNezPhIghC1YsO00Loq9tKR28Gny7TA
2UhmikqU6ANSH+h3gf4/C0HERsUyrCG9qtgzQAspcDX9uhtrfX5a1CxqUZa+qF1Z
1gJyzkKYs3OLYup98HjbmYCJ0Fz+eqUWnf9spE7WqgehLuXQC39DgB8iL7jqZQk8
fbHi/thHfqGkVsbGP581+J+E42t2LZUvLoFmjwoeAPOvsN9mfWRkvH9N43/1otwp
lJx1W0ghXPjmPOv1/+vdeYkI+JkG51jepLq0IXF6rLAEjpTrqJBtrm9O3AeJrKZx
Ed4f+y2zv+BZyV+KGLFcfmZqxadCXggoc1VX186/QRHItRmD3mLqjVOLJqt6t8ML
2pCkWRvQ6y2OY+Ow9kcKnUBhNNs4zF4Q4cF9faRWEBQ+DzwfLK17GvPAN+ClhESg
3ksQKMCGVilZKliLX1U84TZiKLF2eH6gdJVc0Jc9Rw9+la3j37EjGDBzg6wpwJDA
bZm2iP8FsU45v72TY4hVGbnd7Iks2NHO50YieVzHMRsHySKu2Ng592JfyxKLLWC7
UdiyjZlbISuGXWn4Vi+fqAX8V1HyXDlmB3ERWAVGxfipGS3BrnDBYFGgRz6jQXu2
0gi+CaRQt3sVSBfd/iSS48yxl8H9ciwLRHsE84KHvgJCZJeBR15/fsvzgGdLBLx+
AHl0PIdVPztw5ndybjtirt+AIYnehy/HNpFCYem7oflO0010hv76vHi0xCUZ90ft
2wwzaC6l2fQRVbeqK93xnbI+jsDMs+hjDSlVsizJR2D6RCP90fU6GrYmwwSyup9M
Tamw6T8gJFYmjXu7qXRLaVPjO/CXiiJQGQGy3U8ysOMn2hYCpN1lpEhqI9N/QEr2
REwdVh+hIFMh8fWLT0bd+3G3WCI2Qa5L0o6pbyfQcAg+C9g4o2N8o2zlglEnlC+S
k4COIEtlASW895BKysjR38DhpTYvAyvXx9sXcTdSv7ZTtSOc5FFn+wvylFx7oWj9
I6W67whh1uVVNief1CORfV8G5jcwarngLpQHXtvZirZNi7ot54JJ9xLh/YT/wmVa
lSXPT+v8/LfRXuA++/6AgFiKfZWstrLSKAl+lGM4OP5rAc9yXz7VmBzrFz+JEVyU
RzX3KWMWY54OrNuvpyja08H7ri5MdKZfOGWUxu3bCv5snkCTOs9EUF70pyigOjuq
xPb0qhbD0qk86LQ0IEmk40VYZa3qIuk35qItWmyMTO6wOuww8WJaPhNnNKPDducC
SrkqtmaHDQ7cX0FVyClMHOOx6wI7av4yuYTpvq0Wg/FvGo1mLybeFXMhRn8HxSYj
YvQu1W9R1gfmKulAC2GR61BMrM6kLiIZ6FlCxK9gTPzjtQDF08k9qfOxVFuL1WU1
g3muvKiDt+brIJ9zFCML8X5FF6ZsEpcPv25W6ZUTMhCdaUPrf0AdKXdOMyb1dNPm
D4AshQOrGUzbU/9cFEK9P7I2PN/R2zVcUywSgt1MEUGqS+h90pwgeWQVjPq5VhhM
5ckhsyleIIrNi541UWQ14HDfhMKsopi8lcTOlQfotg8qYKmODLy9k7X+l/gCp6vW
UIiwPIB7wQBQAZE6d+R+BxEb+blGJboMPStsyASr5ZBdJ5Ja0D0wTZuq3HWPBusZ
btk8o7739xpDc+EYXAFLnHuvMnDkLVcuJpvaCwXPSx6oqSbhpA7CYg/e+FYouJIY
kNg7k/VYOkKBiQNSb1V0g4OzryMEqdabx8R0u+at/oH2ux28O4/C9SxkxOVRPEY9
r8eVYVuHT+mozR6bXHaV8YfyRfuYtiJa4R+rlg8yK4WK9qi7w8B3myZ0n6GydvEM
vMjqyDIkzSA4TEeKo+nDRupYpZ2xem6JZ5ruybpzT9UgyQ9S9+W0FbRGzhpTkP4I
sROtW950DdACfoecDgkqp58kmvfx41RZ42UXdW6sQs3IwzbPUqrhAhDSq6HuLncp
fL93s6IztpKp2yY4btdIzknOHuj1tlC6we5mmdZ7OIuKeXypZRaAAB7VjF54/Sfw
QyUljGK+C9HBoVsrQm893t8ygbr4FMWR6cZ1S57RpKk5eI0mtej/S6uFwL19QJug
wDL1Pe41dkBKC2eB+Djo0AJzIVOR5jMSDjOWiXtVbwhJzlrho4/3Wq+4dyL1za1F
z5D3uy3Q1JXuQqN2+7tPMgWj8m78FfdhodqsZOqwc97zAwcUYk0IIQfkVeSpTTFs
mYJSZxiC3A9RsO7m0j1tlQDFkf9HZtI6JyJ1dDwEr8BMJgK4Skm3ytjUyYMUBywY
ubMJbXuNYedtKGUMDBdkb/ltSHjIhZLQfteaVHM3cn2kW5xxn2SW8OqLqW3BGz7C
1JI0VS+lIuwpQywamMCClJRy7mfoARnbiYd6w2IhZ9OGq8tuokCdruZG+EQCjD8A
0p8e/3n25PPVB64xZG8qgKFhzoh/nkyLzynMmo2xUTU4G8mcz9V0Sq0qGCsEsg2d
D24DCcusOr9/0D7qsOw/QxZ+Fel3w8V4RhY7WEesHRlcNRjboreCkV2RxQ0CCm5L
NO1T1Mx8JzRA55lh3DutCb2/XOtfvlXNlLEAx5rnO6nIIz9RzShd8YBxLWUxF82K
j1X4wak9UEVK1KcC3QC9hGTSHQQ0iQSUI0SkfC6IbSl3JN2/wxdiHUlDrmg0ghBX
oqZXDVNozQGSf4dBoio5chzrSCLobyFKL+0yDu5PUkIkqp6EwDwbU1g+nwUvd6Ci
v2R7B95S5H2ZxDmjEULw400/ZRGd9UwCy86ksW0bVLT4j+jebmP0+49+1QT0h5+M
/AityOxatVBwaQgLbLBH51lUF2Uo0XRziorfAlt0IaT0mMwu9LPjLAl+zGsytCf1
P+Jnx3UjxcOFne7lJCp/SFvdFInWQ+tNlYsiPlsd37J6+Y9dHbOTNG2K62B70IJL
RMMmu3TxtUKTI9UZTX26L9oMvLj85a5k4eZ7o1TxpLp/2gbCCTg3nRjEWcGBWyrs
AqQifaApxORiwluBuYjZ6tdZt0K2WjMEc+V9cdWQwAdUAFjHVHkm6UKEAGMHVcGQ
wCP6D9XDl4iZzJuELkr68YXTOSiZvl4BDBM0RzrQpOct8zGBUpNmd80b4WvTO1lG
cBR1V+3tXavVCnSzD5KRd8CdV9Y+onIMgn5+4Fipfsduvzx7oJuNbuVAX2A6Gi0L
V9MUiwWPFf6IgrQI8JWkJ/sZFcqmskWD/nVuMIaQMRR73fA5flixQ9AiZjBAV77H
Krw2doTrAC9GpAAgRYKzpQtf4oen3hU5FRu8vmJKtvik0kF8QgujU4yRdriUImT0
kZvU2ao089bi1ol3O9mxNsfKcoIevLNrDK0ApRvLYg7Ez2UbsxZX5VawMo6OquM2
BjLRMie4yfksprPMZz0VuHIx4UjM+chCjFdrKvIP+CuPafCjKvxcPrS2EwmjYbwf
ci5GFvWXhhLXDt06XWX8uWMKIIn8cimatjaqE3y9XKFJPM3LCjjuWk8YgkRJODIx
5muvSZMEaKxi4bt2GHfDZrTuBy74jfQB1JcPb4ImRgpS1UHZ2eRyXXOveOxUgulh
wHAPDosU9ZvlJXcV4JSQFlF50InlMSPCR/3qE4KX+zfD7n1ZNdMOyVSUQZGbDR7q
NiktZ4rjeM8t00cQ3BFsEHfzvCi2H35FCekg1v+KdCxGa1MXxSwvaCEeZE0G00z3
P0dbpPT51ZeVQGg2tO25h4zII1QpCatWzzWpQ7U75VfumTDG2+CFlzhDQKbRVj2M
dV8Pr5a4EVr+pRHqLzihrxIRxmGu7GRx0GuwO2p/hUX3t3/uHyBnBFtV1J1jeZr+
/yz6K7AJUBNb93tsVz/n0zWcUpY2rxPpxafED4+8JY8w4yrZicFTjWAqK/s4ZZy0
8Cghq0WZ0DcZ4SLXxAw0M/ewwYCvQFhxJhkSior0kQ6KXHmHYEtCbtNZNBEX5TUE
qrmBLxRbDJiOcpFd/pWXRlee+eBAr47NSSQCtcon+Ih/g9QmoqhaVBHMXArk2dxD
C1te0GQctI5/Sn3AHHaBz8EXFee0mQC13bdyLZG5GKwv++/NnLc5Ceh6Eo3To3mv
Kbj54larXoODbgNbwvqfPQylLW5wSI1fWEyat1BN7roVcmhp15HO3jxh/F8DAv0M
Eje1iRisoh3UUXOP5eF3ViNRRHp4V1erHNlFNm+6KcqnVkJD4CaA5w6VesKW8zPE
sl6awhjMscFw8J5REUAbE7q7d6PesvAXZvOH+6yYkxiC97s539NTm10Rb39sGfeF
58taLoskShlqh0gpXnUJLlzQh9c8mMku50sbmUDsXVhTJrwzVGRtxKq0T9Bb+jvR
T5I1hxFyWoAo9bl7XMNGg45aHFFtH+Vqe0WxomWCb3VKFfy8/frEammR8rPf8Hdj
Onpycd4nYXYvr1SFxClduXM9kJ6w2nXyHlq2cl907hOjmi8i7Uf4M2Mxnej7xIkz
ewcjiL50IVAvFIMknkyDQGg3y1W+Uu/0t6F0F2XAkdWxkpdE12YKotZi/VhgFjac
hWn/23r5004EPqzk6aLTKYONq0eD9uspSVpzt1ocZTCGn80P67gI0huDv+Ax9FqJ
TfXAHqvqxqaPXm9YwQc8x3aXMoopfS2+snUcDx6g5c+bip2/rIcHYcY4+YEc/zlO
rP7eSEJjJSHTBq11xjoI/uhfuUDCQqdU7p82UjkKWzi1UNLFDGK9jJGdVC4PkBnE
X8VVVhkWdjeU3wV6D7wyW+of8pDsDx697tedy2UlInZnKSE8bE7K+t/nkRfH7kZ2
KBw9w+3pRJkiGcJNg3zRyHaaWILrUZNPukkgP1bUBFe8gq8iETppnPzCxvphLmaW
0uhXT8F75uJKTBiu2L+30qH/sbSnUSDeVBV3S2A/0n6zqEd3kh4QtRsNzm/aigus
yAo1z21zsXgXL2rfkqP9D5aqTU5PY4thMMMu4mm8Vd493tde1uD4fu4G25sHLCiK
lyd9re+zsIwAFQ8e2igKQJU/bUWcz7lunU2SFSLhPgOrrCF9eqVCr7AL3Ec5LP0I
yTsANVSoY0Geset5meqjiwiFgt4SFRQaZI0lhfn2Lbxo3YrntemEZ2e+/9lfmP1W
PhuRmfTuIeCW9f4BycnvwxLswRyvyH885EZv1e3TgsOWKt9MApeyyDagbuCHjmlK
gAuzGYwTGw3YZUjladqwf+Mr2gFS8XCgkR2AKw3lJ3GlGbkg+3SB/nnHc9FHYbeR
QwYm2q8XtIubMY8NZbcJXvLUld1LeZoIPxSrSah1x6sFXJ6nHWQxfEnBb2uo7GdV
H7hjeFXQZLa95mJ8wOt4j2RkgmonXYIRL18BUWCBkVx7uUyxDWVmtToevfa3ymbw
xrsM+pkmzv3Gj7uhvwuxbIqyZWv+iJpa1FNFMeoto8K03463NjQ/IhZDB6EhuZsI
W+4/RdK/m1o0KDDg9TrR3VbynVnjTqvQtBz7SH2oG4aHg5xYVrK+ChjcaHJBMm6j
v00+EYm6IgidRn7WqLTltIy9q7h/CYItHxWn3tp8/7XgiJVapxUnxIhQyu6jThc1
nUp4DHo5fkuH5bef6Roal4LDATB86SycQ/lxa7pAhqwF88+ku0wIo5/ktfrXah2b
luFfg/f1P141eO+oxhtsAsxN0fKz3V96UpYpjekZTxGLAAmlBj13lOSsk778AA4F
Yt8nz/FD1zVXxRqAypbjNKanZhkfFWZVC1sEvfi5xAHP9zKPm9MtkGzughvejq4Q
4Xzz6UEsicAkeCaigQsSOmvarAaGeNfDFzuc7+4PRDDl9t0+kXGwIoGNlq6WzX30
AAZ3xtjEcG5Xythlrub0diP2w7HqBDe7e0dY4Elbj5Qse4DIP2/QizdITjUr51xj
2kwercLi5ktGD7S4AZ6AKwoPGOfAgdW/ylaaRVyBE174XM9FGDVPvGKwbjl0ULHA
ibKpz2M8Utjr/bemOxjxpI9A60jV58cQE3awXMEMwjCT8shq7Gt4tebUidoQv18r
GOknqoyBjNHwaiP6uRHyG5QHL6CvWu8KBRMW+ErX8+FKNYC7C4ijZ1BzBE3I50w2
SQf/PVbkQyib1xC0we3NOs5h5GiWvT2K5CDdf3r26cl7F/OfsTnJCadyh/Xt/Tk0
04llPXtO+XR2O1nNS5PWC6tikLNRQ9Fst5iPIfqXiaYS4RyZXGWlsKVeVecZfu0e
FG4UEDFtkHvwuNJo/Xld+aw1CjW0vA5F0U0hAH6FspwJDx7R/M8pjVojeEovyAiW
TEB8nb3BBBINswSfZ5phR90Qxaruzbq2En16WhEDNa4vjsDSMPc/6fZNfdWZCBSf
GLEPzwU4VeNTmVe0uSqoHCaHfWHwlj/kjgOBXdRWDpF2GwpbRLRaKVZkP2jLuLlK
yYZYtyN83P9NFrBW/v37xt2NVu1wtDzoSx4ddnxJENQFSWLeCJPr/H5X6u03jaE4
EfEAwbXtuzBgEn8xUxI2XkVaqyCjsSXVpVnZQojn5bu2WamRawcQe48KZz7LUrwU
f0wd0cwtOnwv1455WO1Arf8RAMvVsJjOK3FOuH45tWEdWgB+0cIlWI1y/gLSA0DD
Kx9MuHjYQmAZcnJ3Di36HUASI6qvgaGQhUe46KXl66HV6+ODtk/9RRdhKNZPuZ4z
TJJC9PNM3RwrLkHhEZgoEeXj0U8aHtVg4Wvp6+/Npt0u5o6129+gL0wkJpT5RsgO
7HiXaFrqmTVxgCn1PtNCIsrT4qaExtPSRPWA/IkkDdaP1doV/OxNtBV8UvEVJ8a+
aPapSIPfcHTJgo40PUWeNbmejUdZkY0UbHSh0/R8AYVdc4sDoUBHdKa95+KQVnvz
Gr3pvnFPua5fbsl/rGeCVpOjKYTIYtMzyJGfJvUAMQSBcX0K0cR2gkkXrIb4U+lG
rhsOjUSc2cYD8I3/yBLwzHavDzP/fTDEx4ahwMUoDH8qZZ0cG5FDc7j0XHIXqB9n
ymqn/jU57t/gFsN3aX02VPEUiHU7NR1aKk1J23KYuQlIyXYTNds+HmNrtTaUfcok
c8JN3HMe+DS/NxbZkXt7fDmY7kkYkVFmTRe/NzIuzRUY85tyhUT6jw3d2UngdDw+
6pzZubtEIXzeWTaHZ53jglyYhXNPs7QUm4BIproB+ibQBJsJC8XFIGEcOKCcrnQj
UWecm+ZtR0atszMlqr42mWVR9ZLUTYK81vtaeum1dFj0H4cJg7s1GHSzlG2iMIvA
mlza27tloBxfp1F8As4fBfpGz52TqOixQ5CmDptVr6oQviTotnAtNso5EqZ+/Hz9
8F/xGhNzcmiTjJy0GMymRivIZhKzs/NrqckZ2z64OxGevnB0g7tNxZNOUeZiDdTc
88Rs1z2XTISoGoRMDKfBiFgbv/oxMO4n6nAWPX+7UXFJ+/mFeDlPbp1EIbBo7LSi
+t/Mms+4TLy5tHLxAP22f7pNZ/vARmYxwQr2bgRJ1Ol5Ly28ZduzkxX+aeUhJPH+
ghQJ4s9UXa1DlTDpzp6eLnH9ZxwJuIpAqIofU5nYqFMG1pd04z3PEQy0CfGxIEXu
3vbfqTHReMZ6wGaqQv5mctWY7NSk8HJLvH/s3rPySS+uzQ/DGSFcM3VAEsRpVeuW
m+HbufnXN3zDsjfs6qfhhuxnj4oXW75knu5AWxlCAHY3cvb2cgidht7L/BhQdAJ3
ER0GSAfaCN+RxyUnlQ7qfAi4sdqVN8n/X9emt701VCZMhDY9dBqikecKmmG7ZrZM
JzVN8HVm12aRgTTkSGzTc7pa07022LjJjRcvB5zwsJBysWKTy1ppSDLG8PCtdIUp
de0BGeL4Z3lsRUxe8Ld9AVJWIAQ6XvSxvOu6USMJrYl9SNHfYSYdVOj0zWn/dsCY
6nHMMiJNUcY4CwLd16TbCpNlKMaQ03RQ7g4ZoJ+gZo0y8Pqx4R62Z2gTQXX89kyg
R+cZwsmtQz3m+FYGOLJP8q9ELve5CFE9SLONhNMKZadR+xsZjl4iRgbllVj4vc/i
xrQs4lrvkfciPoUo5/MAIsGSPHSat/5rGNGMLTlwHdZjKXHW2FlziK/G8AT4ExSr
EzKE4KTk/4+Rfdc6EOznEPPoTO3jlEKu7Ng1IUGOqAbwdRxp8xDpVmom9jFO75Pf
ElozqYpAC8zSB8cMaSomdvVcjCirRV2MBg+69smdNgBlhu19v0Wl3K4jLvvyp0gX
X9S3qgILhI4ZN7UTztx1o/E1tWqpSxENx9VlfqffnxtfFK/jF2iM3729xBn8wYXz
/IIlCgt6pKNaaoajLukGj16mwxJEpYJOwLEBMIHu1L+aibqZqImJOdNJQjDgWdeb
ssLxOFKrjWu+6dirhKm2hzhA2qjehiv/u5otq+NYLi0SxlnCvx1j3jnbTGQaWOfr
96dNprnEGBbwhPLwJKzlil8YqtDxqq+ECpkSpMZUAguvC1kfLll5zXkjlZEuUbZs
6nvedlv8rST4dqhjqXnezUikOr/d/hHD+cJXIdU2IbUjEJXD9Y7FfHZukXPjhc8t
y2/AixEUuzWHw/hHZ5dfDBYsA2uBlFzHGZkHe0C2mADAYwnHYyJofcE0SyzzD9N1
ag0qxqJpVsFrfTbAybyx9f07CKI+WWZnxLaHb3Q9BePPHxyx5zwUEPasOCp7Wrh0
StiKd62W0n5GlHUJyuzgaSvZ4ZnlQcB3Z4MUTJ4hZf9Mv7tbMn1155e+9YlR4DgJ
TIZcqZpyVAuknltUdKoORpRb08QmVrUrScBU/xD+fcNzh1VLnjXsJ938Twsuzn7H
eBy1VXEZNHe1D6tBrI0D2mGSNhb7qXdeHL1TFD98UdH+QU76QVlSigV/+ulm5Fn1
NPe04RSSJUxDx+tCluASvfgE/PAWd2XK4X/rkuGCEn20I7yaYIqJBrl8GABLOCeK
NfPObfomF4KgwEKMl1rBUnT4e5KW/AP71yxCs0iVHqZbuc1svPUrNXncuf/jyivn
k+BeuOvgtwy9UulAvVObOzQRoAPLmY2KHUQLELwA9JFRGFNYamPKDq+Z3dOji08g
Qd3mXkO6xrCAaRT1NQUlGMMHDurU1n6G7KjK0dkP5fIcC5h3kGqy4n4hgCCPrP4W
rlhslkL/Rv2X0XNcD48YiYTbhLtJc1RiFUNuNKVpUNMSvRLzsO4iCd62Eq74V7pY
cR30j/SLRLNPCgQ6bVFezHd7Ign53uN7Qa5mfFVtLWZbXHsZNXOZ0p6N7bI/1E8Y
e5OCaRREWjclK79PgrCmXySorycPQCTfXEfc0Xk4NqaBZEuq7abrfviszpC4Xwgk
8BwfJzG6OA6AtyCnfxnSpifT/Pq57K2U7bG31UpEfysontTs072Aqjq6dJMxJXYP
O1qAFDf5xk5Fn8DOrgdsQxHU2poA2QwN2GB7xAdiOUi2jzLePdHHaCVIb7dMpf1h
2Ecp3zvKWRxu7Xgh7x7BONmN5Y729L6whcQi9lQI8AuMZCZGTcfo2G+nHJwWj1hf
QdW7j3epMcejyx2b1nNV/tx/iCbhep1xtMZkZ/AejP6JBnPqRXlUuESWMuxwyuvZ
nIdNEkE1FJt0tRT98v6nVjaUbO/pYg/1mCbyRGm7mVvJQLBBzA0HSrorp3yaVMZP
+4eTnve0B0OKKla0WuaIJk+gbsn2XgAaYCJnpYin8jMW7uUjN8nYEu7azQ01ZnER
0Kn5ubcwF8MPI83L9yIXCmCqqK5KXQxxcSy4uzD4Wk6j92VWojxp3WkNUsxaGaxZ
mN2EAtUfcYrWBMNNyfzN5dxCJ4N1U2q4yI0nPvuezhxKkTxnWpDk12jPULlaPKgd
nP8yqxKkFmjAO2TExXABuM36BYPlkWnBW5sw88/dbk95GwWTjZm29z7Dbv/fUC5z
/6XCgsibqfpyAJHV16rtlQeRrjEdFZUSDfCGodw5pjvXQtQvIW+XLNmBH3mVIr2Q
3opTHsnUQdXvwODDAzcRVFpKYk3ZXm/7ZbQL6ggVqiqmgQxQy3sQgBPyO++Xi6Cy
DVOkRWoobPmLmv0daO4bQcO/hqk/K8OzvjP/U7lnn8nGeTploCBIhhYjtrjCnSy9
U97jeAyOcGyZh0oDjbi7m7GByyjZut3Zpj6f7l2HL4rcHiIJ9Ok53Q75P5QrL+W+
2H3z60d/cths9q4hV3LcWg+xxbU2/+d3Yq8qckSi3mD9lDb+QnwSrz+qL+qTb/ze
a3xilXa9MBnLgYCb5kbX90keevGu/kwV7Hq5wFCnC/AJVE0bnx4rpSIlEpa+c4Ig
EYW4Q+ixiYUT6sWCXmiOOU0R4BgxrUYu+zoVgISRs9Y6SEq3CtDc8yyiKuYs5epu
l+XKimTqpdOjE/cEPs+t7wTKYtGHy34xTcojFEB6i7J4e79nZVXMkl5BmATniXb0
1OHuOvZCAHE5AEMb+rPqBzUj8S/KkxduXiJkvL2sbdfswJDaUb+wpL7mkQm13JnD
nXyXPob7msNmwNcvufwpX+8U3dPZjb68Dh2PV8HqCYr+VjgUWZVl6jKW7wU39smt
DPXN+9DXPWwRUe0iIY7xsIYvLiKLBMMaALC0GTgeNpjjJJtvC6tu94AVnMdJkMyp
Qm1iA0Y1ibhIE1AVhaebhlHd8ggXVqbWOz6zW8zmpALLIjIuZDWsdmONdGrgqJmt
VcVtmVR2Lr66j5gFgFRVpvalzrczWHoyzQB7GHQSH4BVnmqXB1pXj7LHMPwHE7V1
jP+YMU3h4OQHm9gwQ/jA1kTt27y7giay/v4h+n/DWhcYGsnOV6AVIIxwr9jCoo1i
Sj5r4BjgXJpN0M90MuYZ4R/Slw1AMe5TYSGm24ogiKQPSf6/ENdv0pZtOh2Ce16w
7eCSe0wf2LDP1iTfPUGqc5EQNUzBKWDXonQ/c8btrWeaKVARx7qIkW3eFcfFptMH
m/kcgDNhVzgirsvmiWYbCGDIgeQb38aQSQQ+SD6qBr+1YJLnRIE4+IeaTCKw25Hr
hD83UFwq/MwHOJx647xeEWhZ+nvh7ohjeZPOMBSD5PbFxTUmU3+caEgvLfMGAASw
VFXRagKL6CHzC7xIZzeOb39KM/vxlCO4NNMFhgtzeqFvQTyrvwWXDnOtfd0K+nqq
fb+0boQWYBFvBTarkyOvQDJydi9wnGKg7kEkk+7FcftQ/5iksuiUzwwYVOWuv/KX
JzAsMcB6nsUMGg2SkD9ESgqMFWoWh+fF+7EEJZq3Xv1W2+kl8EDUTMw6VPxt8EbY
uOS8rDCMYSuxEtHN7d+x3UKz9djD/6p3cJ7C2NNeW/Y=
`pragma protect end_protected
