��/  �l�z:X��t�qu�rcҘO�u�1�O!@Fw�}���c������1��*o�BLA��öog�7n�(�4h^{��O��s��Yox8�UTu$w�a�$�Ї�m�ڳY:���G���͏��ku��+��0����2�L�����*R26$�~�М��Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9��ˀ�]���G�-%W���c�Y|p���םT" �X$VD�盽�Zme����4x��`A�k
� k��!�5����V`#�3��?��nm��������d��Z�IY����5�FQD*�/p��X2��������kP-AK[��/�h�Q3���=��8/&�L_@xD˖6Ԗ|4����79sb\*���ե$��ƃ�#�:Ń���V0��:��m�3��E��}\���]ԯǆ@ΌO�$�Jպ�� %Q�D�=�6?���}Ӎ�N��wߟ��􁨁�J��̻b$![K��^�zc:[׿c�%��M��V����SH���Jo@��R<G����o�q�M�b)[#���X:�zpI��o۟
1�Wr�`���6�[��kf��ϋ��˄���.���E�˺s�7���0�����ڛ+oH�X�Ƙ�6��pA���SC�s��?�x�^B���vSgM}�����$c`����F����ѫ]]ćZ)t<>�3�yb�Nu\r!��/'�7
�c��R����������qef�yT���b�+yD]�Ct���B�2J<D	 �˅�V;}��E�
�U�*J����+��mo�43X9���Ŀ'ܰ.)�9(z>�j�zN)q���w�	���ҭW�Eæh�N����)9
�_��f>[��ļ���w�n����Z��,~��_:h����g"7�>������H�-�щ�� @�N�w�I��@ȓ2o���}�ߪ;j�����}�+*�:ѱb��H~�=ɯ�98?Qm��'��e1�؟�J��h��F���k�"i��m�X�6�2�8�Nw�h�`�P̳������:=�+�k���m�
�1�E�8�n���'���^^�G�
��ʫ��2F�36�L櫢Wqj*���n@T_ta�_Y�IE���Q����+(
��[wC�_"ݚ�&(��i6�強�I��'RջC��qO67$L�0��N���V�%L�"�+��v G0دu\h��)�E]mey����{�kd��{M���|���i���u@H��~з�eiX%��٠ٗ���� ����������Ͻ�b�i��_�}�`ڇ����
c/�M��P�|U W|+l0�J8�ɉ���E���@~0
���B�D�]�$�L���H�96��B������J�!R�F�v}O���U�:�;�6v$1�ET��{>�J����t�&<���3����ǁ~�Q�䬤�FckA`��=�ьr��C~d�B��^n���OLA��9��<0���́jp(7�"�_.�a ��SӖ-�����ץ$�Y��H����n�G����J܂z/yd԰ӗ�LS�Y�h ���l���|x���7�נ��y���I��٣�_=f�y��烱��H�_��Ԛ�v�(	����]��L���o!�s%���ǩ5�o��M�V(��V�z�a���Rypu?�6���l_!��͔q�?@�毹�Ã��Bٻ�d���7����V���XQ�z��O� p�;C 3�GP^�瞃��W8�k�d^�?A����s�������C��2K����&ɹ��!`�(ؓ�*�Z^�cg<�1^��lF�:tGܯ�Q�{xU�-��[�&H�zSf��Aq�*��R`��F�2���7@\Cٜ��t5�Y�� �髜�s�x�ۤ���ms�^$K��qX�b2 ��3���+V� 5h���~ߨW���g�l�������D�_��+L�C,��'1v�;-��JuJ�YD\�L?_Q��u+5���u��
���ٷ�G�F-b���󱛄��Vo1���w!N�w+�[��[A����f�z6���d��A�T�o�*#aZx��淹'�Ɠ�#�Lh�*�`^Z��_T0�Y���֥��lX�.��
>ۣ{Q[GLդ�'����$��Z�|fYW"RM�D��Ђ����?�ߵI3��$1���D��(����+:��U�F��@r5�d S�_L>D~z� F2���n�A��W��
ر{��n��ל�)�|�� �'���> �~����`�'��=�h�n���q�3���mȣI^�}<c���%	��lN_�yѮ0ů�Y��A}�Y�zq�����>^�$��tل������e
ہ]�Qi��3�q��Ѭ�6ȎF�L���I�1����M�9������]����ĤV�0���0���4޽�,۾�)��'Q�1w�Aױ����mMc^�8^,��?�<��g�Wv�|��X1
�!�KR_��Lu`-��#��P�1����4����u]�`zYC��_ b= ���(����HߞV���{��
 h��$DSy�r�?	����Qr>6EG�Ơ��F���\&����7��E���r��R%�
��1�k��!�cb�.-��G��I@b�@	�zDO�a[�e�O�/�y%�S�����f�r�os� N�z6��憸Y����g{�9�!,A���a�bg�d�r����NF�4�p�!H��|ʵɭ���Q�o�w�#lҀ�a���Z�N�zd��_&axtIN�������	�&��x���H�Ĵk�1UL�R�D�G�6���Q>�h�]���?0/�i�n@5/��p��\�2LXǴ�P�d�ྛ�V����"�+�))�t����(ߧz��3Ǡnc���y�:_�V5>�J"tr�Ҟ���Rw��BV��`�tM֎����H�3�{�W��(ׅ�g��R6]p�i4� �B:������I�}�إM�����#|>��0j�lO-͛�~Kr惓e羀@�H���	��2}pMշ�5����J��|y��	�&�[W	��ܙ���(2�.V�-]w����1��d���F����\��ʪzуce�t��=>����9�0��Y|�<�!`9�@}*��!#���_�K,�o�*�jI*��4��mx ��}C�d��	�l�RB�qG�~������*�?xp��� ��$n�e<�ePCst.1/�C�� J��FۦQښU�׼��z:6��X�R ��H9'ڏ3Z'�Y��=�R�&̒ �cp ���%��x4Q�\AF�wb�ST끴k7|��<BM���'i�i�&���<���%/�~��3,��!htH=)oWFY��ge�F����c��9b���h:���PסL�ڊ�/�|8¤H8��5G������÷�K�@����9����W�6�t� ev�����Y_�#��\����\����(���dty�)��Ժ���?v�����2C�h����"����쁬�|(.�[')8���+�1K3�{�vm=Z�K%��i��L �T	�#�	
�+'��-���~���Ҫ�����R�#F�5��p��?kݏ'�+t�E[��dbT}@r����ߩX�9B
�=�q����΍�؝y
�6A�Z�W��|L5�_�r�a>��PHY�Km���|��4p[����Qb�U���O�^��2���9>B���Fmya��������հ�����	(3�xys=�����t�n(�ȚBA�4
U�v��MB����.6T/�A"�ż��.m�� 6��k�z&���+��$��y%zKm��碅&&!��{���GuQ��E���������J�\Yңmݰ[8�=�9�,�VE�/#~Q&���s�F�Yhp�X�K7��Ճ��_s�t���޷	��ZG����^Ӹ�We�F�!�;PS�8��J���?��?	�4��P��i -��:���T�����)�@�'�ҧނX�`��P�<�b�Q�E�W�&5���������g ܐ�
3
�	1�{���U� 7�n��u��ܚ��
�r	���@<J�%��p�7'���Ւq�wK��@E��ܛ6��43�I��)W����^<ڻ���{�~���kH5������IƦ�/���3v�����@��f��>�����y\R	�j��ss�7A�-k�S�_�����Q�M��&t7Ҫ��;ģ�J�IT\i%��L<'�������е�7h x�i�������v��:�Gnk8�a+w��rW�1)�5��dS��oBO�+6d�=k>��naɐ�)W�����|�	^�����=]���d���������xđ��vT��/("1/�(�#�R�S�z|38�gl��K����lecY�{�ٕ u|f�<������d8����E�&ALE!�;^�.�z�J��R��� �yk0��k���-[���t��m�&Tը���h����L����~���nK}1���ӽq���A���Vu���(���R'��o\�X��Swp���X�Y�z-U��p:%�dd����pž� %�
��/���VR�����p!x��7���co�S�u�'Z7i�toI��k^'6����މ@��؊�i�p^��aL2^�;~Gr��׾B�Uz.M�P�T��?��n���4!��P�O'r^�A�3{����B�0r�Aj=(q�U����?ߪ37z���?aØ��'�L��:w��>�u[���
.�tl�r yU�<O�,ɠb��˲���K�8�l�*	C:������P��6h�/HDbP,����-Ҭ��{�d�����Qk!޹��jf��#�&d��
e������@�Ζ��LW��Q�17R �_�?��*�.��,k�#�ĶDZg��cR{b�W:{�5xQ�����6�,�j�����?�Dp+&ƺ�F&y�����-��l��:��8������!�P�|�a��竳_'� VA�;���<��� �!$�>7���ʣo7��0=E|��V�ijn|DԐj�t�r�֧C�/7X�*�D��P�ݸ�@�Æn�Ȇ}�m���zR_�jE��S�:��2oS�L���|�8;�I�L7��[����Ġ�jeݠ.��2�	lW�������-t�G�Z{�	6tg�CZ��^�Ⅲ�lÔ�7o��`�\ti�s@�P�I��oI���(�Y���lK;D�`	\��CM��f�ޱwy�*c�����nW����!�Z�͛��|[��v�DE��.���؞��̿j*IN�V���7Q�܀�>��� ��	}%qy�3[��p}JQXЋS7�G$�F��2��N&�>O#��n��r��g^�u����N>�lYF�������"����KK�6��Ypԯ�O0�ő5�"��}L�W��krW�����	�KR��O��h��V4͛��a�A��t\:dR�d����.:,4f��lTCX�j{�{�2Ċ! vS�A���G�X*�Mÿ�)Q�5(�?�YC�I�B݂k*�����ʍ#0lE8�z�F��s*p9�����r�^��D���{�Z)��>oע��B�u7�i�DG�u���t;?(*�)����bDr��e'�����ͭ���UM�����t�TF\#D?��7�¾Fv�V8U�&!6}S��Z{�����@�*�f_9�p��E�to����è밮V}<:ӵ��`n����z�!Cm�ݵ���T��N����<��C��ϊlP�s�-�/���nG�[4�i��	��-��a5�Y�>�-X(��(f�=b7C䊮 n6
,YM���]�8��2�[̂�T��0����m$-F�r��+%k*f+I��߉(8\g�U��Pq������$�J*	7Rw��������}�B����:B7����E�N\�� �8+Ď>o����&�5�!��ư�����i�w�p��/b8M;7��D2ɘ*U���+^+�Ձ⽱�P��Q�e�[uPV�7����0��v�y�ʹg���a!�95ᕀ�o���&c�k���+ab9�:=�����S�*C�9�۶6�猞�c>�nJ�&?��Q4��!��4OP������aU�5�1��\y�Ҽ�>�QK'�p� ��3����6{*]��M*���̰�lL��4��+�o�������-t46P���R7�-��ynxr]%m\����p�2V§5��ee��)�[&�K��G?�ǆk. `!gV�\Ow�D@ZP}/�<RpPd��#��BB�Df��(��Ϛ��.jGd~M�����vS��y���Δ`ƾ�h����v��o�K��y+$����q;�B}���Is�L��n'���f4@I�?��dC�B=�2�`�zF�62T8�
�m�^�x)��k������o�8�V<Jʆ'����6M�ɥ��_ʢ�?���-�
W����t$�*���ns���
4r+��M�	AeU�����I��p(���	�l�:��W�c&�{����.�x�j<q�f�ۗsռ����s��y�`�,�>O��� tC����k?u1�z��V��uB{��8��i�����X�R��B��?��!oE~�ilŦH����Mt�x���hѮuʯB����E粦��F��E��~��}����t��~*�e	�l��A���c��hg��Ȋ���Ue��H6!�B�A�♤l�᎕Jr��Z6�~����p[n�A��n�/�3�e_����D��T9�6V�Vg�{+�	&�B~`pS��.՗�Ao�/$�T�G`�D�����W«��F���_��4��7Ȃ�����G�����_#z� �B�KQ	���8�)$Ƅ�m߆���� V���L�qk�ks�*���Ц�G]�b�ғR�yTE�)���(������:�v�<�B�4�<Q�4�bX�a)���C�����D-hTo�X�k��� ���`n�a_��m��C�T"�$���@l� -�m(g��RKD���?�����72Us�"�pkM|(3;9e��ٷ^�V�4��{"�0�!�\�.���LU�U_{JC���r�,�!��3�����G=�����t��b>U)�k"�2��n��BY�	Mrbj�Ka�
��e��u������HE,jKg�nA���H�[��K/��b�li����Q!���ʃ:�+.�މ���ז���%�QܖMҤ:�T��O K�0��)?f{�s�^�~�8O��O���+�ߌ�h������+���rcR�I�M�P���![+(��y�oRr��`$���=�*u�N�#y�,��d�^
���=�=���S�?s,	���v��Ic���,��ա-Lʭ�u�?wP&�W=�{[�>��֡�nk��B���#rR©����~$��]��U�P|�Dn�x�"��`�����D��c�W�z�1�e�o��#�5�ܺt8~�¾74��ɳ�%j�- �!lP�N,|�g����BE'���7ݦ�"[{�b�nK\5�����s�Y���G��2EX�h~�1�2���֚�%Q�+��ӈx8�m�2�R!����a�	��#�FX^��:�/��y�K�'X�z�r9ӧ�۞5�O S,�]lq(;it��<�y*�ʤ,��\��%�Y�u9U�y��=yQkN��g��.p�.5/&�"��7�,b`fg����!�Y����-�No�!j�{��˲�����4�j�� * ��0��R�X�����qc�>Z쓢jZL��o��EC9�|��D�9#9�� DE!b@TX��"X6N&�k�QN���T?5� S����?���{O�eD~?-�>�t��0�1tu�溚����^��(;@Ѝ��ò�~,�	z`/���(A�&%��� ,D���p��u��p�j!	�ފ��Y<��v>: ��o3�� #�e�f�Vz�m&�)ˠMȮ�����2��Ej79�������E�o�߻
��؛����!S��c�$��f{�?�]cB�ɑDÜ��S�Y��%"�'G�Hc�N��
@+�\�nTmk�l$�����w*d�H���1tr8t=��@ץ)�>��	Q�?h�� ��-�RΣ:��F��A^Ƴu�ug'�P�z�w���kˏ�w���	h�)����G�#�9�&���;�A�m�z���΋�����ר�80�5��(����(Ka���sz�K:^�N�������03�#��S�@K9T�#���XkR�B��22���2V!��WA�����{��U�'������S7}��BF��$��'��_Qұ�۹����:�"Aշ��������.W�OΖ��jI�,'R�K�����?:�K���s�������)3">�ą�L�0V���v��>:0���z�R��-K����=fy�֎�S��N��/�qx]|�"����4�Fح�p�0��E|��;Wl[��绩��.�)rˢT80����A�`nP�BƠ��8�G��7���0��G)�� ��6��d?'P�!��K"\�Y��Q���F�{7,�R��yr�߽�*4�`���0S��I�~?���eo`���������J*F�����b��k�bo'�+�קsʊ��<��^�>�ư)����ъ̀��{��7x�CB4T�>ƈ�v�"�#���	�K�a���	�R�}f�<8z���JB.\V��B���M'{iZe��L��vr��pV���T�D�*��5s=��o�eqK4�fT����^|Kw�2	�M�����ڈ�#x�9�*��frX��'s_�%� |^?
����gCd�	�hi7��K�4��n�^���*B��
w�X� Y�if�F��� ��'��?�w��	��J�'���mW	��?9��^>�bj���[1/��5��^��SRt��ӝn~r2��������g<��
Ki���t�O��_L����M�Q�*�Iޚ^�kz�-��t��מ���B�i2��p�����[r���KP��H??��A�ÿ�'ֿY���9�B�l"�b�Y�U�yw��
d(H$)g[�t��qfD�X�U��Lë�۲��@ƅ�l��:��,Y? ����}�~�1
p���R����"[��F�>�Uo�")<�0j�d��k���:�xh���p�r�(�@�ڤ���Dw9�8�/~�;����~e\6��i�ڜ?Ylœ�~udr��:UR�O�öL�V\��+^'��R�la�V1�m@$Ŝ���f��f-�R�{�����w�d->��Ά��o��f�1.�,���]Q_|�v;܊�-!��{�M�Ȥ*���{b�7�v�l'i���~���BI&��^�,+3;kse\�Z�)�:��%�ʢ�U����#�IȽ����ن�ܛ�}r�C���/I���]S)�-�g�_ !W�3R&��t9�IĜ�F��Ox���I��5�D8$D��[?�@�mI���L�Ҕ�)���m����ϋʞ�z�+/:��ae��r���s���M{��͗���>Ʃo���� ��.�sQJ����L���g�$L�w�� ���r��m�t[U�]��(�^��|��T�1c\>�Ө0uH���2���H��3�#p��F۸V�<�DT�X��\��m�L�"2]�V�u��I^$�`�1��Sّ���"+ҫ�ϽB��%kE_�rƫ��CD�?���v��<Q`��"�=�-�rc[�Tn�	妾Ư��(�0`S�F�.���F��ƣ��9w	�s�d��Ay�;^�8�q;�ܽz���R=���)Ҙ!Jໟ����@��D��$�a��!��QV}��i��+iQE�P��ȱ&�vs�2�3t�o���NF��!EN3��T��h#X��!��}��Gyǌ�u�`��,�e
�c��͢ $�ɰı;��o�CE��2֣��7#֑Bj�˫<[(�J���hl����w���Nғ�Ҽ/���S̯��'6����"����k��� ��Fv��-`$��Q��=��%��E<uN+r��V;	����QT{�3��Zq�'"V�->��5j12�z��en*�-�Wh�����z$�x�~�#�� 4&?�E�����i���\�ADh��%��NVk_�,���gC��`Т�apNӁ�R�Ǻ'�0V�����tַ��E�;�~��J��{>�I�������M�mבo�ߊ�>�O4壘D9 M�&}(LW����nO�~"��Cp��2{� ���t0�
������F��F��%������찾��8@�4¼&5`�T�r@Y8�^��dF�/�7�j�FX�i�/(@���H�-�%�1����I����u��)�f����K�����Г�������z&��Y�O��4����}�ĿO�*�)\Q����/�����?'������c;�j}P+��@w��+)$^v3��j��Cx��^�.
�~$5��e�m�vu4?���/j�?ݩ�{���]���~?c�@LZ���K���ی; ����o��������S��ď,���S�H����cpD���C��:��H|@M��D��7��W��MG��w/��׳>��d��8ڲ�L�ￋ~�<��Nj���"�pP�>�1���\)��j�^�~���������ߐ�t/���4����3D�&��D� ��}86Χj�P��I&�,�2)�6h
ܻ���x�ؘK��
݁�і���k��������z�lt����kZ���s���=i���D�~۔Q����=�1E��}b0#vq�T�ۀ^�������R�f�����I�g۟b�0���;<%)C�Ot��J>���d�f�Aw�#����[��z��g���x*q�~����%��Q�մmN{ڗ�?�u����J�5?�	�EY+�������Jh)����Hea����C����q�j�2
\-�
t�pFJ��_'<Z���}*B���w?R�n)<���ߖ�{��Pn���@�1�i�Q��-R�O1V�����:�׻>�GmF��yq;�)��ԣ͍��Ɵ��r+��f�{�v_��{CE%EG5H��-%�u�wQ6Y�T�9//yF����̣S��l�M?-d���������A��ԋJ�HUV�����{_�?�ƺ�L���8�UG�� F[X�Ӊ��/Q2$K�e�;,z�;ٗ�L�y�CP�+C�.	1���UPU�J��Q켯��&�w�h?W�0��b�)�<������Y3�T���*
�K�#��QDt-̉UK�3=�4w�/�՞��B����{�a]IB����CЮW�9Ǉ���xp�
����
�i���䵙��%�A	�!^i�3�C�'Bs�cZC�7��s����e%���GK��VX�sdPi%Z<������H�(Q��`uQaR���G��'W��V���H��7p[�Z�N΅�����$r{-�c�q����EB��%���e��UX��O�kB]&Ԧ�=91�f��IQY�3�B	�����9�ʱ�rL��?��ʬ0��~����ٹVgF]�۷k����ed�$�r��/m�^��$�@��0zW�F;�(��3���Y��[�.[��4���H�J ���r>�K�7�`�R�>7�^���`y�Yl��_�[� ݜ7Ŵ�QC���0g�_���d��s���L�Й4c(q����*�4j"�>%:}?�)�*i̒�A�ř���ٓ�ܦ���G0�r�����E�'���f��`�:�]�m���K��y�v�(�3�#_π�m����Ջ��<2]��ȏ���X�t�o�����WA."�XI27?%U3�@�8�;�ʒ(?�3(��>E�ՌZ�w�����B#"���OmS�K3-nw�ߠ�*e$�ʭ v
	����յD���4c(�^@O���GxI�C@U�3�-٬�덵l&$U�8K��668G�2�Á��[fuV�b�s��~�2Y֡y���Mx�|9ĭ��I�	���Pqŭ�o�d}�T�\��xL�H�m��'��V�c��F��+V�y�A$ӷ�\_��99�������4&�dR�wt���;�C� U�ߚ3H�k��D�L'E��P��S%7Y6�L�ͳ�Ⱥ<���G<���D��� ��(��$�����y�#�M(�zy�D�Ж=nm<E�`�k	W��*p��l��������'��iP��) S��֊��]_J�ya6*�c�Q^=ҍ(��쎰���Mc�ޠ@&�����囇�a�ܬ��UƓb��x�iS��=Ց"�=�>T���9�cp*��q�Z&����F�V��Ak���m��HHmǻ���7���_�YmN���M��O��z`�dz��� �*6���3{M�-�ƹmbS k�$]gnx�H:h}(�?Q/q��v"j�ޣi���/��&����K�(�RD�T�B�q2����40\	8,t�(x�l�$)	�׳�`�x�k�ʙ�?�+�Mԇ�S��-�J7	z���:E���P�lD��Ј�Ķy��x�GT��t�ihUd��0���>������Y,��ԯ�F"/Tˮ�"89���Aӝ
�:�hHR�<�i=�_�SF�}�ekgEf��T��M�>��H%x} ˇ�W���TB�hd�~��q	�T��n�Pw�����{ ��Y��٫��i��9)Q�͹�@U����|��(jD���Q�JT̤�k�32�#���\�O�{Ġ��6S��Kuo��;��D��C��Vv���Y{�ך�[����s�9U�f3("�5c�l�[4E�dD�z̰���7��ۡ�55����)�YvM�vV�Kvl��Hp����$��Ԍ��s��c}U�*c��!�۳�-� �cF�z������Uְh�Їm�T�."�8�;�'�%�v��k2�����N�cބ�3���"��a�J��Jdx>�,X+��a�K{� �i���\����ȗ�s�c�<.Q<_�M���קC>���o�O�)㬁�b�M���&�R�
9|_�r}v�;j����;h�~g}R�Lh�Y}.oZ!��b*�w�]�36'l����Q����a&�Dyʪ�)��`^RI�K���B�7�|,,�gN�u�����F�&ƿ\�%�Q�Y�Ɯ� �2D����$���j�s�Ɋ�W-gmI)�{!4�t:�M//x����(��ͮ�xm2,7\d��|���^"t��o��/��)5�GTI����CC�n�����G��Bm%A �+p}����2c�(7�%�������j�l�I�\8k�ȝe�8\YGo>��,,�ޢ�Ӿ��F����X�4��F$H�Mz�: cd+�~Dz�7��B�o���',�:$��t�OUM<x0\mD���Gݽ���{])B|s�F��b��6ݞ0h���~�pԞ`��p����ώ~�Q�+C#э�p6�񏱹�+���-�\�G�K�Ɓ�-
��D��K�Ľ��J��⇴�xQa�G)hT
s��_�9�ǫ%h�^9*�i�/)���&E��>��Q�ѫ���2oR�u�8?�:��0�M�b) ,Td~���[�����- �l(���B�t�H��B�C�}1��w��T�� #�B�F)�8���Ҿ+G�^d�Nʨ����!��38k�d��y˹�h�3N9�/�7��δݲ�?��r�i3S��}NZ:��"�˜C���oO�ս^+)�yS;�_���!E��?B�..;�L;ī����r��0�d���G7�>��l��n���)�֗��c��]� �8��mƼ�A��+�{I�?=��T=����#�%sB����v�ǯh���V��R�R丩N�uj?L�8l��\��7���>��FuL�(<׏�i��U�g4ߔ[�a�a�)���)�E���P��j���%�����Q���x[L��[�����Hi�	��G�%C?�ӻK�f��_q��'��P���=rږ��G����!����5R�c<��'L�i|�i���G��]��z ������uك�Ax�=t%�BmP�*&�ZN7ϒ���-J<��$

��݌z�d:1>�/���0-3�$Ii���g���HڿՈ�ש��U��L@s5DN,=]�0fPg&.��
 ��m8��ů��ig�|�,q)j>�F�ˆ�8�Nk�ֶJ=-.�9%w�����D��L�a�F��p��K���r9�4�/�!�w$���(jp��u�BQ"��B���_c�yK)���Ǽp5�*d |�2W������o�'C��o<3	,��4��ͧ�e���l|��{��[�lf��)��!vD(�+��qj'�4K�����f+ρ��[��/���Ƒ6>v���n�Ʊ��쳲1X�]|\Pq��_IPw�Jy�vT�߫���K��v�&zg������<�V
����_m��&
 E�T�g��~��o=R��(�)͏"�[c<<�~�
Ulb�
\����s�-�4v|^��h���=�,�7[䨱d5[�2vϚ��H����[MX�������A�?ހ�]��.8fz���}�n��Ց���^�{� Sa^�-�j�˪>�u�$dP�1����T�0j����Ȧ	%VWp��rбmę�:�]y��Q�N�-5ӄ�׃���9�<��Y������9 ��tJ������)���'��ң�����e�P3����)���k��~N��-6��a8.��GbS�� �0�<�Z��P��ӉT\���SU�F��p"�nô���[�yU���g��:��V��ЀB�g�]�;���r��c1���������ݖ�"aF�q�H�d�0����'C?���%���'�}?h���ˆ2?#�%�g.k��3��bwzT�Wj�xpߖ;`�H@f*��z�ck~ƹ�.�*k�hW7��lq�/|�5�n�k++�E7��S�v�dmO�ĭ�����%��}��y�Y47�~D�y�����G�����Nȗ���wZ�y�����r;�z����aN����W2��l~r|�{�`�xM/Y��l�+E�V�D���#�&���O�!�v!?f
���?3`�J���a"��iC92Hax���i�N��!^�,QP"�,�p�	v�Ǝ��Jk(���@5���ݒ��"�z�q�{A0��;XI�r�gR����XW�y`��䲻w���"H�J��t����]Ǵ}
�)V_<��n�>���'����٨��q1KӦ�0 ���Ј�"�>���߰aZ�°b`�#l�ZpcKl�@��$��md��4����r��K?����ו�;2�X�ة^��CV�Ο�3��Y+�/ư�~4\�]�ʮF'���7�St�I�H�2o�\c��&�@=�%��bk�x{������hY�.��盖.�r���_��Ay����y	�K&!��8�73u������۳��K���Ru���C��ӭ�AĠNv��4����j�'��:׀'K8A���IZIm��H��n��*J��y��V���Z6�_*4���*���5��F�%���
�s�Y�����jU<�4l����@"_�Ϳ`q6M�q�7�/�n��.��\oYے�!��*^�7����Ӌ���|��ۧ��
U�QM��6j�|ub�e�����"�E�ΞX>Ls�Բ�&�B�$�Hm�LJR ��6�hF�CoK��393S=��8�ֱ	M"�2A����b���Q(�gͰ��:�aԥ=���1�eB�C�)d���Z���Õ�J�Tx>rD�}d�3�ع��T��՟sC���C��G��ꦧ����i̿����(�{@K|n��$�s �iZn'�FFi�;���AOA.�.�������O�%E���@u���s��;ƿ1}�%L�y�W��3:�F�4|���H����6yT��ff��~ȝ?&��<�~;����=L������
 �T5$Ҩt^2#��}���$��V)�P1��#�6e�_��'�ɍ3�9K�r�6���/q� �WE�"0�ù��s	>�)���AL9�/me�K>�[e���ծlW�i< w��UOu�;|��*B�Q�_�X��t�6�����>Y�&Th��q�L�k4� ��:;V��0�ҽm���< ]ɧb)�}G�|�	�F�"��UfeN�Uֲm�ԥv�	J�/�W�4bM�ay*"ʙAj�K��e8tz����Nb3|��SR�\�U�m'���zUf��b����&oPZ�/3k���d�9����r$~6VG$<n@�Vw�o�0:C�O�+���ف��
����mmS챧��u�4B��3P�&��P���f9��5]��`q���~�Ti=����:��YP�(�M��Wo9=� \_�o� ��8_�ޟ�ӄ;vE�ͦH�ZR���I�����x�h+�%@�"�	��[�:�
<6�\m��~K�+��"٬�AS�:lv��Ǻ!����2���"����`�Y>���)c�8��z��7�'7��3������Ҙ"#m����Ŕ� ��@�Y�A^��I�;�>�|�>�霾���&���G�{�&c�Ƙ�P��1f���`�}eL [�x��T�OA����i�rPy��BT+#v6T=����ӌzi��i��[����>��NN��E���=#�jR�-�� �=F��Z$�;��{�Fܡ%u��*$�`��q��������,�(�^�caN�+8��4�܃+�&K�{P��sT��7K�ִ�b?�W]��ʔ����]yҤ,�j@Y�di+v	,�*�%��F�M9p�{��8Ŷ�����M?%�o�:
����;f����N�ɶ������ �Fs�����$�Y]W�v����;3�jDx�)�z^�-�h�S�ڈ��ﻦT��
�3�J��j�Nlq� �'��Q��$����)iI��� ��\`�4>����g���W �Yv�%�1��r*�]�h.�����TKu�ԍ�
���h���$���C޶?��(U�P��<�^A-��q[K��v$��|�(+dd<�C�}����3UX�|gHT�Z�����z�w��z����I-����>�3dH�9�*� )�{���b��z�K$6���#�a���6�Jd��g��)P4D���0��CrQ{*D_�8F��X�J5���\�k��RX߭���ڕ��H�~0��_fU�$H1�h�i�nI�C<�C�$ܓ�Z�-���˞(��հ&-��~W��@�VX�<�����5V�`M������n�I16s���ea�[��d�ĈSE�%!�NV#��|�� ��3T�!m��;��/L�V�غ(3����]�QF��=��ŀ`�B�h̈��I��M�jl��P�[2}]h_�#."��WK$�+���|!���	�a4I��~��9)��i��|u������T��r��J�ƌ�竑]��0�,�
9�.������J�;O�i����êI�n����F!���$mTR�Q�)�K>��O)l�������OAd]�?yX���܆��y\�4 ӕpA��=�����D,=?���[���<��?*+剧*�����l�����2����G��Hh�E���Վ���'"��:������v�����u���:��i��i�M�16,��m���u�i�iK| T~��%��ֿ�ێq�_��+�WϽ����ۛܧ c1�Z�!���1�@�g�g3lk���Ð^K��p�cn�xx��H^W�u\��N0A�A6�9.�q�Kɿ |�jw����ٺ�� X�{��%��y;4u%e/Ҽ}�������i=��c:}n7�za����6٠Z��UC�J���+N{P�ߝE����g�X���v��^D{y����e�[�|����3�8@��WA'M�D~@#LYl�rq-���h�D<e�,�% ��s��9�Ț9jx�}�|3\zL�.V/3󍼚���a>H]���Ddr!�����q��`3�S��C`���Zkm�a����pT��\���3�F�f��.�9�/�I,qp0J�z��* RQ���e�:S�t{T)p;8#�~�E�0��sfs�y1�a�*?�k��'�.1�����)E�\��B r�s}T4�L���Hp$- ���/������PpG���+�~���}D\k��δ%s�| �q�!0�n�P����{C�L{)�u$���~Ѐ�2��m�(�!�bmZF��<dpxg��OYe���S�ArK
8.
�\l2��tZ�
���6����Ƀ��_�e�b��M�D�e���ఝL�Tn���7λ_�;
�;[i^�{(p�<�p��O�T' p���wx��F]�,tA��f.�X&��0�n@R���m�
S�0>���(nWWk��+y����yf`abFU�8v�Ceb���8�n[�,��u��˸)yo�<0���Y��Y%��4wF[|*\+9�,Nưv��4�Cd�/�"��Q>��"]u�QK^^iʴ�:���*]2���W^�+cؾ��M����gҪ�!�&��LӶ��x��*m1#cp����ӊ���܍.4@β�.b^ ��>��ﰮd��@H����3��H�:L,��d �G3�{���!]n3���otٹ~�$���Y��?�o��{v6��%�u$WN9�( ^wY7��'���l�)�=Q�
:�Mʬ{#��0Qv�	���e��g#��y���V4���tn�_���|�X��I�t6���pzQέ��/ǻ�LK,��3j�۝U���9�]4�(�K������;����Di]t�jK��?Wf�z����x0����V�7��	b~�K']h��,~Xbo8���f���я��P��+����� 9����[�[3�~vr�q۸���Qj��sr�_p�f`������]�<閊���WizY؝|w���J��۫�Dj�ڤ��w�0o5@�|�Y1 �z�$��d��cJ~~���p�"h��s]�a�O�6��Fq�������}�?IE0/!�vL/].tmHᡭ�͆��W��C��Ցs�j ��<Z�wЈ��4G.����(��>GK���Ej^��[�T��	�j�N[���"B� 
�~.Qs�@S�4|�.���{���J�t�9D��|}Tr���8=U�0�!ۗ �pŠ�DI�;�}N�s-�_�����`㕳t�:�|�pI!'F��pNh�ELvt��/���9�E ���$�#�8���<zQ��DM�Es4� ���WX�;���ڑ]�@|竇�����!o���.cs��3�H��n|�]5��>���ỳ,[w^tr-��0�%z.�iC �`�M-?��<�;��ı�����8,���ї/u��4b@&vJ��&x7����}0 k�X�����4���j�ٖs�p�8�F��^w@��ʃ;��	��J�����kR	���o>��0��p`+A'Ҁ��[ %!h�
��UK�%:Z����H(4O��v�ZEڄ�l�N��4�۸wú��8�i]c��|zC��ۂ��]%n"@�>h$@qe�CJ8�>	��?_�Q�ӏaӥնv���QN�J�L	Âƅ3C�
���TuI$O��We�����Z���\v试��5B�K���dȡ�sjL᳨�����!*(���R�9 +?�Ȧs�r� ��s��`�3%K�j}��+���u��ԅ���)���n��U��u��l�>��B�lr����o�Ϧ_gz����W� �����R�\9�u��cިp\��$�I�h�&)����m�M+����^ͺ/-!�@��s2p_��EU��9����)�Z��ߺ�D��]5�~��8gT$IPh7o4�xP�����N��V���c|�]W�͌x� z���K�\nP�H'�M4�ʋI}�]u��7�U~��aS"�J �;�Vb߅s�õ�&�VL479����v�����m�i��x�����^���Ņ�i[�ӏ��f�^�Ov�vt�AB�g����ӷ{J$w酊}���Pz��Ŀ�rϲ�x�q�s�GW��|���D�����1��F����j)���@P��թ5-f]1�O^�Op��9�Y�v�Y6��ʟ�A`6S݀)o�o60κ�!����.�dR���Ƨ�=6���D�(���Ɖ�ep��1��v=�s�z�.���&I$����3!�^���#)MI��Q�	��o�md��{���T,�Ԯ�P���o˽0:"@�ƞL%�&\zV�<��	-sS��M��B �ȒP?���ICSQ1��p))�:G���^ԯ�X�S?K��f�}��-���-��v��0�JYb\�����٥��ۖ2b>�R2$� �!oC�J��zÚ��@Y}��mE0�|S���>T�Iy�iUL

�( ��J��̟�Z��;0��%C���o��2�kF��ٗ�����'c>����x�8{����.�Ԩ��;1�_�%�Q����gl�WFU�;��q����R���t�e�0��q���3��F���FY�\ًG���8��<"�	3Y�#��������܂�B\b���䆃��z��|�GaxٵS��:�_w��2����eU }�`�&LO� ���
r�x�h�k!�W�%�A�Ql-�E��4&˻'CYH���7�����&4h�Sչ�#�o�-�P�5]��nw�Z���h�2AZDb��ԇ8�K�^����>���~xIb�wAɓ]o��D������[G�?H~l�Dm�*��>���rnC+�䔒�C�۫�ҏS�qM�~�r+�"�[z��<��*==+�;u��	���Z�l�?��u4�I����~V�4�Ć���^}��{�`�������b��͋2��4f�R�F���πd�>�oQT��X�mw��u���ҽQo�s���$Ci���r����s��,�iǒ�6�����d�ôyC�ߋ2��9-֔r-�h�6V*)g�ڽQ�e�+��Վ��=������x�Mm��L�_B֜�)
n��Vۨޙ�(,�W�Q�S����P��ԁ�Hq�<j�=�]6p��M�=��X�<��6л�p�g�672h�3i���Db[��"Y�Z.��'��_w�s��I�y�A\t���&55�T_Q�f�v��.�`�8�bs�!D��l__2�Z*��ۑO��C+�I�K$�ƛ�������:3 �[7.EuƢ���~���1�E
��w�2�L��O��Z� j�qc��4%�lӭ�F�����`e�� 7�r���� �̈́�]3���z��Q�pY��|�00�:X8�*{���<��?v��H
�z����a\�x�?d��l�r�rIh5qv¾A�2���d�AY鲤D`����?���l��c"�+q�0����G>�AQ��«��Y��bk�/�H�������CM��7�ρ�
�珧�;^�L����ݱl"Y;u�AB�dT�:�����ȍlh��D�̹�ٸ���p�`��n�w3���Ֆ���G�Ix���"���ፚԚ۶��Nv0��C��R0��ɻ��P��B�O�t��;7\(1��@�`5��_	���� ��rq{��z�w9S@F�؅8�,N��/I,+f�t�{U1�P�z�C�jƩ�N�*bȷ4zk�ڲ��X� ��vZ|�D�Q��Y��vCӲ�m��#D��M�4AדͳY&�Yn҆�z��%�Wj��@��pM�F�ɲl�Ҝ%������ale`�;]�r͎3��ma
?�!�$�G�ժU������閹��,�K�u�b��'�P�s��$�^�^�B	���IoA��K��9	�j��E���l���=�nt�b^�!�ߛ�^q5گ��P�t����]6��m�bf�Mv��)K��:t�r�A��9��kF^tz���"�S������ăEꪮ�X�-��I%��$��J��:�a_*�ۘ��J�߯��3�g^v���b!a�1]r����;^E�aլ4x�h��Ob2Ȍ�U�-�
����a����
�������#.�-3���C�zj���㪇�ڭk1E�:T���B;Cfo��o
|����MԒP�}����\��1���m�9i&�]�q�u]p#�p.T:��I��<��E�	
�D�ZQ��C�r]�`���>�|U��	@�s@��|�w>8�kuEw�@�4ؤ��$6&���rV�wՕ5��=�F:����0�'Zj�I�K�'�<T��]����,���G�}E[f���u~�kÂ�
}b3x��̒�� �4`�F�[n�>�����ڋ������X>�����0��w�� ��}t��:3b�O���<�X�K�������.�L��aJ�����"pU�c�s@6nK1ѡ�d��j\����~���bt�g�D����=d���R�O��,&��4m꼄�������K�!{Ka�J�\-��P�Xx�u�B�P�,7����f鬜�-���/���U(��s!�nVm ���_�eB�Sq9Fj%^�l/_f���A9�^]{�E���V�pc��5ތَ��K����,�1���5g7G��j7Ef��/���[R���t��|6�,�ҷ�<�3����� 1pS������q�=����C����|�,�#�e|g#5���	Ȏ^7Gy�>"Q�jJ`���6[t��J�S�����#�4YZ������^U��p����%�G.o::��-��l��V@[�8%Ǿ�R�m��<�&<��(��%��A���������|�,�;K����H���j�{��]@͈B^��\:�`�QPV@���E.�	�)��
�%+r�,��O�&��G��ό������.Gz�l�jZ�vZjApn}ˋ�g��K�o��,'(�Y��=h�������S�*(M�URp�;���S&�H�	���C-��;l��考�����9)�@Ɉ��h(�e�|�Ƥ}?�y�#�n���e�d���:$
Y�&Rݜ�v	S	�\V�߹�Ǽp��w^:�vq\�3| �`��S^�i(��Nwe��+PѬ�@h �;���}�n�RR>��+>�q0e֡���:2}��Vt7�Uwg������S_� ��e�E�[*%��q���փ�NN�3�&q�"�*B������հ�����By��!?�|LhI��s|���}�M�#^�����xg�T
����S2G8��t�9X����1�o=o�BK�F�j�ө��q�(7�*� g�W���=���n�F��,~-��ߝ��#֧�rg���CZ�������ݩ�Z�B�=��F/�p� �G�А/\���V�2��ֵ��Oh�$�5�Hy�� �v�	=��DW�M�U<#P���9��̊�>���]�$��@����2�'������m�#��/�'��_�4�:��� ��3\�b��8���W��[�Z1��Ǎ���κ)Et:TRi]�I��6j�G ��AX���Z!&leW����ʦ���<)aσI���X}_7	OШC�?8�U�T�:���	��OP�Ġ�N�olѓ�di�'ߝ�����U�f��m6��؜$�Is���z���w�-�NӤ�X��HÚ1�Z��l���4�]��4x��d�i,�3U��I�&S�����U���$�%!�b��l�`�a�;��nз��U�0ˡ-\��0�E�U�G��R�gWV���wZ���)��õ�%�\��Yz<�̅r�������5�M�}(^X������b�y
EH�+6����0����
7l���r�GP����?J����ą��xq6�ׇ��}�%�f�,kO*�ф���D�y'u��4͉s��Gp�j�H�S��iK(�P��a���0]1������R�Օ#�#CTH2,�<[u5�$���uoRr�8:
�D�"/��T��H�@j\�\��Q-�c�Ho+Oz=9wi�#9�� -P����u'��S��%�ɣoS=�|�����Z�% :��>`yZ�
v��_��7�	���y�C�Lp����O]�!I	+5��>6�L��^)�x�������o��DhKHKn
}h��ix���x�tT��8���)e�k#�#�XF|���iL�Ra-��M�yR���j��,Pm���L�ђ�n�g�9A�?���OKC�w�h!O+���Q�	?��u\	��6����Z�r�=�4X�g�����W?�J���B��wζFpɀ�_8_X�(�=qX2�{���8a��jJ�wfr�Xv�t�ъ�D��Ħ;�y�sE}=m$7-����c��k���j�oEM�;{�r����'K����b̘��wt�����H��z-adr /����o�K�v�Ǟ	].2��{��Gݽ�Rt�XG�j%VP�2D9�cy&�M�Q m���;�[h�c�;��,�a�"a��ķ��2�6n1��?&��R�����ɥ�eyj��ѱ8�7���g�B�ݑ������7H�u�S��(����?��f�f�����=�Fh]�rU] .�LH��ny����h�JO<D�W6nc^DI�;$4�f�w�����j2���<�_��&@��G�P5��Wˬ����meN�8\o`�)�B5�g����Y��Q���!��a�b.l
rvf@@P�l���'�w7G�P�)Nfz��i��ۄ�؜3�=������v�݊m����e`���uY���ϼ���mQ��F���C�3�h�?x�[�� �h�vy��ĂF&�W�'W�3��h�H��e��ӽ++�8yx�`o��ؾ�r�&֦�1������*a�5ۂ*|���pZ�ǤO�|�T�A�=�r���( |526�˙��l�[G0��04N���/��"�R��a��Cx��܇C�J_�9";���L:���qp	�w��H{��"K�-���ΑgL��4�0�,��n��b�!8̷.+��¿.�y�mD[��p�8��@�Z�6˰�|��h��4�7��7bw���51 �YD?�AU�/ _0{�
��=��Kef��q��Aoq��� 2JCO�Q7/�F:C�[G`+��	��'�%Ro����l������S1^ȅd�yv��5�<ԍ��=n���eOa�x��Pk�mBw�ɀ���Wfy6}Z��^�`(kG8ݳ&�.��mY8�P�CT4����������fI���i��U�M-9�	c��Ҭ�5�d9���������{x�Mۅ)^�v�B�S���´����� HV6x���q����
iva�v5�澁g� �*�2`n�:�U%�fn�cƖ��h����w'�r����1��,�����l^�"����^A���CXR����6�GÐ��T'�8u��9C��1�*=O�UI��m���ʹ;�N��c��b6��~�u�\9�<v��]:���^ir詀$Pd_��%����.�s�
ݟɈO]�W�� E���[������0E��cĐF*�W`9)d1�D��c��i���W{]���!Zý�(�J�>�ܩ�낑n��3��v��e���?h�h0�Ձ�D[�d�#�O��|�:��!g%�R��P���:lO��VK�w�I)��F�ן�c�$����S*��7�}t>�՗=��b::�7l叽&�7�nBlp��B��+ ����C��P��;��J_
�j�AͰIdG��Œ�Z��GX� �}/"�Y�
�[��)���
ܓ|�3��گ�oڄ}j^xI02��et�1d�4��s.�i�	�(�(���V�����*ؾ�0���5��1��sjK��؁�i3ܮl� ۉ��k���W����2�?"��XV�M�A�C�h�'~�E�Xګnm�a��5��I��:=�1;_>0����㦻[jN�\L�7�A���;݊S�I4�LV^��ޅ?(PS�n�c)�0�� ;I��Be�$0��nq@����RIJs�oDi��^����J8FQh �}�x����� I���<��o�wm����j�.}tZ�]�ʴeH��漤�@�Fq�{YC$�0��R^�T@����*���D�Y�5��7C��f��RS���.3HS䀕<�9�P,��eXu���"]Ú��/��Bw�2�!����!$+�_������P�ST�0J�|�� ��g�]ܴĴ�u�+�Q�̾��uG~F��wkifd�AX�d<�~Ix��"�����ol�����t��э㶊�?�C��p�����,���l��>������h�0Ph����W^��9϶~�~��0�_j�1DVM�hvBF'��aP�^�p�k��Zb��X3Ύ3RchΑ>��w�43�o�Ω,�%:n��Z�D�Qmģ0��56�Z��t%�h�r��$�N4h%Fض+�[PX�t%;^:�]����
V��g7����æj�!�&�V��i�\/��ߦؘl7�	�甋�n���v�8�:ȭ⍀Fe�ˀcR��$Rj�dZ��D�8�N��w�ө7��c@�6�*kC�u<�}'�H4�I�!x����X�-zES~�j�z� �I'��c���<V�R��`��kTA��H�pPwL�â���754�W����� J�f(��k�P�*=:������ǵ�� E=dѣ�t�Od沅�
�cS��8*z�qUs@���J������Rc �O0�p��RI�P4,�)6JM�#�K~��4%�dƓ^��P>�	�b�s��؏�4�t�I�77Ӣ���<�)�D�&ԉ@v ͥX1W=nW��Z��ø>�V:�oQP��wh��ǎS]�W'��bw���]��3	]��(XJ�����5\ѪS�,|���QŔs��M��}A�u���O�<Sz��`��b�.�t�9*L���aԾa�;.�Ӑ�F��.�U�������V:y��y\J��s���z#$��P��p3|�j$��K�Vj �o	�ጡ`�~k��'{�n����s@��a�ӗ�0�$�i�鳆M���%�Vn���tKٴq���G5Ya�*�"�#�
WR�j(o�l�s�:��6i�e֔.�F�s�� �1�ң1�!��N.�ッn�7ʟ,�q�J7�� 4�8��}?��%�=�+�Yy���Oxgd:;q&[6�I��Y�fW�o�)M����$Ec;P(���-�@e��NJ^ٶimJ��η�t���J����]6}�4��^B��=��]PH���J��K���z%'ɯ�ge_���R�8i��p|�e�v���qx�Bxul��.b>q�s���;@u�ɶ�s�%׳�ې{k�
�P"��{�./����R?0^J�u2�L�h�ahm,K�f��}�y,�sَ.�ˍ/��ñ%ḩ��ȼ�/�i~8ݎyvO�,�"Z�lX!f@���sj/�������Ò	�8�9DIqwQ)�6����@�~�nK\�9�C|��;ղ\ҝ%_���_5|�uۉpq��0'�x��,-��47g�cVy����YK!�}�Y.4���`�KK�c�D��FSt�3ۯH!U��;b�')n�y��rע`B�:�{�X%SNW��g��)QUA*;9��&n���c�c`�p�\CWK�Ӆҭ=hNo^[�n��g��ޓ���,TH�R�����oF;'�8~�6��f�����t����kɤs��?|��.���]�K�1�V6le1�%�Sml	��1 ��K� �����W�HL�*�?n� il������H�3jK��,�A�n��܃��Zxv��OK3�H׍�r�x��*�N�&]��o��>�#'$�.��"	YH��(�^�j*~�݈�}�]��0w˩�i"0Z��`���(v��)}+Vy��Zhű��Em�r�i�"$pG�?Wf�x5�Md�=����s��A_Wݠ*���֣?�����fY8u�Q�([���y��g��XA	���˾`�ݴ�S-���8�"����C�.{�p8�ioa��{���]��ڒiEUl&���ƺ���[U�n�,p�h�F�OO���
���Y��(<18������&1{��H�G�t޶�*�d����]�TR^KQY�N��T�}���a�����Yw��')�Vz��� 1�tO�y	^�����e����h=�X��\��k���fPO~-�����6:�:��^��#��!$G��竜u�6D��8���´SPK��9(h������815�P������T�*�hΠt{*�'m� <�͐��ޤ�4a��
zl�]%��dׁҔ�4h�(Ekk�8{F��f���-�d��}������V��L�gp��E���W�����G\q�ʐ���Ҕ0/���>�G�,F'=p�ծe& ��L�7t�]�&�Χ�w�(x'z�N'�6�D9dQ��o3��;� ���g�N���M����No����I�&�8�p�-o��@<w9&��T�࿜)�Y�B��C����	�[�,�-`tAq�N�M�΂mT:Q� k�8^� X�6&%Xl.�s3H�1>r�4��X�Ԥ�[Q�n�uF��q���Kvd�i�S��{�� ~��E�K�*q��繝��˄��UQ�=��b#WN�����+���XF��-u|��W�)補vx!������Zh�Ka��G�n����R}L��3�6���+��]eW��G��hN+_aP�XI)�����L�{�	G@���A��J�1\kT������PӀ�P��@�Hf"���d��`�$��N�Xm�����}�+�a��^-�5ңP���и�?�D�~9kp��_~������(C�'p��v���t2��(��g�g��օ�PCX DD�l鍯�S+�A��OY`�뀐�'Z���z-T�Ʌ��$��#�a����l���L�]�}���U*�0۝�iʄ�X׍n��̅�b?��@m�B��b�Z����\q��k��j�[2ڃ�G�9�|��?l�������<�C�e���(�H@�߰�D���>�F����:�0�'�"�g
�Ϩ�Q��͌m��ɶ|��ͫ�ኊ(�^!>k�T ]��� _�7B��&��)b��L�� ���d =�]�vM>sAҷ�$.��~�&|��;Oh���g�&8�	��׎>�k�R���d��)�H�:�I�wڋԆT��Ք�\�,���0ljoR���ۗO�}䁄<U�"o�|����"j����Csټ����N�����ZV�ː��j=��L*:Y	Z�D��ʑ{/W`TST�ЊҾzG�BN�	\�B��>4Q-���ʿJ�������+��e0;`}(�TgXqw���;I�"EF�"�<��W����-�b���e��'��<�K��\�O� :���@�~=%�QD��x#R^V������|;���A���H.R���V�N;��!y&��6%.�����i��&n+�v�`�@=�N-��j!yY]_�|;Z<���f��:k]�R�����Zp<����f�x��N��S��+e<�d�Q�=��5����AvŦ+��N:�*�L���7a��,���1卬&,:X��V�$H���[bn�	[��.�V����_8�8����M�HX$�P�v�ʤ��h��eqP��i_$�H���>d�7�QEP�1η40��+J��iӓ��	h����8��ėctz����J���:��W��z�o��6s>B��M;ǻ�����b@�(W�V�c+ޓ��mIŶ_]���W7�E-PY
:�.���}ؤ_Hŋ�.O���`w{U���g�og&�Q��N�^q7<�ݧ��Տ=�?��J-�� ܖ��a��I��V�{&t���
m0�ھ�`�73�Z�2���
�����U<�_� ����Z�D*>�(a򓞀H�%�Տ^[I�>9-�K�>r�d!Ni���w"�>�M�B��9Y����s�W�$����<|g3,��^��+��ܼ6r�S�.�?�_ֽ�-�|y���ֺ�>�R�g��6ӕ�ԃ�?���D��Դ��h��;!��l~_'��2��j�[�������ۭ��m�$ x}�jy�.N��&i�6]Q�I��{�K�
�g^�V,��N2������e�L-�2�G���4�>���c���3tbβ��(��x�j�#r�,\����� ��@�@v�=����&�F�L1e�j(x���$R�W�Y�V�䖖��~1����'ػ�c�\�)�*A�8柁0S鞌Ѹ{杯R˷�؏4L��h�{6��$�W�����G�i�p�W�D���g���/CB@G�ev)�����V�o�+N��.4 �H)(�4�Ԙ}�KX���C��
(����CzI���r��K����^ָ������]p� �Zk�e���"��4{#�D�C�ƀ���ɸN�O6���?�$۲c˟����M�͙q7$�kx
�?��7��̱���+]������}/��%��PRF&5��4n�R�S�N�+n��(��ߔ��6�)�|�$v��C=�l�|D`�����04`,D��w"R[h6�P�EZ�A�6_~<��6��{Tu���8���W)[3}Ҫ�ڑF.�y�<Ggڑ��L?�Lټw�e�:�c�D��Wdj�
�'L�8.����� ��Z�$F�ेI�Ԁ�تv֚�H��2�Ha�>zO�}�^���� ��� ! [�$"�rP��t�vg΍���!e�L9�^�X���p�g2�����e�y#Y6��8��U�ǘr�[����c���j�/�/�y��g�À�pI��(��抚�MH�@��id*,պ|/p�m?ӌ�v�m�L�	���OX�k{��9�� b�T��Ԅ;j1�.Y��h ¿R�g�#l5�ރ�5�v@{�^Ż�L�]���4��G���v�KI����b�m�z��<QL)_I*l�D'vA��;x��@Y��|U�]y�s=���f� �g�ᖤPp�t��6�P:lpg�P�W5� Xo����٫�yW�ﵴڍ_r�9pӪ���� ���{�_��X���'P�&�_^�@
+K]T��|Q9'����T�8����'��i蠏�?�{�#�^$[���o�<��͐ �?7�V%���J�!(���GZ�ӊ����O�!�+<�w�:�5E�
���jz0eK8P�9�Q�@X^�՛̡��!����A2�}�gnȽ�5��J�-�/泆��/���h�<8XǄ{Z`��i�Eޮ���~�9yu��k�>�B
3\��#ӢF-��!'
�����7��%`�u�ZCBPu�����E3S"�IA܆��AmK�T�Ʀ���S��uvӸ�$�r���-���%�G��
-ڇ��]��5[��\sų`�K�f�K�~;5@�[������E���<l��]�),v͹3�K��#l�M�\T�X$Х'�Ō.-�N�kV�*�$�RT?T��)�x�̹��P�z� �^��@ðJЁl��:����+�ýC6pC��
�l���H�T
��&���~,���[����(>��+q� �v��$�>���`c�h�h~��7�aԙO����sy�%������6ǰ���"$G��L��~�Bi�倏H����17:΄a�ki �<b��SGa�-Q���>����V�ï�7-�� �$�%���)I��}���$ܕ��y�4���.���Ϳ�����i��œ�zS-���`���-���~&w���}���axD��1���I5��M�\��<s\�/���O���B�ҽ���'D�P�~O�e0i���fƾfㅚ�#�9|'�[|]g��@ў��2ܡ��0���uxWM�DT���o�MRȟ�=��|ʉ�������?"��(;_?���`5��p��N}խ��*[��PU��%W�׻��}ʢidb4�Mjib�9������&�y�Z0��^�D�����$��TMj�ՠ��Q���D���N�/��?<ၜ ��s��+YBnjv�&�4��ys��p��ۀ�3��8��9��Sբ����,Wc}ۅ��@���*Cs��H��)1g`�����&%8Lbm9�(�S�a�Mj� "1��.��?6�� H�wE5M�=�Vn7щO�ʂ��ZR]M���)�����@�>&�I�l���� q�����ɱ���7��覂���.���X0:�]������I�z�[#gH;\�-��*ֽ�Ove5��X]��O?s>1
Bt1m��dVg����%3<Om0��|�0V[��{���S/� @�n�y�Ǧ���u��8�*ׂvҁ�'ꕥf��,�WL������:����D��p��YѷƩi�ϒ����݈v���k��Vy�G�ْϣN���7���|���ݤ����X��Y!�`��4aJ�N����b���8�>	��o����W&K1nDu�s�/�h���J�Ni�ĥ�\X��q
XR�ٔ�j�D��w�>>ey�B>�A���;�B窘�M�;�H�*��.��ؒUg�Ue2L��P��� E��s�ڇs��oR�W�BK���*��E� y ��C��0�ۺ�+�8ж�Z��v)w���-�5ɔ�\ם��9!f��-̬�{JX���kV�Gލ�A���wV�e��-@��I��k�].iڂ��n$Xà	��P�77�����nf�d�)���6�ډO�叐��զv߯��H�F=�WJ v/\�}���ﹶ}����m􀓌K���е�·5S�L��La�H��C���ʥ����+�[2\/��'��Ɩ^n9��Q�FE�|�pVtLD:F̻�{�|h��ʴ��*�T}�"�$�tLޅ�"�2d�hT����4�* ��AݩP��:���7��;K�H�K�:�p�ʊ"�B�?�&֦��қ��sp-|�E~��%��H5������&�ws[��a�\n<m��|��[F��z�����J��r��<u�&˪t���!�����!���M}����@�v��J�Dyp��}�M~��K��ڰ�?����bp�$k���/	k�Ẁ��W�v�(d�Ӌ*��)M +�-O��Tag�{����v�;	�8�}��ى|� |\������ƪ#U��)�uS����֮�Ex�?t�v��?�ɹù�����1q2K��7��r��M���!Q�7}����t�#�l����ίݑE)���¥�;�z�n���5y��"�f쵷&b��d�>?z�@�*��t$
E�_�	���>������;+󦃼�5���G#��Vv�@`�B�펩�C��ў�
D��T�3�,��M�+1���=lE+X��/1�>�v'�ٖ"-����_gL�#����0�/��R������ӓ&o]���r-�9�E&%�Lչ��^-����Z��܎��cW0Nv@9'�68zIi������2К�����3߷�l;H�"�^�p�g��V�Y�7�4�R�3�mi�*��EcQ㣤`x�\@ڣ4�S��WОZ�c��*`���w8f�"`�Zy���;��\���k�y�s���s�x� "CgI�SY��}�$_���a��d;��ڊ4=3�l�4�~'�sA8�����d[Bl�>Y0qښ�_`xA�j�@V�����?Ԉ��I9y'`L������~�7��ҬJ��sx?��r���4��o����SSK?���R�	6�!�r:���MJڔ�YG���p�P�Ǚl3R�ZRa��x]&��O����o��ljn�(P�y#�j�z������r"��_F�cܥ\����IH�m,n�t��;'O<�F)0�4y�F�i�Oy�[m����c+Z|kʵ9h�ʙM�.����ʗ����%��g��,�dP�#��K�Ȋ��,�p�'�̢���5�$�k�(���7d�4�y
�v3l~���7^+:#\[�-V{�aZ���"�5Q����_szm��{��p�!�1��F,`�8}��Љ�<�\�����R#�DsGj֩���fS8���4LLAϼ��o��'���t^�i桕HJ���W���3؊֬����R� -L���o�}(8���D6R+��GYj�#ƕc\�5fO�͕)�T�� �a��$�YN��O&��Mܼ�JWf�?fb��M��H>��+*�UH�*]�DS�'��M��,����h�(�*6��=tL�����d>8�mB�tg G�sɂMJ�*(�M"�?ZOk�[�%#Pa2� ����7Lzy��C"�x��U������@$�%���u%l�����%J-�� v��c����UlV��W ��/
���`}��Ɯ��Kk%�k�q.J�u)�cmN�]Ѭ��E+bvyR6{�{"GB��¤��Bw�	��z"eѤ�Mآt4w�h��"�Q�5E
q�e�Iׄ�~�����f���u�3�_�=�&d��S�@)�g���V3MS^�|��#0����tkN�Qp�8��]k�����B�J2c9n��B>�:HF��@N9�p��ie�/�:O��4�YL�/X�u�^���kK���^eKu�����4@�.�"LN]��и�mh�QIj��&�f�3��/;G���̢���dM�`E�`�«�qT�ǟ*Ӱ�.k���������u>� v� @��Xאh��T"T�`�ܴ��~���]IA"�Yǵ��[ӣ[n�8���j�x�(�,P��52ee䰃��M��4�ț}�7�m�'��|�$�C���lwN ���Ʉ��>�pS9"lkt���vV�EB�6�<:#o�gj�9�vAK��^7|�"�����_������c�I�;uE���d6��h�n��5�ں���?ʫ��q�OA"7𩙇oiFUz��03n�HM�+�h
���U�U��g�h��m�Y3?#��<O_���&�	F��'+1�=MR�%}Һ�c��jY�TLK��71�; Y8�Wm<����N- :�w��|��Ƽ��3I;�H�va#J�J���5�O���a���J�uW*C�~c`�]H���Y�\���+����r���h����x{�.�,Z�V1��դ
$r|���w��ݽB_w���]���3�U���/%-:|/v�2��_��"��!�(���܊0�]��Ty��pe���D�\#
(����S��K�N����d���	w�52�����޽ᗰ�5��i���Z\�w���ʯҊ?
X�k�Gv�s�����ZF��	u�ѹk]����UpL������^�8�T�D�#.k�D�s��~=o�G%7���_A8��Oy�S�7��^V����E�yޙW�6��u�m\�e�D��>Y�6/�rJ�(�`��������b.�_ �R �?'�=�� �-���vۂ�ߟͶ�k�R��z?7v�FuW���_���H� 0�B#jcߘ��t��U����hZ��@�����Fh�=B!�l"��=�9���nFG|u� mմ�Ĭ��fb�@�$�k��&�����" ����ܾ�c�GbC�.�ŎLo썋�܅�*`Ht��7�ٮ3����צ�f�?KA�0R�u{:'=��tz�C0"�;��Ww�U��B�J=�G<v�s�W���f�������f�]3�z�wf&中�W�ğ)y1#�d^����jP9,x�݇C�ct]7*�h��6���$���I�-3��U0�I�`q�ߙ��H�D5�-5�}MY��/N�v�G J�-p�߿��o%U��C��B!��^|���^/��Ԅ�͟��e4�H(d���d��iN���R����wǇh�́<���v�ٻ>���l`υUI�V��ܷ�b�|az��H�ƛ���9��X�Ȑ����/�J	�9r6�0ڟ�B��������T���~�zo��;7A#�2
yR���ȑl|G5��t1t��6]�,�9s�fο��x���&��>��@����|-H�'�$�#�7��ۿ	EG�s�Ќ�m}ڠ������ZJ�L��DUU)��`8?��?�$"���p�^�P��L�^x!:� �-|a��Qq�
���dR�A���X�����]�7T����Htg���i��.�t��MQ;޶�w�Sc���T!b���A��\;��<XB#���.2�Uq�ô��� ꋜ4<���\e`^"U�s��Es��9
���0��^�EI>��pe{�jz��P"���J�`)��������_	���V�o}>!~7�J�\�T�m#�t�3���o�
l�sU�;���. ���F�	���"}�~8�Q���y��Sж�(n�B������p&�9�*� ��#�F�B�$v���%}��� �hy���}�C�o)DR�,ڋ��g���6��b쯜�J���v�E�?J��}N9b~M"dX�#d��H���6��c��Zlȷ
���7�L+�&$J=�U���ζ9��g�޵�}L�b�^{�J��ĉ��x��� 9���c�Yt�Ň�I���KӶ��!׺{�B�5;IZJ��}�H�����q��QL1�=��.�nB��D#��`gj����y�4^�c8뱰$ڼ�vW���at��_^]�D���$=��9�Ia"W��2��5�_�6iYM`)�8Q�ɒk�����l��u���&b	W$'�m(!�.:�t�kxǵ�YS��O��t�����_�;�q����.�@L�a�������w`2�`��-GQ4l`�)�Syn�hq������]i��-�f'��yW���:_�t�@�� ��X�paw��+�*��k�5����y� <ǌ��C読|�6�%��r_R}�3�2���m�V��:�5��c���y? �x�w��/�9ɲ���|�$KYJ�����������ǝ���X�j�H�d�x}�a!A�hU��,4��)LF.nM��� =�ۆA\����o,�˔l��c�#d�L}iLyS+ݔ�p����QOw6�����'=�5��+VE���a.&����}����D�Q������@R�-�P{��Qo3w3��84G�!�{�V�:**���E�����"
�H����V�5W��֊��J��0���mZk`C�t-��;sM��;§�Rr;��r��d��F�*�fﾹ�?>�@;��4������P���
�MW�pp�Sb�7�����W�D8����w�ו8J���!(�ā���ό�A��7Zm��%t�T'�7^�)ql#ƫ�L�WC�_d�L�b����T��<'>���3���~D�����#a�v�*��E&��6t'��|��	������	N0OOϺ���������ӥ:o��J�C�	E��𫚒�Y�?�t�a"�!��������K��4��%�Nu*�K�go�D�,a�谵e��]���j�i�\�? jۚ��M	v��U	��h���r7����|l�6!ɭO��-Z��I�/���-V.�6�2mp�Ң���'%�8���W ��`�R����;l��9u߳�h�Q�2;S�Ν�艤�ݒ�mb�$�,}j���PQ��5���}�N�=�J��H�3u���q~ �vZh�t�	�LNRN�Q�s��&c����Ԋ%�S�)o�q�&jn�0��_9��X=X��Г��ѧǊ�n�s'�u������O���ckh�X�`�������SA�BJ��T������24"���J<UF�@Z����I��x�Æ���)����4�Yx�1w񈣁��M��)�h�Pnk���:Z9�SD�u��Q"gBuT�I~��=�@+�Z�F&<FGF�kE��8�>Mq����E4�M#c���.�EGߧ)-㏾��b�E^���P'?@�n} ��������N!L�6���"�1�i��i���|HgNo� ���|!'�0���v@��u9��A�L�O������`��]u��g����nǸ?q+��i�Gα��7�A0��D*Gs����M4Tz�Ôz����i��s��Mt�s���@<+�l�#��{�^eUwcכ��"�S��w�XwqGb"~�a�����u����9}�ȒC[§�TΛ&a�I�b�sK��;0��0^�69��-�����4# ���r���ŜLR��C��ea�"0ꥐ���R�B�2|Ͼ��F��u#�#)f�,Oc��.�( �w�\�@fr��j�{��.#��ef�s^=��)�u��L)?	\���a��@^ٓ�6H}G�t���E����q����c�Hz���!��/�Zy��A��tcBj?�̽�t��L�/WA˲��\��#KW>�`<doG��<���l�~oZ�b����KX�T&:X�����[�˒��O
�=9_� �7/����c��d'���q����u�^� ����ơ/����孪��V�ޯ)GD|��Ƈ%F�)������W!�q��\[����r>���&�g���bUf}8�>��6�֚ ��8c{���J+5�l��ˢ<�s=2G�f_��R�c��Dן�y�ֹ����(��~C�b��e�~ �ˌx�Zߐ��vow�Gz�.����Ծ8�0|+��9٧c#��{[�
"��4IW%,̻�$���NK��A>�(~�F�#%��k�3����%�p=�u���$Ӯ��cA�<#[Ԋ��w��3֣�/���>��O}�y��ʼNG\���dcF�AyU�n��Ή�m�����]R�8g�a�2aT��O�<��I&�;\��z��v)]�=�|��`��D��E./z?gleg
1mV�B����j���Y3�Vŭ��u�{�@e3�1-��N���\#mX+�z�P�wP:,Yԩ_?��b�@�#na�!�|D�;z����~I����)g�)FPXM�v�=���9M�8���4���Htq���OE��򠝥[s�rDQ9��F���O�encܑj_�q���H6҆�`��ݭ�J�]g�W!�Շ���翤Y�P@�M$�+Ϥ��7t��o��Q�����&}i�A�<�D$�v��uʘoyFO�"�5x�c�h*yeܺI0�\�~p �X�?P�b�M�):�-1i�d('4�����v�*�4g3��K�Сx�^0�f�b���/���g��L1��ro�?}�s��ҍ�C _�����~�B�i�]nZ�j{:�$E��~����(R�ڗzz9�q|��ɧ0�:�+���
e�L�4O�T�*����i�\W������s��J�?x�1��c{�ݰ���B#�x0e���nD��A��b�s�֪�:#x�f�6�B����{)�Vc��FVV̒��FzB!YSiysor�l��o�V-��L6�?u��Nf�V�z��%�l�ɇ% �4%��5m���ʳ٫�]�dǖ�KZ� M�x�5��������e	mAxQV��h�>�.���~.�ە��)��Đ���r"�}������%�q��N��_��0D �>��:��&�sI��Ȱ�#��hյ<F����0,��_�j�d�Һ;�X��W���[hT��
.�T���~�h�h����go5:U�G� ��yi��|Hc�Ȇbl��ى����ء�d:�������=D�N�ߛ�I8�sTHt����n�,�e�.�����Ѱ���e��&��R�+Gš��0(�y�]�Bթc�5@���{p�j�����8��~W�U^Gh	ۡ����A�tq���{�ia/���>Cy��޾��d,�F67��&���'ל�<~=j�b'�?�p����%��t �n�:�q��^[��ҥyO�ΰ�A�� *�e޽�- �����ʅ�Я�"�2�M��#)}�{�Y��[\yWè����m�A?�{����.-�
�\o3H�ܐz-���^��ãx{�꧜�V�'���X���-RQa��k��5������ne���WD4���ȩ�s��慒���!I�KA��͘�w�#��e�J�.�1`x��9�ϖ�<����0ƴ�)��O�v����k'�V���L���T�H�����3���1���ww�J�S��6�s6$|��x&Է���B�
Rq��*~]�̛�P�AQ��]�8�d@$ ������t�������5�CNK�܆A% �������.,�9.����7|vn�E��JQ<Yvv�5F�/j�� 0'��+&��'ʧ�d�N3�+7*�̓���_��><L�I@���m��E�$Iy��W��?(޳�弚"�|t���#�Ro�3*�V�-T]H��і\Q�jr��6�8O����C��3�EF��/�4)ͱ|[q�pw�D}],�P6\�$f�ï�����?���o�h�[�FLh��co��^{R�;vH��?j>�d��],O����_�Y��~��{V�d�f�}q�͓R j1o�fR��Q�c����Ðe�)���G��V���\��D�k_܀ȪZ���K ��H�Q�џ�K$2�C�ߗ�g��kr�J��lD��\^����c(�ة��M��[�H���P��S�ü��\�$����]�����\n�)`�OIc��/A37 �����OwG�@E�j�����k�j�?z���)����'����k n�L�t@�pS��N5q�BH{��f��!}Amh�F`���d4����B=1VQ�kE]˺��n��� �Q��B��˯ ��/�뻱@�?��i���~T���f��g&Iv�Z�.hN�d�'��F��%s�ZK[���������qD���� ^���R��6�����~G��Nh{ow!�Yh�k��J�7O�Nn��ke:FqY��(�����~��gƦ,N�������/l�]n���V�<�����
I�(�l�����4/�nWrF�iU�}3��w�"o��cT�%�#D?6�3���=RP��*�%ʁ��/�ꖖ!O����p�./��`�];���L!K6F����5�..�A@�0u֭���\*
�H˒�+� p��nB#$>�����s��� �'��N�B��S���s4,�G�������FC<��\��#�j��3�S��0Q�dsj��Z�I�	�U���W9mQr��
�_����-Z����!S��J`�ٳ4B8��8���+������
�n��VB�u_nS��O3?I/��&b�3�8�>BW�2���a�l��OX��E�!���		 
��ȶSϗ:���&?�g_�
�4b�\,ּ���|�Ku���*�QDT4B?�i�*K�{���V#����y�eK˲�i�X'�5 fF, L�KX�|P7�����7��L�f\#WR1�tz7�?�]�$*�7�_{�sZ��%t�����d��o�%���}��xv��� �R��|F�Ҷ _��E\�U/e>9������xx��?d�s�VtK��9 !�����_��v����SXs������X��F��ӑ���"�51Ov���6�aۜUY�X9
m���
���Tղ����9��P+H�3�Ԃ)l�FChؐ����]�GC�+b+��/1P�,r
A/u}N!��-��!�tu�oG>F��Mt��	,����4������ui�U�q���|qeMW���>��>�3f�=R/H0��g'���/ˣI��_��.�Q�E��U(ۂ����Ѷ���O��W86�
�d����M;�����q�*r���3Sa���H�۵\���`�9����-����j�|�ߍ��	IaK�*4��78X%�j1	A�K2_��V��%:��a���J�͜$߭��˿����w`h�Y�j7�קِ ������o���?-$��8��_��)Mc�P�#a�#�u2B�6޷�r�BC%�y亀=<
*F롣��	�E�����F� 0'��V��5���Cj`�ڏ�qde��&� ]�m0Gv�����,뭊�����D�e2O�I�����Ba5��Y��2<�M�F�R�yR �����0���MNV����Q`��Ow��p��{�F�E3�۞�atY��g���ms1 ��T��f_�L��^�u0��W~�ci��4+v�ƞr*���k�+mk�,QhI+?����ܱ��_8�����]h˲#��`���G�>s�	M{��`�zԞ;�6�J ��ɟ�C�=�&��[n�v������v�ы���cv@	��_����Df�߱n���"89$I�_�d"��?L!W��!D&�����9��a�"y
;��3�n� ͹;o��9Uz�_����tI8a�
��n�6/�r�*�mz�*���c���@����-�w7�b�'�	�'����#�'�� j�*�M�#vi�:9)��s[�͋��ƮWg����<��d�s|�i����O� H�0��{Н�*��*���
�Nס��"�#ҵg�
S�Iw���]��*߹��|aA�j>�.��,��|����Se�4A4���d�O�	nSw�趖�s��Q�!�� ���M�e� Y���o�����Al��[��ZѢg�J���`��3�/OCH Q��|��6��ƩX��Y$�~��"u��1*	�+�7����!��|.J�=q�79�iQ&}�ʾ�VJ����H��>ƛ3�Õ���۪-0{��κ����F�FrdLa�Ue�Fv��9�@��W;!�]p \C�n��!8�h��P~��G��$	�s�O���-���5����fF��5�Hѿ!5��d��z&��o�P<�z�򶮲����g+�WB�q�ŏ�]g�i���n�1}�Ee����i�iuI�������2�)� pl7��f�S+��\{�:3�rF�Y��1��V��A����׋ϙ}����FԹo1�aDP�qo�>�x\�x���P�ex����>��+�_�)�d��/3f���Xg�cB3P�P{ ����wF"���}Z����%��GD��-���XX�N�Nu�$	�X���E5Y��O�#�D1E�n�����V�{O��k�g
��fq��0dM�BcJ�S'�M�����$t�Hh9�ᓏ��H�L�;�c���������.ζS������7	.ᠭU+P�&���h~�Ҷ��%��ѽ�fM��K���ՙ:_,T�O�H,���
uk%
�ZRB�d'��L��ʵ�q��;!�q��{1�M�ͳx���9�����w��2Օ��y��$�	�x3���iv�.��*r�yyrA��X��(`p6�A�+�����u�Y�^?Ǟ�z���э��I2 l1z%>Z�ֳd�֥�v����-}�r�]�2X�0��6��	�u��%t�E��lP��ٱ���1,��d�3�Z�T �mG>�Y�:aF�|��h�hR�L!D�po���vPr��{P:��p��蒝mTC������m�6��	�4���d���#�ffL���?� w^�:\#&�rf4!���١� O��v�-W"��G�1i��BF�-���@���}�q�YgFyp�J@��1�]��'�d!��vE9���*=������2�2)��m��o-Y�����̠P�Wpr�#�'_���t��-T�]k��G�]JP$%|�❖F�����l9Y ��
�Z if>פ�%R@ =+�������Jl��u�A%^�8�ɯ�"!|A�RF
5�t�G�	���]	E>|���{q�^ Iw&rU[s{S!���!���4������=f�|�+���z3F�h8�a?̵М���Sh��l�|�6�e����%:��L|����2��K��"kI7�,����_�/��~�I��Ӯ��
$�<3/(�Pr�r�h�K�r\�]-^���L  �L��bK���.�W��<Tu��7�9��9��,�UM�:6��;�e��o.�%i��G4L�Nama{F6����r�sp�ԔY:���ս�2������)����5
�IK�=Z�i_����2�8J9�rp�	ZK���=���qNv�s9"_;g㴴����l����;�
WO$i!#��2��DjpY>S"s�9f������a{��Eg�.(́�l7R+˞9��˕%(�
Wا)�F���r�2���Y 9LM�#S��M��� C�D ����y{s�
º��������!?��b��/���4jJ�[vH�I�׌;z�t|��=��:w�����z��0���dr�C� O<�
����mb��re~;C��&1�A��7`�?��j�ſ��2�IF�+4�Ƹ���k�I;]�����dϐ��#@;�����'"��=�t�=V
��0���T��s,ip�b9��� K�=�j>,��Kj�p���LiT��Es*!�>>�̎���C4��A9l ~�m 9���:YĤh����W�_��P�mp|�]�c�&;9�)\������wE5�~�^�I�XxbQ,�0��z�'��HM+ک�o(9^GF
ؾ�>5��ª�+��w�R��zKo{'�d���; ����Y�k���g����,�f��n�49�!\9�?�����_���N�v���9��.|٤���E�3'c+=Q{�-m���R�C�����g#�a�R�[���x�9���*�r�E��=I?�Z������/�0'a�trl)ΝWc�%Q)n��\�D6nN��Sv�}�uP���"�5�]��C?dV�!�=�Rė��.�{�W�'��=�k9p�]�7�4������e��ɻO�DĤW|x�ԖO	�$T0O��z�B�ၿʮ�Fk%rL6��9�C��/�Qh`�i��[�U��㛵j�W1��3�+������� ��uEoc��=W�?}
��z�z��W���	���3&Ȃ��G���uS��n`:�n�#�w~ +N=�7��҆������I�Q����������UW��$��o���t�0K��Եf�/@�Bu$��a2((u9��A(�\�j}iz�
��	�o(.?@��Lc;	�~�������񷪎�չ�O��Fs����{��:�]�	P��[z嵫������\B��㫐��%���`�)hӝ�\������+R�e�6��j<�-�[=m8��v�Ri� ;�n�l�{_Z�l���uE��0KC���֩j]����^4����̱t�s]p$����IfK�qA:��ӌGNM���Lw:� �`�;c��Tμ�9��-v<���ϑ�̵K��V�3�_����ٔfv����\��G�=�����gí�ne�z�~NAո{��^�7(Ĩ&�4�]��N.���PZLZ�#)���<-�0�7�k5lc��f���)��i�X���`[�H5�}U	"	^@N�@�l�X��s4c����*���mo15�Ҙ"��8��g\����S�i��U?=�V�93� �Ke�X�B�Q��X���[~�$n$bI��]��.��ȵ!7�*�'�"�5��_
�M���n�ۜ�V�QW^�oΡb�F=�~?��r;�����!��##�^g8/~n�(?4������n����&���Ə��%E�&���t{=�=��4N���Ng}w�^�*zo����ŝIDv�?h��;[���> ݯDa�����i�P��ݍ�F|�]QMw4�RB�-�$�P=�#��=6�~�y��ʈ%1�A;���mE=�J�%�%�,1��� �U1[L���y�z\��L��6��N�1q��z���F�'�����d+��ہ��fLM!+h��T��H��Q�â!Vqo�&wC�!}��WP����+!�k�)/w�a�~Xh�V7�ힲ������}���r+����z,��ݝ��SH�iA����1�$@�k�f�-�I�޶���p�1+�ВBY	&v��V���,�e����Q3��e�L%��Gƥ7Y����q�!���e��#��{ĴV>m>�� �G�h."D���t����AB�訧�-Z��zڐ>̣���,�����^0O���N=����k��h��A�r)�kT�����YB.��,A�Z!A�Ī"� E�"5�3�� #�g�����Ǎ���Ȁ���Ắ� �����bW:��@�%Z�@sa�"u�;Q^����d���V:��U@�)e)��F�����9�Gh��΃��;�k�V�f��$7�̈́[ ��a�70��{��/��[�&]#����m��W	{D4��F�~���� إe�5�ۡ\ǉC/�Sd��L��
���{e�W0P�_��c��뼒cLa���=�3G�9W�:~�AF�;��h�ѝkJ,����5���i6���o�t�H0]N�����T�yQLއ���D��=e��geI���x)<X�������_V�ٱ^*�\�*桅~�
���:�b�����3��yˌ�ܝN�&��E�W׏6|��)a�>Ef�O����#�|�,�^��eL��Rq�Qe����XHM�t2�V>���
�����h�}��w�A�N�Ҍ�_��KP�m�NPx��H�ξR,6|�`H��+q���<�`��>a�S):��� �/qU��`�D)�G;��)�*�dB0�[��{Ĩ|إ��|�	M�n�kw�9kaiw���U�"S�7rv���a߇úd,�/�R��M]m��:��cБx����2�l�<�H��MU9�5LG�н�m�wq�shu�[O[@�H ��L���i��(c �X8���E/yu��E5�yR�EM�"$!O����	Q�-+�v�m������I(
��rM)W�aX���Ϊ0[����zn���6`S�^���]9��,n}S��8�b�K�KvV���UFUF�W����Tf�x�a����&�ng�
*���ո�O����>fTN������n#i��8�
Z,v7�� �p�q�ɫ_�|dDv�I:N��C��Mx��7}"����:D�鮴��<�j.e<5vGI=��_���Ɲ;v�Q���i:�r��¿�C-r�(-Ej�i����8��t��\J���PP��ϼ_��XTE���2�<�"'��e�5�,_���EW�J�M�����}�P^����l�~�7~J�,h?�q����.��1��s�yٵS*�KlQ̾�BB��a|kw:{��t�F-�E��U|2
�ElD���{�&(�`nz�����;�|�dǲ3���O�a�Bvg��J7RͦC4��e,�z(hWV����[A+e9�2rk�WfӅ2k��l� I�08�U��p�E�����e���j���G���}j�����/�R�%牄�;o��7נ,yK8w�]ۚ7�����^*�_����[�~KS:���v�:�m�4�L7
���Zpe0mŃWJ&�C������!/&ف�G���4L��L�&!����ͩ��o�Y�1(�*��u?%kZ�:�88yͫ�F��)�����Eq��&7�3�6�!�!e� Z
!�b(haoc���6�:���^U���c��Z$�J�A�m�� "��AYQr���d�[t��d��yV���O�c�.�'�1�K񸶋)�]Tb�E��N3N���RB�dnw1Z�a�V�N����E�Q5�f)�t9kl�K~��[d�^P�����
	G_jQ0�'��89]�W�uP�Ȍ����ț��5����]�ԑ������4�4�p+)B=���2�>J��-? �@�l�	�7�l*iD޼X�֙�o}�_Ca�ў��u��W>=d�,���:�D��<}�Q��QT���~��szL+'�Lrip���. -f���Av</��B�qR<j�[���é�Czb�_^=c?�m#r��
��@��]��U{RۼF��fI��NS�ޓ���HGk��n�ܹ-�.8���m���Mw ��.�k5$��v���'�@��]�B���O�Vt�����S`RU^ �{�N����.��i���»FY|kUd��H�a�����H�	��$����G;n���7~�4�R���'�}��K�Bf�g.N)W�G,��쩐�[�(�h����M_	��qZ�;�*�;ڌ��+���T["/>Zk�;��,5���h�x�Nd��΍sZ�s��e�1ȿ��J�%������Rs�\1�$/�nx�(����m�
0G��:+N	��#����?x��Q��L��2�"�dk�\#S d��FR3��h��+=��o!���.�p~��'#<���"�xj	Z8T֠��oC�z��{7h�zֺ}���{�O;ƺ�W�Ғ�rԶ'V�~�>!>���^�s۸�ְ�� �i�J2�����e.��%O�N>�H��^����f70��J���S�T��mj�O]�Ry���^���\4M�s����Α�?�űZ�*�}�ʫ�:�-�9͕ɓj�����q(�:q��;���(+w����`&<��̍]��Sܣ�W�`s�n�i��Qg��,��RDDXA�eh"��Nv��*/�d��kKW1!O���!>_+�G �YA4�?{5�BF� y�d85�f�9LVq,�2�������7EU���:[VRe�3Y!��
P'r���t��|\��u �>]_E>�� ��pe��λ���eR�+�4��z,�5t4d���`����#}��L����ƴ����/��K�a��|��>'D��cM8P?����$A���\����^��-���CcaB��k-�@����K�P�����OL��L:p�����[o��?>k�OD�sk�`��F����Nd�21m6�
��z{�i�yk��	�H����AMI�5���0����z�3�W�:o0�r��e/ri��V&Mn[E\1���!�p_�#�fT5N��~ſ���:���k"��w �A�:c���)�C���w'w�ɂ�nk�8f�����zV?��~��~P���ݓ��['"P�>@��[�dٿ�9k�(hn�U�o{3Z�E.�ҷ '�p�KwS��,�~~�Z�7��7�^"�w�JVs�6t�h�r��j��<�9@q�(��L5mޑ�4Fs�sVW�]���F�c�K��<Q��'* ����/ �\�KR9��:���gb�ݍx���Q���˱�SG�-0���p&>���8���2f���m:��麪rx���+�۾8)9\�n�y?S\���`),83/`�=&�]�o�ʁ:��E��
w�>�T�k���.��)���3
L�DA
�M�g���V"���J��8ӵ��l��۽�N����6}�Dp�ɓ��b�/�o��U��C�L������v;����)���Iv������0�'h�jCs1�8��=�Vv���B��[����Qg;>��L�5ʢ}�@�T9��׬#B�+�r�
�7�nȏW��;�a�&��� �R��9G0������7����%!��m����¾_օk��j~�u�������u�껇��`!��fW��
�Bt^��&����R+�y)�5a��g
�M�+���&�|�bm\��=�ͭ������9$��h�(�� $�|𻯗�"�6�n�h�U~����[��:�a��aj�t��!sm���3�gO�T�6Aq~��f�skZ$�e@�L��t
X?S��iwLMd�4�E�>�@�#)+4�����t���� ��-	��;�r;��4�������P���g[*¡�yJ�@�_�� ��z�d�;J��;Y�!n�B/�b���5�<cξꂈo��{������%�y�N+�Dk���e�Iw�uyH�E��l1`�&]%� K�;�?�����Mʸ�#�BG:S5�ыZ/�`�a���#㐝�7R��*�WZ����x�Ҷ-)���^���0�d+γ���!�ƙ��#��'�4;`n��Z�f��/讀1�1!k��=�����&؇-�{f[!6�]����i�o��$Ӻ���w�;7ը�Ubn���͗a�uU7����N�ٯ��
N��0\wx�����XF���h���An&���ߑ��������K.&���Y;��TE����tˋ�!�%NЬ�����E[H��}��c{T�u��Q��u�˹_S�F��#GN�l��#�e�=��87V[�"��Ad��,N�{q$@��Ԙ�Q֠��P*��aD�h���ϛ�l�f�,��;?���]����i���}�5������aj�s/*(�����t�3B��<��Na�3t��1a�	H�����R���IsR�hgΕ�kc�e�'�'�� .��FY�d�~����F����q�/�i���#����\���y��%��Q�p	�ㄠ�ջ���#)�/��w��e��G�M�`S���(�3l���� A���ࠔפ
��=*�q�y�R%��������VEµ��h��R�'�-̵�S5��l����!ac�&���u1��5l�7(L���?kyQ4i�:���_\O�~�:L�QF��-�����U�MN��.��ʥ̡�����F�L�������0\Z��1��Z���^7�|q�Ykϸ�����1�d�8Ş�6$b�G�/��6b_�c���W���4�������V zP���O��h8��f���:��,fW�x4�]��̸5���Vb�,����L��>z��c������%�,yd{[b	�(��	F�SG,�Ε�}�+��G�R�&��BM���K��,F� ��u1kެ��=c��e�c�1?�q��� -nAm>}��$���?u�t���Lz:^�Mo����y����[�s�d���s��?h8g:�
v�yK>�/��#�=�~��G#��[;4,ԛ�W��:k�e%.�1��S��tx������Ƶc!6dq�lV<dI���D���3Zk��O��� ��T��G�~'M~�_��%�%��O����#�=WEN�йŹ_�7uyz�9��F�#tj��2���3����R���#�����Z���t���!��]9=�
st]ހ�t^g������*�d{�o��]f4��*����y*���ǠN�վ�b�@�N`�ھM�؍���`|h��Javf�|�!TD�2�j�	@rKc��W� ��Y�&^W�(T"�-d�����B��Z�Y;R�u�^^�K`5�/##p�մ>����׈G)�XK�Mx�r![�tJ���[!rLac�W@H�-�D��I7O$�����S971��dV�|R�R�X���z
}S}61#�$ȩOP��D�6A3���Z-���L�g<���u�r��J0N>�Ӝ�pس�,#�*2h&�Y���w�~=�E����Q �bb$Y��L�f@~#�s
zx� ��9�q� H�"gi(��b}��ɵ�	������*��Ü��і���WOG{f�$0.�@�i*�v����"R�m�N=̆h�>=���:���ilZ�,\���f�-�����3�!�u#��ص���I��1bR-N3��A��W ڻ��Ix>���,�<�/��+F �g;�D�q��+g� ˷,�f�c�qF��\�Pv�]���M�X>����z'o�Ʀ�4��~d$0u�㺳�鱆��L�|̎��th0Y#�C�KZ���
��aJ��Ve4S�[��3�x�,9�tn�CqY���H�k��y�KU�]+Ua�/MS%�i�����yg���T����������گb8�i��b�K�S;#�J
���+`Z�T���w]!_) �\���%�{@�h���:Γٕ0K�=�_J���Z3Pb�4�����O�����,����+����f:�p���2x}�ՌO�G��X�uz�~�Z���<��H��>��w�.<\T���֎�;]���k�}Z��$�l�0ר�Ck�mN�_�񭂒3v���djwO	����E\�Z����G���2#vºB%�6V�{Y��dH
{����|#��I>��^Щ�N�v!�d��)q��<jm[�M!�%Ll�{@�/PL�P��^� �s\������0��_��#9ƻ�ˈ���r�ɹ��Ї��/�"H4��ז��8��
y�M��GWځ9���Jad��T�"�>��W� ����H��M��O��.����U�~JA��`O >��b����oU��E�ҭ�u�ѩ�ޖ��Y�,tod�ϱR(5���t��ר�
w����֮#d/i���ч}v�s�|r��deU�1(�m��]����*�����8�C��Oc~��mL�J�\m��o���	��-���Z{c�+X������;.��������p,�"ێF��8D�:����"cy��Y�_K���~�m1��L_�����4@.r��ץ�꽔7���ZGuT:D�s��7��Rz�*��oOT�P}����ˊ�-_��%׮#A���lA��ۤ%,n�SK7��Kd�^m�:��GnDI���!�m={�rXvmy9��zy1,�"(T�l6ƶg�LE���g�����~Ѿ9F55t�Ka�|��-B����l��׷Y���W'�0Ս-�?/�ˉ��:�|��a���������F��E�[�"z���#�Xq��{vN�@��s'h�A�͕<��R9�a�IAv���J��<�Oh�s�N�Ή%��޹K��Nb���ښL��2��T=&5(��B�b�0W�u�����H�����aT���D�&xlS%�� ��6*�p~�xd���N�BRt� 'VrK�#TU"@�w�,���
 ��s�4Kڟ0��f�bc��lv�X�8?�Bs�zjd��jW��ɾ_eNSl�n�ՙ�J6(i(�"x?��]���<�#���X��_y6�Q�2��3�ɻ�Cmd�.ܭz�8nd5��_��T,��`͹,�fY� ��)<Z�����&���3�&?�ea�tcP��Ck2��}|��ϖK���,*�~oY�� ߘ�,Ԍ��?���v�n�
�K���|�Rs9JpN^lJ��x3����&;��4�w�Wk���\��o�)����O�A������p;�p����1��e+,�ɪ��AȤ��J�Dv0�X".���,HzX]RV!B�R$���)Os=��W9?c����u2d&��I��L�����Q�f��:/�ʱz�d'
S��hVLR�d�����[��o��,f�7�y��9���m
�;|�9����][p�q�*������U���.@�ΜLd��}���ʄ$���?k�6e<�
�-��J��M9IDX^��h��iF��<74��8�@r`�s���3����m4!�\�z��X���-��'2㛕(���X��]�����3G�:幜th�&�p�G��!�A�����d�W��9�~.��d���.�#gZ�R$[:��?D��O���胞Y�DL�wա�ቩ��L�A�ȶ"�H��T�%$\���o��E+�?����RQ�<&�֐�OI�e ���=��A���.���Q�CqS�jo��8�:y~�a7�7�NsRّ��\~�W��>�g���Y�>>��90��͢��x5g5%�gz*���D�k ʟ6@d�_E<���Sh���.���J�m8l���`�$�$��r&�O$��Lj�5C#ɽ`w.�^�K&�e��c�c�sSj�T�c��LVg�3x�ȗ��S��!LU��X��:ȩ ��%��^�c�!�צ��#���pG��E������ۦ�P��
ۛ�(��b�6�y�I�*�
�Ɯ��iً�n��7�א�B��c5?Iù;?0��ysT�/�=��C<Մ}��K!��8�cxߥF(���ۥVN�s�����JUR:��LȝE�Pg-qY �0�2���%�	h�4Qיֹ���J?��2Nt�ߑ4Oa�)�\�iF����;fxs�Iz��H�����uv�v�oZ��k̝+�p��V�;�F������a9{���^���������t�����.�ӗ�AAf�Ѓ�?�����枝�K�"lp�鮭> 7�ݗ���0�I�rl��|�s���N��B�ÕK�'j=a�GFH�JA���_j�O)!��ŷVo~���.�|��5����V���C=I�L�����Ʌ]��n����s�թ�9�������Z5�@�H:��6.ZS��^��!���X�3�t�t��w�B��v`��,I��ןԤr�b^I������~�����{��@���g�3Nyk���k�����l+q��H	��
��oa�����_`3����.��z��*ty,�\���i�#G��L��:�r=��}W�G�Q�K
~�$sE5Ywm�#`�wNz4C��d*d���@XH�J_�/.:K'����Rt�2�Oj-�j[��#{	uv"Oh����#>��%_ImZ�E���;��}N#���X��6h<ny0LO��C�z��J����5�Do�]l��=A�?9瀜`�s��r��n<GW��z�����ʹ	R9}Et\�-o7#�����;̮��;AS�9�5^�7��&(4$�yc����2����k�D��0��H���E���8����ޓ}o/��@m%���i��Ҕ�ފe8�4'r��L[�[���J!|&�ڙ=�Y���XA�pz��#�w������4�D���@�u���� �����7�*<�'7ir+�� ���>�r�������M�km�=�;*��4��v�U,9(ԃ�G�K+;9��$?G�$K��i�>�ڰ� 4ff$��^�%J�ðE��s8ԓ������LN���K�i/f}��̗���օ|�*��2X��4����jܹsj�E8�w�۸4�0ʄ;����~�R^��=�������b�n���?����GG@�+��hg��4AaJ��.�s"���g)�ԣ2�F���=�m�Y���̨��֖����DF5���:�,dyÇ�iK�������Mi�\_��/0'���4���Y W�3$y��ۇZ+����
9�����/�����0�0�לx���mf�Jk���E�u�lN�I����8l�Q{[ؽ�av��fl���ʥ�����]⁇b�iud��=k��DZ���K�� l��~��l�9��e��*�9���c�s��b�޲H�;C��X���9�_~��5V�N���$�������ooǔ!�-Q�=�-���?J�(Kq0]�F��P�+����n���h<F�:�b�Y�#����3C�Dt�g2ºk���>���n��U��Z؈�O�A]��O��\!�������Ӹ+�#,�=s�ڷ�5�.eJ���"���� SWpb���ᨴ��;�z�LN���"�c�3#	2{CJw�*�O��^�Й�5��j@��J	���T'�6��=+��C��}�2e~�JYC�f=y����h�υ�M0i�&	�;�����aD�OiH���2��B�i�UJ
+�Ԩ֬��:~��u���-�������#�G4��Ro-�$�a9���i!���	�ߡ�wn���K��Q7�Μ�ۀ���i�:����E8�L^c:ML&�i��G�_�_����/��:�����k.y��
�;R�V��i�����x�"P$/���REu��q$�� b"�2$%�~���U_A���/�%�.�9f��q�G�pm����c���܅k�P��s��N&��a!j6��oTl�"�q��)�F�"K�P��?�hj�9v�.��m��w���*�fh�QҍVS1zov��&
e��4H�tM��- ��ЖV�#r��s� ⌖c�[������͊go�⃨#C!Ά���}��U���i����5\pLh�c�m�J�B�u�rl���Б�h�����d��Yݪr<�9/���Cqp�0�Ч��b��� D����]V�/pm��U��ϫ�(�C��Ț<��C���Lfx���x��a�g2tK&�{�zA^9�^�.�s���mT��]VDl�޴�ԧ?`�s��V:M���$dݛ���m�Y�o���*�^"�2��gƾrz��-���Eה��zM��"��̬���+�^�R��ME%oex A�/D�4		�EN�B�'�:r�F��&�y*ܟC>g��ѻ�,<�L�	@ʙ������M4)r�m�ҁ�F�M_MfŵN�����{{�O�Zz�c> M_>SA���
���i�\��i?���DS����i����p�H.�k��R�ԸԒ���2,v���V)A�V�ZlO8�Wq	�@�Y���!�X31b���`V�U��#̀i�|cC�f�V=�f�f�P�f�]�M��x��tj�R%�����U��p<�pL����.	�����T������S�/�������B�C��a�=�gx1硳,��s��{�����b�����Tk����4��7��}z1m~�3R�q�.2����İ���~BR��YS�6�c�U?/�wem64�%�v~��~!y�/{��(���u2U!�'�R5�_Қj���l���`���g��;�B~��zH�/_\=]�U8ӣ��u1��I��I�i���_�D�Э
TuuV½�s��_Q��i�/rF��Y)��~�4Î	���y���������}!�W�L�ҳ�]��F5�+�wg��*mp�(Zb�*l�1��ӟ:2wŔ�i����l9�.��d����.��5���No+����8PP�zN�D}��L,���(��̧Ǳ���������ذ��!�M�=sI�8�̛��Ò�'
	l��?������v���ɻ�c&�$J�f$j1���İ����3��[s�Mn��}���E���T�?�4V�sv�����Jw�����$@?��
�Y�F�5ZJRa���_l�o��1���#G&�7tps�>z��ԐpP�.���]�"�m"�`*���1 ����_�i��C;���&f�0و�5�p���Z��m��5Tٗc��.�Qʄ�2�~�o������0PL��y�Cj	%����@��5]�E� (=1��9ޗ����� �u�v\+��t��8:����=ea�M��U��>���4�����wc�]zV�w�ȏ-xg���
���d1�c���Y�H>j$��ܮ ���+���Wo4⦝Xpz���:y|4�����񱝛����B��R�3Ԏ�ar*���B����ҮԎ!
*P*��O8����Ǳ)�i�]G���V��)GP*vŐ��= ֬���\�T�H��͟]?�`�VB;�wƾ�,�i7d��@�n����vJ7�US����`����%T<e��'�e��� ~�5�����"���r`ǀ�Ռ�xw1>����"!�Y�|#��p��Fi$�H"'|U?��#���k3G'����_�$j���9m�Dz��=���k�U���&��Y>��j�'&	M�p�����գ$=f�G���:z�7���]�#)]�����\����jȐ���j�b�\2
��_�
���_e��1s*0���Ok�]?��	�a䊽]-������V��ZÜHf�&�1��o��5;�!�
:t��/� ˥&�J�%G�|�8�<ӨX�pL=�mD�-g&�29!�]�=d�����d�Q�U���Y�����6׾5�r�O�����DÔ���g��R�F:�؆J��%�LX-;��0��߮@�H�#��=���~�e�k:)�Ǆ��!�@���Qt�}��;8����L���.T'�)�����5~5��,�?��l'�WR���k�T������ڞ�V�zF�#fF�
F��c��j18ug\�q�7'�o�������:�G�\�w�*�o~�(5�D�϶��T"�<c��H��l�A��bl�!z�a1�_�y��<���Y Q���p�4X/�PS�Y��U�[@�G���E��q�Rj'���/��P�WS"��d6އ���A����F�N��Ɍ�}u�dF:�y�R���,Õҋ&B�ZH�	��/<m�$�J��BڜF������p��}�`��y�˅[��7R2�: ��7��0T��W���4�;��!�Kl'�\*ZcK�����y^�ʱ�V��O�i�2��{�8qT���fjѪ�L���80��C�Z=���pō�TR�1g���UK�?����J^�β�����x.��}��U�����p$;qJa�[�Qy���A쐭��}����T���.�N�ƥ�>˭�_Y5EI!SĢ�F8g��̜ �Pc˂v��(C2g�`*�q���ښ�:���s�w"֧���װ�1�XU�IR��+��u�G��D=����(RY0� �c��>3�M�hH�q�79a�=����I�bl},�����8ouE զȹ���n�5{"��ou�5W�r̋p�XbN@݂u�4tX��h5��3հ�f���fל��5�v��v!FFr��!Q�א+F�YNO��������/�:��4 ���a�����RZz)��Qd�z{9���Z�Uj3����{5nN<w̷���f�S$�=���V�F؋~[q@9�ê���tJ�u��2R;1�1]���� ��Fk�8�ce�[�G2��<1�ϝ�X�a>8���z��D���=���$���d���w�w�\J��tk�%W�J�j��Z�q�}�	���Z'�yw��ef��7w��XIS�J�_�%�}VgA���a�����k�ٹ�}�DЛG� ��w*��f�x��N�P�r�c�m!�7�CH�g*yO�Ȅ
�&S�?-��Rk~��]�K��#R�F��n��Խl�by���\pjJE7�G�L�,:O�k�bg ȋ�Ql��-'�u"��C7۫F��>\3�[ٿm��d� 6y$A�#s{tu� �q+�q���	>Q��3��e����j���0�Q0uxs�G�]����A��f(��yK� OF愶�v�Ś� �6�1KI��dxt���46/�Wj @�䝨�u�NC�s���ȟ7�!�!�����E����-[s��&~_�p�������Ѿ��.���U�Qc�nfr�����ol�!�Aw�����+�S�#���$�9�� ԏIj� <��piLiV�p����9�D��/c�ª��j�*�m�"'���l��P�_�p��*�M �_7��ظf��8��T6N�;3�9s��cd��]�BJ!*o�r4��+[�N��.a���Hěn�΅�[qdJ�-��c��g�-]lB�� ���S�h�I�agU��	A:MI��R�'^�� d@��3�z�~*�0�u���w}�*gRZ!��q^�mB�Q�0���e��s8b���8������j1H��r �a���{�;���
�E&�����̖���Ytw!���86jdO�͕C�����9ߪ9뷒:y�@��A�\���[��60U�x!ez.A��*��L��-b�D8wY�jQ��Otɣ�E���.���z?�_����
��:����a��X��b_[�&>a�v6Ffp+W�.,M�U|
\��Z!NbA����=�ݘ�<x��݀}�V�����3���ݻ�ZIe�#��s[�|ZGm�z;�}� �>�j�ل��<Y4�8gn���G[�	:�2��4$i�B�P� �Q�PN#5���,]�	da�	�ҋ�z?�r�Fec呭Cy"���&е���T`��l>���h}>9�KS�|�ѹ��r�����VF�uCɅe��pu5ښR�Y�������ss��1�)_�4��R�_l�Q�m#:T�O�.>Ę�&�������5=�䆟��u�@oGc�̃V84|�����x����O�C���4���s�=r:�5gS�Sͮ�|m	���&.��mc�(i�z+_��՘�I�tl�[���?��h��؊O�