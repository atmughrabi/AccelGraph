// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cMIcigtO8aHgwz6PmfHAA/2R8qsEWEtu7b29/QLv12VgQ5YJ3pkqUE/VNa01XnW3
M8WzbajcLliUad/kRhAa7BKxESlkOyhx/U5z05K8I4tlgQ9jT5oIueBjuxLsLWF8
ZtlUWCdc5jihDiW1ItjGSbEZ80iMkGT0GQF6Q/UaMEI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29232)
IFpkQXYc7mHWtKOWlD27wPTeYh/3Cx4vdRtOBsOFIblICxjFtWMtOezlTN+A+Fsc
4R1VzgINGVM0ta3r+k0GWx0Q+pIRy/kscHelOmWVPU+qX2iwrOLCYpj9U1IArrCD
nTppjk8b2RntNhDKyM/aXdqiZ7zu3dr/Tr7YvbW/hKekcGsrmv6IEs2Kx1yJitvf
Onsdbx6yxv1BnbSOj5vzuGWACvMya17XkxEFCLq2XcnUNs7fqkcZNzVzc7sin/er
P2pa8IjwOvaHb3FjEIOCMEjzOXWD9G92Jhzwzu727nVCRs4RYqGEEhcXN5IOgVg7
xjXLRKAjZJWcmFF9oakkKfG/VzbJqJlRTUoDvtJuhLQ4wj8fW18RCXk95F0bwmFN
3PqwES1MiV3pUKse2hS7YHSbocqBkbnYatleKHlcTxjdXVvO0FP1gnAASD80mr2L
4i5mAh1FZxMY3gdq00qVMCzTdsygEBYng/xBstCjF6kZsb5kXclKJ7DskBOCs2CH
KhZ/052+Czkfw6O8+lAiglhJQk157ACx0z90Rzr7LARI+xgHVGKL+8fgGx4KsCjU
gVlMFZ1kB7iOywlfByNpoQX1XFS3bIvMcXq9LTcAOrUUUFRuGN8OsN8c3Wz0KVqW
X8GhhxzI8TwV5+52lAIjQpBo32gw078X0iR5f/3YtguvJI46gXuQfqg/vm15RF6d
pYpH92/pyQFiNZOrKD3vqDoPWr+1WwY6BCiB3xcdm8tzzN2kWcQP9hnCINHHf655
Oa9RrndrQk6FmtaIa9NN2dfXRfMOO6KvSCYehSh+J+vSjPdww5fBiBfV5rM3+j1Q
FkynaURNiQyvsUFzQhIqq96mDpkp18W7qA4w1CN3dYKfizfyqyDruAhtCpyHJ/Df
KagXmsuyRYwXQRuHtWlc0y/deXi00TBNV7kL6hiAnrJnZVLzdaRPIMwaaAlDwnE2
f0UAqyk8Koo0b+CCl9ZVkjZJhr8OtD0bH/HiRI81quBqEmI4aEIVYl0G/1S4AMWS
F5nPD+wVioitZQ4c2y7bRslxJyPLerD6NFeMlpb37B/6S9++Pi1BUYJhOsHZH/+n
F7c4u4yTpwJtLln4DuAcm5wgIhrflblMDw/T2Y5/hG+FgEPsT+UA3AU3pOBrhCgX
n111f4iQ5Zn1e5Gtb7sCtrfinGgD7fo8TeIoIERp+FutiZfhmmZc14zCkvVzZEs4
5U/RbHby0igBQweHChg9f/GS9X6z/KDitpcOFBI/0jPp+LjdkdF/wTYLV/jlWtM/
v0QfNaqNU69ye4ZxMVt2Z/amgoXeCFXe9JpZjEG24Hc/qiBDC7p9kAXa6A7UrcYj
OUFoVysAeHXIwKNp0lQ7BT+ifrWpjTSeZkohE0hiKbSSdHHBNr4hNEXMo0wvY3wS
rzzMb2DVFyUXyZ2gF/VCddH2TdByVGNlkG5Gt873S9PBJxDuIfZpSr0pHOtYE12E
4V87x8up0mzIy9u5AKgiUM/ScchtndqqIHjRPzYYcErouMu6SJj4VVhUXQ5Y0fdX
lR1G8VTNLCRawbX+QeZQbc12Xx2kzRX2bculhn39ydwy0/gcpc9yl5R0esut1OpM
TV1bQdoOdsVO7chb8YwRIjPnxJ5AhQESpemHig0qfWpsGgyId7G153JTgZ1MCGqr
ptpOIxXPNwvTHYfIekj1VbcEu5yKVqjjNL2F/SUJec8K098MxVX9D4Oc1KnaRGqH
sBtBaPXEjr6SD81Kow2hX8om4Zq/lZF6u0OyRQeSsOUVBpwxf/EnwwXrxHwjyeCp
PmErlpP6KELl52m0BWqXNdkW0AkGlMBtUiOYbvEO+XkW7AfWptjhxrWn6VvsmyMN
Yl7/CyqsWGVNNkiUWqGcKt8pP0Ek3bN0cMNP8LYR3WWPTYGev7pVI9SNz+6Lze7x
Z+U6dVxg64ALPAPEC7mW+phLFK1abq8zCQLGcJ9ZHeAeGepPH7ZrowY4wrSnDfvB
7ryVWybe1JQj0tXUe5N0G1BudW/5u59Ruoh+pfbujRE0ZEjMbjOIexB6RAFB5eBR
TB1OSYXD+PJtQLGLmj9z+lMcrjmUYtKNRpQPB2jFZHIURQF5jF9rJ+RTWpRBT0xO
qDpu9PJpGIbMr8trdSw9wtCA6VWWJg/sPApr6CoB+9r3B/AWWVh5AoiRdkDo4DvA
v3EFFc4V9KabOzWV4YBRPtgyj7X34Zk/gsWt6dT73CWJbSyC5wYPPtjIkwGlh48x
Aij4btmK7AtcG7DQ25QnXcxV+3sINspVn/cMkCDf9Rj0Row+Ds17NESpft0gGxNa
Hg2zGkaZ1e3utD+kTPfEc2lkYPm2l4VV1XGzMF9DhWiKQNmrh7zHMODC5B+l1Lmc
Be3eO+JGe7bm7e/FB90hyWd2NhKvtNMBsyLBAEYeVXFayZ/GUOlcJEGhrGKFfytq
osocihljWgZf7fj894XThMbsZUR/muzCEhSw9dxoEoIbiLzBCytGRGBrfXbTR2yn
HNCfKJHIsEvOFsOUjI6Yiw67Qg9/+HYtUyFvVAXZcGc3T3E1jKI/nfUbqlwt//H+
FzjaS69noxpDIdI1q9q5lr5o9VOxWCU4nSIN8hTIvg/Gi3WMdlFnJp6CPnrdiSCw
GULplSuJo6HAlMa1MH4dNm08elv8LPvUrh+PSB1T47NDPEdT0Ki03BBv20V5wQXX
onByokb7WqnvNm6hs2q0r1FnsLRMKTUYgVUXPxacPTwUQ/eGOIiEBmxQUQYdqCCq
YYH1nKNNpuRrFbBSu/FBkR5l4LaJ0LVjVG1219SH/soWZUfNvyTvhekgLdUrisBJ
0cJGav/ttRhy4HGOqNTlaaIC5r7TlK8nfjgF0Zu/vvWq/lG70Mn8mC3osPhg0Hbu
2PDZQ/CPsRDotFmBMjn1COPVS1+NyNTpvZt0jsmPa/hrh90VggqsEbi3foTygvSP
f6nVIw668nFVlFdAqUcqDPh12ERtjOZrKx7jhWxpyzBN1JNReAQl0oikezHMH5Dz
r84HXWVbYxVUSJpJbBGiaYHGXuSEhdXnCR+eFGK0uxHX/ahjZCkpTB7S1gT+u4+e
PFj5LIbFIDqJlGE+dqDq3QMCQl7+qdb2nJG+RU3yPD0aJpmVscK0dwGUMFsCyuNW
EWwQONRytlcMRZF9d1oUO9U4zXKE/tYgxmURem+H8+ATlTelDcEG3tQSIyfwlggx
quXw8wHOXxRBw57By3jE9KcCuwS0EUFZ8evCp9hjDckzDnDa5V+iM+RgxA7/OXSW
9Q6MfzAT/SUKg/Cmk/UB3KrZvLVZrOWL9pKcQQUELKsswr6KpbDzulvK1m0RZJmG
/YsYzJchdkuSXttUOGjuYhgyTMNW+1T+vxh2gVvCGIIIjSX3Y5sMVxBhyWmqhONt
jsX9WdJvEzGgX/9prQOl/dVlbFwbalQC9cW72fbMHEoH0O7zkV+vkJ3mg0w61sUn
K2FTWijAdhU861wUOZBOCP2RUq5V+uut4TEeJIqrJc5ukuyuqXdF5FHVQj0rYly7
snMX/r2g+Cl47E6i27WULOTbcGRW9/BFZI7pFcTbqFJTzERon72OpEFu7smJEnwP
eutRfis8pCWvrAtZskbcOFCcphsWRex8r2YHr0e2Sx0T6kj5/L5eOXeB1sU8AnCr
SwiwCcf6QrubAK2Z7IX9uQXLwJwiaAaviYjQC7ifpFiCKk2QfN2NZwK9hPfoiLq/
VJqlLsU83hRirXzdpWjT5vgxcIuIHolSWNF6WyMcdjtmlLLFWxTTyVoc3hCr7xQZ
E61CHFIUJTuSJvK+/nv5dqDwpRzgM63DUOkJtFpObMCGJujkX8vZko34MkCkJxAW
Mf1jrXOrX0tJcXXJQmPLxczh2kGIdzSGi5vHab85GrsrIlzYiSMyFhf9o19fncsB
6V+fb8mqXLu1qry5ZNJwT36WWlv7LiuNaMUJNs85vnTri7fr7Z5ZgYoPykdZa13g
Nsq1sCPdDxGj8Kfq/CNfxvFrE+hRSTSa7ir3LOsIYrmU0gFRlLGnuoQushJmaXuB
YhO1HNPzxw5QXlyTq7j8Y9frpE0VrKC7PZWSDTwy1b4kF0xKt7Cer6RAd/ErkFR5
pDNjj1REo7aaSsscOospvy88CiphiC6PYwSXOCuPtSPB+A+/9YV/6rJQ+hKmxj1n
lNYD/XcQ6w3yNEyNo7pycJDg3SukDb0mR03ZZXMhKKUTzfRctJkZ7/079HE7I4Ec
NTUigJeWj/5vB2TKzZHcepU2ZqMCz0Y/qzv/HjEv0Qcw2xxxdBhHkFqPzzC8hH4T
yzEczrjimNFV/iPLdaAfP2/z+A5F9e6UHm7Ag1uipfLHkaSmewBO57dzS5WscqK8
QUA7LqRgPS898YNmYUx+O7y71HKu/BCcn9vvQHq7m7XANq5UpA9vhgt9SZ7IIPSv
twfUCnfvyzFrSJo5UPd/RlT/vqjknft4chL4zX8kGpriJxVr+9YrvTg0dsBowJz/
5tIJSDOTWk2iDPZ7ERNUKyBXzTT48dDBitTqjToU23AtEXeOwLtH5g2/0FpmYBNn
sCMGZY9/pNWCUam22rN1aA5e5YyqGjxnZMDhG2C+8Dr+kU6nP5OxIuwfy+W22eGT
Jirh00vl5xqdsrB3bBVOIpLPp14IQpzk80OBpA2VU1ot0582JlLQOWDtS0Kw990Q
1AjBpPPjQwN+9tTEk2/+ORsKlCiwiqFiAUVcwmkc+K/CxwPFtqKoAkygEqf9CRPh
xucCYqjr+xVFzUmKUwXVoMLtxJ09HoruSiMbVHsBpVgwbcneaf3+D+G5vZiH+JCd
Er8qOcbZ7TRR6Ve2i44l/ffNGpGDQ0D97S72cwm6Iai4VSHcWeYwG/Iofpn6eTRF
BhztEK3uQnnoEwKH2khhIuNM/FE6LhR4hJQj+lk95MmtWBqMVQDpXb5mFEyv2u2w
jTxa14M0t582wg6PODJS2L21sMigeAjLAFuR1wO7F9ERpaokc7CqHnhDRk1vQKK5
R28DpJzO96O2yAE6c7WmaFos50RMCdInMU1hyt7LH2UtRLThe7mkUPboLCFA3c8M
+if5vzJJa0XP64g75AXQO90gDZFd81OeuYo5nEWlBTeM0S92fhQ9c6qzuz9uSjZo
85p/3+JWzsTXnjwjGBqJ6x/VPgMZlh3ad9+C6N5Nl4DOAcRwiXOEZ6xo0ldc6Pmm
EIoyKmMKz3U+P+ClK87848sOZdQJBwKSIL5uSWhSDQbbLMcCiGmHpTifGXEfpuqp
prwvraft4+YCwLIk+nhmo0OlaNoIJIcHTcGH0Y0l8QfbrrWc+dD0gpxByMkOgt/c
EraeX1ApqrhROIFZmWOJL+hiTD2VKbSOXo3Ik1WhrMPc9hN8bkd/+L22ySsBcwv3
qhfUvSzl7whz24VegGJTzgXneL9NRsRR92VyCT241aVcsbyyD5HnIErc+7/DYIHy
qhPW+kn5QE5sz6ukurY8y5HP7aWmUAbVR5oFKHxQkQ2dm8fnc/V06sbUt2yyEaMQ
dt+nRtVVUG1dhnYgHRN+B8e/9C/cA55IwcnlxhvPmETOdGiCyGqZw1V+KgVqWayi
DlvTg+8Ifm5Z+zyJF7Vq9oyy1GJzjoUf0PCY6QAZJWLJd3gN6lQDHlq3qPiYQrF4
YduqVZ4ZhnZNGZjHaldMdWFlVwvdVdcotvqQLl9VdemN1Np9Dxr/zd4Gl+LkpzQ5
1QkbrhHfWSeDHjPDWtHzVy6eB/YCdD3X+OjlHWmM/h20riYkQ+Twor+i8Ddeegkm
sAAg8uAgagcvqaIhxluvBn+n7Y9sMbnjy/HwpIH4nV9rAIUy3MecH3zpJgeFypQf
Lq+xbyPcfslU5uN86hltJUcIoBfW5n4rqKXk1FvMVYyYtNPuIUCuo3/oapX3vaYJ
OhEj99v9pYmol2zIc0YbfYQDIVY6RuNyU9E6h5+6L7YB7Icj4sr2tsMxJRlK+BZ0
CZiyszAjpIKVnjLMAyhfYzofmHKLF5aXIe07Mmv+4KAwRddNuGqLuNyvFHTPioEa
QNAeb+0TFXqERkrgJk5ZprnQykVQy1yxLLanipieou+RDMSkvVC7QC7UtiUtzAid
sZhntnMv71WM8KgjZhP6l4cTWJicQAnUcLTeKoTfqapYDU9Kk2d+tNQzOafUyY8d
jzMdK8PNysCG3iWpPvSDoEyr/Bel8QzI/+0mr+E9AXWHwP0pSjw9OVsAYBiGFGgV
mfeQKQxj5azgH5vb+IY74yc23Ne+gpa6tVDVUna5g4QP9SE6n4FPYrG0fRMtNGIN
sbqqwptl16A/khgIYnsWt6gq0LLIoOiheEb9gFxviQoMQP0ZpWud1sODmCvrawj3
pNCI59ozvODvGRSArZumrPeXqpAcFzk2L4RLPcauh2JmRmz7aKb6h/QouytDToCx
nDQf/VkKOGlKsOTIXij4CNesueFGFXTT+3eYWQRTzJ4PBHKxT3P8yfIO/SVbeEUU
UOyAVEKkWJFxDEgj2WhXEJu+TD0LCj1TGPNofHDVKeUeM/ApUfwxd5a32s76Vy3T
5tZqS9/p/bMBR/cYbkUl3/9niJ3OSvBzRhqNcm4XNkkNJCj3aE4tq50LKH4HwCNn
lb4eOS+vEf/61LvAJLZUXM/zmhDBOv4hCwEkoUsargs+4h9axWZ04BEGg90tFK+5
9eXEqJ5dLVOlU7dV/SbkjMg+m2HIjtArh7HzhsBOmBuHrfbcktthIFJsmpFemNnj
dIbcAdfaqZ2u0kLS2KBALhS7d5Pyg4X0i/tFlV0w0XchmbjR44826/8Li7kkS/ed
hyCEgwBrUo+NCbG8maJHNO3awZVx5q1HnQgtIjEZCd/C3vOslbQCwt6Uj7N5TjLx
7e4We5Emgkn4c2awMJDpKZTy6+xcDbXowHVPjJcp6JPT2ccp2jVvEVmX/TjF27oQ
T6f8yh4JEpUdcY/Kc4VzETaLFMWgYOHUKPWiGdImVtGhucK3+Hf3aXUQKG1qMvjz
ZBgZ+1nvyhCk+c/bG4Pz8mxOc0avI9gg7ACdQA+1KdIpFRV0oyOx8Amz3QtP7+/R
7nKcd11sR8c0zR4W4zSk2JKAs8Vz69X8PT+weQQt5BFn47MSVs26v4UgBXRZSu3R
8G2z5XmsleZkL8pqttBruC0p6QkR1/UhB5ru3CUjdhlFGOWQC+POv3wKrc5JfapN
MMMzy36gdKSTRx9LJxpgGcbAEQ8OHRfUbI/uQl+kO3DVdj31O9/S2/r9VBEtciMh
jbxpPhRgoUFMdf067rS5keMndzOPjU+28ABC4qIxRhuT0vN8wkEf3JI7VruPUUe/
uhkSfy1MKSOntiZQj0F1aqAmJKcOkfheVlHgU7hdRO8o/iEoMIT7uN50h8Rg2Ok+
QWFemhpkh4vJuyzGkHqPiCD6xDhMHuI4ZK2hF9sn+xJ8zcrU1hJEdmCIlSpMrmk4
sFVcoBjrmGOUthKkIWCwj6l8/G78h1tFaCZgkdGNdnaHsYNBB60IbA8/m9oqA2aY
WQG5m9v0+zM4oC/HdkHTkcdFUJ825csGJXmPL1INSahiZ9p+0CXC1Deoj856WCMw
ff3Zo1nx4Ib17LqkeVfuFn2o/BIezhbWAPwT/BOMphKqBFL4CrDaDNgb8vZyxqF3
0i1zmUj7CljK6QFRNINDh7IfinuQHtEG+4s1waKst0RZfDAoV2SvCO2/i/2aapNk
lTRNpQ9ge/NU+xB82xdd8THGDOEJSblBBjvCecf6khmEBi1ftIBlZhAIpIYnWk0V
yChld8Qad9ay6LCLdhooP9xsF+gLACc6ATReILbqN+QDXuAb2/NaaeTDtsyX8g/0
R5b8JDxFBJI10zCGlQZndxUlCzlKK6dI8WJMdsrW4qeTa63jWx6v04j1eQTsM6xK
tFSNpKICuDTQlJKwAj2s2FChrqukCUdh1F4fU94QVMOyYgWBPL/Ker53kRfBf+7K
vec9m6a/MVkOkVPoFws2SXcgqWqwjxjtJZqPEzPss3hACnSPkWKWJmP3n8PnoYsy
ZT3SnUL1fLZnLNiZgVM3H7CrnGiXIrNxmuz7WHfuq9JYU8jvdGr3l1LWleWuUCwO
G/cF9+CeReYSXhKxdR2wvnjd0ZmQf4YupfJxhVl2ca06eBvC01Sd0EppJIQIMuts
HWDcXTbYP7PsxqCto3F7Kqm9FcFVGqq7JP1NL0xQbb20iEcjnBAsqPu1vKoMirid
ncPJt3UMB1GDjwsRuxnzA3yKT3zDmQ72xBtTzYRWj9IOme/2YM56AF6tz4bz35OZ
J6JvjU5e808pqH8M8S/P/5V8TOJoQUzesDmV/rYW0b6Lw+UMaYDrmlEaGlRRImJw
W8Dk8aL8pw5SsB7Eh6GxSVbFYVMZ3sze3HRopf1GdyAWZRD0yeMwgDra0mXWo4Qz
KiBqQgfli9ftqmi0tRBIAJbdwFM50v0yIT9LfQ+jgkbFaGhVw+IVS+R6KCVbfN/N
ErggbTvPYKYSntFoQBTQMLMhYGan8PWSSApX9BL5/aySq75L7uoM7zfH9enoonN4
TquWkQUIDpKmCd/KofphyQKFt/vcbhPXbw9LxbHoIvtG+YSw5XzQXzEmkfpGgJOm
O3zvnDTjvv063J9Iv48q3o2GgSif3G+yccylIXYN340J/iQFVj9VLE8XFTN+SVwE
W0xJ7GpHk9kvC0oPumiP+V5Qd0j7XwrBc/sYL2E80/+rroRIiOizw8Wah0X6ERpU
3JLfN8FGH7IaRen0hpSbmfnhsFBPVZY+sU8KooTZ5N4yU7kEv2v80r4HOUAhRrrM
MBSf1Z+t/G2cfSoC+SpVgCex+apZ0DKkxMQ4w2LOQRXvVbd1J/shc3gnRcXm4wg/
Ro43E/doWQyGa/lcpNFiy4uq+/abBqXtW/MGJxLa5KApXg6vR8R4pT/spb7JVPwU
Rl5lPk+5BtdViV/qEXOYL24aB5XhyLp69jRaF20eH9Yz5RJB8j+3qocWtiSvJDcE
nwP4d4vOwxmYjigaHK6lAbOMOls/F7rrxXTJFj7q0UabKfcfod+faKN3eCWcFnrA
PwrzrwMdCEhtXYv4ncN2n8/jKcEIq3Q/G+ijMqqYTAGx/93RjD2TjR1Wi92Vpcqa
GZ3rX+jhL0jKfrZqTQqMs5G0G3xOIeYAvU7dKLyb+RyzgxUfiPoxSkmCGLWM0XZe
aOeQcgSwRCFoN7eXzKXAiYsHRn3bIP+C40V9GaZjuiQc4AWNgRs1WTkIVYXgxhtn
4LE0j4Yn5+88emwu/LmIQG543yp14kaAX2ljnlLcm+RiMYknWQNt6U5dtulEK+yE
1xlUVYiC+crUSP0cqEENj7/URbvVpt5nGiPlilSRSx/1/fco6AyXErjER6Xc72HS
JA6tFfG2kotN92ge/CMiHb9d1MROmSjT0bs5V06IzbT3btZ0OylGiNTyPnAUlwfv
LV12IY25ztquMSoTRxZSYw8+bBXxd/xaScnKMC7zpWqg2ZHmvjX6FVa2GPfqjfVG
hmn3yX3wUW2onpRnATLqFOYSiwMcAiqq5fKRtSMtAhbMCw1h5MimTfily397Khmh
zh98MIT0vcR63UePtyVh/STxuaUUgBAuHUyp9zMNoatjbh1roSTiI9HwJVA469qu
P9nc7sop/j4k+nqS/PfuxUsjoipqJplVJUCNUYV1n12zsNkJbTQfaf2gYTpx2J9O
TjOOjqGIxmjdTauufCNpBEU26t1b0akdEEkt5ZZw6fNZAABZ0ob3YjeMdt8gGoyI
RwUl5ocd5UUABe5iLLj8/JHQmFaLlzfuFyf/vPF72gjtzuUsOdmmK85ae45koDG8
rMo3HG5OgLju/tekIixKw6mMpa5H9SjalZUSX4mTwG7gXur1KWTrO7JuuT/aEqMR
xerzsthR53nIbkBFA1BYCx9W22dHxSSIiZ7I33F03K5RuO47Wae2yp4Vvv5zYYx3
wOZjuj2ffQI5UaO6M/cL3hTdmkdC3biZE/sx43e5SZbGqMmXYQz+hIXuKYxGztBK
c5s4/Q6pMxeKCwEdMOC0eRPqJxA1zjYK/2Ol/awwMTc3TWNH5y50BtjG9/A86MJC
8MhKJAfOtQcikUjmFjskq0RCmKgN+YdUEUC2vsjao0ZVAgaQEi4tFK1TC89lz/rl
4Uf5S6WkKuetXd52WeTb10fzIlYL5ES4nNOTJN6kDZGBXO6/642s1yvXCrw+HDvz
Ce7nGBaiA0TXmiYgcGKwMsPWEjrrltnBdm3BgIp80SJnrtGsa6qXr2SJaypd5UzL
RmgSb60j1OqkrKTYO9SflrfeM5PqlbYWT8gdVixRn6tpcSVQcXOJKXT+HI28Ys7N
v37dAjlkM9OECUxenYZrmaVA7lLSgP+RO3NcAgNngfb3kvGhc/HQVxEmo3cM/g+a
yVvca3A2xG9CgoxcDVv1WHhEK5zRD0zrQIZwLXM1rxSZ/j2IKGlfYyHaTDQ27MzQ
DDVM3anEqG6zC8PLNAxAS/poMj7KoVG8tydVicYa+a61qvqXzhdaPK9wXtVUiuTR
f7WvRmM5ZMu/GKYq9EubLHg6DhkjIemnkcSM87IvsUvBWIrf5+u1oCvCxrCvDBs5
R0APp9f8KxXE+gaUc4kKt5TEbXOEEtl0Eyvi3nl5HnLBAK8THz0oU+/KpVmqdu3v
o4IGGBO/iBQlEED0/OUzzAdNohBWjvT9e51jVyzQ6znqSuKD0zyjSXqUyo5m8srH
/4GatwjDoHOCn3IhVmrOy8+VI49C0NWuu61XIl690lvzA4axBLFnv9N/NxhNz18G
6LhRY2rYIcEKgYRWnoZ+iFlC72Ew2dJw3Wm4e4j8JDx6XA8TwW23AudenDIbd14V
EXCYomiefAcL4aiKyokRlqfm4wM9NtGWIOLGG7CLlihd23AxA3AcYRtII5wqr/wt
PSp+HNxV5PFt2KqR62xtMoy3T9uQLcLAYiibhwa/oBoaVmJ+3u+btNTneVbicmBt
gBHU9AlyiCjy0BtB0tf3Lg8ucbMF2Ux3Ka2Aupe5WZWyWVBb0+AamuigtirEyX/v
/jZISKyvs/I40xP/M2t0c8khObwhRNFfPHMRDfaDPhKNNffHI3f+AR3uMYOLnLPt
V784gSwUBV9q6BSijLGGS292e7WoOxJ59xW7MVmhGuYYGw7P1DDg3z/do/0lNaDx
hj2mjAYu9717ubGDJOp4OjvFCGZFmuH3u2IqT2biTg7i85SoH1tna+kBIR9d9Eed
X1hPFUQc+/V5J6PS2v44IB42XUY9hsn2bu3/V+pDEOzlwmARAc5ypIp5yXgpL/P9
DG7AZAkiRlZMVe1bDaSAASB3q8iD/9J0czpNneVURotAjWzp9y1nHtmmj2r2OFRe
rbaNSKqEjb24wu4HTAbgT1K8TY5ByGpqABc+oWnbXuk2BEp30C3teEmFCTRlRZnS
XOdxeBqYaIwBzGqZU5ExTfdYOlLTmZlWaCN72km5wRnug/LZdssXeXL5CCDmHvxn
P61fAWEe29b8JVuA3ZjwbKmtiBzamP220we5Rmfrtipl/iXYrp6xomohrw62TPIz
1lhmcZADBSEgZpc3hA1mbW3zV85rvd7EMghCz1GOe/y0wEu2U/sRNgN20GVKApA6
wQ8dpn1OVuEYXTPJbq4zbXrdSIAIWH0V0QqMNLCByU98xZdNe3OcdAruhuoSQiJo
Bf3hdOztGvF2+6Dvtt+s38sKr4Jq70nwLdN0NdYlHdFx3sh+ijJLKhJFBQCvKGw6
ozU41gzfpsxz7+hpr4UoE95IKBxZTNhLzhVed8lpSTxbZd9ZmYJGfgfq8CEvmkcX
fng37X36UHcVeeyTfB1n/bqTVJ4XXJ8iTPG1+C7I0z7MI6gFz753JX4UYVmMjsVF
gtEbZJvki/73o3vkbxJqHe0lbcRr0Jia5Qn7VmQOZ0bbz7HexSZ2SXQ4MWVA1g0b
ck9sokKvg3TegIsBTVFmLRtHZ6k4hog5PLOmjXMk+zeTuND8g+3qLKrsAWHnpiDh
FYcapaqHleDQXICOu2ahqepvZflyt4uolAKNySZ93fN7zeROJPK3iKCxyiaB/p3j
FRLyd3QS30ydQAY4wk2Zdo2hjtWjRXicSN9w3fOC42xZ7uA1V16p93YBWCxR3ywp
5YE6V+g/9SIE+vHTE9s7/N0p5R/qOxif6pFZ7mgF7Xy58z/wp+1rFOG9SyQw671S
XS7CJ2+2HzRroWwZBz9MWuvw5gUvRJxylpbm89hlvfvpQ2pgNhnDtRIDj5Zuhx+D
4h7Uxh9M/L00RHj3lAPGzL86E2DuMx7NJ7xQiuHqYPOl33F8PA84xsALfgbuNMG2
7VsidPLpkn5GcOeklD/ZeNbkag07Py0TKNnNCkhwdm9y/yMcvqHr2sd8SRZpCRYm
g0VjrwTwdsTnnWX94jfRLBgkQXdPjdvpJysulAJH0t4AmtjXXuOhJ5232PXHjXqF
xE6toybDqTmWlYAth7IK1D9+l0OEmOiYaCmfMjt0gTdpEqez+hiom8Edzb1y/4JE
ic1VL6SFT0fPhRvBe4jhBjKH7wSKT3JZhCSUTF8IBXWQfxKdBQWd+XUxa8keCSAV
d+TiIADuSF+t5PA27N6lsKSFa2nIuX0ICICre03xvuiSd+IkqcLysxSur6Cq+8gg
NytJfh4CZfDq6EY6oucaDKB+GQFT21evrVKTHWBU+ImfwKpLXd190p0YhhDdKjhh
ZRlIytyZTIY53GTujgoNaX/3I9Wg+BRYwy7iNukWO4z1hW7z8xNuWIxfiWShjwik
MPy0zNzRHSwqKGnMNHiZzyegAHDNLWdcaMWPL8GaKdaljIcHWFfXWReuY6zvZnd/
EwrqbNfkkeorHqUnd/JEtsXiFCcOXjuLgZU2x4TnOpge1jvwqPrSyzuLXLfydGzg
w+3jsIi/8kbWZ84Cj3C6J0cj42dz3BZqGB8siWUC0rOK+QZDYU7d3WIEYwgWvM29
q04/sRQ7WrC0KZsS3VndZ4yoIctIFAb0t/xYRkcClPRaOqW/Fw6+sPUIPc9xFgnH
iSOWGZJDwVzrIhXADBYP65H8opmNL7hAdux+zOdxaZFpwn0n+uzl7JkgXzAv1Ddi
wBQMmidtYX2zfaFha7+viTISC+a+KZkiI/vMCAi88636bP0dDUqOEZVwieLL9Zx4
7pdZX1e5My6zKpWhSLCSmxfwf8br1JNXw7Eg3jt9cqg6oSvbHq4ZhES0shtppcdy
a4PNDe2vwaCKCiPe/LxIfA22NimUTJlCY0668OrsikuTShonoTGqHETkWoOo1ZCB
hIQF8XWq++eYZeFTq6Mr7QGDhJFSE2A352ramy86dz/UJkA5d3WIERmvNXyVCLKS
vFJkaYA+WUqoK6aZith5RV9nVPf+wt6OeUHk5k7XQFtfNT5oUOTFgMI+K5JhvvHb
i92CfVGx2/2vpcXl4Ojm36nIaxgkU+/rrYxnNfURAtkKezkFUKF7X8uORcKnPJSO
Wr7fCErPWNAKlYAvJR8xL8SqlxjTeocztAGMxzqh5bEZcYnWqFNRXwX/2xCXnhUt
Rl64xcsh91hOkkh29dK1n7JPnNhMUSDFJkGVWByjhP9Lwpa1WhUW/UWZAo+c0h18
hv83Cflexde20usVC/F0H7l8xyoDRWPe89Ed9RDCksIPPDqaeW4mW6cImR7P0LbQ
1Zkz6t6L2RScd+dirAFE3swqFY4P9tQ3gNDWZHRiz3QMnje5b1nSypq9EZoAxxkX
NHFXbh6YAG4WRl4ydUKTUvhU1qFCs1HKVOqQe45PczHNUbGCxHOwZNhSNSIDowfs
UZo0R4cXYkLc1DnEVBJXN7tzph6L772kJTaFhxcWwKAfqi/UuCktP1W/ZpKt2UMI
HQ2wESy1l5MYdhfN72kOsQCls1AXCRlB1A8So3ZpAO80ltgGsnP3WWeWUUYFevF5
fxF87pB44WVNITZhbrkddsZVKdoM+YYK0fxnZB7aSJgvr6FPZE4Rl9/WV98B6DOv
sleSOBkcuE1i4ly1dI37P5IO8UOBcTDjuqZmpK7QsnJ8aAWf/QHsixX6s4x3faq4
lsGRy+Lsa6RI6137QB4yTr8Zog42FAhUSzEioBBHlCwCAqfLS/u+nz1jphMxBQ2l
r8VorQLv/vpjphYdOb7s5pVRiHarmYLkNMNpToj8JvF5yQnqXuBuw6i87so48Uwy
RQYOX0iPrtCHHiBhmDHFfwAih7Q+FcwgwciVGi+UZCAZvsbBMcyvmd0O1U5b2DKj
cVcf2y8I+WoEVxrwfyELCVqoeeaop/EO0cNl4mSKSnrEXHhZxlblny1WPvd25A5a
yPkcrRQuktdCYZuB998ENQixYJQWFaBlGmP8VPiw3hErA6dGMEQ4DtJttcG/dM+T
pGykMilo16RUdVwg5tCFGcQsbX5j75lSdO8ispytnlS9bV+iBlHs4w4EGpY6kjT2
HW/UNFbEwIZ1BC8pK5h6hcDdH5kkwiGCI39l0Xl8no+oqMgOHmJSWg2waNuoKZAJ
cUHTBqJlvkAOdAwc+sWlMIJDhX2898QbDRC/+Ny1hG1NgjFumKpSDGKiZAWt3pEG
VuZNysHn2WbIzgLJ30IAtDf5PQPVTUQwsl0ZMtkdCQoIrDLF8GSfjPLimYE94wjC
dLh89cK1sXJTDXsXU05ZrAkvp5d84EzXxJ7VoTByvHEL+0M6zW6sE/uvDXPCJSE3
jzfvBUFBjUeVDmY8z3vzxp75Pzc57rtJXDT/03Ek5Z5RUW+inh2RUfuHs8zqgbRz
BvYZb7cqwLXGrrFwLFvMyHlINDZgaRRFSthmSitbgfOPRO/gbp4LztLvM6hUP0Uk
xB1NbCIZyX0Ca7/Q+cJv3XqM/AebJmkkPOcHfxPnSeYvn313bqehC7dh9xrkrzOa
kN6uoKlFr24elg7bcwGifPmLTHTu/xRzqBpY3Rc/Nc9Y6CuNmktuA9AEAmjS9Gj5
9RnFNOWnCrnzoy+U6nQLiiN+is1LJAGQrSSKMA2tlcIKIa6MPI0VQMmPmydKEfoK
ma5JyDmxAR0UTqcXCLuxrwsCZKBgEOZ/dilAh6NRwDBsRIIYtl0GLIEZLz7eVdAe
vO2iSRtm0vxRvoXaWydqbFnDfe9kp1tIDxwsLIom35csZeG1Nyh5cIOPTM8/0fcb
aJQR8V8uaOVaD9qarSUc8LN6fGQSUMQQUzK62RPIvt3nlWQVioDwX2/uM1MWq63+
QKtR0eAXGGhJo8N7qf6Wkf75e6hMiraM2atGkSwY2C5Snk5Fdz09gz3D+G99U2QX
dGIr7grZ57teTS4JoNXO+xToW1ItZt/eMsq6unE3u/szwYO0Txm0/sjvTr7xiQ36
nz+GzGgC8PFcjjY+BeIEyvsc5oAbspAG+OXOzU9tlWYXJpjP9yU2xYY6G9yScNs6
6nT9SGXFT2JFYWjO9FyBreMSwQ0OOf/1EcHaZc86gOSvKreDl9vLuwa+m8mIzncW
culmNuukBPgtSfdZlRC+VMdaTyWqzvsNMXcpX3Sc0t0nEV+Oapvq00ZTeXrhUIRz
VQNWUAq2ed0ciMhHEKJ2whSw9Wp1BJz8b/IJ1N6/uxYcT7H8a9hKq75ekjKt6eVy
qI1+9wmevsqxxKNiLsIw+Lt9MBmZAzVBpKNQmUJ5vqXQwIFndWyDixWWlgas4jdk
Lacq+NnGuFYasIyofcr9nhsDsSVCtr0p6FugKYEYfONel9gxqSKmYRcseWI6/Emy
fOqTQMC1xheqvVylX4xnF6J14jHadd7X4wAcsRJlka0X/a9aguzSswlpthPuDKJ7
c+qnjKKkFDjh/zCiX1AwG3NwT21HZBkBzA3aKwbcU3MpmTOcONbhJKce551rcstz
L8RfEwPRIpYNtuZUGOMRF10GzOR0Q5ZlWSsjRw8xtQPLniTI8U1cYKQfkWYm4030
bh1kR47Mr/8qIBKuUy1y4AdRT6gtYu8HHREZdNuRod6dlNK0RolfPOa6EuqwVbHb
vLV3V5ewuiQRv5Fls1P+dzHUDM4J7u02AvkqN4X0dcoQqYYHvLZpdYtGRlE1vS0R
M8tY/5TI2Gyi6Tx/rTNW43dSBYOjCsgITg/1pDqy1as7YfeLBBGzLAUGfh6j7RiR
83ORc/QM3OziyhSWvpdNIvQTYFqGy7ruDT5wxi4jHG+a/HNK8gyV8wcpuCyTHJI4
1vbxc8riUGJ0A5WIuWMtQbiK1hCFqBTo8TM97MpXJcPfUif8iIqIW60CKm5HzXTW
uU7AJdYXXn5rbruwIn+Y3r+v1FYeufCWZqeIp8VGehaw4qvRd6BgMDkM22sySRUg
VgXJ/kHCf6EpfqDAwlT+HNz1RW0KO3EeRVfaVKZQvbPmT+L4ef8qWMs69HU/iOSL
5+gmB5/Q9b2UBmvBXeyqlu6Pj+EkwuOnmjpFl72FoM8kcJ/iyaAZW+JZXNTrkZN9
ChiQ397+2xGxisAkmNXGgUnxRP5VQ8StSHF17FNY/s4rtbhblaG+M7WH2wOv2R6P
frH1GFXMIGD8vsv5O/R/6LN0abYnBKRPn21cqHLowHOPhN6STHEkE8sWRsDWlVnu
+bIkyndEMsIouC2uPJ/dhVHXu8au5JVArKAq2Vxclb7yVGLyFiZn07VuNWWn7e1M
Wff/I0qfX8OUQpjptyN3dHUSMCD5Rkj7k3Ej+lpSC87qI/mmrP+H9UPgRPTVNbWS
DJEBIbuihLRMfy4Sz6E0qrb4zqtYcD+liiMBP0kg84aRNeehu6y1n1EpwguptfGk
NtbLuQNItTnUnMZXHBzrDbGvpDyJ8iNyyX1euvS57t3QGwvo3PztGaJ7OU2KRNGQ
hngIpwJuGKjCKAEkoE0gKdoBMwjhil1QyuyM/pcRo2UdcdWgh60fRbp6toYkEqVw
yRU2zqSZAy4vsTKGYNhdX4b9N2gwLf6YUjUtQY55mNLzbVC/rRH4sRvlI3Ix/CRe
3SCH4brra5X1CWbCb1uVjR+5AZAxit0fEd8OrMwDDq0nOpPlxERBAnyyUxubDHLj
7yC66Dt8XZwvOBh8y6GZzQnRxx64Z1nN+Bon6w3HTyMRhRxAHjLAhZbWXHBZ0fMf
WdP5QSpdwZmo2PUt5t+oLJz6E6Arfg5hpcgXasmizf5nDCug95EnH7XxKVWae5ss
GiQOuMNKBaESzEBOFB2cBOp1a2tPixTSwE7TbSHurPcSTUO5ZPYgQJJJVlgL0rs4
wQ5+CZv0Yf3izdSyf1VLubSZAwmU/TJhu6k7Xss8SnFbwrfrL4P5FTXErZpGQceC
pWXYESdwsF4Q2tI41XtCxw85C4oZg9YrnTOrJSRww1cwEWETNXOkUEcD+UcuMLnR
twB6x3XIuYkBgJ2Glh5k6eefGy2Y5tylC3Skf7hP4NoJ5ZsvDFgg6BrYTpdBReb+
SweGRmVvjPCd4EPgemkF1GxCse7hVjuuKX2hkUQzSo4wIBU7o7Vtl+oPk2IDBQV5
zF3qVU8LrG+XHXAEPfVaWi5l3QKN+4RMXAmj1/R4JOH8U5inLOsFctiOi9PgALKv
wy6E1XV/C1R86Z+l7SZvQPF24sab6nWYvwU42FPiPpmeLM3VznzskMFuisMFBLf3
+tms8c1wUH2uSYob7oyxRP0k27UyA6vfsRptBqM1O0MSTF9QWX5JkSO39By6z9Os
dq1fFkO4Kh4t6IHUNGLLJQGJ1iE5QgHp8eddSATgx83Hm4wyPrS85vT5SCMTm+mz
59WdeuVAsLwVNt9FfLwkuvuWFNjETDmVm9K5GOjBuugqo4z9+qpPKm3WaiPO0Z2+
iET8jY+DBM7lgRblKFU5JDvlbsgTmmSYy8R6nXSWHWZ4pmU7LR71mLp8qytUDJcJ
SJZebC4UD2HfEIHqr9Xgg3+Aka1bGz3MVsnEa0Glm3BSFNiWJmsD4tOnk64H/Czv
4Eh0q7fqJpuav2oR9yzlXdfI++8b7HkTd3O9LJLICwJBxs7+KDknuACl82uKjNUs
K1uf4JGNgydgwg0AAvQUoUKVi5qf2QpeHWd75Efk4CVrLaxqtjWJ04jwaxKVbgGo
30/CYvE0L1QfyAicecLflkSZKfRCBae299KN6FgQj5CPoqxh/LxNuaBn+uY+OgKS
wOfrJBWALj9r5PSjo1uMbCLKI3pI6b8i+oVwsc0UOA69D3lzcfBxPL9BOapCd0h/
A+JTUuqAkqaqKLa6hgE3TRbl0XvUuVhd7jj/P/HXO7/1t2fu0GyGTk3hSf6xAsuV
VxZ4fdUcsWzjx7Ni7W6ne6OEvMZo82xNO3QReT5YQW6m3ZfMbCSVX59waiDJJeE7
fwxvxzySga+RpA2V7GgAY1idk9SL1xlwkzDKz7JBIFTiFBWr7vFXy6uvW3Uvx0zD
JrZMukI578EDH0MhxLyYOAyAQlj9TwxL3GOylOxK3jMLvjX7p5l4PcDFHikbFTKV
VFGmF/Z9glZya5n/M6dVcpOQ3NhLdLpNH15FscE+zZ7lXRvIA3rXHZpzb/S9arHK
r1SdjEu4IUrK+DAqybpEHExI2kbWh+rguUdbfyZsVatnnMsR6MrfGm3qy21v3WcR
0XOpUkgcncZOwFRVSGiUnuo1+Zz4VVaoW+p8+kfQJIjV6QkI+hEcjiBFo8WeOKXt
3iVx2FBCK+20OTlBPZ1zgR26NaSrab/r4XwyS9B7lyv/ZYz5VNWxuq7ONu2faG8+
bMt0uRUa3yxn2OqZSrdcaL3+JLU+1eQwN4dRF2aHo+ocFx7Rsu1oDXgqpKFFsCYp
S8thTgSeaJf6c1OelUv8+UqF6tbtf6V/rie8uGsYnWgAr5RSPTEqrV2tYDTwmkdG
xTnB4vDKjU317OETU7Ve0E/3w3QPBp5Btl1RNNJ/TLSQO3U4+XjJWOaTO9MNmz4Z
lZ4UfjM6Vl9p2MibGObQuzuwB6gqvfB4DIQ18gr/hog6RWAjyUnO+Jy+f+eqxaUt
wURWLD/HZZdzagxYkXhnNN5BXZHGAwJ00lttXqFD/S3k/p1rmB/1Rx/ZqXaLeLnc
cHK2z7jBY9HzcT5sr8my8ypbNmWn6qx28/2Z2f69Q5vahziDJQApXZtoGkK7/7XD
i0sViP6yivHT/eaTSOVR5IL/KL9BUPYQBmJh5jKfSV15URGWAfaZU6p2isEk7wSc
lO+iSB4aH6Qi4M5rJB2Q0QWTdfGk6DbN9Vvl4J5zOMoxLz5xLxUU9E1t793op9lk
IsqmUaRpyUN9txNGPHc0BFE2ozSAnMFOgpuzqKmSgjl/HegOrSyZ80xwz5BiY7XB
apkPLfKm1hXFm6CVNDHp0PdQHH6vGR9fSfWP7K1aYo7XJTyqeZr1mLrmwF6XMXZe
iK5kitD89MIbNz6uDhxHIlFznkrAVwkZF75C/GoUH/sUZl04NfUdk/yYLY+1R04c
4Pzb1+VEsdM9/57fq8mOiD3cWvHpta12O+ObgyOpg7yzrQH4By1EXyyLOW/4Niq/
LP8k8saoOCxWOxGVWkMHRRu0qZBDdi3zGthmjppigaKaKg8iJ9Nxs8dpAWTh81qL
fw35GLMl8kClizTREI6DUjHCa49PPES2C/4TI2LpD58LjhA6JE8POzedZhPZop/D
yxN6GVeDqMZBj6L/mIvo0JpDkwLWmT59OSkj2I4nxOvWTCB24hhvFP1mpv/Ir33p
9K+Y2JNPeLuNA2V6DHwgZJXRqzjAe7tGwiuJzvS6w/GtP66YDNvmLUWI7kl3ECEb
+YRCL8vdxgWh3pMAp6eIzP+vPp17+rKW4mSYRpCO11IdZXEs3Hn3K1pKdbc/qJj9
jABiwF3y0jROG9koOOP6ru/h+aR2kdj0JIymKMf9ph3gYpfqqW3SDS5qQy1OOw8k
35QIBiSb5toGTaM4M2FKYjwVoyKbt6VmfJubvV8MnDp0yyiQr32WBv3iHzsJEXmQ
76PfJuh9c3XK5oMUi2rQz8rS6fIKszUz7o83jPOdaQWznEOkU317YG+G8by+0xfk
S9KfHBkihYIygmsNM9p7ZU85BAkgU7jgIbMZ5Q3dOtTf87xfavqC1tbTZupiYPf1
VLN13vU8B3Ok9Qd6fTT5+uafuh6hdoorIoOy6fnO+B78v/wxmJadOBel70TJhRVP
dz/jrpK8MoFcIRBfyp2AsLrzKsrxTvWz5mpfQHsTU4hUtM1LgGtmkb8OdReywMjN
T+aSDOQskVU/beI3ShP9MleoTIUyo1r04YREtMfFipItWmkdTKqTmdK1HnGn18u8
QSoV5w7BhGUmMyAEDK958NXycxhSwlGLGQQ5uszPYK12PdtpERY4AcGg5MW4XVS6
RYD+D2wVv0R5+kkeOw/gO3xem2bXTos57EaCWo3OAJ7n/As7a9LXrJN0YL0BoJKT
Js3s8bzZ8Y4gHF3IlOQoB1fHmLSeWTswmz3hYh5ayBfGS3COtCnKir82+dcxhIo3
Ewv5TzkfOqlZbELFMdh45h7LxslaCs1gbDy/ddRqBhDGrm4JQ8lk0ZVaLK1b0wmr
N/CeuEL00l/gyTShpCjOWbrWu1X1ArtAWMzXSXv3LC/2aYUt5nU2o1UOa3r9R95U
OVBxWnFlJLFKc5qhIKGbORyuYxB4GGAblPazlMr4cvP0m7hqxIBzfC/4+tNIrJLm
lhlqOP0M4cTQb6qcYUr8/yHq/FGiT87g5qaRbAXGawsc48BQNBVJB99nhGOp/YIi
dlAG1pE2EX8A6UeXxiBiV6IXMK/f/7l/q1KHJusCvZ9+N4+GD2GezCM2E0mkaGw4
3MZb3xHEfkhZgJu/ZxG/V0ZaPmaeOJsh3jCqCqsU1FCDRPbJznn81luzeW8rBGHc
gLzm8wVyJ19hln9Yx5ZijNcXbvCk3jnVTT4Fjuf13yJgKRTV6uHwmducmz4kNCdY
nn4ZOKwRyd6Gd/XA7jistS5YQTm92IxwWrjeJXsnx1ss5C5lLQllbpu1Qfmr5s/r
pO0TDMnj7U3Q1sVgHiV3UIbCMowxs54KY0okkpmmwIMbzaVxD36wdRI+ipbMoFir
z4t+SISaZkR7yE2PFBUqCiggp1bBG3v8ke4om1HagHXKzqGFvP/qf9DjQ1GsWGEw
HcrzxcZS6MoFM2vG8ALv1THHTtLYXc7zaE3KKQfYlplN4Qval982t3Y0dIgjSKwu
9vZRR3bm1xhjQeLNib8GGxN52IxynNbfxvEEGSPfTjP4B0zuUK2dwbcKOg5taHVH
hjTBVBGP6fwHfhhMZcgm7FuzHE3a4uV5R8Ast3JN+E7aAItOX8oTF+zAJGoMhYnc
zxEdc8F4PxiRpkmJoqEcNjky2RTRw0HRqG59cdsSHeElcFGlaF2nUr6WeVq1Rp8Z
dAsE8p0QdszUoZOiguIIehd847LOKAVX0hI5ucvehwKpT1pWSo8/ca4JsCLjns2x
c61g9grfUxrDnasYYwYbM9ICuFvcC6irJwCgH3UxYCeW6z4QBCfwCF3RXHbAWUMm
RW5kEi18AVxx8Fc1L4kzHWncxo6I1rZCrh+ziAZX01AMagOZ6vTcdiFzwwC+tdfV
xlWh8feqxKxtfWsK+X0Cc/dL7l69tZPV25jstk1Jum+xjzKBYip3dDq+aza9Dond
UmYcAwRU0RHTmaTCZeXAXQdrh5OuWrDDx1YFuPIodgXFyNtvqMnR4rUs/iD+zaxe
AhJiV5rZAGHjlrmc3GKeJ9Q3hMk8Yc5sP33E0QsO6B4xH2Yx/MnKg+R7eUaNMBTk
AcgpKGje5b1kRE3UTSKj9puRhM47BDrojujekC8LhkKsMaV9k+rPod9PEw2IM41q
4mI+I1adqYv6MwhC0haCow23YAxCPKnmeQCig5T1mp24qfvfX3gggm0Gx7tEBGJd
X8d2XcPc7/xi1U3jpa3OZDDV8buefnr0eYhqGc4UxAzYvPSNE5WR3dV99zs87/0d
vp8l2nlp6jfNmpdNNWBhg0SfoPT/WxLSUw+4jJ3fg2qkaHJM7GojzHthU+Zj3aBS
RKjm2lmint3I6DXuHtlZ7MPqdS9nChj3PPrM1iKGxFOFviNAQxPVQOl/eB+rfFu6
Y8ScnTvGvvQEXU+VD8lvumWgYZ/TwtIoc91JCbuJV4NJggna9NmGB0pD3il75uGP
6kUq2QUCzk9wFDcosjzvLD1In5DWUOpZ9ZKuzOpCIJvHwL+Cm6GHGnHL1zBTJAKr
AdyPKMLXBAe4B0PvzQnu29ND6c92uDFyrqOj6gf2JSxQvJOReLomADtW1UydNZup
BQUZi1KY2KrcEN3xW1TzBVISlRcSwp3eaNjn3IkVFznC4hO3jUBuXS8tx5gRZQbD
DMtIfqaL4ZdcnSo6P1CD1rpm9DRjnPH9kt6SMCvgVu1z1VN5AobphfNxH8kfgH8h
IaT5w7hgy8uWSbMzQwy3Da1qNkTIYRBiPLI0JzXI+laU5kKukvo6rsFa9lsiBFRs
pKtlJiwnKSSUDEYfPaZx3UvCHy4xVSpeR7oAEAC9dTrORwJepTsdXYnT/CAhuozI
3U+YeuMXUqeiRG/Ii3o07XWSzAZYI5pn610ny1jNtLYBO9QeQb8rafrcTJ82WjFl
QR9t0ZEvbE3nUG6UtMfrtVYZPN/MgWYyGzopqzRQGhV91vyB51FX5nwVFFsxKgwZ
Q1bR3Tq9owBGKfWLvHRPehn7+Ini/E0540T5mkpodRL50Ew6wvneNthSYD2f2Hpy
eMpK5F3aS6/6e9gnOjP1WKDcNrTcFop2XOPocWjk9fZFuqsCbWdoFrxr8Jyls1gz
gQvQgFuvb6817NRME3CSZxidh5R7dVcrZK31VCYOyK+TXLwh1n+KiYJ4sd275kur
do4f5ev0hLshSUxJ23vXaCS14JtQELSGLsiJAwhLlvH7gCnn4ytSzX1QQF4CY/GO
7ndlXgPRemT019iULdZROwgIzEz7dY9cdnnGYJOlWkDKnmpZaKM7iX6hqt6M8vYG
yIISH8p6/N/GYoGP1yWn3k6mXmwz5MQE/iYeGJ9YlTNRytgrDF9mdSpyl6TADG3c
N65/aFwoY6qeDX0tWdP/EtfOkTaYjv5WSFD2o4wGwWkSKC2090l8sjXMD8Ufxvce
W4mTzf7yFXlEthXwDhXAew/3og8nuLqxLzNpSwj8qVBP5JwcNf4fYmE90YBXGb5N
+MyfXscJlTBZiWOS0XQoTRS0Y5cqWb94moW3ckhFRo9sHuSvClqPOIUlgF4HSI95
vCOfIlby2MrrCZBjtugOZ7sqsBsdvMuM4sgSK0KMn99+XT9gz63nrUZJvVg9QqYD
Smttfd/jN8o44nV+fKb7PYup+BwwAxlvw+IxCdzeAJJWKJK1N0azJ0bb09giBh8L
RooZsUNKVUYzmRxwSmOTLxbhWRof5IracTFjbkYX8w5Y2p+2lUQ/s9mYlEHWcvqy
tV8PxArvk0K0jHzChBQ25S8iypnvjBc9smwK4OLzgiIJPS9dTpZnGkKS6IuOJdWR
CFe2nmyjgy/+LZzUoCQs3weGQs3kBXWkHD78hPfTX0eDhJEZYReazsQU3TghIaE1
aY9JO+NoMtVivXMig2LeE62Uw1laPbihYSTNtIixCvzZCC1Qpzl8mUbAVf6PlIaF
cgj43tvQrpy1FYhu8TlAzspBFsQ7HxBP4TQ80SINT3Jh376z2+N/udZs5H1zq/z8
VT7GVkP02jFYucMPetueoYRl/+norfbMzO119p66i0otKZCHqdHU/nrAlsEW55jA
kgc/xMUa7/31SSLXnEXkOMNm9euKIT35w6NKBC4lXazecMSyoNtzjIOombn1aO0i
BfYFlsY3ds5F8oBAqukiuJn8bUr+Lzodfz69biqbFpOaueng93Pwc8a0VU9PD5rT
cDuZSmKaVhzZhSSArPSV0nA3ZHqUVoCuFHrLaR3itMHqMdegB2AqPK9xY1joxvsY
zqxb6XFKLmTZMblk0Sd7IOusPp691e5ek2ln0V6ZRRuoICKhL3cMZkFCXxrj5mP0
EYpTGL59y39fQhvqy8/rEA1kULAWtII5J0azcARWs4kQtgXrxRHcCJGO8P4HEje3
D6shVAvREh9x3p/cWUX+nOzyGtlCcJVq1qQD9nHWLNM23dMtsGTLBWY2k2av86CY
3MJtOKO6uXQlYtCVb2YGQszBjjCfcT7HTB77dsv0ZgNjFUHhGKZJ66NSXYJ2KUwE
4x8OgpBYUE3oEnEGkHPxkHJ2CncTjxDfUzUkvaGqI0yFbAnQNO42pSuUv+eVh9Hb
mU4VgpY0fsTXARuy+p3Oqqgx8mCBUTHC6snhgBiiYEHFLtIxBqAO22Fh/uiQkV2W
xyw2I3lvffeHjDVOXY2frsfXsufwi9l5qqRQda5ZvYyxZdD1kQcwstAWl/vXzgFd
xvF+YFWlOBHjZC+wljD4R12mCu4Y5+cWwIgj23qBVEkcL/yNPI8yjOjbrFPlgRpb
4z87fLtw+IYsv5U5ESDcQj07WVQ31Glte+/pfOnBBavDwBq57AEoJ6xows458bc9
7zXsT5XR9+nIz6BnZsqht6BBreFdZ58b4u6uP++HDxIpZDBDMPCkHwA8RwwAksRd
rXZCoVDUeBXicYNrRaCAxWVGicdVLH42gozudOf8Ixbjgh3aZhx7/kyvs/rHuzod
qnKhlOJltCy8QP9U1ApPSKopMJzAGQE2BhlKOEHeq78+iQs7kGRwVg8eAIUku9g8
SKFmpehsapmcBpX+ajDlEwDrBmsMClbGcK28ZUVLdWGAS/eQoDxhc8HWOKNmiRVE
9VbVLfn5NjRUw0jgVTMDm07ynLzR/Pf6ybOu6/SN20v3NRGKaneTR4JdyGMSQviW
J7dh8wNlpTJsJBPPgQPNkLTtnz9Mc+vMwRdUCdc43ynhH94sfytx4GrI6Eq4n3Zz
1UEPpADdMPPWlNmT57yJHjy8zqOz1ETAtw1EaHATKhC2JMDJ2aM1gWN5JrQG44Mo
QCgNhxYDsjiq0kt31dd/OHfbExBcmdjZrO8eEjDfdFdachdKgcdedwmCyUXZUu1A
WloSWN1+/GRl7X2OETIrlT7SAYZ84TTtzZAMFXiiuXQyZwNejV5aMMDDTInLm/dY
cRJc7OMl96owFfen/J7sQ45Jwsou2VcUyFa9WoQNcosO+g22BFdhSgSTx2dODLw0
G6N+1jheQWMk5pGBpve2YkdRWfV48l4nf5BV00RiV1ta3Qj2wYzXWaZ8q99JhwAf
N53bqdZghpjAm3AHX0fk9GHLahtYu2bVyufVu6rHdCHtI5kI7M8sPf7ir/yqx4Ju
08myfZYCxk+qEL4sH0BjwkoBe2QF5lNt7HUB2x/NwBPktlcVV6J7QlKMdvetPZD7
dNFXqPRZS4D34USySkqhjB2eFZwiu7URucTpVlxW3H/Vjj11MMaKraRJC3CX/XFy
3P8Zb+C/6PdXLVDC69OmDN8SaNUnid2MqAsON8iJzcaUGTFjROuJWZ41Cx+gTWOP
IoncoZn45QeOEOtxd0J+RNoxPmYDRAN9UjaHFA4wYLzyxTc/Iq3NEwzh+F5cazq6
OyVzumcPaQEM6oIAj/XuI9rmrSO90B3uZB+1rha0ZfUh48MyX9DmVXEQiBUjPy81
88SzOaNhgM0BNXX/UAfOOQe7zXx2rK32qtTyxQIhL8LdDMtVGjk8Rot6Yxu7c/rc
MzgLXGYS5rxPaBH+igJ7wS/ZisDv6qvIBgQtQJWNJqLP1ykjNgFfPZOm9DZw45L+
ek89LXDYezHDBtdmdikOVPCdsuZNDbbv/9QKyuu40kp31d+HputxkFbDW4pVyEaT
/b0UajG9KJa2ChB63K0sj9cIAFllqiez1OBs8qGzEtaV+MpuFrfm/8KYBqSgbwOy
XNmDEL5WKkxa3c8PdfKG5Wlur2LanubFLPpUEcN2XZF7q9/ZLj5kqiMDT7jEw4tL
Y+1vFjqFu7e8ciai1BUCii+XB1trLeVHqpvLu7oVDrHYNUI/inEOYTTQwJpCT7so
MlKkFMM/lx8T7Q9y6edZCzdhnmgb6EeP6HKNWHpAEWp+d/m2JHPCfS5MznGnYIJg
WYui5kuT5CSJywST37eUp+3PgJ++gOt4mqcvWRIPsS7hYiKrmfGL2IXuqZSuYlsr
Ae3c4hy9qhTcJI0aqBqdvQRcAKwvZsu0njQvPzHfajZQOY7geWQFM2R72249chFW
bDCWkTWIGjirbQcU7TgcEuL5ZrDvueCwFI65BksBj2jznI34j1Rsp5wBPpU6rtB4
bGrbrXccMKvR+BONmtQSccGPt+aNEVVdWAKFPVWszhRoKdEk6fb1mpcOlGipscVZ
RIEvaATo+QjN1l/1hqzxRhU5d89Zub6mo6CuwjJGWQ21uvRPYxzvosP85Chiyojd
3/5p2ymyyJMpSDBzJ0S2abtkv1JvlXLs15wjIDOCslX0bAsjfv96SjoN+Sex4HNb
2K+9gmrcscZvCGRZFrcdD3d/CvWYUErMoe4c7k07NS+j461KHvRREqs+d6xLHOYq
b2SKL7fDcRE0kCMCool/Im6DcgQAh4TVG+4+zynyxCepevvlJl3aY3/731E5NQpH
8uJzOZDldqQ4b0oEHNvN5BURA86grp29OhbUuOeE3GG0A1AwMK/loKE1sJMS/w8v
YgUOUByJFpS1hPfTzqxof44fm/1Ab6Q98GDvi/ZIuo7vXMK32xSmWFJAVwq3dfPR
ZKmyLaSc4A7zu7u5kMcLxliHwGh46fsR99/HC9EnqwgogOpPtiV7qjirdbGiMN5y
yH967NMZ3OmlYHE/41SNKu+AhIHyv7S+0FFRgzhTObBqiQvRqjIZBLf5rVSKxnCk
H5bwajN9DByk5opawdKYd9jWedBRXRza4FLsIBW8VsUPsxJ1HBQnoZKJF19OWd1D
JS1FaLQCeZ0BTfpXsNgl3lkfKZ5QInuJaYjUSJhboq2FFYDbUNEprWLysy2zjtYE
I95ZcjhDnAg/57lXd6eCWkBtG9fIhEIgnv02rIMvoCPkQWqwfJZ1AWKSN63A58V3
WsjtCTaExCy8hsoRzfOnj1O1EZw0D4TjpBA820mxbvpb7Ruwol1Ui+MusxZa6qe4
jA9noKR4Mujs8xUjmQKOEvV7hgtm/2Qm16a0DOjUeL//miwj63ZqeWvxnxcCS5l0
WIkweP0hpCekg8aSU7Pdl9VhqE0TFT8l4dcNgCaoEpl/R4jFyK1u1LLCuSXRG/de
4mhsFaRExx0HIeopYC6tbbGhxk0ZqQDiNKNVs2m7Gqaq9x/0Lq5dD7v2DrQj8GPn
nTFEVaijwie1YsiNLzafV8bx7Fb0mEP4MXGrUQferaq8QMdX8HiguIAkz4PUkPlu
+y+v7KBU4Nrg1PuvPXvpR7OpTdhUzX20FT5duMKwKItypwTnBZf15ISnnfy/zk3g
dMvm7iq/nMcHsFIzJkhuOD+XMylGj1sb2jfxdNhDgkc/9Ckyr1G976Ctmn3Er2Vv
i0DRp0Q3QokYclWQ/QLvESK9SgDLewIUmeyVw9d/MqkRWYtFBYYNef/dRyC+SYO/
346HC0Tk9hegbUccmjGA1kBM9QyKtbHavUJlDNfdDmcLAbfx4yKC/yOkQwETwJ+4
r1ubsDxqwh5MCh//Xi10R4SsQRHv14YcVjXIyOPDRy7Gx20sSdTK+0PNVamsDGeh
IZBDtqPSeDOnFUYXbRXL+q4OL+5mpLW+/hjM/TVqdUOKBHlXAKD70f3+wRzLmLMl
iyCfJUFlTNniH63xkeL7oXNXdaPiqpsDGFXkwH8Ht6aNUDCWlIWR3Yv/KsJqqWea
JmfrTTMKmobBphjNL5kz1rsBgKE4uPTisOcz0s/BazOaImRwrIaQg5lYiHPE7h6P
aLoknuPLCatnsnctH+XQ82BqlQWprCtV9iBkjcOi2MPgfKDTnee4k+OfncOtB9DE
lSCxL2kJmF0HJr57tjy8m8ZW2OzOEzVRcl+92PnRJ4zTgvaI4qJAnCefdzWRQBK+
prsowmGV4O0oyHACN3lRgL1MJNFtKeLkGz+grDJSIaeK82AC4P3l0WmCrIbLFafE
4Sv2JzQC6KuvvzdemclIWDKUeyCAoP8MdYqYPJdFdGa2fJO5xGpC1NG0Jzl0plIX
q7Ru+aIIhVWTGz23wir5e/j6AkyDiy2h8Zn/8+6TsHc4HUgZ2bbdiiiJ2DnPgZcT
37L0FCwZQHA1RgvjcnOmDmkxEXbjB8/GsVokmE8HIQDCKjepHInMqdmu3Fdq/bBJ
5S0LKdcuB8XTxW2eOd9duwlHgIQ7Ok2li9p/tjVX431rHGDA1XxYV/JtDkYvxskz
uc3miu1xLcPzMzg4302uDOHM5yjQjQcT7aLqtJi35GKYD9RvTCOCC7eSB81kL0lR
EpLj0OitkvP4E29SKBGUj8BMEfqwuY45ywK14eMNG9NGYSISupgYdlYzJSvpaau7
idve1APqpoz967MCEXmKNPgGaQxuOb5IVwIziwk/IOtqSWrCi7+B/gcKjXVocB84
L56KuQtcoJsdF5uSvhe/KI/wuhgyrnMoGdVON0oBgvfo3grrPottPiulQjmc4aQS
XVaTWUIY7c846OoN9+8RDZxO2+8rsujeGAFYU0USydzY7IEE8n1VVwhFbXVtjY4P
cfEJEWlOlutWzfmMkawUAicFr7qZSTVcaGF4qkneCcu41IO7RnhIWW/cTdleipsq
6ybXzFKvm+sS2lyYmcarogEM/LUd15iqThbGwysagiWhtuWrf9/hOK2xX1scOH7Z
WY5NRQUCocxY1uEDpgtb6iGCijxgR0No4R6wmRWPQCydcmpxWTZkUU50Af/zdY82
g40yLzIca7lwX7BS/yatu+XsY3trHzbSZ9mL6BvpUKyP1muoGnr1agG3Oqo2c0gE
S3z7hDuJe8bjhYH4rd9elI9q0bdtObw6IX+ATf/RCEZWDXTg44FnnyfRrU6w+ygZ
WT9pCMcw7L9lLU3X0Asjv1AjBtbjvtUD6TSK1GGF0ZEVcAJXCkBu7/Y5aTnFfDVp
BZmCQVde7hMypM0HYb4tkJeZc0WAKz4cmcmWO+Zw1/YOfbRKlN0wwbea4klJiTVR
C4/bmXvIQzPVld7dBo0VBfLAnsn9OuLS0thbv+nl5NFTbRnrLFFG5ySwhd1hn0FG
zpmsLXIryI4u0sazsc9nRYnRsoyaA2oWkKqUNPoVdm4Fxb7d4HG32Me/Ma3FM3yJ
g/CQt+thWMU+vMkxgsL4VVuY88ABrkmmmKWgxgYXbcn8IQA5DMmAWAax2mr+8Gs3
dB9jd3TwejXYDjsl7f1LcmDktzeL9K4VqhBYcMOLa3Jt4o4Pf4Zhp3qq7qEtL7OM
4k1zPDWxDBr0aUSTj0j1Jv+qLhoJVHGpuInt8KJFu5ov8n6STzcllCm89ZsOsKpM
7/WyO1FSavLD1N8Xd+eCwdyT7HqPvkiClh3Pd6GMhWqtxO+K9Z1UnAyMMG0R5+oo
atIpX2rCFBi6dIboNvScMvWHoYxQeyhbcGAtFJ0v0fnQ0K2uYr/OJuy6Qu682gxq
087ulyQ6QgoO3Y3uqWLZz8NuEgRPoy7iHcwhSzzykd7+C8PU2OS6mzQ+WTLP46B7
t2CsLMsYBJyU8HYshivU0bVSFCpr4VI2SKFIP9wTLVvYmmyETZw+1eScllEBW0+A
Rh4LvoJUxyCjOt1mEzw4zRIBAv/mtsZNA15BSpnaz+gbrAjqeeik+u0AVqvLbanR
hKT88RJa0s3Lg0GvwFRo629ZtRJBltuMy+cDHUwkVdmBEQQF22+f9ZGrJN2RlQJA
tr9fuQoVq7HNFfMFE0an89LTzGy6l3UvptFZwqxJcOj574jbB73PbhsC9OU4gzpm
70r1eo+hDCPHbGHuX07qVBtcc6n+MekNLyWw1BjNvyfsRVOigVoxS1ceYG38vJYL
kvdXmV5tuKc6J91la0e5MKb3HX4G97voVxCXzQtnEGgq/u/vtXeFsS7S7B0Pnush
vSP8RWlLijTXiJFZ5/m2uiiUMmJCJZgw0Cj11pVWCRNuVL8lAZRG87JMunUU/OG2
3pdVfAiEhXlTqZTg/fZ/oGnkM1lD5IUCNyZXHHN/Sjq0QuHsz1I3mKa0356RBHJT
jUJjdlstXFNpQkIEhD84HgWcq0c6+BzrlB25XZ+R9Mq0MJe+deGM0X7uxRFiBKMx
Vl1ft35vHtxOohYVpbRCBvVcNUrLbrA0cVwinLTCUoCA3eOMvTyPHn3v3NFGhL3p
LrmfsAsm09eniuP0asNhaA+qutrMu94KK08iwinsxFBy3TKXmElvVF0nO3O6KctS
7DSQrwleVRATrg11964bclgzjb8YgXhF0FQCXGKxsRy8hyteNvPRiPch9zXx1KLz
VIbURvuFYi+W6IDplAbmcV0RRkrt1bm7x5ZHJ63PJDAyCzYMQ7oG3gO6ERi0s3cE
/V6hRgZDQp9uGwRutSVlRXbJjY9ABNW+27ZukDIB3yUrwPlRTAXykbd708FX6s3y
Me+EDSmydb5KF59YqAz2kPI+wmc6tKQWuvERR6aJUMIhI9TtRPB9/0Uk+Om5PTMZ
TaD6zEXfTjJ24aiWZyWJALtW6PnLYg1jXkLaGCku/NCkUhjileJ6izCJDPrtYRZL
bAQhuNlj45Xans4hgYUOYbDCI8j3dI/4KfAIIhcK+49uMuPiFEg/kLAKKYz0yleD
vODc9cdd9gk7oQCnHMsAcyC2peqiZocPMul+nhAf6lVpMxyaO7x6lxMbT3U7VgfD
0U2ld8KrGJZE5+PNveuoi3LLljIYkll3mKp3lSM5+iq2xn2QGcWxYkFQRnzdddTp
aBPOzJMdRShXe9DuRhiM7Rn6d/n8TmY4mK63NgtEvLDsImEC7uu+cfk155sSbYIo
jR2wTqNRSNBAELEoGCwZskjh/2T/h/Xw/nyJImCUPlLtKBSpjg+IrpXDncW0PS8N
3URlvzYTw5KNH8Ln1bbREYTjX0sAeqzDBbSBlVqFFnTGYTxL06O8ditqbV6+mx1c
egII13pdjyRGekjVghpQJ072fFrhTx/A1+JmV3J+BKH7VNv2U715vWiXXO/XeR7u
06Crtw7UkScorViYYQ+on9jW4r+uK9xfuSMDz1FCccHaHMTFsZkz5gOly2kpgSFD
d1IZdXJpZ6zU1/ZNWnO9uF37ps3elxSTTC7ZOg4VeoYpnuyjKIVVQdMVRr1JCoYH
E39ovucIfrLb9Bv0zmCwSK8F5g9dr5PG+2Be/iN79/m7Xe9lny7Pc4F1+W8gW/g2
atKXlLqnq9JaPlRmTi7GehbNig28gojMs2WZt29b3+E7OdyrHj5OLO2mLZ9EXyxQ
KmhPw5IEEDpuZ001SzwmQFqSan0N1ALra5QpWh4s25na3sFH/u/n+AsXzgYPMRxi
UQN6uTW1YYTK4kSZho6BUpOgt75++15UGvEGpB7rvbswHGJKBhbkdwPRB174pFYS
tycu5Tr0G/ep2ve7D8SwWvU99hpTqXEq6HRM6saYNufLuHFHAj30w5ktmqXxfei7
uiIs/KcNvkPGHjyylXNmsyC+7u1yeYc4suTEVE4F2wHJ40M144QzsdDeNbqmoF9a
D+XV7Fkp6mOy6RQPP/9ZYcqLPqEyulCLdMiSmYI05x/XT55SjfsXBR1K2XAUIc0s
8P32+qHLtp9Bv+hqTL7AWEPtgexRgb/SG4d4rHF+xCwUuL1v17aFn3Zbu3GoEH5S
UihtNNmt2R/euGeSmLvA4HlKlPodtuAdCy5EjvFQ2aNm/uVMiSnn8FXenKtANTCl
Q3Mt5s0VXOYmhTGpuBCGhlX870cnSOYQzyqr06SBuqiWMFbZchfr4QC9kHrDCWJ1
C5DCpF24Q9VeAlZfYgTQceWtAIJWHl2m2FtjMRhA5rWbIdRHJhSLP/ef4cviOE3T
ZpW1jy0/QNfpWs/rCtpVDddE/Lh2JvVFBEzY76gDROSay5YnbcZEm5kCjPL3kY1L
s9TAdvdAOV91h1bKOzAwh/ukMxFezkpWSpmJ2/v/5CKW5b+gJtqii4s0xBmBMVno
MvDclZaWUOTAigwZA95aFNNy/c96TgaJqr0wcvakJ2y016SeuZvadr5sDj8oMwbG
Ifl+GLxUuFDDa6Pwsms7qZQ8+5fRmIjRnJ3IHgr30wDdw34jeUrW4GwFGPHatirx
P/idZwfMIV5pRmFP8fdi9YkhyZFkPF9jy8yd2liG3VAv/gXb6f8sUTDkN2hqzDPb
fcCqdgAGTAca3b3vPeB+KDbInQhz/ASt08meGGiP0ckqmdIArE7r99XKwkhxIJgJ
JVh74gyLvnwBfw/s4mffvl6m1DxfaFM8Nr/t2khTmTuGPMCq8RhVfD8/y/DJ/CBx
1MKcEQr40bwaaOc3DVuKJvtMUnPuNc9adIJZ+YVtDXrN3/dZKIRES83OF5uvQLgQ
PmZmcEoE1wiDhn1T7/APvS37AraI3cz1yQXjDQov8UcH6dbmnVorVK0dO3osMQle
jHcgkxkXiUo/WaXeoW6opAZ0rGlPK2gddR0mpCyyVGjwVpCxT1DIhyoQpfNGYxRM
dRN66oL4bHf3PJv5ljtqikQ1h6aeCxxlItjOsSJRHyTmaDAj2386ByFzH70w3e93
D5qfnBoP6CKyBFn00IfAR+CkuytU+TTF/NRF8WHMoV509ZojqDOGeV48UzOoh/PD
HkvO4b/zrqKTHxfzty4Zp/Wh+8DAUDI8SBpf1nygIHSt5fxOpYDoV+aweAOv4Y8q
asi98wCDHvsVT8j8ML8RpxrKdfBEux34ZmNcG7PwOyPVYlSQgYTEmc89g5ifwZzR
Rabz0PsdzHaW4KjxkAOhL15aPpOQAdsXNf2ZX22DU9Lec0aJ6dhTeq18A5Kewgr+
0W82tqRt80sj/heltpGYBQwGnfcWR22kG6mmn07wXtgyN59CRNc28P4ybMeX1Cd6
raAM4hB2+A0F5zE6qaIsJZiaynGoelXz53D4a50TreztUsp5hgNxU+4AR3W4bQ4c
kdB1Tx+obLO8Bs2vHPuDLaIeMNGrO4A4RF0AMOWFydRQjmj59BeITIm0EDTwm0fj
FzBn02wjfGEgrWNTDDSYLzvqBihhEA5x1NBmTukGEn2oDd6RFh7u8HRfnjDuwW/9
JGVfjxh+ga4sOu8SmlGQLL2gC0dH+sR8HCJcs8sxRFJ1fLDmHU1+pCLh2wr4O5eh
SecGQ0XiNiayGrRHo8Jw1TFj2NMZs8qNxEB7dOCTusonVFCI5pTUJPSWeC7Q7T8n
zZbRH6jBlddw0Ox40ZkQ/oKDGAVQwQuzB4tZpyJJxAFXXTzEI/moFH2SoKaBoZDs
hi4bGo5tgE7XuRND46AAj7370mbUS262AwrV7mIs2n3gDO4BhvSx/edYnOGwANco
q3GGBMkN2azWfaqta7VaabgjtnV83Z1FNR9vm9nwB1KeZV4bs0itqCIJIrRphdzu
02IGCwxaLydvJEaZUdTDUv5Kl2BavdxHHK2Piu2RGe+XGgmh+uJFwrvpsGmPkPE9
cU0v5Mo3/+Gn+OmQWybtRTIj2Jja/mdcka1U7isIpNHy9Aut4OBprbXNHUbB9w1w
xT9zJkX5D2ndGB9IL5H+v0QFL7gXOUFcrads+0ulEVc/d98r8gAEVHtDPiSMqEa9
y+ea+SpWmphjQeYENnR2CaVoDfIHjwSEwSccqWRHy+2esc2QR/Gxafpv6em5m90X
5Sxskp8mbiX+vMoMyQncBl4GYbWlXXmNBw6nAS3tVvAnPo/iZpECmeL99uL2K5vw
ZeiY2agzj+oODt4KPcB3hlr3wU+2RUNw0MCXbj/wwKtgCW0hrRGcph9Gcz2GJRTJ
3CWLhe9lmYbFMBXJfqWNfiv0388tIxT5cEbn3Q/QvahnqP1FgwKsrf9NbVQ+B6DI
zMYay+nCJgFLBztYQNWI7nZKpQJi1ikdmK88EnsXrfIrKP4VAYz5ejroDR7kMtAP
/GMzAwy48Fcnn4pRjYcLW1epi9FrboJzAJw/mjV+Ws2pyOJLVjaSAUVIoNV0/6zZ
o3u9Y9D9LufojSlrcNXReuiF3GvO1+HW3MqZZy8scjHnUyCeM4gv2k8CrZ+xamNe
xksGN1Q11jM4FYfbWac/kxFeJCnPoaILrdP7J71btPsGOB/nIwK5AAsJzhU2iWFc
J1ymyVVmwctXg1YGmX7DTOpoe4S4Env0CIJJ5o5svA7fOpNjBjTqTv/6T7SkpqHB
LJJ5UwyQqWJQ1h4YlUJchx/v4wXamwLb7Cmk3jqjwC2QWixgM/UmD5syOnTMNHqs
BAh6B1/sxJQwyv0y6oJh1ICgpHY0waZkoaKbe1VhFga39IUXzRF/+2vLKKO13av/
anDA/Xc51vWydAkYzdY0k34/AZpfmApcLxlMFewlUnA1eb6wCn1NqxcrKE6s/zZe
3HSgGxYVS2MoVc9VDn8c0xZ9dtIt+dbI/p4Dx+WbosdsGlHOf3mGR9ihOYwUHMiz
pbH3nVFoe1Q9x0Ubx8kNnLQ/PSN9ym9d35Eh9tVvjgoyqTSK6CPwTuRsuieaBmJw
Pi3I7EZDwmzmxRWc3aWKLEX8HdjKTne5P3xPCJlT73bzRT0qu5CV3FfBSPXXwgYS
GXNC6Kg5xomuuRsS7zHJz2MPVrv1tKeKbSwGtijsErE+SqyY1cr99Wnxz0dygHx0
/4U4X3Q7m3zom5na1AWTgx2+1a3gXd0lMx0gPCkqQ1l+eRJrQ2nHyQpFMpAc29PJ
wDjNz/2QUmp853bpLrhXDFWH9Rwd2sfjOcLIbHsk6gv3KsxWzhUzmatjlI0Nox1k
uTqx+6g3Pu3FEYfpiIWGCKaLCpgza5hjdokr4IDcEmo2s+BuEJLn9xzjbBh1mmLl
ptpB5spiRHxqqEchQlL8C73MUrJ4xr9Vg3TuNyf1t2LP0xQIB+UzLQeIBDruaViq
HPVHTI6k3jq5+dpPwbpKHQr+Jf9eWLEgZDyMPI/ct/xbEF2Q+HpNtMb3UoIlgBoE
fUvB6DjTGdAnIpug8KId9p3iohq/wc2O4JMsz9SZNDSo/6eyMGjj9tMtlFXLpX5d
mEWnEMiJeItajBLp/XyoHQv0KvUSyTk8cyBaH1M6ThQ7BP7Ih3izc0/eSS1AYHl9
2DRusbkE89MRDoLlZ1UXU9dhzG3G1sQ0LN0b5WG6IdgnrZGaHUtRovvAoI3l7ypY
FOUwV86dG7uB9tB2rEZw1G558FGy4dwZrlNumfJaby6G56BfOrfHCNLZ3nz2ov2+
/A/v2KoANm0Ae4klOAV0P46C41WxtELXT8dCx+qRLiomZ2QR7xIoKiR6ze9tne/v
eHL7V4m2+2I7DNari2T8cyTbe/R4SXGtvw7WLs6Pg7EkZ7TV3H/LGlt37yiTGw4H
Z3XUjekUEkepkCr7K5qc8JTJ73K58J5q/qd59AwgPIlL21gbcMxF0LW/kiZI34eL
QVMUs1aHwFQtq7yR1WhtpOmWEs8mxG4gQDYpzCSxya7VhgsTycwOr8MpixNZYuI9
p/VLKLJ78tvvARYspU1btHb21CXizTUOu4lExxtxlvdwrLDUex9hOGROLboAaSve
Cj1glGPrrTydEqYxj89vkBSv6d2MSJ4OhpEwKubX1KOlLEH3PKfqdT+UGrViAJQA
IQbkmK5mb/ydKzVt74rvTIgZzpjBHAROkvR+7FMGajfs9dLk/zBEuQVWhATqKek0
GIe9iNXqZzfeb14y8YRrx5C/QML7DqoPQB4Q1YE9VTwWTNrEM9+QrTidd+3XlCyQ
NlLcb6LBHFxrsPV8zSHsvXZT02ObbWDYMZhLQL1O3hDUF5wW8TnH3SQGoI0QmnzZ
faNOz8C1HSmDuPdnSk+6k8xw7JohVdQtcYF3n6/elo4rntDKY+WqIWIKVlaYIaNb
P5hjiraeIMg8ltYDE+gYKmqcSgpXfRjNDbFfmV8hSIqXfMIDT75jDjjBoAS152z5
+RmrgZUpiKHgVGTIvTbsQCXhurcNAddUP5ucQbLG5HDFWgNQHCAaNEXJKg78mY4N
/nB8ENuNqJCXp+mjnieH1Impa5foVKxrTTCKYZHlpZd0sY8e76dBSTnE8fvgNgLs
8bsiOdNZ1vDkDE34S+ISEcu0/EOvtooZcH0ChpfsBKBsFRBvnvPML2WcNXiUGQa7
vwlLv48IszSMgTtZZnfah9dXp+HxBbOOesrh4GuH6ET2X8ci5+6RNN5IlIKqC5h6
OaBxe4ZekE3wL0hPxBbKHbX3pe6dzEgHTxz8PEHzmk2i/Xcn0t8HnG7Ky+0wE8cY
LPCPhzqi5u8eSUJ0l/OFSl6YNYUy/gBqB8cb7ygKp8Rvybe4pATIeWzIwqcIW5pN
KipOfhqED70DjcWL6Lv3YaJVi5hcwLcgyCesfmS+XQ6uWAJAqujENaROZSZOmXRO
h3ssgehts7J+tk1ca2yGS/EZia6gnuJsAD6gQp4kXwi9BFBv5AwoiggXj/pOnsWn
01zSeh0AaAvWcZa4CotZogBcCtc5PzAwrXvD1U1gRvJprIdX7aFDo+JXffgG4NY2
ndJ5rFrfQ/ZwVH4kMsdSUQqB8tV2GRa1aj4qrjwKa7Qr42CbJFMM0nWAw3JP/MhV
HEkRmAFifm1CsoYtCIcIkLI2rnGXyNim6zmic0xK7xvyYonwxE6JMSvHBUJHvMdM
8fqLMVEQVWLWh32o5FwU5h8M85LeK3lc+E8Wuz9msG+WJ646NYeFmxeWC525MJb3
OUihEViiiD2dTV8vzA2SNMIB1FO6R2e5qkA8NCKyn/EPTcVTFxaCL3CbBjfqi/C0
bxsbi/DzZGg1bB99oip+nojgf6/1OpLC70MWSDXHeppoijwQy9KQ1wU+TFl8d46t
+0KY+MPb69LJQ23AU3zGrA7+wGfLfURLtyO5Uvo9u6lI3SNHRR/Ss3utIAiFhgKk
5muXgB8za4JfEAXms5SLPW3TJMSIb5V/QLMoN2gMfoscw9QGafKosi8vDRAgrHGr
WAu2rbZtQl42xvVp5VpMTJof0Zy8Xt+HTDig0EkjcjrRiAq+yZaiEo8b3EO7vESI
qJ8CnDmcYhbV3xl4uhWhbu5DUzHBS9iVPzQJ4SH/5kihdv5q+iPMLNU0ollyhUFz
7/wGL9MWPSpX3oRhIV5bg07XdSmOey98zYYIn6Tff85yprz3NPK5EMpG/YhsQ/h8
o28TC9IIL3Uk7qxKiaZbSvSoKz1U0DGPCrW/Y0i3v+lomwz5CQ/6b/C53ff4RmAy
aZfxKEYKSaveLT5ZB7mVPyaGkYqoW0oNB0H7MRvuSpRsEsQrOVOdACnxbmx2cW9x
MWCsu/Zgqh/pcBeMGgptETtwt1toP5D3A6ya6v6RGgJhuBP3pCHzSFkrkF58y3rn
fsDhNSWsAdlN9hhchDiQnUEmixuivbIQaiBaWMC8pFowO/C+eVNFNnv6iteSbZ3M
gGJC8StTwd7WX6OXnpy7EzfMoTa/9EeaVlhZdP4+sq8FSFxdXXTgyKDiTC/DfyQz
OYDfXzyhinwCN14RLRzBxe5UCA2+Fx8A4MssechBwY3GdkEi+uIm2CiJGIuHs298
uzxlqOJ5FC5lmWhPICXgEYv/LYHDDEl8q0tBOd4DtjCy3AY/buxdjHX+AaQ+bodd
cYd3ZBKDgfbAAeTB7ovvG0aGrys+gNLtgapB/614ucrQLYanMrMurZGLjX0pqhOV
u8CvdOp34gCfRIZpFi3RiRIMvH30nul1ayLghe6iWteuqgAkWAmkuWTw22X1L98S
5djNSSlFcHMFKX97IfqGDN3O5ieVtx/YK2wKl6H8gw8lspgQ9xrJcOfu/Cu9oara
saGd0VFa2wf+AcHh7PZ9HziVTWUwq6MspbDFOCMGjCQRc93sUzymrJf0o++GPg6U
KKZBsrgMkgzOM0Y1tTO181Ws65Y7XM/Iyqinm+zabfeNilmF6XVHXaxdBlg1H076
UsGnc0y0tyg4Gf2etL45whaVwCbE/+P2si1Mi856SdIN1iNesvd1kuuIWuxzGYFC
H0XI0dZKzWituAYJ24OmQ5MBU2xajcwEYFqSNkRrYH3+z7PM8vaYqM5ZMQB62LX1
WMB4qxRNAt8RMajTfZAYUoZD8nAAqemZI3uQ8zMIFgs2AV48Ge1ukcz9I4TIM/95
aQA6gJb1Sgem3Hck7feLdB+fNREMpLBqTrq1HNikg5eyj2VhoAyRZ1prBOERHA1U
/T4mrZWRFLRCOgChfO4JZGw0hlII1AfdZVvc7L1NXx4TBTrZT5KB5Vhk0UUs7re2
Rta4j3kWUWHJ1FD1uEVjAFYV0FPZmu8qZ12zmWnhgJtL3uWFd22pVLnicsPs5m3f
EwUZHQdyuQpxpN4tz72BfPpf/MXcwuTxyRiRluyDCAd/xN1sOxcR7Mjr0/djnXqO
tUGB4XXpSc49BDKrOj4t0/17uOe9BsCJMmo5g08RN5TLRzMpHln0U+3PcbN7SdaN
aXZBgsBprz1zp7PjfHYo170d9rwbFVaAt0eVxPW303wWx6783U2JPpLiASGYWq6R
RiXwbH/57aa6QDV3aT0wpr+l0JFAVCOu/jed+S+I7spZG4DePf6rs2/hLhNOaaT9
mJzwfhtLxERACgSLvN7PAuxkv5IasFwmOjTpymWqZJkSqlToKiQpqwH2akNXrVEk
KcCDHt+FGjxwMOqrkHuERWY4Iolbr+EckYrpwAaTwLnnq10VHao+OBoqWqpD4FKk
jlpZddgBHsQfYK6WHrF6gTYwCbflaQGlMzw6Ip8P78WMMC33+E37WT8og4OFqdcJ
XlDx6KIY9lUpk5lc97qDClDsjhjE8lXd2Dk17OMbttT2E0HmjnJx4GsNwC1waY7H
pmbvZ0MLcaZzzOgCRoqLpPH+Tq5+BWZY7UQhfHL89L2a/W7ml991dpAw8ZDm1gBU
0VPwY6Jar3kW87HtBt/KIknmqh7/Gi6qzdKovLsDobOst5JcItScJJh6IRbHCvV7
EPw3GMcSTfda6l572sY07thCtWQ84Skh4fBovyLocQ0Q4N3zz0j41QYPW5iA/bcU
L/UugOlcAUrb2GFng/JWggdcNKEDYm+DKb6OcikbfrdRjdQ/g5ZH9+T1KzTobHyh
yKKBnhdFv3hBHO3S7Ceww0tnLPJKgmu/PEc6RH+GRMjlOf6iRyVQroNCRzllfvuu
`pragma protect end_protected
