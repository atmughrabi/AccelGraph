module cu_vertex_control (
	input logic clock,    // Clock
	input logic rstn,
	input logic enabled
	
);

endmodule