��/  ��9&\��6�4�[�����<��=~6��/,��>�tSiːn��UXlHq��,_�����f�����!�\�.R!�9��x޸&nTi��jIIw�$#� b���p�(�6/ۖ�2�3�Z���H���t<����b>kY�ȼW�h��\t�����Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9����A�\Z�� ����J�(�_%��7������CA�O6v�A��
Dw��W�,����*��:��.@��Z6:��8�����@=Pq�R���Rxp$�ːi�#�S�&��vS��4j���>͈�7v��8�P4��������^�:m :��7^T$X׍4 "TJ����.ͼ�l}�� ���<{?X>Ks'Ao�����G��É,�>,���y,�v���Mznb3�之�9���&�<�k���k����%sۍ�T�D4,n+�;�����	\�//�m�a�Z?�wq�j�Ogx	z���L�S��OK\���s�i�Bc��L֥��G��6�\�{ت�� ���h��A �O��9�W���/�2�R�k����q�!Z-��_�P �<���Q�q͘��-6��*_CyI�Q^21������d.����kLS�E�BQZ;iI�mc�ow�|�/������Te@���y�BpqU(�����b�p�"Ұ�M2�"�5{�"�+>[�:%���c�s��9&N`�S�g���O�q�Q�T���|5����m�A�/\VB����]�Ɓ�k5��6��u�`�2�[����&s�-��gc9��b{�� o��̰�S �=�V��5���i���$⍳����:v��x�����y�E����Ș6����!�D|\E��`c���o)����y���)ϮY9�(����/~V�C�Pt�U��F�\y�od�� 6�Cc���#2Z@�!$w9�޺�v�!�!�Ʉ�-�}�ESzGR[<��(OsC��p�>��7�<�x	���#N&�*/���<T�������7�O�s��{�l���ȁ+@f��Y�e#��V��t�������G;�����y���w�g�/�v//�\?/6�M���*�/D��K��Κ���C�����m�ln��Ef�vt-�gf!,U��@S8"���|+�����_>aXU^�8�Uz �[*a���]%.Ǒ���`x����n ��c�Lv�����O]�̬H�?����?����ƺ�UT�Od�X[W�
���R�G�n�)4�k�����b���RoP�c��>�֗"�Ȃ�Uj/'i@��D�"�lY����>�w6�uX�ί�=3�A렛_�r�|��SIr-��GH��0]�)[ͽ3�kX7�`�H�QNkj�����s�ϼ#�-�8�tHʜ6�7���7N*����.̽��lE����4��4ԋ��b��Z�a ���a�C��o��528��� ���?f��CA�T�<HY�N���u����}\�`]�/�J� �\׹�����LL���)W��o ̡�Q�Q=(d�A��I��y�z<���8�6�t�(|�������Vb��FYe�'��f��.N�n���H$|/�^�T�(_������Z���VN�I8"�����9X5��-f�uJ�8>{����ԭp�z�����q�~�`tch}���+�+�?Dn��� ��c���6��Zv	m��ۨ�����Ȋ$��ER΢�N��:2��L�ɑ~�뮕�