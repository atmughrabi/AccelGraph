��/  1Qy���D\c���
��k�;�]l>4���e��4C$( �t��e���Q�.��sҥ؍���4/����k�����Z@�9�v%/�ס^L�Tx��T)��m���y�t�)ܺ������=<�E%ȯ)�(D�}g�����8 ������bW ����Ǽ�+���Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9��6k��`[�D��%>ˏ��֯�zuu�;�Cvs��Ӥac��0��^}�v-����Ta1#2>�{|`��|M�����}'�������,9���[^P��y5�Kd��|��L��eP�k��Y�oΗUW��D==����	�޻_u���Ǌo6`���J��=ʪԩ��䬋��N�V����J]�#�{�P؏	�-�~���n���0'#�lO�L��T�/�*�B���@�<�����u�>֝v�b��in�?V�Lfϒ�݅Q����X�b8��3X��/D7($�C��& VP\���\W�zNY`����rmRPl�4�����v+��(�*f*�}�(�,Mc��3ո�1;���W�ݔ��&���*���YXJ���Ǿ�*�9��yǿ�@%�w%�?�v'�H㱇�`��Fc. B�i�-g���SEkR_�X�ω�0��azjNQ|��]�wB�$�t6C=d�������5��o��h`4��铒x��������n�߿a)i�P�s��%���ꖸ�uM{ڛ �4�P$���V���M��sY���V�v���^�ii�+T#��M��������7�ݐ�H{��z֡��)�t"��@�+;��_�>�fQβ�S���O5���� o�E�F+c�3���I�*���R�~;P���� ᢀ\#�(�j9H�"�1"m�߇�xZ�gdr�