// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JQSm0fzUu8AcgY/8hjQwxBg28SCjZ6poAMtigmeLSikXMK1pOrweJMiUAovXRyVm
mAOxhfWeddieN6s15PpIIf3pr0xJT9mn4YMAhKGx8ssQoFbtd/8ekRnfx9M92kNe
D39bORXozbb91Nhj48qa/pYra3VeDA+NDC3l/TV9GyA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2992)
/yEPe8byIbHLi6wKpW5abHhPcynUsmfdiYkjGDNiQJQhUx89lq7xOhOmY3g7lL+g
IP2vqMuE0b1Mi65dOFhgT/4kv7q4GFQErR4FvEo7Bp4WJrJT5njRXCJ8gAPvdZYJ
wLPHntCONUVEYp20JtNUEVkVwhD68wdp2tv7qFszEkrBvQbF1XH/liI5Pq3fnZBu
oQ8SEquhCobdOmcjX9e58QMFgLf0Unb+ByL/gtFKmS7gPxCYyWkcQ/Hy3B8jnEuu
cx758LRy5ToYI2vlI8mvlhGTs0iCsBWP2Wb/HUqXXQQZ379EcIsBDkto7qHk5IVk
mTm1L9YALWZeg9eM2QhLxJatYed9N8S8lyduo75MDPkSqyXjsGz9ZyMXAcvoTfD+
in3yXG6qnSRxycIuCKPwL6ePx+GiPlCXfPemFENljSDl92Q8w7LG/22GRd9n/l2y
vs/UXOU3cENRp3fCcf8PTSe3Ud65YqIfmyban0b9IvauriwRlXlYFSHjpLF2ZjQh
wl6qzjbPHgQhACtbmnos+KF/1iBg5S3uWBRcLXlIxjQMmflvEgtRuRVTfxOzSi6Y
e9JvYRzkH/q4vBSqt6hDVkpwm0JWtyhUnojOSkJUIiKomZ8beLhlPu9UrEU8rmNn
HWkHI8XRPvV7ikm35KWl8+9n7GoNgLESpK/DyROjjDC7SAzPAhbwgCyx3V0hC8g8
fO0gchOqTjKJxARZvD35ufuZ1kmr3SuRUlHf+Rry3vUUwoB5+Laf0qFJSZQYoeUk
ZqlLsmGf2TlvGPMBuweldfmHsRQZ/EnlkjqRNAS16riWCod9FICSQMzc+o2aaTAA
uY2OgF1b8LeFdzQEz7bPg1OVILla0zWNuRuzKU5EQ3V8neKRNChEpc+91RoQ6Uzz
trCh0qex70e8Lj6SLXeZ7gyj2I3wbUjnQMxGX6a8e3T/6RcFvggSq0U2+fpGSPMK
Kmn92Zj/Ut+a4cfogqMYa9nsRD37cgxA9+7A1ivFOVcIhIZzoEl0cEw3bMi+8HXs
nzwI12B3Jtga5JmXcvBOJuTq3zNCp9FROo3HF+33w2bjxxolm3zCAkd0HAWGpQOR
56yaan3zZtZPqCnWNOEjYg/w0IxBN2OKI7QUPYuzQrtg2/Ede/daJ6jzUOVfnU+2
EePy45AhtD0tFiTvIyyUWc7IKVORdq01HjfYek4K8MJdkpql3vIltZrSep3HKrwF
n/bLymZZNguLiWycpAHETbe3OGD+S2YiXNet3UqM0EHikmiG1MPBJgX8x7OxY+fz
16VU/D3Gi+DtIDPKglV5hCe7UwIqPG1or7qbi62srtToSBwKfjaRm2dI+AIqk8YJ
xMK+RrQVVHidtm5bCvaxULhF3EqNdGkHY1cfm1JH2tX/QsCLat3FEoqNx7uU6jyU
Mjsuf/vDwnJAa/PReoJtPNspGnO/LLnnK9fM9brhQN5EkHEK6+PZlaPPkVKUAPHV
RUeWbpT78aWRKatiN0LjMD0uyFXKU5xj8P6wyoEcETztq/unGmN+AcDBhisjXwfC
+rDHp2xyBzEqdHiiDSLnomgkbbI2z96gQ6KKRBV7e9gE1r6NAuf1+0qK2GrXmSFP
X3094BOrIF1GTuN+JF8Uo1NfwqOaH7hgBlyq3uyB2Xy3AjorhTKSmy69ti56pWBu
RE1ugpi03ZK29gu+DHFkAWcN6nElIU8Dz3TKLdofPehKBDiMyhf4YSi1NMgS6DPA
O4gMEWHyaKT5xbaNX4PG29K1Nr2VKtCwbUjaN2ocHN/DTXKN/yUi0Q43UJdKhZc2
2yk3A5Z6hI28ES/l7YmgjGQjmRa1DIwI6aItyM9RLxZ6Swh6PrzsHXoH5AkwEnIe
UUbToudKVrf0ml8JgL+iESaV5b4g6212dxEGU22mkkf/KQRcaRrLBmPidiUtMye6
XZ7NmAjJAPs2kzZoxi+or3ehFMOvnl8AEO4xC585lRjyK2WFqho+57jVrIlqti1b
TzYQISNfsn68w0fV2q2YfOokbjUn6f8edY9xLJDBF/JZ9A7hW4xJE9h/Q//1/Mtw
P+Xr/vDQUQwTiBRFa2sJ/K+mRZEO3o3NfNReejjNbtc1IT3n8FOoVn5MT0lOqSAz
0LCnFtHstavP359qHefA+IPWb64pb9reynGF+w3nhkBylGqaNNEUNQdTXO2xoyov
qO+0htDuR4NihUvVUsEzMP5TNYIXVsudMYgPdgauuRIia/xdxPKO6Iguhcyp4fIm
SBVKctWm5Mn5BUFchF0kKtKS8JYqV/+cn62lGQaj8rSFF4j89i9gyaeUY8i36yb8
Mybp9jl2J7W2lnrT8/2LDxJlm+YFUTZbtruf92dm4ls3t6tnxr09noftLcuN3U0W
0TpFjYJr1GFWPWgISR4zErwPqiXvAPj+uJyHPR07Z9Wbipk5chvOEhPNZ9Q9t7iK
PfjRf5T/M/MtdfjuEWiA5Y13LVXxUuUc9UM1PB01YSiweye/hphAdY83LtZDUoex
MZXjUU3oeEK5cHnbl/ei8mbGOmzXUqBYIygtGUE0zFNYKPPEtGtwm6XLSR4qMuQ5
yvQZ06OyiQz1fWxoMd4bjQhuZZsKuawg1QVAUAYepk8mrkPqGRcHZ24u0O34e4kl
wWWGfOX5tDa0F87vH4G7mApiTZBdTguJ5FqUDZXQ1u1FjV2Dp7eW1KxgG4BCp7WE
YzrgpLhgyMvWa3CgmK/lrhAXGSHvjzfGe3fiRniggGEkcnvIQ9GqlavSuYgANqt5
7U2ubUizTHyKIauAlC5hcLHksx5sqJXJQuDogX3LhXxlZT2UUS1AUYSXBxKvmkfP
hSyepdalAymJtqVVzAOtGRLHuKeSPQANytiJrOkP/SKwfI6lOLtB5gcFTb5hwhXr
k7v5OHf52knhHWbXiTMRsNw0B9BKD4UH05u5k/GwSuZbIFwU3NsHEnOfdM0qfqvq
gXxUoN+/AzzFItQM+rcTx9zvQvzmvR7nO3iE6ODdvuBWxLXHVnE5/qnsqo8YKHJ3
EmV5REo6xAQ960nelthIi2YTHqX6W9WfCQagaDj8wMsO0UGatdzAuoXy07SbSixh
Cvc40xoum43C35hi0Uy08nHFSR3bwWWnwF0YSkx8O/sU/8wO0Dhh44K83QeIRVXD
BMByJ/cCE69UTfRulCY1CBQXKy4CiKSMSRJLLXBhqIxmUfSIfY82dYOkzAlkZJ1o
rn6pjZEfpe+zZw/WiTaloicPSylWDhrBGgwsz1EgU9DaP2WwceBKa+a4CKyx5U8g
t0r+TpgU3D4KoyaGqp87acb+kBjTJn/PnljQ61BM6lBZOA+3yA4o/u4Mlm64OGTP
F9QXxqVvdEFVfe8iXiBwvwtYMEhq+xw0x8vG6Ja92qRE6lqZqMsiKeeWZ4Ye7oQc
ffqc9Rbr8dKpiZpjnRnx0RY0u6FTRQIndt7n+5Ti/vMIm1kf/jnttwUNa6Eq7FI/
ZqD2xidL39/hVQr40ZXsK+rWuT8dICTUqsB0sjr4aAv9W+L2mIeDQnbf3bFHz55R
18s9mtNvC3dTWUExLEBNtsAmHXb40aIFCxCNobJEnFUsc7rowWWQFZEJrbda2NHh
J2duv2zcVUAkpGms89YCrgqxwhnfm/kFddxy/U9NTQSCU7o01Dlnd+NNnE3rL/En
kwZ+Lx0FmVyMU7rsc7TIbZe9K8g8FjA+D5UgDKP1hwDWme0wEMaJEPcBdzSPNbvW
wHbaJc6SBYNsShacS69fh3fl3MoFGvz8opYHr0Kf8HzLd+rVSKodoeSOgqFKg2Y+
ZKJITsFzrEoKXxBbCPDrQJrTa6P/iOC2604ERLeN70xBLBOnSd96+jWfmb8nhOIx
lxC1LTNw1IArskSKW1GKhc4EGgO6ZhPIE+vuR4gPCBI+jFGgzbEBF5IFfV/rQW+j
f4OwaZbUGj0ZkVgIOJYHOcagO3r62+Qv+K4nkW4Hmju7YT5vCcTui0wzRyp4VtoR
V5Juwvxkad3z2SlU23NV6g==
`pragma protect end_protected
