// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
flxO6Gpnj4L7SYlDmqDChn4WDlA52cR/zUGrisTZZH8g3CFlz+cGCuLPv9tyyVmz
evvkI58uB2Rcdcpx626YiOPJnX09+pVy1Zb3aGcO0FEX/fw2t9+0jjvNid+Vsh9u
12XAcRlO3QMuMuwJJhASqUvNvN34MLuLW1kk3XQl3Ow=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12080)
PyDgUWEG3wNrLcIpec+GoSAQV19izCThX3EA5lNxiPGS7wdwVA7VrTFvnkB+P5z5
bVPnSiTsIAN1bM2VV3kvwzWlOpw5i8SuGAmZg9LgbgoUa2tAtSt/SqF1MJPqWc40
ST97Cfd6aM1hT+57ip77PvteOK9q1/XJHSRU8I5UL4PvV/5Zs1C+HsSeU2ulo1Fu
TdC6Hb5XemR0RqCZeBAP2+aoqWAPS5Wa6lo2sueaDTDFXqPcCifEAxGffGtL8st3
tB6yhVMP6fw4sIzkbR19yO1yKIF3gJVw0yCcYilG+FEZ33g5enniV5mVxsmHHECQ
/TYvzvNT17mKhKC6TlN8+Ja/g+jz4RLNPDQAMQEdHnGc+sehr7vd59uuTQYdQc3I
TrHwCuDKOx6XVSxJta8GLTEUslHhFX1cFrJWcB7jy4dq+6t9XDFvuwrmLMEJXQ58
se1GlHuSYBkIIrz1jkyz1NbaanKZZNvL1e0+vTEpCaDnD5IlQUykkjjMBgnDwDbS
A1lhxIQCr0eC4U9VR1BY+QC34xG5vrOdj9w4xD0ZssFNbkX+9NllZR+3vUWSCIou
7K9GKSgI/P65mGxsnQ4wYZR9VAQjUGrH+tsdIqASoJqk2UQfDU5A7NNa5j7zaDql
0oXON/uvqFTWdmSxVSYlLpPg9NYEjfLNJkBCsfeSoq6SCEIs8/hQxvukxDVGgLgd
VW0+QXZwOqLUf8o9i2UK5kcU+m+4T+vu6RdnOS+Gb8H0NgDQPPeO3BkQD+kuc9+s
EvouyPqgn/JpqTzqLosynm5UtdPYczeluHNL/pDgyYWXVTIymanK4asWhNTcZcAQ
IFsH8tP/nqBZr6thYd2ZMecoEIJ1VE1OBZpPQvDY8bWPPYeClPewz1OIhKA8W63C
Pwty0bnHOh3Ev4OvOpWN9MdMXFKhQF1gE39e0vwRW5qzYo7UBc4WJ9bAlFVHuJKm
IBsz8PNBsTTgAvcKDy9f+1RzgCOl3Uyj5ZuOklhOLkjbzXa3cD4jE9Wlz79Gw/os
16AOlnXStozbchCsjyg97Ps5q6+6EfKWsN3dRY3T3A6+F123p+o7CLUklsjKXfAh
YnNFpexJahrhHV5wvXOjVqlzQGpFoIxMi8jOVamnI4SjjxFmKLu4YIZSlLuwu38t
l8Iwr4TcNhsL5H733zY/qG8ObIR4UJJLsAKCIQXk0tS9bFZUZcXie/S2KqBaPYpP
OY+k67LExuvdrlgkr8K/hSKqyJKB6tgfQn65XpuknV477Nm6c/9pwtAtl5qGgEX+
UH+OUI03TI9HBT22Yw7zNZ/K209JabGrH5jle+XNoO2jhAXXp4/fjXQy13wcCFDw
KKLlIYwvw3nZCk2TiuXiILFAPSGBsynxt3xXJTllGEFKksOyTd7TuDc/l7gZPCQq
vp4AjLGQT0/Ra2XtybA05cHlFT2Ep9vEg6vlc4bJD/CsUAtKv1g/aOyQpUxg8q4B
isMW7OM1fzWwCYw3fkZ54Sd1O5Ts1NCtVxTtZy/vlCWng2b943oPSrnVZ/2Esn2j
gbGO9uPcOZjSc8m2n9FAXqh/r06fHhUGSOr2+JSUOY6CwW6+uSYXVK+SHM9ElYyn
zUxobgCT9ffzBDy5mO13jyBBp4Mt4Qrv25RKavxAFhfsN7vMT/FBzGKiire+1mYX
l9fd0bUw1JIQXDfu3n5uL8n+FbJwQBe2xlXZkbj2HoTsrQwKdvLn1e9OhTpS8FHU
mXFxQXTJmjLUEGumZ/+5B6HFC6JoAh4tN49laFE7/n6Ny/gEPsJWIwdUd2z/2a7y
rZwbMp/Z3MJRvqbaj2bUDq3khkfhV2gTGTH+YXT8LnCoFUH74n0y/OuPljs3BEww
595+fDehD4VSmGZlT7ee9Ovmi4woaBkxl1dgxq4VtVyJOykZ+sPnPeNKRXLHLEhL
1sRijsb71rFGsLdcu6As/blUyUsOydA1GrQqkcHZjFofEW8hQPC43t8wlZI7NjZu
+7YjIhAr+a7obNGMTA84s+jYKZSFEfzl6T9GXiHzC60LjjhEOcA5dijNezPX1+XU
TFvMqlPhXEC109sZ7HvGQ9/JixNrFgTsT7AYocDM7j9HeIZsCeSUDrrHHlmgkUWZ
2tDu85bvI2tJtZSceBoctKwPj7GTN3wLTHCOkCz49tLOhZudeSWhuB4WSIBYjaZC
xrefxoSJPg0UhJJN9mw6FwE3Jb8CJ23ttuXcaswkwHAYztnCsg129fegjLNooaHs
7laLhV2Xr8f6nXHtdl/bCOswU+mK2lUt915WcYBh+28DT6awKcoKwRFCO9CPiOOo
3WyM9APmuSE/TzsWNc75aB/GfRVOI/o6/fPvt13bht52JIM/0w3A1ADzG7TLL+eh
nuzi5abPOY6SIJT33AcTHCZ6/XFZvcQnmfTQWkYYDHgM6LcbxepNpS34CD5abIBc
TN50ouIPkXVWUkSH+ajNott43WPJMaaVxDYf9Pt0136J1s9dNVrz9QF2czapO/fY
om2FrMgQSG3sL3I4Z47OTag9j/CiUjxJzryxA3VzlXpfmoOUKqclDryu8LkCscvG
dGi8U6e34zzPSEF5vhh8+uIbqSuBN6OBVNRpMdVCs/QxEkv1k+u9Qwtgq49/eska
5Pvist6zKdCAFT8OuyWzpr5WtivjXNB9ao7wbUVwvuI3w8d1ThsnJwtxVK8KRjA6
sJfDIPsltkEu5QKjRrzgHILku7/0CLKNyoSAFRNuoHWDDhmx0XRAwiIrUDRm9ZJl
qB5wvuJ3h0YlTStrIBegd13v+A2T2lc024xANS7chxStf9Hq8oKqFAy9XKGbz7Kr
zJSxlYk4zZbwy3+BAjJgiaQDLlRtu9t82R4bqyMY1w+WUP78l4oi3vNFu0bikDZA
+0xYIN1OYCsE+rhlHl7lwB3wgkOFDtU6uZmedO76IzDb5xfkeScY1LuTbsd75Kt6
fTWdDZBsBiNme/SaxdEyVo/fnBp9U5Fs7pR4mku2N3Q79NGdKSINxQSLEc2dJOlJ
sKYPLG6M/lLbmzg4n6PNOWd3Vd+HDQbL4YK7WIRZ7P0mr/Xe0SPtpHpU0Q7hYTSU
Bf5qgB1bKpa4hrA2AAJGM+Hb2owpHha1jze5pu4jUUT0K/RsJi6zj1+rURdEs4aD
0Dvkh32agYF+ulfAxdxb84XWecuU9t3gKNtuqb1X9YW/yYRgdfGBQqAJ3ZtiCQsF
Vo/fyQSqX1NmI1sd+tnstrxRMh2CCMqSaltIok6R4XvGTRHCMOLKAI0kOGz5z4Hd
5ZTEBaAYuj6Dx2BWJj78eXkqYHBzXut2ucP4axhCzD3aooGNKktfFYR4VszVMkV8
tsfH1xXPsRZ8SVxdBx4irlCUQIk6CpVJfrECalg/PjsiZ+qpsqanvRjdfF9fO58n
/6/02QlXPm8NLf6iEMvozFx6janOklDF1KQqz70NsiQIZR7jIecX5qMUWI6StH3Y
2UXqjLn/i9Z1OapbHKaH6Vh0HjpfYJ31UPvSezMmr4PBrSIJ6fsqR/eTvMO0fjuL
LpghgH37FhQHBB6YHmWwVrrC//ofERo9vYV4xg4ZSV1/MAtvhdml058atR8heuQP
8oYPjqnl55CSdjh78iwS+dsEysWWCIb5tetDZCC4IdDMONqz3qnSShRESR81pAB5
YgAn6uqurOqZ+0uA0jzX/xqVDdENHBpwCD/GUDRM1SNCs7yPDxq4Ywv1RZg00p+B
Lx1wNy9AASQHB3z0L6U54+XqGwSl6unD6+muH7J03r/P5OUEnaXs42WYhA+DW1iI
hcfAVRKs2Ub6FTwJxHsno6NhTHaYWTlxOqpn+sriIofH+TytaAcPxUItlkrkDX6T
4ETL46r7T1oBnXRvnsnLe8ZXHY5sfJfJmVRzLpULxZPvZY8nzn+qNggw4sziUC2l
kWGknqcB0ZcYYfPtOoegpl4cPtj/p5RoDdkbSCgYvVn3J7WVhwydNx5boPVJ7WAk
rH2q5CCiyZUoKirorfr0l/6rKNeMCxYGdJvih+zsL/IQ7v8GevlRvj+D+r10hOfl
1cc9XvzwgMfwV9dtNN/bmDuCy7QSwZjmtLO4Ez7StCa2bZfPrYBKYtlKgjZii3BS
P2vNQIVIeHgTen3uerIZwsZjTqGhIaFf/HD7255mczkAEioKEJysUYppNBDTfk1c
0Xu4QZ9oxghfZSB9HYKK5OSvhEOwsjXZc9dJ3XrlJHXfU3EeQ7971v5NvOCYeWj7
i2AoI36rOrKPZNFybRRhcvWcNZv14GW+UwWhxB/xq4INLTkpKQhu0o38vIcqT8/n
GBTgOB+Hc9fjW7V04j/OI5yLVOK5gDYFjj0+fbIbAp3z1dU54cBPqJjzM13EI5Ev
qDZFiqHN9MnWZDWrR0YRgVPGyRXfOGJQmSpVCaRCYjFE+RQdmxL5Km2yjDGntILB
cf2Fzoq009hZ3vt+y2FaSl5yG26A0udsAaM3tJbdqeiwQ6pHomGQiMBP7kadolmG
NXJMVr0PRYg7nzdJHBHgOnRsdvIJNThT3OBTSETwpiKxu29SMN3/fLKm5M//7eiF
9D7X6l8Xj+OYYXMa229ltZb0XIgwZKjbXqmJSakQ1CaARoOBtAPULx+gFnU4sx2e
HQ3NuFuU0CL36PeMrPooLTLN6uj0UMH2lO/V/pOP/40b4vttQjDSCSWA3mQODIeA
bTPcmFUnwNlnEdgjtns+G0NkMdt4Ef3ZbU0gQSDbS3wdSVDmj1OUVt05ZNsQrJcW
r0oT2VEJDVBG4bBbq2T2jm4U8RyCMHvoGMqKNyAN+ouhc8f+MY/L2f1nPJpNHEOf
a5tYKasz7gvhiKNmYb/KI3wqnhCCG77woiLyjTkVcFqF/4rAJ1FPB7yAN1oAdFte
U0FBgeV0MZJ8knI+KDQNgbiq/AgpZbQ5J1fNTu/3bkrOXo/Bi3fndYOrMHTi11SO
uNu5tILDAdyfys0+tGWDEyiU+E/uy+YE/666CdHSPvJ5eFzTgyxMzbXk+RDwSzgH
hAfBJMB96UG4WsjKKRHeoCpFvrvnreCmZURd26kXW8PwiLOIXCR1Vjcr7778V6mF
pNiGZclN9gf4WJIAmEgTp7Idi5JNoyLCm95uO4ih9hnk9lcTcE++MW7+kxL+2neg
r4j/IECQQI6r0h6PunK+fH6Eb63tkkLsgYXJqCg+AH9HhXqDgAlqHIRAN11eD53D
w6eZS7RcvDx6oKxHYQq81wCrbl64aABzilDfaoZZCEBI4n5jIdnQoslFBAyWK6n8
kDaOXenBVM2h7+qPDlR1f1yFB38L0UBZq28EWFVoix11/lV3dryIU0lUeF4twyb/
eigS39ajfYmd5E7yYF43OBDHI5Abf3zLvGVFnJNlmfT/e/VGdhnw8mPDYY9w8uEL
13nd4fWjhdlsEmLBBlr9pzDrkRqceomgqLo0wr0YGQa8SfMAO4QaWgfAbg8dvTZ6
T99iz1kXhZyXdjyaQOPTTqLsRPaq5XPSlSHpUVHreybB6mbccmqRM/k0Q7yWVIBQ
g4TjANQyStYlBwzzIvIz0GaO05XJNH1x0HYtJzStzAKSdjvMr1rj7+vtr516mc9k
iL1NeDKme7DLKjIuguPg9mRvS5DoANYxegZusR23hhlQiei1cDM4HGtI/fEYgFi2
Vc4xW2/3FO0X+dmeN72+z8L/LUNhecYkxAx0m8NaIifUBEiMKOS3MPfj1LDLFtsr
LodimNO3mEpKeaQt77977J0ENSMWXYxArccpq9b4vxAfHKb3krmyd7vbkD7RVbHc
E40E6SAJqNsIiKvgFyXNMGyl3txU++Yoc7KPJnWbTplwsSxxdKXMLPoZWCSG5S+M
a0jg1J+yAV1jKrck/ZLAxpgjJ/2G+FxuDd9PqqtD+VFXtwmNmCxhno9CwAI2a24+
PbmEHRNq+MLq4uBNoiWanvAhBNVa9L2TwzFmiTSm/AATBlz5w1+ma0hLvYgZ9iiV
e88seC0iV2oTX9F6AMkAVslMuAz/oTxbLonNnO5/KjAi5lbq69o+8/PARs6fGOKC
bk4pgySZ/hpo+Y1tnGuWLJKsHusL4oF499VQDGhP8/Uf18rGPw20ePgx5cGezjkC
0myFOfNhSFMNpMsF2QxZmPJuTd0GKALIbUU02bbpz6UqrIjVhj4wXdLCUHGAGd4H
hJkDRkVxkIhEiEgikNwFIH4o9DSVSdqhoUQCL55spViF9CHqLJMbUKAqpPqLwug8
TZ7jJVwuyJaE5rIDR0lxQ670+r2Gpd/Vs7p2QafpyXT5m7bEoNcAnJ2bTTycZtIv
GujWe8K7/3rpZGgGmnWEPES6VvBm2wTzOwuaFolj/rfD7GasfYfauzt0RKij1gLy
vgGOYWJi1uYOjcI6ZRLnfT3rJ1pdE6mbmDIFRefAu9Dk51I6FTDCG+PVaFP4X7RF
mcBAAu/zFk5APa+V2A6jKhCjYNV4QzV3rHr8/cSHnKdRe18lccBUgQKqbV7fmAjC
7jAVPfhLGtC+/AyhE4v9NKec1723+34rtvXocqOui8YrCxsX5ZFFPQaLJfYR2NC1
48Wk24UT70FxElrv2Xfyvg9uJxhD8WUSpTklcELt64F9e13DbAd+xuRkIBqVxd12
Tqz0lu13io+gYdKn7v24tC8msU8cCgkQX7Begsi72PgFIAZ75bpurd6WX7JTuwkF
tUVyciJUbGFG7zw/PzDahJt/WR4rPbRrGq3IN6/I36jq7iSZEOdoHfGm2say/d0K
oAg8TTcx0RV/cWPoS34YILqT0NgUWnDB+GB4H9rvot1fH8kR6wKAJEs9vXdt6UZz
NQQFDld1sye1lciz4Bf1d1KVkKvivr3cpO3UGCSy6Fv67kWIj8WAxeHhAYn0VpJY
NUFFW9x3cV1hEjrSc6JdkW4R2OwcvVyVoWjESj6ksHZmSbK/gVC9u8gKOb/P9cUi
RMJB/nYuISBsFGmNK4aJguH1uzvdwL7j1cpVR6ozls6gY/eBZJ3RjbTD8un5wlq8
RtTsX+ETBdAFJzoBWfQ1pS3AdxTt4uOomkFr2KgioueSJb3BKfo72fCQAbFKM8Ny
z4s0PRCEAxd254u1Bmgylm9nVuzeSjTNxlAaF/3Y+ib5nOq6SO21D968nF6N66Oh
rpWJvIDuFYRSBVfT007K4JGy1qoBu+xPlkymAkKB8j+OVql+Vi2+wRBTx/88MlOh
ZKEw+ygy91v/aMyG6zDPJ/Tbmvl+tnhjPbv5DIZkcAmbNL6mWl2LEw4HUaReYHPA
PZbZHsVjjP0dJ87XwQ2AsEYEonrgvsa28gX8GOLAVw5myKe3oBRb/GUYH7hiIq0F
dx/I0uUXJFCTt2Gszx41k8NvgUQE17MKwr4x1KFHXQE41FwJlGs3H1/CQzwKrDNC
7I978tyL6PoFVCWZC4ct0xlRHeCwZtJE7ZOf7zunfjb/jNKdfL1wl2bNha1TXpVD
fL5AXSkFLGzU/zVXQBX/fCiFEoUe2FwObBEhAPVxsxMSvBEqo7GECePyQaJrx4ti
FijMnAjRwMqWfHH1Mpbo2yyh4j9bipNu2CDPJIUD/kSUf+d/rZJt8nnxJ6HHIGNW
QN6ypRIexloEMVygEXuOjBovCnIqLFTOsYbNKp4cat1922YAkdeEVEu4nHxyI36m
SyrFj+XlafvtfNnvL7Ng47+R/bohXysu7q0vEWw5POOCLK531z9IRR7LpqgUZvDC
UJek0WUYY+YEvqg5nRebKbwhHPf9eRhKUYbH8yVnxmKuaZaTdt3pAytYDdLrYD3t
8uZW/xrdhITcuS8RA27tUi58KZrD8zo0Wwvsc7QO9aplgctwmw6LaY4sJPravmQr
Y5btNzV76134xJ81XsFrdoPT/p5xPVI4NodIfRXyeVcaFtCxygHnNV5FN7onAnNX
mhLJKe3ot1fmREGAbmswefAbAZEBeVuK48fzQoL0Lv5UUtMffEEMi3KNvOT0mrCX
xUljVn+Owj9DxH0TZnPc4SzGjLNFqGe2ACt/oE/CfhPnssifjzYFvrZLwbkDYCj7
uD3qWjkGNcs5kzEC1SyARC1TDlu47AgSrd39wZk6WvWQQ0NfyJ4ssKcR5DNfMIxP
OhC5WFApQyPMHmdngrwcW88i78Gz2DfvkCt8DFVqPNPLfnlDlA8zf3keWJosGBBo
ZHNfXskpeg9zqDhozZWDIXTClHCi/+6mtJLaau/MKLzD/8gS2usxwuuPQUBXJ6fr
Ixfid4QDA36CXT+SGwb11kM3KQ45kPJFr9R34GrZiaeVKEqbsMYFHtIii+HLAiee
9KdCpZprg5GX7a8rYPg/Ow76uP2rh5Bg7163yXyR4rPMMn586abtUWYwK5jozxJ7
prE9iFap1iOl8tqD/g/LVYZht7qrbZc3L/cCGQQF3DXF3Sivpwp9qCC/TJm+CYIa
R285mNkAzJ4xMpl6BsOaVfg2CITmRSeobdJIAsIBnqTEhCw3J3sYNGAfjgpSi5o4
3lJh4xCe2o5AYmVc+Fs5NDTSY9WlwNeXwbA/7p3WxgrEf/bS+SPeTcvCH0M5H99J
Vap9GZNRULfuG0kf4+G8zq76zUyK2xwrotror6jglZYWU/ch9b7Zp9qHpiuHWwVf
BVFx6tSi3IX3CxLD64CquVZlikdmZN51BjaF1XrhP119ClSoedmHAsnX8NZ9P7Xx
mqQTY4MHOIrL6fdjNAKAZ6X+2JljI0CWiAYsxiq5dth/+TWwJ35a7QfbjuLBeWdg
L+l1yUW+HTKd+K/rjA2inLidMV7IEDmy5YS9QCLvT/wW6GYBdPx140wtpacgoVeI
FYnPhl1WBTU8bF8LuHcnSdyw79nEycqJtE3/KMnoQbF7rOXBJrLlQuELcylnPgij
wgDGdxCPFar4L34cck7XgmGwHHALNQ9mn8ZRTknb3ysHAvgOa9oCf7jEZd6AQlR+
6aDHuweIW2OuVw42WPM8GaJG3/A31GHRopZ51okSRVLCg4CQpW2HjyiXRd4wugwE
giaeePvXpJ89g6fprBy7DvNVKLs3vgM2FIjDSJXpmMSNfe9jLdG8qYdYt2x11YQx
07n91XF9mDmlt7tUwIreiDx+KGiq5aIY7C/GpLcIBCL2QRY7j+jbyM00C2TOGftr
PqH+qq4TT//G+Bk00NYQt0LJ5JRSuIi4FN7OAOf5XloMbattCUa6ZzQTtSomLrp2
bUgocJ3zczoJxM/0wewr6Jv0ySdEXvI4EC1uUazGjlNvJziBIxEbwcihB29PZMZG
a4GOSMP5sgACADf4gQAjrQEiqPcGRJiDn57qraQckjns2FDWB/G4NY2wPOhVoub7
cnNmidM4SDX2lYbJDyP57vGNJZHxzslculHV4VhYgsirWWSkdiwxhWIbCrFbiSox
CYgcPKMyI0Vnr/Qr69hFlECTtBn28EcdMzYHBzR6wEBqxmgSzaG1v8BZR/bApbfl
gkUrF8qXA4iBdoWfgwmJ1u0RuLp001JEpP8cufzl40pQA2eFf8qlnTtf1GHpUaE/
gv8UvWd+mfWSwcVOS+m1QRQ/siOrX/dhe6V7M7RdpeyshKo4umYMVynkLivjsFx2
DajullecDNIkr3aOah4XSPbthlxGcGkoPJJKZ/X9nhtChbZKL5hiZbDQ7l68nNx6
ADULQxMjtvgSxNEs2HZ/LvfgmAJlyoP5e0AatNLI5Q1pR7gvtQB3weps0vGFiDIu
QsJG9vagKBLok+b65XFNsHjffAZOWTG5ENF6z6Zh0wYoSCtwiI04S+VKDBC58GTA
fc3sDZZc0u0YdATGm7FcyK2A6EkpnZyRgjl1OmVAJekfmja/KRVQ93I0v27mWZZd
f3deoy0dYtty9DJ43e28yJWAHcuc3jw8fmeILulHAuKizBHzre6L/MKDyqyPOtRH
uFQ4XCviRV8Vt6K3v3+dpikDckoZEbYF5R6R/cYgIM5PzOFcY1qLOQwiRahqszId
Y0JwLHwdmRDZGRrSNFLitZLGfBIqyjzWYU8VHQDTRRMB9SxexRFknVV8ug15uDl5
1SIBXsVmW4njTdXocwXzrC5MQ/Ru5J7MLrymeiJo68nIg+nkxsybt7JoKwOKHTx/
MdutdUoMDNpPl5tGQdzfpd4WzHcgw026aTx7QhJpbMAagxw5wZFA5k0vb2W1TpGG
MhGehE6Lzzpy9Ep5zldcBiGlhv1+87nURo2Qurg56OFyF4e9hnmkf0kvUeEVycB5
yaiMvS86RWQNfreUi2OofMNVANl/0659q+8DQlgtB9+aAGR17rE7oyEmhi+PcXTN
vtZzmkO0/q/9lBXyVMByIEb4C2OK2SYv3D8Wtxp9RETDL1bO4WxHJGvW7gwNJSiA
HT6A68uAOo4/TlkgMTyXq2EpcImTMMfM8OQMC9UH1Q56PZfIXz2V1dLaaRe+JfO5
6wXyjD1i+irfRYaq540LZbLatWDAdLMw4DXq9Un4/vGZAcY0WmYllKQTF+Noag4Q
q2hT5NqvaLGRWH7EQWHrcbgDp0T7pcuB6LHKMr+WE8MR+H8KDuujpd2HWqzi9cDA
XmhnZ6gfZ086+YsFyqmKCx0CSE/u6L5iGfTsDaRXNmJoz2J7tbB22etSnyYy6KQ4
EgF/6RRS7LKMsCUeFru4T7Uv7wsp1iJr2WM0aRFcbzRqtjvbZY4qOeimtR29kWUM
G898cdbF7fkL2BexbgeebV1cWStR2IBGq2VNKuJgdrv2OkUsJ0PojcHvUDewIVEK
Fqi28u+nxOmiMFWFOOgRYNXMFT+9VaYf6uHVubHe0aub5FX1W5o5x1xon9y4ZJzO
5yXgPM8k+BbcgklQRD7GM0i2SKWp2MbIKlgSPtuo4DW26xKuo6prvos6/xgVp1av
CcnYbMCraquPGWD0uFl3Z1dd835fB7zobts4rR2D+20EQMWIrVujyzzbNjh7FmYK
qGGTdUA81ji74ALaHpeXI5jpjn+J1D8fjwBkt8Qokysaqf19EXoUmiLp+xkzMVQF
hrGzfUar4VkSZeNPYjzCyDHn9ANG2MjyQ44A9PyMhgcXljCsTTBBb1zCV0i0GIMN
fNrurOB9Qzxxsd/4AoyfWRXu+qqPi2GLs1xlff/6WBT6wOgLiFDJgvmaLxFYtbrf
TEe/3OuFm8FswjENGNT4i2QYZS+CA03tJ/HlPEm9K1uowpLRKhf8uirtEAiJuD3u
m07wKE+OrBV4g6zForxPOwBZiyeREjRodS0+i1VharaLKU5o0MiAJJfQzGxt+def
JRT5N2sHgr8t+xrROnVAmTNBEtDYHiMmczqXnmgKDp4o0uPw0KKDXy2KuR6KG9Qo
AypTjb9GoGANAtdZaiJQ57DcrVl/kYHtsMw3tWtNPkZYJFmNv/rXUtRYnDzDauMM
aTabO5ocwZM6FUB3BCuMn5YVm4nKa1CHs5NlJ4CsS+VpGuPkcNI+5hDh8DMQG6BQ
AuXPewKCtVUo9QuzREITjBdLbnsK5wms4jx7hQ3WF7Dud1aBJh62RlIvAvszQv5S
jzg8Oakr6+gBnvuXuPu/1411aRKhW8vfGarTIP1MrvpiFtyp/RSXQbMntlYJk9Rc
gMKMA9e+sv+t0qBb0YBPkPFpK6xWANZIvdWjtShtVOiaY6hdCUNxsZLdC2adH0Cy
zJebl/VAkU+AAdCUTcC/FzfCA5UzaCQPMA/+Vja8lyJSm0qVWoxDTyHynJsw7D0q
Ypcem5omvYLoR7rUll02gY4Dk6aOSN8yZLsnfOUNPht+m7Xca39hsFCpEWNdkXk1
b6QVS99myTIs4ugvztyTAXxIpFoBiiR2s4O7pOaDeGKXgFm8BVrtlEB/GyqItrHl
EyiJfpfYLkFWQt9LFMstNBLRwBMpyEZcau+rAjey70DjdHZVeOvcOCRe8Bx3jt1O
dSUmXUDa4Hp1jboSBUgy/EQmssKPU8PNPnNLKqkHFw9+y1W/340OcCms7undPJy1
pV6fxA5AwuX3M5CukDz3lt+Ojp1Z3x4bjLFn3O3b1EB0wfgwPbOOPt5N8mHflGoA
8H/T2y2JTI41TLJF1+4gJmL2JjmjnBf28slTAC+CH6iA7qbF3PkGjHZlwD9i08d/
Y00AZdwBF2WlUAtTClYgfSGrAogw7fquQONm4WYh05FmAX+OV4mTXTPDg1GbY/WK
NyCo/PV2DRomRh+mFqthJyfWeOD1EiR9jujZky0+MtNOj5hSdtKknP394xijbTtR
QVgEIaDqfv4dN+jN4nu+YTTUPPHoKdh0uEr7Wfgo8lVibZNIttxeetc+RG/NAOYV
g/QDN9bjLQpu0/621BOAkCE60SZR1RPXrWg1Ycvs8UXom7vTjvJQ7rwTFXL09efR
LmnULgKjYxfZUCSZdNGD4Yqmggf6beTlAHpSb4kfT2HZY7V1gYHtmk3EboMxV3/6
vy4nF0O9eROEIL8c3Lrrq/1Chl5rQjoHIhkzMMSQHEAG3XSK2CwZjJt02CTJo+vq
JD50lH2MsaHxfHW7LoJ+HnfIvtRc+fy7FKCsMCb6vFH1nWxPypoLotAzH3V/5b2j
IE+JmSAiRdgNVK+wALi76d/qv5B98kGeffuMtn3/kmBfS0ioxQ1K4GFMJNTLi9AV
3v4JBl6bPL6eahi8LPsFdMWTK6kGC3ybsj5uh14gWsgkDVvDxgm/0P6UproffB35
0yPHVIy0eoi6dzYySPHKuNcIqsJtyejDfdzGSJ92iweIQAdG5dd3TwzA7/Ex6e8h
KhiJGiZBJg02fad6JQ9iYMJJzHz83jlRNIpYM9JlgYudwcXlVE4C3ytcv/Yavija
+3XSiBAHlPTbZz/C6+qWve4mG4ua5B2fnD/ECEZsGdlsAIfw6Wyz7K/xubqi+RkM
mZHU5rQyQdDC3f9uTASnKMKrTgJ2+nT2rl2HqAoLsjyi616PrbP6mxCuYe4khvaf
jKU4Pdd48T+I5NInkt7NNVL3Aa82TWErg2A6ZHY41nNa6qzI6+KIn0xbvFq40HAp
NLwWJjGZYS82PLWK0OrxWdsIYVIt1sQ7iqA6RkF4uXvhrGeA6qhuDhujnfK9ARad
JQc4vyHgAlgDKPJEdmFEWrX3PGSp+mqFLEN/B7UKbD/GIO7NxWAusxXH5umaH5hJ
n1TnfgYSQlrir9X8OvYtO2oh9rkfw7cIvgx+n9MEBs1ME40l1zOKVZxzfivix3mY
Ved4qHaDYND0u9cx/ILFqZf/VBjVe7xX2Q3iBdSpS4GJLqVI45MSXXTuMdd9ScRH
1akKtn6W9BVoYTORQdYETZ1pjcEpKH9kBKwqJ2jhBFYpw1yN+lvg92f9DukM4dSa
TTjlR+x3TEf71UR2GjVovi23nYecCW3fzBiMKAtiw+zDi73pqOqqyvzBroTRUkcq
VmDM4YeT6oVDpy5mn06LSVZFnN6oUr41Qs5ji8YuK3FM+PVKpW/3L4fAO96EI/bL
j39gSV+JoPgxMz7rbJOuCoSNs+L2g4CF0o1ZvXSbWyVoRwf83a0MHp3BvmVou8RH
ohrYyNsz6FWNXc+qRQDQUzI9YRjeSoTNWQLGeUzOhJWF5cL78KpKblyoT4c5qMfs
pDbYQo+5uQ1MeY3ayXytmwxW8Iho4eTlnNDlnER3w5vTuLhxnrSoksWoIhJJ/7HB
BwexrQpSTtRthI7Hhso6Q00LZBnKYvd84nBQ0qfMzxEUbM3EX1Gu3VYUJGd1ynj1
RRFsl8D1qTh5DFuoR3QB8qrGJbUeusXlUMeZy4HHveum9nts7N//9zIR/Yf15qCu
gQumI8tnN3HekWKg5JH/yvkedafO9ttlvg5qTfuF5wzv4ivDm3BmTONApxPa3XIh
swwThQVyE58qaBdKx5mUVa9I9FrlY6Y01ZYNNIcWPC2obW1YcNZQiwLbr+y1mboR
BScPuXHi3bKq3QYfND4zmwcTTJgr+uZR29ARR4kEAcWdjbgkfNpuyN+DduYZreaG
rA8Fq7OnxPYcUf3yAwe27TIjVQ/X6we0jZiswKx8AkuKTUVkJb+0hH5ozlrUw1WO
mTzRRPPJq46E2GN4lLR65th6d3L0phEvNFreYjqTSNZoYTJv15UA8u6L1VzC1P/F
dgVuqUFV3c3+J0uc3tHok22SbtWIYTEKl82nGdH08zRq1Tj0bTtX1y1AmIT4jRK9
NmSHZvfZV0jhJ2kQ8bdWHkG+D2YG1fqiqnM0ryZDD3UQMP1TzKm0H/YTdP/e6oZf
9s8iQEgqTjyCxzNEF/6OYyfjVj+J+VTkg58DphQZSs8F08QKIPMGNIXoBw6I/mcQ
zU42z+ZPN2DO+8NTM2FctuX22Lj/fvVhigJsOylQhmO0ORH+O47dRPMgzoUhMR7+
w0p/7fFFh68Iw2pgajNjJq/ctlYtgAPZEeTXQ/7JPLF4D1hi5ZnppoERcXU8sSFr
QNzIN+KZ2Duu5twVLuYELrHvMGDOZsgQw0BnsSGKPixTI3u2bgclsiBkcztfuswT
tPZQarBw4TxBXGfPO7y5H5ZPyVRnZzrB7uhLgu9/74eoUKz1gOGvJsCRvNZX7FPh
ry0kkv8ZWfrDkAMto3IItNzbxAaFkNDDrfQu5szjtKwskxESnS/6X4Sd73N+pewG
lL5GfPAQJrgDY9/dOx18H4mn8SMUVKqLHdp974vcuPsSV+rtF9I8IR13g3NcmDHh
+2zUK5tNSaNfwF936aUypvXBh1LJjFC3SMd8pMcplmZMiz7hPFLZGnhPjVU9GMF3
WZuRZdAp5u9eHc+naLF2qlmw4JRhQKrUzWSEbijil4+IQk8GvocHxBr16cfz6IkK
9uxuPP+EWEzLNjPboIOlJ6LQSLq+EoFNnhLZBbBny6OQIV0kutqi4lkOhmK8B/DZ
OmtKMZ2+/icrsA6yvXz/42Isv9A5qBwYtbWWoWylo16Q3Gv1B5Y638k7P9qQA7+j
xO59UzxEDHp0OzDMqn6y+eN+0h9fqgeqnrs5SELXFxhOQNBp9fETF4wBt9GgoN2H
UqzxbtiGc6P8p9XO+HifL42rOwbgQy4ivTto6Qhqz/lDYXBx97OijqGvk/pw5sH1
c0WuJahcDNbHrp6vMuDijaZu696KojDMCq8r10iMvLq/HXISrv2OhMTG5BVaYzwU
dGdqu8lXVP/VMqngOTpqyym/p+/T6ON1yJmHLWTPFxZdGrDQlutbsP2O8toMEW14
6nrMonEty4d2hoY9AcTiUNnYPM+kvdv5Fnzz8buhJVado56nrrM33tRta7bMtWHf
cpkB1Zo6kfkJU6AytfUx++BxVNRH1PO6tV01u9xvh0yNF6JIlgBMYq6IsrPuC6p4
62FdYbUJLKUQ0ntbGDJ2Gyyxm2x+SY5voGt5Vf0Vy6VXZg/ZK7b8Fg3j8CS+k2QD
HnWybu/GWUgA/smOyR9rDIozYUtdkRU0Jmon301wV/au9ZJJYM23OZEu+pUxMMC3
//PABd5W4Sx8h8Nzzxmbcs0IfWVcUqMUsXK1etU+yrvyp5EAEhaNY0X0SPcIcSIY
ZZN+UILGRu3L5qMpa6q/qhI5MhebuAeXt5WedrHEDgXBuv9KH8sATMTIpi8ZdRXA
jVZkOqCYfeWHU8dqAf1sRYPK33ClyKoONUg/RVoaQiwHXRlqORU8KPUpzH3uamcI
KgiAEVydzRO20VUu/WssI4HFXgnrd+VFq1X7z/M82WKB8UBHm35zvD9giJ4aM7zr
0K/bwu73BFlzDZo6XkTihrqkdoA4QvHmNMuY4/mD5aaK4ke2rh0P9WrbHn585p5R
jWP252/qWPFLVd9c9WbrPiVuGS+KdWFHi9Di5a04gHhBs9I6EqVPj4CZIc8ikk9O
zvpoyGVbCmEMvtB/4AvKW/GiFMPToDQePoNMXo32lnOd5jQeKceFCDuZCrfKIL+w
vN6g+XpoUv5uUUPYU3q71cqNaOkFe1HoXxZQARM1kExqelFqc74++Ck0dYZRCsAN
ClkGDDZHb6BBxK1xPAUDDgBWq8bFEowgudyVpDdzkOLdNqOpn7JXVkTZziuCnNdN
Z53Du9E8Pi3whftsfdyNzfut5DJ7XMSCzFAewFRRO6etBeH3E6qgJJOJhh8ZvT+8
/bFoexe5st0XDBz2GjI7m6WKoGFkMbbjpNTr7w7B9lOD0eErHaOAKFjMbIta2Cjr
V5QTXJDX8rNL8lsSL7hgKKMTUgTjzVrMrtFlir6Fh28=
`pragma protect end_protected
