��/  ����_�t�ɖ�
�������t�_y�p^$�/R��T���{ƺ-�T[�@�NЩԿ0�!|�'үJU������kR����gX�Y�ŭ���o����^��6ҷrK�R��8���%.%
�.���Jq�:��C'���RÌE�����(:2=�}����Ԋ����H����#{@��)	�<�:3eE<�᭮��yJ�Z��X^dݭ5W�!L�cSa�&,�q��zN8�[�cӭ!��K��,#�U�������k�#!�ܼ�jH�i!r��$�ۃ7�g�ۇ�P��J���F��dN�[y��Ov�4�eC"�Sd>S�}���/�;rȅ�d�a�e_�Qx�¹����xc�u��S�@�����w��n��M�֮a�G�����U+�e*���'V�!�}W�j�LRQ�=CpY����<��9UK�V�"��	RL� ���a6�]x�_iX�m��rʙ�'g.E3e�v[��fS�@�	$�%���U=l�\�|���-���h�YL7~)4����x�E��1���L�W�L�>F6�_݈�7�2!�Γ�j#dC���s)!U��tY$t�lE��?7�n(L$�3�iB��6��s���˶-7SOg�ș��,�Q5��Ɲ���#���w�����g8o7���8N�$K~SfdI�k2���dR�p�^=r��T� ���P�)�q�e/*=�^E9����Z(��V]�:[.��7��d �N�<�湵�_k4C�oBG��x ���34����|�����6p�8��ܩT��yW�=	�b� V#�����(�Bk�w6���?�\v!��q�� 0+��y�ØVi��s�}�r�yf�;�������+d�Fu����q�s{���I�O�4w�*�����a��n)B+LQlu�(K�J�
�e�o�ʬƯ�� ��2����v�G��n�fnW�� i�Pw���%�W�
�u��Z�-�m1�x]
��1�.te\�JW�e�i=��%RR���մv� o!�<�CD[�p����Su�Ӵ��pJ��3ō�k���cOʄ47vঅ���E���z��لS����Pz0�T���sgu�H����.��Qq��oG�T�O��cy��N���������Q 7��;� �U���*,X�5V�MH��X~~��'��Ĕ?��T�?Y�H��������J6�[0ٖ���M�6'�9��K
���g5��l�:E�j��2��6�x�L��S�Tհ���C��f�B�І<���PәF4�ܦh��3��!�����F�v�S�]^��ؖp�dUW�;w!=5���|�����HE��G��l��ј��l�� ���)���7�L9ۋ���:����̱P$t��2Oux�́�e��!ri�O{�� ʅ�t�ǊXt(�$�m��ߠ6\���YlSh��6/�|Y�)[����
�u�C�A�_��z]���G����{X5!Ï��K��'/���A�Hi��S���P�E��ܱϩaX�����+�t�"nk��<�ݨ�$ɫ��Lf�Zn��\��&�0r�M4!(?�`.��S�~��.�T���L�Iq��č���8�!�'	�yK�Ћm�-ɴ!��C� �2~8 ���# ���� �	�8Q�ќ�AEΆ��cQ�M����e����Axأ���^�
��\�h�y��Zm�S����B��,�%k&�g���Of*[�m�y9l��e��,�Z��-�-�b o�ІʽW<��Pկ������H�F5��,Ni^�%�R��Z�H�Rlb��]?��	4[%p�ʺny�+ea��05�����Z��'�6��|7��.d�,�����f�ݒ@K��Ph_���<�N7'L�U�����A�.K��f�n�-��r�D��P֙2mc���_���i�T�������Dַ� �|s**���7����1��Ҏ��-�fV���[T����ŉ�`�!6~%��=
�V��P��2Ђ��=�>q�xGDY��U-��+/|�:#��Bb�]yt�E������~�9_kmi���l��~*��XY�B�:0��B�t}N��n��K�Z��,�����Lp�q~u����]_��Xms#1��e$����Mm4��<pU���h�GKشT��W��uF;&��M�ސ]�l��%T��`EW�ђ�9�{�_�u��ӫ�!�,�7��(ĥ�[��硣O|5�,�
��>r�"{�0��(���i��|s�[J]4`��s���
�r����������x̛z�W��P�lP8���@�(�
#�ove���A���yiXe.*��/r|�B�V{�o�V1�1p�+{�W�����Q�(M��ɨԾ��-��M�Sj9���k�Z�vÒ������,�L�.\�EJ��F܀���(���� _��!�38�cԄ�^<7t�]�TO RGܒ'���z
&��潶�b���H@��3F1�D�ܨ�;^,��|q��RQ�6��j�9��������a�ڶ�����r���_�F0�i��n)�#�;c)pm��ѩ�< 8�>z���Z�'�Q�d�t+~�)]ĚA�@����r�&?���K��	� 2ؒ+���!��~c��/,$�Abn�i�!C�E�3���.�V꙼L����q}�H�c�7�t�W�����nvV�.���X,�2���u�%BY��`���93��Ȇ\T����5�@\�s�`6g�h��>�?d1�1��D����lsM�y�,�A�P�� i0��ښ34�u&6Y��K+i�.��Z�&�@����-��%�����!!8��15'e�%=s'Ȃ,?�����	&%ږ�8E��}�MXO� cu$xn���jeR��vG��}��<K�����HZr�{W���r���c�ו��������}�T)�H��M3� �A	��2O5�_��J�`|G�5ː�/�2����];}L����~@/4"���k#���\��=�O���=�<U��[�����s�4��qMg�2�Jr*�|�ۀ������[�oh�h	��VRBt&�Ƕ��a��U;���X����i��C��6��ށ 慻 ��U+���9�����v4��"�[LK����V��e�<H�PYt��bhm�p+Z�KL�HI�v�`��P��u�>ɂ���j�/�؉V��	)^����(>|�C��m������?j�vS�Y5P��Jb �A�D�\wD�#2]�н�D�$�?[� ��V�P��V�X�:k5zb)��m�ib��0�Sm`���q��޸�-R
�g��(�2�ÊwG�+��(F.��)cs�h���E�D7H�^���ş�Rҥ@(\y	K�ֽ!��"	ܰ��mN��F�K<�\S�P�i+����t7S�V
�)m���qk��PVК�H���b>��
o��r~�G��,+�#��܍ ����B{$��Sq��S�E�7�_Ŏ-[_j���d\�#�\���d8�L��^���]e����} e¼�ߣWF-�&�>��e��]X�^ۗ��y��<gZ)Љ��M`�W��n��I���{r���
�e��	x�F�θ��$�@�{[ӫ�������;�+Q���\��85���!������,1ک!Y��q3pݦ;�k�𤙩ȕ�C����IG���9�v�����S�7�;�@.-�3`�8�m��Mc���h ��p��$�viz9!(� w����QL]�������~?�~�ҙ�Wmx�G&��f�l�� k���/��x�ۣ& s��L�V$vEu������x����v���gt�4*���Ҕ>z�tJ�¤�?��W5g�l�U4e�P~j�r��B۷:���uM�'�=v��4f�;*�z��deN�H�ۣU�.&�A ��q�I�2�`�(���3�0�i�����I�mS��۞�z5JŎU�I��y���3ng�K��o�/���j�mc���_^����>�k�	��uFd�@��.�F!HPlHi��	���_����xz�6�;��^�ڋ!"f�k$GG�\F.A��y����<l�e��Xz,.H�D��p?��^�_���!N\��ih��y�����_��*ˋ9�L
�V+!!Gv+Ca~ʱG��A�iߨ<hlS�XDƿüq���)�����}�*�jbw���JH[7��)Ø��mZ��G�C���i攞
�^���}�F��v���m�,*��P'��#,4�)���.��mג�z��y|���0M>NI)�}�P�#F7�s�Ov� ]��/��=˳�%�B��W�i&s�x�1��?�0y`(v�e��~��խ&@�ydQt�%N��P���t�no�-��A��U�e��6z~厔��{�J�>"�+�����Uk�~WQ+��Hd�1�`F~���-��&��*Z�5B�P`^5�����7��4�䘲����q���04�$oU�S���8��|��i��Aci�m��yV^�V?n�A��g�u@��U�E��	�1$���ErFzT�#u�$ɬj|,4r�ZnU�7jB�XK>�nC�=@<�P"��)4�7&����z'�m������R)'���_0c,"G`�o����h���pI�|

��=����X�(3����1�&������\y]�Y�0 T�>�l�ࡗK$[���1	(��0'pdr}&]�	<+A�;m�������$��Su+����2��[U�I�{����ޞ#���n���w�;x�;������"�7*���Z?d�MU3�0�л���̍Q~w�����q�Ú�8���&��=��܌���럨�҄��A��;�}w�Ne��&�I��5��<,Q~�<,،Rg<ٟ挔�d��J��q��]��(Xe�-9\���Ծpr���^2te���hS���q����Fp%�BZ��:3F��=��OK�ojs2����`u�h��9���[��S���"�e�
0�_ܣX�yH�>�7���ho��)� ǃd�L2�5��V8�=ǥ���Mq��'�R�?�����7��8��}�#�C!O��GI2�/�*�<�ʯ�oŕ`�(T��mDNk�N��$4�z�F����+
��y���r�1����tۻ�o�|�U|�����LRݡ�����+�����I��	��Ù�U�"+^�#"���f�2�4r} �T��2�K�.7�g����X����ݚ}79��Py`��[/R���=m\����%\�<fo�hz�B��}��W#�Һf���H��Jh=�ʣ���m��Gwg�u�'�L��y���*�bm����(&?o���S�}G�뫢�z���e�-�-`|"#�ګ2���g�J�'1v�)�v[Qp#��RQa@��r0$�:q$���28ㄌu�C	2"�)��3�*y��j�`��@�C^uR��\wOY�F�`-;�ȯ�擛�J٨����Hou���w�w����F'L� ��F�w�]�_�|�޴d ́�W�Yvg��(z����c�U�k
�Dj+���7XVV���E6
�2I#��0Ն� �ڇV^�囊z��-un��#�`�P�����!����~u��`��70�lFfX`ʺ��0S��d@��4��,��L�X��=����ǰ3Nv����k>]�K=b=�?�a:[;���Ov)�v���u� ׵�:���?q��Қ"�o8�p��6���Ϥ�HX�ҒqYF��wؖ�rD���@SɁg�d�~�������ȺFho��}��L�W����;�ʻ<�	����ǩ��A�J�VS��ަ��7�Q�Ʃ��E6��F�?���"@P��^