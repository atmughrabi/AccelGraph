// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:02 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cLtAu5Bk1ChFsXO9njl4FhsG7PfK6p2jljnA7Sf9gLLCg8f4Kk9uLlWNx68oo+vz
jXuLogCgAHER2iuAn5l/j7+3UasHl8TsWmY3/WlPqce+3buCOT0H1vahd+e7M2R/
/ncBcYAMBbV8c9A+qlDVpRUDmBjqATxYSr2NVoxghOg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21472)
tKyHYCptNOEKG4CUPK2brhzxQtJPDy8RTtsLmcVbYzo7C9wVGqAQRcujj+Llmi0o
0dt+kXbVHp021FmNWutTIWDtnzi5BVmghw/ngRTz6Oj4BZwo60rnqmZ9wk8SPlVN
tx/+pmen/BTFn613180oY/RJj5nLZWFuResA8OflV8UYgGt2+BDOjP4Ul1r5ld/o
eKbHM7sglNYdt/myZ3bGmcVDl2mdlFpro2o8Z6SZ383o2gzd0nUW2xZaq/Khlvti
SG1yZjZsdNNfA8KGwvYsyxlTpiWQbZbCpYTJkzLtBX1WOwQMjIBJGtuftwvZi3Ef
8xD65t4sqs8nCRDhKyMTXGbXgmSFRW6NQHCSEdGePwTYsU+XdVVNn4nxC63AlG0z
agtfZvG8Zg9My/SHprTlWg3Zg4ZwexYQEE5JfzjtgkYw9tLt3e8MyxB6vO2wEYZ9
Ylcotd0GAH1r+/jn9/KjV7+DzsUVyrBUQ1TFOzPACPNi00xjOTk2NkQq4m6nZ+Z4
ix2uFJ/5yg3N5Os/1409YdV49VnngLHOer3o/jJLRNiirx/7OaHOIZbPri3aeQ+T
/ttvBQ+xWNzHLqgBOkUBu6GL9/8/aLPUL4Rw3qBFSi3/n7Ut9CKEzhpuwQIflO07
OiwdovlbXdO+ByKLJ9EhPAvXRZ8vd1qet2EBoN3fiu8nf5kbPbfqTxhp3HajFvbS
BlKVjLm7VUavY6vsq7ubigAftXU2rdvQFdV7syRVo1D4AiIEtY6eh5TLzjquP1IT
J0P9ZMsN3XlF+Bi7V98NYrLQQ/D77OXrbQA6Yp+7p+Qgz1LJoYVj8/5RV9ug3ad2
MzslWMBFdkTZEHkHy9YvBF8AFVXl980GZ8grLH+2lwtUdIJ/i74Fb/H1e7NiLuR+
Ezb1cPi+5D0C6WdzDW1cmAsQPGmsVkuYQsi/q7H+VxNu6c8MDnluUP+XiZHCV6L1
6RCkomoUm9uC0eX1dyPRRezuldwTycZlD1Tf+sXtLV5lb7F5CSQUh4kV0tmzg5Tt
7DXMmK7lb2VfQl5jVv78Ozyr4C6FO1xs87kgiqrGSWZzy9RzMhBIGNQUx2SSMsMB
4qDWeT/xz7ho4ewXuvXF7KySGfuYozEbAZBp+LBtdEiCGG8EPtuaX7LtbUHtHPFx
ZZAHDsGQ2hYjNiE1pzd/hfT4I1v5HlbpdQwXTiZmjYbTNQzNe/kgNxaC/rQyXL3j
nVaI2Z57u96QSlfzVaRHHz+sFtYDy7+D42RbcX98udumKBFjgwo1tZM7GX1YWPZO
cptxJAM786A2xkXF6ra2ZXEbyb4P1fXQdCrNnM35xP/BD7p8VrccJ2E72+S3zepT
tAOZCUMPHzoDmN8No8ZjmtfbQ8xXhmtO0dckF2Rpg5Ub3cb908T/Qh3qgwgoUCwy
rBLY/L6LXBTmS7BCyU/uf7e3aT01IyAMbE+coB/DC5M2zUv3IHZFQdghKGpSobbl
sHOo1oRIAJj4g6BeSH2CC87lNoIgyik8ivCTDeF0z5VW4P4yW5fGF/fhX7FQuXBc
UNZqbEBBq9raS9cUxpGd3GPKuJp2uM4uowvkT6xmP7EQJMMJ/tZoykbAB1ResiKu
7kCKs72/Dawme97iCBQnvcT2zJ4rmuuwI8FrHXq0lNZdWJe8lbEnNp/mJy/XKVBz
up4fGlXXiVRco7M3WEBk4Q7uYhMVZEnE4IKtkpGkhje+GYG57DTtT540oLozqdCw
nnI4ANXlfk9DLQW3bNcY7GmuFuGcYQyZLk7rvAP2dy0pZI7WESRyT4KBXoPAUmKA
fIBwwK9PTCJZx43U0+cnzechX8WvO2DLnwFMQ9uVWQMA7UpE5KrtVNb/+fM2TwXF
X04jXuoyeUUhEyiVih/gNpF4LBIFj03EW/CXLFqLUXqt/lsEN6AKrduhboqPWekB
HRD4jJTUZ4CbtpI/Q0JHIDqb6y8waE1YeOL5/8EGpUeXTRlgq+jHaK5Av09wN6ND
wOkEpkOGXqBGbrJhS8/U4fZICWsAuAaEAV6SBi2Q8tZkyyYDQ/kD2a3DPLkn/KMd
mgz1140fLqPOGS5ATdK47hiWLV8rkFpfh2FRlhn6zavSwFNetGMq29JOb5Yv3vgI
v93nWoit9IlCVg++m/yqxbkgpds2NAN5eByDy9fubPjYPfdagtJCLcLNF46aKvRW
PrmZ+Gmw6zlSmDruArU708EwTMF0gTya1cPHuRoaBJ/3Ae9KcmaAFzdKwNYacASO
9YKbe0OxR49MjSIKksDyConHa7x5TQa1lc3MJ8SZSFwwsRB4ZaqbcOwaelN9VNG9
GhOzsb+DKpDlZ5Mw67wexWLvYVlCGEkhNTj6gzREQj0LHK5ksk+T+iKR4gxOQpos
xlh84HRk6g/ozy44E4g5Hsdviuz/wFqj0Fk96CutHy77lnjxlh7vZGwMn0daYtKU
ZlZKIXaETwTSCU+Xuw0AShdmSfD92PdenMq3ChbbtgS3hOLV1JcWJW7BWns34daL
9olMJhsHgYIPpdfVeOtdm7qwFOMxjnRnRE/AOhmS7/ZsvxCaudbm0SUoMs3vcCvK
oWplMF+QKr+wzu9KoaVTXowyoLMRklU8VWtEOVlC0WMRgRrwBttwEHu+1ePlHWOa
4RE2to4jmV1UB2fysk1lYZ4ycrjAsEAm3Iqs1XGfwyVS/y7bq6dSa9NBTg5MC49N
A77c6LmE7VypRnDUgRrylIbYe+nzy8T1YPE1o8e7jfOINm7VyoZ9LpfHkpB/Pxzk
CtDpN/sHHg7hoWcO4/uru5AuurZJD+cwdUb4Zidndr6kzCDOxq2HLh6pDSpfsyl0
rJyVDDRBBzvfzCB93P6IlRZ9EWxeLngpo51JHLx1uTECf8rMrjw0NH/ZKkXvEONi
dSr0f3unmNdhGxV3ZFBlM5Sf5/HN0fif5hRGBGziGfXB16JIHUBl60TkPeI5y4cK
Bl7Er4/shNpOcts/oskogCA3jZUD05DSCuaDwiYt7HzVODQipaUNqIyuJAObiKkT
DIwVMwZrvzbW093SYB5PxeVZn1ZC8bNWirgZNKdOoooELCdmQWsD3MT1B6KzDHuk
aN9THpkppGhj2lYk208/s16kV960AS+/CgyNEXxbiD/KK/GWlF7ACun5Ru7hhCDf
hRCgrxIhRhl+RZAel3SyjwB29AHLVa6U7v4x+3ExwXcTxNMI0a4z0xqctM17jcIG
Yl+3igUTApMQ2B38EDQL9lxNbA8cRj4ito/0XMojBEsLoThVl8HrRM/wtRiDC6jg
wpWezm468AerQs5pyFQ7xGu4IRKJcmh0fhH035zjJLha8sxoW/iRoMbc0lkRL6XA
UreczBme4zLRcmTfFPOgvMBkTPWu7c4OfKvp7le0aiUXSoNxbKAniaHuRa4+eOLr
m8MvG5+r96sbqOMcm+LqBMg4BFJyr1IH2JtEKgQIcGYHGCX3Cn33S4F5pu+JZmMj
yZN1hZcMxEF0qyx84Jc5YzryrHcST1ZoUf2CkXcJgaDMg7GbJipUpyzAuS/RyKNi
AXDCku0aZoSdZvQnw46UN+b7Zq8vFAfWWcn0qJgBhqi2WGSF4SyZoyaO0M7gWF+g
pMGqUrFfVJfI6fgDsWgvl26INKElYsoZtDLWIOyMXWrcmyMEky/GD+kG4bETvfg9
/ugYQjhaN04CD/pTAp/Ioqgr/RWCrc7ooxIK9xzp4MGv5qto40l/n3pAEG9vRDZp
MRffz0Npcq6CSTA4eem91hTCfUnbI3nkdxspU9qlovecgTqaZTVeL56np9rHzbtH
+dnzqExkJ5Fll8onh00tUabZHrtp5oTU/sLO6G3+T4FLpVk1HnAPsTsv/KTGzDAw
KrmUMgBS8DI8IxKkJUJJ5yPCy0fqtb+8QNXhnBpZmsTk9XKyXv/nZwBpIELihadn
c6zX6hngdQUlhOa7S2GL/hpEo1HaPG/hMCYYOkqMIzKQ1WN4j/0cCbd6LJy/VXkl
FaUFyveGAQHQ/JOIlK+I/gZFNyaRRWJbiCQHcaTuYUHOg7Gsch69VXLlEMk9Z8TM
ucXFHXjcm8apbNQOAB+lvWgaKfo4ixauGL1Tpp1L6QJ+1nCwR25dB5ws+lJtJ1pi
l+hmGmE82LVuLR/O17Id8eqJWlDUK4WGEZxmj2jsVv+qcUB5qc2sI4aHUlivBTM5
qFCtOg1Fq4jsJW6sde4lzqGRpz7+ncaOqelad1vdnpBofy5YoQUOmm/u7+4JNb9d
8kRiMMo9biosl3MOn9UzGjDVlACB5S1vQiqWTtTUGszHg4L/RAqRbLaBveosQDdo
fAkSzbPG803QnWvvpcJur676dtEdHaEWjUwjzo6nwjOPxe1sUPJPYiIXtIu66xPe
lk6mHk6ReAuKh830Mbi1v/UZcqrvZPoTjsYLTel5g/gAXHf88xq675EQfpZBTCgO
1NsTcqo6L2cZ/rhlcela/R+u6QxcFbcRCL5Cn7Hen59p4EusEoEUtZEAE9c0eWGL
oYAjPtY9dLoiYx00G0TlQXgO6Bs/9kvKL6MQO5Hch8iQw7UCyuOt+SNwQOUP56m+
3RMdK0Yq0br0WkvdgcKyPi5FlmQL4ltYTQJZQa/i0IIe8gCdftOXYItqYRFZYyzo
CwDPzliOxeXVEPSIjp5OnaGYHnMxOCroQM08inqL0bT64cMXHN+E25OY8WfZzwWQ
ap4LCyFhFhWzytpjVVuk3euKIuD0rKoXFIHEb4MJcQSHClnq+SzFigpMGXPsoek6
qWg11i8z9D4ayx9rhfRtlgfAstibFgwA4/MGb8KHO5fQEIKpX9QuriWZcUmAU3/J
610ht4CrPAv59KPMChA7PPcvphxlPTw/vqFII2BbQTyHJzA0fHW3spD362Pdr5fc
mThvLFZLyARXIUhQL9h3YTcWmWCzQuM8sQxjGOS8E+eGCcuaKwCrygdC24TYXses
Ga+gzyqTzo5rIh2I2dZSMmLSXWqSHZsjbXubKcKSsfsWLtReRbkTq3nv4Z7cbzHM
6AaTdfFq3aVtjvMe0rpnzZkX+GRQiUm4B2EzyFz1pcsxXybyrMxY8rPC3khOThZ8
irX8Ic7tqGA2gwf+yjn5UCF6lcZ3+9zKHTeq+cOS9Ijt8HVWxBoRjZmwA0YKicLb
Nctst3EwXS0dp0OZ/hqcPOgehnuj/94Idllwl/HgrPBwlQKpp1eFUQSyRrysZR1P
vgb9EC4sCLf+jIN9aGqPQwMkCWti89+x4UfX5s/K9vwbfLEjTWJm5CU46TPrYHBV
1PUXZlNzaj9bzAz7hRguqZxyKlXxufIRh6nLAyE+PWEOpy6VO2FkBv/W83Z5Y39r
C0QBm8IBhdHZuxTNN14/vxq0rflHucC8rylkrzosJkhBUI/zvIGZKADSV6vd5rZd
W62E0YT1qArxbdyFXGqHq/XOCxnORjjeNBSPIJQ14HYne4JxFBUnKDV7j09PSPW4
fO16kRiZ504G5aXN/sAM/1V6BdEk/kfjDMVJrx9AXdVWnqDurD3ZMiB38EREeRRo
vVIBw2ukk8EEjBcyhRLCDP9Zs1daPm2zoeIQFFvqBpjZQQvcfBrZfxPlZE99Ypxy
hcoWHDEE2LjAhUKSb9c4jSUrNkzYFiGYyJ7EYfJIBScy0BYbKFsI2ihfSjRz0jzi
cDsCDHKZh6IRTwxvXbOXrmZvysnB6SeXkRIe10WjDqAMAIIRvRPwBaw006BSmXVE
xxBi+wkQC2I5IDm53RspIeDRKUq5qrB7fLz25ZlnDqoIFNcf/FxO2fEMvz007N4l
DhOei2Idc+zN1z+bI5Bjg7gGFA79uqvEqnkJ2RMrhRO+ngWCaJDngSu2VYEbwMDx
fodb3yv+2kFBSuecb2H0aNSmn0JoUDyIi5ysXsIRlPciDpmhYj4rcpPCBmM3IRg0
3pPhm9nytLVPVQDhun6D+5uljcoteXt2oXRzI3PL+jawRHlv9R7Pfyw63ucgOhbJ
82ELJZ8D4G9YzzeL0U5TMqh+v67JtvGYo73eMa4Fb5JUxdbIo9cjoBx+rG8KAoCW
fEZKpR1NwvyP1nFBcBxBhw9LKZtMeqFFxRi8g4ZNESV7bt9cb4pzDeu20pWLiO4I
ag6T0EDPBJNp+yyFqoNwEFLJvL+OQTU4/C0sHtYqN1IOGQ6n+2VCsDm/Nrw9odqh
HWV+i3Q+z5m0WFH2JAsbLKzhS1RuV6UpSnsPghLj7FAmXZMV6tc4yJ3f/t2k67+Q
7iqTQWhVLcDIdMkkPfJMytqkGAxh5b7zBsNrStrV5hkIfTKNKu74B9XMHVIJtT5+
5HHL7cpgHG5WYV5Dggiz3a5YZh/VG0L8uqoL5SgxGxqNXYmJiPXbZ9aXX4PnzGZV
a/hKLnoh+Br7y8fyt6ikFe+pjnXcX85/UPdGwcyNkKfsatiPJsp03d1hlUrVvCzT
4hFlgeYS+fgjAlCKHfPq2RELeMgeZ4kBLMVas4BYKUQtPLrohEeXR0cBXstBM0zT
gbqU4dF69i9jqgz9wi2dP48pTtfqUMo4Ii9UhQwmSEiu+PgweS8feryOyNBmiwxN
OC2uSMsmF4/2QGPXsb6Ld1guYmDyngsoHle6Bgnbp+eDyjXVjZiGDmEdgqtDBvIN
I/Rh4svseU8EzvanGbJ/+yll1PWzbvgzdF6+ml9sHhyvZqhtRc4NHPOLf3owK0om
KYJs/MYq6uEc+2O50QfqjGAS9XaPUCJwuWimkLOK/fVMQ6EbEhSTROZ7I1/+QLoM
qYfnvYx0MzpKFWa+Z4CdIYrwlPvHN3uikNH9ixf5w6527+X+cldspk8UKVDjchwb
KNudk5SqEN1ZNnP9AgygeOUcIV7+vfTtkCQhuzSDXgdCEG7c3QUpQrWNRjam7NQl
35LrAa8Ifo6hG70spWbL+HqeXoOjOhhuVfJtTBn6Jc1C3O5dlPSav5KriRsSyzSq
FjN0mHw91DjlhIyknu8Haof58Dn0lMchcnJy5Fy6aFsId/vJoTelNP7SmfMPP5fF
MKrBHs7VZ2M3pTGEBJACh0CM7D1ZS+WmGeFzkR2RV3cJ4HW/8T9xsAU3GD6CUw+j
b1qXYoVGjar4t0WjtJT8D0zvzcIjdDHhRqoa/wh5Ss7XjbBhKc3Z6NzLksLv4/Az
hpYYJtj56ORJoB3IepPPkMnvp/aCdUI2ejE0g03zx1tYgbFnH+B+h71RU70B4PAp
g7+f47FaX7+zV2Ijw/6EPT2LFwE1AnusZgPU6FwBgFmc1jFlCGh3ozAYZg/Cis1H
IrJob6LBu+vQOWytm/BYu7s/H4qPz1rsp6l4fUViU8R3bb3Gcm5yJNh4FAnMLitI
PL2dRFVTHAYWiLsu2x3hYzRbW/5ZIjArJUG32Nb46W015SKiBYgmK/bNgxA/r3fW
LrAd+LtBla/GqbOQE6rsKsQNxZBkJ4zg/ErEVLcTJW+mOtrQ6H4NG9i48eTzrLO6
eOx5gEXFtAgDLPFOSPmvdsoO2j3UrZuqB8ZQAF+GckDnGTVqZEbbv+Z4nkkfRt1E
Ei/nUhBDvrXVbMM81eQEvEXLtpm9/Rpji1RcCFyIEWeLyMvmRGVJ7i0erXWS1sW2
+NbgJz68EgjgHQxFa9/2vqDtNRizqiePA2A+pI5ckYi1iCoQI43PQ8zzF00AGcL6
cmLtW2SnP+QR6VjP3WWBKhEnvpleUE9tYib36O8EqTZhuQeBEMEPvraHuEyj9ZNy
SgPsB73f4t5W21uZ5fSdzFIXow/Q0ZQKjVQV2eUjebqMvG6GMBICS65VT9TGVEfS
YAfzpYXotPVBcC7LPP5ha+tIT89em1mM5mFDV7VPP7ZkyNGZbC/Bv4cIbydjy3K+
jSnnUTxRmo6CzSDHE1D9hbcPTIrHmyHfWNOxfsVY6CGPNIXaXvGD1tiqdl967rEo
9JlC/6+mDK2yPBj3gTELlNX02M4s9tXV9pq2Ass4CDBDHAGxFaYKPl4o1lWeC9wG
hIKCIeLZvWtjnt1p4kd/t3sBfYV6ucfB6KIGpaV9JevyHrj6h1MHAWLaLXKQM59h
KpAf3lgS86IZg7cOqylj7KHJBlvIwF0Y4m+SHJCgv9DJYB1n+FYUdwcL/+nbnnTs
WbdqAncKpEFd1Tm2dfNtPKnOS6dgVObeZz7vVcEUtmVuPyH0GqFCTBRx7npeJs6J
DB2pBytJcT72NgbYfNCkR9+oim15Rlm664zCWz5C/SdcqU1wRCG68v+aVC08Qt2y
Nh4ThMbcokTgR+V15mPQtNEyzs00dybM33j7krP+FTUkdCpCzB7pzSmIBliNdgE8
Fj3MaY3GONK5KOO+OrUGXXwylt91ZpYD4bP8fJUcyOXp9ni+a3Hcsf0Im+fF+Jo7
+G8+2SbpuKWOymJrk1RunX7jRyJWJ7aCBtTwZENYDp87inS2TC7KqB+uKdsRpGpK
wBtQFKAR2+09YBwkGeLiCS2oyF+xWFP3eRKLtxfcKYNL6QSbtd3nPssuibYY6I7z
5EvA4v6T5QHP+g3zepkObrmbhNpwmt5zD52Sw+3T+wDWj53irjMCA+pvPtCLRi25
uKISutZDv2JNm5KswwlZab0d6n7KFuV0/zI73iaZgj0pH1xICnrwZstoKEcRIUD4
bccJ4LdhtU5c93AoEosNTcEQfn6qeq2K+uCM9mPleZL86g77FWc87JaLSy1rN6iS
h+Q3Wz458eBFizR0OLQvf2mKO8mQ/5chtCxDIJY6boPE/RCZPzCbeE1KXbybAang
3cxXGgBreyknDbBuiR2J15vca77gYY5OBei33m009e6r7ga+425w129jUUAU4zcw
Br99RgToWqKS0FV7EPm2fLC3JzNu0uJe5XQTTsZ+jbL7uzAJGiAWmAKuY/Np1dJH
vG00fqogrq7yrnIS3e/98+TaYkkibPFoJbM8vK4odk2oyokV2sqYPzy1mQQKujf8
K0U61jfRWQ+9t5OQOadJnLihkt2Gjv9dbmsn7zSwP95vP6inRNUGagNQDvFgaLOz
uHrB+G6LbMyj4hWT+ncMDsGRNXfwv7L+CxRSsBubInFPo1MXZgucIJj75NUXEVoZ
0gJ9TjAn0/xXJdY6hjt8mLYcAjq9cpGMfGo/SOGByJSLXzztmlMqpHr3E7NRHrG5
7Az9vc2+ioYd8W+8epAXqw3chCB+dOcrGqB1uu8PkNrM9w7s8rgHF41GmJu69fBs
qjERbps90AE6ucK+BAmX9T2By9oJUQC/tGeT/JT9Fd7V7hj+aaW4Ddufer5Nm217
Jz4jjCy5i46rdlJMn+Q4yKGVayzFdd/prGimiiYmWEfcdAD6rdztWafV5ILmbwAr
y/suMSCL+vW44xIVBqg1HEStCtkS997LOv5bboGA+eCjiDmEcYfVjukp18yxMtla
7Tq3dV4maVjcIIWIz55anEaU1L18QvwonkaANHXNetY2EveBqtoIohj0qaOFVHBJ
WCevdwkIqAiA5zMthpoftYR5q3Ox+bkFmGsKGhA9YMihWncqRza2H5wo7N6VWT9v
xLrcfyMJQL4VMhfjSuZ05k0vZKR1MlsPtJfewnk4peEJApzdqqnkTJ57qK77bz+t
QPRtey0FQqECqmG3PH+nZSXm//6CK9i60mmOPTKST8kAxPuuAvjhwmp+8OzloV45
EyBCAeL/tsW8QUBBtEQpOt5nO7O8ml77a0C7eLs7o04RmoYq29+5jxKHeHprJEcw
dgzwqFGV4W7R+LWMOLJt90u7GbjbbrAgjQTmEx5Sqz48mprddYtwjJCW7r4KavWO
vDSF7mKmGzY4aR9+9XgH9eUo662l5QyirqxjuJkGalb4zulVbAIE88vk0xRAdg8+
3zW8EzE/TgoY8NUjpP1PEHSmJ6oqROnhzPF1+h+Wy2ySHxHu0OKBvyhQaeWv+SQ+
UIQ7VvpN5KG98P9y9WHZ/JMF3kVqpQrK2he+tqjT2tvSvwocUn7M4RhxkcIUSZxQ
aGMwH05aatr7rPcCvuToAhTOekPRX6YICyX95n4QFXPev4JzRIKkznhxa7Z06/9a
saStPXEo/FEjpfCPc31QKV+mcbdkI4sgGLcJ5p0f3kZ8zFtwsBHanC64q4XLPQho
bftjsqvy238M8PIqUyJAAMcqVbTzkh52LBGauuCPTOaMjGZIH+nyJVkXkr+Co2sK
9helhOzvAGygOAWEnkDBTaT6uNjbWePwHeuOkqTpzekeIt1JaHAIUyX7RelBUmPy
Pu2ejZoJ+pLMVREcB7E19VJwDcQZp8N2m6NCH4ww5h2utFmC0LHMJYpsUDCDcwPw
Trl1RGmDaaIsLy8z3+5TQotAPWAA5FKi1duN4XuI2i/hrxRdos1eWf4/8DuE35h9
6hkZJWIcGf4jqULkRCpXB2shOve5NZ5YanXw8arhPeiqZ0soOMMO9PwYf7lQSaAM
A7PtHrcjlKC3Z7H2pGqfS+dWSqdAdQtx2susZTAObtLI22L32QCjyyzY6venjakN
DObYDq6zL+ogZRKZB7zo/WS2ZRESaHyt2Unjxkv7S/+jAO1BssBxjjkY/6iliV3Q
yN2AOAujMOR2WJZYfR4CHNLCrnE/ByE5/IOdRUm03F+R0jPkkaEWf5X3pB+T/glz
t5giXoTNrRcCWsM2jBWTwZ09VGC1ErR+awVsGZExZDESu6D8otWgL26GX0Qe6fZQ
KaS4pJ+5cLcQe1B7XGBuxKru3BowsQj/g83IrUnZFq8WSPD+VZDSi7/HCfFNMBcm
Mu9XkdOmQkmvGFGfog309UjC3/nN5nXCGlSNrfEgIR6PEa6UWQVtJYkRD5cBC4QL
QNQRjgw3dKKcqUBtFOTtY/oMDqftqNrMGTJXfqxM7tt9NOaoB84ddWFAFhLtVeNQ
MrxKLgUFsR3GgpjI+Z9ZUyTGAhKOaH8aAVfyuqyt5CN+roP35UaD+5eO9w9+70iq
Xz04DvDj+MvTJdoY2e+/uYq0EsV6Z/phfWRjqHBx/xCVsYkL3bYuJpF/2EJhcnt/
hpB329LsiS10ORg1iMuyauPVHK5xDmYqJ+0vmsa1pDPwkNqgY3b8YT+E58OvPpc9
0R+YELyFiowqFj6CY3jCrBPqqiI0y1JEnwubkdi7uqTqrmSgbTBEOGTB5jyP7ztM
XVPkjqhe7g5IbpOJsS9H7nVyEbFtnmHOtsIkn3PIxajHZt2rBJvsGeZfIORH6+OH
/cSz1G4ZAoN4y2UAW+gmz3hjZkoePiUiioEs7FJGEjRJK4Df0QoXlL7rpfUjTdAv
trmir7HpzQAmxrO0d5D10rQODLD6GBU6+cLZKObX4Q4Us1M8TeGNcWl4LU5ioyiQ
LRoCMdwnlDkBejKvCkBidCqZYYtr3c5/WuHiEuf9JgIBtTzg4AaaCCFvrlG4m4HO
mEpaFaZYmVv1UN0iCpoQsSzjRyd+cE0CcWOKiqMLqXcEekgJhSlHk6OncjtZ+n9K
RFRuMQmEP1Q+wNE8YJBLe+6+j4ddk5WCJ1ktn4492kyFu5sq4LLSfbQb4OMKr2/L
RVPQxWs2BiNKLLndPHwcZ/ksstQYyfQS1YacS2t/AtSDjY1zw62CSPTkblkGKUFc
bytc+3cNedD25IJ5aGaHJb6XKgE1aLrtI7yhFji6CBS59/zuDARR4EergwcXJVcr
FUQPadBt1xUiQf7m0wN8UUz10ByfNVHK0XxGaqhwR2sOHEdoZIzLSNYWxcr5HQJa
jN3XswyzGgHatXea3An7K7575x1YHdP9e2X6JXrY4ej+X8kqDh2FtpAfIPrIdNar
xr2zToJUe4zBIOhDzysUF0aVffTdLfPHkxmnDcrJaVoVpq8j87tdH+jIdOxJBM+z
7LTko1wdc+Ctnm8zXQNWsHejr8nco52iHX6IKtk0mCcRog4W3lImyOF6DiJRHe4N
bkyGUs3MswaxoTULpLiuBnCR13HIohpTkgJ+L97mv1Sh764iSREg6R2zp6WiUNYs
0qabEMh7jacJTuRipIAZiByEIG0Deyq+KceLReLGRSmsK1skl33da/jTIEBOHnP9
eIxUcxBLzfyxnc6/sP/Icb5FPfivwibUxYgoiASWnXqWXVSEmldiBgGoIK3zgLDl
cXgeRB1hvvhG+ZessdBC0L4LWRFUP15S9BENRgcXruiO4Z/GSvjRadCOsdwhlOya
91Gk1oO30O2b1D0LoRc+R3pQqaRplXIiBvqKEtY2YrZwgUNDWsWio8hQGvsKLIcD
lXR555X4dgHXLB8UtV5oSeiH0rg2qkydcW/FA8hdJSTMB4klmr+q4lPF3zIR7SsE
kEq8H+koj0eadHWKPhU3Uu7D3z68B3GAsaTByVbq72bO3Pz0pBN4QjULkK76y041
E5af+xDv/O1RG0evSLu7M44sZvBSu0SrBXGSRi3DTU0i89rBeu2ZGM/pa8ZYZjb/
aMqmNPOH56ooVegcvxxiSqTsmEdObyAD8IYyUi46V1mPJwBa58V9NITcNAuYavdD
JsRmQbXbbKrQgA+nBJPXcliBl4JGvFqJregEUcrd6I96kZSQ5wSPZT+va/ZBMsKV
o+2EL63vKvelMZQ9L92MoY7idN3R3GD3K+22XyUuH51OnlnVhiQLljobOXDCGR63
8UPHz1MWXnJpfXPYbPoSCdBmZPWRsTjz6FHiZmNCLQzfZESJTzpXXLzBiv6rQ5AI
4PXkt5Yhk5d/eNhciejiWeoJFWXU/df+1cRpRy69uVBqH2+gRED64DfVe00frov1
Eo+tIuo34WHJSOwQSCDV89cDbVaD5M+cySlDjHZ9HM4OYHbTtvwMWaOIn1T5fYC+
ZsGmWxr9lXrY50bPn4UD/SbqV6J/ovVKILLEFlH8b7ogoODHoTX3w0Hwko2Z+0Yp
Nv3lSKWJb76xts9nkg4PVFGkF9d5Pnclvj067cXts8wt4rAsTuz0ZBKWwEtpvYF0
JoFDEHENsq8bUVm5fAV8OePUsT/ag+NoKYZKSjSugQoZkVgzc2PcdtCiXwta0+ck
+htW07b4Qp65Qcgt9aXUpX7RxChwtBfg7PbnNxqLiUsIMOo1nkhPHusKXdjmEEpC
rjB7gyJ3vYY2AIRSbHzSeBZMY6rcKmh59NBUfV8a6ZnVbQuDcqqTDiQ6dO4wjDpR
p/zvPjYvM81mijB094teS4QcmCABi2unHDY06jTWzhXQpMK8y5nZff49AO9VK0OM
eNxn/I5aGulc4FnzUz218Hb9MVKJw98KEB+Sx8aDy1o/H7Ja+nldTkSHMV94TMmI
lx3pTCnVrGXqzFVIu/wvZRRPguw9Sxk7fyCJQcTUUvMRDHU6i1P4GlxW+Oe3YmWa
uH/z1FD/2ZerkNoE/dL0fcT74m/V5HS3LSmHSRPD6aUQRhlJxKqxlmv4kqjI/z3W
d3GHZvLI/q/KUeS1DHYuFAdyymiFKYoayMkmpBsGzW6pukBLJ3UyIoqngyDo1Ixq
RCDs41DM4P8Lqj/b2zwQJnMx3pZ/vXQwbSDjdsnAGzSKkYKcFHreLd8yxCnvgIrD
A51wJqkAHiHcyLy89/LDreuWgiml2tMMAD4c1VDHHtbTPgeF03+RSke/ojj81ujX
8WoXEYAkSOgv2CQnT+JdLktaoAkix0/437YtoW5hyZI6jvVhs8RvnXDMxbgrQir1
aPX2mjSP+sin0ibeGY9i6zim5y9PchYPgawHJLk+Wo2eLMhYpJXX5HYljsDJLrTZ
O7srOqgyV8sMNs5/Al57BVi3EVbcYuy0sljBz5MqaesA432dPzloresOhlfN37Wx
K4eZOtDmMDUBrp25/WKFqifkRv/8xdHLchj0gV8JnV05U6nqng4du4sOUxdabyrQ
yD1zhxuw0saN8inqN/G+L70mlm7FzHJa9G4UldJAUUrnKJSg8eBNDpzC6hc2GIGJ
NvJXvUZw7/PBpkfBKnoTSRIX2jVuwdL/tHW09Ci/v5Bw/wgV1Dp497JY/XZwyugu
8WJ/O/vGZ4ZeFSqjEVy1EPwwWwfK7ak18KIVwsTIhAaK8Jcu/l6+jfiIM6ygdf8g
KtrICv5bzz0v2cd1mVl8qCoSPwXzzQDiRAlhGQ5vWSPr6OzLpZhIPjYfYM57QtDl
LPRSKCqH5uswDFN9lsMXXD6OQWFlERImUXzU33uWpcesm2/PhU9yNqb2yoR9r/Hk
GY2oC9qw5KtOzepBNDzQoXWy3ND6HJWYhlqi+E83XEUrBaRcHRSE3qtzY8gigTHX
NoSVkxlQp9JdneBCLWWMnm60BoZox9Pra/0fb7b6GkN7jOYHfHgvwGCbpVHd2qaY
krw5gCbhCE6Q8gyF9SK/H7aRncl5Hhf+NNnXOnlyw3kkxbN80pTyekXJqzsao+2c
kdOrBNXQ5uh9wYEzmu1DguhYD4P5L7PyJTHDXMLo7ox8GIpVlwEErJIvy4A2EIoa
8PJEKcP/7QRZx82nZrZzUow3JibL0bxdq5juQ2qqsWnHQPqOfy/HxMBrl9Q7EWym
T2/EGJEzHCSC2txc4s79V6iAAgKouBL0CvMiN1pQENLphi8qaCVsSaHuocLxhWXn
ff28eWdqX4q1aEAC/KWh7heG+pv4y6tvVSTPaxzn2xGiqPa2G3YXY8ricY3PMkXj
3nQ5Mjx25l3CGdairA2nHZCszILt6GQpTazWTtPRlCJPNCnVJJq/LfF6O0qSCvrS
Q7CScQhlGimSwNNAdI5dPXqe89S6+kytC/oVoFZoiHzytCV/we4DF1BWP59ILhAQ
rWTicEVBmo9qNH8LSrkXv6aZeAEyMUaUv6sxNcDMAyBHz3Pb+6j98BOykuiBAWyc
oQQaFC+aWbelWRaKciHp/t7bQub8MiUhljIwbW9SnF4PB2V0Vy+qjuJsh829yJZV
W/7lgB8LHfl3+9Deg0YDVe+YJdxR7CtYsbRgI2PJykGN5ip7lVYFTxcOvawdjKs/
ny3LGgZf9QMRdkl6gX0M9P2WTFtF9uD9iC4QNes7N9uGoTIQLw58Z0Nz5R7oLr3q
Kiw0yeJeX7kIOAukUoifFtF4VeBXsjMunabYH2odWi+WUY01ky0KmMIypO+Uo6AC
zv3lp/lmJZAkoNgQaT0lEIiHU6AEcJRV44YDaT82u4LQoXKdR2QvrINRYFB+W6y+
hfcDKRzN35q/QY/n3ChBida+e6ggHyalbY55luIMOocIC8aUAYk85Xlieqq67gZw
T0N7B6bo944lJqwlUk2oJsxmaUyxqRi8N+lrV4uXK9wRQZtFfSJEw9zmrT0gdljr
llOdZ4oh33EKFTcH1j/OI2lfyjfzwsjtbxumZZZdGrkSyEl3O6imWCIX3jZ4y5oK
O48OKYGYFjmPr8WW1OZe45rZEmDBJAEqHzdqZY8RIGRkfQaaJBtQl9hrQ0Q0kdFv
M1rpYBDTWJqJzggYjLR99AXDcXsgD9awStKxYAmaITejFHiVGDCZsbIHRx4TJaGl
gXdPS8TAXI7Kldm4kQee+y9j+fBGVjVrDz3fengkGIcSwrddjN41VP0h/ID5Jq0R
8npgNt2xbMvXUn3KNMmiDj2TXOavsw4SlGzvsOHK/CiiGsSSSU6AInsGLw/uHi3f
ZqTfehkLg6ehWz4pj6y15tw2vqCSJt71NlEcPpOUPUtgHqWgBvOTO2n/ZlH5YMSH
Ao0GwMtCvbIZkC1Cx2dLfF0/Fg7ATCNGxZU7/dw+Wm5BJgrX+kNOkWhSvKNQ6B8L
colvJiflYEBKQSyz7QUvPX2IDhVsJ25ahwwdInV0t6OAtHOj8lsGqHfjX1+3hp8j
mGNOAskVBDhz2umMnk7R2U9PY48mN0aBRwIrX2qVQWAM0eQPDLEk/lwbNYm4di8S
CFGMhVZMVZCwnz1fET/Lbc0vOQ+9/BrwNz3PhjDl/W4V3kk26WvTm6Fk1WzjglUr
pAyQl0NT9yYlGGVU3dHjbXiz8hjH8LDYRCaneDt1X1PmgmSCBcUHKpzLk4TIOlkf
GDSJY2dsspGSLbRJSCCYv7eczNX1GDkzwcSjRmwsPX+4afn6MYsb+KlvakSWbKaC
3ttrrQ7LAHXXPQJtRVfwMO1NcyGiCLSJQujxI8n5PSAIVkw5XLzUjnElw/iur/fy
fEY1WqjXsrQz+iWyFTYf2oCAEw+An+GRftAK4P4IhwP9pi9c1u120eiG7eqfc8um
8Ew/a5j6+LQL4KQ2drTjFVNJM+913DFz9dHJ9kSqkVrxOUJYdoQ7yi5tFwFNSJD9
sCMOWyOB3SOeB3Kdoh0eDwWSEpYYiw/RehTtxEEJCMzPxWkZ1kHY8L/9nnmR2Alc
8xqIS5+F6B1ueSmylQFjrnVASIIyTScv8oegn53vIUiVoHmrf98ABtw3Wz8sGmXq
N+XBfx1udXgVUsY5Xn24L0VynHFPANCtJ6q82vxuXZJcDpV3TS0fWBteQP7Pr2z+
XV0gOamspVEGx55WCJuS2rYzVSOEmsKLS4jx7xz7ZVI6EmTlhtoGM+6c+bPfy8EP
dkbKDwCem3kP+LnQuGiS2KjxjuXHrNkccsfq9582kmyJOfzJ2x+5wosn+6ju79Nc
Pfjf/jG56uRBBgBm0BbApWH3jAb0VRwRViEAoNpzjwZ373OBWgAK50wbBdSZ3Joo
68ImcVNEIstEZ/3hJTDHAZ/G6O+HMBAScHTXLb8XxmxwQvenOV+CB0HvsjlW3cxK
R+1osb7XVXfbB2rcAdhRMMv49x+njZvuJinFF0cisr3WYANGRI5tGz8dmAO1t7Nu
DWP+Ra8A2JEJI6ByaFT/zcRofryMKPat+7BJQdGTUyHH4AYfJ1MUo3z8rpvBNRnM
CqjIlsQne+QwBynFGTWQDxk6Ul5TCu843+i1z7eUMtSF8HIsAa5Z2tK3vxHeADmd
s2ZWxu4ngHALcO8QBd+xH5VyUilnV9w1OFimAX80Cs2YtHkfn0uAOKcyxtZKBrAJ
VgzBH2qGiqCsnW3SsFE6PtGIGba3Xns+H5MWfahrB08X9/B8+PgT97r9RATxYL6+
YoF7xpG973AsUBTItC8QfH2lkYh/t6o71nThXoeppVRT2W3MEv9d+SidNzDREa8e
HGj/xMXMBZrRW4RjWPnrK0Y+7bGmB/4Op/BD+Th/mcFadj69d2qkMXZWTHW+e2NU
7/dgTq3xcTsfK1hgitp84vB1p3D5hH+ecpRsdffAwKyzbFOOVn3bjPJHy96ZTGfH
X2MLybJ3xQHbRuwhbv9SFsZNpgAQbLzPqXA2DloAPwu6sP7qAABlTYB/n62MCgj1
x/Sv5SmdpKUbbA+ftjsQ5DBEL0FmOBsBgI/XIocv2Ug2Qv14c2RJSZ7OpnfkR3ca
/Sg0ubn3mzaH0X3yFPMX+7om5mRRRrnp0oKjCeH/REZjyvfbsa/gxLcAVgOPZRNo
7LWMSWmie8bScidUMPWcTluaNgKC00hsTHS7KZML4LIP/OPhEZSkfHH1M65M5o0D
HlykU0ws9tbKzt0thDLpqJa12m+ubZS6HWdNJpFABkBNh8rvi1bTmBMZe0AUzPBN
Tjq8lGat/BhNE2hHS5fAzcV+O4KMQggn4D1rgcGeiIVk3JpYQkHX0cWeN/15InSy
1KW9vC1CrVLwRkrOBN7IlJEnvTmBgc5+wiZ1CCm04NkmW9U7qstrTSZGAy2xZ4yS
mkl1QMeh7K08k8Xu9JQljo/qciJk3DdjnQckeIwvmbfuHmvNBzbp2VYDCgtPEKVr
ev73lB/4bTp3J4nSlk8DrVrtUWBNO00bjaBI1UX+0BuKFF3zKgSJVgvg3q9a0Yjp
Ig0qAX/lmJYm631TjjZ/iLHxV9f2SEedQFDejHVXOC+0K6s14qnRzQWZ6UFsPSIn
aunyND0G5VGgG1EZ1YeK+7g/GJ5nMMKHKNlmcrd97iCOPp7EJ4HxSXNcNbVbZ/Z8
VBCK6cO04GGbfDR9Evb8SrSlUX6GgbaLUBcLKt+jKrYY37qjTnI2sjxno2w4TYkL
rZH9w5BYPVQXI6WFPcKtnEc4ag+oOGb0VK2nn2REXz+gEhcnUINs0kQPc9boSymy
9aLr6xdbsNTQoctpZEoJUFvvqHWJpj+HGviMZ6ETrC0gKc8UGyaF6thA3ytecFpv
4c/WjvisYqVmlE4EgpfnP+tuLlKECg5kc/zJQg8dScvSH/oCKQP0w1qPVkd7TJL5
elHzGUGCks/j9yudkGIERdZyVHU8mkKYIdy+jIaXIqqCMuMorxD9c+jOE7fNxX08
SnEc3SXdGRIeKvOHfaiWk8CIAPyj/PnNuhsAZMTJxfgItFJFQuCwYgmQlZyetwe6
lvfwpKxmnM9TkDrMmY3E4p/PKPkrZ98OqrsThnZQwjv0z4aZIG2SBlbwTDrXLDeP
4pDqYjWKFvyn8C1qKXadb6qFbkNhj1E6dMwShYqGxHyXTOV2C4KO8+cOckvvL7n2
2MdqI9xhyuZWNKiS1JsMHntVaT2OlwTmDMgecNjo+KPbS9ehklhP85QpREw0tgW/
Lw6c3bsMZn0hCT+MY5TFqqIMILhmopgR9URtXmCEXvPAlOwRaqRqlkfrzzn2KdM+
L78JOFRwDyX7vk0B7ZE5UQ8sB3AaHhJj6inseMABAhBHCpl/AcG56MAV+unpgfYq
9cD3jvmmyvTMne9xvReYPohm5T5ala/Ndig9TVVPBtPWqbG9SbN2TXJIbFfNJtqx
0hyChKi6Eo0wVUvdILHGEqFQ+ezlTiR2M8CApYGeGv9VFcJeYU+4wl3/yqRso5eN
vFue5i/kg06wAMPQv0QydCa6fnYq9fWTIa+bIhfA34u3Ni89zkZrA5tcSq5q5b24
c5UX4sEhnBXv5wg+E7U26hG7Sy29aX4VLhxRQaPtQtUAMNBObS2TbfYazIvq+9OZ
M3YhEN7mAu5zBFjCrUIYuil9ConLG9PSiOKiRMbZ8SSHy3N3PEKplznO72XxbO8h
pVA6Wv4jsIqG6XV0OuU5r1tB0/xVJqy3D77MRw20Cr/T+g7qeYkibwRSy0qxhTSF
ou6/6y7HHZyfK3hnEfFNQ5s9xVRM/hNoLbzPUd7iXnMy8muzON+Z+zkzfTL8r51c
8oSi4yIJHeka6sMjyr8ccvKw68xwGkGKkqsZZSsdNdZJ/0xisMlUTwk0Qx0KIEFB
9rJSCibby4v3tmVvOtpBpObc+DrUkOA//l1/UDQWtJNDXmhhOkMCRBenyeBhHSni
Dy6v9OR3R4Na4DLwfpTa5oidppCQHX36nkfXhQg1aCieN6U67x0aKgh3m+9FWiZq
vzUVIHgDBCyG/J7ZPjpz2pPNhmnUs8yVqYWlz3dcHRZbYL74wobIE4WxKrRQQyjd
IFohd65tLNwNmPEXBhJq9QxYc0LjzZ1viJkoMg/5dnChWR8BFcz8Mcizb+Clh9uV
m3FDVR7NAIpTDKtCMSA2SnK/uExbMNJWzIZDu5p/0+5mQwR6hRkywz9cJqoUrlhg
XvLGXDTP4mdiSfRe3RGyRxAfRHbmdWDVp31+7B8nW72Mlb72djJeL1fowBU/7XMX
o3liaxoDMjiFeKbcn+7w4FK3RKwEvRK8bMSdW4SH4wLSrfL/5cl0HwADkURjNHXU
MP5SXJFwPy+mnwIXvubBbDs8m0MpOHhC6UlgjpV65zys5oQL3EjaT/TmQGdWeI78
STCx5MIhp7i9x7il8Kh+eiHoBMi8iW3ktCgWdSo01MOBzBSYlRxuaA6lr5jmheyk
D0aIK0e7aKLLaD0hSjfE8cYfE1OgWig+Zu0WKgsDjhNEdSBMEqsPKNfeFAyd+dy8
bE2mu9+LaHU+BRieKv+VvMHCXJHo/z1vhgw6eS+p4cjXsoMus69FwEkcQkagual0
4/jdVOOYdW1zAmcQ5WkC+LJdF+DEuIteV0W3+DpVYvoVT39Uq1Qr6IyBQysccWD1
6IXhkhctXLO00EjpL2J5+ub37Y4MbcNmKncN+iEh6rjBRZPoiB3dBAHQS1pIu+op
Ak5B7yb4BiMywDSdoki5wt5IndkhBMThS3OOupRNAan/mxPz/phQla+79ekNRmN8
1tkG/x199KvrKp3rVsDDENCqEI+IVkrXnINP/qjNIPXEAjAYAd+Ak6t/7BEc8wTu
yV0DZCmqbQ9IvCL4fK4h7sZO9SK41xmN82LCItZ0hXgC4YLMm+0XLRVifHKpSTI2
WhPrjYBkYaiwHPcWCfwfjnRkiLn5RjfueUWcSK5FMS9jJY82hfQnko4BeZDaKYzi
P8sxjuoSaKKlwRapDfxlTAng7HDaa3Z8oX6LiUsHNojGWIx17vkOjgYOILBU4mfq
o4hofSh+gtMEM7eizLWTXx4seD4bAJd6z8hACbOCI+2qbQ6+/9e6frkCgYA7f0Ic
UYP0okh1FvNCF3XkfoYMEjIUv5l/I19OISKU8ReLauX8TSTGa7YBuq0b1tqtt7Ll
q6qn04fU9h5vuqI156o4nb0K4e0WX+N8M0wHBLJpC49ZIKqWKFz4+Ep30BORDkIw
B0ONjZiFUn8rgMPSbZgxFR3SmN420TMrGwh9cnfzQm3NacSVIURXyQGkceDSQKSt
4OvplqZOlFesh7mzzp4yXo7Iw9QuoyJPY2nbRc63avgIRqk/8VbpCXGsvmLdof+F
rQ0TQXckMB8KQntxVSqZAX5dLpIW4pv7NXRj84/DXny7YrmKqF90PoINZpilyscg
YJrlcWOktAo3NesT3EdkgQPHngwH6pIHVwN4Vxe7BWyO0KkSDhbSWQmIBVRa7lyC
MAfM0kwdaqQ3Y9pNjmu9P9qSXU9DIBpsOwORZKw5C8f7UPW+A/3BLbtZgIkKkVGB
Eg7fv36pzBnpK7qjyvfX7YdUuX81ryXAoWoOKG+hJYv+iqN2iF8//yT3eaGjH1Dq
tpuFnpNwgk7i2OaF1z+NTT0V+jdjwvzyksvK1eYwrSrzvGaAHl5lhEyj5L0NvG5z
B26NMOm3GzFNGdsv1ULQ2ENWu04iQ2aG3TTdbPuLY5ApVRZGmrXcboQGW6tp2KxC
JohGXPh5cL3lvieVAt/tFN9DcRPJgw4EUK3e2cxrJ+jkl1MPVmkAo8gTou3CSad+
gp5bO4OfyaxNxtvNXRl8ZC5UwYoC7c+ziLPHZ2hz4NZUude/5sydrporJ3yGxfdo
foVYjNI/s7ze3OnczXb2H1XC2CL/YO/1xibhbzUsVEEtt0frsFWL4e2N6ijJM1ow
KMZ9tflhc2kgSxZLygyCVDBPKmUoADqfaKaynZtq2eEV/1gtueTZVwK9vG35UWQr
fip+MlLF8ADdTYqn3QDuVYcqBia5H6IWf0BWap83NAExA7ShZaKUAd39ECcM0kfo
E3d9TBQfogVyyvz9y1cMMuuePxHIisMzUYyHJ6iu0yR3IP+fTdCnsqCCJPXzCFdK
aCrhubToQBTPjzd9AkCmWjTyQdokIsOTsibmTLoQtgj3Dw/XXLXbcsJiG+xuXCrj
LauPomedT6fXy87Kz4GHI0FfPNxiuT6kCgLUJS8zAvZXfP/4wY0LpDNWb4MfPP4v
M0j4OuGvcsRptMRapdfkAjzwz3WdihfPLw8kBTfTqYUK/WEdoOmW1hSAmd7lrjFK
95MsOZShYmtYltZgVyL8it2PKKcK0ldH8tH80uiunytgJabHY55HunwOPvzBguN/
NJUnyFxzI9nHEvdn+SRN4b8hz8WC7xkpZslh8/si9qDlTIE41tShWM8cqgdQ3dmB
9rqIAq2GZsSWSuMXBQ9g3nuzK6VExPwO7OsF3ddFbOqlJ2/IRsS5+iX/5bNNJNZr
7j0tsMOwC2LOWLjy45eLW2daM06ec5gSXfSQ5nx6UMyfvvXSBss0Q+QeiYUE3LaW
MLF3j21Fne/j9LIEkxTDlF9p9zFrpxFyMhcQkTpBobMXw+2krjlWPpQBt/Au2U7b
TwvSTaiAmR0mZjRry3owO1CeC+sAUY7UItCwI/X8e+HqrtyQZGt/8uYwI7Faq3Wo
sMUEHPJDf/0XZAaOzXOwj7JQf725ltrvpyCKp3JASSeEGilEYmwExpW73SyWbUCV
wM14oc2qFV+xjsBR1IfqlMMbxM83mfhDoZhUimEIoJFzL/RcFGk9+IjY5UqAQQ4H
1kGhBxA1xFqbwTD2q9gpq0YWFNJqiRT/ja6Lr14HCtZ0PYBnvSRGgh+RYuL/6Rlp
H9lHQmbL8VxYa0/WxXVYKAppJXd+FXfDz2FnTjD9jiga3aF4MUFvK7NrAceWtH/t
n5sA72ywcBhMzx14p7jsZBFMqd08+VzBJjH0SkSLTF3yTE3pfzngvhcsJg5LfxS5
7VDK7Fk52npR/LCy2eA+oiP+/tyXtlsLuEQ6Rf2U6u9pLuoHb/UtIxBErlQ+oNat
mrnQzHvR16RVyfNqpYsrl44zilE+OVUvsntmcYAItTkENFmhezsdfR2cV/qPYddO
dR2kMJseCkGa7BG28Vvvn5f3tGsMutpuYYlo7ZNOusO7a2DIz58Ej3bZxWALdO2c
5AJE+2k2iQ/TbJKqmlxtIIbt89hlEReq+vux5LD83/CWsOlmn3D4/xRBhizU0zty
38RCjK7nIiFSl2cBIcx98/7HUrjkt8ycOry1UuCWEWHmGk7LtHXWg37+DI7Kv0XB
crD8mDVbkMQIyJNRVfgozlCG5enbz3/Wa3LnrdvWe+K2QqyrFUZOPMxaXQbgBZjp
q/qqsYS6AU/p/yGBGJnO7kdguDLKEsNsV6Wv0543FQmqk02nMnAuEloSZQTPm/PF
G/Xb/sfDYO2laIu9l9h2zEwhEEPUda8xc6lVRAWbUdNEueZkQxljDfBl4aq/iwA1
0Ak1kHjQNKyc5d7DlgcolwrGNyVGX+kr+SVXWtraCqjFDlLgyRVig9eafMYbxbpH
H3BSBFwCsaD7FDvjTbpJvpPmDZJgoCmyVjE5/DwOZ1rdoAYceQxKJByvZMfMMocY
NR2ai15WoCOz2fFvXJgUw3dFMOYVBc8Kb8Epx53TmNwMvdSKhtGvyiW4/UPdTKkM
yGYIV0ZR6JTIUa9NwapSBrGlKom9saMfkEOAKiH8cSD64no9oRYD7+x1AdTAvdI9
EGkJnYUvbiRFMbeeveeiV3pzVl2BpvQ93eC1WqkoaM1hfxmHiEvfDQeivaLpTYBa
Fs8d7nZqccMF1Ex1wcViltD8nFScNgkmmyZ7q92Of3TIfB6awC+yxuPMVTepu6D3
g+EbuYF3L/MGUadwZUqAnRWwjgbnl2eYhKg/oQwxaUCpBChav5UE1K55QOPXXEcN
HIUU0hLR60/WNfSLxMcTdTIRNJWsxvjgaTQKkZZu0b5nYkJF+5fq0KxUHpIZPYwW
hnjCGe+2bLUXyUmdmzyK/lopDpYfORl/xifUbOIG8sWUoLThnguRQ5+Cusszme+F
kE1lRMq5LrQV4FCX8t3XzMn+KHr81AHL2hX7vmmrcNJs2bwCKj+UyfoxlIYM4s2B
cQCEi5T4/fyN0UcR61c5Rocxdh+7+GQQ5pc5aDLRJWBwoAQWKVEEPy/EExqN9cKI
5BXK3RhhOG8uxVNlQtCO/rC5jegHIDtDNscm3S7Od8F6ksMU4qCemFTgX5kxxKKW
fKgt3KTG/vz4kNp/Je26Nwujc6AOfzf+UULm3j4ITJJ/cXZiO3xnGqNNFtHVfIZf
ss93yNKzhMCxHJyz8i42aaB0jitvg+Jiox5v7CRnEVe8zzoS0iGhJKZu5NLh58XA
DaJLXn2uPrqavPLx1RJMRMW1dMAGsQbsBKNHCGdWGJb8VCuXk8faSZvHFYSTrad+
VMbOphXnFH5kKvz3EE5fi3L8hTSJNRnDUt5gYQK7yBZiZy8tGSJDuJoTRvfxuVyH
GgScAlGidwOnFAFmHrrGKsQwrfr4JRak0kxrbPqu1IZV8Qp12Eyjp+Eb6AlBJmTo
Cyj0usYlD3cWUNZ9ALRi0DmCifmlmZgBvSyUPT+aF+nCmKTojtN1CJEiZRt23pOA
Ajydvm2hTSp5LHQbeYsm/2LXgPiFFZsuVqVKkye7iyiTzAIElUPyu1PwAyjrQqRd
d4qGVd7u0KkULzf4t/aHJobEEinI5v08eTf0B9buv7yldalH0HxL1MXtWjAeNYvG
CtPZwPrY6dttoACxQUzlZpAmTJmw2nHFrf7p5whXjFLXOxcALNOVRZtu1hpGhy9U
ECCRnuXtRiyx6f0r1bBSnZY8zH0rUm51rCONQXEkvUklrIRT0IzKh/EriIqtIRrb
7Dc8LBgvGtpDp6KxH6tzAbmqmnWBQyxwEV4lNhwHKpZWA/JfK4UsCtpj6sjfW4Zb
//2EK7Guc8kkfHqnawgOmAspRCoCJ2HVuqvSMu0k/cR+N2HrxatXeLnr1/ilU4Yu
bCFQRd2lf6EOf0KZJmGhZL5O8TKj2wy+1NZVGgdQSAjxvaJhO5hiorAVMuaH5qq0
VZ03VfcC4KonF7AyGU59BghtnNFzpK6pTZXXBp/btmZ1C7a/SjqhxhHEkGqTrFTm
vy6qMhGTetTq+qhT/Jvy83tV9fLT3VSv00lLLF6IWUJre5zbyyr6n8aC0iCXfxGy
gUqRmUWFSyzEO2p35NT2Km5AMZisuCyqOwPbnDchRtULbwaYU0YIyL2lUm62hC1L
W0dcbbBmL8d4YTQz+JVysQlB8YJnknz9kCyiwdoWluxz5EUDNNZB+DymVPWd1s9c
vrIIdTHPoOkvcm6/1MUSVgunIdU+KFNl9faN+IVNrw1kC+uDTA+9urUr7rF8HJDW
Xwg+pCXFLcZdSp1mUyKIarJzJ0L8YRoBscrOQ/wY6Da8hwjHqW9aJvQaOB9vsW4k
uLugFn8m+lvkDqnG99XMK67fA9JRgz6MBrnn6CWbKX84pLCpOnG4ykJMRZEuW75h
eqnvZoM271MsD0unj4Hge+R4iZscnD1bpZh8FGixsU39xNP05Vp5rIGiCQFqRQxL
Bw2Y1aKslDrigb9gWZLESsHDTPVKrp05DvaZay/zjIfO/NgVeK4nTZoabw8X45Yt
knNIKKlNRp/STCXrmUYsQ6dC1r5ApuGGhfrFKE5BDI5XmPynEy27Sz8cXx0L6MxJ
B4tc+pRrnB1XYzAJ+CEpHOC1Fobj4JLCy5jbfEAW6rv0tPC49L+w5mFqbgcPNHdi
2knf3F23y4BbzIGMZ5FfJWa8OnBceLjrxWA37kQEUahrNfvC1VNjdOYUm2YkIQm/
RYvlyRpjuytYKwhg+LZdozMFjp7S1ApVid8l3Hkoukk6pu2G2mVarBcJoWSuZswq
VG8/IH6U4Yj9SNEiaPMRYkYmDpIUTe+v0oj7JuwGlILbcpyfXNK8p0R87Qkh8GXH
gKaaxpaimbPBwnLaiwN2EPMdyMWQoN7aWIXONSVFAR2+Gsqp9w2Bjnvn39iuuRMB
AAM0qnGw6Ag74C8pW0ZJm+lP+xoq9tYN/YjZlWEOwQFCa19Ay0o8Zqmssv1ORkCd
Ai1JXr61VvDwzdOTrFg4goR1knEtVU0dzOyJvrgLNbCal504NdE4TreeLm9Q5Moj
Y3IUNELMVJOSITStznjo2qrXQpyGhUwrrpC6GuYLLJGOxTeaQNFVDh0NTsD1e7jX
uCmCiHyNgaiGs4E1gAiBxukEU/D14LPKJCpczfuspLSvfPJVvD0WO9uAOwbjRDo8
ELMdt+xPQYKv0oy98qniMRSmOFa+LE56W9svdjDY2daGD7Duu/bNZrw0DnU3z/Ut
Lt5z49l9nR39sMAydOlkzo9IHhew+67n0ZT/98fnzVfxzfDjg8meRhO/XZ1xbjIU
EkqTQJYYDt64agUyAKMx0k+LiPaUrvWFCIIKJP9FVFZ6exjymD9xcH13OIzbyKfI
xvpkX+SeyTeSW4OBKEvUPM85H6ieKdBs3MkIjjAE1HKYALbWZswv+mBook209JwG
i0ZJvGIIPVmRGOMFdSzTsYF2F4iEOjXAek7zqKh71BDKoE6A2fNsWtUSZiN3oExN
7MsWZAUGOKj/qd9PyexPSPEnrxXASLzR8jeStWasgIvP30s9zFTjExVwobvCIEhK
0k+ZwK4VtgUsZSqRCRP0r1z93zWbxbRyrt/HSRjz4BNbVSKek/FUcjGsprgjM3iK
qmtsuQIuwaftQ52Rpk8+uCp4l2DLXsxRB1hpWhMCrBSzeNhA7OxJC765dQ0aDV+B
zBDWEsEF5emODtI9fSUeOcKHucmo1GyL4YRjb8Uc5ggyQXBUJNqJjqyTPtD3/RLY
0n4rbU77vuXAO7jglfN079WbSeC9NSvW2Sc2WGH0zod5XMoZ8hnW4VzpbNoTFH8B
ld4A0x+IsATCSGRZmideAMb7Nq5/5V1ZbXQD28J+hXfQTjuzvuvCS0C9gtsCMWFc
VEiNO1J+ajOAxwTEFAXgUilxfmFPxI0Vt8br2QOV0lsW5F223iIcuKK5TmUbAANG
OB5fD2rNd+CO0zHm3AMoWJDsgYSC9vsM6x7IGv474oYj5RIxVGiFoNM0XMBrDmjW
3zsubrbVDD4S3d6yVDBy755dtS1PubK0sKjYLzCfoFmt4weZKnSO3v/92rCTSR68
a2jSU81abtTFEN55E3c9gcXLJ8+2EJdvKYx9/0zRtS7EjD7own1T9JZjDAHRXaI2
g4970pSPHrLWX3W90FGuIPEdvJF1IAJVu+lamubA368+gtGK64jFxAED9YOjF46j
hlKoOb6cmgbeBz9y5rJT3G5QjVgrm6zM8lAAlJJf/sgv5zSU9pYxWjfCDxJUcwRs
BlgxyrEwQvNQh+KfKAmKWjJj/mJEiXlDBCnSicYF5oup5/NrymrSjMVn0+Uh3bEF
eEimkllcK9bNKk0V0nIb6WhIgNvTjqQkAfkEeZhNoKGeTMcA5Gq1sXhUV7wJATcK
RsEu0iVezSBUWGvo/rN3r0gKFWSdPue3oWQZq++cn6cEXhExhaJ8KbqT0FHs4LGH
4LIffcPjThh2Iuxz1xR/V5JrqxiM1JEdlwxWYCHVLr/QQUePg9E4eHBZw736LPxu
wkgM4tJmXL2vE0rpsjkER8SAc0ggQMNPnKBnNlfm0HzaYMDn/zPIXqtUlrXUwc+D
DcfEJwmZg+9OozsQ7IuKzICzpcjYxyoEUKp1IJ92CgxVetSIgkfWZkmT/y+x94Dy
7SICFaYfojkybyFikH7F0Xf3slFSdOm14Ul6nDAhOnCoibzFS8YOWePoqifMWzqD
HJ7OTbz46qBDy72zwMBedkNTdaTwmskrQgnSx+bhAiFEkOu5h3zFGlrPVwvz+g0a
BbQtPJ38zV9AiAc6KpQbvDZJPFMY8c3BmDhxnY8c281D4A7nsHAfLq7uNu/X0NPo
qU35gEzMO5F+DM7FXTSD/QgzcBktdDOkVDbfUqmrE2fsDJUrPD6BoGtGfkCKM9vn
vLKKqDdtmmjbJbA6ePfCWYKv+WBpE6AXt/But3TQt0unt2bNhK+ogUQAbiM2+CeY
BQRXClsERaDtnBq4FAbGpZ6CNuvFw3gWzibWfPlh2Z7csCCH583HIcKk2LyoZdi2
iz3dgq/rcOJfZ4mambvHoM5QQZn5H2Psz247s9CoqrJZu7CejgpYr1OL9+yBcw3W
7nrqCGSI6XgrdgTailIGt1vfe9NlkRhtHNM+vJn6X8g84xbh4xNnUws9cb0yXRGc
4kVoaXpqp1/6H1HJyK6QQkGEZbFtLqE+jHCusSpnE3irIjEBFBNTLI+9VL8E/WyE
msigXgvYD2WPhstdkSnOEXg3vpwSXhMG0BiBnQfInLb4QPg5tELz/DxEeMpgZieA
1qdRYlElS/KXle625J9QeN0hfwBK9diM2Tm22xYB+1nMLXOkTf+j+iSTcM0UEyTk
YaGIHZm+sQIEVbdicIzrZRTqHP0414lmbjQqZ/JutCwTdoYiBLzOLy/jMbasmr3F
e0WxrXrWq4nfPc/wmzi6quUuUjHC0anmTg8YFzQvjDEmEWtbls7GUH3vGSw+7Opp
EXd8n61mJPuMdu1JFogCmk4YnsLa9dJEYbRWzginCARX1WESI6pYW6IZNISvnPUo
NZYx0CvESEKINL+QEgC4sREhmnD6Rryy4+/+IcQk3cxrUagjzr5hudq1+HI6cvD9
4c3t5w0/ESbCJZSv57BaEVDhuT1lMEOpxA3MFyVcHmheImS3PwiGW938iP0rR9Lg
LIc938+gZhfAQ8W5nLHsr30nfUqCYwS6+hwoj8J1Gp9RzxssCAnk97XX6ZmKAYwz
VVqd/zZ/K/DuI72rqwkzAPuzheVQB0zDvv83AEeo3W8vE15+YkouXTcSzziqiqB0
F/zzD+Xfjx8OFvshQRvPrYI0bCDZ+247tuhs2+8wLiekFjyf7fSJVD12l2ehgIDc
pmyO6jZwjFutyfJ+pyOhn1RtL4tNSALsWeR/ILjVllIv7lNSZD9OMZ8BmGP6DK9k
s7Z3qWXKUoDc8DSNVH2NPv1NhagHR11PVVYysRxADE82qe9y1u+TE+yxv1O/R8ea
dqMV63GZqIiJRsq2VeWrHt/AT3DNd51tZJ3tVU9vCW4O920Bu5iqTu+pOupmbeaA
oYU6FzxMOmDLRL56gRVjecqIMgLMa8GhOSZvDCsjSOPzxOq5LVovOrIZJOQN9vam
zSsdTOeXr24vzkccxxvr4vOoIY/SvRSWT4sVTSSRPGjfAkZ7AX5KLOOGBg40Dp/7
aIl1pMWR6pmIT87vgazYZ8LTPRzK8Xe38Cmhs0dn44sUiFUQfKyiVRYjka8j0Cnb
Ot3qH5XCT6hRfUZ0Y9UMqXpm4magNNQJROQ3tWvDRIVs589xG1mIlRwW8qxo+7kL
PKppvYW+VX/CpaxkE5ywYQ==
`pragma protect end_protected
