��/  ������7Z7D]���-@�O�W�b��;܌b���A?����M�l�5�W�y���2D���4ø@%b����������s�
��'�_.)A�%�=�
6p�eڕM~�M��k1G�8�Q>����`� Z�'够 ���d`d]s/��f�ל��Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9��j�2����Oš�S1S�)B�@.&"0Ǵ7E8):��2ӥIA�jP�����ɱ�Y�y-,s"�N�:$�(�<��/F�������\�i��$c7 HGxzryn`�>n�;x���h�����!���u�2G���Ù������Ѻ����e�=��d�G.(u�����: �f~nCs�������}ͤl�[��V71��X��3,W����p��O]����:� �d`�;�)�j�T��oKa��4�*��4��_���`E'V�B:�t]jt)n���)�'5����ӻh�2s|.|h��X���g����D� ��@�t�'wU��Y��1���^�<��J�r�F!��M�Q��C%d,��a0�GpfQ�hF71Ò�阩���DCF�aԦ`�HU�8�N��Mŝ�T~`;j�<Rp��2�U�L�<�[$C������*n�����v�����I��s�T�b��E��h��0$�S栕xw����a	&��+]�lK����=?zk�@Jg:n%zc��~'�$��Jy�m�� ���=}d� ��F���$�V=��v#w8��9��N=|�'�;^; nr[��6/y��o\��X���7���*#�+"=�F�Sc��ΐ�'*]m�հ���;�Ck�{;�1��ؔY�/C�s��d�F�vʃ��ł�����3 �'�6�ܦ�1}ݒ�:U(E�-� �*H���� ,ߴ�d�M�i����n��@2z��D���*F;�l��eb����`�N|�/7���3K�����(ɑ12R'�X��8���GD��wTTdJ���.2�BJ\,�۲P%��H�7&m�R�B[&���X&�/���컟<�L�