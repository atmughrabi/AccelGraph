psl_clkcntl_inst : psl_clkcntl PORT MAP (
		ena	 => ena_sig,
		inclk	 => inclk_sig,
		outclk	 => outclk_sig
	);
