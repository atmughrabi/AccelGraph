// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cULHRZqEG1+REDjZgXewuGryy89NqB+3/KsJu1zpx6FIq/oLFfTCSQEQKlod5ljg
/aer533mAYocRmRZY+goh49XqE5uVvkkMxr0EX1clExaRgq+PuAqyBMmzGDY/Xzs
k16jwmw4SmxoDz7egsHuEybAq1W4i6YJVarTmuf9/t0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4736)
2Gaqh7cGEaC3g4DJujrbTarzX/UCbKoyWO4d4c8EtcfKFgcvuKP5DJerTMhosUHH
wmjHJT0Oipjo7YHqselJ3s9txk+XOdh9yAY22NhtPY4rof6cdqpPMK3gNdroIA1e
iuPa/tFhnJoo6MN1ECcppjlzkmy3T87ykouWtjNUmtf76owqPuQwn6+H4ZDTicVd
rKf4NLTeVuAshtQlRrSkomves7/sr0wUMyqshGTo/wZGdWL02Taf0tR+iz+wkyfp
9kvNlBkR+O8s6HQ46kQL1l4Dg/kpFOvyudoZkytsuiA6Bm0P0LMXqTTZaF8ICk8B
lZzz7R/78nRJQKVyTavkStriIgHD8mPrW50GfRaseaz2DCtW9moE3/8Bi3HeJcnX
5+K4rc3Fgnjb+Fi1/AhZldQVI8rxdk4ZhSIJQBY5I6aBGjfY01j/l0nzybPUJnSH
HQ6vwH+HRE5xGEpxOHI/QQHrxP9lMxVNuR0GWtAK3GDQsVnrPfuQTmjKW85EJhS4
3YlArqr5COpnofmskapuafUCtNo/dDlpE/4oJpdULe8L0jQk2Mk/kcPm4Yp+fKR8
/i6bK4/mATFtbMBpg+yHj6EMQLrCCuywaB/T2lL53whR4i7o2mTSlFocR+qGZ6lc
UTwmEsocZamDP7DgAC94TMgOieYklVD/iOsV56vx4vYVKzXfpsM4xHnjDaf2bNXr
kfSRLoDQ1K8sNyX5y3kbGJG+dXlcFFILAJceFWXmyGcRWk8kY0//+qkTSlBkGDrG
3DJCdpxToHgfIC7K+urpgbEj5pmmdPlS3Ym91VtGkAuLUip9SFH98T1x9T99+mCQ
sTzsUPwGrsJtK6FZsS4rSCWw6F6D4DK3uxZWW2Mm+srCMqqGH1wzN2n2845YXpvZ
AQrUebdde1HfqDOEN8LLcpJCoO1ExryStO2ZOkCxb5/frWCMOXFqrrpOGX/gxOhL
UzgmiJyVx38IAIKVsNjmD3FiiL1Ns2lw4aWh4OsiPM5OMYX1YlAbOvjo8p0LNu8A
quXtCqx2+3WNH7DUVFMqYiEVJkCwQ65jbvlNjZctBKI1K2QllBEdWv2nH+FHxwMc
/qfYQ6HUhPTFxduYwiFmdDFK+83cperturrH5OVi/ZPJ0zmxnbE8Jb9N9YA11e6L
h0JkTjPJ97oh+h0xNfISZo3JP5Goxn+80bWZhGrCg74JFY1kssr5Es29HqeANC1k
OajSciVl4cEqQPjc2WOZOmLlserAw+HO6aM6mxFvBZHvgwQwA6f7Ytk2cqkVv42/
8W9YFm/GKdGCdV/SQvYQ1/sM3BB8BZljH+YZfBm4+spZqdCIItESXKVDPeGhVPL1
aHOjCjeo9D9VtR14xISAmTbGK/NAM/ZpIB0SI8sd7xB7AI904clP79ZGo/GtzNKb
EPHiMS7cD13TbrUNGFoMQvaOU2dA4U7ujSe673w7SOka1r9hUA+I0vcZX/2N+haj
7AGBhqYTZ2vjFRmHKlkWHhGr2HZsm3caPFFEn5nZ3LGK7mXFDx9JthFA8AYku0OB
XA/JWzdJ3FaBXg/W3rR9AApr2Bsbu0X0vaZFL457HLo3OcAcCimK/R1yvIVn7fyq
G1BAg8KcQzEk7l1MQXEoqGDFGDliRpIQqzzvtbl0RXoo78bvyWd6RBGOM6oXTELt
R70sntkG1F5rLGIQYJC9eKJ9AldPUWUByUq0qa2mluYB73tlVn397PH8lYlG3n3m
uj/yUSum8wUBqgHxH+Skt53hINe6rOZoLlqfWhW3fPmcWjjvziurhVFbp7pUDQea
QVFalQ655q+fqmIQDYQe2UdMne/1Jhz47fHmckqW9hJv2NDoaH1A22CpZjRgrxbG
dpGYhdLUzfVq7+KsK2g9HfXwLulbys4Cfeso+T0k4JgymbsuqjSV1NvGo8efOQ8w
N8P7/J4p7I6H+bfw5pfMSofJlraMLqhTRT2FhrxmlByqNPnIYn/e338BgKldbWqU
p869dfSNU6eEjUJTYomODjAG7XIsWHVGa7wtbnH2j7sQki8kBAGgkIvRAbnV8zJT
VMIFYkgdn3+wpRuMadn4jtspmjJV/7KVvf3E7YE3WAWKH7o/bKDzveVBb+k5gNPe
YCl8Ya5+g+qtQWrkQDflxzCpKQaoi6AZGqGH1dypVMRX5fMGbbmq86WqWdvLPNff
sZQarkYzohNUXjK2cRWHLcWgSMZvJUNu9Lh3q2W800yjEUYaLC9KGv0ZT1JszqL7
LLgBXbU/wsdpXX6o3zYnZSwW6m4ZekR/uhyiqqEsspuRMFaEXhidL4Zl/NDWUz1O
IRHfq50MWL8QyGQtS56ydjBhxCgFK9gxWyKKh9oeeg17uXUbM9mXav5TMEnVHljg
GccBj3jLlQNL7nmsdmlFWrAMfUNFDfBHClp5nW/oERO9uYxiul6si5opVDDWvh1U
Dj5ieseYa55gJewgcQUfQ6d0Wn6Qon4gvR0GKJxpuethW+a/kaDr6bx1pys5WZby
XTYBVzzxgNZb6at7/iQ8UivUNiL3+R4SFR+2D2SbgL3De4yCFncMKQK89utEQSXt
lRy26aDllpt2AzMATDTvlR7+lzsd19VkzJHnCqoTHAdGeG6KX8T478deCw1vxaiJ
TssxTkDrXhI+z/UAsGW0756csdWyMb5QKT9YsLRHa5F+k5k+zU4dUeAjdLNZZUb4
BCPRxRe0hvfbShvXZTv3AXoPSP68D6HSAk58KbyKSfuWthZNjl3LI4RI5IYrH4/E
ZdzdA9nzfNHqwNdZOfFn6CkpmjH5HIz/XnN53GVuLZN0QzXbJMREUX2t4bswaJoD
yCBNRs9Sn8DSROIrbnN8KVnlW/ikSEAcKzOpal9UvL1n6zR92DKfd+kAHVNEirul
JtPzDtGQjoLP9DwbsdQHSjmMSU9+6ra2e+QdJRw4ZmlZO0JdRt5tHLijWiA7biNT
J6nfevT3/218oznmNANZZ241Lmmfkw4DpskmrC5KYny3RplNQVFwMzDgm+E8Nz55
HW9dKuZSG4D1wuciH9kSSedvVz9cN9IQzeNyScuic/tr5M2JLgh8oJXTOhfZh/kl
Quzq0hvGRJTYlB6Ax9FfhHDDOqXlkxcbReZFQyq66tKfo3C4/iln/vwZyYe1khIV
Oh7s+oyjI7dE7OxcpGnmZKg55/sQkHIRfO7pMrgaIJ+DNvOcpBwE34v8ZhYHqnXu
AZ1HLguXpZMdyyJfCNJZU0s7fVWumodigWMbJttD0HKsevqzVLsHRfXXbZFU45RF
Mf3Az/pZKUtc9DbVM4v6TpwJqpMj12xpPnbI4ynOMypWH3pWwRZCxub7Jo1CVCU6
p8bgql0fQcKfg5DeyWpwMijdYII71+AwKav+Br1vOCehRVXdnvIjmWavQtWvDd+r
GkiVMvbcUOF6OxGPW27VTGhYaRTv3joB+uZZquN37v6mH7Lu2bFHr6aSDmzB32zp
nOHJrnCbPuCM2aR4efYJpDsJ+CmleUwWbme28nuUqbmo2Mw4g2oTJm5Fg6R+35AF
oo3niWg7W4yX9hebfGyDG7ahuxNb7JsSodme1FE8QnF//B4pEXJm/8yuBOL2OOsb
6e0s0PZEFM/8L7qZmrWkz3kerOm+p94bpQhT29M11jEMwX6y6cvGDMwV+9V1Zpmd
n7n7uWWYLw2AXmKRmSoBp7rTvBiWiMt4+CstKMrL4ZgB/TzVZ7Lkki/816CuMIpt
dBi4FTFwU/MY+fn5MsAAFzadbnDTeb11Av7UeVQ1Gnycs5z2ZKwkMbn35I1mBTPJ
0uI8/KhLQwqky9rmSqA2de8p6pW3wug2ZOZHxtVw60dTnnJBDwIPYxjXQNMLRUmr
otbli9oDZJbR6kFU0p8xXjPCNs9HX6S2RAJ9QR7DbzCuiCQw9FdVtFLSi+H+Po3c
OO4aBX7txFselxJX/8MHTAAszryIXrW+A3B5l6NpGPzTvIei8JtpJjxsAtwP0MyJ
1wHkPphqAOQJvJhDj47RLRuIG8vdBNKXpWt7fr6ZLvhr9KwLjGEz/XyWBEoIm4b+
1lbmHStXku5/KLWq6KFJSdIv0Iz+KOrb0XM1suuL9QfAnRy39gyIqtveq4sfSFiX
4FKH+0TWBUOuSRzEu+v/lpguY1GeVmSW3cdNj9cFCdIFANz+gyY/gUZJXKIAhCWt
Lw5ISsfdM6yECjNEWM4ysgtTgoMwNLHAXnKjAUM4EkGbaGv4GmTA/6oj2jCuKT0U
PXcV1RQhQdFZ0u/u2ho83C03WJafivpBqXy3YP1JZzrn3GsPKPjgVctdt/+lqT1H
5E3jm9gSOeg1SSJYNEB2ZCYEqFH2QZz5MRxBFTwM4WqiGjdEqwAM2s/lAGa67hel
oCspCn1vhesOhjNus5ZO7p1xc3NG9+ArjSron8OsqOINRB1LAm6YEn/yfGIe1i74
fN+g2kgP7d3q5wZMai68zwLtoQA3kalZz4VJbfPHRFVRLo3pGX0WQAfxJ9LdlPBw
ussxVyebKjB9qP8I6cgSMlsFWWl/IiVfhw1lii1Uibass4PpjZs4jzhrLVp0cH1A
xMnpYsgGhDqfpJaAhmK4iVrn7yfEBhvTUi3am/H7dOm22BFBGn3orjpg9YMbpyzH
9br+tOl6Limho5AC9J+nZvJVVTLm3WlehSi60HdEEOE7eroBBqbTpQia585CF1Od
uzjMs/KweRNm3aleZ4LArQekf1+O9H4TGyf3W0F2cIXw8hYkxrNlj9kcS1d2LVRr
Ajj8LrH9ZfUfPBslM04YD+OpXqbBy0KA/37B/uw4cmBK/ph3qbrRoznJXOZsjuq8
CHg2c2i+pTqeoeiAJzK7FgE6C5tg36vcelbmzsQ0vcGc4N8L+z6dni5WZPN5GIx+
FGg6EAh7YTDAJD3PCYx7r4s5btZrkrLgUeJ7ywU2roug9a2XkyRdbLAqBI+Zlw9e
4VYKrq5AKxrOttagV4KI6KIswFRxdFt96U8Vx9JrsteEcIeQDmrMYeugMrlo/u6n
HwkeW0+jhuS3wdraaA1PvNQpd2F+C64oK24QhQe8XPQ2etmvKom/wkXa2lAENVOO
YncoMCm889tfI3froHQlnyjxlkWMZsNZz/jg3etDQ/O12hX/ukj6ipsn/M5T7eKm
j989lANR1tKZ8S4/Axd5s1u/mz8m070O5h98ftxsMgdESetBD39Iv5YVcW/RbTIT
/RiRDu1uZpl+C/zMYr/iJIctDp/ARqrPOFjupklFUW5tNgcsZ/HdHsH7FjIBttyC
9HsylOvLeCJV3g6Vzz8GNLInv40U6YbqJDQiK3UPosooCWyPA60CJNMvh6d/IVhB
YJKLVaQcfam+IjTjUKbWZIjnaNazVFk5YDDCfSTYRnMGWy4/ar1eqk7oy7nDatRH
Dqlt3Bl5PuyBg4a1bqhWMwfmr9F67+N/FXCzVLl0y54fpX1yw2Ymay+k5LBKpz/c
cYl3dXqktIYlFR6Cf2cLgRYGIkP0uScnix7D7P5wG140Pp8ICzVYBdUWF3jvY6zz
gXxyFusTg8VmWfAH2ITDmjCPePvnB3rs1OXldIBnCogOhYdcf8/V0Lxz+yJFaMxP
t8xZjckcCOyA27y2reLSln79ExcNnbb0s+9EVt58eZ8qbEQlRMA3UPgWeg2PQ8kJ
hAJlj5pnWTDu6N9O6P2WBcGRC6JAcd5VtU/CLkICmPfPQfkExdlXxAy1SOL+p4Ho
vU416wgtRfXbYrDEq81Ukcm46BMpINqQq7rB3FHTn4meeaDDDSye6dR5MZKlzOd3
pTIAbQ3TFS2qqj0Da0X1cQYYDcb7AiVyQCP9FCcW2+HOKVZPfIsSEB9VW8L5JD/R
/HFC6yYL9uugwgAlr8ko/iASTTUJKDAvRykYeXukAPSkqAyTZJHC1YR5AUtFRBaa
+KXvk4JCDZ8hdAi7iqhmqTgKsQ/KilHiru0GxPnterPGNARU0iAguBWgs+p7Ho4i
Y321DeccgJc6Smuiett7tPNR4PeM86EDjjrORnEGgGtX7/r/TFk7J17gvo5AmdHL
43/fRu+l17w3SSckWe5oyBiyc3t2adWWrvf5lNP3KI1dYE1RhGvOzs3/fxuozpTb
xzeHUqXuzws/fSrGg7hHQ3U5j38TLynzvYvUonAQ4/s2U7T8townWpsMatA5UebI
hYiqieqlJbB80pT7udGg1MZ1KxTZxP3+SK25YoOMlgHfrtMdpDBbST5mFpmU8d82
R+6JcNtXLobes3C4qKi9ocHnh+PuGlm8RXcCb7FEg/3KpyPGtCJvjOb0622+sx/b
lV1fk7Fmt2B1pq+dV72px88NHANsRGGZPfHhv0YCNBY=
`pragma protect end_protected
