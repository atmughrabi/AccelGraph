// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
W3z9xAGi7dI/z23D6CNVlsBlfWfH6B1BJJ3yWXjcFCmy22QF62g/JyEWtT4jC4uq
ntB2O1wL/c5ySswf1gesBpQnvmB44fhj5nnYyCQVe7w8HOX/aCWst8xE0xpYG3TY
yfAYirOSRFIEKzr6VFXf4sBx308XgCJhVk9Elu4shNA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19344)
9nTOtqzXM2sdpNuTSrAjwz2CbfBeObErrk6QMrk9AbIcMEL9YevwY2vSb+deY94W
Dt5Z5Y3/l+DjllV1koKJfsJWCtgfIURQB9qnr+uoaK6hS8RD1kmAqtdFu5YfpfC6
KZvfZqf5m6JYkx/cPv4UfgOe5nay0yeKyGEvIFFkMvzCj8LmEnOfaa3xJRoUyqcp
Q4k/9IuGVO1kKgT43o/ymj43P1/8lqz7wZC5Hu5JWHk5dlS2D3x2G1jgJRND6SiI
AP5r90DSJhpzBfnDJ1HzWXNaH//waGPRKasdiloQVbY9o8Uj48pVTLgLSjjlOOfl
CuaxHi45yrf7t2UC4wFDKhw/lJ9DyPXPVBm/bpTojpru6W2wyPZ/SgHHh8nSg7bC
GroiCKs+RDZKmmDZ7o3Eck0GU8R/++YwfBtU6S6c2GZX9ljwYLlzyQABOUvogb3d
lmiFtQb5o31ULxTxlAEy3rKfGBZt5Iit77GM5p7EKCnAme9w/ROK7xUUY7BsEo3x
am0dnOmkzvOGqp3awMojnpTY4m1KIvkSxAenohUuTBN2ZG1JUgog0dUoPGOQBnfQ
QJXFpIVt5pDGsS5gs5vq77Mwgv4MkYayL9XHQEcRsCBw5TRcPGf5nUmCat3ze7Sy
PZWwf/aGxRIogZIUSZlIVx9+AOhEtb/7/VbzvPLR7hsRoLUBHxT3bFgGhCQ/EiYf
bib4ilLFDfOtGQjWQlqz09fzqcAL5R0lX8H2RfMWiL9sQoGd+ct716wry3itOjAw
D49zGNmddPhhYKDfY1qM/ij9M5L2s22sE1LzN47qd5SkNpk4oFW5N05umnQ2hPdU
dK50yYjCZGfwhUKhpuSMSutFF0SFQw6HrPcepcs0qR8zVeXgWFLGd6BwyWhwohga
g44QRmBT+Vj5eDFADi9VKYp5Cdedo8RC2YOiOg+jibzfFdjOuAMA5hSqggTSnFR0
jU80H7LEFVY7AMjPz7sIn3F9voBhqUcarTMtD1+dcycqSQugnxmPpKdHYqk/ZKw5
wp9Gc5V4oSsmoWNemZc8OMhqr2XnwsEWZ7InnegEbMMVqS2OpV9oDj0a/zivhEI3
W8HNgZKTRWxZJK/MQYV8toqqjem1rq50egWD0RP6KezbOxGhQWiU+eAk81BH/dz/
L4jwPndvoVXOsC1s4MP7yboczpjs8brJFnguZake5pX8Qpu2U/mm0R01VjdmXPqQ
m1h2KUjGsOcnzQyJyi/Y7iUZt/wnE7+tFTudO0zRrGizeTmIj+GNSegnp7WBAms+
akQcpQJP+eaWuCrD7RVuwN0YzEmkErxqXYXKFUml5YDyJetBbG5qrFX2DkTUUS2a
/DtPbIfNhtTSRpTsrfxkscwhoBA5kqsAuDIPibEzNib0MepkVCH3LqWQNfgzxeeE
T9KqqKdYvP8ku6MCL7G/dLbfMjfcYlWRlQVQJWG+pIntHflcoNgezv/EiRMZ+2Ol
Mu3HaKnuktTMPclrMuF0CXuqqFUeB+cMEiT77iwxYGm48XxXtOGrdkeOZfUnonQv
pK+2t7X7CbN8cZEmRFXkQHxHN+QStBg9J7VNKjScYFFJELdN281PBHFsV6DgpWnp
FToRXBMtu4IVfvNjO+F6LmOkzVmn+B3zfBlAfe6qaSUHKRYMlIgPf6suko0Uu4h3
Cfk5Z+desqGvnUxTsPhGXrWB/XO9zeDDEDxu4DXZu/sPyceEyG+0a1Z1z21R792X
VxKckBxtlT957KrPYC8eTZd6tJi2vwNOlsUK+FOAZfElHf7+swkoKJG/0tepESXH
0MB0iCBE8N0rItMbo5d96gtk/6fdtR5nNmogSaP3z6kQxDLhHXPZJ0FGG2nNsRsr
LBqhKc/65g5UR/if4mL4Lt8NX+aXe7/rsu+wc/J2E6WR1tAeb/+vdQmCVpqcc8Ms
EK/GetZD78jnd5ZtXazyGgFN5a0DtVk69JaZR8/V2hU5ClO0Z0ImbkVdgyWtAfe6
brf3QX1sM/boyMMDLru+jDk3vrdkWjlIJZMlB7ubNewusNCff2GLb6QqT2mNtO1h
DTZAPlU26jham9CkqE56TCvh2gUfb8iLb3EmHrzoZlsuZhmRGj/ekOwWz7F1lxVz
539suzro9W3hAE+Dwe/myFvlrckKXYu3/CByPakxAJE5aE+21k9w2XgEXTPHpg+O
7syCP17IE3pJ+YBtsZSEHuLPBi/m/x0c+K7E9bP5E6ZAWdDgV1waGYrjr7GUIYpx
TWeo5944xFFElBcZ9QGgV9AUXZFl76aOxz+Yhx50fALm8oZGsWSv27LLlP6EoisF
vi+hUonIHPgKEgZprwuPjCIJuDsCDH9TEIig136SC9nvGR/S3DCFBlMQoINthRBc
QTVX6bFnaP2zUY+0CaRIe1g3ZWeAEDXFVBJdM1OCQL/PMbaQaU7CTUZtONzYOICG
gOk/hU8dmrVnFr34Suh2TB99nt2BpEJuIIhQd/cR5YT7aatkxUJtTkvFhoRivQPo
yj6/iIGgl6li/ZF47k5JuGS3XaFloWzgT66DsXq3GyaP9yaM+lvIh6m6xH0iwxBZ
+lMyciLRzoxcs9e1vbaPYaKdwP905pY8Ma99EMSOsF/GSiC/JFyMTWDc+9X7tup+
T+P0AjkNjqDPP1dtzuaq5Z7exYvb+W1MuRo8B+EgOJupaWg7A+FjIeNY7ptjkzDQ
xfsY/DnIFYJmVhIFLEPR+C/A9U0wFBkcZ4x5zmqsoPSGW+IrbIlQS/e/cbSGynHj
wkX/LdfQMtNKbrphN9Ov4o6ycqXGLbZUgdYS5bYYUI6MVdWWeo/IK279jMHY97K6
HDLLfHVb/fvqbmuYmW2Tts0GSTrIcs3N9FpSXiqBo7CL5SHbGcGSvYV/JgW4Um4d
4t5m4sTjbKigjwvl/qDykoALrKUCroBEu9dpXx+AEM1yHJlL74kh+Pftw3MmmfQW
NWjZDONTYB5FB4YazayCZxzprJY6S6a1Y5SoI662mIkrrL2afBg7v66Y6VbdzJyP
+6wYnivYmE9+KYvoRD8R33Lg+0KNIOwBeD0tiCGJhpgdPhgO8g/DoBI2915h/0b8
GjtkesIeQrtyZeOEhyVg1g1W+0jplRiHWF1Uarp89MP85fLS+px3KMKIQIcHOcP0
kOzxpuccM3+F0AkT3PxJCRJuJTpsIjgR0zc1WXM7vFZlit92sTYTJeKZbxXQPneN
RK+sMZOtNWmb+WaQaY0DNvxVR3hnndgD64c4dmQyKw6DBPqwyE8zLzkM7gZOeL+c
XGf4SbmW11WSTX6BplrGga49kQW5jKtXY3Yw/iz/JcMqbB9QRdex3n8mWvrmrdYX
+zLJTEPDHx4Wmjoab2VuT2G+chgi2AySElzqTb35cVI9Z9OL06UWL3S+PgUAFhWy
oeOlDGVQHHRvMrKA+MLut/cf6H30P0WOrKY7nloHTSdGUH/cd3R3ZSudwKGYwnw8
M1t4xA+IJt23xqUB0JLKDOHsByvANPy6bpdAcsYbKCWU62zb77db7Hm7u3qDAnj/
Q15ZFRFWxhMuZ7i/akARJ24/FzlDe9wP8Fs4/WeJ1Y69nDZXI9iJIg3ZUfY2D12f
p8I57/a7m5UOW9+LCL9ReFEPHpU2zIWjKBpbBE2A2XylJ6z65TcbC+iySgWW+iw4
SGgpP7/sTHH+q5x251KBn/kWH8ATJky78UWnMuJuva/5Rvj6ogRHuDJ74ZtyF24+
3iUGhair0brFPWDkn1AsQQqt77r9psaX3eKlCkak3ZBye8jEZJ35sO3iYVUsqAxX
0uXhCeUqgUQWS97ahINHl8r5nCTsjSiPkgO6nwCTySoU+Z7KDORvA1k8fzAfe1yt
bcuvp2GF34bUe6iF5EhKVP1hXJvWaqKyLxbvMVmQPRkAj0H7mnOvB4dL6j+okBm4
ybqxXPyrgDFJedjlv0YvlaEyt0juCt/oDZ+/aojHwQ01fnlKs2K4wL85mnarqE+O
Gd4ZUjsDihj39tKOZrfXQVDWkWMNf4Sb+HwJc6LF2kKB04VgRP3/XQdDO21qUd0i
FNh05zqTKgn+vfcfvilkF6U4YLt6wjmMJbGoTfalo4fr/7w+7cxGjI9cW+GH0Ot3
BsdtYzcP/ydX+uSKr6EDyPshUs8kxTkOZ3FxwLFvVwA3hhWTvHVYwemojrR62KAZ
Db6KVCgoZ1bn2DKyl9M1zgVzwlk96REb+Ec7kHyOwd6QsbwHlf2+toxavhTHBrtn
gY0wPrSGPadgDY+SkM4Kxf6ebV8bwOws9ldDnVsL4OflQcCZpnBwlftsNDnxBHNr
+lggOiDhnYJbEECpMI2olkNf56p7MbAAr0HaAWGUo3e4q3v660wSnf7+JUwl8wwP
r5m9ugvbHplC5UaqeW26zUh6IdzkKhj7PM9smiWHSBcBhufZjJOWHAwznWp6YUnM
cVWcnbMMLAfasCzCgdQqVocymuh9aT/7TAhSEWvb1+8bHjzpSIaNJ/sS92GMxn9S
moOYeDpDYcIUPh8euplJMZHbz1tx99hEdmlr++56WidgpCaG5ITN7WDJGS4/2NmT
UUOATEKhXXpBGmh+Pa0qPhTnTc02GY45tsUAXxpzhaumcMQ+bSXiYUbMcXriMRxZ
qDkGEab0Kzji7/MrN2UVrE0vrlDQYYUW9uhURDERmHV4DXcY6cuo+xyOnSpKgT6n
L4ezLs16z9rHkHsUZ6dPIl7fUHUeUwC77YiAax4DcbrZep9TtKebuSBH3Mj2XJr5
k0hRBJ0Zbn5pqSsjO2hJFAQDV6kmxbjS2YYx1wBIYJsVd/OSCRmknQDClSmlFAIb
PX4fpXepy1+MDCkmWRm/DEnwKSuayhf/cmo/b8+nw69ZfkKR3kIAjigpJaQlfSHH
RtdY9STpgE24g5PTHsl+oDItD9UxqBJwuz7XK7cy3RpUW6pnXQQ6Fk9tefmCqvCU
om3wMcppFIUcxisuawlZTAkNHSBnIPgaUo2ERmuUi8w08wm12WceQ6sg7IUVB/9S
kRe3QDLSt/VVrX0I2CAJdWnpFiJrfZYk1vPOezLkPGj6T50rTnXl0MjnKOH+xkE9
rWk9Fq/gpOs3xxPGsTnxkkhusN8vZiJnPrILjvrNqeZ7hOTSbdyldHZLhBALutGI
QxG04NIbn45dl7ugz1tePyy1WmXNQi9TjmP7/mo4nnCHJdXTN/FYw/CCtrKiO3Ik
azqINDU9vFWwOPqKDlClJycwpWeCyus2b6js8E9xaszBaLERbbQMzXQyG9pfPoJr
vnaAOy3b2d+Z8K5mFiNSDlg2EpqpPJCPkn/MgkNHPzggEGWYhrn8CuP+p86rC0Pa
hKz48ncXWE3k5wZ5Iyj9qFkiLQME4O+ny6M+M6aikvsW3WLIF8VstssZu+Qa7N5z
m0FjIeI5ZbS7xSxHOk4DHHUloByaoNISDDIuBjY9Y1NYHjaWbprXNEX/uRwZX42T
Kp+ufrd1ezDAM3YHwVWL5332+/Y69Pt00xLwQMWjF9i6Uw0tNzwTHsvZNBNt7fYL
ftFSHqm4g1HbGpj12FlAogVEA+vMfu2he5hwA+NZv6PoKguZSnckVwNEuib8aS5x
GFH92R1DRsHL98/oBpxp4MtRAlPEhkZjBAX0MFFZ5QWJBqpmE5kYStE/SWo4oCma
oM6nI2CGcgyaORaFJ5Uleb7rWD2yzU+OJdNvZ9HEcEsTWZVlM4OsEFp/C+5EB0oS
DVpOSQEwfNrWU6H2HAgIeIzCfwp/mTiP9EMlzz4X8HPsaM5qWIe1QFEXrhbnPrjd
3zzBV/ozeGXZ4LpYwfHo0MknlLWBBq78fJomRhoms2Ec5qke8xOm5m+a9zc45aOr
bxrgkuYHy2EwPjt3RRd2f33Rwz9MJSi68OoN6dDOPH1G/6WE1g7850vXNpIXccLa
xdbjWbCQiMqdX7QW0fshKRHwp7L1v2YAdZSCtkvE0+s/BP0rr87CAigiSVQyAZrf
SUugGRk7qZxVm7jV2qNthStTvXUIQE9HxBaGgzk2kmYlPdZp3F6s/kTrXsY+VJzz
cNoHVyBpGoOT1HY5qu7s4fEUaKO5fnk3bsjUxhHEl+Yvsqs9S3FxMIXj4o74HlUr
TwJHc0IvbOSaQ7dfePhSnSM55QHoizTrb5mR8eNla/vImNUX/g8RfBAHLPguUwbQ
e2xlSr2LpsC2GvBtopDzUSdRYB3A43emXlLR92lhja9jagE4cwGd4fJ6Rjbr015N
st1OvWWWACkuiSFIJ7AB8LrYAH0IqOaRsqruCjad2rDGUQbhxEEx9i9Lx3CkpNQP
GNwOPXKyfKEJHx+0c7zz9v4i20ihhZxwSSLBzeXtMg8b5+aCfYxJmXcYP1RlUKTn
5c3c0ptu/DF84jxCp/WlmFXAfEhqwTDt7Lg6Bwv34ag5fnAup5pm/5F8V9oagLgA
Z7yng0LA5HqKifyLBIflN39z/YNes+INUrE+umPhhcCLYvRV7AkEe4AZzeA39JVE
/b5YYR31HLXXn4ogxpsBhehq0WSuMzhGXdGvALSKgxJvY8M0MTTuAtx1crupgWYT
x1nu02vedOaU3JUdV8i2o333fD6oz+utcVf0aGS3b8edx8fJtl2gVMJrdCO47ZI2
z/8M7dH45XQXdKCmflM3BUeeMqJkaOS1/nQQXzMDqJytNq9ty4XlPnKwCLx9AzmU
Y0VjxBbaOA/1NgmhnQkDs1N1UN/gL37LK8FowUcntF/8XAhF1XfgeqJA+4eH1adh
QsNw7nsbpH5QatAm2g2uEoCkITYWWsjwtAsd2KJHPSFn6DTHSCvogQMUYoheEwkr
g9HGg/4PsGgaM0mRhCtZp31wR58YgmXuQT33ZPmK+oxCCUota+K9kNO8veWBE7BP
m/pDr4wA35aT7RB1Ale3b/cMG6UqAeZ4IUWalubZMYH3uYDrRo9yjqmnBQdCzHDW
CCpoq+XYBd5T8ndSGs6Oj5fwkyoyMHMsYXhsxDY+8C520HjmPAJg21b0V9WtCzRp
dxbMFAr50U7KprCnWgzpbnoxICgonaC0crEdarJKunWaZtxtdlOxEY1goQJstet/
lEcqYw4NmZ5sEN/w9ZJCqG4Qppb8OlJLk25TVz5rODZIYAzkMhCr4bXYC6AhB9OF
4jvyzuX4UNMdvCPOV8YSy/f2/HDvP5/uK6yYBO7SqSEDefBpd9orkfWnop/QDCxz
QoQ4cJfoU9LyPDJwMMrjsCOx2KdP+K2VwqXPDlSghUv4Gq5LIncvgu0kTdb/h4oR
N/PrE2DHDFkzrtuDCXCbVcvNlmspTmGhYr/hXs3CG+abbvj8n64GKQR8HdBWZX8r
OjKSPN7Un0d16d814Iu2k1w/4X5Mhql/lLlFWyUDtV0MGIH077Wp13p4ZPoFdkNk
n1ppVWYeBlHIte69xB/yIOAvqPd9VkuZ9zJimRLZ9uiASF3lmUpb87ewnFKHp1/n
RV5DDAgiJxqcD3wDjTZHP8KVtoIqK+nHxSy5KVtZQw4Wqa0ArE6w0kfyik3mWQTW
pDCkmnkyDaynOmTam4us7Oy6UVwN9SN1Vs3WU63sisTuBzyFjmPvn2muVds2K3hU
lOP6Yjamb8VbKCki3JdhOEphvDON5K4EuLcVcsj1aqpvMGu06QQ2IZ4EKB4znEqG
CAp5Ghbq71Sm3xk78MxSvOm375wITknR2kdrTh7Kb3CaYC0QCfeYBT/qcRU2TynU
X6DJ6lAMK6tNY30s7WEVow7MvVkzLOPAN87MhMShrAi/X1LN8n6fisLdICzqGHQP
MT7JtcI2PtwKIKqURPvDOMqUY/4A+cYauz4E6ASNHxRVSLvbqV8AK3t+Eb5IKMD+
3LIymmQHKLA2EkbVfu3KN8hJxv1aQAiSkkcm5avi/1G8CZ75FGUbCFXpsXaB/EaZ
V6Hhlk0h6B9rreeoEq7zAeNPFDvpOZuXbXUKOvdSwWeQmcpgPUHoXJf+u7MSlX+O
/NwV9Wk2ddpf/8Vr2MguL6OxPpX+7qyFhCoRXy3kRsOym/WodtiIsCKKlNwPasYW
TyaNzbwNSPnON2PR7PBgH385+oHkSk+SVa49BTOTfkXciGTVKEO2M4xSumHMxqsI
UDP/shw0ZH+NhTnNwzGwZKws03Dz19Ka1Btplp0EbFCOdZ6eZt1bXEedTypVJ4gy
A4he+1Qph6hsbiFnOjSVpEhJ3A3nMnfitk5SRWzU/v9MxV7UP7ba4LVlctUDxXRA
MOxok4qSLXMW2qGHHeOuxny6CuuedXMP4pnP2baLcV39ltDPhZ2OeYC7WZBpHBY6
kLY1qIQvueNGz497x/AQxCMm7aNEqYyw6B0+ZPoaIs1XNTxM4cZhUoIY+aoJZCXx
SJmmGTfZa6OABvl9WFFtka9zGidwbFaxYO/xuO4l+EWTSvVvyU5sTrWuDalX+lmD
qN7WsNFBOkiviu5wTicyVSHLN4Hm++TeqXhQ77Rca6bJzOOcxWjNZtbl+r7KNCpD
N8QD0E+Q2lgFN6apdP2bSGpczNsi3ZgrZ3qXNT66I14wsJH0bqAA4yvCpTCkAKxj
mN+7NqtRwaIX6Ugm8dc3m9+Z9ampBCAjBT45EIfz5pHCu12hkoVFv4JgaqFxUr4+
6tO0vzS7zrDBiPnUIgS5rqdieHvUhrrnMbdIIEXrX0Z0R3NxfzGNQ1ZNSfOC5mZ0
R26m5rp4EURddIrjnV2X0H/1JCZfo7ujwhKGjKh8l9dM+BSPi/e1z3tWJrOPOFPi
q6STLQ0oJzbrttSYGTkQS10DOwmRMoY1iYXVLsNC4rFvQ3JOqLqltkmiGCdysjtu
WqIU+dwkc/yZ12LZxFtMDkeXSfCkCpV7UdVCi7f/eYIflG86AuQ4V0isz1XpcyTm
Nmo2WpZpR6dkB19V8QOWZAc8miFmOyHcPqq3Ptt7DzaMwBjGAiFNCMLfndmnZoLa
3xlbHhygJAdjagML+Xijm8atJy5aFdq/DSBljqd1AumWDjpNIPcOUcn8Veh++b3j
HSilq2b+INi7rqrxQEGRF/TIxujGJv1EGYLygLJJGyQhkNXpFErIijPfijzpD12z
rEgQDf+64TbjonGIcmy0l4sl4uNfASHe0WBxfA4mtbbXSJFrNVbz+rpR5UNlgoMk
75f9s3vxUiAO7cdy9hpou7eEiyv53XFdF6O/0wvyRoSWBEbKqgOWGhIVutn50XlY
lyiSWJSNsxoTDUbfBf6WAa5Kuy9gqTLLHsn4oZ+i/y264BffbEJGWLpgUD4c7F7x
w4SfMHEtyhI6nqQnUKgqf8pDRNMzDh84Mknj7C4fm/TrdWYprP7hUSFdZ+UB716L
FqmqSwkkjwPHCUMALW/fbzW3zm+OT0dpNxjaUFB023W0cH9qYZylaarEq2wZq+yL
qmzZyyytPOXsFYQo/IZ2foIL/BdPUgpEcI7fIqTUaF1Vzibmfycz7OI7yh/mVK1F
d3FUhlFg4Z0as2tavsfLUEaUT2mUAxKwNk69mmEgkPo3IlrnE5Gns2CUmr+Y/N+W
L9RJ1zk92iZj+fpeciTYhjpGMRzp6oisju+90GSgwFEoNx5+Y0syeg4XzSjSic8J
s+97qCwZmuOCRFcIc2cJXK2Xp51p/FdZQlQ1eBKsqR0EFw+QCLPaMzr/4uR/AyTY
myrmdqsJAWRuTt2U4ckg2o8IhOwORYMAq5HvgvwE5+9OcthBWpgud4gtg3Em7Aqq
KfVXRMvJP/bKXriLJzkLFQSmWYsLHf9p1xebqAhs77XAyltyOA326TddalzbiASt
uBfrotatEskNaI+0nFPCPzA55Sthn3s9EDTS/d+m7ZOU97Dl1oYLL/CdId1gaoPM
Okxlu+T5vLWdr/bRJovvELxOaEDrCtCD3f80/tSW4cHOGIKikywx1R58LW97PmvM
towzenKtBD0M73Keim3hiiioU7ZKQGpXnhgLJrkKxVQkd3jGNH+qqycyuFRJzMne
FhkYjQxj2JukUpKO3j8+tTaOpEpC/yiy7rFMuaWnjMYkGBHovPjaRQXCWe9/9kiN
bCnRp51Tqjw8vKz7qyNeWOcardsTnmZkxjKZk0lUpF6jkFRTHDYLKEHufyoul+0c
yu+HjmTDYNTNyU6Ec5QVamnNB+EFapjnpVHxVYwR+nmCwOAUjCUgwDJKhzSgekik
t9Sy7hx+9ZxJCUF9mj/G3mmv+0d9mRrL/JkLfcnnMBc5tQUIvkrGd65+65gHruD3
aopt/ms0OT/G17JJqNsIYj8zpgsiLZwPBScAC+DpvSmUawRdodanQDIx+el/Rl+N
IUFAsTRG03k3PiirhG9XrpUR2jO1HK1Q/KmBJnP0gT/Pv5P7LOCwpZWVIKTMMPqZ
an+gP/2B5MG1OMLvOiNXHTzqxLoSnH3ckWjIqTLr7DT2M6UMaMBV5trLlP9E08fR
mMwpcDVCY6Lo6apM9NvX+p5Vz+SviO5yQjzTZnaEuJUXW7UgmDOgi36tzGHp2bTY
oWC96ZGr9EN51vABg7WJuRKpEFGqNsS8CYkoy+6prKYkIU1aBAmELZZQswJ7thkh
oobXeYKOI3ZlJkyUFaR5BASVFMKLhcN7TBuzM+2KJM1e0JQTSEgUU/Qhzja6pgk4
KUNYeC2u6t8UkRjvwPkOEHXe2IlEd7xoIzzs5BS1gt2jVVwG6HnzHEty6mPHd8N7
BvYw3LTIaZr/wM7dGAi1CcIwePt7Kzry6dBNRcjgKPPgjFdLBP5vnFIAClREU2VP
DIKyUOTi1VIPKUSkB2+s3gytaZ6q+tehxnZwbHPr0x8/r5Wen2ijIaziM1ESeapt
TFBfx9hgnssYZ76c7t46cQCECo/qiu2y9WRuSStMR9kIpoadnSeIgjqNJoIDac8/
Kjh4vrs+RGld4q8NwIOJ0STD2bpMHMILBGB4yk+FUj3GtA/IzmdeqRneKAQm1lvq
ix782FMNC139q/Z6xW3aExMUh1zJSS1vxz/t4ZVCRVRzmbtMAqx5FNj25Qted810
ZwKNx8ro7h3Ows1t4zlwLEvw2IxoBDtY61sJaoC7XuRCjkLRUKazt0yI4CWjc8xC
Xu7pgWzcImfsxjogKMAiFpmlQNv9dCpVBuKVt5DrwXUU0BZFAzk2yFgWXb5IN3Vi
EY1IrR+MS1cP5Ge3K2k/rtJ7wbJ+UyjVmS5Y8e6KInR9wieykd3yVcQmm3h5bEC2
kkSXNwHlS0DlOXq10xNa7fK3PIrbyNSN+FB7nYZ3ZP9DyCkxRePl9pDq3hVc2zn0
wFSQEwlr+EC+W/6PRO6JwGwFaUy9e3X3IzHQcpq90q7SK5JMVLIISLTUFUw9tFZX
QpEpwN9YhM43pt9nFZB472tLJ00fcoxz8wfIpeiKZ4ioDqkukmpgg3y2Oqu4nCQP
nJJdBR0Q9zqm0w9TNn6zpe16Mf00GamFPEG/6PKh+OTn2r67odvDsz8FXt7fARXN
hUkyyOUL+BYzN7xPzCZ0MTeH9H+PB4zmhbXJBsu4JOQCIBIgdFxvSKvtx+OYl8Aj
5SJVred+iix2OLX6J7LOnjtv5nxA6ZcgH2YhakjxZvQeFk7xSKvEbdFmipvnMpBH
d8CFIHul4CrUIy+cEHb9S7OM2Os5/PhA4nR4VxBhVRUmABOGk7dxUlOSoYRVzTrE
MT9O91CZ7ZBqrKSjLoZyDjPis3pBIo7oyUQJk7yYos2hsm95dov03MqwtOUuhZNG
Qvu63C3m6JRKLgIUj2OjNX5wQ/nWT3RDeCGVvNPZ1SRpDVvO3uZLslJ0RPYEkCcp
ZL/DBL0dp2biynRaQV+CZ7iGfU/cjGsADNcKNvSXJp4AlK6eFZmX0ts06bsiTvGH
4N6qi/440vZ9ZvpDTKvIgA7BHF/uXWu7bBqKz24Ks0HgVFjT3fbI11znc1bWLzhu
UB+jSn9uopwsch6O0eyH/U5KJS0OhSL44ahH074lJ140oS9pXosIbOsMEkufIZ0a
raXp5M3jcUPg8b43gTRq0aorgPBuZ8l0u9YvnZ/zGB7k/nEUrozW99wUiIYmXiki
oVTkwBsVFzmgaNf9nEBcF5AMrczZfhtlI0QfCzjQTrCicvS+mmbZ2ZpXm6Xn8fWB
XJe9o38WvqjDLM4U53GINwU05J9Tpg+b+0wxf5VhdOnt+fI6tXw1WynNoE4ynM4y
7qNsi+WTb0wvlJ3wzrhBm2q20T4fWou7NZo1gkYmZvYoHrCzlumOJ9CHZkEXj4Tv
XbASBsr3z3eWZ63uCZ3x60HcVxy02y0SpONHFsgP5pt+K/Wh78OfJs9ifi0g5ybM
6/CvLN9e1ibNLgv0Gpgknson8t1QVuVNGZx0U6Tu/UiENw8eLQTcoAY/7krrEfWU
dzbbt17XvLf0n43OkJcfEC8c5nYOHsK4vYL+pdq69HH6Okg8h4PQKx4AnUR7W0BC
1BMornbvNd4kQTxyWogYQK47jhNngRLB0wjWbPXpi+oHLzYLoJI4xfpdv9CCS4Cg
+oi6oBu2f1ABMk9MSasuLvmeBYEngY9Z0wnbHL+rSV5ReE4olJVxui+IYkH8g/uK
vTI0fOLr/K4luU3PgfpvEp1lSnPQOcN9EIpByYwFhm2LQosWL0VKaU8VNTqrrYhN
LAHFp43vgqXdhilpnxGOKwllt2hMB6HGgZhyL3w45pVG3IkvAOYsS0TejgOxRof1
vVMAKIOzrBIsKcpKFtz0Wza8y15vVkvlA5ga7w4TuJAt6+yxKEmt/JAzeYezfA6G
T9nCIgXgQMBt6/MrCWFi2OnM5nHS/s1oEg64IkwjWpdMLvtLTaWch6TZ5kthLvZd
tfFiXWhnx1FyU8psTqGpVBsRmXrMQqlYucyauWry0fqi1PotZmO3J54AhMmrijoi
gffj8vwMTHUU0bC46qpD8U0nbCvhfOQKVx24Q8pnUmJwBMd7XFTvf5agMBsgc0Mq
5C+/1S/gKxQORRhAJP2+B0oRsAH5kKx7X44LjtjU0sf1pb5CPSdgKdYvfRu4Fal5
U9uCjc9DJULg+rLnMK6I+FA4E/y8s1V14L7sgZeIfOqjVphZj6et2nqY5Pt+Ig32
eNnq8qMZf5UUy+TTuHaU6s+hwHs64eCB+JmHxa5FDKAb/LeNA2GPQSHqmqcg+wA/
S4Vy9AXClGAoEVYntsg1up7z6VVeFrIbYcUUVb7lfoaRn+DiS8mLWDr5XPrpxQTW
FgP02swY3YfEWMVoIc1vyg4J+1t9FJ/sUprDVdMJA5Kmxobi0I+RsQHC+zHe7poe
b4y/wzGQr4so78KmRn8UPjklZzFaYHF1girKzTc5574RQzC6raXmuY9612FgYQAq
70b/Vsa4pb/UDdXTE9aIXPT4xFtbS2Q6RXSfnGGsWJvJxUrFbxOS1X9Q4SS4u6Df
FrftDhB44UCToE7/1EHapgfv/6SceTpU3TDI0Eb5d7GjRm0QF8I0CwmoJ9NsLpOp
LvZOmjlwoYlUBQZw/XRgUcwBaod/g9w0mygHT5AOAtkw+eamNat2ks9Zk+mrnHdK
ZRZBq74dt6zOXQiR3pEYXWw5RRDU1wqUxjD2fAbuWpAJuwKJIGcQxlCVRWFziYE3
JB9zgUnw2/h8dNfprOwt5gvi+3sSwZBJfntJehEBicYpKQXJvUcmLEiKNt9xzP9L
EkfjjMhPTCGPiybq7wfuxuBD/TlP3spRg8s6V0K1QFBdmxWrDWEPgd0yndm+Swl9
E6M9nUiQDCrq7UDYujBd7hBTimeUkjhU0LKBJ2inzEFJAPvGFni94BFgiWGy+Kwo
v3sjg9OM/JkeawLpgIj7WANwZHKX7R9wlp45Jgm0yfvHCUkuvpS5j50BIMoFEdRR
Mw0KlKwiMmYNQtVJ7OW4cuPCYykuZrn8hgC+4IYE6dbJC2btoDboNPU+U/WkMBDB
tOZV4+sSUPwJdXCusYVpEXKj2aCexukYXQDxJwfkl35+Om18F44Jkm5JJwGyMPGW
jwhSLUi5MQmQWBoMRWEfTRSAvN197H40XPVGRtHQTe2gGZqvA+saVzemrojqrQB3
UOU8bYoH1Cqcgs+hUQUHgBqMXvXGAkT1o0QsSsVyhpJM5Xnwh9qmrJB2alCPmyZi
rajzsXxxra/BlhIMlB60Jx5SHRYbCzPpkJiSA+7aB2uVYGxCIAMNb9rMhLduU2Cn
kfU6oFedn5GTdm9X1ElcnHbwxcgANqYmZPlccYLO+hIoE3DtWFrsRF5SuKR/2dlo
C7vHujf7xwjZEma5CL2CHw/SfpSrTllPWeIrv/BR6yy5S0GmQwQHEWXwe8oxrFKS
4NU88JZ++NGXXffFWXcM9xT2NRM3tpuD/aziewZESxWmMF+j9fAVfKh0dcFea9JX
5XuGGyqBei0lRUnOyLbUjIwGJ8r5brxVh0Ovio54Ozb8mujMDMLv2wgNlm6gSod8
YsFMN/omwbR8OOwHMxEx+ZcLYGwcQTRsDnTMwu8Gvn85dPixdtT3e0TQzXzbE+QJ
4YEIGk3cazRTaAEMEaHOOpiBnOM47ZFc41tNptngwikYGDfBYXUCTWkfdhU7KeBW
DRrZTqrOSvEOaugkInpF+d1D5slf28QR6ulCtX4XZGzn9sncROqsuYUCpkc7683a
5RHEHv3t2pDmnEobw66oetaKbJIeP4/WIUuDY2EbymGuQdt6BIhmBdG9jU2/iqy5
kvpvj5Iu6tBJJ/nMD1uxYx86KTenMy3TsxfTb9mBAmek6frNTSbugYUEQHQWXRkH
rovHiyVYrGmTklfjiaabKKEK0u1JHdmFUx2QbFIlr8+ygaIfqgOjhSMHLqABB8iC
3e1Fl9I1d69qsg198cwg3leCBGwNeUe94tcLcCNR4w1qzsUxqM/25+kpoYL0Eem6
nnd15lee14ADIG8Bl7xy+8oUvP3Gx6z7ZHTvyIppuCjTIhwewNFLyaMeW6heZJUZ
/mJHJdRIRMSsbJ2b8JXbNiXB42po7GH8EnIL+qQiZEcgd0v08fKZa6qsG/sqnUj5
xyvA1gZezJBqdXX5BhWy6mPpLv8cA8hIHXbiGx5vMbtYrXy6k5ML2q36ZaB7iLJ1
Yw0JD6QbLc6Gyay8WnRFPZ8Qhz7sYBlwQlRskEejZThHoCV44Ll8tDlGBK93iYXX
XAcO+/YuQRk3Q9aqgb5Y4Ba+zsFkBLB7/ppve7b6nZSLhh2vdC2LJFZW3E1GK7JZ
Amby4d/7/ryuqenjwKhmMfqpoWilMXSS3FRwpVn71Yss2UIa0NM189r3JApAtemu
ZNjl/UmltC3MAbJpELrXxftShNjPyAEAFiPSdnidGH97XU1kAkJdFB5UQFSyMOyK
cy2XgKApOkyvJWQal6MUq10NFqdjfHqpLOvQpmVsBqoroly6aGh3WXSPCwsCzxO0
u9ARxVaG/lf0AynM/wN3bO59kJd6JGnqbYJTyRoJazvaFZrEwvxuVJvlO4yIcReF
VTXBPdowfM9FbaiXkN3wKqvwIOOzRGJiw4fCN1mwV+fq7BaZxEdEDdCGme65jA+V
Q+OrkgsgOuovVQLmuZqNSdKxGbMxs/VAuUzLyczHLMjc5s+RkbDJfslbSq11lZAT
as0ZI9XZ4nDji4nHirmIVLDqUOggYfH2c6YBeUZRAfWXLZ3XGLHFUbUrw94zufWn
iUygWMwV14zPlm9MMYko6rDVgeh0YgbpVL92VBkKtJea8OrzYJ39UGawzsOFWaUx
BVpQrNd6dP0JlB7dGlgU0Hb0vNgtE9/SnHpa3IHBt8V6Mez5A1fSlVEcKCUOIU2k
mpJyVcNcBhaeAPrUJdwbq5Lxx0AMQu0cLYL1F7FiZEyTV5k8eAgbjfkjPben6l51
s88QVERDcgga5+ZcttoGq2vHyqkjk81mmZf5Y2Yzo1ikXg08woAVfVbJjyaKtJOe
6yaCwV6P8wA0DKJddlR5GAeAQo+Lf3Z0c0TTjQXNrkN/LiPAJ5J0S8G5rZThdxX6
RZ4sPV7Mqj9iX+2+2WMtpDnttrVuEjoRdQkRgj04bJZGqPPE5htbmGdWHABCaXD2
j/BdQ6J3NAnU51MJAM3Q/fPSraXDMh4gDPDlZXAFyzU6i7CXeS7FRS0AcTIjJMTN
JQs8faV2mhwD21iUHwf3HOC3KI7p1SlbXshmfBPUfcjInyIP8s+2nQng0bBhvLtW
AlIb1+3QdUFLPdJwIjO4UarHW8InKRZr+8PgfZUGRLuijIilj/FQHY19IfjtNP+p
9DwqYvulB1yd6dUzLguBc8+l65NBN1jmi8pfK928KBef9GtCM8YQsb73BhsNorc+
Y58mV/OfCu/DCWW22Uir4SkMkaimMrMrs6rJwbF2qNHMiwGD9u6Fvr/V3TKQiI62
W3XoWJ7Uhx+mzfF82kJPb4MEieRv0+UnUCO1loDAEngogjohx4a+v5ODB3hvKjJ5
CIBqBbs5OvEUyOOoP/zJM2YXIF6WbVb71c3AyUP/TZVKmMC1uHmeMYgnauIoHjSt
xH1YmWKSFdQ62uowfvmpw81CqKCJvFbgwT0pYvhkkeHQxQmtsRaRsn68HjbXEP/A
TpV4xYFbWfyDavbkrtUYbais0TAsQkBDuWNRZvEmUcAka10zd5PJpaI3qsgDVbHO
/Iy5Od/xKmMuqVVr8e+tYLUMEkTmgEABBmwPEXGJLKsO0f/AvDDS9ARSqGJHYpOU
3qn+HPNzVFjnUTcoDSmgGQH3TavZvgszGVsFMHXqM76Foo/Y4xsllu2VmCuXln1b
DtmA211xLVUcqmJllyapQECRhPKQ3YUqh4qVvOdRjppM6dWqLwmoNgG2zwfYWJgK
ENx+dgNv+Zjz3oJ1FiYX+DO2TTmupQ9jlHDqimejafJJgWQKZiYfnPXw3gmsV9A2
I8rNa/T0KY+AvtO8qn7xAC51UmQfmyC4/0isuh/W0z2+pjEj3YUXBmlEZUyv1/1u
TS+DnWooabHEH+fnbGEmyHdxEAKE+vo5gOXbPdyeyVwSsE0EeGxUC44KOVYxdaT6
1l5SjEYqFMoqR9L+CdIdR3qxbNmbETDaZYNRGHM+tEOaVOwf0VMnYTwgYlOMGOLO
Qv+n1UFLpbEkrvwQ8Po7RQmhQu4GiOSNLsfFypqiU5Tu0kyiJZ2PbYfL1/BYpOJn
n5/ngEA+71Ralsjh2LGVTB88jOBp8+4yWQDQFpV1fuEeA15pqN/W50nWxqxKNKJm
weaj1fYRaW8Ih5RagOxnF1NMwNI1oRN30S/FQGt/5NQyjK7S8jYuifmMS8+g+7Zh
q5jMWGjYQ4FrHfblPPZotQBfO2c4KAtGDUcJBvH9JDfNG6igCD49kkxoDUb26go5
2S7jzn9pmUBk0posD8jYW10Dn5SL/xYQzPI63IK/QWfO5XS3BUX7MsieJpfgM1E2
kHLdqR1Bb0ZLRjXsgBTdIGJTANQ8Uxz+xJmPMc0VAMDCcyplOIQT3eIHVzvuVJzD
00ALv+yCmBzRhvRrePka5ADduxFhANYFqCgUpUinvQPqASGitjz8hOv73bAkgXYa
rm5cfLmh53GxBYiVV1LpNVC4IkIAstSZN8s68Ojgs9oHp8onrdSGUjIDkbVxsoFU
rkzmwbvUw6JwlSdKRjyZRvKHkLjO6CTU7FQQfl2CfqhEQCFG10adw6jPTw/IdrRI
KqdgxwvVGpksj6lhnWpMTxMXV/7yE60qRtCzsUEku2vR+6P9Q6ypaPK++rLI+KAA
BQnJJvvT8+FvoOfibZHlC7wwbdQ/PE8mNZraeijSd173galoq6Mz8DF5iL0RNeQo
2KHY60gmqBitwGz3MnHTpZYUQevHGAO1L1Mo82HYtu6N8AxisqjZAzqsFtZzQQoA
q/Jl37dwDieLB6ZXR/G3fN0HD/Bz8NgUEuEP0YTbj80sC0Cdrp5SBW/wJRbET0vp
ILRs+J0T6TJuDusbw+lSWZbxgvUWoumIUbnJGpaOZ3ZcRfZXxyxzq57mftYKltTx
HqQNusGBwQSBI2nf/btk1L73q227QGjFcgGvwHv8GvrZe0n2jt11BqiYweUEd5Yu
/Uqs1GypgvtAl7KeMG1HUT5nSfVUGFrDhQYH4say0XLcUd+4Vezd7bQ3Qt3kjkG8
zH3HZcUPA/V1C37rm4Wsqnec9XrmXBng+u8tKq9h1goA1rBVEP/r0lO5yBN4Lhgr
UXGxwGYwxCUHBLI3TDKOxOpNZW3ZhehSulDXY05RxnC3zh738Sobayf5Gv4klttE
sU7821jVgIHTBJHFsL3ep9nlIj11/8blCTCUcCvEERZxFdQZskfcVYUFZ4bdMusQ
+lAQXkwMsKkWRkvhw0KGxTzS+P25XsNglbcn0Iy8GUuHMscBqNdmE4vVz6Jj1ZI/
EjjCiHttv+2I0Af+KwJgjC+HY5av8lZXBrxaXo31Led9RwQF0NFkmi8mJ2JSp0oH
nkLYAx6gGM4rpVCkz5CqLfNuodNV6T7eb0xbCuxBgIHxF8Rx8zZDccPSZHCWC2OS
MzE3Yi1Y1zemv/O648DCEOHQujURMac8XvUcEX8pVkxDCypgj3qp/xGPqzrAH0Q7
JElVf1RKNs8idyERyQD2RtM1Et0ZYj1tXFQPYxhC0EvluG0brq4WqMwMykts20Ga
l7LDKzpepbPwdiNN2wjQpCJOiRdBKvnfYfONc9iqP57+C9qMTFKdeQIKQTdWZF7A
7qmdw7vLN28fxra0CDZSg02WVDLMzsoWfW4unZGOHpgS/+TC6MU+RQysYMDmwSal
ugA61P5dSpuzYP+mMosUqTCzpKOvHiDlgjHwb1g4RGtpBNloBor+vRYptzMQQrYh
MM1bDKWJpbd4KstexMrDJ1tDQePsPTKQRCD7/LF+nJ73ursNsvOdYqKzHguXw4/d
IMPsoP4QtXMYAXaJ4wiWeRA906GiLJClFFXlexyq857rZj1UVqqmB/y7FbKL9ga+
6ptOvPvTIadYbJkI27TDEx7OjhhB11tVs2FaKsxxr2LxPKknIHGWq4VKn3laz+3X
f3DlsEU8lqGp1Moqp1GQ5ed64BprDUr3rbD6IppLWfTZ/kUj21SCCiH5iaIdH4m1
8fYxgDZIJYHjYV+d6/Hz/Um8QsC7m+OILQGeZj2UIYwKukOm6dOfMARqRnOvV2oX
7rHdl9tzWGoknYvpBLpGlLtK11vWUlHx+Gi1xIVpXv7jSz4U6MnIVKzMTJTWTT2s
ODTKud4T5oq0871KTJ+/XOBwAupUzleoDfdg4cWw39GSfEfnotMmdyXxK6o5stY8
jbED7yAutAa3gR1X3nrzsz1Yd1sLTApFAvTvzox0MHKTJoLvhuurhomQZ7Y872cj
Xalw+Ym4lBzTkBTOAqGhSk4xU4hQ1kHRDyLGsR8rG/epxjsm5prPUOnfg/EjZ+ch
T+efmwYRkYvwni3WwKdOPnJu9dJng1l72z1smR5ojnlOsb3aIjz9Cbr3hat2BQd5
AWFJu1yLZvugnmNq3qKcuiQfwtxKG/e05QZezTQDQtDQ2EFRc0Xc8E5sBAcIQG+9
cChqwpYEA2+0WX+kdibhl7kZaZ604pkgvlppIyHkSdbt99/zZRfF0urjwmiMauU8
2ezLjfLB5uvBK2LJbIBEORAJ0PSB49lWpP6I4ZiH3ov3HEuTBzyXl/XV0+ATrScJ
PdwFD5eSjr94VszQT63El7JKE6ETBt8nKrcOyWMLqYPvBdha69tyV59mKyrL1FY/
NY9vGmQ0XRCcTwxde8Uw/txVhZOPbWoZ1jW4BvCqgBZuCPnLKjmt+aYUl4Pfo0fX
gbjj3C4u+1W1bU4ThtK/3OBxoLhkLhar9OuT66bwtzvW8vRbDh3ouKs63xib213D
2sRWq+VJnJv+VEX6FWsLCIFB/eEqL5QRvIvdcdaEfkxk/RHJV8ugpOb5dyScHCi5
L1r7RGaXGDKOH1bj9ihsvnpTPF4o4Oh6XMCY+eoAQpuE5iIrNNZSYyGegzAEaQYq
rhqChtji/K2XHItUXUNiCZZUzDmTxyNcqlN3pg02mwTWIxG3XJAr3c0kBMmJSKzf
qOHQ2EvwpaF9794X+7UQbexzdGZ46yCHQQ1359TkJXTkms95ZcoaApmIpjvHMxQN
FjaMbPHB+wBeofq0jS3VY/Y60jXXzJLKWs7H4fYBXk9yFcng1mQJC88PrYN17rF5
ysXVMYqdhVGlOA2TIUQtv4O2EXlcSOcY5rIMYC+a2ySwa2lPKxXdu/ZUL+XTsYJt
PeXWBZ+0Phl1HwbEWF+O4i6zeIebK/QX+Z+lCutTVeK6s9VMdY7eg+8Ii9Irz14b
ei18Vq+dTRfuhwxb7Cn7XQMk0Pgi3riDfJ8JNXmP5KVYqwk0AmaDRb8R7svtnd9c
gcD3VeyA/eyNkFXRCjqFAOPZwC6p5hqJvhN3+4pKeGjDjIwXU1XHbDujR+BXTNQB
FzBccEDFYy4UmzFuTP1AC/WHWVBiPo3xVtx5Oj3X/S4Ms9eB/SlPZud4/uMkqUuR
KQx520eJDTkuZ8r0r9ZChOIMcULLaq5TdQ1p/4uYgb4sXJjWo0EJCr7gaIzNTfmS
4OqKLuWz58T5Eh/JbxhPZgxrq5r2h77rcmbHfBGHRcnf1i0ul4ReeUHQvu1m1E6M
E+7nk8gl2cF2CTGx4FaJr7AIg2Yl173GfB7bYxfAY//mgPzBsIZqVvZ48dyqy357
Dmj4TeSd/kR5nx4AAoHgjia9Q6Seq5OAO4IIcZkC2+Kfw6fG+N5SeoR91MfIgJW7
hMEtmUwEVz9cAhbL4BFvMWPpW4v6jTt7rK8x6Pu+9zRwit/js4i5s0/zsMJsPzvL
s3Dq3lFftf7Hpuy+cqqFZ+xKsqwWjwpXafPniqe3VyAozn0TSSLOlF4kWrUukVyO
n01tjHfOHOGuWK6UJKv5tPOYKSBWFLtAhlUfsVrYNSWHuqcCgAmScbdmlAzuaYkz
TFh2pGoU527yIehLkF4oWuDpEGagcdJgd0sKxFFVbkkGNdo0JvcsGZaOWNRHhDUV
nKqfKbRrYnMLm1VeT9vxYvm7seagShnGGUREStqsSskSEcPwIiUXnyygnO9OB73u
EfTiX77J6xiCZBt6U0JHx8IarRDN/Y5o96booDQySrQ8+EaZCzZAffDqJMLim94G
q/TrkVLm2dDrst1bj2HD432345hA60C5qJTdTvWTfbyxDM3hNRtiqPSYVp3BpY2t
m31ekUWmspQgM2P7KMGbykMifn0nR70aEkiDABVEg9AjcuTsiSBIVFGeOudmCqaz
E05Cqifi1djyIbWTTTY2bl3MRpyCKRDPh5hs+2AbhF0f5MLpeEzXRzbpVRYum71Y
sOKTcyudxWcwFazDjXYb1bVEcqEtDHItkKkJciJzg7/ANixGHL4mzPgTZFd/op3+
gqEB/irXQy4PqAI0zFayOegvBIzj1xtM2E4FC94RFYed+qvaFmdYuuA73er3oCmp
VmrB+5mNRBahVFZ7CTB1w9H+pBi+HTdEXVIl/Y08xN9hSw9WKkP0KaNQ4VavVuFJ
GmoVIuFfGuCTw40KnwJFMrucO/d8MbIEuggTPYf5m0shpaM/1XhTpYEfd3LEISRC
kT0qvyXnwAJf6J+TPeLPIhlHoUkP3+Qb1vRwmTgCW7Jr2rINTDtBaBzy/yK83Cbv
BVHZnCRWwQtFmozrS4gchYDYCu6+JZrBI9DlTZ/ow/9vBBoO4jR2xDl7Cxb6oyYG
tW/F0wny30buzJLVIRqGZJjAxNs1A0UL0/rsrgaMxLTgTagrS26baqqiEjjxbf/n
Ux3QNNuIOqQDKen21zrm50QkBJLhhvsfOP16c0Y0FZO/rpeqmX7pMYqEWDD79ZBn
3DI7YCvgrLF1N6/HH6v070Q2AzChb5b5ZdmHRfglEv7oH/W9aXRgcvW396pDmH7M
Vp57rD4dh8Q2ESsvu6d6bYt3Tu7YoGI5ywTfOgNaJSKdxgGvfa9Gkn/A4tORHidk
GeK+/j+PuTsOBZJbukheOu9U1OtNRltqxLJnrNWkkO+UfqnZ0b3hDgys3snuZfWI
xXkjhpRsFPn1HX9wqi+udIIvmnIb4TsrgaeKDLlMbfebKh7eyxdrs8VG9PzSGVVa
Yv422I+KwLXz0Nmm+gM8mhKB4FEUgHDLw8B0t5DYgEcjGBhwwRIWkayLI6RR0E0M
yCev9Cuh10pNWxDvxb9N1199/PuOYXqp/ClJ7ROskgU7l93FIyfMkyYWRqS/EiVE
GLgLR0mxaINaVz6WC+MMIzLDRP/xLQDpBXBIh3rpmSPV1VauGsXgao+bkiorI22M
uYoz61+WyJy/wHF2sLc7EK9h+pvbEs/ZVlR03CPuwiucaFKJnItVtBTR4HF3R3/2
kiPPnfy4Rm21edfoGcNRctqiYbqn8bdVmFwcjnqWlgsUWBmBXaZyQJhmdkLYL58b
moQIIzUPNJryt6P/vZ5+aCFCRabEhjUu5uhDWjkZWNd0om5nHcNFrMUL7bZ9i2Me
1H/YmM2Bh820g8Kj/zwCWJO2OMJx1x6/GSQxs8u0SJU7MfjY2JWBoDG5YACEAKx3
OlU+8AI4GPeMO96jHuyvhdfDVaBJNodH2sVfl1D1KyboSlMA8iFN/+6g7Z7l028j
OH6JayjcnW9d7CYe/vrjMDJJellKiWDTyDx5oR61IxR3MXdr0UR59LNAPsqo/i2h
nhdg6Ft8607cN/uLxV+5HEfCcYLK/b31+xWoB2BBFujw+dpbBSvONOUH68+NNTh6
L4hRJTeVfr5ScID4tdiinBNs1zAirwp99EtY2UPEtgbbW3/ItI0RHFSIZkhle6ZY
mUxVdxQD8/TRTBvA+aTAN7r5TH7O5nZI0Z/vs8Z51dMkJvhLH+tq6L1791EO5Lqq
aj1gb8B6LAzWixKP+a8lvpDYfKkGLqiHmmuJbgol2MRk2RZsbOUghkx5d13xOwMA
5BMNO6PaCySRk8F82MI51UMQ+3lpmgH5qD/rJYMiO34g7BClaMXbfa4AGsQzOzFh
RqV2RwFwKAIuACIytNEjl7z1Ir/g+ATNeOXhDGLvO1ptoakrk134m4+DBD5fdbFB
iKdfWR0S3b1oVl2cbhW0wL/fJy1mzQxNUN5eiVd3lH76/bqr3Ys1ZI38QkbPe/yA
qCbfwaTyZuzeknKEkWnd+OsLMVd49ZvZzQGOH1ZWdrCZ0yu51SGWt4pJNVKO5fZC
GPVg8GvNJe4jtgQ1xqxB4SFhSPnARzAOE5ERZJXHhEZ2x+DRQ7BeWhOSeEGf8zXN
mJYdS5yv/bGad0mi7EEun/0wP40B31QVhy3CHl+1tQwMB7yrIlQ96m2bb9NDwKvb
b5jKBJME/XhZoiEP4tL4Fwjo4S3jJCAT4noUwPrf5cAt+wU09NHRnq4NyyKAyeo+
sEESSKquzl1r8Qib9LIVDKYt6Sm13WmgdOGALQG3yiwuoXRd0BC9mrrcIY8zAGHn
6PskG2oPbvzPnCfMWfOIe/DEx/HBr9DTaiZb5QT6v4T3fa6bFINfRGXugPubaxPy
33p7aCdfqN+4mxgfZh/RsggQ4Oxu0Y8ojCfPnAjU4repKur/7hU01ST3L3u1i0MP
QpvK7JV4bdgSF7aR6CWe7VhkF4ngps/DGO/FA63ufjqCuTIUDLRom2ZjxeMYskjt
slV0YmrOcBKnVA9j1X+aita0AoJ/FGEAAEcAAoV8FC/LIP+zE3f6srEvGYP4Cqxv
EvAXpy69s9kukBjXa4mYGR5aF8SNtziiSWkYhrEO7vUDnNPYE+V8jDza83iVbcuA
VNLQAoV2qBU9Z9H1eb0zAX2C3HGTV9mXLTHxYKCmG/5ZYIWlgzbXb9f6y1FDKEpL
VHgkpry+ne3+0dIeZSI1vCUqB0iK+a2ebQqna2uJRFkVBTG62VVjpr0Sx84RsqYX
yAadaKj1MjhX5sowUmyG1cUs9nP0EZ4PKnrveEQ3J7wuZmMBJW8pcyyxI2uSjENW
KcmIYOXj/IzjA5PV2OC7EXN/UwSDy941rI6o2X+L4ObOQEeHok5koOWkFHAgLIGP
BikVgv+Yz1SK6V3Dfvq6zFpezmlzchj1TlbTwqVeRf5Hasn/ufmDEz6KGSfBsi4/
10irIfAUkyrvz7BC3tVL3dNXHXpA5ULQ/LzkhwaLppMFQSq10ZmwFS8LoaG2R2ep
02uTVtsSS+EtIOs+Y8vWbxmS0bNJk/tyaNL24ZCLMLxdj8fQvgwn4kb6xFmAkkxH
QnYw+czUmML3lYtqj6AZLO81zvzc8xEbMZ5kdm5Y0zBLwHL3Xd5zNPSCSgVK20I4
cMP92Wbovs4kU8k30vW1EH1Id+R3MezHx24M4Mx18sSdsQOS5KpMNW76OydxFcFM
S3dm8BaOtm2F5MZZ/fhKQN5O9Ba3mkWjQ2FguG9/fywSpvt6oKPrPuO+4EPreRGP
HNdQ3xvO+I+BT7VfS8WWNrRbgg3xRPbFPVtLdfuLZ1DnMB87Ixr3wgxctxBepAe7
xfOKIYvBzEeV+PSxbGRblWjP67FVtZUHYy7CjZK+m2H2KTsoreyTWn9vZt/LCDzx
92ujCjfxxVQaycJ+s6icDl8Kpqdpi6EZ9kVV/1Fbu6FuKfNnjj5tLLCjQgebCs/h
xVKv0wbCvBlnIc2l36BtvsKrkoc+SVOFBQWPShKZx0coMpJUJSu8ksLtmys7gKyv
NBVWdawHNu3WZDMmJdprRY0teGtis0i3/P7lxQrr+YPwJ0TeHdXQY2rIR3JdRMYE
xGViEZMCxnNcYuIMiH9OMXlgjh0Pa1CEijJE4aMR09DaEWzjpPB/zpfO3cMC7v9W
BHv5U4UHegEt+DI6YD6l+YDcnXnkYQqVGnPCZQQ9TdGdvcCwtyf7WN6FNFiH+Uiz
BtaSP+bVy2cy6thqoXyemceCEDtvSlapEYrvOyGyYGsnqXDz1jm+8yCqcBLI162O
PbAQDjSmziUYHvnqRP0xLjBrpkTvazCttN1AQ0uUvDxZ6YS+ynNqA+SeBIknQOMB
YnRe5A9hGhd0aU8M++bd0A2+ihGBq9hOKN+aRoEDwM2U98kIprCqSGDAN8/PXaBa
3rk3bZhVfNMrulj9gmXh7MMHbkSw7IdAC7S76KH1XtGZDmYMy3cOcvb3d76leeNo
WsMtLMX3oPJxfEFfLBExZOCL7mQVcZeiFB27snQ66DCVhyYnZT+ENrtMfwu5blsY
Z50LR3cya0fxBlfIunhDkePIfwYwQhNeG67oc4YXJ5RxLZ+9K6u8YLiKe0SOlT9O
gl7HZ8MpmD/MkyuSS1uL1lRdWFp6//5L14TDSY3dgKgYf1zu0kzZVnTe9Ij3WOap
7L0YGIax37c8fzwM1zWhUw4n2vhiUwwjVX3i3DMmTQ+/EwVx5vO2ei5Rd1gQPKkU
hg9aETJzhVWZ04RuAL2OsjSBju5JQQgBfS00olbS0YhT1w9mU4TymhB6l9OMMM1G
kooTXUyCSNpWT4lj9vdw6KaAHZIeMy+QUzs0niPphmTTAt5dtxtAjp2LbAKum7fX
T5Cu2Ce/FHeVPLYSAtjKOybZ6Ko6zKSBGmdGr5oBJbgR5H6hSfng0aSL/QHIwBxW
EGiLYOhW1DyQ7N6c6he6SKba+3V9hauYpaiv6CT2oCwtRW0FDDZI0FXmhkJFaXF8
D5pvlSn+maqI6JMQjWjXE5yX7PUkYTSqJd9n6vWNEuu0upwxl6QtW7LbcreEvyrR
f3XnIa4hcigd3WrgynAaCy4SYkoq/Dcu76ZehYdCdOfNSFH9TgRYmSQ6cfKzMQyk
+2dpTHPgBkAmt41DR5m8wADbJIX8ij6xW99/zl8dmGam4wHmjh6+ZYzq8Es9imKG
ADJ1dhU3rB1onklgNYQeVKgBOgUD+IgLU4FS3a5P5S+Ds0vWhzsrHzT1S5BZBBtC
+GuyoD+xgsls3/PYwlbVI3Wis7b5v8mOnuolnDsLMYnFmpl46rO/R+iYG2T+QE75
`pragma protect end_protected
