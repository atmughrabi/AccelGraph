��/  ����T��4G�v0Pw���-aa�}R�0����H��)c��@�A�yA�R�;�f����U<��|�s˖������`��	�L��b��4$��ȱb�6b�>�arn ���(q�t_����:�}�]:�����w��U�?kA�f@�����!"2d���Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9��ٜ�G����b�+;5]�Ƈ=c�gj20�	�ZP=Q��ձa�BN�6�Z�("�h5_�X�(��`�K����E���!5�	����Lh��:� ��h����b���1AZ��C��v��t�}�L
浴(�¡���}��W%z>�9Ɂ��Z:��`,�v���ܫzژ�9 ��k��e^zRd���.ae�S��B��f�o��"���%7��5D���F%��t�*K��ep����SӈI%H}�{�����{�WO�<��{�Q�O�&�fc4�$�]�OÎP�w���v���#+"ܹA��;�es�����3�}�j�ث�N�C�o�s�C��K���J~�zQ��F�ֶ�lF%c���u����%��X���ǔ>l%/����v�O�ܺ����@y�s��x�H�Vȝ�v����r��(��?�(3��y{B���)�ق�+`��4G�������ej+�C��MTz$ը�hwAB�ek��DtZ�
i�Eh{|L�6qǉ��T��� E�G�@��	����Y����V�$�%_�, ��I�CkW�9D��Cf��z�_����>��&���)p˝y� �:���o�_ﱬX���N��r?J���l���9�P��,���z��� p׏B�!���+e�_U�}~@Eh�����p��ЯuD��M����a�BAK/C���м�n��/�o��9�=<���N^�s�E���?Z� >3�d���rG�'���,s������Һy[f���c�)���:������@'�J_�[.�ȾXm���.Y�C���#:tc3Kj1�d�DR\�;4�����	ӝ�㫓��H�ڐ��8�eAV��9�'(yX��`�J��͇8������dm�D�J�j�������%��Jf���� �y_ ���נ5����6���E���y�4,:�\�q�yh�I����i�17�H ���B�=��ژ��NN�ɠ�������\.D4�슌wB�z�n�;��y���KckD�4�Ω�m�@�6|��ȃ���\�i�����/bT7�9D^R�KY�d��3��9��ok�0* \��E��
�n��@���8PY������j�|
��)���� �����~D)
~��2����Xr��msɺ��cڠz��*`�;%�x����]��>PD�y��v�pLJ��`����G�C��E�Kw���ww�����Jhz��4Z`
�I�r��+���#��U�(�舫;��ڬ� �0�4�҄~�:a�Ŕ�s�5�g
]ɸ�󌏴#�2����y�`�y�ԑ�g7dLB<ղ�Y��{�0t��� �1m�_Un�<ݷ�嘲��"�O��q9w�?A������%�+��(�y��CZ4w���v-��>���3�{d�,d��m5r�Z[`��B�T��n��+��l�^�D�9��i
�.q����SlV���C;�5D�aZM�~��Qp����E:�5'[^u�,��
9����T�z�Ѱg�g�/�ڂ׀ȷ�Bq8R}��yu�ތ��O��t٪}�����%�(�D
���$^����f֞��D
3�Mه�Mp�#9�;���,�D�� �m����7�����+�8? �
���1,;j����.��UL��h�
	\�JNƑʙN�����Ժ�G�*�����E-lE�f�VIq9��Tʟ]Ē����3