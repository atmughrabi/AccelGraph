��/  ��ɇ�[�7�����BV9����eX���i]h����ǊʬZ:�ЁAT�8	��*\��GPq�4k� q�%GT��ٵ�U�7҅Ro�<�?o��)�D>�jQ���2�^�}<[�ngO�]Z�(�<v�h]`[��XG|f.�8��n �2����Ԋ����H����#{@��)	�<�:3eE<�᭮��yJ�Z��X^dݭ5W�!L�cSa�&,�q��zN8�[�cӭ!��K��,#�U�������k�#!�ܼ�jH�i!r��$�ۃ7�g�ۇ�P��J���F��dN�[y��Ov�4�eC"�Sd>S�}���/�;rȅ�d�a�e_�Qx�¹����xc�u��S�@�����w��n��M�֮a�G�����U+�e*���'V�!�}W�j�LRQ�=CpY����<��9UK�V�"��	RL� ���a6�]x�_iX�m��rʙ�'g.E3e�v[��fS�@�	$�%���U=l�\�|���-���h�YL7~)4����x�E��1���L�W�L�>F6�_݈�7�2!�Γ�j#dC���s)!U��tY$t�lE��?7�n(L$�3�iB��6��s���˶-7SOg�ș��,�Q5��Ɲ���#���w�����g8o7���8N�$K~SfdI�k2���dR�p�^=r��T� ���P�)�q�e/*=�^E9����Z(��V]�:[.��7��d �N�<�湵�_k4C�oBG��x ���34����|�����6p�8��ܩT��yW�=	�b� V#�����(�Bk�w6���?�\v!��q�� 0+��y�ØVi��s�}�r�yf�;�������+d�Fu����q�s{���I�O�4w�*�����a��n)B+LQlu�(K�J�
�e�o�ʬƯ�� ��2����v�G��n�fnW�� i�Pw���%�W�
�u��Z�-�m1�x]
��1�.te\�JW�e�i=��%RR���մv� o!�<�CWY�V��ĵ�@)����0J���SM�YǩO�ʢ]O�<�vډ�+eKN^�����د~������ӂ�)�?�J����\x��7�V����X��n��Q�㥻D��8�\GyA=6漼O\W�C�ej9�`$*����$� �/2љ�hsE�J��K����t=yVyQ��ˢ�xo�[I��M1"��/�l`�9��2�a������fc��4
r7>І�Uߎ^r�.�L_��2B�kh6F�@�2��O|Xy�I�UR
}>d�#��UȐ�N�'�8.���-�-oj�(P�B�����vLj1����q�Fc-^���M�(ࠗʛ褝�gYJ���[��fM����#�G<%%#�~:5��1g�\�LQLô"�LsP}'�]�c���%ff]��~�~v��_�M%ʪ�3J�d��i($"����^�	𮠠r\N6<����`� P=t�pǠ��}�p���+���V.�Aah������WOȨL��3?��"�CW�!E��W��o��
�^t�M��˙�ȐOX��	�F�� �g��y9կ�p����#�.����6��x^���OE	2�m�n�EӸ��]�\�BP�S�K\�>����FZ<MP��gb!��z�V�W�ĸI?���x��~� ���=�A}@
:1d<z#<�6���S���W?��u��[�c���5貊5U%hL��8M9�#;�x�]��?�"��Ƒ螆���H���XQ��[G[x8��(}�w�W�"�x�Zz�Ł�F̝�M����P���5�����g�i&~`v�����qO{e�MTT��Eq�!i��}[�I"�qC<\$0��n���'kp�ɬ�_�;��0!o����-�JJu��{k��ό�Up�6�xŖ�5��m��N�'@J�pS&��/0������w�L����\[(!bȌw2�#�[+�����Jn��S6D �	�K�*���C�l��B�/�Ӏ�d#A��D
����$E��\�7��5
�v9�rm-��j.�4Z�o��5?<�Tsv�c<��+O����t��RH���t��ȅ߄�I�Z�мp�T0�D�����%G̝k���:i'��{��P��L�7��`�B���C���
a����ImM�f�*��[r��h�nF�:WF���$~�(���8CX�:��B7X�:�7A.n9�D+�!4��^�9���?�w���՛3B.o�M����&�ɪϥ�_��/�C�AqD�b^������	�7$��o�R�]i@�4"�,�O��+�������%j,+��	>
�	ɕ\�X���m�fo�˺L���A`��u��Loz����l1�K@��D��Z�'q̝���VY��`��b0S�͸ 1��̙�k��=@&��9��n���"����x���U��'��Yh8�|�	A�oc�B�)9��Q�|c2$�$�.�yBƑ:{н�+=�q�)�7Ra	�_���<�m��tc���51ڕ>zX�s'$P���ޒ~���P��HN�
o�EuY�4bJ��X冪��;�9~Hr�]z�^@�0�B)t���
��(�_���nhê���L���Ư!�,%��	�<�$��-�5M8Hh(�F���{P�r2¸�����>g/�r[�w|O�����ai	xz���O�x�d���8n�S�h�fP�m���D|�wg�����}3��P�I�7��(֐/:�q�r�	l���:Y��a��F�өp�ԧ�WE�~��ํpHy&�^��gi��_���O�t�t�C1*�}-���9miݽ��/�� V'�d����������M�DA� ���yG��nŖkY��#�|�[Q�"*2�v��*��2�`{�y�?��hUC����d��Q���̫�.�`d�;$t����?/ޑ�H��G��eҺ�wp���pm���IK�v
^s����SK��#\�^m�g���'H�m���[V]�@��7�?�1�K�`/ɤv������c�Z[�GT�2���SK�˟�w�~ll�)ۆ]1!��o#�&;� ���ː�L8���n�e���9��	�awԫe��}Pc�5��6g�G_5y��K��ۭÅh~˚�Q}o��9I&N�>��Kq��Q|���2��q�����d�Cp�H�N�:���4�����쐣���S�-�:кՂ�^Ӌ�x��LJ� ���T�Z~)����Ne��/�$��v9Zo����1���=!]�7����c��H+R֊�������vB(���TQJ.?d�*�Qb��7����G4�����f-����~_!��c_�`nE�9�;7Σ�dr�����l"�i4H������+RQ򸌿�Ђy3 ��;m���o�G��<�36<i�(�հ:Q��ܐ����b92��E����,4-=�8ϸ��W�
�a	�*;X�� !�&�]�������xd�1iG�*1�K󵹆'5�a&!A%wͭn|s��A�J�ذ#Ѹs��г�~��5u�d�e��mDޏ�� Q�D�#.��:����I�n����['	ٮ���.�+�I{���X*f�S�P,��B��L�Q����ڌ������Bd�.tMd�39q�mt�~կzUu�����&f�p&�sB^v�F;�W5v��a%OG��~κ������j�PEb^a�>w'=*^��m�Ē����t���o4���ϪM�}eػ	�/d-�R��d���J-B�=5��ԸVt�`�t
W>��K��i�E�'9u����ǝ�&��y�)U��k1�O-����r�١�2�-���s_��K�{�ۿ�˻�%bK&K�,#�^GA7�s��F#�X�ʯ ��4��!�y�o��hen(Tk'���g������{��hb��y������8ņ��|�� ���d}ŰE���di�b�q��V����g�S2m�7�L�`�iVNvX�Y�GT��
~{t��Ƴ+���"�����$2�
�Ŧ�&�˻d�(q������Wz�57���sn���s�"f�i(�3�����P�o��9��wO�"p�M_ 19�~��%��G]U���T���-S���}���,q�:��w���\s�1�6"{�k������u�o�[�Mc>�~ɓd�I�fnx|*G����WV��Kv��3��ѭ�t[�6��u��&�m�n����
/	�]��%<>�7L*��X�*�P�Ws�:��wG��(����5�{��De�R����,��8��^e�'�'��KH&�v�}N�ލ=u羲DlcN���Ŏ�N?o�+�\y�Ŋ= ���T^>^� [dM�t��{��l�����$��ZY�',C�*�P�9����z��Z��Ժ�ݎSn��.��8�>�&/H�/�1�͟��C���'���$/9s�G$����߄'?C`Xw���X����o-{2��D5� �6���r�K��҉����j��¬!�L�C��RA�p�2��v�G�q�,Ò��u�o�r�LB��1_?��Q�%��b���,�DA|	xԼ��']������/|�Báԛ��<��.Ѐ1_L���\lm�&��&H�&'�m�4�VE���x~&m��'�g3���p�_�w~��f����B`�CFU�T��x�<Qhݱ��2!��e���԰H4݊ؒ��A�!���P�q#u�O$�1hL��m��L���m���@">�
���V�����Jb\�fH�i��v�`x#��4���`��:d�:���Z���\'S�KSҝKl$h�,���q�vU#{ <��ԁ��+	��y&-����&�F_.�e�(��ze��:����{�+"�ߞ��zLm&i!o�R�,���S�˛,��5�:�s�ͤ�r����gGf[۹Y��Q����3}��X�m�o�g�_r�W���I�)�,�Q�#�p�e�%�F����Lƫ��`�'�fN{�m��ܛr�(֗U�yC�դeC���g�2xg����$�-f	s�~��ne��Ni�1��f������	&���q�l������a9�,�I��XIL�n�wx��?�r����ͻCV���EԶK���˪��4M�Z����$!ֆ$��֐0'�y�{�{�dCF-����)���_��Ӽ�������\�в����F&�$�rv��:s��e����HN��������J���h"(x����/kū,�0Xۦ�r�I/R��6R��So����$>�"�)�J�����ʼu���E�O��O��4q�2-���ũ[N���f�T��Z�,���G�]r�b���1M:�/�!���OR���>`�����J�٣麇ɽ�U�>�_���� .{�fSm��3��`�Z/Z��,��?=I�`�؍�C��M�ƙΏ�$��~׀�8��:��nrvk1��	�f|Ix�e��>:�-{u~i*Z�ZB-SXQp֟F����y���A�=�m^�=;��T�փ�\h�Ǵx���o�>4g�+�R�N������f���V҉��!W,ҬG���`�<�JFK�����fEy�Z�\b�v�	��(� �i#�v=ą��x�l�s!u�8W�\ � �����2��h>ϡ2�%�/�ݨ�u�#�p5�xT����ڲ�s�W���,��l��n�����}�?ɗ�93
�J��١�6�s61S���*�j��U�wh�]��k ��쮎���s�_�p�	�z
����>�:��;�ʤS!/E��۰ R�9e��4YL�tK��yp���c�wg��oaM������ò�ߣ��Gǔ%f���+��	A ��|�Ą
?E9c�_Js�g��oV�}���H���~��>r������1t7r��F��7��G���L��:����)��djqS�*2��e���m�aWf_:��v�&���zҀ��w�}˿7���Y���?��J6�z���_	9UK4��cqX���)s�Հs�}#����Z��s�L�%8�h�`��>H�\��U>�l��_�G�{��g�:X�,�o�#�3VH�o�wtN�BF�ħ��r^��&���>m����Y��㠔#��g` p�I�o>e2���
�^��9�A��P|{'d�m�+Sw�dF6p�͘G�IKC\��:��)�m �^r��6�!�;�ݒ�gݚ���-�I0Pmҧ�A����3Q�i�4�vOl���9�c�!��_�W���닆���%�E��i�
0��FV���V4�'�Tf�S�ŉ^<���L%o�������a<��| �
�{�l�C�A|�����$X���M?���Ef� ���֭7G��1�#c���>�ݏ��/�J�����&�|]��q���@Z���Ԋ�#��ᯏ��A~ޭ��.)q�{"ϐ֎����x����ٍ��Y�e<�)u��;*��psj�)˓j�	,y�B�Bq�����^gy\N�Ōv���S�pщ�42�[���^�O�~S|Z��$� 4O�L���7
�L��j�|�BsYS3���2���iӅ[RPe |��.�#J�JsȜ\Hh� ����C?S�n����-6K����h����� 걐UIk��ۿ�4|�7�s��Q�(	��L*���f'��i�;9^r�OH�T��g)G�8fY�F Jq�S�Xa��������"�����V~v\	>|7�>W%�38r!FXXV�����<�?����)xQ򘥉�>�����c|��/9��[Q�{3s{�ǥyTd��@��a��£��|��l� ����0̭;'�W�z9@`1� �B����&�0W12ē�ZZXUM� �y��Nb}��ƢPFl�����x�3���� M��/�EE��!�1IQ���� ��C�SNT����oX������3�JO6lm|}8�����=g�2_???��</�i�<��W-T��g�����+i
2����o����3{���9jk&&��~<|t�E��c�QǾ�F��ﯮR��繆���9'Lq(��f6kJب7V }���Y@o6Zm�Ny��8�7��"~e(ykeh_�Ed�\��01�hҫ0�@T�6��e��6��H�i��j�4��n�O��:����d��U%�$)�[��ZrM�J.2�5��e�����2�61qJ�Y�?M7��OʜL[��$C�?���Ŀ��N8G��3|I�\�ʖ����,��{�k	u'"N�k�.:�Up��*̈����Oj�$ �g[�J����%^鏾{�4��W����Z�o���U��B�c<��X��6�Ƭ��
� ��J�]��%{S�'W�s����%\ڹ�<���k)9�,Wb��:U��Bmc9~�I��i�&b����˩��$ �7�Iݚ�?�7�cz3�TU��[�DYui1�F��HV�f��)/���[
ޭ��O|�X'C�GA�������GN������W���Q����s� #��rW}�~2�A/��L�_!��y�M� ���|x7oKU�T�Z<�������:���כ��,��M`^��"�R�D���]/�e�b�U�(�Z�R��2<����8���z�C�`e����J%P~O�k�구z�x%�,eN�6�_@m��:�@�Lɿ��s��e���y�	֋�x�q;�Jjm%v8e.�	~�8��y�����_v��
����Μw*"��%���,�4b�^1	6v����U�'��	�)��@j�n�$(�aE��	"y��џ}�}62pLi6�������<�3	��pzZm��n̘ ���C�DL�t?b.7�i��5J{�v�-��q��ᒤ7k�nĽ��v�l�f�:�'�W��Y�������fz����hS�X3��s5H���"rc�ԙݔEEe��i2G�*!�\����ڥ_7/�?&�q�<讀��B�͔�gy��|�4�Jw�@d}].^���M٤×�<3�$��2��@NFl�y�ᳫxPW�	�T�
;��B��|���P�tcN�?�<|3yǹ(���I��fI�7�5���I΅�eں���Z�F|��lZ� ʝ`��F̚5��R@nfӋM�+�LR��5Tb�����**:�C�p��P�U�?��T|`��5���ӳ�@x�%Y�q��I%{3�sF��MyY�
b3$tJ������"O=\���1F�?c�%�u�R�hO�0�# 	+ի���E+��S���A�u����IH}@�2�S�x�����,[Ip0o�┨߻��o�-�_Ӻ�iV �SR}��;�pX4���n��@6���{k�NяNy̪$�o��RUŔ{}��*�Ӻ��@�yz~[I�8�Ud�% ����S��i��/��׈I*�쐸�
 	���)W�i�N8�O�.�4�:[��*ǝ���Bq8�p�@3{ܸ�#�Z��S�~g���Ne�䙮�2�R�JQ�ǆ�V�y��,�?L�7�XG��� ���aJ���V�@(!�&�Rk�C�x��M\KqK����t��o%��UE���`9D ��P����Y��V�^����=��+Q����y)�~*$Z<D���a`��� ��:�o�;�t��D�^q��Z����J�rW�X�j+�% ��<(3����	�5!3́��k��V�z��M���d�N�5oF��r%_����4���EL=�Q��SƁ�I$G�@���Ǧ	˒4��3�ηʏ�)�u5]o�|�cׁ֬�m��i�`�yJ�ǣ�J�%��*��'Ͽ��6l�����%Б�I��'�v�ս%/�S��o�Xk:A���Xܸ�r�S!�Mz��͟�O<&��Nd��Vy+��D�	�(A�Vk�`�Y� RѸoQ ��x��ݚ��kZ�?�]�D�6����	A�5dD��%~uO\7gn�砦K]���#^��#'D���.��lb��ֱ�f[y[��q��I���7u�染�5.��(2v��)U@Sj�����jt�hnQ�~�m�i'숻v�.�������mX�X˸e�4.���/�񫗁h7���5l��<O���!�d�����VU���W��ɶ�F����FH4��K9ن�x�~.�E���w��O�(85��x��f�ji����| ��Z冺a�[������C�$�[15�G��*e�{cMtd��W�cB�Q5�z?�Ep��pݒ� ���,���ۧ�;�.�?�m<ۨ0]�o7���C����Ɗ�u����6�����Lxj!���t��PMj�W���y�1��ZТA�H\�� brq/?-X[N\�n�]���@3�<���T}��pÏc\X$���u��.���! p� Q���xC�3o�5�^�hzb2����;�����$�v��k�*&�{AlNKB��W�$C���y+���\R�<�����r�qFX@�����	H���hQj�K@�KA��<j��f��|��V2i�E�q�$ �P]���>�U��|��&aW~�ϵIm/w(
3���<���p�`�)$���?�	"y�Ԛ�x5�9&0�m�;������ d�ܺ6�5��2�y
2��pپc��RrM��+|	�ަ��L�MS���v-��z
vJ]$dY3���Xo��C+/����[�'��Z�x$���
%���ǒg���Y8\X��Y�F���'ϝyq]����*j��;_w�OQ Je��F&���щ�����x�[���� �<��4"�J�A8�������!R>9}��A��/���nF^��2E��Y�i�ְy*e�Y�+���DB��{��~LwGN�������V���PVR����`��3Z�yԪ�20'�Vk��dgG�{�^�u���9��C��o6x�?�?�O,j��e���;��i�r�2$v���SF#)�F\_��5^��+��<����3��D�R��悥nn�5L�ƀx�u�ʸ�K�6n���k��=`I=]#�@!�9b�Çϛj�e�ޔ��5����Ex�ӡEJ0r�0��y��=�E�'7�V%)�*]n}�PA9�''Fqp?CR0��5ն��ٻ(�/ �n�po��IJ�ze���ܪ����bIE�<c��7WL ��aBѾ��Ӵ5e�݂�l\��7�o_|g�1af��{/��������9�r�YRl�I�3P�a���}�Tf��w���*ȅ�$�Ñ��?S�3R���q���D��o���<iG�Յq�X|~7��¼Qy�!�I�����Y'>�R��U�����|j�eeU�:@h�@0)|��6�ĺb�{Gz�����O��QABg��gA@���D�B��R�Pz7�?md[����}��ȏ�o٪n�*ɉp��'/)��:�d����ߞ��?E�*dς���T���Oy.wY6E���u�=���(S͖���b	cZ%NV��w-�h�\���D)��t���~��YS,�
\
w�(����B�j#~�����2a�+���Xny��'���޿�#׭�wJ�RX�O���-��e{�b�u+_g����ZC>_��_#�w��$���7*�}Rգ񄶗�v=6�|�ƭ!e%i�Q%��ddp�UW횻�8�$䡸�E�#Κ=�"�@�*@����E�Mя��H߁�W6��7I�UjBNh���3��ȗ�y����D�Y"�'w*UV�!k��:�,V�S&��9�Jv>"�JaM�j]��1�3�5dU�l0���(��/b�8D$��!��2�gO�8l��{�^yA�k?�V��a��K�N���#^��oahn8�K��B!y�s���� i쑒χ%�5�~�ae�C��Ma��¸��l�5,���}!Wj��b���������H�!��I��|���{�`"���e�LG!b���EY�������� !��lSf�?�;K,1=#�+��Nh�r��s8��$�����!)�*�"%�D���� �1ώ�*&	H��5v[�'L)�iSy�������Ya�\��u�R:�����؟�g��M�u�f���@�0%�(�%�Av����qs����4�ȭZi�s��������[�+��ay
%\A�՝}�
�JK���2b�(�u�4b��y#�n��T�q��_�$�o�䙀&]Ts�-i���]Rr�/�@+�
x��*�޽�M{F��t.�cR�2{����}rbw�~�!U����{R�%�D��aL��U�&��0�nBhխ��}�]�3i���y�����-*p�q`S�i����X�T�mA/Q�z9u�����Aؗ2����4l�U�U�^�M����<=�*�'������4�^@��#�Ac(��gphA�����Z�P,M,iV�c�r#I�U�pŚ��a2�Q�������*JQ��8�/�T�W�'Q�EP��"�����KS��\� ۴��t:H}�#�H��(�vo�fC'E�N�殶 ��UW��gU��� �"f$ND�5��Oy����	�^���} ��H���i���k�f� ���q{U�Č������p�0,���!�NB/ʘW� z�$F���IQ��L�6�>�nv �Gc�0sw���3��ɵ3=�c�惋�(쫇���T�l������>O�\�(q�Q�%���mxi�&+-�-埛��c��o��qC���ڦwE�D�#���ǡ��?��7�	!����R��b5��&�#���(��Tw���>�Q��#-��ޫ�_�h��� u���V�b��U!�e�5�3y���Ä�����Y�c�5����갑�#�\2xq�w�`�l�×�Ɏz�wU��U����+�߽N�W}�#��Π�։�:1��Z/_L�����~1 ��	�`D v�m����0]�mx�	j�$�휁�������)�)��3��Ѷ>���Y�H^�D�n��l�w�-Ht�09 ���3��Sp�%��U.+x�f�]*iVގ����w��*�.�n�?��mW�m�d�� c+�w�+���z������`��x���ҋHOՔ)��o���W��F��$�Eg�}�#��`�u*�y&ў�=
0X�b;779Q��2���,q}��� �'C-�_u�G�"C��Pb��Ѐ�g5oi����|>��� ��K'%��e#W�{˩�cmz~R5������ F֍���@y�1�A�)֓_�NNa����Ĝ](�g3i`�����R�k����P�p��E����i���(�;4$�7�%0߰��������B���^5����P��z�r�i�8G�dQ5� Y6X�*m�H�鄡@�qi��81�f��\��M��ާʦ��J��g#�_hΈ�̌�T����5��DďP��t�&��V����	t��T��kVx-o��i##����=)������p��^��^(Q����p���P�Q�M�Cv�;�8�x	��ż�L�
)��3q���ȧ�`C�i������/��1E�D�b����K^x6;�S�?ҙP���z�F�~o�}
����&eN��Rf�î� ߏ_ϒ�yܯ7v&4	A�=��=�S�ȹ~U�(�2]�C���?��m�*��ӊb
��0S)/���}.G�>��ķ:F�X������
�͕;Ċ��ۘ�d��v(��K(o�h9[]!�pT�������Y�-�8V��ŨϞ����Ņ��8^ښ.*q��x���B�����Z@�xFlJS֨&�|)bR$�1��"f9Ur#C�gIy���K/2���8�44l���dDH��jvY?�[�p�~&�E��>�E��i�x����4��(O( �ro���"�� &f߽��7n�1�#<g"� |��jk^L���l�,(�q������/����f�|�_D4ؾC9pip���|U��l���q6| ȨB������߭ReZM�'��u��A����-aa�^�<�9_ߴ������Ą��+�g|�}qE��d�/n�m0|���<2�����w�f�j�C���
�p�b2j`�����C҉ce�ՙ�ʝI��$^�Z�����ێEL�tELP'��6QHg�E/�,�OI#{	y��۫��r �j8�Ͼ�b����H[��a���83j@0,}T�����&涧�C�j��:�����."�u"|�hf�]v��D_�������wG$Č�jd'q��טdj$�"ܢ c>�����ء�a�rKEҶVٙ�2I�# â<(q��D,��lC>jSa���C�"q�9-��c��h��0
=	�Â�J��4(��g�|GF�V_B+�"�p���tu��v^��=P>��r�S��5N�v�؀Ш�G�Mk��W����r���!��&��}��`a�����:_��]�܃F���a�K�o�o1�X{��Ԕ6�܀�M��������y��B����1�XDx'+��r��V�jWc��:Jʆf�Nin�.D�'���Y'Zq���{o=� =E�G�C�ex��Z	J�T?H�c���+Y��[�f���Q+y��2���x�ɛЙ�{��j�&�3��0�=�y�6�F�W��>+�d�D)\)��V�x3C���(V�@Su��"B�_��-;��/��lr>�7�z�L�7n�o�8#���pnV�D&RD?Ԋ)6\��Eߴ���< ~G$���c�mJ�^v�x�����$�Gp�e &��|�t��.�Db��[*;+�A�:���C�<��OE~���DqJ�R��D7������,(ꊦ������ZB�Y\�Ξ\��Z�(����ܹrPǗ�y�����1���y�Nږ�4O)c0F��R���{����aE�c#��Y����%�,��JP�ʁ�y��G#���oOÌ���	��O�J�L��V{�@XK�yֱ��a�t�c��FT�����1�8��j��|���geǩ^K`(��ӯ0�$G�b��U~������>M�v(��Eŏ�e�DM9\�W��ͧ5aye�����/JR�V�*Opgǚ���&�^]}z����
��R<�6�~�*�z���ka[ɫ���AK�����;~���
��V\BqN14s���4�[�T�˽���J7�Q��Sۑ6<��W1�$�ƭ��Ļ'��bNi�<x�k�-HL���g%�2_�(�4� �^RW)��u!�:Gk�|�J=��I}>�I��t�� ����ǰ76#�ў��,Tj�G�ϝ�d�1�i!�/,�5���l,�xVN���`��;I�����(U����m����M	���~�73�U������,^����V��K�m�{i�{����pS9[�g��{p!�?�S��������~#��Pi��	8F�-#��5��t��<��4�))�E���4�6�^��qy������R‣�n�>հ�,.�q�cN�]�/Y�R��܉w���R�	��<[��ҧ;K�E�,sD���,��<�_�ڮ %����-ZI?��Z�Śx��AB|f:
�z�ն��ps����7� WČ�:x����ĹM&�g5zdI!����z�~�,ptLQ��n>c�^}]�AZ�ׄꚣr�����6ܞ��B3�T��4)}���!�E?��T�^�w�9ʅ���~�EiD�~���~�-5H��y������(��#��Yݽ����S{��&�r�yKBN�T�C��.����g���0UB��	t�Pd�M�u�o�j�#g�ҊȄ[�bd�޶
d����75�mh��'q��g}�6�
�2����׭��;L�k��i;BSI%o�����F�_-skM"�2���v�����:���\K ��&t�A�e~l49�g��	U8�򩁏�(%�݉@0�j	җ1��ͭ)PߗW��\>= �1��^}��n]��"2%vN�c�%t1��vSIV�ݬ�1y_E�]��?Vᰂ �o����Xo!�~��؅��u�d�E��Cs�Y��w��r:ky\�gDN%u�j�`@��[��sf�[��j�@�P[4Xfđe�DT�ҥ�����0�����_�3f���[�h�O�fY��V��e.j3�a��	�ɒy�x|j���'���D�[����p4��r�"�UY�gs{�j`y��]\����.�����ݸ��;�m�;�O��Wx�0C������緔���6F������A8G��G�2���:�>����
�0[Y7%I�tm���o/�7�q�`闻�S�|߶�x9K�g
���v/���M�|�?�v�`�%�ڝ�8q{O�h<���v��1[m�{4�NW��j �>׷�_c�'�u�O;��¾�^�� D�`p��|a<Z:оe�l��\�Ojr�>�U��b\{R��DE�
�tD�H����>����v42d7!���g઼v,*����B@9��x�L��A����뵈���Z�Q�np����h̔`�d���(t�\	�P� �%7�./n���)�6u�����&�į4H"c�d�q��ݡ�Z��"F��>r#��������B�;{v�
�NCԮ��B�y�T�HD��(��Ho^8/�7���&�^"������=3j�z�G�V
H&Dn8{Yχ��~��yD賽_���KvMe0`���!E����R�1�sƘPK�$N(�J���n#�K��b������v�^L�X&v�Û5I��nLi#򢻙��gBt�P��Ά�*?��H�o;�"�zP�j`��&;��cV�|]N߯�hL㿤�����s��l�Ԃ�c�Wj�93����m��ڮ>d|�w������F�r�=]/f�����9H�"�CB�&fG���	�����2����?��z��L+�<`�Ur^�D�> :[�0��y�h��'7w]�C����!�� P����+of9oo��=_����O&e��Y~j�V	b��M�E�@k�(%nn8j�����%�� �8`�E��:�Kr_c�^+?m�xĜ_�#�S�s�1,E��|::���"�"�?�w<V3�*���&ɴ��n�����0<R�K:+)���:��_KR���|�r@9G�~��,Y�fy@���]����ZP&��@��e������X	b�j��Z%�f��Ɯ�p��s�3^c���_GY�b7��F��ڻ^���ݸe9�����*`�Vc�� �{�^u�FF��'�A���q6�c� ��OQ��l5�k�dٽ�v�2&�z�U��2h���#��>����xԂ��6c�et��"����<��gL{M ��#���L�"���14K�0����k���)���Gl�����Ӗ�bS�%����妖b�@V#;��Ol��.훿��g�&���u,ݓ�� c�1˛�0���c�z�ӱ8��M\�Kt��6���O���s�z�w:�8R�o�ҫ�����l�9�C��t!�L��I{�Н7�:�0����Ji_�_^6-��w~�|��<��ܠ ߒ��Zj1n/�C���qh�}�Y�*�Vλt0Ì%���gY��ӯ� �����c Jp$��3�W+�K\�oï2[�=*�Z�z -8o�� ,�{�`̣���# ���1 �Kʪc]��C��c�xCC��E��0rtw�>��M�v�}�ft���""���n�v��q`�}#��I!z�M��̝� d�Zd�Zj��B�j�U9R�����r���z�6a��}-=z}ܾx��������п�`�{�����\��Zjg>�Zj�^`�|\�o�����;�
iv@����j�5XsV��i�X��D4����u�RW1n9R��K������\V��P��!1DD� ��f��	F�v4�B�����E8�H��2G��p�)���eƌ����z�E�� ��I5�M���Oߗg�t���^B��W�--E�!,�v���i�a��۹{��ZP��&2��/+�A�36.5E��ԚI]�| i+t�<�����?��H�\G�&c�q�qJ���W�W��]?���32J�b��ُ#	8+�ů㥺������f�q�?[�!��gP�qrG�<�w�N�I[S	�9���ŏ�B����"`6� �o����OK�_�I�l~u�f�!j�fi�h�k|��b]��hw-)Z#�Ja�����b֍�K�.�[ڑ�܉�:&�5��#�v��F����^�3��@1+�\ed�fv���+�N��6�]�A�&O�~�B�n��D���_������w��/�_H�B��w���о$}��s`F��s�Di#	>XB���.��;�vvj'�huy�6��T���q#�T�{��?� ��y_�f�0���^�Q�y,��Mʠ�f�a5�.9wuA8�g�w�MF��ⵟ昿͎��I��l�g�����Q�udw�����g��
sL��X?(���g+��X��e����i�&rZd͌�~=#�o��e�#D����P,_'\&aewF��Ï�0�W��73�֖QlHg����vp{ҷ`���f��xD�����o�*xX;�#�%,�y��1���,�je���BXb?xe�|�g,;B�{���B���9J����g'����֟��2R�mz��
Pٝ��*�����y�ԣs�u�:��Tg"���R�!����,284�\��.O �l�w��l���!�y���X����� M��w��T���דc�w��7�؈f>�w��U�1���W�~�K�l[Q��<�Ѵ�%�^��5����1��Q�<=q'�wc�5>|2��� ��C K��I7d�1'��2}
YUm�Tl\��>��p�̓T���\\E�2�Y�%�����RL�X�|�6���h�����:\��jjq�B��kF��g�׎&�E%Vj�����a:�* �(�h��������:w�dv4�T=��Q��<�Th������bn�o�!���Xa��w
6'�Fw$!r�z������$��f��+��&�JO�Ӧ3�I��Բfp�w���9"aVq�`<FO|'L��Y�A���0}�$��.���ҹ���@��Z��^��Jn�XvV]{:��5�t���CN'Id���T����Rh�8d�ѿ�''Hy~���2��3�kp��J's�k�^f�'7k�u�}�������1�h=�o`��� �A:
�B��P�t>�<��U~�	^�H��¯2_�r�����s��,��sw�Rg�U��ٙݛ��KT��+�#��0���Rx� ~��j�|xV���馂 zc��dDM�"~Ʀ��1�J!
��)�6�,���N&XkB�e��U�~�.Ym�^91/����.�_���[���7k�
z����w`�w�;�6f;h>���S���+�}���?MJ
�d�Fq�ϟ����O���A{p���YP�������pG�C�!i�&-�E��1 ��X�Y����E�f�}gsâ���^��w����|�(L�N_�x�J����D�]�㯳��\k@W?� ��"�5뇯�a��k-t;���ŕL/�э�	��.mPj���9G՟ �T�4�/&�|��!��b.��T,�+;͋�������Tt���$:�q$�c�s���üvAZ�Ya����,�����F�M�9
���oYm���s�h�&��'��~#���l�Ev�?붌z51�b6�2�(�����vk`�
1�]��&g���x��Zc�)�K_�l࢟��Zy���3�$K��Y�S�өR���P"��6�`_R�H�؈�asU���->ŐHy&~��Û�y7����,�Y� ����sr�p�E���K4;�z�^��ݥ#�-l�݂�/f}�:�9�4��� �^և��pX��QY�����ƾlQݸ��Ɉ�� �㉆��e���i=�`��ਾk�*���^qh�Y}�u��thѢ��Y>K�<�7��_���@�y�P��X^G���L.;�tױf}�G(7��<���k�f�� j�9g<*0�m�&d�c��M�FǼ0�#X*�)��h��)��5�,��4^`�a_v�;q~M_������}�QpOy��:�	�0��#6�3�&A>r�`��`s����Vǡ�%չDVԄհ�)=ڧ���H�}}$�����B��V�O��*�P1��Z�>�����~��bgk�/ҽ�<^��M�=�Y�- d���$A�:2���(�>��8&��S��r��VW(��a'-0ο� �ϝ�f�Lҳ�	 YZC�f�G_��QvJ����Kн�N��
TEς� {�ɯ�v�qwL���ܟ>���AT-K
j>:��MH�����cr�_
��ȴ��-��Ǭ�K7�F
p�� 8$	��\�H�,5�A �]s7�� ��Zo���B%o����-�#B�ƣ>�~���0ef��"R�ZRIYL)gu�g�B����s�!
Q�:"x��wl1��E�k��!��c��j�q��G25�/�A%�Bc�4-q���%q���-y�����=�q�?��%���^�A��l�=�Z_t�0��m��?D�)�1a�VL�G5�&[mˆ��d"��#+�^>��or��b�? w�����p��$��{X+�.Dt�e�Nu�k{�}^.숮u����qY�=�MG�	TX�a��$�K�����	�D�a�&��hSh<����<~����J8�>�@0,���j9L>����{L�<fͯtӤD�^�km��*���&?�8���4�0���0��&���ӵ�%ܔVdo]��]�ʇ}=2`���ޗ�t���ȉ&���A�EP'R1�r�6/tZ»�l�3 �g�n6�'s����ۚ+LǠd��;�ʞ�e��=��%{V���9�]�-�D��_�/`ԁ>��Ʈ6��Oy��{��X#�>d�Xs���$3�Ro7���n*m��L�L�1-���*��c"긱[�������J�-8Xmz����=�;���^/]�;�ʘ��,���cױ��0
�ui	�Bᇎ��ߒE��i/�s<��px����7��!�kmCD����ɡ2̸gF
������?�@�t���.���T��!�(��J�����H�SC7�5�oj)���w���]�e��`%�w93�^=��Y]M�~`X374���n)�T�:FW��@k����]��ߠ���滪N��HGj�@ !���&E�4��3��s�$�"�^�2��3�&li����*�R~���V�+�r��v���ן�2Tl�t��VL ������ڤF����kڔ��T�I���D�օZ�Mjb�2���B|�K�Y��G����$'w��:	����+��������	��g�w'̒�UiO����Ԛ������9`ʐ��{o�6�@�/���ٓ��q���CRo�E�t���W1R��p@��s� w}���0ԉ4�<�)����G �˘�*�
i{F�T%���۲��e�'?����W���/�d����������t~Fq�W�߽��7*�6����Y�	�3�
�ps��de_��>I����� U3(�}/T�R�GZ]T�@���;ss����^^be�Z�8��L2ջ�%��pz��TErE��{l�;�xL���-�̰�vݢ$�)�m����[�A[9��O��S�1�=AR��Ahr�c<��Å�Հ���)������f����{Q�g�g��=�S���|=��] G��F��<���&U?I��p�7�)Rٿ�J��OA8�(�ծ%K�v���8`0�Љ�F�3t�)�o�R�C��@Ѧ5�����In�ek����.�_��X%۲�H�æ��7:~����&�B�P��w�6!.hy(�P+7B��谥.��.�ߪ�g�O�������9�.�+���| j7������l5�Y��o�f��^��eM~�
��>-[�����9��q��q겪�Ғ��-�v1��p6m�|%��`^M�$A���D5O3%�"�w;]>��;sv���M�ŗ2L������g�i	4 �&�N�%��f�Э,���z�[W1E�A,��n�����-�~T�e;ı�`�2}X��\�H�r�a��HM�/���(FkzӠ=Z�V0�޴��S�u'�Nt�~�)3(I2߅j�V�|��gK���P��Fc}8J� ���8��4�"�A��*���*N�j�_��IEaZ9��4����I���?�s�q��׀���Ɛ#](1s�@P�Wp9�BVH��4}<�E��@U.(��u�k�����t2��_��=�m�Hs�����<6d��N��-#��ؽ��+1�C�˘ڜ��Ej����5��Rֽ��M;�K�b�xc�;�~H�c���
��.��YV�q��f�� JQ�>#��Y}�7�26M��(f�e�)����Ԙ�VYd ���Y.�6�kE�r��ج^����'Ǐ�Arm@<���'SOyJ͛��z��x��U��K�n>���1w;F����$;٣2`�u�/$���,G��E�£f��	��Q`Š�5�J|��O��G�K㪿��)>���I�-]�����7p���f��5(���p\o$�~����ZFo�d�z�uyd3�����7�m��#��n���h�3�Db|<z#�+�*PI�U,K�}�#�]:;{C��hߟ�c�aq,��K. �5����l��i8��"�sI+��?��<���]l6��L�n�P_\���C�3�?c�ʁ,���$��	����x���� <���%�]��G3��3�kG��G3ɦ{�0����m�=Q>6M��t"�dy�ټ�R�^zZ�qL+�F����g�W�ᖻR���5�G�D#cV%X��pLX5r��a�ޥ#�O��үl�R�����yO���Zx(T%�q�;��7$��T
D��C��&+��;��0^��ߩ�YQ�P0dκ<GH�YO.CqM�l��w:wè�q!k�f��2D��V�H��IVK��N�F�6�qʤ