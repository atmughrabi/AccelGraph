// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F9w0dCSgFM7GYBwJ+Jsg7QnEWiEUCh2k3UEpjv+3crmpCOJgMGAEcIKnAq/9LIOB
PMPGkmJ2lHvCspgeeSJCwF9+ATwfvCtqdNCgkZI3el4ZzNJJCZNgSyBCWbc7DWgu
mWqDDnGafgAZvnH4W6Qg/d/ro0QtbZrAQ6OwY5yRuJ4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18016)
CNIQsgCL3VU4Y6k+9078tWBRc3/0cKXIJJud9Ltg0UU/hBNU1yPTcBBUNJ2F4Kx4
x3tkUal+1lnJ+Ky2RV9KJrWgXyhM4DXrhdqBgHO/ezcfSqUgkD5qm17IsFoGCHWE
lgy8HpYn0OAeaMN4pSkTqZRE2j7v64ShSEb/wKHxe2Rrw6j+wHKoisUGMORn6S0U
iuHE872w+4QoJ2N0iCZ8jt1Lrqh7hk6YkuX1BmO9slqEfLspoXr1rZdHbbmpj2/d
eGclXMHyOKtERbCWA/+B5IeGMu/qadv8AAUPCv3d5luge4B0imEaEhYXNY0WtVfL
956ISUxnA+MlRtXOq3oskjEofKw7kLKU30AmLJM7YQafe5r7RIPXBbMUllosiZJt
VO/Np8CwzOkwj4KJ+K1Fc3wUABrsoZ08BZAupYCqHHoSzzLWSS2kNCDBdLcB4DFE
XQ94i0UjVQ1LpWQspTCAS68OG/o2v07mAz2eAP3DNguV5/9Mcgh2tg2M/S8mV14Z
dslbRtTTzbWHWCykQDNfxWB6H4wRoya+GdbEL3kaWDMefUFA9czNu9WhySeOwJm9
qUtOqNMtah5zkDOMzCT9CCsKgSyloTWqqo3D3kw0hfpxUmeiiVuwm9lLlCEzakHX
b5jYV4NmIvxIn3+sEXWkxq0DfY70Ba91/3E0KfHbGHmSm79d+tM7dqX41dzAft6z
NaWzP1hFC77+tIgnx3AMv4Pu+EX4CJOHA527kc7n3NyLciYRnG0WlYpSFxOGdJAn
uB+rGFeP5KHkiRXAF+Bcc0NW2XXw+ah9uaKAAoL9wWUPXpSDbrlAV02sQCYLaoZU
XaUpRVLegiUf1kyeIvGlIIVQ2frbOWYVoE9rDZXtNxvURzK8/UhdT4FFfLyKmIeJ
SS0D0YJIoa8zOzPXgqiG7IOga8GGs75y7IMbknAiDAIImfHMTE8DPosZH6fF2kIK
wJqDfrt66wQ3yLRmhH1eA7tN0aZDd9y9jFRfw6uTUCum5t1kc5fG/Npaaqor4SfB
5Mq9yXgz8ihBRwQ5nIKzMgo36CAmfXVNv4boetP/ueHD5LDD1k+AfZskrvbUaFIT
MgSuCwBDk0sr7QohPyzZJmPvZyGVXn66WBio6utmBf+SvxbDxJoXGXcFncgcvpV/
mA1WwxSP3zr29/GBIHGsZJiar6Urt3aJ+VzmwWYQviXds/zPLfoM3m+V9Q7Jx4Is
jZl6mHdROjoBdw1tBPOPtZsXUCofykgw2t2dNvguaBRYvCrjSNXBG7N40j4XlB5A
nfGzVt1c1ZNOR03r9q3LvOP6H2NpZwQVKvqD/E1COxZU2JEBXIPGpb617CJjI17g
3gflKpg3H4SSOcFI+NpmTIbNMa8PPTeAWY/MvIGf+7ACm5MOyIy1gNHSl5oZpb9F
goCxF1VoAkzcyU0da90s7HkO5ssSIz9/votcrRlCWY+QBP73veIiwOvKnjDYQ/8d
mx7DsRiOF1nahK1h6PNanrjtuikrb6oCWOznjlkgnQmrXpwwcL+gozbgKk7US7dR
GnLcQ2i/jO+g/BXwzsETv7zcGAC34mVDcbrIau2a0SlR4RWSYceEKJ8l9QiKG13d
5ZZDQwoaWJqZFiUbAT7N6CoZYFwzaGel+MjXQb+G8PMueNwRsC3GYgSjLwFFiLLU
mJpke3idjOY//EOrb443R5a1n/FXn2hk+o/DUsm7nhNZsAcpwoppRxWI3oytlFEx
zj1b6VmU//d5fE/b0eXYexf8+9D7InB6UE6UGRPbobtfH8TL1rkleJ4hxF6XbQrC
GjIt9Tpj8eOwUWn4q5Wf3gggJuGARM0kFIHG/8hef35QaMiPSYIXbe+EuUMj0pKo
40M3D+GV6uB7cPPfZ24KGecbfX5LkBaxKCX8RYgG6ECVd7OtbaJV2bR1IWIV2ZXX
asBGyO7ayAvIMz7/+b1mux0O5AA3N4FZzQcLOtBzLkTRgmpgwj6M4ZjPvevibmyy
z0FQf4bMtgmPzPUrndf2dx7caY1fxJkhR8OwMv8u0URJLzvBMToZzSiajdNuUg06
wV/EOfKvXXy1Xz8I75fnw1/LwNHdWfssMGmikLy3Z2LvLdaCIrvITIy+A2R/GTsa
sxWET7FXQO0RXlaJbzPhVH+JrES+DlHp2Nru35QVDdiu5gZ4Dryz5vdS6Fh5XpKm
Sw5lvu15ORGBdABf5+9Ar+50wD+6RNS124ZMXGZ7grMSNCwxx89UJk8vBcX8q/98
TkxD00wsVJ70HGmMZL+L7N2pKkb2Vcsiyf9V2eiEokmo3rNmmyz0pmsmg5xXDHjw
/hlb+3yyNwzNZPDnRuLFjbW53uUSKqsl+wy5tfK1w0pDwilI/XXsltEAwj+izmNa
PC8DzXqkN4jrW6BJ63R1humD2AbYMmKsxdz3ZrYVrDaFGYWD8UHGdNKxMPKjHJSs
/CfiYvqn9TZQHTStD6LfIMXgSVqQhr0dm5FSg3D4hdXtJg91NLLkaLhZ9ZimUy/r
lwbDGhbRLW13ztkqen5qEHCADzxpSKr4t6pmSTpRnKKK3bixKCiNkYKVTnVzoQ/+
pG4cNDzyvrI5tMn4asuKKX9VO2qOTZuIGZsqKVSfa3v3Mx6y/cY9WAxrWLOjP/Je
uoIvXGgHDxORgKZLeNjqZuxFtciCSN6ibf/SYTJfiik/XOLujLYmhzdVIegLT2Na
8BWIq9vtoc5Zj8Agy5FLM2QmJQGEA0NC9hsh+U6F9xqn2NQK001aDbscjtS6YtuG
xLaql4ysB/+Q5kWAXI2oVn/GOE9oG44/dRqwCmaH6otbPm0hahe7AoL9VRB1BxY9
w/KucJCHx8Tmrb8wgLb5JwphTc/JlEaNZG1Tt4sxQNn1hkHaCesbuQQO8ZgfqvVW
h/VAlyHvyfp3I0EBou3kKA/8X9r4rr2q8G2QI1DDLzkLPclrxKezUapXnmfq4q+3
pEnKkEvG4xXBq8nja4jCrb1ugD3zoPexAK1KoFsvSsP9uA9C9vvPk2bZfgunrHeq
EYBufiPBQryVhMw6ALCI6wOlOQP+qk9S3EDXG9QBTNvqMH226V894Ewj4GyVOzoS
PZxi5G/uzGG7ff7OKHjQcPMoc97Etwrhe/5DVxXbmo4xpMf5d+warLi+3fJt4gxP
HkAHs0db2envQ9Aj7ihX35AiL36UKZrbIYpKGlreSAcKTOPkTs/NYGuSU9BpeujE
siRRVfXalVxSL5Vs5mDy8zF/RTOtP/el7rF3De206C7wjJ9M+TRvuepfZcsdAyXm
A3agZt/2zPjnmyKZE9DZsyJMl3i4rGFm+flVKZUU3rscHb14eYr/tYZe3yunua8/
yPaxoIZ478ORovsTcjqrcpRk10nnoYT1pJyBrjPyoGTa8wot4SErmSmJzJHUgNM+
V6G/YH16lx7VsShkn5OntQ331IdEdnro8Om78V7TmsDGGGyXYffJIMCkBYCWPohk
YV+STIILBoMrbDlLjzJF5+zDpUI7JXQrE9jiM2/JOrlc+WV1lcSIUb9OJ+LV0LZh
TXm/yFh36gRgKYyGrrS2yysLns/DRs/ls4GvdEbOmJcUm9aSfqvMTuercJWb0SyE
gjKXmUKnNwlE+stuURjLDZIOOEuzoQYSSqZyzEXoSZuZE+K7U9a2+vDXlU2U3Vqe
/n0ev9fPM964zHOWhecnYurSJRnFm6jPIlMSqwXzbKGAJE8CtN5lZ7MwvraQ+10A
XE4PtyIoWsdZ5Eo4Ra6Ru8Wz46SC7ytw3UQcfN2vt18ZLZWyMHpku61JlyWRoZKF
JtAm8GQnkMF9jjhUULs4OU0reem5DHKwQEnaMLJOaOhUQr7b9zjrj0b/2cpbaJt7
4Uono6AN1t/Fq+v766pGEfJHOkLs05C/E5ZVbGCbSNhhYfu41lfO3lKPZv6wLEBZ
vThkhI+mkFsYB5AruksPsjbg33vJ5Eqj1AWfur2cNbcW88UdxrlCpYOrdjcjsZSo
/IOOt2SRNrzhNCHJ+HSo8R5yikK0QABAYi7TFgD9YVT53jxPF5mc4Nr45ZJEyHCI
dUQrBsp6+lCkrt4OczsCjIYQC2gDzwZrX4rdPM4AXLqR7MOO/I8EjzrYhGnpuw0v
AbuMssoim3pqTmSKeVDBoUJENt4vhkKDHxGsb0QZi/ehG3VZ6s8Wv0Gb4cbcCEKT
x+U9U8y2S5mwZlzpKZv0bgyA2ZyarRnmMttpEP3q98slIlNJELlRrKpOyu3A8e3Q
tX5P2DWdkMB8UKrafewvDxO4se4YJtNRen/wdsCTtgrJeUctABZYr2iV1i/RIxkF
vq5eF2cy2YJkHSPC5qi1WZder+fj0PePSUiIv/qYBO0oDfvqsKSsPzgVK8UJJNcn
bT/TPH2fVPa0txzw/uUiKWedKMq+tszEJkvQYTxP3QLx9tIDCVsq2hNoABXY7zZ8
++2PQG3UuNbvXlhNy3I1HxgV4c7Ves7+oGWdbscpxWii1MvbNaI5AYsJPZi7Zn6m
WmXStpins3h+4gTPTmD2pCVlZMAeK/AhQ29xMJw6KMci9TNdQy4IW5+MbZXmgdtT
Tq5f2AwDa+YINTJxPPEUDFKecs76NgBen4IH/QMSpC4LKkQ0eravbfvJtirikXVm
27t8gcdcQUr4DxZUGVlthSwm9Plj9jKylixSwnV/KTItBfNS8IHew+CE3xagPxw6
g3FeAllKf0ZpP2H3LUafCzEB2B8uQ7bdVknG+qWGfn+5semN9JRDr4KlWfN3GWpY
BpsCdyYpvTki2wt9/rsOub1oDFYmb5oYybG/CMMTXxniOTvnmayz6gq5/U3alVpQ
f4H7ooeHQ5tyqhQY+j1V9FQzwEMebdErz+r2kuTSNg9rTz2AqqFCRsxE2WKxx0YS
UOgmWw0OQ20Cr/mKN/ha+wuB3i+TmnnWFEfv915cIA+GIxyQSbkvNggHmHXCIt9J
rogxMjR0TuDcA1uHb17kirr2bGabj5NgbPYq3FtbwUUrkvq0arRfnvDyrU4f9J1x
rtHuiTVuyOIRBd8f2ECUgvcq9kfjiR8UN9P2Cj+zs6WYMZhdtG6WpLzHe3pjM52c
TH6k5goEMI4DXcex1otZhZhDu3lC52P6OrtthpL46vp55TBY2nE8NOPwov89kb7X
13CWqXpBKk3YwjTEGtHvyYPJh+KTma3dEQ5Ds/mQTOoNYB64YIaAaq/HTugiVueB
hdmqNGmh+0Js4jRtbXa1RGLG3svtJSVMbUMkHGGnbwfYYkPUPE5Dda8aGWVTgqz2
InURntEF77IDQY/ijr9LccbjEh59omZhHTXBs8WCBhZ6w1ZsRgrZKoe6lFEjbQai
6PHylX4FiDzuz8hKNV4/PVYDkPIUMnilRmoTaBNop28QvbJ3RObamAZlgbdTEGKD
L9oHj+p4FjItFTTsOVtdR4wYFpbwZNzAS9dnISxNBZzBAoJS+PbU+kW2Nz3C/GLt
sttlI5bAzjyqCesGbZ9MDS5Q95uEId1mykEs0EgkxC4uhXCB7KdNev4gh2WMkpPr
erTe34pqFvFMsW2K+0PazGRRhcjSeqsjBunp/qHu6acbD7TndVeKlzBTZdvJGDJc
S7tuUD8cjJg4pdnF/lmIHG/QrpJahOtpQC2sqn4Ob/px10E5ohL4/gddVcPQfnEw
+51uCKHkUN7ulx1gOnoxxbB6dsc91IhB663o/fODZD8YwSasfWfG/0xl3fY8UpXw
oxIwY5RH74nsk9WUIRcWHnEpa28pc+XUnRxv0SUmOZ+akudodAi9TIy8rF+zq3a7
c3vqv0hJqXiCliFXME8b7Zj5BrTVXRUFj6PrjZ2ZVkwZ0sEwQaBNeo+UT5ekO1b6
AQOrbI2pdRkoKrsdH0mhuwOzDvPhqMwHt6yAZssgS+C6/big/XdstNPxGSysS5+J
tsXaFT19/3/mFZZJKEqAsVZApK0pYtwZIAHTCYUl1nRnOfY954QfLaLGpqhMwJK6
6WnnATkWA0BbJy/hbHBFaXjbcghZUgjsP320hh+w5pgsvLVUwgdaXw5UJLKinuxR
nk+8c0EmtItySbSc6MarX9K6qlHIZ6joVoHbmcQUHAR7mZDnET6HDUDjcV+E3zrZ
A0Jsf89SI61u+k7Dv1wuGlUTM9Y0YM17BqLjfwcSFS7Rzi1VNaDERlTuaIej1zkV
naOxgcKdKqIvLMqjQTuDBRTGjHD8aOvdTr2QYBho+3aoZz2HwvnQhdzv/rASto0F
bg12MY91GAWe5yEsnG5dYBDiD1+jLrY+XIakZh2ac6XRk9WTxFYI/woRaR8FETfm
rZyVul/o+n3W2XH24VyK0dmMIBuXu76JKi42LCW+3T1L0wcgctemfHQeKKHxkd9a
98VKhN4MAEWqlOkvrRRdGBjLIVQagI0fLejK55frq6UwIkg65tgkjy8LudBtv6KH
BWhIZJ1trIVwyhELaaxm6xLtn31KUwhRpnalGm48i7g+eghZBXPrTQZoNERRxN25
NDn3xClL3CFPOtjkySXfftz5V+ijROyd2B/JBrNKydGQyz2ZbbLmklPiJd4DWzM1
bSNiel53xHv3F+KcLmCAxoh4mqMmvfiF1W822oTb2ixjyNA/lBxM7Qg5PSjJ40BG
lHl9YEu9p+Ce66XMyUlxO2vV9+nn8+Mn1JzC8VV88lM2PvmqnkceZQldL+W3mqI4
L1Jk60AhY7lK/FPbcuQMqV7X3mjtXkHCwRYFyjQ38iOLpQ1S864iWZrvik7ZeBWV
ziGCiNi1ktyRnStkgAr1HkCtvCHKT27mBcGsD0av77tV9zgHqBw6EWLdMw5UFWYg
k6281Z3nSrGbrOIqbSMCwCsQE2xxXwVVy4eEWM/CV4fLnk3yp8GWTzRnheEoh4q6
e30qQKBqwXtEA+t+enyDubCusBX9ZOV5/uNKa1LvOtReU5+qarKDt4RCI7ikflaB
XfSfqHjABnuwDkj4lNBmGf9xxeHx12/bC0eRVmneBh/+XKv3egKO4vFPLj2VGRfh
ALUH7uCn3itn+hhFbfPUy888gtWqwjaD+OQZ2s1ItLo86MvrqRMxEeTlU1OCqkE2
QHSG46Gid4HZQThA45MbvvDEqrmYpiPij96rYvSsODBaHUo1kiRUS7f6rjDuxelF
lpN56Sa1Iovy6/r6DKn2An1urw4K8y7PNUuqItzUOgfjJtJ9CbfjXrS7ACeDjzf/
lJUDH7jTj6XShI2sGgauEDeRtHF8N5ufuGfCAObIdkzUVg8rICNeRYTeuRktiFEw
k/E2TZf/yoxkypX3wBBRe3x8B8QioSijUb/vHjD2H03120hja4OZUkRTGFnC/jpR
/prFNlIqTwNOCG8Wlb/EJ42QBtC/RiH9WidipSSjni0Xs8wQHXcPfEGsNX5/7Ib+
oeDK91PhX7bGcSth2OBR8mbv1fXNx4ubyd0Bd7azbImw7TISZIjbESEH1e8E13u8
cf3pim1WmKP3BODjtiPUd14b92wcK/B6g/A/XrkHjDEiMEX9XHbrQcIT9js+JBYE
YxKnmOUOMNPZrvGMrhK8SBhbmoRnH7WsyLOby57NB92I3pDZdwTFaanQx4LtJwOm
fdesjcMNvtGe1Xkm8WtJMMJCmMPqOUwmOAUgn0lmM8JyRr6sugAMUH1yv+QH6roO
aCn4TpLPAFwUBi1MLLdOuslv5TyEOEhWveNDuUy7dYGjFB7lNMPeIV/7xubrS9Fg
pFSKbmPRC2jGReMb4owYBJyd5ZAM7eskIA1BEnFrqI2X39nXJh0B/cRaRYoCO5xC
sO2sUSqjhr/7Uuy9/4xG9Ri5NTXhApOo4JfhhfMjJdlw5SFQGS5nRHysosghI6/I
QggGHNW74e05JjE/FVRrZw1GzqKPSLE9h6yC6CwM2xpsNi/SwUbYxjSQmjNRceK7
JNmubxzvyCgmYuaBpUaY2X+HS2o9Mwhsg9NEud/Al4NKICIhB8M7YJphh/xZ+Yu5
YUK8hyTGCHQG/ll2NSpz+R2Jp7ZzKQo9VGUzH0PRys3JIxP+U0Pae1t3bXXv0u2Z
Pdy4zfRNxb8ImZeKh8AeG9UWujwGOwD7YuOuffJzqgB6QYEOlEudn8VVeYk2d5hj
RV35FQfQbw1C++ei0elljOufB3PU9y4PZXub4mwnNN7VQv+/9DbQS98gCi/Xu59M
H/31tLCofEMRetNuJFiPTtKusiHRvv6BH6rwcjyz1lxOlYZtfOlpOTH1Hqfgp8Ub
1Ba6Uf/aZ/vz5qVCagu1g8VEqKAXsOUguV9fdRnLVWHzwiwkmUYn8vrEmeZI9w7M
V4cI4+XYniTytmEWWOPDseNmnP8UyjXeX1HIs1lWsdxztN+a3eDpwoNjNmoKqCyr
yEE/3huGSo/cSvh+h/I81In5EbIexZZGYahvW9ZhtEm6m9L2tfIiTJhv4cTar8uq
+rU/eTvu/6NTLRi4YYjqK90VvUCj/kBU8zggogC/g27qyUiYh0p5L4mYLSM5c1bj
cB0SEszwrUpqtsyYTdfFecgpztkz/usUfnBvojODzU3NgsiC3sxC2kiB+yjVW8r2
qM2Jp+rqEYNAddRndA2gpCxfjqRf4ZUYL/c/hBa3qVdnkpdVCOLmoQniX/d9oo2e
sN4oHd5kER5KQJvhZrL/1JfIKpFHTVT5MaJYSL2/F9vt5VnSPiypnZcV1xYgVFaR
wQCR4VWfsqbYW9ftbxynsH5PyFeiTRLBqv/iHUINkmGCKRJ62gRr10ohHgUuOZCr
zB0BBu/kiJWrY0duk6Qsm4wtzUUlvmr3m4VDozxYHaZh0R0cpdRKHU2N0Mr7wVMS
MhyciWZVUMWcOtXCwkFzy4IFVWKp9KrQJeHpNixvBq9O1pRwY+dIANzk4Mr7XuYn
nFuHrG7xEjyTRUUyiS/EdABgPCobYOC9dQbOn4mh6Wufsw1RXBawJg4hUvrh7gRz
pspQeSPe28mwYUNHc/2prZ3hDP0uGva8MNtQHHsc53rw4RfCC1XQPRgqws62mnV4
6GRYbFohdttCe+GLylpfWREW/YelandfIFMdhVT20N4rTR7V18ZS0vGhR1fCzb46
DdgEr54dYQjH0p8YX4tfIxZpzkntzWNN4q6T7B6ixz0oKZDsRFMSyZn/nVZTmo6L
ObZJAb0N4Y2Fa5EW6/7Xpt4np5UJvBSFI60mnr5Miuvp1q2kA/02Wd4w03v4EGqI
H9eq7t2aOWkXoSWq2Cf/YaDMnWcCscmkCZJ/0Evq7sveP7FNhi0mlHt1LiA+O/uB
IBxRT4RZcwMlDqJZ7bBcDZEcykQXg0aKOJrVb5DWniwCmfv85lumnemP2lSqQIND
61uC1dyWOdU0ZZ89xLHAm/Ljtu7OKWk2Kh3qDZnQTN6Djl3SBv9TqwlDkSmPbKDe
aCx8VCJ7gl3GO2jcmEqQdVbV3ZAA0Kz9uL/hzKfWlUxOyjN18yuUwWv875YCkcQx
VCGJqLwNK3LHH7VLN5eH6kre+89POqQGxj/WCmM+kPwsVMsc/IFNPgO3IodF22kh
Shoa3uU2h3YD66D8Dy5aieawZntAr2Zl8qffm/A9V5YNIGpPo+WOZiSAdlci20g4
YWXYTxeHsPeRjX6+dT9or0YBwVuUY868hF7SEnnfLIj8Wa1evQya6aRMfKXC7JTK
cWfAfO2i3hrIqxrjyE0dqjuddcUGkhB4wyC4PIMyMw/G0yHK97ooj4udsrV+TAGB
vlFQoK0TNA5DGaqtA4qchObE87nbD5twCa2593wgwYkGNqtZnKZQCA1byJ/+f+Ju
5OGlgx3rpV3OpHF5yAO22TSEVl+aJS28NTUty7SAdG7xlOlQg5N0v9O8iqMZTSfh
CI9CLqkn9pXLyN7Ck7ejpY/z+N/MTsBkcP3Fr6Jm8DMWM2t4H7JVx4pirdDeTjf3
MFC2sB1ElIBE/EcZOiqJz8SK3ih0YYfOoARaLW27agS4BmB7CFH59ZtUrYok7yFZ
NCk7fP75jY31nUCPGR5BZ7t9/cduILvWUPPw35QwSHs6e/LEocRyoDm1dqFFLf8n
IPuxRCdMd49Owk/evDJ2Ip0/tjf2e3gu8yZsS/HN9MoDp+XxJOoxH1OEIEg9MfkD
UmDX/FZVQz2CaBMCT+gnwPgHcCXFkFe8IPt+rjQyJQsQ0dwUBFveUOPFB2r293Ms
nnCGRZv7FaLbyHYpSl8l3kLZbFEyPTEDui6mzGuuXbtEZc27yfvGNa+nNCUxixL6
Pz1jnairylLzqJ4xpt8AZANVxXm9Sfb42EJb+uSg0W0cXAVCjzRtOj7uNbVifrz4
h/hty3CrXX6j/xbHBELELVML9ez9YijlzVsAiGZqeHbJozMzXGje3exOtbZIMxju
Q3Lr3MWaXkuI/rY5a4of6MZyTMrMj5+3jupaZczPT6q3aNZcMIeboko8iGGAOu27
ePd4O/cldKSfUMSnoTUloEXmuyd+er/TrDM6JfVZ68CqpyxmmzYy9lGos5NjqFoe
AN5YPxRGfoylFcd8iExaRCyjhju/0Hf2qQ54ZDNoR2KVC6C0mK/8H0KpAtEVGiJU
CPACG45TcTgQVETv3BkUpDoK2rgKYZV/LCk9z1DZJVRnIx7xI3Ett4IKBcAekEds
j5nKuGTn6dp4vYEq2Bv6gBSfLeEbBsgJ9uRvLXHY11wJuJKV5oRIrSC1Odfpmka4
+XQcegcyEv17gZXvPPWVxa9KKW81pAlkHlTxOJHtunrf+cN31SZQhFPRP/tfD08q
uyY9hZ/xF+wIs9WnF4zT2PbNsao5vcslf4QRMLhbHbUyAk42J3FSXTqS26ABCrwz
0GqIdaMIJVzQvyQDEWbBfV1iy2tlN1owZVY9nPsdPY4b6EvcMr9aVACIFg5MxAOf
wPKMqIRkbK8EMg2Lewe/p7MwRB4Zn0x4a8Bq6GEBLRMHCbvaltkc0u1UMk/NDG7k
WADEr2PandiYb30Wlsc/n+hxVmsbPko2T67nqCufnV8Ok3tddo/oHtn5XjhDAdGN
hMZKop09gSH+jubRoUh0TvxplyzKowWbZ/vaQtv/JBhesXVcWcfPIsefZ3I1qBJY
SCVy9CS3fJFfg5eiQ2AqarVJWdcawpMkgW/FRldbFU8i7/QcwEItOyr2U0aKXNli
4DiK4S3bibBurz1SiCSW7713WvL0RZI/3mJbg5a5dk6m51fnCx905rF0DmQy+PZo
70NblMg16BttBUXk7SEjdjWtZMJyBq9yfvyWrX7XaqLzkAwQitCrS3ZdNwrLV5l1
UA1H/Xkp8fPhbgawGT8cSRdvslMsHvef9xTMru4LBOtta/TeudN8UWiV2G6peoOu
OCmkBslFuUP67ewa6sOxQM1NSkYRj3nIAOd3qUTd8can72YVE06gckPELcvS11pp
ZA90wrdd9d8B76ROKG1qX403WuL0jqgbk92ry6iQq0o09LmnzwpLaXoX76QpTKA6
Dxn8HcxDBxV456f6Hwagp0FcInQu7ou10vbGTwNAzXu8uwq2ztLmGPM0VX6FYY2V
X7Ir3HsRk7Y5k0uK+A/d0oRiNFKIz9Ia0KmW+Xje5tG6doxa4/85bRZoBI3N/mUI
Gs2cRVKcVPAd8gFE/hjC5J5xsAFeAfDu6ZFGLKXC2k+Xffr5L6qigiot341P4tub
9ggpCik2UcpkHpH2a4XKTjNaVg3mkBprcERYU/VOuIsbQ1lIW6qMJRRwY7jSZ10e
XEArhw40qCCIzSqtdrt7qTKhogFXkfwp6rWrj49bdswlZiU2q/uqYHIL1c+fkFpi
/dBoGJJahs2EEOo5IPoyDlClz6uw/0DVchFYjiHgGTN7/fZAOzogQObAVGF+JQU+
zuQWG+8SNMd5uvOFWS5V+/VOMTybnTQCDdTNCYpLe5ciXgCRgCJoAxdVxWrXiGl1
5vCsJMC9Xx+o1mlgDZq82wBJ17IOrQwIuHWZqI1L6zGKSnrQLYclCmAZGYSi89CQ
dWl3/ZjoGbv+3codyVFqYH66iNcMip9eQd8vhw7Uq8cmGhfIkWcEd+M93FLBDNvH
Vms1Cf9JH4EY7FuP+QAxLNX1I64XeoAKsLsMhuw/fBx/La8aJjXwecYPdjalmZgu
RW7DWBoJzY3wrirSjBqLLbHnRcT5CsNoK9iNA6VQNp4tD/VYLXOe06r7LNNrK9fm
ibc66FE1mVjIGtYp/1YxBDSvl1yMbNj+gwzwBQuogp3MMefgxpJ1V7nxygRRnCt3
IP3a5FvWzhyuj/LETdpJynVtWdJqTiTj4fYmMpci8QEglSoLyLpxPxIaFMtrJR6b
8bA/fc3QKoUDiB7hrXCA2u27Xoq+kcHaU7D+g8TSdbmofBQu8RrBh3qfzrvDqkS/
VZU2hw1eI8ypXpmSLaIWxPFeP4CAD5GypkbGChs+Sw+NOY880zjtWmrWptK4a/mS
lWcuIeBpn86YAU2gybFryNBI6Zkwl/iZxIuhrRnOtPs5ZTS0M51FAnfn1SckZY/V
/LaXKrG5dEOYe7RPOb5Mj2S9fcHJW2sY1Yo8xRzKOcmRoQnPmdXjVjmc43ylYiqG
eiB1ueqsy7bmj4ZdaEW7hCuwTGNjaTFKq8OvAAkCGLDgacumkiJRlCSmmBxmXWbT
WwNOyVqe//wKuYCioCZynu16Hn/sQd1p2FDhtcgqUGLqCm91lEdAw9Dxihh4bmMR
HouytAuDkHCdwIxpe1f/kjntmuvpxcEN8SvlkUsSWPbgmZucaTMuNFLIk7PxZula
RjFZ8lGosUygZZjIdi5j9MRWgQp3RKqfBMuarEA8jkm6oLL8JAgi71UQT9FT8REx
hEzO0nLu3H6AHiwUqGaIfOiTt3CIxgI7dPf8MpVi1UuBuKZSf2fzPnYGjUbwFQlr
7MPQEsFzgE8iHRq0FgMcKYcPxECY0adFeYz+j8+GeAP3dkdxfwUg8chWTS+x8yVY
lOSuD1bNrvFnmlgkBX6Ypr3k/lfTfxeQr5lv6+pXYKPMSrM1eSXtAYU2jkft44Iq
Y+d09G1OHgQooeGBnndewiJeIy7P8I2Mbg+2C/lrYxotOpmOBEaOS7H9PWb+3hy5
em/Ohah1f9LopOORq2LqxUZo9CjN8frvE3SmD4EkEjckU5dYIyTBLOnoenAcNY5K
GVL/8RfOJF1WbSNmUar4CFo8YJEVyt4pcCDiEIhU5pt8WYxB6nAR3+AOpAFe4jcT
UoZOkAO+k/M7r7r0rDIA1FBfAwWSbO8fx753ONQveGS+NKsPMs4y64ibomRIaYEq
ztLzWArkQjlKAW4kmOv5oh1pTD02wBQu7/x0Ke3CEpRZIQF1CMFISGwey4XXdNBD
aVvatgOh03I3jO1voGQtjG+axzbfvTjzkNQfzYKKBQPZHsSh9x1w1jvCd0iDaQnc
VA07N4EQaDsbToG7ivZMDrYAiaxnVAOyD4oxxcfcGEaoG3kkoMaQPXPJfXLzf43h
MuRDJ6tz6CBU6kYA/5BXAEBFuwpLOzQvcMp/zWp9ecKS5Eb6PxFlwvDTB+DWGQrI
09fe/zuGFp3Nbtk5ZB2BvwXGz7nn1tpMkF5KB1XBLS0KqTy/6+FvdeyC/8rszcXt
yhoZLn7TAA6DEINjs1zTkoXcdg/1CynjvoeNiVOGwksm8zPuTLL/G6DFBRhSES4o
k+NbUuKTmUht6SFp7dIFYf+mxfzMF3LULqWuRe52/YUHvYn5Yxzy8XnEr1R0XA3k
qxpkh1ulGtoAqKRgXeS4XNAv/604c2Afeo2lulYyQfNxiCbhMcUiJiBwf1ypOYH+
dc2/xJynrkvFa2ewZj25+Fv/JY7728Jveetyna6VRpoY8BnSLZRQuOZ8JxtRs0Xb
nDtF/8Nsb+IEiCaufRgiwAFF0mysFIht8dFkI2/ScITb2ugF5LkxtFI0RgdiTjvx
+WlBsFJIBNNoKv5UWb88QSdX35lpBN3cwuzkfuznwuZHrwzMkE7zURGSGYdMGl3I
cSilqzwwrQZ+julItDdBIamRG8l/ub69RVax1frZ1Y66smIYv9Bwg1UEfGzMBF2h
iLSuOKCcD5+0zk0rPICbp99/FfgvSaoujYKWZQYukC02/ZZ8YICcQxE+Z8P3kEWv
YSZ9HBqdcXHVLLGVa2MXZm/P00krEDnY0s7gm0F7gbGK/fTV7llh9w8o7/GVJbrw
mhWQHfEP31M8cpaV1IIrudMrZWKD8zxybsoUC7hPdKv680hDG/e5JTzPlDu2IYhH
K6DJmWGrmWw04fDIbLhpYJ8/Nbz+SCNpQFNGl+Kqlt1CoxPG/aFSfj+zg3ycajpe
nH//iGxA2wghcEiGM8prDC9XnmK3swzYF3zWZe1yFopkaSRLldxd6hGK2+oRfjyK
3as0mmpxkhUxbthzt7vSqDw9e1tI4FVO7SjdNkeQwdI86qP5dsPScIVtXGM7P9CT
QD0JQepyKU5Y0PyM46AAnMzJ9XjYPDZZC0WgxPGuedyRug8g7RwI3QLJANKZMHdX
JllW7IY0Haq6jizdgJ+3SqQZ7IijQG8FkjwCCgtKIxv8/QPmLe6jdEQjHNwEtlVy
eI5YcTaaQyTlTuDFv0B6vHuQZJbTp5/M28yu1U3Cs16hZnr10sCJW84U4KYx3kQO
Y4igfL8J6xrwvtxSWBM+ARG1sUZvLRcscVn8PuERctOjQFFBnYmDuaIjqJCkyUvx
c9RQUtFuiXjYA7xn4qUMsnqRoqnHUegC3j064fIoNL3hARu8rBhQjYOHQEq2A4CN
c4z7roNI+zXpLQUMnvIfTWQuA5PfqdUD05h3bsFyCAyOJujY4OAeEKNrOZv7gHEP
ajjcop6VbiuHuyv4P77VBRgnRdvwHmIbHy8g2pMyubRJw7L45+wQ86fBwb76hAHK
8fqYfLFvpm+ydI9nTSXuYasm3JdNHx+eLPDIpei95GkMt062O7lTKvRWy2Az6axS
OdA+z5Clt4Iw7x1HuSia9dkqG69gdCndJ7VYg7LDKNdlLLq2tKBzuEWMPW4C5PXw
4ja27UAaxZlCruEhBXUncq/fnHoNk00/EDkyEwQtr+NoYkvy9F4ZaKLWNuh/yupL
h8LUJ845sXEweCMpaRbZcbWGcekm+3TvRKzVPcnMuL19KXMGYaP4GTvieQOPUdTL
NTbUQmzU5lknxWglNo4QYZ9cGXl5kdaZ3blEy4bNinw5S6jU6nyWEEbnq0NQjZOq
T5vjaUvSecDJnHVRFSct4vuzmHxM5xJo+caHJLYvKlcwY8gy2qyQJ/orOTnBvPqH
G8Yn9GvF1BC7jnLdhY/qStokTWZjl9kui52FKPFzfvUqru+mnknyUnhrLXno82cv
/2Cm+qdP00uU/Xx26PwzG/XzsDgUnWDRzFYXPbu9lON2x4cfGrBxPw3V40nIf767
rR1vADFkpRIKHdD6kdolGHDyWCQrFdipj7rTvW9oMLO0/jaLcX6bhHrRsjxuGEJu
0KuH/RgfuBBXkaE1ZF0PtGDDKzr9a6qFxnj/U4ecf4X/JjKh+JDiG3h4efc1FQXM
hV4t0cN+mleZAlJg0VjCPg545tAbxZnum5i5liQcXeMrpBc14YfkXtY2enJUGyF6
+OtyQMd9LlpgPADz3K1DHjNsz2Ngt84+ZBxGqiTuSz2sCgTHzDoZYAdEU3iyiT8n
FEVezRMc/SNXUQ1osFvv9rsQ/irC9296NQNpP2uHsv9qY2qOOB5NpICNpGG109QO
FrutK+iXVMWcZTKglkJA9aTrikf+KmGwxZhsoUKnji2MkvfYGZcPHaG7j9BhyYHB
SNYwoBrOeniM87Fi/YQG6LlwMHW0yz0D+jVXYL+zyAXLl9/l5DXYMH6gjzr2P8qb
OuT2aAEvbrISPSMIzFORwe0prnvoXINpU+ERlsndi87XwrHIUVvsX2HtjMnWDc9w
PEaJBo7pn/KSsbM9YobSVBsApMLuyqGU1o+1YU8pvnx8hMESCMLLJ70yYDNkQ8H7
zVjEfumHKGwrMc/2pA2aHnoaCMEoT+poEPGCDrEfrKy+A+BME5T7zteEL+W+m7XG
3TDZf4ypGl5DhX6+AaAlttRFhCGB5HqEbzTbH+7D8c9j9C/TGQ0M3VzRnWieBgQW
7m11E8Dxzum+apPUgOJseGtMP7ed9gOrB/TQcbVHQIC8YMKdHNSMknQZMH8QGXh7
Z0g9V1vl3IYvudvD83Uxo0GGIDzbjqMmwNh/pqXTVBJeTQUjcEfQ19FxXhUtRUJe
+TqV1Ntmfo/0j8bxdFkeQ50DqplXXsMe29G6G9pnqsOw2SWdWoiDWFe43fgFTV2X
ZR8T0WmFNYp3m0KVvPV4BBn7IOaCBmghGBAFFEQKtKEy8evKSV4ePTKUa40YaXNv
4qpDfjdiFA5/XKd/Hiz6pmNftWhZOKwyZDe2i3KW96SdxVcXqlb36A4mypUWXw8V
/ZDSG9TnFNGwxWw9amhy/830DTqe1rn7y0cnk5lOrZjNZuY9RAMOFApdBcgH2/EB
l7TPO0pE7b6zzKmQqUmClbwL+JsFA8lKV1wNXYeovJhBPSkW9puc7Y41oHk4FUuv
5VFI74L6tUEJS/3ZKWU8zBt2P+vmEq9Z+wzacXchMadEy5jFkC7it4mGWqWYSjIA
lVOgCtE2v+3estyMqUPNQbzbEm7GN10JSox9l7ybnCu3wuqcYXp+HAaXH2Eh4Wd9
WG5kGVgluCPUE1aaU4IV2BEuNt8WSsHg74ebx6AxIc5okSuOqOZQ/O/DUSuFne3b
QvXQ8gXRXmN7PTO09LxwRBze3xZUDLTy/EG0vhaj5ckjQTpJOs3SX+qzzDD/E+T/
z7FsHFo3eg1D9OzUwSE0ZyiMC3suqiAzmFitMx+JFDFhxCPuTBuO+MZ56NlTySdF
ipsG+Rh4J+qqsG10HADWafx28gr6FB4+zlUZhJy5DSFQcxdjNEl+6Y6oKo7mnooH
5veKPvghRF4EXD/XfTONbMzWM/azvxNHgQj0zN/4VVG+BVmBbkSP2HskW0WxtUUl
1omLX5oax0oa6DA4JK+3bctPnTUcYDm3lboY4SN98N+wwxRysvTuZ6sfizTn63sr
U4Hx12pVCXXkmADrZai1VkRG6l4kRWyWHcGdaso+zx1ZD04GyhASmrqIsRbZpu+0
yLqxJ7pRWpiYxTxBUx0rAL+l/+hE5FalVAHVjYGSPmtx3U3fD6IbVTcFke2d3WwZ
HI7XLWNcLVYYiyNTBazadJEyqbGftPU6auvVTa9+08EItxrwKF1I8W/qRNKRzXj7
mARnXIda6dJgjvyLEZmhNeGQTCvHMADVGjRwZN2ysc/C9yGPbHzk1qynR98+KSFV
JHR6AZojjvr/Ei6/R3uE5B32AvV9Ea3tMP2W1AgMHMsImMkiEeKKCEila2sjNrlr
dYWyJTUPqBVb4KCbgI+JrC2U7rSEecHVCnnrRijO5mZft1vCfx1Rs5T5T0L6+/sM
QbHCs322V5DcJbjcfgQXBEVFNHqw3Kkz5ry+ZpeJooUWHjwi4T7rQqlLBvdKUmZb
L1GuGONmIfimaiu4mfNkH3wPqZxM7NReNzW40YfxAJO7TexBcgEUAioA833DuX/4
N+1MhV3LirIn+U+jLp0vLkajzSXIwlFgq/ofpxm+hY3b3w5bz8P9QIppzEiUIFJU
FwfP2swfpXuWK76jwuIQqtw2srrU0jjy6PjhLotyccGCFwKc6FjRzGyie5FIsOng
ZSWlugqNDhruojAuP1maccTN74N2/sT+fcKmFUXmhOAiN9Ptl8WkhXd5OYT8HPz2
KjKXQK7NM3Dhij79YoA6oABWqji0CBLzj6Y/R4LqsOhtMo0BO3G8EeHMmkB1p8VJ
56JK0kb+aw3o5iBnJdIpCMX/5NyY59hWbEqhXbbrYMSaquV6qL0d3Orv8aKhYE/p
johfcUaNdXmpWmxLL6kgy6wZQzV5oLVbSSF4AMYz3j4bAOhjvdld8gsvv3qdHVxA
56TlQAUOEXHqDFYosOItD3gQVGl36c5mhr3eRV/NFeVrgkjMG66LfHqXiPT9aWHD
Ex7JGTQu1RkV/Y1SDQpjnpn3UHprQ0g3gWg16IY5d/sbeRNFPuKLZYvMRgVUM7vs
eEw2oqvhE2Grob+MZC5+n16/nrFmti0YR0zkLixghr1DE9wk8h+5yjfjU61gPSgj
fnMBVUZQ5IyW65YpxuYziuqidFNL7yBlMqvYqLAB4Nbr16yPZM0Cmm9h4/GwrUhz
+E7NlHUvjMBJMW7as1k2oJd/ktmJDORZyhxk3Wj69TUnOri4k7iEQUVOGoGiag2j
4kmQZQvWbK1Iy4CwDt8NeZyQpH8w/IY0vDY2RsLTiaMPzjqK05ULwrpJO07DRp7U
EHtlEYItBkV0pm4zcmHdCRAEym/oHNCqRjfUPPfi+60piSJkTxjivAI5skNr3xKd
ae1DGMoh0K73KzCqD3TKnGHnCqvqqQ0d8ogeez4A047B28d2ITL+15ZAtcv0dz6/
xRGJoIYqAVhkDP+HOUHlTvuYfqaATTxpphcxwv90mE2jcW5vtSgEtoWqg9dFr41j
WMUJzyk8ei/GdV+ekFztfDoBgYQb/g22ynaXALq+AqX8hzT6VYMtcMV2MY3t1G5l
HAl1nR+aIsXXfrevRhIYH3INWxe56dp2fco7cZBD0c1viMyniuTRGKi1x95DANKu
mw3xXOC4rmm5Yxe5FcUsM97+8ZmdURhPvlos358LtBObVgYkQBsjQMs6hqKtp6yU
YiU5ZYUz5HJAjoosUeZZq/qEaJNeyrUptYLfobNR7s7rFcmLAPiU+LAGRcgzjmdg
RjiFKf1rz1fix0uaab68EUjcgeofFFw06Z4xwcmDXOR/RTVub7vPAe7Q2KBhIBsZ
/E5SsmVPvlCxiqpXDEuS52AjywZDR38C5HlNEDAXMh/RonAksdVS78fz3c6gpqUT
78/tIJKQoF5vyrMDEu0TNn6+8oCiYgw7vWK5xt+rjlcrDQjSQIYjeAENo0RoW28e
jaoaP/mmh2DsKpNyiICm+wFG9ED2rC+pI4va/hbhJKFFT6H+gnkjlBLPPtHU8mbr
3MudkImaDN/JB3Ujqx37xHAxqEAQ5ti25gZYiCNsmdYDDZf3R/jHDiJK8L6yvmpk
b1OpSa29wKb+eSOH10WnAEEeWnfPNrJwBU1SZlwUC3KmDtl/PvPfVhX5O4MQOxaP
6RFfGRIl1GPu6L9p6DmKdyqyqaMmCHY2d7QIat4wgs2xmMSWq3F1JGA5+KudQ8z9
auOX899CFoQAPyxPgWoT1Q6MzXkJNR9tzHjiHxmM9D7XH/5HCG5QxD4Rw2p/1OMr
bXfKv/XHvjWCB4z6uNr1bJ5/RuI9LdTdhzO2/YP8QS0MSAFpE9XmdbfWy1FaNqmn
/nUdA1OXQ+pFlrUuLdY5wfJvP8vJaq0F6g08P+WnulY8Vj+buqU+wsiYyeR2nfyM
y3DykasjcJP7EJnFGDXAZ3rlD40m0Fxn5K+Qtepd3j9UiXgwbbQ044umHhllvpay
i9FIdbjFUk5Y/IJsh9OO9AaGoiEaQMpEFs4dS3o4MTDNv4hFcIq+kNnGFXXdoiF+
DCokHXA65wal2FtjDIw9Oo1UaxWtmBtMss9UXKCtpYl4Q1HdxX/ULgVphJVTT1OX
kAP5OZ6BT3DxlqCOS9cwEei1JFyHDsmUQmH50nKgH/qd+UZbCdsV0NWvKc+0kre2
oYaKRFVFJIN1Bk9tPj9mY+uHmJFI8IALodMpngU3DG4Aj1YepVI6XeDSHK/bTv4p
uvm/otDNnDGNQ1CvQBakK6KgIm85jrwj6MkEnILru78FYYJwBqmsha6A9Pdaha0i
7yPp5IaiNW6CMfUWZNDGWExFT1VgcluV6fuqUrlQ0VrJ1Y/oPGWF4Iq7pyZfCgN2
9JMtJJwQLZrRIGYONkXiWHHJF8MOYOrftMpQobPrzGna+iDenDBDzB9/sA9Uph+6
gwoLHQ9VFI8e5tzntq+o/906OidAsf0r4Jj6KTswbHAhs22LiP1uv0wh2FTKNHPC
8ZQjx0A1UnVA3rbgoOvjXTAwybD6vOWHPiEggKtUvDRc8J9Xvs24Ba9iK3cBmVeW
e0mcMM73iW7EaQN1/fGRLhHNqDmK3Ys5cJdqwGMhuUUnoi3uJ1je+M2KF2kJJ05q
5RBX6vkPV+yxORO7QpHTpW/EoyYtV43RY3UopFsMPMRfn8i9Bj1n3HX8kcETNjDQ
Jqy6z6RJk1hDRmOP4GJoWbXtdHAlYYDUHRKjHdXyBrjOtOEl9FsJlliNZXdI2/um
VWlRzgyBWqk9GXDMYCdGyjb0B2HnyCIv0QIWBsf6CEZkaX7zosvpqXDcstnGN3b4
58VjfHo+aCVj1HI3JGO5h76S4qy4TW7o+Qg50DIxt/AyHJP+BBK45kimSgXy6raF
GOooIOikZNdkgiBmgY16C/te6X/I6A2XF9CtNhOk3d3qW43+uChEVvMyVU3DiCNx
vjJIELF229eJ5ObdzGajsiiWPO5ixXOnNIqTUxmh4t7w/8VyBDueAE2hG4Inr98/
It7fijTiKMVErkN3HdhBE0An9mSBJD23mE8bVKIA/8CSldCt5edvJ5ib+NVSSuet
8lsacnOr8tWQLPo7anrP7K8LbdAnQsbc1UlWXDe917eYwOLGaZ+jPut5+kBX7o29
cV9xUAmu+ScJfjbgcYT7ZgcoKYBcgVAKqVAkYV9uDzDtkBiBUVDoncVUoDr3tzg4
BQ2VMzApwqgmVQncAHzqWp0mWdmlSkKI85JVjQEI16cy99JEf076yXu0ZyKvdEbY
AiOtl37Y1zuNmxUOwAWv/fYm50ZPHzKVNZHj205F/QVF7KD4jMExNRbfoYn+Mih4
vCSk0uzPaSCHDpzq1nxJBOJoqDCIrUyGMsKovXjhUzh+hh/u/U+0QHAWofh3hdDl
M3y6Fn7eZABMfidP3HupT/pzETQHgCBQH6/y6GqoRCNPpbYBsEO7JuZH9wt3Bmdw
6DsGXEbZPwBmbny9K++OX6QlNyeUlWvUbnHIeZRp3Cs9/5jnrHs7nR76R79VdicY
PWKfMJj17TC7T7LrSjeAfO9Mwfgjmp8Uk/Nn8qz+/wD903WZH6chAl0ndrXm/Q6J
IMakMufYqoybH2DB+bHkPSnE1yW8HmlLeoOK3oisGQ3kI5IRG7U/F6PyfoqPVohM
gspehwxbizPKbWhOMxg/C+XhjSfhvZiAjE7ngAJt6HDIsFpKchPsyNsP1M/USLPi
GK5xK7mQLxn+eqvq1Osu7bXy+ut2jPWySa/w5J5SZtJomlg4ufboMife0i7JicGb
U4RxehuqTnSazQ4BME8gFX5Z96XAznlJwjJmzvrGXQHpNTpCVWmmsMrE/kyobyAa
vM9MIThdPtWZmxDVL7+3paZguseuxq4CVQQqVwZEI8ZaNQKJiG3kESf15pu35b7o
vz3e07uU9/K7OQteKfTLsYqs65Ci2pn8/vVa0YnwUHDdEr7dpa+c9MjcJZ2ry8He
W2Y9bcpv4Q79GdfPrY+vJEWd2A3jwM7Lxy0okMzBWqWuMdOCpEJvzKCecM+K4VsI
Rd8OXVsrEonFU1eMhc6LWatwVRGDM8k1BIYVQkt1jYmd3VJGm8tQiYKBQ5a9nYdL
efoA8khRDDn1YiJ9iPCvAOlTYgJbTvj1B1SmxONosvXaorQMJRV3gSFbfio9j/Jo
7GV9I0A93rk5OCrz5rxHnd9Jq6J5UZkfL4fVRRj2JPxyjtbAXYTAQZrpb884wdfW
EnQ40kGYUJUoF0NVwbjgaaONt0sow8/xaNCYZ3PQxY2aWIK7Ajb+WwubSsNKk1vp
6QovQN0mJGlWxCJhMM9eUQcBPVeM7wQMnt0SLzLIGM+Nidkk0nn2+b6v9G3WZm8K
a8Pjp3dQdubYim7XaoR31r/BJmB8cI6ZHR3/ITPCuv6MFUnrOn8BBrozg4raeXli
obcurP8LbySn8zg5KkYBVYyMbWaBk7huufWXJz/J7FUCvH7p5I2kC20KyVcUcFy7
cRetemXs5OdycQ3fXVghW3I3Rov5EdCj2KlF/SR9qMKbqz9iaWCyhAmqtaageF17
4b0hfPC6SJhZNU6iiTfBXF8XOCPqcB9U3vCxhYu4TPxHNUrdQng+SthLiCbGDvt4
dQ/nWwn48GU8ARIUwWmXkpsXeGmjN7q4smErrvBaayUiJfGxOWlX+7FZM8p9f3/a
UGiu+eQoaeGo/AGFiKZz3YQoxM/br/1BI0min+URZpnRQYojOTEpbKnhniE3hCEL
rpj0uv/8Ae+AENFSm+CbcdIbepbpjI6Rppd+i2Gd2PD3DRlu7gWeHjBvKADFViWe
nXiL0VgKPhJ+yCcApiYb+PymqTf+FMOcP1evcLpsZcLiX/osy1/59EwZQSOzGzGH
Nkx1eVgVMY++waabWgyqJyPPCZNWscgmMozL5v1163y08K5SN/sXIgkau7drp4zR
xDODyzjrYJF1axPTMYAIIpFrIg8quLKPlZ/upeHGspSC6cx+mvZmfTW6QkT9PXZE
9k88zOxxGzirhSDZalEYfHsdSfUnjLSCqOPyKf6p/cI4YCZjLvml4x/Ty/6vo9IH
gaIK/0m5eJf9G7EJR7J9+RHMIzHXRMNOuCkrdeUx0vZns4DfacTys+gsNPXHCDHf
ETVeHjyeMnInGC1LPMYcB2GDylRWWWFC2g5L53Wf3y+nh/tNNfRszGA0oYsGhN4d
QQhB955BpcOUqgt6rJcIn4b/CqTC6OCRejjRQXrKVlN7aseOTlmzJw2rcu8hZ7Zz
nZDQkvISsZgoDK+C/pXPrWejjez0WPuYWpmkMe7VrQ7vYTXCaKdDbzMBL0PonKRN
0jYtM2rVwU/EcKaK4CVX7rxwOPokSke5QE33zuV3UdVkqRAaaAU20Zh8KDN4Oh02
62oL+ZHpMLdVBQ5f8hU6KVxNNUjpy3koAhJD7KW8ozu+iNfQK88MAiOLNNMCL/HD
6RDKDGv7L9u/jcaf3HGB0YXC3ihBo+1+dUp1TysSdXL3Y4nylUX3zv5crWjWy3Ar
e4JpvqSPC/5vthqU/TCZzWY9xK3cWeEtQJ1A4oB2IgFYwj2vqHhmneqCPIE1sUmM
YzNXLDAw5p8F7muqTk1uzz+ZfvTVqqK+RlSJIWU+8asFpLYb4aryAPgQtT6G7Mjp
U1tFyGB2/sY5UHfXVOiz44ZmReHZHkqUzH+O1YZ7gzysuBBTfeqPpI0oFcngS3nh
WzY78BEQHPDApJCHgYhvcsJuPZbaGhEwWDFRgouYkCjTcbe/5m9KnDXxkk4q1yMw
wnJkTNUe2yow+zbAYcnCQB5RZwFi3373HytliwnTlSF0YnRkRtJJYws1yhP2Fonu
LpAbHH38+7DtXdg66kGi+YZpqySZW4iAzewm46cMeomwEKt+oy4FMvU5qGx5xLNY
soMPVvvDT1lfy14fWhOtoakvfXizmOQoV9n7OSD2qBN6n/Cq6wbPqvwom7flWGs0
PzZx144fy0PKiWQuOHmWw7ezzhROMRzFjk1Qt4ifl+i4/wuMaDq5nEs/W+84+KW9
IT8AqaY4b+qw8qugBqxaQG0EAtiVPpUj5lyHv9XUOMOhotZUcdwZjIis7l+esqzj
RG7/XZmmiodW6Ur1RQclhAICPSty46sNTc/XoZtFEewULLEAIrvMsgG3OAgoOQJq
GmTDT/yW/2zX+uTCwEnzATi31b257VGfe7BVWrve2ezeO1BH3j5Zls5QllfJ/6Gt
THhafBlIXBf+ovHTLGboX0Bux0MAQ2hjY1Z48lCGFoV6EEve5XmNPIFOWuru5xwy
Y1xssItUx6KfjnwXPxptAVr7DjVkEQ8I3Zl8gIOcOXaV6FU3CnYoSAyv1jvxb49I
UDwwK+XlAPW9a4RKL+pgsq0enhUJBHi41uH+B36SB9A5Q0FX7O+iZ/Fqm3BBY6Cb
tdEc7tITcIbpP2hXnBDJ7zr0nXwex/Hyad9EhxZK7DCF+3l2T66TzVzhJ8cMPZpC
KqPHDyGEmLw0WAnQBe2I7IX3wec7hP/L6ADBtu4vdPIf+0MtVdS4WqDPn1OkKmdx
ACVQcDhj+OURcIL74SZFbSgdRXkj3W+Zf00S08pxmRoVl4ljxw4wXphh6313D9XQ
SBGLDGTnriYIv1PU2shUzw==
`pragma protect end_protected
