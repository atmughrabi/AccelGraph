// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ECjriTLBwc+FIt7UihUAdleYhHuKkRXEnV9QOtzGR9QEjIf5wkf8BPxyZ8xClZUo
e9p5vKvr+HYn8iW2lRDHx7abRrd54oOgFLGAztpphn0+QfoGRjkMGbBOvgydNmwj
RSBFFDxN/dc7Cat7D7dWNcDi0yizR54n8GsfJPPaKSQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2656)
/0/27ou26X5WXzVrRQjBA5QHoVZVoKiYBYhqk8QM/T7ccdQKcoRNYYKtBcLYgbfa
rfTwUXh0+6h2LOFcN8sxQ018Dp3y6m0+JDVCQKoMxtD3kUIoDhTSoXmf2DpGKjbI
ZaaOPNwFR8Y8sHrUcz9IV6zUdBdSww3Wj98db+YAdyFCZeaJTuqaaBjcGpmW4Ovy
x1IYbl1lltM0607kqi3L86HRNRc4MdRIm8Rw3cqXkQoKbhDvrao3QcKbSyQOQfLU
7tUtZoQN9Zybs7TtcD+DUpQIj1oUzYjJ+kJWB63sHPs1s7gU81N3P5X9pNt8/SDk
tn4UIUPn+63ebZrSkvcFBMQ3hmJU/+ix2lcmi+EyNj7DhTBuWyJWTtYE4gtnlHLt
dSg0g9YNSCaHca9U1cXA/p8z6BLRa9/aa9BABPXXjdfW4fH5ehW2x3If0+Hacwsb
Ayu9EpMf5rhKkMEYj6Ufabiz07rT144I0By6AKsDdMIPeLMYdTziYCxb6HmUIdqf
6Q3Ib6Z4KO8neX0hNLnNVG22DSeD+ZtdiSaQmoEMEdN1QI9nwUF578OVB0e7EZCn
BNZZrMt0odXW+E27+DTNC/+3SUH1nUbfZ51US8p2f72Na8OXokYTdNjdLzQHj0Aq
ZKmFySnxAVzhHI3FWnGUD7fW9pi507ImWbLhfUBvFTSVsOFhQv0C5luRRBDGQeUf
ONBIQBuj7xo2vTCbMO1QjNQSEjPOysastgReYnbJqhrlP0bYg+vKppXX4vf8F7k3
Hx7wYFQKP7dzzsZDVdU9/dIB7a7Dn6E5xYHoQwH4o+DGxUzD8PE3nY5/kOGrUCd2
eYKXf4+HWkh6/JS5t0/V0Stja8Cq3oOB66pKYRMoiH+xw6HkCA549zDwiOmPSxIn
YZqZ8BS00/oDBJ0UZEUm/miISiwtJvO1QMDwKAELAROEmzbUMSE4/7msMmcRmYCF
+zNJx6VfM4iICZNd9V+AM9rWeJDdPAq0VkIyzseicLE//BdAa7NHJQXugWaXD1Om
Wids3T28ogGZ95C9j4Nrckwp39vqSy3SNIkDYsHMQHqBm4uvAOBDY6wl3AsJuwch
dHuzoV2nvtksHu0usZ0h8IRBnuT1pn18nXacnkaOFyBHlQuHY7dvVRewQJHRn1zM
Cj5ACLUYNUaOD7vOKHsg8Sgd7VCSbqpY6fc1gGtMa/TEXZOCSF/1TgaoCrFTcO/H
ghLTQ1YSQUS494EPd51ndKty5aFLWWYtLSFPxNc+cvqC3ImyYqga0Y4akibNWD3t
KKqbQ0/1bA33iCT6srJp06IxSxlIZWhk3YusE006GqVT46YfqkoOJUuEJUup+hIw
g9zfPig8R0649RIdXFC4KMPPx8MIsNuBaqonrbXLQJjN5Crtr5hLC2u43cSBZpF3
2jUkuGepqqPhr5xcjoqcTwloo8V4FYEGtW6zkWzdIPgDtQfb/lWGDXRcOmVkmRzm
ql5Yv1GTHz/hwk2QPAI//qULixbA08JQ4gT1PCI4wQEYvVer3rkweP8OcFYZnDUI
j0SQRMLh1HkanSSmLrh1+77jV9lt2yK16NWDUEiRyMhwUSjfULzeTBghy6wukdKB
0jUR0MQxhtG6uyKriqKSweIXGfijWrqc77o4gR9s8ksmYcxZ4+ppi1vV2qP5dAU8
OglMhO7LsAl1Tj8u3+3fxzf5oNQQDTiaZhDMk64GuNs4tqHdfLzltg43FeslrTgY
gvFDUYY+ceGaGwDLrvKjHMIx1HKHZSfCgd3NAG8Qi4yIdQhOXqp1Tu0n5/CPmbJb
/1I6qft/XyVfsXdxNv0Z7R4Ib65EY2+8A+f96iLfGG2RWPILg4LBHAxnKyO6ua5K
Bk3pX5Vr220NXTK+uTEpxyjBSisEtjoZ+jGmQgpnainDoAlCyJSPuTuRCt3LsHXO
se4eS8p05c3aapzn6ESuK7gMRlgJgKgunvrs8JV+QEzrPTZpFs4RSK37tP+z11YX
Psv8w7OAjLrVc4vSwv1aAw+73sYOhcuAp5kvpcx6eXp7tipqOCFp4K63iQF5n144
F+epzo2JjZpHrrNWqt9ILGTZDhHjASXSp89yVKdB9obYQsyZ4i/2wwKIPfDt209h
q8aP8WmByHyoQ/7v9Cv8LV0zwYIjh+q6L1Yq758Q7D7ot7scgvRnb3Bawid4CjuG
/siJ+d9T40xKJ3Z/6bCsjUEUCxIMN0zc/aOwshHScDccYzKBaQgpvGb+alzGX7nW
8dGUWgqZsj6K0r7BXAZrhL+ejUHw8Y//EOtNyy9x1sqqIap/kcmz58Jd7IrHsarw
rFTJdmFhmiqWfUb7xVAAHh3z9eiSYlkwG298ceCnLeL6vbfglYeGy7tmlY6IqlTi
iufEfFZmdL0qrhoj/VmQkyJTD46m4EJxwVSw2ZrZUMRECtM6P/9qOqwBumq0jAek
toUBEdm+ACncNflAfyMjf5xoql2KUuDzC2vY9JfvqLAdlSf1YSTYvZCq6tdROwlI
Cnj+OKF5RoYbjZVumDeVoSmarX5fJFWtRuy+hWE0wCyiGdsn414l4nUZBTY3bX5K
cdRMEXOEjA8Rm6evojs9fqWlu+w3+R8IHKSP/CZcyVOasgz4W/sPmbvU1u1kwIFT
xZZQo66YvESHGDI3saW6X3GmqDhAmS9yjDQ1Ud0Vu1BQnRi/wPGwKvEaQHKkaRM1
M9uoNIE8A5ahTZQHJdz26pDCistf9gLOxBJE0joq9SS9NsH685LBBmWEfPyLL35p
HNL1ccHwOSh38BNHBIpiwT/EUf5t35iUJ+MSOZNTA89/2224EHHKZFsCRd+vrNZm
zMy18pLMNt2WT+35nk4vGV3gO1YUggCSyLxTSFsGAlXO1OPtS+j2HhnThDSODoCq
QtBfBtVAZBJBkcMDkOnkMlkrpO41O8TZ7TtlMET5qF1EA+CSURjgSZaiAEXGGOSZ
NTLdt3cf1kVYKtzTvpDN7ej+337iK2elMZ+bsW128uYW39mxpUEy98z5oKGxtwyP
A9mW8GLnT0/uYi+pIeGOJJ2vJ3y+NoEVpgRts/Cgq6LlG/2Nas7NEbnJSYmKKnau
U9E4X9Gwp17KxLrzq6f9k+SXxE+ouyiSoGFTS0il9a5OSnWlRjtsMpnDMLyILzDO
9bXaroyL9uFr5j4V46PD+gwa343iqX5+NzQ47MmzYFyUarhUcADsxrzCV18Qz8dS
MJaWECV3c76upc39/+KktR39a8VW0XaF8ssmouGqzCY5AZ5XpZnaEAz0oRxfwOj5
TgQe2zNZpdYxjEDgr+v+kDpYgGhPyRkeq3ZPSrMit9zLAKZufrf1nxxYL1sXeR9j
+IOF591pJPwREiig+kxee91ArRKGui5fi96PRQfm8kivgmKt7iDcdwT40nGHDD/Q
gx/QOgUUXcPjr9VDcV1xmDCq3HF4pcKmlztQDyXws4T1Kp8f0wma1ZtoEgjzd6SX
BcXagCKjXNPGp0Lv1KS6zz1h43X1SNzDYWjlE0cUKGERMTDIJTeKvhWQ3oP6RvzH
+Kb5re/w9BKgSXt5MXRWlw==
`pragma protect end_protected
