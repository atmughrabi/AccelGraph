// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rSTmxezLxtNWDXUwDs3jTHRPGF4xbQOfeX60xyu7zMHa0gVwSlSGOTN8k/MQ/tpi
j/BzWNbmacFc+YTRZq5p4RsKft+l8ApvRErxtR3rhs4itEe9mUdu/woUbV5iEl/x
ptMN0T08xyu4UmE0YnGv9SwXPxEDP11dTAj9WwXtY2Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8992)
cN5nm8dJ7HPky22rgnrIudiGR1yggWU22hOcTA/Ek4YBfLv8qjahTSHbNqG5lFUd
5hg47mNv7aEljGbodIXvssPKqoioJuA8Fu/4EsNrc5lMe9797z+Mickh8b/7cOr3
P/CHctcMtCvqOr2CgFOBefmKwMnjVyM/xLZaf2C4NYaLSNjdySSGtYCBBu57wvY2
LMPJcr2UfDfDQQa++cPgFXJFaDiUHsSm1YRsoxsrAkt82eslkEcqZPB+wUA00daL
5+hWMGkQs3KOInjO7Gf0dd4C+pZ+QI2NHGJ8IN1hr5Pu249cCXI9jsrxVDNLTrem
dfwjnHBDmkJQcpqhOf+FFsxpS/m23Tm23ESMwWFFMCuKDAB6fJNPPdoLft5FNd01
Uuikuh1Zj80WWuvUfdYi9vQLuewILuO7JWjnl1wOyzaKGJ/XER/90bShSvWW65Ns
Fa0v2D8d+olm4uOskFADmDSX+s5OtXqgCNIoWUPK/W5W+Lm8o7I+3UHWqIaEsoll
5eccvIOdIm0kMuAyUbI4h94wjr69V1+ebOVeVURr2lNtPh05sefFQc4im3YRdfvM
YXA9WZq4Iaw7b1JM/P5Gl/UgXo6uugDaV2IdJLmC5y0R5G1t//drRmY05AKEgkyM
3wpfwUsx2QM8cgwGGi/XY497ulc5+MG/bMVwAib7GzY7Lb2qBThyGtiHa6ruH1MP
yGhFNfRtt2eu+AGi4JKqOYhd351iGkDv5/IOCNDpZ7amEvqqKGI+XObbKfZ9ELEz
1a/WyencdyJRTMusmso5mh6W2NXsCLxOJIqihI/8LWKsmNUsmMP++ZV89rBgcxvI
qW2jvR1aoPvmLjtE8ARRVBoRwcLqWRXg9d48gjZJYaFw2KvLtsYlTUE9GBT0p3Io
Rc7+1pruOmaM4rwRTCujBpY8Nb3V7gbRhx2fre4iGh90qA/oGTHC+ds+jimwIUJC
Gec/JFcSOSf7sZwwmPenG26dd9SZ//is8XfNSgGk3CCMFiAH2G6bUA7xRvyq8L++
f8VsoVK8D/XY4kdsjtmuY4HWkp8zH80RKSoXWZCVHNFNV9Poxh2bw4aOn3CoTGkw
GzWmOiEV61YHtAvKstyz7rYqG0h8aWK0Rv1Kx4gnyfr1HaC80HHSkmzMe69cwSfL
mnn7YUGqmBVgn9yq6TILwTY4es5pb0J/uqBwHoPwuyH7vZrxBvdbNnR+zIM1N47q
sDHH1v0Hq6NoQlzyVOXwsqqHPrtHvTQHupSRQXOMCF7Q7mLY+/FewGYJoGTTKceQ
oD0cOi2xuIJP6qXFXvYpS4wrZWDrhJZqpEUMYse4E3hA0Cr7RnKijdo0a9z8Nlbp
k7sZ4G+2FE/RW3/N8mw8/c4UhxA2/bwAY8RhRtYU35Mr1tD49zv4twcekZqPAIeP
bpUNAlLnS3uFQgichxz2Rdt/pLOC8qwCyn+jUgIFe8UmBMDn8trvYQasXR3FRkfy
Pe64bgC3rNN/jtnBjsVTO2uvr5LKA832cGWySImWBi0H3+hT8+UQGcZe14s4AFFz
N6T3Ie3c25eneedagyJ1N/9V1EDfQUWduqRCcupdChJCSMYi9at2RLFOOb+aQjCr
X/HxKl0o0zMGwU8bBXUSVXNuHQLgF0pcb//x8ctBQ69P96qvD8EFXAyUL0Q4a/15
5r0Tvv+mud+zce2azCwiY3GnupJylx2wEwLq5tAD+EDx1X54AtfQDxymp8CGnsbZ
aVd6cFvOaKkT44tOcF5Wn2dlMDQ10x/Y3A54+OHNZPgT52U3eTMOhWCsTQ4m4xd/
6Ijn9oQSf000F/JWziB6qJ8epeBC+fL1bYK711x2qwjS+/00N7AkViLUfxqiIMtQ
EmmPa+sF+pi3UeMomIFWTMIP8QilnmCS+xNaBh5TvMEhlV1qDgu0VDujuaSdA0MA
qbaQtaI99r3FRi08/JKhgTdUeW7m3+Pgnl58NmLWOuUv29olL+VyjNi0w88V9gbo
CpJYy7v4OfsBmQlRcrtfPE+nDMhg6uqXsmiZRDQNhu5MStWHcMlAbPqZgOpInpMQ
/FyZupT/dg6QkgVG9jkL6+rJo3JRvV/06MCJ+lOTeNh7B8Nu1LBx5El/BE8n6dVi
qrsvQ2IXvdbEGw86RLSfffg/PFj5JtSuug3qXCF2znGtbueAoMQr4j9m0pnyrq5z
BsBxnXPsYhNDzWwlXwg4VdWFleRT8SyDtqbkvtiwVuwFomtD+Ylbnk8t+jKPvkgP
Y651jY0rFiRnlphNVZu8r9wwEo+k8Aecw/w4da2xwSVwLJmzGBcs4FvEuAoBOavF
cqgMdX3tZ/NtDPAcmF8UUiYVRFJXTU50AJMkyPicG7eA1D5Zx3Yydvyy5/XMx/pM
yF7kKkHV1xh1GzagFNsbUFuaLyyRCHZvPzYZtKVGOLvvbX/5+hHJWGKEPu3YzlCU
PpopKyCL9LXuff7IwLMxAnsGnI9y76uNq0Y6l+l3TpSzqUIBOkXCLhFs6OSJmM+N
g5VYCRlAhFq1geE1nX2/IzZx4o8ximihxqD6psFhleiA1+mACayuu3gtZXBuS2dW
kv9DGr5yH4jNq4uj1e2p28y82TriTuEeX1h4GjFKBUY1DD8oRoI62U/0CQ1IDHkC
t4ZPvEc0rRO/Rq7E1J5HjFS10vRsPhAE0RCFBEY+oNBoRV0izK73CU2C9ZH9B2tv
guCjnu+HgqH8Rr9LAbMAx5afA+bc49dGoIVnEb2x0HkOY/rhZv4rjyqq4VsTEjp8
q4g61J/vzwgg3M4RTsMmtShtdfFJPLJ5XriVVpEfqwnllectjDTdkvpRbio6j+oh
xqe8kMxLh23JjqtWI3Ae7OTlk4xojwwvHrmQ+ZoVN3njqW6KNidhONmIZbAxL116
8CKUXc9xJzQtGCeZVcwJ2qOIDHgWgiAYUrP2MGbbiPYtS37NgDUZi2JYr3jed0Cf
nkOQLfY5fQKyrWchVh/1X7X0csC2F6iDDy1m+8UeAOhxlN0yYvUHrzMw9pUk56p9
bsugTMoIV4fgyaIUB6feoWHxQkLvJFNf5lX+r7vlKXXDdS2v8RaDM2Sv+1M+LtgA
/WiqJ9KzfdRt6+DlJ3zaFhsv59JksogXk5IiQLyvt654Jle1fWDKzj81c1Ikk8sn
ZUYfh6LdqeH5m+gmOXHSlYrfMrTjcf1Dg737ty9gPg9qFY9hr90cdNBCCsq3/gZb
hnmICvG8roY83qja1aiuXLgFWIJY3Cb8/2Da+5QU+AYHjmpJ6YomnqxIisH8L/0r
sWPq2FoxQ39h/+mM3YqK7V8prNeY25K7XwKZFOny8nI8xOKbWkAHWrVmQi+HNfnZ
ozX3HrvWcfX6FmapeCBX9bR3Xw/Xq/Qw1BgjgNUxXmAF3GzTrhTDIvLDbitU/RqF
xrzjHqZB7DTVyClKwhRhKx7A5NWvOUFZx+JxbMArw11BoOBLce5a6U80nWVtueLD
LOTBdnyYHunkxJpfnLiLAZMdEC8JFQDrrnDNoooFqprdn3esRtMOVuZTfdXI0dFP
lAMcUunptDoDl4hQKn6sjcPUgCA655U4Ghc9iFAYSnwyDf+Eft4O86teKjD1Uhdb
HBHFYwO37sE/+820skHY0VAXZ8rVYq/yZhFeZBS4YZX1HnQS+8jc1XUPdUz9OTJ1
9xvC/aJbetQZmKMpNj9qBcbuj93AHjBfTxZNt97pmxoOV5ozj4azpTBm02BDwhrb
3Twpb3RWFc7mNUe4nqcm9PCltq6n1HYJL8W9KSP5HxIeS15f/f8DuOjyIE0w8Adf
6w7MAfq2gsRpz4L+WxoumcUNuxBxTcYZQyhYr1Qm+MUIaWlDedZY0HWKQjhCWZI7
YziankrWHVVDEMVEdGoaoyo1OiDOOcUCjjq1hrQkHCRASK+KPj7vNCD0qdguFI1E
7kTAJpNASK8QNQCdnx0W0cicxkhJGHXSyj3LcNaIgQc318JwhGBCASPfAroHp4NF
IlCBrJ+qt0jkizMzlW03w2PEvJr9QI6a/76d7HDrbvMhL0T6fqYNm5+jnmupLn9p
IlzQSZPfwD4amXtFO0DFJYw1ZnSr6REfojB3o8RNsi3EE8yBPu0Vj73VD6077uBU
YoGECpGmp45DrdhzooCz4vjsemv+4SJXzD1FZDctehkHvRXvJR5opAQAEazT/Z0a
fdJI0D2o2uFx/KgEwUXOxNYqGT8zPqvJt/1CJ6R7APSBO4b6PStk9wTG2A2nUbe3
/gqmMV2SUZhjGZqXG15U4hmDLXp4A5xnURlLEoMjPng+aQMiaVRDK4puNHdQ19PQ
HDAcrrvWeyOfvezATKWFLLjPX+WPHSBE2YAbpFwAttd1MZ/RDm6KYLGbfrLWH7/O
9TB/a2cHd5ikAed5ypZQff7WDsDQQDN7XLRtxHa0VPcfpJr4lx7NJLuHrih5Kr2n
pxkWNSuRNJL5MYqIdFWm+Ta1FcL1elcVdAlktcZ5ffrA9XI2AJbkDdZ7RZZ5bOgO
tF1XKDDabB819R2lAtVhY1bSL+tDwiVB2vq2Z0j+glKOwAlpq5/cEIUXlFfyOaWF
QmVD3U7gN9XkL9D2BXH5LuVNlb81B5vSEIji2WZ+U8FLFapY3+50RWgd6Xc/1jPf
bTwpe+XEKIDEFX3OZL8/8MB1t/eByckiW82YH0xoHpa78R5SYLtiN0GSqd6Gwa9E
1cn5OArBohMzh4S71upYhgnT1wTztFtnndzWOTa9GE4GlsJeK3zVLDvVhOA3c844
AFaOwIHapdrToOaphozOSBFViQanFvMzcG3OxdMBEKRNZmy99HFn8xASLlN1cLGo
LlvumHBWikDHm8leO/TCvUDBy00LJMUweA6f5eF2S6D5HGrvXLUDxEK4FPcEX9SV
SWbbfATuTj4iA7tWgswcprR7RG6Wsd2js5UeiXsyCq36XY+aZI31tbuN8/SgMMbA
qRLY9CJ4/1VSj0tP23nnu1iMBxwwKm0IJKPK0L9wz+cFOa1W43dKoXz2duIMy9vC
itgJIkVsK8G1/2s4Mw33T+AJyyKlT6PH85CAOyzkhptEMniE7DOq4X4NSK5LWu4N
3Pj+tLhCYuh7+pdjEea6fkS7GBQOuZ9teg+Y2rfYA9v73uauiHZaaSo2dNnOJizl
3IyoWqCRL2EX+o3yASNy7exUJb/Cwxzqn/sZZdk30UP8xeH0oECGBFCXQaddxGRT
z1udTIFjZpyLCtoPtKGgW0p37s30JaPc0muAM5iXABmK+GAeitXiULNtxjv0sr2Y
+8SYm5cAKptd+3HGwaojxsamS7heHWXtDgD/UBW3pre8E9+JxZwVJrwzr6FwPT/v
U7KfcLnoDPGmWCeQTnHWWiMaBu2E2TtQ6aZTYQDc5vlcAF8qK52oql1UTOcCur7c
vHH2y/s2DVeISB1+nPzRNJxeb51mxkM+E+B7lmZQS9nZnGpBDv8HgoU9U7pWmtw7
kuelrPeWFarCKc3J66X295lx8x7IuI7ySC+9uP3q0zNmdufr/akObUHkFkowbgTn
YsIpi+wLDKt3ezP5VGT0PFUtMsFM0WlsZSayGZ8k6mcmNaLsTqq9cwO8CRWbRh2H
2dtp3nLAoTM98C2V10cWId1hsBPKBUc1Pa2GZ2TZN1omBTjH0vmXoSMOlHlOge8W
V6CHOMX0FHOml/WkX3utQNVmaw7zI2tujvc9WHugjfWXqQzPgNU9K7LDIeVy1TpM
T4vUg2wwp7b/4xAsD8EYF06zIhBbQXDW6/Bpf35W46ngwslw7ffdlJuYB9mCuP/S
7MNndAQ4yoRvv5CxY0zt8zifUP6I03Z+d4oYsnr2PmXSiGVXC2gRPHy26W8Bdaxj
R9iIOHz8c21sHhlJtSf+E8MH6CaB5zo82X7opUcWdVLeNoYYLNdiCiytCnOxvMG0
LuND3thb8MLcTyt3HVVzTMrKEYNLibcc/4FkwQOCQyo3exlXYlX751wWF/urrICY
WAbzw9b6ffBwMz4ChgR0/Vcz5aEfqhnxxnFK2co+4sPJRD6a0Uak1uSLo2dxWc2J
pxm4j+gIu1DFn57ItEHLccygwYKFBVR8zwAXuREFfkLZHMBt1LC0ZvYe9Jng41W2
3vwlWw2hNOfIrwVaXX2RYCwc0ql65JBs5TMw5wCXmgcyiN+cq8Xs8VJGgbXBhmpx
T3aZWHUxf44TpapRStoaNlsm4w6yjMAcNDCsjVjZwLsTw3gmf2+qVLWvtumpD4rs
lNibHM9L6xbebb7K+hXy8cSb55Y0lnWOCwhBICe/gJx9dsfiS9eC1p5BAHUr8b3B
p00h45pugruin9b62fW/nd2FWFhYSBfejFZfZ8Xpm29ih9+furS+VxvJZ/lQb+dv
jM18bdcKzNoALeSWurC3JTnEnd3GQIdPZDbUHx3/6uhAlZ8RhzqLMxOpQdBRpMp3
7iJlpZphLtI4EMXVHQx4jKSuO0Dt8IDvxVJR+3cocj6l1PrIuYhyWwtzMnd7p5Mv
UTpz7EjzpZSeiqjBMA3CnOPk2HSSmcWE3qBWncVK+ylbiZKZoIIJ1x5zbQN74yh9
EsmEOwmqmyuA7mCoUS6HK/yy3xNNLPA7+a9jDFcdMeNFeluSob3UXZ2rwJ8ZKJ2P
WerLdGyUTD4QwdVcLvXNpjSiMxKcx9wHTBaYqx7xfIKj2bbJxysxf2iBdSXQKW4m
bOmVKmAvAENvVwb6m/LQvZoUewVfwaQ3zAQXq3i7ynXlS9i4e5i0Fh8e+iQQxr0P
D9gxlS6pwP2wrEn5cKOfytcq0xD8sLP0EPS4jqD9y8K0DDqGVF2bqVZ+oJ0YCwr0
bAKJHGpw/cgHAgLiD1+EWAhPuAmraZo9iJx3/2I7T53lzjU02oFCyM3AvWYfbPp3
rw0D6+6GvVSyKdQoMEObxra788OrZcRIICy+K+Pg1T6jPTVafk3Pi6kmHrCnFmfH
oxcw2xZQLCf6zQMVhZrrd++/h7c3eec0dw0vVZxgLJIbaevRYMNi5Jsq4WFLBN30
mulAJnJhWL/Q8UQ8IlX+lRQtU5ie5EaSbmpnSK9Eu6CtoeuI4mQw+rRqaBYcFrwL
uG17D7MYcUMOPQmrfM57BBKWngMxFDqWOrNg6u0dEG1y1Uoez+9MqQWhcBC28olx
ONgr1XrE6i7f+snZHRgdRdW+eCFC3IV7kBiSL8SmIDGox4c5wvsvMVpFlDXHxNbK
3OzTUqe2TDSfCmbnGKsvtjYqeOSxNiMhSFZa+7VX+yszwfghDGum/or8NWNp0b0Q
vzK+gc2mXU1572OSzrF6p7C4ZQQT02C2rdW/7aBdJrHn+cba8a2ZfEYgEj80GBNd
QCcLlnC8TBnHoklj4Oyv0YtjUlY2LU15DK/gnN9XUKmY9nrgTtlhauEvk3A0uoQX
1B0Ts4bLSfgDPzvvaZx66fpkyEomSWRgferzdDkjjAxli0OACBrpajmY+3wI3z6C
z4SUCBpocsNnn9G3bi1NW3FpB6oeRQAXE51apkXOXc5PyTiWloM8qUTamhzKeoqI
VZVhoo0MY84WFV0hgapZtOqSLWKAa0X4trRdhTAb9E5L3e5wvQbCfbc9ZG/2Re/7
fb3kJcNFoBkQQ+uHJI8lDs1+NP4h/ay+gwakcWff1LSnXUtc2gdf4qC4uD+UIUNc
rTNVFhGJc9hhSCmtfXuchPIdvWVtWHAgz6Y25RXpD84V5vWugCfS0JyoUGTTvD5H
jT0tJhCjtIUGInhV37TqWVKM47xZHQjfVoFn8hxK3QhHCI5E2VCx3+SORQrnHaPT
SZr6w+lNApK6i0Jqu1EY1ENlyZjYg6Jy08+qMudKib5/66YGt/5Klk8eSLrq+X77
vgFMMA99nO35DwuYD0+fNGwNqGvvFwrV2ya5+4UvXtxD1usV5FwVeibEW/K6PEYv
Wf0p+PTRr0UA6fh//Bbgu2Dq4hkl0LMVOvuepCxg1U2PgXJY3Bkrif6/yPjHUnwt
If3aBojgD8n6XNzEb/xK8sKl1KKfhMim1ybuN+YFWge8jNakKOeB7qwD1Dc2FonJ
p2aYkWu7vnlHj3otZFuqBX/UcsrKeY1sjusct6XhXQZRQChA5EWvAbqQbuNODLM0
BDbL/aAmIChKhZm/6UrqyZvNJS0igx/r4TmrNgJdit/AmFqOVTHj7EtLCNBhQhRa
NASIBH19+EnIrQIUu65dJB3fO77qONjyptMSo0Q4arg1bM69HRQNxowXcY+h5zCR
2sxZZvnNRGpm2umECtjWKTKDg46MGziH0Ivam+r82/M8Cghi2JAcWxa1yXK495Yd
KZlZKPjWePpkXab9tPwTScPWgW12hbIcO+PPqkxHdW9JE08fdHOWukEpQSy29FO5
Z7nDl8al8+VPx2ddLwWWse8e8tlSrRHqAEiqJ9kqW4/me+JEVbWmRE0xSRmKZUlw
QQltNZ3YnHaqu+CqUbS86fUlP2Fhr8o4OwV3YXVcDNjL4bJ3EuCOTOJfclqUK10r
NgFdqT3Erf/ShTYw0Hz0t4jhE2kXKfFXbrv1FvVV1eo4OtNN3n4fakQxv9+98fs8
qoXQFV87a3PnA8yQACkNtM9iX4+LlA1terPpEGH0/H8zv2hpeccStHicu741MHHf
JaZeg4l+r4vDitNS4+IZRO20HY+BQ8RbSRyIpPcrQpknAmRG5iSIo2+pgh+26PIB
AwOhI4isorcTHA/nsuZqWzmlavvBdE1/PneLmqJBh1KAfS67vvLQ6aIq0Yalv1SZ
MpdvUINl6fkPzySUwm4VlOKwGGv0PV5lpugcNU0Il4WIYDFP6j4oEgRvqolRnQe8
4xkNXQFVD+ks97p9QLG5BvZnrYIctjgymKnQjhDw61znMnjOPgLxSfop8X18ilc7
eVFfSvorRUZHz63b7dBFIEYXh8jJ5xAHAba9seC6kmcy7kwPQ3usUN/440J5piKa
X69nUoVZeVsrwUDZhyy2GFbVik3CdaIZFhU6kT418cM5zu4NgYLI26PbIwnnO6h9
/ikZVp/x/vzDOeqhhx6jNMImg39W5sTwfm3jWYLlMBCzckghOTz3VZ9Imji+KwC+
SzvSFQoWZBjfleRG3p3MuCYfmcJpoBFBqkorNdjQqFwo38dWcBm4ZUKRKWv127PF
CrfQRXxlClL7oBiQcf3VQIRDX2stLQ9oYnEgswWiGJYgTqLdL8qtmS7VAfpA/1Um
HI4ItIkPRyIY+woInVZr14yJSi8JlW1/HmXrqIXBOWryvYWcdNPZWCHTFSwbnfRe
wIoAuvpJscZz41e0m5cUTPLx/WVsLQv6wRYdKE2UzybRU+Tt++OQxnp1ccG+RbKr
a7Mxn2HHOg0xVBXbGLAibH3WC9MlU4zo4UXEEYisChfGABYCKgzJQQnJxwcE+XuQ
S0W/J0XqI3Yvzyt5m/gYBHCyr6vy/gzyPa2XCUukf5Ji6kO14a4YG61G7yY+sWrK
qMXzW4HRdSUgwum4q8Zn3bSG0/vUkgdTZirPrOwv67FWdzus5K/jOaopdZj/cAuu
4NfEOU/I1SPw41PeZlFgZv2aF6eLjuoUnTiyvptC9sVUpUnyBBqgu9UH1DnOCvOv
pycCKD280fHXcl4gDfVoffh7i7Dy3C6i1bvxILuQSW6gUpD+dUF6KeyXiLeLiEmK
W5tEiNAnVitDDT9trhvfG4IhPLYasS5uCedrPlrP2BrxOqO/avzlN8s/LLsLroxe
igaYhabqks7gU+Sk+wGq22u9CJULVBWM0/AB08GG5f3Dzkl3iPqiVok5UC+GCHIt
861nkVvAfekRBgbWgT9RrxyBPjmWzDdeTJNyiGQq0uS6B3nL1KnQZ0ZIPl73uyCw
q9TRof3qVxyPw4IRY0GBTD98W9W/HUaphkFyww6ZZ90FTbxgu8acwJxocrUOAThK
jjvvF9hfRC+Vo0OkqGMfchtKCMxW5EyzCgWGGSv4calPwHJR2OnjWBYPEbHpNB80
pdgSXCX+hkSguWIbFdHChMvGWuYBFVV3y1wjnu7I/oolroyCIVepJQP6kdyd1RWp
PwaXLWJ635AV2l+bxBXnSeM+56C7K3NAhHRzjO36+OYf5Mm2zD3HFx/nijldJmfr
HhTgsNRuaQ1G+xxhQyrZ7FpTf5WEIOU7SmJVvuvwlsFMg99dMflXeVCPErhx2noM
apyHJ0akSFv6VBvykxsiABs0Xp+HG6XbQc325Bwx81NWNVvjbCpIgqBddMD+U6Ni
eTToC5MEbOuZcQ0+UqsJWQ0IYIOdaj3QPneU2mtEunu2mn2OB+N4S76k4wPOlULg
mAWwY0swQUGAV9JAvEHH94KTd4nKgmKzHUOcd58kD4CV1kTTejmHROb79lW7hGwK
sIFcJ4XnsBex0pIrAy84HCoYtgbAlx1HSvC8S8Jaq4vt735XoQT4G6cthxGdnL+v
+J95GWvYAZg4TMZ/+PO7e5ynqqVEjjJX7BNQ3D8MhnPjvpj4VMchpWGTHfvwShQj
A0gm2gAt+zYa2JoHN2lvxi8ZrOsqVlmlORjn/uiOIJaDfC4aVrtVv8QAsY+vC7XM
Uz5O3Ub3uOcxcfBDkh3ZEArWOwj6QCuBnpgXqeDe33+SeEqEUgAXViGMnxD/ym7G
3o/L81OZp3gLScwP//B5xRS9Nr78nOahAEfgh0IJJ/7PM2d5gFo81e/7GPTKyG3O
7I8RKBfgkybd6ZKkBeMS2ymoszDBpxQUgCw2e003K9BKZazbOH8DgQJ1n5ivxCDY
l1hWVmQE+Y6x6JjrBpYWn1gCSezrJlnHrN40zRNOceqQ3uMrtNDLEAtspRdkrrQ8
pJaNLFmDU5xrqbFrXIiT8X/zASMQ/AW5q1q8e+NMwdXHWNkNoUfr1LbAeIcEpy9h
lv3VgRXYZEP2/rRxdHe3JhwXtdvjoQFZQcgzyfdY3K7QI2gMS1T/BySsIFk5BIKQ
ii9EuxKjWMGHSkTXSQcbAL4CsYRfpo6GYAF20H9QHZhdEFODLvrD1lBRuYBsHvP5
5XWmo5VSDgtPX3vdgjK1Zz1Oh6vs+DU2GAYXHLTk2D7ayHJCgL0fmF5bTwOLbO7s
Qi6NkKOuMstJEcGeoeTd0Q7exPS60WJFpRqmYmLRksbk3wv0n+xnn/6qc1f25bsM
Nl5KzXDCTq5Y7ikSWTWkNpFKm8lwhqK/YInNHproG808BUQekIffGr2U+ivj/LuK
Fu4Nlrbl4CDZEDHVtft+O1ctvuKRPr6+BLSzW2CKQ4qsIeY/Y6eEbQCbo9MBo3aR
s5wr+Sr7X2GKUxflk0ooBOGBOY3L3nB40zwlzM9T1wnotYnFENsF8Rl/7c77SSl9
3sO+pDGW/GOT1IRX1UzQPnfVqIjXf7yizsvzH4z+nuzhX+ES/o/VBi3rqa7KICxw
iEsWS/N71f4o0AzazEVvTxByxxCSOtmHUbGxbWdIc2BY+OUkCpMVzJnJb1H38Pk/
Lmjpxa1ePD+woBU5GeJnYZu96zgVOL8yzsLIMlqHf7Zl+3EY57mT5AeUsDmRKVOC
Mj/1+wt9vRsJhnFcnarTAfsbBnY7KiTW5l1D4SYmbcqRgvApjkTxY1KKF4p+ZgHK
I8vsba35nmFQOkV4npV2MbylVJhmhJuHyAxh2VdosbIOV0EZ2jIiNicPJjd5xJMc
+lXNJgAyXPoilkbrt2f/n9f4xeVd4Nru/OcuTBziiFnkr8waNNs4B1LHA/6ypEf5
IEkkHKR7juYRzD94KM6dyeLnn/IqCbJPrYp6mrfhmdtZyqF7SWGl0MwjXl7Os0/2
DhkiAKgFB9Uxo4cAoHMxfkG/XzjhgKROhv1bwkcTUEOn9a7t9MItiPAbQ0WLzBYp
eG5MydZliCz+WO/ARH9M3dJDk9vVUPIeb7TeIsI8sGSgKxCT2gye4WUAOBxj2ocS
efo+jdheJd5FzyKuZj0E1OucmPDrkxWqF8TaYQUv1vRu/Z6OYkHqRJU53aV+HvoC
4XrhDxlljthdzWi2NcuMfffdUcfR/dK1tIdu/CVxpmaBT8SKn45GNU5DF02qsz4y
cPy0o7Bm3X0of/euI8sr1w==
`pragma protect end_protected
