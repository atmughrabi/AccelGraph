��/  �Wu�ٽ�;�G*�󤐛^f'R��?_�k@F�N��@¹�:���E���zٽ��
����p͐r�+"��b�*��eN��|ԝ�����|!�pKK0��u����Y�G��U�$3�:
������!���:혍6�7�w���ANkǰZ�UOc���Kl���Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9�㑝ckh�^9.���_�4�dt ���o�Q:!�l�͊���=S�J�8�{�̷�ܗ���X�5Z�S�AD�:��-U� ��,��U����i�
	7���}6�͜�ֈ.ߺ�^ %��F�M0�*�G�e��X�k�~Υ��
�ԖK;
�uV:�1׷�b��d�Y���o���x9�^.���Q�A��6��(ev�����F2�u�%S����zU)�I*ъ�@,��Vʣ�(���|�8��Uk@\��V{�s���Ɂ�j�n�����/�ـf�չc5g#_�-rⅻ$��Noj/ �_���	��`T�:z�-f$B�o�6�|��1����W�{.9�Gv�}q��l�Ǯ��d�ƻxd����i��sa(ܻ�����(b���-m�jJ�J'�}0I\$`].|(�P:���ظ�1��I*�O����Lm*D��ո��p�����fd˅�D����n�%��v�-�r^#h�"���M�D��p�픭~�7�躍��%�P>9,;(��>���$�;Wv�&u/�0.�mV��=��nM��T.
q�@�eFh��Q ��&+bo�*�춎�uJ�+�#Z�=Gί�o`�P��^ᾤ�i�v���|�����F���0v���tN
0�Ӷ�.���=�AD��Z��Zq6��,��Z�!s�UT�m��U2��נ��y�P����ټ��~u,7�"��T�$Vt���q���m:�� �vH�4�0y�<��E���v�5*��	58"�P)dR��=�pC y�Qw�y��3H�����&*RT� �!�']*k��t��^��UV�����Ϋ����B{����"}�D����x���^<���b�7I�%W}j�Qq9M���.��Yn���l�����ҭ`1?��83������-��*�Jm�)���?�hHu��I�jܠ�A.�.�5p�^�C"�������s��9����g;�$��+���4=pD��F����|k���ύ�
�:�@H��`�NJ�Y�^G�jgd�Ot��.�x��2�b8ˍG���a��nu�a$A�d�j9Isw��T˓ydJ#'�_�F�6��g�!����vǾ+�Ў���՞�gI�uK��l'�i˶�G@��?��Y�DH�q�p���|���_>藱��dte�D4O�H�u�[NmD��(Hy�]X:�ySbߙ���UY��S�g J;�4���Gt���9*ԟZV���@��������Sf%�;��m~�ol
�심��"�-ڶe>�0�҅i��΄!խ����g`�N�K.:�*H	�f�%�#h�m�N����i��DM��_��z1���)��u���{
���EuXu�MP�n��m��a���M���/\�.����5����[ީ�� ).+�����d���S0�aY;�#"�N$Zu���IA�4ѭ�Ƣ�Pa��R���Wy�e�X��0w&��0W�����+�q/�t$��/�~i����K���u@'�Z���k� �����=/I���#AW9X<��y���5O7�z��M�u�K�є��ǂg�����_,��,{p4@ZQn�Q�m	�%l���3~i��H����W���}C�Қ���Zl��z�(�A��.x�5JG�hw �xK�LY~AI6�׹7�;��A�����;�s?�Mr|nk�Q�h�-'�D�an��3�X��|¾z'�\:nϪ��"0���|"+�S��)� ��9U$&�)�����h�^�X�u%�wÇ�#����2q���֯�>I��>	��;�o�3RP��E_r���$Y�V������k�WO�RQ��[�^rx�����j�A�B�*J.�N�f��ǰx��#��h�3w�M���V�"�&���O�H��r��2�Ma15��7��n����G̦���qs3��闄������|���	aw���:�]xK�Oo0�7d�u���[>�OFƥ��T|��*�9׽C�����b�Pk�;ɤ�ڜ�1 芃��'���År�V�s�+dC4\+f��
�x�*`wO���I��I��#.�V��R���IhCb����Ϯ'U����HB����h˥J������c��bl��*
��h6�����X9�����|����W�m�.�Ng���$�<^%�Vۯ�^�4�&~[�D��bC�=��G*�bߖ�(�k��������^p�q���#�,��R��so`R ���97ʈ�?��8?���Ih&0����v��w�n�0l��/��8�Q���>a�!7���<��@�k�΂�g�9m����Y�y��7ի��Q���
�S�BQ[�K?%9eWJrz��0u�yL@��P�)*N?9a���X���"�Fm��D�|��J��#%|"pQ��S���Br�n�&�8��чm
��:�Q���.���~@u5o���q y� ��87(����b�(+K����D7��%�kGc�yP�h�_�8�s���4X��<�s�G(�~���QT���ISu}�i԰7�-uc��wi�
?��l���34TuÑ�K�$H�@���FG��%
���}����2���5�����+G�`��T��ԚQEDO�����d-X�,$-��` �;�e#��Iƴ��bC��Ɵ_q��p��z>�§��?��kB*�5��IBI,t�� /pN�J���䊭
�O`��A�p�zB
G$��nk�$_L�%RI��u(�Y�)P��\7���4�,� ������$� Y�v�#.��)�3��p�i#Ac#˟�/ũD�ء�J��V�ۃo�3���ЕOe L�/|�ھ����E��AGj��X�pD/wy&��Tw[�SG(�v(k�ƕ���b�	�Z�����G�}v����H
*��𹵜*��n,��Ia��V��.;��9�Aktv���5��u.��uq�:�YA��BzL���- /��O�2E��������z�E+:�V��C�8yZ�[[lX�Tc��@z@2�S�BH6�2h�Q�t䪏*��G'�m,����4sedX�s*��{��q%q�l�����o��������Xn;$f��u�G����6��Tqx:#��2�C+��`з��)��Ӕ�0<�IND;
���Em�ƈC"���jʲ!.�E�h�a�i����&O�
M���pXz������z��R�|��Vt;���Bʑ�N	���j@-I7�����GC�P�tI�NmǴ�Jo�|�d�k,���@Yq|4 �'�*Y�a���&u`�P9�V#�'�"�l�ں����`�Κ��h:=��m��+��]���x^���b�<Vt�Mo��{���$t�Eҋ���FU�O�mS%7�����3���~0XN�A���PK��IO0X����n:�@��ג��خd��H�s@�MG�N���A�����{��I(�l�}��=-c��U$���@o��\�X�h�0�.S'z�P�OQ�"\AS�X��R��o�B�	kl��[�.�va1�'q�A/@;m�