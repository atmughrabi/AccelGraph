��/  �c�9��߮�,ZLq'��Gq,&4)�hm�1˞#-�hb���~A�]�|���d�g_
S��t�(�����1�q�%\��nBj#ؙ\*u/�)!K$�T��P���&=zj�p�l���J��]\�i̠h�":x�1�?7[
��"����͂9߀�����5\hOwɞ��O�n�Z�h�Y�B+i�٩M���y'�>���X��Z��Ƒ.���^��^j56�u��]�q�|�C�cL�py`,L���eDi�ܨ���=ܑ�uH�{���I�;�S_��(�+C�l8q�����~r�Y��N�h�#=�9�+L!��Ve�!��$�^�f'����vX���&��)������� =��j��ۢ՗w��T�z�t�(��L��y��̇{F%���$�!Oɬ ���oP���-~==�enu �ȎH���^t�+٘�1���f�J���/v����X�����뚪�MS^���P-h �=h4*Tv�Y]kj�>U��E� K^�L9b��:2{Hf�a�<r���^u9�W��i��Au�#a�|���5i�+92�A��M�2h����������96�R��"�$U�Ε�ܭ$��I���$���.�Ü �Bj�@ F_D�'�m���d ڮ=I$���@C���D+�r/�h��f�%<2 2��́�e���lbQ�(ʕB<����d�C���SC����>ȯ��Q�|i�G�<3=�j�{���4��s !v!�|�o����/�`{ee���ߊ8!��c`�g��]'�}�"��Z_x���pǟ�/C��h:��nJ ������E8	�xອ㲚��� �<8�C�ݞgA/�
X��L�W^�:�����܁��z��~��w̫�T��߼䴆p�?�{_j=�����)v|�"�X&����V��+�&؍סV����a$���^?z
!n	ޓF\�I���+[�dB90�[	�X�lgnBj�~�(�Q{�{���a�g�}�=������p���m����_#�J��X��7YYwR�Yk��)�B�����g���|�[����%�Ƚ@5�m�X���v�����n��'qÔL������/ *}ܙ�Bk\�5�JpS�2o�6�����$�o]�U��V>��#p�T@J�k,.X��*���J�E��8K�:�4��"S�F�S�[�w�r�N���
;�<���!Mǹ�3�� g7�8��e㺊;.P^ӓYD�(Kje���Gқ�s��3�.bF'���kǱ�U�x��y�R� �ܫ �X~
 x�Q��E!a-�_b��THO7Oxޑ�9:ֻ�ii���$�WOQ�� ;�{�m~]���= y��i�$b�B�=M���ᶥbJ����H}�}W>��|>��1�0�U#P��*���W	�*CZ���9�h��G�� ��^��p��o��b�UU��
hz�t{sx��t4qs����m������(��9�X�'��ʨG1���L��+�G$��ν>id쭆���Ϻ�n؇��jj VbK�?�N��[�Wr�a�hDX�9�<\���!a�����v���*�0j���·�N./�p>���i�B�i�&��2��DѮ{�[�͡8��?�H���y������2����Q#�s���櫁0�u	����i��J~yi��⳯<!�uk�v$�Z��y�b�a؝���&;��.x��TE6��/�O5�6'%�8��d�.�Kd����x]R �*^�I:34�)�G~G��A¤�H�A��xv�÷:Xr\�%"M��C�ˠE����'wm�<�b -�mv�bu���%��&	�c"�y�]��G�3@m��2�GFC�ц���~l7x �ͥl|n����SH�V� �b�Q9^cC��;��oQ�;�&�Т����{����r�ޗq�W
n�Qͤ�*.&�n����ݖ^��i"��iLa������(�	6�����v�?4�[A�O	O�-kNڪ�	K�*j�D�O�g���wZ�E������rf��.`�rp:�-P��K���O�%:�͍��+>�A�L��@�Y7�a�"��g�d�-\�췎�|oI�m(��ښ'x7W��"�T\C�Ͱ�]�骇��*�L76Z�X��������tl��`-6| F��=�(> �t���L��J�#�'���/u�����K�]�x�|H��U�e�]k�H��Y�)���fT/7�����W����A�X`ǔ ��y\f��M��|���٧����|��Z��ƒy�*��T���p �,�Cm����eׂ���Ɣ`S���%�ߎ���Ypy^E:v#���S��tA��������Aq:�=ys�x�v��FOm�8�7��-�h���c��_�hQ�U斧�Vl-�Y]3��\�r���w���J�k�J#i`�D�@�}@}Lh�t�"�}^9�j|*{>|Ӳ� 鄿/�"�S˃��}�����i�h�9&8�N` ����-P��/��`�<�q�3��`��X�j��SD�����p-�OcK���
Z����{x^O��5�vc>ڂ��	���Ic���O�'��*5�J3�kͧ�G&ʑ���/��s�V��6�X7�G�&�`pA�Ѩ��v[.ߕ�eL���	���q�]��=�֠�.�&�#�A+�/d�m�ɂ:s�Gԭ޽��vfU
}���&�2��]����d�)N����P�I3�4+'SZ��yQ��_[x/�<��Aep�E~��ڠ7X�`��Um����*��%�c�Z]�DH�OY	w1��k� ��H�86�p��[��Bb���D�T��oɕ`��5W֚���Q7l�&��v^IbÖ����=���x�6��q��"��)[W� ,E�h���9��L�84��_�0��}�tF=�pZ�C4k����kC���OZ[�a]��*J
�b�{�|��G��v�4cQ�/D��ޏT�9r�|��H�g���jzXC���O�s� �Ŕ�a�̾���tu��<-�vŒm*�˂T|�@�(�|,�|����ͦYn�y�^}b�:����M�n�-�;�N��Y����ď�Pw�y��s3t���s�DG��rP����cL�ܟT�]�D;������#嶌vr�f(��ӷ��{I]�Y�������W�[�����9P��Ȉ	�� >_Z�-�+�] �:t�f�.�į+�Vsz:�(�Pe5:qט|S͍�5&�C�P8"�r�S�L�ݿĻԐ�D�#�����ae1������Vl��m��y��
�(�\��ZH�0.�
�ݞ�����D�®L�`���>4�K�0%������
���@�GJ��2�Hf�=_%��>���&�����(נ:�PH'�!^3���<�D�`r~>Ϳ�fuc;KT@6/�%<
�Ɍ)��༅3\L!��v��[�gI���1�q9�F��i�5���T�6]�݋�)R�ξ��׀?ݏ�?�"�&ڈƯٯk�-�]�sC��_R��E��9^BCn�{5V��1z��vߛ��`�*K`G����B���/U�����j�R�/�:jK5�ǲ�hp
8qЪ 2�1<r����``E�*���H@c������YfŬ�X�Eg��;�>⋾i�<��_��|BB��jOyƷ;�����ٷR�~AGu��@U~�����Fuw�w����@��i$h���$<K�?O���-�J=�]��+;BJ�g�,9�$SڠӉ�#A�����' �x,J�Nvt;:`�	x4W1Î�(9QV�c��,�v�2�6���[�H�^9k��q�� �q�N�1�-p?e2E�Otg��}��'A�o�${iY��ZdSRfr�G��O��L�L=ӊRa���^����O�ۭ�k�C���[�q}�'�/^y�iL�N�q߶f��f-{��vr&hn��c��z����nUZ纫�s�����
ݬ���@��;xz!���!��%{���7J�MZU����M��6\�候����Ԯc�jw0�Xa��½4��e�v�6��>�^���C��A�2ք&QDx�\/����^A����E���l�r�;�b����Y�u�����H3Mq�G�����!�PgǱ�LPpPG$�{9�$=հׯ�ш.�
y�����6$�%�h66¶���Y��a��E;(�QB��FZ��J�_���c�@�ə��{�q7���$r��:�k�.��p�#=4p-�tAip�?w ��bqxj��#�����1(�P
u���ߣek��A�yy( ��ˑH[q<�6,N^�sX�����b��7��o- RO�\.ʵ��O�mJ��+�4�[�6\r�۟	$���~�'Ƭ0�G�A8���J"i Ǆ��O���I1�F�[��eH`�P�H-�y��+1�D���1��䠒�/AJ`��2kj�c%���>�X�����](��?DW��R4 �0f|2�+e�r��i~\ue<�����L�C�B�y4fGP���ܴY@�C��e@Ll��@n8�KY�x�!���.L�����\'g��\������.n(�fy1g
,�$2�������m��Gh�eK����8�u��ibm��}�[�;�C Uf�ʷ�k�������2�}��;�)t>ݦ)�!��韬�&ϒ1�7��Ata�jq��5��+�/-Wဢ�^Qҥ��%v��=��G3��5=�,���rf��)�R�D=����W��e�%ķ��_��$�����Ksd��Ќ�
5I
=������F��`�"���[����b�I|�����M�*_:3���@m����P�{-ي�D|�X/MC�	zv1��i�|$\X�ޤ2�\�/��L��z�-�Կ��r@���1�D���Ӂ{�-NBJ�-�CPh��)P�K�[�z�+���Y���^� R��]�� R�������O&a�oP.ʧ�D���9��z�**�䮵A������b~� 0%AMG��E��H�/o�Si���i�3'�xq=�V .䤑���	 f������;D��&�J�q��k_SЋ8
5�b�FBϖ���XDKΓ��i��Q����2�E/�?�B{~�O;��YZ��[�G �gC(�vny`��� ��>.�^jX�	�㇆L�4S��=��c���K��]&�ט�B�5�����z�f��Y-��(;mv*p�_Y��
$��>��	L*����Z��\�ڒh�y���-�t�����}�z��9qA�6��:+[�	�52��� t����̌Jj�������x���#���7�vz΢/�S��?�Pa����Cd���45�qf����#����X�J0�"��9~~�g7	s��o�+4IÉ'`�:׽�<��Y�ʈi�Su�(P������tyWt�.uRd��!���9������[��ˡo(b�ou�:���YI�ek�h�{�Ĭ��N�ß������8�� ��7�!���+��m���5���5a��|:4�Y��k�;?�b�{L��*eC��Ct�ϚJɌ]�����ۉ�lG�m-����f ��K�{��PYA�l.,n��ƋN��*9IP�\�6�~�@"�5p��I�N��q��阍��>�Z�Ҧ�͝_��'��ld;!�q~��i!ܡ���DC\@�ˤ>�u[��.��ˌ�ZÊa�b��b��� )~��=���!��_�1u� �`�6�#"f!����r��S��:�<�]�O��6�eC�ռ�BiC�������?���g�2�ה7�$�7S34�ާ�_R�^�w,:,����l�ܣٹ ��f4���o�֛������u��|�F���J{�,r�u8�#���}�q�e�u�U��1F�0� �>q&\���٩��h��c]h���O�)J-p�R�55�,-E�� ��'�3Z�.hk����d��K�ɍ��Q�_PHl�@7�U"�~��n>D�H7���1�]�I�Y=i�`rM�����WE43�_<5K�u��>�2k�[�� ����xD�����7#J�"RBX&g�wݷa����.�9���/���(�!��r����݊� ���Z�=pE�n�k,��n���P{>���7j@��|����Gl��`��Iգ�$��5�+��k��P��>����f���5?Ȑ�7B����K����EX�[��Oq]7ii9g,g/�I�/S2��]�vT� #�2�3��ڧ[�\C�9i�ı̯���A��=��_R��"@dq������
Y����VG�_{@2\��k����
�Z��]�:�ѤRU5�R7�3�������lc��3�CCkԫ�g��a7��RG~<���P�Z��K������]5{̺5Ȉ� %�����Ɏ�p�F���~��:�#M�8Pd��d�bAN��V�_�H���&g�����F	��t�=bHa���w��]��y�����*,p�?5s>�O��&q�/@n>E�ۇ�`��t.ͻ��>`Ӆ��h7ή'��S����7`-���9���[��۪ ��FAb�w(�`G�U-��>�F'�����w�<	�D�}�KҪ��d�?�	O��t�8;C�E}T�/k
oG:2�Ěa�j�/�>�}��~��i^[��zu��&��%�6��4?����qk�i�iS�g����q�|�1�>�ɡ"��&�-��5�j��k��`�	���,Rk�;�)��6�r�9f�:m���i �S@����=A�0��ǉ�6���|u@�!@�!���
.�mQ��\	K���-��ܿM%��w/UԡP��0Ņ�60S3W�B�
��)�a�?E�a�ߠ�m=���%��7J̞�~w�<�A�O��[���Ҥ
�X�9�ɝaN��<ʹ�<S��sG�����
hl�!^qSY�3;����+�n;IK��m�Oa�֡���<&-�o�qCmqx%NL�]��S�ro+��2�<kKI�=��M�F)n
�X����D�2e�_���v,����D��q�iVf�`����lɅ=�>ff�GY�w��T(�k��*4b�H�F]W�;Xr�UR��R׷�B)v�C�Y�7�>J�!'!ON��f�U�� rE>���"+c��ma����cE+���R��&T��l�dH�mO�7lǣ�54��P�P�.�|.��f���L�L����h�U�c�Ze#��M�T�ӝ�cT{D�f�<���L��ݝC!�E���Ī��N�|������܇�wy�#s��m9��E��a�m?���.] <�w^+�,�9�����԰�/&]��QN���S����I��,���#:hN蛑R�cZvB+ki�n��q���ѕ��b���Ղ��?�4�����O�l�5�x�L�����o��ᅍ�ɡd����a\���'-���;���� l�z<ҋ��X���cJ�Gi����j�*�U�(�����}�1el@,�D� +��Xz!���<a;�K�	��?�D��A�6uՓqZ��O2c��jZ��c�~�Z8�y��  ���,T�����(���Yl.@��n\�ʢm���4HA��z��U��B�Bx��� ٩/��.�5u�¹�AMQ���r��2_-���ƛ����G���p�`x���^���d���p#�*��� ���J��[��ԉ{C�)���#TK�MJ�N�qvt��7��s�OXH�E���#|p�����%8\fQ��C��ϡ[D��'vv�O�nks�~�\��F*��}���eA�k����K��r�m1 $Q6��9�T ��Ǆm�	$��s�Fy���̰��lqm�L8Ä��U{������ȧZ�Wɢ,����j�ś]�'�s��R�
�p9��&�w���n��gVk�I1�����
^�1V<k0lnK.����s����������"w�g��9�뾓k�s���N�?���6�'��g=���҉]��H������Maa�G����k�2A���T����@B1��Д1�����CysO����8X����>y�&��A�<�\2�]~{R��ߣ=CvX���	�,�~�!���jű֓'p��f�Ze&���gb��Y�����ր��X@�W]�CaGZ�WHS��ֿ*mA����)E"A��69I���=B8~\�wG���Y:,B����ru��7�L���#��̔5�ԣ�5�"5(�2�ȓ�����9A��\�	W�$r���p�:�3'�n�G�d�'92x����I�+��e��+�W�y�Y��ٔ�����%�I�:4��s�?��x���R=���δ0��t���!�N����n��G�m�{v,T�U�0�-��7�Ń�����Aw���$��<Ժ��8ڠ-��N�8vp'`8��(6ԢB1d�)x��*+�X���ցBzv�4j�����}l��'^���5��ϋ�];%���?:�%��sr]I��dߺi-RuS�a��h|(M2#Z��i	�_H��f:�<�����F)��s$-ޛLNW�aj�,������sm�0/�o�C�,���*&��ýݵF�r��?c����� kՅe)� �sF�2����~}jo� ���J����%.2�O�e��ə!ʫ���xiuZ�}�D��\ݎ�p��h[�Yi8�G���e�o�^m �Q�6�����)���ѥ�IU��`E���΢�#���Pd��;�d�	�R���(}�>/�� ��׹��w9�C`bc�@���Qh_g�#~�&�_�k}�:�s��%w�n�{Mͱ@Վ&.��HosF�D�'a<��,l�?�󇼃��N�&I��U�_��YP6<���1,Q����0�Rb�n\X��m�4�N�3��V̨wP�Ұ��+�k<�^i�o6n5�e) �	�����3,<s��^E�'�-l�1���9к���&b5��
��P��J��cw�#ٯ���2�I{H=�̼��Κk(	�W��jhH����u�`b�h�V072��T�'��1�J�袑5��3���Fd�%o�Dc��̓ɜai<�V�e���,迋�r�`�=I̚���[ks7�Nb��Ї��R��Z�#)�z� +u=�(A:�qn��%�Y�^e��B���`��I��M�	]�h=/Z���3~�C�����xҘ�<;���vD\cx��ȉP�����4R⃊��GY15��E�^#���>�i��>@?��ۣ��y�E^���ݶ�*�C5�Ɵ��݈���}�+����C��ЕEҔ��Zg�
���������%�i�\Bz)��70{�����WD�St���7{!���+���C��qp�;������)�Ѻ�)��F�NOK�	���z��	�4Y��|��I�Y�3x9а��#����fo����S�����O���;�6�����8��!� [u�l�4�27��O�D����U���+c��@�I|dk͊�YTw�)��ߚh�b�
P��PG�F+I�7ݑ�}�k���@��#ֲIK�7�'؛dO��\ݘ
��S�
��o�����-�@�&��'��0�S	v+�C��"[rT`�{ ���Z��X�Db��C�&W�	:;8Ш�$"�	]_��#�l����^�U�'3�T"�_ɰ�v���:1�t}T[?Qox����	�zS����� ��xZd�=�.�2<�����|��>��{@��jcəK�dNu{��c}`�}�q?�#o�g˫[�y��!���BU�i�Tnׁ��f�w-n��0�U�o�*;_�<���!Y�ZA:����"���93]c����c�g�t��I��������'�7a�g�湗�)<{\t.q�
 ݇Kw�M�y�� �QO<�sb7��AG�����&n�w�m� �ȟc�E���{#n���J	�� *�� !�4��b�F
b&�p�h��U�,,q���;9��j.O����x��(AŹ@�W��$�{W,u�#�|�4�1br�(ys�U�%����h{�$s���q$j�����=tģ��ȭ31`��b�1U�$1*~�M�����2�Z��2��%P��K�Տ�43�R�T�o?u6���u��2�jeq��r�j����J��;��9l��,��X��8�	�z�V����ܹ���(��R��t7O��;֋�rEY��G̜����
Znc�)��y��M�L੿�n#~&���.���O�Á�x���UY,❚�w���e-���	p�O{�� ��XL����nK��d��o��Z��#�(u% �0�X�����v~K�P�|2׍>�Y4�D$I6[w� �Q<�I,ՙ��7� JR�#l��s5R��6��dPSXlג0ʔ��e7c��s6U5ꥒ�)ɟi�nM�<�S���򱿚�F8��"��"3}�(�܌)���bWթ--^�nD�?��`����jE"��!�A�W���+�Z���G��}k��:�~l�G��T*�=e!A�Ѣ�i�$nг ���Ϭ��dw�J�w�|���q���IkN�W^k�z U+�=�V�:K� �z�ҩx����Q���Gc�fz�Bo�$t<=�A$����4[��6����F��#��s�MG{沓�\|�llK���'sD�*�
�G|j�H�$n�5����|[o�U� n�1d�t�|����q|��s�s�a� �Ӳ���sgȕc��>�i�`pa�d�1�Ulw��>n�hϥ͞�v��Ԟ����\�V����7�q{�� &��ZFa�H�5���?� 	߳V�J�Rj�8�	�fu	s �&��h�Nf[���%������UF	,���N١��6! +�C��`;'nO����dd(A�J!*e�A4��',��/몲w�����Zn�����+%a*�����:?��vܼ" ��m�Y|�`�B�_�B�����K=
�-⩵�6b��F�
,�Z%㰉�p�i���'
��.�p��.ĳ]���7��N�Ujph�5�BNq<����Ů�1箰���	��}�&�3Bv��1�"���c��#1�3@�ɓ-�O���~��s�0�O�}G2}��J
��c�Z�dZ�T���˕�h�,��)���֡�~�6]�[MN>� }� N�(���\Z��}��k^�L3i�>f�^W���v�N�����F���`�P�\ĩ<Z��!F$b��2��h���s
]m4ί|<����+?(?�m�R�b�ɀO��{�����gՁ#.�R÷�%����i���� I�UL��p�01>�
����\��htx��D�����ن����kuS�л�z�E ��q��/	�aX��@ZVd��u<�b��N�Lx>�\r��0�p]P/~��*�ŹB�����n�oC ���,�	�q�T�e[���x�z�ё���M	�0���s�6-����So�h|��[���Ǽ��g���5/��=��d7��N���h�x��c�A�2'A:�`U��U#Z�J�XI�Gݼ��b}���fO�^�/s�l�o��BؤP{K���k�W�/��2s֥�k� �l�ewYz��V���Ƚ��Wʞ�OB��A"���y�c<i��e ���h��*Q��	�zXcL�A�`G�Թ3r�a�{�K���`/���:����>ɭ�i�8Q�b�A ?�`�K.�ut�x����]�I���v���K�]2��{G��#T��O�ԉp����b�v������G�{P���l�xq%O���2�xʍ/��u�>fRt�Έ��j�V��2N�m4k;2\�9Y��|V��\n���Iڪ�$�e�<��k�	pe*^�W�k��<|�>����������v��[e��j|�lFq���dD�|�ݎ�F��J<	�h١���(U�i���\�Uk�7yH�I&�P�ɕg������"�[o�w�Xw�
�T�9��)�Q�O��������=�\�-����fu��!@��򘕞��;�c޲Ut�
R�b?8o��1�eiv��C������,���uA �0�r��GEYB}s�V��e]�B���S3�^R�~<#��Q�w��Gܶóo�Ib4��3<pՃ('�-���'����Ʌh����l,ˡ���&��/x\@'���� �l��ΗYǢ �ξ��D�+���!���gẀ���D�Ze��dEJg�u]1��������Vq�Ċ�&!��q�s�f�(��L!V��r�+m���6�� ��ي̚�̌I%Z��)îݹ^e��S�#o�^�`Зq(�Ȫ�
Ҟ�F�ш�L���ps-���յQR��J.8'(*���x&=4�s�h�SP�b
`��Rf@[Eߦ�:�p)���ew	N�B=F�p��s�	c1��߇�v����R��5�V�l�*Ţ� �Ds[�u�d�ɚ�_ge�)�u�K�)�	�=A�gA�̒�P�v���B�&�]�i�Y:)�$X~�z�<�A{� ,^x����
�d��i��������kn���B�_� `n~�� Fv\�ߔ�^#��L`�q��T���H�)��Xd/ƭ8�����s pH*Ȣ�ݙ�����*�
�� ���t���h5���ꌧY�/~����U�R�6.�XF~k(
Ē��(��V���/~z�������\�qj�s����'�����
�����4�zG^�O�;,�S�S�F��~�Ѻ�U_�4���ˋ9��(m?9�f*���`�@)V'��(أu�y�&������3�w�O[��9X8	�P�2F<@w ����΀c�_"��g��V؋��<oh [O�3���==�׭[r��
��,��^��=��C�*��6�7�2����h�g1eH��/vv~B*V������E5�#$���~<%[� �#�֡" ~f�v�'t�a,�L�b�M,��v��X(�f�xRٮ\VbA� �O�;���P�e�t�9{c� `8M����dDa��� �h����)\	�i6%�|{}�o����b�ks2^dٵn�~�}FR:)ƾ_�X*-a�3>/��-A���e�SR���M2y��H
�K�/�Zuf�{��{���ڥJ�,\H��;�s�c�J�E)#��J�lr��	$�V��=(�x��<&�4��);3�/���%p&���:tW`m\�"F��l/X5K&B��\��ު.�N��ǲ�f��s��@Yúle�
-����?�k�5	����}KC���-h��T�Uk!;�|Յ��mյ��t�O"C����1�Ў��=��CL��E���Z���������;����/Υ�q{��u"���Y$�Є��{r�J,S����������P�r��+����KQ8��Do�ǰ�(ć�#���34{�����E������MI��.����Rq�,e�z���x���7�y��=e�ꇀ�ܙ�6�ww��O��\Q�k��(?ߺV��2ݴ�|�����]��#�E1�%�6J2>u���E={Q�[���z `ѫU�?}���g@./���<
!4X�_��Ꮗ;�{*&mv�f�V-�-�{���
SF5 a�G��a�y@FN�!�:���Ot@���;������1��^e���p�b�uR-p���ʂ|[����쟉,�\Go���{x
�cH���3��)_���3��awv���e%��G�T�$f�m����]��k0#1̔�%r���*h�%* �O�y
�x3�b��y�KӘ[@��\{�,w�?��m����\a�e�m�yPT����YuJ��aN!��]��5T�����y��_�P՜�T�@�}d�>�gCl�~Q}��ļ��b�qj���]`H����W��;��YV�$��'峔nSG>k��OghO���@oLXAoZ=�TLS��9�j~�u����M�!�?����i����	X��a$y��Hyc3�s}��x'�W4���4�M�*=����Q�V�Q����L�:9"��0Ʀ�y���-��b��TS�����w��w�f����wRj�cD���Ui��x`k�wp&��
�w3ն�`G�xn/3Ii��j�����6W !�WK X|K\�vɏ�����8�g=(����3 �'Z�s�(�������ȹq(�Dx�E��jN[Y��Iq������+�ɥ v��P��Ů��"��id��;���p�\N�!}TT��8\Ñ��xӺH��a$,f�X�P�8�%a�r:sx<���I�^��
� ��i;��vQi�Pt�����ĭ���s��o��v�5��"��C�=L)�97�w��W.��	�W�B��fy ���Z!�C��ׯ�}{Z�*�����s{D��M.�j.\>�;�_��Is0+rT6ۏ�����~�b��$y7�e��g�߭���f�n�����0F<"g��k:�g ��TPn��FP�DK���g�������q�b��}�w�����o�,3���g�N�� C?��� lk�5ZH�������Y��p��2/
�
�1�U0� �+�
F��a���ܖ�˩�2�]��n�V���e���S�F����ၮ��������k��\�y���D[r�6�/	rK|b��ǗY$�����7�5 �Ls?,�FE��x}�n�p�*y�y��9%m��X���؇�nR��nK�T�m|�� 5��4�=	���!ޜ���0�l�itMn��~\��W��Ue���S�m2P1z{zƄZ}q�AI�<]ޕ
ybG�~�Dq�\�4r�FIqX�c� �h������4��%,��l+]s�1����y&�����0҅C1�?
a��׭�$���5����z�LC��d�v H�r#�+32Z��Ŝ?|yK���7Z�4fŶcHb�d`⽏ZQx:��d�)#܁�s�H��e���@��b��i��{��������pj+Px}��f8���b<%&��� {Jr�q��
�K6��*�q?c����o�ؿ��щ�j �_��a��7Z�����E\�}�}y��-%g��CY
����6����B-���AD%�����wr1���&<��E�ߙ��ku���*t@fQ`�J̃�����7��=,Wo��M�h��W'>Xb�M\z1��b���<ǅR���!zj���V]Tb��)2��������5� �G1sL׹�{��`c�um��<O�o�FOސΕe0�i�C� �,�Bt��N��� Z�O�n��A�oz�4N�~��e���Eۦ�MðuT���[���BDX�o����o���]��ڞ�S����`��������?i��n�=�����2���e�6�A���䩀:�8I�ɖz(�?�p���c�b��S�@�M^�/͍p >��r�8��`�}w���t�;l�f�X̙����]���῁�܋������J��l3�\)b����M�Ң�g��)��r��?�[��1�#���Bo�U��n��S��qv��g;ޯ��J���F��O]Yǹ�BR*�.��@�I�N����zbWa��?\TH���^%�h?Q%�Ґ߱.&���7u(jk�!{B}G��Ж���E���[�R>R�:�i�u��?G���6�\�J)��?&ͺ:� %�L.�J�u�5�	Lk�`9��PnoZ���^�nd�ʇ��%�xŲ��VD�~�f��NG<�k�߶q���<yM#":(^W�G& }����? A�o�����8���
�I/bbJ��,��N��/�)�#�Ɣ�Ҷ��آH�D�`�5�� �P9j�`J����ݙ�lW	�!�
<_�k ������@ނ���⁼J08F��]�q��̌���Ynү��!�S��?Y$��WKߤ�7�+�+��g�����#�L�¼��&/��l7W�n���Q�Ȕ���Y]���֞�{V�Q� @*4߶B}]�/�EX�,gD�g���j��l-�+؃��MB&����*���k����%9�����v/K���'�hb�	�	k����xf>��Ԗ�D����݂�[{+J75㰡8���u�⮝5���	zr��T'���l���� ���6�y�C�>wi̍ۘ$��r��1Q+�t��3��A'�(����G"��2�=?���'��,���|�ۅ 7��{�TP����1���)�/�H�K�����70����3)&FG�l�b��Nn��L0Ә��i�;Tq���Ȭ`e<PA�1Z���+�8R��5�K3���KU��=�sG���ҽ "(f
����9w�2��9F�$��a�����R�y��ٛBCo�PL0�>��s5� '�T5m��ȬG��5�/N�T��@�D�#h�������Ԋ�|�C��A�:�fΩ�?�e�����{�����N��<\�����,H��=��V��C���pNXo�E�`VI.�q5�1��L"4�����߱/���F�h����_�(�,� ��'i�S�}B��?q�?Ŋ�Y%��!�P�1g�&gfDb�\�����i�?���a�|��&[�-˓�.r�ǉ��'�	�}p�����ٝ.�e2�&��	&_Z�k�\E��bP׭�>-a{���!�j5��X.`���@ʲi�i�|��[)��t�����_�7��P�R�(x%��eӗ���}���J���}z�0{�R�+l���oWzZi�w��.�ƿ���x��w&>q��h5xiU�L{�L�)0��Wfp4o"�@��ް�g,ϔv�ļ��L�L���=+1�\c>Ĥ�s�Ɗ�%�g�JNa�*5 ?}.��!|��X^=5�ps"Yp�+~\6�/)ە9�M��O
}�ց���p$�l�^m�o����Q ��<����"K�?Όą����W���Q��
 �G]9��܂�<�s�n䣭�d")�M!r�2�_П���"c�����m"�u�K�T������H�����Sǣ��W	N9���Ȝ� 5��	�S3���:�zp�g�u�Vx6�����!��u��QN���Z?X�)�#�pmK%A�I7���3C-���P1'�v��O� E,�9[;(�.�͏��[�EDp��R��4]m!�ώ���o��#2�<S�	 RF����|����&2�¹��X�ZHg����q����J� ��"�M����n1�K�S��2�I����P��F4b��Ŧ3{�x )%F�N��\>����p��D������z�2��4Ҵ7�g��,�WnPj�٘��֤x�BkS���On�Xm!xHgHL�A��R�a�Fg�k�sY6���k�#�j���GZ���_PJ`ȫ;VZ]�"��B��v���$�S>�0.�&�A�R!j���UU���WfD�a��ER�P��
&k�(N*?��:�S56�y�+�R@��tz�f� ˢ4��S�K��]�	�(NTb��n��:���]C�O
�SJ0~l��o�m�ҳ�5�vP�,����E\���~H���|���� 4.g�G�-��)ě+���Y#2
v�c�WH�$����bN�Ӻ~����R5�M��;^"�G(~�]�
�8n�<��m3[�,���s�f�?N���^�gU��rXr=����>}������xhGM�^
��i �<Am�vXQJp���dO�ͪ�`A,!��_�$��
~ڢK��4�k����,U�+!����%�U$K��b9f��su1l�3����Z&��/�L0ݯ�'��d8����y�Y�A�$eOK�t��Mk۹��7º)7�$F�=�czN�ƽs!i���~Z���M0t�/�^�����P�z�y��P��|ufU
�����L�Q�������ɩG��9uD�QH�7�M ��CgW|O��+��K�#�Tݚ�^��mq:dl
5"���d�.��m���$|��O�����~�zX?x��V�%�>���#�� 4kݳ.�(������1�%�$[���\�
�E��m�@5�����!al��Pӎ׺�u��uG[L�a4�d�_=�����Ӕ�|A���������3=f�{��K������i3ʕ &������Q�'JH� �[�
�'�{l���@Z��P'�
@y�\'7��i}����݃��a�5Q� jw
��I7硵�n+]�ơ^�:�om��ػq����5T&�%Y ��.�KZ.t	Y�( г��M�u7f䇁լ�+s�n
=���L��x�I�p(¼x�<����(�	�������_|I�ܓW_��H�Z k�h�Y��#N���?l1�3��cW��tm�"���"E�h� V4��!@��Y
'
�Gq5�)"u�)��p|��$����̠`,̆���!��<y��|r1Q�#��`���~���T�^�o������=��|��3��ٵ͹�z6>��7Bx�F;�������u������.����A�w���$�.v��nS�̰���.��}(�x���}�v��+Zk���P��z"7���͎ �d-.�:��<��	��ʎ��'j�
|��]�����=��ыߢ�
��JU���W�L�)1m��N�`��z�@��L��D�ޯ��@��S���ػ�⬋��8�J��Ҡ��r ���MM����e3��%��J�>�&#" k�O�w��ry�dӘ�Y�ȣ�Ճ�Su�ь�g�@�cq]A�j�>�G^�$���AF�����(3!���t����G��(.u��i ��.c�~?�i9������2��d� T�3�9�o�B杼;:s+��I��7j�h�Y���� �D�:Ǹ8�%ŷ�%�s��A~l���U?�R�y��SV�z �9��%�a�2J[O�ec��+����na�?���,�/�p� ?�Y��F�&�6f�&Dp�&��/~_�eX�����^fe�t��+5�� ��x�b3�yB+1o����^���{l֑�\�~������$1�ZyùX�/��i��5%z����9����̓�+  ��U�Q�z|k+�t
�a@�Ϲrrj����x����ֻ:��se�׷*n�w��C=OT�s��%n��j��������8mAl,]a6����&�9��n��i���t	�G��o�1����]�1`���R_�_����-��O��ɏ.gpA$��d��1��9�ޏ��1��_�T��:�eq {���l��b]�	�E�S%BE&��.��x�u�'��f�f�PrU&���W�Y/��+i�ً���(Y�RЀމ�2��#��Z�}�Z�`z� B:F����C��DV�"Z�/-VA��)'��VP�	�U��-�E�~�	�i֙���+?ۋAN�D�7`~����P7�-F�8ڜ�B�}�i,ݛ7ZT�Z�=m�-�w�lE~�8�5�F��3�Y5
��yфx/�.�i2{6�v����H��u7`���k�Z�Z�#�Z\�9������nKb�PQ+߇xI�:s�S����FcQ?��	c/J Ƶ�EG*n�E�{86?���l`��p�2~��,���"lKC�U�F�K�F@J�Cm�5�s�w��(��\Jf��Vk�wNb�X)0<)�98ø� �7Df[��`�u��I��Ʉ؋d��O�&��"84�\1'5aT�Ğ��8sZ�uC��Դ���cA�����R�L���8iʱw8H�G����5�+ޏ]?���kJ��H��;���'�GN�|IK/��͚���P��`�K�Ė��Ś��&g�C,OS��劂�uZ�.�⭬'��0��P�N����Q��p��&�z�^�46���@� ,b�8j3��Ka�B5S�d����>���C봐w�˔�2�?7 �������:�_�8	��P�0�hc�9Ġw:�DWV	��	J���o�h��=6�R
�Y�4���2ccEIZM4:�i�%�V�M�n�;[å�hƳ�k�T^S��?��(�Q2&��+�kG����C˞�l�-7S~ǰ����f��ʌ깧+=Xdn�\�𭏖��!�rT�Z����M��ܺ-r
���ʛu0Kbe���gk�2���t���L1�"XZ�+e��*3bUa��L��a'�/�2Q�Bۜ4q� �ݝ�d;ʟd��H�JIX�����E-�<#~"8J�����G�d��\M�c��q��A����~B\�Q�����_b�+�b�4�܏�=�K���W�n��`���$1	��u9�m��A:��{]h�N���$ n^�
�L|��<'m,+�3%)ǧTI�[���nIz�T�ȁЬP����Z� �x`O�(��kbH�o�Y�j�A��=L�Q"�'A/O5="�>9�p>��K��E�U�9�8������l��(-�ߟ�:�0`�����V��Ő-���p	��#�j�qX^�n�]�h�H��#�Z�B	ÛV�x��A���z]��)��9@9�h�M����2Y^�W������K��or������l�Y������ v�+rOC��m	WX�X�p��G"�w/���#�z�u�A��\6,�ܔ� ��E���e��۸sI	�����	P�$�n�3�#"�,UsV��q�̞w�4�<f*�T��׻9�J�D֫8X��H�+�y�3U̡��MF��)\t}lB�y�^h�+4f��!S0y�y�i�S�I�k���~�KFwd�(�?� {ꨃ�����oeǪ��Xb(r���3`7^��t�=��w�QТ�������/,�6��ZoB��%�ī�+/��8�mp���!�9.�d�#��g��*WP=a�-��>���i�����F�b+:�������1���ɐ����b��#��-���X�Z�S���D�l���$�9���Aaa���1�B��$���pG����#5�� *rSO+6��դ���
t��R9�w}*đ�ч��c����yFfѥ$ƚ�Dʙ��a�Tz�����#��\�
���E�)�<M��l�M���U�5~+��wu;�bҌd�����7?�p�����UF�9F2�)>$ �
i�,�c92_�B�p�~�d�9H������Ltm�Xd=W�j��dQhu�k~��֓/jD�@Iޢt�Z1�W�;��.N�A�՟$'e���#��.�2�[���v����:��z>���z�$\_����ɩ�G��*�ME��u���Gv��s��o�?R�[�<M��J���H�s�\[<��w���=ڽB��9����U����)V�0 ��/��HW�4��e_(?��i����RoC	0�:v���G�]����1���)��g�ύbI
�+^kH��qk�Q����4�?9u�-�ڰ{\����59f����5�S�EX�јl!��ڝ,-�� BUa��|4�$f��N��Y#������8�ܫ��©�9γ�Ǩ��G@t4	J0�6d!5�$l�_�X6� ]ֳʕu����\:�Η=Vz���c����O���Xdư�<B�SjR�kɌ��]�ͨ̃�$��4.���O�p�s�[�����UmJ`��f�[ʽ�p��m�Wo�����W �������Nzf�a?Er>�}ϒ��=q�ߡE�Z�,=f6
����DC�ߗ��Z����|�E�P	6�u��c�u qvHh,�s�ȩ2q�ԽlUi+6?�l��H����^��Y���-AO�=�O�/W�A�*2|�e�Ɠh+��
ԱRV\����j����*��Sm��o�.�`�6v��U�����_�����YW�a+��s�Q#���!E��c��;X���O}��!��_��z�L^��-q�$+�!�*~GiټɄ�;gdt�����ѪW��zʑ1��q&������G?�
��[�ٳNvc��X�+�w�&��qaą�4O)�ڔ�-�4�_�ٝ_�l�%h�sI���c���7g���ۘ^+�mGNr�ܮ*�݃��k��������n�?���E�2O��:�'嶅d^ȍIO�fQ5v���J�A6n0�X��?�et^V��.W.:�-�εF��}K ���T.%�߼~؟	k�|�o�b8��ip�U��nk+�-��&�/�`
�vS3������a��}�k���l�Fw�[x}|ߘ��|����w���EV�`�A5�΄��'=��[+��4ٜ���cwa�9t�
#պJI�Rh�n7?/+q�
ol�w��ɑ������iH�X����O�+n�Q��3����j���������bA �\�b�8�.=&�����ފ̙U���� �U��6���4f�`��.R-fIR�`��R[�"�+Y1�HN�u�tc;UL�_(���O�Ft�z�s9]�
��Y>/����J۳�}hиhR���Jq+SQ�+��0�~0aT�C
�dξ0/��}��.5h�YQ��ii�-��y5�!�t�V�9dp������<bp�FfX9�'u�
�ݶ�hȐ�8gC�f,}`/�%#���P���ݔ�9�z~�� _G��ʁ^�˫x�psY%�}{��R���J�ō>�����r�߻�Ze-ī��$U������$|*{�D9��g�|�^D�����S��e�¼�|�y{'����>
מ�z�w$�d]SF�k �1vwKnTOuÈF#���;A����0�j}�O)�:�7�{� lk|{����=Jô#j��#���<�Tֺ͐�����G��:
�4~��Z	���J,9}~��7�����ך�,�-rW���%+���*�r���
^W*X�#	ϕ�V�#����ߩ��Z�U��_��	=���3)��2����GT��H�uy����Z�L���4��)G�OO�N胂gJ~���1`�i6[��a5~��h�qr�3��4ZS�'}����5up%"��Ǧ��#k3晝U]&��z�����45u�~��z��X�tc}Q���,�Ѳ��WhCUG\_�y�oc�IP�9)X*u�9�$� �է�k�3G���O�B���K��2SS,�d���Y�(�P0R��e"4[�݇��5�ֻ"&O�EpE'��R�`��
�I��&N�3V�D��`:�s�l���X5P$,��\����>��s�9u��>#M�Ά�9�}���Z�$���9��l�`����I�	�o�˷�?�'Q_��9c�zO�J����p"�y�������ܢ��$c�~�#��@�Qd&o����h���+�c1�5>��H�1T�Q�څ�Y�ӂ�N���{���N�v���^$�2f�T��Ȅ�%Sq<��O�EBF��o㫢f#�@�s�z��:���|��,���q����RP�25�!�=��R촬5R���N����g��L�:kB��[���r�����v��|%k��`2C�έI�?u��h>�<�.�$�͵����qʌd��g\�+��|6��m�R��Ui0��")#���a�ejC�&��WAe�����L�p�L=�OZ_u����⹽��#�3J�%��TU�Q�~T����R���=�-d)��JuLӄ!Z��f��Њ��%�����PEU?�[�Y������=zr�n۴��n���;�{~�8�LV�7��-7
~��0G�EΤ�Um�.C���h�����<�.Gnhh�I_YF��!�뻊|PTq_���6�����7<n�ыT#؈�=��%�9ܒ�#�t�A�Y¡�??+�&��l}��}vB�p���Ն~���V������j�`������3sh�㛎dw��W��^��s��5���c��~��%�6K�-I:�[ �U�����4]��W���Al�R$҃8}Kl����QTWV�d����ZZ���\�2�F��9q#�Z�U�G<C���<y���ŹT��ө������jܸi/d�5X�Ӽf���+N#�d���`�ʹ��£]� ޝ��r���p3]eg5$h����+;��7�/�,%H�'6�K&�C����܃ߓld��x����w�u�Gc�UM!��u�A�(9�&U���"O����6B��J:�i�J��
q�_�2���M�0���{Ӈbz�+j�����
��L=��3+
W���$��1�2c̟N�X���4*1$,%�ɉ�"�􎊍C���i�ʪ:qI��eN	�)/u�����kHu���x��Nڧ�#�d�"�C�+��bGB�N}��
���Dt6G�)Q�e���YDw�9�]��ЗH��c�=��Z#�%P�㽾��y�W�������X���e6�@���$��(�IH��{��KK��st@���߷�O���<�<dυD�w�2�l��ݺ(=L�Xg�5�5}b�#Ϲ������_ĕ�y��a��J ;������U!�!�����$���,F�E��4���/K�WLL�	��'�g�q���h�O�z��1!��y��6&����1[YO�.�{��e{\K�%���B�ϭO�xN��}$�p�To��+�`�O����=Z�z�G�R��zԳn�Z���tY�-�q���ާ��+]H-����ݾIu-Z�U���B,!}*�[�,�}?�i��5�ȸ�٭+s ����Rpﱱ�]ܲX��b����]q�r����Q�%}��^�V��<4��M[ ����|or�Q�+g>O_>�Q��̾/���p�����8�M�k�98PP�8ڃ� �$mC���趥�Vc"v�䚏.�w`BM�-CP�:X�'�g`��<U�)���j����d��d�yr *Fa�����D6)�|ϵ6���k8Z��fL2z�=/�r������O��̖L>�q�Ѷɿ��U cZ��{�쪟��T
���i�׾��}��Iv�EI�����0,�E$�;k!�a�V-9���j�1!�p��p��ķ<ι��,X��}��;OYH�p�~{LG�?S�=�d��&���LP �x�K�%���jo���� �d�鶕�0;��}�%���#��L��/�ew�������ܬϋ������x�r߼W|�h #N塞6-�A �]�}/��[�����8L�����%���&��Q[]�8)�o����]SE��
A���Q�&�^R���G�S!���6�8�;�R�(��M�RdN�HGزx:_�n���;{�p��-T`Ʌ.��`{�T�3�`i��iG��L5�Q�O���\X��� �ge��g�D���н�rM։.��C0]��k�e�,	B��6'��ky��vZǑfI���j�ôb��5��h�6��͊g����?���n�đ��o����.%UǤ�����΅���rE�	�~Vߧp9b�ݲ�N2�2\�y<�|]l_�"l1�/aHO.��m��gn�#XFT,fRK,T��=cx��UW�R�:i�"C^��~"|3�^��ᑇE�E5�ti9rA���f7e�u�v�������z�*��N�i�&��4
#I�������9�f|2WD�>ޫ�	;>DQ�2P Ө�T�:�i�=����W(����b���8d%�xt-=K�ʎ �\\Z����y�6�y��`���2�i�x�z8�bН����D����3�m�[+wpK�8�� {�E�Y���#��
�2`2+���Zj�۵�{�S[� ��������_w�j*r��.�y~k{�v7W��1�<��Ew�@�k_���7]��p��V������n�=p���숒R�֤�hv�!��E;�"�zb�!��&3;�J����nh��Sf���;S>�
���Y�v��/-����y��h|d�����τ��h����������D�e3�P���^+�4I�i6_�����,Q�&u[XPl�$��0�� ���l���q��}m!2JH��U<��&F�I��AG�eT��p56�?h8%���q�;���@�����$���"&��~*�����&�`�2�|)V^�{�A�?�;�$�ߝ�u���ĕ�h3��s|#;�����0�	D`*95�s;���Ȋ�^���'!CoF��[Ȇ�p��*ұ�+@����u_f��1W�(;I���1�R�2=s��,Ĕ��od ��m�VdJV����$	�Gr%����z�@1��x{A����Nj�Ï���l��n�1hy�D��a�"�����2���g����kF������^խ�n%���ر��"U,���t�T4���iҡ�y �׽��Bm5�)cj��Od�:�QO�@@���+פ�F��{��{����
���qB���)'�##�80������Duп�Q��y�5P4va��n���fV�Y��E�"�э��DP� y�h=<��+r)�Aj���/R�VX;o��X�]�s��;���l�4d!�k.-��񥸞�@$S�+�X����A��-B�[�ci�\#�X[ꉗu>j�V����	�K/���U�b� }���A`�d� ����a�����h�)	;��X�B ���#��T�X�J��!�ϐ]��܌���]�cD��}a�$�'���v\zJ�W�>��j�E"��-�������0|�F��"�A�B�^�K[��Rv>o9��E���Mu]������*��q����xI����\�-�����
�Ah�k��̟vFI��Ou��F7���ֳ���w(.@uh2�ʑ��)�)��!y���x����eL0�M�+�pOWP7#ʙN����˫�@B���MkO��wZP�+\��}��V�@F��yCZn����jb.f�x��gD���ryc:߷����󜀡�^m����� ��Ī�e�j5$b¦sz�;��9/��ʔw���� �ߊ��)t����:kB(�\��?�����=�lc%l�?yE��Y�r�uL<��9*V2���nC�5	GI	�{��ɡ�f#�x�\zb�+�5�9��V^���׉}�2�������>�y3��.8�ʩ�k����Zmw���(hd���*Ҧ	W��PE�r`�C��L>���:v6�y3mh�Q�8����i`XG�:�%,��%6W��qe���f~[�������1�j�����u��6?�(�b3�`�J�U�r��'��%�|��h�&}z=���pM7H��y�[�U��� �e���+��̰���jXl�l�f��n9$P��X����m�^���L��zP~>��+����Q��s�wu�&��my>�(�\@�ûq�~��D�3���1z�j c��;t�9;�g����������)\�n���I+�h==s���7�雇�ĝ@a�p������\i7���F�%���<�X$?w[��q��ŃN#+8S��4Q��/��Ҏ�S�r{��@�-�i�\��pP�$�������!����|����b�Ц��2/���/V{������Me��Ƙ/8�����3��� �>\���m�����;=#}���H:CF���r���{��ҿ����*u�U�'!�"�� ˧���G�Y�G����w^˘��1^"�G����,j�h��LT����r�0&��n 	U�PY�6�!���IM��)�}��,���Wвݭ3Y}>�'��]J���`{fn7��@�A�*�[����CgtWr ���%C��=9Fhqlb��4�K�^����nu3ઔ9'�Z;6�)�6<D������I��˅FQ�X���(O��e;��K pH�A-�����=h �^�iTXeR��q�������.�L��n�k�d򷐁&���ў�%�/��_����G=�~���ŕi~�^�^�*ґ�ٞR�?��`hn�����̬�\��#� j��f�`�4K>i���ܛ�nxU��RK�%��[/I㾨��m�h���
�U����@��P�z{&Pԯ�bN��H�ȣ~O][;-n�
�Š?)��M,���M�)�y}�q��Y���o�.5%�z�@G���ѫx���)F.N�l��F����%��g��%�6n�I+��K�%��58��Da��f�)n�wCW��p�)���8�):�:�j���GœSI,�_��t�ý���	W���N����U�����f�Ln��?��}=X������կ���@�(�_eE��壯@�d�ˤC��ȣ
��F�:k嚍(������{4�YG���'	��z��ٗ�D$��\�{������;�h�$*���6Z�?eY�W^���5XX�^�m�}�B��Jw�_�JIc�_>-F\*�6�v�p�:��s��B��@��e�t�Mm���qb��E<La�����]!�i�U���]p��S�S�:��f��$�`uLU 8՜}c�d�䚕�,�ֶ��:BC%bc�<)1���|�s��v�M]bΫu����ج��A�������]e��%�T�<�O�E7LhD������i�/{�-�2�ʪW��q�^Y>];G|�;�{1=����3�c�W�F�?ɶ\Gu��ί������	�e\�b�y�dq�Fn��"��1Y���� ݛ�e>���-S@}��[3*S�����I�Zۄ��=��iCہ���v�g�:���g#]}���*:�]�g���m��x���vt��]-%>���7?�ա�=�E��7c���b@P�SE�g�/v�.1WݟL`�h~�S�H��@MHժ�F�L�HU?���Y���1�����h���#~@X���������9�B?H/{CH �7�Z�yO����i���o�Z=c����P�C�Q*7�9b��u='%�2O��n=�C��4�uJ6�g��q� ؗ_Ĩ�[M ���ư���<h��1����3Ͻ�84G� pΥ�h�Es��*���<m����N獰O��#�H1�B�i���'p߻5d��װGkd+��A��2Y�9��w�*���F�=�� 7Ə�ĥ��	>'�T81�I�m���ߜ=_1c�k��|ט�9zoy�A��iF9��x؁�T�Xu���T%���+;'��qK(W����R�N���TʆEU��B�
�vD��
��EW�U�>_֌(���L�h�
��z;*�f�6x�t�sL��VQ{�Q���/b��_�-:@Za%�Ǉ�y��z�/��)8�d@���|�4XGK�mU���s�'����y<�D�r-���������="B�!�|r����(8�+�\�E�gW��N}�ZCP['_N��?]cM�m߱|���H �qH�dw�F����3	i����a������t�{10�j�^<��z�)hq���KJ��@��.������o7�_)���|B����s��BwX+u>���||$���1>�>�&��p6��E*��ȇ{5.� [�s���_���z�Zvՙ��I�n���3�.������B�]��;����	1�
g� ��ް�@P�s��܄,tg��%yd�=�R�<�jn���U$�N�,�K*�*u���P�ݮ^��'^��HL�)��U����1����;%1�]��� ���sT�r�J
��9�ORu����Ŀ��4uEKc �2�o�.���)�ެ�'i^�j�-D3c��G��K��OeG�g~�ش���\��S���k��f�����-�6��:e��XO?[��X��9�xB�@*��u.�%��K\�N����k ��H�B}��m9�*��Հ����5
��ʘߏ�&I�#ak	��"Ώ�;.����N�j����厷}�w����_����@�⪰�-���J��m^)��)K��
J�)Q����y����X�6��8]�V1���<eZ���겔irK,��a�/�#r.�t�Y9�aOq�UA�,G�9F���\|6/ܼE���+�-�٬/^N��S&B@��7���5�>�9�P��[B���F��z�KB���&#5�ny鲪��>P:ɧQ��K��N,re�඿+A^��|n,P��)/`�� �5XL(}h�Z��t}	t#Y�������Aʴ�����k	GÎd ��$���q�$1v�Ox�WZ��D���!@��U�t�N��uI��:��x��L��L_'�(?�-D���lt��aD�&�r�ꙮH��M����hW�\	�;4�e����\ Blޫ��=��]�-�������Sɥ��l�<ڐ)�Q
��%����r�U�|7<�v�04��L�Y[	�΋b���ħ^l�V�OQ`��^�kV�1�_�����"�F�p��JQ*��T�h�o�B\r�(Z��z�u���)Yh��>f-(a+Wo���1�v���T��m���atf��;���6^-D[dA`��wŪ:҇��b��|膺���9z��� C�I��(���A�sgޮ����n�*�d��.3�<�<��^��N��p����t�pV�!�J�!۸엀Y#OcN�0>��M��F��))b���LI&L;���&�y����K�[ n����"��t^$Мr�ɉ�!��#$��ޢ��� }�1�����"���2�;�,d<
ݣ��;�Hϑ�w�񪎒~��{}M��N d��ë~��H�/A�w��t�4t?H��-2�5���A\GUZ��2�,�>��$�x���^���B#9�r��١Q۫�����T&�J<��㞭Q��^���a�s䁌,���"yB5I�X�z�D��ד�y����e�&
���v!6z�N�p��%��lb<t��P	mx���wJ�]��_�Ĩ���p��
��$��u;��i�qG�
3�.�vr��l�?d�R%`n�g�=�\�t�߇W��p�u�I���G�a�ќW��X��ʼs}|�/���5j�8��c�=c�/�pQ�Q�D_j~����[(�*"=���L �Ye0">���z���زK��:�8�D���.{�8�9�bИJ�j� ���I���P^o�D���>�-3���%[-Z;�z;�g�h	i�W7<#b����]����e�5��mؤ�>�y�f4�F��wA�1;�S[�o��e����2�eS�HXX3i�G�AJ��+�=�(��-c4�Aŕٴ�ymP�\r^�X�&�-�h��Z�T�^�&�yV�9�4:��+G�sw�P��\`�:l��Okv���*Ac�tpniб�d���������wٳ	@ʟ��P��Ȩ�l�R]�߈m:ԔMד�?Y| �@�#���t����QＢDψ���u�I�XO{F��M�4�'@cp�?B�л��M�
��D,�$�J8��W�t���V��?W�r{�IƆ� ~���Ʃ�c��U�m��F,��V��;4^��R �-�8&�  �[ ۗ�ߋ&�L�U��Ѡ]��ռ²A����5Y43@5�:�%ntm.r��<����u7�X��8��]sb���r�3wM��}`:0�1^P��OJ�Q��M��'���?Ͷ^΋�,i�L�j,y����q�>���;X������h��%�L^�L�^Y*j�������!�ޮ��׽RJ���^��{��x�~	�X�m߉�����#�]�A���^�-Ô�R�B���HS8��{��K��;�/ ��n�ޛ�pc_6��$=�[y����g
M)��iQ-ٓ���0�K�ᨺ���"�*�V���3m�(B`͉R6���_��i(����[��X7�d�)��E8AT�~f�2�ٶs����C���|���`����b����
�{� ��C��O��z]r�r�ʚu^�3�¾��������D���	���q�����i����>��>���~�E:i"S7b���Z����3}ӡyxu��Ki�Ӿ�./b�i�"��Y�nv'���a����Ux/+[�?C��Z瘨�2��"5	7ӦX(CD���e�i�/,�Q�t���Wᾥf �,�<9�eF0�@fof"�4��D`�Է��/SBƔ�Z�"�}l�[�4���4��6�,3�����Ao4���嶥U�#��~�h��BV����Z�$����	fq�o�S�g�C[Ay;�A�مTЦ�$
_2��#.��ț۟��^�S.�	��|�]��"O-�_����uO`)6p���U�r{-K�Ū����a���h���ޓ�X	�j��3�R	�Lqa�U�_��8���W�/�ӗʟـ*^�Q�x��Y���B��Q�0������	�~�;1׻��=��{c�:p�[�H|�k�;r)��]��$��8@#����U9��d����6w��Nă�+���J,q�@�o;0��!T3�ƽS9k���&2�j>j�1Y=�~�\Gp��s;�>f�[5MUOxkN�T��A&'��
�6���=���F�D�j�������*iҎ��dX�����n!/]-�ɦ	f����S?[w�=\x��F2�zsC�����ސ�h�'����6k�׮<�̾tW2��M��Bi��寞D2@b��+ih��+�6>�H��<��p9��2Ҏ�p8�@�pz�/*4��;� ��쬐�����I�gA�´�=��0zڮ4��T�C�<0B�D1��"ek3�_��Y-P*O�M�]8��hT����E�lA��݈��ee̮DtC����B<�	�3ߕS�k�[���Z� ���F0�5����Z~3����ل(c��=)\/�l"�舤��_'���&��FX�M.�N�!:GUM��3�|C��,�����&sԚ�Tn}��d:읲%D,�g�=��i�λYc[I������>-��';�?�:���K�C����=QRH��7����u��r�p��@�.jcľ��\خ�f�Pv)>���E��p����>�^�ش6���"��8rTú��:�߭ X~��pƭ�!-؀�1��N��pF��<��Q 4 �fM�lb��v�X��	�o�ݠ�,(91Ѧ�&��4������&��ƓP��Uĺ�|sq(�RG��Z��ܞ��/���m��S�i+�'�[b�o��Ba(�s�`A4�4;[�b�fJ>U�/�������� �7|�d�8`�e�cŤ>���e5m��<�=�r,�Є�h�j��&� ���O�O�K���wV�����rt!C�˰r����B~�j���7�;e�,�C��쐕�y�3�c��i����҇��q=����̯�6}C���Mf�(��I�.Xrz�sA��v��g�����u��P6i�̍��ͱ�F���EyS��G�;�!�ir�����L�	T8m�C3�QEj��]ă���
^g��*��p1I�Z�na1���H��`Ģ�ᐒ�a"q��L�-G/���!�D�G����9��'��O�����kul�=#%���f��H�������4k����x�֤��j���Qd覮�0 � ��؋/�I�]�S��ǝ\��$�����,�w͌)܎�`��V����	X������UE#����n��O��	���Ύ���̶�D�:��wز�z���q�Bl�g��/��.����g��P��TT����3!hxh	�Q$������(kư�ќ���wy	B_�ڴ\M]��ݱ���=��G�;𝹠��v��/m�w�?�.�:PPĸpY.:�Qv��ZbS�W�l���NĖ�{�/�bg(���r�z�!��2�Xٽ��Z+��`�r؟3۝���6z��<<����P �ip�i&|��x��qv�@!	�b�;,r%�S!�]�`�ɏ>V][ʻс����^A�5�)�ah5(�p��y�򆓲�����C���@`�Z1kr�"폩U���~�����S%X�܉|�<KލJ��q󃑵S�B���G1P?F�M4��_9�h��4�,�F�NQ�:>�w��D�-��wRB�ǂPU���`Q���P� �b1"�}�P��e���m	 �9;n{�-`�6h|�OA���]���Q�F�N��m�C�<!l2dU3?��tGb���1r��DF�IX�6���c�Ao��S�!]+6<��6��reB~{Ϣ��X)�5t�b������̳��[�7�a�ׁ��\�a��m�`�VH�듓n|��>o*�E,a�a�t��4tO�7�zJջ��S�M�A� ��z���ΰ��5{g��ϴ��^&Dݴ��ҿ�����1.��w2����IM�����M��:T |u�Vn�)Q�m�0�Y�"R/��IsQ��Ďe�-���.otZb�A�ǘ}��W���؟�i
�:�����@�_��B L��M%<XJ<�di5�V��S�'�)���P�9�?��Է�-�V�*�~�g���v��=�J�����y����2�vL*�u��#(J�Mpх���W�V�i���2��)d%&cC��q�9X.��vhf{�ܣ<�H��WM|2~��ם=h��wD�����Н2J�h�ּv��`�!����� ���m�B���d!�49]q�'7d]�W��;��s^O7�<#��sQL�ս_\����u��L��b�Cy�P�
K1]ms�lK�o'��z- `I�6�{j�-���]�7��ܢ嶫yb�o�J\z:��6��ߜ�(�mڟ����-|l}�q�M���N�# �{���!������}c]Ҧj����0�'��{v�E=�-Dtr��`�r����Y@���4�vJ�M D��ɹ��$ � Vu��`����nUH����2C���$�'�$��Jp�'#��EF��I����lܺ�ޖ��}a�\���3f珲����ʷr��a�g��+w���c�7�\���1G�η_
:��
翸�>+j_׵�qP]��B�s����t��L;�;�A�� �T�'Ew�k:b1�^�IP��]���{�"W����1.��z���\q�jၺ~��Vo�,�����|_�P������[�`>����邕MT0�̏w'��0 �v�o���
����P�dā0&���L�"��g����Bbc@�\]i�(����z}õ���Pwhvh)ߥu=��翷T�3P۔d��!����s�0T!��}��݁�Z�nbPB�G�֨��P#Ȳ�ӗ.���M ̅&�~`�`�R�H�4��x���m8���7ErD:/T�+��>��Gn�T2_��i�!ݟll��B|ژ��D� C��o5 �V��8�N�+���<�N'X���(���ޥ�E�y��&>��Ǥp鏔��$�O�,}C ��wJ���W����X{R���B��ُ?v�s�>������=P��8�P�I�ز��6z	�e�����=��\U�:���!p���������,yl6쳠3it'�@fx��8t�ʢD��4h6=���b�ߕ��Ag0��9��j^�vT;��5qu�Yelm�6A��-�x�d�`ʺQ/��%������?�w�^��˯L��zI�����\�c`+|���ъ��c�T�����=�f�5��6aK�N�G}f�g��Mp4w*
�;1��O�CZ?�-ҟ�Nb�%�f��u^Ť̎�3؇"�������ʴ��EV/!⋏?��4�h4(��9��������;bTN�]8�鯪�S�?�.a�x��5Ha85��ve1�팦��z7uQ�>��ލ��%RI�uד�� ��rAl*�p|���S[�C' x�ˊ��{���R��';:P�mK��F��{JТ_��XL��q<i7M���5���9�X��� TCZ��~lԧ�*e�}������6��C����JW� �D���a��f��6����oS!��hhI(�=R1\�j�1�ܛ��?�U�UƆ���=�G_�n����β�b������n����@�����l{�pWvr�����G��v�!���$O���\\�i�7��YČ�����`'�;ֈ=E���u��6x��Jqth�~k2]�b�dvGVm;W/�%S�x�o�)�b'�ݖ��=o��c0xDq0�"��,�z�9�?<�|\�V�ǉ�&	�)�Iy�H �@��T��e�s"�i�_�x�F	��i�W�=�ɑɊd��b��n'�j��b�'�W !�7�4�؉���Sʷ��ό� @,��yVYQ ��l�� �����Oܫ8�&��a��ܥ��_��W�����* �ktY �Ą{4c:�_�&M���O��L����=3�O�'��"C�p����s)�ȸ�]ƳhD��{�Z�>��FY�H��t�x�7������Xw\
�� :�B�I��y�p��.�`�7Α
��|�4FF��Wߝ<��n M$����C��p�đ���D!����=�m�T�����&�{;���A�VL�C9 앛MA�����I��MJ�O�`��Y8vMJ�i��ʿ1�<L��V����,F֬6�V̺�P~���f�V��y�!6C���џ�7w盅$~XW(>��z��g��<[)ӄ*H�Ө�	�MgJ�8'0���F9f�+wQ���NW�Ⱥm��C_+l&�D�/q%w	hl�,�0���6xMSx\�
��1�G2��K�����<���5����pg09��sLhL �qŶ�(�m"H�����;��Q9��w0ľ'�x	&�nW$r6�5��|_��l�A�	��95�L%�K�/ʀ�f*���r�=��$�h�9_6dC�)������E�%=8|��dg�r�xWa��s�D���y�$��YG����rZ~��b�QoF��኱�����؝�v���0�}?G`$�~DF����v1�, \���]Q��g��1�P��>НˁZ\��-'��C=��@�GD��l�hQn�)�����5�2�۷�c��op{��!�I�+��l�L�)/���|S7�uP(�d#�~����� 	P�,�F�E���҂�+	B�Y�����uD.����:.�L�Io�c�3���Ҍ�q�,̩��\u1t��5!��|�o�da��m�ᑎw6=�G�<��8���nT��Nx�&I��1��0CD<M�\U>��)��E�|R�%L�x�j�r�3x�[�6Fz��������"�w)_� ��RK�P��O�����D�H'��)��G Ҋ�ًZE�ޓ����I�8-�m۵D5¹��Q��C+{]k�&��ޠ��eЭ�Y'�=!�'�A�b��O�G���=q��}m3�m�=r�#�,{kh����8�7.�V�L��I[��T�&T}
(�Z<�n�S}��[��Om�E��n�W�10
r���:R���m
2L�؃�<��g��v�w�9�Ɇ���O�n�e��T�>����CR�������;�h���*s��v�����Q���?`��?�Y].G������H��!���$<���֋I��A����0��]{��e��Qy�t9�؜��TSaa�&�q	
g����ב��G�h�Ƽ���,�M�8�ȵ�B�B����D�!I�~�Q#�)��l̕٢0�	�^�|�x+�+�o��ɍ��p����B��i'7D
�O	s�J[��[�Z.�]<��6����A�-�(�*e��r"�֧P%y�RH�ښ!RCY�8j�ݸS+4h�fj���.Gؠ^��F����ʱh���/�a��ro���s'D�j��8��Yz��%�_O��q�0 |�rCN`�iӸ:f�!�t��:�����< ���Mk�|3�~Gb��K�ѓ�d�����;�le�M=�
9C���4M���n��;� ל{����/"=����c>0� �wWyM��MP�	~+w��h�%U�N���g¬�a��N����1��!6إ�,|�,��l52~wW�P�==tz���h~@��u�������x'V���"�-��|��v@N�a��"z��k��F��" @��O�:�JLUq3RN#J���w�5��L��^ ��s$��v�Y�D$��B;�p�J 9�Tz��KU�<�{-1I���Nx�rZ&���Q.��� ����k�%����g���.)����f����W	��H��\.a���7y}o�E䕧0�նFs�Z�OH�F7�$<ޝ�zz�g��S�UQ�F{��!���%���`L�2ɥ�����g�J{3���$���\]�0~5W��)�Jq�:������@�
�U�c�]�	t;�n������Ő�q�Ŷ��8h��]����<�u��N��*�z�!!�����ݛ�'b?h���j�ê�>�5�=�ϒ�@�׃^��T���V�@KM�t�s%�����a겐JRi���n6��l)�1��UG�VFw#�B- ����E3�U��D�aksU�ś���������c����yR#;��;�m��	����k�	Ӿ��;!2��z��֠�F[�$�U8��E��:d0����,ڒ%�M��Lr���"+��[� �:�!h�I��Ѭ\�} �Ɍ�¼[+x�wI�%gTٲ��Y|p>r����J
�@�n&u�#үC �{�R��j'�6��W��N�]/�w+�W��H5�'4g��t(�5A;˱�^�l�hcg������r*efx������öݴ�?�B/�k.��O��P�/����Wu8y����%+�;3�(�]Ij��if�F��W���jb]V��Lݔ*��IP��� C��AS�>�+���#���eӜا>2�~��Wme�h�T�f�M^�X�����f��Y�L�җ�x?��GҨ�����w�~n�8��sY�4���ևn���|�,��\�}�� �&�@�R.���nF!�\E�</�J�բ[���L|J������PY�B�Iڊ6P����}D�z�՘�ӂ-�n8��%� Wᠭ[��H!y�&<z�j�<�<*�j�%��B��O<�$�pJ����#�
��
�u8��l�����B�G��i�r[%.u�f?�1�w;��c��U*cʺ�O1��p	>��H�2�}�#c�D_>��N)������E`W��!i���ǜ�V����fnz�z�5^Y�m�t��g�u���}�y�Y�j!�k�M��X1�y�S�2������ꂺ��&�8�MpD�G.[(7@��I�)|ҴPd)?����A[
{��k�� cef�j�C�j1�j3���t�/�[��L��q�x��8�Uo޿�=p��4�6>�q_�~א��SV��1ck V:�((+o\N�D\�\.�zS�4eCafR�2y������[k��Bn'̼/���)��Ʉ�h����W�^�:_��`�p�ny�+�&��-���̸�ҩ�S��T���
"6T��Pd��� pvB����Z��+�� IM�R��?�`�6K#�"�������yBF���AM�2X/o9 Y)@�G�Ӷ�/yw��{���2����05�b>n=�@�蝝Ϡ�~|87$W�:�I���aVv(�̌3\�����>})]m�3���	zi��S��m��!aXBp����@T��2�/4����|��v�`绹z2̸A����|���s�j�˻��C����r/i��i��GL�����������N�Gl�'���h�b�*�qj4�'��,�[�~oK�k5=�̼��S�Ř^mv�l�2�����V���ګ�����PKz�4����诼xYGW����UJ�ܣ#�¥���b���@V���"*�8j/F�v�u-'��y�Ջ]E�,���d�U�:�N���Uǈ�ftJ/��/.��h�S�[�N��1x��0�H�����AS�~7S�=�?g�n;��tؒ8uy��S��c�K��
�.�(��dB/���?�I�W��ޫFk�`�!��u�ϫzJu��J�ڝ:���d������x]=��GGM��A)��%�L��N�VŜ~���f�j��r)բ�@2�%\��R)ZY��D՞�gm�Cs緄i2�Oڮ�3�\?\[�&b&�rK�f�:�2�%�MӀ�\M�&Z٪6�_���`~Yi �٦��������rC����B�~E���̞w	gd6�0T]�,��QM>#R�&����ZP�9iHr����E�}������ n:�\?/"��L�+M�[�F�e#R]�(P2���돣үj�`bl�50�
�*��|E�Yp��P����'/�)�z�ܼ����2I��n��ay@G(@/�Z��%n���J��H�R=��ى�5�WA� �e�����O ��۱� �0*����,�sR�;UI?*��<�mK�T{�.y[n���32΍�Iy�����5����W���6�n�xXo���s�!���dN�����tP����믣m'��馧`�K��2�VFk���;gQS�EG�UZ��#���ą9r^E�	C�-n���v��|�O�B:4�K�h�y �}�Jez�����YI�*<e��:�V�}J���[Pg��2����&(�0 ���6E�ܟ���?�j�@&k.�]�`�#t`�I��R�Lt�Z��/E,���q��{���0�D�8s��:�ڹo��G ���mQ��`���C>-w��Q�<Vlo~���]�ڂ[�Tɩb 	s៽�X��9M��*r�WB��Y���"qJ�������c��8�=�k��"ѭ��3�����{�x/k��,	��'T�&��Ibu��y�h_��R��O�&�w��vg������1[gq"Z5#NP��o��dХ���g� O����M.�"��ؗD�妠a�#acp�M���Oٻb��JF�R]�tH�,�R��}��F�P�ׅ��x>��C���T� ��p��� m6�꧶E�lG
2z 5�e�b����nY@������G�}���ٶJJӺ_ϤX�3�ɂvo9���a衏�BX����c�@�����m���l�_E�O��_v�5_@\8�ޟ�j�'�8��EHl�,�"�	�.ʱ��p���e���^0��)'q�V?��%��ͽP e��A�;lլ���4/��T�)�ek�*�L�&�D�~瀤vv��1�g�x�Yq,����:my
hGЪB&A�5r�ucl}�JЧ���ޯ`�>6�����*�
k���}�SpA�Ь&vqB�x^�/�`�����LR���iLc}�ը��k�yM+��M��v��υ�/C���U��*I������������/f��#&*�������񝻔3K=l)�7u}`��3+��w���uo[Z�����
����gL9;���E�Gh�\͉q)�3��8�S�8����p|�F� X�tA��k����q��<����H]��Y���Q7�IX�	��0�i��z�p��2�a��i]����r�?9���|ћ��BS���$�_W����R�tΙ6��L����B-��a�itr'�_��������x��	z��Ԗ�z`i
�}���*�_<�R�f�J��Y������B��,]u�m�xή᠞k����2�w `Ny��Wu�E��F���-���_�[��;�9�Ur=u��z-��Z�Q�p����(%�����2��$`�	C�Ua]��b�N%��:�c��5�9�]=9��-���:�(��z�� R�v5���Һ����B(eXb�VL�	i/#�5�[8��4Ez�*������C���w�}.��_��-�������E�v��;�`Nzi�M¯��ݧ�UX0�O�B=�oc\�y3�A�{@~�.���/^#1�����h�w���诏=QL;� ���;�'Dբ/����a�l:$f��*��x��2Z����4%�2��#l�����;딩�s���c.��'�*pr�|�����Pn�is eֈ�� �K|�ۊ�Y��⁵�hܥ��-���3ԋ������ŧ$9�H�!�&@�
�P��W�e/�0l.�&:q�ދ����������oy�(�I��s�$LD+1N���������2���=a�.3��#�\�����q�W;F�eɃ�U�;��6����Y�[A�����i%�#�У�-9����L��	�� �,���F�����}g�R�7�$�P���!ϙ!��hVE@O<��zC���ak&�BO�޻1�"{��B4��LW��Jn(�)�tGBς�	dT�nqͻ'��-�mx��Wz2���ziK��D&G�b�J9F�:��t�C�h�!�]m���m_k�uc2��6�����y���)6[���L;�ݾ��rbauW��]���+P+��T���X��Xlz8[9�G��e�!�!�	��[�&��<x+9tJ��|�����'�Z��߆�^���%�����.Op��v��l�����tC��N���#�a{�Gmõ�4�V~��A�����f��y���c�����=��+`8�>�����/pfªn2��cӿhq�%P���n����t�1y �+�Ɓ��j���H��k�P��y��>��� ЗQ+m�I�P��c�0�홹�����Vx�Ϥ���t�{�l����7���AA~�uj�#˕oM.����9�t���E���<�lět�3�1��k�=�[�Ƿ�Ƨ�����C���,c8��6̤�et�\=��7Q~�vjƛ�b���4�ԏ�F~��@��a�Z���d��eW|T�feK����L�:��(�7<J;��9S����k���=��m}����'�z4�'@- ����K*��3��~���:!���c�>� #3��gݸ���s��XuVmbh�X�4T�}"��<��|���`c	lS&<�=���}g�ㄚ(���Ϭ(664'��5����EuQa�Dnq�'��K��S�����0��{�`Н)��^L�a�Z��l��tϕ 44Mh�!�����(�-�� $Lk�Z���X���$ ]΁}�n�כ�'���N���m��<t���P��m�U�bv��d卙�s{4a6���ʍ�;�{I�9�*���	���n@��E����s=S 8J�m�����k�o�u�|১����U�[F��A<D�9����3������ ό�k1�T��g�]��VK� �U�wD�[��K{PM{7��T��?	�e�8o���z�J�zN�/��QiDkS�n�x�n��e]_��v�a�]P;���`>�WF�o��CN���-��1�'HgC��2V�U��ӱ��l���+���v��%پ��9D�y�o�(qO>Z������,��*T(g;<���s%��'X{�g!�7�)��'�7p�q�<���z�W�o�࠱y,^8��;�����"�w����_��58��R0*5���m��"yJ��7�S��z��^|ڻ�|���mg�(�����d��/���0A�?���X�8�7��t�K�-�O�É�y4	JSR�"��d�@�w_�^㰽&�����N8a�>��\�^#篸��q����g=҈AOºQ�I���x�iH	 ��
��f�N�'FX��l�b�6՞��[�f�m�Qշ(�`�\�a�?u�>h��(A��2#��bm�XdP���wJ,�U�X�p���������a��E�!�^o�r��v��Y���ך��Dル-��T�:�U�J��SCC/�X�G�y��O��<�u,�`��tq
gI	�Q��/��Hp	0H��+=7|������қz�q X!���0陝&�����q��(f(a%�Y�<��u��M�������V�hx�'T��2�=̀��g l����=ŨuC �1�<T ^�Yq�X�f!'��i�8���'#��ݫ"ǩ^�H���J���FC<�G���6������d�R+��놮�QR�J�X,�\]��:�f��,C�4n WQ��Z@k�Z{�KmTT#�E��=��:��Bl���l�@�G��B��W�u�[�4'�H��0~�Wd������hS��� ~�����{DΛq��-�u�H�@���7#����wf���\���v�_�fO���[��#<����c�����9#��k����O�ac��4���6y��r��mA�y�b�Q|h��v�$�rp?ҰD/"(:����t���6{'ʙ�b�Mm�Mp��d�)'�Ȑn�P����GrtQ�򉁿��Y��W�{���L���m���m��j�&&����C��7AW��1�w�i�����=�G������.��g'=��q"oLk�����b���c�˸�4'�R�fb
�,:�n�e�A�Z�݁cj��HB|;=A�{$K�)�
��~��~xɨSc��y>�&�O��l�y�(Zht'-����~�δ�W�N��,Գ��V������o�
�����Eb����8Cd�/f�j�.�Vx��j�ԯ��ikL��5a1E�u�.;�����S��{�eQP�Ff�$�r����l��� G��H�m���W���x��Y��Dk���>�|�f�����Λ�c[�^�_s0�8c���#�k|�}G��1���E����@�1�t�E�rE��wۭY�ʏ�?����G!�̷��!�*�[c�G57I���2��pF)̷Ǔ��싻��B�*z�D�Ȁ�'5�KB,!��g���k��H�/���t(m�%�D��";�z�`t�f(���Y ��7U���3���A�r�������Y!6�A�N���j[*^�����lJ��B4��A.�M��K�C�T$�����YF)_��Y�7�;��kI;c�~�V&������9����&�V!�묞�Otvg�d����,��{���B�h��آ!��e�ʋ���)r���p+�� ��6� Ǣ���������x�C�בX�`7Z����~��d�+�P2{�6����������IlZЇw4�Rw|
�7#+��ը����ف?� ��0�}L ���lX�=��@1�M���S
f��c�~r����^����Cꓥ����@*�h�@H�!������^���۴!o
]���P��c�4M%�U.g�>�P��u�1�u�oȉ)#KT���4�p��|�s��S.�QS�\�
���)��WS��i�R�f�U�*�\�J����ۑW?���G��R�*����r$�E�~��c~��Z�V���|$qe��fsv��-Շ΋�M�i>^G�A��2%�~�R�E9��1��:A�]������2j��²�V��������;����kڵ��ï�λ�S�y���C��{�x�e�C���d��@D!�ȓTUR�I�
��������C�B�g<D����eiq^,�"�ZV7���)�9|�1M2e��%7y�K0`��;##E �v��0���Îo��me��jB��nV���5��l}(1o�u����P�k������ٲ�3�bȗ0�V�VNQ:L��L$���$$�`��2|��� �SG<�3B�QCd�Y<����Y�ü�ҕ����薝0v���ҕƒ��ů۳=[�[���.߃X��8�p� �L#H͗��j�ҜE�I��b�+�����Td<�E\f��v��re ;	��	}g�Xئ�D[x�<��EBׄi.Xt���7s�teĭ$��ڈm�]�9US ��N7�{��#�S���x��^��#C���d���G�RPK ���Ti�Z];�FyՊ(K}�Uj2Ҁ@��{��,�r|q?y3���I�Ū�#Qd��[�X������؊�Y	eE����ŵX��G��6���Ja	Y�9ݮ�qj*RɜQ,t��	�z�`�B�$u[c���DrE�S�Ъ�X��9�k�*r ��?���$�D���1��C�Ǎ�D9�ĸ��m�&,���'S?-�*��}%J+з�UMK0�ք�)d�hJ:ѡ�ܪN�KCQ�"f�rSj9>�~�������U7�l�ʼ���Q����]��Ì�<�҄�����d���Q�ZNe|OS+�yVĒ3���6u�Sz��}�ߟjnK��F՞��P���'[��±���WU\�
w�Jcu�UE(�--���AY,4k��9�R���oC���O�����%��,�A553&���R��uL�lyh^����9�
��dN��E}��|O_�/Žq�b����v�٫���S`�C
��u����\�����׌������m�> S+t�l B���{	^�Z�l���VO����	u����{��-1A�������r����o-��������L�'��%�?2��K�.�O�@���I�ʊG{��R�w�L����ᤥL�X��[�Cǹ7��\�5ŗ����Y�X�u����j5�����'d-�&��q� ]iƃzb��g��Q��>�F�?�gh�a��
����Zo�x��/C��G��Ć�Y��O��ACїpCF��D+��m���T֋=�����j�tI ���H��C�����tt��t����hs�O��F�Sٟ&:A�� @��2}�A�ɫ2W��t��Zyi��9t|R����BSI��96ú���q�Yww#�6�g�+[E
=R����>r��$;���}�z�����*��G_8iDc���u���k�A����f��6�,'U|�{�ZW�*E�ڔO��.�$�W��9e|@Y$S�ٍ�Җ
��7_i� *��p��_�`d�4t�S
�
z1��:r<��#�ly1�9�D���l�S��oҟW�n�8���Bݲa=A�em�W=��ll�Ҋ�o��8�B[�=�����ાW�]F�n_��L����7�:�
҈B���Ϋ�C�<Lܘ���"�y�ɣ��+f�N�C�9�¨�;91	7 �:[9�|��t�1�g���*��+ڍ�~ ��_���:G��+�U�61��-��	��G�e�k�j����J&N�ͫ�RL��L��I3E�(��D%�5���"�P!�>��|LL5��`,���0��&�5�����9̼�*��*��z�����͖D9i�*=ud~�1䣮�7�:��O�I~��3���=������2ؒ�4zu�2é�Ӊ�� ��Nx0������BI\F/�+��C��5.4�;���6��(�!���)�ԃ�*P�+C���+8���&��*	l�͘�;��T ���2�C߱�vͬ�@-�2�H&盫���2WS�B���],�zJ&!Fwv	�����m�<K~	X~��y��n�ڊ��������z	���_��wAv|\+���k���&Bo��ӊ`�z�o��F������+����T����{)�n�<��XM��1�n��T!�s��z{�"4\��)�J����3ř�'��e�Uh��2bK��&��:�lw|,�髒��J�:f���m�w�/i��&Ƥ�9��#���c �04�7�<���.PKY�//zU�Q���9#aV�+q�nRI# �;�<7�=��Q�KmywH�y� ��,r�:V�6t)du�VPG6�p1$�G��:��qC�v	���1'5(�.	���%�-�8m�|�@��Oo���Oc��)1^4���Uv�n������s6�/r'E���p���ƴr���ܵ�F�?���v�����N��u���4a� ��+�t�mӎ�5��AV篅޳�觛�ܫ�4��'���sý��#Hp���p�;���b����|�E�~��7b�(t�s��=p�#�;������j�����&�v�B�l��g�� �G��Gh-�$�B��ڄ�o�;_TEͳ��r�_�m܈}&^�����h[��3�z���%K�h���jo�~d=�ӭ������7�6Y��J��o���w,�T��s1l\�P��]�>)=2>�vqȝ���*3Rc���P�j'����0i��)�*���#�$��
���>�#��أ��V	����[�����Q^�ȋ7$�} 1	��EL������xyᇲ(5��2P���;�Α���-@M�շ�E���%sL�Әö����`]i+���tH�� �1�qg��Y�M*T�G?J=Z�p�zۧ��&�$�
ӌWw�0���i$������y��$y�����P�q�Uy��i��w9d\�;Fw���=�;�G?BWȕ �U���
�t��鞓?
"QА��N�L��U�K����)PwƩ���*�ٗ��p?�//�&g6�p��*Zy7;��й���E�9���2XC�+��Q( Zw���	z/�=�c}W<ˤ
オw�n_�np�=�!������h0-nv�i��86��n�v;���L�!|D��3���+<)'3� ;u�G�d�N2/�3�FV��:w��cRJ	Rs�ְn�D�"$��T�)��YVO�R�)>J��_�����6�t�d���yE�C � ]O�:-o+A���$���w����5a"i?�]�ݱZ���QC̃�v<i�8�{R=/Ӂ��O񻫓���,
ﵬY
c��ՠ�����Mp�+�m�+�����]�n�CXwdߋ+:K�DO�B�Fp}y��ACjpAq�ӊ����x��X�$*��kNe��Jg���*��.H���wM���q�P��s�I�@��ۉ����ԕ����Y�S^�ߍ,cG��W
��5�p�y���NN�&��pb\83�Ӗ�}~�m#)�?,��	&�t�6�D��P���>-K�G/炂�R��)R��ݿ�X^Q��\壩Ec���e`�D-�
:��Y�;�����E��㝷��fn2���:Zo��#�x]	�7����7���/�؁DՙU:�/��Z�������n�֨�k0���N�\
~���G�p��]��ul"�D�Wz�o������.����k �K�,�����h��5tP�\���]��'���������X�2��ߴX�w��D�澑GO
�Փ0���x�7"$S�G=3�~U0�#��Q����q��>5��*O����'��Rn���}���!91�5���r��̃�y���k��I���_�D7=��,��Й��i��Zї���S�ǎ�x1�}�3
�;�}F���E��ifȫ�nԑ_o��ʴ`O�4�m�T��<sf�O�G;�,]=��M�%�"�T؜��1��s�B`�.����Rh�u��(��>���K}l�le��8���y��vy�ꣁ~�O҂i�
Ӡ��x/'�����z�=5Oj�	S��4W���������?8�3]!�
8تy���䮤�� ���o�*�-"n��*q�0���ɝ�P����:E���m5q**���T��f�=�v�j�Y�b?k��3���oĩ�W�42�o��ݓ��+M�$׳k�ـ���)1_���a��5G#�X�}����c�z�y|:{fM��u<؄]$���>�h���7����qM�]�p&jVȄ�٧��,�17�zE
B�<�s+�r��i�]4���P�+5�����Pi�{�w^� "��
�����' ��<mW���KA���ta�� V���j�Ƽ	���|����1\L��8?b%����هo\�x�y\ݜ�N�+w���A�{7����d��j�����٢�G��vl�3�``9�9s�(K�P�h�0g����W��-_��� Y�:�C�nCX��]���Gt0lz8���m��/���)��>c�3.�d?ڗc;?��*�"��@�٧5�@��ϤƼ�V��	�R���V�w ��'�t&�r =U�<�b����l!��=}�0�n�;�n�N���lW�SK��W3����s��,��+�c9�����ݜh?����AO�=Zo���Դ��R'�Y�!�M�h`���������4��������৽��̿�򁋧y"�	/#������!^P��%`�(�{����*����q�
8�$giEqP�� �C,j�}��sj����£6�	�s��ҥ�ue%�+�-|�HpR��}����>óh�n��0�v
��/�:ϖuS��GԪG��� ?[=ڔ�"��3�0J�3���װ�ֲ�ғ)�Esk�]c7�5�%.�X�΢�������,��x[�|{�AR��V��$����G�n��d��YgC����T��4W�aB����RZl�����o�7|�U���C�3��|���ɨ���/ ��P����ƺ#�Jc��/`�#B�É�Z|�L�b�R�xd�˝��;o���W�ؔ���fb�%β)���$O��,�%��j�|MU���8�i=!�V�e��n+\%b=��g��ߧ����!ҍ��Rż�ݸ㗔ڞ����8H�{@�G^�I��7��H����@��NцQ-3?�p�=��&���� kt
q�x�wZ�ø���e�=��ب�1$	=�0\�8SB����	��~�!g�ӛ�(..� �Tߗb�C�@�H�0c��_��"�$t����z��,N�@4��9�9;�ZZ)�r��fe�1q����̠�{L�8�BJW�і��^�g9UդB�A��у_�NB�$Iʟ��`n2x�
����&�'�y��#�]��	5�l͈��Z���o�7�T!r��^݆«���|fu�t��Z���B�Y��xƇ����m����aO���J�k+����
��o�dĘ�DlT��E��m�nK�ՂK��ˊ�=;�	��C|_��e7B	�V,5�{"Kf��w��ǧ������4	WYwC�1y�0`�w� 0�}.�3;m�9�Da�=�9+���j��bw�JOQ ���&T�dM��ׇ�� *���h�4�X�״�Mvm������*���暕VV��T�V�id(��qZ���E~d�F�
�j���#��*��/��k�l~��
e^R-�,����� X�Ř�1,�ţ�oT h�e4G��`qu̇/��CE Oi��s�0��(�Lx�A��w`�<"-*J�1�I��9hj�F����	ׂ :9��W_?)9	Eu˂Y��m��5�o�����CIG��`�rg�H�Ͼ�_^�.�p�)I�^���p���i���=��`���O�B� ��$mH?�Y�;�'� ���#l&|5�[
O�;�����}�.wQ˱�m��߉`�5� Ӟv�Yn���Ay��� V%��E���E��~�H�/���At� �y�~��	�.�@��I�#���lSeU�~��4H@�6襮��A��F5�t���C�T��!d���:N�)|<����@=������J{en�ǌlZ�6�*�*��,�%��W-g��(kT^�s���8�0�iԜ;0K[S��5>�9��{��30v~�$6��|;l�9>J��c3"��3�;�⑲�#�u�%oqR؊?ء���� 5�N��a͎g�|���}���� ٚ��>��kR"pL�k���Q��e��9�J�b�b�M�[NDh�8qh���p�Vz�%�Zy4H!6�2������$�B�b�-�N���;:�PV?��2���9_B��mۗڲ�ώ�`�%VZ�1S��5�nx�����!ë��w�5wb=Y�2͚fU��k@y�"��=�ZPDEQ��hmѱ��"V�h򢲖�����{TU�˳��?�oA�}�d*^ƾ��\�{0��� �Q���$�m*��j^f��$z'�t=쨽xߍ����;�I;�ƂUt��O��s&�١�����EO�Fɼ��z��H�MM}�6��Q:k��x���۸�Q��rr!�RD�a�1Vܪ׉jL��?�D��ثi\C�\�N�*�҃X�3�T��KuJ{1(Sj�f<C,k:ݏ/Uy���&�z�<����'�����L�zʴ�(8�.�*�Hq�Ź�ҟ��9��s���g1�� תϹ�%.�DZשn1���ܔ������砆�!?�~�7yV�����p�}��hx"�������K�pIy�l4�}��;��C:�)4��r���! �/:#���,�&9���Yi���xu������/��[��_~�%�������<������!8�����yu0Z�S�y²�����d�tv���#~t^<u�e.i�M0��)�k���]��]5�PT����7�h����Qd[�Y�&�(6�tX1o��R1#z��`QSOWY�*{_g?�l�)��;ZM����7	����J�A^�j��{��H�~�hl(Si�� �%���ȯ�$D1���:c.�W�9���TT,6�qb�����;t����y�ɑk�ySD����W�1�:�����ʍ�n-V��t��ыNB�!��p�Β���3�&Ϛ0���*˙gtp��5�7?�?���7���s���,�T똇�G�r�Nd�S)՜|G��`Ep�݇��D!�X���H�UO����NH ߖiesܑ.ghJ��P�I��9��ne�k��d/_$HyXe���(�jU�*acFyBx�f��}�>��)b�;���K�Ў��M�`��({K�h���%j����f"=���~ou��7��Mo�g�H���э�!̺�=t�c;]�%U��.�ae�D��0�L�w�~6Z5t�:���*�>�g Hu��̮4�-�{G�K)2lF�?�y�Rb��	p��͡����Ы����Ѹ6�V�r[�HôΣ���)ȪOI}���C��� ؔ�c0r=?1��Ǭx���i��Q���>���^�Lw�^��H�ׂ��R%�����9�����:/Q
��Yuf�!Ȧ�pk����F��n �@��*�$(�1
�V4�Wm�p%Q�n@<|���Scba��D���g���#��4e���,�o��´eͬ�-픕��Si�
�]��|1�
,�CZG�Q�>�����/���s�Kڊ�|����]:��g�6M� r�'��w�s����� Ö��z���ݓ���2��C}{t��{p�k5�>��w>_NO��F�NBO��@>W��Z�z��Pֈ>>|N �_G��!�-kI;�&u�0�%Bp#�L
P�+�a�>4���n�g�y�����J�Ah�Wy�\AX��S�lnz��7˷t{Se�Έ�ƍ���`K��ϯ��*,z��߭b��m/�6G�!PǾ:��)�lFV�C��ȩ�V(9���?&@���Y7 ��ۋ�$��mu�hY�c�d%��d`k{=95�����в�`�]|Wg�q�� �=���ۀ9s��S�-Җ�d8U��VH���?��Iȝ�*�%SH$�딺䓎���"d��e�P�#S��g����q��n�Z�Eai�Ż�1�c��G�3��[|*���{bS[�쪦��1�F�<j)�H��ӲHf4��:��g�J�]�-2�\���oO|H�8Z�7��V��o��v⪪�cS{"��k_˰/��S3RbG�g&�̗q���U�d�M��*{ʕ��B��]'s�F�[��|&Ʒ�/2$���0;'T�V���&E����,��hg���،�޾���|;"�ᆔ ��,�7�a��&٣q��Շ��̴g$>�:ձ�yHڳz	q{�V��#6�sE�E㢴J�pI�#���L������d܆V���G�gJϑL
�n�阥��"h#G��-#Jע�J5s�#(a�ȹ�7��\	��a&!�{��#��G�!jAqQx�6��Q���(�(��L��C� ��=Dp���'X�|sa 6`=Ycs7��4�{ni�M��4���@Ki��{�ȭO0����2��j�ǗS [�)`�c���}a� ��N���ݖ2�8�̎Z��M�p~��l��VI��Ea>!�A7�XD����"6щ*y�-���]�>}�L��STŬz��
�S����p*?���2j��� ���sb ��/�0`%�Y�3u�9.M�C`:���`'s �C-�GCY�y(z&�B�v�<T�E�� �bBx	�M���R�㓋��s���|L��-�%yx-{��u�?G/��Cg��6�S� ����Q�����[	 UDq���L�6��x���!�x@z)�v*�@YKL�A��3�ܬЗpU�B��{�$(�)�s��e*^��`�ƓF�l����	��
�o�ց��wHd�i�IK��<=Y����}j�E��VQ�Z'[���H�im������`yr��k�c����zo���Nd#�R[uÏ�)�CJO#CadԨ#��"@N3�;����z7ά�ًji��&�C����9�v�x�z�T\��/��7׈G�����a�kuV{��D�.��Yx��H���7K�;/�"t�mv�,`�8�\o�H��h�]k'3u-���̟����E�M�#�p+�KF�idm�Ez�	t��V�Y�� �T;ٺ�c�	ᔥ�B&K��z��������]��$���;$�
�2Ѝ��^o��j��I�λyMK��6��H�f�j���ڦv
��0�yl�ˁ�Y�ST��k��bC^=��]��s�3_���%��J<.ɥ��k^��f��$���>ӵ�<�P%�Ìs���_�Kw�����}r+Yy=�%�� տ	4��tj�cS���ݬ�h� uS-��KE��s����6�t�)O�d�{RI4�F�w�O��Rbz�>�t�@��DH�j�����TV�ƈ�w ����䦻���յ��U��~ڛ���w���m!���u �F��R���q`uXp��u����:����Iђ��u�3}�$���DH��6����/,s
K��2?Z���+���۬�@l}���4�Vhv�xE=��@"���LCc^�l���b�34��X-��UD����Zd��u�,�U'�O������c�m���&D-ɍOذ5gL�,,�-�������5y;�Ή�7���s������Z{F:�l��O|{B�8�0��]��5�g[-���N�-���;���oa���o����BX�����o}IF��f��@3M�@�T��j��6��C�~��D&5Ѹ�C+͏k���q)E�4�l��@}G��_2��y�֢�����v�M��﯃�<�-����3l�E��ܿg���������`�a�)���u�����X�[�mHaf+�M���[*���s�^߮G�1P�f���v�c���Mq��ݮ���09��B��N�>��}�.t�1�@�`֋���H�I�*�WdVD*�UG���e�E�%Y�'��tZ�ua���~�G#_��U��3o�D�B�s��$J�<�u��QM��������^lx)�?n/�`�l���[B��t�G���?Y%���oWg�8�-��+��t�)���Z^����\ſ��9��>1!�\���i��6@���0�0�e&���}�a�C�gb��0lM��S
~���g����Ȥ�
����X*�*ី�֠M���w��\*��;�=��m�������H�=��C����Z����WW/���а,����ݸ_��+pC�qLp�����^�"�{Ȱ�<DVNL�D,�,#��
v�)e� ��Թp��K�뱗<_�b[��0qک�V���k�.��p��/���dHaD-�~��	%O1;р;���\Ar�!��3��k����:�k�12�A@79~���6Ł�z;�����"�)`�V�p�ho_i4+k7�Ӈ��(��z�K^�eB4ڜ~���ſ��3�Z�MZ�'�� ^����(,3�z3٧��H�㡬�8��dn�0��e�[�V7�8I6���p;g���)��q�k��lN�儚��6$@X�b14���CsAn٦�X ܜ�s<�J�x���=7Vw����1͂���r���S��=���Z�o�2GZ�1D@�bn���� �iSt/D,��uc��76u'��C຃�44�R�f;��Y:��שp��Ųc�ͪ��b,i}~�v�d��.��?B��¿�͠k�F���F�2q�~#���4��/�Y�&�=&�@E18 �L�A���0?�Ou���+R<��7�V�\C�q�ݻS38�)�:��^�L��Hh.f�,K�x����2yB�]�a����W�+< �/�_������Q%p���6\�<)� ����5��ޝN�նh�U������tѪ	��Y}�H�w�Ҟ�䗚̽}��̲���'�>9X՛]�v�1��
P5���3�,���hd��*�d��݌�Uw))i�\�g���]ٷ^&x}s��,��P�a�G�O��U�$�囹�����������s���X�u�Ͽ��m3��U��L��0'J���z���v	x(�2;��)+�s�}��r?�ؘ(W�]UzP����>�-�W6�B��� 85ڦ��!���;4�Y�(-/��B�U؈�[:Q$?�B���=,�H��%�%G�����`��8�T1A�x�WX28���G��Ö��������{">�NxZ�;bZ�t��oH�`Zѹ0?�������}'ܰ��/�Tz���/��j64��t �b�{s��0p��"�K�H)#x�#2g�w?���.��i�֐g�0�L�P�5<nBF_�;��z�A�'�`-�� �[,���qJcaI8OG'  Bx 0�1��e��$���߇B3����v]�����?(��M��"��>��5q���u�?��C�[5�����[��9t��m&���P�����4d�.�e�)LD[�K�W8��r�J�>�D����[5XR}G����B4�"!�ߞ��6�l�:�������&�S;ڔ�XT E�z�t6��Y�Ly�뢯҇��t�0��S��E{y��y����k��y�_���^ˌ��֕Lr$�eLዽ��1o�U�S99��!붐� �8�e�+��Z���_Ks�AL�v�v4%��ô:��֧a���|�#)���Zl��fC��.wTUC_�RO�}ԫ��*�'���\��d!r�N��wFt�yG�&5q���>i���D�+ jܕ����
���>&�3�]AJ�N��UlAI�!��8T��������鸖��l�i.�kZIj�g�y���ab�1�������0�z���8$v����ȁB��6�-x���%�����
/���k�m���D���\���;�v��	���n"͇$��O�T%����`BH/z�Z}w�|��~���z���U��8��[��w�b�:���dA$��seT.3��B:����}��#l!�I!��#�b�a-��������n;��qf���@	��H} O𛯡o��V{\�Rl�^`��B�E-��{u%����U9���R&�?z��{ ���'!�GU�u���R��J�����z��e����>�#�h�ED�3�';$ޒ�j�
`��$/ˬ����@9������+7b-�t�4h��XŞcc����4
}n�\I���`?L��夬0K�df���_T�l��e$s���q[�u!�&�#6�mm��(ŧK���N�}��I������%�4>�kx.�A�B!aX��B;�e�}�)h޽v�Gdd�0��I���^�q�1uǓ�տ�)Nk���}���P�zy���[�v�R>J��\o�&�#��|2B�>_�]H�l��#����u��Lށe��<*E��?��@�b�n�f�f�j`�9R&���Y�$�����uQr�������F�L��e5��Yu�'\S� F6 1�6X�B����i:�Q�d��P-l�oI�Ѫ�P=�#yp�N�A�2k���1�c6�T���B��c�]1h%6;+q���]Wxlw\ۆQ��q�w#�h��}c��g?��P:Y�4e;�p��x����f+�g�}�l����(2��Z�� �>F�h�XfM���Y��TЪ���ζ���*4�F+;~�GZ��1u�Ŭ^Z>f�U�u�T�KM�Z}�P
+.��$��+� �O��_��a�Xh�ϻ� ,6�(uⲉ�mu߬��a�����Y �"�FO���]�T�o��f,� ��W g2Jg�E���]����~e�B0h��ꑫ��1B毵&㊖~樿�oZM��r�;��|�T���ut���s)���h m�h�ɠ��/�,�"�Oz4-(0���}w�p��\���Nw��Q�{%7� �qW��bI��JƮ�~�0����9��hF�yN6�g⬄#[��P� Pn3�`�R��Y��,O`u�\/�9�3g"���\ԴEV��q�VvA+3���
7�,#��I���%)�:BC���t���S�>�]���`�;��U�pV��8��5�Cm���CB�L��=9w7��;m>v	/�XT'�I�˒L��v�ao���q��s�Sn�b��(#�	�w���KM-��S�(:�%~Ũ�j=��8$ǯ����2��y�̊�%����0A6�I��_GA���]?V��	�(��1��h�ֻw�z~��lVS��#!-}��R{�!\D�.�Sd�,!7�YN;=�.�Z$�{+/���PGN"*|��zE��֞����%d�v`i��s����LJ�@�-q�o5{~����{�΢��v�&[n)��`�ɩ`Y��j���k{�9���m	��?��I�.Hqri\����^�Flq� Sl4����z�'���N��>���ܢ�)�wdS�H���d���g2]IM�[�5���d�-�ssV�f�\6h|�W��+��)o����k�L����VFL�Z���.���������`�M��R�C���_v'�Z,������2�?i���9v���f�e�t�)��f�1
��P2�B� �������!���q����c+9J�2G�8�h�60d���b��>ik�m+�
f���7��,!�V�� ��̙���`��~U�W6�Ј2|�)i��@�Ҹ%�}G�;X����k��Ɠ;_�޽Ќ�v�%����yJ�L��K�u�#����tD�BG�I$�d��~���g�Y�r�i���F�:�bFG�$e���ż,�M�wz�cJ������k	V�"7Y�v�Y��x�S��-��l�L�d�xό����kzt���[��oW�W�8��'���I�>),L��ԭK��.� %n�9RY|�#��#�q�PĊ��H��p=���0WR�G� m"����Xs@���Խ9j�4��h*��'�R#8d �<��H��G})���ȏs�����:��t�X�W% az���ܫF9����?��`+�y��kc:V�$�b1���Z�d�E�>e]����j�	9Z"�g~I�I{�bN+�� �U8�7����'��A�G�����Z_��1�S��Y)�vt���݉�N�?S�ҀN���+ִG��ӢE���%��������ḏ�O����yq*�)�n+{u+���7˱&����NA؍K�Qյ�*H,^�y#7��r����@զ�[���H9ӼE̽��aC2�N^��r�A^����֘$�$ 0����x��'���٬E����9�_�Ml������֫;���� ��VA�B�c�۩��I�?�"����⅏q���i����������o(�h5�۾��û�+=8�����V����t��|��ե���k<�Oe�>L�@`&~,�w;Fq�Rf���j����IĎ#0e;-&�]�����Ӡ�����t�*e�(/M�X\��G+O<���f�����1=�r��e�Bz�$zE�����K��E�Hc���ŵ�Xq�]��C��]�$|�x�ntsP��������}���<G�R��A_�ɇ�
;A)|�{���(�Tʩ7y{vez���V]j��������s�dGR��ļy���"���&�K\E#N��FY����uS���z\�+c�K@���3C�Vzh8)�z�J���~f����":c�[z�\z(���,��0o�Y�~�@�4�AO�~���j����"6�bA���4��8�62�%QqHn~V��w�Zc �`|���B��p�����Q�9�'?D��Wf<��q:f��3�/���q�/�:���&4�^�o�8�ي��ʺΆ�_=X�$���<�|��n�q!L=���8yn
=+��5�tL�v�oN�_�zOu��90���sb�vF�G�*�TwN�6	��4�7ִr����V+_���Ӥ�X�`�V�byٓ%���z�^���V<z��U�Ԍ����0Q����5���QЦK�i�MI���6�sQj���~���ʥ�t���fcҲ�pɥ 7��b'C��x��c(#�ی��*��S[��S�-P�b���b�7�4���\����^��[8�m%�9�A��j�鮵��XO�K���X��YR\^��ﻶ�A?�����7�F� �gsK�6��D�ۻ���}M���BTUf�n�k�~G�ǣ�<�Ve���mC�_J����P���.��}U3�/�G��@Oy��3����{�J�N��gTd��^9�i�bf�	Z��r��
X�H՗��k�\��b�������i�Fp�b�`4u0�	���$�+QA��l�O>W4L�y�z��.'N���ْ[��=z��/D]7��壦�ď�����6CP���x=nf9�#���S���Q����X%�`�l����A)��m~͗{<B��WW�2���v���p�q�h�=nOk�Q�3y�����	F�Md��D��84C\��J�Pd���L��W�2ğ�#�ӌ���He�}���&�G�)[k�[��&C�p[u�4P�'���g�cbT`�Ȏ$�=��y[2��u��?ܖL����h���Gi��_y;��N#�G֟��& 8����p�n�Ў�P�W��` �E�a��\�
��ȅ{��՘TF�S���-8���i� `R��wˤ�Ioм�
��l�^�]��A ӳ��T$����a��S��c���^���_�l�1�ؚ�����nX���?q��l���L�Q P�L{d@*!g+r8/̺��l����*]II�}����x��1I�y�ǈ�
l��I�G��܄���C��Hw��l�U�QJۊ0Q ����WJ����(;�F��{U: 
�-(�G�{f�^�m�]���a���_�mB�����8C�8N�`:�U��%+�z�K���4��x3���.�~dXUolSX��k������n(�.r����:4�z
��Xԝ��$[�ͺ��qqn��Y?�;�2�p����T((��f�j�d�_6���4(�?:BY���4X�ea:K��f<5��{]� ��J�������N%��$P0~R�ؠGk�X�o��0�j��0֔�'�R��^1� �j����żu��#��ç��H{����T����|�3���<ҶQ�[�#�P�X�$�Da	�MH����?��$�*��"�j�[��E�yN��ڟ���gR-��:�S�Q�1�e;��c>���\k����3��M�'�㙺Ԙ�c]R�������6t����b�@R��\g�QAٔ�(�V��c�X�n��'�D
�^Ͽ����&��B
,|��BS�(U�!9��ӓ��n�A�~� z�C������-�i8����7�>�,x ��oF�HR9�ݢ��7uV�M�Uf�m�j�������D�m��Y����F�(�D��xߜu)�O�(F(o������Gΰ�q���`�ff� [�mA���<��Z+F�{�a�؏��$>��_��L+�̋���_I/��=����$�}f����;Q��ut¦���l��X�/r�
�2�?���&m�4�^���M��	�����
�,���`��/T�R����u�A���O��m�ۨ7��0A����j�dϋ�d:`j�")s��*�9{.�n&���/���t��������[z����[�yOn�6�Dz��Rޠw��ӹ�&!j� 9܂�u�ěf�{A6�v��A��<W[�%�r$%,�3׈c6ћ����
O8C{�l�S��x�#IЎ�z��:�����Ms����蓈Zͯ�au'�� ��C��;���R&��O�ҎI?'??���~!�x�=���R(�\�@:��8m1��-R��RE ����ȯ9���{�%�UA-*0}��	���&�.�5s��1���sT���n{�5Ӽ�b�Fk�]."�h�WY�0�����&T�s��N�RC��z��,�y��al��S��q��\5!�U�@�'�?7�ݚ�t5��t��1�L�5��n���#��=n�t�L$�����0��\�����<��\%�� ��7BK�?�klf	�5	m�ۑְ%X�e�j%�n����H*C����p����w��FXv�� �rXA�B��z� �O�2w�CQ���������8M
�v��X>�����J~��;�V��)��8GŌo]M:χ��h��g^.k�t|%}��V$�/�A�����Fб��	lRc�D�笅���)#C4�W؄p�3L$���R�bE�T�+'%��&�]A|_��<��Rj��c!i#1����r�/�Eo�A��Nx��}�P ���x�Z���|܉=l�z��YC%��L:���a��bүM� ��t�d�Ǭ��v�˭3x𾥴V�78_ �a���}}4�D��>1���0����ʶ���I�֧��R珢���y�NW�Ԁmz���&t�qi��Z��}���>I��F�n�`�:"'B:��%�}��ݓ�S����X�b�ޣ=�B����{-�ùs{'W�Ío�!d�2����N Ҩ���� .�>�/�	[�O/Z�m��+Ĝ���F�z���*Y;S�qb�Τ$s%��>戇s���������@fe�²�!'��Cf��ޓ,$%+?��#����������_V�����%f�	�8�ȱ�b`��BK�U����݇����A��&�f���~�ެ���� �#1hv�x�q�5Sw��S�e����>"���YFJ;!a�S�D;�؋��7�����=��*���<���5}��>"�R"9,b^�z�xU%W/i �� �����O�O��%Uth5h���:Mf�WOOA�9���P�2H�k�\�fF!K؂+���]G�<aAl�R�q�����pwVl�����kx���O`�e��������JO:�=���9~��m��
R�q�v�1�Q�ԍw~��x?��;.�~�JW~un-�np�7ex�[`o���\�����'���Z�t_k.i��?E�GP_dƣ��b�Ƌ��X���qV�X�E��R�Ʋ����Fƴ���~*no6�4���&v��L��~�r�g���+t0+��@�t�Q�S���� d�%N0�]�IJ�L�5M��g��
m�4n��`��	_k��e%��=8����!�G?Q�м��K�G��ĕ�\�A�6j!#��qɟz���R�
���p��,vX2R*Wa`~g���'���Q\:F��O�]�Q~��'��zI�;��t��ٴ�U�$��ޫ\��5��هg��pP�FU��ָ����ҧ�O #�B$�jd�������f~�����+��ٓ4;�����|�%P]G��j��ǌ�\�W����i܀{�c�_�2@ey��ׁ��p#���]����r�͖��pSB�h�*��6�r���y�P�&���P�X�[���Pڪt��vCcէ�,�|QT8i��u�!J�pD3L�﮸J���z.j���_'I/�Z C�D��b:W­�^̾��tƁX��oX0��mY9SSe���ԧr�ğ3
�*1�2��^#V�K��E$��,ĕN}�y#<��_�V6d�ƥ���ՁO�L�`�~�K"�$(t%�1�=|�g�B`9��;�H�x�X��X��[����<���b��l'a��H�Ϋ���!���Ä�-����}c���:�{��(ǟ���[���If��`��ŏiAyG���#��ًri]�x7y�6�i�A ��}�޻�g[���ރYK�nm*��P�-��&�r/[���n�Vs��GC{�o��B\!�Y>��^3�t'��5`�#H|"G�j��!�jD�mm�~�̹�p���a��o� F�3b�~s]���.�I$l�6o����� ������l.�"�֠�g�d��Q,fG��Lm׳��Fa�U�x�H��Kj��&*a[{�L&��,1r��)�T �<�6�u g���,��&p�m K�<�6���j.��W�'5���|�$><�C����j,�ْ�[hf0q��ݿ���d��rj��@*��@WIH�y���߸���
D8��nz
�hQ;2��ʳ[���kS�A����,Ӯ����+�rI6U���w黂7'4�ܣ;I$��z��ak+�0qZR>��D9VKw5{$�||�+>��x�+�((��q��ҭ��r���B��)ڰ�J�k�?{� �_2
'Ϳ�.[�?s��H�P�h�2�^m��z|��
Cr��v��ٰ�`�ϑ�
`�
��ؔ�L��KN�&����W��!{ʈ�3j�wK���d�c��=������|l;������&�Ԙ�"�r�W���R��P�o�Mپ�ݳ�� �K����aW�3��9��_K�==����#F|���r�װ+�,��l\���Q���:>ǊJY��]0��U��;2,�.VԎ�~�7mť��=R/�^��^nb�%��d0|~ѹh�n�Y 儙�b�31���@1�<�]i-L�6��*DP~�xL��Nt�C)���we��:�����j����+I���X�DX�x���*����sO%L�TLT��E,��w9$v���,{�%#�t�lG�|*�4��4ת��5��&l�5��*����F�\��u�G'_yf�'[O���~t,j��N���ӎ�kpO��S�86�������
\����:	��\���4�u�\(�,9�<�e�'�C/����E4�˺:�E<���5�H�~�LiH�g������x�z�b�Q�C~���[�e���۟U�XMlkFu#J��cmG�Đ��M\4�I��a�kf;$�����k�lG0R~�]h֋A�	�c�;?)��!�����D7��I�+Eف�ѐFm�{��FM[�����5�Κ[>����= �B�x�ri����>1�d�Ҩ*���?�oF�L�M��]���_�Ӆ,#_����#����k먻��ĄD�h�<�����M
W�!�K&��e�i�u�T@'K�me�>O�]��� ���\��h��R��rڼ�L�:1�J�ai<\�v�'���Jğ��J����-�Z���d�o�cd�&��G���P�1�_���%W}`��ڌ/�S
y�?��a��B+DDb<���/W?ii鲳�3��RðWBB3h;F*/��h�sC��)%�����	����?�����Y�v�XV���7_��� �S�L���I�:S���ru)WIZ���T��R��u8�K�*]<�&4V8�1�nm�΄���]�l�������Kw��m�����4�`ãkA��S�dQ0����r�ќ����[��S	2@G�3X@J������I�em��f�NL[`�-�L�hV]5U%Z<��H�(�@��Ƥb"�W1a�h����{o�X��4��];���m?�눁������}�[l�]HeDdB6���0��@k-x��>Bn�P�1z�����'���#^E	�^��$�O@����d�n�t;b\>sUHnD�ȧ���wD��C�|�����Kp�d
H�% �L'�.g4p�cr*?+\f�rJ����R���rq�3 U��t<uC�}["VZ�õ˛�7�c�#U(�ݕ��{��z�P�>J9��)iP���?|W�γ+sk�f�ī
�=��� ؎BCu����q@�9��r�0��е)H�j���s���_c�������&#�1^ؓ���<T6dʄ�Ϧ��|������&���;#{�{0os���#�`��P`c�BW���(F�َ�]H:b�&A4�AR�`s%�Ǐ�����{3P{MD5}���, �#�7f� n8DF��sX�?��5 �ۡ���S�fЅ"O�f���E��=����b�"����}9QA<ˤz޷��u��=�\~<�J���w�Z���[z�޹��.�0'"�<~'tP%�!^���c\i�}��.B(j����q4m�.�
�_�C�X0�$3~�t�~~��P�;/囇ٌ�EbJt�;=��)n�.�t[w���j�"�>�h ,3s�h{�V�,#�$��τ������:��>�z��Lǡkh�K&;���r*Ll�g�;J�1��m�����]�X�H�K����);h��{���2����I��[cD�`���_�Ӌұ��}^86$�ڹ�@�1���X���b@4=U�'���hvNx9�(=�/�$,�NlA�M�Eqi�
%�P5v-l��Fn�1B�w�����ML��ICj���������~R�B|~f9a&钤����k<�B�N4O�+��^����y�ۊ��`9�ik�*u��@<��b��E%�k�tY�0Џ��L K���p[Yd*9�d�����I���k�ƷCi
D��9 ���S<�`o��D?�	>�S�V��O[Ј�k-��*�[p�,�v8�s�\ߘ`ՔQ�Jq������'eL���#��@#+�khXK-:�E����t�+p8���h#k�����t���٩
VrlM��&�����G���"�Em��|&��ܻ1�i����+������/�{�P�H��
]�LUm���]Rk�w�!XAd��EM�zF�{B����Ds)^v�Dv7��;q�bWte��P|��)@�.�GP|�F�ϕ���w��Ͳ��"ג+i惔$.oM�Q@D�Ճ�$V��wL��[8-� �Г�8�S����g�P��>g&���S�@9i&W��W�	a	�m��x;���/��Y	���;�(L �Pj?'0]�79c���9��kA�+��p�v%�We���E��gf���ZyV�S��x�j�:������S�W����������??A��d�p�*[�����%����J���� ��S�[Cӝ��i�.qva1��ܭQf|��D�Vw�&��,T��ːf��'a�|wB�s�DO^�V0��(���n7������Y���R�h�˩�݀�x<�m�0�B�x)I�x�lB������6&)P����(Z��+���:s+3_f�Cbg��e܂�R��'fř�mz&X�)�X�&��VT��Ü����r_�S2:!�������>�
��+X����� �+4���y�Fz�h��knoN�~��D�?aMO��@6���b��h��m)����c�2�F�����p#|Y�u5�>�N�/ng�Mo��e�ʓ��.O��)O>�d҉�&��>^���.u�f���TND�W���g�Y�C0�	���E� �l*^�r��#%�h��H���c�'��LˎL�ڣ���`�Y0`	�.��d��Ӷ��6��E���N'��Eі;��4�S)<���N���x%×Lt�2�;���r=�ҟ]48�hB��m���(c<ޒ<X����t�E�H!P��j�;f����[�&�|�jg~�vS��d�U7˂�Hb���h_x)֟������d�t	ڟE����.���+����4����	�Až��3�;�ԟ��b���ax��&O,c��˩�o�6��j�1��{�7e6
J�@��$b������S	��Q��j�@�!rH�y�d΄� �g�L ���#���vBC�5Y���7�J�`�a�e�� e�����6�󯝡Q��ȡ:�6w��ACX!���E�L�hy����k�T����r:�o�9�gF���~��x[�����M�N�^�ڤ��`�O}���*~�>�5��lh��Қ��}r文�+6��G8^삢�]�8{vƿg.�7.z��y�&��"� 
4.`�ܢ�4ہ��\�P �7�f�y����NW��P��_�kf����U�
�z�h�t��F�h�����i���x-z
���'L��a�܍�y�ԅB�ܑ�Ïp�\�?�-7�C���ᔪ��ޚ�����ړ�@ں�5�r�2It��9�D��_��f��۵RW�$�2�XIbU_A+�8�a�m�n�G�(XE��ּ5�U*�ON=]�����2�Y�F���mq��d��-cE�j;��2IR�����	���66��v���z3�cR�d�x/�!^_��G�F
�.���-�!+���diyH�gC�L����7�w-��fNμlK̴|m�����p��G�(�R@�s]�%��o�h���n���������6�T��Z]t�b�Y���J�����-;e�"��{]Q]�P�)�T
P9�eXko;!��xv�וL�*��M�,:�����ƗfB���`�-/�����ڈr���D*�V��V�	r�;l�1�U��R�	;���Gb6ޣ�7�]���"O#���y�yx�	��L�m{���wS��Lp9\D}\@��AI��[�ɼ�y�3�y�i�@X9И��h>��X}f�C��y/���M��̐'� Ӣ3&��؃(��d��5bI�6Z���5��{��%p�f�;��됝#>�Kǃ�RŻeU�6�̳h�u�o�~�B���(���}�'���aG�N�%T�+"��O2[+�1�=G7�&���T�j_��W�{�����;�0h �9��-x?D%̈#џ�XF��t���/���5�s"�lj.����!���~���M�/�Ȯ��NR,h?k���v�:a�ހ�}��!��#�~�5����g�L� �GG���\�>L�ׁ�iW}F5����Έ~$)�
�zF�ޖ�嚧�8�����~|Q�p��A�?ȯ�C�Oh�s�+�
�e��Mm� V;|1�k̬�s��-�z+�(_��lx�<��0m����I��f٨g B�j����/�x�3�):��eOI�.tl:\�_@˵O�j�bۍ�b�Df�x��Y��W��8c��o���2�e*h�y���5l�uYⱻc(n!�tN�l�M�����]t�o��I�D�M�ިT���Ŀi˔�D��I�!_4��"H%{co�No�I��έ�y������G��'��7pM��i�*��y�� ~5^�c�Ħ���z
�-����d�?��_����F�4�L��N?b��ѣy{F�d��"] w���*y���خ�lo'�!f=FF�@��\6�ۤAX"bҷuBhMZkŧ[�8Rvx�I{+_�qX��%v��_�G��ݹ=3͈�3$ډ�Կ�Cd@�F|��P��n���6Z�Ҍv:�Kd"A�எh9Mf�-;�ka�҈J���q���J�8�n�ѻky+�B��AnǱ��IK�6m�c3�<[���c�q�ټ��$�1�?���L�V��R��,���[X��,�Uw��Jm�c�O�
9��g&��y4����M̃Rȅ��N�`�4X�;�e�>{���H�O�{	��.�Y�g���#��8�h���~9x`fC�NM�I��}"�=A9r��J���1�*2�)6��Vdy���9 �$�~B��W��t�-s�ad=��[�}�ٓ�eS'�(Q���7"ǹ�M��_����|�&BN�gڙW�O�? h7W������6�L��j8gY��v�S
����&Ķ-���k�W~�˦�y����y="�eh��䪜�4	\'A&���s@B
AJ�фGt�X�ҚfЏE����GP�4
����N<P�G��E���Wy���_���>��Mm�BV(0��t��IbΖb�xy��	�J�߽�bgcMe�j��qJ}(��wăX�Mhmm��62����K{[����2�l?M���R����D���6�D�:2��߸Z�����7��vxJ�2��}p�B�0�� �ɰ�Ka8�j��]p���0v�`�x��ֱ����^/�%�\z�ՋpOH��l����Co�o�Z���]���L��^�������] T��)��<�p�~P�M��<�v	�t@C�P;k3��.���NR%��Y[lLf�%�3@ۗX��aU����c2<KL����+�4+*UY��)f4��Ac޳�:�"�kN�{�~_�V���X�=��&�3Xn@�wqx�vlC�[�$��hJ��*��@E�N6!��k7�zٰ�U��e�ܔ�x��j��j��h���hw"��seC��U�K�]���ٜq��Ů`�'����to�*.^���G?c�$�f��`��p������E�4��s�f��D��hIY���t��Iz��.�ҩTb�!�y���*X=����>\�����J+��%1���e� Rh�o���\x�oʖ�xw��8�FtJ%�\U�vBj9���i�q��7o���+rS���,Ye��hnpxf;@��)2Q����Iϰ�^�eq� ��p�C#n�3�K���w�G�������dgc8E��7X��vy��~�?�,��߯�
w����]w�iP���.�ї�:'2�@�m�;ff1[-�eC� �@�>��w
.�F���'}o������<��0�;�[B�o�&�ד4����`+u�V[���f�v��w�C��m߂N~�|�\ +�5�YF.��L�G�{��fK0}�ۃ�r���Rn��ۨ�Nawk�Hw �������������Y^�6�Q�P���qz����������%,q0ɫ�84��^a�	mPB�,D��V
O�4`ۺo�5�rh�n��	"Yd:(�q<�EF�gK��%9�T��(m�N'v������D3��r (�.��N�7�2�|(����˓͙��C�
 &���'���5�b�H������'�?���C�����-�q1C��$M �ݛ�ƣP�����6�VV�`,?�1U�i��h�h����g�r��95��MB�6�rm�����`b�A��d�:�����v���z=�H�!�����PU­�Oɏ���'hS�;�cR̆�x�S�U����m�&���5[E�l2Mh6��sŜ_�6�?�:b�D��@!���4��â��u���,����#��k�n��`�F��|�_2 4~��o߸G����	���G�e���w��Z5�i�]�Y)�*�dw�Y��߰�M&0��pK�3UNL)nO����JEX��8/@�W�j�r���j2�fȄj����M����q'aP�~RgX�6=oJM(\�/��`�>6�W.>&:F|�I��aocM��ɟWpބ���3r+��i���4�F:5w,3�E(�>�O�o�u�*>��Ɔ�}��g�l\�1��=5�hL�ڝ0�:���EslB�
�� ���?9�dI������n�K5�Z�+xr��62��~�|߼˵&O:��1|X�t_��oA@�=�TƈG�2�~�P�O�%�e���N낎!��,IW�z��'y9V�P�����ň�>��2�0��^����&�RV�[�+2�A�*��LWt-݈?i5[��M9�?MA�׎Yn���c:"���U4�O��3m5��X��%�K����*�]|P`*���p�5��\V-%R���L�W1l��ec����CňJ��E���X����S:f�P	���@X��K�ۖ{��YN9cF�\qF���0�N�ܒ#�T�=�r&�D�����-�H}�'�q��\��N*woZm�b8eN!�V���]���I�r���:��DJ"�H���׹�K�������t�:$�]����a���,�wML�o��<�V���U��9�s�7Yt҃�u�w���j"<gTm[�&�Kyax iKE��vj��Y��;V�ǵ�������P}!�_�u����R���7���è��Cj虤C�#��ne�䪧�si�}�)��Q�vi���ʺ��r���h:[$&�=�u2^Nࡑ��"V:+|[�0�`�y���
(�f�Wߣ��2��Ӱ�{Q�Huo���	�ZZav��+bfH�Pl�f�G�٫̰�^橑�eWq(ѹ�Ѡ�I�"I3�?;A\���������o:�AN������b�� k�/��0��m�޺q%*��Ѷ�j������]��Á�5J�[{Ξ�B8��vs��O�X�2O�A���ʸ��+�|���-ؼ�)G�gl�w4��ƣ����������0)�4A�1Z�T�.y(��v1n)��F^IQL�(�K��k���s!~�F'�X����DTe������<����9�i�����^��[�f*	�� �}�kg%T����(s�Z�r����3�*�W.�Q�bM��S:.Qz�ȓ^�]���? �#��nk��`�|��=P���-�����j��=�����J��yU�c;���Bȹ�sJ�+���M��I�(��~�4<�b�$�eu��[�Q���X��T��a��+R���FVJ �;H�k�ٶj��v]7R͇�D���ky�=y��;gE��Pܹ�ND9�**F0�Śi�4�*&�h���}�1~�mn %�5X_��D�o��&0�*�v�NS�0y�쿠�۪K��d����/��+Y�u�����]��HJ����D $s ��C�|�zj�t���T�݆�S��U|���{�=��57��7�פ��š^@ޅ�R���:�B�G]2=V�4��.�8Bݣd�B��B3g� Y�����6�QL���=��A�G<Y�EӹCZLZvw�ݿ�r&%�\�^!w��iݜ;��9�R0�G��Y�҅�Nq����`�D�B׿ p>Y��ᜥ���R��%�z�"��G8尭�7+�*G)�l[`�j=�*���C&ސ��
q�SS�a�"^V^�=1sS����չg~�I�I�^'T�>��&Aϭ�j�UN\u���#�Γ~����Q���w�m{����W'	��w�,���
s!��|M�h�	o	��k��B����V��z����vO�Zt�]^g>�{}�
��"jMD����e�dDԾ����o�E,�ʣܮF��r���x�ȼ�m�Eޫ�o����p̰)!+��R	6��j>l��񳰈�����V���NHF6h�j���R�PH�.I�U�����A�ɲs��Կ��J~��[�A����g��}������	��;�Q	
A�濑tzy5�kT� ��q.Pn�q�p���%�O�����$����(�W�>���lq��jAo�"ы�n\���Z�<���dK�I���R�Di��li?��@<���R��
dr��PZ�1���LLC.����5�����`��ťv13�\Si-xwyu{���m���ޚ}��\ˁ��r�|�MO#��>����/���4-�3ǝ�A�<�l��4���ډ�����7ٮRڥN|l�ΑF��	D>3Y���Nb�Ÿj���QAK�Mr[��f�u-�H���`Ն/vY�DX�x�j����HR�c����=^|l�K������#��sb1α��%`ոs���+���{�P�������$0�C���&����K�j��J1�W1x��S��
���H��Kz��{��ޗL4ywG�eX��4����-r���V��(���B09SьE��!醀�ƹN�����V�9��q���7C�2������$���C�yVV�+%�-ǲjGG����}_֑�{Q�@B�lO���-�y��T�k>7Xg��-�8��[�&��1iX��5�vC��/�����Z�ֺU�Q�Í(��Z5��/ײQ�]�{@Q�d�Z�]���H�A�#�<C>��)�9�̿��L�
j`�#UL�L�K��E��D������1�J-å&�:�%`q��ჷ�վ�8cX��&� #Y9��i�Z߈}�B�R�ݣ|�2��?n"��;�'�͍�8[}�t�n�$.���_kb�0��Я��B��K���+a�6Hw@���L�эv�`��b�)�[NN#�%�YC�Z��q)��w����)��G��G#V��\4����v�!R�\0��	�Je2m��!�/���މ6�y ���e�ݜ��"�Z�%���`
8_w=<��������s�.������uD+�e�	��f>=�t�Õ��p�IfYaLC{yv D��H�
3ӡK�L���N��,x��s�?��{�Z2�{"v*���%�rwW�h�v�f�u[4�|4��t +¸����	I�!�䘥µ�� �Ĵm�r��m7 �����t~���t�j`~d:���z���0{��h�0���Y�� �E!_�+w�<�U��TE���>,2������!��)��{�ӫ@��*�ɱT�(��^R{ z�jg\��d`�km=�i��D�_b��P��|N�y�e5�riÛ�Ӥ~/�1�+`J���S��+`d�F3�_����f�z��c���Gɂ�Y�1i4Sy�U���W�H`������=���0M����cw�>�Wz�e ���0Fe�;�ڄӾm�<P��NyuR6�������4��GG������N4��1j���>r	ׂ�p�ku��w� �{��4g�,�w�i<V/#�{�;���fh�j��x�]��Ho����u��22b�M��SQLnyI���}����=�"�G�H�fc=r�vj�?{R�	�XTj���;/�X���������˺U��S�TV>��^��������,x�02>z�`�#t	γ�i@��y�s�dl���S�l$M	kϺEH��-2Y�{Ӏ���� �)��W�^�M^�c�	�<­�OC��<$2�d�D�z�&k�ý��pyn:r'u�/���֋����9</�&_m�Oh��e�c���	��^J���#Z�����ռ����|4���DLY\�J���:�$c�܃��o��5�~�0�t+I6&�'˵w�Q� ��d 2ԃ��O.6&���w�ǈ`^FyB�[]-�s�xĐH���5)=��Y�@[n�/+����B�@-�a��d<T�)A+O��{̑�X:Y�K��hw�_e->d�^���~��	*���Ψ���b���}O� o�2�$�m3@�Z��y�=7��轄�P�FB٭:�Ci+m�|�.���(�t��d����u��U��S���!'��_җm�2*�7��n.q�@��%��I���[N���_Ӌ��rU=�z�u�b𜩊���J�\��{��E+���
: 1��_����װ[�G2��!4���=4�dY��)c���Xk6��Wױ҄V��޲�9V<��&f��n__O�=���{�738K�rn�w��9�NKP�){���e�v�� ���K�+��y`�]UU+�,��G+D�O*g�::gD���FR̅��O���J+�� Z9 ;h9�.���w��G�̸89�����mRz�EVC�����u(Wж�����l��� ���?��L�F�N���Q�s�bYgjfM]�z���D��7�	�?��椭"���EПU�ב���R�Y��B��f�n8rq�H��G����vij����g����y47R��e^A|$� '�_-���������G�w ��(�|�¡~#s��٤v�4�x���k�_���ZM؉&9A���7�K��'�$),�d�k�Rư@S�/�7�
�� ��#����4r��Z��o���k�9+[r�f���n���3�� 1�����p�}$�	���kI:z+����xA;�OsL-o�%�i��50E$-�R]��}�0|���B�Il{EK����qд,����CI��{�啊e"-n��R�v�~*�ft��PH�Vq;�\S���z�	%g�{�읏i[rc��V��V^��K��I8`��R/<e	�b�<p	��yzrZׁ�/�E����Ij.�0�M������� �E�=�� �x}�^����S��r�_p�8*n�l������Jd��k�����i����~{�2o��;u���
�ӊ0�4�.RR⻆-���&��u:��HK#���\7?�@�6��K��\�Ա]�w;���c�C�U�C˽̱�t.�����ķ�j�̗}���L�X� ��汈Q2K9���I�F	)=�19)	=V�$d>ك�ԍ�9l䛟�`�l+{�[�k*�m�p������--��yf��#hօ��n�`^cWƢ
h� ���D��7�_���]Μ�+�0�/vφ�Y@��Y D#
���>ȗD�(������a�7Y�����7���5��{���r%�D�0��>��7�--�?�$�F	�B͸�f>�)����ii>T�.�)�����[�p�"�\�ծwҔ��FG[T�֫Ӡ(9�Ӷƪ
<o���^*��D��w�k\ Dk��N�ߋ;�BXA���!�n{_��� (����-Peu���9q�;��� �Ytڋ1��Kԑ�:��*:�.#��-��uN�I���o��7����OUDq_���%K�hA_X3�E�I�ҝ�ndmY�^��c�;��;{��}�2G�G�k�y�渙��X�H됫b���Xc�0���!V�no��OQ��w2��(��?Ug�iP�q��-�X���;n�FC �p]}!�Y�T��*����މ �<�+�c/8Y�獜j����P�Nw��;r�?� d�Oޞ�69|*�nP&+�i9 �D�Gv�	�v2!ۚ��߁j�t��2,$����@ w��Ѵ��~F�).z����eM/����� |��)ʙM͠�A��]-�!��MOb�}�B�����/�؎T�lY�~(��9ޞ�
��ӛ��8�=㣹�sj8�O�Dh�廵o��w���Szz�ő��bE�K��e�*���W;Y���9em��(=�v1o���a	(I���>ن���TE�T�o�<n�P�6�a��Pu�}H�Y�������Q6�Hs�R�Oj_Z(}��鱺
��T۸@m�;��Yl��.�Z�YB��%T��C�8��?�����V)[�{/pf,Q��<�����c$��O�&�:@5A\�F��	ݢ�	1�Uɦ��|����3��y����2=g�H���4�n�u�@��5�F N��M5�U}�J��{J��n�i�\`ک��p�;�_�0"+/�X�!�ᩂ��^}Ɩ+2Ԡ'��F�\ݓ��wRU��V��Z��������&�O��w��`�W!�t��^9:�C)�Xoݤ��"{���g݆1���(;Q$C"�J�X%���Џ�~��+f��\t�UX:������KaZ�UHޫ~EYm��vU8Ӝ�e۽q���r�(Xܙ�7�9ǚbʭ�|*��"%�����$o)݌Y&���İIp�|9F��㷻��|�-��66t��m���*gs��"" �!v"`������I�#;{3*�6c���9:9���uj뛍]�{�����PC��4z�&wz�y�#�L���>�_��3a#���7�!a��Y�a�M'���$!����ْ7��F��F+�xV(1�S��A�/�B ;Ԑ&4[E�I
��=H�a���v0rƸ:�לҜ����Ф����)to6$��g��~aè<[`K�\}�~�E6L����ow���d�
@�?��肱�oDV��� -�vP`��(�B^��_�����3dh���nS��MXNR�\W�$��m1�^q<d����R*ⴰ���x��s?qR�n�0�*�ʭ;�ZS�O���f�:3~�|0�rh��e�f\T�Z)���o~�3j}�Q��|�V��(�z���8|���TqّG��-��*yu�Ҭys�]�m��n&��l��YŨO�z�1>��wUW��-��QOyp�(���m���ޟ��'���ܺa\��X׊��
�嫞�����&noX�C�[/��C�K�?uU����1 ����7J�XL������UI!�8u�c*��&��Q��j�%��OSL�r����FK�WV���^�@�-�����-�j�<����iP������W�.�xi�|��N�����3/P����s�1��^��������+��X�-=*gDMR7��nn־��]<�6�{]��I���7������B��q����n�t������˻ʌ2�kC(��NC�繢��&�IU9����XE��M5�fl�\r䣘A�x�q5�V�;`����}�H�ˏ��B��(}�is�>%b6�I���c&6�lsMx4��I��iN�v#��17��j����t�sLᆅ�w�PM1o�z�_��uM�î֚�F4aX:��W.�������}ɪc�ӭ�r!��o@Z�j~�e;����f�=m�CT�1�VD}i}��=,�� %��~�(�鬀��GYX�	�]�w��ŉފ0����r�93��C��ܒ6(P���mqL��8�\�A��6D�0�y��n�F�v�FFus,��e�P�Q����,������c��z7F?�A�J�x��'��^��S�Ȯ�B�r�s�W��PX�;�������¥Ҷ��ì��m�nI�6J����h�'f?�l�9H�[S��>���a8�F�G��|�����,���0"ɓ+(¢�Uj�7����뒁#�u���&Hu�T�T4 ��qQ�6��Y>��3�k��&2�� %�0w�A�P@����T�?0���.�4�W�E4�������5J> ���[�o�J� K��$�~h��(�3����R�=��H1m`�C�#�nD�@���2��~��d� ݬ/�?����R�pd�n���RH��k��Mg2���1��*�_��th,j��̌�o��z����W�k!ж���vV:*�uTZV�CX�.0�>�pV2�_c��P(�M[��11L3�bE�"x�ID� _+�?�w��6�1�9ȡ_�<�[�+K�d��Cj��3c6�%�>���eکa}ǛLČ�^Gk�0w��X
���^�������E���!���>AJQ��h�G��R�q����>���@��g�� �+�#5��.�BF�Cȋ�����=��7��$���NZ�:C�*pn��:ӗ���%2-���41�
��N��a�� �ؕ�Pn�|�~��7�юo�&�˨��[��:�f��kxT}H?�<-�Ͻɧz\�=J�����[��T�|`�N� ���ɤl9:T8����@�b���
���+j
1.��<W�(����K����woY�����	�|���S���\e�^�<�&n��(���{ד�*�5.Ţ�l�9<�2���!acPǬ���OO������@���7A]��|�`�r7���j"�ۼ����,���J|�5~5j�8��J�MUJ,T�l���$y�s!��_���@��G���Ag����Ԁ=N!���h	F�+�g�h����8���{|'N�7?7�$O�&,�/mi�W��Ty���4F��z�:;�K����]��q�o�
�+֓�1�yb�H�LA�F�^I��T���%�6/�m;�g�@N�Ս<{
����t�w`��mQXW� 7>��|����0�,��U��1�/���R�D��2��+��A�jJ�#D)h��-Wɼ
As�WԔW�`�5�� xa��y�M x��c���a�a�b:u�v�5+��
^�����H�kc͂X;!ƹ�����-KÃK��S �k��d�{1b���񍈦�X�L�u�@����Y;��2�"�rՁ���ZA����ȁ���`jNg�4h�J�v .F����\����C��v��v��C���)Om��}�>�X��,�f?��.L�j޺cX�9��Z�zF4��j~<_$���L��k��a�Vu�9Y��4]P�a����ǚ@���x�������F0�oi��W'Sr��n*h�m�;�<�3o�/���'S�$m��.?�ڭ�O�
68w�1� ����4�Jy�~RP�B�p����|����Q�N��D*Lw�̕>U{���T%Я��vg9��p���9qT׀��f��l��+�v�.���Xa8�+Cꚞ�&��Xggbŭ��x���׭?-�nk�ܳQxV#+�c�5��䡔��Tn��S�]Ϟ5�����9�;��6
�m=bt���$3ň��%�N�����%�E����=X�K �,I�����H ��g��dpvT���>��P�G���ZRL�2e�����x?��o�S�P@��ȴ�W�E���^H�	�!&����9z̩�a	n�y�?� 6�E,ڎ�?Z��Nq'�[%��L��P��K%�_X%�p�un�����G�{A�谜N�n1��?HUs�d3�T"��g��
z�f��{o&��u���Y��e����Oy���e�!��9���T0WY%���S�5Q-<��)7�ͅ�9"?���(�MuT� ϓ��Xs��w�_���	G�>��f���6X��u��P`���C�9�;�e!v}eviy�K�+�׬C��~{����3�( �	�ܚ�;9�	�\np�� n��JN<�m}����̨��&M��� �
��u��6$�I3��%��z���T^�q���X�&g�(ȑ�W~�� Vsj�����,�h�ԫ��E=%�q|e억����s���sŚZ,��}x��w,p�B)����ù|z:?˿���w���S`��B����-��z��@�p�!��,���+���/wo*M��/�7����8S�u��u��G�r���} ��1��K�����0�.I$Z��di�M�b�<�}�y,�$Ɣ��r�VC�X���/C#��3�4����y"o��B4Fy�Ǥ�Ο�������eS�ݿ߬�>te�.�`��.E���۶|�ſX�,�ڷ�h@r�bnIH�����@ø�/l���Pf1a�i�&�62+��#�7�3$�#��&�z���u)^z&�a^4�<�3��ȩI�ݮ���Khar�����k�.z�N�p�~�/��/\j^qb�>h��e�x��M�2�� �M"Lt��7��ZHZ]9M��DF)']��g�I�_{��Ҹ�x���>�Д�0����E�@p�%�]y"��e����UQ��݂ �yhi��L������e2^<9Pޓ�C�͑ٲ�h:�D�?`.r�O��,�O$܃fJl������,U�]����f�ң���'�&��Z��#���`��Y������t�7��b��
�[�<�3���cHFʄ.N(�g?Z�.�V�I�2�r/y��=�� W�h�	���`La�,��Ė]:��Yč'�%h��[=3��ie긼�[�"�ϽkQPq��8zA���)��*6��-��e1�Y�}���(�
��
xZda�n)Q9�#�6��ռmj�D��]���0Ƽ�q�P��چ�oa͎.Qt��j�۫U�����s����z+���~��s��i�.�K!L�[��n�~�rK㭑�E<"қ�J����}���C�R\UB�,-�^d��m��9T�g���P=B�[���Q
C	�8Չ�rR�誓6-�%_�7s�C;���p���K#}� �t踼�L�!δ!ƙ(� �=9��an�1$N�J�����Iy>�FVv=]�v�IK��I�b�\8ݻ�f�_�+}@�������pU���+��:��?#K�̫�d�5�����+��I'��e���fܾ��
���o��F��I��༳��+��(s,6H%2�r�= ��>X��u�(7�"�Υ�C��О�'URS�`ƒK��y@����1.��/F�1�G�8Q*ױ����ɗ7yyZ�Z���6�/7 -J8��:�7zҍ����{G�N�zZG�XQD3Ի���y#���$1-�녑����NS�c��.����X-��҆|�j��o8 �N���T1%����*(��H�K���k5���N�t�>6�΢`��RsM�i[C��/��������9r"���T5X�K>t��鞒�܌�CC>�(
��in}X��T>�<E{u��)ލ-�~�u}�hk� ��
`b�e�|�� HG�D*�:m4�V���%ٟ�{c��)����j��K��'�*�2gr&2N���C�k��gx����������'g9�m�|�(_�?ԧ������O��e��E�2�k��k��$G�X�d�j�V��?9�΄�
'�"���(xB��@�H
At�>�2�F�{�:�'M��ʚ�]D�|گg|l�/a����Lٻ;l�nKh��mM��Rj�k�J ����`�j�>�X� ��k�i���]<��Xp�M�r!�r���T�x��2a@�N�H/:2F��D���E��׹O����K9%[��=s4F�Z!��{�Jr���HR�R��l;Ƴ��z���ÞsW���'A�z*~t��	,K��R�`(���E�:��ֲ���o`Q)<_���dӓ�0�'r/*��p8��!��?��fS��E�p����X%\�uv�1 �U�H��n*�m��V�z�౴; ��+�!���	��슑[+���B�(�2Hz�Ш_���Y�ͅ��g���	kQO#Æ��r��#ip��u��M��_�eE�/��~G�B�@$�I�P�B��������*5S��e�5��C�/��o|�4������-��Gﶣ�0�(��q��hV�H4��:�=���7u�Ƅ�ڢ�C������~�
�oM�L�S^�a�����oX!����o�}%{�<�����u(Z^x����8`��i������Ԍ��y�Ъ��0~w��Λ���_���ׁ��~�
��0��0R�u�7�>=�TN��p¾�/�_<��Ml��~т�ߞ�e�r�(0鴉�snrg�{5�)�t�-�iY�:�P�8��V�;d�p 5���Ǟ�B%����P��*�K��/U;��bC��Z��&ň��ĈEE{Cu[�-+9#�V ��e�$VƒU��V����<��F�߼i�%�ʂ�Ru��郸?4�����߽Vk�,���OX��$�BNniؘD��6*VV�_vTs���T�6�B{[ߗ�^�:ӆ>?�x5�r����>�I$��
���D�Uey���T���7Ͳd�?�9u��o��&�g˚�]�L��o�˹D�����_.�I��	��'w��T�x}�(C�^������9�N�����7�SM�ZS�5D̅�Q{�C����C>��Ѽ�`��ɗQx��3��Ã`G�*~E��ot01{����"�޷Tj�v�/'U���ӦQnNO�B�\V�� NI�α�n�2��Ƀ��/�R�6� X�v�}#Xz�$��V�o��c ��1�z���a_�(���vZ�.��,}�s��ˉ���{���|�`�/�ES�ts^Ǎ�ނ�-8ԩO�,U�r����6���g�`Wp�d~@p>�s��"�pE�s�����ȸ��lH����r��T�➄�Ǘ  L�+R����SV�}��)֟I���Ƕp��Mv9q?ț��G�ȧMG^�X&�R�A�4<Ԃ����V����lۦ́� 3�[暓&p�a�C�
��o2�蠭l]�l�=?��@��~=�(c �l�N�h��PV
�Ig���XjǬqה���Q���,�<������l ��K��]*�Ɂ?V�t���y���$K[:k<�T�8}R����(��ɧ��i(xrÛ1wn���r� ���e����0�@Y4�6��gD�IGw��U��X��9hs�lY��kDFj˄"�"d?>�`:vV���q��8�Ib�6Z�\����e����x�D��84�L�VPM=���z�5� T|:��WZ� T��v��ܸ~��^֣`�T������r����#�Uh��_�7 Y���D���tfU���@�E�a[�B���X�|���ze�* U=��sѭRT ke�	�+^;�}�7x�i������7�\��	G�0����魓9�u&��1�t6���g�J�#~��u�G������E���f�\�q���-��ù'1j��&�|���Ƌ�=0!`K�Y��tBP�����9����#�{�7����c�B��i_F>�#`�p�P �h��'r�^��C����1 ��z��G�LZ���X�U���	��u4�нu\�ws1."��,�.�2��tm��������F�y�̉8�_'���Y��g����uX�XA���mt��ĴTXJ��O�]��	�*P.�8x������]�4kV(V�@��ʄs���AF�Ԭ_�S�s_���� �n��3K�g��ٶ��k�lP�Ђ���SK�o�WM�ˑ��{&�i��j�Ŭ� �˸5	��m���%��ۮ�"cm��k�U�
+�ٺ���.w���2�H�:���Px
��)v�.F��Xl�]�V	�\��b�rF{	qj�Bơr�� >�"z�I(��X��+��>8�����7!���<m���O���u�SX!Z���R	���y��8����v���@iΩ�M�vؖ���$	6`��X���$���:[�Lh:jP8���H�����Me��g|��{��iOh~i��[Ł�$��l��%-�.�����>I�R��P�჻����k��(���(��6�ZMR��!wh���W��<I
�!6��]�B�t��D#hVѤ?��-@��&X�����P|A��~��Z䊹���	a	�"�e�,�?��ѐ�$�f�����?N�D6���'Ȥ�P�?�Ϩ�����������[���`��YB�ک��;�	�#����7�wD����V�5��J�;@��LZ�_�]�O���, }�}�a�voXޤ���z;��ϮC�Lg���!A4GF�i��`�貨��K�nOx"|F���0��b���s��R�3�vY���C�V6g��x���1��e?�O��^m���:BRE)Dg�(�H�@PY�g����M�� G�mx�`�mgaloOɹj��#k��Hյ�N߮���^�5A/��0�,��9�	Uybj�֬��_����ga�s�B��H�S�K���	6�F�ɍd�nw�}A�&#��]�?�Q��z���~mm�(Pw4���-�)Qe�,��g���^�3��Ys~J�Z7�Z���6�-��]r	��p�(|�L��f%zn#���Gb���d�$�q`����$㳑�"$�*���c�ㇲ+��ƪ�R��?��V�Ӂ9rb�R��&s����q���~'�8�i+�e.1�A��	���Ʉ(�i��%#��)���KEv>%^I$r	�q��*%Q�D��ڤ�N�=� �N�GT� g�d'��@���x�:W'��j*P4� Ryb�XH���\�_(I,��J�d1��L�C.��!�i�0�^�tb�I�><����P-��Be����"��'�ie���,E�UmC�h(}��
$!�/h]Wh ���?�h���>0K0#:V�L���1%B�=ٍ$�4�66�c���ۙ��ђ"�T��"=k��[�J�Q=�?�����h�Q�J�
��.�<և�ț�U������_�*E�0���첍�R:cKd&\ڃEkx�B�~.Iv@Q�T�����tc��ԧ��o��Π�Y�9��&����0�؈U�Hwh�vE�)
��D�֩o���i��
M��|Nf����jN?"�����5�-��Y{i����D#(�/d~`��^�(���hH��x<AS�_�e���a�g�E"��)\^4��Qe+��Q��okD{�V������?��:U�K��a�����������a.���i��Y���d�f���O�|p]M���-Ⱓ�n�v��s��)v<��T�֮R�^��P�X�����U�sQu�.:
b%�+D���pƨ���$]���g.�:ěy���H��Ş!�J0a�����\X��jQ�j\�+O�Q�p$J��?���2i^Ȧ\�ӏ���s묝
����Ȉ�+�Q��*�%|(x{-�t���`���P��#H���,8�Јp%����F�Z��(V�A7pd�h
�ԧ��������=�&���(~l'�D.�#U��J�CB�f��/�I'�Q+��I�|#���/������9������?	���GN`6�����G z��!�o�p��;��!CAV��)N�0m@Ƴ�I��_�o���E�.�ے�����=�}�����UP�m4b"�Ǆ�o*v�S���8��Ѐ5�>h��&��1��Y�v�#�Khyzg��v�Jq=�)}|G�ќv�O!<1�BkM�����</2�g��2z|Nk�0�w��7i���_zH���`3K}%���
��I�K�^�H��ZK.X�^��m?cH��6JF�8nl�>KEܟ�^V����\l�)u	�{�d.m�n6��5z����@�Ҧ�ֆ�R��BaP�&�:@o�S��T��婪S`O�t����;����N\�T��NK��ˋ���\$�Ma�<15رOC�ǈ�V�\|���:
������32s�[sv���V�lP����hf�`�4���W������f�{W�U!��4�sbM#�S�|0����,aNzb<i
�c���_=gRT�E�ZC�ߡ6Vs�}Xvrw��t�
hk򌖦olr:�����)� 
"�����Đ�Y&�҅uP�3�-��g^� �������by�f����YkW���>i6+�y3�I���x{`���ڥÁ�C ���8Ș�HHӠ{6R�0Mu�Y�i@~����Y���w��K����蚙���$QA4��#��?��
���ܣ�NS�~$�E��kk̏DK7i���>�D��ޕ� uhb��^��Ad��+�=�k��팡`����= aGv]?�Q�Lf"������Ƴ�L�n�����o���z7��,��X\��3��_���|��g���K~���&h��`?`θ�}T�ö����d�^�϶���\�C�	`!&B�^�v�
d�P�O��Th��#ㅜ�l�>�0KR4h��8Y>��gs���N͒ �n�ާsL��1��  �a�S%�8�e�(෵�^"�&���/r6y�c���/�Eq_	�.>�j�1~�� ��fk�H���RV?FX���	,��'���oS�?�!�0�F���%��3�W�M-@�� ��75Ȗ�U3�Zɿ�'?2��������{���''�:��F�k�zt���;-��?�x�˒��J��.�x����¿�?�A�!H�<(�at�1E1d.�6b�n��E|�__��w82�R��x����j�B��`��O�*��l���N����
��a0�"*����3�����9�;�4 �_4	M�ɋ1���-#�K��/�S0�9P �ca��n2��:!����	Y�B$%2VA;5�����Ķv-+ª��Z��5HJTILp67C��4(�*IM�7��������{���/8������X@� U��'wz�_�h�8�h�����D_^0����n������Ixo>^�a�H^;
�VJ5@�X�L>���d�:K�6�#mQ:�CKl��/�'��pd�ׇ#��64��{H[LU)/���O��P����z��N�lѤl(�4�Y}L{��`�S
�)ۓ���'�a���B�h�mZ��%�l�`�W�_�:�# X'�M )a���P��� �0�V{g=ĥpV� u+��$�1�=�R�������%8�l����U���/y.EpKj:�{��{vӝ������'[S�y����P�0���t�Կg�4�L�'_&4K���j���Z�T{w{���.v��:�e�
���T|?��Yݕ���9l3r Y�98=�-�:F���~���Oz>�1߹o�!t`�3�|{3%C��Qw"Ø��&��O��.�����DC��6t���� ���C9{1��_K� ��/:��OƖ��ZH�&��r�=��f�<1�jc��]�Q	�.�uH�9��,p�6 ,�7ED1EIc#�]$[��d���7#�M��$��j�}L0ƃ
����]�t�3ܥ3��a�]C�S�x�7��HuhVd_ٱz7L�۞ۤ�O�J�1�'y�K��Nn��V��󸍉Y;״����u-�v�aũ�8K�s�;�����{�k�.�p�~3���@�/�����I���'����9Y!�61L��囅��ʉ5�~�zppx6u{	sw1H&���A��3���0	�y��#J�5t��*{�QS2���ѹ�7ϣ��E�H�[��DD&0�U�7RZ7Y�r�.փ)R�s`��1R�-�c�w-2�3�=��L�\�|��E!=���!%H�H�+����:A ~��պ�����I�$��xgz1g~G�'��\%�%���O�:CƎN��/C6&�����1�G�|�m��$�\�:���Dm�B���UciϨ�)b����pw=���A��t�quzH��ɛ[(�0�I	���o���� w�� ���'��e7���^5��+�h�I�f�jJ�;�Jh��6�O2f={ʷ��Ҟ��xmm��]����y��e��~�'������}�$�\����hU2��Y�:����]�_E��a!�TPO����Z�ui��3���6%��T*��/���΍Qq����1ɥ]��Q,k��J����������,����c ��<
2�u�ʝ d+l�Mm��/����C�Mx���)^z�7|�j E�7L�u�M���}����^�<��OO��2���,"z ��]���H�t=�N�>�%Fo�vW�Dx��P��u�9� r���!�u=%\meIZz!�]����$r�׽��݊S��h�Gm���yc?�l�z��pG��X}�X������Pi��1Ȓ���ރ
d���,�59��6�D�
R"j6���05:�#��4��*���(�R��Ĥ�%���QA�o������2�� �@�\�#k%G��t��ԩ!�qC�8�iu℧[�+��\z����1�]Vn��� ���Nئ����s&�#�j:������e���PfF�&7"��q];A�`x)�
�7��s\f�R���y �6���iuӟ�����`��ƨ]A�:S~���@3��P��;�8���ᙡ.1&א�Smb�3ʇ�t��&��j�O�MU�Z:I�M~mw!F�.4s���\>�z��2�ʙ�l��6�Y�럝}���^�'�
$����^��9S��q[�fB-����遲5�,#%���ށ'�h~��	��
�j`��m,*�O����i���o��,T�Ca�x��~����vM�.�W�O�u~?�L�/����Hs��!���jI��f�v���� ��G&p�58������2��
(?�n�H(��z"F���+�fP�q/�7�$����#н�.��?!��[%Х���\)�zY.����#��qE������/�ޔ |���{� �J��G��,��u(�.+0]8���5����:�Fs�l�7ô�%�Xj-��Z2� �
�d:/���!C��A�h����N��Oe�\E�X������*������b�A�>S.��q5�I�r�.ǚ��b�T���C�����@����i�E3�����a�>������N����uGQ�UM��w��rl��Ήzz����q۞��yfǺ�*{(#�"Y�Pz���)�����[�C��'�*��2���h7�
�\Q��
���ah�{��.�@N-�RV�u��M���N�bo��+��L(l����nl�'2:7�;����s�-:#tº�A��N���' ˡ�_��e��

��������m_4V��Z�I��$Wߎ�%�T�3L������w�Lph~#A�l$jC`z���cq�a��x�e�e��~�ri��Ñd�.�h�y�ݳiS!����v�j�,uc�����Vr����1_�>��&�JхO �*'� 9���B�gJ�\#���?_�p9Ar��i�6F��KDD���U�z���(]wc�����a8˂a��$��&����*��(}�#d�2iH�?�]��a��O�$���������{A`H���2əto ~��ME�p���ss	�GڒTCb�ŗG��S��pձV�-P@�)��o.ص�+���f�JD�rS�9��;p�R����BF���Wht��)[�����1'f�y�#x�H`�Hz����)����;~L����÷μd����ߠ>�.��;؊Nz�$��Id�S��cұ�츈LP��୕헤�s`��-��|EFF�2Iߠ(�Ҵ�����&ۭ��܇B�����8�M)��Ô�j(񅟆01��R���R�J �+�S�������D;�D�eF����\�����{���/��fޯ<�77{ܿ�CA�P;g4�Y>�J��t�CP#.��Ys��� �9dmjf �����n�c _��|�6=TU!DX	]
��w,u(����]��6*���"�C`&z�u�ʌ���qܷ�O�i�I��������rMpfmv2&L@���I])��o���W"���;,�l6���gX��;x���h}w q?^�J�f�;=`VX��׊�p�0�b쩣�����3�C�-��c�j	�HFt�}u4�1�ۗCp��^oR.隽�����N����c����?�!��U~����r�A����RÂ�ƪo>EB,������:���Q�Пf�Xm�ˣ��~��M��B�Y|��yf[�0�"�\�@?|N[��.k��T�:�58�l����[ɻb�z��-�\g������&�r��$��j��j����($��d2���b�$�r��j��*t+�n����1�V�ϒgα�#�ٳ�EB�Q�Obm܀>/?���R�h�6<�&���f��Fc�#1G�\�&���U�,��_��g��P� H��"����J�uw#b2�i�[��Y��i��խ� B�\�% �������R�Q���쀢Y�l�"���w��� ��R()��d���l����l&��YV��1Q�O�1'����Q�D��Hl���~:��������PE�I�0 <�$ �Lh4�$j⻶-�V���<?I��?
����'a�;���	 ��_��my�!�d&��`&�|�JMH��:��C�v%Bl R,M��	�i������S�iM&O�&����Á���K��L������|���;�s$����V�e�Hh��K���k�f�5Ru��-D��3ga݇3)�V�����~e��.�i�������ٴ^����<E�xqW*a�>�OћF���\iY��|�sf4V!�:���0k�n�3gA�O��m�='��{]��U�Y�/b�vx8C��Ϧ���И[O~�u�����Zg�v�#�(G�V�QxgN������ԙqޛ;}p��'��{����>0���4��a~>�l�n��LO�**@!�FM%u��:�o��@��,X"��*�xR�(S쌀"��o�U���C��Z9�;���" �Tvu���H��>e�"&�{�OJn l�����nC��\jJ�#�V���˦�q3kJ�!8br��<����h�11���5E��?� ��@�^B;0	�Ce�݈I;b�Ѕ_I=|j� [E��ÅZ�,��PX ć�����ތ¦�L?��X����`Dݸ�3;j�C���?'(l��$D�8����?�.���~i$�V_^���?t,���']}s�1Ye�W��|��:N$�e�ц�C�SkI� ���<�(�{E;��4o�I"w�q�a�DD���6���Xhj}�c��x�ů�h5�������<�2����p�gp'3�l^�v)J�#Ů����t!q��8ɱ0sFT�r3̓�2>YSf��P\h�Wf���Ր(bG��jfA���2C�	R�ƶ��Բ0�	��T
l�GO׈�a�)ԏ��I���~f��@"l�AL&E��t?Ui�j��^��e��0��� �c<���j1�������-b�<�m�sCh"t��ڟ��bi�T�:Cx�̇Q���g����yP�$��"���sc%P;�4�)�O�n|J�����V�{��Ν��̉4h&�*��PS��AV���ϼǁZ�����e8f��,p�k�j�N���@;�����2e��ܘ����6tP>�6t��=��?�.~5~�+M`�Z@j���|a�C*��q�-����g�U=T�+�5��;=m� �=?���Gx�Y��@�BoF��K#q�D/tC��P�;	�[M: F���L]	q����cS �0�c�C�Nv����7+��6$˕}=��6hI�x����?0�2A��Q9�K���Ȍ:�>�ª���)g��rE4݈;���$]ᮏ��?��=s�5�����0�O�P�d��|mp�_�L>�^�����,DIc!����;W�G���J��ߓV�[�G�Vit}���E����b}y��9\K8Z���-u�}"�l<_�m��z�z&�r�Va���,�E#�6=�
��'�-��D�9�A7kӯ��b\`����W�)MS�A?!���T(9yyt������E��6[��Ax~F��b@Q���<B�5�8S���r"�G��|F���2�4�Ua����J�c=���7��f��K��;�KEF(Ok�G���w|�Ж�ƋEw��i*8�i�,��>�Cr�FݵZBO�O!�n}ҞJM�_3K�OBa�8{���_��uĨ]�2�@/�9Y�]��6��6v4�8_�Ƞ �i�4T .ȥ���ם�RI�H����<�V0�l�1ې[��0�E߃*���ǃ��x��iH��y���U�Ew�Mj1����E��R��	v� A����n9���#���;��~��������N+��;�S�q���Y�;P	��͙]���1�l��A����������?�&!	�6-B �.�*l5�c�K*3th��y��
��E/\�8է���c�,�.�$����'��p�J�%PTQ��_���F� r���.��/nT��}�.��/��]�ƢF�b�RH�f,�?�����y�l�@��Z���7�h��S����f��'f7�����	�͕}� �N�<;���ˊdG[C�ڊ�:����Mo���{���G]O06�k	ѓ����+�����kF�LW�1�2��۵�5�۟-�^	���q�2�ϭ�L��JFi%Kr�R�C�ɧ2�n���}!��&��I �/�z���Qt:8H���x[��ӡ=<����p���W���e��ad����S�Er����|�v<���3���`"��g���E>tY6j����L=�o��⡛y>�"nQ1�>'�Za}�G����C�Z��Eo8�� �q�B�{��X�C��7�Y�q�E���Z���٥�r�H;"r\+�~��̉��6
��+@(?��n,c�4�ݝ�+g�ME}����� $�eym�Cx�.X��ɶ��Ǻ�\�W�@C&*|B�Z��P�n5%�$�X���1�	��@7Á��M�F�1 �ަ^��Ê��.w���el����Um`�˴�l>��L�|付	NLmy���Խ�~�i�����?ޮ3�U�gm�&����h]@�8��`�|#�s�1[�Ɋ��\�4 +K�B��m%�����X���.?}������Se _/`�6� =*�U�8q���e��c�t�J�~��t��n��8��g?)甆�{�i���ᝆ@����6(w�1�A׹���?U�L���U!2*�(��1l4w�@Qe�1�rG"����qw�|����f)���ȝ�uP�p��ߖ1$� ���8�tݶ�s�n�N��$����J��Q��y^���D��C9� �*� ��L����h�';�隆��^��o�(���{h���%o�p`t�Li�67����\=�[�	��4�ÈT�6:9]<�m�I�N���ܥk��I0�/2w$S��-�7�CI�;�U�"��{p��%�i%�f�]$z�'N	�C�o�4���a�,s�_�-l�#�x���F��{P�w���W��11�"F�k�M�,��Y�V�?�l&���(��!���mET�B��ɧ1�Y�\�6���AQ���S�k�P����~���`l4�`���ICN�g|����O"�����}���^�Ik�����`X�Q�<e���͠W �ߓӅ?m�h�c�<�fJ�9�4�(rM�Kz�?0�i,pS���G����e���1�0�ח�F+�[�A�<�A�I2&�tyg��U�Hu$�o�ܰ8��
��X0}|f7���	p&���W8��?�U�0�&3Ҕb*�"��[�*G4T�4��Ά�:�D�����$PI����&�\��~�)�[��SÂ���у#S貺:����Ws���l"M�C�Ui�P%��Qc����x�I��Ap���M7��,�O`�C'��7$]Wa�;�@�6����7+k��=L_���ן�ls�#0�����?��ǂ�כFB��	�l��=�R�%F�xCF0�F�zY��m�3q��&�c4��V��z���� بt��j�4�`�в0��)B�C���ƨ�P��z*���x���<А��7�f�=i`48�;J�P��nX��j���{@��/l�W->{"�DI��'U���xY����Ã�k${��]i�B�V�Eg��[g��̇�x'q����ou�e�RmU,Sׯ5�U�;,O(E^�}�A((���,ftSwX?���Ge<�ws~��P�A�S40�$��0�)��T���P�G�}�
��>4��fpf ���ۢy�ց Ub8�%��ǀ�������)�簲�Q%�`��Y�'�c�q���šG>��Ǳ�,I��whq<Ԇ���N�������M��.*o��ٶ\:�x��8�V
�=�kb�h��p!��b�6&B�_B)~�@��;��4ZS4N�ة���L���VI:u;��"�U��E)�!�{٭7|�X�9�@��n��~UQ��pVU(=�WC)Xyz-�%w�r�β�ylaO�����9zN�B>&�����
K�F�s-����w�1}j�����Th�f\y�s�b"�	���*:)��fŪ�;�e*�-�G��J�x��8���OH�u���3����G�i`��L���hՆ���>����lF�ն�������+�~e�t�j;�B�D�i^u�O~FO�fdO��_;����4��Đ��+02S�����7�o��6Te���E��4���B��Jt=�	��s�/!w��~hʷ���������8B<�ƭ��0'l��Nr���Z��~@2>��6�y�6�	`�E$� @M�/��ʹ?�9�YW�ף@��x6�<l�*Y5�����f;�g�5?��5�ة�S��޿��{Q�����ԍZ�7��S#7^�e�h?g?�#�����j� j[&N�HXt8���I݋�s힚jUR!�R�j�%*_����= ��VR��0	>< ��.C�X���!S�
xG��i|��l�Oϼ�nȝ`��%@�߸�=�u�siu�p�H�>vu���噒�/��hՄ��'�a"Կ�Y��[�#�G�!�S�֊����+Z4�|�+թj�+i��E�÷�¥���2p����a�k��1�,K��p�;�� ���ӈo��\aǬCd�x9R�a��Bt�Kx��e����-N� _Y�ս�-�(վ��A���g�6��t�n��}QK�9l�����_��9Rč>�Jp�����`��R��H�~-�	��T���o��^d����T�V_�m��eS״s� C�E#�wE9���aQ�8W��(���9~-T5i���~;[F4��[��s���nؤ�@������2��bWy�+���vs�Z�}�����cCÆ/�H,�[��W�u��@iMh��<�7k�Z��l�^�M�3qn,J*��Q�Ű��
�6�_5��j�b�)+g-���0�J&)>�K�z�W���}o�m���w�Y��%'����Zrp���z��-�����B8ر�g���kn��L�Ҟ�]R:��{3�X8���r�8#���Σne|��)e��f�R��K��t��W�Ky�g���i�p���'�]�$���=QɄ�u��VҊ�R�;:j}���{[�4� %�Y 3�iz<B����v4�\^��
#���Y�� J>ʼY�+��7�H�0t�4J�>u�:_�"T@/��.�c���>si,�j�ކ��q���R�s��H��3"����:b7(���wv�qZ�A1�5��?
Q%
 [)z)���}�d8��Є�L|�g<��)<
�G� bɼ�����i��5��hW9�_>��u��է.���C����zdV�뮏3�^C��uq�Jz�AG�#oگ�µ>�~��i��Γ�0"l[	�y�4'Ũ��>6�J��K�U:.��a�F��w����{�QNH)i�
�*��4�*�� ;q
N^���(��E�7\�Ą�L�kV0ʹ�q_~?�y�@�O�,�ˇ����4��ڐII�Fc1t���h�T���:����P����2%ԛ�����UK�0�C
�������
��Hl��W1'��|m&�Nxx��O�>��_x�B���E�$���E*h�]��u���v`�ʦ�W 8�D i�xQe�g�M������,���t%q~�{�A���O��|N��\�Ի~�$f4�N�^���Vy��8&���K�Y�4����F4���	�S��J�������5���8�Q����	?�{���᚟�!g����?;v��dqN,���>�qC.9����?qZEųl�~Z���3p��2^}ߠ�P�MD4G3�MW�6�u`mQ���P��#�l��!�1�Ac�+��/����
�aǶ?\EňZ�b0� �8-6h_E_�o��k��)H
�|ʽ�?���e�FH�i�Y�^����u�GF�z��jFH޿&X�o�\���4�6���h�|~;mG!H��VX0)�-S�e�3߰�.s]:����q�.Ts�.
6��N�����3�C-�2��r��U@{���D�����T ���v��ۏ*�9_v�DmB�U,XIzѬ����B1Y�`VI�%:"�U��_�L|m����F'��lm���nl�������M՘����/8��
��t���H�i���S��ٟa��b�ڹu� ��`�d�,5`�*��d�:J|ެ�JDK��$�s�a�ܢ9	]g#���4��ܫG��g����Kl������v?=zs�rЗvQMÜe��k��Wk�Afg�d�r��/Z3����S)W�U�M����ɺɥ���}j�Z7놃O���8S��
�ptXe�K��Q��8�����3�^��8I�����)JkB�n����ye��	�ۅ.�,Cs�Ѝ���1뇁�	� F3Hl<��hs9���7�*�~*f�̈��B�#O�ԥ��E<��I2V���D�l��'g����v�\����R�V)��;2:�$�x�N)�(T���d'�p�%�#�4��v�$H�kRh�4�7��&5_F&� �NWsItKNԳ�]ц[:�����d�P\W����Zz��l��k��X����9G
�Ӣ(�0| �$�$�!ث�5g$��m)�g��!�]b\M;��<"�Wݣ��x��ʇQ?��#�Qz�`�ٟ0�	���Y��F��{�|n��N� $/bA�FR�h���Tm�z}��jaK|`��"���D�lQL	GLt͟8�v�n��`>?�Q36���B˻C�"nO��t$���sb�;]���(�l ��Ӕ��x=��Ȇ�6���j�� )��{(��XB��7����E�ľw�K��3QZi����+�o���W�@v�VK���F�A�ܯ��{P�5�ֲ�ЩK&U�c���g��!!J6�A�g\�yP�kv"�ʻ��M�@�� છ��N=��٭�V��f��E��5N�q�(''�D{}~uѥ�ьN��������G�&�6�Oؾv�;�[��&��ʓ����x�i�D�X9�N  �a��XHj4r_�p���sz��!7��`68�%���]|�U�>qw���>�P�߆(�/C�"���\[n�F�����2H���z��s 
��Vң�9�,�Y�"+yAU7�*0dqΌ$�^�N�o޹�a������֗V���TK�
YM��>�n7�$�sf�DT��q5� �X���8p����3�Y��N+=��aga��lʹ�n�~q ����40��U[I�j�����{��e�h��DF(�hp�ڮo i/j��
J�֞Q�,�@QTז%ڛ&6�ho�a��%ʏ(��)�t�4 e�tP����7�yy�q��Y�d�5��ڈ�Y.�	��L9 -I�����Ȩ�Hk� L����9u.�҉�yV����}K��loG�r��j���i��R53ę�P-�B��rDh��D\�@:����ɬD&�"�����Q�w�|���Ѽy�WI|X��V �� Q#��}ٓ�ZW�Y�z`����Z�Z��Fa>DSn���JX�m�s��G���`��脉�.H����=��b����ģ���DՓ��3Cd�R�vQ"{�+;-�"�q#��я�g��t��qjXЧm����E��'����WZ(���qa��aᷢ�d���aT�E�����^��m��A�Ѩ�XH� �L����|ѹ�l���ob���j� V�-Y �´�\�G�E�F�?(�;��x|�@ZH��IA8d�
vUу���}�X�A3E7}Cm���;��U*�D��q�u����n�k�����}al�.'o�>1�����{�G���I�$��eB���zp��~��?r͙3=���)�Ev�z���܀�F�*��h�Sx�k�;H?�[��*�
Cp�!1!���g�6��l�<w=X���cR_�+zr���y���v#WqN��W�s�3]�ÝCm��qe�k{���A�ye��V��w��h�|�
��ҝg���3x_�<�
�A�)1�ko�@�7������yY��)BlB�?-!���&�MB��� �T���2���&��F�H��_�Y��r�Q�����O��"*-=�7����^'�,�}�l��_͜���Y��M%�U���7�D.&w9�p�[�cP+9�043��
e_^و4����h����c���oj

�cƕ��_@T$��2ά�ݗ�|7�y�;9�=�H���Թ��[��$�**
�w4GI$�sÐ	Y=}]�ӈ��x2��7�{�v��N�ŗ�M#�b༤F��-i���7���%�<g=ڣ�:w���t?����;� e�^'�)�j�V��uR�Zb6��Ÿ���{{2�&:܌��4Ԅ��'��~�P�Lr�^��Y����l��uY5E0ցH��]��<����nl�9��.��MM���yh�.9&������9�<]�C��TH+���6gf�68�X��й��[��<a���'��[d��<����L��V:yT�N"o�l��y�ᑻcцv���v�6�u��E=�bW�����9>���t������hi��9n,�ܩ���P�F �M�
�v��>7��M������9�*Fr/��1��{@�0쭚���Ӯ�t�z�e��Fך:�S7H�ꨬ 5<N���n(��[m���_k�w=\wk���Į�2��f�4v�(KM<A���:�@ب��.�^lG�(ɸj��Vb �'�l.�6�_�`.v;��D����_粠w�O$ ��5�6pp�m���1�>7d_�T�]��ufc�(�G���Ozg��e��\(�;o�h�$SAs��V�� ���M�z�UOׯ#�����%�����U�wy���B���U&�ܰw����rnQAЂg�d�)TCA[���kx]�j$iM��or(��@���Û�G�Yy�`LM�f�b<6㽏ݓ3����o1���]���0�w�z~�s��p�?5��a�O"��ka.�Q�1�A� ��� i"�p��G��zL7D�PO"A����J��z!����g��@����W�|�Q7�lȱ��s��6�
N���q�\Td�*WHJ���j��0#�Nh�' =K�f���b z2X�9��ߎ�Ԛ�8r�CWI���u)Q���y�S�EJ�:��lp�>��}��\udP���7�`�c�8����C��h��_5I��m@va1�7�GV�Rn�u�:��G�����K�*2��yz�
+�H?n��'	� �lѧ��.��"J��AK�^��D�a��)8
�:~��￥ӆ�ҏc����ϰ�����\=��"��pQ�3��̝�'+p.E��+�����gm�g�݅�1�qx�	�C�5�j�y/��P�[)���y�wרB�P��Wb��*��*�P�<�hi�U���:�e���{_6X�{�$G�^N]$BoL'|�����h�zj��D�Cvuy���W�3&���B��(`��-;Cnq�o�<�P��Z�'k3�N�W�1q�2�N�T�^,~ѝ �mٕI���L oa.*�Cm�4T�8��2|�TD���P(� �@u[�M�}p~3�.i��sx�<����S�sW0QD�>�QqX��Gd�YAx$u������X��Z����$%%��@m\�`PMg����?V4�<��ʪ8�6+F��^�� �'0u��M4�(�����0|J�:�����Jw��H��T���0+a�y�O[� �&Kj�6����-D�����ѹL��3��Cj���j�^���I���2h��E�3f�z���й�o"�J	�i϶�����˸���������qF�]��L�̖��24.q)�!t�D��@�Z}u�D1��4�%S9��U�ңM�%���:�4X�z���1�#��HVwa9̝@�7�ț
-�a�}e()���8M����[ ��,8~ƛeEO��~+�d�{#�\Hg��L(��=�"j�Q3����f-���0>���av7���(#�?�� �KX^"���6+����NP�}we]�n�Dm��F�/�� �(�������Pr��p�����;�����<���"ز�yF��9U���(���"ʜX�i��Fj�n�����X_2���-���zN��N@��i�E�1�`_H4;&�1}t"��m�F��ݵ�g��%>���G�]�7���</m��Co����� �|�z
\)N�f>�L��̟[}������'Hqsݑ�!��C�Ex����yYhWЀ��Ow.�/	�]�q1�AfOY�S��I.�h(2�F�
��
�A?:>l�������������T�e�H���������T�_9tͷ��>q��Qo��m���7p(�v+/��@���~pI��,���,+����B�{�� �j%�L�h�k6A�nR����;��Ϟ�4��Ln�0�]1��eU}��6�
��[`o0���8�.� C���T�Q�?9 |4�2+%Q�3L�[2�BU?иA5� pil�������[���[�8�$!�V��M���l����-�ߵ�P�'���O4(}����'��T�q�WD]�N�{�G����˯���=s/��la7ȡ!�`'(������J�P��z��r =�	Y2i�j�=t���N{#�4�.�,�p�����ָx i�Q1{y0���D����X5O�����Oׁ�E,���<�u����(��
������8н�h�I?"����]�ZӏXE#jҎ�w%V�oO�5n�+q�p�U��?�بK���F���	�-c}�vK��rT�L�ۨ��]ނ�H
A�:�n�L4�5��~�#Y�~�R�5�����qy��[*�����r�W��s��45d[�T4��i�sVR��6ִ�����U�o{!���mA�Dr�ɟ���g��7� �I��=�Vz�J:��?�q�����
��S����i�F�aW]�(�|r�0�č����Ϭoz��sd����5:���S�Ώ� ��i�)E�ɑ�%S�`v���_�.M��{81Tin������J\ί:<2��(�S!�:��p�A��wXḤI#&�3�C 
�"�
��J�!��h�83M�� F��U�x��`��u�׋&���jC��O9\���+��ɮ]�N0�V��q���1}�!���Nۉ7|ש���`��8��"���2C�Pn�[7��Qs�^�����+`�L3�T����?����rK��6@�>S(��"����HnH9�Ok��j� �:�v���
�0L�͆F@(���}��C8~Z��'VI@3M����	F��˓Àk���S�o�A�ЦZ�u���w@�.�s휕Y�LS�H����3��4AaP4����vg]�{0�P��:,B��,����Pr�Gma�ǩ�UR��\9�%��;�o��û�K�:m�-����'I�2�U)�nx�?�۷�'�G|�;ͨ�u��s�^0����7h��/%f]��HxV��i���h]l4�\ꠠ�g�VC�����O�=܄�X�7a���Z-L�A�<	Ά�#⚦H � �'+������1N�:�l�OM[���QۻG�T���|vpt�!R��l�a\:��o�3XF�9}��w'���? XIPh���a�f�V���Zb-�\L�j��qx[=n䢬�R�k�8P�}<ږP�Q�T��k����ɪ���,ֶf��;K��W%yꀥ?��T;�(%���O���t�H ��˺��cE���̛ ��ϖ�v k�'��<��tI��8�S��Ք��h������S;V�~��\R �2Mh�8~�Tu�KM�s*O����M�
��wF.s��kα���2�Ib���a鴄j���7�(�Y*`���u?�tw.l�7�~�c�r���T�*z�����>��<����#�:8|WO�`~��	T�I�=׹��8�������m>�k��rY����FՐq�T�ES*!7w)�������yӲ��8��|�����95F�C��#H4��d)�e^��?*r�b�9�O����b��xWY���`� �Q��o�w���6 T�?����(O9>$���L?*Q
}8�~ln�A)�c��>p�/	xr�v�G�" ��(مY���F'y��SQ��,o��aȲ������L����?�!�����7���/��9w��=)g{墋��7�O�#qZi��v���w��ny�w���ߢ�g��\����}\M�2^S����Z���/�"�z�0`C#�8���	������v�a�5�mg󾅢����e����Q��{3d:�y��=6�K�5�D�_,��o7�7.�I��+taG��f�F��8�D_;K�<����-�/]�%m8��lJ������
���!\�g�8W(���ͼ�gT�$���D*l����ZU�gN����!m��}��%Bs�q6iC����!�Ղ���飏$ywb�P,$�]���{2�P���c�/?���íz�$�ZV�L�3=�yd0B-Q�F�,(����L4�f���k�l�v�R{��]0S+��~�)����7Y�	/7���D�����H�/����+}�y��s=��@~.�9cn��6�ҭ��D��2�$�~h��/��tJ�À�L}߆�p�ۭS�l�<����IZJ"4,%��s͆G�CQ����'��#��8�-�9u���'�t.��e��6]A���N%*)��)á�*��jZ�/HJ^l|��+��_%^��^Â' ��.��Se����==]a����,W%a->ӧ��*ȭ�4��n�ژ���I>U��b�Y��x��8��|�OuOn���
]�A�C="���)sMq��)��)yl��ĮHo�|���Am|稩=+Y}�c%6��q��t{�&2Sﻨ�K�w���cp�~��h�����d��$l<�Y���/iF�:�	��͢)B4ǆuc5}!	D�⊹��M����CF8W�WS�`뜎p��"�#:W&n,�-8۫6����bl,Zy���/w]�x�}˱��ՆY|��7'�,��	w��4]\�3��P���a���,抛�^��O��f���5*8 -}8V^�"�*p�I�/�5autΑ�t����S�4J�c��0�D�����G،P�0�i7��k��i�,Ym�����k�WҬ�¶3_�_xz�*%E�l����r�@�����gw�M26��:Gj�ө)�b]�`�y�tӎ���'�˃�b�2uD:�
�� 4#-�JTV�I!ø�*K����q$ov�n��2�KsFf�j�J�1�� �캗J�Ă��S`c���8j�_1e����V�M�����q�_)�6�40i��7��P$,U*��S�6
$�VV4���͠����G%������,x�B����e����t_�Mhx?��N{���[R��
0�Xy�����7�{M�ՠ�	����z�p�?2D�,�+�JfD��<�n�ϙ��*#��_�����\)�8�i�~W"�9G�lQ�5A`N}[	�~�xމ�h��r���-!g6��ZhV �?cM5k�ac����g��Z�r���=��&n�@E���?�p�p\K�ʲ�̓rO�[y�ut�Q��:i�5ib�q1�&�듓#�o�Ux�T�Ϋ�²�\-f�,g��_,��K[���cj"t�)��jTV�� Y���H:��e�&\�����l鶆��0���~6��`��4�X���mjJ��q���^tZߏV\�b��!K���������{��k��� +�&��.R�3IJn����P$u�F�,�6e����Ռ����4t���P�v��-_f7s2W[U��� ��ѻ��?S�;�a ��<���W}A}�Q�Ϧ��P���<f���RGz�WW.��cT��JA�B�1
<��e�����s/:ݍb�>���z�#�&E>X/�\�xC��n�$Z�Q�����R�~}�Z�P��K�j�o�JuL�*7"�(��k�/��)R�B�$ࡨ^�ë����3�Q�w�a�h����3	���q���.��~�r���"O!E���V��=w@
/���v�ԇ���`��{�m�@��9aIË �����&f�~-Q�[4�ϗ�tYΎ̮�������P[\E4|�u�� M�e�2�i��D��Ѐ5
޻E`����g�-��}��L`i��XJ���g�2a����@$��.�P��	��'4qq���UȜ�{s��We���Q����Y�=�c���X �W��ZZ�b��gv�.Y���.*�f�hv�mO�P�~�n�҉)��}+8�SU�%�IV	����۬%�J�Q��^����}��DB��_��lm�by�z�2�}M/��!X/�JZ�`(nK����y��x��^o�!�3PCZ�9n?32�c�����=�%ؤ����_w*)3��sG�pX�4�6F��+",;oK�IyU�~j^���-QH!�����x*���jӞ�Nȍ�J��-����A.eo��;#'!������Ȇ|(��&�ض	�9�6�h�N�M�}
���T	E��M_�-�tDB� n���4MA*\P�Sc��/��Λ�RtIV1�d,�����sFU3W#��ODU1Y*����zC��3�a�����]�p�>EYy�%'��{���/tuâ�fѓ��	�`e����}�?��`�����ɯ2t�Z�b�]�mz�%�ADHH��oe]����ufKg=�ݷ���?�A���!�K�:�oQ��P|�J���6֘`hݏhM����`o�a�kH?���f�V�ܡ�Z֒��P�<Zl�9�W�@Q��w���>��%n��w�b�8�C��͒���}Y���aA0��둊�"eqs�-�߹T������A�\k4�1��(0:2�ۡ>����M���D]@b+�C�OC�:Q�c�n�ڷ��!�ηJ�M`qǩ��5�Ƈ7]����ﳑѲ�׌T�tE�=Pw̳1�Wa\y�:(��
r�<D��:�R:��W�m!���~�ȡ��fn�I�\΅hԝM��W��:$[*��)d�.�W��q\мx|F�o�l`;�&,��r���A�[�ߑ����в�{F#y.�%����v��$]��	|Xӣmg�~���2�Y�|VF�p'����E�$IMڍ'E�*k��]|}���gj�Z���=0����ĴjK{^�/��N�ra�M�Z�����t�K7B���A�=6�׆�����n&�Έ����`)��R|	B��m=�ᝯ��Wk���7���=i�(���[̅N�sf
.� ��롅|�Ҿ��n�����Q������0�u'uZ0et�XmĿDZ�sk'|�HŨ� ]��ˋ�aL0znܺ���H#O�tN�&��L"�By�}����kL�'�b�P��͡��\�(�ج=@��l��`����)�S�tMΆ6��IAk4੗�W�K[��#�D�R3��ig�קL���$��<8���D]8�T0e[�a j���C)�ho/\C-}��ht�[8$ J+�kD�`�>5s�����z��Z�AhHV�W��zD��o
l����2fI� ��1����XS�R1��S�=Y`��:�h|V�WuʻY��N��g�&,�Q59_E(4�s�.�m=���`�����<w�bG�e@�<!��`a���[u��v��JV�ˤ�z�J�E�R��jʑ�T� � `��4�f��a�4^%c�u���t�%O�sB�ԕ
h���?8�[p_�ɟ��	�ބv�;`�?[!&�md���
����;e���@&S����
��BdP��8N2d�`Q �O�,KiT��d�P�J5���y�k`_�