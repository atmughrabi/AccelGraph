// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:36 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ywz+3iKyk9dvzwqEzpGss9O57WgCZ3zq51eOPetPNgl/KmRn9UjrkStk7BEO4hTM
2b3wCNd12R0SJYZ0MLP7Tl39YVBxmlPDhXq/pzU8ek33bmfmyBxKUNOkwpjdk6VN
w1oAAx0Bof/1aI5roP3U3rek5u5XSP44XgiePkOUhmA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21968)
fZ7CVkyypjSjF316oOjUeLFqTzjiY28V6kgSWC7/tf2dsMUH9q5JtVXc/I5AFozT
/6dTdTiTNfTP5XCDmbB1oSlkk/GtN7I5AoljWkWrv1zweLPA0dB3GBQN/kKBy4WX
H53PXXsuwG+dIqB550L/aNkEwG1vogYulxaywhu8K1KGrXVu4bU29lof4R7IqiIw
C0AA13h6AwTz/BuIFWKV+151DikY9q0XcRli2AdQYpyjWVPQRA1JLB2Jc+0FFjIh
5Bgw0MbTkSQ0tR+KKmz56+skYyJBIsgFVKmF/doIpi2NYCUxfNf1VKmP3P7ltRNk
p3n9jvXlAYvr8Cyz5Kkx+c20iaX+8ftVy6AdD3q3LYSj4KKdm+ILuH8N+Isswc4s
yNIXCkTrptZlHegx415kok3ZnuF8bNdTCA78lc32HS8qR15EE6xmSKVPJNIKgL53
JXXgR0ZwcTF8EuTNNXNIw6Ql6H+7z5Fn+uTvC5RGE1VZBNlspmIZ9Xz1v1CaHfJW
wI5WyiT1XTrvO9SnIloOrGcb4TEq1BxZ5Rbq00R8EUJXDppaSui+sqDmMlQes2hM
jPUxLybjZwAXTi/8AQ95UOKmWB3G5V+IYMLgf69VV+RKWCYS4EBKhJmJLNLcFygP
D/nQnUEjAmdJEQZdtNOTTDzTltYHL4Li9UPrnsWVc5j7Tff2FAFpETl2vb3NNmz0
i4DP2/fi84/0VkIWF5/cIgymU57BfDNCv25euPtwvo6I5X8GESeFhAj7uITtWLrZ
BWTmiciYRCtEjxE0yrMD6gauDCnIKGuzLvwpUsMM0p18Y88CgvI5MdOze/2yJ5NX
eOv41doErzV5CdQsMRsZTGFXkab6MN4/o96dySSqCLmSZtWGsjMQQP+bES147Zps
hH2I7vwxH/MjgzaVV+rB25+OauFEuoevaqlMH7/4W4Z5a1o0ar4zNGt/HMwDivbj
PAWhlDl/R2RJHjCv534RaKAx2BgZxPDaU37Cb1rA7c/Qxeisxf72zF07kGiqEhyu
frDjgbrdFYal8lI8QWc1qLXerCnHCBNHvmYxnf3skK8IZY2L6kwdvC4zN7HjP+Sz
HvwD0BeUyoXqG7uol4NXzAXtnCqMYmKSAwDH10J9OMmwxQi7FnLbW+ohr53BV3Vb
ywCW0DpsIbLrSet/NIq24r0OMDk/o65W88Zl/I+mj6tgZz2sWsLcB5HOM+OVsXBD
rt2PWrgiluXLp/KPE1RtEuRioPKn4No7xQ93mHh6JyqwPQt18Ve01Iy79xXxDGHr
xnHUxIcid36Jy5PtzPJZCp/Su8B0HCq5wuhZEjNcVD/MG+8bjKlzVJ7ONbcPiOfA
fp61kJCXhPBQEq34DvX6dbqQv3K4/wCILm3rSIYvwW57jJxP/hxF4Dd33O1G6SCu
6eDX280EirEtyz9mB4qsgLvmAgQa1JsfH2f13AqngJEPguwz+64qs6+VsvaynidC
UcTJWxd0hly//KfOdJ6jH8EDs1MacP/Y67BBvu77Bn075Dw6foVa1CdvAKX13FTp
Mi44pmgqU2H08lL6NMLt19cMhk3upJ0IMYDobBgrf98pOdRe6ncMZT93AVY+Fayz
NIbzXcmd/ctuMTv4/PmUsOD1RhGh3zvhO2fvZiqt2+6VihPMF6c5MjU5mgpd0a9u
ZJHgl4YbCCbfJmVibHsV2Cr+nAp7yzJRjy96JpBVHtLT16zrO61N8aA9z08RNsVg
gO8T5vji6VAKmRhBXeE4tWH+KWbbFgtFmc3/VstipLt/d2/Oq7H/1cS6AnS9pxcY
KrobyTNeFT8hrxfAQbOvaHSbFBcnH/UUOlbTiq/sjy5UcSv+kW5X6G050BXv5ELU
dTAiJbk5gXIw96kOBXNED9b1zG9BZaxbbDPPNEZ9TObrMyDqV5RrU6NIBqJ/u6IR
HIMJ2RBQUeltPise7VYk6Quj4qThGeGr55848R+YqofIL7VcHUCN2tl3+OSIqtdQ
nvat/HTI0G52BgzlmxO8panhIKIxJnVT+P8+WJRao0xggwDpizFxmvKaetCRVYXR
5DKwpeUE7dQYStiA5Cdm9CrduqZSa3mACfh8jE+2+ZOT/JwBtuLarrcETjyqTVSY
c+GwwOrE73gOzeEhW6rLwCJVfuCNC20jiSZtJRXNiRTURoowyHjEzW3OXVOKCfSr
aXR8u475CyfFXHOr4qicSInTiwP3EiR+Xh1hyMbW0AALsIDRs22+/NmyGfrBOTul
8HyoKH4M6virsFMvRf2DEQHr4pdYi+QugKX6/2XGJ5h1XqEjI+D8UrvMzMz3Rw3W
jV90L99jiTmjJmD5qL+5UEJZiwpaPRubqZJ0Ege6uX9gK2AjKWAkWQSUvYWoFFoP
5ocquLXqmV3KZUbBeLon6dAu7FQNg4UkVXDWqaZkebT8H9DykMgGXXGmJJNNB/hu
DxX/XzAwNNuo/gcyvi9+YRRYSQJ6zAQacLCo20oI6YFTJTYplWnWSXyI+MbCBhKq
3SzR6rBwtQEXKxNCkrE9kdHkI4Xqbc/3sNB9qZcvExFLHLm7yHmOdHvQc5LDd44Q
mDx8Z1DEe127dJtK3BsxZvoMe8rkDpJW5CWhOe4QFZuVrC5T2oAwl5RrFEfKC/eM
Ktt8fPSi4Vy/+1GXedTg2+0pTR51nduqhdbfB42ZaAezjsBo2ri5XZ3SP+LdCZhK
HkroLKO1yZqtV4QFi/Rn1utITzyHIQNnyJzBYs1j21+yrvSIXXF/96i4VN0ycJqL
8xYTTUfJ2xqalq1U9pG2E+lcLzK+/nNdvHTGlRHqXf+m2rIEeZM+0AIfgeS8+27f
/4KaBTpEXVGc+ept8J3apl6VA8lPaItt0CNye4UWmOwOO8+Q/79X2VduiEKmPc0g
JNPSIllITu8u5QpVJYecx1JmkVVFKftfVO0oLGTrFFl6Ar1gFkK/jXNE98X2d/3K
05NiL8uJbx68ylB0MNylAsA04UpNchOlDbEMODyHbSN/SiEaIjRPYUGvt1rFAOGj
tsG+7Mq3FeLm2s1F61cx9Ef5d5RMUuEScF4si9tvGMH046kmJRuzTnHoSFz4gCJV
Iw1i4Da+OlX6TwiHN4fJvnGUodqkjdOoHy9voQzhdksAKlkjtHDhFO8TDX7M3SFs
UKrOTbtcj1ZL3vRJUcW0kuJ1mNgrIUsoeJKqboR7FawhSJAyjgCVefANg5hkjVZ2
7mOiJNQ0/DXKNrWqSttnzbWK2eKlpXSjnVUQ9miNLVj0FLuU9r81At3ar4/vtuQX
xby8hyto85riRWxWJHRMWvJ4D31snbwGAWbnFY5J2jwds9PRuIK0wQtTrPAFcKLb
RIhnjZq9Y8tToe5zmDTTykJa+ddQOfsLwBwpIoWipBcnUIW8UH7T7r9SLzJyNDzv
mdW2Qs3AexuAxhCmHfYhFehJFHKVHGFYUCNSFiyy5ZJq3HJ5X6lsCkD53BZ7AEAg
we7juKrgxoXKhs0xq6iZtM4yPYFeViIJyK2nzLqGVSH3pAHVZJmwjbC2tD4CTumM
E4c3bhaJskle5NxHkwaC1r3IWDDgZEYsh5PyQtrqzXJREI5Lj3kby6bz/TrMVAmD
fyKVDHAKcyZgcWcyCFge+h+1xjBaVTaj+H6pr/bvkuc0wlUjZWVlh/6LQZwXunGX
XJVQD23Z08SDRAuvw73AutLUqRBhyPa/k7TPXbRhonaIm/ibnoZY9A+7dw6/krL3
3KewzTdHN101F3VzSKaolCkFpCLRPMzvdFjGijZ3Yb01t4q4FgTy9O/Hae9I9vsm
wrd25vyHlSa665c6oxekBKgfcTJ1rKgHOmH7EGYoYUxOO7p/u7wItowDhssMGwH7
RjxOB2GNXE8LE4Z+9CwBXMDt0UiB3zueJurTYuQnP/j9Y6XIHXOeOdL7LLRG6bJK
H3fGyrtddEjVLxTwhkhYbPtdyZTySh5n5sfJz2A4ZfQ8FXBRRCI4nQgeGtVwOD44
ThOCZBJwHLbRRlsZpUzPOZk8Gu56bUAywehzn37iALKbHa9ZBrWPOkvCjQUB0olL
Kjb3ubkhYaJGkerELoADddd2rZ6VyktfyFzSEOC/flldH0iBJDpi1UK7QP6UOj00
pqtoPnmMYqS8quTmAJIc7+frfN02thApzKj7MqLDuDxVCHE+9utkb4hs4AWBJrSF
bPfuvkXrsTpih9ZaSTmj3UZlkx8NcCYBS+zlZvfCoUQp9B4Y4XfFxb3Q2hJDh4nS
QFS99bHTAZ5Wre0LBxqVESEFwN4XoiIqllCuzs9/hy2DuoZ+lBsXN9s9v+OKdj7K
XjvBq6SQEgMn0QGlsL5sM9B9CVe57oJOGCofllUbMocp/T7rNo0UZU35Rdgcri2b
SeJBf2eiADcmbhXsQpwsrSdzgCbGR1+SDGq7Pshl+L8qm4grYRjHhipq+sjxwbgU
ct86GyEx2jYKg2FQjhUsPfSSO1kwxtkEbJbBK19W5hjRc9gXDAF/bAaIFJN5Kw4E
L+zh4ReMVn4QpNwAPEtJOQCddqLWgx5hcm34Or9JrToypt12N23SVq+JDg8yimQY
B4coew08u8MhtDrkkPpOuOhBLlJGiaTjxLh9gpSgiKfpBZNhw7gCYyKGkOUNEmKF
f+YHYLcJtS2d4PQsWJ0fQYfK20kBr715B+NE16csKziA+Y4j8thvkx9+5v2pboNQ
7IxrtQY1jwgvYU68mXTmROe+8I1SPclJhwYfu/mimQqVcMtNMJscPU1Btcd845S0
EMXC6daKUm1/lzb71POTWyoiNjrxci9ZPl8mkGIarSW00G6txvSkMLkykwGAhQfD
+wAARd3+5uAXDC3Nr/D+zsfraIPjmON+lG0BaL0FwL4EAGTX5AtJ8cQJK7TJnAGd
nC5BI/Idj+F8wktt2CM31a1FTptEFM6HpkKmX6gf8WWcVB2+2BduKcrryMiX8E48
qzWk0UzcwGblDkMdLsk90y6AFS7nxhnESNv6y21yZ8EXC7BPBGNo6vTVaUw6RxOm
fADp/PXVhfhl+zKt710eEFtNYKO/MzjG7n5JOWzvGI5At1Y+qnWItiOoDF3Y4BMQ
rHJP3+VlQopZq+uck6kP5+YooXMQQLi59cZhxSZkrjLZEtPyi9URqjuiImE9B5Ky
gLv5nbBXgpqi0PhqP+Q2C19DgVA31xeCgIYIni5oJ2zgr9IBLJd+VR+ISkH4FhdV
H18QRUXzGwYsjnb6/l1SksYdB8nBZjojgFPU8eQuR3aVxlP0QI9yGMzSxTbUvEzk
zN/07WJJWYncm9jUdhTKK6/AQfkvh2VSvKbu4YoCXpFFEXPADuInH38XdC5+w3g2
uSfUvmG5p4RtcA8DXFEV3L8K+/jsfs3FKQykspdikwHl8bFVgStc37HXdi5gCAq9
Vz5DiZ3ScKxp2plK7bm0uorN0AJqMncGhoGUZEF7mNHGJ53IKGdIbWt4pnm56pSb
C0HpOi2dKcLreN0+sd6Iixr+dt7NR49BzUtY2Nnc8LTlYA4Ki6B+Eoqiya5MU540
pqNcsiedI73cLoDaTYpICKNajXlvANs9TK8/GgrCUVO4AhwLl7N8eiTE18itbiAa
cp1V3DGRCbDtzknUm7pcFJiaDQsm6GijB2mudQKBOZkVGfLfWABVEllF/jUrNeeJ
TLQSOV6xTXkhbrwdHrLlsnozJ0E5deSj3jjMoly/Q4ZfwGIEzWczW+tx/iWz1j9G
JKO2Iul1Jk/7JTnzXS4AMwX2Tb2394/q5zdJFivlrJUH5NRw10Buve+8Kk9XncfU
acMF95KYt1gvfAY6JL36MFZyV5xzZad1SLkRhW9gmjOPoIHNNlE3jrw+55aDRYhz
cN04YStcZv6Lz6HQMuPBy6/8xONWMyQ+xVa916YM8JLWfh9BDp63hSwU+DLgwnN6
0wUbZdAd33DgvfleaWhyKT5BtVkYpJYAra7Pdu8MXBCr+SM3vr2dkNzYICxFZh69
t/eKG21JwIHnmsTVxr6clwtPjgaVCYY9pq2BWaI7yI8xV1pIcBFJV9Z8dkPUfP1I
mw4Q5XWL1Hf77RkURtCAou5zKMwkdlAEtnxt5atztkqKPK0+FJ7Mqgglqm5c/2bg
jzUkWuCex+N/UEE/ZQP8G2Hmexc4NwscwtOp0ZEk1g9S4r4pA5wLlRWxLJTxV1iD
uxXukvwg5k97qSmw5qDq8/6iAiSt55gdBNw4SdAM4ZW+Y00DFqDcEcxU2uE5PL0k
rzozrO7cLUQ6wFvzG88lkuHWHtQw5GHO+lCXcNlCeQisbPyc0LttZMXfE2T4gaUd
zpugU7JAcdzj9vf1bIImsA/HIJGDXs5ghQVXwcYyAjwCICfWuNuL5tZjyUj4bFyV
IZ1nu1nrbUwt38bpKebVkPkgS7KvR/OrORm4NaSZPCkRF1B3ws8RQymZIT7tT0DS
deWMsyFV9h29H7H2Mvw56WMsjQ5ODqlQoIjfU6wh7o38jUm/2hOA1m2pJ9Y2Xry2
zBFsRvnK461Ivt290c6rYj+vEi9sCJoyVJdxbNCUU8+HD5xBkCtqC7A5iZx5rxbx
WMCxdR8xFG6S8MVGqf0nw7XJcuTIJyDHRMbMwK3G7zCELrIELu6Txf5yW9wqyfFd
y4c+TllRs5lPxJK3gQk6JcoTw/JqKXh7Rc3ksDjtzYEy5l6UBySsZcaLWwwGcMi/
UF1REFfw4iHVnFfe4rkbYZIK5aYr5aGfzOVE7HQ1gdbIZXP+YleTf1bgnS5SgQfS
uWw3WO5OwxUqMjGK/le4zDm8qdA3ajyV2zl1MAACOEqCF4QL6ARZM45by+LkbY51
cYQH6qAdZ5sfsIdQojsa3Zwt2/n/xwTxi/LrH+6t0Uh63A3qZ8+WLPbiMbE6/t2z
+AuytGg/D0845iEofsJbe1oB6s+eJgUcvdrgQsLn4AU7nCHp/fP2FLQjhwyhKtYH
iFCl3Que/+5yR4Faqj7egBCBYwmfxzP4dBH+3nDD+4uRMqJSwb1dAqjKctkQZ8H9
aeGahvomWt7G/picdJhw3kMu6LPztrM64XgCXw1buDbSxBhs7FpKYn7ZTyU2QXpI
voIXRlF9nEYhyuOqmhPlTY+vZVDIXiPp2k4FeNRNr1PNCjQC7c6AunKzDuXCPfDj
g66sQKIr60sy15kmRar9dDui6IUAVMW5GaxYpXwjRDubplrPGAXq31oiQigbI2tp
pTrARPJG8fQtna9pEgytOlz9tSIsNu0tXS279rpG2le86eYiiQEbuhLT92qnLsJ2
NBG02UeSVHKVKanRMbYbjLC6RVo5F7HgXmv0d4zyUYw8uhC7Qsh3xhR+uKeM/Aw0
mXs/+XsHIIvldDyhUNdiP76FoX0auagVVzlnLRhTETLt3ToFsQh7ctwO0WppQNlL
kifebh8O96mjfb1S3RP048m02ir5PBXxGYgDz3d4+yPrmME6/ybvcZwrcOuQyupW
C2OySFWEIV97ansrM5yrI/qfxYmz1xXypLy78mAGsCOxAMS3UNFZLMzbLd7yA1IZ
onk01VPPAjxnlQbBb/zbbD5Jst1Os8A3HeI1oQu2Py+37VOGVlRKucvgs1HEqZR0
anmKsw9lmwGpYgytr0H3UvkpjY4wNIMC0SNwWXjiFIzg0qPk+S49CiEA1g+zu0ZS
ytcSLEaD5JQTg4/AM8muNcvCSGxpVsrFM3Co/ueQw+8vGUV7ZijYCrluwb19MtKh
RGiyQuM8WX9/vmUG4lIDQACmNPjjVfwAsBk2N04SHcN/4Kh9/LiztKnb+5gOcEs5
Xn1d0xhpj08cE4Lsxaq1jV2kR51hncG0Cl8j+N2LxLfCaRiQnhOeMUDgfBho8v6d
0Tg/pHrir1YMJgilYcX8/LCzESqnciW4c1Qx33I0Kowk45AeeNL1cdb0PbA1TV/3
9OGPeUphRqHcr2SJaXIj2PXq4KF5pLv45looqn3+YiqhxiNaumZYqkBUtZyiZox0
kFAodkNNkO1A1F3O8yehCMTBOeb1maHipS8XXH1vgLXcFhP5qenqtEXLZCDN1TyZ
FGIZonAf+CZmN45RVKoBmpYQe2lXOpba2mA+JUU1UOgjeVHmeJzYGAgR8sSOqNPK
NoIisZJJP2P1WjAyWBhSyyeIsCh3NnvVUsqVDJ5/RLWlp/pjySTNwoT9ZfbMFSRq
vzjipD30VEJBjvUhhe5vWkplPOJQ1AjaIlEfX+/i2XqXdGxVXBrOBxjABufh3yr1
Mr0HmjwU66GR9n5EhL4qAJoW9HA0Md3kZ/vznjDSG1MY8JrFWCwKNgt74hhTeDSd
8nZ9tQEx8PYBq0jJzx6SYd37qQ0/dkH+5NvIASzY+KVJBe2XtKXJf1+8zYCPZVFB
7try+w8mNvThD9IX00CKvv5OM9SS2S7V/DjIZ+j362oA2H4KGzhzA91wcX3bVOoI
NpAyzHOcrcKicE4w+ZeEBCCzxemTw/u2TPVdEa/2VqV/HX47HOwXpLs4xphpcBhF
tlAzK8Rr2Mzg2OLHTX6aOJgAKnaxxxSFD0SbXAGUMj1S2hhs5FzPCcsBVjp7r/Lc
8FPsT1K2juAUT/sSB8HQoK+HSkbnloQq0iZ/yM1ZK8sF4Kc/3SVSJJKwOBw+GVFq
N9PVA3c423MdCJ77rYfY/YXKyNeIjYseEgboj1uQYjxwOj1qTyyeoIy9QQJMGYpz
oSX46tGFAK2KBP3dGnw9RqtAO2HaEDvOn2pXrgZJbURJwGE0ozvE1x3W3iixLD45
0iuPb4JKIIMeBl5NSHcHYZGmBb9dkUtnU1nO0KaQJKfo+/xgJ72E3zfbjEJvebox
H/OxSPoDUxMF2ZR4URTH3Pdz7/N48a6HEf4P/QaHef9d5N3qgZgNeEF4MnLfg0zQ
p0rD338/yIQ8lrtt+m7BRl+h3FHsAhszBVChRQdvJHzZz/YYu4stB5qcLiiJAEdW
YSuWMzuMz2vp61SI1tB9CmkPz1VNm741Blc2vRkync4//kGoexNDFHjXLYhymEi1
3igSQVBUBa70N14O61fjRZQHY3BSOv0UN7934+ACRZq+L1iIsUXwoKC7aU7SqNrO
5GN1cV93QtoTYzDHyfD4eA7+NFxIuh/8QbXs9kDjyXjTOl+9LqCX6HurxzcoSoCb
5izp8pJjfUZnIkEnsaLN7SA11adON0rLtndtgI+3fX5OEgGmp6yejD2XJ0um6kll
OnbH1Rz1KinVFszVzoe2x45PnWdTmbvRILeffUcWqn3Qk/bUQ4LQaF9xZU2E/bA8
iDVM5zVvzu31yuDcxMS9Mh0DF/7lMAW+fpNJ4tL/p0ODXscD3hRtgzMP0WzffPBq
HQPd2MjscMje8Wqc5xSqpPqN8P+YN2np9sMvEVcA/oegJfn3kYT0ZpIYS756r+Cz
DLL9iSIP87JaU5tgcKWT7eOJt+swBeSn6eXaH6fWAcIo8087Kn5HgvjWDn+7Rc3i
zg6n8MeK9ZshriSSTLCCMZZTSrFZcA/+K6HyjOoN/j+Rnt+u026NpaL2UsjHlfHi
6GT8mA65fIUgtBV0XOq3LX0qSKsI6HrOo60N02Vf381ADcvzRgf1yEBWwFin5F79
OlTuuY8eEzPG/Mq1SGj/u0ePJF7jM63ayqwDCh9kwacAv2dOUL+5HBb8LVIRNyWP
gLPJFCOPOnoc/ONqXMmqvVYjQi929Mddbd9oFNkvOfkjR+teMpnL3uOrlwVCJl3Q
DKAw5QbUEgUuiIyPAf33IEwD7BUZtQ4xIYHGMR9yWWZ+zCSyYnLCCHLu1erds5Xf
eWJU71BMIkJ/7Cy7AHJjS+hs7XCQ1Tidkcwt4xgAV/Ib+0xkw6idxRELIeEbrQTs
G1tAD6W2qIpLhE4dVZvBFqbRuGUsfPv5eNLhjBZTpFW6j+a4lwWnbOtwkjddlTs4
0X70fYE1LT/odCCcUuWbb1/2jACEvPkceluAVpQzDPbuZDroxbpS5rv/35CA36s/
T7w/brq6hno3PlNjGC2FwC0yZMWKy/JT6frAvAYQc9w2AkZ9d2NWYCXbk9DkqM8x
T6ptqOPH+oT9tCfWIzU9ik+CkTHxRgz7IOA2pZiwEvMJXYYX7QVLmPg7DDN67mQJ
71ARLSBxY0LMV5tDNkNnaXAJS6oux9FltK1u2lbPmAqAiJlvqGRd3SfL6oJDwkIQ
ptOJ8bCjBOY16g1tmMyrxuo5dI7avSpI7JDU9pDcCz1VK1K5XxKVZNs3PQrSFTnW
Br7Xi0smiBuPpmYPi1EslTeXalQ34tpLCzwTa6OWuXhlqd/EGOpDC+NNKuoqIVPQ
xSNNL8jA62zZC+FlrJMrBUbEEn54l/xtM5BAiDTEn8zfpio7bEaj8WTGFZjQ30nP
h6L73tFj9EaRcGSqeaHZMKPMvgbALvvBrNp6D/ByLZ/92HX9swoMa7JoIRWWXTlV
4eLT/ZFyj88imMaGw9MOVR43ETWClBInlEt9PtFOMYcfd8AMPfXXUYRQRlPU6nyx
Df+z3l7VTxQtWuslY2nDlT7yV+Q5oKJoZzRofHReNMClXgQntaPEGXUbOY1ASoc7
AkUu1iJOz5amJRkOLadHBKLzixElfGBYupiHFO6XCVBXRjvj0su8ieLiYtzoIQ/k
lK4DrzUTvpxeJNzkHCMz1dlRuQdTAUXMqUlD2CL4ncP++sb+dKIAI+m95xoLZiak
ThWGR7CENPdH1cTjszyw/XzV34BSIaxXn9gCOZRZpy16IETjLXpHqiRipzbvN72g
yGEBfuLjbmo4I35ClC+Bw0S9pV/exoKf4bt48AwTIZtjhUJUCzPYzn/USoguHttl
y/o2fR8noYBNzqu67lAGCy3hB28F528v583PLOHqiBHO6tie5UqaqS+aBezr5Y2y
e3EsZngnnmkls5D9pCwGC2ijnfcAKPMQO36CfjfGjv4ijTnyKaIA+jUgxyCOxk6c
A14C3w+SiS+h1pcXnL8iycs71Sfzby9yPQ4AFvl5/ohx75t3GVhd4LCuOC6+BMvh
NOF6hsII1UnKrACKUjEaaBoprmv58HkPRDIgPilnmZVj3fwYWyw+Bcavg2LhgOhu
tvNBjx/mBSYDzJ7rH2bnFeHFX9D9g9cxtfBAEhrbIBfZ92QY6FLCo7E1457X4JgW
Uhy9fxVwDkg6WzHf1ERysduFo+Wd36OQuRYwdifvQp6HV6uN8YSLs38obU1yhEQt
ue7PoLNgfK/vuIHN6BnLiU8B5VBXLCk44mGYkCgpQBLkfRiHdiyBNlc2yT8l3VKc
r9LwTof38MVrMtrowCaWZ3vGQyvQjopCf+hdSVgKMC0mZb47q7mmGxXHoxbBTdFo
LIIfVkyRhTIFMFNEY8uGKaCxuRueEVEBEpCE7GxSXBZi2b/hQpgjVqjqUBWTDKHs
uIQLZbTDECzFEzANEYOx1nH8G3EozNiaywpZGw09V2OCYurJIIOBa/oS1AkjeU8f
eWbJgqYFpDA/vhk/crB3R5Rc39ACAppDFHB6eQ+1JcR7HlLFXdXQ5Y+Jf/zoDCk/
I5/iqdHzTCIusvPKffH7iSdpLjPb6yDHFyqTGudIliCj2U6YM1FmxLPy+BXsp5bn
RfJ6ja4K/TAwrvkB4YBpbkaBZ9qZFN5bghxSda4MNflHiSp+zHx/ugp0Vl+4id6V
B8SPzim3/3j+lqZ+XjBNmY7ODIfpjYzyPBMAixh+e5Ry4YK4wU+spiPVOOiXqmcM
I33eBh7VTS4cDqC8HHTe9h/lIX4MQ2By+4Q2FW28liP/OUX+6fnFWnB8ivAK64E3
QilDBC77RFy0+Fmh/hS5caaAi2oBnCZOk01Hp9EAA/aq2Z3mn9wWsviFIdSxFoHk
Cjvod97uTRZocUzplnJwqwtmCs3TuPKrh8J0eUx3wFozDoS/OHBNmmo/Y3C0RMO9
zkETXxQXQB8on3C1dmN4nz5o0T2DrmLsho1g52W4HZV1gcKHJD32Ur0N+FVjBWSs
vbVzsR1O9/zEstb+7rrJf0LE/asYmy/hNpvbQF7iBq+gNY5/GK3vOw7xn52d/Oy5
i3MCkEs1EyhezVyNTQSCtI8UX7fJ3TwRx//neTv4f4gPZC04JBG8/quTMvqb2SxP
8OUCCPywQsEUW7k2Grx9KEJhK2OZBpGONPnOWc2K9nIcHYu4NXVKeY8mL8T0wsHZ
hCuizrTCxx6UkH4TucFJQ2jheBKWM/mN+bGNTqoVFMDcvMhD+4+/QPTYAh2V6HM8
fFeYKTbAfNaz5ghDnEAs283a9RKc+wCnyAW6+aZfI+sK3S0H/jyXw6c4F2jByA5Y
VkqrR2tMJApKc30K90HffS4iqsC+mLMFo/6vRRr02XnfCeiIt8uPwaagcYvAmWgr
BEJoiOHLR+ozbat2627fO5G5tQouYKJ2gonVrqEwmtHofkoQ6ztQrRX09AgIjIsS
+zcyEzDcNOLlh2MLeAU8ph6jEH+fRkoRRVDFVtgbJkDx151uDZtfbmRrBNVy6HgD
BG6N55u6UwryXZ6fgVwB64ob7+aEyhy5m+gQBY3H0fioKsRWRlJwunogtmxIAVF+
27yfwqC3vzWvW0k+dJqvPovaaXJrAegWmideRMevFmT9zSMhdOCvXKO6hkT09STZ
4Z8XW4yAmQFnvdjyk2IPPKz0tWPZInf5vZtWBR5ghyoAn166qdiWqtUq9KhehKQJ
930ANZraTYqvzS0EvNAE+PUoo2cDW6olAWulZDZNwe4yAqlqSUNomYhTLKvyvG4w
967hlbFl5F03D3aBGSX6Ze5eqklRRy4HNLmYWNB9oUhW3TMjuYFmI3J6TjKEBaem
L28ROaQh3E1VN4xyQcXvYO1Pll56q2ShIWKvnNDd5b7BF1G80Y6GdHbVzOkuYT72
Ac0o4+SOIuWC3lhVoP1wkREemy4c71fb6nLpMNqvMuZRLpMjNRPoLH/0LHNdzuK7
atnIi2owj47LO5kjA4eS6g8G/7DfT4pCNORTk8K13TXw4RbG1MOTGi8eOsfca2iO
1Hw9zCusIl/yJvZnp2FL3wRRWF8r0z7/AxuyYD8g0EUcFoJxtgCNaQE+CNQdK6Vr
zfrZcnHboVqeJEjLikesp/P2RYfG3dIf3O2giidLH5TkMGpFyOUPKvoHsHqygl9Q
m/W9Vqb2YOfVdlYZaoznysEhe1UcjbLuvRgD6ElWJu2dooeYZUIto2DanaXXsswz
JtTrPzrMscJm33TvoI4qCeKX2sS6JgGCEOh/hoZhurXUWmebO8yyuRLJZmF3yTxs
xaRaQL6bgK1YRgffmCH5d/SNEKyu2J+ej5T2LFN5HSlRsX5qVClbQTDQsrXdG2nR
jxVTvpbBxoaZvlgLGihPZpyt98VReV4ML9GMy+JLPTArscONk3toQAfChyO+2BY5
wy6zsR40MMEwNc6ekujlZPjErjQ9HDayNTi/92HSgBa/cBntfEsnubRLpP0BEPM4
QjPiLq4QtEr3f6aINYkBUksrRpOKmOITnaZRxDsE3vJZpnf81wFLN/Fp2rP4Oo0v
aIy88iDYNybju/6VSe+oUj6A3OmsimtUfhnBteEejMyd71aBwCjvtGsLSIFyje8n
lT/awDI0jSDGbp7PwiymKT4w+UP8IW+Az3WYC5uNMBo7kvE5zKejPIuhw+eyNy3A
xiNedrngp9e+YNycZm6o77oX4rpx2P64Lgtrmno0ELTQbCVZGNY8v2JDIp5kgl89
UTQmhGfjDFaB7is2YDlIMGHU/XHu8mQdpDjXVo/H9w3TqGbFYLRVgXaAw6Vei/8Z
KiVRdFPBcm84GWrAi11TvnBW4hEzBKBoQLq8Ka1y2HwqivAz8JNT6OSym4mDjP2s
SRBu40tu9FyR6xu6pJN0UXZMbZGwenr8o5U+O97P3UBlXdGXBeh5RwT7rFHIhqGI
z5Ecj2Fm147+knZOYoy98IRacTd1hA/8APgtNjdPkPAB9Cuxch7NwRjhZw8oidb0
W48K+yBqrEizHiLAP2Db7gK21slYM6YeXHz8QjhoRwOi6EN8DBL2Fh46nm+5NKRr
GD9Q52aWQH8uFl0DbecBg/yrjirK0Q8CygziF/Gd1OZSjb40Q2B8ycNvnzKcsF+2
ovbg9CJv6fr+E7lYBmKGtlwITaNtVxj94AqHu2lcx4yaVqh1IQMUbHJkAyy4/VQ2
5JxPq3RrxgoHx7if1D/NxkaAT6lOwLnmR/oXHUb6n4duzp5P6yT4m7tTCBl7o0Sr
P78tUThK1HKLbCvz2EIDJqFsFnJwaY/YZ+m2ieronVh+kVjPq2WlnMvj6CD4bAcb
53iwEK0eV5EpM1MKy7e7QsMeNxmyw7JQL1vfvQPwnl9Tp0NT0585t0bOADNtin1w
o2CA/SZrZqhkCIE+mwUZ9iG81iQPMfjMOuUvstGdJUWKJvHsOurgZ6IolAFCuVJr
xJXjMExcurMt0BxofeTNOzMqQ7KyyThc21gE1g7X1uIZpTMSo8J+qIGZLFCB/4XU
zGAeI9u1Ja3eXTfdwEOCP/WuX8ZYrKsaAmfNKBwbWexjI1WwilMvbJj+Y7QDkQMr
PwcHTpefyt0hWTa9HvgUnmwPvZ9pcgbD+s8QzuQfxqI0MzIPu6AHNr4rGML2FZrf
TWSoSGmAa+WAUbJ0XQKazlo5ESU6KmpfLS/uYIl4bhUo332tFB+brVyiFr9XB1dS
urQx7JLl70jffL6AxU7Mbr5opboENldw8nbL+a0qcw7R8AXGq+kd2cMFgAvQqDKY
IGpQS84dQYtEqibohjTGDMG+wIfdoa+nJWf4FZB4HX4izZlLz2cmhrMyPiIDhUEb
d8cK57l6XZm+0Le1Mngy5NiLBZY65wmCwec4G36tx1DBiDIa5Qh1bCbKsHTfggTo
2dUOfSxtnABggs3nhDxPFnLkEMUuxqvGJPvJr4ajPpUh86l3gVIWUpCd8+fgC/YQ
RIDk6zVqjw8jq1/KyxuJpVgWhXH9JY03zIwFlLTFSsSu9LqdOvhNc99Kqslb16yq
OmDjbr3H77BBYp7+PMYO2Q8VvuxQcoF75NZIvS+M8IyvfX82vfnM3EMqH7dIY/ha
OIg06medGS3zgg45mKyL1CL5aiKPwD6YBIOqtlAOE8kzwivqLYO69UfWPNXYV2qC
O4f9CkidEYJLq4BP0GgbA5UEGMRsU5L5rxWrG2zuOJ1WD0cKOMXMeSujdwdxGLoV
AS3tihzUB0Ry9Prxewcmm64HKrSM4UFuE1AyWnFNqHVRhkT/ouJoo39QJ0p5K/Ig
nXQ4xMVZi9VFYe5Qi+NPzBQIjxiSe7ju3totB5cEX3Xn+BqyB4Zqgh2U4xcVfQn0
SZMbUcSdktljUeULTDsHRlbJTmCq6prl7yyUwf21lVCuWDRMWuX4vI3QUq2MICO2
0pspJoJ9tTnOd5f+TzWjVUXi9pl+a88TpqZOdxtxa7Bo90/i5483TcGcusEzzkYd
Gma7HFDtPv77apd5ZMRyD2RGmEr/r0GDm8aBxc+Asesn2Wjykd5njBCgTXqvWDc/
oKkhXUwY2IMwxz0s7eCR/SzIJu3RvFbPgeiwUV5GXFVAS+xpKSTJQnZJpliZ5h+r
AOQABzyDgnm8R4kwkY8ZT5orFROpjEBfDycJwWTigODq+yRpzBcsAqlLXNXscxg7
/a+BQ0eoi12J4ZmJB3ZlIqRsztL3ysrbLohJKT1dAv0/pIqtOiWinRam6vRaY8fy
mBynrX1JvlAfQtISwM/YpTUMubgOabRDKradJ2Ro1YnT8g8DL8szta6ZBdVlhWrX
KrTErlBXPeH+RHDRu5hWn3C9yv/wdszWITaXU4q2zBC+lWujdDCxUoMuZTYxlSmi
+ppUkdi9Ahpjnip62xesU2aMNKtmtj5xI3iUCxMjktL+w3ir57PfUEY2uPHkKsph
+382foz4rcyXLdsMTje8m1OPFWrkAwAZ0AzBcU2ReGXAlqtZHKKPJKMJUXnU6kIR
0RhQSHfFE+W5TFEvXOvU5sUNB8ZtpdxEuQIm4sOuzTbTZD4bQdcijC7uhwcVjNIm
nPrFq2+LeTc92BqdCo8LRAIFzh57SBUXEfeXwLx41fyQ8ojBUsHcc7BCgjaeZ3iC
qNDsYi5zVMX6ipO0wla07MMJZFjo4OzJ8RQbt/HqTXhzAfIRCgIgvCoH+n5p+9YW
Zuu5lrPMFU7SJOdieWXYuk0PjxCsIOt25rd73DIi2FX8o0X1310G/GIoj2J6O2Po
a/dmkOhv8Dk51LBqTdkxBxjzjmxQVy1QelKomOgFlXFPdhC55/MNVicSzD+mo58l
o2zjIYdd9JFPgCT6XHXScMptWm881+PLl+nimATL9vZsEJs6JmYsJaXvzsvMhLsG
GTvFjuWWL6EY8D0j0NheGaTE0XVlDS9gl7eny14rVcqFaP/xSkaQtmYtjXB8oNJX
yg9D82eAvNC4QDSViei3eHpovalu5RIRDBY/993N643dDeE+JzTIcehdxwvUXpzm
UDhW83qF7zW0Oz3ZMct9YbtnB3bIMg0WUbIu9IAIiDaRWLci0X6QT65ppP6l6eHi
7W2GXppkU3kNiaqOuaucE0jP2uIc3N+852sJ4DJUfH3JdQnCnIo7O6pwLbeMRCMe
hO1JcCbbDhxfXOlfx2PUHNnjkIUedS2HlolHFLwEvEPsLt2oXXjhsBKAi2q4Gq51
jwRXJXmsgNZjYSMajFiaew4eO8Kqya68V+Qe3CpjGdWrkxTsxqgp3Qkc6pVo1p8o
bnQIbRY9f8cnJ07XPv/6dWJdywQ4wOoQO+yodAUGfoMaXOcKey7SkMy5Y8qqyIiK
FBzXKBz9wBsCIw440DrVPK9seQsqv6osnyv00SzC11enZ/L6aiSQZHBgdV8mwAAw
+rHSkasul9pmEHbIXvhaE0WmZWqBHZDcQ4vp+VL7ne1fdGja1dkHXgpxkTFqT+LP
vQXXJuUgRNmvZfDNX83WBITkMsZ9hF4eAq1sXINROtqTruGJ/Nr/wS5w5Hu4FCkX
CLAHwAF3PNbYc8ojbixtmHfT9xFtrIZiSQYB5KawcAK7k7JnhYeYWAhpP5vv8z/d
mSq8veGx4QNyYvZrz0O9BzUdCqvu3DJHMUbGmHRynoixgHsrEySJGPw9UvscJm/A
AuZgUjq6u1rBIS70jijLtAwKSyrzV/FH33etgbi6q5BRre/pxytZaWu0khTDvckz
z7FSJjV+Z4/zr4TsqrAvcPix4hODboQ8JySff36nD+SdE1mwjfc4rYwkcbH7Rd8I
61PO/M6Tyx1opNFOtllBEnjZXyx1ArUYWELCrM2FkQ1AyeuAspq4bbnc+ojEUoCE
1dNO3lpPdottnoLwgEdgT6IOROyFocA3asIVLtYuwbJHJw4ya2vfSJjTRphqWKo6
JMw2Sg159Wx5QpoK79yJn7OlUM1eaCKnU52gdbIE1sYnAZfoDnEAbBrFRLEgUdGh
j7Hiknl/4SNTIADLR/axct0O4WN1PHcm8A9SzvWWSHKrC66F+OoDIpvZBlqvB0w0
1zz2uMJ9AZ8bO/hxByhXMTJRSE22m7m5KvB3AG47bdH3iFgd5l/xKo4799w7+iFo
2zPdD5STAiK2mboEXkWMOYiVRsiZ2O9qnqchj9LaM55C/u3y7BkKvllEjxJxlQqd
onIiSaylW9Tid6lwchw+BDb0UiTKv5WXteCy6X38ro4FRp6CS7zyeqjXO8lRWJ6F
mntg9rH3mcCt/XQHWeXspOBBLpqmEeqJLbqjT0Ecwos1LKD013ah7ZA3xRsO8L2x
uW2hSEx5UqhHWiDSWwAndkafhNctLaD51Y5IsHuobclnA79WIW06DqzkeYslL3R/
j0igzjM1GoY4APBTcqxDwIJa7kV3Qn97knKMEJGc+hBVhFcyszqDtqG2pV0srYCy
aoDC4uVjpgkwygzKoJUamNf7qfAig6WiW7t2nWgKs24cz4APiTtK77DJ8O+rrfsm
oLt/Y6ytW1etyGt/WXAQMlzLJ2OU/pM8foVEwTNTGxYtavMvlCc8UjzXlOjQqeNJ
MGbmUSr2kYo70GNDfp2g+HMq4RU1l1uUiG2NVQYLyMOr0pwpr7Piz0mMvUNv3lWZ
rlzxttYpR3ljb0calgbT4KFUb/PmySfHMlZwU/6D3AkoecuFEnfU02Lhw/p9LtLh
dEDRl+1pfMGSAGeJ70ZYgbmrDQedQjJId/SWKnUlKgq/moXEcbeXYl+r0MbZofA/
MWjHqBBMeBGNNfO9yut0jVHRDy5JOPmlE8jO3Cl2+X0BqXla0xXkYZtuKJ3XF5dF
fPauDRBPdT9lIkYSHvnfs+fvhtRuvfLaF2jjIBVmjLrZm53FYGGIJ48tJUyqVvo5
7qC0R7FrbCYnwTO8SGe9wKzZpdJ1qw/gb2qoRaOkgSMF66N6fkzcdEFSTc+3yht7
OARIazrtaEFTe1u8ydNPbq3jo/8JDTpYeibBoZE8BFrePjcZ7hdCbB67T1wsajt/
qqBROi3dIneFy417G1pMcaVjW8L4pVhml3JLvCBIu6Ze6FGNXWxwYfypFfICuOiB
xWuCbxiULkgE4hUTlEx5BT1p8U/bvzZslNAU/RkbY5AsCQ8O6+v+MItAFddP+637
f45FrtGzjCCcPl646+OOsruG4HELl9wOLY5QEl5uaxcHEZFq5N/QhopdH8fftOjw
GyVtA2cUY2Q/DwZNNY9+oZLDvfcmruxr5EA39eljmmULMYma/oANSvyqf8EjID/b
FaBKM0ymTj7bi0gPaLeRYsbHHqplbg6tfiK7uqBNojcK7UWYxOX7DWiJcGJAZcku
hZRE/ce9Z585Qr4GmS1o2VNay/OvqQO/Fg6OXMr+06q7mQ+8ndy3CxNEqYn5ja03
eWOYcRMDsv8y5eOO/sxAke5XbQhWScFoN3g40EhwZaZ3PpqhDiQt0FS0FjyIVmDm
YX1glWena6oCHpRXF2+w7VGqHAgoU2Pe9JwvpvA4ECu9SMZhyIGEJtnNQDve7Dox
HK5t2/PLgL0lYmQ4zhdPGPlu5mxnHHyFuQhlVHyKLa7EA7MBFp+iXJJ8AThgEHwQ
NkapMLc5uG7QFdCMRIFvYwa4nWmM2K2bVvDAPaXUkaw4DFHlh6BZp1ZyfZncXdeS
tktNhoXOQtpsjgGILhBpdvStXU+mcTFZUQX+pxTYA7zaJ/20ftVPmheLawcXEosY
/sJHyxnTiYD00znm0k7oNouQMKjE0vpeCM/6yXPiNUeTGZkZU1Wt7OL73twpwkoe
2h+JHE2NsjZNgDQKrWt7I/kt6SIHhdEgOqRcy0ZfdfDZsunfr53hncCvA46u9MaA
0UuDk3uyjNjnplbPQyphFZ1weHtpXm0EV02OQ8ZiIMkZ6rUG00Gz1x2C1tfIWXJ3
TYCRC+ewBcEkQaDwaNQTVTkWlif7/O0A+JzZKvnSZcA0DdTCsmwqmiIvZglbbyCW
CaNULYhs1UHIyf7Y1uxVp3rf3cvlp0BdmJK94GTo0vqtCZRxQGGAg47QwXhYdk7F
RLm6eADbNMbfP1YdX2YqyfL9tE9AxnhfbYKOVPd3Xtef5wo25ufDxa62nu2yTdfT
bDtaklU1ThgiXI6Q50svkkzXpITgerzucY7Ipq6S+Uzqydhp0TxBZnoUY+HdQ6pU
PawbjvXq76+gVfTI+1q2GpdUhYjCV60K9PWhImdhbWHs9VRK5EJ48mQfSla9Q/KG
l8FFGfK32VNJbQXRT+VIkz0NV7Zp4WVTe+8GFek3kx7/5sOXo7XYu9bD5N8CCy4v
1BKAVyhJqQvG+SaN35qIc8PUqvCHPj8QjDNH1NZCbxh1P5nyL+ppUU0/XfULiDVp
nDUaB1cdOzBm2cBFQnv7R+eySHrlxMECGTej83XJt2CD4WDW5ZN5/7qyB1iRBARX
6XQwL+1+Y8mpKv3SVsEJ0hC3Gm4FUq1nHxZ0pAmxOzSV0nSQgEp3A3sAVbVvVTvQ
pQIAHKbaINddrGOM8GDHKfoHMfhkArJMSjtAWr9KaXCPDZTbK4dvf77ka09bYK2m
WbZmlc+kMf35lQ8+vDkaNuUE2orGAIG3xm0y9xHzLy9K3q7Cr2goUJEuL3vh6eQ6
zKKTaPjLfaAjh7vpMpiqmKhFMjhjeELLhhQCVDTrbsTu9aFTa9eShxZ27c7L4ozN
Rz5hpVksrFyr3P+vD7XPaZe6oQvjodOMTJUfLukAy6c8kNDOmqtrEMEh7YOBxbC1
3V5ljLvRgrvaSMm0PxSw/JfFXa5TSyHW59nGwQVfK5e7IK8YJuoQymlTHx2aT7d0
UEsKcEjjJqKc/ldLYtCeSXcr2i34MmA+GYJtvnBat4lV7Kl4GgJcsIwUpj4aF5Nt
RA7MzO5WTT16gE+KBjX6NKLgu15tUmU+Ch+lDK9ZtYweJy5Y6H2THln6r/1NAQCQ
85q++PKA4k0j3qkpiJzEi67igFE4gHaLVchCbd5Xkrgg1m3F6LzwTFWI1uV985Sn
5f0uruc0r9LYUO/l7YHHlA6UywXnX8i5GbAER4pvU/rJUTrKMB/BJ5lef3YnBU5h
6SikIbUDHVu8m6raEd0Ssj4uiiIxmnh2Mj6UheiOvVKFbEO7xrsganb1YIVV1mUW
GbtsW9DbMTPoILTlXF1c3ZZfUvyKVrnifg99SWMCkd4JK77vprTOUobAqQRbCvIu
Sr6LeaJNfR4HAM1RY6VrypRDux2NsYt4KGeMWW8qZN1oiEm3tMeuu7tUDe+2nNru
m+j1WKqARsnsba/R4H39QWsKQdH2IJXqH/j6Hv59wbkO5+XUwljPyvgOHbrFh8vw
y45FkKL4ov0gdR1k3BjoYcBY3NtsVjLXjbMLjKEB9dafoN2WFQyajpKpGmDnS5JL
raxbL5G0CuwyBdReqdoullkdsD+MehjaBnbnrwz5PqTICSdO8Im4xsB27hiIxBdh
GT08kcEz458DzAG81t/x7H1HD7t10ziGhwwoxLTLn/DqgAgCwkbaN42d2eaYu1kR
a6dd8C7fjfi0ucE50JDfLp5CgOwdQsE79Uc+GbVdNSXzmUbJ2iZiB90eGapVQTXd
cqbP/h8Yz03qzvdJWdVvAZHIx99hTbHH4xBLtg5iFH+xDEa7puY4YR5iTpGZ1yiS
L1SIk7fVaTHEy58U03Tw548dRckYkB93LZUZZMbjIO1yq47creel4zF9qbkU2r1m
2BKkAWHG9Sx1EcYEjOe4XUeG6ueRbtfHD9AxSo+VD3kRxvrEOI2osTpTzexQdeuO
50bbyQnsX+3zBDiYjAIjRo5384PuFRjf6DQ9ULu6fdVMpFeGgv3vXhlzi9W19IiG
VMEyKmShqucwoU7+xG1jLSDbG5q1GzVjT36xg3ffwlnr7rou+TWcV0WuTmx2/Jt+
scnls5+Nzhzeb6zXGc5lefXu/0e3BD4y27MpLIQ/dnMWIzIckQb5pn83XdTIwJXi
dndcbroC+PL/5hrJmjYlk/zW0exCprUcmbAWWQHxrQgN72fJY/AwV250Nl50gY9u
VGHnJuBzJ8H1DnM9kgeQjmsfJYOzTlfg2w29T+1NNY526cvsrlFrR0k5PkXmJlOi
b+Q4hEe4v/rd+T3fYuMBgMFkZLjv9P1gn3QBuGw1UCoVW2O5B/MgLyiFt5szUTtx
X1AecfFq/248U8Ei1xyWyy9qGE9J7cMFk9euEtFFZXYt5TJutiWfnFz3CeelaWD0
8oLBD7i3uHeQR+VgzGhNfSP5gNQVa/Di/MP9BPQhbrPAK/fm8VBoaZMifyFqIJqT
h6CcsT15iMGFAM4whTN1HQXlcoeKrdTHId4AMT9+LVZbY3oFWj6Hpe/JgKqBqW4K
4cSlOH/sxciMkU5sE7O5D3FYLJ49VJy5XeeaZyTrFvY18K+1Zp9Bx6DhESDT538H
4AC26c5Pq52ZP2dumcC0nglNrq4qPWTMQ1UpyYcnBocftS7GvXhWdHvU+2jVGVuy
YAxZug9Nqqjm4O5AvhLK7J0O43+cOTTBFLgW6vpChF0eWhG4mBPRRpbCoqPWkW8Q
Lfj2CyctySPikEaUQuhXLDS2I9PMBOKLUHxfwbBbVHn1D0G2p7qRPCPsrfoTw80B
TfW0AF66OksDD2QIrcoqZ9TlAHO3+rKeRtnlykzrI8ITmAO7TcGbjD1dEmbD5Swe
qpVAJsMqtEuZKP4/d+zdpDLI9SpF18Ab8X62UFOZWhjnaPJTceFpPLqpGAYCa1lx
wtvsKTTDNL3BWQVo4XGJNWsTw3UoYJ5TMuQ8V/Ip+Y4flbzQUG0LeazYJE7qj26r
oiHRUWO5Ywx45cv83Gg2H0Vx9MvKX2IKxrt8OGDkdK1g4O88T8u5qQy3bIlXnCQP
xYyIV2aSRUtvUbK3wfy9/NDLJDG3/36vRNpk6LOhw5P+XuSoVda0Itzak/WdYxyh
yyLGcFjeMwIJqIX6ZNPlp5KFiyvT9iQtOqqopRbMBX+Nty5zUCw+BiFA0P1AdIjU
0dL6wz2jvT7dPvtGxO/f5Nh9EItnTLQl37Hw3PnnF5Q3ZuBW4B/zsS9PLaghXfwT
pdJ3apCWTGkyXC5NxjvvNgxkqf9atF2cs8zHS2G5AEUMCHp+6y2DSYeonNGbmzf9
egerNTRlE4bLVeXpCILiaswGVFAp1Khoi3Hsp4e2Yq6QQHH5LL7t5eEB7pT918b3
aJR1kaIVXJqDx6wWGfuGAjzxHlat08/eJx7mPOUGWibUenowdwqHhmriCAYhM2ab
erqUX2drcFazid7SEl5i4KhSXSIrznbj27yK9JMkXaJByNe3C20PxxJxH9bOTOUf
OxJWWK+GOdBv9qSK0DOG0lFLRaCiV7FWNJvCGdJoR2tTSEQ8O93zEiDCM4TVt4TN
xK+6165is4QNiSBWNX5XQnvxVirmbjsIDohu6CM3QuRXGbNs+WOpiOmgQu/ysyK6
9sdPQ6i6W92JZyJeYqVSAtsm5Th4a92EHcNn8IxM3eW7d1jBY1KOPjpxjPaKuFVg
orecSdMjWrpwdwDoLJfB07gWPa6AQeut/RgyhnEhnQtZEYdrTh2ugLbjMBGR8YCH
Cm0eoemTIxHje3sB6oKFEYWx7Z978BVjwlfryNsXsbaOzYY6C/5t6o7k81OCxFf1
7CZSJCdON5Vi5JuIUNKS0yWWIdVpDjYws/91hBVA7aIH2tRmJpr2v33eR8ri1Q8m
E1SQsB5ROnDf42IKehBY2dv3JTZ8l4tt7dMJNDCQNMxooWKF9nnGWUY5rmeSm6RR
IRI7IdVfH+Jb+W+WJS8a/zcmzbHCEdTocLWrAdE2BcUEv/ZLX8nOWNTnpShwpMtl
99mZmjJuVFfTd6869GGYJL+2oUlQQiXpyu6WT6qbm2d71CUzfIR07npZOWpGoOCp
oqKVpLWJg9OaxlfGOLvrqjrJWjejOaP6gEXJlRfthxIGhNZTSY8B7Y7gYFjQaTE3
YIvstOvG46TJfALL6htV8mpmiyeEe+lA/QKUV86e5jZuRLLA/oovwgKELV2ZdHO9
AGteT9BAfqUi9HaheGxm6V02JLQTayv32J+oLbpySjKUxwuJffn0YB8qKWVQMcAu
prOvoGb8sRwMMTYXN6vkj2nYPVkijSKe54RlpPkp+f/38KiCERb991Br+UOBdPdU
LZz5fQiHsvKJJfvTjUvnsH5+Kowf2CZPni4Q9CYtwUbo4wQX0zry2zV6OQYhg0CE
kRe5rUHAs5zG5iiTqPsa61li3lwwTgcNuE3Hp9WGgFmcP7m2+OR5lWFr/Y54rOH+
s9O7FXDJVLj/phXTXx319jQTcan8aviowa8D3KS0VxJJmNSaPI17yECaxXIPNaIm
nUXSNcd4q47W/FnfJlDoxUR3MI43pI5b1wMudAQJcVKmZm3drqXnEuzsRJKrbuj6
hAIZgPHQkk08g+1O6YjP4kYaYVajv988HECKmynAQxgX/SmkbnOCgabBjTlm3DqB
nUCOw6uqNRIYNKGM/7dsG5XiH/HGy2dBOdUqDIT5TDU03CA96y4uK1w4TpJzqVNR
fUjjIYItKkzBm91NhPzgLc3VwpEICTGDBdJaIdeCSvzbnLIaMiWnbXr/2hruuecO
gNanLIg8pHL+pwtwihHgNprqOPGskK93RohVC/0sk8Sgcilfmfhs4oyWI9Dkewk7
l5hK2X12+YZm9Iq1LIsjH4J37JlypJ9FJykQ0MEsztGn8n4fxTmjPh+YDUrctoDX
Uk891iYI5ZCRiQ3sfGFch7YFDXcW5Biu6kUoWvyCESg0Iiw0D0JLay4rVtRSIKYk
plCQoDWMTPT0Giw8q8QB+TOUFyyrCbG/5Bu5N15LuR2l+sYRBOc/sKfmv7bVJ34q
zNqMvdpolHU8iFi15OZ9FNYDBW4J+BJO5ax0Vy005br/OetaLEsVXI0nev+FXdTq
qUxz2/g1Pe6OcG0BF6SakBEm3wLTZ3/SA/VsZ/AfbksXRaxrPqlW4YfMt/+VMgWI
NjBir+KsHqAkNwfEpwJsc+nLTecXbjMNl+e/fkuLus+HT0TW/chEP0sVI0YS0Gfb
4osV41kY+bqeBH7Zi47sI5PmajoTvBqrRZXtDlhRXJBKX57zqrXPCR09+utXv8PV
tyZ7HryWUT5IkVSL+4U0xhhhyQisw/U+CEYOE6ft2MjYTK2l9f0hqktBHkoEOslA
M/fGKFN0g/juSJACe3qzZiJl5UHyhwoYb8RouiSoaiqZvlm07M1czqhx4Bd8JWmF
3cnfqEAxhB6MJCte9fc0w8wjhl3nf8DtuLXwCb8xF9oEBwn4dDjKJPrvLNsDdeWb
q9Qc3PSZQ5GuNEUc5rfYiRC1Xid7bSnMTbpA/7pZzahPnDvg0ruWW9kgK7iB+BHz
ElEWwQw93nc48IqR2liI+ZErRt/hHXSoX6XPteAqtHVad5WA59q1XP3NRpLfnnEm
/+de/3MiGM1soaQ6weSGWH8KT/XOmKt0/WvibsreE/EhVs1whu8RW0NHqaS5AcTZ
RPshLY+phTUTkvqlBmJ9aqqwIuULeJzAbZs2jGlxDn9gk0CG9ehX2QxNIEJxBubp
2FMZip+R+scm1WpPF015JdcrSM+tE1ThjCZTOOL3mFOD35UCG0D30tMCKZOjbU+t
/5eRxL0z6JOdW0n9ZRAvcb0ZHY0g2SrGdjKS/vWgiZlszMctnYnxNSgA5mmcsw6e
h86z30jF1+Esnt5zHEIT2JK1Tc9X0tNins4jaTVHD4nBn61maaoT/C/rpCwSxpJD
pXl7DLTFqWQ4dR0VSnf3g1oCljo0Ia4Ve/fr9YET0nOV8qo07AY4UWgobS4Bbiwa
02OtPaZq8bwu0lWLDenvN2kqxM5P2+OtIQ3aklxYXJ68MEo39UJWqIS2V0oPBXfA
6XPdrYuqzQDFlOSBk7SaZly4cRvp89IO/aE9nvbTDc0zaZtIz4lAAqGMdBeUSN/V
EZGdRcWxQfSRftz/L6bTg92HBsCwGHT5VkXYT25i9A4bGeGya62A2gqYUNe3m1am
2HvZDkJinN2XIBE8Wszo0BgHYBYoaFUb3vbIDCnLQei2Bt2HgNyijqEEZxUm96IM
BTmO6SAveiumivV3kAgaQZPsnEPdP8QoHMS/0tLVjFeCUcQNrUPzxXyxwfWPwBz0
ww9UadZ2/Fu4+iivBiO3ytqvg+Q6BpaoBwlzsPPu27v8jAh9nKFDN3ExfVMhILbu
1QI2XXKYMuB5z3CeRX9AjGy9qZxxErUjP2FZuB//ShvF89laBKw+hx2GqRiif4Lp
qkdVBCKovplJU7WNb33sud0rXp8OUhdFVvq0i3/dU3pLDw5+BkiWEsszPlyNBKc/
9LTMyKAwHDA6N4Pm+W6Qly5bBaMzzZR4fI9UtkmWkSDfsTRwqSxlkvxoiW0n3Pyj
/r48IhT8nRm8FpOLlfvBmR6WdFnK6yiApwT/eefopE2rxwz2t4i0k6sRBeU2O2zI
3r8nk2h+worF5dKzPY4U7AB2IGUrAgZG9Tt+lu25foMVrVX0OatIGn7fwLNvk98d
Kx90WHD0kz+3/ot3IhWgGVzsxom4BgsEudodOwrG8Qd08JclixGi6ITAs3o9BSoZ
xFAxelkwiJTlHlJ8wALHWHE/c85KcP9KoAkQk4HfHxoBUkvXXKPO/3x7lhzFI75Z
EPJS0o1jzNzyy3XATBmJgIq3JUb6w0AOIWKZwTUgTNueWbHVUKnAc/XT0SpNUzKd
hkuVoLUmQZvAiTO7ibfBw9nRx5PSXAle/h4rPma9/zUBDPNQ7Ez2J5bRQDFXNmOV
kCGbAqW1+mb8tzwSvpYS3dGOI6+VixehcPhcHfasZECa2ultGnBEpsuNOdP72TQ7
PrUe4kR4MHMUVpbpQoZIjnTTYzrlAn3b8xscJVArTbFBTIm7xTeVRkimRNUs2mW5
ni9Q73Lozr3tZRfx0sI9i5S7dOCVyg4asuJOwa1nSgPIjnMOXD3Sn/gcrbCIAbIR
YE2raM15uHC7PSSs+/OdZ3D2ATFhrBT659/NY8lDgdRjIM9qiFhtlfzpD67B7vjp
P9XJRLAHsOv2+EVNF5GBAHr1mX26hQyJfog/hj2VBNiKp5W+jQWxNDkynyPl3zM/
RPVTcWInzQxPueEqtRMb3XROHwnnzhk+e8YhgcJVVwCrDT/yQf+gt9m55cbojPQa
LanXhp8ve3wVGq/xRDyEzeBFgA7R+HHcFAyqeD0ofyfxTiBwe8jhgVIVNUbLE8Hp
G+Z4wX2mBO7P7XeOrI9+IwQqJz+ddyArZxHmb97M4KPOPk6xMBCBU8tAd/a/km7v
ElRtUbV9Y8zOSYR3DpdFoK306sUlVMTfnJytiF+KZ+rzQ4C1kXItSnLkE4I6e19N
xdWowDjRjrSbumMNGOgrC9x9yqCxw+l0OxreUNOJ/iwA6YJsn6q5L8AKqIYUq77K
1UTGHQUnfyF8lxIKwf5A57LADvkjHAtqhwiaxjdB2I9yNPbEumYkGuJySGU7b6nz
e+12QO+iLiNMVOBqdXqUhr60rYsNTZ4wUJePMPPuu1k0MTk1brLsJgT6M+2+8WRr
VSNd860MI6gTzvv1OuZQKK9kKpSnAgH8NwgpY/OtwYmT9aktkr3hcQjB9kqqDQj0
GY9Ca8o8xs1SLQY4KGMaYREAvJCOTsmYbQIeByJcH90TX9MywPv88xUxzwAtkAoy
SATF/SDeSoSxwhofI+n+/ZUo140ciVf+3FC4M1mccU/FLGB8D00bpXt8vDnR7PQF
zzFu/ihvcuN+SR/Vlf7AwToufHT4RUcEimarfEcDAtdVkxb4Yihhytxd2gEL7mCB
QTI/UMTe3WoqmJ8gZx/Bzztmo1jxqj0tH1CRMSI5rZ4S5EtdE+lA+VwS2h4d1LPX
ew5s9hu7cSNnSExb4XNQ12wZ+9C7wUD75RsgjnOtFupOjbWRKdLa02RJhcw89dpj
KNRmowygxM4o8Q49bYD/8R5/amPS3N3RHO+Gs192K9Gr2TIUVjIWvJ5G5o46KM+O
4ApVGoF5eB5iXf2U7rptLKoQ/HIB5z/2ii4RKLipeAXn4LPr7vpV6iCfdtpgF1oh
qIjfg9Ngqcl8hQOqcx/pHGPbvNP9OXJyZcRS+KoblLDT1VieRuM9GyuORYoNVlvD
x8Box61JF2ESaGQlqmS2pyHmFaHFhtB/4wN6M5EdjI5bZbcRVhCQgf2C7ZuGvsPn
/vC34tmJpj793v9+FIytN7b6SVkXX1YVKMXCaHjUeQSdS+oMSxuDHWvOf6AywrqC
cXuQK4sUZ78NlKIlAl3rPW0JgBCyn0WbcRzbcrPitlQDvW0AdiddQD08XE0mS3sD
Lp4DKE7GxFVFDdqElNH7A9mp56iATCxbFEXwarpjaOTyRqYVJ/Y26S4sRzzkZU5V
fLCeVNGz3DCNsKDlgxqCTz8eI28jvF9aQtVNFd6SwS55vLQ+gwgZ0z75OXAQU+GW
ExnXYJ4HKtMQ+fk9XRQWj3raF5/H4XUCZr6V5iduy6H1tIwlYB3+ssw4DgxuR2PA
eJm3JC2vfdehmRCEwxvPnEterTqVyuDqdjEZgu3A7IkqGlebBYCj1VYhy0Wep/3v
qf4fpslHcHNbdVU46Tj5vboN949SvoZqTkcOyZC8YwHy0eVtQSQ8wNHKaJ9m6inv
L5SU5p49lzQz+1JaUUKkJVM1779O//BK4r+NuOJCaTuxNV6KyP+mL+MdbuItqSEK
1OfcVo4ivImoW7kTd42LK672Sy9Ptc8FMCyYZIHrCkCogo2Qq7Tq+JMif0mbAgWB
GZpPkthO386k5R4hnyQN/eo/Ie7u8sNBkkke5nvodMxOqb0pU02UsP9J/itdKzVv
KTqqusE2joJ/PHDckR9DEu6PWkQ9HkqHWX++9CvR1PGoiW8M6QpNRYgyikpe22kH
vcuR/e7ArHAABPzfkBq4gP3wu7hDfLD45XUZTsWEngc7QOZnnHedwKdpC8T43kKH
cyPtivqMspWD8BharBYopbvOsCFcZa/CQLvPuDmWSx0j7Fd5bLrMSxCP81HZbKVb
ueRdl9JXU0WjnX1hPcCsBp+rwlTqcf7HxLaH7F6aRuMihjmxx0loSQCpWo20gJ82
uWPTmoeIH4tp+TdBDW2O5m650Z+B8m9LKhtsIm5jfnQLpqaqClS6rdz8uj7H8/EE
LRGzObrOguu0Ymxtso2TVh5k/mTH39FIAvrytU4e09Ds6U+gJMq5pHxRmn5NstCy
IF+0C8AJx5BPdg9b069oTO4RnIRHKz96hTp4yFZ9hAn5kUPFpDmPiOKof8IAZS/Q
Ag/aSeF1LGnQCVhdOewD/FMM5yo9hqMxo6MJ2bzf+mc5EU31WaVsUhJBbRF/khY+
NEbiQkjX/NBzIRsIeWQQOOMSplf5s+YAaFHoIWwHP/LRcZwXCG0lKDFAICdUVbAs
Xhkkvm+JAImGOwDI91cPsB5boK8grHK0pYjj+MzOGBQndVsuXR7TkY9LA8okNkHb
ImiO7SoaawiiSRCH563pkaYoN6NW9CIJDs1Q1Ec9IqgXFzFlqKPtZx75bfvmD2Md
s2irYxKh/QhSdQ/Uxgzc7QEWK4sayOP6Ah54/mMXALRfJIFgQOdWmQqADL+SCCEw
Y7ecJLl3Dgqb86NYEfuuIIR60/kjrlifmTI79to1Ba5H6kKrPl7+qw7jVAT0NajS
f1+xOjBejsjf/kMueNG6FKeqfIGbjEdJjkMgAGGij8IyD5YWKFb1FSOagg9rMaBc
7DTlxm8D6VovIBxo33wCv463BgAUve1E0b6caPDHNK0QcqLzRrPJ4T0J4va+0W3R
AFwj2qJnIMvB3yVCRGtwlfzjfU1k86wluKo4ouS8ISTVSkllKn4TD7d4yoBr6HS2
yLNaDn76ydCVtqBaM6NI2V0VtCKkKlnGXI1+3iDcZEltuy7a0UH9JHUBJMQmmPJS
eaZfiDcubZjXbNMDk3h9TSyx7pB1m0fwBsbSPfdnGSg=
`pragma protect end_protected
