// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kAc4Iw+ClMXxC84p5xmMzEyenO8/nGBNdr3l+/ucpsz0m/Uhx1X6uqhi4nM7wjrQ
ubPqqzVbx3YYivPxLWzpEwMH1lN01qFi8o67k5gyut8Qb5vLxozQFTuzTfulfmfQ
my9NU+7D48mZkXKIuY19AgMsE6s0xh/BCV8lc1vD/gA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 178448)
bZzAYJ8W3JMrP6+rjQfcoqmftnZ038trHKpABg5Uy09kJnSDjsdH2EWTzJ1ZBb/L
+kpUX+0rpFmyM7N6Uny1/sOxB8OwJ6QbHvecF1AAuZ+hFHQ1Yomwidd5+hwvH2YT
lag0oGXbOdJrOm+tiVd1sVNiRDqRStDOKAgvscslzZ6takFUNlYZMDvRdfCUId0W
xJYRsAEnlBju1jqeNsxmN/z+vrMy51u3soVvTBBNC1cXp/dUmCBd2/lDTtyS6jNl
Q7AIRYJ8u1dgutECQw7OfEF7XLXkbt+IL5JljbXmSC6A8fiScfITekv1wuumDPpT
hjAQw9lakBuQ0EhBsLzRspv5PS2HL74nNRZumwbsqs1vAe9dGpY7DOTxj+ExcRv1
t2KpBwbiy5NSfpO5NKibHMDltsfhYhgPJfKzBBmpK/L17/Ht2j8hlUJSGKYHYZb+
VUyWOm4JDK5p21R00ADnSHqkYwYOeUCY1ciNvGjl2SdIDfHHRhXqp2TEl0QoumoY
IKto3XU4u6gI8fR1U/lx4tYFhBcd34/6hCNQIavPxuoGRTh5FArPQZnFZttBb0/F
tEgi8Tg80nVYCuKK3ZvCHLg3PeHgncuGGykt5bFQDkcKOO0zo58N/I0RyinU5jLM
F82qfZDCH3g9txCwIngFT1osUm+u6MfFC90uvjRFBnLiX1X/TJi2M5ygllc73M40
8ezalywwKDpfupHOVK6G+HW9xEg6uMjbhEO8R80bHCaPHBc4Ob7+uoRgD03mXiGp
hJkDPXsJFKnfDL8vdYaYRABFk7ktLuM8JawluOx6KmMgfy2jUlYAtQxLxIy+j1yU
beO+U622t4uz6f4Zg0mZmRBphr4XrOBhpXorJKLBbhZsyJVdK+V0TKBjmaKvtOJY
1FIZh+Np4mYW9ceX50G+hKsoFbi2ouasYRw8Ri2m9OmoYm1kM3eCzc4RxK2SoV0O
hmCce33VJAD4z82HHosQCopmiWUM9oEe9wzfMMxAnUGvT+w63BBiqmmhetzaNP2R
7VlJ10A+omHjLiHPRDgiJbtJ52yQbGcWRoXwlc9wde4cPRchIkc9fhsGhg2166lo
KViE0iKY5FXYFLhBB/BrWmHi75wXvv4O6sYSVdU3uFb1nAIeTfS5OPJc2VhlunDJ
qXDWh0eoGh5iPIG7yRU8br1qQOfIySQCtidHVz2+yQGeJMEmMTksj0fSZfBGEMB0
pVu2liQFcRhDSxSLeU8fgaQ8Vzu5G2u+2iaCTKprxv1BLk8vp/S4noZ6ZCLrDM5g
mvzG3wSFJAvaNhAjG7QJytQvjEDPnSoKxH3h53oYcYd9WY57HbwlmRdDFzFnv4Ca
pIN62vnQRl8MnjFplGyvgr0klll9r5km8U2Mv0VkY4o/6jX4om5RkScx5ZCD0GGD
YScX19sfVsPMNvquzRaH21wQX6LC5BOCJHWLyXhbM8x+sr91Ho76aKystSWGHerQ
m3jd3GIoqr5OCXmp8IwKI+TNguz/lqdP8quE+28BP0/Tpa3wCb/M04FpzfvR0bIp
jp2fgJAttb9kQfis1hnFqXk+yMCFbwP+EnHtqvPY8m+Zxj8GcbjEm+t4W1go86Zm
aH3mJWPc38DRxzU8pO6M6mTj1OaATsfpYjsQR1aCy+mXDjVEnmWnpecf4P73J95d
7LGSgejyb4k72z3rAqeSzvcV/EZ53H6kGLS9Z+RxO+8whxb3cZg1CThrbyzG6B9F
3q8jA/BzFpdKIYZwDiDVZRWtay9tH7Daa/lhUQYqEGQdJb0r+Oo7Mnx2mSuDYg4X
2Okbl1BRZ2lrXPrOwR0o5Oi8PJvrfIJQzVlrriBTxnL2z86WMYXQ7YvXZiW8lC1v
NhuyBbUt2rsbC30XReQpjX8IpCko5QxOzFFj1dosOzINSz0n4TcpqRntDIgKF8Zz
pdnLnGmpr/6zjUoT9H/bBfu6TUNAZw4d/cnvbCMOfXDtOZx9H1QxQ+P8CWUVWCUR
sO5OmJ3ez7ihwt7ksB+7fx12wV3w7rs+pw2IX2IhPQ495jraYS1v6VUsIcJcsb/g
zQZAFlRSPSP3lqVN7LUzJ80Hh45NdsAIX9xozSmhWTM5gbxfass/5w3LddWNoTcJ
WjC8uSaib4zDtOXg9Qn4xigIq/WHRVenHcBiKQpTcJg9uhdrHS463SqldSpB7VtQ
g7dNnAWv+L0ihjBlJYWRHlZ3r5XkPUDlkPmfgvGdnNs9ZtLolLpSTqmFjyoQZEaM
jtKKzqMJiaSoTIIFwBL06mk8Y4d2GOHSIfY74YbnXdmN39RVjHbkEz/DmzATU57a
L1w002S6ZdYFX1R0eV92iywgpWQ/+HUv61ID9kE58aYQdWDyZJIkbGclvVPuCkPj
X5OpTxwy+cM00p5KShWDCwSGkWccgLRHEoSGZHsb2osdQUYoycUQBjQzW0Bnz7uY
tlJkzxK6CKWZ+R5MxiGiikSYF2K5+DRiHqqA432A7gFJeebeXnGxX6KFH+gtlnHb
g0w4HmUfaGbi1rA41Pyw0xZGcmqBxeckMzAJjEUqyP0Mbh2GMu5Vw8coH8mZ0sHn
aKPD/4Pi/9Q7nVbUwhE7rFyYlM1mvuId9IF/I+oVv5FgmjDooJR3pXwSzl+U3N54
Ee1E4kTJiSNYowuqMyp1WEiVEAiUYKBOlaaa6BoheYQe5pK7H7brJ+yzbNLbJPrq
z08sdJ+YhPltuHKcYCnyRnlAzE8eN9Oe7bL9mqAUDgMnpnsIp+DPRbdITYtcLsq+
pDt8YZmg/hfnclhRYGKVIQVKzTwTxLlwdKEyG6LUeyjvBl2Cxp+s5sF+ATgxFNcL
iyfNFiR1XSGW6Ee0AGSiw+h/DhzNBfojm9q1KkwzBU3JQ4R2xF0XRER6MKXnVWq5
0IgEC9YjcT1Os8WeHN5XfsgVKvQzcu+7p5+lvN8vKEZkaRoJxmxIZXRz6CyEtSOc
k1ucnT1qCqlxkAWsZl2bjI3oo1n2tt3MxzpUCq0qQ33YNBoJGdqf6VDLobteyhox
O5gEBYHnuVdzwk3CxKoFcfQ77Se83gwXOTMv2mWg5PROx7kv1lvDJu6naLSdWoY9
bA+3lpU+bsOjkd1UluOKPkoAC2Bts53bjMTLcycVyJ21pzg25+BpVzhGJh87+U7Z
wwYOut1NiDZjohOeuw/OHc/OvfSqFhVyKjHS6IaJOysmM4ly3E/chbV2kYnugNr7
w8yDkrvXssEL+ZIiMB4oEuc8SeuD/rjEZjBRIGdc8Kv5Y0gSrW9CDoO5uNo4XDN8
1BZrju1zr/wD87MKTqtt1G2VJTZYnJG+rlm3pASEiIslieNXmaSjC1xixGWgWH3U
rABn2dRz0uc1J0oJyorR857FhYP3+2tl7NOGSuSv4JvIRRWE7K1NSs/iTzl/T7a3
Ys7hPzGVTw5rMoOQ7Z0zeZmy9y7MksD993bnDWD6z4Z1OHvvCmBBZfd5qIaaT3Sy
EI/bwN7sS6qJr2mSEKlH2JKFdHP9TAsvYEyB9xaNypcOkbfkHBWNF4nnme+L+YSq
n4jA9n+J5ErC9RQ/QK+BSYrrRsbU97fmIUwJQDyPkAqHkIHXdJdllDEkH9L9dPXR
AOiLqZg0SLPUxUmMvcZPB8h9xj2X0lpm3IEFsBir9vAOoaRWcGIGlsxIrda2hfQ3
ADlcktIKVY+t6nWTsIrNScQlP78xjuuG1WyxDF/PPeoNWN25QImiraF7NLe3LJ7U
Sd+iQPXbwvoqZZkpTrybUkOZdSWQRKRym9yRp1Ev+D6XNBFq0H6e0KQ/fCoqvyJJ
t5UfZHLPSCX668O+9zJt+KFsDF87xtMWaIsZMaTuLmTMQUqfIQrGIhFIClZsQnQc
bYmkCT8xKiayO/4qb20RDaV13lV6jan5jMMa9i8U+JWx1urpA4dZVtlKzqAqVosZ
2qWAb0td5oKu/Vb/sqVWwpFFxSy+ERg207r0hefogt1+SxzPoKVCAKRFLzX1lipe
/Yf4tDjSRr5/Uwbra1bRIXCRKKD37M6M3glLZKzJPnynEXcNzxa+Q645FsYjm0cI
AHsspfLFUuN9u20GUKq6ZGoFuzHwyk/9dfFmPqQVgEJ/x4qNRjt25EOo08eQAKKY
Hx/KgzKPnh0VQDFSppUs662TDo0drFfYr0m6OQzpSY/B3r/Xaq2h1pVcy3PBfRpd
M1ewxu/ef9ThnvVYWyEr2sORsjA/jHytM8mKwpk3EXj2Q4XLsErwkf1rBd//O58p
2VYdnnjUYMzRyNVsnxoH9XRM8AEDmHu3siNrQD/Sp9JkM+EYz5JZFSKq23Q5I0fD
gT3oqsdBugkRPqUtfUR88KxEZ4U7dVI7bRM+oh2yeHi8kletTH8BVW/hFNxvXBhQ
GBZTVSp0ER4I5RSnH97XBt0nABYDC9kwzjFVkaSA0v1NBHIjSdpu8q1nEedE+bri
F+Qi679l+Chdm5QxfA4HUvKqvd3pxZ9nR9Tol40LKtmfFTJsbPktkU8Ung4VmQ2Z
NcWNEgAIx271ow+W+pHfAslCg5FZeOrAFXCgjECUrAN6w9PJX+YuINrHLIyluIC+
FEdGFobRzGjfoFPTiOYIZR6G8iRzPLqprmFyJL2uYQVfsDLbdGAC9Hko2hmvY0c4
VQU8/tel9yGsU37ZLD/gZ0mXYTGOVH8YPMQF2X8mdR2RmhSkMLnaFj37dHsQAMwR
dxqG9SIWnZY/B7ePhjfLLiR8mW0yd3/ZD+4Ozug9nXTxlF5hVz/IzHsHXVNn4Gw+
qX4e3840suMdMJfw30Y1qDM8qSKDhDLMx+DAh9Qd6tbpX14+9tFFxAbqAQ5HZ/0i
fYqIORy1w8x2fT4q2J4ptQ2ujDVwq9CBRrTofKgzu57MrO5k2Yvje2gAZO8nEVLC
zatWgbhucMJvLvdyxLIPpLfCiBx4Wv+N02BYxer4Y/lAukjHRRLhgh1q6pMQXF0U
wztSKzaSalwySEdiFtKl00/MIfq/W4BPJGhnd8Xp/ni7crcpzFOMmIaXabrduZcC
MscidxHlpDvB4aRDXIlkYrjwuMWDBWnkYsOJmrS0rt9uMDyhuHTWomNsZPPHP3/B
kQwCpA2jKq64Vb71WyGNCNyUnASRgbU9DdUHFRi9VMyFRyJvGp+RhuioTZfihoou
B10sUCYKH9IZ0fMBkNA73jElfRHH60vFXiI3OLl8SL8HFGpcyhHgO8KckmanU1ff
fZROR+iz9BZLod3nFA1xtQBrcUs8KfZEQTnL0JjIZdAnjHvaX+JmmjZ4rr1DMSKF
uKBv2v2JdCiMy53P46+OKryPiutSaWorHs1G0PeNTpUuU4ymxzf1tb6vRV6WfdKY
/3q5YZCxVq7OK0Ib4CEmdz9uNsektR95N6zCQ127ZhKfCc5LtwwawaSUyDajUcIn
GnIdIGpDq/EHw48F7zvO/Z7bw84VEP3x59hB7MGH2HGpLOb9eM+qVsfcyCkHmYbH
tLNLpgzaK6pvVbR1TOHFXF3cpBvNJW8iNzAsaVkPiX7T7ULsRv/MoXWYUtw3mDz5
ThxiXXEvQpG9WXTvcJVY88thtWcfe6uXL1mfioOSWptsrhWxgRB1dCBVQJ/KX8hz
vKgXE9at71JUMcsDFxcQeikQlubs/fcBa9jAEAtsEpgQS86r3+S68bzPi9TyOZHE
T8K3FNeNqZEzFQl4so/xK1/Xd4+j9I3pqEwhcTA4OZszGA6zlxt/CvuO2gc23foL
rkaFS8y1MU/2wiwtGN0T5H+MviiuzEt9gU8CmEBl6sKpuaqjXP/NUUiNIsqspVXn
D4MeBk2NOatmwlvflEaqC3cX8c9mNUZAu1RgUYSuLSk/sou2nHl7NEFKfa/tqnwO
AF0CY1zHT0PEDBIjp59HrQqeNUhHCt8QrbLk4s7epzskr5hA3xbVyvkmAxoPUYfs
0sG8BA0czjjTpa0hR2309sbzsvN8eG+YVfsDHV5RSEuWWqbZWawRlDxuW0f6pszz
n5YqoqH7RmH9DcV9BImvJL2Fihoa1/sRIJtybvg9DDMicH6hzgheJxSZGCKRNIRs
YhvC1BTDPBv0hq4+VZ82edX2e6ZDdCGD5POqPdiq0KgLG80K29NXDpQMDUc6ZIfn
SeH4ph9OenTuZH2xZRpNfkjxXNjIsF0Ly3KiPKrL5dNu4zrZRbG2FfYVhr14qWPV
qNqlhZ5ygdeNeoZMutC2LqyJVqGIuFIJV/THLpSAmCW/w7DBtKgZM+8UuAJ1rwte
Cu+9GcRQAJVDXNloNa+e/tELVu01/PM4Oxz/DtS1DpBLh2TDCcaiMmfXLCwFenig
X7neMtmO/72TiUiw/wP6sDvLJHKzksDsIq9Txw0HnXegYYrYmMGmewR/bfv/SQJg
r0No8e/gniDbvNCJAwdrl72keNY9xC20XS7Ubh7mVWOfF45J4r7hX9QBmv2NcgnV
pVLu6WjM/iiB60GQn0hIJo+0+QncYaR8uSZjB6OqisGrQlhAGEag0wgHt5PWCQPP
fAFCUlko12OXqyb68Jcn+n3aH/Q2ceUId422pJGyg0fMilB2AUrUvof5qTenuS9q
pc40bYoaIDzPALXyQybwQ6DdJzis0qYT2NMwBBJ0hjyQzG4cHBEISplOTGoJwldn
/bjlmMbklse0kTZEtrFeJFJ3y11oHuN8EeE04BH0Gd6e5zTcnfaHLsZ7CtgcmSfC
+YZa3SvMVN/8TEu4wEfDTRyELs7osziVRfkOVdsD6FrosF/PMdpUcJotohN4dY3J
XorCu4MGsWAvoHIwvyQhcLB032cDXim7IsD0Gmpg4PSfpInfw8AmDgkTz5AY/GFK
Cz6npSLOhBSdaSNW2tDt0Aylj/SlO+7cO2UeVadkYQ83k/xYJ7jrkHZDQHcS3kfl
kuHqlo891pdJ0/6JHVZFxNDM4+SyD4hrSnn3KfGw4i9+VHdhVKBZNsTeBrwgXmsV
cz5du3mo1hg1TVPblr6QMORr4vxiJyv/nLOV10KeqlLOKRNTYdUHw5NlNC7DfAD5
wBFouIojEP3pQwgj2w6KQ9lFjGr0T2RfUxxIQXQ3aMDMQM4mXx5hzMztYiGhRdmn
7jQB64LZ70KVKzpOPDhFuUVYLIv2Xu0IfTGi/08ManQudQii8hNc3TOV5Zn7mzH/
PVQRqPr6LseFP7YfaFmyycwOifErMa/JSM8ye5drLZS8GXNLzo3J0iDd7i38HltN
Zx5SKmScYAlkkGZ7INjvadJxwtJJapDQ8EQNdAzkvIoRGRXXDjipx2u6oKEYios+
/lM7w/abA2GBiLYHavSGkcfSrDgu28W1Bj6ItxKq9KXj6gY4Fr7wdLY8UQQLO5ke
hcodMCyeoEpkNMju7oEVoZhNayJT9sTZkx01PVJcsYLsdEnyYTtMCnTZFyo+5fcY
3S6fKkosJ4OCxavVfe3leH6xZioyU1p2jBjWO4BcoziZ/6U+NCi3Al9ITrgp4fC1
VfpTBy2dBOigxNBR2jmWxyFUOBT6bzy9Deq4HoziyF+MR2dExXR9uGkNRnm69UHZ
dpPTCl8+PHVZO+HGVHSLhq8OYsaja/f9X3lMxDsc+a+47WERFSz0vS++QvyO4McJ
xgW48v6Mmx59veWuMZFRESojoneSDywnyU+gaQzE+LanH8VB8qK1yTF+HI6lkiAF
VTf1JPxWM8nXUpgKD5WV7CSGVuEl66PL6zv2jQCZXMnst0Wcjrk/sRjdODL89N9N
QMksH2exVBeib4LIutB14vn4VsSUv78N2otH4W922G7pSpbMri98nwKfxzdsawmh
k3zj6JXUa6qQ++pedkgtXPgy28gJ4MCWtdJrK4iOJwaqHyn+zz09vaNrW7hdEJbZ
5ge9IoSmxthFOmI6DH1hJypjbXx4PrBWxsThIk7HmY5q7UgcwkMyJ5ItVtHcnRjC
I4q2CfjSNXcc5Hpakvw9yTvLANIjEEmBLA9PruYb24FcvxaBPgUi4ATKqG7+N0cO
iQ2JPc1TS3IifkNM62Oksze5bzQxk7Odwqnw6fUtYLn6z74cvgFMNnM1eCVcR6ST
THRZ9mzzcVGL2VUmymIJw3rwkaREpqZxqRmcBG/IB1cPXFLAtJsyDsUvbNsQvadx
hFZSk47ehpBMnogUgU+IC8DV9jVKou6W5g7caxLKspNpkD5AkVbCiGpIaRCWXk0k
66cVzkmJfRtC8V8vnTmwB9Vj6xa9Z6noQpaYQMDoYmoxTuMMuwS2yddrBu+ZI+Xa
NP7qw8bzPPYfnzHSfOZsX28RGQRHsg5tSJyoAovKCK26N9nqSP5vWPfwuDxzknp5
mtsCVOWdlm1Uas1KdRJB36MQLxOxK6MCp/hE7ZBCg/GZFVWUC9UWs+K1YrRHya3Q
mLpD3lzWertpytgfRI9aeCD4J9hx6hs63EmoJrtiobflRzmeoaECO4sSv3XTLqiS
wn3Wi7JFsxnFbcqnjTtlfT+7V6g8SrvrCJZPpOzb+4DwYc6RmjH2hs7XNLyAwh2B
UfaOjOuBWTJb72DUHmcrTeFCdcJ1G7dbCGoro6KyVhbLAgva38y0b6rVhAqB9x+9
BIsMdBy4IjUOuhXnayK7xOr5eLBNcIrlTM8eZct3+FPwN3xystmaQPvrRINGy+nb
STp+Qr4LuKWEeLKQoAVgRkNwX+6XPJOrdK4aZ0jMNAGfb19CUlid4rIgEUdrFrzx
k6y58LseeK/7iMQ8KxXrIoQodjnVmWo1X/JwrVjblzEDX7NCc1gceiVNJ4E+Mz2Z
+pWdJ4RJMgyfX1Qw+8tFfeYZ3TjWGaHDnhgtylRhmX6jkzm0/JdBoeBs2V9UucUS
95qs7ltDB8oeBAb9j7+sTqhWBErBo0SyYfa7amq/6r1CpFN1k8FgC2cmGa6ENG3E
ypm0s0TQgLk0tNvCFGqWW9BhfD8hD6F6agopvSWPxq4ZPSBuNlC0gunDE6CiMd+O
0y2W8NkX2MeF4dg7r1y1IgSU5M3+V8+n1Lp7rQd8xhh2bf8CCls1KztAJCo7lMkV
95m2vA5pvkKvoIqqbhM/kYSI8pMVaZln8uknu6VWvgjN1yB9f5gdiIMGiOYEGc/O
cQh8Azx1HiuNgalmDsIezeLEBSppBrADrHQdqIWnsaYtXdlRwDQgUOz0acMQWlC9
IL3m7VfIMsIopm5EJ8dpF+y4u4O+5zNwJiiqy7ECdxaGlgss4fiyPb6zDx2aipJV
nuz9fGJUo/+LC/PJ5hn+NG4ffwsz96+g3T1l5YnmancFFebCuZrsg1b/wynS7b/a
eSbkTFv7DGdWCI/kydPOJsEE8RHt9bvT000amkXcY4mNypX53o39DCXmcMdOj7Jx
zxq7Su2OcEOntXAKGye4J/WbCPXqkkzQI6w7F/tCAcrmtmoY9aIkYE1gVOEyX6Tj
Hj6Qe6QeE4jKAwsYY36TYXlVpX9YNy76mDqpc8cCr7i1dcbTH74LVZ4PfNF70z1W
8r+DhYIJuekbP6ACEg3YzSPWBleyPPbHJMNeug8ujNqRVaxYZzWwEFaLiLIcjp4V
T/JLKievIrTzxRzYmvqxVeJuD38mQDxYNek/x1MQG2ApFih4+4L+FEN9voGq7/9w
osIzCPz0suigMhIl1ehfS1yrXokDWTHPFNWA2eoR8NLXEBn8wzNw93skRADyk2KT
p5bs4QvSh3EKy9WAhhf0KqmcUc0hNpPjwITYUzZys/s6KQoGBl8Pw6Inxd/UxUG0
Shi2gjT7K/K0KT8khi7+RQE4JGaqHfUKH6LAodBK4dEQI5a4YYFnCg8SxM9jvHil
2+aCBvci1/mjebC6vfMVnU1Mx3xcumoZmzKl9u1Exnrx4GfFXm97lZRwkPl4wwYx
zH3b81lanR/5aadsVQQgOJE9piCl5kKba5arpKU7LMzLFxxTvOe5G9QBa9QxyjHs
lyiQb5XAFoUi3DdCzO4ToCqK11GEjuTeJr7DnZmXrATnPKUa3vQvUjUc2kXFv5y/
qIbqCc8x+8U6Sz30YJWCNSk/jBdLP8cwq40BiPnaQvaF0SO6ollI4Z/vMw+CajG4
G7CXxXanS0UBVshkSRDWb0jblyxufLGszr9RfWfviTr7BhZ0AerXOcZMDDiEXdX0
2WbWgdrJOLuZ45ky9udp8QAwN3KzsiFpLdNgOGvhxfUkv4DPQPis8uMIqQOfnsPo
j/cbs9TyTnggIhztHbfxgSdbbuv4qVQ6rdGhwS86a+Mr2EnSBH6T7qVfuvZ9gbhP
RfG9D1AXpE6fJytXX2soKQtwH+1MsnTnDR5WBjwZWAWTr3Oy9ICesWom8fbIm0q4
KP2K6VpQnCpaHznB/diQaCss7re3Hd0G6yXUEo2GR6itO74wglBGw2r6iVfL+p+x
fmUFWISISXT4SaG7wjT/r2ShEo5ABXmtma+ic1lgeJL2FpLDsm6TVIUqAXyt166R
8zY9NX3WKDrwXXGgEv0w8hqCdMTKDKVHNJtk4xudbSUlNd20u0YdrfI3CfM/Mx8I
qRXMfdlHDrad9KHsvl36qkpvbbQjMR4uloeSUfYSSSNGB0AS6efgFIpwh05hP/DJ
oUH8nUgJegCXRkaOTmsCbYbZ2w/4u7V376fppdkJYm24TWQ6NMvbFfYKEi3OSJ8H
zHyHdFhNWBAdzHvFevdP8LsH8x12ETsxRhpiwsz9pc0Tbm5pdc4CbFFyCoVB6bWL
6LCqzRmhL5qSSXwMn76FkVbN3UzCr+YNFjbwVWh87tBawkXvGcUyQGHc+yWE75ui
7ruexza4e9CwcK9NtQ0jv7wsSaOs1uFRtNTkLVtRzM3OeMXr6gdzS55ZIK3PVq1M
l3rTnMJJXekOw7l5vdGW6F1gsJ3gcqdecISVscl8SdJ2TAG1J80sYgRaCQGH/D8U
+KIrgIaIRmXU8GKAbjatAmD2AIr0Rq6olAtoIBeEsr9BASjwfANlv0dySSjMqLhd
v8WfqedhbGvm72SP93/1nK9RJj0UW0pn8I9CSiej+QpIw15XBBudT3Qrx1/OSj0i
ri1JX4C5NAC7Vvfh3kZrxIm8E6f6KE9Z5YYQOorjYak1gQhoALhDSWTUeT8te3SY
0iniiAz5QngnvaGbWDTFYP2oA5wafkVTM2RLa5oDgOAS9zJ/5o350syLoo7zSFAa
Md0vU+eX0Bs/9nv+g787EG+4cAS5fVCNOc4QLHoqIfIyGdua8UuvKQJQu4V7Djm2
fw0h00PztJbqFX4id+YvMaCZqFAziZWm7f2GDO9T6V8Ochv/r2irL59sfUnYo3jh
9C2QqCxnkpit3L958hkhMDL/9vHh2Y+RfBuqTGgibrQbNRcVwCwvZ8VYPUJqe0za
0FWKeDYtDxMTkIDlsujXUATSnnzikqcJdkumwfI1o7sxJkleFVvH1sHRn4cTiq5C
TwYkA4LWTOWnd13RsA3nipio5qSlerShvRDYO0hM3ifswJzuPsi61mISK3wDZt/X
CGW20nrjbkNOfo78R2QVr37TElmMHjEnv74ccWha2r1aSjPhD6PL6JmYLiG9WjkZ
NEIWUt7vnUDv8rzeYE2gsgmYzOsBA33Q7neAmn8kjUmwdJI3M2Hl0x3ydCQkwSpt
/Na7ZNZKoFuoLJdUvbTkDmJtXhNOenBFeeAE4o2kB2PyezCb59+VnMdmWg5Uq4eo
ZSM4OXJwDNoPLuhuVxfoAuSFJTDQ+Q2DqwjT9fLbImM9wUx/kf6dfaef3QHxRkZ7
aZzXHxrRIQnatF8Geau8H9w5Tt/JWXCKT1N9O3zzTQs67MpeLI7UwH3klHs+Myb0
AxTF/aqux2AjDmWXlMgvB8WbMtE+btxhUUKGCAYxw45/f+VKWAJrtcZDlLVsvIUh
uwY3zdwEhWre2/TWpqFFeS+wXGaK4MuuOdDtfjyQ9e5aRkSYVgYzcGBjY+0ok9mD
zcVLCRZdnr3L7XYP58CVkoGJJ81rg0qOMI14hzlNPCEZ9UPO6baTFVDABDHtm0g3
ocEO83SnobXApTg1RtJbl2TSZr4xCd93J5K+L28oTaPyLJRytFoLzDvYWg3kZJWF
gq6P3eED/k1pmBL81sY+04QJhJI6CrWB8bHLXAJ9FvZTLFHg3p88GCRnAAFBOSAC
ALmGxjHm01NDhpjauCCqc3EoeGL3iZIknt+h9qYO7bZ0i/3JghCD5CuzZqd6QpTF
MxN0mzIL09xky9hTqJbXTP7UnBbyvm/e9Y8Rd28S9EbovEnp8PgWTQ9p0yku4vGi
lwgWiseJ4w/6lZ39pfkp8YB4j2U5TgFpv7MQF0yTJgygWKrxEvvKkHz0X78ELivs
PNNWAVQHjVa/FbO55TUIFeBfkAnveLxTIQNR6wV8wSw7jRBXnJ3ovjYBl1OJeN2Q
cqhWvCdrcGieACs8rOJGFr1fPFj5k7USrL9IoPfZuV3G2zxNS/kA5qgB72m65nFd
z3AHeN9i7NPPnhOhsiMIkBkEuKtaJAIKzbOna/+K2/CrsA4eTTThBO4tqB+enWDq
iVAYyrWM1QZKaQwYoU+EeXi3tRg8cFxCphuFY2bYckz1bgvgVplpgi+qMsO/suRE
s3coUoB4YS9Z4qXc9p0sjaP4nFRVeWZgEYol5WpWqWczFaDCZpV9WkVsm22GGqOv
WHsNI7KNte6E5wx+0Zjim9K0PDXkMlJHU7Clr9qaNF58eAZLf59jSHkJ4+4vfq9x
uFl+KvsYbMhhke7fNKbJyOYOcop/oBvXqOYIQokObKGHQBT+q2CSvmUBQgPzCMoV
GNtTDjY4ZtnA4THxSsliQnMok+bgTyp/gj3P0D3IpTYpNNISd+MZL7zOase+nBSB
E2a47+HS2sI0a1e51jQ4yxlHs3dLc+BfUyfr+CODhY9Or3zFJugIE/Xv0A15vkZ5
0OFTfAR8IbNkEJ1TqaftBcEs4J3cN3iTvA3+vk5oiwgolz2GecYZYJcMyIS2fP3j
LX6FnNNomNGL6e2DFfT4xy45M9G9PXREMKWfFAOGtOEpBtdVVFNAVhe47/P5UGkE
ds7oxB7BoEksTOmDwfjIgrfPvGGLP0qMy9zvo2HnrMVG0n4GnvRqUmYqM3JiGvR9
PKijpEwQW6TCpj9z8J2F85wUvDjMjYAa2tzBFtmTjXvhMKI4BiWL9QL4x50IAMJE
m7MwAL+6zgi8SIBZ2dbOL/J0scTbwBXx38UrPfB/WIKB4u8vVmrLimc6CAby0ovR
czYdagHYHAmJ0G1WXjkcbtSAih/2ZP79DPJbdM8NI7mgZCMNkon2ZtRfL4/3pSBi
rCZCNaRe37UaRLNyIbZ/JDvjoGMg+utaawTH4SwxoZUDT1QU1z0cChtCmsTmDk0M
jwKhDAURja1LVAn67JUU2W2YlKlgGk+xKSfdVK8Pq0emLuu0VOPtkNRGc/d2JJFT
GOh1OJPCcsRZQCWEDPUexWiUaqrzeOfJQoEo/Ndp0ejkaZXdDWYaXjVn2FLvxPX3
1I8VnemzqxW5hSgWc2EVRZlMvw0depSKsHCVnzxbpoSux+eNsQ5qGv+VYSwiAE+R
deIRy/RIbC3DhWOeUDcBPNcA9KC723+Jd0dnfSOimohuaGvfqC4XXU1CHnvt6JCs
bdHNYaMKc1vrBkiM5fPias7gE3gseVgGbNC9JJps2tcQqeUV8smC8GZ9CdM/1Ew9
hQVKqv8foPcc5is6thlJ+cyZ2RpeLAupVxayfOC+Zu78OW1/bB+yZxZaswiDwQ6l
SzobXo3QGh6rJ7gGlxbs1Coxicjl0bFI1Gte1dETeXSidtaHEDf4IS50MI5TKmxk
Ezp41U0WsJoS7MtYKSC6AH0ArKLhlknEtAlAJ7uR5UVX5M9cspyH3cjK59RZnZ4K
qZPiQOzMR+7f6new/rBMS9x8xtrc3m1IXQ/sZ/yAVUI5IRW6zCqKnqytWYffQSgX
sFV95nE9s6mUIVYucRNLSudC82dxDwP5YmjF3N1lZ3cqbp62VuAwZ8KHDxhWevMO
v7u208+P7TzNOPYGjZRYN8zKF5Z8Rkcn/eP2lgyqT/K3DaxFO1fNz4trquWlVKLO
q1q48VrjTeGnlQVVVF5aq35+N3cI+kkvZIOQvGbNEQnLIezIS00st50EF5TZAV6O
jhdA84aUK5TUi20Q1bLDr7Bjp/uMFdlRydQsiH1iwmUyVCeOjcrGVZm0nKEp4/Jm
P7eeiAqXBmPcL5SDtaSkv9Jo//FJFH7sb/VrSV682wTGidOK1Ubhjb5luDUWoEdg
V6VSATCrTTTUYDZl6HMzaTC4zlesu81IDboq8mcc2c1/rNmL19xcBHIBkA4Gzl2o
2qi9iaXaEMe7Qr+DuJW1FmnVBNdcScJL00qmsVm7e8AFcWiOmXX3Jy+mFVSu1t3K
VGGs1FIADjtFRreskKhYIm7GWzUG2Mr2ym3nZJEwXuKAniNRMAAepLy6okApeafp
uNqlZLdKTMi//NX7D2lTbNP9pwHTz6TkTlkOsbOqDI8Tcam9qhPJyVi2hcJ166Yi
FlH5MYm/+RwmlhadDSp89yS8PbSJ+XrVW9coJVGptDkImC7Zl32kqRVwbdKn674c
/rrBdUbG/H8kCaIlzhmgVmSL9S2IqlFLHqeyLZhhISwSB2FIG6MiwzurkTzXOX9r
n2dSPoB3LE9Hx845neVPfegf/U0PKO194/paEUz5tSAHTeGpe89M6w0C5X/fNvHY
cTJI13HMDlgEsxDA1ABnLzLuiL+wivgy9d2d09np2YrUrkVlA+PXxfYDdUHs/fI4
tBmJjFenPJs4Jz1kLdzib+20krpCcdUJy87DjhdQkti2DiJPqsXK5/QKMN3F24Vf
kqq/9aY7dE1BbedIID8GxZf3lK0RCnypciypaKnubNtNoxFnDpByJ3JhnLf3Nw+7
Vmif4rUp4GyvQe6wdesjUvw7NdDbJMjF31iCxulhc4y5u1MgDuxZRXLyM6xfpuSl
Upkc0mhVWa8S3eJpzSxSClMQ12nLkmM8Dxn4YDH+ohd6SXsV2HU10tjLZkMZf6dD
DS1dpM75hKbXAiSjJ7QnzW3HJ5ulKvwkDrqLMs+T32ArVfHfsLras4RHvS3SKaGd
Q725OgN6NF6dhKA1JfR1B9v3uklsHOq0BJ3Ixp1JFFHZ+79n9q9E3hpMdZZNSU6W
FGRWroHSccy49pMYJqBLWVkg1klc5vcQ6x6Xl4Zii1Fde00UAZ+ctho8n/UbakxP
TkOEW+LiqbQLnaFWOi14dTed5wZ1lX7q1D7XarEbTn3U4bzHQRJohy9ZqSPMlEf4
HH3ROMbNS/ZC9aaLLpPkGLFDSVq92BY4zBGzgLilXJSI9SlhfRjpS56JWQOnQuD+
3T3/fS04flXmICTmrFlKL9IxcbnmYzjM5fn997dHPNpBOhxIP+EU/MAKWZX6EqhL
XYlVmfljyUgEHXx8SOp1PGseWiEXUIXrOcQgJ8WYD+KowmGWJrHKunCjjt7E0zA4
AHVRs1XV6fmaoF5LAwZdJxVDhOPYIDLg/U6FNMBnWZf+v6MPD8TpQGrAI3Nk9dT3
31WfMGlKhoJZdmwltrnqwZb/CgUFnZvrP70iKHkg0qnbQq3W92ZVCwFomTgKB732
f06AhYArhk/2RD4//sZtKcx6PyGB4InznmgLRGSzBWjXKHc07cMPpBkRpKU2j+Oe
QkFbrGd5IGJwk51Q4dJQo9VbP2JLiX1cHUBXF3PyJdEIwYO7Ya1luMAbQsEkhI4X
5FFBXirhFn15TlWYqLeAkSTvnk9YrANtoV1whOQVhyRtJYVBtMkRiK+2Q0mDGChY
QD5x/ZOBAO+OmWhufE/DX3FS4e+ZaxzcXMyaxAXOwVXPoet+axiZ26WnxX+HSk4t
I/dakqb5GQ+H9NamcmPA+0iXQk1xVSvTWd8dixN7GWF9DjclvyYgKFe/JuL6VAuU
F1R7Kgg6p8EISF9RHeKq2z24DRRCv6McCR8ys1qAShAWMupi/VrZmGtgMMb/4dYr
5ZLf89n7FKB+oywo3xQvtPbCqrg1KNqOaxHpR4Q3Gmf4KKTJj2roicG6IUrr3Qdi
cALUZr1megEtr5QAoLmcfqQ6ff2OVirQ/Of+84gwUUsCQHC67ij7Mvi+vv6P6KWW
/XurUYgrved9nfyVW0jnLjnyE3sFMhJXRejciaSAY6SihK7rlRZVJue/MjC2npH8
gwUkaQfm8G79rcXegJUVC7m9B3YfNmRpm5SDxupKUPfHRKitp29QHxI9zGeS8evD
oRe7B1Q7iQRTPu40UtGMeaCmTDc7KXTIJVpa7NojHTXbFIcoiYtTgDo2xrobHuin
vn3GsttubaZLKj7tgMbCBlfV42VAt0g4az1AzPIrOYRGVFwTzr6vJss6xdm+w2vL
juqDSQ3PT5toXMiBR9Q6yScd33eBALVwVK78ZEi1bKQXmkCLq5wjSGl7QEzThcuI
Xmoyw/5ZTvP73VtXMg4aZVoS95izYgwV266kwILnqwRaPdt/ymD9naFy/dzsigzN
LXzUZBIy5FEw4s3PwL+6w5ofa/WXtyW5WRfu8AGyCC3aa4TECZuz5piFE7siYVoM
k8L/p+xEMnU9yIkR2YRw9kULpttC3G6+HZ0HpiZ2pvnfzmQNYy3HU361CTh9it5E
Cv290dgLIK3W8rarVbnt2CloMUukA2Zx61j2ZZQSPuZd/NaZ6L45U7XEn8hxAqXa
vZPp+ZOHd6VuFMuCyPAbH09oN3j7m9rmdHpKnocFb3oE256xqbnAn7M2wl2XQq1A
ry+fwd/GFnY0l31ZfPqAPYPBgdM9tIgfLWM+wtGHADz+LQYRVUkbx/hKh4oRhjUF
liQbL5FdnZBQhKt8WugaFNgWjXB07nWFrVDouVQu1zKnxfx4plIdjhHTOVtimadJ
yiennx7502OrwINvIqpMQdkwfvrRMUOxC3nHw9etVbAGtdR5i72orChq4ia/a7xu
Q9jrkQ2ggVLxH6ta942LFovQjgC8IEOa6lhxDdODCwGTBzfpAFJZJcg/CiR4F32A
P58MCWxv/VLgCBlCblngzTDx7IMZzeDMl6/x/dABWFyhRSyNDnWpaWV8VjgcML/x
peoSTtwipS/1ZiC7wkgYNO1HU34KXF3A/XAxOf0FExHV4HdZMBFBITgj03BPktsY
Ko9L14Rp5qa4yViIe06+WifbIEUhBV18GtTHeoVLzVyqqKXrUNHPkLNtec8JWVPD
4lSMmM7uJT4A6SixXT/w3dzIjE8ejfIpomFfTRTiesAVniVjcsr3ZRDlW8txIX0k
uP7gFZKjI4looXPcwcz7D+SeZTNY4u4k1P8FKQdkIpUPtXa7G5WOF16nzYuLqNmT
BVSPw7IEdE0AruJn3NHut72VmFPCyi0x1WVEQibowFdKRTWB3HQicM/BYokldDUK
jPXLrW1FAbPZAg+aAp9jgbEjiFzOWNq9PH7mpIQGNqOSf8ql+1A/jnVcG+k25MPT
AnHbQEPDo4i806q5UVybld+zh7CIcOkgocpcwQql4napwPw7EkWi/1U1RAG2ceyK
7MSmyzX8CulpvJraD+/c+xTPjtTO70jomFjKI1WhqmWkj25DcvThRfzYHN4DYIaZ
3wgxuCyUcbTCwgOUmjW0oKHkRhqzITbsV1DqKSL2IZIapjA1Y6xsWTtg1fWMp8hp
uEddd7EamTDiFZMXwrpJoGqNRePo/QlXssOSYiS5WCMW8uSIgcnJDExJWf3MErFV
33b0TbTpGG0VBTAVzDYde8NIyaBIwakmXcqn3C1vg8Mi8Jh11ccoXbrjNzfFHQvu
GdAUHuTeQvqCGiMUWUSB3y2ir0eHHXhCpQ6wVR4Ta/6n+VVq8mdou0VjHRrxMYhA
pSesVIm6HFFdLmOcwlFqo1mOf4j2INm7AIwf/7/WStC6HfSqT6i9TWaxDbUaGhwY
YuTg3PWrUt1SZ5kvava9Ix/fma4Pr9GkX02Ja6/JI+bQIyB+qW5CbiMYV+i1fJH/
FJffNm5MfGHpIBR/vPG0yLxEsigX7UU3nKHdBgYquW5EnsqgMGM7DmHmejoSpbXf
k10MKo+gDLKv8E9FCmMSpZuXcIVMrlieewgMdH/AgwNKz8T0hJwrLwa4Rj6tRCLn
f3eQ/+8EB5OvDhtXdZl8fxA9ed4X+agOPLvPC7ukRbW5I4aqZ5vzBXb/AvZrZyUP
DgX8Di11AxF8qvfPTZPRUPMIxm8yPmMBjaNLVhPOUxP0NX7X0iN7TFxD3KaPIckC
/m+TTdSq+4SOJG7MfFNlgbOOIM0giOgw5eea08RGNB5cl+7wAE/+w165u2t6qAYD
iJybZ2FQTaAHOXUX382rPXTaPGV9Uyea8nG/GJVo3GEZYd0q9oLYCnXmmQEVA7jW
/9u9Rv8CVwJmsX/mqLN0EWOvCr/eQGywaMNFpHcTY1VX/7rXaigKhopfuH+BaSLq
YJXBgzc7NxfUFET9CCiB1leGYLd5g0NLSiPYNkVGDfH+AFA8FOBpkyxEVycGu8tQ
V3JrwdsO979CMnhwZ/P5FYiPyflkyjx7Buvylc2bVbTouFnNzzoG/8xPtUFiIcAr
a9sF/LrizwpiTI+RK4GARTiV88O/n6GALDnSJ6WcvPZLB7X9dXhZPIsQUuhDRmzf
U/uTqTP2HIu96EwDndNw+Ndcfls1F+zk+TEwL3KKAjZQRxRxUj4Q3okZMLhMUC0t
+D6rVQz0k0BpbYrG75ppT9Sup5bIM39m3VL+cBY+28kozo2dmLWGFgZiWjoO0Ps8
PJIm5KFr0MZMcMQ74A/8ozR7yP9iI4u2f/+fJABp7pD03XBEF7xeGDdjzOz14vVY
hja99A6s6Zxhqb3dCpGSfj1fgbClOpe0EVhV/DUkw9SCsGJyTT8+A81j/QykQ2CW
bXbS/VcIY8kgZQuJhQtrqFHEnTj/G1NVwGCLi1zXKgtGjG5zs67zYOluutZ8sX57
m3kY0Cvthe+A9ph7HeJuNfK9nwhpdQxZEwdGBr4npGOqrfhnP8IcSj4RuWeSH/NL
0UhMDDZUbR9mFQZzomWX+5OWn7w6+7osxZqVLiCJf/B8PwPQ3l/qSecUYxxeZIKj
wrOXtNv5Vvwtt/vS4vKNKgVZ6ZyLQJlqplyMKrf8ACHVfzf8us6Hl8UfnltQmduE
A6LJdDH39bMuvUwExIOhXcUV8V/YoDdyaHCdyoe6n2zqtvSyhmRzYaTRMDaLvBkM
TQYuX4elTE41FM1DfNPTqyl0MavpEiNmHWsfLgGvXq/il/9mHAVnsi5NJHKmaT6z
2oY/a4/np5cy8S9kv9tNNmpUZ2Bi/aIAJ+qZxuZnXlADRCc69kOhEB5pK3iTUHfu
B/I97N8BJ0ztB/aJ4WE6ePgOq9C0HPKjAUUqztwFBSFj8/pU5ir1Y2GYbRlDfDTJ
F+G/4ofipmTlAaR7hf2UUAKBFqAwWpqBaBPlLBFRP4nGnsZd0k/TotYKf/SJaQeC
pTWXqtOm12fz3IQrBMEJW9mAKoIVIBQwsXBAIIfX3r44Zn+W29a8d8k0oNLf3HTu
LCyoYiYUsS5Q3aJIb37oMxo/bLAsif3lnVARQf6zQjo4dvOeyvFC/GW2Mlvbod+V
Q74ZW+nveYHkrOv6DRtmryNT6nxIr2bW/jYl4C8fLEWD3bfVO+myTCcnbSVGRj7F
od1AIOv9EcLHqUNkkDG9mY23jdtdbX5hRBSksR5Sltdyde9TISsHAP2UoKtJm2rU
WQKO5rYFny2KgefAjGAogml3hOcyVQIu76ih8kbwMcfJkrBHg019sw8qlcpa8iKC
j2J3UxtJYw+smxQumCaTeZDYVq/jfaBr6Xp2ClkOzEelPbN2GyG25ePqZh3E4522
jGrvrjVsXgDUQboLgZENlzKqIxM4wZA4SCq/4KkcZVyl/LTPSKU+00bGNx2du+Ag
lDIxyLyxfcokjiItwfPAXSszZOi1y0z7u+W6MWyEim+BNRjJdRLQ+/msS0/AzbO9
LwFwodSSDyWDUC8rBNPhxqpylMhPC1DItTBnBfvYdiThvotfHYZ7a0z2SHBvALrs
jXPduxQaTSm23PYJ6ZfiKqEK//kxC449H7wYEJDtpxH7JxerHY18V8yHg6qtufDJ
3UaRelmNNTZa3WIOjl5tjkNiimhPuwfRB+TDXigesesAXq5u/M2SHaOuvxLYdcjP
l2HjQeMse6FqEFx+Ab4zYDjUpFxrYBQxu/0uD7rY48axsh33o/jCtTl6nHK1Q2Qt
X2Ix2cXgIxMujy98Enw6cUt3/EM6CVebdKgVrcF9fRB53fEDAHqiMUjjq54Xe83Q
Pv8z/aI3V06ejGmRQWmXyNcSSRcQpuGigrobg/USbpQs8ecdyqSKDi6sCSXIuxHv
mdFsUpg9gWmH7yywCalo0C/4w+y+LvBheOH+wIAOtoeTgzJs99bMBqkues9KjBM2
yLyWjtdvzjukZpPiRmIUrKcW7xd9ZM1diXbDdXFWRaKbt3Du+ZT6sIqN1pwMQkoi
HDtSfFs55ra9I7gLsOEDxmsRB4rXWNEC0bDF5GKixuzu02gco6wV08MrZZvxIxMh
8yL8AyXgFMP1hW4UkSviDUXXhq9ETj0SGChIHvmNAqz75RptL+vyVP3D0nARZkIk
iWzV2qZT06j0Yk0XOKbmkoazjGA7XG0UwUf3aqT36S3IF9CFnR8MVdJOk/hoG/xr
bTWRlg1cHIXQvA0VwXOSpAzzmmRR40hAaM7MYwHe4x/5KWeJH6Eju5LdYBMvTNAZ
xoQbKiR8NnoCc0TfEsS1uLjGmvTluRirjs8HVzKm2VR3VQ4IpRqwdSkBVRcOBHBS
Elw8sG3YFZ6Cv3dgDjFHfaGvxjzBD6oDOChAEkoP4X7eSTeZcVEN6Uf+pBB2QzKX
dwq11sSjTaYmnPud+dxzadzXkD/AWYG7wMZfpNGTNXg7xFVyvhbGSe8wUHVcADNc
SrTDxSG+q7TKFc7zZ1B8Qid+lK9UGoC7XxORhz01KyZ2Jmp3QxbZxMIMIKEpA3jU
h42N6/0k5CaEhUEHcTsxr09OWH07s+6+vljddb5GtSGHY//2/UVV6asq6Et1BVwk
zYo0Enshuw9pQCVlhuxyjFA2/X7qTVnjTDZPEa9wJfEMzUe+9fhZ6ZIh/1UqGZv5
feFXtljYgfajZjKzsldTcJrYZWhHYMRzIJagzHDTKBw7B+4HgrNqd+o6ZFSqlIoR
fprKz0hM2rrFoCn8gnvmQKg8RMLWj8xYKAeV6cFx8GobK0lNbgbaa6rD1eEjVEOe
FH91CcOmcib8E+FygUqUmkNHW3qQh48KUqusuDHVws4upyzY2NTWTr9yhoyiFO64
+NlTgk+w/QiJXv4kpre5CH76jzQ8Ugk5jVKGxjQu3sIsjpaCDM5QRTgCxio1MOXh
3iopMb5ZhRyssYY+pwf+OT5YQQ4D5jCOnJ1GAlbmXDMuDcpEASv6z95ZRiZsc+8O
5qm2sjYRTXbHgd4ofLqC5OVrO6P4xyvYfszgI0io0Lug+AP8tNMmWMAY908B4KST
65vt5vlmoUocO524ethPnVLSUd+L+OjN7FcCEoDDYzHUp0hrNotFvYzsAUReuJVF
BqZ7PXG7Ti6daxi1C5AzU8yTiPjTV5jr/8ZwqNaL40xwJQs618Yz8UO9atMCbFQ2
QCESjN2WHfE22eP+PpzrN2r1X5Cryn95BYn11giV0sU+KsFMqH4J5vJDVaW7L187
57AFWygj40Re7JE/Ak8sMud3Hpp8zGG5LBk/UYjNghHePWFtBNFZyk04Z1nWe8Gf
iMjbvu6Zv+WE9GQ2nEDqUkuCgLgpuCMI+XnnExangKUndQS1tSwfZsdSd3KcTbrS
NeBu+kZnjaPEftcmSMWKFrINiVqXRX/dzAhKsMYvnsIIY9FfdQL5PIOb7gPh1uxh
qtH2bdtLpCZrYUBaOTXl4slvliOB3rED0cWdJOD3XOR/TftbRTkJHF/xsTqcPs5C
iZXpKgE+LIo1wGO/nrH44QNMMiT6ao9UkPBSOzpC8tmohpgawdwq3FXY99/+Gveu
JmXNe00hC5wucR9++61i74ijE69meJm+yU7CdcVor8CXesgw8CVv6llkwiajRWZa
zuPvoEuGHW2zpOUstq5iixjrqiz9UBC+xlACXxtU7wXzLzfxR2Bym/z9zk0LrW7V
1EzdRfZ8U17/rPOXe0n0sEEeLDAyftM0N0QDwqut90CuEJYCz6uMzQep+21CEbjr
VrDx/q1k+eDvSkChgQWnQuRQIK232ZbQhlGc4dDsY4X8bgFFvcHjpgshOprAnIOW
fd6uyFjV6l3+fUbrjtX5pUDXXKFW+6QNzHbkdoKcpi70VFDYAwMiuUOvvwP4y9N3
iClzdzaIcKwDRFTvUujkZgMaDHsJwH6eAjzKve2R2TcfYz3rZKHDpyMSubgZ91KE
1G8qTYhpjE/pUCikwycEKnylXOkSGAsNFw7nfUIykBfaSJLV4QuepKbTgFUBTEek
fFNwWbgs7qqlC1FMP+4khkiygqpHhAmxWTD83W+/AaJRH6ua956KxOmqWdco5H//
hMbLHODmIetH8KK/6lJhzP40B0QtNJvYH1jdSiSDMY9VZ3VG5Ng+eeOcBT+a9ado
nR6k4w6mz5TpO60FFg5EQlA9M5NvfXu+7FopfMflXF5lK813retIeTRPxVzZ4ZiR
DLgJa5bgAmbETeXVpTCd/K0p6AMxhTcHhbwrQYecXTNuVGCed/zMicslhGK1hJCf
U3ZEk+NUnLZrOcAPWpSqxmieIGCXzB+9n22sNorNeLkkflSGnGGRNOVciAUgccUu
GJONhqdJ1FiBNPh0ctyAK31uajD3es/G0r5XIcO+NTaIWN288XAe07mN5PmBCw/y
UhLl1VGksy5dLkXit7sDnrhXZILIlNnlKhDzK3YseyZayijlF98fNpwAhOr0551l
2Ie47DpBAXzZwnKZf/NVatf6trrlbP92a649rfwMJuTZBuVFC5lTGGvUeRHVINS0
FEbuYLTtlktc/QI0uwHXYiUBrJ/ZxXEzqfSLX+JPRulIvIMkEfEPuU6/ksYKvfQq
46tf4mhqwYTIoBHQD2Yf2FiyXAJ2bu3ucKlrjSU0dY1mvuTTw9KZUgm7p1Us9hlC
iw1lcoMQWTYwAFyc8YN5xxRlZxAR9k6AIY9cW680ai+9DyQKEPCqJHpzfRxGgxHQ
r+EVm110/+aBZl4nidbOaEG2w/1yl9WaOBrz4yUKBLlRBshZQ7TPtQ7Me9Xy4FaI
sCh6EprEQN6NNBvLici2vbIQ1xsIIrpHBru9/6IXG96VZTN+x+1js+63JWnfN/b5
9JsnzX8z/HeJuG3Blzp5wI8suMQWiTqJxnBHuQg/K4qXVrZU5ckrsBP0s+FTFBn7
yURPBNTmlYNuOTBgquFO3kTMxSFkdLC0mBNBSWr7OaXoXZ5L3qzhtx+cl3jVbMm0
RLC+trsOSKuVqzYdh936ZPYptP2XXJuLFFinaxQcLqtjqPUsD8DjTT2fZ4gR5oTF
S/sby/WgQBrZ6AsFVdZH2enPNpB9i7YkVwj9cc/VoN4OLjgqw/w/CVUsPxio+JQH
mrrQsr+pVIRqLkzKjpP3FcsofB4CbceYWNG37plTrx6LrIk3t+O8/ozDCWtbQjkA
xTIn9Cc0z0sVF41VBHmP0sKOp+BaI64t2PUyyJGjBe0dv6Rv9qG8II0epXXVwmf+
jIN+afDA8kWEfgy+0cgTFk9hJDa5uiWfR6vFzzZRHhE9AbrHILse6N36hr8zJYPD
WjI2FWBdAmkU1/i6xS7zrWG4XbXC9gV7wJ16FXWtdG5bY/f/U5QqBu9o+ooVJlfB
fvt4M+cTEUCTMyQyDmP16lALNIMPe4gYhAYqEaDu5sDfyOxFZad2kevIsCz4x3A5
TapegsecxBAt9eYnhGaivCa9/vCy4/hAKMNjCWHPunvrMonveX9By+Y7f6L5OuKr
9m5eylxzBG7IVrl/B79H00UqtQt800gFVe7dnR6dPr4BumovWaKQCJoCkjaCdNiY
bmV+kgeGGHiA/l2pmPEOcie6VjkVQPKZ4dsjVLuPHXRxwPsqfjsLVQEJNQA6Ibay
Uj350LpOYSZmPVBH1tGCfNI2fmIrRO+xs29qkSz63C9xh5fhlhX+qCp4vCP7rGb0
ady8sfGWLsYxhiwkyQVvWce2zFur66CMCZDdDVRQtLg/RnYtSMj7JAO1xmPZ2qhI
ImaIc5Y6Ue9u5/qVlwks4zrGjz+jLsLy6shJFPzv6kj4sdKkTxy8dRFmYhKYmTJ0
6vVvc9EIniIczRIzQDYlZi4RzSmLNisr6yJ6SWd9pLcvoslBC00JGidIOL9R+CBG
a1zkk8UOatj4lvNTpzgcAaNfpU17PySORSAu33p06WVQBQ6S+BTyZ2qKM7tbW8gH
eLA9YBtaUvbgtahic9PkqZE94teZ7fZ5HVCp5b12Kznxz836p1OY/7zzQpTBZ4ov
C1gcIKroEyY9zifMVojPGKvNTfolydE60QT9hoRp6Nv/gGEDHLSf0U58DGvHPMbT
ucCdF46H3Dr7/rHceKgP9qipZbZkfnEkLqvmrsqeMmsEInXZqWUgEOoqh5UgB741
uR7Ffd+17qBEKYA2SAvvahPTSDJcbbFXgNV7b0UhDwj9dOlGqi6UVkGQRSPGAQpd
KwpYGI87b1gHlmdSPerxhqsDmODV3z5/JvYtu82/tAOX3Tv6gSW7VuEXma152YWQ
exxsV8w+7ba7knfR9Dw15XQKSrpAqQ53QqR2ZfL55Ub33mjktEMzM41NATo7bk6/
lSfL0Jo3Xezulc1Rvjkv89CHd1dZg1TkCAjhVJFxVOudoHjUfWDymiGxcvZZGK36
B7KjGsJmpow/NCKrTRnJlvZCTpnqZ684jayrVJ7XCO9fq0JcE/O+FAMyBGhbu3PL
2q8pXwT2xtyw17+9LK8Fc/gQ342IpXHVvEzGeo9jkLYE90Xf+w3jiCXqXWjgkQ+f
DrthspGLDoVOIaTo0NoxXRu2pUhiyz58CR6488489IAQMOZXuNahVGuibryLYxph
i3lX9b727clZV4Xlig36aPUOb+u5S29uFHgWDNu+FFrjwke2vUdHqiqKXVlLpXdw
TVV2rqXoLtau5KkVPLPVXa+Wpa1nIPkN1xR8fzkC6RUu31jVaomaqb+IgNYaWtEO
C7YCkh4TRca0zTbAvHNN4BJaoNtJXlK71htZNtkZhW/lS1av8u2zAydiU5bLkzIV
UkpffkUP3KS++uEKNIrDzFJWu1ZUGl13Is8xOu6ZH7JroXYGzb5CTLcbrR3eIkYa
+Hi1FYuaKHGzwSESTPu2VdUIeoxeThiLoDEdEOlYyG3pNM1roHZ3bSQ2tzUQE3ku
4gYZBdP7vJfIRrqvIwjON6fL1zUIIzTj8G44Wdqnk67i0sFiXRjef6izHmgX+SBM
NLVgqIWYJVvWRuC7R581e6kTsQVfEmH4zJuAZ0Lt/poSCGD3ZOeMqF82XqVSGTrO
zfDm8gfbrKdEt3SN5B3S/uHbaTC0GIjK6Ng0dYv2X7ivY//ODcoWK7/bdta2Lbwa
yzcE0aoj20zeuJAU+HvZRsJNtDuHNK6cpcgRVT8ibgJrK4c6nyLkW9A85MP/Mj+k
xrD4xN5Bogr9dsskAptKZA58np89DUh0wQ5sHsghF/R4xW/jhseWOpJ5LOFkMmDS
MBwp/KTYBbCZ1G5uShvtIJA+vagA2f7z/PyLtTjeOcikG0fwsl7bBteJ/ZYOTeID
qj5cjZ0KtS+WX1RVDRw6cRYIDo6qf4MBvviroZat2AE8IZe4e41+c0kfuzbsQrcw
WzyFew48s2qIzntAa13gLONXxODSa+XaEk7it5ktu1+zrTLZ8May22TiHZB5mqTA
0mZ6qiVxib+yGo2Jk9HVZSkupht8tAXSKEOECS6hU33lMeeEXDorN1GNsy+Mf4FX
YwoI80Q2YoomT82sobNhcNaMGN+e5tJ/tdeykKCNiaFVti+rVBEr+9xGP240jL4v
8eK0Bg67Ea386S9gi9Lu7G0DkgbrUUF+M64hV2CfKFMvvT7yUEGomQ80jk/dWQ25
Rpq/HyJIjT/BJH7Q2sax9N7S7Y4aldFfFpplWKugdAZt45MLmyp3gVkiwWoNRqvF
J/bs4g/mYx2eh6JI9ECh/SAtT7iXUVL9K7G+wFhGJRaDeU1QDKkj6KUjGxn3xWXs
EDzT3PU2wa6fmkYgq9aqkGXxcYLQvD6fe0j4Uu/n0IkcQHx84ldOhAO9GIUruhpp
Frp6ek2ECLbb6WHap2Fi+ZRaZLLedaX0ABDbPwuKX8jCNTCwOm2/fe0hydXlkX7W
tcMbrEZJ1LvKq/vePJ5eChvRENxHGOp0sb//POpaPvRUUR5jE6pFxbaq3lnRQiFa
YqR62Z0+lqrLqexm2ckm4YRdwxb3l46jTUQiCVtVsKy7NpzehPXpUME5WkcSSXYH
RSgQIVYNiCcAqitR45vsn7Jnd1HSUv+bKfZ/IlbCmsrzA+bCfIDEY7NGRSZELgWJ
VwpvwDDrzS6z2gaQz8ftB+sXikGFHlETdbFsq1elfKxR3rsO2gvbYaHsADOqqkb+
aY0w0FQiRQg0On0wC4tZnj16/dmirYNutJDonWhCfLSj01OXbgtWppx9M7P2LZpp
wmO2+t4u+/jgvUXkLzag37/h0oZpX/uBIks5GKvtI4gpAT1F0rby3bYwUZbGdGoW
F935v9Wgk2NBSs1jnvoIcrUroY4yMuNG09VHPzMei+cW+yP5H1deYiGY14zVmb73
H+BVN+z5WjNewlA2dDxZWkyocEVh3jMCT4LdljdgfcjX9BfQjceHgspRAQOVZYJp
IGeZucO0XlYO6nbox+Cy21rUVQtOYwszTCjg3EarEcnk7dY+dTtS5aRMC1jUvg9s
KHxAieoAgaehl/XTulFpNv/DhPQE/tXQPIzmIg32sWh8gSyoKiZQEO27vSnSpnuV
STxxeAZtVE6Sny7J8zG1EJ9GzW0+DV28ehr+POzr5/5Q5K3yUsiv9dUUpWT1a4KS
l/e11dQsZElomKWnRDJeRiq0/b90dmjjnNyEn1PvkVsBX6rOQFUKiZNJuKmiouCg
7fe0kdncOlu3Wp9anLrVGfx1VW/MPiulJDu/WTN9/kzTn03g1ke5wpI3HjhGuUHg
3VoEbp0IHkhA+c+kLWphVfe2+Lq6d3pXVvR5ksOFL55tZjjFoCDT4tmHkK53k0Gf
lXM0Jzlym3PrjIP/F96MS2DUqDz5xD4Mk+pzGfGK5gYIh8ovfy5Gp8r6AnKfL9kL
5jhF8VHR9KkLKZlGeWgaYevHLvAvwkPQiqN/SSJCIINOz3jEQ1SXzRiy5xcO4wjO
wNaH+kK28fLYWkCXHHCso/Gk2e/3Xisf2VBbD4HxUQzLFfKM9UY61i6ZrysNzAKW
LtVa9tFM/ixAeuwntlDaYMAf8Mi2Jk7QDDa5Y/0FO/N+v5R7+gwECnwUoDJVBlxC
J3NnwwgeE753Ftbokm+ujgnqIFVHEFd5+L54bTYV2W2KPnkFVAKtqVIx8xji+Q0G
IDRrpSJaWW6nFrvgRvP9144i+xmnYM93RtQ5OlGmhpd5PjQGQiwX/JpnxDKPJlKq
4gZS5TzlpiSSd/q5q5XtN73KxWlm3abcEQnxuLoQQLLaf1dHytfbINt1nWs4OkO6
373rXCCEUOT66zvkZ5CWLDibiZNt4itg6wiwKvmygV6cm2QAIwTKvSvbbEGSeA79
eBY1m3DupzK1l2qm3xT5QMV/cfyekLJcNOtQmwV5eJshgRqhv33p02lUCmKg+oNa
9Q7xxVqFj6w3pE6D9cpjbrJA1FcojG2pBUpNS6DDVWe8WbgDckzw14igUr2V4LfS
XggNdH9ZZKioKqWn0tVgvuvtPOh7qxmb6M8FkQDA5drHez8mfZSjpLB11YM5cWTi
gBGF5jM8nuUW+IUUe1nMcWZ/mUShKA2oPaDLHlgN5y9Vbo4j2H/NXLNVZGFJd6jU
D75FaF4NMAmfR5DGmAURRjaNsZA7H3P3/QFlr7sLNcm3+7dfCnIB/fviDz3QNLJL
YcveUhwaQrFBTN5zweiIxdWO+El4tjxsBpN9t2vR9iyQiykAjhD8GsyzBq37tVzi
zNJtpO0L5NYzErQclv3tC1shMZk//PLz9j9jA0+Bf/V0TOo7ACzXKgTrvPaQg/KH
TGGNxTVtQ6Z3SN9kMAoHisCWZ5z45wtCQlBWyp2oXbkwdSV7TOrIBBu1R5xH8Nh5
z3Sd66O9WWyn4wHEbwJzgFiEe67V729nKmY+lCeTXSUQH4/PJCbmsKpMUeQCXh9k
SH2Whb0GBkfUMoHYZXtAqHWJlRbWQ0PHq7ViGp8n4CROUQoQgLOhlibOFfGYDyJM
xXk2TAluMqvJfh9opqgCcHNuGo36KGrmYUrNnW7ucWgHMs54ZljCyyTVeSyxs7Vt
/qxX2wLJUiaFQkkNFMG01V/5CZsofIANBHKLSY+B3SvFKmqpcHTmGOWBxUNNpbfM
9/XSgU80pUNP/0M2O5uGYZVUAyGD+aAo5qh6ki9JewToi3NgkJ6xSlNU6croc8qU
/VKwDubyHMG2/vtt49jGdSfWcBiPpSwYGQWdNkvOZ3tyIkt62vIKS9t1QzreOJuA
LZREzh+2WYNR6noZtWb4R3mNgKmKN7lzRqm6OV5YmJV4T8WMI+/noIZnwDouU+PG
GMHxsflZR32Bxvlt+r7ZuPcblAv0Hz3PlgOa93bLwAMKP+PNl1UATqgyVgU1QowT
FqkpGfOhga9kd5G6oKcEKYMh+7RbkemZEZ4VSkfbsHGMrxsahOutuspTJKPCJlcl
xo1RPrld66FU3BpStyzSMDoroyL6DYsPlH/UmkWHpcyJ2GC03fBXvmNYf5d6+Boy
3kfHHZ2QAlvmNfDV4Wg4UnKuEjI0/TwmSpQ5wADwwW7+Wc84FZH4mDUO4qfGim/Z
pI7kBmc3TWUkVBSCDh3oLwbuSHLZ/GSDpGg8rcYND01GlhVQf+t7OmtEG9/ny6m3
6MFdJN22AEQBEeNQOP12zGk3vR2dn7jTAowX4QaDYO00jE5hDhsZVAlrwighf7fc
2k/ag1InsvopAQQvUfYo+hP5O/5W8IvZns+2pqFoe+rQ9trgAca2aQBu9jzkw6/H
slLIKE4YNbkpAjDensny4JmYLHAtaZwoqL+ISezrsJhvZyKmnY8IWF/iy6CJIQfY
Sbvum+udxB9z4AShSzHIF1lpRjn7ruwBIP4Rjt83iowGc98nthIWwFaXeC4/DZlk
6JlQ4crzdYhW1vD44sV37JI326GXegwH6vSdlUMHdW/13jgVzhI8vNkdcw6sW48J
CwQrBZ9ZnoE/orqwwkusxJ7G4rfBE0jrS+n83nsjczz1021XOly3HfjPz4csZJpG
Y9/CHQxSZj4O8V+uNizs0IjcgCzsfW/rapPNcSUWPXJUu2zfXyyqdd4Dh9yaq3Fb
sO0dpdk83qfIgyFg0mxFTj8F9dth3LB9FcNTeSDig9ozOgV+Fv2yMN5x+VziQEnJ
1uk+j5qQ1V//lNLqtZE4npLY40EkigRAsOZTzyAgscj/ujdLwjHfLZNJ4TlxB10b
33PQNjtgm59OHG1UA9NmyFOPa2+pSVLy/UYtWUVbHL4/4olO5WjTtl/ZchP9q5D1
DorJYRMjnv1XXI1DFlCJUUIb9FPCxGUmX7T3sD5Iv7X3T8URVN68Hjr62fzWeLZb
BKM71AcPz3rBr1wgob/76QGQeMm82rp8RmNX2Ro6QMW4n/eEhOt6QsEpRUqDLonu
MJtyfaIwmJrkT+J4DuOU2WqAq2IZpx57TwSpXwnl4VPjT9N9fVPrcE3CufobAqzR
rd2hs1xvHc22GE+YZCvuGbnWft5MsfUUGw/y+zm7MBpGUDVdK7zwXfmOTEsz/opS
lvV/gDdqmBGb9OJv9lhN/t/+RWYrgVus6CJ7AFVFrR0LerAMxKL84fHyie9uIQOM
qBrLy90xdKjog9qhGi9ADI+NlQe/YE2icmBFf3zhdL50Szmpsjzi4bnGqPuh+Xh7
L5vTjLOs5FgTTQL4BYM7ORLRdnUjcc/GRmAtRBT/9+Vo5x3kYN6xtaJbwYcd85G7
UdWoD2Vdxo2LgZ78tSRSOCvrr/f0tWmPEOcm88rJMGQp6OGeo5JRRMvs8BtBAYCm
5umXIwCH1TTcmhJQQRmIjPGYOCtVVPQl8+qtdo9zB9iRXwCfxBbOalEwj+lM55uW
CbRKcyM5moi9tgtcyktoEamRRKlj0TfjB1PnkpPk+dPt5aid8+UDOAzkXviru5TH
u+fQ90KA31KyDiHXBV+XGyAbO1+cbixy4c52GTrV6L1Q2nVh1YW1jN9MPxvnmOT4
9Z8gEpr9rn+etsdcJ5GL6kT88/xq8pG3NN5C1GU0AI+zV+ZY8SsCE5Unl4a2W+/z
dQWzC8k8shVmBjBDHj02a6hKhFb60mDdBLVuBa4ilElkvfrY299mKKUlQVYjoudU
X5CSFYqb7tXq4mY+3DkdxZeGeLNl4tVba3zPKp/cryjXz1PjZ02dQj9JePApKfIB
a8qQxHU/to2+/IFD8AkFLM1w9xnSGP02hZ/HZ/6PHKIgm/lhD3iBe1bdz+xoblVc
uaa/ZCrmy6RJk8L64C3bsSzumNSbXiNTj7Y44W3FYVejux520LpksVE1kdHF0mOX
2R7D9VOzTrr76l1dUHI1qe81vo+ZEFNM0R3pgeG+iIRqwphwP8xLBkVadxjpTG8M
uugDiOaapfIjyFv18eIEIqRwyQUuTGVOX4v6Eh4KHOE38K83W5txHEmer/wmvpYK
zayNbKbTlXJstyTGRWx++dCNN7vQ6RtGu1CmYLbysHpe+OC3tN70X3zpSyT1J1kk
trny1DeX0qjlGZugAYxk3bEUjnaZ6acESgSNpK8M5R5UtfRPX7AppRf7t7jDNqnw
KqqaZubBub5sy1o0uR0Hn1NX8+NymDcRz3Y07+oY1Xdlu3TDUu+LjhXCVtMdXLHT
lcdDe0KSULALdtWL5IJ075smwh9bbIixY8otf9puw8FG2ajxHMi/+1ag/miIzxyo
HiTBBaA2QaulIxvLi2IbyfpIBoppK7cmuB+yZI8a103xW2SUT78o45mGVsnDgfHX
2APYw6FfWtopCCBMBdLc7ZyLozvlcdgwT6fJejoQ6EcKWRTdw1vvjnLKO0IXD0sZ
IIgbFh32TKTG7OCwY5uo9sdp1c7qBetAYMUT+jPdv904Coc4g7crRh6nDlEtaLG1
Gamtzsj2ujjEasPc1HQj9GbnDsSVEMaFDQd4xkQV/Tvs/hsEdA3rSjwMQOTG+NaH
+y2ko/X6Tj+XMpCJguAH/T/ZUIG9gzqYAR5lIqYB0Z1KV5RzPrRKrRRxriEVESmK
8/uOacNfY62D2tqk7VjC6sNe3ZMWsKi7aZkgXAwpvbmbVTY+Bzss4IZZqmpFSI0B
L4db/tX7ZIlT+B6ZGAA04jXAHlxP+xBAUfBFjXppWvUY+8Bg/s/sFx12yeYLF/cy
2ZiPVFYxlbZBo7uy/4QC3GAClin1gAhlbrkUrv/17FDQ+A7ccbTHH3b+CFx+vCGN
UL50UaQSlRqvSIKEdoKQV8PP+cyz0hMKXPfzbDs/utH0Kn/lCoGXMzD/5kkjLyzc
+lEkApZrI62H+AxiI0NwGID8HL8/hdRcz2cMnI1Nmt3JpRdzypXkY9CrjWPUamAd
SnnSh52Ikw6EzxY/v8kxZ0rbzPclBeo6DcpaPFm8Gdr1EhtlSM1jcTPWAVuEbUwG
lKrYJ+NUAwlk4GXK6uOUQYlytapjR+PpP3LoQfdOPos59flpm1b2QzHsrr0RR7v1
LJJ7p8vU0MXvW1G1qvWmbgJgkTPqSelaeVLza8A8LHbnsc2iSSC8xw0EqaBeQws8
mE03TKn884SSGntQyLxlfsCnKrdSxrTZZKwIukSK9T1LSF6w1xIEnjMDn8YwtFxJ
zTXRnpxt9+y54TrDY6Xala4kEguUWY2aO3pIEL0O1CU+QfFToSF1danqPRdQemtH
nW2u3gR+NSnkzvPU+NjAj74/fi955/533mQWxLdApL6TNqXoTruUiMkKPJ7nIclE
B+EoPeR2yvdrPRzcDzLTZ8ujmBlmHB3q7RczOnQcjKowZqmHPbpRlKd/ICbDTP0K
k/dzygt09wEw06j1sliCKa9ZnRrn0ZMBWDk+psa40AN+KaVBOBK7fbzTvNKhjiEO
nR1cP2/U2bnO2IgPYPnwgEvnjLv/MfncrOyZoKOTaL+2yralvkyCykYhicBdXSKK
KBZcZqp53j46rZQ3S5iSyjSMGdkdZABY18LJDMeNFDxlo2AgbX4rU0A4jlrPspuI
VD9LNQaOL5clEkQ3HhLUJQOeeTw3P3SGxKWEzQ8JgL3F9ji6OVX6wdtXcCeD5Waf
0UNhCbIIlixqOBLSbbP14R3/EhE4YrBQFOfVV52lgGWmxNwi+qmphidBYKWlk3wH
76LdCapB4E07mooGTWrZvTiNnivGwpe0PLVALc0qvILPCx48mIyi7mYsX8FkDYQo
2eR8naeA0oaps1AZnMkTghnSgbWW1/z5Z0jIkptjTccNtiXHzpSc5Jop6mVkXefC
9saA9ucs5yCWgRCAXWJf19SPxXYE6DO6A/Am1+n78ydtp0SRyZd+me5I7ZS+vlkY
6RKNjofbm7rLHgfaPM6G1mnGhJbBtiRLfCjB3vB1DVx40bRFbXmiqonwsZEF/WRT
+jfqi42n5BfoZ6I3WUWce3EOD6jD4wyj/V8zBPQ2Y+rT48uCFnftqyvH+j7n7Jyt
dQGD8bcdrMyGsmhSyrxUvZjzL3NHszY2OkS1FmYzbB78DnEQg7OyU7F2SwnTPvp/
LNWn/8HfrfgLTynE1D81MSU/J7jw4K+2/zTgA83wKW/hqbAHxeGHSBcjZ/rYS00y
1m2lbg/vNVrPSGZcaGxlUqRqN9QUwF+gqWaI8tQkesAo7S5tktmbCRP2IBgCz/sq
w3TctyAn42UceaLQHzs5Kt27cfcf9SR85wq20xOQxaZpP9Ke9v58Ulyy4djKxRuD
hSPsZEGOouse+I2FoLSlpk51QQnlrGSPVl+lsxkPJuimrALjzIGARhqIa84IQBDU
oEcto9To+p8PijCdu5iaDIXnqWAXp4N/tCVNsgB7HD7Ojz3Udu39hBCzj0qv/LBA
6+OnOJ5sD8baYGxB5CWYzhmvBQqFJtT3tK4lMKk7tklr0+zMbybxoFFRgT5PgsFO
0fMpFuqQF0tWzXOBpkJNoNlZnPZejDR8rU+tm93up7NDKpmpl7prIUUjmmwd3ZAi
TxIQyWsdAx5Od4fD1K7k61Lk8BT5V2M07VW9IU2zlw72E3VLgkd8v+klRZlzDpAK
ISURWj+Cy3/3ozUw3/zAbkIXg8xxAgHtxXpKTeQpUbJAGx382Uon9TXsHdY4LN04
xOy1hih01Z2n4B8zxR7rprUGrA4i8YFM6pKZB2kDY631OYAwy2EyyBvswjtv0fQf
8nXw9KgvFcNOINCCg2dZQz5sOdMsOCtTTOyFkWGU1MeX3gI0Vfcmg+dp4SqLJG+E
PsXOYpDy6VazCl/FEIhD5HhufaJCKg/s8L2nI9iBvPcHFVqlA16k8PFkjDtLyF5T
caqk1ETadRuvF/93Zf4yBT1mSgMittd0757Kn/rpfm6/BWQ/k3hoRgqMFDxNsytZ
SQeVT2KG1QnzfJIecqEGhcYpSENOPyAiccuV4zAiR4sVKyH1uXUzGXlhF3YFxc5e
rMSYOQoz55UDa8Gg9rFE/0FrG1OS8d99cSuCKToQRlbSQHvirNrOfue8Pl4xWKfV
kM7WaAe7VHnuPgQY87wvZ9ZUZ50fdBshKtKaa+85/JCgQPIo+CcYSoT3vxi+asK7
tCwqoADnJ5oRN4JcRyQJ62MG/rPQn8Vc/DTavazc2yEBUwoQZ50y1Pki+5pBfQdT
AvovTaBI0FKIkbv6u8mbuGV7sS4hNvNLf6Tqf1o5RmxehWteMIBKb6smaFfzXm/X
Gt2SWwObLUV8teEgMywm7IVnzHreCo7+FUIX/CVQzGofi9zwygb0F64nfJnduFgr
RieTxVAGM4OW4o96oFySB9gVXA7wobwLwF/He/6VIvoEpWLwAl1I6Ax0MLj/9Nh6
eNXrpelEvLlmMl/8PaB3LTLPLvfohgpC46JkJkx1CN94hOcXVI3sNRAD+HvyVxd0
RRm/7jpXERc+WK4/tM458Q2ngjCHW0Nt6/9gRrpEWYqdueh9Mwvw2C1RP/s/RIPn
RsEx0Lxu3k7h5YXrOzU1CHE3hGfZdmMaFlj9JLS1Rny2XvvECxBy1nFwDS+OqcCg
XhuK0C1afvzCQPEUUjreITapi8jPFYOuH6CvuM67KBJhhG6I0Ai95v4ZtGUMjZRr
btQr2LGKT1kYPCDlWQk0o7Fbm5Vtx6u9VBhao8L+/xgZOdiF8xGF8KQ/QJPkYw1e
N34SkcTvnUDfrVHaqHL2e+25cA/+LNIgU6aHR/kW9BgQO8CyaWOUambMKvivwsif
zJuAI21+Wuu6xwnHFd4jUTQiXqKXrCjndnvA7rp9tKcwqeDnYp2mGrAPfRNR2/g2
IXqpCL2DOftkJ2AZuFrEDSI9+QcB2YVyyX9W3zd3LmE4WB0VcOZNwVJJPgeOx5jk
2PWE7QTFcKsAdwWbECrvjl4noiV78oIwBVRrteRh+AQfCbW9vJgW9jPnjtCnDXIz
6T+ha4j7X7DCPqYzxvw9Z5dNOW988OYl63w0cWXrdHXbocRPDm8T77vnyio0LrDn
/s4mzyLlH3Atyh1shj1K2YqLPGrUkUl4QJEyYIIfeD2wotjmKcaTWKbYoYTHJ4mC
Jtr4JvP9VWg+gxu13Kv/rbqSKI/cFzwOMDTnfydplBIx6jMFbCA2KzmrH/kzn6VP
hQl2pAuUkiaLy6S12TrVfOCBs7sak6JijYHerETrTstaeXtkfcvBJt/9h4iS8Mh4
05sxUhd29BFLC8A7dEIY2gnYONBLhsDtD2IzdG+SwUh0JTQXNkefADXgpqgxSldg
P9rgqK+GalezRkuWSw3oKBJbO1VbN3NhpxQGyKBKE6OkZmofFA0qbOG/TcdgUr25
Z9zBDT4Skqu1GKUa38Q72jQaOKEWmChpuKfQlFwAqF+CDTF2kCV2v4KtxLoP+lQt
5VWHFZh6MMfXz9mJaE6ONro5hxXEUHHE/5JFtkzMaIOZVuYCGkdHiLqGlinpyMt3
VYXca8AqG5/AEhfiwe+l7wVPU3Eoa9FIOOT1IEDui8yqKmUwMlPw6HY0eeYpF/ZE
XJDJp45Xt36faeXejOWiIX9IrQkMBgM2pQNpJX7qvlYvkIApS002TGaP876eUY58
y6G4h5zgFE+nNW8AxQbbBg8f4t7Wm9xYXfjwbhRw+V2rK85MNwcN/q9oPHJCStQR
/iK2jYt6Mx/qv0YqXbzKDJcQvwJ4tMPoSFKYt1zJ1m8XGiBNUBmOWLLHthI5of5i
I8xPxYSr9BTvGQnGBRRpkgFDegohhIlXJ9LmgvH4J27Bu3E8lnW1fBxBEelrlvAj
APQh1IUCkzXbE+E/yt1w/4TlwM1bznvjC/S40h4uGlNhS/Jmj9fz2+86wTShCThY
cxrjW5V3HY+jzJESNPnqAkJXsJN8bBObEq5nvoOZb83931fvykOZTbDrwUMT2Ta/
6yfsc78HLPC9134wM4dnhD/Nj3yVNbInK1CV83rjUnHUbMxpZZOptJcVsgTFF66y
x4TUeaH5x0umBmCCciERm5CaukDdPU/bCbMB+SiPDV8QRsvgKxWCXt/ujtQHGp5S
jaPFDPC33bauYjI1YCc3uPLPtDdssn8/N1ygbqOmbW9pO5puHRTxKa/+bdYYOYEg
oNPDnbDid/VGywNu8876UaFGYvBpmREfArpgBkIeZrrUZztp1zRGgWFDV7mLUp+K
a5j9YWWOVRKX+a8jXq3NElJQnkBJ82v+dv7INM+TGIyMctzQ8MOKLuxNB5hkaRbv
snAOqm4C9+oWgTcHQ0//YdBOJJ8GMEg+Gx7TzUg/K6xy0xCmIPGAZfXfSjr+U3yr
WMYQU7ySvv+QOdbI21fEDeIGvtKvY/+QaAH0aElcCbGyJ4o8VXWjbJXjpPdymEPp
lznksCIjvrmsBbHO37DVwR12+25czM9N3YJeFfxt+tVpCh8KwXCCQGGfgR9v3N/A
CV/VNbLqR3JsjBDyz35xIeTbOJYPD/OEScan0fHqZQ/FfdA+u6TZIFsOSn0C+/S9
L8OSok32LI/q5AhdmrrAldfWsGJRGLWmyTgHzL/4Ufe9cE1XzQcyelg08W1EluSy
s/KgEGmekR1Bq1Oi7uFrGHCILtoU4rfcRuZoRNmfhINaMKrCx/vXR4SfWvqKnYAq
p6QejY53+2cb+DbgCY17oYJhO9JsH7x7IGFTBtKuLyfVtV2ole5Cy3ZaVDFQ/oFa
ASs+5lk1rw/Izftn/miHk9LcqYjDTKj6UZWeSr5akqGxnSGxWc1RUj9tMSBhvWmt
G8V8u2BsjG4HFg2N68UjVvW3jLrlYSfouMNKQebMG33PPEjKrrkMDkrqdKESfygE
z9+xrS4daeCkRTi8M49WIl9B5608HybiOjfroHSTcGAiXFm99h6LGxTyhlIZTk2A
aTMqtMBIR+0rd0xh+FdVcTtwoPuslfNtREXP4K+17ZuzOyNXCR8t/rdhHMo9UuoL
XRhz0zMMbeaXnX+/iLDujEtHVl3b8KKtVXZple8tT1U6suCCltjhy7iP4n/Lnvpo
t3RZ6o/lzxAXqwwFJAjIyh5NYBOZS5khSuT0HwC01MWnmaaJ4SmSM5Ytyg8zVfkF
DL7vKtcpyidavgjVBTAJlalLSn4oXoFdNyeGDuIDLAu4bGxf0rTpcs9Vo5RryUXF
RYYR0lcpovqy6BzH85W4wSypJWMK7jtCUNxHdP+ZJVhbnyS5SpM9NGYGby6p5eAG
36jEQEy3Ck15knvC4gZ957OuJWzAb3GAbATmadpuQ9oUqIUv9Mg7WUmLN+KNjleC
ak74/aPhgSzofn+o6j13Sj4P9Pr3zw0Y0rfO5oHCESSlEHX8Cqbyg641q5lGUd1H
IZQp1ed9WUxiTJE5B4q5tkecYb6IjUHVZQSp2lGPbKbjFlKF0adEOFbPOelxfrLX
3pTqJKvywMF3epK35HnHkU8Hjv+EKClKYFlTYLpakhOKYGiw7t5C9qwJLbwo4Ehn
QTzjzUGNUAwWZ1yMMv/W6Ha0rZVh8uYpRffw1feeU9wWWeIB/jR218zaJxnzgr4Q
OtjBQa/q4QhibX+M3vQkLSvB4dlfykiy8eQH/KvzvaKHbO4FWJEeVMnfzqdXGx15
uO7jzHv5gPxi6+W7mjqlw0X+yJ9wdQ9NYDNlTnuS2FLkc5J1UbM2/FZFXJ5SZP9I
PILtJ8oDC6DTeFgdSQl7iJTTjbH8+a7V4HGAgIylbU+HjfLcSZeML3EwpPdTOhYi
GSg2naRMQGsoTdBqNyDTAtDJMsvJcPhbkB1go7aqjQCE4zsc8E8ZRK65CTd044F1
PhR7Ca9PO8D/t0rxSBsaaXlzpQ78QE+sBw6fQCm3TunmxzHiI5yCellYBUVPzdPr
mFU+VmCx4nuFhVn/FTDNAA8OJoZ2nfued/3/FndgI6Pyx0QF/QK++qYK1a5FiMbH
UvDQJvSuytrabn2dURw1bf3ePuum+F463Uh4Nreq+7qbpvo1Km+Jp/UyIp9ulWSX
CsjKEDE1ELSvKrAl9uRlAwPukqg8FgDOavBRtHHzcl1jJHQox8x/xklEeh9IGalu
QjWudaTiT5rwWR/eHfvVBDUerNkaYqpTWxaxobNma/XdtLgfNyk7vTN+08QjgDwb
sQq5i5+ssdB6j0X0NVJK5AU3TgTNI6jPS9qJTUA/CvglydVJqZLSWbuwaA3z9Q1G
lOfecc6R8lttrjHHU0JP9M4ocb3tm2A+OOQoKQdgUdiB4yEhTn+1BnvrtBl9BfL4
73Ul0RPGejiWZSdwANMJxK3EvCzSCStWQC7GiN3YYEQ4doO1rYMST/ZPVO4hz8s1
22wjj2QxD0xDgcX/gH2whp3m9rqhHZ8TSZtLhWXDgqp/c7KMSfXJhF7NtVuippOq
1lo9HAVDuGU1mnGS9jHocpTm5NKE+2r65q0ymv/LyQoAimgnw4J2ieOgmdZe7M47
HZ0KRvt0FZP1xkXdPaBQcm78dgQcsuyIY6L+pzZm0vAFo5qce9qjoyfOZ8omLw4H
LakYA1DIuZh4SwtrFPCVwLWyx99p2qmf1mgh4oh8athVMHtOci2tJfkztZ3bqqcR
0XwQarQSfPNzYI8C73LUTxo3DCWAp+kgJDlvHUAQuImiUHCBm3r/4qOXO1gfFJYi
3W5hr2uDJ2F16KXlZk3TIRhQ1NZ75nkxNiQixXzsAhwSUiXjmfUPn89iX9P4EN47
CggK4nBL2m9XncWpfyoKntddUY3f9PC3WhFyZ8EjbrVSiq1p6Z2AiWauRuh0Vil6
uoXjh8YHPSNWZ7EyrJLwP6uJX16qEbQZmLbsvVk4DbfCzpzroQExdBfcoa3oR3aI
3WzYrr6Z1lC2ibEQLaI7BC9A41zxQ0H/iJNFm/lV7hFKwuvpfITn5SX5MnvNAL6Y
JhA1vjdJCbnseA0Nzq7rpqFaotwiycmwHWh4RtQbL/N9G3Rxp+US0yzFyFkBO2o2
r0l5JO7MTY6UVWAzJESCtXve5O9a87lOV5/jM9qTxaay4VA6y1XOFXnL0w9Ldft1
+F1+Suvz37C5wBYTyAT5iJcrdfiVy1q1xW8lmoWw+VEUTGfOdM1fzudUPibQ5aUG
9rkGUzO0bmu9INcFK2H5tVeon7S761Kxy6k0XSftncsAaXqdgNWRqwiDyEzuxxcc
DwqHjoE69cJuZVPkk6yfIkZNF+FdJGzoFJG2yytsMvdxGR5kOD8hEteDmTgwxJ2J
09yblmYDS4KkrIuc49jaLAZmLdAq4LfL/6/sLI8pD+ZWcpaxrtqbPaxy6SJg02Iz
rPCgbo99tLO4ObFfA3C8ujTe1GpMFrPbWUDKaZNhr8EXlC4vDnb2H6hySQVBwhqN
mi3PvjFS/dAiJQ6GRvHHQ3y58mL2GsF06tbKN72PAu7Bmg/YQJM9zZb3ZGLtEit4
qmuALUlrr/hxnjTNWR7aTSHylYRWSIC01l3KkqliN4Ix5rxSA64LVa4wTveYe9Jj
mAzWY0CizVuO3SUr9r5ozgvbRGaLaMqW96DnG7ptN/OQaJdUeJBdP0SLJCca8tvu
SLG/8ZCcUQWbDVekiowoQjZH8IBESiK2aXh8Q6g6q5hD6Usso1G1XYsSfvaMy5Td
62XCRwRH5WqeIgz9w7fUQ3B7dIRBt+zj6VjQ573lD0f6P3M0k3+i8OH89/S7mc+k
WZctHc3ewoKQ+cCu7iUJkhkPy5u3AeR1RInaaX5Qg1sHzbeCwnPVjK0Yj8ZYF3rb
ua96ATlEE/Yt0msWOx1qXwXqEkjVzVNaE/t/yvI0UyoDWX+WuJNM0YaRjtV/Y53B
qXHN+or0LU+0s83bz+k3Tz7LdZ1fM5ta/8pII9j2HydS68q4qTVdEft4BTR54GWg
YndLRLesTVqokGbLGXaOwlok6IFbacNN84FSmNUkPcv3G88Yp7L8qh6CIZ2AsSDY
kN4eISmS9xFDJojWGtQiJqpmnhzz+l98CEL5BoLWaobh9e/LUpNTAt3jwZZGhnuD
vaDTCZEXvpJJrVjieDoa/Fk5z6E0MkSeh+GMPVD7rm8GQtW7qYwtfWZT3ej2KUJR
fuh4VIv3KNKa39La9wn++51m9fJbL1MFXlHqjVdzLsSjdhJUcKASmYNFXV1fl2z7
eSdeBqR60yP/r7cacugsaZRgDdXFgcn4xr/avF2gI5YsfL/AvIgwdQ5l14c/g5oR
o3OtmjVyJX/C0gC8ofvaTsGPWzweyy92TbUY8kGQCljRGXFnCcZy4xvRKjDqzJt3
McbaMuntXu7N8CqOLFMq4mKQ56armtbK3LF2kIfzZj/xJMsO8gRZORDNA4SmW66P
5cBJ5bg1giwhnfc6AX6w6916xoSBgk+c23ZTUk2D8paIMmt/VvF/jjVOgye5PBoQ
r1iIeoH136rRmxKe65hwO15yjSPquZviz80sFY56ZfWY+v9tIQ2p4iw2kxx/HF+q
l5QHKv2G1phVCfgADDESjRmy7a9xFA5Yx49KNJ1GKCA9b2T6lFrX9b9eqib9fH3h
QANyVsDJWzq/7wMci2hIdEJ9iOYiSnaTQq0E5W7LeBoPgwInaJkB8iT1py/UxqUx
idACjEc9CJ5l0vRc5abjbxyuuSTG+8GINCpwGXxpeWrRNoCAGODxv3dGTB8XDnYt
ZvDfYUTrRkEjjFttzOsbbCPWP6OHkyM6grAK1r+NKcPjdQPhZZc55B2zsr/HK/ap
h5V9k4k7Tz9U1ZQAcYZDabL9XSPFjzHjNyOx4kYZv7JzB7YSShlmT1/8YvYp7vJt
WF0b+l/BPvTvtkqCG0laI9/bmkOOzuc86/XRN4uCAIPl6+Ep28a27Ignn0Q5uMdl
lm9obpcRVIc9KuRGT774H1ZkPVjSRo6V/3znDE2PjN+cLV4zaQitqw5LAWePUU3T
UhZjh23nzBdFghgRBOfhgWpvjRDzl+nKWTitYQeD1e6e7IdXC3HRd+IQscTZc46i
ht4mu0WreKz3/VEjCWW/m2i4ECdt4CRA8izXTY1MEVRH6TYPkrSpQc23gI7P/ow/
kTD46gbH9BUuDISbpAhwDnbW+L9lcrq2G/Ekte5iGIi8AIXa4QjkYGu5nG44Mwyx
oLb2H+tcgZ8c4shbUUUYX6KePRZJlTjQmF6MP933VBVcS7PJ4Z/EyAXPN3uF2gKi
So8l4Wj6pG8QVV3mRgzDCtD/tLS53b/z+MBdJZJriazlj1KSlPVDz7Mn9iT+BilJ
vOYEnuGxzXfyIxJWD7VIr8Q84JqfQiyoPn11a+7rzTWil/cNpbA00w6g9+XBJs0a
f2THte24XtcQ4Sl2VR9Thw8zRNwzar51DZIegzXlZf1Vy4xVouE4ByWpgPLfsTmj
j+zqWza4sy8MGwpgLG1q51/BVOeLqdtqRceUR0mMGgKFjgW6K2hUDa1mKM1Nw+8Q
rpcwe4brVdPkcEUFPGPmUk9+ShCGAnuWYZnPJhf0cDhD8+8xMa7Sk8sMTn6bdLT6
P/394HKjddeXy3Lirlj1wT78RlyYKSPcF2iNdITmPv+fysIkQe+E1ehV4fYA7+M/
vHeFj9ht9L5O1G9MZFrI/HU29hp3W/nTo5nZc/MLatMMXgkcJfXdmBFyvSxjlYt7
cWImD+bhK4X82wxP2WaSTFUV3u33rHJRWRrxXjeEVwrVvgb6wf2sCKU05g7fVdOR
/DZ4M02AmSnniXk04T/Y0xxdq1V92ZC0exPMfQdNzx81Cc/CdtLeUWrvJapeTwmh
po2NAlGBe+sJI3dOIQuMJNJfnV4eAswCxSGfqPLuYnXlLdLyYmhIyLGVAtdQ2Cxa
ltAv0AhYHhdLB9PhaL3w0XniCW5EDf0iRja7aNOf3xV6Qu5edz+KZCM/oMQT3j+R
fY5rKxrKQ0qLM2CiQnY0av9qLvCuY8oS4VWZf/y6bva6//SdukdiieGiWmYLEuW9
1WVqod0CPxlfySVQFqw4UNGRXIOTra2UNbvDyV07KGPwEiFKueBMMVkmj86Mr8Lh
MXZikXYLwrnn7MUVhs+IYqRb02nFzsNi2rekjcYKgGY73LWRP+PcRmDGGJsyysir
WrsR2oLG6hnV3MKKiwtt06DRetGvDf3ijtFZcVLgzMTbGXexHBuNwHMv+IpyDW5/
ctHRYM65LQKiTkUP5dtiwuSgfLcjXcwMHOxBtvxWpJNAQjoPAiG14/iBmiBIKNFO
SSH2qxjZnZzxJdjqFwHxtN55HauwhkyqLylLpPEhaDes/cz14WdGzbmqs/xcbngV
Z9hafD6/tlllkp6zcV3bcC7OkDG705OjofSQ52x8fNpsaJC6brIXKZwM9lkpPhrE
YqhDqXRjXGrPMiNPsHC9kPFVdyv2Semcv1uvB0UFLZzsRqrKh5BVnAyErjRKTUVP
yyL1xpzb4JTPY7kVc10nsetw/+w9mNVQWruPbnyv0B33DfQa4xWeFbSM0m/MfQ85
urVSxQSBpHyat67ce+lTpE3dfdsFey6iRy4vK4TpucQtWJcTJli8RusWZglVEO0w
/MWLSOkqizHMbmyJQACxpVIRFggH5+k/zzASDocfvggf1imibM6ovopjYTdBE/PK
ECY3lwsARZYbTpzJmjexCovNAoxa1bXD7PSSolzp7GWBkQeMa/HyVQe4eTuY3GDb
u9usjme5JIgUwNdpHIEpj9cu4TkPjcdpdbIOivGZ2c6fr6h1Pc5hY7oQAUPBqxTl
1VGv9XC4vylj8dCd7iwWkDLgOSvR3caohE7PWrCOxe6J5KTDhGHJBoZ7LPSrcCl0
IYEL6ExLRQG7yYWdjetrmXxh0KbuQNUTBc5aEkdHTgL5xpX7kfizdyhec8BFZgok
qiW0raq4F0yxwJg7Fi+bxBC8F4F4Cz3DaRBMXv51UfOoTiAYfnRnvxMPhKGHz7GM
+utydpbSii3seGUS2UUh4LCDRw+EAPYmQ9f25ELbBgo+9KkDHjqCmde26q7UV7f1
JqzHB0MFB6EMpBi49lvG5QsKQFn5E7e5Y6NvcpZIXXT07g6i5yhEKN93IfdrnbsR
l2lEQY14tz7+GtBS5Lg2cQGtmexhrR+I4dYu4TCHsN5sNphgAw7w/0hIvOdq8itS
R4dxhrrheIcw/mypdTo1MCVI1nbDKFB+q15KHISqKIZGf8MvUJkyqWySieXeBZtp
M+QAPVRhERFJROcclhQkbWNbZIGIIqTYPn8SL1mDJIH3bIaF7CENExBWMFRo2m97
9s4lq5eiZHTP3Yu6Rpa/IMR8lK7eTntOtFNn6RqFVPva3o+YvZJT30fhOGuQ85Ve
4c8XRb3439Dxuy1Gx8Tz6rgmLw7ud0ft+B45eORgzD5j2NfqVr2XCitF3pIBfF/U
Izrnp/M6u3haWNgHr2fmkcpeDunV+EW2w1JWwfwE25Eq1u7jF9H0+eAbhOJM6fEK
htW3bHDAwfUXHXqrDt+AmLldowLvl1qqU59/vXaIv59UqXdviSaS3DpJlpOe4XaU
A7SdchH/0KR7NduSvrSNCR+J0bdEJxMj0OrsRwCnGS1OpO9SlwZsfaTS03SXlAso
R3dZCaCFy4DuHTMWwN9D4i2pDKD9Za/rftuc7mNjExZMDXzTSAxM21yQ+M+54q/5
n2HIuFwIN1JGDT0Ekcgx7wi7e/e9KbLHBuUi2mXTBqCkk9k3PU6ZADGkG8q86Rx+
k9uy0iiRkkLxyhO0vId4hoRiM6zlFWL+P0P0/ozn+nTdCHHmb5c4wn3YuR2WPxv8
usZ3FeGP37YEcEZovG/CnWdOViJOEKePVFbdwQdI5+K7hNJ5AvSiDiuDx0fgvhL+
wDRJ34kkf4Gv6X07aORI8/cgGCZsemeNjYKJODOVFCoXKC5JOMjWYluSDoRsI6hq
FBSMUo8Pt/vS9uyraA1Dt8zQgyV/yO47Q66Kz1QhfDvOyF4sAySoGq8nMa7Jiyuj
yfFl4b287Gu5KolO6Ms3Z091pMA0t3yferFQ229yU7fOsIqEVwOR68wPylc+lkWa
CfB/hvZutEJsNmW7ks/7RsU1+tgrOr/lEaMPK3vSQyoo3uMaH2TtDRkzpgSF/xuG
Zq15xnDpzl7XpKjOxDO5S3vpsnVM8g5GOP0FLfP49VDwzsWrzKYWo42mDvQNCtTA
65lP8ilWtCSArQ9MI2L/r4ut4CQmisfz5ORowIC70croyLyFAOplIjiN4Qoupyt+
05q2V5fTQr56rGJyTU1NcxOfibkMKqMpMqd1euGKAbkUvR3CVNtqG888h6MJE7EK
py4lRxSH5NnEc7MdY+SemB19oErpj+m4Az6UAIkInw7YgpfvecW3ze4uppoFlzUx
m02NcocJSPebqCZTxwGy1gcd+MOlIgKB72k+Tr/EjWOQTtbuuizk1cdvh0CLxbol
k/lEY/AO16LgeDgmKkiFfTFs6y8hGK0KG8SxqgJsZR871n6UmtNFvhjxB+o+sT6R
Wt1wokMf5Kqw4Rne3wqTfiAMlGfBMI2H4fr9jjYmolIJqD5qVeYbcp+7VSK77Bub
ejPr3lNhGg0t25O5DnXvGzhfUfXq40ZRbeIe5ZzVqKeqlaHePxhRw76ZbZQcLB2u
S4RTD2oP+Nscez27Wy3VihPnTUZUDxWUSFD/jMU2vDRi1AV2bh50eF7203eGvjcm
Ieyp+AFgCZaxsjxIdGhW0sYtIhWuQoGLRmInAUtCsiyywG3T5tHia8Zt+GHdwiCT
UjhS56QcWtkyjb3FqRlWCrW2pOtM5i+ueMZTa7VV5AUeMcekNQoQW/T2affLK2Ea
mYE4IHvlH6zQGPZ5Cpacz0vEvcR17a1VTA4faHFU47FzTzWiwzLmIjKj6ccfLcyu
fJSN7Ua86hLEcywltbvFmSxQT+QHLQFNwUAf5dHgsRP7VAFOkNDRexkjJdn7tYBK
3qskBk/LfvAhp1PS5R+TI6rXcodFt0Q76SLowZgADLiGla5ypMDTkeDD6aQB0DXV
UkWB1+PgnfddnK/bLCtQL2UHu3Zo6AhoDWPmN4FFLs+9fiBoxmgaLFwrYiFVzixn
SUTN3eTwqEAmLdya4jeOfiSgMh/qY5f3PlvvqEK6x9gqLYLJyDl9qSXblNaEStRX
Lma7XsoKKYsMhvK0r62GFhnB+x6GrRAgdITrR6qBATgcNLjzMIHF3FHgy7/cmYzr
jpHc4HYIo3PCRP0TCsKFKfeFjSGRWfyHLnA09wlGEHLq0EPzpqAUPTWBGdzpgTF9
Jn3BQTA++nqkXLAXZuw07nOXVoTPQj/i8PBhe1PXzWKUxzGVChLiVqqSSA0EQvsq
+giIaCmwSh/+pGHKUJJuhfJQP1w708CoIGhik3iOIKzXlrlbV8duvGmova4txG93
qMzmiUdDc4yOysuU2+QPiAOSgaqnWY0t8Gcw47oIlqkH5CIjXz0Xo1T6pidgsnBe
dOk+N1aTp9lWxO8Mf4s4tSw7AWaH5QmwXwv9x0YZjOH05Q3Vy0xd0tzO8HsmtcQx
V3mE7x8Q9z3+SbeB1GdG1adH+OeV3fSKiNs6gBM/k9xyqDdg7vY5jNCcwFtKAtMD
F6DzriDHCfliF3tZjh3FxC/sEawZ/RjHn6u5YGen/J5UTKjNKr3OY+13V9uM/Q0b
v3TUb68X0+7HBRwDi/XQLBJpDwPyZ2AQ39gQTx4hV3sQRcmxCR2na4vWDfjtkm9P
zj/UXgxi8KM9UUQAo+N3hOqW5ILKfRHASC/EazTlUMpQqsp53Ev7g3kIhHe98LG+
h4kKU0uCWUopG0KtcJrgw5WBAWtyPtWrSWJzRuJnjofDJgmzHuJhn47UH6E5Mm03
hJfwAUIRayhfCT5Vj+06YvHFUqzTU8sS74RydFysoQmvDs5IcdkrRhzcJHM1rlAZ
8iufBvcO5FrPoK+Ar8e16lNuMyAIIeF+mkQtxTzroDzThHpcsz9eyvdDjtILihi3
fqB4x+SRxMmnVM58mhFGW6kzLEY108lRxS2ci2hT+VCjLFJc4nZlDrZ5ixLR/QlK
ztCGwzhe8Ywbc5ESqb+P2/ggdmOhksUchqbcQeYRYiFl+Y+/8YoM3WE8Ae7OnMGB
+ER0odXFW7Ba05+YygE5FRdolJLW0j7tC9DOZrRq6WjFiITPSG+/a7L2N46XBmzI
9PVzZeuw/0zv5MwK5l7eiYYcW9zC1GwJ5pdgPv8NL7Q8FqtXbLl+ug28JqByDVmH
7uxw1zWiD+Y+WdS9eDBRuUtAB0y8gfDz/KbO7Iw3JSWLKtpKQ4yWcONEUHEAVJqb
9wi6KMdqD9AjZUIcwPdzFmaQ2LffdldcN+HuvTviXXVewB58HpdM51Oe1xaV3ZsN
utnJzRs7M2OgGujLan/JQTJfX4FjSf1mccFETl80Jl7urQvAesS65OJnH8iAaw2s
OhCVXbf9WdEbvltdw82KSc8StmJXw5Q1qMechSklOhV2/zAJyXZjGzvPu0w2RJtQ
jhzfBdEgdPbooAJq6CaF1nWp2VngARQaxl+ZUXJvB1Td/x5WXgukNiaKcACphUT7
jJ421r9fBnIPbpMAjyWodpvw+EUJtvG61XiS2H5o/8wGColifgpZHUsy/L0Asxb5
/7Z6FBqLwTdSp9A07krvgtCaZXGsOFBVXlPOPrkhWWeVhwvZzSrMwoovuKJS29Bl
YUBYxIrWp1R4A0XRUetZZR1tLAGwqWnDWMysU/Qr7IdIaFNayckzv9qxi/5tQ8Gm
CJF7xyFaz/trgZQ4TgP948FVn6OZHk+F6vg0pGI58vp8XtkN6T6CY1pN09/qyR5q
U8Jal1l8JBPF4ttJNlh59hc+cXk2GheGwbuSMMSsInVkY3eXXjA8qIWsh0T/h2zz
KYxQLXCXulLpdZQh5Wu9pzkN/nBXFMHpUX/jmvzAGPEvUlZHypySwZk8AeTbi5IY
v16r786iQbzHSDAk2QNCxlKPS4XwU7MRvoyTjzmoSld7epm/9kS9lyYxYz7iiT3H
r5EUk0BT5sKTRChlTs+B4hGccXnTa+67XSR1Vc8L4WnuoAxbJJirxNlNRMTKlpwP
X8KTxkXp6Xlekqhfo02FEMFPLhA1JOgRuk2ZAsM1fohhumQYWigZIHpvow0nz4m4
L+3STm67g9SbjdVMpK3xgV3ExxNh1ilEUYjXbzbnI0CXcdo06IRpYbN6Mc7OBbz5
iJqchQrFytR7leSKPrLQU6cwJpI8uEcGRe+QWtS66xck6Y2dqAT2dgJqu7wruu+/
6IrWuCpwL+WrexdHMF3co07yr9599lmdGj/vb2N+kPxhCjwEvGpeBje+h3zaS5at
st7e7nKMszM+HmguxRyKEBgX07hkQ4YPmAEcMP+bCoi5unHQ0M9mXdwf9N4HgDtV
CFChcNxt9FsCBNbvXaLlt1m+wNBdH1039w3BKPAg3Un4UjIRw2xskQ5N7u8lWc3s
h59mRNT1Zda9Z/pccQVQwpF8kvW+TyYOBjaM3nm29YmCnvMkWU2zCE7SrSB4j6Sx
hHjIMGgylAQY1cE8HmRB1R+PnGf8H971fHpQxShAxXD05CgeTYEAgsRqWYd2+464
Y6WqwSjTKkUdw0yoPPP22/va7GemiokTHEg3Iu+O+KmVzbj1IdtpvrQS4sfhkwr5
vYOUVDeH9OwbCcGI6YcPMGb9mKXv4O5gncPeMiT6D4/KPozuxMfDQmWWPGV73qqa
QNwJRx8d4Io3+ucawnR0ODrTyy8ez7itkYxw43UikSN6A9H3WxjhvJdA8vKeO1lj
KWPViQrrRPgc+VWRwlYSPEUxbSE5p9jxhpD/mEuDYJ5X9etUoLv8dvuX1+K9yfSC
Pls+ON/hTmyemthu9rvQ79hAF2drRfkm3t/IBy6uQmjzEfGiutS9wqKHTEAL8VA0
SyMOzWfPFAvca/U2fZcBE4QC7vYIhgMp8b3dkG8KfAjMg8JNYeJnIf1uyL2J4yBq
I+fmDVlAYEbGNxltvvykf7aLodtiiwO/N4FoyGMLOE+4+MfktZtTwMXfD9fv8Vt8
KJN6giynZ5RAcQM6OXD65Y0VSEVenOVcdenjlxXxPWLm7OZjG0ctVu9v0BwWSriD
XsnSCHdOErM5jz63G0+HHqO/wW9HwKWY/RNUOeHbPdNa5l/fIgHp92yJT+LzD59g
e2JvGkSNDCIUPV5oKBx0vCp/XXbx2XcanfuWTgf/rqKCkV6d7GulIbIjIz+123Y7
4pgpBSDJVgWFdAOt1txjirXQhMTZY/1wmjjFqYNOhxOK6t30E0ko8AXwb97qzfNK
3DqCYykajXn+ZgD0wKK2ny5QodIW5RZyfPtyBM+XJdv7A3aFEIdrfrljwxB2p9mZ
vusdjgLXuUBo+z8fvVi0Gi/qEwYKrwGGKNGwXNid9i9SKLFSFQ5BJvn1ebJP6Fl+
hhY8+xzAcTiBqiGRCmSaODt92gCpultkiV8RPzc7PzAAWh6E4d1CyioFnwfsrGTB
IerDO3X1B7oMl5oA+t0JrfD45NobXNXt0TYAHi4Dfr/xwyTN9XIYFHINSXEHHHhF
ydxIi5HBSVgWXF5YJAT+GjgYDWayesjhP5ZAugxWn/7gwvuCCebvu9CMkLIPaPoP
Sf0r15FqYRHwb7whGxDdUfkWKV330kz8xaB/TrLqI7tlf0A3043huzTfVxD0IpL6
L8M4I+cZUXBLS8D4JP2mFdo1dI69ERXi9AcAcfB3m+nYuULshmo+NgLr1E0rgobi
FmQ+AbX3LrtLiY6I+lq06jHDrnNAfXJ1ePSRECNKpx6INqmZoBtijLpLgHUUi+Bk
/gVwwhasVUWctV1vziiFXm2Z56iqVBA/twITYehYZOccmh4ljQsjknJcLHaHi6HO
1FGCDdT9DAbekm2I+0LRmJolmJBXl0iM4LKXzMbgUJ/twz6fBpTvnKKocgI6HlKL
etvaoOyUoTYpfWKuVBsLIGa86G7LGl8huVz1+xwkLlaBoHbVrULprU5za36Ejk9s
4nIHe+41IzmsktdKMb8shMHwXDaDk4RweM+1x2YwzsMZIs/8F8S1ehcggJlTFHME
jhIGnzZvPrwfU07EIBlQuom40cl7QEX+T2KN13zx8qLwrPk5kX1jqfIieB4bViER
8mHQ42Lqkt9vqh0zrU4FUnwzOvcMb/z9Kvv/KxsDo8jLNtn3RqgD16ACOWzy8Hxm
U54K+Iy6s3RyLAl5OaCk69u4oq0GJDvMVhHpYgoGwjbSoYn5f+zB8VF2n+jZFb0u
+V8m8SksUymBAtCWpuY6hIXyig0wWYhZ7a4SK2G+P4INWQ5G2XbJbM9xUaLTnsQK
JUY+2+Qo0vK28NvU6mddk+D9VAl7AzaUvrgKxKsrDA675aHEXs0sy02sFRo6PqAP
v7ZmBuuhS7KAWF5pbgB3iHWefQtXmIB7103cAnTExPEZMVwpRqZ4m+oKjb9SguLb
+3+96PVAjhHT9QlTM+ZQs+7E/FMnd8f/fUUwMgtVDxH7rlQwP5GKyGcG5JKfQX6I
BXptaWLlut6bAl9efOyis5aqtsVTKpcaCkuMTifw9cg5MS9Ogy/CJ59fl/fTlGKl
SicpZ1Cftket3GD5z0w8l7j2b83CQmjJvqtHCXzlnFr67Qz3Dg35iHt1y4l5Ok6W
jbF+FGB/4dskLXJfPz3grDzr+7lpS8LkX9eEW+fqVJvtA33VkWPWWKyj7VawliB+
ZAVcxBr7VSfgoWT21qqnNtVcwdNuunTTrii9Yl3kK/HdOP0V0SUBaK1TesVEIygS
YX33BDrr+H8KpIwN+w7LiIKbBntzLHQzxj+cfO41hDiq9sBp2P8YddT/XbiJVDeK
QH4qHJHAziGSrza7ZqUpYaZcqXy+g96d7bGmCsM+eAJJ6Ud/041oJhL3jfszuSAI
uOCqYd72hg0keevseMkMNQwguJQaRaZpRudGxqR6wNux49LjSJH2BRaayLtxPWBZ
lTjBaKEnOLbg+Q3CY6BbxB4oxlCrBnwgR9QhleFMT89rpvJfkKQUb2ryz2tgLxku
L1AHuNgwEwQg2cs1H2nNVfaUy/eAWfegYMmmpDBB22Zhuwe5Nqta9P+Ooc3q9ttv
cP71Oh7o7Ar7hCMiBp2ghWd/PnKEmhFcO25BKSPKU4F30ioLrNrzrU/bbp5T68VC
ZhhgCdePXyCrJ73gCamrQtEj7aaWsRNzS7+ZWXiqE5mlHyuC3zGqL34Oy6haV+hW
Zm3gjseORK5dSpph3H6qrYZvitPqzsmOB2c9uXo6SZGbz2f5T63S/gjfbMFdv8Ki
M1UgZpe1Or58bPxq65/X90jiuEObaazbMsuSsleN2teE9xjZm5dColGBW6scdmJr
R3k5YmHf+VSJz9aqA1SpyejcQTsk2af7JD21XfW4sUQ0i4icHtuxW5wBibUp4ha8
6iW7jAX+7Z5dt0W98/wo4PFvxfWsYTWeo0cX91hAiYzW+gDsSS7FNQ9ypZZpQE1A
xszssRVwEi/JNR9fT5hRoqwnfaZJ5yk4AFMKFi0B2OcAUw++3hhDCF3l6I4Rq/dk
pIcz4enpBQTbj2AweatLfGwZSR6sobVG8TIjtJNfzOiSREHvUqCPI5t0mrh+KeGI
oh5sVwWREMnEJHHgYsAG0mtrYy99jyJwT1LATbDfJxybUx+q6na5YjX4USKdkH1N
6cI6h1rX+6CCM1auKtl+2aN+txYI4RQ2+9E9EFH5ZMb6oAjB5iebcRpwGgYCD80h
KOZw38bfufO6XsA4ZlrG8/HY1KUcmVcsccemDVyUHAuKVutlLn+dQJl765X/O/6k
sCl9aLUe/dc6LtAIV1P3DP+JuwBPAsBMISdT9MkBxSi1Sspf/AiBxSowHii9ZfTU
UpSz5uIk+9bc5uPSXUoIxUZwDAThXlmkwonr/N2pBGPE2birpjYmzYoUn8IumZbw
IJguAs+KrfshqCC5YRhE98e0Q3wT8OWHbiT5dG2/geaDT8847e9OUK2lipcOP2u7
ufzsZuENNpAC1EsQTxJjF2b/L532IX04jKW8Ec2eUBFKiK6MYcnffTdPa06YU/AF
h0ZGolz2FRhgHY/2BgiZsw/v8KU5+eQR1wRxzvNMkCiIebglFeovVU8RftnTptRT
S04hZf4CYUD7jh0L7SqzABPwbXaVC8HAcsy8bmJ8qSpFewT3wGJQ6iNf+zBLk72g
iikJjXVXhsDidl27FvKmPpk/vG42x2DQKFHm9o725Cz15deA+YlEWUARYcmUOE2B
j/u8Z3j5127xGe1BMZefe79l5HIrFk/jQm/pWT95S9GePuaBiPGfEmWZGCUSHjOg
YjClpvPuwLDe8GfBvc3464Tpv7shXvZ8dqGbpgrZTyjZQLjEzQQcHiAS2EXtzTYn
XKIIDzeOM26YSoKRbeKv9XpFZzu0gihTcSu8Cg99t5Zr7YtJ1QQaPkXwq1yarVyH
3m29vzxHCsWGeokh0W9fZbritNIFYAqJpVsRHx4v3rHOGf9Q74grVIJfXJw4JM2T
0LAIF38VDu6qILCB5sZecjOQuDBYNFVAQ8hwG4bWTnb++WwbyqZTtoHvq1gzwkAc
xgbtiYFSoCkIHN3wEgC0N37Ksd/dx7ZFgxJ5TRS/vWrDQUt83zrukG+DKYOsDj2w
6JslEZxDHH6cF1wDRIoJaHv1SwilNJqtDMcUYp5xkSXTqiW21Eqe88GqNYy/cG0A
Xu/R82soYsGiTdeD2QWJWUdUpz0cpYo3dddxIdBZzDl1Bpnz2+FZcv+jSm3Nruz9
TyhyWA+6lpVvHt1yxhMD1qq+W56OKSyPifjTHCHkQ1m+j1LlCcwWK1vbw/9LOT4p
P484aOmCFVAahI9ac7RgyTuqbZz2hIb6/D8zrTXD2cr2FbY7JZsn1OtXojYB4hHG
SZO0B8sw116h1I7HbMqameKAaSt2uAR48f5gNS3kVpxbWnbvjOMFKwovoaGJpCd/
7n4aE/0etsWm9AvlFgCSjjlpDRT6YEnacNIgNNsjFODL+6FpKSHd6fudlLjH8Y97
f/fGDL4pDUhsAsGFxei4wpbvdGZmOfxnwJ5Afkg44KNuA4++FwkrZiTP+QUgvDrb
KeFTwEk2ZTAbrpCM2DaJ7W5mRigrmi4Z9YvmMx+Hg1yqKB0PaSrAy1Dqz8uyL5Mt
vbK2M3bZ8lh2BrwVCqk6KQtrEG0sd1e1XEM9sHaVeJ+UPjvwgwLzkE5gJhlY1O/2
JyKzlRySo3OTMwp9Npdwdcht9ORuthkNl4esRe1zJYnRNM3Pp54pjWcAnlpR05Hp
qJm/JMNI8RXhL+KP7IfdY1M/I0ZrZZ4sVvrIpsvzYlfg4PqQh0g0hnoEbsFQ3bmB
7XywwZgi99AoamHLhPc0EPRuuukSPEczGD7RqgLFtZTK+5lVusuwhAP4ZKwKKqGy
c/sfbukMpYQI7Sv4g0uhL6UD+LcQAqvanxF47QlMlSsa+oi8dNdXINTxnFMxTyu2
mF7IKw/bA0OgHB2cnJRBCTyiKXhS+c7lcj0UfvMJaFlBnAlPNOmY+jsqde/mkLta
LUcqOozJTh2Yz3ObD8OvWovAbBc5v5RvE/n21caEc6FcuPwMtlsOLQ5jT6b3S/1D
fmSKZduasR4M8DMQEY0E811KuBYEDCGZjw8sDsNllcRIT/lLb+X7/Sj2EaqR2lyj
lP1tp5YiAXbO5MM6Jcgn5U2f1nj/IU/78RoVVPo9kBfbGtZIX8NRah7Ny/koPztB
5jkqaXRuX2NSQVnPqSHaWexOzHQm1rYzQ2BOmyP6Qhw5Dmq+zOzTnZeAerrxPlsW
oex13x/6tk/e+trkXSTF4lMGpY2kvkdHqjs39DpHzGLf+5KZNz4fb1LO0JUW/G6o
iOEln3M6YT+47gE/NCt61P8ub0V/swMXFPI9RK8gQhW66Onppu3CYmc95CiIu35E
yg1toxDveZcIGt7Feg1NKgGPRodw568pi9vNRVK5rcKfJZIXH+a5vC43SutUbs0J
sU5PnygFZeCCD0NFdiWCF5HXLWZ/euxKC4U/vWyj0e2yfUjV2gu5HHuxe50c1xC2
kaNdUs2TZex7BEJalvc5Lld+WJaSnZwqzeY0aGknGu/AtkyTOMssCN4B/0LH73Xm
VM4I6ZrQ3/OMtLMyX9W6vf9nvhUNVaUUA4r3NCrJbKY2afpPTz1DQz0CLzmH3UYZ
BkyeHQc993fKAeHEzNI4EYhsjERzimeGZzD0HGACqCJHajlwToL93NmK7VEi+MSk
JniXMu4Z4hpm3H/UX7DgFa4VmUXGPH0TcfSXaejLzpmXigkIbtlXjzUVaziNyG+A
mdqKQBhWwW0hJdf3DeBiEvNTo0Tp00gMPYy5bF/G2UWmVqAJDJub8mFK2BhGeFhh
122LcFTGq9raxxSfAhGDTPWtUOl4+U1VBUvFZfcjqeF/gVkGyqIQH5rdNAqK8WUH
2+oDh7H3c0XV70kSXY652TjxtgbMYHbTZViQKB7bvv60/KvRjrNMsmQC62zS4Wkk
JeL6MU5TvBa0tLHNeu4stmhF45xqEeqoBiOa163P/SSbE4ItE5YQuDm+aU+xzJpd
zBX0oqt5PmfLXcudene9fFc7i5LvUd6FLqNI8oYsAOett6Jv5+GtRAX56AtWwCVr
X3Ec2Cmfyc1rRz42vYUS4EN35MXEHbsYfTDerCriJbNCiiV8y+a2JvSnTMCQCHUN
7IX7Cfgma1j9FsVaatEztTird+XGd3GWVgaLOJyxPzXsluy54fDkz3NfYCskROhN
Won3KkahQrcLSkf7xJ6lJlGt57597gtNHwaFNfIGn9Z22faR27+9foEdOndsTtVw
YuqAayLWcx3jeO8p1huh1PS1617WQUyegxy4Y6iuNW29WcqRC0wNrv8NUAqtHdBD
Byrwph57EkEGv1FpupC9SKqYLNXnDEJZzpa+N2ffkoX3ae83yPVzWyn3hLqROx1u
BKAXytgeRlBIT4q7n8HzlyhkAx0X4hr9HhSlkf2STp7opsTrNfLLxKhIhY1vBYyS
2uZDFA8I9eP+JfOkC6ECnquI8/kriTp/VoqE/GaehCB8U8xePhjxD89IkMcPz0Rp
0Stw9bbwHAHaWeSBnavYdMae5mhejJl+wM3SvHLEWdaEpcPSV2AwTx6+wtoYKX4e
iP6pqEaVeZoEUg6q/xAedCCAmu9O0sbLyhKvYex50Gty/bOvYhC5rnUbXIlcbsRZ
b0s3dnLQBU1FHqGvsbeHI43oSzbVExijezBK9bPmg5IY5ZYaQy2Bup10HGq4zXiw
e4F6sakdYIxtmV4d2HdFk5F0ykItENrgiW044pGqoiDGgVjfBYk2ESRH/ysyguIY
InjTyeeoT3brJXyqLnVaJGi1dqPD+sT5tCJDttt8CVIyqDe0mHTCTdcFAzQ5Lusk
Ob6pDv3+N0r6ZGU460ryDddmjxkjz9jaaCQ10/YNZfGH0xX2pQAMKsW9VKGdW7QE
eQvOKBnmfpyHr3JJ22d9DNQv2OxdT4wDegAmykVADkpQjkIlBxYz1pZbHHIBh0Yg
gZbexs/WNK7deMvpdpAGtftipBoE4yX0GzfpFu8uUhBXzWelReXIPUqpoWbjNPtA
DNFBL6H2y6ERYNbUNwKSSLLT3rcVWqfmtCJrH+nxkAz0bZi2EBR5jEMRpxrpOlVf
+fheiXHd9/UVjmV5O4bzdkk6hjvHKswPZNBfRiFrN5oFTnjhFP5vHhNJs8iNUmNY
gm5y2DiNCQMyBynDP0Mz12sbf7WYjVowAXjB8YvKiDmo2jFsVBuZ9thCcvndlr3R
7WmO6SQSwWnoEcJY/Y4UHxM3YkO7dFIYBvwiG3ZEXHEqfnSV3UN8k60rJ1TrWtXy
I1Le65G0quqsByJzS+yjK14nuneb/ieUD8Yl5CkWaZD8jgo+beiuFSB5gZDevIRg
qJZk+kFfdfo6aDDlF+B86NX/nXe2yfvNuF3nWtxx0zryr3rOOf8+5iITHo+gmfLU
R0vfqAWH3qEs7/S1skIq3vb4bd0oiPpNfvNqBgph3hqTdlddHsbp+IhWWBrIt6nv
+UTL8lNsfh4Nm7eRguvFZCGrwykhXiTYDBk8RC79Zguo+M5K9AmStIZuT0Yvco9F
pzj+pL158HiZkIwlU6ELBKIpaOFEpeNwrG3heOREnDerbLdoTg5iTFASPnccGmW6
lsw7iRuOARozJTwrTpUcJuKw8246cAwjgiabqU+y8sNExAag71i3Q1QSLwrZEu7e
Mjl1+S/Zg94AE7b6aL7/e8c0qFN9brt37INyI6f24/hPjTbWj6BwjXLxXCc7EP0/
yQKN8myq6fBVXZRrc9B/iVCwbNKWuW5H3GiSP4+S/j/WTYym0p9hiutAG6TjvhO+
YsCuf4hEQbtuJGMdw3Fmd0WCzWYJXQ07MKPmtget8Z7uwAdH+tA1SoSZYM+Q/mL+
UaOQR9pcu6nFDDTJadaxw/QYreBH73YuC8V0KoHwVwCmnq8RCoK8jkcrHgMEdM1W
vvLu6btfbllZqXG3TqQO86LlEjz/Lr6tf6Sd1M0Xf+kG/BT1ySr+VyIkoJKstJRZ
bbd3kugCNdCSpOFCHfgGhYzL1YQllthyg32elKnh+WRI22FagO448BJVi0OH1W++
eNSwcmM8vjNRgL65mrIQsDMmKkaDLttZ8Z9e7gQYQFURuASGTDVNajlbrIltpGk6
a8ryPkx0FG2gwnkmXlHv2BtIKLbirzZdGZSbdo7oQ8+NncaXJFBrbh1PVy63ZJAQ
21g7OQWealROtA/HvxDrPp6S2z+dTiMf+DUD0Zr6m/K2ZSHb81b1ZkF06pVWPYgE
AhY1WGr2+9Dy+5bPdmovow9Zirw4zFm7apMvYzDwpW6nSjjWovB4G2akP1x++5b8
5U2t8QAJg9v7kjCq7j3Gp2XDsCsRRBpmBh8DAZkDPMNI1F/7yV/3vi1FN+CDE6EM
SldbDU8AxGskBuCbVBAQaioUg9TRJp5wE6fpSGFgx0UQ4za9iqWXt0TYRey7xcZQ
LOg8YF30spqEvBF5mvd6dDIJzJdVjnJjNSVhKLj5egNzvJlxawJ8QAuHt1h0J6PT
qHoFZkhCKe1SES9Y/S3rCEcyR3BwVCKXzScgzyKDkqdSVKkGnt+PgCE/BpGXI2GS
FicpALOSN+AF/O1rVtrIC/ohEmiq9msmuntwLXfU5EmvTHJDG4/HJAD0c259lG8M
3NooBbe62sDpIhAjJs64BBH7IHtSUxOI2DfYSTNu+k1IkHfgklFnEdNc2nsqCmDK
NV7wXeraruK5SY+JW7bI0KO3H+qJ1ceKOf1xhoSsn1ltNx/p4W4hPumDF9I7q3Eb
803FbIXF9FAVdOJc7HUTZuRTXWt1qZRxHfGm3QZn2z3eicJMm30/4XrFOneugz7Z
tKOeUYsFQ1yQxCMzKVgx8fYMMT9yPinkAl2bex85TKHnO1r2ElDoj3bWXHprUAFP
cNtd+C2jFgCjfGhb3y9cUyZIwKmmQ7zWCXhOnAed3NPAZY+YeG6zEncpYK3Iifn4
b25dVFUNiLrIohf9tfhvt3KXJ7NNHPFgWLxY/b3/Ow/GNh3U/aUREP9bo13e/Gmr
cRWlfoWiPrO342CPP8E4N+rC83wNOO5Cp63beQiqhCTh5shHF8pFU5sPTjJ91iKe
lJ3P1PbH0PhvCeSD3m0kReg3TBUGnzjVRl1bjghtkJeLp05ysGqhfxXW4Whbg+XL
crwE54eFogC0GbXq1j4rNELfMMZoHIzHhgKH9JUrPymBgUvEamxvEQovD1vyFP3a
cWTipkm49s7hc0hHUTMeRF0ARoRb/xx9c3f6JNpf6Jrk5YRQJi0c9LpHUh+ZRGt7
eiVSVh8D8ojCxik5hooCPxNSAkaoX4Ht9/iyFOREfZPJ47i+2ZsQlqzisI3lwSwk
gO9rt+WxC/5ANFK9mBS2fw59jl9NJr2n1h+amXiKGotjpvorMVOTdNFeAgaLj2f6
y8j7zcLMhvJ+wPWE6QHTUWGBX7ITASosU31YmHqxueNxc/rEqnF8YkA1rUbwo9Ek
C/+0iXR//cgX+3kigL+T6gK3STAEBYkQ2gHIGORDdoKhqDuclFB7esNX1QLhVRKZ
HIySBEyZSmXXk4X2LQBZRYLQZDwCYc8gFU24UC+xQM7KtWB+MDqdIxcIWb5o+YMf
b9GxAOIe7IGlKaTZJfjy+IVuy62beNs/vbx50X5ty7tD/aC2KcwWb4wPK6062tTA
w3mATjrJr0nqPWgqMdkIvyX1NoBFQmE+XqWCxPLheKw/5jPq0ZovwiRd8X/ecgmt
YcDuOWhnPvGyL2O7BHPP8iEaQMS0zW5PQjfu8ik23ie+TVotKviqmsM71q5k7rW3
JZcFjKMvU9kRohbgOZ8PBYhRKKaf4L90zIR96L2gv5HqliN0MlKhFHemgd70W94K
5s5We6Vn5mz6vE/6oLANO8/qbv+WWJs9dU5bkexJlWl7+q5kaf4mUlTJoh3s37h5
gYzjcN7s+495Ag7uhHRJfNUphvTSIwgkUFN963GX13B+4i6DXc/tqlIGQ+nqe8iO
OIjn9ykyFtsaBjUOEjhSPDCgV+s1dcKzBTMoz6ge74q2SJ6sVC42C6RWyPqR4Fjv
uZM4qxyxtJDJQZK1Z5NneqyoHbW3cRl2Pk1lfZ7jRnc4aIbXBAhl9UPTjIpl1Ud/
8ToH0VE3wlGHkf3aSywoekD2ZoAsfqZeXCkrX3p5OND/YqUHW47gwF+UZNjGJunp
GLjjg+bsI50PN/AZ2d5zk8cMMqS8O57ToEozfkcWnS+993neQG6u174+2xUyvS8V
xG8X7Xav/62kda8fTOWxyRQHSf/7ya5RiZM330mOgZyELtLhg378h9+hnnRcbLcQ
UJugWRGhUBkkkQBY167cyl9q2f5t6KA282YuqTN3CHlmr45b2se1h9fanqs1ZgVG
33UrFokO9vx2NjRaer7LpezkT0ey2McS+V5k7p0SgXO4uU9lkWLxI3N9wbQsOp4Z
OS5Ke7DIP67NcR9UjxO1w9Br9gxdeAZRuFSBrNkYWhySp5tTroeNuj6JdA6pG0vT
JGu3OqKdxuM4725p2nSddunuDNo+I5yiFBmiFYNm/bvS5PuKWraMci7dJhrMMbOa
orC2R3KFdA99DknZdBcce2DQwdeHdG8b9kqZ9FW7mXMqhav5FL5heSDGO6f4/H4W
li3UMhzDXFYieuxiW3m6TR1cTBVUewzL4weS6ptKEyPEOanbYRE0H+Y/3JhxKJsq
ucnVEOTygDr1lg3+qRJ/BSzkbVQRTPI7WJVNcjmw0k3Nue5wxQKvELf0ZG+NllxJ
OeUJ92kOWueIo+JgQpCM5MzvMSduwnkOrKmREPfmveugMT9k9R9fFRGmEignmA9y
8mO5eVgIlhxNZx2F5SdCFvmXqJ5gLvkTvBJJSeYx88ndfNOp504kv3E+Lk2dnWsY
wHi/Vi2iItZL4sfS5x0nVpOMsl+A6VZN/oOLOW/CgsnQJUrQHxu/9vyjbBCA1sD1
MEnovAFIU2yXCUrNw1HmHX6hE4RC9W3e3CElqdeCCUTRRFJok1EFciyOXe2J6CLs
fv+XTWh/TVOkAn1/K5+NukvWxxEq4qUhJ/10b5KGdnyHYkkv4roplI+6yZhR7ka1
CZ6l2NoIJyHQjzQ7ZpsHnVlnsof0wk3+GMhnbXTdDhY/qIrj/kEdhQC7VDciG2qB
p4mQJkoUkFihX4jM6gCbT71lnkymT+lgO+Jbw2rSD2uyqsoiWzcLAx9ZOKIqu7ZG
BMfHT/F8uKvsY6IYyITAjQFLc+U4Q1LojIPmHtWwssRVZCMYBuOFNnpQE9+JJ2dm
z4rkDlAOYbniw5j/hxTroKnamgddgyVO+O0MKnO6tSZ6HCtkrMCgcA0CNOHyOac5
eBlwG8n5C85eFI3c0ow6vSiSL27lEkhVoGEV0AYOhGZ3Gl17eXtXK/kc1g6ejHvv
4/GhQYnmTGNGq+5o5Wo8PZTXJxA+UNlP/gkmcw4N/CukvcHaeS54516yILltdiKG
gQMxnb88331hRxeK9htjHgHqCAKAnPUtln4/bz/liwqpvWfYdF8Cv6FcvPg92sw8
3DEH3IlH+/r+A2DLBDavE4Hv7OpgMiTVccVcA1JW2gj/V8alIkgPWU9O2Jbui7/f
RLECLRmTIjIDXTQEoVFu3u+DotFgK9lh7iuyxpLD4aKbRrhbDj+mvKFJyo9oLHVK
X5tZ8CyONXZU6EICAO84ytEAEbfaHoT3Dwp3Z+Az749EY9OOPpDHeo4gcWI+qf2N
MOp8en94vV65VKXxtTVj+OQMRss4D9+QkGYrDuGebFuqa0HH3Mdh3fRiQ3FTYRkE
vzAY95lUjjMXWN2nMVEoRTKxuL/bs2nW7zNHagdAnvfpWdMXfk0bOKBFKJl9VIqR
DJWBOJtc20+4RccrJEHCDnD5LAexxO5xApKCTqAJQcmWSxKBP8CcoeFtt62jjDCS
aFt9eYX3UV5XYtRDU99uEt2NicNyZyWIB6Jut/JSGEPs+rywhl65zhTm6NqRHhg6
pSDarcCuFvMjQqUyDmc/ebP5StMdSzWC8g5nY9Yy+eyAGroxxfybxeTZ8at8Owku
QqznyJotv6ABqbgQu5skb/LSiComs9v0x/zuzMIFDj93Om4Gs78ra8PPW6QWITfa
N6BCQ/kcXOf527pw9uKhg2EPVPA0hQmOgmAchDQR8tkynWgJIlATtwRWOTTEefih
cXQ4C5Fe7/DpcQLHe0gSde1BYU+HD0O3k3DHQSZVLAAQ1k9+VfoJaYjaNXdWAA/r
c7whRYktlGBrVWATTEraShCpibq2QXL1WbGTq5zIIQsyrVj4UvdSsAVSJA4ocvCj
hXc0OY5ihz4d2C2fPA5loXA806ZXd4YTdnBeLay3edE9+exVD1un5hmwTIsYoLKQ
F7GYGzPwbrSBt2D0/3G72aflPRtQX1Zy+Y8NFbBmcum0jiz4RrQKw/fxwHbIpf9W
a0Lrmer+pu9orR+TBdPxgIcC2iBSSZtHbRmfxDOZrbQAq7y2Iasf/QFp/BolJxig
cxEo2PDvZX9LvTb4hMlAZNDgzGXXgdFtPhUaEnu69ao5IbOsAteLHpnHKBTH/KJ9
6Qb2LkoE85KtgHm9D1oxXeSpWlU/RMAWAFLpnXs+RdEBevKB9Mf4S2R54B8uo64/
a1I4RGLllQC+xfoHHHc5wq3w2K/VJfzwS2qoxmrtndBhdmxChdyDrhfjtXYMFRtf
IHymjzrzuJLHbOUH8M6UqVv2ou0lbHuPOCFymhqRpaZB/vVWtcx3fJP46md1j4Q0
44yEz7IbL4kV4mHyYJr79+0CAbJAvNrEQzkPRIcUm8P/8FYMjDMMomxynZl0//aS
zH3wrFutJR0c3HvyPkovIzLCBjcEMdgIlZ/I80vXMW16jKUpReP2DrjM321kTiGD
2Soh16cJDF4MbPXRneUvyjqYBAs/OM1kGh/3/br4spORBhdTPSE83kqtPRQDN2eh
WRb+iBwIRERdebiobtwMUjhyTTR1AWJpY2hly8JjbBWlyhlYSkrCzgIiizpqYVJY
wvM7tU70Bk5DjQKrgCkPxLgXAbyGWPJOcRTIzEcQ+J/BE3o/onpOeKbJMgO0ayeb
H39J+dcQfV6tHnfhKe4vaY+NKioAALJB1yZBkLgQ6KILv9vHA21RESzx0TIYRZie
BLgaGOaeN2JnRilW46W4m8usNhsRasMOXgMNPfEiSCqQMPwI6yt+dP/cKburWuQX
8/qocjHC8gU6F/7yTOKhu7z7nrYGS6Eipm6RdpdERdPfJgteAAiR7bGtLeAfEEt+
qgEGCZ8UqkxpxV+8epPUWtADun0mm1ZiG3WPm3dfVIslvN5hAUR0mojoV5MpWT3t
9ObKSViwx2CqGk2UvjemDAE1ItIlPUwDFAzr6n4OCOBySTNoRRB3Vf0FOVUwWAw/
z3JUjJOUsu3JMCf+Ab/Z61o5ckJlI+x28XXlA27WLu+me0UqGo37oZp/cl3PZrsA
0obpGXj38vH/5HCy2MIIxyE2r3DvwimUpr/Q3+P1YUiwwFggcw+k1xp/lTrM+81i
a1KWgjXZGjmkmgWchIj28I+i+96P6bjgPKIDcnA93ZYb9xnuJSOzbb9Dvdxs3Bbf
iRYNBJx/aVjlui6UOU8clFfeKJNDR/vDEMwDa3nhEKTOUWBWjCFlP5iyRvXL6OXv
7pJTEfkmjn0EEUKAcjuk89ucMfw/GAed9Ibvd7QZyvA+L8c+GWGeUHv8v6+CeZg9
Rw/k5IHYmfyrP7y21ASc/0VCHm3tXLXoDdQDEGpUNEfdTuI9wYkwMfl5GrIE9u4N
99l890plYtLI9+pQMB9pLWifd1vWXfgVvnPVOyPTDSxyMDn0yUr22gg2TQBtG2QT
zKB3SSjViYbpUBRgHcUxpQbK2uh6gP0dvPh3HUmylhpWZMhsUael6mh/bIL9CxZ/
418yxa00/BbomE/cmE2WCmQPmnh06jF370gMC5A2ogHIkkJgL2xSAow0kiKvHm9r
ENepo0tuYrRSRmvi0PjcGcJNVVNTfWw5PdiMy0AmfjugcjDDDnDv2wOUsMCffYNE
M9elFs63UfetHJCkwh78nvOx4EaWPotskCJaF/7ztsroKjtwGkAjJug4QcwXHoae
8U8AiSN65siPY4irHd34o7j2VgSKVZxwWOdolDuAUA7LfCuVYWSQ+KMvtwO+J+kZ
i81aa5rBT846jabxKNGsmhqNyWPtRSrGR7mkFN0STTWZpn3uHN+z/Go0zPw2Xjep
bUE1VtWe8mxMXVlb0/YsaLmiRlklaYMrNx1blB90+0m8y4benicq5OnyPzkE3S8t
v+3V9dwG+vQnCz9Cb010JWqkSO3fo2WUwvS0BYueGgAbHxmO7jJXkpnY3InYYU7n
xiYUi9BsRRmA4ZbL1M02InlC1lmPmOMAkO6LZ3iItSHQIcxvA2WiA/juTfTmJD+q
TgHm0CC6i0zj289jOr+KrdsKWOyMDaY+oq5MXp4f4Gn343xbck7SgmeeYXP00rcQ
gWHl6F4HbARR84qqeslb29GqKV7qGaPj44wYuP2dmpRb/ZIH+pYviG0ECeClONlh
/o9+NZ8tJfWDROm4Br1Yc/Ja49AuXEkl0yXrXCQZF+ci+iYOtF5DutqjAc93yfde
sfhgDBtSQB7gCYdxh8RQbTsMoZZ8ee48YIaTNvBS7l8kgIc3fhQZDGjar5vmpQOy
nYfYEiDwGKMazeBdPevyJSnjfCG8zAeK0fOo+RvDQgr0lMiBbjDDdJ/Zmn/8eltP
OJjx7ZsIzbDsvD59fResQXACGAZVmOESaX3mTEA9u6e+0LuOCSJqz9EnanXOMRET
k4FgOqi0xUJhypufSL9qKJXp/uCneXqbZFwKyestrGRMvgIFS+009vz0jV+TnY8L
miMJ/P+Z5gaGh5RGKFmSRd5jdg1vpq0W+AJk3m1YAePu4UeSTV6lX6zt3XCPGKRb
wA+nfWKLTAde6CqKn+m73gZnhP26cQ0HJgHhX/3qK07TYr8lOTjDHPLofQHuv8ZP
H1Xf76Ji28/p3xOd9kfoCd7tJpHXbcd98IY9qZNp0ReIC2RkBdCE1i37eRiGJEVr
556Nc5LGgy5USUVSawxxy7mYCXHrsGrNHNr5ruF0icxXGbVKEjOTHWseQC2yyS8c
8HP7cKjqoUdXfFI8z///CysTuN9eIWBIM7knPU3z3MvCs9ql1PWoe8TJkunCyys8
hjMqP2//R44sQ4NgrzVTlGmSCBKMw9FBdZLpTeMXwDiQ9waeIwzQwxmte8UEXZss
SDTjqJ2fa96Lb0iEk1RAkgWn6fgLojMdvZ9yftpmJ1bBhL57pgVHcGnMNgkN6nhU
xdGASlkPIvC3WvwbIKrGUyH5IeFnivj+cINaq2slAiq6Y+CzUegTJUr8eugdygRp
04r6qe7/fYpwaC3yhUqo4X5+YKZ5CgY3B1E/QdfTMKu10AbNPvTxGwB93SCzTKSK
o+fqTVRdpaK6ROeyPPn+dJrm9soJEX9vZkNEXKAmsxe4cnb3uSJaTBLDJrI7VU+X
3nwrlz7KD/IloQ69InU4+2Go33iLG2J5cc+XK1d64nSlwsBqc4iFsWSYgOPti/dv
uNvv8zS0mcz/hLYTMtUcEOeI0bnwNJqZ30RI/LtoBp4Sa+Uxf0mLUs44TKRX+EYw
mWJYoDw7IATW2ARSVcgamH02q3GAp/zl2E8uJVVQ5mcI3/+3HFu7Ji8bEqG7XjtO
Xx74ikDNpn01USIwixXHg+JY5EK5rbq8fHDVJ/h9xFGtdhdWBLc5ZU/HIIm6W6p5
hJFNDnlWQz9ZyIZG3u/ZSLOFoWh9l5vD41pAnZPQusIySHInHXA/qD/YhiqJVy+U
QcdGKc3Wq1sFhxtH/xVcYumXf3JGSuKLqc0V80M7VWCJ2CwxqRn2oDh5Yka6UqpY
Cph1056uLWtlhucWqGmvI1Rc9PDSeWiK1KkBOcWpq0ZJLX63TiX4ngga2xKiNpX1
1ffQu44mKtW7WyjyQZAri2R918I19LiJBYmhZfcNHlocPyKEZOZj4Q7CYwG2iHui
sSG3TEJXGlz3nMj7gfuwzmJzpMN5rbkNACHwxjujUzHJcvypyKVR+BtJyg6Y7rBJ
3SS8LUdoFuT/ypxr6Bn1zmz9EpzV1I2waCCvdzb8NRLG006LLnwQnG1+y/vWCkXd
RUYVOAbIN72P86KxyrF6edzGhvvW6daV2Fw5FnAuHSHhZory0CYC1JcRdYakxk9b
BZjKugiLj5bEfz9MX6BAwhw4OX3E2zyz/1C9qxHdqlMTFbcJ89FDNln6CI5kMKyG
jSkNbRDP0qbjNu4zDPzY9lgeutyCFa+jjEWgGrNTM4irAxYpuebA6NesYAPfFuLZ
hk5/w9LrsUOU7DuKODjufDIWbO5gO/qQFbqfAFVnzRcwn7NXGut6F1pu/59Mmk4R
uG+lK0K27RIGaJKONsEBrm1s2l5mL8qEZxoLmDEWzKbofifuz6YaSb3cJtT0LxAy
cYcNgdpx65i/1RW5mfDKfnlwafHSkLlwsWAzc2Zd1f6JYtxZ7TcE/QBDy4GcbPFJ
Ih9JAnmznWblT3F9xfEzHvENUvnuB3Nmf0ntlpFC3YfANx8IYSjnIT6FLfF8ssOM
gzFJ3VfooIn0972zBJ0t8RuedAYJb3liAkaQ06Et+tx2G1yQHKmbR2dMOUOkPO7e
KW9i5oycsifOcoHbXGaz0Rxvy9cod0YgzVKrbr+CYET3lKTnlW8S9SWiUJBm0Pvf
Kd8eqURhJUJ83t+XQ/q9Rc4yephW062y6eTu26lP+B2KcMTTsORcGtCqJWCh37hd
2PKSgUMkgPWT4NUZwj2wqKDUMwkkxd0wdbF+kxe99YSsgcq64UZydbFDJe3jjzcb
QR4sBWssEojz0kneglo/ULKwDw1Q8HzvOt+Wk9OHKmZec4DaKKSWpoR1+6fvLFx1
Dh3EFBGRhFj1KBw0AB+2SkqzvsOVQtriyK20tqwqYh6vBEGqxjd+RpI4LbqvSegg
6kDa8aYEhIVJ0S7S4IiQ3jLYy1srHLOhE2veWb0C8BD47EqPtuMRbE6o3K6ZjCfx
qWob//Lpaf0feQXqKLs61m0gJfl3fKMZqWhqsJZG+4AHX9kqAI1fLDgs5fypi5O8
PdqBIDAROWW3ApQnN/G0/63YS21PXtbhwasj6+/7d8u0vaitnuf4b45Kouw7f0LH
XQuEcc/1d5O1NJuJFKyAkoxflYZiy1p05FIEMK+yTbzAa0s80USTB3KOfODa0SyG
sR8Fq8YlMziO/lNDY39j4Ssp4/VmbUGQ6hFfD1oDGtDz07kHRVZ3jLf6S3fx30LM
WnPreyI0qdnoSVOgRhkgnOs1vv5wgE4seQYD7K0P3jRQe0MBjJ7pcqjhKbNkZgt5
6x6n4jrBKhtR7bX0DqnTpYSfK97y+YWVDAismv7ikgLmokJC3ZdfxCe4C7D+99fk
DNmpE1B7Xl8wqc9NC92niVOuf64zFcjhwnYsYbR9paSeAK/BQFssGh0ZPGsdU5Ca
7TQ2YHw5kMINyguaRuvkVbsI/tmRsFiJEPWXNik7Qk6GlW8kYtt+iX2H21OWkuRt
3BMtr782WfJ1QDyYbVtaZGHTjtbpG9FgvFNlk+T0S/w2LLXFTcs7BvBcEF9wrf0L
bulO0YwsaMHBaTACsmZSpotx8s50q935Ehib1ZyNhzFtCmK5XoyxZNIq72PiPYMy
ij5FqEpKtd/NX85iSGGtOxvrkvzwj/DAJe5hmWrVCM9UtIi98TNFBFbARxu6wkES
GPTV68QTi2VFEL1r+imMD9qePmidIlmIHo0rxRR6ns4AuNg3FqIcBW25OccJvsfe
ivaeqtaydKE7GMZ8kFSRMxO3Q7nVtGQe55AsCizr01uWoGCHRDpz1dLQLzVEtt6N
xo1ByrOh28Bj9Qlx3vr9j6l2HLoHRFGNMk01kGNB2Grhbw5yAi9HnhkCr3yOrFZF
jvyOn8EmGWIn28sC57QoZfT6aCf8fXLyOLalSZIjV7qN91vK5LR9OXo67ug8TutS
A0YkyFNC/wWm37y27bPV/0a91iZwtqNPL4accQCdPIws+ssCFNUviY9Stu8Wf0yp
KT5M8/0ZpAVoAhDreUUC7zDvTx/3/etxt5sZrLnqPLuA4+4lXEx1ux6JMmtJPa9H
Au9O56rCkXYTexzTwPZMhSgPAAWacQxHFBChbaQww5tWjJR589p9OU4lE5snWKbS
tSXK2bwifPtKeGvQFvYDzADeysoN95igtuFD5D7glimpvXTSEqFJ9RFSxFKOOBah
cfuefOsrJ8Y9UsFQT+BHUivc0DIYQfzN8+G3gCkikEcwiZlBgvzaJmuSQ9vGRGbM
iQmeLkMxSy2108ebOHH0Zgv96CsQFFzYzCImaZKwhyWol/8pBOdGdSPPULHv1zS2
3BxciucsJvYaxaF7VVf9t3VGGFEYR6TYBO49Y4JVfk+8Ar26sFiPPhlHzdwhtj72
Ag1uIhBJKOmKEJcBtPNH1iCKDGZk/HtrF0Q87oRfr80nPLeze+Km/Wnut+wNhmSa
Ka7tQ+6B5t/FzragpiYmK4ElT8WPWZA6oGo4Mlr72/WmTBM2EmLzDxY3snLx1/bc
v9Ug10nLZ3Y4KgPgSs1RKSrY+8vIacJieVqTHVhf5+DM1JMMALJ+/nR3wQ6teYIF
VT11SqR2si4eBqJZPC3K9dS9Pu5B58QJP+4N0Sl+7dDCiSNt/mvR+0XNju1r7EnO
kREWc0G+PDwDxr34D772QZYUlb+1LikpnkD19foM7pSwSyoZf9f2AlcP2ZDpdLma
rl1WuboGtY+QDS0G+5Sa6iW0mawqAj+ycSbncouH8kwBiZBRr7C+0ArswPI5QMw0
9zxBLoFLghngW4ebGco9yeT/0GLRxT24Vh47BWavNp8a+PjGHDxNn2Rn3O9fVeve
VVENKgEn04jyyoOzgUb2guMNodJ8u9EJvbJWDNgx8mHh+hHWHV1lGcpaJZCI3vyb
+IkhSxqL5tzelH1Pp0ZtLfJ328907WM/C9QnMrwkXyRQ2aq+nxPkbi8EFBNfao2i
Ub4MOlNL2nqVB3IbesJB19peCh7GCvKPkr0WatGDnyJ/HQns2freVP2nSQr4qmAc
626ULU1l4RluGy8cKE/PZE2u0/HNDt/ZIGv190gacUBGg4kLXUp/+hK33opK5cQ2
OOekobk/OPEy+Xy6hiEsJZl+zadACxII98zD62uWlKlcbghbGIE1RmoBF7JP44wm
h5U31wRPdE4UqbFXiDvBMCDn/Vao6Sqjb43y5s05Hj4C01UeCGoHD1m4Ff24ChB2
rqX+/HfIVu5J7JnIq9rV5H6rbH9Db+mpIDMRDMrwBavkIUsvSITtoJe5XRAvBDxK
BeRrz/Eqx2GstS+6ShqWbxs1WCE7Tr82gIRt+gbPdh8WaT7uIkntJfeg40gqPI6L
jgilIFcl+epLn1xnWQPDxFKQjwD79/so+mlIjYZwWv33dWWlVt6SraSEQtkPG3zo
Eo69rMzB0AQYJsndZyPE7tUkwApjhh78dH3Gjuwn35NveYlYNiIoSiplLD8UtnRd
4aiEOuV61VFIKU4OydFR3+UOjs92ydRyA49yO/xXPB1oCqwLEHvBvFPZvlnTz98z
58t5ewUyCzqgKXUdlce+59JDvorfGpeSLfRiDGRrvqQS8Sa51CFLxLPnrTzGdxyn
Fx2/sff3NMWsLAZQCSIAZAqUnY+ktTM0rH1m4OkopYIfKI3Rt066lZoK3xtv5mKX
79k08/KhhT0Sz24jZ88/7oB9SLv/dQLWu0pgTpuIDuUPTw/d89Ar4G/dW36SNe2/
BENOYaXmyfKo6Qi7VFQSzcuKxQybRYXLl3SvDU6UAm6612ZYS5QREPec1W4fCAcN
KZDaG+as2PikF6evMCzTWmOrA1swX2eJO9qegRBM5BLChaRU1heoybGmDqGMTjsh
0sJG391LUxs7AU1PU4xQnixAgp86V6dcfbXa+oSrJY0XTaYahKfLAfB+627jeGm5
8JrZcGLYFy2cIDsBMq1RhR633gNTGMPsk+UtZGozMSAubUOq2F4K+BTiw0j23S8W
NruCxpbd8ZImmaHB7rtI07Ok9qREfV+O3/62r3dWiwV2KQHl81NVHWpujYV+i7Q6
xH3xNy5ER8fW8s0U7FTxCec0t4/eaa4j4O+r3xMIUGczDHiND2eMUB7PfFNSdEtI
lnhBc8zQDPCXVSVApXRuJonp56Evv7BvBlcOo0Rbpu8231iCzpHR9uMptIwl+s/S
ggbWNAIzUPaK1TNu5smsGrGz0boUVRQngN+XwEfsEJLJPSHXBXLmIAO+pAPiqd47
vMguiEbNx/CYbpYywLdyHg2E6uaImOGgukLLrsfWENHf4dqNXHyul8RMVoeBfgYO
jZwnpDyz2FyhWQMij63rJNvPKl8/FuG2CTMjZZsrIy2fp97+Fr1cGOF8WnTlbVmG
eRY/DWjQkGP9Os5pgAYbJ+VMEHCEZqzVOJ21b/nT34URW12uhuXULttx0mlIiUlR
TtaikY8WhpgFKF3j0HIsBNFP+x990C8H0DoxOn9JKKdYs8qSTtm/6imS1odp6oOS
GkaBawj20tgaid2ELefT4HhgbNT3OG5Ry/gsvKfZ8XwlhzzOD+Yq5wP/uNqKYhAQ
9S5GkhHtv32bTV8fqmoYaItvrda64OWadEb0TNt1PRS7j17iRxqkgDJiqblbRkku
bFMwL1brtjGO2w8xBt4a0ive0sQlMCLO2/Vk1U00eZK5zLqGGsw9xxpKxqN+ev1X
J4TTdB+RLIdPmdBCQmRf1WMQDWtas8vYPStHPhdxWgG1ZlZA607yqb3tIvPsCxTH
kRSGg0LiBGklb+NseJEx7Dq2R3d80WAlmFrsXMUmmdj4WVFQ2UbENJ9D7WYH7HZx
q8O1WfG6DVhumnQugv9cNQJKfm91Fi4zjher6WGnVCUF0iLBzFT5rV+R8408qiUw
72q9p+kY+ZwU69VV9tlzD5SJnG+u4Rijy2a8QhXRoeUCNT38XcK92sEQ/Ihb7U+p
7wroLsr6Yrq6UMYL6F4IPJ0rYwgcT5Ot4Rkx1Jv/5zOfE53wu7caG/72dCssa52F
ALU6jQR9VooX3xuqvDB3AC8Bc+t7QqTEnAebTHC7N00Mi+elaNEChp+n5taUf+bY
3w05ErQxL1b75DYjM/qeivUA/AcXYaG7+LeHc8uPF7ji37EivXQ1FrcvSRYPsejm
96kqgbKtqfOyBuuv6imtHYSRe4z49VrAmJdk591UtOnS0VN48osFKk0ekMw7/RIb
LKIbWfWrqqj5b+XFyiCW41O1efQicZRNiWeJG8IPleXMRrLzV9wd6pFHk7Ej0oAh
OVK+aNMjSfb9Gc8rMSqNQJQ/4iZ+SyiwRpsFeFc8vCrbAbvQK1Pw1xfF78/Qex8z
7JN77KGlNsaOwjEo53TvzJv6/pY+3CbzNyOrBPxsVwwyRp7+NvNNHETdv52z6m+G
lRWEbdNfx3TUZnJBghwHE+zOLoQ9Qv+JNlz9wH1H8dKtxD2+kGjWvPuedA45vEnW
loIXRlvHQUez2HSBdzUt8Wt9va5IqP9n34bSl196798yXwafAdbTsr8vWHWyLuk+
SVRy8RTNbq/U1wXHkFFIWrWvovSOFjUY+h8XljLSrLC+v1a2LPKQ0uCAErfeO1yd
XZQcT1zZNK26xYNZuy0pXBZ0LJBmdJknb5H+w+iLCiLAu3mdAuvGknndJ+JV1lDg
sYARd415HZrPHg0sOwcSaxg4eVFkngSe+4EJ4HLjHGVftJmUD8S9nrMBJ2PZa206
M5ESkGVL+Xlcdbm8aiVg+fuHVwPRB6NbJJDdildwNw/wIIu33s5T/TR4ezdozXeh
jeTzosajPcsfn+RfxkZKkESKN1RxnTaK9+50W81sK6sjU1DYOFu0xnLjNbneDfUL
cbIdPW+ORPYT6Odqop58LIBS8ZpcHy0m8C4XiS7pTKOkp40lf7Ei6JOGZ0w++gUa
NDeI+Sm1B4MAb2F9FpdQ1w6OsRhODNApc9Kysy09NGG+VO2+HkAVDOWo39PdOyN7
azOyFw14ZrR1Ag+xuSUXVyxRzzuaEtK4fJ4OfEdaqt7gU3QUHIWpL3eMZJJB5R4X
K5O6478Rrr+8AVQQn88ITKgBi/fFGaiRetu2uM+WKJ1kcEGL8v5OwTnYq8Uli+k3
Sz9jGEkB9guaMNwjIliL0dN+JOFAdeP476t4Gmd/3LBfBGzOOwa1MwL5y+9lkG7I
9znG4CCKMkydyf5yo12C5vXOypKRP+9uPssX4EGWHGoo5ceXCDqzegHhM8KtEgLV
2UQGVQ2Eddulr9aFQiRVzRVcBe/rE1TKgR5TF6+y8Hh4+BTmTqURgl9akNW2bb4Z
8rERaEqXVHjxZqIWrRL7u8oxLcNz2KA1aMs7dKFD/LajAWNLQmBCdGtLCJb6oiyW
bpK/kSse5ecdjRWA0xSQu+ujG0atf8dBenPHXzvHZIj8OOIMgVxfb2IVhoEZ864C
IdUnNeWFDRje0k5edYgKj0w0wcK1bYNQ2lUh6EFRIxW7p4/OerxqR47x5+V9drD3
1gcnwO5rGoaTiptgdSrf9PaU/fsLfxsN/gZvKyQnxDT3PYm7bp81TlwUs+wx/P2J
PsCBRMCts/PJYhTiw8XkgZV9g/v/QtYYL3U2/nYw74hd4HlhxkoDfWbpT1mrhcmz
dhXBJPoenzcjbQLcpUfWdTxDUS1ocWoetqxvMqVGPW9zNX70+yLQPAs1i57vkO92
LAJ1BN3fybUUlcqD3f4mCMg6lVBsMl6ZLGcAtTczD7an3wx6qvalhwZ+enH3s3Qe
ZpOO0Ey6fFNwaTfRcvVFQ2W/hKPjKYF7C5EhGkDN9Y0wkrJTLkbGhGbtby+MzCDe
EWzr457jeyZzW66cNp1lko0SrQus+zKqVYaBLnPgQYsMK6cgKXc45XtOd2ZEbsLF
zEb/zxCCjTuYQ6v0/+UZ3TgobM4stn+biaiyepjFB/ookp9I32bzzOlZdjgXyM1t
eX3UuyimI2zhXQdC71/p2kNsAksHlAUEoAMawrGn53tozmye/dbH1yzMviMWZMqg
2S9BywjDsyztpih6yICtNefGnxFpNtkTknB3OB5JXkxfZjw555A9SSqCZ80llVFU
5BO98pbycOq0PsnvNTGbIVod+NZ95jyNaIJgqAgpnPV4d3L7JbpLwTalJQXTU0cm
z+V6zAhbHyugivkd/lVUfUr16NzzxcepvvAY+LiyOadjVmg2Gu0Fylcaw9phHVzl
ERQ5n/as9xIAG8ZweutkmwzxJPsJgleRU68gdfN5UlIs0KYOLqrqwVCCgT8SH7b0
2Ly6eh0nxHzaFeGp6j0fpyP+KgpkSxsNT98p612HA6AxyJT6/B48MgfPEpjg7mVf
zjf5INR3iw2fKolc43Xfs5vtfG4wwr419+6V/UC7N5wTWd8lsKLuD9VDs+rK2J4m
dbBJiIiMPjNpJxX7jbIo4EK7J3KtcLXgoTBejnxhuREdjJGJe9qvAcT3wxzIXE7X
kok71ob7/o8QI4OfFCnOWME55TTUp22DyjSPEnt/8uEhn1H0f7mABRQRH68vF7ml
Pz7W1iR4kjVEZIY3bvl/4VGh6u3yubq72E7uZV5FOabp7PGTgPqoluEjDk/89LDA
PbWCjFzvUrZx8wfTroOpHFb3H5hZSErVvy1huHyJmAKWh2CNtcAtI1BcaLcE4+dd
WEt6gl7vZEvKrsHEv2jMTEOrWFYyXql8kk4zpa03cqbMamGvl4taUMCLfY+af9Zv
PczJA8cE8FgsPRKeGE9+rtdtM0HxsWNwPEpIirQBfXZ49wQKGtzm0oCf8dxWkzUi
Dn85lPhUBIVUrQhsb9jdfpCLVUxe5d//+gJu3E6WnVk2GFhv8NUqYlDcM1sxwsj1
7FwWSc/mz9uePoW5BlfomOqlikGaT3eNLUnVffzkCrFOzxSUdH5+BeockIrZ+EYk
1TEAyQ+np8TVlWJBsYcWPWdGLWtNPjPIkpp8jjVoEsSmwOwE7jSp5MnfEihyKXgT
vf+fwPkgvoz2mEFbNPaxIdGohoSYCJmiM5rPWXPbRMKVqfnbubDnE9TU+udbgJir
NHfTgWnjyrVYJA/LFnA++4qM1JVEeOj95TbOnY7OLLhvqBeujXvsrIcSyNs4NKEW
DJ/mE7Jy803sqPf82exQGB1CK1arWZwFjLWsq6wjCSXbpPWcl7rQanSpjaFSllkv
2aJvBm053Sdk1RNtBwenXWUpDq7qOjn251sc95vKnC3yvizTZ2IU9VckHDXxeOrA
MYUtwEbTDzRXsRTmBxDLVtFXug6KJer5R9olTTJ3132A355eK5I5PzLZKTj2hWBb
7qIj0yx0M+j6DmKneSVNvpKi0vgAvMf9vwMaNQ9euK+l9KnNQXO5BfHmWOccU8AR
0iHSpQwKVWiJK/4EmtmI1xxQz0i+gkJejvXxxcr8Zg3m+IgCyjnwzng5nNhVjXqq
qBVprQX2JcCZoTAQq8zTTDcTQXoB39PnGbTKdnhOpov9uX9RRbDte+xPl2CiZciq
QhVeYf5IxJczYjJnjdSm0SbCEdolqmKDdyoUwPHf1uUmeseBpFh5X6QXlodyirbH
LbNjKTMV4Q6SNHjODQ19UNAJEOo8SpIXFnBtY1hhjXT3dBUomJoLa9uqG5EYKch9
KM4jj8SWlgIuxaReZZ3XFft7IPPBNiSqPuFMWlawtX+7MlIfHyBPJ0FQRUXtRHfm
XrGlQ/btaCyJzYbxudXZhcILkUK1kHknLgMy+NLH1Y22x389x2fbP0Y2GLmbe5IX
C5nPkOg6i0+dIZ0qnD8YqY7qUjy+GkDGCnElokULCRR1AhCjef+EKjAIbyyKJpfx
8QSE12kn0GHYUaNT9O4eAp8S40KEO2fLkhl2kOevXybqbv3JJ/abFAJue/j6JVUn
PMEDF3sQrXz/BaipIgWScfEa8lYrJ0Ii1+dHafwHhyD5iYyZf65nz490+1F3J24o
CrPZmzF5xdOU15EKoFsxFlvvo6hue5m9WxXpkix/fMuc2DfIxhj/amZddrLuHKj4
eW82x45yNccP9pib8ULx5q7cKbkQ5IqKUVto3m/zZi8OweRUJK26/8tQgylCEO/Q
svC4C5NF9m4K9t8PchPI7gP/oZ+180L3bbNJPE5NJHYO7yIzkcCCQ+SHcq7pn76u
7S54cIPLjxy+/qBUSIhjOWGKU/5oIQNVN+eK1od9S3Y8jzjZfM1SUGFQJTfbHXp0
j76Ao+0PAvrSAnjFJzOl6Sv2JVF0bKn9jmdYN33IwCabDemObYs8DJuX4WuygP0f
fjftCr/WMugfC+S2d0gYmsd3Va+K/h9Bl6WBHrmg/hTBLrnP/67mLJ7QK9xAaZ0n
W5D1WleOWwHTVNUk6zZuccgUee22qeaJftul9mheEd6Ck6fy+C+ga0g0VhB/RPuC
gczfU/p7hZ+fVjw9cGENxqjGvmUiCI1I/mOgMNnqHWh9UB7qtRwE/F3lHDmhYYzc
zEatUCrT14tqyw+Ehhl8ne/i5mlw327KbnHdsyMpt9qPW3/NF4bxYPH3RoNWJlXG
QkOhBayBuO94nKb0wggyG105XqJtCmbBDVtz8INJtYLBNX4c/OiC/BwMhT7kIhAs
jzmKD1dYuw/uCrYezU2/MECUaIINB3KKRshyFx5RU8EdQEGTGe+L4horKchat9V4
J7YBA1qPTZN9Wgizkddgx37QqPG1tN1BJEB5qgHU1wQgai2xli4UX/hEfMvwDPhA
xVUNGLKkkvw+Jom7MWz+26hwlxjDDz7f0kSJkm8p29O25dZMV1fn+jxApnHAEOA2
r2+sloPNE5/PIeoY6xhbpLA0MYUXoaQwL1asrE2GwLOKF4n57W1QyiNtzOJWmBnf
WJGvQ4hgbcPj+0xYz4IDvSsbLIk5TZI25Ph2/9vIRaj2xsxpHoCukvbeWllu5CRP
isa0b++xTw9o5SVwJqfcv9NYwsOWltw0PNo2rBgt5bEFeB/5/aYXTV57xZKDgAR9
zdnkajnFZxjKP7llDQme8OFFeWnFCL0tdWJY4seghA4Mwf/2awAeDK52wcXwX9Mw
2bG85Z59IMcctL8FQsNswsfLJh2yFLQgvNB154VOteWtQMHQ8A3PPGw0rej5Z/fP
FMpA9RGyLFMzjUaBraLhkGIaFO0Zj+1TVdpq6noLE2X113F3JGyJFX3JgiX1LFRD
JcKToewzcJGsTD913FBNXIbY5TqSGUR0XkzbMnrh7feGjzuldA/diUoZC+4vAorM
UujMpkf6H8D9H/UIxmjK21hYXzG80pOzZXgyxqo/7oYM0e5Y0nRQA3ldT36KzRHW
uxZ6kR6UH89obfc2wA6gXroQqy4MIgQr8kX6pRljOySKiI3RdqFXKJg7zt1wbZCf
EpAaQBavrJzvdzlLIn3lHNETnEMYi+IqBMLXM3BVIfVg3qHpvRoKMQD0ScRPr5p5
ODKO9vlAS1ulUF7GTm1bWeUjn9FVb7Sfn4AFxL2c5rFKOzuCxY8XdYWdO0JBZhlz
XOnnHU1GQWWLnCR55VpqJl90+udF4O00AX0SbBlyWrvUmyGlH7RN1RzS0z64Ohvh
Md4zt7OSRG/TJYI0DotMamJhhRBtm23QISas8YPvnTTtTjupEzl9joHIz3MiVy/1
M9P0Z4JOcBlC1/Lv2+fFDrDV89f05ePT43i/KXZXwdNsgRZK4hOqd8eWfDKN/Tdv
E2VB/4wa3x87VBSU8Us9L0/gzgymjwL5iGfBpKDiqobDqD3T4HJOYQ+rsuRnOFHT
77HFiqmXKtpeOorxvc37OhM6gZooZgjjgXhrBV2Rhyc/Zupfiz3RnbjimR9GM+50
JS57ZQRma3HRc3N4C1LmXJ6UpCX2QsDvXYVkq6KwKaw2S4W0o5qd6hZbATXhWsGE
+6nx6tJi0gK8B4oL2Rq51bgNw1X1VjX2kzKk1ntpKFMVzKnpgShz0TKKcoJ/yUF+
cVR2M/t/paS+f/pzHNUFkBKaxcdYPfPObD3d67D973YVohaN/nm+VLQ/bHB0z8qN
2l3zuvLJVDgCKD7pAgHzzm6trqfCvsZq0JG0MEld735Sz4sqpHu1UXaVFFYvTtta
uChT0+RD9R1jxotrozrEI9r+HQezuFhuXCwGn+wH1by/XjGIvL2Cw1AL38Ds72oc
eYfTEbLo/YJ6Hryab2USo+1ifP3xmzL66ApEannlItQxuPmuslscNd3iOczeZxJP
cpq54NnKSBEyrQJ9C0xT2pigtwyXm+CFdl1vyQ9GG956xP/xiEtwVeJ4gKk/3SG2
dtXhABUfSHmw9BLfMqCleKkQwIALTyifOrCb3/LIkXeDkLO/a4Q+/oPLi7P/r52w
D0AE7ZNKy6whrhAgXTzveRGQAaUrKhXG4frw0HHuKrXfKCA2sxQpgi6H4ovYHbvi
NY5yOpHIFGplVrPL1bvIGdOAKQEjq9nr931iasBoSdygb2AoP+FPWqu152jZF9ky
vTYKtH9hxgtsWqF/6VnOd8M0maHDm1SYPF7UyJqt8cdzuZTJGitEAwTOPzG5XFy0
ul/ql/upp3PV4yWFresog2K8SAII7JfdqvJpcUL99VMaxWOAt4bM5O3KVAJwpQEW
W+i0m6/jCi/RYiKqsbSOMj+S8LV5mzcsDxOGMNT+dZ0wLzuoJ8sP7MOcr59vWO1H
F9gNmhW/pKm1be8xAYOeMB1yYLjqklenPKZaJto4g0UkYu6KLuD3IVzQ2XrrOnRY
3/Nrxhtt/pOhHeYoUDR0H8/uKaI12FbK4F3ue9SjN3nD7d1KQRrCAKKm7P6f4oBi
TrOxN3DRiP/CxLrECXwcxxVbt5ohuf8NuKDLeG0KX8b5qB8I9kZpm5H1c/lGxs+z
G8QyGCdSs+lZFiDMUq6o1zA21LMSWKZ6W+c64XLHuIAQlHtWwF+SwIVtFdf+fkJc
xR66tdh9uimCxtTyIIickyBVi0C6S2ObIP/mowGO+xDuCKTHOE7F57OhSKf3L0IO
D/Ubie1N4DY7h3kU7KwQqOII9M9ifvyBpq2uT3HTsI8jZmg4RAC75AHRF5MuWhtI
u5WpjyXtxkPLOsbRcEwrqemTuLTCef7bnIrSrWF/zkgWthhCak+4maLMwhz86Exx
4XocB8q7lDgzzLr8wy2Yig25fxcxvKYyVXX4zT2JWX+5PEDBXV78QE21O/0ilgn7
DqlcWpCwSZy7bqVN4mZj7v54+MokxuYyJJnxBgwDHfu1I/rcK8F0RBU+ZXSc30r2
wGiF23PVg0xz+tdoHoSATS+xpYVXJQX1DdHGJfiZghrFIQp24zH52zFYPPxDe6Ee
ybr6iSb8CxCrp7R6b+EdFMFjpsZO1vPE4pN6IM3/TLlaC/fnnnS2Ld3cl/anN60W
tAzc4/Dx3Bo3DVZ4hpUgMmWecqCM4sWZadu/0GZbHe24y4ngMZEa2c3lYkLI0dOB
StlVI3Oxh72q0UfXggFdxHEBGsYufZGN2S0erXN2h11LSofBCiMw/lqm9eFqPku6
x4JKOLhZWcXopOh5VsElRr1JqJ5xDjTNAR4XQngIWVEqmFTvT2IfD+AsNP5skEty
RHFngIhfhFdVnhbtoyaG8imuBffzg/Sn8FSKh14mulnM51d5VIVY0cznPpWXDZvG
8d3p1Jwc7NfV0+EIr0CPigMqleMUgdG00eu3p4Q35qlx8QbQp5DP2eNlsETNDlXz
KamF7nrAmt8n+CPlQhXlROq6KnnqIVnueMOj5BrkKzn8wR1EI00Ye0OtVPEfeOsa
vNKPNqNyp7kZbbXn9H+tp0hXljdjibzkvzsdiN7dRj0BxPydr34zSQXEUSB+uQww
nYGz7sUhk8cumqqygEXw6eI1sSEjjY3j4tcB+nSIbOqLzZgkZGDkxjn8QolADH5e
7OJGocWGmXTrIbJyMyeRIzDT+V5aWJ0UFmfelsZLBc+8x7BWPgV0isVMRI9it9iq
qSP/VuRq9LmU18WMxA1K383KUzh2MydOqoIFLmcAendxxHpxly+xBPnEh+DI63cW
+VCPL7FOWOlGGdueAhTb2mTr129+sZ3lieypUhVdaGjXeMMQ1EhjMvgaGeUA22Jz
KZBBX4uql7b/+ASYoKeEXKLb1Vd5PZ/WkKMw1/hnbxSlAfBQXo3fJ6UYUYP46OpF
EdAzfGeLaDJi2+ttuMueoR4ECLFRsP0i8RTOeeIU64e2+EkD5YWTcn6ndLFLAy4b
YH09gGd0iZ5IUdvNwVErMsBd9nsMaeoFMiJuAn+YmrR201OklmGEHquTwDUSr4yg
BNno9oH/NYxumhctgqY6vS5zssqXFLzjIvIhPk0qKe2+ssqsgpICv27s3Cvi/Ywi
TlOjNHUr7TK6DdkNbnrZMF13qaoIB1hjUruLiC679eRPb8kYlfZcp6bjF6D7ALM8
v8+AITn2XwAVFkwaNFnaUttq4perWoMly7Uu5O54GZMZl7G00bZ5PFDZkckGEVah
VIx9FEm2ZJCTQbONaPgLVgAqNeq4sB5Nl2vF3pJBIF/F8dyKZsjEz4dzINPZgHBB
QyAhIp+sJuvegXdFfvBe8sLdzGtrm9WxEwjY5xiW58sjFSb0X14b1oVgoLSXPvp9
FcLvOzQg1vO1avZaKrcbfrAY7hW8Gomln6PHuOSjjsHJnw5Rn7Jy6F75FbTNxI9r
YpC+c7LDh2309ZYLuZZmGk39oxgel9OPiMDAYzYEw/7aiJ4KqnSIKQRa+o6Vr3pO
geEguORGhc43HGxEkMV1puo1G+Th1fdJ7zBcYiw2NKU/pxXplmYe4gIvVYRDRA21
UZuUg9gvHYOAPBauKCApbwi9AAokeAe5uH6uZIiU1jRRXdCkHDiK9Sk+sczltMu4
NwRwBiJD/CK1m/HPq/y2S3nYFWDtbyKkQu8i3SQuH82GEkxAHulK3tB2k6RYCdlL
C48qczxuGZnVQ0xeTILWcTRVgNLnb+o6o0gJpz5xWbT+N5bBoXTLssEL5/vIlNVU
Y5+ktHKv2toCEMcJjEFBKG/g+XHxbqWDWJLs1VQZggf1F/FKrNbdf+n/bghx+2Bn
XBkR/+LjywjbUK0Sshb634rZ+qckkFDc7UHzlpMmAoBzGh26AwORIIijrhQj+BGj
aijVw+okJtet9IMa2/htSsvK/yI8DIcvJC0eDt1lb3LfmTNv23Ni6c8aDC889UNE
JXSM2L4x7+6g6RbdNmd5w2iBXddw2Syg7ZFr1p97hlsngbj6oBxRGNdMzkTABQHf
LYLgA1v8G/XicSZRxJMWhUvwYPd7582j6wNZS6LOXo1YiAl27l5SjEhYjsMRA3oz
W0Am+uVJsphEpwpLa7Zt+qN/aq5PwGB+YjinzkUXcqsqYdqwD0pW6/6C/BMcWIW2
zR76+lkUfGhCW3yl7mnC3JiEjioXiwX+/txvaA3KktAXzPXxcTe4U/+sTIVH1as5
NlZEbVxkHOh9pzHBIBUPzNHnmx6TjgL+u6Pos8RT6BTFeYZyOgDxKdayn+pmX5XF
w572KwBOkLo5UB+x6VGmzHjat1hBH2St+Doxblqp9VJ8VOuZcuTtf53er5tPiUM8
AbhNGnpnRdSIcUIbsYp5NqhayDyHl2F+cP0SQZaIC+5Ny5wwhIi9MHVlJjkYdaEO
TsD2ooFet6Hf5Nz/zKgaTFKDmN7PkvuPpEfzLbIIsYWjp1yxKbt3wCPaOg43aIPR
lSvIP80lV68RKODcjH7TrjCdBnA8yPX7AmoEOU0sSitnMDRoQdnBebA/bcnFMnLv
eiDkagBPHa1oENj+f/L3nelI3kNgoVkl5yBUF7HP6ziFNSXDlvshRRvLNCn9cDIs
0+46bUTL9wwFcRNcYur+BaFRXV1NEvM0VInnxlDzXcwGrinwTN9tMpbi2oRFzrqR
hj/nAEFBOL7dtyFEdVcCa0WuFBCrft8SjWkYmKkmw4TlcySRLYCptjPVoeKVn0kd
U1IoC6tFGyCqPXSqx+guXed2VofXj/lW048stoaZWi3sVVqbg7GxxKR9s/hm7VAL
KWchv1+6tpPZZFytxSAtRWRurdwtvHU/QfiYM07nlYdJ4A1gkqDuL2u7v7yP8Uts
0djnGe5Ez+scRbbIAyj3IJb0QnmOtGsZEHqqPZgUaw/VdcisyRR5zl0O7Yb9ct0v
dBSvYlFZJ9RfgSBHkj8kikMH181eIsS9B3WZd70HxZjTcF6FfAaRjCUSosVeatqG
IuSB5m2hlt5F9MyLveGEcLJbHEUCVzK4qBhzNf7E5vGpx6dfAjFMBUcmaSpVXiJm
VtOOrdLlduU1Umqqi+b+rLBSBbP/OK7HqCHEV/xkOIA9oN9VR81OTv0Zp4KDxB9J
S07TZmwROpU5RFDbTlCfo91euKVz2pJJ5BCzCgDRU2vZyKk8yL945NwLYp17v5ET
x7fh0IY+eJ3kAIyhETgCTNqkURkJmQpjiQBLmq1I59pjCtBv8oTziedBYrPdsjBX
4M319zm0OE4oCpQ02Q0Cdg9a1PVWfaLk9NnkMawWaMP4ekmcmx3WgJDdnNyZtMKQ
SnLIgNIFEXf1iF8e9FpV5Q4IckE2Iyfabb52f4xeIg0/X3c5kgM06ootDHTwkkil
2DBTFxPO/meWxu93WoeQ6/1W4B6GNLAgmvtKgGT56aJciSfVayu8vlactRwmbaZi
VKMMd4U8Kri/QVMjSovlo/k3pQfw+Z+0CZNcKxF7a3pLOmKlwnR/GXEDRpG/ShSt
UPu6K+Z/WCoXc2aQfEXhyQUH5C4hfC4JiyITqWpMZ0m+WtA2xavhbgHiy+q+7hxO
GijM4aZIhpgL3O4PbeKSUJH4R/+E1zOxWOMQ715q4O4hWgw7CUriKp3YCBRmMHs8
ReQfxVCI5X6HRgBjv2u6Zhp521ZBxqWa36+dVRuccHHIOv4ojx36Uz/yxTaKR+JG
70wXNRhWznfY/W/X1mweWvet0DaOPRaPqlqxV3OfYpdyKbJSzEITARmGJWYN1/Pu
VA3x1gfNlen/+MegFoRWpIQm2QNfa0bGGg/ubLiN/gKLcE0cI0hZ+kL3t4cJo+72
+jOMs8POU1ybw2tWoOBpvFhaXpVy8dh1HKsZwlxEF2YUebAEEi75KgiX44vLCoTL
y2OSgT9fTDvA6OQeAD/wLqXUkojwxiBvpaJW41S8f3OHcKHy4fUKHyRqNubbehsk
3i9y2/qmeprfe48B3tZvy1SZp4vub1Inpd8Wu74pc+uAiYPzqipcOpJYCM3eIskq
k/Vx2Bvsf2wy5NiTII+JqAurgCE8a7bWsuJSZckWhshm1NGq18nEPh9QyoNIvJ+I
1UdA7pW9KfHnPlkIBv3LI5DnFROTTPgE5rsIl8aoD4feOcVG3Tv6DX4mlUyPic4d
jdv+/GNqHQx1cYlaD/SesMCiyAPptv8VAwPVEGikkquSATHfx6JrPqzS8ucR1OHN
12JhHW/30Pp1gdQzwJh6DZJXmjn6xcMPCxxeqLG7oZ39oStJfbxfK3bsRQm5y2w/
Na+9cwDSD0qT0jhoINYDUFykIq9pKbES+f124O9+L1y6vja38OskqAEycm+9kj6b
QbjlxNxT0LWbzFJKkTu1/yowMBW5tJ5+NwqCK9xJdXZXSUO3c8HSxZ28HIU8uvSH
CG96dGJijr7J3AGpE7wxdnhS4fiPhDt/67QS3d+BfVyafdz375e7/oyuR1FzAT5k
GPLtRV/mlSB9Jaj7408/UJxon5dB9gFwVwesgZk/BCKK2WWN6A6rA7548BRDCtxE
cEvoo1pClKLHKTtLC830BkfgkyLzvS74j+/f7nvcJD+78jWFweUQtmT8Wt29vytJ
EYhhrM6jjTyBFvaa+I1VwFALKhyhWWdAox1FhvrUr3X6mS0qh3SWW4Raw5SYwE7W
GoJjvNbsMXKRrizzPlDQXvgrvOtxO9NCg1kb9Wmm4PFcvrokRIp4utdupfTigN0+
fWgKzJjTimCBwRyYilsrDvQX6ICIgPEOo1yWG7O9RNFJ54QDIk67etuTZ3+kUNod
7ggf/FV36EmZDeubpb5q8lH7QifDlY+X20tq3ql7V2ZC5BbScBq4n2i6BylPOJ69
vfqr9tgiqyqkktee7bsENTQ2vfqrHvh8tpVy2mf+b5dMIsZcLDZQTbkb7rOMNYXc
0mKIeSWXDQY7u9FUeNbX4dZ+u3U2EoGODNQvDkOY3hPpR5JWooVO2Tk1TouMWMRl
SLm7G9w/gAM0p+itYQ5bmqBfp1QYKhvXiBdU2wze4CsppGup2zl9cjez0iSV6cUL
8ln24FZrkBSeNlG7i2DuteeCBfM9OWxGPjEZnPvDl6tnW6MPZW+1f+w1XBTtXa68
ezMLhcvc6FZ57Ny4sDax3vYe4/UhtqWfWjua3tU9IE+/7csy9UlEox0CvRwibJyd
9HKxGsHmjgAG8j/Hph6YsfAC9ecXnxS1NKhf7/d3+5pz5Xjjy+0ykSNwSaCxQ6YI
ZwnFvMl+mF1V0lwNoTbIvpcbNWUo+erzGsS2++93ceLLyGaWkk/l/HKnlFso6E9H
6xCUmnLNTqq0tbt88Jqc4a1nrGIntQRqX6kjFua3kvCNztGsiigClAqY546MPcpw
c46Wg4+8ruS1TexfS4rQAtr/3hH12KCoNSh+DjinSW8t5Ti3cF5rqBMpBVp/xIjI
ggiveWdEyCnlMFsGMFrBWw7tS+8hRNQwghG3z3ruVaBTI52S2mGEB1/KFJPDDUjX
tofKIDIhL3OcBo6eIy9cLhPG0BwsBMtSd5AkxnxcFzUkeSp3rKjGgrIdIwRB4088
uwKwfTVaOBNQyX2Jw5zd+LBXq5amqmkrcKBZA30Ds+8TDVYhWMWgSFY7Op8bobOo
YtQHuf0/4GnW+oHqDKVnXiv48I+TNlEUuxJfaSYFsE2wUDA7Cw2hFOxr6Y76s6T4
d4qQeQJpN//48BLf4T/7l7alSsUUH5FGOJCSfXvXGDtCAlkk9nyxvoSi9upHjwU5
RDiGMmtZDk3eICZyHS7VujcmMN/hTB/fgTKI35phQznkRrV0GCf6Q2rk0fbfaVup
IsKgCQ58aCets2trzftTKXpGIeMD5J0mrKLV9AtxmQA8/DAIJ+0aPjXH8gVGFetI
wUj55x2oeUnFtQUvVz25K5PO0lh2dg6I2+G09Q1gesldYScXBQLG+jMtZHl64VGS
8sKrC2YRsfx7yHfGMDBNf3GXZ9pDjkMnCU6zn/nCvOh7+qgt0nmToYwhqNR0ZMPs
iEBjx0WM+kG/MsnDTPY+8xgiPSDN7VEQ6k/ksiC/XeTdyCdG/x+23vKwr922pekx
GEM3/5K7vghwuNqcwzTktO/iyvbVYJEqicKICPnvf3k+Uw8xgleFbYK8mR+0AESj
F7MIl+ulN0OCVyIgYjBCBw3fAjS0O1Zaj83F7ZkU3E9G7qtclgw/hKhoukH3zh20
vvNJpyaqGXZKN1ybMnsIZiG1PmVKPgGsfODtysOE6S1IJdGmBUO5O5m2z6MYdCHC
dx0NsgZmJPHte4kXVg8yxs8SMF3HJJGLKrLWQ0lREGNFezqD9VY/KhNojGmCndWF
fJDv3hrCNmKqrlhRExt38KOx/AawHdO2IX2sVcGcZWhXmF+FHQe1hr4vTmrWSBo9
Uu7IbUjVoKQUMBQ7IKqG2siTf62eWCIf66cCgi8FwDKllnSXIewerXsQ6v4PbKxv
2amxL9sUV/h8DeCZP76JySxLgTAdEza0Krq3vRE7ay5dw6aAGXEojQCz4IJFlAde
DAiiZ9FVeRoMd7D0/HUsdavlWxsFyQ6gS2PJvbzjg/VYMIpRzoaFCR/Z3wDiE4Fm
vDB25XtzLwQNosmG8F5ATABxyeZOdT5fkzy6mTjOxKqory2vZysZyzrM9QhH8wP7
RHHRVfLQVcqvX/sKwYGuhxKIn0joyM03kHez6Al+Cgi0D2CFCNWo7wNEJK53CGDQ
UlmILdQK/zdc5gnPot8oxaI1bTPPAZ9CwFOWzzxMi1oUmIBwHgfffiXF6edqJZ09
HXxhHVeyx/hUpvhCl1qE0xbULX5ZJK1ywcohad/2EftxFmdUkQGsBjr+RQgVDjES
LDocxwsoh4vgExB8Kqvlb5eT7boiKaU4hfxFKMEPckG5x3Q6vJtYjpLthxl0d54T
c/SQmFsR5UJWPVZxtB3A7O+A3c6MxdMl14vA9LQa1SWQib4hl3OInB1fajw5YMPi
Y8KZdQQk653kvXp6rDiyd4xM9RZy/3au14Vz+VwrPIaApYgmJ8Un2XZa3Qaasn3E
8kK7fGQkrYXvmdnxRPPolqwA43qvkagxYWWlIYru8XxGx869/EPYRvMXMu7TuTRW
U/1agQaCoofQHBdQJLnp6pBFief902AzWdetWkKxlegtY7kInUG3BvanulisWfUl
8InKTSj+rl27Zp0i9iwhnM5CvQ93FWJyT536wL5w9KBIy0rXspRrbChGqCnOPdib
AYP9z0Mvi0vCDy/YuKyYWtu6aiyJYJ1iKtemIyCwNg//pZ3IZ6NW2OEPWS+SVgQQ
hYh1CxESVQOtOdXwm98WC7KUBu1zMs4cGXOLKFox71V/JHk2XgLyjEb6K+7BnIA+
PC0LmkorPoQv/LA430tuSHGGjbMV+GN5UiBhjezMMeDdffz9FsDPUyuDsEx+n9U2
BAw0H6Q9jcUyjqqES8Jc0RioNKNWnSQ7g0TdsLK1co7nHkQt8B1QPqm1mSFNpvvx
9EZOot3J00l+pE+Q+hXrxz9BclNppgZjaMcnWNTmzF87IP2bd4p/ntBb+1jDSe3R
4qqIg6mnu3ckwDIQvqK55qOl2Ycbq5DuJEavmT/7a4+w+L7PzA59T7PF7BRMyntm
Cjgf83e77Snor36Sw+3/C52tQ0rpNZEdhJsTL1FTzC9R0rgDfOSxMsoQbghy93fz
BeGY6A1KfPkX95LsZy902N2mZnGkF8bSYnsqD1+VtPpb9cGCs9sd5sWMydA2mUhq
7D1Xaq5LUhPoFaoQpIcxccCQmkekeoxl0rAp9y7oimpZGs1QahDlIoSeCm4fIR5F
gu1krxnMpqpynDsqeTMtHM6Ro8najuYH9inZ0UaxJjdyOT5PSATHSb1kZOmpTKkv
pscbN+vhbPYVYrBH9HgfjcPcdr0U7EdU2Kya29BI4CI67wZJNHxcZWBKTfrnyUHU
EU54fdDe0ELAlVMrb3nDINarNgU6gfjll9MCWlOj9NwMV9kAfxKfcOlFwTNeOcGQ
M1GiBhfQrWcgKlZ9oGlIy30T4tA86jNeYGyrnN3peSbbHU6BCQHc5Um9U1XD3ybZ
z2jCLXJ+sVynufIiSgNt+G8RNdhb7336icnUnpxlkUtcWSVY5RhikBvy2lUgdIq1
Wa7Vb++Q7VomnDd187swAiN3eaY+9HSqV9kgqAYAc2DQRul00GTvqsvbWEVWAq/Q
Zb2Ep0ED4XhdLkNO0Lde0BF9sYYLCihXt/pS2m0nPbrbl4Jiu91qESs1v6D9O6WN
bCfG5XdLf/qnb1inAbg64Ir5NmNEcBypB1SIGInmKFQaHHUNE41zUSLkScQiR25i
ltyxAm9qx+lscRlLoNBIxH6iH1eG4WxpUVqAE5uAkoG4B+1obiPwM8Wd3FE0Q8BA
hbdmbxN2acW50aVrql+tHrXPELR79XScOkf58p1str6cMzXDTxYNjkx4PPZU7+M9
edWJDxr+C32ed2+R/eXyv2wqyXN1Du8HAbFUcxFrsSzGpiwjlmO0UKEIacHrjRPb
ilRc1rPb7npf1BVGtLFzm7WM8+rTTYpB5L2DnxOxLNaX1XHwe3q6Wu8N9e33EKr0
R6S1G7GJekAv8cRxtNVvPj8oT/MwVkYLStRjKfjfnBAlckE7I7XcUWrRccRcoIfv
3RnKuPA8y67Uyona/ZB39LJztLOeR1T07D/akU8B5pZOUIic11uyo1QtKwBl6SC4
zXYa9fcpwWeziPBLIHEYthFxLP0ePT0ohYKWFP5I1zQzMYm0wl94cXFw+rthQIv4
ZzesZOfKd3Vw3jsZIei/hayuip5Mh0URlcD+i0RFluRaS83aj78e5rzxDHu5U6yv
bPVyhnRh2PmI3Z3jmisujWXY196YqZSDKtf8PgrzJC1vU5g071LSJuY4P+ldQ2z5
QBytF6PHvvUQKyJVBd0GiMRaiJejlCybwJMfTBgtIUG10dROXNtf9MuCFaurPeRx
lgzgFUgZGLJPuJgV+PxM3sbJExjgj13dbdHlWfpHRp+2nUQkKLGz5XzYZIyOqFmJ
GUUI7NcnAxkqBFPnFllTJ6BsIfpHyn4OzCYgQWQv4cMZ34LdhAq2r1d7zINQA5oi
SlY6YGHRLFaPnbipvFIUxMJTzaTWEBwjL5ZhApbxydLDmaGnCr1FEZsNmoCRV+vV
G6ojnYsJR3mZwNS0Q44BwL3s08eXHELhrCHyTg4u9oCu35oJTsC0YvrJnkzX4a3W
J0GaxoJLLXhIMTLCIcPBPh5Mye8a5x5GmhgcItDBANR6jpMhE+rrHNgGXaFZ8oha
/EJdw4IIsQUQNA8RhpdMCs9IEmgzL2VHVaQISl/yQLLdTmjV93nvLax+yUsf13zn
HSlFw0esbQEGCc139wUcIjAtU19B3kj2GABy/IRKkb4NmhnaZIFlF/v1hq/TxhG8
BDfPhVrJunMUkoqNoyZfkisMhfN3vg7SMHsA82JGoknwRqHWsqW6UDT0YE6wsJti
Vg6sDTzcBpv6HVp2kpszQ7YpOQZirejKorQwoiqcFDfRDTVXCc5i7uTMF2hzKDzF
qWqN2Q0g+N2s1EMijYuWZU6aT69br96WtQz4j1GxzR8ZOipkwiI1v866V0ozLGbB
brncIWIGeT8vSSwO1T3vzPASB41mFHPE6WykUZnLa0iOnFHXBY+lWZBTIhnFM0cj
KTSZykhIZUIeiACbb9DkuLeIORg4qI1nViTIhbPhH0E1MEJsBljhxPyWWfb/Js0H
NOJ51aaJzT4z0/FK/qCalH1f6SNYLPTUzwjy0AMq6H6ZTS6E6dnvdJ9YZgcICAYw
iAXIpXOtVfyh8dyGfrFlAK0BQAGoYlJL8d4qVPyZ61L3rCyKKmYgwXUg+o3YuCGZ
uI049UkeKNQORcnXnGuuNaaLeBWKj40n/Pa0nBcOravcjiDYVDKcmdoHZX0//Xqn
qQLfUx6glX1KJds74MYI9f5TzFkVM5qTQdrknrr2iesH8AcX7zE9FEpw1TIitVk7
Ld+RsW8nURLbLaSunCMh3vPcpCFpjv01CdR+34QBm2LjfkJQYIrxDkNRS53uvdDU
5FsqBeuqV1jjwylNMEc2HqJPzkrKRwfVmRM3nduutpfLyfmBA6h0WPghJKLSZ5Db
4zbukXdh/6a3cqbKPi9Srrk1rITk3UTI/wC/vSDi/NajVvMFaCBOtcl3iPk5auWV
MwK47jbnKMf5tjaHe18Rtfz01K1yAiYCnp0pPo3ekI2tgMzPUZqJHwKpkQQOzA4p
qVbfIQiB9fgMXq8cxFdLZs50/vyRzvrk7qPlQ9OBFt2bXLf7G6AxPMai2BGqseyT
Aap1V3Q8VMhvr4hww7U8voEVg2vNNiXBE/fGlEg5jACA+mRZGyQSE2FvE2sEZrGp
hjs5O5SmOFVe19fvvpb5psvDGwZnvDVOEHp8oqNJskhmxTsHX3JVvYSn3JsX76L/
2/AcUwNKzpqlyHsBSKgbSeO/7sth4j9vclky8K/LnF41/HOnHSl9gz1DaQbNWDxn
H1r3Siger8TE3Io+Lfl3G62Cl/2auAR1augdsAalL6oJTowxFWOZSgO5EK6T6FSZ
/SfF/8aTFnRIuIqkOLSCrMAyZrsrYura/2dgM6hocwU+FHyjVAqL6hTLg1iClo6R
ETG+VUItjf9ap+xiNFZVJ0UY5WqaayssWAh/+uVwFoEAFE0l8HNbNy1kljq7PmDY
sD9WHBjMTGqwc38vfIuPqjTcydTtVblYQ41ONYBqCziyUarZ+O7r91jp2fz0OARq
iab4Ergf5JMwPK49Y7wEq2T7jEgYBrRaT7PiuOdChEtXFPsqq/rtFbMOi5HU5FSb
gAsW2qZkmfTHRdfb1XuY76T5ebMPMnt9eozYPNAorP5z5vJ5zKEy3LBLMyKlc1Zg
qVB83GinxQsC7fe0rqOhyLj1Jw3SP7IIl+fmJ1BXb7/2Qsa0YVXj2aA0xEusoUE5
/D510p7QHrxVFhVJmRNeoUjz70fUO8Co6ZF0iJEgF2qXV3vXyvm6McI8ED0+2ZfP
qesKMb3j37gfCQLK5anyjU2yJyFH/GMO5HGnJSF0TYwKt7arG5x6BQNBUJTJKN6O
ZP6OD77Y7dVzqRW6zDGf2ReEqNFAYQYGyHwp/wQGexgYZColwn3VlBaW6O/eGNaq
RwlVpYt1DJp77EZ6F9P9MbL86t7bLxMau6EcbNGBk1ylIHr8azSQ61ctS+Lo08IH
QNKOe/yt3oZdJDJEB8oWFC2nhGjflVg3eONLG2Ag5GrKxX+OuxSd4oJGccfPgmAJ
kkIoFOXp52wCCOrFjxi1+Ss4Wk0Uls54+cq7V7l6l5Y9ETcMTgGrwHN5wORkdFMn
5G9+faN3jmHEALYDGq7x5ddqdmgbbknZbjN5C87WSpdnfyovM3XQuJRhw55I9lNh
46erFIJc96c5UyHaxxYn1Zo6dOlkRQ4kBeDcvfebYjEI8y1c0P1eYwWba/55CRvu
y2Df/8qk/3Un2q89+BoKnGfQ+PTDrcsGKikUeT3MQDkGAOnmybehbwP5miEgykue
TCF8es8DMm8wIvygqEBVCSJ/6HJ0olQypyax5CZIGMODGo3OkATKPdhAeNwlJ4Uh
+fDLr/ad1PJGv+lSV6Fuu5OyGyrmnT/p2Vr8zKEw9WUKQCz76B9xCuMkzRIlo8yG
jAercqF+gd2jhK336aQNAxNXHzaP8OfsdjRmFSDVs4jhPUx85PFOv+Wx7iH+s/uS
+ojWIFb2iby7Hp9KuTt3fJqM9Cp1cwZvivVeRfdY/xf086cYw34/Cj8ai++60TmC
E+Rc7iAAWewOphG9PFDwKWk7ST180GdKnO0B1n4B/2w9vE7canupXUXpEBUGo+23
ZTAZBL2PNOAeFy4jloIvp5V1I/1Oxo4T5nEFs1ISin9bSLNG9CvH4/SokjgjuydR
OSK5JaUC1HrNEMbaFtxXkV4ZIIqbfvVRrHRacwUIM5donPqlnqZOwLL1qlUqkBdw
ZWe1AP8CjXbKWD8QigZKo6N1QjYHQRgdhrxjuo0lkdxdueQT9hpGuEtnMgWemVMU
x9YR3ZMRyI0jxFEIGAiBOhBf68i3DviR2QnBCYeWmA/yJRb7UVMuXiTA1b2o2a9b
4MwEMP0YWE0Tqc4+xCLeV3o9DvqzHEYnBums2DszcpK7LZFF97awhLTAJG4GleKl
aZk4++zG4mdpecLDO1OIvYdzqPVuJyJlx3V8OU6cNGZW5q/7ShC5eOm1m8X3ObTL
U2QFneRGHcmlyi+xpwHY6PlWummzlyuKG2XrFDhxgdLj4isp/l3/3uGBopr8d0HG
f8iNBTWCE1NVflvlFx/LtP9Fym8FIvhqfEjXJ1uOkPKh9xjpgxBKsDn23vQ88nUx
/tPo7zJuZGFObqUusZ/F9aLQqheVZPdFemM5K6FiRl8ymkZSZm/L638mo3iFxVxx
kUzM30hc+93/BK0ZSOAQzXIVC4m5L/23XBU0eWwa9lPmWpjgG/ulwa2LpqbQSIJu
7pcz9yJxcjuNWMTYZv3pZIQ5FdOQCFgYUhDkqrZkL4/N59yR8ZyGMcnR6y7qv5Yw
7c7Xw5dIzp9nfIX9P7HBU51RSBBMRRBvycPKqgvCIaSpncbQjXa+dst4MTTu3oDc
RcLgSshKnb1KzmB6R+haoi6ROW0jb4plKzIPU0lj8hS6lb63qMiRg58Acy5KKh8r
Si/uHoijApwJEf4BFI0wWyG5OKRyCAdMc3OXjTT6yxJ9zUoqcpD6BadzNy/zlf0b
ZJbBx/Zx1u8lqEw2OeyfOQftpzH3E7KYdGXOdiJkFh+eDCL+cvccaFZI3WWbTf08
SFxsZsOaAAHUBiv9YxCxzS/RKg9vl6LmgN3yvufHT+nBh6KIYg4Rt3xZgq53ZxRN
LdnpPAwtashk5w7dojllUE/S00dIoAC321vHLpPvkvs9ky7eqq2luPTb6JtRl3cO
SGrYNM0YdldGujwA0gTKF2eM2ZpUzJ+7TRg/gy0df5Tg5vAn9NFhw7C5pXKzs9GZ
qH4HnT1HB6PdyjvIo8oof9HZoGs5pe66mn0YLkhp5tImzJHhOw/N/pinJcGQfuS9
VdbjtOyOvJxhkJgk7xslDvTDnvqg/9233s+drzOljzTTLOIGiJFshtUsdrurv1Np
XscWRmhHgZ2DBLXasVApVvIGS43bSwVQNnZUUouDNTDzqqrrzuCpbYntglLmhZWH
sAP3VM4aEIbVZmw7+68OAeXgOocRabZm9qh0Ky7+n+46UAA+OBahi72ekSylSmyd
ajNMgN6LqRqOMBSp2tDeXbD/Wpm5Xuv/rw4Eu9+vNWvBVt5YXCB+4vcbr79bx6xJ
m4kI3BYfK1p2iATTqCWgeLWGiJwlH80cJcysIYceLKTq5Jy+gkaPdO3gHpDR82f4
cQE40/+5663Hpo4XDFhnYJon4i+Rp3ZfOcJVKsv8DoKfUlDLOCDBpy4wguW/SkuS
z5z22qcCT+9mlTLAhEQNGj21OVcZM1h57DHLZA8SCxHmjvzhCeyMBO/h4cgDjeQ/
tpo71gHVfsy3euuZEsLsI52tx4pWTM+uyzHm1j9FC/EhhkiYbBcqjtEO5I8Cyg0r
C3SjIZVPbC/JSUIuOE1T02wDC3vhi9nwxP/F4zJGQLyMCeq5yAeS/YkNqsSyWSPA
bLcMM295r4tF7wQKC2yLbf0S/pwKtgZ0V/yNof7RXCuz9p3IoHUrSvtj8LnYCHYX
NU1zgYqOlFcD3BiPiQgp1RRt2Nl6pzMZGb5mwt6YWFMdZPXP6uYmGu2SfNLliLwT
HgmKqPEEE8L/+tJXcjqHYlmbW2EDYQwF6Sni8TxWiCBjz4nTsYPnw0mLO+/zscos
4Xp7e/vZs5LyhDIcnRp/FIDiLYY73CYAdSUYyqu+gruA/7pT1BHQ3Fg4i8oI9Igh
83DIKDYF1HE6jZfAZAqhT6ifKQbVW/NkNID4B+Bf1heNHWR7tNO8ECHw9LGsRVhJ
3LfYs8TSGVIZdlsdJUkAQu4VzLdTZl8XzCnRyfquPkXYnzzDRRlmCn+5iQdHMy5Q
7T1gt4DKn+rjDw4d+4CMtoIe4maZSFs2FG3FmNTuhN9VmckHtJOCYfCxI53znEVs
zm6MyyqcScNS33sL9LjYJabV6wfqkQBuS+PwlKcFhUff4rxmzWUPRtnW9qxhKC6z
W5qsRBwfWJKgv0ABsQ4KeeyJcxoAhbyqmleSUd5F0H0sfmmVI7GM9Y6VJdKnePwi
wBkW2JxuZ0RAy3ZID6gixmvRyAYB6jGtzpTC1bd7cnK8eiPgfUYJHh8fXof33oPg
pLE6xn2R9+/QiIJhBoHX422MCaCpV7kNojbKs2IPZjYUYbPjLq4lGcG68K2nSvio
amkNCrnbKRwFYxez/JjExRRjQiJnNdu6AS3qeuxuxo1aFnMy8JuKy9LFNKgwgl4m
KfvoXimA0D4+/b+W87+ZSrQukmKSbQy98y0B9zOtmJK42jYKmILqrhT6rapfYBpa
aIbROpHE8fXsiVrUYUy3eh/VXCauHpCX8vfEPtCdoN7TTqeULdTTiHcapLh6P/A/
lfeneQSHYTA66vsmOkYZxqyeUVNK/grs5pIowR79sVs4+TfEJTsRcl2SlZIDu4n9
pGKlR0O14x53KDJk2PRLImtV/iTwBjeRu5qOn46Gw5fKX9LoUpggMr+Htetf+/n+
0oxhGU3oqHhIa873+plsUyJdfLPojd0+NJdYy5x4KLUp5qNiRkAYreUTmBaUnmTU
8tqeQH0itdf/VctdLDGpPT/qzyZJNFVMxVhSl3ABw5IJBt/uanjYoN/0ISMqsFY8
b+5TtMyXRoO7AhYZfVLTKszTYmYP4YcmdvkJCt6ZZjZSNHTPlv5mhy48ZVPiwVuI
290NHx3pMWlafON8eUGTg80eNCIskERAbzrmZGifGWpEAT+LjSBAhRwAFlBgOqgO
AfNhW4oWgcoOzQTpun0JUS1bvrpE2B8kRcsXIs1emBuLgwyxIo7qVvi3Dd8+0lxa
kIi+BpJGkJ7LGlc1CAd8XJqbJ3w+fUoEXt0sM/gK2b6klxGXJtbg/sKOy+YEK9yj
lnQ318nxPvrxjhKB/BOyjP3Y7KLPYW+26uADhvQLbXjlHCl9YbDdI+sAMpKHOPQq
gmQRkIfVYatGRNse2AxpxFWk9tWd/dxDKlmBZjmLZqzL0ZaZK3M01nvLmg8h25dN
nzsf7ngmUp3qQLUL1rc+2kK9qovb243o/IiRZ0AGk2/kBsdgfCC8MGf3L5xibeUn
b38eI5aPP9/miEBLSwowiBc3yki41GbV7wZD2jVd/9r5XbifpVhefx6sg8plQY2p
jczzqLOqy7T3nRYw+OF0FefstNi04K5Gt0sZyKMymSJU2nsywEIHkrIuVPWjMyCs
e3q2pzAWjOEb8GQju5fSD6QjX+KHNeba0A2PlsvC7QqVmCstrnfE3z9Cv+7lFd3D
5TFbbyimd6Kn2jLPfkbhZUCN/q41kVhYmv1AHugw19afPCKi11z7grzOu+EDNLt8
sq1VqR/nmRt4t6/EDacuM0xQbri5TPyL4WZs2tDFCRc3+7CkZXdfhn9qbgI++/0V
/mPL5N+5ymCwVoi/PxcUM/9u54Rx6cOPL9viZCpbe9vL2ndHXXZ2Hk3hnyChA5B7
f1Uh1rY+TO4lEKf+TyEQnWi0KQOqPrg+SaxJv+lfny5sZqGxWQmw+NC0Gn35jvyk
vW4CMTW6I3M+DRxYhhBft1uy6BxLcRSKqvVa08YPgDBcwuVk6k6KQKJgsZHfUYEw
xdiQjwFh4VU1A4vSIE0eZbuGF3d//GsOt/Pxs7lMD90fYYo8FCEhxZdzT6KCtCn2
d4QAdjJPeDHlu87XvwxyTdYoe37t4xfpUIElesB0JbHavq5OXqHvpSDvnH12tuFf
B+VkvERN+8yaGmJTcbyh+IGZXk4k30oBFU9ou0n034B+QJs2psxKug18L2oj95fI
XEp8W81eh0VU7/q/k17v//MWB5ao+oDWg0vicOgyxQfd8cL7d5iBRa/phQ4ChuFl
OTHcEQZZvQJS8xfNHlcIDh2HlrMVBKFJ72rWITQp1c4ItM3P77siCIX5cQHrqdle
6XtuWy6vF4Iog0Xix70qVEcRIa5Whbu8blBEvX9QJ9DN1v5LRkS2m3aoayxOVj+p
yjDYkW2o8Tbm0ym1OWfP1N6W1DSuMAdqUGnRkn67Imqp2LQZ/nM4URCzZcFP9Cr2
B4KrAvnkvrQoQ5j7lyEGMcUNeV1zfP3WCtqI6SooxwUxEkeCyJ7S6VQpsTMnDdy3
r0025KUqfsPqGuDOu5sgPxdiT+Y2piRDBaMktLFRBWXPheCG5CqSs+W2odFdpR4P
fj2j8pvVRyp0gsWq7XbTwJJXwIzOB7m01zLUG9BL0N7R3pNbxkPx9E584hD2ocxC
iqqngc82uNimuMNCcxTfS4BFJoY4tSokH+fWmfpAxWxPAY38ysG2fXS2GzDDtIgj
Rnnrbl/5GLsu9DzJrTiz9ES7JOul5lsyUxfKTk5IY4hbajZCnxXUxGsOBwqDz1LX
NBIIKiqQSBg6FFaDieEidwiKiB6fK8Kz2dDwDbtezqO0bTMAVsQTdZRauMjmDxwl
AOq95npDLWr2a+YkT//JtZAryPFR2HUXDmyNyk1R68EMDk2pYy8njWjk4Bxjgkpj
/+osutB4y/ec6NYUKlA9H4AOVms6UHWmD3xhsQ4oNzGuCZ5uEj36Eq8Q7VZj4oG0
8MrANPCVEZwdCdXfLR1lUzkr/b0QgE5KNmBE5NKkuUSldEn8bgShBVTS2gQIHYMd
27kBxa4nPG5RKFTimqw57OAPc8UL84nHiWZBSMl93hcGL1foRJT94u/8lTyXbheH
nvbeHMSG3cW1KGkqgWLKZanE8dGYOoCVHRDFy2hMo3dmzDWbeT0YvjJvzGLGDIbF
cH0BWhgufcYi3GYboZI2ZOTZxJvelYwQeS+t4h6PyLfx6Xocmm4ntzCnbszDAmVY
TP8iya6uV1XzMRzQK0O7KnwZfBokcDuKcmmtu1tQnFRc/7idwThigt/uRKBrFKvL
u4MPuQszIoogj9eo4QsnoQrMX4x7Q9Sbu+gIj1SQvBgTeHHsiCf3QmdZCHvavH4q
rZjg8PT0dW7RqBJzLmcpTEQwQ4DQdZdrK6IuRawy1RXZYATBLQxv+OVuCQ00pRom
tDOsTpZHCaulFSRFIsKrH9tEkNrJVFr/+1Y97xzeY7L3QQ5EXxxhCowGCCt8noXm
9BYbsGGfEFiCojIkbhiYG4rh3sHCsUHX134pP8n03PfTmUii/nRCcQKIC1NxyrQQ
jeHnRca68NSfB9XQEXAHNVptL4+Zi54hNQkkZ2VzonDNkd552RLFa3jTKbaRhhWi
11B9ixeZwvZ/4oDM6DNyAmgS08p5u63qJfxkKNKRfgRu+SaZJEPkiNst50c9TAGC
ZtNLa2BfGcAPFSejYMmILtw7MOjU4D8kT4JdNNfDo9DWPVAc748ZHqeX2gP3jCsC
cuebKZd7j5WrS3fcbUllR9g15RhzXV2Y1O2nd2oQTNepycQFtnRx7DdT6mHC0WJ7
3pycfI94FGZpMTjXpP/zUt1FISKcJ2QLuReT8z+EEKUxBUpcEg9HTiiA0uKboD7N
/EJi5z6HZRzAycMqCRAYqu9DzVuaTgPiqXzvS79ut0wNKulQS2EtahZ06W32IoBH
NzU4Z7MIIa+RGM47ezmKY/yr+Oju/TpUo0ZaoJjTGC7UrPrTu/m6uOF4vs97EXfd
vs7dSM0VEmAITpe0caEJ8dEr4MDNe4kgrraUlDXJEmzbMbtfK7eJ9Nb+UgUYqhV8
6UHc1OggdHox5FaRPWWH4Rj6qjN3/RIw2y8/2JKsaEJlfTswmbnfu7JFJyGojRbw
l+G/QMItS5cr1yHg5w1cGfA2wNDbkXRJCRXvyxzS2zgDdI98OzlgMMsHBaamhix+
gnjkhx/drvOXOSTHevdpy+8qSC3kDF9Mg1RYs06o3gt5IM1E32Uo0CMiB31UjwZC
NGTv9OHHyPP8Ypne2oS8xwMYO+paX8YwIIy2qH16PF55g/7Jf9CynWH4PG8hmc4k
RTgQa8Lcu50//03PHtJc4O7MGlODGLguSQIwZjXD/udsmLqP46fz41cF7XZgkFht
u/TnqbPCKV0D1YgL1ZgMbeNvT7qR8snwvZgkjomnsa7o4oq0P/RBam0ssoxlGQGD
gudkUDwtuIRQjN+5ki8Xrg0OzjDFcrQjoB5CpFY5tMNm3rlDYHQ2dr9csIHbIaq+
Xx2jyRwIXdQFqjqRIPT1bEKpqSc7qPAQyQgS8mJngUnDP4aWy5Rx/mldL/GMB8kc
8DzhgugfDPVPJMjhqdoP0qKT2qk03H2UYn1kso5mUNzA1sib6zGgWOckAZk+UUTK
1MtqqOaUCwize3DPpJOTqdO7Z7ZLMSRS5SR/v5YZvhNGUTSEQHrov5H2Lcsh9ogh
m6iOmMiG8BVJ25tBUQSvC9LvNnutMwvpbEW58DsbS1Nw2LbX1/A1jhTlzSvft/t2
cyroiwddzURv3C/4q72E4VOcw6F2xhCxOKSNBToVflEnlTT7vOQRK4vMYz/Ktn17
QxyfzEDvl2pXvkNQMdj89u4C8YWTHadE9mAx44AM+iYp1yFyxEumfGXttJ1Y/GSj
Kf5l1QUROYmuCJE9QwM3rTSvXAxXLsLprOkbFG/uyv3fwDfjGcb8D8r8FyB5abZ/
MVRcm3/gSAx+IRgxXm84T19A8xAl910dyBHGYtN1s1YW8QKV8JN/Y6U8IvQWusGm
+Kc+gtz5wnqwpxLL4Kt7vg6fQpmqzDuzqe3vdXcj+yUVGdBQrYscYGmZ49Mbi+2D
GeTaIlfwkFYO5Nk7EDdneJRixUHXvqLj4nuNK5dVxzosbcbhhfL6xAsGkjluXbKW
CiTWJCa+mszhCmbYLRIeKEDqHBZHn/TVkdtFNFwJuEqI+pzXJhUKZ17+Mk9H3/cE
tHtdtMa2l5/cpQ/0RJGsWRuYIghwLpFo3ars2K8vzvucfQld0jHkBZpTyFUe7vZf
7n2Zee7HbcS9ElGP8ta855/iOHGklMs1Gd9ajTWTvY8gDydXIbH9ovXJzNDzYXED
hfi1cI/6ziHw6W95AjLS1xjNbO9h/OJGqJpIc3tteCN2oczD9lZuXt1VufimPv1R
AY256h8BSiPvygSYjVROCYCM+ieOR/l0/TBc961nkEvxFSXlysLnN0sn1NgwG5BP
8i+ZkCdqM90DlSsjBIJFrROoJzbK4ibtnjYUjNzEVzSepecWZNctZpYxLSalBSfP
8Gr9lwBssa6kEturtCBKJtgR0ZiVGF1kijzanFy8RaxI+H2BNifL9OS6953on6QI
dVoiNu0fXuzHoFWThfy0cgvg3R8nlwEU50KVw9mcD9VHlIXggMJhZKKHj029xG7b
PzDUrF9MOa2GoceA5ZgFkjf0y5KjSz8jIt5mjcoWyeb/JlIRqZUQ62Bdq0tYMbGS
ZRYqsFltaUbDCZ3jLPr9GNuXx+C/827DNJ4ot9orwwj4K2GPZN3EawOH1jG2wf9l
G4PPw7ZCNgYAYMgCqZRyBIpBu1aGZkiVkWopZKvK/nTHYMHuxDwXHPHMz0LXrn8U
tbSax89V8SvAXtL3XdQkFcjANFT/Bc0hmiW6HESW+aaB8RXqZuZM//z2v9ki/itk
9RYb9ZnG0NBXpR72SGmEZBA+gg5XZ/r0lTwyDNAO4FrHtPoKejZYtldTq0cZmj/D
h7Gr+MGHGUEjjjbOZ0pbYqcJt+R2rFs/o+HGxGJ+Y4LbawYjHYucw8T2UMY4w7ic
DvVJfEOj7lDjhAHJkAs0yGKt+E+O5TbP2OyWrpzuB5ao03WnA+2/bGLtXomro6c1
nxP3B65vHJq5zVZ00iJrF8oNzCD9a03dqWqWBkRLRq9yFKN3gQSK/rygro5LxHB/
JOjU7ZbTmcz/Bawe+5A1dWghTmYH27fnYFvM3txH39p8XWTAzeo57g92YsL4ZLCd
0hWjqsWOPj6Gvj+EO5+SK7Y7KwA8BBneJm234Qdlp5krsUXoOe/CumTsCBEn6V/O
78bziqNHx4CT2Cnr5iHbOdElhSGS2onBzRG1hMQw8+qVOCnk+4bi8fUDIAJwluq+
q/jQnmqAHdbGv4NC0rVg71evTSToYtclrULmHzrl5KX4EBYfREmkO9zL9k4UNwCm
wYWpVlPmkBXzbghAQEElu3MEG6dd3Q8LxTFy0afVY5Ap0m7zJ0194PHNgPyBkdEa
akYkGZeDOCPXDQ0ZcuL1gQvEll7fttIli7rGun+cfX54cpZ+Y7DwjgnHgMNjRoNY
zg4asW53FsWHZdkFSQKL65TA7AdGqvsnpjIqGMWafMip+inAmdysEP87maZzGiNF
fbT272mEeAKukWsE9NLz8SxI+9/5tOOB8wyMw08YbP5YuiVpHeQjho6cm3PawwGx
Wz7OHl0zaXoypuxz58MsQgRWHQpsHYwvWEG5aGCVGgrWDCEHtQic0jfT8DUoENZu
Fau8E2U/Lmg48hxom/jcI+Qu5EJsScW5dbktNON0NjdLvYYlWmuVbTH1+DpFox0P
FNoDRG+uO5Dk+obPghmwl1/We2hrxEIbvq/5l9uEn9m1hib4QyhGqq8TqrMjSe3A
tXVMPfoxgDzE6gz2/xAPbF4rgQO2myFOrVqCXy9WdLDCKh3AwOgKiOCM8Sos3pY9
ffsXaCz14G7/mY3twFQQbTJ+rFQZG6D2ubUaNRDHWfq0wlPUfUK/5NiXyiCZdNTQ
zv1T6kLShsyNxpy+9Jax2muOPppmzAv8YcUDHs3kmc1yxyunenIHRsWVvTQCKfWJ
c5srPAmjWLP+MN7QhBulHnM+Eb2twAStpHGYBcac4abVTrDAO0IfoekjsqctrwXb
Bl/KSz1y7t+T9TznQVhIivrigbhh2qNbSo6W+lMCa5sRk360r3cjRVwWi0C0ijF5
3R0axPh4mKqNpzI+XYOVuL/WE9KOUIlyXrPMYTKjKkvcsaSYVkw8U3UkJl28ZbA6
wrRlt7n0yJl9DQFA4qlBYfLRDF0Tc2kZhwW7f5g9E8zuHlUWZr7AL5BJpN3y7qw1
jir+yXVNOujoAj3yWjvZWrA3fAPmqnPjvPVRX6JT1PnAh4FPrmr9vywFjObIJqyE
UUef1Ud6vKDEZfMsNc5OegcSYGo28KxLLgkxVF+r6B77/0Lxst35kvvxuXTWlXCE
D+NoQ7cNDE1OHQQscww9LTDatusKQMjajG5btLIi4zYBPc4OGMVbqQ+i3NfKSX3w
C7AjjP2fSeGHNxiUjgqIA0eM/FYDMKLWrbucv1lePcoNLTdtO9YF42BwN85NBYw2
ojxw7csklaip4WdLb5rPWV69qNAgdNTo+yBB9t1WTEPhLGoP72TnQCdxvTqStioH
BfE3Y8Y91VXPpTrbFzp3gAU90wcQgMy9Kdd2MBFv9PCXkCoyX6HpzckSPtqfEF7T
T+HK3bi8R+rxhM9CfKNtEhT+fmjq+C/SFnz9qWSRKuff9pusTr3U3AntaOMtly2D
Cdntf32DnrD2BRS+DFHN2MKR8mlIXgkYBwh7xJOLIlummDc+sWI6ikKDrgBXJumV
v4FyEKaPEU2VQOI8RlZG815kRpH9tnP6TLUBUYC4vZ/oWZyCwdmRk0qvhh+TlQNk
bU5O+ocK6RsCiIEnPo/BUPjDJgt2feKTrMQ1udDNB4oilQajDukYOcB2zEtWOReZ
c5qdwxpKHq0BgqOggnGbVje+8PWeDCljQtdA73X2eG934OJ/xHLtu5NKKS5g9wHG
PXl5x/jm7kePmkZzw0bin6KJTUbiR8spFRQ2Sdqglib2AqqasDZeVR5mqv2Z794G
AZBNON0D3nrkolg8fWr8VjiH+TFyyShd9eT+LSVNvVFSyKDjCJsTNwOWUUnpy+oh
5XJUcFrBujkTmb/TUUAvjJV1rC0TcotvKR1uqpPjsMcuiUBxC32OQFXxYJjvC3f2
9ijYroweH5UaC2Ri21bl0/ERzavrLjePZChXWgEB2G269hggF7vPu1H7dIgovn5w
00QOCpyu7R0Siq1AphJx3LlVgX3hOfuqG533YRy/x2HREGwm0B17a2Tof6iBfzDz
deD2PwP3FkpLS04TzB9ZfaZd3icUs4p545eTPW1H1P4fWHyi8QB11VcZ2QKKmgOj
+Q1beadGEoHiX35iRT5nLaGd0nhtlQ/xPOOLAF7kGIhjp9sM8Fful58vUdMyIabe
Jmdf7bF/MLVGjwYth8l1PW5nsMdFvbimwq1fjr3Ws6QTRrokeZOTEd3kgYLe+O6i
RbVee5ClVyyKNmXiSGKLVewGYePZr7c/rxZX9XjCy4xcD3AoOkC4jFi89Vf/NVhp
QrAXFbVoSJLnUhC+RdfEvKGePcVDcaObPsO+wbB3hL2hp1F9NE6YKkHKx1m+w/eX
uMWn6prLmoYvUcsNf18VIkVv5CO9C7xyxO5zHkuCxjg+owcEXs1W6ftgBZeJm8WB
FbmqnTHXiU1JI3OejwqNIUmWOqgZcfq3DkyA8VZ6wY1k4Utr6V9ufbLbnD7tYC49
pB1hOM+BmImwidBAtUobBJBAUddhLlECSS8+R03fNC7CZKusWKRmVK8AY8HpKSZY
Z4Ty50c7d7n1ir6ZYwV/MUUtIlE892VhMoqz95Pq0B0RTXkA4Xmz6ToSG9u2BT2l
DmLZyuIKvBE8euO3dQFYk3g64xgtbS3mw7fwendA44yq/cRYpuuz+DZATxXX3p3p
XpTv8eDUf+G4lwLEJZSHfrLqmZSMWw24PVnOvlqmcRpSz3ZPQzkUNyzI8X7ve5uh
93xb0IiinjkmcyDOxcz6SJIJeaFDRGRczrNqalWWJu8YMkoXBjVXyx4e5Eutof3k
vMmZnhlYCDg67HTy9QdT4AzFlA3G1V3Ji6udufkWDqXFQJH/VtFoe8ydGXsLcwjj
bxPzsSODek1pdIrNYM064YD+YB4lIaIV6BlRMD8ZIbSIFYzi3JXHNh8hJI3wKg/V
8M/6To83yni7Pinqx2yrAWAEwP9/+lmdex4HTg1HOywD5ANNDpEIQlAop3Y7WcCi
L+efU/IVogwvprS89AKDQo1GpLgUcl/Emd8IsQVTMeBXFfkohMR8zdMx15vUuTJM
Cb+DpestfDXwbvRHwld3sXdjdLHRnmk6Wow+ZLj20wa/wh9fyUL1glVT9XifhL6E
BEqTyaxzWR1pz0APrwu1q73tLLCY8f2eqrh/m2gGtewKcg3iGwCLwD9C/nxSoXNm
Jv6isX6MuaGdAiUn+4+y228rvsPNOgioGKRgmiEBzH4e16IzD/FW+3ItK2DYAg67
vwkV2m2Ztyied4TcsxtqAFzXydZPc84vj7ScntJRAuFJKupzTTKAUFb7h7Gr5Gwp
euHG/kQUgaYrAqQdzFu3/SHOYg+1QxtxTI1S4iNJWkKl9R7PQMvQtaRlZDt7R2t+
/ptGbvFfsK01wDx8zBNdWZ7BE85XMPnR8fAH9n8yTw/md3iP9e1OlVhmM8xtUtYf
tJmp2q+9IsjZtlBqH+u9Tb2fe6620J4iWpwST7quk0bdiDA1Iyw3qKBh0meVvT/Z
83GM23K8zheDs4Nfm9qTQkc9ug3wFKEKdctlL0QSFPtmBH1RxjXIgMJz9l0PE9xp
Kn2HaRJM1C5UCCvpsKnWGxgGZx6zab3P+1ySoUi8JYuC6oDY31yXnKVOwo22rVN0
PsCz/BgciDJcGeoga5q0DojylebsuBJgrlywpJGdM6lFHlFNZy59K4lr9vddTipp
UXZnKuE+K7tMVuGxuHGRwbkN2TsiBCvFSlauKO45XMEMBaFxM5zo062aNUBLJZEC
k5HdoJ+qxOYJJ1BYjx/2VZh3r17ITft/vNzTygirXC2tvtwCzx1+yzqMtAwjbFRl
LgzkOs+C9ZrugF5Ooo8sgG/3DTMxZN9SONocd11K3u0i0G8vAQa/XgzMdwDM5naF
gbNNr6Y2OAIjV2yYTKfaCd/azVfm91ORZEeg1LywaNaiDxMcOVSU3Lpe2DCVxSeE
shVx7TymhJV+U00jEdThKeZ8lCLPlVPKj6lqFMjC61Bi2HZHIws1srwzrkruktTM
o65njTz7AasPUIQ413awIpmXj4e+Q1iiBdsgpJ/7rsAqO0NlvIQQYy9E4pdjFv7d
gtSwMZBTvXWQIj64qnL25hARpMIOPzDP034zMkEDYDZOsnCbOU+ZWP6gZih/tkVK
dFnkusI9f3LYQco+wr7zxoiz6VFqrJ9FIsPv4VoBZOPdjvC4hsxgBwjyoFs5pJgf
j0lZfbjM0UWa5RW/2tg3+dK5vMiWDq6rkVQau19zoG2dQGSn4M+ai8t8Blg+VzdG
ZP9sM+2wS6qGSle5SOS3+WGmYYt4kkzFccV8UxunaXtEt6wRFx7uuwG+dpGKyK9f
PM+ooKwCK1eRXOMRvtGyg5jnc50f3UkAqaqUNpKRnzM93XPEIlnF+lTrMSpES8XP
7i4rcoLZmQCIaCe3cZLj8DFKV4/C1DsxiJ/TilLLb4xCF4pSFo9qyonCoRBTQmfy
ots3RjXkMozeK0HolO2+ihaki7gWNAlTAp4xetG2MbvkjUUP2+513xnYsm7+AZOp
Vi4g7oPi2Xd3CAX2kvc4r/bfyeVKYb6Sq4VNAyobpvS/PLJ6ctLIDAcYJ4N9u/6/
CBInCrU20DcpcwKtOoV5nEqZ9nKDMpJMLxpxOGE8PwLUunJO8TW0Cf8EMK5lP17q
TVEvzl2JJgBtDf9nh5n4AMYiOvhsIsZNXg8q1TuVw64cb88BEzNte6TGh9O2HSqf
2ZIKfneqom2sOhW2170uQNAUrzrhyfF1bwgk6YtCy3KGIGY0bb3kUr/IjacKrEGd
xUWj2l7h0apaGmf4FRT4aoStylouaTLQOvdcabhD4CdM6C9BRRR3vCAfbatbbMA6
ug95YEAGo0AAgZ+wbanQDSrsqJybPRDzgqbYw+LOy3nPeK7EdcJiHg82z20C3+Wa
eg7X7CwugoIyvrR5pxziJT596CxZGbzYVTMsJIDPl5mnqQBYbZHL4cCaDOS2vtNw
OBnoTujG14zSKv3+AlN8Xn8zKaDPjz0M01YZaz+3lRptWc3WaFC2hURQ46GyKZpo
cA9Pwg9i0hzfD6ViwBlDAC5V9Rd1VO8Oz9Mu2gqx3W15Kygvi/dsDsKMsEqDEnY8
yx/QnWJ7sCMesh1z4/tm93hatoo1uhLw0JKGtC1ID49kf71ZEzDDnq/3tUnvy8s4
8K1G/cyJUuNk6dvdkvTsLrCcrdeOIECnYGtu7UhQaHQAW3E2dEigcak+LA5s3Ycd
M0iTMTKzvsgPt+3C6QNCekTQ9yi0dZiROlQmTdSDtbYqQGJyCwBazoxb19T3IYO9
akYfMG47pjZCf8oudcPGYdb8MVPC9eBy94BpFcBXznVHc43v7gCc++Y+s3GxCdwt
x7AZHRXtyajmugdK++Rccg8vyEfAz0HFV5M3k3Nv2T+RUKFDObqeS4tWxvLRwWba
PyscnbToHbjuKPWlXJ/yn1UuLCyr2/Pgyi/C/sv0nevuIC0xXcKdn7QENjNPkMMy
+AXHOFF919MKfkwrAKm1nuvvnboilxoyHkWkv/aF8FORFjdyl+1MkfdcMBdRpi0K
I9LEcO9wzuvjngsNRZk7hTFQpumnyLd0/KLlQGDwFgjgUFMdLa2v43rId0tMrn+t
k4lLgKN+5EqjGKMf2R9pkmuMnmMnNyz0HP0rFl1n5feVu5OS++f9VObHUbDbAAID
u2HMhCclPVAnvLyITu927kh34L9NYmvF5cixkcKmAGipne/+sBT9/R7MYKtU7g1k
VAXhk7RusifV6c2RE+7x67K/oAInmOKDBftWhgG9IH9ty5oDZf36t0t5/O/tUVIR
vDtdraErES4GIJM1mDJ2sG0OTCE8ZaLz10fly41wuatno1t8KOYscQa8oj83U2dO
2e2T8r2FcTwCTG0EjHWExT+S24axJHu8AEhbXPs5rc7ntB1Z6MY1Vb9y6Z6oILCK
5RMMy8GF4IUCAKsImrRCTKVFPDMlyj60sTssoTT1BJXkRCvAepKN0t0Q+7UCtU3u
9yaNY6dlY2nFaC9QhZfYR+Y4c8dW7OMpbyyACOAXz/e8RZl7yCwL5Ikks/4yxX6C
0/pbhlAhgD+YDSF66D9NGZMtJBT8eZHsxKoLOhlDWoFjP55j1klLspvSZuJBIOqj
V0Il/dR5A0miqM+zNmITsn6OJGhNaRi8Z68Rx40tlZM7+5cK4Zv8vZVuP38iwMg+
SV1jfxFjfX4vZ5PKB/3hfNFu1xDdptnQqwJHWxYjHWx00chm8NJtalyLeco+wPsq
kD3H1FrfQRgHGMz8aJ9wh/OKs50h0J0oWdI9pUhHxbruFSN2zlhsXVxudP0O/AfL
EImROPApiZbCacQtZD/Sd4a+cLieIKQLaoAxEF+ysDXbsxKg3Z/CQ+IPgcFTlSum
lC5viJJcaV1y6etoOHuZuToPUZxp2sTlmrj2JulGyqVb7KOvjSi+PcbRSv8gRgKT
jCXJ9fJg2NlxyYUvL57U6BTnHv0IEV6XYtCLFZvjc4WHEEFpWlakDSbAO3rO2vCw
k8rZgCqXN64pj1FqEc+Tp6gn5a6g54pHGblciy6SWFxQ+0qj+uKCKiAPrD3sLcQA
OHtlDd603fxAHgAfCXlHVzDlRL8rmLjJqOQ1blXtT2g9C8T4EvJVWU2Glb6g2f0r
QduPOIHFW6znA3xdBUmKYOzpOm0xEOCwnvqMY2w6bqMkpAg67FJOp2RiV7/e9BEn
xc2HqqEf50Z1zfMMLo6alv88p0d5iNkj59OJKkfOlRHzY4mDhRDhmPUavDe08dWu
f0V9r2JWzYXl+nWdM9edefVO4BY0lFjVwRGr7MN4eJq/NUbRmHUpG2i96yvnqpjk
VIJqaK9nxXR2bXMrPcu0h72un6X0zWc429AydEbK1CgqgHLvuk7oZQhbicRhTmZf
3oOBdT4PxxfMyIG9ISd0DzMsejuHLoDGAw0C9YZaa84jHcTT8T1r/IAV2rVSdsen
QPfXu1CGop1vGbl5JPPOJKnRoPAjPM3EKgfbp5LDhGXzge6dQ7IkB3rBBfD4xj8E
Vi7eDgOvFg8GvAq1+29zUXC4j3ygVbCJGYIAr/qKQWqPIDttknLVcpuo2O3sQTZ+
VF0DuB7gIp2YB8Y0sKFY6ptaO8SdLCwhuAI3KlcIgwqcXFMSU2BHollqbV54gCyl
zw4tiLK7QJ4B2O+f4nFFrz9z+YBEb5ui3TLm7NBgRFGKiGTMfEUdR11/2xayIlqX
LaD6UiqVxwxKKFaSA5+m3LoSpO3wnkT8nBNVquQSsdY1Ls6AyqR1uHMMxLl/S10r
o7SCqlENq8wZLI0NQwlKQZ8DYlrKXLtTs5mWzyB0HIjKPBYPDUjF6d9Ru9qdH/u5
6Vtt1g+yugj4Eh525PkjUh52thRkFCi86Xo0avQpPsFZbXwr7z9lFOZXb39sxFHS
iFUBL+G3La86AIb4ktup4NwQDdDU1ZBE8J+yCY2drWpm+aVPtNtS1sJ+uMpZW6y5
bvZGpbhf+l4xvEXIzao74qN+bDM1QvIloZCWEzXcJH5UKz+02xdrVJ/zC5wTQ4fU
w4yWWaDckr5IDFMq7F4N057ko9ifqXj5Ua741wc2SZClehLIlXaVB/rvopXVnb6A
T0F/MQizEENlprpWeabDifZdvBKmQIWLfctj8p51oXJiPscCbEUUKWaoNap8kyv2
/uJsuO4AkWn7dgDvJ64B4T/tx5rzkSojHFBMe2q804Of7ZuIVvkdDsnxjG0jag9c
Ir0CjUTOzArT6NCD2fbiHqoZfnoJTF5HGCDSrebUwl2h5kc8nLw99jkwfLZgrnwq
Jkx0VQ53Sy7e7scmIOznmACKVd9b09tBg1RDXx40mmpLiPcjx/sSjHJZmnuG08SR
4OMoRpqrXMGDiUoTnziRZIpLetIQqIbs0Rr70nD3yjsMG15D8VjqYi4Lxh0k2VVO
Sw5uRts5lYcIySi4KvjwPFe2uF1ZkTIteVIJudwm3rMWEB25EHxGVQpENjk0HgbQ
/1NNy8KM3F7gOP3PAgcxTBFhjd4bLqkgEo0a53eDQcs3eW/ppcEZc+ygB9xne2ig
iYu2Ye1PJPd0NZ4dlZrHKQxcN2pp0ws61PVpsm1EbGJvjYV1Ob1Z9jy8YgtXLU59
IjGQ1pexpa0+/ogTqw3CLiOC4aJAT796FxBmr/1xsoHW8A4ZXHXjJ6q7mFnNaU36
OVJI4uVbnJaqrzpPyV42Abj7Co94O3twCWoZF/Fo7AZZPGK/BlEYX8Di3qSRmLkF
Ug7r7ltQmSNkUVu0xXsW7r9nsfIPbRehjS/wsqQTJqSTX7+6FWaVHXrLLSuwR3NZ
4NX9RJo5ltyG9cfBf+4kcSfAMyKMOSoh7+tFBHoF9r2zTj4ml7rFk6Vlfqs5sLXr
9nt1n6DbEepuFa08BcQrt2gWZ2QFom/BsLkgQqNXqIHFqerUpVPtTsCvdR3sWYcp
yNQxHDDUc7Cml1Ibc4hKvAKPWai+oBIpisZs1s1zUmAvVIFXb9U50wETgPtSAoJF
27Z5vNPUDsWXyUn8GNEJ8SdbmQNUVeosaDIJqlikvCB9qCudIVoUlEFr/rlgz2hp
KpcrxiXMnebY9r31mP2a+inncCtxEDrEf4OZdXAUDoeET3rzUXjxtRTR7H1oZp4R
qgb+eOANjo50fzl9S0l1jbfTbEUZsQkOj2RvSboNghBW1DOWnqwRhOANXb6q4XiB
fw3XTgY3wNuY9dnoB7rQNQ27zqhN794WnuBiC3Etp+YRhDMADVv7gLMLtyZBVqAI
tt6PpHGegUO7JCbi+0xQfVlYyp7q1o7HSemmj/awyHYhizMoaeiAwJI3XQHrTR9I
ViXFghP1CSfx6HF70o3c/RHLwEsrfcDEXDtzn3Ax956osZX0SLTNItwrpA9KeCpD
AJfMTHwI2In+BJi8s0LOrROrpkXt9jKASYl9VNAMftDXnp7oUjHbh3fA3zsEtNRQ
qQUkreoMjHv28Bn3Ab9c3GfgO/ICPlwoB07C3rzBa6nesIWEBhBV5OkVzhyCpuPK
qvmympmhiSFKz0mlt/QyZ8HixYKjT9KKC6kMFqD2ufO3/E1orXaKneGmtt6f+nhk
TB6BQ8Jz0cdu1IEZ0H7wnCMaiey7SgvoRY1/WokTnpzmhJJgy51wdBuRtmRTjMfa
7Blgut35G2m8aTHdRrvqMY13J+4YUeybzJ4nSGUGGyD9SxbPdRQLoXBwzz9d+Zem
cuuNXwQ2Y4qyJgXQwJ49aUSQy1GqtxjFRtV8/7M5/dSqV0YCrJf1ZjdxNm24OODQ
zZQ5Ch8DtI16OQBK18g+dux17uX5Y3bJujPnqV+yz/ssY4xriDw4KjqRATste025
sc3nQbrBWuDUPCjYhJw+p9d7+2LBcV3OglYgYUKcDTECTXQjr1q+0KZPt6yJyw31
dtnp52cqfRrtHASbv8SUepS/09xaVt2HjeRbhjMwb73a98LzpzTt4JqxF9ZGEU4q
5Y8qet/1TTiL+uZ7sXow9LFIdbJtiOhJaoEGH7S1C19NcdBziSgKs9yQstsKo98o
7a/zk0mzeUbBOKgyqOw/eVru0seeplzbefodgbrL3iDZGCvEmRm/RAHLo1h+aqOl
Jt/bxuofQUcrLUmaHrHbKphQ/SpGfEPvLgNOTzlbH/4QqHSVtTqOyN0lIzmAOH6m
ksdM6VFTO54b22XMoRcytuLoyfbp4GAnG4+aSrM/xx8vWUTTRfZWSKIWXmMWHnCf
/BL4/c4s6/yusKHqKpg5IUJiIwFbVrL3GCvcBvPTHgtbrVRG7IndztOw22Vs6Qph
HhKbQjyu4wJMxBkhv1YUVdo6ENxL/2QoMTjxlgyJ5CJ0cYFKvhRcy2Le+VcsCXFw
FMd5WGmVM3KLtUTAPPUdByQ6qAk3QN32weWom8dhOsKRC1CoViEYT5e5C/4SE0SM
XTIxUNDK3A76Qq1WYbc+hJOz0lySaahxI3ftQGC2GoiYMnOp2Oaz+7fQ2Y2pwLyk
bkn/SpETWNr9nwYf4HtOLCcJo8kLY3371zuUk8TYg5EqpDvMr/d2KN/nbn2jw7I2
gRyuw4qAuqzUFkSFG6JSSB+PV/ebivZSgDk91988D/eO07d651jvRVW1l/5tfsJ/
CZkgJS5iQSd65hPP+FoU4kzUy0V3Kwp40MPIT2vYjRHvmwkyeNAe40do6CzVtwjm
+nq4dzrfpnhRpXqHCV5kTDwfiQRXjLCMsFsEd1yeNN9ehhzjbnfn7eoQx9V9fFkW
rVz9f5CZXddOz5ithqapg2sK0C4t2aBV2d1CreSeL+tdxQIdUjag+T00v3g05xJs
KHco3SyoV37j7Pm0hFXj1GGAYOT1Su4Iv/7Flz25VkSnyGVRXgq0R0F83G0B1wvh
ayS+X3y+KxYk6RbsKEbgrcGRr7NHF9IPnPneImMFlmiV7+ofFgm52vpSHIOGUhTl
JGgZdbMoHhLeacNLXp9LfTTs/ce471lc1tZyTVQFpGaEJIrqQorAJN3DpgsUyAYg
SwqIFoWIIqGQY5qNktE+AAZWj2YvPrueG30lomjEatMNJx7DRt5CQ/KxOZoVnEeo
Xt8a6sTLnIn2eiUfA6sqLE3p3giXrifubymEB++etiF5DrqHfC9kCoIcxcIf/rbI
rZRbz/hw+07UVgX+JYwq82CQYbQPvDLHwDdoVlCfu2dUoBEfbVXAM93/7WUN2wY1
arlQGWh7BwVl67u/Lz1MmM0boaOjH1vYu1BylAnok96N8+aje3lXQNT+PKCssmTF
KSHyfR4WeUwjTy/ttkGoehc4ONAQJ1W5idDqZmmwIYlFLyreFE8nQ1tru5aql70Z
yUf7AwxD7x2/iezY6pS7TRFQv1pvqhKUKt/MR4r5lCD+WAxjnF4GCIy8HwSSEjnk
a6zCmRMvNqOml5c6jmssfIDfZcO/TtQR0JURRp/gp8wMva21J0kzV866zx0ViOSz
YGuQcLbv79/B7O5xfdIvF6Q3GEJZSYrjGPTZwYuqzRCL8k+xSZYcaMqD1YTW4zlU
KinioRsdIb2GVYcnJpR/hWBK2fMhm2GU/vylY+D7zLZ03geqasdiAmuw6RbnqIJj
HMxqOfLvSaBhLO0DygGZ3tASJOtPviMg5HRSa6ykS+t8RqJvxTfSz/AeUK38I+uM
e4iUJWUD7LN+c84WHQa/Q/rBJiMY2vR6Li4XlBUDqx0BoF4lIt+TLWt5iM5F13NL
5rSnwX0+KtJpmS7XZeXG/SB6UeDWwy5juytfILXc5YScl/OEwshy3DdHjGycRA0z
5MbQW3L/LpKxKOx6J/8cMILVIk0O+YrOkvdwgZHd8WtCm5UCI6WQxqaONFt79Ijq
uzbBdgDyByGLBjUgeGAKpyrVHWDmRgdvTAg6RK+ovv+WG8AbGFVeaXo4NTRcfqlW
SDDMNraOxMi+suaGLEqHuDe3O/FK4tb04rgSIqqvmID6StCHw/YeaGSEkhGEQ/pU
mD+lJDVdcZeRcbV1tNYHIWu1g/qGl7un1w42rjvchpsSRAviEqMSFxlqbmE8N4zg
1oWoJUNZRSg/6Row8ulx/MYa9dZwCGE4ChpUd9lkw67VMUBHB3J0T55yJWClfJSr
SywggGHKAMQPW8oqdIFhFGWMbgfGEsksGUFi6NzlQwjJfslmix6iR9wetdnD22zc
r1+YZ2qQHtWOh8wejsokH5koskjWqf91+3lW7su330bikFFbceOuL2P/mWha6TJ9
NewCEMWlXbahzzYEOk1sl+QrrUwLdlTP8cxvPBcPAc2wRDyyCLjklALbPhgezmfU
MsEVtc9jxHM831I2FEUFPBVQX4CHGQLrUoOljgxuU30MiV07hAMjpuOcg9scU+fk
hFVGjjG1lVumqwpwXKrtbMapbMPAeRj0lTdU1MKclYHfssulv3JRa7uV+s2NXPlE
x8qx04FY/sheb4z1P6SJ/uLo3BE4nt28l0X33kNUhkvK39JaEUktElCekwQKClj1
IfE7O66wSiNdrhe5alr0QjzrbqXB3sbV++uwAcrgOdr38/PuLxWh6fHp8mICPmIE
isfjqssFT3dOlNxz+xU4ZReGyKIa18z8Qw68RiUxmJpN5O0cnY1JOt1gOnV9xJMO
svfj2rlhsZFPmdGOPA9Mmgxkrv0VBejlUrmscZ39SuLUM6teBMk5kILvWTEHMEYT
LBVOE8xPsbivCI57J5sHW/12wnErnYkF8oDlIzEPW1T2P69uBhJvPXGOKVITx7C4
WVzfaFXl6/+U3B23Qc1/x+UUMZ/ExWc28Hqo0d7I8sGNgJ72AVgQOLq4GG7P1gWJ
qs/SukSpK2T19ezo467DneoeXUeQKvyOQZYJhldIZnlsF229STJ6r44rZJ973hkn
8fOxYaDOmWtrTYGzrjhVrpsOzTV8opWa6MQCi1bs/yJMucvrELAafxhd6/bS7+Kh
kX/6xzRdLJMXG4FWv9y+twMPTYm4dunCw7/TCcwUGuho6gBgvUyOYHGUKEkZlITO
JxCUhufXHsyTjsm4psH8Q6pNnPnHtKzc+GysrNszoorTwqyVGAtqH76F9NjomQHA
z7NlToT919cjeDeyUHWvopoWNFFbjE4fTmnWeHaeWgbKLxeZlUc9guxvC/3k7p0M
GPG5DmE84K4lzpfGx2BXUy1JCw/tNTZthKr+JXknAZvBsRWpZuzeY3HU4HOwXBmQ
P3srUuQrqQffwQbjkFjZoicDDXGblEkXNQNU3IvwpvibQjMl/p7vPy5PWdgu/qMY
1i09QJJQ8y7s8JH7TTqlhnVgHfC4JIKWxm7VVkXNM74KJR7scSW7ud5pETiY0PQw
lNo/NK2mzVEpuLEILAk0N+pWP3ArkJ0q/VCNRzia4kkarqnxHp+YnuoAyzHFzQgX
6lQnwdxDFNn+VRmW08oEPbdcM51PvmnQRmkKldxhuf1CbQztrjGOgflO/UhvTJgX
mL3tY3cADqHE8qvkI7mfL1o2ym9je3n0TGg+uDP4FXFMUASJd59Q9xTj8o3dlw6s
tAY41XC/ecTSfQEYmNhLMyRvrOIPdd7xDTmRKaPBiaxoBwH9XqxTkCUlLLYtKm73
xFONjRVP3QeJKfPSo9EV9bgAtLsKYBIHjBNVxUgM5bgIx5YTvNhI5tgUQMANuARD
VNh/sRSnK9anW7uKsGamXvUg83NV8Y4neMcxk1fGgl0yib0pp6udIe5fcSevwMNs
OUBvWmrnBPrIYmp/AB9Hfh2UzzcpKahAKvJT25jNhIE3BNneSmGhCJKoyonSk1/S
VURqgg8FFSFxWhQdlZDYYDCQWnZIXxUUovx4q3L0PXN2V089pNwMlCv1vj+Oj6IL
ot1oDFm7tfWYCzPgxfauQNTjDI5PS9Ybpx6wwLPiOsOZ1R1buW49UJLalH+BlZc1
8KVID3RcnIAtYiihg5D5tG2JmOvjkQdf8IDLA6lIfHjsnW3pVA1Ogy4KWR7ZX84m
8iVUBZXzy5PrW62uKS3AvyHQ7dwShtBjsYLAQ4KX3sSsSXZZy2TqOHpsLAzlq7kI
pG7dPr2RTp5gVqRkTtY2O6UpigwrEewOxsPRPMCBUc7WHSUrvpEqbTHIvnkKjXsj
U4QFpJQlhCxt1DIyvIwG04e6T7kkHX315ijqejhG3E1sVS4pVhjdiSP/NW7mBmMr
dO/oobwGVXZxpI/Lj5Qo9rDrncNt3n3Flb7wYkoERAINIgTGjweunnDv8BM7TYdN
joTmfUaR+KydYu/NYuyhJWLUeANMbLXSxaogB5R6Z/kvIyE/enMaoDNzn8ssYSll
Z5sks1HgGa9ugSm/W4XckXX9EvWB7iYKrBhvgniLqW6Js58O+d/eYm1osMO5K625
Z+UMjFKwR3W/QMxOcP7XFJt4zUJ8x+mSV1ly+H7l+OIX1opyGMZJLV7DB5Uflxxh
b2D7glbIrP2lx+NVZnHzGMSe/LdfGAB3O0Hu8SrmpVPl7hc25l/DOwCr8TcP8hB+
foFWhjBmNz/W859ARrJJWPfKCB6qr50Vu82/psMXWVvJcE39n86H8hKPeeS119C+
aeD0jfRoiLRjJF8vhjXwFfz3Q3RojXBGSncXz87dD4zozMSbQb+9j67UZFA0ieWs
qUp8ovM5G2HxncgwgpQYDuwnUAM/G7boIuWcDs2RPqJZ7bstnizyW0JWwO6kM0H0
N8pWnQ2o5aKr5sUVl66kqOCjvCgY+ebSMXDpSv/HMoU05izAVgdQz1v9YlOiKIlM
+KnXiYSWCdsEbQT0eOz3cGTYqaHLMGAFr8Liz05QjexMqv2zmykaSQ7/iOCDwt64
S1Jn1wa8qAZzQH2Za84M7dFWO99fYMQt3+nNyNbtdUlOx6zYE79CqJ6Ml2vESg3s
YyDHUQzqwFFJZuoDUi9Edx2MMca4uuRmJTfx+Wnj/dKKHKtaet2+pGGuFq1DggBq
T2t8MiI7my5P8a+nF1+/BPmidrKRaKmTlGC7MQMSttlOauDLm2vgtOC11RQ24vri
Xbb2bDvPesyhQUO4eQ7tyCmgKol0j5ctcrdQ63UEJ7Q8mdOyJQ6kcro5ztQ5UOLC
41MIf9iQs1AR9AtrQjBt5VXxQw1oZpGCzfokCzocWBiC2kA0JW6XvcDVmi4pjbFk
FuBM7rX135YAzapi6jkaClfYC5sf2vns90oJ+xiUHBQdYzusOt1EOrdQwUMAhJ25
GvbgPoQKuJP91VHZlr4bbfGDsESLQ2dpBMGdtGViMfcxBprD7wxDfl4dSPDglKmT
u0T7oDSPHP69TL6ktQujBSwFUBZ55qo0qtgYw5o+KihAdrwaoubyzDSdZWVp2HIp
n4HhBa81K+7hJJw24wqkDuUZxTNe19c/xqmr9C7HN250ub+Bd0YrJH/jTHYydAmw
zWFDUNxFH9qxlqjajpjYT4pOrPHopU10LH9WySvnhxF0JkZGZEs379Gr+QCOrVGv
B0eqNND74Ucory+8L69zLLaPbVp0kU9ExalMwbh61dlseMsPGIKDwiWffYJj4WYX
dVeZmafDYm6fTpf1DYbM0y98jUDfKXQ2mGa2oQEcErrG5gjd/72Fjafl7L3xe4a/
FPRlTroxjlgPO+v6Y22jC5Twkw9xmL8fx1bN22cWEZ2J1OCYsPIPct6j8i5khz9L
xqQWAJEu96J1Ig8UD+PY5nuFyaIaS7mtBzKmbVVXrgxbFw7CH19basX3qZ2SFXLj
L9zwml2p+6uv4Rh/aUF/P+H5R3lJH6gTYw9nycy3G4xG9wWY4ShBwYyUiTpIv1gc
1fCIJgI834GFQZFsQ4odRTVAlqi49KtRtGM6Onb1E3fbPGHtYiCRWnzi3MhoB3Nf
NQDhCukQdypKZuZHPDZJTRpjwMo2DfR5GxNnhKte4HbsNmcmTbFakwpvA0ubA4qu
tWkEib5QZXmFLRU7IAxA7VB6X26qgSJlO/EV4GGhPaJNkxrQ0l9IbGjv1PzuF1Od
9poaY0vT++EOxFhcJz/sBrNYPWmYnwryRTSQ8JLCyLDzD1JtQ3yiGQ6CrfGdWszH
QXTmD13WYsUlTu6rvo4MxflqcsMUz+QGE8DPhTVuNgHfhFdSnE/L7O6Dc3RVtHGc
8RpsWqtWBzQPGuiQz44YCNTmGteQgdzpHEHj0iTbk3EyAQ/QoE0xnX7kq/PCbBKC
biPMqzv2xNZD4G+uMhzXH26VfcVuTeH26OTz5jhPmFmczpUl66zF9DtEgmacK+FG
8gPGAtP2keq1U8km1kO3hQojqyxNSqjQNybt2Lm0VGoJhze9IfZ97RlIYR/rC8BA
M8J7JjZ7wnKkhZH5qEsZvpLG3R9E389NZ4jwvdAQ52TCZDcsRAkhqPMAQgBb2hMr
hSASRTJtxfS84WecBUItd0JdMN8pGflhlDpIKBUT3Y96VzT4sqRzETc3xsp4OepT
9tbLln5IMtJ/jHjpcV6POPy4SLl+MuoK8yaZWz5KDeOkWUrskSsdU/giE5Lffvn4
f35Dgq7uUmZ5oqOl8TGoWb2EQWAR9dd1mzEc6234BcIko62LLrsLlQ5VJ3mRvRNE
sJDF2m9+HXsHXIoITLJli/j3k7GdOkBCzetZW/SaJyvrXh+gfS4duA8B8dSC3J1x
3cBtIIrFFYgnQTKByy8Gkn85VM/EuvD7SIqfCzJFLOe/fKEDHLTq7FXv32eY59qx
mbnTD6LCNUkxHsyt6mfUWc7rQVAmh2LMA8K9QO39HY5b0mXkDlekRXIHFdfalNCg
0litv3c31eU3wbrzOsSgRZVmgTHA2v1gY5kR0X2QAHNORyQ2rf4TLs8gewnAuxoh
Z6yoptK/o3HQkeXkLDxyV87myZzlShR8ni0UG8oaUv/7dlTBsDyI3qKgXAUqrg/g
xQ2txZqGXd8R4D+Xo5KbSyYtp+AaoQ0vdbBrwdLGArsjd2+wJdUTdUM6IiaUOhz7
uzKkgPDR49agvax6cDCGTOStzVHNgQ0sTR32uUaSrRHXc916bgfRM2tGcF1wB7e4
SRtjZrlFLHvBwlEqi70iRsj5y/VPEGBgFY4aIc80yQ6kcgrGpnFJ5bqcO1QoqxA9
2GWOCQQWXrh/khb+bNPsYeDO1sdlHFClkonVBSCtthGkA96yi/pByUyWiSX8LssB
saytA7SqW82heJv8tmMjvmAKeUmpXDZ18yREmzY7coa53hbw4fKA4l9zoazBvo4m
yx04/qhjoN9fLAHBQY4hUU66Jft33+Bh3+/aNRRaHu/zWkms8qazuoEHJ+hoMDUU
uoRUf6DqzPNzjyRkgreooSYbcTN9A1SxmimysC4QLiJfd4aSr6o31Qj6Y/hVN3m3
yQtlKtyGgSpIFRZnL4lhlLUk8nwSMALqDCzmhw2iTAML2RIehy35NIo+azvuQKnW
vfTa7W2k2VlsiivhN7Jnw7s6/wU87MYdkD/2a8JSEyTJ28i21yQr+7SgZKRfyX7a
5MtZqhvzGfxewff3CHHMt9bABGBy0rz7gN7Y8uH8ydvVrhQ07NrhEJyh4kyqvWVT
vhyeigi2YKmSbGDesMPvBxbkp6ydzJMB6ubn6FyXDoZgagcHqgzg528Vc/7CHKSw
s5NyH5DDeobsD4q7qlmdMTR+E9arvcTehY6UZDfWpAwMX9zedUmx1KzvH+SfkPSW
eOhRYQj10Ul8u8ixQFUvove0Qi2kMDxrYn2W34BAAgg0gqzz709bVTrn+A0lefO3
KJ1aiAXXbHWSpq39PisArZjsuQ8HqyU9tcTJfzzBdIb0AnBOMRlyuQNEb/fSRCYq
Ohuk2bobZhXB1vABSR8Ok/sH9Eh1QK0CoCCUINABohdkjKebrTVkRAwaXgIwhk4s
ZRLaMvlsZuj6r2ctdiFmSotByjGyZ2wx5vHFcBa+PXGEJ/LjPUPtOVSdgU4rsN3s
yulmNDYxgTAYc2XTRdcgENkjK56fWxXJofCmwGu9/q4PtUE59La2ErezNfbyiVbw
s1qFzJgOZQaAHyNQCy3uVhMN6KeO/V1n9x8LlKReSnhp0Co+Qn7YkVogXJUr9vNI
cpBWyHPl68LYpctZXoa/LAvHv8IUn3UASQCMWivIZi/oqn0FwBRFWmRl6NRZvTTv
K+cf5DmbiaYjVDyD6zeA7IzMuhsWOxgmBda/R+r5Rybsy/55a79tsapYlL2BgLfn
EaiAXBp4BnAIIxd0gjm7Y/puVoRADFeXyjK2jHg+FBQIkMxcpRpJyHttE5F32hQL
P08eJoQ0NlnMnpUPS7ztRVxxx8LWHFuLxL9FkYSnlWqp/QAejbEx63AW+LHGuD5I
f11HGnRddzbbFIX/co7roefoBe/enhTFZkKKc5d9vDEuBCi8WkbWlDNEYxzwItco
Xh6yiJYcU/qAxu9iO6SFr4YAph/fRSpCi6mgkCrXO7ViwJsPiPZS+VMDWB0+HiYc
OcKHsjkwxnW6oRwXDZ7D/JDFAS5orNe9VHKQ4pGtvm3d+/rCnrODupHM9eXCQJBb
IFZn5vmXeIaRdrRtJJ+Sf+DXGpeaPgLvZ7RDXyxZAKHmRN0dJiiBt8nG7oaX5bD7
t1IOuDldkuKU4oubEXDcs6ZwsCyRKxpXHmiqR88jp29UJ/Of8rgPeIWvaOVYY0Le
Bc/UHqPtOs4vesbBCbH7lbbJO8XGMEfLHuSI7WG5IsI6AavBWm0P8Zi2rjbL/8lE
8Hc1OM5xpV2kKIyYeWkbduX327CefPhUMRb6cT9iipbGhdk9i7G+wRo+eYUqQT2f
GsdHvKX+8wdzD4sm/eOFKV0rDYhQkXsYf6+Hq6dNMfdJ58LQAULDCvkZNqBZaMY5
uHBJJYEDbsXckMFgiJ676hcJppsXLhxkYiSdVkxEByBTHolagvwSJ+nspXaz6QOi
mx1bUCeDBh1t8ToN+ibIzr4Pe4OnowP9i92Er2XDkMOsUs7QX4635w8MLECZzx+L
EsLqMz4hbUXUaaJFwDaZpnbQkFXigyAJCzvZIwG+S8MXen2zxzohsLyynVDeCKYK
JQk6Y1KLUI1n7R2tyewzHkcDgvuX04Gl29P7dci4f/eCp4hu/sVMu4w01IKTAfyl
0ngwX9359C5sV/6b6coupo6kkeNIPO8B1fD8EFzgLE0Kz97CgqJ+XfWQlDmKIQRZ
MzaPYL+0f77t73NYneU3qsw5rSA6BM7FOwOltnY3GJGOI+60EdIQCPM57sTACtnF
6qUSKZpIfbuUbiuaQjqbuWge1V50FyS5cFpdtY4RJw3aWPUSUvJpHWjd0XCruQID
HdLoBo2FrNcUVYw2qfIar261OcszBzrczoH5t238jcb6QLyr+fDgTPAQ9oJUiwYl
4iwc3pnvv5Cy43kwzlW/tAtriKSNWJtJEMxiv1C9E8EI+hUzEXwueB6xqALGRpSQ
7hionZd35FWRXfvW1Z50LlLpUVsASDntxA5kP0JjsncGA6h+qUhMS9pLty/7S/t2
waf/CmPjxKgh027xO6OhImZvYtJb1Cf/NjiEUM+iY4hOuxTuS38uM/q/c91TjEzr
e+mfI7XQbOy6F5bUoOfFnvElOAF/qofWjPXIk1DwY62f8WSYPXnmrTgm2crIO2uk
pgSUkXe7rRYHnRUWIpX3NPksh6WubPcpDqVjEu6/4c/KiwKhPlerlP6d8lpgnCqJ
TFjbX2ykL82KzmqQ5mrI90eqO7dzZCPjTk123AxM+vT+HnQnVnZ5eHCiURptOoTO
K4QTwV617SrXbdnDG7hf0gMTyMGLOx6WwzjiwVElzGmghtbxKBpiz/rlJ2yD0a0o
yWUYzr2j600+kvIe1ZK3qcKYepey3n1NUh//4DQmYgHhxrAnXNIG7YkTWIJ70WUt
y2tCa6RICjvg3B4r+E3Ka/Ly16Aw7FM/EGA7YLlpYc+0qh7WasB/KPmdV09KYoi8
+CnDsaHUzjT01JyvTaZoZrcr+J9XjzWYu/Tw/366QK551WTY2b3n6MZH5TxJISpS
f8V6oBuUXslosLq0eEvPJNY2jICftbzFFmZmvP/iZCC1OeFR2PViHXTcrq7mGq20
4gQMGFqNooGsaSanP7kieJ7xVcTdK9OZKkQaeCFLXk4+eY/a6jbZPipYhl/cFN08
VXHsdhMbvWKvZB83y4hlO1qAE/5dtaW4qmF46tnKnGGdbK67e3sSeT8HoRh9I7W3
hiYy/6BdI/WPAs1USW+hopOATFbyP2Fr5Vi4k0+++mvOvvuxmgt7eE5u7RGDEMiU
NOagDWpgvLe3dFTSTr4TXV8eBwvfZZBr43bFl9hm9BGbPUliDSevQkJ/SF1wQ2Q8
3eJ4laQnl9ik0poMO0vdC/WKhEkW3C/vojwrl/GEKmHIgZ00gdKE4HU73WhxxgOP
1vhzsZ/lqXIcy0xAEBCmjS9NI4zQZ4Nl9EWd1/iw6O+iDTonfrXpXSh/cJZO6XHV
VihbLRfyd6/4SPqgGzJ/lTjF89pV9aHUcdnGs8sUiHCd6BbrdJZWty37sOEDuKXp
FAd2tu0IjssshTj8EmLLJwS0z78Kw8hAXhGLQHt0ahdQNlR4P9BRAhJLm+Dpm9oQ
z0zFvuPI4tcUUSpUNuOqsnu4nDrT3k/blp95+QZjYnajRGvDy6Eh3oJuRWmOnvvz
AXkbsUUqXmLHzWdXqerTjk2qqDUkc2oJx709awfx74JEPUNQWtzacWSqBltxUv2+
SxWhJCTiv15T52vTCIBCWf2hQKnnGS6ud77W0yL0434zNjquj71+Lsgk3iIegXwR
R8OAg4ebTCRPjxRzQJJNXUZ0UPw3/0b6pEvQzI1PkTOi+suxdYKxkTGxrKxl9mVb
ZQ8hpR93b1BCNz8l8Nx8S4qcJQ3qPr9MzbQi1glD3h/vCMj6p9lo1vaSUvk+OXb+
OG3zfqgd+sP04/jwlxjoadlysS8ABlChX3JafDzmJNvSc6OwH9YWo7LsvIORkDjy
j03VTUfhVYuK77/p+d/xqDnnGEFX1bE+KoMBchrhBl26L0c7ngNoYCC993+YI0A9
XfSS6iuUpte9CeqmPbJ4MplRIPbhWfCSjfcOQfpymdsxU6Hn9yDZBdlv8cHhNBVH
y8cf6d6DvmxxZbvn7LvpzrFI4b5fzhoVpZqXt7dqjaXRecAh7vb0f/lIc52ujb1I
IoeHeCKwMPuNAhqDzsR05dxYdQBfvHyv59DYzlOyJ6BF6DdYBSLZuoLsFYRXmHrU
tH3Q/IX62JWLVXT2URN/II3PlGQivkqRRtSm3yCP9JGB8i6e2jExPXBRZaMMakqU
7Ekm8ItLSx79vFBHdhge6h4Yxk3uteyMlrEj/qCV2icS8oLrF4llhl4zcmF+0xyI
T7VTi5ZJy0ZAZ8oOKTzEyGrrhrtCIvvc2mYfa4tlOtDNbFsGpR86VwxNTEBnbjbm
65NEZPRJJKj3oKPXtPFbtuOp3RBoJZdHtHPsffTLN6bgIKTrQM5mwiS5JaBDXsb4
0zT472zwrWXtMbcKJVO22zis93wqHGqU7bz2D1wP9rmIbsvT4mMJLz9/Fvmj12ZG
tyo0Z1cLDCXWTAipBSZk2PxVFAlzDIUHuANTYYpSRmY35JPYFt1o7j9xzrpJwE0M
G3yA7xfWMrEkPhVzkhyyhDprgASfabXlcE5E844kJk5OzG2xqyF2DPkfGKLhvMFk
jPna0NsIPy1eD+dK+bFRczxM3QmHrrrNAX7x0i4YbzvY/VooJ73jlRYPGqTPhePu
mDCBv8I4mVpCKyFK6ZjAIlDjooJuUOeRyqSepsnY5ijkzrfVDi4ilAfUXhQ89ar5
lpmcAoqBVSIC+lWaqmwYnkJ/gho0BDRzHP7uymtOtdQlj/wioQfzTRbiRx6i9TrN
xLXBCDlsmXfFj3lNMQuxhIBZttVYytEfTOIrAiUjYmRkDydDX6Ic6fFdtB4m1kuP
B2r+FUIbHfMyBdDpNxQN+cEpovnjr8KLBJMjt+yCu6JHuN6TZAOb5mK1V7atuXcZ
BjZlg2cPywtTgwu8qjuFlA6Xh00hHBqFLpmU40L859H8VDRjmlnTp3EU9Yeoj30k
BD0MljgZHZo2F7rfpLdmGQRKax5IX6+5KlC02roU5Kr6iFJq6k2/cB3P6xXW4CvC
8QfeELeCa8yFftN54c8qtJvUIxwRZIzdEVbusbEfkDpxq1SZlTOsFf4yZOm2hE0/
UR7xLtNztvp7DpT5jh/EVwk4mk4w3lzbaN/t9UD3xkF9IISf6Tgjr0Y5J4VupumY
KdQQ2OFyYNJdCSGlb8Qh6a0aChLm1ZKfa6Ey5NwWVr/VunyOoMGTPOP4vDxHqkGt
lKL/XeaEsWhphUepQwCJYklu7YLr++qUqca+ttIiM8jmXGEVYXxFSBXPJhJPz6r+
mnJs8P6RYequSs1bL0GzaZEF4+LXvEvxvlysvOU4iXXYbStdR+95En0Rd/41gU8o
oWfR//mAqGjNWHkY6qCr785tRpI9/NM7js3ljY2d4ykueZpgoIUrWRqqqbv0IbEI
+drpsovJWQpDFYDTOdeZooVNI1wuVpeZjLsLk11q2bGGgwbjrV/D0Vxqwq1SNWku
qtR5+uLr5t3vsGhERCY3V4MdZ6XooO175VbPGfweXEgbQ39cmqInuscG2+dq23z/
DB/z+rMa4pBcGqaOM5ybV5jbMZY/HzPyfYI4tFmA7S3mNHjT1UBmxQWFE9Z/toZ1
e5j6poeAKmI7A5smdmtrfrB+vxMZC29/ImXaI7MgwDFLWioFuyN4ZoXN87cnXjry
3ohwZfFCVwXiQWI7sylzv7KeZJiwrmPVsKYSspUoo/yi5B5XNSvq8kGFrEZd8+LB
PVfG5Ddh0Gn0/6yTngH17mLjzXdvLpuyFlw+868jpu1KIiLUvNcFr6vu++rvSAE5
fMq3pHwXICnf1b7XnJBej3WgxfPJmfEOw32UXlb6gPfjYRLL6hMlYCG4K1KEaZbz
U/kbsx9Ogp7NHQhw1HQ5m+SelQ8sxdOnza0ATthqxR9/Fca0IzetPL+M+fjoRftj
Cn09nxhExugiefqty1jtR15v6JdVmolphniKm7JWosZ3k1NTRMVISNPMG/iFEXum
vcXx6wEoovbQUTWd8/X/AXDa1093xWZWQv05NsZ7HiKy6QJ2S8k13xpCWGlL+Oo9
IHNfEEI0aJL8rTSbW6XVZiUK/OGaDo0kQBgDjI9cb6ydlNfD7laOmh4i5sW6QwAF
V/F/umqbI09JM4YkTivcGAYZVsHHIqRLRUHZVOLxSQ3qBHMn77zu/VhBpbMBLUyH
DQSWBKD8nqU7Z87CiUt7RfVy5nfbkJ+LWkGKkZ2E3DuAT8BYt3MAB7s3D3dM9zCy
hY7e8bncCbzm5yOuI7xNg4d0qgYmzsLBfxx6wZci4tsbLdxeIML5Ac5GR4x6NiXw
IHSIjXVb1/vTBFZDPXKoqp1Il8Cl8JNgZJ6a1pQd/t86M4ijcf3tKHQrfCI1GsMR
nGPu0OywTk0PgknzmdH6s7rHOGH2OTRABOq3qyupUmzcuXt6n9Ld0T/+OzW53hn/
E3Kgu+oQNRPQThtyT+uvzawD1dDvG0YOnaABMDfzxK+h5xEKDlBKmmbbvK8OCWIn
ejDrS9gQraa9L1kH0kBTn59SRPrqQ9JJAwaukyxUiuSm2LjhsKCibTwGHdyIZoDN
12OLjutIRRZ7+lCmhYjJBTGx9WQXuGAF+L9TnBwHQCGltUkeoN394j7m4U1oSEa4
oTgxQrYgDnC6YF0PK76+liC5KsTAEAOY7rZdwuEfpAT7pAPJ0ZhL4MSU8PsaMtgs
xL4UYMxoDcXfRhWKbGS00J4e116Sj3k3QWeR1Ip9YeKV3W9HHicLEbxQYr2QzhBR
c3evoUOPfaaufDN3Xf9FL3C9/R8xKmrgOOOBWZdlxSFS79EvqMJo6BbXQoValjTH
K2i61vqTGzzDIwO5oWQvaoWPTyQwKBoqO8kuNXvaPoeGgFiUt5yry4kpwAERjMUa
+rF5NspffDPtNItGnsNanZ0mjp4FtAa4lNQfpEMrDbstnp02nN3UdPVSeekVlExS
YsVIvpKUAWvONVBbW0Q9+sXJDEhrQl+FmSfEcGQ0pNcvp9sAz5yQ6YUyrruUECXA
eipks2jgZNno4RoMBfNTm2oJv7Lmv1ah+RkQWstITi+FjDWCdrYewP5dXBg9blaZ
SbZ7WX5QS39fuzaIOqFnPz2UHsW/cD61JNHhgHxkIJEwfyMe4Ys1lVcJXnxsuEQk
/G54QraH+6SfPYeCvCMYBXIeEsFj6TCcQllSKOUapn2G55MIuUzbB0le6GEl4XIm
aH4TEA/NVpeTfy3b54QNPBcsQ+7zxu8OgMemrBsWpUZZxB3P5oqov/qsXpOmMiIJ
OBB1XmpcAOvbIa4w5W4FD8OZoi88cDpg5VGMks0vfBoa6tnoG8mOnic0MaQIg6m8
WklgRCJAK5KyBk3M/82nQcT0s8av1aQgg+pA3KAcaRTqi8gN2b4Y8iiyf1z/s2/4
dJOGQLDMYXntRkTUqhRZ9yPRAJrmO0zDR7EfG31/i/4XVK9OsMu01XKErMXAIhfL
Od8hvkToiEEpahiAhuLVlm8+V72tjFyb5fEmONsMAp6hJ9sciavWPUi/XmM5XqKa
G9zk+VR4Sx22hL2PRgqMqrIu9L6zSlxhc70JRI18avf+1kGdiQVxHcRezsj9YyLM
R/HuaMSDsCX9zp8b7zkK6NHOm7RRe5a1mxcpb+gbKE/SC3eI7u38dm026TiOukcj
X8MPpJLPn4md48jJU/ol8MdWmwSTJAMV7I/QXGvXpf6qj6hPAcoJTrkJDD30J1IB
eVfdUnl+b6PW4qBXNRwEwv/DII1ygVWEbbpRfrFSxBIIvrZjsy6/ny815YqV/eEM
sRkReBHnL4n4zoWQJUlMgtbMEBp+6Wpx8r9i/P5przB25iuTna7MXWnN5qe0OD3Z
2g/V9z92fAugsullbo9rKDfirqAnk1SkjkhKKThpJnUihDOoOaCsfL2n1I5gQ+xb
Sp3XK+fRU+tge+3J7yHNErvL3+YgURxc0Ido2ZvGmVW0PZVXqm/bydMv2OOrcaTC
xKcPlMxBtdHckKOvIGGmtSqlzZNDFL5rLNb781OkhF/ROZZJbbImeKmmfHUrrNFL
F8YuJlMKKte1VuZREb2keu6kmvfCq6BZx5E1Aqqt54+NRP78DRphqEGnueN3A779
4ztwuwv1ksDWF8ALbNFfr+I1wx13oR60B+SjH401wV4Hobx9iS0rPGkA+ncNa9Ws
RwB2r7ut7kx6TWXhDvTzDHIWPuLFRLDId0nFNm3fqNm42aUyl0h/ePWmAMxzyybG
y2Hq5uquy7T2RFFJMT3Icqj548tayEWs2x/rWnh3KFGlv5VYNnDRciuWdJgJ/xQH
XMbEjKmikN5b1kIHepf13pJ8qrnqzY43MVetNjav/yXLl/ey0/y59nRQi8CpDRU7
4dZpsM+u4/wbdM5jh++Osx6NuPBiR+RHzrWw8U0gu1q8QCLXSTqNzANibdIln7LK
sfHc5sqZzslsnKAJ4GRvIuyDxEvNNb51w86gMGrTtAEsVW9N64fHZx/Lz5Jq6KNn
sQVbGqck/4jyJRV04WuB4XX8bJkCFVUI/KV++LdrsKCgbmwoN8Oxxo++nN/W9Ozx
top6T8aTKZn7SaepP79beo4P5na/e7w1qEcHRqmXhpNAQBQWLw6qKk3JZ7KPHJtE
ZOwnJwpYA5t9xEahr9Vi9hpm3v1Rcf6rMeSc2h5tP6pDp2wIFj0znlmBaMXHse+t
J171PgYFXsXPVBlQSw5rDxbaIrQKVTKXztgBFGy19th2/CwkwIDCxJcoDLT19g5t
VYONGSOxHXNhXmhD/mq1tyJo+jaNzbd4B5RBR4jl39CmMwZAEReRUY9DegDGEMD6
zLjlSdixpvIgJRM9DONrEnjHM4eD5YlE/z80BBgMLC96fRA6NNF4GE7/9nDRaCPO
GV31mmKl0zKWOnUcQvgYLoMz1ooUZ2Js4XmYuk5i7oxg6G9rlmOF9bW+TsAmBkDG
4lBB8nGdv5266SyUIusLfTtol8QNTheAR+y3PJSPAx4Alb0QC+UO3GMlxF/reRHt
sFJayvH6EuHlzLyCszhcL3rnm7ARNY0vkD5o8LCKn9Jw0twIs4g4MRjxp6Ey3I2e
tGLPgOhHJGwvsnTkk6glSfjD1ddTT5VNxuV9M8FUSyKWPN3hICzU1oiANHaCEQti
9MZVyDuCVC2l1aB1tGyPuErJICs0bm9NRcy9BHVaYFs0sPH2VfNRC3MPgrr1a0s1
hWDE3Bzdwz5mYVZ/M7sQRF87b2PyfPadh+Ks8uuqPfuziWZVGuhdxZNGE5rP0dbs
QqkoeHjqCaFfmsQypLSJZdQ8oc8mZijdTpveh7T5MmSsd7T7aD7voJJD7oyA6x1f
x/UOsPhYDOBBK/hPFst1tARIKPnv0EabIURv48NWAR1LAZdqFbtZ9ScZbtiOOavJ
EYFHbV3IaCFviwxfp9qoHzTc545mz9DPzPLiYL96uT4iAyZL3ypS0zDeqy22c4W+
NoVto6FjE85kAUn22WpOGZH27RTPI0pVxHWVmnXA3q7Qczx1wCalkqsNO1LAcv2U
EzNpliF+YNiUcKH+qd+7Xj2pxnLan9GvHIkIkfn/s1BZEWYiETDRV9TwcxHy2qE3
saoVljlPZbYr5taxqKBp2hv52fnNKf8/ws6SMNuXUFFoBgkkvN/eZSPznYJcp6AU
ZJsWrggKDgvUMyDX/Po+KgACgTcUkLvukV2GCnClM970EDcQVrfkcKlICjg6/MkX
ZihELlgR2s8ElMsf88LVHxHR+remeGnR734jHD5v6sh8FBFwi1g8QmPTLs7xu4ef
X+4uDjmamNrROnuKNTaH5n8QIpdGkeLXNMxlJ1ndm6NbmJPDst4Fvtqe0yoMG6K2
jobADnYC2sNOqAD5n2Irq4s5gfIqebYf+p7ZcNNy4F+2Ci1kwPX7wGC4TghVzNTj
xDaEHLybZrlbRy97/M7zROfGlGKGCW08mNMzMqv5HgG+gWGLqU5aaNkRl8Qnx6uo
GXZM8SvneXl7YcYQL17OXe0gATPgFt73YmHpvmUWx3ARxZTxoO4GIu/OxmG96ZEu
SbDHyDHvlooUOj6jH7/jwAbURZBAGrBPZUXXp3Gyxl+fuwp1LM/e40GECEF3+zsZ
V9iwoTYBrq8KT49MQ5urejXqyYBWxES1wNTCc05VmHfHAli6sunFNXIAvUAYFOkM
C66gTF+twEYZovIWEY+daa2cn7ad4SysrcilPBCLcBx3DsPigKZNo9yRtRKlPQs6
3P5oHo1ArRHJsXWkR9l6/67lbLMI9/6ekX0De/hLHwZi/w6OQ8kn7UC2Xks5eeNf
XVKCrSLQ6rQKeIm8dliwHsEEv7qWtBneGD5SEdQSUpZiC5lP3N38b1/ROm8s1fkv
WTMfysXwnqaUnk2kKt9I51t1J+C891YYGpW9YC3IPAyT1ialGnQhgjsfg+FB4Qn7
eA1lf6xwkz+FPyUo0xbjIfBlI8a8M21HxcLQVGEJMK8IG4sTqOftRww/n60Qyh2S
N26gq9JyQ8UPIGgrUvN0YSazGoNIRhatNU9uOTl6XGiTSNot+kOyMVkim5CpbR6i
x6IGu5Q9PHd8NuYjYdZpwNmfU5ZArjUZOel80tBxkVJN2PrmEvUb2uR7MoNSk6UH
l8CO6HbJpqtSPz6f1/H4pMYC91mczrv3sL9j6paE7X3eWMWeHJzjTWfMCH+3f3Np
O573NKD5qXY3SS4j2clhDmhmrvvQPsbKqKSyemcnADaHejysX0EMpdQENjShTG1Z
A2mOG/1Rscv5tX4hK1WN26BXAsJGqfvM0JyAsaeGSKByTe8v0NX+NW7uBqWM4U+P
fqgVxHHt8NVw0u+BNBwdUwE9pyT6CSKwaqEmbcTBrPX1PzPRBi6HtqqQ7ulJWsb7
m62RKklTT1NG2gT0a1c5++kTfBjPSQoIt5LC7ByaOMwOrAJZBHWG5NqfEhPsJpo7
RXeEZMAc4blm8lNrE0q+w7SlKZ4N0suJTXNRm+AiwVfC7YDPCT+UgRpuW3tEHzCp
DSwrQkNeuiNiVAVIv2hE0lVMBEt2y64w9MmibArQ5+cxYrCBrQqKCd9PAUfNUwOL
zKKlv1qzC1N8tG4TY+H/8o/99zHeOafxsggavQNXrnOqpNFKQGB/TPWzJ3RMZgXg
zu1pLmHme6LuFF3S7dqt34vrzUBX1r7H6a14mbenadRKltNnJ87ibuMDCWHLNQ89
B8+fuPWbO4lF8gwzv1SLjJaed06AORk6Ekh8RxADmXBzKKJs+UQydvtC6QNLJ/x/
YPiLJ1ovCjcLTammI6L1M32+DuEKbBuWHiZlh6mqFHUxPBz+FCXPeEZ61eHmGVyT
kNz6fdX7v62DK/X/NW188TNl9rFo80QA+Nndqh9C2CVwca5Zkwhgtu96U4uEc6t6
MV4nyyMvwYkHvv60M3M6FeXIUSUJ+bZ127qBTsp8jLBsFR1DWF+Q6azvfHbtUG0M
ON8Ien5W9bmFpThnqT9/o/VOz0pc30aBkv7sS1cV7QUEVzNyO/Fx04wemsEYtx4W
ZpvI9qiE3O2IByW4u60642XsquaKE5p4EWcQBR98WhCqb/aUk7jtHp9pQAZcLU8k
qNbVSbAkOfwiq0tLk2Mmv2TK1dKscXKYr8V0aonvIy/E/Yg+ttstOJjlC6S4eQ8R
F7xnNHmnnzuIh4+8aIeM6M6GVrRkxWi9mIELP+lt4Fs7Yd1vSD3lTzDaufM3lOuZ
NjXZZSP+uAaKK/TAI3uFvL963MvOVhjUqtRO1xuTLitNhAYt9SvMwhg6f2V/lL8/
2HLzWXYY41mzaBWqqA88QcrzDbeqjlcn96FnKOnbYYWvH3XU6e5x1QOjfLGw1wb5
TJegRyY5t+EAUev5k74GrPuvAWkCZEQx0VBFKm0FX6cok/kJZLJqPc1QM/u5+r/Y
8eA3+6oeYjQYeKC4P+n9cB4dep4Qu4vPVYSKKLwoWxw1eyW3KEAUbN2os6RLKq+9
Fn31BB2rhW9BAVPEK8aqGyBK0YAvbyAzw4bnPu+qfjmmFB6yTXigjlv/dDMWXukv
ys0nAgTT09b4i396oUASAiV7u15bTjlzMqgCjupMh/2bF4Us67uRu2YL5tlETxlj
uSUNKeblSD9l8+/yehcbzbsdQwi/TYAtXwxIRb7WtU7B5LpUd1E/RFh17HvCNuM7
k8VHgWKviSHHlgeqyqFrZCHKvOQ86Dwbp9fsxo1UMTyvYf/oBQnl5K5bI0PHVEgt
lJhgCJvzpelC4BwsrNnnPuJA+4aCbiUYud6meBYN2EcmQ8UyV7OLqaXUjMks4itz
arG99KUCiDTt6kyXvIWrCo2Zva1YCVhB8O+cOAeGHmjiAODt6DNJ4kGVfK94BRn8
bGafzliZAJqVf2j244t+okez5K8asaW3pu+PTIroroqtLlLAMkFrB6JY7jw52SXr
MwIyMAudqA3xoKvLBV4kaxnG2yPDKinXmzaqm0mKKkPuWpbSIaplkJ44G7oxGL8C
Cd4+AnhxKH/ClzJbGDqtEkjT1naWt4wJwWdBZp8QevhLGYJ8xT5FjKjcvPGCUV7s
Jjy9ObGtjLJKY6Y3yt4GisyiJaVABo2lZbu82EG/xfLbeQVuyCHodasrHDN5k11r
coe76XxjS9gYocanq+DrKW5uGY9IICQyTKDUFPWUUa6Y4KowSSUTqd8DaQhAkZ9k
ODzyt9AE9Z/qA292YiQgR5Lx3rLKezlP9bfC0Z86qb90ueW0gQf2Buvx6ospeiOh
E/jomN35fowcS0QoJpVezVpFc+K4wyM9JsSJRY4dHZT9Kz18g3AZa93OXNuqBObx
Iulozty8o9ck5Dfk6+AihrDoz0m20xJzVPQTy6EjqLT25FVRDCGlip5lScR7GxPF
7nGnlQFI2zs7wceN2CtGnjnF7uTuJf8iZmotsvZnClcR2eiPb6FPnNURf3v6Bf33
OPiuneBK+aBQP5BsMsvEpjhgwEmXKvzyomAWXko8Ung4NKhLZVsm9PSveA4mnh9Y
6efDtepsZ3iadOfn0vtly2kIUTSaPjGAEFwrV3FYwkgSkLVj+yx2k0bjKLkACnpQ
wb/ZAP6hfaNG4COZZQYKaXbJsfez0O2/dwRf4XYMN4mahGz9hqAseg7xzLo2NyJA
7cLVBBX4KXnlOGMZQ1+ym+9IodUMH4JuL+PLiyx6Ui9b5gDciZWkF3iUvb/czKYi
5V0U4to9EZ+GcGRmHKR/IzxXdimcSbyprJxFV9TZs2eAPDxGriLahErVCT9dk+ya
QdmSqxtOSohdDaBkxyMAwPAGQ6R9JV9nkbFb041GnK52TleQk4cNHIntHEypHdUv
5RH2NAc6errgndmpDR0/YrquEUFracVzHhgHdI5jLfZV+bqrK3PIuXCv1cb9C7tg
me1MmO4sufam5DLtU1bUyMVCYdzwXAb1V0QsVooKNH0OhJJTpMs6rEKJ/iVXIEEq
EsJna4/MbY9zM8G5FLHVdvVLpzAEtMfajj4DiAgd70tdrJAyDOoPzorGvBXxY4QO
qE1rkT0guyBFnN6URQFoMYd+hmplht9QLxf95PkCalI3wWI/nCk27Hxa8dzEK4pB
klw1PuaLRiNrJxGvnHpLtKrKEaaS09QHLe5GVs3xSLi37kZQFKbxkDMpRzXxOp3Y
yJQwEbQ5+xjC+IZ72DcSdFS5t3aXm2Sh6q+rGlCX68HBYplR86sWVzlUbrULSETZ
+ve6aw7ECPYa8aC47kMGyMdrwBTgp+V3K0GpUfBGLpKcsUSTD2KM4rydwhQDWUNL
DEfmwWOzyYF9qyoGQXI68duQdP8ciZ7MlnjWe73rhzuciEsgynuBrmZbXaFVIHwc
oeVfdfpJeuw65cZJRWZ87Ce+Mv7lr2ZJPfNNaxcdG3Fe0AeVM2SSY3akFoZGc7mS
uy+eeL5sPTL6tiCnLl3PRKRAE2iB47QA/wS5K5N8e7lhXr32g6lq5cIOFruY5wKK
BZmhe5e96nnDl8Go/9XjJYmrPZ3ausC0znoHbQI6t8n9pH6wU4na5Xkr/VDNhaJz
wwBU/BA6oVh6vhIYpVs7MjVj5Z+mqhZnZBbi04H3WJbvuIHKask8TOiH7nuYF/u3
vOOFpXgjG57EQbVxkUK1pX5f7I5YYZ+NZvqrEWK6dkY/gHiEErWixhsd8pnKArHJ
scfhEhUCjWKM60QA+4kXKWLObm7MamsROuUhfyNLAUcgmCls3rDEPGQH6i1j86F6
bbscvgRISYvHp0HKGWiTDpms411+qkuA+IqtFszV87O012gEwOlVHoSdVceg3gSn
+r+hIApYhAQMFoB3WqnoFj84psF0PaGsEzkjT7Tt5jzc8lnTwpm8QdgtMLob4rDn
/9oQfsjUfLGJ4n1vR95wRyj7pK3se0IeWwCfCrWagFEN2IQxzAM7v3/2lJ8arVkQ
0P7oP77Mf6tlafbzqGu0yQNMo2OlKtNcwL8+PNBrB6Myp7XF6vkFvfycmMAdPRlk
hVGIw8jldindRkG/A7bYrHEaWPaVlsh30sqg1W5tjDN0N8O+5P+iBydmHUsKAfU6
gQxHxvadzRAVWFYisccArhXhWGKyvAPwS2GD0Rg0VSyWOBPJxfb3xhrYaLeqfYdu
VpPBCRUK1/m+N6aHPGAdrvvvpYt7bwptETIavKAjCxZYsj4Dtxx1S3OnP2etTjGb
JtifLO0jX084shz5nJtb4LSSDu3XuWijVPHG5iELaWGwJhe636Mho+Duo1Sb+WLN
SLUAzwHa8bk0g07dlJcnAk3QmNPEdEmw249xNt8X450AMj5R3Ccb012Kv9o0MO4A
SDjqvy/oLQulLGNxn5s7vC+Taoa2093//2ZqpZwflnvB0sox8tD4K+phVez9Wecp
80JXp4Ntyb9cgOTlWZ57oNd7nYqplma4vBkBFexdkyArkHRhBueIbltx9jMfHC3Z
qcYxNFaRhNLgCdlIXKuqvjbAB6mGRTqAkc5OMiboXEpBlAyKDbbg0wvcFsoeohO6
B/gcuM/LjWCAWoVWgEBLHyV+hHLhLtUB30PlBdVCv1hL9RCS1weKK5JPFWFXZr5w
VWf3RvFx41d+Dsi4jFh15v2xtltwXvKNUxtu8ogGFqFi7UNGsW8R0YTus5KW848d
FDD+fX74Y7iTFbpJB1hCsOG4yrdqQJIF0hBZ4jetivTQh3HO+HKnLkKCVTbnD873
lEkhRzGhOTTk2K42IgtdNXmhME0UDXykRwNnG6A/wHeUkNg1ZSj/ARokj8816WS3
5rlDYrBjaWiQa1K4FcS6G9OoIXWJok+CP168u82LGIoAXDSXBWhnOTMY3SKt227s
fOGMmJgzZE1Uu9WGoSvH4Q9YGgzOrFEbBQCtEZqIIN4ggkN0813qLPcgV+xGrYFQ
le3LYyRgz3kD4j1cDK4zDKNCJ+DxQrrFX8Kvjhk3vjkAQHHDCnGjzuKD0LBebUTP
CMzdkveqjLBXEF5OYJy1/Dr+0nxkrAk5iJJkVCmS4lol5l84Fh9s/M6qLgKfRaPp
k94zffSxF3VUfySQW+jpssyZDmPaHnoNEK7b9CZbbSMmDc++Hc6EYaolcS6okcmZ
wYx7P8dfwjkjboIhGPa4Ju/Dyx/F4Aa7MdAEWiC3GZD+ppN5fXrEZrA8/arD2RdS
HDuScz5vYvgNKDjPxzgqvwJrgnmSYMQHL/UyksSz3H+e8lX6JCa6XYWdXUt0g0ew
GgWb1DFZqWe3DDZxLBz8NiDA1kn8q7iHfzrJHNm/S8+eDkTDTbWE6rrUkCYT2sRY
DoUO7fs/nvujUKGSKZUHvBAomOdrA18DKvRoWhW8cs/ilhYS+WdmfWkkOuxmuJ0Z
OhRpcKBhLEdOMYWLwl1BvDAPsOxTc0LlSfcVJ//8xGsQcNHe8gak4erbPA16N/Ue
6KDsi9XpQGQg8TTI5d2WX0HcRfBGui0Dic2etrJM+lKDCwjTh8k7TYMltiRqKbXQ
z35x5ydRX3blcZe7pm9TWFm+R3CRdq5iyHCx9r+zYGcPbYp55MsqCT4bA9l/A2EH
TCs5q1io4WohstNxv+UKXu2AHgjMJwviMg/lckLm1b5/DGFhXlBPY4AzUfxQ7Xel
FUgO+dutSS5MX/BszW5A7xGzybuovYgbVp+BtWUolSsIbO/rJw6N3um2PoNgj8lV
+qRc9Xz08eA6tQ5b8ycyuwdL+tEf5KJhHSkKr8Oz9k553zBK5NhNki2asSx4b5zu
iK5oguWwt7WjGwvf2TkQW4pzvPY6c1A04m2XyQbbDAD4xugzlLc8JbPHLcjPe13R
N4XFRxUISZYhd1AmehqAysyiv3LVslEdos9n0jui9UAi5vWp6VWn0LcXIxL7bbSZ
KxUiLtFhXIRFSKUBIBcfBXXu/cA5l5E34O6IcPz04en71efAUe1Smwzkuy2jNRcK
+kr/jgfFCY4gLyzpBd4XfjiOo7QbpA8jIShCuRH94Jw1Vzk9B+WrlrAMI1GANAFD
+yiRxy+CPQTnNPv2kQAy0QJckEcQL19mxOZZ0Msah9t33mDBdNDb95RtSwDuz5n/
LxkWy+xZzKZVoBpXbDVLGPUyWf2/pKd2omEonSIoVztNoQHL8n1H49NgbtjIrngF
7cmzXjPtcP+gdU4q4EG78d2JeTbjbmjpJMXccqRtyWhBuBZ/Zi2wAJTLm98FGWex
fZB3iBuG3i7UcMAjz4jb2pkq0Pw7wi16ByRNsIsqHKjLs08dSGGQOrCfckvIdmTM
Od2Y7NNlz0UmX0PKKFxDR/u4ofrzZ1ETpFL863YC0kWjXuBQKun15Pf/fxI02CZH
PylO4X2tlNoe22grhOfvPRYxzetZ9QFB71KzZXCWFHqiHbpWbw9Se5+lxIlhzSXa
ZnBWTDNvBrFCU4CBbj/qFLD3oasL6U7JVpeI4QQZNuEXzd08aCkA4j1hSb1aiEDX
1NRcTmGhbA/73Zm/rbi0yOsfH+hQSSFWbOwCB661t1fXj7Gw11xbxweYzjJjLicS
zsJCAIp1+sJyjf9C5TQoCNDvcnO/yEbQa459ue/ZA7N0z6cKPwXFhAnCjC6bOLd+
hiEg2p7AImZOHsjrI8SzRQwsPe+BzQ5dOjk8dQt9UA+ZUYfw/ERnjz7LOh+Ptkdu
FYX4ooHz4okXC8dA6zwJBcqFes5ipk2NSAk2JUk9iKbiJiYpINi58tTMvphMZkX/
ZXDzvm//JXrLDxFDOqYyslbPg3mE61gsFUozkJ3NsHYmI5lv9jR6tLSesTkwIOW8
xQGoLWyYenmxYnlW9XFwZnZQy6dGGcRFpdg29/tOtoEKt5ZNj04FL9I4tcTfkzk8
b1F7R2/KXkGhkmBLzLz/XbRNq0nhFEghTH7phV3prgOzMeBzQmVUiI+6js6bdigh
eJs9qrg7onOSV5oTMjL+kq9mKAEFm/fSFmnCFifLskzzSPZksdX+XcUuKvosQtFi
Ej6vVQuFQc0dDi+lxpttmqcVPosV2RJTzteEqFczEBR9UyGcYe4sC5GRjinemdW3
e1aXANqK16Yf0LUbF6/rzN76s46mmrGxd1fQj77BIPsI0vPk61UpzjJdnrJb7vNy
+qd168PvglYuT30cudTRJI9VQ+4DmofsL+65jQ/A3qJp/fg9KDwhLtVHCb5VFzMb
J9vSUpgcK5s0w/yBbn1hGvJPKOQseoN6yrbCCWFzOd/h149c+5kqV1Zxtc+KgHB7
vDLUz+nn5djpbOIZ/Q5fEOFxV0p2ChTCjh1r3WVgGEHuk5nrI8C696s5fY4sXd9s
cWjz2z1u7cwu9vGX2IyTzyzfRpze3VgNf0gahxrZ5UDsTFWPcxGlgiDsFleWU7kl
ysnnraM3kLJUs8aYC0c7TV1VAer5bxQ2o7Otn6MaoIR/hzCVYuown7kpFpYYDpHq
4+sBW3a9zEkSHHCW6v+hMM8EnibM8FuJYM7sOk8c4R9FqGf3QLnIStdik+pcWDYk
KBTBGuwbraRlBwbeBHKVVd0/OMBQl4fVHxbIvudyzgVjQyq5loIbMLMlBtCg4QSl
jl6DC2PyC4gY/S9njplFUWSkR3Xb6fXbIfgPISYcM1mIY3PNh0wFopLV99Hb84Ba
q1GYw5XA9UhPpbb2w3ik8oxvBE31XprB7JExtR8KTFuVR9BlCBq6bmjKsbO2RiVS
4bBz4/XCoLZ001jNSxbqPIyat5+0nsb3oXeFs6j9YJIWv9IoV3AyzdGf9i9t/Vb2
enaxGLo0Irg/uFOas3Eqw2WNsA3ahbFgaekymeShzIEqQigLFfePaEXM/aDx37BU
VVtQU2m29RfKXrsLQl1dgN+v7N5+IiGOs/6ad+6ikl2VFk+Mo3ldUD4O/KeoXgxu
I61SOmQquvwiz5l529NpNvjeRGsE2d5sjik9lTu+8XFObNbjYH1o8PUiz5Z0KnUi
MaVHPSY8/HyOGAMe3gcRagwLVgLTW063RwIXBeg10UHHu4wZO8Lw5h2EXMdEfhA9
SFwgjumEesYYMDgVmAYhxBYGpC5UkRoUGHHWxMcjgtZo0oD/a/szfDZCJbCxZU0T
55AdW5K0eVrsJZGN0M28o/hbaPgxmq2QnRcyv3yoAmC429b6olGgkcnmxoxrwzXh
xQO7th83A62fYdSUGpd6XnS+DeJr5tHPZzR6CvTCqxV3ixFZL+av2ffbjRfIwYpJ
7zqDItiY58LpmDdCYReUu0mz4a0rK7pc6cBYs2bKfWibA5etjYPpcDnMHrQFieeI
pBT8eV3EyxbMpw916qZFL2hEk00ye6VO9QFvSOiVZ9D2Rt+jUrsduZ2JrlAXCyYg
yJNbeuToGGho4G2qei0LGNHGNFLfipoi6DA1CcNMYoFNtoVDf/QvvHQDhHrZ0hz7
Q8yhaj9J2xtbjkT3hcpzZo0wzcvbJVLrH3OK7L35lkaI82qCY0458FLuqZpU2ElV
ndsi/gsWcIoI62SqeCyuXPrFTwXqae7y6zmut1JQLOPH6aXy3yHkiZweR0iYUqPp
RPetLNL1BZy+pX1XcVYZBpbXSx/ORSW7g+plr1n3AxZUiVgi+XIMh22cVzrmD83y
+razECNWh2eBL+18yGxjyAQ5k4SgeKp+66J0/DBmienVzgEtVw59nw2ReLk+/1hp
wgwm3z/A8ZeRBqWxzEQVcGsQxCSp8EFRzmP8sWkz14ScT+JaI7YC8NMjExPAtg/a
suj0ltW5KtZPd2aPMi5o4caGM0rlUaKb7n0uFKM2N+YfiCDOu+MQV77eBu5ybp5J
8WmZq/S1q7S9bVql4x7CpRj+1kQexb7zs+cRMVHP3jEuOnh9irzLdxbiGqCqSePU
e+9NgL4IGQHGLP1fFKa+KXmrmhJDhhA6b3dYDHROVO2MDDDslDBbbdgqVN6C4tWc
HSlF/jb3wSLTLpAMFc3ZxhM7d+5kdp3KQ+z4GwmZuCkdWNqw/fpgEvA5yZwv21ar
lqMOVv90t+bisNE7r5/LmRah9PCvU65bCneGp2gvuDz82GFeQ084Rcaf/tOnw7Su
uPtubIZFJvLdbMSTs+mc25897FAHQaQVyIIeXiEuFGrJZ5g5mEWMQ1jfS/BfvXsW
WG9nW5bRmvTEW5gCIckb8PO6DMwsGiiCKh55Xx2+W8px0KEtK/MH5Rd9Ve2SMms2
2fWxZt+lohqmC/eEA9ndld5/Ubnj4uPrgdAxK4LlnGjqvpBor+yIIFz84jlHBIg8
BpD/onlMz8aEM/9FaUBQSpHpXYUkB8OEBbrSPE/oO8ZzZkwznGcVDAdGTGEYMCvt
NbP6BO2ggoiW38OnGY/y7gKB9zba0pIFvhc8OrXe3MQnZm5R8QDghPbWo8JcT719
IA8SpIC7RVzrtOseQ6Sit9MFpKtCcAg81QFQ7L18d8+zRLuW17tboLtt1S9LMrSY
Drf1vzLkiKGqboHQw0IufsiN63O7Kd1CFOA83Pyd8vhflwD1KATa8JuMjoMSo9In
AljAm4Mo3aUKUy/4JWkoFd/HvNHmQ3znsNvEyyf5h2OCEPjia4RJwIZypdCmb59U
1BDEY86ZpFwhK+lf8S6xuo2JxEdcMz1WYLwAjwjNW42ZnHBoY4EC62002ZwqukAn
KF3wxcmPx50VO+l17n/w5mCa9gBGgk4HuWGbQpWukJBOeFB+hKOb+AP3WS4kM7Rg
J6jPceIojo/5HzQ7+3Tp7J5c2Qv2Q2RL48H9jU7HihGF+Pz1Yyc/gf3vQyTI4uWL
kNUiEyV6jNPTctllNOSkQ9++uPH9UGomPm77eOzHuswXGtzRi/IvENprRcStMXij
dl4GazCn6SY4GPA5wHI6ehM83judvMMXfs3/mQXyEbfebA3k/R5b51dxc97K+MtF
/TEzhe4KHKqyubCqci0Xd0KG5E3qSBYm5nGSOoAmr+dQ91ZxCYBef2FSj+yoeVBM
Kv+G6ImES8EL0Flr1xE1BFpyg6ESw8AiZuGYPSwfAITH+W2cMoY8Kr4cMZV1kD4S
14qNJUHXNelVqoZ70TKLa/YYjUcqdto0CEm17PKNtYibpGnzIlu/5yF3JoWpetGB
VuPWvidbpGJ+8l1APIq9DYL4nR3ZeFDSQ4eNIaHk8SD5KZ/nFHsvivlctrJkGdLK
MFMEX7/Y1tDxcfPZFEvShMkNtYH1Sr174pSup1xydelB10k2rvkvSesoLQuXgF6/
P+CX3g6gZHMJDkVuCMtDT7r8xYe5HtulucDX2/s1c67kZsqpr6HBv1mrf7exTVt+
mvGUFJCHg1Y/z2ObOuuWeEKeliIxp3GVoEyYYVepXMT8CpXTG/qa76A0k9Fx16Z3
NQeAoLyp1f7JlXx/+7hd2mgipc7Zc+nqEtoejxZ1jXO0ksDMNz/gqmkPLGodyMay
coIkWSJnDEAKSFmlQR9a2ffB7SCOTiL5hxLK5gPBjsxOiONg/1w4pNRddRXMbOUB
xCCf38GiAt0y38lV4N9JOF4kq1gHDY3S7XGsnMFv4LyVb2sNR92HljAas9rGCIFG
TVC2JhgnsyD7g4vhan1IhTc/uUlds752WUHXbbQ9BFtoFNIHuEXFCvOsWkQYXMLk
BOnMcB9RYZaEhLyXBTsNdKk3umURZ6pcJJNVC4QCfei0e+lmUw6B7RQL00eiqI9t
CUF6gXcZPSBjFinn9rIlWS7BGaB/TpkiwyBJ0a7E/gbCaZtmiipqcnT6CoMCsdV7
NXTR3xDjVpJmWAmYViKX3bSvsF3Zn/7xaxoGZdHJLHLtvYegxqml9OUvnPfKXzKG
xwPyp+xrRI39+sd0t1J0YIOWHdOrSQaVMbKTWY2J3Q8EN5JoerVXhg0vVMidhjAM
BsWspQ4CMvMO2KMbd8OGpWvJjB1aX/ecexCgucpk34f6Wdfdy/G9ttrvO4D08Uhe
UkeEnbgFkjAaecuGAWxrp2tmONVAQeV0XXTvRYY9i7xAZ2oncgP62vV7YghrYJpv
eXcD4FcZVE2gVJf44bRllG4yp5viZcB6/qjMHRmmkNfHSK/BdpkvxaAh1SaGnMzW
xe505dRreb+/n7qZa0dhRUDlb0mo4qTkl9hPNXynIm64Qrx9k6/aFoRD2QXvwAb7
4LXv/cNTFE89OC92tovp04/F7GrR/LfV/O2XXMgaPPuTFfsWFQ2QGSf6TkTDQski
c1NwvrBPMvFr27gH5RUguNFYnuN30tOCaxTWpRhkD9s04RAgdd+kpWcio9+yuMzM
2zOkEyLmvLGBku4q05fiUXIbpuN5OiAEbI+N3K+38+IURiWb1e1PNM3wQNW7X3d2
HnYidug8I/+AHY9PWR0dgZkxIXhqQBFPIwI86xq+gCdEH8buSAcL+51gcA3IoBtO
GF1JqudUXLJeeT/rsY7Bc+/6MSUUNO2MZLk/EQ5q4A5YpeqTjf+SlE0jWk88axux
GhMrJ8wEm9P1RmJDzGycc/BXJl9x4wANePFUFl3UE3KPS2/chhDhmv4ODM5D8hLE
EHcKziq5+EeJWkbg4OFnVCR4h1BthlRFerAPUgKzKicYSWN6yvJBrg0KWoo3FA9z
0efvZNxF5zSzHM+hE9MfGl25uSwgYxS3OpfabB7gsVTi5WyPDptMQueKhEsN9LSx
cTc1jWv132JUwXyTI8cQQZMNKuu7RxcDt/qhYZi5lZjaOIoRkTnvn56mZicD5b0x
h1nBfldhiih1NqrhwN1XtaizqYIVsidyizVPB+uEhxCGgl3jEAKueDXhQL9aCUcx
D2mhuVbu9engJWtq1NpFtZzOaCIRbe4WZ9welk9JVBDnx35YKtVddSg2+jdGPHqN
JOIZ7iQj6VR6ZODdeBx8yELRrzFlQoLko/XOs+XVvxeJ42X9o2pkCaPxf3vb+z+p
1vReHzftHSh1s1gNPO2Zv+lzUVKESz4lsJdOROyc9RHOWVYoxp8EVQH4mCI707B1
RezZUeyFod75SiL+EVu/hvdCg/S6TAs35Q7zFCrol4xwFRVKLCQzQyIH7JKsNxal
iFMohQvoBt/fwGIsqgDB4dJmQ2Ku+dO82f/vqkVKkcKAfC54fcCxFBIh1D79mkMP
Nw/3KPUvz62F9NuPEp72oqMeYHzd1j7nBiR+YQhU6fSDB+mStrax/GBN+g+SZPuR
PwHrg279c/CaToz5Xuv7lk+Vsdhb3khFV1GXxCVppNxV1JQnMdlspUpBAUWPOGAs
xSKNLMNyBNNDtRJa259otaWD1WXDP8MH2b5ATfEOR+vNt7p9xIQUjO2BJrbTZ2U6
PaLJ5XSOZcZinQTKqOMAzZPN6NCyMGDg+xFtGnYQN+j7+iNb8LJ9Jpl5oc2ecylq
iI7JQSbu9pTfNKQ2y+OdRzwHXsNNpXFSMOUerElCCD5RqlH/6BhIOKdTxuuCg2X1
x/zjwJxBnwlMxnfsMDi5KWneaM6f+n8+pW0GrtwMFGn8KoODCmL3hp3AUywlJSiP
rLOWKnbohYNXSSCCdz+T5syuakH3Ssr2eCIldexBfEToGefHYoFfF6taylnvTkjW
vNgG2DMc5+55B3scJ4+SIpa6lSI3gR1NjIVqScpe2/hffAUudAmJ3eE9QixJiqnc
YO9FU8LCCJPcFxBcKzoZo1t6cbpa6L5j1AwRR6UMPF6dPOv9YfD8x6StpiMjCGBA
2dG/sd5U2hFBClITcTotcXC82cRGwavLoVVLwEBVGubt9X9bbuDJNaQ2hCNN4Zv0
oltXiMSD6sJ9pMpHB/NF3awNbgsJ+PrDvExgvoNTBwX2y9qalMiYZOvCSD6CuZw/
nnCr5Ls2cdk6QFY6ucWLaeFJaBHgycDSylUmhmKmd5XQfHITJKSef+mQHuH+1FjC
Nn1kkQFvB52I6hVUMxTDPD6n8HnRMSICFIcrXHmOlBml6Jny+hL+zy08vx/L+SZ/
yOPQu0LABrnRMTd1VyORa07xom2ZP15NKx6LZ0SHcFn43r1cp9DLVP/q4b4cMHze
yfXUA+wSsTRvuiw889/cpuTgM+GEr2VLr9OfDMBOZnhrGWDygFWykCCqfh7N3GIm
fcXqR1mNJs8HHzR/VF7iVy3DxHqX2XjAzykRnt4dEdrhG2knMLL5WGK7Z5Dz5d/S
Ddd34jh8VPthsEt7Q2Qp/WCRvSaes7yZ3fQFHztSELPUvRHJkuUe32KXGppR1Apn
T/FXFJ2ucgPfaFAL//Ri7kiYNFUUg9G5fvAH3eTYlTRXiOVa9OYYCnMD7Tz/XClX
kSi5af5dhnfNlBejwwjJmdiQ9JMy0GYVbNb3nBCRinAjUjysyC4k1EO/L7KAvWlD
d9ufqaTmqdbK1KKeata2yimsJiXxpqojWo5DsEqLqqeFnUKeeoOQkudCnJf2xFeU
AMxTrN6fkHqNMU+be/S8gpRyXg2O6JQ5G5aVoc2R+Ytt8+zMlT8jl6WpOWNrT3O4
wc8k4iIT44ku7TPe+DlST0D27KKMk98W0GRrSzhQJxor5e3yrALBwKLCt1rnoY1W
LwdWEIsyr1NIC8JGpPR9NDsflGhKgoCpIjbppeR/NnhVzwKKZZ+9BVkK/B7giG7g
leW+a6833pIJmiLseQNWpr6q/vB5fgMLsHudde7F6Ku+O1+W7xqysomw4zCGkXBh
F1gniPFx1KlEvPSSw3q9+Kej3ZyO5nh7muQENGHgdwXDFmCihKRFEGFH8YgT/A2l
S1oSkT6o0jqyA6Abtng3M3FMPo8aHi2Tj6WcoIJtVzyybuCo9/Qf1hIFpIqFoY8q
GkSy8jusjfXcvZRUbtuFZmoBm+2b7RzN1fLiSqrKuiU54pw3Kflee0JivuhJSE/e
JcQC193RxQ9qzLH3da29NfVAesePIgeQpI4vAFsPAZpcm1GPfenGpkuY/tziRzBS
qYrJFdUnm+fvtD1082HGFuSbgtMuIxL65Ak3FB2vir2PY6lEOTpa4Tkw1iCBw3qR
5IwaA0vyMpVoqFGs7543uruFmsQfM4PpXKDVTb0QUyWjky1MBk3QgN9ubKaEvZIa
yq/FrYQa1ew3vGDdqtEuQz0AURO7Bsww6AAvPkT9Mvo4Mb2PBQ3TrwSw2I3j7Be9
joeWcWHYNAK29Lo/2VX00CMrq3KRBMG5/IyAkqfB1SDM5rWLrdC7KKDBggfs4oxj
Z1WTydv2EXYheER/qjwRu7MM0wCQLZyOr+hL9BwZt4twDRS/GD9z/Z9Zgm6WlNpV
FCKtQw+MGSCeXhonSoE46enFoOhU19vVK6+y7d4xf3cMxyOt2KajvkPu/wquJwxl
LrWQNkGiJ2qft/le5dJ/N9G+NhZgEKpMRAZ9EqzlQYlMqK1jqcNgmgCACY+0KK5i
twkIeqVErnvSeeo2c1JR02cv+orwwiROgFBSj4sE56KlLiuMevErHj2czOluSQSk
2yckbusO9Bqsz/SFiYXch1Ld8f/1RI6UhEqsfeV7JTrxLrizeTBnqA+FDqm24BBp
LZYncJrzJ20dK1Vd+FbNcMTOduXy8vokKmJbxB9LxDURK7zwWPMYM+PybEIg8BtX
VhXBQZ22kLSEAtNpF6gZdZVRSC+wqaMjaCGkZIi3JZh/Shtpia5d0VXqkaxCfNsP
CdVOqakHC6u3c1CR+nu6zVeYbYvcL6RIM5kvvre/jHdXgDzIcltP8ZAL5zU2Gzbl
Z/H0bZW8Uz9KCMpsSBJk1kHeZvaYdSX5hOAxDF7j8iW0MNBKjYc5UcTLVexCvnYG
zPr97jGHkLuxAWW8yZuZFzwz1hv/kFc79MLZ/gU+u4fwLOxDZ0AGzbqGR3Sz/uOh
InfdvhmigQkQ7ODXju7ArQydis1PVyZ3Aw9N0zRVEfA4HY0lC4/ryObvMIMyO/Se
lpECNqQhBezOGUzWUqGRrqELTb94sNL21JVlrJinqBO6tt6qh8Lx6bhEAIZWNiDQ
mhr2biA6TZW1TqhaMH9fQk2tOB6mDflfSAtwXzJ4HdjVy4+t775N19v9ctubPKX+
SFjMqT8Tr6hGdOhRbOojU3eXahptyyLsjl0LNdFUcYCLjUpNS1jCQWxlrEw43gq2
CIfpdLpagYVzsgjEBqM3uV4tUsY16RBLMohniZ14/xd7fOVpHOmI/J2n+Y5QOktM
Lpfn5pqwE3dUXuhQTtBXDNthYZ18+9f5rGJc2n515YTqwN7Tha9JoFwYq+NVPdZU
cvXwKep3p937n6DiVMLKP2ZyduusstcfomlCPucxbqE3xj9meYQ3yymZaCTNIwBR
+ULgTR9ZRucEdJI6OkRNe2Cp/Mt/G31ucIJ0KwGL0s/n74UGTaS+idqEwwAyI8nj
vLQolsP6UfpbZFKnfZ7JGaeZh8Gwj2zMW9SDI15wVMnCCLsVyl7thhaFzDu9c1JW
7bbutXnqtXIhze9gdlY28WVGre8D90wCoVUD43NSPcPzODZYiGmPTIQ7RNBwkd2g
MD1aRFr3eQ8ppnWTCJitESpfHRtFTreZaE4M/7ka/pHxbndIpyBr2MAh/dAlRNNj
X0X0LDgThZBYHzEb9P0GupQ6685INQjpVIJ6egq7gSHyBMr4z/vLcqRwEcDUDKc6
uIjRdvjJbAE9ywbSXUP52SvXwmfGi9ZZnrIUWH3gHO34dk17YUd7ZZllpLCuFUrL
JI+hA11lx/YBFOzlr0ab1csFFXybJBESYHjbhbO6yu6PzYzcXP/F4v0DQk+8kiJZ
V+NcaRRK3dQWunx5ZuEedFsTsCNqRs1mdjGYdsc3CbufGB1vPjAZ3cRkN/lMpHz7
sKEzLiNNouyS0CNl5q5fYPFANBP7+9sStN6rew+L8EGeyh+ra9T44zYVh7Gcu7Hq
oPuXCfAAKsK4E/Hbzc9EkXVW5H4eQRhDblFwg+cI+Ho4v4AIJ8bHcSK4ML6Vb7zf
MQxvnYLzolM7Y7Sn8CXnCd4ZDCovN6KESi1dtpQyX7Un2KbRG12nmv+HCEIMdxa7
7lRq/tP5EJTPx3Cvn4gzVYbQIqwBhieMjZSxrz2V3r2Z740ySW4EO8Rn2HtqqCCE
353mNw00Z8RUWNpZDje7TomA3CcgSnhF/lpXCc6nAkDWdCajwrzNlHkCOYpW/CbU
kpUpScivxvCkqPe3oGFcob6hh+d7QEys2k3XFDS+213PYGLq9gHeyfKNf5yhIFl8
Dt40abPNI0Jifbhgk1V0puheRUhdEhq905LqrYFDgsrHyommrSvMAJI2p0+8cLaD
loXquzsSyshbwoc9w8PRs5krMNCbAt+NqwIO6syR/ZVFHmGUNa3K3hKV1yi4E4dL
k4EAaFiojIFgb492KjNJU2MqjjZYQNGKXKu+a2WNFZ8heFhQdrM0pT1ax3hiy0TP
45DeQ25IoAChVoIcM2TajCqaesYLYHn/51PQCy/ePYpd+PeVe81OMM12CctmlZSP
Kh2Ca75d4Ifn5kZuTC/iiYQ4PrrbhAAwvgqTOeh625L7/MDQ365+PmzWd93T5cfy
KZZYQwnfC5gTl/U3xnSHCB/vez+OItxuG/wcEFgCf7sF0SuMup7l5+6fvC+mZXJW
Q8KOlO5piJsAz7VCIgdh+Ln8os3PjtZuY77G3t9RpqceO6BLw5LFBytNhSxfajf7
IvUkgQLrur6+Ip/LT4P/iKt+aaHVbDpaz6xiCbqNfPLergcx6YJC4u5ykw5yZODQ
Y5MICNK95kHdN6qzjoAjgEWotG3fpZiDOf+318w3vOiHOXuMpFHPvwsjuKhvevvT
ubRfHTQ5klx2lWOAB/n13h8ghLC9fuMDhS2y/KPBaZiGLYQCjg4QPnSHMFZU7Jly
85AUVpeLk2XQxGQ40nUpJ58W+m+7WFc54VtiCavINWL+u/1YzrI2Mef9GcLm1gyS
03NSbStPCTuw0lUQk9jtjx5kBOThBA596rJGFGC4W7IATqGjT4IQi9/5KkJq+qUL
9W+b7NtS86AS1s+7ZvRA6rrF62lZ26pJgl07mPnXt95/uc8t87HUSA6wAqg3oEeQ
lYXF/UvHFJdMilOqPIcKz3iCOygxDbEcy8OcYIW+PtUtV8LeIMtI3CCqEy/fOR3r
f1UyrCGT8Zm+PGsSlI4sxK0GUwUUNf39i6T4ZQTi+2eAm9rgaA/Ptppu2BrJScmY
TC5kNv7s/Nw1UGuV2LyI8TTex4Kis5MHS4drLqD8AZ4tiJSOD/nXrEH9P87MZ1kq
iCqZsjUy25k5qCgc070TKEq9lABWp9fc/5yoonoO7eD5Jrwr9GEAkRvpOzzzkJEt
OSF89CFYASW2T3mduhgyZ43G2rFVkITuhMSyQHh0Ugw9SQhyehiDc5A3F+Jao+fU
ZBkfN0jjs7tmfc9VJ0bnpdLNV1J5Y5qXAgO05C1ozrn1v5Ko7kZ29P9gniJZx9Mv
yRyZhlWSkO8+mInaJuiZalXvl7rZOnVt1upJvw58kcVfk4vYjy4+UM/+hiTnMFv/
BkPLeLyjSoMHt2RLSRkjUTliyY4KfLMY27BZTKqsaBIfq5Oucl2l6ElRbGXTWEcK
LfgtrIr9OKh0gKeivDRyxkhPSv0OzzBHLELpbkPAPRFf/w5m881C7I7BwtHrK8RL
Os1+Jfz8VYHyS5jtXneinS4w8BOQl8htoTNQLQKhz2hksQ799zszlQRIpmLprPQY
guQdeCyvSu3TH2JuGMajKsTCRwO6BjKgOaNn+M9eblNL9NC7YMTqq7EhYPIyn76+
vI6Q/uel19PQfpQ8rwkuIfWXG0f7SvWJOhTHOjGf5YQRy9ZTfB8elwVZDa5kjAfI
OkkNpnnoJEDfcumP6wgkqtmXm1QiOr6Mccb6IYD5mkg7uhjh4vlduzO4KMT9aNKC
462A+3Q7Ba7j/t97oKi2rRcUSNy0Lb4N29SWGvqmH2+k+VaC8GFvIYk86lb5Ioii
2gLSV++mwIu/eIw11KrE5e4ckscFwROPk4G9uXpNd2w3aS1Nw958u9H97hB7T3FF
VCD873k4kYD+HPcNOOBwgKuyYd2MF2rXke/EVvYuFYD3rCqNFfuKXBNGYLYsxq5w
94WyzY4YaXSfoIFVlnKWxqSkp1vyhQdm5EFXUTA6uN7FUWUNhPjon+6HkREF5S7k
0Z6VABYriqxwQowV4vnuRrFKmG1C8gepfFH2KLghiFuUb2Rm3T711hCoMz5d1lHf
q68jmwMTCOvBK9zWjhnsgmMT1ap6DjZVF3XiIWlPF1CmBNrWp5vWXqnPl3Fg7CFH
1MxxjgzWlvlDL7qgy+ZQLCxfcy6cYFd/XW70P/p3uffPEbbh7bWenxBKsXJPaYQo
nLbwMCrLSXuRBE7Uk20PXQLhMl3efSsOvriM9MYSplxLMdH499iRxyKbfC2W3dha
357mQ1cWJ7nfP89mKnlNAX/0IFUSFCNAqoMO7rwqs5r0os2a7Q/1ygIJG11rpBuN
LEXnguGR3WCw5RU7Uly/NS1uX7jEvCorG6NdTaXLS6pcAUCuTUCjG0DYVPXrL7Nj
DVvRhs61sVzt12bqqta1STArJA5/tBlLTaTzYJ9yZ8jqJutaRHWij5njHrZKbec2
ToWAqEBlRfjPKS3AuXpc741ubrCDHpk8HkgsJ0IYkdFcKAJNWutlu6AKLameDIFl
skYKbg6pbUC+wVwiH1aPgQWWizcwLb4NBSCC5veOSsUCH5YfjUpaZKtMT8ss+rle
LsUnUXuUKx+jE67QLK7ZdYeFHRFDHwaOvj+Lg4UXUFvw2/ZCW6HlpP3t/c8Gkvdr
GA5EUruihHfXhyB5jS7sW+9o3BoTU9fEPFt9dQTK2e5Xa5qc3rEWnBlMD1aH4R1y
E7MRLsOW46iR+NAxOPEFr1mJnn1RBrBwx6/WwmA2CbRnZhVWG8p/JQswYGmHFlec
Hhnwt32TW4JPDSesBYgc5ukiSlsfmLbxuvFYUgG8+DNIPrlmIIs9/LTAcFW40aqb
5v5BJ14RPmHiSeMxdRp0uzbcXDWSYoyJetsUyQDOX5xkhKr/6t2SiXhC9GFo24vI
yvpuUJcArxmnkH7MNbN4hqZ8q6FfvNdNLZPFuJf8C68r2pVGayB8X4jieCllIKRc
UeE9e7shJ5el0RM0wAqqdE5msYur/81mjvFGvQ+HpmRqs42PzRpHQh3fRLrXWkac
zh3fx1rYSWIkaYEPYR2uMzKVRgxdz+WI107jdKSuktZgBxcB//IP6ODonuNiimGW
gFMBsu1MX/XttyHlTli0iusSoI9T7enhe8NSkLSYas5X6EMJgIC9Tdih5v9ikDD5
YDjq48Z/M+eO3f0Fc5EW2EDtDCszb34Tw0lKCn+vVFcmSzVduwAUVJePaIXuhKPI
opRSfWhIpBp7OMBRtJxWRpBSxyUojgD+r/rXXlaD6Czv+8mCLyAuA4glPgmVIfXt
jViyeSVzDD4Fv4U/6UmXjlDRvqfojxaKUNG74PNkVCnkLjf3jF7yjzwGE3cdVaM0
TaKvrHiL4mGyHrnX+7+c88E23+Oy9QOPnRbWd0qz+TFyKazriOEzJS/qjRX/JlH+
fAGnJ5paFFYtrOLOSHSDa4u7JBE/yN0AP6D200jCUXJbJZmjFlQxlNi1i8LD3kGD
PWmdwfdJWzBS/cKsl2hz9f9f1G2VEzsnJXspOVHTaWPWR+AuUSisFq/+7YCRlrl2
d3BHuiHm8TZ40XVmkjLbyIDatRoCwITgqLlOfs1Z20psaKYKi/ciCc/LpsDP+QKa
0NVHLkHAUmwAySi1LmmWp9vzRs/ixJlW48UDtFwtKg3UdNBCt435V05foPR9HwLH
H1ybZ7+U620Dz5LryrEyoMk8voraQ6+po5OdmoIhpYxI3xA+Ai/ESrtA6hgAwaYI
zHlwPtroZm7Y+NmSd+BBHP+TYqt43hAZfiEtKUoHOcNNebZJ0ZHeZsQmFRTPziX9
7hceGLk2KxPRsm/vRBDl1Uw/BcVpjiO1RHc054qC8FUJRoVbZouW2repNjF2R+S4
uGtBiKNr8EKe7GaCkDs9d6OnntxojkIZXpi7uJBd5xr5MXEIPD+CEIxDuwUnieYt
l8sNK7La6RaBew/Po4X8OynC0W526ze2IquZ7CyUVh/42Dzf8gFKhfv2q69osMpf
C7lsuapEDcsGW7v+Xjqct2dqMsI5O6ZDeafZ0jdo+0/AqfJFThzrHbjurxqU3GmY
yHkh8AG0u7nlpVHBrDxQQfWsr3KDttn3ZC7xN5dFdUrnUYGbS1kw541EpXZBK3Ed
+WZXSGTkd6VL5udIuu5aPyIGoTC3Y5X6FC9ftkIdYFYuz8B/Js0toA1v7ft6w4mv
4sheYNiEfFGXKPhcgf6XBTW7nQPTU99BFLebxmqejk8/VAQ/1zAmwZxDhU62dpfT
insd70mpfl0F/GolBsAiK4noI8m+l1688K4onu9iLkMa0zl3nMvpHXEuADKnVNCd
DSoQxhEmm8OfZis4YxY85zL1sO20xalIHODknhWnA8UYjO6IRnuajXiNsxSsZi+3
0CCP9G86k9fSAnNWBLLbbJnSpyPVdPN4kggMbOCtKTxzulL1pqwsBklfZwSLCsJW
5kH3Qfv3NAmTxMqzVLeg1gayDk8dobKD8dXCLO+vvLlQHI5T6QfmNDM3ccq5we4K
iNLu2ZWOYhdBrFGik24AOEobB5UGPGGOBoszLRwcLbPeWos3UwD6HsX+F4jnQmiH
22zHnhtAYrpU1A+cLYd21RRiZ0kzFyPQyKaSkJecf7UY3ZVkNr+lzEUEj/2ogCvv
wV37ta9T3Cwev6DKKRUOk2n460nc2jl8an66zFA/E0z7AwoCDTZVkgOHgv4c6V1S
k/TdR7zvC1LrmmuYX6zKgE3XymcwCFl/RbqgMurc48U+QEWQwGR/r9m8EKgvbaGz
p2KfvZ2Pr34q7fnu/3sXyEBC56gIu2jpia4+dWD3AaEw+XT5CQME/bSCPcROlNuS
fQJ3V8dBIzNqqeNr4kSAH1y/mXLeMmG7tSMPejkoP0gYROxIru63sQP9EXCgFDm9
tTwSLulgpi41I1T6DW92puzFVnHwhkg3iCzpsldaTdtAllwDvhvjRhEYgiERKnx0
Nl4MYwd7fL9erC7RZAjElaLRlvR97ALrDey96jgw+L0iEsBNbOsMPaOCn2DY008X
wc2eRJSCQ4WwVPU7Id60OvKGaVZ+XCYFyoZNvt6wIM3sarPnX8VliVbV64xmOq9w
tFztmzSWfVMZtc4AdvnwfXS0eYwO/dkcI/SIQ/Hg4yfUwkds+p9Atw6RPRisqLwz
EOOJC7gWr35WyGMuPFFAkZMtpvq5wVIpR/7WuR51P8TY4mflI+aJ25kztwPgoIWb
xGL1Ep8W+Uq75/aQ9IoAPYw6f1Unmq4PBIg6fi1dnJh61ztalzCzafRuagpfJ9Do
pMLYkmon5xm6ZpgnVcj7DTjRzgIuIZXuB0ugOA+hQRhXvk36bN+kp8Tl0wB/mSe/
iF/4NeA1HQmNoTmUEJThFhFqekXf48gb8poFWrDPJNCp8kAwRS7ZomajVwNMuFs1
yJPAoHYbF4eD4elID4dvbpJFzo7PFItzlbyn4VvB8AkZA4Ko6+nrFbU9tUPldYCz
rdPM43Wmxn5u8CvIPRmDH7D+rU5lEMKwq1J5ntsX+U4kue4RQMaIs7g0Y3W2cZvJ
dspTEM44AthdUPXKI7dyGqHLo354hVAI9y/uGCbC80NEoAbxz1KlcR2tTTzhKpIU
dBAxB6Tp6LqApt4wBYa801+KV6fBCCnjb8nw43UbtcUlNmhwREXdpPm8RN1Q8eE0
J4JQPYQ2Uh+mQu6xecp/CluZzO6dJMQi+4ILuL7iVP+PJqPFkH9Uy0U0DuEAdkWc
TeknfTUlPUk41prM7VTScRUKo5nJCKqU4GHAWmQhtlZEcp2pEon8FLC5wG3iECXR
pDgH2Xa4zbNPh/Lp2mpqsTWfoRYCL82osbGyk0guI8iXqqkbVqDBGKMbWKNcuK/y
BOvwbm29Z2JbrxTN1cPmVVgN74cTDolSWfUc8i7Y20vaFIFBQFwH7TWkLxUU9T5b
v32AVOXZVdidgJ1Q36D6GXeLHieP6sUMP2pz93PWn7q5WIDvQiCSHg3VhVOo05W/
hWwOZapliEr9A/acwkwrpBKbeQtf9y90ilGYGXp3ExPE8RO8shi3EoQEsFN7jhIP
eSIDxcNFqE9+5wUatCkcAHzWLpjB5PtkwBo1gl/w7eRjOjT95VON588rMPJb+Vy/
JIn/rvZMRL65cvqNr6Rzw/hijVzDC4PX7q/oOe+LQDdGHObgBHN3Cd6VBQB5KUyX
yAKKgS+u7tMZv1uhI3rEyKgejHqFuR+0Knf4svsWTHzbjWIm9xi01e4cuRyTtFPw
3q3Dh+e50JwRJeq7UWXtAHE1eyKlsUC8tBNoCxh2lSclSCcPqNCiHU4tNm0hIzyD
AT9PALNz9ME4A5yqkHgbIEv+0iEo7pE1leCHkNBkuRHIJPKqVXFIfhkzhKgUUq4K
B7xQx+ylNn6uK6XvMmHm3IIIOO2/lIQBCHJZVY6ZfSaEydTthlBQH9zxRNOSByo3
QcfS41hovdHhbSHzkIg0jtRxu7lMsaGCl5mUHQLUCGMDbv1dTwwB3vH9dZJxEror
sG/ec2kRikii5fvw0aTF2UuAiaHv1iayXK8+DVRMQ0O5ipsTGtxAhy80D/7ln3ry
svVtl7EUlQQQtiBTyW0RJnXT94fOkJIV8zOfkV8NiZRLPlkmNzjxA7YwL47FghQL
WJhivLZqvD73VlnBNPRK+eTpeBnGgu0gOmZOyvyqQzr5exPtxBzgqHK+vDpE9g6y
iii+JMO6PU581Y1fnGUxgHomUXU2Ju8eIDFmkiD+GgZHj+/+F7a4S+J70gbr26PA
nxroPWU1suDhibzFSZl4pVadW1EbS1lQue/vjGQlVD3/KRZt1lDDK953N9UyHGXy
JXa8AyohcIRqDub9O9XZGSisMDIawqps0dPYYyayIwP9DFUpuvXmBrK+Q3zYW1MQ
jFm4fcZ9GRmV3XFI0hFG+2zArya9xfaFtKBQiKz4G6Kv9VSqdHGN2MOngBF/cDF4
2oTTqXB1f9znucX2SSCLVfVtyGoLREkzKAkS9GlR61JfkCSofcpLWKIHCETxyQqD
EHE1cJNnmg5MKXcSf8tMI2Y9NOC5+4dk2a61xDxt2916DA5noiAnUASWr2cRCzdT
OpkQBG8uHKEW7zLMYNPxgXjfM4yZeKLqdhIh0k1WP9I/mgtmPG69uNO4h0W5Rs7M
YShTTqzwnaH/6noC6Js9dmEEk6MV7gHNMBrhoq4JJmUk0rRV0An1oenqH1smo2Bh
qyeJI6eWLfF7PLDDxGZyuNB0YaIeE0Z1qzNIOZspSEPwzBekFJlHliz4ycRbAKph
aDs0nEXIYapY+m27irUap5LcYBMVGxtpP2JaVIJugUjCqUuQf+KV+TwlYgJeSfdv
Z09zDsAHbWJRteEyuTqB5imipTzdiWkxT/GvDOzUAqscOaRhYYF+x8K3xD8YsMm6
89+sJgBrYm2wcfd7rDUCA6di1ENuY2qhKVhGaFFCjA9I7+uy+0RTAKPqMTdE+swW
iIK8OSbt75hNMw5lcFSVwly7d9OCvdfdczwfVsE+x5EYBq8x9ABIrhbKydvhcuPu
xDZOi2tEzGZ4SCywlGWgIXImUY1TSl8uf+ULlVJGPq5YvHIuL3LQfry7m/L9GJJy
rsb1OeDfbbqDXIgCgzv8Hbiwx7nYOR5VC6fLcbkbO8imXS4Q2o2Vt47oSLbmu/mD
Ux15rwC5be9vJKkra6TWqcA7AmgzzPZg+6tFs8a7EtfaGKAcC4szWv6aaoWnjXcf
YXTkitpldn6Ib5Q/+13Camz3U59o1EtlfzvzLeJWLK+R3Fn+QCSgNaksEG5TBN6H
mmbQREc0yBSueZD85bbLOAe998RuVr/v5I6gQ2dmeD4BfoQMtKOjnE8x2IDbd/+7
d0+FSH7K6Q3MdXI957yll7LoFKjIfL9/w07zS5RseKpw73oUzyBdIRfyrV1FZ5ty
3GCt7Q5GXxiMKxz9y7UG4rzgszfXOqGdfF7duQ3/6hePNFBiBnq2Zd6AUacnwVXk
AApnUxW2qjRb1FbKhrH0J+uE62Q2BXVKBWGrzQKp3lLmXnjBcMcje5DfLG1/YAe4
bXx+o4b844lNQ8Fe0UEFrd9hH2eZbhVMmig1eusZOjShjFu4OnAdxcFLZkzfJegy
Sdu2l7oXVlcPNV/TEtpsbAS03QECYUXNe7Jk4n1S+XMtHhBQK5aFORXVD9H3JmTA
YiQNkTsPHutAZ1Xvk9A3WREkWEiiJV2CIoSsAChZ6SZ5GONEApc8VIdLrlv9LK1J
KvY+7x4HtDR/wx/m3GieJrULEGOuHX1uZr5fpmJoVSwyacFmGDv/KvpZne4zszwK
JD9I0pq/hxI3DyOpR2MjIYTHqxFU6QUJrbp0pW/u4KDf4Rr2YwJMnxvLD2zCWFzc
JxE4lDpdSRUWAeAMkzCHMYcFT5+wzrhmfCmEMVtBh4EAVMFqfE2CBoOZrmQeRXXH
SICg+CypPLcOIsY6IJyDsPhsVMS+hHi3VVyqVeyD3dGNVscUSQFELyQFE7imHkKo
9yWZJKIpX4v1VKyrJKn676PECXnF6TlVO1SvpHI9//iffbJB2TUFC2RO7tDGv2Lw
/6pAgtNClki9W4QUSRvrLiLt5Qn7F/icdjCTe2hc79dbFUm15W0TMqx7M/CS92mD
9Jsdl8G7CfPpl3KZmxYcc9heSYTIPjvtNbjaVSxPtv3TehAjIBywjczkWxPckqdh
JcjzkW3ZzaTvexilXf2WlkYBXMoJHeyfAgcZQC/eJFCtoQlvImmnRiKWN/JBj0hl
dgVeORYAZqWci00piT4t92GiB7IxbwaOF8P9JnylwJ/SQQMpwn4JpPvY4DMwJwbo
04tD15fD1PNX4sHQydnA6fY6KHyKmGgzb/md/mWIanIDu+CuXafHZ8rDu9FImvPz
nuXWTqQLaTWJmzzrLe1Tujk6vmYbuTVvlRUyKdQmjYOsK3CQPPC/urHhI4/Qx6N2
nR7kP5Xpqq8l9boM3QZRyZ1LEKtveDGZljlVXso50yKUplQba0BUAbeyeXTTmRXC
18jugm50ahYPGKxEiqp64ZbBaOnEv7ulnwADbcyNZUAHWMzGRGWpuF8hC5gYF+G0
HF0N637ROA2UvYqnXeiyYbtxwAei60KUvQI8YuR5WIUrOhdXXrdEt0FLUsFv6NkS
DXGzRjcPHCXnPr7PP4nrOMWoTKNZ8tR0leiD62V7AIsbSmHzmIJp08JDvWRuz9Tz
YDybP7H3bwYOF4p1mVqVlHbUfM+j/Tf8su4Ae14y8NOORp4SEi7lk209QNkxlTtz
Q7nsmtZSfjfPStDk8vQPbGIkDmYn+T99SxNMgw52ONIFkSytfZqcXASvNF0uTMLu
wwqSUPt/7rlTWyzlmH1XT/P7aPry20EenxT0kyvo/x3KJQtyzjajPWLaJ028SPhM
4gR65kvqRyOKLS1gSIxEyvncKY+Zwo4WYQhwwLS/1AjhLAk2q5zOmDjhZAtXi8ov
WuBRgP7YcSVShK2GqXvo3cJmKj6YwkOmtnWZ/9lnNktrz8ABhPuiL4dDoWQA9W9V
3a5HXCf+LA6dwXMETFBHbtUrra63xDU1/jB/khzFwllcxKcfZmw2l7MkVQBWNeT/
FwX7lEgQdX9eQlzxjr9PVzgfCxZP/kmRtcDbctE/3JGRTSl+qtP9XhqmS7FAoSMp
D7N3BEvAy/UGXYhs1Co5u9DAnuYC12sPgDYyNWQiQkPkBrcwt6HAZmRDsouEkTSK
RZrOHje8UyKT6AcDAbTw6wZQht3mgbceSljci5S0MJRL4aHrcBUyfABZDY34WrM0
2iSQawWy2qcSee8bh6dtpSYTBgUBJ4mZ179ozdfplci15ji2P13KSsA3fRebPZ1y
YTKGmwlqYw4IsdlS8Q0UuVpWybyQF4smF44Dj6jBoXXvt7rSg4L+4K+bUPryaOt5
bBwtB8qRRUEoq+wX0LiBa9lCGPjMy3MHOu+x4EiNJSivRS/wiUsVfYpz/Ng+UbWw
yxK79r0YxY4YVvtb0rwPCfKzONVRedN9ir/LoWQizi3KZCE7REq3KW8xA+OMqMjp
RufOi+LxXy7qiaHO+zut8au0ChFeCOzawZ+EI1KD8o2tmdj1KEYUphe9HK/K6q9m
KXzIVPAY+E8oeg4Ok1F0scW/6X3T0oCCW3bXwAXRzOau/EjhR+9Y7MmU8xPZtt7x
8esUfo1wbiHLteO+rGefk3Two5nyDy8gpwymb8xWbb+E4RTz+UrSjbH/gJdY8RkH
3piKajWI2ZRu12kHi+c88mffv/L4JsK51PkknLu5/yAMbUT5TIFubqkvTTtjtecF
+s4PSb4iJ1UxbljZyCcJTfkypJgVynIGg7LVACgHJiE6i5auAshRCfi/BKqGqkIq
ztOJNZAWrNiOqb8/WtcNnqnMw13ZsUnL6YkDP5qlVxxV4W2GNfxiMrZF5FhVL2Al
lpy2e+3Hw2m7fkSI4F4RAw3+oOAeFNa4n+14MNcdyGVr2mKprnF8vGdX+2+2MiqW
t2iTkz2+2RhWDikQYq0LpK54pei+3Nn/PKAivu0JK4B0CmvhlviUgstfm3ngn109
fQEy0cHypoqrSQzEJ3fv/iVEbu3vZzFe2/QMYONdinYoTjzIPoAKHBoHaA8BFyk9
auFw2pkNok0dkCB0GptgXW4zR0I/iEgN4/GDD9jYYXT8U6Kc9eDXlzQCLXtP7Xet
w9xFm0zRa8IcGT8D07ODXrtOSh/T7o96RkTbpHqA7my1bULe8uyQnRYLuKh2ycO3
o/Ylg1suNLKC8j11v+A2C+uOU+X3W00eubNQkOecgPE9aDgN3sUzuM6luLdadQ80
uadMh1gaQdrc58JVajvdAavRVhX6Wp5u90MtVT55idw1zXcvtSMuyYNcTg+eesSg
CtHBkZUWy5bkF9eNrOh2R6GC/PW7Seg9NCGZFO7TqnRtQus7G3L7QU94d4kNCyiN
Aw0JtK4LwPs/ReNt3A8YQl+zsmrsFBA6hoRfkjkVgSZ0smco7NkiXBr2DvbcaFLW
ovItzVKtHe3HIps4/l1/k2YQE+WbgzdItNBh76KB1LKtM+wvIK4KJSkUulyg8nW5
t/dckUey9+qe5eoLwZbvWvMV5XaWazBllpJe38lmXZoydjJb0JznBOE0KmQWwfzA
uhsr60xIY8+L5lvMdlUY0JmP9xj9ktCDK0Q7Ysh+qdFU0MjH+PsCYcp6RF34mYxS
VOAtH6uEXlJ8eq5VWv8wcnMduVRYco6x07lB9qqsbtluejarG76Ey7rEtJE7UXhx
+1hQrV8FXQoWnilMtT/5rrq56iacdYqbGgkTvutMiIjJBc4lBCAldrHb6N8TmZJR
8xaWsB+1ve2M4MJzKZWyQvJrTfooCj5Jks3MVSv47jkrJGtQ/rTtRojWeP3qYJwE
4bcKR+UFIJRvPyCvRAjG790InNgZnIKsMtAqpHoq4Jeqc+GSotoVBXM8gWHIjh47
Hkk2UbiNF/HOzRuWauvvpJD4Lz01j1t4Q+46Bu7ibzwqhuBxLBH3AHmdTcas0I7+
zev3jVRu2WVVExj96IlRNcMqa6FJfXKmA2tKpGxpIFwyRJ0vqhjvFa/fsF1vEKH2
NaHIpcJ2AyyfiIe7TK8uDnoTlQwY8vFCKHi0Wxlm5J0tO4Z/GQczvKLSuxyKCP4q
JraZ+AklM44NToTDwI32xeRAZQeOOgU9NqN0QMJ4EgQelZTX1MNdVhvK/5xz09Pq
V35sQWB9A5nxbsqoxpTGL6u34DW/LECmATddEJSXMkmkTHXbLlG3Cpfh1lSehkob
1JS+L2AU+Ce0dlfq/DrzhAEbeSso0iIe0e7yfSMvkVgBTilZmGEyfJcXFWqXgJAM
G554YC0jTDe6HXG8szz3CNaraobDl2Ez9KUWO85y2jHYv5bfdOiTsrJDPnPkb3Ij
5HGZD3STYH8utQdSvQpt/WjYVcsxBfIg4XjfQKh+jkq9Q8n7hgixG5eiZtMZCDGf
FmUoQeNS0RgRqFUdbFzHZSZBVDCSnbWlRnr2L2sMrag/htb8uQZgi3likwNpQKl8
rVmfb34RdZz4BBUPHfjcsTaRBIdN7CTbmV3q9fNbjk/9N8P8NM4KwkO0h4d1oFPL
BQFVUM2+Ub0ynazMLHs3fEk4dUVCH9sLHsdK/VbBZgXLnm2s8F6rT5wjOm5bYOlp
OlwD25S/VfKUzhRGElLcUxqbcX/IpoW5APzGvY1mvpqpkOBC4S04gG5Tn1FLG4EQ
Mjz//TGK8cIHst4cymsnlwQYLbPQqc2cwYv5sGun8+OzZbgi6HAwIEtQV9YPhGzh
Rb0mC8UUoM4jfc6f2gvXEWrkh0tRC6wMQPSu+ShdYdc2Ym4iXNxcttWIrZ/Kmg/1
k1z73Z4CXsf3QJQ5JOlfCBJbl72SVgsZGJOcm0UgrvY4L8eDrh0aHJZxKP80I7Wn
U61SfMaqhplCOma07+RzAfY4vNtyhhdaPLBzMEksl5e3L0ljqwBNOn/xn7rH+KaD
578Dy91SPiY7zomSZ8rRQqQuIQh/RkhyzSA6FDDYI3zgjk/lx4roOZCCAxV8G4Og
F7syGsL+pWWUWCNxtx2ZnwYcrtHJcPQ4buqXkFQpYGc7WGLy6ga03pL1vNME7uXW
WYF7uWAOezhiltXu1r1cGRUiqlZi0Ufp+N8a+VIidn83i4yrvf1nDuODBr4kouoB
WUhRw0EaslrP04a37TR0Fzp/6awHQUkJL0F/mZFfOiRtqR9GPCgorjUNioG40gXZ
EF7ucLYi69Qijrvh3K5w+ExfFxPu1EenD+vtKX2vQeDtlJxBVm5V2Qa5ubSbojS3
BpKs3OXvqhtF62DuLNrhEzitie15TuOcGaYhbmel63Alf7qr7pwJDEo0p7Nft1oV
arlAK/7oOkxDDUl9KNV5GX3PlffP33uz5jbbFZHabqY8gB6zQuPtOIiWc1VfbYj8
7xNga8DZ5ckESDC5YnNLyBXNTHnXcHdqV7iL1hOl9MVTk43+bKrDejLWpaQJ0QD6
zzaj3dZzSk90VgVUU6SMuyS+3vP7luJGid19ZRPesAqbitd6Pf0jPTZLtInyFnyT
CB1fTAlwNAwos/HMqccPyf/rB9Ma+h2YphHOgv907gjU1MJZImp28Hy3O6PAGCpc
KeSINzlF5v24AvxZ/1RRMR9Ex7V8hxo/QxPetGYA1xncIvosLgKB+o//7ezBgy8/
gJC0WPOM8JHASr3uN91fnURInZ7gibMbwEOHQLyGFuRUEFM/ZxKLkWCGus3qOUic
fbks76X+9wnec78/JJ3SgyAUuZf1tLb2YjhqyxySpryeSkvlM+8hmGB2Xqpz4qev
UuPJ1z9X7qHHg0bYclUYXHpTUm3yWQY/fIdi26I7oz/2gk8AiVR6jDmPS7odzA1e
g+/hv6M+IONpFkoEJtnBUliwIQbhhutMS3aXjAdbyFSOdETC5ueu/YRDHIk6jBoZ
SjTeyEnBQXC5cReK+DkOqM+OKkp6lEvMMblqEdzO4dPtrmYew1R4/RLU794AiTZy
yJZHtjvfXWwfN9LSuLqS8mFTcvewXTQoACmlCsuCbFauO29YPVjz2CP8rSs8ffww
/fM7mZCV7/0vDje7vL53sOtjHh7yBu+EjxOVL23lI97YFcK4fKfQS2k88NjQMXOs
mmlpAq43aRHW/3uUZGo/9xHbxECwsbGm6IDwBve/Oy+5Dfq7AREB9VAGJLpZ2zPc
ivkyznKxBVoHQQWzUEgYisUYnm3iLuzlI+OdThfgXbn1JjQ9TNgfarQMgGIYf3E5
rdtEYm9CS0qLCDhmq6WFiM3eJEWbfWlixRGKw3HN+S/WAO3zKkc6jJ5cQ/6Rf1eO
WKK5AaqFp3FHoYkiY8ah82r1SsQJr9DBedhC8XG4WPPN60urOEDif9AZrrtCjx96
a1/7kUc4XhQKuYSAVqsncrbWgVGzWAhOnxCZxoJD4X/ywiMEVYKJ0sZ57hUro84t
wG+VuQSkT4zeCr48p7pLE1iIrgXaMo3UgUaGuaCK9oFiF/U/9WrgMRSj9inEDehU
YTHqw7Cm/icch2RZQsOEsVwAsax+z02111LJKqIsmIHToeIasOvTMAXgEznAwE67
CJ44tCrlT/uKXuDiMFUYve2qSplweIp8u+TMKkd20ebZYdER8AWcFaZA3VDIKUrh
fxVCpmdJiQvMlxF+H8zHpzkQL5gdaOltsGZDHdrQZvJCQiYJWSf9cIVa+NM7aO7R
7awJ0xAEk03XYhGk5RUp35lZQs/jyROWovcVQTfb177rmCuzcxdPvOFtKWcGKb16
8J2mr+MIDWU1TSU9SYrbj5AbHTlhPQkoZN1vZfYRl2CXH9I/gFBXSCXcQl6+AUoL
dGfF/T/tYtpOSd5cMK59e+i9kdHhgJ6hIaZWKsFwtIL0811j1EsKtfGpVqEeJ+3F
+dQjZG8gtUdupqZUfeWvVLqu/E8kdj7R/tyk1BLyZ/7AUqSBvQwQGTf+N57JRdIM
5y2E2VkO0roHXIR3gzQ6HPLwcRy8h+BA8AnKdkqeJVH/5uWbC+BfNbgfqoZgiy/6
3jIyPs9TG1cppLWvKqu4EfFp77MrI6moitXhla34SshsqqSPmq30wd4Ah/6LYFSV
yGlq6tAJ4e57BOKvzsCVvPXG0y1C84Gl+D7kOjeexvX7wmxBeysIVBawvL2hNBPs
OZsRkCaGD1h54trTWeUcJxVtz2E1D0NljpyamRwCQm+I+ovka+kV4xbwjHwfMDfz
cSZtL2M1LSt0sl/Aax+m23zSa4x9MhoqI60RiKe80YEqNxxAm/6iT1z0iuSFlA4y
VYm9VdQDibcOKd4NKx9j/m9v9TYWXG59E4+w7lPy58Kl2Qeu0ep0Gpyq8HIJypgc
45IFsSVImgmEVeHZAGQMmPwRHnRF+xyeHo/+QFbvZ647YIEhX+/omz24QSFO9VDf
d6eAk3gXW/7/zgb/u7+l9GFYS+Yvw/A0j03198oqwDtpILrMrd9ee9eoZLrpr0kh
QSWBL1AY8YdumH/ZRMwzmSm4T1tsyxbL9Hbs8FMgOCY6MBmU8nz3uk7DiR9w27RF
UFkr2Mrfmt93vaeeo6XLK7KOspS3cQ6bpmfsBxMnZWRrGvmpsB6KR3kv4m/H20ui
2ZUNM9wpFpouaQbE0/oX3e7f5K91i3t/AoElivQMklK61riZxgvWtt2Wl6VMErUI
AW4lL8KuVcoMaqLIxA6qbWoqO9RgHcBDCTCgQXWE2S9UHTtW85c6wUIbm0kVsU8J
gQpnh5ABzqQCfTasfCbYD2Omz3utaTHLEGOwTi9QadcQT9LPFqbp2W//Cja6PNEJ
B8QmZcidQz1wwNcvi5epkXLNQAoa6WybEO9ThWF7+l/7FK8FZiQo5Tupv6AkWxbQ
TkWZpuvdh+VqU+lQcjN4Gtf7si1oQQwdQ5O48Zru3HK/SnibrWRB0OKsrM8EbpMO
aJ0qqpiG9l0q0R1XTf1FPvdV3c5xmDiPyt7i6thO/0s4jDGGuyiuq3cRP3HgZcYZ
ph7WGoQXFazBjhT1LVbe4w8GaHisJimrKvZ3LtcYc7RzsdKwfYR0+MqPw8JyQgoW
Evz05OoBEL7GLqybRvkXEcfFvlPH2y9eX1y1b2LMOMeEMWLBauIGt5uS6M7NrLLP
ecjcNC02Nu0pfg5tCyt/p1028/eQOE7WBGj8Yk1/mBDGSgDcGYdBeInTDanL24wy
99CP9HsNAsWllRSLfXbmBK6WPbVFnHHUeJkFxchStJNLL2C5t6/xnlc3DhJpMLyw
2TY4i5pKh6LkoSRD0HgATVQUhY83D88w61Ez2sdrTm6XXQUDm9127aNJZqg3zdDE
lraeK1/cC90oPj8HjrcD2qiu5R3vNSHa9fdeJVWjJOSNw4BOIkHbiIWoZDbrf6jT
gArGRj2r1jxUlRcYYwxSQAosSvdyWktKEuouX2rFLgMDMOD7onwj5EI/BdfPI7Lv
/epiRCXB4wl7n/+OPYjvZRY23HrKBH7Zwn1dIuu0qKsmz8HFyKR4QI+l8llJGFWK
1h+e9B3Vs1ViEB5UkrUPYLhPSARtPvZeu/tRYmWFlwY49vR5ZRG9ZnoWYOODfPdQ
X4x9SlrHGhKXeaaiwh0qSCFqmX3r7qX7Ap1QbrgZOy8xto71QE4Uk/pXMPiF3RH3
Q/WNOUtQz50UfeKekjSpb2VJ2MsE4kpJKSO7UgwaHfN8pllD4KkEtj+QRq4ndato
Q1Jja/0F8GcqH2WExKrAYmtwU5NHO10MuASKZiS1t/RjxiB6d7ebL/ZRrpHqciN4
UFJk3kHIfBGlvm3/2VloN4TS6BdtGDn3F3+b1hpBTpGS9QiF4lmUPuWwns/oK8zp
WqvM8v1AegkvaEgfd7gGi6gUPq9YW61Hg7mMaPrR+/KZ1n9aTpJsVdDKg+mwkVoP
xFrWc9biOMbomB9BONMZK6qdw3XVDGHgqvElHPC8y3dxNKMY90Wcfkc8GacuFPf6
42N7ahi0vCYzJj/cf8s8TAMGMthbf4nrvnNO5Hu3DfppyggoOEERrh167MCe6D+a
+MD2kgR8H/nJhTYGCuurIO0M9cuZf+ATzgg+eIMWQghMzopRSkiKAnsJ6nWhZUCg
DTsXphi1MEW6287C3vCAc/QnMDSxrbDSd/une4HmYgM943Peh58yQlg2ucjBZUZT
bVjiHSLI5ZnjwYxDPUraDdBMtNCI8gBGHgQPkdyS0FYp2Bxxf+kiEDebqDdTLmf5
NZVdWZCGDhRoSv7TXbn0rxf8Jv7nTCIr2LwSEt+bf6IScfxhIuFr/2C6AsjpTMpG
PoBd22lIGpL7PdmW4SrKSUVBAYROWKPAU0HOYU+G6lD6+9Vc1Fsp6EMkA2774MeU
M4H0jSGmYqkTd6eyzeMDXPKCYp+AObJT0iRxL9ikdxDwvPz6H1nQAUib+TlfowrC
2OtM6FrEmHxm7HQreHVl8Ww84N2HB+axnEekpWUBTBb5LECs4iSpFwzSFy9QBBSw
rw12C4Z4CyAXHovZlDvXZVsuInI6MQGuUQHfLMastVoJA6yXhyi2GPQ/Q28SVdHa
luqT/3FMWuied+TLT3FyP3BQzv8bJmMjp7DVjImXCbHi4OfIs9WkEYzghnSvGjGj
sLv0APHYQHeEOllSxnvNDyanFEPrz25FkaP2IqZ6JrTv42LK23sMQ7Zwznzvw2zJ
Es5HLc/FmaW1pweii4mI3i0vVEsBm6B5Xw87Pq+Y35m0cVfftcpYaYXNDQM0mAcU
NMY5fTUAnoO2X+BRyZeV0gzGeNHHOoakM4JftDrlIJOChQ29Hq/IYbImRxupoFaD
IcBNvokkBOuK47f52jngK2ldDoKYNSvkT7K3P+Pv/PKzpzse6ghKzklnruAL/688
nmmsmdiBhs7zywb/M0l8tHZ4kHcaIQRxEBIs6y9+1rA1zVGAJvuXzMt5fP49WPes
vzcCRDfkG6p9pnyPwl92PCG/0J/PyV06z6uBZMEeCuzTO1lTI88JQKeSe12IUg+C
D2O5cA4SQXFgwsQizGgPjWcZMUAkcaggg8ZRHkcZpH/FA6F4/BBfEDJhaO47yIZr
1k0fg0l5OcQB3VqpewswAruh2T53O/t38atfIKQFkMcLg2gE/aBu//mqYw2jy3qO
rGxycSRS/goIjz129Sgv3gGyB5bwxl2cv/TEfDJVcOgPIdEOYjzujqUinlFHrM1i
TVi48zrsc+gKC0p/vEfI0Fr0+KVTFnb7wyGiE0ITI3yRDPt7Vuh1/9wjN2dkwc5a
/niNZjQHyL/CJn1crJIF3GSkzByzLAw5NnTHLbi28Otwzd868+qHADXjB0ctbJpa
i/Eg9zjeaFE5/57XNeUWO6gJ6Ldf+ZMM1rsqOTlVKs0VYpFhtuxNl/JIacDbCZ90
gCzZDMdxJIcp53GDDJ4OH8+9NaboV52pJdFagEW2NDbWuzUv4lAK6tUmzGLZlVq6
I/HSm3nxemKIqdlWU71KPAShSUrBpDB35TXLxdo+kCB5o9joAVLpcMurMdtDqQTp
HsPXsMiQOA1bg7QQ8Bku+c120A4f4hiMISPDSmoQ77R9dbs+zG7R7c8kxY2u6/pn
MA/nu9l6ypEkZwe+w2LwVxaVGWB6DmO6N+mXgp3xmnFhOz7f0KT5smrypd/Uqu3G
k1WFZPmubdFON0EoRWlnnI/vb6tInOd3glheGLTZMe2/a7qu6C9S5R0Sx6Zj/g+Y
cAGbRtoWFcgIT7RUORAmR0wuptwTa9+6Y+3gpOKJgUeq3xkpPNBh2ZWKCPiw21Xo
Fk2Ba8R8wM1ly3w3EERP3X2JowPMfUrRc7ooLf+gSLCE7BDEaAIohpvCMCtTbhot
HmJpPHei0KnuUNfwJ9J307FAoBVnxVEMIdsWULPeEvSfTcbMDFhiCMdtEOyiDq3K
aXCnKnJsgPGVxn19V6P+PiiknpjxVLA+dcemd92Wl3lJYcY0rLmCddm4HFr66/nU
YIZtknlJwOWbMJOApvWJ89h01dnBoNiRPmbNLBoazyK6RJc/rnVQa4Y3v9iqDM1O
SYj5ejp2bfzwNFWXbH1O090gqOSJ0gawggLWdawZ6YK8lSIk83vBaKSmxKYiLsB9
bVDRkMLTcqBRc5b6UbmXHp1+oMg3BulJ+ZqsK+ljO0cxdsNHRYxd4Y849OVl7ya1
XmdaXNSVZ5IYt2Oh1++rXObZwvvQMUjNmr4DVNy9ZZ7DVHXDA8qUn5r98Z/GMCc8
oN5RLlRaNXjIAahdeo0LutBgpW+/+D3ER0GPOzsA1zvANf7eD5BHucnh2gNz/gmd
kflBZBaHdKEKl/pPbXZ7Wfi55mPajFAi0NEr8Fe6Cx9BvcZNNARZpy2qOn3yE2ux
1Vq9Hc0PQGOAaJri6NcxJNkIF0Tp3Q28H2sMc1MMVTpl8AUppMXnbnBIDcdncAXG
hYTp0kBGxlohl2alqBoShLuPM7UdQDcVpRraMDCzuhCFdtUN5G6zXl/bGaUPBxgN
YPLKAmSfPbJi0G15DhI9c4b3I4B/wbP36pUgnsnoJL1+9HUtB/kfDBT05P2Twze2
kvdVWoAoWlRoHmUO06wb/sLl1iEEmbhg2VLKiC3qpSaGfvBasrK4So5GJK09F9HQ
di1aZwmdGPBVB+CvabR2n99zpu1hiR+95Kyd88wZUgoefse0tVWKQTKeIzl0KD/c
RmElXme8iz3sOCURKp+lC1+F4zfxOU76mvAP/itUytZa6BQvfdY0K64J+1Phy5db
lMjF1vjttb/kxiaNgy6Fx7M6A7sJT/6HYGsOEorfm52BYg1xqGDK4pEbjC12g9vS
c99Ysazysoi9p0tkzS87F9Xku7DlxJ1cCEdOp05vwq4RGZY5u3GANnggoZ5rh9FR
kumXNViDw6LJlLV5/xaWGqNnOFaAHgw1WtmSB3KLrr/JuGwAjGSv9JAe6J2rXhGd
KkV0hV05MTSlUUT+hezwi3gKbBhQ2rogrRk1QoYlgq0qGBMRp4qyPASDzTo9yTw/
R2YEFGHOI0HTRP8J64vcp7WjQhioR0gJ0ul2OE0qF2txRn3y+103kJRCAoWmP/FM
qzei3vs59WovtGPUvzF3ABNfVbqOsNMNGcNoU0oxlhzzBCpQxC0cUK1C66V+IVhK
qhc0Plq2S+9zZuv2CDVLCjkQmC4inL8lw8nyXOiViW5JN4qGXMgXadnagN0bQ+u7
9y5sFnrzNl6hV+pp5YQdDsGqJNT7/QKSzbHcOaE+SM9Kn3B3xI8yt7cA+ys2BwyJ
gvuUD6N4+TKfWRnYwzzNCA+RXys+PDmCUxSe0Yo+bVOBPG1nofXxgpMAvA4dz/Yi
mF/uvH6u51Xv1GmPUEcZEybf26Vl29YcQ6o9U92xNeMTTpj3k3jJ5TxYFQJ6UNhL
gDnZTm2QFytxBpmgzp0eTeaznvX/uP1C5miIXk9b/9YpZ03o6Ma/6Gi56iFnOWZL
mZeSeZOaxurJi/8hKFAzf5SD8EF2k2jx9OqIj2Cavi91w6ZuQFTIu+9ktUgfez1V
Xv8shqxZM5ZoYWREUyS5dnSlJzxZqmntQaIQziy5ONQ/b7G5xnLsOwsRYocLCowC
KLWtW2/FzmmlBUHo9JxSw8Oq62uZu2O8AIwDFL5gZ7jBH4x9s4PEywkKKb27wWpM
MIMzcVEpGz0nZcvU8zGr3hOwlTLwLch4Sj8pZGvu8n6nU4nKGPpm3aSIsVVrXXOk
6Y2EcFX/1w4UwSZZALCCcGi7fJzf/Sh9ooHnJMAi/mDfLZZ1r1dowtUgQ4U3CRCh
QkTR0AZSPJ8E2yFgkv594MhPrdmwcxDmBnm1GqFGBT0oTSBeN5YcHF0w9GujyFiO
eXZ5rb3iL5x1az59jteOCMxVHv6qBjdsUE/SOLBQLWrw3VEYhc7g0vZPVdXQ9NVd
DxytKW+hNZVGzBbKK1U6dQvKh6Wch49h0ajbtNgtSOwrA1jQrnJkKeBEdNwbubAV
0Gh1pdtBbuAmnU5+IBuGAvgxi7lo3aotszIcQzy5OjQqLs21hdSCobJo8Wd0mz45
MRKQqXqLwWKxrLv6IbpkzRy5i/Get7VSLplQfPSnEN2UriW/dAjLjqMl1nS0pAZD
AwVN2aTRQAf2SfURfhJj4p3YNO0kPoJ0DQUK1BI8qguqC86MKB9GiAqQvTKoQ1jR
Ys1VDF5Pk9h7SSzQQAlGmp2urrJOMKiPbFXUOeJT0AMdf+yKWE94QvzjQH4HPjUu
N2w5ijzfMH1SEoOFpq3hMbidHBo3YN4zmY1Fb4d2+BjbuSS57JhtBJWYma4x48aS
MtNapaG8svdR1gP9+Sljs1Agcxpt567JUOmxQyQ6fIC/h2dFrNdb8xOI7zUl2Fsk
OCSMENp/ud0LchfsX0b9L83v8AT/lhjQe1ijBw30Y/5N9aUPO+g/2T6HMzJ4NQcR
9Ff1mUT9A6n6DpXyHEJ2OBwfRxZq+O6jpTcwLFhVywBG3zW0u+FzB3U9Ryj6knqd
FRiiqI+wu+R6pMWdJGhUBzjUf7BLip4LX0ZEfJSI/UC/CAZuJSTbKI/VWtyJ2EZP
NbIWpO8t57QRHNi2J7e/Vil+CiXUDEf+DbBx2ZShKfhS9iRI5KxYLbN9C31lL5n9
ThcVTha34HPxpiffRDSW9osF6/qSHTxL/rB0z9uAM/i8C18GiB1/ESStQ1eoYEbr
ucTkrVIqtmhMcyOT2pKxzyYJvFYkdIeXOBhORTgJR8NDarxAh8miPy3d0L9Gchc7
Ya05Tk/ZQSAKFIvflHXG/ALViYGLMmW9mWvir9N7A+htKXpuZHUBaEDS9Lv/f0nH
8ap8QrRHPGZD4X2ENqjVX/3L0Lx+cFc7gg3ua9UN0ZXpIArdGbU6udXegSSgBxWF
GMlhiOMie3TMdZtDtF1u3Hmvhgb06TeE18YALgc7xKVNsHIv6AnrSmKCL8uDUC+R
t2p+dnuV9cz6lCb5mLJrh3uC+Wf3xbqkUhjmmb59+IP3w90X8c5tRoWv9XRFS1Ji
Q4CcvuqKsFIh28rrd9kEkNm/1hiPZ+wuLrOk6xoQgye1IgC8XCeS84RALHf/3zB7
qOs3MFgOpvVRypFtm2a08P9/DbOFdH8IyS63/nFiTP8gg3Riw+gHPrU9GSUPQ+97
+bwgtSp1goPiV8IGprt9gHESMphapxm5fxqOXkIQqeiWuxPvFbuTXfiC7b7a65EA
MeKiSmf2KtRCrLaPpgvHhSEmW2l2k9A3X473Lw4Hv5Tt6KvFTwzuqA7Mx8OceHaw
9EYRpaZtzQGG+YKJheIXJ1Nz8iNrur0dmTSjP6zqjTKcg0SFkB9GJ/4euFTz7Vi6
OblSwsBk+PIhGM/kuBvJOB+L/CzVnPuOlDCTbSLh0WFBodPX2Xl1r0MNo1Byd5sI
j1Pw4vOuqCudsMjWCKtr1CaGAJR+ccotSTEVqFNFsGiiPMJkmWFNlnv0xGqVwLcP
L01pYYEZ3ZvTgOtLxCDbLJ6Mostq0grRuxKUtcG2cH9BvrHqZCxFHWb0lyrNvmgq
WUBc0nE42T/DwqVToLzOJhd1rsiTU2AZuLNjWayNezzasWQsTfRdo3C2mTBYZ+QZ
DkA2d70pLdKG1v+Ovrx6J3kQ196IrXXl9/GEzzzDmyP0OWym5fnYxv2LOQdqJysT
mqwCZMpsL6Vtp7dvS4J/qfubvRB7i9G+t7SPAJURxk3QPlJOnCRtLzkunAFKz7cU
Oa/33aidMwUBnHYUxPLRoKDM5t5jSK5K+J0hs/6mIHlhBsfB1jeioI81DqpFi4sF
0ebWheVg/SPkI4hk110QFkdW2+VPAwcvolBb6SQeEMT1s6jgXu0NDrSsC+XsJgdI
1HRFiIIVcggvntoJfx7WjF8ABPReIdXYFZzaSUiQaEORdwq5VksziSUK5AY3tW3n
2CshihA4693oMVeMRUY6m9tZaASIPpSFafJGlzWQnfvmF0oJsRS5ZdkVXZswCjg4
hZfA+SIJ2Ce9U2ue8sPh2A62l61u6efdXUI3ljLOva8+LwO/l/gcJtt0nHd/TQpH
mDov37k8LtFKe0jKXdUGJEnp6dxSLC0ynOi9EE2Iap+MPjoIFrsLzJhF7dyHhToC
Y56BEVmY2Z6KbV5PAFkSe8+0ocsqUW+FFMq6P88xi/5wI22B3UbY9FC2xmJ4aiQx
NfedzFRhaTSFSRdGR2QsUDpCA+A3rpRw68xb6dnNuTZyHXolr8bi9ijJNnSWPhr5
+dVdLJBtul5acowLAPs6RxNo+ivuIxOWEWL/1bjH6Cs3RhZgHs7qSZg9LVkosetD
mH2uBhfsW4jnRk7bMwQ/Vosm+u6Fmn7iSM8oE7fI3JdPw0ZOP6bfP6p/Mav9nIIj
FcKqwTf65qTTlVQLsCy7fAtnHPcXTHQR2cMugXMODWvuedQf0Ent3XL/jg88f63G
HzXmQIFiGZLG8nJl3cPBtjl0S3DkFSKupGvafG42whMMGnaj0QWZ8BBk1Lt+Y9mt
+R0z471in4aakOxH/epQLiND4O9RIq2IppwibiyF/5wExvxyUy4yeVbzuwYrZ9HR
rGGZN4mBVz7Nvv+PN5O/5qijls20DJdcgiJ55bzJmpJ6RFdE9vzk2a8HtOn+ODEU
Ar2hDnVPkUeJaj/vgMPzH9CUUb+WrIz+f2PgOttXEMOx7aiPR27090KJ4l0SAcsz
c2U2urLOXKhVL+wEejsr4N1jZJ2Il6fii/ZnucppP2FenFD+OgNjrjyrFXSSVmeX
f3NDsTMyxE+exa66gsmvvwJURLNWKFxsKUM6dWPOF39vZROvUmMwBc8s0jiRC1+E
TUAxzlrOuoK3xF3i9G2Lrju03VbDwzzS+Wc137JWjgg+9MqwR4L41LEqbawQ9nOI
z+j+XTYR0KnIK8xvcxLmI7BLLSnr3l3Q5JZp0CgSmfXlEhGH2GOE+px6ypCaakum
aVcT03LARRzfO+/1RYfEArlotJE7C9TrANaugjVt1TVdLJ2E/dJ9OoBwZ/cM4clu
GAvj9z2c95LzORR1PoLz91WNczqnnT5PrT2eHPDZ7KHqAcwOo6eKFzCLDBpfipmZ
UhGZPF52NR5DqAoc9P1sd5NJK4Vk90VVnG31IrCSAcl+aqtYa8Ryws4cXT3FqCq+
mIrxS63Vv5iYzuPbNodrvQJHmp+x25OjAAp/jhX8ALC/uMmejPAoK/Sf9JrC9Dvb
rKboTPZ6EhguUxY5otuWrlGvn6r/VwTQC0AO5PHRa0TkDII9ymKohe+0eyq8MZWu
eKoXzElZ11Ra2snUx+hRfwsM+uYTQOwtVL4QRVgWeLR7efNSIAhPAMMnyJ3OXE9c
Ej8eGowWuLkIXVJwhDyguaSz2+7sufvcONCQlooBqjwHKAkmTZLbWpJu5ngFDg5K
c7REPdzL8kVlrVjVUxbmolbW7SH1xqvsVjBjrjp/PbFF6ENCN9nco9kyyDBeKGfX
i812p6mPq4F3KCdVMRapqVMy8kCN4vNrYscDHEp6PY1G5NTsu+btF4617vETSyoH
RbJ22XQ+MKZ022uTPuu2ezr+O1zVsMJwbZ0Rcg3fqJYqxzqTMbiOBINY3xVT/CNj
OImKKltvSdaPJOd9i5Tx2GMv3oJ52MxDSjCyZxaxJfinAGMdhUcjcXePn7uP/7FW
IrlZtsTOZnqRyZqO+2ikmPQrpgubZhxmIgBdClrGgd/b2AXg4DPglqmHG4bSTBQW
J5jBNSVaDeMSyg/Vllmq4+eSgPiebdKlTJLzFMALY88PQJEz3c73oDI/vC0yb438
LB5/pFsDKuIiUUo+5l6UJYC5pva6e1XuLnrDAUMA2q6SPTVd5OPAzTOQTtHLziWr
1jfYbAuN6vKdJDo9dq9HmqGebmtyiabBAEPmT/LBSxBP84Z+yHLDV6YHlYV4WJbg
nbWGlcpE2Q8TjGZqmr533ySj+weqJFL1TYApL5VAc0wQqB1NQOruA1MFDtUPD1Wf
KUbXy7SBQSRA8fXmFhyaU0H8drGBGjygCrKg7ZNBm6c1nD9dsAB2QzJA1DDK4Jgm
HeVbTo66ilpZBbnUG2AiRS1V4v22SuhdSxjCfkt558OiOriBCtUHkteAQRVy9D6m
+7ZFH5Xtysmj8YCRUJJLbxwTT3ss52yw5pDJGKtcaIE2VEwrcRvHgapKOKDZvFvX
9LwXiXMcKlZ0bgWqpi/OLV36ZbjagYpy2UbnQUPUijLY5oiPfgyMesVJ6MzesrLe
Xdcz8Hx3QmxOHNllTmU6RV6cDGEAkzhkYYhJDNSeE+DTPBCF66zG0iVM8jgrx+3E
/7jCiYDC87Mt9Gr/T6MGExHJPmzPGFHbgjI8djQVgqDhmMXLWukT5jXXI2UFOHTK
Goirvapv/8x9EwckrfIF2ULmnKgLscaRvEsY3GAiG42gxgRRtLFMHxUdyoaPY3Nn
8k2J33MJPkj/3nY+dSvmYMmuOmJn8YzO+HuST9kdQX95ubxOvfAqL4os5J2grCMH
JsPsHYIYCR3YX+QIXAaigVZHUU7C4C9QV1ZHMAWYL2NcgWSrmQKeZrYT+ugd0J/P
Cxrqy+OHNqo4QWjtindRLHKFXeiT+MIQvF4KD/16xb8523GQ4ttmmq7aO837IGFs
5dGFbbeDETWQs+v+YwBoG8KJLxKYvZcoD6boNluJzyVOhv7dqFb0VxQW0OXWRgmC
7mOHyoF14KP2XutQ1HwyFdEoed9p9pfzez8Yb6eATci/+kNkPGj51nX13BP+286L
gauDbrTG0IuSIk6zi85INmHOFZ1lysBlqiRCgKTlGxSixNDFWbobDeDBP/znVWjs
7LRsvQ3tyXnjXsju3B0qHBSsYKTxO06GUkE8cvBGWO0F/sNA36dMDlkofFwzRChz
GO0y1jUjpv4T3JFttyYYtdyu+HPSCG+RR9WINr86tHUze39gB38au7efDLMJtHQq
oJq7byEeRI9tD2nZzpZrxG3JH6OITduGfILJSKaNxjvFXmiS+TlPtsCHjdxf6qhP
qJ2E21TCp0zeLJX1k7Q0kFQIiEQUaKS6uwqGnx8JX3y++JKhcS9VJvk+iojIBfoK
Jwe2CvaKT/X0SnsbMRgslSqm7bVP73evReijsmjxnDp5BRvNjx+TFO75NPbKunzX
6QQpQs5xiCQD3+WsptXQHkETG8liYn7djRAPgoZndFWiSbxfWltS+ha66jb01iW0
BdR+ZZ3tTWXmix0gqkE1o3MS+N/q48mftKDwZldh3ZDdmO4QfT/vpuTHSQSD4DjM
sNJ4Sr2VkbpAL23moAYlPsCZzMOnPIYURKB5oss+lznqz1tDkpcx0Selr045zUNN
5M4KNSKkmYlm0+0ViWViiMlOLCXZTG7rt2LoYO74Xr9qsnuYxaug0FMiCLazxzyi
J/X3BxpJ6tp1OSxsesG3yYiwX5s5wyCV8L5PKwTiJL1hC71ySUDLm3ASmJBWFkZt
EPlpENcHA4zLjSsmDKeq18WnbFM5pLQznz9L8XoXGDmLR9iKPgr5KkwxO1EmikU0
vCzymjIQaumZjF9syQa8cJreiG7pvziVm7iLr60B9Zbvm1XjoB4cZjFcWi8pBjU2
gSOV8c6gu8pHY8NKmkh28luZI18TVOiFzFdRLuN0JXkYhayIc1j4qsMYSq58jFr6
XtGK/PuKVBZvYEtajiBACTT1osVKWBTbmai2qnTJi1yqanzdOELjVmEgwKV9oPur
+jk1RsDlvEmHfaY6rOp6mWiGWcKXKfW0pYUnT+paATh68RayYrbMAsbjHE3rxvok
YKHx8Ipc1xkZd1WL/4IYJzBILLmatMDgH0CO2JBN8oMSRwwZRGQF3RxJ5AKWKeAA
ov+it+j7iQCc5hHeBUQL7tzXNzIou2u1efLhIA5yIqE8oN3BhwZzpf9AtNEEwMtL
gs7hr6RrNnvuXdo1QIu780/Xz9+JwEqbdI3EdZlkWsGyTdCL5+P2vR2ruJngb7U8
ksDhUxwEFUxfi2yAuaO3xaLoGuu+0p5Vc5J2lbFCzWJv91lIF7pu/XZP5yhFugkB
cS1pnI3Mkgv4E1fWl8eB2Xa8DlE8/32MjVUnEoCjD4nOE4HgOdHQ7r7cKNWUY10Q
HKQzpy0Ap1eKTpfgGAn4NczHqygfwD4PN3iSEIAsCX0UuFyKaaWmjD44VGZZn2s9
ZN08a8Sj+oyzAikUbrjtaw4qNgg19tm/U/uM3sGQaaeJuSVNvH5APHH41mB5OxkZ
MAzbAm/mmqjH/v/cjIvvsOtBzNKGlkI1qILRCmkCjzhLAAxhbGyRsc9Vz/gaDpUo
q5lPjmwl4YZhGPq9nUpUXAndJw0qA+HdyR1hrvCO/YqSEGvQtGZHjfHTgeOv8thG
qocmpodybHyWf4J3fmgjJJyAZhBis+aMJ5TcOghnZAVkJYmStwKpkmI1zGvThYdX
GI2h6bP/PMY4TGG4pnE04aXNoWXJ5h6aGJuYXgxdnOGWS39dJjU7DH1O9MiTtLi6
2Gby5D/wYeAiMuVSMNvzbN6YB99Yt7qtYuv07QgL7I6S4ym78uDSqi8ve7lcx0A0
YxHfOJPH5s8T+P07UEASvMkqVu2cWaIHWzCiNqhp3EsPcqv2vGKZFN7TFaOmawUx
ScfsBy7kOVG3lEtRocGSpsEYW3gCq+m1uStWKDxr37ZuGb0+GyLFNU+HM378g0GS
tjAhkOiJJVgizwzQ0zrvA8OmliSnQtQMcrdPNV6F2eWvEUEushE/ufilJAjDBmoI
XnBayBtpUM2huCzx4KQhsERurDMNhh/zfKnam/TrO3eZT8yCfwsIpMFoMpxLCrLH
J3+tfC84jAOEyFUSq1y++jK29n8kCtITFQYFTiHsRgno5vr8HrP7TjDLi+cFvHmk
8KzAcc5TYWXyTJWfW9QRuvhkMY4/IttS5bNXgTQBoV6tq02Nk9jm1Z9C9kro4MDz
vvHh3rXt7U3mT/iX5lOSbReAbsljLs1MfPYcIRoJ2uTOrzKJ/N9OP5Me+BNK7Tyl
s+WpoE8AjhO19rGxRizP6DRE8PT8MAYYXpIpe0AZwOlWfKHVuzv0LDDBWFNlHL/i
0D8zZOtDTeIOfrwBkH+vg/J/V1DTOMaBDiRlxXo6LTrceZhYrnNSF/u/iWifg2F3
riT1xOhiMiJ9LkWIuFzezN3h32a75Bq8Mtvb41ECpl2MpQpOi9vtBd0j2S2T7T6G
wZVykr38IktC3w4lWre2JhFRIxc0FeTlf/j7FHV6a5jmFsLXNz3NbcQkOka98PXm
enAsz+m4+LXnVb4HsiBMipjATt7X+XsPCBKcr/WlmoNv8z0an9Qjk49WlV0BRAww
hwMj4HtUvZdOEoZ/7rmBNNnuoMN9W3160K1lH1f/wpuovdrfthFdMGSJXjJST5wE
dBzYCGtqAuWv9UOxyi5XTTzjYWLGnrnunNS2N9QKTPCcW+XG5EpQFa0jLULfcn1V
M4DerIlMjGNf5T9P95h1fFMHV1LHux7diukuI0MteKQf4Iiq6Yc7pYXv/jRtYAmy
5BXU2tu648pIm57kA5ZLi2CBtinJdK9KacicUrcqsBt/LD+h9co34aH+2HGGFfiZ
CgV8zfncaRnVmOEIQuRF/C/cBMUXbWniumPyKMOTQU8LytHinOsGYK4OJPN4THPh
Ph/rfEb7gnQWKJsJItwhQb8rUl/LnnlpyMH56E131pNcbRNhMWYiCzlw4/RIcHpI
e6Mc1HjeNTra5wyhXEFItKzNZMzEQ37jDrsUlGHpNVp72DmEGGUO9Ht/yldr11wn
Ul99btwvOCeIEHRSFvlmfQivFxXINmopx/rCyAg/VmFck/qf2xmV+dSmS95EhWSK
/e2469uDwWWOHUqMKxGdyNWiiv5zneP86Iz7SK8bEn+Mg7j8bmr+3brQiMSmyTHb
TyHfaiwD0jqxhBFLwd2nw3ptDflhXw7yKkQHNSNtWe05aOULY5ZV327HUZFM4gO6
+YpXg33Jq72+5k/r1D3L8Wb3RVi+QuTkcpMtJB623F9V/JRYKFl412tJomQrmPS9
IMw7oD3LsN2r0lIYF4p7NGh9Cl0RXsvWzTS0DDKX3n83sPzgdoR56m7S8Tj//Mp9
oVglK9hsFastK4nm0kXEH8wJ9gURaD4h5uIgAbqgYZuQTeTWiVrO/nIToyzoHv7n
OcAK6BWfJkYb7nGwKxtGfn27mxX7boG8fqJFCIVnNCgYdaix/l5B4Se/pHuQBTlN
4VWqNtr15tCw9hH0stypxwLxY5tqVUW6UQWdq9n0fv+b2GJhv+a7fOK6MyZSpuuD
ippJMQzdTQUTndapUwEDUORINOpscHZ9SOY7qB0Vpd34osR19l/oSb/jry3plSx3
GxJ+vophiAnVFk4sCIu7NO0aP4EDMp6qPO3tHFuz2R8pUMTVFmHJ1lONB1B3i5RB
iExEa5VwjmZTOhvnMIZWn5fboQygNY7SfcE/HoWEWJRGT3b3bCqHMcBoBI1zeEuk
i9qDpefPZBuFS6sYEqYyDHh3NJcFs3hEZsve7eMzBdLcQ50pkNwG90uqm3pbitz3
4CgRPmKZ46O+QwmLX7KC4y1cUtpMpVPbTsSVHxv7EDWwVZ625eXu95iRw9DL78DS
uQn1BhRZVBzF1pEiuBCm9L8zHzDygb4gc6dy0OhkLC5KMfkJ6WRtDde3tHRntsvE
2jPE02iI2cDC9Q1XP5fyaCzN+4dJBr73vWFAD6p5bz68dG68Kc7y+JVqx4cTH6GV
RKPFPOk4L2B7EyL9XbqkhPIb2cQtaLqdqsaqBOVyshZIbkUE6EgzjmJmuDi8cgUe
nFxRi0Hoba9rZZBtqCx7/VK8XQE2aYmBiCFaybAB81HFZsnFZbOlsfMAlKB0XGTH
I8ICSoqily2LJFEZ8yFX1BdPV5Aypb8ujHSwbh0DgSuCubIeQLGucP82+Mu0JBzM
3y59akRIP1Z7ZlnPCJjUYqCyocpkkz2yv5iv9k3VqPec1I2/ey7EHmhL253quBJE
9eKNvcwUwqE6NppNAgpGYAfoo3wsHuZTFn42T8F0uJrBsrQRTcu0aJvXCvAqP751
ArsN8L/uP0j+u97z641sta7Hpy6YZya0k9/fsZU5dyqHGbhOzczVGxzwB18wvXgz
RVfczCh0RsXF7chgVgl5TYANK74iomqdJD5vtr4qy6lO1UZ00AHgzIbqClnAcTo1
FVHt53z5WeV5ZjRf8TeKLVdiW4OTf9SKpBvk9loaYfXrV+bLq2VwolRR5kk47GKa
Rf8xZqx+9kOqgJvS7ojsYkdEy5u+cNFzowPTDWP5Q1YejyP8LhRXfuPvTKVowQ68
kdoTpWo6n9VEpaiX+cf0+2/43eRItn0XUBQ+PRS/2qbR515Xxg92k05LW0C5XWDC
gYL+lQm8/3Wary4itPtB64wW46XNeYbcHSo0EdgGWOnqsmoDMPDcwC4kbknN2qYX
Lcp4rW3+7BjJaTUDojFWRYfz8H5Es+13tnuYMUNCaB0XOcrRbS/1G0ARfZn7FGuZ
TNXHRUMwTPNid4Fq4R4h+bo9qLHid0QmhmuMBQ/Zc7tibJnsiVyR46HKWtvdmW5Z
/LjLnq5gA4maDPrg01Fb78aEOjuXWTUHbco4mZKnigdUJxQSo3aSArh0kpFkR6MY
U9lRzoWiFTZA/qwNbm/HjpVbKxNpBef6p5CknWbLmIZV0YKEEJQ8D7SC9iFdzMQx
NjWgB9lWRQ/rId0AP9Tenx8WTgD/GyBk3dGutejE54sxdh8p06IFHuU0UQgmKTfx
GKsB4AdHUIyrLmdC4hQOHgnYci50kcirbc81Z4L4fbK5bGi2gFOoXe4QCAuYnKg6
EOuMvTaHH38omSmnGMOUUzB4vFaD5WCdJ+6mB4RVCyUj3H9tUcP68t0OMqxuShQa
hpRP+hQavfiqWHtdFuO8wk1Dp6m7QsKFsGHaVn7Ygopob1z1xdGsTwggJqZ4+/Wi
edtOyy8fFDvucQG4ZNpJ4xtvzZBuyRjiKLRzNkdRTZAfgQjinjlZrXjb0T7M3oY0
m71RIz3nI48quxfiW+5sAIHfSA7UxAseASUHKp3J5NPhEDBxU9moCYAXwFU/YP9i
2gv7w7hb+qiMRjLP1EiRjl2eiKmRaH3PxryrQ6346SwAJOt+hFHw8pKA/yumFlZw
xS7sLYSUbu1UttrHOWSJmcFAdlRoxuxsMnJt4u+3rsZjijT567cdtOXa/+5Cl7g7
HECcVhd+35w9RFmN7Hw/ToeCVzgTQ41vyhGqP+aBgMxzTMj2tcmkZrd+WTlC2DxZ
26Y0T/ndhMUa9/X2fg+EnspK0uZ433GFyTRl0DlnUB652IxfcgvTtNGqQcmAQJ70
pKUGo0uG3SZGd4zeXkF4Og1Ppvna786ActmcZRO/vIlVU50lv0B/vZGlFlSsgM15
xvmx3Nuk8i5wCafd78YC27Z2H7r3517TdlJXqGPF+dgixFCEvOzXsfkVhCOn7vYq
nHA1a5jDNCTB0YFKnsZ3b9HC34TmbErYF+gMmhQt05qT/xYUu6AzK5rHbcdx7fJQ
PKorFfER1oU7ZwVkvYagxYfSBG7UX9ebjynfkUIIwkmEUcp/UySxg1/NKWyJdy5L
9XfI+5Lmx1PrfufezP1qhehaP944HHvgSo4cuEi1XVjmRj1B+sS/CCX8rBkwn9jA
KyQjEpxWVloserzOlE1Kzyg/ODnDizkhyBgrhBbUYqeRr6R/TZOQHNCvji5UPKOe
MZXoOcTuVpzuvmWi0X4xB2U/w4dFm+OEiM+he1OzDq4oA0IzZyHq4hb5di2Q5Udx
sAqb6zJgJEqC/FGsusiGAN8g8Qjfn2FpuRxUAZj+0+sH7oAKLeXA5eKRAptO0SYh
ZnzPsxfvcpnCRvU6D7e66+djc9Tc53kE/n1ytZV5GNFbQ2p0/Utz4O0tP8la+up+
hl4Ka+XPKJcf7qf2TmuIL0e06OYrGRLs4cpGh6JuWAhn09N6RPlSCQBRwTXkOG6T
g19lVw1EO5VglzZmb6e56w8NCs89+0bIx9g9vGkyAB5vY7d8VD65jb8Lr92ZUFgO
mGeL9pTofnfENpSiH8H3GKsppiJ/EgII1xHJJU2zYsxYOmgion5Tt0t3NxTSO6Nq
3ME6Ypfc6vUwgb7P74l4PkxqgEr9vUmtMnIJXkYU7QwUF4GvHjdPpin92GT0N5+N
xGQt2F7tRXQ+tC2dlZs4F0WNKoexiNna185N5gaHrBYRtE6H56uY/+ENN9ROKBZ2
uWchP/uztfyJ8zAU1xhiR3azeQCoU5r4QgJwNiqPuWMUPachXGQ2vweSwKCtAgVV
1kWZhh75tpSZXruQ8KP1hz/a4wDjrsvo0EntdDk2b4edYM1P7POoSqw3//joCHTs
a59rjMybSLzDVkX12mbtZVbozSQz+LkP6kCbEfOYnZq+hRjDLGsMbcVcURiex5xB
BWcplA8Gjvo7ukQfMnoNutn4Qp2rkOi8QnDEvlHfRH5CXjWAB8QxU834CkRmleT8
i/pYYVyykHxlou4uqL5agKfcfbntbEZ4o9Ey5z2HvJkrtbGkJRQuCeTskIDSpf9K
AslggH+w01UA1bIflQYaMrcZSNjpeexhHcX1DfV7AGmqe5tS7vVFJRaLa573VzLM
FhGYnEHPdTuzMwrfU/JItGSU8bS/6s/qvvdrIXgAzyGdMpKIOGuKI4gPIBv6i3Qe
5Ig5bzLQZHMGMbM2PmFVD3f54uIJnm8L3f8vGYBPZMcMR0oW525GQizN+YLNYNqv
3bToSqxVeTkRUNnk8azb+CJqnb1kMolFtMGPXIvLP55uuuzMXUFbGTeg6rxz9XSr
68/Ho0JVTTomin2Osy7YDlCOA1J3ev+63JeFrlbOikRqMwZdtvTI8nWcMiE/epua
y6kFxaeVRaPy5DrKRKMXemP+AuAwvMB0dO+QhKAK7QEwKdr5ysah0dNkErwunGF7
XfJ3B959IFDspiUdKxLFCrNbJipN45mp7LfurRbP/1RBBClAGFUDVAiRKzfs/yug
YKu5Q70M1O4AVF4FxtaPExUVyz6KijLOF3dO4lMEhIr72yLgKeXYdFU4Fmd8BDGY
fgVATLMW03moGeNWdwCMf2+1Uv7bltGgwreEmDWfOQ29oNHj5C3769T8RkfPU/gg
tToMKhlAudTZssjhR1OR1HAEypf0WD3/VHwmJHfVETnzAJ4Bumskfeqbj2Up0+aH
rYmgj/xcZRbitsfDSGP6jQw1zQyITJyEoSrvc8XAu8PvSZEJWjQPW9UW5jhNVWmW
kOtxTEJArpEj/kFO7Wh8WQq7aOsaKhrxBkbAtNQGjrUId58PLJCnKYg9HrTVl4Ue
c3YgJrnICL5LxkRLPgW9RXXZj7XtweMRKcXpDAlJ1DjJE57jogm7Elu5Gs11Plai
QEBr2lECnj+xV/IYNjKKrh9GhH555RO6kvL8xFWinPL/ao35DMgBEq+7XhK3tnxm
EtzgJr4jG9pMCCH4yfA0R04xt4eodeUAhd6GmKtq8YmHjnNQ38uV93loVYlK0hF+
54KAzVv9Un+Nh1rXI8AuiILARxni1yUa9yBAusPd3/69bSrfGJ2h6On1/9lP4zUT
SMf2BcuzpL6hCxtVsAXg0QkS2ypGvCZLXnC01OpeMmUVmdiUOvdfqhvPUBKXbGTx
l6yAHtp1W8eJXNogiJuhHghQiec4GBZzWm+gfB9tgXw9PtABrDCqehO00jVbCZf6
7s7qwfSHbsqd+GlXldlzjHYr/WEC087lR0cAXYAlGtWOjBmmYpudqkAA7GUiqN6M
C3wGowqvLrHDVWRWgMxJVXsQUm4xG+D/LvHyMofU7pEpMNygQXfq4v/BxsjU/bzY
JznOw0L1NlZza4ArCAyE8Nrs7C6GEeBJhmhkxuGmjjP5iBYQwdHA9/nj0e0WcfXX
6sXMJ9e6UFkpxsH7CfTrK4KqUnnWTfyk3wYCA7D/4J/mZZc2kvcC63wMPRD6Hn6M
WvXhkPuW6DeJ3ddGZHheMJyJeLUpF7tbdRCT1Guov+gV47x/F5hDTtCZgyivWFu9
XxF7gWMWUHBcsroBGgyr69johLWzpakehO4q8TWUL0jFmFSZUvYi/cmX7kQgWB4Y
bHg0BwSq6G2zU3kAqWfdg8wyPwKUilS7ZMbsC1RkxydxW5GXcSQq7HEhPbn5YgW4
Ea3oxjCBITOs0uxqxi6Kv3aCsVws/CwpHwdbe8ePK/4EdhoKnr4OWMDr690DRChb
BgHiL73OwufBMeBPbNlU7+8g3oCoytwJLajhv43vHNbKIHlq3g2TWx0vJywnpza5
6Pu2idLOb5as90s8fXnhYtoeMU/y1FbBMf8958GIu2DjYotD5iJB2x5Sd4OY/FUG
MRZKX85Eiv7kQAuxl9jDrqzNy6A0jZbJO/ZKCTRvDOnfpe1xzXQ5QfoObrBjC3cB
MNwTvdVr/xPf09M91mtmGvtZH+TtzPScG7XwycdQV8qqeLVbCFT/rLHZ0tSnN6Qf
E4rOGr9O6if9s8nuwG73SNn1oFHrcYMRGA5CGdjpQzpUL93NhgXbzbX9s1qeebem
4UBHsdHvLRZyzFy4vx3CxQwfjLGXbZISoRu/ydfIGl55vYq17V1TBwhrypFM7ejG
ExOaydr6IxdUgR80+RirSBGOdK32L3J6pt3VJ5U+cQoOzeLZm/jumxtBab2YafAO
KZfXm8ORKI2JnOsC48G3+zq8KZMXPqB2f868Za+wfSVqyOKoB3DSlPUfrjwaVann
l7jpf5cM6ek5nKDuTCWoh/hWStrD+eed/etpoHAE5cvnyx0V5GbeNNwxWVeSrSCH
MHZ/Du/CgJLHIa8StM3OAaLWndm7RGis0RQGgTxVrfz0LnS+IR5h5lJRao15Tvio
084nUyWA/Z9rk4XiBIFcIx1yUasVskDLDs7+M810HwWXXucSp2aZxwWET4MzSw+I
WSV79h9BjqAZq/TBA1EUTQ4ZcePC/1kkj/XDj6MRuqXb1WWDDrBtEd4mlb8mRqzj
f9jyFtLXgpvVDCVH3bMGcrxIqnJ/HKA4rVPs2b1h8CEuHojZqThUWpNvZbY7U7n8
R+yK6QnEGpCvNNxvqVJWYKv/XSHeTGyXcEEI1+w6vfr+75Sxu9O1sX9hXIKFpFEK
Zb0tUJ0M4EHxfrkH4ZcIq2vSc/2Hdd4Sqka37t8f8s3vdSsG1L7PEepgQKt8ckZZ
FTIPr6lXf8l7B+yMzcCOUpUifcLnu+gx9Kzkr3kFVD6kqq/kjM60cQ6Rp7easJpc
uuoJRuo6s68zuLQGWV/vALnPmd+Db9GzzzuJvo5KoGLfV/fS7fMFmo0eobJj/9wB
5ObEQgNrM6dElR6qkoc2b23TUZ0LtxCmVAFCaWjyR50FtUnwzg2t0GqDJ1mUM9Ay
yOE46X9OFRcqayxIwp4VHPqRZN5Hn+CSUtELkCOowTMuJKLGropYY3piOhdQRj2i
UqHR3aOSxuxi5JHu1uaR3OpyI1wWSyM/mqIankv11xfNEVyBxKWwvVFzaFrBuZ8E
Am8PeA7TJifFzp5wtZG3LctpWJI10tUlR0ubhXNvHoSgXLnNvwc2O8GyB65S1OSB
SMPteTSpMgv0YTjJrizBm3bOBsOah/JJuA51ACnbBZNMZbN2c/UulAoCIYmj+26K
qPIDDUCzGW09iPnYn1tnpGW49Qjh976wxFFn6GRrSLo5mSimVUkVmE0aKqRFDc8i
LU7oMju86M4g1kLVy6KUgi4UbUWE6Km0+OzT2tm55Xp5c8Wmp2kR4i16qGnBSXaB
eBobLX4k+ZQ8ncSia+xKOyYUsQ1lWwim1vSAy2lyDPjzZSwnIw8aW5F9fZM9UNYR
lq8Bg78XItDuXHGniEDvvos1fmGLLXQdP9DzH5BHOrNgDSihfeRnQvyo99e32wOZ
xgU+8JCHa9t9oNDYvXcMgGmrUIPrAhsHPReUjnRS6S1Jz8qMfFxRGMm1zNrnYzC1
xhPgsZob1fMYnLWzXdM/qSpaVMSjV8Yr978cLabieILmxlF9ZeRisjWMf/3H6Osd
XEMvEe2+dUR7wvCdsDrXrBuD9A0duk/verfqzpeSlZ4AOyaVJS+EIKrYSlNrePlp
kqIKJrss91smvLRQFGTZ7/jLHiBLsCzmMZxuHOSJF0nSRz/Fa66Lnkz/XL3NIn9W
c9baJvfwm97lEkheQmqxgMERXV1wSFyHuxGNslPVIZ1Bqcg7dY9jWzlpkB1O98NS
lGQZj88/5Kk7bKnhqmyQJbHKHfU/VEY8uE1dc1HHqgWwtyJjiaOOSPdo3DNYIrqz
Ds0aTltgDN1NkcjJc2cg68LPcs2Y7L5sUteNGs06uVTVF0SMb3jXG2nB8V/zz+3P
+9PdfMqlG6xnLg3P7Z57rWD3PqlwvDZra2b8oMe+aUN8yQeihUD6omkP72gvmREY
G4t+i6nJ53Jolg12kDFH3frEEB+a/ie2YO0PNDfXYzMSl+5iwDykX3r37X7aSXdd
sZCCCUnhZixKI2ayoysqBSpn4ZjvFs7NPC9GulzFfrNXdS3kr8qBl6EZEJRdlNPS
PtH4VYxb2bUvGSJbwrFs8UIpLCm2C6YlY3KOdN8SfsFhjT0IM5QDasBW1wrVdAT2
Geo6RuRr2OaiPhVik30xQA/rEMcylojKsEZIVE4z5B5ReIGpJ6lzOfhW+WrZcMOq
QnrQzDxsapbgPoY+vUQj+1uWPGsQApoNOo3OVmkRObhKc1YDXOBsAYBnCbfkuSFR
AyVBLSbdHouHj5K/D59NubsDSP+FOWy+WAJGjZQ7ZgoBB4aXv9UBiJNOcaiAa4WY
deM+c6DKHvNeW63uiFNid6LHU4Lwjw2QkuribwXJYpZi0IPH0iki/czHa8vV3yak
vJXZYpIlXJBnlvwA4ZsIu/3ESe7UqsGeIinakSxOFEieOtVXgGczcsVySbc9E6rU
NoZEysVAhZRP+5es4zJdkFOnQ7ysIW31tTS3Vva1a50YFORLC4iLUCWiTJGVcKTf
UlkhcDPcaDqoBbrsa+1JEyNHW+gGzrqEBPOmuieyileDasC8XW+PpqgzB5NnO0Wl
X3LpgJvGnjPtWcLNgf1B1nyWf3eenzMLwSsjY5yn0wvgZmhXnW3q9LYQpHpAaYN3
r998KKCH4/wIFqKs2VqnKALLTThgTheAnp7OhrCf8gDlenVzuVM9USs9uAFD9kJ0
BzSNFkZFzjXwjtQjM7vnv7B4EVmZoR4QFh17B9ujwE17bOWY3gtAiCQ7rfjb1oeb
aQ/eQL7/uG73pKb2Lo/Fn8VAaZnNBIWyekYT7XcAMzD1JVjtnaQmlM268bGRk0sW
uI8S3XnWoOPo8Pq8L+ztGsnAVM3M6cdKhKMTV7qCtK2e87mWjLQJqa0QYNQz5K51
i1oaF6d8NOYNYdLYp1u9qw0I2LXzHX54YGfZ6XTPeBx149KcQsp5tTlm7NRrNkS1
9UtT8YSigcyeyTEALXHsO2Fck8I7iDQLIr3F4E6mB7U9SiglkJ4ddsqXlBavDE0u
zKL9eqMpiJ4DdDv5hMV3tJzsaH1P9Zk/wvaLuFXLUXWcfa1LnzB+bGoxcQOtyfRh
OX2wAdAXfMX1I1Fg2AnvqvvoS5hh1YArgCxdYCtpYmiKGSzki7rI07lfSoa20jQH
RDle3t5WFNUxXI5S1EVFYnoCjpxs/FhJXpIefQSI+gHYnh/ZwjK1TaEtXUew0OdK
lxqh3nz9BVdJy8Z2G06xbRwVWX9lTcKKUiZp/XmzSconb1Ad9rg+y8zXkLUWHsFe
OWpEFRyihX9omCyE/00J/8wAJDm+9E+yaCSfx8wYsZ6fW0hR4URGtdHz6+3uvFr9
FUq52kw47XfqNqJTZ/lSPegw421k6vGT2TYe1Oga20YTIIvz5Hvu04XDCtVuoFzl
xGyIvIItlIzTaODEzNpGrPzy6x4NPgkuJZwzOUh/kw70Wa+pOAGP6eygXU3Se5up
5YzleXmxTTcJGtTR2f2zCX7a9caHgbDzHV1UXt3tQ5tpmsDA4yKsaF+/KPQUZtc4
lRzmlQUolftX1wMUQFvTklXaR5uUTVIAAZJBj1Vnp5zCeiqqqcREKCEt0Xhi3o6c
2b27nO1YxRw3vBEzIGQ2IS55OIrsQo1HBFmaPUJV3FMQHm4GakbV5LbQOYUsvrRM
tsGmbZOknNNP19gaZ07VrdPjNRWB6R5K6KiIhQ3TObj6fpFuHtZk94A1BoZWBTBC
JbF//9POPRHWDPpPvRByaJdBFMYASiQUQE6AKEzW/p9+1Cwan1DZsEH4C6Xnd1QP
MI+KbuIczOgrlZsMC2aLcDaOxkwhqRK4wujA09BpM7cvShe8H2uvcbgjgINx2+Tp
e2QK1T2VhFMY+0v8tu6XmqB2g9nmA7RsinGl+vjVKLhPg6F2cmiWIEBCjuqRrCvx
sJ/joyqxwrgkBLafKoz4zxLtgXbX3LNwKp1xJzY0oZd9tAFWiviVfAStFHFiY36f
wFbYFb1t6ir7/qMzNZwR6iiwoYkTIFiXTSnr5S+qbEA4Po9nv/4qeGve+awDy8NV
PfBDYKnWQR7gmGXl1wXYFBu9MX4qPmAI55thImr0rtDSUsdwgeBIOrXfc5f0LwDD
qyIfQ4nanaNGENYQmkb6lXLGf7Nt4WPY3ffe5KhUlYTqnMPjz2t/b4uRPSs26AKG
hgENS/q/K1du/Q0YtmwfMuDYIedwXKdFdAVeBunH2haYlPtGOJ6HipZmzjgzD3pV
7rhZanIGm/zchIiGnWVdPTadnhFy0i4LyG73hAWuqcOLBtaMxIHlHDpRmWkKEB3I
KBXdVktLbtBYy0A8Jtt5bI9cJt67iTo5/+ylJw0prxg3S4VTtnz0GDqvTnxTUav7
b74wMRzqnipmPCfzVmVyXqhhfW1hbALMycd+VCKcVex6shcmmffzCDjZtFkmMU9p
odsuuklfuZREX5qq5JKD7TK4wAecXGN28tjYdeRgO2ft9P6oInGwSgSj9pK3H0+B
z5l2YmgGGaDEW4X4+4elXOTWjceUfWTYTdpwDiNYKgLH+RTBINPCblmk8tqvsiwM
3j4r8reJN8lwltzAPvwomtEQF12Aj77/Wk1gp28hWUF+uDIb7TGbOjV88oKZjqCD
5g2AXovDALm163ZwiBNm0twGktYLqojv9NQzUEaq2EaXUE3ZhVTY+veOPuNjFDOs
fP+zrZ+qgKpPRSIqAU0IWMrXjjhNl+Tb4cd8st2pVZH6hQcPyHSOWVY1F02Jittf
8pA40FFtOQXCxq0pvpLkVLPRQOcFP1Dv6D/gCJv6nLD4xx1ocbj/8POlpXEa3kvd
oS8djC0VAlcPKEQvt/CCgGroY+g0zKkIVuu/rY+1wgVGXtjP52ueUYELh+POsYOo
gtFf4J4Gi1vArOqo9e+kfQPG2QrZWX5MiKYIASUzcT8bo95/J/Db+23ZxuRIDIzF
OR71HBSeTs6s8ModLh4N9CimoymCrbtpRxkpy7l059p2uuDwXsDbdIoBspREF1Nw
JOqTXJhPrerJ0XeLK2u/g/0iqbyxK8cap2vzroH9rvsTOI1A78iYSksQ5TFW6KsX
9tYmt+1wj1ykCOwwda28FptFTvAn5H8JHn4bMwrNlBnYzJcj6WFxhTOt1o4oDig4
U2yOGzJWO/bxtKhLridtqiXRI+hKh0yTUUudX9lp2pHRROiai2ATL03SVNSp1Z9X
YwNflnlVFtcTp28UcorMlrIL8qazaNJ3TwdowyJWaBqU66fDSOG+kgkisglv9U8q
wwMgTz3lomr2Yp1UyR8qKDs5++xiipzOqTFUEp5Emos8SUwgnf6Mi3J+Q8C61d54
XKisR/qKCT9Yjzp1bhUuV6TSpI8WMTTh8MPLubv80r2PWumLx0pGsAJezDpoBcEc
TDM5+zYnwWnYkJuCwA5IUo5FxniQ7ZVNkGDgp7Eg7FIVUZrOKvpSVDS/KhYQGO+j
dGKYdX1TxWo044oW/bWC5lPQyVVDciQ/l9mOa1xYC+ZwunENlGuQqbmvaizzr/pk
Qha4yl9rKaBzTbp1zLcesT0C1tZ29ZV7pQfTrsxl4kYDO3hhiW/C2OiTFAirASpl
BdDE6bDmupCvLoIdsoIUrp2se/rUILm+YL20o+CBqLkpHVOo6dqda+Xdp2HRZ/C3
hXghFOVC2lJSimpkaejG4rvtfCzf6PHtCI0sy1GRzl9+7at41uumJ9AbmU4KGf1F
wUY8zS/INUuvpYzUGtkSytZ6S8xoolrDxoK1t0WkXiyLjU+Z9FoKdwB45pLr8gUF
gK2DvZm2/3DdHGiCedQ2PlQCOAZ1aMgNAmQlxTrmHOscHsV3egUfByZvqwS4zA77
MYoBTNN4Ww+bg+iiIKsqXFFVA3ZaBpzgsJEx/hzm3r+2W26VYWdy9V9GZHNH66Pv
qRJOAbnSz9fz4tEEP9itHbkNVISbExff/S9cWHYEaapCNtD7Oaxizshl6SjKCaib
hu2xl4WMhPwwbkZBhhl6ZuS8lhpn8g7zFbCPqcxmGT2vrAnF0kdZm9g9pqjtmALO
DFC/UEZHh68LUZtSN8K6lIw813c+vgWwnoGlvi+xQ6Aio8X6D2WFadtPGdQTepqj
Cyd+Ae4jgSZGe1YEMuZejz5nU9bFT0XUp90lMuHG/Imzqhqm3Z1hu8K0ivNp4awe
lpH5a40zNykm/5vFUAXY4reIF5B5RBTcy+VJZDK5HUbOZO7PcnAP4qXGPXLvzn/O
WsIq2n4wx1WzFWGASjW2kA0v2t8ZrSMhqcTAI2UUVn/NYlislI6lnyEYAw5weW8y
cgyzby97KHks1wnoVAv4EFDVoYffFxJiB1ZmrTwJCSbAf+Wh4yqqeZTqzzc9m15v
zd6J2Pky5vY09VRSGy5f//vZ8VkSE92oUTTjE4LE9Q8K6rwyp2AcqLowW7Mp2kCW
3OliP+dJ55BhN5jdqs+bYxDu7kjzhJrD2ZuEneOKYnO3/CIIEoSHFN4hlgyMxo9H
TFvG/0ac77rfiNUbgwoSsW+ck9kqAlysfPutCwub5bpbhpKi1fCIJktRrptTQtGX
XplF2ZaZV0XuTrqZWUCCZTNBdVVl7pzpMeWIj4gxw6qhxWpegwuqmJgYbsdLbYKE
nEFdhhyK326uadFHBORAPLRpXsXNCdUkHg4wpqiTF0f5T29Aq7J0dIf8VIXUy+O3
LBru/VGO8goBMcfhw1fby7ueDcpVgc/SDO81+cjILF6NyDltrBy1grIQzz0Pel8E
R2YyR6aDJ/r/FJOrF9YD436BHo8377T5+khCsNTMtojTOyQbW7Z9urjwojsDPE+e
oQzMGZQY2xvuvdzA+q+ZZ/j9ElKAAmft6ukoWRQgPrZTLYqONrCUJtl1M2kSTxJV
WwNLnI1fIqPj8KKzTyrH3XtcdA5KQcAyoVDR2UJQTV+q7WoXJ2GtUUFWkbVXLd6K
1+MltMipvszty0CkHY1ItTRQRNM8BESYDbUbEP9XZftwHwIwtIZgWR9apjs3icUR
0GrpD2TMbsBzntq4bp64bXKLbI4hpiOVMhPdjbwMGqH78RNvyY5O//q6yLwzaPO7
2owkJvpWVmk+CETmKMAV7LtE3Is6b/bC7UNbEbT9WXUzOZlsg5j+J9MRha5xzIkl
UKpf9hmuhDauUAHZCyFsSxw20pSoSHZ8DqVvsGYj1FKLexDhYhh+9Cihp8fcmJlw
B5Kqsdrpqbtq1oiLftVQIT87e2jGQaHJ1KrNoyAnY6H2W9NVA/wfarglPK3RR2vu
APFYA4VaQW3jokAXbjgw3Yx5H9I0h9K16r8pedBa/P2kklRvs5UYsYsl0QHF97RN
CAmhhZR5jdQA/riqIegIR7x+MM57v8DIsxIYd6M5wJsd8upEstUFnn708C92ZOI5
7YXVSrU72DRJp/XW7ATnYnWh5hHw5Xrn975t1ELeRkiW+ec65iSnVAFMVCYzbydj
peDRwMxn/1kSXS+c/6yks/c+jdR7C1a3HkXhUr0/pSNth1vfbXFMi4ijZd/QYw7v
9rdov59zRaPLFotNrVK5FVxh5764+bvuGn6H9e3tHIM2dVKNbYu1Rg/AMKkI693a
cGCpS7XQ0M9m9jTfiwKYUCZDBtF7ADyd3cmQ3/+UQwIh9lj7u8XqTr0gA2RrV1/n
Zs/ZhjYtmbGIcETYR4Evf9lt5sISAkh2IRXDLwh/jzjEpMUwt3f+zZPRTWWTMAvq
hnV/O3ounKNL+5MzN0b36ADSHOVT+h+uwQ3sGRwrhNLl2FA8NSn/Vq0X5GAryQKR
e1SeUwVIHMIXfQzCbpHPyTvIa6Xs0g/Uz0qp43pQT10dfWN2B5u18fUpa6DIsGuO
BZp0HM18VQ/oyoAwmvcdRe4eGmOLDW2quvIR7vOLx57Zv5mjVSxekf4gwoPMynNB
25xFkI2LOKI/nYPJLRdLjJyLr/hrnLDP3t+XFfmj8cHUvbke1TVBO7u63+h6NCyx
RMi++aysjxdBHMaCQ+M3eqo6AX88rhbKOcslkBVBTUC1AFM+SiwJzuvGIrMtjI2l
bXOUNU5ebJftGWhE4msQECQIsuQPIUXPqXa3GIB6F3qqjw5twXkLYSnJkZGgGY9X
/73SMA0Vnex/yLDf3dQOGN5NaLE0n35S67SOUy23eopb1YAgl1vVCdmNHbboDbf8
mT7HrLP2QnB8VbsvIlsbXZJDGFFRodtK1qfJlITd4HNx9w8b2TYg4wQaNvLXizt8
EfVhs/LrB/d7f1YReFaL+aQ+PsLZUHNx7ICN7sX2N/DkgSNqTTUhPg6KuiyRyYiw
SgD32WVFXsxpBYKj/m+KB1cV8yznL/wZSX2a7fzeRWk4gIkEaq36TlQkcYseXXSg
tgMd/LLPIb3e7Wgb7lU4fj5MFnzYyWGvOuC24cPVA+jrmf94g9ye/8V1lxArpx6Y
deNRTojJkvPxeY7JeD2tYRSG6ZfmTkYjB0ytUns5BQyz/t+PUxTLIlIftOuVYUpU
K1aKMvjYUOTzCYygtqRo72yc0T/w9DJY7tRzIKanyDAluDRNUM3sQwzGYQ8VNuHS
b5jb0BLRgy2inDYFniTK1bl9B4Hwa2EvFfWu2c/VYHdeOUjW1giHYVAOGEf65f4B
rr2SG5jZmbDLsq3z9mTJko1wADhmIisL380flOnHr1b6y9YVsk80iqieCz//FYFg
K4UnU84LOVkQuyQVH3+AQcq9dxHXy0XBt837qawTOPb/YFFED0mWN3CAGy3dgg7F
2+mVcSr7yCtp/COBZFSuqfDKVV4t9fQ5f+HO9gsDdW/XtJMTpdnYcbruIWecguhG
6tPtWVHRHa1+moy/rtsQI4D5YOnyJ+eMvNgiVdpRKov7rtPkGhSLT74Ez8t1nRNW
8KoWm8GBMBcRganq3YiNdyDd0s3pygPcEArezx64CzbJY9QwoPo62S5bYjkd62Mn
6ASQZ0/2iP+QFpoh2JN0L8YGPn87ue5sik4QokOR1EOsZA7Q00GUur7OozqxrIdJ
FLMISK5pQXtaW7zxuUZsf6RRy19Bj3x0JVvXMbNvLP6lyNd8urghAZA1queQUAe8
ZBRDxKZR2mMyx7o27ERysfDNjoKe/6FgXjDQbU7jkPsHXxemr6IVp3TPQfGHLVMw
ezKTefbSgzzx1u2hvkBIRxFjija5x+3p3RGSoQVt86yx4pjuTcsQiU+P2G/kEoC7
SGfvhsRoVQ2D/mUe89HbXSRIJa8wlIAi69A/XvG1FFgsbmLm+05TgIfSqym9wGxM
yOe/tIvOt5UruWzD3EpMmxJj1JID792Z6RqNyk9ahzVWpMwBDYLv5kCBIKFuKdDa
uCUt+zCwfco2x1/y0v9TGB3VLW+Yedx2UYut12/Bkia9MgxhNWSjVxSGWUa6KDzV
xxKBJsgf9Fes+KH2kpuoBPVyTIM/yCHyqdAoMIkb0QV+eo66Fp71NSYPJLejHZcr
xr50i2VPxXmza5Pz6EguXh5+HJ/YzyY0sJW1hcVM7J6x3pEHH/M9vjyqjqzdz0hP
uXQprabD1yK7+foOehoB1pd/yDP4/ILuacJ1rV6T5kRpXVV3RCpLCf/8XhNXCznD
gcoe7DMwt87l3Yaa+EJcRfwblF/5nFuWLXflIgWZLJUXMzBhwaJTubZMUNqPd8Pj
Q5zRx165JCpiAdmEahXQnlqMHqfq9oifpS8K9J7hjuciVoyi5zeGiNQH7l0+XoCm
Vo6b3eUmazG6wUuEp6xyZEJZlvwXaKsljoZeRSgkEzDK4va0psJD1nhQZKTaI0fk
VHtyuy0rUEbUf5Z71k2D/40odwxoKXxxx5xA3dnggZE8WN0gx4X2BPgjDWHoI/d/
ATMAvTpvo65FX/4kI3JunSN4Jwtuv9wm21WPJPYXUZLUDlPyh3GPuHBPmZua2vuw
XKVigoJrPc8m5Eoj/ykTonOaS3zucTY97aJmPhWW1OeYpT54AHa2Cg+D0Pocl1iJ
KUhTDoccaHDm29uUDmz+/LzvaLNjYt75MSHUdQNROyweUnddN0hT3Ur0Snw5omKY
YmoUGftTScx/SgfNTUgHaCOj+n7dDDElx61uUFLfC/PeBZBlm9JoKsvaBKewZEq+
/xNqHSKLjt0veQqm+0OjRQ4uP1ssZ5DPI2qP5XWVHd6LPKAowqXP2kDZJdI73QkM
/EHiee1HXz45q1r8R/nyS5a+LqRrbQmbktHPwVvUMUr6B/bBZtyFY5JCt4R1HUYt
nluWE7+IurvHp4X85VIZCA8vOR7O1U0pCdcQgTbg2CC7iXlQ5gVIc/g6XS5okNMf
v2dxmXyKAsPr1LrcUGh+QrQvkQJeN2oawPr2eXUJSn+FRfy0cANOOwhfyciuaZ7e
ZGw3mjKacIYnTkstJhQUBmL6I+waXWts6Q98TVnaQPyJUSKTFt4AG4ByHA7tv+2k
usEgsjV7sCxfmq2Xiz6qMOulGVAu6EKFE2XiH02mUBAlfuQdfUH44fMc2xM772h6
kBDe15vsMkbTVsRWZOzYBmq3KOqtCibgbcBZ0rW+7zeIjrqt/vDVEcNDSGuzPIj9
UJiPQIPI7V7pywKE7VLxwM569GT3ihd4ECg8OaxDUylKSj1yEyKlHIYyAAUB/tkY
ANTiAdd74fwLJZaKTtZTVKQyMWOKkCawbHHmX4AmU/zhYh3cfVwv/mvTF4MQhnhr
CEOS00+U97RB0jf6Kudogd6ZJ7c89/sbWTxp8UwKiA/s+/Wc2IyTUPyPdzzFMu+W
PjNXrGWhw3S66LKxyJsxmLEmf+kNJCXhpZUjAql2Bmdhyc+lMSO7Sr8/yMhdqfEI
7sU1x7KkR+lI0mn/DDDclYRv3IBhqF488JyyUkOa5Cy/TtZUhdlLoTnRnStuQIwA
czP7laTOt//HhPcyOGlLfIulxl7XxVUtsdkPbhARBeTCAYa2JEwiGnt+aa03L/iq
XZ72YwLlUr60HFi752MGQ+P3Y7uvZi1PLiq2UKhq4EgNTIUfX8MLNYYizy3oeBwu
s5eZP9a9GSaSdw2F0Sqh5Ntj+0OtAmHwAKB7y+CAG9PneAfFdmqqteAoe8ZJvp8A
Xn5hnMOsEtZpQKWsqjDNVY1NCcy7ge2Tn6sM+ckxcDELkejdEIl2ad3v93EapI03
DxaDgeNQW2dWt34OQRCZPc2LsxLJDoSKh34VsG446Gz8zwPDkOLhKuyvJO9iLWzm
vCD8ZyxRudIjXxBRFyKhaQYQw4Iu4jB5O3JnaExy3Dt3HxRtfjwcWnSEyK+11J8g
DMJeEfaYtbQZ8gvOMfJQtGM4Ak1imgE30UsFAMsVhXWgtxBdNHjh1apUUGPT+vSx
D79c+jk65+LpKZ4x3QSI2bz19tpFtcBAZaZshQk3FWWlUlciQsrxJglusjfQUu+8
BnTGU/5fNa6UJo5kJFyTGX5888X/FXN1aAPVSq69qJ1CtTGIiWFdEzdKB8/OKQF9
p1grfi/B0wDr3B5Rhsdz5AaYkN5oO+k7DTIbRbR0kkm0mo1fRMLaL2PKvEKbRoad
I7i6CkylI6MIfvsRgPT3Y+zQVnYgFGnaGehbf9IkKjaRu5XzJI04F9gE4j70o1ss
I4kGoQpMpgOfPX4wNSrefNgWO0KONPLaHo2eJT1eIWopS1mZLeyvxo6XqizckJkf
+Mr3MhdTGjWuiY3SkcqA/NJ6pgbOLivflISSWqLC81NUUqVoQKhCWhAQU5bbiiAj
jsGycW0XKif6urbsDVzMP17UBjB/hQJevctwCan5wxZFIx2IG/MgW+FV4i5hT2As
0rwkYKnB/JH7EWyFjps+Y6QuQ3ncSXEskAS7o/DSn1q1DvQJdeNULrc5+QKN0nkp
jXDdGwHrB1Pj0qmMtc45Q5FtmvBUHtnMSZF/edddpr09+Splmakf8l8utQszjSq8
ZWIcdq+tSGsOB3KRSuuzOlSJD+AYSPeJW1yltQXhhJfhWGn9I2WclWTm2dp3GiM0
+22jswN34EcDmGqy2N7YIWG3lWlumbgCrFdCv5FkkfdzWVXWTG9GMbVwH4MlrfsM
OgQaXF1a3qnqllIqK9RHrwxi5Dyc1papywyg8yiN4Tg0c/TJ17eNFRrpTTJBFj1T
k8TKIzeUtlhZIFQpcOnY9bFPcCW7jG3cq37nY0MvyJq96ynjWHOGIDY3tgkU1L5Q
XcmLXv/MuXg6yw7gks/uvrsJwu2nsuBa6JGWmX0o6kau9/ZAt/GBR5gpNK8lGRPq
giZLF194BuLmFtrD4uglhLYx2G1DcEj+aZqA0UXT9ldLba+QSlfTKLpWgKH7qH9M
0vwr2tk1Wh63roNG4hn7A1CISmrERiWraO8eWFSMEIa0ZMfb/BIazI9x3CW4NgUN
ZqcEiyZCjSqb30wleZtKnlkI2kDfY7mFC5A7+2voU56MBLORgpK7wsThLVuRtYj7
Ttocg9uBDCjQP+A5puMYtP2hBvo6ZrrBtc1BRRKPHM5JA144p4xhQA72RWpwC/js
kxMP5cfYIdip4JNvBYDNgcn7WiNXKnYQtBL9V0uKvD0R1RD14fK1juCRSr/jEnjX
IeNXvo5bRQwciX4oZwqe9MruvY7UptCqAZ23Xl5aW10GuvZaEkXbeR4j4zpl3bDS
qjMAf5cvAX3lXN/Ah2caJaU3j0OSM8W7hH2BGSbIv6j6+BzaaJP1/EyPDxkTuLzN
LKYItSr0t1GCOli76B1U7OtbP0VV7VBy8hyVLLDCPi6aZRxhcGCPTk8RxoCKkcjE
P5NVjtk5EGcptnG1EoYiRUH44Se5I9UnBc0/rxhaqXhwgVVsI1wURrNvq71b3SNT
S7VT8PxpNuIG2Y5vtQk4ua1EVN6blgLRXJpCv9CkLTc0GD488UUm9gYYYihFdcC8
1c2IOJHiypkIs/kUv69IFZZJyeGGi0ZG4XPHf9v2WsiLp2Iwvv+c8i/Esaq8ocqW
93qtzNpRD/jRCwExchCAyVChGCBS89yIg2knuOLV6nZKmarqyxSHuAQX4TKDSwMo
CxhHiHm9Wvph1tNdNfO1cD8TNt3wWeOorNsur4yYJ4ErwsBlX4HOKliYltwdVqXL
kLPw8AFyrfuS2hZkkbSRAyQkYFWJLybA96XRSQZUNR0+eNrSDlbrWLJJxsUKa2rC
vynlCrODitQApkhSb5Sr/YjdNHmpRZCdNOOfDLp2zQAnDhb0Wn6DcnUqQpO/rsDq
hm6zMSGhaUt2FOw3+E9aKNdnJmpzx2bdkaRxYTdLEXAG79mMh8T1c4eUJ/2lH27n
Rmpk8lIIaJTbkIVXA2FPRvmjlnsyZBYwHj35AmGJXEWrrXxqzgRslESPvfj7ko0J
ejRhdoEWiF+siKdKWs8qZhgX0rrgg7f8Ss7U5kxrcv28SrrfvYjTQ0tOBacwc33B
F/v66IKPILMyVTO9IEu7ONAg9mmRHu5NbXfU0NmYjnkhFEfBBlO91mImSvf9UR71
hnz8EZWheVuwwGhHU8dkmaD6yZxjy3vWV3Hr9c0yASIS7LOaAXU/dyiXrw43oSZI
yhCgveBDbJYL1ljbwkvM5eaUIvBJ0WlKBJUao7xpUrJ0bvAhjZTVFyB0rOwMuqM4
ECjiw6ucvX3DOjCVVZtm/XQqQGEeAKbKbeYY4PpP09n3ZRDClrjrMnr75+SP+0Cr
8HkuhHZFGTf/bMRR0c1e6i7/6asK1arGnOXVx/ZMRFxTHd5B04O/4Y+v7W2KmqWq
nMUaIKUVwOiSBC2QGa/7+d+kyBawGEXfGFCTyAkJoveJXfPM1anu7zSIQPMunb2o
LmVBGRnJNrcEkIhlZRZ/OS+y+sc6NSOmrPIe8PZ2E7Umn52TitUCRZWQpo6I4c3X
gbnp+aaZjNiLfFuSx0BKz+ZlD7Voi8P/esAwuYZrYWvtIzgrrb/PNOH3PUYaotyP
Ye4ypnlqn7taBAjo6JXvt3ZsjVZTEAV7vwsFszOAH3Mh19teirHyARvIq1GTTLFD
0BeCoNXJtzTGihVpHjw9FtEVb03FTk//WKFERNWWuPH64X9ao2L+dQRhA9mCiPHH
ICUZ1lVoxZmIrNGsYlwu/D2mQMU01B85LVBZHRYZU1sHAgGhJC3c9LR/v8+94x55
Jad9Tht7Jq6PTZ3g/uZCnQsyyfrVLGhQbbRdz5HEfCUmUQ7Io0mbD8oW14si0Rqa
4lGxM6LXccUtAgTOgU0boKxNfJ4xxEV9zeVEr2koJo4rJ4bYN79giHhLx7HEuF0g
lll6BdExzqZW6SKvbpMqXNLHdxDzzUqdtoCnglCbNvCAUPCryU0katUL2cT4uxAn
wwbmNgvVNOA41ITBnje9FffTbieWW0NOPhrcVUuMIYzo5WEm2dC70QiMMii29XXC
z4tRm7V85hKnxsdM90R9V6M++8UCo9GFcFuSpQtMxJM4yTiSJkHlIefXkA80uwWg
4AcMeuCZ2nC8v3LOojWdpSlz+pbHLhWzzcan/QjNt4A4KWrJTh00orZ6JK9MaDrv
ht+WFNiq1yU/zC7ivHdc+4Q3DyNYtFXKgrdyJ6ABw+lNzmGIk9BXXLcl2JGjQYgb
occWfVMnIl3wsZxa7UWELrLrT9qCZE1OZgMPFD0BEPi1/5cLZq6hDMOmCUfgcYv/
K26a3JhocwGQbudAUtRvbVxUYY0Legk0ZGMnmInFMZ956hCdmGO569P+j3qnQbIt
NtiykGQnAFivXwBuQYqtuCM4a3qvQZRrscdMc6SvIAdzn7LFjCwWi+KxYo/Z6/Yb
QiG5Eod/qyMb44z4WZBRu+AM9polFbBfMUKJmYvIVGUJ0G4LoknhSK7RCtwxiU12
lB22GODd5pDJqHxm36SPIArwT7/FEfFciNbRvxCSb4AcymCsBXjiq3y0phQFFbXL
u2EODnEuMXdymYjC1GVilZj6mRODv4l5c4/BjoPzV18eFEGdhGyYgiKji5LUlYPd
eUpC2T7VUhr+IqbP2IivzicXiAKeknSwBlGT3y5Q03gtZjHu/Wt/W5Xm+A8UrV2T
+mTGkOxGQG24izeNjqEyP2sBCR+RYNkIg3W2vyiWmgQVfkRmwiPJuDOuStdtt9XL
44FeCyL+ZAVfwwpHXDEeZ4KxP+s5K0FgsS6pF7f66xDmYHRGP6svY1CAjv+QVFYB
V8sACE7PNs+lmCbbiTWCiIIDY2zDsisEx47EdiVTXoMUbsmIRGC78Mi2JZWzucuu
U7PsI2r0R/QhuiwF0ti1ZWOb3Ojs/NC9Xb7irHZsddoCqgBbCECg8PWmaAaZFupm
nCy+y3ORo8RIww0Z9PlEORBM7LrMDzBwBNtdf8QGRHU+Ine5dLb7Yj95pPcTN2L+
WSG2oAo3V311GHggDTWPZxDEsK49gq5+s3nZAU92WOEomC947KmMRDWHMxriZes/
ukLhljVevJLC7o/37RzOZKtyQeonP3iAqQKiaODXQ5QAc/aSTD6ouK0M26eD2mEB
iLBo1L0GPhng2lv4gD/BK6v8SiLqiF2eErYJjRHj7eLJgsPw8GrlNRc/dtvtUPMN
FJzJpdRBj3VFyUwDCIr1o2qB/TXYPPcNSf45MgFQwsYMZoKyGnuAaXk4RJrj7jtI
CLqGGKmoR/6Ts+e9hSfwJ+HOo5N322zDSM7oXzKoi+azBiyASk/LDfE9+eKChIlk
dJx/wR4vWGMDMi6c7UkthhNSwMvTloE1mncnqBQb8x+8QvjXSeHkIosfCKSAJXT6
MbFPuLjQNwavHhYbaPG0ICrKOmgBkvVVGoTjBUJsbRbzd+SqbXD7r9dGm2GF375J
RQJ8tMs0c3jgaTIboI4Y+UI6VLjNVw6XR1xqBk7mcsqhqF+56QsnYe556sKJ3yvP
UVEL7c4XWMDfA0LFTzyUYJHmRw+krfGXzZw8nw1/0oPxV9HFdXiZXAcOusJHIppK
KlY7N3G+14IyGiQ1TQeD+/AibWisuqbKd+kXsv0Ea1dMbAgflN+n7GFDomQNLLiD
RB9TICKfI3RvcZ1FAbMojSHMSXWDHbD2PIWm6vgf5Lh/NySHj1/18ZzO/2/+akh5
oqS4GFfwo9wOiFOeGU9YLvdi7+jYKO5dhPjqYJkiV7X60iDIkWcSTs26+TE1xMDB
U3NALsNY9PgsHCNB7TJKdNVStLtIx1FON19wl1m9RzEK1RFEedcVOwtDVoAzavPW
yf0jRB95c84QobMGUYix/Cp3B/r0LEdn5ZgnpQVnwc87sSS+ZoCuipQy6799/oug
ZdJu/LojjvMPdyLkIp6RGM1K+o60NTCzs/lyQkGMIDWFlgcyydRFNbLlFxEn1mO+
fCkJ8y306sNCGrIrKNbYCb4rWgh2lKjB2wMSwvlOVBs/2QUowHvGaa7ccx3pwh9S
o8e5sLmUGCAxDoSscZ11zVIi5iLfZDFx8hLISHOO2b+41+TKNSB1nxzBZUnf0kvW
rJWMCZ9DvYOFi0ei7kc5QUyejke3VpRvAo8hz34XhNK++1ir/79ov+YcFEb8v1Rk
6hDvep0uHDeAeaZTx/BRgKK0YniArbcPdEh/HcvS4CGigeKM+dMVtu5BlCRJ8n+M
k+ugJqfioMdeLAGHAluZSX6wu2STxhkObS33HWGiT3ncmCbd5k2M1Z73gDbhjLsy
+mYlsZFazcTwEtDl4xZImEFI44ThirJiR24LyYG3RBJT2XyvsZSlmn19bDmXeIH/
XBXQEIYly38BqpWi7STOYLWqDcHPnOVaL7wnVXAY3XHPZlx4k0bSDXmeybqReMuJ
RJfxg3hgfx8vf2hAKaq02008YjLKjhfE2EUxmtZ+EtW2NSWtUg0knZvMEwUZcoFY
Fx3hBpZSPoEmV7QTDS3hvkOcov8+943oKOWBXPHeVwnme9E+8u8EEmuaDzEKjOus
emXpu0BaEZizvC3WQ5AdHZQUgeQ6jhPCUN7uSa9lo5uTcU3WtF0MGK+M8rqEs9Rb
YKJ1Sw8snUaEfFubDxGu1VkXI/uDHuRBmdvmbjWiEzeSPsQqJpX/zSONU2Qp72Wd
TnfolX2pw7lCh37yBQQBZsU1w5m1B9/j6HrBxJXYIYa3tIy5iR3YW+GYBPDTUXmB
HHaxUMDqThWGkeQcNFtgYyG29mgp6i9LJvhyRLPgq6ffd0tskzgCH10HHzOntlgQ
pfCb2h5LTdkdNzNRDu8eYVZI+yqw8j8toyFt8o+KTu/3HnvxhklSXXkqKvr2jlNj
tqHMSR7AVjNnmoHibOicY/90btRYdY+jcPtYKOuYXOKSw2NuLkqj5+/StVsrv082
+e91DGpMB5ZQD5RG9kaKRNxxrht8usbh8f9MBMNwPgyfNWXE7gIjHBDNsomb6k0M
c5gIp0m9nyKl+wBXoRHTVgVdEzo8qCvtAk8R+WwWqvZ018QTsBDez+X6puiao4p2
n0ojvJRzav+Lf6NOPa9DGTiMVzKA6OJ/kt9MQ6oXuIjJJZUpLOpUdgUaGnNUreH5
oE7SXr5wJUCsoYoGPGzEaZlO4XySvqdqmQ/lkquMVd8HDtmarNBjpOAZIpTLi4A/
UHNkfBoN4PuIntHe4yi5v3K0SkzrcTm8omHJnDig0nhKM0/8gA7U1PjIt9Q/M+RY
TkSc+QbouQ8jx8BlmUflGiyZRuz0rFsBJOOMMFlIXG1LkekKj96VmUG1HDbT7ANu
Ps3eb1b7h2KUYPq5kxXxzEqg2hnorjV/OJlnjQbYW8mLXQFHZWrog4bUQKqUUluN
BfIx662/B9LZARm7QkzxjfHwwoumslzQCIX0iXZiX0zdxqbwiAjKOqSAyw35flmm
zZo0sAPstbTMqdVxssuR1JJCTOfxdFpgNtGr7uhRiUamZunqrJgTixtSOvGr0Zaw
Gdv9/1/xUmBQOr1FtcmEzret27w/81Cnws6OW317RzoTpOCDmAOmK1t3Fbws2B3v
bX5jNH6lSeRgVCa25oxirXoNZ6GxJcYfZLA17oLJvJUITjEXgxJqYCdiKo4uSIjq
XlEepUpqqZaCYB45GGkSLCc6jX1YDHEUZXATse9IFtCX3VcoCQgVToHtmyWQBc4h
L9dWFRLER3OPP2/I0YmI8MWR2tWoFRUS3Kkwa83TGp9rwo37YWoctxa/QU488F3B
dp07UWp776soajoq0eeakuvQM3TAPsh+iPuhcYH9O4CNd6VS8GsvgKXCwBjz39rL
XhxZ7WkdfdxPqugVKT3jIzPf1u8l1dzHcdCA9K3OJjjV7hrAym82A7GZx3kjPJzE
T8OicHWftWYuiV5rldqPnSoSieI+jPr/34isJpr1FZ9glyyRaxhPhSeGNXv6X7Af
oSZR/FxN8k7UV0Z6h1c8RksbwD8ldj8U4YWCDDA75gqsDEkkEDJ0V91h3ynymwls
1sZnhM7xZZc+Myl3ZdHYsPMEP1vy7y/kwJ61/o2xWdaO2/ZSuaG5ciAwNThiEWpK
1gL5aekdzTD8SiJw0Qt5ob0hBJMzSmULs7yi1amoNNEVJOOy0pYN+DXfELBmDPKU
Tr7bdDLWN04wb7MHc5PSwtLQ9Cll3/vpiGPehUHuIIfnRU3HePntDxhUZYVXUnkz
70YO/U5bB5TiVZkDasfJS47B4m3P5Ec3AgI2s9io53YWEKEmF50zvLcPcZ86K+Uj
VD3z7Cr4p9lpGjgF0iQh5bfaWGYnN6Bgo1Gn86vxBEA75C/sGHKNxyIlllyi6/3+
zMw1mAMEtsQ17nFCeuRHbvDTceyIWDGtTbYReCuV4MdX9qwv6V68MlRq9S8uhY1G
pkvZy8k5Vu5rTGTesa5Mi7nQXLZ52ufBFKYjFjoKG3iKqpoFOzJLz69efP6YpFa/
qHz0sNBoX+A71iLw7f8jZsTMgKX1qQJ+z5Hs8ouPzcCkaFjjFWiLaLE/O3NqdVb4
TIp5iFVMcoVRVOM6cPKXhriAX59Hv+rX5G3GBGFz54uzOIncflOCYqeEOj2REuu+
hyb6cEDZVz9totms4BQCq4SpnVbVOJnn9JMjd3EHYzJHvJroPa3yaiBObqvCgNuq
Nta3xFnUCP+WZALse6RpH6hkcr3d42q4+JaiXPFcWl7kFHktJlkMYsbcy54Gcjkb
igeC0DReXvIKY2OT5Avxv9U0VtKiYXmrLuRmzedB1k9KRJWKK79vkYs3dOV1PjD6
T4b7pHeoU7vJ3GOO4RpM51yfCbHppKGGvJAIyXp8UmYpj9Ax3qetC+x8GM/KkqVm
d7vMf6O+/J5Uwq9UblVaTDp30vDisR/HXxcocH8IC5KUZrkehGsjhdtnvztF6PSO
xI95Y2zSLwRJkOzE0qsB8ZNEzmZFViPWujccdedEFzTzGirXSM931IagNM7o/xkJ
IxrPA+lXgzpxVtanE1sR1mEWqjze0UgEcNi5biNKM1GSn6uIiOAHikQzgcej9U6h
1YRKqlCHkMoCQUfjCLiZkmtYm/J0W+YkMroqzT0VNZ5S7fjD3wrIMNM6qkEfgyb/
EVP5/y+cv1bzfKyZSI9909f9lcwilcFSg1a6/fAKgJYmyevv904xFB5GBM61XkjB
TIqM3dyVKMD+WYwlN3C/G8dIS/RHlFt4FJA6SpK7du2QlBrPNC0B76zxnQSCmH6g
i6u4mKWpTKvkijCx3WgU0YVUWD9Mk8+Dg0Ak25KyaO3Ek+cmhYzePXXgEQGsMCNo
YfvrF/wV+apcqFK4ySPZRaqahA86sKIt9tqmm2MxBzkkI86881TRa1OPzk63BPZk
BSL+JiPjf6E7HZFDVMkHku80NVIZ4KpuAiYQ1Kh5ZqhHo9HMtoLYMRfMHJfCU0JR
qb5LLJDPgoD7Qml9StdqEcLS2tXhm0XOj2Nn/fTkSGA3ENSryHepMu5u4cNhw+fm
HaiQu/uMrQ2VN65OetmldrIF0rd1VxwjDOFny/ed54/NAiX77ztesqzDvxIi0S/f
cEEphdvxC1KnzhWP617KUtYM/s9y8DOZ8fjcNj2/3QRXR32cpzGmle/naOyUwcMO
gn3g/335KKFlBqOZk2wBqa1w0oFmW0+LKTxXvkCYY4/VEBagk35NRx5Ypu8XdDPB
VFwnZsIXAclMc1nGtqjx/oaeyp24Y8PZVWfp0/6fRwyigMxVCgolcEtqzwkU8Ehp
nWbHnFYfYJKwtIZQmuy/Dd/dYpQfUugcRyJrIrm28PusOMwTetgvivfBJSsvCqFU
ml/S0mSZRSvMvnbtkzyKn+7vz/F03CxVgxVA2EtRheKFL6GCHUVpjupAKBY/1EJj
pDg/NZolhDMpHpSRt/B4pdSwM2nzSWC65Hp43kwba7ZTRe9RgZ1G956talfGLG/a
ilPSd9v1rfYdT5Ad0Ni+LSt+7nL1trb2OvjC+4OLcwqveC0Cdi6N3C153oGEwWgZ
vyBk4XrTf2q56VUnUUiTSbqH/HzpDQZ14k/WLpVPN+dyehDxubdRjtXEbh2N5Eax
y4DFQM5Gl8+XdiccOLQ0q5yS+vC89f9es1SHuRlpCN6UeE4xMyYXTvz8cCKPyggK
j402YqyNuk9wfONGUSg4fC8xluBdo3yd8G9unEcRTpp6j4lelZbd3UKBmxXp/15L
DpGZJpOI23TcAEy/O6AaZYoVNo+RZc5tWEhaiFctf3Et+NbC75ig0YOKYpbtFZEY
mkfpX6sY3r9aXiPb/PZ3CMmiUqgizzZQ8JgfYk1ezIz9g0ul5ANUjO7KTEhKBYen
qzgPHVh3BmkuOPUPqT9sw3Gf99tmuqHLpg2jQQFuHKOmTBv5zL7gnFBEwk4FPV4K
4KQgUv4RqsQydYYWf5JnsUm2MAycy0vrIvU7iVugG0LtybWXuNjQdFvMHTjTQCqa
OSHX0T5BQp/8dtcUXtIgsxtULVuQ7LaYBMvFwT+QXabEOyEnwxGrPkU5uUlU6Yxu
YEFkjQi48VXG8lpJkLiXErG3urB2RM2VVz7c0HqosFPC3Gl/nuZ2B+KR1tQECHYv
bZ7kZIOHcwXfkzM5fmCmuAjJ+wo93mqwam5vwhKpXLxd5kCl0mpvQeb/fAR5ZCY1
HgrHeyw+gFjSoGjKbCLQbp31NfPNQyWbG8/NoRvFw2nouxk2e8PKgMyigLcfL96F
DGUSAdi5HLt9rUgoPxaZVKEDle8smva06Gw4mu/i0Vkn2Yf4PgKYNKXX0sQAQbdt
EE3zg0df8zo8edKbV6Er12xhSCbAhSYRlstesiQjEGWLwON3Aw/0wRaNbM8z3Udb
gxWp4mBLNHxQWvGepVfEScJsAXMOb1y3aCkPCScT4ncNGNz139Vqsj9OqjwMPc/E
Zia+luORW6KWHiPDz0ficl/ln5vmAhgHqTBc1z/5TbcAnJsvwEql1zNpLNzUFM+t
ix7dSpzD8/4aJiLi+hXdickTAVhDumg7JEBUdkzktovfEFyv/BmrO47cu/Gg/EFx
P9MHkJf30mGz6kO1HtznHdvGGJOGl+UQVx1sr4PiZhXAGcn51DLcSaTOK4avEc91
EVeS+f+dK2LAeyP6VLx8Iw+z8tyJX8dzrQTsWKb1mt8CCeiVWTWgKRQnSvPfmafW
prxweIi8kQ3sM5jCwRKSI+9r//FGx9mV4IqiqEZbmYoGMT58LBPk7dvLvc3X3Sql
HiWh4rpst1cQksbeZ7Ir9VlW7/ut2Q81AdpmCMjB+/55ocHkPhsYvEDh/JHwT9uj
eUJJHQ0uePLGq/jJ3q16JRbpzehRayuOz5eY1dc1YDfN3ZNvYRqiePGawe2x/uI6
NN2bnLy9F25zEpbS0VC5Cw/uj/1WpNvXP2bFL0zsv84jcAIDrehzjhsh8AU/PAz3
8eXN+SaiuaWKvafm8990OTiGuVw+yBOjQ3e9FGrczvxJIyV1wYU1xP3qGKbtMw2z
BNc1bx9I45zL3A9xi5UkieYbtvGKxkzlDHoKRlMO9HTD7VFrEbfxbRaudMe27SLE
KooxO5H8pLgeHBBTWIENXN+AixsmgOIyFmI6Px90bTrcow7lyKUAwanqxDQukizC
jUxHPC2CYSHwIXJ4jEELZIc93h+nFAfiyskVLAVcvU2nV7PtPIG7q5L712WQIjlw
gQpzxBKlJclw7CgZiw7UXRITPaos8k/5r6TlNGlYPJqvUIGSvl5cNyMvlnVYvTzt
uaDLL06OBybwkpMLji83S43RZRFyNTEEvtEnDSvVv7uHW6FIkRndg5Voc1HH7Fqr
cGf1SKtVFwg3HgNhPipMyxiiIVotLdik4KHG/pWBdDqSE/kjP1z1CXjAVdd4aapa
lK+7FOzmlat19fBkf7FSbVBPV3AZAZ+oYCebSR+4u18iZKy4S36yC3VT1JSFijeO
srD9G0B9mYBP+Y8iY8UbqlOuRqK0oe4e8zEXIj1/xQ2uSrP28AmjvfjfJ64vxsdz
Pn59IcwAaZ6ANpPBZJ0wrQrSeB9YAng6arDJ3H8sVweUose7YRgk1qJTXKsBxSru
FrQorZSWPFRcR4GI+e3x8OByV22N23iRLuePI++pBECYNfrAMN5SFiafoceAOAIo
2fOk7iJF73QsOFqvbRv0x+z+YcZesLq46geH1HlHbCqKOeKE0McrCn5eSCX5FGLW
kSB7UlSVuEsvULvc2aB8GHRq9VhwJL6hxOLcmo0NjaW6e6ehA+DKMvcGS/Ob9+0E
kaeY7ANHJSKkgwIjAq6mhKV2taWsPxuOJNYCfaCCqTyiwfsU1wbuSq9GFZ/sANi1
nvaEem9c2n7IjzugyfGvrxk1DjqhRHY8Hhu7rjUkoMub9YkKNi827Jl/oakU+w7u
Yq9cAbO/nP/qA8cbaCZLMp7dcBLTnJ3Duzt58fycIYlvbX4a0jTwfqmOm5jjAs8o
8ICrwuRfcmAlc79dRgxu89pZzFKTnPrAwwYYxXTlwJBGPvadRfZ6zxF68GRnBYPP
gu2hMlojArgmw7cdaIux9d8Zv8sS7+TlUTPhrVGxdWp+o2OeyhDCWIPydwuDudsA
WCnZNcfRKD6VOt0nEe72VMc7Ky42j6ICEoKWUTyJNx9gsvQ4pCiHStZaUdmglvmf
x3uWeVkE9M1gT9OXEVilqvNQi7arBABWIKXrUED2d+Zf7cBjm5iYQnGfxfvmHHeM
vhcTbB4H+W80BwLGdCVqS8TeYQca4EIeNnT6TYt9cwXfQQtGP/8GFipq35gpG44q
h0VYCHQ03x3hdMJlaC0GHfBcIfKDdS6oVwIzC2/d1be5cgq4gX4wDbRdH9fiq6Lj
CCBumDtGYOruqxpKQPpHnJUYLxWlPmKvXgBfBKD40nyHsigHj3QldyQ466zZ1BQp
cgMCA+2gWbWH8rt9Axgz710sXy/HJEZJ6aALxl+jb8/nEfOZXe0xi96JAzkgw1ON
g/UPOw8Uk7wA/oJMl/2/y3Dx7GDnVUb+bpfeJgaWt0q52mtDB76/ydWty16OHrvA
vC/3KTWNniv59zsR3eVZS5HgTl4iKD2n4hZ3riVVge8dVtesMukLJwipJ9DcxjmP
psz3k+/pcwzAqaPK7YWct5r6ZeQMT19/nNMFIkSdr4Ax3Bc5HEB8/IXqS8hhX/sw
ZOFXYYozniCwWRJh8C9oJ86l3ccnVZRorTmyv9XdId4z1p+8Dq8fepmEdOuUgsbM
FX09fsC8RYE0NdUuReptjhYy52wZ28EbqcEjaqvZxGhn1upFdnCBQe10kW/lgh6B
h9AohRAp5UVY+kVe4GBrqKlJIhA2kTztuCwJ5PaOEwJX7pDjgYc66bUU4aTzIQWI
GT2UH/u0wCL2KFmy50ARJnPxGzChD0jGU3k5uJTBpgLATe2M2e78hLokjialiGUZ
4hoaXhYU9jBaev6ukU79n4o1LUWvfd4Y+ReZYX8wzfWRHNW2E9FxGNWVDfU+uisv
GZnfyaoiMzbcdwbFSc8QuBIYgBYRSEjijQ1oBZUNZrxESU/lz/ow7HKQRFWPKXDf
aBhmvrxjNP94xjVphlBso/jn82ezME/jB7mBvKIhdza8DE9sYIJDgBNd9uhvc5Se
nmOSZiE1GrMYjrFWWxH5itiPbnNou7PiwJU0+em552nzLmy+JYQ5m7P1V4d4CX00
4rt6E0GB0fq6ShwHYfLnabWdBPT3bDRwORs3ex/T8jiS1KbPNA4HBt4y/Zsmt7E7
Dv5aTIRsb+Vlflb7ePsSAifNVTNH8yVM3oip7bC8EhFUCWMbr3kgg1MZFoLf7Eu3
iSAYYr6DpFZAzmoOQnxqY5VUTGBSLqESJGZCnPWaPC4p3CLTAQu0jDAZFlyVpvAy
Wa0I2VPRvjzqqAOF9JVL7aoAiep4Gc7mdo/tfMbvWd9pA2qOFn1kfMQvueFo7LL/
v/cD9qPzcIYkhFtrRwBynB/Hpmg5gexpfC9IcTpx2veLsZRf44YrABJNeQg/f5WN
Ju8Jzk8m0lLj5eQc6WzLiCV1XsqD4nIoJVaHHiK1FupC1uULrZPx7DO4Lm11up+E
615Rd33rVwrYll5tNT8JInuIC2pEc2IS0mqPQRQcJLBcj6OPGF9KxlB/k/PtVhO5
RlJvZOC9bodDTFF7MDja5Xfww1a8m+eGcPZvQZTPkev25Di0JRj/6zNPwicWXf5g
9Zg8pUfIZGvROap7NULNxdFrHpMZ1QlOVr8XmPDDtGgceyE+39BZKS2J9ujxxtNS
zNwZspKliNSF/t8+OrHcQUG0KReOeNH8/E63gouV1yRuEFpYrdqCWU3mW7SEt8M7
dZ2FYaKivPGtk0aAw1BQN2be93Dl0PPCu2t+u834T0xhsTsgGiAbw061xG8Hi1GP
JxADjKTZuyxMlxShMQ+odFJuMpSerk709zp+0XY9W1nTVGvB7zumLTcMavr0ojEm
qfy3TasWWwhgufjO967fZlIq+dbmVBPyIrQWRqTtsI/YMF+Vl30oRVBhJdhXF3YV
GR5ZJHSI3P6if4dkXBaQZLHz2XOuLGII6wN5/40OASuYu0wGO1KgLbgp1/lSf6kH
9rqr0eemynAlXMnkuq5gSPnbSQdZ0GcFi29S7T/qW88MHjCbDy4Z4BDzUh+CPTLu
gGK5iVxIkOwcduFhvRazKfOzN6SPUpdXWy9tSjtdanUthDPFUhvx/C/mxZP3BMm9
cr7j1tz2JbfyHQIwpC8VNnr9ljhgWGStN8sys6RB0C4apEwnfeDJG10/NpJ50BsY
iI/Q4NKL0CfF7+QHkc0dod9r1mD1fCTxHnpUaM8dhNhX3MjsO2DGToVjKarPncqB
q41DDe2DNjjWLiSnA6dRlF9+QQKrslCm3g0sOcdAfGEmYUfzNbdsgvO2SBhQOiVe
q+pgWckM5reV6qAOjlkYh18y3hft+40Qh9ABBielr/Ib8RRpM0ErDGuLiQDuxDSq
4CImi3bMBHnXWHQD372352ZMtSR5iiif1x1UnjqF9tCwRJZZmfQaHH77zXQZt+8a
wWaBn9ctVQqqLZGdl4IiRHbcZ08DoKuntADh/FdLt762t7Yc7AahTAA5l6lZDUnA
ZjsA4B9AmjVva/CX4TMmvlwpdf2kOYqmLLc8Oy3VXfJcO1cJOBmAeyGarR/eNaQN
ig+Sdy/foMxZfJArsN4dmOpCl8GQqONI55Xt0W3dT8ArP5USKztCG2ed1IKR087D
/VdoPc2taZ0aKczbe13/J04kLUBQCJw2AyfEHgiFu/13lkdbau8DYFcqNiiTNnaG
Bpk5662lK0XMWTBVrZKCWDtgJNYBo8dFwLTDlj4wDBt+w4jM08LmjlerrdGXEihV
7JkFE188eiA8ESHEvrelQZPrGLBrbzjv+irXUtBrvQMIK3NLu0N1W6TeWlelx145
UgjPDasfSOuFAwon8ne2F3MBeZT4fAyenVXfr/B0UkRTjZEzZ/v8o8xQngbM/3nb
kCPnf+lAfZjpMRuTGVU1/YDsi7K4qsGqBiCRBGCNQuGFZlK43t3rB4Mlh0Y7b1Ra
y9cDeu+s8zBIRYBhthtQgI//bm+gqx1lYT3KeiGlrDXBgqu5nFT+onpql9fQtPla
rkU83Z2pmsLmgR/vgGu2F3wpw9wqqFddurPbAjLNN3mPh2XNpqmLykUpfZQCAXZn
ow1HSfUlRmAgrXhL8VSAc6kvl0zgf0hNMqsN+AAJFHns1tF0s3m8Mr5XkYL7fDlW
uiyM75zD5y2W5tEaOqMnu0qkbtgH3X032QJrVA8M/q5TqCZANq9CDBW6eHg4PETg
8sQP8p7+dUgbJKRRv/smVBGLv1L2uj1DJo8cQeTncHwjb0QsWe8hIHwRhOkm67EK
bQhxtQ/3AGaTnGiNxtDq5c76VRGD6WSFe4LsIJ5trXATlBcawNLqeDaGjBt4arsZ
ANCSLG8iQpD7ZBC7w8F+YF/SNjccw65qUiaQX/2iRTkTsx7Uz/EyAcJoDZIYhTTS
DrfgIsvmXlscCzLRwDzivhdzGQwwb0FFyiJdgkbcyi0E1fzZolJHBqqec5X8qm/S
sFsnTQ9iUbYHUnuvVCR55vO3ewJki7AiUDw0rx+jR439LufGym5WT+NhlLdO0C1j
C3vCC7vREOSE5k4rEbbCz1R8uEAlP6g6G25RX1t3dl3Y5lPqvVOtqpHYnaHiHD6W
doRlZpdnjRNCVjW9GafKX+qPhC+CWgqmkYB79jrvlfeXqxkNP/QS5rKdAcKTkxzP
c1Jr031LwbsD8bP7aUxMsJl1xUKRn91pKrbivUsfGjiPf7Z19SvXKUxcHEScGXNW
KSIzDxx69LkeHc5vJJCk3++fHpiilh2Rup7Kw+kF1KEkJy6qLMXfEhfrvBBxrLTe
02bAG5ix4IcR8suEE6XfWFFhMXSjOChc8IJYdGkHLpLPpe/dRh1hOhl5geZgUMUK
R1nTG34xT/aIZrBe/Ox2+5GG6Zl/7uS1T0tQn1vONXxgCI3N7QUY5rWE3t6kRQw5
tqbZG/ePjMn/F3NHlhGEXS9i3wXTbaHNtwrqrDotS6nZq6HzimNVw82+qrlPJZT1
zsknifwQfY2NgBpj12tM6ZSGOM0EZotf2UaVlrhq/aUqi2+5fYWc7DH75aU6cAkc
3YgDOLQHNWghvnD8aHTueSAjGJSGHdUOCZgEriWPx8aoSsmSkBh9O9B4EQnd6hcL
d6W/cJfAyuqc0tBWdAyeq1b+gDn9aFSBjakBu48DddcyuX6DXnEaTysPpZoxuB9T
GUJSZkRV0NzONn4qdBY7mkRmj4FTL/+zlIAzp50nTzNg9JvXtt7QKBu6/S6csBpS
b6PSg2plYhseLlOCv6CWFTrtzhpc3eEQavAX6O7qmvPhNXOI7SnSK9uzgyOOQYmd
yNC0fd8v2/s1SiA1z+wS3k/unPtyFqCjfT7JgFT+1u2ocsFM7ViK519Ty+8jkkl6
guTnKcHNNaRaMIqbSgXySImHSIF60yg321hGboaIhxD/yrCJpTnAfWS7zUrR7MvS
NGXuwfV4nQO3goxxUwyMzoAFLllh9d+DzU58aOhJF8Ih7n4HUcOiU2KcXsoAjZCN
B3FTOJeItdPp1D8S6rZArUuZrQzZxCoUByyHhxApY2o/9Mlqyw9X2WapViGMIVnd
6sETajxrmCIoJpEE0V4dpKE+37+Wt04e9fJeWKIP49RrL0/5gDbUDLu9jsnJ+RlB
3oWkEsFyfjaWulmX0XF4pUyNL6wamrPVfu9gGiw8im83SRoLIeiapgmP3XAFZOzX
HUigAchqDDDFeVI2iOaRpB+RearwUbAu0nNolmrqYorqWGL8yRi+shmiyPMEnwLi
S1dlAIe5lCD1l/Xom0+RtdsT8kf749Tgi2/qEq6Y1zGHNFm5R7ZE+t+FCTZzjxgz
6RP7a9coCDvH5uPSoWwCROMhexW48Ow5SYy6UFw4xro4OJ2ZbLN/xUzYqg5HIVGw
E0ZjocHrV1XWmirbHFF/C2ju5KJUNJUQhuH0CyfeZ+iVZwRyXpLjs8sLb+lS1uPJ
MH2MA1FYtPscnUqtLFpZ+scyHxt6ZZ63yetLbEac6mdY5sUPuGqXu7901oFfdDIc
BJS3uH4f2nShbA7kq05CYZLRfUuRaMs+xZzIdNREs/x5J7ws5wixdRLEO5ll66+K
JVZHvZfIbDLxSFvf7VHnVR00Wrblj0cRGcTcRD6EZYcdr3A3RKdwykMCb34VvKMi
2pgAlB/vh4yZdKosTC4KJX8n7m/x85wTieAHclykRUsgYxH7fdzgepWW6hweVc1T
NF3K+zYpXnYhz5QiOK23A+ClrQBVXVXHYMUJGXGb1VdQJvhyjeDv4H9rVeIFbEaS
ZtwDUxh66zESAa8oETJ+qyLKUfLSpbh98n+pI/LGpQLKnS18ImaM7JJ4J1Iu2B7l
BDyP+wJN5gyGcqAlI4guCUFgOi32PCIi+r2tTuFL5v4EbTaUPZ/V4YY3VfdfI6WG
KDvo5HtokBTFbNxXpajaLtJF1kDUS/4khQyF/ZThEvA7hFM7m6E/lrRQ83oVI/ce
xvqSeXzc0WmhZjwjYzWJhgmTd+tFvfaVVWzuh3r9bjmaODwREKXDMJ8qPNqRn7mi
+BLRND/A0+JonpJiNcpTFY9Z22Htc4bNGF2nPFGOKn3d3cUNZkMPKHCcC0V/lmGt
U5AihTN80vdoHph4v3AYE9V8GevZci5d22UcBPsxYvdPxVY0N9ojboUsMG77uKSj
amZMvriD8NZe4mIAfl9L90tJB7RW67TY75v7EuYGznYklUTQGqCJBOKArj/c2w6J
czAnzG5SNvn/TvMiajp5OgfqwviYtyIcAxVHx3dPXp1+82xfoONwYnDhYtYM28Yr
M1hx5MHsSpvKfY18wOmNczJCY+TbS6jCGoNaTJu4lg7AwdxMhxE1fE+WdEmOFyCV
8rtaIqKET9U6I+WBt/YAII9KydcJRhsKbjsEaH1IJxgpTLtlzUWwWRpd6sZleD1u
C+TrGcZdRocrjxgtNUfczsuEN60dte8Z8sTEwAXJA1BkIe+BVAAO0/QdEgvHE1N6
dueJkQ0dOQpES4s2wIIQ8B33MHC8q4d2Q7O3s3iebwJAy1kg3YI2yVaecP8yZ0iJ
5zEfiiV1MkGLmYJ7toalHYn1gQOCG6ePfHrDgo7uVSqJKZOo9hP5YGDtHhwPsuLr
irA3Q0se0qpJWYQYEZgQyxFzBUjEnMuejP06LTrjw1/Ox7qqKhFHLVLMcfVYa8x+
zaVhsgBPJR7WRp/q6ZvUic7rtwEfleybaX1gLAPBvFN18X2jTt2yENawLng3uIjE
jitjkS+lCujcOt13GyYUtNa0jlVRfAsfG+0/1rVuwa0Bks9OnFX+NKpbCSv3VoHy
G6I78a65awqvsD6STBkjJoOI/8SqkX+C67t1+bpqmgwJ0wINfoKmsEW7L7SxsXQE
cyPAWTShrShwYKzbjpcwFshu7VTBifgf4V8Dr4apEIL7+ZY/Z92j690hPuabTBCr
IkFa2oJ3NhHeMQiI4tmK1AUm8zljnW8KLfTs1NVJzNQ6XdXfBvfaAz03NdnWoRg6
UpKsCsju0S1MoOZPyKGGOrrXrwYK7HlixoVOBtkWLlpbNMjrjA8XG87h+izg++uB
UGSjMlmY3J1a/d/barV2p/tGN68cdoTT4jMKsc4/M9A77VEmzAQqzB47ICln7kH/
umNcL8dYREcmb9pdOAL7jK0+8+xeZ7aV3KcC6/xCQ8deA/Sbw8/23kUmFdjofzgO
N/7RvFA8X4ghOwzfLUB3qASCccVdxBc6IRxxgWw3fes2VWMXZK9npegVHTspIUqn
PJ1yXso8MxD5HnNCvd3LX2q6jz8JCBP2rWvMZyisE1BS2IY2macMVKitZB6TWLju
ndTQODFbSuSJjQk/J9SHwsjiP3AeIeBvSlEOM/GxNaOVZS9Gt/MoDzFecpno0sXh
YRtBpy+QYH7NLiZ5g9DHVMMYoL7qYwRKiBE5S55YNFtWzEsqZxvzF7C2B6zubhKN
pQFyvN1K6/apSkttXhddBmO68CiaOd8AIyB5Enkjs81IQ3AmS4n0giui30EoMEbx
K3xdob1nfJjLS8CnlIf40RY2Kua2FbyQ+s/5Qep155VY6QW5jYC4j1gijLIEjWkt
tSTEGTg3FogPUGZJAkSzudbRCNuG/B3wTFURdw3o7S1AGVbni+oYIHdfcssZ5NM0
DNz3ItJODd4svkXMSF1azsNQa4FEL4V2q0kD3qqtJNw6//6bE05BIAnLk10Veb9m
7kTrtepfUX1Q+1F4g1PlZj36t5V+VTofKzLaDAk8BPPj/b/nBMeQObrWzJ1KFcvB
BOO/rnp9DdtVsnJ/1qkIta5LeZsxAqAD1vwN9D3z9Zg9yQICRHhjS4/FCPA9nJuW
rSSDdS0AVBZnaq5bJqs/9Rm5HvxgCp8biFsBX/HsCOMtbZNtcogqCZASr11twevb
ACRyBZSiak292Hi6jwsjgzNDPPp8vAqtKOl/wSQO7fsgUCC/zYjw5Va50HKGkySL
9hlK/fDvWuFzxEDi0KB3AG/ODKHnhLnDyNakDj3GDwQeovqBl5OuCj3CURtbm/p6
HKTTSInosnFn96GKWV8Cxbnc7kSKqj4z60LHMjD6qd/Vq0oo1rl8CQkXdv+GnUef
kUWAoaSfO+ztBt6vMGO8kl/vrLgeunis15TdSGVkn89U4CJ/46JLUATHPPM04Z3p
MmZxTLQMmh0gvtbEJU4Vh9ltq5IjOh4n6EaWwSTBZo5HXiIpIr9e0Y7g2p0nkcCE
+8L5sQXrMR412NgB1sbMxKukB+Cb/+m7Bi5YoS7BypLSN1PjH7RwFfW0onYfhVxA
1tUoPWuO4mFx6zfSVhg3mJhgxgqfpOQe4XVicS9gNxehQ9kDxGGh2G62SaoxQt6G
v/gm7j1S14u47KnrIycCbIC5xbboyLWQIxI6B5hL9+E7JxbcnIDZpzl04pAHNQiX
meGahCW+/hOiPPFkn80iKjlUZ1dfVRup+FOd0VNFlGoqmd/q9rdFa2Z+0jhk5vAt
duZyfvx3YmaWP9N1jDPmOcda1lTrRbHqyBggc399JEUSg7BYNtq2kJq9rLuV0WAJ
JPJdWMB42sd66woc/Rbz1Hy6o9nXy/llEFBou7F3JT2JkA/EWxbAtkKeLFq60Qx1
Co5DpcMz7tTNblkV2gKiDR9diXci/tkYHgbnPsz9+Of48h1N7+IWk2E0DhOt2qgC
o46g9Fl/rjpgnpfs/thm4VdGdDszc6/3EgU6kYc29fU/o3eRKaV+eKzOBAOA9ZfL
hCi2/zP1dNwhvo3V/lHA80XVC8ugGt1ApJLEXYeEmR4NvqcTK+MUfkhFfTz6Xi9p
kGdVe0QBCYzek+x9BBrZqywCcFQEoWGboIDTdkd7jWKiEgEycw2tDmYZwcYfqqB4
Vljqb0DviAUMyPsN7L4HA4YBjfii1Kc3H6OCwKerCSnE6F0l9VNupVZ/aiLc5aPa
TLxTMtcpE9O0bJucViV13qt7iKPmvWol+oS2dGQRYMPWOHC/v7hC7sh99Ij9IIn6
65J83GQ9yJHeFFHPq5zHDEzE2nXxz0aaZ5vSDOgSyc5Ht96NrEO9qHE42jjw/qyx
nm447WEwX6/GmfCFIwRRF96pToty7jrV2wzjih6ADgeiX+CiQjxnNcYr7pbpXZrC
LQLGaSxakFYRW2LGu1xRY158xtsa+eaKT8Iq0c3nuAIvN2kAHfnBX5tvMULfyawg
cFV4yxbuWImGTIlhnOgBETvr6vXDsRBclPOgMf7WIYN6mQsjjhx20azPOZFh7/t3
BRk/aWmaJdzW8APa5RA3WNUhovucrCskAVkU6zHtfnrUzkupu6USITDU88jH26UD
Qk50hCPYZcQTOI5D5d0fLRNIRcUXNiIYQ3igE6501/AgrUEyhmGauGzDCOqjZx8j
XVr14z3IFF2loLGUSyJ/rxyOSbvUw5pA2f1verUkVMrocl+sykFtMArnaX+uvdCT
KBzdNno5bORrC6kYA+Q8SIaeNdZLdLaBF+Dxi6ZZxJlK+FNEnIn+0bCY4HQxvL8Z
zxalR5GqUgF4bNGIi4iw4Sk9/FVennWElO+Z31vj4oBbdDBy7mIslGdy315oBA/i
d7vRoH1n4itf3dtWViftrEof0HQdcka6kuGWnUzPpnjAS2J9/L+9MJ8R4XkZikjB
DC5sJqa5qDRCvHbl81vaDAX5GiAHdB3ximgfYzwE5qkWmnPgjZT20HAdc2KpG0E0
A0ebWrIMOyKrc4xRXIEIA/0+Obh6UhvL4VhBoUA8tw7w/JuYCk2Wxhygkgqu1MSh
wnyTHSIIOJ2AItzJ5AeyFkGSn9feSpQMUFwxHzoLPjuExAyOM4BEslWVWveiJPEO
BUuhHlR/GB41zHE6Y2ApQ5HZqo4xfgGwKHf1fpb61kbdE3jSCBpT61+zhSN5fKe5
wTq3p8YZ+0vqTSau8Ac4pGCrGdXdds8ziqses7wXbylnlTtwlMLzoYoGCsCSCBAZ
D+sNZZcUk5MlMFxNhLqK5wg+aAloAFyztMPhcnfB9gV2VvY5VvMi18StaPk5FpiK
YMT4m3UAlhFsBgdXL78A8/mkYHBi5T7q8ZZsskZA0kICuY+ptBQ8qloXlQVLg9B+
kfu9P7AVhew5erkM/st9+wlbaz4m2AwpP3XvTE12y+Xz4N9gNgXWYPvS7nhvYwRc
1MB2epxtKm/K7b72ZloTdl4p45BqDqN1ax0auPzxkfYVjtnIa1Uz2euX/GLlr3Na
3/DzRr8L7GDAI2LSUgrtUhTRLPhCH/pjwmcFkDeoBVA/3gYw55oeyqDau49ZHKFK
N4xMyl+C+dxArhyMXZSoqJV5oL2J7WyaI+aaSOGloQLdsHpf2PULqAsTuVHoT+dG
uNNlAtxfduWGV/g4gVqgGVbI1X/L609q5+sNMhTKwsxmjvwtCucH7Eda4DCHRNi5
PQRYqkWdk766zj1VnvXdGsP2B0T5w+pza5No6fRpd2KKpdjyjFlwCd3bvesVgWoe
sQs+EcGm6fDCf1VlqwvTtMdHCnnTFMP7N1vr3J/Iq+i4yBBmyDcdr6TDSn/10EMA
ANlzc/jRvXcH9IJ8z7d75Ga68UM2aGzaLmvxHtpb9mwbZ9qyABSCP6ahwRvDQuq1
g0u53HUGuG5Elj8Ctaq+PMiJBvu84XWyG7T+1LF12hOETdOH2eq5CbZs5t6/pdEh
WrvzgrDWJTqlH+w17b6gyta6KRwgCJcgpCCso0YvaA1pACsYwalY2v5k/hD1dexz
NwziCddsmk9SOl57funioAbuLlUDtmAfcSoI80+BjAGQ1A+HH+0Qvl4GSleoz50g
bsKnrFSGTiEONOYJQp0gPCAbO+XMRD+Ch1VhJqpNh8VRwNV80VmWz2bNT2TWZ761
n79/NV2Sbpi25GCf71eoJdfFISOueOurcUDOhkD4te1QwaIvsYgFnZ6LeT2Qdg7I
nQ3Nxv/fogUViDV37t/Yfbvaqi3HIV79Hix8iTnKANJDlWV+islaIgAh7KDCgE7x
N7nTn5JxaFW6U8kG7quc3ETYDKPsUTr+HxHGfTdzWS9jbqBMvdXsG/RdoRpnJewg
NFU41PwWewa7QZZ3tE9snoRCeeExOJqxi+0J+dvS20HnsqQKVcZM4S1O68UqYlnp
fG7yc+8kQN8gkH5X9pYK6ldSV+dcghqo3TMxMET6b/P6H1PBpLxOrpPJFYorJ0yn
RnISnCUtVPnHrb/ibZYbFv2KqWSv8+lztGczIDQicQSpGrs22MF8bnat68x2eCz3
vfLUgsbZijaLY3hFJjrSTD1eiOmQ3TtWWOkYuN5W1MRnIwYACPJgW5xMPjUn0kNV
74pkLlwI4srBKVGGbTdvPpubI4N3J5/f3DkynUayCObuEhSNQGLMG91rIJftrs4N
w6dB+xML0xqYBdulNRpoWqrLTeOXp60kI2woT834QpoLO/pw3Cn1vAjPfzpOG3Fg
7SImpYh52xxPg1ASzmovxuAqV2FYnH9P41sjjjZtcGS7pDET/B7lDAfA5iDMP3b7
LOLlF5I3BPi1A46p5Eh4JsumhXuakzWdpbpISL5ybbB2QTSfyHt/qTjk0leFWqB/
4/7yikj51s358iKjdJeENm4B8+Yx+0vIWoDUwVz5PLhZna7Bxa1KRsT+Y9EYVfM2
QH9E5THqhWVsWii8xrP3qUKJVKjlrv2S110/iXh9+lt132L0Ck9jByDBk5b7y2jp
Xvc1lJxEizpZvC4mFGOEZWhp7wnFY7AG271XB5d3DY64b1kJn35wv0JH9oZrSlja
/WQIHUzXNEM/Gx5Ox/6q0ZYRIpimmGmHr81jK9lp034RZOin7uqO+CA4PYAyHlbf
CWAnY/Cr/Od6YIVKUPKRL/m49ZcL+Zj4bA9jFQKI02omEqIV8Gl9G5LfdDu1ycLl
U4QjJBWbqIgfiCpV0JmRSEI9ymHQumWLQbUDQpR3S21V41o5hMrretJz9LCEcLOQ
ZVolI8zJr6Pi6VF0EHk6vgW90xrjdVKLZBP6XoFUltBZ1euW0NLAgasPGrxo+I/v
NbJKaYp/ygDGv8b+Uwq5QsgYaf8a5lKyAc2jhrxGTMYmv5TvrqPJApNXAFbfHZY1
n3+uH94iiCVonAlE9qBzAq1E8Z0haY1fOs+ILPzFAIBYAyTePZmbwchsZNh9uMUa
DxlEv39agh8UxornlD53wEeoHFzc1Ir3U6iL7T+wZVt1jmlMUghxSQPDmMnjfMkY
dgOLfWXwGCd/4Ny8t86ndTvFIohBNAYCnxGaUPBWdQj90U5wj3FihuXupXex3SmN
MwLCdeOHCKiy7umx2YPHzg+LuITCdBxJd2r5PYLekv9W5oaQmVZyKnm60empwVDk
528i8+zzL1RBgovrRTdYVJy1JRTk58qNOEmSlFGChxPMLEwgI8xfxrlaaROPc6f4
B6E5knO2K3sarWvKflBGxcid08tYtI6kt6VFa7QoKgCK1zSYsj+SjeVToV56UgnR
zGGy5PjDjjI1dPmpLB5rM6YbelU9zfkh0q8rcGquVPBr3Hk+LTh8AbJ85l0NQnns
CpX/9S1DsoPhneaJ2TiU9xhhYTR5eSB7Ir51S8FhVmkQiqbtkDLuyorRa6dvLTzb
KOQ85OHFrluWqyoV8Ypg2oS2/VhzwU51+sZSfFWOzbkKUHuw6T7XSngaJATZxJIp
Sdh7hLxv8sdVjhI8C7yyGfY20HgX/krmx3eddj6fWXN5gPKXoGtd/pY1KuwGHEeo
QDv3RYM1mWBtwiDigdwwpEwrTFpxM+3WYJ+s65WPTAqF/dmHclB93qGbYHLftuSx
gC0CAmVkkDY4N/KxAKnNJmYXWwz1POVJs6vO7G2WOtdSY2CGuAYHg5YIinBgIVYK
xUf8a65ovpx3avfjML/BZCG6mwa5rm4P5edw+hW4IDmWhMvR0QzyJE512TxuOblv
SdpAMYwtju6s6vx36UELZNiS3rzw6CcpV/2eIRWW+WMIE1bwEqrsw16c9pykSS7D
t/p2+pm7+dA5zfZgGov+VBjqhvn9btJlkYcy6iwJedlg2pFtD8edV7DYp2RkvyJ1
+tnLDbW5EUzBvTfcX8+xoKQbRMBATOuthlbbcvc1gkS0Nq2C3ZKzw4N8NG7oe+o6
lVB1D97OuUyPjnJOIEdeBC1UI8fi632S/1K66c2E83CB7IlOjde+hSELS1PpBGd+
mE5vVmDdXz3qqFyLWtEDOtfhRZ13FmW7MZMFLcDNs0FuNcR6pnNQw7puVzATFD5a
ESBbScrGRvXeHpFP0BI8kfQEaec0/HgzqMz7cgD8fQuUDdxtzTspUelN10HMz/WA
fGv2iMplzLAKPgVtfKJvehrPaZHkXZemLrN+fLTvkotN0ioPBgu0Pcbp3K0cexxv
zroB6SwHvFkR6uOpQTFfTPYOIc7t6Jv7DTzxuaLBYmSAEGkWVqIaEhOGUrgI6Kg6
mVzmRxt4BbEvzHbLUuvq0fA+hgY+kO0EzrgPbp2YCeBO1j9GGTk7AIMZEkGgbbaZ
upsuBnWLOuS9+iEMsDfvTINtPCqJtteN1xEMSEzSztAn423R8KEdQir5fKEI+V+F
z+8yPMj/bTGvQt5Mf5/KluOWwr6q5XfIMBQitFLeYCubE7HSfwKK5MSCF9owIGBl
U72bGwUDDmphwYZHV6xmKvu395C35oOt3RJorvTWWyBX9JialgnacRw40sgqwaYT
CXytYV/T/Cu7Bhtsave9LvpSqP/YwIRByHWt+2677pVUVoQRVYLomslyksbqf+Gr
KjppK+2YAjeBlA4wbkFdLQKWY62imcPpL4gTAtzmasWGsoj04NSKOGu1N6LDjmQw
7shlJCx+wa2SwbVkQl5y8yZF04DpClZJ6sZD9f7CmARCz7r5HfFZU4Ib2UDZkhfE
tZTfJS/wcgnYLNe/cj3MHuAH0c0offG4fHEAJT4TGe7g5zBZxBZB1eH6Y3xvTU7B
7txOGTzK2jZlIrygBOXYeAS+01XMO9OHZf+nWNQIfERsyfGJbGZRBa6niVTGhaa4
k2yiv3c6y4AX7/9sbO8IPQhRPLNiW/8IE30z4ggNRq2TYIDjx10kQ17YObDlSB1e
U8lVKwXdZe9TuTcmPkMdlIV7M2hiqaPcuS+qcOJMbSso2WRKGLratCoQskXeIwWd
CoANKyKzqRiFqWrHhry6gKrPUP3+95nrNvGvn3OpD/Er+Px0J/OGVDrhjofIBxtE
Mv/mZ14ZK5e3d1lto+ACcYuHhUZhJs3sApd19aNozjk2mpvi3JHmBPz2hWdqTOgM
wt58ilY8B19oXMT9CE6dghqMIySvrSMerxnGmxJvMnsSrUtSmHCKFo/pmV34yyw9
keudlSzuU0Ebs1OO1hI4bFGqkKgM2zivR4x/YtiG0WRrm01DUTXq0g3YDg2ttWbd
UPWw+VxkGKC7bbJw9yGqxv/z+uG7sf3ZTY+EAbazhgNwrniIf02kQwW/PRu+I+hM
+N/qiFXYtvyk2R6jJrxMzMHKutbxuc50sovVa0LbIXANnRxg/fPMxPtgjnmlRvcc
BEqpXXEAJHwEh+x4N3staG/62YKmnhJWChvaebsnmliqOq+0JA7ZpeVc1rZpuAD5
N8oHi4dZXjSAUT+cfKlCVJcF5g0Xzd5KfUKPpmzyOyXQU8irO0x66jarxZSGYQdY
4H02WKemWR70BDfxGYSWTk/EJyuWHoGfGCbdcuUbQ77QLikhdI3U3A6VdqeYRsq+
nVaaBvlxg/YA/8pGoE56X1kRE5YudCF7ZJPi1B0Zm5o6bK5ts5Y0VY6QKPV98U/S
1HXmJ17NcMXskE73oD6uKUenQt+X/3O76lRgl/R9PMERHKJmjazkaGWeyRK228ao
uFVoVLv4SY+AWLVCxL0H/qGMxU9pEwjp+KcNoYW3uhQo0KLdBmZ2/n2v9B38wH1g
bLjRYEMmC3zU5WAsGySz1PVWqQMd2HzHu+jWMYpxpNsAo9SDzloEmJO4MXoZqg75
oC7D+rXAj8ETgzr146zNI0qC96SeZbzUDKD5Yy+ANEfIgei/W8jdgWtPqHzgwogW
VrZQF3Ydxv2rioKI+caPUuoom72wBQuRp5h/8ujF6WcKQkq5dNt1+AKvq9FZ8zUJ
MAJ9kx9rOcTNGhDWYPGoYD4KPOO3JXbNSB2cW1SeTDZwi0TH934TllSgD/tfM24w
Yl50pkX7fyAcWXeOXob5G5LdpbPAH3rVdoLDx2ntfUIJEFuVCk8T7mnk5kIkwq1f
rLMwRJNUByaX8x6XEOstPqc/B1Dcfo2x/u5RJ18MZK5eiePDxzghgfp2FBodp7HH
sA/03Mwr095SdBD3RjQ4MfUr0KBqZayxuWKhUdUVDJOKpZtphIRV94Mk84t5BMFY
cYwuy0nqepwc0zZTzPv5LFmZIQsPA7M9CcMCrhB6auC/9b2QeDssFzqM4KY3rAbE
LuvOQ61/VSIOrhuqf7FnoQCKAq1mRaVNGdnUMV6A+CbbPdasFMxvDE5WtkwEggBX
VUaFMWtWl4p/fpuRJULWde5dXroVLiFQ9hh1tKZ7jmPOBlVjAh495vCMcXg4EujL
IPgQgsmtJslp3Y9Lx10LT4tcU5r800a8k57Y/OiWJR5WT1y3ur6k7ZVwPt55p8a/
RdeigQ+eg+ZQEHIGPnkSrsTlHWnubIaMvuqLLKna9RSvweY2F0dyFpPzbzueKsR8
6fSvu+H3L0nv+MT8PwHKm3FJdDW5NCZQ5KAsY72jPjQvc+dqUBOQtIYmBcZqe3MU
RUX/rEfJSeSRV6w0VpTdcDcCIBKY8J5inU1BJ+Euy/yYMQVawihwX29T/xWxiiTT
2CML723ax9NTlKFzjmfh740AAI2ZLskvV37zqKWj1JqkZMbyIYHFgGawQC45Pd/Z
VAGcMSXBZJT8uIX+4YBCMX+jc6M0/+FIN/jS3cjiPLgruLshTbhklfFaq05LtfuI
bgE6QQvxKxJvjNoCbeLQMMtoP9/ao3AtvpcfeX/P61CLOJ9jKYl4s6od2tNpGzM/
vicTzc0AzPRQPerystKyqo+39Aam8YZ6Etb1t+vpb+QVi5yOx2xAAx40cGzjGMWG
Cjx+OkUXECFstsD0iBKzoeikkb6/LfjA2HVVKwhYDQ6KLeQCCD2BetCEj1ZS5+3Y
JudkmJoup0x3VDS0dv6vylo7HRfzOGtRpcrY4VJYimKC6P+4GwTosbVzRo5u0ql0
AiB9+iVAeGP9iLQyDf59iNEYfR6PTgRamKZA2pBUPBSI/TaP5hErWaVJleUGKV2H
r4rnQolT+HEGpG3Mj8mrHdWCIVIdkW8NwDqTwCUswSeLZOzChPtF6ZqETGGmA7wO
U6PgB8SU3lJMA/2vBfqNBx0ChPR5QCiJXl93Alian9moKNznLEmtHWY+3duGGe14
RgXP9pOplkeivRPQrkLIErAg4EVXsxJgzV6RZxOMnhf37Hrv0kAxaHtyPgjMxaDZ
jk3A8mez4hYmZv0+K9ol48GdbBwJyfl5NcwmQxEUGNY8zJkmMkBDPXJtOYHTF649
s58daVkIPKWGKjP4MUXk/HoHJowiuypvtzXyNBs1tCzZJpH2YPsPljxTd42HW5c3
7hUt8FFr8Z+6URkNFzqtPOY6nxXNGxAU7x6vUu/EcECvicMTpRAeV9SlFbEpNOyW
mjKuqoAaBaTE09tR/DEjnWBq1mXwzsf6PGKx+hQP8lU9bP3KRJsd+d5TDKSqNmAA
jwAHOSMk0GQTqsDxu1efR0QWIfV8ZW2lw5Hg3320qSD2GkXKPXX0AOSh1+RAxYnh
g+5oozwdFnw/f0ze99tJYpgT7pApgOZAgE9OSBrccHZlcz5IS1kkVf3YnKglje5X
BQudkg7ThKTeDY5n77uxWUeqXoDDt4M4kEP/Ps5Vm7GvCPjGDvHy4PWz/RCLyfg6
YLnz7Nq+OL3Yk1F6b+ZXkhzFqtNEMVVQoyi+uUNjtToMoFI3EmCEwYpAdP+2SY8/
XtrPARZP/wgPKKg+L9QqRsstLeHl3ZbxCt8MEBaRmy1yZv84SZw6qwcSx2Ck7MHA
5s3prCxfx1LwQAzHX3aiVa/NugNUdQh2RiHzKFEooGOt7CnwNZly4YGFe3XBDdQ9
ZX38SxLdch/x7kyczaFLYPeLnGl9RBj0Qg3SoTrY8vULNao+qdJOA5Q/8W1A+tyr
HOsaLYjcsFxetT9Y+eyTlMjUbOhkFqI23ZfxiZF9UX4fXnrqdrRtVYuToQbkG5wn
7W37bpSFvvLhNA1ysNfspyi7Zdss28mEiEHtA2z5sEt3wfxLE2jotiPLn+JX73Xt
26+q7GSdicM5CRkZYqfbPTnQYgpEwa/NbkQHIJUyyIf8W4Hmy21IzPHK420I5PBU
mzRhGJh2UZnfb5zIlSBCmlLDjPYncBvzZUTcNxvCAPqHRre2lNQxN5XvDJxg/9Aa
Pw/GBl1eV9Wiva/0Ys9uVVrJ6lQpff4VxGaAhj23K8zEpmhNO878FozVyJxXnpFG
BgXN142zK/vn7lZxEh7uC5n7sCw/baAtjkenErW0OYb2nTraBBtt83H+CStDOaBG
eubbT2fYpZFQ1DL8AzfN+dPy8Pn8RH7mg8B8Y9WCCjsGcz3ewIVjFFwCRebNJme8
/7L7MMGVyt5KZJwlbqY0kwIs13yjr5XHPWGzOj8k4ttKETOLpNJlw5z4e0psrnj5
Zj2Fnd0SeNs4VHNM+cX7QbKKTRS1WQh36MhpvrBb7AOBqiIxYJHJEp6JwAzZo9dq
KAli7o/ru862Y+eO0bCE8ayxaqrOioCRUDy0wh1rb1P6EXdgzKqpWNFYWB5bat0H
3RBbvmkYtXpTXxQCQ/M3/+qwBXkGQhwpIClNlKxmHGlsHN3Om5q/UonNChUq5t/Q
bpWQm0E+SsaVW2/zj9HkEnOV+Ga0ckp6VbmTwqnDr7MPNpyg+EqUmi2ywyBOkrh+
ueg46T6S776/CMkQxqqk9aVlYC/HIKw81Bto1F2tCZZG8PTo5aXYnCZtPJzzjDGL
IOJWaSRsIE7SvexnaDSl9udaipBRfNJ5/N6MD1SwFjrbwdFE7flXPWsMV8hkbW+C
j9F/IkVgZllCQfkkN5GQBQQ9QvvfI2WGani1PMP++W5W4rnAMxBt7OXoulOhk27m
zsUGjw28WG0Dg5Iqm3xBhuttFBruMUJKQfkUzWbOkOGB5L+hqjqkN9kI+kC550gB
IfH14vhbuhIzwu+nkLrWkMUZvLJucI/4c+q8e1fyWVnq+YlMSqWPFdZ7g5rQWs1f
+LXpuDrNcYEF8tB33Pqb26DR6bhplseuJ/yvkeft3wN3NNCb1FPDvdvuQ2AGuBXe
07QrsGcaZ8f28X5vdGcVpItpecFCBelf1fyUwaTGET3/QbSKY7Uacb8xWHE8NT7T
QyvhH2LTfaWrZz+HAhNwBvK3/qbxFnuOdJrEhV5cz/7sZgmwDsoiVc2BouwsA+6P
J4h8YHyJnW0ZyRUc2ss0WTG4ON2b9pBTZnbyr948GKdYvHCR3HkB1Sp5r09AyBJw
AH7+zroUwIEtFFKuvDOaE0jCJPpz21KFzfjUDlyV+truVkSzvZiQmCWxSfcrTW7T
rlaB/rPiswP+EjfVf8+bXg0ugYRQnphVClW5DoI4jgdfTRRfCKQX03KhnAM7Rm94
cEIFeOini2fPUcfynSAylhO3LrQPK1yGcevWdmZrUSLS45VkmGLE+HVOnNeFoXOq
Y1ZwBDLLRhLKA1t/i8OEa/lyw/QhoQkkviAHkHj4u7T5aavmuavWbAirfalB/Shg
+YGXz3ODL6wNSnoPpOZNs/niHux/k4OKyyLOhbQbNBEFkee7FVVGsNTmIX8RRDSZ
psQkUB40K7rxsswdhFfkwZtSntEJNqvoQt74bQTCbfB9vXXN0YxXaJUGSlSWeS0U
OOlT8g/lRp4xEeZgK7m+3wUDT/Ce1I9KPb9gtnxPCVdvmq5ncs7gidgdatpwoL9H
1Xu9Xy9EE1kvPnsQ0oCi0I3MPITretRh37LJy+cR8VbC02HSzGGQf/i2oYv6VNcd
AqF0XfHvingb48ko23r2G9JLVC7UQ5xTVg9QGCw6P3zip6nC8K5G7NGfMuNwt0V1
tMaXsPszh4QGSUXHrwdKKckii6Jn7Nk2X1u5TTIPzReuFHE0N+KsmJr0HoNvhinj
4OJRtlO2O9DH+4qgS4hIkwO5u2aa5np9zt+KOfMxg0tj9BQtdr5e2hyETEXkUQNo
BjMmKYtEZlBP6BeSkyeEqigJJoynNSpP6hE1KVrfO6yTiO3+9oU63Dmz1b7oRlTw
/6vOgj8xrhPB0N/lpSyG/KSrZ9qS2z1uvuoTr2PKLwTLJ7FcytPszIXNmCscOYK4
BcaWIq1JLYItnZn7tLPzElGgwwhlmlDXxZFWYGAsag1DVjmJswGrUZ/7coka2qnc
0d80twpKgUpY+pd9R1by1Oy3UJ0V+gfN3R0OchNaXILLi1g55mg98dV45iQHXHby
VGx3bG5pk1Vngw3Y0CicH0IUHbezlODL05t+W9F9/xBrd4KHpdY+wZCcJYYfcldM
KTg/vPFhzwk3T3ssJQI6GU3LF8dYAblfZ2eyTTCOfj77Uw2cyiABwfsHp0ccmzk0
evWRstkDQiU/bqS+x4osZVJayAslTpecVMeTFcA9wNfBS+5dqO+b4cL8bh/EEhAu
4uYJ9MtstHlEYuIu6UBaHZ39zNkNOQHCSMr7PVoh8oJuwoi1IKIwvKYdAXm0Z16b
gH3Me/vE06zJDw5j+J/geUeTevOgsSbPrhY4OVUNAEUMLtjmODACVW6IR8Q4Wa/p
+tN+qB7OcQvU6P5exzsLkGr1vd2XFRog5d5JHhvIA52+83zu0kBRa6ypcbJTjNj7
gYpvHv+sCCxQesQmG83/O3aSYJRwijZe4cMheOl3IZY7JNFbnldtCtIoRKWI7ng3
FrcknYBpXPiLvPSWocOa10KYJz/V1IG6wtH6qCBmKk5mVZhMvuS7KV6v8HtOsDUy
JPnqXxJYxHOHtr5uTnCSa5Gy7Cu6Ygtx5O6QZDShiAiYVfN+5h4lZc5Q9W5XxgBH
RuuAeQI4Gv3Te1H2XYiVITwsQGdJ0C5ZjM3wu3lvVNEHMRWo78VCZW7wJeXTsFeE
hwINEfCu1HJg1u0X4Ije9dn1TXPBMI6VCo32jgwkC3mKErpg0mV6XZHc0gMcPNZC
HLfWlWm5LHRRcCFrdiAA/84vdIaZPSXkYHWTFp5ALB3FcHzCZ1VHEOxV0KBvYp7t
4oszXGeBxlmZ6D+caM0r3Rh9wOk6zPIrnyU+hv1OyBSlrMh1LKyBotD6RUp0fxrb
ZJhVNlYyZeyMTbdJuQ3Tr26NDLS355ESXG5aJRATCQN9FgS7tN7AK/Emwdqfk7Va
3YVh3KAAmtLyDFZ9bgkcupa9KojAYBfnn25aY5l+zUZBL3KK8SijtjnGZnOBSEIA
uaer9hR+eVOsNBEl60698I2DJM3RIHsYcHPf3qRMwr8lvyFSzlErFz+z1Yt35D1v
0CL2MN6m4Lbg80CoSqsUYEnvDnlZ2YUcZpIUiI0StapMtMQVu1/Y/vc+S4sis7PU
skpvgaUMkB8szJcQEe6yIv0vFuVftTlKWlXhB64gQKzq/XpqkXKNbZeAXeElzQ22
KRIhPjzN4/JmdCsRHFNSqftU/HUsEAXedGQKzgaFJHl+EadpAj2mTEZcToSCcqfX
Eexqgm67vyxQA0c5INLaBg/G1VZtgeWHAW8IGIAO6M9AueFONSBSTa7w8h509+t7
zKae10wRTac1pqx57tBX37SNBeDe5up3REJ8y1aM5HqNtae902kdOhbtuljAex6w
U6HmoH7qYJQQq3DRrYmJhPDcVeSXnIWKKozuc5KPNbG11S0YABeMOIimlmV6T1xC
229yx/HZy9rMd4C96CYB2W/Q1Iuspp1upyAAZKeEtTLH7ari8oMA7pOOLjDYIcBG
Y19IDPrFG+eLTeRV4tullm2V8dvt4E93JoO8vI0lO3OQ0b4Xel3hPfCNXXWHHNJ+
rRneV97/UFjHfFdvlz8iHxR7TjTXGUpli9XGtJy2W7hiYHxv12ITlxTl3V9R5wwb
YHSSdHTCG5PppFZzDA9uDZgnW44BEFahPccCZo2wn2JsslEiWkwo7MzkWA5jjmld
7v+SiSkGux/0SEDJpW1UC2hxGWmXW3nijXWGMxS1Iy1iBk22d49u60SLRitYFRdY
/RwImjgrVjri3FOAF4YcYQUhXvpuEu1QXNpRn0dg/6bOmqWKs8Ak3cApYWutdDnI
y8OUZWjcvGbUX/rSTI9oi1GOeeEwWBD6txwIvWiZM9BaLQf5d26wMpHFe67pra0B
IgUcCJ3ugKQJDFhbOj1pQscAjoZyDZiqaRMoewKa98e1jbBtVoy2TQkK6ZXxD38C
x9cex4m2HI08W5jTGXfE4zdsZNymQm05EmB7Ud7W3EqmhhBplJ1oPaLVuGrqGeg0
tWrhNvnodgjz3vQfT2eFv9wy5FPaVfTkRkAFxUtSQOsg+usmLsUFFYjAWKxiCSzK
rWeF0DKDvaOidLlm5Z4/rX8bN3TR84iidfT6mMbt4jAGnFHaADrAWMa5muY0HOzr
CDNQ3NW4kLRYlTlwZa93cmsSoyAOsB9eJPqpYitPMi0HJGS25w1VlxWpEZqHydkA
q/IZpsmkl+x0bEiqcQTb/S9HG/yEoXz3s1SuWKeSMDZvld4HGXKWeTxw8AJaAIQq
a5qmfRS7eU+GN40wkKlagY3aNNfZpuR2WeptIbZPbl7wZNX5iS+bsta9/L3zEapX
sppnzc4rHox1TEWH2VDvT7VoVUU0jHhToE9ukpBGWpecqsnMuwjPIm8zuMg493be
r7sD9yOSDSMnrok3Aq6vwPkaJYY5P4949ohBATg3ypXPNe/EocpZfgLM26a8AeL0
1q+oNVhMsqwmC01ShAdFmeFN1tfj7JosWc3P6Dea1aiyIXAH7qU3ytVNwd66915M
Nk2YHAqvu9NxWI3GmZz4nho3akPVvLSG/jmlwKEs7M4eCP1PNOasMa0u1dM9weos
4I+hsFYDmO3WI9Jx0wroqLzSWQUDjYux354wdgclfmx4R64BKzp4j6OtlZ9FnsPR
cQRrbUScurah/Pfh3AVMOSD4SjJNOCfvYyK4PPvc5yZk0P2xVzLmpZorgowu5oKA
9yy5vuqrTOqGb3Qz+xaXUQ8MxPB1ylFdclucC+J/fn3ujEIGNYuCRsNZvvQpz+QV
/yNnETnRr0m9LJMflPfb5wTFX4mTaZQC0lKPdXorAc63WW561JeRdcl03Ca04oOm
bDsIPLlbDI+cXI8RgGzzTn2Hu79Mw8hrUGnipYSzqWvWeVHzP+nY7QsRZwxed+Px
hgUEGPdN+1JyYSCLgGXR6+GyxA4EOc91aJDmxw/K/VjBB/LMNa6qh4HeDfSnJn+f
SMdVgo1fkcJLl4PkJjsbxYffsoFGJmBnsMk0Nk9t8Bn0A6ZyjV6XiRKKcQYWtAcT
RtkB4J9Wv5Y7te69Jm1X9TqL2og45ivAOmk2nkWi3qTBBqaNkJV9Rs0qtpR7tB53
17HskLBeF9K9OeTmBagC6DKvCngcITKyzEqVrdsYUsvNRKNWzFvN2gQO6Fk8aJzL
YGII6qfXVJMnGa53k5OWxf5YhG21Qp6oSK0C/NQUWiPPkgundFRt/mDuhS+nen8B
W0QyfUKUMsLDd+LMi4wZhvJb2P6OTvuNBmccku7vXjIr/h1RETErOTgKSU47esQI
4lHD0+Ydms9s/L1Ar/MNj0vYEacxfEptQ2ANDAg8aIOH2lwWlwPFWSA7PAMn0Rq/
Kuo+s2NXhZ93il0Ps/ILzJENHZbfOlNnmogfgczGXwO+Bjk+MBx/slK0Usb43G5H
pVRPGRC0fLyIAZDQjKq/spxs1xBGNySzGQ+cg1pp3lmMszGdJeodK6jTMUtgZoNk
B5KI7febtWdQAmW4X0Lqd8ber4IttFUz0RDtwSTSZuw2paOHY2XWgOLpb8rpFVTQ
mJwlIziYkJb/m2FsCC+fDxXrZgX7AUvKpS96kzDmmKgt1GMNi3bEewD8500HuMdV
s6lqkqRTncbugqaOq8Hb7bspqdkvsKK5ADeNPRZ1xdTmko7VZ+oBwaH7EUDymds8
xhjSfKehjDdNmtQn7/O8GVxi6fotirxCs5OE8NbNxJ381N0TVvLiVrqquUDwD/U7
PuxdddwXjBsIQYUJKIoHerhw/bLNzradg+PyUuLqYK4v1qBvMftVBTHN6+k5k6FX
Nm/xYl5ufIwfetMTo0YPOn3gBIXBJIzXlDQctxkjnAR+gwuzTL4d1+OIL6PEA4DY
Gw1FgGPAqg+1V53c22El501rrlpRfkXwlBMLYjfSFxjcxFMwRvtMGVdTuf+QvcFU
nGYEGBKRVejlNpUeZpcCQE4Jf8DlnBSgzjplU0QE1wyVQI694txBpbppSYtGxKyx
PcT6/zzay/dwz7h6io9udBBRjCtW4pFUdTCWLkfeP/NnZB9j8yVTkWxZr1ro5A7S
jVl5EdjhT+EWSxawXVYseRJG1KG7zERwctA3KRsWYPqU7OIkGHJBRxbJrzxcciUy
N2KMxp9fJdwBDiuLDhm6K0lC610DPu/fd3janORRuFcQ3CCMiIbP7IlSTMzI2iV8
GNFSXjbBxrH2k0lsvZQn9smeqQk74BxIq/JXg1PpUb3gZZ0kpdDSw/egMRPdi11K
x1O1p0bzdPh4dLXJdEK+CXGPyTtl60r0yAxa2KLRV3Cgkhal6goL2eQbwB3TAIfC
bMlXwRFqRD/nccfj7o7vJqS3ckusY/9EaInkKBcJlFURhisiByAgh3Yf1d1+p4+6
H8CybltBuuRtPaqIx2bFR4Fii6WfZBYsTXloDkWH4KdqWVmsEEe46xiNaYIYMe+P
w+0sq38W8y2bCVU02s6/Yasd0CT7gR8iBYkxgz1Jomr/lyWaTxfBXmCdDDCTPL15
2/ytsdpZscfjK4jp1U2DVmr3OOLENdyH/cTLfapG9vamC444ryBSVJ3mmAORWvqj
mRQrZ5bS+o95pXVnfaFs0HVpdPZCBhtcSQCLM8xpFr1JAPKMc2yDn52Acna/lRtp
GxriY7nigJFMigqHgcLkaz/ZkJLiFQ1mL5RL0anH+bU6iMMWr+ysrFj0mjCPayl3
IdiT717NPQUwQcJicEbQrYsdvMeSXAINVVE8cCvx94Cu5mLqv/9AEnv+mva0tYqA
HY/m+5eBygUIeFfeAkuFlFFehS0AeRMhCdA+C23XC7O3+apw30ml+PgB0TdYKGTB
KfbcBmaKD1p5ZYROw4pYUnKOFv7gNOr4mwRKIWYH1ELFP1nLyVkegFgHVLhIT51N
utxHSQ9iqaVa0gOWZEi4iHvVAS0+1zmDiMapuTANGxkmeKISxlvTqQxAry1XxBzJ
wMun7NrleWlmAFjj50mvo/qrfZglpE7Li8Ew9p5lt9qym/juG8UkpfpoIJHO7ewb
+TbJ2wMBnSiIFiWCTjWktQxGA8Aqai851LXXjkJ0+jppReZ27TYRxMAnb7WB/C02
meofcD6lf7o5Ofs3SdEEIg9nVZLxW3P/hQ+rz9x0upawhgJ2GUWb2b3twAxghdZB
3QNp8vgYZO9SNBHNamAKiVTkGvl5Ur8A2qxhmndF99Out9x7emteu0VWwYq0H0lq
Nh9HOjTdff01I0FHI+E7KqyPvMP2C/GqzW1JxDi27lB8d1AwtjMeyD2USZK1ePLj
16NU/FMSvTjw5MOQOFoijuQH3k6JcMvq4BK0zWvUV77skkpp6UMc0IkdDHHhNL63
XW3utKWRXp8xm9S4fwpTKUd/HiH5S+xeVwNjNEU8NBFcPdQMBWboN2VVgZp4l0Ip
UQDWO91hAV/EnH15iLGVStEWjtsLDsqVMj9OPef+YwM+jar2a8ZfnF18VgAZ9Gx4
Zl9bJGKkxfEOReezu5bgeItOdKwxKR+68ngDb52J0jrnX80nGmhtMcgYdAjhHjtA
TTSzkyD2Od7i9kkG6kFbyCkkavMv/yjxbUJl7IDs0Gf0L6Nxog5Wr9XM5E9/8034
gVR1dAKGXozVATmlY9P047WtB2k4nMf9RMstqkx3HUfyu5uLBqAfXlRa7e7rBaDp
X55Z0v4uXfqGcIJrjkgHwAwIb3//w7ZXnGq/Ff6vwHvv6dU5IsNSIJ44sqFOW9GA
rjT256GCzOVBmD1e8rdprzfOMVEBCC8swaYixHbNRihPRvxQQGhpaZXZGCZPwiph
RNbXZLsDUglMbmkC+xlcqhiCaz2VBCXjRlsPvs8Q6M0SI5FK3BYf7MOe6SI+Qz1d
HnWPyyJxz3AY8gl8kFwqgTNmcNcGKnDPIweYAjWBMALapRhRaYQKNHwAbLahbm9T
xgzv4dmE71bQbD5gF9Sx7RsHW/RhN+OYtZlHpI4wzs0h03BkSBOidM2dRaJbHAS+
W1EqlRw229yhq5HtsF+n7nCWFl4WkWpjHr7iE2MyxgEYvOsCew5hpSEkLChSj/UQ
sX4siTdGoSbmk9iK43n65YpeadLdo+G7W8I569LdbXpa8Vp0+TrqOPcw4VNllw0k
4LKrTg2yVKAOe5dFPelg0MySK0QqCgMw5hyv5hGKiGntg6rpbTLt9glkx9VYemWE
uSqX8gU23sMb8pVMRAX7wqEGOAP57Hvul/bBVrNRT5yY2Smw3/TTYQX1r7j0z/Rh
HQUTnrdaF7F4G69Wevk9cDZxN3f2CmAzZKvG5r3xNTK72bQLc8XeloxgYFCNEYqL
CJER8KQvvsjaIxswVU1TA4iWAHJIFEvbhFwpTJsylTwbh+BJXCNu5XG9tTXQmBEk
yK3Z7nGCo3Pa6mYlwiR15i21gnORYQDhvk0HAubdukQ68Jz6lFw415oYdGVn0MWF
T7foH2Kd2SoG96oiEy4qyY7k5xp7Ntfxp9hf+J4Fv5xmLMGx1gN7JsYdv7c1d0Tl
d8FAl9/pBrnvbs0ycwnXR72C5lFrVcntOKZRu9Kmm5Xf1ip3g6JdVvyo7NJ2gSaJ
1MxcN+SF/ImB1c8UKqXdFR2e+NP/C/wbDG1vsXz6HNy3vo/N4raMZGABPcgfufLh
FL2BTdLNynlGQwxkMAne1K0Yy+Ie2nGebS6Fbrl2SgOVG8Sq0kuL1h8tw+UgUao6
GngMyX5p558yas4Z9v6jO5IXAquoh696oMGMhWwwxmU/f3niVUeh/Vihjr+ZuidB
scsqBY2XIQ8eZLBLFQMc6HgcswCZ/iMxvpI0T+BCTJ4hv6kJRsUBZ7u8APSJECeU
O2K1Oaql4DY5h6kuB2YPQ4cqLfNP2mBUa++0ei9skqPzj4Y4tKZ1dyXeAzeUachf
W404pALpSuVQdy7WPyp1dhDIrd62lGJeF11ZXN9rt+3su6fLr7Rag2jI5KnrB1lv
fe2mPnNzrk3VdNttGkyVmObVePAJQS2qdpMbVH5MAoIUPLx46cii/1+J0SEu37kk
IwkDo5kFe8lgRa/kru/Z+7RX9f/qyB6S6fSDMCcIay5LmoIwjZt30sRhq8eL9JZJ
PBRL4VmB3TeYfL8xvGrS5S+4Yqzgl9enSM8jC4M4mCAxnvgefkCGBBqYtskivj5k
PLmWELg7VVkcH95JhNGVtGIMzib7a5EDalHmZ2wP/I84f/9Qswke0VTRUgH8KlVt
wUDDHrFOmOObNybnWRNShMLBQCpXRBt6iVcK08IRxOcgy8mWJc4ptmsqp+blDf3o
IvEIbNGLEA2Qn/OiLwdPUEMLT9zbiLrwpL5Fli87EMb12PzBJOdbbk3C8GKmWj//
JzCknI7QDCqnJtGYAMiDiVdmtor5L+XhxD0qeGKcsTW9jsf3/94wKEuMUfHmoI2g
rAGy+yTY4SEbCLSsYGpIX9Pq+chEA0xW+PQcmh5kQujcgAEFCnqwG0Zj+kdwCJd2
/Oluu6IrfrvTP67vv+BPAevylCiDpKx/V/XZbxWNRNnvxCK+w90Sfa6S8/f0eM3/
oWlFWM+rwHlnTLHOw1dCEz78ZVj09KwAYGR9C1W7pNjK8BowRgen8L9bkyxsIXJt
geYWGV2X7QyY/DLnGUpgAS2D6XURa/fPRk7WyMDEQGVqXNG3gGjUNMe5/48IqXPK
cysj1OTLWZB6bB2QLHFSVUGQAtBxrDbL8CwpDjv6mp5x9pme7RyCWWP/xcuJkxPy
0cHXl3kJBO9zNFTBp0JL75AcJT/iZ2Odh2LcdQsx97lBwmESm8WbcoQ/4z4zk4Av
duRmnGSY0Bx2pSHQHJ4hpUf646ZVCLb/0Ee+M2l25Jdgvh7vKUNvUL/MnYEmyer2
4pT7Rgmi+jYaLu7/zSyffo3LgjH6I+qbVC0gbdKNCnEOQs9gEIbUbWE7XbVur5d4
aZIWDDFSsJ2yDLG7goEbOtP2rDVWNE3b481qC9ek82ttRCpi0vOSYcWO/N3uk7Eg
m8G+V+a6fUF5fmVsOmSdxYG1oZ95Nk4fioEF9t8EJczOp4Yo4vXw4R2rUve3gOE7
Nccs/O/MxuEDl0nlKOL5B1QB5ABJeNjr5QqioW1DLOeBWtIxfSLppl2BdF8WeiJi
CGiSmHF8GQHyAbQFrP0myM/YnwqgF0tUlqGZWTORHHIQ4LHpy6eG7WaF0LB0qFkf
hGPheLWSiPY3Ls+tke0LjZ9PkE24HonWqP9VW7De+8SBgiGH3//+ifdi6Hqz8af4
tCZdsOo30f4DNoq8Z3chhGhvna09atlPFd2TIpT6mdbwuvvhWuDvJWuouHbkvu1/
YBrvKa1hLTk6tL6FNR5HgodSID6t+jKqVJ4AYXfr1Gv+537zqVE1Oeejd04ucPtb
gqNCA9cujPXXOBahPHBtfpDWk+nEVHVia/hGOHJ6OI9cYMi0GFjBMRfUy6iJYGVT
/51WUVGljcz9OaksFs2dh0XMp4xlaJpNokR3UzkcvEgBVRX/fRgAjaKx5B7jzwk+
NQD8F9IbiNLhoFXm5zbHmDcakQJJYSPrRFXipOVWT9x/Kb/zgJLqotJk8ljqk0VU
ZkkGhzGalza0/I2iOnO+0hypSB1C0v3d5SEZzjAmLGzXQTdtZGsk+cYDQy0hUnoA
TrPH7PA1Hwn0A8ganZ/zj5tKrpwOFcJKkTbiXgFF4MqcuWuIdZfHL8Zp0gQsWDUA
BVVmME1j8WGrs5jBk5tJVR8dCX9MFh7bUbLDB0XLOALwhT8B60L5hdfNCRX8ikAX
Zwrc3guN7k3UVfgc3C579XqNagDIC1dE7Y99wKg/373nU27RKElIm0ftqxKdlwKa
584/k6WIVnkcSy0dxwAf58M1TalWYgQgdU0w2dPUulZBynC5mQlEHeDF4Hu7r8Tu
LzjIi3UAbRpEhMCf4HRzmDTb/i8yTnCIxSgZ1QPoUCVMsoNDGUoSkb3hc/aQKZ+8
ukoBr1G8NvZJwCrCjGXc8oTBfe+XgAC7x1dl7d9ZrWzt9AypHXI4mmKTbux10gsk
DRYBQeY4LFgPY6ZK3I/PfjyoIC8taVuapreGIM9wz5/BtJERYll2es4EhMWy+uLd
dPHPUmPrYshHbjM+s7D2qVD3Nc4kW62YTkEvaFulA1PHpqpaNf7uS9V+jverra9X
PKO32QHkWybSkKwXN9cQxOIt6dJLAJRRHmL6JpwUkyydJVhoMKLEU0J1YEiFruCv
Fuonnjmho9+xDKvmmUQGiHkknHuerV0X9pOCj9aJHxJycailb3wXb+atUG0As4M4
K0KyRXSgXTdmYdHWKGpcGYUvurwmrDPYOs/jYqEv23HIBqEUJZNYDbKriZMxbKTr
Guik7e5H3JUfK6YbLP2WQuhoECsV80HdFA22Jvd1J56xYPNxWyQTZ2kEbqbSKuXb
oIF+MNv4cow1CgdCLag12Nvj+iG1iVbx6p8C/l5IRn6WnT+bWw+74qK6Yhomc86h
SrjfYSuTrhFUgk2IcIqCwcO1xQw7sUECz4Ge8xNs6d67nGfpVdCmRMkXlMc7AZ5b
ZcSdTk/jiU3IP3JSs9oV3UD2HnpVHLwsyVPT/LMGEFai4dXoaBDAN4t6wguLBc4C
AHjc3aY9ssyOTSyYb8eXkPWATQ5CXKpJIjbP1eAOn2ju+iRStMfPGsFg6qvyuX5P
T8RtKVt+IRzInWr9DW16bri8keChTsSG5v4WEi0OLGhPHEgcHpHJts0RuXhsr90J
WhsNBRBBjsTJ1Mqx3mbWzHk7aepx8e1wVFNsoHIfN20Uq/nCrqE4+DY2QCvtvN7a
Fkc3y6GhluRA5AXoBjIUJ1wJNHdVc1W9qydPLqkydMZep/0Z1xsMlBNs2P6cK8St
J6UAoSWNovCwynnuOGG+3mut/F62pcpKCkrK4avJjtE76wa1kjrmpSugBao0efaA
unGzEs03yZy00OpUvmfPFZJOXgDCt7Hsnj4XVdGUQMUABCxehwacZP2wa4eF25MX
ZmICCruggGWq+meE+hv+AveEAvKcwi8Kub3mjoRAWD13ydFtdI1b3r2cP9JiT5hU
ax1VRv6iSHhwC/CIjgRZS4VmXVwfP58e33wl7R1/DHbOdnjeOV/FtioXcCLwsfUY
SuRFy7eEyrMIXIi6mait9A2bixxua3uBK3FOHjC73pK98HmEzm3gMAfCe5B0k2OD
1Mh9v6AdaRyRJnc1H8kW4aIs7EzuMUuiwQcp11ZdwQfz6MtDkbKe2vAoyvYNDsV/
pnfk6xE4sjcMuJBo2nF8tuRHtLcthK+oU3Z8SrY8FHxH7ouvbek1MyxN65ZcgIy9
7zK09NtqiqfUAZenS8Ut53N67rFJHHLnCOF7S5Nh/CnI533s0c+FEBj8nZHHZe+y
tEeEVf4Po/DR8lUYbnaja++Dv3LgkDg+f87bAx3xPivIFbB7VHovdWQMqQ26ARR7
dSgxtCQd4q9NlDcwHYdoc+u7SaeVp/IUSmysF/SD3KnUaPPLYm8D64qGLMSHAyRC
38WRot2ALet/i2SEDf9dYxlz1PJHYCFUGuCoTxmGaVE6B+ZHGMd/vyCIzBEB0hc5
2AwBxd/E4aMejBSf5fAZr/Q95gf2er3cvkkW6WhZTLqhvqsI8QI3I2he4LscL7Ph
ZuDbLw1ZXpakaX++g/1eUx38Of61Oc9836GS7m78KP0XKD7qAEoTYHXbr4/PgaSd
t2NclWPApcMPrL8eQ+IWCF9Nq9GrIWiX9xKg7cr3/1JYBorYq7ZvsyHKVkuJyvAk
BLKkM/WNCKzdrenHiLEp7WNGg5GirNJp0WlyaxERyehwiGsrjm4YRzDcAGocUzLO
NmlGfmPb3tQKoQxiZh6E5gN+UmT0tBU0soAOQWoZvnIq8QlDfWs0ZqgxU+Sk5cKG
oVRp3lo6ChQMMYzelLfyUe1eLAn1o6yE1kXIgPqYNBfxJ6+y1IIPXcZE49YevnMO
BfK1gnzp2zBQlIsRDfH0XZfgLppxLKawFZ8s7L6DUUYorbuaIoQoFQgBKKLgox16
tExIS17u4kT21MUI0uCVrhRVl5CRSzLgmhQuWBpXiwAxVpednd3yIjuWgo6+q/Od
hXxUvF7bQv23xhkoxN9fJ9H590d9/7JnetUTUP1I3+CRE9qY0Oz3wxAQPRk3896I
tEM7Ya/d+SthFaDtHZmNrk1cU0Oz8NhNxZrGL2mtX8WfGlyqoW42IS3Zpv10LyKf
8IuEdSOZP8OYR0ni3a1rMhuQe7xff5JZTRrEyM+ToyUmnSNsr9A3JVOs8v+emZHM
kj/AkWpJXfG2X3BSDCPtD8X/iMUf1UOx0LTRZoW9j20O1kkLUPP0eHNgiEwZMUKm
5aq7DnkEfG0yRRGLMuOCTsJewWU6z4F7VCCyw/lNzEYmCAZVDwwoLTCqgvSWQoPe
mlKYoIfxrXPXn+g2IdOHTbczbBSDXXofQKicF5ZaR5eANIFpZVm7sOiKxoxjMc1L
kAInStUD9u0ikqwqfxYF2NzT4lGhnpA1zb4n0jZ/4LbF0cWa5fyzsa3T245ZdMCi
XZB3toADp45xHLFK+ZF2mNE+oZjuy1oYL5Ioqgapy8EHQg5LU2ag5UvrTMKH3P+o
FFVDhv5Qvoe+pu21L43rGWJ+cpP017FhuOouyBdGh1OCz6X9FaC+EiJGwGhpfzWE
d/FeUhKrXz1JrMAmXVfhEayrjzdSzxl2WMmpvmLkIMx+wbH10HmiQ+axvJn+ChFL
op9Qp1ES5GT6jgG6psXfPqkVyIgkOSFBZiOC3RbT+vwl/htzJ2LHhCA21ZOB4HRh
EhK4cKAOsTqx5lkoSNbntqlIa390GEvVxgfbpvoIvGa8qMrvpSlfePqqC2ikOJbD
UxROljtO1PayCzEt2/OMcyD/NohXvD+e5B2IEJcYIQrZh1LOYjBSZHt42iLSmNZ2
mnDRKbJMY4HHRMIFpZWD9jdMzMII8SIiVKokReE/UyhOD/y4zyrHJ4lFR1TwDEWX
gXRzH9CpO0KCG/PyTmrC4PHyyvvXAgpp84w5SL/LGqPG0qSf7WPDqSntSyOpugR2
0Fp6uduiFSJus4PYIcaalS8QNvJhxbbgvpgwjiY06vl9+15Q9NCvSc3iiLnRl5Ck
1Swt9rINTJRjFITOCQ0PNV6WglVITiHgm9VuFxH51ADAcWs39JIS+vT2Dh7RUCfz
RTRZlmnFmFqN+LlBh1MmUpon6Xlol/5qAS6zUNv9e1E21VF7IaBzwmk8PcIeXHx4
6V8Z/n7Q3B9cmX4XyjRG377TSWckEvs/zfzsX+B95qW4kbK7qmWbum2nmiQB3nwF
NXfjdmdz7YvVV3CoL7dvmTD+aW9wNhJuB5JBux8GxqMtJyvPPs9/mQWyAquJ9IXv
71CSIHqUcvknnyIRr2FM9150FtaoVdaTiIvwSN0EPvw7ovfK99I8S3iFsu+4k48n
ITIq/jaa41goOQiWUbO3ZFcZAfYygOY/Pr3neKuluZKospPRKfzcFlRi/4mOc2Fc
ZnlXcIqkwW1Ndc3eGHAsIjqRHZ4shSxLaz5Xm+9g5N/rCAI8/0Q6dvAYx1C1K6UG
7wD91DCIeVqd4zAeTIGgjGW7UGf917QjSyb6gTkDV/p/ZgIAQvtRIMfZhBifGVTX
/vvyJVeHQWAxvLA8A32+VJmuTpvl2zCKMBxTZ8F4oQaFbJuUG5P81dlEy99qOF4p
VzCQjbGjfVP7wQ1IHnUm9FjjexMEE3dqfzkwhbCEWjyBIkGbg2kLM9BQAGtFh57P
Lo/VswJ1XJDFXcVsufriq7Nw48Ni7J1szyhkCrh6ODzzfWfY7TnMB4fdLh0sG1nP
dZDaSRAbxKMYB8rqDxSzJRUQqEDWNdKiM8fI63it+RzCAoDb3dTepDdyA2AGX5Kf
gm6Q9L3KIeNZCOKqdanTBDHhGloT/n5gsI/CxjzwYcHKi0kNAgbDMC7U9wpnykK6
wd6DSAPI+uWmnlPW3kRPpOuqh3yqXquI320GuVvXjYzDYtjD7Ehr+STbdChDZYRs
XnXc+BbGOaOgiDFjU3CB4KBjP0dOrIYt80M9xPwYE5W3ovk89T6hOe7/kF+tyPjI
0SKOApc4C/kw6wt+6Bl/iHg4U0P07kXl9CCbhob31De1efYMrQ0ei3MQATP6GAa6
cfxhwnGJK+V30jAChOVWeqpdbOs0wMdpXVFBZnuautQ1pZV/LkAGCgiaMWYUQMpy
2DtvQz0xi4YUfUT2rIOI2+qwuq3zzNvX0XaaaReOy2fdRtp8v9ypnGcEmrUwaF0d
msPRTRSQuy1ZAayhJIjjU4GUksDxOL12PUDSPlZrV9EAp3eTSkRvQo7B/kNDqeiD
FBP1m6ARtXtuK1lwzR14jzfo3jxmoECICKV6xNUrjI+Re4L9IxoaKHSAoDWk2uQm
KV6ZSq76YLzvWeJs6j4Y/UGhiUrmt3fhjAFOAM12bDtkyqJy6KRMnM2cmhZq5LDY
jwcLO6zmH3LV2F6EX6MiojalD4jg4lTQ5BQvKduZIMn0WWU1gf7TLDgPLFFyzT2S
2s+RN/0T8vAaQFknPi/pkhYbXpJpJV9rtb+bygZatvFl/Y3kw4zQ8gxG8r9jKDHk
Sj1jErZW+JIwhW89YKYQJw4S929NK4j3NuiRNYFNo+xQUrdf3MiPsx3UGu7ZGZeK
PBOGqoGsBRp8lrZFoTfjegsMkB2KRCfTB8jYPel1lWSqBU4awuyv9T3hfHER92GI
5InU5P2a6/Z5A0iaAgqe7gWt1ARNzubv5c6ZxmauQxzqGdvfNB9WXfMi3Gp7mQbZ
q3ZJaYzcVmke0e5/PPpMvNf4jIMdV6mlzODav8+1Dmsp2m1E+sQp3J8DFNa+4GsT
ZaIZGTdW0qX8tCHSEX3DbwLVKvVtprq3v+aqjYjzwLat4M79WdQgWVSuxVo/lh50
7fWOM8xtVjTmU9h4PzcoAX/ofFBtskHEoJS0zZ9SZ2L7xeWslQ7pvU0B9ghLFfs4
7ZR6iLdEyDL5xdCEWCbmpIF/MOanWbUK4o0qInOGMusg8Bhlzljh0W64swdgnsPF
AtyrBJBxoHba6cbud4HBJrKJ/bFUTcBs/LcgW28WXv7XSBp+wrAdtIifDMue6zbe
j3RLWd1ac9KOqZ0tC0dKiJujX8KP0gkclX5wUQwPcgtZe5cPmk39ClOEok2pBCvo
ZGCq0Q3SC6d9irk6VpolanFPsXiI0/+u8py5pIMEaJq7sd8TBQq8Kgp2bwnHktDc
VuSeBjBZjsWdtk3tFIEzWlZvVpKsEanBsevlj0t8skTERKh0+w3cyeA2coenvVGb
67Uhd6GQWuGat7cseKK4FW00grl4CX5gkEjsGKVmh0PS7hN8UsiDOw/yKpiXabS/
rYm3qMv8TnsBkf7saS47PWaVPWnGXcXswChggVAvMRdlp54gBf91KLhDkZWik+de
nGfB09IncbVdEM7UlipUtJGqX5Hq25+l1Vvi8HLxpLPecL3xtEA2KvG3fhXjnoNv
/XUBa6EhyszFp1RqieydsCThiRyyTcdcvPHp7QXTuvlO1FeGgvvl9qAoTANcuTsn
pf0QKJt1nokQNVB5zncBNrxWWlRckRE5jSegb22l+EsABjrcGd8D3Av0hb1NhFLj
F3U5YLz+8v0TWbAOsSmFUzL1EwlapGdpozpNTPsvCndDm2nBACCGNNXp6dEiIHQC
LMAlqMmXLi8xnukRoSNtASoRdEJCam2aWUXb94ZpuLfrI1q1/STnnhp6Bsc7RrqJ
SR0wVG+jgUJTtnAfaycPuTmPyQs8Q2b9v2tS/PGka6LswUIe4rK8PFkMa3Ab/Pn3
tSKNoTwfprxbLhfCzCY2+XErwO0yBHmoM9rVQLP+zNAQj4tDC79tjH2a9C2p0Yli
4VQqH7k1yu+XKoDS92M5bHB6J970V7lBgnxAo+EyH8M2yi7di9ls560/REZgaCoj
VblbLQL1SopteFARpGh1A9N72WdVe4O33mG4xZzLg1uSyKiRw2p7QjiTiGrW67+5
l3As3SRCXongLV7ILT/tfHstPEif0U8+KNZTQk+a8Bp5Sg2zUno5cJQ5mTAlBImk
UkGGY/omv11X1aYV13SdQbipH/J/JsjTmoYjIj4aTvMoNXQ99TmCFFwfWiEG8QMN
7s0eRy+Ipsej1cyhc1DJ0x9Nsu+06pSNKGmFVlDfyh3KtTdk9th+Y7L8HgMffSUD
pmZkSa4RIoD5wfHuWPYhgnCFqggsHEjNK5vp/DzkqoyS1S3Mbl14GZakGGrWM0cB
Wp8imhNHEXd78HyqtJg/amuJT3/yEbehqhdcm0CFRGXLqCxfXeMMlEJBybW0sZ/I
v/x76x2LFt2BBb+OfFY84gxNs3nc46MjP7TbXGVTWjnDmky2hQjsS/atjDxT5SCY
dLqUjcELMysMW3EfwIzajt5u0BELdLV2VJV3vY1Gbzg+EaKoswcRDOiC+w34Jw1y
b9T6L6mwmL6K3TrNXMgpckcSqo4KMFBK+DBSc3zTjTZbnUWhjzC6KOgZCZ9EzrtL
6ijsRYGBMNbrVDOhUocnHCDsx9+KUkRJIWSor0ILWvdZFPinznHZ6N2lEO0T0SPV
3TR/Hm0EkcsygbZKF16SNmDHCaRVHg4HxlvrHtDOGCERG+4yiIUcC340rp1wdoUX
J4BZxYZBJyL/B0kWicFiyUzABYMV/Bj03KPSKCJdG+MJ81eRLlhDA61djCFwu43j
KJWBrKzB83ayT+EFXkWVaAoXZ/IS4TxFeVdy4i30iXH84a/o/xQaqiHznyt/DSzO
TVEvFE5jA18iSK6Qh4O2Wuo4skVxT48woUtantMb7c2McXHRaPOy0MnFY9+V0w34
ddemU6Elxp+jayJbZ1hU67ARhsNzTJEtZw3PoDluY9uLTCDLmmfDwt1r1Gn04gM8
l5oErBCp7BkjNgMm8lbMANOMDluQO/mhnjFbKcBf1Qgz/GUFzuI6Ky+kTxtrFbTP
gNENIxkWUWjP+EjZRXg6Q0Hp+S7GTDMXyHW/bD7VrRmExt0hV6aHheLxlw091wau
3weOmeT85QEDUXSXe/5Vyo6hJeo1JQwp7KgoXEDMY7ekKVjfYUF7Wieh5P4oRIpW
VStSQNuPLTLW7h6M4PA412J54Bkk5QaWGU4NZzY8UJdCscDZqz5aWWjk6+dU8A3q
TEEzvVkPmIOgCQVVGf3MRhlS8UWMJ0Gh/a4cBWqdaP7XEuECFjiPBpVmhRi4M3IS
sTm4yiE96q0Rq/H/b9T8Gxv8lphICus+UAFErmA/BE5T/Be38U88X7lysvO2ZSEc
xPgquu6+KoijEVPyCfOV5i2EBaLfhgXuTaJepoShTTJAZHtWLmCsU0V06bk04mQ7
+HRek8lOS6VJvlM9QcHs3nlPMSb+jA33ZQq9I7wgDW6/LfpB+eh901ZYhjc92j+V
xbe966BuaKp1tTp+9K0Kx8mKXtZwVvoJo9Xf8SyQyU3qDsLIgci9djvAcIXTlqyc
JbqEjmppyz0xM6Un0/pRQn+ZtUPWUM1te182IMNHcWNA/lAgrgFi/ozMUUXhdQFS
/r/E12TE1WpjeOx68edfteNOluoEzJxBjnxFFxN8PElHcSRFtya9gzUgbONazUUR
aMgwjXtvfPw+1tq5Dz8tbr8YrGemzJ/xDZlN6CN56uR4tqZui5WKeCc05iiSFWcg
C0PX364Pjy4CaFsqzFrFE3IPCL2XP5ZPS3J11QItgOPTNvDG8HTnAleT92nvCGc4
CWA3MpShLhMLYTlElhdoNItxmc/G3Cs3bcOxNLcOV4R1GNqiK403kvn1tNYqs7bI
YBItCtkVbwa8acCOhxoNkRl5rC1aFPerqjr+rL9QTxw8CyL5R1oE1lguBFbSurRc
YahlOAeKh6TZU3HSfiyUmpwLIkLILbbLz7h0aN5x/DeLoGAx4KWhlm3bb9a0Cpe0
Jb4/J5MTRaOEgOepF2tijhMF+zjxDfz0MCGKpuIPaTyXCr0NFhG2atR0ctO5s85s
qniqEqzPIj7l17ikNmB+23lfJXQDFnuPm4MioPLuno08dJRvdR68nMGoZ839RIH/
7xk85JXv9kPO7GueQOEbUgD+TBLcv5Ju5PR1eh3mGxNkMjsx44dj8uZRU1OiJlXs
10ve5yI1+JWBH1j8WEDA8bQwCbvNxytTHtHpJAZiul7P/fLzBuWHoh0O8E4wiTPE
vFIUYUmanMTJt/vAHx8KQbZKjZfC4uBzKmrafVFYUtHS5+Oe0WH52xeGJfVNi/zQ
ZZ22k/dCmsvA677k7FKGv6E3OfxY3ZZD1xI6g5LORLyVUyCUEUillBVZPlpbvBdv
Hjd90Cec4M0peyVSA/i+AzXW8xQzNklewcZPRM+9EB12jXsPa4ftTpU0HLA0WPwz
pjyj3L1t+PPcIRK+jE52RtFljpLgqTdeBO1Y0fBYBhddsHZYHDSP32PTJqTgwbCR
CtJAe6/d7zbO9e4zmUmQxepYe47jCF4RCzGL+rWAHd10f64MsO/qTe4TH7P9fN7X
ZnM4ITABpBtX7FvsPH7TSO09/O3fDhfPLtzY4pbtfGoIvmZUOlO6WL3y8qkvgdGY
LFEXMOED8bOFqeQYemBnO/lpzpiA+ux13Y7jyyLsxLUgT/XBjwdrfkEQbqNeVCso
Jg5SHnZ3r0+6Dw7DefdKlXwmGt1eqcgBtD1YzTDC1PhCwVyYoNcHGTZbBwOS6Tir
dE3LBi8871YXAnoEgEEo2u8QA3uTauww15ErdOqpYXsVgDwLrT4JhIwkiwPrEctT
4Vwj/xyGGk/yux6mYeDKFRT4gjo/qY1KgrJeelcscK7FhqHu+1TuU74+eqVixOOZ
TZNOT8Y8c3Qdwj6iRiyRZVzfzQdnOuThCTirZpjHfBsIXbDTUSz+WCP+LSbrlqE3
S7sWWOsKWp6nDjd7n+peO9j6N0PUZZ6bFkRJpMP9wkXh7krXaGqyfFCZzr7UwBUF
uUuv8sNtR46XjEsoCfwSdLGJd4r6KSfPmgq6Qr4GPQikNzets3ly4a/6gTG5BiGF
HKaXXR+qiKfk3skWTLBbty74eOCu8p3uJy6V9Nln+EsDfiyjy4ALpNV95MVKh6QH
5+g6+vYItqu2A76LWmeJSeHOEwjXYlYGWExTIwjTFuVITuw63MLrLGkbADzRJW3d
oTJsYk8s4VmnlxHFr0vn2FUymKpUHE8eEPii1FPgjFFLU9HjI3RWylV0q3xyiVmp
/0GDNEoqVEl21a+Ps6KDUTn2xJi8VFWr1ij/T6hUF8OHowYqfmsEjQzSLoQCyOA4
7pfzo1WmYANWutvOp5tRMv+bBiNjgHiGBiFhhgqbwuNcvGnr41eWZGLQRbzB0RXy
I3lXQN9ZJlnor+bnjE54XYDS9eYfPA39GEGqz6UEOBWL2I8e+ObzeIWrMxKcLH31
ZBZ5W96XNUco5sTpMOEHhQcx7pOrseRd5XYt1ixzM8qVSMzC5WPardMKD+bNS8Hz
gtBlmr2fRnwQZtLbKIRRuDdkncjCQccmEHQPaF0Pz8Xk2JwgBtsop029N6Y7ylNd
pEP1E8Y2LSSV42rcilN+9yv6rIeAgn12Gi8kBddSWSAamsKOIx5yiYmtEkdxbm/j
60ObB6GvNWzTBEmOwu1sjcJGMA/sy8adWfAIgBrNyVwBFb3tRP95An3Coh91LAyO
qOsfURyLXzrfVZmBOQNYcqNm4CqVAhuRrZ+UsVsoWDRnPLso11ctZ6d6POgnuLMX
ZgQKEV0ucFw6WDc17xaV8I/56tbImpuGeOViAXGH3OhtRsQPzIBmbYPyKcSu/Bxt
CKnVckTfsa2Mg9a6Sj4MisMlki4UKPbt/3FkECJVz0jbZcuDzpJll5qa3tTKe3G4
GNGa6urxWOYTkvR7LdWplnCXvZqJu0JfUqPzQPUgnCDew6qmPjDtyNwEI+COj9Wa
tHiH0tZAwIhRfJSWOwwteSBB9MdgvAZcNHvJajZRN3RtIMFh3nw79fYmO4aSNznu
ByHNUMzAuZ0RahVENQ37HyQwJCIIXItw/flVxgYaF4qER9sgj0tZZUSuEgXcxJKE
CmdkBrpueh9cdGRDL2vdvmLMzgzTIpzET8rN+4Ugv1wqMrAUuIdfCS4KWlEa8oK3
Fnj2ra/3wgufas1PXZ5zKgQczZ3dxjVVCzvBDXYD7euBaY2sAeXF/MaCgcWvZ2R0
7hZuC2sAd/A+rz9nBrQOVjElSQghSx84Cgr/c4yE4jpqpvPz5pKwc4roj9XAqWzn
1d+4L4SvLcmhABFV/aHh3IAWL+lizSO9eQKjmGhXZ9Ktbs6FkETksmTtdv9FhKIn
a8FILzNbW42wrbCrhOXTZbiqQIvBjisr8XsDrwCI502NjgkoA4mWGo3IuhkOKGaO
m9c6bb2IKpSPJ6NCNV83IxhBb0t64KPqNJAokIgYHUyQ5CJtXlEqOljJCc/H/bMT
Dz99q4/BdDRdi0PskDlWRAayxMphvUIwfSI2hIKbdSYmZGnO7lNHl+6XuY3cFYMK
fIj652wIulzuI4xsTdb6Dl4G2yc8Sig+bYRPtKrnaLAe+cCXfF82oV05KhtrZz/m
SeI3MNavJSZ+SagSGvagGFuyZ4h65c/QHGkjdIYI/NUjNbNlR0PkTqp4/npVKq65
UvisNKQi5px7e+6flCgafU1hdQb6Jwy3Jfud6Vvtnw4LdWBN69GjqJUMaK2+oa7T
IqJ5s/VqaBajJ0xZsJGyIlkKLgrsmbnwYVP3RSPxa/hMgrfS3GCQCDN/8nzQEkJn
9tbrH/o+oegbfUNC/8RT+4Ev7LzO3XeBu1XKBImTtIWxBbLp/8/y7R5SxnX7J0UX
pYFp4S6y5+i+qXkoOOY3tAjh2WODedsw1+h9tsdCLcO6PIWbxziKkVldKqd2nGd0
XznRhg1v7Wb3zaV6TFgaIyRlZqN9EM9/ftsRqar1sGNsDszDWNIc6mwdiCdNn+Iz
UIxK7MDfBkDy0BUwlX/mb9aiThbNRVYEC7Hh8vVlK8IwTsLLxCTjDIHC85dLrQNW
kQMYz4SqXU/4TB/QEGRhd2lbd15m/4q1BnJLaUGGFwWfA4AFAvzkLdMhlEv6rtUv
Fct5fplDDBzP66gvqmEoA2qmbQ1s8yy/ezcqmE1BEB1+GvQKoP1P/fy9JR7cbz3t
CxtDrhlVlPEo8hZ6XGzLuGLi5BpV4B8Uv6yITfG5STRI1R0T38ZonrW83ox8m/Mo
R5ch3xd2UncmW50EGrM86F29XoMY3E85zu9gFLBBtHxtsRO+bhJK9vTRYJUb6CcB
geznbGWVWbkqmaEEXq7U9XM12l6m4AjeDOR/FR/5BCPEOf5db6C+cMQo7TdRD8at
EOH9c432ElSnLdeFCLDpq2srLYL3nKqKIfRIubK4YqxJVx+eaCB0Qyvn82pfvuFZ
I0u7R4NsfHKIhVf+pFaqb2neXxIkDzMTgjInaX7bLJWCT+Fh6cQ0XNLI5VGLnSmC
hL/+GWRgnDl4d9kL6xbsPPXbqZvf0J+g6/CAblOB1GlUa8Ac/UvDY79T8Srwwsj6
8I95yf4crTT7z5UkXQXId948gy97QIPattuhmuiErlNImHmH8jY+CpW4AeaWaX59
L62SxGh+/TRoFubMz+3OZMMzGfJCdhlpusvZe/Xxzb9RIuWMwclobh5uyYlmne7r
1aeRFRXFuyM6pUX8GpPyfMkcBnt+5SDDb/UxnhKCGdVnFpGpSECQ3787nLarQhLs
vj+hJWM1ra4D/GxNINOiu1vd58XPbk+opPmLqUsewXSFzv1yXBasnwH3WyGKJWYZ
m8uYuc0TA7YKOSqejA5LCaP0ycvlvy3i4yxL7Fh+WA35CMhavlObMfI/6aCPE0LX
CZAiL6PLGI04SOZH8Y989m84ioxnBOb/X1xMc0Kbtqu6b36uTk6owqIACwMqhiY0
7YY7Fn0X+2hWrABSbrr+mZVKXZfZy5MGshGWn4vMTSuDH/PC8X8MLjmbP6plT0fs
WVHMVQDiig1uDyBqsxahgG9MkHGYylFLbdfkky4E3f3AOmQnJeqKT5MzZG3FAVcm
VcE0rPiWlNKeBqzRap9ATKr1p60rQgjnGcM7sa/omKJyKf6a37tS+bQaXz6sN+oi
ZaiNiAy3ojubageGezP3FOtBOcup2scHk9Hz5k3sYaT6sSwob/K86or2BYdZyFSA
CVot8aBREO9DnEA8lzn9QveucdvluDCBB/igS5ub21vMpPmVJ6lRuk0UZAZwzVkB
sVPRU6Jkjj/hSVfdQyhfgs3286ASAtRJFVZTyHi+FHJL4sWWnGORuKkjTQNYHAHV
EAKH0CJ8Kx5Yym5bplpxQyinWcN2Y9rKtUmZwfk/N1isA0t3tiC56DvWvO+lXf0n
1ZceCLgk60pfQJ4gfJh7hiHn7V3HTxd4p/UEj4bVBAuULMJQd3DVaPfSaIF40pAL
kYiq8WqeM7W2/t11zu9Iw5LbTfirsJVNZovGC20Nxs2QrMkE222ujhIG/G3rv+W2
Bl22d5yL/lgo6coDTNN/yXF0uxeHK3fzsVH1gOEeKsSYGePmRcyz7GNm9YJoYc7f
ShoJ48reJCsCeohFwVWPrHLFKovBTGiFSTgXMIQ9Rwu7vHMGZK8hGKWMXv3LB7Nw
I4O3WsY6hKiEe0WHhR/PSsU7vOW5ZlXC++PDSFbUrzIQz/FdyORCYybeFEKwABp8
gYFS4XKJiXTrjfyieeY1e8jd6+A7ElZMRXh1OxY8Qh5nzIriX/IrU4EN/k/DG4ow
mahhDZk1J4zSsBhTbCHCHwIQfN6EK247CSe8xll8DalRGOFeEIAqF6beDGmy4j9m
7siRziP0MDYvx4zEaaB3rUgBNh/a3e4iC0zBrjLJiyD6J8VtH1OipuiA7wz80ASH
IFpqqwCUGCw+dzx8NKR0qK9Yi8K1er2esupsUcdHzKOnq5zYXaS1Urw6QYeP2b9Y
YNkT17jK6sBzr9P6dq9vKbmcsFa7bdLeDIn6voUHcj2nxwinALyBEiiaf77Dja4A
o9bManffC2gsHJ88trg5pXvvZe6cimH6EvEgmhCBygXziRD/5bC1bWOnTnprAtbr
pKypbj2a6m6bSM0X2Ivt70izLQOmrDuzuEPpvryyFMZ9uEUa6xNfLz+FdngyGWSA
28Idh+xq3g7xbM8uEPDBidA7BoEcmyFjC5NySvDfrhHCCMHbWxRJTCx8AVVJpQ3c
vGPf/xxmxNA7+WNQZmYYuOQpFCLabZlukbhlnesYBr1VtvUKqdpLvebN3vd+oYlV
48aotkex/xvpSsN3qodzz0Bsa6B8DhSZEBckQxI9WHbpJqkR/hbD8uazWShi2Vg6
LQN4tF4DgaET6b0KTLhX+CFykcuOsfmM9esQGfEjmX0BeDe1or02aqvme26+wOOf
Y1Bz1EnioP4YuHbPp1rPMh/v/4ONjX2eLUkMQ4k6X65lkSECh3uCc+RjwbxsKk+n
jiAWjO465xL8ycobaNgs30q6jSLWvbvAqPIVU3R7dvNw0oNmal4aTcF2KDJQWCiO
CrRvnglv0lJmoVCI/B9rOhg3hs2zGpWWTmS8ulsS5Ndq7oy1nrOTirjr6G9r4ztP
Fl2gfU+kF6O4EL/vZ4COASJzLLe+lAcXtDXBETRMgSzu6QGD147VM9uApVvRBKCE
2JhOvrFbYxx2d8ZGoGHqRm+4vL3C15RV/8J/U3lTY/IV5i35wr4RG6LNamT3bFoN
uTS86CIfb53fkVQ6r+JUlvy3aY9FT31JnjnMa2jDGMU4zavq1qhiuVtoWZjkgd/z
/+mRRU51RuxZYAHsHbqW6LVU/SegSaz607VeMJmq+mYWBun26B+ntAanK6LuAQz8
bP02qZ5r9TOJNE+7fIrhtDlWPlkcSMe1hokTdeRaqFMNpLH4IAijVqMz77EDqa2R
2yVqmE7ll9kNvuicPYJie0kiNMYO8aCjVNDMGANp5Pi3gbvnsK82M/+dPsNn9QdF
ca8rZUUQ/fxUkvfN+ufiGK+YAT2ni8opmoT+8qwM/P1K/KaUPMH2eJfyfPTtGLUQ
rMO2hkDlaCQmw1XzCedHtJo1PCAm4JqIQBMs0ah9PGWpSyKo2pXR1a6YxpR5ogqC
oij5s8kI0jxBy4xuMZuVqF3FRDrMA3sbcDO6H7cPQ2kjQhuuQX006unB0u9BNsCK
9+MsbVY54wM80WmTFJ9qyKh+lTRf4sW0OCIMgQ8ezkU/y4B89RU46Go4UHFiMM9q
a8bt/VAQhVJ3TI/latoWXDXhbRRVMRq4mkemntomS/kKBcOTdjdhAN6JuZNddZcM
2g4DJtNiyab+t1s6XmN20GsYcP/AsCl5TEu9Pt/sIw+y3AmPUvwI6UzIOGgsvBUT
aYfGdtQv6MwRs/vhBuS22bK3czMBLroNP97IenLULrMVz8ZnMboi7cmHp46WeqnN
imoqQn2bvU+M2AcmlrjG96vEnyvJq/c+PqM+8Ph6FFSVsuVGN1CmmuPxGmXdsPry
ng3x6UKOvoX5VrWCNSJ6il8xhnoUCWgjsLrhjlluP+sJA+Q2SNdpiDuBmFZCg3XL
QocYmNKy5WxbO9o2/VZJGdpivBEF6exy/YvZI3uibvQBpp/tQXZfqDjnwp9O/rYs
tpUI1VBeo825k4/dT93T+8nLX3ONK/T4aGsKZ6Aw95ze5+joojE8p7eIEggZnNOE
hsawa6J7C7Dd83ytgG7bWLex/TjUHLz/XbqYZDvbKODw7I3U+ELu4d5VVJIQUzXc
rIBmxFXRikG0cprL5r4MZ+eMHBz8dQe6/EN3o9YLSBNRscqEPVu7G7P4IO1P9gkB
hBznDpwc1kPnlyEgaSJoM6p7FStrPI9pdLZ8/LRQx/Jz4M7El6C7W9q6EC/4oobW
guUAi08it7ahn0xyY07qGcvxpkVcre9kWnn4CalLgPelbHzmbMoXxYPHgINFzjmk
sFyn8Q2EBFx/WcoBpZH6xjzFqoi3k9aQREoEnabj8CHaFuiXdAG9SCvpgceDR0p9
zs/Nj+Bg3d9//mfHTDXiIl+HPIDuNUz7roB9XoK/02dTXLrUBRf9nt7gv71qSrAG
DLR8d0B2d5uAu0wvNReIrKbVUfJsjByt767KCZeglRiiij5FxkZlB2D07zfQcOb3
O0cxNUirj73XFPmWqilePD5B3YyK5VPr56jCATeQMk04Gw1xIqMMJ6KbtzWyC6Bt
b+08Ge8CV0ABmuoAby2FhlTOR7ruaxnTIipWHUGa3mACQ3vdCYlIooswKbcEwPOi
ZVqPE+JJHuUADGUl5T+W14Hd5GRbYzolA9nZLirFVItKQ2Rtfy9UmK9QlH1HdVgQ
ghJ8VntXmufV34iNzMKrF2niahxCZhAcFHNqomRMWq5TkV4rdx8S6FIIoDKNrMni
btA1Z2L1/UguBslkIrxrTh6mqGSPjwSYxXnEGeGsoj+tnAPFReYtxyeUijkd6zkd
hwLxJ9LJI8xyiUstXmqcRtXn1T2cebi6EdX5K73Eqi+i+B81plUjr0l/pBzDLlbC
mmPsvBiqM8pmIhWfuXUl0S3dfJ1hhDAmRhb+lPg0ES4=
`pragma protect end_protected
