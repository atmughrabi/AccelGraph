// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WJWZevWCm4MR/yJ6rJ/TjaVAfEiosnRztIySKDBQnv9UnbjV+9jra3EbmgYrf5gR
GOAkUYesR1wZK/QMmqhqRF6PMTDb4T/iheV9AJYxM9KE9q/y54w4NCW0r6WjcDj1
UAXUCLcT/FKwpBX8M1rwAYkucEtNx56ofGCp+ZWYCnA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27312)
0KCkFHYt1k71XduDgroTPiKxuISt++3xvryG3t7MO35R3KK2tv4cMXYLRhSMwZNi
iD05vVXRLaqyFBGWBHSAUiqYdso5GSbHcDOFv1uNRcL2LRS4X4f2Sgr3zZs8I1IU
cK64JR5VhqVl7jPVBrmtmxuhVlRFAVOr+8rN6l4G4fF8tIKDWjFOpkYlopuEfWF8
hwD0Bjb4ooFFQzt9oaPStDnZUlnvFrqOP5i0jfIzXq0jEeEFrXVsGy3CX4puDkC8
uVQapxavqECsHl8zfFtIhbOJB9R2CauvLpHLljLxrtKXIRFtVy99FFeCcHnrBGr4
cPeDl+v9ItEfyyUUkTkKhfWQz5Hzxus7IlwKGirbkvF0dHnL72OswQSEcJmPbggB
yWdlO5zcsGLwtUAM0cAJGfbH6qp8ERS/iSwGrQUPzs51TytyX9VVegm/RKtXJvON
+Jtziyppr0sg7Ng8bQXchpRbHKOaNWyjTuGJeM8FN/esuLvygXftEqamN/OHVDix
m7cDRGwp99NEJ7P10uI7E0m2wm2V+C/ItDswc5Ke+mvkCg3iYLQKdh26blNseB1o
PLQKOTmOMfXxZ0Wuwzj/FkSjNGEhl1EgaOaXFqQ0S7x6rPA8v7UGr14MNVAtr/TY
lSrRA7x3fqoQfi4B2OxCgKwUTiSOT30nF9jZTlvMLGe7vu2SejR2rdTgHMjI7JED
2g8oki5ZninjNsrV5R1ZSit15mlcdbSAqw/OFgl9ZV8XzuOEI36TjqTVSb27I9UI
pVilqTi7GdfKvY+/zX3Se4dSNwiYiJBXQITRVs7Uiyd7KX/Vjwzh/BFrupiekh5d
pcJqKYUJjka8NVigFAYocsKp9fi25hHDQbRlnBWTRTr2US/6kopS//62bOjW7YRj
pZ7OyjEVaaRcVuxtLwr0/n67NPIfJTbG4rUUhhoBX0+Ys4H/CGuyCirZyRhI+Vk9
4BjewMzeMPhO0bFwSuO38/KQAJ8wG8U47ezvjGoHtd6VEYszYgAfg8547MYR/vx2
OFJ9B4+ZYh0KR6Z45M7YFvrE7Ti5NTQ7eLJBkF+64/QqWeVi03qlPXB6C/KZEcF+
AoLwOkgel0PC9oV+1RXNIYKBG3ZLz+dDpEx13Gaw4PzWzz07JlNy4c9HHaCfKsPi
FtdycKkKNY4w32TtvE0TBvsAI/qQ7DVCVQ16mr4V+fj6X8nypnm1x/jnb+91tkar
64DEDEo+ZjsQep7h8llV9tq0QE44HQ0DR7JozxT7mN/Y66+eHl7pxPcFRfAt4NhI
2tH9Db14Oyqzd8s73MKKz/Ee3sR6LpvW+zPNsKDQMXyySAQqyyPtVOLbNAj6QbpZ
T87QWFRuPgJTqfDMouzHScQQNDXCBHkQd/TnGt9S5n8fPi/DwiL3FebxRaXgxaLR
Ue3HKqSIQDkt1kNeHDRk+mO5GnoZNDIboR7TbgAM0sgEGhBTDgeb5LvR634sY3G8
30bWF2K8gfCl3cgKtzqn8ad8SxYimom7MF0DMqZ/nwQscKOz/bQujTYepiVNt0CM
Os7LjyR9ntRcYajXvF0Ysipl2fpxNA4rUipx+6mLxlE0x5MpVgR5uiW2y+SDXdH4
tiviNUt3dt1vk1eW79pIJ94DB6vnKJDFZ5LvpO5hW4V7RbiMzaVx6N6ccQN6bViY
qxsn4d4pp/nEviIarWblrxGyt9HIJzXnPby4PC0A86IHzibWUAtAQETi/SSsRhfa
QooJ7Dp7b8U0pQ9zbetP8t5sq1iOB4aNHnpQe/yzn0H8p1bs76Q6v4tjlhfvuFjg
fPWgf6n8iEY7kSwA/V/gHTW+5GAYt6caoriPkunkYSgfInUZXBF74yyC9KJOj2xx
E8c+F3qsWZrdU7EkvP9kC+HjsTHyw3Q2SolsgyVLXQhBU0eY8zWvCA1nvrp3noNp
VJY0vbUJNDDl1X86k8Mfju175QVKSCgHjkExx0x/T+lmg3JcokUazeOLTfFsLHxC
QbLqxDaiZIiZf+O8xYM3GrpeZ5JBp7EvUcySXQLQKkEMnVuoh4BalvmIJavwee7+
oRRPJXSssKFvchrjZe1tsmBTCq+/HKZcrEDdb2992TDtU43B0styAqs8MYPhbysr
InEYP1zsuZUJmBwux6g3pYh+SU0u7XU+tbIOCtzhgUa5PB49P8Ar9RbeZ/YcUTPr
4iF94sg0bYUQUonYzyj1NNCCJT0saNttanLQ8KXV38zib/OND18bdkUHTHteHvB9
I8AOlLj0yS6lY/QltyePapaiEOgI8mnnka8QOrQZQ4mbxZKbNrIIuKLTmPnEONky
LzFMvJTiBsTKq6sahkciHaM3BjlYRciujfeaTdJgOyT/BTHeoowMeQYNc9ggCV1j
h2G7Xyv2xcaMLvPwm+A839BhclCweIs9SpXAxdzBTYcyNqnmDhf3biD13MhrLvTO
gInXQxR8BPD1JRn5bguLiwmuYiCjZ6jyCREZQsuYM7hloLjFgk5+qS/aEudXqMJU
8QEQPCGbEHZjQo1U/i/Cwgd9robZigw4YoatVNLA7UoZc87k5ZYnVszum5+SHoXV
7q7PR85ogTcaOdqtExdn4in6qyHICx9ReIxKGMOcGE31VVZ9hxNsIfrEAO75i+SW
fYjpYhpkYeoYgAeMLr8Ryeh7Iu8QC1AlCJ2p354uFr04TWDs+DgadA1rj9nJZeGA
MQr0n2uE2+pdTq/Lg9iwADQJuI5XYTxudSKVw2XAPyf43yKFmneO7qx5t5Z6Kke3
2Hya53MIp17ic2j07tQl9wxegIT3brLS21InSfobPPs0WIbUR7ht7b+OGc8wU31E
7JYI7/L2V6yD/U5vlwvMyZQsenKgOKnTzABmMQigozBUXEpR4/0hdAhKj3K3yEJZ
8dFkX7FCaSZ6xEQ+KJfMULoTr08kYxvIoCdS1Ny6APhzVffepM4P4C1pxxje0lOS
QgeD8Iu/brLMRwDGdMVdhIkfyb9XjRSPaPPWraOK7YOPB1r5UytFhy5VVT6T2ZrH
GXUYEVw98qnzgElorR5czt361AxhNadmKQ5agk83IEKie3iB0Ut7HoTlcTv2uZWu
PQSOsaDupy9vTyDiswElDS6i6orf0uvjv+OH2s+8seTurZs7apdxYNGGFsI4nv4o
97gW09AdAznFcLwDJAt6vFTDaQ0eVpEeNiC/t16jb/3giFlTgdhIcPOeQ7CMo2zQ
TNevB4KBR2avdTcPjSXQDUY7siMSkBeoH5YQzmmdTuJiMxLnQofptOe4L68tmOej
ttbi+6wcEAeKk90UC1STjswJsFLbPe/wPg/YuIJo0a7Rkh75pS7EX8GAugCX0m16
c22LTE8RHuGWyw3lPHcBPxx6wY+iTVelKgRQ8lJcN0UE3STqWDqs3P08VSaWt967
VdVvVrBstoUOL0PLluRd+Vdrw0grpCdegxmukG/h3uXAgMtYneZiYyhFUcrJn3Xn
7n8qPmVNflIimq3fuiKNGUHMq80DRoAa6e4liCycZO6fVtggeTy17ujWZKPfl7fm
kczVpAdQNKHDYY9/ApknXMuSCB+G5YfqcvzWcCavc+t/Kz1UVV5OHPZ1y9OthKSz
RzyYc3oIaxuygXQnqSpo1pw3tjtRH8+nt+lP1z/moLwN34OY8NKTPazHbrO4vAJ4
Qs4Gm629aptoIXPc7AsMpaUG2Xr0cT28ygE8PT5SZeX1GeDvzYlEhaKPr0ayklhF
ZBCc+cIXfvdiWjatk5fYdxmVaC02D3WWnPDzsIBz+pwL4GK1I8wrOJg2+0eejpx5
yGkZxJl2dQdlU/3T9pz8b2H/ufFsvL7jUFcNJOtEWEZD8Sjpgo1kRnmW8MWxP0n8
GbGsH0sFfXGyhan4/VnyXtrCICShICvDEApWGdxBXIxLcHYcrfjm6wDaPxfA74ni
AvvU2dIOv0Smmj4K9NmL+Zf4PfS2Rh8PkryEUU3N7lglESO52kPJs9IZmJb+vkKp
vA78yO57HqGW1ydO8NArr/QDoDUahj0Hmauzvjx5ni0uysxeKv4UlCEuljnEK/yK
vb4VQGSDnl7DSoq2GiI+LaKKvfPLMW9k1bsNboevYMtq19V/lDoaftEgeXU7Wcb4
RryyfHUw2XWTrP4QGzDTNpasKKHR/Ifxk7MmT/nMCBkto2BWcDE3bNvYOtq4exXN
iHh/zoMG8sRDfYYeJQoMWBGp5oSZkIWoV3M6jLN5w3hT2UvpwLJwicRiz4cmGZf2
hl+WqovEncxsju/stosDOa0QwoqN+gpGdqzTfbpV1SwnzWQRvojDQS6K6PnZz7Uy
Vxkhb2EsBdObR8iqjGep3nv4FuglCCCHxss6nxRyN1IUMPcv7i8UdOSu9sPPQ44d
vvz7VsWdrNSy7/PNB7NOSOWSnugD88ybU3x4ecxnu6qm8iS8LDjTzizKZqarX6O8
1EG9a8yrwadQu+hssma6bTqVRWuu19eTtvcBaOuRBsVQU8wPAIzqsbrvAzbzOjKp
1KLvJgqnxW1UXWZkSEegdx6MUe1hLg4uJyM4KZPDiPVWyS1xnVXOmn0oa087lvMi
YxKg9Xj5Nr4LUVGKgIjGvEHauV5IAY6KTsH3l4ZuW7wutnKPCsvewG8rJnUgl/xJ
GotJw01epA1HhMhWujmwxpdWD5CZrvKiy1odWj4OytLKNIRh1BbJjHnhalTNtJbS
D18U+fKWNHTB4mj4UC68ZwM/dS4EHQTwFZritfdcCZj2DDGFcweSHg1KwXecBL/h
WWndC9AUohor+K9U3lW74GjSFu6HuXj8EFUoEGV6XZrwr81tkJqnS6rUOAYAT4Y2
yItkRSdmMZoRj4FLbgVa6wWNl23mocJz+Em9y9OTJbhCkEOj1Fy+TRFQ/KZLcW85
MHfC3DPG5HjobXB1j8pFa9TdiXVpUZtWLyjytpElSfDfvnR2RCN/VYGD6xkJVU1H
wkwFRduDJ67l5R/5fXYwJGkrZT823VVzRglZ5lei5ZgSn3FTslZuDXtzn+x50lu1
SiyfFASGeOZRyDkY5W2wQCIJzeyxdYjEViCc/KHnuu1xa8+p60LFdVA2SmLCGSxh
bEDnyScbSZAgE2TqXSMjO097vJj88e3WMJ47cJXM3PwyOwQswWgcxbEIWW4LlwKS
t3k9YPPesSaEB86fR+2E7SbBCbKdgc4clHoOr6MoQ/2g8Rx4VzWEcWrjClyQ1n0p
/Fhn+V/ePE51Ut6wQol2oNISC3Xjzi4ewJ7r0UTLzMRkKKvzr4NuF2lN97uxApsH
WqeJcd2vHcBBGoplPXc0Nx4eZgFxFXoK33nmuXTJpYwf9wJUjMWbjyJp4yYmTWZS
vxi36Z2IhQIBm/GnOnXbSygDi3XVWhkmfY2XOhUld1qMC9ktQTjRqjxrr7NuMjZf
8djeiNGKqc3TMSyNXQKqrY2VCeVnf3YFwyrtyt6AGiJUGv7X/4er4LXZj9lu2dPM
0qJLEZMbEzXuuDNLyWM6rz9OjOuMrBlXv0UG7NVZEe9mJI3vqMPeRWjbJdGQ0f+/
JcrzNutWLqyHoousk37oE+QcOMzp8qnAm/lQ0RCEEgmompkklRjtmb8L5OmUr5RY
qOXnhQMdnnmP6PK2T6vLLf5NTT9zgcArL31CIMweRhNJfTGDy9Hes5oc/ILxJp3f
0t+/XQWWa/juYDiWfJyA/VSOlgLkJX1U6iPDFeMKNVKaPcFn5ORy4MK8QYVDQ7eL
pjlltCp+qLjTFum3coXDi9aeESiQlx1FIYxroh3GVAwwlfDb0vtjVjNPAbpUFEG1
zG86fZRG4s5cPKtXRlbZUMXDPaHEQMaloKRSbglt88J4hSI3l/m4s1eu7jivqnRS
HxJGlbM4TN0VSvtodIhwzz85JsHVwEYL47A+7ls+hrB9++9cZSSvSrxbEiuEYpxH
h7Y0FT9CjHYK/881GhurT6r+QLJzcWi1S/eOE5iJa8IdTBQNOyDMAlwbzvlg+dUV
0qdfhKDI9/o00MU2bExfcTmJFve/NpOLXDRu8Sx2yL6RtGuqcJ7UZ3eHkBm8+KWy
esFra1XMEzYWI65E3E8CZKygq69zgg1baRye2Rn6Rliyi7t4zcgnflVawsRMS+1k
gd6nI+XlIP1248ZDEwywX5bDUM8uzTR4/yuu31egJrtIm8lkqlSDv6cBkHUznIUU
AU4QCUgGRvedm0tLADpQMei71swxs5ZamH12QWwvu9tf9jD7iO3cmojlMe20qUD1
hosieslExP7AOyUzWIhnzGKJ5cq80QgfzZbBSxPBhHMjrh7/nC9suVOKVS1kLu0G
0qbwqoufXzCAOSxdPW/jCmmc9YXRvEuLYrQQvi/bP8YM3LHKFEHpKJtXjcoTTZoP
oJdcDx3J13pjw/CHhtesx07rurmc24SRRyfpB0S+HuknoYT0F//4nkuIRMT7dCbB
sBn3PzbzjdTnf/WMT3ogT5xRCxpsQFl0zT2oQxlo1EHFWCg2nhSfoRuskBGOj2K7
34qjL4ZQjwkj0sr8cWZ0zWHkNTn+Pdrs2Dct+ivSFfM4Qfjd5lncjBkvXxgj+/Mw
12QLRj1j+zJuYIUFa9SRCKPhppeKD0GK59OH4J+c5hUraij7FRYKbIAnrclrg4oV
Nh18bjQVq5R9KCsyyzbCM2N6ugWXMH54/URZSzWDWyuAXN7sFaz3S0XmiWqCT1Nw
XSO/zEB20u0rn3iL+F3lX2OTx5J3mwuBW+/rPQUpjo7uZCzG+4xDUIro+ANXz9Ad
E771D/gUnMIXGbHr7QteUqGG+s8qJWmUAc1HC+5p6pTUyGU9jwDakyhPVImIU31A
2DwkAw09O9y6tXVBWjuDByafMUJrCfUODo/3D8+/B1EBnliWukylzFVkAjTT4fug
TunUNSD5WJ053IflZZNgzywnvnyeQPol4m+HCQWH2QBEDJ+Q9H4URNnNP4OQjsmS
sJh/pMFun5XWlo5b+/H9N+RMkeY9/HZO5PnNPgk2H/JQ8WNS2te+TNJGuReP0R8M
Ca7APQTe4ZygkU6ADlF4++EbefULTkErDwbpySF5ANNNCc6z6teCyGFSqHpblVNd
vv3500p1wpLNGkYb8BqOJdB9dSqwHAwDVBvB5Llzp8Bc7CwR1G7NUIBww7uED13T
fKPJBfNcsNyfEa/w9LnVDZm2tvQvU+D0ZnuLmLgvjHNRrs62VFoHeY68SJ0gb36m
tZv91QndQPO83iAsorQwFCLm4iA7/fdxFHl8ms3U+Ibh/c+usj+4Wd0qq8gqiIH5
/LeCGh9x2P6/BIvfvDjleFIrNlgvO69Gq+10KSyeRv4Jr2MlXOV4LT/81oQJAKst
LGxY681yCX8W1LaMOVq9LmLdbO9VtXzWQ4OIfew2h++/Gpe9ur/zVFg3b/GElC52
QE6zzwimyghvIas4lVv4/36RyUvAt8iiiMt+kfM4vW0IjuRQ4C721iz/MHZXccT5
WT5BlCZXIg7PXZTZqlu8ldYVXBU9N3kTLPS8icv+Ow/w7MGLZvWtktonpJuUz7wq
x93j43makHfP9VucS+Ycs0NWFx26FtX5q+LnOV0YXDCV/+yFfX81KUHRC/EA/aj5
f6U/p2NLQ78dDyk4a77HtzF1mpf/vNX2WrJIVlPKT008NvCtP2jwN0C5SU/jx5js
9ckclIVXPMCHlqvVFXlGHfSlZ8DuPaynsRrDSnB43scIefyEBhWQied+78vP8ky9
hljdpvjRbEfkdB3+gJQowA2qq4HFcabQD2Re/RMgZxn96REJV3lxIVeeDGL/a1aC
SjhBhI2mIb7lt7sGvYt/jP/fcdcvaTRJIW+34NJxKaq/HWc7DoWnULBZKdmuf2jy
P6zc/dvD+SZzXi2RrCF2oabF7cRM5pmS6S9+RsMVKR1kB3umSwyXRoZbnW4bqPt4
3jRENYsJXIjfIi6fVgLYt/pD/JQIOywR+6uJ5TXMvwhNz3syKneMU3cdWnOSb5ZW
HeQQaKRQE933P3rAZ5823nKJkn4Ap6H9xGa02oky5guYP/lgcExH8B+SEX0k4FEK
z1svOHA1AXq5a0gZ8nKbigieEGSi1A/utdWJ6wv56wicZpmn9wVYOcVnmrlH11aD
V1Ett8pP6LH7mS4s6dG1QPUdUCK3rP14StvECsg7GMcpl1j4bLbW+3aphQ5rB/dM
K+Yu1DV4d85LlzIpWwfjnW8DS3p3MBwKwC2kaddpYouzC6S5zyZB8s8EMJbK5RjC
itTY3rjxFIEjJDH5oScTUUr6sEoW8YhAMOgsLeBFlIfY4UQlQrbPqbrB79fbxqOy
dxzPt2D91OWXKmi5MH6sHyCi8x0ww9WdxCkzphOHdxzoLHDeUG8uem3ZqaA0x7vh
pq3CQFa9HLY5jbDjEO7IObzfcg/1TU6YLm8J1zICKYYj1iNkE9SwFU2+j7OmiAMU
R+eqSxyrcmDDhIhMghTR723v2edIS9US17gIxG7Dh97zTh0YKCoQk7P6pp/FWj5k
uwnHCZi4ufk1OynKM+IBVbiGwaOQlPsTJZMpDpS7w8MfQMa5E7dfRYY0g3c4dFy8
9IPxjDWfb6G0nL/koONrb+hG26uh7PQRHkUTzQ6rlNUvY33RS1C7HYW6B92lBzlG
sLjWvAcdLxxOoGRRwleJ6gGGSJmXdbNNeD7+B8thK9VRpQxK6gy/kQxxaIR5/53T
u7Nn2OXhVQvKThG+PvLu95pelsJH9vA62A2jrhnWDKjUilpMwptNUIULyrBVZrNr
GNA8YQCTb8MNjoD9+VxFNJMCYQ/FmvGikeu7YOsBs7XSSXuGmcCzclWeTX/5CkGt
tfhjjDIMq8amMqV4NrnISuLFxLYdL4nn3JwwzwT5+boxehcBNFCSyne6mLTmnW07
0GA97FZumn4SpfxT7Hiec+CxXyFk2jO4KwTmmU21g2M0520bYpRP3oK2CUZmQYMn
rABJmHndzZyIjy+G8EB5aRRlERGUmsOjI9MXOkXfkwIKqUT/4Lx/vFEruO7Ofs9h
OWdz0jEP2r6RU84KSwmWWbtio9cdTcLecSTU/JnghDcGk0Kbnz6j+498T9obX6jY
ZW2zO52/7nOP2vFPhXqlG/d8eCji0+y8f97x0UXgkaDgq7W/9a7hr6XVAqH0tGLF
C7WzTgFaXVnzHxATjt9SNd6cLBPycUWDrUKhoNVdy09YosL/PJW0ATDAroKnreJE
s+YOkcG3ign1pM1F+zzH6J3OmuvO3FhoYpCwp5DNZT/CmewSUZ59gfQr2ldtnO5q
tfSdVQT+0HuulVQZ10kI/RzaxeexJhtXI1znR24VEV+zHWclR+ESg2GKkbg7p3Uf
U9fC3nUDqT/9oWcdYnAusHfC3dSsPfltSfhGjgMdxM7xESsj9Lh19VmNsXTkaiiR
vGLNf5z6GmyHKXAqrL6CYyBSl9TaLzki97QZe8dKPftbOW4slS1WEuNjTCPc3rGj
Elv3pOcVHhqosDNPCBcRF6iMFkSDQozpiyuJwRkOfiiyZDgvCh/f8TPgJuK3H9b3
US5Y8Y1yCqFLD2TgB2J9klgr9gBuxexSy6hjcrfddX/wOevfY8MumDGvBlEYaIS5
AuyUFt15WO8BFr1+H5dIwdz49ob5dRgr5qmkOG+/GVFrMJOJD1y1GzaltqM/H8gW
FbwBfqgZhvy8OvvWqgnKvRvKCtctrLc92NYfi9kN6M3Z3gfCkSvzfCGSCj6xyfrZ
iXvaLTyZ7d3IxWXcfGL8zN3JmijWrBjYP4/DpZk5x3ciRbXZV18kXSVrxvCcC2wC
YdVZsGdOZPv2GXNjIs0YdDjbLaBC4HHLvVobR0g/pZHxyWgUAE74vC9wmeHRk3eI
ysjPTCFmWmI5eHBVSsVvf0lqQBU+1JGuErjBPxdgahFBXKWcOO8xSRriz3dzjCoA
M0EfLZW3juUQKqOGEsJuaSYAR4jz8jMUrPj/X/IiEql+CTQHNEvyEoP6TOOOPt7V
nOfUAOr1SfSLCFf0dpOiF5ozC2B9/QXQzQTv/IhuPeOaMyk/nyCgmqQHb1JZLVTd
4fJ5UO333uF7a5ATjqt53f/ApNOmFNfAN99kCwTHBYkWGVcwrZSTD2HuERKgkl52
pL0s2d3T+wZsCPUT81NswZMBAEttc0FrIQGD5aVE4/0IWWi9o668cHAsRx5TRdNU
Cilj+F1LkWJSfLh1aTRb1KcLaVAfb4w0UPTvAHPjNJ0e8OP5u0ctjorystZStBIt
Pe8R3wpdqZ117QAIRY3TFHNc5nI2vM5SzrDbWN/1Ua3I64gMjmUZ/tV4/AGpCL9V
o3Jpavww3jOmj/EIKu9cy5t9S2fyqUghekA3zCGxdKNzCUIWOHmoBsjtj8FXCAAH
2UG7lhln9oMR2IJKwzzYLNBBn/t27OHo74TWtc4Xg3AUs3UEk5TxNcSKawyFHrVK
6+uyXSZthlPDb5MiEQdzrbw7gC2ZPNQrTwcInOHe9TsvoCyREo/5H07imuyl6AbK
cmaVFUyLJyVxZqv9j3o+EaIDmz8jjfb6nZx+5J0ggf26q7so1Jl1gDSegrfJN5DH
noMEdsiEaEkZOiRAlLcXs4Hh0jPABZhTmbVLf9I9odauv48Uf2tnTdOkCV4s/lt5
D9zhUKcDDxkveabWV6vPKAxJafmQzy+EmTIzv9Jqor6hs53OPbBphPf13hMvKOQa
p0G85XvmswKuDfn34u8H4L7nlp8XwYZLVeqNQ47Ly+3Ur2Ik+HGgzldPPTEMb6bI
6IG1QJIZuNUmM4FHszySydEw7wZebQaTA7wsTXThfWZWTYDC8+yN363QCdEqswik
cyyEKpGdYFD61Fk2z0JFU9UnHKiO+XT7dup8M5aePla6BSkwbyOwmnvjjnkNqHyt
ObOvBCYXNVe4W/bjAxq6+6Ir4ieKD3besyny9hkRgMgA32Ff3tLabFRO4wRWYrQ8
7Seo3DoYkd07ieiTjV61TM6AybHNA5pe1F19nUzA91CAfc+d1meypDPd//yuwvuu
9fM8TOKTs5FWo/qPjdIGpTevwSRUV8lsGkrzNbTH41bhJLgFYPps8le+TI+0s3O4
HV4G5Mr2kGMskplhq7HqDmNsLOROHhEboyY9I7IxMEEoeKMJLQc9+AehdUabZKeb
BgsvD7vbaVS9WqekQ/Q+rpd29TAQltRZO/PgLg7pb9pW/zwpO7A+tKbpg20yfnNT
xTrqWDPjdiHMOH262DO+5mIpg0J9FpS2V2+DIsxoTxIOQMylpOrDkldRaGEksV+4
1BNoWIcfhtP9mPXhQKhzh19S1aYSFZZNfGZ+mxOsL4YVJ8yqko4F6ivkbhM/RsVc
zmvh5uhIjb+CktUrylODl8YJvwSzciJQTlnd8qHUQVAVY+DWd9acw36rFZl2viZz
NJA0WyuYHKjFnFjRsmuLvgyxfVHzXzO2EvhG5RzBW+cIq6pcfyJlOHMNSKiwgHri
v7n2s6Mfpg9eBboeY5b8AmxKtg2qnEGW88II4xu5hAPrLQthzpG/Bo875nS8wtp6
cSj+EibYJYvBJRivIrW0GoWUxc5edGGq+l/8r/o7Yr8j35EDzONgp631usBW+0QP
Mb+c/F0rE7efZaqvAWvVUkVkqRUmFN/6TxZ1xEwrdUxgel7dvnqlk7IgthSBPHSj
lCeFxD4hmu+V/aWNLOx4kuUFhaTtSICMB3ZBrUlnFrf1wxoaclX6xiDP+Lgf/M4G
6UWmLFHAzbAs5FXkKYcHeXU13vDt0I2AkBcAEdEwD6AxueFFOkHsZP+kVj1eg0zB
dZ9xNlUVY10mksMZgMDxEUWkCvg0LS9/se15ePoo/MsbJFUvOdOvRdIHAA4xGCkQ
5rdveVgjY+L/lqJrtMga42a1nS78amAGAqtZAfF94L3fRPhJCrHijpTBmAVbGZWh
EqmpFth2D059Y1XPja9UHq9ik2yihM4WLQ95CNJ4Ln+wrInnWLFWdMji7EmyWcwz
xnNIg/6Q7R+l7Er+Q0CafqBORy6bjufl7M4d8LC77YaUfEBsKChz+N2QGmbkGqwg
qzC1dSW2dbFYqpsFT2z+YVYn9nMJTA9S+9U44pd1oSB7OeZAlqR5U/0R2DrIrw3p
tFzqRpxWpxQXPcc9FVLn7pQ3OLH9QgvxTInjbdOfUea1nZrYlEmD2Pkb6i96W55n
naikTE4hie2NeyHMuEEBe1shARdcWfUpM4blWwBCdPaLdwyh6TPlEwKWroxacPf2
9/zIt4VeS85kCJVLPGBW/ugPj1IFxDmU88sTsATMv5km0DBB5ppgQKPKB2yxfZxS
dWI7fQtMdBFXsWHfX1CRkrj6ermhXHjangOoqG95k82kdVopp/1JvFtzE0pT4Sfl
j3+u8lU8lBhX4WwKscM3YF2wEiVNBSxHoeoZzxK9GUzNxGEmpmXeqAKV6aAKxZOQ
A3PWDS9F9Mqu0Kwc5hNtch/fxqP/cruOeOOKBQtCnPKUYtm02gHnNrcEOZm4E5Nk
MS6bWbfbD/73E/x/MhVu7++hrZ7cj7NHRBYPmdLjlWkgpk00aZfVtb1KQSOQ7Z/B
Ci52po/mrbz1KhBUg6oVP8uslHFEWiXUCmhvABgFL496+LuFUwZqIHe1sncVMAJp
wsdQpsEl15hJiYVw9lcbaUzNAEBXmLM8SGO+DoRIA9Pid8FGc2GuGu0ESWNlynFR
PXTh9ygFGmBQ7XaP21QqU3LEPPpFilEpW5hzOMBFZaqLzr9COWHq79W/iULg2e0e
0wWDSwz7PvUdjYyxevVajMfl9YUNgdHi8DatvePLj1hIMYfQtoEzc7IvwNbOzDzt
7Mvan4O4OPKaEkG+h2LPqpc5RiG2sYqKLSEdvIG/UUF1BtjdDzHX8NLoyTTOZQ4S
tTZwjxhdfrvY4St7/d6QlTrksRop89rK27PKanXY6YTvL9YlGmSi7B59TFbJev4P
PsWm6wtthT9ikwkvdTl/PDnYB1bqm6jNez9SW6yriADhFW/rzAq6A4jEZGOko3b6
K6g/KBjQz9lyAfHWcltbqvfKbpmZMGMBfmGh5qHgmRPUIFH/wJiwK13b4R8BvbXq
nZAFNkERXeNw7Po+WGa/gahd6mI1H2TpYMpeyX7O9undFfg1+ChaXKQt8cYCoiTB
c9CeEfNfOhGpCpYvu5e4v1Ztde2D/ZhZbT3q44uKRQFy2k5sRiQwGiU+G9CCkBd/
eE5uJsa7DRbj+7+Q6jtd7UA8f+Dg0/DVJp3dS+O5k9t7Qo40aHklwlta9zL0fXus
dOx13UdsiAZTQ5XxoO99BA0ySZUpgwwJo1BWZ9QY9TsjC3Jpv/huBKKuU5Cwfo76
UBfNF5KQRiyvct7oPALyqh8bZNs0LLQrdH8hTOFvY/YtjdGFr8UAO0wOyouGfBus
3ws9Co+G4ZP51HltgUKvB/ACADU21q1ER5UijoiDoRHP4GVngMRx1ox5rRRz3oUb
RJnieXjdtPPp8Yy3bM18snV+ZFW7ciPnMQM5PX8C+Ttjcu17+FV+FJ62BaOhMJzy
oOf2+/YrsGnAYN+WL2kLDT+fBikb1uqNEmxDlhnmFkenBPPzJ1FMbOnM/thgLAZ0
tsDmibKoMCqGmSy5xBOAtnVUFjheGfDk/9KOqW4VYP13aJw9hnn12J35Y1qcEOXd
bEjsmLq81HjAQExNIeU9/oNMhLtJMnuxelfqNKesmQ/vNc2wJNRM0zL6RmRemwHV
rF/V7qBNspB7msqDERWP0KpZFwNp5m+l8Tnrcs9TFdPChFRgwWMf6HeDlXLeY4+/
ON7Md9rQfgIVQwAayyOqH0hH1NNjN/linoxF6RQ4kn/z7+cxyYboa0p8e7EE8s4J
xt9iFijeWH+I/MUQH72zcgXTpaA1YGoNxEU1X1zO+uPJ4mYVZ/NfVBT/byL/8SLR
umyrKPp92A/xgwTmvOqgPKUBg6LBKxRJk9TmkyOnzIVRiji3O1x13kFdtR9TNUlM
SkPR7ogGqp2A+f1JzyZpOTqtd99pJ16503lpqlr11oDsNnX9nh166Pd+b8hr7zrS
PFimQmKD4vnTNVkPu6NsLqucs1g3ZyC4th3wy1dIuRjOJze8MEh9EAf4Ev5d+WyX
DhAnUt3dlC+1oUlDEIUF3sDMFGq0OAnI3+Pep3d6OZPvnLt9GV1VNNCtmJ3mIHcg
aXi+v+NtIiMQS2vC23pwTkfWcxFSw5oi7SfGhB0EVkGDO8Wuw/XkN0jW+G+eJneZ
HceEYxd14QSqKuw+0qcWV6JtcSDjnSemwX4TXQv4vBpRxHomhcY4snithU1en/or
BPpcGozrJSxewQToGbKdWfn92VkW5SimWtrCSN194Ug9JFIINRghkkkEmbhD7jZq
cUAFoNa00K98oA+a41r7JkLmIJf5D/ubq0Z4TWVn0xz/1GA1LbBpuqocyIzg592T
GVX8aui0ZHYjbjl2T6+t2LOThFWuaY4Tggw7+EE9g6z+PDWf47HbSdFQVZ/gQVpF
J/HMvRMGyEMDGS5AjeqJGOEkvfU3bmlmhLImndzo2wDM3daZhN8rXrTlIts7TKnR
am0pXjnhGiAueFeS3Z0qnt3jO5wU09qL6P14hhCwqde2ltzvVpDdFsqVUaxDrzLf
9QiMDYDywGAjGu4PS2FwPjfjolvqtJrZcP06VLRPf76jkH6PRoKRgaR+5k6T6g8A
pPzZUvSMWWvr5wn/1kbjTyHy8fFo8001WOnZ5FTNnz+t1/7xcGqQMHK6Q0yHrL1e
jkBRIPdvuADzkfKvkM+tWB0kIJ3VMSiMrWJA1tnUpY3rNAFsjOwHXnSw989u4emQ
IdslwqkdC27Eb6qFPQmXD9MSzLQSLiIJEGJEtuPkAeGOciY2yaAu7Bf82dPiVufP
melTh5RYtL4Nvxq4e83juhlJ3JAN2pXbwAAh6EBDJM/o2tiOm8HiQmMzdETFjxsh
pZoRZJ9zBpbDxwUUybm4xi2Q9VBYdbZBB+0WjiDtJR1Ix4oPO7KrHsInXtsAmrEo
OHJyT1a9LcLpOBQFrz92QWfz5AArvklCkoCpdJlQOn5e+0dMS54ayGY62aItqPmQ
BVd+et9c9Sn137gUoYgvBriCQ59tfLJO+wp3EMhvxYN8l1hWIq1wrW/OXahRp7lu
elzAfdmtZsmdd2CQaSgvNRpRMqwpxlSyDlcu556VI08gE0skLVrqvQdiNiRkdad9
t7NRSTDKRU3aU5k9MVoy7R/Vflw9rHoiItXIQPC6pLDYQIFwI9meLeejsdXy/8Zk
nvHIxvuKLbFpz8H+bGn0mggVdZmMso3f52nZbtq0oWHQpwC0Dkh/xGMzo7NpoDxt
vSffacYux1Y1z5uHP0gmcOLT60E41osoy0ON6Q2jXK96x38/csE1soPmIrT+0/9Y
24GG/pEUWum0C37WRcq4elVynDX7JNRUHxz6TOWRie1EHm2T3KQonTg5YoaIkFx1
qv7i1nghDv6AlyJg6b7eDPXTYEFfS5WgHwdl8cXXzyCH4p+ed4pIx/Qgov2HoqB2
4FiPja4BGTQIoWJ+9qR3FKwa+itkmgJtCidsood766mtgdL8OolLQN9uPXT9l4ey
iFSFKDxFcuPC45EG8Hoq/pNmdmvyUjNQJ6mZAXXgLWpBka73CC5LliuDeW6DKFNp
v0EI2lnydwkYKWjKLOamIg2KIj3JiEaO52rEkJO6OCD17dvIqL31pVMuMgBJLgQD
qQI29LyDs1E/llqk7UA2cW1OEbxpMd7ak6oMqopY1wMDDxvKU11TrUp+k3xcoeI8
TBorW5tTGdeaFzPNWlERP+5yZ9DgCmpd9SlHWXAQycO3AihO2ETvsMS06CNXbMGe
BDwHIwdxDwAt8iGGYDBycnAuB9qzg8hcQIaqOopCZzpkn97gZnhgHU8ukApuFgbz
4PhlbvG4SmzL5VVRvVzBkqTfs8itcU8VA/u3rn3n3g9fhlau2ein7L55oFvO9s2V
GgrebqO7pDWteGlATOHg5aYleg6w+JTGMnwyC7FEzjPHCM3rIZnMEnX9Q8V/6/Ei
cq23z7sRUhNQoMklUvjYJKVMo/pj3jIcXG9wkirn1ddgzU533fuN4iupywMfJbtx
NrGCEwXnJjMupc1iwFsnqKdXAvb70Z7COfH3v+ZeOiA0NKMsMe+10JKPFK404mTZ
ZYrDSQFb74YPUgRhV7q2GjzzSBUprWcXIh5Vgl+8CGj4QT815eB94HKWuzr4LtuX
6G5EtZJ5qBlRDzW3hPzV6NK16gNKUek5rcgSungTM/k+hM8ULfu5lxiwYGlqQeXm
sg9n0wcvF46GbJDCBixw8TCDy+FwJq53cZ5LyqqDeFiI5icevYLak799+MAxOnQD
IbebbPdjXV3ESGb/PtK5aTf6pj2genx2F256gKMWlRn4wL4pmb7h1Ly1ByuKtoX7
L+aLGD4Vzw4oCNWczl2uWE2mGCEXf/C0BgmU7LG9Lxazu3zxjOvO1Awtc6k0MwbZ
o1D7PsldlYf4/8muIMYsJlRQv7KoGGp7h3BjOp6Llc9vfsaSp1ABDvAQxD9rtj7j
kCYzqhSHEjNC2C89ePHVfPuV9xv4VfVkybUqwnmPGd20fqNhdZaCfotyU7rWv5/M
/XiC38QEe+0C45bnMnZMjOCZfnRNVQ3CRnqevrWzRsjjfYLyGZCGdkyLqFQrEBIX
RGyoRtSm84EnblaQqEtpjHDq0ozds1SDVIjZq2nNnWvELCwB96TNjZaqKjQq62SG
7GJZ6EVjkN/W2u/h4rk89VxPNYM1u9fkxOkySTfsFLrR8McepEQkixLz06Ypd2P0
y705hCzVFRNGyKt2DCuhn+SRql6lqbdnJOxBN80budHezm6MZltiZuylbbR7yRzC
GivA30xx1C+523r58fIvIoRfcop/TYkfg1aMlaVTXSzOj7RWp4YKQNkAU1qxuPLr
5yEOQI5vbZ21PZkMvDG4dCeuJcn6KKDH+kKo/m3srhAhrZgDlcW7iDbPe7uztoUw
RlV3A/NoZ3S/UhJB1D4XwWYo1dHKyQ2TeVtUbqjUv/wuh4563r/XDkkV9Edr/pN6
KOmqYKsOd6AYG0P8hEqZHgpVSk5jLdpCfeo0qSsI1IyLTuWhkAEkyzvK0uWMpw0h
kir1EoObZkpn2yeawq33mvVatGMetSoHrtC2dAVkV9Et6mO+OVk0WgMfcT8nAsYz
bVtlU9X4OUnykCeywZtltVik66/7ENkip++0j3VUPO5V2a+6rxa1xQfzjsw4XEig
Wk4GUgPF18PuD2glvqMoeFhAOoTCBAgrOZkPIW/8d8x41zZXseyabAQZlAwJZYEv
1Wwq4RKKSOahjIcy8z9yomXzQKJvjHxLP37iqWV2G7gft3r2F/VAH9bnv5Fv96HA
52SmZY6VPE+KO9moOjf0Gon33oPS4WDFGJ2JtAkdvygvoUSbUzzxKnPF+9dL+pQT
YR7rj2p+URBTt0Css/ZB03cGqNniF85WgtPPJZQB43ESsAM/x9XmRRpv3hApjeHj
pH+Vprp9nlvWuEwgZqWTtwx74o6NrKEduZJXqQtWjZ3NhQWNWEgV5nwheNdzqPKi
PEGY9POykxfh+hpCexrmscekrnbzZCjjbrYKdqygx3rErlkXsiOcnYJiIYHW5Y+L
JfnnfeXSoWnmpc6HbIW9XDmqpwrN8osACAy2DqkhEYc/j+UudoUOx8IMZiDhHvIJ
BK8Xg8FQVyXWb06owTJz6UkGnDITtzApKp2VRrGzsxIf2Gu/1A7kV9kCuvpQW2Se
5nb5M4XwOXAa8ucCtX2SOxXpZb9yHM2+Kzb4G9c1E3OYeTj1BtSoczc1iZqq2BMU
m/myM5HdCvpbNUzLfSjG/odOpCqxNE3Fh425/EoBf+td9uD9D/X8HyEAOC9W0/A+
TJaqGzgi5kwlCotHeCfqyZWlMi6SCl3hOAQCbHf6bJ05H2nRLBfjvjaJ2HZWjIdS
wcHS/YLSsmxUmemPVRANaBFbYxmnsMsur22rJJFZviAPnrNMi24xzSLbBOZDfRvx
/uBDwBGnBP9HJIid4FFJ5d1Ab0tiJ0hVdk6f/xZSj7t8f1pJnlev4FLnziyXzFcv
8z1QEh17J/muwpmC81OyewWbwiOvVHB3z6QX7V+1FUtqqbWYfpI2Tat08PIfpCW4
ERvrAkvRzewI8FvMf9ZDORCdADATjobG1FEeB6GChoXcObOIG/LDhGUCfvnL1BwQ
jUKo2v1kiUlEKnfW63nWGAnux2cnFY77r/wgoNDKmI8fHJVfNv1pskOgc8bOHBqw
KZb1vU8Fy5759STWUrsAU4qIt1urZdigE7RCeTE2kj0U0J3pWEgP/70sLM58C2sR
E0YZsiMCaWRb0loeBcSRQvke+uSML/Oeljwtw0+xooRK5y0tWxyE815K5g29J7am
iGDsJ3IlDxUW0WkLPy/Mg7ooAf2C6diwNk8R2ipfEKjx89XT2juSxcnZG+fTF9nB
Zv7hpZc/+EMKbIn0mMylhAXHOB41v/rbKY4LzLHjP0q6MET+jJBWFGwVl9m+XgrE
4R4UOiJrd2OAwCYrOaFIrjo//DWgS4ULUv/55gg0Jw4Ac5nij3X3jHHaNmvmdL/i
tKZLckBvHytR8TzhxqzZxE0KVWqmp4yqDx+XIf0GyDRmOM09fxA4OPt1DNe4Xx+x
WYsXiu00tb1zts4vpc74xC7cGzxzCYQzbMNFooXKjeyC/kDdCZAkcSoQ52TlSXGk
eNGIJ52cGc5LD2MaMzv0WjgND179NRmscurhLo34HF6ucnZgwEjsIAni5AtRUR17
ezo9WVKhQbFLZu8GFvwuerfEjRwJlMDi6TjoZet4bolRraPgP8v1nzW/WCO6M9+l
Wy2dJM6j4lxHZlfV65idTp4PXd2KOqKamjcZ+JVIL6kFC/TAR27nAuaj8RhlZD3l
x7yVDrDrjiJ74+yoop29neDJbnR2utOMQcW+nrEgmym/WNBarGpLOeUI6sL8lfL3
9NVFZeKrTaxpGpcUamrAisO+O0Z82zc++n9M07OsrJYIsCOHvHySJWdjRxhJPemp
PcDVT96k30AYtDhC8KZxAcRnIvxNmVu/EH+xVRq9iok2OREDk/I5y9aPaIsAucT0
o86IuVLQFEq61rWtbLCmjJKreXiVxDyslqpwjR3EW9car/CxbNSB81ZDY0D0lRqi
bj2zkYvnPbFtrrJsDObrF5cJtCCOCelDcbHBcqQjgNDbIP9ql7cat0yvNiL65zgm
92mbVAp8mdTs98XZc+6E6zDj7UPxHr6VLoZkC+BbxhJ9JqrLuPhTc1W9Or14wtyZ
fPRHV6kBRP3pB4LlATBLuUkMPr1XMsskxVmcYyJ9yMnoglcMmPcvSDouKL/NXGpA
aQwB4VBTMTXuyf/8zkZo68RiPuo6a0bRMcuTDS9g/pbNVGn+ltJgwgYgx0nsLWY4
TjP/Uaodf5xboepqbQWZVWJy32tMJiMmi2z7kKL9gCQ7zKiB2f7r31boRVNMLozg
aSyqb5khFIi6LRt/Abu2gak9Uonht4DpPDnqMmdIqjy4zWlSOMvipgDnbsXibxWM
Ad8LLTG/SHp1o7wZgj7hrLhCjJ/WnATIkMaidrKkLzz/RJw7sWzGmgRZREgRimVl
T39hMzwSXF7rBnATGdGulHz6Bg6EOxRtNeDrFnWDmh4y642n/4yCuPobImsd4lqq
nR+qwLbae8oBgKVqPp6mfu1AHO4Lr/x/CZbdswVHaYd0xmkR5SUpKkC4fgCFcLSw
0RP4+WKr3F6h8ou7H3RlaaSYWPDARX99EZyQoYV9sQ9AStaFkGbzpyiKIeiLcvB4
xdyXer393utOd19e93CM2lahiDpD7q5xDzdf7h2aoPRrupZGDPPeTJo2L38miM2M
gU7CnwUFH1bkB7X3ZcipkaJ8UgbGFZ2PA6jHjv1sTj3/sSvME8xcA+tm5kC9Q9+y
XnKXthK/OgLFDVKpdkugyjCq3zEdvPb7cN9JYmOHs7z48bJ/re1FlV5awEgXzSdE
hs5yxxVTo3fyGQ4JgmuCO1fSRlwu6ZT8BWw7TmzzsgeD0dpXGcMvFmJtFwXacC7g
KTAgFyPh1F4Kmb9+8uqyvkDTZliw2DZ+0xO5uMnROeob2nWkukaWEC3pOgEOfNSI
O69VsxBom5mBwxA1R8Ur3HsAiU2osxz/X8lMULsqOIHdPFtUCHh1Ob+MEnWkxDE7
pSooY3nna89w6LTcywhm7VWCdX7lxpM0WhUM/xiiEfvU18XTWPuOr5Sf8RbwuCt3
jnegpSspeQN02eLBK6SanTPqs9b7exeE587MfNMiwQYvkitCswr8ic7Ry8FJnME+
uxT/BFz3YtCo+82wMZ07a9SmiWucsUxENbfMTKSsWSPL7zF/KokgfIZrcrecpXSy
InJFzUlHWG0ndmHNz7BBhh2wQ5tqqx96k6fZIqwoiJpf+cc/NpvCDvzhk81GnOv4
R3f2+piY+Pf7NydPqBKQcUmrVh1bez/uqXUktKIGYUD8eb0ZGlxDvpDUUg2/sb5y
IBDADqeZi3e7+zLAIsxflqJQ6HPc/eDNs0mxBItMHzhVBD6wrK6ykgI74l0EeU44
Wc4RxGcTVyajp3ogTz7A8voB9+JJtTNEYyW1WFhH+NK2xDv/gb7Np/cesvCU2Xcu
XSLQ13xYcVEzMcS9THeFuaIhuHI454G6Gl68AV8aEgQNvUeT3ZJ3a9w/Shd36+jD
KH+wsfvjiXuDcXtCeoA8FAWVHbxYO6+VpBe0wYXfNUx7TjLPkrH2Qh2sYmQMlEHa
oiSho/1ndZRMVgolifwjVqBlarspChLh12oniXCFVEIEqsBhl44iQ0OJwOUHujfZ
/FbpnomQCmBOQDL79m0gBVa74BGkmqGd3QsYpJ8mIyXBwI6Sbm9z3iM4mAGVd06K
GQLmD1GRY9X8CnoKJLN3cHqvzH0dET5YzX91VjJMnD9nBc34zCWVLo8UWfV0Dp2d
xFBoPvF59ADOn/IVuuLi8dHoScTC74jsbeGKochhOq5FXSsXeBw2MfSmT2BbVtdQ
Hdf0tHXM6LtZJwUW3Kk8arDxRKYzxAVYyBzS+BUrQFXj9bvOWPR9/VTf+derKMnV
BnQY0jqs8Fp29IxpFTFocBhuXdg/yKQEMQVO+Jf2T8qz+qhYhUyXDR2jx8o9p34V
mPnG0qlYoC4+A0MV2qknpzpUc+E+7/q0oQcaDimAJqbl2Gk13CYmQf6TT09ItOsN
19Zc1ZsB/QlOvXGK0Pep4JOv13H+/5B2zwBPiEsZx6LohVBRwCKtRXyszSfaYNJp
7lpzXSP4OzGreYeOHt3OJ4qnDXevy+okJJMTgYan017YxsYl3xk08UEOi0wgaopA
G95iAJGZi3VB0iIbg+ihqziqTPB1zT8I9bMHVYJNWUSnGEg0fCPCeqpp294GdVVa
lWD0T9aDDx8K382fZChUk5Csxr1bEMWCYKq72x8Ee0itkfkqo7bVmo2Sy0rh+0BK
S6Zb55INw0v6aHJJYINCjEN40fhUj/FTjPhL7i7DDMO+xmqExTCRVtxQPAH9ESxi
DExV/yC30kgkIK6YMTg+csX7k36xisnAG3SC5mQaWuHIpUtDaZ2oBeKMtpxkxqxi
hq6Taf8YIOJ6LjZdHaeTaokE/PSX7ztHKjX8G/0/gVqc5QoR6AbKAysCwuxWY+HZ
AETNTlb/e3jwQRIH9N8vArXYubPGp3I+f3yqf0zMQhXn44myaGsjWc7M0/9wRPeT
/j9PSGrL6eXJXQr7K/os7R7xXMpRjd5HYja8p9y3Xb6irSMnXsdrTjamo+Dbgdx7
HB/livkC1rOHl5KKoen7wBYLMvpV094Tgdpc77ocGi/0lvcDWNzilvHCDf5XvaRJ
hhob7gdpPD7hffImu0WKgKiyjY9m7bxCCCz8Lesl3tS0KElRfpjYdzAE6k9aeRlD
1kS8QbIkB1VOHrapImyB9in8FSI3iIUMw3mADjMld4mUvD7OP+tudBy9KvOLLITX
iD0QFr5kSrc/qr7cfMxuu2PyxLobJxgVZlavxva8MnZqvDDmUQghQCw32yUQdPsn
EL694gXKyvhzVzGnw6/QfaAjk5UsOAsva2atHii0T0uO+PAER//AO7eFqnsNd6ub
9L6fffsv1aft4RiHzJEtYVqtEscF/4KRa0EpSXcOENfG4/2Ky7jy9ZYqsZCWc/EH
5AkyLnTI9l2EkHrZr1nIPsDSWwdEdK7AO84EXpdDx539DAHTlNa4Jg9+vP5uU5Uk
jBEAnCz0jyR0wr+TjQT6TFnwR6rbBIUqcX0hGorohJLcnrL6S1J1paCAhrhlcEX8
5HGr3T9He70qYfLGWDZKISNDxQqvEfibgSt5h2h8+ULc3QTQDhR3ekXeR/xN6jzE
xD8FL7u5ngnjwSNgrPdNxIGpPqujCxZPWJZ5WpsVki0NYx61yFDaRqSfAx5YxDtN
BfZxZGecI0MH/n0MvRtm59JhtAmSYjLGr/6x4oTFL7g2MFMXy1BHFt+BhxERZmvI
VHD7l8kCrnOSpcBE2R28hfFtb4rXa36DRAAlsh4RcT93nI91LVkblcVlbL+PyvdD
760InPqPjaufQ5jlQmQJAXwLfatiwUZuoFwJr02141LuSsjriQoRFCP9P+h/GjpQ
JH2+VJDMVfTWGSjQE4xhyYluhz9K8xj7MFsAbHCHO5qb994eUufLBRvCmYTXV/OB
eMS0/2zhxJMSDh+Rch9TJPco6CW6LtGr/F7bZH1RFWZdLlWIvtK5y1vPlDhOsTCF
TlPCQFXooEn/VbdvkYtwfoY7bpoFIwIg0d7wnyEMQGxhBU68moeCcrzc/OA2y1ln
4Y9ryV8M08FlL6FEoSnSJ9sHk6Dsdd6UDABRs+B3caihO5beTcQ9qUPDXGr/NBsH
pqKONtKrUjkgh7X1pQM2SMvVn6kGh28Kw9+8hhjW2vP9RLY7+aiZmR0CahWXGlxb
iw0NXvedK9VxLk1RGGnSh4LmmWpavFDPe6ldulmCVM7y+EoHhxykjesxFZgCrO37
4BXMP35tfA4McFiU5+LJRKPRSwsGmJ8C6QEmXTcFGLjfXskqPCYL5oLsA53W5Xh+
r1mbaGAu3toHHkyG6xDEnA9gWKIDmHZwv96birUWudwGYUY+99XDsBod/T2rKgEZ
W2k3uShppl9nbS084dbP4SBJsi8vvOIgECNuaoiyLfb5Pt+vb00WTL+z3/Nzd+nd
XJqxY1hh6+RKzH++mg0Ib30+nkQFINI0luIgQ/pbATO6B/Q5r+ARkkXnfg52XDit
p8L5bTgi175ElXk3XhhenyoWhCWuJETtEgr8WH+nk/a8pYi4IK8PUYeqMa8j/4vy
IA07nSZ1UF7upS7uOv6Q0pNY1pyITDIbvUs0caJzXmPQTpziOM57/8naaA2ypAaU
RhEC1Vb6hl5NoKmxdFsSU9JuTmbXMRyHIGFbRssWhUacOIPyeYO3YByqKCBMZUhp
DwVpkd20zVih7eiP9JAx4iRXai2k60sI7wU6S8RMEBaPJvIwDd2/RSLN357QnNFk
KQCTtn+J1ONh4k98pfBtagw0h2j8xG0Vp3Cjyl96vnCGDcnDn0yDF4LOVGUxm16Y
iy6G9lfEFRzfbK0GA8FRW6NErqsJ8SAbpUVqLUAemEdfegfcD9ikoHGgSvrF05MV
I8j8mGuRFr624GF8PVSc3txOnWgtnVi6za8DmzFVnCiY5cR0ITXOhLP+AOuPTwWf
JcHPURHJnjFT/cO7BmpumX4GwR0IWVJu/FtGf+V8+igQiRNttkpEQe4nvZg7JtsB
pK/gPwfwgFAZ4zC1YWoz8orLfLFt0PQEOnco88k1AOqMQEoLaLMUdnLC7+cpHJgS
zSlCYg4zUXHoDL7LbGNXND2hteEuAXyu7bdjTjFDzxkkZlrqjOW4TFIa1jqTpB3g
E5Nc/tiy58+T+rR8642YlAjIlnc1Nh6rglpelZfZSpH7w9QFcMibsluo71/9m505
/UlUYDYINDDkpad6YJTpwvlqFcxok+s4c/5YHhmzWnJvzs5rRDUB/gLD9vgbUIZL
+esR6FGMCT0Udh9i7CgUCIMtT1zAybUXe0i1I/hUKQTXvv1PP/G46luqbEabRu/V
Y29XOhMPFvKecG62yF4dAB4sIzcUOOPyU2cbETe6xxAbqCyYDmRIdj1R2rwTmzhw
D2hNK9L8D5hOJaXAAnTfYNIj6kd/whNN2+G5MiRNNjnFkrR0eArFsnqZRUV/zCTW
f7/d5hF4v3jnU8loGhYz1KfXAZtFYYJwrvJ3x4Sz/YEdiuMAUZqREUcGlj6CJ9fT
f5XaqfQ4NNwj5l5VNQaY12qZPDbp5/ZY9JFFgRliynFtRwZF+qBPq88DD6uhzQrg
iKkKS96TAAYIj4OuOssquTnc/Q2TqDzrv+cmglKKcB9e3BrlyhJIRdNSunP0ERa+
oD90QaXsNJKmBkjGqxIHRufX98/YwGLEV2IOkZQfLuAjCf8+ZPKM7snJrvrZGhDy
NKiD8y3nN8eGXveLZ86NcS7fQVspbD1ipp8AqEHmCNt0lPOn4mUCK/xb6XN1ze66
3MqB3rS68oxlbPT9fyyJmfw2uGua0XI2FbK8MktDLFc+0YCbl7f34HSwkDE8Jga0
eyrbIEEfuyInP+MzTKAb9gC/k2Ey2L+kY83YHcUgUN3k9kpq2+5z1Oqkm5cKvjCa
Ssw8AWnWsXfFyw/Kh6aSZ5B5N2yvReYcIEHBRQHP592Muq2XSjnf2ITKS+nhPfDv
3R+CY6rKrX1/wn2jSVIeLsVj3UkMMHeSlmVOt3ABi74NVSlCsSMjhlPyc6CjWzHP
uJGRssV7kAebkW9BPHiA3uMByZc31sA9a390mq27XhBrm/+AJmRPLbHdgzNlhoW0
RDB8kdT3EsbeFrz8qCsPGBV3oE+gP0r9yd1D/T47x04vcr5ec2RVge5md1Uvy3/r
sv5DW89/CC5oLBhjjqmkt/MH+tUnwgFagCewf4DzzcghjY85ArEzFAY6AY3mm188
UnOuvZYtMIUzx/SVTA/lETexHERtPLcMqBQE8sDQYJ3SskSLgxVmy2r8Umk9Ybrz
51C/a2YmiL+zchr9CjkRFXQaiGKMWFjRHwAeXslp1sJHIKrePaZizX0TEyt0qLbF
PGA7ZGGA5zR00Vun50r6f2hzgP+K1kV9ku6IbINsX2RLQd9oe+wLRb5UPqPITUho
F+SoBE6no98YeSseJ4OmWLK5MshoG7Cx4z1Z8i8ViwYnY8Sww43UfVNOg8EciDH4
3CKDSovwf/yc2XCR27g45QNxamYI6XA4oKZJH2hVNygNFtUEsts5TEXmeQR3+Yam
z7xBeZ7LSx3aFASFbIpDYmeEXNVheIQwP9/S2Xh8YMfr5st6E/dO3wk3aWBi+mP/
rbF0NF8ptVaaasqypy/rcKMf6NNmprnNEfLioo4rrwlG3qLgHzs2OTsDC8RHQbKw
2Ih2Hy7aCZGXcsQCmPK6fBNu+hj+TrYWH7h3Zx82iMMZCpqYcNQMmyoWBKjpiRHZ
wkTuHUG6f++Bu6gBas16dl2gsP287KxZ2pO/aRxq7j7OflWsISk4UZScPbyyEJod
UHPvzfFE/IUTJZ8JDG1S8iI4OURs6mRe49QcB8J50IDOyFt2mDOyP6A0NE1AoZ5I
bNtMm/NKPp/OrCuOXuf0xaciJ78yoz4c++ysBzBmrQRfhen5UCNzPh93n2ZPU1nJ
2BN0hNbqfYXLfm4YQW8FmwyNLqMI2fCsyp5kAPEBE9bC3pHhjG3DpSVfRYFqVCsL
fZc+PZdTIBlGWXfdAMLflDiqZs21/cEsTjAIVj9fhUt6BideJQjab/WKSPUgUBCZ
EpNQuogqyAfd8fCse1f294VgNKLYhjAgeDViYJsEGRdk5etlsdhpBvTTH+Tv+FME
73NgkO/9gJTyykA0ub6KIhk3/Bok+j7PWQQ7W2Eb6HkTms9oyCsZeEFRVv3XrxNj
328QrF0gzu9NsSAfECZS5cTmCg10724T/Dvp8ERCoZHudB0+G4ylnBZZTFHvt8zk
LYg5I9mfzh5SdsPUEojq2YRIVfYwwmfDTJupJ63+Oyau+me+2fjBz0Wv3CmCGySQ
54tFCm2NdaVB88zJMoT2RfShXnmVfyYglZkRwFlATCh8tP9a2boHK5kxkSJC/KFG
mynntoT1UZmCwG1/KQM8rdl6tgG75GLXSMmtDk70uJ2Ae4WL6aG+075G963Bb+/K
h0Eq74iFSZ8losdZIf9EQgPi49BOjx9skQ/0ltEGalXo2tKInZHRm72MP/gM2tPT
bPyM+pYEoamjcFuYLtMwPi8Rd93DSCR26j/34aJrWSX3dGQiAfA3ZNppkmIqocSp
yYWyRisGaVJ/tHIsoOoMYu45dbZkSUqVmojA5LOWdgM1/I+8Zj6EgY6zhfZbiyyp
sz4ffdBvO2+bzYFQWfAHf32w0pSZHdT2DLLyP2k2FiImg3Odw0LafFGEpsl194dX
kzlbflM9HPXn1MG7ff8lP7x+E1kf2xLFomR8D4hev9peL7M2neXxF/ac2bHcI9Hq
fO7XcWmXeKCkGPG/dQxEeITL9ouuTB2E7Bq4qpg7zVGD84nzDhhzj3fV48fVS7Ml
9hMpCoOmofGg/XGrHvhjFm/b3OJSDA0ngg/pzQ0yOTubNOj7jso/v/+WOumAsQCH
t3cVpdqxzH3u4zULtoBQtA/iW9Am58SqS193NTETEwGgqm0kLRc0IsbpBfKEnxSx
h2dBllxPWfkFwqB6ESNXkdG33ZSa9fNFZkmDN7U1+wX2kg2pOaEY0Dde3NiRzWAB
QSQ+KzV8TrTa8cJ9KIRktIDQAJy1/YdPBXTPRkvwE8S35sxdzMo0buFctiyCLdBK
Q1ioBhY4ZfvhVRB3ttUX2gsXSr2D6xJTsR78zD4XW2RpAMgZxdu87NN+hYncYcmM
+22RNbk0QOLR4BKUUA2s/VNF/CEOUQxuG5VOaS+ghxJbTpgn+X5EHrxBRR4Tf1u8
6pW47PW0xNRjr+N/RtxYVqpWC9dNkUzwLtSqI4twAxm3H2L5/7EkaRX8OUqiZX+i
zO+2iF8BKjrRGBfYqWgnCOAEbGnZhqUsn44pj4Y8TSMBnWnYsEEqNSEPuKxRt0q7
UEZ5CQucDfaVC+UIBqKTsTUUcSinGumH9k774dRF6HZAanvSiAvZ9jKPgc26QQXk
gmU+Cqmgg53FOuzdLtYQA6EcbZECQn8XzeBg4hNwyxbCIw62Y29JCiM5YTpO2pmY
3dM+VrNT9YZcez9ceE/qi+FCHx+PHt6UO9YN2A68g8CVMQ6HgfGNrFmbobEMKFqy
2VBGWKl3F8J18REkAkIkd/0vwaSqHKVeBx2bzSBpu3OBod3AHXftn/2MUtAXmPf6
Eog0mEnE6UsLhxx+97xSmJPHIAWzjSDdQfK9FEug3Eihu5VDZV5hYz6b91yQg0VH
fVVfPCt3tnJ4gQh/nhsPm99edPVoaPQPlxOyRcfbaikMsVI6Mf72RQz6tr9tc36x
SN8FTrtrCPV5m5BnHPv9TsmIVqaVZKzPvsuyOrc9GfzYWNrqUf46kkfatoujbej2
vIJwURynoH+U8/+qlfwco9aunN7GoJ78ycck+mP9dM3+30r8TD28j05999RAQ6yB
DLXseYvhW+FSZnxscE7DaPBfNK1t5iqjESg/K8niYOQXLTh0RJTkSNooxXqAgWcz
CTQiccghKn+C2h2onse67piBXptYqh858HvdrMMlkY/WD+nCBo2TQZ1Uz9/pBIhO
Ud5vKvfKrm0U3b6gsJ5EAJE5AA9wFweT74IFEOK29ycLVJuQBIQal3zmgXFOemsC
O8xDu4NfCzjJ67JiM+BcsQtpVePDwo+IN2lImvDuzywA6xkaB0fbKFaW6lCdTWyO
dW0l9LS7+xfnsK/6Dbex5wiWWmTIexvXr4IaE8qxSiqtp4GyuV94btSTSxr2Cg2b
pCNeuV5qF+H4JIWK/pSPAkuhK29AWUMSdjQronCOSPYlGG1YgAU/eX9r7+Sk8QPX
NvNXHurMGCVpWoE9ZecP5mOBVgdIkZsQEhocHCTFfV4VNceXZjI7WHQiKmLnkj25
Pfeqy0lhuoIQoabVbmCE/cVfrSP74Rk6mcNco7R1mcRnnh0uzpxHVZiH7njYVOZg
9RaP6mvV7Gr1zWBSixlgG1HOqJhMjizA5skZeljqIbsyIctY9JoBXwv9kMeD7BjN
Mi4SA/ve9AH4jwFUZs2SdzTt3tF+aNmUWQjAh6zXvR8Wz5ahwfLB0eGMMyqfOWB8
C0QBDByWHJosdlpA+ZjgOLzfHRxzAinDbfzFmbAEsTJkf1LzeCurUyyJnmzwh2DC
eBwT87td6zRYiY10YWSXBnw4gnnbH0D9ii0SwU4EWoXjw03cIoN6BsVyKji0Q/i6
PW+xxirRzR+Tf8t4M18EpFNBRWSjOYuSnQ4tQQ5sFSFkWV/8V3mdQlrmr+bd7i81
Q8kNzapYuWD1HGHiqV+Ly9kZXiiGZxc8M8kInbFYMyH5e1tS4uY67eKbuLVDl6VL
2Xk4DcuVe8PotcFt4k0hSSiBT742R6uwW/7zIuTxx6B2V+XE80JCagmhr2oxubns
yocHgPvfxoG7XbAY5VHG/W0n3saNRHwtMO8Ix/hjRKOGvSSO0t1hWPVeCs6yxZlh
3dDuPOx7smnsp3p9F6RLEEPbjCdKlAhqBGdvW9epUHSJPpRKyEg7DotdwyMMyAJk
UkADj76I7gRchzuaBijDY8lfv4iauakn06bb4znzUqhqYThEGF5vaEOnMNd1M6Xc
wauR/CU2Go2+mq16KLYmSf6PAcOrLHOoWQQeOBOji788WJJoxUTeffQADVfBDy3P
ciDUyh+dncPrUJyDl0H4pxO93ka72xwYep6Kq+GsV3QeGB8vrZD3mihOhNfmrbi0
BMnJhA+aCvU7iZ+0E2IyvOOscVy8nqKq5IVNI1zoiychI138uwFjgtZyT7j8e4Ml
tTPQb6otSKUiWj4cVvPGyRQ82yS0kSPaJz+PFEkYQhZOQc1H0KcrQYWevqjgUPNi
Jcg52egUquIqDTT6R3EfYTaHFVETJiRTob6o+3PRNCdir+3zGOYlVls5j3WHFkxd
ZDty2cRnArvRfF4XceGwpJD7xpaDTq3c6VybhvpXR6v4lAUAc+PQJ/w9EeOf1d9o
bzlE5d/SV5cGdatskJUp6qGdHGMg6t7tttk6C+B4g3qrsl5WM6VIdtEVOh/dMpu8
e6tSUg6ojAblyJhvemFaj9Ak1h+xQWEhDC4AgPZRXxOAgocYGu8WUf5iRdakz1NG
6GMofXNpR+E6a7MlW1UyLsNxt5zcpEkeHoEm6a4DLFrdLFHEQLbH3phLtPzeI4lX
+cCwoVLmCyrUPHr5PuO3kk460XQWZrG7+anXcJ0V/+9xu8afhAU+9EYzw/SMcpGw
JZcsTAPWgGlq2D/ki+WGq4qjCs86Mic17kubM7812XQV7ZtxtLhzt3bUgEbgpuo8
iu914oovRVirpQBZt6WpJgGKkfqRp1/Ykq5T5+NciV8PbJUzd2wTmHE4VOPMwcIQ
K5vdJHCpw1cx/b3JhP9E+pqoTwqb56bSodKFQy0BvK0exvdo0A2hGfb7PZLpFsC5
6ZcDGaqf5i4QlS5C6Bz6wFyloNgQUVPhakGs6/vINY8TpYspsPiwe1HFEiL7TIHk
gLThQz+n7y9LlopCQ+g/Rzqq2EIGFlpLAP6i1eECszGeiAgGk04oPCmHZB6hJs0Q
sos0Hb/KYDI86+IqVUmHRlKLC9OupIWI7zUP+472hodgsxIZss2Rg67O+sCK44pP
eswTd7QVONm8FRyVpqDJCZtqph/bKkxMqkxu/f2R2nkCYATrAfc21SZ3UOUUqefD
botV7T6fOAj15bp7hTIpzvu9+bAcKxpy/mRf4vA78mjbgoasrRuTvRXc3chWl56n
4y5rl3PlR32n9FYvMWhn4MupY3OoL23RYpdYyFFqvYvjHBkGhyO3tL2qUGvG/3U7
z/KDvu+PfZcrnzbWHoQ4ggEffa3eVSXmFpgOuJQ+eKBGuzSs9oj/ShS6r5HgfXeV
h+A50ufWLeNyC3jt/BoLCAw3lcxZqUzOakSa4thP6VRHMDJAcFvCRyrtb93XkEtN
dVb9wHr78EVfQnQ3WeYQvMyO5vFA8ckljcT0SfKk3RIGfIvVCt5rC428ZZJ5Xs93
7bUsNYsuZVMOuyfTxnbJl/FgT9vCkT4L8KShfsDvCU/nJlNfUHfFGaNXs59JJkdY
OU0mCqqQNNjK/zxwQhqbTltVPqUyJfUinKt1Wca1TWS3VSNUv+lAhxGZl2Obe77e
QLUdkq39MoDyIDpwB2b4A3LKduxinLsgG3tkyTpnQ8GYr8c9GuL5BXAyboe2jyYs
VcTedbU7hAQh6Cz0SiZ+DDTzOtdT6LfR/+zwjFCWrjf9tg8OsD2SaSIBBhU3uELc
o9HHLUJJKO1Y3ciO1im3cSCiJS88YzWsrkCSczUeSSIgrM7q2G6qRBIVexAzWJT1
wCxNJZPDgFIZzjmb1PE2Vwyt94FZ6q2pspCjO/CWHG3ISLElLUT6jHLn4MgtFfB3
5BxWWVXb678DuJKOhqMptCQaM6F5b1IAhtch7uPXtEBK6TNT0BS6xIZXavEN2G5e
ZH4Cr30kgbePNPZF2tCHWNcsMOFjvHPcKpp8L7rfmL9f1CJUD9mtG9oyFhTtyvGM
GoCcZ6Cev6jZ3s0sHsyvUo1CraEyidK5a+Xq5R/nN4S2xmjefaNk/oyaMhIOMs8g
mB9TpZ7u8EB9aZqWUZyA8mVgjLDvB0kIH66ogm6uUdOEO3LRnkKA7L9fH7wRa82F
xnvx0zrhmZV36+8TVoFGszaNEBpGEHeulSD3qM1ODm9f7fw2y0oKHbu73h8WTe8h
fiWn4FtoL0luloYaqXOUo7DboR8ILKFTRsO4swlXit818VoRfcWGEct8Tm3NEOg8
N3usvLUBJQ49OnHVD+wgBcVAmAOExktCnbKfCqjzqmzulZaD4meZGJkQnKMceOT+
Tsp8cofKu9qSiTPkPgNAMwlaS+YDHsttLqk7k0E8ztbrNSY2LKhxzu9jTmX82aVL
Tb/k5EAkevcVS1csPHa7z9LCQ/zwf4fV9ELLS6hTjAo6dBJ+24uw2HL5DJ+KsGLA
U42cifNvB29eBdUUx1dEyhir+mjyb/vPlE334Q/sgMd8C2dEJcpGeW8sIs2vDnZ8
8A3QbeIjSkxsoQ0P1LWHsrclpaByK8zlabkgBvMDFTXSTkXPEkBBnYnyeAzfAJLd
zyR6eQJeevvNVGsdzWBmbJ88YAHDkna0LAIimnjsWFaGin8XwrGR9qmjV5qGx3C3
KJza7rWTAcDpuj4c5x347m+Ojwe9aKyvAwCpDTTPTus4RdIM35Wf8zmKRthNgjEK
fU7FdAzb9cHgYrpaWlq1az4FNhvsvDvXYX6IXmvl/1GCtdF7SiFw9lKbrc3afDo+
Ydb2ced+xQ/dbP+iThtqooGCx98DnXXQ3JW7meVH4cRvcCAc5DYP1d8FFcTLJTtg
j2X+m6nx3QoLz3+rmhgD8eZ3vHpZSRv+ScmCeBBwh80wIriFVx/vL2cuLmo58M8d
Mt+vn0WEAO88GOGWMzjEKX4kAeKPTC5RhY9jxw7w0mc7yUJLfmksCeA+Cf4xcS9z
LmCeqZUq5PWVoLXM4291y96MJS0H0J5om1eyVZeUSXQiltjnUn9ATY5PbTq3AyO3
H+9AN7BjN/hJBx6QQ6EYUm9rhUIVrlMqczJGchCj1bf2Vp5Y9JbmHvYYIrpcd2ch
0kqfsus1t77vXnid91ZIfHXpMG780PkmlEDxagkPF7bVE1Se9HOHbwfKM16XHcFu
kBMQ+dZQd4lp7WlaEp0UivxDqGNp0dGqL3OeLr81EJPRNgqfMQckMmFqTQ1BntcK
J11948TVA5NyybxEWzTC/D4i5StcQHR8P9q6G1h3Exce0ZSjO1uQrjwKgcWuVw47
I7bVUesuTSxj6ohl2dWxw3k37rJJ5mcJn6j5VO+ycGIqqdD9xhNB0KjvyvQLkxPS
ci7xbqKSV+knxC6EfNzwatdu1s3/nUu59DcTsj4aNHnPZnsCYJog6ioMEnzfh5Qf
6mqFyKS2RxxaL6LmPwYpjjbtFYbAFchpo2eWLAruit30jl6FcWmlRkJ6RJq+VdFy
X+d99NZ/ftiwd2l7qMUkr0VjeaLzjDGlOKTyaaghyDkvqisWILS39Du4SrDDLxAq
gBlv/nPsOBKuXWIbkagPMMY9LLEvCPgUzT8vgBwqNLaL6hNqFFgkzz4OuA2BIC89
I61EBJCxhAOU/8AESRycoVwNbAG41r6f/lWBKgg7U1de0/ErSEfN+Lihb4Ks4+aj
7vE+Q0lXsFIGQa00+TcCY3pBLSNNQrbvc9HMoI8B1r/pOo2anFPwi2u3yxi6dMbD
oPHjvTLTiPduXpMYnKvkXEWPfiyrapy9iLZxKC9iGSqjN9yBBodTechSaeiUOg/K
1C3DKh5/ys4wb+QQLcUkibklAA2uapQzXcoyFlyoJSFWYbXmeYOYNAd5/N5g+Avz
JZsHQAPs31LGzj51oAvrrzCzEDUu4drh+5/b5hNVs04YemmmojsW9oj+rEgt+ERf
KrKfkbNczmztpIRxKf2kOZDAA+Zs38aP4Z+rXAKZUHdK77OVwKQOXyMteYqaPJ7J
iIfdFdbkt69zIg5HwiFAS5/u6D6xXNmJJNxgUsAOVuQykztiwffHWZ7i39Sa9Wi3
+H/J3NtlFUgFwVLM6O1Mmm9i9LYaXCIMDSfQCAfzEr6YhKcXC3uDh7xKLQ0uy/CJ
VQ67NoEV8iU79eQO7ARyGzYE7ghtASlaFwawkfSvoB0dgcNR3zOEuL5AAwIPj2gn
yej6WYZ4WproqS7w+7koYzPEkaVY9XyDuv32BY0/w8empTFBTiPnmYZV1tWf7Upl
RnRQs6GcLutNZTaCgl6YgqsIQVSotuCURczIkmIGrPPOq53nkF+cxyYSHE/c+eIH
3dAyRPk1Adx+JhMXLVJLrHTYQ5BCOyRfHI/D5nmCgLo8oAXTnCsXeTFVlK0xOJ/d
CAA4As7HH7EKdLS/Gby9MHqQeAZtxd6z4JTflmBs/z4DBz+Usf4wrT0jM/uJ5l1T
xUQwT/ev5klmjDd89FAVdjPafkJB8k+xOYGx//S+iAcBcPU3rEG/hswcRyAMqVn2
9D9KO1lhImDzGCflVRim0ubF5BHe93HV8rVQscanxDVXTWi1O92oi18qXui05qZl
r6qw7+YGhgUGc2tgPjNELH8a56jwjPU+GN7fWx3fLvRkmsKq9ZfV1nViQUhN7x/w
EHHlnGh+pifcDNowtoU9vvoJLgQ5ZfsA9lPS927LE17mi5f8dIcrS+EVuPMOF35h
UjlZxDI5oSmtsVI8gOhuZ5U2ok0hy7/M4/4wYgZrVyeKlOv/rLF4SN0dmxzjTd0Z
d51ZGnUWH31mFGtmL2FGUzbXnWecSO6z3SrydzGyXWI8ldInFyPDwz4YNXT+CxZV
ZkYMvnvZSSgHGA9AbKIs3MM4+BV8rp22GvAk+wRE6dIXlKaxfTYPbjwyhYscLQwb
2/aclQbEG9F7QxieG3yY1rpymYlFnwJjTELNE+rOVmoD1m5S9IwZlpEReSGjN+4Y
y75r4Sq1CizO/+5CPJJ02hIn4bzZi8+WbcdS2SCTxtiO6wPYM33KPPEOBcFBPE1m
1ijHjO2xySOtPvH73tG265adcq26B0x3jIEVh92+iv36UY/ptNKQTTTClCe9RPMo
Lkkj/rfVccHu1dbP9h9CnG+zrbDT8XIsJ3XVWeMEEF/Agiv4Tg/BnwWk4U6a3UO7
XUZRHkzCezgsM0Y1W/bwIeLHw1qiHM66Z+7tQpZpIywWFC+6xqrcpqm+4buWJDWA
SWX3Sd/xEtTVOGvT3vgk244HoInOy4Tlp8eQZ1v2+aio/KLfkqFUyoS5xrnAOHTo
v7gEohNWhXXB3ziFmDBDsCzvOjW5JbWxshLqvErr+xdZiLrOMQ6a2CP5eUPUIqRf
+FycYx6ZbhCSfIanbhE+BnOIH3vRuLuS/GZXKN3NNrOeEjsoD2+yXojhIsuFbmWs
s3SnflawBKzw+oPx4P8st13GfZsWhs6WaqR4fnvS/dK4vdZxPjRE3UYDgcEtYccX
XeM6qBXobrAY78aIffcQbS2+E/N7LIZYJHB5IGYMokaFNFcGNux/6aOJQoPYjg6N
1GDAu27gW61H/fzm3YVPDXxeQg4w/LY0HAOQWFQrtUOEAqaT+uSuoOLSrZmJ5ZF4
e0qTdq/DwQItWAOYQKinyxJZDpv73RbJbMgoU7tSBf6lfe89x+St0Lw9pYl1DFEp
G153Zx0qSi1OFu58RnFQk9SyDOq0mhFNT1TJ6V7yMMnLf1U1ZrnugwdhrkUUY9Jf
InIOsJ6SpMZIYhGzqLxNjg/b65Nr7ng6z0KQnbJ5Eg3VcshQ866Hu0/oCijxi6xn
taft/8n2humypr9KfnRqegrJ9Ue0jpnK41fbW/rKa0EmMjpLS6XpAalbjsTJGZD6
QWSg6LmASDiY7slaj0g8GGfjmRC8LskaYvo/0Ns+RZniQMCIwTN0XLoeciL7DV33
h5hRrVzkyfzZyfzqpZqLd0zd5T6oZW4HwGgZSUH9el1VO8lRmr59TlLFPN0WbizJ
7JsMQo7d1zG9MZslmX+cgW1meGUT107hAss0V5gpDussgmNNQnk6+k8xkGC2Q59+
srRtg235ipprP9VINtXhAUWuILQtGq1Ni/UfLxwPP+zhMew7FPRfx5UXV85kAvBm
ia2WaputvKj6k1E/UEU15t1oV62IVijqxuLwUmW4D+Q7qkBdGxqgRrUSxvxmbOvJ
3HoWnWJnQK+YnKad6MGLvwI9b3UYU6pVJqGrqtilohj+TluQwXso7h1jGzx/WgTh
22JGDY1YJOI/LvZ34AlsHevc/6zsr0gUL2kShM1R/sSfRZpB8w4laO1Tqjfhg9aF
KYkYQERlqL3srdsxTPz9m2R448Q3OXpbpKff5w2AZVbLi1Qlcoekv4Nugs37ZOsu
AAlaY/6iX1zLif9V9f3B/fJ04Mbf87ZDoRJVwpSQLnnsJgH+k580MyEmsnwfcb5/
B+IhdNPJowDxXqoPXOVyfvZziPUp4EVcd/7KY5d61MjUhgOlyREUW03ZKuYioLrd
P2/t8rxsLYDtnrWuMEzinTC59DDnFeuhK7YlIiT4KGtNBMGttRHPIYiz4xuGEVb4
/SkTh0yPhbRaDih2cNku4qAjG0lQ2iNpzzH4N0zC1cviQwN7p5xMpqDCsm2d8jGB
dS6xnY42tunxQ9dwzOVcEqmpepoVVVTnuA5LKREwjplNC9zM7O8vvab6N+i7MbBm
68etwwJhOM8dyFDRIHmf6H6n7btg4so4znTy2Qop+idE9yVtj5DhH5kfYvhU3yzj
zKsA4jQC0duaAFgaw8ah8LE2suMaBva2q15CvK/ZVvTvvcXcvzq6kwWwPQ6SUUuy
Wvz0Dnvurb/7+odUzXoVqTnlxSj8TG6bwd5LZ9xUytWIlWvXgGn9lEBPfInONorb
BUIJqqtBt7C0AMQmLes/G5Qd5o5MWFEWoQkabnq1C+50xynjkDJUoqTe5OZK6OqT
PFFsKEUTg46uPjIyJZM3PfIWrfnEaDqFLU9tiMdhSKYLuzkufb9yWUhpLBEKuzHf
uyv/QugwAlVF0iDPTD8t1/ItsKpmdL8bDV63nLP2Z/d3R375L/11PqDbZCHIaazN
1lU9lWIjlT5USGi3pOE5F382k0ycCGf+4QGwycEzTCtJm58qzLdeVD3PtYhnrJH6
hNGUgG1L1cCJgFEMghzikSez7yz7vWMNvlhicEiOf9hxrqTGCZo2PtAoUz2BpimU
JIoXD+NM8H6jAWgDQoNfHEoiOvkMZyhmbQWfK/MJDrLCjFKSUKRrs4K76mG/wqex
qJQg5+8jrRMJ0LLD0x2kaCFusIxXA08lchSaZ5CHfXQB+aJVPNI3VFBeXsalfzu+
SLtR754SwEXfW3b9wsrYmMcn4YNdVzmJU5W9orb02C6VSVhnX3u++FoMU7s55ggw
8xBHQO2UDbnl1+dTokLkAP+B+ed8UwgIYI6KBheffekZM1tLIzgyy/P4Ggpn+UcH
TvfKCKewRip2H2gKvJXzjgnt53qTZpO7b6evvDzjGIOMJlouQWRk13xaUN7BfAYj
w1rXAKn5eaE9wO02zMd1uhfpZRXJdjew1cjdzcbvbXRV9m7OzDQcS66SOgt7PRNF
MPUoMg83iCQfgpNjRCoi2RxNI5nCbfk1TYLfzyrXRNM7HJv9K+6PIT+f+X5bDfU9
GQW/Gm0+Sd8DEY37AEU6scCUUZGv1oZ5fz/79aTob8CtXnDqxK3sl0VEJUrq97Er
4ppOh2d4BuT1tXwv8o1a2Q4GcvEI41RsP5MbnLTA2apmboRA5u4fm1Red3CPk7UD
dJZQCnU2XHgrJDlvgBXHh9x7qqJ3IFGWnBUPKJLRn11K3KBq28F4VUvqCNABHde+
`pragma protect end_protected
