// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
t0rhvGxgcvjdhSsck+MC/vmQV1F/FRV5cyurZNbopvRjMdrjZm6Lhgf2+YoK/n04
E1cuA6l1XSUclUwb7XMhF9KzkwGvSwflfH/PFuY3lbJlwT3L9+uV8G0EKeUxr4Ua
qn5qJ7gP0LFHcfl7yUn3wXBOZjWCDbgH4mkwcUy9ZGw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17504)
GlcxdmlbUDQhZtFV2E5L9otuQFUHZZhqXMpuqCW5TceZSR8AoQkeWT1N+zWobTXc
9Pw3iMiSmu9lM/6EO8TMmusC0tiX21y/PAr3mHU0B59UNylG1wkyoTxCdqlPkXmR
D0d1/JiO35MXlLXvxdTkL4YqzoHxc0i8eELlzj/s5ku2K7CyIWfD8RBkTaXNnyj4
KQuiVVGTHMvHK/idwLWqUZEPFnZdJN7UH8bpIV+ydddPTXi/r9/WfsBRfIRRNMy4
8vU/qDxPsfPSBj3ESy94d+FFx1O3YeXmA6q1RguL87n3exiealjMPu+LBEl1B1cq
mRPJdmoyygr1Isox2QA5rm7sPsyJOAkwXduEuWUVbIi1YlKSB47FJb9viwaB7m13
9rWHxHDdwvWT4Hrh3ZM1MCyY6XPKbBqwBvmCqYCAEIXFsbafWrIMF2RfwbW0H1Hx
A1/MFAtcphigXgQboNOs1vqaUz/pzSYpogc3og/CGM0b/rmJz75GNj+V98NA8dUh
7wN0q7uOm6OwM7pSEopXDqJ9VOpc7tvK4sM+FXFoNOaJopVhCk89SR9DGs4uwil3
77sjPm/pHgC4FNhbIAyTBk2z2m9bhYRXq+XabOcT+wyEOr9UkahioIQ7KnGjm9oe
8Y3O0Mpt6jUEvy24PKjVqZsEK03/4887ytuk8e4RuIZcb8crsx6I3Yzlf4NcBBm8
N13QG3BEHKstojPmpniXoWiAR4GMsmhxusJOeDRlcQ3IKw+Z7FFu2+Eiou8kkpSU
+lYEsNGs27eaudp/Mw2qdzglFRNpRc/3Ep67t+NRxvkPuXGiDRPlqwhc1LfztBun
zTS19VgSQoq+0xWLyGQTC2auJzBiK+SrqwlF4JdA5/CJ+SBJpWxtW/UA4/aSaDG4
Xk80/8Kg2WmXsJsejcu/GlKh73v4OU0E2AdIEsSB3KLcIQWOyhIZFy58v7fgtIYj
3DNSX1DGt5zaAF6cWFeqPokv2Mn8lXMaxHuq8R/HmHAG+RteOhKi7RCqi6Wc6dfl
e4zluugWBGvA92fxG4debIlRZpfxjKozBsVPGXNL1fWI8GzPl+IYhJEfse2A/Btj
G93v6EPQlnPTUfp1hmOI0WkmL3Ym+WfdQmTafEhTF7CPXGLPvvLYZ35ZKq0AeVBZ
MDmiehdhI6baaDS10KEP6bGb77tzrSxYzg6FgNAJlRUIRKso1ydKGWqPFkuVzKvp
73+n4wD2YR6nU2c/sPwdfZ5dLldyxZ+Yyzp2Gthe0KGQQhMvAoZhGkt1xUy5hvPk
ZbDn4WjizjvTSBAoDD9jzyT8j+sKwt2C1IRUovBScXEPx4HUYgOgy71dtBeZpJ3p
qwoiXhLgBoKL3Q3cn3Nq/sx3HNJEmZIY+qoo47GuX4XQo3nmXBQmar6PrXudM6WQ
I+CRh1nZ5EZR5cgeTZuJdOp00Wy1jqgOMv126Joy1IygAH84HajdFTQKG3bpdQcK
4MAn/Z5ewJG+bwXBMAAxC6FKzMhG8Itv0WN30rNsO8UPCwA3KTqIW99Kyx3n9ErZ
Mc4Zd/EdY5viIuswXB/+a2bfyQxB8BQck5lnJOqkBEGbn4xOPGy8H0eBdWdHyWQ0
8r/WpMJStgfEgTmoi6gaEqLhzynU4ycg+iSC94taHQ82bjkNmyrghibIwo0ORzfG
YhtkRRcjdLozTpS2iRHaB31K2hZ7Wumq4ZPe6yU4tthS4oN9XlljHwPjC4gXP2oa
yIMxxF1AE6M18IUUMzepQF+NhQMgsl272MskCQ6sta9XIVHTxVoIxWk7m0s+F9OE
7w8XOR/BBFCZ9KeEPG2/5TPQ0tt4UWpRchu2miG/CJK/TpUUeEuaIrrvZhS9MCja
nl1CEWry0O85L69c2ZHMml0KinHVyBdb65NvGKzpBQKx0a12Gc5jDL6V2+qwNr8p
TkTDzTSzV823ZRFLOL7RS1qlvyWnVHcSp6RPxnwUYRPxkD99NYVLq02QuwYpcRn6
lCbYPcXK5RmuGchJg9HqUxNtUQnzsuTK80vLNXxDOcXWy1nLH8AOlWFT5N/DbW2O
upKQlEk8LM+q1VKcFQnbokwM2z096bgs5nyHlJfpDYcqyRo1q4rHfvqCPCNgVx7Y
rZ+tZNdrxGslGOhdPJf9YHC+ASW857JBYqmPn+ectUtT6u7QSOQkjkrVdV49rZXN
Ck7REpEjOxqIH7Tp1u3vhbgh7TiACS/YJOTrHkv7Vl/akneXYva8ulPijZrCQI5p
rmvzOo6k7PnDBCQm70xwBbyz7xBKEDstl6R9SPmREgW3NavSmkxlY7dHWey4+2Pr
aurV79UuLKMhIA1dX5SS5oQ0TQ7VqigmQXuEIUmfcSLDyK+ga2JsvrGv+9TbqyzC
EXoQuBw5sJXw3VB3J89Y8tSUbGovy52yY3DREzy503FlSYGFiy7XWC/IcQ+kTbVm
lWUtCXqs2H9oTWrn5O9bYizAOLa6TSfg4gGnunQ033j/z3c1DFpDZKh9Zhqps/4L
O+H/o2mhP0g+ljBhpDfw0dVAbO0rntZZoa33C7cUAk6bMGEvoUlKd3Hp09LJ4B6V
WsW6WuW4IU8RkVeHehI+ZW3S7RZQZIvyyP+xxAHK0s4SJJU3zq8d5OTmLv/zuoT0
sHQaT0hC2Cz6oWR4u+pF9DsFwcitFDracnMUy7R4tI/0uLCvaTSziORocncawnAg
uPDcz32c/vW5FEvg7IGvGkvmfl3kO1aecd0txTkjlbPc9HTF4jSzpgZf99GQsJvv
X5TujfxwvSq9PpGcBZnJ+rZMmROCqeA/mvJTzHWoZN1P8qijGADUVSxP9iSsV+Xg
zlM7E2s0u5x2A2nB20tcE64Tb/hgd/YxzukNjeqS89unu8Hkn18ByYCpkM1IchRa
d6HZjoteexqce6+YaCbJtGyWTjcujKcI1QTf/gYG7C5SBSq5tP7rI1SMZ2IqUkfp
/gMCDpEp+Li+CBXm+Adz5rocfsYwldma8bV8CtL0KlcCo6B8y5xe9tWfr4Hw4Hj0
fLnDaCoOlWoKHDI3IBDIWGfg5quZC9imZjLDC1c6D4MkgtGu5J3yLfA5CWpqd52O
PoMy3T/LaPQb5dfMf5YiZiaZ505Bg888JWhAYs7oszISBD+jsyLIYMfPi2nmU0KI
JPd9OBbWZs1r6yVPq4JWE33OeGfTB4mVwD12ZgigBQ9IaIMTyM+cPPJpkKFhXm4w
eSyyHEad2jUsFpK0O5Ku51iTDz1SxRwj6BXDPXiamCxFela87kGWpXvOHwEN+0Y8
fcK5xRyNaFmNQVAJI2VJ+unoB/C53vMRLCV8YtpvzNKBfXwm+J2CBtX/lL3am8Qq
20lnWFj/vkbBguV2Isl+SZPyoJ30lFvU7mHsmxo/YhrRPr5mTT5Mgumrb+L3s89x
qtw3Ki8FwilbhcyoI8Wgn24VkJRD41bB7IZV6+Sy86eMRBkOs7xF29XZAwawJfL8
NWK5K33SS3Ji17vqkbPafIK/jS1XiV5iHDwntRwThRSjwCF8gp4wBdtx7j0gkxik
EmFTuuY3zrcCjN34OKZkDGhaGBtMrU8RazR0poArZ5PUtmvey5qmDA/PIXHEgIEy
0OEU14YznzzRxv/m6X4giS9+lakKOGnL9SroLJRXnTzSE2v73wUq3qZZqdNzCr8U
+1bqwIkPNLXTDDhPmbuA+NsuqmcWTcOOnzHGnF0XfakRn3NQeBKXIJ7kkjHZI9Jf
hgs0Chz1rRThDNj8wEs0S53diTYC2r47Cadft/WNiPkf2sLOWfbrjcaqGsBYqO+j
L2bwUMLTs71lInFCbZvUhY03GWg5FbKsxdxcPPSPu1HY3xwK0MxKN9wD/1YDZGMt
2x9Kq/5EivlC0/8wgJb5lDf/ZNCAtDsjZRBSMbEZstAbrP7HY6hmygaJwNfa9nib
LIrvmvFdVxBMoE/awhKqmAcv9uC1n21JTtpGi5iy1sZMkzeFpfsYigiCM+mWfzHZ
LlMyGP2wuMIyTmSmScH1/OY1zBaTHHsnrdwC61pHElUmqbIzWgGymNa9BYjGVC9e
YC7Owi6ze6GLEJmIHm6t+0vm4FzmZtHdayWC928FbZCg10h43zb1ISl4EPu1ooG2
dCxNl9E2ka0/PEs75dcHRpiT0xOl8Id87Z5as5uhaIL7QKNttnb5WNnThAa475l6
VYA7leGigat9sH5N57CVBnmw2Fht7kR4S4t6Ubu1gcP3Qt2bY09xT2PfAJskmiYi
WDKFLDPbixzSGtUuUnu1jcwPE441z24qUSHODCy4dvwt98yxo2YD0plBHK3Z9NGE
iLY/JVI3gwCCcEJKhD64vOIb0r3EMIYcBnbCc5nf5lFPU1/JmH1m/ig19NgePKlh
xrR4OmbxaCsq0EzTYsWNDLrsxeT8mxlWMrHY1GzZyQ+uT0x23Py+o+HARkm7OGDt
W0zignlNAsuYyC5tPRr6MRl0I8lGiz3M+nfmVJofGMPJt7SlemHgkNgd1ffXlBPS
VGHkdjAJLQrWf99jd21gqluXOo5YotWUPqplcKUnEVT9Je9eHNaHdfQwi2+JQUQ7
eXdpMtlETqG8xWFSjT/xhSLig2etUmMAGRa8xjNKTjdptlYPN7ppY2rNQP09hMLh
ZYMfYkiKqFrem2Pkikla9kKCvspMPs/4azlFky2SN6rECFvwELJVOPwxrphFUHiM
Zvgh6mafdSGZ4Wi9Gm2TYsm18an0E7fhtNE33T3m4Iow238gtqqWK2frCGSw8lVb
T2HZV3fr01hrAz42OR9aMUe7f3bms/vbN1Hsb0wlKjLzc2jKQ5P+OyVwvP7Eg+6w
AU5IpDHgXOIJq4b8b26o/n288sUU1Uj803pytZUG5lLnCH2VDJjy9ni7who+NwhF
9GuFu7Wq8HanExmgkPVPgucDZUJC4D/zna0MlZNngERoHEqpUYYA8bCSFZzRqLD9
qkYmRiNb2cvr8LWjwk6fUsNswYc6Iuv80ZgOm2mQ6Y0/sN8dAlIF9U9GmnDSCDyT
7zN0Jqmwpwgai+Z3ctE9RHAuEQJmXac5LjUr9rx5arpqGQszy2iwGChm9IA+yogU
ce24R4wHusIErgdCty3LcQn88eGnvBgCuD/vIp8B3Sl1ciAD0v8qK16Wzo55xHeu
C8MZCTmIAN4DBtbEVUbjyw5cPz59nYD+uZBTvhaYReidIgCGIdFp5TWpdQAemxRM
yHwsKPF+yy2W6wnhtyOebk68EalOR+Woi4mzSlpe5lWrjjOGvZ9A4NHn7PCzJYL0
F+nl/75CLi7XIQ9Y5+nH+rOfFVs5WaqyDsYHdPyXVlgZJ9dE0QlCPb2azypN6Xs9
+cdySND1LOZ1Hk8PJ1hRBMtC0222gtK3Y7xqijI8Cqi9wg/R3IBqnFjPVZ1UQmA2
YIk95VtQJc691n9lThcWh1Ei51l373eJTav6uVYDACwjq9yI6AXm0/67KDKqlymq
YfNG/R2nUqUtNCvS9JMMJQwMyvtF5d5vuw214yUe5ftiFXB9zqBlrfeD0ex2R2WJ
6WtywKyZP4357cMHxk9Ppcs7QAojBZgjuhLkWeLxA9FcOorStlw9OFOsrkB9WitE
3cboetnr8VZHVuRt8/EqvPhTFjp3qLZYsFP/T4/ER5qyXVrKMF9TOMlSiHZPlRtM
Zb+TuptitmQxj2zWAjdaSDDC8P1r23JCvJRfakPNLA2/IRc19cyBGBcOBf8G6/Wn
UELbgDo3A+yyXzZP0Vw3+ehZNFaPm40+qtjQ1Es2ypKXOxI6n6yZyfZS/a5RJTBb
OSo1EruNKSNBOrjrxuaP5Y4ALXeXrrgJfCZOUstURaP+5BpG9Mu9sMx/h5f3xZQk
ep/3YDBRJZvC40RSSSEwIaiVjl6xYvjrmPBuO2feLS1vny4bdYtylm6U8s+ZlC4Y
GAse5c0JBpK7nXW0cb1q25oAOQA5r9p9arz7MctfQoOZYjzbSOS3zXOEnxt53K3G
zAQ7NRguXMcQClZFGoehNZ+mSG6kanD9ut5BSSbrnMnNcMfgebrWKRZu0J7zwhw5
HqFgmjAM754oP9i0f/8LJUWULUbP2+VF+xc12BtDei2/CzB5p2QslD7pIy+LcWXT
MoUXrQk3Sylvj7J3IiWCV3zv5KC8MJSaNfboMnOxAuvj/s8Q+q752SHdhhcts3Yx
U1I+rIvkJcPFN0vpYLBRI+hbQ6njs+GDuipQh1dApzJb881GLXMOEfeC799ez/F+
EoEzR3Hxs5+nlKkFg6RoUAvn4+Z+dlO1YVybMdLoMwOwXCTzF8GJTn9+tDnDhjQc
7qzHd1m18Br1bv//P3vUMheepp1J++8PL43SGlHqPrfoyQzCCJiSavrPdg8LS1h0
uf1EbOiESqJdur2mWi8z+LZWhoca3wyeFWDzbx/2dA2MWGh/CsjvjUzJ5eaOiAN8
Rlij/8w2C/KmjJMMqfxBFE/Hjn9H40CTxKJ/uVhgCoDg3k1sXM0d4TiFAEO6lird
0ggU08O8HQFQiX6JJJ5dgw4ZCg5R1sE2imU17qTtfoPLNh8bpr3tgAKrbnQgbrSr
GF9voS9/rIQ2C4w7RQk6FV/UQQn72eQg3kDuzajINlHwNv/uFtWIQ6OuE7pCdc7N
NzXiHjor1FDzUn0GgV+s8PODLMNumVv2K0Qli28AfcFcyw7gSKKGAMBDFcKQ/n01
nulBKnTfaYTNl82cquu9saPMEkkBfDMfrEgOg9ndaV50RYbBWRCRtcriFh0A773/
WS85KuBTB6v7LnXbK426dmV+My0jpekxqWv4nYv84obAdXAdZDukviQZ4F7ZXtMa
43k+tgyqYKeNw0LXzs9CHdOCRAISpkGBlN653bKW89RgPtMJ74qGrtdPU5wKF3t6
0FSW/atn9dYxMfTvschyNgR+YiwVoQlYY1s0/d8P5o9xSPQBydr2qAzaY/JFIuy0
Rc83W/GgbOC9kuLosb4JttvIBVBW2ZzM+4HAwk3FkYOOR6VPqm7/we3G8KamsW5i
7Ts6Z5dh56sgRrVrXuSfBxapssTVSNvzLljAQ3j1jR929+xgEzKRVVZBOE0BBkJC
TV5tM9R63AtMIC97R0bVCyNz3Av9nELZByo4CBWkedBgBEVKktNHN2bSVEZwuxPw
MbAKQeGH+jl8pFCLN4iKlr+igQwr+7oa0XPpTn0Kkg0v84kctHzFjvL6NreG3zna
ym6P2NymvjYzE3Igw9tj0mjparRDjKBXKSgnD+fMC61hRzL0+B7MZf9QCGQOH37v
WWCLm9XqaY5lNNdiwy8ryIPsSVPh9w12IS2zfJTiHglBVAR9AK5v3OK7z09kGg1Z
5RlzSTa6vAD0JP+9dsFjRjeyGB5s0MPXM7FCyqG7cEISUail0DEq5xxwkBJAvkrh
6Y+SdnYPUghMCIKixHNzkVYisbUAHMdMuK5S2RZHonrdFGH8ubF47ZuMsvnXvtOK
BjdYcBvRdevuIJJGYKgBRJPKh5bpymaKXsvHmdG24c9dxvYloj8V1xoQ7qDoPjTZ
SwH2jSVbPi+JjBsGF3OyXp/nMW2dCRaxLNGWt4uBprIK6QeNjoVXFXqIyLLr30u2
uPA5/VP9G3sAK36ZQYkydzhGiR/lsxt+J6Z8trpVMxCHJa8VFW+l5FHj4Ns1s2fw
TSFpP46XnsL49xRCjd5Msv4nzG2JyzbdfeIwRpAJtvwYiR83bOCIRHICxiie0ju3
6ZZAkieui95ZrePsM+J8J3WiiuJSVInni63jYKHK5UiP+D1WtAJX0z1+GX6kIvis
ab4JznuKZS8eLaqsuRDCMiYOzZJ/eIS4gsGoHBOSBHZGL7QNkiuiRpbpAGNZdbut
OTKTw6BIvTmuBXv7d7s42iPXg26Xpsjc6mlcAGlpxuc9Hd/QZAFJnbbwDN+R7tiT
O62OuSS7gVyJlKMejYPadoALWYwCMLVtia6TbOvcyh+lbwSRf4j3OZVnY5pq3kdI
lGrPgA+q9pvLpNyyjyLECYjZQDVszXojKit49/Xy0VUotPn8s5jQIAbF0HYqIv/C
UBbbgLmqaXjLL1TSc3WMrmJ42TORgyJOq37sc10hgbNKlNx37ImwlY2RY5w9zAtv
EGxz8dQS5EiTgacedwMCNqjpA6xV7S78Xthx+8C4PYlwd4QCKvhaV3q7c5ik88VG
0nfxh5cpSpIYJwO0y1USVK1538aTMlwgOPz9g2gIYC94Qy1KL4wRriGnXYMcLllp
ufk7mXlV9elEENrlb5CWSWgh1ufnAsYzKF0lq8TiQUI7SVVpQQsxzk5WP+yTNCpu
NfebcxXAMP56CgQc1GoeBA2sOdAUVZQOIkLtFx6RgnpyPLDvnGpQlT9IYtoodZgZ
EQAohBvhZ1wlHqVCCH8BTmH6XRrXNic8haZ8bDBKw1RywsmW+WA7WDlu9GVHJHSm
70oVMygp4mrIlfeyxYmEAX/M5EGlxaeVJOLqCLz7AjCOLbQMHUBatY6AQv6uEujW
jQkVhbdvekQ4zk5UPCS46DpROTbo7zb6WffnwX2dgtp1rgnXTONibHkzm5bCvx+j
sp3rG455nIBLldP4dI+OzQB0ArcqIIQjcz2IG4Ej62C6YTPWeBOkxwP7PnVGGoyx
+ZbZrKk8KkzeodoeqH3w7qzSwkoQBpQFQiJI4uhNkxLjChjE3qUty02Hu+izKfGb
0vItJ+4Sjxw3RyviDEUgR0kvqVOf9BIA8w9BHmp2LqsqwRyeI4spvh9GikQj0RLq
/5QiWrk2u1UKQgII2sAdMZxd2cffCXtY5SDLLat4HjIkZYAqEsg2nIvw/UNXJa1h
TBd7CKdtQoYLw8D/t80v4D/VjMPr4kiwR/8VWTt2paEsev3fLbKyJrlM53F7cttJ
iNzGkS0260pb5MgCc7JE+kqKC3FS5M7mBGeGyZC3H/ji699Pl8ePDkTUvl+ajkaa
XcjQoTCkrIlNHcr5oIaopBs01k1l4dZImLzHQYqXIpL0rdkM+EK2gt07WlcyJoGO
Y7ekjRJu3+6Uqc5x7uWzOK0YwbnHLffq/Hrw6YyGoC1cme0mG2VAny4sLoAARtN/
J2z8Dvex0vUWYWzVsaWHzyvmKYFHeM0OMu8/xaguRMAKdYFWLMIc3AN8xbHQZgi1
sH3bYYdAefdKgNa4Ckr+8a/ekBaset5PmuYp6pKaQJW/iAl3wbmXgrA3N4zSriLD
hQ/6tIxqmD6EqGguWOmi9Djk07W+vdTys3kXMfV7VUwYnbi5ufo/lXucGt8LWTBv
pfrhWnMDyHEV+Sub3mapPtPItWzq7UM7/1voW4EBjXLZ7mtfvGYDHfIAjWyN7QmC
dV/OexFloo+c0QbbnodosWo/kLI0vCco0TFy5hF/ufSDz61osCBI1WMgUD+NSgMi
5nGR/GNTD8F+6KnshIJchRS5wgmTpSDTgi41vhiqw/4OTfsl1CD5XtibboSnd21h
2Du0R9Ne9QJwNic9i/6ovIXrATfkjxeVOwohmIlC7ZyP89Iy3x8RQDGwP1QOvwp/
gY5e+SJwOuecwp2hiXPiyhF2hJGEEfAF9VqEOV3tWNyuGPSCZeSAtjOuUE3HV08r
CL9vVWrcujSkH31jRtYXPAhNqSDKaXUFVhi6b8fScsX80v0JClUOb60kxY0Qfdh5
kaFtiquAFAURWOghGfSVC0SNnMHfu68p6j4PaFPUcAz2sHuLv+0r1G15YAsRZCAs
Nlm2nzt6xLIwrWZ+O9mgpt0SCDV1wynHvZXxrn1Hw9wxyfB86+6C0NiJMsq6hCc4
vUNrkyNGLkIFe7m9FNeBLe/sWCf3Aj8nHplXXoEtqHUizvbmkH6tIqtO/vkslFa9
PUHpN60TUJdD2j3n/IrmAiiA0BqVXOHv+2lfDIrj6jLLxE/iGNsdhzvoTUYervKE
pyFJ53ArpgUm6tk6MIXd+5woJN+JrsRxeU834jkW5Z5yB/V5FujyLcM7HPvWpWPb
VDhZFdGBTsIVzsaNmeCPFPU4wjcPb5Q/c1rfXlS6zK4AoMKfIkXYl/cXPykaojhU
+rZZ+waq8nYBd9BCuWU9/WSvwYBQXXcceqZyHQ99/qNqbptDA+ksBGS2r3Gx/IBc
Xtq5mPtI+jUNau2bH0TaPA3DBb5g919rMy2tWQ3A7/4/yH8XBAIONwU6ZXKOKwoP
WF1Ke9Umu4DQAsANj4cp2XtXyPnrbP3OB6RtWrY5hENju+51I/x29CTTnb/AiDgb
5/yDnSCIKEteqTpQPR7kEbWKf21hdMp8cKistbte38e+8NqWjJLSY9VikkEVjF89
Ok9aChU8y2MZSBkrEvhKDntqabYluUs6PqE436A9oZ0TlCfsGp9FHpwe/1QZYZZo
PBY4Z2T2QYaEiKP55fF+oFSPyDQRbUFHGd52yx6CFeNcxh7BIZX3f+tAQ1Kch2gN
wE2qQg6nkTCKkuBur/hWGK2vvyNDj+PV2JxpaD6b85qFI/t5Quz58nb7zZ1q2Kso
qUiPbPJBckzOaNe9BKhiLSlKwwsLlnlTLgHvtIoIuN1YFHvaBslc1WV9q0rCeRA2
Wc763/ruZuh1fH/+0u4XafBPVLSgEPTS1uxfID+CtsJEUp/aUP0Rz/fW6erLT7Gt
jm0By+nxxpfXxVQ65XuPa8xBwoKxHbQ7SjvSkgOYqTh0aBGj+7mUBLixh4WculEA
jpIdPjCOPgTIeh2nIRQQJ2HR8oB4E9K3S8Ngahwxv872aZtfBErDD9HSD65b1APq
AB5S9AHXjtdTE8x9sl7fZLpBjk7pxUKdOrlJhNt5kJrvMfJwsdGeproe/kPPfNFv
c0shCHN5TDQaeSZ8MMwrPKgCx1/fu1i/J+pnMvY+jXE/s59c8MoXi5DgBk71yJ3O
MsLD95Fu3s2gSRlcNbhXjgs60BloJq/xbu77pa8pMf6jFO0OC+pXKh9XHnj3K+d9
J99GhsYtR4y5vCfnSgYzyIkELWO47iIE0dynfmirK0ttAbX+VOs9Z7qglhWwEIqG
Z94K558Cw2yX2g4/+udffNbNsh+2DArZfEl/OX10Xazv6whdrc5H64GhqQH09ex2
BFgO8qvjqQNwy8Na4muhEsLpW2MHdRgDCvmnwbTN+P5kGYXXThrdl1nug0zd8AMW
H11raUfieDTU9AFf9akTbqSPvP3p0QmMsONQrdsh2aPSCP54+M4K+kNyEdr7seqq
hKjhvNn1IVezLam44KPcKRXcETboorh8r6nUwqAP5LiBSdO9hwEScQJwF+yOdXyP
cuNRziJKIt7UoeOSDS1lK8AsivVwAX6kyFYZP5Zzq35ghEfegQIKZ84CWnSYLZBf
VHP5qJopayjm4qaZIz/KVSk5o/dBKLoavYyNXfmKdxEsIevtV2fGVQr8/XNz9NsK
ipaU5ChOWaHO/yVdqQScOgxfU+ta4+ACO6EalW4NP9ITtKl3osr6LW3myyPtBmnH
kWk0AIT3hMRlv3kNW0+RRmG7edKQJ2Ro34X4wgZX3XOI6ek9vLGe3HtXgWu0YTEJ
32bRTwzhALvVXMa71nyYuBOLrTrObIppmKBnBysmntW/S+mOMomCIBVvQbCFIsyw
P+1kA+opJ+W53NyESI94WCoksXAY4LLlqWaCghUF6SIUuZFKsnytNwGz2f/LtUTR
4zmiWcKtr6jqRYfvNmDhllQbsXWSDW/+919OF4KmsjUl49wBt8AORDRTPvidDI7g
w8snq9lwVZG5IMKGpeKj5KAenmJ9eXGA84++P47vYrTly6RJkoZZtS/dheJHDP4t
Euqh3NjCC34v/98jgSMmOHFAHjy1FQG74MmXaQ0ZWb4LYaaJRCQdAqPcp8MIbC/P
lqEr16foKj2KJ9MvijfEB4n10PMasCYM3CgIwCcMB9JgPBtZzkbG8ngZdZxCvvQj
wJzLPsWSHu5JeOV4kbdWOVAWIQEMKFWdvfkihjgGyPIJ3QQCPwDxR6Soe8vlz68Z
4ZlzEfFDDdFMy5SIEhSNM07OEXH4EOdjHGuiHnhso/NHxZboTupX380y3X6UeAPJ
jEozrAOHa3tP6231FtdjxC133K7x32ZHdKlA7FFfjeVl+T0uYvM/XvNz9bccuoUQ
N7GP6zVHk7Mnzt592vaB2QQxnbUqvnF/mlpBkNrjSMzfqrCoz3LHxqX8J+GRkvuZ
4jRIMwsczYIfvGPsfty0tNTQymqciXZB8lL0zmuyYYu5BGTzOrQ4EKNiw+scg+rt
STrwTOKo4d6n0nvVfzjAxfXxrz0HEpS6iM+U+0BereSNfto74v2Q2z6X1zjErMxJ
f/6sA0vO9kPIWc5y47oDsYkrPVSxkqokqYU+YCGPovAUVwdgIhPmwqZd6etiZzjh
1+udZevl3mw8pUCCoAOcboH8pprX1OFGy59CtBJgSrDC5ocqE6KsmcJMbgb9Dw+L
6MmF3rqVKA3dKRRacAvzs85hMj3uQBn5z8sYV8W8STwji5IFcV6lfVjeL1e/WK4h
prAjaP4g8T9SRCtdEbUI7N03FSKvnqCMiR9etl601+AbuAt0iWSB/vhz+qcF+9BI
AFbr4elWOR57ENxTfvTgKFnkReSQG1YYq8USRWcgeGnkbyWvYEEx478DQjw8aOoM
u1uJgUOWn0pJDBjXDR60DCiv5x/K13n9v9SevEIP3S6XvLhtSKp6kh69KKz/xOYe
+GkEkBvCXs1jY7ThouGT12hOO0Mtem/nRJpgHDbsvkV5bzTjZYb3izyBScFj75pk
vIh9UoDdmjlhxVcgelK7zKYBewxInGE5rHJBQYUe22fy4mIOw+Fu8q4UXtw2Sqm8
tm13XxHAZWelf7W3OxyojcJRwCpzVpSqnN/3n4gNK9X67t06hsGwAKihZ+WS/ZJb
mw8Bd7u2OiWCxorSzgIpgBy/mEhXvat5ZZGCMYo0TwozLf7wNu7T2a+iNYsYZaaH
vZa+DKx8fzB1AtZYyFlTEWqdpwIcCYlgLMqw5lTrPcfVP60lXGA/E2nMEHiU9xZx
qszDzORjRwmsTKvs/YBOSV26cyvBm9fNAhMIf24CLJuY98uFnp0IfuEt6Rm7EApU
7ZgfAZjRyr6BDrI+e2GePlXoNtUCtuQwnhndHWaQSCrIa7z+E+SnGopRi8HyJRxZ
3jh9zHjfeAK7QM7kPvlChRZI4bLFAUMfZDD4CBAtUSI0yfgdK65mblTE9FFvJXMs
OZR4O/yNG9ngjT8c+I5V6jHoLCF0zeLqVQuPNHccNLdPNJAsAmOXP3xTg0etBaQu
c4P1T2H5ubcaHMKnnzs/y1h5TpmKYAp++FSNrwM1E1Zv6w+mbyX8VB/HT880Z72f
8QN/F1LDRLPiaxoEoSVO0QahcyIL9QT2baTslyth9VgxdpvpQM8UKZ66GkBpExeX
DgoAYskC9RpGlqxEJsKrkCJzpxUexzQXBbpkZ14ZXIcAKh1JUE7ILGrSKskRcSfu
0S1d4JCL3BdwkNFDAN5BdXZ0z8+ufEJN3AUAPtpfyteoVlQ8jSzoC+QIcyJNXG7p
xNzQZCDD40fe9BpF2ILbahsgmJfBh19CCgWZwKRgpR2ASz12PndMMlUJOPAwR8aE
D71vxOWpbjO3TCGHBPLJXn2jOrm4qmx+znxioD7dXZ0EH2VEYxRg0uvixejDvndv
3PQE1dOyhDcrRoZjo31UR+Z1kN0KpEqXufKGJXclaaN4wYUunTRF+en0ZkO5CE4x
8Is2pH9VZSymB3C/9UM3fGwN7Z/AbsCYRMH0sdiLN4jDKoO0g+V4cERIlPmnBsPY
GAYR9PxWPOwDqJWAwWZjDutj0bfhxWjwr96rDHiaehZvLSyg0N4TxhhtgJZWvQut
0DZLIWOSgDSR4Z3pZ7Z/Wyy+NgzQzpYt5EluoNsXEUeNRiujJ2zy9a5NPMGNOGEl
smFXlr45NqKJwpO94lA4gGy0EzRrc39n0SDkHsnnv+UztF8nx2EDmliAZWjtELfE
iP6WdCSrhSMSXRuv8631I+hzKrY0QQlQfFn2/lHC9M8Hd2ZdJx6XyPbF/ShYbqKh
Cz0nDV6ErWKuq/c2fcLWU7OUcd6hv76In6XypyvbBh05owi0CXJFlc5Zpg3k95ZC
iCu2iQhTsNusNX6dBQp9tzK+LhcKyvyZ49VCmuTPMimXANo8jAfUqphH3oSGKF63
cjZNTFjI9bTtbFYgxzeBmNfq50YSfZ+nSuAVksaSy/augnlWEGuP3hdd4nAL7hGe
wW67UQ5ME0jcDlX4YAcGKt/pYpyGLseoH9Ci78oeFuEV8rwIWEzkpufuSxkpiwQA
DZV2TPkTk/usk2zQ++qghggWXrrByVu555yFCr2w0pGDpQxXqm+VeQ9cAHUwBSGV
aE9/hhvYWPHJ9zttQgjrDKUsk4e9sSUD9exNdb+fqkZgiiOMjwMBhv25qiVMH/3a
wKjBlv+hfj6xI6SLCX3e43vua3ShN5aC0rahUWNaeaAbas7VHznwrPpp8IcCALeE
gPR9INrOhQaNJB4+pFOzJm/BY7hsSVigJxOjrS5gvVBtMci6UFi8k9zfOC63X7hr
PD1NfVqtTEaNFWCiuLAXwgof3J4mfaRCq/NrgW60jdh/wPKkZsKyXdyND7SU6f2r
TK6+WSe1se6EvIkmgI+28Wf8K3QmF6U71BFvp1GQr1TcNhVcnL7qq509f+y423EF
zDZHBJld9lMiYZrxli22VbEQ+6KzgNMIU22aGWBBCxwBLPhncwW+jdaJB8/H8zMw
K+VeNxcv6hWatXR4l135UCnXljZDDseaIv2o7jTLZ3pey2ihpbAy4LoD+9MCw/eH
qZ3sfaapDgBFUCxmgjvTrcjHBca9mGohboXW87Z1yBIJi6IptjNck6WXDCPOA1ny
XmnchSfb2R1U0P9EIHw275umgt6flsVDMwFE4d/ZuowaTJQhYbZsAzRWo6Urvj5T
SscbmHGbi6DdnZibpt6dcz3PSemQZUD1xhsBxu4k7FG4J5iyOModr2y32QG6OS2s
xPQhcyYSJoH+AX+F0+KsG1laUeAuEF9EZ+pwSoEi35WEBLt+i9E87w5eZiqOkW2n
msIr4KD+y9b+FQqbuJK4dvalWdsNcs5sjhU+8aWEzP7YtjTh5iUFynMzTWrP0GOw
Z35PC2t2DYCXx7AvZWWaWdaAPWy8es++ik89A95Bi7rcPUPDrCsv9bb7omE1JBRL
iwq7Q/zyUKQYSh8mimg+5sD4ggV5AWkQoI4e3IVwHr0Yy3s2AULSxY+LOyNEXtn4
Zg+9ZD4QRl5YcyJLEH618NFwWQtDUrKJdiGOv/8YPnOl5YkyV6/Z3AdTP11sJwJT
FDdbDjA1YWBrKREFsEuh/BCqh0Kq7SiTh3qPXG+nVoOKHyb5uVYQNjnx0ZIfdALY
8mA+pdV0kWqwfkaHobFuMSM7SRwXdsj/NuoBhKjqtC2m6tWdzJ4H5fIBImpvev+S
alFETVZqgBL0v9Dw6rTjCuuq0aZQdPhUEjVhBz7CEbfadWPLs5RQseHbuND13sZA
S6QU6+CviV/tQi91wasI0eTv7hhmrwQWbXCusvjymJl8+fZtPxCFmEcT4PSa/hHM
/Nrl54fm1fo95zW1E75pDFxAe1q81vxy5F3K7tt0ruFHF+bo1G0lvuWfI3pN8n5T
UTsPInMwaFirhU7RWsmjeW5qirtselQB6zZjoJTuDXeYaV33gQlfTr4kMlJs8E+u
5JqKGm5wTPynHxJyzX7ARLkXlVIIFeqGWQpHw8dRvNnEvvsH2VDyHAoBsMJ/NQqb
DvITYKWmCduA+ZZrd4NS1LGZLtvBDkzUwhQcBGda7u1JVdJQ+tCk/oZkzEIc50GO
aOrfrEVgZnqB/OCqOwmDA6g0vwzdjJ0fqNbSEZ66OY6JjrJaESUFP+6lluzuLFlf
2wYys+bIbJ9GIEhnBhukuTGwQe7d2Q1doxWYTQlaT4VVsIX6LjGd8MIVuWQbQRTT
OyVQgkoboLOnd+wLqUAOe0CsyQofnOuwAd7eC2mlcCQZX87rqCfJQDASJ83bbYuE
wwKjAQfQtFPfH9wFaTbBtK8qPcPC/sdAHIkZAkGpJeoI5Mi/kvn9JKPtF+Bqf2ga
YuTeP+0VFqnyfUhlr0oIrLLr/12aSKoPBCu9kgZWCRajO2NaHsD8RCxtMDWeJpXh
FCV1WNqIEpehfidU4RytL5BtB025eJd39elQxB3C7dGaNT6hpa+vTlkxiFhB+sHL
VPgr1e6gBJedMQ1tQJ1VAhHj80U+o7dzcj9RJ6un+iDLJHjsDYnzeirUzhydCtEx
03DYJAAhI7/KlPcRf/lt606kBYYauqvuB9I4VG8pQXCGdKx9Mf41ieYdIU41FG29
ahTo9P4cbh6ZziubBBbN0lgeAaiAJ8f3SHU8Xw8fPm/8wfT6xhQ1hNVxbbH9FFGx
UNUwV7XohtDA5K9uY9xkiFW6INHLtP8fzMViHSk+wRcC/VyCCUqBCzk3FGvcmWeE
kBzeF0PLJwgcV8usZKP3nspb5mDMRKqT/SEv1RntWfvXD6/ipYlTCQg/FBhVX2FH
gj7m+U3dzZ/bMlfjfkwqRwAGkasVejOnH17puobZQvMwV8ofzxJD/93JAqGXm8On
OqPGTYrbKkK0go/nzyaES+jR/X7ET11g4dEHvi2YBeTE2tk6CFG7cNK8o0sfM2vs
zhTem4K2Egqh/zUFdOSal1uPTNoddL2tS4nlm7K5rZ5BgZfzxxWgMO8ueHa6cJmp
BvcVSwiWj0TLnANXR/R8odBFYuzA0KQeKCnUXcW3GAurMEFb7zZQerlV/TeqeiTY
FSx1QzluYIdPgtvWB6jCFoTNZKZFZ95ywcs+YMjJocfokgJCFvd9rX4Mrb892Zoy
RC5Do4PbB1P9Jh78SG7+8pBMU7nniyBYFpxyOt8jk/S94ZmigAEEerjZvnx4VVPa
G2Ty5KEtYlIXLwngvDfwrSThWZjXbLN463P3TbkEXZVcCvQcnW6WdOJehq1G1VxR
I/DfzShf/83AtDTKI5CBCBLsZYTna+wdEJS5/dTRXiE+eFkS4nlfN5vWR4psbcgM
bgJiNEssE986JWeKaaZoZwiJG18aXNEvesJFBLcASILm8alzAf4y+M58NX4PW1NX
eSbaODED3IdqRGvjxye1bfMR/RGLeYw0eo8idB3YEWRQpOD+u67gK9GJst2OZvaM
H+jAiXCawfmF9s0IywNbHFnTvzYy49yYsKlg07/KkkYENS92TfOKmqgW0UVyhJI4
f4mqFLA0Y4biO+llDUcCm4w5TZZhqhvsvAS4dOqPmHofgTx0pjY82GhN9CTRvAyu
YKTZFEvOL9mqJOw0929XozsQCT7RU+8YbuSWU2sn1J/KR+53yu0pIUc1+FfGeimV
jgj59cGIBq3RkRUcEZotmbw4+skH6fXO7YkbcSFyeeTpGacDTr1naMj8ULIO/iYH
tDRSwygUesoatlxBdi293vftHF9LBFSJiLS28itgE3ByjjSha8u2WcPWk0mP7D/Z
KX2Fw/7e9Pdml0kIZspAzvBUTOkSRUVjRHsVqfHIkFACZUl1YEEhCkoIZpB6sJmN
Tuk+zgcheKmkw+ZGq3t2g6QzD6ARfv0gZ3nRH1uNEHWZWWlNKLvpnUfVYYTqekt6
vV7Pb8aQ74BjtZVUfoJJE3i3TUAkqMQiaFa74xudyqCTQKqi9AgDs49nl2rNUyJw
+WwFjsnPRmyS6uBfYHpwnF/osswUfBq5/Syx7UfwNhrqIy2sXoRQjiABZXxT2HNn
rSX+avx9BFoJzQuvkatHEG3QksKg/55nqkOOFQeBZJnDqh0VR29tK//6ZM78z70N
mb8ZsYuNvTm4Xj435NBGcyh1ise1cToGgI+e/JkpLcKcYpvFV/xGXIf6ksZFYlQ8
T+0wtPPSWVIZzWxGpDFYNd4Rg9ZQZwdJBtgZogbf/HTWByna1qWOSj5Mopg9SLxR
hU4ttg+p8MWWcnPk1j3dqjgZUHFFhx+Xm7A0oSzyovtHYXAL3haPQEuiQb4RZ99V
x0iwcxgyyj2gmUThpJWlS4YaSkJgsYf9D7bq/H7BYN3ofiPTcrGe/Npbb8nDoFM1
zhJNFkgwqz983fM5Tr2Q/Mu6Dnlu342F4gAMI0F66MMjrga0baJpTKWbU9ZhjljK
JOuRSR+yLLfxOC/ZQ7BmMzjjHhK7ZPuV/pMzmObod8aBaW+PzOiR3zNbMnfoJe0f
eYu4lzrzu0qQb5UTFaWWUoeRpiSkSeZpL9m7xDiCjUA779GobVUJBhRS1LyLQ2Ki
gFO1G4i2MPeI830DhPQkkU/RnTpNqUvKGPrNEUONgpEVNFTaV4H3ooIyI2+u6lzk
ag5OLczU5PY3AW/94bkf8Q4AJLg4kzv6SAm40tDJXUpGX2SRG1HaRCMtdM6ts6KZ
qtyN4jLbc2zyX+4H821G7UBDyiODGpEZcWmy04DaWoyk7cDpWm/E+xxewD7cv8Zr
0lbVwC4EP7sUKTM+tKKKkC+7LW3OyFZ3nygStllkYNmm13CQNXlInmoRBJLz6GEQ
XREcbN5J8Ccs+J+SYf9H46QctUo2Rhs44sQ9fe6vbzhqKykK294cm6hTGfHATLB7
omeA+LuOxy3PDJUnXl8YS28Y53k8alhTHZrwCEkQnVlkG43uPIiXTVcUrDQZspiX
1pb/4LBMPWvEi+SzdkkuzRqRDlfaG7+5Fzne+Ulch4bEfRMOTeX/MliLGlQ5N02E
trq2JoEkBLHGmSHF4uwNlP9gCrJvTYaToZg7mGoOtcGY3qI9ooy8/BJ6r8i6Ak80
kT6e0bv5WprCbb4kxnmPeS8PrhkIHpC5uQt0W3tKbkcUgnNgyIyk0mw0I8fy5ich
+FlvgUMevIQszD2HsF74yk3T+QsuNU3ZKQEk3PDSHBBe1dwkzILNQaiEDDqcnJJt
UfQcsStQv733xyKoZpDGtO9ESKcBaJHM/EozrXoIYviCnsHA6X7R7ouVTpb/GxOv
Ml0gmpp4XL+Sz9zt7ZH+VwMdvusxpMgu/ntZPf48HxreEx0GB4ZDopwkZQWIs+3s
R37+OBm82viK0JiT3Q7K/usItX1jB7bS+5xoYhNQ2nym1ISsRnQYYx7WRjKM8U5U
RuyrHvNDiCT3kJwoBOv98+4eiyH3ZHSR2SdlCHmQt81CpLwk/Wz+QjwcLcyCv8Rx
e03AtLEuCsczbA8tNBAXvOxNct+DEBU3OU0oWHZi5HsRzky83djbSklsUeh8qdXG
TDtmqkdCQoENczcSmXmnRtudA4DsZkxNRkxgwxpzYcG9MOAw69c9qQzTnyO7AfFv
xzRN8Dy3O5f57LoqtwAosWbOpfVX2ZgLr/ixMhM8sEP9LVZrKPe7570g3VFJkIUq
Q1QvLrLhS7KgFLShgCm7s0U/sbYCa8w3kI5hh65YWvjjovG0O6aAvYIfHkQeq9Cq
k0qz8+mB356XQr1/PyV7VqR/DX2PGuv6auuYdB8idgnfMbuDYtIki8gZjhdoxPZN
FRiuqaszNuP0uPi4NZT6rPFVzw3bpZTs9l1w/PeulhwFJAKV8m1gvDroVXTF+8M7
vGpiqzxQvTJVPTRxspdezwkjrIec6jfxGnsBhVG2Mg/eQkHv3eVeDPtc6+fglUH0
iAttE8810J+fxkOD6s32D5iQIbbdR3W4/xnGK3WeifO57dlDweq7Sf/4E5s3qysP
e8wVeHe5RwgAD5ftWVb5rBc2b0jLuiiaO5xX5tImCfyqWtJSLJZuudN7pcoS0gNX
e4zmRDGGWO4rOTmoeq5zGJqlbYd62RCuFzVJaXDBGwoRVsA7INEuKbMnPbQ5xlw/
7CLF7eH/0zYQjP/qfrIyuGlPn+SebkPq+V6YoPaoeMkrH1kCbII/KEA7tcqf8V4v
/AdMpNFlNP5BeUuHWxFeOOcoEw0fVY2FGtkrQQP1xnjgmkYScCJha4PVUqeFqbVi
MlgAeLZkc9Fr3d0TGWdRl9zGCkUGFTgNV+6R7S6ofQU3HjjOLXIMTg0ehC1TgEJ2
NQIuzgDNTJQooD5+9wVT+XQjQ+d6SjJj6+JmmPHgxfw2qhvprDDlmBgjapl+8NMG
ULvjUQEFsgJwPXW2N/zffBnOaLv/YYdyoRv+d6zD1Dki/T0/Tnns1kq5bl3XfcIc
KRk9heGQTVz1mBWo4ppzg4gFmOq3BIUr+gKYyDoq1RTCZaJZn7UUdZaZ5XtvffZX
ms27yz6jSD1YZPlva9ze28RrLdBwpugCU4dHvhaQ/W1veQEZXTHA616C4opQx52b
8WONRxDvMtptRfZ3ju+aG6sjj206McCpDfZr9ufC2t/cM2bXD3sZSMukraf8biLc
3Eucdnq3x/gBrrHlZHHNjTh1Xw+EovMQBx7DG2Eo4sBTXJSAUAL8LbpIj8bR06nN
OicWXC6hpCAF9DMaga74CxTIzkAj+hxA6LwQgQ7NcQoxwwm4Sa4e/mW86Am08PaB
hSqHw9x4JL8AWiyaAsjLOqaExtIJjgmX4zGEBf9CRsin5EtCHrf9Tn1AHmHp1QqR
Yoyo3cta4JUO4O+VTDPsmokNMVFBFxYnCwoIeqEjPbbtNpkZKcSc0+COQkrNz4ru
nF0ZMI8x9mmqZIrxUIx1UZf2ep+suOullF7Ok9e9U9qcsNQ9edF7ELpu/GylKdSa
6r6wYDThdMVdBSWN8bC2+2P/DwfL8iC41QkOCR50aZ5j0Z1wcXnbQsptfqqzfEZw
mC6nNPXnf2ypsSqS6wbNSIX9P7MAvq+utLNVq1lgJoSiIHL+FvwL7pNLm4af9qSd
Ac11O26aemLfG5QbVMU2VYcxO/opUmM+YmkDccR4sv5FJ+1dc/MWcKYazT30JY9m
7l+6KKg506uQi1jmikltpu4wGg2XELLcKeiYvSf57voPXw5/52VLhb+KeBHlIbJg
z30jKUGhDw+ChdOnFkGfizWEcYs4XXJjThCilqfWRyu2eb/9riM1e15C7lW1z8gN
0mCnqpyz9JoOkLDlPqVPeBb5vFWK2vFBIJWmUvaRBLNwDgY7JbqxQcxMDGuRparU
ItK66w4/lDXuqj9F8lDqACjHT11Q/v4KFwugEIKQ3DAqJdIFshBSX6XJb406S++I
ERER4sUHg9a18b9hwRslCAYcrvcfsPLTvGHWJMTVYlCitS2+S55VhZs4HfndfZrD
6kGVZ1KF8tpTSMnhkh1Obbd0/pv5+T66KFWekXRAnrIUY3LCJVO5t2kacgdvDEKq
Qs6yqpX/Y4eaWhyIUiAfYcG6he501FAMO6ieHvaSGkJwdUhL/HqA/Ew448HfEMAr
2EEhRvwTm9Y/0Iy0L0g+aczHDyJWawZ5woizhRbamrQzWkdHb0oCA9QsChEq4BUm
Jomk7fYKw8y7A3IaHglX36nY7vXedXeerf5LnEJ0GY+o9O7OlZ4K5GzEYZCF57Ba
dg+baSk74XPmbzbQJYpo8cF0tJ8kQ/eaPhCEpI+OzIwmJ0X8H3/CEx4cTG8u4wB2
X7bHxF3hX5eOvJ2J/KjmxzHfCTNNLYBeMsy4DNPSPGcoP2NJOLk9nIIrOIWjJqA1
E/qFar83pGCSTinkNqeX4RGCn4tQNIO3Jai7MuVtOw+hvEQWXnqCSZm6VPdgsT0z
mdkxazTsr9RRVRGOFVbB/IodOswp0u3TKm5yIreFh6pIieZCAro2viJzNmBOyNDA
3srSRf8GhWx32l3IWmwmiiA5VcsRhLPIREgK1+dvaBDx45LRbdWWUzVBlZDys2zm
EBlx7N031SM3JRNtQzHThmFP9hxtxKsewoAio+upSH6xHzQKeTchtJYyDnj9Z+og
27uqopqKklOe7ksCr2MNLO1VPFfN1Ik7pk7Pg6I4PindqlEUDazC6TuP0kIHqsUC
18vMSpmzzYMM1W54k+ni0anyvdkuvh5sXBGDxXB3jUQzXRSkxRusciqnYHvah9PC
dUU5fgID9svAhZQhEqjEbUHzE57SI5IyjydyK4yAzbGJx/6bV/CBuKmsNs+L2iEF
6bftLrNDXEnk1tYFsT2n86k1TSVTZQI4Ud49qyIfqpqQ6FsdSVojnBMhkHrDnHB1
cU2Ip3lj7HiZ+R9EvhNsXniQ/g/YRwr5EziP3PQh5iovQIEY3CQkmHyaNK+IKWZk
KzYM7Mf46exXwBnLkgCkp5ecIQS5AuORoDJUm0hhgf2McaruwPjd+z0FHDlNTSwm
tXM501TpI+B+NYjjUjVKn4a2sBx4aWTQq0BmwDBs1vGbipMCaTycS7KCkPIArAUX
RA24cHLgSrrzxEeoUgihROk+J5ffPuaE5WQOWLpyCHsJEGnX7E6v2YlGwqbr0FeS
rUNaEToCj0jqPHgq0oxwf2vRYcdLtJxipc6kUBILWhgQlOSGaDrNRjs6Lpbc9mRN
wgdxvETyMaO4Hnozv2C60wJrxQjPcRiZEB7xJMkkN75Tpjhu+bFKtdvC8Pby9wWx
i573TWNKweXz8BhoTthbnvhtlvA0ZiguD+WGxLeK3Lm191nDMqOxELY3MCzMsELH
zfMXDwMxUseHpO5ZZxsZqgA8v3xV8bRAa2+P/YxJbLO+wneacKqOoghiKXkI/Ixk
JrYAJOYCd0bocRtKaSTceL2IuKyf9IjyQJsLtNevu6z5kFt1JDXmCmWKrXEAnAEJ
15z4p/uTJz1iWTVgrLvBoPowJxLHbbu3pNnKzrW7gtM57XTG03aIY8JRS5NS0LmB
tqvChe1h3VP1F36xtO9gKrND032jLXk77Sd0L1damVHLXQTFN0dhgjkUuUdpCxE/
C6W83IDMFV1BATKIF0BhMS8xevOT/ncmgULSzM+d5dOPplb3kOY0/FgJ8Rniysbb
e0LKB34Pyp3K/LKHC1gdGk5KwoMmKRcGlEZvUGcMk9BoNavnhuve8P29k2KRV/N9
RtP5yIwfrm3Poncl3YtA46l66Q1pAF/4ejTMaJwbDLhG7NICriWbyYWzobSZ470a
0OFX3PzXpJEbrI1nnYZnOFjSOgL4NCD7Bmn28++wiRel6TXB/PNqUcNb7YxmGBcg
YO8GGqnxW5TkmSHaINzsFTqwkCY+pgnWsq2dpUzGDDN/+axai3h6lDkVpmPkUsSI
WrKq9zTNG0NqqbewnTda3TvMXz85FGBf5+Tp1lysJxxX1LbHgnnf1f5PoObQoZ/l
RqIY0JG+KTwrGzooxmEvpmOcz2UmArfIF/0x9QE+YxrISv9UKiQAdEXcq19NHSxw
lvVKct9tYZxS9R1Oy2dxp/2xbidgH7cx+WiVDbXclsjQy4QzVoy5s4iGUXI8adky
wmHcVQYedtWO/TeRW396YUK7Z02zxk/3wrhR08CO9ZAuJhhcUSkj0lZhtw/QPk+3
YUGWURDBOLoNFEAm2v4sHfKijX+Pk1XiQ6sLvkJr2yRoj39bfwo6ySCcVrfao4Oz
ghz3v+zLfkbCIVGfzGshby3oy6FjZqEVfXstI6faolg=
`pragma protect end_protected
