��/  �?ؼ�ǂ%�*���H�%l�`����EPn�SJ��������3���9�ͅ0ɹd��t���PY�2x�a0��?���Ŕ�j��i�,�E���������Mj����ĵ
h�̮�
2BA	�/�h���(��Si!3�xm�D�\�jC�Y��Ѥ�}1���Ԋ����H����#{@��)	�<�:3eE<�᭮��yJ�Z��X^dݭ5W�!L�cSa�&,�q��zN8�[�cӭ!��K��,#�U�������k�#!�ܼ�jH�i!r��$�ۃ7�g�ۇ�P��J���F��dN�[y��Ov�4�eC"�Sd>S�}���/�;rȅ�d�a�e_�Qx�¹����xc�u��S�@�����w��n��M�֮a�G�����U+�e*���'V�!�}W�j�LRQ�=CpY����<��9UK�V�"��	RL� ���a6�]x�_iX�m��rʙ�'g.E3e�v[��fS�@�	$�%���U=l�\�|���-���h�YL7~)4����x�E��1���L�W�L�>F6�_݈�7�2!�Γ�j#dC���s)!U��tY$t�lE��?7�n(L$�3�iB��6��s���˶-7SOg�ș��,�Q5��Ɲ���#���w�����g8o7���8N�$K~SfdI�k2���dR�p�^=r��T� ���P�)�q�e/*=�^E9����Z(��V]�:[.��7��d �N�<�湵�_k4C�oBG��x ���34����|�����6p�8��ܩT��yW�=	�b� V#�����(�Bk�w6���?�\v!��q�� 0+��y�ØVi��s�}�r�yf�;�������+d�Fu����q�s{���I�O�4w�*�����a��n)B+LQlu�(K�J�
�e�o�ʬƯ�� ��2����v�G��n�fnW�� i�Pw���%�W�
�u��Z�-�m1�x]
��1�.te\�JW�e�i=��%RR���մv� o!�<�C
���bU�@A�����'�|O��~%��D��q�sB4i��Ó+��a�@ڎ�a�����t�+�Y
����;����uxY�zo�9(씌yS:ff;�"��M{t�{��Q]��(��g����e�M���"�,�(�z*��Hg�l�wa͠�Pai�ؼ� �[.�a>6�W���J�¼���t�/�4��#Z���&��M��z����J��'�e:=��tiZ6灜��9j����Zx�v)��M��%&��B��ʆ�Ւ���`�My�f��j,2#`�1�u��.(��� �z�|{n%�Ap�`M�ޜ�z�q��	nj�G��~�c�	.��#D�����I���[0�/6l�p������tyU��<���j��jh��֩�Ê \���6U|���U!DΦ/U�1,K��QxK�)�{UGbk/Tn)�Fp��
t/Kp�����L0�c2����Gг9b����2�o�p�q�|U�I����bM��
�P]�U=���z}�����đ(o���*E���2�p�����#AD[����υQ5��ނ����T�_-ii����Y�7o�c"��r���u8� �a��D��!�lR�(�@䛗�\/IJ`kt���t!v��m�~�}��f�V�e��tt���������&��)�Ib��j9C@��$�#JS�k�'+f�$�okVt�D*Q�X|�%PB�j`3s��m�G_sם�h���#?(�O��;8��g����-ܿj��d�W��`^���z�c������<Ѽ��/K�8'�4i���R#V�9�Jd'�� �KS`�^�]���Ɯ�FP����C���`��`{���C� ��s�j���L�Ks�Y�d���^7.^7g_�l�mN�~X6?��n�u_(�&��<�f�CI��~�s��#�xE)�%� }���18��Փ��t�A����AޥA\�ra^%�;��C�Y�l*O��8
[J��<�X`2�S8i��:š�b�?E
���sE	��b>��GM%	\/�=θ�l7W���5��**�Y����YP�|�E2S��}�:S�eS7t"�g�Ŷ3
�@)�b�u� �O����e��`��NK��B� �m8��Qsz�=��)�\߲�GV�?Q�3@�M���R�|�<��3J�Z�LT틺y,'�T���9�]@���P4D�{�jb�6 T�AY+���G��z���].gmeu�v���W��� a�����K�m�Ҕ�<�,�����2
=��Է����29��P���0�ôb�/�XP�y���lg���k��v1��]�7{��,�v�7��0����	4�({��4�٠њ���V�E�1�G������qy��ꤎ�a
hW�ѩ� ���G��ˑ���`;)O�`I3�_*������t��x��3�FR �/w��"�T!z�+ �l����/���@��h&T���$%鎁�N�wM���H}-���ĹF8�!���i��i'�L���$[�)
LP�x���+-��q�����9;蟐���눂&Uo�3+�F_#2R��/�l��F�R�a�,�}����j�S�d�����7H�0(�A��@Q�� �{��+"k���_ăc����\=٫k��2�)��ѨG�)W�Y�X*����s��P�k��I���)��y�U;�JA5+F��E׫OY�ljU6����&�gi����!��}�S���>J�`�:,4�̼������
�U)'��ɼH3b80G-�N�{1��<���z�fQ��E�Be���U�=�������\�۾A	6�,�F$��e���y�9KQ��;\G,���.�^��]���c"OtT'�+��y]��;9}r�qS/ڱ�]:c8�
��lq	��և}V��X�y�+nyl���oH"�O�m��OD'�J&A ��팽����06G����	gB��g���$�{/�0ɔq���c�l4��}�1db6��:�"R܊��_Q�p���h>.��Y,�{{9)�xc������!}Z���O�~&�������l��2N�`���f���6W��[����?{�'�Et_Q����@B�(��k�mln>���=؝��"�Q�AJ-�b{��Н�\��OwuM�6�$��$	�hŊӜ4 H>,A�_���j+���y&\���w�TXؑ��Z�*X'8o����.��K����A:-�f�㤧�lB�|��w:�F�i:��*H�l�p�Ƨ�g���*����yQ�����P^6m�c�qq��3e%?�O�~V�5��??�����oY�td`��&��C�E��ag�v�~�Lje� ����#��%=du�R%����g�n6���(Mvу�ܨ�"qF����vG�jY%�t�i�_[��r����l���8=��V�{�b���<o���w�%Kc灷���Bui�Y2����њy��k�؉�?ܠ㐆j�A;mf{EXQ�F�
U�|GΆ֝��
ɬ}�d���x����Y����9�G�<E(C���i��OĈĚ����%��\�s~O��$�/	Gy����
􅧌�p��݀�_>��@����5}����U�	���D{O$�,�	y�.ڠ�T��b���_Sk:hl3Z��D��t�aB�c��H��^=A�8@0F��[����BU6�OH/-�?�.����[59;�I�v?��@:��ufLݭy���pX���NL�yL��6F���oD������X�Ī�r��X���q�I���Hb��57H'`�{0G�z�3�\�-~;/t������'�8Ӳ4��=k�f9�G�i�Y[94�|,�KD���V���?��X�L,��ܾ�4�4�y��Q��2��nF��ɍ��Z��J;0��񬪈��2���a�ͣӎ�S�]�������{�MDY��.��!zÍ��<�x\� � w���s���h�%��owx&�`A�&�_�	&M݇i��-�l��컒�;y�@�<���Yt�F��H~�P!���Plg�P,���3mx`\x!߀�侞P�'�S�%�
��zO�X8+���rM��NЛD�~j%��kf����D�S(w���J���U�2�e��c��!�Ds�«G���tj�Ր�������&�kd���<��=>ŵo�b3�����)j��`��DT�뱺�p��q���eb�����l������6�p�h��V���Ԅѭ�e
r��Y��=���ndh#黹�k�\̷�>�u�4Z/���޽(���!���rSm'c�Ȧ�4�3޴Xr�`�ZAE�g���@�7&qT�4�H��re;���j��zvU(5�=��S���P�E�Zo0���T��O_�e���aٽ��>*�bY.�[�v��V��8c� _J0g�	ӛM�BVK�2f���%x4c������6�%ܑSR&��-z��3�Ha��VK�������,˲������<���͘�C�7�M\ȴ��Y|#��b{Z����۾��9\G�o���9�D�����9^k�*��~�D���H�lB<9�ձ��<&tOT����$s��7�#Ѭh˵�f���-�a�#Ҡ��@q�U2�J{<Hy���#��I<�n�m�����OZB���|��2>N�-uƘ����D��b��2��r�7��S�Ɨ�R%W�c>z��<�~`�W�M�"{�R�Ȓ�&D>+\^;w�(Y�D*�5�����ó����-����b�L�B�-�B^&���|�rc*9���˻� ��~�mLQ�zQs�ݞ�������?���2�~X�--H�Ǥ"6�6���@4�W�@�WTJc��?��3�:~�����<T戮P������m�a������� [#f�T`�pR,X,�z�i��� `�B���c�W$yΦR6�� Y!T7���}~F^/�:A���<x���x��14 8�!��i��	Ҙ�Z�[�&��]���Ur���uU�m���(�q8�\eTn<��6H
�}��`��L���G�_�G�+h����6�����\E;�;*��`��@2w���S�"=����2���[^�C2E�P#������'��zÛ'�	������~u����N����i��W,�Q��,=����!�z�.�-Rj
I�s�a����	C:wa�R҄R	6յ�(�G㑮`}��A��S@�{�D(�*�m����'�X���c����`BD�+��9gܴWq��SOABۍ˘�wb�O��gΝ�a0&�]X��j 5^�B�Ԧ
Z����<�ld�>#L��qIw$J1�A��Q���*'O�4�kc�j����G�m��$��/
�#��1���gԑ=me\�q�Fh��;'�E��B��/<��Q�@eo�6���.�S.�@B �%J��ɰ7R��A2����cA;U���q��u���bq��A���T%B�v�j����l�]���4�@���S�+�!&��u �9��V��I(�`/+1Bܠ2�5��)�D�&�U�Fwj^s<%���A}������qݯN�_	�I��oΝ�:5 �C���E<Q�(���s7�q�Y��I}��yi|1��f�|qg"E<�ب0d���:�k�m1�����1L5z[�P	N�5�ݲ��ɗX�a��m{��ވ<�\��-��C�K�0��xY�`Ĩ�JC*i�y�%N��J�Rl���rV9ǐ
X|M��#���@�����Yk-Zs9ަ�g�檟��j��� ��n})3����]E�$a��$��٪�A��>{˛k�Qh�qo ����bEGt�ۏ���kCL����^��ZǄU�k@��Y�k��v�����DDw��
�7%�#z���Uw~J)y�ljO�R	��h���փ����`��rWm��J��T�{��h�_%���_�6�c�&)��j�X�����%�"�h.�U$��g4�Ƞp�pL �1�3;���r����k�H����M�vܒ�;��r����\sJ��o� H�ƢJL��E��c)�),�e=�^Zq���m2M:�:/�)����n<|a�/c[���RR�A�;�Cɰ繟ڍP&R���	�{��u��C5uqh�[���;�:�}$9x}<{O��CvU��EZd���nU���oC�Tj,m��2��zb☯_�MX݃��	]�z\V 8l�����x#���U; Z���!��w����w��<3x t�'��"�'����j��m� �kp�9I��Ҥ��T1���ʕD��f�T������ϒ��q?u?��L�G�=uX�([��>�Vp�\nH�V`u�VȮ��_S��יA�Ӂ�ClV��	����UX^,#Fp���V�J�ϲ=�˂k�\�A`x]����̍��!�t{P�^���gψhɮW�� ��y�{9�(Mo�~jDW�~��>Z_�ϗ�	k;�%3-[���������/��[q�F�����9$�ywZ��b[&]���+}���%Q� �[��&��w��Y6� A접uYu���d��\|����~�k�bG�ut?��顛G�iNd3ۜ�H7��%Z�V�� �WI��H������l����#�B��0m6��ڦ����S`�?�'�Ixߪ�{�_��b�$�dIyy�|��Y��Y�ʴ���4��Z����NX �cJ�GKu|�ÐAxӋ�֓a\V0���� 4d�g�P��׶Z�Wg��خCW7������#h�Vf��
޷;|1��
ys x*O?���0^��-����!Nl�GAn��w;�� P[�15��HR`"�v趔�	4X�W�{BC��)�]�co�~���T!R��|�7'�|#L���������Q��HѬ�oт�j�E���l�\�?��Y�Ǡ���'��dyqN]�Ӛ���eO*ȅU�6X�����γ�WF�՘N��fy��&L�Q~�*~-'��'��H�*D5��et6h�;��~i�o�f�G
�8#������Z�����<7�+8�%h��2:థpmc�J���a��W����ho��$�ܽ�f�=c�Y�S�����NW���UW���-����lU�L'��d/p�����59����Q�Hȩ����x�I��Y6nR5�!�½X��,��G�$�z�AN>OC��|�)��}0�^�B$�R�ů;���G|KAf���R����^���C��r�N)� ��u��
�a��جy�+�H���>����S�E^MX�O��h|v�
�Y����c��
��Q�Z˒
����0����i���i�'pL"��6Jf�����%��ġ�"Q�`1�R.6A����uS���'�9 cQ�Ù�ɿJ���'@?E�j6]�6�V���e��F���b�v@aCD��uS�R��}eX[�Sw��u��s�2��]�k ���3O�J�X��>A}-q�0`G�-�d��{�Z�@���N'5~s�/t�9��D�ELeC�?rQ,=��q���s��7H��9�"���� �sý.��]�V�K%�Z�󊥐{�����pi�3����s�%L�.ٺ�╧�q�r� w3�e3���~�9�L�ۆG��C�1�E��P��U:�� �	\�լ�;�b2_!�R�+�#*'6hg�2�Ked9̟9`��Lt</���ޣ�2R�Z/^�B2�JFOݭsϽ�o��F�I�M�ɹ�3|=���S�����|B�s6�Ys^�g9�\\}ȹ��h,�)��'����pX�ɽ��@.s��L˸�7/���<8ȍ�P�L��}�Xd�lGѡ�W״~bhi��pB���*��'?X�`X���7-��Db� �R�Hk|Q�y`U+-��m�P�s�i�����2�#��z����u�	�tK3�2����w��i��Ŝ��vKV�ĳ�x�pIC�k"��y�8.�c=Z���ΣOb26�R�D:iDI'Ō��0��ˣ��H
oߨ*C^2x�S�ئ"7MM�g��7��"�Ӿl�c7�f��%8*|���V�'n���?fM��H�}����E��C ��J��7Lt2��m�����D�PW{�C��cz�VuWnh�^����?�6�lX'�V�J���j;u���}��`I� ���=	�~2� s!�'��f[_Zp���Eu�\a{fxgWi㕷���sH��SH�jigWYF��st�m ��V���D�-��� �a^x�N��rM�ni�z��b�E.k������нٲr��0�@�);���0j�w3i'V�ӄne�s�݈���($�'�rdIǖ������]�����;�Gg&�d1�Z�!�s|��*e*�E��TJ��a�EVSf�i�?E=��g��|�t2���)�N��gL�A��:4��i!�RHpU�N:�>�Ph_�E��&�ċM����I�l�Kj�A}4�������	F��B������G<��,�*���^����ӒM��Xҝds]�{�dsn�{�5�(��_�+���Z�J�H���pR���f��ȜR�N�H���47�!B�Ҳ��p�Z۝XU��43���N�MH:[�D˛PU4&���a�'8Ū~*8���4�a_��p۽u���8J��s��>n���jZrgtoXr%ON���+��OwW6�,���p�Xzgn���H0wS����Bd~D��,⢌�k{�*��I� �Vu ������-�ke�6S��}��n���*Н�������)�>���I��� �
p�O-��x��/�>䚐\(���G<���|3����tWΡ��^)!�Sb�I�
�A܋��z�"[��V���@�ζ`4�l�����n��Ů�k���XU�A�ž��"��(S���҄������c��+�l�S��[�o��@��8m��?�8B�u~h1#��J��9��g�<�u�5`���[�3M��ӈ֊nv}���
�F�eq��6����sʋ�9~��װw�1)1��|��kՀ5�5��ק�*R�B(=�>�pu<�K��3���4��[8i�z֛�mZ�ƹ�,�j�d�F��s�_�#��s�O��pɋx��Z��q"OFE��h�	@�nA�sIn���ԙ}���*L-�����=���խ���"(��w^G��pvO㋛	��q�]�FkE܃ס'}�~��0���ٔwzhs�p~T��}:����>�h��<�`*�@�,�t�s �z^���*���:;��t
j&ԬW,F��>I8��L�n��,vtoϳ�OW$�3�Nq<� L} (��m��b4 gd<��Vc�<m����_e���@�ڌ,6�H' sV)�����K����YN�s�R��S��X���+1��(F��_ҞҘA�i�3Jѥ?<#O��Om�\�5��6�����Y�&�>����:�B<��7�9�̵h��j�
��G����5I0�6���r��i�_d]yҘ���K��Eq��"�b3.Z���rll�Dy�逆����xVC�,����Rc|�w��ȭk�E�$GE�,�>뛏pG�
����Q;�yQ��L�azH�L����Bq3e}{��lm�L���!��{�X-��)���H?ωj�[�ݹ��V16BX��_fN�A�,���񟛸�籀_�<��Dؚ?(P��q���t~]�+�k����Y�&��[�L�^%b�2R��9c|�5�=H�S�6��zdO�%�s�H��(ױ�1"d\`N � lJ��<�X����G���10m{�� �p��8�_�������dA���r��^�9j2���7!E.<��d�:�!w��M�*��z�ܨ��e�U�q����X�ªN�ʸ��x΀mc`.�����
��A�Q�+^��ze�����#3�d����{��B ϧ}�����}�y`��A��L""z��.}��D-���R��s���H��-B|�uOW��C3  �j  ��ݯO]b_�6�=0����bD��j]����s/HX&���i8�lbXp��^)�2&F٧f��M���w�p���+��\�XPyt�XR�+�3.�Y<.���f����h���~��X,`9i
�����zgZ^�#C�6�OA�e��XB V����LF�,��tle	,��Զ���x���G���8�3s�n2�,<���VJ�QޤR��8a.{��j8�g�H�6���8vf���l��
��[
��K������'���Y�3^��i1�[��)gC�Q��>�� �{Un��W)��(gN3Y�����5�vSͣ>ޯd�4��O}>2��w#�=d;���,���+Eu5��tY;>�fA�	k�T}^��ҳ��o��S����9�<�/��D69WP6��������D�[�
��1��@�Ov���N)`��R�a���O��"�Rˏb_���G�ˊ-l`ֽ3h!ŘUC}ʟn�m��>&�j�Zd]��2W�?-#p8U�D!������]��2��ĿF �mޝ��d$�Hzu?��Vl���N�7E�)��)�a�)9�<���:����D�-�G�+9GD�.�1��u�h]�8�"N��}02`X���ً���K���sV+H��~��g�Q�$\����x�z۪����?@��Ej�.�a���D�Ԍ��a��[ ���TJ#�j*h���ŕg�.|�dhqƣ�������.�vw�p�oa ��{�:�5�\���L�<p�׮���*��֍8��U�H����Wb��^ח�Y�l�}jK5�X���M��u��%��I�����=�QM��26�<���ωx�����1�
��hm��F�Mʠ�?ײa����W�>�_[eEB�ko�g)A^��9:�:�*���,]���C�#\�1��w�����W/���+5=M|�vTDz�XQ^锚`��:vnR�g����W�t�{;��:Kf1�:X^s�2��H�Z�Kq˧��sI�eP�JB����r�*�>ģ����h>�P���Ǌ
�|�����4�f3K��f�����Pŏy�j(�6f��B��r�tM:�Y������1L�?�gI6�7�T��*J,�����u��g��x���!���Qw��~���ñ����q���>�����8Ы���*�)"��s�w��k��4\�g�M�"f>��ȪT�WP�jE�Ec�L�Mau���2@$�lC�8�u�<�j"}
����ժjK�3'�uW�e���@w�tZ�f|���6s�F����]Ү��W�:b%ݑ�o�F�T8I�?P�Qˌl�ό��oPwCA���)f���n*� Sh�ھ�E�r�㛨�v7 �Ů:e�~b�)��Lh���Y����P����Ѡ�� >2(���kw/䓝}X�n),�����b돛������{��I}=s�ʥ=p�~N��eD7(�3�"W���ޏ�l����E�%N�'㹞U*
NdH�Z�l����am��h��9�����t��h�t��e��+�Gk_��x*ʖLGf���[EB���Zu�������wR����|��]oH������pz�A��E���]`=J?�#b:���z�	��\�I�K��Lc�E7����i�g�4s$$o��Ft��G���g�L�ُ<6hr�
eGd�}Z�}[�/���3����������/�ii��
���<ʏ�H���F��o�\���N7��l��_<yox�v]��.���L���!����lO	��E6�=�-r�v�u���͋p�E��?O�Խ�Ⱦ`���3��l��6����m���r�-(eCK����Ec�Ʒ`��)[nTimO\��
��:ԞD�!��}Z�w{ �~o���b�7�\:l��v�Z-��)k�On��d�,9s]N�d�i;>k��`vI�Tup�G��b/ұ��I*��ts�i�+8�m�+I[N��X���N�T��Ԕ#����2�����(r�[�`݆�Q�!{�/��&��&P&hỐ���=�k��5>)&uG������p��;J�^�؟�)q���i?V���%|j9���/iU���WDx���1[�l=�#0�7i_mr�/�b�������v2m�}?���d�����+��D�Lĉ�z"�=�.��iVLw�G��M�����C2������i�Rs����Ye/���@H�o�Z ��<T���I���UE�4f1��(#Ԯ�&7��%2��-L���6w�P�ܭ+O�����jxAG���x�4؇������Z�BS7�iʏV�k��Q���2��\-�Qo �NT��L!MB0-�`��_򑁣t>��Ӧ�DB��S�=$�_��ࡐ܈j��ͦBӜ�$�K�FW,�_� w����~�u�mW�/��ִ  ���54�]��x�d��M_ؽY�+���B̨pCa��ұKD�[�įG����~��ăge�Rty7���u
�#�AlAi�_���j��۰�pR�ξw���cҖ�q�07��F�Č�E�� ��Z��Go�J�lT������ID��i���$��=����Q��.�3B���n�7�Y��p�D_������p{;O��G�P�q�K��g�L�Pم�]�m�h�|���D�}���A0�$�jg��h;�eNf-�ӭX��Rh��o�=��-w͘g�j�x�C\�F���<�kA�gp���|$Kө�3��j��ա�cHh�������,�d�+kW���y��ӹ�ri�q�@(~B��s,�֏\�r�^;��m��3��f�WO`���E40
�����=����էc�P���J���%m��md����H4�jRx�c.�X�LDc,��`_ �À{�'?�D��u��H�;�k��u�]���*=h�ܑ��2�w~�X��r�F�u�[/�U�-���Xo��FwD1R�B�g���P�Y/=X0d/UCe�N����4Bj�!��d�K�)�o�������13�G����R�w��3�����f��+t"gS���!�¬�I� :���4 c�H:��5a�S+f�^=k�|�5�d6E��.�ؓ'W{�l���,�c�F��)�桶��W�����ơ�R`�B
	�hl��1X`62�k|�d
f�n��b ���3_HgTWM�����O�GlD�~��#���ƮĆ��SXR4�:Ź�
��m�����QD��+�̠ ��Xe8j��U{Z�4��⼃(~J!Ϭ' 1��O����Ö=f��̓�U+�%�~7�c�a6��E�@R5��$�?t'��/��P̭���Cӣ�=\�^�QZZ���V�T��i�7R�/���@�t�Վ��׼)&�h��*��=��ݏ�,�!�I$�L�i])�dD����P���H�0ڟ�?��l��b��Xv��d�A��A�9+��gE���l$�����r"�k���Ǧ��P��8(0Ŝ[9�0 � e�3��8qp�4��\=a�uK��Fq�\�V���4g��S#>!�7f��#׌�줯.��t��x��!ϭ-�K~�+����Q]�����!K�_��T�(a��p����Btu�kQ�Ί?��cC9?��D��+�D@������l�QF���.�T��e [{$|-�ey����^L[��~����p�>��e���^3�U���cl�3y<�/�I9�����R�r���pH���T��X�"�G�13w�)b��O�����s�,j��f�[���r ˓p�Mx��y��2��`��i��NSc[a�m��I���U�?$��1G���������i093O#�x~�:IQ�I�|U,�E;唥_3a
��E���PI��hCŝ�Ȳ��W?�% �����l�<�̮��)�E�n�T�Y����n*���?d�n&����K:���X�Y�\h���?����rL=�B��6����v�aP���	o��E�k�9d�0n{u ��1��dP1-:��f�z��X�ݷ����P%�>�Շg� �6M���3)/Y��@*�c2�H�>���7�I
������P 1�����s����e���`W�
α�˦1�H@Ɇ�q��aֽ��ʝ�i4'J���-�f���!iԽ�T4#��勤��W��
&]���h�H��C��$�2)=I�v1�W�P�<!g17��q�Ն�'�@p�ZŁ�@�Ԉ�f���:�7;����`ڵ��l�)2�ǚ���C�p�c-󺷏�q�����^��|~@��ɢ{ٲ䧠^���#�EE�+��G@�����^㋝Pcy�azTS"y7�GR�,��1�=��p#B,%����H~����ő���o:��Oİ��Ժ�{�S��7R���f�+��t9���  k��4���khWQ&�J�Kj�7{{�X���cPA�;¡2%���Pн�a�\fs
�5�.������H�9s��y��d��KI�zw��)	\���y�/��+�"�O���L����α��Ś;;έ�c̬��&O�G��#��ᆗ�I_2�̸S�}�> �:?���i�^P����W�y�Y��rZ?C��̖k�xiUQl".�b�JT�,�s�O��U�)�����p�b�~�⮳��,[Y�9�.�M���$���yz���U� f�ђ�4V��A+l�����y�Q��Bǹ��\���DȪ�x5�$��Qޟ�E�{���d65v�	��)�2��&~U%��R&���������ei&C�uB5��5���4����3|Tl��Q֗�{�B�
����t�� ���y]��]\y0Pi�߉�PJ���>9�6���-�Du�b;6���ɢ��&�}h�0Q�T��Z�����tYTl�n¼�����e��N.9'w�6F�����998&k�<�G�{e�mbHͦ��$�0(g�U��Y��@~3�x,Q�� ���^�8��-O���\��Ͼ�H"XB��Vm[�3�D�����N�ގ�!�'�A��?R�$�M<!�k��̣��3����������7;���`��	���NE��Y�sM��q��<|��a�4OV[ga"Ă��vE�dӔ�]=7�RJ����P-C$���t	����-�����s��ù����E��1�TL�{��5�K�5�d�/���IKl�)�W]L }���Ѻ�
wqfah��Md8m*�紿�[��\:��5��Ni2�b���fj乶�#�1������ڕ��[G�Й�������EH(	r�ot'\�1 #!�*��ii58���n����v�-���h�N��~>�!�RRV��p�5�`����ɼH��N�>�RKyF%�CP� ����ţf�sI�u8u����ϩ��g��Q�S��cqrgHX�s��2��d�|��,W}=c{��(u�﷠��!3H�~�uh�Ҕ�9 K��3y�Ra�%�f{ҼKV�U6�h59������
����Bw�	fp��W� �P�D�"!#�ʺ@M+GDZ����2��j�@�98�C$@���B[�_tA�������F��k�M���|O4��M��,?�J{[�_Y+�E^�m~N�8��m[�*T>?�I�^��rR��~�ղ$P�1w�oŁ
=�T1��8#�t]���h�Pf�,���.8p�����}t���S���:��~(��|��	��Im�8J�΃�y-�[܉�Â����^T�HX�/��au��kk����,�b�x��>��#� �_l!�PIM�D�F��uk%1�d/�pZ�%���
�cA�t��xv������D����6l��r,7<ږ�0��H�&�Ԁ�:�/X��޼��I��N)�ޮ��vr��#��A(��������g��8���(N�&����C1+���|����\�"�T�v1�mB�3�;�2�9���ᛇI�a��yi�cb�y�0V�Q�\�G;;Qx�i�@z����|Ƀ�ǅ/����.�KI���q4���w�&��e�h#%.
j]H+���%�`5����E��L[Re������`듿Q��MaI#�/�+(���bIO�c�1S 4������uw�������e1�[��-���=���)��]g�81hMF)i���A-8�ѭ\�
��IL�NZ/�m��0�vfІv,q�e���v�f�J�J�,���`�t�dc��8��JT�,[�eWy5��$�A	����O8<?���Lȧ��d�Q����r��Q�����o`"g�4��[I����O��F^��.��5j�p��M/�Ս�8s�* ���/e��������f���$�۔�_Hh�d�,�z��!%!6��[jJaJ�O�~<���u"{�F�|�������C��NzI�Fp�M4�J�$F��P��?��u�}:F�&�*�������o
-7���qbH���'/�ϺH�4F��͒m˩~_ZǨ?��LYеXڢk@ty%��{�1B��F�M<���h�`�`KS���V�L�^�67��m�����#Z5e�" �v�mѩl�|{7��T	@�@����4�Q�6�nX5^�@o�8;9�����4�f�Cj9P:���43����ĬQ@��PM/���0yvz��}�s�	[�YB�Bl ј����|�,uHRI&n���C)ќ�[J�j�<�e�i"T��2Ţ����@�Ԅ�Y��������i�V�����n_��������^�bvjtb��,��8eO��0}�ۘo?��+�Ԡ1����:&M��B��Ň�����`�7M,���d�=���@��_�?"6�a���M�+��˘8�YW߼�z��+����8�z������5�Ɂs��!^�n�/EW����>{"�Nn=p�L�k65�RP.4D�×u���
31��,O����b�h���Q�DN�S�ERa4h�j�z���~���脪�P�����Ϟ$|����+*Iw`*F��t���_�\;k���%d�w�Y5��^@܏<�&̚�P�8hs�ny��ΪN�[Zɽ�w��R��~��"O���$UaE��c�y�7����x�ᛂRpFď�~����i������9lT���+oH�t����EVi�w�s���D����4?�l����X��-�ȵ� ��ۺZ*C^�-"V���Lf~�O�=슠�8Wg��e���v��������l	~K�I���J��R����-�%c��܌b3= �hDylq�,=��k.��z��G!b��p�!�]hF>��R]e�������ff~�*X�laSr���$�5ǁ��/+�٠��"Xm�Q[�9��r�g��@�ȃ���E�A�����>-�����7�iab6���u�0�f�͊�����~�ߘT�Π m��۵�h� �V@ ��*g�=�Cb��Oj��WDX������0mk�����o`��wL�#�P{�6����X2gD�{}tإm�:�dM��F�N�eC�?R��/^��/^YZ �uo��Q�ٲ"4�M�uj9�LW��;2.��S�zv�)d�M#
!����JA��g��oF_�`����m���.F㐎�1<WS��?02;�*�1I%�B�[YڶR`���[���d���ɶ�`�	oE�[9�w��un�i��ߴ��6dj�P��2jxts�1��kv!�hG��އ���{�We�&��⿸�/�ހ�,"#O���{�#�'�)+!A�
EJ��N�{�Z���;�����f�}q\L�LKEu�F��l���h"QC
 �\l�.'{Y��ܣ��1-״H�z��5$���{ؑP��=fr?K��"��a�^H�Cy]PQ57b���Ē�j	s��M��;"[��H��>FF+ň=T�5r"�3@7 !��5���|���m����c�/I�l�̆2����/�܆�<�|K��7�L�R�����7�."�~�80�:�p�X;��>l{��IR�W�խ8���t�
�V�u��\�������jeә���g>�����8��P|훧 �� <ͻr�/o��P����L�����%q��
N��B��>�X�IK}U&�i�KZ��"N�@8 �}<�:�x}���#��N����%���O�XL�4Щ����<���X$OH���[�+!�aR�=x�L���>�ʢ�P���+�L`�7͢�#-��.{�P�\���L�QkI�^CM���XBt�kj��O9l�N͗b�d�t�O�i�����f�����S�F;.^��N����,�����gTٱi){���$�8=\�H����x���{kV�NzYi/�����_r�����q�dg�����H쿣��>,Ҝ�{E>����z�L��E��E�{t�7�_l\�=�x-�b�Y����ڝ[GRS���m�m��iSJ�y�4a�R
M#�S�"���yzE��DH��ɪu������Ȝ"���z�sl��&j��{��J�Ѻ�H�P�<�Rɣ�7oz�)Pg�9c	�l�ELS�jW}UG����r�jº@r�.`{H����6�~]��æ�r֝�U�RE�ҽi$��LS���TP���b��4�F�>&�X������Yq�PFF'���c�UcV��1��8Nq�����lǜCdKg�|�E��Q�˄[cOЁ�5!�?@\	׼�%0�'�3��X��<��wL�����8(�Z�7E*˪�	<�$!�C%�|�Pr�����ՙɎ�ɚn�����G� E(n�� ̓���(�w'%9y�iX}��
)��}��YR�`�,��]=����-�
t)��ٮ|��D>��^32˛��ۓL����ם䧮�d)��c�)B$�2/}2�sQ�g;��C���M(���k�*�	]�ς\0g�攠W��C�D�Z�7����`}X����΁=���}g(L��x����4�o�p4<�Ѫ�~Z΂b�}:�K���p����^=+y�e���H-�Ț� (B�.�Ƣ�0��C䟹Y(�*�x�H����:�ԑ��$Ȃk����r�f#�3|@9�!�a\�����w�Gn�S�q�=w���}3}�SQ�-7��y�.��m����`Glb��iF���B��N�<|#�S$b$�5C���t)�w,����֏��lOp5�Rc8D���>�v��ÝzY8'HP�[:ǌ�ҁ�ws�y���\���g7opLPZ�}R������f�i#�Ư���%t]��M��z�s%����V� �*{/��K��cl����Q0ӹ����@<�pF�Զ��pt\�-��,��M�lA��6a�+�P��䟴���u�c!'肭`a����β�� ��E���-	�����o�B%j_d�d�2w�	@5:�*��$D~t([�aV-4�t������>$$)<��9f�YQh�.��VqeQ�.E�.���d�����%�I��T"_6�_���W�LU��e�B˪��C�P( >��iy�B8�Չ�"v�������+K�������PW)^9QL;Xg�f�+��7]��`0G��sr�U�¾PF�S�������t���g��A�2z��CP(���ٴ#���πf����v]弚�������v�EY~�Ř�G��B����`�xs�h
mZ s���;�c*<����!�5����8��+OX��^��<�E��c"���7��va���j�~�s��u��$�x4�+Ú)Ub�q;������z�߇&�ކ�O�`�p�y>1!f=�ʘ�	�ȸ��5k���M���}�@ݬ���%�D��q��]�UN���N���?�zP���h�C�ur�5W��O���6��N3,�?���&|�%�ﬔɢxW8`��/'~��tr:�kCV<�Hʾ�E��������\�����S �JIr��u�%.ǒ���rv�p}�+R�#�����Q�ց��\~��a���r�mH����7���n_�t�H��)k��_#5[����J.Ձ� ��3��m�C�<}���4�=�C�-�Y�M��p�ˆ* t��ʩ$�{Db	*�u�P���8��W�ؙR��eQ� ��Auj�ph���+�i1�^�C&�6z�3ݡ�`�J�>[�Y���v#:#�
�!�
��Uȧ�Y`�\�6�FH��_�>Y��!�i���wպ���+�k��<�H��r����7K��3�e��JV��5���	�J*��R<�*U�yzm�>Җt�q����_�1�ThP�����/��+���x��� �#�6��D�d��P�E����D6��8KUn���J�졶�S��c����}�F5�?���f��9c�ј�Pc��u�p�2��X?����U}�po�`�!W����|�S��%��*3b��3��!?�"Z̋�S�鄎.���8^��>g�ʝ�Id��#\��p%�Zs�.)Eׇ��S1l��C3f� }4�i��dJ���F�>�J�BE�*��vY�?8m�{��e�c���!�:yz°��]UQ���� ��  Ż�d��82����� �R���@
ڲ"!˕}S�D����O��K8F���킠[��qt�EN���6{4�߭TN�&�v�\��nB�e���;�l9" yl+��J�k]%��
�-Ϝ8f�N�y���|�2��������?�I����&_��%yTe0���͡L�0yk]�ژ��R���@ă^�U�ك�?�c��	�� ��BԴ�\��.`��^%3��:��oe�(Sy��<�dM��H��7�cA2$_�o��W��a)P�ת�c�d�́*=-87��W>�1�2@������������W�'��ѽ=���.���"b��i~B�0?��i[Oq�ߐ&��?�C$^c�q�v�{�š����iW)G��潄��u_��G"�Z�F�����i�dn�j��'����[�dw�'����4�G�<f�gT�0�x���BN�`��Ol|M@����O����Q��ņ')�pq�_�09�R����o\�
}ͷ
Q� :]���Et
8�D*;�+�Eˎ ΐ��Q��'v�JB�!����/we`[��̤��ݑ2;)�$х�-�Z�@t�hE,`´I&؏�Eוtډ1M�4Zw�E>���e�7CY�ݤ�B��kz)�v+��ZQ�_��[L���}!x�r�t�­;�܈����(h���v��8I��椸�4;�ՋJC��*42�ʹ�+���#���y�i�b�eG(��M��u�_g�O�٭r�O���h09i��޺���G�.-jQ�W�[��d�E����)��5�c��-�5������>e6	:>�nV�勪��B���6U?'�m�������ںd�������(h��� W�)U��Jw*;nW�bg��WTwLqݗ���4��&1:���^���`�r٥.��\�	.��#��;;Rz2�]C�|d=0饄կ���h�^��9�G�A��'V���mZjJt��|�-v�VH-�ʈ��O0�?@E��<{��?��O�|�W7x:!keV��ĸ�Y�G`�Iޭ�Ws���@�G�;��VZѝ;�N@�MZ��0:�#4 ������z��e����<��cqDyA`�c��v�����Ӷ�=t^sd��;��v��y��3#��9e6���b�p���b�"��̃$�86���`��L�;����=�L�N{�K-�O�Q\���Aҁ��w�BR%�2(S��k�q-u�/c�J!�,�w�V���'�U�����љ�Έ ��m�%��:=�p�^���g���鉵�)E�D�k *���h+r�O�������c+�;��d��H1Y�H6Bp���*����J�pxL9F]�*0p�4菁�/5/��D%��S� ��uwMx�G[�T�1�b��
����WiA�7�OdV��J�p˖C�-�����:|N�tQ��[�Y��G�����,ܹ�Y�NT'��R�bfE	�=t	Nie�b�v�_LBu�[�㻒!��RZ�t<v�l��z6@9�@�w����=�-MI ��i:V-���~�2�&�, <�(�tنyL%y�K���fv,.�?��M���+�W���jٹ�Z��1L��!��'��k룍I�uX+r0��������o]ndMV��g� .7�[Nc�1�F_��C�̧)����,���si�$D�ОUֽ�p�P�����)?��"�����n	�J����^�]�|)����`�no:/J�[Lql�0�_x{)Z�n8�s�`5�czx� ��,sI�31OVYt�Gb�b&8S��GZ�V�x(��E�ț7�%N[��c,>��|Vo�t.�f�g�Gp @�7nls�L`����b��Z1�x"*﬽�e������!��3�����$@A+���ڪaE��sܕ�`1�ش!B����j7G��r#̂@��V����7տY�`O�wC�����	��2s��Oeg�[��
 t2H�`w�l۾�`�c��ꋫ�,c\�*u���Y��/�2�8��A�䠥~Hٕţ�5Z������4��4U����X���.����ii.O��᝼���I7�N����#F���Jh�[��}N���<�݇��IӠ�,*�(�jQzf6SN�6arB��|��F�w
�5mpt�<���W��`|��֐J�&��U�$�#�}'�ZF�+&�:�n?���:_"u�K�0 �~ۺV�iL�$��CЯkj��^�)���;�X���،��.�o���I��j%�zU��d����\j�B6S	�(ӡ' �<��ceJn'�v�j��K��}F�J���j�"��L��1-�z�\�g�e&����O�i�"��'��U�'ꢊ���c�l0目��f��U�]�e��9R`�cB x��R�,�zש�s�յ_��	\�5|�>�MSź�KuU�zb�Ȓ��K�e�_gy�M�=M!`�m��|�<�����E������f�'��hR��-�y���k;�A:C���d�|� Xx��'T�zA�����@�3��6�$���P'�*��a��C�`n7,���a��K?�_�Xl��5�ֆ!�ܿ�7y��助�?x"�h_�{�c{bA�"�Fg6Ka*�i@��^�Q;Qh���VŴ(l��	�#j����͑A� y�?>BBX��+ .,��;���h�h����Z�U�+ʾ]�G7^�i�Y�W��)��v2W�6�*$V�~T�<���D-ںj����A!U��S5nA���G�ԃ�ㆡ晳�'���bF�GE��0���I�X�@���9* ��n�7ߴ���>��p(�d3H_F\\
�E�|��.��ϔ}�l��+	JmRw7��-�]�����(q:��"0����i����B�.t]x¡)&�~��am#,��<K��|�	�-R��wӷ��!�{7-h��a����2�V�_B��i�
&�aS�D`�wH%����d���W�ZCTqHQ��Tx$�늁L��n4��h�������8�M�[�29(��)����v*�o-��R�!��@h]��мsr��=;KIn��<��̯��s���k��e��R1֮�
��I�ۿ�[$�p>��ː���O��;���w����H�^1���~��y�&`��0NqZ5�4^�C�����N�� ���EW-eN;�j�N��\���'��H���tD-�ֲ®�]8� ��4ٹ�M���}�������ʕ�-��mD8���dgC�3)�
��<��q�ؖ�I�c�P��w���=���,��C�G4�C�K�#����W�縰^% ���Rث��.َ����Eԥ��e�v����~:�ig..�;��Q�N���W��a�V�� �LiT=�^-1p]e�MV�e����]/��|���"�Z�En����7)�N�(	h��k|#���+�����Z�jUţ�\�����R��uDi��[����Aeo����n#�v��Xda��%'� )�����K�BѠ9`��!�W���Oe��ݖ%�}K�W������Vi���cA�.�5��`��+���H�TA�&9'RPJl�c�إ53��D$o�U��K�1bR��h?1��x�����{�}��ăd�qWXV����:�{�q���x���W��%�D�B�V�ۼif7��^�`�Q�τ� �澇c		/T��-�SO�OsG��/y���c#U�����c����b꿅,������]��~i�l�{�I|�N
��:Oj8�e�.�[_j`�0��4k`�+ܸ���s�+!0l����)U�׫�a�<lo��y5Ie���F���
�ڽg���}ߩ�M��QE�G�{pWY��k7L�1�$�6�7-�z�йIYUy�Ն�O%Ơ+�l#���}γ�r-�1q�tF��$��&�P��1bS'�|�Ѝ;��h��fw'��X��VLby�E�R�PaF�mSu�� �w]M��<M�m�� �0T�/i��T�_
@�[^]���W(\� `M��|�@�)3b�Ε+"��F��A����%�s�ٰ�	
����^-
I�|�BZ�@�Y�� WS������ښ���BDC,����W�t3��NP��aݡ�P'�m�c�m���_<�z@e��牤��ž$�{�2�ɹ\��\]��*����[@i
�458J: ���U�ڭ�4[_/��֑j�X�����a&�M�@b"���𡋞�z�@����7Iþ����Rs1[An�=�n �)��	�ю y�-��xV����8��w4��_%�?d�1hw묁�zѕ+]����/˜emЏ�7P'�Z�A݌��ᗇ���Y�-��v��wD�w���e��!���5�C�X)��U�W(�03����$~�����hѕ���U�O�.&����ci���z���9���/m6�q��g[�35--�b��Ad �<�`�9���.ҷ凢u��t�}]|�p�ϰf�)MQ4RY�*��Q���2�p�A��cD�f���X�tn�\/s 7��:�!+�����t5hZ�G
��#2k	μ���x.y0"�YX8So|1YO<k��We�@-7�諫T�uZ_����ýA(9 ���y����C�i䈚�����۰�57��j�Q�׃��*�dm�>�^�w���������=�BS����+��j�^��1�\��O�=x��j�����DK�U�H���*¡��f=d}���p4��������S �}��vQ��ޑ��1�
^�nZ�9������ƽ��'���z�a�f�������U�ʶk�F)r����d�=�^@rugaB+K�ۢC
�u�w�z�D�m��|��0��B�WX�i��`g��!��&D^���l#h1�,�Gj��l�F'�n���\ۘ��?�S�Mmh��JH� %:��r�.�yb'����;]�d@�ɻ���˲��O����[u7�(z��.���8�� �.���6]�M7�;;`[GZ֪��19�qj���s(���}��$↋#b%��� k����r���C�����{�
^�A���7���Y"PNK��~ ��+������a�A����X�7,a�Z��8���QAD!�Rj�N`GkI2��9�!��;1a_4�I����u?�-G���(گ��,�ɽ��w�<�,�[1�X2�*��(8���v5�̺p����~�[��Mc��NvS��ӡH����X�u
pEB��_?��+��6���+��2�ӕ*.�RʶW���-r��25~>����³�d��4P�ߏ�C��e��X��kM�%��'P2b�x�ﯺ�(��
p�@�p�ݫۺH���{w���%��R�|)���ȣ��z�����o��x_���ڝ`������9�~�W��B�QE�ڠݔ�J�l�+���kH.��O.E���ǰ�l��;@��
�;���/���V�v��j߹k���
Zr
���׏������٨x�tzIT9�
 |��/$̑��AW��N��?�s�`X�2�m� ��=}|>X�蒟2ԩ�/��r%�|�ᨆ�g��d��PMêA�Nr��6_#��˕=&���	���1�rZ 4��G�w�8�9,A	pg^�����M��hZ���@��*<�l҇�*0ze|Es�ϧ{~�����Ky8�xX�8D��u�,�j�A�ao��Y��.�Y5��MZ� 71׵�;fŐ��7T�)��]T�ߚ��s��%� �87+��=����<�/F��6��-ҼZ&�[��x��,Z�m����qB����]�����.#�6����xe_����H���J��
�6{5�[�[�q�rQGm�!���4���>ڭ�Mj2�%ޜ�&T�����t�D6���G �����\���A�����ܑ� �3��A��=�JY���N�d��b����rCkA՗	,5��U ���lm����Bn�S���E4��aE���� 6�w�B�2/�VD�@9[q U���7�:~�@�X�G8�N����풃c�j�����,>���1�/Z�\����@'��i̬Цɧ��`�P���� ��hkg��PA� JF�i�֋�J�e&�A��(�ƣ�%ҝl��@'8C�W��8���(�X���)��\���\j*ڝ��9Xq:�z.�6A�⛭Fq�-�U�FG�BȻH��3�����T���;������]��>f��T�"�8b�����[JH[4�u��U�+*C�4�f�:�̙�Ɗ� ��J��t�`���#��&�sY��Z��=�ޒ�ǳ�
�v�0F2�Z#�P���#�^��𰲘�5������۾�)P.��(F�r{���4�i��`�Z�h+��m��-�C�5�A��V)�G����]�R�5%�dW��<񝱧�laZJ|��o���&?]���z��ٯ�.r�mf�#�Z;�삯o�hȢ��$��h"��aP��y�J�U���mm�'��f?De��ʥ�#�W���!z���_%����!�!hy�y�ɐ|odƫ���	T�C�*��*F}e	q#��oY����[�c﷭&�4�#2��I�Z������QJ�"JN����5���]&�*��ч2��₥�A�bh���n�vD���� ����4p�4WNɺ����k3,M�jv��0�P�*i0ڏe�f�X��5 ��F�=slߕ~���qt�����������5`/�ێ�;�$�Y����I��ξ������ȿ����h���]!���_�}8Yi����>�ίnr���aŇa����MrRu�T�����s?���P��G������~�*�~��B�aych��*!�-�q$���9�Ѧ��|Z2*[�WE8��0I�뤑sb/�o6�-f�}4=��w-�Е./
���g��K�Q8��LE �1=]5e<Rh�ฺ�:�׶X��h��
Z�%�t����Ԗ������wQ�&�J�폓���.��J	�,��)����&*i�D��ϓCן5z�Oy��Deoz�ၢ��G�I&��$ @��վ�xP8���^^�=�6�<���5`s�U鍻s��R�׌�tңz�/����]� �$P���_^��_��e�"聆�(�ݍ�J��`#,���	��z�}���i"�>t�<4�r��*(�b�V��8�_�"�߄�a��C�/
�G�@�gU
�޹XA[�ssu���k M� $Ł��u�VŢ.\����j !�EOʓxc~g#����$�m_*�B�ʌJ�"o�C�y]��岤�	�,@���Z���@��2�dn�������O$��k�e��ve�_�}��ܙe ��v�)FZ�JۅO��Nk�����#d�q���ǜ�Z�)K�oO�u�I��W�t��u�I�!(�W��;�������/����{O5u0U�P�t߄�м	����I6mx��'<Ԝ|ڮ[��_(O5a�P`M�i$�؝ҙ��ȡf!�ؗ,|�XD�X�NX�R�ح�������@��GL]�)�wɄ�+�:b����m^�r%�X��J���ֻM�f6ZO�WX�	�!#�?%�b�<5ʂ���h4�6ក!Ӯ[,�o�q���Z��5JD}h8W�E�(�T������Lg���Ծ
�t��`���]���h�ƪ��8��'�� {��y"Q_?������	&Mo�o���l(]+(@��<�+�Y&{q6�a�)%���@	'v,?�{��pq��,�p����n��V�J�A};�M����^4����e]��3L^��"9�;a�2��E�ͱiQ��_�9.�y�v�a֮�џ�z9]��-�.^~�o�.+�$v�2a�~���%�����)�+���	��ٝ��_�F�+>��.�Mj/q��uV�%Gl3�H����Z�J������كE�x�nzL2,vf��epș>�u�KUӍ�v����:n9��|�2���8�cb�B�u���!?�y�뾂��8r0��)|�� ��O����I5{��a��W�a�"���u�5{��1n���=��FR�r��Rxr�k�R���u��`K{��4XUP�ܨg"٥�i���l,\n�H�N�'��,����6�G�Ҏ�
}����4�Zɜ�l���#�v�n��ԧO���s�$&g��:H(b/��?��9f	%�/u򲮼 3~[��5�NZ�^���s�Z���X�9���aƵ/Lޥ�I���/��r_�E���\r j bTE�Ƀ��A80;���<5:+Sz�&�;d�|?��{��@�*���jn:�?��F���Y�f��xUՌ�Wd�`�?�zfJ��Z�7�hz����PSg��1z���5�7(`��ԒfI����F��h������.�bQ���M�.w���x"1d��*�¦<! ��6�˪��}�P�y� ��.�N���⡰3�;cl|�z� �N�ak�S.q'�5�=�{w �w�|�:D���S��X�0��쓳l���}G��'8ۺY�@g�<�O;z�!��za��X��?�����
�CӜbic^�2b�Y�m>� D�������r�.�T˚Q�?')���'���c�V&��1�ǁ�]Oo�L�PPm�5���P�AtB�h9%�F�I���V�Z���>]DR�dtIi* �5�P�`<�:�c����ف��D\�,޴�\�2i���qqj�����>TM~Rt��a]ĳ���1C���|����Kw9���|��}�!�;o!�5\ʰ��8�U�}W
Y�c�������u��era�^��Q^6:�|�8�,7���/�a�� ��H6���2d�6G�>��vדtHѱ2I%z##���,��A�;dF;j#�jSǺ'�Qs	:��Ƚz�u�0���,E�*|�<�f=�N�-x 's/'l#���6\�������#ӠR���>
 ek�%�8�}~��\e�����c���?US�)�S����� ���]���"3�������<�MQs6Vh���	�4-�+[��8��1h�;���u�OC�i 5�[_A�|Um�������$5h˪��Y���@l�Y�m���,�[�C�9����+�%�2�ƀ�_q����q'�m�"*&�B��sE���E��~�.K)G-�f~?z^`�KջՂżA������Q>�q.f�%�ou����$��-�X6�]�������q���s�N�O��<�����צ�E�Q���ʺ˂�3U{�B�a�<����L~�3�NO��\��p{�E��@�(���b��w&�O�ªn��Y�ٿ�k��Y"���v]���Z��vX�@m�4�����_��t�\�$
1�6V՘�\d�U;����xL�ݺ�O�q.���i�
��������rK�f[���
k(���%؊��x@^����e�?��N�`��0!=	��#�s�z�	�';K(l͊x����N�E��tZ/�`%��p�-h������հ#�%߁�	^�Ok�yG]�Z{����i�����+�&ʧͼ�;re8�(�$ Kz��P˫4H�A�{Z�}��@�C��e�"���1����L^`;UV�J5�*$�`;lE�Ī�%z��kϫ-d�#w�^����m�{J-[^&��s� �N}�=u�o0z I@qX�#	z�9�|�@���`ޠ��@T2#3�iI>���=�|�����~�(�4l+ ��吢���i�/�aSK�^͡�������F�3ﷄ��[������')��yႱ?lh>��b�f��>�������.���O�mԪטe�Y�ko�3u��䝒u�^!-�;�U��B�K��x6[5�ܛ��9ݓcu�̒I���7�ÖD7@�Il��C*ݐ�������LΞ�$2<}\>�f�
�}�b�%iD����0���o�#����`%-q���$fD����H|X��dS{r��.�$�#��0��	4��1�,4B��26�{43�'.+�tX��~��L׻�!�zԁ����`өeP%���!���F�OV|W����0.t��H?x|j��ۯ\��q$�6��#������W�._ޏX��x���}$��!�ˊ�f-��m�Z����7�U�&Q�0�^Y�}C+4�V���8OFv���PIt���b
N���+sE�uo�"�-)��*פ)t�&�/�9[�¡s�����jF����Ҹ"?Lps__>��hE�`�F�l�pڅ��7l(к�@�\?;�S��ˁ݇���hW���Ba}eG7���U���pŬj��� ��j%�'~D�Cj��LX��T�*/�t �U��d���S�v��O�E?#2�����ϵ�'��UD˝75	�H�^�݃"~��������4+�	#�3��M��|lPq��&<'Щo��=
ʏ����_�J�T��B���ۑ�c��)(1��%U��(�H�m����b������6%`�jQ�#~����5�A̓1JE��W��5Y[S�I6$.Sђ�Ol>&��@*�l�*�C����7��a ͞��+J�c�`r�{���a�ҤFgpj�	T�3�/����A@÷�`?T=�?�4=ǧ�-p ��9 �e��N���{۵�3|<ށ����M<�م��,�*����m��[�	���AX5�Z�H��=L�n����*�l��"?9`�wl��I�j�gA��BM��H͵�W��C���� �gsO)z���c]����Ƀ(SpcyM�3�*�;Af��!<� C���2�h���3��êfBh��^��vD�R�޾��̑k��A\�\�ozM;�F �؍����D�7�I�k&/P�KX�������]ۓF���<��Y4?���1WJf�1}n��fwX"I��?ѧ�ѹ��4B���l$??�B��%,�bg�ZC��O�厐<*\F+#O�?㭴��l��pJ#�g��4S��:5�<T�pC��������9s�����0��<�y���Uw�΂%ZDlX�C7�^��RÙ�y~1����z|&&(�et�m٦76І�ğ��)�x�Jl-�	@�&ᳩ�xT0�4B��ӈ��H�����ɦ����-^��ٓ#��:�6����7�����4�����u\�l��B��v�����I�%����w����m���T�'n��2{��STJ��Qo#\����.W5욂��� A�_�d����2?�Ң>�.Ӻ<hv_������m4S��S@��u��@~�9�J��=�65g�Ő{�֕��4�&�����;��>�$�N�X�����S˪�uol5D�6�����ә��8P���k�W���)v�m��3����|O��3�;���C���;��c�;X���������e�7�C���PE�)k���"$�t��"V�_��bɊ���rB�� -�2�S6����"\MQsI.@�����L���+P� �;޹]w�h�����Y_Z��m�F����o��:̽{W��Ix��z�w��e �UXq=T�%~��ĄU��*�<�y�Qok�� �>�G�>U&~[U���B�w��L�Q�]�d�M�f=�maxS�s7E��J�R_%� ��!4}�>%���PDf�C�`_�,SB$�7x�IN�����u�,�Z̩|��Y?�j�À��C4R���n�h��G<P�W�՞l�}�Z�`����l�Z�^s4Z*~�?2�e���!�@k��O�J�h�\����A�RN�����V��~�.M� �D?�~սZ�i9��A��N��p�ߏ�A����s��5l�FW�"<&�V54x/&�f�`��	p�q-|yVAAiߐ�lt_<��!��l�.����Oo�w�l�<$�׉k��8?�i��8,A�Tؽ�03�CֽaN톪����XG��H������U_�*h�m�-R��R�Cx���;�*Z�
܈�ŀ�at�P:�N˧��pf]C�P/�\s_��?�e.i�Z*�	s�Pu3 ���\a{	L+W��p� �!�< �Rd�����d����=6g���%�����6���B�:�����e���ީ���5˱P�4��F��
z�Hsz�w`�z2�aw(}@��V4	�P��h��=OI�9~,>U�ɉg~�Ym�
WN
��!����8K	Ɏ�n�/�E��=��E ����4��3�L�z�R�J���;���FgLc2����#���P�W~�/����78\�K�
fT��r�H��
PA����!`B��Ɤvq��CN��$�Awϝώ��'�RE�#~�[��)#� �d2��
]ථ�D�:g���Cw����P�<�ꢴ�A��$ĭt1��W_W�\3ֱ@�hu��B���lM�DhO��S�=���A�.>��mHPe��D���cL�ddV{@	����30J�5^f�*���+��,�Pi(J.4�������yy��e���h��6���H#߿Dy�(�i.�cW6U��K��<1�S'_���*�h��Ë9m�4/ò	y��v�i[�1��V�����)��>��J�9	��B��	�m����,��6M�^�(M�/�ԒKR/��O2��>���2K�U�Ϩ�
]�O�#�ڸ�
�H�"6;%��0�m(�Q\��vG�����:\Wx{��Aņ�7>暺*�=�ŕ�\�+FGv5.�T[�%m ��E��Ãs@Ȗ���{e���Q�|O�&�AY�JK6A����!����
���:90h@i�xfa{K�po���2Mw�]��͞@��}5a�A�^�dX�$��F��ru�:�V y�e�g������ۘ���⮖�Q���@�qx���趿Q�U���Ko�茘��}��Y'd�}Z�I����_���e޾��s����d�4 �Ĺ�#?J�����YMÛ껑uV�#�suۂ�~W����DԤC�֔hۚ��V��T���\Ķ+����?x�PM,Y��֛Y����ɉ�-k�y��Wnˁ�CӔf��I�x)کw�6u�%�4A�/�yc��P�!k���P����i(0&	��g� >b$��D�+��׾T�6���(�+�,��y:I�`�D�d3X����3��?���^��R���\�$e[�6I��A���OH�b��0A��~�,���@�z�C�eeS=��-��ۄ>n��I]��̋��9��n��[R��j�sn��>ܶ%n��?M϶:����5��U��U�=�Xfr���F
Pp��ج��$���@f��g�s�}�C���C����m��