// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:30 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UM0uxB7uScUab3suD7FSpa8B/EtTLV3AY1VqG121spPr/Pd5ZAP/HU9KP2nt1eW9
jESh0mInZ7VV9tR5lRzlKSPpRNNxlhSL9+dvzkogx+A0aF6qYfBGU4CHEdyy7P0Y
DHmwi5pS00Rdh++9HoYVJO03+Y5Z0q1zwcQCMRrclJ8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23104)
AVgimmqksEnfkbdg8rLpXKsIXFvzSx4ua7kAaaMtaoT2DwsbUgIGF2hifMjU3tT2
VaBIkEYVP1EioEMOA0ZopTygLZf90goqPIzSXlbO7xuhC52Rwy+X7djHhvpz5fg/
1qqfmjERy7NghI+NlVgSYxI+eNFD3JwxJBfdTzt6cFPbGKHDEHcXhtNxvoHOT81e
vxgPFyXLuhQe4gZxS07c6z8paGb24Vxt0cnMaTr4dzyRD1UpxFX7LTanjF7fFq0j
1H9MJG11kTqsBcBBfda3Yd8RvTv081v2IyGywkVy94pw6tNc1dJjrrK1jHjNrjGD
dG+irb5cUQQsINCbzGZCO50XTxyQ4iwijDWY72GKpABb13rC32fG1dOIVO6ggBph
/Wc8NfHkmIX8+bzeqoV/929+eZ7OVTjV+vODLUMgePXrOWn6CSumXXBBSBkdg0jC
/9xBlGkqsirUQHTOn+QDF6k2SYS82R/NKYQfAsDdkhJM/CmrWNSMhAZpWTKgMInF
E/hnHdXvrzM4YGjZyv/P8isJAQcmrbER7YYqLgMYRN5PFVFXgWg8fHrLr+h77qkp
lyzzpfBqXrCUN95bsk17ejpk7T8mKW33U1pi5tIRx06Zn6EzsrYPd8V5lIZWkuZf
5iyaON7IcuctsFo/knL9We3hTnwUmSkC8HjAE5Sj5SFTm25MXLKNcLtja3dOv+3J
5G7dgHEHu/BY0hN1eDpcnWvAK3pV/rBZiPuz5JKrcDVM5EQYn5t0r2cM7bVCefd1
XG3o4SExMyrgDAdyXE9Q2yb+LJh02McGBlP7m1uGefjVCr4gCVlzcL6ZZlM5CRLV
P9PeiYPWWDBFI3/+nR4/BzcOoxvXPWmoHejQS0ZHCpLjQIxFWwmuA3GimxTswWB8
0vMlmCjHLi1NhzjbHIOTwCKPS2H3fBhEBEuDAxSx1W4zLEzp9zAiseKRzBNi53vj
XGa31PlaJHEQ0Xkr+ICKd3YzrK27UOgYIeXCDDCv9WIoqYC3NetjmJkHnrP/wYxE
PJTi0rWVvDikQfOQK3JvRIBTkTnguw6lTPdyJYCzHzijTjruN9jeoBIYYksUxPXV
B2YYvKahGvxn53lr5hCoa77eHDAwQ+M2DpiYvTvFDQOZ4vx7kRQIuQcACIzlFw2f
xRrII08ovKUJ/b4FlpYl/jeXoRAI0RJz5y0fh9Jl6+fqnVmMhZhwan41Sk/CT3LP
Vmsp8vbX4+Ck4eKbQP3vETK5vyfGIbfKDFC4AsIIKcUW7hYVdlysOQbym0eoKbCY
NC8m7iHCfBT9+z4Ij98HGNIYomRylxCfJ8O35hAXZxmXEX4poMkp6/EZzS6OzG8e
L+1FxJHSiWwlbIjQDpVBWAiUsXsh0pz6KtWBvVkHhxBESn29vet/J1/xg6DL/t12
9f6SIajSB94hvuO/tnVGkK8kbMqeS7Ogt5vALd4gmapjm66WkpXZn7WDTFVIL2FJ
hTBehYY7BaAqvvn+r9E654QL6ZE1eG316OUciK4B+xXArhKWvomybcxuFt59rvwv
KwbCQFrNvVUzkfdovGQ/nuPFM8EeRzzKPX5+Pe/6qfpH03+IDWMb66qGGzd1pcRL
sDsKbsG3+I6U7JOysZjkIhL7hWYm7uiEJ7wN5YRYoBUyTfdtnC7tO3i+SogrmmuW
+EjxF1nfIDXloOXuuRCSzlKxEdfY3zJ2XV+uhPL9rCZqf0GQj88BiMTCCjuBY50f
5iELJn9VkX7ZSWKaaRSHw3TKI6mqiNNKxQRgDX+8l2sMq62o5KTmnbSVspVU5tKs
4dg5MWxtvA+ZTLSSH9ojn4ExvDmmiKkozpIXKiO7dWq/l7B2I7DntFBy15ZRqO+P
xLrFUsplATXqZvasOpydbWzCnamSHQVd0t2USiARcgKnDqTL7lolX6CjJWWkq3wI
3b8guN9m2ExTChqmBvkSsHl6RxIg6XuIkrMYL3kCnVv1J0tmrr8lJD4oPbT7o3W7
TfnvAsMAB78X9//5ZLkyN6Ygde/RkvRJow2/BljYeDqjO22ljAmsc56rKZnb8UGw
9NRXyMjNR00Yql1qpwThHTW3D6q3Wgx9btOGqU/0tyOiAKZNbdFDb/ouisdkXqbE
dK26u3koiTAZEuVjAvVc4WOLw96FhX9P8x59eAUp9BRpHvK35CqHmpo6Zp8eaiVP
xwHpZ1laIC95hqZNCZdJ34QgXI3JOSiAcuEvYw5K9/NYrf4Rm1VYMlNpK5GUdi95
FctDaswItCqnXIuyJAr40drIs4knsOj9Ls+1dzUPX5qjqUwyofvXwN/Ghraaes8r
CIovqIscdu5JH1aws4Ga2VhYgHHWxfDpZ+OnK0XBuZc0BE4216l/uBMr3zhCPQrQ
M4GvFufltLTEl/icVPtJwTHzSgHt/tvyOgKM4jZ4dDv1NBFKoFXGgDIkmH+MARX/
PB3S4LTOO2C3DFIGkO+ODFzaKFvqbF6TfV49di72BDwfD5ivB656JynHmVsUfAed
4q81V4jn/BNKdcTokdL8SBL5+nEmS6Ilia1dCTro/fBtkhwtpX5RseV5fzS7vZPO
4SwGKoE3HwZvChwiXAQihBelzGzm643I61iX3Ys84TUOZqOo8qzWLMT2enqtU+MF
0xsyo6iYg2n9mTSAVVXMPvNOG0twCRWbdnhBsLPjmHpeLRfbuyzoSr4AKsIwzJaS
+593g5vdqL+T/H9BBWUh0V56+03R7leVKNWkCa7pLi6tnV+fcBXLs9IFFBQumEJd
BVL124vfr+wsaZ8vsdrrrEu+ltcJcUBw40V8uUOivkyhfsFWlCe4ecEuag65DOwq
R2N1VN/aTfBKWC5spNtebkcDlOOGxH16uHZi2EEG/itUus5HenV8PlDtozgxWwvN
JowmAKpcrDQ28aIywMTZMGlUb1X+xuCImr0FENi/xV4ni3CB02zd7Q8P3qbMe9a1
PISv4dxuVkCFR08HDpUAGeYg3NplOhuqFnlY2NuKaKS8OFGDe+tdJFGVxgzstLDn
KJY+FNdbDdQ6lDhjVYXWHm+if6Rayo9wXgtYGU5KoxwXto50X3mh7Rejm6l6Jm0A
5yiTBirNbXhzWyRVNh/8YDvnVqMJJncV0V5rELIIK0zup85X+4k8kt2LrChzSz+u
agyfKX3X7ADY53WAV/01en9pQZtjBm7pKqzKrDStvYocEqMv15RnTE+P9LWJ2c4z
LLZBuItkS1dX3eMd7HCmnOhYgg5KCY79zvAjtwX1ncL6Z+ukejxI9gwvf93uP8c8
7Ew0EqpZKH1QkaJr0URE2v/yiMtN6pAH5vVDMbrClRF4qoYNkhXmKwRcJgH/1zdn
Z1g10nH3Eoto6fD9ZW+G/WmxS2xGVU/+JMelPehHV84HWEw+HtH/vja7NZ5M78oJ
gaaiy9jwl761tDlv6XaD7YEq4craUBmd0b2rGY1mLqJ1Ei3nni3leZh9ODxrAY4N
wH+s55qLxu1Y3+2vcP8451l9m/yHp/ltSj+riUFVgMSgXtHgoqpZNPwgI2GOX6aN
kN0BD3zSEr+eHhT4ekDxbt+++BLovOdWGy9208/BC6YoNsqyTtR+Aa9N1a240R9n
qIf+HAO5p2xu0sWciLzBiIqZR5T67+jYQm34jmHDt4pG1ZBH2pLbKDdGnqtbfStP
S8AA3wW8plrZmYPxrRRA/UQFNQuUu90qxCiMcfQpPVPRVaNlfYszihAkTp8OWNqY
PVAx6hX9AeI4qdFupkL4vWfW5CipF/1RQMDobymXcwMgHE6UEgbmA+1dodikBzg6
Cn5sDpr65vWQ4Xh4r9c3be/dM1g5yyjy6N1gJ/PtG8B6lrf+M1LhUGTqgm7UJ013
/rVOCe0MrJ6rndOrFrU3JguQq44w1bWvNDDg1S7pJbCCmqkC4NDs576GfN2lWjx5
GtVyvzcaHoXV8Oz5nwdH98GgMnatNGq0SNh1xq5sjYE/Qy9RoDkM24i+QpC8K1sN
YfmX8c/pkz9gjvFlGByAqPVmJ9F/Q+8oMrPfxwJJXJS4Y1uCGRodcpWTCGWa0V6b
xM659s3jdIEZebOwK4A9bRko6OerOx63Lg0KZoUVWwZKgCTDAk1UkVIDiLF4YVYo
k/rCQC3xHTrd4KRHxU/6agNE73diVTX4m/4ENlqWKrM8FNgat3NyEMiDoMqBFMOe
dQdvKMoqK4ED2zLwUL1K6U7NGNc1eWIRoBgANH9GApusLzeL3cNsP2WR2kD6K+AP
dTYJ4uMS4dYFlbIge01BWulA5/2TNrirveFnTigPAhFieAgPnxRI9DEl04H0bhmA
dy8vfHbLO4vD+seKrdm5i+hY+GVYo5R5tti3FsSe+1ROjJSueiif+gNWjXFqV9OF
3bucud/IUn4C0KXxWjKjOXFpEJpWVbYZ1gV88qLKCkhvJxrL162BbX5NObkD0hcP
mGpTaisVOk6KGL55t4fz9aQ5+iUgQmQfSc2Aq2zLdHXdbeyB42VsMXifb/CT6QJ3
yw6yaLbhzEpD228wKOBTTKNT7Ae02N5rrHrGiJtORpSeEdQTO3QmI13UUL/hM6el
iwWmezWdjzhx3K4CjR1MfHPMp/kH/rxqu+wUriXcfU1I/86hF8QRihOsMRJ23ulO
Vcc+6QkvvCmCIL85KHLqvv+tR+DnQvYX1ePc8Hsqztp38xoeWJQAzu1HTH86zj1T
PGOIFpQsT53iCajv/SvRXG70/r59pFRM20w/jRI5Pjx8BExFxa5flFecxcI7LPB6
TDLMf9Et9C8QivuHSfPbiNhdzkFto5psOqM186rpEGLeZNZ//lJK9uuGPfdn3/fs
0DnEgEgISgVLNDdJ/Kn0jLHypbgBWAzWE+17ET+f7CpNNP1ThJ1CWkIHJvQvLmgi
8TZC3wCDShHYhZ/d3MQWgkZoqgOM3cLh2EzkUC0BT5oaCvbA+R3bdiTNXWw1z7ot
LwtGKnkoZ5C7IRVvJSj/l7MR5xFEjMdEyg2ZNqMxuEe9Zk2te5Gph34Eoi8UDHDx
dXYIRenVtmHoLJbsqVg5eEy7tRBPSCY3FayVlFW8VIA9f94oK0iWt87If7+K8LY2
3g+HJ1BcDBMMC1AfG7qA6jQa1ylStT6T2qAATJS342gVlzxrIoSMIK0uStGqnJGi
0F8QGq7iUeMbuhK6pDzUS/fk74ykRK64ag6ateAteJ7Cazf75xpGn2hTmbwtcJCu
5Lh3IE4ejZWmq1j1riPDGiC97KgveRGUg20jVktLDYqNNgx7QvhHA1uFH92DkziG
O8cKy+IUiRrZFrVMrl7TBUQD1DplJrOR+Pi+DY/2janBsx3ny0bhfWtkGrGAi5tr
WqSisBW0dO1JCcQeBSkujo4makPhbS6TB5qVwDS0Ng9vnt0bVOXWvFThWaMIvFq1
HQSHeNQcfBd43RLhcs9EOwG90fjFDyCYNieLFNkteiYX6jyQv1knygBaAFiKRa4c
cUiU0DCkdvFnwsKBDy7hppj/WrEi75VvFc9Xpz5IaN9n8EWmucwYc4FBtpzBFsZO
cIj4FN77pHPo5XldVNj/uGMcQZEWZrJCggPqRPXQFCTAvsftLvN1dV+fLJsscHqV
+I6yBHiwbZrkBBl4qzAevztyNeQvR+rjL2VwjCr2HwH1ZV6Ig0+Cm2NCaA0Q8Q0Z
XybwPHG9pjytPRFMEbwvkTq8oXIYsHbscvuN5J/U/G9kWA0o7oHfPiJC5fURhvhD
WnDIw20U66+OEjroR0syRHTMlGoEEuCeaRJrPctVsQXa8zSZ3GDiK+stN8vyFRh1
KNA2lC+zvr7Lr3pN2xiwa0YnTMtiRltlZXMscBn/+Fw8rAlNj8O4dzfGdNmNZTwD
NSqPxuH+6vXCSdc0zhhPj2ldtVBek5/BW8t6JLVOu250rAyulqooM+7Lv9LCQb2v
JnFhXTfASBZ3kvqsmeHSQe/VcD0G1ByqgNWNW2kf8KbURe8rx4L/LhT6E3G4oO3q
t7yvyFZ5M5+WPsDE2uDrQFvn2tfOjzR3kT0rssWiVDPuxoDXxSdqayc9BTxPqFgK
MEafl0KAsIEtPdLWlXKF+iH4IetZGJNCamz269oBvOWqhVlhNCQTSfyO0p7zD25x
J8gIusQleeGFy98AvlZL8NoCDbDN1kgkAx0Mey4qipvqsw7L20Q+AGfR0tqDIunI
id7nnDNwEvWhBdnPl98t4CJLYyMyM5s/q6pgm3ZDuxk9NFDmtv8d3oBrDawmcvWA
rqZm+syQDn3EC+HnDu7H6dEni/3vduaD2YTYQi+jmu9Dt79eEFSk0f4ZTttitQ6y
9xjUPF1OCdIC3SXkHtUcphZCUCbnWCc/cCck6nXn6gnOmGoCJPpAVW/zaFfqdt6p
ifvZI0SEvowUfEwhucAXGEZl7E4ph2Qy1K9vN6+XgMt+ZbEcflsjsfG74Us1MehM
50klG0AfIqn4bt2EhdZkJyq/uVrc/JWq2qc1orOWIPtYFH2xZKpOJpjhomkWcwSW
Mzl3KWCLIur8U4Cb/uZfqg4DhdIU+zRo/Dfgy8f+yrrVU3k8QHTX25LbFsuacchJ
z/C7WB+FFK/OKkrguTIXQ17VurRUakGxcQ88Z8hSlgWMLUp30TZSMk5cCz11/732
SUmtiuMTHexJhVtY7mzivyHhWM84YGnBByoPEqhev3FzxudX0tFP5omoO6t7d+b0
Zw11+FcEYl2d/0WjYQKNTpKpUm862S/qo5VtR6pAMy6VmDN+xLI+54M3OsEmbAP3
88tKjAD5XF7dC7pixRJhK9bPiKdpwD4AwnnDl/UX7WhtRLt6klviTjxVwitqwKUp
igos2ZuNEnWaagQK0NKLh4YgDy+a+00kYslGmXlX99wl4+ofC9cWZd6DpCLzTPwN
7Z1Y5wJBONCHZUiv7ylaLP93gp4q55wZiI3ORH4nhQYYZKgclS3iJZK1TImu+F+O
9mwSDltKqPsQYfiyOgNSXB2j6Kx8AE+9oB7VFz8kxPgEjFhQ1DXoFLuSLpkoA0bk
CBVnok3TWEeq1VMACo7yyq8hlVfhfuu6BPK2vTOPWsvFpqyMHFHdN1z3bj+cj04E
1uRV7KX0x96q9OFx67ZFjPoXcrLqNkXVHCS2NF2isMSUjTcrB69QMin8ayGjoCAV
xj4sQ7jKRdWLFiUh4yDd5vTQ15qIhUhjO9+FnGtdut2J8YCFvuSbUGxaYI9YW0f4
f4ZrSBHUCHwmzUP6MO3M8vzQ/KyTcEv4dgH6aFtn1F9HCWLnn28118tW8AwReyiY
4YcZPWosXuqt2C4aTPvtAaleAHzPvM/UPhj34dJ7g722wwE6MOs2ha8ElOhFSKWo
Tyx8ERj0pkyKYWT6ds8yD+lNYM5NIrmT0HsmDFkUC+0ueqcSy9NhuODahKLmBr/O
XH+0+KddMOgcbj4fh66qxgTVdBBOxNCsEPk8UuqTeKcbNYVymyB0EY0wZ0VuTLli
+m7OdH/nFz2uLPc7Vmjfa6Iy7sZVvjV9xXhmHVmJw9gfF01VHOt04PYre8S+RDTU
dTBH+XgdSBee9y26EZl7t1T4VUcks80LGNjoAdUJ1jH3oVm5t90x1/8N2qQC8VeA
NQeN8cd+wRIUu+UaJunoG3aUAwmT3wJeBPH/3+JbKT0X88L7fMZvUOx5ra4l9zyi
SHPjZtVfAvDFj4K+83nBjosmklZH2n53shtVUOoluvsSrC3b+KPhtC9NYsKDwgMf
IsrhLrw7boFSVS+OvNW3BUzqLad3gnolG4dBTqXubnbblx9fftO98eB5yF/CmJVo
t1LVljYJH2ougiEbDqhnRAWiYMpZHe8qwh56e+EeQpScv7Moh/OoEumpgsS2ZA9q
OkCAtWPGGIzQCNa9wQ25eACw0kUsQdjTAU52OS4zl5S1NFJBqSaw9T5zbXYqX4rs
uLowcHOQTUR/wuzlMgl0cKKLX/gH35ZUgS0TxX4iD2YgxQ9xQyNuwTgv2j3kaFjx
ZrVFOT0qUo5nFXqhYrVMRoyXv8U0b82w7ylESudFOcTL4tHoTn1PtDiLw4deQBYS
f3WzbxmAEcKrV8ANn8Hj1pAs4aaZsAUJhAmHd3pcMpb9rAMIOfxtXFrGXsTIzyOQ
zKBCHqu+mnD50/9+pCIWrPpbretkQQPkj4+r96A/yWhhoRu+YowOaFD2byMslkYe
9n3GmvP8ymQt+AW70/uDARXIZB+IyqWzXXfJlnAGreDtVWjmhoqnW99swjvIp3mt
hBQ5r96noV7MWxuK4EeSrUzXFsqh3J+bzwT5HNuHaxR+qMIORWceQfJ3OiAaGX32
5bInTMZ/RsDkbjaG/E+rLHmO42+sGup1ANBu5oz28PdmRX/bkgRmUwi8xIWm+56R
BkODsEaSxH4lR8bhIQtSaBKtf9aVZcLTdH1EMpPiNR6uEL87QIeOiqNRwdZ1NKzP
uyXioUtdHhffxGIsyXfV+YGfAuxNzQ3G0yP2gwavLVHelrQQVXFi40CiZwo9lf1r
vpHIb77lmIKEaCI7Bq/yftsEzComqnBBKMy+ifR1qCrPJOMDqeUAajAlMCinqfq5
bdW/gaxtfqHvwrFFU686MpfQJyzvdQmPKIiPHpO5bk8n8MiCz2/+1skd9XPxDRwY
OqsTy+tADrOrlgKRa6lFk1ezB+JWT066bcQtkazza77+CrDc6izqrCdA1ZZF6XS6
Cfc9XePz6IHek5zqmYiXdlPyQCFRtkDn7niQvmC/xb3YqkReB1endtS2AbNWeqrz
UfzYigneb3202Sq6QGw6DiSNMFPiufgxaUabxbUWoJljuhcJySDooSVIR7C4r0d7
kTuiFACIAYRisZK4qM7x16qUW4Nrnovpe1+43DDWShtq5+cl7CleephJ5Jt4GQnQ
G3R0+jwKDTI299vjX0msKAMWDKFaXUEd5R6t0ZeLkVk6lr3frvbZEsWgqlTeQWF5
D5v8F2p7WFkZ0F4INE/VGoz7Jv6LTUtWHnnFt2IkKGI5oni6TGS/0mRv6d3Wo3MS
/sMIebGIHfQAC2PEpu18xC095EzpDJwMgdC/WLzPM6l3WHi2dWQmejlL/jFdyX8c
ObcM6kOqEKsFsfIPxJ8ZsSX5qdOv36iO2DEkcP3+5djbishM6Kq+7QpRYDpBXSdD
0QxHMw81zSaxT7lhUbu5sPecQMxkkgrWzyo8s7oKsXm6cyguhrDuJ66SoSBoYrHp
dPpS1DlIWWKwMSiWNHU2Tb0Pi4JHwajfSUqCkUrN2qSqPtoKvCnbP2C6sZHJemPZ
3d7oNKcnUgRngtCcZvcuwPaxP0V2WPaZRAPmerPtIPdRH8mgXCkXwhGPnjMU774s
FuyPaHTo/WQNu1H5BvVZ41S7PanbPteZ/dpqqbPROnZ4chgIWtJhodD5f+zwKfmc
2QruUjgTimlaToCI18+r0Sjgq75AR2sQoikOmOOngSSRJQwjAbVX4CTkREKZbN/g
mFmoo6s4RsKftBbF7aEmT25hrM52ThLlkn/7aWy28wy+DDIU6kgqOKWT5SLZDe53
2dD+KnVQ1VYOsVUZ78XbkBb/KuleYFdv+9+pE6z42KrIpngJFNAyavBAxAI27Ult
3M/Xe2cPFdNVeBjifwQTHLzOvh9MDdXV/kzU91x22buRGg1UnQkWuaNoaEW2Rtag
9dG22KoACNFz1A/lhJ/lH1vQmVLkPop+GkLTVo5RS1ugF6UChsUriq+coV3T3dLr
NgZGB7dAoVS/+/Sb2XCD8DmrpBY4bDK0FokoB0o/rp0ER96BSDQp1jAmnTvs4LYP
uFCuMDlXBoPAiKo81Bs9W8lAocurhSrxMHhhvmtEndmgLWBbHi8dNurBlQbtPzbt
4UxE0DjrcIfLRsflJVApVdF2DXVIRpGTgSPyItWvsWMsQHGzDx970pyDC891eWiy
FqQA7un5dkg7OVmp0nOJmF6Uf43B19BCqXSVzWixvIfkfe1ZR7LtdgRX+r4Wf2ot
vyHKf/tEKTpI2SOT8Bi8kia9MMUZZsA92IZkcg3jKDZKCovdUzzgjYcvu9XOBe7T
dJd9mohwQIaDATCU8qEg9RyK0LeD/gjVCEnzIvxi+dFind0c42urPWa/Nb6vAQSt
4DmYq9v0IP5DasXzhy93FipAlPqWODZQ19OzZ9NPQixgUMl4e8L2FQuVJXGDzz+V
3CPOW3S5tQEyTvqexPp3l9438kBNfXFYdpicmKMUuIeNLpMkduB6MgyVuLTVwLBk
eg1umulQea14yeDgEDQWQYVtAVe+K5enA6N6G5739yhUy1JkNnmtWoekEFe7C3cs
OiX5rclUEe2rbyQ+N/vPsoqwI66kLfOX34tAD3IQF8kQarWx8BFmRC7tdpCAmfIz
q6U6H3dKFrXB0EZU/N18u836dgXSSDgGpbh4XnKXdD/Rj6/wQrM/wjHa7gjZtpeM
z/y2MLkcHPJvzy/5S+0D4gyws6fsD+Pj7qfENmdYbKgLj+pIa2DXpYM6TCeM/uw+
MSxfn73I1Kphcr6CB9ILVGjEHllXFWA8kf86WfC5zPI/XHy/UQKLZ9DmdEtOiFrf
2J0Xi5f4PjljxbWPh8+hwGcEvtV3p6p1CR7HFK7ARuPx4OI57UY2pxlxwinrNy6M
CtpwRqetUfMBKtOLQ9ka0TPSx3BPs37Ofi55u0CODBgULizDdFWXDdHqIA9nLJK2
rMuDpEvNk1sbk4u0+Si2hqwxJealuLrA3+P7m0nD13t8QtYoW3+sdYcNGlgwFqjl
eZGTTfvYEsepqrACcJ5NB2234mV/tN7kW5IY7V6g7mwzNGrd8i5RvR+77GjrRCSZ
o3O06u/XRJkMM201807M/e9a1z18VWIWOFBRRKbwHTZZECXLgx4z9wI/G5jui+hl
0DIrgc4XpK97DnTQurkTbfpCXKlWCdbujy3h+VsheRhI0DshCyh47hpQpOkgf6Ks
QzfWNSiOzlPwNTPtLvCcTdhVN/69ebuzpNWxCYmyO4s5utUCunDJN/Fe4u/9pN6Y
owOCGXxQ01rmpTo/BHAilUy90PWEG8iN7ltkIhQec8ed8dcXn8uPZ29byJkeIoUK
k685rmkCwh4QltQ2Q60yNB7UBTxsWGHRDX87EOI/y899F20Iwi+wGrjHu6CcpT9s
FEJrxLEriS+Pd43WpFkerEyK8cVbM/Au182CFQlN24+KUo3XkCQaWvtbodiESDwy
71Eb7gMuuXHwPMV1LNU4t43/aojzTGCso5wsxw3GzSsqwlG4RURq/D9jW1bc8a02
JWMke92uTJd7X7JZC/JQrrhivcQD1Ckx30WYFLcGn5fw8VZQ29Itjt8g10pA6j8V
E32n4EPOSzoC1UE+lmjpitWLI0DJBjwM9jBQE0Cjpavu+JsVNJ+627cGb731JXs+
DPu/2Xt/utVNNeOlUk4oJwiaMbVIlVTBB9LKa4kzn8V3QuuktFFxivyjxumtZmMY
i+s6+uiCMpjyLx0CxxFXV9jvKq+LhfCX2HoPiZCQv4H+ZF2h45UPJfEnJE8YsJVS
vxogCCbfmC6ITikNRO3qflqFxtjS1pAGDFFePPWVa3SeTh0JePMVgzLYmSZAq2rI
ZY7a1MzdGwyzdJB3tCzMrupMx2ldCz1JURx6DHnjE4/VXbC54cfU99FX4gPlSnoI
TxoXT6+7D3qLjf2cuzLXaKMCUioAoorXk6aTH1WCdWJknwMxUYdZpmvXUSKMwgpV
d+yjAEmp7yL3MMswjwF5WmClVprNVbI/CxR8fRxP/RvFWCZFgluJIihT5hp4xfsO
cCpTYqBe/z/GiKr4etOVCdBWH0mC+r5e5rW3mvGj5omJH4rSb/Z/6H5tWszVUlGk
ycC+r50uMXz+MQBNZxl+ky6k9Zk8l2xA21LDJEetxV4P8eI5Ybokyu60FlNyak07
RDLGmStf7UnmSfJ6YC7TMMPU7koNCi2VC+lfTUPACkSWXgAltUULXB7a5OoR6Dg3
8crX+Xv1ILeHFyUpVb4hWF8bhfONcMkPt8t81r1uBLnfd2WERGZS3dmJNg+Rvzhb
B1iWA+yXR2dzrQCKPYPrwvkkpnqN/HW56LEfu5JS+MvP/AhWyBS5SRaQlghyEK+8
mrEfBWg+CrR2+XNWWXup49oJDnsqwVXTXiP39Xt7/4Kbw8ZONBvX5Gm7JTQ17g8G
WboIODmUyiLet2AyjZdRgIL6ddP+p3PDfFQO7YtYYct8cMouCx84pKHRec0/cffu
nEyxWPmaFT/Mmv7Mowlo3yMvl6wG2jZCIH5tXS5y935h2Z/MyYOB+0ZQOXFFK+GN
LE9C4APMbF2mEn7Mg/mKAu4vX3sadOZkt6amiaJvEdN5OHKpVFenpSusX/YaeGJa
3WeHJOlU+LW2e/0lQooV4KWzWiWRy7BcB1D3xWeIdQclIRTl9gFdHSt5LE7WxCBX
xxgSdgPD736OYoM16XWODflvQFTy5T2GJwK35PW5U3RBygjkwzTjcWkU3i+QuEz7
ALVn3MrrQYVjb0Z+mUXmyRazo5Ejq6EuJLgB5t1DedrJg6/Su00dv/5loPV3iCl/
2ATHoGIBWHYvRuxlbfZUyvgSEsLwDaZAGwm4z/74URjFoV4znmnrsEmPgWPO+YiI
xUwrWhMSYMGVgbcftyh/T5Fy1oC6rsVMucRaME558cGq9395JiBN3HSD6TpsP+qY
oDk/ck6d3eHRUL3/8nBbrLWCC4WkWwXrVbIpnJsjgNTAK/ZAug4MeFnOZfg6eq0/
Qfl3cEWhleqFF1ZcBwqVpLESQ5ol9hTG5ugknDIlcmisNBv+qt0pAwdeMBS5QZEz
oey529zjUYYXiwRIoY3FBgwYGECf9a9KG7J6YnHOrszlmSjiByaXa3kikVfa+2lU
+/BmgwUjfE/FPc5bcTF2kfcTC5AmLrOGksHC91PypBqXNVQmJTNyyYml7GASCGHC
5Ey5Mg3Or2T/TBFH8F9+Du816nVfrr/pK71XBeZfFnyD9jLYPT7tGaAA4K6ZcZE/
2/2mK21y7H3VKhVn7N7PTXOYGX11hHWCJcJ5o8R9gVW7vPOMetTsHALB3bP7KIKy
EyWpIZ2bUBnuepgdO34HNII91KwxtcStuXxn7qxLfltu2nPMtEAVSPTQTYLOis+x
nzs3/8DUhLX9KDAMLm/82KJMpluDTraL3g4aszOAKGH5F2VE/KR9NsCgtx/ICS6x
0tLerDfKYpFEpUBIcNuLmQlbiQvpAQKkINCZa2suR5C8MhdN/M8q866vt/VaIsMq
qWdGukhsQjrayDJYXL/FjRY466NZwAF6sUTfd8aW9nDI/RogpgrYPj8TPQPhpNCc
FBVv02C4ny7fE5mVPKWJctN+rPCCsS7hlL7/0eKTympmUswT397El03Rb0vxrR5a
Plahu4y9z4PvYsyxkSUlbrzRVp/U+thLk5tgwilqxIf/kuNR/20p9bLNpG1NVTg2
IesHQUGd9AGc4faehJEMaiXkuGN+W78EG+N8mg0f2PLjSLPRblKWG4cCx87YJeRu
j2As0GCcJGqalP5vzXFlmqcI3x9v2fbi19m1DjVnWOlCUtcxDZWL9Q1SdSGJElJK
0xQm0A9+Z12Wa/s25fCiemlkv9qcQqr1uBHAwA4hQNHVk1UCJF3IA/BFOnpz2qgg
rKz4XA/gAYmaV9EgHGYftR4ppSlZoLSm9tUyoHOAcSgSWuN+dla/Cfj9HB7UkO4v
DeKdUGoQLkuJ0XqzZQpJ9jl9jlcLryi7yxQNoqx8RrXQStJ3mA6hcKatt28Dy+4f
Y3sC46POFKC3yP1PdT5AjH+R+M3Y2PaVA8VTcWrc2Av2NktdPGx1SyMsTdBTdA7W
K3Xmi7WPYlKVzESUEgyYuoA+bLDywrG6tiJgQUmlfJimj2GQkeBj0cCSXx01PMPA
GKRElkhVKAZReF6gU4uVZuijD85U9KgrBlxOGWXb4DNwo7zfs1Tj3HXff6YZ+qqy
PnYL/zdv6GEshgNspQXR2KuDIPq1lYAxm+7b5uPupKri/AyGOX6v/XAdOKUJuCTI
exNLGaJwQQOIt9+PT5nzbvyDetsqT8TDiv8t7b/LukrIwdhWKoRqLMwtBd28eNgH
+839xXayNhCRFOFE1EC13H5qpmi1ahrLXauLB5hP1CbqXFQMpVClkE+zA7WLdiZ8
CRhdGlVV9GN2p1qkFY6KL6hAIIGKJOIP4cIcZ53a/fLJraMofORamr9+0QhW0kVc
BaNjBFpgbPmMsKm+5tb60M3za0iMOKagXQgLG1Ca2yDOT5nnvxGLQYp5JFy7CK8R
PDLCLRpht8CfltY2dmWlJh9PmzX8RHxYbXXvAz3mibBFBo54ffqrLpJnn6z9LDv7
AI0szyPwtOUBglwX14nsxeJ1cgpP5rRhG+I5PD0LERcxs8i3ST6jlEyRSt4ZB9RB
aUKrBT+WMA3x8MLRZdxD8nP5x7dL3WMiPLnQhxWxmhtzjB4YKEds0+iJNP3ohlNK
ZIksToB4wRQy9Uzl2W7xZy0tHO72NkQ/foOaeDMyO6ENoGDENUQ8PPJmG+rKnu5o
McAbbIEsyY18Ij6ttk8dpMF+E0GQCflFMhlZcBfemYBb2NtTkHVSZag74US5T4s8
a+iENoyDw+E+G+2OMgOfjFaihQudvVhGzCrkdx+qalcdGvND/ReQc9so9CT5ouf7
60/mNXmujbdFpy1Gwj8O47jJDQ03uhrX4DS99pmTJVHxVZ8u5K0gt1nEEPgXrW3e
5LvifHUa7/JiEiZ1OOLrDakcgu+ODXnCxPviNIFtfMUM/aNFZwlmBXyk+S98YE4s
PSjNcnPqCmWmjfJYL3Nkwd8cQUj9yemTpJ5VgGDbr0aXVMSqe90recqPMx5vog1Y
7097FAFo+UeOkh5OcC4FbHHoyzufKkm+Azl1l7q7yA8HFP6pSqXhS6vfde3sykWL
pdMVgaPwQ+x5I3JQa4ZJpJe1L9cqQGOZU/CJqE65qdfnOloVzcrNTmYi8V4Be6ty
6eTl/Ljg/HnG8SlZkygNcPslYytiwaND01odKi4xBWlzs/ZGpv4GL7l12ZQH+iAS
AmeWP5anvTEOVLcdL7aUgz7jvfWY32PMe9kSehiwvdOP9IRHaZPzTjwyxTBcszpu
x69QbLf1FGkIbpU351ilFs9icLhtd8CcX8gODun/Rd7BM9Pj4bLNaixwxeH38EXO
48EI2rUY/2y4i2efUStPgBdf3abkLPXBpEOZkDZpzCEcf7Qqdsfs9Wc3WiBYnVQO
2x9DthiQPJ2v3u1zQ7yzC++0cvKtTTcFwLl16OmmFc+qH/quIRUYOuhaoGvkwxjx
Eg1qsj5w1JHivNBcwoxnBhl62As8YAbgOhVb8LjNTzu7FNWmJG40P2NVW82M8hZ2
kFfWVDHLel1Z/gI94JfqNrv1c9ixUJlzA1xqUWr03WGnFwUcprbV44RMV+vZN6q1
GL8Qt6LWFem5hxedMUXNSXdw+zHl3de3Xqy8OEiS6f4NH6Ip8M/rTwMP9afrc2os
RjKlADV32/1OVje6DGb+edEqwuWuoB9qrEGzlxNrqBGq3BBDjpcqq7IZuKahNvPN
Rj+RH0ebxRAEjx1O2Vcl2qk0BPRb/4jRQD8dWoTwba6GTwN1c/i6h5DCKi4VRtUy
5VhWETkXtK3ozPfR+mgkMN46G35ZrJ+ldPfmajgyBTxIyCvs74cfskVWiLtsAi4X
Stnjp0N8lP5utYu3D0E4YAEyyNOKn1/V2yCdXkqmwNuVgCUvF7Fh7cM+cHkI9DIy
nTkYo5D/mgpga4Jn/yuLt8wuGC+iE55n9DfbFwOtREFwPMiJQKryDiOyhsdunBFf
p5S4jqAMYWmFMbDqeB131w/wmUE2FThjYiVP66LY4OY2KkQeM8tOo0owR6lMp2DG
jyOmFrHQ8VxD22AGXqkanTu9m1yPXaizJQfRfhupaVrQY4ow7xR5Ei0yFo5AwcYZ
XSN+PtEl00tAAJSqsF24AK/DR7A0TPYYJ/IqYLJ05NI6Gx+4JypWf0Vsv71kxEzX
ZdNQGPc16b4VYyNYjqd3Qs5wnyrQ+C1dbssPvMx/IFc2WncyI9KROALR8Vi+m15I
9/6imGQSYj76bWQITmUfvFJKRb9+mnmwRhBW7Oge5O1vqUf+9TK2+Xqi2yLKZZXf
senNz/lmoS/znoyGCU/56tJV7zIafb+Nbpk2sy2ubzk3m1TqUZb7WTOtPvTqLz5D
mMSx5NVEtrdeQ/HCTcGLBGbZ8oS2uMOCNJTGoSQGoBcinxYRTlfntWSLXLYvzQ7V
AcDwpYe5+t4NL4fol+EYxvqbvsmX5I6+FhfYNZHau1IJCZTcFbLhoKRu1p6dwhgx
1SdPmhgTy48x2Xb7+Ckw2+3qeFCCyYAdfQZTE+mOZnL181k0eJMbIoiBh6G6HPA2
bhgaCJxMW01urGroSWi3BoK6ZIQwFL9C2xYl2BLUJPLYtUZmXnHkvJ0CzdbZRBi8
2lODwHeJkcJkoV5f5Srpruc6duD6QSsMrppRx6AKL6Xkrmc7WmnUeQ+G1jmZg9MB
LKT1+89hx5bW3A5o3XtDKIvPtr8i9VHbjsrd1iKxHjJ8LuVfJDZd3f6bqhogm7vV
oL1HSQjEC+Hf48tZT/Zk/ha2zBBtdJ1hW3yqRlSa8+TCR0LBPG1YBeIDLDvi035N
SSEJ6rl3gxIW85dFNY/48oFEYKZOv/kvPAbw1YeeZwy5bUxRlllDo5Z6H9DOprCE
YcxbB8d4ctwWvOoOzMDh/Ksgb5+E4yJYhNWbYTRpjW+PtuTMUH+03HDh/0JooPB5
yjmdK08bih3WroDFGFnp/bGtpxhR6yJt9bKsiZCLzgBH9L6ZC7BTjhnrXpojG15U
sHm1f8f2efrpJl690A5QJsRu0WFAgmQdvbOUqNaWjF6Bmz4Zg/TvuRt5buIsGl3r
MiPsuU7mMPLPRDXeh86t7uTcTXWAbLhbH62ctwL2k+LMtInnD6XtPCmGivJPZdEl
9z7hjhfifp42Ij72WKaik04nt06ir5TMkXO+BuKzDMpvuAZm6IrzhtnQFDveTc60
zpXLp7vVTn0+rATK19klcLo+QXScmNyRgmxWv/bvZSawsvRNr4N/EZryVKixfdU4
9RGVXH2/2Xi9lJpONfP3ontgA1q447id7CrmOY7mwUDBuVCbtPtFfBY/OjUdeCEe
OVZr5uzDp2aB987f93G1+QyuWp8nGfQkFrwQQmMYbVokpyv0R5/9PrumpAKyyAbU
VFnqu/i+9dktFhAB3jTBJ/zBqLtQ05ZkxuIRxC3ii8MZ3trHfcsphm2hcZWeH9zV
30zwclDHKyyS+abc9F0hYrM1Q/CUl2bhCsCRxCXS2osCGt4bUomputqxYKGfTlt6
uNgBcExLiWiBb5Ves7wvhpoJ43eGDvwMrXHm+g71qBDKBLiQRY2q/eotn2yr0ZJE
1bxv08V8jGm7ytAlISFinLAVA3xZEowJ1632f4XhMaBr7IoV7PSStGHuhCWO+x9n
CYfFhzQSQbcAcHl1+TnGXgYAGvFI+cOGwHO2IGY0DOVZ3vaSOgS4XpRBMH5GTMDj
HRZBrP+3QA7nwYc7AQ5Muliz3/5tIz6Bj422/wz6+K1sroDiI73TYZTMbA4A0s4E
lCofwCb+CZJRuyy01Mr0pQK5nPjs22CUeV77O3B0LO8AEUiafaxfYrDt8LS3/M4u
zwxJGAM460zfK/YG0tVZ9buvcrPBHQwZzWmtEJfpBLUd/z3k27cF5sw4YDQnSMms
oxVl2isOBiOIrnM/AaxQWFZlzHjuR/HM26w2+A4wgLXhYzx+eoAvW9LtRwDdMTmC
BZavzynCy2UWNnRQR69uD2hPcpiJE5LMgQampv8neVW8WPSz1Cdvk3G7LXvkVK8F
U5Bge5xL4dPtZ11z8PlLgjDcUeV1U+l5o7xv703m0khpyGQxqDgpACX+lSJAYNFa
fbxxB3MuvcvE6a1qs0seTBohjycSggFKFJoW2akyArFIuCiOQ+n3AfoprMitKr5L
ulOvbM6wOFLc7ezHUYQ3LnRM1Jzw+2AlzG/yG7WO0NkgiADoT4yDR5nscbqdfvGp
iZAMhceIAD4ubI0rwisJ/yxgbbLMlDFQMeVkQ1aNrGqXcSfpNrpSzeFMmmGnFMA5
DjuewrvMaq0rHzfAJYv8hiMoZ6cIgP6vLmqA44cM+3kc0dVWkZlXGl9FnlNeoUml
kRdJNR44PVEakKfaCQ0+voP3RLjoc9hQVXX+BkuxsouZp0r0s0jw45WDqfJDpUSJ
wtfG0qikVQVrVmcFn4kv5X26X9dQaxq5DT0xred8nkydEoWrbzXn0zL59mevnyEt
BAIuzFFvRTmNOxuTDwixvWYGk80AwUNZOTLMM6xtAmiclMUi0JpfTBTi+z3/NEZ5
jSR2IuXuBdVjuz6ufyqaBmKIKWVeUXwLtW1QSqVx85rAEcKskSKKfUEDUCmW99vt
mxJVN9ZWmk3Aei0llgdfXxrBx7Ri6Kn8cAdMVWQ5vzExhlURAIL0AsjX3EgTkpGI
lHfON4lR5kk8kPY6igf9iL2KtUndrYUFBWZaJTtH3Ydk33RH+/syAzICiwD1wlIN
4wPVCAaAexvt7z1PBV3QKTVrY0PkMpPgnL27HgwfwVCrp46MGe56zvVMOGf+0bQu
EY+l/8BG+GjT+PVu+z+IXfe0AVHbh91QZx8KqzZ6Ij08ey3cyAAV5zp7YuDzcen4
K7zWGvU0pFcg0RLsMtnBUiNMDerQl8s+m1QcY9IRSGW5qf+eT2Z+siXhDRFt+sfw
VIIa/kFi661F4NW0d9Biq+Ram8AAGJ/fCuVUiemgH3BGBqsSLZrj7RG/AaxqzU+s
4NzOgvtj6K95mrzvHLqzoMuHoSC1vH1w7DeiFNevchHTp9AEjAGYldg6elgNqc2U
92nvmimw/tD3OaC8zhrYWe66g534DhZPkxbE4bEcVSxLGNJ0B5VMlovsFf/YPT9S
o2O8zSAOBqxipY4mt0d/dTgDK3IuScQEq1icR9oEe++CWDWaPjG3rp0USje6BcYL
9jG+R1wVKYgVGoxnx4LrtGgYnZImSJsxa8A99Zs60UNdkV5Zp3At1Ba00hkb6Fnq
Sk335k3V2sWGpCI8bI8ic9pHamG8V99cZ5bSuCIqwsw+YlF8Uyp211qmHhIl14yx
ol4xoqHbQFaBanB4b2IAvMi5D5IiByBNfk0rPmn250c5Lwx2wiCv1oNrWMBwBHOg
JQV9DHM4C/vCY+zl2teRyOg1FETHIWUpDThLIIg3/Lhnh58j+msPjja8jq6tPVrC
4gEBou/kbYRy0ZyGBIWDSl0/NCp9owppgAhZJob85slRR4gZLa/u3nHQhHoOkkX/
PW6AqphiHr0OvHGTBQe0geKJPk/3HI11WcIf1ENGpudKQfAV0pf9m99xhLfR2wMZ
xhmQ0oiUSfHqiYeMFixU63I+kKN3Wmh7ATeU2K/gKcuPxTiy/SLKeWs3uSmNKDCn
iTridSMdqN9Pc+/66KN8wm3I+w6OQyG874c+zNlHi6v7uIG+SV9nc+gVPokfctDq
oSN2690xv/d7oE7knBmqtDt1jxDrvu07COJCjsh6M4N2Hx+Dtz4SQovchEmqAWWc
dsVkWWI347NX/4WdupM3WgOf5D8+Amm4htQ8cveMW+rrnJZ4YD4jVfSUkRelFaTM
CWjx+A1tLxGoKKyEVewQhTFJYZapv6/5DDvAR4h313qyvWW2JzA9nf5eNwKxt/6n
xR2SRHvVHkn9Ga+xV4O1Kb79g5vc0hkW//ubLi8IKYbBb6XBymBnDndgsOhgZEvU
uiRnte8BPiSEs1kguqtx8NcjGO6nfNqyHbQCGKAf8oWgHwk87z4tveyCk2uJRrQL
NvDzj7Ddqk1x3d7czLe14WAiiwicDbPR1amCS2E1YkhwL9SaH+15SkUDNm6pNOCN
R+ZDJPn0E6EFNQx4I1i6EMXKHyumSKdeRQDQSwwZpWpHWmVKr8yQ5ALXgz9bHqhy
tIBlhO+fkQNEK8T0VIYOGk0ckCunK1FSNxuokuXrUzmbc7Vnz7LUwr/qNnlrewoh
VlwfmEQl3lBtDv32KfQpCN96jql82aWvRGHiHUfTWsxw70/YbDm8l0ii3HrfC77U
nO2OsDD5GD2Aa9JobBi9BHhGkne0tv9M9qYO8pjlqwqNpdIpfZjx7EGljEcmyLHX
kode5Pp6lHjZ+Y5zvGZBLyQecu+ovEjqphBmAi/QYUkE8ISWGLBZIsoYf0rkuYvl
0xTIBgRZjlysQzPM0L/JM4wmLQXMxIFu+79x7z9WoxJ1HhZgWXk6T7SbgQOREGEc
fpB98Cvo6LrMdUKFvWliXe0DNdIFhCA+sw1aHrnVlUflkytGUOURKZBxV2vpqrJN
UAyuaFuBUWYHlwnipnNKijSAvhK9+hUquZh8fxp9M5/u+Fw63DVBcua6L11+QJ1p
m8Hcy/7lChzAIycWknG/OEPJabPCBkHK1ipb+6M10HL5ulCqODpsCu/68iUdGxSg
8rxtZGN70ANZFaMil0WdjuoAa5jx7LX0E9Q2tIX2UflTwrProk/BGPNffyDJosET
sRtC3rdWpdrHX4YGhLZLT8gKkGeyP/n42SylevGkWs7/vJxE5ZoqWrpaejL7f/8B
9OgpAP5NfndPo9TDiFSYBoI8uIiaP/UlGx2ttLZK0S6HJVfAvL8mayWQPG3BSAsa
mGUfekfXvOUzJ3pPudEHKyhVySRc5y9oQV/xESqb60JRI6aX3ZWuBEa/J/xcc6vJ
Z8Y355XM3e+JhrVXiIgNGyxFmYQvXuTZANkrEhfcu+ZpNZe6+ahc5U3NDn0tsnsa
CxhLXSUqfOXfnz9Mp7Fv5Qj9KH4qGZ0C/emPF87/sHjlvQiPKjeSr85dZzr+/UJd
KTU7j265lb82Baxat5TdGTRv+oa6hFK6aEwD3RX/RyXZB771H8KUiIPFyDIGMWik
qqKh0pc8Day2RDMpbqvaF9RnLRTUBs6JPE6SxVVWC0Ya+Awp4GLf5BbNfChFuSBV
hHewqaT8NfyxmeuvhR0ulqPBR3rzmwg0d+1WGiJ4avLtWWNvxZx8O0kEitzTNXZL
w0ZKdVEqljvEUtsgot6+zCJYDSKHBaMnOa0fik6enkQiHWKSWwCDPa7BLXNLvQkQ
j8eSpgWQ+AcrOdzCA50xdT8CfF1VVSDkKyx56yFXIb84deweiNxgM609ZfbMiVps
JUmTzA+5MAwT4KLsx1ElZLAf0GBshpZwq7nUd07Pe1OU6p+IMzM5y9WZ7OeycPrF
O4fRSirtuDSr0X7tOUdTIVilfPkKxc17Hbqg4dEH1/QVQg+avqqtNoj3af6l8yAS
b7k30YMaRn2XazBX9a3PUF3LLkGQ/NkN2zxepuCzTc2WIxLpEWjp3Kf/q9EZEQUn
hMVwDYwtlm/ZyoWjqy/Ppnc8KmbG5r69UN3FXSLyYWb+1jsAGtYp/Hgm4y5rlCYc
Yku09KmzAGSrLWoCxrhmbzTtp3KoxZaEixgc96Nj690OzL63RyIs1g7FsJjkX7oH
HW6i7tVnEyCk1YBX6ianLckzk7wFzbfH7zrHNB/N8EKH8Pq1UBo+mSqvln2/USUu
AEAoud9etPMXBVYRMi6xK9x5g/bL1EuW0D/olAK/BLZ8R0grnEDYXN8T02vJUPBr
z6JkVMlM63XWdGfmPOMkzEl9/+JqTF+6paIP0tOohTPC+eZ+zhVcRsfCLbSSxCYF
espeGD2SOEqJOXcSDIm6TLpGrjJT0+T0VhY7JXTagSdswhHDkF+1S8wUP9X6+uNU
XurxFZqQWRbsmI1c8l3bqD+MTl+DBSvrB27sC9Dij3ogDLNvNlyk5bnog2syIBvw
xuPKEYtBfmGivJaQFnmcstFfPDnlTzGtI3Hm+BS0psWbwOa7wfGZeTAXOcnBJPPw
xwwyQ0/Y3arrBoUROoSnJy5ZCdocc0P7TdyOiETeX9EaCrLXg/Vx+4T0MUhz/Sxa
CNR1oFETJAGYcnbZcB7I/5qMDEYmDmhOJeklphxQqmH9klvxLkezeuew6KKfJZxT
gd8zxEEKHq3Lbf+DCoc3flvQjElIj8ut8TNmsMXe+gS9QUAIf+HYJaz+BviKOtQe
BZZwYxKDbxtTMGjuGt1ljTFxRaKDNfO0CV7QBBf4A+xUh7jPYXUeIomdK/N1VW+S
Po2EoD1O3LiClnMH/Yzd+uRaJ9OjuBcTPtzH/8WgT6zQXFDCTTQXABu7w8pHI6bR
6vzMC8Lx1itqIhQxRTCJVleoiGiOZzywmvoCB+wxgpNxgxj8cc3PI7Lq9WEtmUsv
wdHUy0l8WoMlIAyunf6o59WC3iDy/zsYqpF22cymMvYhU00R8lhXoPFiN7AUAPkc
NLIrBvMUSVwmMJrozUlKgrfIldDUzSFSd/QcLMMh8o7cBLSkqzT4Y+vXejjP3jbC
znHb6jUEOck5CrOSoGwNC+dOpiBJ0t6SqNRFAj89pFTbLsZ3qJI/zC09aR9ZtulJ
CmHjwReih+UGwF9sEqjn44xRTsDje04Bumaf1hfHk42+CQQS1HBz2PgTEc6szzro
TtxRXieb6CY+laiUPfXXeB6GzI6lskTkUSFUx2sE9WfxEfjqnbFrwqQvtSM2JbZX
nZ2s/D1qCQV08nvBXqb60yTh4s5/JrhDrjgZ9Hu62+IRv6olxY+sZ9mUXCuHN6ND
O1NQugUs08Lk9I4TuFKPtauJ4GYEZEUWmV1pymyObnamZfAgAVP2tV4Wtx9I02+T
9/NR8P2snPVE6pneDbge1D7De/GaSQfF+MsGx+/xaJQggwx4rrpG+kzLzFHQo4BJ
nYlKT5zVa2pDMY8KyKRUzLYnSSG5Apogvf8QqsP6On6VMXuDvC6PyNkTa2uhKyrf
kb5M/7ounEXKyDImL+92CikaL5IKEsorsK3PrgSJPMDHRXDD1+pAxJqB+Or+8FR1
Q8Ov7sQ8bZHu3Voa3aUnSKOdqe1ByvaZQ8KeAGLzAjPuKz1zliN+l94cI7uuT6d2
BlU9ynhDwN/0ZhhDFOIFEZDbIrifnecoMdsZhMvmk+BTVvyfhA6K1Oac+lrW2/E3
OTvakNnfsM5PeyW0+2rhdXXIHXvxzQ1nv8SqBvO/LkSxr429h2l8pcgH7IoVgvMK
+YCjewhTlKCyDOfTS1yWM7QXk6lkpHG8tKl94LKKcpoCRY7+GnJOY3yYo4kTfaoW
8xvZ1nbJTRP1UrefJEeXdYhiG225f4cke412CBrHlqB9T46Mck6CS2WgogTxzJDa
T4OlFqZ5YxoCUZ7AFV33lIXSNV1vN078k/D3hyJnwjLziGeFahupX3HQ+ogs7UOp
T4Ch6ch80uOxM7deZxRa5zYR3w+VCmjEDEcv1UWBUUfMQRsVP5E1snqMR4nhJ1Pw
192XsmuinHW8NWNzOwvb78Vx9Jg4x1D1zJ6zqXRmmTjCyAJxrbf76RQaS1KXmbPy
bIWoEN0S6bNWeJ4Bvmx+i3ObbjYvRbiDwWRFRM+5A5/Ej/Mv7WaOWAqU1BsT8bA0
NiEcfnMiFsZCMm26wv7V7+JmdC8A9en35ZoE4VqZdl6JEuaPNFRdeZQai2N6yjXy
B6R9HaFYLc6dMzOt4XeXqEXKQmWB/LAgSDzZwnq94Ih/reMLpAOfsAbP0yK/nUod
BDwSjE3/4p5PAHLYYHldwLuaktylVz1X5+i4lb3TLY/XxEKjn50JQyWeLv0BT0JN
wsxXKfYpWeSKO+qnEKHY0JWBp2NysibsbMxKF4UiH+1gxwHLVagk3e+pvHPzJhSA
akN1xCyhHijsdvZyW5xkF0muH52+4DO6EeP712p6jjJ2nLd7SB+evUgVTpINWof/
ths3cSg7Uo1jeouOzqpQrORFKYsMCX9TZyQyFGmvmiKeYJX2Z8uqbjOqoJmKzka1
5Dcv5bXHha+PmX5yom6FQr5kqjc4q3VvE78hsDSBUyEvAE7WrTLN/duFSLppyC+x
GqPkssUPC1j/thbUfsslfCqtjm/29DrYNuOcht6tvxLB1CgM6Mu0lY0Mg77F+jE2
fSqhQ7yblkQU8fkKhBMd5DLZ8c9n4DjpTX1QapDHTr2mZ+veXu6YDSN2Ne360HmD
enJy7aeDAy1iTBskFoaXM6mLd+DPsZ8sM6+vJCcU06GoxG0QxBt3mtqHc5a5MaZY
fCV2IdjiLu1ScQ70/mxP43kxLJ4UdmoGVhI2pispI/x0Q/zeyM2FOekRu5+t7G6p
dZn+o5fN7Kldlp4J1h3Mp1byFbc5DUPw1WlEdEea2qB3cVEugFeX8ZpCXlaWBLms
EMNIyMucu+S+D4sd1zV8lQ5TYXnQCOL6hKs84q/PUzhzYjForvTqWiMQ7WuAeksn
XI1LbsR/xXNZjNrzlN+ztvEnRM1zZfR7ADYtjoMMU0baUXVcqMth8zG5Z4PJYSUo
FImAtY9LJ2cFrOgky1kIYUA3lMoWFawFXmRTb7e0E0RCpjRD/sw5xD5S9uZ/R08O
eTzRLhA91OWvVUKWtJF0Bd+1y58Rr0ocM/IImj0cEJgBYKUCFsDO5+7Kr+w+8CGS
96zy//R8IxELZFZZWR1OaUzoLB6I6o+UXWlrl6FphQZ1vU+vm3CKv1muwrFdo/H5
li3w5hFA2CDSh5+o2eIf83WU1Ox0RTB2fM99kRqBn5+Ffj88SMhET2/KSc/UBOfI
E4DsqYLwSf0qwrJuos4ZLdIRMQEl1YsYBFXja6Iw8qBE18vjTue0miEBMC+//DHC
+HnM2BJWp585YOKx1g7D9Ez039ij9F4xkIHdH22m+PWmyJsIoA1hewLXLesqYgmk
/8d9YXOt5TjIJscGTpgmbVV3V8UAbeL9M0RF+O7qe5jC1YADsf1bwK2kGQXwZN9d
G5trq5Y9AR4XX2cWwl2iVv+ahoHi02h8w4N2Hut55XgfqVGIgdE0DTOth7PYXdJ4
bSSj4IF5h+Bim+5F60vY/K1FKWb6MUjIj160gLuwrA/IsuJxaZN3SPPl/+aXAqoT
uezZoDofSz5EvOB0cOYmtU7474Og191tpqJF3A+wAkk/kBh2RhWWEgyHawTd5fWs
fT+RFHFz8vSV5lA3sLb32Ds00860UcHixgdRETuQJ6ykbTvOP45f6OCl9DC3zPf8
9/q2dWOEYuE6l+D8YvYEDAE5tEdEIafOKwAH4cj9sDWUzHK5kO26aKyBuBXhoLx4
LPzMNukcHUMVjvRaIZoFt0UfSOtn+4kI7ht+PSblRrexznIkQMefyiJ8bjXwkeSE
pTaSRaQHsMeYqnVVBlA2DpDH36NLeEoY9K0zsJOeuEMJEN+Zvx+fqVzZM5kGp/M1
8+LjaaE5nGTr5oNkMG0RnHDXcEQPm24D41mTjMdcgW6dpbjCm+jZ6uRO1nh/sz5e
uSXQyLhOAU5KfJw7yGXktqutC52rJTfQ3WTWI4t1iYRympgVSfMb3OTK18WrFOPa
GpgBy8WHNVjddprpN37fjTYtxLpJlAt+OcT3O2QBESHuLlwk7CxykXi0ZDIEElWu
xW9MAV7XDgV4oIK1XQYr4ZLqp3JThdbt7UXP5GwZmB4uElLow4BO02kSXrHVHt4F
adOjEQ223Yhim9kaIoLLWf7wTCqNghNFugsAwAt8hlzcbK5CgF2C7KZ2yRJf6XCv
DPZkrKY15awi4y3DwM5PhETZ8J5J34O35qh14n9IsXzpGehFGnm8duFGfnBNc4c5
iho5jEnhZKUj4bLZpwUMfVtMcxBtpI8l1NjBhsNpnc9ryYtSCSvQeRTJrlv4SiY/
W/UX6AG/2U9makEitvc0XcWxMRcpTQd2fpX6wKToUMT02sorxJy9VUJjcYbCYoxo
6edjwfCtPCN+Hn5H2Cug51nnhvOQGt9p5z/gyPyhRQQKMQ/YmW1omM8wYSX+7gV5
MB+HDoSxAq4Nxwoiv0269zln/Jb5w00FV1vQJVTdsiDLHh+mfC5IekKdvbIGVuSC
T0/nT1swNQ0E7gpJfuC96WwznUjIzouXsMKsmc36YM6JtwDFaqU5mfiNKbKNPkef
+VQNni5kRyN/Qk92PAScPiO4+De+R7FzwAxCcO+CEPx0uvhQIU2wHhYzuCiFNI4Q
y/KiEk8pPNhhROaLeP2xk3QNnlGtPCFXNYhAhhDxCy8+njy5fMbWRtdku+r6gIk3
njx64niTr5Z4tdpvuMIw+Ioxw6Qbi7L847PC5tFTRrFahO0t7kuAFltRsJvT0YZX
HopTql6OEaeQkadcupEu7OWrg+hhXFi1OLBis5Pb01mIV0eHmBT+61zGaGpXfD5c
sMgUQ1BFdfJrGj6R6zc667WYGpSKNLApnKuuqnGJZVE1bLyOkwBZhcfHcuPEG1BS
HzqnAVlMyIuhpOnhnlCRKBlWRogFOMt8TK2NPhsjRJKOYGcsArotPbc5zzK8rynm
m8Y+NlRyA16Dze+/aKqGBtn2HaSvrjaIW93eQO0FegizTaFJuGFwN7w+qhXfIzHp
4MSoPactApOmXkJvLW4aQpSRacT3fe2WxmY2jhAAy10Wkts+sENjmyuFagsDcc2q
axS6UWgvj07O5o4UZDEhYlNVMZql4u9db3xuEe1BZAjrj37E7HCRJm73suX3MBis
/s3prW+7uvw5uIcIuA6MyzM8Gj9UCRd788HHksDpDBQnjC8AqleZBBe63olZaK5q
E/vCekCAJZEZn1Q3WGpUOVwc1A8n5PkpLaOcE2RXcGS0/Dp82uRn1A+Y97VRsgwU
tSLy0NaGdBI8Tbh3TCERXx5uSkbhk7yW0rkPcGnLnQQn8XGoKFPuYDojz0hA0sVl
Rda2f/M5xmalK2vl6ZvWHjMsRZwonp/0vGmu2xusZm5gm3qFvkgEaeVdFBim11rX
L/OzFMRX+LLK7glyCQrJvNRCgjuM8WUhVMFqYxygggwnwNhqeMNuumM0fnQMUHTg
CntwP3yIndxhE1WO47EdGDaVXpu1/ZLBpshXSnv77Y4qArPo1k61tXG46MeHm3Tt
8/apeHV8keJiRosNICCw5uTrHTunFXreMZHwTJR2x2vpvMQRoWHLlqqASlvdejQE
r67pS0wgqyavUPjFu9p7oYRGhy3en9vZ04JsfOlT2Q9NDAz+B552AEhxZ/VF3nT+
KjZ9owB47Wi4OiewdoeTM41ydq1Uzq0a8sp2q3EsQBlQmlGKX48jJyBjONQZQ+2j
jqh8+NOelah63RS4dA4lZb7pz6QVC0t0iwcJ0nip9gi8guOLDIUOo22QbOqZxf6j
aOCndHAhR/kXssZW72XxlgDP2j8EFVuSpg8ohKJACD/oJzKKkniT1Q0faWxhMnBh
Ic85VD8hED4gjzcFW3x9mFtsrO7fYuFAhWk+E2b6HTo15yWUoPs2XfI/2jMJOfBN
G4RleA5U9wr5NjdG4gbccwnEjoc63GCIIioBi9z9hyBHpoXDgwvtaZjF4h9pnQZi
0mkd0L4vEOMml6p0CB8oxt2H5+PQMoQ6eSp8jfiyH/TDdOHgHEHfaZLMoMlfjPb8
ptAxLpMDlnL2hX1YubfqteVq43/6w0hu6cw1qzWZF3ITDYgL3VauxrsXGmGWAXCJ
RYN9jXU+dkQJKTkzNDYobm2DK5HmI84lipKldCr904SEpS+W0MzW1a5H+OhKYKjE
KdT0xxAw+RsasxU4dKyA9AxLmB06tb3h3H3taNFTkqkMly4azAvnmQAkxA8m6e9V
V53nh8pIoHlv1r2WbbIacbusY+1yTDz1r86LA6aHOyMJ0gcgvQTDxGCoKOducn5n
tVVSdzKoSljBDE5O/UhC2OMoqaDibZ0dGbzLjn5BmMGzWiFHaJCBMO24pDJ9zL1F
kwYkqPICrjEbnQQGTBTJSROiAwOmR1xnjJrUAaZmhrwCz3iF175it2bwN1uvVJKQ
VoogBnumLsyEUrhFexxp1LRMfRRU8kJHx+JNlCJv3mAuzseXbo+mwhJClNuwGJgQ
fcK2KbR5JwpvxJRJcrMAX7V7KIbDtrcwfjoitTjUmuTrgbFSd7ZPW6am2AE1sJhX
6eHBb2CqpbeN4dH/0qP687zlZjt4Z0qH4Rh8M5EDeeG1nKnrMnkVilrPS3EhP2BZ
EDF8oMkv6JooPd3rmpP8aIKlZVYSTLZHWkqASlyv5WkmKC7zYOX895QQue1qcLB/
0R+62qD25i2lNdkFebkEkCoi0EujEIaNlDfVNgrAogisMTquYsYRbzAVAg+NXXsa
MWZiUuZrmOEe5bpwHFiwG+DcQruXaKBU225SADuFW5/WIfamwQJHnwkZs7mkkFO4
87oZ4R0Wp2HyZ97aFps0Iz8L2oQXfA54e8VNJ32YlG9nbcXPCAGg3U2kRPdOhuyJ
MvZpfdMJrdCKFFZtFlxthZbrQyVhmY8TDnmQ8cygparAAzDkGn0Ks+zNqxhoN7x6
lifAiEL/Q81LgbZ3E+itaPxTbTymqoM44EQKiU7Gi/zrTY4Vn4P3OR3D0XzpPIrn
GxP7lJCyTXqJm8nQGaxsWdoYUViyJes6gxuZgxq81KOV6cT07W+tCuJ6RdDP4AP1
+zc0bFN1CqKc761+QS3vLdJh/o0AMbIGuhoRuRNte0aqzfbSrvfsR/zjz8Gj3r2/
Je0t40N00yvFu/KskPNsON5myUt0Bs0pwzjJCJlbB3m/VqKWhYGMYkx7eww2pZ2r
rJRczdYMPJKxdmFsdKgyceT2SCRRGShZAvrkDZl1g1PvsoUo+uGJZv6TOnIcN++r
xi3GOZ3Le2ywnrcembpw1gy2/4t81MsRU8wsyQnH5EN7y3RT2Ymlqmik6P51pquK
lyAaHm0zPt2pijvUK7bQMUNiW8nImDXBQRpn657ynuvOIv7pp+1axGc1dv0kOiYj
X/EVBXZgErDeEILzP4b8euVPuUH0KMxM4tdMU1CLzmPpz9j+e9w0sxIFDVIxo2ZP
5QJonlYYzNurLqx9wgATCp7spd6zjTi51zA29VSXnjeDkU2tSDNVfe18AnlkS1rS
i7L0CILY5AMscQx+rzjhO9+evsDCeUxl73f9G3Z23qeffTVXZBKsAPOHU1EYWMfE
xHiFH5p1XjemAUNWl7LrAOdD10J9ZzyNABo+1xqaOao/6cv1UGva2LB4qJtmnMyg
bIFB2ptyPPXd/Zw7PHC8pa1h+uJnkXJgK8p3lws3kGH1nwi04zh3Oe9ewrwW0Wb0
gBl0Tuz74rn4SDFl6BdLqKU/Z3FbH21lraHp/wG1ULVSMnam5Xu8ezSHpg0NQfJ3
BOajlNsr7CAClQna/3s8X6Lfwy/jvYo6gRbyS1l0Ocz4PQLmfkrY28o9VVTlsw0W
SXS7uBKJWB3PHe8fQn26kevZvZjpLXsKwvOX+pHjHp95wKlKy2IqCvuUq+l0rd6e
vm4snEnJusZNAekVZcBD5rjNF/faWh8URawf07xHdoyoiQOboX8QftHd3hdO1k14
x1w5ysYElgJFPlDdC+EpIx9ByPmAQLL8aAswIjzh8i+R6o1Dvnka5WpF91ZJ7GLb
zQpjfXthb2lUq+DrdTYYe738fzbmr1BkRdPAGoWweT4UjE5U009HENpDuvtrS+vT
IdlpPCX9TskyD5CJGSEu1az9mNTV2ayGdQ7f9NealFDuk5TCR27OZ5S9bkEiyN/w
/F++40oqQ3L7lNJu34qfMFhSHQOSkgSjQlYUbH9t/Uvku+4uBRH/cHyZuJb1+4uX
cuptDbI55u4KJerlfdAj31yLyjzWsYmMjqoBlQkoJEMGM+sqOp0R3MAaQDlfQM6c
lGCe6Qd2t7+Xz2+CJmHONcCr0JHw8sBA1vReG0cxjUbLMcQPb+c8QJxSWmuy9Ma1
vGnVfA847Pp9L6OIHo1cyDj2oKVUA02K3RDd0+8ASqYK6VqJOvGFA8OjBUUfT2pI
k42C9d1tTAkHI7Gk18INBGs2JVWkEwUx4ac6TD3RZ0WmEO4RIlLyo5hLs9XACz30
aKkEqqP2FBvuZrxDOQY8ZJNLcYxTcbZDn4SjzQIX12MHb9f27eDP7UvBv7ba4qHu
vxN3WBgekVYyXHo8rwvE25r5mIscIpmUI3bIx4GaQgLUxTg2gk6rkq84IF/dBu5f
Mw/2LKw7tgUZmaM8JfeLzXSbHwO0bBjGuS/XoSAx9rBwGgv6p0nRySZZESFJHfP1
oZ1wTottA0pmMS8YNn5ohhXDpQ9wXzHFAFL6zpcNGTeAA4eZHMOEWD1/lfKOEnBw
0+ZoZ3cOLTDWlSd8pSurwyrI7AyDOoZMqL6fsQnRIxxFL9hOu03/0nPlFXW6RQzz
AjWVuCuW68W+6MSEa9syAZ3rHGbM09RyuohD9XqCdgl8JbyBewqZqbK5XBLMAe4T
81ceGMWIOJ/zBjsZ1Lnh5Mq0VDFnbEuLOss6YZr9vOQwfSlFIzNc3PZRrMlF87R+
2DNl83Usvt/If+hYeZOYGB0WMC7NrE0liNpJ0VEpqI8la81+zhEA2ATHGmQPZLcR
iliOQUjruAIkQzaocAAjY0PLW2xAO3QKeLthmvw39tit6iiZqjz38kwjfZw05vIX
2YwIp8dfo1j7+SmqeHivjXTpTr6dyLFtdHvWn2dDQefGkcdJTpQH3HKZIpCePnOU
oVfjd3ewmxRvrAT6BnwqrDtLQkwfA2fGJWlR5OgPnxDHg+O22IcmYCaxOLgs9vL6
wHaG4/tOSWbHDHxVDV1RQH5zIMXPNW2GsULAp+Apo8C1Dp672IDP9nta7eNLDkBl
LASl+EOqfSrIoEPAluiwxT+ajpebXz0BxHoJWZmolqVvVM2yOPbB2TaGZ/xG/gbK
baGg+ts4SAmnCAetJLYLRB/nBQvODp1HOwytqALr2Ek6N3xYhcMagIfmfDMb73Uj
IU+ASkvSdYL9Qa2zNjKXw+3da2KWGAicyYZe6e7KjTQIOtT5k1DwBxOuF4KJcWUR
QAMT0C3pYWVysM2sHTZTyw==
`pragma protect end_protected
