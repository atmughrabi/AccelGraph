// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PuKLIJa6+3RO9lXM0r0AXtzNZKjT33dq+EW2xAdjvnj6/gzh50M/z46BOhNlIYdH
8aVRdkTovyXEAFb6hYQhiMX7H4ntjyiiJukSi9mIAT4GCc/PwSJUk41wvVQOoSZ2
Jc0cZERnHUIUvqxXc762+7CjM+sa6ajDPSGD7Af6Yso=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6976)
ssEeIZZb9kstkH3Og8D+8HpH1pdPH+Uy4FIxrV77v1YSJSbQQmUGT7TIfbhn1oEy
nqSxtqEolepPraCvUH5/eJgxr0NVa2VhwIDLe+FWg8TJZ74IbnRQajTnU0eOHzoL
h/cyjn4iPTe2BYSOiL5SG3u00nG87266csfoq0IPkliGx1xyAD8CnufKUvP+b3Bj
Z/lm4wVPfyfBCtxlUNHbAtCCI5qLcr/MfFzyybKnXx5BWYwG8w3T0t/BqqU67EFp
tVrNTUWPyFMXBTLSrE2E82/72Ncicn2HnKQ4F1ybMSfIPot9TFJ5ZMW4+jKErvce
d4MlneAJJrI3CDIvamutvEhXW6JDcql7HxnzwWxh+qcMpJ//ElVaw0cs/YJYl9+n
GBjXOjKC1h4GlhjLeGeIUB8YirPIbUhLxKAOjqnEXCeQj/qK30fuAW7iwSdOybPw
ceJk4s+ajcqkgoIIdbZSIxHwMhHP/qUHtuYkMk4GraFBO/tNQRhTVuuPz8TDUlHw
E3pbSW83jM2xV7G4eY34QU5F7geO/7lPvlh4LeDOxeodoo9Zqxl0BDmvrMgJPsfz
fXB/UqDKQPLVL+AIW0/tivM3bkOHGb/cxsy4pboVh2S69Y6BpN6Iso9p0cyj91IJ
6/sldeeE29n4aIjTlp4noRNUtcoHVytJZW9fMKorW4rFMVZIehLexOlSGiD3dFhQ
cxd6JNnN4tZdX/Y2+fTU8zl5D5jjkwnlNQ+3HogBPr+E69frBhreG3ARraEtbL8L
EpLwBXgUZcW1A5tW+3xFXcTKbHg6FDLjQ5lKKPfOg2jeOYiP/mTtTXWtqVR1g1zs
aEteDYQUr8XmDMmpPon2+wK9ME63+Tw3J8RCegFgKtYpq9XW8kVkRjKd3UhTto8o
TSO5PKratTjzZrj6noNZqDi8NUltAg8+7NlCWxvY5UfgAZZB7BeJkzSZ8gIeginO
GVWZjsn8LqfhsgCQcbRJBL3iinXmsWohd8ot0opwbDX2FZGNo6VsU80yJ+AS0PLx
WfdVmMgE47H4LSeV0GoEpzOBEh5Ahcmzy7G8a06zXB2raif5GR9J3xa0hkVkDuCz
a/Q3JQZr92VlI/ki3naLpK/JldQ47PkFNl1VYbR87mRjwqY1VeHqXt3VhD5UVPpn
v5Ia+pA7udR7BT+Ms5T79UFZIjDujAHevmEl1xenDDxYmzBgJp2hM/5LFFgTNkP/
X+YrZqsl9ZaGdc2G1419IrrWX7OG/ZuiyV4lMNHWd5KSq8yEIHYXupG5TjJt8gTJ
EtBW7+udrPTPKYDl2ydlmlW9g6s+kM1HRdnNAVA88zAuawxXEYoIAfiW4MBXEEaF
2z6a7zgf0iCa7iSNytLQ8MWM5cMOIwOdRsqyz/U/4tSQpf9pT6YKq4xgz5hmrkmW
05bY18jvw0aBm2DgGduLi20cZQv3ov0i1fsSU/8Uz2yN9DfXMFhc2rFOz+gcmamC
0+NN7vnsfC9vEa4XGI4/VErsBtvygQyK9m0LYJMWl01Pe8PAFLuGs5DniGjaTBOi
L79EJg8QkjVLNShAyqr+nPkGEthMT2h0uJWgfq6zQvozmg7TrhU4kEk5fScaKcve
0IZpQ9EuSg31HD3g9O3ThLJe5kxQopLH529EdBh/d5/fZYRo9FGcw/QdCyz1rP7M
g0im3q90K6BNl6WFJ18hdsF+FZSlDCCQrP+LMsYx3DTVcXOdCbR9PRHa7aVsN18H
xXFJz4X+DEVIxRuRKcR1PyR6h+ps3GBLjsUwwBy737CqKPnH1XeoSdSTjsDDLJCY
YDVU3YVp8j5o/KwqSAluifGkg40Fny1M2DYJJhqKwV4PpY7mdlNAOAUskl5ykDs5
UFNsaYQphQlCf9hpWS1Yx6B1bb8easAdXrJGtic2/uBZbvTwqp4o+61b93NYE8cN
KlaIZAf3hGmAVNoFDGhlGinwkI48DnXdMHaKZTMxlkhBfsFcO+nMMtOODbS2SfXu
s7ylK83D5ChCN9BgT8/cQc5a2dEEYWoOkt+aJ9zxX/wKmYYmyZvsVgDxhboX5T9C
QEzQIcqfDhI5VrSsK1yAmkhtVeyiNPPSxHBvwOrQ+f95Ab6tK0DivZdPlAFvmUgj
VD+MuXUVE/hofSBQ/ZXUlqL3cig83mHY3v8SzHbVdNK9mXVj2wdoS39Qm3EM6/vy
a5XuCKJGPQtMlsDN6OxJdNPaYnUve7bqxgmMBVs4xulnmN7Mg9UKNTuEkioN8FGv
6YSI9BsOxmilkFUQBIHhP0XdlPyF1JRui64pI53C/0zuF8lbQEzikn7tBqml3rv5
y6v7XATQ+XnHMmLkZMOuuBwBq1Q4z7FUXjQ5OtfGCJIE+K8x8prHTILWB582b2gp
YlKojyVcE5Pde6e+Z/CsUGtH0YFDFZPIH3iG8TeIDG3O1XQVDcpjo/t/++iFHeLt
acM+mwUMT9OY/TchdUc65fHhQ4dYjgML+sR8eeUjbwNRTWaP+s43V9cWnmaOZf6s
lzxU8rBUPUh86JD2S8IregYa/jyELK5mPgD2Afkx5AFheL8uK/47811nsEXwewFV
ZLGETVxz4VtVZgbB+B0yu+M8xzCj9h3f6UExV7QlEfI4ah9BaEGE8Gx21m0CfUcl
oKkEevc8ls84YyqKbuLT2I33Zlu0N33rMt+yjDz1QaYcRQsXRQObOKfZ/CQiviSd
u7tAjApBoQOEYzkbqVbfNELExPq8TqqD5ekz+IxY/T2gC9PGgs791APxQ1fMJDAA
Jk7u9g/+6JIjl25NH6LdABY4V0hauu6YNxXom4qteae15+IEqebbaBXGFVPesxHn
vdON6Gdg/L24efu3K9p5QQonB8+6cWsLyDZV1T9Og3nMyBdqMwy1Ri3mvYqX44RL
A//nRaGBI3UU3O2oJwZHpnexfkjeoX4qsDwD5ojxK1+R2VB2DpAu/uBAQCBjwm1D
3dnMpz3WuxTIGw6Ga+ZSn+2SY1LhEb5EAfJ3O2M5f20j2HpffzFc7H8r5rI3kYHw
K459Aq7sqKcbJ82kLofk5C1nT9vnYgRE4hTIDM6h9qYI89JRlRBnfJYzMWQ0sjjw
YhYTAAtQlJqzSqXcrfa9NdGub02T6vG/Zlk79Xt+Eji8OBWqPgqr8NneSoTG7NKB
S/GOpwJsaPh+oD0kLTzggrB89GhMET1XhgJwmSUqYiTobeIfBmtyAB/Cppev1kp/
d8rwxFawAubkgCUdOrvOkI4imJ2+1jBRf+C1715PCX2802gnFDLaJs/QElDCABeA
gj3+fDirus8zEiIP9jiYZsXmwi4LxbDxOPO+bcFBefyP6cCk+Gy8auDlYelPL9/a
KOQKK+kdTmGOehQjmR64D7G+2zI+OHzrfPkzcLVLUJjEZUZfWazJe5IF7iRFmKxF
wG5yu8laMRyvVNY46U1EjaTBCcOnp2+YfeUxYK5SWyJgKOBPMPgY6TXvGlHbCZQe
QWu3UTdeGLANAkxRVtwe2MRnpxxUaOQ5LS+9Vrel4pG6C1VjbZPzOIqLeY06ZH14
dGpaX19gi8tD+fL98kevT9K/x0TEyd8fK3hLoxVThhwPDqRFlCbyk5Q2xPHkDOQ3
5d9KkV7rgnqbtAr8FfhcQa9/Yk/W/pUp5uSjGvs5Yqq8i3W2RajWh0mG3QZaNxWi
uPXzn7y9YC0LfYkih4LXCs5lvFu++5CnXy1TUec27y02wOqM8TbEGx2zgCuaNnQ0
T2mUE+sWzq7Vl+0x2izH9AeIW5z+2KwHOCM2EXGJZSXxLp6IwpdvoWfJVzLsJKgM
vbucbyk/WIR6VJltCqJx0hp700U7LjoVxAkg+ePc4uDVI1duMswnsrnDFR3Y9P4K
owU9FIv+GFe5/w/Gi6vS4mRukeU6TZMy4ixF1N7envT1fpiQrTHkOWakK80NPqln
o7xsz0HwgsaTfda6Ehs16ilB4cLb3hwI0B7uDxFf2wMgEZRbZVqxvnvIZ0BzTg7T
8S364DZleYypBKs7iaArfy+1ixiuoUyNj7nThQ0mpe7iY3i6mXccfM2YRUYgTlkP
6Cqi+2em2vx8yuDSTrAF80jdjly0MKAwKd58b3V/HDhVaWpORPnzhyErP4YQhDOk
2neSg8qlLYF8KpKKGgZUnsGsrL63Iz6UOcOeqcQoBaAGngQjDtRnBt72BlCFj2ud
N7FWnO4ZlPcspuQ6PNIkbYbztNHR8TYK/hr/YpjpBduHsz9a8qCkksdVEe7SvhPR
bCZ+GIq0t8x1Vp13gIF0TTzkuW+tfhKnXsmd5Hk7MncsffrW+bwN8ABegXpquZAk
EMFsDJnS753va6ckBcoBqHAs5BszzHgo37QlGvoWLzBYkVFlgg9ycWYhTSyqzIgH
/ptucxMmdqvBdB+DiZA2oW0meXIj40ByrBy0X8IL9LK+1eikz3MgMvHkjQnTgSLa
DNrWxLxuM5pvBAKmJSweu4IUIyATQLK/YS6ep3L81Nw6tb4wdePn4JAH8FJ71sln
u1Ny3PhWy5q/yV525HvsV65/dxbYbc1mk/PukPLfN6uTr4nCDWWYhqhNlboOxBts
iWKq9cH7SnrjTmycHv13t4JQRCXuXTql2vDs5oCKSOMqCL5AinQ/zO1OiDnjZbaS
BXfyR+iRDPjZphxS/4LzGT8Yn4IEkOQz3RN5z167Dgw+JahAaBrTpiujpamMivZv
u/qjmtxEtTMb2dxvAWDhi3Gr9mNHq/U5kfSBjA/iR/ZThO8s1eii6m9Xs8L+fhRb
X7iG7IY3xmG4lit+6rwqbR/6EUxmHAIiFoIJO8TDc2ybTcJkAlURwxwb6+lsUSRi
HFfbWbe8+PJa5k1pi78sdIEMY4J/knWrAoKdkrsiAZzKgYRnpd7z5I9JNiaVQwJ9
Om3gdJ+AXIoF0Yz00ctOYYk8ZhyEm8cK+1Xn9sIhLUI2yL28s9IVYLsbpRMVhmGE
Gwfn6NBDMcLvAo643MSwItU7yFSV5NBnpMCWy6FKB6/siy7Q9RDdOlW1pEoDeXQX
f8E4p67mah28H/miROlg5z8uqIT1mkR4u0LARLJPBLjyiudU7cAel7e6v1L8qhg6
s0GNcm5dQQSJkfxzg2LU9frd1fezNC8G6ZoA1J+5QD0B5pVfIufwPtXnuvH+gmvZ
p7WDLleBchgFELEJ+0AzT0TFhsKlsRp1MTu0YpTDJDS7o84ohr+jyAozIak0LLvQ
0iVDS6JViLAFnn6DlvvuqmLDYK20X3sGVV7p0W5/5pmww7D59CnqCgsZ2zhbSG6x
Kw31OUot93OKMplGDsbGOJwayVsr0jkxRcETB0PMWuBN4miKcuKUpgYre04x50sD
WlUalZpNfuaW+zfi4tCyvFfwgWs+1QzzfoyHjY6G5XMlPKKTflp2vam969B487Dl
9Yyfs8wiitBMwHVKJNgrFrYKexFRoWSc7b77eawLZocyXTL8KA3unONsi2RyWKIi
bXHVSXfffUuU/cRAYl32MURqTj6S/Ols5UcZyTEP4eCz0fBsJs+2Enow366CHP0/
u98zX6vLhaIXf5rR3UDtV38f7cUX8ESo9rdlm7UvyN07nBeSoGGp/sF9BioGiNTX
eISZgmxObsOID1HQVD9LoQnA9C0YQp1Ol5wlvEZsE7K+vy3Uy6WVTh2Rns2BxWvl
qGWmIxISYqpsejLX0D1d36HTBRw0xMLnVPB38kvgK7XxTtL7mj3jsajSFYUm1dOF
SdqcUwVDLXLgZ3Kie+aPHW2bjZULBv96RAUpBF6RCGrfOKTdF3CL36UU2bh5cT6h
bodIkB6DbcZTUgfx0/tByKKC4tirCS+72nPz22GijkM9gftXoFCZzRV/kZPYHMgF
8lduriXS56DvIlF4K2LY92fclghrwn9g1HlTG1EpNyeFDQiCye9EXjk6fCuCN0mW
N+aZ1IK3gPXtYlxRBaRJ2zVmhR5VdLUPv4RXTqqwHo4rNzWunTq5Eq8bz+tuFYcV
SSqYq3OpfnypE4fLspCdp3mbM26PMmJsNt+HWHzJmVb0unuancV5UAe8x4ZUYbRz
+Leg7LwXY8v5bvShv7KIL5Jr0z05tRXu7i95Y5DkufqXswhEibRx+p3fizSdrl8l
g2a3idszY/GDtHv5wApYDzbm0JBm4y3WS1og6nt8Vzjg3JEZJIwTs0i9XLoaCti0
Q9QWq1eShobankkIWaHmsjqOYipyYdOBRAS7qT/0VgfsQ/9JIuz4PkI9rznO4or4
G5zfoWQXaVAM2wmwX+PLL+zHs2XlR0qjm6fpwvMQi0vGrq4wowrcM4zpKfpbYAJe
rSxjw6ODJfuYBnZLJcPHQRGTbi1fxKfT08fFmBzm5lnwDpADZDrIkbY7IctjGZCM
lAp8j+9gK+A4zQN1IoIpOvtLq46IW8G/+238mm1YLhj19DTW+uXjdUfiqyrf8dLA
6bWYC6igjOVfMG2zL/+waQVGOespIsjFLXZhf8sxBwB/0qCl1zBAP4YcCIaot/lM
QZOyQvAZW/I8Hek/Vf+eMyA6RUqNUzuExfBZtX2PkjBmJzRmlxTB5cVIjxO4dTb+
Z1axrhU1yr59u0QaW7HGo4ioEfHko0N3SNFbPu51AwQHdQZ4OuLtDnqC9b9I9kik
tYwSUZXa4EjbeM0/2oXj2EP97mZp8lULRWDQE27aggYhTBlf92WFIhoKx7h4fzYm
1GEsL1IRk2efJksS/XKS1n/6wcKAnDkauWTv3bOrURq2VuT9MXYh+i2sju6t8H6E
GvHn+HUYM8m1ezGOR8YJ4COOs6tTixLiAd/qZEsz9X3BoZH1IVycdi5RP6UbQcg5
/OvIed0/Jg/yry7w2CMmaNXDBUBXjkbtFLilj4f8C8MFMZYRUYuxjtXE4ZObDefj
gOtPXluaEqzRM1vjuS3bFg2dCCDPyBpo3ur1OFWx6myscs4GWarPKHZvRct8Gi6I
q6mFRo+1KJlX2yOU+VRAfbGAwdAPTS0Q0Tl1BgcGmomSyuwMMsaBuS9V4Om1Ta6s
QjlrsfBwl1quW9VGMG97aH1bm7oNH9TO0M7jV4Axd9Xwhpg7YxPhUPowvXPuc7pt
yA2Dw8DTqcIuy0uERaKMyzfnQeZBebKZQDIr+3SWvndEfDznu8LiaCvIAm749nfv
urTxBJOkux1N7wMkwm3AvHpogBIBxiBDFG330zZlmJTBfd/PxAIZYI4dSdsUkdYH
H4M4Qi+PzyWD+H5Kd2SzOaGKrcaRGRDBOT9amqv8iuxrwQIP44Xj8+yHkBe8spWZ
1ksWfxeCM0AYOQVvaRofb1ldh5yiWJfPE4YesdViiaT+s5LRQ4hxuyGOB0lSfjxB
tMIPSZ+NRupoCVOVrqApoDAo8m+zJWjfECsK+oG/WDcTccZK+ZWpNjEwnDP7aBlz
aLDdQ5/tMfmY5ZyAsycJlxd5JCbEum2soWaORUuQpk0/YFeKY9+mSU+084BOKAX8
7AWoHdF5+1f0gbtHh3tjzjobKzV/wVZlZ0trDHztXUH2SrOJMXsN46y5HxsiiFHk
L2OY19Yb2rXlqofMf93HIqDcFUIPzkahmM74JJOznCs01wPlwDt3gSfaHkkp+IFR
SSCYW07QaCo9qGl968WLMD4P0OSpAboAdEL0aF1c4G+/XLj+oMkF3iIjkf+h3kO2
pn+giEy+8KlOGfxrH2su2Re60BAWFWTwp2dRXPWvo10nWeruJcPXDg+tz6O1U3Nc
bV/r1rW7roSZEBLDk+pbn4f5v5v5VmrpjJ+TYYPVDe+MqGOO2PjTJbcBG6Ag4KQV
7OwB56gD6jEXH3+AlKIFRj6PU1fhzcc7bB78ZvJ8W/rGjGQkNWFfnZ1o5SjEaxRu
np311rZdY37bfSeK5fm5F8zb4F1HfuQwEm2xdbK1zEyE4ryV67Xp5V9RTBtQhbTG
QbNHVQ+3sMJNv4kJxZ0LO+RHJFXsOfTaaNERM0JiiQ6/U9KkyU7jHeZZj2CuilFN
RVdt3iSTReXMzcE605ju5MUoE8G3uYEtrdonglRxRoidOYT0kxdzInpDrN05saw4
lP5RFP0fHhExxQAdIALGX7ps0I8Ka43GLexrsJXiLbThdgrpGFKtdP0uufT23PWt
C5utDVALQGtA8PMKsKEf6ceFqYn/xyq64lHNpw34rUlaziSkgau+BKfEIuzGjBfA
095CNo5bAmLoCN90knL1IpgwmnSUpeKj/jaMCDXMe0fyKfwMo0lD5dhh4fu9BNYf
Qge10zzm15/G20JR3tg56L8gPJcU+kSngFuVzG3Lykn1oJ/NV3unNYVrSDHHAcJ0
PK7qTJsittAvvYDsy4NjrUYiTaKlQ9I1CTkXxchth4jopLJXEYyPy3lt08BCmUtt
IYtKU/jaAWCGZkSZda6QnVANuAjydBNBBsHNnkZqiPqTJ9CE1qLVppivQGm5+oof
+wT/m8T0V/jhmp5nNQ/tJ7c5AygljhL8SQUvQMNDbWZeyjSX2oBUD9UsUo6EX87W
rfxF7LLP+OP1TDteCQY7Q55PjkWYVsEIATCY6oZcIgSub5rEuh/0EbvikvIXKg6w
IrmXz2hKVOLWh0dXcVnLXak2c/yYKrSfzu/Ztf7c/6avWsMNEW4GND3wOKxITjQD
iIh8b7KQcl+hgDk4tBy6W1UDe413utRMbtF0qXj73nqqL2L3v/4PWx80GstCK/0n
X+QOs/rx416ZB4Ri0HwRljJAvs82NJl5HgEoPuhbRu/2oJEsUUFmpGzr+aUQW3fd
oUAQrb/jqv5bGgkTjKGicM02quOnub4MVm69oW+2wnSKzIQvutY2wyPVvYywCP8g
tSpzM/j3Ikl44A7AVrjl4yGhR+ACL0Of4mNODSx9JjiJlUWO4bapptCq3PuIEST1
yCaxV2XfS3+plQJy6FBqwh/g84Q2fQa2xkQkZMZS8M+uWMryL0xcDiqJGHH/6nfJ
S88Q45BTqGqz8pp1y+FWrtSS5gqkf8JzW9MBbmwOHJcNe9XU19zpqxOyANAA5R2F
4zUvB/G/G+bLRfbKewF670ddvWtKEH5Suiu1/5REVOUNgNFwtyjWcvkZ4UmP4dtz
wm8aEAI6axG2scaNMOxhKhsi0BhD7RQshaEWQn9EG4oJzjgyhOh2hh/0f4Q+Eafn
FUpSGnZppoHtVn78XxPojKPs6xHfeexBzXXP5wkMpaXxK60otppoMe3FgRVWBILd
7APR2fzmJbCK87303IPnhqJy7RdhjkvORzVCG3vPuWIMGAeSJIR3/IWtjsVzxLef
VltEk25h+vfVxsk+oYzb1hOxPE3EWG2Rri276de+c5wyRScvd9KryD407zoVB0o9
QzU7O//JL7xR0BH/goNBxw==
`pragma protect end_protected
