// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Wg8Sh/CcIxvjeMXqdf7n306d+rzHP/Hc1M7Hv9QAetxIdoMRJ8xggWhrrIu7up59
MHt7IcFUFc8dWPNdYqZs9UqEaB6hNyGroJvtyimMBqfSisMXEG0hromzi3KJVf3K
yc2gVNoAJVmFwFqVLQo8BjrI3oZeD1ma+TlIvu8jYdY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19056)
gFxMQ9jjavDlm0AZJpBIEgDWLSLW5kFbTJJwJo2zGZ3/txiVGWANMWo9Ny2K42Bt
Cn7DGOBqMSsih7PK1hm1xSTqcO3qEQDJdRZmo7+KYxR0FdQxmQQdfzdBSZ7jNRTu
o+8FcBYKcORCHHVxHs1AmfHfDO5SDWwR2/fjKVy93aHLBhzElwVBaEY63pw48OYk
MbQ5dCGp8JMkvsHJdczCgpWI6kLsc11j3ihd50VsX+JTKR3utmFlZZNDdpv3h4DA
QE8bTexyiL9yuT+M10aBtjKqD9aaRFUSdnQxYkPMKFlMOdWOzaDEywX5jm4gUSaX
CZIkHTGfWbOoAWszRglPGgNYat0JSsCUZMSM5GROH43xmLwnA+N9GxZx15LCcBc7
LCwmAADigxRh7Z3NV0mPebxuCyIKBt+zumaXZ2F6pJKkyYSO6wXch9BwTniI0jen
DQnqFcNxWxFMu5tGrDNn+ZNy+wmdyC5or25GjX13/Q5zq+O1Fl/zVguQ6T/5vWos
jqIY/Vhl21RYBT8ii29w4Y4a7uKIRuWmXAICXbRMw6b5pG2xS+eWm/Yr9nn2ixuB
hTkjCs4nXIoTAm/VSwj69LRwac1w0FPDHrBKvsrSV1Qs+NVXHNXWynjVUb64kzNi
ie7BmT5g4IAOzX5RDd9HnjGV2MSPZ8ki0iR4FsdeJYDrkVwSORioDxx0BfofJNrF
vXBP2pRlGsRim5LTnYr5f4s3o6Y74wqepyPs+aT5OeH7rs0LG1hv5SEkqUp9x00C
qk8S8qZpjlV+WR6oN+Iu6LLAoBS5aTwSipJQKseYdnXnFBgcfnGrcEiZdwhey9Sp
0M64126RJpeVdO2XUqKMTuinLM/xLGAp6s1iC+ehXRuk8lmYOHSaSf5vsbDnkV1x
wW5iFNSSMLGIgp4+B02jyErVnM+3dvpehzLvwCZTOQIOMh17SXTsgNoSw9CcJPch
caEhAfIS/DNJOr34/pDGIEB5Wdv/JFx/FMSiufBXBMCHH4UrJe1cog8JcH+3OVt6
28hol3jLGnF4Gd2Wdnh0nyw7X0fCvten7JJlw0bLn5vmlLbsXPCuWQEvalIB97OT
wwz3JUX0ftXA73P+3AjTGQMOoV1Xycj8haJ8+hmtGlzMqjuFU/dHEdpe5hUOoYif
F3E11+mUyPL+k93p7ob48haZbWxihSCusG1xVfg4hzHFpRsqyB9j8zGiBdWIs4C/
Cm73XKupXeyKaVWmIWxLdaaPHRZ14I5pgIkBR3A+srUXSBZbHyQpyBomm9G5n65w
cu2Y2PmJRwABUfUgZD/DHT8OP8LR24hnGXoOGHzZo6VvAvgAgyhfcA/cGuCJUgNn
8t6O9jK4+s8m9kHLtV3msPrVe9+HcWrZzXWPKtmj3ZKJzD9DtEdXjh84IxoqbSOY
YpgXiMGPa4hl9V8Oe7cYR+JwewTP1p2LZ66JpxL/Mr9dbo33cTSNE4vHO4bIsarB
/BYUSyAAM68ojFoTULGYGZN8HxwOR7H5WiJnyjqIW6AUQNoYSgFvnmRQTyL+nrt0
EBid5/wIsqZSmYTXvaLKTg0CmOB4fcvZvzMwMmFUCuuQWWoT9LU5ya5/vTAZuhSx
ZsLzpN7MqZypkKewl6l8vL1SyQ+aeoOiEe1ZIKI674EeCgWkJJQh5U2LlarVgb10
6pJdBNDAH4XENiOn9JvpebO1Y24F3xbc0aiVcRpMoIb6Te3mzOl7AVKfVEsuJ41k
lenvdJJP85+LtXIfnFmnUaFUDs/BA8x2eTAExGbCkZ+2OFXPSAIQXWzhd8oIARTr
0KB8deU/jAaWejoa/H+vPZmuytUd3nnaFhqYyRqZawkmaPlWzi38odWJd6wV3ycW
DzAl3pzC2DHOwxYOUNM4eAGE2hJXhlnYXE4z/wWG0j1Di2EkS6dYpxa1gFHuX2MX
kwY6HVtTImBBoqiNN0Ghhpvv8VjJPshmkdIr2up1SvZ5/LnDCXaGuo56fBx45bsO
7F0b7OIaI5ifw2d9D7lSCejoojiU76ynTKx6L6gAOsxbXsj0an31eG3smxfn28fc
gQay9fEJuHm0n1DW5YF7Kn6po/z4nWnAUL9KG/MGFDlTE/TYA8ptq9uZ3NgkRqFu
/nGEDkU0C/vKsM+aCz3KJRX1AuAvddtlxEsd+WKx6NRqX189XJZ/2X+efBuVXVL1
o4dAkFwqSsXSAHfC5iVRX8jyfVPjwNyvHfMqKVMUDfytECXjWxTDtq6dGxGnk4cl
gmRVyRapLFPQH5px6VHp1XJSJtcBUFh4XPmd8Jl62zWc+ByRdiDznpjAmvsbo8hC
PRRxMo+KATMqpcJ42ZbXtyTaY1/0s8vRi9wPJNXGqMmJnubCFBR9JF6RHNYREMj/
dH1HAfUlYvWJgaDn519uJDXtfS6rjmBcAxEZc+SK/iYkMjROWnUOs1NNYvDm7giy
hKFVjrbPUpXUcntRSxkvJ/tQpqXw1L9Bik3ov96/q75TYGZk1aFsbsRwdAvfpWde
rjK6tRn8efX0eZ7QVGzL2cl1BhffxCHhjFQhLUxDfBkFj+d2pxvoa4x5oDuhq66C
xWlJzVdFQ73X3vjxunof6gPt9tj35aVPmbGbtg79lyuktfDt36iXOKkmwd2507xe
Q+kHubUlJqGMrPO0sLarrFr5KgkXIiLaUSSbmLyyKYKTxHTfeZnHWNWTPEC2Uyjw
sqUKLMLiXDq5/1HHHk1/xuFB/Z9erDJj7hLr20a1WYNIkseGL9kiVjaD7VkN0+wg
YXP2Mese9Ch0ozhjy3UIsNDR44lFwMIEFkD2gBx7W5zrI2oD+/7iRSzqeihCd8+Y
CrlD3ppdl0Fp6k7YLHi+FgcVqfYX87nvRTw04gXdlzLYAxqOzzgHrgQ9WQW29rIZ
EQAl4nKyjP9KR2EepxYF/3r2GBGESD0koGuVg/HIg+jkD/OL3LefsP1XZxpCQV9t
GvfJupzWpysJlSYfdWA2VoGsdbAgCRGUI6w0yJF7OU9Q4/u1+WenmaKxt0/6d/S6
weJzhChpeNPuGFMtk+02qJ5ve7pdy3CYtylqhiFCQxLtbUZZDLt6Gz5bip/8fyh6
xKtGfk9pEAdft4z9ET63rV2Y3xdn2sX0pMNFTYM4IenhEFiwDjuj1RuSBmYAXYDC
s6xi8julqzelENnNUIhEvOhmlezCrqICsWFb3bbCfoWj/gENtWEmfG1adTJXU09B
RWvWbPDrCXKj9RhW5ywyCwsd6xLW3uENDkw2RNQSy0hY/If2kUJ7jj6UevU7x/Ts
lwRmYClnO7RmhPQeqZT72nFjtMGu2vTMfWQ/1Dcn7L64t33WIq3d1hxehsvLBYUJ
hFI6jgCkmf0J3Ozs0q5kPBZO5lm7X8JXAdzjoRoW/5QKSbS60MK+PEa8yCmDyXhf
YjJl+M+r5mT0z6WmV42XoMwiHDQKL4bOMoQAzo6vEg5muS3p5iy5lcwGS89MlDtq
rDCD3msvAtDyBq5MORjP0y4Jzc21bdoGrRvG61mk9JNZlwWQOnvESmFrB2DIAzlz
QuUvvw0ezw9LCs19SKpVuPM41LqNjIw5V7lsnjkAqlB667iri+zmY+8lBzO1MGgq
C9B3sZDqX+Dc2bJa5E8MxICDU5HWqIOqiT+hQKVeCWEh2zplphMdQ5U/FNqa457/
r2Odqu2W7Kin5ixv1M2Uhl2yq7Mi53cXTq5KimKtUIp9Onps04iuyMJcSAoyx1b0
5qnK+oinOPslOoSkd7nli1VGclrLfZ9UE6BsuVEsxwnDVJY+2eFhMBy4c95ihtzB
P81PcO1fXy2XSj0aqt8nKpMGkOc7XAMIg08chKSHyUXtGuPoq47sWYjLaZA452oC
HZ+rSf2KA/pOhJcnGWibA4+UuT7i5XI/r09mWCjxAdSfe1mPpBcLYO0pY5ofUKV6
8QU7xJIzbXaYD5oIqYGuVBLdXyjooKWs+qDoYj62czSv7TQtX2zz1e9hYfcqC/l1
AhbSNFKSJABsZonZdGafxYxqe5Zp0QpBInp66plDZRBVKxQHaQ8eYlToBhen+UlH
6qpzhWk+KE8rwHbhHiBYg1P4FSr5IYpZIzP6eCFujowr9SD5Innb0jc+VUFu59WV
yc8mj3Z9nm2vbIb4uee2jJvDSfg+LMMx+Z9bc0Sorh4UHyVT+LUCIiMpkssesShc
fC2IlVClN/8hoDPL9CWWX2gnBw/puXhflYS5Ly4qIdiCKmpj7gXBqzgvmSdYeV2e
DWHCzMVNvXGofKrZ1Vt004d2DWOw9a6Qbfy5jvzPFsCekd3IXTuc/zlHzWZtt9ZU
VsxD4xzt1DZJ5v9ub39yycHlEYu54Wsv5plnNTeTabbHuirroy0LEBHBlS7UJroI
l+a698BWs/jdwW67EWfc8Yg7+6f3ROZUVuyPzrIlu9THiit3+rs8UecSoTjhyN5i
tCgExaF9p90D/e0sXxXLxopLV/REZgKXYZjOWBrIHkZavb+m9cavPImoPB81tNc7
hrI4NUIxJAwRtiE254m07LulR95EV3ZS3PNTtgT1A4IpzZyekKEgrWjOQGSoHug0
dXbqI7Dfh8mptdZguuJWTPAmixJTC3YrLkXNBHiMwy7Urg5OGcnKb8iIE4P5iu0T
R3pELulaTSNavlMnAXrRbh6XKuYJZHwMpfgynoCm2Y1qOjakcpHv0IiFWxlY6Lw5
+otUP20FmDXOe+zooLHmxiVmwUf7LirJhOLuZNUctWuHBcDCNmEvl+3xD9PaX1F0
RYQQTivfFToiPsVZsVZCHxFaBxBpA7J/u3SKrYXBIWW4K/Xm6AyxGqKmzj7OMJWE
AI8oFjDWGiws0RQ6fgcm3tFjJARQkbJBJnXlZ17OBtk0+eFnDOgEtN9LOYjP76BW
HX677qIDzsVdqBHMLJLz3MwZ4+M6BXbWbbRhtkfrCb49waOnOdSDGc6VSh9yfx8l
M47xo1O22ris5bOLHgx/VMM3Xu1kUlTkuDSLVVAh36/UJZEUfrwyQVHWJbrCn4SZ
ndWziA9KUr4e9cDCVllHBeZbLm5sfjpC2XqHesp1g1tUcOyRIh/oDUIQg/WNln5C
Yvu3b4cLQw1+QqAA0H+x4UNd+E3ZD+Mx3ZYXH1PEK99BMajwcN+nrTKe9T9Irm0b
nUXijEd7CWwdjx5rQYkM9Tof5vg3cX4Vt2PPk6Q3xHP26MZYMtGk+YqfeWipDQdD
hiYv1g7OqBN9xdXFlOmRkoiKa1PqF4CXG7Su6Mad06GQEBufSNRFiEkrRqHwQfZ6
inGzsu9yulUr71+lKa5YEtt98URbyZLXtG658X/wnrLkQrk7PTLn92HTdbY6i+uD
s1PoTfv7u09LGaclsxIYU2Mccfb2RuEcvGv6yIIkwO/jXgZj4b7JRqYtqzM2YY++
N8SViqCnJXfQadvRQzHEnirlYCugTO/2itIcbMLvsF51TXW4BnJUcZ9nHWibyCZ6
SsGWUR0TJCCpCJJndthclE5N+MZCUWSY2EnrEZFiYMZ/3625DjusmZ/9wlwuW7+S
Cu7deBmbbXG2wRFo9kTB4MnwFQswZcnf6+x92Ue+1b95lrZyDhMeWrpRP9HbvJdP
Q3x++0UxnTZL98XA/H3gV0/NcXta4CPYqEUQT2ITK6EkyRW4o/ntdKEufkBtkU+X
TfxhkKr4ydyxykbOGoI+KWa8zDiQTEYImDFWUbeSsFTbClDDNIS4SgDjyqpuclMJ
nJFYRLNmJRon0JLTHcYjtltkPk+11VakL+dKh6lr+IIq4D42I28m2kzfk5CLfWui
JoAv6ZHjup5eeRPqjL27LARU5CbR6UHs/A0VRtYbSrDOORaHmIFZ5wcqUKYp1WyA
JPBFJNmlw0Qcqomb6KTueVMCOaQBNBi0VA4LXVvJA3QeHqii9q2hZXPJtKdKS6xL
RTTbI503l/JCGyRMqLt67oDLYNu4760VdMglrQ6VTt573qEMTcjc0T9TkU98h62N
ZIvywNXiGewFfVvUCJHrLL4Xx5gt8bj7Wtdk2bC/O89127fA0FMa6FeHW87txZSF
OHy2BzMKZe1FI78eGEcnue06azA7JQgzu82pIbtlI6WomD7V2pUmvNtZgHfk+sQG
Fp7vjuMLYUISMiYB+iwvViKoGlvT5o3ZaeyczrB57BTaUnMVh1phIypXwSHl8Tim
0rdPgeuscK0qgiRFyRMDV9zqFHBZDLGYS5/mwv/PxKmHGlOvOwio8C9GfPfZx7VN
uJiMj5rysjyk/he3Z2OnJK4HA9QBcZ/DIZp6ZzHLr06fikyBYavYjoWgikVTXK6u
jyPejLSyvR/fP8LctUfa2oEO/MVCHWypPQYqLpPoTTdv1/V8LlQEqt5N5Akse8aJ
Wj6wIWqRy6YGYcRne6ndQbhF6pinsvsctzgqwqU2DPSMFAL/sI41wmuvkLn9tRwl
N6v5Vhu7Oh5GqqauU796o1ZESdf/cmSHhv1Nhg2MkndCE+XvhVYoug4Ue8epkAP4
aVsYkTvGXq6hIU8Oe4GTJF34tX485OdLn60DVocrNyZ8OppLFINL6JbbNQvNHWG4
bBc9b/UX4O+v63A5eQpHWYkbRJXLdAQnezdmdUSadHKmOvs7l4qjTJe3r0vnhqnN
QkFrwb/KpPhQA7Ut0N3MYA2vxQz0sn7lAfFuD9/DUBRmR2HVb9wLqIAf1YJpuZeK
Xz6iT6qPed3G9Vn78pEyv+ufsiKL3cHhWHfgxnWM16udu6GvxEwwe71VLuggIg7I
S6V96WBtdstJtztHfz7NxH69ZsakGbfY8wSNDbynYUYBtkMG2yHMfXqWT80dICvo
U1oT8pChxvlMq0tsOEqt9PjWrd9N8sDm6/fuvCB5qi9a2xSkY5/tWD6+8VaBuuzo
wFKeeBf/R4/kvZDfjdbbGdzzPgjQw7RjTS3AwyKhv8W+9SWOS22aj/DFTP5nPYOC
O/dDimuzgsCeJ+qcKQ+4JWamSQhy/Bvs8gT5bQoRX5L+EFeE31rQo+KfPhGgq5y5
U7INJSYrDGDZkh9f/Ji9ukJIfPe8Qjwmlt3ZHMzq7VQp66MDYPIFqtrJZPH3zAtB
FN9ZA9ZEJdKySvTzUxjoXqEO3+dDb4NAXdEsJHMo96jFA/tKEfhD/JgaOw2fPYXH
Am1yeCW0JceJK6t5nGpmwuB7kFuvNyNB6HUMUydFZkiQiRrvL67jXvTFlYkVwWai
P2igFTQt97twQP211EPs/+Lh4QgPohqPG3irhFuu6rsaCEzXIHjzvvVY53OPcTPR
/uiQIZCuIbNv8jOpqDqvFZsvyKusx8Vj3tQjvKFx4wddU0M1eVrhH1UWU4IEttfK
UJDK2djfI4HffmgBYZcXwfWVkv4qIF3q5ONGT4M7nsK5QDCwPYPbCJ1cDiLLDjN8
Q/3FQLWy3vxHcD8cKGsSUuYsMJXRzCi4G6KWfUjMPNmPfDCljyj2YeyShO0Dfmc1
ZnGQzZngbBm612ODH1mzz5TeJiosX6wPjon9goO9h0XnAUQWYUCrtuDHazEG4vo5
intASjIivLdcsXfxcJ+HM1jYu52ktYtsh4Earmh+XRfhNsEnZdCLDM2zJVuta98x
UeLT+z8iQFIBiewf0opQ6VcfU5dss20x7D++OctZd8dqzJVlvJ07mMEOIpUtvuWv
11hzV25FetNSlbdY/gpi9RAntCDp4Ui7vC2KDemXAHXFyp1k9bRTjZLXJDgfj0Oo
B2Ojs9z6NruQWViyWqRX7LIkIfzxRRlUWIWguts+cayZoCQG7+oQihoroAAIWdcD
PG7QB2xf8aYKtSNnc4rYCYfHqwkFPZwbihKZtBQdIeItLQVi30p4sOBBjHXtEk3E
grWkL8HUm0rrG6cGZWOEW4bpIfr7KwXiaNdGE4okIr9Ln6ygZbLARVw8l+0gU9UO
QOkQhr/yjcmJmoLcL4t7vbQTNBoMYbQm3KGMksfghG7J4XgEpukfq/LXxZDe7ZZc
BlBV5ssqPLJl9mOg7rEUxR9ZWpRRFXRtCedUxjZVIb67pNx+4Gtqgvd6b5RsOgzb
0QVgSuGTLU9c21a6hh7xjFJYh1kHWHW4Tny1VdB9sWe7itGfBC9enRgNjovwov+x
jUU787ufSnXQDOQ8xE907pA6Uwk652QGGQtDn9mZiT44G4pnGrrWEoOhK3mF+QOZ
ZVvVtGlIIXpbj9uHROgObBNoSAZQ/sqRFMFLsKUiPLZmNzLNqeQqaiTqZ5yo/SJl
2lmfWImPaxPtOGoGeGtB4QgxkO/+jQdQWnZt73TEEnqMz3YkZA+E38ZuJtAVz+jn
3zLcgTiverOJTKEZoH4fFaDdo9JxKQaRSOJle4qFsiU//PgQ/gOTIziVyTuR1Eez
Q+zh8Jd6priSxYzL9bQ56mYfiTNolzDt2wr7029W79N//JqKcmwzhIlMMoYmH5VN
KUU362JOtdICAtweLJI0/Y/tAuC+QTEDCT0Xt8AUUdpv4oWxrndg3m4N72KgeOKE
lRyryWNFDhG0K7L4tHEfPJtp0t4B+mmnhfccbcsNarY4pTvsog4cIX/7BjujDsa7
iR6Ll+l0r3UIxA0oILTpN4lENfVlXyZMJjulURax8GdUwUCNdjsC8VFNxEuV+i0V
e8iJ2rTQov1pZNRcC9VEN76TnrxL4U4/vNkoGdBBYTrM5QJSL3fGkfABLD+qRxQM
Hxzrco4/72VXd8Lo2SIJi1xgpSPZxjALLi/H50fP6KIr6QXZYJFiB62EOsdWHH1T
oU87SMWD98tKNm7WhntBxbwx3CK0PiG4RJgMApsEiUstDj7sA+4ltTTwihep53nU
+ni4mgKov0lh1atgNT2hTlwSFLV18+CL7VZyzVbScntnUeJvfQ0Srb7XfiJxLzWx
eYIH1onF7JCckuAxunDIdPwf0NQgWyZiDDSSnCyxzTxYadiajQidnP7uIj/+kOAr
ADmSV8wmdtKZhZnVHravUXlP5yvgLhDsaeiOKkmJQji/SSZCVtu8vchVebBA+07b
oAFREAzMQtfc1Vb23K7UDETYqi77//wfi5/HVJtbEvC7/88NChfMdQrFcu4BMqAU
bbjxr5OA7i/wY+DwBMUh2AU0nkxqzBnklW/LSpxDZVaL9ieT2rTFhNhcsFBm9A8E
oSXOW5CXPCZbP9qPNY9pHoplZ+Itt8wVX5TZ5uGQSk/hHWpuPPW3Jw+zHHDSrtIT
5ggidRcWxWwKY6xwRzaGxWbYDxiA4v+ETv256YyN8MMNDnpiT6oxkaXyxfGN9C9r
JWFEQY0W8A0U7Xz13ECi0spuQ6foFKq0WXaI67Qc029VbAhO6VQODh6U/yfG612G
vriPhabAFEKq5QD8Ok11hFB/LUmDCoPP96c0udOdGMlfh3/ikhkP5jf8SPt4kuHw
zOpEoaNNnJrrt1T/rMhqNopGgZpw4hfvcWWnknpEwkTqLkLV7vbWWwpft+wPouM1
6NAYJcgapr6NUW43+2YjvgnUKHFJKsemgUHqSpJIqlWe+VgY0+OQBzD43EbFmxD6
thIJpVdB2D+dlVDs2uLtefzYBDMqJZZmd3uIbVlN4mY9rXiyg1DkvwPQ3d3uEyCg
h+1yeBrBzWaEZZfJ1xpHjko6tZlboIhES/P9B2IGPV6Mr9MwTfmEsVqGUYIsbUEw
7mvxHcwUdsSyApUuynZzlCPGfiJxOOZZ+j807iYVbUIHd4SNnnfYDjywdtSIHtfb
5SUvYWMBMWb+HBTyJFb5BHxGZDaytJiWDLg5k00sQE3Jzn89vwtbl9Ac5/ImkX2O
EV1aVhTZzWX0803/fl1jHwv78+ZspZs9f+1VfT5jGDuATfNE7Zvy5oP5VU5YCGpV
QGK1Saxi2JaS2PErN1hxCQ+XymLAuB20CK784HQ2PS0tfq/dipk9HC8vH9FB53bH
MQGsrRXgIetCCd3CVI8VaJBTs8XSnfcLj3D9cqBGqsWJrCzloNTvS0xWA4ZLqzZy
FZEKPeXrv9hfIxTEN8esDsgmkj0vSaAmdqStLmwoJDq0w6GqEmyanyVUkL5e/2Sl
5TsjzEn3IATIxAeXRFzqGgyK+KPrGdf5MnUB9UIXCYLAbxcoC/Hg9H2nivWdZkuQ
wrXiAhR7p4+HFct5DnLRC7oEUl2ZECCSAT0TLCgsH4QTaNRSXyDwMaHYa/20iPJq
FJ4VygIsXg5Wqt0y4Sd4UjV8Sb9iYQ2aCPSpO0XAMYt6Yhqy7XmiBbE9g1fNorN5
XT8e53kFAeycL0qrSw/oj+8V30qpKkEScscOSD/VpqX5u/GY+HgqwCULzIXCEf8+
tjNgXn+Ya6u2paI5rVyC2xd2bNTJwHu/PPXG2zTgZWNs/+4KXibBQnx26gOirqW/
8jTkSy80W4SxWQG3MAN/LUeuWWk8LbQeY7wso8H2ZvhfeZqyE3TzseO7VITUHVLZ
IvVN2DQ4hwkQthV6OpoiSY3CFyS2lXcFL2cu9tfR+r4/Sp7zgUv2slzZxcVKTELf
MMcCPQoG0wqcbK8sA3nledvyHCUoKporMj5bES9yP5EHlHWnlWQNyIZeUJ1CFqH2
zj83mZwflLv2SLTv487isKqsUnm4zoo9r3YGC/jspGPd9JNSgwKJUhZBeBW7v3ax
yIJF/Sfex0oD/cneBKa5js292YNeEocwkD3ZYiD0R/UP43ZdnExDg/ouwyK4PECz
S0m9KOJDIGgWZXrRW7s9hh2Hn6UKRZ0IKGoK7nvEyy5ijrPx3YtKq8p3KGjpBk53
oTsPGkJLixT+widyXBP6PYTgEOi5h86QUpkxZugyAPnsOd9XDyc9Jd2P64VsAy+A
qtoB26KTkc4PcJD7iGnvhh8s5bfH8OurnOxhNebgdkLh50cNbCUAZmPhniF64UCs
H+1fmqfwatRC377jpPEpcrlc6a2L1bRYsD5RChqEif/IWGG6CyIip88oqUvRHsWg
/d628Sd8y8AcnzQVma9Gk2D1XNxauKLBKBixflM8SURPuWQxzQpm77LlIjUcVaBu
7PnqYC+6k7pvuiPoB9CBYmTJsPCYzOuDnLC9ZqjiI7IFKxDfU3HmIAWMBxE+3bJ/
e5T/mu44U1XYpjqPJ8bA/rjU5dAKOi0Yr0Suq+zsT2QT7bScqDtbhUddJaN2jIjP
o2ZVki10w8VkOdUElFxd1SNbIfQ+psP6yAlg/u8IX8qah8n3XSgrhnhkKPlxJCNs
a/Yw+Ioh1aWyhIm1HEIn2ZRbmTjD64kIHjd4OObXVbg382rqpuHTrHVPdmUy5x5B
hw/+plEOLsphztfxSYnqwSWFLR86wYcronYLkAya8HKs2G6nWpYsbwiAsxfWPq77
5ziFb0UDgGsKal2sGG0LALQW0VYLsCQo5bhg5uD6wzuJWQgzsjByNiL4vu8cQtnV
wxovWdPjM08JNksZgic3mPy0/j1wNuTQrL+Fd3xB9/vSHkTOYSqjGmr23eKerAJ9
mVgOsCHVxtf3zK7wei/XohuTRT/OdvEBlRCmGL7ITp3dquIpXi4G1FwTY3bs/hA2
D/zajWv06gahIsRb2G/3Ae4KT1L7K9OrqBEFfjhhRp9t4KlOdaReVs+vjrzo8DZF
lhXXb0yXLcITCNHCDGC+Szfz5jARA59yKiHh8c3LxJrdo+39a+AMRBSOz0EyW8FI
LcsPOQCvz1uU2klLrBhxbeWTyyuFjgAUFG+fzL7P5YPnUI068lOvJQRwtZC2DKWC
zkgBVkmaUs36AYCAjdTAkLbiZ35aBfMkrl9EcZjlKeAMfX74WMgsv237PhRXS7ny
el4d1AaLvfMSKYvy9t4IvY7lLAMBQarA2zMUjsC0ieyCRPVcsdRogjj2+ggDKkeS
DtFzdQEhpY5RbYRg02BJqoXrUpRsZjpM4tnYW06I+z2zyAvyFj2vPU333vwOXQys
kXGdiTxPY49SPNwo1xcmoM/48Dq54B3X++OtyI8MNW8/azOw9O/VowEH1BaLOGPT
dNG5SI/EDWL2Dbg2laferxwz4j/u2rjCsq3wRrz1gzdTZFgDDx6ytp/0QXNR8m8d
lchAgJnoVGrJvf4wPIeay8mD2C+CHyq4bv8EiN71dvw/+J1YaC+FjnaC5FH4UJ4k
2TZg2F5dRJEkMHzvbF5rG7Ar4sTFR3HhclBp20ivc7iNf2GdiVVKIBdw3mODlPV+
WHEH/dH9odZgxBYFcl2I9jkYXu6YBikutAhHXdBqS2ibIg6CUNs2G3DcTwEMIVae
uq8Q7kBuwQCCsu4ksGSbVxGnyKtZZKx665eeMELy7oHpBKPAoqPQGM3YjOBRrTWz
VLcg7J0E/vhC24On7zEoe6Al4qoEuWRYfCAIgnLtysIFq1jkyFkcWmFZWfdpC9vR
562dzH1w133XDykN6ANNCRkw1CNc3PArJWzfAZQOZkC9oYijbTZkjDT7ID9VEY2o
jCebz3nrnniJP3I1jNajsEDQtja+U77vklLKXeZ9P4rMvUAedCMYq3oLaGsIy4jm
sHXQniVHb/uxZtRweVjsJC+ojTd3SIQb4kdh24Ne+YwBbH8luDoCUlBDLDCGrvOB
b5paHu5VrNLzTLUpSPO2K5aq51HqoXz40XUoW82iJieabgYXUbxpUh1OtLiKILeY
LPNH9kWt/Kt8UPfWfF03Pl1+KPP+rOcHHxbNbd3m9YRw54eaA1WUzvNUy5bi+D20
gDhIcQ6rXWFKfDaoww8wIBS1ZUbnz3MSvLHXTxZAmlEHkb455hchbiKqNu0lh9zF
MCx3dycq814H4H/SXrNYM1Vsk7Q23EfVhnoEWqM7/j4AJAFdfT7MLxiZMzUTJwgj
WFTQNpFwK0yTu3SB/7uqLhgeuEPzEAXHltTuPZRjXis72I+nNE+KDltUtnUT6Xim
sGLSpVn4mN/brXQ9mzqX++ZqwRMGKOn/DF/3Lsg0OE1lp1lpAYgTa1LG1dpPQZt4
yNd5S6nhLg6UNT4ariID9QONWmMsv1uzUcxiQR010iA1TrmdDMvHjt64aM61vq22
9+gHChgKSTjrthUyGKKUWqjTNnyDVZvNVArqTuMiArrMYV2xPAKYG+Ns7jntNaRG
Kp1MqtYS560NJD5drySNEXNJjxpx4W2l3bVAboseWdYfjcS5doT7t0cbS8U0sSD4
SrzIioWKKmB0dUkWd4PguoDB1IW6L9mfqlDbmQJYqKJe9oYTZaO9RWj3zB0Ks+IP
VHGJWE7CVajiyY7LeRUUOYwpNiEw406o4LyrkYzk9NYKIkr2K2a0+dS3ob+Ol7lU
Q+c/ENMx2Ha0eRgiT1JousbUWcmwdRi/3JnMg5nNJn4WaC7H3rY1RizZJBSuInYc
IQaP3hA4qmwP/rvlyn+bQYH06ZuHkD6IEpvNeh9MpryiZ+7TT2v2qvbmCAod3rkN
9DlurYTZMaE5/HBKSiQMmiaYXRkvJQi02Ia9f8Og9azZhcRZjTOfSZZiKJdpoBHm
VZT2JH2Kww+Z8+2mzODV3MWBpg2uqQ+4nZ2HBiiZly18/ZVc/9T0DF9D6PX/TEfn
/BCAfPxwN3pqLFmSvULceDQeTkrAL9szTN/MKLVDFVq93OOzMhvvVDRB4nzXDbFf
3sV6f8e9y9zMwkDH++VrOzqjtOG0HdmJ283b/6Yop4z1zlzuNpVX+8cBK9p5zvYe
P+jEylB0qDwYO7YkYwX8ZyqzLK0yu68jXcIkUxz9T7BbzmhC43z0ak+dEJQd3PGm
9KpTiAMrVUPjRobUfxPP73txBLEYSwIFIuDVk2JtXErLWlq1/HLPluABwC7SXsZw
aOWu7kfcqW74SyF1iyJD1nilG+N86QfYLopwmIJkYC8F6yjnewwAbeGhWLez7bX9
y04/Do6xVMmqmbrE3NDzFnGL309Fq3zXMShakw9DcBkqDSo9KiQJVLTo3cVsqAq+
zDokd713SdTkX9XXOhUecMVmY7IDFuwkjDF+Or6ELKSzjamxzFiHKrZVsDgWNB0z
ZMomyd/09Xg7vzc0aeAEphz0812x4tZGxvRXMnW7p5DPnyEC+UxSBJfwILgc7Pdv
E38NLX4yHQjrEFNEOGUOByB5GMWr3fB2zFiGD1NpSdR9IOPeP2yGGTNZwWwWmsX7
pqatkZK8k6QvX9Tk6/vx1lfmM5/FsBAzEbnoGc+wApa5rXUq6FJnnX/2DiOBpI2G
hJErk/XSgKelvcc2Ye8L59FQSyUxR7AQSwGmiYkkLgFlbPwu1yt2MN4Yv+eYGKj9
2dl15CY8CM6mDheAZMnZbTXnpu0efPDALQ7lZl7SSPzC0nv0ReMXGP+h1kn2TlMz
AhEuOoJ0gnJsk25tOdqegSXj6hIM/ZePiEYIvS8yeiIxuw8z4KkrvXMbD0fbzfGk
z19jDRjP52dCwFZMj/Ha4+Uwz+MvkPyP3yVoaAfiLxCsnfu1YNZ7OO5s9eDItw4G
6IMk5oEAy32qFRDBpFDBwLMTS3z8orCU1jBou0I1xpQdPwF8ewycdPP2mi9quiSE
R4z9lh6pp3HW2Jq4JTj9oGiYHP7GN7oDIF9l4rfxUjta7f1YlQIvQ5cIa+piXVZe
dQeHctlrzrUM0lMC09cubYRXsNGdSMGvG0YfNg4utS8HyfZqoKQQOcZmTinSBzQY
gnu06hNv/QOc/B5K6DkhjEftfVsURSDMDS1PqeXR43fuW5gjHEcSPua1r58c4T6u
b03t6vXLuqlTfPErzjow5kX7Y0veNWlT6UpEaC4zEyPbDFTqQeqPy4cTaM1ZU1uL
K36KiiV9kuuu+hQh/ZqtZb3WG0u0wYI97HQUeWI6OIACyhDV4l5ceKAES6MzR1cR
tnvpEgCgwlvQWhSu54vT2O50LgVu3B/aSXu7OcXNnujcGrzDslU1q+TSafCW+QvE
yEeLfLT0MWVYoXZJM13gldAbTfogHbpYycnGsMVRIu4NARf84yVQ8HP5yk2nIL5k
KcJTosXU1fOd7CV3Ibhq8X/HHJAmgdkDiuPY/QZFGX//EEp/pXsLtG5DhwzALGq3
+Fg/zPq8oXGRKeQ++7DSAnj5NaKxtEC5nqCQIwcYUtzO5oJYnu7bBYHousAKojqO
cmuGS/ZFlH/whVXdDgeFVIfOdzVBunt6mg076WwGqPvIXDrxHJPApGcxaV7/k8+d
06tG6VCbiI38t4pDFMBucglIKFyPE1Za6DnTasifiVqwMBAtWBGAsfhB61HgF+aW
+GzYPpv0kTHL3zRcE3fPEqgZ0FpwR7GDM+xbQkeXGl15bQdkX8ARQUWAYXF+Mo5S
yj29YYs3yA9lo2dJ3L4j281X6G9EU0UD0C3iFossRw0RBEekWnikjymiqqL1HgZj
GQeahjlpYBHLKuEb2VcRQOEAha8Z7fMS8Azpo/Sxy7h34wLz3wrzCRgCpxh6nwMN
d+HzHndXHYSrRvitSOt2Kh8dUajLqX1XysavxAbNTWxuTW1DLrvfOrQuJfhgn9wi
Uk+nsgPTQP7yqruSlqi+hkmC6sHMH57tyUrtd7zuBoTniC75bNCuF5OQjiXz0oUB
JUski41XG6QwEMb2pmibHv5aDWXEeydlbbqa9PDu0UxP/riTsaEIiyUQM8xGD0Hj
7DLSZB2gLH6B/RtNMjyBHVg9F7Nkns7IRvGeud/tcBND+TSL3XMq3BsXo3zSmf8M
ft+kFhNiHL56RtyukSzagtG6sOhVNXkwt40Shg9fatYj4rp6Nm5IBM6F6hTKHeDd
UQ96+LONIcB9G+DyH5djonncneyqs99AMBn7OSMCI5l7IQrbm16C5yiPeFw4BcM5
Pjc8mBgzcioBE+CxrMKkfSpHEa6kzdLc38HqnSN8qw9RpjKfHXnqtUryDukbzlUK
/nC20OELh0WMy34wLNRIKO3hW7vFjIMjH+hMyM4yMTDExvNycPw/9FFPdYhUzARh
9fT1kRmw0hkDd/YUnv1orWjp3yv2GeFkYYKtF9YuybP5I2p8T5H48Txy1p3EQ0YL
O15wZcKrrIsveZ+gpMnz5Zcc6oOEq/D/eoGs44ZelY8t6Xh5Gb0u3WY82cHFZjmp
kuo9a+4DZdKkRaUkQXjLQImfqG7NmbcZfql4bJ+qG1B5Hn3XVZmNCLKFtL+NM5j3
1cEdTurCn4fHlEotaFDv0IYWxgrO0DflImj5zPhd5ywJ+Arx20/+e7UiltVWM4Sq
7QUnw4G4/8FtBbuxyFBTPsTr6VBwE8Hl66GNJsuwPONYQoBMA02E7cs/aTaHBmtv
S6RSKr7XZZ2DGJdgxApyZbXbeXcC3r/N5frZKNXoj3dAsU4c2Nhpl3POfx+cdksK
oJz5E8e7BN9uUiDSyE/WFVKzgnZd+VpzFdnJivCGQ4J+eR6ym2rkm8xlPY0wCSO2
nLC97cbBkkCyCaclEubtPzqQQvHihtgLpyHICjjX2HneyaSGttaevlEUxWs7Zc1v
kxyb6JeoQe5vH/R1Cx1oedMfc1Wb0LOZlXX9JRK+SEGo7NIFpU4o9F4DQiCO7S8c
Sm/glXDgM9hPoDxZ/yOxwRHsqwfOZpitzTDDrlsXzwLjGDScMrMWGXVh6JldDHqc
szE/UzJWHDkJ+RcRVsa3xL0gEs6p4PGmS1BQgoXd6sB0P5MuIsWJ38QoNaKOn4Vt
IwhOAhUvwr07+DWDrXI18Bf+yTptLNH2IC5F1MlBn/Gj+K/jUV9dWIVFezQ0mJeD
iGiEfUcj2ls0YHlRNpXlSrMNPxgnp7/H+CPxhfDS0jot9xxIzBMyvS79Kw22LM3B
9jNS14DT1mTUmwR0vDaJfJr7ldq5P3bd55adut8/SZ97eApZ93YwWVr+t8kbeGk7
jHLRQMisMZVKZRAumQhJD2bBRtYgqOlyHQLnzEnA5rC7WGOVfB6pfprYPGmTRKUv
mk1z4R8PkrjDuQea1A0YlujQySjdaOn6Tt5xmIn56TpbMzTEzjOoyNmitVzpVM8A
Y8Aur6eIONvB9/PNycH+Bi5MTpd0Eta79YLNKFaD9GUUEn+Ja2h+M0D13VtfUCDM
JtJ7VdyUVQL3iNWljPr13MnBRZvBcY7VhcqnqDwnDrCb+JnvjNJuDCqoLclhxzgO
uecoQeZI4iSpUmkelGjLbFTBQbJ517Oo7mMd1nl3YSxxyLZjrNeDfUP82yZRnprM
zXdNxFCC48Om/1mrW05O9iIVLkGP7DlA1m+N4U7Qi0kbjJ83u1c7qMhjeAcFftTI
3UTvuytDZ0rMBsVuTnsVUeF/XxZ+c3KIjtM2H3ilCcybeVbL6bVYeOJLSnBiAYjK
N3kP0/VASxXV8dx9KuCRc51rO/msCYt9CH33uzzPC61czviFv45731LYalp7Y3NE
j9hM1ln5O1OLeCmiVSSoReMcT2F6hjo3AObHHu5uUxkKFlmRnCtUqlQ14ZyxsYSe
tKqVKnk8oBvvgyD6zUkAzM/mhZkvGeYsj+CYH21nfo0M5w/9whVPWSq5KPGrjJ6z
3Wv9kEzVGUVgDs8unq4LKC4RTL8I+AcFQFyq+2C6TWdYRCcT8kq/k9yGA0tWXsjS
EDBdG8t6aNNtF6nM5go7bLAUGvZxxZ3hLKR2bCOTii7suSJ6WWx+jwJ8WJeaUnqs
GYHYS/5t4HFf6Yx4xbU6S1PeS+lNiOE5XYdNunyv8PLzkiEVYFjG47M9ygSGdwyG
9JSc8463mMdYWfbHZbt+QT+LliwucmV2jh8XyQQeFuJbb6wYigFQi/pEHs5Da8fp
p+dWw3pJdgJ90Mn2fv2IeOfghA8bzPI8N++gaJbt41N2eX4iD2x9qCp/mltJ/wIy
bz3u/9whej23C5e9vx1qVJzg6zJ702Ez/YnxV63squPi9dezDh0SpqSXhVBlA3on
P0g8kEIIax81xNcQEM02rFrhZOCknq28GnZugCJ7USiHgopy6ivOx7LSmXSLbkqV
odVtgsy0hN9I5zbsKZxSLfrWSgeRvO/BLjDHv9dkRMNJxMyvnsdudVTMKdBws45F
p8tTmcJ6ssLZTobMJ1J/WSgBH63MRb9toHfDeyPef48n6YZzcu0T1qIvl/m6njwX
mpoUNj/RWrx8fggDVbZxxaDHiZ4YcV+Ab1TeDKljH9bVnf+I7HZacLQuStnaqvO/
sin6XAKaCbbQUBp1G/xmG2HUFMGZFDQiXNeIG8EK7vk/7KpN5SoGX7qCyies16+Z
4G22hKFDv2jauhEz2Hdu2tCOQ/Gxmp5o+yiKMEROfkUq1xK7E30wNLHRopt9Iigw
mhfHJSASyg/YqqMabBjbWKzrmCYsBovJiBRCXJ2uBNOIlAwnhFVzfWyv2aWTp5H+
00dpq+4pqR1z7B9Z1ocxwozwhNiNkQXI1S2+nw7h/eLXXVLpgCDm65Ls43H6IX1w
0HOM+OMh73rF2O7UWyDsXIgYqkVWeUT1tNv008A7RJh5L937zzvduoMB40aUzf9a
9K1Cda4ajeM0pNTPkH7mrvBHCLGREwwg+Axw/NfVMM1/Vmnhi8ZbBLzfg/2jZVGG
3rE+Kj/iETYUZ651dWSCTiM7CaLITEexDCukLRADy5Q/z3smwbc9D3OjZ2erAdC2
t55sJgxoUIjXZC7iIOR/4LvI8E2gZMzVE5VqDkYoIdBRv9fSO2+IvdWVnZNbaPho
EzIXiDOdFYQYphNifODtg/n20A5xRJlzNSCCRddK5MYHH1NdRPlo55+BHDLkBcBw
kRC/PiLjtQ8qBrgx4GolGDUhpuQcBrvth62y08gFqklBXHWNOfVXFScb4GdqraxY
LQlGhbjnJFNIKWmkP4cD3LNIYsmsWtNv0Y+0Ue6Kyj1LQ/XE1JgUWRUdW76M6Mj/
tvl73Syu2AX2ThAhwX88JFJmckwYLxEp362yJ1Aqyg/SJ+gd5lTLMBtnbP0bOea5
kXGFB3J0BJvc/fKKIwUxSXgw5L3IiT2jxFiiJB48ohd2BDy6KcSDrKHI93lDMK0R
oqo8gXzNyCgcDMCC3o3xlOep/L+YvXENeFORiaTlbYRJQZMjnHZnCFTVdV5iqzoO
qHbnLl51EW2otO19Q0cA4Msq/HKIZM353ysXrYmIvJnNPyBB5Eq4uyi8gXHQpREu
uEY3Fd1i7hFGoyAG7Sbt5fuoJDhSUmrwrYQBfg+Ui9FB+qwEK6Mso2ZaqWfnlDMP
+qtV1W98svMN+S2v0oy6euMIDeOISAnLh5WvSI6vuCJO3zXSlBU6gHdDPSqyMQs5
g6EEqZDgSfU49zQuGOwnLf5FhuKU80O1mhaB9X8pplg2pO9OFRVMkYhUTgeSOMq5
9yi9v944a9zhoUDkGaX5FOfeP0CXP1S7wQu+pARTu5C6oZVyZXOlCQKz3k2+zTCw
g3vVSll+7kWLzh3FiWE0kU1yOuP9fh3SZmi89jSiWGo+KB6/Dbu3MAfzUsw5Z53q
Gy3gJdSqaRwrEob+iPcHohuZ3fnqJlN6AJVF1pFDJElLYouZaqR68gYFwQ7WXYzS
tZGMTLdA+7HfHLi/U7lIY/R2sf1UxSppmOw/+qMbKjFVb2vMctczs1cZzukzA8uW
MPpCw9SKD7XZA4UZJxfXBCOsEdNTBVH1T4iyNQEUmZ0EMPwamodRge4G5483JoLr
DIgu+YhoBBbhSgx8Mw5gdlSsgJ7UE//ok7qLVYwkG6ep2oncJJfS8rYZURKyhrYv
59SnvnrXL9KLPTjy2j7VhnV3TEZUCN/ciSNcr0+DMQQ7DIVH4nrVL5KBik999CPn
J4jLnWbQAgjxyxyzAOmaGq0YXY8EayzsSeLnMwuroy3og30a9pRqH23WjKyjGRFC
1MVWVlW2wp0KMFXcxJZ8BlDozGjoXK4OdlaMse2uVjEE13rUHOo8WiuWffMVKXpa
TPCYe7Q7zbuY/iE1YYSUjFjdjZv0Uxrl1j3gcA/HsvYrwD1mh2WZzcu57afMYISa
AlhLjiHGWFQMULmCFDj/5v1Xef4DmQpvIGyrGYN1+5ONCNvzF8awyMQyBOzQJh11
jRJsg0S1/2SJa8fv7N1qX56XXVm4ySOe9nhi2pOAZcMITi4rOcsILnuX+OcI4KvJ
G4qOWQrq06+lTMTrZSpdjdEh1Vfu8TVbGqQgrd1my801j6iFAN8uhyU66DLo/5We
F39cKmcTD0kCsNIuyAJyaRrtsEWmqpIkhehmLnhT0vkcBMT/bdjb5XjJYAN+MsiE
hhpXnbaaJ+na3FRtaFI/SVpaAqvOsIGJ3Q0CUgviLtoFhrRp+Yq/aOksqo5d36/n
ugapRwiuba/SwBiqS+pZyIAoBQiCheEJsZj5Ao1G+LXIItTHegfY5VQq+Vc38709
2NWrN4b/l2P9uJl64iQAFQWzvD19YkEHyacF/s3hDH0Y1kxDIAb4uR6j3dwXy90c
mkvls4OPnJEi61dd7nKp6wVgcHg0MXFvJk7ovTryB5iiykhKkdTB8UWPxKWFQJj3
X1WEAICU+B0joIWpFrGzPoNj0FBPBBDH6BAlNuuyVLu/XMsRI0EvMZ3ibKq1lPLU
eajtWupevB3RQvJG/9LEZ1da/J+TKOWTkI0NG66xI9cr3cDTsvc3IUYnTolfv9v5
cXiEE/Y70HzQuV5fcNsENqZOfSlw8emNObno+FZyZoGP/UQG8XbGau5UjavloFP8
zSdHbIoBxeCZHHLdXFIOhnzGQRescrL02NdqQG2Myi5lS/woGUYArTxZyu9rrt7G
khDFuw8TIucJdWGkNqM6eKx66nsRyCEqKtPsYagkfYMlHxT2cnFk+qy8Mm3nFGie
BbHH+mYF2dUb9alieGHtsn+d98Le8mhO76Yjv3DPFxm9nIOTh6X3Burjz7pixBYP
g7A1i+a5gzQozPC5lRAolLpSnVfsjAXFAxWYl4idf31wziM6xfXIN8K78KDzB/+e
aB4kZoxdO7XWeBQmDtuxpUbNHLNzXBzmuBoBopD2Uzlp4kiRS55UJaR2dDYZTc2K
NubruqNE8x1385XcLcbcdUXBTHm6/PVgSolBmaXShp8dZ08flNvSsNPdzkxs7hC1
3w+nDejqan7yJmaAeDGiSxBgTYQFeVRbt+uUasTxYSdGzY5KbSbbCeW4c6PFNi4c
Xq3sDU7aX/PxCgFweoWtzgukktU+kAmmtbZBDSm4R0FFrvL5MyeIxcwvL2d1yVTl
O3LTvITHYkX503IBkzeW8vg1GZMdqDwYSO9/leQi2lPo/zeZHxEhtU9Hcgm+stqX
tNHqkv1CUc86Sljf31R/RqLTfH+z79wLTqP4ofP22K0x79v8FVQx6tRhIfXb50ro
4x1lhUFjis8rvSOyXxwQ4i4SDg38NvUmcz2vlQl9p2eFiyE6taWT21gKfCbYrSFo
E+2Ba2aQ10YrZghMJd8JTmZ9y3Mum1LqM0nB4mdZldMkq12VQF5xpFRr5uM5fUZ8
5LsZhGLjNBRGk36YcELBpDQaYFX7w4OSYrGPVXz8fXOxDhbHNA1SC/wNA9ejvUQu
cCekLV/3NbGoPaKV8T5kED8rBQDsLPmFYanVvSxPiJ/yQftWQh9sQeOAZ6hMpVAB
KUk5FBMYH0MRYhqsqJRTBO+b2bkiunRUFLAowxD2FZhRhwdHX+gMq0wrLH3Nicdn
5NXyV9moI++86n35EjroIs0xBnM4saNpG2SqojfKHpHcy1he4x3+A4yW9NkNutHz
SGlrrLFjjENK4niVT2jnACd4xuj2lRRhfHZRDyKNdnpXTbhnvSl49KLfZpimyNjZ
uh5Ycgyeg1ExDtRPcHSSOpDAXJWIjSDE1G6is12EvyLY9nu3hqWWQ/IAOg6P6/gm
wbwnLA4M6TD6NPP3STFLTKai0rLURC+LXKnA5Tzznjdtyk+JBFmZ7sGrh3c1uMiv
t3ZZV5ZHu/3+3QJF97UHfkyucSWGMfBA+BKfNysmTauVV2OZI+B6ug3RS5aYWZPu
JCciOcq/8jdO+c024bmeWO7MqRwkJ6tXK/hdfUFM8OwCBZe5urnBTCsEebfmSKXU
FnNPAukyUMU3P4py1k43WMdsUxcWxtuq9ecWxanGZUNNDMQ+W3YAED2flpdlzmhm
V23UNPsLZxAr31ClL09OXwYAs739kKVpt+tjwrNMSrsxOtDECOKJbl6fFJ3cyNGP
R2rC3jY1zmJN/eAG3cW1LkQ+zk8iZzCZuFkRMJqv3fzUi9lqlmWl+FQ2Sm2bjGJP
XApn81xmQIEVqM3lObtG3uw7gXB8lvyOM2RB7X1ZO0oSbhhWxjt/4YSOsFq7+yLU
ZCpb43pwuj4swjHmS4NNrwa0gwAQKWuFdKDEZVU9BPUQbxTWITMDAOBXa3VFdyoy
5lUFWQ6y2mJojRHSiatAokyWpPQgj5FqpVxThKg0UdyNLMpFt1NyuvzNo3ftgGc4
u2m3iHpoSf6zryouFj5BjbneV/ipGnxqY96vcyHFQR5tz6C3jMgfCJRyjFaJVsy+
c586qeiT+CrUs3lG+UmaJUOZZu4fWApt0JLeZPxIqI5rItScriBR3FgTnxAeYsvH
THWkWwcXAhmayE5mx1MQa8pdHRCtAMp1rzMaXroVzy7LZFTkqfWlC1IbxDO+QBsS
alSZEzFcDlOIjMlrbRbZ7IxCW4bR04W/rj4JCL2+wGf+t98ifFA4XerFatWrTgVJ
iPYS907E9R1Pj4SkZan4MUPvZkKZW83kNVJQ2WF17EeRU9QF6i/6sFCBPW3T8PVo
iK6OUiA5ATtUDoQ3rDoucsaM2G7QK/9uElbnLhlX/ruz0NuG4fEDzlE48G9gKCig
zoZp6TOABLhWWJ2Cd7v8Ay8WprzqMbOqEwA6fD9fb8eH+uE373El3RFN4HQsZJRG
DjTmWZdowSOl6XjiDdhr07rjPpYzjhhzC9RGV9iLHt7edX8QkUoO/ChYFsr4DxNI
ibG6prrHEB1q7QCdkXvV3z5FnlyRRf98KImmH4gR5xvnAEeGGk2JBPsu56n/s+Sl
iw81TDzXfmMaPttDgfArPxvMWQ6CnQ2P5FUNsP3tI+j05i+LTkvlFaOsWo8G5G6Z
gpbACQ2KsLc6y28BnJWF5CGGxTpXimWnMlzK78RV8EL4xOG+lnv+TpXl+k2V/BqJ
XTrgR7uapa2RFJYjwgZFLl64DNNoFkhE/emBtZIXTNGua+siLbx3aIQiwsRLgKbD
riZlvdE2grA9Hurark2hGYtgUOSijqAeIhuZWMltwabLF8j84QOpKLnr60YQSpFn
A0C0I202I6sEjFwYxO+F5yKGxJrOaxpgMy0HS4T6pUFwqjx72XnPZfW97A9QAFiS
SdoyLXk01vmCrsz3fCwYJa8fdiyvvyEZI/Pi7An0+qn7481YpDbjmCDV58dLggSt
tEN341CIC9wiCU9Aqyh//rpZV0NbeersFcO3q4Xav48icac3wtWUK5Cf7ead1CEA
J5QkSrul0LmHLjJP2oIvm7OLwtcIFpXBCk8v2cp6tYMLv6/FsyuUQzSFL3TuRfv9
bP5ASG1Ojjpts0RZBTm3DMhYvdhiNZJbLIrIDCfuiHyI821GOhMG2/NlpRMR1riX
XucOmtC/ZnS4oRhp8/cJbpj9oXjOdU2hv3LIoPbJEqtCJjwkHNc1KKdH1QTRHiM1
50gMaYs+YXO9wBQ4kN3VpHHeQnr68hf3b+iTEjuU1829iGETR4bvS359IlsYxtK/
JTmRMbQovyIf4LLWL0dgAtXWXZ0b/ZQWJDi3s2wWZtQp/UQe3tT3hqZ2kQ9Hq5bL
uwnvhDAeuHIbixtIoZ8M/a2K7ly52Vln6W9j9beR/Ri3lxrcfjUjWE39hBWAMzry
U17ZcAbI+3zltXcts5p8Ft6hC4gVeiSleKWlGGd9aeC6D5xacPyrkyI7uqO7qs5A
nP5EBYpJ5eKdDcgh/mDRAKcy81JuamiSIZu66TVIYlxVfgkEiLnsM4eLAYK5uspu
lCsumjYF8dIvzmYrSJjXhwXPIDKSzyusqKt1xy5WidmaxPkBH6NsghrrlMub1N6y
qe9Y7ko1kYw7BBXblC0r/8mTL9OFSK3sMW8KDhfGgmvCrVUFdXK9Sk3slOPgOEMe
lk+RbFBPnHe4obO3FguZ3T7JqH0/+2+1dCd2wDw0U38u6hifJIFEmzQinVOfpMfJ
iynfPERGfBIRb4r/XjzWKCgtsBQfpP8igYJgZfxXr1tBJioIhwi7oa74RgAz+zDu
68xF8cd+cDRjL6aPOGmtphG/l7hxFv5mF3L2xaayCyCSCE1rlvTz1aWwiJ03gfw7
FmpH37WK/wyantwTRsX6HUpzBCn4sfndB4EnqgaP9M/HwbfGOFL1gzAnT0c0uccS
0QqRwghELgNK3DlTSSSBDobwdWf5u9Bw1Klf9XA3nZU/zimwkk5f9YLuIvgNMqko
Pm5NW7m314gH9ggkWmrWe2fD399Rec16J3y2O0UoOf2D7iDr32cHh2HPOJ+8iA8N
5aE/IpHmIPciBD1tTnPEe3PndMnO0EU9voFr3FzR77f5+9qMyxVifQxFKzr/XmSV
TH2ZihjrrySDfjXFfWizMTJp+//3NRNUh5TPthyQguyofBZoP2Ioa7qL4ZFu6U2H
R5FsiKufeZm44qZLJEfAHy2bASI81epgykoEi7bZ1XnVRIzOImWIkKYlBLq/M/X/
vGYCN7YQZL/CQixPTdtB2DEMh24SgbZpoK9SeQbpFq42ipwJcEi5fIysmM+q1MZb
spBkSKttu76/kF5l5ctaDltY2yLmQoSKeBHpk4KcMcjCf1nm7ToGhXCcMgesRaSS
SnkTynEzKSbYG7ucq7aurOneJcZzlpImik6Q305PPc5JWcgkIEmH97t4BZidsAEY
U3//6XZ9pN1YxJOQRR+uve2pCrYrKuYJCR3ZunIfctOZ/u24EyWJL7xnrZzDbqYf
j21zgIHQSGVRF7VougkvK8PIUWP7GjDKA6LuwUhFbQ9cehojWF20LbZHKT48Qpym
Jt94JcAziZTUCSt3acguV8+aDJK37ftA1u8KfvZxNttX1f/BZKmxtr795TX1WEsW
rzU3ZbNTskJh6EVqu2r1MVQix47IPvtyBabZOruVUePT8i7uQVlgqZj2MVm23IYm
gblJyU2ZpDuUNFtt5PrgpioK87CnU0pvcPzpRU7q7j6TRxGqieRsycvT/spKq//o
QTiit12Ac+uSrFp5FpJ/VCF0dmcWITKkWqCiIQqGrhr9XQWOy96ArF4x5b/eRLeN
zReU5w65NEmvbvY6j8dl6ybiZREr1Nb4gXETwBS2b4NWwha8ReJA8DVesewarK+4
7vFHFaf2iWu639jI7H67ZeaSLhsxua86Idt06Kutxp2NW1xGHuFdCdnfMBpq9Nfh
4exbYRua5OlQIB5evYfUffsGNiA8ytTOv/oEl+t9uY45xI+k+uz1x+H3QLUH8zLl
xiZfh6nUvTMlpzFmg+xXMp34hm3M/OwLEmABH4IBN/ZDNXXiafzIq7B6Wk2VH6uD
kY3GRPOsxu4pgQE5yKBvGerPN3JbVtra2j4edhLTqk48yZN5d1lNnLZP7ucXkv7/
8Om3XOt+eyzteNH88VwpimDi+1kCD1FBkIpyBzSrZnbD4terfaq685V8J0PdMoP8
`pragma protect end_protected
