// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:01 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YdLFH88eVW1cIdLI455uKw8rPm4FZ/DRQ7Y240yGDU+LavKSWKr6FQ6ynOkMUhx6
uct2SdzSmummbSMBMkHngq4l6VNrIT18Zjx79FA69tsLLBHUPvjhT2pYcNwa6m87
98PoZ9Zhd2IOCz1WM1WIB9g4G515Hv9GACddcu2Q56M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21952)
QmUDVRR/Xq3+g7wX14J8xAkTKnYpRDEIOnjA4o0rRofgXfrV7PERDz5MKhmGamrU
v4QrgxBoeghp4TnTpqMqcXjUuRtj0bIzW79YHWPd4i9KR6rk42ImGAIE/tMs3s8/
m4Svk4nIoTRMwW5UocQlFBzg2+dkpk642FottBhyCqXQxWTU0JrsnAvJuwqZvDV5
M1JDc2Y4XOZ+VR3kjLzISW3nh/Rm0pPnFh+7Uu75giTOI1cOXR+tKAhlHDagkL4H
elyETjOa7hquw+qDaxUrAFM9UTDesDn2o/NZ0IM38WP42Q9b2ynHqJ8/Vo1vxucu
mhOlYxwnzEck5RdOZhvSnP9BR1Ic5KO51r2SP8qjltgcY13IP3jUai/gG86B7Uz7
ijHi7Oe8DnrGR9bWElpO4xFAOwzzQYFTEQTsBVkNrR64SQpTLZLhFAd5hM9eLoht
DrGQs66PpV48ERlZ+hdv1tbje01OIcelqFd5Q/Yl+1rCGF+fGckuszdSg3ha95hh
5MOZ9xcDhNFJl3zFd6YHQkSrp6kYyGViaMncQurtQPMy10I0X1JEOIY7bAFihBEM
F92Aiv6Po/8PM5EouCdqN8C/WkYBKa+SnuktALrh3qO1W6ngEk18d2gi4rhQdTkS
2NBY38qEvO3UiDpq2QYsm8wOfH+vRnrKiwLEJm5EXzZcfSFYzx+I3pBaDbktNVUa
SkYMvevpSuHQ4vXaNOurOTz78w/nzoiqpKpqXcuFFRva7JBkB2PNtRotdtz/Boqb
3M1qhX3l6xpAXxg2Fp/5zRzy6x/tbQkgSKC8Wy+0raDzuKKgebvOnyvFOTy+MMsM
49iYBdP5HnutncUFZzgXLxKXDlIdPvSMcjjAia6AAQhldSrfnCYNzhddI+SdMLut
YJdw6Ax9LZndVMjXI9aS2TR0Dqsif6G3ekyo1snrmR3CxuMvsInXSDcwJD4wM0f8
ooimRcUl81O4bqf8uYyqTt58SVSBwSufz/aRvMtvUAi3CbYDvErTzvanPE2Vnay1
37eYXEm9AupX8zas1IvpRYkl0en1FofaLz0k0YSe7bBUP2rGZlacETUDgLUAg5HJ
iM6sAVFedY3DRZvJUn3AZsxC4DvGjzJ4rqMysN/gvYGVqBSPbrkkHzJdmlfskGPi
YBI1e6HYu3sV7x+XlC/Aqgn7FmmVbCRQWkXYy5Zxm82mhvKynV0PxTwT10g792Vp
g9TAfl+c8q4GQvuGwRmyc2V4kGjLJdNB1TpCS7UEpdadmqAKBDOXZAaeuT22MQ2r
XJM/lbHrrZlAVcRjzTxuIR4Vvgu48hFZtybay8HXzuh+HiXfiM5F7wSTmUsgr0YA
uK94YCa3pyC/2TR/WMje9jWVFfZA4//LEn1r/l7/QO3PLoVblHcTXc5pomhuMfYn
OmFOwlmQKHSknARJqSnnc4LBX4PeqOkdKzCBOta5VI19Ha4qpjj3YdJ+SYtAF6oj
igEjJPjazx5rTUfoZvcje1ZuMRW8Ph1hOrbKK0O2Dqoft7LFlhmLsJ4Ot0Vb2y2v
/IATyFAbWtDDXzr7b8D0F1QYs/B+/7tSixTk+TeLdsXoJegTtOBQMcoW9AdHt48n
lhZO3YOQ3JSqWYZGhsbPazTazdEkCSS3cD5SdjbKdgJNy1RI6qsGvIMbK+btOAjL
e3JsbzJhfvT+VFgtoE06KjfYfFeDFArDGl1N0NciBKm6TXCrEiMa3mZohi181EUs
SPFk3IYVyYb3gI4fGpsavuFJL08tDk7kV04E9tao5Vcik49feWSQ3H458OilPRVP
Hd7hcCFAC0kmp57LBKzLbDQiWFwtUPTkmj7FAhy4c9PqmlKfupIPLXy1oLWKzctK
Uep5ewHWN26QDbnfBxRhfXPT98hRgtfpiBgJglDR4iWc391NhE1Co2lY9IiXYhrI
xbjyBZ2ItCCYRJiOq7y3BVs4aIGosMKAi+r6T56JcV9cdz0A7sYKhaH1KwoOdBgD
py0cotUc3/zSczH/GdkKdJ+lBJF1Avak3vYRx6iMYYNxa5FXCRssh515GIgN4nx5
ZHyVJy9jKYEvgkfxB9ZVdyRcUmbGoASae6FjRGHX4ffap5BZJBXoh1IaHWfMkRxx
Q3inLMsKwR9Tl/TxCy17UCundcVsOI/DQIBuMlLq7KVO9z7XnrU75tDEX4/SMKTL
02aP/LWQm2iEFdGHhONV82Lm7mZWFNZdNBeYuxABmVFP7j2YZs2qnVaakWf5a9v5
UkdOPMcS2X7NgXRArrwyVQ36wGk/xSV7WYkPlJRuxOioy8mIJg2vuP/eHV1wZY5u
ZWxCRPEdp5FSc/5tB4aUBakiFvaGqmk4X3/f87DUI/tgyoQ1bW6r1RpvcTpc7N6I
kWz6kaIUqokzfzYnXaF2B5iv+sJEKEvRrKdyn0XI+Jq+/ZCSmf4/KAjx4p70kAar
VgNBAn7Bta9Iofdbzk3XaPyRgXyMc5L4kQtRiqftnIqFLdjezieBVQSjLZL/MGXL
sYdaGVLs9I9MuQCVDjgyjBWJ0d+uuhTkkTJyxmAU5IUvPeWsnyr6oCe2JPMDLBAK
9kT8MPZvllSLXB3SarwBqW+oviaEXXLNPVUXqJRPmoQu+qVbEprpCROoPlGlByvB
IUWoXYA+duKAhSUMY/yp8HcABO31ZkCP6Z2lPs9S5caAmBJonm46CmCxQ/MDyd22
sk7i0Ih5ERSUW3gTqBUfbXA91Ft8mnujCad5X/0NnRShrLPX4L4aXiGNXYz3ocbr
hiXmbduQRhOpfpl+Gvc/MQks8qpRuG0fkODDSEjCElE74aUmqQRod2fA3Lra+SI2
SFHVyi6ntMIHGGqoeR+XI8Xx3UZ/+wZbG4mLE+NKl+XAIXYVMZlnYjb0oJ9O33QO
u9iwJtwJ1EJBhMMEtO0EdjTIIZoK2wFcpfgwwa5MFBh3Wn8PDOFG/b4JAwBYq/kC
KozdQ/aGCf1SgmqMDglCLexEhoXqvBIK56TdTluQ8q7yh5Suq3NJxTOFTgC+sZcf
OYBplmOEqHKg3FHGZiJE5L/RJ3GWjXI6N50l3mmDpqnXrpZVj9hAGqsIAxO6gAil
PoU+9pBifTTz+88j7yei1FyF6BgtM9jY5cioP9AHuSyOCjoZsKkXIbDMNmukybDn
Fh6FNTeRusJ9rnFewFexnGGGjZg8j7FemJ1oaVb7QaaCLV8DSbAD+MS4VAcIVmOa
KrsWkSg8NEclI8RGvRCFBq28AJ2kE1R0v3A0SR60oOeWZ1iyOqWPIODP8gdGotYY
YvRo8C2m2RjXAc7yMWLbHO5f8F6ydnWC0c8Up11EOSGCjc6vb5zZZhDqIeutUqez
wP0vcKEFtQ215veransln7X7T07ezg3ssGeOuz1+oxAH1traEdCeR0LqrvWmKMFr
xAQL++sKTsq7PSxRj1ZGQdo8ZITYkLXVjp+igQvdxR7fgP8jVBKyvN4tJRZBYDWQ
4Odl0SgqXqoKPRFy8JRtgopHzhZdPZ9Mf+Ov0w/oZ4q7zwJYpk4d3ONt4Ry3buOU
EKO9sSN8E+79O86mv0JyTs7097277ecH+Adb+g4577eyxlmeUYAjpT4xrJe2x6c5
mHQqKRderrPRVZkbNLWZs2E4MPyA9+au2oeGqwN5ohy+n3i8qnJnnh14JoPHJvHO
x65svw+DLnItQqw1PXKIEy4xYkFVRVWYbJp3wDuoTDDQZ5B/YQpN1UPp/StJfF9H
pb1zX2RL5ceI3lse3DsYt9AHT5lem9J/G9NM7HJ9pYxYt4JzSCpGPj/h1et+Sj5v
lpCTL1idGKBi+2+vhYSpJJeiRgmNE0wR15Ttf8JoSzUcRLuSSsOGxpJD7aXzQRco
0c8twVwS0luzvgBkyXm/XDB7aYqwlOsJ0Pod1SSZslnmlsso8xKVr/PwkLQuEg5N
kBRFU44u8ZuMmgBH3fxtWZQwWTyAuqZnN1Ws2tj5F98rBpE8tm+eVweostlI5/Vl
wVECUxl+GbrVGpjg+BxWMuQLv8s6ZrRPgJQVuXtl9Z/vF/S2BHAg6BpUWD7JP2XS
/n0CNTErQkJl0xP3oK+snV7pYOJ2Moqefd77ALAnTHgvZWJtALPzAxbVNV1jnf3j
E2fr+5uvMT+y07wnx0n5DHz4PAalvVP5VqfHRK7KhsJheMwj/5LtqASiVp5zXSQP
xkHcVtJ3vtfd9I/SBgLUwW0mSazJsNqTKKtI3cFdHXui8NGCgWKwXdreZnQ8l25q
uUBwqrbXtWc6W0cHXZ4DgJFH+sDN6yAIFfmNCs0hnqTDSsOLrBN5SNcuvCAY1GGT
Wr5tibWXi0vLTVZkE3XxGpMWPv+VHWkKERIn7zSIw92eBBh3fjgS4CqPykIvaO3/
YpEsnVdJybnJ+a7Uy5oy9onP0DaxhGmqoiVHwmpofpX1lYNGESJXYa4nyqC5Ot7c
oE0rwk68i40ZlbVAx7i3M/Dmx2lMbLhLiPO6iIz88ZyPBxOcazMpKvIv1ZPXrRn+
6LcDnLtw4ZeOjXaCjnpaDHFbJBriGr0yUpUp3IniWhwNf6QzbBZRe2XsO8r573bd
WJx4PNMNXkgaiJ8RtCZofbqWygGXu5w+KqjfZZMQLbEYEtHsrTCVYtREHcctyxC8
s5BpSECIclOHFXgym8om97AqZTnG5uAlMB16/j9QIzqbvCCW+N6tn77y+dR4M2T7
fs7XcksoK4Qlq8Gvm6dmG2PmTAdrX7lkayHFkUsYTbOqQRoiXsslGa5QMPODarq5
UUg6PvxdNZ9H3hfasEnGOBMsBv82y4alWnF//A5+CON/1mH3qTmOrCpvbHkClDJ8
/DZID52XBAQG+yZry4ht0xOkRFzVoJkHUemNuFjvhFT8/Bq+8rwMei/kT9Wez7vE
GdUdmABype9eyScEnq9446rdpQVb4/riqwb8BNO0CV5uQZ+yVFWpNsG4J/UYvFCK
3ogRu5wB1X15YxnYFiVsDKKx/dbYcoWEJfEmE2Ypj9MND/3TnJf5RJqNH2isTCOT
t879tm3pqvVQdXcnfV1n+pS8bVr08j2CU9XmpGJ5FbEqmS8gGEphNViMEjE2ty0Q
wsy/xPLmbO8dfe+8V/T0D/b99bTNQuzCsFupytYYKpG0DeuoDP33eDeKQebEy0N/
9fiDTrT6o/IX2IPfp0Arm8Ak5VfvwlzLojPomO6MqWu12ZJK34w7qWhFaFMDTRAz
HIR8MxlQWivrCJiCO6lqDbz0xGr1RPrlKiGzucGHH+QTqjYEJSs4JkPC6tztLwR0
U1B4JBdrzvpo9Yc2iWBYnFl3Q+6akwxDcOFN9W5RvVTWN+NEOVaF1BDCTj4gtNnx
e7/C5lTOSzvodZ6d3UgXD8DXvqE1rdLUqIXb96B3pmdTX5aaWgw/xfgk3z3ehT75
W/HT1N1k5hfOtUw4HfaWu0CVXAPF2WNAyBEbuIpxUHRfW2c0RAoAJ21OmBVl7bWd
rkCGr8zUffHhItnYmmXdNkgRVY1M2Mta0k2pftB5MobcRVrVlrxEkqo1CO4nSvaX
CsVmpuNr4ZETWEYZILb2AtQ7MIssEzhkKsrkSl1Rt3Vu3x8jKONnncmpm34o1CxY
272BUm3ggS3oLo3q3niVX6ICPfSqH1Q9Q97pdHRdqqA9FJaeYIqW76fTkwcy5F7p
bhaiU7eh25fPVjlDBkmNaHot6OCULaCJhYzj6rx4v0JZxzwTMxJXoPtv1ReiPHnY
lXZNqzS7DZh8aOvKU8lVi01QNXNtVTH7OmrdSk1o7PKlpJ5FtOVrKp1M2SQWio+J
+i3PxldQUQjMBD0haq8/j6SvVVHWRfCDXzD0f0zkjLWIEkXi0VSTJ6eQqoAjw0Xf
Zp1FBTc/Y+JxDzfrf33YnQF+vukc3TY0LpAaEqncb6IOcRar0zuv0zRObv1G2c6G
Ef0Be5+Hud8mdyhw5SXvzsQZgnHJ1WMlg+vhKORBNHoGQpJ+DBi8bZWUacNoJplP
DmyaI7M+TLAMPd9xJuTBXnvAqIyD/iMjwVsG3dRupSnOA3kUTmi0jDtuCi9pDeKM
QinCsKSH2q12WPnr7H3RIFZQ6q2C2a+bVL9nudTl89EjC2dDirJslOirf7Mtf8Kl
FXkaOtve+7xmGswUR+uhuQ6LkdcJLFl/ghrH1Zcp8Mbm/It0Q0Mp/9FqMMAYYN+B
dux4dYmuklhSLZ9FaecUU4WsUao2Gp97SlQrKtE/vXKRiwGRSCeWpahWqG2liOZN
Kn5pV9U9GpsbQR9fzOo93kH6NcyxvV4507YUj3Pus2mA+P0ryhEbNZ7E/GDSlVbK
io1o7l7r8G2exDdBsoQD4Sdni4Iw1nb8dWpfI9RzgBPrT5ac3GMI93JLnt48HVV3
uI6JG6vHgC+S/J8hYsVa5T25V1nYBCGK2Q5mNJWPJNq/z6uERPpXjAEm86uWypY4
k3yBt+dGb3yxIv0VM8ssrjDI1uGFGnBU4tgk4L+q//KxE8JlCl4ZFqYJW5ANAESp
nQ04kSeg7wvE38KuLwh0T3U4SfqMysIv4qvpO5cheQ1W40eY4GzM8eKOSg4CIyxp
DT5iScf2VLrriUvUaktL/Kt8j8NGLISeyQ+RYM8ffgDu1Z1jfKLDM5P3Ph13K8no
Ui6K/QuHf56s8GKhQHC2dmJwAZbwvK/o0wdXhZclEDEtH5GPd+2cBpio3JmeJ4Ha
X8icTdNVqN8Ljh/GVg9zefaq2Q5L+Ze+1t6MI/hslg4WuUmSS/jE+V4t8cKWYtNN
nVm9RU7aOJz6RJJCsG61HwOhii2HKqupWJ7l8gYY0jQDpHXu7Ewyhi4aFfHOywoU
6yK5ZOzofuzYYDpJsHWBqH1d+byNJpwu539JFu+hkd/MIeUakVsLkWn+u9HyY2S5
DpkDvCJBlafWOMexj49w4YwZ+WKs/TKawEr4jpn5lCx0bccVCl5wh1C2g/yRd9K1
Npjla282lRGAKWuRB5klCXaQexiqPvhECV0X8DM+ggsEaECE5YrQDg7pezqDOFxn
aDitdkFGPMxtSpYNobpL58R7wC7a80md3jyQL1vhPtxBgMDbPHDpxxWZnaDfKG8y
Od00Hn+64J8N+vgB+1AE6cU1o/Esxu8ZG6yu6GfReXjjWkqVjyCfsDZOYRExUvI2
Bn/S1C7affyhV+q/v64MHBKnFtHCEqDawqiLNmx7TujgUc8MdiyAIEMQQX0/jHRL
78dCNRJUi/l5G0v29+OyxsPu4mcgOzpA9xjhqmJmeCTT4Ffiwr+3HZnbnAjVt2Ry
KlR+ZyTJno8S8Ni2oy/HlkUXFhbv4c8MIwAtV6QSqO5ruE2q15m84Z6wVSUGtNb9
xS70ACXr/x3oAKXTri8NEPtYDFsHH43GAiF6yat3E4c7k6JiIROCSPjMS/9G69xI
Qj+9q/5ZTsTw4F8yGPwMEPUOH3oTqiGGtxi4mWYZWi27zzblWzVWs+7CEcnT/vEL
ZDGx6ItY9DDnKsvQGcywP9ZxiCwyRJVBz7KBrkohjx01/jSspP6qIlWeOYmGRXv/
SpB1rX8//+jJ0EZYzntEYt/gFnlBDv9zWOI1mEM8vywFrgLcjG6GA9ogHAAtBm66
dvwCe/Qozz+erWmL0lfK4bR9FlKHUgKEDl6N0dkfdTrVpx9BwbxpO400uKbIZvAB
UFgzIXlSefHfPoPQoOU3O9IKxmyKWLx6GUB7+2hf8st0byCh3tHSG11lKcagx0H2
cGw0RXpUirXbufNjU2rEXQSPsr7s60iqqTbN0ZzO+W1A3pHIEvbbNRcXYyyc/u1I
CUKgC5suoNbtU6+2foKiRTlx6MpvqNZ5tt++pm8miRKaSQXszCBn2es/5y+R77du
8GF3518ke6OboThrfVZbc92abf8Nay6NKwFBmBLoWmdbVg5gcxy+cq2LnPrpIgjU
tlrIovIr9GRKMf5R2CbPytYc4kvksgk6h10OWrhSm5Tz0Ce5LF5iufX+vFwGRkIP
xZiwWt68ageZou3sPJ321x2w7wYyfcNkZQEzWp5f8yn0ab8scDVrFAxWfQyoXaNb
+oth7Lt2NgoULXmP4gJZIoaebZrXaw55s1J5y5mfXdyGbUHxAg5pp2PiPVbMuGfS
cGD28dfDtJ0h6oJROFnT0U6G/8lWxPhA/wYlB3N6ArWAufSlKWoEekeNe6ZU9CxR
JUrZVrSFK278WKgEK8vY1uYu8rpmhlqeJ4KBkO6DM7aCMxFsTJR3YhEV62hoHO9Z
HkqORdChuk5wmbvtbLRPzp4PCxYdd+oIQ0zNwt0nB4ywH5T3BDoz2byEAxNvmgLx
8lSvdjUI1g1tfqQnYiwqiPWgOFi0aY6kdeDqE42DbvZVp0X5HDeXB/77vc4vPZtm
3KUm17WXoLKQu7KAFhX+jgGfg4FR1izwKcHgpXijJW0KjMr5FUHKcncg8aUzrzDE
NnR7oDipAq9okhxuPtcxBfDA3Im6k3QSu8JKxDGBxi7RApx6AhjbBqsoto5taEhA
zk3h9Zhq1A4V7yHxvZ7cLtMv73epNHCMcKHCTEQqqFv0GXHHxaL30ngDPW9XR+z/
ikkOoLnmklMquuRmS2sWL6YjDbJ9Jgevqf67nHdicK2N2VcC5vKZQKQmNTr1gSGR
Adov6w9LJDRQf+zpVt5vzaQdEsBRh4+kk9/WspPokyx3D6jbFHYTUm9RPBsTGvZi
wMlXqdFSSK5EZRJUl9A5BwOe8l7ABbd56AhJ0IeuwmMP6/NHPLUrGQqoIOPVlE4T
jO8vrJLcS9BNsQyYIGGnx+8Zbf5W6GVLtKurdlBRw0P7gKrMmHVN3JemcZI/xJYd
o7bZK3rdFXS0gW0eVwUwJ4cGye3uWo9AhpcVvgsGd149Wdfj+w7K1uiE8RyMBjBD
6rIdBwIyL3rUeE9AYaoYc68wL191mu/5VETrXrFoY0Sx+k9y0ESj8JjLEIOKyb2Z
MhfdZgQ5JEpNVGYhKrH7UiWbmMKYui2n8Y00OXVh5nvKrh44Por+E2tA6qju13fV
BmCyU59AHxs0j+7RR/V5osiAcO2nMGVwjzEppJCe28xumBbIfhZ1MICzhwil+lnL
hI03KuGc2LprVMYPeVtsR+z4FlVNdYbr41MwEQj8R+iYVkJ0W3EXlB+MxY7t5YRc
meMTaGvWxS9xqrp6CmEJ6rp0tzUxwcQyz/eitPqxdBqn52PtipgqAQ/4qYW2+y0i
JWLpevQrKOxeEV4yJxwETUJKyXIhqe1FHyOi43gPIsriDsMNyhT4d+EVUornmKtw
cMDJoji8r92pfSfJEXHCzKu6jD0ogB0sUSK4xZoczAV1WPpxpj8vCzWB/5F4aE+M
5q7afP5TFXXYyLSWg/ODxfAj9dRpt+mxXvMGQ+UakggGPXxRKakLn4QZ24xUAdVf
8prsaED1LlLrMckJcSDW9kEKg054ZfcCqvQPFmfbqNJ4iDtuHQhOrEdM2U8jcdfb
n2JRSEpup6gut/KJhKtH6jjWYwpA8A3L2ccteVh2Fg8W7LeDtHCnUtsRUbUhGAS6
Sbt0MKAEDZ88ih0QpzC8BMfrQUz6OgtemDBTjEoR9ln0/Ciaf6aUOMCBPC6IEqD+
OLJ+He6JhNFBwDWwLgtx/DRzML0+O410FDFzlV4JLz6AFmenwWK2lP5eFLvvWFcx
Trdbt83V/ZcxBQxw4vG09KomkSeP1hlpgIhQqf0j7RI0sfGpENf476hd4mCp21sB
cILjyGsLbTOVVDrRs2f/U+0n1+Fga5iCCvk/RWh50ioDT1TcuZyY9tLlmsGhMsBi
k2SsznWQ1iko29SMVyCFoYARvPBH6SHq4luP0tgYPjzr7eHVXnk3IL9o7tLBp5VK
bILN3nPlgysKwDK9F9z7fqhf++k/BeGHTzDJa88FU5JQfPgxR9qBCk8dM8n/A2ht
OefQB69B8SYw36QqUvHzm3JtdvZO8dSyuRmjGpuUgHEgjlEAv64TcxFJvQBPYIcG
kF83os1XEK+DM2NG8Z+9ZTrgM3EYa+KF1twpAtEkGDCZJ36LI/gZXYKUYX1w+xm/
fdAbpx3P6tqXsTiwDnqNL125DbyItQ8kVFyp1dMXeTb+UG24BhDFyyFneThtucl1
u9/t7DVSOMsP2O/enKHmgaWnZPxtX5krUg9I+8U9UTIxqUV8ZkCs5ySxr064LpSo
pQdaRxMlGeI/kjoOzS2X7TfDw3y0zmYcV3dvXwEnmCXD68L3hHOIl/MTed61FD5v
sU++ORMA2xiGKCjAjmPVMjFgracg/he/xjvLZ4aZcAWfJvj5mI9qblnSM0HWrc3B
AaM+CoG0x1X/oV4ulRX2NXH5xvyBK0zvP4cOYhVuCG0CFJJGLE1iXVo+NiCIy1kD
vrtBAsTyKulWL9bzodvLLGkzDU78Ksj2GzpqvC0L+4nLfKodFKjhn+MvaYnHS2wv
CaD8x4gKgT5aVmc2L3VXxR3yPqp8Dsj2swdnOvHdob9NxmvIO+rnqve27n9SBGIr
Y2wmFYf3h6piB5LgsirX4aVHPXVxJvsdVcikRXntpfnkkVcUJnzKDe5IFOxOtUFN
PniBppV6ThProuPgHSs9LqDZ5x/ICiKnBCpxO+NiqPj473vVra8dtPV/7lDcuIUD
5zEkTWjuRxzykWr6tCtdoRws5TAZsK13QwNz0erMehe8WVfZEHi9baktZ5gZv6OR
GIjhYu2XvQv13O+48+CQYl7TT7w0/LtUfmu2j8mZKq+Vv7yDDYRBd/cK5ku758Yu
UhuH0rHX/van6s9m2kuqJpNYed8V84Zc6X9kRR7djhd9tEidUJhKIaYMdh7CWuCJ
r1IO/bzAoCIWkGWB2A8ZD+VuY4WbE3Ujr4djE+fiPajIk3a4LQzXAuAHGt+e+AmF
tmzVX8XcGJ9l1DpZ6+9Cmi5W9KuSyP7wSv+x3YsLDn8urMUKf8jVew3eH26Z383E
n99TF2tF3m0A90k0AN7G97O5WShUTyzSyY4TzbB173GrZyUl+DJ0PT9q3uMsUQjG
1DO+pCat07bfcnhU/VNfsOenOMa+DZtYjZXxm4ktvA1uA87eQp9i4jhifVo5lKcK
WVNsr8DLZrXbMbXxNPo2gQcDfAraxy06Fpqj+bleQwvtmxNdr9anwQLIA2kCfhrN
wjgDxnbiEajoK4tcuUEobKkmNd4CWHuvrQxUEYgw8dCnmVQ6nE7eV8xIvWaj8mI8
q0kzuyTVvRC8GAKUjTVipvviUasM/tuGDAsOPasHW4oLTbaOQdlgKP8Qa3Y+MINN
G/G8VvMsFpQbnNh38ezpDiFW72RAEMmOu1dl2QIVZRQtOQGQk6rADa9fzmkjnh23
7DxzuLW69A0RAPQxVNF0BXdWq9aWW0kPOqSUs3L/u21qB/DFlAv2pGtPq8Mru0F3
khjOKbIQUVuj1IM6vChCUVVmizE1SY+Z4swwJcqbjqwOCVVDXqHRmTWClYixXoiz
1Jmb4StpQotDqxhr/JwAoe02tw9ovkFtM7ySAVAopq4V12w9UIzAFtmlrlrMgXPr
6SMKRUvDprSP7u8N0YmgmicwOktmBguRHUQUnji/IoAs3cGBVftAx4jjXlx8axjb
oVxrXbpPDQ3fWOV6zUtAI1lKynM60R+U3itKvogBx9Bd94T9qgI103Yz+9+wXeb7
FGYjWHaHY8ItojNr/AQ5BCXSuBsdN60KpLvz0RL8tXnAbRZKMliMpub5lnjEg/DZ
ji+NCtAiv6l8Cmt6LFwvQpOnyBuZNaiO32DM6hFM91S72QznLex02ldd/t5vyS+o
ilOUFiQFBZZZA+M/95RbhmxNSCWguqx30cmFg8b0T+fn7BeIs31kLJ0Z8Qbx9PLd
qbySWkb3XlEVyEkt/60G0+HAzK3syJd6f2w1nP58KpOBh/OsB4gZlIgLE3kpsqVh
5ylSLDEycYHyBcZy/n/o5PcAauHaJAErEhUZjnTf8ArDAJzlhjR/S0Qo45TO1WbM
+VHpfmCaEUH54qaAUTqsNfb1e+QsLZlnZkqv6pCrckJEXZRDpc6kxRLEOFKtralf
rvWLVaC4GblxGMRKKiSb6X9BukUs1fowFvNLC5uJ7+GX0wAM5s1vqozhk3cXu+B2
PY+nWbgseANJzH7w8/E4XDP3aHj2PhAdw6EfmCyA450qr+3U+V/KJRKA5DCXoGfw
D0OvVKOvI9rnRgyYUL547SRTJL/OLn4QoFXjcAKnLUyykFpH+JpgTHhApy0Txhqs
ELK4h4Lq4snVxdqNdXb05yv9vf7rCdYeI6W7t9EXmWTtaSNuXwDecJG+REKvY1Z6
kG4RX82nnXFmVXkyEHSTkbTw2BlQ46d0krH/i1iVYGZ6UU8fiQWRaleLwNoPS6so
xADz8dQa4U8PC/PJ7C80FLn+Byu5ET9pr/BtZpV6iZ1ForNlxGyXfuT6jN1iFUlG
8Tr5wXqn002IPA7YfBMqnwRG972rnjRH7MaCbOvWTqNJGceqEeIQtP6+Q0ganx9E
R9xZFiWa/eVyWsz4M0vkNncaWqS3aJU3rEnDa1K0b4vOnAVQft5mlRbuT5kriISe
f7/67Hzu3kQVgj+BByxbCti/zC0iyRo2q5OoP02WxMgPh7zoDcIJxQiqy65u/FlR
rsH1/G8VQXI233lBk6yl9w8ATewRqOrTx7gz/5OfOfHK8vcM/JUnnpXOl9aJZjRF
2hwYDVw30c/2Xg72roV9GrIl4oVPtPDiC8M0Xgzup6vsZ31PHgiR37SK+0FJ6m3p
BRRn3IFoxk1LhNVjkqqZysseyJt8yD8Zd8A8dJP6EtcMOGc0+gP1gXAvsy4DLbEG
zPpDwJVj7R+LKYUxeFJwpGZnug91M0btGbzdFGPotxxSYvPutkJKVUCipHGYjJ1/
BlCIE1BOFeMhROaTDjcKhlwzQovx2k9HLs2U9Hz/eypWsn7qTvaIzLID/FXrRZ0b
2Etf76wAQPTWvT8BOglJFd+o2wcvs/DENwLCBSo7/pR7bSN5lUSdbjxS4zBe9l2r
htv2SVz8nBiIXH77pr+H2xutiA5+7MQkTF7lA+snzeRBbgWWvH6kiZbIVaW85Yat
q2tQCAOqr6nCpDiexJ5CIpSsXWYmDR6C3SPTDjCdAYRHBCzE6gIMToJrq0W0dplh
+nWkazVEzWR8ZSW7tYbSry063aoa8mrSdpPIfGR/WsZeokcPrtG/GmLczPRQjhQS
lABsRI3ETMXpYHUwsn3np8VWCha0POhGOlaLEtSaFe1ijsjVQn9mrnGIzpiaScqZ
XeQr7uZOQVpYhO+0nL8etuizhLon73OBEpA1k21z5kLel5BKNAHaIqAo16EC+mZE
JpL8PizQ3h+TPd7GxAupO1nHQ3J9+Hb1yXmUkeThthqSMw0kWfqRx4uk04WIRT5g
cEpxReBlVHQCh0+627OBqCJ2Wv4ztpx5ugPI1h39fwdh08ILlKheFcy2OQOvIYou
Lo7BT+OO/bStTJhs/y6MRoRgScV9touCLMjqyMCIz3J5xRibWwVKFOxW16ZneQTU
rmm0a3jaotoM9oEJChblLi8i0BLNR2b1kbNG47Jv2nH0sBHaY6nZLbqH+/GJpMbX
8ZKDAHnVJTCAx1f4ymALGnerMurQLYvY25X80/TcM7QlRcb1dcpRcv4IOuo8sI5Z
2fGuyWH3/OmgNeg1uByvtcBetBDCDa6R7MTivsvvCiFvwBeLU5rPxbDKu/3G204r
dF7/PmZDFelQjccbf5AUei0Sqzwt4w6QnfGr2fwDzobljBlOHIXS0j0M6SLIV0si
ueS5VMDf3aM9N/fZNmsnTDVZ7/dj8oOIQu30c4Ou5vDOTaF7P4oZ8jw8+BRuLcFu
d46VsCHeJEC1SA79vtWxHpJQtoSe1EEirYspViAscrrHfqzmI6celUGjxvkZkpYo
3ftMRS+6qy1ix4f6oqSTkqC0NmG1LnGgxz2wZ9pRnuEETqganW0DEX3V1l5BFxtq
MbCu/reQeaJVTsGRL5bkdVyE89hvr0/nIs/s4GgLVkeJSu9JK0OagYRoRJr1E8cT
WYk9QRlCeBSO6wf6FukHI7WT2IY7441it+hPRczTKfLXCX9PHaoOBPofLKzZ1Q3d
RBfXiomtAIzm854jLsDhsTaPXs3AuoT/h5HSFGVNJmaw3+2Q1e6tjSH0Cs1MfZ7S
iaw2UgMpVLThflP5poyUJIrpadTCGUt6o4CQ3q0qdvyxybrU+v4g/dvuaESHcdcf
uTx1GeLPn4UfZZlH5Phs3LtfjodDf/UpW/pLw1+skuSRK7iTXJEkanUGnhAaOlZO
nrVmxwpKWcjToiNnPUqPr0T83LrPaua3wtkM7r3AE6RGtzlhy0onF6NPAa8ixfhd
8q5HKMsgD3AXqiJU5oduP4sJvZgxoH/fAdY6G3ZJJUHg4S2uP7Vn/lXa/pXc3eMj
2SwEIp1UmP9Jt5ZTibU7eqepUPloXZc/bKK64duoQR3qDtJDZlhOEvXAse05ZgeI
3H8PJ6elQX13KkFe7HTyWa0lF92a2uR+nEjL25m1aPGWrprj/Dl6FDWx94vtkOdv
PPoesDepIjPiCWMqv5W75SwTMn9P0FrTU7sOKtmsH0zcAolf7RE1eABy12AMHICb
zTejdldUkLQ5qIHcpf7h4KHEYQsj6rVp9T2BgaVuXXAyq9myoFmf2es8bSeOq4Pf
vBcNzdwl72ysh381JKqmWU4F89+JM5xlWzuYkE563rDa7K38Dm5TWroso5yEDR6f
ZUR56GMwxTu5dvpGQSbHFkKqOr15bwIoJCqsEiNKChvG3taIj3a4JN7J0IsqyQrw
k5bSfCFjwG+my67oUAjiIo3rYflcz8R/x1p8IATCrisI/92umo/0HGu6MqIs606I
pF8mNRUmAQvRZV4pj/AARc9GKtj6x1JwSTzcrWxNNxV42mSXGfxcdciCxJYRZBLs
n7u1l0pg6YkeAuVLBvnHWpuvE/C/JJE8hYQYxtqIrpxLb8n6zTWdofZ+ns2GNlAm
W17YAwcISOtG2n/ASLAaWfB24mGBLSp3XAxP/mlobZGLPXKqSvLAHG49pZZfX0fB
tdMi85wFYQg3eQQHQ1H/LmcuAPmhYGopFTs/42qK0w9vZjs5Q2dYd3oX6lwzKcEt
SqFjDfT9OJFz3of8WRo52rXsl8nv9kBp+8DIcUuRNig3wHWh6+KbAGCDJhELEA/L
GJaUtmeClubVoz5cHJuPHqg5MniUhnWGHajHJB3r742jOedOc5QXWd2hOwdL0YuA
hU8dzdtq4T8yxKhtL0Id+xZ/ZwOla3C75IoFeiLt19yNAPwH323SRHtK9LygtYfQ
AbVzmGJSAKbn6OmU0N3/xXf3/uobq5kPF9VvmzSuJ6PesiEaxHz+iQM2n8CIsCga
ckVxdradPMhwym2KTmDvWDyLsqNNj4+dO7NU94Yp3GY9FvOeaWhtx4QJ3vmj6hDV
9f8Q+iPKwnTROAgAi6lvb07YDDQ9SEF4ydFhkQaoxpo1Z3xC4EHuQ0+PQinX8TYb
1MXHkUWMIVMVv2Kgn1t3y1fozrI77+5zUoenzhCRm9m6qASPZBpQg83kYZGAExke
4g+wC3JoaIl8ozKJZq5or1/Oc/XuNomBepBtz/yelMmuIjGYyo3PrSmWhZ6e/biK
Ib56hbWrlFPZ1TwnCL+vQn3Yg1AKyW1pu7rgr6A6lgmGLPqFgsu9N/9mki50iu4h
wgzcKqIQFERzvXb6BX+65DXR3xE+/27OZLDaeEcpynnzPUJd+huSXXAf3eyYlE/R
PEUSpFRSH+XKdaFn222k+MTKaorDNZ0OPbjX/uiTZ+XM15blH41ahXvUvTD7KqJo
Cc1wYCXq/ga4RsLI3lG5dT8c+FFBlEUw95Po35vHNYXo0fhZ5yOgWKupryevWvLv
tYef0er7r8XP5E/4ChAL9AIruF+buGatBTHWBKpyUeTcmruMJuK10LgA8jDlRJoF
eKXOl4e1c93SsTPLbbji0KTW8w+KDjF7qYteP8qecHw2NQhMZrA1SBnlvcUukSQs
Fo8T4n/IYo/j96QgFHNd911chyYpg5o0CiK7T9Djwd2CWwAxiajubFHR/KeOQlk3
9hT8lTNfFqbHEiw5iQGqnBpY6TwihRa1Y6y8ifr2cPwmrgPfQm3GAjCqxPY9itfT
JPyCeCJv0x4hrK3idjl2XakyPcLQ/XkUPXDuJxdVf2xnaE0nOqD4P8YVvcBt667m
yTRWp99kf48MUQDH9asgVoJcklyQcyYtIxK3UPZLfol/IYRmNvkzF4Kfc9UAUIXM
Z8cWpw2KKJC/mJuRubC0rYa4xr58/EU7t4/wpmuJA8HrmRGE+7MKRNUitA1pj/zL
y7JI5Q2FpFcl5y5ItUOuFYaHlS5NAy7mcYdiV/ZDYKW4grYUSSqJ2QAkEdMg06SR
uJKrHovsoPxDJRahy7G0WMTdOLKhhubhUeQ3t+p0iWqvEpY2SLiEqTHiW9pmLp9a
ZNMuQjewX3mKB9LbfwbEA7vLxxyMZurHPihRDRXu1gvhNLiA7vtkDyWkzn2S6mjH
w4IeABT5+Iiw+EZ8coj6FK5Tjxz0+7F6JJNZgCRHvkf31/dZs14QeX3AfBmijUdT
GCEknTKBzJjpVQL/HchZG3UjvWTpvrtCYyzE9Y1yGKP2Cmgj2aBNgw9wnW3s4M4P
cu1DnassmffLIT2AY8Rnw6cJWgaTSqjO9rkWsZEdj62V+goAJXlnmsR6i2rKLyek
5/zmzHGT+Q4Z12UtuCWtkE+MsSM8fZOwZowCDskGRU+XjCEhD4Npwv9nX528s0cm
O15yw8bpP7mqnTNk4BWLG9ptr5v04qLidnM8TiJwbcgNwpr4Jm47aGUZaKF0Mc7r
U53KZiIsbtzxjB2h+YcA2UImbfxanzCvcDZ+aksrZ9ifFIMMwn6qFDGvf2tlpyBy
J5EUGXsNuNsLPFO/qnZ+Ryir2k4PC3cAnjjjCoY1kFYCocDMNAWb9v0XirffnmLf
ipogZGlZOyDt7wD2cV8h0/uZI3P8DjgR4Qx53P1g2NZp0Emq9VeUZE9YzvqXUswY
RYohDqhJrpuzGpEtltNk5zR7os3TRqdT+MFfypSMDuUFJPgzyosMuF4ut5vQbmuV
AbjxP5RkwalsZP7mMbfH7aW0ycMr/79Ch99OOf86nJhQnsiyi2i84puZPgDA2+gQ
jzNUap0J5Y+eodVrCW8Xhd5bECCxeRm0IBYRdafAS7RpnV7AqF16y4DJ5TpbbYPy
kze8HCxE+ZrPy0Mn3A/b8UU7ZYW7MlSNuXv/jLrD/HxC6vrRmAKobM/9QvvsiNzF
bRti2F18HNMoS8NRW5GUGEPa31XGFfnWEvbGkyiWpi0TgIg0COdocdalGd52rwON
H61WrMuceRTQrKXnjWF2Ng0CQ12+xM35u1DBc2LtvXm/LoLA5jEAwkMyqNIfxMLr
pCX+lvm7U4VWlPXPgsD1kglNTnVrfTpCLUfysMVFSxbRAwtddtVgfWsRWJlLaiZ5
NoQv64Zf6Pd4poVVtND2EO3qHVSPQ1vKDY7osY9Sp6ptKLJ+UaOW7FWrEhLxZEVu
hUayOvDI9MvBxuO/szm89EneJsq7RPRQkE4otNmkUlXsJGG7WrrdKja2HeQZQJ7x
APobLpg5c7iBST15eT3AmiKOdib/b6pRHESc9yjx4+6KG+G5KVrRX/WeDv84uHF0
QLd2XR5MVxhHq3u1xMfHayASBAvqllwlGIMDYVk/gCjwMxynKqh8V6QhorB0Su9j
Hil7BnlL9NU4nutqwK912XgtTb+6/2pwzGjAm51RDZl9Q1npsZVEbsyxx4AqyLwp
BsLEwHlY/g7vZPVV6t3dsgnTxxHL96I8ke5hexLIKzhfJtiuq3Vi2+Yb0grRTJlo
UMLKgmPkMmVR0kWeU9dLoqG3jVq4acZWnAgDGMGog39wdmRy5uFgcZvlT/qYMO+1
q+P8J5c+bRRP+1LchLPh5s17DPjO0RHUCR/bpRfSQv5u0h6qasEI1/SYu/MAnTpx
a/yBkynT3EnLELDSmMj+tFQihY0CRlWH+UbUM3v9x0F5CwWv9WPN2fepTMvB+La0
D8mweOMCnhF4BHNPuHkkMhPh5NVoDLVmJLupO5m5EoyoCtkEaO9iQyX/zmYD76+L
khInFo3on5BmFh1IpGA8m5jBU4irARiLINn1UNnxvGObNzw66YzT9r9ux0qP2FwC
VAKCWluqPNEHWlQmSB0HhfWZos4cLkGzKvczKKpl1pYWpCtBYM3BpIb2LfD/EFld
getU4pUQg41wgYgYC2/8C+59EQKksAwjb5x4wYFJGXfHYPBv1BwLtsupgyQnvnDY
NNvV6wf4nKVa8bPvp3RzqlV++P41doplC6HqAq5r2o3Qj5vkUh/A2+k+Yl8IxDxR
pHywGwXrX8Efgtg2wxZf01h+Sb0h6uXbHIH9HBxhxQKSfF1465VOtW95FQo0og+t
Y3HTEoybTmD2VShQbo6gTTp9KN98PFHqNboDCrEhMt5b64tpqnvVkpt/4Pe+9pGN
oPE57VYNxjP21IWCuAMBjXrpBKUBYVeEVDorxSJaWfOJlRhKu3GCeHy6vYkCdSyo
ZU48nugC8ttBp5FY5wfcpTIM9rZxMJgm6Cni7xwGLsZCemmN41arYeET6JsXs4zT
IBZSOQTavIxcu51dR1EX1mOtOtcHcFtW6v/ZgJVdt+hQvIQnhT+ePXKexyUE02dw
JdnzK4Xj0fv1lu2tn9dp/Rtd6yp5LVVd6ms10bEkmiCmvTHeTO6mrIR5WFxEoojy
TOW23cjE22nenJyfc276OGOTMVb+Sr1x+3nKBPSNGOJadFttYoA5KlviM65PgXZt
P55nWTgJIkfN6Ie4Zbb71YODPh0HFUMgRuADLv71Qt7zWP9O9rJTW/ZgJmQIy/Zf
D13czfEFsOHD2dLSGiyBHQVtcruwolCDa2Al1vPFF2F74usag6Bq+yahM1tY8B6C
nx3MklKmPQ5/RMFTJKGorOSrjZEDc5BxRFSL01I9IaGul455jDrTnVM7gLUotMEE
qiArVfHW80giY+9oRHUOmxRPIFBcpe2nWXNnyO3fXwrMb/UTXiIXlyxUKrH9SEDX
H+GlbkqTpiaeqPMDCBjXknAmI8VtfZzUVvexQO98EM1NQXsHdoYr9ANjSZqhv+P/
bqFQNdv606VGWbiGKan7QtUpdESik2g28a62Wr0xJWfi043rREWxnT45HlmNkg2F
3e/glb1fhwMlx2s6PHOqxIC+7oHib0olw4RWUQ8emYfyAb/BKfA6Rzkdz8jgLBWy
2xSrxzr9SYTU4p5oLj0JGB5y9v+hmVL5JjJDYyYmHqbA5gHPDDSzp96Syb2l6Cch
aztdUz5sjjnbPpnUqBNO2t3dxTPe9OhxLPnQEaSfMbUNE0MudD/y9LLdR82WVmZC
VSaJDF9QRuKkg+LYSWNwqQCLXn23S2KujWhFm67nAgCUB1kUIElc8vnKmoJTM+L7
0TkwCd9WDVFjwVi6yPzAfNSQzDS3F2RUfYYcNBDGJLM6mfgL6tJ8ETykeArBhjlH
gbitgjhO5kHlT0jIcFgwzMjPvl7T0oDYCwAET8/sU+X8AB7QglV7FRRAK/P7OPOv
ItrsVZkQ4ZV7sE898usQWizqpHkCZeLJpNMR09jLiXHJ8OSlIbTHrkXUJBpjfm/T
/mC3/MU8dLW7ogevDBGiXVCIEQ263c9i8+QlhQeFLs2C5wCxfugx4H+WGHxdEcA1
PZLUCrmYxsLHo/oxzjnUnsn/l/XgxKzs9OlM66iCg4ujEnLPNMWn2/gki84GzNwO
IxlTEStpF8KZPqhbeleQLwuV6NHdlu244AV5NyrTTQvLkyEdul5GTamieSIa/KnV
v+TodbFUkMP9r1KhJY1Oh+bSYEO2FPSBVJ5jjmuv+wBo27GR+uPL5MJyGHsozFrC
Q/D7ZwF3O5yn90J7sRYimU8x5gjjCdkni9EM54NRcAb1DrLGzT/vLY7lW/EZczC1
BsQu0inW252kS5xAy6sDbxYzQvMpAcKsBF9nD/S4lsuP3cN90FFI+5kn1s+F3+xH
1KbGllN0dwBcPdrEEppaafzgIQAQg59FAOkOT9O9MbVGtiJq8KO63jcI1p9V8fCr
82vPnneT9U6EDcxX7H0kCdqk92GMdzGnJsOzMnQouT+LS3CIYazioL+AMKO59SS+
cknbY7xg/KvNtTmcR6yB1KwfsGtDl4X/KMajTavGACwFIjWP7yHjqAwHHQg9+b8c
OFBOYQSBMM8XGzulF27Zluxgt34xB1M0WhA8E69e2eLESui00Y1tAkwl8jC3AfYS
i8xOolv9GpN50pFEidgF0zTJpTV5yP5EoHQVf9zX0CftYG+env+SOOcngF1MuAPJ
ipDrz8xAbK9w+3HiZcKEJRQNE1+Jap6xuq2quXZXuEAmVDlsb1SPh6nPGPBXQDIC
KZVsoggH11tkQhSN35/Yr4ZV0i/QR07SVHfmW88IqLbuy4r0W5tLRIVrncrwcKZs
zoS06xoDOjZ/TDcuZPBXDW8Ofw6yB2yYg3rZarS8T3viJiXp2DchfJomyxy1yVki
WznjGJj5zFTqU+yuZxTXC5JHRB8NNkOmNmUWOa+Tb/cMzkh3gxDKDF9m9Egg6CjC
/UjXV0JYcr1SSLbZyLrmL2CQaKjy17zBwn4f6UCzDTpABo+oeMI5wS5862JN2X/7
gqZzYFUxVgctxZgKsl06jV+s0UnIGE/rj2h5GTEsh9tULLf7lJNsn5HsrcPFFlY5
xbDxrp95oXFfweZjGH0mtY7SelbOrJSXQSw41YUoceLkmrHrPFyMOz41sP+q0Z/4
t76JO1y2nOwxsX/ZkWeScqUxTvRnpjr6g4mTgawXr48YhdXnvaXiRBaHOp9qAwd8
VdQgR9DWs7fSdCVcwNp5EjJkgo/QRKtCh1C4KCgYtgHGojXAVt8wb/kAT7Ecwl7Z
Umeah/nTRRpjk6Cg2HSgC3TjmM0pCC1hqw8ckXAiuGk3Pv/gkBv6VzsGHKz9slWf
WtWQmTWZfuwEVWyRcFbzHXl7jKqWdYFflXNDe6PIcTDMLGKWq4UcUunaso9Vt1FN
GG+sv6vnf56Ntlyr4EngYUnPQfeFP6m/b2P6D0ysYXYAahhDV6AC4eknb+WYV/s+
LAca9Q3Ao43XdyOl9pFGM7BnTbjmihT2Rce0qluBZpMvcaT8Lxdjsj0Ii54ckUpr
9WZ0wylufV1twG0vjFMROrFj8XyOoQGzWZZHTlOBgBQWBguUhUb6MxKZFKJJW8Ki
lvWfZYp26Yn36AL9H90VxTINmZ4o7+gXfrRJl3uNZUmUJjR9JfB3+7VZRL4u4nZK
98RZQ3o8+DXfOqVYcA5Y8wXvbUeE32BODEqpLzkE6ZFYERcPgqC/5Ts2bWrkw1KR
eFXQdkvoriQgvv/aljqy6EeN4k3T3rVxBd1onxJMAd/IO56Mry8AWeFlYh11qwYE
4IvSCF/c+4x4VNPUu4kQitIj16dKDP5Tuq8ZwZWktvGFw+6/hvGb0RPB+3qj1uRi
WNBTJCK7n1MIwRaUnhiWA3uiwOzccHsdK77wrFB9JqtUYgAES6dGj/G0lJny5EsW
JyijXI3kR5fWeFwd9Idg8RiiypYzZSnPUhtrLe/0LC9HiTgIL7v4qXc/HEiqfIyZ
GvnXwd5uJlypCIG6BL56aausshRS9NSgmS3TwPnk6MP6U6UVXMlGywk7K53OEjzF
uDGoXyls23ia8qgo4K0mQp/pyZgDSnxrDYcW7yjhBNjccY6u+2H4ofnLBE9KwNEW
Waeenqo8G0MIJfM8RGTLeJiO5A51ZDQqTO1Ou6T3OgDdYzLyDiCrdUlLgssYj3L4
ZBJP6TsAUOayREuXV2yx7SIMNL9SPCb4G3TbwludN2Y0L23tJF/9CbU8GbdH9m47
IPXVgmpHtVb+qtbNc2LXiUfRhB3CrhxDv6hSoDmdEygMXvbJQ4BabyfUrW6PE9/m
9ybgZT/6l5223h4ho18IDkuKtdWwo2+Wm4LRpdBtC6etLbDcC7GcVJMmNovLyuaJ
Ur8bxqqWxxlMTg85bjvthmJLQ1D2fKVM397Zx9txH9D/tu2+gFWMpX3TM1RzSrUD
NSmCeEGzXN/WlGpMcNYBArSXVyeoTCDJJc+waNx5bT5Tk4HTEzF9/plwbAru/XC4
jJn3n9HgP1LwCiM5VWE3erNR74QM5vX5/EROktq5z0AXx27Oz7eIBMsFGUIL6hH0
4kAzttWYaT57TxEYwex/NUoVwzjSR31gYL5lpo9W959LEZaXR86jr1+AOGt/OV5I
alRioSmw4N+O9Wx9X78A14+okyWWwJr/r2D3VTE00TXG6/GzQ6fc/w6djN4Xw7nA
grt15XOenJziM713nHZGdOMwW2uYtQDGBUujedbkr33kf04UR7VdsJZ6OHNU6qs8
P6ktnp85kn0i32pNUzXbOwbX/kw6RgYfEuFLUVpgsUBCwGu5TB6/1QYo3gvI0msG
OMiCofJ4+At3P1tiC1QWOB07EvCxQArFnfXffDm1V0TBzC0fF34Vb9QyrFHW6KHC
g9W5dG2X1y87Po+RpJzlEM17G+n4oNTI7kIAHyJJtWqtsUspryqQQHmDaCIdcMpT
edPlLIiBVTigxtY/9FVQ/h4ueoyp9e3/MiVYTi/sZCRryvKz11oV02bf1dd2ES1a
focbpP2LxIOpiNnUFGHMf/yKkB9QrXcGeXUCQ3wffD+jWDvX95jCrCM3MMnh4AQX
87dHkA4EvnEbOM8MvE6D5hCTRnsy9F9Sv/B1zlZws1h9QR+3XECx5N5XlyDhz9tM
Zd6HGcdTdOuTTD6QdgTZbmfG+5LWYgwq5CvCNwpfpD+MddgADX5D/YdFkLlWG6je
VfGg7namuHJphlDMv72hEeWuIobBZf6+MavFzpuIJN9aKXahPl4/W5qaGGEtnFxR
4xxBLm3jrowGGRUaEaXilOhX9wU7ldOZ+P36kuYJ7Q95wQ9+GvW96eqHmvpbXRiP
q1X+v+QRmXoNUgeXE14KWGugiE80b6Uf/5558VUtcksHcGgqg33R3zi7UF0udcYS
IOxJkYU4Hv3S6IO8NmEH+MqTbUJlItSM4hkPwCKGJUww1rAo/upIe1SYLcVej7Mh
kWk0gfIfJlC1WWRRjF/KqT8rlrHZEdRYkRv7tSdNFIMeZQyaa0TSsbJuLs6aruRB
pTsm+ABo6ctPB/RuWzq0XQcQ/acsOo7siNSlxBxSoIcoIirmXjBEwJDarqQZzygS
XOTL5kFUcRr6xbu5/VilURFduHMiq9sJfWKT3IMB4pnUcjCy12wJLFz1J5wi3toi
dQaGU5ARM1F+2VTzVueaGoGbfVUE/bEZjC1ajhWofjQ8Ix+gimikwM/ZQPnsnyqr
HlpTQRcRNPSCORjvX/o5KRmkNSLt1Hac95Wgha22wXNwzQstyrg7/FggTiNaa0RC
sRAnpcZeiZwy1imsio/R5Rgg62rLercaxNNuwLe6DaoWrvLY//xU7dmOI0yNfQEh
jJpz4c+7Bc9O/MxW/8koHmCbsk0mUQOpdy8cHL8Q7xdigUc4QdF88cGIOpGvGRuX
DgtBjSBoCf1RK6GtkD2f3fY2R3445wtps2610q3np1pDmiwCp8mqB8a6bBZHcuje
KTq4cTy+M3bwD1Dg41LSfJOAGpt9v+ieqGLaUOJOHgq0FI48bAyxKyq0HZGQoJRR
hSDD7a7RHZd03xUzoEOY+6ki8vFc8v+PQuOEl2HGj2BC9lb+QP04TSOleURLYWs7
yNA9ygBZS631JpjgVuurYiWjgzc9ep4SFQCnePBpomiK/x+9+4RmKsxDDSE1LmRV
Sgdnxc1P0wg3tVEIQrKn+c3VNX9LvD02PGMfSaeoAI3uqokBHiNP8JXuPVBinBU+
H0mMXY9P9/fMGV6RX5aAyhCQRgxFE3QqsuJI616jaCWjD3zgZ+nUxe714IVQiwy5
yqodiFcKJtWsoK5YcrnTdYurUFQBreMiqvnXaLz55tmIWpQceqc/2l0I2EHYIB4f
uKxu4h9kJ5qkSwWhwQYyVwXyZuOztaddYXJI5cZKeoFt0juQ0DSOnFqk0BVorHpu
hZy7C2zcXHKH2fhenteiRrOd9uA8e6ZJknXJ2zEWgXbnbDywAE3hFztRb7ZUEPxX
AvJiJiTMvGnCgHs0WS2QKGIH7cxuxN7DKPeWoIHC3HSsN0redPWe3+UjIKoGmFDS
pOTkuQQ2wKRcKHwVGLk75Wq3o1MKiEqNc10jVrMD2D2gFyotaRc1jm+L9NP7j8Hb
bKNEb6cNaAnWVLBNuj3gPKjZBwWuaLoAUN/3P4RAS2jHJ5IaoAO7l2VT6eILoQqi
5m9Em3loig04GvzAbZP5R6ALMjLLsWodlaqPfRvvs8NrpMQoDilWZ+0Vr3WXCzlx
2biibMvB2Y0KC3WtXKIFO4RJHl9ts+lJnMF5DoWI1FNUcGRscN9chkU3uecWT03k
fbpwC0vUCl6dd3NuHg7DtXUJ/f8hpNqEIgOnm7lycliTeS/BCYkWGWI7n2hVCAGI
cdDH3/rOF9B8jVZT87ydqS1465UJpRcvwhYynNkMkE2AW6OD3aF4QiCV3Vbf7HNm
e6FV/HJnPW04ZE0uaV+qM95QUKERp77aVjfx5MzsGGKqFPPOf3hfJnnyrhLi+RHK
EgT3cHncdLmjBI3Iif4nvTrq2gbZ2+bG5NXSkdcIZvR1NldaTE/1RMm20JysZBtM
CzaK1GRAS4cZjlE7f6JCkcBV5W5yS2dAg8uqe8C0y0BnWfj1+WhLjhp20Lx5+JSY
RQuN/JDojZGYPUbmUYluOJCv3y9d1+rCa/Nq5lgRBmbF/mSFKqz3hvBOlWY1PKFz
FDvmLc/1A4wL7+P/qxTkBhuvxsxI476bHyfC2sSgO0ZtNmwtW542wOmNZ0L2VM+4
iSYcalhYkZEWQZohISkkeUUETVODqHypk6mw8u44SF7+z3S+piV7cylY65Dv9Q+l
obMbatQZI5xrNI8uDfvjc+eNNw/QM3sc/x6tcR0+7+7HGB0Luu7+BEOcU7CQg9Nt
3nrJpVNiTXFZxPjSCxMvt3jnAHOpVNdHktavuSt3T7aeTKDo22dWOIIfAwSwlXcB
D/V6NHXfmAzI++pERHXx485olcl5DqICgOHZsyj1qb2uPSyN5o+m0MTMNWyQoVrK
9tQBeVZAVsmCD6vcq4NnZs09uVhL+aoMjE3rZ8ecrCBK+pDnGIWMTFzIQ5wjdx1o
Zhcefllop/3nr27ThQi9+RcHQ8Na0SZalVO3YNiR5jSS7xP/KE1UKhiSyjIaeH7G
51gv7FKHXeZ2RI9Ta2QOVkzXMb9PAq9UyzReu7Jfrco7Q49o4/jxQ8tcmiiKOp+n
3SmuKvuz6kYAWOBCgi9vSYmvwiFkxQG7xIWidSCS/JnOz/lNHGILdDRNHe3bLMp+
8cwgHu4JuFHtGl0SOsbKA5cZFrFSPEd3F0LzbcadJlITGFFxTGzsvsbARmteRySi
GeE3EhrZfs42HJb0JujQ6igzmgtFFfV9y0rSRebFQalSTe6hrZ37UrJ7qKUf5Oh+
B2DLEdwrBmEo9Xrq4qpLMs0KSOfANKuBfEz4aFJRhWYhzWQFLcp925HDA3Q/duYx
I2XiKAteG3C07dv5ZUFL0OiwaXFXNjH+qxzhV5JnOWGbQ3rgi8ueiXzIg2BvDyRZ
kN63xO7PDMm9lFsndp5pvyJqterTPb56zdb9CUg9isgxskcyl9Yf1FUqWBOnpHFL
1BPzFCmeHFGKh/fl0jXC/ehD4BBrdbYaDB+IXuo6eKAqev72KFhp+tTK+nU/50/p
R2SPQ5SJEzbQUKNRM3Y5ZU1XIwT3az4ScaTVotw9Pq294KtywNZYI8x8B8xfyAeg
q1ur5bzCnU9AdOtB3m/5qny4At3jUaIFHcTEzv0YLPz8KlpZCox3g/M0bi/TIaEI
Urid3nQ9aQ9mooRyynFAJiaK1/FXq40ZcP6513OM1TdV1gqZxOddj9C5toNPVEAH
hhTiLqYNLaGQc2khW3Lqa9nvjjmQ+o/reT9iq2VoRe/VkgtsQFGUdel367l201BH
XES/QPpQ7n5MBisliLSZYPyA2EhiqVCng3FEzFVUveJh1k+hKWSg7FD53hkSwt/O
mCv+sKZVY+3sDQ4zYG24Q8olkAM8ESrw1FRUM9u+Ebnf4djUih9YrztZg1Ib1SXh
tmUiXITEB6TwEpTPsCEHKRnueW4X5iF1pXxy5NyHDCMsHcgX3Mo4U1ie4NGBSWHW
KCjzSxyWc0lI+Vv7rb2d7v0kMOMBYArRVqvp1QfYfZ8wOCMpXbBHHojfd+Blkn6H
fHUvlYpydx1cOt8+Umavq/t7Ifbj6Ugac0bxm+H7lpMnaFuNAfIRZ6lskKE5o+l1
s8HC4DE7WhRiaruKz5kILzlhvDQZDWj/l9g0kIewZygKn+8TZJBKpmi25MC6GbFu
5kmt7O4HbLCa65/E058mWOi9DZKyCFlhXRarwlao2RM/32+RPoRFGT1NpcjzMxW2
f4G7ineYFCIBc13MvFJxoh1CGDOguV81rb20fcQVor0k4ufRmD2nyJeLAWVT24Jg
KyRfhX15T+abOVQshiPX3wsXhVicKnxKNjmg5tky2Amhw8HgYdgvYdInlnSCuWNG
tsHMGX8t+PKW57AAPJ4gJcD1OhuP3GYk/T/ebnf71zRxbTV0WDLTaHQrYN1AvI7Q
OVQByHgpikvkqLSJoGEjn2/oXxPkFwesLYq4b8PUnUnZEnEltzIgoWt3l58zwx2E
r4+WjmUz+JpOGuRqpvDV2LpfEsVnwxD2KETJlpIenlsVUcvdoR5Ce6ABmvOKR7Hq
TnSkpDuuEL4RMERgIftJ2fUmSPxMFT9avZO8yB2u+K2xmtE0tm6l3YH5ELMwd8Mt
OA8dubHlF9sl1WNcepT2vrqDAQ0XOesaW3cuypLqA0CQKdw4kST4/O1bkxftOgyI
CWqa8cehgluDMSpXcK3sch8g26feBLU/iTptAICGKlE/zdJaF9cOJuE/NocV861j
yb7LT/orwYB2tJYjo7jQ3X7KRYc7xGR866xgBoJxisfcD0m0F538aHAzPvs8IcIW
YkBpspzkuUWbrr88wV2ySPTVPizqiPK3iAV9aDYUmeVP5VCTG6aE1bN/WNrlGzGh
R0ln+YzsXPbsu0Q5saDLq2165lrw4d5u1L4ljhARHdYgBxRlwIrX8fijSMnDTdp3
5iTukDFR+5fR4A/38Xo9fdJyBU8xrJsLZf6OvfmB8car75xLGSiEnnRxUYn9SAYf
ewT5xsxLTkAYQgEABrtLsqaOt6SH6QUejagrTMDWkqsP/QWVg5bqc9nifRQ7GZ3P
IO+W7qeNfEM7ZIsVSzLZYhCPFAD3LXG12dP1O28/DRcOsWVJJ1LIxwvGJInFoQEb
sc7/IhqHh45GENTECAI0COL4j1T01lqWj31AZ0ymZzWFpK0J4pn6y0GcaJj1P0jk
VZSFGu88VAaT+LL1SQ/0kbXTPhEE1zKfmrGd51mZ3Yw+9kIFugg65WhCr3mXNoIq
Y0/qlP+tZez66CiXP4wjLTcftvy2nXmuIZn+YSCpHpDILN3UvxC0XXAcU9amktzg
XjYYCnTVcLDwXv+9of1MzwIJGQCpBmhp2AOsCr+Hrax1YvWlBQLvmj6IM8BXbhrW
ApD6LUKRIQx2sm0PVrXro2UNt7SAK8DKAeI4QmPRRxZuphI4PfigEzSrkb7e4fLi
ppxuIK7eRx0kfvOnxFctcKNNqoLonW2y2b/ifalKF/KGKJaI11WTGjOU+srdMUWJ
lekacR83r64oP8a66bsNFJJUvIQUP4UjTiBXLavToXo4J0+mUrzs4W5PjVVbUhbU
rnd2h3Hv/7HKgm+bJFwteYouEu45XP4myLUygWWwUzNykjqGPL0ULy0Agg9GwFA7
2urXPbNyH1zTPDjKEQe5me8wsHz5AdV85PxT7q5n8hNwbXR+HG23Iy1vLxubEc3b
wHbbHa2aXO8/toGeCNjKsLB5hYu4wx/cxYjjOaD2yi2NaHaTuFnQGuut26B5vdZG
XwGk3K4AZW7NP1U1IJokXzI30uCmRKSbEZAbJeCI/9tPIZaq8UMXfh8YMM+Phzzi
raYc+80o4NFc4G2Ba5raUdbveXVSpm2r5PqmfxhRtnj0MXQ3x0kUXgxBxzUamRAe
AV6dYEhdQ6PtZWoSa7x2+GeETRL4J/tvOUuvobWArSzz1IdI5VbRcAkiXIxv3pcw
IZcarIeXWvVvAzv7LgW125qCzrc3o/EMjOYfZBauaug03PSR3nfZ/Ot4+MrDs2rx
XVw7PMjLFOTNzSBE6dBUWVaRlraxhFlqBqnxGtsME/qmE5JFWXV+bE0VLw6ghwgx
MKLo9cyknXb9+Ccy9KbJ5IvwDkxksP1Es8y9wuHZ7aJTcU1MFk++UG7+IVHTDu2u
bMR8yK8URtVQo8zOfcYwdydn00UNBgXc1CL1R1pgM94/EAN34KRF9P0gKzsp2CDQ
B74L0VtR9cHJgWixYEqk1ixaoiJWukYXAuRS7L4U9Pig8uvm6vp/JOrxaDKluvB7
Z+5wuolQ5T42QBQUoTgG35KS+JwMsUvwl6VfV3j/jUHP4gCjY0HX4ezjdrLphZF0
NIxrsbOzktUT/psKOy/+KOYjxmyY85ZtCKGqd9AH85wwRf56BUHCvp8Qjk2yK3vA
7FV75XHEvykpzLJNyS5JpozqwAfOWUMYG3USUx2VzA9vo2sG+hKmySfa9xtbuqVo
6LdV0AKAZNg+GGhBcbE/nYqm/+k4cEq0G9ug7mpPtoXVMVOKKKacsN2wFgoiAzj2
8A3iMIyAZLEDvVJSqG/sEK28yVNUbS/LZOjKPGUhofRf6RUhoWVSEus07LkYuGv6
WO4QiT0PqmGGj0nZPtUeDaPiafouoiO1Kll2MZoL+/BbFVjY8ONvcmFV9htN2V0G
KobMvOoO8lPQzN4Gq2cAfsMQ7EK0XwGvI9QNqElC4NWsnWFERib8cN/H/jYe21ZB
daDvUwDnjUe5e9i0+nAHLzuVXyfN7O1tEip98kMGgQtZrfcCC4wriE88BuO8cDRC
/0xeZFI1Rnwlk6Z57NcKMtGny1Cy+AaWQXZR976+opLyUA8oXPfYJxPkkOFP4hUy
iQ20NPnW/k3t1A02sqE3zint5JlIQGeZs6/hs0oTU8DQbvHG0gFmF6zRrqlWbX1q
E2xUKCI5doIAS17gao39usL7/IX6zB/ITNnvpHbDQ7Sofu5+jjj47DnHgeXDcbiw
NY9nXOGVchIYGazzcg4lZRxrsVGCX6uKCAp+ZhskuPLjwAyYcmYwt75NEm7fI745
QgeR3XPEcdH4wIiJrtq5+A==
`pragma protect end_protected
