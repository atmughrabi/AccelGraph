// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:01 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G+2aRwiyquBqV9MKBU7RfDNHC2SWZYoaN5ih4K4KZUVEyD95jAkcIO6Nj2V6+nel
WQZFrXvmCHYumLGln+cJJcw7f/NTjx3X8rFx3h03mKOzU7eEaSroImDVMn0t7jhg
22VWYmaQ4raHHmI/zPgXeETRoAc2OcEw75GnadKEWjA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 54032)
Ms/B7LdewnKClkJtsL6s+nGEO4cnZ9Vv+5wLhziERU0/EOOQbGDLZZpSCTMmH8Lf
Wl0xjMbcjn8qrkDzZGJvAJqnuPIw6DZBtCVgWaMflF7p7T/jn/CnEye2ZUAf4XVY
sFZyeDCx4a89+O8dk2tq3eJxDv2RUoAnnOgJ6r4yM3CjIHs6aWAnAn7nuMOI8j12
Xl8xc6XG/PJIw6pWk3YzS84o+gl/Yba4oGmG9VApg1NYbRpePqe+G8J6shxOHx7i
OTQir3i9vq2MII2oQpaHG7UEmvcJtmM/CQxRdU9QzubVnVsFRhS+lhbPecirKazP
Zyzu8IVPSkeS6eQoKYWvb8DIdj1hCP97TI2TyQqKCqgzfoo5gy1oyT02zxYpONbP
gxJiGEU34p94hNW2KCrdFEVd2xZkYCrBVL6IAG0WjlukXikEpZRu82f10qafJ+ou
AlvcP50RUMA6S9H9blk5fvc5Alu5boXcZ2SWsmbbjOP5u/kiZHRdr8im4IdhSzVv
wi8MzxzKeGJYiF8hMCPUK6exHojf9wbAOj7ZoLOK5hAQ0LCGz3TcxN9Zub5hoq7h
wMYPIf9MZtlSlzVihaZuBtcZ6ct+1Isnoe4Ll4AMckcuT77Tn84yjNopdf30lAww
UMDzUnM65ysiD1EK3la99Au9y26BAEa92YpfP1H9ptk3WqxO3cWD0/c2LkzS4RyV
ugragGTJcZtfvasgv+f3mlMw2TJUJh9woVkQFo2LuiLxdApcPXp3TMk9WAhNYRAJ
Ae0zESQDb6Af66Qou5ZEpIRIQJYs2za93UynCjXd8mYLYctewuT1AEJOCUVEgoDJ
Yd9aeX4yrwoJFVDlRgVHQ4s4pelIYim3V6iBJwthGReMYaxQ8cNFQnMDvVO8ZoFm
2XLaXSYpdJGOEvaj/pyW9qP9Dgo8XrDzolyNmR9rkg5HL8ZjoPpvQh4PalHZTPKv
/eekG+06QSd3KEEeCM/Yv3Sva4LckyVulydqKUiWYKvV9owy0ggQIQiGVNjpBP2U
iUNOIm6/KbGKXGiOxAGTy+u5Hn9Vu9+gtoS+CNOCqCRKUOLQz0BMMScRGqt49Jhc
HBLmFSeCokZKnQ9EGR4RRLh4j+NHfpXnBbjToJ47IUhh7biKZzObHflFQx0nx/Rc
KmBTh4EErAPDVdGnEVcGY+A8Oktt1IRDktEIX9h+MFWV+GMn1FG1SKYvrtDMYYDb
5UshOmNOeM1H0AMT2mor2+zeFfg3WEDEkozXp3gIN7oGjR4Ecea1JbehFSupFWQn
sRqrAzL3cAv2+A9Jz2vsG71bJshNeKBdXufRYwnRRHNmeghGzMD8D/uNQGC//8Jr
rkXsXCnf7N+vF3ehbYTG6KIruQstMZdoDPyTRIkt01USfVEu5XPLyQ43nxAG9HDv
9kDHWsfFLCIz/8JfLn1Gyy6eHOtb72vjtXXBDWFYTfK4keVpCKm5+euWXp647ntc
c6s0wn8fsYHrUmlkfl8jiuG2FfI+x+/HiXRVCJTsoKZ3JsW30Lhm1CQkAGxIEJVI
qikzBz0DUPZ3edGpDqmSBoHRfrybMpWet9zzXDxs3YrxLWlCVlZejKqBE7yzpIEO
+AHc8AKxIR0XdJY+ET6jvRvz3q1TItn4S6GJ4lbz+TNKs5BjR81642s4H66kCPMG
WMztevLHiowniLB3A5eGER1sR1F1GYJIDz7enhOwBypFQyMb13mCgk1MWovjczTM
uyWjFUAGH4stLfnJA5HtihDDx3o7SVP7nXwiHiY4Y7yr5I6eyvYn1vZJ0cubLEOL
umD44K1vkR/IFzOlMboxmK/HWjJls5hBBzmdgU60HWMkwEDaztD8osmFWiAlecyK
8/rAOWry9T7XbRgxBzrBbVIWIcmAn91TRJ5lSEaRP90I6JPZ2yhxoaKVv2R1Pvo1
LbuVGEnfTkD5d/JTvTCfXdwuTwZD5lKWrKCrWZGKHA9FruBMos1R6vgfdtZ0nAnJ
y7Ntwd2EabeyCE4nEco4Ne8bUN6i7COYKOhEKR7uAUUE+Sg9Vv0m7Itu/JskjZP5
rONRVpd/8RQm2HPeV3iL/4qLLfXD6hslG+Uq/uOoni13srTrL6sCaGhgzZGEd+Op
MdtqVMn7MfwPgbC2MIcA/+Ri2pyHn2ZryDWQ5jQuudC2uZ0bhBnS8zXfqcc0/bt5
LtZrpfy1dQndUXVcrFptVityaFKPmZ01lPwyq7AgA4hIR652/PUE8g29NJODU3L5
xPLJwuKvJ3DZr9YSxN7dh5vEW6bGxRNIovoQ57HabVoADFu4suYux2xPvASpLX49
4hWL7CfYQRcfKyhDQgb4oR8uTp//W3pA6+yiSKogDC9CWsUDUpBpik9eVvIlZqpK
5wlmvvveoAsolSb06RzjLW47QOTDqJ++7iY0CVBmuJDDp8wJtItsK22grYqXBCG3
Babdmbd+xOBFqS8cww64IFXT83/IK/DPTgK8yVFFvcfLQd9mhsyZBJ2v74Y0ILAv
ncPgIAjHkn9UQQjVrNtn2+mlanMMxmHP88KANZe7Fcs9cMFIg07X+tFWjYhcWqFo
bVIbDCh11Fmh8uWuhWmlyvYKbcgb+Vd8+M0Ds03A2jvIjGUfGOG1cGICrLbOnHem
FhCGKbySIgkW4ux4okN2hRZZ1sneZ7dPNuAUC5N4ARkqiMKdLs9QeXaVPmHiOszY
WfVQiOPxkWWpwnPuv8epup1uwxFX7TICTSiTzaWJbLm3yej6ni1aPp5Im5lFSBVV
/Rb/NgqhEsOmDGdGiispmuE8pWoZEL4Tkfmno4vcAVzJgS9SzCaUdTnKd/zfEwwU
xFfCijpA5bnMuMY14i663p9RQhS/kE2WHq7exSQcx9SaItbCNASayhYGW+E3+0Ly
LKGLTeyZMzp2GUZRn38Ch9Cj6jV6dsEf+5fGIFEmD2r0JZ8ezoA4LWr/H82XuWhn
HudrX7rUexm51PQAFMJGWejSbJGQ+DmS9c5z3lN+cdjgTwfs1oYxeoX+x/WfNqYK
JxJ89R8R+TWHL3M7iigXgnZ78WUzKKh/Evrg6zXBWANHC5064d3gRCYIkzr4ecMs
DdTOsSfmO2Q39Z5gjepPI60LIKDzQxT7c0fgn2fkpo2jLI/DSfVxGxFL8k5caJtS
2aP5JwU2s6wp2F78n5etGcl5sDYqRONxd0iUkbejma9ELJS8RBWZMzCiuZx+r9cJ
nwPBFIeh86GYhHYgdDZSehTXWjfhEJ5xTvJoWRJdOp2xZDR+taioWoAsmJIbwWmI
WA6tYEoCFe0eF2lzj1pubfpI0QSl2gyJi2p1vJLsUUOzdSiXYRt9yiZV8hMxCscN
xHmHxMZdiDzH9ahfrEt+wUTRr6gNG9KHlOGeMKZrKMfBToqwLSiftzpCoxXPVCzY
Qwsljz/oPwSuRKxRaqQKaeJI5hEfm5R/sfNQweDUPqZHaOAIFy/aUPq69yoMNwLq
6TmGy2mxYfzqsekPnNRretFuVBhHuVTM5mlyh8KnXbMMFpYq8l9CXfK9V5saeLtm
O0TExNfm42/5cxmCga28mC7/bre+TbWmasl8Jw92qJnd7MOCPhSwoJs54Dy7YbAu
dRcqlZBcMoG85hgq/bsckJ8Q1dE3/OnP5zPpObBkAdS3/lnM36jXvPJ1c/OUa0sL
aSZ2TKk+XeLkIp78vioLe6VK5cShHfa5h1yk+xC6WoBfcBVjmtVXoWWI0MiyHhwR
YPzY7rpcST5CZE4iifnveaPcX6gU+/ZVfRfQ3LagEFfrBPi2p/LarR+IwDxXEPPj
G/QJH+lQTBvk5m4gl8Lh28APkCP7ps4KCCJPMziEsq23+zHfHqSSPr6SpngZ1non
uji1s9XFQQ8NKFNPuipcyf6I2B2L2H/PXxJzTs7aqvTi2//WQs2Ud8qa+u5AZjzy
fbKk+mh8JA/cLQUwBLqYdAHKXGLivu5LUeGyKS1mpazxYnUObGs6daoqrrEM5i31
yavTfg1fV9Pjqe4yhht3Ch61MK3fYcq1zcc2gK2v++lToBFPIEdaoCaioRJyitKB
ysTgmhJJmngjQz6GIK2ko024RPt3x/0mRA/a4qiEha+He5QCuervfopTov4+nO8P
IaXtEywS23PaqscZ3Gm6zjuIaNjdPTNUuJuWzt4Axl37/saAJ+arDKnGDH8WfdVm
oSSbEtZRVn6VcaFdS7BbY9x1lw7WOgvN5Ti0d9MmlzIYwwOiu4B1FvJJjAGfjGxc
JAlV8TzdK9Ylr35Y7z43z9sHat8bAssCLASHbAowVS/eYhByZcg1lojaPldS0qte
SwqAHer7ZdtaHPJYc8Z5OWVDUXEzM/MCy9wZ8bb6utML2iQH6Y5TRfqCphR1ufd6
kSCbp8XDmPauTzEIQXZKHHxUnkN759fDURwz6jvzgwQiBM5KBgbGtS/QaaTNN93U
lNEbgiG0lGij5d8WYEpxBgV2LEI6iYHVKZfr5lG1LbRUwbjKhZ8x9Pjanc4c/JsT
Bxjl5ufzyXFf/Inq6TAO0bLPfAtBskdrOYbDnNbW2zugIYciUjMva/dECih5jOuz
3poCKqmPmwvUPK6LUNvSRewe+Ko99J35oyCJ0hSGKPUAubrKPbJgPhpciQoQnUFK
1xUsH7rr2N4jBamgS048DffqpZzJO+uWlzqmdOuyKz+G3U7aGVSTlb7WOocELW4L
a4x0s9BLp1QRvtHJszocZRYUAFwRaWOsOEUFoQ50vdTZfiE1b0+L72yjNc2dyzdz
HNAu0K9QeM1Qdv5DbK9CfTeopSMSN7vvW/ZKGwG/NePAg0zFRUj4qsfeoWotWQqO
mQt7LWLEfV3qGc4dDbXHITIGFtRxPb9jb0oCyW0MpdQmyMe+vLDvyHsWt0dsbEZk
3w4P4eIQtsjVkYcmjxVEIkAWuHEUTMK4vFcCUh/Ou93fKunbxkLJ8I9q0xv09qJr
Ms6/VXNHpldbxCOXIG0iXqCBDiEZ1GBIXo0INYlgk6bc4OpxcYIBUP7r0EIXE4FH
b/a0rPoHi0Uq4tK3eg+MAOqWoSsoMNO4cpE6cw0vlnFAKjkLybodZSS/0lBttiAh
ILgczrDA7IEAwZslk6qgWnciSJI5isk+JmQJ3pGeytFm+baAz8gMpGVqGesxcIXK
Voqaev04xkd8YcJtYifTIokX/gw1fseP2bK3dKg20TIq9RyF5lhS19scRRi18q/7
HSfA0AaT3ani29meGditwL5WsQz7ZxDLajESoLt0Li4NYgVpnQ/y+M246gHv4waT
vDRNCceVLEGNAPiYABWpms6i2DIoJCF8WDJyQWm26K+YwZSsaG8Z27f8/H7rixoO
sOgFWB2gocB+ZQBVBj7aVXGFUKCpGQCf6BodIF8yd9ETBs8xpU1QQagyHPxlFOOV
6syHw5N905Qql0OPM0scVeZSO+LnA06i2OagqKty31KGUat6siM2a/TsHItan1cn
8h8Ft8+t3G+vCGQk7SOZPAGuyqbmS3ti8e+HYVfWPZ32RdFbhAuasNhiJ6qTXtti
8IH2tSFmwqhPWt9gbQ2Ur4/wH3H2JPwzKsiws5hStHH6S+BOvCmiWAZvPyk4wdvx
4QCbuYChTGSEUQYo3MbCSkH9flAfU71bjQYbMdrRlDDTWYO8tbhw+R+HOfIUO6BI
de9pWExLmWF17H5Ow7f3ocA26qxZPAi9Rva3XssrFHW0qXfJW/+T0SlwcRnYEQKe
wTHibdibpvWLZDLXY4LvedOyFqcZp66uQ+wCfplBHD0SxNyR7wxDTvz/erQqJFvE
bqCYoQszDukVqnDMnYo4jrtpzKoekvQSqXj7Bce6UvONKlRdm4WshDjjnKXnCwIX
igwL5WbnvQcsTtIb/gE3i/4UJmT29+0jTaW9yHbz0kDdBqd23/EXpuegT4pnpK8U
7B/i7WDSbXxC4u8d+f3kRoi7ZNz6QZvA42z9azPaADEvfgZINmM9Tz80JUx1f6Vq
O7B1HLZtZTsbYa3yHMbzlM+XWU15XyMGrW4VfLQP36g2qZkeL68/LVXIcCWZlZPq
NPaZCD0K/KGa6W/ZCur0b4RLZ1ruQFhX32n/4aZOLTntMdwuZlc0pHKwIjaHp19t
+YIFslQ4uucEPXlZYT57dGbNl6kjU/z+D39zEU+AHBd1sNptbgDaK+CoZONRbsts
hSa1exaKioY5riFzMZLSSZZDrtsI8Q25bt8m153tMuaVUn+niMUkyN/qVrvbB+XA
ru9STAdU4m9I9odiZqM8SrTT2U6qpiRIfXF04WJHYGAZKdf7bNXgINWYAWV1ZA5S
dlmXoNzoYcI3bHORpB4n4636iEOHFb193iBMc5viIobQO4+fsk5BA+XUa4Tj7OZq
KTXmeo9SFIr3FJ1ydpbuNsji9OrocpqvKvKXI3PTA7nIgPLN5hjszFNMImEzfnzl
OMNymh8nGHctFg25z5ld7u8pyqL06/XScgHKUPte6GDN6mzYgJg5E+uosQgUI1/1
IZ6D07MRCHdBo5dw+xnswfOKQRODpj58mTMrDKv7p86wEp98f9eS6/3z4tcrSqn7
NyIoviXT3QnDwfYJH7OXO5rRFeMWeLPtH2PrEDUWE2QU1GDnV40Bhpv7Pr8SF4dW
zgIayu7ea+/I9PKdML3hiCK6kb6zfpFqtt52piwcljovV4NHVduMkJbB3Nh0Wlwc
O7Wz3tcDJkWqQpY2kFNSjivGamZD9oIrbCy0du+KSsmTZimfdOX7QTASh4azlwpP
VwWjnRB1lhvWTx7UhtmoRWh5I0EGwkGn+wka6+FsUPchlnvAenoKvvJqD4r3f4du
fBKSN40JDOiEk/Zbtjid4BriPuL67P/9K5MD2yePSl7pJvruhMEB4BCESaOySRxm
ren0nZSE/e5e7zLP+Zr9d8CUck+h4XJ7ypqDw2EXBii6UTFg7WbaRbQPOJvsAozd
N4m1udaXT0Ba8YrF80wfbxR80M/ZDbcNrdAbH5Z2dP96YptPxZ0xb4FBUExkAr7D
/XG6j9gsdAmmDE+IP87QNl14QoLmNo+QoUAstaD86fvKQi4zQbrdtsyFJDqBNFjH
5KLF3Uil9v3OTpAqfYZUgZDb4uZpMJefinII2jPpa5nIEPjTvqEucfpkuswF/zN3
iJ0hjsKf70TyCacXSs3zNpszw/xnWfeayufeRGupaZn3//9g2piFUXedUgnNggcJ
gqpfGFMhpROgCwefPsEn4hqzBi0+MbLdPE0kIFQuS2oN8kIRmtTIARemwCl67Mi/
eChF1nKNij4qCy35wrMF01cJrUnf/9sJUWzespzzqIoqh1UaycTf7l3AOP30MA0T
ulSkAW3HOMtESTytvtcrePThdVuMu4/6fl0u7Y5/lva2ICx7KIfHOm/BGHfmgUCY
YDVH/5hzY21d7B+qiEjP8n1+UlSkzzq78+Hkh4QJkGwtbyY780OtfKDn10/9Z5HP
TLOlYJtmKYZSjfY9K4L5vOWoOG6R5qfgiB5TbwlSZu5d74q/kGRtr+D3F3j8NF5e
LCfQdklNPpNibOpJMk39KHWy0dzKzDKYISFTxdOHEudWQqcGNQTSrRU/UXFDe8VX
NK79e4dKI3dU+o6R+jeAeSvvpOvsE9rGEtRzB48EiRMZu9hKaWale3jNzA+uRU1c
B2vIv2dz0QKEbmVpJE6Pa/m9ndsJPmG8SYZGpZ0uCNFQR53QtRYi9PeTV17f/fTX
OVk/Ce2gOzr3r3+EQAi748z7/w5lAvI/u0b3wltq7Fr6JAwcVBrkSbtGcuBRK7j7
0u7M2Zd725M7mCFRU1miiPhEMrJP7U/spVRwvRwDf03HJhSrtDXK87d1edATMbFS
NfWuaG243DpO18T1PwYMGBOzpJhcQIq3jNeV5TofLkg9la8VfuMFMvOH4XYNwIDx
o/VrXDDP8ePhTcpYlwsLROSMRWMmfuLwA+J7NmJY4Z/OwtGm4HNWbKgrovuf8h8I
E1OYCneodUDZUNJVtPH/zp2xYh0Af1nF+vz2lP6eeB+GLUF5zHFdZ/MxZcCiJpan
kB6WJqUnnYGYWTyxd06FpZvRsmBqsM7juAfK4wKxrvbjqPXSqD753FlHOXneZwk9
CuHwdDUo/6mDuJndosP/jXOwjhsDEEUYsLD7C7bQI8ay1AJKKhqBsNN2qlPsrO+Q
PwPk9mdsvIKtBr9DTTdHdFsyIQmXb41ASyXuRZmxjI4p+FLUSkTLex2x3iXndFwS
FvAsnRwuprxF1beQQFiysSQQ/brM5JKbowLM9lBXH2GM+2roCrqJ6j/Ey/hKLnaV
0AJD65bDtb0UInKJBk4s9bewPe8O5eU+245i837LVV0B4Yu6WQu5rKftABujFhDF
N1jvEXxwuhqhLcJsj6NXU9W4WQf+j4rScMsJa8vBMg4usmyiIg+M8Jsd0yXXhVOS
FXvRMi7QRfno1DJ/3DxlEg4l8Zj5KOFRAYVgBcd2bu7jRu83unBnktfboXS2PrS1
6YeHzgFQKpeuXOJQBsbHeJv9S9T2cPAMlNfvCzRB7+62WW2wSPZTbJ4bA6jDpaV3
2puz5JvsR0TfiYLNx9tAFZZOb+HZCKT+WG1wH2msDQv+6aCiv8F955ySnCdS5hlF
MGN7Km4C+MEuVwIWbnBSS3NgMXVFAPqFZN293rcsNrdqzuMVZlcdJQCKoANrti4z
XVKtBjYJW6KRtJvxMXRzAx9E0wayot6OlysztF47qxnMuiDWa0jCWOU7DfBC0j1g
AB07fUKCcD/dFQCg2o6oR9ET4yBxyVOBa3jCUdN9XaJmAIP7DdEHGR/LI7V8qRx5
iN+Nb2/S7TZw5FHcEpsLve3fGREsHkWRy/Ch/rIhcVEQgQEsDHwgeOGYPpGGUJOR
BPh4b07AwSJRnjrol/bUCSlgoc2qVmBwJQ6DoINyxbPehgwzJsbfkLsrD9kP6LXq
I8MPUimQKR2JE5/kt5UKtVgju2kKV+Q0gJxybR+f567jIKr6PGtNnhrDqS9ozD4D
jrSKHJrPkoapW38d82s7qILSoTlVss3mHFTcqVB1rFR9MYLpctHij/BHtRcR7R+G
akoWWhQSkNgxq3ofAi+yzVcq79NFrG8jXEE/HPtyUrvO1wfdRDmzwnlyFsNSINWe
z4FoipqOE0Vr9xbcHhqKYI0wRfm13wL5U8B2+7qKFLBV8skq3BQJFQV1cQ2O4LtY
lcShJIwlSYIi4TPvq+qrJ7TSPx9Ja1Qv42RRei9nS7qA+F/yDJV4xXgHAr6acdyw
Q2ZpE33StCqFqMZyFjKd4Fm5csDR2dH1wz4/rIWgDcg4Vr8lcXg/QXhvO4M8ln5k
A/elMJyNMcbdEImeAVHwyEgvVpSso+kcVwLCdj4zZTUrniXBCiOcvEWeO3RBoTXa
Vzk0tgI5LDbodm4zuwWDscjgVgSyOKxfP7LkPVATDq9H3kyFNP0yAGK8vbK/77FE
HMMJhtIoKzfXsLbpYmz1W1pwJHToFwFUW4r4Rdf8g8yd9MjQ+pCbmchjugq81K2V
7fNFRIpiqL/i5e9ZRRjSc2AqYRiaDx7swyKaR6WluApLLVVXKDEynhLfnhMxk4ba
lDeX1msRtZP1x90myogF/+HnA1ZnfX7i+ZkzInPxruAovNfOy7KGEuWxSmFl/zCi
wjZFET53OjGJO7yu6PtX49nG4hYlEv9Hstl3Ge7HuBmfuAYKbyvpAH6xRwVn8JMW
A29zNnHlTGksj9HfYTmcelRYDrlsFXX8/fFl9Kez9dEtg9iZN/aGn3JEJRdmtzKe
gVzPUD6dMv+4HmHIlwvnFcjcTlcGRFoUWtBes710+ZSoVDNCboLlV0HbHUPhSgiq
NFp1Rq/YvSnjGE5mVBTiMHij4eoQr3GHEhvhW8XIczeeo3GqUit3iwGZkxDxE+zm
79jTfYlNCowu6VJpIXVdoHP3jhtMqDw/a63cWny1ywE401Oujr9dww/xnLykStns
5IDmjpkbC+U5s3exBhuZo1dpfPFjD/tQyQgmlYLxEBxSGGrr9+JrFI7+EqddFTot
z3kwGrcbfLIXtxD83ecWMFDLXW3SSovTUjMAG6O2udJ1UKUBj8kByvE3ghzcm4IS
vqc5obnxk4n2n5u6BceOP7PuQHcerHLSX7Dq4xklwt9yd8y5GGf8DwsnOI0sMSWS
K/WjS71nh9KSLBiHtOPBbxEOrdpo9iObPTdnZxXsJzi9u2e4A9SgWAnSQRRrR2Gw
qnKI1x0N73DXHJjdAyPcPVVbumlXTV7VDVD4Sart+dMKOC0I2hA6is3iiFY34lIi
3wE7KOi1GqC5yaGXkGws+NwrtYwLyRPJ/XF7T2hdcEQMYIKQ298hVs2NkF7sL015
k+D7sOj5idlgZuwyZpSNhhQlbo4vQIPtqiwn/X5Bi07LvElF/qeEeGqotMeOWpKN
0/KM9TyBViARG8BtHCW5gSbJnGl4TDDW/ZBY2+ei8OrRTKBFw2X4Fw2CJjZn/QHL
gL4NOlIvoIjxCxLxuIyQiG4wR9e7OewwsXJPypST+CK28xt1o5UxRNwHG3jfF9wc
t4Yr0CBJQS5slbLt/CA79Fe4a+lT53F3naFl1zc992hqp4WE9RUcPZIjkmxct7Er
NoF7f3ARJgNydCApKwlkRHxlrrSF3BWc71nWG5hPv9Tgx9lOJfIJ1Bwt5VboVVA5
Bv0l/VHhMv2qETD92CR46tRFhOUkuR729hVk0nuc1kvmiN2ixA7q43Ut48dlUfPz
k360LLT9NmaEdDJnzO3l0KMyEtlXUtK/jGfJMy+hynVhGYMgL8p+eimIw1TUIiOx
5D2sQnXg9aCVforeasSmB+T8OzqFI2t6OkQNDTY5LUKe/VEZISnqqoLKjg8Fx7Wr
urkX0LhjBOGE9YKM/k24C/jJ4phZOAM5ZrgmjufSKjTyggJEQHurCUiGQ/eSzeUc
1gCQmsOjuTg3V0QblfQzlbdrpYMxE7M88kuVDR3845Aty40xhA8OI7nPkiXO9ovY
GzueCcv30UaCjqnGtHqyIkmum2IP4SPnD0b5ji2JfCJlE+hNGIs6oJkQfHSUZ8/N
if/1fBtMERZ2GW3Kio0QsOSUZV1F6UPjcrQmsKN/TEmZ7DeurlSAoKD5KjtqHV+y
JYFGpKMrLZs2BEqF1TEVBEVGfIwgiltTr29VWKSyzQ/XWrlQEZwhOFw4hQYFTzXR
Z/+aT6DCu4vVFZycPDNqX2BdcezoKP/hgQilwM6HIaPjQGiI1SCiIR2XApYtwliN
LT3oGnUanfnFQHgsVd1ScyuI3ZNPfxFB5SJOT0GhChaycFt/b4zEnYejkUkYAjoL
3SKkKc9wrrcSWI7ujyrN/AiiuAo4chrhBo79+V9GUL8PeGUvvl06QZ1QkFD6lOJ4
o8dNOKFdZwvV3MMWWCKhUObSqrQLQ20jwfgNxlIlWixIkFEeXV+7GvKpeBRVq9G/
Cn/oK1WVARrEIIUMOfPoV5Q+EClFz8oQBKvC1GU3AMEihKyWcYwEkNxX8bBiOV8Y
4oYywpmMOsqv1Kxuh21qOst9PAJAZq3mDBCVtLBNGI7C31KtyRzMMUUSwcfkuF0b
rlXo7oszKdmwOEcrnkpWviHmS3KDdpCX2khI1x8uTHGyLNu7mjulz7ds3zA7ktvL
K/fRvItOfV0bPBZOgO/hikJWSQpMvQWNNzg4IrxaL9YgXWFtKSTaH06rEirwVjX0
M8Wx/nwFZIAi6Y/Ybz6a5oyRhlzjH7BNB2VduL1BEw6yyks3GLV/Jnm72z+K5zdN
263ybktmcziUDHcaF3vDhIEPzU+BZfMDsjLYU3XQyWRSdmioWxIBH904RlPAbnfF
W+G6si3fwmxBC5SMQIOFUGQFalz9vpgYbnRvDmlhl8HiMWy7kgMGAxLKIiEqvwZk
O1oNQgFNn0LUG042XKCmHO+24kSEeBFGMyg/8mEYGHNCUkqiVPMfeksB300G0QeA
VTyseM1Wdom/yDemhFBz97Xw7VudKh1oladZHHq3g2LlIenIVf0PVZnyBqtgR8+u
Igp97RZLTh+Uig78Bvi6jFtVFCga6U4KvkDtij755rAAzORUxt2x9WHvchEhUTC/
/DccNuXUJYO7vcmFFGnEzbN96iq6kCi0Y5sGy1IWPp14y4PhfPrh6T1nn7z0bdX/
FeY5EVT2GCWDf5g+K1UPUQ6iTsoTUhZEE0LSTV+vlRc0J0BJ4IIxYOUTcgL6kwmt
mtaL3Eoy0IBXjT5p5oz99EStx9kveC5oANVjYT/qe0j+l+6djfIwJVl2yDCE/FNS
HSZ4lMfm2VIc7GSk/4G7quO9MkPnQElH13Yq5ecVD+qqtizuDEYrTqme07WaWOe8
ZqnwdsxmQrdRKmIiHFEoPJqaOl3vITlIwQfdePA0ea9f67MAwB0vHhpX2KWAs+xU
19qgNTrwJ7NYfzFBVa2RCjYao1VNm00LDrV0xLm1KiW9rDD0BBe6eRXJSJwWE/EB
9W0MATY7P1vYnWx8NI4zsKeJKa/AvEb/NSVSEpFQWE2vUuYQfGV5s1SV3sNH8wJh
E3XcwCzoLrf7ik2JxBeCFcvyvC+MjRRWcDSmr8t8D5WoeaQbe/pIwM9pXjDvSTVo
uD23nZtk8FvbinofDaie7svfDvNWasRodKsMI8xWY1jgmnre40sM89bcbg1fut9f
2ZbZnajqEa0KkC75q9VMFK/NjM1ZG58MaV73vzULoNEG8qYb6QkXiieT0s400n1r
zMH0s4cMGFe8MRlvac3mnFx+RxNM8CG3Fbs811qlxCuQf8olBiN6ei0es2dTIuHt
66NvuPHuEDuONLtLr1D3bK3xXbpUMcj52d+PHSfj5OsuZNqoe36QIoafenuIacNX
wHOs4dvIF+pRl7NqYgi68kQcluDGG8RRJMm2tbPJGEmyhcXIQzbE1VTe902U0lFP
L82Fnu3jCHyRQtGIGlDVumGCWINo0qGHCAx5JlTKsepinh5YiaJmx2cUVT1VVt/J
xbTxgeJBDVCfJdRqR20RmWWOa+imMaFYuBMTMcFwNzIG4o8KEl6KGVP/2HMWhmJs
btLVUPmFgGEab3Us2fYKVCoSrFwWxSWfjlGojnPaZE3Q64yEzuV9g9BZjVt9YD8k
J3NDDdDPHGsAVr/caQ0YI80hzhNhihNOuNdT4CjVv5e6frnZfmE8O5dAFch3RYjm
YQCza+nBPkXsAMX+wK+QSZxhW2uVzNEknlheL72LOBHfTYBz2UMXZ5u/nlS1LJeO
qPjblIg7fgWUMXDREqZ/duEdbqsLHlEeJGebSVDEg87OhYwZh+41dkgk5wW4g59s
cFurvMgHIfZzQ12MuTrgMFW0wGsKNzPUztav1tfSYZvNRkoU6zRJ3S+uObwi0zjq
dyBTzPbA1s5ac9iWCzywrLQpttV1tH0WiiajP42OeEuIcW7HD/wR93tkbGqp/0sv
961cESRrl/nD0B0+kwHWvXgamt3zYJwYbPSX8xSRBAvoLAKg7nS33w3QcfyoCf0T
r6pvR6eJet6+sUeDTCXOfghsDg/ceJfI46XhMAo1cbvVduQE7fI1djzENkTVmdAC
tOGD2DFtPw1UDecVrFPLCrk+fPgrCnPoJJoHZd7FN7bN4WT/e3I3uT58+pHLCGgt
numOc7+NDyCxpUdCKzrL+b/P9X4F+XUFBVXuXChY3OlyJzefS6Dj62kS5DBxryEB
QbNWEyVEuq3StD0j5g0+BNM3kYmA+ACeZAbgqY84uKGFHPHKFKDiDtI/9GH6UZ82
vltIQ0L74tpD5F+jbWuP02C09LMVLE3yvtcmHo9CWVQdHwWoeq5kxK9cS1NEks+p
C8F2g5wF42Nmx438/HAosOLvK0PFZGq4loBrgqmFCjxnj6Tw3n8uebz8mpt8UCO9
bddNuUJpbA1ftInnuOpNDeqHsCu+4jgpQuClDbTWlcqTbGiOsvs199yk+5O0mFRO
sRluOaXeWvj+BYycEqvURxohmamZ3bHaSU1yUWMToT6pWcRriRDYDdQoBWJSCyqJ
shUPq74iPkMEJD99Sm3+DngHAQopjB6uRbfxEn04bjKJN7bhk8uRDIFO0tl9YkIf
zE0gVEXfwyC9cK3+2Bfn+oAkcbP+AsZynP1RApqXLLbyJYQdAsqck2A/BEeoTgvc
NHQ8UOtbuhgP0b4fHdl3OPfizr2gbvAiD582ZHOsHidfgcbD8TWmA+vIHkgNyCjk
wvt/HMurM1u4UfjpcwK4RzLwgxBJsGXm4j56wsXcfPN+UtVxMrXSTUfh4OGWVvpo
zzbHswmNZ8HilxIyPTDwDtPjhyGSwHxhoAhLj9Mx0iP0T85SSv9ghZ7fsq652dzZ
xqjc0TN6wIugpGKnWXZKRKDr+ZaZQkFw6S0oHQ2IzP+07ksrGIhvKfgJCwxYPfBa
oRFzoH4XzMX9yBn+Fp5ejriIFrg4o3tgHPqK+rKWr2zRCbGU1M9gG1EJTp++SMib
LKEe8ZCEho+WszLOE4pHfFn9nQGHfn3YtgN+gHVqDdaMSwALj5RuMMAIUBG7QFXZ
hKzKSnp8Tb0AM0mZKXLfl4v6ag4020QfekbaHt6PW+M18RpWwIMG8tl8UrC8QQp0
+EIT7yWx2WSNNbwpEX+aVTGweCyFttlZ2ZMUpIuzUtRgLzCKAPJaMkYjp4m0zYjT
lhUHJ9QDiL/hlgs1NEGvJA8WeP6A5lHrLCeNd2R6Ym3l7nFlxbRgSgQxICM7lsKx
//rQd/5c3vOdguy4OSdaBCBQQD/Ze2A8NQ/ag1znR9t4UoKvyamX+Ibdn4+T2oNz
s0nhlEmlqWT0YZZhM46BKGLy5oH8dXqKzyQ2fMNrdZ+aV6nQqETc1TUixoOsIWbP
9gazk8j9DsgOoStVZq7Yf6DZVSpaFTJO1gKzmxaVIzSMqwOAA+sI8NqenBD0NNRG
Ekwb/YvuTX+WTITshBd5IITotewWGfU6MrN9nXjenl+A6Spy/N92wqrmVskb/3pL
A95ggXkZB97dejDqUAXv6/3gnG18HO33KXTVUH2ahCwbSQsRHYaYRJQYELsab7xe
5vKjpH2eBdwIpHAtV2D5vF/mss2IXwrzzGZzS/Gi6QrJyFp4batZ+CrioV9yyQqK
HB5hOIcqsUFyIJ1smpTkO7NlnsftABvCIRlib0IAG02Iep1a0VLYGdB9cGIisxfd
qFb76LfyEhLerb2XqAWwGvKDitn3NeckKtlNThKdkECtlcfmKP3DenAVJiuwpF06
ZH4L2JL/54W4stEWYV61zkXCgwpmBjXOel/bHWnfGPZ7ddr1J+WWEjeIAv4jHYRl
b+kf/D8JDLyPGk0hXHjU9AqCI00rLnKVvzmcU+82I0cyVkh9YQuHRMBmuH7IC8KA
sF4/LNw4Qp+znNPBfW63/DeTUJEZlzDVHPYT6hfTKed0SkNTicL2gb3hw3F2ONUC
einss0qwnRDAJA/JSjQGhF5CoOJ7WXvekaHuUrUCKHeC6+wFXbYjphxeKoN6IPU4
WUI476toryS+OKImjQsaVq+AoUiP1RroLGP2Yv5QEq/ldwoQwfEGXBpZKAaSP4RD
KgUsdmbObYPHd6pIhHD94ICEB0D/d7P4xoH0XZflvKbTE8DszOK+sTltgRFJwtZK
cndcsbatT4n0fC9hWUs0mlc/4k4tS/IbucBP+VjAmWJ8F1St3RtJ2YC3OjswOyib
RQNqauoHSBVBnIs3odCBkv/VV/BunrBP5sjbnStEm7MbKdfbB1jhpJww79XsSm5q
se5u9XBana2H4hxm9y/3ZJs9HwTGcRte+JsoiDqC+4M0bAm9Rv8WnrZhDUiitZIM
AJjn+QTzAr2HFaSviw5X7Cz/cXb0QJ37d6fYntei5uhb16FNcT4ec++N9/Tupl5p
m5FC1aYwNPSRRApo4b4Gyzq6D51pn57HeVVP2NwIq3/fEh6m2kC57dp2tyHTiPCK
UGToqRvAWS/uCbQXTYWF1Jgr88kzomSIgj3+9dMOMctbAoFGtaPDFTsDDiqCSIO+
qsLBxoMoknWzb1Ty0G/6FBkgM4F9eNWyz69jPmNAyv96e9rMpYthopOjF6ydktz5
sXP4sGgO1mFeY3JDMHXozyiIAY/DknAJUoW+Vm9gfgiUUtjXzUyYktbRjHzfAz02
4CVjBjh9cbo8gf7WT4QurallhehA58/B9T/cODRJyJuQqR2dk+8eeQYRas8wbdDf
VdzLGMEvv9MV9IuDYwvCZwVo1OZzti1CWfbPdzisFE3V9qwtWWmZ/41X8Ii6ViIi
tlu39t1GA3kQ5vasVcCsH0HAqyywLfJjlUxrQd2eMNLdAStjMlSgnQ/9lkFkvD85
0iUXw/vpZchTA0A9FASZcwtQS0yfE3xruRw5CYbWTp0Luie0zj4vV440gDkxNUBV
SnRHE+BXkdQKf52naYQgbYL8faPEPbiYGDa6Rbi0pRKeMysagujUcXXgSmyqMVxS
an5D76KOdCFfjmjy2mcUa/ojBdUGFFtrWmwseAmDumowe070B+97RyYlTpoeFBjs
AzsgAEmpvPS6wEtBSpn6KsXZbmXcLYDTBGcYA5Kgxs6ktVgi/UR5OQmfCEPv1Za4
kKHiz6SdDGd6bvzZBegI9+ZhnjtNcKkUN8wb+D0P6s5bWHnb7TIGbv3939UF7RSD
euHFsGkkdC0euJtnBaD3Obf5K2UfSBfyPjs+x/H4ASP67apMUkiMIDHbJ5Oygtqv
tS/JsaVNiSwHq60P5ujCE50I0m0b8uVLEQCFl9GA28/v2Y0KSkChho1iirLjswDt
3NU4A6pVLiMOirmjZy9HQBAIZghVgqxygbTUn38bB1bOavbmkQ3tLKArilL3kQbn
xYxlFw4Tkh9u/y4L5x05whzwuKnEe4+uwXeJFBWZVfxbkCMS9svTchv1yBzNIklN
AGAmw/pSCmqYdjv+2tqAkBATJlQh/s99vHTccCQk48uU4vzsmANqnQu+j94y/A0M
qQsJhnnfj2BUF8GCLIElW4H/1GVaa+j/lhGYMtPPv+GsT9rq95XI+HdNhaeN0pou
PTqxh4XX/blC/8+wKkVte16S6/gMINxWoJaGmUWpBtwSQAy19nETtKq79+Wuok8F
VtHMn+gWfwSfIK8LJgQCkWkFf/10oth2xXzXi6cQaX5Kbu4meCQx4rNgLHkdBJfM
+eLWzw1nvSJfUnnd+8NniLgM+vcRbJtO9kuB0QFOmSMvH0XnDjonfskHRcLpX5cC
yyZvUjOmSiOs2EPB5t6Yrtt8txCbq/Y2M91KYcg1NRKYkiqmZxwtNj877TEqH+D3
VT2n1f1vdzeS+zMaTeRst3ao7Yoof4xHhzUYkc8pVKAK+jNL32XwvFulLOaLSbgn
uxxy1AuXI2nZ4w159YMv9lDmVxsVshinGloda6u6wf/8ivGZO4slIys20KZjyetV
0OWyBOI7ktT49nbujRKDBX/CAOXEnWvGZn6NqEf7OmC4sDMNGjWAjFGjYM0VFl+j
/a9u/Juq/JfGdjHtYHu1cDeJMe8bw34/M7ZePrhIhQpz46WQM/4N/ZdQGpzojQON
ICYE6viENZMS8EFZoHUYzlr5JGMQ24pMyk6D2UfbVL5L6IS12ZkGP0BnmEUAjB/M
W27MXmXrBi+6b4t2t7TmgXGVsTNyVirvxwcwcJoa6GIde6J3E+2GHyhF8WtcsiOH
C2oe/+/tRXDa+q7wHpuWePzKW3pC8ExTSAbqO6yIwoYpFrrsFYfnDZv9ai6Vb2L7
MKdNXJ7hZWKUWaS4rqIFZLFWx8TrZZd1sIIhlin17wtF3SopFCzjCEkt1I+tehwt
zO1R0zmDc+j+BwIP44ndiCgX0rPYN9tHdlRi8bxP2gRSfDFWbewUaWRR4OR2lQ0s
Hy+XcFYcpl+KEK4P9ZdwwLCb5KdAlcaNlXf2B9Z81OhPhG7FcByhdQk+3tOih0EN
/Fyv9Bji0t8NpofnCgLS6dHqD0oxbgVYlz/Apzc0oCfeF4bxidcnkLgCvxPafwe7
0JFm9iMyn9ma7vzyvU+E4ddLWtWXijcpMDJ0/1m1MP0mn+5M5dJgEmTkzkiRoez+
NpxcRCuaw+UAlTIofT7uc1CmQ0RHiCno5RL7zHjFJPaO285IaaXCb0BXd+v9SRIh
XNDJuKYIkker3AuJFFV+Dphoxo9udUImEApPVY+LoS1coSXQJzvMV/cxl2R5LjaI
KWkrLPILHKIm7j5eAQFDHQ9gQsL7ioMtbi2zLwLFNuvjQ0BcEjqNsVSFZMgvWs5A
THi4ZjI/8uRgoYmW/BPJexxk97AZfiZAcXVVR7nqXGv18gIBDGfBcNtPJLpP/zKv
3ABHAArqOBENBL7xUpukHJPa98dwdViHSoECxBthGwC2NoQ/KWNUx6Ec6+Z+9oFW
ATjsa53NR/LZtC7Ar9TjUHyCOWhNcx/KVxOok5Bi/n2pCVTZcJjOWMpGC33qyDwO
SDEebnIzMGHH1QLCgmSyBMDaLjgA+6G4yLXClGEJCYIl2g18JtvfKbBpYfLJ99zt
l3jQwIsyK5Az/jA7s7Pl0WtZLZSQ5GVU3lpJ/k40Qt2ulJBzeRpTrThgCl4cNCo3
hD8w5ipCZEM5bxJ/jIJQxrTD0YgxcZNsKwfEEO/aetFbPHBl38l+Q5Voen3D2t05
eLnKFo/nRrFvkO8rWwVaSBAqiS6v3g/Li413j1BtYM7lzAq1GY3SDTdG2rPS7q2Y
udgmKuTfv7JXj67+KvOPuE7J5P/0CMmKnHTIxfa/YgQODvHu1/AX8VHp6HpTPfu1
aHl0YxhLfekNvCJPPV1k/jLX473EFs+MUhY5/IkSFvSongcIWeu0Lvukb7jowxeL
iGHTcKvmRcNHfH1mI5gyA8rBQZvP6wHgwZ+gMGWXf9M/T9n64GxqJU5KoGp4Dxbg
WraFono+xq7YRSMVjmbRwEQ/yKuW/LQSs4B8VSbANIn8HUgLfu/wjEAtkrQiEbB+
/jKozcYgTgGMj29vyCkrGW3VJPuXNpm4ugKuEVhkUJ3/BbiwvgUP6rRP/5pNkP3T
yGZV0rjVwMQpcW24tCqGylwyize/LLIaV7SsWkJQGv+7XREBlSwurwKjwNhtDxWv
RmdBfhDC3UQ6a9/B4CmWvPLO/KFAmbK25QDNYdTvbtjkCt7PmrvBQ4opUbBPm+0W
PBj5Foco5x9U4xYKkZKODlYVQoZUjIwc/23VbsMDLiKmhyk3yZ2H0U/ktL//0Hgc
T96fDbeQGFNqPHJ6+WxyhMtlTXoEdkpah4krILI+o9k9XvWWur+cKNz+oK6O3twf
G3Wd/EcZn12DDCVDdj+1WZPG7aZXtUF239ZEpBMlOycS09KEr5huAArZsKzhxk4S
TTlSwz9qZ5LFpa6dhZP8Vdr2Z95KFlOX4rgryBHtNSqnLJcJ/rkVuOO6GJM/DkfX
rce52MauM1It/ATuI4us0OX87sztePHBbk3fDYI00vOca4ib2sXOCCuQgDjhReOB
KsKHrLx6p47rIPQcZsvVCq4eCL2l42CvKVQGN3strNAuNWnQ5lmzATcAhbOZxTNt
R9+F5nwSZsQ8cbNKB0Bwo1WD458yIsj7vNN5qiwEKELVTgmoqYRWgKncOkZxRTcb
WsOJaOmsy3FrlqWSpVpc0PV7qh5KsutPw+q2V02RjD4C6qEogfJa8T6/b26E+gQ/
XnFFoh3ySuYVL3nGL89tAcGW3uJE67NbqD2bNvhSKPltkHGqB0VttpNndHB6oq9u
0jvglv6UqigJH0CSidBplOVlodmX7WYnCrwijj3dA1k2P/R11ChZvFgx48KN4fqm
t6o6k+Zf/CqeakQPBOAfXonNH5GIkWgZORY2HAiII9UeRQYQch5kntV2nBnGsvNT
5ZrGRPhmah5yexcKwlEaTsDzQ8uLrh7B1X5gTFa0cGua4leZTfXnR+D7MvgbPF0D
FxMX9BCj0vCiqoYPs1I/Z1iE3zbeQNrsqZM0R90rsmU3pPTPG9LPRUbyMs17ByLZ
4CeRxzGPQD/tWwZ6cIS3CYySGqh66nAUrSvhJzhjt++u2TevXOgpbm4u2N4etzJw
VctnC8BqxQ8/wDCrcKI+ohx19NxTF/tmG0dmgMos3n6zK7p29KGUvvsmKwLQc2vf
hM92YPh7MFlx/KlSDSSFhR/NNHFjffbtQn4tHzburCFqGhF0c1krBl7+eF1sdEre
2iM2mVkI1GQw18XN7ylnTJvjIampioPL592TtEgI8V+RYwLR2Ao8to4eRXfm8uLJ
JKZgQlVjBiu3T074b587Bsi6i8yHZuzT3RwFtx0SJJH7PqbMga7Qc1KvFcJ3a5hR
llZ4lIGllDr12S9iOrAeaXjVk3YZV0b9WjbIGCaH7MrEJY46IcoMLsy3wSezPMig
7kqj0VQxw1Q26E/IUKiZejV59dHf1M+dYrvK4MyjG/irSwde7FmMylEw5LnPdbYe
PY9C5jDOGfAlmfMQgTsqXwWXlpV2wxF/fzb6r6Zaovq9PUSvxYMh9D9WLBcJWzEG
JqayCZUWLHgi9DzswZSY9mweW6bpqrHFaSDbjxBUHTkpnm22Tnbmzma58pg2OH/2
WTRhyfocV+gzNZv9L75ZiDIpRMmMYfXX+N4YINRNwgHlUwuJm7TonDJE91GwuoRW
zi9xAtKg7E5kxMXO9sOumcB7VWAfgq86GYL4Pkmq6cJv5+5klgrrB/2YkzYZFOur
QUZfB0v0N3i6FMoa20lor1DLVj+6mQKCYCV0kbfBX/b7rtDrBXFDEFu9fU+WQp6E
/mod89Pf3sxYHnjhNiDCE8wk6UM8qmqovAhUOKxnXZTIHfV4h8P4HnmkTVfbGzyB
K6t7JiEUcRhiJ7fkup2vXDG8JssbydMUvXBKLuEqwKPMnsl047jeNy0B2qavdgIP
XdlcBNvSGQ5NzyfnQ8a9TDad/5b9epPs+HloagSIW5mx265eZJ6mBnqM4eBsszbD
cXT0xuJoqVUYHKAaVGSCsfyo2M8iobYJn1avW30SGDlMx1IWsLLPnDE2LjPsGBU/
bhv9/aHewFcZvMS+d+WiL+mYjCFDMfCK52Z0xi9ZvvFv4YNkzMdPD6lyZbCaG1+B
CGe2UkaOowWALIyWVNB35rxK8j7grolEbYUeqawrnObEWhw3V8f6Is1n5jhhe3/9
SxqWnV50BSfWtpTAZmwTnqZkw3ilcy/Zp6Bf4Nfpo5zsqTLE7Ua6/7eEXxaDdqgx
IOdF4rws1IGLKqxoQzrBrZbjo9bj5giBZ71oInXsVp6dJzOJ3QB4sY6iSfYFOsJS
PkZG6VMFYeR3tvgP0BLR2nwi1pBDA1hc34iqsjMjSlPOYNusl5nzGnaMI6mG5pSY
SB6fbZ8BSNEUyiJ9g2l9EIdvdTfjrvpKHTuHX0ft33iapvx0y7fPkB/t4a75pqEH
H//O4mErqN6j2mJFVS45QPFBp64uMpSpduXjXh/3on7s8bierOVAizO9Uh6/GL1e
wkl2GyMyz8ulkGbx4Ad52/4bwIXQs6OplnmpKV3VGqQGsXEQuYrQ+QKuRRZhcITc
i00t04UYBrVSzgXDStqtWMIw7Z2IsmdXw8wefWs/54KIvA0rI44nqdsqX3P9k/T9
H79zbkijIUCxTM2iCaf0drR2Vq6TVRLs7ZUNI2hxLjG8OEJB+7eLKiY4gnt7yhi8
Hga1WJZ+anRaJlMHTqhD872HifnXh2waYMDp+mpLTO9fu3xhsxeu1RMe+0NjZ1gT
uMLaE8rFHQUcGgQFgpEyUdanUlvWU6u+btKY46Wo0RTpVb8Gzt/V1544gmi3eE+z
V5CGq0f4qd7EqIpAMOn55Jg7RXu96OuyPJ8T6emN+CsU0yrQV82719dWxLN2HTJp
rwF1edjz3UKkO2Hcy6GuO1f6fICM+g7slAc2kUyo7b8noAC7OcwRlRbD2Gf69/Et
a/25l6SV/Eqdgc6MX+6HdaJG2RaqHP97oUtGI74D7r12Yvl8WHegyvIaVIXFRm7S
kfvNiWzZPIrZ4k/K+eH/U31ckMsI7PtVitlymMqNDk00Guq7HwyW1L0DJuWfmr5K
+KTtTIoZoZZLdh6NFdzrvGFrwAMW29wi0JfxH8uO0yw9ZESPWgCdyC3G4DBNB9Xe
gqZic/SzirjaiXIgcBnrckAJU47I/9ThmJdEXQbQbMgW/BygmYM9FFa63/q/m4Zb
cf5502/JGdlxHC+AGpVhMNXSYz5yK/mPMCsDA/z9FZ2fDqkrvWTAuRPWJFcmniXR
z/aZxBMsFF0MKYun6GS77WvTQs7Qo5yBwY5/Wzd47i5Ll0P+/L3UnJZ+3ZMudu2s
oYwbDLPPS1IV/0925Erxm4YfLPcklxKqiE0QpljGZOmPQyV+rSmXv36G1J99uP1T
7GU0/N58E/gZFRuCd4UVF1/lYLA9gjMkpXqiXjq5HlIIuOU6GStS50sKNY2m3brx
7yOBOHT2w0s+WTfD423mPMjhX6mC0YX1PKdXBlBrykDUQR8K/WJrq2QD4ZZjGKbK
XPBeh4yTBjFMVx+QbrgtuHjnoFRwS43xYHDmW/v7GmsszNJHdXiaK1nOg9SaEo3F
7+tgLo3S/fJO/P3YTsp455QOdxkIT7bLN95BEv2HOwc4fWZJW8BezS0M5nJHQvYs
/A7zlkLlgoGFQc775FmZMSjJWtLa+J1D8T9P29V4n3ZDG5l+TZheCLr4nyvawTUY
45YRkpi1OtFcucBG5tw370MhrUlH/8ZvztPUNjwKzB+n6q8dz6hlVHu6lAUT8QLm
1khbF3ULGW8VQ/AwislZPRL5FkD8g6h0dy0/cTG9ZUqIEoSOa8st84qhSSdLHVO4
fTY6ODitesmRZdFwZYHCli8UFadMZeaqyvWqrrzbfFIJIEPNw7yXlrL/npiENwdC
OGpvMcD7tc0QNZHA5KMrEI/2RQSqFYpMUF2fOsxS9FNVF7jmMU2iFdA2LllKLlKy
fBnSmwT1aC89146T+n4UXOdl+9IYATuD7Kxf4X99BkB6giL/AISRdCfiCcj+W/+I
ZQXYT6doEeoOh0EVIY21FTPIRnfkLq3tL4/WHTwKgTfgpNN3bA70n2Fpc+O63ydO
QkGpyByrObyMjkkA2TBnfYH7gZOM6A8qDnmm1ccQDonYEZ9SEdocyYJHIeyRvVbW
cSjfJZElILjedmLcrSsrUh14zqviY7Y++XX/7u9qVv7f6kRdxxLyi2oJX2ZR9REe
atw4Kw7GROxrvIsQGKHYpKLnLBpEP5oyQ767n3XsjtAcMy6MNr7eivXBDYSEwuoj
6uOY/cJyQZOHe2rIUwe2mxY78dxCOhYx41hvlx0h7AM1ZJRV1kyNwwAyBsB+JIwY
uZutxC/0I1NWuBK+2nl/9808JtRbM3zA9bvccNzf845hpMSFZn2MlByBXkNfcePS
J5ohQ0AEK3ZklgbTN5FT0GijsNJ8qDT1Akd1UBy/cNQIyRFBOugyqZchgydAhb8o
sFLSs3DtU419tQuW8CWcHsHAKqIvFYQvHogJtJQM8oV83NS1xGm0JiN7olObfuJB
JsRyby8czBdZWWh02a/908TSWAuirtaLvQu2CYwrA/p5nTDajiX5UmB1S0fpEkwG
yryGaoACGoLaQDrBvmrMGkakJt4b5T+cJYtW0G+JtCbbfDB90NpcaEa/rSKzo1js
NV8597UXyvTQAH7b8yBWRpPip2YF1M6FpT4JCegrGNPKDTh8xGqe5scKFCn88n8C
aPkyfODvSyCLS1wvb9OjJzYKvUXob8h8+W/p+0dw24Eqy4r2FmGQynCt7OqNpWwv
4UwmyfJ6gPyCiUruVLXu0TrQRR5DV/Pz2rndgR0r4sntVVm+vdes3GYR88zTAa4P
TkHmf86JouHN06vhu1gJCR/yU+QBltSJhD4VRfYGEBxK8KAMTJY77CX3IRXFmG2f
oTWidPbWTTRx8TEK57IFv8HMw+ew2HLTko9dR1XwhwOYxGnUokgojjkvYEY+4CEC
lKGv/k4b3bL3C0HBoB0Da6SIyaW8cZf0pynvcw092oAhkiQDz667TVjLU2yDGrZr
QunV00txqRaoJa/G9eQNJNgtNUODToQt4U/St8RmicOgAailbCkgCTaexUZ3HMD6
eh3uie73R0SyoJvMfmSEQqC5sadW/BzjnhnkFjgXiFdvnHgh/7BiEF30MQqKqX/K
IEe5ckGPZqflfLLx7guVOK+rY+/2PMasrgZuo3ddwP6NwuFUeVgg0eKqinKwCael
TKJTRA5sx+xRswxXiPAmjmgDiAZdz9lhRZboyZdDSOLJyUYwcp2CfgWU9ugUAUyj
T8zBcY+/jCny2dBeGT7i5R8DsHZEGfWA6X9C+oBfh6o5S8XWZ1dSbkgt7RkU2Q1w
QBncAY5eUoQyD6lSxS3trAYaDtKU51EESV9HsG72xO1OQ+rktdx71VyK4g38iBg/
H1vTinmm8YtfMwSo5vy6wOO6R+8dM1bJMbtuT+j+Zbh6YgJmbSh65ChO3EKDeXGx
vIlZRSU5NWI9GPP5vKyExEK+EYZY/5da1xWDyW2sBSfDB+79GdrQDyHCM4UB3qrt
9COetB2QwKAM8ldEaZ0eqVDqzUwaiC3qal71FEiMmErPt4j6H6URqaWTHYkNcF41
Pa3FBvwMWgna/YUeUUjc/3Yyxv3jTWnVFM+8ly/fxwV9gBPHxHS8vFLBH1/YV52Z
hBsMs9yXt6m7ktjnfR7LwWorXEQuIpy/e9un+K0Bo1+LBoRRiPJ5S59jGYsh0jga
h3uGUEOa1EtVupwM28ImVVkdAl6bCsJQYZpBR80U8r6JTLP7t5J6jL/kR28aweI7
h3bZEclVLrdr3OchmXWBZSlQY81clm0k1wzomHkpb1+SO4UI+YdZhA0s8hWVwOM4
qbFCao8/pn4o9lsWhhEyMmZzy7cwLzmgUUXqL5dmYUzHbsP+XqiHDaOJWiMe6jZK
4Bhp0L9qmVcVsrbIzDu1Ajw6BZ3zEgHhudqjDwvn0GlUOOGFLQvSQQUSxExbSVuu
+Q9ZKLSZ3eh63PfBgMflChfejgjcdrXDNnhjiYm1xOsdD/hCyNdB1y7K8KS8Iq4C
5IWHkrR3MHSs7/YX7zj10Y+wG2ATELjrpdMPifPJaun5KsZJG6Ich1+6h10d0pkE
f0e4ZXKUllGeRpe6tDgymHsb0XbCHiUCFpP+Zn7c+iYiirU+dd/eqxC0QyLsvqv7
1jRYWWV6fq445AzVr6BDyuNIzoB77Bzy1MNscuexiIV4SG3A/WUYEKlyQsoZ43nl
V8tn2lI/jGw90/kTS/uNxCSVu6E94mqK3On6muoLN1xmLXcPwXPYrdYa+dZD3dr3
YCelw2OuP0Syl/vALAhyaUOPA2sUDOO2fNkLkgc55ZWEyzACxJ1BZN+liZvbQ6OE
ylCWoSqlIxqvcvis0IIVqu5UtRdTCEb7pqcswgVKfWQSKglCPnP39sl4VCXOWN9H
6ZYHgmYaYwU3HCxSPi30NZjMSPpGm5BjKh1kXX2TlNn5vFoQd/MvY6ZTAMNcvwDm
k10djcvcrJF2baeJ4kifQGe1AsGq5GQ6iR/51JRdEzpJVu4f1eW53qtI+m17Vqix
8PWcB4QKl8tZ1fEKQs4dJUPHmnvguZ7+hhHEw59kfEzmyY7lhV2CvoGIlOa2M5MI
YRo6QQ4IwkNBYbIvT/TIYiROKdYV/xoxMNJ7nwxPkrFpe03INio8AwV9pqS1A42L
kMQItDk3v6JL0PyLoLK1TddhNCAlI+V+ekYvx3SPp834+TJvPWunF+zgWIZOskur
k6hIUMHRfhu4qfsjAl5GShfBM9cZRuA5wEF+uS6RhQl5kRZqUAjiQvUUuZJEAaYy
lstzM3ZqxE/ws64fjxpYhcQOx5yJKVa09gS87My+1GnPkfgSjU89D/ltdf47wdAe
HRxru4bY9LIywzI2rRR0vcDOOOmYl/jcWIMT6dJvTnbS6fBd4WFb2FIfbQrWD9zo
Py9H1cWtQrKSByzszhYxnAETWG9EIJwci8RIfpUh9ixcWCj0iwjldnqzv3BfvPBV
aKzxP2DBmXVo2/HUa86DuBAh1E9xLYMA+fJBUl7iOpOpycXhv0imO83DiD1fc+yt
5KnRBX7so6hb3ZcnINF8aGvfjaabKPUGJcfj3X16ly4H4OdVZNxb3Z8GvTE9Rp3K
f2+S25+XY7zw1zSz6Q4nfOScgdP02whTp0WgAe7rF8MKGlJ4I0b5p8OQUcxBsyVL
PJ3zugNLVXt/4918JmW7v5sAZcm38PNPnD2m9l3YhRwduEKVe8ut99GMPNAM0/4J
mDOVX72DF90BOINwMFRiTmWHkDtVnN++d/S1M0aGiShwXcu9dsCxrjVBOjuc+YNE
vaE0oup+iH/r3B5dfwev8EwYr6EEdC04ORnn72zNleAVnpTVWryCOnUxBNv8m34J
G6S+7M1wvMeLdyDJMki1QahCfqIquh6ZafXvd+6Bv1VgQEtUqLaz5gPD+A4FqvoE
TGHP7gFyVBeDbDY/fjM1YGSZrvBFwMuVOsWuOUsVBRIhP83pSuKoagJkAUo1+KEI
ADt/iDpv19rTDQZ0v3SeNsm8pHDmsUNyRtARI4744B6UAKycdYms+m3LAsukotPF
OXtcAOqmbjQWEvSAR392+ULV13MyXKnLPNBo9hxtTlVZAc8WojgLkAZLihP+2jh3
PrmLgAxG41KMgdBuA2VFC+Opc/L6G7RZXL+BzdTgQKg1nhJekcYlmYE898Wqq+eM
YdiR+k84D7MvzGkSZr/RXVZqtFAYjL4jqI4BBp0nk7gEVjgydgE1zJ17oTPM2BHK
XRqIPZpGJI8+E2XOxNrIx5R7Nn2+Kw1/fG6/jy/T7TWee3zOKuqfQOt8C+OYYL59
/QK0XV7y/SISAcbmErRTVUzCUQ5uuywL8I/z5Qrfvi5GnzaOMDoYZKYy69gRCvns
jCQsYjGpwg4ZmaxI/SqCIPUPsBuDWvf0BsVwZMZH+zS9sJTnUhkcR3uMtAAr+tym
9wZen9aRMslZjSMUEW8cYyVtLM3ngIKiWLLCpNdVGCkOo4Al77XnFY2GaOqwnV8M
CubFu6brpn1K9SU2lX7foddVTBnPXpNmF4QdLfzc0CxHDI8EtxIlmy4GzvqXniyp
CmPsUW3yMwJJJ4KsadQIaYzgMZfK8iOnwvxx3rXM6lo2Zc6pFltYh9U0QVXhJU/F
Kd8PtQ+HdT9dnmEShBN6tSFgiot+E7+PFWFGY6QJKZORuNsbUxwEmwV5XdWXGHIj
G+aiWt6hdRoVHAQfL2/YWruLj0LZnnJ9pBPpTDT/r4LZGWJAZqDlJ299sVAW2JSg
7Zia5/ohkTupMSSSEGGZ6Mt/V2981o1+6xICUyDBiCgLGzTw/Z0/aYSfYyEKaVJO
fIeDYRrTwudvXegH2hBJ18quY+uhRJuussNfSQlM32evLiZSJZQM5aw4WzWkIKB0
NXp1oR+ONJJ1Dy0e2BhGwyVGUptJSA9S/dychxcFGyDBzO+LSZ7r9HhSmup8j93l
3EuPA5X/kVDcSfIW1d9yWTITW15xcNbCCLCH+Ed5j3coh4GFgXTE5/FzGqRCsNYk
5GEQLBZ2mPQCtE7FSkzXY/Rj6sBj+/laIk8InKkJ3iQwQ5a8LvBz+Jx22OZqXOH6
BFhvJcX5GsbhuisJasubyJzPSTaisKwGnkXOrI6q7tOhTFAfTRlpH0LsP29eLJX5
H6GG/5KKXvX2xMaxiWhnnr/vB9TRpv7tqh3EB/69ZDuNgIFYeWvNnrNhMdcDAqbZ
0SRYv1fAqUcXfGQK5HskCrturviQTGgjH75hhSrM5A8Fz5vLWwrV3zpqtxzS7O8U
0SPqoekNDUox3BaoI2cVkwr0TcYc22P0Rn+liOpOrwfkaHz+AI211yRM7kmfZkQn
lV69KtRByj8yr0vm4d8V5L3BRccTHvW9dX6e6oBNfJw1cvvzQrfuoPTnil96Alna
1M5zza3orYTtJqhKK7oFtPJbKkPlupsUQ9htqljnU2o6YWIGvG2KvKAFOFKReGI+
voPnXrPMLh/6mQtF7A0WFfmk0GM8WZXQ9SrEtdYIH94Et/hM9dtX9XjyZtdCC9md
a+vpIQ02Li41YxElWB1uVK7ZZ82pPLKci67Dz7XD8Xl21JzkD1EZALKplXX3Ojbm
f2H5ciVyGvbrl1OZt3uFC4OBXHynpQyko6Qvn3U069/Po6u5wL3gbo7MnKjW9gcN
VgMonl2GlcGMNzCO2IXToHNF5h0EUuf80P2QkPAgGKwUfdpbG+5XHOURoEnPNtJo
FhF3q0APmBNM/ctfrOlZAwtLAgm0PzmlAT4AyUToPhEijkQkxmjq1KoekHwknPtH
CpKQmuJWVBRBDKpx/IsHX/8mdsVUSQ3oHogBTrqcDW+f59BYjnv0PaekTURpQmNe
Ylk9NsiME0BWrDt0M4QVg7AVdF6tMNFbIQ8eUXLtDtmXGn+pcuV/BALaDU1Ad8nt
31RZ1BHTODpv2CHF9lz8uwrxLgpcVMfh8jWNmI3SNTmUJHjdbhPTQI7QJv6UjSA9
mGx3cFADAH8pCrx+s7fFf4C7kerRQz2+RcQG5Qjri2ic7NetiojZYMzFRRlOA7b7
I5qvflg6HcwqeRrVBLHJ9MbqMz98iRb6iq7LP/oSei4o8OEJtVhwNaRTuc6qPTf0
6Y3DR0S4n0Mk8QtLHyzU6emH15gFuc8CDlNWVNdfPcDft2QNvyD+jLfHyfomezCh
Ow1EoiihqOFEWXfM8QeoHgLD6UPLdRC05QEyCd/A9BlFRi3Z+rNtSXhuxZW72pR+
e965/ChY5S7co1bdoTn2D4Y5UAsEmvOLRiU9FD17TzYLE0ckkbr6SRzrmo2+OaE/
EJmOTXX11PZojbxAypC9OXsnAOxnvZ8Zt6O7HyOTA1XQtAEp7IjupVViVqWS0IY5
D6y68g5O/E42P5sai88IMFyX9QAzBm/uRQC+8y1zPA5AIA2EucIKA5THX0mFe9Va
pt2q6sVEueb0ZyouD9wXTrIYicfujtBduFlAmcn69apPgAtJ2meetqEPrwrjqPLG
Jp+ryeeYqcocsXR/sonk6C8FksMj2d/I+9sHk9J3tccAxVHKFzKuHg6PiA7evr7r
b+W988KqpWIP3T7XraaUtGFUlP4XSWxb4pfceDzGBK1Fu+IEVXpY6mlVPD3LQgo4
LAyraa1hkD7cT2numuj6KwKOgm9qCfY1qWmT7+Y1k2FWOZjKxDx1tJoHNgdowK7v
mWq6nuGF8ol5yMhLM1d0MWNwAry7guTriRuKP2AnI3vOXtOHFn1w0n4iKKOOaAe/
5VY85/iY1BweujmtpyprwbSczN+IVRRN489Rws64Q+gty4FVn2AZoxp6F1W6+vcd
1tJxKC9rfSHxYek9R3CmqrTlDchqqD3/Jl6PwmQB8hmd8wvmBJAdm7fgBOMbt2by
kv3F76nhB53jyS6VRzzYd2ZC8soEDXjOgx6UklIaN+UsCNvJSBk3meW7N6cTJ+Oy
RV08v11bFXpd/qVRtEX43rRmnuFli27xkIiTLkPVdBwiF29ch77f3mHukFhT1+s9
Ndd01JEyHA/YvUAkIPfCmmYkrnMHSsncR+H4FlMMYhRgVEZWYMyYVVZN2cjcah3+
XeH/o12D5sPsA93sd1l7RBUd+IpAP7YSjWQaZUzNjY59bQeTb1Feh6ILkmvShxtD
7SMDYBAqvVtDTkP/2yttx/Vix/U8ki8gCgTIfCYmZO+o9ARDt0HJUcqRiaKNOFXn
ZJp1/rB6PWpAw1JDvtvW/afoJokviR0nHFIuJUJ25haxZNlcauDNK5fIxBAlwFQd
u/Aorwm5ivGybg+ZS9Ru5IVEzFMnJSOzfz90yYvYyUdIihQUOV1E3dOL7P97V5nG
AhjpZjs6Qxkewt334QraRIwPdMUvRRbL6Zkf/Vv3M78NGll3piBKC4HwUguIA7BN
AFEZm07WqkmKv0L9Xgu063HwRzTVbJyORNZmWfCGdUboAauaVs7u6C4bl0u3NiOG
j6HXmjaNEN9o6dmTnvVoFBf+FClkWqmdqWDkHhHhJfuWjwaafEuTqt1He5II7ERc
/QgGAHpE0pzWHuVQorOyr1owbvH9qd6zfRQl6vg1oPZjvTNk9dE1yPtIbdR2AWeF
iYR33SjYbOKi3T/CZJA/fNDbfizFd0ReojI/KjH1NNDq671q+UBtcFysAASDA9Z0
lJXwUHuAZuQp7Sm2NPX+m354QMm+GMrEUzIOOi/qyK1xCl1YpvYYlT84rZ1bMYAv
JfPQ/0yEcxomh46/BBJ7/y+115nHsx/mT1J7c536vihvJvqjz7pPMOIhH+gMg/cn
PayWO5RS2pbI6ApoO7z0mpucnCaEcXpAiDTglb9Yx1VazJ2Zb/KzV3kcQDhF1nTt
uTdeYzq++PBr6o5nqM1Xdz5yJvK3ZYiSy0nrcxVOK7X82ZARYOLCdXJTbfvZ8b68
lihPAGW4JrveLyxKwCuzP1Vf2h3MiCIbYGKXqXnOX79fM9ESXxfw6Eps2Rk0Ltrj
n344FxrLP056wETXAJRIpYKZmWOkZtp8UItbAV7e7+zIOuG2870Gn/MIOhWrG8Ao
YDifz64dsHXeMlAZuST6xp1xsL6m2hfHTmN05TZL4E8w89CBc2Ibs3SVPnRYaJW6
shVjOH6aAmqjp87n1Rc7jJKkgDc3h4rKNY5d0q+lzTbdBNMC54HdfH7rjC/ON2Ds
I7K9J1vH4USAgfUBnDjU3CdAivXrlLJ6FwnRa5cTqEEmWu9SQHdKPBlafx2L1oda
xuO0uiqC/4zFmiktMf/JgV2ozKKhcH9mR5DKxspE+bxMsqkLCNBf+6wIBG6sBEnw
KgYdl/v17wotbEGqJBvud6JRdV9yDSwdwLBm2juD4RQkI+DnkQcoHAaqQ8zzD4SR
XKBcRp/+/gXlKRro+N+2UrQqCBrEaydFxGMb3Z6KEgQTRrdPOOVLJc2u8l0nLpQl
sTjTlqI7obn5DTDu9j4c29Eg0MGB+A/v0MFv4qmPwGE+SF1Dmc0pcegkjKOH54I9
lCWgwipOtMXtc6HhUvtTSXQ0JQtQzlbawbbWvrwSsPtiUKh7M/Yy4EjGnRp1/r7x
LO/3EhNJyxQ1DWXnL8VjQlp0SxwB7ZUhRGMAWy8vGdbom2EORAFvOfb+QHwe+x6k
y/yJqyzofstq/S96sNxhdNsN570WMFoeHfZSRJrkHSp5RWrQD0cfngTjd3v2+4MX
78vnND1WdZ/DUk6TKlRoDGELO5X5qfZaCl1rWNjVlb3H3NYfqRHF05A5rJSuxFSz
YlNQIG1aPss9y//1n0AffW+2IWW20QnYr1Z+imzwouVrvOmx2sahjeoDxtQRY+wX
GNVpu0lTHO15shwOsFlHUXa5eeVNuOlQYb3PiYF9qxMjSKmoOUfIsW64/Op+Og4Y
5JT1e7tvbV3q44v9Ijh9MDdrpUjhIPkpKVhlGoG41oCsaf0m4xroK1urf1QkmcMi
GDSlHF6G5QKsQlHzGABxRDroecUIEJ7X0/ll5CRfMZrWNMov1hS7hYil9Tpa1CRU
mfVmCghZ/HJmWeB5xEM3fwyV7+qPjsQUr1WH0Zih31IQRPTMT5p2wDFqX8cclFVs
ubhBum6yJcYU2ERLj5dAlXWXF/nkBSEhstyR37ETEVItLW0FIW869mHU97EZq7j+
svPkb0KCzH4xF6NmzFCleqDP0f9TI6E1jp7GczT0nLh9pp+uzMmEUKQv6PrYs9+K
g3yi1yL14S9rcp9z9zwKBXe3i09JMYGNbizGwNXXWva2Eo6ulyYy2B8DI7c1lLG4
wx3JYmtpI0V3ltDH5L4rDHLSOxTYuvC4V6RD5HsXduy4DNN6LB22xAlHqknYLWhd
hziZeA26Xxg/e8zuUZ10FDsAIC1zcFPJEVN2MT2Mh/xF/trc/h8twPTz+s6Lw6BO
Q7PCo0doRgJI/Fpw3eFLeIwTHGmO8ZzZd3vLCIsOUnWrUrGRYIw4qGzeNjKQZFM3
OkhY0c9h/nYIX1euE9ZQwZqPeJUmm3Bk6j1ZL5/hvKrrBXCwNVi4iHeP0OVPnyZW
vU9WHhzQZ0RF1oimKVqj/y4vfnM0u1msrEHuWX8Z8n9tSqptaPvuvC9dm7RVsQQg
DRvT7Re8xeUofhPm9A2U9dOpyhGvGDwcmlGumIu2jLi/T+rtlHTE0Y9CL8heBz0+
7oYAfZR2/xLn3LIKA6I+aNW3oBf0/XXicnd429rtaB4kMkClVTB6/D1pIp4EUzRG
6pAT1HVhlA0HmrWYanijXdaGZ/NwMoexbl2P3t2LQRqM4ZfANLANtHJc77aa5j6L
JeD82JSpxLhZPIHsCS5HSPd22f//4WKEUPS/LsHqYapFlzKzmihQhtrazhUH3rtB
CK+cq3LWWUCMPXr8H5/Knf0HTbh+ypura30iOJW5Lijjx+jnRqHhtCKHR/ItJTBL
u/iZRkL7PdEHhZkPWbVvBZahAEyrYgWfVSjDbKokIlV5Its153g/IRmXX2g3GCwP
cJ2wXykpQBrY6zlxVGGutFJty/lLW0IfK2No5TpL8CjzVTqB4jNt4B9NG1L0w0hN
DxrysL4pLo3vorPXCSxUEb7/RkvWy3T4gQxVD9e1+a5EvdhM1gFkRhk28JFVWx42
joIzUPXiVPBPv521esmHzQWYe/GFi4V4AXMaKZyMvR61VFsomZMiNwi1AeoA73mX
d1xlIRgrLpGFINXGiZsrrJ7uE2GNR8kfcACF6UfoAgFzoCIpqqoCC5MGqqG/C9QB
BVvdhdMnzZB57Mxx5vY21m1QLSoOkYD2jaACfcLXhyBu3yvaiVkwxNIrZJu6OMLu
V9VeFJyTv8RG5wyEXQAK0ovOeX+LNEgUNPFAD3c9sWAf2qTWOWTs8uZTcOiu5BNc
YlY41tOd84AIcHfYjohq2BqEV/RS3M4wzH5Q+3efaEFTreMyhamE7gW0S9BCq4Ly
OYqZ52WXYWXTDx7vDesk27eeyZiE79czG/VC9GXBzC2LEqhqWPvYOYaEvgXDlkBV
xPWw4aTWOznpu0A01+oVVGF+v+rI8TTTG/wMfksvNpJLMIkSN+gkrSAnit1oiLXa
Ez/tLCun8+I9ypmZOSOAR289QMf7O9+ITddfJ4EhYtZgvGzG+o/Gm22ifkRmjd87
W/onqbu0qQuqjs3nJm6xXrsFc3yeH4STmGMXpkRnuacVUqrGabNTlyHIOGG+75lN
WoQZRmOB6PhoN/MN5OZdhuNUqTSt+74+mcaytRDFpv9nDJz61wYqn466lEfF51QZ
U4cPYyPln+cNoh+C707o3r9/zGDMW7pCb9PbzEuu0ApT41M+jM9JJd3qPVMYX6rF
K8c4WF5TXxCrZS6KocZOE8wR0ZERBApWmvtePEEBtxSEW/J4XPc+f5oZgnrlEUyS
n3dD4vQLGnwtJzN9LSj0kZlUGCR51yISNJvwbC3yH2gKjsK1BVwXNVOXjNmoifZ4
rsBalCJqhXF4wlcZOPO+tZERdNk0J1RcfFxBSDGef1QZShi/IIGx33Krrm6a0ZYT
Zhk1xZZoMTtla/rbjIzQogayWNi+Q6rVVM6UZxWvmwi2AMbr8VAclvWC46BveP2N
lEU6ek1GhFi0aVldCs83rrqJN8MUDhaDLwlMeJyKok87abRByeKi6IZvD7U1euoP
PyvRrgqfmzM4bwCEPevWIO9JwG4WHsVNPFaMsYgpvPR5kRS+dUzJZlm6QVabxXVY
eVjZThbBfpnz7afbPP/FiJKee9nRF3o8R0/XTJhMh0Gm/OjtsV7zfN+b02gFaS5a
SJ7k1Bzc3JBa7rmtFXybgPl1ZW8iEoNW03/Q84Am/YLcm1//70KtnnSTTzifzi/E
1eHpyCAvyyCX7PqM8QLMIP39CUjFmKQDBjsCcaoTl9swfFENgXUUmEY3Sbr22GQn
OfH0s726BaEUTvqhW6cU68HThUA2J/bRdtLRwoxHEry8h7Fj/HZGdUQts5yKB8ec
pqmjMK4j2DwcodKWvWyBx4i/4qwPy3ukxv/7xak8Bkxsgs8XfoNvYaHec70Q3tSM
/MKdTa2r+1JkQxWOsKw+16PEL5h61+fj0LOCGXWmgTpbs1drZVFhww4YYZgUsuTM
y+d2sLH7VdeOKmd3oKUgOrqr3lrtkKIWzYLXpRwV0fpdVbM3Y1j7QzADuaDHpUWU
IQ1B8zWqLr3u40eMHeQIT8QJI+v7HoEoAPxl086oSu7ab2UWF9S4j9SnpUgh9OYj
LNrIM6ASRFL4TcQK4pAFGJts/QfLK/3GRpkiH+TNEJBPforiV8bq80JoZJBXZFGr
+mOizT1dPiT+1rcGFmqS9gt/MJyTYW3V6HH0l6z2dz2kuZJIZ0IvY9LuXq3E2D0I
VlVQI4SlYAewaLfrRxkZrtfFDJuDnGEbOG5yR6tIewG/Jyq3GBkjShRDHYRZmwa9
13h+/x47BPJIF5RC8qdefsLb8V7S7inqi5mzcsywQCFxrFd5F0oFH0LYPUhdLTRi
rQSS3g3V+cL+eZO16EdcCnDNFcPkPYFSme/ZdGGgE0Vnm1qW6NMbtAMHNP4feWJM
uxMgV6hdCUcIog+d/VHcn9Qfw8GKLuK/mV3C8pl3DOPZScTCw7B4/YO1l0D2Pw81
mW/UiwnseBmf5E/CubF/yr6jibPYQHAeXgD0cPYquQFKeRpWENNq27b2626DLRlo
RTA1w2wJNFMwLb/3Qf6IV1eYi1TK0TbYqdrwlbRZ0KJlCA/4oCpcixoL2kbKdkF0
n5HsijmSP1cFb04R5RLv/xcBZisbWcDLn54F1ZKIlD2arUJG2awzN3u14tiFLuSx
7YSoP+1IPoLA2yCSAlVH+xQt50ULIMFXLckAxuKwri1zinYFq79qGO8k3JDJZGJB
AqdqIOPjWKVzdGMRn/mCjy8O8yxLCg2cVIPQLh8IyiyRqs2ng4q9XqrD+ABZUKlF
yiP46Skhy/fpco7h2cQCoiCODOkaZu/9mvqxDSkY+gfSrCsFbOL7YoT5V9rruWWN
jEzhkPMgQAGTUm60iXFeWx+7BOvR3YqZiHYR4EnAtloZDVD1ZcBE3ymFYQ2zhc6M
YQKc8HsM5brWlY7fWLldqxppNXeDjhnC+6O3KYVQM8fABiUygEOPax/TnknVzbYO
i4PheUMo+Ole6Oa8BFNTn3OT1W2BGSYK0ceK/+dqBIHQF4sODhnBzxsczvz8yh3k
fsQv85XKoN/pvst3s8f2zw8+Xz3QSh610vPFYI5c1XBN+xpbCooBVjcKj2KZsQqG
FbR4QnDhUWCQKuCz4tZICSrP2iF3czZamrAgm7qOcM86GFszcK4YgGgIy872/1Rg
0EEOVdYVw/JhmBztSh5Gu06ueilydvrH4I9POcy4EXPxygUI267uAXsUhw7XgAza
NvPOKTvcTDdwzj4mFrQsqAufEQedlAxMu0PII5uuXGmYBYIPaqncObz2sCgpPccK
fEIAc5t2qImAgOQpWFAPHzFgKHXhZ7fC+jb3ttNfhNUvNCJpkaxQAzWdKJaarkuZ
V2xO3Ay2c+3CE+db/auE93LgFAHZIcWPfXJbQ+bBz9bsRIr38PewWoW3RWo8CxI/
zUqWVRWFMZISpB04I+uUOOIKOE55b+ZmaOWdyaaxUKb4yVEkTdjNna+T5zHbRFx4
1PKTn3G/J/GuPPeYqbmYXNARq7IKU/zn6MHv0E8JJMreocAxygEVLlGvQTISTFD2
1lrAXp1akxSsUHEP+NqnFyl0qt6oOiCd1eHFO2stRro2x3OvRt5EOAbcAe32+VZV
Oq0IlqDQt0kiu6tMH1H2GvMVpOKzLoiRcOG6xPwhEiJVOZHdnj3Me4RW5GT3PZVU
XmMs45+dnhLX7RQgzrESoW2gHehybv2Nz3cBuQ+m5okJE2s2+OtPIoz8/qKe68D+
b6Yo2RXR0Dmj2IJQ5z0uoGIrtxCwJU7XxTTkaxhYW6bjVpk0OTw+e0yjDfQtNDS1
KiJotTgGRWFdnaFELMGHdOjA//82vTBmMOhR1jQtGDd6uj5erb9N+IMqZgya9D0A
WlIo558Z1Vd9MVmjTHRqXZxSFHY3j7igTE9PzYiVqdifL9OhknblXwaIUOiMnvhH
n+Fta8tVOjPijGrHs24PKs1O3u8XG9Cw1mSRF9CSXs0bGDkjWlf1LqBQrYofmLka
DLas7uueFqnPcM+N81CFElLpFOkqFTCVMaGq9t0OjkMXTbdA6wSEbdGtwvpxn3Zs
tl+8lMFv9ioO/QegGeAxn0GbyeYuuo7BEyP2zW3Hnys3uzdzYtw4+kR5pDFQfPg0
7oLX1DbxRzmSMImqmnX09y0SiUyHkseuHzq+R3fWjGSK7Dgf3p8nB2aGnaUj2a3V
M0TaTFGILRUUjbQoIqVjT74wIZjr+hfIJMCXmBA936KGpwLR+wLIe894Jq7MHoXh
2ssWmk0wlY/HRuIgKSuLDsic01EbzbzxQ04Ef4BnocF1RGXzS+vXf+w6wYvgV8Q5
mfHSW1dgIM9seWqa/9vbBfg5PukMlu1uJlcIqlvxTfVqA1qx6hdK2537RycDR7dR
tSDa9Npv4ca1MVtUlbJY6e1GhHnII2a/OPefVttcrGThEEIiorXm6Ewlr8cHqG1w
An3GiR2NLPW641OUeo7NsvSiTb4/4VajGXcgoKBsf9kI8fU+IG2m+6atC+Gvh8eO
1RJ52E3j4Ur7fj0L7L26o02NGDDKW6hqYP9LgRX0BfXBDwYZKYshGS+u5E0yPZzw
WgIWDnty2W+xyjWuHcyATvFBMf13YEm5J8HlSfotkzPo+EiRCLMaASbeAx3mqiey
H65CUMkOcBuu5CTYtre7wCamIbnmEQJgifen7NohGrXAfVMu75jYfZXPDFicRJTI
RHYhwIdzujxUtmT5JRHaDSg0hrEC+0Nxjt15nuozc7x6x7UwBW8Yt5jovVyzd/35
BXc9XG7HtKRu4u3UWSMUTJ4khPwrRhlq0KNI0bZH+n8XOSv1PVfXCGYytzES+ucN
3sZsBFmn77VUEwhk2gzrMs6I8ZDpzWmIYS9RABkYMAdcQMeKXl61jYBbKiCl3iKo
1WCfPdNze7k88xLzuHYeRa0uO7hEYx05s473vMGKd56DG1jH716uBBCg1pdxb6jQ
DCnk+rYifjFX6UkZ2jCVQqBtRCKeJPlGA6fk4n4yIx0a29YjT11Z1sC2ibfVakTu
9OX8lH62vml3bmkWkXxTfqxUXJA8DnOrq3tvrM2LEiT42BwX6x6jSYM5E9jpRcHl
a+URJfG7gknze6y+YXFDmFxMxWUSxvQdxj1KihhL9CegQLJEQ73zF4scsXSfSc7U
2nn1TXXspAav9vlJnTCzEUwy2K5O7RyYLoELHucfx8U6+XPagRNoEsAnQwPPVXEm
btzB940+MMGALpkiR7XwPYKXEHTmPJJT0wmuEVZIJIw/FsM0xcT3FbMwBIIQzdST
jAzRMeBug9/8lALwBOih7n2N7OsqqsuayTFJAp7Qrxs/UrYEXdnnWl1MnLcw1zM2
/xMsgc3w+4wLyRIdU0/KqczDWQs7ep0bDrbD8wzEu4KEp8ZX143iZKOHkeBk4EES
Wtia6tFSKqnkwVmSZm/HKMfyALyeBVn7EXsQHphedLlsDbcrk5a/Hve2Z+Xfg7kb
REBRTih93yb5xAGuvcs5ao7kK9F02v0660XnqtWpaSSNkS5xY3CaZL1wQx5/Bu3a
clMNCbk+xyaEqtyXxB6SlOTarX5ansxvBfV7ykfwVcw4XbVQdw+PQEOPw4sKT9M0
jovzkUkTrcdRtLKlVF9yr3c/XRC+tDuUjESr70uMI9g6XYcfR5D5RULkdnNNzePs
dBFeLa4tDC8nAqNoRdtxpkQWn1lvyffXSYqj+HlLZou3RiY6hdpw1k/9VF/QFreg
+6MR2sNNz2iZbswBZvKkx/oB+Wh9UeuUGcaJesI6BPRT97+oJpa/LmNhn7pSmSwr
1ZKZpvlQA1ckeY4XBLwpf0Cj5MQwdUGkQtf2rKVMkcrGzwisFreuLQRHKaLJ2p5T
/8Yiz8ceIgVPYIJTJZc5dHI1a6JwIdFui0apT1ihURt7rcRzHiqFFOG2WAOm+JSK
38jsDDeiPxH318aQHe0zMcbvSUPcQh4mmbCcvtw0vEaTrxp3cnH35sLmo716QZAJ
C722KMjmheEIzszSnQVVLTUf4WR7iOhHfXdTADAt3Ss1fSgnI0us2b13BnB4nlGs
Za2syxWkME4HRu/6JVlIWWb6eMdQj4pknd9OQzYyURKNaSuks6sLGODDll5hLkhq
+/fvsdY3I9TNdU5Som2ykpmFQX5j3WeHoWtKpC73LSc3L9e/Qff3xqTHgf3eIe/A
3hGxC/2WHZkZxHY7mnUAG6q5v/XkZMsdi3ozU0KQqqloWzc0mWIOM9OjCW2ndbYs
mrpcQASy8yZy4o17riYFdqDGxxghY5J736uXatK7C9sGOGBW8oxbFoVURZDGY7tG
h6XMXOuOGTWIcXLmWYqNo9+Irp/mz3KAJKEAyOlH1d3Kfs9LyDX9OKm5BHp0RRLi
vmCtlqGV5Ti8k37lB+p12zUqUXDPG2Q2YRK4ZfOxNriSzyeAEPuF03g3uiWdl/cC
M6z9CbG+T1vpxUktUxq9exs0mUnfN0oq/RBASJCogM5sSvTHBOysqwizSGwcTQZm
dy++hCzhHq49y5b1/QuJmRcAQtY+twBfNMtDr+LDy7oE51GQTex/MuHcb/3EUq2P
RRnXEnm8AwYuJDImKvi9hGgs0VCkpo1MnROrF3d+nQKHbOZ4a4YoLHjjV7nNmg8k
Wqtcqk3JvFwkLuTMaPWifGnmYWFPnA8uetKWRslMLM4/4tju/84top8aozsVSQBu
lgoeZ9C5UpJ/TNjPzVIvhNqL+0uNFpQ5o131lbd+Gi6B7DR5vVQIvzrwL63nFvuC
dxmSUgL8to7a7Uxa41y9S+HSvhxYvFAjp45l/nRJjTCb99feqsLIi8289a+ai7zK
fWEvfuTF01Eo9EwgLRLB6DEXgrGD/ZCVvqcqO/03qZQi7KxEohdunAIbD3dWW06y
CknotDlz2xDYTr9WLBizj1BE7v8ZHbBFA7x98qWIlTPvPpMDZhYkDRr7HMIB/Yr/
6laMa/CMFvtrVONJSZ+tTDysYe/Iww4HL/SXY5peSM/FQPJe6mFOnukcdhYbqfa8
fz3cZswg0I2TS1vZasK3F5lC5BsJvmKbvpOKSV5wcFvdnkoWuwNSCC733fRamu2V
MXUy7ujsTjXrm1jQXcTA+JhziWtyWInoNN8FhCfPyCOwcgUIx2WA01jJnKHF1VS/
iuawI4hQYAHnBG9Ndf6f3FPT6q1OJlwHxOwCwbg0/6JZgEDQ1zmG/maFi4ItTC3p
a6aE/L6Jj8jkq8PQ7i4xCg/govVurXk/NKhfz7NUHJAbfR7cZCuOO+DKhmN2o3AA
yOqZuO3LVBPX3A5tIavCGCaTpUfcB3KrtmSKnBlY/4/hXRrbOLHGAFnA6Zw3iHtD
gUL9kDcEGiLXKHxLyN9c3i/Dmk5xFdpoWk/oRbhW5u0XPIr1Q/N15ctgY0KUu0Ya
1fa/PNi+SZhixj/qxroMoy1zodiKQzvsgRvgiOg8cPdaipoLC81Yie8BTfyblZ2y
osTS/Zy6ZjAVMYYq/69tBY/eFw6srwVgUw2tRacQqSMYE60qoNMPYEoXv1lGnv/y
zXdMi38vxEcvXsWPSp/yNJjrqCZsFpwaAe2e6HCnJFSmONJE2v9PaV8SXW1ogbXv
O9Au2Jxi4k3wRebeRJcnN2dtkqG4qxdPDUJ8UUhQ4bkEb5PIM/xh06pTIighTT5U
lmNox4Cg3ydvjflCSCx2pMHue6vurTWlh0CY6zEg2/amCJ1a0fDyCgrtT8GuiGnT
/PKTMk9uHjlJ+2mtJz99QHTxXmxvQyGYR7EQafjvFW/GqiahQpW+aqStuL3pHNxE
RK0fXnGe2ws33EaPnG/YWwzJ2O+UvaJ7H3iGfSmiCw9NRs6vL+6kkQkFhGo/qb1j
nmanMC2Y9qySF8tIkwyr5C5hqRoY80WfYQ4yVEZRpkRfz6LnIj9Ng4vbrgi5VNIl
HohnorolmFQ8QUrnqHLSC/Qt7SV5MpdCYTXDSfe+GE/mioaxqNyiNdLKC9KzhK0V
VlxqwhsFheIMlkNYEw2NxPUDp+a4FExd5X0ZDFlF4YO8L5U8mTno3Z6oa/TkEZWs
IUj8dwzLCdEZ7Ds8Wp0fqbqN3Cl4iLJtiy+lzQKMspbDTUfpObhT2JQh3TG/X+ve
xXj1bNXwd8rr4j1qazgS1gdZe230W5AhJ5Pm6T2soBFS9fhxnP/BZODcmLoqDXhX
7QLyf5oiFN88B/W3tzWzKmsH76YWtJnI5GJrb3M59FJFgSJ9aQK7dTQzBBw2txOs
1muh94GPpvRW6W3cQYDMZG7sWBvFM9B804hnXw6I1wY6PvFA4FhDv5or7nC+ZmX6
rmwOKT0TGO7xfFxJ8O07HndnYZ36qD5WRVCgs1sh010xUVCDRfvagAE2BH6G3z02
26btg8yqmq2gWq9/IOBB0J79qGvaPrdt/Y/jFqwh3DLps/1V7hQYzaWE6m1G4lHe
DorNspDgqMJRZFt4FAaI8OE6sc3UE61wBhgz6i0cuqagyBb2b9tNbtt3hNbNKdYb
8ePP5JtBJIpqFf9zqxlfK3itFPrP2w+de3pAAo9qP4R/MmlkuMY5lHBYjieS51Ps
mUYR3Qcgz9iOyF1/B9NJ56mWCbx9s68lmeo80kolB4qUqgiFmpu50GlhqvRkXT7p
kYNpfGK0fUEL4YpwfA6KB0Y/9henu3z6WWte8te2yFAK4FAbsihXvAl785FtK7r7
qgx/Nn3gKjnhFvKmBm31HCU8I755tBiCdsBh7zaRrQ5sNHLZT3J1OqkgJL4xl++5
Xb9ghmX/0j6vkeiz20rvRuqGw6SzP2Ru1wKFtRMkWt+xmCsG0V/AfhWo62vmRtvK
PtiY7YKKYBNbp2oKp+4BJBATMSQCVF73PXYsE2MvGQ/VEZEuLLEdj9RHZrDKPvdw
uK1DgDNqi1gWv7Y3xqt4cpqpqNUFWIV1dKOPiV0h8xNYzv8gZnqnhIBQfIYMmSds
DWpvuTLVVKqxc6DQvcqna8tBUEwhqMmv++yvkrwKW0fudqb2wGdFA6E5t89CCyja
X0DAZjveGsgu4jsLKRhpjiHGtzJFsPvP9LAcoiVYZRFPjv6Gngub4jEVWzyl2XDd
uFnp5Qe0fduHcQU5MFuLUJOPiMvqiqT7odSCbnJnvgM2U3NO+bLu6dRwrFP87N2N
TDGqXOSGq3bg89cm5j9XNNf6MUF9R0Vk6v72EPol2CmolXevs+rMiZ9Zot8yMnRw
750fgSxdHTfbX6hoJhGBpqdqvxQa+n3P8uyU2zZA2C79Vy8tlqeFV/L4SYvYaUa/
kYKbUHcIf6n4dazqQ773keTotJrdDpZP0zXZccKltQyvWGOM8tgOJr8HBKBYd3jl
ZDt+FEmfAprZ/tvTbBHj6MNhC7HLjz/rXXfFo+Jeb3oKXzFAmdOdoGmfT9OZiRvx
nJG4m+JXrVFKd218oaXvA0wsn5QsBqJIr4tNh7h0Ghzp4ymdlPG/VSUv1m2OaO29
gq1uYSKNXHj08JYqc+N/U3WXCXWDfRSCI+VpPhM9IjeCcLwtuffgXlHemnL92t1j
xW+SLgqNjGN9ujzTstZKzMNQMfNzgAi7nn/I56/JxOx1YasWes37N8d6e+2mHtL6
80g1uZlfSFxFI+5aZN9qXGMLfg3N9Jn4hBIOd7I0nUCHcmKpUd4MC7jHl0a0dsrA
MzAUAoZJtvzIypPfuk75mFX8prb/+AEqqN+TyAT6YL3gT2auW8PXNiDJL7f06CRH
tg//bs6fhlZ11z6TInhCFkM4vk5xUVXtasGKbEFu6hGoSPcnGpwoTbIo2QpjoaeR
XwQVSWWXnvoQgMBHiY5wbaMpNku5uIdM1vznaH6QSOUDHxZQWIKea53BLZkB2e6g
rTF33hF032ua7neIdnhGry6ZUnrUyByqagYSRFTycq96UVbHAW7rcgiYQ9GoNNh9
KnRZsgxdQ4HZ7H/YG39QS0ApmrxRokjaj73nMNhvBQ/HaPOASJz89VlLTid9n43E
/QfrIIK9S99tZpctveNMGWwGLABRjxROiXb5f5hTo44vurBv5CqhW3o4MsBWZ3xW
TJvl1s6dKwPmXX7rLaYpN4E/Fz4KJMw10cxJTqBEqBo0M7qFuZi0qx5nBubY6AFl
KEVZsx0xWogwwr/lc/pTjuVEBJl0fDH/DKrgibjWwIC/g3tcESU7Ej/OqIxzP71b
P13X+Do2IW5JmsKopEDQ1TkzL/b45hbvsQddB1NYhcsMNg0DuwkVh0T+OUCPjNII
1a97lsLT3ogj537Qx8xC2X70Ty4QGA5y0FVyXBF0bet+joCMwO/2WhM9dHu2OrsL
k7j8DiH/RoexgnMPMeIqp+7yvd0k4SJpcrk4dEGn/mNc1r0dDu+JKSdG/kGJM/o5
it4rb5Uq9mXblJG8EgjavDFa+GilwHIhvmUlWB7ZKIE5F5QGH4jLZuAQVKhap1vW
UsIayGez/sLsEm8c/FMT8n9kp/LlsAf1F6vVd1fhWakj9DhDNJgEF5oq6IhcH7WE
cqx8kO6z9gGIo1ipT6cekFU0GVTkKkRL2p98xYbrEFRUr18LhrByOmHzxfyx9SqV
ey/0vlOQrozK/cRZUDbrB9D/8baIjLTBw8ghd/Yno34EzBGMgXEkrSuxgEGgFOWV
DlF106gIkQf+gmx2HGkrXc/hFLr932J5vPXJtE+uEe9ql0vw8eQsvC/8DeM+yT02
8Q6XuWiRbIVT7CIwGQAjbopV+8CWVYRVrf1IvjmgSrBSHRpdVXsZJXKmV6Vt5rQi
+f57iJJRjNKc6AiCz4BxVTxbWgBON3sIKuOCCezyjPMkowwZP/CVsHE/LPtdUAR0
nLRRYreRQiSBfQ/vp0u3RiVIiyX/bosMp8dqZZV0di+qjjU6dIokZW2up8EcgyHV
lxhE6mNpOr7M83W3irpOjAI8HLg1HJePDx5kOYfjjsAmM8sny+7+6kl9TYMUAlw4
48Luv+qpMla/owxrw0T0c378PqSGGxAuXsD4kJPi5KwySEleXQo6V0OiMYDIi7r+
ERZizDFWyGos+ZUHtYz8cS5SYC+/oEIZJIRhZjrUzFWgXO3fZqJu3IBETWTHZVXr
OgjCwyQd7OelMFU8QxIHOYRNCGYxvyla5ktDJudww4m0QvQy00OV2scyGUNaaa4J
NQNWpFhIfBTVDwKcR7QPG/WT7GE+M64xnlHAgWIr/u2tmimfizweQw/X7sZC8+DJ
XgqDXyzxJTTP2Q9q2q8wRM+oJbOfrJpBMx056D1BDCHaheJJAX3J2V4j+nnfC6px
o3b6+NTA+jqFQb+CRQEsSuZUXq/GoK2EUODYa9D1ddKHp+5oz7lLrQYtFY/fHZg5
VP1bt/vdYcYG+YAiLneUOOZxDuYEtmvFxMEWM2dapZGkgUbHO7an6mFbAWR/IVtE
MaqjguwuKW8HhQzKp86CGaG6VYWjt5A9wZXTqLP+7v/e2tiHNtrMezfxqd+dUKBP
Alfm93kV9I0KZWT65q+jsNXN9T5lgZ6S9NGJXT8CaFXxaRPsnbJpbVrs+ZPvYJeX
G6jeF4xQK9AmtHEhzZ/k2nlZu9zLL5d7Xh+nqvyWiZou1US8KPCixm33bEpULweu
9Ns7Qy7+g5wYIoQL731xOovFGMkjg2Cek8rUuEGJ3XRVtmCuTfv+Cg/90IF6ocze
cPoM1wQ6n7/s7IyewiIjPzuHcrOQo8MJuUHQg+PUcfnqCKwZvosWLW2Aio23V+ip
ckdTcMJDGf3yzKvm0afXQ/FTymxqwRwHj+lGi06RHQv8iXhMp7Orz5++RejsCg2e
gQ73AbtEdkGMvFI1gzhdA9aKfVyiKI+H5dFTgsGvEhcnAdMmmMaJ0PYm0fbqb6u5
rRFPJlhuFyAu/gtKkW3xvLO3z+izEVYxVK94JYLCWNR+xBPk9EMLZD2aMMcMWIj5
7FFkS08+6mp/CZ1t27AX4lQGq2/MDg5Zw3pGJC++xCLpASFqdFv3jO6wYnb4+f3b
Cb4bwuWj8YvOjly4wdfdu/hGwQ3JIq8YuzV5CguYWYu5ONsJHl5AKiTnHmpDZd2P
pRZBORs0NpLKNFluVZamBql/nU1hJb45d0qhi7on2GxYUNZ3mDx5a9LjPYZ+UtU+
sClZWoYAyw3QvONVGN8tFoUhG7U/ArzhCPjrQojNIiLUt37ZIDo5bSq9qzidsuBY
BxV3yjwZXHsw6B0u0Sadqk69rRIXRS5m5tOhrwotYWdoS+UMMiHjlfQNmd4kUOXi
t6uOjBXhEYS8pyP6w2WsZw8pdfxUgvy/VSsUg1plgGHbGjmCETCq+JHjweAUtj3g
kT5MGRA5lAB5DRq21JR+6tZeZHsnO6Q8V515yEe5fALGmOZAESEdHSmiYz1WCvGi
9PJJcpvld5OSwLmmFQUcPt3QqycpKbwosNgPIGMz3ovVWTmKJG8wHAdXbOdqRzOM
ZsEQD4tV+Nw4yo7oucjZRRAuoi61hvEL8t+A7zfJhk9+IyAE/QMOHlcUBAj8k28j
eHyXYkLymF+/ddGVsk4ROxyqva/xMDGjhPXVMqNJZCD69jatwrizejW4Yrk8Tcex
1kHfgDPsbLDzGQEc8/hWTNDE4xewB+2CH3Uaq7xZ5rvoMIKcuHyIelucMIKoLYoa
mfu1/Ofe68YpmFTi53+AxOtGNsFaEFHq9dMC4zWh2NlXKWQMO87pf6nUSy5/eVjW
odQS7iUQ5h3jRGUi8vwwq3or6ucmmDhhP6egl0zgeBDnUzrbkEoum4uXWKxx4rlR
HO1hORNLtIhIL4lgEC+maK6LPUXus2BWiCOhokV6xCKN2fnEPaChvQAn1uayBGGz
5SF05oWdAcoxOh1vmPTVdH7HGpb5tBNr8UM5H6P7uTVwRQelmy0adqhFriklwEoK
DtYr9y3KkQUfjn/CjyP0QYLdWdsSriQJxAnWWoidezQmPIjRjKrrdKKaTlW4lRMC
45aeLad8Cn3pksEc5M6D9+WnNdPKI6C4lCKN6pF4yBWM0UXt+fcH39SkPAg/u2US
E3gbIOJw62JZk0VQLO0/lBL6Dc1XyHTK31wsU8LRSRAdXdhIqB16LGRxrlAH6oGO
eFQ/Eyz8GHVsvCzJHdxDySciNoEqBIyWgY0rcDkhvqhyiNaNd3M2VhLA4Lj0zEAl
jXic1fMHLuHAEfGYGFH1X5u6plFSpJ05axJGecHs1Vq/uvMIMvRTdkEa2m6Iags5
a1d/xQ7AdFcliLSqvxeGsqTFuWK90ESbGgVgcIXOvDoqWJAzsTg4V10ThoHL9nvh
T8cvGcfdgV63fmAY8e44kbDL17bXgUNnQnTlYJI6rCwNRMDFqgWwX7TPcrJ4L2nc
XBiYyuKjSqBYzHVH9AMdKtMlRnmO4imURJDdbk6TFPyWRwARE9uUICbBOFHbDTLY
uAti4BBxYzZycYMxmfcvLqALFIK7gcVJ85UDgxyMMJ+TeK7+ILS0fQ/Le+EZg56e
7jQgBK9b/75CtGW6L9+SkVBdhU8HIbtwMB2nXLUXE4/QFpbt36TkHkQ9BEJeqqGY
QyMbc40vuY1vRGoNNTSonvfKzuO96X4bQZG3dkdZe9OVBpTNcuctPKRdOa08yb5k
dppjiWgfiom3O25jipY+VMaR/SF2UiAHvMs88/39kj8EXn1ahNk9Wv19K7MoluTr
/ixdc/z9kQHR78Vbs11mJDyDvhPQnX4tRzgYf4SJpcwniOjqvnaBVFJ5awiV7IIB
d9NeYP7hmUH87+6f0ROxgpncJ8JJWl/KID5W1b24sLI3iIDNTw2udhCiy+jae+82
kDmJU/KjScnbayOGN6SE+I8zwe1wbMjSIBC7JsPy8tJ1MZt4srVoXzZQMdxczUEt
k529pCBC/HrOK2yeUczjsKBbR0wX1IWpFiXM6deKoKVGZyEKxhBB5yYVjO+VYdJI
hjwUT4qPIvi22NdWK7cfGfENoLf9N5gP9c5D6anHggtt59VS1osGMeP2OGO6fTar
nJqCK68GWzsztlyCVvfQ6Ik56SDHptcDjWmpOTDENmGLcYqmREkxGUne2t0/K1MD
Bf+Ib8R2QG+qC6G09UumX1R9ys5zpogzyI+3ytYgaNYNtMt8WxK1bIp0ari6xel0
BfUncSylydFzt5CsPOaFQcQMspiv+BMDpJzhogaHp1iWPzA7s0wF/8SqbtY04ttv
irZgyFSwHO/GMipjJ4EaL1Y9279X98RcErnDDyK22EYXymAxdk+i31lyqo/ft3sT
lOyLeGzJv+zu8Xdl8E5yS3uXVjQPgtTi51vSJXQPLB0rgMrFYDaMtBIjDXyVVAzI
V4Prz7QjNp4esvV4EEhFsAltSv5QOKUNygxMB1Klsl6t6qcEkT2pj929CdSzBukh
u88Mlhnvaa7fHbPo8ATBrTV9DgVAZwLXClzWmCit9+Sq7S9hYvOiLrXCqpCYQaZr
bky68VOdny9hx910z80Ex0BiI9x6PExRQdZCvRYiWLfyWvQRHZVwiJ6P4eiTbLah
WlXtOVHioyFhu9bEgRM6JcJOPlVd2vygqzoH5bJL90mqXvAUtAQZZNhxvB3vY+hh
rMWjjHyALccSc3zHX754X8WWvSvrAmfOolz2VBGqf0Q+Df2Lbpm8xnE3DgbVVXVp
wjyq4l6nvecGOXPyfgDyKglgC2A1L1qJogVRsWwW3KskTQCAWmTtYmgEuWZIPX5m
bIJrfn2uzFFWTAo1LpjG6/tMRKp22kSB+1J826u7xGxZZfmCcMKwlVzXJ7B5RBSh
QsU5WvPu92Z3x8IU9vs5ZxrHk1jiWpJXKWLf+pISMycmqgovq0z/6mFg01k3Qk+M
JIPtp4o+42gHiUD+eMx7HuulaBv8tVmW0sySif5cKHl9E8N53Tn1OK9ZGvXyUVPR
buG8RmMXtDZayKHJCDpFBg3fKYMWD4JKHYt63RGtO2S82BvpWFjncF8Q0ReRZnTd
nCeK8YMx2lFl4Ank7IkcqV95KmL+Col4U/PmxlrpGA2mpr7V99kna+6jfbm92z1d
M0KIRD/rsFN9l0gR+oNpklUl3Ly5/OPT/BybKa6EctxHnh9uQ19G5QL7aoZvi/kO
pudsEuSzJHMddXD+K8qCRirlZFBG9s93EA2wWaNsnRtWYxHWUoL560esBAVTtobr
vwTxjZfPd1SvGqFPc3R1pC9mDoJwv4vx6sbaW/hZXcehVXcRHi2B2sQxrJrF6LQl
BOyaxPDxpko3I6GLkan7lR7GeJD4plcmrV5G1XECtOjV82PxOfwQ4HZGhiIdH0r0
1LNYY7PQ7NGl0Z57Y02OOMjGSbE4gdMMgS3lHHHa+KE3tmpMVQEDPPJyKR87ktP9
WPqqKmarjPv1DwRwdChr9Dyz5UDZnhgSiAXo3Zdxe2qa6Q8vPLVWWoLQYEsD7rjp
M5Iwx6OpokAvEyT1Vnrmqwt6zYUEykviFzihksuYd+RUzs02mWOErYzsZpMYnc2c
X7ktwwV2pLZbxD7f8Z4QlOYrtvO7LcGagIRsjCNyBlpxsWSMKtATP002jnZ1NJOs
ISPSFBlHf+ObWKFEWw2WiO/2QT8lJv3aeoLneNsgjqVL8rQUo2LLkL53TTHGZPwm
mQeSjaycI6v75svHeyTuVIc+0HXD8u8oKqdPbDqlwafTVRZaNHL+GESfjWVm5Hep
k2AyU45/Q9MVo7Mqv3kUf8Fe6pEHLfP6kJSB8kqdsYDiLVmclGFpEKtOfBVns19J
NXCcterO+flV+/NrpgBAVhgAb1bFEb0sHCIcZeD2+xszFBfG6kTKw+k/5xWfEwrO
80Ibl/bq91dsNKrHK6KMxy24lmWmki9ohsxJpYWZhmTO+cND/UOvy/IG3tGmZX4z
dI4Hns1KJnIKJugqVf3J0jQZieehQgBZIPP8x9bp1ZuRjxhfCHVrfC/uDwA2w6nz
68VA0WtGwpx0c9wrDc242R89tHiOoUWrwbXJLPNKudYlIhjzFJHcuqpeaURSBAAV
JY4vyxH1f4smYVR6Pyv/lC+wYesGYJAWOOND4j7mXNFHo/x90MDzwaE8PZIHyjAS
9x5sH0YDm851eCElZk0P3KHL8QWpbWSy6LUkiRQq+vW6dgXigeEU30+Fme2231qX
0oo3K9E4MJJbYL194+MSxH2FkA4oKkuNW9uwvcO78/fcpegzpVeFNJ/F9JTsACpx
ROZghYjPioEk2rTOlj1/0FdMkfblfVtvDhjrtCQGegXGlFdnyoW02/2LZ583ei5x
stpJODA7TYuSialgKJfF7r10oGQrvu6jOH+8MudY1dqXYfLRXD1OMN433v/HU/gx
q8vAD5TCk2V0O2ZqAk/tZ48lG+3KQqymnps1Ax1VMdgyX2OMHhwBRBHRftjckQZm
heP/Ko2yXIaDtQrfu9GEz8hebpms2Dcr0vYYVlZis5+gX8M0UxuGXXKuey2dYk96
aRjKwUSGw3uA0l5uTz9imjzK/0ENV/693SY+icZFogBv3UfnV2YmxYYOVBUmqKwQ
7tddaGfLi+VyXdqZ7p4wTD12HIAHanZ1J/t6+rBfd9kzOPuj7I8B2Ox+QRks3Eku
enii9yW/wWDctrC+Xb3spfPK/M9GzknEtpQiIGaoBU1Uhq3xADBjMilHo+5kBvHO
NuWB1llcty5K/0Mk2VS5C0jukh++KfqKi29VgbagXObG6+gnZFRQnj6+fS0bSsut
9P6S2jwCKyNaEHVKkzABGnhIeW/Ui/Zbxzi+qhHiLUGUW4EM4FBEW7mWrkrTclhn
3a98DMTytzavWb3qcdef+iOhH91eHrCTnsUJ9I+KyXXorubPD1FIUKYbYZbai/le
ktAYX3wpzazIz2Q5dNwkSret4uyfU8FiRiK0z1EK+RuVrj7j4MgSvCiED7Vs+G3Z
rvjs2BXxZq47N9IOhHXUeEVxHpEGaVTNLsdGQmFHWOXi2iR4HhMwmmO2HqfCafuF
AZEI09HAMTzJTOxyq2GOOxHR4Z+AdlAQ6FPNQ7bFkcvcaJkAcZ3DHXyYIrSN5LYW
p0IFPCg1CkHF7QINWdpTuGtzMkKji+SHMKFDnIV2ivjW2vln7CQwVtujYvKtJGi+
kyMGRko/Ov/RlAIIyiTBaFysrkI70r3ptnms/L7vT/OSgwkWbPQpm843V0qkiHlA
WxKjNMUtoqK47Py10YKZheR6WFa6pDwjX33v/jpXxegFJBNh+D44PgfT63ckY58B
9vJ0jENsU6xPe30YJG3cPASyTiWIfqL+7pdY3z5qwvJ6xbHix2snr94bil1MiNrh
8jE1FvL0iPXvtsH00dTbtNRFepJN41eu5wGGpMYHS3NyiO1dvXe0mqe9BE3v9R8O
cggR43Z8TLa3birsLypjeLMfpBb/qYXuNFNFfmTDHnMWJqPIlu6YS5b32Gqk0Q7m
1J2tBiQv/qjpkYA9hwzytEOpl/SiWYQp1D+Et5SmW3GKGx9Lqpbknqvz+UFb17Zz
MCVkf2Wr34TAEIjQH9voaf4/73zEvBKtBBSA5XYZRoIix64ZrJyUJpUpqw35kVeW
uxVIsGrC13ffFyf3RPwjHOx9UiuAg7i0D+7jfJR+uR46hjTr6cB1RH9WTjeTi/Ev
f5IzJB4TG9m/IgyqqnYYIYxBfBgdGGKzrWPriYPpxSMh/NGh1OLEF80AQ6wNI5Ee
5aeCLO0O2RuVDpwYXaOd46yZGitkVlvT8RML4y7nmo4HeP1iygnw4gW3fd/k8uJj
82oxRYXpjkpgjT5ptPeDohvFfaJCdjYcgT2UbfbHGsyDrxog/EA4iEjr7Y4DXx1E
Hx6wDzO2tXbN9BGe2Uvs7fFPW+YSinHFz13sTpmzBlCurSqLCL/63hbVMReo4Lku
OwJ3+jJw3xfGZgw9QRVtlE9Ui1uqCZsfeu7maaYlj1SsRpk2/jX6XDbjHbLL9Rh1
S3nF/0GhPj0H/XEiZXoIClEeKrQ0Dp3U+sXBpVuCRWU81iLo14LaXbOa/4j37vfw
iWa19SY+uH1qZy0stTum2HJ0JudvsXLJBMf/XWWohgs7DkAHAzMAK/jp2iX06/4I
4cYmQkOe/l1fRta7pdfO8G/M8P4vLksT1w/TJPTPAQUcH1phMeh5X3aGX6TmN2E1
ccRi9LKGXCwsLWnME0burqUqQCQ///JcXzfku7l8qVqbAIRCZcbLDy1Vb59FQH2d
z15znpUaw5hJk/WhKc/z48X0o5ASGceADWXkbZ+GUWCVC71q0QHN5SJXP5aq/ImX
D1Rgj9ShWQo61E9afDn0JNfQKUxVhcKzwKRY3z648rb6NVb9AfIUOQaRjCTUsZNM
MoxMUOQvY3EAwLznWzvjR5ytZOK5cKavlPyM3zyYLDP+11eLcOULfGDw9Grvubv1
r2Radt7RKYv5rPWbdQzO9HWhyd9KBJeOjc9tZ09kL8eJXschcyvJT4NPh97DX6Lm
wZEggVXxzNTpOZ5YOHlE26ZWYHDf/hFyyamWx7CCQx+25axaYMFBEHz0W+AIB80f
JKeDpPPkX6UB5/TvcDHYogdS9cPFdPrIJWcvy95vlFK+a9y2wYZrSupvMfunjuBc
B8ZOf5cS5kOHTjgsENoAEFl+wTiRWpSdD4e6xAS5g7AbDIWMnDiCfzxX9w37e+UK
ZTFz/AG4WD7pNWlzKCNISucm55yRoO6AkTF8z6nohAisk3bPFusjW0/xE86Cgt5e
Pkb/IqDQDFlah3qCOWs119nTH5qpH7Qu1rp4vk6RXubt9aHiIGjxTF6aXcX5uBkm
XVobqggxTUg6CnfEXwl1VbYTlfT+fSA081+9K/TuLbJSRcHfzh21gXyqJN9xmlOB
buzjPQvsMRyWX1Y7JuV/qhqecw8EAZTC95frLHRXt9atYQBoiuVRXiLXzzx8mYwN
RgWtdi4FWoNFyTZxRGuuSNYt2wsvQh1LPpBaGk7S88EKX7iyFGGzOgaZJ87xuOvD
PPwVReVjihRDO9AxOHuZzdXmGD+uzIu4WoKUz9z3x6e6FIRdQddIkUBQTgsPGz2L
KHKzLKZ6NRn35Zne6x/dXzAvAcZke18riHHNL5tfKvrNwnj5wKHB3UA6qTTVEx2Y
M0TV81aCnjLPyEHgRWhE3Mu3FK5Dxhx+iVKcoFZWfX0tm68L3XIMSW8d7Cf896Zj
0Z2wjrZgPQIyQKOeWtHsAZC1tcVHt2rhhcZUgB/h0ypT0DXSCh7HeuZvAdHYExhB
tfxJkKTnwpobVRj25SytOZFnJ0RS/mKLsmCJNpBj6ELJMvq61AYv33oBPbYbDHZ9
SgZKVuvxrw7ZrH4UO9evcV3cUhhSqsQhgaxHnaKDNCuvbT3CXMW8hpY5pEGxtaWc
lZbhJ/rwL2HLSr84KIxfIUHF/42bQrcAMScGoqSzWg10eSM+GyfU//5jYsSja7N8
Ge+5esDFiTjB5+Fr4lAzjW+JYOb2Lc6FSmPLWJ71IEwfEzo7Hq4rEKvrFWottxuh
Kg7zdVy1SQZDz+q8Anz7En3x65ICSJOmgW5xBq7rpdk1uf3GPNoVbaxysKcmqSHC
gwVxJpmq3GSZnBLen4CdVsiIYzORRMbxGSk7BdLKxg+r3zCkDtCU62dAlW9fIwG1
wpO3ycjvzjQwbxP0pQhCwJSW+2jzdaBmGZv+D22h3Wt4LfDs4a2/DfYS476QAh1a
TswIyJ5/Se5M5zKYQF93hFLFLIuz3RuTx5SMbAcqyL49TDR2DGcBggrxpQoXR2z4
F0CoyJRScHxawVj3X9Rj/TVOIO4GD5uihJDZtR+OUKmKQ7D4/1RnuuMQkeTNU4RD
53Vl7p7KqLtVG8wsnDmTbkM5urlqud5wDHC0opWRFxZjmeD/RF1393h2BBVkSVLI
QLXfdBR5PzIxKxQknu8RB2GvzhAYXpd7VlENy96SKzigTQOV3FYO4KRdCr+zUi4o
uhOwaf5Xlkcz+Z2qiqlio1t16shtiThkX0nydwP6Qvq6B52D+D9G/Vm+QhmtCn/h
MsxwIslzsaqnXt20HdvJ9fHU5AZk/jgQPq063uNANj+d4IjO+8fq49uVZfNVg2Gs
OgmzR2sBa0XL/A+MJgKxIqwgtZG0OS/ZPZFCwOD42LHgW7YglYWLO0LFNPoIIK70
l3SAD5VLwaIq4kVnLGTmkuoruh7EdG48cFxeL4jveC/MMQMt2OdIXzFJ1p5uJ0gK
E2kqMy6niCdqnJorM9kDOuNp2DaBxa3EAhKnX7ZoA+KPJquGplOXPPwrH+M3ThIO
KBWwU5ySnDW2YuLbE7ADFSO7NWbgrQis+QcRu+5UF5NlEEo+Wcvt7geGdN1iX6Gy
j1eIEFRdySmq8y1/JCdsQIXPuzLFGYwnNkSSny8mzfj+2wprTMN57HzWDljWCDTE
KhB4qcZaU4j5IIyIMTSSQq8qcXJBQKe3V9kIyg3L5+neFLaB00Zc6O0Vgh18F0i9
bPZ2hEgnto//d02gtnlBmRm5HnZNFfkNvNwKhPZ8AAazm0dp+UPfbnwsh4Ap70Fo
NK/u/r/koOmB5d7hfR0j0Ezqbk8ueeIFgK112QI6jCX8Hbv2FFFZc1zkIN381zrg
IggncDWKIRa5cp2cM1jkQiVeeTO7lS6JVuP1gJi2ORwE18GUDZ8tqDu+lit1BmW7
GrQZS1AbkHmmXbEZk1VPekDvZvkGxidQ1pAj1plrGonGnOkFFnkS0CSUQaJtb0A9
BAec/6OdbqVJUKRDOFF8gTdfq+CXP3b8jTooJCuEixRu1FwTGS7Tqzw3PwF+rVaI
iF4Op5JrGvBe/1HQms9HYn3dwcj/jCuF1coEZGy0jlt9zdw7rRpilRUA7EtBzpno
W6M22JHxI/P+5T2fU5G+/FJfqIyJhA/YB4hSROip2fg/ZThJXGl1zRvjw3KK0QOZ
o2gSSKsTze+uOuFbuqaxyOinyGR2r4uBFUERTe20sERAL0Sc5ETgxB1OBovWpRIx
u9pUGa7P4+wUTNM5DsFzTeCo8KRMURrlkBfJssLJfSpnaLUEdsyPLjmcZqBUYg0l
ZyseRx9fPARcHXOqEhwOXstOb97THgXZ8zV/z19O4AsgL+VJaZncstiwKTbrG0du
DnWTIlw1ht+zY28SlFKdbeQZ5hFVN3NTxPxaIVLnMWp8lHRG4LIGRtdbpdj9kaHm
ViX8s3AunZUhcuoHMk8h+e+PBL0yH+PBbZAzicCtiLEapXFWRhsgzfC/b3UqxSm/
L3IL7yuwZuOPdSxkP5tVSqltZ7Bn/2Uizy+WFA9cmWMQKoqajAJ9S6Z0c6Rl9YDN
bN20YtDjhOYG8cZ3luJq/n+1LQBBwYg05lz+aK+3DbQjNpaofEG2to/YSMLXe66V
rM7EMuJP3QU0/rjRqEkaT6MLfcLdwdzWNU32yMBjPoSB8wWUkpNkmbYqxwqBbZd/
/aZoYigHbNNwW7D6RFsD/m3BldjQORz45+1/cL6H5NJ3VL3ZHd5+5lbpdVpsUX0Y
qE7z4xdiS7ZNRhoHKaMfovffkwWDQHo21XxdLGF17Nhc2NjCsEXpb5nkosRX4gUG
YmfMtWyePs1kQyEVIr8f6174ExiVKq9uqZ6n3VZKhYhiBXX+8Ton+D/FA2XA/a00
w9WqsUn1eCqJSq6vLBk48r/rnpmiBG7Z/i1ehTW0A2PUp1fUxMTdBd01RqvM3+l1
Daw4AUboKj0SE8vEN/zZRvbSOB5vT868nlAdBe/tD1mL8vYlHZc6rGg3eWJkj2XR
Z38wUB+6s3tviu1ORExBVdWKBhhxf6duXeXOVm0s0Xf7yK4KW3TIsiVArlAz6BWi
UH+eQm3ba2u91NSE+NhxrC+a+rSy9+aO51jJKQ9sk5MN7FzcE6ZIniooulyJ01RJ
LPEo+3UYDIIT1Rnq5Y2MiKMVzUBiUHUPgWBeLoniCI/jeZLEkDhcXQ3MgtTrZPyE
LYkTVeB4sOxTVtmpc16jmiUhy9AVGNSp3Kn0bCZs+PiMmRIPAbgoDZjPeLih7jfU
t6ighD103W0EDNS1+R81dOIsjK1eN0N2zXLOrJ1LTLGw4QVLHzT9UqviJtZ92bG2
a/ADuqK89OPjAZvT4bTPm29ZsOupgEhm69L+pdiaFeyUkZVIPCmNKPBPbH4HsG4W
RwU29ZXp8KaqEp4oiZI0v+MSDM3OTcTjNAMsRxGgU8T3RTfyom5H5rivItDdZsj1
MfxN5qwSlZS0gIj0+pX8eMh892CQqiQGf5yTtGW8H/fpjQZ7TKfKgQEPlZbU9UYy
RCOB/68nx1zPsRA0oco4n1AuMRIZfaLKiCc04o6zgZxkFGpU7O0zQj9CLxy9Kplg
Wx+46hPvKHkhU9MoM46bflwGF7O17ZQOR38gY93R7JJ9K/cdsTEfvP6yGlm9g3iW
4EBJXb2mkzJ3zkwKL68U7Ht67R/KoFGFYYYAPW3t/bDl+q4qgNgWzia80MG79wsd
3TUtPdtOaUgGQXgDzL7qnc2UHuWjnni1WKsMUwimO39tKbUwIv0dzYBU0IwnZjyi
BbApBa32Y7uisn9Fv25SlzZQcKzwpBGmpe1OUw6BFpSAF5N5pdpVRBu/fquUec7v
oLPhH0lJPLxj2Dm98SeHBj7aWvcvDONr9roq4CxEFp1HQZbInQcxtd8hwr/Uhmgt
SueVd2WN1SzTQYA+L6u7hLhgVz82f7cPr8pQu61yUCr31tNkQiGfY7HBITJm8bp4
Ic+oGBNhwfnkb122CFSUrJ9uKU9xjNanU29ShZXVRvXKujEaVKjfNGgo0kmToCsv
LmR1OxHw2ORDmz9hW8GgZlEDilW4Tf5BZ5ABeWW/2zBb435QdMEqNiObaVTpeinB
II9mWeD58i8gwRGJfZR75jKqoX39JUqE7v45BzlWqoQt8jipUh75ihXFULLaqER2
5UnnLP///eqKtaEBeqHYG8t9S4MVWus0lKO0fWS1BVHhtO46OeyzHLwGyWlnlIRf
jIo8sEt7Z9X4Kgf73cyFlwwpxL3SRHsX6BpXprPH86zgzkuWcBJx2gN0TXcT1lu5
H6ttBGINRIvRyxW04ghsz+T9Yxj+ZZ5UwLiow4rPBk1erSMkqHA+byZHUkFVIw8C
NecZ78kc0huJ3pUnAG+xgJvd+d1ntYDcLNVJWxySEZoPqJVBddhhPxwNmtxvOr6A
4EbaczmQKI6grmqZxKGOgphIqU/uLtvym6VAPc7MxfkqIInZhZu/H/xRz7fWPAQa
gSkEyl00h0BBF7kk53TszXC6dlH//06z1oADgmYTo404IKRsMzommJyQ8P3ZEhXp
nC4wiq3O5FiSbBnCK+bKjnkAN6aUDYCcKa5ROtSOVLhypT5NODJZ83rk0P3v9FDQ
pJ3qHrR5b0D0e/9Z31X8WtboEJTBN14fpe3bGLWPktXzZG5sd2OyUVmvSCX/mrYo
j8pEWCEDwisN3oQCosits6JaiPTitH5aTt+ncZEVmDwK8zfzZ2/liV9UAUy9BNpN
EF1KoL2siI+ooqnRwZJta63sVMA7R6n47cs7Zk6/H846NCOBL2ukjpkU0nAyKPjO
iJmwY8kn8yU9s5Rvpa2w5UneQ7f0X1J4qhaJlanUwAY09Nf+obMg4jdFGb3PQWhF
LOVUy4vZSfYTmWRwOD5Ijk9P3Sn4wArkmnN/UnwZ1zKYyeRve9wZAXBRDifljSiv
DX92IkqZ3bbj3X7wQ3YnGS1sILA4SRn+7ADeve+cq311g7+pzw2dmy/gIQbswAq/
pwwrM7QlipNnsYIbpm+kw7rkAaPrhWAkmdeeFGHHkCQAjsEYlcZC6BfVh/Wu4/Ju
YsFK6OKAVKv2P3bOnN0GvsseZYKYT4zmSmFK0RydW5Hn9vnMJIpscjiDOUNHtsuQ
0gP+omRwMtHWIgPbcH3byAye78ezqGZ5X+S2cxZUU+haiXvyNBQt3cPlT2hmtNcp
4G5AcVLtNdzX7VAHkeUGrFbUS51aUz0yK3aMGQMQcMrHcHeTQaKHZPVy1ZIbaRA3
f0T+GXN+ufeQZuWghiF+bcDGwfx22lfkh8Jd/pQrGrLsIZEa/jmYaKP8iEg/USKF
/+u/tge4Qai8wTf17GZ5SvCNL6X1U1xxwackPjdHLiVNVvoU/TBGAnZFYOUpmXiz
kqJIjVKu8WcWXw9qWzN7H4N2Ip6m7RpjOP+61LK6anYwmf4eKi51sfNyFXZOjUKu
tUQFHLxXBa5mew2jfjL3OaFawevz7Ch8uFXRBDDPIHj4uZ84/1yMMcujiedEU/Os
AEdzPzDfvMHo3brRm4gqRpj8wco1yXO/cZ0Ds056uFuzsOfZAkBouKbsXjI19Qq7
/I/3slBiS78k7IOaQVje/GGvyhBTP7q2OxA3yyLEQevkfWCq21oP+GYiZJMoLdcT
v4vOgI5gd+VV9hc6VB2cwEOCBW/YbSoE4E5NeLuo7DYW+UlB6SBpT4tUts8AKJhg
M6HqO1y9SoeJr7x6b/L9QAjvQDB/dyZ9wVzZ2KfvaqmmT4wVF0SZf/aASXlkvkfj
LyWUrog+bOuPXqeuLIxkbzx5yD+Oi6rmUeayGnVy4FpUqp3A0XfxqZ26hDHjWKnA
3UCD+KOMlhZnP0nw2ZIVOuM+YhO+KQRHdMBjwCR9F0ki6J/8PEijj0mbfMrv07uK
7MWbWdODpz8kGnYRVA6tTy1th5LU2rZ/d94E25gb9GogmVso0mCcUhwKO5q7lWGZ
uZeBzndpdzfl86EYl6DRUpEosfyclj987yUuLwsZK4bj31PlnUWEzxuCm62QFrzO
esnWlqIkkBC1rzRMYfXYBaKCuBHpjNft/wmUasvqZwb7AuCSt3o/cyXaILRTp29M
C32jnXjawFcM6iQ3/6tT2EndVV84TUYCVJKHcA6M5FQTrg4pYbBSq0m2kaU7EJXP
qJP//h4T7KHhnTP1kLIcI312CUTpcWLH6vWvz0Qfr9DWPR7amACLJoL8yDs0Iura
5CGWNGZRWakuGBrtPo3KBlVOVd/gxIEEGJ8wE+YX1I2beFtCYQI04WeYQjQIbZwW
cno6oQazujXaRwpSCogZWv1XUcofH1B6ti2213XpUHMlp2NVjnn06ct8DvdKofzg
nudVFlzi18oCvHGNtd5ZMsBO3gr4QsHQlbjdWra00BH6mvhcnJAkJ6BA3aL3DUyZ
57VGCgXJPJoxqEj6H7ZrGkxPf14JaH4cdHFpMSOnBz2pWjZgItqAK+FazqkxnYDH
dD91y6P8gLa1E42ZcrH1SeEpL02XA3ajBzrvsdDPsIeYid6VEgu8onKZfosZ+40p
g+FjzE/QAQIqTXL6uso/vvgqXCAeeR8VOYlMbPMrrI55qBUUizHABxJZjmq8B+LM
Petq90asomnhuCJaA7KTSgQbJVi0hmSDXB5+Gg2afQlNX9L8q/vrRg4uR/oNnrsS
WhxJauUi5nz4V6M2N9r4JOdy2AB+sUC/Fm9u5YmZOvlvWmeSaABI6kutdyGkx0ek
L2DTzH44CbvVnjuPpPfrfsLNtnNvjIv4pi8LjHBWf06wJuj2vFdCxCdxhBvNqT+N
YnDKzEzhjrFEm4VOw0g92mhGE3OknrF/dJ5uBF3/fx+KGwymagrtKGduOQMu1MJS
xTDQCsUXnnOp/r+sT9ZyWMJc3As6jJHASOhuaozmYb/aZyI0WRmmDrHcug1M3/iJ
TM7N01o+n+SrgL+SNmxHECnCQRxqtGQuATJsj9TFSx5vTvOWXcGYpg9w3iysO5px
IRWsa4j++V6z+9NNZk0MtQ74iyY0czkiTjZhrYU0xVHppHIHAjuTu3EKrFvrWvon
5vr59ClGauRhWDyQnlVb9EBhQCA/05kzfyTPPYMmfT+tFx5K+VDCgjXdLaFA9p3q
bZLrvl1pkf8YjdikZcR8IXU6waW3rOSRRkx+ZnfnVeWsC5aHwPW4GYIWdz3UBnuT
6XfDqMjtXKp67dC708gPZ2dPmD4f/MJFsMoYW1NrC8p853annKLUQUAi+OaohpcM
L3eIUnkTkwvL9Bn6RXCxtnjbZ+uFe3g+tipI8xrSk32iN4im6VF++yb3FgakN5bF
AJJcVgx7XXzCFB0cZfqpN4NU5tEBheyUty49fRRVp6kAo+3qxrtIgqofUgYeLUi7
BSEkBsYh5so4BpI+8vPg9548e5xiBX4p6DcmidzzQWQ215Qex3aYHWvtOeIDC6Ob
t+x9uAAhacaE6Bkp9pHcQPWljXucT1fvGrZ/t1+F6YR1J45RPxMDBr/8hGwH/mns
HrgvSiE54xzCkWYFFXfWTCLenLOjPvXdjJPjmstbIb7a1Anc6NC5WcENf9Sch4V/
tluRgHQ3MTXck8MD+0Ywhn1s+19m4E5g0YVeQ69zRoDzCqcOf9POmm1G+1PID9sT
9Kf9vftzy4qQQV1iPa+TxTvFCoO+l2rvVJwMmnE75Xd7aHR2igBppnXX5Sl+s9M4
Nk5gIaF/aPeV1LKlK+j8pMwf+H2VXhqv2kSiSnTc7fa1WRbxJwhoEzpaQiiBaYsn
OSWGfzEYQ4stnaR5yt3EvQjFPJw2e5GAG5LGyEz3r4r/RTDdariXVOKv41Du1wSM
bH2if5PXngMcRSCQgs2fjpCHS9PbkprLC+hKxqeyg217qfruh3aTteyt5Z2tXv3Q
yomHJdsqg0GObHz2XG5Y7ZwjfBLeIbn7VaNvF7GrZ1jgTgqU7RNywWyOy5erblD2
MKUzHmDmySsPJP1OLXT4J+h/BrCMiFtS2V3WfV3SPk0YAKA/FB0wrUPKygSbKTMD
Wir/+cdJ7Kyka1UE+Y34xEpvbL/J/rIETR/3OhZ2qIyuR85Coz6kwBA5Ow7hR5Cz
YLNPggQE5yXcNrWSz3mmIf6w2iREgfyxjaoKAwXfxI27MYAbVJVjLa691pFFxtpo
fek9zk/es6sMe/G4dxtLEXqo06Iaq4zeSkYEBEK9gr1RtQjpoZMjuDK6n0f+6bva
C2HsGEb3ASyDdgR0sIjNvDFT8CLafrz9uabLd9Dl9mIA0eaCNm3N3l0NJ62Z9Q8K
xIElAkmTGR3bwVxyYXcooDOU8T3Yw1DlqQVPzGrfWi0PshMZDBmeDpaIT3sF3Goh
pPiKvs4wjaUatI+Uq7se/fmouNIevZ6hau0o8kbOKHLzaXUWKsHSwxNzKdU9QruU
0v51qfxa6veF1KkUPYcyC+0483a9sOuTz66UEctU+uma9raOZ9eVX3i37yKiSd0f
+tM4VT2lpCxOYLTsyTb5vU0IRz2n/bhII++7rGdy0fEcFy2Fsbb0XwPuurihojmX
XX8slbf5qt74JYLq9CzEuyVuv0E5hu1CGrhEmN/jhqoD5/W2woV9M8xvR4nifmhK
hYaUnFLFPLcI2k/CQaw9K/Z9tW6QgEapSEu4kK5C7gDN9z9JZtJZo5l1drSO4upb
j34NbKxrnBBvyF3pm+ZLp2bc+h6tdpzYc85wepsQu//uRSQYHuTafgGpOZC6bk4I
7drPeW/lbxWWIqsgPddu6nf3SRnXoX1DZ/WReqTcX1ht9nXnR8BaY4ccYrdZtyQB
UW/z1mDobLLVxoo66RFsri6r4URxZ0bwE97QennPOGNj4D7zxnJk8voIs8iU9KMP
CVjkcGM6m9bU3PjYEdFvf+OfxvDkfb5HH/z7XzdomMaCz9Lh8nFzsnW1OQPqkiPp
g1xp3e74Z+DL3dSb0DTX4nJamjVA7P5bO7GUDB8mFkHeHoPNQk2CYH1AQNsS7LTC
rurRwnrSxmMd1qlaesI3Gyw+coGreLYgNlYEWLYL3e3/i4SOwQBkEHvwqeER/Tl1
TAxAVXpoAgbAm5A6jJSVmQ3IDS2UdvHjPHGD4J9Vt9BDT19YYjqaabnFCvKLJiDY
1rt3xHEZjSkuY/0r0UhE9GLV4XNoAMpThu6m0k9pNhgzb3bSaB+CvNzCkBgxnA2m
iv6bED/HyVWUm0o4OXjidpqIP4E2lmSt0EXbK8ZlPj6iZelhBdBcOLohkUWf5uam
B4rdaI/V5Ts51ZQ/eMOP5bTwlfygoQ3G+aCIciOjY7nhYxGE9gac6p+3EwrSy8M/
6JyEyI9VRsxQZw7Zo71L11Ab7yP8qy6wsBDhCB9GK4BffgRuS+/OEDEmqvh8mte0
ultaeyEkTlRIGenooTbpyB2LrSp7pz3gdAhmK71B30lK1KTSFzq411vCPL5Nv0BY
7BZtiH2qyyAXPErxbiw5o2zhw9DnB66r/tKwO30ZwmQYn3LqpBXF+cEnJqNP7MoB
ifleXx6OSz5YMg976oGCsyrWzPsgEzg2pLzdpMicvtTBEoLfb6H+bo57WtwRbU8j
Oj5xxmsBBpeZIjJ21zxTpJQTw7OwKz2wGfNGluq/JPYodpU9pdcojOrQ/UOCpd0r
ZL8cc2SQGgPT/kZ3EBHKjTZim2tQ3ONK5cwciU2DjcOLp/mv0q05I7XuEvo2QSYu
pL8qILF7YX5B2lTWnc8SfSBosS8hKEzJRY+t2SuIWQM3iiGpp1TZG+uww+OiY19h
g4MQHfp2rvnofjS3K0BhDqznx1egrxYKGAn/wPZFzSZFQtllkIUBYnR0Tf82vq+H
4TmFx5oGCi9VohvSD8xqShqcqzty8LGb63o6fS+887E+Col7V5WrR3fPgH9sBhdN
qpSRHUJTm0nQr0U76irbKsfLwOPf/EpWLbn5DCkmMhEOQm1Oah57V1jQ6xiFqCno
GUfe1pRrFfitIqWf7U8XcZX0d/Bn88qcsWqesw7U3l5ZqTh31Sol4u2eoKTdyHsV
f0D3HYHQyNDeVq57MAlCEVOfltW3OmP/8uIYLlvii5r2E/Wf5v2i2KsnU/GuMAO+
W1y99qzT/kl7eh4XYcb4p+bGKD0OexKEpdVA0cdtLOsAWeGzg3sNxD965Tnpq0Ip
iHJemKacfYwmC4d+HOztF5jX3fA+9FZmpdJA7DHSIp4e7uAn8l7Scn3/MCCawtOC
LoWMK/Wf49HbI3Ra4Kpntsi8CdpREEWOHoT0641KK9iANrx5y/IOOaVVW7GD/cbw
aVXdXe+Rv/o2XeswXIxt0Ya135UMkqwn3xiWe0qxTV9FI1tt/SJyJdpU3zvEM+ZU
vK65zlJlLQGlFDyW/u7ZpU3VCtd1eFZdHaQlEc6x1mZ0N0HTSOwpeHywDXrtHkLh
ge1WJN8+y1XFpmhsOyhRVZixgU1ePgZeWCELQjvLHtncB1NMMulqPrcGQv8y8Zsu
cOVDv7Bdkw31b1vy0L1fpOnZMu/WmbLrV7jw57ckq4b91g/73tPGWpGuZKda0qfl
vpiNAYMkEYMEmeY75tsAKIA+tfJG2f9usUhv63wgQgacLNywsbNh/19dgcybhMX4
BDwSt0vA4V0DS+fzB9uP0mfkTh2CijQFXpcbpP8igJRuH16Q/sEXp+ymr/H5vFKC
a4LOhqQ2mNSpBgImLT6sUfBY1DVWTK3QFAFdgZk/lZmETUf7EeJvxN0Ja158KeLr
wpWf3AkITkwtCByuYLsAl2LKmXX6oDKsoCwotLKF8Gtm2vKL/RlyW2IKFwK8xjxV
eUbXPuh4aAlLlq2a+B1othOZvmRq2PLKsoUECrFmDus8fsSqsyS9QH/wk18v2quS
g2OJC5N2ipapLy1x280RREeVQ5DoGYDFRXANXz8LCvmRYUHGMTTZGhGGctx9VwHj
mqxOENtuQsBy/ftB0EKgFlo1GcB+3ss9sIekEjaSMsIoe31bvNz4BCKk11SYtGK6
AwnPCZ4wPhNYKwAQRYR9OutXvG0TTqExzbcz3wQ7UKPaTqJam3a7yQbYH9diWBMo
ywsYUgctYaLFoz5ajw/eCrWOkPUnDsNl4GdV3/hF1LOUabFSLnTRjr8dXtl0kz39
+XJ8OOu3gonS5LIHvgwjKfE030vt52ykXS6jgasDugRQfLD/gy1+aVSY7AmoOpP1
xRbINMmpT3iM84NpFRItlvhSh2cEtFHwlu6rCsG2V3p2vQMt00wr4wtHAh2gIEoN
H6xc7bKu2bcPN+Gt7pltTi6kdsoAZoaPrSWoP8Z2BtlYiNe0laZ7/vQatE7vnWzZ
WdYwXL56vkhSj9RZdkp/+c/+fqecnLclZqBOpiBuOfJpB4B+yGXcE2fecyqeNZ+l
/ja7dcFsA1tnGBa6Xis8v1gIg+A2YBOaXW9UFrPOropIG3KAgEw5f58OAkWOfjoZ
GBCWrbfcH+8vpt0gymo7lVsRodl07W3QH1a2D4kNmFw4dyjG1Qe6T4TGSA1OJg1o
LbjSLqObBNQemqOpB262JYzmElCU3/y3NBrHX58+PyO4pX39kRXOyBqfiuRpw5lg
Sib8UG2BkYShd/8kNkE8mtRGFG9wSYmZqYr0Agc7yR17+4loqp8Y9OgASEEHV+4z
k7swEfPfJ95cJ+P5pBcbEgmmrhtNH4Y/4xlezIYCno7LzgMjx1LW8XHtWGusiT4D
HnDItYPRvSkZfKEMcaaX3ZqW0dlENibwyq2eLGXzV8HJ6+dDzmfC2mRlyLbHpAN+
RwEtf7RLnYe6OOmHleIbiRukEg7blh1OzDEDVVPmcdtaz3bDN+gSIUiCl5jJB3yZ
5jHtT+Xca53TPc0s6GXDEDxFm1BSyAjHY5FSmVXoBnFxJDYqbfhrg4Gy8YdCtKqp
UrQwS8T50XVNWZYg2Yq/CP3LK/ibYXt6o/bHaqVdMMFarGr97QXJiCjw5brECmVg
wR8Eqx+FQbW1QHdcC3WmmMsHQ6CGeO9fvM6F/X/QWrkJjpciVknPjT88wZKA7Rj+
s1K2D9Iobzgi7+b46QnfGUjP5ypdNJLe+YAtx4F64iA5buMWbq9IzKLjOfEWsA7I
66cupsb2Zf8y7fPrLxunaXvVFcp4g5Ji/BWrXwOsUOrKr0xM0gvYC59U7/eegQfh
EFoJM0xTPQBWYgvy3zDk2tJL45B2qm60/gndfm3GivBKWSGrTKqoK3CuuvjKS6k7
NEl6+gAVBXJWldk6eT8mOH3Syedw1qej0C05uz3QnNLwy5DBnpcnqFgc5JPpkvsU
JOUeyoCBYEfHo3Q/HfZefRshDROlPpI91TKZcT6ntrhP54obhahDp5p/wQ8MB0/Y
u60CMiSxGDmVok320E2Nc9MXFXPXk6mcdyZYsNa3tfxaCCEBDsYcDDdL2BVI4Ngr
HpMnbPRepAfpXoiz6f71ttImhgdcwAnKt/R4/Y2v5OR33vTMwNMdcabziA+mwrXe
5C4eJHUqzw9H346COEEgCdXQJ1jFk9K8mm6AY/YQdyxH2I2ePeBImRk2bE8vjOm6
2ymPMFbXzv5/hny6Y81qU0eVry1iQusXQmnt4kRXtMQIHVFMSsxe87vxgn6mbv+P
V7/dWln2b057VkI6fJUEZSuEGyrdHA0dRY3o22tlgdZWpePsR9cQUxfhXAbyBS6n
cbmAzUVdikaaImDNTzxNPiy2pgPD7jRyZP6H2PnW2zfARTmYOiJRKHqBYzfZSPem
PL7DdLCYCfoJdJR8yJmUON4jud8d7FN8X6U0XO4GtztARbBmYslSMrv6fESp3D76
K3Ywk9LgfTLJ2/NPm7dH5amvv43IpudDSiHnp44Bs/vKk1/JkCyprWYXcvkUV4/d
EYnCkj4UR+L0qHbsFnotdskavTu8VLF+HWlfOwO/x64lCe/HDkAHG4L73W0Ol3hv
xzpGvby3a1tskBE9aRGs2pSm99Ip1rBLYlwDBEVcrN5GH8EmF5/1Pq1BXRy2Pzz6
IbePWs0WopG9a54GfsPpWLR4qC3CHiIZWLVSZb8pJiEtTshfB7gYjEd/bqUv6Lbf
p7RUlyAKalC6usGrvym/OZ8Z561YYdVa0UTO14Sng2lvKcoAtI6APk2dOEm6DOPo
F5RUzt+6TEfVKKx5+UorS7liK3rA/f7UqZBeC6J1503wzFh2wxXsGUS9SSaxSSBH
6kVhnjKF+FG4CKdN7U/iAyZwg0mEyqvk4H8FkTP29J4fQKEclyE1oRDHGKU31KE/
Nk9O9PN+vCHARL1GiLXUBIZH5lXWioe0u+mD67ZGtSxlxLNlVI1ogGjCupHPZR7G
V8CtR0FlaKwILmLAbPyFestQSkZyl2SfqNxK1PuwkYGCIiby8apjYagJDIzSwjtL
Q/363aeL+hUA277N4wzm+FE/7NcPbP5/UY+xfPrK2Fx4Xq0bFDgB9zapHN4FFey+
z9BHmf+Q0nij2lBCBIk1Ff+qc/Z9gAJbSnUSCkuFf2DWhFguWZITJsCJVFC1aVaJ
pIS1QVwVMzaoy7OHmtY+PTmqK8+KGPnd6pzWVt3iILTSQlLS3+vZHK10nxM+GjmT
r9QquT2tvBAs5xcmdxhQ9VVFRabGe2+u2aVH/4Ga5d7i5n1fsDxjTYdalXT8w48U
BKeMsnLmZwB7uY9ok1IhYHatOOvN1Cop0/Hlzqf8ZWFGEtISmDKabm717cVK07CG
bDimdZ0CbEJEdiMuZ15rrIHe+lUEs99npA6sFou5uunzy00lB209Q4Er7G8YKRaE
nrt1Zec8E2KRn0QSkYPKz+AAw+0osf6fKncdQfAMnrTPG/YpC3hYWKPS4/gtIzO3
I3+dAhbAHaxBXksmAQzbUbSKzg+AXZ87gB0yjM1wAfa+gxA5Y9eFAQASHtIZWI8r
lBg4M+EXrlE1L72k8UBf/wt2oZYsoMqjWvyrSHm1d1tgI90R20LLkCiBR60TmtnR
+7FCk86JSZbXOU6RuQuVyh9KWblx3UxtZG+lapEKQirZyojAvXr8uc8CwDkxkRUV
oqxiWejz+81iYMXKD9rGq4c3NPbHl6cEC/2XkoUjOi+u/nqZrKn8nEYvb6vHy4jN
5cKRhMM5p79z/zZIWaYks/UbozdXpD1KetjI0+sMF0qmfk+New0+gMqKs2ce4mrC
h9e824GuEA0p/VxdDOR1jf8sl5G341AGol80iRF6OYvO3tbTqYKzGT+s1EYkXbz/
X1E/21nYD2ZId0wmkl8mjb3nZbQJ855/MY6GPmBDp4X3+e4iMvviXk54d0J2AssI
47OdcALEK/7N+xQYEdnYB33cg4XzmCx3GQxu8KNLl+m2l8CF/kduRzXTEhjG8bYr
7IcAT81shXcMmy7CIj/IXhHEOBTXexPRWYbpkAVcdTB0F6EFSQwKKlnlvRjzNnxL
jVDRm9K1S+TenKAuq6ak6XI7YDctE0BRt5nf1FMMqZRAFhaNS8ABMkNA4Vtg8oMO
IoB28QK38WNS2MfCy+WUIPYdux/u5SkCJQGfKvDEFbKGszLQPUxVDmdruFVoH8y7
xvX3UpumTxIoBtez46QsyRjI5zO+l+k465f/EJwjNbqGw2++KodRbPlT4sy6YpTQ
EoY0LzNwMIE4MqpfZ2KtcUQ5xs80p/5lVsOCph4RUHVUmr45VAP0xV50FDVRp2ae
8iIFO7waYW1Pe9TahKFJ3pt7FeNXLRzbhBNJIi1BzB2Ml8I9NH/rOXx+tP7JwAF0
sK6rb2uzoCk77c4F5cohqqTOrzOAVEdqve64VksiPbSaF6heH1g1nZUWNYxe29XX
3uGR7nXkq+GmhXjMob5qo/BsMz01fnDuSa8J6VZYJ8skDJ+fNQc1vkYFI/CwfluB
7gQcArHIcywPdfBM5NFW91VCPNcJFEz1qK7vzffVuaCsl3DftI3Ys1ZNfXpqyMx2
ftVJshsz4Mo3gekQFsaf9kaUyPZj3l7bygwNWktPzK2xot/ahiWdie9f+X/o51YZ
r8sfKlBS6DjprDPmjgemFxLZpemBqkZZO9MkB7kCWFvNyHlDFKdVVb9vmwmobtSu
StRyQlHBNgSKphar/7Fqeo/WLfAZWzNTvQ3GstHEb4QLeFxsh3p0/2JOGti9BQyf
kVkeE6QTLBTyPIvmicSdtuwMHOTCLRhzaDCgKsPkbtkXqy0myBXCnEq5OZ+3S7hL
cuHdgomLYHJzOSCsMQ+SbMBkJBo9I5wKle8DkbdHMZdgqSbjobKjFb+vd6wln+5K
psZzjli6d3F5EfL29PzH0uibfJiZmbe8NyU6jiDXPvdxbL22TsgwP9fZ/bwaO8VH
xNISxdinI/jH3ihDb6MDgQoYEGPR4XUfcysKI3tZ1qIVRoXn7diT5XIMZuiY+g+L
cUIqu1lohFomKsYHC2DDpEowHrOC+lrdV21eioIlZXb23jpGtSWAmOf9WaF8jVlR
qcBYedsEytMTXJdyq2xiSfJzDASn5OxEF/d2YnX0aAdN36P7s6KevpKJW2vEiLvK
Wzxcxe/+/E2BNZtWdrWd108eyBaji5qZ2dC5gGq8FzX2zhCrguMkyVlNPEwYxzQA
R3iTSPIkjoBXMDLjCJfYO5DTY82HgEV3kyKJJNSUl0Pg4S3Vg+VEwm6Ub3QM/I1k
/r9T8NPf3xoXJpadZ4mJXWci46KrAd+F0QoggwLVgZUw8c+XtbvCvht8weBM8ysq
+GRxsP2RJYkoDUD84dYUJlTeXvl9izSovzCJcR8ppY4K0C1xYLn4kAyyzXZ0Mzv/
gkOvrCcJNshUqA5Qx4cthmLCO5j/tf6UKqaQJ9RXvpQIUqUTnuI/bh0P2dzIDtwi
c02wCjbJc8M0isSMnD3cULA6ymgbWqYvroxs8US/C0ZWUI1z+5V9P6qnRJH3735I
w/zOQkvEOB9lZxHAASFZHinyFjZXx96kdLTdTWaWYwIipJ0LXjNE6Zmx35FD2+cL
cMavXw984a3jIvwac1y0kJAns8aqo9GKudYJpEMlozIUvxnqEz6kQEKATyGRSy/t
kb1EhvQJIdNEtI8fqz5cyylu2Xl3tGAfY0zHATbzJ77m9Tt+ceX0+gnkdzPHetHh
AafBaSMwO78AYshT85SAWj1qHAsm0L9URmL7tdaLx44rojpDveme+YoZqLNE2a4A
euy54HPMe6ZQ+YINlc6mFQGrVOIgrdV9kR2Tb7eWFOyhvxm8Tv1+uHCwmOGF5yoR
Zt1caucMPjqOtelj85/MZ0CY2cIpfcISgZmgqPB12vgGLnyir/O//OA5p5kncVMN
eqBg/AbaBnWBgYUV1NlnZagdX6kFyF0es0f/hODqGf0t1ZgT3qyGfBFmZXAxRb5H
UHV869eqmSU3sXYS6+qzN2MYKek71XB2o5XgMaJoql1Cct8KCbwnexRYQv44lS/9
jdFjG0MEFUpsXD8St7tOnXFRaXM2sHcAHhtujG+8eb5AlHxUGVnsvTAG0hJF6CuJ
1FKvJkbYEEL4GUzEKMWRiom/9lHqvByUafXqZlsANCTqTyNZOi5ON3c7Xz5AK18V
e+tkX3T79RUE1tuTWGWIRxWgdF4nYguGcMbhcyWw0ELNN0Bzj3/gfQ1VAPPwyPzf
RuEPA14qC5K3/xJ/FVBGdcBH1rVRVazHBLDqQ/BPw7ph79J57Iju9A7u8JvBImsR
KnB8/m5OhAY6PzV8F+XOYzRh8E9BpePcrs01Hw803cve/epAsdzvyUvSEcjYkU6/
bbgef0Ct6gEhRgjRtbPNLY6y1NDTUYL3BZkRFdKbpfSm64NGvo17oy6258x1Hv8I
6cvxXWC+U/WdIAXZPDAA5e3uy9M3NogCdnyiEm17/RZgtkCWrkF1bM4yhJejFJ22
jkuBmIHDuKWL2+HZYjyXPad+l19YXOdwc75G+ZgK8tYjCCjM/GdwD1hrMlv+DOmM
ZGrK5CZHpVN4dFEh8Y/Rbi966hn0ZsvoBZqU5PJ9UQ2ehFA699ZhA/x4ZKFbAcGo
pdByq8zVBnwv4XbTPGoE8k8TBs4NcVZgkI794h6DVvc0vQsb69UarINXkhR6Bkmi
5FTwi1HR9qu9HlyOh6MaIPJkuOhtLze7nfEoWhGKxaAu3QAqtf6yqEDqjZvGQ5J1
LZwHJ/Ll1kqvz9nTkVFZi1L0jphAPi/iVJoKi8tSmMRClQyn87tggOUMpuyQ6tWk
KiyaeVA2pfuglIdWc+LF2FR6FBhh9Z/+nEMdXdNFKgdO1Z/YE+SLa+7G5uQ9y7Bq
HSJI1JLYrkvmMxrTXWM/ZICSLVi2BGw/j2CpOA+oBrpU2xz0HGTbJXyjsGvbfAwZ
29SjRagKOTsZx95KkTfIH5UuiAOJ/Trq1yp6t/lcg/4qUDXmyAJUs7r3TcpjqOTi
kLpuXre/PCr5x2+Ri1doF3qufXnsUgOI1I3rV7jEQ6uHShNWhHXCOE6KpuKAUops
BqR9cMubD3DBo59t8e3T+f+bePC+AEN1ujqRW1IAdL7DCEkYzpJCZswBfZfVPES6
a7Sp/6bMxF+QIHqkCou9wgLFybCSKocRNpMxZwyP7wlRVwY3bMQBH9T2GN2cGmDi
sKmr8eBr4wN4nwQ5iFrh/hKV5mzknXRIhedDCqjf97Ja4ACRceX8xSpyF/6aQZZX
GlwRPLJexR3PbLyeIdkcC+b4yAkjPz7b7X71IUUBjjHe0RDihdpVq6Lb/OdWxHKK
12g4wKvnNizBbHRAN6hAxBxzKZTS4nq06PQNKBo9JYYd8kqvQ9lfthOheLmH/Fdv
hvMkdu58tHNVmzakcmeuiC1iS+rM5Ej3xmJO/6LNEzUUigRc1XihyLLgv4m1uFzG
LhrQdDVWNF4MZ4bqseBi2PPS1QexNlmt4hYfnREauieVmqfCON/Uf1qfYC6q1q3+
nfB3NjTtkr1AKMNwMzJOBj7sL9r8GyT3jmmYkUDEoru3TC7AYwt1OWQdKFx9wnAR
Xq3C9ss5Ng0+pL9+sRmFyr/qeSbJ3eedHci7VjaY/K7Je4/yb12YMf4dXf5bpS2e
zvmb7RV0wX12ClTZKqsq4aPk4afflWTUDUd0K0hTYIjbBpUNkxh3M0hTx9/ZGT9n
nlXXQpUq2d/ExF9/CDdtE5UOMcRKC8zcSosqLgJekW5xEpNXkunJCdI69X8oY1XO
QEKfkRkbF9RLGHr7sNnaR1HPH8qYBslTS/VJn/PZ1g0hm4eGNshED+hkfDKMM1vr
DR2r2xun6rEPRTIaUqZQKz/Jfy8rHj2+78R+AzPas1i8aQtZdDJFBT2U9+bqa+bi
DY1vdXdpp+HCP0jW8CgM0/bgrBpAnXxKZtozXu212O5RIqPGq3YqHLPKiPSAJQbF
cb+nzL2lUB9km3stmqZOJXDeF9jquq5zcgRh36uR5LUcP8rklv05CtsitjNnesc1
bZ5c0ycpVnqny3x3xhhJIa0qo2uuGhMu3J7dDVlTyzOpm5Wa3bMZgHid37Y/8LGS
Qc3RFsuY2ODVxG6S2qNTgme3PEm2Gc4rECtrGP2JwKCBsHYJvP8oufaO5YjSaEKK
gTsZeWIV/lquCUibmPzrLrFxQ0QvZaTKphmvxYfmMhNO5+jc0+yWBn+cnojtcLZa
vCJV9uDETIYC5hp4tihex6PCiTtbgUxHWuM8zoYZsV0FNBhJgJbLQESJyKHBsYjv
DnmgJ78NJGqLosfH6aHzuuSw4PLnk1S0NXIW/DGkJtdA/cPrr2HnPpNOf3VKDC/t
F4or9ZlPYjPvmCmiXlw+oUEH9CKopq+5/SisMXubQJPS3reCGcoBvgwD9mqROBOB
/F5EL8NGX7dODTHKBo7MtlDHpNj8UCZKk9FBkMitEF+a6LwmpZz21EldIAusoDSp
GY9fEfBa48asHwb7sH3AtrCx7pQJNMicK2D5uY4T5G2P20BRnUaGyHTLAzQWmS9M
ZoqsdxJfAQXc+XWY5gIz3h6KPcqNMjlyIpign6tiWwUbsuypZogoiSmAcfTeXZ3Z
ofDksa08WpbRgf3zjRWiN/Is7xiY/6NNZpBQIxxDsdh8PCY55ESXF83OgSdd6DyQ
Vsg+cuo0BRaENsroUFvhqxcQ2KXOCfGkcRYjbX0yqzKNLSPM8Glc7W5etmltHx79
CeY7zbvCCbzQ+oNRUuA6Gt8wd5kNyjS/rZvC3dEU7qrsULFj9ZCkIkfBd3wLMhxS
wmMBSWKbmrFIG6SG6ALDvyfOZZNqXN5WMEhd8asxUuk0ahnsRIffg1eE/wuxxVpE
/V13XcN+k0g5yD/nK/c1L/7TEirJ4sD+M+esgS7OXdL3L6X5uxd8ASTPaFpR1zmL
NipeKxUOfsXjQNWF7rm8qZbAFhboyX1ByRFizZy3mfyfelu56UHXyQN3PXRzatUs
SefAfURL3e67/6N6pfF/3wOTY9NHfdkueICwBq0s4ACEzWGgn+BdNNOg+pc4CDvG
199k4B5AM++4ApbrZgA6EJJ6S75nQyeTB5FQUtzJRmtNVPdLDmaMMnz6KLHxDu7I
E4D1isJO7lH/t01TMCY62UnRKGjtp2YjGZwhwnaeTPnUBZaAMMKEXYk6DLocyJ56
GgmT6evqmFqNMIrLvxtIQ9JrhlFCjwqWdSYjwzBYDTKkKVFGMo8uNtPtAOhE72H1
O4EyS8amtc2wdzGMmMHHN3CGmc/rvnI7CCmD7+4gcuKHd3FKKiYfTPnv9ilZMbs9
XIfB1Buj6LAO+y1AsEd0KdkhBxwaQ2B1z9h57NIFeNgfzIm4edlTxw9lGHoxuLjj
zrDy8dZGtICovniT89SFuvUiKzWd5RtJiaLPILBoY+I083h/Gg2+AEmqwSD9ZFKq
7norvxjzL62jr33bbj56M+oseCB1BNX9onxR/ux1kzcZ5xe5IHfIvlSGSc64IDUN
z9TtmFia2vZckJbg1T1JNKvpm5pCc3uVAlxXGVdfLc80L8oeu1r4WU0QqAgN6Dyp
xq1AYEXsxPH0WmRNpibJA3rqxkhqbUy0djKKhIyLegRCUdIAk5IY9QPF4SjyIK0A
9/MXVrPot6fe87MNwiT9tJECOe3EzqF33hkeoRTLqSTVmhFuXuUlQK66U8UxstMe
VZ6r8XpK82TYmXUksoMIG3u2J1SB+T1W78At3t3kUbbssyxeYUHFwDH5djLMYHP/
BxF4JAx/I+Mttqw6vxCfWd5VD9E1Z1gjW9X96BGICyQCHufKZRV/kLT9lX+cbNvL
AjRYmldgouh2jARBfsXBbGU+0vEfq81xHO9jkrlCO3j+DHaO8NNgk5IbrQqjVWFl
OT7MRoP2SP1/MRicasRPH+NQU4z9fQO02QWX/JBySFD+8p0AYdGyW6ILwGYmaMW2
EyrdYeouur48k67KI0OYkUp+Nkib9lPWlQvaCJYSRkB8veFGLEzlMMcm3jv0Gzvh
NG/TKTlecacVQftIl9ddldknUPdINd+OyLtpLS/WAw7XJ7ewrskPc9EvkEqidexn
ijNO1ZgzRMujoJCcCQtobWjSuxYLCAAtbpcFEpX0IhJseARDWSpmzrfWXfNAcBqB
7zK8rEysyBRhUx9xV+GQdVvm6JzHaRrR6vtXuGURr8mruIO7VaZB7BVeQFWYO0RF
h8trwEnWUaa1PrckEMuqWTaiEWO2Y4GhG6X09q9/3Rk03jC4k9vFCv0+pIckNVqt
N3VsSfljRLLGcfAzN15poXnkjxuVSpgq4CZyBgK+lGygllrysFDl+aNj82nKfwRv
yD1k8fYRGkTLvVHpncpmS5/cs9YE4pWcYwmjKdsWH1AtT0NU6iGJiWMawTmVqZ76
rQAunlelxZEiq0T9O9Bhtw/0rBzXWmNyI6FCIx1gzehUizMzBaBrWJ+W6s4nzheT
F0hqXxJrJaqt8VaCpjEHjEhDcU879uqghj28c2Oqg9Czbz5vHFBP/TjREpxhntVR
qytrtHfu91jc32EIpRlEc3Fg2tjBfVupsqdKK+Pf06BJRee/m5V/g41oy/4Mh3lD
KCj2d7aNy0GGoo7jbK/8SSsJJIAKRWP0PoG9LhNQaFrlLOievUARgtTrijetnCqW
LxlsHqIhE6fBiK5FXVCgLbuJPQD3RVaxS/82O/l4ywgo6fxnwsWrpRzgSCCy0h5q
y7CxWneSCe4xCtv8jWexOHKoTRISB/B95lZlr4WK3YiygxNutjje6q+++QSJB37C
nsEfnWtEZ+hDs6Zpfz/l/ayZx6xzZ9RR5GALD4AUwhw3lmnL89uz9SfDF+S4nc8/
FWmiNogLdaGUB0rIVLjXoPji89zQckmLoqYPVHOoZApPLQhvfDiWEn7rpxrhBH/I
Twov3gCkc3lH1mav7edYhWlhANXTc7WtIOi/D9OEQCwltNJbbNcy0dD+sfMWMw66
eLHjY1/t5xQh9bIi77HnwOL+qiWtuNo1VaPyZBn5vQLTsvL1KybronGPv8SVKZHF
Ux/ikg9TT2RhJ6eutLeVlZ7MJ3taTZBzHiC/Tsp9SiNIifF4M2sajbtTZCR/G5GF
ZObJMRd1DRdz5w95IKtlnPbdGa+coP2EU9m8vbT+Z6Y=
`pragma protect end_protected
