// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BQlwVWAeC64OEA/03h0NDsyKAxQXiHCNtruh9ky3gLn1FOZyQRFNPsBArYlGtDfg
cAtuJnSNMZSZwYNwUQVv38HRm9+cMBTgEN0KV44xA51OmNTwDSlg4BN6m9XsMy2C
MVW8LA69lccGLmshKNuNfZs3MS9aXee1OreCxtXRy0M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20016)
XcyXbx6iQxhqFxkgddxCv5fDV+UF2Qxy7Tfc/lDv6EsnCJRJaTiQg7ZNsKUTGmpM
wqkVm6W4pbvtuf4vomJyURGok0XYlPVTC+Cl+j8aWviilRNj4dXH2lOHjrN3ZJXe
szDCRVgx8B+ZC5gjF46um2rEMVRiVNk/AebNOX3a7XbO313XaQUkDpGKaZyKgXZ+
n9ihW+HkM6r+uToBvliJFCU9Rri5Ela46CYnM9q2KG0qAFzJrgw+0UYF7t9yL8mI
L0BxIjpttLHE7uM0U7eS7t+nYPtMdoRCHpJSh0LPSu54UeNrqR6nZyZuJZNZRIz2
b+0s0ffGGapfFfeSuDpC4+gX97j2r9dmWnlNFwMHvj21w3Sv+89t/LOZ8aPgcNNS
ouDLBhcUihSMO8aaw630yhpipEvkhkuu/0fk+ArF+kUU/2dqrHBjGcnM0M/kBoNd
YTszE3I1MVfzKiZy2rQuR7fY81GFvxGeGgB5bjunxKq1abyV/o4/xebKqnlQPipQ
0g2a6iqXr6k4FKpDrR9Uorx4YdXidq5z/z/kDyfM++HhYlQmc0UVQ9eyd0LaqrR8
yBdbQ3bg+oLmxxq/NGDJBT6WJMn4osj1/BvsdjbLmG6CG1ZejkuucTeJpTZjqA+M
iiBM5nYcBKx48grb01bVSpBq+zw7XGRfw8/YfKoECW6N+v/6/0uJX6iHNFiw+k6q
5mpsAbx261+ivUGMGlJvJs78CiFpPnAKOsgF0cQLi/cgNE/BBTQAaeHWNWSpFfxq
Lupuy/VpnwVuo6LsFOKdca0+iOKiEwcsEClC0UEGWp6MqyVgH3cWo77xTEbW0gXq
AIyxNNGDOaWPIEXLOuwq3pX2Nu2H4AMsqyDImoaGHQ5TPQ3R9vdtqCAnc/AST4jk
TkiQvi4/QHo+Dj6u/bRLqU00R38Jqsa5IaG8BfqzfIgD/4j62gC5hfFtiSxADI17
8swv3JM+/LlUNLOz+RoSH03ABjw75Gqof85krXJkvoaRw1u/Qtdo0nvRCB68TwPO
pflUinYwWyI+r8I/eYmtLUW/7X/2LGvHFk8sH0+6hd8dWuhwbRMxfM9guaAeiNRq
la1DRr6O1vlys51gD/su+pVs/YwW8eYtMVyrFCRKVnYaGV27bnmhA6NW9qrK8W1/
cezRrI9ZSkwLxEdOwX8yYn/iwl3mg1J3/51uJ0+3023PPQFCqFiYUvSue9mW5PC4
JUQnmkUv+ehbo3pjEMWHXi/CI9Pq+BqJyUz+Y/augH5gU4SLDUCPb6CpP/8bKcxW
qXcFYgRj6dWfr/AHWYj83RB32ZQQ6WenJwYEEk32dQlSD7eLdcYSc/fKKnz5OV54
ydq6eSLIqMLMljM5iUgVZOFc3Gj34jo7Bg4bRucXiKfjaPLroBAoeP3n9VI/sZWh
1P/9/CXYHpZ28MsucHFKCOXbu3uL0op8HvG0+2nBUMItBSeiFYvbnGDj8BMnnSR3
zuCZ9UNKvkIVd0OnDJsmGUuqr0nGiauEQwCeRh62sPWSB9/ThAzXxsV4AqmBDkyT
1iBJorHIQE07VSwKqmSawfLaZ03/KEQqWy8eAFlaNALtNga/DXpGHeTXWkFD30t7
vTfR4fNw0OKjt3drC6TCOJu6prMWuOdBSF2Hre7POK1G4toUoZpbGkaNSIgxIMkV
TJ2uOTJdaiLGJceMemZrVF5TnUxkPAy94J/mmHNbumgOrxwv0rYejnH2QIXF5XeT
ucC3zJgdMoLfFesihAOfgYrg03lR/nkWqg/uJM6bj5PlNzS3ZoxFqxtfhaE/hFY8
mLLWOCpSO0RoIc5VXWHxJKUlwRJh5CyC5y2r9jX87yJID49yZGlfdMQ0vZ2c+res
TUQDr7B0mNDdAcKx6MKvz9LVAx6IU3nEpwmaJJYBJsENGokjQ+PzTYH4XwX98Nwu
+9PPKun23R6MuW1ToPqRR74RPfb1C0fve2Vvz6+yHD4wcymBwFbfTYTCZ22JuXyJ
5EoM8Y7fuzgKbtbbR/jkXn7FkjBJrDkW0utGxYGUzIEYuhVmWV+IlP4tqN0d3hTG
nJmf73nkfWP39UHr39XeUAmrvGkf/ON/kq4R6Kff8uvgqB8TWMdld93RQbdU1F3X
YusVfDbTADlUqtHa7bntiKyZ4ImPDcZvoQmmS/X/oZnV0sfZlRMsDt1zFIDFe7Qc
ZhWj/yxrfKugmsjgI9If39pvokLOTDai0vPUZ3D6KwR5SBZDSwLrInGV8kNqTzqA
z8EfH8Avv3D2mVU8CjFH5SRg4tU2Me6O4zfpc02GJUD0ix8LHQZzuYvsrtk4NkkY
kxXEXd7urucyMiFpSvNk1VhVOsD0XEZeuoIfeTvT/5/sgPvznT9zDmyh9lRfXotk
MruOLSgFNEzaWRy8Rk1zHzQ9gdFPpR6I3XWbShjzcGzzo8Psa0b28ah9xN+wS48w
1K27dvTLNYSjZSoW9I9UXxvKYKhYiIaXO6X5UttEUYAnUoYplKOrlLxp0t8la486
hHikzXIxComv2CjGBzpi9pre/OaSe1lKJTApPma0qqwDavL8MStttUWa/inrWRTB
7gCgmVIgvQK26J6QF7MCOB5K2DV8ds9yXw98hzGQagVyx1nkQ6MJY2qIXIdlfxPO
9uVYD2hcs7DfL58C6dyygA/IkLI0wc+5WbdJdIqFK/+k8VZ1m1IRVacBAhJzNyc2
i3kZi0SxixUUSQsC9c36PYtdB17ca7sgk/MRQZAFCqqOHwju/PUKgWG14cjrTmmR
Jcg2YTQdiqoUHviL4RF2yI2bufUWt+A6t7Zrqc/G1MHxRcwkqpQc3SYzZ473hISg
cPvvmQxmy4/PnMyjkj+HkNAPWigwZwbJHACA+guEnJ+2cliqn1apuz2+uSPWh+LA
DJjRvTWL6bIan1heGPqeQcnaYg0kW3bFCWcrBn21eP9cFWKkJVqAWKLfMC0xG9KW
RADvLgRllMU4rDWqY5U3GcHZk2vqJX8mIopfIb8bDqry9cA0U1ZYauU6xOIViRuM
HHAy69jrnyWknZXjCgQtlt1E3SyozXP1eLjVGD1QfCGLo6skkN843LrWDisqjYPM
q5O++g34vs6lphUAXQE4Vbs+hROX06SK0haJiuUE0BPwQrCtfZze0GM5v0wMo6Oj
ivpBL8NXNrpQMF2xn+26OZA68nOCqQiwIuuZ6yOdAGSGd2+BCh/W2rUpnkE5wtd9
WmDsvW93fYeJ+OGPD/PGQWAwP+qOwjrL0az6uBNzOKnZNdimIty4sNzdy+kzFTuN
1u4t/QtRiWhwb50DqYFQNShzxx++XtTKj5HivV1cPhX9v2ePcABtBWZFPJHbYgwl
BQoIa0kgyUiOZl/bLZBLasEP9hl2e8Nmo4k3H3i3KSrwMcZlClPl7BJBefQRMEQw
kflRuxkEtfyagiUV/DqRm90789psNpykyJ98cIj8d5aHilGzeP6gr+gT4DFnm958
wtnvb8nE/kkg4C6ddurvNNCNXXiIQsBcEec9DRshrQJ6E4sV9z6+RHID8bsfpYGU
Dv05MDGmBMbY2dDHZ4i37wraLS4JPafkpO8fM1F4OUHh0/l81a9UDUiim87d5LmC
0JivlARa0MsjucetREFBeg4MsMxRUH2VgzsYYQa/joVXBcubIf0B7KfmXHK7NtFC
BJmE2BTt689hO17qZdNEjzC6/k7U5OuG9JY3KTGmJfIh0Lm0ZveRHPuDnduvP7kn
JUMLUt9XnJ8nbRCejL2nDV+pPoNvbaHdEDvKQrpIDcT0yIMhfWujAnl4Ezqdhsxx
NnbbSwWMal5ymvcG0h2ZbLOP5CDLISr9uIlqp/mc7nLkkvUG3/QeIk+wMwmTSKoQ
l7n4u2AknF9wZrI7x/DyinP+vsZnuh7BI8JIDX4yqbApt4V2lXR5QmGFVhpjfndk
ACt0JsM34yPFvNQjp+R5oUqDHHPie1QmjyAGgL4/+8Q6G6kA1nto9XfWcbVmidyE
TEddato099bPdgspypztgYVoNAbpb9l83wrTn5ZX4z4sQoXrhEjg30L8bikeIr0U
F+2Hclq7EbN0rQwMVP9OJ3lMnKUdfj8FIqM2oRsslC1jiJvXx5L1nyIlYxbXzeUo
NevbqPXYUmB2FJuGG5H+WLjZXKhc4iBK+anv/jp3JYhsMWyf2Cr6AZnOFYKaBzYE
YARIXGEQFaC2nOepKAOLBI0J/GD+UaJHUCbEAR/biBR7nUVOm7X8lIuF00ky1qpB
R8OYsKuoWr6P9f5GA91aZm3ewK3oxNy6UErOiwX92iXGSVAsyzq9zZ/yyh8dNBFP
Lte3S9wtmEqt8CcHcDdu9R4cvr2bva07f9ziEUfwB3++qXXkL7d/td4BvSuJPv1O
bDmZoPzEuzDPSSyu/htI1eseVe0bbpKMhd5M1UvArho2CAbePRMfvjUKsgEwKlrZ
2EXGRJztUvxxRNuGradweJC1JmbMtrQ9MX88kVOhy2LUHNEuPue8dBoI8q2lLdj4
yxQxPKA4ko1LKkfrX3BHVst7wURtVZtbm6xRsadDhlPoQJ9vldBCEMQ/pG1sGXbt
MRl1h5Ve4lJWXjmtAeSVIBCBG1YM3U4Yqh5LvKo8ReMSXQKdqifwVF2Qh7TF1c0A
932igqaonEQ1car8OW1T/pi+daAIPrVKuSKah9h02gREKB4L1S7SAkviTeVHZ4qk
sXQ29pp8+RmjYlWqE1QXZu8G9ZFVGn/k6HCdpEprqdf4XWuvlIrt3yYnCRbDJH40
oqRkS5lzFl9f9Gcmjm/I48tM0cWwwTmELvKEZ1A8rsbtEEsYg3dGcRNZwenv4LqU
z21bS+P7EGeT9J+D/InFwPiqVkEsMgMXDNUxA9GJW1UM3/yC9ip3x7YmjCTSILmL
wjtJtNK0G+87KDG5IyVAezsO8R8ZmVAu1lyVfDamiofKJ7XEHPHrLs+eTZIhdDJa
qshCwWaTdFdap/OSoutLMnkDwnzdsVGP8J38FrwL1YcsXrAZEjBQ1SKmmFC0cMe2
W5wpKzL7TBifVfV/nofF0IGfYsDpfd//76rpE4h4KHVI7TNO2TMZ8cPSqw57SYWP
NsceG868qgyx0Uj4fXX0sWQwCF1WEl082e1qMlmtaKOOjeCVzO+DipbEs9dKGnRK
sXDJJmHssInFnEfrxioq/mse2uSHD2Sf5m6iIe253fT1cvGkOhCfcUPHGBVgsCjF
imfX6TqJ5Eg1254Byam9stMvTshYinaJR3Kmufjym6TzYrax8vREh6AV68pzpYCV
WKcsV8YiFBPHGj51eCSqDirlRaFNi0kZq2LAyy0pBXcYke+vlcZzISyL4PsYETQC
Yi6K9Gz1kOhk8B0QXQEhnxDzSpIUYiVYIhQukQCj5AuDdMBjGXK1rGVdqqo2lPxY
//aHuA/9sWZb3Aqqdwz7W4LmNzpjPAgzj0N+1NKhkB9Bmhuaga4fasLWBpA+dCNr
CSvYAiEb4flG8wJzn4BqJkIVHBP/GNbHOFh47IpJ8ZdBAcwPOfa6HCSn49I1xlyj
IoDVxwe7wKckil3zFfcnEyYjA7J6RcK/HqCeer7YfbE084zNvFyPOPVUT5ebYf+O
on4ytWE00Irj/zCRONNhDraSn0ZKK6UsAHUA5Pw7Ouf6ZdtFcsJ+l4HGtJWGTB+Y
OK7Szclqweae2qPRfVmhnc4qMtMlUya0f4IbDFz7M0BhCntadajXfKqur2POeAF2
hPDXxQxgXBFf6c4KM8olJoJ+oU8RK7IT/Mx6ECb9G/sEn0oaVmRuuEZOLMpD3Iyd
lyIiDZUIBs4RMpxAuz5yQqcvKqzsouuPLozfFECuLqETaLJN2Nb6miIuYZ+ROPyA
dP3vFi5WDAIzjtNVDHXQOEFN/gJkIjcf1u+kkzfXHMmR8ZbqsZDL4hiCaIAnmVKx
Pe5q/ll9/mTNQoFdo0iZWuNBclYYM0FrVctTYKRAHE7FekYSuePpPZJHcOG6NbCV
NPuOGMy/bH3EtDDwg9IeGwvZrfbtd2KgRou3FnLoOYz7bUNbiSkdUJKrBbFBG0uN
q2RJPgiaAfIdJpWz5/sfyeu0zrtalrVk4Jz2MogRCiHMdJ+AweaFlMCkSn6FHxPz
VCa88SCtVg7Au+CEJn1si4rGyBTeJbLJKqayEiAqR0Ng5fAm7ZWlRPckyRTM6SWI
YPwULggYU+VPuDBXnxLSqzPsnPWaR4hmVjTnV+kY0fMWzXoLM2sXnaF+gGBx05OZ
cfnaYsx+03RwVpeJ+61iZH1vzBw8VzAUi4nSko7iJD67UeI/kFIumr6poViidIiM
XKAcXP8CFDtxQo7M9p9tC2jv2tw/EC2/CBwYLMU1u5sTuB8BidS7B60yWprX939X
9smi0zFxfLmrh0s35vWzQ14/AIxQ/OKgkL+AXj8AAX2vSKwUhY6Uev8BxN5a71pb
dmOV/naGoAQQrB3czG4/rujl7LAWy/Gfbrg4HFUn2B3XiCAiAIB+J4A+FZ0Qve6E
xtX4SdBwGBI88tSxR0k8zqs4lUTbV/bZFRIaEbUBaKYHfmAVU2OY0mJXz9urKdgz
/fG7jrN4nVGYMN53PaGEJ9KxsTqAOXZ7xQdzZvucMwHW/WqjlHUJmLzLjmC+fuhj
XeDtjccEZijEdIrDEeCconze3Z4bRt69tUFAw+CrmaiXzj2MEVpXSOZ2sDydcHkD
jvae6pP3J6q0lThTfmrq3pWX3TE8mx5iBb/MtBBgP4TII6E7NncuN8AvwhEO4b+r
vEeVnHH+rzqB2bB5VKDwzFYj8nd9pmgewcwY7VlheKX9/gg8UVH/iinBiGIBgy10
u81s9oDHSbEsd3pF991a6yPCIwwPgy9Sts3vhRNTB2jzKkxFs6p5s8zX+3jtexTq
vayUqtU51YaR+75s2O7mIJQMoB0txw0r1u/7+FxfbdjJHsf5seAwsrSXGwo+AbrE
igrCJKllVq0k5/uVjCuSJxQgqkSZB9lcYqDV9YzNFKGuWu6j7ZPdlTkkH72zjfy9
3fs+x85oC0a7iMid/LrRDfCUudfUCgGMFBgL4L9SMo6GZfcCkzQgaRRPFcPgDMoQ
ZjrjDm9XhYPOjLC4PlIfefOxSyUwXQoxCKrftLIa4X+QaF5Xi9jZhqTBTMckSuZx
fXSiTdWLoysYr6AHqUw9XVNI8vtYnDWSsBccdWAMf+FssFFBGUcMfOemzlCuBoNd
vNMw/BGHZCKWTValvv+pWUV0PK6DGYR87Pi+EmXfnSJ5ILuyeGpQT5Fb54z9glYD
6C5kY/uBF0F8sZvFUyCLvoJxXbNoNApIkAXCeQ9MlojrCQTlrwrwYTOD8yMOMKHi
JvaPkfnUGErGa0DkuxAq152FYFdZTNbl54KfFS4myqivaJf6tG3AiMST7HhvpaWs
/hRDuHD2UAVBLX8HXV8dQi9UcMLVy+x9I14Y6F7z7cdwTaj54pZ+zxVYOmNIKsuJ
LV8LaBJc3qO56edqImFwqJtZQi9u2x3hd8+mLXSGqg1DQTLqzGZBeILXoDB7H1tV
XiELDyO69zGq+6OExgrWlup2JVHwd4lwq83vK7g2wIEPdsZq4d/vAFSaA4DQPm+U
SQIsAfNk+8dhPHEorQyUQfmb3K/YsjyIc0E2UkT3ic+28i/D7TlYkCdwGjvFqL7u
agk/8XpkNyxUjYGwejoBMwFskEyFuyX7DbBlcCE1p/ed4RE6OQMPDb6A/bEPQaBD
9m/7SH8CJc7/q/KZjSGBgBieF5+MhtMq9FMru0pCpAcDEv3yyr1DJOGVZ2MvSOtl
BDWKhEl9CuzzeXrrDioI2IObuFc4/WVKf7yeWv3I7zeMvHhZRW6P8mbtZhRLai4j
QlZIm00RkM8dyVli3uRnO8JNftQq65zKR+UFkA6BHo5HJ4pb8f8epxuD+DefPl3d
/ALXy6xbNyQs+6lG3rJw3CjKAkBcaubWqx+non1IElnhjHmhWRKoxB4GKxqVidil
pwYaNFpQr+JCjF3YKp8FmfimwtgHd8HRqfEbCHzlyVs45ilf3SGlsZuPwun7+JB/
EdX0P9WLRiIR0z3VqCtScbidf4tUIyzQ0fGqmi4xz1eYVE9P82kxurETQnGtgpdE
DrkRe6bLKqd7C+4TSy+8celAikUZN3D/q2YyPagUUZDmuga1bDY2mV8BStaHgC4Z
t/TNvdhtq/ZvOrNl8jfG+ICrpW5PxdS+JqEOoKUNSaMH+CiYlR3I/F9dRHEhdsnF
EASznQf6q6iGHWzsuggKXNWX2lkPv+wgyxmdvXzkKRFrlhq9EDP97hVmoyDLYXpk
8xYBO+jDlYXygmkWMyTBjhrE/u83dXwyRDuQxTX7WgsVOe/naUA9zwNTEKaDSJjB
/SQHyF+TI7eRDR8KxORzKrTzOqWMij26jeyUTBTCwhclPDQ4RsLXvRv/nLZ4ELSJ
li1PcUjosuH8Y482mLiaTY1LMp3TdMAqooaYOGin6UC55aOjpDXrae1KzhAzksVt
ZKFqkdPBwIqvScOZNjE6wdoFud+4VzjRzVir0fVcwmulH6l/ZBTqgwYfUfCa/aOU
bs+FxaXGPHxh+FdsFMVuxoALWe3bj0RwkfwRyvxCiQZTqJ4O3aevE/9QR0UrObRv
RaE80Rljx1yNBHr7a/6Y5FOZpQeO/xThdqjwN3iRBWONpxSzAMo/xxP5BwnqApYb
aLO9TBa4lqq5EIQ9gpXu/1c52tOP5PzFuXo3hLTzQBAHtcLdW6nOE517iH4D5jwC
AVmnW8ZS3/jDy2oESAZ8tyH+Wg6J+YdmTzU3Mhic3X+QaJg4ApOmz5ps9G2glcfE
IJ4HsqwsdGQvLUJZexi63gqjmehljaav7nC/gyotmf48te8mbRN5WueqlYp8hxES
YKonxNr3fdt+GToAfMHZEeHBLNNq669JGoPntdWicKmqw5oSKUBdsm6GcA5XEzOW
8areOgvBanDZqC9no7kwqZWkyyXgjlcvULUUSOuUAKndOuaaqY+9d/sJzkCicXxl
DOchaQAClxtB0N44kGIeLqisDUse4xbmNGPe9Z7BRMJQkwpW5TpKXcgYdS7sDDfh
2/2Y29UXnHwGs8ftYkgI2xgMP499EC5md0HPOgfyjLjpAQLr1BmJovrePNIkgy2V
dt1XGmNt0EblG+fcIbt9KwiR3MYHHl/7Xe2wkjTosD06Y3lbv/2lQ9RF7SkTVyLW
Ig0FVBgnfaQN0DKyvV9kw77IsPEGv2a0P+neBYCABGIn6QROPvMm+mcXIyeXY5wY
n8TiLV0OpvHX3/9jRVINfzr5/zg4YZEhKzaLq/JZLTPBz4Wnv3RuuAXfRPiPYoom
Cq44VOHnvudLpb2L3ASJP6HZHpWFVhp3lQn4XVJScrCMRaOXYxj+QMSYkSGOer5f
GLHpzcZcC+ggGQT2TtnGIQ0VlUgYFNf3+Qiy1irQzAEI1Fm8aoY6eOCPVQJSsKOl
NRjrxLccNjliqX3HK71cpF2JngkzVyk+1rYz42a/jXKIxGUqlYStl8xFD3EhjE0o
8lqVDtmhf8esM7RCD5UpKZrhwTWOSCkO3+dmpV42/+he3GB+QD+OsaavfM/5QLbF
1sKib4ZBCs1CRzSkaFnlo75KUA4QEJccUg8/122auGKcxZI1wSj5v8Nc8t5KBOk3
G7Edh3DhJQCvft/fM4aWFViknfpPJ/rrnhZ+yzMXaHuSUp75E+6ysKVJV0lrAWQr
hbbWE1U1zBFJKgvwKyrzVVd+eUQYsP/6J1GjNMeTF/bq+lvPZP+/U3B04Cwakl4O
fJNt2phgyE9GV9t7pIUx7vensaHtjYmpZDY4jdSESngVRUJj0l1DPy922oEuSXHa
AzTT01scsDYFLfFQxm0jVMcr16Y7hCGqHEH19Pgx9tLkphfGOhNxNvvY4cLxZ5LK
DN2iVocpK9yXwnvW5UxKIReTvUagplE3rwgjQYMnPW0UMeMz1UJ1yavPEvmIPN4B
w9+3axQOfUK6+yvQBM/NDhLTvoK5peDRDK68hBldwJ+Mjrg5HHwlwktWERM291n6
AcyxDlJEUdNM2/r0lOrth0T8yFRQzwTzGg9EoxEF0h02Xb7xc/WZaF66F5dROClM
U1evwmkwrA3Q2GZFon1tVWWxx5mxTc+Q0KJi6P9jZoR+e4leT2arPaJZtpOnKHI+
G8PIQZXOJBoSDbHNnlavrDpYwf4Z2W7XWXkMnulaVmd3iLc5e9HBOlVr5npprtGM
ntvrcAx6QtPWIzvjAd6BeFNh6UpbQw+X9kualYUT4Et1QipbnLUlZdu0Y5rSjQ4G
7tFeYt3jbJ5MQ7GmWoxmd+s9b6U5Exj0IO0Z7Kk+D+T5umh3CJSltcuTgwRpif3d
ftDUfLTooHMXorE3zGJYUXJOAQ7wncJCpiM0Y5vE5oei3v5/IfOhxSl0DoC+MquP
V3admpD3w9sBldYBMRsFO7boVNnJ+7z9H0M9d5XJcRnQ97rrO7rrhcc3+hVPMTbm
pwCR8VkLVJ9ay86COP0nQNJSBzYCtaZPzFFboCz9W/gtHLIBUl+tSbJC2N7otbiF
YbxLTj5xLMXvJ2ocJKuyGuWqB0r21meA/lfllwkvf335uWI++00awkHfOwGp2XRz
1juT1ifqEx3Ob8ATL5SgBKl1KFBsY/MZr+ka0LyKRS1kTTA0YHisPBTyCIQ7Whgm
VTHiHHE0G7UA3GegX4zDHfNq3hiotlQauqSrfbgOPii05FjrOfv8WGXRIBZaOrtO
xU+EE1xHHYX4IvJT8fOT6imw5ioUym4nq0taL5t1CiRD6rYJi/rHMLtLG+4nZrwf
GvoNwUsS9S3fHKucPuyFCU56b7XCpasDsqVyN49EpJ3WFSEiEYbZXfWlcgwZstj+
PhsaTgmrKuH8bENTsSVrKUWQC077naYP6yWptMcG1b/xDIy6s2uAKWi/1AaISbMy
194Lj2LQnLHyQ3thuo8LPv1Phc9a2A7mhkQ769P20jLY3HlNT9ruh8F7B5gND3B6
Z0XMEL7RE/iN9ICFnVOMDn1lA1Fb5mvqbtqHBWQTd34NZ6vqbdna7cTNdB94PbZ4
BflBkjoy9bD7V+JqmYKHrOIMHciqCQSvR9GH1K6Paxcp2/5f89bSNnIqJ+aIS0VL
KRv5HtNlVzJnwmny8ap6oucLMUwBZ32qF0Q3zVI5FzMFwOX9+Y+6dehZ9nLh6keK
IZQwS9DqzZ8VzX4em9VZcLDMy7kEk3anwpIekqlzHj8Syr/UhxoPkDW54a9TjQ43
H+wqIMmbkmyMSfZ64Oh6zO+/4aOY1Cs3BCrVu5H9tvTL6fxWc+MoIAk/6qZNRx5y
xsLSc1qGppy2YpRXeDkqjyyJqYNZ9AIVDzuY0kb191tSnAuMqLHe11QcnuirycFa
A/8uV2KuqdSIZZLduI4aYZGL3CHV50hC9Td+pozg2tufJakH9hf6IKl63NsjQflp
/AroqO3Q/+kJjjjqI0TreX0Qe/1ytCgqhqgVxBNVJu4cnE6TsoRHQWTems2m0VN5
jE/5AIszHL9FahAFFBoJYxPVWsFvP3yj988H/RtP7Fe+9FpKjPnhNMVHJUBdE6cy
K0WpTanSX97EYAEYQVAX+UqKYiWjBW5fXXOhaubZwgy/f9c8+Mf/K4tOoH82fWoR
JH7XtpX2qqt68ncOOCpZ/TAZdnPg47lg018IbXJJ5vtnWZuEPLBgEU5xWcKnTvzr
6ZqhCi/tfryzCV/k1TDfg4vLZQRFSHzDVOv1OisCJYzamRrEmtCkZJmeiAdsWS/o
H0bR68Qrsy+VewlrXoDYuLte0LO7nrjDV9sXurhvyU3CBKPdgp1wiFUUlLiJcwDP
R0JQ8TgKy+3O7ZlBjDrArkGolQ3UCscXgD8QWq92d7iCGLenNBDq6XW/1yClbqM9
glRik1qD/PR2H8w/62D7/9XN6xKWmefBRkpMDlcswDWDwvs4ZF7hZ4/eXrDEBgwN
YyXqBhthDm4HGlAq9VYCx5vNsWitaPdccb1FNDlYCNKvEyugcsp7cUX5AAr11f38
rgw22VzS8MzomBgoY+5Usw6ZBDZBCYCu3oO1+c0u8qfGwyRO5mys4nMSflwj1P8q
k+k7sMizqgzzrABwhdRHSQVwDIAcY4iOScMuSIsAOz01w9zf8HvgdKE/QcA9zAMJ
77aufXlHAG5hCKgTaumxMSLNv4+1diYIvzYH0J5QlX0ZA9rKZt+JHtdNcnamzEzR
2MyiY7MGUrxbWnCGJ8ZEVvY/kbcxBBFZRudWS09RuBEsxl5IStbzG10L5d+TBQj6
P/j3PteDU/V7dyB6BpKT94nVCSi591hhlF2jIMxQpoUFrqf86VfRYPj4N9aUl4MG
EZkVDZsUL6NnvLopFn7vQ4X7EOiuyoHCDVlmgwQbdkY3wfz5+QsRKobHjl/mpS+R
YD0PVpmt+rA3r+LIOucCBrHQLfBdb0a4zRvfgDHdbPpuftNnIDDsQQ+Ygd/dXASb
ORinlH9G9zZ1inAy6h5b6I5/zpwpkD4H3IVWcI2246Pq2me+AIHsqb3oljNPBe+N
fY0tL6YtmLtjeojKVMPQ+V+tN6kQ+V0/pKWUw6GOMLbKqv+kioMO00WWaRcgn4nh
KXdz253oy6DQd85IO9RVfAplvUMYn4s5bKRBePD9IS9A3UhclyuOf+3TMAVKoAcR
OF22/jFmpK4efVBh11vM4JZyX9KUqaXhiy+to1NoBMuopWQBHzz5jNcEzZZO9LWJ
kXIpZApBKxyayouGF0lHM+meY9c5lu3h/rViz1rtmNfD/sPgI4b1cEJkV+f+lWeh
G3/st9fL1U0h3zpL36uPj8uf8ns1D6FdG/Vla/3OPUefVwyzU4aboSgCog7NfYrZ
Fsc1qU5h184bcm65nK9jRwheCB5LLvBxD36rjHMKmwZgUWSUuKrWWfmDIFqrccRl
8hic76CPa4nzi0nOn5sdPK3Q22zffYrqqS5ULeDq/IAqtdKUq+APjhiWxD2uAdWy
36lFC+PbOBbMcI21WJYd8LV3KqqsNd7LVT7244YFReXVZgdp5t7tS9BNaAjHZz6h
e7wIikvJltHgcrk307nmO8wGflQxya3Iq2ojN8uLupgOwhnUb35XWX7zq79K8iKW
aJxPDW462ePIp0wXEq+svrkJA9x++FKdLGG2qJXS/3YXwhoGc6A293OMV+XN3UVe
KU8ZXBhkemYpvHPtCbMA4H29NYaEGJjRvnodGkZiwxbT2VBsrwlvmk5K8DmtCrO4
O3BHK7zIJwhQTZKeAc7LAss3KmY8aU2Q+kWPxsOj6CkA0qksw/uAejfo7z0QdMI+
xmOOVMCAijZwKlAoprcD3CDW9Xa1TnzuAesNxeTOhA+/ptPsTtAHygtyUa+ZgcWW
QTnC14DZnPQLiqsDdTXKlpT3xIe3gowZHJiHWHEjpmQjtOmrdADD+lR+M0YljK9p
AB8qTvVH9QMZJe/xAnF26QI794Gcyi6GL+cVX5Xu8mBhU5HrTfukF3BcPj2X37qI
KAOzCql//Su7FSfLpqkK5492uSgsFjIMrrPTpSzpuuN5u9dbRoCHWbuwG/P72ZRE
LeukJ9HU1MQYH1GXp/jS7McyH5QmYdqAeiKXAHNaxnbNeQK36O3jNjz2ORD0Ge2K
viDuiZjzlfYc4Pi9cTRlBXfKumz/Owm85AMbMWFmQR9EcSiE1DQYoebJJFQZvVil
sigD+1kdI4B8fZSkkdvZ0OCkKXzz2C7ebpC/qbqzGDXbjEvD+j5f3lL+9Yikrc/w
UwiOcMCYKTlurADyoEbcEtAbUsRvlpc3RQdZLxJLrg/n7uwoGv3jcBUhcO3mtG8D
dJiirYhvMyhNKJCyETu4L2RQd0biY5ipZuMQ1IoWluqB3vzYYApEA0ZdjX9zpSvU
iG5oCQ5HG/QLGJRSFwRvCUD/80H0iTSMGaZGs/Ac3IbGHkhSgKLG6BI1qtJdxzv5
6yLHL7NDt7knQnUjbpmzQQzvhQTpwIPWHbqc20lT0JOOmRqAg19MtVxDBDZzASNW
Hx+WJgeQAXMbmgEsNlX2ovMvVGBZhhWR6wulj0akhrdK/E7/6OXvEmiVNLYprmqB
2WAIu78KwSZ5fsNKmyM4KjgY2uL/IN1fR6N4LVdl/+zjbcvapnTSQUKfnema4A/s
Sj6qJDcyUG/aOJjrMOewXcV11xpVcXwUD/CPluqADie/Dp/z6Umgf1jfmO8rWiZ2
S0wBLV8dg2yLSVjvPh4ycWniWhDOeSh+N9kmdUbagx9QYV8hxTrm4XgEvSCdmqgm
hhyyi3mGmCF+gpQOAG1fXIDnA4gxdGG9eN1XGLPXGLlYtmVJJ6nUpIbhS9EtA2a/
iHu/XhFSKsa34j0OG+a2WONSVyl+0JTBFJA5/2OwsD919yGP1dhJlCCeLijS3M8X
MZGdn7Cx0sa1qpTseqY5u7OagbsLL5kfhu31/4Nh6ik4LuNsh/M3NIKgyQLKi5m1
W+EhJXTujE2/4V4sgjySw2tzHlr0FcW1enwdvS91iIT2Q2rfMaRfK1zJzhWrag4U
ov6YsNoT/kIptD/m1QPxB7XomTWEZF2FtkYTZ/wENEGOcjAoqwVF84IDmk8oHI+M
dKnhb4m6EZo//XaIbvXgb/9ecriQrSz5/qwNL6yXjJ+c4JwywQvsp/KdVvLs/Scy
Xal7OplwXrxeCz4MH94SmvMrpN1wF8i3PkXuz3ysXs5+H+5m9fb6N1fL65lWQd/e
sz1DCGs3y2vUcw77826X7M1EWGb6bdI8jv/Rc8rhn96cZJn3eSMHlz60YHOZDNkY
+fTMQX9KG2qHKLlghn1OS/rqshIoLaLgn/6u+7HY1eT3stMiR+HqULMxKrtYuo9j
C4UxkuD3mRYenoWiXR8AtK8mJJ3LFNVxnOxyC31kbDzYNQotuOuTXXldLL31V90+
UC1tErRrTgjQgVhMsuWofyQfrB1s7aqRvU1QEBoyl3SW/LkyG5U5Eqt3nziG+M7g
ZDQmpX07VirHKCsKOYFOFFvCELY1vxB1AQW0QHZgAS+e6x/2qRCiFwhRpTEf58gz
bHwA5/9KXrh8/Oq6l11vTfPeMPgQ4QWD3crGU6zA3QfhwNamQjJ2h/7+Wc/WvVGC
9XDPNZ37qIA36Gao5eB5Yr74JIJbeRQZ/gh4zvxHjVBf+uxL+nKchwwy4foZ0qhU
XIXofAeoplcZybmzUInUrbxpY5IWYagYM5Z5NLZKNHAmGR+JWmxFo7AoJnVlNjWp
DjoLQ248dTNN24xTLLMMNaRK+H+pYxO6p3fWyD3/TaZGl2j5bG0yWIALW/+m2eN6
o9wNoxNjaMfTI88lIhsVDazit4T/A/Iedlu7RHM4kj5oX7vawJ5XYa+mOW+oEypg
o8QDwYLQ4awIflSk8qNHBD99BK9vArRrdYP8r6768xEixWUptugnnyueN4Y20PJx
s9FEJRdALASXR6eK1Y2D0ujLM/LDEEAgs4uxrb+j1QIYd5/Uqwkh31ySf3QtWStO
ZJfViCFcWIBL5nFamVSaAXP3Q6JpKUjJCnurIUaiWxdnxasuCoh9joHBeirqPtCM
dLXLl97mDt86NL6IAPulW7L0ALpogWR/qpHVe3uZO7olqCk051ZrMoPWP2FXDOc9
m0/mLbAlU9IFUjTTt3yGkdDsMlxkbSR/2w4lAiHDKwqbVIX2tApcCq4ayArZ4DLq
FzMYJnMw5YbsT2jbFs0bkHzrNWgXbl9ctxvORgas9E3CBnGU6+39ujDwjsv8SUkW
01vaM/ewBLGRWVlEEgRmPSO2e18LiDPfHkt1chJqBsloPKG5i681guIQ6PIr6BVQ
IyiF5W+bJSaxMFymJ2kQscq+Bgnpe8wVTAI6FSRHfvr3utHBDTXUw5jz/fh8YBwH
vwvHheNw6xeCfufJ8B2e4EqKhnzRkV63AMQGm9lGFLv5Cal1IYF2UfxFHQAj5cDc
AE/XbLy/ZDojgSfMC6Lh9gBuDaxTJgw71ZWVsnilVauINkvD11IzvTL1pdoKbIOX
xcihhNgqkWPT/F2BC/7GoGmBn/z8xCK43z4F7o09BY6Ck8EFk2f2hLOssna9IWP6
1m2kwo3bAd83HaCCiD63pIEJhuzbt0Mly2qdk2+ELVcbs08RxHPEdryZbGCDzSrx
Cuud6eW+aeGpcpmRfn0waUXocRLTkRCY9taZ+4CL7/i/SOzKRf0MBxh53t3HPAXC
+beDYxSSRQTzOpaAs6ne420lxIT5Kg3xU/bZB0y6UULN74eApeNpNoR8z+uE0Z3d
2Qv2mTE4o41A3NXjvCZBoCou4hR9MonnoRZqPOuYh9e6MDdms3t0jIa1w/rtlWid
4DVURQQ+0x4al94LsdAKMF555puJSusOsS4abKzqVMCQF5LTzWvvbr+kh1+FC+eC
yuwqUDJhPgSFV2ldNW5vo27gxvT0qNn9KZNpjMBOsFrn/q767T3YLFkOd2x3mg+Q
biCsi6ycbsUiY3i+j0Gna03DjBf4zAiojnf+zuzDrlzTU94k2bpnmkBjM+9y4zNV
LK0ZtfGWvNzGauHQ9HMGWlUP5/hC8OW1yz/LAs58YbxcBvOs0IeqvPW0QVpgSHKs
QeB260nZxBsXgbDpy/oZM6TNmE76RwIRUYwbYAseofK0GfEAI8M2jvjYsLIsa9oa
f7ImDLe2do614XStAYisk2QtV1eTV4R7KDrLmuhhSRXYE0yQ2rSIfMoTsnQ5fsPU
Djyjtj4nVBFuqy8EHIw9Js9r9o60QVg++qmmLWjc70kYSqDRyA0Q1Cf0aB9S8IPT
iy6JpeX2m38kF2eELRfNw+S1bGEnjjOP+1Ntq3iFGbQ+QREidrw74gnaIHsg7qMO
HjXGuUcDsheBse7ch0asYZgKQpZ3Txe8lv3wXFJECCytAV4SHXfgHR1hxxDcw3+u
vz554H9oZT/Tt8+tK6TBScvPAcNSmBQl2ppqvTwJMRztblEqaqzDPBjR7f4tAiqp
ABbWLeqFLwq9n/R/xt7PnjmbbuHx3IECIzvTDk4NR7CxpwHWH7u0v+6uO1d9bOQ9
lfMxpFHSOxqHDbps1YCx0iXpXuevGPQc6/hC5FU/P169rvvkD2kN0GYPG9zxy2qw
s6ssyfYEqad7EAOsIX7/Vild41JC0wni1ieGkr69irijhtHMeO2SjaKUKeNRmspE
XlPOBMYpcyRg571+qeKmQRD03V74Xn4IZy4jvby5CxKs6L6MqZRz7yUThIn0ETA+
K4EGrq3+p+c3bKGibQRVbMUSX8jooacdxHLy6Xghw3751sdhUP4ZjG4dobz8uXjz
E2C6bOsM+LwbxFHQte2rnmGdcAjHYw4/+CS8RnIOIl+pW/exRolMumXUDbSzo3Xp
ahxmFww1s7KtIo5siQSkr3dh4J/Xi51t5YKh8t6OevYwgeHBRkXFv6yRK6NFGPVE
mmYpSNHQnhfUdAbUogZQvHKKFMO5NmFp0A1GfQktKmgi4zCZX2vkhGFVz5Sd41yb
O2c6wMQZHktG1cIAm/p3LWYRUWCStCdFqA/TPO/bsXOXKVQUuU05bWyYgkhAse64
pQake4N95wXeWSqqEnaGyXkm5P6yZIzzpy5d2CNCpsy4cC3ta8Iktg325PeCyRs0
owRomZAFwIHYN43DYENEgOI3Q51K65VrpKQ+O294dugLp+KyevZin9jk4mUo/noR
YK483ycsLeBzkt7i6Jy56+tXUJG/siGGJtz/kzBEefI63dU2/4ztyi0peUDZXbUa
wZ4A+8NSzobTWsr5goKDuO1J45TE6/gVfBs060eQNudCrFaX+MF/d2sr4KMIIpKE
7c5ivRffIU5LMVFnSKN9jvkS7lnD1xJp1IraBu+0a+AWRmHJIVr/RwwE+50Cl/qY
/JqXPtpMwRrRPFyE3MVyCnL7v9BGNG4Xkol87azDzHZ9nPa6EIncikUVNT/jiSRH
wx0qX6K+ux3idcytBsrlGHYhLClY3X1t1nDooOAwQmatL8cKQoRGSZXcRgAe9Ep+
kOt+73B5Hlu8I3kpwbg7ZOePRduAkEwhg/RSKGvVVCWlRMC4o9QuZraKNCavuPvc
LuuP5GFrsDJNnKTW2/O1KzfZElvAjMui054QoJgtK48cbEmoUboptn0avodSE4/q
ADtJ4QRxzx502Ozsm+aer3gD1V/fqmdnmqCp4ppoitgu/HoSHNm94JVhUsWcYEih
JwAoa4ijdJBHOz2WJwvSASObDeA2ZrgJhNV2XJbMXv9xPecZUj1hKgYOgnoQxaBu
C753l5aPVq7aigDYa/Rz3r70M/t2xeJzqOQ9L+tOsHs0bDm+kkeaVAppJp3i4V2B
DcWXrSyvYJWIbfBgKiO1hKa4Rt3LRaco9MvbDwoNqXsiKl7Ery+TkzfF+uBwN+Je
7s/KdkSXJqz7WKBC/axhnO59+oLWmp8uMe9DMnWZL1UiB0zZiWkvBQ0q5MdSXjiL
1K+fNtT+0b6M9DbGbRIjUDioHPs+4HIscbNzV9/UwqyG8HyqzGA/NjoCaV4cf2J9
wFeo6gAZAbDqAHl3Cm/qUTG/omG1Ac4oObmCw6zkf/WT+ubIMqOlkoUbT+lZOUyt
EjKsUoAh3+aijb2qlfRJHMmE+wLe3BuPaIn/dosbxlTg4G7RgX7YtUpxIKoGRwz6
apX0kFDQbU9dVx2EAbj93h9hE3lKOcmcXgh5rCWoKsFJaJkQboF1YwIXA2TKr90T
4joH+2Ed3P4LpqCVPs+hXNeUwXiWsYpzXNgNMvbfXzoNGx49kdqIvrh7f+gqz/Ve
sWnvVNt4N/wPZGqU28EnGgngitTzzUbac3Wk4GxK209ON5I+aIfO84UwSc1mri1a
UR/mwXbd3cUTW627lKiojPuSVXE68U5su8Daj3EibtULzR/scy2m2RWhWwZCtgHG
tzwOzwlpvYKUbovx9EI2DKiVtTJDJQs4lTeSAM9wV0nlOY1e41Tn8MUZtS1Lebqb
8G62pQt1n6ZhW4TXJrqYmIbdLbS1NKFyXnXeavaZQOjBL1O23Tg7lwTDcztfULPe
iOYe+AI76w788p3fJBQ6nlho778fQnKkRxgg7HXpFGMkeT3rxCx0kkqwi3vNLYHa
YJyM8MmxMq/u/gKN7bAmNjd+yz76pWdmu0wiNqfXCx9ykaDWAIjaoAnNI8RHELgk
bsW3i2/6Aa7OoYJ5cbhAc2j34ahcV37WSpTFx5jWqHZBC1d56lsUPliN6iNtcxeC
fk23RW9H0FStiMyF5mX7R4Ic0W4R5bkE+iGV8fw80jQDBia8pwVJtFum4L0RDHhc
e7apMGvtx9tljFlOKwu4uF6k3+yleRfmzwCufG0AGUjnosqdzSYtQ3+5PhcEK4JU
0vMMWnyAAGK5WdG65c4pkYhqQY5PMcZj+c6+5nhZWslnpTO3JeJNRFsRT3BycB6B
3oUh8VHbSQToJcCKRhs070Iv65C6kDLiZpqfWi+3PLbpEa8hK7HNkSKMQoxU0O7y
1cnU2AlvpxACJ05MYXzhRHqVkvtX4NmCjSmHIgXSf++c/nC//uAB+cxoqEAcj4bP
azEOy3n9fjLLvhhlTHGh5IhHBs1fXz7ZhRBiBdBNVbRjznGDwv7ysUppN1vgHuS7
IdajHXdF1F9wr4tgK50DAq+9oZPQJV1ZW9eZVfQAd+tDzPrUFcdcL+4KPU0N4g6t
U61qjNdghfWSWJEmWf2DDxTtmJrW8j5v0f4KIdxDeWFuwlHLDH3CAMBrc0UMfDAR
O5VAAw3YNqJenUeqnLhk1Es7o2Wz4hVcispvEUnhiZ5luhqfb7hg+SGY5Ac/Dtcg
XjtNUYGPTAI2/tZP/n9A7QVIBExynFkajzl+p4+T8qMQEwA5P/HkD21Qfik6Qfhu
S4lZNglCPXjq/+BS3DRAOrXCGYSlOVa3+1jZwU3ClPdkT48vbyNLHdl+a8AroCxc
8KT0HcASJUW7/NzblP9pdmFmO2oU/5PhBWqkrQN/BFR/Zgmn17A81nJ95Dq/rCCX
rCX8xF2kr0NNyMK0bsYeccsg4hHJwupBuYALcC+DB5xHBdshX307tArPrMnWvwTS
kVN1BuTvi1/EaxtMi+RDqQ9xq1KLDmMPRCVQocDTXbZlxTT1z3m6Jv418KW8qFaf
51vmFtxucknWcwTXzRYAfjrX3IgL0kBpQHpnLRv6SE0K+KnQGvhtslkQUCt+Nl6Y
K0XmlOtTyZGPZfcTGUfjVuWecUdHTadBFmUi85Rq7jE25BYpyFjLJIpCvOjGGh+e
KwAENf63g5il4/yWMvMAhjvULajtbaZgccOeHoVyYM7xYjN5CwZXcF9B8tX5s42l
+2gyqmUHRi3XdtBUIM/Ulpv33m/lPi22hvPONp2lwQ4b0XrdWu+7m5ViUlBgy8zE
ExKSHJK4KKox7CceMh/qNM2LJoVdpcMRaQ3TZfqSUwTkYunEi8ke8sUVkmDtWuHB
ii9UrSnsbsSamUNy/8gQzQswxjT7LW6XpKsdWgFanmRhOp6ABwFYagsWlMRGaqPT
OaDhI8kaeXA716fbCHgmMb/wtyt9DkC4PubH5hyESanZ9ooevNebuBaDD8mnm35j
J+Vq4GS90v0Iol2th841SD3HGgyc7HUu4rIDvoD8Pn7/y7AojHyRwt2qCrUfb45c
bxodQmQp3znkT2aIDoGFRM8YchQhW4GW3Yfc5GrRHJBcwdsxIl69J7/l/mq+0hsM
Xy7Q055ivJDmn0vKQjsX8oZbdMPAwR/G54J6RE/EPScJt5NwlNBMOYXm7sKb7XpH
hm2kuZPMgW4Hn64RbzSq154RaN8FmK6pWPaTrOD7hkGgQJbUirD/KAOcZdV+SeSS
XMu4Od54HedV9qiPZ+WXBGaH5s41LUvXeUH0aZOdByss744G9bdePActMR+dRqRV
XLaoghQaOVKQnD2/1EQwxnXfDEJaDq9TL7TdqF6ngIVLzatxvgIM4HqR01+mcHMx
sDjD7iCZMgrMyWhY/dZid77uG0tan+Okg+NBSyRkgGZD5/t/8b3PnmC79B3xthDm
Qd25El9yXMcItZshQFpBZTSLQVYxgHqFt/mhMGHirXPtbPiKOr6uwJ99QEiyxNhS
pkdOk697HsCi1uCBiO45Wywp4aK97yNvTrwLHvOmYwjC7a0p4uUKURpdXLkfDE/X
Qb1KCGRdhB/IU194c6ehysOvfy+dnAVeWsH92+8Yg4fnlr3WysQsVZ/O5rtjMSvM
PR3q5pgP1GbbLyWEmuXc0hTtrNL98LiYFDaBmp7mKH7ZfWRb59WaouoJtACDPnBm
MipCtzNQ1wXB9otTB/MMtDrXvK1LPXMs0HUtvSRE6A7x4wh6128N9N5Se+55hx0L
HWmiIZkv+5GeaiklQACXujJNxZoMF8cG4/MoW78ih5DUZy/yxo2xAIx9v70jSmMG
xpJ47Nq3bEgyT3o9iRxaHN+WXBpkNBNO4ly1svqbOXyLZPMzcSzmoCWBr6EZopco
cywL9l10nbzYSZZ6V0SJOfMhX5UPxG56+n0we7G51hyFT6raXNEqvphYkuIlGtF4
miWZIrZyhvBW22pNAYbj6ouN389s6b2dp+NZQihJY7K0PQTl1+TpNHnWU/j9O3Rw
WjxndU767AhRnwT/WPIL821NmgddeYZnDuYV7CuRoxtaN+b3HWgN1LYI4LCKbp8D
A9vjKyy20kedt/4ged9qLyNhtjYtN8iAPtU5723iwSfAcZBeas5uxSq3+gkVgXcm
AkkuH2Re8nwUjtJVdR5pe8a0UmAbhxJAOSMzFKsTiZyoYJsQrgdK9+W0sMNCzFfK
ql7ZjqD10WXfZgMWUBm72wkxX8jUod1n77+pQ6wSmhvumeQjIu0ZWUtmSQgGdUOO
BEcfiV0YWSorAteRfKO9T0gcA6NkC2SjVT2lUSw4FkvPo7i5/h9ItUWP4yNWRFBf
CFs9SaE6Jc1rsk6Jj2zlhvWe4HrlG/yTV6b4SWlCyFxuPtlTkYaqRSjsACH0cU5d
mob/E5437zaNgrU4fvDm04b+whmXUEM961OmzaeOEpPfllKU8SN0dvHMQpdvRN0E
vCjAfLZshvDOo+JwAfuW5tDWMn4LVICwriDmPgrn6TD0/+x4ywJPJMF4zQNN00r0
3rI4ZCo4wK1I+RWQGWVV59WlohID0yIrIgvUAVmdU1DUkFAQxHb1BsydTG6tHWb4
VLTXgR9b6PVW+Jq8uuEZ4v1xk+yaIN4r84FprLryVfIkCiTk3VNExrgKk8WQag5k
mXBCkixd8bNVg4DBh8KdZptgOMrz+hvWb6ClyIGR/9RdJZV3NjtzG86qlhAKxnbZ
PwsMCsmjNwxx7nG3A2B9BLpupxDdzWTDLctELhn7XuBFoFckXk4V/KAf1MBomYZ+
CteKpJPOrhEx+yzHp2daIikRLmIEt080AMdK/qPuLDKuO5Scu5qACi4WQ7MfFH9K
7xEeFA20GS3I0qiurYj3zM8/c9BG0i9gJbdEow+UQjZT6EUUlv1slhZ/lCQlUytv
/tcx7jcwV3XGx86xA/NPpfOmOELVvXui1619CA6NjI+gsyExnOrpFbTfRdG+Ghkc
wddwFvQ1+sgwt7WMNuyyhCMbSJmlDoC8oI1TW8M91opo7d+4jBX+pKz+ama7lhMY
CFx9lAHuif6GQsENFsTkJMzJKljRW/UosZrbH38oaM81H3fMD7Fe8xTjlElmiBSR
pizcctJYFtpHExM1Gi2YEyqX5xhXDFFgOTHUC4OIRjoxYA2k7svJkvKkAPIkYN39
9EGlbGSpdx+j9HnG0Lnvxs6YHnUwW/8WOckHngLndzZJ68cjVJTQhnigQHfvccX1
ZjvSW4LgZ/Wwm2Jd3kNHy8+7gT9HIsVRP2T67xyCxoINQwdPFfD7A4gPnN7RbG3S
J4/Kk8MLcwPST0GGi4KuPA2w7khHqCfGx4kYH7s9hVZr5yEGiFOFPfTtCWWmqMh8
jaI7zJTdj+R7jOrd8cdUkhIO7W97beEh7wlUGvrJO06zqdKWV62+s7ltFQ6C5ur7
IcmtHy1QhMN4qQPDHGzXhCHDG7zo8hoaJBlDZwpHIlI4fynhsBfgEzmE30GZy6Di
/upPXtSoAfyh16z8Po7kSR52ncYJpAPVyPv4DRsWaGWQ/UrJlgjiponXyKKaLe2u
F3xXED9a3dXsrqvBhZ80TKvSrg39kDU/u3mgorEAjpPtSAQkvDd80asYHozeqQal
K4Z7zFGBgqz61qPoyugoT17g6hFzRHsVezDAWwocUig6Lr8i0sGh/a9UWEVZ8V+R
Hf+Zam5nh/CmwpPwIb/dn4nIPjH/+1lud+dGcWkLgeCEyJV4gQF0sFEwKKr2+/vR
3uScYLdGLcN0Btw21xPgr7T5lsKeymjUgmSNEhjM11YhY2eDDzxBoLXdonDTg4Fn
8AGiesSABWzgQDFAYz3mjAhY1XMsMxKjfRSiDu0STJUVE+MFSPxBvjYlHJzV7weO
RHRYFi/KFu7TxNUrM4zzjl4qHkqgPvD/nNQ9Ke0UyYjgCCIwnJ6BBN2mOGKGBKhJ
GJV8dbD+02cshXv3YsR1HALrCxGXwmCTyQ77bLUtz9E2UMXzIJmBtNHKfXVtnsos
qv834gk4TpfhbcjxLzj3niLjRzxpRCnPwZyeU1OiIewnDpvIA1qtgb0rUzjbhs5B
SnzrMCwHQ3yYNBr9Uo9cbLJD7LYQAK6KXB1UMC9k8h5ypDIeEOuZO0TYf8nkAzo3
USsJFul3uWUS/KlYYPuU0CETBUZ9EnCSdUL2hq3tjgL/AiDxJVJrPnbsUbXwVqeO
vgUFonksoIE+yx/3NoK+G/1q+FysUzpmarkEfIaCx9tuKsmnjHQt83qoP8t0yYpR
Lmyj2Q6QGn3+eNbEhXm8XskPf+C5334/3QM4lDtqJOHt6MuVaULWL02ocXpoJtGf
WNcy12I1IdewwEX5TRsZ2+8g37e8+qxlqtGNZE2Ou7lmXDbNI+7Nw0cQLpBjvPcE
Zb8yXSI0UmDY57V+xhHfZpOQjrRfkr3All0fYPZupNkxCWp1ftYS6On+U0Yzju9Q
Wl71nsVzhzqe4v956V3JPFq8IGSp8FHsEFQUvEhRqqR2ROlv42s3Q9jCREsI6g6g
NkhjrwzOy2VXMCU5ItqxSqkYt2gLGnNp90DCrDWdI/3Nom/5Rx6ItqdbtPoRIHKQ
bqenc5Rc2SNnCQaYW0wok89pvuEROK+99eM5tF6+LbeE0FORNMLLJHMK9wS1xk2E
M6N7OqyxaZnbz3VDP7UIQv+z2rzXz5xVEJCAPKYR2X3ZZ6e9ac+DA57lx1qozRtM
WfVfFEUCdsPceTIwS+h2fiLSJpqQqNtKWNwIBv+tThVuPSOWMNw+43RIy/9WXd/y
/VoUjWKfquJiDgB6vK663NRdkX3WEIAkAv0l/PiG3NE9sndhZX1E/lyLNzlhKuRs
xdTL8mdsPvBMzlVw1h+KiyQDFxaEcAxJ/SptPjAZ3gbkhkQwwvgIYHOigXXPSHCk
Ap4bNHT606DQtAWKJk65D1YEB1wc7tHSIv5xZ2gQLiXY6XN8zoCMAxFqHCKO6ETF
NFTjzpf5nwtGJ9Mar3YSj1+mI/ersmd5iqms5Dfq/W1mzUu/fFSyE3aDA1lx5Ctk
bzbihTX13ADZX2mzUUx7O/jo2i+gWVMZTihHhuTbr5J8fyQT9H47EOJoL+2Rq3YI
F9Came0CwA2kSyorDNFQ0fJ8ISNbNiI9nHBL0Dr/wVGyh5ZJu5rz5SAsJo7iDjDW
FIDLzyKpTxuGIKm9rtPkrdqG8VEgnJwGYWa3m++DGzbRE5ncIoIUmnxovITl5Fy+
6M7ZniJPiBln8Z+ihQL93z5FGrCtPjZBaS7Oxr0wnBGgKNMWONgJekipHuQu1ChB
iSl5ICSTesf2/O6m4Ps9/Q3Muz692M+zZbXyr0SUsFCghpo1Knk8EKjHEgtfRTWm
gHTwCGlJeZyq4jAWOaYRYbxDhls/qjRGRhYuHzmvtlspkxkLLN6D9hJdTpFNBnd4
SXL9JbUDKWgqhzjF+KBp3oWvLTgsw8TwmMys5LzBPEvpyrIB8yM3HIHzf92/VVj7
wa0dFQRT4dpVMCzPjkVX/K9HamkRxjSASwoYTueGSrV6bdBOBRf4hMwZrpfg3B1n
Cvjf+yFiazB1WFfqfPyuOT+RY+xGYgILv9DumQjUb6mDQNyjbrdOr0SjfFEAkUe2
bCrDrT8htYuqvn4yn5964w+Yz/5J4LEeMqbEPX+4s88iqy1SGMosuFhF9IFnJBvk
v4x1bjd2+GYJwP3ZhlTanOyDiNHcnsxJp7FP1InwlA8yLlkSZU5l7/Jz41hWr7vH
m38rUVvfdm8LKjkzsjNloU2sYCFKngy9Z8gTLVaOAlfnw1zR6uLX8J+vk83RZ5N5
vvUZJVh2JBH2ElL2jb0uDS1LKnW9GbPg2op/4Qv4xzAOY5pqbP9l9ml1VN1AQwjU
dk4Pz2/VZTs479xz1dY1e5d3j2VDD72HqL+9/eBXD+FKPMpsY+qmDB2P4PJ42pUx
4r5rBx0bBoE/mU3TJkMacls5Z6ru2rJChDs5pg+lm2WH7TVrKQqftNR6QNkBDmT0
vrGRSoz6qaXohFC+FiHpWRucLX6REygWWmKTcYpA0qtFsW/X2zYudsQLUzcRXZeV
it0HX751vpF4vJMy5u3ZZAe3Cmm14Q5NZ/8UACh5cRJJWLM3yUEh50LDOoq0GZAp
+ubiNg0oI/bzmjELPf32KeD+YzV9wLsvgYiHn1VE320yK5jegxVR4m1muLJtcp07
C/CM8MdAq5eGzkEM0XFcTKUMYgCnQF4vlcuN3o2bISe9sA2H9Paotv1BYOntk2iq
KQDkERwkFwY9oibH1S3zq9iK60zUS3pLiH4A6nkcES61z9219QVu4OL+/6o90V+M
oypuFPjIJ9fjDyTG9uwNJpMxv+vByQsXQPJimOtYOawo5ujWZMBdMSsN+YNLINte
mb5ykIlnB+ongRwXvGfNQ5rJ9ZzeHDanZnGqm+s1F2HbT6sIo/xUll1YL9gFAlAL
6yM0C1/5Scmy2kWxo2rNmXk99vGHBNmhsbA7BZ4oHI7S3WD61YaWcBQMzIcUBWnU
Jm187MdZTiacDN5vxd3vzMkYDTrB328a4UxvG8jGHFejJpPdtEh811qMLSTOshf/
MZ3rQJQTue/2y2IhkDFi/IrTd23FV/rM0jguxb6TuO0Md5/GbWEVU1TtMgA4SFb3
xxtABnwUDNK+39wHCXl0+yzk2gKCA63Jab8ur7DYGl/Au+5W46Wq6hKX9X73/YRR
0L63dWeL2jxaKr9v3mFnPfM1xK/Mhaj3M6QhnaiwmvDAGriJHf4WerfafB8tEIT6
T46cSYqFx5UT1MmUPnJDS6bqtJkCZEccuD0+GBvXfKXSNguAK/IrYjN9wtZ3H1lL
3/uBn4q7n00W2uCdfQ6F+2Qg4HyNU0y397v732wLvhuV+aAhmZVMmRT6jh+YmwYi
mDDj/VcLVNWqWTxL6nnMuEZZBqVd9bt3KEcFrgXlFAS+1ESYcpdQ/I0mswNtMIhf
lh+7ewbmq5PZRvjuaDx9wjEQcuvkCuxG01eTXtrXUHLFpa6vx207zglLVYqtOqoA
w2c3/aeARgXa4pelLHGN6o5qumc3Kc534u36hFl1KYPlobbn/F9X4DxOIAA8Gbkp
/KBqxsy2H7FzYYMLaDl+DM8yg8xu4+Yds1MOAedeseWBRf8zsMQPXiHYKIqIOAAe
CK4WyI82tYM77sFySw3SRdf2ajPW8/AbTfZ7IUDUIWcOTQxMeSqsJ2uxJDL+kc4h
`pragma protect end_protected
