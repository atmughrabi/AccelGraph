// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
baKBjEor1rDi7yFcHZsF9Q4r638oKQV3SDiUu4aB/tI9mjpYDNJlCOZfx2PDp3iI
EI7G7IOJD+tzRoDAqSpaaBBQE4JMo3rU2/upCDMo/aEk/VXJfnZvskxyJjzGiYxR
vWwDPPH2mahXVSlYg2doUpwB3mnXjImvXf1m3ldBHHg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27296)
UOJyLLxKbVPtmre5TIVrflGF3sOtgL5mWoVUPgcDEqr31bRio20BeNB3MDe8EIyp
rbAXJvNDi3rk3wMsKJYwAbSyU4lh22LzH27zlGW9JVJJlW7wEwW4Hq1gnOfZLpFA
wpFTPEDHnQntkml3eyMC5EMKBCr8HiW6uh7jW5DlHqj5ply6uKVnyg44ZSp/dZBR
Gj7oOiFlWpG5QdFr3Wr05WUcupNYCIvsjsZ5x8AEzY9TlR4HYH7cE7QlcDxx2AJ7
c1r5OZBZYVWoW1Qb4yIrkXGMoWYxVMB/yplw8Yq/ChZzmbHdSyvm5xZx5DoZXTOM
2prnDIs6Sbmb253E5uzxaKN88uOr8m3iK2Tzgd2xJiQxYg/ugeewsej8HYvLws8B
UvShYnl+SGHWIcZAUAKAriu/vq8OOh/wRJ5OTVFG8bLip4m0GwZz2nNGpnUWa9KS
gfZE/WgYODSlrBB2Ncqg5NLRA2GZi1PObk3192YYbHdLwkJlBaGPnmz3VRZClQfA
9vFhLFdTpyJjI1UFs++0HseJf+2z2jkYfF0WkFDUq8yB5rGpDVsyvuYRuWXpX134
w2uTvf4iVpnPLX6B7JYktHCsCDd7o2M+mNYhxklC0+H+gU9NAj2wWxI4y2oa+QiR
ihxkHm7n8bncPDqyAMH55C4cXlomr4axA18Lw1rerFIw2gMw3xxKYbSemHOR03mN
xa2Ig++B0DHgpUob7U7YHeiMWaMQQoFMYv3AplDFA7k0vB/1Z5rjyyi/oRgjupP3
PpB9VVll7mU4yZSOPdHPXw0eKVTgVrKeUSkZ3Ecxp1N79TNBU31HPwAkJ8NHE2nJ
ahTBAJy/i+oUckfDNdA/+JlN0YVANWFWgi3foNaCUnROgHN0TOog8B83Pw4GmijI
wIGVjQ2f3LFt/Ud0Z8PohylPoe2xelizfQumHTVHLZ4oaRO0VgHYu/7oIN1Grwpd
kIVnPrAv4TYlOMFvaHAY64oMFiirQuoCWHjwIMif/qgwY17RUvze0nppPKGF+FF8
9nYnRS5cV42I0qwtkBPGqrLQj4vWmTEs9m3X6SpmFRmwUntp29UnPlfajm09zVnP
2LNSfhlNGV5yiRAPrS+sdBTUFQP/YKwF4VHQpuZDNfnaHnFEQd7FJd9mOUyWzgzx
77BHASAMY8jqgbp8GbTs2hM04rIZGbkPecEo7CUAg5hYpI3VP/2Vk8cq6dKEoBfa
8d863kwItYw0MCzwf0JGQMUHojhugQdqQlmNKcHUlv9aaAaMmyq802OmxpdPmjQj
wMm8fTu/KW7zA9shcpeQB5PshMiAi9aYSXVqpNwgX8sG2xtfSjLusi6wCt4V1jVz
6Q/by69KIJyDuhbevbg9e88IRKL8rk2ekbu8nulpy8W22bqfwDGKz/w3Al8hNJ3M
N4YTYiPjxDNT+sfFmIwMpkFdmo2MdXYyMukU4txT4v6NTxLuekGGjVTEMWHSR96G
ToPGTL+RA4vfNlFy68WIEp8HXGJjceC9WCzaH6IBhcwEqu6Dq0kJW5PeyJse7L8M
9kDzXxXDKHoxDKPJRuO0fYhIGNezbxDF6TwdWwd7xW/mWBOjHVJBySl4uPJMYYxR
bY+c4s2LSwyvW7uGNnhIYJETy58ZzXfWWGl35TZJX0qx61ZcvGhJfUCKxRJS49Q/
MDyKRkepHgvbjunWFf1BLTKwKblZXnz4AZ7ewNnq03ccphwUdwbGS/ZnDzIwv4dC
Tb/A34pm1ofxLMeMzAYKPGB0xgZH/NxtUUOoet+54X4yL45TU1/wjd/o4+3w9ff8
W3cypueuFfFqpN50FpfhL8iF47j6h0k+GeJqkH/rcop1RRD/nLwVA4vWpZ31tuhK
9AC6h+oSmbI1VNz7qYjZgssG5ZpiBNgV/lwQepXpqKu3TkabzCp3IjAP6onsUYEe
TNyM8Y6IzciYPLgWirXugzrhfTZQYUkgy4ne9uF3QIsh8iTiXtAGjUXAoqlHanVa
eFV2tWcl8FzllgY9bX5l1v7omPLtgOc3TAKB+ZC80TJH5TGJpW60Uo4RdXoZRaNJ
hnJtcXO/peWRqi0w5meovsZ0ItieieHM0zSk4bEGxsTvXbnK2YMK7wo2uAdUbhKX
4Ae7C4VSJ/F5WwXrcrcQBfhg4k0E72GoDSFz/9jNsLiKJ57zV7Kz6ZMxZlQ9zpkI
yxlycCJmnsVy80+OFk44F5fIQEDuqO3nNRw0CjZZKunYFd6IjOA8YhyHAbiDJeZy
FIh1PtOUuP2FDYyJLmUUuI9avqUM9B8LmXFxs8XhSkrQfaoPD0NHFNA7vEFtlH0n
u7B1pi30GUV0C1HqfB/4XaUW89nlHTEM9PhIPlQfTt9fmUCZ9GenhQB4lthXX1cM
dvy3X6h6O7SYZeE4n9Uto3vPXeJX//493a2COtXtCZcTQ3evF6jwtqaeo646vsSs
J8FTAYHF7EFmukIsLDtrS39MfIWidSvrbAVB16umkpe5zJG1hKXiaK+W0NtL4MeB
cGFmEzUtsn4ZIK1sdsRRPufgxuGgsu8ZF1uME2quQ2mYZx4Us7WBhI3LTRbuK7Fl
Wr4uwDAVJotOV7KU0ih+HZdws8YNtVTNwNwKsqP8hx05moK4M1bCaupWgoaSLMwU
92YhnLHTqujHkQE+Tjd9fDHMor0IvZU+Dpmqj7s1HioZhLAkVz076nyg/2Fy0gOd
+/hD+gx3bD9HHxA23Hnk0a+lTB1c77ec5YMFNsS992/wDci383GLaEZGz8VZ/Qoh
U1jzAJeokzBq63z8+6UTaltOB2K2dTELcoZ3CRJ9fOpJ/5CP9mUsbp8RsffpsDDJ
DNLP6Tyw/onk08pC0PYx2Nw/WeQWrIINR5hNPx06BVA8AHtpvoeBHGxA13k8N/1P
4wmwlmCbuaJ0erTBwUhfHPHJT7ErWa2dVIRaaabJcu+dPKdBT+hUVeK5Usi0Pw/s
hF2Mpj+EAa3FxwKO2LX8SCGS5BVf2gqvrWGmc9lItJmbyJI8kKx8EZXNNOX+QkY/
Cs8aOYmegdu4EIKpaU5LqN9MRBS9EQnn0l7KuSarIK5ZJzAgRQ13FMZcdzCuX3de
bK0GwFEGj1xRgItvT5J8KkRhz31bJCQix6bMpHEYYvAx7Ov3ClLJUWczwKDlPNvR
toSkkfDVrUmXUVgKDCH2AGRWh8R15pRzDW9NbbK8SIceOTOSqfpl+oW6Gilud7fa
P5m8fOl713gDjSPOHi6tB6FzIXX2DqJU95llbgY960kfzITc3zIwgNTTU+rrzwVt
P9jxZUTzzX9ua0FwFm0HlPiDaz/eFozHcB1Vh4NYhAFur3EROqho57+2VaEuxuTc
nrPt9uC1Du6MPUnXpAmNnL6haumDt2f1DWIuJy2v0QRjmyM3Wy82Hc8Pdvl00OoU
ANpJKaR/PeCtaX4PbL1jYYLIfTpL+ebThmpdiYN9UAVGU61gn6oyjK66gq8DNZFa
bZNBjv6Ab6YpkkV5g/ezeF8KOW+kEyLJx/y/HygCq0U0XFpfj5HC51++3E9F8Ssk
qTny+g+O3lMMF0WQbzqwQOQblg2JWw+owrOdJYaaUXYqITgodnHV+XDTfpDYdZ+/
gZzgWiNAn4SxA2mVR+oTTsJVFfqrvxuEwCvZSkgoA3Xchq+bmoLiC6hct5xzXSgZ
LbVYQlmqvfZICH0eeFwyLf+lUP22dUvBIWmCfBZWHlMekDk0Ye1v2PIMXV57Aas9
mWxL/tyyLXaMYBcCXFXUIliBaCMHtVKb76BuVtm4zMqBqAtfjzZmFN4DYjUbd3+T
EN+ZKf749qCYVQPiQ80rPgtfnRhcC/iQWWuQs21phpuwZ4im5mmK16mbcVY8auxL
PuFQG904YTn+n1j+eskNXT6qyPyvPsYCuAE9D66o424wcf4Gq100okIxR+9N2OCB
dbrZaQFPfJyMvOU7vyBIgBNFMmA3BikEeuOVGUdoIiKx+qz7LN+vkuhhZoaZ386u
LaeW5d67bKnbuMZ4/EBZUmNIlJUcyl568fWh+G2yBD23lM8EogKFWc4RYI6OSX/n
F7NX2W8ZWqB8C1sbqF95CNETioJJ61obDfcdXdQJTZUEEfKtDZXdHTQwOYcfowQx
UkpsCV55TgG7LBigOU8IJCaqCH7cU8wJJtzyx9QPMLgsRMQuX7wZK8pyorB1vS7O
01Ir/RO4ZMYsFVeMI9ES7r2e8li/+Z8//EfCP8+AvIvyPkVLSBVpFdSDFqZFKpXY
IUPqHWbC/osSyteNcUzes3au3i9JnnutExg6cnFnaG2hBenekegZ5J2ApOzIICz6
RsFS+LZRgGRzhxOPs5I09bXnVJi6p/3FEc8y78bTAbJ3oea6/hW4dV2RrdAqUPz5
hgJWFMWdH6jKQDDI06Gh0OnGvHYgUIWKnNluVWxUNgH7Qayvz4syek/qCEj09Rsd
2GFN5ILPc6qjd73G7T20KpdDeRDg5ur58lohtlrlTDIGOA26zmko89jGXdjgZw/5
bBMMDM3zu7KUXorlyFwGfjEY5F9cyEd9hcQ8LPVzHgZmMTnriCnjf+nkYWgv4tkt
xdHPKLaPOp6XhPpzur6hxj8uP8UM+jKMClmBqqyBHQmjQXNEKaRFu6oJNdxMKkQM
CDLLQ7lLISDYcuJzW3JjeHxe6clBMIoigQXGM/4wqEKgqjvag06DZ1ncMO+sr7z/
qqiSjOjpR77hGqqGP2b4bO9aRbeVhSNBrXT4W8dG+pEAkBaxdYYJTPBRK1gq1S8p
bc24NbUGsUV1iZU5eBgzoHG2W8FWNlz3Q/pMiCQu61foXMWwK5ScNeGeMVbezvnW
JzLr57lA9VLN3awGEzyCNhzr4+qgKhN7vTtlnUcNhoS3bEnuNUgCqNfib8kTBKTu
iEbHzOPCm3alyOWpLy9I9CQJy5LY4AM0BjPn4wAPf5kGNiUZ2V6rdE9G0sCFjFGx
mOGUyRE7a+SvfE1Tps6Rpw43nfoymIg6EIXTnDXokvIeXj9wKJgUTilwjOrXRcsA
jpa3u6eXb06c2lOX+eXzBSxzCIjxE9YkH8qxSqHxWjkQOEVAkicFVDfi2iODNj+O
H1ziTfvg6Ey+8O6mTEl2CVpLyhn+u7l/fkAKkryUXgV6cCG8kZ4TnrF8T/eDxNqi
A06pJOYkDYm3f8qHkZqS1MVW++AUFKCbNqDuHXBWO/mEmBI7S2ln5z0hzkuKFVxX
5QsnoBxpS+YWuUh86j3G241YcuKZQOeaFdMTwGj5ChWQjY9UEFhTdV53842PTRnA
iZF+2YUCuN5JbA4ckQHYDE6gRX/2tLsAocSXetJPWBavB0eHhlK3unoM1gN9z/Dx
rvNXEBNZEAY3EmsKayy7ry+UZHfP2Q0pxN0IfcHdjm2EG+mHOJTy6w0WIHduG+7M
o4fj9dqPAkYK+/bEI7opWVVFzVNBHVCSJjsaOQK3CfMvRXBQge6Xd40UlnShd10d
hbKNTFCdufe/qY4KUzhZyNlsf2uSmmpl7jthGhvxDpLCJae57ovfa+0S6l2VhOTy
YQnGI7r1/Ebtzn45l9DUCBsiqZHxYAw+zVHg/5xhxpTTMtXQYoFMZsHcaX4BWNzb
rwGhJc8OH9ePBC+wlsuDiyX7zJ6U/RN1ITASmJDEJhI785cjTvVU6oijFRNLDIwf
Z8SPHcJ5zIjZ7AimZ2krBzW+xyDLO4I+8YMXAmO+UHkZkXdP5JtsHRqVukjMFa7y
0SixNyOaw6KizAZ1LWvzWAGocTeHbaJe8a4yZL1A6U6sWWkoP7XS5aBPkqmHyIG/
0k/fSJNlO+pAZWnW7j86ZRMgfnUZ36nVHZLhXcwL9RLgNJIHg85MGezFrrz7LKRP
tZL3V/D0BfDSksf/cfKk0YOAdE7y6+uxAHNDQRPOJCKJPpVOdFwz/dpTfzdsqFCc
iw8ipaD0J3zsYmq0IAlOttjhef38OPgnK89JEIZRaJgdqiodxNB9HGCOQqiZDHPj
wPxTtJjJZeys/f1S/goTKvAeOZZQj7Secc8wkusgdf70YAQWXbnvf2LTf3sGaUSW
l9C6aviXXLMWkhuToRAQDfbdaWdH3WzGXNrNYClcuqpCKUJdpKFJrFBWj6wFeDaY
G1chSdxFgaQzGqunEA6TCvWWfxTclKN4ddCXgvGDUEY6XmbAjJMzPLb6KwkO9WBQ
J6IcMuSkQxw3/99ZQmRG2DHwqSEMsH4hfyduBTx+CyWgr84LrSCwjj6SIUcNLJyp
YMw5cacd+QYrgb3Ws/JK+PSQI0Uzp+A4y7KxQbWPxwVs1nSArgYeNeFXHUgBltm+
o1acwGM58L9Dq+Jsu0cPee68iI0gmxVjS82k5BuDb/YfbsPA6wtOPq246z0K1dZP
dGUl0rnVx0nR60wduEfkJl7y9vat5o/F38k5VbrRC/mqrJHK400E9f9uMOXhpZwO
OL5M2+lYXqQduYDiIRLxYBLDF1AloOe15YhpwocL3rCR+fPiXTPMMeoR+n0TIVAQ
j5EbcbSC8vEWUrOslRhsQ0hFV4YCs8zFYwrHewb+gu/GscKLMkc/ntbYzdh6/UaG
qI4p4eYY/uYxly4gesw2hXZ24JjQWQu/Okm+w2tSF5z4lP+VQNiTd4TJq0p/5ZlO
qC72o3yxe8yX87OJhB8Wun1ivrFaYdORKa02oKhFzUR4/HGIYRRx557Gn5oANFec
nVzuAgpiGlALdvTw2IsrMpY286pAN3S2vV8hXxMiUWEiVkp2aD5t0Ey1lSBEY3fs
vshsjqMhV0HjPPdqZrAOzFtfQ42ulLjY2CfMfMWZM6CEf+z1ckrQhLaMj1fpurx0
pzuMrMdpmDI0o7VbpgrC7PiD9X9VQ+6eVg8bV8QNunWwAgh2iw9G1SKEWg8l65kt
NuiIlgyoovuD5JJBw0U1v0UBpPOnD7OOxbvcm5Q596bIgSTvp3szSf4BKi+3Twtg
TTbUvzqDbAZvZCBdkgwxhBQI66IlDHjeQj/x9+OpAx+zFgj5Uyhjvl3REV3ykWDn
YozYviPgVYzOHggoXxtaXRXJkSjXZ2++X6jRAPgKZn8kPwOe+3JhF66hr8eWZK8B
iryC0iYKrNoFFey2e4Mq5DlPV7/G+aR192QWDYwzOgDymMme+T3HAi8Bv3lATzRE
qOVfAgM9abQ9w75cb8Gprg09p9S1YfzFIkckkVur6oIOqwrcp99RtewHwyy41BXe
0dsmTS232yLYzxGO9mVpUIXSD+5sKIQBxmPn21WT8f2t86w/veXKkVYveLesYfA3
il6YGLX1aqUqkraVOMdEkQlTf5ZsGStbD8mT71n/VkNZk8hITkSDYpJ2yH7r1/XF
txp78L2xE4x9T3qTY4mttbih2pFX3ZdIFsXqH4/c/paxzk7GNkuGFFAi7VpiNXyo
AIRc4wHqdrKx4Y3LyE4AvNsAetw3i2xo9sRRBP2IbkWIvVxIYSok9vIgwBNGRpsY
TaXlJzl2IINXGmbl3imHnaVS4sQcI3TMEHtyYH721k0cJyneRLXId4CHdTI0zpfz
jC++LqO3ZyuBPjBosbOrAfTeli22Lu9pM130ryO93XSv6YXcK6Zij0vDIsuml/eH
RzJQgjqmD/EVimB6bDZH0KXuOdCNBnTA96GJ12xWUr/TmyWRDDUzUGFFeSfNFLWi
AB06cruEEIzX3Gxhy8ImZ/E8Gn2y7u1DVc/EkSxyiqXv74zL05Smr9lZiSZ83vi8
/udCfHjs21YbBzADTJdtyGH6HyK9NHfbqv+NKY+Vo4DoewdbiCAm/MJYkFH6deZL
ITXNHBJLLY/8I6P+2KZpwXGvutA5Sgv+RidggJO08NbXdjES92u34kID4XNpp/ny
F63RYKMeHBjR2m/uf1VPcEhsMN+2qPLYdHRz+shZ0Wg+cEq5DdC3X4WesEYzNJyp
B8pV+fuV7bD30kdB+Kfbl/fBkn2yJ9TZAVYBBktfduVz324UzFRE1uTAt3eZFlJu
1+yp3ro6HPRTzmGfWB01IksQzj9HQp0x7gxkOT9wbC8Y/GxQIhYybO8DP2PI0e9W
qEM8cOOEeXPN/YPxt8YcFtn6NNWRQjoH5LkVtXQQ1moFAbTUYlruXHdcdbmnAq+u
NJ4aoGtjzjg/4zKOBPEYsVVxYGiA3HG7JwTQ2MPsGeAxgmE36WEmNyiZAaDe1wsl
ZgB4VmlR8vDE7yatIJ21zLu/i3LrZ2TjN66niJMMMd/Bh0p+tZvr/J8U5XWXNCz6
hjyGWTv8PAHtnZ2Sx3d0EPdZhnsB21rVxNSrBVxRyTstu+lgHfX5CFi+wOzmWkDS
DWtYD7RJ2XWhezqTESJVYxFXGf1oxhz7VJtxTOESCj3P7wpZNfVeU3ll8XAhm7I9
WgoIgFPZT0fRfLXTynR4oMs4uiegHn39Hedcz2+0MAisYEpOX2or1gFGLA0W6S6T
+MfE4fknQO8L1MDD3WUNhb22oPTeHd06gWuBSimh0GHcZROqK6/ALhaHb3ZRw3Lq
UfpKrRxjpcB+lBsXQ0sNiAk0+rgHDz9OD08hDpKdQO2TIe2qIubZjM6AUKIFLB9I
Gm069hJrsN0NCAh9rIZF0u063VcgIa+WyFdpeW7UA6Xf1Uq3hU3U6jkB8GJPvj9W
8BuUnddwCIDMpeiMFDIJPmeEDv6z0YbXOZG1sC8PvlyZFQGHS1x272OrjvXdj6MO
HVqN0xff8/rdR3xFNxj+n6pjwdJp2Dtz3x6fB/3gIB8g3a/VQPks9w0QueVmHH+g
JuM/paoPyTQ5kdJ2vzIhdliYNhVhLrZ7BoGOLFmKfv7Gak96dCrvVfpNlohTad5q
CuTtuwHuLYI6XvlHrzbGSJpTugZsGwcS3enssiBwoxwdHgJeJ7pwXQkA4beQIhB8
r776VcQs0IoQalsKWVE/eYyeu4wYLo+koC6BTByvpUXVCR3sQDAx9trWY/Zk2qDT
h0et/e1GSUqPF6YANdmGbEB9cjZ6kWldeLdYKJLsfy+ow1tGJpRXbepjzD9mJYYD
Al1uOWqoxtM9QirQUGvoVW7q61E89KD7wluiX03PcHyyI0UcUH/+OTtAkRqQGOFE
dyNfNViVRt6Y+ua1O+kyt8yX4Lqs+NK4tjv4O5dveZwHssTgEPPFTt5T3iPjuFJb
ru/5aZYbPnHYLNdkwYG06Qca4ZHrHkgJYMIH45/HxtV0gBldLz796dsV9mTq5Oo+
exboiT/9oJC4fiMgkF80PFTs3XTGfgn5KPsAai5B0wb5PGsxPGC3KEU4kNeVuKYj
WkjWuo/gkYJsZxUwLbVGStnEpMaZ+oRPzb/qGiRtAZT8gXYkgoq4aD5S5wsTrfCS
GXWje/SyssGLhK8aPEI98usH1x6tPeRjtjfUQCLaDF4nHbhgMRj75hNpDdhL/a21
jEYV99FnFpf93m6QpIkQCQdWK8IR7hoUGlA4uyB17Vtc6nrF4Sg3j2YmzIH4bp6i
Ya6D/cA8XA88AFbkG6Vebsy3WFj3CfjhrJKr0PR2M8xXZHIVrfexzxqfFfJpjuC4
ywlFt32vtJjccmBLT9sRUWI3PWLJ2bRVSOfbn7pPHfETSeaocQtT3aKWMNjECBzc
aZZzo/lB8F5n3H/WWdIBm/IRCTQa/UlT8cEgrKiHxfERJNt1zek5rNQiY/TEbkcM
Q7A3KC1NDRtTKc8kKttjF9cJuvLBb3PGTg4nwjWCXKYJKSB09lSGU9PyCkcQgg61
QyUMKraBhNClQSYQpAstHc7VKa89GPhekJ3A8RjesVEs+FN27/iqdEyJWJL9u4gW
p0uBkC5QEADCOwYZKDXTXHjoQKjl69taP4Xb15CMKPoiHAeEV1Lb/Fj3Ej9D/MtN
bFanmKyyRgBUgHH24ld2bhR2z5Hfw3NGA5343OrJj+MJtr7fDVNCpoab+NiFGGTh
OiJBgmIAoCqFc9Vspt7UfD7oGmarAQqKsu5NoChIRfkmMJob/FAAhJFJSzwZRVcQ
/Z+JXZ2GjyCwUxRwVqq2ZwJEFg1dXuN74PEAbLwzTZnVsnPQeKdrFH3ksB1I/OCx
UqJzswW1rW7GJpY2nODHe31XjbvMfrEMyOMOM6T7ZPhIHVM/SZko/Dfksb5oeuAY
NP8wU869c6UmJFVEl7jL837Y2gIgHfTJ2BpHEaQH3Gis2YD/0vXmsLbZuZ8DCFqO
bKUNym50/oYh+W9r3N45WEkHVtJ4Akew/yA+E8uqyGWWLwDR3pH662yAlLmHVdNU
UtBSFilrEB96GrvRt67hbdgQlIMkUzHtaayrKT1qxPjXaWIyaqWrUtab+PYWUQX0
Ag/0ByJg7O+OpN4nxb4rMPTgI57CZFNCGEOCMFKu6mfBWYQKPS+1GZko983JBQcj
6HXQwY/CKYrXeNrRdcj1pXICOliKoqB2neI0Tv2gx1knKiZ+XpOOFjwAFImXAbOY
it6tKQjlc9p0JZX61vdRootLPDb5XjG1m2irrw2QfEIVnDCSQhQzFSJRT4mik6m+
8vsmjgq9gzQraiHycjt4aUfjaLPohb2QGl6G81ccHcagTIY3NZjZTZjgaYoNERcA
fAcYNnPs0SDdeej6FOGBF5cqQk8g+p50+pHekKKmlgLkwf+1hYZw4o6qgHvuOzZk
kfxYBuffSeFtQl5aPR+J63YYHSvL6ZBIh+i8usmmARmFTjdM0fZlbQiWXj/UGZQ5
sUCR3BrmJIJtYd17iNf3jeLLX0b6Ad410sPa9yNYqoizJGGZTpEeyfEeh1hULpHq
Kj2v3wPrtPPGLFAEwaQWH4EKYHhc8FaAcUh13fz5Ku7Bxzb5mEno0H7NtpIQKvHG
Eo1t/qbVqu9kY1xn+ouE63R0CZKZZQZ8ur/snu3csPhymRLfL0JiQboOujJabAot
UnO4q6lDsbuwmdx7EOfGSWR3zp44wTzCtM0KVCjr2Udlzl77A6UJb6eUjUz3kU29
pMbusiefXOW47rZMJw0Nh6WoJWUyq/15oV/3VZUwha5r0nEBrJpNInbFPmLU+i3b
eInGxvTlpolJNzXrCuUNVmFks8SN+dSOQIp0NIRnuZyinEuKr8bviQvoqHAdwOrh
xezEE2FlCfFb9DHXSWtRCcNBUlJXYeAepvp1KgwMyvIIZi1mugASL5TMylPiBLr7
h8qUn8Sr2vIrWrXe0ueA9140wUPVrpBkqZ3qmHJls+uw9fvpbMue+ueBifkEdEN0
myoqXsVHMqjlj/wu3iuJBTslN2jpFL1LQSYPj2u6WWDArfL4XpMcprJw8Ldr48Vd
QatvWYPouS6pL3z2o1+BlSF3+qXmO5lS1OMCLl2vPy5bDrUTRzYzDLeORm1o0CrA
L9Js/11okJrd6IBAN5K4Scc5NZnUNHKZz/1VhUbZuc9wbANe79Jk/dV5aqBykven
/l0hE9zWLP1PYKres/0+gnZTRRujr8/XYPcymgWDrcVvs5LC1AQRWYhHNHCdEQ2J
D9xw9Y4rwkIc0n2sv8MSsdVoH++MUNIM3whge2eMJT9IE8+sVMHZHhbLGEZuexw0
WjaFjdPZkdlzwQSUWzm1aLiBhs4ba4Sk7tRQy9NpPHA2eiKf7tH5jB43DIddLZr5
ylQ0BnGrMNH8qtLipM39NWjO+kUfMnRlFQW9oh3fTVsu5LISOly97wNWQZqeHvI9
N8N22Vl2XiIJD3XeNslJDv4O/vmnqdLbT2+bhXF+F0Ql36vqN6wpLwpNCQcltT9J
WSbvpJQ/7aXa09U0oeoSlN6eadNRqC+Y20Ib5W+DjQ2fxS91O9s42hnMOoLPV4V3
n2zfxtz3cBy47Q09TdrxWOLYFkW5JKftsgZYGOK5i1YNBnkuBwmUNIaMOeY2JyLq
GQBpK3OkMoSPekirRQsoRMEOwQ5vRUeYYVd2Axh7xLWIVmFUMW03ovC+L8zXWZy9
goslxiNeboEdhJKcZiNzrMrf5nwOjHHza0zhCuQsZrnNh2an02APYICbmb8qWHTz
nZt40FeZ81rdiDHSdWXdJpMjJ/iO7zxL/LKzpXtrVlSptDoyG+xOx5skSEIGbKG/
a46attgQGnraaJlT4JXBhAmKj9pTqJ5Kg/8GNdAVhLyQIz4UgSZSVMqXvuaeBtn0
RuQJwoj/p8CBd/+yTwNfOpKt75W6oZawJXO7O+98dLNfzRBqIFPgyUyyisQ66DAs
3GWXGHeIrkvgYvZOy1mBtPYG3V8Mrr5osB9zb3BunEUW6kPVwrZ6Qg5PyREhCmVJ
bWnUNO4a6ncgJPAWCarkJGKIZmWmt5WFg+Z0rwzCvnj3auCxP+bLtSTqAktHL3c7
AxDrPq+fA3SvRni604+MfcbvVVsHXIN7fjUDsGL+gMk2LsMluaLmhWZcmBx4/h+H
9MKNaTiD7pIzwWiBmAjOdSNKpkIvDTgr6M00MK+BpVe91vPHoJGoOdef3i9MJ2yL
27r8LA+IFeFUDD+QiYPf5ebLye4VzlsGkGIokpMkWaHaVah+/33Ca5ZwqIxlncQG
5Hp647VIQCymYUp5Qoiu3/8mgG1K95P7whIj94AR3aPRugdYVdMXaLXbcKs/TTG2
ylPqQ5sn9CswkBMLQZzIxLfn5z/3e8eMYaelj30wQh9Wz4dTFzuzlUbuS7uKGqmp
GmkYUm+cW4DoVnyqzkvHL/YRJzSfWtW7lzrv4OjvG1QdkAwSdqf0fXJEHvPUfWUn
9NLAUFGQ7JslCNePc7QJ9v0Y6gwel84Minnld/6EI6gb4YBnqdfJkLmcGnVektuF
VqVakQkuSiSNvCOdAyC/BUYK6/+XXwxse1PiJ2nK+LMSGhz1qMmqvbIt5uT//bDG
mOrN6yi8gO+1ZCT1r18ttvnb2qdjmsF4UvyQJlEvW1oWoa3eHGwiZFeST2idCllM
6/OYlAmSWiSt1ex+JJFCCLw00yNev+1JRwkvw5E4HNWUeo5RB+mkUHGRYBg2UYkR
2N1k6WJbiKmAZisF62TCucn4LfZQRDr+D85NsNblQrTfNjJQG/mXXBo9t5fbf66N
Ogt5PkdCfa4MniX1JrF3rUEGl3l8asdZ+oeDKa18lFEuVBOlSaLgrL3+tzkgM1HS
hSFGFAX42O6B104nXRuzRaLQjBmb5ZwiBD1CnTcawIhhcou1jVV4S1R7uJavfLgv
+THOTYya+2iHmb3S1PKBd5R2hdJruYdnm+v28V+W9WAUwmJvybuXEYjU8DmH2HaB
SSI43AJn/8LMksl4CdT3zCWRJGsQxI/6UI0eaYaawZUGC35YgDQusW/xJ6gWq+eM
dPk90Yb7YS+HX99hEBlPaAFIWr11jz+YvaoO0CyG/CycH4SAjygUshTcgRT2IFiX
yf0rooQ0QXelhINYO/6RF8STujd3oNPqAGBKAuIVoenWL54rlBE+fBK9/qfsXXfe
qlOSUzHL64cRGPDuGJtXzhKlttEiGlJWblNsfpLY0BtCx9sXJwci6XeIMGF+ndYE
vuZSPuRoiulQr6NyYKw4NhSt05VUkqEAzfKMa60KgRa2x2lcpcCv6dyiB5b8HKQl
yyrMf7IhTr3XGB/6ARTo8oAral3zS1cUhAFZhE3HgpNDOpcIkPX8/4+fqxibTdk3
4pDGjEbeClJjj8tttAsFdduKuTd440zh1X7uJpqmxWZNH/Hc4siHDVx+bMgxR0hw
kWOPc7v1a5DrVP7lX7ZsliZJ/N8YvWM1EQdCuL9dWtsM1gaxSTRiEo3nWEM5d7oL
UOHWeDgoXLacubDkn/KXBjo/fDrfRR9WO5dZUMd+X5ct0V35/k2JqwnJ8K6uvDqG
rPhifqQsT2XulvldAScnos2mEy/lmDmywWxHxbrLyVQ6QwrYi2GnBY08P4kGstzV
bOqrQrfFr2sGPSZWHdC6G5mPAzvHfYYfuCGMuyfqXEAjl1e6muZDf5Sbqc1TvfPd
KPCICIjHYfg01E4DXteK8H7E4Mj7WIiIwPf3nL8c/NGsSn5fLJEdJkowPH23/bYs
epyWSJHN0MUmhnq+hgVNaPCGDNk8QGyMaylfPwGJcfgM4Fm+aKtog2rRL4aqNlLp
BYtlynFtOUoULxDA6gIezCSlBLVYQ/WHe7lTR9HU+/QdcdTdarW0enAln9Ndhf/W
SOykJJ7EBdiHrKbMxPEVi0Gvz3bavVpL+phxrOCUoeWmald2mCtqK8c7Ouctbl8x
8g/HZ4SKrJTXvsuXJz8VSf6QUD1/zyURlasn0eaY6isEQ+h18481z8MD5CKT4YSp
Hdm26ANyOmL73zgp4stZnBnwhhQJ1J034ps8rViHxXsd3Kyfou7iDo+jf2ybuSUJ
37F79l/jgyjM0Tge0Z9K6Tx+shSegD/l3R9Hl///0+gyjgfJFXHq4A/RybgTwfdK
1tvq2AQuZPBkQX1EDkocIQbVHzOvBz75uYC4gHVbjl6egDqPG+KL3KK/T0hIJY+M
jDhp2qyJ0rbn+vG85J+zvpPWptuxVPMlwUJDtcA5K8CluB7QtthWHIoLx1E15EuH
hiJLBYhNWb/fVwoY/Bk5aaiZBXPUo+xKTT23EtOjjeVBMU/rD5hW8FFmkcPF/a7Q
FwEtWJm5HQ0F04k6W//DIj4mYPgcxsguRso/yGnccRBdFfsMINOzzlnls1/PbLk/
MWdxmtCZRubILp7GGzL2WLWbhjl4YRhXuF8+uXKwrqzKtJFze1cKUixyKvr7zBPe
a1qvtsjc6RoVV9OL43NaFL/rk5RraFgvaClLUmuzgGlLvIjhlnkeCF0IajYfw+/3
NzmBl8Bf0aJ/5DwW+8/goBiJp7ZZFaLPKXMq6Hu5xgYlRnDm5Sr2VhXCejKKr4A3
mH/uF/oILr6/gYjbb0+4ei5jH/+SudIWG9q4Q0/XcIKzXmikr/8TFvb3V2/LaAvL
ABAbFmE5AxwgTYyNxSzLOmiwq/qy0hhVgFK1t3qTYzq8fkfXdzxCYodGu+A9DxYG
krNZFQqWocHrVNpMYbbyQbG6wEn+WIa9LhWwGMXu9Bwto5ycEtIYHjY1/Qu6dFe+
e86gsJG9KosQ/l8Zwfzm4pkQgKusRsZ0DwymoqR39c30G+b+c3VWXVOED3JwZI9R
LEIaXPBGBqhcO1dhnFLpWk2omutNyaZHdx9anFihv1l58/2QeGQU7auAUJOHFnoi
hsWXpTEw2AQZbyRpU7A7IOUJFurpS8kz/HviTW3Mwnrptel6qZaNl2sqcK7k7gdJ
ew/IuHpEHJdWw6jlE30S5opRxPq3EFd90Mja7Rugw+I85pEIwzHFj/VoBHZ2QqlE
ERkdKaYsftgzFFpaGU8ju4soVW2Tqgnfr5R7sBZ+rWgkMc+k00V3vCmYFxXmvC3s
B8kPGaGCiWOiHEMl5DRM7+JyrF+Xlaa/9lG30yvn/YeKCSDp8tHfDDgCJLfFWn5H
g5whoK2zdIiKkmYHEehYgQjp189g4fGywa+1ha8DybRnmAAdjiIFXXMcPB/AVBaR
l5IUu7gPAULQPfsGO7XxQMZejEpfVZGlv1RMaEloRAe9u1n6UjIOn/bKXu/7twHM
huCsYy8rY+Alahj2seHiN9sLSQwJvKh+QN5IYnSQ1mUPAJTI7adTDfi5dHk93MQj
n+J6U05PRhs4aOViy/zIBUYU0lwJAMDugPOFzeLXJidKwNAXGmj5mxVigrH+SEG4
vTxQR0+12S002Jy3Lz5dPrJnzxW3ffyMi6MFidlzcb636uNNUJXeXDAC0CeZhELy
kqBrMqT2YSF72X+q4SlZ72k9zQN7t7mHhBQ7+5tkyjGScVTBL+idgK8UjhyNBoIX
btHxzSCJ29G5B27VZNVrCKQKVAfCV3MdPC5xSoJoLm8jnUSk2UsHFdo88BTl5ZGY
Av8RK8JlYWfpmB75FRqrSam8TxVfu6l+aukFDc7MNxRWkAUMEjh450euZhbIOq8G
PJ977jBFVQ23QNJC+LUZu1QXzxVS3GscrgYCNfakKQQOK6LoHphnZeZAY2i3L5rE
jPzxcn4qC++phFYYTJEZe6PoO1bVTEJ9nJsd+jRUXuFC8EgVKgp6PNeAqeiPaWGJ
br4OV53nkYvR59yrAvhIxMosl0DKY0VaDFwTQig0Euy7qoJoe0jA1UiQ89Cgsfzz
Ri48jxWhYAeP9FBvEiepjEbLcg752UyN8iSJJhnqPZonfIkZr3RyD9YLQsfCwCZ6
HRvjwhcaIkbih298i3R1fl+Up/5MlApQM85QT7f8zlOUfAReoFnVBOba2TaIXUKX
EdNeIYem5b4DA7znIku/bKqTELOly2fHitusCAameq8EkmEk7E1eqSjaEIwpnbSJ
MqlFuz+FkDUzdyzXvBee9yHT+GdIot/2rrAZwwqYsu/fQvS5vGEK2Dug/23Kww/H
fL8oJkkOBNisHOKgQOETmyWNnQIGltQZqntFE5J3o+bx3Op/TB1CnoZOP48/FPMB
KL3bWP25kToxuJ/2+w9BpgHx35voJ5loNcnsF30+iOah5jjf9xpAH9p7Aml5t+Xj
3xYfbLIYH1cIYvlefwaA/hXP7wccIDmW+/6SLdmCehtWchCXCOmUZoASNzlOR27R
+hPMnmQUSEMeAWvwOM2RGe9gSRfiQ+/qk0g/0P1+3JNAt5MduAKuuD5b9vHNURRM
6NzdtpeZ1CUhlkgQDX6+3L1R7RZfZJN1nxdYXwcG2og9fNLPJE0TspmOk9OC+P1S
s6dV8BgaQXvnHcFrOQvB6dfEvqrwyLUO8KBKY7Po8ovuPFP3sQ9vLgKnJODee2NT
J83rSp6OQpr63tZ3WlJ9N25c5cixhXSSBc55FCEKLMNnGF+HUH7VhjCQEJPx7WRL
Ld5yN7MFtSntjdTh0NxX4+NEvr+Lo9tt3neNOEtna2sjr7Yl7itJ5yGQO7L9rPZ8
s/95rwuKUjxf71RCjKwnR5bJTGeWC3cnwNpFfzBdXNk7IWbV7s4Nv2sGYG0k7h4K
3AhDcx4a+fIS/ea0ALlUZIlRDQi/QM9SL/H158gyawr4qbAtcw5g7Yo4q2XUQogu
fCt29k5XrBLEeOUDmgDp/jWwqCSiqMePqktqtf1qfhyetP0eWsPBJhxfgOYx9F8G
ncgWTB1X+UVuzGQUyJkURuM4+ab5VTnMXhAuZOttFNAF4mHlU7e+ZfKzNizN5Bbg
uIJ8kp8W4s1ERaR7qPyJqSy8QB3XqWnoF7zw1T+plStGXp7KSWnPGnfqEq+YTrWU
62+hWp4r75BFcS+6RKnOnRCGtkeWye7ApzOScDNfJzJJWiraBUx9B5hFzSYFiEmb
a4oKBJA6Wl8Eu/Sty5i2aQC4yxbvtbA2cr2uj9mttxFH1N/hx1vT3Rn6hajiRcvK
ElFcQIUVHyTlVNWr5fDmkGMq286sN9LVDbDT4Aj2pjrzT9UKtpip08imrrNOEP9s
7ZDednV5y/ndZhIJAmou3lcx/vq7Xv6RAhyaKNPpuB2daEwy4f69wbNK2Vg/afWd
RdRvPBOkKj4IBgBKtT+zngLqKqZDyo/DHYYEZXdKvLS7TGK7Qb0Jzm21YqTlHmv3
ez9uSGC0PKO2zsxby1tGLaxVjNwfiYzeAcbsIMU9/FT89ix/XNkUxUZdyjW1M493
LqBPNoemnBrreGFJm3cyH3SYWtRMJEzkns4frE6vu92XfnbboQGHk2haY/2KPq/8
SAxDEjRCu2lk0Yt0Gc2MO0xQyzZYZtsOzpYeOUybTQoUvqr1Om2WbCWkM294gVM3
PKp5eUIEb47kYa4u9h5SJj1nJYaBAC6XzmnA8CDoR6ZATRCEX72hEzipouQ8yGXM
+2Hmu8fz/tclZi2YzqjX6UkAIDHpqH4/NkkQomdSISWhERC/mNphNInbMRGvdPJB
xBrPyWs5PPSuzjn+vW5EqMqqqD+H6St7af852t58YxgMlV6nzELsWPdGR6vIm1UW
WDPIgQ2MiOdSdocHtBeiS6DlCh19AFw63UDGtgzFRDSipFwuvLBt5r+3mesoxwxg
jYpeY8XpoRjNDV8oeV3K7/pUMFn985fOVi2LHTeZiXMHq1UuhB1q9Sv/7oVuKOue
UcTXKVwxyy0+263dNOGeSwjbsuuY+ff3vOWk72yXcN6EZJYuaEvky95yZ5r8mtpZ
gITemZlWdVcshbkGLLRssmdwrEGidO8ABKxvXNPL9MwnFrLMGxClvY3HFsBJJiLk
GSO4mo3cn2zz4L98NtNInPHgm1sqbsiSijdhbtpbYL6EynHb4rEBRm+qLp2pXuJb
8NIwN8zfNXwyS6ut68j/8G+UInHBzRW+ml/REYsys1mB3/kkoWMNr+mslNnI6qqn
wKvhKZi5O8dykahvCx0nTtaFh0sBCKeLERLYzaLMiJKsKddEFebWaEOvRS6q6Hbt
JMMkciOgkYt0YlZGZeQILSCsZjFiGIEEXPk5PAP+ZQcrEBziSNq4He+EwUDOs7W5
Byp/EoaI2SXW9QIaoT4T1qHDjK8WbdQyzQviJIXx5kMIXqYvi0mlGbNZTqkzj+Dq
dcwsdU/z0fPXdylwTCrmb2wleReI0fexxfJVcXLcSsw2vHJlvPHqe4Hg5Ji5DXwK
OAuMoI8KHowr+P2r7sFS+cyd5BgeCUQeChyXGWc/wzMI+5ob6Fq1wzdXtOEJN04m
OOhNXhNBKmw0gO6OhZJWXoKg/evMEhUpkU4WFBgFqo5GuF02limDKhrdtlkvs9+T
wLJKl7UeyoypnpQ3C9Iwpu57nfKoIiJ6GmylQe9m5TqWBTOrOoIvdEmGaQC4ALx4
V9DwW6KgIUqUWRwLf+EdJIUhR4su3lxspiwPLDmQiOCTF+DF4e1wVqosiAbaRaPy
gcxNUtxkrjcX5Lw9MeY7125nOKe3gwN6NqEMiA8xAd9aULOM0rHv11VZSxlp0XWd
+CUlbx4tTLLy+5H65K0DvuVgpcqPzgNK9Kb/2rMe7YKnKFIh8b6RmrS39xUFyCoO
06plTXipWAZqQzLM1ZGi60o5Ax+dfOfmgzqyxZaMxHhPlsXf0PvQZzJmQMfo8fFc
T+BSAAjZ1Fwv0icL6o/tIrdauGNFVyB07yydqSX59+QaGjd3bo7AU2c57iQ7CtJQ
WB1fGKohid6OE4v3pBNAHUnEi4ce4EIG3SBpfWN3KofgSA/X+HFwgyOZzIfQQelJ
vWcI02zKBis5or0rZdCGIuYYGSyU9o8jj1MUNp94oTJ6bCgFuo6Alph794NV5jQn
eF26moIc2Lv7YNyZteCUMW/AFL1b7dHpJa0Wg5e2EwGHRynFX7b59hbd1+kcO1DG
iubQLtnp5R6x+Ir9ES6ncIWlBvbDDMsClSb/xRuVWgENRUgvxST3L6ZzlJOFawhr
lWw0I2wzjWaiTGubDy400ZHBa4tU7jHTCgvim7TTV2wGrycvxhz21NJ6k+nssOG6
Caip/W7s93oR8QaUuUfiTBEY07rJ8uSvxzYU2WmqqyvGI3fyS2BpW6HFczCrqYv+
ufInonyQw1jtPA5xuzM290LVRMh2n6NEtq3G1EuL9+ZOVnC6SzroKnR19EwlMEUU
B46NN4/Nh4cdg88VqH4MgDd9vcymS6WHlW1Q5NTPlDCIZ7EwjFDJs4rM3m+8MH7d
fE9vZn1IWfIdUOA5czDVbtI0hPlhEtwYZiasfecbZz2ddtV2lG9AE80yhv6ow+9i
oCu8lJb/Cmp87q6hDPTQKNfu5TsF9W4lWxyHPbuaRA6dhfIyoegW2FcGdbpao9P2
LyBRiw5WgZt57XUvQMseShLHET/JIaotlbq2IkxWlUSRQpwfKdxFs9QMwB5h56G6
rASu4ufACGknxa+897iiiAN3vCrkjnkV46LYjQHne191kqqjuafu0+d1weHyZWTb
PT1XNrbt+rRAdxZhchay3jL8W/mTBX7Cwv9BXWfdrXLqmNmB9kKDwrJdxxV7SJxC
Eg8Sni/kQkEp/3FSaLLFb6QmSls5pvpnEBnRRzGBxcsE6vlxa1ZdBo6nIW8PGvf7
X21A3Ml+Lr81VQ8Kd3/RIzrLXVzFoNwP2PFCFnZRBf+9BOb2fwfRrrFBpRaNphJl
HIpNdrWXs6bGQGj9imXAsHajbXRYHZ4LkUI+gO1geKyuy7WGvizx6Z9Sd4YQxMGx
iV+bxi9XFLEOTh8Es50UCcqT9pO5TKZEzzhU1Iscnbg8VcMsRFcZi3FiFkoIps5E
lt5TECKUoAP4/7hrx32we1mLJm7L/B1C5y+NtlrqUAmpwXwiknigeFX+uJmz/lXB
ABijHHZVy/4/bVtsPivFnxOmQMvhJbE6ItroU3O+HbCq9BIdOOtTy5QvtvmyqrUV
lhPlXN/snAyrXakdL/zESHw5xihIW+yB3zNsCDnq8AhWfOOU91VnxQivtHJUKUXO
tdB5TiJS7HIppql3MuxeZkXdTVbR6b8/Q67G0vaGrd146ZgjUeVaD3MzAKMGNeIz
KFwukqH1HVCWBKP2V00ewC0epJZTA9pkKbOM4WLOoMH29OCpXv3jHAjuJaklngTX
ow1B5yH/VODSN8obg8K/jNHB1YJq8GFM7cUY4k07gg+XLzMaXt85SAp7UQ1dfuT9
6Zlt8SmA2qhf4k9HXuc5Zcn0O6dLPrn5ry1ijPcd+E/uVT6xVdY1nRKJRVzeid7+
kzTaXkFXVuMh8A36/awMjtpeJD1eOEGW64M5a73LkJUpautm0NfGdmIEYwWtYBdp
XBKBQN0qDf+PaJrUdRhyYpsXIKF+IVuvzcZFA7Bub8AmbptkDG5SnnAwAjOV+L3W
ZuFOs4USlXj6hcbhEFWCfFxz1wTxNS3nfBrlHW2UdOLA6w82M+prgg5r4tmB2fhd
fu+UwlndOts55EYBcJgDY7crCbF1tOK2YJxuwo2Ka70VS+dmmHHy4F0amo+vDokf
xiZ+6r6ZO2C3JjiIz6oxwSjnd0Ilw8i9B2bfVjPtSUXpii8WdpaeVxjtB6WzrSzB
esgVDHBV/oGqtW9FEujgBe2zG4QfHaQNuSKHhoqbsXUWRcjRmuYXhCrJejnmkGq8
nVWv2h53r9nq2KxyZXu4Ha2Hl6K+ChnodzVhS8N4T6iq5CNijOqvHf+MptTUFycM
+IutUEwF3Zs+xe6x6uLfgEDvcabnOLuRR8FUeYcDQi0U2Ym8gIxLA5vtC6IWOY5B
s378fpPdoA7tOSIJ1ShmlbIYX6nV1Y8DGK0v09otUTSF0xHKR/I8LvqrfNlIOBJG
L039eg3RK6/ZDMSLsriXlDdTkXH/ROpAFy6pyGZBimYpS9S7cyWOyKi+pJd+sG+L
XwsTaQ+Qndpa7QVvqvB/tul8sM9DAgOnm72vIyyXOI1ro/iQHtNCqEWJj7jDCMRg
Ynk+j8ljofqBngc48y71RXz7PYnVlR6txugDcXNNgEfnAmx12np91bg3f4sOftLM
4Ljhd1I6QW5Mx4VRvmkWgmRPp5x/WfwsHHKvRpuzQeD7LwrvW+ibFs7rxz29/x7X
zFoTUSv6jLnJ6A/pLapVXOIOE7WoH8jUCcL16XaQxc1lAq4C8Y6u6p+F8gp7G9l6
j81sFnE1J+n3ES+3sJf2zX0ZPlcB5jLe5Cr4Gxb74inEzPdG72hKoO9ToaSAyWZ2
lW6IiNsyB/sIuRKrU47Mij5ngJ4hHdXV1I6JXfQU1QcGqpDnNByIGoPIqO6kEF7u
LwpFphtEj6sc2RJ1NoqFPkuFhiZ8eUZoRT89uCnsjyFj4WMmBYJTYiDnswRjvw8L
uuKTOvF9fGLH+3c5H5cLb4vFWOVYkO56ECvK2TPrRXt+eLjFeVOgzrBn3M05/NVB
zCRtaqLFZ9boy3UDrzC8LcGmoXHrs6zrl9dOK/cLj2y5rejUR9rB1ZYDY9/IbbVf
IHy/2CVQm33DYPawvMO9rY3kJW4vYyLVnuWIdpYWPbzr73iWSJjUFneFnvj32eX/
v5klk3SjnkpMlkUwLRR3YIWQQ2asRNexNxBWFWRx0yjKYRNacHed8+Yz00tenNih
sz1MSgHs3sPYSEpUlSv2khUgA4eKUDO8Ush+UjTxpMzeHffGQ1JIMTCJQBvs6NNC
gjhEEYhRvwmD7sqn+g1SiDCS6/5MH25TWdG8bQAVHgt/PTksFgzY1U06wUHIuTwo
7vREc4+tFsyw8/CRp8xuuGx/1CtPLmupuXgyoNb1+UJ0rgRzjt2SwZlHwM+BUHT1
kCrLctkJQvj5JNCINd98aBkfQ2krOzLTU71NRlk4ybx5fe847uef6A6Rj3wd0N93
6wLNYJTFtnNl+GuJjnrosfO8ma2JFo5VKyOl+UowFoSFvod1wgkquLdnXS2wpWpI
f/uqcLEU+56abhNH+LWfewmf2lIu9hvG7CsYihZVwF7Iyzch9lCyH44QqgBjpf6F
5c0NXK8yISfrZ3alvci8u4Pf69pOY2fEtg74k2ohi4k0D+HHt09+q0ywOsUzuBls
8cU2ieHORg1ZKhzbZtOowFFxaQV0WS0LPHoA34PTfM8aT4BD2ReePXmuSdcSY9pT
MBqU8zGHVK7N1MHoEmv7qgVq3uNm0qd/AkYONZZVXp/778kNAj5wM5/izgeEtGHT
YqPaE5gAfuu/BGD0mo/BPBETmrfuUN6LpS86/VLq2sh31+/Q5MvTp6gU+kvCEFnZ
509EpYC4lEm/cNGy+4WEi7jG9VKUie+n8WtNTY+b5Mjkw9AlY6Gr3oiwvP5yrG0v
HO4xkcR3SD5HshQ0ql32qCPA0RJJXcMHAGBNPTJuxyVkxG/NACOTiqRZOdSZxXPl
mRR5V7BcuwW0+t/UPM1HDleQ8ebpba0fxCnP3Go84WZudVsP6Q4QfIpAJnHYhkQr
2pXBI+2cDPgAdV6CoYeNgf1Nh8WhLbSlBR92ygbNeYoUyVWUX/nAJr5sZ5f8Wd/y
vMLBaiEdzwWRhSM4HertP7006nAeStyTSQoXknCJuB5T2p4NFDOHCOnJeuX17CYz
m8v9kYvoSmuZxo9YGe2U0FWfEoJVPJ0PHvMyrrOXV+SHmQw/Esdi1/qQ63CUTqAv
L/k1nG1YNjXgsg5qxyYIB6vyBpM3cQboaDaT6BGSsq22ZmAmyI6KahZu5N9OxHoW
XW2k1nDaJ7YOAOhe05pKprXgK8Nm1Kul2+8dyDjv0VGUPkpC40Bqdsebx7jxWoGY
rTQZvs3VqwonaYaq4pEQlYMmWA8aKXnywQLzGlylRFCcPJay8l9QiAHaH9KN2BXM
oGcZwD94mIl32Gni9L51NrgMPnUBF+6lcJtltTn7dbWSVuHz60ji7fTDx2VUQ1Wh
OEKIbA/wH+Tg71bkMOuJ/PAH10fx87Zo/qjB9Kc80t0YkR59UUo8gI5v5vOCCS31
+X7oRKNzlUWwxXZ6SuWGpTCOZudaBUXKwch0E5IFEC3ub9Q8tgkDPXnE2TwVNNBq
1z2bfOTgT+eQj1JfaLNunb9WH92vh4XQ7h/nOM/5Qdp8Ac2lW7DwBS3VkQ7TCa2D
a404l02Fv+5zvhWeqBRD35uD4OdDFwLhWE5mKpr7bUTCKcpjbEmgq0QwRl+4Xh/Z
5HlFIXHAbUwqsk2k3T6dpjpESkV13REG/RNfJj414ZAaGX1UTJTu4+/Tr1McJzAm
v7JW5ZB8ye9kWIsPQn9SNeYePjwootCE6TBquOg/iHL3fKoZ4sSc7Jn6O3z+mYD0
JAoF6BtWISHyVqxkGvujMgm4bZStXI10ixa3efzC+bwgob1Vre3aHGixGCACpZnT
WMuTpjf0UydGoGDfaqf/+RrG0OfoYfKkfw9Ei03QEXZWgxUQ7dqo7bEBD8ZzGeJp
GtSwrUJeo8huxhmiK7a+qFTupzUnX+C5omuFW/FovUwD890CU1+u1kuQBEkPbE9z
RmaspU/a7jnEh3ACWPni0iIYXiow8ls6ANpDQKxMjN4Y5VWC2+BCJcljdOJLnYAR
aNx9nk0YrrIx5GO+1/q+nbekfadcwJ+xbfOT9kUU/IgFwQ7KMRF4wr8uPUzItTuN
Rt7DO+RlKpB4bTWkZG3yy/OGIdCm8bHMxDWAbqDLRwPGYHoL4Jt6W2zrqy6xH1w8
XhCL2VPph19WaqVY9wfMU+r/f5qiCdRoiDNeFsn+l8Sn3NuS+/fTZZ5aPLgOSVeg
VYbZywQGgup64kaSwT73lSFTOoWgw5kUhcoqGL09UrZSuZN55V6VJVqKXvlMogrF
z3rgyGfLv9H2ooCPpCwKlwZrcVvdG1r5ojUUL11nv71WA+Fgr6reW7hxxfKCCqzr
mle4qyJRqEOO/SBJlwj2gJp15gDDmWK+anr53rthgOyAUHKvB134mNULKiYpNFpM
aVVH+39CBr7J7ch/z/zuvdQfSU7Q0njP8DGDCQPTLeH0rNBWmHNxAdaqJFk1Hcna
w17k0rBkhAHC49MrNL4/H9GK+BrptE6jb+dL6jisgKKVY1oD7HfHkNC/ZUxuvRq/
oArihyXeVyatVPnPwBtmru8MrDddw3sPgBrty11TRp18/wtK1pUYE1lrYuF1ElqT
IUkm+YGxKf6TLWf6NjYeYnZU9fFKh2duFju5CrGsFrYW4rhVyP3m59NGHH3O4WHQ
unOml2SzBjLWTzXLu+BWdupewVnUSe23lGK2f3Tlu1rwEkccV94mCP8n0e7gkXyU
Sz8ypCoP9RK+v4+q2V/RDyT4TEl3Av4ILe13pvPo8J/OyL695CwqkcPDpGmHSwdI
flBX23e1GpsAYfmlMPysPNsg94KZRB0lG7KOMd89y/mauwcIscQJwL8iOpGT9PEt
a8jT6d01VF/Ko7H/Hx4rmmizSgoXUqmagVZZgfPgkTr1svhc9Sjl5cGloHGpjQdK
/EYlCCEPl0ssQeI/7YE+HboeirR8m3xWsvdzWmf+j/YnK8DlZdyvCoWhhkdhCtIb
KuyzHDu1UdWvKReRshukzlPpcGoBPeNvSVBaYXikVAlcVw+dp5dtjZ8mcueRFyax
ap/FFlONtRh7wvg+8Xzt8pWVJCo/WdtzwmnKc0I4ywfMGzPVrxX8fGNDUdtuztHh
+ckcUaNhcoKV2k/tqYnY/uATISpdU4obHEJsikw3JOiAadGgLzKfkWwwXwQoOa8X
Gc779f1uiuDP8GS3lleB2PI9SjD0VTcTZINaro9Rvak+Oyg4ACgG95rFwbUimYa1
s/CBvFMcyA9GmuowWn/m9IlnPeCkWfgZfZEIVTs+F8ndB+pqjIAJU/hX6cn38BTW
oEzZ4MZgZJHXfTuJyEe4cuda3yzDxYyixAlq0w8UDQLZDXLOiRqYbGsmkZzgAjuD
WzanZzsmjBl/Prctfzm4qAuyKHVDKeCpw/Ph1WEbF/QzxM8cwhcghs2Khw+oSdTT
rpC8IHPr/QZGcb8PZ9duzmAortgL0e4mtLBgq9MgVGXuSdEGoWfl2KdJO0xE7Z7T
/su1auZBuvGnKoRYfZURc7ZLu6Or/3VWD84eF1AEQcRCh1ghOGyy4bcY/IiTR9VJ
EDNlUB2IHwvAz4ENmvE9ByxKQAgqRTN/6bVShF7yKLwR9MqailA8jiWYa9Ra1kSM
ORIC8x1tdXLpSCTX3vsUoh1CBPzT0y/iA5aNCMbPj2ivcJepwOQZ61rJqh6AhBV2
WrK+J9DyFcyG83RSpDyuF4wYdCOb0rMzfcZprGZL81CEpbw82B33PGYxA9eC2JJu
NLtdUNtwu7VqcpzA4dFgMP5UhR6qBZGMrjG/H3nyXeAwTuSfJ/OCN+hdLPkbtDk6
Ut1vXnhKDu/t8MiJgp9suamxlmw3+NqHzLM4XwoiJWuqpA6EfbpF+uIuwDeuNB34
zIzYSIraGQCQ5DnzMbjYGw/NDfpe4BwMTW23MjfJpsGpxLIomP+RE1J/JqRqjlDL
8C016SM3v/Uxhs3x0K6RRCh/Ca9Kbjdgk7z/LHNSJ4MOgGD0Y6Bn3Dc+t0ogU5T3
jPNvmSJFVI7dWfythpPS76pFHCwBdMWaYPJfOaMS1608mpsmY6dTSqBbywL/2ayb
S1jzIlB6MYK1o7r2jEMZqizYlsRbs3r08q1nRu359YncJzvC+7zgani19Ncu9o/8
+rq83GW/mHdanjx3l9NyNyGN3VkMr9APvT9pfeMUfPgG8zpae4Jv91lJ4xoV2sUO
NDaBpwQq7wRe/QUqOUa/qhIfWQQj35FxvcsSPoIKwROQ18FwQFby9sjnYrojsHet
kTzhACOdL8ac1HgU/QnukqAiKsx9v3imYPeKX/Tvq9+ceLT6VGDTwES50AeFTbOT
J0dn9K/Dtd03cCtejonML2uSxbnMMtkSOdZ9Y7nBLaEx6blCT5hjSfRVFj+vsq6O
dfoltUScnagmLKIvX/OYY6wVZGdevibmzBMHznZ6dFPh8bIpQc9DuNx37eFRNDsu
AJwtZAI6LazJJBmCskxBRQqxjPzXHGHwfkzEA+hPzHspNQqLFQQWWU08hJJgVzN3
uItDw0RgZQOSrAAPU4SQfSYC5kcfXmwq214GPfJa0ibOLA6S9ktuqrSp3mOPBUN3
Wh3txq2n6mN+vXfZHgxJhIwqIqIX4/gf+5M8lfugXv5XdkWpMQD7zgHiF1n7F/Vr
NfUvaSQ0e+Vfc099ZLbCB+dORgu/36pu7Ys2VAKPqCNxZcGj7PwxLypf34OFY3KH
bLKu50Jy7Aw0rYnTcYgtYkAuuJXY6m3g/yw+fQMZBGA0yyMM9DgcJAbVNjt1oboO
P7HDRUwql88nOD7rwbbcCe0DNL24zqMRgMCytH5DHECAU3e5Vg/a/hjnrBVWo41S
0gLatvKxYGMPhJbTLGoqfpLnRSu/+Z3cYmu5G/niGZ3+23OHpiaAk7SOHuPP80FC
ErtiDCQJ/Q5sZWtJZiAwd5v29oSi22eT8G9/M1DMzm4yaRjSKtkZdyrfNrRv/WFt
lf83JnpJPUxyTX96vDm90AYgSI39XORwXDVj0AJmdms+CqmphwXJ9tsiwR1BYGk+
RDOByZ1qkMdCKwWNH6E3+JbkeDypTcAzpiP872D09jYvPMeAL8gsQKdnIBBnCnni
OAM9m9BYzAguNcFliexuZqUOBpcZ5bNJCTxWGdNcqGun2rwGiDSxGYj8UyvbtQwt
sk9sS483N5GYH4Us0otElepgH3uluBeuNzg8W3oEQnS/XP9Zz0O7z6ZH6acpAR8n
oS27cGt/syHWUb8v7UCneLcJhfqeaj6JAHmEQyNt2kAnfrAMzdDPxz1phcjOuFb+
bAgWexlwwScZOKV+0I8CrbfYSnyCY3ksI5OpTfRbVTsMabHWtsLDqyks5K7lM3DI
jPTZSO/Q3iJKA1QntTbwlhnvoykSYldkOa4P52ENjav8HtFqOoiSfqr/2f+vwzxa
oEdXCY+urrSmZ2s8g853ZGATNZwRLid+rQG2npva5ONYL/C8u2SHjwhl1G2kze2x
un8q85CFgwgLZ9E6Moqb4yRSxI1/M7sLOyJYGGYep/uqEy/Rei/OL3DFotDeGGOK
0WQzk1gcJNOSbNG8IxwMWN/cGLUmdryBTmvb3hHhfV1v9O0tAWGFXKE40xDQC3D/
5iWr5yGdiMDk0JvxDOQQtJpZsY4sE9QQzhDGvbXf3NwsYhcC9Ay9U61BXM3uQRhN
pZG+iDJxa8uQzLP5TAKnSOmfKRzgkIgzPLvUSyStNrcfw19YtmkvyFUx5Ej9K4Av
KCdqWZBoGGiS2xYOyJqDqPoAC/R0rvK+2JM889P3jewl/+Nd7nwtMaidlClPQxJU
KuY0fzCMQSKZaWsqGL5EEMG8kkKAnP5gaS9WBmNQd3TJ35tUuanCZpWsW9KNBphb
cp4CHfuf794VHwn7sa3UaMEdd0Z/vCLkB62KyNBrWvfYwRp70YINTKKlKsz5fvLW
AuybqASO5Tr8QEoFHR1WGX2NDxgpqELF0rpWTOlkAJe1fXP+Zr72kF3jA63ejl9/
+VicD+1LBmBTD461YLutLAYeEadWOxFOBJLbSg0nT6Rs/wmig4dIYg7JA8IFZIbB
wGgFgdpyFvc2AoKc8HU5atHxyueyu3uv27vZnpR2BOiapZHSf6GqPJmSpsW0o15a
IQ2BXqQoeQ3RhQ4e63M7iFD2T97MVVfF6P0ZAe3t15Mgc+MNrrNopuoa8REur3qB
e9Hhy0O/2A+4zi7pbGd2fqqI7UBCTonoXwVaFb/N+0wXrJBrExvoMLzM64O6riIM
g37AjUjThPqdRAU5SLohPjIL0ss0+/TnY9PGdkrHnX9UpQ0aDGmxgl0Cxbbtlvmy
r2SBCbMSfB6G+sx02hUhJhRp+DOvP9Jo7GNf9PTVhkrvNzWxo9ZVXp+YPi2piZgY
kfv2KStxBcraccoxnvQvnNDngu4wYCfx9b/8ES/vIKJ0ubJeuRdp4xZglTAt8SlV
8CDGDxLUGafLBUTfDyiRX+gWTnJP3U+9mY/OvJA4y1Yl6NHzssIPyVWYJSL6lVmD
545iPDDd7pIesYkpeJFovr2iy+PkbhoApRrjoLS4xzi9yje5AUbQaAJtwcyXVqgz
7KCv19mH30FpiJxpkiyOEdXHatiftDa5i+umJp30CSOBxHBmIFISAi/DObtnozsK
Rv66xlXhvnJ1xJJRMM5AdL5BCk8OkbiFgdSXRrv+TqglhlZLTmio9bPDS/aZUmis
adqdVtcor1E/6+Z8sm9d0nTg7Fv3W1it1BHhykieMJyXTB4rH7swkfHoPAnJEliL
n2CFfNl4IfSXPsjNFfFBozEbgObDTNZNS+CDPSdXq1RG9XkmoDlluLNiw6Bo0AEI
aHytxYaaNYTDn7O6sIa6Z5Z1ZXV1XIVcP49A58fHdO036GsYsrJC/HxCZNJ/1P6i
fe/0Tz8qap4yARzJcojWPZrjQPeNWV0wqu2PD31koCvaLa1uj+s92jBILMFcOqMN
cbhZZQty0unfnKMVxlTvv/pWeDyg6Ez3ocpUNXFsoO/PiRFltfvBSa83g1gVipSQ
x9qoRFSl5Mm072BMINNXko/qT5uN4sUmKiE9zPK0+6EPGNT2tTRcALl0/rTwM96r
WpP7IEhMeK0hIBDv0G4g2G6id2yBgREthE9OwrWi5jovAy8MO4jZ5dURujoPjud2
SbnKTeSC/AYiVHpbqQf7WaHPZALMwGFqScyDhYpL4uDAVZiMgugnX3kvKgxNf1vv
kNVvSfZuwxGzOSTHB0ZZVDeBQ9LSCDoglJjut8h5T5pA8sqVqHzFCpIAYktOlgJR
wEz5qOd/L8Gd3mg0nnXi857PWet209osW8T+G4tmi93qOC6teMbzAO0z2PiU6p2I
FJinjvUUAKbpf+dp0pAdNzrWS5KIeyHXof5FkXYqivcvHwWhCIw4gK9RU9RSN5vZ
VQ/kQ+WOOpcqzYBpfKayIyMm8+127I18g1mMoBc892uJ8QIs74XM6ooGt17a3eXY
fIyJtclEGOqcYeiEjGIZSq4pircEEGwMGpj2IRZS8ICRbJJJGmgpLoShIFX/uI7H
piojCDSjhIzy37AYSs0yf/qGjrnbu5aetyr1DDSb/7Ite6ui3sFv1reJkY1K1c1u
ahsbcXry/9qw7JqSjopq8yRjFZzsCiX0eFWv5+xzw9aR4F1ao2h2LrRJGtXJlVsG
Hv9hgPS1ZDlREW4gt/659MjlWVSiWcJy42kchLGGMdb0pzJe8zD1FQjih2XFSI0V
/lP72WJQ4EnlT+atb1O7WfHNT8l8LAAIOtlcwPIcvHn1WW1SWzASs6Uu7xAnpoRk
TpgQL2nMAXfk60N4kDZNgR3MEBxdG3OdvVIFlGsShBhJb92lI7FQiFMtEXruQgqH
qYmDQjziHrEafaj7ejz9SnS+TkQX4Nt6d5JVFvG75Nbo3mkxZxJ7NYBiREaooS97
OYb/bh/GEnmGEuyaW8deI/PqTa8PTbadWIpbgnp4qKnkiplMMnbNKZAIORYcRQ6Z
eFO9DotbqjwWdbS1vduMwFTLajwp9CD/hSRtozjp1EXe7B/EPFV/Eii4EQr+oa7A
huUbUdQHiUV/dnSwCf/eGlRctEAYgSuVbUh4ncYJdf75eA/4fIx5KHm89QsR5nA2
CqasmxtCHJgyUKbFyrCFJWEeACSxjVXtigyFYh970RfSCzPBDmObtSxJCMceZ0uh
iGNOGie/6AP+MVqmxLuB95VqMDqEAOc2W8793qkiSoipas1NajO1eI5un6qT94iW
1I+ey1/VzrAUj8iQMqCk6Uahvsh8afS/HRXQxTLT0FMCt+j3Yur35rHAbMqABX8K
l2xDQj3vtOYeDccdptpAyxmJq7wrNg+RiDoA2PluTt6qxo+swCW/pmOO7VaA2Xn8
PqYFRht7efCnSxsfwegnST8eANRztsCeDtPh96JWCpeAbv5QpTQ0RwIqQPpK2+f0
We9N8cB+Fy5VXZjjSgawPoUulbFvxGy4YpJFc1LeMZO9/7oerog9g5mkIMAttDE9
+9BaIsIWaWOzyu78fGIF9dO5lRyr212zt+uBjEvcbpUu7gy36CA/am7pyMDGC5JX
I+eMhufB9VHfEENqntPn2hdNPswwSdKGHwdSNesVXRF0rUzfk+nCw5cGoYaze0pJ
5Eyqq+jcmHSqTG8m+yW9rAXu8z613g0MPSx0x1FIs4UscN14iwEnjVaLQ2915yKI
59z25CwJ0QQ8xoCHa4eX+ck+YaA6HL4RKvfch97+uwIOfd+teOwgrmaT5O06Wnpg
Etaw6aNG+6eRFJz0o9AeZ04g0QxlXWpQ3miTSoqTOieyRKzEcSXHyPbjsbA59Ohr
ddPB1SzYVm6eJfhyqtluBX1DuvqynWGSyCvPp38UGB9AwNAgBMTkKwxfPKMo0js9
x1hoiu2/dC0gQyyuHRuabm9Bpe/WcqlfWpCiVieAIL2ZmdjKUQlYTCiyz18vhscY
ikCFetXona0HJzmnvsy4tRG3BQAEMNupvP0FmHmOk9VgoTQ/ehJjlDudm8h/2YmU
pn2uVy40CEyrnZT91FRjKQ4tBhoTJPh+Wm+tOIiCM5soH1BCLC9Zm6W/6Ubl2ZN9
+ZLWFryIVKnHDnLgIURi01CrOvKeNH1eekDTc7EckHg9inWU1G37WT9xDXIThg5E
9b7t1WfLGTlcxP3IVKbFenBhBxzZM0Z9owkNvPXB2XcCNVTq9lMos2yO26/dlGX5
JFO+/3ZlSNBIIfedeRVlFWMuYIrr5BOLIiHjWDsjHN6l9UniY6sbYdpFFx2GEueF
58uQwP8eJUw0uC6hfF5k9/P/K2n4ev/kIifUrhR1F5glkgbcISn7P07PVTIIetBY
WShAgVImVmlGFnR4elfkGvBLJhIg2HnWA/5nnbnqWgXPESVQgvIBDemqBVnPICwe
KU+mBLpyxSdogI5ifyAkmdWCv4eyRECOrcNwGDtcDuVtI1XY7DlvRt6sLdYxLCen
1HxQC5kidJq5mAiCv0lbsQejJ4DEEIq3VMVqgQ3NnTw1h2eRsiN6osFt0bY36TBc
RdzY4P+R3w0DZDINPlqsgvPyl0nU8Gj0sMwWhDtS5cHWCdQuBhKD5kDRIX9GWHdY
6KSunPXXk6Ak3XyUS4HnQwtmK+wwI2HGNgnZamDomoE6nOvxDP1GLQ04/YkpTF59
62V0cVvR1IatEhysxOEYorfKhip1YbIa2GbpPZCLc3ONoHeChXmbzCByJIdpmBkU
BvcsEs8/kvAFcYOFtHK4pcorrfrta/+JyIsq5VEW2dKryU+gBHRpS0w5YQsrd6c6
HTvQSRN5Ih+cgN2KV8Qt6JOeBeE8M/OcOyNnL0l4miGjWocyaAVItbA0dmqtjYIj
DxsJ+HoOzbMq1oVgdG1eRpzTtYea+gIP8liJKQ7RlJ8P7n2zUZFqTuh793eyyny5
SDl7zSdBzYwmtzn3N3Enm7onxjoxbbZoi5vxnkb78AQTBLgXaQKEPxCrDwC4//Cs
7v65ZWNH9QuyWGzlvPAeUVt9Gnli7rNYnQI+aHlrBzWhjM7J4wlKR+sMt/Ti1ax1
5ns3aPh+s6ET6mMOO/z1Wr6goGuxmsQ49WhAd+AU6zAfJq3M3mk36n1CiVwho4tc
Lyg3kzx/FuNARx7LVdWBIKgh6ZNzQn3RDtGWzicfwMlAQMUn2BvZyej2Q9vO1DxC
u5qeHsSJdDPeEEQRbqsxiQfmQrhIh9riOYVD33zwLjsteuahoepv/wtJnVISb4b4
GJ1ZaPC7OSUB+dWnbAYFJZ2ecGZrc6co2yZLiTVkJrweOBnOvH9PvlCc6bP8eYzH
3YmSuNfGd+vfticixAgEULtcksgesgLrD46fFvTKEY8l/j7N9+N50MmuVBftus8Q
0Qe7wR+60NdBOr697uS/LGA7T75kg7boRS2qDKJkGfNsvgsqyQLfYipXXJTyunxL
oywHxLebyBs1YaTr7RRLGm/wqBksuEegjIKFFHf50Vae+uzemb+u2RTuAjsF92x0
6w3abMYhNjHKKVyciPW3iVVURX73x54yTfnSHch93JN12XaOlHmaon3eFkw1Fn2t
pKn2IhT+W1i1bEL6GTXmDrQmEnMjtGcP4yv4+nkDtZdaeRtOEM4fASwDDIHrpiNy
vYJq9mrd5xGp3IuB5ku9bhvwEOlEvEkXxOMYa1KCXCw/jNbT6VsNxA6xlNu6uAuZ
VOSWTVitjLLIOO7ZkfWn7vKt6jIFIlN5YotdAIn6KBWvGbe83OuQa+Ldp9KZacC+
949Tjgk/i7W8k7h74u7BxU8spHNNh2OfdKf8P5RSmCXR+0Z282FZWIrWkaj8jCzP
MCyM3NGMtL94oydQc+ZrrXFMC6LJQ0bVnZw5YHzmQ+nRHzBPz+ddUcib6q5I9MWf
cRP+Q6C+u6s7YQcWX8kNAWhPF6fugcbnFGpgClgJ8o3iZmQx3ME/VHn5gb5vKI1X
7LxoDcIdyhYeM2Jjggn8HatEpds9FK/D4eh/+g7qvoxv5kiT2GIQsk3QNSYj/dtd
oN467Id08weVpI/nzAmxsp27NTONHsK8xnSLKopkeOs7wtZ3oWbAhDOTgfQx3uQu
bsqsOKIUpmJiESIAUt5i/cq9g+4986OzbYVwCrzC10zceEZuCxklKJ3KyYjN2wZD
7QX1buheKXiCe0A70imp1I50fHsyP4WLABzD/ZFRGPbmDYo3A1PevUQrfVaEcKPs
xvXpbvgOCOqdSWGETCzZfR1XYFQ9HVbYvmOGNHxrWpGEi5cdwDk2oGFye4KU1rZK
bP1w8c0t0bkCqKnulUlnlr8KR9D+GCMdkiWgm5RIhkbmL9D2eaK4Agizcq6Gg0XI
dWd0pB/IX4dBljOzR3v+pwgh1Gg5oAb9/wu9w6QekX+3TNylDMN1Tp5ly6tIbMfi
9gahQ2+XJOPHTcCwhB9F2WAj5wd3mph/GUmA7S5dI7/mzoJ8WVh6JqImcgz1P+dI
bu7GFI+N/VpRO3gsz+4x7LgNIVUtN7/oLPVcWVwFivlZX37fUtKXrp5rYc5piTKO
D4KLQ0nKbevapeybAzidL/kqZ87Um90cfsrQZvmZ25rC0fAxsBd50hr3HWfO2LiO
5zzIwq7tkk5fwfDnsuhHKWsdzzCEE+emq1+WUHzlW1svzg8RpM4oSwL5XjzewWBw
KjC6fUykP1wv5AI2pJFNL9E4Q0C0tgoT8yGD8DQrS+dw3Ho4+nCoVRa8fileaJeW
9MFMIIYYBZuWB8jyza/gCpPd5Kil8YmgE9LQ2HY+6apdyhWM3Aq6nPi6qU0mmPbg
SEzTG3QiEJIQOYZz3xpJ5mWBRFRIRECnLoLmBbYwdKu/okFBumjKjob1G5LLhqy9
UaGpkmewMgeF/kKpI6atm2VzCTZXnxmpIxkV0Ggf+T4C1GyiGjBwv5nmt0qegHim
k0oYOiika00gjavtKlIsVH6Zro++DCNlrGRejeZKFwMn02lcUB8K5HKsf7sp7/06
qOZQ+PtglMrpQNvxryNS94pxk3glddcCxIdmuLA4gSC/xJOXO5z7yYDam4x9O9QM
tRUpkiCeoNVrNu0DWY0eslE+gUTUvjnTNjwJCuW6e7QEtFhzKAtUkjBvaj1sT/Cd
u0mWeslTY0+PfsU/smGaLzXgt7Eu772s1LqsSIIego4JvhKGXgb97/IO/ShAzbiW
0/cMWckFv0SJCxfLXzY36y5IHA0Ba2lVaq5kQybn6/NgHm7xPL6xz7T203ud556j
bVg0ybjHXQHIYGapPMUjNOOIGH66Zh6JC7Cuoa+Gjszz2rL9Wi5fSVecaFEv6g8w
tMlGUU4wj73TCiMFb9mjSeFLAQwXby+v3xmmfyJUzeXV2SMy4Kwez5wDos4Oh4rx
FBLEO6iDjGNfiaE6XDHHa4JTeNyxmXyLggssYKHy3eR1r2KHJ098r/rhVogGkwpN
CMHvTkMF48UDPTsjdUBTDKh6+QydyCZ9ksEna/twf23a6J9xkzvL5kC2MXxcBsIY
pV5du7A9eJ2VU27zVzecWOCnHGh9hSE1eKf0FQ3ofd0TBF1zsYKMqJaSqyH5v4s4
PiNLE0eZfPhLqQWiY86znSAzlmUAPBDI1oB1xDiW24KKLI5xAQXSP0PykJmvLv9P
RAggKCZ0R60S8WrWo63+8jQihTHpDVFLn/uYo5dVt6kpSnq85QgpeTB0wo7sjYLJ
SEonLGc2OcPUhbFXb9xGQ+pWKHqAeLe0auSDt+t9T4B2YNuAeUMn4bO7HZWEAcTL
IkJsT8EyDMvXPY/Nr8isR8s79z94K8saFnZ7F4npTtR6SipANXpID/Hp8B3fwNwY
dT8e2BOlESYVejytybVvlONzkvDbOKgkxVw0B2L42n0r1w0lTk/i0t5wcW+0ZBoL
EVXvAzefGcxMbzZzwkWgQ/fWjgTD/6ZjnK2j5PvflVREDRXfQkl8CNhpHbTOKAe8
csBZSbgD6gvSA/Jrmr6AJLDpVV39Ea8u5BqL3h1zkt72B0UCzOQrvMwn5LWT8PIg
2pYz9gytkCfIAc68VXwNViGGef5eipP6jckcWZrnHnAzn+uFsKQOBxTerXYp9BW8
9PiFd+rlAB3Vn6Pp9yuMlACXjCnZAnFmyR+Pn9D2axK1RdfjwwyOSB8ReFKsSttr
/ysou2yZxWf359m2qKoG9wU75CtXDErxhK5d1pXUCHKoRgGURFK2hnqg1f3LTm1d
DNu9I8tTNL89JnW1UdWVT6dn1ZdOLYWCdow7D1KLjUBgj0/m41k11I2p3snMLniP
/BVxGEohrm+BzIAIhFUwWKRcKRs+MUomWc6ShNofffi7vYoyeBJgPh5AVpMXYc2C
LeYnSKNJLgmv+Jthc9je+YJJNBztQi8XeulnEA6D6YFremma/cnSCKS07IY/Utwo
7RmIRxZPSD4fTM5Fn0IqazHAcN11FcdTwNITyJm0R7lxHIWiidTu7cpC0+GeTlHK
BKnaKX1ShR6mFPkMx/I4kADfZqNw+PptiebY5anKxjESgCgHkS04MWZNHyn4tB1L
9UQP5pQ6e8dIhpT0/HSlP2t6410+idHEo1cH0V8KOuwsRBbZPMSW6fpaIHiHe1Zt
upZ6c4WPAmUgv4eU1BqOGtgriDbiFCyFSBc9rqDBjWtJM5S+XY7L6OObdqNvWbn5
LCa8OzPLew4IAhg7QRKfylet1i9egZ0aZKUardbX7tt6RszWwuE2P+cvBJ2h5H9R
FXrRD2ZUTT0uM3lo5fVF8s/2rEqJNoT95Tj3DCEVaIHM9Ny4UjvdMd0JP6+Fiwxh
c88zehRCDD7c5wxHXYKoc2N3tqvxbw8mxIRO4IuB7GNOdTY5g28f9sLjxjUBsivA
tlEOlDllc+0YGTo30tGt7Ra47dUVay5J08oM6+NEYvJSERqSKVKK63sxNE0VBONt
JDnxQojIdS49IdNPwnTStu3FIQkfEwz9qeXkb0M0To1M2GeH4XkO5WEksCzvtym1
mymu3fi854W0tpV8k2+g/oJuo5GsedBSv+hTevtXQamL/NIxUfkxlOr7dnxAn+gf
oJs6CxHbbUxFa+iZNCjyOFzjYEiYQaG09GizX3uaBqiBEqCVbe4hSaqzc3tOeO6B
PE0fE2ffGcrJVjaZgiUPWHNJvoeu+03GsKfLBgaHo6s9kjYcJke8JXQWK+VwZ5IV
Ddj1nf9a+uaHdEVd9AP5Z/RWajSp+8lPUb1g3u1MD1seleLbK4sDl/XS9btSFs7m
GkzMTYUMxQruiCwHHEPdoit/ncz6f09AhfUZq9MYTg9YlCzZNINk9+rX3LKt6TMy
Y1UBeH3b6kdEmtABdG/hr0YJZZxgu/4d2CMxzSfzb1+jyyeUuhW8J/IBoeTuxSTe
C2zIDdKSfxQxWv6XtpCbOvp9fbITb2simYFsFmWamIHKCDAVeQqLMKmoMHZK53Py
iaz5NxRNcuYwfsaXp+0XhoNwA25Yx/H7HpPzdvgCBkhTydB+glsjqovzRI5u+Rbp
IuLD9JH+OV8CLRFPoNUBPIb33iN5wgCLP9qibcMEgK4pY2P5/zczmLAH4IeYDmJv
ZE0l1vuGCVsbRBU261KpJCE00NumDsgmpGEF/LZ+F3ctAJGfxdUSEIEyNDDKTyv6
NUzcwVOrTjxI9Fk7Jjl4FkPJQQKoypTxxERygPaI2O0mZVS/lHJXP1xoG7/2CWnv
tsm6tceB2ZjEdo1wfeUNXRBN3MvrsgIvwVshYUnG7G0=
`pragma protect end_protected
