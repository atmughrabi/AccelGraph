// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
atfmrquM0hShuXZeQH81bqCWovjuKPjTzeGuqjnuZs9Rs/hY6/QdaO/EwnVbXGf0
D13NOk9h8MvLR86DPWyKLRtM5sX+e7izmDwWHj1MnhoPc+TCBumgpyG39za69YZD
+P9EgktLdqEb52ZBk/gFD4apWFu2dXz9soPpIdByGHc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28176)
mMGMBdBIDRHz6RcHtNdZMJ69k6Wd6Zhm7riXjNu57kf4h78g+9/lvTxaSmZGRTj/
guSTp6t7JrtsYAhaZaVSq9sxrf2DIBEGO/l+d4rVTTiWJtfMSGWP0iiN99vDD0zE
6FfSaEV6tbOUu+hP4phqW13fHYUufdtk5MdXaQDwAVzhmF7ySvg2kFXE6CRfFwCI
rScECGnn481pxNuY8PnBy+RF5+4MQgUZfe+qESPQc3G6E1XYpZaFS3SqJPQDoURf
fnJEHGaLWwMxjSOUb8KvM6kNQ7vwTQd70Yyp85qslCkxcgznZaHAc+aomhgwTNr3
/J+INZj40ZHh0V0WYi1teWbgTp03GRm8Tg3AsrYRr0l1Lt1FZlfDac0e8iSydXQu
WP6eMo7HlQa3gOpy9vWTK3gk5TL0nZY5hDq5e6TToxx3RvvtwIR5wbBHzxHSN5Vi
3XY+xzKnkHovIapwrwgrQcpBCmuHgnPw598XSoSJskjtIjOWMl/8rYe2rpIuoMTs
JabHZ+vZIC2dj3QzdSKy8cTeKD/U33zf7+97hWeEnsYDpwKjiDXDQa9aDS1Y9gLT
hoVULk6RxvL2RHwYA7QoBudNvZA/jNPtZsCnSRogcqRwTUEd2pUa6QTBP23QQqsY
Rf2tNN/8S78Mgnz5ntjgpHOg3HMTIQlkoN7W1chJICFIln93Y7E/RaWCJpK5rg9P
GUWpuYo/ms4UY8QBGgZrA8J3pY7qNJviYLd6rOLM3VVC6xKeC//8gfTql4fRR0uP
UzI8qiyW/55w2mV2A6JRP3iqi1aMScAUM+moZagWSpqWmBELS7u/Y6mCN28fVZA6
sjDnyyWkuLK9f8QnThYD/8dgtbAQCQcyDWPy0fD57k+FfcdbLgiKHAtXRk94+6+v
Yv976bazgi8dEJkOGiJIZxeBHODL5oJ08ln4k8fRGQuj379JNLmIWki7mEp8pOf5
8PP5ow57psHtZJxvRNyL7R9s3FQspMKTqtMM3m9wjqMBQrrMdATzXb8Es239XOdH
Lq+fCluXNsRll7GfGg4wGJhTgHc3nbGtt8PjCSOfCS/bJwVpmpDGnXdBNgfVrG/h
LFXkhZGZHkHxIMMI1NY4dd0V/sRj6/5w+VoDfjAsuf5FOULsSh6kk/1ffE5nEiIn
cN6kfhobGEg4uS3JcCrK3CA15vjJwxbBv9OJlSrfcf0EoxicdV9DRYKrqVtb/vnV
iXiQ7IbSbZIlDKt2lXV6pPT0B2G7nN+KaOwIG8KA8P9A8Nz5K4XG3EXaihaum6yy
hikqCnzulqcrsg7cGK2oqG3YMMtnGE8h9wrg7o8hX0/weAB7eDjP5mcn7BNVHT0P
wtGpdZ49afLc3Ee9ekg9TiwZsX0Te+61ohod0rSpa+YuPD2e3hVWjWudWc4ZlKWR
cjk7AEdMUa/i+AFSFE7kI4AKlvv7uFEOX8dcJLbRkFnW1YvIw0NxY35NNXOSnLx5
hnWPpPNuegj2LIdshxOfOKsZ1KR3q3ynQNkdy6oHKHU9l6xxnq8M6rYtxm0Q+rZp
V3Y9yOvLrDZ/wKz4m86oG0xS+TH92gDcFzqqevlnhG+fZD/Y7oaPbhhticu7vwJM
oWvXPpcsSMx5mNjEW52jjmNABlahGAnGcHgjEWkMjWk4TXrT2Tg5/Yi1vL455PAI
0hKdoH7pxX6fWm5DiIw4hUugxiqQJsxu+ILppvpeyvhztD/UJqWyc7JJJYukkTAD
SJ2LoaT4qhaNn6AbhR7v9VVvl7BP5Bl3P92isZJ8cEUZ0ktP3k+22K4fDDpS8ASL
KUZI57lmhkTTZYiTULbSYeMlScnHI2KFWho2oFsNVHWf+DoNlE75IEIFD/k1hW45
KucE9LUE2zgDs3GmlrlcdaCNZbPcrPwrT4oaK2SYG7Be+82798ff3T5GnHX/TOLl
f0hwCJPd63zZQN0SNlhfqv2X6DwmDEurMIqKwefPasvsxDUnvbSr5Pt2Cq6qGnd6
yKo2rl07y8JC/HYxw2OdodKOV4hQ+UfPHBDwBacRicbWwUyDTyA6yMlE44W9lwJk
OkK5f76b5rKrHBYFmMi0trpCNL4bbYHyuju2a1JCGxXitPprago/SaKSe91OZ+xs
2TvqYfiPsL0sv8Fktj4OUiRNsNeaGI4J9TS7vwL87Ok06M1qLvr4YPXphlB7eerE
y3U/KKZ7t/4Y/yCnb4DFDV2vc59VzDYGRmMagsItEQsMpvYPNknNJAVrDgUa1jad
KgI4ex8/oij+gc4dOjpUFXulGLVdkw3Jq1lS0QrFUjQ5om1tLtuSLF7dnVxin66c
+FRr5L/tdKp6AGovRkWg6PXURcO15aahOS7qrczuBukfeBsT3+zQtR8g9zD+U1yq
K9mu9ZJAH5I/c3gxyn8KYL0vtPWqMb9dSm3qi6dorHjhQl3LQHU2uG7Pru7M495/
kOpB/72Q6hhZLOd6jJXewhpKETeV7GsOrXZn0ynYUzrM5icHzNJorMbR2Koelal6
AMK59ZhA6gnQ+Nu8fyqkCS6r2J6SDz1ejwwSuIhKp3bAJeImv9kJgYI4hnI0w4ID
7QAMa3rJeRmY6bVYYvnK0FlTK1ggcr2SKzv6jxdQhvTK1hiNuzL08NGqLatswLtR
k7D1+Rrx+bt6QvhE6yrit1+sOv8XtmVw164cW68qZxWfUb3r8V9T1Cqio/ShgENH
BRjLXehVpRsobkzQHl9tlhJaRm55tG2X6B+8hf9b336V7pDU4JqknlVu9s8LxtRo
oGM7DoMSb2Z+S+TTYtFTNxf5L58s6bp61JC7yc365kQAkBHgPxIJb+O9kek/qMJE
u2FBaiuBnnv1kAyfXf/Zq3idsfWEOCDjKas/JuNfGo62MARkuvKd28tj+D5vjozX
6TJs12M7XPdU9yCuDGY99rZdi5w7iXvU3pLxbQYYb74HMQ5TmwO4VRobtwO5jNvP
sP1CmJylNNLX7uVbSOGjOe2YMjNa3hX4CAwPL0+6UcLfy0EZA+tzAtwYZUtPcJVk
fq5nwsXEATQlCQ5lV1OdWS4d4PDR2fcFZ396CTvCwUUto7X6g0RHVo4BrlVuL3HT
lkPUA3TEXgyYpMIua36bT5ysJ5xu4mInb633ANLoa0DL6GFvsy4vIfylyKN2DO9X
Q7icqpQma8hwueiICEZy6yE6vRQjUcTGNkWautWo2qCmsOKidpUEvphCSV08c0ra
MVZ5uvDpRFRq9lcNEq3xPWIJnfQ2T9QvA1qKsJJKCYZ8GBHvG48VrNuGLdn4NJ/f
pxVSA7UsaBs7QwqZHknHfizIqb68fjPBU+GNl/qxWbE7MOiBXH21rhmzq3/jTgjr
A5nv8gqaTYuLpC9o7vLaZi6nP9ODIymqmsWNaiRqy6qh0tNfZVpJXQlyMHSdAeE4
nMZ/aL8tPrvEI8s+z3aIY+RXj1xoxrLJdHjItLSrzv1eTDGLIU5A0kYsqbOJmi7V
oVE0azG5H8IF+Iug8QqEdSxGUVX1vCO5k97ngK+BkgyvJrrxNi1vpDQnkqO3L3Rq
aJ3TngwR2FCh90eaRwb4svjBNtIjLQuBvinu9Mn6SReh+EWkpMOs72As2aMD65uz
rfWg7S7y55NCkvHcYlo59WnenMQy97v8qysnzpEYhjv23f557heT0ZyMFMV7ZCLf
xwKgAcfoLhSoR6Eym+53736msqmlXhtwkN9kmQrTBInEnfPYCTR6VCpPARhoFVir
WO3ZondL+N5his3/VqUo0AAOyi8ADQ0HkAJ6hyOEjh+gkSMDVPsTYR6PqDcICdPZ
Pq6YaSbUPi1cOTFoPIVDlTrkiztlK9CAb9mVvQV0Tm1dJJ35yx2U3nmjbT1eCbyZ
Xnt/s1hNZiTf18ZNpZyRoqq9G5lBzm4voHpVWj1cTIAO4z9r0sPNz7u5WfuBjlsD
zqHixmBC/ncGcd1KeT+/T2Gh93C9f2mH4KNCHhxBO25kaIiOJJ7lqpv/p5qO353L
/K/y5uF1KrikaYl4iea1fngjL8aaFN26OpPwzTvUTFbMZl7GBrheUutsWUpw0dok
KS2Gu31XWDt+lL3w9G0RBoUvMLsDSXS3Xh3iS8EbEdaKM8LSp+z0iEivLWtGQb6J
9gbAMfA3j5P6jw+utLBgGchoBncQhebHaEWl1KPbqzTPIFoaG8g2adUsjhKOK+67
JyavLM9Il7N4ADS+VNC5wi6la8dLDzkvfGWN1UVtbB8WTHyFLmS1EkI8CBGuuBr2
hx0Xhz2LdJhfhneR+ebj98UJdyK8PleKlk4vuCoyivYVMGfObgknOdkRUDM4uL9c
Jv9zFRqIUGwpuoI/lC4NqJmS7hKgJb6RD+lVipHziZvkifRFHS+AGQEa1WWa+tiT
7ioMo9eOZ2x+UoyF5glAz13TOL2X/t0qf+/+Fp7lPSScF8P1amFl3tjeic6d1Ctw
mBv2M+hNU1bYeSLWu9qO001PXECIgBFtF6DH091MnoKdXKIo3zbqc197sMlvoTGs
/D/eweBIDIT2Z3Y132RrYGGUMaWiywa9I0LnUGozcOL78V27IJpyF+yzi8NyAfyn
d11X00Z9jTX3uuUV1McmWN7efTZEaJvZ/uFSyurF3v3OdI9geiclSevQItCQ+dv5
MiCF9l+LSM6/DQ0vn8odZhUEFZWOBDdn01LpaIXS0IN8t6foEsMj2LHKISUuz44F
iB8pOq7AhBzV0JXCacLk0qZWgtpxTwSgl0UR54rfqj2pL1RiXxL4nhBOALQfMKQZ
NR7OE3p8/AR05a3+DiIirrNMBVCHO0MCS1dedWmMSzPMtWL2EjfTwvEPOa+EyLzL
f5n9/dr9k3d2ScCvoE8Ua5u04UCtP8HL37IwlCE4OOMtFGxiUtAVh4nkxSoo1Gjn
32hgZe+HEtm+ECdIu57/SzDk98cSb7HVFCu20PMlc5a/lCOwWduoYf84F0B0qvc9
r6VbDlAr8P8VVQUJiMlWuAzeLT0B7qldZs/Xc4oxqIGAdP/fsYVcDL52Vxl4M9IJ
P46xzyqE+Gfd14pt4zJ78T8QlHZT4UhiDGuR24wtWz16vyiIF4NSXbyTpKFr6J4j
0MrIiHh6Lhlp+R+iUY0j06iQaqTZlE2TgXdheGHj0WT/D+XQ3lLGbAHiapJ1XK9m
zq2t2S5ol/4fyg4n2gLtRCEASBX980K3FTJiGdL0GGApfj/8KGbWGP4zhTU3LvqB
U7imC/gnVQIQsqiaEVCsHP/5eYgTWRL8WZQvlOvKD6QwLBkrrmaNTrP/GZlFIorV
/nJ1oFL1bayzqVfqueR9y4MoMILq+ALK8m7y7lr9ZdpdiRdcBtWA+l6M3Q+M/6a1
MzMQu5vfqCQwC67VLWtC3q3Xt2ycDU9WsBqWm124RWVHl2Mfi8IdrvQTXWWJx5OI
4QN6nQ/g81PhAsBrw0v1JOiKxk1ijbL/w6mt4OggVPlWPxGhwh+lHFkcM18PzOG0
w5vA/FtxaQ/1eHut0EII7TvniGhrtReahyor9Q+xET9ycHBaDEm4NMyPnZwzIZXQ
0udm4t2E8GOKODNU3aH47ced4+Mnm8c91LpaTh89zLZROMve0WKyBFVXrAUcSWwZ
dmJI1VOlvpBVRUD3Xj/MJKMLLDFqGNcMf6VqWQioapxd+EQPfPo8zOLdrXAdzfIf
q6yUiOZgVKTYkIx0HRQoN7CwGoV15JLHGk88WXXqM7e5dee/3oy21tocxMO6yezp
BRQfsoYyNUFv9oZuC6o2NQPlDxGXFq5ArW1tFkpFoOAy4O4BHxQsQUtCs2WAwSj0
ER3DagpfuvgM+0S313KH8vHb2QGdrP6MxogVZfkN3mPWtcb0wvxdszVXbIUVanpG
73e7yrsRAtTB2BejAspw+40s8cPndl42GcCXiGlMIJQUjhxB6jh2bLD73tf+Vel0
SdT1EMvSOPgfG9HeOKdHQICTdL1ACbPYMwsFjF4v4HoIpkm2yE5LvgqpPJjpJCOY
DCyObm3FrIRWc2mQt1Qid4shyF7pfnD9Yq6KG0SQqPt0zMcSY6ds1A5MRNmqveiF
cnGe5KO1f807BTGAMHedHnGKJdBV5j2aq0ctCuc0NwOqrlwKfe5l3/NVbfxhWMtU
UtCgiRfvi2b8Oryc+QVOvjgw/x1fOG2lsvzWoOdHO4zQ9/Cc9uBUgSFkutAZ/TAM
EjCSJ8M7dYCtqYy5Vm/r+/lhxgu/FzZRCwpU0roDWwWVvOqITU1HScQqZHmUKGnT
Wl/TKeX9/caB6duXq69oJCPnu/fHauRWdcNRr7BmqCmgvDUXMyIBobA9nGvoNe+n
3HSpcZBHNer7gIIIquumug1+tJo4FbsODH6Rnm5V0mM1752+Ky8r0laYm6wJrWjU
W4HRx/KJrOTCTxKLHv8zEmxGxvGzzpl5QGiNwzS+0d4hp/lP3u27vpfLdLF4+qxe
u3X815dA5SgcVgJO0RsVwAt69eEzUvb56qx5gfdgLVswtMLilgnP7iaBeesgzNCC
f29l72eMqarZ3pjnMXV3iRcXlqIQDCbiwWVMv1lylTkFg+Qx6z5hYmo4RNMCMO9v
NwEZHnkBeFmcDjhxBELM+ZEDTexk+wwEvkGndOEbv9tSGZRRqvEBzChO0M0d0ot/
4vy1U2JY10Oiovqw70DAbuPi5Rn4nwfkgis1yRzsKcXa6KF+quVEzc26M1nY2N+u
peawNPIKyXGlsD7d6z6Au+eJm4sie4h7V/LdVEcSmVDW4fFu41D6xmUC8CLfgTpu
9A5CHmb0jwXTAGljAvSuvtoLtshYJkHiOHyTwWeakzzVdYgVx7b33oQ3bZmfIlGc
E6SO5HUVpL2wC3KT6FSUEEAtYVeXrNxOVDJa1vqkaR5/kOpxK9L7XH/YBZ/I8mOU
s/SFxBOUAWdzXwIku8HKEjIkx8EY2LDoLvq6GCVyZVgdlmwc7ITHhh5gga9mtVvr
6TA3Rm1LUfp6pKWlUcPyArmkOOPakaermjNZ01rnxq1u3rFyZmNzPfRupuIlBTzV
umcD1wCpWpmzuaIev9uJClrxF6XBUDWTT458Hkv+dtan7nmL6UZPTI2BBhrOfIIV
lUl7k50dOc7gn6jhigzghU5v0eyjJNKnLIcNKFBa8KsB46bC0DI2O2KHk1qb8qdE
rDzVy7GSupJ5Ytc1H3v1kFgf0DqTW37JKPuA7o9iJuu7HnCliGGHEIGiNfB8/1Aa
RzuGUT54gO6SP5TdPrU3PqrDTYxmouU73gFSkzopB4xh7Qt1Rz/seErQzQVZBO9s
8901Rh1/xnCq3i4c73UplQNm48rtffH/nSvXLmH+NBngDkqkyDDmdV/gEOIRaD4T
F64krm8cgatYT907OUkPkuoOI7PZeFJlO/Kle46X2w5GkV5fNl9VPXk3VUlKiayB
t0GLc5xy5HEWuDAzfIDLDevLDvRFZ9/mOjRJ/B2K9b4oBpIIkzPFLrcDJAKHhK2L
mFTTLB/wfpbYSfQato9T8fLv1sRNyQ38+cBEZP57IBJnz5xXHpA6yeqUba9x/UPh
OgRdZsX3WF5RKoDkrn9dpbA3cHJ+PJsrMftaV45bkaQatTKRQs3XlXvGi0fA6rNA
+4Cg4fzDCDLB3F7nX3lzvM/fV/8iCIgYMB7PdvxNqEm9Fo8/7WRkUsUmxiaxyFqM
jFGF+DzCp9E8pWQg1Br7WXiP/WcO8RcLp6xBsIrOfaXQxvgLoP5PvieOTM6EPVsy
nRJRiQ0+IvqQF1aiiAtSkJ962/B14j9Xyl3TbjcYz+AKsExOuRP3gP5kgWy8Jnxq
SwForWsNrFuza1zcZMAb3YQk4INbv/+B/Kdy/o0uZWWs38JvrWIQLU7sg3JED8IR
bQcriY5hdk0p69mD7H4LObow1fqHOlcYSeOc7iwnNXtSKedecKjM2xEK3k1bC+gu
m49oPi8QOetcRdLLZucMKg73I2vG/0/ItrFLD/NDSpBTh68e/8T08lmcv5KIOlZr
B6obhyJK6+1/jih0F6wOq6Cul4J2zBDAYraV0RbX4z5EGo1mLQIK4N66C9dIVU/V
3LrV/eawlLfYbd0012ft/XpNF4+V1BJvcizcTEXnKWgotbXqm7T160soJeGr1gtd
+l53GfonddEpS6LUM6eH3x4y7mHYhRqwhchDVuwizCE1JD0+LB+LWft9grrAjY7F
hlEVlY7gKmobBRE5t8DzAPezsTXmt+6ElwR4lDPebgoSP5H/jOC9NF4DRn+DTHBy
yrEJUtp2MCI8/ctxF4FtBuzgySkYSlGz+G5Ogpf13Bjy08KrVuW6Q3p1G7N9lpXN
gGOaReN1DpGha7pIe7cUJNBPAXYryPcs31bs4umMCgBv+6l8FiCnCBitl1F6w9nj
S9KitYfJMMG5UYCEbgHZf6guNoG6whUydbQdCPLSOvDHUqKWhHj6lk8a0DvJHY/Y
fV9U++K9bVyaVuIKR0m+HYU+uZflQtc51ZooleS19OPuZFDipzCwfe92p/HQ2B7L
H3GK5/Po4nw3jPICM3UTcq+z899R6BUUYMF6EUgw6j0KwJZlh7SEOSU6im4/TpU6
aEx5JK8ib5NC4MSOLqNxyCwNPhZduRx1w7jsWSdcaoJuK7+8CtPJ+aCLQyOKUPRq
XnF23VfVEFSJs/Kf0Z2uccBVjmFfQUDICMjLQvxP8De1LuyRq9SZEDQJnAdtjJhg
DqlKNjbd5G5s1qszzHWjimrm0xJrmGIdEIele4R+p2J1YAQnTrY7d173e+5UzklB
vZ5RrvZRtWf3ndnExZcvtxF/DkqveGA4jW0OviRBovVIQirlBxFgfeUw26sZUFX9
HM+yJgDVQNYMrS3Gp85bHDZAup31htlw8zlFRSVgs6hLHwGMogKyUnFLhAuekpkt
s55DLLKj8b6pVumYMus7JWuliQuB/P2rDGC2vrtvKr4fahFnbyy5z3KrhxtdiWIW
XbFy6VJ8zahBjDeUnoxNPoRTxBI60mDaz5WvOKSA+QtnRI7puPl04bxopmowCfk+
SInr02j/6Z3mdEzAsSbxb0vaNIggL1nvVohhejfFsde+Qzt7sh6r9xUc0dhrrp2q
lPKNDinEqS6OPk/mi8fP0VLo16eDplb6j/D0dVT664HVhCIzFB2LrO87/Q2LesGY
dFAP1NpmlkWgzl33mYq3m+afVY7sfw2HxQMKZqfFhq07Msbsc/0BzKClmGWzQvxV
cJPMFSTS/GXUwBdfvzDI8/Flh1bQ93k3XvNJQHsiVu6EXbxBL+DHEHAEPtct5f3u
aa4M66AuNtPaJAYtVNDyPoX16pmo8NpswQrkvMhY4yAwwjMCzPbMU02iwfFolht/
jIvehG4Q76MGxfrBVCQWW4ntLX0qNKno+Z9tJLgYkT7YwTv6FUiE5L3nNzmIA5Gi
TIOVlL1wk6eEuPbib+wQlw+lY7CK70iexWxQ8MCW29vTDXUT5MG3A2DYFkSNRRw/
nM9wvz+8QpquiGe0Xyf15GsE8Jpe8L8tKjFggrlhAGhaANeG5nLqdFZeFRpRU1Ug
Q3RYkZy7NaRRpwXpCXiaimcDSx8guzY058/0IADISBrE42Q0pvkhPsSXMFa1MJb4
94B1ECNVvJm2rLawiYkqHPQEehq1Dg2lXtPhUde/TLjZRzOa48K4vRuyWhJV/unQ
Cv08X5yZRjdPRM3W9j+2ff7fHg5eoOcXf9jDwf/nMPaNI8jpLsjN6B/PmaJDYnNZ
beP24RJf40Tfg08RoNy3PSDM1vcRtKZGJ/FZ2X577uIsJMEdiPCtOCto1pPZoWyE
XQwMRnBsFeUqLVP2dehcRNRt0RB/UZOSNC+yG4vGXlRFG22MMFby7wwr5zcDbbkz
29b+jToN9lCcp0mnmHL574x/tiHUlFTP2Q9J6A2cjVNxePhsqVTpfxfb1DFuwW5S
I/sEZsN5+iHkI3tVlZoVJ3R0kMSpvIEenhaiYcxpsw88RYczmUB73PxABfAI1fLy
+DNBbO20r3ICynLnPNP7dOqGHcYqgLHboqSs0PKCOoelLByGQ+BR+vb0095nEdMa
J744HjKwpgLZRyDgl3i9B4J2qeOLUEDLvPfN+pUJWn1q20mnUYQB0M7fjgkck3xq
1eCBCnWx5o0tiizDIzD6KFcZIjfcK8dn38f4orrnmCAGO4Z/cDK+xyGNCT44Kvg9
IAZGUK9OLbPvXW/StbefGoVm97scAPN+igQmfcBQeTIzTcAw0MMq0m0sa7mdtagr
YDuDqNql5qbdhUCs7RBSnHAwqbobYnzeNZEoG6Ccr8XRzAN3oYsUpWsc/JF2jifh
3FDpq5RkBQ0Gd+z0YvekDCMpxT/ULKue28QoKdhtcDShTNG753gpIaOrkdcTVfzW
hEltDhfoKvldNqmOCftZf9z5Ze5Hd5EZVkQWBlzDCiKW6A24heJiyGObiG2x2P0x
w+bwSWWjLuPRI+HUcOuDcE5I563fcs1nIGhiFBGGCDZjepbmvkDCTWK6C8kqoBSh
nu85JMKidxiG/lhd6T7RA4TKqM3F4JuWdMKke5gvPIKmOtrTgbl910mTksA2suIT
KgGsQptvYo091jAmWwtMAZjAGU4AqbmRd5kibCOMNHyB9ZQARwhghJtbo2+XeTUW
YQ7odkOPNYMgLjqS4iby9DTl/yrfuKurtHwFTv8exuPzn6IzJMWDSleqhLdah32t
klSxLMRQ3qh90QbM2WoopVC8cvnSzL9GD0F2nogt6iN9z+OamQl2wzUjQwJ0dLjg
pJIBrjvrYiP6KwSPuH2t1Uh1J2b8Ts+SfAV3fq7hGHuqKu4n2RNJO4D8EA5Bm/4x
dtzNwCCCoq2KDWMMl3T94WoZgh2sL5JAa2z+4HVpCSLQwpLwommarXMQA5pnnzpi
Ud5x+jFZS6HXpzU5PUcZMCjFuBR3B0o0/w5jQjeVVC9C7bqLXjYT4l/2CHgh9czw
7i4hr343ftPbG6AaXFJiIlQlPmTmzlVwr9r3ljQBXJLKCxSqGqnonMsjp7NlHbpC
fEh6J53KZCCXR7ZtBB6UIdfCh8/8gs7BAHcm6oi0A0rsVqB3BMyMFXb8hv52bvoa
T/HGWZTglA24fIv6keRjyuywEOPIldgfKNmstcr+7wlRumM8VDKcyQWp66HggeVE
gbr5pBVcaqND70sNcViF/wRS3QJLtCCKPJSblGZ0QSurHafkeHlb/6nmyCecSBre
eIcsT+tpg3cQlySX/CHeRXZN4Z7ycV8yg19uJj3X++8aKSp8pu+9CvzoSa/16VVg
YKihrwOZ/iSiBsUOo//PBN89nC4mzh8R9zreN6+uKwkWLnk+sfVML76NSggz3zRp
NFlmd0PxuCaQCAdTxUcahCq/PeJkBWovHpbYyTwAh39BH5ldE5vG3PNohZ37jd01
2kUQAqvyBKnNR2KOFt6oimozo8k6TOlp7eie6eeBKkQCWL8342uuThu5H0GpR4YV
9WPQaQQtyuvoRiKtQeoMXnaDGz6euM61abz9x1mE4LWHxBkgF7KssRSMzEx604K8
C/8k2xf5GlnOap2ZlRSeIQcDJA/GGm3mMIjKchbyLQXHlwDrDKXAXAp42sjWkW4p
wuDVRqT6xQhI53EIqGSBnWmgFGoAuCpa8cmb3I+/gHEzGWqHzzaXZL9gXvZIiA1W
0Ow+pCqCULnN8RquTwpoBtwZr/KDBbPL0xhlFqXBJeY2rbOG91RIILSazH3qLo1g
SsYhv4sU3434izNXlHyDWa02P5zWzhGQzJCkJS811LE2atEaYgetHW8RXRFN4d2k
B7B6lYZmwzvYDoz+GTWnJr1gjhLqB5+/4oEOmGbHopL+rOyHz7tC0QK9ny9tZSeG
VKJ8U43+oTuQxTmsHJTx5vS4/fymXyTdIx4PdTvn6aSJHHrwih3ak/XyXmlnBMEl
Vkl9YYfDlxoqrSjKMKHGy6r2we8hAgf7F2i1WrMW+QGftfA2JXKGiJ4guvfO/PwR
v/TuJoPfrMVmh/WSzoW0Icn3+15rY7spenNfeMrshXGszG212iSe2rTP22gkQU+7
H4f87+eTTdbTXUOSakojIzIx/dQ2KkyVa7h8JyKTxQGw8W+K1nk1wnsM7Z9GZZsd
6rysiTAAZDtFzIc6WA3ohMruwj8RGriVYrhIeMMwLIxfHqWuxH2cSLkqhH7jm9ry
sDVgGD6BKPV9EgO/C0+/A6IoAcJtX6+N4AgHUNT4xqWYn2rslQGgCyIzzN7nPPYf
9zcWiHxpZdRMhsq8rzgk1TjJcFrFp4BeTbUfGH6ovMA9RU0vJTIyJMNwDNQMWxok
sKn3MrqamjFvYoyROuPGuckcflzlB9Txpr5/4O8KZ4lE0Mw9aofDEihRoaKXikqn
HTAyo3kKRxL6l+aNZG9oItVmUxSNiSOyKCLxhL3eLXwFgzhD8to2iG6XqRQjtrAF
Njn8J5wemyqTa4axbKk6Ikc592k4imA+a4PxzGgQLc2qYkczCnTCURg4hkk3Slvo
qRyXLLiQPKPP8KEBk51mZvOkK9V20gblBC2fS1uPxLycgeBZTMlQV34H/gjTx3DR
gpZYWGYuEapNcc7VulwqvvZrI6TkOtu9v00JjucsEvZFr48sDG86mjEw6n2ZWMeX
S6MQshffuS6IRD1SfjuBVTdrzFXrHuqR+zFmwzCos9Y/fLS2S5Q991GW3n/tlbRt
Ahc90FntFK3QznytW8MPGmOj1wonCmFRLU0tG2ZnGQkva0wDgivMdzBWKGAidAbX
6E0qka6qg7xYw9DTyYzzvJAOp2RHi9He3WkbcYCdlYevOeTa3yOqp+Io2S+hYROI
LgE0HzWiVHwLViEGG/BSqjFgr8+Eu7mnsp44zIOotI4QJdxcP0oPUmqlhEpO18eG
gFUnUIxG54z3D9SFJyG2H2ZuN51MB/U6kjjfeTpHb+gNZH5kmqBESHG+D2EETvJ3
c3XA+Rz1poHC8SV6c937rg3UA7fw6BVgCXHpglr+qUwz72/vEOj8YOwN5OJUdWHw
fTtKderyZZwI66eRDuoTvIsmuZdt26T4S+hQU0e8ft56BC09kwvwBPmRp1yvD9TH
RlOWTKIK5Q9EN4i6pMS4KTkMDiX2PUUP4flPFK1gkEmf93qHeZCOy5rmh02uuSG6
nv4H8SnF4yxENnA738mPpJ+isChFchH5Nm73YXPs2eFJruHwgTOggr4WakW00bB6
PTY/isFB3OIV3suwu9dl/YeGaFPCOCWQJt9coeDPfWW6raCdLs9GAWz9iBWG+Ts2
3/dOwmgiQmib+Gfxns/fhvCgfeSVzsNRNYtz1SWEXtGzNTyGlKzeSL3Msv9FUQ9Q
KRhmDZZNlzIgpCcEcu+rRB7ogVgvN9AB10hkhgAYTO4O+P0JPt5h+bkCAuUzKf0r
myyT4juO2uN9pVGjAoS6/mPHjLSuOw47W/TFft+p/IsvchzapjLZEsFjoubhdsCl
r2gkxkbvSVTij1x1vUgEj9Phohd5/CLXGGIQ6tfkUhJffLBwGCI/08go71/sz5M4
4V9edGvReHMAy0QVDcdrR+Vx8o4xc8knMttN89G65pOMR6k1qoK6eLdm57mk6pLq
6FIyMcJFLE8TibihuHVNu3JPcyDGDKdTAzq+IunuyxRmEm/grYgie/bzCCX7IwYT
AaYnGluyRKPw/OweCGKUvO1KbdRkilQSCs4gIVtWaoBrr7ZFl6ceEvIz92oWczZe
dQpWRSoN1JkamTEU6BIq7jWVin5ZlxYCW/7fqEkh3UT+++w0P+DE5X2DNrZSyynF
y4MET1Y0GuKC6DH6pXH+ORxLWsV6BuZUmBSPAlteWJRU7UZ5hGOgfUN9XEqXeToT
CXtm4ZDcVHpJnjG6xDEEkTQd8thwV6kQAVw7ziUoW14CriH1TQ6yHNVPUozRTFO/
57sUmbzZV2yc673rHq2WAVSN8xwocq1C7VEGja8TRSVceFSgIlEmX8ax4ljKlYo3
76LHd6il1oUPWIgmz7E/VyUUuOg7C31RWSne8BEB8ku/jmNCb0YEj1708ZjWf+Yi
O86+oH+24IBvMQ3K7YCPxkE4a3iwMlYDQmrtTPCyUAEL3OsGpDP139SY8oLp1rYf
jLSI7esm6q8MD8YL5EcVnu1h3/T7aML27hDytKlNScE3Bec9tNfaqAcpTlVi1r63
ACAdbgWHd4tFKKkfFLa4fCExSSD04ZxTtUYjftLp3eAmNK1BG3gP1G5IM7MQf49/
7Ogxv9OWlr9zS9Ds/F92KD+/Sg6mAz02ZRGXYeSUZEZ+Ip8WzbxWyoXMn6aBcYqb
YJ1/VD+KIRV1pW8E8KwAIjc4mRYTRG8Bu/QKacQLD3QHoms7tp+3ohrVdIo3RBdH
CMW9iobRyNOi5Z/qVvpd/i22S0zZKLjpnoHsx8tMhCer26qw8i3ZbG6f/2HUwlQN
osXz7fuORN2Jx44VNtgo8maoEw9gISsuVf40CJHVfZEcCG0CUw3ZUJd/nDHcca16
wO/cSfP/6MB9HGrJMbVmh+PPssJW7aZzuiMqJD7cEJzDt9elfOwuL9fM6JmUiey5
2CplUnG04PtCLWgv2eM4e4mjzXkqwMFrwOV4r0sg5WpFdciHNmOKbSceX7BrxpUx
8xD+PVjzbjnjCP1+qkxgL8F2sQx5XaA00wgVLDEXjzQCzqzljNj377h5GXDish1C
ewV1lFi3RoKTXk/sCGbejCC97sGmtijenJx4jejHjKA4290qdX95kknIiGt7zb8U
oYbv5o39SEN4JqgR4cCowsRwEt8HPT5UqSjZ6SP5SCkKfnawhkbbzCM6C5NDql1v
3bhxC+qgWBkWrcZnOQILazo7rtOtbFzV170hy1yvpcA0qQEHS9ljbl3KdAPQNuxB
ysBfpJxq5DfpzV31P9DJKuCvb9FRxQRuSyOE9pUDa2xbzL/geEX+EbuqaqYtklZf
7A4FhoSRYy08BPKodHxb2KbHHLQY6J4fEzVAPW6iRuScdFT8KgsxNP6UfLi8phM3
gfesapxEG9Mw2WXgLlA6dJUktK/+3t9pS2jVWalwY6fPn8WlzBo3Px+vtGRB34vI
uECAmzhqTr8+4Y6f+pb0b5BtYqFwmllSO+2UdsCc7ZHnWGnTz6MT3p1udo6j54ve
1VEAw0HnS+DXTSfZT2F/9J7GrHyP3/hf2cbsm4tnAUxVLJvaGbfWOPbw0QBg4+U1
fU+7A6TZLnj58aGShleJeB6asogXVnw73JZqDJsmWtEa+/MdvN6VmlBxMyGVDToP
tgzttmEDXMe/jCSq3cvWQKurFzNHX8dizP166T2U4Pz9SJcc0PEnxHzpsFxHIaq7
hGWs4XRbegz78bCfYKkR4Nc9EQXNlkJCuZUerKqPImvfrU7Lv8cV87xnx/sncgDR
pJH9uIIAxfDMEADf7d9GJDru8BzM47BRJUxn1KHVebc3XzGqMFqCyS3B7Ld6jX4s
ZNdnvuxMWppEB16ILNPFbCzkCckn9pa5/a1Zf2zzX2vx7IiG4fPS4QDYRYXyTKm/
4FRz5cgZqMgzEaz35gd7v6YsIqWcyvao4SIJ9rhgL75OtzPDmiAy8mFLqCyqRPH3
KTHqdHZh302znjT7ttk8BdM8I5A/BW5Gi/RgBjbB8IWo82VNT44J3bauRKBJW0kd
T1wEquGZ40m2HFNCiBJvucIAsDP0SgazTf4Eq3p4S7HQVyZzqdNALy7Jt+O8DC2J
zwdIMZexu9//35PVUKitwdCGJW4ACNQKlB+oK49KWAhJEOwQqiXTRTzg/iOFTh+V
uw9KNbVvIyVHHF7vK3QeI3hv0hS0Mc8To1e1mwT1XwoLcVlsq+7P85P3PBIgPNpZ
Y8VjmKCfqEjIUpB4UtjqRE3fhvPGgdf60ViwXSHi5qdn3eDk9NFh6nQ8QUT+G0Kn
BLedGHRKTG9a/EJHuzxdoEHOpXMbkCke3k9ADAQ6QRVTiLXfy+Lu7k6puaWYJvOC
+oMRlVRvzS9rCFhMWdQOdt2sK4wek2ra05BcHlW4s1LfyRqLXoHkpMdjmcpkjKO/
PrZCDPqU9yVD72jX0KVFu+HdaYnG95kfkPfSdNpVe0Qu8dbz0oVfsjVw7YKmGlWR
schOKm01gvMkdlBxxGpZa3lXZ99INBuzHuvLglVsCushsPnOOcDrXFNppHXnEuWg
oja/mSGiQnTuBf0NkE6RMaPJclgnvwTZHRZuPsNIIrcl5kLHES5aeP7HLflYYTt9
ncR3BT5dvWD/wCvTb1+lXPgwGokCQ1MBcYtB2BF1BgEiVaFbcE0SLbFqO1l+ipJB
sZPFDtq2T3uvD0j5b/fg0AdPswSLz5CDzgbGo91MdcmOKgFGdyHApSGV71TaZit9
G/mPmjiC0EQ201o+jBTmc25Xvet8Ok0WONvH0ChoQx2BiSxvoGlqZrk00xHf4F2j
XNio8V2BrGOcthKw2bblGME4ZDWJUv0s3eIN2KM6U8Rvt9K38wcI27INCbnfK/Te
IObd0w/l0PRxTCbhQndz1jyskY3J4sXTHEjbwyZcT27lZePyhucCapIgkYAgm+6s
u7e/peJaddxwJVdLqqcCGAIpJL9TmJrsNQG7oo4ilbQEnIuUTBzDAYjI3UuRn6E8
ddsgQOAU/P8j1SNICVEhtqbmkS85vJc9aPoMfHW0qoOlopkuLTsP0PQrunz2AUQZ
htPhaoroFSkhzWb/XWu/NI3+9CQNi3sEa5yG9nvnkTf+I8YQLPvP4BQ3nTiz/OVD
wg54C4mbjbkHWM6z6Tydh43krHYnyBOOQKpBb3wwi8ESU3WWrSi9FYuuEfGAGTr4
AAtbj9Szz8YZrsr5AneiNydVJ1G0Xgyb3X3LfFtrGWGsWHlUA9fY0y14JqFFUXj3
fodp4thgY5SKxGP9up5e7JG9V25WUKBQOcXvAO8BTE6OGgHCAo78ojJCMaYBnvid
RPCBlOg40vO5Y9RYQrKFB5Gzo0Hg/U+vShfKh9s16j/YiRsCiuPMKe+zcLz+bPyV
bqzQN+T9hX1UqEqidaBaU7pEzL7l3rjqDjyf8VEbW0qBiV/Nu3Dq61y3ulgP7nWU
a3fHhMa+XureJ61qGnv7m8R8jwkD/c7WlhR12IeL0wuItcrRy1/L/F4g1d/T8gdE
d29lHe2yFVRlQl3MFMiWT8OETmgXs+H02XT0Yc2sYuVJAeSVWXtsmlzS78L7LuND
vuCL4u30wjtXqmMaNKIwG1oxNF8oTx6yqj1QaScS6evJ1C9QIWKlv1CbI7ej4XBM
AOINpn3a0YBvhe4+HxM3Xwbo9ACySuEq/f8LJI6RLiBB83SpquUyLj4JT/yTkcaR
YCPHC+46iN6hi5mrj4UAtulxLM8LVhcH6tNxeiFouF8Yjw0X+kkaiHrtDOIvEyZc
jNp+tYMlmBczkX7VTydT55rGIzUFdlrCjgkeD+IauISWMDRIQ2PbEPgUPdqkTD+4
ycb06/IFA4y5LQ4BfsmuUVXX2zhnLkKStj5s41ivNAhwDeBSyWDZ6vK3Roee+ayf
jctZjIBcRDWyoYm57llSI/Z7iuZZTNHqypH4tQvcGz/fEkkx3xLUAjxbRHGsvIBq
BoHJpsgLgdIA85XiVGfTK6N+zZeIr2+tgvn7CTCZG/F33P5+yFDerpW/rfZdtXH1
9JHl/ZpmT9IIYI4Fkckl9Z8eMDHWAckm04qovC8y9Up0tP2QTW5d95lBeClY7n+L
FM0e0LWlJ+n94yCPKOIFBL6P+dFjqJKuRL5Ly57sYh5I8xCT7qYxdJg/P6vZklNH
Dt94ZpbI/GSX1W8H0evYvG/oAEOAn/MviZNKdhQYZHV7EWeibNiiL7TNNokY1DQQ
0U7zRqhntwxUMqPx9qAJHN3h7iCTIsX6sMTxEDLyELkOSlOlz7CN52JUgw86A9YX
yGXCU3yergTypq3WF+4vUntj9/odvf4TUN7Xfh/wZ0Pw8A121wj+iash15xl0HvH
wqdJJBGYLiS4dXY7HtV3YI3dQ8Zlbv/jVChjOQe/eFF7sq+i5zbo7Cs18kb8zsFG
ysBxpmexUqcKMa1snZcdm+DEsFmGDPOdP1yWR5nA1EgECPl5aNpg/QraGAQwFqjD
T4s8+fjpEXwzJfUBrCKqhERnSnJAOi2dzps+hXms5bQcvu/qeUBSG7MQFSRLoSxW
h7Yx1aNWk34774epAeUeRPm1JkMPNZ2FBhQ8oWNdVYr10GmL7NbEwBjsksPoExHL
OVgOteupQmHSmFTV2Fg1tBJnysbJrEuaInRtJcaA58gyTAUobBBMkdbwFKm2yjaR
6KKNeAj0gmI5+zhSZ8eOHObT0xWIDtVxGcmikuzf/ergURWXTbXY3ojKHG618rxL
uT/q8zXSUySkAPtKA0taKytYoCyGKJ+HfI5tWsNe6JdRyW+K4Nzb/4Br3i0y92nc
BedVHsKplNWNnTxVAhVVks6BVsVBHJTWrc/Tu5xt8AjOLqwaHnEzZoqMPAf9lYGZ
vHJGe6YYN9wyNFi5M+x8DZ3RW+9357/Os8TLR36ESCVcrVlVh5NewwHuES3Y1hFJ
JLezA6cdOEOfFEuCnmGO+63h4fU7bdxp+3JIV0LrPaYJ5hTMQcMaJLb0x9Z4X/X/
2ffrhx7cyg0LqKVLt9J1lVZcYWKo5jDMSAmfC98sShE6ATRGpmuGRb+6d9W2MnGQ
QIcYomAVmM2NHCMrT5FZp1JZtRTWr+Q2lmaVRRVEq861kXm2odcxQpVqp9jtcVB5
dIWX8HQduyMuPrcqkyPJcEt01WhQgTy10EvDikxn/LNih3t0Ommd10DoRKHKkHqV
H+Dwn4Q0MBRK/bMsRTjAjhs2XD+luc1BoI3kYGxGrXDCa4gXxoDjudn/uoRVgeJR
zN8mT6Q+FwObYNQNkJWUWhTzSmK7eQhCgLM872ZW87thY1X4EnkBqsbPEbfeBpSr
25corFgtJ5BeSclS8Nk5haF0sjITjjhQHddq4m96B1EEsWVvcwRziTm92toYAt1t
sVmnMfX/mGOYVAlIT6FDslx0v3+8Ihr7eKurZQK2FfKVQ3HdG8qZDMyE3lOqXaqz
COV+O6POvzhc654qJvw8z2oGDzcKQY4SPdXxihAx3LLRlDehwXy7UQ5meaMmWAWb
GpVbZJhvVU+j7ZhraeNb1UVkzFY2DdUGw/DbKKcXJxSs9Fbz/yh11srsaF8FBDv2
XZilQdyqI/CVe1BJ1UL/PUzug0tiQZFDHw1PK0S7uqXh9bIPuAeQflGAVghbyV3C
/2plNUBnYUd6/Lp2dSiVO2r71upjew49X2Rf8X7mmry/cvbM+RRcIdtTo6f28jIS
zLOqVJxDaK/JEIRYNOwtgbuy8xOzf4/ZDMAMj0PVTa6WnbnvLasKJ0PSra3SKdMu
UnAJsBmBT3UkF5+OrNyZ95AcUMSPbPIBZwGESm90PSfwoNFdTKhj2iEYsDUQRjKl
3JKYqtBTyiL1WOHm4ZaySib3/SBt9ELxzyalJCS4zf6PujvwAh8J4q16F1e3lT+J
sto8DwRX0vYcWCcvlCvBFWSUP+90mMF/SPiPCXbV3HraXmcoTo4pdapvvTJROEpB
nSUPpNHws6zdaYRByHlcFpEWNUZ9dfjwZ3qiBu/PbMN0j6NuxHRSbjaRH7KC00b8
LnbfAUN422WLxk75RyyxpiVO3c5xOg5zTQ8wuOCG9Gtj4pL6C56UeloNO0mgRZXi
kzf7B4IwzecfpVhrkPJzVHjwig2CVH6Ejs7hSOGjK/4M01NmlYnIWTFbPTH0mDUh
pJv3HHmX14dKQRCMDBDgO37u8qH+hfaML9o+arTGgaZqdsMbw/ot3xr0+lT/Smom
ow0bgtHIZIq6Txps9T1vmCg4w92K1U/VWjsa1COFxv3JYUUKz/rgPmDLXIYi0NiD
jPHWl8gCq19O9goYbpiJwinHDwJaZoRHmicbonb1O6nu3Qc7f2Ssb3lLV9zDfgP7
akyQX/q5rgeur3NA5vu3NvLN01i/NBK83sg8eZ9PtLB2Rc9bSo17Gl6knZ1gzJ3F
DMfnWVvBXNBjwsAPF/WBgn1zRhDH3PDuXhh7Uzxdifet96zGmNAQV4FGnPj0Jryp
+ZanORwj0ZBc4WY0vbx9Z3ZBKzipLTyYrCozc1gmaDpxcP09Ws39IKd+DsWnJ8e2
A3iIRZOzGkDR8SQ2CeQoSX1huQ+QnCnFUqs7EYsKn/kpVEl/wy8adHXpc8kDYgCw
AbS1rNsI+e3Nfgo6XZkjyaZvpZeOB1A9Ptoo2crOO2L4ieiyOdPucwrBNVTWSLH/
tryOCH9u6/jN6UoXPuNdVapkYQRCFdhIqzDj5TMQAUtKTWZcYXP0K0IsGj4r438R
6pAZX5N4rgssnYCTV7VO+/htJ7PfkBa82q/GqI+pRs/arhbgVfAYeaiJEOT8lGYW
frXU/OQBEnxj+0N6PKhzrd5yIBDZB3Qhv81KBijD0O6vcoS1amFKa7Gh6leOcUKM
dsFbWgbB5y1aQ2pLPeFbEwCcjS+zUeiaOOz+x0UTDqi4xFANPBX49vPbKqk8mxPT
Rp75rrmxWkzE3CPubrya4t7C2ldsWMbyUeNtZZ+/duBFNmVsY+c8Edihl9D/YEHs
htlkdtny3j+o5Im4vywKiqfn4p42kbU9/NeQAWf60PpyADJkmaj8NVnw109CK2UD
QpOppM4gSlg/DYnQn0Qm9kMQwW6CNIg4B+qrJ0Mv1vR7a8W7TrCQ4fuDQcWeSe7O
qL+7NqoCG8H/FzKWq6rCB9hmMX/LnHbWbs97PaxacMb91KypW9ih+7FnlE81Uxv1
3xjPDCVPrsIFFNtBtcMJ+HbSr7HhVvoxGs4uuJ96Kymwx8/LdNPpGz+uN2A0bEtH
W/CVPACpcF+Jw77y7a09acIvAMNanP21WPSzDyLDRBCLM5AcPmg4uScgKF+lbcSO
oXhr5tE2aFTNLxXrBHtAPr3wDzVJQZg99xzs8gyB7wE6VR9zvItdhut0cE976y1w
s386zXhkXCxK1KbxFLaK2gBJQy930q+QoF9WNl44J8OVloZdq4ulTa4WgE8eu9Hs
MwOtPDmh0JNmpA4v5E/yS67UDtshn/hqFeotDHbq2J8NAHj6ONw+yITOvfjz2mYm
i4pokTmD8J7G1Uf3bT0OhO7nSkZlX8EoTlrdI2EdDcK4Wqr0s5LPVbbOxB0vF4V6
IwKJyjsikgMxikblXGUpegqRWO4jYYMdEvcqQdNJjxNzWJdRchLGkcfYJCmOhNf6
0ZzDfm/lZay4ByRVNQLCTZJckWhuQdEouwyJBCxooFI+gsTIZfCb1z8oRywlqP+V
KLkB3gGK5s4/lR3WVs15bcSlpXOTQufzlSNb6r18mQh0Fqm1mXAztpzz8BosZz7U
DkbVIhw6q6YlWhiKnG2dseRHIHeK9JAQNyYB9L5ef3MJFSt8ohlAIRusIcgwE5Fg
61z3fT8jyCHDkCN7lY8k1SpAZeFwkL3xL+3KJ/Rqov4Tt9zGULQXMzJUv8uzl4Ui
DosPl02byeEy5oj2assLKRBJB5X+xYgnQbhTuWkeLpuHK/i3H7smUHXMoaKZlIJ9
4AV8SCN/FilN6nppiLPaB1zYF5/FE4EV7q9S79QtVFhWs9Ql9ZCPzBbApxccs+vf
9pBzV99WeiM48keD8sOWh5qXXKm7DkCZIuCwdQLBkdSdqQ4QMUkT0wciFKd2IuRJ
nU6qyVjGWaQW2KShw905UjVi1/czJCnjM/knSnF3O0YNDT6X9G5YzhhLlqHs2gGL
VOulqIrrJ2Dnmi3FD/N9lto6YAlKF5MKfpYCx8iKt+zikBuYUemXpdbmGCmG6PHj
wZ3ZS6Jgf8TowAio1tFNKPf6dmW5EqjypOlVelLY2wyAXehQqgc/1MqQEQZSDR8K
ZiFDJ+tZjHI4FmZyvD13eR0VDNkyRZG/WY9pfjcHc+C+cSxQ61P5IJIZS/gx7Q4E
NSjgH32r/9iLdAKAd0JSJKr219lmnIBdHrGXPTON3M4h5IJR+Lf5+b/8KjbtJfll
uEzS3KgTRjMJMO7M1At+5NhP1I7Mywgsa7wSCOpm+HhAxt4h/XnyzG68sLvNGpaH
eKJECRwOlg0TVGt7dN623a9NDJm9dwjoq+jemHMfTALcVEACoOvwxkCpDzsw2H1Y
U+vltn3II2zXch+ukd9hfqym27H0OIojpowVjscjvs8eQOqdxtfdXZjpBbRHRbfF
sSNwFkG2MK6RqMVHMF2cbHYw1UhIWMjmku7TGh3v8nmWstSK7PABAZdkScU03m1F
jKat8Xq5HnRxsCoifqrxZWlCOT/rwXDdH8jJnutA22gSMCO6P4Qc/pb9cJsphfcx
iYAJvH/JQLIXokTT8+IAyxEK9Tr9PoL58QkgR9AjG2xFEQ8siHFTl4JaENL2ZkI4
lijETizJFFTNEAr1jUDsvk/SwhWjN/C0vbHt2pOTzER5Czus/PREq9hd4ajPrQZR
OUtiQaWVK1P9uxSXdRfwMaJakszdAY8c3Gk5BQRcUkXAufu7b0MwSgP1CmWPJ5s2
hlCarC5dL9jAgGf9muvaxqNI7mYm89GGFVwmsw1v/HbNutS7Efv9mIXhLL2/g139
NLXOdo6Z+Nah7PZizLJqxKhTs9H/dNd1DYBF+JLSh6RrskoiHbO05jrYvIbPuKhJ
+M3p6lA9apW3Uz/g6t4ZhfDzkwvrWq/Rhz92C+KihBYf5cAR2juGyMkSWjS/XBmr
mtjVb/gE6kdopkAbFkHYc3W9VjGKBkzXvk1jvHEXJuWWInG4y0V7gF//BfFSZTV9
WiUA7H6Ssv2qUo9IvfKIm1t8fNfs/9gPCuRbAy7BsEBcfBssxO6RQyyJoPXtg14M
OlFAtfuxYWxoolDC1n85jEsiIDZSOuvCO61G8VGK5D1tSF70iloTcVJMpAfyWgcT
vNs22xuLDhKJKCebU4t1V0O5S2LQgt+FLoTfo2U7kiERDjN1JLn2mRtfPjwjA8Lp
YJTWLY0TjnUmezyj3mWoidLn630kXhW+YxappBiBedpOCdcA8iqkPdADQbOcZUrT
V4M6nLqHm5zEQir4z22boKt7w3Qij06agJ+ELCKjOGOU6I24zLNziaDNB+5lMBwm
zp2K9bWg/CT9Dmg9R7VzNvMsynuzP+F6hOkv4XKB/vQcn2QMv+zJxlDxhMXp8Avz
g7d10s82+7Ku4G3rFzRJX90M55zUAJpf+9Kx2aHNqvzBgDaKpOhdrcaAbhijiOfX
4KrhHMijzYDnIv72gVWSeXMgPiiuOmKqoNFTBa83Jp8w/2kUYdjCU+1cFFycF5Sv
BWxbQBfcw22tw7i4yiKO0xATy96eeR2R8croh270UzdgdD/JyoOOQ3BDn2Gmq9/6
gIP+7jeJ6LFeZRscB5uZl+mwKEFcHme2v1bQRuW8vfG/NFRuVUq50PmVaITdwL8A
dIJJ5ed759aVFITeq7Wtlmk1MGBFtZEbELIZF4iPrm1I+rpJUjJbUpSlXzfqTd7L
++Oj7/SZf/H0RsDj2NeCFtjkUdTunYNR1dX35MfDpsFz//W89gNwkswlgstlNDvH
9Z0fHXBi5jIaYSGS96c+y/Ax7LL8jMCSMH8DW+BgD1sQN8RugfSTgxoBfiWjnYE7
X0WpH0TufZpeNqGadsFDcMQZ24ZwHXGLc+e+srPm4QRx+yngOp4VoncNhtTEZjW/
RLWuSi86uxv02rrKUw99tTBGq+XrNKOLm0PSXlzQKWHDOLImWDC7OHlo+O0CQqQx
qj5Pl9oFldwR/zvUi4ugdLBUSqhQIQho8dmOjiJqR/uicV4LSym26YKeArJpWcy3
u1ZOm9vjA+VENLgYYpNDuGkbASH2lejYxOi+iZi98HBN8gm8BOWv3lr6gkPDhhMG
5/grlCmiCP2qHX3+zp8rRxF0qJY60AaJ0Q51EURdumfueVSIXlcGAZHDsfVLtA/u
fIf3JiYLT/Nc8xIvfJCCadcHaHQ6JSLt6V49tOttOvCeoM9o7IFS2fiG8o3TGyRA
e6ILP4E9IXLxr6MN5cumyxUNwEwffDYrbNa/uRFtRfT/J+HuyFfiTo/VVx4t9e+w
rh39Bt/eDQ62CxREMOQfuk1Ekse/+33ib3wwGODDnqswSXf8BTkhPOTSNPImwds8
lkoiVN6xTqlX3RiRooRSo0CukraRI+OPud0vcj185OZPVRpbm8JEyKZPNLe5j/ex
xwySw1P2UVQePnQkdCWiyvTFvVMXVnVeo6UEO89USF6VDmsQ6DfLvcSqbt7jtWT4
qKHWg1amogskr4KIje0rT5yhlBZ6HjiBM4A9CA4n7FILpKqWTmbVBEQHFaoHkMRz
cb6vCd6B0gUUIGbrgR/okY/gac5213cX1F9sWg3DlKIU75Kby3+O2mukE9jVTcq3
cTAhiuhYxp3j1u8C+nLALuwl/IhMo7f+C+X/t/VvwFe8VvS9aPduqM+uauPM3xoZ
tpSMvFbeHRkZN/rRqHkqVS4xtr9XWAwyZq8Zb0F6CiU+7fZISFugQAa4W4fTDyYY
+YNr9q/VcFyNKsaWFTue4wNJHrJD0/QAkzArxtlkkjpIhWOaLduFpUktS54fr33v
t4gCvWv2nGEo+4paWPJWSgUgpTYzPxy1ZH6sgolftnF1705Xq2ocSYsROoZVRqk3
wj7rRJV5bM/QPhesLrWF8m3eh8MogkZ4rYRP2gCz3ChPZFr4WKq7KcPyVuZYOqO7
eeYPoKfsifAS7DcYF7p3w8vVLYLAYHPYwLnOb14wHPPfj3opNlW431sjXdqyG5pf
hsISM5u4fIo3TetgcI3VPsLQN42/AJrRDv0wl5O77+lm4cUFYUhSQ0qAkM/2FNHw
m0AODW55qyXx/Xqj9epG0UC9dvFyzmikwQHd30NBCSbXM6dlQ18VWmQlCfAEJpCK
HrN3DGBp6wSD4lF1BFLwPt2vq08sQJNszOGhQwqU4RJp1LgYy8CfMhgRLdi2sMVQ
UawgeVuVJDl+fmFQCljqYPlYtMVhFMtRnRLIiXGQYXYSMCrn2EvBUzcTxiIQF5BI
q8WQKq9E5DgkHPxHoCsmGbSyeBTWQYL4UIGmX0DZBfX3WXOUYchIsiPlLTIC/cwt
6zWlDfHe6LfaxVFuXmHMcDGLl1seghtuEdb8HeDKT/GOWC8WbY2BfKBU8Z24/KCA
bmYfWDNtm73rNRBGWyK2TDzPDbc2c/fxfjTdQydQCCblTvve5QOfG355GE4Oq/8C
+K4S8gHDgONUuknCkYvnkLUe+2fZ4DN4aqJOxcTf/Cj8WFaAa+9fxnsQhF89pOv3
AZTZ/L1QviOGQYmB23sb9QVM/WYSn/hUHvAcxooB9Z6Rzm+zXuNmWRbuuktmJLIm
nhiJMZ6v5hF+JOw/1KUDGjDmH7IooXk30KyiGjkkyadYrbqgBug6K97hSHzfmDUu
EbhJo4Xi06dc3S9aCpOte4q5sDxOHQr4SSgEOnXlAGYhtIfInIoqsQsgbJWr88Is
d8zm67FXSGVk4mEBqB0enk4p3hB5ahsjmqWfGDZIooQxg46PKsBmikeG5vAGfwnL
Uh9BYo3OGIxtV9p/xyU7LGMzMlmyb7AZB7+UiPfWQpx/DMj0debcE69BOpnbc8yn
Bse+RXFFTollqE+3OnsuQjYckLsHuaHeSZv1T6fd1sJTCspJrwjehytJ4HbCcKw1
VPBILVPpu87rT6FppCwmordHORG1948QRY2jDGwSO/zGhK4XFuwSaGnlS1WT79iA
X6imuhe7x9xnzHFBeoKsWsxklp/EtIygBGvVIGtf22ypC6PUefoVJzAwQgWhaO7H
p06rcZMOrbu5IgErCM3HrynvGS4H1DB0DJ7Wh5BCfaJXap9+tgCacd80iuSdkRRl
yREbiYqPsaQTH0mCbN4AKQKyEwkLEhoTo9Uh2u5RwYli7bG6YTCx7d98QjIj4RWi
1/B1URdQv4av2cA/IvztyhUO2X55L4JO8tjChagzcLHfU2voQT0SrJ0i8Z516JIj
D6WCc9ZC/5sEwT9v42BGmGg4o54oQR2G1IF6rscv7CxsPRmgGoG7JnkA6kcM5AFx
0oRDBUs+abt2zCmXZxA3V7HR7/EkIa2YCzEJwYRNjP1VrZkzguSK5RettRupXUHw
L5W0MoJNj/UnkXCLWcIRq52L48CA8PfGTfsaU4z+hLvTIUolAyRe9LkcPSJSdF5Z
xbXxcyYtP+opIAUTjY/yBb+hu13/0lHQ9OZK3TBDqwfgdrbUqWOgd0FPrbMyFPf6
q8tbri8+Hpc78F87OhO0KcNPz6/eKVn6+TB5TOtCwigtCnrVJrHcjXN0gKr60H5H
047QzksNhHnM0JCYULTXuzhERzjNK1FaUNBXRTP5gUQcnjs3pW/9vsOOJts1OFle
ICPbi0pntDthsWg1QZyDQ4Y38rx24/+mwmb4Y10u3osahzNUv6TiHiTJNxWTJk9s
qXeVo+o3I/ODFmz2vlaU8VXCuUO8RnfaLImmUUYQ8q6fqIDd4XvBsbhyxnL6+3Q6
ms5vLoxn7K3cuClhHTaTl59jCgbBO/IQCnpekh+iCuXwjwIL/h3kx5narmGrC2YR
gBfpanmtNh27wIUGuK0Lyi92n3dAfnNhTJKYDDZJcHva7tSpCnqJ/iKbn/22s3Qx
HvLwi9STtrmurGHG7zGuDUJ/7fPQfhl5huFOJC7fdyXxmzgPiy6GGH9TNatGTHkv
BYABdQvAwMZVaEYsQMRYJajLomqpZd1oiMgrjxcaAwf3ppIG/XQqeruIrQDyyRNX
8r9hlQFWxI7eos2VtjHvw0mURwf+bWlGJIu2sO20uJiahM0E/JG3wRFFS++E1V33
8l0JacFZC7bAgYb8cu1Orl3MxjI3yxwZ+Yc/1s7HoPHJYoMsak1M/EldYsQYSbvz
KoqzA3ZchmrfEIk4fRLUP83JnLRlRNxlmks1fspGW48mkSx/D+TPL7YlK5U5odYg
+GyXrLBpi6aXb1CrBIDkvCdk6q2tDdWXh0AtjnGrR8d5wADKJi7r3qHVAk2Zbm5k
sfkmOlz/LbXiKTJUc9JSk4nz/X+8z1n0mk1z3kc1CJKMuAi9AOnZy72ua53CTwFQ
6OUsnrgiV9xWWsItKcJfY+3D/IyXHVUCd6OdC6k4QXtR+9F3sWIzkxz/gHj5I/6l
CkWOu4OMdWoML6bA/VlQDzW2vuLADcjRHYYozQGpIVWsAa5UJpecCEmdBM+VtHOn
z0K5ht7TRjtWZLCPxKzUOAIc1FfWhCbWpvyxTOtY9mCU4FGcpMAgLFaTU1Ik5RyG
X+RrWlmpxEtsuWrYBfWI2mLXKxitLEOEIlsc5Zto9LuX4X3ow/nMwyu78J51qKdv
9nWj5rmQE+lTpW2JGOnL6RRtOuH8iuWYLCxsugYmDOxbA6dFpbg6BS5Ykx7SS5BB
sy31MG56QvAQ+papS44XdlA1ujvW4HuiYeALIB6/CpFkfjA2s/jVdNIUVPfsdF41
hASVdgesFG+Mc3P218AH9rxcXfxd3IYZ9LaX5z0Sg31+R5UEex9NguffMGuxTkqj
mpzKAaHYYUEk7r7S4gxpB3ppfG/7NsU1NmrJGp68deBEsEvw0nabmo0CYOspS2ut
Ik3ehpUJcjhN6SApXU58ORgEXMG64R2NISkfc6mZcVCdTCu6q6XppKKgWGwkX6ir
d0fCsBzWdYbtj6tTRouRD1g25aUTQtmS7WpLyw1L6D5KxbSdyAF+VNOcgdOVstCp
dMpWOWnEWWe0F7kthR62EWuSIRWwhVkDYBpsqzVW0qin0CA4F2PAOID/qGQYBGRm
LfH3LNskZ6qViL5PjMkqRorBGbQdpyBEoc7WG/0ebwkeLkLiTYlNOU6RQZscLjhI
slay2IjGsZ5Py4jMrLTIijwc5sC0w+vpQLKvBPZ5jh47DL9NwkVa8MIy+s1QGtfs
zjky0n4+H7E4XsG/02IE2v0yHhz2TfLjlhPxycZLqKpXgPDnJS0l7aDnCL+T4u6R
Jslq9AxYlwVMcaNr2NexlUdbHvbj583qVjuRzzaxrT6RcMBKwJGbBkgbSQxHOpK1
Nr9pewSDJBMxUmKa8tWQPu5ggznw5rrZW4Mz/i693szEODb6yOLvm3p4ZvKT0ay2
/g9BYwbtRyTWBnoaH3uQUmHaZyvH42vho8HLlNSEQdPFkBYg0zgV85L648L3SYRe
avYbDB2bv+OruxyJYs9dhQJl8VHz4cKJB/F7HU6hLxJVTRk0PkVahchGyHCUARCo
O2HiDuxyoVbBEKoSSsXG45KikceCKgUTkGv1BDkKwIMoHdyNsRnT7boNviqvVTnW
z/14kwp/Warikr1Wg8/HgmW4jTxhcsluCsop07sMp0xiEpV5h7K2GA2tD6ikCtd3
kpoahon9Ibo0hVlC986+D6hUurcHecKVZJ7kY+0J1arPH8dl+nxGPn9L6+i49woP
+Ry7niiEG0gIb/+1DO/6d6Lub4fSxjOyTLiuACTIKnFYC2jl34FI0VZB8zQbByru
igK3ncm0klSrjyKR5xvuQOEFUQpDHwFp9Ajsa8qUdYUjoumeyxNZ+N82WAZS1hrY
YZCd9DtBWQeJc5zXP24cq6lCbj2sV0dmz7/gzDJTmwJb/6OOunyNPVzYguY/vMay
v200klTxcMWKdGFfUFNaRu2ZaZuuNkCfTpW0d4/gjDKDI3hzEEorB5ASP2ZXWC1b
om4M4IUS9E3pA/0DY0VnqEMLdpL8vqorI+QeT0B0E30WgONKwnkq4NWNGhHtKRda
UK+eqj7tlZxUFnUqL49bQk7agj3SZNzSfNZNO8Gk/cIcuBAjBbbjh19uUiCb4CER
FcOd+7QZa29EdYuQ4wrQ6M5eK9Ulc+C38ykkQK0Gh3lem5pJG4EJOUqTfSBoPWNl
MjdqBR42cu5TRLthm0VKWuatB3pzyY4Esyd9Sk2TZJi2tDP5DA6ZO0x3ismxgosH
pnDD/12Y1t3tRufN33GRjFr4ROpxUkhcTZQ9xqurBI404KITWCXna/GCEjfNIV0m
c6LtPDE8Dd6Sjx0qgZKx2IDk4YBXhijLHcC7vRTCMJYy6wF8STKZl9yloaAizL5v
xV0B2VN3sG84XEwGbfS3AmMrJ9L7j/ylgs1OfztrHg+NRqD+hKWSkENIP80/gsua
su7gK5ZfnXEJlPUbcyCqD32t/5I2ZFlJyh1fEhR6Bs+zi7wgjGinL+qV3woyyu04
nNcBOSIjxXmMv4lit6q2fZLUcAxwItUxzYjFnraON2K6BToW3v8l6Cx1eSo6G5Pd
exu5epcFZs/MTdvZXRw+ASDZaL7baMxJqlQxnkR+0kHCCLQBHo8cqZzDthAlWELD
jnJCyyLDATEd9ND3skmylJJxmjrdMsnWUCEUSewHh/0HksuF8+dqZUQ8sqvV6KjC
Aaj8Ef9XmneNzkLz2Yylru8cmMOHT0X4iBItfGpslnF8qoxSV3lKZ8Q1qcsX82/2
a5NQdBWim2naBvm9W11dXYvF6TZRDwHK4Tgzjal8VAs4OLXTnkhaNeymX/df4Al2
DU+wrkPQB46zPcUa2lJ/cl0aMejgsFXCJNhIyjo5TjAVOK4oPIQ7M02JlBMNnWRm
S8VTuzcp6nQ5bDLCPyv3TdnMRJIOX0Rq+uJEXEbfGW3ESl8scXGUVqW3HblHC7TA
L+fwczLohrf7+RxdkRx9Ebmp4/oI42Dpp5mH85czMke1YJ7gFS3gMImKuMAIK1jT
uN+xUQu5Azvckdp4nizPlZvU8Ihes58K9hNq+0Kw0i69UbkxqrKVWFhGnokKzs6T
Gmr/lWR7YaosYlpJ0x6wGZYXF/iWGh5oKcIFgLyT9skwih/Yvz1U2An2YIGu8RXo
dpgvwAHXKSVNYAnaMCqvf2VCPExXDS0gTMVkZkjtgvZXxZ+X8XJZMatiwvJNR4pO
Dll5Rnc6ZAqT1uq8t2Ri2tu4g9/lyeGctPDhCdAfPXTg8BaX1XHC4KoG99MYLt52
jwt7gxbab41Ib5hZ14EI5Tu2/mFLdqI7cU8dEj7kP355v+msGks3ltoyTSs45gYi
aClAKAZVNuFu3MSezcjOxLao3Rw4mK8V9ZPIRqUrUyRmGSCdyTz7KBvNuKOYA6NT
laCkWNcLy9qvTVYY3msvdJTPJi4w2K5tTuzFTbKOy/ap4Qe6um2W1cxaWSUSxdKb
k52z2JbNtySfkiu5TcbfyrdZdzdf7XcnrugaSTz1Y4TcbHJe1uR08HnCTRgT1Ive
TtTTSKo7AmtfKK4rGHvniOieoCT2jDoEWop6Wh0EevK9/HeaXmTLFYmL84Gz6Ser
cF4vQLqi5ycd97kTi74JeblKERcN+LnoR1WnoJTJEYwEU+XNjbtExbO6M6S9yA/M
QbVU4cKlchuVgpbHjeJwINRu+TCxvwedxKombeX3xC14o6xrQwUwA6P1uXB7q0Qo
AlYImdjgmwazSfr3x/Y9W/FYk5BxVpLSsi+ymT30BSHb4aujp4AbZYRY1g3nZYpW
F6KnoItMJ3VR+Hy1DutC+xBGK5qArjn6eZoB6imE9sL/eAJICoCOeKa4713Cp1E0
XQP5RBdA0FUxhlBG44PZdKSze4mAtKfK7F/8Kn1uqojnZVXR12z03BIO79v04/Cd
0eSNcl55Mi5ZXE62MRE5wBNALZ6XaDGGE0D6womuSxC1YeKC7kVgzOfPsawZfaVn
4WblQoYeRqzltilzd93LHymxsrFOemI4yNlnCA5kbd7rmQGLQY3ojqelsXfgWwVe
tauVtq7DI1B8YglrJiH1cwnWruJmKmDjLyTavWktxRICuWUNc7a5xTVZwhponh15
nmHBQtfWYRkcJ3ZoFU5RT/AeyTQ1muY0oC3WzEd6RNBFqxIyoAYCTzvazEQsUvOm
iq/Js+ZdbGkL8fI2iSBDQNOr7PBvBFOqFgkZNq7jBWteQUawnyLcaUf8w/DtQAJI
6rboP9tu5OrKjNP38VbU/8LgWZrNPuWpQuFP+KwfpHRBm7ksFeuU9iD1Ws2CMUbu
iPpupFAVpqW4bPImQPEEBrjaEnvYit6JaCLdsWSx70P6D+jeoWeTDsuwo30B60Zu
IwIon02iQYY8EiuyfNWSsxyMkuFYodzz81JYGN5bi+26DO/kx6uLrP+ydeMNogu1
8Isr/U0PDn+LrdQsz+BRCB73/2WUeeQwLwugbPvJn2+llYFygNyBvoz7tL4OMPcF
e4TkFKJOooK/pkghX+/mKE0sV1fpKwFuhdY0Lc6PgE8tcFO14CxlOMDb6hvLaHGM
W8PDnJuJOMFmxIxPqIIYQXwh8i0w+TZADndT3qVx6dxCQnPEJ/QyTe4Ayh7xpZxR
8cgXxKSBG2vegvJAShpejnWtFPAVIdnP8Wnk7GXd11a/saSULhD7WwMsjCAV+eY5
JJ4N04CJzfECylgnt71fYT+gax4y8KYeDda5p3oUHuVMNN5JlrpDmyn61ogp42iT
LFFQgf7E23heCIjXqARa27+scyUMyh2PJnUhH/pHQBee2Z0uFpQ2UoVcLaG53U7x
dKcfgAhrBnzKISLQtBTrwRe3hz9J0m5BRNT+He5uWIjkof7Y1thvutdiP5yA7UfG
XTMcVLti/y867CopvYGteW3yx4UIDQex9UI0VDOBJsxD147b9arjeoNGp2OmN7hv
wI1OJQYBwqAjjEyaa7MSOkgdRjID2N/4W6Qc2xIDj62je8Do3P2gD3at98aL0w5v
/ODzBMahTnYvEj4HQgukE+YeZMw+r7AZmUeMZKX8+LtfxvuSO/DLqunz8s0hHFCe
gZGeBZiUH36liIWOPRB4//svcJOO2N4vhN/ViePprNPSHKD8HV0MT3WMV6CFmORu
Arco4JgKFHpZ283RNreuF4ZBI+chwn/qLfX9EzllR6R8D8tlwCofX5RkTKZn9M2r
Zu61vbJAm0RzsBxBn+4d8/ocyIfPFR3ePB7nMsplJWLCjKXeiyScUZO64W+AEAWv
pZFz9hZefzXLm80wbmKbgKxVOGSur81oIuXlvH+PmaxjK/wW4XZmEBwWp61828cx
V+8O1alCONT1HHO9YtEvoOrmTbqBTbli2QIp/OADS/FrlXmmDzWbW+ASBCHoIkUN
c1W3sFpK9kHE+1hcF4q9wlPDEElaiwb05/aULlrLxK+mCjIlYVF1htGlJAqzW1L+
/M8DMowZ7eUWgKOd0EU7AC+TsX2WIvILXGUm/Wk0W4YEC/E4u4YSEikdnzxQ05/p
tooPuhBeUsD0dr6VrgSaKzpR0FE/mqzgir2VrjmbGKezQrMJCXhhEaGp91VTEyZH
9g19seB3HaQxed0T31MNFpnAAs6FjPdYXW8MhRY4orvbRdl4GFVTcfpK0kE2OANO
Y8I61PDBBLdl3ehVJ6lE1IdK4ULMVS3H9nplNX/E0gCw9602XlA4izaAkII+aahW
UvE12Jlc81ZuYniF4sNby4xAXSFIv+lTYy+mRa5XvzBeMnJlVUDHnKI6ufSlyyeD
DRz4zI6T3XKhtrlgS+8HsNCXHYX9HiRBWT8RAqhPv1m9jcjh0ITxGwBH/U+ylkTh
WkPx9rWBhJl0Y6xXE1HiJtnNE1/HfYGErdXYJ0lm+WAyrxh/sQtIrHuYEhqKfayb
OHipSahs6AYkhi3w72nyWoDC5b41/HlwPgqL0SUMibK05dUyJbsrkmSNIu1WcZXg
8gAA0V3kjCYdtSRP/DTF7GSyIO2YCYTkRjO3OUKzKM8DVV1hsPCTBNqF6lBt+YNu
Aol60v2U8LTRMaX/Xwsf2ypBwPcP5g1kA1YCeKk1HlDxfHSy2H4UoztJEaVHBjqy
wLRxtMo1jTFBE2RtbN9tq55QmmfhHBpBsPqSQ0E0O4N7m0VZInRDZMsMRJ4NgN0u
oyfI/WeIF1uZ+id6aeqSuDe781MnexW12XtRQHEQ0t+yS3XRudKQ+4HO81zke5qf
DtR+8lqSzqp7N6p4KgxAD0r0Q/EB5YpJTMpxmUBSOEd2CFJDaErb69MtFREio3nw
8dpMfSoGoUdjV1ph1iliCKQC5t2Ag2ohes6pcHyplUUzFaAkCA9CQA7XTVZ+Iv03
YXBmUTXiptScNnGicewbLuvjVNo3PsKm3ukuN3e8w6IAMeHJY8zDQlH0zwQduoaL
qGzGczLkKOKnKcZJ3C1lT0W3Jq9HigoEstdlDQxFxzTn4ElEl4XW2Nlce2lcGgJi
Q0LXMyLPZwVU4L0hrwV1WO3qfJmcvVMb/o4gkkesOTOxsi1lHCvzJyxgYkJIEcj3
PhL5uzGwDfLHX5tUP1HMCV2vU1pfxapi5lvxUVJ7vi0vGaXmq23fq/SoZAMDLW8W
hnpnDnZOX3tSGb7nYzuA7Jqk42Gv0NgaRiSnCYvq+XM/Ym7Nc2iUGaHWIqEktWgs
aQprxniUnliP64G+mOj2BL5UlKiZZD0v4ZwN+YaQqUVTlf+9WY8hbJogy3V404p8
y0eDCnsKUMu1Ikg4qRnq/Ecuo0I8ydi/C0XPHDULQt/uQ704r4we8rZlPMdXs3a9
7a7PFfqg2bG/KBfoJXTCoJFqUcJQ4kBWG+LLWJr+DW/nCKLSCqMz2Gf87JLN3a+B
kmdrzKW3BowiC9H7MCKjx6KiDFihbTYwHCzBEqtAiv10NtAE65gUpWH9vfy3v4t9
V1OfeOdlukP/l2xkDrcXn1uzszGq0a28pn7WncSN1xhhzi7mOl9HfIIwUevw+sbu
Wy0m2WCm5VZPzm4izdDrGVOtI54R3HQhOrjKC6VKvTT/M9WYbSSTgOccoKsjj6yE
flDwb550JX0Bics1XGW6EAauC9De1v7u+w8/bSL/VqT8r3Ec2iLojfUUdyk2MZdY
vv/UN3DwqEJYdVCr3rJPC9IRjLK9mtjqmOHiHqsuXF3QqDhV3s4k1z/md5Ed4Icy
43TTnzSaem8OMX55HpEYt54HAHActzNx6TQHjTAKRL3+Us3Xq5kKH/N9upMUSEMx
kDfFBWnzFRpMCbWWKCSeX+Wv0QCdFGDRODi6RS6ik6ASR9mE3vBdC1PS5DQkLhb5
Z0nhUSOY0qJeqzNONBcEzNGo+MIfoEtJU8JoPtvJMMExaUUL5JuG5iuVTuU2+XSH
aeagfNYnmlyO5cJ1d2OFCTAawGemF+50rH7LTbaqIoFtJw15oOro5w7T/yR4MEO0
XE1RnjxGfyunulaHQ4QU7LmNXSxIobJeXp7fBuI0mqD6BCJU2Iw3ZajKD/bvxTs0
KrvQsVgi0h6vF87N3FxWjuO5+1nFaJ4YpNr1H2gCz3vMTOCS2UxtrZE+xUd+S2LE
ZUIZslOZDeutXAr8ritADBGqBrsw/R5bsmQ6TabTBdy7gzEYYmLwYsSSUSx4bXU9
/lF8e27RQCYRQ3P34gUXKYpw1yWr3rGkq4d64HFDkW7gZRday30VQC/OBlmTyYQk
U4fo6aThkJyrErosz9F6eW0OS9Ax+Wfk6QXbn52EQ0sE/fghawhQGhaU0wTS2Qpb
7S3LmFbx4np1f5gt+CLWJqxL0/RxtFoHUjK3/eP7g5qVb+2qUAuMKq4Zj9k5R3iJ
VgXXQaGBb04QKKSBQkCahxmtVmSzgJjTjofQ12Tr4om/FCXYTMoUnYTTVDYV7OFY
A7X4tt9FHLZWHz5zVFe3hSPGaaubXPrveQVyi+LVJ0D51Z6IAyuSGBVn9og7T8x8
QOFjyAgC0SZ1qMfF8ABU0SP8ydfbZOW4LO1AAILMAMcSdG8JNwZAvZVsYKXeqQEh
E+NZV5xQc/R9+/nU989u4Tstk9ceTOaM1p9OxGijCySSn48GzZL21/K+acgy5do3
aHYvXPWDDz0zqq84RaEpnLgos1rceJagHfrkT07czu06+z2JlFr1StwKkbROxVHX
H/2PAXuKUOIaAtAoGmbhlz55fKsj4hJCieWkc6NDgkdqkI0jPfKRRugFeGZlpV0y
V5DnhEZH5ABQ86dJBzl7opmmnnIXNVlB4S4/T4wKlN61/63fTqHaYd3KtDfiJZzs
1qSQYrzbQXlmIlrNQcukmU9yUzWCz0d0a78ahMNt2GXc1j9miR7BSIe8KU8TDP9q
cEzYJD6xEE7xjHCLxA+0c312qjSDWxz7jPCy0lc4aBsCPFwiNOsXwH83Go0vBRxU
YYsrVu2V4ZBoUSkh9HuJNza1YstsUDX8zAH5jlxwzMRrRh+Ha3Z5FG1lYMZWVyP+
IhqT+0/8Dwnrj/+UPM4gFMfRS76EgipeEjuHgxlavVJe/H14bTFLWmFCidwQI2YW
xk999g6+VIWv+/NwlFgMKoyyELW6LkLn77BsYJN55Z+oKp4ELiQqSoAA4B+Hm90E
8SuqkJJ2x0EGy/MCk5O9dn+EM/ozXlhw4iVUBZp/pU7cCSx+9ywn6b4K+oiyCjcY
n/4zpDkHyZUcnbC6VWzto0D2kgY/qGpQGB/USt+tBIB5NIcHkVHmaDTtCf47NHaZ
dV+8RpsyjE8X0s5wPodiy4xBVsdbHdQhkgIPiSb4sdwU9l7zsx3UYkCR6wo5YS+A
tmVk3O50PLew5LRfrzoEoLapD/cTx/qtMt0RiKEvd8J8C2nXF5ZCrODA/uwAZBgs
jp5Ls35yDSQYm1jfDhEz/OZ8Ha+fMMkN9IcaQMyGlvB4LH/jDSkg3HlFYKoWo5qe
W6WbC7j5/2HLVIlgWD2BOD0p/mT5ZLTgwUgOioITAkgvOrqxEFZKu682IHYu0kns
Z3+m8m7Y/epz+4xdoxWjHuDNRvuB1CpvwnEV8KaSq9sk6Xa9jrfhI1QS7L6VNc9c
ismdGVhnWVFPDqZ6wI3je7l4atvaNdhvHB6jXHhmElFpeC98GCvNHccgh4aCOnsL
iCqW9pOw/JJcpYENavsrtu7NfUE+u808DwxLr6TXOIbMloVxT/3zLwOygCmSZcCI
1EFmXLwtPuzzoCDl43lkrnOYzNNjf9ZihDZKqiQVasXjuZETBRix/XgXd53Nmx7A
5/HaaX7ru5K4IUo448z+w9UO7BgP7FHYafk4gGYzHEMz1zV6oZVDGhXQNzd9W4zj
uf/NW0vAy4Jf96P8koypH2VT/Btpwp3P9KHkU5j92U1F+LxYNpCfFknpeFBqkWXD
bQWUMQ+tqQyhOHLkoAmelgqpQubgjT16/4sA1OdZ8D33gqjN5Azrxb4ugPgLv7SV
406MvrxLTvEpXRwNsZtbFSqZQCs0VUtFbWUL12JehmFCjiMxhpqoAcw+nhxaKY7W
zFLEPRd9UPFl6ehGc987dHsiTG8AbU3iTFPU36gpl6eJY7vxzsomgE0bKZqcdYP3
Wr4CCP1xo4axrVxQBBo1zP0hmQNI0GCmm87iP9Shh70n/v6oX+gA7Wz1qIKkIpB+
2Z+YFWXRsbOXEQin5Ri9FPwH3VO+CQq0+TbzRgdRBuT/68u/Pnyhf+Q7/Q39S16y
yCPNvYZ3K+Ro2WloY90Ksh8wQU5eAwJgQjxlmC4VHiXbivyxmxFDLjgmSKSMj49f
xmjjcQxLZu0NmvMbDxmQHagJCYdroGlgpvIhAPXIuRpF9Eu7pGghiSwVutn2Ekfv
lB7455sYFLSXaDGD2zo6ki7c3YuSwxmd41zUoSn6BtfjQ3fjLRnccQ0CUDMvOcpo
xQjhgvE0du3ox6GQk8M9TNTHpwwI9nuiMzojjq4Q2IjkGs+bfVeOkVgGBNs8vqX+
HfIgQLPFtq03TH4AgBcZKPoiR1hnOgpji8sdbByCBTLmEth0E7BNzZ0487YjIZLL
tdKf3elWkWTIQG0Puu93+FmnW8cs13adIFg8WNxXWz8EWWlq5c6YSh9Fm9MZs+pl
wMYm2BRzL21NRiOS7FlZZINKmkRGeqhR1JVXuhLAVlo2MvJX7ksD4m2XkTYZBe4S
0CGoSzE7LGqHUOUZv2r+tGUoK5cygx3nMui2z/xA5cyC7zScXTJvBYSE9XrKu+uR
Vp4/HKXKVCHozHKYcIqYKMV+tnX+q0oHkXfyxpucTtci9KboYcn/SD2G2z3AmNIP
iXROYj78FEzfTK6Z6y0f/2z5jcpsdX3Z7nyy4AtYLK80kzHf7mks8SoueeJke0Tl
CC6pkFfEHmJI2dFPUJ0UPg7ktEcyOPJ83znC9TaZuUZAlluxyHstm8H+p2fj0JYl
xQIG10vgPlVX9TnFvKO+7WQxFxwUaSuNlE8i74SWpVDPZZIk5WlxSDSHLwGK1wxJ
8Lhqu/YdPlFmWSfQx0lfupoccayehYpVCI3bPykZNVKDm68FDF0UcPYI0Ej+ESZQ
+KqTw/4YMfRcDEEc/KsnlahcoDbQ5lBC1vw8eK8NGjWAEbd5LJQQwK8vGgxbPdjU
K6j9OUHXOcQo/V52yR0CcneUZuG5S1jwXW1bfMnw6zurpKbLIzbMLhGJurQeRhNZ
pjIOcJaoMlIhV7o+N/ESKpQ92oZTlPkglnhouv8/RAzOLKB6MZfawR5nkGGkJFfG
tmlliQWiizQzznVmCTcXJNwTwfw8bRwyj+hKAwENghuHYCMi7jBrdW7/6YVKZV6+
l3V2gUuGhBJhD5nISmE/I8qQlMwPsjm3X7+9YM1PfToQ+8pw2xp2OdWbjAZhoBmp
huFbcYDED+8oOLnG7dBU/ZjwdZ8fMpkO+drUpDFBjdXL14+3nQjGL4VjJsqp4PoH
/WcfbL7EcCnT3fxT60Y9m3HmkwYcAM+yZIfoW95yErKkq/dTXQ+bsMhlErHdy28/
JpVeIfahv+Ktw+r9CbQQGk4Nt6H0n2alXldFgjlWAwBH9T87YkglAgP34LP+cUV5
`pragma protect end_protected
