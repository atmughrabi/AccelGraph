// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
+5kiGSzbEM5iKf+zse3SGPMjjQP3ip3HvgifEa7saOvMiCJhsq12Daw1uq80pHy7
tx6TwV5uZxjbmo0pHOIzZxkyyGLyp+unBKZLGbVv0BYGKxiG73D95gFlixt6pT2c
bt2U8PDx1yjgN5MzEerFdfUgH9Dkv+mK1UjREE+Hau4wYYeIzwuY7g==
//pragma protect end_key_block
//pragma protect digest_block
npP70cTpEhc4P+eKwXloO6a6kLY=
//pragma protect end_digest_block
//pragma protect data_block
qC4YvD5d7L1NqUtvH6BlbQvLXm/RvFltthzz/tJzQ8pDK/jddyXKmUj3fHoUWubo
unW+MRhn4rlkbQHdSdK2bHqNYJMvNxB5eicbEKLY39BJ3r/8Lp0coZnVaOg9U9P/
AxOyXAx8qcV0Xq85ZmxCSkfqPZG4zJHyS8raFIubU6Njsg9LSv5Y1tmzrupP6r02
s3HsehiA8cl2PBCDHZhExOH2zQ5WGe0lUZ39nyZQ4BNca2k5xRmOzVLz2fjLmm34
76kig5QRwW2NhodOm9x7eyOO8PJ069VOg5R1W8kOO614Mne8su2vOkB/4OoTpwQd
E71/wzHvdXU5D9lckLbaqLXL7pPurWkG2ZogatFYE8YPVs4O3D8VDCtaZhfCI49r
N6ah+Divf5VzjJBBvzdG/VX42KIVg3SXHJd6GMohSyRsttXgsp7vlxYRxvtPEBi+
FQD39SVJ6CprraaGmedzHCuU/toRzHA9IL3TELTE+OXKSUSlYllmW97CUz8BL60l
2bcAif4qft4yTwOse98oasIkSiYwdz5gPbn5xbvAiwaWV4OObVi5AsMRVAU3jHjb
xJ8U9zxU0//WRBkyeNJIXjb7D4MM8WMVPN3ef+9SHl5/+xkd7tWf4yPVofhEOLIc
J58Abfj0haGTvu+EU/uFhX5+Hmcoey3nXz+FNZL2m5k4NMODTe5KJVtUprfxu+Pw
hXWB4TwpQeGlC5VthR4b7yaEwU1NNsbe32gzLRnIT9M0IEBnUlOhFQdOepi2hKNB
DMuCPqhBtog//T1vW64zYiopJTaH5QF0HUmJgoyuBnxMDHvJRXqmuUTzGbTc4Kze
KIvGL0GY42Q10T0mQFKdGtI6+uhFOkIpGASTf2QHsC3G3D2uwYpIOxRuVVTrJzqa
fZ2Y0IYaR/6scvpx3sQ6xnF6vdRVYw8dyZd8XUC3Yh/sg6fh3v7jir4KybIXtp/h
Awkf25c1WV1Lps2NmrideXBWTLHfZIBKc97MeBAWD/2ZNskDTK16Kcm0RbSyny2g
RTAPuKZLIb4ZrPOZbpyWezasi6+CQizKwZFw1uusRAQGV5TrAOP+J/LrYWM6aBNx
4HO9PQr9I3Z+w/WlL1YtNtkE45LAW4JD2DQZYZhhizW1LsZMYIydqn8fTr3P6itr
7w8MnqGSL7hqVvyJgPaeBK+izowefiJNdmCq+p36AfxYsTYukad97tNHdgHuyEce
HmexIlQJUG+whpidQX7rvuzE8sZXe3E+QdlBB5dFK7Lbrl82pEcCFGfViYfL5HJ8
MgnpbsErOsmU4GmW8p1sBd8QxH4vmYxWtq/V1vqq6eYbrsYKM6D/DZgHR4Jf458o
qIbueSGpBjgxvXPbNQ9igEUL9U8TPhYpxGdd8HztlyV1LIH6WwuLcS4dj3nLwgkK
p0ZHPmgVdSmkI8cCxtw677SsymtnfxLrNWrfJTXex1AzUxzHPW7muErI+AcH6lPt
yotIClc4V9hfVt6pav8prAvRYzy7tIqqAFz62d4VpzZjf5a4p2GzndhONu+iFIpo
f36dMSOXkbIZKlo91qE5A2Rh0rWh+fkXJurOVd7Y6vOnDSZGUremf6HuHY+J4f4B
4q34yxKIiyJW6KaE9Sd8aFugng53AT+Z5e0fQSSxfITya2pcHlI+zz8d2aVDy9Gt
EG6vqyCbP7a1QwmDGtHzh9U7/xYOGFT+fBvjwWCl9/9RKVeO9SrQKw3/IRixCuRH
79ked03qK3N6VxOXHuQKH5fNhbmd52r/2X9JiUwhGHtTxbOsvuMzvF4weuf87RKc
aSerRGXgaPb9Z82XGoWF61KHNtWs34Q1MRIhIEKFrWa/b+Z5PNJ1oTdQ4++zW8kx
9XrcLay1MhqTFDkisFhVR/kg7Wss71kGFMnPAxQiw5/7ntfWZ8ryWGhUs/PwJZJx
8bxccPEg2/OZXdLX4d1ZLEEMIbCexYEYO4gJHelXGAfNQ1rPq3tuVadTqUPDAZP2
CM3JUa6CV+KnoI9oW719+7c+EyXZBHfYil+HVVtV81jvRFj/b6QLHRsGa7978V4o
yd3mehtwZ+PA85Vo95kI/TXJ53wlQlBh/aEqaZH2D3E734iIIWfkF3E0QtvW5kwp
FMQjAy33/CT5uSM4jo5eF8a02f3xiqhLIXvjbT+xjWGHG2RNM6ATiLMXFTyBuGaz
e4LD1qW6JYnli5pvcAp8eSjfnFQLiynM8XcUFoznJbj5pch4yt0limhvoZ0+Tf0+
+CflynMxgPX/6uyQfburXRVQRaMIJ27cQWG0dbxknwD2oQVDdKZpPUOtIrTWpaPB
G8XxNjsIAKksvWZzvaI2Oca2Tv/YZyey+vkHwk3JVHrs1db34/WCah9a6BI3aP5i
2s7UpgtC4fBS+g9gGV87rXNHyHU/ATTFZcOKirS6BChs8VmomHFwQVhGcoXVfkf3
Ok3Pqq8IHp52x7GkwLb6Fq5NE2fqf6xBB1rnBO9XtAlnrUalTTxjYfo55OlDMjsD
n9+ub0du9IURoWYl4HHtI54LQoV2DuzsE6Zm5+QW/UkoZZm8EK65lMHTifT3gIh1
rY9z/qYOaF+ife6Rwqfza3aWI3lKjzLx2ISHq6sYMqhxAc7h1+bKjkzuJ1kUD9WE
TuU6nh+Iw3XSlMW8vCVO4IngA67SVx9JyVQSF6vKIh3/ryLaaMMmj6hQAu0EDA6j
miblDKQPT8zfpbXV/MzJVXo6oEk+uKLZqX+Nj8cas5EXQQ0wSvl6Ge1DCy484b63
tGDhJSztXs1G/vbi6CQ0rsL8s5JV2iPUxR+2/1fA5le5JcN236Y0HREFch6p7aaH
6+K4qsCqK6a3eWYay6wsXN85xy4gkYghV5RG4l2KspVIUqyw2ZOILmd6AyEHiIwW
nAiwwhvzNrYmTwLBNtGxHdYLBFbKKm0t1mpa8NkY0i7j940JdanoLGey9qOdBeH7
ev1ydLsVP+IjC2l1sMJE5mR0d05ONYSgW0atYHlftC9h4eak/mewu4u5Nm4XtrH9
yT2JllanNjXf/wimSQEMSXvpSsR3a1RFyV4a047LjdNBY8aYjMAKirJ71TNAq8Y3
Xl0jnLu5SaZBbGxRyg0ciNshT40LU/Km0OOCwGekEXFhFzaaFw7MrogtyWawHD8N
e1rt7BiwvU8+X1bUasVRJ7DaEKI8pvMLzgEicHihUbhM3xYGVGDs3QzhbPoV9rdc
fAMPLkTeoC2PS6Q6hmx6PTxDFmOnHcQUaxrg11E7v9cicps44c+FcYvssxCpzPwn
dz+TQW7aOR/k+153iGh0Li79XE1v9P3froXIPxIEzitBNBpm04w4488N9UIBDGOu
kRQSIzZ2WsEo9HOGNoTCN/Cp0B98d07f59xQyO6nNXVpaiOEheQD3wxqdJMulwN0
rA7cgAMls3/nu1As7Vw0X72ZB4R8AgPwj8wdjItQ4RYSBqfHio5IAEzk1EXU9njY
17/qSQgbiJ72Eq5+FnXXfFlpio8uPlSqfhIh0OH6A0kgNo+Kqa0Q2eLMplyln0Gq
nMbOsAH47dzF93dvU7V7m5tYLF8uil0kmbEp7Nr9lvWIhQPI7zFOaHeplZexsprs
o8fe8xPFJoWjUcgTSzHt14lxwnuXp8PIooGTvYIK3XN2m8vp5ezW0FY6sKJdvvve
fainmx0lsND/tjLBJgI80yqPNlmCVCiZ3uARW9VEwX3dm82eLefmfcuFEuw8CdV5
bv+ZzT+SSlM0KMw16ChO/U04pYdtWvcFcRLM0ku62oOSNy+MQ5Wng/cHCrbKK/tx
nKOGYZ+5kKHbj5E7WCbjdym63Lbms5EXNltfUVxvO7JWh3KtCtzuEHWDu67xijJC
BbmV+lWf6WOqlLxAJlk03GLz2lLvN81C4lSF8QzSG8VnRe+gPsy9zdgewe4e/9OD
qIPGBRHiwLDHHC+fPCnfCKzoqFxDzg8PqIHyzKddzBkX88s3dtdKypfY+H+tk7tN
x5pLx7uu1JJvoj4CUFhoL4v9mHT4SfQ4i330aU4l2U3vs0NJ1ql5Th11taq9S7yc
oJ3nzh9kOFhfCCqyIgHPSRPYO/a/0EWPn++Nl2T98FUHZIEYCT5znseEwLkVAclX
lTJuJxdJiBwZrCOw6HLqPsjKot6jIBJtk2pQkjyKfcIViSlW/u/B4Ky1VfiZGOl6
sKFqW2czPE2EoLmbYJaKNnV0PzMyMKQoA1DORne9CTKViy6UhbeNqt32sNiLEPTA
B2hC4FbDyUP/blw4MLKCYhO6EMtx+PDLBHo0AXRfhZmh8KDz8rkhAPQnuJWIjaPl
aTipo7vcTjbjN9gkfyBQtJLv/6WuQTjwckNMKPGjc020XpWvffhj9Gri13H7Fgeh
QyxCa7ynkhZTtKv28RqIySHFtwy9qhCjyY5wSx/dXXiuq44noP7zvOKpzM19A/zB
HrVjG+DK4ZE7yUkXyqIl+gHX0rA9ZEKZYjRueNS+jO0TQdU5yhc8lQCe1jps+AX/
xtNmb4efWWQDSBYaJTjvIgkV3m384LrO3MN1g7/EmWluXvBQAwvW9adicM4zTlip
AmZ3xv7Ej9LMKIivCGFX28GQ4QkKSL38fsYNK1q824hYsn9X1E0GHt7Nt70f2E/e
WFS0p6kaK5X0mApoGZPdlU34RvDlBtU/ugz5MzxkNfCL4eRXJJr1UGcOFLfqyrjh
ZnfzubXgGwRMzTTQ9sXmHlNt3VIvgHMQd0yYxc9uTB4WzhyTpvks3gIZ9MBNdT8X
193J5Hb4MrjoRZP8/zdso0ENuvlIehwimo3hUYcfeQfGb12AsGan7dbEVzNt/Y2I
XAl/gvrmjSEodn5p7NAhCdTTbF/kygUEH/yPA5O5lakZ4btkIIxeLIrbgXxo9Ofa
fIiONkRYF813jFXbQmdZ+0DA7Zb+ooZIxIoUN+fZvlnu1QTR4nErQEpFZDlBPsqH
3r/voa3OWx9UTfwqfeRApNTtJLNLlH/sdCGl/IqZoHUUeXpb6YtE5F6BjyomQJo0
BI/xI5PDrjK54lB+i1ECrU5PzFfY7maX5L2A9lf6d/1ePQ8YQVt8Q6zOhhI+VJu1
/xuq02bsY5GiwZ9KYOxFwQbrNEHldKRk2OWEh3iKeIgs+PKzn9oi3uUMGjHoxm6b
36Xgvixf3NZimPGm8mRG0xX1lFvdCf2B7UBkQK7VhmXOKyZ4gqDfGKGCfWv9Pkp3
uVcumZEmuiynbaayfnEWrufjArbdrAlAlM9TQtPKxGIl0/offgmmd6abqbJEPevk
ggvL+Z7S1gHVngIZw17kUT/XjKPAplnX6ZkwpNlI+ptjxm4iRJ++c0/kH8LWe3x2
T/3CQRkSctaAA/pBVCK/NCbKOh5LCrDMsYNQ05oLxvtEncoF3/ul96z93G2qmpLJ
0ojblpkifFUAb6YTv33n7Si19S26uAjxoHmR30ut/J0eQv+7BrEgwn4LHh5CE5tc
psXApfYqjtNriR7y6hbYx0TkstbcdXqneFK+rUe/FC9rIDmpQenUykrMmnDSx7iX
raaiwxscFmfPdegyAp8y3rgo3Boy7LUhsFrxboIHuMTF8bsrt5FSyg0N8qhO+2VF
ItdC3atpjVxvhbqRv7yNmMZ+ZVLr4JlgTxYbnky2j5rMR7qUYi3GRRG44By4Am15
2LaDfYCbKBEVJ+roXH5XmUbrI8C9A8zTeuA5tj4SwLonBSscEEMCuNbJaHhsBd6q
fcvZuDfLtP5RAU8seRTC5tRGbYqqUc32fPtLcEfrrajn3xo6G2EaiwZAWxyqr7JP
jKvhQoI702LUZ2JrnEW43dZWlD+ypdFuP3Jf+26dAtQh7x/aYmwWndxZJsr9FAAy
mbYXGKx/LSWKi4h07yRCzjZiJTw9c9kkukMQIJjlRfcz19aZ3prfPyCzM5QdfYi2
iR9rIs5+rAOE4URDyO5I3gZ/euWOsm2ewj09BLjIQ/y1HZpEmhh2+/edZXYBeTTk
g2KN5p1/iNB9X3yELoZWtSAsr085JKdieQ8CgaKVI04yKxWbBkj8jxcLKP3G88Qz
f5GoWvQRX51mEyr7o4s1/A30JfcDCowKmV2kzjZ+5Zx8T+6X6Fr5MgOG4uGCUCh7
nM2dVDVq2Xxs7eUciOhs5OWOKYydfDb1ReiT9jQFTr2fySXPt6KqS+dNkT2WMj8y
4D3QfHepDFLmuKOGgV1Xu04/I0AoeXKpsHkJfTcZUFwWFh1LMF3k5Molz40nWoSX
mBgTItTTNEo42Ge7/AThM3OABRrXCHr3ulRrx1/df9pphhXPTLWoQRm4YOIpwWme
X2ammPgKUwXLYWyzDcIW5bUB3RjJ5834QkotVQyPGxkZRLUjdNpQQGxnS7BK+sRo
dtEjL5fmnEHdqDyp42ZnzRttQmd8mVFUoVqjOB1+JFgkXYHOeSHZ6VKOB2CZIAoA
A0SxUHekV3hwqQ3CrCFUEC6Hw/Eiupd+/PkM3gGZ1kEwd5rRcCLQiGQ3y/sLwoLl
rGMDod2zavMaLb+Bzfrg5c6iZvwB1/wV8VENE0FPyR1Fqxqf8Fwfh+qL8WDMj8Vb
7ynI7jQIdUCPoo7xWR/6KjjJGekrcuETY0gazxb4gqxsvms9ZXlt5uq5w1e6Xdqi
U8KgykOO0UldXoQn7N2/wnbOEVer2MmuFsxRpVQpz8l259lfpcbLtRhs0pU7V14c
B5zFmcw3wI9RFt3el7M5kgG5hZoiukvxgWI1k+hWTb0FuN/Zskhy4YjTjTE0CMO1
f6PZ0FdPcZGz9M5/YiBTQBje+lsiGyV50PVBoCTu25IXeDID1aqiuuvxJ9Lbtw0G
+aWLG13QDaVI4bXJyPKFV6FzXeyiqQbnvv7/3XhDav3bMH0EFI0KA4Uji7LJ2LrW
2gKNtcmfIqKwmjT2Ly2RK6FguZof+IN/MbX8vEbrtDGwdfblUfKBxShhg1zT0AiG
OmAfWttrFQCSSIHUsP1MIGbIXhZULXqh0ZEqwrzjj2wAEbYluqNmC9JTuCRuzm9y
r1TAnhKXRRo3ZU9QLzCWotqqSt0JBO+QW1WOrMA6wzVlUDS63r+eiEM4XdV5Jntz
5N3SJimKPSPZFdKJsgbNXDcFFUtf1qr0JFNT60alICJuKbrX8TIRyaazswWOhVRN
flUOBUrSDvpy8BAZz2Dl341l/bt5zxgodLr40rMfI8CVaev2kjhq4gDIbT2AvoU8
CEGHuuVSTz0axbQkf/doVRzoMEjGY5Mi9AOKR4TRs8H+uZyOz2lDdjRBodDz6bQ4
kiiW9/HgOO/QmdsxuukLyyhn28n5mIWOZjIyN5XQeOxIoYFtBTOt55+Kl8LvMsCq
fGn0EL+87v3ZFhn+2ywK0sLuAZpqIiRyBhBVP7JEEkkHg8y0PnN82e4XBz8PdUWQ
h9qyjAG0vB3z4t9vywzzie2JVGtLFxELCVWeIGgG12bd0SK4mD74UwMEwQepX65S
7UJWSWnH9G0lrjyLYMat86qeNck6ctY9quLo763+9Fuf3T3S4/wTYSPDfcsGA7ZW
5CQRLrLvaNM2OphjTwxVlTznkjx0FJc/NJdtnykwMB7k+4e4ffxUdSvKi/5/VMmm
a51LcSgOQ7PltIiCopXBEpCYDEm2UgDGQ3skqfTgvuHi9PBEiYrDUhYLovhybAfW
CzQnd7n1K67TZsJOSS6Yzi/gQYYGN+nAPJvZMKMSRQAnfbTQPYP/GaRjFIGPcPh3
ePtzjYHiDjYKp5/eVLSmX/0gSCecSyV2H0Q6+ZyHWtC9L6043jJaNzRCBfoi7Vhe
HXuq58hj4jeYyMVFUzvXy606dUHqTIU58b5AK8Cu2IddbA+WgCYMMfKg55byd6Lp
HWt6n2crBDhR+QWQm1gmNJ+GaiLS+PxwrhdggUS9b1Q44VZHyqmYP+nHIdPqFB2B
zlmeeYG3Cc04dFxHlho+Os3Hu6iLMO3sc+KHNX3szxuGS70pqfAxMgRv+YQff9LP
Gd3MvO8Kx+RJb+DgkKIwAI4nwTxc3F9sBB7Ju+FL3GlCAadeq7sSg+rZKghpqxQh
SHHm36SyRbqoV0aSMOCVFBotmdm08j46mOjyApk/RG503x6RA+oMx/AwyY2EYdPq
PT8wc6IOUNf+xEMv9grhgmbUHWAfJKRRON7T4KSIT/3SXiB56fDdovAiK5lkiMZd
jm/gZMnZVbYATX9o2y2EfHLwWDuq22sxEJ1HXx+qZ1GG/xg9bjku8avmOszXfN09
DwtlTREX/ad5X3gtfMP++i6NvlUbFIsHYA0h8czMRwQZJ2s+bbcX/g+SXWw/TV8w
SEVBrApSTJI2q51vLqmRRRCX+30cC5YwfiT6xLZ1QRhPvC+k2plwq2dTMz9M99oc
OBBiMVYLd/489PBpTxIQw/d/zXzeYeIqgaJrqiGhH7Ax7k8t9l2NSU3ydZ1WdZ9l
zA7fCOhexsnRkRV0bk/vMPvzkVHGmIE+ZKxp/2iViDNqyo/Q8nirNGIus6Z1UP1B
oPDAZpkjS3CZdMhy3GwUtNgb/umtxJGjsPGmPKZMGp1AZferwJBu5JW+vD+JEazh
6hYzt/SKCD1ftARrHcvQMv0Z/04/qsb+RW6c3ZVrp4TiAwkhTy2awOrR9dXyr42/
M+V0oqcPwOvLLgYaCheZ/NCOCeskMRtom5B1Oa0nwCbdJIAYFJoR41Y3TxFDvjrp
T7UWDxGT/VP7hApHd7KJbuFKP840jnbyZq/wErAxR2VnRMeciZN+IO5rVj5GiKa6
BB9u/FPy4m8Kh+gI7a8LVTleBkxN9CECPixDYT4ttnJXjyclrZmlEMOZLWqNJ9uO
Z7uEFnyT6gL+wSJ7/VJHtUhNJV43cgB7yOLfHIn9gTih/qmQ0nX2rmSDNfiNxsfn
abS/OlQ2yJVyxjIMwsYd0TXBOs9gf+qqifO8fxQoLnnQ1lLk5pPOPRft4n0L+cnQ
1py+leVx+cyCcs4LmjqzhBxTp4ltplIjeP4V2Dwy5DwBK7AEtqDGwOepzix1Fpi0
gIPEz/WIRLV34rF1FhkGFovjO2E6ADi/m1MrDcNRic45RymPkCLmhN00AbXn22yr
A598cszKOFgDmiZEFo7ds5wKZnNj6F904cp1slETKKqO9SWZsWqa+R2umoI4Z4SL
I1kuauQb4WGmTg9dVTxo18ksLU0yTcmG73N7lINHsPDDkPNttusVS/aOnb5fx7+e
BrU3ei3d/1k6SeO+obsoQtUE//08a0VEpKPezFr0dJW09rOUESm9BsAglrINnQTs
JHB5hXqWMymaOveGqyB924VnvjgWrHbGMhE5VRmAR0+3FGF9cbu4icQa0OiyMe0T
QqSoMZ1MnXH8DzS/f1Cn4/zXSrrdpPYEPViDOdqBISYcMLK6Thikg1jb7o0wNMTf
CYqo/+EBo9cY+zvktt07EJ8jaS6jcUjB5ccr+uBkcMuszedFV3yfO0Ju7V0hxZQ9
nxVRRfLETqCucO6CgwCY/JJpVIn+weg+IOljCwEvAlmeQAUyeY8zgfL7CKHnq9vg
gRuKGNX74TIihgvPe00jvqLyrph7Z/kvTDo9lP27lyDarTRtLrEC3X9NX76pmL0m
lTfPFti5nNAfDv8FyEUv0Si06N0322v4ghBLdBzbuEyY+u0wkIiuMAv5PmmakzOh
nOSFuku5WyYHBCYsdZCHeHO1jqxdZXSvFzuWI88u2VOP6lxo7IQgtIB/9KacAb3B
T0CZ7+rzhBttE4/zFCds1ApM8+WsvGt95cGlbBdUnhQvsTpuk8D57Lo3kBCrRxXG
HGF0SgPQk8l738mVaMNMJbJJMGcQZlnaNpdwdg8soUS3I216/kYTrJdNJCmYjcEt
sgUcKiSkunsTy8Vdf7FcccLlSzT6vKQlxi9/PMq+3qkTICUIq2KruAsdWb0PsbcP
4wAizAxk8wyO3vIqoQZ6MzFAcd53FSMr4JifAKUt4fAtWLrn0F+fORuJx7YHt5T1
j+4sIwpDtSviq8r6jk1l+XcfDpTk6AD63BKJyO8oksLQv0MJDbvFMals6e4LJFFa
X9leDobVjW/BbTtcRdwgT3S1L97EF0J5Gzeyrtho5t7d9qbvEqRVYxhuIGKjnDb6
ppG6ps4eOhOhcodTKzbECxerMaaEGqmRNYr8ZM7yQqvTuYWx30ZtnINo3ap4Mkvg
CtAQaPMFktCtyM8draeVXljs6DKypP+tdYJcq1Bb69M/3TvxCHRLvvsyurLmPe79
svqjNjCo+I9Xn92UYy3hLt4b0/xuKCb14LCEmf0Fpt5UJwWI7rgw+Ii4LDj1FZ4T
0fa/ZEARjBGGq0VC/wxYnOk3dqHpTE/U946T9Ggjxl3G+LUg/ISAY4fqXdytrVwg
eMnLsFVWIUXckElTeQBxNELP/kubbicc8e7pT3D4t9nojCKorVVnXHqOcylueO2Y
iG0WOZbSt2YoIfQVNy7OkNFjtQfidzubSOgyJAwQrr5T6oQgOnfwg3jbQTAS8gI1
e8E+iPGstuBQR98GgDi/rnJymTro2AxmZjXmAQoO1qMxT7iApvj2m9PfCtvw2lvy
/NY/do4S35q1qnNqSk8fxnG/z20pnEvviVabdl1D1/hjv4g6sYKmuGlaCTZjprYd
vr/IP48PaaRcC9kTDxaVuoPHeXqjSlsAb+BtxKhksgYzpi8YnacpcUy8lafOJx4/
nuFexTTlX0O0k36vIp84YDAzTbtW7ynDcBw0jnuctixj2YKTy7x91zRcrA9kGmNv
f8dey/IE1jGw3Bh0991j9a4zzfhqefs34DGz0FlqRWCnvhUFBTVPrDwAzepsu3Te
E54s7U1r0P3StvCFSDMm4Vap5zSwEWup8tZo71NAVMkZwkB8kqKEQUU+xDvQdaVV
yGOHyIbyWL6SIGdwLGk6bPvI3dn9NZzjusqNCaGXlCUmXlgj9zBih6osOzj8KhCQ
ZPhaVF6fLoP18Zm8w354nRc5yZU0iolPjPNJl7pTUYya6o45VPROgQBVbYCmFe4S
FIhVrqwZg6wGgCbxPU8CFotTgB/kqhpxiW41AvRDk640jFPgDurEyuQFAc7O4KHz
LPMGhgbAPAnzI2ohIjb5ur0Rlt42MibPdgzU+v4w8/un80lYENtV9fSfmjmWCEIx
DU1JpNX7DkbtjAc+9yY5URGC3VW6Z0zPWot7c1Y0mKzKMsK08TtFYNBj8ORe4FCB
3QfNomk31Mv7cQpYA5rEnrwU3K1WKXBFrS0vWwCc4prBveZkUMjvNHn2vg7DZhWO
QDc0aB/VOIv7E5pNKI0TjcupauTGKlArZWyDLBJZeUS+nHiN3GM6lDK9ROJx4YsT
tkX+8g/wdtudLZKhqL1JP32XKUnvRt63Vickh9iekY8PQXHK011ipXyzpN9NBDn8
amDui8ZSML/BvBrXt2VGxw0W8yLwfzLlxfspI5g5vXLxl8bpVT/klzwswWzN594k
K5UXX4lnCMKTjyWTqfjnYcnml4Ufi2aJ08V4V532+Rfc4QdYjAUupeYKobfdfQFc
glyJU8bBoTZaHbAPdem1r/euYpwtqvqtmhZzaGWTMXZFXkCgNl3IQ5Mjqr/kZ//T
HyB9kA7spHRxfLCBiitumYhqHG4WyWUri8T6VOSRzBe+fzaI1FnLNO4xU3dSTjHU
zd23IkAazKXDqScRXV4EdhDCEEtBD/sIUPaVTFUdVAAXzlRTfC1iVS9QAuCZjgOf
hF2PDnUGLIQAq/sBwRIgQ9aTWMfh6zhtSA8iXa7RzBqu0T4g+wGieSVECXRZ/Uqg
ZmpTYzZIMbLrVpHS4mcKzYH0D3NUa5anEB9LyWKBoesP51ho/uLxEsj0Kv9bdoHl
i0aKkt8MgzuJ/dW2o2/22RWgkwf1wzhAYVC5f3XFJOhq7oPy0YVUtk8y+dO7vlBW
Z7U4Apw4lpuSBmbg78aZXAvHc7yngGI1bomCVYTgmhPw24gGAc64QrmSC1eWuYJg
tacW2FvQ+/DykcHWRiMNqOYYN/Gw7/f4CGof+jlOpehhVjtmISCo52r8FrGC9GVt
hFL5ypMIMAaQU2L0hJUJxWhwFHAAdGm2M5u7cgq+e3xmH0V67HlaMdQ+F4L1GRdp
1IPhwEsazfVWjVHNwdE1osZoh+ixrAVsp9DvPnC5pBLSLgvTtWdstWfS3xw7Wboc
Wmt79Ccb37fxix4s8dFexr+I3ULrG/u8vgwK/sEp2CN/zoNFMgoi8Xh+GmSXVj+3
Wb3qmxQFvA52bWwyxoKmK2aUp7ibMLAujIDv4+9pib060rLamTB/aWYprdKa8XQI
FI1FecXawUsIQof81Fk0K6ftIHrdhc9IKqYfvhpVACS7pl/FWx8m5AmDzUUjtsfz
KOwJGMa56CUM2R9o5pHhiwnL7eDEzxxpSXfpuv6AzE/yc+1Xa5mU9HLrx3E65miV
gnkueFbS4XV7HBBf/egFx3oegWfCFA9c51tuLbiR+0Mpx88xzDC/QbmR3n7FBir1
4QiAsClythm30pYKbUg5LLq0Jq2FqP2AixMN4HWr15gHKDNGjtAwReNS95eU0eUz
uMuT8zc89YM2uLNRTzxjWKyp2An8z3dAxZUO1iJPXQEvlVQFhUNipnInn4wUsdTy
c6UqbUti/jKaWV18U5lWr44KXkIEj2KmqMRCBD2WBHCPyyzjwLJ8EQe/aARuyWrm
34aLArb0NssPcGc0IwLCr+uswuVlKKHhLLyKw51hUnBeHK1XccWiDXrKQvFHSfLD
F8XXusgvFgaMfPt1RuLH9ERjqIvA5tvUCF0c4sjtEj0JmpR481LlLkaH6RMzhpFv
r8KnqLGTVJD/+6bBziFlWrUFrFiJzW4CI7tU1F2KnMnmk1nqT9Mgn24QoCRnhG3c
lDqBDQL2+svqDORnPg+RbhO5iqDPtNTJlfq8rsC0wDpCWrRksW9u/LD8ty24hPKS
GHpbLtXvrGsbObj4z/9GWv6xMwimRAO0E+vO2QHh/zV8jVBvNID3cJ/DOxjuHHpG
aDJIx/EYapBmb3yCkqqJFT0hmQPUaGpvM/iHJ3ub80RmOxKmZHDdsKmbFlCUSHRX
5rbEGfEG9cSCkzYOnHk8O99baNVLeXsk/GJ1imc8gFllAJjZFAII6XsS4R4h4oBZ
ONv3b3AmkjxXlN1puNqBy2UbpKNlQP9Nua18sAm1JIJZB86cDP6uzYz/c4ctbEpu
sDmj4+KQ49E0RD67wD0qAzRUkIOp13u7UqdiZ9fXApkTd480e1i3UL1wpNkQ35iD
EgFH3N2Kvx8veJqsNF48RQ/9vJrhvsWqLnp03XaD/tv4x6fMhch5w0XB8pM8+Mib
hfWhXzTVnEpR+2idsb7mbua8Ua0FE9bG6pBh2HadhJfwB06aG9dUqiWMrLNZX3IZ
BStn26b6UWx5WRNCWYgnXIRypMCx0i4VuLrnQxlhcB9IxEzRfyz8u1IWfolikCam
k6rYkqu49hal5i4B+Yj88Qm9qaggh7jEN71dnmUxGAZOjO6m5t3Bje0jr/yfwL8R
/pz6mAnE5fklQ8jHde1/JbtNVgjctB58XrAQIxpf8V9gsMM38nWJYnfZGo/B9OZK
CnuKjqGNxFcixXT5D1Gaej/T5dvBfHd92HKhcUVvKfpji9Q6JGU+JXDCPAQYSVYl
lZWvBgZfyhZCoiKI5jQ8EdHBbxJ2XNrfHTFRF0Vlu8zwMhUH3Lr7UjQOULnrlaKG
4YA5s14o8aUq/vdin/6pbZPkg+USrw5yfAOyAM8sG4zzGs+KRkMEeSmhrQlLUdGh
ZCnh0oiL3Ew0Gzb/dYi5alZYgUFMvqyon7FsNl3O7rNOca6EpruOu1CbmcBVa8OD
gr94FMvDz7RiI0vOyY6kBmh0idfR35h18VM91b5Q0A+TjmDPHOhuScSG3hfPkQZo
OdDSRxfP0iFvpM/Wk/P4vdVo5UOqxJFftTUXUkNciB8cFg9hON6pqg/tj8PA5OCI
2FZvrjnxA3eD0eER+LRxUmTC70SgyFCAosBKD0srUsp1SJtElqayNY0oEbaJa3Ys
efhgZP3KNXZUN92HOkuxDx/x8M2eotYq8+O8imhxN+RXVRMS+vlYFUwJA8RK94A8
zK/3UUEbFAjYqU+fd5L1nndzR9AABGLkUNrjkPqnLQQdNuhptH2j6Jfwb/ddtVCB
0PPtPIaWX1FuWZJC+UO1CH2DZZZqLkmFfbUS4hiCyXvUocStdfIP+b7i9+bQKtSr
VWhpXgg2mYKCIMSI7eN0LlXExxgGRSq3L/paI+sTD0VwPeqJZeKFk5QwiGMA8w1t
kGYNiblLKWCDZyVR2376u/dofHr6Akojs5v4SkYyzUQea8Q1Hysoz/DKLSQTCK31
bx3JIEfTnFKQSn3NkvyeEEMHAf+nZlmUP0/FbwTVAqOD5FFHKlyUye+tmZeMz1ni
1fi6GJWdGPhP8zCVuZzlG3geFaUkVim/X94XTjc/H1QG9EFCjWLanPumRl+YdU/g
ivZ31NZJT02a1dcG4MC0mRrSHhjYJcRvp6rrEfOgTALrls8EzHjSRHSi0oedh7Ax
1SW9JCEydRCzWLXyfhO09G4kIirtgjwZ8FjIzVF8qWj/mXkGzkGu4yTktuSIlfvW
nYkvNthWPUiWaxSbD8ADZcb6UyjHLnbpD0tSggPKbQQ0oyz/UE0adbwCFJoLcVO1
+NVA3yo0wyCEP1Fnv6RBPD5o/21ChlRSPPfDhX+Tw9xgASPOY4PHBZxTfoXCnG4t
XtdKc36csZTuSToIXG6kjX+9gH1MyooAVDptKQwUA0uAy8BREmKz7LlqIbGCgkt2
stx9YYd5iVpqBgZ2tHI6SJHdvOpCbSWoOrZBeHUhlTzznG2tb7HG/3ILNOjSFsDN
XPaOiTxTOeADZie+cf0glf3lkFeJB0w0ZcJTRDAk2+1zNVP3akRsJFrGCRvZ71r6
5Iw/R4Yh2y6LHtkAN/s5/7+s1JRG6VRDJoEJ3dJ74Iurpc23K9TbDyxzCq79FPSO
lWVn7vBJjzIkRXXGcyUWo+eCAl4GsJbMefwayoQNEawWjmWZweSsYZFyo/cZClnu
EBzhd/oUVLzpgm9G3hE0OqxL4vz+2/K8khPdzwoRuXbGQrm33wKiFSwN0n0BnCK4
+PQ51KXz40y146dCTTE6JAxfpS57u3SPj6af6p7GGhQZlbfpyTVut2OWRcvXPinU
RKHSJULYSA+S84TkbQtfDQByiUiJOwPB5sMgF2sQNqCWP1g41ekeLWnAFgz6XJRv
io/TVXgxwhdXx1yoafa3SzSlUox+VfyqPkcVlLH+F3uV6iYmstLHOOdIANDZnN9/
4K3KZuxwCAejKtDHcEiwwAqfapGhQopiqEqseaZe7loiimZv27QU7SRXq3Y3Pe0r
FeraR+AUqucjLPWacFfwPb4vid+wG+V8oBCODO9HRiDjxzakay5kxRDHHo/WMSYx
reMbPOGrDZSUTlIQGyRZBWiqn8xUXKVY4J1R8ZTNWTakH1U1uKOBPlZbf1ijFTW2
VxHHqe9zU3Xx6mZXJFvh9gLaeYvcloGVsMPZydvC+XOF+XGIIb9x+xK/SlahC0Fc
axSEAMnYuRzUtQxqs39ormTBHOsDyUY2KfFDfWYuhNHYI1R7cZAkywuntiWuBCKR
tkeA9k9CNC0WktXUvYdgDVWWyLott0zJyhZskEyUhUzwMOuqjwhGzWTr/DR91qp/
wGArY00199lMT52jyUEl6v86Wf9ShSMCwPOhgsfwTlIVSZIek9I2NtHW80QpMeJh
yVRltNwovMOelXRoU5z1E1hVJcPAsJANQ7/JVTNIS4OaQJFvbWGbuSyIGrcGFwUV
SJH15hE2SHLS27UGAEbDUZXgCpF4+4PRSqd8JYMOMPmIF1zCNqm7131HRtxLysX7
WM3u5KW3C9GH4nC0OKsR9wO9TR5TOQCAZJnSsJyc/7W9mEhYCRTLKlWoNsaFRDRM
/CzXBRn1rBJf0mks1bMudAgckozUj63lAZMpIHAi4bhL5jDNqwlsPvCDX012lvv1
5K4SZF4BTHeqceMq9yzpSCtUAy3z7g+2Qz3WckiT7AhDREfXbR+fyrFBMdBzIkcq
ygAkwts0AZSrvZ5kAR6QApCSGRkb8Cu7zbeOyfus9lY8ICTK/2CZILL78ZM78GL8
Xj4O/KihSVzNu9gCNUuuGE+8QfeiIYSbc4kX73DyvsOpYCgNQVeC3/iv2WT9+goU
nJUL4vhsaQCILFPrY9qjjH2AjFFwVWwMs/jRcJXpKD0kH+nrmHXl4lmT1te7FZEx
zNXn/GgCv0qeAyFZ8bJqr+NrgkhYkE4F9LSkgvBNIAvxW2VYAHMPmyUAhixw90nZ
aNpeNQwujS8tWJKJZ1yNl7kaawr1AiSbPaqdGn68rO31H70OPQI8c0YgcHr1/e7Q
KKYkhiGAGfOUgKZOT2iGM901jnvdIK6ZJfbY5zBLQWpuoM9sot06THnfw1zaRP0W
cVPMVA0UGzMnzO33hOc63roPgMasrxwPNkqW3maVS+rX6z1LWmv/3OZklq3Ds4ui
tP/H3dUyMqrXpebSoDlBuTTD3/xZkB5zVlzkH15Uk2by/k0hGpQbgeCVaXl92NBs
fec2akJEpmM0dgvQAVP83UsUsfI57rg385tcNUPGwDCBAM1YTrpMF1xh9T/phy6/
LoPokROk5sG6GFle0SVPwqbzyLAF0CiVP82eoTX0p2aL2bnFI7nC5LyXwSIitpJ0
t0cLd6wziCVtAMjl9Lg3y9McG71q0/Xs2cuFki/x9hJ//An/QTgebt5ugM9gmiQ4
aEQJ6p/3uaRbZCGGf1OxW3m9/rlwNdhiyV1BpxnukzMuPZUzoFDlL8MwvATYDnjn
sJSxsSXqbaW2jpWhMobn+xJmWm8N/U0wBYAbegXmVsHGVt7SzIbHzgBt2AWkza7n
nAHC746ibNTSPBf2RbcfEazn0b+qBrDFoLm9R2ZvAWTCNgHnOUq5uGAGo+ptzxgs
lGUBoEXtWQLW5eofH9cPC1N+a2LLv+9mkt3ua7kO0huyYRmHrBfMPD1l/EeHeqE0
vqVGuacCcbhMeLdOVi5x4ZxEW5a1tetLujdKJhgwztBwl98JSSMNRO6a2VFqI4jX
OTS6y4Yioa1xDAHdhdBVnz9zpic52ykl208Qr8yOqPgRW/vgAv0eo2ikM4VOFBE6
86A2Ltto9ha2mi8N53am6ascpn6mX0nxyQiAO3YcDwHwUpUfY0lbz8iWRdh3ZwP+
2CN7gRnX1i/zXSP6sSLVX8gf4ncHZpoWeHX/LwP1YcTtgjAShNiFZueYqOadAeX+
iBO/cv+rvCg0fYzVGPiyC4FWt3aFIc2KFOUib4wJoKriIaTn6WwJOO8MRcHj4X/t
TPHEA4lEWV3YnY2hPkYAOfpDcJ5zb9cZua+/f02ec3/FRQv4NaMmYm+leN/dMksf
5FJ4s98PzfXmV5aNLRSpNlLQkGq9HYp35SPqAIzu1sCaXSJfAjEEDWzZAcn4Nywt
M/0mI9qv/szo4jebKUZ0MVYjMF13FDmyKFuEgEJGWzOhIjFdopeP7rGkvDCuKZqi
ofHhI7xlMAN0scIWmFgsJu1h44xQrsTEiXXdhIQ/Q41YFZfUbpH796fSvzGcKPjt
eTQnPd7PdE5K4uOyy04SQdtYodF9gaPk+mWvbVF1aMOVL/IgnlFDc+/AYF0fCwmH
W4Ql/+Ljj6U2rtx65hynFKA5gkeYmxnWCxR6/uwJ0fi9BobO4NK0tMCQuqf2k7zF
9yx/hnQS7iLvL5zflU21AsfW8hMlk22W7ztDsCihkNjFMcqhFYDmGbOa5qpeIJhQ
jEpg7toAuDuwIdX/vtJLs5Ke4uH+aB2g56HegOkeHQvvFkWs28Gli4UOCSJYngCu
6vhDLIGHE1LUnRoFSjAv05Iwlz+IqeZkv6ZCj8mWlLeykeu2zjQgbO2UVh67jEYf
gAcAKihfVsxLjZhDfKwhOnY8opJ4SaKByl1mn75EXtU34I889+pFG728jrmZCd00
d5ntdVNtzcH+7E5FV27b+7gaJUGz2G/iXlcB/T5/aOM+gmSltFGeyGkOAFvEm2VI
cKiDJ8AwRC3oHvJ68k6r2bxpRTdU4qCTjYTBS3/aMOPzdig3hEIQA8mGrIhhz7Ta
X1WfoleY1oOKWSZhqV3Ev4W/fGGPfeDR4zv9P5dnD5drY+rmT1Apvwy7Ye7CuLqA
viycLZXLhwsOBBypYdh2ChpfTcqSdI0REKbOuqMaa+GH7R9CtrBePMFQMztwxGig
69RG5JHFKKMQhAyMIxcEXZxYx2PtOZS9Mfowau4codWx/14+HFrNaTSojNz++9N6
VqX5ID8iNq7t7aq3XT9BKsAIMYvTizb6B1l8JibpM4czLN8xStundeqMVAs7YSDA
jMHogHnn0nB8eeupEcsdyF2Cmi8faemroLmqYOe0AY9d/IaDWlg8AtJcyFk/qJTb
yg5e9ECnNN+KDOymBfRC4GRNIA59AOXy2OwKcRQAaovj/AaeDuexK02p37BTDGo/
rJNUoTVcQkqBDdAycYCX7NF13nKMylfvngaGxHYnUEoKP6aoNgPpP3/OfEPcKpvT
ufwdRQRnEvKSZLYBjAYP7XmPXLlgqebaMdYYyZwDDhkLDLCpIy+yqmPCx62yS/18
EcRLr2U8ozjKLl+VbmoWZ2GWNsxjVz4lZ4kXRjp8TVgpENL871j/5ZhHRiX7lOBn
IGi6aQQ7wt28kGSucaGLyKavwizCzUubgsyIFI/Ovxq3H+rom+S6VNjv3FOnhCVI
0HxLZUWpka1wcmwmUy69n+iXrFNCC72yI18cHe7wMvl3/E2+OwOp4mXqLoUqDQPe
LKrnCpv97abXqALCj1mbk155iH/8s2mBK9zNidvzmLysEvLOZoV8H1oiQmjaIiab
1Ry7vK4ucJsX3FxnR2WfU1rj+2FqZ82ZDK2Q7YPnW7eZrGdBCT//Kogc7VmlSE0d
vDClGJooxtH9UFH+2kcgWUHcuVaYpmCIsKZd6zPRwd1VXG/yRM8QYJnbn+PswtVi
cmmcCGVvz0mu5hoYFgfHSNrigodJwmVZYzt+8hjIMsVW3TZEtnhjBx+YiCd7MQDn
5X0dUq2rIJ/92oUJF1y7Yaq04N7HLnL3+lrlQOIv2/d9l6nMNIH+Afc2Q12Jk513
p4+MqAyc5CV3e9EmjEvypvQlNA3jAzr27XwGNfvsVS2wLJl//1O0aJ7UxAd75Q5+
SbZlDv2WEoQCd2UainBtiY03tqMKSnDUQEOQYm+emVVKCbrQah2JPwDHWF5HBeJS
iD9LDbY5CNN2HWzmSqjfxyY8tbbfHqktj/LVUTVuksQQlebuKRA1ISU3upNZNQGh
SGo9yLKM54qLzfVkoS8bVaDgMBG3opCg3l04g74MRPcOFfb2CslU6SKemXUCpkM7
tffDZ1cLLR0aV5rNRvgZfTL8t4ZxOHP5sR/ekHDsbiBFphiOvjH33xbX5lhOmfgU
DqvoxhoQReiIoXB5laurqtQXt+9FbfFW12OdjJ2p/RKC+8F0qJSF5ojh610/96IE
H6TvPHqNvvjdB3N0czk9v4duuHM4G8WvcqBTVcIimZMB53uF71dpihde/j8Zo6d4
pClz5FYebSxg1Wyo+Ny5J/IbrQ1pKiEo+2y7Tuvj44F6ZUqx/ZstTT/Em9uotBhG
FPodluzcCLMCodIt21Gl4ceCs0kXW30mvJ7H05+OMtq9dR6jEF+dnSabqIfZlmBI
m6z2Ggl6oZqNmafYTFwbIUKQ/6MLsLFhYwwVzddu1mJGMA9d5zgAVJCIYxizLKRU
b0O8ihaEG7zVnhrwkUWsHn1pyjXqGyukMCtTbsgncRddSEAxgVIs3dXkhwKCEVpC
T9tNWKLApf/y7G79ALDMd4/IL9Apc1gKRLkNpT+oD474K2QmU45x2jgsHGvMV1QT
d2ceyAGogkbBFFxWv7qrNknMizSyTMF3kaVrP4pTolAZ8qAfEeR5LkBlKdZVDi8Y
2IQ0Pgta2oK2aJlI0Ygs5pqKZuaMNv2Yeksm4sMcgL826LI/vrK+4RWho/LSRKm+
rmHMRRzGdkuLe9srNX1MugnqAcBO5f9Xe8X0kAuruPzq1enea9GdZp58rfvYYU59
l3mehjW0tBL70O8sAPUuLMApWHjQHIsQmyNX+teMdEdXVfY9mrEwSnFOPWBj9w5t
TiWyF/v02y8NAjLTuqQ/555aDW5j+ZXbCT8GwP0cgOfAczT+FYm92Qi6v1Dza800
JLneC+49Nx/5rVhFkgPFI3X2xwUUnHwOU5JBesIRi+ozBqvBAiJFlUU3MHAEcZQ2
uCaikdx0lelB3qWjn+txu7EzELMSf60uBPpLG1wPB3jtndUxvRkI/RMbWH6q19u3
Q8OcFNXZUczdHpJAtI3tOeLBFyAavTN2UAnTtFj/TEc/S8bBPrAB2jzj8UdN56VX
DWJiCjyVYJl2fu/TZOmWfY7z+m8CxDtRI572ypk8/V0nzG6VZySSC+5ZTNog8RJD
Uaw7PepaSBq6mt7uZPYcJGi3I4Zcn93xa2y7JxqHVkidBdi40wkev+92MtZcfkLw
Ii4E+/zuGG/e/ouThChqA59kxaiGoErJxZTofzJq7NsNkgU6Y6gUwrvcOQAyfSvK
8Y8TwhEAsQ0YOg6fFglLAqQSZqkc1rQI5YSVqMI0mkHEsIte3k2jZpgU1KrJIzk9
Jih6qeqLcb2gmatUWInWVr+N39X9fsZV623MputT19fD9wBkeWCYHHFlv2BEHwDi
tWxwZY8mD7TYVB840fxtT+rFglYMsxXVUEIhtY9W/o7GvF/4KlR4xLIK4MfmLRsA
T4NDfjnkYOOdTaHGdhlAwLM237h+BNSz2LC0J4rEgOZ170lOxY8Jv25og6IiVamH
NWgbCcXq66nnGn4LF/BkS0YnAgykCFTXvGg99Zgu9cB5fyo8ejRunjRblYtoCo/U
aRweLInkyZymHHaTNmWHmh2e2c+F+uT8fa1bk0u1bUlSF1OgzXrEPNPlDc/CJN3n
WQp9hHq546Qz6ALutZ2aIhCJ+wJnY8yBfn+/LFHmS/O5QuKBj8Eq1GU94k3JNbgN
84epwDWAk/Int7pU/LjPEg6cpLsar0cyoW0hYyFC7VAVDwLqUTqJ7UAaBmRDlPCY
/ZlbqIiSViKwVdEo9qKgwavudmeOffP/gJ4DHaFYvjtvGfo9ce8/lUhByfStStRZ
Xo9WmbDU396l/sWpB4+nQkHojamItRjRGC4tFNzeyzx7Av7vcFiZ5fYAG9buFQc9
LgAdFMtc9WpC9p4xyHMg7Ij8T4/CrF9leP+BMDyqAndsiSPHLAVlmkYWWRkKzGOi
5fZS104+QCaIZRNkh7qhvpNNE0pGVLTFK3R7uQIGemTKzjRpofxjd8xLXDLTp4Cj
nak6cLYVozXaOrqUK65ofnpvyjRuXwZ8mwdIXlPRlOFDyZTrlhuR7Sn6Ez+hmuL6
kdUTDyYlxYDNfOXMrKQrb/tVmh3BVMp1C/Nt/SeZMdOOQa4JXIzLqaoq6kZfzG+T
um77nvz1luH4yOH+7RbGO6IulqEhcM+gBiYP9Qfbu+asb6hFtc0/D5yctcYld1wz
dJ0VK4HgJTggikMeer0QilHd5OQJGG1gtaD9wHhjI51sRVKwRAmmgdOJhsAoql4H
6gaqlpBxvee2PKkv6nJrQb8wpSvjnSbPE5JbM13lBo+ovMz/xaWbf5qkjV3VDQEa
3WaRGFWAUFQDWYVGzuXGCqBtrBiqWsVpmzxGRPgNBDP4i2VI6UwrG2tVLDZg6FA+
jO+/yK0SHJGYx0dnEduPr8So+F3JI1I7cdzqv3+nehJ3T7xXi84ZiWc99YMbt2Tx
AvF5CbGIXGXDTc93Bw56UedFMRNuN+JkxVsfhZoaOe9J+XF7We6Td7/ufb77WwSY
cEa2SXdJqnn1uwzw/QAzUHs5LzpqTSo/wBCjPZt364IRtcbmWFd46zuh9VmAv7lV
SQisXpFHGdz+Qbff4fYVrJK6tcoTXJJj6Cr19+gF10blgrbspbrckW32nEvR1rmj
N/GDlIPvU/wyGBQLgdsf58QHtdPgjDl2Z1UdWun7B0Bhu56P7lDSlViTlyLrGbHJ
0H4qweSnp2XFkw5WP7M6rL2sp1C9QafIambn6qVwQSFMuXhPDwe6fmQMivWT/EHm
BKVjrY1OWgGc3SlofNEMJWmazgys9dcsTzrLq/J9xepgjo7T+Cc8Ry/DBOSS75Ok
QBKJd3ak838/ywpIn/+sBl1S2z3N9igA6rNiOl4eHs4FuS11ia9Q402DVgAWEABS
ASdy91oTRUcfm7W/axTKakkj9cQvTz5wYjzW28UmxfQUM+8+RF2laHBveh/HdF/W
pBLVxxn7wHqUK2yRyvS4T03RJaPIb21KFx8G/qiUgBG4E0HR/UrWy6RYp0CKt5ra
XI0f1XGCgiytOclqrON0FEoBbD4K7C+MXyAgomCX+aF5oru98Fhy46+9URu/wh2D
ErA8YrqR9ry6CxurN6t03vbiErhajCf+wXWo6QoVzFUO4ipNqF1UEl9JWx1B6W5g
DF4Gg+YEBy3iC1vPiFCT+6cmXEZzJmKA1mL8DcQLFaGsfnV2sjiMoQMAzQyQTnL8
oN/fhEFyrahQ0Y9J+D0tmi8BmOzJTU5vo1v3uzXXEH+sEi9+jO8YBaDhUy2L2ran
tY0nlHTE+BHwc4Dx5FF3hamlsrinnGRXzhLg9+K+gNfZbvsManH+xTP84t7vElH9
nMiz0y9ICqJx4tC5R6OCG9WYBW30mUmrP/0YFH/CtPxb0HdWO8Uynqc6wJXPE5ix
srLHIaFpznYeTPVM8S+TalqeqEEddreQGc8IKfMRY67xt8hj5tcj1MMHqP8CWB4X
75i4SOhkGCNSPWz7LKoVwrOepeJrTFL+EaoUozp4zzb5zwVu5fbuUUUBGDwrJjWw
D+qDzKPskRONHo6trZoo4O4NO19ztOVOQ/NhHaseC+RAN9OmA5VS8v5lfVzRKtca
cpzLm/xwDlStW5oU9iVKNrnqHxCImJZBHXViA9IvRyEZ46vhheP9WPlKGAuC+++I
W3PdAtMa+0DscyUUXWT/nNKxC5Pg3bjh3o+DWyrRceHjnWOcNqq8eBl/j/8vVfT3
RZ4XDID7Jri+uOIyDw64WXzd8GennVPXlFxycOxfNWHjrOzPycLZ9VCKnIQfWcw6
5bY4wVeqiimjiWBjI4PgfmWeCMOhGzXA/CiRc+HNlZBM5wUQ1y00N1zq5RMzyuBz
UfnWTlJZgBUIkJbQVTNxZyV/kpxNuk6fnwnLo7wqs2m5q7n5fE9o9RlpxoIRwdWO
//mhmNVoF689Y3TAGHWuAmYHIhk6kuWYawXMGvd4vBkzVNjJR19aL7OUeVA0bp5c
QonBu1RdZgx+xPXu47Cb5DOulKiyUYLq8Fa9fOXLlmbQyhnUqz5VU5SwwOiWY8mT
dT5UFlpYdk5p3iHXv5OJyIb9neL+5JdIUR4Fj3mRUgM/OnncylQm/NeByAuvZpt4
Ql90dknhq7M9KvtxtfY2oc++7gM+7QDGw8EuEm+V7A+ejlXV3C4RvM9r+sMmdsFF
X3oSarnJ2hU2NJqoz2MtyxfpeQ95PArbWBTNQP8+jc9RUAIVMifvO23p8mdWt4HE
R38YayebDCP3BGOdeQWgG5d2Ts/LRIxmHQ7BJGXa2PTrDuZrsIjbafmqdSVkLgSf
hNtBOjEH9TjkS0Xuo+Z8lR/RnPgLAfR5pkJrwfVLglt2DqXCvw4NaVpG+dELqQZ3
CST80Ias/PXVQ84GEHlFuq/YoxewRFBsjZrU4R85RM+voToi41NXXrfZOVH5EfnF
NWdsFPPWe2llBibAMf5zLzpapVr2nObAOZr5dAi7KG9ksWFb64XE/DvfECERV/2E
aGCEu0RWhc3tVgDNA5AlbA8mIMjgJDAkn93arX7ibUafpxVQVs6fEyd9WNKujtwy
HsTTffABcq+uwXrHaVeDwOBau/MK5VYU5CC4e0ip9tYAkGieVBoTV2tGRdhBbuTW
OYxwJt/3KiIUOnarvNiB0YDhXUnwgcHDhsbR2skkoJk2nvphgWOWiwxQcBkMLJe5
69zBXiuvbed1dUnMxUnRLE7DmFFajR2gNGXByxjO7JYihO4T86KmdDOVgES+VpcP
3n0yBUqh2SeXiAPLK96jLIxfKP+ByGarR6/Tj5uENqcq+XDdcW6ati9QzakfwGuk
5KclOuhQwaRMPPeSc1prPVzbxRaN/tUoChtibLYcbRYK1wZvseNJUZtF8JFXn2fM
Ea2D4sNdI3+iB4hCK3Pr3aoYO7Ayjxnbgu0MHs9bLeQkcw08nHZxW6ZIddJ/FwbT
iBkXW6EGQqp0MBWrfTsb0dBzfNANnyxrURFHdwbWaygbUQTBxkXvrMdQu7IO0KlI
tL5SUV7te3nfrOs91EAyrIembpGElgHu6Diqj8vTsjpB2elT35fOpQHsw/VcPbln
KoIwTmTzEviZae6hnfdlW4wD40LQF0ydRFUnwD5osQ0UMO3REpMYCnwqzwZp04JF
nSAgo7tigio4sVOwTc3nLOdJzNbim40kydzZBiwUW0azVk1uyRYf89UBMmiWSGr3
2MnoBELZwXzL8L46J5bcCfuJrXEjGS+iu44UF0BJHvayZhuNNyMcHaWpuZAIaWzN
PyYE52Og64eXnFNab9bTNKKDOApHYGmuLxnWau0sRo/7zNoSUbzVlgSpHqBftb6p
V7mM4keO8hj5FZqOEhMmjRSzYZ91EdvwUYbjUH1za8vpfhv4xybauwCpkZSksqK/
0HzoViwtn7+oMsgXiwwVGALf6P8i5cu9+6u3/f6OdZyfvwVLd/MIoGZAeNM3Kr2N
uLNSPol9WLApyaDlYKcFt7FVniAbhz5QPU0jhZeHEbOjdevFuSy4O5T8CHbZznXw
iGzNDMkprSfnLxx2gawC7p8F+L08iqUyFHGag/8VUR9O7u8myl+PBtIBskk2D2lL
kOopIqVgGZ8rAwUbmIUWPYhAqkh8om/VfINXM8OiGaC4fUzRwoPCIYy7N1RKaKTL
NqJgM/4yqJ3rlc8u/HEBFzqBBGz82CxEqTu2tWKalE+nuh9Jyp9vGmIHj7uC35p0
5DbnDu7tYSsAVec/AE/Ubme6pG5Uqza4889cpskr+vzPpqR+VU1N01xYm3cbXM3h
ISTh9ev7G2x199nMPbUVqcRyCEa5pltrB5Fxm+qH0OkTpYTiWrK4dd17xUeQSXBi
wo1jqUFEuRl7w/X/S2qlrtFOEhre7IRrBjye6vNhkrNzqUwet010Rly7f3VwuGe4
ku+2BstEJBj63V3uA+0NRmb59573amwISnb7MWvqJfEaA+Mu5Cv73bMsMIbPfXO0
pM2/08D18fbQ+jKF2URxPjEsFW3bcHApakVrtxbaTSOpj5azyl9yCjl3ppCg7IMB
k/lAEEELlq2nczkMwY8YZDtjT1K9soVHeqgNCe98aHcSvttRMjgyUWAI94Wo6DZ6
yaTAAiQyl4z0SLJuT7IUpPbxRTH+uG4FBUJOotQFxXfAOsbBWUp2n4Y9ZKB5YPbG
Gc+t1QliTZpNUjGJZIfYOY+qXS9634XEb+vZcN0PVJMqkCue9ASPeGeNQGAsjqUk
Y5uq3Rdwgkt3ds/esQKPUDEy0uVUKNu8RazCjIca/Rvr0492gJIdMa3nfX2V1aTA
Pofe7YptpgoliwdS20i8o6ziD66stpVYs41NalOYXPDdwDafwRqZdbgFHmReb+Nl
70E5Z+TeWDWOwUzRH6QP5xzfo5cHrP0ny0vuK9u4Z+qrMz+ChoL+Pn4kb2cXO+U1
NXcjA3Zao8Pt+zaPWYHXp9bZDA4qb9jmqthSRWp1P6o+tl2MP6jrP97emlO1+0LU
kYIegoQ7cZAk2xXkmjcKoLgw3k58RXMRFusYr85E4zoL9yfEQTwhQ31H3tI8g8h2
9cJKqISuno3EXxYKC9lwuuNQG4R3RuMhCeVbFDhMAGkyA0eeKsJ/w4k+ilSYsP66
iS370MAk6eNFXlYSOH+QtRq/B/Wm7mKtn4YdrxXCXl3XbDf82NIw/xC6Hhn9lql4
l3tFqZyXWArMLj+YzyZjeMgqOrCO8pwTng5llvNyXyhRkJe9iwKuQgYZNIh9FJh2
Nt8/PvlTLICg0DdnCxmKXvfUnqX5B/M7e621KrIi2YafpBZsPLzLG2fZ/Ig0cTAK
vU8muptU5VNm6YaCIJuEgTuX/sFqrup8rqQW9I0rXMgwKSDXRJWuh0zAr6G4/2t1
ZjLtCuYU3AQF6A6zZxhQkwC+2QbG14eb5IvIkvuwfpT0UIl6KzzUqdaCRv68qxto
CicIeqoQRnd48fxVxzbdIxCOSk+PUa95gJm7ZPGofnuwLfOLx9suOPzb/gkxFUiv
/dZx9O9mOINFzQ9qXvWGtmAK9rJED9GysSzL8LYw3YuRXxPQ4ynGTtFFfDDzHBZz
j1KHcil9dvkTaktwmG0CinYLiyLK3d4IoiOskqTc0r3W5okVhptj0vBU/C3Y1p6B
pVGcmUGZ77UTbltbcT7z/26S4cRKimLNgmvoDsIYNLr9Wo7KE8JkuU3Gz3I2XeWo
bqiyFCYQmQHUd659Ya1HW1TU1QfJ6v33j8zzlZXIQ00XrNekMvlVy+LZeH50OnPb
CvydXkkG5eQLZzK7vAkq/IYJRL0J3mq68rUBKYKI2+IGkocEfHyekEHnjYjT3C0/
5KQ/S39u9bZMecBC/g4WW23B7J217ZnzxfGXZ9RG9icC6Fwk2HhO660Exh+8n2fN
++39tL9v1FSK2WCTAOMeEwMbOdHAtv9UkU5f+vbiX6wbWNh/sfzthEEStC9jlK6V
tUnw/DFZ9dn1M4s9brWKy5vuPPiXCKQN+z5gBKNPssI1A0NM4Q80eySBxFckEKCW
jnkkGZHE+i+yNWLSLeo6Z3X6uw2Wde/t1ev7Hh0GRqY0U2h/F1NQzEgykMCUW1Sv
9pLxIOZEt047XAIUzqGXrjW5WD3Ha7BVXdq7Ha/m4Zc/ySrWZLmjjT2zG4KuQqkS
y0GaGHJc8QQR+HQ2+YPY5kn6e9+LN+vmURvvk0vORBlDnSjw1oIvq6x2VNvNBf9Z
wvJ799CAeBllhNTlx/6OwO2llRfjHryn7Krp3b4cwPiF8kht5wDmfnIyAH3QcfMu
dBmaPg4ikn+iMZKYOeZMTmtQoTawNb5TO0f0Wjy/HznljIWH+GKkQrXU3OXBCkgm
zw8KMrzUXPG5XnpGiRUF/EZxNXFHy0GGxuy2c85kXJCsXjto/gyN7k1BhGbyuFwl
DCD/Rxh9ldpqEMdKzh9AW3APCj4Ek/ab0RCuc1av7BEYTK2upcNuZ54pu4+g/RvB
Aj0XD4Mnj62NOk8Mc3R9TLp+n7kprStqSVq74LWV5cInkbagAQ7z72OhlRJmGyX4
ns2sfiCzlBY/cllzxClykWGTnRSjwTixTtzy0m8/4WwS5jlYbTQxVaQWTFmnIRik
FmiZh2w/HEGoEdz/oy35EYb5akXorRiQKaGJYMtcESMA6PZUQ6zYAWU4GuDzS+rX
6gp4isjWylRPbEDER3R3zgbgYd/rZwno42mJNzswNpxbinHgMTnBzw8dAg+qZbrn
7+ZJ16UT9kgoLkx+nAYT80DVxJNMQmUk//qH8+Gpuc3bjWK/ZHK4VC4yXPjrWz7Z
URfGnnyC6jfSfRlIbSfB9732rp/QxRAzK+37p518vGLzkRo85J3wp44gwOcB05Q3
4Lb7DYPWik5JxaD31/PPMswJKUgC1cSSOQyqzI8w6X9iwHtAitdzHZDshuBO9lqv
6AsVAhow+8tSY2mpG+nvc5+Iqr2xm8UPy/5mB9ZQ8iYi/T/2ncQVDpbdMzz6hDkn
kXpGc76TXotW5dXslLb30hWobaSMrOgFXfnJzaGZygWnaEB0x59J0LyA5fD+5L1V
kteaP3fJTxSDN5xPZbFLBbbGXM8wWAvpe2kPfXkeBS5mP7FP3p+cXNmulKt/Qefv
mK1GZaSDdTR1znTji49vTfDY+nGU1Wot+lopb9kiovPet1R2hIh7dujgMkn3p6Vf
AD2KNbAKJziBHQYzRGdIgqo4JCl7TeqxM+E3wusFo2+AFM0c2z/o32JB2Yt2TrPq
CcNq5/u69m8kQ3Y3UYwgyi/GLmLF021fsoBmGeM+GFoIIfapqvsPaVev3KkSgzag
x6PESCuye4bGbv00edolNXLfXoL46iU+zHcFfVOQTnKjPrykPj3XcMsHyNTxKAO0
IJofLMT5f5uPpGPiE1XYJfGOkiqo8YK3EeuB2qHnEzsSUCz5LzunkbXKv47ADzx8
Wh3vttCUCXk2tE51pcl9eRYTvBeddUXAu3c7EDrC7q1bFPhtKfR6PKoee6VpFYF+
eYWCxrVsFr0KUpopY6/TTZ22ZqcjuCAGkbOsqOaqt/x/Q2NBpgU6hpgWxAc3gdh4
fV+9kYMMow0MAYoHA/cq1LTWGSz1Cw5/5Q1e5j5WmjLtIXD1SPmhLsKZ7ISizVMD
nI5/j8A3xDLpIju1EISUcCRg/D1SArHSJdB3ShgkVmMvO/VRGj0+GlpR6NZXewpt
OLEzxs7UFCZDxvFs+xvZx6o/p84Ft4vitxVjC49A83vyWCwxBbJ6D3/fMvTwRA4b
bBHRcCNP1URycFLEnzfRClaR1sqrroRZjAvFJRU8RHevuN0CEqSA9ZtPGP+JrfDo
stOTonWv/oKIoWLoMMI/DdnvJCRHnMb8mv6P23G4c89o8RkYMedg7knBZ19X5ZqV
ROg+y7FKnkaUtnZ9OCcTV2w3jM1A3hMFjL5QctXDMR7fFbQxBU8DEC4ARkQwHFCA
tNZnGWlpey5OE3ILcUZMBW1r/v5HWUL2nt2CLtCH+TteFIH35DJ7NH4rNqEK/pge
1G8/9DXXTpES/OnyDT6T6SzPUWZogyK/YC41yyvqaH9jLv4F/O5VH1YBPkMDJTqO
9gOBQVHL7fK1TX8x24k2f9OGNKPKNoWXFud7p4t0oOg45mSZYH9f8qaaFhQaEuVg
jDyh03lyzxhx37AihUk1e6fn4SFeCjaR4eK8yaHQI0gfUAK3XhOxv/rW6s00R6Nq
5OJFFsDus8YIYd2yUivFB8KtouY4zh5H/duztk9fnFG5N6H5S3gsxV6nh5m2R3rl
S7m8vnOKKfBlgFD7mFeULf2qcye0upuwWcp4D3++JYVBmjMzS9pxBQELyw0XOLVk
PSPm1B5f85sjcmzVHy7ST64qrQSs6O2tt15Uahl3kpe7lg4yml4PbTq8Qer6L/7D
oFVZeSvKut0c5g+SV05cuhD+OoLySoDro86saVWJBfeW5WZYbNmBMNSO1M2IRPgL
+JNncupVQRG9zjLp4BjtzS3z8Q9wrgYeoRMxRo45nKtcYF6tc5esW73QvT6vfF34
cxGKL+HFKlhLWq11Hho1d4Hj+nCvkEPOj0VHEL00CL+kOQCY1wS+iTjDkeCmajwe
guXFQ52bUzreWVn1c5ihte6L59FQgD1wolVwIX7GDGadDScSr8K7fo1qTQSc1o+/
X4VyV4qNnXSj+QrYtjSOZddUOAOunw+COZf7fjFK8s0v9rJ/XRtR7gdgugmvD3yo
ySn0B8XKTIynEK7u64RlqAiw6kJTtTAQlOmypImnOEQT111wo7C0oWlSUaL7rcTV
6NwhpYj3hMnBXzkrPyzpSuxsCvYHCDCg2uoltSACah8bQtzyc65/SuMFKuPfSuyv
Iiyrc9BTsh4Z+RKODkXVJ0Txkx+FFGluU8ASL+oCWsnz/fGSUZPwOtOw19yZhUJP
KrizsqD3o6c1RFDRJD0jBR5h5kQ/SSPp2mVPRvrvGcOAU/fJaWfrNes1nTtqVlVV
rhSAPcwc/DnteDzLVlZus+wz5Ocxk3NmsT/VFlKENpLWfQRg57DBMiKd/W//fyIx
X5vQOA45LyesPogCv7QSsfdc2PovPRa3I6pSoGTiEURE90035p5oP0khIoDoNff+
6ciLTXNhQVZFF7PgjjzcmE9KXbxOmHwluSUGlB9WkIzYPE0a/qdTC7t5g6JLVpnp
hu6wKs5eqZw17DSmVUsJNYqFEAhS+4sI9kjpNpLiEKiRplJyOjhFuUqNyc93Mn3b
E/gxIVPCAMuDM7hCF4Ga+JExRZOM/VfCE7Rv0UJ/EsGQnRXjWZr2RNcihqPds2um
+WoEYmXOOQsWj/gBh3fDyQNAMF4U7FSK568Ewo/bO832/u1CO7RlTnCvfrbegXiV
ABzMWnKkhn+xCTJf8mgyOrNZwnpY4IVOyv5xugcSfS7T/SeKPNHdX8uQdGj5WhEJ
yZbl+UB1akrMt7G47wa8FnQYPQLHvkH3FJ3NfwtPhewuIlBT0NvhWJa6xblzcIGE
SSOhiLNqSdnHXgJ48BQIrlBniIlkBNTGC/chYkvwoY14YxgSoDY6Gzqir0zp9iZs
imfJ+FaSXeLauhdCzEWSmiPpkRS0GrOJ7+pXgtFMm2Ns/liH1LIRlvZ/ns7ZF/O8
wp7QrEiQqX/Fj6/m79fwDVS5MnfgdMpJOQrncDpfkBapVp+gB0L1XNh5UgzuPIlx
kLgEKL12rNIpxGX/xPhh4MCpWlxUs3EJY2knpXdpVu4lyzTk6Zad1fqLaYPjecTp
K4s5/NldWoVyOvvd/8EJAICfJesSqgFUs4k60gMLyr/5tUXfkb9D6+S3q8aQenLV
UEFJZXtoeHBx86pc6IpGHBFk5IcPiqpaUIONmVRS1GtJRI5Ydrr1+ZwLn+4sg1sJ
cb3tAGvYqIM96HWKwg2xCpSbTTFUsrDNjgy3gVVc98tYOLx20WahfyVvzscsVIWD
JVeB3F92BCBojkY5W4sb893TZ09hgxXeTneQOL+Yu00HZaEQV+UMBrYUOw9D8Nu3
ssKT9wmmEAJlSQiBp/UeQJq/6StK7ce3YMpT8cnxxUxsaMuyV5e1kdUxIUfikcLf
Z+P5AiASNCkNQQNTYSHM3PdgcsfZYIsDhW+8RrgfLkAS3slGt7gJmE4yXCevzr1K
3jB4wR7GUGfAx2W2DfviajyYfQySzAedxDweGg/r7LY7UyCkiQ5QFZrb7VOtmtPE
O8tjOi6SjxrSuguW4GKl6g==
//pragma protect end_data_block
//pragma protect digest_block
22MiDq0jLY7ZD4W4f/fndrYEEKI=
//pragma protect end_digest_block
//pragma protect end_protected
