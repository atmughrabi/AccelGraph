// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gNxlya23Stoi9HtT7k28+R8G+kSnN6s5PYWgpSjoLzyfw9Q5+DdXyP7CGBDDgvbV
5xyHwBF5jUsPm/COIYc6kSAryes4K0mI2BmkuVK1mpE8/YXWPWv7gqXRXRP5evS6
SOBNt/8NpSjbN4wmtspClD5NG7mZzxg/yahCUYNq7dQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 58016)
6rotvh7LR5CnvZ4Ir1R/5T6HOzZFNCXwJQZcV7cDmiB8tH+c/hJ2gTmMgoRzYrfZ
mzGD9x15999TpuSODVcSyFvhL5oLmktkBvkBQhgNtk3V/FHUqngn/Z+115OGUPrk
QrozcWWchW1z9QwAnvbX8oUvTyyc9ndzYA9MDd32J8/xSG1CvYU22nJY1pMr9en0
qAoVaZyc7imA8JuDd7RtVRpPDrz07f8zsHWYZbX6lDH39ykvucWaTudp1pLEv78M
eb8yt4DqIyUvweA9YvYopHIpipYFklRZl7SYxcMBai3YBS+6sywVDUJ/X1oJh1DM
PtBpDevQ8I2b1aVix6byCVSqEwx6p4swTg490UXs5WG+cLqrHfWW1EGGpvYuosXN
9vDjJlUh7BMTiwBF91bfZpmGAU6gvxzGu9nXKMRi7nzHCEdGsB97eO77fYn6Tefn
xi5ro+4nbzN9pWGIqn3qkdfD4umuPR73MbM88CR66quNLREfSh6pSYegvNmSpN1F
fbWICjes5sSX/hVa3A45OB9Meb1nAvzMu3s/HUKT/KhiUh+jWd/apBPzbhVCeiya
+jaxV/Mc6EedJvnbDwxxpFfNr2DD2NvjPKtTHUusI+GsfUhh66VxyH01U6XRK08B
ldHM/s8s6qlh4ASUOGoesRh0KZ2yyH5+Hy96ildlDhnjSa5utlYj7JgzPVqIwqut
flFhw4wBgWCU2KqfUSq/PvZbUDynbbgKgq/ctinUp9BP6m679qQatJKwwrckz1GK
zMSfTWk7UGTCvzyRSVUY8wGvCryOhRog8Vl+TFcvW9xVZEvusgN3k+yOubpfPvkI
dbk1598gDnKW7v53e98jMBspgyKwMbleEY8iO+a9YQ8ldROx4+B5VC+U9y/4+SDg
OCkba6dXRAAUR3TKyLnQRAJDnc1OaVPFHQysOyA+MwWRF09xrTNUaKGLdAAAeNo0
tdn7W+DPw+FK94KsrcSi4EqLX8afqOZdRFKB9iSK2Sfp8oSeE5gWGg3VW2IZzAY+
K1yuL0pO1kFBwEDAqxZp39sFLAYj3GayIXxybGYTogKICOQHzO5WUheKD87guQ2N
fS3fQm6gWBKuKEAd4Dg79VnLKNc5a9nq2aXBMQj0oXTk+ijvbuEFRRvEhTfbbGzf
oMMVfo19LaTrJ8WOqQut9072d+fbjhxKlfLOiBQvwo+MEvAsiYAJQZlvwRDZPuNI
vzgUIdyWkeD9AqCf+NnOXWjustyWm/kpj1nfFUUS/IWxSNjHSfUjM2cWJISLXzi5
05hcNtfgAA2doDZtkc+fAf+la2X6lCP1mJl6T6/c11akrKEQyRKaFFRTS3CeLqqr
GrpRRQFRyJL1tssIzzyWef8Fw4HW1TxhMR1089U3uDZCSlghdvQkJPREqoAfwtFh
DB4jB91C4/BDNlzNWW7G7/VnqyEGTHgS8x/hgys7eTo60A0ucwAlfKrWBqCZ9SGS
YGA4pMFa2e8AEOk0u9nEC+FANAEvkf3F0V5bNyfcX9e+DKgRPBi+gWBu0o2Slc9C
AP3q8V5BgzUHMQHiqD1Xnt7LpjhrCtCGYxNzJhHsbHlYgECeMK/RtkiPHv6AN6fT
UOgiCreRY8csXF2v7/yTVrnouvKZZ+Z4IgDj6yIkGqYQO1fsosTzxSaIYpEoywLt
S6irCwnDKv//01y1Pm7qOmdfkivnB+ZMnoOzzV86Qoc8xYP+4CzWk3iVo6HnqLWM
WzfbN4xlOOgD+YG9K9pSDV7S4zSAShl/ieBdV4KBL303xNmt2qr5suuzXv/jIcmU
ShBGydvJMotPzIKMrIFgKbmbmidBnopEJkopNt0xcTrNyY4WGzSDxw7AIm7TmPfC
+paQB2C2Q7IknymyFw/09H/YZTPojBscA4uV5u6SmCXiE+6+pGvaUz82qHNpMKfI
C6ZMRpkd7nWSRU+dsQ9utA5NubkEMO/YFdahhVofIFvUQpPNh2jx7a6UqQqFzMtH
YkE/qzFaZQ3BNGhirvE635c9NlvnBBl8o+7UUocJ54A6AbQvonkSUk22QCNkT5TD
UpNb2EBjlYL1B+6aKi6tA2U7fmoiMCBrYqzX64T93b3llZ7WcDCq4dw79Rij5Ldo
I9rBrB4Q47eV2fmTnG7t876zaWq6gET+7HsVN5s+B3lwgLqipEf+vlWLsXlAe/1K
Hdzwq4WzgFCEVA72KA4ZIhQs1IX1CRcyQRz9vCdHOe30eaIk+8l7DSe+E9btmeeX
Le9qkHLtkBwIYZZ/zNJRdll8zbvBz/bOlTyqnh9I+ihkb+po5G06f/xgnMxdGdQ/
8Qo2P8dorCJ9iAdwB66FgGB6/mFGdp9VgrkuNTdgb6PvMB+RBgtoeodQMTnHut9A
oag78i4v3Ujc+OOrNVH4p9cfBdp3UqmDdP6wxjJU0Z6eYcHDDHrAVYy2/HMZqo0n
9Zg4V6q2oAnOALY+G7c5SoSxYYIvVJAEy0yZLWPRa9RqfVhqkOuy0nVcbgf2CUXf
u7hfRdeDjnzzr9vVyEEif/vSMB4CZObtDbXx6HKSBB64vu3w483Ha1tgF2c4tTTb
mScLSfcJgi6fufhhdO6naL8tFRr/tj5Gs7yHq8Gq5OjdtyHb9lUiJS5Kik/JF3tr
W7B+HEV/9x4ShN5enbtehGomL99tMbh5XLG0RkEbcEgf53ftrSwj3A8cNgUvZL+m
h0/Sqz6ugeTmU6B4edR7L9ApoPVZ82mhh2HsYwXPY4X6szkiZIYCzerS0e1J8TmN
b0kk9pOhnt+ML9lJ2gGnCJhAie5U3FUx7fXuytcT/ppzE1UB8Eh7O5PZcT8BS/Xq
kNdKHQPqr0vSz/fxW00kYK/sAs+/SKR08A6F0AQjPQ+6DK0oEeA6sgs6Z0MxTf2e
3foasbfvuxcHzAm+uWy4mbHn2zPejfhcwcJooBYU9tzF9NUCfZpa/E1fatrJfCBX
YjbmrkWjsAND7RR+O7nBlFi/+Fcou0TQumEKZi18OVaa8ww6tcWE3LYCN4MUs2Xi
giiKm50o+nkdS40BWM2t62dwX45PlM8SxfZ+Vll4UleRYwHuXIsJGi1AZQTSF1h8
evTUVLnHYysf5gjl0XTQDNVYhWL4QTizChraWcTDqWhr+rm4DGC2G8VwTH0MmL1r
6IrUbzcpEOn/wluB6RraZfOMtkwsX6WLHnX8pqMjFKzEFO/Kk4kXaqKiF0i1ryFC
yUFF8b9O/ypCxrw8xTEtUqM/5BTVvHclDdPNeeCleBuGWnEcuI6CrOqz+s9ksjHU
QKk9gLnw7sIDuF9/EddV2+JILK0mSEl2Aiz6McyMLX6fzoNj3YBXbJToG3lb2GF3
Nyk020vBVStiMfSNfx71T0YY6Seu8mVH79rMpNo4AqxxG7NoRCqoqnPM0WKzDpUL
7feybWh0s1sDeZr+YpX8utNLeMNrlOJMotP8kDjCT4H7bmCZ9AHOhUGt8FerVmEG
m1QjXZMr4LbxGCW7RMDV6b6BQe+krobWsrUbPcDybSvJ3tI0eK+B9XzBUk6Xs6sK
HpuSBaGO8/zwMmmP6cFzOmjiTein0qvnlDF+4DmsE9PZUZs4NFbcxhuMEdwpHZhj
bpbPPrWa0HJcOVegg1erQYKfMdArOgHyAXJxHNwL+yYAujzJd8xDu5hZu/+bw3eh
j4Fa+snN6/aM6yt6jrZ5IvhOjWxkkUI5voGwqXxQYzk8sKivcMV7lMcwjxsHTcZS
DrlR8qsv4hO3MIMcwosweyVYvKdVHgJ+7hJdcPNeFwhguTOc049loMW+vNJzjmx9
atgsf9HdxeE9MH7yYwYtWZYi4Uw+jnulCNSzQ9WjXViN5w2445ERVMeZBsrEhE7p
J1WAn+XvUcBqfbulXSOiSC+3ZvM69mbRdETaUjqI1aYoVar6wuXiJ0EiPugE8kmq
1ZCjSMaWbQ4i3TmT83anyxFG8e+dBq2WNBDxv/T1hEnUj+Gqt5OpMgNKoythMEnk
Wxm9RARIY85HyywUkWTaxoI8oO6534cA/MCC8abcrmVl6U1sBzHfA0W+U2mEK6oE
EuAnhRADQ5IVAFhGc5amO9vqynHYTd+TPukIRtWxgMs7ywQzw07UG+xba5OdHwX+
GWpK66EOC5Asac5Yao9/l97jUXlh2yr06GOqz8NqBNYUvnkBQN61M6/abK2PC60C
KiD+OqyGWR4J1vPlM2VwSsB0ITjL8jBrBaE+C8ScSH8V/kNMzLr77g8jKLLJbCpr
kw4U6/3k81Yb4+XH1rOCBM27OZsxhlFAh/j7kTooqSF/ueImW9iA0V8oVxjqGuK5
mC7M82gzd0YHZXH3DoPm78YVfHLlSoak1oC7RN0jxo3Idsxhb8w+0CX9liKOgwJo
8qwIH+dUhh01gqSFF9alKF//QhagFqda4riIXTUvOHl7V4LG/K3GS7hNSSxawYF6
rWWVUgrBKy+WIp5ARBvwEy/l7jxjvbCTZ3KT+jCAB+jcKpua8rw5uo1OwbCE20kG
X7ihou0uVgXvbphStjMuM6PVOsTKyyNmR/Q0bKdhiQQ5EzMF7pGd48ZYIo1GpayY
nijWa+1cZyBP0XyLEurIqidfcqdEZmd2JlwypQRvOZU+xwEKQFqVOJwzUFW56eC2
ve5svd/685hFgJK1YBlEE9y+mgyLtMwbkiyJcuxpEQ9nH2lt7zB4i2CqQYsWc3mx
Uxc94JXguJn26mntiyZIoFDelItlq62SJIvPf9/+vSOc60jSbwecVljzzCukBeZQ
iYUBSAKeGEOBeHaMez4hItGzW7ssihP7RqEfY6eQZ7aLVZI7WL7hvJx1Vqi8ooq6
IRd7/JB2X0rVzC1MLKtikrdKNKfBRoDOwm4iqw8A47VaRIblKfYYaHLplkRqfn4a
m4yMMOUmmlgUAbRjDxfvjpb/LzY8QOR2UfZQoL7G+Za1QzQ67p28ijwlh5ofzKci
v3HX90dD7Z8W1cUGuYzYXli2vIASj4kS3uQYXlj4ryeO3krN4wVcBQxKPgo7cQ2i
bxK5tduqE/MWlDLXIVZnGb5lsuR+y2qHxgFlGvmS4KX4EiIScmNyM8bFrvcxlv3i
YoFEZpdA+Xk2z0/TRPmR6ueq0Tx54HzQKiH0I3y0EKIf4Wo3Tq80rgLhNsUtAtLU
qugk29JJg5IHNPQvXwUjWcWrP2KjVp8GY4AcaAcmKckTberV38oLHuLwhwsmuc5r
WroSk4+IxGPpUe4cKbeNInl34x+dZgynCfaBUMVbku9eyQe47uLUQR8Tc9e/0Hak
BiGhQtwDfBsQTkWLYAwJvB2A5i07rbDcyE/30zvH6dWIE753eDXf8PHfC7eN2Dy3
oTEC4cVHUPj3TdHnslTHIZq0AlYyzLBwfyD6gadfLR1tYQhyZR5K2rIZFZHpYgx0
pW0gfd2kSA4xLcQwYTLjgwsWCHqKPT78SbfuD9TpzXEdd1fimLr2MvXkhHsQaz+S
c/TIJj1OJ+K0kZtpw202m5VB09IYpOmbPKWfS/MfP7PYh61bF0A8d91s7XnX8hvh
lQtgyq3rnWQ0uIT8giOXq8anM0R+Vk1kKcAxQlVisF9y66CLxt1CFeF4IjnSApkR
WJUcOe5Sbv4ACLvUxyaMUHvrfdW2HUBiNXkNaOue8tnaUjeFj4dzUn9el69VnLTN
ybhdOY/PjIQNL1t5kxcB7zQwgdNy40vv5riWHwnbaZBLPwZw2QiFnoj0NhoOG7XD
yUfUq7CP+CFnjHdX3vpi7JqIsyCDvaZp4njJWmBarhjqOJdIZxJAP+OEvy2pfWMr
VDTVqLlz4RM24SvyID4/2ejt04sYAKcY8b6NuCyYRsCYeGVmJLMFf+vXlI2t1JVB
F4jSEvwoaJHeoT9pnYfWs7jLqkLykulzVEtDqMCThh1omJ725Fcc5N23NLLZq/F/
VkTtilsf9YbJm/da6kGCHLeC/luzx4Mh5O/746YmQ2YtoRu0dKPwu5uVFncEBG/Z
vizib3qGlIJqyfwhiKVbwMblgU76CSbrP3/YUuVSiHbftZqGyTaS7/hQe4KKsn1D
XaJIv8KfYOpsY+s9Js1paQOQ3nN+ev94057NZqPyT4/x9cizlRa83YR60naDqVZ+
hhEJjE0L4oEhv5SNXMsIuA1J8kcVroip7Qr2xQMUfCbxyisky14V0PuoUX3bS/d7
svFMUhGwXB1534g4Z+ONKwS2sOwe25WHPDs5TVxXSGRmbOr6yR5p3dGUCoNJWYgq
SsnFcFML53UsuTorz6dQ0frK98LxIMHYWrusArJNwv1pWSffwKoNA/Ml0O6/VSAM
CFlKa1tg4xx77sIbJiG41VOH1eezZ20Af3My5+lriVlD+Xl+afGn/O7NYPfZFUEL
VuNLfBaSu8iPh6WJofsgNrAUGyQJlIDx1IU264WYkNQNU5qyZb/1LXUTfP0swfZ3
4tPfkQDxrV98gVPDSl73grts+r79m9rLillpZxr+ZfcGZXnNGmy98+vNgim6+O++
Z2yLfeZaLUGpBZot2MyehTlP9LH8idCj3UMDUnap2zWY3nSdSBmC284GBCE/8VK+
mVEPIo0jPpJo+yLe6C6+LvhPAVUesgNUsLjtLVOU1YTJm7992YPimYlU6YxkJqyk
3joytkI2IL7rrI78zKIt7P6uyNJwo96nK5+nC2q5rILfRP/4h75LmeheMnVACMPJ
A590eO4hnCgykjnpwDFlHiRpnB2jQhWDIHM8KVxwaku7v333+GtJ5BdvJtZXaxzm
9Jyh/08T26b2mm8cTsqnL2GmwyNGh3du/OQ5Mm/wu1yX4x2IVTOlovN4n/hfK1mW
a5I117yMPI63jS326C6bT0RDhchcto9JS0cueBod3CQuAiWURgheYfG/oWz+Mnza
qv16T3H+33uOfL4nunyUOZO1vgjPAdd3sOfjE3vNwIVDzYqyXjYAMKnewr6EoV1v
14wFToW/JEaS+DmHmnVf1oeysmg5zRsXZHkj0zQennlVpdDqR7GdHjjl2ZExlwr5
FiKNPEe4SPB5xdf0zoCNXpCvSGO3egE+x0dXs8bBUjLG0f5pTSCqcUU3YfETOq19
QoJWXDdJA8nE8ekKC3G6NlQkTpzbVAsEUbLS4X6SdP3NTQ9lPuPzExcK9i/SG4KO
Xp2kfoNpDJHr9iJY8o/mb1MTkDdp0grG51WdCAkVNnkqokV+ZfDR+R8Wkl7q5hNc
NrYilVL3IpYHB/i5KynrY1RAmWvPcEJfrN44mYqSRHjEMkMxqK0XulE7WFZn0bqZ
/f7ixhfCyWutzd2i1Bcz+SsK3Hi4igrF07VVwvNvLPTEZDNBckwxeMwfGmKl3mIX
ch/fbmZMIfSBxGySnLaJ0E8Yy56c/zoquREgO4tEV93QoQQzt6yRFlEjXOEMyPJD
XSvTGF96BSh8910a2PJ7BbuOanPUIm2gMfUR5F9z6oz+90ghG7YVeWw9NxUjImcw
/sIK8jZ5rUobDHnd7EfyJDQ1NyNLZ/tvzQET3kbf41WxXv+MmcAH0flLR+UlQYby
ZYuMiOXmJ5WYcpQVHvZBvOXEeF0aLgcOEVAqNT0iBlL1Y6fvb+nl/aiYCW1FI2N3
CR5tHLFIR8rPHlLw0faRBR3A98MGygNj9l6D82iKktJv8KoDZYBIcf39+ZyUwaAD
v9CiQn18ENooUcHzAXC70y0ZcrXhQaO4oXG1VxSEw5+Lqp1oNG90chsaWFwB5RmD
PqnoUBu2kIL66ba+4VBp6Z4bKfah604S13momvqi+nvgSMG4SUs6AA+p9XLEhTDY
cIqO+Sz2RtfcL5pYDzKhUdvLWgjHbXg6v+O8AkIfqI05IxOQ2NlQ5KXeyevJqE/6
YpCZnPraVPIp2DEpWVd1PzZf34JKd5HFhIBtmxjpuVppMlBZvQ7XejmzpsPG/wlG
bFmf48XD/qGE5UIRKwrwh6yaXroegcGrHcAbiVLb49QShkDyOCcMmQOSpCumvUX/
TF7cGTYYCYtOiX8ENoji1j5CNeu5dPZK4ufsngWNHvOvhanCxNcFYzro1dW1Ciy+
E9N6N8O5Xktlt0z8D01acBeOAjFC5FCk69eGLNWsBjUUZAPV48nz8e60ukMfxSBu
Odf/NwE2RlDMZlzD5dTzT4sI070anlV/8e65+90X3DANgpYgXWmH11VDXvETw/l0
uwnIrJzm47xg2omnhpKKdoiod6YpEgb/kSnwkQIG8oZ6unK0+mWvYuJGfgJVCnXN
N17vQoYiT2m0vbETx5JM/8O+Rndh0W9e7Gu+RLq8d2l0N7yXX9JZauKVQi8KNUEt
jVeFKVb7kSHa8GnNA5CoHdCNYEZbgTXfFPXbMAHpLZXJHdEvZsBfri2XYaX4GB6R
i/mRblxVY06YlUJqASiwtdMvIeaJ8T97LLG7CuJalNmckxlpErzk0L1a3AM1VkaB
40g6ucaK5PROleCjDlgtTaONQYF/0yWAr44M5EwMJJS98/Uli0o+zZI6HqhheJ3G
3zqRtwO4RmG1K27pXA8Rt47N5caFxyp7Ls2Zr6EqZJEbUoDVig/eaqOhqxa73FiV
Oy8lIARqNqC1k2pjRROBevxTJT2DDtf9VZc545yOGvqnLfEJhk6Z8a7RZi2zb9Uf
tds+9dTLFoHxJNF60RPUDRWi5uejvYlb0ljtGRiiLQ3KPNzL96fEGnrnYWS+S/ps
LVrZSXItb+vdDkfrWa5FHJVp5dwJJ4Tksc+capvfIgYA9lPMbeP4chCsk2ULuvKN
nia1fefsUwfPw7mJG2Ua5lGmLsFa2DGxN5MnfWpNiUKvIq2CWgSMYQ2fTfsJQkW1
SeWiHA7FvMACnHJg32aLtm3Ks26opIY3hI2/MlHbnZEoCnsm/dQsNVBLpD9aaMXk
lCJFR7VWv7qwL1T7zJSV5nejByzGuPDayhUyuXbuwZsZ8LT7pKg3M2giJoTzyNMh
ZSd6P0C6Yjm0HJZ7D7EJTZ4czQWw1lLhkB3KwlViOzvJXICWdydWJ2qpKIxByZRX
QBK7yke3UnVXCHv92yE3JBW1Zd8uuxmKlvoULu26P+sO8P4lfDzSEm8hdwXC0/j0
e7UZbLtl+z3We/yEPe6V2FRDYtU2BhfAxCD8RAwmLrYVtRMgFWAaiXzjeC7Ozjul
pcryCHEP/eLuymMlXxKLCSQXykSlxYcH6pVQ5+JRevcs9aKFocA3eCzIGI2NZJ+3
+LUM4ypV/amcZS8M4JHz1WIG46APsGDf8OYYvnqU+TMNneIRq7JNGQdhuIRhZG6D
RbIOY5Kb0AIAFwkkvVHGahjkO+9VWWegmtaVkwqw4tcC8fkZNq8bN1kZYivq6wUg
zczyVj0e6Q48VoQiigaxkwZyWSybYz8ZBvphD0mVO0cRUuMpzDpRJyFVXGz8T94o
578/BrkdjYekornTqA1YQBdEHylut0G+485mO4erC7eDjjTXoPTtCdGhUsDupfRI
2/p6Hn8Bx2lbJSV4O/LlHcwQk0CzirRT+GvrptPxE3qPadsgZh/LkFVYn+QSYyBI
MR7lBAPUCRLVeaCdJbhy7uJ5VFH1BoXU/KeECwZMqlYhRyAsim+FacUyPI5TPP7m
taPFIbP4taA/sRYa2hJzQ3W+DvrSMlYVIXfKF9KwYevHp2/T27UlK1isZGfL+2xW
P2Zyvh3zg15aF4dW9C5uyJ7LU5WOllB0239ciAduMizi65xmagboADZTmWruIkYp
HtbL6pYRDIG5SbuP6zIWQhwn0GCu0Qa9VkgI+CI8cAGj13XyWWEKhlq/Let7jMrQ
ZKYWYkfmRtdd4bz5u5QHEEHjK5tG5vlZUK8bggpGHwYNpg5T0wRTzC1KDVuwLv5G
y5xkaZrsN6U8T02tB0JpqU3X3GQbXn3qAIFmYSDZBc7FQIYgiqr5tGV23YtUQa3X
DkAy70iPIhg6HRRiv3VzGLu0RDwl4bbIgzUNYXu0emwXX11/dCu09VKMRuXvMqDi
fLLerMdPvpki67Y10jwoHLTyuXGad5D/RLz+MEST3W5ZU3zgftvhvlRJBcWqd/oa
sWrS48w3F6KhNgufVuAw8FfuU7lSBNx3KDCjOnzp/jJoYQwCsgmmz1/4mRpLQJZs
UDBjtfzX0S5I4uTl3iUEKBTDmZ+Rt8TM2Bticmafe1IZfnTlJbAohvMcct6c/z09
+ZR2qFAjs4YS112S/07+yesrGfpBFsQgYodAuYGdWS5HFv1RY69YfV0/suM6ipUt
Cvn2A0eOiz9A2teJHWWcf77EPuBbT82s1Id1ssU7z84wEPeblSQUylsHljnRMD6f
NxWSDs6Xo5It0XsAyf/BSSMiE9vKfioY1EtXuqtCz0ejs0d1tzmhgyQNN/fu6yhY
bBFpRy87FUYiCIEJ1JbaZ9cHQou0sLy2uQMv+7vixvzpxcBESan8e/vpoLFMZLzB
b6Dbq5DpSfj9NoU409jplnavnjJB39djifeSH/WSasoe9XyFWVMTy6HM3YQ+b4fA
8ApNdcpAFg2ZRLmgY//3ZJYCo4whjIBU+n/BLDgTM2Gh3W/mgM1txdRDqa+I7/qR
/eOOqXvpyW0IKPTvywlKFGNM0FWMD7bY2UWtiZZoUsaKX/WJOzyGA5PEux63M6/i
JrsL54cjZCJi0mBm8CO3sn16yZWdl8UFEKoEbXvu+sHI22UadexNGyGhyzFJdFJX
GhRjZqqFlgvQGJvmt0OlJEpOOdkg1v+NCG8Aaci+UfpjY8FXB+BkIu3K6x1hSHb9
FPqeXQTxHrya0QvfZiOln9qOitThuQmBkYVMk5FXwAXPoZcuPur5EoIwHjjHu3Gi
LUOt5c9dFzQ3YZJc1t0hWMd0Ns2y16Q6tTeNkNmcUih1bYkOTJ005Mhc5pLFzKyF
nfIvN41ToY5IlBVjPnYspToTgEWIE6RBZdNnPXLUSxZmE0gQbNbhn6vwsnvU90c/
UO1Hk9bETBVBIH5tGBMCCf/wmYHOuBTWuNDtpPGBBBlnIZZrCR1LJeEXFEGLddrP
X8KHTXPZOz67V2D5I4jiBy+3OdekFBpCCBQxn8C/32UM4ObAMBpKQSrhlpg6fZ5l
CpR5Ay/fEuAKsjOZEyP0/lupxtvLKZabFMqcjMeh9Dn+o/hCzwDFiRNk1f1YoG91
OsIZLDuv0CNpsnQTapIDk9cGSPVR0E6ugR2COnF68BBw4XpnmgkaJkYSO5vOQTv3
YKIJjbUorUO8EucTojQ9DuvBINmzEkJpX9tYoh9aNIDatnsXLWz93tfoJMIX9EIi
DiMocHYzoF9efZ4bgcu4AUHemxfAxlCviuz/bhaEEVFXRFIvO9NTtp7kKG6Yf8nJ
C4dUoS2MnD6oGkvv+PKveHgdyAnXLrn/NOXNVHyNBhi50u9BCBLYyvEsbabWfLwJ
uRNmqM6FjBWZFlTvm479Y9T9tm+RqTDXjeTvpAG/chsEItofgtY9xYTKjTaTJwfb
vYNE7v8m0droc3/4xr0ryVI51FxEiFvVg4+013IPvMPhPEWeVcdOtHaUXzdml0vH
4c5Er57E/nZV1oGfX2QcljZdEcy96fEgiAiOdiq275BqWbfj1d3D1pJjkWVc0ALa
ARzS1pHp0Cw26bR3KOGLw8GcOHGh2sDS7sXOgTbwTebRqlpCms8M+HCI0nVLJ3kz
1D62QMZfszIrbl06nMdkUWHvL3Ua1tK8L1QMES4+r8Vh++xNHfX9/nnjrA0lOKqC
veeQX1FdtZs0VnbiBg4ZJ4CuYuZSoL89/TICfAJ2MLwDuXnz/xZBXcvlInf5ABSd
PQidrZtNzMoLbtp/VXVqI0vduYaSPUoy+ETFJe+yGI5Zl4AnmP6ovzKDyhuRd3F7
asOuaevFC15RjbuMxt+sIfR/iYwuPld54KeBR+OD8H2tAnNnL4RitLJ4ju1iGRHB
tBFdsrPwYafiV09+GK2rbP9Paf3DI3TB1VHlp3HNnx4RhTNFT8AfnPS+GTNuqwdk
gYkUQfpXuDmipFaAiwzu6xyXqbXdMfsZmhzhUtas+5cB1bK+XAjCG1PfeX7MbTNL
eHTku4RMok2/h+kNY86pVAQ+p49bcXXAkoU8ZAU8iB1qA+PuLTx/cqmq9LO3+GjA
Vftx3umZPokGnqPQ8fBiy70Rsvim/vLIk/haZjUd5Co5tZGO92bWLi4SqurfhBEt
92pahr9NqeCthnAwfk8cqnDQ35vd/6RidUxgSm+LCZstGkhxi7g8hvS0bxtPpo/O
rWk2H+ADClIq0nnZ/FNISF4Rg5+ZZ/BSjOV6rmTunB2ESiyzeuBfBqBiefeuxjqg
A42QglGZLMjhsNlNdEvGhLGEfa54mQC/1I1JFhETN0ENe+c365GSwGlpdIY07qK4
ZvTBg1kxoVMpsKYKTYTBJ33JHmlJuU/XJ7v7oiL7En9tkjpCFlGEk9mjvAby7QrD
OP9uhh3udyVSMnhNkcqtDR3UempbdGKDGwyu8CN3W/I9rhkfVO+HQ4bTdTqGsj1J
PqxEgY74+OpOq02N8KlEILnik+ni3pnAtZP9s+pvge94jNNwoS1qQZ0zxdlO6RYd
iSYTiF+X+0Zuyz5mogkcf++VS/KKai3Z0ijCHrDemNYsA11NY0nUsLvAAjV6hZl0
7ai5pw12ilTfsekBoK8uby6FKcb5OQj0xjF5/J+ofMPCbjTIMjE8YMFngqLCfD/p
hdeLPETMbDZ5ug6XqcOEQqwf0ClXmVxl4mxwxKm1rCxMKLPjOjwDuFwTwLnKRx6I
BgfbRcH5kskH3PLCFr2m/HkWVhatUDAryCpyo5bdB+cPTjDgrdIOyBBhWpzzegcU
ZraTIpo0/mQ6DmAwI9XjWzPo7loU4hwwS14FGhoc1Q3Gh5gNoJ49cOWLhDLJEcWP
Md31s8wCMfrIHL445dwoUc3DHc5sADKjWcHZPDV9ws6z8rYOxEWtzGNhQWsZWpdg
CT0Yqw6RdkJfCxSFr8bDH23li27doriovAcULHTLMWKsHtbO0DsXb+Wmz+Wq5cFG
0ZjowIzznwsWiS9aYijRLdTCUCERuAiHd4xIcWXkszb9NX10x8e9ZhF/7g/Gc5T/
nhiRfJDhKfsuJc3XM8eSRBr/MgUTRKDAId2seisosiRq5uTtlqayE78cz5X9PxLz
9dMjV1W4oD1roqFnnqE0VxPy/tORh5iLApzfKrj3sByKnxLjh8lFHrcSV/ijOC81
t36fY584vBs+E0IutfVwm0ijJINKSJBQUnaianFVkgwG7fQkTauhq6Bd1XjncSC5
m1XQNUYPHTZ2PpCakOmSsMLHIpBiGIddCsQmOs5U/ABkosxWcV2fcghmlXPolZQE
b+9s8UyMVpuqy476S1D6FQSQLjoBAM/BH5uSVz2VsW/0qV43CW+EashscdvRIeja
g9DSar7dmcWLDbBJgzep+xQN16eOgHQBG995woVGRd5SiXrxecXxeWHAPUGK9bZT
/FZ6kdKSjNHYwqnIDDBBTi1V33hgZkKGxEm8L22csbKY8iAdkr2lmcfS0T9k8d/B
gAPVzloAtqGjJAOTUNifEwJfPq+hU83WKnhsn8dVFEvrVDKvm+UsMLYjwt8W7Wf7
y3vGLO9+d1qohQfgjC29/QU9L4sFsOEG8J7jvPBV66zsI4gekKdhR/kfT8VhBjj3
TZ14VGGQ47L1oJTh+Roj/dqflrcWQwWRJjQy1w40K96XFb6iMdIAdpCQV/pwWxzt
gyZJQE797Z/Q8UEcphVJP52j6LLJPU7Fu8jiewEjjm5CUChTwGC7LDOF7MZdIdhd
bc4D0VAMK4vOwp9IxoNhp6+2sVHZbFeuNUZfoUrqxhhiH6ivndEKO1gp65CscSFo
r6hDcImkC66cVKAYbj2/9OYOswSVdOm4tYur2OtWD7swJ4i+EToqvWnCtV24uGB4
2T4h+aerqL28djPTbGolEcvkbyV4QtysFOlUDVrTpj48UjO/gufILz80J/iDkFiq
Pm91j5RKzdQDJcvVY7LQ/eW8EVGAhKvKdZ6sb0cV5KtsJoLn5f1zkwpp4+tRTLDr
NlqTDN8s+Iwu9nWGIRDVLzt0d2ZG06tvf/VNtDOuns3Z1bGpZIiv+eayaYwvSWov
ypmFfNac4+aYt7vIMEpiMBnUrxMN5Ew/atV7/tNXBPCa6ZVLuj+LCHeCismJL9+c
cia9i5cVGu1lgiypIAaW9xCBNGRSvjTbRJ4/4qDoYlRRV19tW2Et9tECBty9sUGU
yULZD5BTyfGHxhoUecVflU1foDYYGxlBUuZX+KI+uf8ctP1AvcaWx9jIY9nXvR3F
/S+dYLhv+r8HNXr5gvIp384pC6F/HERsfVfE/KHD4EPQ8gWzuqt2yKx/rYNRaRHm
Qct3LXXwegg04abT9seXb6+fm/GkYdXiNCwYjlsyzrayv82TfEqELezS0ULFbEUJ
ddgH0iekU+Wg5n9P6ODm/g61f2SbjhQDu4/epThvdCsdMWcWTi01bBvdSsePl36e
yhsm7pCnNei3vhzJYI9X1nCoXWbYBzyPY7EG5mdt/1vDdvCCzhEjpRay2SvYxPCk
/x4B43NfgSGKKI/l7C3HGXmEjf9EX5AFwb2EG4rlSrsrsmv1Tcq9SbWzxkKip63P
7e2sw+gSmn+vCj9YsW9STqPU6GOJsQx0t07ennG3ezanGxHtW7Xdo+TBdvJdeEZt
Qls5J5RE5LeuDXZyyW5h5QZg4JmntVPbiFnBO8acWhQYP2ubceDauw3BbMqKLOLm
pYC0PkWiLrKQoy75neyt1n8Qt1gbx+CmCfIkdwBdilH5jbZsrr+LFvegbF4jmXl/
rt7eMDDSFgp3TnZBBwgDlY7KTaZMS8Bvn3WttDh5to7Y+PUutLGAfhCScTq+5C74
mnLk9aRWlwTPZHtT9LR9djkOjrI8BoV2v/nZSAQameOQvP2cE/iDedzyKEZNWwwQ
gbs0obTw/v8ruoluN8tuGqEIOn2DsB//KLchqVq5us8dOieNX0/jSOIe68t4Vd6V
1E2ml47KBXmmLYebxMdtRX08y9bkuaeYub3VjOec+52BmtTeX84GgwPZk+CwNsDR
7kvdS+W5Nyt1LTwS7DakU4IH/S46cbdcLeLp3PUOj2PEksuzljxMRzK7amum+of7
UW8s3wdylo6Eg5Jz5IRtsq2OL7mfWZEDZOunR+Q3cQKDq6p8MlThCgOXb1RPkOru
H0rcg3JYqKSGWjN1MQ2L3oh5qbIEfWDOd9XDNDmL85+r0k6tYvaBXYw2aFFU1AS5
YoO0FoJYfNQJjakGboExbAXOc/UtARQJPrgdpnngufbp1Ulpgb9tXLTBdwRvQzvB
GUgOL2FUWrEtN8eHENENqhu38LdnDJ4S7JitwxDs/oosXqvFBDCO5DsuiiJl/L0D
FCIQ/q5JGQrpkcwb/exzExP9M//2peoKyObwmX/iFNSWPKyYoMsp2LCBx9hECPlb
6PsXvTxSD9iMJiIcJ9957ZkbUSer83udZzXwMAIU7lyZE87zziK81fjB3kCZqrOd
ftcFIM2kT+zvdjrjEAWmfZmPV6cQVSRjrjTjHLYLv3uDcXWU6O4xvxpd8AM7QHsQ
McNiDQ6D+fPOyjqXBlhyU9tQ9pZGgU8VN5OIRKZys3d9lTyKkF0gU0AlLtJurcnr
kULahkqvblvR3lNhXnJtgcghnUA5a5r3Hpj6yAWGGacWG1AmWWT4ekxm//Q+kaYv
K4rgviZLK6VicIoeCaDXTWqS3HAWMcBC8tLL42guGu4Mt2MS1NaY0UkzpapJAYJw
atcR8+J6w0wUvKGFHwJw4IwJtA8A5FHDJO4WkNxeEAdGetlytvvXtXKpWxc6XWNY
JRNcg2dRpSl3B+5hCbV8HYSACuKD9K9vgvGHjW3IQHIMbaE3+yehYgT0hhG2DxUq
vGShZ8LxlcK9NGq1/Y7wIl9AtAfmyTCkdEmEdU1yuZ25oqjM3PqdVBBeLgb7hoYq
//Xr7GVsFUXtPf1+JfHIxJCxwVd1WJtbc/1jcxtKJ3MAqrozdOv/iaPEN42kCuFu
0QmWtT5hs2eMwwBqSraB+tNhFB8dm3Zb8TVJCjcyosyurbd1LNtXX4yNjv9RSee/
CuXsbyvuyYzMBup5RAJtU/4EujqiRH6EDqVQF395prBSjKWFxOS3SYEM9uYmbFZ5
gj+fuSwvh9ZZtiPfuaoegEM3BW6qLG1+OlHwi1hCQhGnotZCSH00ziy1USxMiUan
ANz2aLEN5uQycQH/TZhgOXgoBvi1iSyDqX3S36g5bnasG7ir8kwMZCgf+Vm+3W0J
gCGZbJq86zp+brR8VDwUFc65bclLwqUlsRfMkNdB4tE8XRrrkdW3i+0uiAxTBbk0
6dJ3SxCFuBt7Qo8HHGu0Z8KUAnb5GJlOYGFzsAg61hqx9R2d88G/tNV2oBznz9EX
REKEm1v+CMTUOvDlDXAevr/0LVZuGM8DHS/dYeeXbyX8Srrq/CRdhE/BuYoYyGQy
rabGYiNqaFQcbpwd53mpw/RKkdjj/NFtASYsQmn0tP+3EubX936ssVDVhzfOwPf9
sp0xMbDcI+Vzoib8yB4Na1nplJP2wvWlpUZaonNTDOYIk7QGN8PNHAmXZBSUApKW
gOHbtqS58hhhh0mSktb75H5szPoPcS3AzCliv7CnjQNJ66QgqxQ6uNLaTTf34Aor
+CuytlYHn0H+A06V5gC7ygKGG9V69u6fxaa7+ww7ibo9uc3mRQ7GFyuqKZAS/eKZ
8UilEU9BqO0R4AZeu0OxwuDbDhdGo+KsGA395ncMy32tqAOfIa0vln3cTF8/uSci
nII/gSqRBW9bMUjH+YcqcqoCURWzMEtNUCZVlOtS3TqjVvrXX8opzhk1yhfQ7WuH
RB6TWunI49iGc3KRB6vfcQGUtgc58V+1UMkAxmxDwwtjQ9KZU7UArGBr680OOvKF
+qm3NhMhLC0r260wfM1b47Fj4obc1FkJ6FRMoMVU33Hf8mpUus5BhoEUYUEbPfyp
6VqeskmMV5UAj23hfaCG2QoP4t2HGpX4cQ57Wuz85bTnDh4ihyQTVLhI723QIY1P
XQWz0VoSuPqFM8oXHz8DRDLpnU1ozz+zklirnDY4wUGiRDxiC9ORGyqeviFI7kch
oVQZGOe72N9/IR+wbNTWRyNGALKy+AGsZRDUw18NwJQvdTq/Gupq9+rliaGGMrqn
j/b7oscJtyFDMulrb9vMf3H7LYt7yE+r5WTmZlRa2eq5DWOEp4R8Zdf+buMjdqce
AO7gUoCenFo35nYi34BExIWXTNMwDPxRHwFigf/BDDMXYRlOHJq4fWmjJUgPCrVA
Oe6IM18YoTNoU6dkBiPH9JiC/k+a5TwlHNa+3pZ/dIQHQCirAeGX5c0OyIu83Xh5
QJDy9C3FH/FPBnUe/ahbpINJqZTjxIfesxK87DfYDxqSm10UwYI7u93hUFebbztA
2gLHTDg3hH9szGPkn2C6iC6n+Zg9buBPXOyTmUWtK/dvA8Wx+HSH4+W+BoWA2rWs
26DzUCy48/lKsXAU9mU377R3DEBpM+MivDsrbwJ40dermP60TSEnWHptdT3npmQZ
HMM722l+aGFPq9VLi2vaBE8Bt2K6xGuN3UAdrfdwNDurrd54ikB+At1iaLyV4gwW
c46sgOU5KHy6EvKZfV0rM2pzQlAmLQccewNwuz21ClpyFIHaf9BDfdP1DXly1/FY
EAd4z9fnDzazHCagoRfAzlHpnEu6V2gyAdCbTWYvrhbT3QL7aHYCKLrsxLznxljr
yU9UCEElgal05l5chkuHKLbGwPtaR+52O0anREq8PjuJ1SP/ZyQ7lfRD484gN0+t
mrm3DXmGPjewYTy41nmYgTKM5PkGGmt9ouMJm30Q0HLGuQIRvz03HXcL2j/Y9MX6
vZGZgzexp5LsdhDIMqzzRYGaEDMsV0qHnOnDRNzZmHS6uyiB+/Xcwd1dBR4Iog/0
QOEi6RBSsLDKYBFdXkGJqzeLJIsZVNRBiHe61PdRvQxL6m6uDud2wKULBrZbRSIV
xJV9UImbpcndNghzee5bYfd8QOQ7zsoze2HNAsXvWTkRQ4Ve+p6huDHLlCjjbUD5
F9ZhqpoyE+bcXMJDpL1OBbU17RMLrvBc3tYyjPTQXmz2AUGDYfWvgCwnCb25ExYk
hvAdC18bmPvSa7/0PtQ4JY6ty1/oIeywxiGrJrOuzv53QOXw9lIUYvGIynSDdDtu
e2zYeS+Upa7LWgOfGbRkXUeky14cyJLEypnHtxQchpYndORe96qj4uAl5Om6dwtt
hGwyhA5EPaoRJfXPIY4yD04OUb6QGZR6KE+djQRKZbooejERZjKmGoxxdOlBPQCZ
geYXrKiYjKgq+NPgFHRsOeLrxUO4nKQ2WOObs5RKwHpgM2PWGXmCRPX2FLbgNMLH
6qJQEhFD6hMdUD09R5YZkE7VFwUc9oqLmKtLgDDLtqc9b6oyC92cF3g/D1xKbQbc
UDZT1EasyusHr1PDVugcusJ7BkVsyJhW/VgFhz1u+xQLpDhIFQKEOggOnL7uWNi0
EpQ9iADl2Ohivhe8OowNcy7RdkuVgpJbL3YPRzq6KvkNmGcaGbva5yp1Dz4g6F4q
3DtFzk5oPVgSItoukAMp/q+YZRQw/z2LmPQO6DBKGfz0OBhf2Zch2pq47FYQpQ0n
AO9cV75AJL7Myh/MSMATcc81dW5ATFLOVjmUaPLPQzFijI5rdTOiMZdnG41Z6gh2
UFbrV/rJu526oMg8sDUhVFya+2Gxss5FdOpYyg7hrlq2y9HOdaEH0Cs1b5kUyxxC
gqO0gdirLCoOWYH5oD8nGIFHNZnRe+Aa4QP0gKHctBrVrGDYOMjC64kPWTOM9Fnk
wUO1uvtM1xqaLubO+NAJ/KuyyDP7ENQyrqTY/jbvM5pnm186el79+CW/NthkMGnd
dFDsiiuSLRDRN2MJpikYU9Lyd7gwdFSbrxgXHHeFKDUBwh6db6iFOZKXOnl78XY8
/qaSGa1LYpFbRSJ96mqRI7kFIRtf2OpN4k+zNtZwGTfWhZblEk7GXHeLxv+WZ3Da
C+yE7OcZhhgnfxt9xOkff4nlIuE6emeOQU1WHmoaI2Rn3W8p2q67VuVXS4yoYoXo
gc9ecfSkYMZfRG9rPsvvCU/5voIm6NLejT0cXQHpma8UaaGnYInvtXV5Hu2hOaCr
X9SWsvVdJMxFNaSftHo91Ha3aDob+nTPOY5fELPoSqxtD11Pc9vMY292XLJ+XCp9
NJUzW1KpxwF3QDQ9jYqfWGfhqBlVHgnD7uwea7IqWBDJ9XsjIFbciIUNm2wPZs9W
uVFprCfBfodJx/bUUJfAGkA/4R8Q9rDWvPc7xmBP4L3b5l7hZ5eboHTtKZBhJC60
WdT8MUBwu7hsYO0qYzEJEij6ypKrfmvWcyH3PWVmCW3SVFO1t/67nnq0FUeNxjdp
nCNlrI7y9N3LVy43+CuKRYG/J1lZtLPQsCMdJ7KiTdDZoQzQH1p+MNvaM6BVHHIx
rDid1nUyazdnJN4XUtot9G0f//wq2fXiwV7hIN+foZ4SuUR9mM4IfinGNcGHiIzf
V7tPEpzkHHy7A1tsYBd5c8kvFjCu6MH1WRxABW9ZUPB7e21+hrJDuCoVRmZfLeBn
3Kh2iMyPzUWROxA8/GVgxlkL1Hr19oLCvNnSUBruwiwL1vMVRo/IcEMh5L1fq5up
BA9ECLdQzc3Tn41ZcDqymkb6N3ZO7zpQ2S/LwLwvjpKkY3NZ5cFoTk6xcxskvnCD
kcW9rtxLWS2uzT4LcRT32+A2Cby1OOoscY/Ov5SDsZm9RwYJvZwZ7vMkXDTZUz2f
0MtqBVmxRc0p5eyk1XfQcSYOSqhO/wSf4XzX2++EZ258kFRFAvOKXT0uIUjmEk5J
T2zRcajpGSW+9Aq7cuCuANeBxvKydFsULeeWt1u8Qn73K10CIGop8xAk61FB74nL
r7QD+9H7kd6u/kpwHxRnHqQ9f4z2k+tRPYA4YrFG+WPp6OqZGMSkf/kUamFjg9tF
4R2qXebCODzeFo8jBXmJHj81kHd3JdxH1pJxGT1EQEmOWnIy4voopVy9uceeON80
xBwD40URi3XoNx1hgPAkfUjIzOE2yyqIxYTMcLwwquwLbxu9GeKYeQRldv+QunAK
orzvXOCsaEHiFcaGbUFdRh41D+Qz3Hyw8s5YqXUZ4nWjQoXPD2DcWQOHGE//8xs7
/rDF4SfNRiVyYLEPO4XfW06ITdd7C18bnWcKLGvadw32LrU7tTCdbfgmlw+tnO9T
AtAQWLPwo8KqLc0nOIF83MVNkH2kxf5woG+WLfwtjIGQ31j2I3R51FVFGLJL5tyw
0qqavvIbIZKZ5TW31IlnVh8wdLv9dZx3/8+GxY3j2WUb5AypLEAJl/zdlTxagmeY
l65yNAq8m4PCzp7vhMX/aCe0PIU5RnYs0UTPbefwfzeJKi6mk1iAQNFaB5OHv4L0
KNJyD2KL9oMxZMGlE8oSBRBGpviSQZE3g6MKtBnAA4tFyNs9NXN0JHUOy7vWlub+
kPrdMcPooj6t9GT+8Yu0OiiwsiLE06yy9w3RgkVmzSBsg2jN24TVQoJ68dt+YZzC
tAaj083ofrn01TddWTIMmEYEMFwZxG2dFIiRJ1UumvG7fmsJBmSi5jyu0WTzq3ej
l7fQqa3y63Wlj59YZ7X2k1077933/sydQ0M5lhqa7/u1aF8JbFhgMAJyFUm2TjcK
2nI3tE4LFi2WN/K1RhZO4UJA95SV5ErzfB12Q7+lKU6czidaYWov4jSkYemFR7YF
ziu78SHVQvj+eC9nC5gBKCGSYlUwJdq63r2KlTsrdzUwQbmJcInfJGzWbtgLxyL1
iBLoZ0qPzW3w4ItzS/lFwwXWXcJeIVv94aerl6mkQUm+ewOGDR1cTkjM61BA9D/G
thOi4enltuX2r0ATSLioStxIZ07IGJFxBGX6szynG2cdLWmdhs2vncYxY9iZRlbR
jyE2nt58EfwlVOZspAL60EsiYA9tUAk1Tp4dUpp0F5ogBFLGu3vaFitxvBwDVzV5
5MJeYtoSTE7hrZVi1xaJutCruTZk3rMP1VZQniotR7HE2RMrr0jah3aXMIfV5D4F
bOuFipdRvtjyUqJN2BuVwJoTE60rDRw1NdeSrsbMnUW+2FAhHPdUlNAGZOMKlcO1
qQR+yMUE7vTgjYGRDU4hEVsbiqWe6cnTdvJubBHOsaQt+ZJSxVDb1g1e8REftKbl
osnX4ZzfoQIyKYdNEMlfJSHKGzX8hhrVmZsoznk6yCT0tO6597kJQjv+dZTrqM8B
3UXaj/2MdW5U8Y9h6dsvO1Vh0Q9C0K/TK3gijNqyj5ixNOdeiXygCvohMw0lYQ5+
6aauUHEew+lkyRKdWcubDbYz4EKYY2TQaD6Snzp3sPiJue5El+Na4X4SCiNLQ9Be
9BPYCwjlgoTZvefHdal/sOl0NqbXUS69IxkycrWAn/vxsx398R7Kpxq/EuuSIHRF
/Yktrww8mFqKAZxEkWveFq4iVgJdSQbJUSuOu91reUEmY2rZwFIX2XTefg3B5tJ1
WeAh5fGXzOPUm8/yRtdFeb4SQYc+eCS3hi/aQYXn/aLeqhLR7TvHjqRVMzMAUkqK
114nQdXGe2m3Zyc68edvVuXEjT5tuHlfSAxG5mqc+7S5UBLc8GVIWLzH7pgddHZK
JAqoCkOMqFuqPM2b/Uf7ka/VS6z0bf9Rn8gt6Gx/jUt6TCfAKzWFV+vOJNgO55RP
aAujfdDIU6bCTr/oN5/xDKEiTDkQXP/GkKzczF4AnUUkyWh/Q+KkawLHvKr+E9yf
IN5MZGKxBo6dgPAbkhzc2PuMPa+u3SFYbZlq6T2ifsXmzhNHvoEx9YlQ21AEPfML
xQHuMG+PJsnJyIhA/KagRmBwvRYf0LKAS0/L5Q3Z+egKTr6ODcGE0JCYVGYO4/yH
ngPma+K6R4hkVK//Lr7x+hyzJl3UlIwxRdJCw84J0UHH6iIGzjOgcBjwECiwffjK
6Oxo59QIJiGWJf0D7QAT5adeO/dT5Fyh9Q49fgKWL3vBzyVQ+2+uF5eIdxSvXXkv
VdH6Ljikk82kC9XRQsZmTJSa0Siz6GRR/DljfTJEVsMMQRFMJpu9Z3I9Tud8yojl
PVNoKLqiGs4oV3cHIRyXVLEzLYqF8sDbpBS242WbQOFsnaV9WiztqPt/GKRrZr18
CKUdJywUUF/mzN4CpYwzbkiU6sn7b9zmI/DvxEaKDRx3X8kEYgcByN4sqajecri3
sLIzNofgZiXsBqskF1kcXsrtP0L/Uki4MdqDfLKhSDT8EKNRi8iqLla4EuR8D5R9
DJ+LqXPvOqq5u8/5jEwHfkt/Eo6aAgbzg7GV/Fr76p/EpSeAHmHdEqQ5DER2MrqE
wq/3Mq0v/j6liUX07jT6/Eg6MlCMoY3HU0j9wKehvgmDy3JvW07QC4fwTFchuOIP
kXzn+708RIPHsjzXvu/kLWi2RhAcoYGWhAC46WH4keu9PSQcqqFNp95uS07sdsQF
G3X5eDoLKpWO7RinhfOPvY6HF7kiUt+xOM6VmHzxXMAtUcShpun8EOXZBvH9E5D8
Bz8OcFmuQR6iejV9Qv3RoULIuIqY5nHKVovw4QDpX3aQMHq4T6GPxih79/u3y9pQ
O6ZYfBAIYACMrncx5gz7PvAXwvco+/u+9/OGI/GLIKt8Wc5j3e3aeZK4oOJw9xqZ
uwA6jry3M66ilDsLMYpOoXwhC8OIBUBu7Dss3qQ4HIXw1qkhYp09MfUdwonGNs3b
hFU8VyaDMdL+JOWdP47BY6hUizlwNiLfPyXMpUzIpyXb0Il301IVaO++cr0pWKqX
QQAmoOeLFHCWFSAXuu/kQGQleD0pGzQPhEff7p3sxT5q8eHll5908lVO965RlgNE
PMJE2rPdIWsN5Qrb8qJFUag3wlSPg40v0eKKKkl/xinyzydAVPL1HfuvUXwCf06e
DGjixQUgJjXlRCiGKOejt6e2F7AtrQSLHilzloN2aHCozbzBfkfZzxabQW3nS+f8
RmIpAbu6HDKwQO/0QgI6zOc9YuPFdPE4zhvB3YBx+z9+lCQcq4ByROQVN+ZFTETU
JqmLR0sCgbFEGy+kAHpBfwH7Glc7scd+YL71jbJb2G2gsyMCEPYlBoNI3x8UVnps
7dDWkfu9IFQbqzBD2/vUTPO7UKargBgO6rRdhhSHBD4Aqbf1hWkeED4+nW876ZDO
2j2+YExNWHxsMzuJ3Jf56655LANK8omOcv5AWB+rNmYrchAceSi5wKBHKcbbqJhC
YURRfe7y0h1F8923mlTPQPoQCScZLTCORb0ZQl1GdmGwsE+SXFQOB09P1tEFdiKl
vGZZOqFAnz/N+6gr1b7SIklWb1Pu4MHuL6Iwg0XyIyyMKwaluvUU4ddFpvGB5tnW
AEgI0vYK902JKKirdy6VuQ9KY/ADYuOOJJ5Mpc1eoiYS3z8Dc0VRgNoZbtgF+Vmp
2nBaCS0vpACSNd3vgAj8uY1Pwp/GcO8CbuPD3fmNoTLvphfIentWKuZSGQZKrxrT
5cub3Wfv89gZvR3ZN5a3tjkldXv4nlOUG3+EyOYxRGmlq2a9ZmSMsdRj+oj1cKN5
WLtEb06wts4oQr2lNcBxcoUQZfU3xtUylF5CzX9EflNDDfE4mhXz7DHnPgehAzU4
O1GZaLH8OloTijDwY0DliHlv8f6O85F03HMPVejIJgyj/1D/QQm96pYRnE5TgNsF
gJKyk1PUcRQSYChM2cX2dJUH7DrW2WMKisi5Q5I8mMXIv9w5ANuqtuh9gr/gBDKa
TeLMwvQM5wcOTp1zhMjIP8TmwyeTOaFYOHWdKQP4fmDGPHJ/lg8veC6KP0VJKXrv
ZcWt6lw8DUEA5473UnMXQevJlsHd/hljB9y5gJd9xSyK+fYzHjVDGXAuzL9Laqdp
m52sxoCtjvmoRuFZoNpRNID/BM779KXnlNCJ+lgtLIs+0Um3BQ+eAWNiO2foE8wm
Je1VRXuZzMRMGs1v0WYeFgPjqfuuWqmwhzZX9yyHHcaGWTPVJEfDz8kwwI3GgNz/
thTISjB9JAeznuvGy+GKdVDW1P67AogliKrpC8mbjGyLYkxcwfXrK5ESAzSnfx62
U+q7rEYKX4VuDs3mPc5s3BJ0xMQthzHWfMwC1iWTxJCuQQCa20JSsgrrzG65qJmC
KSdavl7+TyJQ9mdMmssujLN5wdgsEORSzeuRUXLThlKnQxNz1zo8XyrwXh0ml5Hj
nOIJL6taJ8T8b06Au6w/PnSiFSx2dT8L6lDbsDDfvRCJ+VgZ5S3YBejyeewAP2VW
Y4t+TW59HDkhtaNvIn8E2iEWobWojyK54ZqPqT3yoH6Lb50ymf0AbN4MrkyVcWbL
Cp+EzF9iMX+i3iMy1DqD22AA9C1d1u5WeW0QBmhKk0C8l3YB3qDiA9ZuCIQNcaoR
CkKRf6kduNmdF909UkES8lBX1djXZj9hca2qnx3+aomVdtcvPtNU68TJ3y93H1z8
XxPklHRJj3ED09nvM9HCRVPRClWErnlm40lJFLxpfgfM+OxArr7d68hHlJu/Yqe7
MbbJqDmU95aYWk/nhRXdIIeHsIg7YLTgjz3JnN0lA89MZow2vTct/a8HUXuciMBs
Tta3TJ2/PgTCKB5z/97DS06eVWOmWXBVxbTqbSticOgiIZjriabFr7GxV9325g8Y
9AQ0WAoen1zfHqDrfbtVC3l66lE83qKG2UDvSvSQKe9OsErc+/L1i+6Ve6lW1ece
zvT4PSL4shO5/0UDJu3ryeoxVyc4+SlGo6e88tjtkVG/sukYb6OgpfU7ri2smMdC
a3wKyxbDaMHkZ5/hSUJCzXBp/qe5guIScJ6aOJpBsNYbsaWl3O/VFiWM3OWPRcBu
JstvChlE5T6wNkXcxUxlSlKN51ZFK+whdeqVXlRNQ7d2GK8jBbVTcRCCWDxrJ50t
szfGTFtlFuRujfzz62keispBc0jqfD2UCF1hVNhpBdAO+YppdM3+d0e43hCohYqY
qSizuqYmahpOMrzZDKk48vwJucDNjLWYV71wnu5ft/YXPn1J2h2WZEXP10jQzyJk
0H1DEqpN3BJ4jq27oFNoYIDXPcN+hXVHNZO94lv7XUpu8vKPYVTY8wp4kPIRmMZ+
BcXwUc6fORZ1EEytYxrGrIR/biwy1sSVeu5OIUG9ibShTkyvaRRN5U0GEMtXWrOt
5G6YekGLOp1rQsbil+Olxki9abGzWwgoIpxB1Yrqw0cEyZfLfEdKnimG4YwXPClD
xD5JpqQX+4ECUhf4m2N19g46WWWNnFgZ2RN2O2hJsYurhJA78xniFUqZYm+xoCQW
xM0Fgjp3yNEDtZZS9XvhMoDoayzsGRVzOlwcBVJEn8FSFihhD/5ekDFN+rhiTT2w
GyG6Fa338d8MA4LAWNHW+jSVEj3yzlnAKljopabaTdkILnh/+UHxkU2nQgOhI6Au
hZKln6l451osd+7GYmQ/Hqb9I4Z2ylWBgNdnYJYqfjIToi61tr2OmSeK43/eOdkB
2sJnB8qt7EuYa0gGGYd5d/pPO0JMwp+saeZdIm2aoJ5g/phGJU7zUcZD0HxRgMMY
VrQTWbGA0uMK1R84zwMfWz+zwtnMuwQt0NlhU0HSp1TwqhBpRDs0OkH9xCj2fbSM
ueBY+yezLgBFpqeqaC01eMpx6pZMbqAsWOHEgPEp4BfN3JQ7seox6fN7NoT678KA
Gu+Jwdcgdp13Csc2e83EdOr46dIGYVFrKKirO2BMMbYeXbY7KIFlpBT50eLBpGNM
KWWn5cNw7/k7JT3AtRbUvnG/jbBFvqhiHyRX6atMeBYEczGrEoG8qaNrTRoFaYwT
nHx3Am/fBCtpqAeGbzCjrC2fpOkhcAT+RVPOAOi0WACiBfGshmg9tWcmDv9IMQ3o
cWJ+x3kQAD5dPoI5qyGqkY97Hs2wvVHAuKdQwupIXOYdgJNEZBous2pbzVN9sbRK
DwfyjFS/bVeFQCrB+OU2pEd8AkrgroedssMyrx2H6TbZiYybtwcnRM+InPsOifC4
Y44e2W3dMZTwtn+tonx2g4Oyq8vzpIdPKgAPo8BfJmdvZ5vo4vs0kLeM4wAvfikL
0yI/T5uc7VUoSo/mFnCMuqPrzlNgz2hp7JqUYQRGu6/ApEMG93QIA8rcWsGGcBEd
lWs8oRDfR5uG306aTwuawO57UvdTdJd9OchIxToypWOD2s+Rz6WESCk3FlwvI34F
r0I3/DiwnPJ4gb91FT+VWp1I/8VhQYnwwaKfdYcWTpYxMWSJZlvwDWCseL/moN4Z
NAD9DuUs0eC9WuerJVrwNlj93W/w0GTlhH+c9SicUt+4oYWh9gEVDUey/aIClm5W
+cUWNvHoG4xSQm24AykjoLfFsjYJ7BSXgd3EGGWW3XVGB6VaqluLrx8HYai98lIk
ZeYbVRGyPoF47MuvTRSep/X962+73ElVaWSoStL15xOTq3MG6A+VYSjlMIOcUB9B
839yO5pxKB+ZLL0RDdxfpLIOan5TCzJQVHmaaFyDMwdCi2mklxo5i4+ppNnInQaZ
LZC76FNXar3ZzkVVrFP7orYRvpZltxzUvAi93kFeVySrIVazx3XGSAIO/72jImGH
PampnvEkIm7/L38zGRWw3gvMJTAHb5KjdjS/nZKzDu/AabHEN0rroC77toobD4We
NVnyykkBsr3XPnzCrpuQ7qox4Dks8DL4MXfgHUHELUmtE96n1fIk3SjugREpM5MN
0nGwCE2w7GmwhiQtxZN8bJ6yI31ed2i7N4WmZ/IZwY5gRsbEXKEIwuQN4xSZctaS
cTbA2Xgm7V20n48Y/EPaFAcxFKyGPZ1vz/McX0LFyD8Whbhut0Hsp7Gd9ZCb9a5Q
Gxu9smdRafQmqBHQhmvMeXWyQAbLUFPDAoGTp+pY8kxOA7uf9sTRcArNjiYheK2i
CHYBWBEkEIoD3qffaNqBdjdpXYTsY37Na6z/8FwlO1+sIASLdx95YmWJo40IY8zw
6ZpSfm5jogmyxCUz32rvsZ5DecwPv2rKVUj2CHUblC6F9O2LsqXA2jdvxR6rzXlc
wceAXdp2+ZBvFoOLDubVlUokr8x6tgGMGwt1qYSXPhLYzN71Y8BDv5SGwqowYT3r
1ur1ErO0MFdIAakvOEbaaIxoPLd3J/KXjEPrAS/xrrfl2zIefgt3D3tepaSh9gcw
wGuF1ywfJvWys0liDty6Wh3oQXYQ0kILEcXaynK/7u6K0K2VIXPptBdS+RMRy3mN
4YtvT+nXvWCuqX4PAl+AindpExGmJDscWHlOKYIeL0riHxkvVAimZjN3VhUPm62W
/7yl9a58TY0ZYBoJRwIV4F3NG98ZhEoPYEH3igVIr+t5fBjcs9/AAc4GYb8vXMen
tZUc4iKl0HRgj94PZtcmDBRfSnS5bEGElACavWr8seelcMHAe2C0YbtBwXNCR8Ox
LG3mdBniGc6Bmox9hOaEs8kNpht4adddqvZDS33zPatsjTV1L8xahlYUX4etOQVX
XnGslJ1/gtQjHC0xIT6SCsrKfQ2IgCulosdSVu75ns+n8Tqm/U/NSj9dViQO8c0u
uCq7Yjhl5AHRg1zjUJjsr5MPSaftKU3mZ77coWnRkcqsANESNRB+ftdAcKwNIWlg
E+eFbgs8cYkZWlj8OOeI/GE4R0gzWgZ4phcE5tzJgy+qGsKEhZzCjEuhxWGhtFj1
B+AGE0gFe2h8dhM3OLO/6cugT4m6JgTSIG1icCsrognEX8zycWQJaeeTa4jI7Vsk
CjbY4IOeWvyHS5/4InGxj1AzHBzuUX1bM5kQQOGu1VP3UM++A9s6YLSZJdML55Dy
Z6DF6PdkVPeUUhoajTUmjYDbC15fMdpncFXQslXAz+pN/GWXyOZx6MxUt4GXaQV6
9w9q1FnbFpZj21IxZJKrY+FtBBTSYE+uLvijhFvvb7M+n2KO1++T/5g/VcNYFQq8
RBNpwGb+ScJLiB3/SUnSrjfUJ1ijKzmFNBxOPOW6NEwNCMvgILpLZZx4/XJOdEE2
E7ohqbYCrxVx1GAKWRqKtXyRHFnLufsnl5feLjENb/AHYgdsjKsa/FqUUCjE8YN/
/VJhc4o3sU8eAFUWcnOgeBbqZyatLo1qbBFqXo6UfQ1VSbjWID+7G4QwjeGUNo/y
0gKWBDPIW6qlzwtT4uByIMddHTiJAzc3QpBPY707V3IwzmSj0wg49zL0JqKGdoSP
/ncfnjIZTZCNdQq4G3taDFTKO2yLd3b+WSktFeMLc57lQXCKeCgi5uYargoQgyba
qh3osmtefvPYjxXyHb+tO/Ksk876lDM2YtqHu+rY1bJj0cQ4/3onZNpeIHr09n/w
36HoLG/fI75jpen8QDZ2dw8sqyVobM6HwhGd+YFa/v4Rb/n0RRrqYAzGRQPyD4fU
f5S7cYIvrvTmCx2fFTY8w+WrheASzOy0rEDyzRxe33mNcEJ3bShxwzYW34wfnmhH
tNONYl9S2nblwKbMbGDY4JmOLmtpK1N2STTW5VX/9U2SND4fDjlgXXhymyj3dqoY
g0h7F23bxkezTIxRlqaOvMaT1bhaJg/AlDAArWHDoWiepmMOz3G382v8hiR8FWxR
NbOVe1oWd0MNACwAtgVwr5TnhQyNBSrUnHAolMew9chMKZY5tHFaSyuLyjrmgiYX
sINgNYlEOaYTj4zqt7eA0whBJRvBJQT8czyX0qtLkMKzk4uysmrumMQPVGbKofM6
klbsTt8wQlnZL0P1QOdaUMRgUZQYVPsxqfm1W3cP1/8tPaB+pqzt5SjgB+MUfsVG
NxLBnI1/6LGhp6HcJQ0Os7inNPr72hv9pqTmlzoj7+ZxseaE118VTOIIhGSIk43n
nJZnSuZAmUpDHX2MgFQxD50KYGFeXvX2lmnJ26Z23/AJ9UjvHZ4LbdvDWM54oYDm
V3vERyX/GV22kZCueTMFgjvBeHQDZNFUZn7BxQs7qC1eFUbpVsPn//I8CW7P1mkN
/vLrXTZayPDOZIkVFetBEzZoTQhAKQ3Pj+B3HN4eWmqCAkjLLv2aZ8wS7xW06kwn
kxiL65albQIhHxbcSgnnUy9Tx8pOXvqRAnWtrm02jctSgAKHEarNxsyy4qtotCzD
Ror7/Ov5KM0XWlRzX9CtsVff4hXCkYvd2r0J19JwXE6NO76e7NPNhdZyS4OAkXT6
EDYVCHFDb5H7Se4wccX9uU09bvk63x9j4k8zV1b2afqwGotfVsGuKNW1lBORuNUs
tyUYFYwaKWMM9WtMIH6A7qX5EU6JDTQLVe0cxcTjMWliNULUZ0H7YoDmXIrcHWKH
nGqZtmTXoKWGjXQo1NaAD8s/F0HLG7FIQ8FUV8+LD2YZ/rZkv9glB1jMT00ME43a
LhXEfa3M6mRHFKEpyOJQKRiVYQ0knVJACgl0rwgiVXygLKxUtNNPvBkgxrgRXsi7
avSoboINk5m3+IAwzYYaYHVTdSepJy/rDmth4SDIPaL/DSzsaWzbKwbWAT5luF55
vwrLzkGf1RLyQzNxprdo+78CfqcLAGhlJAdL+qxqFjgsml0mi9JZ9t6W2xAhuN3a
B7JPrqOu76tIoPHsL4p25aBcTt2tirCyzoLAKg+kFqsxEaaCcMey+UY7WqhXeFiL
ziXRPTljmoQt+BkJtzYy3tqusPDDDipb956JyPvyoauS0+ETwIzUkOSbtJ2Nvylc
mqvtfQ35Jd4lOZese5Dhjbb9RrxqE/FX3qUNNOQBtxjkdh8rb5jR/6hzRsrlyUQl
JEIxR7xh8Md3KNyjLzO8Jt5c5kpfmHfVBcFAhMCveVFVavwpu9P5EGLgWPi+Pfck
9CyKCt4b0XyvUtUoEvjqnlQ6GTKp8eEZ0M83BuaVeBgvjZK0Lo2NgGv0VHs/hIGN
V7XKI59W4ZeOcMi5sPIEZwVPzgOcpchljFNyuD+MuC+MZnfIsBZ0iV5R2PF/9cbU
7WWV1ZDayWUGVgCn+FCQAMpItn72B0gR4VZScXqSn6BFEEDkXy865LrsIUog2Pb1
ANgyVTERxSaM8LCmBj0fkoFmNdWIWRAMDlhNSQ9lRuDZpbSo6hZazlAXXFykbGCI
5Gu+spxmgKKL2T0iCY3IUAvEEqpWHYiTNGShAeFlykaApj/G6gbjgK4Gojv8rivY
iB+5k94Mzp5YQPIhci7bKGCpO8KYnVB/prZow2MNvGiv0rNrkwPv2fWpCM0rfT27
lSKvgOIHUHeEOpcyZ4u+SHUE3RtBsQOerh8yqAdotgf198XnAdwAxiX5FU+i+CSo
3Kl0WFaru+Rcr4UpcxuhE0CGXK3zK4oFOJydibt6Q7cauTSh6y4m9ZKyo63mMb5Z
1nk4p5yOSRNDU+ZE3znh2Xb0J5tVLrpL4Rtus9rm8NhmeJHAfNR2+A3oxPj56LjO
3sYJNBe/iYt9n1IdylCCWEholMh6H9Ir+I++36J0j/mcAZ8v9t28nubDbvSBHx2x
1+Wtus7UtQdWgfX5l8lL2rjZFEMpxqTOvXJg2hGx9ZZesqaNEqhf8hUcdN1StRlk
vIL73yY/cKWQOUmhpxoOFBgEGJCX/mTeeyuUgtJJh4hGUzZWpXaj+E8zhqrEwTxZ
l8NNPRb/4yL9iMyyfx/H0q9GE65ptem3owBw9uU3GbehnfJx+9ZIoLB3vRcjpy4J
PVOZRYRxXZe+KEZd9rjFhr3DIgLN1/bJlk14oxydYiH31OFZeZflIRlWzDItDRkf
eonb7qvpaF2GoSdqeA2SFkrR3FEQkNcLCXUv5mD1M3hq5AMqc/OXXi/33jW3LcPt
lua+vghh42pTfp+IxPGMhzT5khSSK0uAwPY8Zpyory/MiYKtplDHfRYTT+EQ9qR3
7gH9b1dxy0UdMvZmDx66+XqxZe2R+kaiKp4XMRHeKINZp60efgC5n4v84gchj+tV
AL5rtJVXxcBtLpMfbuQB/EkSaythXYCSFD3we25LoV0Bp18exObfSWSACTpZH9VC
Ohsw5+7mcAOJaD5o0Mf7d17wNNroJT427jSh76rNCGMcqwhsTR6mnnaenNJ919ov
wdOk5LgsfObNsPhLIudZejsJH5I17C3CvWs+5qIIKWbRoQCBk8Y2NNCxG32RI6Pk
k121bXsBl+v3zNp5Ql09/sbxD+NkNGWIDzcl9HYOUAIz1Okce35QrMn4HJiPdU18
c2zh28HxvhBKc2ZsJwlVWa4yD/3cZ1pBkeyBMInqRTSImEe3beoGwyhAy0PR8VtY
qhc4cs4aCdOvzPv1xJN+UnyndjXzNtogDZxY5M8eg8Rsgjzz21ASn7aKKaNYRGE8
kW6UywBiySKd9aRHIP3C0ifrbYGks7YuQ0Y2jFrUNDrzzWTrmxV/qKsTK5TU0JRW
mh7YTmpuFOMAIGFcsBeb9YX0VYjEPMqhSt/Zfn5h3ChZ5uJi88oQmXKm9RgncpTu
mFIKOo8M9ktusJZHTwTqjoLHZ22OMB1D7Kwb/QQvvWDnFavw69qVu+JsL2Mrewy7
bsOflbp+lTILEVXVRsIz9LeD42wFSC/BrQiwnx7AROrRp+PUH7QQn2DTVcb/4GTE
cZbxjtzwpCHYIlmehB8VY00eRDibMEcz4DujgQvHUPh/+2OW4LO43EOwWEH0tXh7
7Yj5441uaAN1l0venzJXwGM6XP8W5W8m9FCSZ4XjIxx/ECNwpfmnNCdvB+7wbWJ+
nIE0KSFGdYN9gVJ/5gpC5p3iOjmuIOhwDQnpT/Ts8xj+woUVVmsxLsjyJdJ8IoHS
g0S6diFuKtFiyp2LRbHTqX3GDHz6EDMTYRRsA8jTVAE5wv3FlZs/iQhoGPWVsnrO
kXH8qUK8HQYKi9o1iwFC7tH966Ydjucwi3LFpOnZIkiOLxNLmE82/IduQq6OU4W/
6ZvZLRP2SeRDdE/boUJPjF3VUBRPMQhs19pLR6s0GwMbsEbo6KdqIQeCGoZMS2aG
K2IVHZIiSQdPuIuoEG87hIh+9KJ5ERv95ojH9NxtPSyuf9d/Wy8IkzOpk0vL7TkG
zGrkh2sxDnsj5ytkGTW5ZqLbX/iJOHnlFy/jY2QY02R9FHNl/LKnCL+ibYeUeBFU
h+qjW/uzsuW7cZYN/dOyGRcUVveaukMESzLaAliTz2VWqOHEbWFxz+hXTG6A8g90
og7p1SILHcAYAQhQbv5HX6veZUEBoon5jHiRj3epQ29PgvIIre6p83cgNdUr33Qn
oaMFMrq/DsRMmsWdSDLRsykPq8z/66/fuTaonMIqAydOueVq5/ugtcVNgHWpHEq3
KDfJ0sopVy4i3wmoZskDZn/wns4/sL4OiVVvtRohGoVnmzxsZZxc8Dw1148HS480
sxh3Sz2z9vBkjXVLpJmx3bOK5ILP0uzylZcqSybRq99XBgrzzqmA5hJBw1NrE8Us
V9JnjJWEyQs4H9PAske6Htcjg/fzVDwhRkRZfq0m74pNbnm1IGyMrDqanhBvZBSD
lKlt74ajzvyhGPigB4Zg/8vPQKegVgQB9vXKzaEhQ1gsVLj4tpmGrx0raV6FUD3y
KVfgsl5k2MnHjTncW1+LjM9xwjcHE8jeuxfF+1ry5xaQM2CjGT+qWVlsN8Dm9MB8
0Kt09NAhs6NgdLbu6vaHT5k0suD3VkvpSedXw4nCPBKJaBBdoCGoyRuTeWXtRNs6
ob7RyzcEjM3QwjLyY7h3GwqPfzhV/VQaRz6Orm3s14YoG7YZmBNvfZyw3OimSr1R
COT/EPzvbg/Y/ONdW8g9jJ4XrSwqgLnqEKl0kYnf/NLzjXjwTr8JA0hMv4eueDAB
bP/5b9iyknc79przBblFG6hjJ/hYaBEjBgEuaGNMZJUiifEjb6HN7Nl0n3hafIjX
f74W3Cu04oVS1Qm7xHyvkI20pwytoytfxEkkU23N5ZEGJ8G16KMivMWwEYuSp7hb
Mo6D4Jk0jCQiWc2bHZxDwxWZsz99sMcsKkCkE2oUshVVtgHOeBx2FFykjy6xDP/r
iPaiZcqia3CoYbNF63w346/ZdItf68TMXQhEgW8r4eO3bOM7uQBR8Rs3dpWloUUQ
5LjCDmLhWNr9J56tBxSDQ1uAdryrEvGVDSicZvxgNPQCS2gfYIOBuChdZkXjiJy8
kQAsOMKmuWdVcf+y3hm/oouAeT+aFBbkoifSKaKKMeH+C+g2U1WpvZxTcHOErtYC
o/2FUIHn7brPYCbsHT7gPSeyocpvr+03Gv2RdJyZM7hF1cCZe7Ka3o9hZoTQGAiu
9jsyYwCaxsVHKM65L4rQc1Brl9p63vyDPlLxLKxQA8oebv653/alcvHl6MS6rMmY
YgtCZNU+4zrBAOeOqSt4hC80fu6uGZTGmNz10UKE4gjpNeQjz1r+nS/xtxYxxB8E
sLrdjun93Lj5uNBMIeJfvv44DUbBUp5YavYjbQBaI0tWSQeEwiPhO90hNxBJ27v2
oaruYg4R/kYPLItHOlobRFaTrEIEhODiYZzuqXqCSAvLdbCoGxssS8OF+y8ZFPzU
BkKgtxMfyfZylB5kJeNImW2VA9PyRKUWImIr4CApiJfniTYxYXCw+HVjYmZ990mV
xJGxDy641tauiFw+a36LkwD/BkKTy8IIuvGO0HeetrtvUWqlJjmft8rhnmIJZfcF
ujXlQao+83btxPEQxInCG/EwH4iTrgvUE24bMI4L/rvHbWRFePtq2e1tNpvzXEvg
UcfFX7riEGBCDcmtjISw3gG+BZoQFnk3GZVDp7ODE0Lsrua+rfFT5FTxX7UieApc
Du4/rOeihKS7hIJQR+7XafEj3RluPyJIWFQfMoJQdwxWvaqIMcl2G+BOBiksbsV8
38pnwQ8xA4+jTcHJ8+RMJOMqhEydPo2XzApVZcbURidIhCDrAY5tuCN7e80eHtkd
IBXvUF6wmQJbmoax3KftOfqcdOkMZFPrH7ff6ZYFid0G1cP5TAhuNJcQ99eT46XO
BCps3j5V+41MXKI4qo5lh8jX9UbH/IDt0aj+Elqjj2XKJpJSd3TmkFNpuujAzqda
SdvpfLMD/8V/1XeXcv8AyGikO+jK7XWEMEXc8IG6ATP8PrCkDILgW18zMnykJIAa
CAgoscvtRbEYjeNE26/iSOUnbzCCy4kbIfMbRWamggBFf3egnMk1Fe4GJIbWRTDi
eRwMNC04dAmfshqHeBDmeaKwzJhC/jAtTLbYpaTYBA1TDE+2H2kU89pEYNuwnuWR
atICV2+L8SMIijFXX+lLGQzsBrEaOZMdWADp1s/lawu/9P7CrKNFEM5EdHvRgZPQ
aT3rItFC1ejbD3Y7kQsiNwYp/F1srAoXdAdM0sptAvjLxnCK84miE2123I99RgZn
n10HcchjMoVC1C8SMTLTfwhO8uFmBqnSQlWyOdmuwXE4xgTJI5/t6RXm0P4pNlB/
TQ6+KvoInqzVPQzq8v6lrtG8nOkFlJEcWjSqpKGqGlWslQqU2PiPvCThFB8pKcJf
crfb1Gs2Txlrtfo8P+3c7Fwj5EVueHq8OY2ppeuTpX8L6GTF54mYcjXzdfj+uPc5
miNhXIfNzBvMc0BHmAICMUkWCGngfPkfMu875hdZN6qfu7mbBTuZfix8U9W+aH/t
cQ+HQJgdZdDDwb0JTcAcFwtSnigUD0T4yqk+EIvqEgbwn0u6Mr8AzL2VWsNIyJPP
RR2+hZAUYsdedsK2LEhp1mgqipHuo9E/pE2zdQULa8NZw6WaxZ5S1HhYOC9fakHk
BBUWG/QzcaHrnWzIRKR7dnFfvBSh9/LR1WJI2dOON5OsrkBuzjTcGHEKq+fsBM1L
Rwjji0mdSlghgTltpYXgjqn6aepufpht7cLqN2/9ol7wAtcpgyrtlblCF8MprzEk
AuI30ndViFmCbyCPliBXzdWtm/g4Qt3YuMH6yIhVhUaRw26P70VEApV3V5AkSUaB
GZnuzQCPikA+mcPClzfrlGc1yezZ6hWgNZMxnFjJ5l0AvgdGeOhW1wrlgueoeyLb
t9iPAOyYO3Jb1ByzsywTF+wczyVwmIfyUkLlr5TxyQxKpCHZW8p9TySOJom44cyv
3PGwEdlBDtlOz6wQ0paG0lTvPpGhyeMOh6r5M+BXgweK2Qrgf3l4UVwGqA5buMYF
CwAjg4gJY0MNw+IXBzra9J+0zhSmdeXBvIS13RebAV+DDDODe1DPFVqgDGRt/bZX
qWWBAiveovvwVDBKFExVjqVP3YlOVTnfE6rpTlUcQMbQM/k7i87qrB8eWaTeSzew
pUasEDVT31suW4gdFzlcngEb1JyI1d5/IeNJzZZBbg7ZPTQHpXeUVxwHH+RfOl22
mHi+O2k+C02LWkxeccD4tZN1TC0vsqiuK4D7r4TIAM0QJwOE/I0psdVH+yHE4tWo
jWqss/EptFDuOJwS8hjRQ7uBosVctLQDoslj7ZccVmWgxZzRuBRIL3vshzI3Y1tx
tOg2r8/xETU7qITnXbpD69w6+hDr/3+4wwAJrgy7PcnYMbRf87oDizY6G6EYVLy2
+CEUrqrBWw9IsFpdp+KiPo/K2T56L3JyYBPrG8g9FRFQKHiXdQKVerCKEgwzbec+
mGxlEW1cgc0m/dtEkNJYPRp/4mQW7xvmX6HMFKbE4zrokLqQ5mZi1DwKBhTtLCQS
86v09quckqip55t01O9ABDR3YbdiAPoIuR+izMSMN45dJMCwcT4Ghn2tb2OZoLtU
7ZeW1P4wkiFQifCv/GUBx+FwlC19osCmX+EfuyP/LE9+/4ApBGKjKlPBnZHEJyhp
Tpu3jdVvf0hRuaorVnpHngd4FT62N4lip+86k5bZaOKxWyxvs4dDvWA1JdSu47fC
oM5665JDJoc1aFt4vbZqvyYszXhgBld/c5Vaeny0BbyvYsxhymTqmGJnacmitZRR
RWa5ANf39N5aDrbd6i9RUbWRcBWcwAZyr4BpU7RH4B/oMwep3Bax7gB7L1FzUFTB
GR+QAK5POA6maiuSOOclvaKY8TKhTNRpr9wg1ea8G6hmIHa8unuTUzXZc5xYfHB+
erU6uY8Wilf7Z1V+StsJ+D+ifVNrlnBZHw4i7rhPiYFWcnZWcAhT9K1Ndg/u/MAH
Rqg03HPPvtZnwi7RdYCyIq5JGWWPr0RAO6e2lxzKaTeM2LY96amJunxz3ywcI9Bb
HSR7y5ak8q3x3vPj1XniNFsekN0GBTa0YX7Cz3Y8aNGBKqKXXOhWyVjASyeXQfNy
65TQgCaNjP8QquK431eoUm4oTpri4b29fo7zjHXLFnIcx/1/CbfymXuWQpW3iKT9
U+7SltZ0CAthBIL9mv0gVEY/MCrHMFz1646VOoDt7r7MDq9jzKQgiC9x7HSfL8Vh
F78hCiOXGMT052ahB0FtyQx/yHWKPFZP3Gj4jhR5JlGvqXME0X7kpcFDvM7JtyAF
sqLGZt/vOQ3OPYl/dFmt9JJT4KiLfyMRcYUtVsEq21x/xx6xQBcG0n4w8l4mU22S
11XAheKrCYYVTw8K4IiU/mKG0kI9trcbHxKdUSlzXecqmirCFsvv0TGRWMUL1fgo
VzwsDEQiYQO2sSapIgt03SN7LUF7+Jd7OMe4nTMj0eeYdTFV+smtQNaQwfzVOxss
hbzRQSaEmekT4bA5XGKCOlYoKKB2Q4GIIQJ1Ejx5XpPW3tjcPB3y+XH2idWYfudp
kFTaWlR261u1xV3QApf69ot8FlIRrNwoze4ufcqeQrPO9CQ/KDjdRclbBcGlx/7Y
NpF8GjDjnLBNoFETPFiYqdNQguYxVP+Qys5HKmdlIInUXG8kSQ3uITcJftXN9chO
hMwuhe4Kym2VvS0D3lhRCNyaXqGo/diTtPUoybRxs282hfukXJAp1DSLCt2byUTb
0rdVtpGX16l04yv+yE20Iw3GcWjUuWlLD57IuYTpkGk1UsDLL82gLvxD7TaVXIXb
9W0DZDavh8hGnOQrN0X5D9TdlMIhvg7Tm1OUnNOFs43m8EJYoqVp9l9KppFVVaS1
yBTPMXG4Tg8wOPMMID3cEZouaWv7yLx8e+dnXyTnq4lZun6eOpafYf8w9ZRbP67z
fUN8orJDUhcijalUITdv7kihhN/BNsNZ+eTKWcBTWAzZA09+26iFYSubMXp85SaQ
XOwvv9AmdyFjWb11k1gBL+zWzKwC+RaQdkQY5+86oj0gtFWGQ+bAjta5/NpiGoeJ
jragIC1Yr2BzhdmUC857WTiZ0W86kbh7fIiBa+ADoFvJdshr3TaZ1o+IWAsUDraK
bAVMQ6iNRxtHfOh9+arkd1Kn/DXYA9iPtOL49SvnyTswnLUE/G49hEVFRW+BC69t
iBrkLXPpmYlIFP9Fa6jUCdmphsimMtsIL7+mDex2Hh1aXFn/JVLim1ErJ+BsOQcw
OIcM7EBv6IXXMLS8ei1cMM1RUKADzKVunKwUEiRPfQDyNBxxuqxxudATrtD2qfQy
3CQfE/83+jDVLKreMLXtamiMT80EHpbf7CKyAwtbJJTwuTx2oRRKI6tAtyDCWTAR
aOVXs8DWxssDPaGWYMtWdnGFCcvEMRNFfRB23HpZi0SH6a0Umv8UV6w4o6DUJHrW
qyinAhXwL0FdymffghmSfTmnvKHmNGjIqdDXloTmn+c78k+a8dwj9Ea3cNW3GWlg
g23lOjFOHVhps3svsMIgR7mA+dFn+tuG4fbJZ4q6knLG3/D+8gQQdkhl801tOMsD
hKe9pKH/emrXg/RcB2RxkN96fCziKauG99bCTZVG0X5wHme7PRlhz1nwnrgIDjLu
lZMqIvuDVTlBhnM9HtmUsza7a33cO/NzozynEKkjjGwP2xrPbH+d5Pzc1/KvbQxP
pyo/rKZTBILYqfBKYAGKPBqHejMkfJOSgZ5DL59O6M7POcWgFmGFR8VdIw79gKZf
hh3Y7cE8YiX/DwV9zhCddTkS0GJ+yHwdRtdBzEssOFXlu78Q/GVvxkQuB+id66Br
bYDURpq0QeDRVhbMYTV1smF/t6t9QwrjCd7LT7IFmtWSt8/1ryc/L78RGUauKF8W
U9EFVxhM1L3gFKETBWRQvQCoFcpVTuPJnCVZwI+7lU724hWXWOLT2lv4/XqRAp8G
0PWPW0gH68ODLtiyrkH6VmK5tKivy3ANDNOaJGkHylc+jTyqvzvRK1+XFCZEOj3s
WNqbIYQu1WdxorUMzBLiIw51/FLfiySylvtOQltqH11sNJSS/hyhu1cn+Omt3QBj
IUsD2wmHt67aIMHfQsatUysER2eOqb03HtGge3MeYf6sjqx2KSu8sYBazz0XCzYV
qSN0pxy5e/8/AIw5Dj76FHCzuOBgkyBp8HQIiyD0c5rBLTkTUY3vL+wv5ecLmHzW
bMfDBeQ0DcYHO5LMHH/T16s7cGofXVyvtIfK17Plg8mCzKG7rGDH7VHfwyGCwqjX
F8GRqqdcsDIfk4C1OngAzmijpn/qfeNgqehK7dwavlvi3G/Y6lliOVNnt7UVm8cH
ElANFdnD1FUv5kUzgnxCNI9AlLCE/7q4jOeQUFdOdCKoNc3vBYdT/NIeayB1LtLG
GWsBnMG63rOYSpvqeX6HHTMpN/HosrUIGEjCgx9j0DYT9f+gwAuChPw2W6OAO4ou
mqnPSO2xFFE6vHKobXAqfQ3CPe3tb7WZk1sFErGJG2DkFtX47ZJEKKvMsFjEJ8fV
X7WG0Qu6ahQjotuuHs+VyOaobh3PESzT2YRWxaI6nd8BjEZ4LVCv8pRYOGwdaTA8
D28eewUrUdES3ifeANZ5YAcxInqN0vwearqV9FkdFs4srSNrA8EzZCS2Q1yNJSYM
zQE862foZg31wNl4h5AzGGULIaXlNPsyQy/+JYHPENt9W/eYDAGXxSYTcn2lCDd3
eB6FKVJ4PIcFdhgoWepetAstYgoqgeqNW7q3FNyb0iXoOQs7bLNB4w+yyL+mNi+C
2BCdNXbUOHZzCx+PZMUxJkJlImIL1s1fFWB9uXlyv9wgfh5+Y6O2cUnKX9BBQNPG
d1lnuangYe30iGGNaXAoh7xEt1btiTqaYEar+LS3gzGuATymS0DHXjk5chjiPIIC
OzgcsfKv3j6BYhD62gD3WV0o56FKSO+xLn0TRowajze+gVCFZV+IEszwCqd9Nwox
shfM7us8vx+shKLf5oatn5/y8ubeICOGRiQlCTROGyf2Wge8TjcXXFBdp2tuStF6
uAyfhkvV7vWvcx2O9kyXFkAs5aEH/RvgOagGgnpK5fElToOoS5hCkc6pX8iaQQ9y
F/Ulc8r1CYXgH84qKjbI+dta5n3HfzPXv2D77J6jWuclL03571H5YHHvStjm/77P
WGX7HXEJ9K3fW61lsSE5SHuD9EisX0tdsJS9ulcv9dQjTOy1BMf59/kTZUMypSEK
cm5DwRpa1Han4MLqCxj1vOifcD5dU1qXQZ6+GdBMeonROwrmhjRNQmLq8CfDV+Nb
vCytUCqWnuE2KvrA07GxDkv6HO9mfunCTykXHM8ZwNlFDiwi/q67Yy+nEYetgtL+
WkEhTzSuifWiKpMNQ/qmNfPJJOjb4jTe9RJ/q1m/7vGf/tygAeddX8L9jwJJavHy
JkIr/kDbuEi/zKGZNG5oaDkmRU+j70S29/BepuLc8JDnzEpvvASUfojaA8wsqwrX
CMpL7eX+3iKVc1zV8/UsNRtPEHJ8JWgUX4sma4t4hoeMEqGBR6C4lCZLHZXKGnya
0TdTkbxxSBJx41Jbw981Gvb7Z7i7whOCtiEUuritC2Ub1PN7+x+34teXFlcEktIo
O9qAraswn6OKj1v6gBHm942Tj4KB2T8a4OI0eC6n4JRTUmURRV0zt8uauVBFoDRo
v/AoB8jVlEqZpuquIkaYTWJZe8iREEP2lsxxFo0OL9re5VM2Y3Vux/kPlmk2qqpy
ni80U0yxU6Hapssgv3T0lfMYZkSaqcSUwr+/6YuZ8eV+ktMfZxBL4iZIRGm1MxPz
WDUo2ETsatWSTi4jjgOF6HPDgsW1qa733q3CjKH3eMPmwHC7BpQ65QM3xS4MrpNu
WDoWmuYEAirk+7n7+MMmFqb7/0BuSsNqkhHN11Bi02TZrnF2xs5pqFGJa4QCOfi7
43Ni37WoRASwnYvA5ZwIKl2upRBe/ZgTqj0L6xHvkpvhSiuf7zjtp6WfbuWQ6JPN
3qt062VeZT3WhKvolnFIZy3b/0Cvw6URZYz8MiJGhHfanEIiKxNdkielEeVgzfJF
1dBb6YReIiYZyRMyuD0G/nYnzN/s7c/EsssYjOC3F01I0xiYgQSahtOzOZKCEcsp
2eeENPXCyAiGlAXyH+VDfy8QCeOnf1JM4GYZxO/1T8K4dmZ4PfmnjceBD1OOD86m
+d64kjk/6HD1SqOUdNQoD4iF70H2nYMKa96Shrn9PtAG/3YwS4vuWFYr5hILCV2+
WYHMEZHdRoVPSkPMrKvUsq0MkNd1j+X780DqldzqOH8Ltvq14ftgI9GIz+eUiy1g
W2ktmolvexeevBk92z+eAjKW9YIQ702uswhQIQQLxOPg20xlamgb4GYRat2ONzcF
wBSv+FFpBYhos7nEoKxvCxv79j0LSi9wLrbVTnvtgJkgiG2DoMdVwUZt/1sGQJ7I
S8P79EMbcyDJY4dRcqXfqasHBfjg5a/8rraHEKP6BbxvRLDm+mMYcbBSGqYH7JsM
ou+ujIW0H7OjtKzI3Gw7DW9ukrH+PqTK0WQaORmSvsm2cLGX4DHeyQCCNEc1qLg5
57y+g6QwIUAT0XQbx3to3G8qIsdqshIPNaysB+8wCxG16g2b3ekmHbktM8frAuPP
HG7vsMfnb+4uzTpNo/80K1esWIQD4S6dkzHXALHjqI8kDy6lYVxz2trDsKkz9Q/y
X9ZrZsw2s5BP5EQ5TbuIyLU2uph425+tL0xWWNx0Swk/KE3cjk1q/DIZ8YrF5P9t
cIFeUB+yB8fyDtKYHiZYpTE1jhfWWJkH28DTx0rHHaltxrCx6a6ZYac3Cv56ji1z
0O7hvwyJPDwCNfQoUW6+a/TYMTrc4d2R/RIjbsS3PdHvnK3SLEnSLc0f16ZGlsbd
6l2Cu2eiFH1N9Cnamw+snHEjqg8tF40grx6+1CdNmDt4L5JObXDg5nJX/cZmuweW
YnFucThaj9NEK46fci3LIIOStA12w4g48BPebWbQ6dUQFQ8ivRT98AxawJ5cNabE
edupJLdD4Rb7yDDEii6k9FJRORyXD6Lt4hNAxWirhivKiduSQP6q5ZAngszkHxGx
Fih1MUtf12+6cyyVuyorBx4MyxjoAPoZ7wD3iNd4nVLIJyZATh84iARQpEpmGnjI
knW/vDhqW7J/pKHFJJn+sMJ0Ek53hx3uigIZW10QjetzGb8f00FjPJno6zv4rjaO
g5WNBmWoc5zasqhsWBPEcXTYUwhlYykZxHqSKT8Xeh6rMPByoco+KQoxgAhGbCx+
uscxpCDt/DD8qxRN4AP0qi9AVzSjWEBY3uU6ZYxFKOH+YS5xz92cqth4G6yzRboV
FlLGowPfFzIRd6FC6bhX/JV1/BI1RaWJahLyrMA5CBA7s9WmbgVThxcsyruHCgUZ
usZFIwyw100HRWpOdqxnFTFzNrgznjsJb1VaJfpbbsLcxJeH+ZfEb1+w6bvv3rOu
qTwK26BWaeENmmeqtHNogR5RQ8ldNs5LaP3Vuh8HLmE5+0GkXb5blRvkG5ozeMMs
trcYXN2qdbp+T/jYJSES16LyoOKQ6TYxTHsK+DKtAde9BbDtAOzi3VXs0ZgpIv+v
F4kGxjGXoSX7du6P0DBrSd0j6W7BcCfMSJn3OwvUj1Zk3ojxEIxR/2VQGV3J7SQP
hljqTZS6Ru7HJGH5MAflru/X9AhYGJCTykI/CNv5IRoaS1DryGud4Xo9Az94Ip/u
RqzHNJBzqquUYX5QUEgeft1JAitpHVKysfB3d3lOaFduVi2+tt25EYdvFUaK0K1o
TA+7f4FZhbUSPN7XvcSJGTDMv/XacTI0H/gkOwnagI0cLTwH5P4sU/Se9iycyLtY
8vXKwO8V6+mYMHZLiq8sV3opReOn7YFFTqIb+88W/xuig5dqSFOtvWc5PoMCq7rw
nqldS51UdR/l9vVl7m1Q+0iwgKPS3cSbutiSj+1VsBb8e+EQDcyd6vgZmllFUSk8
otDcSCpZuTMBlJ6XiXJLp6EYv+bti/piol4RnHzNDwPQTTTUzs5wfGDoqD3wKEBp
ibNOFHEtJrEc2RMxGMOobi/Vn1fsHHdmedYepktgoZJjn7zbvhZAGoO22nbuwbQP
OPOgpJcN4+zP5yR8WSTZJLHUR3R763h3oiY961uyzkw2qiX0TkTtHN5tA6EyPxmC
CFseoP9bhIjffYePU9PG9530WtZ1U8bNHOkwT9HXJUPpCyPWC3hbR8/DsvPrx2Gt
cR5NG3OHZOAkvpHrGoVS5B0DNsiwS/kngE8CYWyYmguOkvdFaprXRchKoQ4QtXS2
vS5o2G0Be4KylEwRY2oTuM/srJtqSHcuT3y5ZFzrPyG65/RyAh58OxIAQtC4/+Yo
qQU9ix0zfPtzW2mp3OvVznk7fl9xULJuIf2LKrUxCpm44UnWmo6gLPZgoxj3TXjo
jAtWTC5X7VdKk1aVKD0H0bMjfBkoMlNl3IY22HB86mYsXvC3i+YTbsafP7jFlctp
pp49XmWLcg6Pu0VwVyXmben4oAWvZqky0JtEX776ZAx/vFVA4BYwxgPstjLuoe9A
2/vXUAwKNBOoa2TNHxj7P4ptY3NwcF2CS7y97Ff8P86eOM7Gq2Ym6yVB4BTHnrUD
JSxyXhncpw+oQktHAX5YP16GuatJzv02NT6w20jnE4pEnO554oRT3twp3belgAzD
6WpmwzZV1X5sNlBgiAzUtPE53XksO3SrEWVoFe5UwV3LkyZvNgh9LJVHBnNmt+wn
+BtlAW7q5Gdr87wnBbl0eYgETcZFj6DV63z8TRggk/RG05F1t5pLxTSu9/J+yiBQ
8Gxi+HGtKhc5GoqGDx3t4fH3aDUd4wWuFGXnA4NKvpQrkUb45iCDn33xwlAuPdBj
pNyE29hg3Cj0q0OFh6c8VC6piZPU8t/+J2uwy1cxER4g7AxSvu0gWKrguDb/2rkn
NbLPipR8y3rgO6tCa8uOy2GrinW16tNLyqS1NskM6LzUGpeoTsqzpI1QaAVS2JbT
rVJGwzG0tjEcaS27+wIjAOVn8l9Tibhq/xmmOeyQkGfsIkrI8ZXmgnUzvr1b43Wf
gWRwoIvagD7F50jUhWo/nJeLFjQkHMslCdZ5TlkLRI1PtdLyUFzbrqQ6SSfPLGVE
cBfnd1mzLJ6tnYMOrUUQpDSDbaKi9lcn452d34jqtQa0zX72TNGeD3YQoQoYIQJY
MWsgr7yXeOA0MFkjHNiR1hjPa07HqLdtc6POaj2QecXEoZtk8rY9GK/+5vbj5N+K
QqJY0Og5CX3ou0c7BRzO9KMS72RNAtVPpc4b0kNqQGCfb6lk5laorGTkEQf5Hidl
x0NG4mtClsttPq2XeP9bwPMavN4nrgapq8yHZq0IpiKdUtnTwo4AFAHbSfbS4CcF
Ofzyf1oQXqaM76pj/M1S1lp1AN5vQkXqB0/syQ8DjIGOdckcEO5Y9JvrAl/r43wp
XQY2eDLsxjmPlkt8DXI966zyxsf6YggB3dHdQLgTpLifP3PIRhChNVwV1TcetrVU
6MwAM3wSsA7dfCXm00h/6WFQlgYdEszc9Mks1EYidv7PnB2XRnAl+5OShRCcEX1V
frNC/h5msMZaIov7YMUyuV50opP3UPo8eH3f0PSlowgnTQYF2Tg3dkZ7zxEEI/eA
bCNDudDaqfDfaJVpyQAzSDUIFiHtYJa1tqieJeA6nOC4NILjBpf/lCPZgUDRcf7L
7VBg1WTv+AoR4MgaoFZ3VV+VmEoJTNBTCEIBJbbG8lJypXG9Ua460YSZfgrrjDg1
DD4ohBsDoC+l+A6zqYTyg9oc83MjgYZdmxM4srOx8YlzvA9SVgqEjcg5uUpBu0rW
Xh7/BIcou15Qj/HpaAVKBvdcdbHieGLpXookaetKfio58O+NfSqPhEX0MNBeg7hc
uTiMvWxz7a5Vq6jqGL/RQ/uWS+7gvYK4mSdRBVeevDMeospqeTvtNo3wEyTCTAKY
W2TPZi5svfNVFTRiz1p1StABpLaKoRXolGr/ysl+Nh+ecxnWBN6UdgmOXqVf2ACA
gfTBmnzBPf6hBCRRLGqtNT4bY1SczZt0oes09WKl5/uohMv8fCOalLWIt99VrG5e
UnpK/vxOHvN6Pp0TsxFIH4o/W0nWF2nua5UfBGgSRkxVmcXahqBgQhXtYBEtFROs
ezjjRUN1RUeWR7d9Z6oRyQU6QJFgHKZ7GPOW/5Um0fsfxqIx5xYpPBKybljsLHaj
lGF8HFhM4a97lVnfD9AaKoSSxfO5YkxJkf8CDjvgYmy3ecIxlJdhY1RJZHpj+Uid
r8aiqZmap/b/GcbRMBq4LDFETFt2ajmMbQLS5W8RuTMwgkMRMmHhl0/zGnaemYP8
vR5Q5gZf1asNSm0xSjFFGbs5PJu98iaRI6xZjE7XbMCLFIvGzcZijMHnLYCiH/mV
Loq0YRTNFZ1WdKHyRtDGUhZGO1+ZaxEbY4TffCxcw2vRVo+vnvOFn27XelOSP/RX
Qzggv9gufuSQqP1/NcfUc6w36Uw0ePPIaPVUXyS8u1MEuOePZpLV+LHpR3coF0/o
zkVi7Tb4yAdMPt1rEQZNZiKwJZcclmXpoeTRgjgYZK9YtC45rXaazY4w0aNEEVbM
FfQHSnHesGpS0Ph1iJyu5O/rlCj4rvOzThba9Eru7bVnvWOoQ8nnPIgP2M889qC0
wtWOtsaFDqntFvOmZ2cAFPB0k16DSPD7CgiS3hAUSItr47g8hvf+K5bJBS/PXOhL
JVV7uiNGIzQONwBykvKfDoKAPLJgFR8NvjW+OOwnmzFJQ9FbfxNoCeglSSIjyAFR
pr3LzAZjOl12WV5qs49D2+5ynpjiNzCZBFcoYbsNYb8+WFXciXHTkQQgi7KT3xg0
F/87BcgeqUUe+4hYO8baAGKXkh40qhCijHKbDoaK90qp2gcotqPhyfiVsz3h83M1
hUCjR3oqhIMJbIRiltoRuN5Xjhb+MGoCxhifVpqkN8T5K2q51jN6FG3yn+HmbajG
0XTgq92pkFnvCyLvBVADUJDIzSRJHS4rLIHbwIbyuYVuAI2DkKxZfB4PTnaXkJip
RoFraMpjTnolRTJPfXFGbknN1vCZsgAoFREyqkqog1Y02NBci3Lj9Mb+UsVxtuOa
dxzuOp/lzeREZbUUjIqydRgSje+JpxRb2epR2wLnVt16/CWHj0MWTXA4Vr60i/4B
D16PkRAC1nVj8w500b5l7A9VggusF7Jw7YyaXp9XPXfNzCF0QAQgUWT0dIPwUCRp
ADQaOZiAiN/l6E+fXaHWOguspRjcl0ACX/Az6PeTfr6I17z4ZA2jTa5NiChn4+0i
l+DrM8WTowQq90ieoR35UVtPrehb7Oqo4eE3M+dUpLL0VHDZ5Nh6U/BO5TVx/0bS
IDezL+/ouX0L9r41jqRT+IPus9+wevoAb3chskh6zikwqJC9Aa2WrdMa8j7Fiq93
G8nre88688CDEIc4OyyxEnRTDdFpHiv+7ltpQieKx7D5eXEAq00j1HFSy+2E6R4R
fyOlwxRMHz9ZylPCcl9S768yYC8zoFSil8M0OlgnhJ2ef60xe0GHWScPa9/ilYC9
MnyV7YztvNnynH4nZk25XhRgjoTTfak8JMRYWZLGBhg8ezv5IQzKFYj1707OVZHR
ZNB1v8kNdnOhV89NTiakCkFnoOieh70VaPGjOP6BmI98pULu4QCj0NYncoGNB8kP
hVgkfu6d08JX4btThodYcH34vn4Ldm6CxHdcHI3hpIIOkvlbRcwcDvt50XWRQbdZ
GVu6L7/UGmL3w7ud2rOtkiRH5K2WHA82PjIXVU435vFadEviDrD1rSBr4PHtuAhd
wKxkFWawqGbi/GTacSEGERCu5eLrXAfZrFjqi0XntEVDwMuv4Jme7ZKPoUyHEunS
jXt60MWi+ZAvUGenS2uBVyoSoJne4aYtfZ8Bu+RAYcSw7HPCBlp56OQXlu6OHDL1
CxVsxyAbHismvQQduBCe2Pb7P5WwiDh+F0hrWWq/t0XSDJVxUcUzcnACK4UZtXtS
TxvQqMc1q6kFA6YJXqPIySmotHwj23kot0TwJjL1uPZgsFHYPbZqCVuXFaLJYKst
7aAjr08SQoyl0BOpDuqCgwBin6JTq8/CXziqXQF5bYYjC7DN13yCEcKskl4qSvL5
9GiSSTSv1G53L78dA1S9m/ruDeBen/CbpoFr965aNmrBdInjtL2dSO23K2i9YKW+
mJRjEFmZbZDLkYd/LLkZRh0NVUs26NJiizIpBiyaNhUjhar4Uyz5zdZvbZSyPYtp
q+itFj0Dr+VkPPtYn18YUm/o9KkIBXCi4a9KDJhqtJXPPgex4TNcMvXPc8d8bbvg
IckykKCs7HDpOj6ps7UXfgLdalhe1NnbU1l/BUwVlHNc3wr/rWcaGuVG5TosoI06
oxImuzjjFfNw80q2MwhKLkOStHCswFBkPpLyknBJiQTgQ228N+QhTGjrt7Zkd7dt
eyB7JBejwHsp0hgr2hxJu+7OdllVa3x/Gr9LVmaVoEqCjW7GmXaHlP6JLl8DvDBc
2U+BNCY+JvQT0gJcDNbNaj8buH5o9w6mwiI/DRG/hddmnq3JYOLOmyMgogYxNKea
8QIb5cnjdz7I4RAYOzTrCAZYO/z9JBxEZZ/iCe/t7MUF3VxSMJrVKEgqS6NVxdE4
alpHUsGjYD3mSEXuKzF9PBtZQaZgog+KK7H+QnM0L9PaZ+pKAxa28dNHW3yonsW/
gWoyMkmsIKKAOy8pYaGSBuc9c/mOmkr7MZpQHRnOZqX/BVlCw91joqZ2Uz2MxT07
34wzVfqSIN1Kua27UdM62ZTCN8RjXlCbTlEeFYVsubUbJ8shGuZ3anyHozqe1TZL
qUlKdQzDd1wd+Osv2BBOWZ9m828Zk6K5i68/ZrS0cf/LYqtBurSbGM3XGQfkOU21
jHOsZGCspbcRcyM7my37FL1iLcGJ2XcxNuRQJIjk3BecbYyVA5FNQlWGzuAEmujK
662CtfSsxby6jZYhP5Rde0FmJffT9SePdTFcuVcd37JHCF8eppQawqAkTh6SEDjb
RzKLYzzvIIn8WyLK1kPNcXUye7mSd6IXlKFcXr1dxY+I2KNd4ToKmOgbb2mY+PlB
6hBs55oEeTWo2v5jPFeYHXJrlREeeBlfMXwqT7u222efRFIb76DQdfIoMpuzmtTE
CSwBli00EpLS2nYaSeolTmZUuIS4ADAoOkBlEuBt3QyN1sngI1kTIautkmvlQ28h
F8QyVB6hfbOu2KzBj97CEl9NAaVDDvgMuOn2emuKPGtPDQfyDzQqe8C3d0WThyfP
RcOvcS78WT0eWz4+UhXCxSPnnMfF0b/U8Vq5Ki116mCvuz2Nmdq3C8YBpoXaGQhY
L+bQmPbC+rMJw+G1YMwhn1J7rLQm2ZKhOic7dGEMwXKQPlAfYanPH6pBJDi3UvEz
rxLF5y8onG1S+2Q17MOY/Hvth3YWLBq6R3xBCMASWU9C4kQs7ROUsLd2VgBAH2HY
3dEyL7RzLdQrreM2Oc5cHEJuClanmZs2Szgc+KoqsQ0jPxiR0+Kt63NKmHRVB7OA
oAxiUFK4qKbkFyozQm7KvtGLRJkydCLzGuBqjh4vaIcSdLoM0x/m67/RoVeQxnGU
rEE8ebaN/TdMboQTACZ+/VigNDFNJmIqeyf7i0ZvxKZxxYBP1ZQPcpZIHOTpWkxe
7KW6Xo+yP6i2OiFlRb9RApmonhFQlDNSgk2Kq8jyFHj9GBAGKu82ktcAAYiYanVS
jPnOB9q+uzUgzkPh1BNeu8fXq7FH9z/ttS+xc9j1XFqzWnMhzeAaHD39bsSJsr8v
sainoaLDIom7/RPrXVa9GdPEL9TOlSieOAN1Be2Ix7jozIhYg3NTG3SFm5sEeEiL
+gAzhg6SyL5eN2WH3u6WVfpMfyHo6uzBC6zksTCevoV8kCD5Z8mC2TRDNFeZBXF3
C8K7VU+CRTAN6ISbmtDNG1e7rpL1t7ZBlNcQaHLoiH3fEnDCkaG1U4ipLRrWSo5n
IS2u2XmhOQdRecPFTFmFlGxud2/jdcL6+1oX98W7RZQSis52FAVmeoK6bL39bgyW
e6HmLl8uZeXO9DcsZ6R62YplggM3SiMKMsVUY2odXEz8EdrwmdqUaV0Q+zxmZVWU
fc9T9TsTiJR/d1PxC2E+1BbOoOf8EoyhxmxApoGAoJygNJMgLSG4ybD++kGAF+qq
1WHW22Y9InIhkSHCJRZy6huKuk5p+bZ0OZL8XEoG6oNjd3LohIgWW6HHREhFH0Cp
dm6dq7elcYupDIEjOk4iKNB082k0Iwyhy5kCAvS4k7cNBOPbSKv0gK5X6desAhzu
b0WWhke09YXleNm7t6dpL8oG/uGtCYjfQEB2QYF19ZkRyccKkySZjPMhOE9SnB7q
xKh06kmG2DDn6t3dubxHfhJCxcSVt2gEUCuZ7vgpbwK2u/bJMJQfeidlRRqoa6Cx
9zsySqeGkkgfKjvfywbkGQ51yStVzs3MNUQwEIhKCHilb2C0jyNo2Ih6aYDPv4oR
SJGqSFpreluRJTxh3KdgRfq9rmCeLAXTaE78led1okP6lVzusr5b0FXUk26UJ4WL
cgNzWzGn6R2TZNvtlq8E5d2gXUxwM3gCpz36taPt+AOO//jsbF9qnOhRmR23oz8J
ACh2BT6BYSEOOg6i5g0GJ53jOsgWOZHvum+rlROSI4nOTsulhhRoPGDnDpKjIwrt
sZ7lE7Tk5vpRWREP8n3PlVEmjgKnAqrdci7DbMwgwiRpEgXN+zIuGYO/WfkksWGc
05ONPipFY3p442tJkCdQ0UCa29Y5CxiiMyxsxkPzeLzegF6ubCcwr/TTyrV3o+/w
Ref6yzwjVZXUczb6XjAuDVi2pxg8j962wFLXuglEOXNy8h3FyQcIUHWPgf5HQTLQ
RVNszrNDyBzvZJsn1q2oCTCUAX3LknQMxwPP6945XEVAhL/k0eci+oM6jE/Hb+zp
xTgFGmAFIU1BX299NIX7CgbrIFFew4qPhRSI8fKoMLqEISjPuvTylkPifwD0RQ0l
zbwDlE58Le8N7l/xvvBKj4UuMTuQ7/gB43KpLfloGm7tsTFLjvSc4NfHPfv3F6An
v+TFpbHd5gF+6PV2G9ECGV94FWWCP/Cs5xe+Yp4nbMXGXh1yNt/01sWrN+EJU+H1
Aj4/nGWn6jJiBrVpWWY2BKp+6fUqOg8fTrqzyIqsYVZQjJ6Cv7Q5J2HYqhC+9Nfu
ysyQh9yOEr2e3BQo0K2AYb7/N7BrtsXeXrFyN6pXSDDAYYs+Ly63pHiiVx0MWmP5
4h5nlvkGRqzzK8iT+e1a1+Uo0YLuRCziMEwlmJ3C+2sHnQyY4Slxd/E8LK4nGTdq
NqjlvxuGzgz+3izMJn6PzFe1865QEfwat1HRS55ueI0hjfdXLOt23/J+fUjlOMTT
4q6mlNHPrF7boplmez66OGyYBw0X3UZiibbOGuufGywlaXAF1pXiRUhgxBADzpNL
K20H2sd7BfyZK4BHCPHurDzVJsTGJndwCUnVJKg2bna7Cxf4RG4W0bUPDrfzRJMc
W8j8bEyxn3CMIUD5y7oZX3JL0FACxZYe0AA2eq+x1zSlRQuxRGZaPAfisoZ4XMov
R8Exho7Lq0pDV1fa5Ti9VYxS5ul3CmfCGIZUnSvaa7b85SWbM/o3UmetSFH3y228
mFiljcRyv9sfk+d7AYPJpJ5FeF2jqAs2Yi+XVXAeXt+hznDOsfyItZNoa3agyUT6
S9g/xyii0BjfVYqWDkXk58uwc2vgoCojyhtraalIfEIH58xuM4q5ilyfXurCimzL
rjrwaNzCmtl8XKhGja2Y2gHPt+zL1GSAJXEmTq2wuOvx4Pu9/dM48lNrouZ1n7We
sJoQgG/YVjpJVqdZPp4GTiUU8G9NPgTjvESQ3Gd/xXCPng5LiGGevoKxeiqsFrmn
v3mvtNNBxhBoS7CBJ9p1ikKKIz2UgLMycB5AhVbd01DTQi8ErZEJyXkYpHb7YCGd
c5THKekesWSutadW1OVxmDoWKGdKiXzVEJX9TqW93VOrW2i4B50tFa9gPHIFaKlk
Mv6NrmX90jdmevddOQlG07yjJYuLEajdE3PTzkkAk/nbYtohBjIpcF/oTJy+wc7k
rxYarOrXEaiD1zsdEseJC8JFyFqSduZ5ejBOoEooR+esWa+KwbphUl9U/Ih+8I7+
5n7Z9OtsTafq107eeGa4BaH/1P5NJYhhT9ZaPqmvUTRJvu8t/GSyekh+cZLLHySj
/lX8cPJ6QS1PKqk8DzyZqZxTbYGiYAYn3otmI/Y/U7hXtlgzGbAqvOwk5pTwjN3J
aDzOjOOWIzRbauer94+I6NyOzPs/cAGGLcTMOkrjVL1bSs2AAwS67yAyr07C52cu
PdKQZ6dXCP5gtzzpgJo5WiLEeV0S+vD5PA6EbRQwEEGlfGWPNdK7vk+CfVi0lYdz
bSyoTf7mNAyM7BuYDTKSVmTDdTJveawKQU/pR/9VR/acJSa4V8IZRqzbDvQYX/QY
cOhTMww6eFBe/d2tDWx7WzCrX2mg7AhpuzWL+M5iqoo3TaIDaXJFvQaoBcpzYX9d
nFmwaMO8tU8G8QPJHVCEA8MOAC3kgwBwJd/JKOOJSJFdxa/KoQVIBCAsWHgmdxXQ
7GfgoQwZ5wwk6IMBR8T0t6jhbScVG7uNp+P5cfiz1Juw9yb3kMkB8dHceM3b4BjL
P9CcLmUcgEieHuckFcoKppB9xbQaADNCFl1LpXUiCnSWGsidiZihsWEld1JTS0x6
ceS1h5QpKYvH9/HRqKqwVEucUqw5/qbtSXsova2JfQb/s9lJiJ8OPrGs/gfLrhFP
qOfoUrA8FUlNs9pmeGJsc4G45Sa6wmtY3dphLK6nsqNbG3uy7hHBPm6FVJwW05K7
bUr8u2EB1F7m8+gXWqTSol/6LhxOvLwDENR0U5UlrW65ASwWvnUt5KLAJpJQ3cou
6bv1B/hQxiBSf3LE+Cf4KvciXKzbnxLiCJXaH6BC3sCB0UJJbfPLkHoBge+apOkM
j7DKR+MrhBoAcNNxdc4m0YtPTrovJOlvs6zf72d4bzqGXFRHSPf4CJrI85y3m8ih
PySRPvA3OMBDdb0vgplpMym3XC05RAY2C4uh0JHD4ryZmZAthVTLHA+bdqR6kVHb
pf9Li33LtI+jMMkRWLk7M/8T6abLBDteyPA4Yti+/HZo7HGH7kJZ+Z7K4nM1CoZB
Gwpevdnf6EQ+LKGbcBGIuS30xW9othRl9N4n7I03MWBRWhbz1Fu2uM9a/v/pSfE4
5dh8S+oJvFs/P6+c5X6oyPdrQ1N9BjVTxsgUUcud2rt/9lMzRqHO8vcxM2EvuuNN
P7FvCLLk2uKsQW/UnEsnbdRw7hgDFYwihT5jV7USFh8loPdq1uPjvyn2M5ohR0YA
+LsyLY1JHJqBE/iPU1k7jvd1jEBP5cKh4v2bUbq/hF/THlyev8LB2u5/Yxaz2foR
eN1yiD4r/TAiWF0lsmkDgCadG9jz2vO/A1zqB1Wv3+yybnt4oEepsFpDzkR/g0Dm
l1JJSMR5wBePmcso924pJfz4vSnIjhjZJo6mc4ElYLuF5or7ZTX5aM6tgRRmrf8s
M1JL2lS8zvzRsM8TwR9XUQ/EVGB2PxgOdsgpUPI4CGRa/vpoDcdRS25IrbILtXDs
Llft0XEzfJ0yGtr7DtPlCrbmy1syXXEmEBdwJqm3bTOc85tpUGKpmRJcZNu0EmQr
ZYqAz/WQBR/iqdKa5mTy/R6K8q9LLek1AxL/vl1ZKKkIFbVeceZZkIh7rlzMXb2C
0W5F2UYs0OImqi9zslI0A0ZwL4Vmf1ChO19Ab4xzcQctGYzHZZSu1zwb0tptjgbx
nvlvHIaHZV1RX7FQnWy2Vl0szsQWcgGbDV2jM4Ws9lalCR4SkoyUcW/lPXYHBrpS
h1XqZGdhQD9DM5vRvehkz9YreEwfVWSwwIKcKIs2oQBVO95m7uVevJ1E3Cs7GNV8
TUSymslP3pEPs7/XnE3QuLYkrFd14/jGXgAwf1OwIJqRMn1TLjYXuHfUitzoedVr
OGCpoJrlgb2gOEz9soL5Et3Us1YU7FxV1muYbiyk2aZQMro5PT7A5h3ALaEs8qDs
nycA/7ffkIXK3CPaYM9Pqr5F96Lgli4I1VBL34DV5127Jk8UcRLZSbTsJxyx3b0n
OoUa7O2R0AnJqly/nRKgxXPXPggyBb7y9YJkK/mqUngBY52BhWoE+fvH9O0/UpAb
Y3XysrMJYx/DCCA2m7FoRPU+bFHxmcyFn6dXj+VqGLh1P0sneQJnRXz8rDrI/imR
UebiFqGDC5uYiUz4paWbvlGibvIP9zl6l7q/HaRlBMxjN1oySlEP5RdFxeA2zkcO
AGMnZ6y/YrUi1se7YBLRH0K+0cnZ+qtKy0xsoli6IC186NbVxRlOfqBNaXNz7jDS
1KwgPGx5Aw/oOm6OZQSpA7bzNfrs06YplQvJUtGIUvONWRBMcl2l7gLy/Fi87IZl
anYnnwr15PD0wtsB2RQUHdsgTXcsGCI9BnRxqWLrM9COCwmRzFpTZQuGPQKFGcKS
1WDIqw18Ww0l7/Ra+X3rpezr/XKQWfuTETNG3PxCx/Oq/kbkwggc7bX++eF0E95i
kqF30YCt5EiPAL6F55XD0FS2HoNRebHNZxqYDO+kzVnsKX2YTt0u2r46jy5EGzXo
0iclBfgE+x/6XJqLS91gZDVIZ+Q+24YvUfpFb8scO7qlwtMOsNKUBVAGQ1qtH4kU
GX/+P29TIlj7BC72bpcu1zA0qqWj5TADF4Yr+gd2WwHdcYEMPTmBayY62aL0mpSL
I4qIcMihxpmoRdjMMG1nPZnhpfnm4VPiCdrYtACAL490myb60CnhxVmKP8d88vMd
53hW/th/SQsu9E0gZ7PqJNuE1R9cBJ5fRKUEcd9nrp7DWj4POYHUAVI0+cEX+5np
kMKy/mekqkSHIDTnlg1bbV/kH1ZjRZd7QA/qPjqv3B2XfMM8moqqNZDyMFnrmTOy
TqCTG65qqkIObH1w6LtR/dh/m9vxRd+ELtj6jrKd2RmoT5OswFvycC8EO57v3PPI
7XqePnMxP5Xu3L/+pGzl4XAjD058TAADINdlYPUVIoQO8xgEGHlNa2zaXqvPPNpy
nvffN/vkfv1B73DR8j9NPZfWDxkmkzvkBUNi2GEoGhtZpjdh6s8+bA0nHKavTPtY
9OW7n4sa1C/WQ7uraqDFRMucgMSTh2xwPshARsFWdbefwpPV27Deo/WsyR9Skz27
cETWC/SC3ngGf2JwDmWebCweZi7M3upVVqZEPClVamMxWdkxB/DxIm21jb1zajNP
19zM1CsYwSrED0s7z0alyipLYgX0va/wm/0yTQCh8WoTOKOQ7Q/ntHDZW+4CwD23
EkRiGjc4LSaJw1IHOrd8r7GG4T+AlzNCWlpnptihpYgSNr2Num/ZDYGMZgpTN8O5
b/esz31sf+O4bNN7RraeJ7oG+vVpNckCi6Bth/p1xI/iiL8ik9tMKqujuLs9DwQD
HErQKc6axaqDU6yvpRvv69jBkvyooZzO5uIcctpDnfJv4XD8doc7BeA7TqSmZnZn
8krAMYuNow4UbhOgRxLr3oEBXsfmSfH1ym7/R2z66tp+9Fz56X4NAgP8FK1DH2Pm
dLGbIPYqgVqSAVORPGUJAvW8J5v2FCiP45RVIj/HKm5Y/ZUGCIk2m1c3fIlXFQqx
LvgEqIqYul+3ZjmsAPfvbUfE7M8a7fs3GMkwnXzABAqNh0+IDIZJeowY4hfbP/o3
AIuIkgB1gDVANHZuy/gDKN7hEANIDNNj1PySyr7TFJVXq4uPW5BA50+juMH4Nahn
/co4zHoZIw8PtFUewxjoAORNhO1G75X7wMuPJDBj6Ofh0l3y4rIwEM2UeRp+BoZ5
G4MqWnisWg05Cm3Ih5aN7Mc9uA2U3qiObShh4UzrpZMDS4O/QQaMe9rmj5k+iVDT
tqwqQSpaNBneAxCASMr7NT5bVsR2DBOkTEs6ufqhuHTkRITm88Xf2do+d3FkPpmY
RyxKbIyicK/ozrbUCR06KvAymMO6NiT+H4dSSq0nK0FCl/0NB91e73rS8EoUstLz
qABKVSibCy9H4RbneVHhqnTZ5xuLA0ihJW4KcYyMxpTMUrCs7Zdr2vaATuPhX2bu
O1hIxPwrkzVDUOowscPhYDsUiwc0191N/MAFHw0cqpGMR3vxAHbspi2V2nkg8U8Q
RFPE32zoV6fvKVZU3zQVx8ZjR3u7xmI1vGIQFRQiftPwNzLugqAiH1w7SBsuxC2/
aBotFMS7mVRVtcW36UUrm+foC2sbg4B6WBfEs5xP7KUfRJxhIwe4qVpwqa6pdK7Y
h6N5ekNUPnZ7YaH+0lJ5ncg9tKdisOpgGM97rlKuWIFuTpO1Pwl/I/s8qQkAAgsN
c56cJ15crXdOZNAwOEfC/MLuBP4GGXzYtiL513ppjhFvZfJxCS36047Ouy//JpiI
9p8WbV0PnUb/9vWLbavJ7CV6fbcxR1678pPkUKwXe2fAXLrVmUlbxwDabhAFAiUt
TDmCGf5oFu8ZfP+Pd9eXaISLWq8xDr+ysUt2rf9mQD5TpkfMpcTm00niJThT9H55
YEC3fVw+A+mgZc1E8rUFR9P7cSSW4GI691h75+miOFfZNJg56Ew1dLwiNJk1b9v2
DiwuzGRdawbRA2XSf3uoIq6LO8r7P1yRMuwjZTYIHnFdoqVRJeCcR3fn0QYmj/xh
BvrdkrmrG23hWQUC3cSRyDAV6alvyR5ZqnBr+gTBiekZENnYptd9xJq4sWn4P/wf
a+FZGlvvt55cZE9dY7Cb82uyKchSkM4dv26KW00U+y8t02QH8XLX7JONU+zrw/FR
o5Zg6ut+noto2BGsHb92s44MimWJRua423ogsgFpLvTmh4AqcdVKc8wUUHyVrfCx
uZY/EIUF2v5CdUJyVhrjutvId0blwaR0sAXX4Fh/B5QYocOfP7fTu5zLCxJ6FSgj
k/kJsTOrH59UHORPLE8DXTawUFffDu4j9i0QFsfSIJ2/ZRX5WTFjjsA+wTMoGwns
kUhdPp6gq8wOb8Rian47QRyBrRYV0HtEf76vq3fVgsAMK7NPCiYMMaoZ4J6G3Xeu
u5TlS8R45Xe48q/qydttSqy+x/NnxsKExeFsaO9caE2pCSEgeFO0eBkPnE3/LnVs
LmUu8ThBLnlc5DsQuTaHwp6o4XsXMaxThy3uzxj4w8XMxIXStYjCApO75jRDhUHl
p731geGOG0oJa56O0nwP5w/YuiOMHSV4Ceax7Zjk4MBGyaQ44ighddum8T4wREPS
pNY5enX2N7poA6ZYWFKltLrANXt7wJP4JALQAuV1ipWnU8c2NxLDA8HXlGmLt1cT
EI3q79HdAt+odeIBC4YHD43wThx5GQ/yzERh8geahebTs98jJYUjeaLvzbHoS1eo
L0HaTX1lrRYU8V3Pw7hzDfL4nXSraAZLghhjr7/UgdxgDgAPKEkQiqQQkEauST0j
8bxv0iVstid5Rl6wO6f+3GfFK31kkeR3u8id6VokU76/5rxEe5QB/QRjmjvCHQfJ
Ws4/fw+kpITk/I9xD4z/CRGVDisRALjAd61+fr+jC7GHrY8f1+zj5JVSItJ7n83Z
JQPpiLKTyxhK52tRGxcQFVd3D6i2Q/68cvcAVwntjvloKDNY/IDd6VGWsFkJ/9Vz
0pNRcGImXym8kctm5YaeCEFqmWE0ZiPO10g0qX1OJP9NjV//rgOhenYoB9i4Ip0I
gTIlHDUXNNs6Iz18qVtAM7lbTVaibrPEv39Uqei7kof3dZPfi0FMYLyNUakTYMQi
Ka2NASZVe+8wqdHPZ42XR+Nq3HNsd7C+0IhzMzolNC1ldpg1ePPSoPTlLeV0qpwA
kxeGWbBFHw/H0yamRCeuH5OE9Zn0Eg8QdAe2Hj0PlG8gvu2bA7S+BA/dV8tqjjJQ
tiV7GNw1C0CAwVm3zp4n5bomg4y0cMULBK/XpeebfWKEp6isMfLIyT8jPBXkaNQy
rToA4QHIoUSJq1YgcnRe1DpL/nltLS9P3YJLLOfMvFSIi/3A2tprDPVm+YdHhBOg
v/DKyWmLICN3911zparmUhxAy+Sd/K2lyPWH5sbsoDsj3Q0Jn0DRo5fJkzSc5dvA
9KjYqSwForljC9kd1ZCgCQC1gKXQ3is+KvbsS3RFt5c1L+1brdCUWwIjgxnaMF4t
y8weCbnlF5OLCmznYThxw8qotaFa4cqzJW2rQjOLUrvPz0F1iw2aLBwV8Y0gxJNT
ccF5ZSu4ryHr5uwhmjPplDMGiL/M4qchJqwrkVqadNsnnM37pAZK73JkdtoUI3vO
u7bCfoRO6jryyHFyhxTI7ZAxlEWDi6efmZjyioOBZXGAFGyWMCR/Y/DqYnCFGjrJ
29b0bRU6z+hdaqe4DPTL1bfhob8HqHr1M+MChNEe81PA7G2UROXtcvCQTdgQLIwY
JgZxbfAa9xic0/oCgHqSGUd7C2OE6VzsSEwwUb8MggpyDbwWKP9RtbTw0WLMJlKb
rZOKmZd641JQZ6vPNMS7WbFI2VLs7aHWicfENQfj5q4kvdCQg5aFT3w2IC7AH5y+
ka5q47NJONWYg+Mj/bdbZ61cOH6yPOawTGj3gAhdgnf7ypidV+7DszQNC0xUjIcF
3bRTXfOVy96lITPCEZ2Q6wKxCVP3A3xZZVIXhSY3Zl8//s8Ms2H9+8zWZvblhRJR
ZqFd1FDCRCIG8HHutAy79SWFNG7ZeVWM4Fk7txdBM/HlHsDt+6RChtrrGPPArko2
hvylvStJIlmP6JQ/BgUPrPdgfS7f9VkbZZFa664xL4Awlh036Zntpax2fVgiVM0r
N7bnjK1CNZ5tDbTB5055eCZCi2tSgrqtVcnwKkbJDHb+ZKCb1X6ojLAz8zA2AH6b
+GdPqg8BJARo+3ZNA9LVjYYTkd+Eh8nYmcfIuBAY9cIR0I4QchMAYRsCz3a0wUa8
ItKogPq9SJqcGlom7BkexbeV3YS0fzcCesmw1ZLUKTKePuoxX7nL4aXv6L+amAgc
RVsaUUMRNoTwLWg5MThFdGgtbMTUWpa5eFrbNdAXzKwvdKfFbkARQbImrsbAKSLt
p1jmCrI/tR50zENzcH/bUKcqRtB8G3om/+pcWKDgiVXQ+kuPlgvyjOh6l64EqGKe
foHjOgrgQ/rvGKqCHqfZcDs/XpIoGmxV6HVG8Yh+cwHwH4imiNc3MGCTpJ2hTXcq
+UUADrTNdCmQNcy8eataAi8/HgKhm5CadyfPq06YqdQQH7Vk7/faWY/NpAG4W4sw
JAv7qc6CHeuX77pEyx8XgCdv08mBrU9R1QOtDCBaojnM4js7sVGa+Z1uA/LsxYdA
FLtSWMGH2yJcP24W2RJXazcHRHOvGxez4K/yhGy2YtFAbAFvU6JKgVuoG9VtsScN
+YAOd+LlEB2AuRFs5/EOtdHmOVU4rZ4STftagareWmEIp8LcblVKS1mEMPzsnfz5
18j7+HNU2sGyHKM/u0gKwkcFY2zx9KTOX4RarQgxPqX2GezMRfkL528j+Dz/eUrd
+1KxPWlA0mDms4EZffD1uEBRYhc6nXbF80vM+72DHoUxECLfMwZTPGFioUuPY4Yc
zk1UOXTER3IEOuTbf0lrJDKj/pNyWGX3PAzCe8zEaO3jLZpZeebXcA37iuFPc3Ds
KrsZXzQL0CjJGnw/HbVIzCCZQE8BDu/p/8LWCetu2/XmnvPpGbplkduXWcIGQYZe
n/H5FxI1Nux0blHIfvLJc3myXvnuoONfR5Kwh0+CHdPhe0m43gwKElSGNSQ3YrqI
T4hsrD04ewn0VlPelhfc5RVcDTfF9usSFDJsQqCHvp7Q+H7j1B2bmhKJWe0B8bIJ
av9YBQhSCDYegZy8l7WqGIaGEHVKySBbCMMDbEpaGWlJPxJxY8yfn1KLNkWc/fVn
Sim5H5tC2dAtbCCwiXmSw0JrU3PeaMzCY9gpDo8d7FxvukdHnCSFOE950minUACe
jEhd+Eu/mP3g3d8nEbHP9xPkaWrPATWbWGXq23QjqVm6xQeK83PWwA3V2pfDRAM1
CrDHfu2dos4arh1OXhMAz7zvJUiauARbA3wMzrljK0InM+iFSUJ7olt9Qk6yHd9u
dnDDtnlxPGgxyu7z7D9aGcfgpGhj7ivG9HzKZ1A3UtXdpDnAlWG3A6L3MXSExAup
eeKuKXUFDOiESMD3eddOSfUMpgb09empHBd/jFJcYRg4hjHZyGaQk2ghW5vByzeb
X6zkHCpqRTqAh1UhabNwdA0KJGTFTH34Ei9hTEOqSUnFRKvhPl1MGlQh7HHCkPJt
M9xFuzz2retx6ytitierNiGbqwbsPJOJkCy/j8M3R1+sh0xmPwTJ8+dl499rZU+N
M+/2sgkD2h6tYpAJF0ZU8S2u4vlaltWN+M7NxPJjzrBJERydySogtKzzmdfprw6r
2CKdAhzeBPMvrREFG2aExRW8sTTJmEPBJEwMji6Q6aDG0KblbNocmDddUvGPKnAM
5dmgh4r6QUdX6YyABjOSVUuwV5hZvUHyoonS57V+1IsZfc9+U9KH9hlg+IPHEupy
ao3F+X9hkjCavPv/HnNCfMZk2Zu+gWiqJc0HKNpl/QKSnVq59ZMYhIzRiHyURbdC
kS/+z/G76xcKF6RfiZnIF+lDG39/AYblbVmNCQ70IBEbU8ZQPt0DHlLbXsVrHLUX
Q7hD8Tn9UoIZ8vePhm6guCUDV9nZWuT0kOu6uMRvQ4rT0jDicohDzUGMnhf9FXbr
WZWDFsf9xU+D9JY/dsE6L/MrzTYUE3J/vycdR89IzgJpZwqDH1GyhTRxMs1Lqtnu
8FTDogSKpFnzxLLTaG6QqhNifCg4v+5PQVJ4LBAlhginLQfhnJyQlzH2f9Y08EyK
4QcXlqWuAIG5zv6VlILzvWDRCLC1FYrM3WcZq79zqOgXRB8MzgisdbgfC1CVzuU9
6rvDf2/1yUX+LX7Efoqfl140NSnKVX+WCdpXWxRx44JIfRZN+gXT4vw0jGjsZhWV
esiiwNbJUrzQU5SRLvoBQuY8uDni6VHnqNRyDvJ00NdS140YOYXBBtt5g2MoYS7E
H08pCqB+v30FovSt7ZUaphZCK001YTHa0A9PQv/i0yke9YdPA++DgQUGBvnKjU/A
hT1V3qpoIksJtDGVO4Pr8vKNc2Sq347dAlnlXOnhHSrC+YNMDeqZm8i95i3hnwe9
SnkM9OoErAztsFKehdabaRCcfynUxRQ43/5fgzDFc10lw2k/xgbWvau3l+Z985Gz
J6YHkVxdI+v4nf76dKnf5d7PSkXCIMmjeFLlamjASkAZ5ARSMBh4e/9EOIb+JBNE
6Rkhv30Oasod1J7ZYwi2ppQYbNEsYNSzyJI5gUhIfWOVO0gSodQHuxdajemsoEci
KCzpVeDw4yARDm6VU9A8RzgGtUzyhgWh9dRhuBZzFzKxYVzRuBzxGYM5Y8wT34Aa
RNJGrinhrOtMy4iFNbpO9MYHyf9p+CUQYZoy2CxAi82YYRtyq17Ll0iXR/kPt500
24CYDRF7xt+QkjT2GNWcDkQM9crYWNfczuOjPD5WtdjobMiuxTZzX2SPWtkEOjyZ
ujIXTfXMgGvvqmiSp5M9p8Cl/IsWtxxNj8kQxqzDXVWNIEuiGnzcUTGWIXeKEUJd
sbbesJCpqFuvAu0CtBJ2FBpkKT8rhNx2AH4VtEUEdR3o/vrG6O7LvdBfSAU73VsF
1PLyf2uxbtirqnBcgta4su2MKrRPpslN/8dIef6gR8UlJTiQczCHxfviuHAiS9Dm
tmy4ao5En0iSJiHDsivOUa5jPFDWi6I+s/8OiczaVCd3PQHiyyUjx/c0m+8wEBJt
wsUh8nHl29fTqU3qFo/gQq7cISdqlzgC19fMUIMJQ2tZvsJ6nTsaRsHv0VNlGIWH
GBwDjBssoKxlJZbCFpP2bgm2BXkEB2XP9DOg/3PqivLXBbrYmVqBaSFjtj9VM8DQ
NpUZc9ErlwXPJbLv20XOej5J9Ko58WjNj1EEsaVoZb4mC00fmpJEwoBvR05eoAu/
U8cFCpu2DhOgOdXFdT+TGszCghr1kdYmTL4iBW6lRiQrweqJZFjOUOIV/Nq6iBpr
w1ZlVFUQ3AlWteLr1wxIB4OO3XXkkpnl/PgJC7ux0ilHCvJh8AFSl0HIu56wfLF9
y5/WpOFW2bKqL0Ml7Rti5cQhU/GzipBoxuPreUIw9bf5bvCLAK+qfiB0C/0n2frp
kPl0BMby36ZtRUGbJIiolMLMe8ETpc7QDU/1hsodyG/pS5P2AvtY29AGebTeAqHW
kaIRkLuormgYILn1900pABKiGUOjwNGCj8K87O3Xd7AkTpVZTSbcfxj5GO50wf4b
trO1ktCw4Ar53WEWob1DKcklk/lgV/2hK5YTCQFnyFH3Vl86un2NPsutTgHK4tay
4hHS/yiKcLAnio5ND1jUZjFdMXsGQY1l3Wld7O0bIA7fnW0S02mQXKw2k0r3OqZD
2u8wLjyBC0TYXZCqnmmV0RrOYkRAlLy9GHssz2v65a7kFuNtNcHvNBj13aV++YuP
jo0RS+8qgpHm88dvIjSS0MJJ0PMqLQ7XfPFPxQ+cgOauaQT7CQE9yrdqAPqWySpR
ulSOM41ZgDU37vLzZIBTMxSMjpftylCtnxPTkbmXkZqXb2Ju8Z9I1xDF7h/FoiUp
A9K9XzQT3ORnVLAeV0r8Exa3EvXDipjvKjv8+63fyn22oErY4Peu4fYK50ef4T/1
I/hBJEmUvgbZNda9IEEhZ8J07Sh+YowyCmdNm4nyHBfhDluf+1hygjdfx+hY+Oqo
fhmeRLQjcOynf4F3pdiSqQRtk+2KbX+aX0fOtLZdo2XvhKrOtxDEbUMdbgzQlgvo
4tM5SFK7iOBn4FOeYJo7pF2I2HGlFMc7VPNZ5YsMpKn3W6ASJZQkb1+D2HFR78FQ
d2a/74k5UVK9R4xHL3Srb8lbFmrPIzYs1Bt7vZLT57miwEoGbvHpqo6RMUWZJTTm
sDASWGInyEwBn4mIFoNtd/Pctv//OHBEseJW17+pr5K5+s+x5Qtp1sqFJ1nmxsSb
tduWvfTpqY2OWLDjnJrX1v4Kx4JdCgDDSUVq55FUcrQConSqFtlfp5adntFy+eL7
CyohPfxOXtE8MWsEhE45RFquE9CXe0YKUZHgIpweInVuV0fUrkF4QRDjF9GJcGD0
HPekbze1V6iJJIHLoM3YA8IMVbdVvvWT1V6O/vG+cbfY5+ZqgHJ7gGQSeXbmu0JQ
ezbNjjXSBmfp8PViuOMt00pGa9o6nYWDYeQ7fGEPO0H27NGoYmZtkWlH6gPsdief
5KHG5sphGhg8sPrtDNEyILtvtvZ/FmF76j+6YyR9sLXGQFAj2vfCrWNv0eEs6hBn
WxIInhcWLi1bdaIJr2D2u228rPdajwxIaFswyHHINXOIAMlJl/QEaIVTE+w8ACcA
5r/HTwNf/MAe/xh9w+W0PkTBTT9onRw77B0NFbpJre3/O7h+KnGCMp93cehEc7ZE
Ff8Lacq1FcUvMvVjAB7NkX4IfVgerNR3MRpgUqtN+GEo+8M/gJO0Muo99006Rnrv
vgDx/mpEVDujuZtHRzbCq6qsJtTZ2V6jFN2O13LzJz+5Bf+GOlgvA/5tO0jOlRRh
aq22fcSvUwvEBloHC2W0kHc18+zPgYjlStE8IIGSgMkrPlF9ri+qdAO6wz4iw2yQ
lfVEu4k0gkJrpqIEKrxVBeShYHjQBQ9Yk9XZUOYH+EqVTCrKstk4biH4ktKa+GJt
b1TLkZwFnmsduEKn8BB00VmwXpwmCaIxF8gNeoMqGge5eaC8kBlzEPOfYKk6Q2l7
eFntxFsY1Wa7z4JdzJWR8iqcrZ9hCETOvqLyVSawt2TbExKB0/BeRuhMK7+B8rrn
xZMX0600hIJ5bznGKfFKOqQxq/6JBO4q07gNtyYBKbp8d+jL/gVM6fKpy+ntnJMr
D705/UnhbTfy9gVNQtymP283kbKGuiyzwLB4WDRZ+lAfmotW0R3Tr8XSajH/kiwV
Z9J4/uWouJD8qKi32rrNF2Qax5hZblj5ssDNO0v15BeEoNHl7L71O4l7pLOYhsc2
zzkJcW/eWddMUSBMRMkKXE+a8GdycDVwQoKFnqybhHiJ5yEqcKcU71YQXsBI6e4p
crwvA3vCBoB/fR62ZIyDpy4SYpdRnikUKRkpMkq3f9ccOi9/kHteXoWhMZZEOjCX
aoE+618hWQRqp2JUcrM83pfBKmPMUp9eSTlOOHLAU5+y8rr0edsPsJEWWtsek/i1
TYdrkqNmjvhzl6EmsmO3yNNmb27i6IN8CIcOZZ2TBXVxzbx5rSS17xjpdadk0UDt
uXSiU6Q/cYQu1zjdzfh1OTt6GDJtKUm8C8RxjNRsQdowp+fajxm+0VK5M44ZLK66
NTh9cvqzQ2I+SdzfPJckVdmvEGX5MachuTm6xNe+s24gnfGH92oBLeSCLOJsOQoe
DwE5zdFm6Ked78VzEFhzfRu8lunNqW/Dwij9i8lloFc/Gfwe6wyYlASyYRZS92S8
mQFpVI3x92vA+nMkpEUXGqhmrlic/k2MCYtyEMjmhtwR+9UGPn5CygvXuWy6mAlC
lr6RDeFCPypDIaByw6lyJeBXYsGtrSnYsho/J7HqDmFeqnUBoS5K3KMXTd+2lOw6
BI47bReC4ClLe9uELhj/TtbECseXOjXOJ1AJ0Eaj5qP/b0dkBzpUBNUHYVqRrNxl
QD1hDIqjaa6vfwlOlE2R7JZx0SjmoA05HhDXtLNh56FpiDm3r1Fo3Xz+5FG2d8CN
Dh1IOnHey2gqaYCXIF85KX8/2vSsChCZRhp0P3FAp5mMFqYOq+ZSSA2h8RFrU4jI
XL5V0+99Ouxa9TCWSp7e4oXHH2IlbTmHt/Jw+ZxiXvYizBQXC0Tqc7uCmfrMoRSE
mXfUCOZo5vPp/kK2Zc3xIrCJEZNMq/6UrQYjwQ50syjOusv1I5nEZViUuPtaviJG
p0hIc/bCFs4nKfI9Yqt2O0993VMkzz7kaLdCI0ps8+xJSmh1Ib7HeC0Aa9xkf0GL
6UF+ksZMFGxwJVvMTe/g9582PoGMfpWxcq3pcUfe7wLhJy79ypVdI4+fdwd5kCG7
/Fpu5j7TWCyDpFN7ioOjwm41JDp9nWNG8gqekR+ihHJ+FgaCHTTgcbxhxottha90
b6CbW+ohmTI/9vTIWpurG7AJtQcddh8F0D9AtXSUCwZXmV9rMa3o62cKmFYifyXD
Ehlhg/sHwT9sdWGcRssBRoplee3vciNnvYK5MXjK+RtOeB7vcqkCfQb9CWrorspA
CNqNgjWrMeJUHgQGCDYnn7X8A2MDMRJZbSEvSo04P0z6156m1pOIxjLickSEzJMA
3imebfG+ee7oHlLfkHOVy2cTEGXz38eVFgq2TstEvGKUZy/4MIEo4q2ffiK7jPlz
Pe4O0ZGYui76vTWHkQcgp0JT2zaVQFMy0DmjraEp8bfHgdYDemv4L8njtosqpMwY
oT5htzi1+bY1L6K01RMOZwqDHs6h/Sk7vRfMREjO6JL6RBkgcno4SRrzQyNJs0Yw
xRy4zJF3LnJ5fUGZJFOjCrTm1DbrS7eNKdh1cS6AS1w8iodiyllybsxmV0KuvYKe
Zh2MaJUxmiQZDY7NgW4n7haKv/qlsdTevlIJ8HnpOw6abMndsX0RCHJWKqdwUPjI
4zrsghPOEIiOww63OUq9uh8s9xYJBDdlLwILIQQDpHzDYDYuPMPElef3JmJg5A9b
nFXpQZM4Ke141SjRrcS1khi+Ll19qfvj2vf18qycZ3FHqXLDaH1l0AxIekBaLqNA
KMXE5+Z0PoJfZvHQbCXlVCOO4b9TKBzElNiZGKzapGi86L6/j8Q138tNCCwbeuJY
YpUk52ZuTQABXHE+7M8EIqIIvBPN1z74ZzyjhllrARYJRDvBjyMeKrG1l6chkT2X
0vxE6sHBw+ycUCONMcJog0oRJa4vuT0opfTQs82LEc3lk6FsFRNKTeJDxN2CgK2p
AUnPwbDuzUGgW1UtvIOFYLdles4u8xwsA2pZJbIe80n8ZQvujTmCp/fjB3PUvDPl
3BBELKT7kTmSVI+ztyyPN+sT6S37a6D1ayWdYs/f9q/zYS7KqY7sHbHOE+3rmhBB
sNojRxMt0soh3Y2EZmDWPL1WYwQg7baQMrGi3S+OGB7/tfC828TmCgoEV0dUopLH
IWQk2M+IUuJlfc37tu/J84p783y8fF9BUurZAaZa09cDd9BAabReR6t+yW/xGJsB
mEZVc5TgsINxaFIMq7CcBx3pZkD7xZt6HHrYLYp/Xp6jpJhHj5OtRxL5raTnSVOI
cNcGsbCAnZiQ73q64myEkFEryTdn/NGplrc6aE3gtNkBFaNg9pfShmlAuT0GYWS/
7OPJuLam37bCmBu/RLXzcnffHL0Ftwo5v21C/tDsGhYRfbfDdnDwnb5UHFnBnGfG
28K4nrHc/yOqpGOkR2V/smP+z0IkD8lDw4G/Z8j1vubANn1SyNoOXx8PIM22PP6Z
8C9aOpGnpos9ZiOIRy2p9kGFTnrkce6uU7X2/oZn6QFSsGkOViLkqmyiEd5yLZKb
wZ6Nf/xO5PsMdsA6Q6kHXTBZqGxPygqcm7XD2A7jXTdowrO1BVUNN51YNauYgLfi
QaOtLOvTqmnQEbVjRIGCPdEStckjRgxVJr5/iWuWrRdlaT63cLXvXKDqXZ5Pr0BK
1XbdgH5sPzpyao5TYK1HsXKwzGM1pwoFIteiaZL0sKu5eYooPVI3ISw4ZUzWWCy7
n8Mg8L83KNwGonjiv2bzJ47xLpvQRD9oZrtOpc+tW9e0xnNsBsvBHYlMDDnTRZxY
Ipp4iUIQtoox/ACRMnNC7H/BPWVWwAjkKTY4DKDRN88Hx5hhTGWwiba+pyYCFqf7
Q0bjQtBxslFZqvNUG99NOSIt0JPd1qFpEF4q9jmFVp3utX7s6Id7UU/XSGSujR4y
FAyhXB1RcY9uskGzdvBUTCCnpsTPSb16vibAsNAgZxjMWt1UWWuctDQw9UaytRkb
Hs43hbXdJRDawU3uk6mxMEvcy8in7srz0RwY0RS7PYGh//opC4vpOfMDdR8nit1R
2nQw1DEVJWa2LjleAvdGMjUwrzH+GQ5DdSLbdXmWN6z4No7p4KT6xGKCbyS5et6q
oawp0F11lpLy2uHA4c/lq+lptXof91XZirj8DITaY/UqidurKuSAMHTOsLi0rKN8
gJ6nD6L/3+pdLfF6JkXQ+vHNaBgrq8lTxq1Y7hFfXp8ZUCEO2QBXrQN1jeKnWkqr
INCuFGgVQC3RAqaCa2Vrz4BquJSka8etXgK/2LGuwxbFZr/FVcPnWxddz4ImNq7A
q1GEjLfamBvH5Ejwr8ZV3YR8+uMKy5pLXRXrOcTQk53AHGnJZygc6DI26geWdJWs
apUm1GD8DfyDWofMtS4vKVuZpiNTpyZTacU7o0bfo5gliEDvLEuY/l8Xt6hsVLQP
xPrGvt+qQc9QebE6lvPAfwm5zCBSyNxA2va4yTT1wOkmO4b+gdqhDiJbBe8bzPzc
yyzW9srVaZhIJsx1zkYN0224L6fgmKIGAQ5GFc3x9jlL3AyXytN7KkmyX/EKk24J
8AyLen/Av+MXgTAQsYb8mfzVqEYHaSIo42QJcxwzyVLeLwylL2GEgrWjmGuPh5qp
m88j2Iemtf2X5VbvvBjyYiPbUHDDAg0wazGnCt7ODIRCQvtIHLDedfj/gQj0ELg7
La1sLTypj/d1POWbwcdvRILeQv+K+k4exq520pxLNO7Rc9WHBHGwc7jKoE+EEF47
HVDAoo8vMexXtgrAGl28xBEsXqt6rPwk2cgVTBs9rG9RdO2SPRTJ9CZzjpyo3hYK
tbPuG/3xQ3CVy6+ssOkFaI5iDkkkafp7BbQo1NF5k4rMrKV1/HbavBRH808NLn4A
tIZE76HsuN+oQ/kNoBfrYLHGz/QFC7qVM5i3+IwFDHXmI4t69xmn9hXbMunMRV7M
UMo/G7GRAzjOhkldtrjVWhxHyoed5sndc+JrJcOBeFszGdVqjgQHpj7vnsvk2H+p
2v3EPpOYCouVX7ZdtbdDjxdu5Muu4JnwD9DujYyP77P/JqAjB/bNbG9RVJuMsoGS
hMSPxYdR1q9d1rCQxTer/KSEyrPU3x8/S99Uk1jLkvFNofP+dsHLyY/vzX9O7Zyg
FuadsfN/AXOYRiDAfKpopt9VS/DJnUq7XZxj67cpLSflFwuNXVjkPcb2rkwCtCf3
r6qz+rxcmpfU4h5CRgiAIcVnloyEz4qDtSIeumZYdJEQph9XCf4H7mTKy7r7xYsz
AnerDGgAOuD/76xAFHWkpz5a7uEU+l+Kc/2B6gvw2pkoaCvZAlhSAYCGtZYj2uWt
AhBmyVjpDK6z9CasNC5QiNVyGxmpO+twjH2KTFSQXOQZp7TMOYRZag+0c6l8AheH
BqNHatoeQW1/Pgt1l85ZTbRa74DppgE7KG/4FPO78vcMXRd2Er5h/ur0DuCe9QIS
fi00wev2EZSMMi5iypQZpuEWSebSwdT+nXdcgQpELZ0F7fLXg0DoQM/Ed78kiScN
qITn9AF/Fp4NoI/owLrCKUl4KaWUDBNL7ps4i/0UI/XHYq3h3YUXK/5zwYivl3eh
jY1cn5lH/cUL7cDh7CBfvitFAShu5EnAl/Qkotzp/LXR6qr66ZThNtLe2icIEu8P
CHSx6LjTmVr6zuiaFgCw1FhwwQqmgjglToDvW5wLT95iC/e9/ds3Zrh1Mzzoi3vS
o58MmEy3tIAFj1IjqQpu0EiasQF6FEmnl2/eAqp1F69577+8BQnjA2ZadO+Azv7F
qlvAHfOAwz6AMxhPqKWHmmW2/SsTWXV/q5jP43mXZHJxALacsPFR1k1SvkGl5VoK
y32POLBwUkAjls3Ys7rZ+e503XX2RjDPCzO4Rg326AoRVFilZM9opKToF8MyfCcL
fzGDCohm/7jV0ZGaAnSs99nXbb8ngdw1wZp2YjyhAKgPM+3G04T+rfckpH4nT1un
1TKckwC3Vbr/QlILqaYR3zB8fsueYi92lTejCQGwatY3krcwB8tii3eKplWmM4pX
cqry46poT0YIYemjNLhW//3T0Wxu0VlRaLM4OY2angpytRgZmlOkWwIG3q+VMbTI
2sIUa5h+nhwuRvCJ1HNCXQUWOgWXwYK94jwx3/E4WOXpvZwk/E5oefETKhev2oXF
/RdEGA2QOUoVyyUfd3+3YopVFbpePgDAvjM9xxD3IPDeTAq+HyPc+qgqBLJszcFE
XmpgwuVdTi692NCbmG7Bi2mhInsylTbw1v+vztlUwlC68+6qPP6tvio6Jb/e6Kks
tx0UKBlycn2sGDl5v1ecqPYFDmzBje3nGmHsvwnKAEVc4DTFgtLuD3rXSl3000+9
hPDlDE7pzA1fbG09jou4VWE1Iavu7q6hoQBaHsAG25iw6zUPZz+LzjvhUBBlj1fB
XbXDnZ2c5uuTF8Gn0h0TiyZSUL2ZR0x0JHKIpujEy2NWqmnGU3rcnKaHSwKyOYcx
HMZT3D2ye0stAleuL1Lfyx2FjmsnlU5eN+YvsJGKylZD7ev8F7d4KMEMmxmCqSWx
C52TnFJ1D5rtnW+QsX9uRLpn4+CdNcyOwNveLNFVEBq9hFM9rkLc8B9aZ0VrRKz0
cyPwKOv56YM3wTDY6mr4qdu0g24YvhEKucyQ8CYLmHVlurit5SIHcENODVPSYycA
oqpn9Eb1mtLGvp50pmv9FnbU3iUuo4d6H3dLOEUuW6cIGseljBJRy/tco52gs9ap
4WRV2jZY/bvhHfc0Cv7Yqe94WudKopb8G96OHrU+bi+DQ2xxdK7LZo7ifejNKD1I
vUQXDtoW5MOzEWisrMQzBazX4UcoNuxFBVZvGzUYmZazLN/LLOepHmLVF3xSwvfk
dIKlTciJcMNO/x/4zXNDBwehSFzaRgRskIeGlmM5JKYB/+Lep0hwfJXdRhazJU3O
1qYwLfwfxc5kGYdKOL8OqPfN9Pa9qLebGcU3YDrKyhlfIw7Nx5mdshGgmWZncqao
cn1t4Dn9uxT9WWOz6k52rr6oXb3vGsDzYegaR4sfcOdlLwmaA4wHwkUiSmRQo0Dt
If18krQ+sG9mXS0aqQ2ygEfnlv7+CUb3OT8na3/VhnrfJ0y4GT5YW/nQvK0Ykz2L
VGG8ww4zgkrbhBiHFJx7ZOHMqEmkkGSSJqCYR865xsleLqW0+dDZ1RSWt6WsQ5AM
oFu2aFBdjz1901o5mlF9dkxZxABwY0La0g0xricD59tL3gfNKF+dyX+ErFW5FgY3
ZQ5Lw2SP/nAv+ozT9/rz5MPk9lWeR66kwBvUJoKQ6o0yDLFq//o3bdb7YBXKWs87
YSYtm1cJ4TemOtufN24hTVvHU4/zXG6LLsYSqQ1k3ynKjtW9Dfi1rkdtcXERIS14
PrXf5eutFsvnyE8yB0XTSPriQzsEFYODKVgnes9KJmGDLRqo3ukGcw5vVh+CTiyh
sj0Os2R1gVqyPOFNGG40Ztzp1XVi0S3d/2ZPiOCw40C/PLRLGZoQTbFvYMPNsrzx
lxlR+WXA5u/uO14O4WdQUx7Sk/+p846m+khyeJgZ3oSwRdsE6zlEyb13GJkmK2b0
s5SELcI8R7KTZejSYbaTUo/EC/5mk/sx5s0vIil8UTN6kT45NMYzKqY2jzjXrByl
CYjL4dGx4dvn1NLRpmmsvlQlOgG/O3csbUq5MgWBZo0AYrjOjdytMOftI80bDhbb
WL8ROM8Zwqxej/S7RLLumgmU3qhwy5s1GwiMuZYQ0Ysw/ATXqPBR7kLi1WBrCHjs
5WX/hGMTv74XAs5Or2fSW3A+e7tukDuv3EQFszmJUaKi3d4oqm55nOJPBQeZOAla
5nk1LZcbhNdRyfHV7rNIdr35CJqYwagceBRmIw1fsVfasTBSlMzCLrmd1qUPYzcZ
OL2QHuI2PsrujjT3Ea7rXov2aZ/76JzLDdU/gKP2b3QM2zFe47nxs410KiiUh3dL
bqTxecMUy5G/jNLlsvJHZUB/ELtDWP0uJhDK7jnMD9xth11XYRyn+QaOcp2C8Cap
x1CME+7in/CMbETLvVVAOta1/DokDOkCl1VeMFmtLxdgKjiyksHNhySY8iDtGZjB
8LIaB0Gg97TzaUi7QC5BEQsZG2tJWirOApKSXLQQ2SVy2E8l7IifVGR0Fc+iNggr
aZwywCYL5od6gT9HArQ6KlSyiWwi6RJ2uy5GxCfJPwNbsOwwjwVXQqTsQldTwj5N
TRN+cyW3eq1XsW5yrGR3Avzr21NohkgORAZKVtZUa2kWx7G2gWXUIc5tNHFZ45oc
A5tfU2adV4RKJjVxAI17vvFHkTZb2H0X83O0WZlZqyvHyFlUq1t8xh6myzKw59Ew
QErq6TH/weS7Gy/y4Mo0p0CLP/Dn02Lac6MpDxMDzE91A59pzWUY4mr9p828s3Ah
Bspm4riwjNmywaywU4tdUCeM6hgqrJAQHEQMA1yAr5OG0SNxiZdTQO6ui4SBT6Qn
YmBMBoX/6hD7lH/azuIXZgKeeeyakWxixWO/Q08xF1X+pM0Dl0atL3yc1Lla1/GH
jo7ZbGurskrHGZN5Qev9J0JKBYq2W72/jJvzgMrRkPLcLMkm7bjXIYeSmbDWf7cg
MD0PxzGqP02yqQoiU2RDZeAypdBQ4o/RfQsM0+oGfgNYQoXAM/G1Uu4iE8KShqNh
6KegCz9G8+ZprVnpbrBsKgilOSGGemw4m54/7b/iBPLgW0Sl556uiJCS29wUlEQQ
/U2HpsQlw2Qpr+d70hQ2nE+wb6i2zwMaNPqWfS0PMz50EILxrv2uFaUOhH6Tkp17
0cNhC62sm+OgaJDlIY2ijsAp6FEGLNl+FxNdnxREECsL/P/2qnfCui41Xrfy+hxj
8qSjYCKkbdfcSuLKPF+nlFTTV2/6DLzLhbWrfrJ9bAQadVJm0Bur0XGMd9X0PhTi
4vu4DDyLcLKvj7TfzcLguiGeQL6VkcZ4327qVRpXCLR4pK9cNQifrKeM1W5m2quH
aLQt9RmdYRATehFgl4j4MYY0ycs6DwZVxbKTgUcPpZ82+joxUJv0IIECRd+A42fm
NSEuon747uNLs4vDiXpNjB7m9+3sXwI3THVZCcwbQEuch8HGvqWszTb8diwAnWGR
F8QvBhKZm8wdUlkL/fklbhcO/d2GbgIjBylOwAdQR73fGYjPCXT86Vboi62YPGNc
V/ImTAL+yuEDrvikRQeFRjoT1FWCebzK3ijTy/bC3e/HeQ9+VYQ0/AfJY1tD+MWR
giFRE0GaUJFwd7PnRpvmi3ShQRHiNDAaHZsxt30aQ+eTypFyx6WgHlLyT0n1NtbR
lS4605hZ9O30Bd/9uxb1S4UMj/jkmH4tcsBxhEzW1SG3TVmLZ8BusufuLQEhSNoe
nDww7hqb5xsE5MEQ6EyFSOLVXCJKCVhD3x6d8h7RKexlMQPbDksNEzNaNmD2ashZ
yPZ2Z4f1hyJyfzBXfm2w3QVfv3/GMI8Kl9xP1ll5HSVCMuqJ/1lqIx0PXwSRQpFg
vhLwie4sbX2f8uZ6JeGYN+l6mL2djWuzdeSctVTRf2KLJY7J6JENtAQgohVlQToo
WHFrzbxZ8DAkZT+3OevmKR7yGGi++Rk4YhkMgBvQxjRKajxUHJ8HbTGLJhvOMBhY
IfVlUHLKLN4kpLav5ubr1dBe9dNT+BfI7z0E7jKQYvrebf1vs+EwzMUt0NscTv0L
jg2TfMomwJFfixgWfbxg/3NmmdLVi7cByA4e8ch7X8YKk4E8zz7rMb0LBE40KtFu
qVOhrP44F4xYOEzGZxmGTxg5tyBdwm/pbDCrZKfcyTlgfAWx0hK/y18Lkd1nK7gL
x5rOLvCa7l3ilxZF2+TWQ/sb0I4Hxg2nQhTUeE/Ia1OypGmND84KHACnn8mBSGyC
EyqEJd9Z5W4rY0huZe7DZPoQyjzrJpp7r4P6NrMjWr+XfRwTEcG+HxaO3yP1xmaI
4zOUFAfMRYmq7T0LJnl+8gBU1yJTgNp4xLV5Co/zA+/eNF6tyw+QHuJ5355afq0J
kW74W/ktgd/W0dcSA1NJ2s6ka/DZzXRvuq4ALAkfHt0OOxbjmbVJp8JgODP0g72i
vmcQlRNgiEKKTi/I0GoSNniu0mFOgzfkiBfqR0++N4vRSbQzzI4gmTt0ypL8Rp4G
MJsyFcdznupTcYxIE0Ssdj2FIkchXV3QLMtJeKz9rkZtKTUzS8QmaOTHzJxQdHTo
XyCGyfVYXa/kvfN0lD+Oksf6MrssqaTTN1i1oh059Vf5dtzpWN5+mwxemWxBU3Z1
xfQd5hfeRVzUUO/GtXE9Fw3uoCtvGqMNLz+oA6fG/jPVmnWKKK/AUQk1PAQub7cn
xuHyBig/80mcujS0D0ARjf2Nk6DKbl5k93GarAh8zkSqUv4VnxqIPUiXVCUZKC1c
e2ZV2Zs4ybJfcN+d0zLWIhQqrz7oZxa4ksAwDMvehoL48jY3ffNGsbNPObS2LEHo
3RS9U2ChalN4Q/Qt6e3ILS8tr+4rRpTUpuMQ2AmdQDUiXQOqOkzhIIkgkE23brpB
Ng8VMiU3DNsz2MXeYVmaNKVaPZsaRm24qvM7jLXYLE6Cl61kPJeQTKOGtXKuuIlP
ySx55VfjMWgceCgH1PFd1FlyIhUlcsIzvREP7KaDup66tm2G5wFq6/MhtAFbhhmZ
v+xC5gOmMAzbwitCcSsUeAYcPcBDPvR9ebf0LJpy08TO8eveRTRqS3NQ2GxWC4cJ
fbdBt7R/TmlCIImMKZ6Yf8uvV4NeiymY7lZOdxje47rlJihzCymB65Kdb6t2VjTP
ekg9SZ4QDMeVkrk76Jd2WDLwbYUEvHU1XCcFi54D0TvNH4dOd9esP+3pdgQOKBTa
LoUkmC0qd0ky2JKcHvClWLKPL0kD7+VTC5x55SZ8C3zajT4uty+95a+SOw7Q9VGI
HENuG+KR+9N9A7TE/K7gZBWR7csQdrfQ2+glj2rakMuNZBuVeynzmOya+jvGZeeL
ZsFrwTy45l0dvoztsp0T5yIBuFvZNMGQbvbq7vCuRha71KqEsceNvgwma+cqyqIS
bOVpDc7q0zY7bPG10UiaUDR63bKi+qIV9dGxog3mBFQL9bpu42iQTX4lxAiBeWHj
jDvOfkdWhgq2ZSo/WT7o1CThBOK8/k7SZaoexfdNiqZS6MGtr5T4m/JQqWxhV5KU
7sOBxYhQcWsto03PC8zhjDhnhOBvZHVNTRUJZstkJS1CDgBdZyPfBbQZyrkwf2/p
mHU7RUHR1z5UXtg9Y0Pfb6TBe3n9F1F2vA16tUaE++auXCDgSUE7sHUdk6WG991X
gHX2Hqnzr0t190FEOZ5aUCEmXDde46JuV9tB7t02sMm6xKvboKkNqn0jh4ct36gC
UytqiuvPnaMwzBdMFdqk6x87iKG2VZQCiSw0ZAtKMjnVjIFXCLcSiXz6xCFQzTnM
W48Wge+P6K3VvmjcFJRmfBC9/IN5jJz1J9A3ER4imp7fM2PocsibGQxnNdWBUUEP
FYV+EKxThtFDT1vlRWVbxsP5XO0vQjFb2mBFSyuJp1VxM40uNC0lfImMYBARAdVa
DaVCx8sCPz72aSOVyiJRcHgB0YF0dQvweJ2HW/ofjvwU9V0fb8ikYjQnmusYWt81
rqsdRAvcbBWqxK1Cs1U5HLfjOi4HENJGCD1OW6jl4SEJFcWhlMZ/49bYeq6EDYRu
KijxaLWNOJNCFyWxevFJb5hXKY/PUGerWkhn/0UB4aYtfev31vP/yI5AZf2trcTc
zw+SI8CiczgCBnksBzR+AP2EfhIwM4nyWhSsju7tdI1VXsOaTICRITNel+5nsxBm
uHvu0ATkUZZWDBKbHKFNYaZSzztbN7pB8oVsOplDLSRdf1z8xIIkwTvzwlIJCpVe
I3IsG3aDBa2lgoSlWVm7ft+oaHiiU9ok7UPsKNIpqKqaM7TI1PGLpwaWDC9Z/euD
BO7eNxnEq/PzQSQNVzhotzSNvFh1M1l9vXtCo3Cly3JKTLJ1zpU6UERNQ+27Uu76
8jTGAUGUmiw9OmfyBAKGpj2ug3zrKCtZBFn/ayfZIh4nrCr3HRt93oYZMBWRttL+
308QoTlaIfF83mBm1l+vj6JWRWV+vvmKfBJGbuYG0uq9J5EGLwEn/ZpovsNV2Jvp
iKlmCAqrkUhrvPoU5l2D2eDsUENRFqHdShglmcEfHee5XYrjaUGfHpru650DzK9S
IPrj0XNPqevzo2vb9mUsqkGujalnQvqqOtuFZQ+cLXoxd68xkH2WXoW9CDphptvE
iWUmCGSDeiYhQ43N19iTrqlH4F11MzBR200ZA5rqh6KmibJXZZ7N0WnHxpRlCBuz
GNNZBq0OUjAkSWXOf32Y2lLnpw7YjYkTwDXd+u3Ok9wreOKIdE44N1gVmwqVCQ1d
kZQjGWtYo9IA0Hv89bMJNruJvTf51BLD2/ZVN9HGr4+kHMeRd7TarPsjbLVffHZa
dsyjrHqkSs6rqJ/PjVBaEj7b67offGyh0LfTWgwao+aUxSFx8LX0F4E7z5i74BmT
YTzEt4p/AwkwZDJY3hOm3eACBN4LuwmSiSogNXkU0n0H3mI4xe0y9DOJkJd9TLGE
LU4LMcDgwpjKeFCyCAwWrsLmGKMsQrkA79U5ESArluIE0MUjt0ANRyF357jckrgR
3zg6gmLAoQn5yRFT+C/3O8rNHnb0thT2fFhbXr9yf4W/s29vS7h6R9M7apb/b0EV
vXjxcwk9KyeHWyR/eko5mI3PnsUWHuob3c9rYLmz8Nu/+ezGiuadNsH6Olgv+i7y
HWXOfjnd+VDo5wyHiDKBkf3NIcX1vRpQaJksAK61B92vnjJ3SQsdZLfMZKmCNnFw
IAlfn6aR4VreMaYdwH6CPKC5SZ+WwDDUwOhkgz6TYWE4M2afRXR+5WH+8CFs3S+k
s0yqcyyk5CHAhy6ao6Tgpxk+AP7PhnfZaAe44atcZV9AKGknYSQ2nkl/VV/l3pC7
AmSmGzB0zvs7HjU9jhvjJ2GpopNBpFrd90Oxp+KLit9s5UC5KWukh/OfrqVu4ufi
8w49xxBySOVjxRo4pXD+kbiLlRktfqm/1b3MR8PYNsOfxYE/e4IxTfCdvnBd48qL
BoqngR2kDzb0FWPOR4f2jfJ6cwrmICpAx6cGd9Hco68fFdEYZIuu5PmDsUicwOvL
oqSYgeJZvXUaglFzvGkNZ4S04U3+g7nclm9ohX01AmEIOTcZoR7YuNRqfajHkJGf
c1tr/Oie+9ZYl0I8vbsvBrpuWnVsYcHXe/rseROSHmmgoUvxSrYArWEkkE5cj1V+
3zBvk/3H+k0zV28FFXUKipMRhDGZsQOOsb2S0ouChNUiy8rznGRj/Yf/EJk7mw+U
N3mdKYCXJScyP409RSyUcJ1tYTXqy/oOLDm4yrilfL4dfxeoaE+/Ro2uL/j6kqD0
2OKQ75KaHmvFHPvbB2Od/FJkFjGEIBjSsP41BD5B6jVGDnlRKzx91w8ZbJetirtU
ZBQXlc0t0lrN9rrFR8lnEZfFkBH650XnmWZUgpDmImyVZzMrXD53s7UWVmQah4NC
xowPanXFUSTFK3EsYNG5Vm7UnLdLC5dDUUIWblVF3rj0YcBuBcU9U3MxJ5+YslNU
00/hiqy9qLmmDifaml1bMYBVrjnpmWqYA9PjA95Y+VJLmZRqaCNxThc3HVtFs9NU
8saMs3gxf5FK7vbInZQ7FZXpLi4OYEERN/Rcb/7vNJVMER2qYogKk4JnxdrbZPHa
rAPBqw41/MAp/6T/OMPi5NlI/IKvsLTdw41poEFSj+cFaVr4zd2e/VkXU0hzRZts
JP9WS4DOmluCF0H2J8mP8pSHsvOEK/wW2rYdXPNATAccppyRDXYBKE885vTVYncO
kVXnSfAP2ID5AzCt70m5+Uxa8xi9TXVvQDD+hu2yK143SLEK5l1rakE4qs7S6ENR
lDM9nx8/UcZZSsloVf21sRsrmW6P11wfhi618yCT3HH9d/gbqQYG9K8qpGCv2ei/
gRoAIbcFVbmHtRGxK7+9SoXZfxgmNqEj0Y9oMKQuADiq2IKS3h6wq9zwcZ7+9iGR
HXiqZIZ0HvjJEEBKHO/+cs8fOByJynXVLScpRe39m7KlfVqOdUdmZGZxTuLKfHeT
Q44sWs05bDt6d0fPm0tnXiWsacRvvZzCTptkKlBzy1+J4wkTcP84nwKPrtl/eDf1
0rcNqJjo/swQiU6Cq6xbbp4nwnEh9zO1ueJFgvOS87KvJ3Uhs8uUGZSbw9MK7yLf
XSmhyghsNQcl2106lwDIeyfbDD+UMt/r2hHFhK7R+QeLhL8jj12A/sCTLAmNWurl
v8BvZxLywxxF+54G/3ehJuGtQSzQs7dBkxueG1OYbdsFLYNBPtrWWObmgsuNLnMz
cELyP/Fap09RC83oi1XmsEYOIQQK66AZBVdb0zvBopVjBPICY6UvJ+IK9I57emuk
VcZJSIi2/n1tpipEVE/3LCybDK+GGkCjXrd7M1uL8oLJnBqEYlZaTJf6OTD4GmCD
ZCE9jwLQoTM4qnRm3GeiXRHLpsKToFUynCJ7x0s0Z0CJHu1z7isCuEXMaZk5Jpzu
8vAMn996TllPSX1cI7u/E7A6w8yY2myLL+RYxxbDCid/ug00/sDTMkzIbf5i0+vE
7wh96f91y49u8fAPgQ66D5+o20FXeYtNX+AC8iAqhKSZ6zgoklCMWT6Hk8d0f6Gi
Uy4d06IdCFXC8Nk6Jtr6IQDjVzjsGLlxW5UCLBYKQgOdeNal5tBuUwUh2DejY1LI
qS5XhHWkUz1cjCNc6dUziOQv+JwuIs5TIlSeUiR79EJmYZZ0+BZqAPHuK1eaUg6C
yRcsgMv7rhgN5y+RWlcfwlRq+ukVEZW3+bNZ06P9Q1t9EiwdR32ZZQeVWz1F0s6a
p5/QLGsz7cFeWXTO9A90sX/aYfh5JGuR4HEYmENyWlBv/SZ+N/b4id75og+Juruw
SjCQlUnewgcrUL+W5sPhhEAWQBOFPF4uYIATw3CPr0kBV0ZUhFTyNyJWzx9THW/b
PyX5DszuWkvlUSgcTRPljw2W7HUIrAaUN0U5i6IzEtEenBQOJ0T4R7XMGH478Pmd
kRTE2S2KOi8aRVvjhn1HlRo1V40yY4qOGSu+oJLifklrczYZV2BxpSVns+YYDpJP
Q8CyuQq5ip8kx8HexYj32NIQXFC2hgA06pVZeQrKj5qAy9xPsSBkXlpCuhUial6C
KwitmQyPq49l6h1Pn0Gq8NGdGcZu70ck3+3BkMIfvN5qxWPS9elHEnMiWyWwWh+A
Bf+Z/aqjRkXzyokYLF+Mohl6DnnQTXhf7Uk/PY+Kj4K1+GOtt/9xR5L7LUvbKGdh
HToD2l8E/5O2QRDsfSeubL6gogP+ko0W8G8beBRkSJdqefhuyySk+ipHVzjTCTX0
0fbzDZwsS1loCBXDN7LksND5UhqmKez96iVxvfKgBcWQ5GU0S9Ta9Q3z+5NX8C2x
cgJ35H59+abuya4YinvbE1woKLIDPbbUq/9Cp9E0j96nbBVuvhEDFzFlZGSv37AP
+vt9fo/U1B9OPxOVbLdbzp9oPTQCRDUckjGxrYHhQ8DYcN2bwT1HH9cYTJAQcV/M
rC80VWckAOhNKT9plQUgUjsuVDl+nzWi7D7ComivjwyRBAo7sZXAbz3QrVJdi2c7
FXSgyq6NrER8sot/6isofvxo2Mxs6awVbtXn7VQOAFdeAESWGRymrtSaTTzH1XTC
UCyJIjbteYpdedrjOvdQyin2nU/6y2XzJdu9y4/PrILK9j25XCAvK1OB7+wRz0lB
2frUl72UGMg3R7DwylJtZcwwzCUs9gUwp1oI5DmzJdgEIYCpAPvyTy/dFehz1wYu
GTeFzJGE+BCCuUSSXjSpjZ+ZUvCulmBaLXrs5zuc2F3TVikYKv1OZRwctf6SsPZT
F+UOprEiw3Q9gGN0Am1BBpqB5DZumFhTD5oIzB64IiuHZe3XKZcmsIL2Pn1ec1eY
JbJ84A0ZKEfOrxmG0HmEK69U2kZtC91mDo5Ub/2NjoE5dVzp11J5osSjceVIMOiz
XMx3ybVYq7/LKisIP4TYfcC2sujVRXZXrvsIm9aWJ/WkQL7eD1eYHNES0ZcgOvRW
2jnhZvBzBrVbSlrvn8ZreXRmaxzyV+zk8wX9/rulyk+KqBEXLLSj3/ir86wbyPs8
kKBZV1MlihsTIpBfi1H5TbL1MbIQ/ya2gMI2ISRuFCkFmpdZyq1LiV7360cxy95F
oJM8AdNEnp+6scj1ija+/E74hW9CiuanxMw/q8FAJWsb23//MfSlULmUhe+p/tYf
InWflMjAHJ3JVS2T3+/Y/TJQyl6ElXoziJD7rsxOehevz5I79U5CiirRDydy1yOE
aejIWbfWfL9ZkBPOytaip2kKfbmLKQ7IqH4Ua5AP/Oo=
`pragma protect end_protected
