// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
amX9ubJVi8HPXLHN0OVC41LI1zdqF0Kea7+7eC0SKez+jd69u7pdCWWBOuREQENJ
ja6dmaqbb9mU4nMQNUFgLRVF7INi0E7Xw4hkG+euGb9dcrO9kUhVIpQW1oM0NxZO
CARcQuf0j5ATHDy8kCPX05shofmAdg/lJGYWUHBqq90=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21808)
G2MhhDwvFsL9kjzx01GHNy6v4QhMtO7RjhIA5TYmzGXhEHGJ2Fe+lhZl0kvmWZv2
9KknkO6GmqOJSFF6PiJ9qK3U72/QAAqilC5FOmym9RvKNdwoM1OzRiZL2F/uVwR2
35klhmMbI2hitmyWhKdrS+C+1xtuhZH/ufnkZvy/ObqTJQJwA5OwFtCFvTiOXyYX
0kQFFszC/VC+nJG8XbPcUdJEDeJvufE0mzTWw3JRqrcOEilIhNqoLd0D0UMOnLqB
ffSk37k0Hw9DCvj2dBBtJW5P/0q3JKSllX85FcgVMssrAAw7M2CeCADAOsVpEWUe
CucsYECpOIPoc/xgLZDRnkoIdbQfNMIQVcCppVDfQAD6z5aXGSY9dn0I7SOgrCK6
rh/Nbn9e38DD1BDFNqejLpyRcYyPmCOS0n/BbhZmjmjKPfSNmQ/q2hbR0aCvjyrA
B9WF5jYmn6B9eQ/pS56T8uCREdHgBS1Mh3x9pb/jRV/loBRRGy2mFHVzHdoZzn4W
U+pLwMCo2wzxVThuHx4tNlfyVZBqqGkiieJL7AxQcjDpsZJZxhqtpOpIo0YRgbCi
tjXF/DhbXzqYoFG9vcVgfwukFZ+FWioDYQlWi9bxKMxV5ez4H6DQ5Rh+hBTN+2vk
m9YNlAEXQHPJYaRALFSQc3Ngk3FcK+unQL8j7CK6XWvDaTUUY3YOWg51jVdt+tch
pNXYC9XrXdA449IR7mmBpB1ciEtlUCkyiVRrR7cPAdlrDbxKWffp55O2gwX3gsbS
5MJg4UxH78lP4zLUrS/zl9jR2aFpmCKoNvf5MQUGLC0vREp1Ees88EhwSEPNUgJl
HOQRtavAvAOg79TZRIzo1AFaF4+XBC/0pGq721vXCw2V3ANUN33tvGZHPced8Nlt
F9RswC+J2A3UJYjMvFEu7sG4Jxd0uPeG0mfpaKa8Q6CAfHhzQtISbRM3LdeGHeDe
yNF4Jkd7V2DfIezQ4GhSH7n9MHp0ajSTC/bglH4+fYZyO67oxCVfKuRbuuXkfosG
AehI6jT+Hdr+hDrwkc71eX+zMU65shN4mgbUxSUvYPqqEAs6kCA7vJjgL4Jkryjg
EiN3ntgnkuFHq2KrzU0Pn5zmJ7V+JEbJflIM5RtafbCs7EOU1HXAS3Gev+/wH2I3
TN/v8qdtRd562s/xxUM+VfuwqJ7IySk558/luIcmTWBXQBrNoqdI6lHoCMhp9/GI
Fs2gKcUJFMhVJZmBGIoW0Zm5aQdP4KV1+fj1fmHXHhSqB+4JEthrl7t1MlqdHQI4
abzdjGq31XLfM9JrG5ChFarnk8qCxxFJnUoaxcYNd5QAmXekSINNX3TSUNAfh5pl
wbyPdxetJL6Bp3EQu2YAQNRAOB6qpSPG7P/P5UIO6C3n0iQ+mN9Kpk6iPiA6skiE
tfXY2FN8RxOt5ZOvj94ytE/CD/SOOqDbZ55vgNbSa6Q5AwQiCGTa2h+C+25Q4Jw4
FD2HZFq9nT3Tt5x4VpBGtbPBcfSpWjjPBztXJfpssUYLrdSohvqJKO0tsHt7aL10
FWQ33qPPT3mDrjtUqv17ZslBNdEDDOOsjZ7082UmfeE2orRfixjllg1dgSYS0F5r
j4zNWarjkueYlqo1ouZUcREzKcIJWhEn9BI67KTP9y1lonqlAPPloodzwztOJowr
VGpv/LgLusU3dW2kIdGrz+bR2gSxqOHEw+omQkqgJQAEO84L6NfBOQFEPdZxVLQl
SoUtbLl5PJV6JNTgMD3N4hqxW7tFJv4qtecETaRFS8OlVcCsYud1Xpik/s4ehoSo
KUXJH8LQkcUnvykPc/cf5NRV2gSJ+VVmxXrfSaZTTGv4UC3e2Y+BeSdHT7jwkyb5
fyD51LJ+oKjNFFVavDqG58otSW1N9HFPoHKyjgTsIaKhDu15/SvjyxoPSJEw/2F9
b8tleNRjouGOatCEEGTD4uDZ31YW+A9ZtUYDyUtRpNn+L0iP1b3UxQt0RPWmigWN
VT/2cilOrLGx0TtRbM7EvA4g+iXRZw6IH4t1BI1VO0xb+eEkPVccR+mr+owUSPA6
m5b2Wt5jIjfCSMCSIL2qyH+SnLeDI1lmra6THLUFR1CifUi3Z+0B1JhTOUaXibBw
dYDQkHyKPq8wIjH/UEhOekTtfFm47ZzSYHNAfNHlePq6y1wlphtzQ3VMIbgQCZHO
N+pE7wDmqDq2IFVJSiZZZh7xFi0+Z4BMjEoA21EySbQbAZ/rZx2+5IBKrBUGDGTX
pLE/AUd3/258rGE12Crv97ysnzuDcIAfRXgtvmqCUuzQDeD5Qiass88zIIlgv9wV
cL7Rjr5rVSP5FLH6Gih8ay7A2I4gapuwgrgLvV0AxEugnwfK1nC6xBxvQ0FtXzsY
341Q2nMbTC4kIYW+zenkXbtCWMT9KpFSpyctfhWqtb2xbdf2rc7Ki6i0ZUmyHV+P
mohET6wLNtwCHc5tjTJiumabNrlRSisv4AgjdsMJVA+e3tpy2Dl3pQ6m9h2tUoC8
Q+zIglGTY3YU82uNPFa+6IWWeS0XYffxTN1W32rT2Thmh2jOu/W0WzZM6E9iy3z2
MNW/kkOm+Gll97KMvgxCc+/hYLeXaP7/1CLyR3U/QaflBpz2Qyeg+Fs2riwZFSzg
6Jp2wE8XRjqvwZNrxmg/8ZKZUFp1Keii9WNgGErZnOnPhuRCAQxtqsGYPjcC68hW
+x/6fxJ580Aw2pNivgjM5/bozxMVpPjgAsywW4H7fkjJqBwaemTzhET6NEuXA+Vd
2JcFz5+AsmjPZCYU7v8MfzD4YQgyGTRPYB1Ht23KGRg1J4d0IFtDzYTq1leHcjzo
A0HQ6aCfRKtkoOzhKbx3pkINJC3UtsdB/o/F/RE0wrLQpmSnOHkIgWq1slSYOXr8
cO//E0IHnochlp35X5Goo6bN2OZlWr8GuEzPbI78KTlpYUyj4E8dk1M2frfm/Q5V
fLyx/B/bKoEccO+iO8z0E33NOxmzVMMm32iskhGfkvJ6+4rQmGtIVyb4/cRhz8ok
pb13dCCZg8PpUZMIftqHzQrjluOhss/J/4+ovezLiyfNnCmSRD4K4GNVyQBLTCn/
1DplYY0H11XPPc1ssoZ2yVSF1kEUqdWdAhKAS6fQBkDkFBm3PvApAcIC/7618Ply
sapmzuUMb3B75P9ZFMFl5+TmXrr2aC6J+dTCxOrV9qOscNG3qX7zsLyHcxWsuAxf
jLtS8skopUihUMNoQtSWihnjJXR2tqjnldUy/FLPGmsTPZh0c8sQULC7rOAWwkw4
gSD/k3DIkNjC2DpMQIUv9lLpxFeQXYYDkbJv6ZQpLtc83eNgxcQnXOL8aCXFaKfZ
kHpnNSSles3Z3seM/p7zFVgKUlggE9mFyaovcdhdWpwexwmf8JqpfvrhcjYg2NIk
GQwIBNELQ597qn0AsAMk7ECF9I/rw74Khy/JQKeW0IM+jWx+Wjiu+x48JNA3O860
vP6QHqJP2qO5KX3hIE7VYZjYvWGX9gdnJcOvRCQ+BHxly0wju6aE3jvN+IY/eXfN
YTi+slp4HwAX09bTN1uFA2YeigPSFyoXDFkinE4f+6PHc2wkRrnwEm2o0/wJUy3c
36V/AyH5ioKw52EHfWCXY5IN2RDeMqlW5Hj3IM69zHFOHBDyG+bqHZ6Z9prt+kfy
HufYDq4WQ2+JH62XRxVTW2FbhtVdc0atyI2HvvzxjKDM7GoGNwRF/6KE9qY5rvbc
umPJ4XWng/ezuNXucDsEe6Xpe6ISdKLVIvgYKuBb1gFd1CRkFXe9hH931kGFFAr9
oTwZfSmMUxWzN4H3vXVa99bfnOQR7V3dU5X9GwM+hIv+NhQwyRfa3N9mz9py5XEg
XbtP/POpJa5UqEE/ffvTdUzPVCF0ZQ4v26BrZRwmgdZam8NWLPePL4SGAg7ChP0H
L9TxNyFcJFVY9z9cLyFkJmQnmNjhTYHpsyvcPlAY8pxCGUlGHrutFfFOlOxLjiQ5
G7V6eepSQmM3oILjrD70WKwnu/hUAYLR5U40ApniaOMCXQ1i4Bp4ZdfRhlOiIhFx
6/ls5BumCe4x2ZYNLxSfq9l78g46vbTtAGDJGLY3vrp3wcJu32u1a7LsmryDX49Z
tSNIuZy/JpZUPu7FFz9Lqli89S7WtRSA7G8Su+Vev95eqo+XlFdjVZvmeLZ0cuDv
qdgt4gDYT/2YzplE0theluLJH1dFBsYSzEKX4j8pbha32AqbDmIQIWvwFK9fDW9r
w0NgDepDHRuiJam1q/61HsTBj2DfmUkpmFTxsq5qWDQ+aGfWsI/CSapk/JhNV/+4
CeXk08GkMxwFJo9qYkc4PaQG5a1FMddCd+Kou2QXgWUAh8i5DsP01nbKZlRWm2PT
3gnEmpFvYofBOxjKHQkYTrwVfnaJX8SKiDw8cZpIwIrMTWGDLd9VY/adAVZlXCFf
M9rfzTFtzl4ZY6N+OTJn0UttkWBz0E9ROFkmu5QFjHWiN1rUKA88U84SwKuNFkLT
upim7tDFMI6kiBSd3C3eX361aYFcHjs7DhE3frp2IPfnxT/OGa7gv1SlO8WtxIhT
wjKaRaZNO2r+ywIaLD87nfRunEKJoXRttr6z12VWJF4asahfIEhIonxMnyjKbsIA
xvIS3EzrF1xJcWtWAOt32ZS4pvFZtPB0ZXtOgmps6An8lO+Ba+9qKC1Qs0QN+cx+
l5VKYJ3TqdChptwveXp8EUonfraNQI2yVB464x5mEvLHK8ZVAEq/TPREG66L6Q0C
roQrg4XD5p4wPUpL629PDNc6MtZapPdqR6kYYbRBQuJY3C3iva157YZNybC0w1Ih
gndhDtty8NBvv9yKktla+nKA9ONqNapwEDM85dx5lznPN+OdM1gJr+xMLiFbZTc1
XiCs28xVuGd8C1Kc4RZm5ZJGkWDvFn0ZaZa9VQruul06hh0+zMmqB2ef/ofgUydb
ihLIQJ/BreF0jSB/DLPxbZI+5xGhO9amVGw020ALmr3wr/PxaWcvLqxFzNFa+Cgs
/vKxNJU/JCaJQWCCdp1Ui+sYtg5LbbhQzdKpP42QQX67jydt5VvMjJ8aUkUuPjz6
5/xO74+4PyKu7afBzeRfc6PkBYU60fKeFOH7w68fjkSqCXCtxBYTLfXUT0Wr22RS
AE9w41CAvFSZU7Zo2vhQ7xRjoePxac+NcpvuI1czOUqj7z9nbQH0caCJW+OJrgZz
F+ZxTKZYpivVIx1D+TmoZ0ReLUzSklcHrT/DoYR6mQTojIUM1hn3qQxuO/CP5Q7P
vJMXTmdJN5E+rfyw41kHjcjEcbBun8oSd9tTJv5pJw3J+ECUkvhVXpd6joaGmUdC
9dlFvrM2nPh1ZjSpq11f92qpa/GASGnokH4/X8mcQXsQ42lHZ77vmf3XmLq+yA+l
Ag2ijfufe8OLoBrJKQ/TFqjroJoqbw0AlHhFaRxs2a+uYsYwcxAs6ENmaWJ/fp08
lzljwet4nsAsFK7QJvSPJEkc4dJamVxUs5dMGI5Km050RFY3Ehs2GK/Vt+pDXsAj
rTdQdgTjr2LrXqwaIZSfgqkxoywAVWClxLwX57XjUV7ac7Qe3F7oQ71GAuNVpWtS
MXbgERfhB6s1Wx+Pvjs+TskaZJKML4U5GaOo0UgXYeZ+L28h4vY8bqVg9rgfd+Ae
G5mEfVgZsFwFR8FuxHxoiTIBuSBpWIfU7hbX76tI6Csh+/qwExt4FV4Z+yBan8HI
8mtCj7SQjnuvwAf+2qTGUR16w6o1j/Uue3g5yO+5mWNPe77TZdD21k4tw9nuoy4Q
ncEnvAE0UhtLq4NAnoyFLMpu9f36elCujvB5FpyAeqOHXClaVB4fcZXVh/xifbKb
uJnPX1t/696rGWaAAVzp5n/cVE5lMjKEii1mFFg7K+MxcOpBzE3z2eGgm9EGdM1Z
guxGSab/AndNTc/mIaMexiWOn2Kur80wKx7WzAOvdilQo/TAus6scd5pVBxnc/is
t8FhWFxhOO9Isq4FR/SxaAKe4uDL6dQTClC9EDuLdekYRDjRzHJoJZwjKiCHWUjN
Z7wlRTOTDe7sjEbmmFdfhUIIgmikvm/4V/g+tzdxVC4IGpiDk0hZDnXcsirGWh34
bX9d3utJmKYycAYHPygbqy7YVnAt9GCM41LBvgaEA/Zfs4OlU01J9cMnLxVWezIP
mVswFKOF0x2WqV+dljL+QCNAfkCUHRjzrrTTOjZBOaMc0tKosTSYeAnRvBoJ9wN+
r61AoZeBmNJFMQkJ8jAod/LpjIV8hO2XMYsuI2pMampboob5PyYIvYXV9OwZcwwL
biQE4PRdyW2tVeV3ekZL48dGW4KasYTqIL76MxbwHAj7UDvVAdu7IXKl5cCks1SQ
Yqq/hhbEvbVi06Ucf8B083qDNcUetN4VYRqHeGOpSDHWan0xzkPCtYVT9uj2dPmB
27yuiY388UxYaC/aycDgSP3I0hXAv9WUuF+vnArLx8feg4N/LhKl5CMOi2aluCXK
aAqjEBvJ6U3rzKLYs0uz5A6JtEloAe5JYQ1oE6jPGfeuKP9Idcq/M3a8nXN9ciTz
YyNSf+W/BsM4gGCKkSPil/vPzC5rXlz4DLQGKHjuN8dhEX71pfCgCydAcm+qe7E3
U/xMS5R0fPm0mCltXaWrifatMxDEpi7pMZwd4BsqlEGxcO36XQqP8BZxTlVArPs8
AzMAHt+i10ERIc4iDkZLwUDRkSKqwNMdhLplOirFsXWY0s07MBIPgrKeP0Fp7KbW
tbC2QqvrDcWpZhX0SihRGJBGUcBnj21OmszkJMhWkjknOCOzaLARZ2Pw5P61PijL
mwb4pql/lxEqs2jHKYb/u1mMJGiWGy6SpUCCmZxMAeGAlk58jU6STcrygMtxx8Bd
Tz/r5U5NFhprjxnzv7dq5ueBb1zJ8x+28SyZkhjJELYf3+vCgGQ8IVc3fCsv7QhH
epkGdQr/4mL4GWmrvNuvorjC2NL+3F6eUwjyPNcHIAYt8OZMkkOmTbklp/5E/1hb
NhtLHKZhAUCiM4Y2nTG+PjkL4rJfq34aUX9sVie21cmtZuzFuawOfhpmuks34jU5
qysnBoysScxlVdBGhWEhkYiqHQ9tMviegReXBKxtzHeuKS6yRHTql7lmeOLsUorH
Ih/3zMFN2oWSKQ8ASVt0Jd3SGm7ZT8ATwpvIJn/bkyZt8JQsSo40KtFU6//cWOLW
YUkhM7SEdHgI+WRNZUEKqxHIyxkHMK8PjavR581gR5QPwB5Gvxrnghk/bW/QDUR6
A8z9UwX+VCgmw/IeinGN68zv8ARzrjDYq+uTVjsM7TkSq3+vxXXwToMgMDY4UYNI
+nYsvb/JKAOTGgWYTn3jt0ZfjWXUBW7GppBKF3+kMD+CobJ91QmLZh5L1uBOBsG1
yKPXbC0Yh65x2QQ1HeixGGLslBVZF4+pxMRkeXGFE+HKho87vgEisQu6ovM9XXQg
vfbIny2Q4jEo500QJfpCxye8o0gmfKGUMECRjaZHKIWQt+vczmo3ZQEw4AJ24BSk
uvdfRxK+OaRX+Ft5822hkmeYt3sby0/lm2dHGPo2Ji4ZYjdZcwXewpZ7VA9KOrWl
x1+0I2NwQsMxV5Es+oTGuuOgXdEI2F1XIE7D/AR7eIUnedVq8l+tIwNn46cQpBd1
orpQcgiR6FrhSGPOaNHly5DgtQ+J4u7gWDUwJgyIOkqgBK86V7JZvNqX4QMghz/5
U88rzIW1qE3TZETBSu2/eIrTMupXAuFUobr3CnVhGxKGXQ8/2dFmA0aV+MazCVBw
uiFL8UirBtMDX32BBs2ldZiXT8Iwg6dfRYS1F/Is/ZgG/GrR5Q0ytNsJGHPW+ea3
tEyOLHFbIp6kgAnD2aifls6O1U91Tva0/pOkNsqTPPX7JBmbeOrBLtHERj+9KYEK
LG5gq4smAhJ4W5tOXmn7fUHqXWiT9AqvUb0VMJH5kkZaG7segAMnRNlbBFdWcLvZ
UPmhWlXAFBl1VEXaROYBIxyA5vcPqWrPCrDf46mGiY7DPyPSlTCaWhtnWZrOrV8/
o9QwPDXLGxiMOj4CawhqFk8M73vw8PoW0+Svotm/bct3UYnSjOybHMRM2xOXHhq5
ss3dqjG8hqj4Skmz1jJjpEyE677GWlI2tOKXeLQQSA8UC8cXgu6781uMmSv7mUIN
DRYP4GiOdiIEajB+pMskKwi6I3yWi7K2nh3CnUpod91FoUu2PD1PupvpNm3T+PdV
ITeRZ6wDGcE4KyajWCy7q2VyGFca2jV5r0FLXplxlxmuvtHj8QEd35gwhqHVd8s2
I3QsKn25Oklnb+7nPuPhMgCfLNuI1xe794vDNe3Nzzra1MC3HpTPCdO+m6BKpRGG
weJrPC6hce/VT9iJAtLSJhET6FsAbAKjTl2aK5YXJOfmmINnZxUNEVmqwDuhzWxO
PcwTAWEiSeywkVasFmP95F+A9NxMKV8CE8ZUQKA+tXW09Quheg97Ikix7Wq8fJvE
6GveUSeG97or8XHNY5NwyermJhgR0EtY4328HQvTvsrPR5bMc9B5f2nEFxqTZuhd
LPkTBiYg1XdhGSEhmmIk+zcuoIBjlLpIOIK4QumOT4rL5fKGugJDw2Zab/FOmBhY
1eaFZOiLs32CiAuN47APu2d+BOo02SXcgBnQ3i5Lwzg/TMAauGJ3il6vD2TYbCEA
7Db9cb0/CjqkKTUZ+CIOkI/oh1XrqA8PiheLkNxfPIDFw8CWnr5cc+dZaxR9XeAv
9Sl+hSXCIfmrx193lDQ32Nifw8GyzR2xSI+PN8cMwHm8v8wMxuFTJVrb4YQ6Uppt
/YFYZ8m5YFq6qnX3YmX7m+0pjJldxGq+h5bcXEX5ezJKk7CGeXM8NDgk3Enwl5qg
eKALEQvzJ2AfO7+2pm5D8OmEN1C+sjB4CNCBnAVxiUk8LQcbVghR5qAoH99JSuhM
C1Myovx1UJYBYOEqOKo59eu1SNAve4d7R1fZ68EHvQ0HjimITu3EOUm/RBKW+ffF
k3knPihhu+MlcnBrt8pIyhELo/bwQUzr3CIao/Y7UJt2wJrxYO7ofxkKrWd+tce+
445nW2FyEvZKz5avVVnbA+NNWWrjmCxuKmFp4IuUNXuwu7YsfghN1+9wkNgzxEr5
NyrmyCKlvgI4//Dk6RGDlcscfxNoxyIEDil1RYfKXwgA+s0/xQrO953GXIj2ZHLp
4O/vXbQtmXiXMRIYFjgPkbg+YKAnDsCu/1dKOUKRFGHjupv64SlS+Mc7uEk7s/Y6
3nerOPkrIjFQstNqXoOrJGrPzerGUWlnf/BFAtntNSOEAo6W8uUb/nX4nq+4nlvS
VVse3fEE68WENLRA9fiWCPyALG6bXsnuCoTlSZwS5DfpmRW1EMrGhx5YLs0o9dbD
bftkv6U/xuMzOP8BmVHeiiEqZ6gNToFNsYoRcLI/q4cJSSPgj0zVB++tSnY0xO4G
eFFC4g1YGaEYnWf4+Wb2afyDfRfbZxERx5sYvZj1opYqeMhARam6Z3LTxVdwf6Qm
OFN5AlWld1p+WYlTTNHZ1XVpCN/3/tXGoFprU2+GUTTbwRwlSyxDBo4fljHT9pzS
3oeWduL/q72M+NWDnp+4bRia2ORiPe5GUNo4z+zOeZEOV4d7M6BX0OtYHwg43vQo
DHiSsjG5/R3aATllE3syuCWKh4Kf6xAAn9a0sN39Tc7NsuzReBnHWxAhL4fvk+e4
O0K/iYclaTmjLsnJGMVtVciouf+BDo0/rJ6Hn/WTtzQx/hUgFYHN1Qqi7tMjy+yR
MjxBrAwp9NQZCE33y5Sgln2uy5Dnuq/A4JZY2c4CKiUZX1bnodIATkcwPdRNiEtK
unaEXksnFjUYcrK54J+EgycADHxjcQi5+h7sUcR+KOXg3CMAweohECL80u2eOSpC
zyb8FfcXOlznrSIss4nOKFgNA7JYbbSM/EQ6OUVHVSm5pqKYNRUZd8kJ+o8wvF8X
hraL5SG4hYqSJsSIc4qZ2JNXzzgBT8bSTpXEz+XSMoV6gJ2K1LSk+zxii1MgXzbJ
Mtp7RTakRB6fnFbZQscilOgYlBmgsyAldJAn19wvvc65oCNksNZjga4yceDjaJdU
CXyqEPOT7VjSzFygBz3FJ2uwcQOYPqANlZ+4P2K7XNTyTYptv4JeK5uSzlHZmSiF
jIzM5VKAG6bx87qG13FtviZ6hdYU5bjqBqZCCqwz1/i/PndNMVUUcR/651E564lz
ydgNNrO71GMbP7TIDh8/k2mP2oaBCJRPlG0m+Sxv2gveXgpCzIVAQ0JxaLR66SCD
eYhwduhFIYSKtwxk6aRNJWNbP7k7rgB0c7MFeiNTQyEVDTTM5mDmCC1yyp/awQ6c
P2aq8qO6lqweUdv9cEjW95rYcjN01Xc4Ih7pV1C+yiK5DMHE2RIU98icxaU2r4ul
0rOnGU1mys4zrv3t8TukJtovWqDzy/5ehDmUIhky2mx4Be+bkkai9C4y8Ff7HKxu
79dgvaa7ZMY4HvwOZqm1rSPdLAvxKWE1SkGLOKuhq7WpaK4xdbVCaEWd2JawPR7c
M3tac5TgWVhQ7K0pvwigqH46sDXjxE/nCtaNdqka71zLkDF2YHn34b4lg8HHsieU
qjYNbi4vQfCsGAfplF5WwANCXVAyR/NuIaD+zOauqT2Shr+bjN7pWrwq2dunckyC
UfCQUgpbDlDQh7Yt+tbmlhgOxPQSn9Uvc6t9Z1jRCNSIcs5P1M9k+31EuBmvhejF
7iavDKrLOPPmhlQQqwim9c/Pq+rgBqbSa84h08DTYalFnQ/dgB0ZCb/56Pd+pNiD
opIKR69qj/zDfH17/ky55njF0AzgbEE5pLJD5eNQmUEPz3SNvItR23pUSJnT8oVG
kJ7wECd5YeHgtjUl9n7jAMvYe3CaK4w0JcCwAUUR97BMFtAh+qK/OB5sZALZoEJc
LcA1cjNgz4ajO8qigBiTTN/klapuoz3PH5+VwK0/KamcA0TGKX7RH9fH2wWJGaQo
k4OoYdJ9wmYI4UIqMWc0IMHzLTplvyCB47U6K8BghTKtRb3Sr0diKlJJDkqyIG/5
Ytrl+xEMdPM5kC6PcUmHBbDUnxl1CBNr5tf+tqV4MSv9TF/QiLRXJyR9BicVbS6Z
PF6JDCkpe61f5weMZu/Ch6msTdKgSiNnjA1oogWBMKlMZtoDpOMBEHAm3BNb4QRe
TTlh+JdpVYMcJ+caVwdxk5MITqMmiDyaNe9XCQfCjy9+d2u7QTh+Li3rirxEEJ0l
maPcKrsA7jSeTT+bZ5qYs//o07XUUzKOxnXFz0Xqrp7WK85HC3gyo8Xw829E4Hnp
EfcyuIVFJc3PoOT3ZprZWxZ5nNf+VOS8Mc5+m5bsy0osVM/llZkuU3hGfAMzlsfk
8updzhReIt6EQGFTZnCGfATOcjNQLCY1JX/SechtZpjlZBjCrBsoRGEXTHoamdnb
H3w7ncdxsfYJfzesjbv1/MyunhOoY3j+SMgc+v6qNwYiQG8EJYMuRUtmpujflwdD
1TXLgeu9OQtFeMgbWS+aHGceROXhwZLonaVWtFP/cAafJL3e80v7V/m+aoAygDa5
EphOotr2KvgBDDiB+w37rN4HOpEmfFU7CJV6VS46guA8Pon7S1BuLbIIQCxndlvz
vr9uuV/arXaq7yKarmNayRqayxm40xIw8Tdi+CjcbtFoAHqY4cq701H+hram0d13
cy/7JhBXVK0haN57HI14WaHBzFfedemAAKSR1CJnBhO/vbDg7LvvJUYbEOTpnyZR
YVlXNaWLsfSc1d3zKvyv6HoGtSdMoc7yqZwbsQQdqwTRbK08QbxLAm3crwN24USq
0ok+Fc/QL3yjnSW0mGSTMXhenkTsOsdKZRf38dsDifuz/jgPjbqzxmjoH2C450j0
/KPBeqz2rjJZ0u/uLr73BnnRF5TDv9YEsJcBdbbvTblBIYV5RqP0XeAddLcYbmjv
lfM+aM72lwF1yQymk+S++NdZf66inP0Mw/+71t+YxhZV3rL+P0eDOvKNrDKRdDR0
C/6kNXjalXwawgu25ZyX+100SgCTV75xNkcXD36kn9oQRaNai4KdBNoZAQUS3fl/
inEpzWqzNxBH7xPsaiuSTPsip1BNJUW4oO6wvtJrm9vWeoV2MJvYSvcgEWGgEvLP
a1rzAGQvPt4N4kV+AGK6tmBistU8IwaspzdGewk61P/tFeeFvhcGHmehlPeVEMhc
nxh9ll9069nx//TQzdtD5HSmBV0cbRAbhb1ja4+yeq5qFgoZvmOScZVRaVF2sb56
ODcxVBdTknrRhKoC8AXsAE1Z2gx7C1VMcGDpzpJcSxWvT8Xw4z2pLEhoWkmD5j14
W9J9WWRCqBVq9j+N7kkBe8lcg6lGj06DGIy46R4fTXoA2NbpqdVPnKbfDrhhzeKh
QLRpORpUcIV/1ckPn0w/JLgCkLgQRnEYWKecVbpc5UOCu7B9Q00R5EYJrCyfqC3H
SFf+3DC/V1UUjZPc6vJ9VrY1yJ+m1GpbDDS+wFa6iMPiZz95XavnwkQQaw1chUTS
FqBmlMNQHLS6IebnsWKsLXRj4AWD5v0IjBSX876DELiGlnudn0a6k5tyNLcsuNIZ
4pFFC5Km2AITolP4fnrlaV93ccULTEHVHLno1cXGbc00+8ZS1vbGs6EpZlvmaUU6
ERrvY30LW6RgUczEONpJUPJOoZj4S4jYJdoTcXdeDFWvMv27ek8vAk1MR/hRoTQ1
pw42eCIcAHO+nrjv5ecx2KGso0/yhksQ3O59cPVmKibio7FeeJ0ZsNCTh+GZKzeK
Q2P79wT1i/RpswGBN0crkslshbMVJtc35GdJ1YMARr9BlTwydtI7AYJV+Mvrva99
6wZueLFOVmgR4eVIVUPLzcqBRk285kt4Q9bMmfyDaz/BZA2LzY7d8DTDeZqPOWbI
E3zt25R5vppZ0hzgJ3/18AQPuj7eiDJPEan1Q1n8P0tY3FyrW5vu/+OXAsd5swrJ
yztcByQj74kUV6PIxfmgoIRiTzhUH1E9dX/dFh3t9SGVpDNYOE1sfo3/wYvKDLRh
UjxipR6D5WRU66hTiuISlRFZ1GEka3hw/5YghWcudQcfWg9QCuz0KWKg+5COXS4F
41oT1efY4HlC3T4MUVamiVOgCxXDvkvfYYBZu+jxafsuHCFiQIuCQ9LfI6oREf63
8LpWPyLpLD14yh4b62OS16lBIa2MXNLo6Y0ozQZzTK9Twfa1YRFqxGr+FQy0h5eP
vGSdey46b82K2bx+fazinvJYFeYvND+DnMu688RgXXONQ9sMIaH+H/yp2K5et1O2
ADPJT7GPU3YDJvMbYZ0n9cq+bxvipnk9MD6ngd0GXM4y4v+QJgOT+9q2BedGTwHC
7Flu2UMVXnU80Rp6pUpsc3oiJtu/Bf6XVSQAe1ojfZTubxiKzWsr08Jo/3yx0Jcy
MuoJcC5i1wLNPZX98Rg5LFyD7I5pmF/uI7ErYR+VXQVIskwGKrUrD+gSjTV7+e2W
9QV/xYmFCqQ8vpBtCNzEvOkJlute4ZodM8tDdeyGuRBKQC47aM8C1eRHCeV5P39U
IFMLGV/aOoJEgAc6mUMfKQ6JM7L33TxCPa76xCeQg7CaOpyEkrF6G9dhMZ2QEnFx
b+ZMxDkWDHi7hCasgD6PSI5c7qr6jqVy+3ABuRJO9Qz3L36+l4io4Y3AulMEzRBp
KaeaYbsdLAIq8K03G4HZcvfjWxvoCGhDyleknO6IaY8eIj/rCVOqPU/Emh3N2Qj5
vXGxrdrVR3ZW764cm92jCnuGvwhdyYiXCL2RhkCj8DsS6ay4pvRCEYQHDJ61dYsg
cQAkXvvtcFNaY8/y/zcozgYhnkq/4GbgKhEQ19HF76bQijmxfBaYxbOJ4JH7sIOn
pObOGZ77pYFkkap7ZXVdbi9rxhS+amwYpdm1eSB5obnZZI4XYkPbDxgihkRz4MHb
sljIEtw2xQiYhYRT0U8omeQ+B1O1qPJlsAHph+xJCIUzEBn+U/lMJK8DtASSBeuK
KevywZqF/syvmj6D2B/QhrNKUoou29t42DTD1TcU2zg9P/aHGmqT0y0HjjVZ8QaP
8QmrF/fkzWtNJ6LilfBgj5AdOP2++6djACa2jwv43pfchBakyzOOaAWhmaUfw3PE
ISN5DtcjVym0BrSZ58S/e9BDTHc3AccQDPFoN30Cy0j9ULY2Y2XU2Mrbdu3AFQ/v
Rnil/Q+fnqrYz5GBtfN8k+RxHlM/n1r1mcz3eh10AvhvLa/YiI8iVG9uTVF4gM7M
wOG5ahgFENKC+kvk2ywENR9mHHCzJBBilvwHdgw6w/OSk6gb6MeNq/rhv1v4DO2q
cxaDyQkedjCWEjd4E8p27bgzOGxuLfiM4wybX6TNUGpt7sGeEyqBblO7wAqNwPUY
uuec4Ky9+8GbeeK/K9rRGi78E7Y5kgD+U+vGOgmrjJGDwdtTy+We+6cSMB5enFVk
lXmW2PIYCz404WuZkaa/09lDa321AvI7TUk7qUfu8DgVFhoII/IWN1qIKdL72baO
jxk+SzUraKNf9a6Hy1k1NuoMw/znbHa2Cw4tJFlTOfgzZeBQ5mDAkFtNGJ2h1xOm
9NEclCk1vIP6vXOc7/4iiQJO2MWQsClzU/XweqHwumwNHevVDqlYL5njHGqe9y92
zw4+RjDkbzU7U+ybPzRrusKTE2DwKn75nHxS11h/6Pb/09TwOWCdCDvYL/oKehYx
3xV/XoGUBJtoWu3nLxdnViUu1H9ZV1MCr7jkv9l7arDKRiKDzsdZtp/F1Y5zykN/
kqULNIsyiWGIPW7tVWF+feuM/CWqegESRyrgt3SmrEESK/dkjBh90ibhCxYy9k2W
tWIldfR4jD8kTo0jvivXdQ46jTihSmMzSZ6F+ormr+fBb8LnAFTRTweftTFVtsAy
prlRfqcNAmbAx4fGWdNZYjdVfRTbGPPO+qj/xQFbiYaBGNueKUy5AzgU7ZgVYtH2
duAbKa2o4cIsNVAddoXk1SNDCgnYSRU3lCmcDGGFElYZgx8cvynuiunDxEA47fgs
5EDSMgFFMMGS1af78uy7lcDA4TacsWumESisv6peYodkMKvk6XlE1wzTxBRH+zgq
S66PvEZn4LnV4jaUFQsJiQVsXdIZiq90HUjKehgY4346Ba0P/2SVIpGQs+bZzlPc
dGEToQUozJEp3UrNAkVrgMhT5Mpxx0BN8Nvjc+du14ihaj9P7s8REIYsm3JXXitY
dYE0j/2tBRpj4c6xAXlw/0haHLhnETamsDZvE96JzLA01EMcVhi43Nh26OlEZYwQ
VqbZLpdV/XLgA/HJUoAnKIQo8OKAkapxTwHPJmi141IFz3EtC2CicvgaEtPRZDLl
X8w/qhqSOFQT2RI1GdIsMGyVdC9TX/HnP049rVeJzGkbJNyrQZ9rJDF+QeEW8P6I
K28WtyQxe9kPFl43vj40zgE0+N4nnNDszYLknlc3795KY8FUz+dsSTDNgwb/RimX
P7gL6aEVMMIHtqroWI6XQjCsacIQTblAKe6CL0huqwlhLteCD3T5gGeI1hnXqiuw
1foI4FX5Vujs5qaYOlvOUzE2F5wV+rNg1gXCII31jBtTTa4ASEgjRqg4ZuLYdHck
rQN6vCkE3E4sBzku48jKHHxuArW9wXRypX6YRzfJ5cXMo5+Pak2S7pnnlPk6bOHi
SU9Af3Y5BqNx0+sB32bl5LjHd77tY4LZZPl5/HHG2DWiVlXIky+EaJY8C2YhZVrL
QSTKUm0mybGR/6yTbCsrxRpGAN2KbFS+7wUYVSV0jluqlc4g8Zx27SnJVVyknj+k
VHJ+jNOuwMni/rQJ8VSggYjeudvNmBHIc4ft5YDFYLwom6sWxqhWEDiXn+SkH/nA
e3ee9wNBBZzWY4pSwPF3WBwinkey0ow9/Vf1ZUNZQBZXEMmQxezEnEE74KCw5KyA
pZ+z/R/Lfli28l8KbdQo9Wqd6CvyAmfirACpbGmUM+9BvZzHWQ24WKOsziabgiy/
jt1xIuX6szTB7+SaJq0LYrWRxM7z5ovV8SzHUqEmPA+p1JWFH261J29F88tB0kBa
/ZYeYuME0+SsKz6xSvFH2X2pcWSvNNumg0sZBdfyu4J3jmTVCRGZyr4SraNkceFn
ed+BJucSY1LsvXAQH9rdchp3FucFAsy/AgS7EFE0gQZitiA+T7oIc4FExiRdRhgh
yNi0R48qrgk0DutawWK/zvs8Uv5PwGg0/tiLXJZdULz0mg9JxRICtl9PBiKBrOxe
SzSBKQJHJk7qIDv8uUG9gBDKPZMq/tgpnQuLmtPZL5YTDDvhY/J6kU9VRYN0LCYW
aZ0EjgonXfDZ4tCwNmtz0lxKA0lr0FvMzccILwUPZud/Pp8RX7n4fDJ2NEz8vtV4
N6XVQYr8uQBIyAUneRLgLxbJYdTxPjqE7yIVIWEgg8l1SlRqMx5TjniMqaV6PT7K
3u1ZXmoQb7f+3TQls2gU/ByqqCuVXUVGVHHAO+OsN6b/OJsYC4uAwcf4zS8dKdGY
QdHg/pe5VnolfrwPl7oTZbBBXptZ0IkEZK8PKi39uoIxz+eaY/M9QmSLBYroP7L5
sf8mIOaRfOeeTMxx7i4nok+Pq/V4rkGUbzJTLZGiUUSl3dfLHNZSSjQGhABY3t0O
o2eUxGDsGcSPWWWsTujZtsIej33hYlL5i4SwbTHifpkgmZoHlVE4CDMljTlVE9F7
/w8y71hJ9DnTXJvJbwJdWKtCvrobXFAUri+uPDJPbtTaDxihX02MO2sYO8Ov39Qo
C20Acwfm6IvQCbeu53W6HDOWULaziI4g2nLtiaB7tS4E0aFd/Xs3oWla+6nSyFHO
7aet3ut53UghKUYphJlGiUFY8dz392s6gZhKF+V1o4z35Asc95pYFbPK8eN5JKHQ
dWuCXm+/qr5kgbefnFt378l+x+WTsBu0QH4DRKOKEOriKDf62sxfqw1yGk1410hf
xbGrqCpNq42jj2eMd4mUsXRChdnD+XZfmtXRr6I7xN1zBcELY9qR4/j2csbZn91q
nwHdbiQTXWPBwr39fQpr4FqeSQOmpUJEoFJlXqwHlkIb6EAgNKJbX71TN7QZjWKQ
kww/96x2W68e/xEFRu1DiPQt0ifxHqFPNEz3M2pZdgXLc1P0ltN38HCPRbW3WXY0
BGrk21VxkYd8q6IVcyjNQw/YICqropdk9hEzNvqul5D0Jzbkn71zPTOL0g9238ya
BZlELKdq4WdmrpB0fkloFZ+Rn4GUQc/IowlULon0ytTwtVlNWNDLC51TGHo6cZHE
Rad+Q9huSiYZNDePTPClWSjeZknr9qPhlFFTL5AEBTHCGwSyG83IRfJbC/3+iYp0
PrJ3VNWL3Xqrb+2FsEcKhoWoiT4/g1gg6T3hsvKDmRy0M/8KgFM963Od9nNGGh6i
x15fpAjGa3SvsxFyL5RY1ezb6Qcz1nJZltiYD/bf997aa8HxQC77Zcq1qnStrNFo
4bHZaRHcSn31zLqxD/tvwBno+ILEZfXgdfDSzw1Aq0VKRu3G+Fc3HYIEjsrWqSvf
kz0C7dvMhpaeCuBjD/svBjcHoVEi2g6fVF3dUeKmXc309E70p6V10SbhhZCWaRv1
+SyK9nFsuK9hMlFYtnfYe2EHBTQ3Q3bJ72Wmh7vxD38jnvnp25c3oMGN5j5SUcaD
+RL+qyMnbEtuQmmMCzp+evBpa8FnfL2lVcsls0acvPb8FT53eEHOayOsxG9pswvt
ZsgrTz7K09IdvmSr5sH7WU4oqwwDJvipkdJ9Pifj2tpW0d9bRHzNjjeNtdcZ5Rnq
vXuvBNP16FgL/tmmJN1zXFsIdhx/qcv4zwu+jFal2xJqQ7rLK39Gnw6B6lpJYgYw
ZuS0YicSdJOaUS6EKssBls9Av3XT8G4dQmxa17wed1NMuBhn71+Dw6GfVApyGBzy
TpyQAdB1d+4CAczH+rIw2y9nmrANpkD8xsTuBoStsxoXMwdFbsasiCclM/cv/CGC
gd1FXJRe/00C4CG+/0HBaLOeJv5uGQTZ59UHB8U2EXMf3FiJL7OS26/4yxf5Jjrl
UfCh674KrEtNgpMd1uUDftr/SO4t06h7ynARaY/kgPppf2mcIEddP2B4fbxIxcs6
ACdmzjofvHCRUIUPzySzvK5t8ThejYiTo6jhuKY7cgnoENvwKQRaFqMXTcHantTw
2hYnGRTxIhPZ5rJXQ9ErwjKZyJqA2lWjSXm1JYpqYwKWWcG6XkXnrBJTXclbFoRq
RzpxwNbe1EnW8fhvCsql9l9nOUjq06FjePQ2eAPMEi4fgXOEOWEKodeIorznSV20
D806TA/FvwCGrwWuR6UpPApDE0DDLhawQOPuMw0+G37EdTwT0/HvL6vIVhZUJc2W
hBb+u8y6K/ibwe1pthVtRtl4HZPvxavySVMovnhihSdU9ZAQyGJGbrNmWWpxj74E
t1YvAOB+twgeevGYvhM5AdXWt1o++JXCSmNmMlIHmpev8sv/pkhYo526OAh3vu6M
IzkE7oFTOLj9QyRPKMylk5PF1QRov3VAEeTGOuGpoxKHs2+VWUZkTXQGFLkQC7Rk
iemLIrk8ksClZmDfIfJcObQkxrpoLbTR1tAq/IWC1BshB7lb1cK8IF60geutdUfS
XAJlAzwyBWCKweDufFjv7GGFfC7KJfzzlctPE1PiGWVo0M3tSE5yUi0g6ld/LPnd
4qzYgIWG6L9jyynVIFx8VbqvPpfSeITASyHm1HvboE7U82tffpllIPWffV42jzck
8w49FaCeYJ0QAxptLFMZZ4hmytIqwYweWT6+SUXRO8I8C5iAjMDQgaE5sk9TKAmT
mJKoStjLCsZt+ZWgr5AdSkN4ITOIHcBTIL6GKJFixCaGzu1G6SpiecWe4Duiu5Df
xn6B6Cjh7Ak6WjLj0dSfZ3GOB1pqJ1oC619nEYIkvbZANpuenRbyNFOCpGBKCWod
S9nI0s3moDQWRI4aJ4kfuyHW/xJ/aYlObKj9/nceTxo9/uwr+3WzqJcpROOVWvD7
WyMWMQV3HKfNUcn6tRi6djhPw2Jp5XSqdaJJNHaL6dRsv5Dv+Y5Asc9ippIFwf/1
kcTlIFQW+8teP+K6h92QDlc87QDl4Nln+/8Yqukj1ocOtnJqNScTL+ZEgw057jJZ
yvzXRmkLWDulkkfk1vBQtUsjX21fd4sJVKN9GNQRk9WjF7rIox+0ALpudnrYUG3m
9by8xgr1OM48ejrpE+wUxlFdwr/rIHzEQVAM6oqVOiMKKK3L57fFwJXdt1qhU2+J
0t+IgwMOdwCEKQxsMagoWi3mesCrZ3SE1lOO0Nx4LilCd9yXWdzbkr/pxpBLP6aY
KqvxAt9tpr99OSmS2CWLUow5AYQuEUrA0ttoY79pKOEiPXtMzYfqk1k3UT+kLYzA
O2D1nEkXlATY1U7FqJNsePDd40LFwFbo4f9DHSX3RFg+HSies17u6bXM9lNdLv+O
pcrF/JJOX3gNWTSKOKxaq8zmlfdKKcu/nt9BS5vcd5o/N6+HeYSqHBdsKCIeNtDu
MQX8Mvw/Nnc9R6rBvAOfkwaptidcue2jmLObsxY7Li6pfG/jXZzunlc8/S6YVOBX
Z4ZS/bAxUBxFU8mdoetSCFXC9XUZ6b8QPdMOWzG4imnKAlQuQVAkqf0GyvMBTvsF
nhAHjMpVnD2mqFPIWWqFn4JwXJIIJYqwYp7g9If9TvDRqE/VNqmLlngFU3MZHzOa
MDfT1UKm/SGwyjmx+efJ4Pq1IycCmPwgGeTK4fGrr0H7J9bAyZ8KvA8iCdEHhpyr
YZ9xKLhT6UxuRportqi4AJQug2k8IVw2YAxyg6vy8RH+ck8yn7lPgMKqEYz1tlVr
yY1+4QgeamonxvMc0BifpvDLEfwO9mwu/rsJAPR1aFlD95vGG+8aXbsgK6YEYfA6
OIizRvJHNM+c4nT50IvYvWH8YosHqpBcU8frC0Xxoc2lHLQ9HVdfgiSywLNlEuwr
NINB7gAHm1bL50IQPcerSjjNUOb4vH8/0NSJnnj1Lza+iXZCt6qjQxhCbZdGJG9m
clhWzftJQBfJTY7jShAPF5NYg6n/lXu/bO7v5kMlzOtJjkktbXYUZ3kMNUa2synB
gn40kaP1LJjQ2mkjDpsbebMMzl4kCYKO2rSj+vD79/W58QygHtGHZERc0EucrIRf
H/ed8snbeRvVp2ZMy3MAkOAjjbchaLfgNxSeIzfOgZE3rcgEfKX7LyQ/pRpFAcuO
pL2pUi5QR7qG5ijI02mrA3i8jIh14UqCbHG6HDRAwTEG86fGbFEsjMIiQVU/bF0B
2wk3ZRdRyeWeSLm0HoIV/byDS39RWJtJDxf8oXL7isn/Qv3QNi0FI/9FEcW1zXzy
QsTATAxqrYHcAiLy48tgS5sSS1D6I0iX2U1wc8/PlAsu/jF1V42byv4HPB97BH39
lAlccvj+SHgSlqrIiE95nFqYAOIouIuMB04psA6uRTWNX5bdzmC948RxaYSBzkuO
nHxrlrleC8tDG99Gd0feptJoC/yDCFXD9OzNHQ1hfkckRja8OgpuXjtQz5WWI89m
6aeSCHXMaLG1aTeLlWHO+n5JA0HT9Ipkci/SeqnmnERYkwdnjqw5I8barzsZgrHF
OfRK1bLmmb+ONcmsW3mkulhuxp3c5MDsCxF7LeyFsgBnnPofGGiHM/HsWj8efcMX
qsl/Yi8jk0PEwFgKNXdflJ+ZTIroQmz1vDAkwPgs2AHv2RsgKaA/anQ7Wt2L3+vj
/AU/nbK1ZBattXhPO8ShpK9+7O4KqrSEOksFt+zr0HhLXsUqaP+Cz6HeUEoyJ5LK
uy7L3LkqrvRCYE71hyE7mAQhOLSQJAALiqo/v1vLXC+JQHUWvyETCvq/SPKF582c
Lva8LyLFY4vJ1ed80TLKgRAD6yLoYIDtoVBh+NMg2wejgFswSiErlp+j08HILJ0T
OZW5kvBQX8ad9/PcG4cstgvtlbbx/3WWSIJsfavY2/NvMhYD9/UE1DEfg+LSrHak
G0/4eagMBFW3T7IA+XwA2a7C3YXEHblgQOqzirkHCadKStXhIKDmBvZUXlHhBZrm
qlA859Lm93rRZGOV8vegl5myanrXUyicwvdlvRbgy4dYIHrh0qamr+PIYWFjVd4p
LMWIyhVVw7XKAT7wkATsoWaB7Z0raMNta32e1z/C4czHzJ8uPoj3EVaYWwa2qtOT
qyHFBMHN7fy0odkKDMl9Z1RtCtjl3Y3hpemKaaSkCbbZP75a5i8eyg6neUQ+SLOg
5q70+DN05gqe0O35cVpBTZxI3SvdRbejAvV+1wOsCyIh37JCkO+8jDHeH3BBMHhi
SCacS7OOqXIoEzre8cUjXdZs1z00mBaRCA6op1AaORMzyFT0pqVKhgQGH/MYmzIE
+SbcI7Ne+WypOwrJ4W4GO9+MYAkSMle8Rm3tDFbSrbHTMk/U3eJ8M4Sjhtw7JNDz
7xZ2G4ZCs4wvYXkEIKCTGmBYibou+itaxaEUtnN4hN+jssQrerBrBsAOYdIEgRoM
JzGcd0J6L06ORFHyjU00bOLIXmtAi5eN8T+IHUcMKxuKkCCdFlzdVrQmHQneBBae
SdxQMHJrhF8m54assLhXB0kuPViXwIa36tL/TcBwBYZn5D01t59MpdZM+X9PR/hg
EUrD2lHej5lsKowWQwKl4j9zdb21A935qICfvpcyS6qnLY2RsF4ge/2H4cXoCEud
J5WRca4Fze/w3x7PiFaNn+fcTaxo9w5iU3jzVmHdLXKTTdS0htW9zaYiGgOukRHy
Fo5Q1+JVmnm8ZcW1DVHsfDnb7/Rz275c/bZgOp/amMwj+Few3YplF9FWnZvDeRcQ
UNX+5kgcZhwT/E2vxE8eS+eQ1oQNf1RBmBDvqshczor956AX9JejZPW2s3gRKm9d
zc6u1DYqm8Cg6jtg4IVkJV6xs7Oic3tJ9Ezx9772YLowxAcavZ8ly5jr/hT395Iw
YpXE4o6EUbu/elolr3xoVxMWqzhAQG+fMdbCywh5pp7oXMnKUjX7tza+PHNf2k4X
BDguUmwJPd57uHY8089KJ40emRlh137rN1J7V4D8UK9BKCb3bCpQMLaA2BXTjMhK
38PF3nmAhbJ0cFD6xe9es606DKmo14WYh2ZvFooSP1whtPU0rsvs6ciVbglLzgxj
5S+DEbjSvstc05E/QXgcG8vATVvzxv/7jwDrTIt2w1Hvt1OsqWck0PQ3SBL5LBfd
QA7Y55hECbRnhWL92TClo4pAeng8gIvDDVuOUTcMecVA6MUMl8IZxO49mUVGZK0O
fzdqSByCBh0PLdGu41Cu1DvDZGOEVgN6PH6WBeLe4b8POHSAziIpJ1xINuzMjSjT
tjSiOYEm49o1BQBK05GCtAJtCdIjP9+dbT40TLE278XZ1SMa2ChQvTMNcS0HS2JO
L7H/W+9Jolt2zPCSMoKihs0g8OF3R836nK804J+wYHRpG1rQ0dJ04MaZAxSddCDw
sh0l44i9XJE6JnnzeVBxpGmwyaK/gC5SAgkOjaq7xSeC92IO+Zh6qxRR/hordq6Z
xhV+9NfB424Z12vhCK6Q8wMXjQTaPB5y0lqVe4GZhZslbrMFL0MQioAjPPhG8Uyq
ZQNJoBCxw1q0mTmwywaWMiJpt3H/K3S18jQN657syNZvMDgOjG0/K6esOq6eiHfc
V/w1E+EB3nI+SwiXEChRXqjtCyP66h1RqOGNWlrYt3ZKavk/biJgDhkaCrCvRt+i
dljDZOSD0nO5PaibXGFDbO9JICo8kfn/3L69IKWveM3vp9FO+sNczTvldIb19PHs
MDYAC5iyw8+Ptn3iGuKD/Kzjrg8jMSDwcPy+E8zjWWlmFL+Sob5F7IxspC6l4KGT
fVhJPJTb9Zx3Tb/D8+CbsSADOj4q99XzmUuyzO+DLrYdVmuWjnyQN6+Qi0NSoU0x
YXu4D4Y+92aUz2ZF1/ZCZQElsvIgTqk9LLPvhIV0Ozh+j0kJ3PJhP/CBI+yY24cA
keKEXn3fDRlvm0rK4CDwIULvcfsFM/CPeHrMFps3ZmN8HcKMo5gdxO4wnSgtUyrR
A494l66wmcErlXyl3XQyZyTAr9FNgmCXcgOu6XwshnIdyjGh6l51Kvu3N2tAiAH0
EiHhFZdkLvs8grzA3m4JZGk1eVZ5SGNhz8Bp+yucQbesr6aZ5YiRGxvREnT00wAS
aFZE7z9osxsZpw3NtmF97mFx15jAI6WzXO/LTtMPhB6scGANqqP0fcbkkmfD0olr
w8pWcniIT03bVXr59wY5eK6rivyisnF2+dZH4XxYRfrNVor29FRji86cI26HuKBX
/g3SCMeGIKvRd2NgciybXcOiTiF/fNsIpO2LHjRb5IbLVnGjbJ4Z0z+slQlApDkV
EZ7+3sVkujz0jwnQdZHvftJ5HRvzsxqmntsF2E5xmR3jiPQkTWpS1Sx9lVDMxS7O
fYAiB/Dn42jZHj2+sSROE9rI0yWujONCprHoR3Bd7Y4lpHFArgR53by/8mGI9f+T
XHD8qyiu/lqfmIAkhwfkQUZsLC0ZMYu+Rv+p7LCJz2Zhv1WbQgU/Fpsnz7Ulmnzu
xNr0XNlaF9e+bO9vOVT2qalVJVTxRnyFjqxF6NajrP5aoLkAk4+pLy1wOcwGzDZ4
SPcQiVdKq0Jb4yLBIJUYZ5/J5cGCkcki7mjzGBKDTRVVWgHf6YVN+nYwePKO7ORf
M58VZEOz0FVsFvDiELIR2A6LRHgui7UJleP5RljCLZbbgMtziGYzwRBeLXGHDrS2
2L1WRAUY3Mrc8nFD2ifKddYs+Ua5quw1ZDTiCoZPrnb3cwZsm+Gn+x/kggTPHr7m
U/hIMlzIAQsaFjRLtjqKScVnZhl2VFrPEu+SDXlp36UvtHbtGZI7cbneHhS0HXlr
tRhNV2v5unWHfgs8i5UGQ1GCgWiMrCWsOH+EEbeNyPnTQ9b4Pzu72VJr2NP+QI1o
sfx2Pld0ouuzad9U1dyXkE63gptwAEUefBZi4dR9RyBh4GeAMeEZMnv6/9mAr2B/
hjCRIhLjtCHzbCFUNoW6S6o4WhYnAisYlpQmQZCR9pLc7UgaHdNm5vGqdFh7pKKf
x4SyIcFgr8Hu42YT6zAWOD9aGPCuWDcXAB1DNrIRA5oXiazgj33MYmPW3eWeIFQQ
zZqc0Avieo9jeV1Vwj7tjclij5+zS0Q18Z0noA3iOJmNiNR7RdVcGL6hS3TWZbb+
a4EAGLk8tR0S3KVRqlXAYqUtgScSCMzY3F1UFVu6J+ug2pkjb6TAwcswTkvILcH2
PizL5HgOyLXwR3yetEmmiY/hVM7UTEJ3yvpucjePdgxxbr8MAVi1dJiA+6/yrxbv
DjqkwECRSJxibPKuJJom7acOCOKPCRZE1P9vWPPPif67oFD2uqx96ye96BomBdXZ
PduCJuXo6cOQ3+8reePHO/WCLaF5Gf+PwdfGr+zl8kpBKdyCuqQF8bLCOUzfeEsx
nBs7G/uNDaX264U075r1b0qFaWiaGLLfA1UMOZwGAS+I+naA4cFvViYmgThbu2QO
JX2OHRs7YmURM6gaOD9bGeAQJ3f2iknFqYy6XZImtXCVSvV1AYPFH4MNU3FMrlPA
r5U9/ZI4AFKXqCQ9v00Qy2GRmmjgfRwjIlDEoUWE8nbNgjEfGWO9FHvrO1KNDWuy
0cMTH452NDoeplE3CRvPUkIAy9VxCW4dQWvK8QePXULqIu6o+vCQburGp1f1fvRu
SzIgXNCIQDG4V+v5/xadg832vNRcgBQK9GPMnIb4Mgn/sIb0DbcsHbgmGZyEBQT+
4Ukiyrfd/S9FcsVwjAqoHBmGCfldoCkLPrfVyc+kYuo/bYPLS80GqHFWLi9sdCRN
GcxH/X1fxwXKCbwsxW+2bD4Dmozj4ljMv3v3A6yKZbyHjNuA+FmNJnHd7xZVhMJ9
Z5t2Bg+t6jQFtiXHEv/mP6LsQexpFodev9edfhaEXGvLihm8WBHimZqguKyTBA1Z
VcQKkoZKIQROyrp8teVPUavGXSbd6abRugydRtfOuE6yKu6PjOdHtPTrEvTcEafC
JWxtUEEhSNLjm0XWtjRUQzojUVWtN+2EjnUEYw0grIu6xBRk3VqZMGipbCzMVb81
9KSYu5O8C2IU+yj8xyDLEwJm92LD9+KscfO9xOwy+ltAD95idzl85baRPDLQt/gN
bkiFZrIM5hYSvsvOkLOCDQekRmYZO1LF649h9fCP9JYqUYdItTIyw+gA7VbGBFti
YcQApcgks7wXwe8GQffiNcK0OdFtXYcrkgeK5Ois1FvistJYY2gAWAwp2O9eacjK
UO6gvkBEwy504uqIVb+Jv9EZ6MGgFqJp0nCbKgmC7IOX+YvE6gEf+sqZTL0AvlAg
t4qGuKkETMWiYRHcFW5Mh9ciREvh+/dszUDnx/W16owaJ65YDptGrOWtDYHY4YY7
hVRNUiBuCdyiPXzLmD8yVOcltBs2KamK0zX4QvVBj7FXoumZ04sS25pZDe1PE/J+
kYKyIwS1jYde4OujSKm86JcbnUTHVHG5Y31bm7j5y4JCslq9QBJpbT8rQ4lAw1Ok
qpOgMRqpVuA0mXwTs7PVPTmP1QdVafx+eOdeiouoW06EyROFYk8Jz20eENTWxms5
aJUmiqop5QOtwlkhAAPWqk2KSfhZTJUY5LWFNaBmGzt63OBaF5Mu8tCxCx1WZ+OJ
hrh5l4O4hwtdnrZtBUExYLieaNCpiTWZuM8rKp0qzxHAXxOPL6UbK+ZrYZewR5pa
mybxXnd0L+TDvwmeO7lL/+LRZfiHw4g7gbvuJKo/pt30nmoHD7PJWlhIGa5m2avu
T1bAa46nbKkJkFxHuQBK+xGkIFcElLtg/syHyAKjgm3DVqcX97e5X3TVpvEJbbWl
KEbyKO2HUOSVC84slFz6jHTe/cxcoSwOwBtrmpJce4HVcz4+6kSzxYvs69GRHox8
tOlVnbDM462nKBPb99ZcXKjQ27uCy6c9y0bzgGKl6Q0Sj68JzlSFc1wIA3ZHbVdV
8yClu5BM8/VkvjtT5OXaKQCp9qt8D1CuTw7o2yAKnLEYqmhoWiFjJ+A4g6aclODW
BXAijUTL0GYPvoRKh0wMV2ZuQqhQwRDwUSihhhLUHUCfnXEZKlfeZfKdQ8lgUGO3
Lk2lzKS2c22U2qHXxfIyWqgRIr43qhMGx0vxh0r3UFbTI9Ll1GzyY/6tLPJAXcGu
6jdvB1v61tnZsi+Pht7RO63YemLv07FM3Pv/X3MI4cNarP6WhHvUgmOfjtXE3JHl
6jeFf14HNAAnE727+ggM/xLIJwgbYNV1fLznli95Y+bvFoMFiU7kycWQ8CLQ2Nty
DOCRiWVYI7ragjRtZsHnjnVd9L8e/XH1jHKWMJycqKW80K+3SHFjQUVhTOLtGAt9
hpMuHO9K397ZJZzZ/cT4DAmGuoESK6Jr1HzBck9MEWqgJue/R2sVGNPlnfSpIRZB
7pAXc/Z6BWp478uVBCw+vMWq9bF0Xeo4cNUirkmKEkoBwbARgBDvAGpbLRv/XQUd
6SV4W4+gBK0XrFo4MbA/Jm29RRE6Y5+rXnP1X0/0YIXx2BKZQ/J3pjGBbJvxcWVG
CzgIfY9VpkHldgEMv3pKccEmfe4yzJAOrsJO5EI95Qrwyaj6mZSeCmJur4+gFDCq
ZMtoqsVB9oTe1ieT3Tbbq+W2ms+Feq/fpWjX9sEWfnyJhMuoRiWeQ07puA3oc2RG
MIcj+3Ogbo1iw2WDnaWcAwPCzndfpgFNUOCXfhT5bs5IWNEXCzVBe30IkQORgBBX
b7aA/xM4zUAnOGxe1NgX4MNAfZDC0WjfpE0nTqH/i88XzCalpumvoNkJVzbXVJDN
3+V53aNOsyT4Wk6erwlAtEM/Q1v1lhsiaEjqdeJThdre+9Ck3jTAl4L+iAkWppTU
GOM0WKkJ/8qafc5aGwr7Oe2LNVpWQiC6DResG/0xj5LVdzzjPzKppEJCFVx9VH9E
MvahTFU4E/QGq07Aq4LhJNRi0Y7bpno/8lh/QtV4Mlgu1KjAUKlqkhUJtn5f+F0F
1DTACFxL6R1mp4N+DEC9TBuKThhzghT4uNWykhBe7vlrtOB2M9LP1mqw40+Ax9uq
YQt4dYJ4BoWLRf2mqNlVDVYqkSsOnm3BPJp6aikLWy9tlLtEE0cYR2j2Nap23rJM
Xv/2W2XcD88qPuMwj/Y/NvJBppHS3tD876diPlFiptEcF6i6BgXwTvzB8xURrzKA
UrtzJGPFn/mhscHDu8u3bMFN1XP58YGV7lJ19vtwtDJDplzynf2sH2kvc24gTH7s
sh13mDLD5mfplY2rIBVuPv24W1ye0VXvZJaNm9JUDeOstcJduZlmZiGF/VDt0aSf
KDc3Vx8CnwvbtV0oSzdDT7NARWH9WVDIGfH0QaeXf7TWPu8Ujn74kng/bnuHa9qU
mVI+WaRib2RSL7QMC+ybE98A8ujFbYOb9whgc3Ko4zaqyFOEWPexcYIYK/sZmTaP
+QUnoLwsCfdcs9KNgeS6Wo1af7IJCcIbtRmmOjsdtrca55Sw7yqxCtCfMcEtUTb9
/dltbLasD4yClSLfLzTXATDsAZKqlXMH8zRT09+1vm1LFvBoaLdzdVVs2ciPPVzU
1eJa/e/Z8Y/bW9vgUWk88D53yhOrwGuJIONSVwTU8pyNQTLv8Q7rwN3a1Dzdt/ZH
Nhn8LB/6oA6NMG3EzLehIWsrJuGGJAO0H5oMdMxWk3UVomtvtsXf84UUxgQylvXq
EVgb0MAj5btE8FRHByJmZ4HKRUO23SmX6PWdSyiQGih4PKVOI0JKHfe6gD+cHno0
2RrJyJalTsBu6ZuHRTnE67Iuf9Pj1iNQY330jzKkWrsOKEPPnFGoBiRcrb1tqTF3
aKzaJX9dLix2Js7HLSN/DJjP2NERhF/nWwGYaUPBRLDEgj4C4yCDQSEJWKZsV69B
b1Cw/b9OuMGMuW8Gl10QZYiKmFPSqsSDEqBXo3aKjBDZBF+ynR+zV+r11LHzchUg
CyiOnC5ptsq/ebB1KDa+AZBZ3rV/dyK+DKBMB7GPE7LuDgB81x5tcOjHDwLSuqb3
IyNcCqp+XiuTNEP7DQ0a6+S9XJSkZOOYN1AdR0O0bBx9u2JCvyeuWcWzrK6hv2OL
YxLRovss6iU9uk+oRven3Q3EgoQ6OPEz6Dgixj9KNRC2Y7oV3zo+Cyu9fTBqKOJj
oUcod2S+zqPGjlQyIL9gb3QE5ixar6o2g/xj3bqcsuldGSHUeZhsyYzFw3sX2eTB
lmOmDozfJ3p0v+82KsITAyv3NxqOxU/qXM0BqILuxeK6x/JYrfAg2tJPIYCqt5Cg
tPm3CAoTxvSSlPBa9YgA1Db1EbA5R2Ky6Zl5MZjsBIejNYLfl3WeegZrUEczeXOs
UxNP+NVs64PMTEBlAtxvwjnVBr8sDJX9uNryfF1J7MPU5xmWdMb4rHYmEFp86rn4
GPqMkE/lftfNDPVhtHwlOiWol9sgPV8lIdx3MS6mMby668ISkFYrEwKXN30wIUCT
fYrgfwVvkO2ldnj9+zbMKoym1gAl9WzntXgB3KwURbsPoc+o8vSFkCKGmbUke7+4
Zl0oxxDfeXhV8sB4LYvLqkkF8qWc7/f+Q8JB6y4MnoyqGWFqVrCr9hCB1GuhEnU3
xcSmNnf9yfCugcUkzS6TCEoyyf0MGzoCDLRADAiWMr5KyrfrX3eQ+WN1P26VM8GB
QIX7iKRbj9Et1MbJkcepVlBY3/+/FWgQpFUjc9551bK3wfy8AMkThmGU024zXzHj
uGXMvnMJbJ/xXb38dGJxutZTftyoQmhMDy0BBYHhhPZlWngQNsdVAbV+EHJk2ID+
WzzVlboQT0VMMPRFe5tXttVj86fJB9QIsIwHIYYpKeANFnKNjcNdzsYUSNx+SILE
g181Vv/menlIszlwFCNSbN1fS6cy0TpxDdkJu6CBZZeIXhT0IF/K9catYK+c4qjj
yV1eEyaxyu4zgkdduTaF8o6I7TWlPtyE89LhTrehufvuNv9ZDOXnFVBbvWxnturn
VFvVjag6IDKyJDnRgxDZv6zl+oniKel4n+ZE+mBo0vo3/9HMxzO7N/JhRLE5QvV2
Ly1je/nJ/esnUzBxWSPC2XLt6FW0rWD2oRj0Ov+2UnXR+4uZjfGH4kDbx2M5OIV7
i6gCIIgySR0u8NeesJJjBg==
`pragma protect end_protected
