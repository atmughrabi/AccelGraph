// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KiG6apfrRUkORphGqCNoDuazv6QeabqdzIN8pHGkAhXt3eRH9ya9tBeWwraML5Gx
VBD1D+cVaac7fMHVCsYxCr0qkAC8FKkpu8kZZjWxM9YJWiglwSW94Io/6Giw0tuV
uK6Zh0sL6NfX3fH7ClWhLACIVwV5BICdtMz8y4aOfy0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7616)
UuWU8NpNxgsPrkP4cz5JZ9wlTbshvGFLVoHqGoEWjk/LyGBB9rM8cbiWGdCO423m
3snq/E7Z1XQCIkX7ghzfq9R1Ajf/Pu4auaYFS5301tCAe/q+8ynw36kHwht6YFHt
LKswS0hxdqaIZaqpR3cP88JLyOz+xqkSITS0PTvlX7wb8c6J88CswQ6OGu4SvFI2
Evash9pjrZPuzLsgrRp61HuWAezZLmtEh9EOgj7EPDABe0UeSDGoYY88qyFbv7Fo
9O8/xqXpfa9/NuWIZW1Qb6l5tXuxepj905EBudZZls0C0vDluSD89+czGIbp5Bvg
nWNd/sbhf2+cQJh6DpteIIHZAbQuH0ZJ/3O0DVPClG4cVjIagpJ3aShTPc7sJ6oc
1D/LOFPpbnb6w58HkoP7w1xFo2DS7bdJW0QUVJofIiwmsrUbPP0l3vAp8WS7zCjm
mOjRdGgzVYdpLgaPKYTqQ6IFIR7GR8knFgW2HfyiNoyz1W8fyXUF9NWr3i3vfyta
f+62omae0bvLaKDDlAoG4VAfKRsGrHbokHadZyZB/WWNZCq0viztjHJpw+bS5qmD
9KDnXy1sHAi2RiSXxhSvFJn2e01AvQU7sQhhFKV17f5uiwFJa+iE7eDeLF4Mte+s
qs8+kyAkGqjpM9lwn94MIca7LfxPJjS88KoClbEu96Lc9GNRmMs3v+q//dT0gZHI
41ZJAb9mqWv+Pj07B7igN0dsPaVtoU6myoANJfv+ZX4Xm7yVjiAiNETv4XpYg5Ra
9F2iE15jZ2Xj2RCm+xqxwVqCwiud+m66Z2AATVYS7vDa4h54c7hC0EdFvELlw3OF
PeK4mHUI7D8Id9WsdlH+CtEAt/cxf2omOR4RzMDf6WlTYnvjqwhrLdlCv6uPJnVK
agNvaYrmIr41+evMOVotIf77le2Z3LKdLtSOVNJTLLSbACqUO9WAwOMO7cf6TabJ
W8XSzVJMG3mUa7WzV7sYqM+F89KGFccX1fJyKwZbcATljxNOyTC3SVQOr/EIsRSY
wsbSkt26wjjfRCivZ4ug42EG8/4LVfFTTiIZsdkZw0B1x7USFOe7o8SKt34UZgp4
7O88gWJv9cWP/CjRbh7/2opzWVwgsYyHHGMzIDIo+BQDfnqcVwZfZ9F1POmgN2e/
e6Sux8RTP2FpNeOJCDpidJR7AZdaxZs1eILeDElqA+VNjNA1fNa3lKihFp+JX6FD
VRxOvVkAuqQ9HFgCsRBPivGCzF2fxPcNqWFrX4knZbTBI8nlhhGyQ+JFrHgWfVDd
5X2bp3qNa6VmwtlnTo/pxdETOT9mw3XMgPYADP5Cce0bj5DM+RGTX4qNclKlCbJ2
tY6TaEEK/DYe684Giw2lrmYpyD3UOGwefYaP/Tg1bTT/Vzze1lN2ppxKVVhDcUYy
3nownqcUo6wHlFI3e5g1OMN/RQNYyQw8/8mlBnpqh4mVj0Z10WxWnDBbUK2HRya1
VqLJw6MAniJ7Jlh2nONufCfNhy5UcpcxkDMKgxBBaRAH3iPQ/2WV2YZNFyG3J/AQ
CzVJQRmS/xP8Vd2kQkxPnsM9oQ/pHP/CVMPbKas/xC3yV48kKE8XaTDkG5aCJtqt
JlYtGdcKJJ78zTJfs0+ho6NSXE3ioku2C+yyGf4ixEjVWbCMb3ub2GvqtwafdbsC
npjTDY+IHEyT4BOUbD0vephl/LXhh1pDpzDDBvuZ+IWPgfvGzGnFYJjR6N13f0cE
ar4sSv7A/ELESg/sHfHLMGovbQjCCEWXAlJFi/JFG2+WMqFZq0x0/0iW4lHumSvj
vqGQ1usZ0OxIm8UwmsYSExlp0A8ifiUnH0O1ZkW8p3f+ASE0SSja3vCrNbxejnMI
Fn2uzMAd1Q8K4OGS0hB7kQZc9b9IUMYVsC5BZB9kgN6a5vn9mCQm8ar0u4lRIkWT
6/CbfRJjeHJ8U7P2u77AzKM7ZmiaBqhvdDFVesmWqWlu7s93nGiWk5q+eDayrJCa
WHzHBbZr4FnpC8VKYhJji4x7sWFdgcV9VtMC3/ZLNBiA9GzhsxKv8YLQC5p8ib/v
3VwReeCxbyDTyw+mY+Jlvlh4Bura19AWotA5NJqiZV+PZ+uQAGG7Xz1oJChqBstP
eqf2PYdr4yvOYk0NRjENDg2GUIpJ9+KSk03ldow9r/ptFsr5wOHYCyJ+ATB54zgO
LsRtCAWFW0bxWXPL0uyhbH0/6DYUOHMMi99d4q/AnHHmGc52pL6aqJiI8MIngqK8
7SZgFW95VT4sxfxGD1lic5nY16HP3ZBXSqwqm0NhT9p+ztjd3fo4fLLk1ORzVP5M
mtYrODg0vg1QB31zd7XnkRF267Q8qO4hftDMd8N7DYWoaF5jW4iDaE7WohUIVLPZ
hLl7O5tYxp+8M2a3NJOfLdTZeO3KfTp6vBEbEvi5pK40lMfcBiOTskVCxy57IvSV
MHrFwN1w0t1e7cxyb6RD2qm2dpi7NDle0u1+RwVpciH3Wq35SBH1hVS8EvXdI4Lp
xzpXdK7g/qxibqcnZd4E6iMSeZOXCAWkq/lPMzv1AYtfQC5lS3fUdfp63MLAUlx2
qbDOmNb0sz0q3jTKbBPU1dzSFEWwfTnBL5g6x0bLTDKBNYw2EiQi1onRt4j5e6ye
i4CibVwF/qUG7JBErBLO/b7+jgQj3i0ITVDCVqFpVhJcPxSE/D+L2Gm9epuhW+If
/1vyBy1JrgTvcfbHhXTaWP2GGJg3FeqcmEbiD8hL8uEJunyvBekv1KyJ9eEBvUkx
ZGYCu1fYn+hfkdvb+4lx2Tky7uY3xvFsS4ig/rqwxkQtP3oxuk+M/pegVSXOme7r
FmwfodFQ0w1pWoXsUwhtc61GV1+2mJRAgQNB/81WVALySLQQ6HyfxDc8nzr2C5AT
awap0kpUxgb4JV1SCFD1pCZ5llPZTOb1Vedf5PXJ/nZACsQ2CUXLhhD3UzOrKggw
yMmdZ8GNQMN/4O2lAgtJgrFCmbrnmrz2axwjdtMJIMTYgFMfG6Ivs8X4FaIs2ku1
xJk0dK3no9IJD4EUecWN1Zv23yImF2mWwbtI46UC3Iufr2yo3VG1VtEuxhukcGYk
620rdWfU6fB6a3PcmeWqY3XtBRqXQFY7sBbkJ/olmvA4+mtsGJzImRg4/Q3NYEKl
P/QV6oAiBR+sMAOihCO72t3o515ji+sJ3eaOLTVlaGLanoeWobAjJT2EnEo77R4Z
0TPOCxZf1wIl1nJNf36La408JUvJ6q2A2kBoDSo9z/83Rh2I273PD7ZpNyrBD7ZI
vh/CsgZRzbJ3qFm6cQNJYSc7DlYyYLrQacAPOPfxYmXHneZBxhyBRR9nKSnFQuk6
HBhqNFfNhIuPgVQfbDsMZlWiSzX9WMD1OpA0IpfAvvaT0P+S/u4FvI04w+10Pnnx
FsJRY5lGXhRNvFASsa/rtkP2Z3tizOKqsgq8rBHLL1Aj3twIprmBw+tISt4tO3fz
d/Cr6E5WzVtV3Aq7DDn7yWfHOk9LveT+JTevBkXpsX7aJtMRE1Qxrq2y0moyUoeH
pNiSRo3aalAQCXbM3xZu1yhzvVViuI/xOm0rPS3/KxW1tZJugWQB5YOpNzq3qLVl
ZAVTGoiBCSt5Gb6OGVXzCT+mR+9E7OflvqEctwKqdCwrsJTfoPR25wWjWb3dhs+i
1l/soJfsnQN4kTdRZnRyXoU7jbIMLA00xxmOYYTFUG8eNA7ybG/AN/JWHCkgUR+9
tZDA+kXDST8UcRto8QMZms8rEFi0D+PwB3iEk9d7OSpPgKFWfrZVvB/cLyUEXgVP
ZzWzHy5w5DjaCQriBqJaUpIpifcrFCXQsl9erL2iBVwVF0e4PfW8V2XMw+XJiqq/
AYtjy+21bIRh+mWsQ1OpBu8Guf8mdlEogGExZ9wcb7Ss4YTm3pKA64mwnn32T20S
Gu4J/Ivo7ItgSIDuoNcvws5jKTmb+R4eRCi6qQQgWufYjMeUKlF+UUYww5Gorg2+
/+dxcOsBPxWxoB+8mr/dPImkJ+R4+YrHeLrY6AESUCNrswmVUHR9tqi5logpoqRu
7Gh0CUYNSaEEUT+K89K0IKwTC4EPTTPSmt9DULvxjzjLvcyjQdC3fHiyOmZQKacd
oBYVuhDvPlx0oBJle7E+MTJmnTXp+FO4yIGMhkJ1pv0gyk8/UVh1wlbvoqMsSWLY
08aWEgFdnDbuhb3QNUUvPb+tDAgNvVcJinP6qL5Drie9se/t+yV+IJhva+L5sDl1
5ryEosMX1+p8eUtX07cZahO7qH14uRSJ3Z+mdo/LS0wDHtAwPN8Mrqisg6wv2MC9
5VW/d1KEIs6w1IynzoIrnxShhSAgYPato0jWl3W0KPdGU9msntPj+PruV3pBF9kC
9HpqandreOxH/wdnTHiThxsy+uf9snUQ7afaqx+zMdQbBCd+pcV6ARGJ3eDNnFJx
nWXcuyYly1B/0JYbd3WBamkQ4vOlyyc2p3k0xzNipvOFkw2YsuE83esMzKc0tcdP
WAnhK0DySJPhckfI/ri5qnCR5hlcaqvogu07h3tMgCnsyEm3bdRWWpU+m0IaKJIU
/xJDZZ5AMzCvgyS/OrTNsQ2/BPPAUSJoQrn9u/mAOZqKjd3m8DsBhAOdUy/5MZTJ
oLr6LK8mmK3P84PsuIZRu2XuTo0CDRNZtjX64K2pjlAVZJCermr6GZ7Sqbi/vl2D
O0HwaNZkB/cmlW1bi3FFeTzUsAmrEl2EUMhAZqqjcQeuqJL95TcpxTAK8sikXKDg
M2MEEY3GKZYrBAHjZAZkL6cJE+fcJ3I2Z+F/GOk9o0dVK9557dRlE30jpMxfSTxG
IKs/4/EZLvESd6PwZ6R27B7Hc6NtdLsOSuN4zWQ8hgWui56xxchKn/Xze2LCy36j
sRcWWcyOCvRfaTTbWhDKTIv1WMNBKiJZ3DFsC4LY1XC0TlosluzjCMd4bwtT9syu
dP2Tvz3LmYPASNAiqw1t+faOEqN5hJHQf8ZokZwaq/eWLUp0Xu8yIs9+oNGu7cn7
7EZ1EpfbatpF1cXZy2fSmNKa9DHJuhLLjIetScmRWga968azP89ZkY6K0YvdUGno
kPI5+LbgoWSgjQjJ3Gdm003nrNXqykcAAdMQEUfe3y3Twm9tpOQ5qMX2y22LHglu
UeoFud2hUlC4x53kk6VTlVeNWlVLwMoTMKbBEApJH1oPijDM+3ZEUCvdLPkgzqQk
aYfZ2tU221EOgFX+nUmvFU29uXxwL4x8aZ5ocOGYPRBD7wgL5LlA7LyaRKBzNeA2
mrGtOt2FrO+Iu88+vtvsBfo/Sxfy9M++DRybW0BVis5cpwm7GcYIOGWj8fqJl/f2
UgIjXbfdYzaHXwOLqkCnt2gJZxwd4zv0aZd7CkWo6Hhv5j20kJtV5MDwNrud5HAy
9SAGLNhSpn4zVfq6lRl2jy+ztkqdCLWRF5LRPzQvK2Toa5w1g0MqlW0slcWQmpQO
8vR6YcrVmGqJDlWHJe+hh1sE61kVBhlofHAhzpn6wlkGOKb/rZab0yZXswVTfmhO
sDpUAg5Fx2pqrX0DYntobIY/+ByQk3JxmVyXaSkNeZUGhA68i13Wb9oH+jl5A0Wp
shOAADr1EGnIKVnjA2BQoaOZTJP+CPXlHLKyWsHLA2i1IYEO0Jaz245+zK6ZjtJo
pZslwUQl2QVkOvoGdUhoWxO6wwTjRQNGwo+vAYy5t9hkUgy9Df9snz4YgQ7et0SI
zy0NkFEvgzmKmZedJ6Ln6Zq6V0Rg0yWGHprBRf+RNAlS6X3OJpPWyAWhMRBz3Iwl
XhUepN9PIWDQA67dVOVGWIF3bK2SvKG/VO60DficMa/IV8aJYu3oXmWJ3oa80mAo
E+1dMZAsuDPgr3K9WVQ2/nw5iF6YMDFegS5HgqTGAFEA20g5Z3dW5HDrFfB2athf
sBs1b6T0b2T2gosmmUl2U/Qa0siHkSDYTWOr/4wWpyaWasaUqO63PhFniDtrMU1i
UjmO14jVDY9FADnhnfgNXJogCsWbp1A+nVSNxW61/r4gy31TZ9HkQTZq+u2GwXC6
6sXBfKOduKIAMxsOMo6vw9DTGxvVQDdbSf8hIewGPlyY+aiBL9k3IXSJJUxCnZon
ViStmyOu1RfBFjv8MgfZdTPetx63aIavMGiDCWubBNbOTpf5vVPU9KZVGc354525
2IpApZLLKql/Gi+Xn5SrAMAA9NjUAacDNyDdbdxMqcg35oSfc/34bTrbwRj68dMK
1VvkOmeVpphnNwApeifrKgQ+XWg3cPXjhI2a1BHEa/nNp05AO1ZXB0p1KURIzEc8
tQjv8d7cPpxtC9qxD23sdf0e0wcrJzp4e8WyNlAlEJ31GUL21hxr2wMWtdlOgBlh
iDwG49B3vnXsOhlcwuAb9Rg/Ur6xZ9BB/wEgiAi+njcwTGeVO9yWAlEJ8npfgam/
QY31F6V3Y16Rq14do3ExRzevdMDs5f/GUnbvMMqDnQVL0uGLgOjiMS2e3IvnfUSA
Fes8LDKHgBtIPVMl/xGxen9AJ/c1NbcixW3/vM/Fs1Wtq3iau8kF0+u4vHvGiDYO
p3JV761NjBWEmmmlPb0I7Jy62qKM7FSvxwydWPH4cNQ51WSrCH00jTbqNVvhlnvw
VLPIyQQgnIocri/kuart/ciFZLUAi026KaxxjW2AmTS/REqfna3uDiaYVG5beiNT
LwowR8QDY4WJXkZogd+5xPIaoQAVGxV4QC2EGCutEJcLmUyXftpa+RKZ3Uu7lCHy
z3T/845cIEfvgU4riW2HKwd6Ue+Y/elApu2Qz8t1xoNzVXaUesBqbaJ7wCpIku4d
iLRt+h3arUgPCxIzv05UXfwjvIK/WNvbq4KvHfuOO9gAYehvP/kDQdhkJHUK55JT
s2nUk7SiQ5MCA7O2L10i4ugFd1bbdZJajndSldyTqRhlyvWyCldGECUi12+BPglp
ypVQta6eMZ+a5poV3p0uOszqKupqbBdvQeru5BWnmMCMnl3ImNbcdYWG/Gbi6P5Y
uhIPV4PCPfehr58d0cpl/7IfLTWVOEt37BMmUl4o3P5sYXdejy0D6FPcYTOLMjB1
CfXprGvl4GqkP+Va/joYDBtEHTRKxSE7txEmeaf0gj6zSGWwAVfpOaERujtPAK2f
8mPweuqbI26LMswaZaYFbVXwl9TpoL8KxT8o+cI3c2hnRk02L3hSWPN2p3iHEXaB
QT3AtMmUOdjCiDsaaqaEhxqthnA0+2JORrMjd+lkQQ1mtI69cXVLaNl8pGkSLrT6
CPYZBqtTOVRUonqwNbEzk4wPJCjobDYfLvjXy68LTqBYhdEqjNCVqe0pfNjkp5uy
0LsVrM18OYJ/5rusL/DKlgd4NQpeZ2StqPELViL2/oe4lnpTOpcHQ0bApUyQexH7
VugmBoCuxFa+yUUacJEdhMUpbcK8mp2t1AXs4FCBXMsynyXYmH1CxWFE67i/ayDO
Rmt4doqEaJRTfIN/25es0cP9bppQPbmn3vGBNkSWLF6k5h4ALoP2Zxw1wP85kXUr
Md1Lgxi/Dzece0HvhYgWt+MPKIC4auzcBVMF9UD69cPWzK09G+PbJagsOZobtLV1
tBl4bM4jY4UvZ5XFT+GtKbBv0Wofhq0GrxDKFDcXiFqAL99O4VP3wfOav5FeLazs
7n/BAVLq/XoAD7IwCC/r7PeWBidMNyKqjz+0VAAhdoVkHeBt4tj/aiacdiuOnize
k2VIpki/CdAnTMEQ8Lv4L0XNWUBrEPGfKA5LkWIw8SSOZh5fVf+kSyw8mbXh5vlC
RdQbgY8EoAE48EJQf+VjdO8jy6te8gghvW35ZC4X8ejUw4YL+40vZqd2BYdGKXWY
GTLj32NmUl4oguMZwu2mY12bm2n4iByWWKmKQp1mhrWy5852C8X9XEF7EcAAr6rM
MJ9OW/ldY/XAb6xb9gM39uR9wFHwy80DE/TYLIBE/4/6bxyWmIGhwEqHrDGOCt7c
cP252apcL0FPfoomTox6Q+289zvF6oykjldRD3EUQKAlfF2UClWUqCaQGDxnv5ON
mlonAlVrYZ/IePsI0GXMFZX+P6DDY78JoxHP4s81bq3YLgBTUZ0YdmyqDq8ne1R6
ypSgzfHrklxpC9ekUZHrErzwChF67+z8CQgQuYcqeN07fdzi3eupokcyu9Jo324s
CCMLLQvOV0V98IjefITAe3OMAXLIs//cfLWGmfMMBt0LjPSXiG+GULPB7uU46+MN
rvCzJNO7Gi6zURGOXpcRK2k4W84bi+l/IcaqwNyI3BLYs98RRCrehkzIvWqhOiYt
vsMUi533jxU31ihPwuH38lXS0su1YI0Nzf14nU5EYMPKsgAx5L++3gTchyVKbpWu
48hMskL4h8pCdLbRT3bQm69Rgdn2S8aTCqlJ7pdxtjTUb4gWzGOe9o8YHhuJyR5h
d6jncpu4Nz5kEj+RRjtbu8NLRgGM8H9q9SROaTSfmB2JJUiKrLkvH1dZ2epZLpc/
477nNr7+5ENTZQPIP8rD3lT2NKYxwaBn3AekiZ7i07N/wz6Zlx2OOiambCbTX8Xk
f0OVZxRZtN54OoLb+UEZLbIb7cdi4r9GkH/Boojpe0yNM8/1Gf291V/vqUIMQuME
dT3nGOCx7OKwBTOLpwxJCGAj9RDT5f4pGXGP6Vp66afqsN/UFh+HR4U4Lsjcf1vR
sEftgEotzcvniQMv8AR26g8VR6j6F7yjBSUARXHuxANGkDYQmGgUgFyfn6HBOpKO
t9IR9kl4YT0IpmJqqFTvB9lvzvkGJdImdgFaKBOa+fIpEVlcnnTI9Qabgv4PSYUx
gWsXjsdtRL9pvvEnrtNVz5CderPB0karl3bebnxxm86tU1wfVAeVfMU01vTcQ6T3
Cyxi1iU3985vQOkdN8fI08zjisdMb2OMUSOR+W6W/PB3qieWztrIiqwY9FRlWRR/
ztpAiIdCpLVpaMz7GLFkXGxkdCtLxdtEg2QTin18OLF2CJTwPXXP1PAy8lbuWHqu
MT172oM0v99YKkxbWwTHW5Muyjo1Obwbv1PrXMze5gNNJSf8rXaobCryIpNJpydg
4sxwJO3n+uD/injRHITZAp+yUHDKAdkS5aYZy20XP9HKTqyjxHygsa3Fp9gB5cFx
a+9w6TR9xSFJQVIQ0edQpesbogLt9S9eR1XXBQVZjgyPtVkqAwBV/STxEu52Bezy
MTAgW5BVdg1xdF7gBS8pv/eM88nz1wWucRu6Ai84WfxILnVf5xqzNYWiAKdsyicB
T8cwiPVBMm2kEX+J1XuGQsxTyszBmzg9jzRDMxbNS+FueTJsk3ER3gM/IymTO8nk
lrKrRHYk2FcQ5QYCptOFIVuRPpFeitG8whP5MyMnzXTfs20irJ1lwd08HAy/+vaY
qtkFJh4HYnlcZ0wYtc9+gj/cq6uQz59o2B/ChretKHp2r11fu/BXFtuLCWUOZdFl
7L5GYPFpoUppzS1+RbmfSMLz3r7yISeAEFHjDTLo8BxlTuR2gwwChsaCwT+Q8sqn
aedUB5lRfj5P/hON7gNaqvq0Vja1DtXl8Hwb/aFhppbEYj3mcXkyrnxS6cClKUGP
zZx3j64zQBbRMnkn4Am13sa1RxjapbmJW3+OKagqbbynzwRlPwukb531KEPKCkU7
whTX3/2ycI9EoHlUk75y2KlONBzz5D79c3YFBKMoH6dGHS4rE3Fxwj1PK1aFhkzn
MvQo6Bp5x995NGXELCc6cMJKKLCXPNw/EvU0wKNs+KAn1iTQP17NUGLFdumaQycd
L1dYi+1s5lNKjcA9d6A8/KPTlL+7ZGzkHPOrkyVDtMOI6WAIwxdm1iawiNiAt56l
1nahOSn82gDKPZn4TNU44VqO1T9BBcgVICFy1oTS1AMLT2GL75jxZaV1WJSwLN4f
pE1slwasko0/TxE9dWdR9BUUffE6ZKmabT4hxLKVxpqRjD8rjDoCCbxWCQMvKJP2
oyMcXuXLkDTOJdzgft7tRso1Zx6MRjvxcSm2COeYFuauPWOaBuvkvpxVzIh0fDsp
UhLV7gRcnA2SngYgG3obS2qz4sk9t1Yo1qwWFbhrs6KKus8/gy9LJdx8zRadOUSv
MWi1FLBC20YZP13AuV5JScnDmxQK3bR7PxNWFwxrY5ReeTghwZ9EC6T65LyGk1mf
1tv6xYaFVTRUuoCkYKlsFuUQZ+w1WMpj+V9Oamtosqw=
`pragma protect end_protected
