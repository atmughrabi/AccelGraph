// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZoyFNb6RAyUAeIiJlHamek1YBoSgX4+jKtEovhBKLFRrWeVDDHzM7RBhRgYsxf4J
7ht1stVZTgdyO9q1+PvCr/aFPpM3gItvb5W42H7+zkIMj+BoqkcvQN5YZ0M7UdFm
3iKdxe+AzO9GCR0IdgwLaBGUJit9WLDlwRoi7vdvJDw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2304)
UTk2I5NeveYZV54am4Cnbwo42RltZ14QTijY3cSUEnVtvNYAHVjV2hHLAyW8xO58
AVADRvLW1vwbGV4FxMCLOF21NVr1Jq696hrtl1ZiNfJDFDpNBQbA/yNseib9+k5n
IhT+LwvGbFw+3dEQye2tyqH/rPgh2xN/AbUdoiEKrogaRDkSbkFNHKcvQzt+XBSu
7UqgJz87w1Ak7ZdqDwjXl2AyzQKnPA/TS0e0rzQFPpO05dJlCI/vQSTIx8yud1wN
Nk9QVH9g9HBDbRGXAAWB/rf9sGy6rRjsV/KdxiEMez7gRISRAFi8EaQ+fWi9oCBu
cYwy0NOj0iblC+pHFdA0Z1wnT/xSNdZmsp7Mksl/4mRBZUCI3G/nSYdA7tE7fHew
I389ZxtU7fXHJ3eNESCH2mbINCSmpBARzSb5OiSyraRCwoEYXxCGvK4sEFjB2UKE
OlmYPhsk/zKY6DSHQ0hhRnySTKzhY9J3UM+C5AfZ7orgj+bj/Z1t7/UGofLv5Czt
4PmLfrVAYwOHcHzqXQIW1YdCwUdux0xLwon3GzZUbfzDpp2Aaexd7RWY9tFk4YPO
uQow8TofkEWgyBjDkk2EM0umtSscsCBzwhYs3Vj+kt9D1BCTbEslpLjgTuo4uDN2
PubQWR8ssVwLhUDJTakEURH0dCIq0dcDJGxlp1PmurljD8uiq+vgnym9KlXOkx+M
/i3M/vVhVAn++4SqtBSbHkxszMI12iNG8e/k44LAunw79KBkquUCLJxBpz3qt7/t
0XZWcKyrY5Npg7wTz+8l8RTichTgff3AB3Gpr69xCGRiJmwROTRYem3x5ZWiiwnA
pQKCT8eCuRKYeoL4nHx6ySkIgawijM2oIwdFxCH7Xzp7H1gPzfOdrZIRXmjHB9Bl
Fx1FngOfPEFqEXMoNScc9/rkuoXxhglCWF6BnroeZtzahad9Bdi8rQNA0cQt7Oxp
KhqSkjIIxbns1TYHS1FKAhZkfy6uWf/Q6uf4pfOfASV0pTROESzEtxfDOFKI51V1
GItCLkJVeUY3kdc83RQ6J3pQ7D3grZ/8SD+osWEAAxvH408CzsQGz+Zn+dW4xpDY
ELX0pooyF8Rnp61jha42OK5HS+UYtS56+bjlr6JmgEkk7+PFWo3ZfAsncQlgbH80
1qp6vHMARqz0tGCsNKJS0jtWjCopab0f4ThL6J8o2uU3R/nLPx3sh2Lpdfl6+tNA
CFnm9SLo0kQbPPooKAtoUSV/IJr+a/OTiPAW19DWxnJtdcYh4WoC6jsBS8uBXWfi
AfW1KFPqeslnFBpapVsKKr0NT+NYheerFREbZH6w2UZlo3nGoVPwx37X7jCtR/1v
yV+rolGU4/TbgPx0+NOW68BVAU0Lb2n6Ro4C8sCHpC3tPs6wGuN+UQRfASL3nXpi
we3v7gAnjeI7Ogz/gqkjf0f2j9RxSJQ4L7Zl3+Q/Cf50xp9yscPrxT6LbRonjPSg
bgsWkVsKMEEWbGTXG1MAYhUYIMnvNpEBY91CFvJ4X7xa/ucgRT9dT0va3Lu+r2QI
5v8ejl8qluPEgB5FpLGa8rdPUdLZDzFKINAMv+2Y19rGvc02BauXzK4HohGbESKQ
PwIbgfiRa0M9Q/dk64bU4qm5pVzdjPmHR1Tz3xaIqN+k4evQu8soAY9S8SzJGjZ1
x2gWy8Lgr0uVXWmtbA43Ke7qKMfBjQon3BJ3s/dIUcQVNmABI5uOF70nxXMHFgIV
kPFDQLirrsvY6ufkMWfQQPuJlb31IuOtYn40g4GRFywn1E0VJgdosuBPawgFqgE2
VM3Wjzy57qrGbPirlKCxNyl3NrTZaI2He/rCQLx14P5nckdzaBKbkogRmJufMfjF
yo/uevHPwYoD+NALI4g2+HIflc4HK03KF9ScVnGv8wALf17Y1wVij4NRYHPNqdF+
K/veIBrkvncnqiiyR+8xjSGFkNyGgv8wA9NS5b6jdG0y1Q/EtiA5ddjVJNEIz28z
jwq1WC00YHeDDup0Wgt5q4SdNcmM0cpAmP2Z5xla+kQRWHzTCMy33gJjyE29kM79
J+ZdcWSUFcJMD1Tkie0kI6rRRTeL3un4LYqiu0W4i/Y+lplE2iNa1ZmhKMGQokbn
XXBpHKvpKe8lDxemu6dD5MBPbEEuRdFUIgfWqSSjp19I2CThHRK2SKnq6wIe7ajF
HYw6gOPiMqvFSNbYMg4OVWrJY9+VvBIL/M4LxYEbTCpvWld9NPBOoyNaQ01i2mHH
9URM0Qgpb8lTSJfbrLJc1TaO9fFzFMo7KGy/W6kIk1OW5H1eYuxW/o7jHPrNVPeS
1bwNfXwb7Kkv1Pg5FUDbXhEVD0vP4dAe0yApxy6NXEiYlcSH7ghyTRDSFxYC1FSm
BBCcAkP3mW3tsodT73l0xOeKSYc3UugT+prvcjQ/OZ3EwkjRkv10FptdwlkB9j+m
VDFOrjWNWn9b9rVLqeFa3DyXZMTrS9fa+OlZIahHcVj+oWqFu7o482xxOHfOiJST
oQs6nzm8o2auBzh07iqpxjNs8yIPTdfWsiICcIxpJoJJ2Aqc4dDlzrxto7a2kEYj
UoPjPcBqNIjealP2e7QghysVMoKVJZQnVYS4KfE/YjdFKLDqHrlaUd2cd1jDbAJi
icznQlLaehYqkqhC6WlkZtXKvNc+M7E+QTJ05vT2GTKSmHnR70FF+a/4BVnvPddr
ZEeefza2UECbLdohGJgDXIbVu/oO9e2Q3D08UctTuIzX3lfrDiU+QnhcdoFo9+ON
tom3n23fDTT6qqKC6eirjOKK7sX2wXUhShJJCIFF1HROy0N9ytZgyTZoiZFYhF48
0qQce7ZOTuKFnWsgzIH1cV2cILTmpOhuwi/1Q8aK7317c+jsFec2FZJRlVy883zw
P4DjKHwcBL0j03ReSu10DJ5VJ26xIaVKwwQRW4LVel6YlJjIfSSw0jno66z5zeo6
SlIFbmhYPw8EwUZM09M5r64anrLxwqh7488Dx+Brv1Og1vIwihVov1aGC1wsuWdo
XGBnRNvaf/zq2XNT5yeXHeOxoRHn70D2cpwm+O4TDi9IeMRp4NfBPNCd84bLmksn
`pragma protect end_protected
