// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mW5qelVXVD/dZAU81m5XQImQyHVXBA/pIvGP+hMJsSAIIsSmTVZIXysoX9Y+lQSa
nq2Q/eKduB5Js2l8Wc9uASnYEUy8BsK9srQUDPdeJ1rXAh0O9yGQK/uWbQgivyit
aZRormsyY7dHL7dNnH0B/jgRflGripdbt2eJxIrH4uE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4112)
5iYdh1HBRoIohvg7wh+esMzVM0e/J1mc1f+TpJxKSAAKeD6Ez7yw1H90EYEb/U7z
4d9PcYBHvvFkBDV9gyQlG8CUxiGJGYenuWXx5jXfXFnsz7Gf0F+FrY+Hjod2rTZ5
6Rn0p95k21bcIvGfRBsEzxndHyLLegP+TLezhtbowgJHJ80hMFbekTFe2Totpdyl
W97NzuAkKgLwyY1BrjmtqVEgoIZtbjj8wmAvPvxhWFp4cGe6R3YlCFyj91fxqkrk
gNid/O1mWKEq/TdTaM1+pDvl/KcAhb386FGGreLDJvZ0wDkebBaE7uxxDaVjn2MA
+MnJ8OH8rn0aAmI2eHpme7TMZre9EFhoFAVLGABHTIsuNodL+zdYIIT5CqWB8AWr
bolu0MrHepSN5Y4oESAsR3K/b+4h/OCAqL2ANc/OlWaUIQ8ebYIv1JV90LbLDYaY
5k/7dN4oTQdHZzNGV38n8ztKjoOULwzhf1dxzcpblvBgVzttizN7U040IwCXsl0i
SOT3b2bRLAa4v2JI7wfaqMyHZToBsAN3oLjI4qa4/hLJBDp//2R+nQkD7hoVH6Z8
+m6apduuvLyxi3/9RloCwUi3/1WbOiutvQFe7+P/SrxgY7LVoEJqwUVtbfoF/BG0
dHvQbu5P8dmgSV+8IKcjCf7OVorpzMNubl7KDvbZ+29+QgqTMsckc3XPCfCU7sVU
K8wCsblM5GHpdg6fGkq7ie27lFRBCSag+YaQjInyAkEXfV3E/6qpOSF2UjYX+tr4
unVOUAaP/riB44SlXlLE+8HcTWC/Hoy6g8z9GljFRJL0we0fw7Q+t35+QpExC49a
NwYAGj2DDYyghK2oXr3hHRaF55mLi5e0IZ07jwhk/9zZBmQk8RFSH4Tug7hscZpi
O7Sk939dY6YmV8NXK9Erd4QBF4ftboq044DoU3FtQ8FCjzxNgDMB5eOC2GPNBnsb
vLQ7+07QgoiQgXNAqBaBfkN/m+02bmQTOlWALL1GiMpkPY5rx70vU/n9/r1e2wMB
GNBdhR5KaAE49A5+vOPdrbWp6tZ0iWWIKIISSs+XGhm+iA95F+K6fKMLP24CLQES
TlgL9NhkbKDyWfM9B3nKn4bN1gFu3bEy0DOAWaeTAqepoX1HFNmo8SdQMJzM/NmC
qRQmX4D93xBlYlBx1Ir1/fW4qr/YVeDfPp9anORmO3HBZtawlXNczECge2ofDzW2
pLMBBdyMK9tyVP9eKxAqjeltmCaqGH/SOxVdBS83u1zal7IIbjOMMxEvW/gAwX9R
H7DPHKbGunnWWemv5dmnD5NFUmF+Ge/OelcrBa88NQh0YsWfB2VLU+EC4uSSji16
pixjdTawLmcmxe/zwjCLyfEBN1Z7cGi3GuIlzGs4SxeB5jnPpavCvGo+55JL4FBN
HoEgypVMytMhRFlyAQgpNOqwrEhd8v8znsge+ByDvoDZ4iYdr4KLuzNM3shYXJCA
V+1vjbYKpaEoa8MvhXsJ9HY0/f7Ndsd3gpomWgMBxv+Xy7A6eCsNJZ8YKtLok7oh
g1beLsyh3ZFJ/UKHmsZdnDOQXijMkXwz+dPTMXtLOFOzeN46EWzRm0/SKzwTXgfU
VrciD3iRJ4CHchc72XdPZUfpVYzzo9tRrEdM0Iy3e+mXjev35aKxwD6EE/Lcl4ju
KgJhCJg+OiiUZv1tUgJ6bqlQgoGbptmLWK9fpZB9OY5vOtkji1oPtW6lYuRrUgrX
jf+dxLmXLdvyzmxlfhBObjrFO6nDryOrtMCDPqcysVwI6fK1HuDj9sF5r0ibqSNJ
H4AhfuL7jSoWuYmlgY4UBAK+WJ+cPf46U5SY6hDHXwFPcQnepuYHf7c3Hccu5PIQ
jHI1UycH4gxl8v5mNIVVge+2LAOG8+DfVHBJpywQFCmn1H6O76Xt9MWoMywkzVof
xVYYfFc1a6jvIRYDoiFnHPHvcPfIb1qS9/vQg6YnJbhSAawx19DwlQyMSzJwF0/G
4doD2w8gYoUnsvjexyyz9Q6gFm5eDgpbrj80b7Zvkj4ljOspiF0HxbJreN0p7Urc
PDhpPo6nwIbKQBmSHIYi4E99uEtycvttIwm+9HOHJyuKT4vDxlepg8o7UFhqj9Xs
FEIUFh3OqsoYqS596snNAXv9FhHRInficri16Y4WScmcKhhLauP60RGoJrYx8eGw
cXiTCcHvNozw/u+HzMsM1DtX4Quy+L+ADXw7cqaTGsW5+0luajX7QunJpj6Na4r0
YndhZ9B60D1IqaH5i2ukp+LkSKJ08PuvoT2kCYf9AfmracCj7a6mIgxwnbHp29wl
ZqthNZoXMtWBu/+kMdiJDpyyxlc4UTZJxQdzrnyom2jQM4KztbxfLTqbczcU1lpQ
yMAREbJAwIqFa2c9yZVETQx3SoQTWk/a/gJOVTXDuk8rsMZRlRcYjoe/lTXYlEoW
CoXAxC2gHFqv8/gQXz48eIP36ZA3yuGuXIQoWsn0d9so9xtQgBltc7jCcJ99MqE8
b8fTl42tSLao2/7NY+uk0FOQT6/gi0+zNQ01TpLPY74z2ra7Uks9cdMEDNjsMSXt
BXtvY5UKl3iIeEfwhrE23TnUvOa0kX4ksa5GGu4PAawELpfquiqh3SqWhTxSw0ch
STTaWveSG8MDzyAmOYeyYdKPZiEU1TtkTwT/G9KvaA1jBYM2vDSjykHoInx+APOY
sZYidjGXoQhaQrJ1l9Nh1gFHvrAiWzMjOO6/8KYMQLuzCbS15qEcA8mB1rB9/F1G
2SDlf97NBhXTIF5zHJL5RdNOMsPYIW4UpyZDgdP3kgK93pXDlCu+Cl9sZZ8lqXLz
7CITo+Wnb0fIRDFO7s51BwIui9hEmGlX+U+JTa0sTFJlkfqoGOnXIQJpwJhfAdPs
6oYFXzZmCdlEYyMUSQOH+05eDSlUYyVJ0N0/qzuzzrItKBKQsnWnjgjv8p/4vQZB
/Yh2rXguz/jo0GqjAp/c6kAyEOCzImAv0NpOpnBEuYCZXEpl43JWC6j5gTVIFZ+f
KY6OBCkfUYJPgzsoHe1bFq41zknoNdP6YY2LCePEqgDjbDjrMCMmv1kKw5rV2J17
It49pNlB0q4s04Oic0v2p++jcQF1DQr9oXyyHXDd4NGp0NCTO8cJOq0j0pUHZzYQ
AiBKYMCr8blNPTiTHrEjOucjUaRt3MOTUNpZhBDf4uLJ7aXmKibCQcaVpEq54dJq
83UNnGw4pwDRBXyT7icpmoTuOnhu1WBXI0ivhwNWJSRYqFp1/pOjg4/AV+2eYQwB
b8od1yWDbnMye2nA9g2UYz2gyrdO/c7TC6mDZvyznIm2NdvvCAVDL0VVbw8q3hlY
0/nORUEFnJ8R4Ua7yJ3XKbdW+MuT8PPWYEmUeqXtCcbR8wX0bfiaUN/OZI9iiEOQ
+R04T819r8rnaZsfBOdLZAIf9/E03wzBlhcuQeYmWbX9tQ5haS1C72Fjfz1FOhe9
Q+uoUYkSkjU90kKm5ilCbNHSljV7EdKTehsQXN1rJbenUSWSFYCwXaRz5Rt6Ld2T
ly5zlUx+Dx3t2ZT7HtEw4Kv5OXyrmONiAQ1czSqG0iEsYFyci0gn2WNUwQ2FGMfR
55YIgbW/oqNmovLmM/x1kt0uzkN9eQXBbXFYKJKQaWiWu44JU7JyWDWccUkNtG2R
yz7idyYffWqwFChrnIrdPfdYQxiCQID1VYBgBZC1ucj9VPgXJvHb9/LFB/YhQWWe
hH4ugSME9ZYjcpee/LGWfKDjUpXwF9FMRkEsueC5To/UjuonKmNT0uDlMfOYpFaD
C+j3oc6hbhjW/lcR509ZDqVpllCrxMUN37fRfTZmrBWcmYWbry9cevIDSeZMzUPa
O+6qyzbN8WRAjTVol2QP8lVqlGp9XqRYVm7dL1DXdKgUkf6jko6OJpu4zXhSmg5r
rguRAkfqX+sh6XXxVf5iEHCu1OzRsN1T3Lvx5J+AF+cYUWyAG1cNnTgyynwAva/V
hLRJ2dI+mIEpcY9syT1jbvVQp3ThZoboEppfEyx2Y4fvCVqasbTq3SxNPzjy6JJO
ZvjR1BI5REf4fjdjzsrCcxZP024RbtOTZmtUT8cW7a80UrI1lwOHrBiS8aRUg1sO
2bcB3KLywQJhf69k6dgF90muniVfPrz0ws+/vvTFLjAe/yVJ7XpWCHkt+PkZ201j
C38hm2Z5iZYLDSVMZ3rtYTJWgys+0xbcV0Yo9wZIEtCG9hV4fLwnk0XbtkolZvGP
IoAlhOuySOhJnWgLSDWszyZSgaOU98lR0Nf8iJnWpGqxU2Z+hw1bK+fZThTxap0u
wSXQbDDBFsuG2HjPEzN4/SDAbM+OEsy0YLyKlrHhejXGvChwZ2mxCS36jiEE6pmV
MRfmWoN7/qaVW8VN98ix7CP4T2t1z+WhzqOILEozoI0oHhDBEiNbEeuauE1HLfX/
EUaYveS4Ako07Xd74UWgS8dTnfSrEBtAoQAOAr7zKQq7JuNfU1oHlQ3fkYXeM2wN
t9AwM+ZB9OjWgzHHzGFOvpqAM9/vRFn7iP2FUmxWNVUF3g3VsWVeZXejBAyTAGjK
MhseXrZQ7nJ+9DUZguOEn8sq5oN4iuYG1bhLPFFceoeABghOI/nkyTeSt+ZWyYDa
pGEZDppYRmR4QGzv5r3HShy/5LRZAjjJIjKyduAEzZSsn4m+rW5WdfCp7tLAwP77
703Yd4HSQa9qCFdsXsidvnncEjDpHX2FTpLJaQFowzbZoH79cbVMYp65/RzpRAql
hIM8vOAwO92Aa4glyDslMzW3d7cNrX70Xq/U0yVabYDlO3268dbuAGvlkBMm+pjN
gQezXeGwnw49/YzFC8rLx7hIbjJDfNue61VVA8Og4luU0rFAzUsoid+s+SD9nMGC
JtKChPwzSjKG4bzo3qc8L1xafyCkZEt57bhBE94dO8AX6mRvMl1ad8yLbzgRZncp
j7K3qM2PeXpb+R8vfpJzn7hUPQCaDdFDlpmlHbd+abO5HhDxp9UmSqQcMzlSHk3d
NcvKX191PPpjY2nov0LF2YOd2zYHLiNCg14/3JrdhFJQSl9uDQo2JAG1mgTNWjOD
CHOjHHJzLeEHl2U0IUF6X5E7uv/dAJ09C9PYkI7ZZCgfmAJmMr7GSe1DlAiAl7oV
xvKUV7OtXE+rDjr/o6mQm4HD9Fm65gsfEyVw0Fich3XcFTR2AhikQfg8hoE/c0KZ
8oVhYt/fbxEc8G6vWpU7h9y8e9QXvQ4Wn4t0RSH1VcStMRN9tvmVwvXo/o+GbAly
lPAC2R3C+AuuqbPy9w5XPz6jYzrFiMvs/U76Fuwb+P6AlfqP8wAAvQu8mc3iqLO6
/WbOTey7V8pQq10IyNEOd01BgdNquDW0ZPkNcoxNymdR2cLAzRYcFQlEcuKrnaRn
UtKsWOJEFx5HBsa6O2rLBt12ucebxu2WyX8YFAfjrCpoKRPmqumqiGHUHINU014f
WarGfcJNZNMCshpc/W2f1FaotbfPXH1bj9WlfmbILSA=
`pragma protect end_protected
