// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bopRFJUVbSuQp0ITAmNGAPGrHcIqnqh8YOe6hSLB4tqVV7Ddpz+gNZ21i2IqY318
pwxseWwTXT9frcapYW9QlZXihHND9PbLe0lEKQ/FK71G0SbL+r+Qu3JLC5GlRFGt
2FFsL9C25C1e2v9Do9Uu71s+XsxJKqjMq8OaKTH9lbI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15472)
OUkdZ8sLDjFDlL61v8/akhchjRon/t9RI9NL55AWgjC1NeLFoCiuNs4rIL/679w0
Sa6C9kbFZIW6sTczpzGbjQjb4YweDbGjZ93ZfxvvxXGh8tJ+3V9fybPfIe+Y4xNn
fv133FKCN23diWtZWw3HhY0OPybU9yEL03xC5km6h+rJiCNvXQuHZ9OlZRy9lv8W
TscvuBgV2y/zHT620O9yU4zuJXjc8e53EJScqBxEIaLK8+MeZkr/FAOmd3w0p3vB
mxol8mHo3NGJbH5bKvFJkTeBoQ1mAssifdBpRCB6u8jyccg3gmDk7VVssu+wfpwy
w7o4omNYtEpez679VGTWsP9FgldQWy4p2NJNurviDiIiRsjXkEKylkBEDVg+afNL
WWKav9mPX59x2qC6kfJIBOFQIfO1jM2/d5oIBf2IeEEXY05VnKui+GvgCsZ/WarD
kO6x2+EtjNd6+EqRoyDLl0RjJTVMaNm9XcCuYIf42P+Hz0dYB0hmHOmPGVuo96yk
bEJDuIb9j0QrMkuP7wGk4n8QE3CX3yAcDnLbiqwsdQA0spk96yHQQsGA/9K5SuVm
90Qmg4UdVLLPhGuFOKyoDlXJevlL/jccP6vpvWNrEu+IJ/4nnse3eW0hB/Y8y0xS
3ng/ULx5bNP4Wc9APlLOD4bVaqzGhms8m+fec4tfFJ4jr6BjWU2ReQEbH/ZRHsRV
PBoP5F+su0MCWrHjtHC47icXIBfOTiVY4qXnkqj/xu7H2J71Vnv05zV50sGfDK/q
wDrIKh1AmpjR8BBcVQnUb1XgwCPQBDhK/WkICgcnb2/r5VlVk9yN6lhByDO4nRC5
1oK9P99QUQ/MsnTPtDH9hTYYlsqXlzihSCrxoRoV3t87nApNJPdFRVpcsyUQbi7J
0ds+8FtdRa5AXYtTGgv0J9DHgDpe7SnrVAMUrwyLAZ90Ss1/hUHTLcFgGVcbohkJ
KfhWtr5GzVb/SELaYzqB7zyp7AjVinOOfyXxRG44bc/FRNVQXB+GDoXqcJHE+cpB
gdZe3KpCO2AQRYzu76N2JJxqEuMAbeUuA2ZYNxu42aaz7qSrf3FqSXd1ezR6HwL5
vrSFXHTzhZLo9IKBLF03f6eTSVvbS9FjG17WdoDyESUCziyBfpaFeezcuQ06PdrM
ShKefy2O0dPSXmAx46FRy1sdMGdC0wKm+1yQPymOCfEWnsXQ3BIjAHFQco5Twmqf
cchegE3UlLXpwwzu6l2WxmcdMV4c5hQML91MUAUmiM2dHfPhoJqDfUORZOnhs4l1
4XurqY1x9K1bkTJ79PODf16jVMUkE6S1ZU5QsNNQkvLTGUM5W5n9oxNjjbaaWbSD
id+vJkA82oEoPhLJ7e+1DpO5D59xzM8MaVUhahd7b/K9zwoM/vA0RDWX9xfftl5J
0zNmvYZ1af3LDLpQ/PAY4fHZL3HiOJZ8jh/NeJIBZvsQgYz/xKfqmE3FKji3uG35
f/1ewg1+ZI5HAbj7EtrmorSnNpJkcTY5y7Z+zEWIO5Zq8hj17eUdddAQCdu+CnGc
XBr/PPH0ONTTtQTKNJ9KTiidaVSbnx6ljJHwDFv72VmeQJ2ARf+MlkI1tO4c2/CV
uycKcvc1veB3dtfvhGAU7v2ZPxvDAjApcBCsdOEpAfiDuXntd+PAhD+kErwXlALD
9Oal/yvwfJZQN08nsQVpzn4O6u7Gf2IPya9tXINX0/LMBzE8VKbSiB7wQUQfuArP
8Z/LONuP5p/Y9ysYrVLbdM3eY71lbVMDjY0h5066Bmz04tdbsfaAjv3ukoOfQ4L7
T28dKY9X4GXp/Hcy3HHw5ijBXT/lnFOWMKb6gG83BhSJH01jZd2Kc2Z169fvjv7F
JSn0NFTnMk6PS4WGo9JROaqWL2WcS3qQ6VWnxoTcirb14l4VjfslqIA3DrQG+lU9
4yMDsmYR0eEdAxNWA1g+j+LnWGZDM4j4MjBGRsk816nMVdZefzOi/ncLgVThsPYK
gqozDC0oom4S2iLftvhjtUaBBNthJNW+Ev2evMez3wQ5pJcWzyYDPB3MSgSkQ6gQ
Ph6vFGX2lpDRGwc5GRII/R4BlBA401VBDLRATfjUgNfzhM9by/khY/WAqTwUYSYc
5hLQKCEpTE8PzSY6J+xn0RPNRdLsPtDGKOoQ5/fSmHWMyoB8zRuHX2QxoaXMCkaT
l5mDnIogdfcn1SEqzdk8cYPDsxvVDWWLGMYF1z/8eVBm0hH9RblBSxLXNgPhGZ26
aj4jo8Q/ziPAK9yKXn5LftSsk4Ougvn/7fkO/Awj3HatT4Yh9VOnKxFDf3NPcBAD
ABdMeJGLXZgy0t351zK+kgH9dOcqrhcjM/P3E56OtoiB0z0pQfFjiyzONFDDRfgQ
zUEidt2TDvjIv6vrF1ASmMyx2+ZNCpdzPKhHfzc4wWr7noNpHo/gZcY+qZbteWAr
FWEYyLAtuu0E8ALKMWJupqltJ0bGgg4a06gj/4KyVLk+tTs4cMA248JGLWoUTD/E
qGHElEhYEcxI3MDzLBEVCI6AYjOAtgvxGdrRTkyJI8NL7MNvkwnJVxWrfvhSSFTb
92uXcRbOpt5VGn2lv+12vyrxSWvMR+Vdg7ZKFEbQOvGfm/SpBegv06qZdrHrVNZ1
byd4l7wC8n6hYcM5v2UTSMCrYSu5Jx/BDhBgSfT5BEcWJlS3I9vdF7V8Of+tNkJW
EdIVSv6EMQ5y1lWP4SlTDH+hbF9TjfG1i10vcUfVcOhwdMoRPoWt/z09V6WSMAKA
G1GsQHDNftL5wfdLtjG3f8CcckuWWnZA3W6bcEZJzERuG4Y1GYVVhTxnTYw3oYTb
31KNKvCRJqr2zfZOkDNiL3V/aQeYEh9Q0CJuixjmdCxymJl15kNtmvov5asZmYGn
JC5QwXPk2jgRWY8BoSvX1X+CRgozc8qWcuKN9GsYCWFrTn9psuvpkvAiaR5A28G4
yg/o84nVs8LS2XjLQjcjObER0jCxpxk6hpJIia+BJra9BkGtBRIjKZIdqe42mzQP
U2B7CxSni+qOi+Bx+UcMCMEI9FGckvB0/jbA2RrOcXm4CAX2jDQq9xGLwK+N3nWo
+CVs3VKld2a1C3eZINVb/LAD8hmfpwCg+8fBVsm47UejXm7TTkvnWAgtoLSs4Yb4
W+fjDx4HUp0hvOu0dpf+4A6GVojva0G1pNMkzci9DjtCpw9aThdlaziBdhTE3NNL
OOCEXW+PH6uZMmWllJHCMTOEcRBxVfruJKNmZV8MghYrf2tX1myL3aWFrf+J3Rpx
H4+zYqY5/C2aS0B18H0/vb5I7ChZsowlsuleQWL/KOqIZSDBLRTiK4SP7yK8xmLU
XaIvq/H96JRtFFX2sTCB9VVbLIdxaEVVhrG3JLKQ8JOz8TEDi5nQQZ6ldUG1dxb1
qqoTQdk6NEKD/L68q6rBc95ycl4sKlO3GIKanlk3Ep/vFDkjVlgn4pJuZ5InbVW9
f0EpNwXw1ZYG0oicb8IctTFVnHiHOy+x2vrFIR35TthyV/pYSCj9FN1rGQKIV/6A
pSKjq6cQlZGgkzmqCbmguIlR/8bJXiv+n9iJlctgRcTKCuwzPmbPj3oUv1Xs66+Q
M0md7DTiXVAUq2te4+V8DeHz4qSFFXDbLwWHJjT3bMEXZHNofLUxym8jZXzoOeet
nAno9ZGNkNHmzNgGNKqgoZXOTp/0fD8nAsmAAr/9RqOJIFwY1wsAGrLZFVla4p3E
OyUyOr2l8S92YumNlnAijIyNNVnHN/nyvMQS5T8FPdUDH2tBDTNsRP/ZKvgAw+Pm
ABVIcxOBbhoi3x89zdKhuO5Z01F4//LV2pjntmu8HsJ49ocADuG0Ge5VqNLDNaZT
45uLeGCvdjHVyH8Jsb4cq17sUkCDGQ4wXvfys9j11fwM4nD+fyszOPlgbg9HqQMy
IcgbnO+MR2Z/eEpApDstc1h8BjALOAY3UGF/GvmKiB5AL++Dpe91zFPp0y4nOq4Y
9cDENrb+SH7/I7rkN5ThAL1TPeaG16hqflRJ6I2r26nKkGjZTzzySSCNAvSsLT4s
xAwVztKaMCeq8OB9ZJu485L3dcAC5ivqoioG7BN1wIcE/RK0ZK26nIk44avqwYEQ
bbvvN/ppyJzFJTVRxq+4fX4BaV4pz2qR8ie9A6e3tGmEpKOgHTj5p5v4SU6eygvv
RXogrgC/mWAmDXhLLjv7KxFVu8HVZs8yK38eIWCSepUOECb0W0MIjCmWEchx7ios
aqgG1gNeVLyi669Ui2gfuJSsW8/snCp6sozJ8r8oibWXmQbBgyFLJvS68NRxA3Y1
LJTRP3PoCvyPmpKo5WMsROjiFh92ppwtnsrf6qigMzcQ9kdPsIKjAx6pymir/P+1
Ng1P65qzl+1g3PHzptXPLNgEv9vT03qdwQPeJLAau8vNahFDWgLdG6NKemYHI+SJ
ZQlJyitaIx7pKYFTyFHI9ggzzQB21oKbRNWAMw86XoVvZ0ZoYLzRyqhsPuVqOq/e
a6eQSSaEuE4ZOR3QcZTVAuuRhcUoOpphU6pieTE2F8LvVLCoOYfxnE2kzQaFx+oi
SMgNDDv4ekK5RG88WEEE8Dh4LjeEjfXoWZTue/p9ylFxkI1ZplNEqX2s4c3NHesW
l4BmX0rSCqRkEOKfgfHipb1i6HblzwnlxOp+q8Qir7ypNSohtVy66SHY8/b1xs9t
8cepJxd7WUluKc69cSRZzlBPT+6wyv98dpcQwpKdy8vz6S2xwcmEKQCx/8/yOp73
vUeC8/wahbFOUFmrCgJ2nnGpQ+yhLxg/Kcadd9UzS3jXVln02YhUs2qZPUcH7mWl
WnBQFwCergbjlYWuafM8dM85OQ5vo6w2SCuiGRqyHhMln79tUeo+HlNoMz3n3Hp2
1HmFEyOxyr2WReYyUA7rgDITdqXkWego+LWCgEilp2fdy9EDsaKE/x9w8illqEv1
/wB0ZDGZpYn1qsZUGMy0ynLXphjl7zbsIGiY+OoMmKYVNvob9W6HLUCTwOYAf02I
yEinhJj2JJFUTJYZpwVAky9vZ5ReLWm95m16oTxE3ahthN9130BAhnVkIL1qJKzE
k2mfY5jvMQZyoSwT2yIfyTqtdjra8CYKqPtnkkdqpIRIXqA3sEdZkUSX605izLUm
y1AFPGuzFEiVPwoSi0GXpaGrqQt334H+RQK11C42ZxW5FZ/ZFRKy+/ftSB8xJCb5
LGFLYVlNCtLgDQlYxDJfm8fWVTqJOplTFargpwaZhmbz+j6bMB8zBWAPmAnxXrAv
shg383ujAZ+O+QxYDebiFQVe3yfIEKlY8gN42Kyzb/ARraZrVj4+lfikJMtIzCQ8
gmmmixbJpuGZknoXkLncmII2xefM4ye2bntT0/8075cM+C1twI4tno1ohi0Ikzt3
l95BiAuBxPLXb54XRrjp9M4BU4KXA5cU3mVxK0c8AVq8uFwjK35BbkrmsQrhvNb7
BhcyMfO7GEf5HmXea+ZYkDSYgjiUXPkKAFjGM+LQChhh9KzaU2TZVRcNMwsXwKcJ
5GclhaS8ClK2LmCZJuJdKDLn5Reku4ZyI5SVqYLzHl1mT/t3pMM/psTcRoOcsnP0
hBXXPsVUNyQ7UDVKR7XgGezwbT0yFbgXGPHQftKU6zKc4+ePbklBUOtn9ZqQEKe/
ODA5ejWqatSqK4HpMB2Aa0cpkuctiHihHfrfwcmCvp08F/l0dAaQV9RY2iv2l/4w
xLoHxtfUE2nAWQngB/Yy2cJEJAvkDrOP+B48vgS8NIrCmuK3Ab/1MD3J6kOifHxY
vTkEFTjoscvefRRVQqCUkXkVcSXeiUEWZI5MEt3Ox3eopLaqc+hBHYp1TuSRmUmE
At79bRpXrevvQIv09RB2ITDkEkU+d2fHbfCzmJVjyKKubhJuWYH+qTvYDv1rQk7s
qIzCXpaN0zhFmYksHovpy6+SsH7p6N/2gHAyas49aYjo+gpWeX2aGNoQPuos/3tF
UenwN2qajhKjgqBmogU4By4/4LQ6aVQjrww+mir9W0dcVHgp+IczoUqbhhG2VOrq
aH8g5iemmiJtjeR391QZ53G1IlwWDrm2Xk57h/kn8fh70JGGRaACA5fEJ3WNWtUi
JAvTvQlIkOU6/ZOmlI4Y+hZSDVptnc3Hog2Uk53SYZJDXnVR+CyZJW/L2pkyEAe6
ycUsJ++dNMmcOooAUCpLWi9j59t4S6hCTyiR/EfT687Z8HBEs599KqxbHYFKedas
vga17wQREpSHF+JvquTm+tTmXK2jduyuJvx2cVEB7XRtUm0coxL182XJ/8IvVSUJ
1O2ykjo917ckGq68w9dpiC4ETAVObs7bqbM44KvM+PbPG3aKEAjxIyGKCAWpHQBD
urlmYXd365C2qUe7IKcinqO0L3s/8kqfn17RIGeTn8AzT6iVXQwZRhoEfziZvgT5
vt9PnblGr+PQjdlZyrsLAMigqhG3FGsDbd7xir/bpxSbVcysBQxxnXofwO/4dJVn
IByhrDASAGO7y/XMBh1CnP8TSCLZ0SU1eypRXtwG59HuVbfJgH87RkUHjQun5ex5
Ymv3+W8pZK0bbX4fWP7uLarfxyGjXnW8Zwk9T14bCDGa6Hv4FqCTNHeIMoc06inN
CifexrjQdDpJEWnPNOXCTejKJVqcG3o44t4WFJaAxixPVI++GHVqfsJU2oXDBGjR
+LizSVslLJnnFzCqBJ71E4G46Q5JBt1X178OK4uUIkdw54r6VUwhtRWdmvqdEokY
GXYargiW82VipFBu1PqmX46YXHb6oGiYNf6OO+6+m1zY9rMKf3SxZm6JRjMuKnXd
DJcBNVB+36BxdCoeS/k9/XS7/kKK0GQ226+qTSZgptzie/x5kSHv38hTm/9JfVx9
vfsz1wEUjz6g3EaR/wuCRjGovOt4Cjj3LENXXH4ai4Ka2C+70dZ4kgDHtAzIuGqO
hPzdngE0nRUjhfLmBjd6P1MoDdhzOfaBCsXNpEGo3f4szWogs8/uRhsPvOVGLr8S
eULFlvnjpxmbReNYj61Qyd5SCnkS3yV5AcjxECHCT7tgUsptAtetEEUP2vn4p/pO
c9gxA8a/lraefvdBNl+cYn8cMJ79qXPo7vN9K7wnk5V8gG6XGAQdfbl8/YLgDIvF
ehcvKW/rXDYuC7L81M8ZnKzs/U8WS3/pXAOZaihCN9SIFwRKZEkZd/Tm5DajUSZC
gqGf6eAzyqLQlunOqz1+fMUxrPyfW+8C8sFFhyx0kTv/FrijYvo7fwvFhwni1ce+
UNHF2D48543dyc+MeSUx0EQpK94MWLAB7RNmc0dRJQ9XHMC3jVqgFtw6usdipgL0
U/ey7AVBh5Ge7DOayE2xRYt8zjeZFvNeoWdSC+r68NAoKZswfAp3ucfw6o20REYK
+1lfRPfV0yw2N4Dm3srUOp0yIito5JGiZpRsrjop8VVVYedCAjU5ifoy3r5VzyuO
bD0q/Ph5GLCRPfdMBIrIUWbsb98vLHPqO6GskSLrbhA9CP3sK0bxUHKCUAihl4Dm
r9rGGV5lJbGoACCHehVz6ah9knfOLxX8YLYyoKYrAS4bRAMNAikK+UlH+FAfcx2s
wTnBWoGC5eHwPStb8mGp2Y2HmddPDDp6pOAe42hzmPTi14+mfP5tMWBW9r9WROBo
eLEjbWNhiQJOI+pUlplBnbbEtCD7F2FMh+hbzE3nKiUY3qpVX8dpU7ECjrPEP5sz
0XFGrqWTXR8dDHCFUdPksU/8BFEp23Jewjj82kvuiKHeHYFzaLvWrm5sBwJnaTnW
YAXP/WijNgJQgbtFeWOZ+w9AEKTPk8WXf8ew2eouvIbZjlspiRHy2L35a/No4bOB
cR7/hk8au9ldOWI6r/cxQlIjaQmrEsJ3KW8OSsz4WvNTJjNMyF8Dr//s1kt51Vu0
6qt8Yk/A2IHpL+XQlQX+4VP6h3xRlDtdDCiDFygSZ++3/7ihx43yDSKVRAXz2aVN
O2fVXvBtrrI5D/UkqStnwgt4gI19k1d88RHGSUhKommQAiA0eo0KWBxU/qf8MR7n
EzD/HN4YU8NlkLdAwA8viARv+dIspWLD4IKq6z0XzhTlTKHCCKM3RbMfwm2Rb2h8
YKKWpVJFALLXQQF6W5C+3cHFhDnlFeHndIVarGM4YsTnEnSlnYcyq+BZiLUw3dIk
CU7pVPspeoD/qtApU7sF/UT8C5uuyPSGLI2esUlHgA7jDKjU0/rda8yxGVW34Zi7
DA85C+OHa3PFyW7sR0D8o/3TPOotEsv88cuO6r5R73llA+J+9nHuB9uWdd2WmQYT
YBDi37c2yI+6sMy1TaUgDlRgswbI6KlQTNT6Q1M60Z1ZROzgyHoRNvZ4IuuoawOv
iKmqzNut6M9ZFnRPnpjTM2tCPCraLvlHrBFI7M+SMRfnZFpaWUVMSGvX3cCAxFav
5JaZtoM7zjndIZYeOJPpZ2UoabAQEkbTbNDSXoLNLGW9P2s3rDXENF6sqYBFtyVl
6y7Hhm5DAVltOJgae+IlUvW2aD6WGcAj7RStLvJwhIEniQJExK1EQkmVknmtBQe7
pTFprnsMGDF38h9BuzEbbFug3UTH0gaVRIigd3fqNDh8EQR2L+Jtv+8EBSaISBjz
NhvShl1ZBqaU3QLa0VGPQHWIissN8ZNOAL0nQetJxBSdu+Pha3DpCYX/DQRcuSUN
6hSbykUTuU79m5S2n41kXh2aAMb7gpVvqBzIYB9Fkw5W1bKE4nSPDBbCyIZVmBcx
vuiPTPx0PMRG/ZUurn1PdWbrMFYLGDLO8PKxuWzSQupwhr+x3FjbUI41RmpUzhJe
GaFk+O8A2CMUk55nCsCt4v+8ioMVZ17aT73ldNzPsgWG2B2fwrw7qMay2VtfVSDA
IwkOB5D4jn2Eqen1yPAyYa1el9Y8eBGdRkn9FbZoOpKQ2rHzk/K51cgqr+jziC2N
fAq8gXRNBuGO3iijXKQWfyjXr1Wa2T1sBPG6KwZkysRy7YHDwcsMAhlraLMF7q6+
bsLoEr6wsYtRBRq9sR+to/7pIlgkOWJj+2v/zscXbGw7hnobe9dPXyIxX0bsTvn6
3FiffAvd+K4ehP+d77Br7gYV3y71CFU8YXAK3bWBBT7++qUMU1EbllmxwkCPVton
awMWSa+GaIf66eet+HwPkO82LaSk4+zaI5iUb9CdXtdXCgvZhWBKPH8JqhVWywpj
sNZTsvByeSU0cD0kg5YjQE/NhTIsVi2EGoVnyzlX1iE5GAzHC1BLjzD737DrPxFV
wf9GwZ84vbaQh2Ij5Jygc/2gLyIpTcZOO6L9j2acJIzJROFPryfD4BiVlqoNdW15
lWBnDK8un4lwJouWd/jqk6HcQ/ZpugVCI02zI2rxu6Uce628/g+jgh2lGzcukgNw
0nYS0kOzAmRZ1FkqKb+7/YhSRMkw2U9MZtTVZp1tFaIbMMnWqcVnt8ZJCWwE9o5m
kuB0u4GDMfZJ6+2P5OiMngiFcxyWqlxfNCi8M/91NsaiAu8qZafNIIm6I/dKFBg1
ffHfSL6ZAXKQFNXvwPqfNO7j3pIAfELPpOOJ6AnCb/qWgymK1QhmBWpQiBJplixd
rleJgxj5tfS7hvGjbNxa3fA+DQZ+MXjeM08kuYcRJCBQ3mX/SZffpKewgSYBWIiO
fARZTpDN2zFsMNDD2VYbXKxPE9xiSbd4oWDYCRblMIx51+h853oLQrelhAxs2JJP
y95lmzdTSXNNR4wg5DDK6ETj2fFYglMPhICLueZwJZ4B5m8sYFO6f7ihOcERcdY/
+Ofhg3R+R19BEOzmqbNUu1vl28Qs6gomVQW9wThkWgdoDHz84yQo4cGmJH2MXMfq
ANd+2iXUjBI9gnqpUIIKeQjCbFeU5d0xqUbRRW8rV5QX+SKOWRah83WlFa/9lTCy
uQJsowsl6i63ovzobY9b8S6TTQRsB7rWZJh2mDAaMCY2USR8gjtLP3KHwValGyJ/
zLvYhj9mHdFlgdpQZCwgawcUZc1yWLz3nJAPzrSv0dbXtmdqKnjc2rXNZRkCw9tc
o8r3Li9XYv6nN5wa1Mb0GV7A6s3HmMn7HNJ1BKJXLOHaWw3oJtXtrhWxaInrEsT3
kILfZqdM+50EiKtYZYwGUhLC7nEujjWJFB8CQLXHYTwZNasknfX1hL+9PpmhZRUu
MQyRAfpN90JYf8TEtV+vTS9blrqdmeo2vZYOZH6orCuzIY69ZpmU90L6Xg61vCyX
vDeLgGMjbF+WQNgt6yqKN2SYaIgG1zONKlM6A5Ap+0cjIGAnZYNMoG8sminoZxo6
9QDkEcZFUepJ/ELu9ZjYPC4IaOVzhBAEejNM3n0OSqRI4zMlrws+DeMyu1suapTa
ELcQqhNRJd2v0yagkmGTr5pf8249YG5cQ8b8qRBcB998yiGA9UlHXu1JLDr/YTne
uc3FCZ3PoSiPTWfoWLKnS/GlcbNW3m2gAqxtwY/ABHaD2igK3HI/qx3appwA/GOU
impfmPY9iXDTz3Ej1il8r9Mqo5PGto+CbTFDfMDkpjdvs3ifAyTvUNVjlk95HtRx
D3NhK7SDV9Zc8bayU1mee0Ss1Vp1Pr8gxc/Ta/jZRiBgCHLwUHzLPULp/BR7X5Ef
7Yu6ceyaW81xDkQrWmkHuPCbOMxEz1U7e0TSrvv/+S9Ye1DrZk1XQt151S7XrIt1
rBJ5QzGj0wtg2Kh3JKUPL71pfMl2zOhCfH4y8NIFKKTXmyT8qIe8G5P6wHyyUXLt
UUcye0j1OcbAZaIJFr24kxSAt0ELfTKrQ2WhKm/e9dH1ExhfwNbKILgY1DQmitnE
u6SvfrwUmCVb/H29T9Nf2zsD4ObdMyWhI0C/7X7ALV1/Fj3DdeSqibE7lgXonTVR
NgSF6Q2j1Fki38CVnCxUIMSC+d0fs87iMcxzorHk3Ivit6yMiU3sln/cojuY7rhP
qh4o4Z/Tt9oPtUJ3wAzQcHjZuEthGLOZQk+Bj97/K/fI0k5aDQ4ZNwUYBIS092AI
uiDCu5MLsIrI630233TYtpNjehBWmo+dGfMuk2ZlrZbl1VhpxkvTXneLi8zA8+Dg
eh0QmowpdZOBozvKl0yuRgm20H05YWiSbnSE7F38/5BUWYMBuDreS3p+arozjr/C
NgIEvi4/UDFlGbvqca+zhb/ZTyPoQVLvjCPFNFJEr3AIi/LeXb51K1Ef9d/zcn/c
Z50U+dAIztpbDBdG+FgOQ9Idb3ahsyBrL+NUMdTcdNw2oyUdznI6L4MLOuZDSC+X
8lkAEc3/SPLv4iTsJMjg0Bvr4vGsSjqFq9pYQrE/JEVwAzZVMS90cdatZFnFyvvc
vZMNexUSbEsJx21xLtxVqjMwALaXU8wAXnTJHiRll6q8OZR0sktjTxywTScmhuTk
kqfYZ7ABhG+s7W/q/h53S4OH/zxj0pFBJoxwIUmXOcfM74w+yxygOonVQq7U9TCQ
qa0EZV7eyjiqviwuHexuem/lGugZmveF/UTbN3WZpcvVV8hkQ5ytysV6jNLgdSI+
l0broYY3sWDt/XTPOc4AODf/lSezvwpKHFF1BRgRwZ3TfXGWjRqa/SfMMksW95k0
9gpUoNBg7gH9cuE3n9Fq2qVQC/PAzsu88byOYftf//2u1F/7gm24kxEzu8qKLIYm
WI4lQHUpwWyyTosyosxzO+40V2mumTjE/y3oenfJZoyak0Ogo/4Ryi3cnBgc9dDP
BSHyQkq5b+dcEtQl6bvcvByIJwQWkbb98H3hIA6eH+3Z/fa4kuG0bXDctBOmQQnd
GN2bCZz62Pzrg5Z9IjlrlQVDSb+NsftgGIazgvMT+tAe//ofQZJ1FxX1gWrgrK1m
/iOqW76iMQsVqJr7yIQW9mItpns0zbwPlY2vy58PFs1HTx9btKkgh29r/oxWxSlF
KLasFkYILWmTOm55FQ50yijski7/gFVJoTSKZ/TVwhHWJzJ8ShrwSjYINvLNrKxA
zr3WBaMToDcuhsG6stT50OvykoSmBYFBOmoYjzwDJ/vlzS5zwGj5W6Vo2nLv3wm7
pqGnbEoHIyUm+Of9zvbMstjfOw/FTd4bsQK1KGtBJomcuSaDeSwO8BZRjAEgtx3D
2iugHsSqjXCkf2QKO31012SJe7Vp3aI4WL0mjqKYMI3EhWbaYQf8wV+IJB/rKmDL
9+xyLCC+Z/MALU9zEjYS3kTK5qcWPshySdmZu9JsKXB+AQHoLGPdqQ3lixF3fLEy
EQ5EO7R7VTq1lALh/jewvbtUIvtOJvVavD5PDiQLltWtgNZ0Wbf4DZiDrd/yRKiP
A3LnJZyhXyvuMjeb3hj+uCQcivVcwU47cJcIyYe0Vm+4XV5DIherTPHy/ltuJsWG
Ehp4Bd/TTf89VKSV/OH+3uywTCyRjZ3teyZzXBVo9S8340wmlv6RGeQClcYqA+EN
vCkwQYH+RZK701GHhIxho2MDU6OauH86fc5/oxKkfdeIrIUQtB+Cig+gxLNiiSjq
sTF6304Lx+vkiWgCo8/HmgGkJ7Nu4lW3tYhjSfT8f1Ik6feC7lmMMrzpjkglWUBY
f3Bks98pUgxwXBKtZDMHpN/V5g1xy3z0XHQejD3lxjbX3Jjsi8fRso/oKD49tGPG
3a3ADg7n+rw6GsiivETDnbeFTQVmj7u2l+zlGDSag4hjIE3Xs/ECsjWm0qBkQDHA
/4RinFJ/sqI8lhXmmCtt0UCCBydYaTnvx9a0toXKp5Og/YA8uhqRcx5N5umJeWsB
IjnARCdPj/jvK7/nlI6+gS2iWy211tCnTqhfQvDsIYa9CSxZocpd1HgBgNmhwuxr
nFBeWXO9I2m2U3MDcpO+MsJiqC8QJzH9Vwzo9XqSX59os8pyDgdsgGkKL9fKh9mK
L/MuXYFsgnukhpIVCm16nau5fRwddAbDwk21AQcuEyu9uxXC2789CTJX8v9rYAgA
ZxcLTVKjLsdjimxratLGQcO/W6p0ipMMquL/uGjhfySic0Iic/ZlHBi5i8BkUI04
iv45fzA+tnw50Y8aH2Iwsok0m2jzJk1J4q7IN0Vci3y0YFl2WrMW0YkCRTfSH9hW
eXK9K0IJbKt/IvLoArKOw175NZomY3VCJKtRagk9/itJxxzsj1mV3C8dWBx7Ra+u
Z3rW3pHg0nTIwFZmmPy4WSzpDP89592ifHIPNmj0/JXoUXMId6hmaQnZ7/EXVy7C
PnQY5m/UuxqsnBO7Ni5uW2X00sASxH+O0rlZhVdBEJBLy/GiOToBgtaij/wIjouv
qOXuGK1mzaZjOWNVdEPHYIU+KMh9FK4Twi3/qWPkMQjamUxTFZi9vfT1fak6vTg5
df2L5934fQ7jWkZd9xb/JqP1KdAyLkt62or44Ifq84vrIN9K6i+++XS1eoqduj/A
UjZNWpIPWL8PXWY1I2zVR0hjbN1exL3kYlav8alXgEP/KrLeWq6XVvFes9fhT5Lk
ZcjlVF8qMxFY0RBwb/s6+KAmi+jAzE5touiPdOUIp3YF9aK9n/GkQgxBenuGyg++
2tsZLU8bKe2Hmny22FWv0RdwN/vlD1Pp+PCyHcrp8mziEmFyfpRGQjPD20OUqZMG
5qUyPIHZhnjVlwHuRki5B4511Lai9BG36htK+dhETliE4izDWwXVr63UF6yFbhrm
4rkOCCIXdWda9lANbdg2gwFr9X0M6SwETIprU3EEdYL4HdN2RnW1DQbyMyRAupop
WG/Cu4UQuzq/aTHZUMdo9s7F82pH/OmGsjCLHs93wBzE+Ecq9RdLwiVvpBug3BqL
EBtoyFQxGFTp/KyHbnwLWf/w6OherYDhPpYldchF3BrU4eynNRIMYD/4zbVKLoRx
UQ/qbHxGCCg7dWornl5gCbhwzrInOcHSg+IvS5eETjvtWIJC1oUFL8FmsnM8XvIw
S5Eoxfn8aYd8sL65WabQFIeIeMb+y51+Jwyj4W9qhpG31XqVLomJcy7O5JG/Y5v3
Ta/CiFmMgVtlYLrCssT61avTeryOr+XKn+HDsFJKAC/QMybrEZmxRBUY9a1g6N+l
7Wn+mxMgkr1pr2xGT/qzjKuEwNvzQQBIkQRyRnLqLn1b35KR2cgHQOSfnNCiPgA6
8ba10LIHwTmdmRdV3QpSx0ufmpQRddTjAtBE7juJSWZb46PMCEQ7+dDJymMMN9Sf
zg/oFsCugukxGaErTHFH9KRgpMBKjMB0D7WsB8oBjeTr0q2tUsB+llzuO4PvJhrg
OYD4bbc31Bruxd61F8hDsz/XgOIUM51iFqfUgBlPjRjEeX6QRg3ooKKgJjnEPzAH
MoDhm177zPKuMjDJQnRpyNJuMP6RBlFSF6hXDVz6wwDbHOVEkaeE5OCBN7TIOPH6
ae5XN82v0U2RLTms/dSJk+LUSDDViWOiAhCj2Z/4m9So6CurYLH9bONax0ghyJzp
Usk5tWOQqHXhsZmxBV614ADorgWHV0hrLMbZoLE/hxkp1um/cRi11SbLxONbKGqe
0noDfYD76v0XwapljFUoPW/xeeSBs5CTLWnrJE2r5QrZzy1RO7FhfJiyLYsXpOt3
/sAsxr6xnzbPGeT3oO3jja6Qnve6yjQilZmsLZ9JNdU13RDvL2lGt6dyXoUUG/WV
IBr7VwvWkCZy1UYDhNPS/1MJvMSLGHKMnAS2LPEDCbACS2FYRndF0u5PfT9mUso2
fXK0w7dIwJfjmU2oEP1TokMMJGVoYkQaOPzgbA18me51nTOEpuje88tInO/aq83S
aXSL0oNUIl1ICwrfwacV1kiSMDSw+4t5NJog0Ez3mmmnjMipdm7iI1ZoojyxsLBO
QDc8cquZQK53sN43n5ikrBZ9heCRZIGpdUeeFT+18bOLjdYRSz8joQZ4MVd77EUX
2067EoUN+dYGHLl3VsNAlYQcxZYtbNaSP+aFI2evtRb4hKs2I4YKlwB9Vr+9+E01
4m32O4/GRCXmigpe04bg8++FD6iAC/IKlw53wXYcXUpz5PmQLFBGXOjGHaa6NOrB
abAKmDzZnoaTJ3Jk6A7s7Hrz3GStONLfxPhac+cjS+TlDDMt04+WjWFnFLcOORmq
WIIIBUQqrccHcXMBm038dlpZHsDZ2tdkgdq7/n79dJ+rZnGo29FdrTdeFj0Pjbvf
YIh1phdwNhAOjrkjJHzEXN6mvI2ILn9kXs0p3LgpyKku8G/sxjMCVrMClJG3AM5R
xLqviI/pijZ0DDPRF0SQZ1bjZCzCXvK3FzqWmxM5JGmMb7wLWXBmhH/fAawm4nzk
ZUCZqBMvWCqoo+8cMyJkyj9V0N9Aljhnqar9LFdMoDhSTO/GIBRkPg5agpNeLPHZ
yGVF/61Q/sHAWKxqcRq3saNpaUooZ5KYW6eoytUu8FQRneTWT82KO3SVeSwp9LW1
UoX5EfF5kdURlQ5ffX3wsSy3p3dkrLpy0adLpsN7FRLqaPlunUbMwSHapLSNGtEq
f8TXH2BK8swYPD7jGwnCy8Kj5v8O5qzBrAaMAi9mIWlcQH358yi2ZFPfuMjyeK51
S8efy7/Rg5ZiYA1bsb+6fZ8VRwtmsmgJHB+LypggBtkK8aeaWGNOt3CZDxkOuLxu
CKc9l11Qh4h3kF87iC403/6sthKgy5fS8wPHTMNcyGx6UmZ9rLUrwx9DcX0WyjRp
r4X6ZIrX4BcXNJ4ek1zZzd2q2cAO5Ao+n3vouj2ORj+rw6bkJhMdkMp+D9UQBk8k
1q7AaAhVhPOlIlWyHGXbQGnRztN8PTr9FWg5+kUV7CM19uyBpnk6WU4psLZRuYd9
lYKiT0uxyq/OObW8uO/qZDh5gYQzHJepX8omA34kBUciqItit3eTinw+9k0miVMU
KCSdmQSGko/Hzxp0gZdc1/D/i7lqkEOlY+jhcvG/u0F497qsBkuJAZy8MpH7SBgL
I6cr+7WVk94FeUScMG29wwJx2BR2udRG0g43XmenJrz3ZEwiPYPg7fmXMwvYF27U
/5r+XTudofl7KPjQE5XXY5w4bAO+rZ3PGj81kD4Jh3M0q4vxry7/Wkpmk/+d1X9w
tpQIdmexEJ9HFegqF44Qt3Q0KIrUWIylHfX5yAg3tK3VnQwzHJNoEZxgvKdBgPYU
ilDRQUAigzsuDzm+mKjYk+/5kQjD1n+kH3m9NJtMHIRsdvzWGB7jkoFWygqCnP1R
IPRdM4GjHsz5zs6sJHJI8PT3zpmYgktMnntPMPEURLOeBOaHelabEWp0PjOklCQd
ruXMkCIxfEprPbWubLAwZptMzWvk1yBcFPA1G3c8BiYdznlF8sbweySloZP1ZB+7
RQfKzEXsL+Og8Z9unSMj3v6db9sik6uyfiXJDQ5Q5lRy3/wqnWBj6NcfdPzoUkV1
2MW9FAm9Lcqzm8lJnWqTGqsm/RuPPZidnIv/rds4glPc0UBN1cm4nFKSsjAiTzW9
vjiz1f546Jrt8Z2aXODV/0PXUXwAE0jYgbEaCi0zBkeEcZ285rLQjdZM//7Y3rmF
wUEuFCBrzwrEHMeCAbLywEaPj2VBrBgSSuS8vZPglzPwFvPe2su6tjHw70uVieC8
JQALRocw/+MgKYbfBsg7Xmz/GfDoRjm1iS18ozpWyuVMaOmrcVnZyFogZa7h5vij
gWnquRU3B4Dgb9Y9CgBjW04qwTJtwax0Utqq3U2PgDAr1I2eErPprLRfFjQ/4EAc
9DmGhXUrTpdh2woU+g8qJRDkWR/dzczpUYrL0zWlHnQ5QQRYbcTNsbUv3T9m/kO9
514sraI6tdyFbAW0TnRVCece9acxlzWqt86GV2eTBwQ3kSS+nKHWSMbHVmyaHVLl
UWvmS9tUH2BOLs7DLwwhkrBvUobrKjADqJW9jPmFKNfiDRkf0ZQ7jcd72DqMgP5/
7VQBz2xFOMz8hqJ1+vOVPZRYRolgWTCMVXaXo+2TxR9z54+04iieydwJapp8+2G+
T6r+0sGRqxAsYZ85lncxE3x4nW916biilRTN/elEzmDe//D/3bgj78Yc4+ypf3DU
T/ts5ENfRocWiI54jRmUdi0n8NhM329ZAT3jwfEbSYSh+D7NWcZwkkpnAHdwuesx
o7A191S7wpoYBXRWZZn/Tba4zgvm+L+m2KqYZmz5dr/+h8CV558dJcHXSysncA4v
OM3cCmIiy6SIf9kHodhXPLQ4jEoINGSeO8RujZpUprV/oMHgEqsdmpQ+Do8BsaXk
irYu4CvlcXwijm/gt3sruQM4aIuiz4L0jmi31fHR1TdkopMhPp8DnqrDzWVDwlEr
Zh5irYihvxjT1JH3rt9sYtrz3rTfMzMiCCKU4c8Pssj+2c4uoj5Q/UaQoSl9L9Eg
ui+6Y3Wlqnp6Doal+Wss6N2OO49U4Y2V1EwhbXTxqmJDQqyBzexb7AxcdiYwpGf3
mu/NPR2aGKj0M35BkD8qCNkU2kBZVt2IEzGPi/pQ5V2ZxXBflBf4wd0Ks+NLcND7
rD508vD5Nrizid17M2yZLexR0bbm3fybVwZkIblS101sW0v6hnqjbPtVSYgFGEoE
R6Ks9IZO4uIum27QsPyZLzpooxdnUJTsxomOHNJKIi6gqXYJlTLrUn80bJMXCnrH
ocGcg/9oWaU3Hj3V9v1m4VDO9VFaEC9WUsyAALgtDLEhT1LrDN8z9TgZxmUlBMjD
kAJXwGhFWYAw67ukRO18GDyjlhxTQEqmpJ+HeYRoiSoqcDzkXF0p7k+PsFApPvuf
Zcy5cNBCiI4RHAeA5TbcmxKxGELF1kO36zVlUZ/CnLvPc8jfstcDX5hde7FKcUgE
KTRbjLqRUdn0gUT71BVfocsauR1zqEuauN1qfm4nWBGDwYX56oeyDRDwy3eB614W
pvDH8dAKoYLZV5gNCT2VvDqjwSm+/m/dAeVLYrXiiIT+XoiDCyLPIidXVpHSimSS
fwfkZolXD2d5iiRcHBz+ijXfJaB322BqHO7xsMKxniVrMO9QSgaBDJckfUbL1zuB
NRQD0ZkOWlfs5o/Qcfew6W3K3XC6lkou+qmx9QWzIpeICwIeUOGGNJZ19u4040pc
GTt3uLq/2wXilukixmGxArmhysHKEOn2fT8Rnmn4yIjD5s7OEf/IXbokRTMzjGcb
aLyQyycIDb9G98L/wM7uZkwyUg4bx+j5IKYEuxI8dr4u5LtyfgllxQI2n29VdFKr
liCC3hJgiB0tJVEodGOH7/9UqFECbQBPAjRVtgI4BIeRCSR17lfBdwCai4xeaWsz
VnmooCADSSOfiFbZDUDbzs3F3ri3iB0aj4gRlf6j7I8vAgWXlskYbZTADs9GWcPG
nlpD1wngXHSGGgaEwKMM820G/ZTCE6I1E41nOik8oeHIrsgYC//x97CyLaPBTRyu
WDy4T7Q8qvBJT6mtv61Q0VnkR0ZJ+HN9mB0tKN/l7xA4INKfp/TD5pS+swBgnG0b
B1/uIf0iGTRa7TypTUcBEyDRDRqBlCt2GDbHrIwKaLgK9jUr3iev+W227aE3rGBQ
/pjeJNCazOYtAWgzU1h0GUp+c++edeySd8ky+adbeZQurOePXp61A9YL8vGWnR6v
wd2CujIFJVaIuAQmp7P1TKoEfyEFHiLsuHq3toJqJzXPClQ0yZKJNz+/qoF2ESIZ
9tINKXQulsYwSPJgCm/df8ZjhAd7hccVECyiLJijzYll7ij3lnL+x/6Gs1v/cUY5
pptEGVwLIcLiwYHjtBey1qbUAaoELMg+m3nHJsUiCS4xVucJNBnyhmVYbA3bKr2Q
kBse+mOOezsBz5KNPHiFAZ24egVG8rjYIc56TUfJeyRH0INV8ea2t1OTOIpcQ6at
Fg8zObE8QbRht71/X8CnsCLCMm2EUmjZW/ga+Rds4hC5OG8ZPpfCZG3EZsoWuAfP
vJWu75vDR5UEbqk5pkStHi3MMwf5RyET23F05zajHwWytAJUH4cN/2aSCCO1vXQ1
QH14Ig/LaQ2YuZ9ZtxuCDmoXqvv84pNkORhfv1MFNCq2SU+peZmP9MpN8yBxVxpw
XLM2dyARWneTWUF82F8frfm5VBIwB/JPZCWKA30K9Xue+2Rx5ERsIO7mi6R+OHd4
tyFIN+8dyll7X2q/+wQQsLduoQN1RTblRcsB0UguD+/BOxO72RWvVFbop5UKYExP
bPxjH+ebPdi/EtRVYjzv1jnP/kf8gNV3/refdKp0zS5NC1Bk+JMPUeRuf8U+UFoE
M2vgfzoIMCgDKu9aRI5UaOE2G4fuGuQ5dWCDR6vzIzJGq/Dh919xy+RNmoa1+16w
cZvHeQBDYT0BulA0aq6QttXWE1QfrpNrrX/rQKdN7s30e/FxMbk3E4EcmIKuIcc7
xkjeOoR0WXg8/xNNwqWDnLSb5iq0Ty37jOYQBAeD8eE2CKKb1C+XeUuUbNiY0Hcl
qJJNwBx2ehYKW/uqNOVsrLG4K7O9YKKgJEAfSYOncX2wP9bN8bO5C3ducDbuoDEL
o5uQRYCFAngc79fHz90F2EKRIaBOTjBPbCvCd1pQtwhKOdKsib5SNe3Jc24eZHDd
VjKZ6ei9e21FFzxw5lctO91Eeyb85527GLw/FHm/V6KmcdsJaUsPnJWhTG3LeZIl
BH4sThtbXlrTFpZno7HksL8a7RMwlDcwtjQIyBCV2TtnG0pGCHT/42JlHQR6MLUB
/wtRcVapH6uKYp5NOgH6w8LE8VSRCCkJJmS2jWtjLQ0xixXG/MgRvP94QpDTYmSa
8EkiM2B1SE4Lte5PqiYgoS2N7Rw2d8mB8sJw8jfEjT8tpFYSbvv6xU6l23lP4BdQ
ASau/2VdW0WuKT+rbkf+E6xHyisCRAb9ncokJJtp8A8JNopN2Kx2S5hE8FQQ3FxI
RFGpZ/x3z68nGLz1scLOTJ6pjW9h1VkZbXqiwNYfeKx3WY55AAQCgTxMcm8avIb2
8lyzQAMbnirphjs9hOXQP1kOv9DpZkXou50fnGdWVA16oGIowS68++43m2GGIrhc
nXKCtqK5XBjj3oFQOS2tGHVrHbfotIKOn/yJPXqtfMn8uDJfHFhyRQoo1UNA4OF2
S3Pev7yF0qUK4ePOjPm2bEWuoyTuCD6CUjD04myQgCahn1LCPsZqUqnZMtzZUs8E
XvFzSNgLk/BGOuSTHl4Ic35fLHUIGzpHT1oUESY1R/HBgnaS8i6qLVGLv/szpOAm
7io9JdaCfmCmSkoOYus7emJ+5uS16KTrHgBwl3T4AvLpNWakYuk1bQd6ymz6lNo9
chMgkj8StpYT6s0Xr4WKb8OpZseAyiXXGFkdzLLE9MO39pLtTyodCCOtQ8olhPoM
FlgJEx6wr+K6nrdgwBY61K61iSp/CFEzVBn+729Dy55RFko3QfP7Qp2j9Bg9ZVD0
VOY1UUIOmJ/1e6JCdEhfIc0aQPsDVyrbcqeoSsjGesaQdyxuDfKeEhQ3PqxmmTpL
7XrVN3MWVDfW+BhEQOIf7O5RX2QxXdb0yncl9Rey4aceeQaJDTDaLGC+yJ1LrHhr
/XZirfMn3YctrM5o76zsTH7nt3QmVz2HBd2+7JIowfXW0WlwAG1yAW9BrzJFVtGb
5YbyOS4O2sb1wbvurxBdiq7ObYLjC2a5hXkhtlCaJLsvr9vPnU+BQa5Um9V/f1pu
SS/pLvsFgn3PcybmDI4NN2n1yGn5Ckx0YJEjyLN/QsP56uCwhOAUe0k+dkN+Cujm
X3aM4/oLWwM08qGz2vjD96cWXzSyYmrXM8ia9MWUKuVU7mTprFNcYG8UrYoGQCx/
DPBuIH8JkXuIxrt2GGC9sw==
`pragma protect end_protected
