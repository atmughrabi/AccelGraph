// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lO5ZyTM0iDgWT9oz9h082K1tQoy+sWf77OoF90YKfu4mfUjV5mmM3eYN3qYZZa9a
PSnbO4TBba5BpWid6vmECpeZ2vneAJosNWXTDv5L9cxkEnPdk5sMLHVzaQbka9Qb
9Z3EwYTZqEUO4++ZquV+w0ZuuLfMWOd0X76ZHDycYJc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17488)
z1Z3YlDS4YtOxGok84WsowSH9TvS+t4xSRGVcNbI80H7SOwYlkoKZU2VLa2QXL8e
RDxpSWv3++GNYEj9TbL2TG65DkeL72Jr7bX+IIRoqkh9XWFHR+4JHb/kslE7z34y
OclCsTfcF6/4x5xSGqbio98uS57hk7CQIyE18wjRjwipb0xayTKvKWnMKlLNNi+o
kFPLikg15sVgyg6doN8WVdjXLUQlXBn04ZhL3Or7NFh76s8E6cBD6fpXFmdzaeDo
1xzAwddJaaA2wlIsPScXxlISVDvllu9FvE0UTp/0t+hEtmv7/8O1gNgBPgfnwyTH
v/VUUVmJlHmr/ueZlrIqq2WnMD654Y9LrXbacn5VR5NA+3LPEMJOC9BgH3Qrfic8
2zaEC6DgEi7ymXaiE2Et75Z+z1T4feM1HZsv1+GYoZfNmSndRYO5K45k4EeqdueV
p8ZkbzKsmw1w0x4mCmS3ntAw0gRzKzMO9VHQMgbjg8/St1JXK5SjBhaT5ieBxKlf
vGDgPC9buAFTD940dagYvvbChxlQsLK2nxOHuwBFMXiyiEQ7OGycByE+o9CifspN
Ioqcy3ILcTNkZzOVVpdnEQsQCS18msMkliS3Y9BiIYfRIhxmPz3v6BECac/9OnRO
u3q04FhNdGeGVSz0Ca55cRecIrkA9s2UKoox6TJDhd97FMCVifgh22FajBGNWQTz
qXSaq19sIe+j/FhnoBaQK6cGxFuRc43RmOYQa5mDAG7TAWM4Q4SyUsJxAWqDAiwt
rrLgN0d6Nr1cr3bn7bH3p20lbmOlw2+H7p3sd78OX/5Mu+IRi0AfaCK4V2WdEflt
NGqQ0SF5stcVJtuk00O588kPu9sfBFP5Xpkv6wR3jbLapMr7TIcCVv/zSRa0dXmW
KKjkD3ruLrHh2putjokd2ww2+MhmM9f9I7SGbZkNVXH5Fl3aJeOZ2IY2QjEExhVu
33pC1P6m4XkqhU7KR072nCLoAQ3h3B/+7QoVmSP3Tdu0r1/dC7XmiEzm1WvLvPOO
H9InxxiWhKDDIHt+nxjnYnmXvA7gHOIgWr8lND0F5HBlH38tJlk1j5fbZzait1ha
/sB7pSl7JbDKdAlw9v6nsT8He8iHH//LgE+/ZMnaF2PiaVtrV6CEwnFskmail+2A
AeC761Di2sJ9nLdQGc1a5gMvgVMZZx4CtEXUbbDooMsg7FIFM5NI+URN2lPqgtjQ
hDO6p9e+a40JMsrpzfZ1PTpXx3ra6uCyG5pyrq5+20lK4fu3KSW9EBuyQaQfPH2Q
yqxccAu91q34Fkf8tBE8+PTCCtK+mWjGTrBAH6ZGNvoaj8kMTBWAT9x6cjFs8atq
EeKzgWXJ3emlOSFH5ymF5bEemymEjtvrMR+p+HqbyKDVn1hxkjTU9ZxCdfo7EejG
LCTh7TGrENDKtXdJi+IJey98HCjZaVZgPlI2oxbPvSFVRZNpryf5PBCiSfCh3pv9
9ng6+lRMp1H+RrdFeY5VJGTVT7jZuumI6MQsYnN3HUX+VVGy5qjyyz0MrmT/tuWp
h4sD+Se3tEzF9+EN0uLW2TG+IaIEy9kEF8JppJQt4AFL6+U0sp2AwtxtI7durouH
jm+RIpVs7fQ7a5YdCgwJh4fOwCM9NDnkp/28/59cAP1fgp5gdva7BbsBWi9R+3cs
x2Fvapvo8eXy0hnHdqQweTM5pmlLu2X1fmZ2/aoWcpMEICr59ipHEb7EtB+n6dXN
oepBIYNTe1ezMZZIs/smMRfz3yFve6nNcSHZNiRORCTk4gpxk+YrgZF2sfk3Zqaq
y4EJE9r7g+42ujr222d81MpXB7uH2VAtYpyd89YVPwzxRHpFMg4H3OF1L9N6TJpw
kRQargQL0GPXtXbi6vF8MJTW6Gtrm4iEUH6v8A/NuqM0zJxsqPgHBgDztvCrSwTJ
Agftqt/k3MFEFr1b3f7Wokr+OHlYnAYhf6+AOqwo+JRw2evIz2Wd3fv2gAS2do1j
BbpBDhywdZms43j398x9PB4C3BoXKKZK7/JU7NaLU9tJEEw01x4FeVKAn4i/2oQY
dGhrgN8x+RRHJr+6NiTLklE5ZzIa3hf3GOFGPz9KtJd+MQNnedpoBtk0qg6kUq43
J4HKxqgvFudGXcvyM2p7FApYUmp3WTKxYVv12edqR1E/zTsQl/Jc7EUg/wRH6aDq
Zg7BlCtRa1qLHAeoki/9KgsU2slNiTyIQ18HCA9fWdyuqPTntU1q596FbSI97Crh
RQSiYpRwYjUKz6p3xaCWjAI0n1u9MzxbmSFrR3fjsXf6FsqaAs789dGjvMvShVJm
lB5hGm4VK4pM0Hjtg6CsPy4WZpa7FRypBZOBLS7NcVq1Twj9eh83f7M13VHwBWRG
YfZ1nf5CSnxJG0FFZrOLtUZSeLU57AqwoXnY4cRbb3jAQ6ORD7LnqCS2dxUCM/bB
c7NaDAl58YwO/heondLPV/wECGhNvViFbxjueeA/r+zvRJbTL8ROHFUmWOX8gb8z
9rHmKx2vPdvVtx04KeG+ePhed5ncAHyo8i48G8diT7n1L8OVM/mvd/U2kO7a3Mdt
R4v07XZXjzxBb4rLTZa0zh+kVPX6GSdmF/4ksez1qmIWmvI52Ayyd4JO4Ryou+yt
/nPEwVUfd09YnAK7MGhMnFCe7BTIgyubVIhY/gEVDzPLYAQBZYuUFLgPLthQjuVp
QvHqPaQFkN7m5ou+R/1qZ9V6/SfqM8v5jR24T6V9jZpomeO2W7AmnpWEEJI24+Y1
ZYyPgV6aCqsAGBoZfoB0QDBlemKtMs9yzE79xAAvEYmakiunNS5A7Y4Aapfkg9to
KjL7u723sUM2cI0DUKBgHc8ZSDZuOQCn159u92pAnp0CgZi7T1HuR4IhQUFB8EF0
RsRIpteKINAzij2sv8JfM6rPW15Jgxabqq/7QDoJ8AwHwKJLxwhCyoCV/LFf0WxI
jrCBJgWF0SgOghgEqJVAWL6xxfC5pSJWLz+x0j5C0V7Xi5sSBmDVdicM+P8osR6H
PXMAFZF51zR77XGmpGJWpz1z6xwU+wKj0cxPawgf/CRpP8+fltwoMeXbtXgXZAA0
zedAxYW+R4b41E99D/FX0coBzgEoFcvx85GgTCiK6jdyDTuz9MGOm5EwRw1EZJQ1
IZgs00sAb/jVHGAKn6VakjzYtIxDYfUs8TvwnBGZQn7BHegCYyyyUR3gh4oVirba
qKg3QqE0BuUcfMuly7OngXuJGrbsm0aJayFzJCDpfSajqzt8/uIht3womWH1oTu0
nPAADtmGZTv3ubOmjLE0vDk/uK8Yzp36kdwZx/6rvQs/If1oJvapD/C82kPt+ujM
VuXGc8TJ9qfWvmvlG0WNtnb6dflvIYLMUWZpzgtlCps0wDha/JCkAuXCcOcJep2u
cYQVpmJ7sonuoiW+EErwZRjcW+AP29p1TN5KJCGQPD1MK7LlfAIhzo4wvZu2pXlG
t6CL41FKvIjLjO+7olxtA5NKAn8pGNak5Ug2aTJakDUX6JMpqpKaJkbtlnnIPDHC
h0MI2Hw6mbdmRgeukw/dccrpxEFvMyYv5vJjqw3vZ4fpH/VT+XXXQSAnFzVciI10
0/vxifr1swC/9SWdBJiWDN+t2Rc7DNla7USUsJfgLIO6e1OfeDLrQIZZSMqjM2Oi
NhhmSCbud8PLME6VSbPGYOIKNZGPSDafKKxNZEffQn+iKSl46qBSSmXkP6KPATAK
vdnd85LsYTEysae3Miaxt9AeYYtqV6JVsOby9x4jajujbGfPJY78tfHCoWuQuxQH
vInvPq++AihmpW+m7SUiHMUFuxZc5vPtZcATSowfiS4cg1buxyNbvnFX9t7Ya7hI
pdyo+ennDEgmRUeu5YaNlOrl95Dc8+a7En221nmpiScR2k1atgcpJXkPe++xptjm
Yos3nWRWpnu4g0YgJOlKRWT2Bh6ykoI+Z2yIUo9Wbqab4rFyfwwHx+zS+ldUs0Os
6/11f/yCMSO7jQUWucStSjve68ovVp2YHeC7clJ08uV91ZhO7uRzlCyWwMOj70fQ
dl8seBcatWm3g715GQMvEpoSRXeXXFLjc9TnqSltAIpu+DvNB62+2ulfA17CP0sf
2nMpBANVQZ8oJ/GDHgf5JHyMdokOmxZU2RVX6zJki7vg9zP34SKVb+obBfYmSoXP
ItuNoEPiaQiE90f58cAnWReGXf8FcpG+0LxX8DWr26ATLVKGU+HLO0pPa+ZaXvCX
hLgYOkDDbJee4lyGZxI+9r3mwJBI+fQfzV7Mx0YGiBk8l71T8vmD/sDxQDt4ZEsm
IDvOme4BgPxynayOt9shT5IVKylNft7MzE6kToZjG//7sRsg2/ka8JmJWNeX56K5
lKg4+VYhSAqIRoeEXjrdsN1jon5GbRlgoukOJWHJC8Hefb+fzkyD7s4ccrWzfYt4
Faa25tuZ0viQ2WPi9R8o3cfT0R+TdONNKi8QDY5/JRAMb77/0uM9c4o/tY7/eQH3
fPyzM0uoo9DKOiT/t3yra83PFVjrOrij+ZyeiyFjGeDcnAQhWAMXTxfwBD0URpR6
ZaDfXwn1dTyxDdUK4BLIcszOYY7YJUOP/4q2r2F2JP9JUtHpQd7ArtbKG0D/Kvhi
9nCw+RODTs17RqFw6O0l2XYI38qmPBj9ZcbBYTVExZA5DZvo3acXS4ear7GtQtjs
9jHB+7LqwWWDrJSjN/FrEY6pGiS82eMjOMuCkB5QAXI0jxy6wJsHkabDMY8xnch3
qMPkjpm/ozMCqOvysGQuFu0dRDV4SfAZTKpS7LjZG+NcLSF9Rep03CH+QucIBlkI
I9Bbn7NeG5cbEYB633L8MHNC6Fuv2VnwrZW80dadZjQEu9it2td6O4i9WiIQussG
TupmSU0gGvuQdjxygFza7Xx2I7f8RdMkuPD68+8lNGp7VsVQv/GkGOAMaRnkFVog
rRLwGZdLKB5yxQBykigbwv0y+A1a5F1QZWSz8hXBRN1SHRNW/0wl9wYjG9jVcPhw
nfW/kr5ZEsxJpK+fkm22J9sZeBcidt+pLmAFl0pwi5pm7GufWvtrXO3UmxQ+G5j/
opAfKzlqjo3AJ3Pqo8sC9qXpS5yreIrZYirFCDU840EIzuk99CqcsrppluCzgS0i
2640Vr2WCROnuXhZtF5XjXUBXyXkNT2m+4h6ScnntDHAOHeeJhKx4OGx2GIGgi/E
/i538Z6dSEh5wrTmDKz/GaSwJS0C5I6OKkZjAEgX/fo3Z5l2YdKByfehmRT3hHfg
UZIuJzqQ/SkJqUt0chiRqbCeYPtAJ9H48QjDwhLbQEmTfKnu7+MCxFfnFRRYa1+J
/f3wpysXO25e4b4ri8+rD80kJeZlEECE3Ak5tfvFMkDvRxGJsOH/hzq2ekLpi1lk
tyTeIIsTqtlZuuOXAftd3aulLfbwRs2rD9Mm7bjqXCbUMOBQXJCvnw+a9oeaB5xL
M8Yc9eUrWttHcDZ+WqTwOVwMphipl/oJQsmZ9zVL1VyX63RyDFSz8p907y7/mJbp
7f7Z3SPcmHTCFX04P0ZBC/NF6/62+PLA1OovLTAbIIfDBoKNdRRwRmnvhfsGc4gH
xMoRg5UKOx2N9i6mjkW0CFQb6AcvuJ1zNEQT9/Inhkx5Cfewng19bpmk1qwef71H
K1cOI4SJPflZsoC0IhRGyyh39VAV3SrmqEMSvtuIThFha0Ja2k8546yjjmWWLc+k
H1ioe9lxnFmuQEYemdHOPqXJYIV4P73naYLkGQKC5OMHtMOyeoFsyEFr9lfp64/6
gq5ZVut66wlfhc9LXiFdp7FENVJAUvkuqVs5RVNr8c8mOgxRwvZ04LtavV/W4tBO
0bjT31StUyKWb2YXtmjpthcawMWnXzttPvbqToBasQgy/uB1GlsCVWRaLixItnFK
o3r03YViC+kInBzFbBdoGwM/GhhmvsLByMD3AaLeZMkKl2Dsx077CNfu/sWlgKRB
hwjmo7H1GE4xlVm7YAfH+BLbWscZM0aaxXPPbNEtgnM0jYKwCJZV+yCUzEiU8CpT
XhHIPU4wFid/nAfqb1DII70BWQP+kIloN1FJFq2JHZfWdBweMMwPRNo4BWW3mxIo
BPN95NdQnVIQvmmrx+5hE9GK48F4h7Uikqv1cTaGZNbErtoaeSKn0gIhGAOYwxkZ
ym7AqjXhZuV7YpSZOAYI2a4q8K/8F6F7GjRO3zwd7V4P1HHrrkB/KzEyxbSsnxls
LQGOF753tQ7K/9PDeO9wDGhbkh5qXyv01wNFGtOZtFC6UTgufFfqVWvltViAJfvN
zWzyUQ+Kf0+fKDJS27IGW6znIICK8XF9cJgBfCb9DJK9IMohrO1Rc/TSFvFqEW6s
HfZDUBVTRTCI4+7GZ8ZXHsUuq2PjKqQ+54Vm0SSjMIsWo+85A9yQkQKwx2Tsvg44
Fa8f+5B71GS0hkvlotgKM19iU0VzB7L0sIU3SYAsjDDVCycfOKWjcyIfH4/UAyAR
uy+luqETqV8h7yKd862e5bviP6SGXuqUwjvpVylFdR+zHDQa7duqadkz7JKP72EK
tfzGJYrfSU6qKd/H3gHVnvBcvp3z7eImnb+GOeO+ZpyYn0/DdEyyxByoh3sl3MfY
M/boyk5xjktUbmzkFrVFZWUJltIWJzcb9Wq8RSu9pOvJSm9/Q0ck6ThNqrQrXZdk
m6v1lh+3BLtb076M6/YIUayOzHe7Fz2SPtkMIsP9hhL/Sdc/6LX4yTU1XRun7h2+
vkGajeOQc4CPzja7n+CPOW3tPVViiXkAU31PYkZ6E3PK/spmYgWwEwM4oXa5TCHg
177jJvCiuvNBQ3/laRc0Y2kUkY80lU7krGyWXAWe7vNovEGkrFhf9xAp5tBOmsLB
haM3SuU8w6R9S5ws2kUYGFx1efDpbhrr1e28K5Y+09b9XGWIfIiq+9N4sXYr64KH
DFpOG4O99zTarZfOWz2UenGP6JmaXb0f4pqB8jpurKABacWZK19jBb+kGoQQ4zqJ
tIGtKCA6mEsjqSMe0Kvi8urFvXQW2+bxRWkwt9YcXi9Gb49pxUiFiTK5Ps5f3TDC
uV3GL/9D01dCCoIwvPqY+EN2pEOdfvMAG9rVoTCrWsNLTLzpflqgku3MaZkNFUkg
3Dahza05wgBa339zd88TcA4SwfyVWkWhRYHfkc6ia1DvHvLypS6Rl9H+dxCBDX+t
oOFakApHUxAzSvZxoOxuAc8YmeVag/Bt7iQh+y+2kCwCNpGj1NZBHYFYmkWoLa3R
99P96Z+ok5ETOCFCc3ISgAp+hj9/t96JeuqRKA9Y7ggiavi+vSsj6Ud2cg1o/UfT
k7UIPzMjkrKPOD/p1t0Kn3jBx/mPyqmMg+qrXZ6tZtmAghyVr+eEv9M/HeLrT9rD
ZnNXMuXRYGKmp+APUCHqHFbekMEXMdiZ8STCCZ+PGod6MwH2ps2byVIpDQfhz47P
JACgGDnUpbsoohVIrVXOzLE9VuPpfA4aF3eOQGh/XhIFsOvhbdR3RYE5nUI13+B5
ewSHqv5C8H56IehleX/g7m4bTdGFLt/5F0dshWLX2JdOQ9+x1pHl3ortXBi1/PgS
svKryapEAE7im34i8xgTN7jXxic0e5vcOwRoPBiJGJzZVrc0tE/IOlIAXprb+0DB
mJhfq4MseyMTAE/Dai5iLW4xCKzkxqjMb6z2saEwZ5b3ZdjTQGYZQZlDPywEgH7I
0py27dbmJxpPEpIW7SeD0q4EsTmO4RijLthLUA8EzKBP6AsWb4KWB+TYsvBT/ns9
ZnRXXeutmq8LZuNUE/Qb4jOJBNycfXh8zCwwXyKvYVhgCuHWnxFFhhG+Pe8lNY6E
cJr9vejBu3Si8fgD4L+waEIgw7dz5o9S7hzLQvs4DJ5puTYHVFWUjOZ8qQ9CGIKn
g2rDU+iQspl3msTwSxKEbIotpvxxPF0fpzNIDDdVckJ9CdZrAyfRS7eEswyae8QA
Pixc+Td0hOc6hXmoyv1oyZCjotI24aZn48ynIE2iSYphpR+6XmpE9TD0k9WHTggx
vF6V8k+mVCrx7ihnju7Ds2CuaxgqY1oyIJt3LoQQHD5yQbTSpBZIbf+ndiFdoLkh
TmnR7DQ0mq3Vc9CTDvqz/ORWQbMlPfOm19l3yNGyzLV4ZevJq2jqLvKJKvZG8CsR
nxI1XmY6a1xEYefjKWsBDwnqSx/7umya79b/QMUHFXeZ13S2QNmH3jBgRD+WCmU/
qa7FSd5BOP7Efp2dhi6/UBsh20BLttS0dIjvPCvch/jQIOQW3+3meRzHsUlr7V/T
tI9anvfcHCB8SfyitJFa6sLjqyWJPqrubIouFel4UHcDhPHiF3B+9buP5A9/VX5n
1RHDE7KimBtEWr6/BoghIIVLm9fxODpgyMLMImRoH9GyEGaRHFjOYQ4adCi05SYi
Tz1TOuKy+hGCuDLRavLLdw0b7x1J6xfIR2xhdmhzxA9M+xQA36SZVAA+07T6XHAG
BcGYjyULPVduDP9cHb5Y1bG8Y+2az+PRHaRqhtWQkjc4RvveouTOi37DhhSfN4nC
OomF+9ZYA9FTTobQ3cKg2xoIQ+Clgn7MPtCcNXIHP/dLImKJ5cYSM6ZehVQNLVsZ
8xHe1YyN7xOI57ZOEbiXI5ipVuGf6hhNY3G4CUytxEWtdRqiz5EZMOiLl7E8J9l6
X8PJ98/HqlbI7MkzJO/LgNMeNWLXFhojmUj3G66yNkmQuwE+OJrs2MBw0WPfG/A4
vios5lz+4C73JyIvmt1CNJok/TvldIetrcU5MRvt2lOetCDGl28cA4tYPFsmKuKH
3TshY9piwJE0zNmnjWm4YPaCDO1+8QixRI4XkpxwYd+xSuVWWjmsN48zfA6DAfKc
P3z1QAwfLjaHTsNjQdUhwwkKgo/TIssb4OPfWRXXHEPfNqmCraHmrH0qLZUrnFbQ
W1jNzhJ4034ZrTIGsf31NsUCytxyzuWGPsvJYYnvfdieY3NHVsRUEQaXFilYq04t
zSYj74IayNMGog05nWcrxeghkFlnU30R2mSMIFrzszOU0bULNRbx79SmGYfJ1CuF
v739TfCWRSWqDPHW48adY7w7Wm0y51IcXcRhHsB6VK2/Cv/ANLPnoWk1pC+T9yZy
BZIdL0p4hL6FldHc21iWecUYw1axiAcdHryHZzmq5xUXpSqL4RwNi1leEDwb/6st
pVLfklHuNUWSfS/t+XUqu7y7Cv5rqxzIf4TvXBaU99AiM6AhpiAjxmICQ3l9fIxE
HOa05jI6xUe/YPumd4aex3PRi68SSsHloOgOi5poRj3mAJjFJGKrqn9MTSW2VBNz
DX3gDCNEazfnjOYqgZR9pYe01szUWBGMR9LoejqZMkTKgvOOPT03rMAL9i8ndOHC
KudzeU21xmXhO6OP2DS71QSm3lovHRlAWsn4pzTcKPx5lvCc3R3f67ydtRKAv8On
ZHhUSjpsHbZ2BLgi5zqvGkHDkJDbZjV/PiMHldN/C+Pfo5Wt90W9xXgGBuOSNa+B
Uh3Oelat+6R55+0IqpGGCk+VrHhpbg1gUlbQLbwauf7uJT58HsKTEZPzxJIK3jWL
zvqNqZvtc0DT7uMLKZOY9QuB3ipVaUm7EeoyibRoSYfxjMDA3wGwnB/LszTN5XDP
SiW8lDHTZBc0G/zfD7ahTZRvCFWOGVIez0z4M1XQKV2uMXW8UD3QKCfVTRgoLuhP
YkuQZ0y4QhYtno1LuFUiyRnaaOiEtxzXE6OovJiIStUNraVdL+fRivGW9Q3K+hyo
n5HrKg8z6svUlqQbvGjGJgI2TpKISQNS0KIuQU3FSsNS/n0vYOmGCsKhD/wl6kuf
TD+k3KgqSU77Uf8hVnlH5gxgOijkOhiZufDZZIbV3dWY0bj2zg9U+8QsFyBUd9N9
VE+95pdWL91yINGqNxS9ClyeG8ePsBO/vQSvCyCjd57pPSRsqwGCn+y7On4alT/q
UEsdY71SthralnxnwgUaW5gqOUNGlNCNF0zhws75xIF2dtbWO99zs31zfNao4v88
H2PWyTtv3RRp2mOA8ahfETFr8/albIEdeWtADrd6ZpFjwGof28E8XvrxLi/RhCV0
fwvl7C0lYEqjXlzqWhmT3VkUHooQVhKZtxS12kVOVK9XoZ7Kx16uGfqc+h3bB5iT
5GCIrxIK+dp//q5irj7THaq60Ebk2+vsJhinHDf8gapwX4dVcbvrMxOSbWNi91EM
WaIGWL/FcDlivn0iQJrQMOAp+l1CqWF24UwNBx969aLCyCcFUQpQsSnPPzFNQR7y
XrGVdiVBFLPqfotT+GTsXDFjwKeTdDhANAQllDLnGrK9oEPh0bRwgzOxpunCHAR3
ui96dyU4yRzb03QFxHkPjiSIB8L2aqophgfQVk2Lo99NAx498kQNTPXH9uaR1q8I
0ujuYdxrCSwZPS919c6cc7IDKZYSbi+hCf1w5jlU43TgcEcw+5++VgyimYQoFSo/
HfGS2Iwe30/POmTgWrJlY7ddifhyQV0BTHZKohHB5sZayRbHsqhOH6qK+bwdS5jj
y+yB0FhlxvaGxJI8RFcIjikYaWNfOqM3DUrZtvEJKK3Il9/Eq68N8Wfk3wVWCnZw
k9U+Ys9KqDiIzHUTODEwf4Nqvot8Q33iBnbjfI1SSjM1M6hf1Sc7nDmLt1VT8i5D
1G2eOK3fnvjS3nLT826yTPCilQ7Tq+NcpQFTwjMsrkYZBBPLhxz09Fq095H51PLL
fEjU+XBtJdBG+YIijuWV7wLhk6JyFojsIrivhKqAKAbnidwtEPcAXbyKFrooOk/0
31rF2y/sa479UTPIBAaKPmjCNbW+mhwD0L4usek8M3cL/YAJU6SsPPhJwVrnhoSk
AQSCKLKh8MDP1tk4PwI5MhzitEJl1HTi9WV0HI7n1blH32E9c4pERqV2WWliRhsV
ZJ309zRd6f4p1ooP6m+TUUFWX+O0d9ehtWj2sq08QGlVtg11+vafHgeyr4x7pizv
J0+GC7yhbkz87g7/SO1x9j19wyTqjBJHsstfPXsjdMrLcsh20n15zNrELEfdaArf
PLo7kfqxJstk+qo4RTzYgAUq0JD7ncLzSgXBUorWejXxj5pgBYvUaMo2vG5wvcYc
3nkCjAmkEe1FwWgAG/GB9H7YuDdDsPxVQ0v41nc3f5fvyHHaQGuhlhIjLd4dZ8SI
bFGsYFw1tTJTfMwTLg5AVb69OH8uwG8mBr2LcVDUooA7VkePItYGb01qsBTgGLp4
QmO028oY58Wf/V+uctrEO2qECnVnyV5iWRnzGSeDtSbwMGpYUFLc1/OFIeJj7K3v
1ITLMoYTCvBj4MOTPlrQV8Vq8HtdEyIcstuzZ4BQdp5LdyB6mKKSniyizno6o7ZN
1jic3QiRZIMyvQ9pl4PCEjCa8KsGo+oZKRklUTE0OwZCOsskGr2rP5UTtq5jprMm
evDb3SnonO+5RW4H85Sp2XVCA89ttx3kg8hGOwHZDlQKojpTynxvo3uJUvsB1fAK
Kg+FH0T4ZFgvm+FklcclbUjkO4DF7OvjJ53UY50NmgdkFjF51a4cq0qL+ir1xY8/
aqiY74M/AGMF1VwEyrJI3fhWCtjj5F6czPP9DNBFQqj4+shcclpYpRDWFao3V6j6
6n3rGqM3bFXPqLcaE/S5J+/TeMtuIIBQj/XFcT94B+MWl5TQaz3A/pvFzgHbEvSW
weoAD+t/DwJ4Z5BDYNCUO44CHkh1EBraEEievnyvv2fk01W0vqmk9zjpS5/iMlk9
zAplewuoFdvROLxYp4b4dbprh3d4w2FTG2ZjDzqT0BFdoCX191ziV5Eq4MR8MTTb
KSjYZtgy/2D/rr5/vq8dE+leQP8QuYiPrR2GO43B3IMmUO977oCzeN9BkghNtutd
XWVu9a2r1B1eRiEfRYFLPMrrcojkpZ0njh6FC+o2+dxv5xB0vUIFWwuh1YIE04Ts
suaGzJYfINxBasoA4JcZ7k624lcYBMcSIFf3OcJoZd1hSOn814Ln+B5EUs3iZwHK
Fgb1tD1KGRrBxxTTWHO5u1vrAD829CTbb1UIUyTpbnD8zotZqt0Mi0KFc7ImLZ3W
wTsq4SL3OLICxcgCYco6kEkcwwSeynhV1LpwfEj5KN6Tb/gvY1Ta4/PE9z0L6bug
ntjFlWEAx7HGmPJyQWJwV+PNGgmrYBmYZZV92VDFOk9nAgu2UueJXB4VjVd+D8nI
NDjrOx4a3qVgv2ZvgWPz1WNhfS2aMTJL36wedAT0LRVV/Vl8YqKNrk+XYNUPref9
7PDLIeP5FEi73kcFc6En1FzsVlIij14gOrr0e5LMaI2VC2NgmF0ZhNVc71KZBNtE
yB0RQsQJofsEteaTthviE8SL8zsHtUR9bqnR4E7nbzJrhni9xx9osNHlXijYjFhq
QL7TjGN9AmMUqg2WzrvQ4M2ekUcAmh7PtKOPAPRQwhWtZ0paibVk2D9mlxOVAK8a
FCjF3sbcBYG+gHRQhvqttf6Btx3J5FfNyf6A2WevdbIYgYsTzKwty2pLfagJ4rYW
jU33DH7RPM+JIiz8Q02o97QtWM44u7GKkwgC3fpXsVKtof4e/rlm0dOFucE9i2Yd
lbX/t/8jcIRJzPtulhAtEEe1qSbc+YcUxpfhhtuN8xJpsATeCVGj38WRTpNuvIIt
Rwv6L69V83Z59envcvvd7UztiY/GB9G0FvOjGtmivAoFYIqR1BxEN9h4GjI9CoR/
UnJ7HruWBKlxbANS/bLDYcuogiqd8+dsfTtwsy16vqqrO3Fj5goJK/zsV99RwyDz
e3XUP3FahRoKJ9560lP6O+3TKpIQiX3jHjorWK3B5oszOjL+5ukA7FRU8/Ua9Gdx
1LMCDzkmafKWKwjOLrX2+a+eNRaEsf8cOTU3bNn5SwnomO0ySxHrqUHvDhreyugt
KJ23NDf/9Gl5ipGp9Q2XvFN37O675tKK1GHOxIUXEjpQWiQ9ow0J8fuHGyEVF0XC
Qd42D9snCsKtU58ZKN1xQKn0c/icTuxkilUKPBZmKUjkV2iXLnvgFfJ3qqHbF6QY
+8ZMl3Ky54B+fWQCFIQHXFQkkeO39MGWg0tarPYoDWrAvUSMsSPVcO/5LtwOs2CZ
lvpPTicbPjgQ3NUzUbzhvPFsTz42S+xijTNtkGJgubtxtFVLtZ/fYITkLDQWEPxp
4qNBVu6LU1NKuINAz4bU+g/bro4Vx8l1DeZL4cDP04xrHLiciTN8ZJkEd0kMYH4a
qO7/Mb+6PpUrV/mS7l9QHNeIISttaMf9QEIxq6CYClK6O+EisHxeqk0m9TdZBxfz
UFIZL45dn0ZPDqq+IQ4UZkdaQIRAUe0D/Q9wrFqFJf8t/S8RytUg2nhORpoYsABA
YJj/Zf8XBzwcK4Iv7s/JTNXuDVVA9UJDHuZPad30M8aqUyxFA+NDzRocC40UZq4m
co53/z4aXIImv4cik3CxTRWc7tWI3hgnoKIQLRGHFaJwLdSf04zyaEKkvQZq+Zst
P926h4tIx6KMBxwNobSNNhQSmAmOXMUfEOc0MrmfTtDt+J02uOIuK3JPbgc/cVfi
hmfck6I5lmilBJ4JCUjQMEjkOb7PKpfWfVWANA33S52H/4QpV5bXSDTjjRXETzsW
pAZW1TLmCprX8mp2h+02qtYLWnukwkP1E4+nE0rU3ltPlqORgqfZ0KhkO+PM0U8b
MFAHjklNDiwELDGrCHdmSWHaFS96aEOjwkyDmNatQJUxnKgS8bTvq6uL+Fo5mEhh
REOhbNBgI0QIImztaqH9dGbqqJZZFLl0AfoiPGTAZXqZH7jv0cHRwSgtuowDaCoO
Br7sakCQBunDPo3ogimk7qlvhnN92toYL3WPx8ydUi3Y0QNDxkQP0ZckZYGgIOpr
osrVCql7RKVDJLkOqrIDW7oPRDHv/X+ioxAiwAMQssMnp2rQ/zZa+gdEvS7yRYta
SB3RTt1SsZSnouA3rHIC235BLAe2EFk4J1dwq0+HFwxBwM+IHPtpiDJpDoA+pe43
o/uK0Q08nTgz1VSnm5XKH1KnoEgxOgYIRSaqgy+FpzdjlUYW/4Y1VwYd/nhY9m7Z
WK4QAg+pqOiXNAmvYCyiABfNZffowFDRrhBjUcaoz9aQzfkLNelgvWCFkQGD7chl
6n5WyHC9Pf/jdq0NZ9yrSPQd/aCvbDcfsRtJC51+j1fDOiCXnSh+VhyTilYUi2NO
TaQhicSjZjbR8D6Qb+B0ZvRiTzdySotOB01hNOmawHh/d2mGpw2QUghiDCqNaXlo
FO0FjchfgSKBzpKE3O5BZtn3Y0tRqmVSm8pBktWdt6/GrBJaT2NtnNns3g9wEnyf
TnWB/o48ONEB4B2klwmqu9aqljIrLIgNXWBNtwN+dbIY3RMtgwjjZJ0S1GXh412m
5DcnIpgA5s1nkljok0PkLbiOzpOtEVQUjngpuhVztIT9rKM5dLclr0JJRmN9rVI8
NPIzP2jnGyscpwwEQC8q4swQwiOYmFh2XGKt4q3zW4G0IfWAmA2XEjNJrMjzBdFG
1Z7HaVE2IhjZuvVezw7oDRkeTq3F2ng/dWU+oO8FisErpRniqgz76hBLwWDv92E4
xWIJNVs9oGIC10ukNpkIiBFf9sAvi9hPtS8tKS1Og+UQk2yfqkjP8FRGaNccPKTU
5cpjRYDR1e5k+HhmTCHF/HM4C9n8A4mw1HsBfciQynjL2s7+5X95lUQlaxNrd+6f
vHNqsOre9WEjC+Fg3D9pvcYyKgNWI8GnEZIuAUPpFvrxtbTD6oP6jXlW0PC2eo91
DCkRwPTzIJfBMGiv4mZnjvSUny8agwkvNz8LwimddScz9LzfKo80fCpK5AyQTKYw
oSmclTLzTHBrr24CU7pTv62scJfU9PYEpHoimADIUD7tKBiuboU72LY7jv7lMMlV
Lh7WD9DZYVLE9G99RT5KAaJjq5+JA5Y0AL39I7u+/ZlA3BpBIB1ho1ZjdBv9c2WY
AXspgCVQlfR3m9EkrAlhodQyFCoKR3Mi+ucMdMKw6a7wsIcFDq+scDNMkmGFKKpM
S4duf5nSK8TECwGIBubn5JWnZpZr+2mRCexF7p0IyCaLv0p2HS0XZFdIBz6Y8yud
2wgFy/bbBFoVLuMFzs0OHm9i4LoamGFvYo8AusaDmuB/4uMOxeA3amNDI3FBT7jR
6VuLpT+Rf0IjQhhbqhSAa8qIH2E3jO0dnk0i1CnPeJ9KvM0Mt+Svci1GsQu8XKBg
DwxoYRKa1n2bkmz1ecuqBAH6bgo256nUF6EquDiNYP0XzMw++RS0HEwxEyuk9Kgu
AXTstLxzX7aA+juwVX3UBAfga4vUZ8qZHtD/m5VGt3G0b0+3N8OR22uhZYu8SsNw
frzsXh4Dx/CNTZxGwOsiAUMUDCwx5yzG7SM9CdOcQL9myfvs9xLo8e/KRR6Wc83C
fD/vDx+nzGlz/SO1jDte0xE/8HG/+B7QwHXKwFks7ieXG2JN4x/uqy6eFCf2sLn4
rnz1ODhwLyeu7VxohWuKI/zqcS4zvE/x4PUNaUa4cjYrNXhlg5GmG6KxreO9s0Jz
vIfUlrds1qC4Lqe3N9q0rwBXcYLZT0jaXAU5CvnByercVAIXXiMygd71hhiqcW0q
KwCb1zZdZ0e3PtMDuPL4v3iC8GluJHRLRvbHlMwrPS9PquQTrQlRq7r6LvodWypZ
t5NFnMJB2/DXQ7glVEeiu4n1GuGoo45QUASiXMP+eDQnRlnU/CJ+8XDF8dUtlqwa
5tpjpog43j9oYkYbg4keMkuNnEbfcpFDqEpgxqoVn1Pq7J6MPyGusCO/eNFSJTr4
SS/YrfToq8W47TzG+ghlMm9y4GLN+hgGKUMPWQ1tiVI6LGFFijz3MlDtXqVJb9Y8
WrLPaj2hddUeYcy2VqMP5RgN+//nUdDos1KXhwg2igHSmgMMrrzGql7qfkzFH/8e
W9YWj3/AcFQiVvy9zb1/6yvvgN6I18Ef7y9P9xccpzI+JNV8cq642rfm4YATCGNU
Deou6BawC3k3xAlkMF0GnPy8dKvykRciMXXqVNqkcM3W63AzAaseu3cSjqEoOdXj
nMu6Qy25U4oYOTater0enrmjtWzHq8dcbOZ+X/oYR+Jn208ww4D62BAqI+w+g25c
fA5taFwAWwvkulROoCG0H+W0o2QnJRufpYmr/R7moKAJ+H9OPXRwlDtfSYW+ij0k
vzCp41+kcG9VcUzNTSP03meCWoGUgomkIng5xqtdDwLeXxmUxdRMhRkdXnNxJK0I
NXrC8+B69dCl7iP5HuRVvCqichnHK8vkWFeiDHyHO8ioGwtZMLm3vFnrVDt9Dkd3
1RJGVcheTenswbPu8MuM+H2c7OX6bZeQ1IkyHm0YCp4BKZfM9uztejhTOcaISBed
DkvLiaWfwHDCJCQLJXmBcET17obDrYdGiB5qGIa8BVvMgWAo33yPC6yKMzQACwGd
ZBCbqX3IiWifPL4Eyg+KpjlNDFS3nf7s+PP6WItYsXg5U25my84BOdN6YAal4dET
ktyRWyjAc9wxmZgBLnW2Hx87SfRpQ3GDRu7t66O/9JrsZblqLQHcU4trBF4GJf5I
OQ3QwS3SVy9DrD8wvG5+0Z9zmyWAA/xmiAfk5TnLZdGL2Ty2drgUeAATjcc+661A
TiVWBni3OnwKRvLiH1ktpB7ulSPTeOeSOr77U71EqHotta7AMAPEGDSyL8vScjBB
ExGjCotQffON/4YqYF+sl34wzeYhnJYBusDBKKHbUetqTmNYGGKg0WBXkvUL6nL+
2L1h556Nu8Rrbf9VM3MVDbI5kwFrOqhDGfCPvBKj6stLurUB3zCSednykfjmXwLx
tUmmP2F3uFqRZzXSZ307MGnLefwsa9wNu7M482CWB+AuDHVC2je5eXlHoR1Lxh2v
BlriDiZOEq5AqObiUeW1I5uyqDtT0pGG3jIcJHRMrahWqgx/zgLnRYikrtIChLKz
yAZCNL6pu76b5sltHDCnHTWIjSOABvIREnUHVyKRU8bv6PvaG053FKowySWSuwaF
tvYbRbwBIUWixO9wvWln76AlLkq4+YU/XsZCQKWF2NK/+b5RLWYMFeRC7lMzBkZI
Uk+/IQz//8tovvrYYJov/o7U2KXSNPP7sSZXECrwFu+gLyut3YHJDOw3JoGny43G
v5STrFhZhl6H0a7a3zcGZhzRtWz+6uzd9eFl4WPfm+RlKFWGvRzbcPYX4P3NBmQF
2PHMObsxR95rBhyHU4Askw0VOSyXbPVzfahkaYi1zsEKnl4dNcyINgQ4AaAWoZ0M
s+kMM2mwNddVRYjjiX7UiSHE4EIKdD8YJg9rmtB6hNH050prQR3ofZc08Atm67tW
g/oeDHVKSgArh+GlT6yMq+ofIYB6GyGmRFNCnaJJuQZPVgJv2i2Pd0Ms8I0rObih
hqSxrZSJ+1PiIi7CuEcfhEfKtgwpHpdulPJ5vwQg1frN25CbnXmT5GBDuTblnZcz
Q5ZGQd/psoxfjENvlmeKksmYJyl5k8FGOdcOtdfG6lcPx3xYQXNa3lQgfgkC9lGp
V95Kbl5271smjT4lhtUdg4maMn3HKsvOgcdZVKCDxpQYxofCE0ZFS/QD8ccCtxyL
f0M2DaLZgYjGkGm2cHE3qlrWhyJBWA1AqZ82NfRtlc2vJ74Nlb70kqRQIDdW18+I
y1yI0NZxPo6en9wG3nEVgf/R7FNQ7tTsTL2nS/2WYrA8r2CIVJTtRAgvvwqgMg+q
YkyWw6df4bfuqg0Y9yjjttGviRWH5129WGqnjSLVL8J/PHh072GQgzKsIoB9KkRy
zc4focxEP+HGI0EYRlTmkTEc9hQaV/224JwqAt4dlMN6gSCz3BbM6bn3pSEP5l2k
bfNdOM1z4yfOAbB0eCWl5sLXN/NGKssX43lZuO+XlXZksAA4yVg1LeVfjrD9IoJD
9utw02mSJ2dfaz2tH58d1OhXX73gFZRow+AMsNgUoFMg1zzq9frTm8EAYO968cn7
PO28NuwBqbatQkermunsEsP/uh7r8t+sFfweQh+8RdfaZI2tVU/73+9QwKDEk4nv
A8OG/SFSnAWDSQGZBOq4skl8t/fVG5L84IrgrHFDIFPfAFblo9Pvpfcfd5wjnKqP
jOIFrZRv6YF61whvsqnSgGqMmiCwRDrgrz0240O54E/jK2Y9KOIRvuy3JC92xIwP
d5SoBkQbqfcvAr3Szggqe+6i5WdRFTUOg8+aka+eshsIzvJpFrSF/s449jNSuURL
24UOXg6WeFJHP1KKpFCr1RUtiYoGiQQBaEQbJZm4sbbj6+Ut97OUih+yNl/tqYo/
wycnw4MlVAHuT+pZGSicsKSQfdpiJbssgDvhvSj6WGeyRLSLLYC9v/vdO4oX1quU
4v6I58BKexClK7ph6H8MkJ9Caq0J5qCNRyXu7CKhF12FBbfZ3UO3vG4xpTuBnLA0
ibI48CLJoMDJAJHXh3dzdAYNUNTJ4X1OoUEywXyNGn9B3CDOf27DcpYK7NSJGtgV
Ke2rhcRe6Rf7p8gut5d8cNUpQdGf+o4vhEUvJMxjR6IO89bhPkn8yPhsNyaf3YF2
iaaniqYe1qy7Ig+3VgtGuRg7+rZJrDu1vYK+9AEHAZ9SQe3FpgJQlyiaTeY15Um0
EWYtwUs/KretRt4XRqyP8XM6S83AiOxAhyrfEU0UqC31+CRFSnTYy6kJOFM7XKun
cACHTT+bxjYi9741/oF5IEsSvLGK7NS+MDhYGVrXaYrUuVRAfHu1ztiow+pLNrQL
w5RaR5v8RLSZDDZeLbVYBkOftCYvvMdEXue3ddObQSGBfVUdpn20z0WzpCXMJfg2
W+EmbgRDUsqIRjat4y68+s7pHix8J9E8EUlkL84g1fzrE72Dg3HLI36c/sqmGN5q
9+VDUhsNnef6QkKurH8NaRHfEo2EZEQJSH9W8RyCu3h58kRGpVguMmb1MM6w+B7r
0VRHdHHPzgkQwX84AROgK5i8h6ptCh9fYJwrFJnws+An+w6+xxKnzGGpGKjcE7B6
HohFF+iJI03BOCqkcg2A8l/wPllYu7BPkbvMrRfprV0J3zPpOoJ/yO+4UAREdGRg
rpNpiFt5Qc05ionEnAjdvgLBOSZJCMadeFvTSZ0iEL4Yx8UnE+2Q0bDgOl+3x7kW
z6O+4o2ny0XSknSRhRmBcgzrjsWsbZTVKzOUuhMj26ObacXIhFOSKNfGT5P505nk
j3Q24V1GeC79Wn6m0U1h2fb0hpJwiRxd1uTqmkdi5d/gDZmpvirAhPRII5I3wfx8
D0NSij4nMRYk3jcHAUPYxAlk6TFnavqQp9RFX4UxyLg9VH0E91hue09iA/txMePo
yj7kwTBPO/Bb7qSDrsPA9ztlaiBPHKUFphtOyHWk/IUNB7BU/6JWgTL47ITIKlh8
rJzEZJb6i3oXoYARVCIpHtQ1GyElYv6T7JLXgX/ACjxqD5408/DwEC2YrsX0jwjR
vg5jO8fY30rn16TpXE6QM8hI3YcY+ELyInbsloy4eb+ZrSZFo/IOAdcUTS7SoT0H
xvoKuSfhlawS74gpGPPbt+GH40kyE1YW+gAMqgginI/pmfiI2sLHmirVvtCde5BX
3w9i9glKUfX/XcJ4/C9eMZyE3340FeGSeCkuZmw54SYSkcx6T2qijaznamJGGvK9
/jTzjgTs+HrJ23DJrKINcklkcg1YYLzjcKxxE8I/VEh4LK91ZAFXC4VazIi1aMOn
OVB2fjF3MfXKcdkKeN+pDRbO7X45/AmmELuqU0pWnLjbrcXDpAFdEnrqkOEwXJfC
NBU/I1StshaApbONTCL8HTuey9rD78UiV/cYxhfoPVREJMkYbvrq33zeLJBiOFzZ
egnavDNkVODx+9zTpHsa37z7oIsAUWy9jeeF+ek+gtCYGg5uuUGCL+vk5FMkg+kK
AZVFrZrPXTjMxL509W8P5N3sbS0irlUadoV5ii9jeoiSrDr+ErFT85sybaiWP4z5
ZIpQlNqm92MEYe2mBrcYLcAQuRWO1qKC8hnI06RlnAGHeuLLMvFV81T0aOv9CyOQ
3Znh9eQ0xEO/9Y1Yh1h14gY02ztPD2rkieEzxUDp8ILCGiJ5RxaIHHLq4wGq5MHy
0qABuK40zJd5Cw789WCvUbQHHTUTYFoQpWo7UkI9xiB3seHEEn03hYFHEVzIJj38
XW7blsRa5Nvi3kk99OXFl2MRLG6Ju5cARVuy/IQ2PlXSvTA12tWGCmPr1hU3l6M3
5VIFgxMu4RP0JQor0USeBHHuR6QGgMGh85rNGqQ+DDIahIV8wlskcn89LUpOMYHh
djtYJ3loYxyfXSkjgVVIjiztzXwTay11TEb2K3vozGVCZG3yp5AWcKkv1Dp0qvqg
6zVt6l4GaEpMChhysoCTGIh5rZnN0CQGmV7VIvn/slsEVOublAIIQYGLs3GBVYJS
nGIHiAxaZ2o8OgtFdGvAqa8FdoqNH7PBipbtJErbeBwCgbfPgn/xoNbbIQP0c2Va
7iH+bzSSfEsZSJSrBT/Il8uEZvZG/eRYIsTfi6RYeHZr1KNPUlvUKnt1SljcG5YI
ZFnwEUUepPA3Zvzv/w5LesMgoH1wvKs6Uv9fEWt2T32Gvd88bk8q7RpNTZicS1ia
iG3XVn9Q1zDZgCkcsfgVH631MJRMVdd14i6Pl/7qu6x4BADD1CGb4YU5A0yVYmfq
Ifn2MSgrF0n4wgd1p/hz345s6DR904y4kAK/Q5oLGCLgaqW56MsDT0uGkjpzUQCo
sl+So/PDJCSxeU/QEEUhADtuv/IeWAJwZESLk3tP2UJ/V13x4l6ihtzBi+/buhUn
ZF5ye7DRxtm8++qECk5N8GgsWUeq2Qjb3/KK2yvhYsRO7RxaVsFV6suPMv9YAjee
r8VQyf3FBZ7EQxR9ZuMrjkHnW8pFSe5ikvBorNO5VD6BjnBBFfrx4dqrMW32ngrW
Hm8Z+//1GWIGi9BKygVwitoLVP19KY6mCj+vuVHW7UtPk8LuhJC9VJ6Gtlg9Y3p8
VEBkOF3v0Q1hF6Krp8NA8sQ52Z2vjjVnFbWHJ8NNm9XrlBBAav/LfMur+Di0/j4i
nSdAB8CC/Cp1WZvCZHC26x6EUP1Gq53sV5BNsmltCTlU2bTpsNfimN9+UaCM+3K5
brJE/q3TY7q+N9dgikkz3hgbxC61qwyVgndy7/RS0/g9wgoZBxdAzz+j5l3V9yby
U2MU9wQ9endsFy2tdpp6wXC3vxSWYyYraoFQtAGuM4PrtBINbqCA50oldlm1TVuN
jnTlSO9y07shEOtnBDdFcyn1rbRTcs0uPM5qC5yliRzJ8mkCGmIEBeuL0s8f0vo2
au7pDwsGb07dMXUrv+ZeQYuxIkeXe9Bd/CJP+voJEnkce/ld3mP9VCC/1iNhrQrM
AAXQYsGgbOOLj04WdYcYBosuvH8cG0L84+8HKtk7q2PAInpmUKpSUUenOp92MGov
uPOPmI1dNtBgtpPxgSZPyTMwA0qTSyfxlwc39eFMa4yvn3DsOTUtCghnT69rSGiv
vfL7Z5T5Ra3m8wYvukTGpSBAyuQPOEwEjHbsxN05fGXzixlCJuBVbQWj1xhq4fbI
xdwbsWZQjVB3FcoYXbSfiZA4QMyMcz8jauoEeu7XgAqp1dtL/JA/0IFlaAha358d
KBFCqw9bkoAzWtUzyNMBigbZsqMRvDR0oA2nHZ01b1ZEeZ79iRKKAvEfYvkbVX1o
AELAVitBCQwHsUHZKDLFLuelV0KVi4Udx9IeVqB8hzfShFfIDw1EvGVz6wAWMzov
xhTXg6cUEKRMGeY6CUnC5cqo26GyUIBtwjlvEKbz8MnCSHj2AxxiE7VxkDviDbr3
uuCBrd3Ci5md3fv0rcNOXAqL9EXKVWgHxICfs26c6ZJJ//n46mR2Ow5smQtk2CdN
/5wwXFlDeNCe04a+6NuSnKqXeTpdyjy6k42pK/le6tYgA6YbjL0SzdlANc5zXon8
akN1rK2t9jEaAbN4m4tKNtloIqB1u1jO3kbYclgOWirQFOkP5zWM7VaMROfoMwWI
IW1r2nStbuvmVjfvjKbx/qaPUcaHBw9i8u5gTcUJO1vCKzlk6TN4jfPTNSG1nyxB
hLTsHIfDDyM+Q+mqALkZFzResBuKuX5LEKcyCjK1zw1ir+oP45n+/Ga3pz1q9Qzo
j1hYXDfbCTm6hGVjicKNHzOtbksDKt93R9u6zt5txN688OBdgoqlW038JytEGcZL
pP8yHWRBOiVt+bwZBSiEKDFWEqwBf/sl+IO2SbrcRXk+x2XiBWrbl1DKVV+aPS5b
E0v/WsK1Q6P6wFpu4w1tm/ijGflUdlRXW1BauS03NotUYQocY9D4o2M4EYwvk3nT
jbBfvabn7ZFmKxwKoXcJ8IBDGS9z/o3h3rtiCLfkVaBKmEkF6CRk4aENvqUIIMD4
Z1dQv8IW9W3lFHkn5DxKIlkTQ6qO9RKnLPFZzwqiVwr2Qv/X9U58DsqrdXy88Y9O
2whalODs0wqiQBPJv2WpzSrzouSHpkj+c+jYYz1EBjmTtPT3+5prjtMPz6+vQjik
AQiP8q0dC+tz9+FEYnl3piSXDdKnJFAeleycq80vR9XJ31jIp+B7abzFqCJTX3uR
pY1NjwrxjK/1/kgrClYvNGVqTx8nwKRiEjjNhZr2bP++TLeUioBiEaQh2IwxwZLj
pszGOAKO7aeOxqF462rcIjU2c+opUifJc8EDO2j1deS+rVGD1ec2ZhjVm8jvwKiK
AY8BPzLL81BcKR2TXvjCE56/qoJgzYU5U1X0Sl12FRCLfuK8ot1fwYPQNJmP3Trt
D9y6bPvMQt+Xt4EkToAwcfdknqGY6uZlqwyGU2fbY/VrjOOZHZw6D+gaI2AC2zsi
lYfOF8UeRTk6xMZgoK2EM5tDHlsUfKbSZ+6HF9re5BurERO8deM2PtrFVKrrj92N
kW5xUGbooyQkjtjkGP/4agZBlOT1GTeUA30gLsKeDUDvRe819auvXsPYCKI9SKXA
pN753+/RV+gQfoeFh0Kzvfs3tKxbvEspNjLEAhVQwGGa2XSY3uKbC9SErXsX3SpB
x2l/4gcL9x2wQnkCovrZJW/WClsO5aRadPCpsbFIRDtCy9i7NLlH5r5fRm6N00gC
c1U5IODI1ocybLH25pC9ELqDpFKQLWcnSjPuFbZbO6Yt2maLH5ubMvMipLjUI5rC
rhpkFe2SInWGNWwTDgJfsW6JoBYiF3QiDI3aqklzfOB0Ulws8hnwSF4POm98N4XV
kZxj78gh46RkUgaiM5Af2q4qnaodTCcEoEwc7x9uSEzscEVjQ/IKh97j0wWOq7R6
Pmpb6Yrk54L3FroBRNd1yFQvmTZBUpektlngKxBSJPD0uwzAPim/RMwWJ5xpoDuN
0f3+/EBvBZAPdfC47/p2Lw==
`pragma protect end_protected
