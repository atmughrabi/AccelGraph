// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Tgu0FY5Z41kXDl0Im+Q6lHTyIMVrLgQwFyIHKtH+ufl0hzPr//Fgdzo605eG9V7j
dGBebve9kWd/DrrBtilIS5eBOqwuasZvdKR5eMViv1LmlDTWTQa9QJ1Ug4VToieQ
SWaQF9Z2uUzg/tnEd6Yz/GU2b4jgGtLLkpgIOBTmv90=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29920)
fyqn2tiH8QH93bXayAPEOaNC2+kHukadKaqjZTfpgVqmklFyFSjuYqgPwnBWsEVB
iQJE/EmEU8HH5d85xO4iNd7oEwxeB0Q/ud5WqEVcq9OVWLSoioOfI1123KYNRySn
QUZIZQbCXwSWOoPFwbTUHIrLpCFzPrTPTbaJspAn+ktqltFwbPryHVldq9Q970iD
rAK76saQH0dUD40rdt+t6n3BzFysTpmY/8MPgLq0WJTiEUdeBy/ldFFuYaI17RVP
ulgIYfcti/JgNf+C7egUwIWvjCaMwN5zZef16BtimCagWav8K3hW6jR/MEjTg0lL
J+tKmTYcTEDtcFEbX//z7qXPSV4TpWwt9MqBbQ0ZKygcC8IZ0jNpb7dK7JGQuBGb
1p1XMVGVyzsqYq4OdGNhGvpDYSYUV7p+5/F7CPZEwM4i2tqOF85k0JQ2VDoNkM2c
ITRyL/8bmXWxmuqmw4FfiYEXq+0tve8hDtfFtbQ9X2h+OyF42AR3ET+dttinMw8J
OCTQBd/PsCuKmkBN6+sdonMtrhxS6aNguJldMuCmRQPislykYMsqahVtqXaJsuM1
rHnK+LRyN22mBJFRUkfrrRFcq4c/HTbjgSGjqwwIrB2gyAQIMw5FK1uWwAdDp6kf
8u3e1wamlscQMehr3Onu98grU1QB3uAAfUtZDNx8WNiE1IDM+O3hQMgdxmxt0B/X
tp+bh8yaSf5oCnuVnmmfsngkyzLjPzGVbXtAFrl1R9GOfom9Vu/ljk/obHtMmmN+
zu7j6ieTh+J8fRbuHEDBs+FMhMYnDPxJCT/qbOMeN3hoTdeE4tnpAYpRlEki/GpP
H7EAAbSMCnwQNdVZ/SUqdnfno2Tr3uFi3prhnRDyBaaBVbO3+/JKcKOs84VTESbw
tu783Krb/OQ74fOrdeP6NPH1bazV8PzoCXi9wiBFXFRTGzfivId4X+2GDEMN5Vdk
hB765VYv4aI4EyNdkNt1uBhzA5VwfjDYD0Up21/mfsluO7D1hPZ0aQFQB6HgoYDq
L4KSWMT739iHK4axLVwbVGdc864LkaJxpihn0bUI7WrQ9IH1V/UJoR8VMXYl2PwF
if7OUeVZcgQn7tlIsJWxfoFIiJV8t50KaA6Wp+AzVcTUcfgAB7Itr2mb0LOyiB/D
g6uvSaN+kuef2CSs/3mbknXl8SkFR5ElqSXFYdUI8O8snOx3yXJn0OZl9kQJnsI0
0BE7CwqdlJBXZt5weK4h5nUnio2z7hjqVJBeEiXfC+XAE54pdsX9s275glVNyo8m
hAIPSjt4od5u6yyTVvbecMbjgiZMt2oXcuOn+7KRGpsAj/+CQ/BkHgufSBmY9AVO
5o+yG+vpa+srBrXjq0sobnmbutGL93LpkFKj73QnASHTJMHNLCvGsgQZr+wq0v3m
4tsIbDAAoBTosQdyWKjRTsXHbfu0JIUGFNmUlI3S3M2qrRlQukV/QsBjdHW3QZdF
2Ri7CfSBliWOkVYCjoHXWLJ4RsWllMU1SlZMwyPa+QgYauFW5WdjVyrjpe59d7gj
lP4BIzMCvf1mmbxCpxecgOD1ds3QWGN6eA5d4BG8rTHCoSDrVE0ZAvnBCswehAt3
raaUG6zmbqwBWgSBsRJ5vRiZQw3nWAUG0GnfGJ0jNqk3cBBxnmXN52pzQ942NSUV
CRqLWj+jv0GLitCp+JfFRYxum3oev76sAU45LNsxqXIR2ZAFYkcCQAe5uW1WzQxt
SyN1hA/xb0DkU3WwBVyYR0kHhcsjOXCZcKjW+ksr1tjJ80tm13vtlmuMv51wmk2Y
f0wBE0j7J9YXjA5ZzBHVDk8J9WQHEHg1lfqc1bi5NTD6oCoDnxgc7hwVV1I+3DwP
LZl4+RZn8Y4Bs5k68eMEc4eKVVIVr8FBzGEo7CVNRkBzY6p54oMKlkBf6CiaQ9ZS
iEXXXY/XKGIHBb+zVmL2UYa/ERSH/8yc2CtjKfxT98pNb0b9BM4z7tkNSi76EeDb
gPmlh6hbRBLe7qSibwKc3s4uY0LtBMnmcN4hf2atnd4nMHiMJHdnJKN4+nDiCYis
Kkc17uBI4GT4+cfEqSiyYHA1nIkZeDcB01LQ7/PSVQjL1McRHVWQhjneOt7i2BGe
+qk6pCA3QqDswnasbuY9Uw6hBJrnAsJ0QPypkD7Eu18tBdE32TzRBHYTmh0+CH2o
13YGm6KWxtUUA33/eltb59QduDvIySD4nsi4jCexhNdvnWrdhxWmhrFNoPFbQwth
jMwBE0jNjAgnXd6or9RPWeZd2RLOKGd4g5yt85ZOqXZY5MrBiQueDw6I7yQyx25R
GyAnAmagGa5Bzn7Znfa3ZQqt3YSHCzJxBf8z/SjASXa6ZH32/26uboogMvNzc07f
FfO5rBg9lwPxuwr7V8JUAYwJarAIKcJgLW40jrusMglhBi/+Or9lXlxUj5iRJnAC
CcB+kg3N0rN2m1a8+IEa8LyuCJLKod+2Fn6jTsoew1x4PjxUsVB1XPfJbt5vLaxZ
FX/ELVK6RcKMlaTVdlTULT6UoE91u9m7G7+VkgLk8KaeboNARAX6hJSJmySBN1kC
UI0QkoXbTAvUVY0Dmt39Xd6haDHtfe1/+70N+8uU+Jy6yrp0HmHZlk4gON3ffPR1
kbuB0r/ha6DuCFt9is7JQRzkhZG61dEXTSLE8hXh7Aq8cWkIsmQMnIDERIuAaTE0
YVI4TD+G2/TqY+2fcF6IfiXzctgF5c0vqKiBfllWH6QKudSY7hnTAfEmFznikary
sF2HI1t3qEp4RgmMq2Y2CbWxfzh5YGp/mzeEAaQW1MC7vzeafLpeSGkGd87F+cNZ
sezwh9w0TWrN/PtMUPw9uGDr2F45JVVG6lWcTfD/lNdHZ21JYmYb9n53f7g74NxN
YZgXQysGJaN//jEWNct79m5X0LqDTcjx+2VvHdhbCryE5vhDhQt6tZu3IX+NZVei
9EnBk9BuJhAFhrMa8N4hMCQCCTyWM4MeuxNfuuM77wGavPnKPWr8uTIH18MVg5dk
HBo0/uh8g8nzNdygX51octgTyF3CkbRdFPk9lSFKTNAzr02f3VEkSvCPNh26Frbg
dGUNifJWi/WR8GoAFfqlc6/YpLfck9vyEiMng6NYY/XviLgZd+r1mMCnflR4IBGe
LCO92Qr/TU/E8juHVGSwzRTlQwLR7IuBAVGpkGvqSL/d+bp85rcuBQd/gIMWB3B7
Bh0THxNgddIveF8TKtHTMTvHvlfWMMENtiXZnPnmqFrTePYMPmEVjdPInhtR9ard
G5d+e39wATl/saR7vojrBfXF6ZMIPdWSBL0e3vYhxBfQJrhhgVmbZEPGOGy7Tbo0
nZqdFwES4fd+yIhbAvupjKCXaxDkJNQvfw4NfFI36Ddvd0cj48eXCn6UFdTtZIB0
Sm62suVY7Q2ClydVE78Z+ifpSStQCqRR/uTiZxIjTLqYgnZe9gb/CuEsukGnmTBc
oNJrh4rO2KQX4JXDnvEd44mJyfVMy5Db7fUKsIreJBJgG4a1fyi6Jghv311KG+R0
GeNAtoDhys8f+Jjg/gugbwqwYKoA5xvTZehY4x2laXuIc4LlWlg8jLPKLSsvatXZ
x/KkCXr+k+67jDVY+pzPlbPPGojXc5JS3GGvXmrAZSZk6pxatnB5s1zbg6hPZ82M
wHpfMWJeTKBC0Nq0kBHoIjC7NFQKHELL7Uu5XhNM/Rj+1Ct43EZGxF+qUe2ZyeGA
L2vryyAY9UbiJBBXuAtcN6PY5OP5QVEpaRHQjXEVYMxgetrxml8PUTyekgmx5gK7
AowPC3+zs9JgSEIlGb3qWqzyDRTqldayLgiG4/kAX4blKru+8gR7q0n4kCPVe8o8
UrAg+QYrqzjhr5V+iVWejqSNAVr+Rvknuep+7FTRB8kgM+dTOmVPFJkXjgR8wEDA
GtTVSi9ao1LqhrxAHruYdwMtIJim9Im+ifmYSykQeuL2aR6GhijnEUfHwTpRD9/h
yaNN5gl+khk3ZBhmMdARYmpv4FaKS7qq5sjVKSWciI3t1deg5plksIt76RYotjp3
ZFckXWzd92b5EY0f9HVyFWplmKNkDi7PTHKLYf9OpSBSSZRnpfn2JEhgr0ttirRD
rApYDzgaZ6zXRtc5amw93si5OkVJBKIzNiByaCFn/l7Z2+sgTRPVigyKmAOzMOkW
vOtCrzQ00x962eGqr/m11FM/8smGo27lrBFMTtss9w2M/v2XWPlXYeCXylsYPfbs
B9C0z08+z2TGGadFbk2hGK8mSPiMDyr0OQMYAguO6FAVTd9SSdGrpibmkaNhanNd
NchpuIqHRV2qwmrVUts/0UIwMNVsQ3OryGM977r7Fyrh2Km8yZbJhWjb76jnghD0
bgXU7tGYfhXe5Esw28+IW2fqIUTZs5nz/KhPWyugIRHjNtX6ab9hEZEzzW+sssgm
0xozgBrT6vAQdoUVt1E7Ki742isQQ1D2WCEALFrl5ytewcA711NdNJoQGWq77pFY
YOegr6uM9JtlACMFj5Fvt0vyqvZ0yLW/BFM4hbyZgNxJBFDLjzetdJSNRPV2Gkhm
9PhNbzIbeMOXPIwMvXVMga+wqW8G+A6vjE+qVWQbnu/E0kCD6Lu3CaekLBNnowDA
Vcw4NDBn8nKYGLF9DGAEV99mS7aHjtJPIueODYjiW3hvsafyvlgZm+H3sSgAEfy1
fY6qwlCc2twR+Ihfmb9PXqUIBYvXdJ3J5LZAbpP7npFFp0FdQA6H8131qnokeDL1
x1MopvZUXoxqrLIj51yI1TYidVKsb8NBmFASflH+6uSOwwi6Y98btRM9juJc/we1
OJu4G4YVX4MBsTWGS69AC2RYEAmLS9nWMgv3Xxuwq4sMjJ+6iuOW62yhPcdEgLum
DaNIPj+Xqm57AD24alN4mfECXrDR55wfl77fUuTLTldDnehFXnW8lPYR0PyJyib6
0PfYOTyw7MtAoqExW2bd4pm4mR1es1Gaqw0rstGepTUHnsnzdDp4UM0voGO1Cg4v
2j+DsBFyvX7TPZPt5mVXuJF9Pv5Y9gIL9vDjUv5C0utQKAP295k7gH66AVf43WWw
o9Da7yfAcZ/3FVFnmukuPZBgSGNwaIy2yh+1jDt319qFSpA+fNaJsx6kbgg/eEcW
sLv9F4R4bYLFz9GuFoFkEG96iNpOQlv0AbuP0OrJC0ZWqhJHl7k3wpgDOoLov7bN
ZkrMICPuxgJ7P1McAYVWeC/U8bcK0Vm1KAIVccZtKk7R+4RxxI/EZoe5IwT7Tsad
CuQlVKOp2kGELhk8f+C3dHZIKHa5T0xJHrZMRapp5qQ3rJd/kC39zDkAJnkJNeMN
5dVgRa4QTUOtHCaQfdX0iD0HybEVcSmPchcmwBnRNcr8UDxcFbpplQUu22jn8P9S
xOudJZqieE6smelnET92YfW9BbFADMcAdvFO7wMFYs0t+3MZSH/5PPBWieX9Yu87
lQIn5T/OwYZ28rmXDeg5DgkGcvy9uKORW2VdCST9enpJyQTUfr4GwId6hzxJ3cvQ
MSmhKGqlaZ6SEsSntqT6iCkhYzjb0uJWBE5I0oR9QBCav1Xxj8IuKEU5cfunxgKZ
ydKY0YONFHW48aGpsLWP9SfULaY7YeKF7HtcQfav7Rptvz/GjN8EZrzsSlPE4YSi
1MBwiBV7PFnhcsCGB798Anq1bkKtY0wNdap9SDXVRYPS9AlnlMjuDMOH/5dealUj
l0bNxdwBggZAvoQSrdvBpBYEw6k7SajypBo+KaRubN/Bxq8E1R8maPqIjthcSMI2
A6fmHG63WHODuuY3GiLaxv+DLWgNUaOSmLd8TYPce7efj6R6QLM0g5gdr918vPjJ
N53x7Cn4ZkKIvAaHpORwcj2PkD1iraIHPFclyKsf1LZ5o5rx9PIYjOzsaFlnX2d9
wQ8lp+xBHCoeTPFRHa0k3dTCB0rfgPx9vDMDAvduin6UR1ejUh9trb7OSDyLjXCV
tyq0CC3Dm+4W4zCSEGJ4AevlHJBbW5/a4y71XLS76LsUKbWdLxnrExtYa4oiT7Lu
XgK7UFUtL08y9dwjwzJZI+fkJmAzcBBk+Xxxc9J7VRpXwwMaaL1F5HNZn+XQ+1R0
MmU5zEoah90X4zmLGMaecx/NFxgPnAKrY4mFvQfOMfF25m8JMWTL5t/JBZ02tMEj
Azg1WyHUQIlN5hIEcog78so6weSRMUylh+H0238miFqNh9fz+YxSXgdNjC9RmFr1
q8KYmFnN6B+4Gf0U3ZvETvpaeyAKg2H8k4EqkepMo4+fjTejxy9HNjX9DdnjtcU1
l9ZZwSEOIkWdQUjrOi/IxNxsGuUGbljjiXucRemzvF7vsJL8/r04P9A2wr67Ayrn
mGfiM8PW/wWrfqXGKSP6o1xv93qI+GcQFOKsp8FudDVHl34sSxPOJV9m7sV67+P0
fkO1t3DUVrZ5xjrLHh7YHtMNJLayA0C6Xw2nZycu0Uqk1DbhPRE+tNuGiV4MEkEa
cJ9ijb+6XbTYzk6wsJuFWiy8nq63r6GMyNbDq2kU/+bYcTps3qqjKHxB+WBOEG5J
wfizfuc3JpomFU49Hpad/qzrW7yj+b6gJFwJk1inm67jdS7i3vVQceCsAA7/kJuI
Dnhx/r/a6+LEctXQPMdAHEv1+EZw6ItbhQLeJZlh/u/P+NWjhpzJ9vaTkNsLhnVQ
qLHkLip4TqwRxF3PzzcmD9glUcdsGcbIK523aMHG/QqE4NU0qdJYytn9Zo41p697
fd41krN8xOxO2lnSPL8Zlk5NOV6ipHlTGXZba/rKoYFhFqIG7PoJoKofnNYKV+Vo
LA3vBneLkn0fYaLJ+G4vUNrKf8yff3UAKQZLFTSqVuXHtiJcx0coqpSllvB6OolW
f3HV3t9nmROVb5iial8Fn+AJOS5/gQsnZHy9AsOaBjj/+mi0SPYJPpY6JBU62a8d
dZYMMIuacY0jiL/GDpOn3PBhnMQXlZ/DV9xqT6P45ep8o+FYwOyt7IjJDi0gaamf
Gg7oJhY3Fh2r671NZQJetKXxgz5a5mj6EEaTtCkXllfQVb1FcjEWrqj/VARvPKGG
8qnCldKsMdtJd5KoletUyB7Z1TUZjOPNN2yMCXdzA+PqWsC+FDH0Ru0I32pRqA7w
2TwFzzF23LoMIzeX96rlH/qUgzE/KrN9qSI9W6DybyNidckolThiNdJFImNS7O7O
5e+9aKuHSlqGaRaTNfscj8Xt9st843M8ztqD0KjG9msuUzjhPOrN1lHNmlEzlYP9
hFEPKHBxSSR2JNq84Ab5VrNB8o2FXHNnFJmv2Xapghb8U+sleHU2FRDttYLxCLMG
r7RxW21RJDeN+OQf2mZnvwICUvp0dFXfXgjXo78J09e08ugik1LoDciaOID5N6ZL
sK95appKbvJXrUjzQunZs6ZtXsIYW0Bp61+GiFz59hThGc9HoVUPCG9NgrEZES++
dOZM20qxE8fjTiHSUVA47YNx0Y8AJ5f8n5H+LcZRNAZi5obeF+9xTHygJNdUlWm3
SV2o1n4vLTsf58XU6BCzeo0cVV4Cne/Nk4T1dY3IKcrMO8vBI6IM0rCEzlAVPfSx
a8nz0s98qgVnL87DnY1eMyqvu6IX5V5EUp6NtNMJgUIJBd7DlM4J5Xe1G7j4ji0e
xl5DByF3u2Fyd5HRxhnJCWKGIADOkAcOcoObi9yfkDyeE8opiw1ZjobdEBCs1Rbr
CRMH1CMxUp9VwxFBJ0SRbaCXnJV5SxcrpX+5oWFVCJMOfY6yLT6RA0WcpbVwXGKv
sEyXtiZuQbxekIvSP6/1uv88Lum4SqyzjTqehJ8UILrqAIaSIayPPk5PkPLsDuN2
qxh2ziHTFi7cuVYgOpMdzawvLaIudNdifI0lhp7CE9OyLKSAxAAI4ruCkux3bdwy
XVJlZ1fsJX3DHGygdJyIlP2GTlB6eT41Fs7z2uEgwmMRFiJx4KRqcKsZGoJbRZUf
o59pj0hBrmIwqwrVRiUlhr1Jfm1j2eO0JWYz63OApXGqoUbnpC3p9CmcuelH9/nV
Q8l2BaP6b3hm+VdkTy/3ydJUmEmKg3l1B4UCsKpLxyftDhDb77OT4J5F7xWFEkLv
dyxAguDzpLXqlJklE00EDHA6pP5joKR5mfKgghPj1DNqJ4p0+6xmYHmJLSmSgF/X
kz4H1/Rtyxl+bpuX2NOQl5usu3v6n8wG6e41pQ8a0Iz54IKknSovoLASas6cxk8Q
7vfCP2uB3QaJRVIl4Qshc3m1XbnnlRUnZT7ScDiYUzOAJLM8bRBneus3nrDlRZ5n
z3KSbCNcodCqnW1OtE8S61J3t6qLQH1YdlFcRsi/TKXdX7N8lOnnRGT7ngJBxSiw
p8dIHHq5j/HGUBRaWqsJv0Ej6dKG5s89q+cQ91ggXAtZJXHAG3OMaiz/QjS+KB5R
klMoMsRewlkqsrZyAaU6XovmlTdOMztB5/LrZxpjJtcP0+dGjwJE37+Eq/h9G4yN
enGdNBhY/0UbANzxQhJHbR9JURhnNCb2aT/ZimBN3Oph0VK4wEyQof7EKHEqLgGA
OiLOFn9K/CuPN5g7TojS3EaqM/bdjEP/ZVaxOthOlSJJtuMdJX9186QC+IXXp0k8
6elYYngcKLQhS6Uk/WFFsf9ytYaZ6Y+DdkVIBtAkNdFkkZBd/VtYjrg4Wr2/X9k9
xVoLh+cKJHZQnm0oE0HNi+JQ22w7D2wmjqDFQH0aSrA6x6PwTnA/BU1vR1cbgNLC
iWdMqU5NpA3NhHm9gtH21pFoPDDGZjf68N8dYvmqs10ERf8dnvheDjaNqh0ESxsV
5AS0D5VYknvt/6VPzEyao2FxNZFfpCNRoVm/X0p3lqN/NBOrb2eLsN59RBO5dlPh
vTcDKkFYT6yb5WgEID0iGdlU6rBPg4QxN+RG86mLA8r/8unISSKU0A4nCKfBeqL/
IWVfpdZWdK44RuEu3g4RzMpm2061GnFUfX2IGYVF2ZhYRV/WZIuSjOQtiP3aSS9V
VH5bey16Jcnoab1DW2/NgWgNUzQ2+79Bh5uYTXsAyIWWHbDnGfsGlBjz5vgkrfHt
nsR0YJgdjfIQ2i8cNE22BDcnKAL1R+S8yZvFAub9CVF30iJQuiibeHYaECTAna+K
Rq5qkfkmDYwmcMsRTP3nzf5MhwtZiY0Nr4w2g31aCeDPGjs4qb24NRfrTtg+V+93
3kKmoEFdbO6gVTQw0KfrVvswLKA2R0w9dlTx4HIztwhO6ipISA5tdQbdPklO/kCD
dI40aOQV0ML4Q/jaBQ/jlrP+02y1orfNnYU2QHf21cm/vOlytIjWAv+S9xepgE2W
qYxCItuddm56pXOZGc9duD6Xq+TuVt4xuRM1JHDG3SX6+2LoidqWDMmX/tgT/9GN
3iqHEODm3vdSpEKOCgAxM94x1dm2qtmnFUrFR8kXlij5ivTV/71ivVERukvx4f0O
EQ4MzAu5CxLWJifiXAy10dxBqe8OTWz32MMaz8DCoE5TCZsDWTuL1n1pOb303Mui
DlcaJWsRjJL5ohevVwM8jtIYsHkx/PMxf/1CVoGbhTX4/h6XE4JShvY/KZysergt
poGjZs/FqiIhP4IKjahifXOB8w5w47olzqPbeKIeEwM6I4wusMchC6ke9wKl3XFD
2DHd8xUzS3sn6x1gAZVLRoS+fXi+5hZhbfEHP0SIcKc8oGbaqhiQyhxZhGESO8YN
DVD3q2Ehc9v/Cc9nuRo3wYsv9gnh3I3UzQppQnmcS0v6LXGaCdNZMNUGjbaTDIok
Gschum+uqfXk8Ofg/LZRAKqjLI5Xod7Qmf2fJ+snPZb0kYiMq9jdVNVw62mWDokQ
jY2upVuPFR/03OyN6voOH8VXddNo/2dsPYPMtPny1RD/gLV0HMSW9l9O6F8u4QI3
EXWVPNseV+Ki6eyTrAaqGc+9jIyROlivc/DpJtZsX0Ku22+F51gnAhCaAQYaOVjK
TTDFKqCu1J2fVpM2StoUD16BVefCAqUUMp6vm4XMrERxD/pJu3m33WzK4oHTJ8Op
mjgLjHI21ofntc5GCKrJmI0E05f+K0Ew4H6U4ZAcqAaXXhrfyawQOWvKxYzG7GsF
lfUzLHLBJXmo/67E2nkTB2o/xU7q4juF7FFHY3c+B7APcfW9zp7o7Bq31FMIk1Tk
/EoSUHCRSaV9jpRRgM/PPFuwoBMzU4N5Oia6Q9NaXZW86gozC56Y/7eVeEVbsnbM
g5H5UhcJLYfXHMlBclr2GiCvalyK60aXoY9iYkkIv5zGnQqjhL5xJDSavYp2U9po
oebiQqGCflXyX5u0ORaHjQCdw3msIn2++sjzSfUApS2G3Bl8+O12lXxUC8aKoULJ
pMuRoWWopdIhRT/qB4Ut6AX/IHGosXzcYRe9QWjp4IgTNnFgRenJ4I6dSuuvnAW1
/pBCV1tEM3GCUFIjMxN7HHIEUY3hZw5O7R4ioNDFMBxlQm1c7h2mPkJG6FdShGLB
tBgcLqqd4NdIw6KnaDYnUhh0Kh746EqxMzI2vth+czCTzrnbfgmFn6Res4SVyoko
YnQsKd5f7FsVOI1xK5zTii45fcrvucyVLT5EYcY00cRgz7TIGX7v7rQK3vBUc9fU
NxlrO/z4mqDrJxC5xz+1Yabaz48mpBu/qKEqxOMt+gju89LFreQf3RlTHcu+RDWz
xfmm4mw+YNd08Eld7aeiLwyC6pjkx9w8P2y1iPkLmbCLpdHmCCI+nTLmYCdl73sd
uN52Owb/Uit7JmTwQcU/8YOCPL8SObAEZe3X4f5Py3Cn/D+zBos582hQjJbHUKqG
U/zAjKLllXnVKA08bRXtfzflKxA6IN384MzEA/JlQ0nyTfEPB7JzC1dhrOgxzVdX
zBN+hcdhlqfxHJDdbgSs6KNH1hcBM8u784laqwC0Vmn8numf8RT6sIf82dlEbXlU
9AM7LdO2D2U9JclmKevweFUyb8OO6Af9i6oTKzBvxpoiSU3HVK57GLq8JeukoYds
DkmjE/AR2XzaM1IjpaGv0/ZdZkEguHtylZlTlNot14Oeqa83zaQCpIBlF80cuJbw
Kkr598jcipDrQYA8qZH+XVlaMHqpiFera75d1LacQr5SIoAInkL2XBt4886unAGo
g0u43pMI+mC6WcPX1O/gEEoEE6gOTiwutWL/7EapBIyJ33r+kgXFJBLHYK+muegK
GCMKwQWlpSE2WJhK87wsIzUndMaCpTkXbVJJQ/HbAnWfhbsHA2r06I18OqX1Nn7+
NiyuVhiNwUnDZ8ntOz0x/Qp9nCYP/zwtsn2lRtQawmsLx3C+azJSpqWChLUIUgOm
PvtuVhFWcjyp93dpRE5Q5R/eDEPUn0J5ZCGFPyprsfJfqRm/2XXFbWf+/UV9MgyC
zwDYqJHk9QZnugNz8xKxkXdBFDRc3IznsCw8reQ+qA5wOugO0pxEJKQ7YMyDApX1
kvUBDlesKTWxcmF+zZlsQn5jHm7B6eeriBsZ9EINGiBIIsQMA4cddmYmFO+3LDjT
fS7hVVBRgnRdoF4jGuRLGlMA3wWW2wfMn6Lvbf6dUh5XnukrI+c/AQ0uAMR9EOqK
XgGthHk7kdsc41DDBcd6CpfCiInI2ZHzFhxgei3oy9wlUqPULWgmYConZEGbTSXu
RLrRSRAc9G0kiukBmBZsP/Vnz08Fqi9aJfqU06XZjBFoS2GjHOYuikBFegCvvJ9t
0VYfXDVxv9/N7YS9bDBt+MEhqAXshze2pKAk3AnH92NL7Gpkb4SF/BG4+tOjJf54
73rxz1SeDTBQhTZOv8cZNh2YXaa2/kxeddRIC6Md8rYRYB3X5LmlmXGm9n5bgjS7
Q4NK6xolKJrqtIvvBNxk1APkbz3zfJvas9pWG4etmjAO5tGAIgfmWvzvsiZkbdEt
zvFk/75vbLq2xdLEudxXyqwIiC5nJdDm8psxNajaMTXYU6SrMv1Z2I4rNg7kjJWj
Hm6q4QK4I3wCMB5LTqK2HA+sX/bqViOmZBqVcpVuEL8wYDAkzkOsyV/e0vd1v3Lj
2BtnvNtxMI/juiFmlEEz/0ZgIAFjwK/6+cBdcWmQHBmAjiAC8714/lf1jTEW81uw
WQb8MwZ4q51QQkkZz482LInOa+oEYq3PzFIHyvAgGz7xaCim40DJ2icuNhIwDit4
jDoO9rnVLjLYlQ2jhSsZAAkspWFcOfFU+pQV/46c+FdDF7wMWQ3q33KAS5uQP9j8
z/2TmjCdl1jR96S+40iTCGVHVg8CnZgWdFAUnYn7M4rVMr+oGeKaN+jZqdHTDTWR
zGVXxINMbEPi/f1eARjhUXwW6oOBgmg+8FnVzjVZ6Qk5va3KUmmlHtYy9WDoHdJk
E4KOMwQ6UAQDt2XOlbfq16UsTbVqB0UA2UcJwRAvzUgjcf42wAq1hDflWr7TzJPp
nevfVxUibwtI1j6OM2RENvKgFOEtOMetA2SDEjZpvQ2/Wn03UTUj5c01WKll3ulh
Y7mvehbAdNN8GtMAxXTM/8fr27zhqFLp2Hf9QLEan+UboRpNLVLt36ZtzUT3AsIq
hPHRberRjiiTvlzVJFL++gvzGU7O5Y4USpFFxg39qvj9VdoPWIDIp0RuqGY9OYPb
7H1B2yJM8l/3TTVcaorAwHIQfLnELz4RBH8yJAmf1qEC6AE3y09iCUp7sdn+Oyow
Ua1Gy6fJtgjNdcuEAEh9abYJyU8FpcTbzb0OOlMqXUFLeyrGWPgkZKdDkpqwiLT9
OwjBHxo4w/KAzOFyTswwTkzwldu5Ff3ZfAWH/2HvCmmJRrVkSCskHk+c9U+3/Ztj
JUnqy7sYGJWbAaGM4n+4/6NSrUIQ4mS0wQ4jBaLHH8xfDVlDkWy3AX1Q7z0b2VbZ
XsZ1L9O0JlINYcsF1AJm0UOSEeN5CaK1NLhIWdNKit7ATNa20qcigZ3HVYmVRVkQ
fIctIWfz86bOp7Z+mTQHlLmfeSwYNjikCV7OPVXGDGH81MJ6w12ym/TAvLL5sOLN
j24/0n/T49a2lN1oM1D0a2ULcEuXVsf8JGNiJIjj6LYlpo1c+b2/ZLYFo6yx8lL8
97e3rLCLHozQXXvphA7vLHnicxajCsjLikUk13aUkKsF0BO38rYyBSfDwKt7p2aY
vROwqf4QiA4LoMtQsMqqAwb9QGXwdiPgu+2HxzvdMgjfwjRJfb5gqdc83D45mO1c
DITWy+uStPUWXqa61AKz2NKJKkHqr+ZY8KO1BGiauZGVmACfc44KKKCPKpkJzJPE
dKckadczaX5GnY+cLXiyUwowImzI0zcLKE735sH8cj7YkX0Loi4MMnS4H+9vm3Qb
bnPYq2NeXUO7YSdR8ngn+PiByI7p+smVCNcj4XSPNNq/VPPPGXrOH4HUmw7EAanH
+hJCSAXT6xVa1VecZgOHB7sl5e+gq8ljOc3MJpJl4XUhc52DsqkGapU7KNauokqf
akN1FSXa4QELoZ+fR+4a6VrPRuvaS0sNu8oVQMgxvFpgEfVbGBxNV0PmvM4Yw6yB
EKiM/xClSAjWaz2ZjYtlFkVqlbDayVE+iFN7A1R+pPJhNyXeNAsmSLVW7sIJ3fI2
FU1w9tYLUmHcHcWu/RB7VJMni+t+Dg9hoHSkxQgZVING39g2ztiaraiiwn1d2Ffv
/3FlHEPI31v1fR355O91rLVYL6LZZKWEu4pny9funTFbxCq86vKl3SYcEW34f9Rg
S5qR6eYP8NNNwx+Vt8o56SY2T/d1WeE9ETIOu88j/fM5BRK+we2vYaBaiCK9dwt9
llzp/99laTjIZqQCJ64ZOqr/BHBl6EI/4+7rIrD97UBIEXRxltxVHpDRkEjjZwqF
xnNUhOgOtpe5r5ncMXOrvrFfkzqcaXTTNZngi1GZo04Ffd6D9ISen+CgnyN1yhWo
sTRTXzYtsNPzBzNO6LVEuIe73fStwH2pCuinulRkSTPBZctikOLmPzUmv8J0i8w3
MLjzSQH8wri+hMp5/viiN9p1NMGXeFgh8KbqftiSZZLy3KI/cdGi2hkAxY6gZxxE
VfHMEE8VbQ7UXMaD/ReuxFExc5fjkz1QkvLqb1ltkpftfLgxxvPo2DfV5nM4F8G2
YlrNnp6HK1UuIPcVS0q7IoyCWYFADftW41jMglpiOmmq3C/bLqrBKwc3TvG9/5Qe
GFbnfNm5nAbz0XMdPn9JWx3vp2Vj4jMmU+UNGcVLHnuz1y+VlHKfVixXhRmvMd17
zKAz3s7rW3VlTDi5t/fTpjv/fo4j56tWObMem7tXTqvErEqBHM8o2EbjTSol+FHC
6T8OrO6OLa+3W4YnVATGnSe2yn0R+Um6MVeBSdeg1KZ6SyL7g25cBIWaP/F9nLTd
656/vbPBWejcbOT8K6rp1Hb8Mzn4l7mFEE9wgSy4KQtudeYMmQQ7eP3MvqsaKjLm
omFpNM2TGTmUAeEzpBPWDsu5RlaO6vgl6YOgUsny9xxbpRooKpWkKo2y3DjtBVaV
B08Tn6SXiIvS0kU9Q6m6yHAGz3mUqzfr+KFrVxIUunxCPukPIbGY1hcNAV332XRA
+3QJcoamPcDGGBZIeCBXqW9nojJlapGBuPrD8yqeFLjFOoEV5/QdtV7v62JAfUra
f3DQlJhMsAThU4WAunf/ZHxj7b2mvziWEaaYhKUHjQvqy0nx0S3iK/f689V6iXaw
GcGz09vjAaElKKL+8Yf+W+FiWjIIiu64013nYXe3mGkZI/JLOL0dQaoT2++g14u5
q0Rydekupq9NadjPiIVpsnN99YFvbSrcziqAEXSDwQlp8xziNby5vimgjKAL3Vnr
NSYQo8AKmNlA2lRvB9xzoSYWdr0sUQ6/cKqq5qrJyGq6SoeCYniNSgutqLiozERS
pR415bHejLAVK9JBB5X8kc2niz3/xbD7DS+RxZT9Vi3akdFBravKYovuXJF5sapd
2xOlYHyo8utWkF5HwkE9g2DisGNt3FYJvkP4UvlYHyMfsKiU6D6pOU9PnCyIG/Ji
Y1HTKVNl5MqnOGJ76jv7xkfU5piLSNRqKl9GHOfviePaFRw3Xiuf4Tng+m9AM2sL
6adJ57CF+ZmXexhUmQKlpqwAn7OwUzwH3sTBkmlmdWthZo/q5pwBw74S/76vnccw
s7CjhLXSMzEmucfXC+rciu/MpsYkdNtPDXkGahu5/DDN9Ttbg/gJxxbajIlEwou7
E4NDRODLwD15RyOC0A0947g5XcrUEuLmvXLym6PszlmY3x3YLrlVSADuCC+kewkS
ExaqOid1PGPczXTRAIHZnzhrNOc9VlbWr1dWpSR8eXRVhxlRdd1VsgTIrDLMN80X
s2ipZcwYCt2jyFy3/Xljf0nQ5JGaNA7S7t7v5wqnFZIg/oWdR/a3rTN6R4XV/H2r
Wf3T+gWQKZfLxKgdder5S9sr6PLSr0ideNg+rvtDPUsv2aVxwWOxQUCZAKkFGBlJ
ngatjX4nXzEq/idvj9/pIab5zUF3FUMdKcPwIsz7ybnzRpTvEMU8ktJVAWeVxn/j
IQ5irb7uvJxRODYbwiNrGxC6zF2zGevCxyvTQl1ABkE2291msHumpOucuZ9aUAc/
o/bkKuzh5pUQ5/i5ZhO9OtXyfZgxQguYa0d5cWB0UkDT+ppeOVMhgEUT6QnxuJJl
WBpNXeCMPf5BF8xRCQA4bRgEIMlnTdtzSA0cte0ZKlsZh60FAvKUjXdUVxfjVyJ7
kezT02x1TTUw/oFcnCk7S25EWa9rThfOIqYRulf+B2WrESyRZyIQOFMLto+TfM9q
cl7Yv/EWMTK02/HrCMt3AplxU0kB9LXOjJnCD7DQiyvxx1QCf763ze7xZKgzMHBD
7hyM/cB3bZPRMWrUoZZGp8+PZuc0paoM91rveeKsAvzOxq06PNwzRvgGmTuHNoQd
e9bX0AZbavTgzursCLbhrvzEYuNYGm6qTxlItGVDG/GnNpTMqF0FP0SFIryhd0Zp
lfyR2p66RZs9l8V5TEMKOmTTAR0Pb+LIL+KxvUq9dK4NjfpuEebnAcIEjZNXWkNl
nPocgv3v0Dna2oSf6MUs4MlVVnX3VqlxXXBWNvQo0FkUzxIZQHowuHC2I8gbaGUr
wSvxyUUm5cILjDLoX1lOopIqnI7V1Gl5Hhj/pO2v5KYtvhZE05MBob09cZsaiTpA
kfDfL81yjheLGs/kX6VzkdYR5KH+5RdJOZb5l+hA+odlSCk689qJxM0fPL8poXMh
jM97iyiVtFq5OV8bg4MXxe6tlchdrjKcLm8nJ7ntQl3GspS4La/f1SXoy6MkTcA+
+mhiLXqMtdGgB5/fkeZd8TGkenzr3NG9MMN3fn2JzeBLtyrbgQRA9s9qDDqsxy2P
7lSsYdxqTpiCVc7rMVGhOp5Sty1NOHNg9u5WjhYqb4N/+Fhwj6TXvO2X4LhpNfXq
5J6DuA4C6Uov5K3rxVFK6o42WRwmANlm50p1BergMywu4uB49SPm0hM7LpRLZD8E
eI820i3sTmvcUQPdiFcP8iaYvz3jhkxn8WAwS2lo3MQi8Vd5FEBW1oSUqZkz6Z2A
6hwR8XKaSwdf7sBUtdJ41krUomp8GmFTpJKBMlQxcdzkKnE4zbrm/bWl/n33k0OK
DGkMmWbaHWxRp0D37E4v4WVNgzTRaIk//LgJVr5SubHzZeqzYOQLc/j4zdycPEu4
qda9bxnV++XZEyprXmeNcK1+ImtR5TVKqz+DwM/K8mT5i6BjhYLR0ZmHtYcUlBE4
rZfz11o3EfFcn2oy0f1wgVqsM0hrXXq3MP5QBeDrb/Yu0gtSSTrFavqI4uooi7kK
iH6VzgF1LXFUloPXpHO3TAgENyQFPtEdtmpbPhQ+xwF8ZttR4Schssq+S6uA3zNv
PhIto2bf0Xb7yE+VqATwAX32WmaURDb0ruE+xspkhsVAkjAUUaKzIne4msRsmRGz
MhL2PGL50RtoZfUxGkqJSgvgsmEbcd+/k9p5HYA8yBpvCKQyXMSMFwZeTbrasI1l
RsF1l3xErfSESmuYgQwWTVlqW0omOuvNq7bIJVCNXXGr0uIHa9neu2Nmck2oBxCM
N8GqeKkIcyOVpaQFc8dYEoUs/ukYyEEHHWitW1rFsmkXuvh4K7/O7xDyOzGViYPR
VSrI5mCThiA7H/IIHQLAiWTXzqvxSSEJJvcEom0/bCptbNy5Q4/4w3VJ04/y7F9g
i5ZJfTBn2kXYBItEQGAwO96Utb+269IzEm6vrg5cnpeF7CUIDoA1gwYMXDw4CMRe
BcNwOmvuo2xDj6Qyg+a49MT8mAdFBi9Hq2B/iFT6FQ34z/rHr6NRjmyn8+mhDGYo
UAEam3g9SBVazgyR4mJdst0USd9qxJlnK1lp1lfIclFGDnj0NL5mwHRjKCOJcV2S
ZVOUvlVt5Ylm0cyI0r1EMGNy1xmoUbO/nHb53DESK7bjr/yZu47jQJ3O7WGAv0YR
1lxDy9NH9BybIq6WqwqoMTgs7OvJuFLvEguMqQeypTNvy3oogWTkCgDum+WiJe1H
OHYI8ZDgbPTGtmslOU3MomoGNqNAY9b4OVngXydlr23swkdLaFl8uXrPaLFKC16u
E3rXizd4bQhDG/4A9vCMShy7dRzWpGgiEFlBpg3UiyEB8ckvLbankAVewYTAVlxj
+LVduod3ELioH4Y4S2xVZMp/0ypGdKppWcRlEgMUvLeCggdKJxcZV39E883Jfjzx
ttPnvhX8+tDKfhkr6ZSdT6TB23pxy0S5b5wfmw7bojFoJQkatt0KHTdY2kHLt5cf
WoprIsY+o/ibny91NVQ+ed3SgsSrQOnpcRio1312PKkRSoCUZY0DLWDl27hGDm2P
Gwjmu6+UGGUnEJuZVNp3uHwsrJfwfQnO3AB4PIl28Qkxel86JYH/HCOx7SrLAQy8
qM2dhJFX1GJoVcQvrYf1q4qRZgoeQ6ujZhDxGViWbg8IS6XQnzh/vbL6RgOl7u+x
TiXQEHPUPVzVDOjmnxr8pSel+4TGkbHmkIRE/QWDan2ZYMTM1T5EWHPqoXWmdarG
1LLdhqxcIvGLYVEvexzBlkTjrCyYR2beZ4gJygicF0y79fT7rZICvDne6Uo1Mn0Z
tIGNfIuSFesiwABFv8txAlP/czxZx6vN83BqczCykZNefEP0atXFyRgIk51xT9Q2
0HaaBNMCOlVBkzXv250P7yOMFYdPDKSDhtnHAM2QszWEkpAtYeiLjdl0MSkCS+Dy
/Z07mJ+lIivgcoMv++/S9tbLKM4Lc9zLbP1u0DsnskzaEsS5Mrkclq858yEjifpc
X4uBg1nVZTen8ytdjWa9P7zZuu8EM4J6FBiPEGH9s+YMN5PuGhEXHafQ2yXlFPBL
vyOMIWEOLsw7MOmCKu3joPwN3JoQexXNGgUGxrgfTlmoK/HUEMZZ66140HqURwCH
enh9qvhDKScEO1UVW7XMlbXM8GtpXWV4VozTQAXI4xUeVWpoT6r9lGUNVa1OTRot
6n4+jAThQF97i3Kk1JQYt7EvUN7+LWudMiTPepGffAOsLrF0qMBwd0DhcegqgI5C
D9scSGcPIyFSOx5ZNY+xCeJMlDPkJLyZWLJLhHI/SnEIPZgYTNqib7pwQzucuZj7
pqSpe7Fitabd5iI6oyd8CWl+HhmNb1GXYuJUgG47tdo4mhDQbFV/q+bDoNBFQvai
EPSgjfZk9nsBy29GlxYdU6ena8Vl1f+gX4dDOi9FEEzaqqLGuqL438nDvPs5TK3a
Bvpwo0RsW9DT53RtErYZgNo9s4WYYP/c56JTnqlzVZkABXYoh8o5EEQek4WEnrxl
A0IAazDSAEbblpWZ2ioxlWxiXfVhmvr8JmgzXSUeNdCR/bfcArcJbX+wiK0WvFIS
F/hsE8dfUYtbBL0X3J3Bb329jfuWpEMTbd1Q6Ha5PMCVdQBOPPcqhVurYT1otjd1
W2mHdcEPV2Q2qVzhCZ7btrZHNaj/yKJRvOlOqeL8N1+n8OrL5XOmpy592vuKW5kW
WfBH1lQ0TWmDiufVmV+w5YIG/AqAT/kwJCL8YKNpqirUNBZUDVNvs2+2XpDJBggQ
n70Und4NQmdZ8gPeJxPIkBB+8hHd5IDrxxoC1Mv6vogaRMy6YPdMyPRsyow4o8IY
mdBPtC/NoMpcL0hXTTR2PFd+/jmuB8+vbvWgba7ZDixyntmmByKgk/xG2uVeieXn
MbPRp6nGJQmUPziB2dORG8WXzLxeqJN1pOZb6/EtZePoLAZvPZvUcXPahU9UgqBn
4tIQUMf6sji2J9QHjHm0m5yaA+PBZt7z/Qr3GNgGv9BR251LXJO1iuqmySlc/z7G
9Ul/VIALr8OPn7q9w1x3YcreLqcGNfdbWNF6xkWd2QJWPcACSFe/whPqRcfgnkeY
ZW4spKYbn2USz1v1UPqzkM8v3rohMUCmb7hSnajpjtV12s0D6IbUg1CNSAdiCm54
jDNsM/F3xNVS009+Xv4NVLjVUx3frT70wyNF1tEgAub+6ME2AW7gfRXgxBdhDTWn
Kxbje/UcJNHaEf2apUE4rdvG296/Kxr3CtW0tX25nAIFSpS9boC+uKCoGqt7OVVU
CQleCjSI6SxjiNTl0rRA6Rnsse/BMG/q4ad0kROG9QKKTCLtKC7BRF7wfVGM8H+N
G4GM0hXIYdM4plI+L0ppLe3AMTezAas5n5cpXkY53njPhywZXNxt9ug9MCNpOHsL
SdbazSvCfsNM01LtavpSEf/uv83FvbprX374OVtxV42bu5AeMBS1PqtnvbJlwDTI
XYXOZXWi8QqPbKB3hRbGN7QvsgQmSC6Gm8o0TVK9w9kChJ5WeNjcxT4ocaoM8v1S
8pvFGV76M1A+Yk1rP9oBdFCWFcnykHOLjgl2knbhRd5C9ws/hHvHN7IbfqgOh+PB
0IUC14Y2jQOXKit34MT4YU/nC4DnZmJAEEFAdYoIrLQIhulLjuMIBtpClAzAA7Sw
FfdzVmv0E4OlLYeBoCpaOxgtfda5Xhgii0iCnPWzSvz3VVfM0kqTYgM4W5My5fSj
xSj6KhV8MscM+lv1inKuGHsMgmUmMuuzGnYQxcZl+AHAVZjxUA0Y9nb9yxKbpDD4
HzG60vZv+wzxQX9AkRTTv/Cxqb8nniFtTYZPncimG7ZeFcBs8sxKvkTSdW04YqdD
+A44FlWUkbGutkMXncL8WvnJyOD6hM8j3nRpAn/eHRIGIO1ylLhesrqKYobTxiFo
8ne9fc+WmvKSjUFx8m7KwGsVT7jEu74uX+bJqqokaLAqEC9FQVJdK2DWOJXGEy9E
2MDk54KAmZ3izuezfeHCIjtjKYCn88XXxxHu18MK8kEKSTBgNCZ/oMaoUVeuRv1l
kt4wThzulJXu0vbIojozVizDvYC3PImhQU+qQnly7U4szXrqKQVy3LspH88wC1gS
e2THbGFKHyChpTr5i2phMFX84/SWI7Cq/izQioR2q+BdNEL03/0MH5nxFZl9QslQ
hio0PHGR5vBJOdEH3gujts6G5jh5Z8jJWp9rpBkgu5y7O2N5JtMIVNIEv8J0+cH5
Xc0JdHF8IxZHCzYWuDGdo/VjkIYOpO9UhXVsNdakH22wdp9eMCiNP1P2NafwFt5S
uoSSpzFZTLIUIV4E61c7uvGZkentMUGrwWB6gnu3wVeANQ6rxStgAnScJceQhKVh
Juj2dBAiCMRFaTNluW5dySDrTWW1MkY7DGYwaa267SmZkVQuGt6rX5zo6BZ99TDg
bbqKpBEVKN4LUALnFEmjXtL2WyVkgeVABghjxO54yoGOln6/5MIIUJvyn4DNwDO6
MgA9Mf+P5Tp/agTxOq2Ul5IB3lAtXKLnlFHDGk8vFsU6J+70ruEfdhFs59y5faSc
7OmYQBEZ+n3ouX7Mzp0nFurn34YGI6NmaGG6l65HfBrEYujOgXpGTG+sXWJNqZow
Qxfq/K3Q3INSTcN0iE/nduNgCpyEXo6Fe1P01YrNaB7UV9ObutwEhjk3Ed1vOiil
8P3ZUCu1HuN34cFOn1cfGjXcHEl+8ajGvxlaHydynHGugiu00rF6VblmsAsRCm3a
qEv9/Hl9IGFfcsuMpbM1TtcmRBK0gXj/y+ODO+plHMKO+UmDceKS+BG7WihV8ZnT
9h4UrC9x6I0XWNjh7qMaXTbWXPwojBbkzTEfRdq3xT6zr9aC4qlPg8nuzA0SMf2C
IqEYuOjq38I6El4Q9tUsILJrK0Wjbemga5Y/DlRmcnVp7DABrlzs0nlZtvvkliYi
aYKq/wTqwot9iNiyUtDf6GxyT8w0/yOdsqPTryokaA+l+9gpBS7dDlfNHsiRzreh
4yVUrHPM5DxTFXRuBICeNlnMZzl66U/4iu/XejDQ78WPYqWMV3Ra22hYdM3vQwPc
sBYbClgHP+iCco5EDNR3HWfdUBE2x7vSNUkHkrjUh5kUTKKSaCVjEgYJYX0mfPY9
YCRy9/r9RN6s4XmvZMVuDqBtzM6SirRtIWVJ6SLl01stM80REdwuO5MEt6/4BYwZ
BHHUmSChPP9H0hoWMtLniLcP1fWMkYH53W9F9d4vY+uLQmPOg+8CJdVDIhVSmaMK
cnB1d4I5APGXoGEwsaDKvneCmRriJNnYvG0dg6gghHPnLK1LPM0Hid4FBCLB1kTc
2tZWqMKmAOD0AfHxvgijjGSJIxtO4kHsk3iucG1LN5ZBt1KMhmOdyu/HLV1t6Ojk
EPxkdK2GjPgfGqHOkGesVPC2PU95KnX8wR8C1DoJ9usgNQVI5CmVZo+7RuoKn8Ur
rHyXvmnjUJaQiIE+QxPHOdRXJDEuWkF8qOc9d2BmflQQ/iVdIqs5NamsMZ5yEkfO
hfFUxm0HdmmSb84b/oEX9mc4HWLYzju4GwGfvZ+s2/Pq5ft7PhiMFtAO8bW+5BEG
XCuunsGka0ABpu8+WtvstnkbcwBkdM347YNl6N8TgVFmc5R0iMmxymuSickdLXrF
lxu0zzdlwPl4weD1/sXtl4iB7EccJkqlJtnv/lCubMiLVDneJ/9hb0SZZFSu35+H
rc47Fqe1U76aHxhuzDtHa7YBduWmpq2rE3RfCa+WQYc0R4Jrtvtkz30moBm8WUTe
eWQtNFLqiH637wkBV1jb3xQaSgV3GBVUaS8qoBWx5yK7h7fIOzZRT8k6rVzKysaG
0GbF7o9Ap7ubBJtfKivQo4vA7ZipFVW0rfMtzM+kcHILxt5tmFlpM8IKP1SEQZOS
6QcSC1AB2a1adY/v7ZA8QyKyHHLJVifM5oWgAee2oa/jl8bzKBtwpXUAbo7eT9kJ
RYn/jt/p3OjrsXdkqyoe2riZ9XzJT8xE5iLpW3g+4L4qk/gc30ri7bBgtKYqsW5g
ob8EbBaxztUW/UotQGweFijWUGEZ1iDB9J15s0UwIIP5lIcsXwuxS49Rwhzxqhgv
oZn9aQAA3nDw9LnyQv/Vls/wcI9MP2a/UGPYyjU/v04YYprVLVMeTqEMohgcHv/N
9FSQsYBqJJhhGb/kGBT3Mcqqtc7cqUs9UCk/zsFWf0yg/pl9A826I2z71vv0Utd5
+WYV+Mk4TkOpumprVQsj/fA62rIoH3ytPtmWEe5/jLcwgPK0mwjAxhfWEUodnZbw
lDRyNIRiFL4IcX3hFkrgvTsc6+3VoHxexF/Nxn2HY1jS1afZcv/ETrnQKHYMdhYH
9E33rb2h8HYjddT1+2ve6UqaCWi+K59vyneKkC2hkS+g5T/Z3UqaGagxr3hZuWFP
TV0Fk8PxDbUOaoFnAyXFYu3YESEj5/t7pygMdgXIxTbC0Srn3WtAEhZmWJ2GcltB
OVX/MhQmMvfEek2HmpJ7gl1qY4lJGWLVpyFbtBgFUizEPLohH0+bm5NTC3K8VbSk
39+SRsaDGOD8dGovr3C4qKuWABxok6av+uUBkA8ycb+Z3pHHnmFWI3VkG3YfW07x
ayzsHT6iwvOHnIUCxD0uDNSD1PEouCcgGr2vk3nBrvFzcjCOo4ouMKmefefVyiaD
cUoeQR/AMqrSBeToIcodOSXQaJrA8LagnrwYPTFqix7Cj+2nvq0pidIc3cqgjDQc
mj2AdvPh7fKrz602BgUKZaO6sbHRSiD/37h3U1PyQe5anf1HhrjwUcCW9TPKojXs
Pwh7YfUsSNalb8+mohpAllKCpR/BqjpSetftAYCdFraBq6bwRSPuHgtTwXi9J3Zo
ySuv2YaX3gzXb4HefDOJZoqZcPbMmb2r5ALT4tXiseNw2qU6bvlXrhy9kUQnx0X4
zMed0g11pUg5okO9dLKiZGt3jzuCNPWFqk2vHVszBt3iPNVOL0ZWMAkY8NcnSZu8
BtwP/PvwjM2Ooz30JSv1jAOENOsFcMujlCHnEzpCN35BQsPM+N3q/3GZhXtXMvro
5t2Ig6SE2OuqJL/AC5B8TmZGeO0XNvff4AMDJlrSrMyHLhLiVgOrqFok3OsHb2PZ
N2fOHokG6OwhHg1EK13+JmlA7LuJdiJg0lP+0auorKSHXssLyL17c/1n7mfQyAQ3
GMwiW20PyAdBcrb12d5eiaCqZTGjdpkvUHSU8nqH5rMcxNCJronMgFUQJ/pbTML/
m9dQHnOQSWr0MVfTtN8H4H4UO8vGknYnT9LtO++q8OTtKLok6XnZ4waGSWDEh/Ep
YrGBmfT3pNi8PfYTSOCyo7HPST0qm6DOHEICdUAcDkEz4YF1589l0s9w+Noe0WI8
MAtsen5SfYKytQy3yt6FjqU6BG4kufenJ4kMLriYFYUM6VCN6mndKpDLJXGCZ/xH
P4qDoTEsbQrbA/i87uECRhcANWM9S8lNIKPP+qTFqKrje4ttYSF+1vFqQC/WOhLU
6nB9Vq6lPWMH08+icB1n/bgU31AbaCreBV6rF5kUKtmAjzFFAJ8IivhBelE7oR0Q
ODzJyZeSp6HQ8rHW7f/YrQpMIokWcLGSMWyBiYkgeOo8AQxzILLd2lxFv6/Ikhle
n5y6wGNaNFWlwBW1xFtl6+7FfgpUi9QaLZxhwzB3SaSJHNcyt/pZBr3fIaz2vyTf
hE1eCYxQwltywUGh5WU5EKJR6A7kD1BqvEeDtyrSzIOYw25pgr4zZNQHwgGyzLJt
9U/5Xh75IsOnGzbCrw9EoErTflh9w8QY9SidJXIDONwROIqGmHvCiN/4UVfbUBZM
pa+yyom511Pa+o61rkkAQpKp2WwMDajyqo+oCF4iiqiPBIlN/JHh5LJZ9rQNxe+r
YNRnZyFul6D3pz4B2ZIvQpWM8eHmyMcSznUNTZNWW4uNDx1iecuoU7bg0fH+SeHK
ZN52wHhBQ8EYkCW6TQUMcpQz9mWibqf+FK2BSOYu1e1BBCZpwSBkHX+7Vx4UhQw1
w+XJVKT53oNGqIIBo4q/Z/V1UBKfYU6S7stnj92EG7rhic527fjFzI1KHD8HAxgF
6C6e3tS8V32KIx1szs4KvLFQPvQze1ObQqlBDsCULkBtzgfGNNq+TXzqj38wm6Gp
B55Nwe3aLIStyRhXAerCG7w9ZSc+sjYqK8gHnb6d1QtAyaYSYtVaAAzi+22fG8Z8
pg1j8DjXGycnFB6E58XQaNaiPxs2nrEVni/HxStbf5Tc0JL9XdSSo4HV6dLoWjA0
EsdkQXu1PQV446i0HNsCgnJpEm9sbanyQCByX6LCh93OnG1Sga6nOWGRUk+z48iS
x06PQOvBqxu0d9ij7sGlhQr880OR5uY5AFIR5RUjMR//ZyeAM/ohh3XWvIWgvXek
H2tj62rF1kc83+zOSsKbuMi877KCSOP3yUtxF4qgDOMRLdARe9wTVGRSJ3VwPJR7
UX1dFYxSFky8Ib0tN3ry84+iUt4aFlUa3F+vau+gjnCF9OZGVmUTZHT3xJwdE4W9
TaXE7pyH1WJRuF7BpHdi6t1JMBcZxu12Iy8EYIgYLkYZMCySlr/lrgsfKRxgc1/F
4c8M6HsNKqdKwih0jd3JzMn5OjZ6WRdF7tRbQvV6PWlkOR/DtuYuVPcAi3SHp2Ra
8Y3bEHZosPtnzBpV5je6i5d18u5jpcVfgeC4jZl+JgaSpVidbzjYdpI7GXVn6U84
feQpkqT4cp74FVUx0htbFeai8uxjOGXTea+smTnTMwcy3hn0fl3JwbHpTnHbCAf2
8Nc9MCjpDIF1ql768Dp3OFnsvWPYoorGmlDJj/CjJQfX+vxQDSw/BvSwG9LrGbgF
FABjbSOupLVXioLl28vlLDWXn1opvppmkmVtHf/if7qsUhID+4797TdQTm8VWsyj
xhpxPsgZmlok//EIoVMvoBvSABFhozoU6C5MA5bKagMvpjHkFD7IpLlDc0omAy8s
PLJeySugcSoZf1CnWgurYYehFAmDIzco7SgG/8tMevR9/iNznBLFREc1y8cGdaMI
4eLuToTIwO5IbTY183YSsn6oqKoe4L8B1il3mF1OD/EcNzksqy7azfwqP2J9dkKp
s7hHHE83m6w8cF15U08s5Z2fRl9QIRptIiWO+oc6F85YrdjIcQjiv1Yx7tD0FOQE
NGz9HczSMBOFvi+t0RIu5wix8SQ7QJhQacb6MP4UsRPUDh6sQFIJDULD2PizvubD
m5KWH8hthBfCWT/sFMoWE0uwvoFnhP9tZSWgnfFwEl8iz8UEfX4NQFvEHV+kayEB
TwNJ5suDkYSQaA2joOEtpaCYy7iqLnXzykDE4b7VtWLnBHTE/9hAw5W+4qWTv96L
4hHnTQukK3kxg79cHxwcv2+MIFh3kwpANPWXxEL09LPv2DRkojB77JI/j9t5DyFX
Iop973bOpjMCp7wQrQiETJjjlj9Wj3Ah8fbmO7+don7nexrYs1kp5B26GMxRGZZb
mI7DDmPqf/dISS9wSGk0pLyBdSK4I+ptXN3bTZAVr1F52qILEtg3qUld5qi1/moW
o0QPrInXzWQegxNa3DWvm/4+RSpSwiuauSLqkbEc254irwT7a7x3cawXL4XwI0uT
5OGQTN/bwwCRiET6kAD2aix7dBfwyJryadAqa+kpmh9logwdlyz+1k9CLKewUsfn
v382jSz0noUVlM4GTZNkSf+oGUyqW0OWvhy14bso66AuLPsUWHHnE6Lui9Fxo30h
GXSTpMonpv4Xr884TtfK/DsfqcesUrvGOlxZfZXJVl+egAqOnk6QM740223Bjt+z
f/711jMFugYnJEGshx2xFfH8b0VaGXVQP9ntgP+jUa1lMGfyF7GWv60mzc9b54FB
GjhM3Xv3O+GdIJ0iwMAkVD1sgJFNs57nITSqbqIxXN4GrF8VHEsUyLuzHEYIqJzW
aHPTk2nUsIwoZb+Vt3C94RXz480eam9O+xkU4HzX7qNKNijJ7sw2ArjMVV++hyq5
PCBjJxARYyBnU4Gc+eGoPgdf2zd8UTNksWEH3RwyF9yqU8sNuG00nZhRRLWV5PY/
UR6lJ8TNXWaurSqFGy4H3eq6712/T4BQt5QqV8QO5jnNXb5giQ65zeIeFbDuU7dR
YcbCx8AM/45C2qlAyxHOHNAyPtq0CHdh3p4B7QohWaunoZXk/FV1ui6TxIcFLHP+
B+L39kpEnSnfAbax1l1IK/iKHofLJknrktJI0qhA67fs8Z+IIZTzn4QvC4htHCC9
p3rG8PVYSqBrKvyQUuDTVp2865I0X6SHexcs8L9ggRI72HbPyV3RxhNx9b116LaP
ikVGgx+lVoCGlpi4ip2kMUdBm/rL2Bb6o47OeqTGDg5YmqpvjQ5b0WLimCtfdLfx
mo104RQCUp3oGfFntCo+A8xtxZ6pTzqQm7X2nSLoGke30160pz0GRtrCgniEKX66
ElI+W/e8QVBhoAjtsw+PZ78L2TNcrp1QovG1MY1eKkdqay6/vjHQKhpNWFrYN4uY
brMrBbc3fJne2PD2VmYrW8pm5ClsETngbE/MQdHzO+4BA+iJmwKLhq8dqwP+EtVm
zo6rqGjbFHF+BABQCFXH6a05fpL1LWcQUiujJYK+VuwkNswjBi0c9nDoGqyu3tAM
QorKafCaXHeYzCISa8iAlxbT9mwdL3osI7BtPSTsYJf64pddwIiQItB8S79GXjut
7K0826WGjbl11GMvTrn8Xye+6omkr/qP3c6IxGEM3nj88/Usd/Uf1gSsVfH5Abk9
L1zO8/oxi0zEgHY+rvsside4Tm+il5A28gioW4bcecOYm2Rv4dEpeJhy+BZbsjJu
hchsPq4rXkz8jeaHmjgsHjvthyYo0f47v5G/JLX+s7fs72UTgyIGtb63yykiTpq/
plVXJCZGXDOk0Fl5jYlaP5MqdTtr18/AsulYU8N8ohpF9gcvpV2LyHJA7idASbQt
lJf5fbbgp/46r8D6blnY46rG4giOk8hYtLrJL+tp9kSpnt+yhxZWUDvByj7YvKUX
06M0BXn4CwDlIka5ZdeQzCTIq2h3jLaISLXd1voQQYSLXWwGy4K7CQpgkZUZ+B4+
xIZ9ppThQBCkf2qRQ+52EqpRCs+yodh3umpM5baHQxg2ujSEgO/EN0PEQAquBpxv
ZNkISXDmwyE69yQUZCDfGmf30mDNTlTnsAcOOyMCF6FmXKGOlWP7solQQa+zMSJT
kMLEGhquoJm4w1qEzICJLLzouYQrOdq/FtWdYmfrMZsFjjMvxTLGBZFg0OBfyxMA
1mETcDQk4Zg5N9bm7j5eVvlmx2+3x5Y9p00pjUpwMVcNxS4tL04GdJyeBMQY0sp4
/CdCKgbCcShi1kJEcS9XJbDP9JxWG/6+bzrxMSBhofknahmDpgOsgSfeXFhQ+Je7
+rEi6bjsXXwmntJxPtfBN7E/4Uh7sB8EYIK6hv3t/uA+1BtSR5e9/BW9jcAlerhc
yC+9EiHTPHHVoD6mqVwhogl2VaoJmlJPdjjOnUPdM2tIfJ76nZTcHGmpNIIXP3hk
BH0eyw7sslPr89jm/Z2EaNuU32XhGnGrrsq+0bNUPYJNVL7KaRlIzQyp34CI3QvJ
ZMMiyXszrp84JaOWc7IKSnSXmMCN8y2SMWoQTdCNTzJu2ZKYGBkSm+l5NFzEP9S6
eBdNRa9iEZ0Bsxe6YxstGJI7o7SwESA0KWMgoaH7zDFlDPiyCVCvIS6phQZWTP7h
tlOxYPDOABKtvpPRdjS9Vk/HSMfRfgGI7GjU4FRxrBCddeX3Cd39L90qxWUy+fP/
SmwY1mRuYJaBR0BC9u2uxE3wY1jHi0h07Ssv7aHXS1EbmIvNY+3CM2RGkgunKplN
Ux30jsEaPuin4zpCDVrKEKGn1bcqG4P1t9shOC27OhUKP3kNU+o5QpkZ6S0nb4cs
iKNBVh5z7Ti5aj7c6SxCEH4rQRlJL5xfyn6/3hLsA3zQBC5ooaWX8k7dboF4rvYq
6kr0JWi0crQM7odbF+OGX1b38ZC9JJpfN20a2NhzENiEsSxMcG3O/FETYSm0aTXO
vyU3S8THkzaeGpIdvkH5mtN1JLq8LeDQd4inOUn1r1k8b3eWkmt+ROYtEFs0rQAP
OEo3RGP7BiYKj0mmfQIcE9WNlK9vHZ83TBgBwazOrNU+ef/ey28rc+PBf0SyaCQ9
v9htkElXW7gyF9kGCTD6enFnsuNVFSix2FRq1V/7SXXe92e2pGF6/V9Ab9aBdCjk
NRsBh5ttoNp8eO5afR/4DOT2779VNr3jXYc/km20fkrasSDE60/JY3ws1V4j/OcR
2vw4Xg1nUNlDY0yXdtzLDS/AkZtrrGDQefo8D1myNhPVujTu3jcgWzrJZoC6roJA
bSrz7A8xsBnB9GPHpysS7q1c+NB529IyV/TVyjaxOfD2de5VH4GsSm8/aalIiQKW
7XJ8er1SZdEWg3wSHnF5DH3zB2JJBiP2bhreiqC7n/Z+Bs9pagIyw8and4kgqrGp
eCOlV9ZRFHl7abi3miZ/q3aJYFcBv/uWE4Od1Y76aOK9U9ouvo02s1GK+0ugNHKn
yt35gxwTAVO9RCZPDNomluKkR5IkmVgyGCIF+pV5N/+bFKPjbsLyOs43ziUjbHjI
23HjypMFMcHq/tlrNZWn54Rh9z6hFm2qQ9w1wvbWyj4FkR6aUhQQGkhH+Bx4Hmr2
1lM2M1C/Op/K1jlHoOvv7nGMny0Uf5dkshZDZCBKoheuqf4kYGYwaFfomm+QApGI
L6Ns4gfrQUWOg3t4BvsDd4e1aFISiYUEY9Sb1LkZG+qkneMBJvJiHY8LcygPQcrR
5F/pikVWK/w8id44SJcDRHDydwgnAw9LP59NFyAzvYua4zR4NacMtyZlOf3SXm2R
knS2NmOdoKxEGKY/n4DvkmG3giv1JlfYBNuNP7x9/XTIW2XjBZ+lHJE7y3clzCvf
86L3rCoBMr/+8vtTEnnldIepj01LjifoaYLWSi0TjGjT0GlRtvBM8buXGjDoQBsp
SLxBkLQRUF2c8XA44Y99r9uI/XeLHhr5Pau3CRItlhk91tW/ZjwjEjA6ojiCabcb
fFQtSlCZvR0Z1kYsBwrdkeYfZ/xRRTcxJ5mVbAl6fOrjdDXF3zRLUyC93mz5mbuN
kkx9PTeexPyLDAO5XBi1FCtebaUA6VRJpAQgBuvwSkkoFIsizordsaSWIso7tXqK
sL+Y+hKbLiH1wtoKrjUPkRZ3Fx/F1wTSXNnuGpcVh2qefghmhU/Mgula+sFzk8VA
17ttNlGrk8eCQgOkS0hChrIt2eflPwDw+EjALRreypasQrJbD36NUUdqRYfSpPFD
MqBv+uzXFq339eW6Chf0RvXaH5ZfS41JR0yovexegEM0ZtR8ncyH9+pPtPDGxtgi
Wx3XRPbH5ohdVEltA5vxtQGcM2QqcRbkg0ekRNlEt0SkRQoLbFiEvtNUw53IB4VO
2oiqn2OaqhpLVl6lKMpK+LJYPmcA06RkHXWuSbO4xJctGGGoNWKATDwyPG6PqIzD
pIEDdt89FH9NXoPuWf05Y37lL8UoMUdFsvlvbLOG5u1sxxQ+31XESUAEXpiASq7p
/k/bNXtVSZsMIEHrUHEmgzHtu3QEGzbaEG6N+slLZvRdTBHeeQplfrnBQ2oN/EhL
V+ZpqQVnB+KuIlcsTuYyTBHSdkWhgU4AN3Z9iBenHWEoGpN7fWjoQZjIOsLe14CX
uHOH9Jlu7SaK55LkKkEhbmhUvHNHdv9FdtoQ2cTGgDgJ1pGakjryUoHoSD5Jj+/1
JCbE/IThVmJobbJYqbj8Xd/sp7CpZhiDUfCG5Y3stvB8a/CepY6F+oESPZ+/ziGf
7fPYPEcIhZL9ry9QlDaz6L9TxY2EGEkuomQNC0wqymokJ3jNL9AY+ZXbluihyS2E
ErdjjrkGKfF6yFxzzUKVKUdi1sth85vZET9VYxNtBceR8yxiclraP0NxZAPRc2VE
UfB+4NwT/jnGsWgfmC54f9cKyG3WBlDWpN5LXS7QCqRAUVDd2UQmPBGoD+MkwH5P
eHEuAYjvESujSaYhWgXRX586zozURYD0VEv5SilcRR11izPDTQUWzB8HwEpnHq5P
aEq2KlunABWAfmCo2kCrOPd/SoWqjPsS6hJJf27pXKFIQZfWNI9zuPAdZQQaGnC7
s0C3vAmj57DEdhnD3VVxKHWuO9KZX7kkURxq1MO0lPaOYTnrI3r+eLeFbV1gDknz
TAO8FiOv9kYKXhbrtf2DR0OfDiKU+L2Rw2z5k3ldnqNYaOgU0g2ChFVLlZ2zhxSV
MFILwCW/xc6nKjgkYRvQNE84Xkcq6hRT2semRdEwtzsbD16pl81tIKoNPHxkRJrT
ed46kwcOOa9y5rtsos1rbe7Pmd5rdMojET4fS0903gGwYi2IPYt9jXioBiecYeYR
l9XqG1SxpV7NWneO+T43pELppQ4Vq6gJ3dZNmpC9p0kQmv7irJuCAI6YEBIGPy2n
Q4FkNwFCI0g5VETzwWz+rgm8ew6eENcCHaFJQ7i7cck6hykckBZzlmKTLlLZY+Ob
RQ2Adqcm5MO6r/kvEbpfgh79Usj1xLMGfW8/Yo/uRWyZEhz4pqI+xiO+tKxq6stc
lYH/I9h1iEzY1kgM0vP9x2URcmseR1Ye7Z1YxUSZRMPTinLC+jD/N9+LzK7Wh0ZR
K0dU+7W5EpLDmDZ04MrBKTpMBVVj3Ku82zp7ppJO2ZZzXKrp+1kOidTAxm9W0S47
9UiTFnaIwcXoHr3QQyRSmV3jDjHWTzLX1meRQ4+iibs5vQiqsmUvX7pcDGqOE44B
K0Y/06olUT5v1Q0XUIF2t08atYfNQQCGqaRysYmRoUOw2GpCCwGM3bvyr5X86tW3
RwUm1aiYLRfziT+5b7d3B2f6T25cIj9GGyxB/wX3ByStj1arunZoI9X4tDZsVKBF
t2d1txe971bWsVFZMgXR538sTWzR191LzGsD0I7Ref3U0HLAzBAHqzPzO9NOmgaw
VrjYvQWH/ufR/FKux7X6Rxd8n2BmKHlmgNbLRzuBTcgmcdRKRn9AGJBLgvPNHM8d
qUUaGBTAcLD3wok8GZTGX8p0ca+k/KlPFkTCzKtk2SkBYlh2zLguc4Iz3HCrrY/1
bObFnFFXAFnwNEazEw7wvTWMumsaYEftXP84IHtgku14xjQbLYqPaVnx+FIS33At
M6nHVgAXYuOPFpzSi1nKfphKEe6fPm4bns168YXAyVcoQ57kqexA+bWXMLpNbelf
DxJmrpc9cT+zoOXWroLXMWA2tzN83UsE6e0MmBIq75AcNdAUSNVnWzI+/bb8Wx5H
JUy09zBIZw1rQw3uGVxLuiPFLyC4dOje7wYIK6W/Uz8iNl0zo46FHlVl+N3fScxV
uOJub8wwXjii9DCgv9lwUGx17YPyBO8dlz1jRLkzHyDLMfn+NkBLygoJdEbSTSDT
R1vojrLb7oRvgAJC68XFId9n6E4Torfc8fL+MGzRt1hGc3lOyVKge6FGHss5pul3
mK3NLGAwsU08jXyajfm3BRO0OGa8W2ifCnOoqh9X0v5PoB9+5Yyu0VfrNtzf/yl5
zFaNtGUAzhj0vuLt3T5eWVi2aN8FAaSioyXLD2EAX3dHDgv5ASRl15nql8h+7QBS
UJQHCg1J+/MxAveNmShrPTpq1B2nKov2hZjBXVwfEaJNSNXCSKPWdRECjZAaKY9c
0Ut+Wo5yx/sCfqLsX6/R/nSls7Y0i3vokBYGWcLhjp4c118gl9WsNYtZhajSEI35
GlgQBhCLQe8brKpo42P1B0i7yE2wUh6/Jp+wKbC3RLTZlfW/aneoC4v7uBbeN01o
BJoxfloCYVvyRENmfrPhdKCJpio90q61FB6sEZzwTZdAivfWeTeQoKTP1RyCPF5E
yE4t/ZIHKLG0y9S3HIdNhKmoTFGKgbcxC8Amh7ZJnd6CuaoQRItlgmmdZHHR5/QL
l48r1TvOWBqk7nWYpw+SrEs9awwrpxshOXUWWbsktSskzr9k0fbrYGwSfM2loKkK
LAvqNi87iqb8xvG295Cf10xzxEAaBNrOkpvfZPFpYwb8lEpVeIkigZvJ/smYKO//
KjNRw85e6un1e2wV3Jbzq6P5PYa0AM8I0fAviPUmrptUCzlI7TsK/FiW/R2EabqI
eB+9XHyzDX8tk/NJwttHN2cyPNvgl9HEzvdy5SeKnXylXtEwGPyMsSQWNkB6wByC
HQtLKMuT7wQAv5PUE4rWWQbKxLYMJZHOs6yYxTG8QI+ehOXEr5/p+5wmNnjiICk0
P2uc/tlHS9M+rkdAYIie7ioH6WDyUbAeh8z2WqE8+GQGBYDc/a+NrgenRDSzPmOV
vwi84dvmqlS/bB989DiGOcyJfzKEfKOCQjTaBXe8l8UGlMDNzbPHllJbzUWHChF3
WAQ2C08JqL/4Kz7E7euO+MC6F/eKyg4wCDb1R9I1EP+ubOPCJsqp4/sENf41UPiz
dn0azJM8H5nUS6u7nS1P2EDIPNRlPlj4nhR02fJ+n3g21tCxmtPypEcFrVxJfxc7
2mOu3JjKi8azmp+4yL900tcqWJWd2nAxIoS6V/W0KBKFXrr3PLWEIlTlLkbUTNdS
ItI32Hs7yO/ZJ5jpNx6g2BGd6AQSjM0ANTB7sA5nJbmSfoqZb+ZQdjApP53aVD7k
ImjyoPMM0kD9tFRW/10PaYx91z0xt4Sq012hc+TRjU8nDC8vceY94nuHzpmovc9N
hIiX0+XuqFsu7I+ieDrLH3XX/61Vf/cGXS2oruaCOOcu7DWUDLb4Rhmro9WXOrfB
D3IHYka5r5PtMKp2aGl1FrITcFzaYq+yORvOHB3WijhSpuU3kE2DoxH8nmjvnWtW
anO4QkuZkiUeDoviXGvXoXAH9FhEfW7lLJCsPTbUBQaWsQYQrQS9vHCTcJ80ynuJ
mxy736a3ACHP4sqYcwnmJ+R2OsC9ykMfS68MOUCKm9TWYAEb9ZYnfwfEohdYClS4
sYovicSVtjYydP9jJa/+nJp75MiGw8Bn+j6xqw2V+Z7yiC0q7H193wfb+jQDHnua
791hm5nNInsAxmJ9VBXebFUaxkdOHkGwfO9BKl/SRGUWhAtLnd/M8RBUI8aQAaJ+
rwxA0SYeASR/Rui3dYFIUkBLsb8dd67/tUeCEQ9Cjw1xXLxDeQJpsiFm230tC3Nm
6lmbefC1W0HbNQZuwCAWshEiiirmW/UE/ELuKg/gbIL0P+P+Q5TqAYQx+Eg+ZNd/
xdsheJqSYYpKBZgIfemUTBrFgDwIKquVAjMzafk2Ffndp8ruBBaWiuQN11AByweX
7u1SzHeHypqrcYLOVFT0MR/wLT7Eg5kvu0BxvUp4dFKJSgHM0yPTfjWjYJ4DYMOP
zH6daUMsyniIzbnRhNzqrsxYjczvZpPGWglQQ8e3GGOVg3NKw6vhts3BFwMo8Ia/
N8Y8eILATVKNcDtjkJS+fxmYmexPRjFPQzHCHuq0j7cluF+0Aqz+P/5LPGHpOp18
F9DnIW3B4wsOixX5tN8QbT6rzOf7+96Q2zefxvUw4OMf0kD+yCsO7zXa3tV9uv8l
JJOMOETOLnrSOIp/yjkB5kCM3EtgWIMpx6dGuk1disuuV+EJyKgX/R9EF2IYFFpR
0JGMaFyi4ynkHmXt90EpWMB0QxAz+GlNcWEMIl/moxXAdkIkZE2izzfdERIsZ/xR
hok+RZyZvaT99gaaVCo9ZucvvMpt+OeTl5n/V7BEqxn8xwmXbrILW3+O8RltEp1r
0FIqT8dcEt+sNWR1xC4Oic3Ts8eIiZBtd0dd798sOsy3VWvZX+fNs2RFy0bC06ZH
SuvWLd4WRIarVfZvHft5OBcdKs1l6/UXdNjy7L1Z5xcz8j6RPC4uAVCromBIDJ5q
gbZPaVursX2lnqSA3guci2K5XNZ9jTk8ZSXRg0WNmsyr9WwWCT5zaO3JUoKcAZmz
tgyv/mSTgUuXJbccNU6dR8a8Jt2pmvqszt32HiTVlXAVfJQFUzGspfz8KPruDKQO
sEJI7uGs4/GsiSBX705ML7l94j9hXrjySzniWHHmMaNSUymKYaDvFA7M8ubzM8CB
Uh5pNhzYIVbOSOiueo9OAhk30HyeGY2fFhXXFINVdS34XxyzWwNnoq1+7oDullEi
4FnEOvOFaBISF71NxcYyCSREDG9AR/pb1Ufti44YTPE/j1fiqDcHkCcgTTm+zAsQ
lVrcCq2c4b3nZ/tTDiG8QA6eZUhJoyBWzlzvBdySRA70MYqgJpBSlhy31Q7I9DC6
OLOH2eKjYwKrBsqIC54Gk7Br+GHjyZGDITdDHOgjM36eEo4vlej9YT0B1M5Ajsrs
1o/2nr4FT5rHMx3QIu2901bwhB3nHWzUeLCCt5QwH2ME/EkrwVCDM3LpHrINnlhx
3nRS/84JX+mb7EsrZCOsPcAZQt/bsIKfGgknajUYXDhjfd/OubVbsauFeBCskGq+
pEMMiA9bniy9rq5QnG69RKGNeVRquX1CFvFD79hLirCiLBw+7rF9gpYCG0JNTNWQ
MA+K15pJ7KsC5yOLBUJqyW9WwQGnoUm/wyNEyqOnEMR73FMH7byXNkzL3OIHbE9u
WLQQ8fZGjDid5gMZNpnJLfE0Pw/it2t4WY+mPJGq/+pLC8zua7WKsgmnoMWRF5YL
6bb5JZSsTmJBTrqV7LlhXES0lTPa+7wjfnBwn0A1Cm8ykFOR7JjIpsL7F/GPim4g
HGWB0Zl2hogN4I/FTV7IW55o7SGY09m4RHrcZQVrA2g9DcB9qVr4RwnRujt9+sPs
Tcb/q/nxQrYbq6mMZcYGdwU/aMCbwnBRWYuRfQdSTwQVmiV6r8Qe8MPyFLvib5Nh
kQYHDeDCU9037MXKL6WLGpocjidpF9dH9gKRCZBYmEi6zkJjTUqyY4JGRTkyTtRT
5uNgpsn/l74Q5GfaEvP+h0eW+NJ9GRu0cI3CuhVeQRednhvlmAyZsrnenlR/WwqL
RleVu8jem49eoTBFOSLSFSOwhQA/cdJAuZfLdZRFOWjji65e5JYhEmQz4sCjLwhz
Jz83hsa4M6JlkGIB38NqH7xw4yFMNo6kAAi/jaKwawHG77TKRCFkQLYWWSwTuL5R
lAAn/dgQr+4wATw7/BqZdPDVHOq7c2Iemx2G0Bh/c98NH4EzwNYZaYfjN61lBDAv
XDQoxF2nyVzkZEr1czS6JPGOLCJpq/bEmedFw+4YpO/8s3xw41CbyP+8SjdNX6Lz
6UyPqagkCMjqqTwYp/JP2MioL7i5G30TMqLkc8HHKTa0O/oHd1/nvqiHlTrrrOyv
aIGkafopebPZGd6KdMpaaona8+GDeZtVr5TUmsf9u9VWjT4Ah4XoWjnf2cBeaadY
guDANDhPTIxPCfLWRM95nB4gtZ1DER6oQ+1QVCK/7ARpBF8uRw+Z43U3veTp1em+
FT6mAsbVuPFVlUVeHgvnT7tD8g8FEMz8DmMH0S9SwngvqYWGEQPCilpUUcjnT6g/
qth/fKXRN/1HDEMFPC/HlUy3Ik5VUcDvakZEKYIZ7yuykMX98mBz4YaZ6yk1h0WI
ndnqfLbuI8CrDOpcmwjI0wN1zdFsGg3IBVcdOEwcK6gr/BXjWoJpO9/isGxmG/iC
508ySmU6+YrfqV11M89nTCKFJ0aXQ0F4S5xUHCqSXXnGZP+Vh07rAw8LJR0yb3BQ
jztThqBvCemIuvQg4fdKKtMb/wkKbNnZKtHM/3rkHYiANiOdJPsppJ8/CUmOHHwO
G+N40SFtSa7bq8fse7pyERejgKxsv4fYkihWnMxFMZA+SgysUXT9Ki+EG+tca5Nj
utMrZYu0fDFykOSbKnI1qFFDboJ1FwEVfYcjIOR45OUrQSngk31JmJ40nX5Rub0i
Pl0jidXHcdEK7beuFriuuJI+izm0XFx2AVt/+Wwy46/ogcujhzqAM0mr7IrKRoLS
4RoM7585WVrXiEf838MyWG+tvYx9r4bZE2Y0lMnTkeD5iwAQV2EW25qu7+a3R1Oo
l18357gTR9iczCRqzxSNKAjwyCOZQYTtP78HMdFHtXLKzdNWE66j1xd0zIV4DbPX
QKYIzXvtt/ISWy12Qx8henhtd94cEXBAIFmXmo4pMngst350p6et2MGAF1bFcgfd
a1fieEDx75Odnkk4wLbe8lsHGVr/pbpxavf8RbiK/+Wyrz6bhnCVyMwUwktpwQvC
Tkh19QP1IPIea+D9K2iefQ9pPxYUpNGF0acXyb+QS1ypGFoEGDactsgGDmmqIvpT
7fwNNzAtx38PbRkOkXr9PzIzLJkAcnhCSCqYZl9mD3TXuJvOtKumfNmeZjBWEbSf
9Cph4dPK7P4ODbD0NjAitwohOrp0G8PJiLR3WWgToyF858vfJ65QV2f25vP8ccWR
sZQnohksqWGtggAvG38mqc2+A8BNo7bkzJCGkvelxqG7UGYl+zODwe+UFEFCpgFG
T48Sas6DmCrZ9UTh0n77wfjj3LnXMyX3qkMIIFjUuDl7t7lLGNPxE05E43d4rgVy
Sequl9fkZG7H+GKv1j3sWRCHExYByQwDSH0BwrTMpQPmnTREqlBriy3rAmSQ2uIP
tuNzZY52oC91oWsKHpAN0ufn1N9hfH7hC3m4oji5zJuIbCFbIwCffbkKLHZ5QPJc
Zt9XvEXQSrt++wTtv94LXlsLcCrP8tWsb9B/Zs2qJOensDUkd9hyZQqm3EX3stRQ
EcpPmNYOpeBkTlDh3XAyfNmTD8CA8C57PeyZyrKv2zP1+2Tu4U7PKPbugk8RS9NA
F9xTYP8o+C1Iv7ba7+KI+9IW+MZwd9yS7h2GHUIrDCtBMKcJJacZCtP3g3oVTw00
S27qavEFFgIyEkFG6VMTqD4FrLtkVoA/gs/fD8NlkOh+AmdNPHomIQB96CTkQC60
xDHJPgiPbO3CBwKBb9Gs0qDUTh32hqDrAUw8RS5Qm961HLaa4yvyiOz+C6GdRFkY
y9HUvtNFPnNCo6PkdefezO0cn0Q07Jdl8vwhplx+RpzKNkmWk7eT4rpLJTDV4UNK
kwJ5apLTpjmrdcNpjQDr1FDoPkhkSzzssEihBtMHyWcejMzKe+6XY/9zjccIZvFl
GPZuMtVtHfAfomEH2esfrxIixrhyQhxncMp5YzsE0gKzAtZe6p5Tcda9Sq5eprrH
V3j1RVJ8amyi0aKYpYu9zPmAFNlOEP/0Prx+/rC76+lg63HguvO3raF84RABILXO
olNo10k4wWjrpBQ0DYsoQ2xNwChCxRL9pA4ISiBvyJ+idUif4570N+jz7gl+71L3
GlX4Om81WtybdpgJYi7ui1dtuQUIeJaaItktGTzx2Svt5DtQr43h6FjY/9BD9szS
5b+v24GT6pDwHbLNQQyoRk6k49+xm2e7V9Yjc9d3o/djcZ47mzEhQSpzu62wNe/9
Nd5//R2oEMu02IolwE+vMv4euvzO5mOe3eLQkTEEIzOxZjZqpIKgN/1o/cWavaHK
3R63M4I2tYBmFmLv84CJ2YJJPfFeodW5WcMwGq/AiSGfxrWIKwpEQNlmH6V7e5/c
bIdgKVGB+TP7+G7qA9I0yQ5PpF8JFfiQgx+CEl5iNozV0yM6XaOWZJNSyjbhlUX4
XqA/EyAQbA4nHUqZjm4rw3o2teoLqInj88cMJtQrFf56wdhCFTBtQDy+zP72NUof
xsW1IoJWwJreLdDWy5dHff5d5meDHGMxtzQnzE/YmqkzjI/ONMni4bEdU9ATn40d
aOsay5xj/OOs5tlOqFj2olT0zu6P42Ujby2MMaA6ssRjHDoC4PlbHdMnbGhLu71W
5RW8TQoRNFrF8ZWZQbr4iIJykI1cEgbIi5HOzQAx5oztWbARzEdAw5+ZXS0HQAos
9pig/ixv5MysmK3lO9e2neYT8zKpz2NcIQjXJLPY0qWpwznkEgM91wClZqVmbpu+
HA1KRd8czSg5DlvhJ3P/JOlPeaJ33aivTw5qJZmpznXaNgk1KnRuSLK+twKXXxiQ
eWJ/lNmdeq5AxH/AXgH5sfdTWNZTtWLaaAcAnbAm7DadGVEoDfKQWui3Ve/AtSJe
8fIQWhI9X9cBGYBJJJ0qRJuadhLLIcKOP6wHPWJnWufmGvIkBHGy3C1IxGrJpXMi
4cpnPnoul+Q14otUnlTHEPrCBRYWaMPhVM8j++Bfw6kBL3VISI2MH+h3QK5EhBrs
Wm/tNgUeJ1jaQUCJEuG5RHkAlkqZPwRXoIsXjdXfAd5BDHsUfmx5du32iJCmK6wG
habwNUppNHeXJWJrq1q+nOeLwwjgApeYQggnScrWjRqj2esGH8WTGxdde/L0OUqk
X4gyAAbq/6/RN/YtpxKTUoZzB2Jm1KnePTd0VgwXMwxAfOwkYQf0t1B8Vak81Utr
G0nm6oku1ZsG80LcF66DmvOI5qpi9j0DewAm3n5PLzOi0ev4HxKxfKFaU8mjOcK+
9pJ/dn+o7wU7Dzi6QmnG13z94aJHTPCbhsjDr9t7m1zdk5h+7qNGNQBhETWQCcNo
WjBsT82O/WcjZ90ic5wSNFoPflG60/kQZdxaDNzollngqj1FBB+6e1iS2x2OQ6XN
SqODbWUmEp9ryHQBZc0dvjbwMBuHYsImyp2Wqci9F2OZkcQjtD8PCEqWApIi6MxQ
WQ+LW9nWVt/2NRx+4C/wi5RBpMTdvdLkCRhN1PRIKQl9nx0kJCQqUkFIPqLPm4tJ
hOWsIjFRlJ7VkoYus4bz3qloyZa3fAzlt/2DnBvVuRXP/46wdLiHNsDC3FivKG6O
ayiG/idF3l7lodu5E6xJN6pyhzO2y67Lkv6UxkJH1F3MgItkGuLdU4dImFNMkTpS
kp30vhTs2FGJhU90KdhSno/RAd+4JGMwMo0jnzf6XZsdZKAUzBSnCvtkRkGVqwqj
XA+XxpDWgGyRTKkF9sWG1dkDF3WcOmMxSuhRp+TPFjktqQQDOqBfeGDbS1cUMBEz
JqYXmgYgIWopc1Kqcu67453jQDZ3XBCU/ArJwI6ykQCbfpRtKN/UT8i3CSb+9U4l
XHjPsg7oMASFQ4XMfksb0Xw9U+BIYJFaLoScKKE19QKpop+/kb0pdMi81syxPWZd
VD6kJbSKrCCgxUTds11zQL7N+5bVo7YDYwjZf+qEe2m07N6ilzT+5Y2fnRTPFqjJ
ze4UHWCsnUFRgbRLd41yTW+zdIZNPfCXGCSE3ck5RKCYMWHyovh/bvKCBhxyYBLS
Gf3pqpO7aJndZn8K2a5b2h7nslexTZwTPvCJQbP2+1DXVrjUik4hoeCTKcHjs8EO
AergPNuHaqn230kisrvViTmI3jqSM4GIDRyxaQ4REytDKBTBrtSQtp8KaB4EbV17
+wEN5W3rodD2CittkSUPxQIY6/eDGWs5q4hTVjNQgNxYodUGOFdSoglnxM2tY104
flIXd7TgHk+jpooCMDJW8OnuE1pbzZm64Ryt7c+yi1MgfEVfkuI+IC520WuFK4dn
5i3SsxBtTRtLPNLp6xZJ3b9Vx1SzSdOSQpOIz4RPzNHBgFUHmd3kSYeeQ+Omsmq8
NdURivPNGDNz4bA8um54t0upGwlZKytv2S6yllJwukZS8yQFIPQlQ+q5lPpa7NXX
5PokUj3RjgBqKL6GaUpNQKdt9GS/CHWRadRhu12a7SbjJuw0oE+Etfp81sGghP+f
X8PnNi9QTnrJaKsCPyNjy6QxhYgarbWBMvYqKu0tVvdpPFJZIeXc1ayZVvRQvzGD
YZhPnDk39GjyFto+J8RW8w==
`pragma protect end_protected
