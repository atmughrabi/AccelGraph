// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rk6Ywm3zB6VtI/itL24u2RY68crlH4WFTKIwQQD8TLNBbtQiYPaBF7PcS5q13RQQ
vQQE0JdCLFSrPuuMrqbD3rEgjhoNfVSAIIf/vDx4HtGKbjPbUKfrxyS4BLmm/b06
K97X6xf6tOMfuM5B9m90DKEvj9jwphRXvQqmPZfRX0M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11056)
1os4nO5efab/FT/BnYKHNCwdRHqWkSiAetZCmyDWKLptdSbDFOwNdFjtFMtos7c1
ViwlAHnomd3TXqXofM57D+MXkAH9HJbyF2RVi1Mz/D/QDMfCp3xHAARmA0PuKU+A
wwPwqFP8YhtPYoNLoXPjX67dUURAWf1ifi/AnbwMGjx6MpUag6WwOG07e3Z6rfBh
gAZba6gu2dCJYHhWYDcpmxqOnIEMlEAM7TW5IGeLkWPvg0chOpdQh7CalxaNY6SR
VCzG7QWoGhIA43bU1L9GO5f/e+UFwGEAyCVQzKsdgJ8sIVSyNg8BSNhfoggLxr3N
2FYDV9nReqz/R5yxZzoMEsCc0V7W7//NTCAzq2B1V6MidoqxRmgP6kGTHtoAi4ev
ysiNETRUoKmIoYtl2+bUlDS2GVZOWWwazeUCsy6iSVIJ6zXYts7DMPaUwsNSKi1g
GLeSvWW2ji5a6nqLbFSR0ZZRlNtvWl3uPUA9tZfbWM27n/JtTYb9/LyWH5PtqE8W
pJyzUBiF0rHqY9N+6HYErlQ+XDrtV/eYKbjRVanlyiux9h0luksrs2GX+hRPSH4l
gJsCWNu7WPFeWUD0gfa/8c24DidO7hIm89cJrEMX/SXtwav7GCsYQDKW/TuArB/x
t0ps1ZynbGQ1OHDdu1rQrzO8FrY+Vesq22UKk/cPO1JGqJiAR39GsI5xBn6BEHw2
TosOv6juMvRnFeaBIGwWgfaC0iaNzLGOH8DbE4MMfA7Rv4zxVpqxvL4igJTMyzhw
f3KrvLAK1zv2pbYWbD+/29c7nLMZueVXg/MVL8KqU0Yd3VVkyUDI5RdA8d5TvGCw
XEgv0rx7XKSTaqqa8Nm7yrlnARhtenwWG2SfSODxLUaRTPyDTKEUylZcxpkq6ovA
UtxkvU1KeYtbLkvBZkxL7pULe+VCiY/p/LlHdzlhBqWnxBU9MJJJOqLGj4OtR3Ed
WZ4waOg/asYWWwT2AbcEXgNHqV43bS9e7w3EKtUwnOzmwWq79I+lSi/fbl+NtnHA
1mBpQKHgu2ssqxacq6e3/isqa68ULKxCC16iHqKz2tKwVKZBSfdwkLOXB2cy2TdD
xwd3cShV205yZ/t09cTjD4ybPy5FfKW9KaD5MtzFH+Rhjilu/NNbLNsQy7yI93A8
Cxwf9X5aRpfwK0Mgnh3ObKKVW2QNK33x76tJaBhjz2KTv9OYdO7V5qxubQjLtkI3
bdnNJ97guB253MJu2PSUrdrnkF42o1q9SRt3kiUk9aQnf5ALrrkXDen0nBbUMpR8
5doNLkauyqy40+gD63um7qX4MAgZtf0rJBx7hyddER5T7UlutgY8kj5kGUE7YFL5
slixtSpPF0ZjI2SdHKflOv6UkvzEQZ/7ut1QXM9vdy5BKY7wld7OL28scBo0yL+L
KiJHmkEur9Lmg3HJtzlFLN5qch6Td9A7O9tI6JLcJqB29Dn6JwjJX35tPGxfX+2g
ZJCGnc3U68nlMF8YcZNbHKH3NcfOWu6BBUfO2VLBgwC7IU55mQxhR5TUbOuClooj
q5AdInkv+BWiQXhFRL8wDF/zf9jFQSs37ySYg+BSW4NYgLb+m344+d2HyibW1pWj
dfvTIW821ExliDZVktfTHCGLyKmIfHxKqDztHXWS2JWdGEymg57wu1XD2vXu89vy
CAWEsL03pFAIRMhPuk/H86obAE17xGBdIt2Pr9WBdkgimtHzoyqVmkj84sTEqgyE
89UW4xp7KFdYI169/i/LtRVX+txufZopuXzNQXSmsBBJ/73E3Eggrcp1ynOjyYXH
bxCGxTog8PxKurKkPM6HJ25DJPFd1jDemdDig1Ai3Nfey6ZT6iOx/g7ikIPxMGum
jI+LbVHpJULP93SU/D6ChxQzLsQNU/gQxd1dLy3J8sq4ADNfUPGgUnbzsUBN/wX9
cJ4JUOoSunxWrEHeLQFT5NhArzN898y6nWFcJDGjdfsZys/4oxjkPMkrw+uCKyDm
oXi5YiPIzmypFaBZZHPnvzaKbAIrq24T0vmSPVXAQQNxUlVwSA/lEXyEzQoSx1Jb
KTkIVudyCwdU0xxmKSiKJqyFoIax9Kamnh+ZHHvSdiZJNNe8d7cWBZh5oyzMnEjU
zx2TrDLdcP2uqU20DDVCTBOQic6wTZ4E4nr35G2kaLkZ+12vVraxhhwPy4NifF8z
5Y0hii50cV1Fak2rKx8+FGg0rwB4YhYh21LETkfvFNpEHeHIsiN3JHjc/Z8fNyDH
4AXMqZWDDktFhF2hU2tBfKNLEAIBqk8+T9arsvI/ucrDNuhMY129HgMuCL1YbK3z
K9+bSbCG961I8pnhT9SSTs3Jf+KCTgOSnLOS0aToEnT8X6px1xlfrRlQY2TFOHDD
LDcsOn+rySnsTZ1gsgdXGPaiKFKwEfKdlZj28e56nUKi83+6ujghMXwqA6wEIrLs
lZOYFV1ckqIPTxCoLaMPe6dRh1COS1/WcI4pXD0gARbYkU7Ev6r/FVssoSBU6UK7
na0B4MDqpCRFFKIm/5fBcp6+UWLd9dq6jWnphLmdwxC6GOJP8n9cY95kKDqI3L8S
ZsOh3qrtehsI1TiP57bp8GhLi31DhySdpXWokxLbmp6dEq7hiwvB2n/3yNqDy6/Q
vUHvHHRCg1LnaretHlbNhSIVq3bM4Q8xOQgWSP/dilV+ZvFbEHPu/5ASuEEkKPmF
uZsK4YuTOJe2ztIES8jw/1tkWUXI5oW2qgEaiCU6Nh2pyM8W+lyqj/UJ/sgiEqne
jYtlafShfpYjwxOJnhLW+omWCRwibMQbf6O5xCYyePUghG+4Yhotg7gJgnEZi8yp
B9mk4VuV+1FlsSopUQ6NtsJB16HRqK1dm6Ucl0+jU90s96uW+8vkGwuVJ8dJUCn3
XQkSIZ3vjZSwCmfGDh328pXsw5cU6qf70SUXNCkiMaXfPgDqlKo0m0ARa76WJbL+
KjTQrEpw1lbd8UeWUwBll8GE97UAgx+SDRExSsVC+SvO39FfsFXVjvQC3j3Rlp43
hHeYW0pGHoDxHKZ58RzPlVYy/x+x+VHInJc9sH/1qc53kmTFH5URifC3B6ooH2e7
T+OsE0sLxs0P090h+VSYUVzg1kltehVW+6eM6qJVuovQhPd26SCZ8tfX6miABztM
k5lB4Kt1UsTtdlY02HvkX/s8/0GMrBQ/j1s8PoyOjH7DkIpvatl2RJCVXBItWUkU
xJaUDwfpmQwtn4BkblCLK3NFfQCugtLx3mBJ/s6j84cyZKotNZpQTehh/OiaJOjy
7jolDQCZ6LTR1n0wp3UPaIt72gOmt6gBYbNF+0/JscbSCujyNGOi9CWtOseXZaOu
YgMB7yzPh56c0MqfMrs/qNX/PGW88zwwic/2jzi/q3kc24nU6eCWuPon6hIqgm0y
fTefoFvSvccvH/MbYResib9DpoQ+9ZR2acpcV18NfOZLHdoMNe7064YnjAUC0VMx
bHZNR7SBDeCAc1Rw3c6i1mAYtqKftdkyTVs+WWsXr3vgM8YpBDqY1010j+QEhSCS
SCP1mhkzbE2172mRdhnJVGGnj09YCnro/ALVlhXDiR4TT3ScIa2XigKTHN/kUSaZ
o1sIREN7ZDZjWV1qpaWImmZQcgKIrb+KkvZ7ENhjhCyyDqb9qOW5fxMa4/sYM6Fm
U3nr2+pqJVEHp4N0GWBUbWkPG6esTFQtzbz2u5EjkMLLI/a6g6kXPHKp4Hy0ahnt
HAg7gDRXbMqXMF+7f7dTJ0ZsBy1yIb/uSqXP3M5Rp7n9dEIRd2Km/Z2twGBvPfOu
ckpCG6kFVlpx5q8CMbqncGQor2YrP+Zwbx+sQVlyKaI9NaAJ7mqOzz3eaAwSMwXY
YwgIzmxtsmWrQNgA3n0R4GvDdriOvUppVUWe0S1n8GtAhKLKlYixFY6o6d5kR3TB
UcwCeZXS3UCNVRJXwihYKOvBYFoOGwqXeSAexksuFpKJ6YGuKgWbg+/rFbnXVgtk
M7v8vy29s7lBh8TCjtzYLr/VTVPcKMW5Ba/OoWCD9DavHQWLQVjeQduq+6FXIfCO
41Fl1hduuH+/pdZFNLITKLXsNPTdANxvF3VIdI+KhZwghbUIBjw5+tnhXkK1gGrO
J1bG8q41e0OMCXGKxaK5uJ2+sV+QusvNXeTIGKQdllOUQHNIbkaguUaryNStlAah
YGr770YK5ivavOJLvH/JwkM2ypLrraQyCLubOGvb9PvGWkhWJWK10oxEqgKuTeyk
I9LVs/d8l0zrSrQ4EHU/G6NS6WXK7qBBMoTGeIhslE1WxQRW7dAF6wnIZVwoCHwI
JvRA2imEIVcM6kqihll5+9VE6iOjgzS+h8G2x7Fidbrst/9r2tCvVaZ0ydUAUklj
I8fNft2U2a6icDEUFtN5h5V4uRDCJEz3BWYmamsrjp2IHbnUU/eIq8kesmwJO3eV
0uIvEGDnixfBajmxn/vfOIB8+XihbBw3/jtbmayyhWhoBnZ3rKC/Q7AlHlkSsjMA
OsPBc5c7joWu5jzSMoPb8oeoWMgD6AHL70kfphIml79MUYOj82/hveBdOIotcgPB
96rtEdnCc2MxSJkqcyBI8/yg1cmj4H+9Z1B+F1enm15k6j6b7iN6tb2B9bWgp8vr
q0fVDT0JvWkymLOVstemDDdHP5Hjxm+pwyGG44pfxuquPX7WvEt0GgP27RffhGp7
mNz70ZkfXCjQ96ShTSFmNtrYdeeMtz2v1/j3H5rfTu9pYoRUvYZ3AdKDm0/JzsB1
kgIvg5Kd45CiQoSMFekE/4t+mGeax/DEFs5IXYUOTXf5UADaj0/IV9T6ejXgRWEJ
l9cRjkYsJ7IIH488ADv/J1uoe/cYcYs3Mqn1x7+8XZBcM2fQ6/Gwngj+VNdFvXfl
LPydL0QAP9zSZe9SmuZtC5I29dGadVBagjQroXyBdmJid9Jfou7IUNNZPsLD+piy
4BdWZZNSu1V22KOK7+xu3ASJc/6QQu1hIhBAcwmw/F4qB35o4r5TjEqlguuYb09Z
3ubGB4NHS42pahJYQwGV4SaEieGYchdnKcNDq9p/WMVpe11oQ/JW+yWKluiCvwqS
f153KDT2e4YEAf+C2Fv1sI5pCfpaJhbhAvtW8kgEGoZHwi2M6gajGxpu9ta9Idzr
55GY+jaKGZSRFYnUt3JHCpqpKGk6o3LQd8+NkWXt6pUR7qb7PzqAFazVLa0auTkw
xUrpisgQjO/yW+wOWoU0gRjYnhrqExexUfltyYuA5+TzSeuEddAGg6h/YRdCOUGv
hgHYoEJWRGKjGWXv3QmTBd0/J8ZWQ9GGBqK8IL4A2UVmteOv0/nZnF1Ox8AQlyrr
cr5U12lCVQ1FuUsfGclIbHqsQP//k5rE8I4ZCeyKUNE9meKKd2F3sc5v02Gtko/S
fTHhvI5ZbdeUUHRYTj2cOn3hHnnZ+vbGTluaiZhr9TnGTvcfVZfBgtDWe+IIld4h
heJQ4B3WRx4DDgS/piNa+UVVs7h3BQXuseHfuABTjgOgXFMi9fMOEFQ+t0u1t520
nG2ukNZzt/Ikwfz6CmpXsdI1o7CqvInVqFVBfY6y8EuwzMrVy8CuUivR+Ya1XTcc
EeypSX2QzJas54ST0UCnFnzbTsQ5r5IVTxqAEt8rhaB4fl8xDhQGSdd9hlwKjxGd
MR3Q67AyQ1iqV8l8TFPKch4w/cmcqUCidgKLhp4sfyWHlbWGZNiE+Qha8PZ4PUPs
/CHnEg6/GTurXTA8A+4AIPXHsoRYmhR2tCSGFaImJdffmDTv44PAtX1DIQJuHbpl
ombXF2CGiZLWLLPordRYQfbJAlDk1sFuDwQc+0U67dNJ+sFDmn2ULgtDqKFrcJ8o
s+HZiyNOsSOGx3fLRAzVfE4daP3F+J8o8gXBCkQ11s4YhA3suig9dIsOEydWOVDB
8X96fWBrjHNniX73r5sNO/ZyJn4P31tYZzj/cnzIIfLsY2XxheGtXWEiAXGTUqBm
GCFkMpqGKvO0igTeBhliPEioatoNqjiPyfdLOT57XizojXOLOUPSP7P12sqsa53p
sfnZ8p6GvNSWXl1hJTDyFKL3olmgRub5yfrz+q9TcAgQSJsty0vdI2iDj8Jm/tT9
5ccFAe7PQi6iJEvz9VBv75ZgM4J6aMwu7Wv5oHpmjzJoEIb77HRcJNP9QH2GzIKc
lkv3fs4RmKo5FWUZ2c0H3C9+RnfY26fWUYFEDUCTRklsyihwjouEY7ZC6q6OTrOi
fdAK0tLMy0bRVJo+4BlcN1Gig/ueVUcUkrb1TFG52i29n/eXDngnPwg93pJYIRHO
hIfOQrXWPuIgU4TIoy3FrrSLYgzAXG7MsL2jKTU1DUNI8kT9iGecXSpPRSdhVeG4
m3uz0ZWUQi8txhaRMmKPRCzoAgtrs3WPNbgSFuTpL8ZLndiRS04mCHKcQkYRFrOp
r4/73nNMuumy8YrT5pqd4E0fvkGDk3bOvTuyJe7gGSmlWAKvnW2DCsQiTvedPojc
nEfQhnbmG2bBBkdJaTsYn52RZYRIBUPM2R+AsUgJi9Hi+hf7hUdckeFSVFgu5ANR
7VdIyOdv/W3wIxMcNj7s0RMPfD3b3yYaDIWO5NxBLlyQ+MQtmrHc5MzQizz6kHHg
GqsjbMWc0iwXU58NwAAa4Glg+EUsYRIYQ3aGOtjvIjVLNMcLT1BNekdMIn+rt+IX
zTW6a6E222I1mu+XSJvxreK7F69uZknYnB7vj1pObl0TXc7B0lX0z6igLDzn/a/0
6SGtdidWJCvRGy6/Ihe1xc9UNgQPswHn0RJTKimCVYAxESzHGbd0R2p6jNcjharg
2gCbwvC/SHyWuS3zMm7C0+dJV6U3gjG8OagfrDAdRFr3tNEL1QBbb5C/KPa7w0Pi
K0E+cLtLnSgeoxJSCX7SHM1eMoBixITn7wBa+z86ZI3l/7ZLGD+6RvX24E+QXp45
buZswJU45COsDfJNExFm36b5JGjZxUqsitzh/fe3eBYEPUtkfeuhhDup5j+gzClZ
nUK39k3q/Zby7uyTGn6RM/eMcDz8g9+Z9mL160jfIzkw3iuyM9440mQCMVSpXnQ5
WrTTSRgU0LNXV/kpaEPrpv8ZeEiszFjqURyNYT4aN4bxSDHTfFfO5w67y2tGoxg5
rjazbGQZLY8rTzOIuVk8ydOmO2yBdk8Z8sdFzmPQK0A3Gx4LkfOWy3YSURfiWBap
PmM4sVrTWbwCCuXxzm6BV0X8E+ezNMf1AZkspYaxsLBlTTlwDic9xWAU+N/6UOWA
iiYbANBjdhA6Mt/1de6m7gnpa/L/genuWgwTYtZXKAxhDIydSgZjJImWvt5BNX6D
/NC47niVJqf3qD2cdVXM2VctjB2e0Xh9EqpNEtHEweSCiT50FHRNkRXFLhfVI494
L+GqdRvGfBipvW9zh+KLRD8B1Ps1ZlpX/dY4JxjY0+TXtn0/IWb4fWpcgbgnICch
Ms+TQrlbA0h2cnrMIz5j9mbSOh+EaUqj99eECH9M9hGx7fQqYSZqo8AXM8wUteda
UVY5hCrTGE1v9M87nqIDAtHCZo21lF2k0v5r0H+qI7oahDWM7mrjF9iP80VliEq2
QK+o4h6f6LQenJ2pMTmSne4tFQFc/zg7GDxk+5QwSIlsMmjlBPjaaCzphuvQpbua
XwI/poBdjmKPihTqQdkYjZI+uOPWH8N1P5+ZPjleMCQX1l1qwsSgdklOEio8bx9j
4YvScLYdjMttxc9e1TN0bqd3IF7+0v56lR8yAKryWnXIQ5Mo7FyajX2wp4cP8RtB
GeSo7q1ETePz1TcJsud6XWxBFVND6xqxNNp5scgAZyomUeC9Cdsqo3qiP6U1OhVg
5OgEgeeyp1WVu/rmxD18XjN+NkgnuYrNn8tXlJNzdKRMUqSxdMPZxPJD60IosiL1
+zsJMkDG7ulOG5cCT38hcHXnTOTc6mpuRLLqIM5uObk2sZyph/L0EPNbSiaw4ir2
srGvXfKk13CzC3bbZQfQ+WmhgNenDc9b9X3zgonPw7AZrDJwoH1JriQdAm5cBf0E
WrDPxCOQYfgX9ewQdP0e+9h6ryhA22qkOs9oFrFNXXyXy4grBezUSFpeHvmbnJeG
hX5oZG92C9TeOD2G0bglNZEZf+H4cPxAblB+7fPoV3C9XPrbZzvDiEns+wzk3Q9g
XNC4+Ts6UDorvG0axdRq9/rIIEUyfjXwDd7HkBDuBRzsIs4WyKwayjF+IXgQOe8a
vMEa85vUlU5LAy9yx9TutLvBDpbyOjzjxjoTeL5EBcjzngITR1ObbOLzArheBEqS
82L4qYvB1Mtdx82/EUHLW5GyW23JQS/oYPnAqSvd12PvPx/An5mjYi67ZTTsEH58
EZM3CpdiHFzC1h9wG3DqW8m7vkP+ZELzT/mkJASRXWlj7Pv8kWi2gnlajcaIjSo4
ubhtN7TSMw8Ae9Q96ysbqhqz5AqiU7wAA5/nopKIEiNXDuhpFv94rSuTbheKfwEP
xeNNGkbIXtYHAUKynRffOf5zPlQBN5iiYSt3XtBVDqm1LFBBRzXkAUPwMQOpdZs8
RWntmQU3iaqvCY+wsYhgFOj+F2unvozbA3ykG6ngvtZYizymfeWlcpRuid0XN7IC
Sbc6v+tI85FFrLfdF6bR9tYrVfDrEG3XJ+2ThXt/vH1Pnxont7yJJ/l1CndiO6W2
DzUy5bHCAaWgAr9ycUWWUrVaj3ITVMuCpP14SvHeLfbC6809P6UzE09e/7fg5Bew
Mq7PHewYnJtEbmwDjTWs/gdqVpzUFONwU/m+vUJWoNStorcfOYLk/sJT7xst2lEz
u8jjGvcDs4novthXRTSSkbZQilXCFKRbDwkhaJffE7XbBLTuYoIQnBa/t1O+F4iZ
Gp05Tymq4ZM/J9FU8D8eW6WlwfdL6S9EbfiMRecP9ZMKQVb1R2dfSdGFwbmDZ7pe
d1evqJDk45r0UjEpmYLY8cNQjmm/g+4VDZ9UmS7qfOhc4wdNxiaqKAnVVhqyqpsZ
t+2yONTflekO6FSZv9DqeP1evHeD1bILmeWnXgcsIYSsIAtw/gjdiR1yrWeWMl4i
34BYwUGQPzx3X3N6uPh8ogXGBejqQsr35UR3VVsrRqw7iSzLZ/umy4g6Mn+4Vs5w
F11qY83BmAD+SCofjpsfVrkzt1fZnlxZnmFt9nfRMjTjwv/tXYaPfRVa2F6dRhn9
SlUdDm2by0S0UuoLUpH/B7j5NusDnmr63W+d7d2DQ7QSnOvmkzHR8s3csxUzuTJt
WtH/1it/cbSX8ascr5xut8Y9VZ2gnLXD+a64Wx4EAT2kXxAn1e1Rfolqkcgp/tdw
ZpmDkXT09UEac0xI9R3MBZ8buYsueb06R+GdyI2AeAbJe3QR+ZNTvFDSwfC6uy1d
O/1NbNEyjdYNkkSRu9PZzc7CKAq3JTKM7ewkA2AEpAj7EZUUVbGW/AlPvIXrBGNa
fBrv4EUrCInLNuBvZrRxOdH5DguVSGw24pUSTF9pmCxzFkTSUtQbTMaHp0lqG3Tq
8g3ZoW+UhpHvCVvqZlvLFtvrf27LlE34+H8BqUzilleO2yo1x22X4VHKL0+2Yj7Q
AXnBYV9fvbdxGkqwui/6z5H6vf5Z6j3KFqGL/nFoxc7QhsOE0Jp7kYndrMP70XEW
UjxgR7eG9DXjI6yEdR7OYBE/5MkHGpmQVb9KLwn6PlK7gbZV0XXwkP+SfuETY5GT
cDMQFLLpm2pu9JdVzM+TpLxiSWJTNVpIEGEfxzT9AjzZ4R9rBLjl3zz3Wq7oPx6T
LquttgisxhaZDvIVKM6tBtAO6tO6TM1vpqarxzxKNHM1clkxFtIdVp46R7xTKF3z
/sxApUniCD7q0RjxuuT1y6p7OskPsT+3vTiTTMOixnrgl61G57BzIX88BXAQ92zP
CFSLV6+xPA25kCIAvaHb539LhjZzQSpMdhqkwGRzI7PoqNR0GmhvG8uhBUDXEk7E
CVf3U8KVYsytoMRdG/l3/5xJsgfxuR1oybgD5wImOoFfXdryLN9Dr9vr2BoJ38Dn
A0xd8/tAjfSE5/dL3U75BIC/Vc0DIam7t/XNvDzD28lB1eygBHB+NzybJQQcqGhE
uxmoyT0Mp4GgEPmWXCe316CX8r3zzSdb8+jjB5d9JmZPSFyp/ykBYZsGUgopKyNc
0aYQRCqnIptL8CWqNOUVUn2a+/7qHJaDEQUFaN3tSmA7uM5hru86OTA9xoFaT2Xn
NogdRPHTjc8TlFaNEbJ/UIy0zt32EQn7OsZJr61+CtKxjSe8WrCrkg4bD52rZZ97
q01bWKJrXwth9efQh029F61tjhYNfUk5UH/dGS+X61+V7mI8Xb4Yfp3LNaC+mH4K
h9cCl1L48AckTjOrLCQVgWWYYMuTJkJ9DiDAMNaho8wiVeXyPJDJtZoLRCJ0y1Xq
Qf1MlNnoQ6KHvu6QYULUQ3Yid2yZkWfp57RXxJsCb3fgUJWbVKB3/l1QLqsjBHY8
0yNcIMDrkUHZNYvmxqxGnuT2xvZ+NpiBN6WTYCxvTaJDvyGEJaRKo+GaWZxWULuP
0kUJJuHboBspy1Zbv3yYgamOH1LhSqSCShWeb/cGo+bPgJlWciiWzYS4Uyc1xeaD
4aosTYI4bSQByCWh09a7H706QPny/b7234YvWNAsi+kyQyOV+ZS9BwyryinCbMoi
oicoVc1Sw5+7Cox5ZEeZUPBlMGefC8OnLaD1sVoWDndxUv5U8tN3Zf4ke3PnTS4/
aOJnhs5poyfkWGdkgLUT9MihYJbeI2hyuWXXJ/0yja9Cv3hvvi3Tm4R1jATLtpSj
UK/GiYaKECFjkwMYVxuJr9K7sYa01bkRTnflvGSt4QtBYe7dedn/q71Qzpnq9e5A
SYMK6Il4+zGzdJ+0PbxOagLbhoOjexTDstVI5+XgZWlcD94NFY8jXdjHs9AnJhip
LrYyLUQSeOZHMi4PILxvGJc/a78QRtaDeIxXhWoE4gw+68X5gvsIIB6faZIf+Ro3
LUKKdK6KJLRfn6t4sTpH9NSFHzOzlPLzF4vgXThu6S8wsZmK9psJkNjumEbQrvBp
XkwAL+88TtRluq3dLEC288DORai+NBsI/OUMjb9/JTdLwtbjsqMveKRyjfbdjj5p
3Al20VOzw62RpEfZtKLcb+8YtePPw7VseYrPspbcMSyHemdpf5iQSlsDe+YbiLzv
f3Pi8nFXxVqPjcWE2PQvl7numGpgr18oCTtRERFCpT1GU0VFPNWOgGZvxd21bkEM
TZPPEmOMtm/IoFeYLKorlFYQWIBe3UUf0i/MzEZADVBezizbUqovDy5cvP77O1Us
6tlmUhhpGrTvLtghGGSCKfOn1KRC0d+3mnsUVpf8uxadxLwEzM9C9CSNiZ7/eHYh
9M92YLY6mOVo8c12bCe1AgxcLaMw4tONIo38fw9/Jsq7jmORiT5cnW/LUh7dZsq4
afqnBgxvLB3hdQJecWP0GQsSTXKDYmyX5y6cBt33XCZRmQJpa2nq4wNJ9BY292Q2
GIcc49q2OEYBgLxBfYTlO9TrJY8EqhXmHZ2jHXG4SbmfNRdLidnmPGiFMv262Dxa
5NwE1qCkzx64kCaHY54DdwfkNNkLHUu7LrqrZQlCZd2Ug6B7CboMzr1auiybV1Kv
1MmE+guhebM2F/KAtMad1HaE9Sd/7NRkPqVbuhL75mxdGlKPf9unF4Ou+I8EMbUF
9Q5rYg9Vvil6h3U7FOIEuSA4Ge/LrwgoTZNbFu0J4i+nM1Su5WGaoRACho8vt+jB
DtJURk8GYcZr8T4oJUPz32f6CQD1Of+B6goliBYSZwiTi4AwZAAEw4JH3PLaUQ7j
gfCUnzlSxXewjm5XpAuobTnFneWeY4SScPJyJa7FJy5q+3qSq2MxeQMsbeuzVOQQ
ss4kvPvBlkFWZtz75WoLA7t9Vqic9sBwytySDItsJYPcSY5o4ryRqIPLe+qHxo4l
SVKjS9DkaIIQBylAU+QgGla4ZAmN5B4slUgVKRdphtewgyY8umjxlqJLqPi7q7s3
ZBQ1Xni8kbvf2xNtBnRwQl36z/9zY1h7QbKGaZRy7TK22+4mPv+BkETYyfkBk2m5
eSkYSD1CRwLWlILB901UJRfqLhSUOWVDUg/51xJmHeqGDq/CY//0EaffW0JRKWcb
imwAkNiYq4t+1B68QymS5nohdCVtjVDxwRoxnNohOI26z0SIsvB4TqvTZ8DNjBeq
gynazEtpehkeSnBfd+TJqRWb+yOltkluzljNRPtaWi8/6lg997NVuAwdh8LFUDzU
l+lsns/pP9HF8M95eJDYg8cuBsu40UEif8ug+szmjOUPzy5EWELZ30lqeLZ8/WDL
MI8XT2WMbxNG36rSu7UA3uCzTkRafeDZX7iGx8MUL6C9sqIo5h3UTVIid/zembbE
8jVKvL66p/MBUQS8daF3a8BYwgmqnYpg/0c+U299h994DcnMjn97Orh06RLgM4S7
lz2ybTSV+CM2mYhkcs9kxwS/MjXZkf8ErrZ+E2YuJ4NPUg9ReZJqD1uF4r1Dv5hK
BC/ffiewniEslwWkkGyJTI/UGUoNoOJsdFdkB4G4hwvgTjmcdn1cCBUWvcKzpRRX
snhWfDskOLjGR39cQnnzayE3s6oPQ2TZFkVZXgkFzABcxZCxvtGUtX+0NkJzgIVl
qXHLzF6Rph7Hyv6brFN1gr3R60vVxqRLIDKzZMSKxGWs/3VfhMnQ8KdlpDl9E/DM
pcPDSpQFqDcoZyvK6+wOxoo6hfqyu209GilegEMrP/oie2AMHeytLA+77Q4KTbkC
mzoWYgq4tt7vdmieKJtweCNeNv0CjtxP/NYKkq9czVQQOfRl9Y3V2SvtVHUWo0ba
LqjPNXRRa82LmE0OkMc5nS1qxJ6zJklagNPqffxJr1vKhrJfMglKU1TfpsLLZukd
hsFdKOjBFPxIayAan2atRe2P4lUOqiMXQcd3rVMWw10qi+YbW7HA59ull025QQvc
RDMg85lIX77G/d0PHPnMs2LIVyw8k9cAl7Kqn5HKgPNrVEnNXvAAxqTnbhp+nzIn
9iF3VPio+P6fkl1XtpUJKWPJ77o39RA0w7v3ExkZ8ovbo7Yzqj7AmVOpcfvNqiuP
wF6fxNl9z2HW1xAGCstVA73hiZYF4TT9AKJnzLoPRsWSX9C+B/hLxgK1UO/cn2eI
bAP4txJVuEOaWhWeqXonq9W7E/X8a7/FC8cBTuh86V8WuPwGBFkMtdylUkGR4ElH
1lSz4uQPBH4R3jKOrdGjLTYlGia0b7ZPFgGV2qkTQaWB4Ty49igM97UfCK62YXNn
9Dgc9j5xRy9oAJNIuxHJkQAdSWZRVhZHq0IiUFSqGI9tDD16AnnBeO2CU3FKTgls
S9sE03V+3XPe8epS68h9hds4UoS9arEbrQzB/2DIV1PFggnLlJb0vpWICWOkgiXq
i5Ya1Xmg4cEZrLB2vygEo5mfyzIv0p/L0TAIG8t4N9YOmLgmmPRC1VFK1wvSYwB6
ml3ZgPa6rMs6lyI7YFirB10BOcJro2AO0SUyOY+ZliMWPEusEhVOIJaBWkMGVUQE
YT5vUCoEnCrp2HksqLXMw4ovgGJRilhIRSZrZs7ggLlie3y6cCEPBuyNXz7/dSUr
UkiRT5zpTBlOvW6ctifchMNncFGofpx4HLV9yuFLxVtyDnqk9HZ8gJTigxcZWVIp
33wEHuEc4tx9QuFusnVVkW7SV3YPxh7PtYKHgTlC2xH5MeK1U85uwmWOf1TTHDXQ
hmenhd0qleFguoBnQLVDOO1YrlV4DzFubXxXoaADe+huxSCe6luCNjOHdVMQ2dwQ
C3/OkDCPQLAZ6ZVcYWW1xfDUpTJza8pVBf+HXjaZ4jYUJpvy44sUM45phwvg5tcI
NTOWHziVQEiHxVB8J/dQBeILyKXaiE2VTDzw8uuDQOXpb6h1yy/di2Znlve3UdcW
MLnxTtUBrIT7hnFbDK3+0Rte1d+QzFEptCImljnyAs6fKcJ2Sf3IfYW1VDY71rKg
TL2yB1Kz5gmL1vxxBhUQ0OlHZZOEuNgDNvMMcl1kvvVy7XoM1YfDPmUZkWGSHWZr
V8QyfdkT2imkHcnHASk6dgjgfosGThDo4kWHeXZAnvsLbBcboS4iyfhPnh8KHkPK
APFcFhpNX680NCGLHupDsUKIKsn+3GRne1jE3qCtSzOtEodkQJ0yfZwPFrkZx2eC
1WsxfNzCaI32GE5l07W9qtw6vyerxuKqL+Xd5CSlfV65NytsyDAjy7qQReR+FdHX
GcMbtbrWj4a3WwEom2DtIQx9sKUBP8d/90zLbW7YWkDphRvBNGa+P4qYVFa6Osyg
Pi8w4uaNGGM0EcnQjP7yaNSWYsDAvW5yUG80lEpWWutanhGAAtWmpt4Dl0rfinOq
74j3ebfSlCjm7MfWmQ5gu+gwG+3qSbYiD/vG5Fw4KU4DSLHuKIUkEXC8fuX5AE8H
RDIA+T65U5h/c7mN0mvmfhjuQ9YltnysYkYv1tEcrYTQkkjEA4ruyPdR2kTAlQ/Z
1VC8D6Iz2WEmam9hA4tWHQAUv2q3t6ZTe7x1hfSarKSg8YImKavTTjaK87zfPbRJ
6e3DnlwKHpVbwkYjpqGGE0IVclLdJQg0ZXU7k2ZvWDfovEaPLP+SogjMO3Go/rF9
IAevajYBQBChnD1Z/IBUx8PV36uxumJp1GZ1o+ssYNt1wd4DUQKNwQ8pitT9g56u
iG0zxTymFLhUwavyZ3f4nMhct4IJ5lVlcs13MJ5YuD3k3LH7Hf3G5kRWyVF+Ep+N
wbbJ5sEetjs32Udc9AGIVg==
`pragma protect end_protected
