// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e3AKRtvko06xAn5SRC0BCC9OzrHRCV42MCb4GFS3wApp48p5PPzFAIBv8FXWt9lu
P/QsJCSiSFC7svxAVxg6dsmukn+N6K7IuPMiFven2ciFQUo2tMMTdQXXIGdYJaNX
n6rMtW/xCt0rk48/QFbhn8AFQnHcVX9vvVZsQu6jMPg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 180912)
bESUnIdr/vhlG0uLxgcg2qNVJJ/rE4bf7hmRoK6Xa+UPFxpp3+XFNQIe5IXRVXCX
PJubYqdYNLlSFqTCnjIGLGbN+LHQt66b2nTw7HjFcoHu6Qnz6xcodmfJxJOwyb7M
k0hrdDh5mfChXZ4Khrh5kdyMdYyp6l0EoYXgtcHCIsfaagd0LGGbOyaVJT9xpbQv
wxm7iqX46STp9s7drJKegQ897AL60CbzfbUqSLqBDzdZEBdlmqbOY1sJk1uzyZaX
PQuAjRUtWRdn+1jFvntDjC9U4qhMHsROlIhc2kAJtffk0cHlfkJ0kB7gIB+/xsad
3hTIJPEGmC0QZsdC1LrIWGcm2orbsDMLi1+71TlsbZYoN+6oEeRkeZVQl2ypxUKt
Fad0XC/q1YrF5FnAC3Go3m4DXM+4yUPar2iKjggLzfTyJ0mJ4KnPaxYhi0enkpuN
3hyi1M87ds3SidKUpL48p8JAqEZuYazZWfFaIfWHUGH5UcyJpgz4AyGbRaOpsBJ0
IogrMBZV7+nG6NMlJqNY3IY0Jsp5TaAkYreyTJNJA0jRltgJGdoDEPCye6ioHC67
boK2RYYBgSGiPFzeQvflw7c/scExnxSsMUYJZ3QeE8K+nO2jPSs7VrTcW9alEDG5
ackMooD61RbRKhXSeC+fk7OGQIOmLsdUfgJiO+eNVEi2o6NWMyhv60ImqP8wWPz0
wcCQdjzT0+R3EQIgbtVt4MWb1ZcinSrfMJKm5ivfzUonuQhj0J0NYLTsrO1NLwB4
JsSGko8dNuaXS+NIg34aOUb4C88Un44/v8yrv7NehnkV5D1K8N1C/tPfVhVRF7dt
KT0iJV8zcfwGRKsm0d3LFrVDxIC3g0XJ4WDegEpa8S3NuvPdoteL1z2oHXwFMLgX
5IUvITre8Rb0gQDG0t7dHVno/EIHYXu3cdN79RqThh37I1kIGEZCp0EfbNirmx6W
zZOZBvViH6vCI6X1GJzIIn4CX6hJWxIwNXPkiy/I+1UgaZ5uV9QFmiFZ8RBwIKrq
ZVT1v9pxf8bvQLvoTUTzb2akABi5jZm7Kx7e/ONMcVagkNSWS/XoPsNNvao4TIBu
PVLcAPo2Q9HYU0He0Dz0YgBYryPBCb00pS8NeJxXaD7usC0e4KsfrnBZUhnYLQFK
Xfi2/JrIHE0XzJFSPDJwLQbL+RIU4TH9oetnsfoVHXmjv1I5+no/n0sxHFoI7ESv
gnVbxdrCimXptf9h1xcAuzsbfF+C+qWHQD07P+aJZ47IUigC2MlFTjijCqMFGugL
3rMg4MVREvF2HdeWtBbNmHY/Ap0x3fg1LiqT6vwd7OeHSjITjKHC41cp7nYSpeLV
Vt4hn+sMwi5e165/ZzmrhiQKgoY/LlS9m3eSk+ALYJOhuIqCPZxfcLJsq6toiTF0
egDyW8y+S3K/2xURfoPEXdyaI7nGNTBHiu4r+XxTIXbpmo42sgOljX+SoX/CY84j
wCjPIwpLS4f+oWFVZfp3wLQ9c1a1z3nhWjBDqzM4y914L34aJBKiHmBQdVndg9fz
gtvgCZa3QSrxydklNImTXSfQg3pS1FqDNLccg0nfMD6iV1i2y1tW02f93htZXlvD
dSIj9DZQpFWauIv9N6v5lyc0qYy51t9FLAWwDIvUdqzEWhqdK4zXTinaeeA33Xsk
LQxNmsvK/t7YhBxPTUQGkiRi2Lvtf4hEyBGPJmWhZVizK2QhiF5Oa2/8HZ0a5CWd
Vj0fZiDZ+e8DJ5CQb2hvOhpphlqRCKutsY+0oEnnYHslwoNtBQJz/NdIXP084ePG
g5iNPCdd+/pKxA+qZgbXqz6HTtCmJ1s2fHggUACGgNdtZIg500/GJQ1RBWmKLL+d
IlSLY9n9PVj5o96Yt8xRzAgUQVRqPd83EehYobXX2XbrhHtOOXJPLT3Y5INsrYpm
w1BZPD82qiAEatRhYn+Chmy4JDZAAdgTcJOoBYcK/iqW2/G2FM5p/6nDBYKBIy7r
ovXh8oeaeK6hBojGXHi2dzmH/HJ8ZZKMaD7iRgxJUb07Hdxs8QzT//AyXxvFAHfV
KL5rTcuiI3zTWRWVGj39vzroS0gKlEazengSvqa0DniOIVxQgHo8O2PnDjdnG72P
unLVJ8Qxo5yiRaUXTlg/obmrsdo4l+/zgZQAjNxUWWWDPJ1mEf8E934XJ6sSiujS
EOarLWNCtoZHIEN64CAVo3vqyANElulZjXepLGeNkqttPV1ZCUJQ0s0my/x8dfQN
Xk2dg8JX9j2DYS9NK0HYnA98Ey9XTUU4+0b/6TSWelooHUx6+oqLLF3UadPMu2Q2
00D767K741vTstJ2s9OqXJLc2cXoaOT0pmJZtZdtpwR8Ia5p7L0wvKrU4ekJCL2e
z3JttDUP+XC1DPAr4dmUWi0/j7iniuvEmAj/G4Rwg21xkgbrMJgOvtuHK50Fh1G9
YK7wzgg9eRP47kOXaGCf+qrF0zwBCYCVhnVtaUJ+1C4wTjkmy0665kxPcZXW4leo
uhe7Tf6ND+Fjq2ABnDel9Oy6WqpOxLCH9tF2P5w3ql3gAC3lyUKigpq2A/D4pQxO
YyDxhIIrVVFCNwywp2WQNLWOxoQiQSMSpBrTYkChUIZJWLY1K9B/UGH0CxDGmVZR
D9N9wPUhIDhE308v+q2aQdPbB6I1cG8WkFCcoucA1M/4LGJmamI/B6b5+YAVt0Uv
QcS1iKTyMz0RDkkjDMz0m0pKg1229uL7XK+4jPtuQtnuLNXV0mIGbItVdjVGlhg5
Nmq+D0rV3fzC6YbIdPeV73DTz8yS0oGeLbMhs47ZpW7CrE/006wXYGg8H7PpeLn6
x/UCdwhyirF2ODMiRa8dMTE2/M4sUHQ6Np9RPzG1yyGq7UYgtviL984ULNv3BYxl
iT7mZsHYWfhsE5V+hsS/85esfq+xGzIv18C6lyCtBtpoQHgAMDBcz27oEfq0Hh8g
3WyjLmDS+6gkeUq/WnkHCAc5esPsld5H/TioFL228wI/NYg+a5+6FsBcgrjNHwxu
GnWPc2iZq2j2FSkHa4M5qW1m3hE7+2LUZgt7ccwBYhs30GUOtesKle293506RaXO
b4uE/hSJFvPayhBfVxgpIcsW99hKmq2H+ky/BLLs3bGznxRWPGs6hrf1GJqcriCB
IOJHZ/GzO8O+2wERXoTVV65VuFoSYwdF2edtd+gy0G9xOXT/eYDb5NsZzlSc0xJ3
J454wPNKlzydlURXjb8/qv7yqQ4lYCWse6k9e+JvrzBas9GhAm7chyiHXPvoHZqn
5oeT3I/ZShfj0hRnDYhRKAuwCdieglZKiCBlT27oSYP+0xESli8W3jAIDpjNSizU
HITVZik8TVEKEWx6U3OkUmI/frNq4ZOIT/SMmvajIbTzIMRa3fSYSoRgL2eVsERR
fWlpVQ1T7L5UQ+YHgs+kDSzxBSCIfpKhS0FiAeLnLFxEDsGqMMtvQShOjBYKV2yt
ZGMo6Q+Oyh42FdgyRjTQgsIaKNeMF/IhuCFWXsjtME5fi+hfyJgvA77qCBVWsCHe
EXsFcXSgqC8LtlskFHnSHhHbr5JmYWQ+UmIKJx9n+R4ewJdETt2Z41aa7cH+mDUi
7u3ArJKmCC5C1vypghp4WWe1R0rbE3Eso1+nUuyyiWaduMFObitQdHrz8wasdI1H
pD33B29APg1tqlT39okpsRx4qMwCJE1emSM5LF6yahPKTFfJyHY/BEmwvyyB/606
RUcPcnp8VeInl8iuXR8Dxz1D5oLQMdQ2a1gRHKFJ5JVe4fnnvGJuxWOazOQOVyRB
YIu6+NIrE5QQnoPP/Ikz+dbSQbt5QdeW+gigaGbDPnKA5nDUX0LqYbpv7zF0NMil
FX/hi0jYpaZGp+wIJz1tE+UfZVUekWnUHvT3UhqiXvwxlWPudNAu9Fl1MdbD2Pr1
CQfmiXacKBXbh6Y0MyfCpvAZF32f5T9MFYE4z8+Cy+oMDvNGb8pcSeS6ZyJnZ1aI
i72o7AXVoS65tYIq6FzQGWnfR4LDZop+2sJJNOZqKxqLpUif/Yy9S/FuSs9XzK0M
sGyAv/JhJrwXpQ9tPBjPP2AiKcQjjHlrc7iDT4KoMZ0lFHsq9eTepHL/b1Cf6twp
C7ladQnm/vpkUb4DKW5cm9LQPC5qP5hfPq+7M6T7m/ZzAxPbDshA2TRifCU8kBPn
q9qVvvv1dkSFqXK3na+pCX/kt5+M302970cUz7dsNbQkmw9rvoebdGefR/7sgIpg
Sf/2OhUe8vlqqQ6sROqs1fjqlRoPB79v2xef3UKqe7Nn1AVZcqikJGUAuaReu+aU
5NU2GBQSry7XywzBrQbDoO38NZHPst5sTki9Lb0gbExPqLdjW9W0ng5FAUO2CYzY
E4SQhB1Jowqj8xDjHGjA8qM+pvi9ncRLlE8Bo8JNcrw0IyT9EoqSfvKZP9tNrVvb
2mE9GEUI07ae5s5+eMq/3+nl7mAIKeBNX44oQdf18w1v6CLS8zhy1OzKTKTihOJy
JvaRME0UFGtSL8nLwDKsMvyW43xYq5KVVhvF25OtewXV+gkW94zIB86noNywOFLS
HoKBfxIPQDP8U1mRIfGahk7FiuvDn/rzQmpm9QGsLD8PqDu/YsfzNpuky1lzw1lF
wpxG7FK61nPtQyAT08qr7Gda8aLtnK5a0QGGWDXDEhprPKj1Gb10ZRrGvYfRCZp9
phAlNDW0JtCaHV1rbEg9aQscmLU8bjHXna7TsyQ06fbG2oZxdBRlxE5V3JyxHySE
pwqURpY/FNxHoqNF/fWTw8GwrgubypPHRzJ1LgLlnrLKbk+yonGzSDGA4TQOeSFr
am0v1eBOkxqk/b4nfWK8VP+VRnb/P4O7BmHy7pU7pOxQV+HsVes06KikmC4mX79s
sginjiixfKVmLhW9sDava/MpF70URAM5CmugWxcu7TI8ZmxXAVbJE5Sw/Mp7VMLD
miRWluiy2BPvI7wrY2aMGKqIWdNK+WcTWBctcTKr8cqhLX6seq8QP+OUxjP+yahy
lvmzunqohFlzcsS75BtbpfjuxdjrwE+uHJ6MV93hF+zj7k3ADSep3/6oEB2sOv4P
Xyg3xlzWg9Lu+dPH545bAruhEYelVe8plY5RVozqfAUG2PywM3L6Lp2Z3iOruSOR
Dpnvo2Ruqvu4OeDnVlbR8GP0psU0fsEHZs0tyvhJGZBBjb/VlT8Q+/17ftw/Xjdr
R+UWNEkRksQXcygyhqGQhXonvVcNl1g7/e4NlYOu0tiRKXDnCwIBrXd4YFoZcAei
O+ZicYHV85X6hydi6zLgP572rW1Z7EtrwQfg/i4AUpgVVCssNHLMpZiLlaZDE2G8
TF9EzUHWHVY+6iYb/plzbI4mogvP1t/ZjsfS/L+J/TN233AXRB/zzAjeUiQmtqbc
L8VNFgeKhhh7TUNPp2bVz4NH6etAZIiIq9DJrghsnZfa905lfoV6BWtU9UBGzKsY
o3uAEA504vupGz2ojgkJpVx69e35qPEB0mdA4zNno4ImklbFKASXh9zK8PfC2Rw5
GaSmPqAEICCgrSojFKl0RusWhYo9Y4mDgmdLitBNFFqQLxAGnzZlJmL8mT6OMUhy
G4NHnVAQ0FxW6OfO/JUzuQkUNeIkBt8GP5S1OgWoBjSiBHigO91JH7xUGJzgHcip
pfvSbUq+1HZaJBwu30yLo/vJ0fsDvUMOEQ37OHXk2pOt4MxQGZ71sHVFbbACR1WC
FgRHfAou0jifb0WNqMUuQKlSpSDtTQo1jRpdSnxr1sI37hwT7lnRZ764sU25Uxuq
YC61qiDOOSGLEFKZOdZSWqM4BQUzXnNT3iIe/MzKX/r0smNM9VXrMT8QjwTUMrK3
VDtDkUrt3+jADporYWWc23XZX9jPIXyzswoYO0fH5pOuX3Dbo4zXTvaImTSP7lHc
K0pdbfoPNTQNORWV2B+XKBdN3Tp4EuEDUxM+KFb8RnNGlhPi8RHoP8MOiOCLirH3
N89QACuze/Bef0zGD79pW0dFRLff1Yq1Iznx7l8M1n8x7jQ/nzHNAujJ+Q1EINwP
+0UQexZMXJXByJWCBy+DfeaV1QMAnLY/OdP1qr6r8npMvYHfuDSxwGjO3+fPfI4s
warT/j2XLv8kg+deiIPVFoPjlPdetjmHzrxW0v8i16Nz/BgJ3GzKIlvbmVthqpNJ
4MXOuTiYxamRr2TpUQPdeGbg1wsI5XYY9u/Sgi+bXcVq8hwjWCKFVZWn8jnMujIu
7fPnbXBV7Fg/u9j/W6oDGKgWwE4a/VPBA6Qa81+/SwP7kfSgEwy5ObnNPVOdpbcp
ceF64VWTE0oXreShlNtkBQS4+bZbyTcYgQ3E/pkrxjyXloLhhfTzOjOJJ7Q5KTvf
MT3ZXLc5rj/m69/vDCcaG0/6ddyUJavXPFkTAJFbyNJ60iVvGED4kp3ex5Ygknls
QoQSUd/BV4PBok+q0mwFKA77sxy6fROLEPGgCnvkXnONQuzeHG4tfYRaqTbaga5H
ArEfEUFgzua6olG2fiyXKWZtlT+pdns6/228vhKt/djcxZ93fAoJ34PI7H5zs85V
pvjJlLV42bZJekhO9sMimIN6WtfcJaPwMz3YeUu2HO+1e00Cf5NTQe8+80BFDs3L
3VlDMPak0uYxQcHL8zQ4UQhsWkvY91QmgPBBHIbA8ssA3am5LkkmVg/ZdmoYLy9a
RZnmBHjquEA0sNHRhwP9sIe2H9SZYwIEvoFXYqWa51w9dmCdtVNn/wMHsYbtW4Dc
4h1IGWon6iAgHe7pZExDcpiYJ1QSfMVIaAWxJdxbIH+Z0bu+P7sroTlKE6+z7pq3
zYHRTvKJWTuPyhnTsuCpq8wQNhgzoD40ocJAnTqVDaBMBlkgJ82DZdj2CxScBJIk
WpiCmEd9jiQwme2nZdV+ixV1SzPpfgoxSGzLp4XtS4CZjqYrFm9ALW+WaWjWmyko
0B2/6y7QGikr8FNclznQGtyMKT5WB9+IdTo2SSFI6bfPDquPbX7CYWA91gcDE0OI
PBv07GnEuXuH3MuDkrRrR/FEygKYI19bNR7LSTEJdrr9va61EdeMpGH8GeShowMp
pCgELs4poGBft2gyd2t6dO9s/Ej+g/G5rxCwQ2uSFt5umv1FG7wIh2SLuIALnNaa
uPj/rygpnKSaOjaiWssk8SiFbAmTu/xoez7O//9ailPlhDLbkzGbYoIFeCm+rHdi
WZKXhfbyhBDjMGUr92IiHnKwG8e+rbtNlKYOvw+DivTZupBv37xpqq9Cms+drDTY
/+WjM0ddLp/wkHrlAvj+HkLXuzW/0yl99noR4mxFohSKx252GcPethktUg3ZWvsc
axAtXZoCP8Yy82OLdq9FqXM1peg0vUtjE50ebXnCYflpvl9LUrlw9CbCJk5DJI2/
CVsNTg7bNu9tvQTScZsXzh37uKHpXuyXn4eFvejP/Fh8KNMB3A41uPNQt7PERxl5
Kc/wTRp0g9OKgy5aLGyuA+WvsJif7P8vSN+PWPpH9ytyJdOqQn1YKwaIudRol0hD
W/r/1xkVQzzdcEpS4p+7esBoKVkxQgRNxIOejiLZXKBkbh1TOCT9eslZv5CPd6Ze
nOqNTx1s9pPHp4Q6OaYt9EZihFEEuL9PUI8t3RgmbhP96g8phNbJWODw/G1zPiEW
dRXvT+6xtGBvMxJ/0YGacHwH1sglIzNoL4HHNTrj7Y9+HCa3n0aaSYUpyGFbphy5
ZD4xRSYxRzD7pg9Fa5VmD0paXkP9nG1ntWVyj5XCVJ6kidDY14RRuxD2GV4X7Ww9
9ndeEbrChdFzjbQN9ynSNR1mptZ3Tj9+DdYBgT9WSwFKswgQXKN36DG3ckBbFUDr
sa0OOhhmXTbeF20wA+kfiiNBPV6Mlx85SmZgJGxKKgQWnSA5ghyH5rnffwPbYSlV
MjkGTA0Cg6HwSrZ66D9/0ztUfH3nteNran0oQc7QUIflfsb8mob2c2ryaBhsltct
lALv5zOnMsUv/dr7bEYzE+vEBSNqiY7zgTjW6++P9XpumLLE7mjUT6Yatzc8HVOS
W8RsMddng7cBVNIwaxih3wmkNO5tjFvdjNchM3xiYIlc4w8J+6Rn+6L10LEvXd5f
gSGtzcif0ybGIuaJUAlzpQD+sCrhxL7c4KnCWJNqkwQ+MSff4pY0ksrY0i00EuXF
bVIdx+2omS0QzrKr+7bl5IEBqvb8yD45lrLLR7WDrGhzadMTBPOLdfbzuJvh4RDx
qqnWFL3ifz+9YRLSmOOiaJaYyJ/8CqpOYoJBaK+vkDUyKBuIr+hM+aaRpDZDVIFi
4pDtS4InleWhqWnmVJOrV004uG1qFFpnjKR7hTqWjsV3P3XvOYqsW2vmybzhZWk3
OhhNlh0i+KUEj2ejmh3TFCwLCgEcizbgNXB9zIAWbArGL+xYXtFqNi2ZQANK9bS2
Y4XXfSxA3326O6Zt1S4R1evv40n5Q2AXSZQnSTaCF0CORDtUQvDTwH7jPxcowHrl
pkODY9ke3kmN1QkO6iLmORHC0K32ht+KCHFf6UtmPoGxtphpoHRuwnqtlXAXtMOg
F4nMVBnm1KkC3N74KoK820t3gguonQfaHuBoEgzM3O1ZT3e8w9NzhfB+dTqp6uaD
4cFcz8Xp1CvHo+YX+ZtTfXh+Z5yRP0Ki6/1Wn61W6gGm9jFEYIYc/Jkgs+BUwBCf
WP4n5NVlN5eh9YKV468j2Aw+FGeIR3m48RMQxs9uG9mVFmsd2dIJIxv7AyZ9hTOg
Z9CaDa9iTIllDdJxzjeP5tkPlrOOat7+KnO1DfyvbF8bQZedRzGgCsM71vLgwYup
W4rpyrbBCcX4DxYtsZX1pd4B4D44qundxcAMor6u5bEzFvXrLORNsNTK/+02lCse
Uq6nBjseFKIAnLXpRbG3sIM0S9Y0yDczdXDJ8NHbpLGbojWu8pkyR54tvL0F9B/B
9DPNQipw6bW96IKfSarNGQWyQnKa22Pm62dApqNT+Irn4v05a34UQvbHu13x7yBy
5V6TPYHVS2V14A5LIeqEaaP3/HYVwP9xUUIyFnX2woJDTnhX4Y2JxHhXfo+yAhBZ
w8r+TSR3ixfLMiXvvLSKa+Qkza3BaBuR4rNM14s63EX6AOqQ047D3oTLbAqH2eXt
nTjDQdfWbTxyYbBW3bg5jmaOC88BBPP+jjyUoEiak+RnQz1NUlkL6wtq/gUNkctP
XmhuDu64ntGoKwmfpgDw22/C3QhjePitI/Xi86lm0epsmrHbd7I0+wL8sl1g1Hw3
ljPfqY6vlGNOWgBWhJrmXXPzUvuqXhMhfRDl9kHv5jH2MshyQUUWSJ9u5GtiI9y/
WxO/e30cXIJZfq9PAm4R96HDzAUUuXHyI4yPhofpdP7EPNB6+3ZiqHsJcwETcOfD
e+BZBpe8N5XLXYAJl5WclOOi59QRCBqIU+Cwljyb2byZVxR8R/24tpUDxAc597aU
vvN4woIiCGNdCfkHp3xJmE+yuyA9zZneZYv3/VeA15qCGUomKrz+VgrN5m3mD+0k
dRAe2tTdy1GbkzjPviK1g7p0XxzyEAOwpbEkdjoi8qkGk83Lzp+viZ8oXHxEZtRE
AeDGnrbJfS5v+6h3BQ9gs+nkSJvJvw49ide/hp3H4OTCsuHncQD0wO6gR9XyrYjR
Zg6AoXtrv5any7ljaeHUEYmjtHGh+Uoh9Mu0LpwlVJYHxjHu07PUsVSLEvPm+ety
MFvhD7rKrZYaImTVm2XGku7XW69PEbiAwsC94IWupvC0RszEmIgqsq0T+JKBcTQj
j/thU+/hrJsc3wNVSmuoKvNAnZitaHV2b2ZufmAvaFPjLQ2skHszVJEXLY5+DjIs
phEVyyN18Ur0QDDJVjlQsjs2MCIVVu0Hw838RPrazLSJlW70EaQhRivvqVmB9gGj
Jr3agNDMM2oAw7lsRUocG2vOzUYiYrJjQPX7hqfOOzeIUnvGG7w+piCXp8nni9Za
LFUTp70Bb4so8b+Nrdbj2lbXswY6iUKiT/WhuGiKy0//s2zNnfjS4w60tIM32Eiv
Zv1dVDdBkFosv9waJthjp/vYpnzQXU+Dz5I02/WRG7NCjhAqNFjdDq1IEIMZFJNF
WX+OP74wh7JIcdFbXxN60O4VDMatW5rQrHrKcBDtIuoJuCpioaSLd4KHvy0roB6N
UUldOCndW9Fz37CMp1Fh204iYq6v9LogVbBNxIB1/pTR+msklTpXPAlqY+LSXoY4
d61cISsnApYW7SSGRXGLq6akArkZnTB/1rx/tL/jADF1YN54/CB0J8vAgYE5ifE+
CfuP0k2D8xQdLk6PB8ouEW1OMEzehT+hbHjXBu0eb+ZTh3r3BdsqOHCTGdZd5sh0
bFOaJuW3SENyBXIdBvIUvT1MSPTE7HfXnJ4MpnUQ21J0g6IxjZEjsbNHl2txaMxP
1A4fuaahg2ffV3412lMiWdM1pegaZ+ohKFodO74YDr22qJtuIkMSIg2beYeNgCyK
STLG9mmNjWpW/ddQpDegEbKbnfuuvBY5zc+GICOPJp8nGwrLDaucsgb6K4tGFsj1
CkoauTMR2KTakJTvYyyvR4/N1nH+TPLLywYG+3F+Qjz+n97B8AdDU0z8WhHLHHTR
wVdlwfT8U59sGAo5eHNPmE6MapAqkihwo1cHWO0k87OdCcfYDzbey0RaYyBSIrgI
c73Du+guYrMPumpkZfLsFnirTpzIgBjJDS/J1hQ84kD+B6T5mAKMikGIu3Q7564T
CpHlQv18Ij/+x36pNs5/XTnlf9sPoxV/4WvTMaUdlrLxcEOyikysfk/q2+1O7f7N
3M4qcZKxQ8evsATrUcv9P/VppLpG+H+l7ejAF2n23sQ9xRliKQlYVQbGO/Ku2/z9
BsnUZp+V7yk/jQSV4LS3wWyW+3MLKSW28Aq0JqicFcaIkHmxYgu1XphGcDcJQJlx
Vdw4rboeP4H4fPnNDfBgksCXoSuscnfOvWG3iarhUUKwfL5K+PVgtlhBlLteceKO
JvSsw4586G2p5W+b+7miH2VSymtkpS4xexjsoQt8W1jD+nLJVH07YXRYpYgZUsfQ
uU5/QamX5rwdQDnpK3jMZ6IpJcgWYbRN0y+yQmMC3Kv8g+UZkJp7gXjKxC53U01G
jFWk2IH7lkLOiSZ9uiVRNhtHcD3zQlqL4Rj8UzQOclXGFOBMhyhoGP8/gMjaHHRX
vXg8cyHwf0cBIDy/fLdANgWYeajmz9qim9/IfqJcOOXrjM4f73zt+Qt0uD4cidp/
BA7zfoWAAYkCsxgVCNOEL7Yylzs44IES7QdU7c6nTOl6/FFyVAXgJndi7OqEaaPC
IS+33ReTKe1OMFd81ODgzyuiS70Xx2SjBo71W5P4fx0z0PPG5zckYYwUvtIZIA8K
uaXrg5vzlmdC3rAo+b1V8rsS8OqpZMnsK9AGXxmDjdLqJK1/wqChELberDe7S9kq
2Bh0Zz3FO1g+BO+qBUVgKZryS7vt9dSGqVUF6uaNKBQ1XUg2f35nnmRjnBQIdOV2
k9p8u00uDP03aPOFi1HEWdhSaVgkH+ieBerPTItXBE2aE1irJw2U+03MdsvFHEm9
/aU7sxwTH5oGHejxBDNUFWOVf5gZUao5mVQEw/1zxGPlNJWbwHW2hCCrNTatsY3M
f2wNgkTSpIdv1NAHrFCIhtUp/Vhm4hhTdPWA9WEuNq2UbC+/Rhb7sVO1Bq4KTzrX
En9rRGCePFHmtBCaXbd8w3AzcIgOLnQLdROmZaQmglfjjktWrB3t/tWCC+vdMTij
5pVxnx2ROymMaef/ln+WXcl+NzxnmeJbYXP3tAj00q4gGUh4J8xx+FhNwvvdZ5SH
kDNqI1p8jjkUu/XhI4s60K3AOc0nn0Y4YyX6UUfVuzeI1ho5q4p3WV4SsEjq2g+H
vqFFi9XsxdH8ScdKMnEuXdqx6VLFWiqQ1l3Fc6b8prh1FFDH2pK8xJyJc016yE9d
8n9y8eP6r8SQoruLbaNBTdr3P+R7Kgyi4OQPd6YC7EntiLue2lA+tStRTwVcoIeL
O2aI1Xn31ajb/jnOu2cy5AZJ2E8XFXsC+ST06Q2RmNfnuD3te0xOS6KwpfwM8qRE
NFzPMe6w9cZVzI1Vs/dus/yUPuMC62zU2wCPOFny7fmojR5Bx6jaOpOrNUmfFR28
mVB/QFpQv18K6ioPP+LC54+GZgl/uP5+yyGWlWa7G6vDErIyTmIsaXsUOZtQyXFY
SPgUB37QkmYBFzlA7F3s7AFQq4dRqufHnMaEw4btb/0JfqG7AagXp5q3qolkOS45
tLmRrjR6XgQxc7EWEHpSPv+trAWd2dCjWh6Nux6F1sOKQKqd+QiFg9BgsPjcls90
vqpepNrIq9rtY/y1d0q+kScKCgYCZ+GvMWzCOGbmFZ27/BrOrsTFaZ52pwjJHtga
M5ETKmSFV17KwfSrKrVON91mCgzw9wMEtHd/+KH1ni8tm5/hue6LYWHksW9Zrqqv
ZRxUAulI8n8KjcOPQzc+jkB8jvb/tQ2yZnbRufSrfuJ74DwzHBdLOP9tzyyVCh7h
ZMOEtqMQubhVRImgNaiY8dx9CSA72bKVVlvLblIWj+jMRjzIcVlm3QP1NO8XShxi
1Akmy7U5Gr56Qs1GU++3wL3LkIn2tmbVfo5w+NPg1vNt76d2VeDo6gsyV4ICs6vc
GHxHiD90kkDwmhJ5h+nHmNNZX7+FOlMsQO1IctiYvVkT6e4p2RkAbBxyCrMbiL09
KDDuo2Uh3hf0NDcDu9UDXsFbk7OojMBjFuXlfk/yHd4VAlLKgfy0GIymmJ+c17AS
5BjB8LyVvthcsY5/wB8ZRXXfgspKqzuaPY/AJqHnqz5S5ht5ujW7VF+kQVhvLqAh
MPR+muTGY1DuIQqQkpi5+jnH6MYxaJdZQuhM24NIX5KkHRkPkl5ZMHOgXdLjT8Ob
8lPZKYpNS+Jo2t6X4ucDgQJMhD5DbS6OiA96ehktUK5l3qZCnAtRaXGkB3dkbHKs
HDWHSX5dXOXhbeHqSnjFP/s+PR15fMRD9DLkxVzwhhV7IGADpdo9mv/fP6EDnl1E
EOzJCUra9PbLTuF3ZywFdTHeDJ4jGuQySQphxwP3B3h/HnZRJNhSIFEJEf8+7aNC
X/hMEyrt2RKelzdQ5aRiaW8jKrj2UW1z+PXPV9qH6oagCNbsu3pqM9zNJSuMn4U9
NEmg6lPuxUdw9BLYOnvuyJdjmcEALb5wTvFHxfm9exjUxd1v0vNKeGZ+gjV2AumG
9hkTm4WSncUt2y/z0LImDbtQGXhNMxwTN/8ARoOd3QUWX2dllCOUFKeELAlG2dG+
d9XfH5A/x3TmLLvrcC4CFErArYMadWVJZSxxV1LOs4CCdrFhTqWwbsI5JmDS0R2d
qFjdqnEEYpaOjzGlckRmaMwPk204IUkxcmYkEK2ezGoPDfES8jUrbHar58UiQdtL
lvMCBQagmrkplhokGMWh0m2gWiCYxpzUo3Ae40vEHH5q8FGmPRvmXFWHDSWNg1cz
qFHk9a8E8TsxdXMgtdQA0lBkdFUexpOqCOhWy86yLYqNYrlLoKk02P9lI3q6dluc
pHfa6lukQ1N3z1O+kOnv/mzuUDEIRtj8P/ey9nOvukMAF4h6AWAgmZ2hqAHADW4R
6ZDLB+zOtkacA2qCV3LzG5kLiTd8OAv6XBSG5qz4MB1yat6jcnjJUG5zpIU7GE3F
CFQgnyxGAK2BtAHl5bidVnSlAVjpNZhkcxrKlbM1lpNR83TBF0BU2e6bgff+rxJW
Gr47CH9FgAg5DIwCvCJV1JP5PoBTI/O+PWu43oearwD+q155RFnIt6FoYieEagt0
wx4PlyME+NU6ZvfVCwFVEm3CB/Rg29dHKxtEXoGhpuzrfIi/MU3QJVFGXV1Xxtb/
hU26EpXOUnU2Ao3nTqQ5nRQIjmLDSXqJtoxKW+/ZCABdkYjGRrYpL+w3s5d4ZJOQ
mz7eJ4JeckWCW0px2Z11EvWsQSOYWtwuwcCXBb5ToXOPkrW9Yg3ApLcJBCcs4UaF
DMSMGUP4gc8JurA33bMep5Xh15moXTBn5NOlA+OC4TEkTjIUHDu+y2qQBFCVx04k
LnNHIf6AxgIXA6Cw5fXsYxj1FkoQIoqghK0qZDUnqmQK15fcJ38j/ka1wTblpMdK
MoY6ZiSqBkS0dPl1FaLoT65jPNZ4/kEisGld3/FqWNwRx+6yqdQ/FaXEJtArWatO
97au+oGBIcHqmKg0eoQai6RNsST43I+tpA6BkltQtnzXzrYJKEAurWSBjfKhWlSK
j6PgTI2kCQDV+BO13wgBGIaWEpncDXjpJnrwcW2Y1bzQrNmHGw/AA6Trg9EFiVMM
frLj9Kki4oEO7ynY3aWrFpsz+owk4BOrWjMqzaXgXI+6r6Q30nQvAPhegcpyEYVu
gWeyuzuVZ14w2MDE4RyvyRO+r01Iw6qFy+ONkujEuwUzjyTOgNsTijYGf6dsXXOJ
MF8TBl676nizmAIfYTOE+hnSXOCjXxKpDaaJQUiUFJIR4SuR7xPZyWWmapaGuqfY
/FqR6rIvDx59GLQj8GB+ZufGK6abgPprcZYzrGCZjHBa4cTJiidHUTNypyLUPbDs
pcKLbmcS4JdLWXJv3PPkoX8MznCw4OCJ55suzYMQVWO/lJ4CtwupMEDlmPGw3aer
tnUxL8BU+Qlq01hZy6j8J8i9SMn8LZPI6eoqnLP9DK++nWgjl6QDidcKaa3B7Sy2
KhNKLSpnUCKCHkZnpt7aQS7gjh4BZMMQ7Dtf2jWbHkNy2AcNpY2ergv4QVaOrBAY
TuMuZAGmHVCWntzaLSHnM6+bC5JUUu2XDqoeJniLkA7zRPxBVMTWqlQt0lDlAgXp
ww8iM7iTGnNFq6JI6PT/Tc5YBITrBOjaDIR+TfKcvtojLPw34h3RG01eW2VaWPDC
AkGHy0OTi41WoGwiDk1uA2QqX2CTHwpS7OcNJhp0XBwKw4vzlkZKsw9ML6iVFEWE
kPhc0sJYVkvCCnJluMXyA2yoP1GLiAEKl4uRY0T/batrLW7kGNuaCpZCO1z/x2rD
noXcIyUTk5MQP4H25prdzbM6/CADrNRlj/Jp/FDJSLcph/XuwF23GHOiKviAAVyZ
25uALrsAQalTii5C9zGhJLp68Z8v9qa057tAPGv2Gh/WdKTk44L2ItwGj5Cra5Du
XxP1qqyVsiRFsRJVrl5cLP8xe9YDLHVryF3oZcCr+KRFehNi9PEUHCqRhb+OJ2xV
knfg5h3oLw42dXDF4grHtlV7BoP4xIab+K8T0qUfz0ACpmvoE8WiVzGDPKxOPxjb
INux2GpJcIt0Mf/fOkssyYj7cTCdXVT/vNQ8h+9vkmTIfe5bvw2+t/aARVrYFYpS
zKAJfAWMarcflyMy6u5UUeOGXCP/+eyhwnjtk1I8cld8PFiDeQCpRnEKPCZnIL4t
QMDlWdLcc1khsDjjgoWhwy8bF46kDugeLou/Z2OTxJBbRTzLvv2O6g9/smyZSSW0
rSHdkdvFj3OjCGlss2o305iL/NYkJkCIV/P/Z9ZZkhAbXzgGISitaIvmikmIvpbF
t2o8sQizXUzOEZLImKLQN8zChMnVcfjXumkoCAgoYrUj1e4LzZQObqPmI/c0CwKS
c+Ya/MzFsgi6pGa0Uie0kM3GEW4PbgRJba2ZosHh+MO/jrLxI4ECdpOcwCxZZkv5
rpiB3EqnFHbWNxtgJd+B2Hwv2eUSCBBMujnygmB8rkMqNnQvxmEwkxqk3O01jEJn
rqybswkC9VdSuM+JC/8eojEPyslyhhLfLxmlB5E0YcBJIs6Yi0Fvohjfcuw48KMf
KQ4+uvozAHEyQG3t7Xz/1vivLkmw+TBTF8GomVzihcf0c6d/eHUaNzdYpOGmDyG2
iWlSrs0iiVmm7/HS1yTA5PlVYigg+UnnpuqML24zvXNtxp4YlytFSWaRgxaDIY0h
pIQT1+JvmbwWgy+GC925xyx4L9EcCqhQWaR8s9aejRrwOWWASbaaXjVOQLkbMNaw
jo6obx2mxPtOQGh5spOBmxVTgvbgRGFOUaGcKTAivW+XZJu0H67g4NNNS4b0cNOc
AlFQfUu5AfZd3pH7L67xNcossNmpTTKtbDNWg28CBsxFHZtx3CfOAtd2g86VUEVk
NxnYq7QJzZq3+MDbmKoU+nd/z6SkaFPTB+uYY9nC+R2EclZ6OOu138EMszw1IsoC
7TXr0/tYDT+1kAwBgZjTq9nRhV7YsaeBYIyGgtFH84eGjrFkqPeLAeOOawdA06OF
TZECi3ehYZFsVT5bhpi6Tfg3xkOHPZ2stMF0Es8l5w11LHBGhkqRC8sZkft7M0Bs
5814OZc8WeGMdly1kU+RqQHNfxdfg9VilmDk8U97lw2xybulvmdZKnuuU+FWf5QZ
0mjqR6TZlIDZyDi0/u+sTEKEhdDXg/DJyaWDkxQR8hEAxAUfOGVcFa1MoNb6qEhM
UgCGe6T5Os2IBZuIo8NjYToeJyXGvsB0eqZiZpgqNhBoBX8gJDuRWWWJF2H0MPNc
Bwejf6RXbdiUttreghMD/o0ZwONk+kpvXIjcBIsKUsGlY1uP24z310i2Cj6u1mOk
1bNtEurBPk9jvQ6LF09uC0fjKq0AsnZQsy/JXdFJUluReDTKh3K0Mg3Boh5SjC0G
uXOmWCUAlSi4GC3ywKY8X/jL4r//eLqoTYM5KOxhs452taPh82Sf9sx6rGX1OSSn
TK8WqjKlGCai/hUvyj0Fge2zFNtuRjRKUzjrH238Hi4c70G/5iCmfnJJRhpesx8i
f2/qgLc+czOj58X0I5FWn47VHQDwE+rNfiQaEaTbsX4JcQZippHx5jvRczFRlFB0
7hI5rvAL0gyz5xNXd8eK4X6CbBfRcWoNluAPIgr9Jd8KFdF6HeFu/5c22CW1RY8F
WHglcEKCdTVER6VEeYZv3KVatxbw6yQdqD9Wr/J+ALjShCiPOKnplVd2IBBhNhhy
zQObWr9GgA1N1e1EGhmmeMbcut1CkRxfnMl+eqAV5Wd1AEmxtUV+BsF7wcg2jhOP
e6jUId0hyOrpQgsIrbgiUN58/yK90Khqhw6ajchwhvKJ4ND/VGTYm0QwC/xSsmHe
9+rMk3Rlhm8Ry/KORExTNY3CTfq1s84kkrOh+Y8KeCd5SwbuM1RpbK6ZDmZoOrIE
f6vMFe5cR0U0O1WyTtm/DhO2or8NYGo3wsia2YeyI13boRWT+C3HccM4x8A8kh1B
WbcFK+XFDNeqnU5hP1/u9OFc4sr5VEAM390yOVxG6QG+XrbO0HeOmCqzwsR0i5jt
DunawTNjrWaSEwt0GsU+K41umd7fRdKzKUwLbeKIJ7l9XOSbkaAXDxDSXDYN81kY
ne0nRp36Btcs5GaTLYSz/u0sZYr2VRAKQdTrA4YnI0DPGcp95T6yxPf7tyX1+n4C
If4vgXvS0H/Pexg7wG6G4YXodA57Tv4vOtdBR0VXxg/b+dzLFsLZmSxbA2dIFS5B
WDU7IL+yfatBEzjUvnLAURXstQ3d56O3NSTNHc8Tq9H+JVVtjthrP7gw/aVG0iC0
HK5/3edoSM2IfSCcC9uyibY1Hoql+Ft4ZvJucVQqgcjT1TAjTQxSHUOM1kaBZmf2
YmV0quqRARiW9UWpZ0kSsZTIDAHmgk1xaI6q2qyYWm+5nW13HiHF5C7MIwKV1KzV
hPqKQt26N8f7ZfhDni9wg+9j3XhdKqmV7FuAlbXi/LJQS4G+vTv8pHU4mXi0Peiw
B+ocrGAJwUeR2plEA0NUJUNiP4e9BjwUcZ4G+vIYRNzUhPmr34+9JBzjUi9eR44v
zFoUiFoodbV+7ho0hS4Ls8NKX+9Dr7rvz7bHeiLQrnC73GKmOq2IsdxpemjWBv/7
PxEQnrH1QX7CWoRujh1ANo01TUz+aXdmaaR1Pl7c62PIyikS3tABgcqLOojHrd2i
KYqsnqS6hUbaypgILc3swy3FBcvYZqtG6LsIEZ8X69RjIKO2wm6oNHkVnzZMhyTs
Nrhiw8/L5MvKVMdzwdPH2TQTF9+SaFFzPbTBQ/o3U1IMx4RxEvU6luRIyWu3UI/K
LRwGXqKgYfxWvhnzsdmydu20fcYZEAr35OmmH96bAwISVLiqD8ktNd1IwuymIYt1
RBp05zp/W6m8ZL794UV6peKlHY9aVoVrSSj5l3UP0KszMDO6TjFwW/MDbohzxw1d
/QcvRPdj0vqjnNwdg5HPqO0o7HcvkZ9IZ1DtFOxkKP27Uqny79Xn5cGCaait2u4S
EzUjZgtEAP7vy+BI0Tn9sEW5b4/pN7n2ayuEmE02OPL87s5OCWbFTOFnDtiOotpM
PuybaBfsRpTqSnxuDRay2HGd4Il3DBSIVMdBFlYVUT8HWayKXzQu9R46MKhjvjBB
X/tW9WXWqlU0VuKg5kPwhThdv4xbTsGx89P/6WBxQ+sZMVERIfz13hL3BvfMvfHW
xEqRKF+RPpNvyUxSHgjcCh68eVP7+ScEsHOw6YKyoocuhrpMDtp2qDULffkv5flD
0up36kGNBLt1SkITcYo1/K9nSF7vdFs44lW5KVIP4wztazhVFrUEQtfDGoFyjrZw
wf8lFUMWZFRgc9HwIVrE+5BOZ4CHx3dJ+9Au0CuggQJUMFNno+uBMq139a62kEr2
1+GurEdHR/ezzo6UYHq80OoB+OjefvmapB6ifBWjjMFtqKJLD9Xvi6WEk2juxRbf
OGk50Z6C2zxLOiK7ZgrzqIS4J3UIJmLm6nKGnWtc31fUF/3NqWXGnkLzOxh+5Oqo
UnaAEzSyNv9+A18TmfxVE8J7VDfKaQrJiGbuIQmSzvEHCbJmb/XvvAf8sNubu7XP
4bxW2lF0qLrg3pPiw6Q+H2HZVyXO8lsnLFoxciBhMYN+J0aRXYFOOEH1vOPFOwhd
95TmNBlQZx9icHmL9Wf6ffS8rDyVFQGcRrmKXUiPyghZqmFsiuQmU79wFEWOagMb
KyCBJnPbRM6EvdpuP2y0epIfP1e7xcJdOT4b8p6/3oMzjzYXmv8yRV6UE0lVuwIp
R0ZwrIQlSvqlXA1aWPjsVYPYRRS3zgeuQxnkibch1TJY8jqXHW4+SL4B4N3FeMfd
DEoU+comjbWUjAYakdQJscfMA573kOAfSLeJhYNiPmPTveHAePO6Tz/gCENCHia2
JMmK0a1YNM8Ss62BC0a/sFTqAQ+ZJExpoDHfXfSlADwlP6c2wuDSz1tPofgBvr5p
3LKrUi5WKMmUeJItsJvRNlWRONs6y0pccIINP9Q2SQDKIv3YZPwDc7SGoU8UGqY7
bPtrphtc5rU9ca8j3Up5s6UPuTLpbyHLb+5tVjG57deBTpw3MfNHlSQbmn+OFY77
MjnZvoZHIMVy+amv7/c7u/fjMhCX2b1UShaj2Br3rO/9ttCPcUr92/GsqCKwjn+e
+P+rabIWP4cKz4XuGGH6Pe57AGRSS5rA7CS9bzuVHhZsEfaNj5o11lUJkZ+AiWJi
kHuHZm9I+LS1IiVrPrlM+30xG/XhtgVKmLHPFl2IOZWl4xW4iH61MDcnlwti4B4B
2MBPUnU5sJzskfPbg4Gkh4F1g4GI+Xi9VDNWyu3gNzUNaHtXMVXybK4312bpC1k1
vmeMsgWukm8eRcG42DCspYAyQSLOszFKS+ACp0A9LQtSr1Jogt8YYi8q7DYjf1Rm
1kqaG4Zww1tl/4QX2qk2WCwhI8c8hACqDjEc62AQs1sTyHLVZ2RAjHNFtlOkIUDC
d6JZdZUVGldR/yeSQd/TqSg7bf0JgLBjjFv6DiiSe3FmvtM8iXNHykgjUausoMLU
MCbqBcVWq3Yc+xHeeYlnKPl1KcpkWv6W9eA4znoFwFFPLWG7MEhfQbITxgyQMYVS
sRfuFD71QO3NdyYzg8YS94D9pJxU+QvQM77oWJokpSvq3RmXneU9ltQ71b0NA4tH
ztfulf54MXDlSEFcEqU0u/apuIM0mPJZp451Ml2/N+ZIp4E6brF3Gp13h8agUt0a
IretYPRSByUly9Hc2eyZKbIAgaIg5dgibCbISonCZah4skSXKabeGIg4SNRZyMCv
sZujfhpt6NZmNnNfyJRxkJiPqq3TnQq9JbvWXMKJPRj25noShGD266dyJgbtBhyg
Reapr3fmspvS1kMWVClfv2rnXjl3X6/CadGjbObYMEfOh/4eohOQPKJ7xtNTjSLk
XQ9mNK2GjNmoqpTTOp87RFMRfVqEBF/4vC6XYZHHI+xpONt6nYN3iwz8odl8w4Yb
bzLeM0kf48BNqFRNj6PeUAFIiGfhLDdjXktra8XtO+yke5++0b3+UlGROE/dZ4U0
+XQT1i19Djl4+8bu/lub4XwA3AM53lC7eCJQnFJmOT0x/7glqk9aW0kJEqsooXGH
rmXpHJH89UVDs9syCIYPkBMRnpsSUPowzBPznqVFojdJjbKLWdYJHgUdzOqBpqhG
9oC18nMxH2U51pJeiKH8ZvvYJFg4wGlsAxIIBqilk7r9HND6kBG7bsU4LKc4VdE8
nnFAGBdpux4LAP/eQG0jSMbrpAjU/weQLtk+36CBy0z/pXMhHPrASTu6RjjWy6mH
EXY11NLAlSmxbhRXyUaxTmIHqv+ooe+y8Tlndxajp5owHeYBVsaTYSyng8FWmG2l
MNCHJ7D2jwyNsn1hSJ8+nA5QGlzpgWu0fa+y2qvskoF8kjOoEpe/cCh0aVGJYkay
sVoiShJSWTPQRTUPNijqOALPv6lx/tzVpqZmO6NsASQJHzlzmT0qVGJoN1IgPJYV
qadTzMO9JLDlSd6L164Lq6NMo2Hnpqem4t5+ozmZYAJPfUimvxpyzDXl8F2WtYJg
WI0Jm+qEcGaxGVWetGVYcPmg57ZzJp6PuydFg6CASfZbebQ/Oes6Xq7vjKLw+bhI
NojLc8qmX+u4o0RKESAAd1Vnhf2Ys8So/r1em5lSDhftKHOonSNsR9U0rzma68Ub
wxV8NW/7Xw+3y9+RPJKjoTh9WPfDsQSh+G5QIWQIL8dC6fzh9AvL+zj3X/wFnrkC
S1ICQDvcGWZCoGQcknxYc2Bujp+ew4E3zZR/nzycqSnd/gICeH5FSKTw7ShGeim4
VqaHFNY8Yz/mv+WRQyZOdvzt2QjcxqyMHRSwXk04iLNKLaVQEuuqbxVNxOFXEtG+
JyVqsYFD9EDGXJU/4D/encPgpoLu1JerZ+HR+AIYLaYqRZnTVii54DDfhQ1uotil
HhXRz/jr2n0bKl950Jxkds3T5SDBVjqOzWPm18Bzdj03+wkAqiLw9n4sTIdd5wU3
vXDOLIygRXw3EryixJGt4ikVUvqEnvHE6YWDsILRhIXQwtvFDbbK7adLJotGdr4Z
ZObCDIWgqe5AXt9/VRkvKB3i9kmsJavreBZU4zBe3F5es3hdQNEAUPjou4fGpcAN
hG9CTAMLS+fpfqWd/fDEcqYxIC36DvHLRKgjATNMEHGC3kZycEtExsuV09SMSI3o
IAM9sjXwLIlIf7iabG6Y7KhdKhO9f26nTVeTWah1RY3bo6VN5FyuJycNNZEMA3/3
nWuj4+PDDudPCiFRsWsc/Tz/Lsc8FYv0ncwNuTW2om+SZLUpPdB5JukM8pZBkkea
sbipfbtxhHAQh5RhQTHZdHwfmIYooXpuUDASG704dC3FwyLgfN+5zWG3EE7YX6j4
YmqBjYCtzbG+Lc/vibHLI1nBQJW3Nd8M4JbX+A0/fbuj8zUn+GYftOGnWLXW/Ax8
wyiNhksI4fkkvP5OJdAU1mTzGnjna5o4FmqahJh6OzcoXr1cesvNbvOUMdeVlEKk
iRXDoH58cRu5Qd8CmEufRi9CqnuHWy8r5vnI+EnjyLqUe13LRPSc3CwFpP7wlFZ+
7sStw0aBtUvqr5OARtLt3PEF2mswbKhB4dMvAKIOAC1Qj9mibQ4JEbOWzCWxF8et
D5W77anRscm+JKJecgkDO7wainNaOqYXVjeiukukpdG8SB1d6+MOPGs5jSIeKaI5
W/qTQoUaejefqCILboxroDLbqwhKLiVXhGWL62tY6Dmf7YBfBUh5SQwQJCGLPWzt
8Y1xI2aJSEapYHyXF2A2mM87YckkQeLHvLG3TXdFa4kmnecRSTAhQUT5n/uZAENA
6uDcTbcxBChlrzqSVzPj5trqQsSpTllBMkBzc1QqNC+9EXqzHJ1r57k0kvfUYbw2
jCN8/H8AcQw1SyQrpPa7m+WSVThBpl3vjSatHRSK1ZDrvamkzAd4SABvyvYs5kVT
+Fb3JMxx1odjCxwQHjpupTq5SIfwOjrRNPeASvMx+l0c9T9SCbEdu9cNjw42BzLy
a9sH5yLrO+TAHHfWt0WxL500REhpaR3lYzw6ay/g5yf5WJW6BJVwMfGWowR51QSq
Fp0aJgsF1PKE8u9jpOLG8RWio5NOKlar4jGqA+PCy9jCaZebgVKt1By+cx8yPYQ4
hTAAOizCfj5M5hpjOIjlR7K8QKGDm8Am1/sHkBs4Xny/8PiogLlVhmaYHn4cOzxi
EZHcFqpXiKCDUsSKVdpCKObLlNypm8/sJFN5L1AKm+EV3Hr5R6qrU8a9HIPIly0v
PyDDcaICLXe3EGxFLgauaYkrryWzfZ78q1hI3OpAm6aClniHnlHkcPfCtVok3MnY
WwMg2fIOSFo0R8jXmKbF3LupzbinffN1M8QMvgmnLiS6lOnBexpkLQa+EiKoyPpl
4m5E4nv6fzpGzLEQIen4xXo6k/2LhwCVPHO/Ol6V6Z1u58lY0YGSfCuX8bJ2uzLe
IcXjQB8A4gxCjEAffORT10Ott6mrPr0n5/GOhCYKuuIBXc27lVPioXEwBjshhRcL
Wb775MbMZH8GTvVAgxmX8Y7OfwBa8/7gSmTYpot/V9A/0f1k6NXLgGHO07yBAv69
5Lu3QC15M+9M3aeaDGZBf9TsPKO0FT7LCLAhF+8wezViQHbzTr9zyr0zctq5Fp3o
trz04Gjyhpk1SydDCi59uY7U/FMMZas59WMnLrOgipejLlgxjw3KNHB9SLG4WG41
WkjmtESlQq9qSVyNEnsoSh6fEsP3UpYPS5yCbje/R+xdtvxj1EsGtJQSf7gnBfJl
/cmG+dSoCRooHI6K/LXcTVASzYONkPFMcAaXecwIK8CUnpchT0G4AT3PVBvAOBp1
QsIgMMzNkoeIYNktP2VeZK1bs8rM5KnBH7KOXypt1vl9ujzQXZ+KuCCNefZUlyhg
5hnI+Rwg6mTPkcim3Nyh7BwLqGmQEH76//X6R7DYBYJiVfC5Ju+8o+obPAi7ikvR
u95jwo6wvlshnKEUbnvyVyToQOB6YbAkxXvUKhoPZm8yeI+LiyT1QH8fr8XXVLyy
5I4KU3S1wMr3sK5AcBeyEa9RPZGYZAHQf/PPQ//GGGU9ZBf6SMdxq6U14lcpSp3u
9ZR0/yA3YxkyqWqZBMK9m2M827OsvX3eu6Lc+O66gH3BPK64+hYsMckc20p54M+B
z0B9DQ/UTitKg21TA6Aun/rGR1xo0QznYqA+rd4SW/2LrywJ5lNGQdCZViEV8Ezt
JQyklwX2gplGyAFZmZvnNOXT7+vYPenntGOZH7AUu+SlJb3eElTqRYavmG/I3QDR
B1YhJnlNPdPu4BMwtmNnBpJX11t4oH+UB0M6TQsZUD9a6Mxn4LkoUMgDCqbSFhHc
9orHgjeUEP1pf41nB/YV67GSHkyCwBkOzq8F/2987WniAHMSe2dFiSAbK/VpY0F5
mztCzTKsoQQ8hsRLuxBvJCOtRlQUYH4DbRLqSFV4TBUx1oLyWSVjXPWSyAqhky3a
LdPBmqMUv0j58gXew88vIvZvfjDYpbO64Y0Z07v0v4tTRR8+ZeVruYSysmRgNz1e
PNDlDyqev8SO+XamRUmx7WKlPUBInTk3aNZiqmz+bazA3Cn4wMWBRayKbmikHSzK
xWA+/CCaJMHLzBvxFmNduO9rorOAyEYZpdBfwM1fDq92uddfuVLOXiWMSE7d6C5J
t0GCesLPj8NTg74GkHfQhw/koZkM/ouZKj19f91g/dZsZ/Hc+gvI/5HFQBfaeWMR
B1/bQStOuVw0Fo+hJpQ3AKsw6ITUDqScNDby/AwsDiYdigQliXUD8dXl0BprM5BF
8yGgxNhbcS4usqU/1oSp3cEIK/22ESZxd+5S8dRmJlDvjibCrHiRDtRhGdtEaVXW
M3jmdspfISvfiFFbRzpDhEG+OnWQvfovMu1NfzQpXjyBa1U5J0bs0oI+SbqkDelV
EDIOr5skSIMgRs5Q+wxtlTzgIZnoSvG/CeqItgFv14FJ2R3tr/KSvIWexC1Nz3Co
n3qIbxLQoaV71ofLlejzZ5ceRTmm2iLH0Cz6fEQAgwf6pDmswVl3lRKJ6n4Z1zst
I/uxWVMzM79qelomHeRajpLC+L8JgRmlaD8uI7RuJfw9uIe2AWywfejnD9CaMyTo
i50SiZrY6sdp1VVph0EbPKJN/QrWGzbcbzUtI9eWBzhokOktIv+byh/VcpjVmOHd
+ZwL8gu2U28ZopZ2/KB0+WixYY4YDrRM0twmSrbcKwBGxD5EndtIkZDQNUjt6ikx
JQuBxa+mXfJinE+Ut3n9Nj8vWuemhHOuKiAjTYkVDWdgaS/aa2NxMm98BTzMSpQa
zGg/Oelq7/E5TSobByqAjSoOpbDug6efwODLKyy8YZyfvYGAYvtaWMJjAkhylf6T
f2sIrNKcVWWdhQgLIGPW21ao0oR2UZvlNH86ewfXR4m9h8jxgdrsfc+x9avoNGxs
b4GZNr2iIjzoa5bD75s05aRk0WEE7irzHuyrOZlGIqVWR7D+XSS0BUMcAY2/XpT7
rrQXgnrhFqKjHnIYhXrtn6Ncc9TpcrAqs7yxJlczsaxhaOTVRdLVMFnfASCUhk+i
4W13dQHpolLK/mSpebg1l+zNm96WgeOMOniWn/udHny4rFMMHOrJnoKSxyGn+NhA
rX/skU99DP1zI8whhj3RqoW/Lk6j6RqZUJcB6PmcC9Q9eK5x+BQjo2vjIJXqCgTy
Kp/aXyT6IvKzyXuQjX+eZjd0EwdllWTPjOurbYOhtKZGQVciit/asoI4CsjM1KBv
EM6hSYKR+Z3JOcf2Vt09I4khOL+9Jhp6uCx86Ar7FAJztkYgmjZuF83HnMKTgvLp
bT5gm9t3ZKutoa3Imakgfq9DoPJUrDKBh1D8UGqmkESHP07AyUsqC33L/TsMzU4A
icWJkfJfVEtlmx5yX/1KMWfimBjuzA4OUfGT5kUZD4t07wrZKS5hpF1S4oveNqAc
2flj3P2dhZpJrDnWjOQLgMx7DPNGc6Rq6rUiQ0GHEdfa3gHHN/ujSKT3Oq0VlPgG
iMUgz0/Lwnzm0dp/yD+MjCfOKy54HhgKZxtrVh4aZB4jtTtDm/0ORT49BKmVfJye
qfwoV/mCT4mxpV7SfIHvxY9nr4YpXQEPr6njZtkYxh6lht8exUOvCYj6esyT46Xj
i+hxiN0+FYaUsG9swD0Io0DVpk1FAPO6VaNgcCfzRyfmym/T0Ir7AG27nF7gvC+z
R3mS2ubh+TKkTaHSXH0iszxiuCDAH/szKzbZEljcstQRK/d2r6opq6LheYc09DYp
fPJCCUIi+2M+7EQZHHX31ePTpSjJbCnWC/bElwRCDJph4TcFq5w1YchAv9u/Qw95
B/omqF1j+QAeI+c4dOabgGk3zjaaBn84tpZKJNk5rR4aPo/jEeorrpbJPkIp41g/
/Wsgpz1+Yjgr/uFROzWVS8CM7yRiAysSuz9qk8w7pWTMjWxX2HMGKjVbcEv96cxL
qYhv6AyenxgQM+5SP9QfyeLAbx2vAoAvyO8vJPixJfH3CxilXqrVJRer8uuJpIae
qLsH/5VDMoGNPDbKoReInhgRnUYkGQsjUYKxt52vj308YF6utsh0DXlkV5u9pPzi
kx3ttt6sYuImy/bsQhQwCCr4lIfPGxxMEhr1dNZgkgcvq1CSBRgTlVmGjU4B7hqp
w5fcPTSMJGR30SUeJX6RYlNpp1r5+3RfCKeNk8pAf+3WHz3wJ5Jqsl3lEcz6qbTR
kQMQc1iWPlhmoQRWQA+JOLvXWwa4yp3cUgnMev6FoWqy8xDoOUgC/DI5FcBnf09Y
azC8juyvYGHIS+6VcVARZMKJom460dD+zvO6/DPuWloCKqVwC/0HgBbhPSiPQ7Dk
tpbj/twyEs0WPaRYx/4QhKBcJfiBeAmlaslP1HB3G7xVHzjantJ70wCGQqZfXqr5
VYzm/gsRm3WCTOesC/z8I5I8zCjzpSKlMIM0iKa8l5+AhPoP5dzf8AqXFq5tZ2eU
MPL2fKOaDfxKdXtelgL/d+qxh2yBzNx/92pwvtLGDu3edav5fiMwkAF58jjjyCsn
jzDKmCfo4tA6kjsNDaQtMuMDoisZ/3cs0xBQS7MpDaucLWbvHa9Ark8zj9t+Zf9v
1rqCc9Uxlryq7c4zuc55EdSZbTi0Ico1k5RoAdim5S40V/OzoawgRxgCxMHg9JWY
s2YSh72sxHdEbUUCddIQb/ZjVyVBi8KnD9Qy5ev1wCtxI1d3JK+orZtt7yz7Zoco
MOmypIphWNQANn+nPjsA3n7IuPf+Exo+QmFqdSyO1tahAVd5L1vLdsF9WvAgS5F2
bmdVefgTUhYsg2KVWLnsDlVa+ZqN9rhlFSRgizDWdTw/R46vI7lok/3yjIAVHSGk
zAlOBq2ffj5syZsNh8jyNIJZrHo7sgZVuZfhh4MzX7i2qfX4eD1vDOxvA9NTvfKp
wI76/PmTjqMMEUgEkvCc8Sm0YofL7XWTThF7yviDM69RR/B9hnF+AiWYiRgvrIKm
cFFDIqEaDED68yspUnYPxxjABUf7u6AfnDKQY8DzwM59NHpNeIrjGm+tOhxjt9CQ
b4zjpxb2olwUAGohcxmpqEcgDQTKy3hukdOi9tmzsa4ZvJtsJ5HM+SDYRrSZSwkF
Y2xQBur8pYcJakoQQbNioIRLDTYQ2l7lptrhrriy6+0pEgRCuaF4VwuX+UEfHexI
9NE7zC180OsIgEFj5u/TUkAR2/eI2Vr7HvToZDnO0TZA57ynwLsj2p8VhK/SCRbS
iJWSBGdwSvaaAn/NR1WcxRnYyPsqtiMX5IN4RCLHRgxWbhyOGqFKpYn402ltk30l
HZu4TfaxV5aUYabSjGxF6tnvAv3YAAQTfGY2IqAgnrle6SVTbHpjJEe3Pusf+rTm
+isnX7gTjRWkkOwLYEdmiZwLfFe4ZSiCEiatxYK21JLNaz4JxBIxmfj/HGSpe1Rl
GugmKB6bQPuqPDbTJwuq9lPetqMA0UcPpymdQcLzO+guX15l8MKm1rbhPkjx8rak
bT1Rk44d1LAG66bKA1TGRXqdiygWCiDhF179HtfuYNolxOWIXop3KMFMQOfxEUV9
U+GSJBE5ZzQtSqaaFLTntLo/iBbwevdm+GqGEedheB+AGv73IrK+gwz6z1mT5KSI
rWMvdokJAtBsuwmPRlb+xIR7MEvsTef2ASvDkeXXxOaAue0RbdOkdh4w+EmjKsoN
jO9Sm2FVg0+WSfewA/TNltpGIB1A7akU6foZrMm3DJC8hB7TcHkZPRLi/qta0o8F
iGkX7tC6gAwpukk2AGBao+tN/TdOddKvd9L7IoS3ZTValjf9VSY5aqQTyLiufPP3
6GyFfH6DvhmVRn9GEyRLTIXNEbakj1zN97B23wpfK80mnK/KcmRgm5ww/Zjfj3hG
uhGUifFVD1ZRiLlBmVmSJ98LuyeMd+lpa67TEyUaxppRvTMsO+yhOXXk/Oll0UPl
LRX3G4yzxyu4ynFjjmmfzvAwlhFC3gRW2S2r0z4myY67438ConzXeqHpPblrqOJq
+HWXgybszhotcOB0JVk54hnAkG5beMZZqA+aYf5zVF5jdN8ddAmoXrmUC/zsy/zL
eQ/12+q6/G02L9qeTuawe2wslYA+3J6txVxmHPTSrUsevbeUCrpVFGwWnuz+oIYp
B1itc8dWwC95Q4hDdh9ICwubFwaUEPj7rbCuCgWcBsVcPA/4aBBuOZCpFGwYCAPQ
MP0pDV1A+lyp7Gv9cJev2b9XmsfExvFgUsP/EgZ2i9swRL0Hw4eMzPYvPx4AeB1n
AYr6DQvKJftuimeoaWtLYsezajje9k/hFfz35HAvUx0fVxubnSq6d4YwDR046H2U
VTBheI7hQ7rLG6XiQeVHgTc3JnOiPkEncyUNnU7UQYUwygp3NinwFw/61udSE0jb
3tVWAPH/gRiPC8KcSXoPir3Di9ETD19suLG+WkaYMsIdsJKWZCdJtWCWUpCpSem6
yRZLj8e8ipUknWCM5Riao7nMtJ60/EpwbmM0dG1cJfMLb1cUIsgaMDOzZwamcEjn
8KFIFXXnqiIzfxzHcnRGy2ECwCJtaHeRp3jhSc1TeVZk3Me0G+zYH45t0kZZUy9p
GSaOTWrOTShsFNiIhrLBCUS61c2jovEGx5MbpLqxRKy58J2T87onh+ACMUtQTSYZ
7L3Pqo8VAXsBDQ+IMImpHYgGxaxpR2jxGnFsyCSlDuK9pY0yH+aHT+0sC3KmQz7A
XsZ2PheBefSd4gUAltG/LwxJ+75uo7uOpqkJZIiIw1e70y8pTOJ/1RGIcamVXsYE
Gc6ozw0U0R5f7VcnnErd6EQ92QHPG9ooAirun5FBc7ufFOI38SuwMfJqTnV3e93T
5El5QZtTBtR2vgCIym54+3Q5VlRPX0IlJlqP3SEHyDG5jrG16sYyKBZOACYBCfnn
moHGi3lOlhcprmMI5ybres0/8th+3PxN9TpCuQcSEughHzqtK0gMbf86NgMpu2Ej
/sc/U5rtaltRROv7hSCSSMkHTIKrNm/qhzZAzVK1hurZ7m0U1Ezv14FfQvIZN4GZ
gTW7QlWXRP+/3n2rnHY9kUM5ZjqSzquyTV0PZ4+iuatEMtNHyFUnEnvmIJgMPOKv
CgbkHGze16jbF8wI7406dNvLMsaQdd8d//SEtQeKXTxazYjal2APT65v2efWtpK1
aDJqphU4LFfXDCsQwo77KkkQSrXgaA8lMiC5Bk/AgJUQo41UWJiofTslbfKk+Tmy
cEvotcEyCyLeT0BD4v7GNWF5VHB1ktwMthIOZW31R0pJdWrjbvFoUfYu0QCl/LPD
ntrhGGWLjJF1NR+EtBFrQumQ5GTx1RKfQQ/MnwiC4ridTUHeEQ9mbvDK2DIH2GYN
7sP2hVXqE8Wn9kSVrrEef8dQoD6iIb9IE+oMlHmDsh2fDF5YfpUwJdhLDUS1SXeL
0+qsmhh/G2DMjy0Hv8RtkViKOm4qRlIEZBBRVaF6n0enqc1qcmSxyFlGmO+KPa0I
TEAIZXMpKYA70s3O5zPDAMu4py5cxFAijZt5NWDd+1LU3VerIlrFVIdSz47TxEEF
cic8wRo2Hze8TsYZ85GAnH8aQ53NPWZ60gB0PODnufMkvygVrTRK4I2qJ5piegjc
MkvB6TXzivuFfoQP+yyfIGXeSqAP3BlB+MBO31CTm2ytVXrjq86bMfHDfqCkXRKA
q66W5y+9jK/liPoAlQ8a/JvIjYv+JhjTXLGGkn5hGGfCzwgmAMR9eKq+E05M7qJD
gvDVUBbuNch+6Hd8uHawYYV2R8vzAB/p+BpfHQDav8oChzhcLmuH0Y9lHHIdzXne
3bjfZs/onmal27K+D40Jq1qpZYPccAgSyn8/TDzYXjg8rGDO/zFKku0MFvcu3PV7
g7ZvRAeivxb36qbnU1lCvOSdyLnHc1jS1tz3jq61X8jow1S/QCP8Ir0Y7A2rAech
8lh7dB7LDfes4cLQHbUG5DYCMtzUbrlg1wPfCxW4c4nyK2b0NEJdjN/IS0kn/j7H
Vf2sMi0LpQ5ZlPm0MkDRMT4drEhq14k/q1rFAIK7uVZd5VyQ6jPLATmtcSFU5y4g
xOSrJ0e6bQz/WVgP3sosXj1dNJNx1F/UXR56c3rQauiMsvIuzQJMUCHtce+qmi6p
etpIcmXbYPiVEbq17iX85gvs2HnDzusQkbQeWd3CHCOItO4KaYJuJA6zFdytHnfm
kg0v6YXj73Aek2kU0jnoH4YNeGZb2SQvvDNQb+d6p8YA3kAdfGh+G34INAioNXgk
IaXnLoTsIxtzyqEBr0OhXp5P8x+yN0D7Wk+QJNpl6VdDHlavM0desrkufxoUTtbt
SBpgFxSe2JNtWO0rNCLqJCDz3KEdHEdO6AW97tMDxFn7h2XexbtK9OmP42ft7YRw
w11Q4VXhT2tHKwA5pWQVkSJJlz3fM9fhuqb+I8ZkqGSavByFpP2HXUQyK4TcSDHQ
5UzPRH/D7i9ooNysIc9Y95VkqWUzQGKUxU9E0YUjfRpXIGykb9P881Ii32gpNy5J
/Z5IgeWjbbtxN+JGcRn2DHP4mir0MvchfJsZWijXv6OEI056f+HAjipR/we6z8p2
s3dN/gC19MyZvzmvDNZK/rSoBg/3L8+jrhF5sDZzNbRLHbmqWZ5RiLsKZK+NuMtX
AseUg26Rgko8SYbuQfQplyK5ciXCARGEEbZ6s5y5Y7DGWvTjN3Grgqv9w0kZt+bW
txg/eic/PjChZXfkc2Y4ynivfNu7ngXwki00WsnCBFWGzXIrr86zoQ3WlTo7jET4
5QgNCXuA022pSJ8uJruEE5uMio2+TpIzpZ6WE5jXMayaN1BNBnjEAszLBMGhDDt2
jTJJ33DjuxkVNrPmOShPbjqfjPuPkKcYm1OC/Kt+o+nZLwqx4mfZv/kurr6a7Pn2
ge1D7eM40GLDUobtKtMExQjydMLKAfLfKf4MNTgdd0jq4vo2Q0p09TJy3pdmU1hJ
8ErhvnUqJWLysD6rYWeMhXMNpZFmomXJTYhIteDhwho79QSL7/i+b4AJTZLYluLe
ayM4s06axEM0dn7BxwtmCqTR8AJlCcgc+167d3MfoEMkoyG8xCigYVWZ7mLkegqI
MLG/UF+4Do7H/jbPIdXrUmEAiOm+51pwfOacwzj1mb5O6bYorPylCAT0xu1tWteE
wbRfLwiCSiU9cEUVYTRVFcWUfZIfpPS0XGndwgWj2R3ezuIjuLOWx5M5xHX4w+Ai
5vi2wEQO1/qp1VuPmatRnrOuCEQ9E2D/moOkPrzMK0uplvAmuy3beGZxH26Yi99o
LP3zr57TDm/CXWPgkpxtLrrnAfXub54EB3F9h8DU5wbHZJYiEgcTpr2awJ/us6Mg
501rnyCVV1cnU2f8rlgCKo6e30WAzR/QhOQAinW8WuKTu49PvQTF+pCtyopp2gB6
Cw/SoZUS7O6dN6fDUOQCmLcJeHzDDq2fcY1Ccu8ge2onQpZeHOyAX+6Ak/1m0gyp
M+byi8F1nyWliT9yUM6gEkzKRvz9Ko+zR0OVftFncYIGPKlRYLggXV6mnUDxOKUz
KvfCURQMpWJlZaUKGHuxEJxN3CCMaW2HxttvzATHcMtNkszX5xOWeEjSYxJNNjJ0
sVGtZKUU2rjLzYQHx0H5j3lgNDfnLzaMJZXRukYcdLiqaRByUBeewjXFdCBq7WsP
VTMRzyk+aNW9PAS+oyuhCTKDcVKOVlY3rJkVZB9ePq0ihfm6Wg2NSqiFfSSJhURU
1BgGskklUrNzSclmTOb9d7fu28R38WF0rHMFNXnSe0BSTMUeY2O+tOOvwTicb609
xYVcHJlIadDyzTNsUs7Eo92rEX+74dzHP2LJcYx5iGqijrojHjH2gEHvS/5ZFQ7C
hVhih8AyzQ3/1P7N1BYJZhWdlaOXjqhDlctqggCvFfNCTkMyXGQ7mCpPSwouidvY
/VlXABN9kJzTvCU43Wp10Ccy038cCIlRTCT9UgNGgpookIbh0TjbnTof4gOo0psh
BkBr0o+k79Na2MiLqVyJoOMrrCzNfmvN/NTYCAXx3bDxLtyuqZVwhR/dMJk/X+d6
TN6mfEvuhhqv2AaGcKco0QU/01GlB4KfefWY2j2TdksjuP/ZJCvfVMFLjCnKgN9z
KvcMUch7CoaHHzJavb4Q6dTuMrXdO3pXEvLeZCf5QUFcVcrPobFgNGjUymA8sK9I
TonUKqohgYJCfC0vR9CWMUwmDRAAyGor4XzoDFGT64yBnpkxIHdvyAjhuSGmVqOM
Tv3Po4nPUuLw8KwBYsvlHf40YniioK+fqkJGHWbjqCbwDcfqQFig60HaD/pGZinb
npAyyCHvHxaqCkgljrBMUP9cIwE4+U8JsW0hoNb+z50iuSMp6ZM9jHxW+qAGIZRK
WtSknAufkdrpFImTaD0UMeMR/QJVAXVL7GaXOD97w1N785XCvAM6ybCyQPx8cNjN
bYSOaxjU9+nIVsujAM9wXk7wlBXAqOVZqstFwVNmWFHcMzaHH78pauqQ+PecAgZ2
uLcOMBGVLyq7N+1CJQEswPT7lNmRjDwLlhPLQropAB2h7KmdPddYcEeBzRjSSBZZ
YeMkJPovcZD+Z/b0ntyDi3uzJGcUG68J05+debRHWUodOPJ5JLKSB1YL+UyYHPkz
9w3ZKuw1rmhYzhcRaYGsi6YzrAcR8D91Y4iJFT56Q3mJDBnZrINrZco91Z5A+fpz
CH9IYvyQ5Lf2QGgrLfjz0fG8vZ4B4MK8USnBqGDMwjmOApwBAHT5fUupACqoOatl
zBLagHLjzoT7pfv5GSrnQV97NQmJg/+3PPi85tplLrLdr3wU6C/joKN8+pbQOEv+
IMmZLtgMU/bHbumJPFjLEGopnhbXbWqscGRb0gt9vsn989N1Ak4dnI5s4yxG7a+P
EGAkeOWukDEki1a1c/AEJc62X0vEcytZhsBse9lk2MM0NfQWFZzFOcOEcdWsVbn3
kRBsOBIeiNwr0WVqLJRqL50/Mjan/CpUImL6f7gf6vvictKvFFkDeQAX3GuG9rp4
qnjksx9Au5S0GlgJUnHJlIYpSPDlDE1pYYRb1OtXvyivyt2so5hqMhNyMohsF/Zs
voA3yFvy/DeB103E0p3qWWdT0BPOgSMjX9zBacrlT7elGB4kVT0herlijUcEkfZe
ANuhTvpjfVIIgBZiWgl1vgXeTSJg0cDzhNuIDLbKZLh4ckuFMYql7Q/NMOdWk6pf
yQesWgV8rSw3M8AUlhFJOswshwzGmxoshiubVt6z5AQGpAv6hw732VPTgsPI9uFJ
cqFozCFWuskZQSml/kLmI0BDTtTuJQNtCvsc1Sr9W8crZ2aSa26E4Wi1hUmNAyW4
to7d5L0Txm1hs+/jk4F9QQhuxpgh5loxjZhYGnbeJZn2S12A4RNaPI9rFeou0SL4
HZ3z+IPefdZFXxgf024e9w/QrzDCsO0FyjkT8CUt1gb/7eGwODJ/s8d0o6iOqhhq
Nco9e/Z97S/7TrpdhJ8ZlbKG384F49zPjauYhDolenZKrhCMdSscdQ108nVElDnr
Sov84d1WGTMwz01kkYMJnhId+Hyl/e3spPDBJ6+6G6Il36+EDJnWwzlkOZ77+/Lm
DWW6O6QgbJxUie/E9LONFw70cNsu/mXOjNAEGgvDRC1LqA83k/vkCqeScpyIhFyL
aKdxsnotLKBWF53z6vPDtWCKs7BjwMAbvLlKW+UknTD9tVVhDF4MPSuaP7cXVV/9
DtJH6Lrj4Fb/gd5CzMtXEeKHLT4AsFB0ohjfzYBjH41QZ4U2Y2XyrcGW6JMqiXzk
zXptuPn19Jr1RTuWQ64z9QKwCPCkZozoJLm9B0G13p324YqanlBj0X4FWNeJxfk8
ujb1SHCCtn09svroR0h6muIQQ29rANXPn0mXl3wJbtTy2VQtpYT03x2ETDddgoU7
n2fgQvnmf6uguQfYMRHbGYjXMB5S7L3Ua/Qt7JJwEzSjCOfAEeCkMQLO+lQpjl3n
ZZ3eVZtWzpXlUIerhr3MpZk6PI7AoePRbAO6/MItV5Rg1iEKWuCL3RW6TVWaVVGT
1cwM2qU4bMIVmopUch71otGqxN6TP0f9Ot/Ftmj1nfwOQlbtfPBQLc4ik5SEUPXM
dubxIvPdcmiU/tyTL4IK5Q14PDGkyEdDyRivPJc/0e8PcK9cBFUtcgS7pvC6Uojm
UCrKcy576pts8HqSJBm55XtFHANP8Kje8v43+dwE5VvmsHILzbtga4f+rFVo1G2B
0HT19HQMARlNVUHLRy8wjUxO/bzmB8JOLkH9B2FSGOEmWWiNDu98Sol35FA3ZdK1
+coqmKYRY/jacFLzuwbiyXqgmKf94eTjWbT3cWZOUc/z/n4NR5itQgwKyvi7Zwa8
7k/TABnmnTl47FSP9h35u189Q8VcQB/fww9IRlcECopwGVmUpHJYp5BHJPAfwM6g
vFSGJwYDmgXbDNjQTIR2Izl0l9/ALQ+xb/5SLv0nYFv8bQbEOviqpYxTD+t7sEaN
r+AgydAv+UrVuE+vHda4vRoijYQU0CZoaAaryaOFfgYpSQhjcsfZap32d95mTxmb
hDqnlaXSwbnwPaNVhvydcdDfAlDNSNBWehWjY6mJ1bPls/ATZV/gJWsTSilSwhz/
znZqqDnr3qxqxEULry5ecVQVoj5z9eR4xr9uFUcXREDE/4+vpZ09vnI2nNUH+PX/
EhZzHcSP9G/YyDt7Q8tmP+n5L0h4RI2IG1IYEMAX9Bh2RynDZ0M8RzMyhqOF+/1L
siTuvGJzRZwtWSC+fnsyO0+KtR9tEn5AwohshKqryBuLVK/nJqawxtn3TmfvDYGl
IrQZlUW2DbzPPpBdBSQJNv8XYKmhjJvBtG7Ss4xSDTQdXOFeCVXxIJL9HPB+FvsP
Hoq7550jG3MwEHfsi7LHP0Czd+0cTs9DNPr5+B5QwZ0t2YoyBS3qwjTikuRuCQju
Nm6CiKwlHPyJv41B2gMb8YzT5dx0MSt/WJ4yKMyOW91X2ulEnSG/N4IjtuaqVqET
54wCbs7o2ybCfaUS7n/iANRXPBrS9zpk5BFl9sdAHcEaSXFb0QSKmUwr8IoP/Ixo
+4pzlQJPTT0mCIap2gJC+9+YYimNzY8mXmPxbtVDOmdtZdul1XOBDVqkCwNSFPw/
puuI8vmq0FaUn8tdrSehR9rJRL0xOJbCIAr43am3oHrPbDQWQkoqrFO1hCXZHWtK
WdgpFV/fd+TgrBjgMUNfOd+zkVOhgoqMKi14YmRjU2XnYRRkICBGM8AX1s+wNf+D
ybS7V6O/sHSvIawky0FcKuEZ6vkYcoSn+d/wysmLxDx56VziSFWoc79Ur2E2xFaz
fDZVtbres9Ub9+0XoS3P8DKT5fjUDUooWYHFjQLC4yrGK/kn3+RYwLa2ZDXfToSP
BtDYejO9La965FKC/N34p7UqhRqWzFL0FMbz5wi9QH54ELWs3JOl4NqGFft8VBuf
4LRezYvjWoVVl0DnaAginD1O+tOXx1MtG5koAIck15QbghR9tah9X4pEqw7UslK+
LBxJhE3y1+kJRVMYzifPuPmuzbKIR5USfS4ngNHa0YaG4NKG74bjmwW5lomw9hQg
LCK8wfZfdvr4VEP/0PYbnQ81WO9wa3uP6AbINcf1H7qrOlaAcZoIAYzYJqGf4Qcc
PYhha7Amk/oa01Gczur8Iu8e9jINFUeFCTLaeNYqLXn2KvfZjF2AWMNfXgpqscyT
FBT/UbC0y9D4TIXhFeWmR5KuWDMR3xgzGZgsdgg/XuwybPkVpn550lNsFszXj+DM
+50T3i8h6sPzg/pwunokcVCSxPO1eU+4URW3J7+h0pwxZwOVK1qhgFVywLYTf4TG
aIhwjcZojCCOdgT4AI0/XpwSbhBSD+YzIVVDpg2OoaSerIsKY0QiMsbUQOYUKnso
GH9qJ1iEtuXjtnS52ZnZISB8gtzdUb8TVAsK5upJYGeNUgHzybTAcGZNXWsSWvVO
5CduSdXSwfUGpDgxn8agBIhdmdj1sGHSHErO3JAoTkNOVzrX1Xea4NJOsFpxPh7u
tzSJ7rPRJlhPIopsvgdBJUMJdJMrOkMzscye/lWGMu7YhzmitwsF772AiIvkXHf6
b6VIyY6v/xInYjXZyMGe4fSwmAVFQh/5PfC5vaz1U7uptRG83P88lqyarbCb1jOi
yxZFrPgPOupFTNjEHzANeHH1IJqswovpX5zktKWRxIFBrFO7w01u+Uh01TkInw9M
WB7GHwJ1/mAPr3cufLKhDt0Tts2/aQ9f0vivp7rrUVRSvc6VwFqjjD7JqYAi1eOP
1drMCJ1/0cmZntFzeWpjfTVGHCgyQcy6axS1bLIdg/W43YzaZy/SJ0K34qz/2Sw1
bc4UUu1ZisLqYUY+gIZJQnLQNSfYrtcFGbWrmFe5HbiD5h9YI+5ESQ8wWddX1i0h
sjNOZDYxw4mWfgaop9wk99SQVYGqHtndToUjEwbEEyOyl9Yw7dQPakL6HoT6lnb+
aDiYjRx6984rwFNVz/x+IzWPE7qSmxVYoG4AaJDPzeJ7h/JzFM3BJerwPl11DO4p
X13agTv8Un7WIVKQJu3Yf8MdSbeUP725WOx3Ji29ZT6rg3znB9Lv1f6KrD5Hx+Vn
4+TzUfi+n6VxQO0DV++kWIS0p0mAM06KNlplTRwuI+l4uqmyHaV4jwp2V8D7FwMd
u5dxovk72FfvgFMm4XX23/Nbb6Hbr0TBkKab79JQDr/3WtkwA/NiBZfjUn7R2vXt
e89HTEtxCxI3HORCs+qLv0zXKaIo4oBw3s4MVRN5lrJf/JR9PbUMV7vgCPgis87x
DufTxQgy5JHiMlxY/qazFK55/qnjjKqlbfcXkeuRYJ7qHGAr/ZiNrMuVexiepI6u
VgPd4ALkOK3d4xW1ZVXglYVCEZ3Cosx54TG5K5EPqvJ2xjtNgg05DXaWcBMYaQkm
Kt3T5oV0Y4xKEScQQqOYIOq+ia6Tmdq6nZgiaTIJAZQxGxSbat4RDLmpsUJs0E3m
s3jfV24OYEuAr+JFG620OtLunX/ltV5SkWjsSzp7/p54bhePahHNY5SnO+8uKeKu
mYeTjUMUvZ6d/YGlc60yFMmwziGTls/gHIsYvIMeWu+h1Pjby1xgOD0Y/bQVjuhN
bF0/7O2aSdYerIDmc6TNhGUjcZCHc7NlblE438Zaz55lz/p4LIQOG1d+fAk5MBkY
aZkz+cx8asqyJ1lC+oOn08WyzdJZXwVfABr7cSYXkPrOr38Gmtfe2/nCUBz1D0Eo
pfmViUKP/vroqFyh+HUVCMfZ0pY8h4XG/FHUcnBJy/6i44PX3WIW2NnT5I7B1jyc
OGXY9rFFAuQAF1iRfJSYB2rQMx0qfmPH8MKTUPo2pjBTNKWVj0eyEF8U2528elsW
DFvdy2cvfSLL8bc4tGREPo4laCmrN78YtCgu9iFLoy45bbCajcFf4cQQTLUxyd07
NmJmd0Qs9MLei+ue5vjbACvFRe55mmozNpM5nH8rGfO5ZElt027cjKxCf0SD6JF1
5bkV6S/2ZLDoCVgBwHuLN86PJYPF7lYFC7/hvpv7uloE3eahXRX6oNTkieDNS/v1
opak6zp7pY7ievKjFZSbXNfGj+oGaIRDfY3ePbDYBMmJqqDY3ZQ/ZiMDBuxYlreq
ShRhlcH7SYHYFkLC6NQXhImkv0fNmwGKj3BGdlBDc1j1BLV885IgpO1PzitHxrNo
viqmtITKQp98lltx7uCr6ed6XSNBcRNgl9xaiUlJ0aDikWrpALEdDYeLvIBpdf72
tnnLjSTMYGjGMNhYlR5dp2+cyqy6xzzZFMILcOy83va7twVbRTd/u9T535ESwqoN
rw8wQxxMUa9xWkVLfeUN3vQ4b5ksqnHHQEznI7ZZ4Jvz752Lq5GBNuXikPXD8A71
bjdavpto8gniotmgVyfqdL2qXlfRuZYRBEFSGIJzz5A0ESUJwEQ1oXkLDvB6RGqU
y3daAXvixT1BPJvvru0mnTDBhu9pJ4crOP3lZS9SgxcGfrbRt6YAs/rsDZ28zaOv
ZxPSVBZiVVSAJnxGNgA6jpU9/2rR8RcKzONWerVrhELZJyAO6e+qeeRII1pep41P
gzdQvm1Q/CngpEbNbo1DiE5rC4T5aUf3DVGJvrfFakNduyQMYHwgw1CXGemxUmFX
7Uoj7qdiAVzae8aswaWBHxW8r/f51YOmqBQPrOLAhihJmVqqiTr3pgyI7LC3b61/
gr51uGgSyND55VDds5trLDVU7iLjKN3Ms5MRchRtwSnKejyiQ49R2pfbeftBcqhY
BhBoXcM/EmXa6cv0r3MZoLa377ScmyiGJGaqOQ9aUqLzpDn2MB+jSE6EE7LnscJk
DfimwTxA4eqztIm5vQqbcFf252UnFyWBiCtfHLIvBVGWi3MgIOWeWsJo8UnTPlU5
MmQzquY1ocUxMx9VyXTu+vfNnTW7IAVc75FtWtPxTn0IBa5Ag9cMHlYoN/Pee4qX
deEEk552F4Q949tzWy+I9BIWr4DmQRiWZJOD697Fc2+beZH2qmcEWFxdE6S3bthR
KVc9Zip7lvtDTpMrUystW2t7f6KZe20ITJC85deC0MCywxhrAWmO6W8CHH8rUQ6T
QxeuT3Js1U5+bQhFy+KECNHBw+wgou8K7aD1fFfUG5gK7IcsHNbPpknBHKZxOyWw
372I9UtMUTbTRYwOmhy6kG52J3E6y+/eCdyU5K3IjViDL0PFaO4Pg7ZGmTxV0I6k
k7MuL46UMjHXt1vgZKJfgM8USwoKwOAyp/D2urOzOvjJ2101ywc2aWmw1D7dxIQa
esG41xMeZx8qLG2U6C1C2D+jCWRwF2qDtOB264+3bWQh+f5xCd68tSzau4jxxK+b
Yq5yc4OfcgnongF8wlcm5gL0QH9GUkZ77Z6L/HWb0P4PRcuJubiiOJMxPx5dqtbK
9pP4I8/goAsh4MJnz/CqbpMvBcpUC4qdUgyrNzYsDiHwbDmfCct+8qPkXl3VxttU
MTbW8SSedZ5y2z0qk8qEfZ4rOeK2Sd4FfiJYsE1wDpMHCzjUROD2aQJWo7+j6YWL
8AdgbfwjOntVZY8S3maxEMHIkDaAL4e4PEIEsrLSA4t96b0ZKuGXRZBVqnXqTWqs
ZM103twdsAF2VG4O+sFqRMJlMD0EI0PSubnoXmYM8afW5aW4CFQqtiMP+no1ASgR
dZESvigKwv4v39VMNF53ydaVoguRj35WVq3rR4j2jGEcaZk8sqWdRx8CzCLbhFot
mWu8AK8j5hKKB9RgqdS441CfFkLcjpL+wZFIQ6V0UAHh3CJprqiahgrrNoisYgTt
Z0yMcgHNHkPwvlzMumr0JdGArvQPpooy5VhKwSQeKMrZbZfGmj3VhQd4Ie+Bok+K
Qa5OY7N/cMWiaVEUqZvIeFJpuWXlPod71+EvQsixTFMvvAClPTOW3I9BeynZoxwi
Ask8+unmdGJ6OJm45UoAvp9PHI5ZoaIkRRhwUtS8JtllbEn4hVgPef5MRj0cUYi8
vV7h1cDW9vePXWkBvWQGfU7eoewlohGszj219cz/4KS7J0EuQ4A3taXkoXZ9ICpL
PpsQa+XKWllB0pnmiUOLJz4hLkihbrXv7SE30jytQKv+PiTbYhHwOUg/XuDKJtU0
dJ+ZqJeFkMvtAzFLTxxTcQO1Ixz46JspHZyz98UFSD8i5Y/8s5UaYEvXe5XSTD0s
6FO9I6m8nGJ/0mwFzFxQLMq6f8rLMkalpshVXxmDpMELV5X0av/REaHCoB47ODzH
ra0nGRWyzDjd/Xgmw43Mh/mjk+al8I3Am9tTzaeHdfNhQQNXinhSGNRuw2hjw9a4
zoyGg9e7xKp4Y6rWZETU2Tr9OPy8mHjdsepkvAxx2lkCNi4ZRKX07Iuk69u/jaeO
K42D9gjK26snZZhglSv6KxTfHDWIo3Fj6daGPqoJBtou5Guck+qbcQVQ/CnyhkDK
wpfEnXfMvQM0KK+LSoQA5UknJhH1EuAyb0m7ZwJ/D8KYYSsWMbbCTy0NBaPZ1O9F
TbUhonQowwjpimYzp3PTyc9PxM3S88ytnEtAkgzgOdzPSSvGPhXZOnpKz2h4iOXS
thLMuR2mq0w0E3q9L5cWvqwVQtYQEp4hCTdKXvnh2ngbu787HId3NDPXQeqxgVmQ
t21QYpKwo2CEko25ZajD/veRFO2976V5an3uOD0xIptbpHcdScxrjXEwm3KGYf82
zdMzmLktkxOj5eas9TL3YtbVqXCojYee5VnTTkqDufXQhoqxnnN4m4zpWklkO/5u
PnCK7lf7lR7g18Vyj9fCZtYWpAwMi05zN85bccsvS2oOhwucexS9N8qOlbvWA6PQ
iVQ9QQmRwO6nD2KzujIjWFaU+5DPf4A0WiZN32VOzUW04YUVMlegpencF7V2TkuE
kvgP6GWwo3wopswiMWR7uk2WWUmP2/Rho9PGB11zYdzVMo9AzPwzz6VFW1kurJQb
4sBJjrfVsQDzSUeHemDizoTbQ7dgcBFMYtxzdbTrcT7xAka66OUm3gB0v0AUGePU
mI8HJxwckE39928Qk9B6JCSfNsTEPanw+yH7n52AHAnII2QonGrhL11cOethh8MY
cQmn4ed+bd/RcwAVb+wLyRAx6S5e6VM6PWAoQj6alRy86GfetSUFICVuZHw3ipTZ
hyp0tMDOvUtJRQHhFKS6K0DugCzoLw06ClVeKP4yAkSbu4Rfk3yA4GTqRbKVUgqC
v0/5fWPeyYAcIAjxCQIKzNpjexBmjo6hioQPR83sIaER/PsuBSnG73P9T+rBbHDT
Y5lSODKVGCc3HaYB3slUACzZR4qKt0ySbORUDYK1cXWanFzYrXJSj8SPi3XDtOnj
K/At1OCtN6ac1hrHcJDxEb20ze4SqnyXoN7rK5lnXok3X8jboLZZJaZlnxLzGdHi
OPGPeEED+xXSzodKeGG6LXr/u6Mp1TVHPg1xqPTWx5bUFv/uBL/F9Nhwl3iw139e
EIE3mDkMVbjFnBQvHRP0ccykMAJPLzg4MIJqy3kz0XP/SthfqIQN/WDntwotkZih
qmasOQCoGapoxjhy/Zdke4lEl63Roc6z3DL8q1Ca9wBWyImwHRJIMGkFU4Rmr5wR
3ZkxWYN/39myx6tsJLu8rhO24Wws8brvKsZmV9ZU4v3JDNtfEdxlNZncf1mrXkx0
7ln3aUm/VAqHgm0PkUdIjDF27eGwGk8W+b3dChRUozSHv+ykwH8T7V/r7KR8N71y
mZVS+GgOnXZb2wPvXr5C/wH9pVoS8G4X64j7JKcq1fRMCX+v9C2N60mfpTHYUC2a
6pPGsH6kCmsO1JpHV8uuYZS1tS7eNnhmvnKgj02IYg3CjyTL3XIGgWXk2YpaJtXt
6EqmVgTlXYzmwtxOwZCtxxwwydQui9JrfSRgG4O0pCvqyRqHGI7m0l7uhkhmyGQF
FIW/TMh+h3DL41cT3KI5pm7/RA0dqeyKfal+l7gPmjE8tQfsUgt7ZrM9QyvXRMzv
Vu62ZBmoHa7mosSoZDGjlzYh9Wb+ygJ+pNQw+OtCQG24JobwMQ9KJOw3dPlbHZCp
OOD1hEqOmNb8eo7R8TdFh3BxOyoPJ/RC2OyUlFaosRhvLn/5S80pyB0ccK5CtYbi
KPGTFe4hAVxr/J5t3gpiq+grp6I1hK0g/9NjPTNSvjsBZD/4CvmFNiHDQO1mg96X
6SI1KYWoGd43V5Ed2gPOCVnQL7N/z0Ys0/DtJ8rvmDxtYuLnMhUc/n53pWBPWN9F
ncJEY39St+zvWb5r9D+6G8+DCv4cRCNd1/o0fz7dI+bk2BUsGN570okFYBrIP9Pf
yNfk4Bzggs2nx1LyvQWhRgEeY7kqPfN0GIyDNXXtGYoFg/m2vmfloV9bvEISEDyd
LKYBAY6ynJzrMr3INjZWpyTQPDAsrQFlllSihFERLsanAyLONlQktw/0ygcrZoBp
OH5AwKLd3A0/uJ61zauKjYBkUa08bwrmzPOPe7PNgC3wvbRmdLTxchJAhzGMkm7X
LaeH/ggtCWfGLMQJMjkgxDGnoBNYRuKBt1eikpGl42LlV/G2NU0foPmRe4eL/p/b
lS5yYb4KNpUgdOXFDLnadGOwGYR79duetwUryA9beaRV2rkeHhVyffcZCvw/fiml
1Irhz9SJRYrvNBrpaJ+aeW73vxAbpR7973csvXgCjtChzNFlym6p0+JXws3bLYPI
arkXsmXOwk1S0yr1aSPel3/4+9u6RMgFN5iKPtk+OUGRX7fp0OuGO+EUVy8W4Dok
Bn7DQgU4vuZfNT69Gw2dHQY+IhTTYkRN2qCxITiwRuUXfz5k4gWb5KjREGw2xuT4
XQOywQPLAIvrDmlY75sp5klX861rxmY3NfcnfWIFmUliDyEwGELlOZVVlDw4Snyh
vOu+TcWZ8JF++5pyNuUAVC2LddtVZZwBKs5b6T0HIjXt3pgmAhB5xmhTiPwb//vT
14GrgTp4Q3gWkjMTbVXHIZ7dvdehoPOL71W9EKN5Qf1W1xEIg7/jrDi4NljQhvfW
DSWGC536qNs8jHF5QA2muD8hT4SWx2DLzUF8koKTIvvolYJTKql/Pu10t1VUx3t3
aff5DNEUwV1Bi6JLyedu/wnlsU0HDsDcni0gwIz0YxFiYQT/dnSm8D4V5oKanv2f
fU+7XWvY1bQiWQ3cuqDBjssB8eI5uU2K/v9pOZSUwEn7KHLB2IzX+3SJ+69u5nsz
qM8SYPHUIyIoPmpTRt9bPoLxjBQ7mHhrL+D1ujY0+BcVxvg2VqWZw8nlSwL5AZHp
gSsE9PuyXUsfr3xWOToTeLlTmszc4o+MsjziyzlbpdHClPWagESTtSEYd8rWgjSd
r86R0zXNJHr0EXKBWJQKuY8/071alIo92I0nuXOeSAEMMqi7I8AB8syAmHBBNhmZ
9gB8j11A/ucLBAcey02aK0W9WmCXmPHXIqIjOPLWfGBb0sH2+PQhdtMQv87aNlDu
sT9s9x2Q8Q3AiuWaLMQweY7U5Ow7rZQnZOctC1IgWYA9rhWbaiYbtlPIsygjQmPD
XomKcXEisoe8DYYh0rYdK/vijsiz7Xm5RQV8BB7eReaUMukXrhjVZZop9zbuZ1IH
Z1Yx5D5kUnvkkatxE7tRwSubYkfz+S66C4QL21ZXT3jqpVhGJEcNIP9l+pvffgfV
Gtvgi6pwFV3qNsd9c2d5QISOBl2tV5Y/eLGqcoEGTaFnjUtP6rI0M7npw2pbmMTv
BTdiGwO31yWDKLEQ8NcfPds+a24216/13MH3tLqKf224IXdbvMxa4f96PHbjIpDF
KcVY0rPN4heiHRInY4K0jbVuQpyRE9NfmXp0D1/Q9V/wl+A8yQGGXRR9Ojr+9jp5
hcfWJFT2BK8BEG8F2Zc8qQmakgMCwYxC9x+UJ3dI1EXmjcnrYbY9M9grq30LzqNG
HYhgKPZvO7R3iE30jiuZ3eDoSUTy1a+l5Zm8HYu+UhfEXd6iOtVcypNxuUERGqtx
M1bxZWw3x0/NrdQdLbAWYmDjUHWQ3GCLfitdXcz9plAgdP17igfrAQ4kDOG7hEJw
3OisZv9T32xqoU7TDUsySh2t70DMKcknYO5/Rg+7DoEwWTwCFvHW/vdXoqc9lqhq
LI9Gn1UY4Rwdk+Ew1vgygwoJ4dEj7NhVXX3Qfm92xAoXyl/MVLUhPfaUxJCLS/Zk
nSlFC45tTMSddyhXkS+Fvj6y3osx0NcAfOcOuOQyxWHqe/R4iWRuTxu9R3mz3hDX
F378VPNiCl5XYARmHaPURqT5ZM03/W6ZeBHYsGN6AVAnQgaeDg5QbIKm/40XkaCA
gY3RAeJt1NKjGGWZw2rxUTmdrAk5UBhWBlcOBU4BzzI1u6QBjR7NQMJ4HapiuXCZ
PmJZeq4uZ0uybbyYHFiQrBMSl3DUkL4HsNizYgBYXA4MXQnFQqCEfIwOE8RWqrM+
jJ7EP/ZOx0P6V2d0DN1XyvXui1aoXzUflAZRaihSEpuzyZq4L/vTAF3i5wf7/Au8
L5UvxwzdewRP4QWBeEXlsFDbODefdBAN6jqQwoxbm/SEzQ8/aDfPrlaznqHE9Jgv
gtib3yFdWSYcCMVEYfsGbq6yXWRPWa0P9ZB9hXBNdbKlVuv+NRHx6r3ohzQduR5a
G/qsUzWNVH1xPWgVy4K8xmKkmikMnERxH0FKCiAcuHxAWiqdoHdWnts0W5yUIF5U
gqIYNnYzQDcO5V6MwddhEeBE8e4TKY5zJFcD2Hpv9L8RAuRCWc2Abjb85h1bpEAQ
smNHS87BhHa5rBOp0idHmcfdkRBTTIC2nGCtHvD6zxwG15iIuCUaqXWoefnpXJH1
eNmy9rDAwSQ1ad9gGFkluqShUpcrKG2dDqUKFUX4xsZXAPxzI7mArWu2QAExZE2B
XNLrFGCMMScp6QNvr/6CxPK8TUUE68HXVmRwUiFRb5NQP6kGs6aTwvdlOAG5paEG
QZr48VBC77l2Q93k+J4BvwCymryP2Vt+9m2G0gjdlIvG88IVd7tV5nRMrwMUvuqu
t1OJnNwOyxFuDKQj7GG2wv+kDfJw7uNzvLKxMf8hVstStcQ7tmbDcNQ69r1GwN+T
G077YfhqA0SpXsA1zjUzNZKPFuapZcJf7VkY9RMRTUUC0DmvMRepLwIbbd7f+R20
2EYb2oQC8/3FU8MyxxsdHzQ7Sjn03u16PIhh4WqUf+nlcE3joFZ2bBt/z5jF7/lz
zvnfhrIAVpFKaCeISzAhc0NesCBMdpeQc8wTu9PVt8voEg/6LFeu6QVuj8NIisdi
2/DW7aIVrqPJlUtEdO+fIJtfNryRXMo9rZVVbRuo6/+NND9ItFDf0gVltejvas+N
pWTiyxAjYWcSxvtYDm5GGoLDJqYafo4fqpb4mR3ux4QF9diYQjYjlxRVjKMulWnD
FycFhzWK8+bH174D4El49v2/P4BEF2TGPBI3wGF+yoiDQ/9NtLUV5uPgo/5jFpOg
YH0ihwqeAxlM058EdPYJXCFoRNyy4MTmB71IuXznmsgfzWGIv+dUvqckgxuo64iA
O+4cuaJWbEGYGGThUFJOy+Fgo5tbpWT5GvFHOO5PNvLYsc75TchNp+a0fORDjYec
avek0HbKxBeueLgh8CRV7QUQj8qh4IHi03S+Laqd/HiwJL6Inc0uYLdgGcNH1ihW
XQEPihtD/uLXFw0JI07cmKfDRvB6pH0rZKCFdpLa5rpys8rItXVHSu2t03ajEEeN
OUq/rtsuaP8cww+rG0/QcE+T+d6a0L2q741FpMDSH67kmQFAnoK4udUlcvYV2CYJ
j2gZ9NKi8B5Wc7NAyGcm/1TJcS2SOTU9pU4u4GTVGofym4dlQ7/6JNLpr0GYdQeH
ZgIuygpeX0bZJKXa9I+TOp4SMMKQHD9doeV1DqiKmzKH0J47l18mcKlH+dHdb9pm
QFS/pcMpdwnjRJMPa21oRN/lTvxrTIu7OZA2OpbMww6ey88tDkm1KDdQJdnz1NBJ
enEolAA+oEh3SFzAudpabQSkB+IfU57Vm40I2/bCx5jPNe/VwAjVDnzzbSNPGfmI
hFjM5oweXzFOgTx90GnfLCf6lkGhXuAXMDaTpfhLI7j2ryL0of+t9E16aeadJzcT
OvsjrgBD19jBXvr8lB6Hyl9Rd/TbpDBwQ894HFkU1If409KX5VoyEGvirS8odja8
LAozItNaVwZ9WFQQAcJ01eNVsi6iD5QudY25AHVmk2rfKODV4xBuLwPeTQ55RhTU
9W4FnybJspy/zbenDJ3Tp8UyUGEKN0bgDvuxtFBG6qeQhyjBSujlkgciV4DgN3Zo
iV9bxD8C81L/77gtwdQaA8+a87o0aDnYuBxWLdT7rN5ZGAhQrfIZMjAZvTKCOg9x
ptvOsTQcBNMx+YhNZUXtyfQXr/o3ee4OBbMPT8pOmEDGY2hUJemAK6jkyFdiIhej
2gX6qIYBJ59YKTl4vZBPkglWM5zHpU60wGyxRjCSXntSqdl9+42Cj9IfTjWyUTvF
w/JR0wyCE+QtpaQX+1Pj1O+KtyEiJj6eVnglhmz9QJZgDVw2Rauk6hJxM4F5oHUH
Jn92dPdYqC0W13wtqertsJUWJuQuPBBLaj7R/DwVc2GdebKf50BcXe65b6BwrNdB
FEGIbH0XbZZRti2voXcr1+ld3UenAcunw0nZZx3DXmlHDDlnBqbd9Ofg4W9yFqS6
g+4/f7rrjS2fKKSxk5Mp3KPvgbBAo4rIjJeMFVmkPdkm+O87kQwXWbXsDRMPrSrq
GJ54zNHz74ud1QaxEUHNPfjiC1hvrkiGPspRAojTiTKM9v/XByGZmM7BNP2TLybp
hX9W9HzBghnB1lXV/1nqK6ssdWt8eRATNaSRFp2FnJFbExKrQkTrb43GD+eGf/kw
3fr5ycSjx/wtYq/vChsCt7xmbbIMR6h6CgudSUiPFZMhUUL/s2hRC3HeMDJCWuH3
dikEyBBFH73WrONXio1VZ7Hd5E2ZPwXgojwdZawNOe6I07bZ98Kl6dFw7HelLsmP
4bkMZYjB0rZNAUyOkxcDsBF0OkP6Oxz9N2eL6fH3BQwEm8BG78CEbF90z95tFjWh
w0cAanxQQoX4rbdVoz6Rx7ALsbJv7bDO7uWMZ8Y3Vj9diwOvH1kj5VFXgb15VkGd
4xn6zXRPub0hEmT53dfQ9+t3GTe9v0s7PwrIvzqgJ6Piia52B39oyyrK/a5+NKCn
g5FyOIhrJrDs4gsNg3O3dke7i9DNYkRBt9okl6o42wAj/7Bxj39aPhmzgPNkMke7
MCeQnvXF/1eV9jVac8of8+Reo7l5fpwpFMSxsbkJZhph9fNffmaROzTIiUV2J7M4
E0L+6vmBexTuZYo3qT8h8lx2olX9BLAJ7ynEovUeBAlNhT7D6W5blRzp8xCKU0OA
XK0nlwFXiAFnbdROFAZA+sHTU96PzJEaZQZL7AYPFZCGPURl8hhNMhxuKXQ5aQdl
lvC+5SKAt54ZKh7q+assiCXKfcTr/nx/z6UODIIR74e2Kqe3lhZ7pphNhPAt+C7O
tWMg14+pkvHbNeAldA8MIjo8WyIWqpQjrrBSnweVikXbnBjnPT6P+D57vGstC8eZ
3Osfw6zIUmqtAZhOMVXY6iEXrctvROxNK/tI02QBoz4Dgo1TkUbL0UJkaWnyFrLq
edsTNA96/FRraQXIOY/3izR/99QxEMS0QiHN+vVjK4NKgeUwwgu3wBMqz+Mc5lvT
pxtXO4bXsa+jxN7mPA6PGISLHRcnv/YqBt9sP1LbEKZ58AcAHYyEHGVnJmTMWe5h
JT5ekRoIiGnKuGgn0HPbAvJDoyZEBDLKBstfYPqph3mivBVaPAEFcQVSfp+Tcecc
Fqy71cHJzqosvFufgbOQObRN8xApW26+9ymnXeM6XUiWEB9QI83mbyh6UAN+Rhgl
G/VWM8NAzQIiauxkt8qQnKvjiI2clSWtkyK5QGClWwHzCbm763vh145jzfZpcGJt
LgpxGRaYIPHJQ/Y4nwezieGWZngXzC4BcWs38y4Hw4tTTNyg9hCuPkxKNqbZ6J4A
cbB08JitojNCA0z7hsGg+Ejk8XPQamMWXJEsAv9OknXLZez9dM1Pz29hakKCyZcA
QLi45h9xkwWpwscbK1EuWZb33ltMBsbn60D4TmM13+NLD3+k7ExAJIU9XUocg644
ICJvvfzSTX1mylYLVHhytrH66+03OVrAZjwSLEI3109asFV2C+MPDz2VfqHxk0y8
BVKK5U9hLRny3dixGqbEt6gOkZ4lSSBuLuTW+7NO6Jrsscb4G91gpSJdqNK9N5Jm
RFEVtSPapaCjgh7RQ/J9SvU+P2nHyTb5ugC6maxhYv3qKR2RM2L9Cw0Nx9dupEB8
dH+T/BgtpLZ94gLKaxrc+yIb9fJPzG7ymypjJsqHtEEaQjhdp6LnXaauB7Y5HDYU
Kj/XYMQ4XnBSQI3zy4rb3odvRsCHqU+jBIyrQzyoLwdVwtq7nf39KOa4g4VWwXU3
GqZ460jmBKX29CP9Py7Awf8NSJovJGQAfADLQvDuplu7xYT+XPIsmVVyZf4CPNsk
3k3ZU/a/2YXv3A/nLZcksMdjDBPezqsz1xtDiPQsKrF/uI9lkFP5SbifBy/uzHh7
/fHPc8dyd34FlJXtVPp3SLH6wsAM7lcbiOSxy5VyJ5LFNG5AfFl9SutgN2yeR4HN
bwsm9WUNzZIOgwQ1Gvz7jPbYa+C5v5LWQlWKliOJQ6APJW6vbUSb70jjDnigeB9l
Ox0lgM5v38jTszhclJOAKwdJBFv866/piJTsfdUGBhf/HCb0Ai41wwZ93CnQpuCX
d+9OQlhXgAvcaXSZgQLwhoplwl2hyd9eX/2b9x4hMmFn9GD238hN2In/2sEz4wKF
BxlMPak5JhP0wPTdAX5+7E/AauSgzuNwpqepdvmHnpI4DlNEfe+uxttrmEPlA6g5
zhEXEhIxPPqBb/eluy5CKkZeJXUBm2bfv1rGVLdf9YOu2oukJpOrWnaGf7DgeqRt
yxVDZ5qjFxcNroilarmgeYs1JiZDUBOAlc1/1ksa35lEYdC6zFWv7NxFa5Ku/vxM
WKgJtkt4dbaodqcSdan1DHFrj20TpLyUFlHd8t+7dREOjXT24NUyJW48kERNCjRO
CRZeZ6Am4e5NNSxD5vsM70HV99XsO/0Ex3QKpmU5/MBkRMYaEZNYN56lN7Lf6EWt
9XFpePywb9ew1l/v2a60vBV9pct0NvLYH90N13cGA0wEqZTvJ00PoYLT/6SJR2tx
V8e4mHTQz2erWqqz8/dIu7GPeY0tdrfWYgl4GFo4eTg8ejPmwlETJExf2bEsvpyY
kig84D5k6CYuJ1mZ3FyRRSMw0PG4OrAf2A2gcSOu9sUpiDKOHvqXR12iS0xkVS43
ppoBQb6UVuMb7k1KaoXdyHcBM5ZZbQpnwvjSeCTDUgBUuaOo7CNMywYmTYbFcEty
vNLErFMc7eBjYB1oHc9imSFi3tqN3Qkoe8+jWOLAWDGnic2tL/DyRntOqAbgQk6p
XRfFwMLs06GvaVNwPE8cIQl1/37LBpJ2Ovki5s9yNsRi0ddTSYpGjkCG1WvQeP1S
ZCtAkfmNyXALrdplZAnTg8ooRzwyIn6EgpoGrBtEJBhGoXcJvMZsoKOfuWzW1tZo
YeKf4N2wHBh/SSWSYXmrWgioleVbVXx7xGgW6uqZBWPNUtv3PemtmruHlgX6Q18U
UkaACr+zpX4Y+5rkou2JvM4aDmBVsCfzcjxERfEfmgnbSV0LETdcTN+msu0KHjXD
yaZjZsn0SemkaJTF3qjQEfjG26VtpCDClRLrz53IyyeDoTCYOowTL6dFj6SjcV5Y
8rax0pJq9XcFEBZ60ZgpKipPuP09krnphFxSv+g0sMzPBSmqPGPWDltQMtj5v3LH
KfEJT89ytA2vOaZd/MhT+QdqsvbYFGczVHgO5AhJNcKG/zCxta34cJyFzTbPENlC
AcHY7Huug0YKZmzs4n0EKnqEYD5kwhVOcGRK25eFlK6Ar5s6YU0zcwHOvDkcbHY4
DZJ7VwDmHWInak1QQkn80ovxiJqLvojADd0SfvyGTpn5mi5gKmNJjehPvgiuphRs
PTsdYCz0GICCNHIdqQsFPvHAaMsvGDSP0popDfw72eEn8hvaXbafSvhbwfoseawU
9ywm/fp6eBphXaCpsotQvxGTyG+tb9nuhOBZXzHxSHJgqYrkDw6feaESa4Y+2G8s
t0JyreNZmuMUbEu6TxB6R0eFRjhQJdkfa7UKXqTt0GAwjFLhEeC8lMvZo+tmzV7U
86cZoulY24SVHEq+Ia/L+ZsKFCm/XSnSYWHfGatGNkHshVbsgd4ktjUQT2BqTaLM
kUnZDoQ2z1NQh+BSfn9NsBcXMj51dotXNnMFk1mi6KhMl3UdzW4vR4ptORa88PjF
g0/IjeRav8SeEGzuLb/VIJVMwmRQsP7i4hU2cdqiapF3UtesWJpjQ3Rdtcc78DtE
0/0BzJgObtTnaM/RMn8zXITM5A3hPwOelBXc/PsyZQVPqx5zg1fUSuLYNX2PLh1H
Nbs2jGG5W/ATzfpiJ07NyS6MXD7snfVr/uB+tu4l+CJhPjTzGW9sZitvohSo1Xwf
biBiNLyPwyOzZQ1oYOBOItBP3wZ2ZJfWdLgwTIftJQokBDJ13dG7k7+6x9iekQQM
x6TPHO3w3NiTZl89XBG1OMo+B3dAjqkjYugIP0UYuLnnv9H2iphxjjcqTpKsSdNS
ogq+YZyJCrQG+6ledUEnkwdMSWqREjrBaccVAVz7S85nv4FWM3CjZJsU3wpX4Rt3
iU3IfFf/WjNMxT2lUTTI/Jp3pkCtq0i+5fpiOwpvMd+jwaHU8s2WQ4/kPgDflzER
1h1NlaFU2mZwlrVa36PHer7VSW+nNUcqBBJEMdQw1wHVZGWCcVJdzmSrzc3bwnzX
zPWX5XM0txNJj2YvsQ/AhTiDE8q/7qq4NiNZ/cYGTqlXHP/2MjpdbtVDl5MdsGrx
Tcl1JbXXKOZjW4vLVLVs1cYYaEUnr7hhq66XuymZqL+khBV9OKOMyTHCkdpOJ/m4
RjFA1GuMB+OspgTRUmF+KGJxq54qt4LoLOcfEit0SVBhjIqtGmZ7xBOjFsP1wuxk
ED3PQA01s6TGEG7w0Fxopbi318UzdVWhhg0K5vwO90Msz/KR0RWflSmJPHtnhDNJ
UYG4ikPo7t3Dvh85EAxk2Ni/+zpFBYNfUh6f6wKsiodMIbZ19kFHomJ9s1xBWOqS
k6LoxPeDOqB7EvSXZ7/QHE82LwbVRTV5wYw0zgxDGMNToxHkymULkV5AV8R2wU27
ky1QEMMe15PpiRCJ+xPJCCYZ7B6KgC2dFwfwSXQMNc6SzHRc+KLT6kvU4CvfV/jk
XBpYEi7SzAdVP9B35MK6Lb/lqFbMrx1ZyiwV0J8YnNHYh+RrbeFyyIroVkvqMEsw
7MgDceyyRo53HBfroaZhxFgNxltMxmMedK1XktXUpV2a1wFP+m7K/W7suUWV2qar
6d0aIsGlCl2EmP6eNozneIvYcIkRMhYbS2qFQWREWqEirqpWSzOllXIMI4BmElLV
AXTYVF1NlPeNPnoJLuWbl0Is+QrPQNiUHTLTFDq4aEOW3uxOGDvXBtuUuMFHQdsu
Bi1P9UwtjT7ZasMTMMHVi+nRVV0RL9zPYu7N4y3dOJ7OznJKeiDVRYjGmpbhDoZA
XRYgWrkZx7rmwdsm3QSZxzZJmbAtqxQMwvKFe58zMLi9BHnZZMKTrzWPk4HuVPjh
b6pln6nif9GH7flOOeopgNt3gA1w4nfZ0bZVYwnjaaTJ/Z9baEE+NvqyglC3c4Jb
M4fCuUGhLZ+EPGBtc4GoUc8T1FuQdWkG5mbsf+xEUcm5c7vxDOAy6S6JJa1wTjVM
eO1XpjF9vHSGGrGB7viqTKOC7EEqkbXelHCRYokTRQH+xC8Dp6AO7lxlE3eixSRK
j0l7DCBoPruauEiJZbfMZ8BiZCSn7rfA1X1yy7vokUMdJeEKIcj8bdtkg+Vi06L3
5NIV73WZszQFEMkYaV1ieXgIrQvaTQqdhZ7a3C5qQMPvwNBUUAlU2Pf6/AqRUGtB
J26nFDUEqPtsUeyPjxD60tccU7KU5g57Jp7MzxDRfgrZB1PrkxPLDAjJnVgD9O9o
CC6T4cI+Simp3frPX+S7w+SgR02p6fDI6jTKgd5+L+T+HWAZmi/K3t/UtSPkReY6
mglaEhrFpxQowHjZt2pJlZmx8NpQLp+rC8B1dIfHGPiUmve3aj5Jd7ipaKvvCPto
ew3HDqJsT5oXczo6SgukbMgefJBrj4ISFzf+s4mCHiiFqJBkUIlA7jHRqtytIzt5
mpHNEfOqUzcXlu2YlyuR7e3eGk3pSt6SRs3dwPgiMWwF1qOLXwfFdyV+pYz8Ya9K
YkLVzfGfRkj/5X7BKwoq8JV0YGPh16OQ3HBcqGY0A+5zxkdvn6p4F5C572RKO4SV
8+zIfI7BEB4abv9zkTCbsoMzYQ5//qFlySOAGJhVjMtQFixz1ItjQBaAwUVxTrqR
C5Mfqo9n9TGE/hW2zDfoGNhgprd1veJF6Oo6oZ7E8SwUlB60stJGkcrVFVDgwXDr
84pjM2WuyGPGJNDn6fhnqw8EzDuZ/zVjsdnclZ+ylIWHyi8cAOTYEkYwxPhLvF4w
i+UTahvWaIvNk8bnqUuKXeL77Z6hdbwqReN0NwobxrMwOg1pIoOnq8zPY3xjMs+I
fh5o60tH/jCDrdvJBUW44Q0dEq8EDS1DOXetoPlZ1kXC75aPZv+uoC27KWyrvUFs
BzKFFR3dyC7nPeQXbi2TBN4T78FHSBm4ZQ23mLjQi2QG73ld8+QriD6xLu/AWrOd
gb1zBuv3sCCSp09L61ha3/m0urs41yRUgf3XW/EQOPtaHIK0zlu7wUkqYjDYjfNd
ugsNilqJBVmXOzbMlnI+V7pQDZPwyL+zD1O9iknGvtAQyC0BG/pZ/Uy6/kH5lFed
IJH2/ufybVnns5OUnLgssBXPJCOHPjn4QLe0STjO6n6RkXgBDtTQdwzhDKay8TAU
7jgK8l5w0Iy/VecAUtCFupHi7gCmyrrtBzVg6LpQL/7qUxOwfIss7cEFSPBxSDbR
xMezAVriw5IPf9pk+Rd2U6vk/ZXKNwO05gFszYit9sz9/3tjhZyYAFnHZ5TaSNyW
imxnwzd+hC5ujbr7Uet0gMmo0R/fJNOcn5BX5ZVEipKEMAOH3YYZs62CL6LyRl2k
DcbTxW9GwhMVDhAK8V8QOgKhsyrXo+FaqGPogOvSNoOeNoVcG5k7V8qy/cxwz7kA
X3bbiAxGN+pT6MFIB3qOV3VAnREsDjBWmBuoJlfx2HFBUEOUMjbEEdo9CAfugLAJ
tRfstI/zFIYCctAWNgH2m4cniqDURwzSAoqw9+sRk3h2q7/59WSDcNgk1WEAYU7X
zefY3piG9uiHwdcgMRrxyKnrlI7P3LN91Jd73JUnoe1awM/ToKP6PTZjxuUPAjfV
3kwSkmXOmA5LXis2+OibYBpAy1vAkN3q91Gkv12kwooG8DBxk1g+PTyyPiWsunVI
9rk0lU81ttUOR7MVGhDZv14F9hf+nxgnVU2L6zgkTf19ZEy3RGAo+iFBeOZPqmG5
6DMf7SUJXNku9QQg7NOs3rnnjYszMC4oBTqj8ekods8hP4JJx2+fAXujrGobXr8v
jlgcTF2YOHbLKWD2Vv89zgbLaE3nWMCYlyUW5BQrsJBbqYrqLF6a9Ff3RovbJUl6
uw1D2GM1WASiZGTIVUQF2YL25Ug3t3AXQtxRG8+mgWZ5t68ZRVb22z7yxMVXrypK
uxMo28lQoESbLSm+7zl0oBXOs9+opQidr7SRKOy74DZfJYEQGczAtdXQHCFr02sn
0rkj9xTBll4aWvEvekD8IikrPUtcXREzc905H3LDatIjXcuZDHkWmzvvmympmUsY
g4Q6nyChSQ2decKrMxSocXlrh0avAoxquQV0sjGJGeu+dxJDpYNvJoUHdfeTtGcB
szXXtiKTCzVCWHE419zgmRGhoUDBirINv+6MP5tvvBLF9g5IGEHmNNVDQsE8UsTP
GfWhRhfqPB6EZZ9BgR4u1x6Eu5AXKKyTU+okWhk7eYq3JETdGj1qrik0PHrE1ngB
s7I4Y1LUXD0gfYHbummubOiP95TazuurSUQjFrmOfHAj/mZuNHryPaX3r5W2UWZJ
K2ANtnLtQY4cqzY7D4Z3vnjeYt6dc8S+aEQwuqOWRc8P09UFnfv16NxtEJwppEpp
Svu1wAvnYHOIFg0xzxFOrH2cri5M1kstRo5yZZHuSeqxwKbqBzyl9OYtPb1SGG/v
DusvV8atbv4/On6iy0IsgGfjsY0Hthxy8g4xtyZZc1rpapWZ0bQy/tgb12tgFcvQ
6tbznVfeu6o4Ws64kDCtaEg90i+ZxTUw63jJPLwFbNX6eMLLR8/RyejTDqd/rTeA
N9x6vyvEghLxTyNwJ/zp/utCEqf3YUPhI5xb+oH8R17I9zYehwkBxsjQM8ks5Ir1
YlSOTuZXp2QtMOZtvYG9xaOqtn4+BkdIKs+2y4RRo6GlxZtdcu5iRHVu0roj3zD2
1lJg4rLK9HYLHz+qWns2/aAlFS976/h6wfYmeuh8ULdBTI0ftZm0v+hMswFdmQEN
porHjPVxnnBTQl16Oak7MF/uxXYdxvCmCpfF7eiIqSBfkMfvLyms93gx9+5EoU7+
oefTJplcyxb2vk4VVanktlBAcEsMfVrcWkfH0GVooM+TcNW0z5B6Z4hDy95mBF1R
oDF45Nsi3dsbppDk3+vP+AFheOBtOFzozIM/W+IhqvYDOBwxJWtOx25omDlu7V4L
a26nR4xUna6xhZhalCwSneotLT4fGNM8CotpsiiPAVrl0y0oR03nzgdycPbMOZ6j
J9D/XdDWmRMXM8At9WjRGIwD2b22DIzeaZcbX8rNiyHBgYo1XD0cPHK1q/kOuULS
R9xDC2i2+fZMFnEImR+nfdKn+iLzeTC84wUZYKFs+UGdTNScsF9SOUv7LSIaoksc
/XWqvQla4Dr/lfH5NGNBpizHZw4XXhB3MJPYpobKgb+wODRrXO8oMG3w94p+6UrM
tXb5l59ONMzgrvOhF8SCFqfIee2E6C+E86gzP7Wwrd83UOFobCk/cX/DzHn+7FH1
WXxBsydCZWSuQXMMG7pChCPDShYuHCstSdcwx6Fzo2KtqAcGTBHKdIexRLCy+85h
gxguIYG+vI8AH6Hls5xzmuumR2opkBTAb9HKkhk+8uXnMcwa1eM+6KyK3iFbeHfQ
Ppz0rC26GtrLls5+FtIIq5XZbo359QZbD1yS2lj1is4ACZtkSTX2CsmVxo5lv9dX
6gGdIY/e0LZ1ZSgmKFbG+MtMW3TDAd2Al5O0LHt9gryzh1+VqBIptEwfhJIiwndY
75Yj4dpknhxVHS6TKB74DqSih3OFWpEINCWGWcq4Qv3xTQOy9yozHxw4Jde41pbA
K1fQCJHw72nyjR4hvovzdioDfvtlAlAmXf230Vq/sklB9uF8SWd8z0aqkA1vFYd6
FNc31vc8ByUtqQubNVuUAfz2T4uNOkndAN21FGIkrNjk4lvNU36l8bwDDlymVF+w
8rXkIEMMtPD+vuBT/MOdFqn7VzeH5le6BUZ1sKaud82kJavo3CqBWjdd63gWuiGk
cffy9Ve+s3CyLUXCDqKbiR7psrEkc5/gOU6A8SJQPgTJol1lQph5NO6KrSeFc6a7
cstE/vEbZ9PHwUpES2XKeA57lBbmN3SZn1NForuK+kQ0juECgKmlzM+RxJUGArUg
vdVLh/RvTPwIgkJ78clTTxJBsmyuFCijZsWztx0AAqqltvWObF/xCr0EvIQmMx6h
rEuFI3qMt7Ykkd/NOsFFPp2mF0kAA8c8FBBWYsdkIOPznCKCIzq8odP8cMr8Rg31
oDSTdUE8EyrWPIvRwVU8tRHSkyvO9YkEl2Fvin30kaNcVApXCd91lIV1nRJmnf6Z
HZovNxFvQHOoZARFQYhPnfRSwLZP1aisY+kJd6FrF9MhivOQIJL4lPTEaDEcZle/
oHCn+WnI7t/oLaucUpRNfJrfw2+p6qUtZFBRoF/Dz/dmUstX4YvFQKnOfDLakl4a
euFZspM/hR/SEKO0pUIBAn7cUYqS/+y0BFTZsIFM7uxOQM9j6EnztA/FSdlT9p1W
uvzhmoGH5NqEBfWTr4XWx7Qb2Dxq6xM+AFCPG6cTG+w4qrQeICbEoQo6IPvwk2dQ
5vG24Cw1wTBCvMin5NtUWSBuWFYQmv8VqCObUIcqtspfR5yp03zDl/sqkV9hqtk3
jvUZOrcWPPcYGalh8zfxCXwidWrta7Pd78JbuRw01kbD6Eg1AVJsuETqPNwUiYK9
9f6DSa9/UKOIgTHjFxyfLYo66e3xaLSbaU/ZsteGE+JGXhOTNubqGjBZsYaQIa3p
D4SfP0R4JPiusvcQvdLUm1bivPMK0rQP/aA09jOiaqfLB9joo5Kcw6caHCKE7IRe
kf0h59hcpBL4v4AGdjv6elFCz8Z5h4vOSMcnTN4xrA1TstH120Q01UeWnq0oj/9f
/Y6jwdmyNoE+xNL+XalYpQWqKwdoMShyDCPYxXzeFxiyFOJr+41P7k/0xRsGOY2b
gkcJzDPEQOnM6BdqTcDcy/JYtKK/q25ei6VQONYHX5Mb0jb/TBTln8YN3jbp5JhH
OHxPcXC/O7qmqLiQ+CJxuG4U95TGXwZKwa5X7+rBa+BErIBfVGD1SzaKyMWd9cWk
r3IafIRFaiqKV90Y2vQNgg34YRSlfwypQJcGPQge3S0mcDk9Q1VQMumGh6D5duZn
Yi+inCB/3xFlxMyGictHp+KkWxnBJh6OpX5zSaU+RMjahxYnAEuP5xX3ydtAd4k8
ZSE7cAJ+v5eIKsT/4Eit0QAkDRsHgUXc0o/8w5jDYkduNP4+jmQifsBZ8UIs+CZj
NfQGE/L23JZlkPSkPAAaA1rwjahwPPbve/L4QJjE2r8qAUEYfhChtl/V1U/VItQd
3E8HsLXWESsr0JP2I0/R3IPjIGnYvtXKf4MLVzT/7DQ9u3nsRIjjQo28ihFC51Xs
8zE2cisOLVgOjkuF9zqd52RSJhaomxsVKcCE4ELSMtZW4yO6nzgBY2HdnFQFZL0L
D5ZmpgLD4tC3CwHkmpZL26W/wMNigeRVpTXtW8woP5BDyFmpRRiE27RSojNk+Jr0
pknPLafOchJZaK1XNBvHwEBNKXOPphooYAABDfTMbK8L9RDXOSs1RPz8Hles3Fw/
CNzkGbipcO9USEJbDT5w1aQs4iD7OVrajRM1Ac653Vil/huzN8LvQYgYVUVu66sn
yal0yvdE0XLtm7+QxlUl1Bjg1CZ+tuFgCT6gmTXOjujCpUDoXzs4BNG8r3kSgf2Y
1xVkowIiSv2pyu5AeESDzsgCfCE45llZPkO8Z6ri8zdZo0CBAAAIgLoZOaGpzlyR
skJs2hVul9E/NrnKrHod+OqZRZtgY48oJnf00wIj06LnTvc/P58+AyZDCaGOpDZ0
k0/zkRN8MZck2Jvf/bewKelOpPq8bTtTMZwNp0atgqXJ9eWdZjY5sY69oLIoDEkn
UqK1Yhndn+BRE38djYH39USxc/t6+Fn7hFfQkIOIDEaFY4J5cYxo4PnSeX68SI3n
fW7/fGYa2U3LRxTVQH9gu7F6Yuwewo5JvqFbbBuyoA4FX76YTTMUw609tlra3RsO
3KotbsFVoXaBptx7IaqDVptEBwN4uINvSK40ZlhBC/QhiogqlqjLyuBsbJsGYhq/
0vuSXWtGwsFPK8o+cohwSmhSH0aXSn06OJMx4x9F69seZcOOG2/zMZwZAn/XxYPk
LU9yDER9zdN1UMfQETGFIRHLohTRrtCgUZCRSilPk6Q0oQcEYsN68bKEi7ayOVmh
EHolJUlxUsaSy6ZGF6vPeUTEY7aAA4bkMfcjkqOw3AeYKLeslnT5VqtXFc8qp34a
CVAJK3IB9Vkk9dlmaA2Pl8ALnwELU0TMrL5VGtf3hhTjKFB3QzcRniuoyo2X5icn
XgYSaiYeVkJwq9O5D8L5/Xi07FGwqK0ajYu4d8CcRsPO3UsF5RTxR5s7dn4HhZCv
e/bI2hSzPCTBcN7ZZlT1v0fewIvZG74rtpo57iGab4mqrhlyauj76ORgnLHnkPOW
HtE+xLTq6ieokJHqEb6P2uQ9yGxIw985WcyrjXHflUSpPkP//4oOQSgPp34AFyoZ
8BCnHAC07t9J2XQlX1D0nr/FmZoxwJz+6ga962W1oZy2yKRwBy86jUapgnm3MvaF
QInxG8Gdn8XS+u9iLFcYWmJNGLjER/os/6B3okeZAN/RDMErg40tDZp8YXGuG/bb
9LCpZgRw6DYgaWkXZXxtemFiBV4lY7f/200sBshkbpaAZR/fDSFjI/0zi9KFnOsP
kQxSicG0gUMO9gSbKtKiJXH2tChlQVB8h5yI1I5GydJTmire6XC4wQtWJw06LRz/
SrI4jcN1X2p09bCrAlEeeaXrDfQYZWDYoTdORpYwHSvqEYBK05LqyXPICHss/6bx
Eq6FQDyBdnMFEo8v+0mo79tTDN/QD7G6LV5B5Q/2I7cYxPAhwvYa+n1OaP0j0BDk
hOpKJPk2Yp2UChiXRSNsfCGdJow9CxWdSNd8HOWAdQp9r0E2FN+moYsPWsJaN7e9
b+Kn6FShBExGnJqgG3lLSfYSA83Yu1XQSAOHIXvWIidJZ7IhYE+HwaQCebBsVT9e
fkvS5DPcQiqBAkgEUXR5oK9X0t1qNwYchnWLq8s1dzPm+zHBL+U2LBPx2cLmTuvP
J1cj75agrpLymesSNqLXVgk9WdJ3lhzQbO9fmTHzXfT0xcKjpxGwcd2U0rRzAznC
8wjE99BSolYwJoaAFIcWkYBoiyLMSKI77m3TiJ3GQA+iK2894bnv3mGhjeIW5+4X
NI45dY0Z2bh4koy0q97JOs95d9/RyKZ6vJRwdfs2kgU3lRfDrbSZiXzJpNdAgHt/
xqaJWzHRE6dDW9sXtVYSuJuO2sAKCRsUL+KNp2Fu139D0C7CoLaVncYOA93fnBrt
j6SyarQvNmkixihgjo4wKL8H0+UVd9Esg8xEv+p29Vmp7Iq7xCWUkXwpx2/SOAL+
3XFqDMCsmCqcsNYg35z8mWcoqyLat0F9TWrM2GGi6EYti9xU072DbRrqJLn9+KIw
FU4F3mFRofqv6PcWPpIHD/w1nFF7eTethyKRnXgPiZ45CeXCpQMgSZguEizTRFl+
CewS2vaRiRn8gjhSD+voeevX83f4LG68ZzsFM+xJcSMkOHCqrDVEGXp8Rcrcm2zB
VKAB4eW/ipY2h/e7GdD3tfwmcdvs8cFPrzH7qbfLyFRe0XHPm6bIXl4O5TrRrec0
shN9WOcshDiUl6I2eusXXtSYt1wjso1aBt5btrf6E3znbCwqIqPgAT7t3ABywDsz
rkwvm0gNB08Qz9egCbEVSRc4V/aaziq2jgtZuWLwvHvml1wPIAv5Wv4r9F15tzI/
wAlPHM8tWUdDyB+hfpn4jnEZqODFJJmId6Eh02SVdCcuO2ftIZwiNTYQMC7mNxNM
qsTU4ugkL9xxT/y/mgCqJkt18/4U5/2SYLKOwOoEeSHxzuQfFXG3c8TJ7U7I1rt3
IoAh3csJTzJ4K+44WYF1E1C7gA8iCmXqTA405F+jFZTIzqyrHm+enBpA+mCh0uy6
k4s8yUKcBK6lDjAaPPcHfmBWam11L5KuZ0ECDgmdQtZ2mJQdM0iFu4Wty/fRC9Xw
wBFZ/SnBayka1foMHEdf4rDPq0QOP737YN+69jAp+EklRFlOL5UgcuvrYqd6W6AJ
/Refxc7DK2Wqq8fXyBG2VKD0lnRUxbR8D7NbfmPwNu7tFlokL5ZtA5Muq4qneN48
figKjVX1MR24spZ8YlH+VrEVTIansh+COwxieLbaxLfQHGnDWB/ozeo2uezpLrxF
sx78uiIvXpkzhn1WKfnEY9QVA03Cy8nl3EMhw1gJxvDCtphyLo1lSeDYNDzDcCOW
U5YuS+uHHsPW7NByNC6/3ezalgn13FBlmfJ2pwHprpIoWrXbqhFaupvmILcbCc4n
4AETuxiB5ckbpVy3yPArS9OD5hoCanGFNefoJrd4LdVbZ51WAhHi1A9iB1JZ98fP
iWF0PIqTINyBpLTyQ+0W/Ab8/f1mEt8YERiABxu7zMbmTS5b1R/NDoVszOx/enUF
bbwkmFabnNMsk+EBPiDCl9JPi4fFRrtcWQ1QWxo1d0JnL5ygLz5UBYE0p9C4Wbkw
Kju7G8GAiG1zU83ogKprvNzO9BuAICHplOIz0dcZBT00owG8Oqdh0ZI7j8sWXRfy
AN4L97q32NluoxpB2cgLXhQcRpmhACyM81mU9hzcsTa6tm9e2IJAw++ZYgmHpjAo
bjuMoS7ACuVnjxDIP0mfllp3YfZIIm1Hq2N9LweoLCADX6+w6eKWf1jedZZzlKkT
1+KAl4du9F5ctgiDtqMt1BElA6+or5XqW5XxKbWBF2iQOC3wOkNpKd1Pu2HnxtG7
qJxPkwx0x2WwQ6ZMrCYpNagWSNiywqnQdTciWEccHlVmBcNyGBQY/4ngH/mtfDl6
WQwraMiuqr7ee8VSYVN0cp5w6tObzPv13udwWj0GIbkbQNtY9Dyo0yRa1OefxEXn
5Zri8R/96q8kTF3cI5i4AjjpMGU1CBMWYFc4bcRWYDTxjhMq26AI1SpFZIi6pwpo
kcyQD/RsCvt2fcWdHh7QxYWn8jQqiUDAL8nHsm0j0Kfw630+jw+dNI8g2ZVLSxOp
/1KUqHuuaiUYLBi8QD7LW6lzJnLbXS/vB6BigAjzSCd1DYWzdY1lGlJMdIuR1eIX
Cs2mu80w1lZByAhp6wkkKyC0Ikbt56eHgUEF4E0fNS8Z+WXm5LEPeUSVqs8gdeYo
sh7KIsG3kC7908wHWVVRB1k46XxUSb0ybx/piZnGL2HgjAL9Os8Frd0GQ8CD4Zik
OyaZXWWS2aXrgLO/SXK4sbFOjGFdTKbQ91Eo0uFV7yxySpdl0i+bM9hVW8xZeD/A
UjHt38cGJHG4v87PWYRssEBpuVWx460aqqlmtatB9G9LH0vkIRGie62HLDvK9zdT
U7QwvQEQ4P3dyrJbIaI0Yo1EscabRIEGSZfKju9FuxxgqWcMW9HG99L//0JObmsi
tum9P5iZUL0/NT7sgYelSL7XNXYQzWdKSH4ZwN7AZKFT8P02sV1J9Akw/ODApn4C
TMQzwQGf7qKVPTHWxMYQDoiWuKMpEOvqvP5A46PsE8S22WcXpavHwEV+tCG2bGjs
HR3vnCZqQGV9Q2It45Dmd7mqrh+fK+7Q+RP3WZMmT0cDJ+1Pml7CX9HrDZHpZ8sN
U70NTljT7jdLPTtbVRnQcDW2bdjb6LL4pwT7anF27p2tm7WNmQrbSMPtdRhzmWku
H2caRvK4CfdUsgFooDoQb/Rg+nofGVF9sveviXkRSmorCUJP2JbmS6PyhU0bw9m4
eLFsVFc45co5hebDeIKtjrEo81rfPA9dNn1vqYZKIcVI8j37JAuB9ZEQa/ngSstl
AQKSh8ixPjnY219doD+W4yL9Cpw8Lz7AbEVIDDt5tFuzqYriDxu4rVv6Lv9xFa4K
wEE52y8qoiZU17slNGYelUegYArM1PGdFSshmpTlir5GaDoDfy2iqKDzGxkiYjuj
j94rvB9SZDkzIDwMN6bbLOqDiZDVy5WZzCM58ik4K6CZpXcz0NGgqR3ZU2TjEhqW
8sU9sQnv+qr9wg3k/TmSSu06bFnpZCgJh3zCzrqZG3nPXIMadHZPGKfk5j35QnYt
G+Pycb+xvGN+7WoJQpirzXxYMpfeRxlvxVuNqzRTZpx1JjzV35gCsb5pKg/pAvwx
gwcI/PjJHGuBGLCZ27Ss51yzhWu2iIUXUpzF9BVko5QZT7P2xzRt3zBHLU1NFzpk
+5nH476wYTrPDZaqaM/f2utRoVCodmazmZVnP4PaU4PmV8Z4yGrzam5JYgMEwZgB
3D4VI1uwS4egxNdrA+cVE2XynWhDxoiD/vdEzX4Q3f2GSPlz2PVMV6RYOGIlhnlv
Ulq0qXQbS1Zo+v53Ylxc5EfXmso45KJ/119tBhnmjuBhdmIxbWoIG6VaPPGy6RHI
on0CMEXpHES6p6n8NpzLqt4p8C0BIhfI/F6sPHhyNemA01i6nVqJraZevXcjpvBP
lQw88lbf37zdejRLHzKC9KBHrMhF93IH8gvo1ZXjH4C8diM5q63sH9hWnYVM5I0r
ymQeBX+M1nD0prGGZxJBmVXwVAor16TFJiL4GnmDvyR+clAlhLX+lWtDa8fcMD/V
eTLLnidoOqqjYuZ4iYx2ZFyTysNAlqumntFSZjDlPgMcqFIfJxMK1+AfEy3tFnW3
slpPJJp5MZomsr3cbUy1DLkx4yZiJM2s4MIv4mqtYwGMsWa3GIi6M1dYCsPwMF2t
9YuAR+LJ3TGDB8mPdMWmKnUvbmY7UHfY+Z6GUh+GB/EOC1JzuSmSQzrJ95GC8lSM
pWSpW+i7LYCFFKShOebfGUe+2dSohE9RWMl7+6pdYDaUOF0Xwz+HRhCbCxbeZfXt
YKoXGyKThTNBWHpUXfNeDgYAHhFZ7cigwUUUlGP749cPpMDwI3D89y+YAz+1Zey/
84TOUtQqGybNwiFutbLHR7oSPYDw9mUb5W+NVypBbvt716sOKUQXDhQKujJzgVqs
TguX8jtq3tpdOuO6q1O+hj4h5R5vsmSO+aLD1IsnYILgTIuMW2fXwcqVqegFDOTn
IxJJ4xbm/bBr0pM5rFXMkjvYSeoWpjV9fepEBhnCW3uhUc1Ogsi5JIg3Am+J2rJh
OQw8f8P9M47L59rHR70Mx3fPrM3W5waaFD59HDt/e3bM0JzWpVHyrVexN3zjz9cP
FsAIlnBH9fUctUu1BKIyPIv/FUnycgCr9UyyhHkfHjzbh3jlBJQmrtHaV7inlgPI
9UfJvQXnEynrxoknQjeCrmD/D5pQoch4zUs+qtaIwaRsLLnh/qOa2TyRO12QvSZE
YjbaT2f+iRHIX8r09xCceJXDd7cLQmzyNEtlQ40xdKIkiWdpX2Zk+iavJo/R41Ie
21kQlEi75mB6foED1zRZ2ulL0ff55NuSx69aucP2XmpX637vukAtuXZXLgqWMu39
lSWTJIMK0hl9S5fhb6KF5of46chAT12pUfEFMU3iUgia5WeK3HPN2jQsKD7sBrxw
eZ+vYeUZHum8NiUz3/rywN0DE1FJ+8oqVrgLhL0OdQ+WF2ccGZ9uppEuYJ+bjv1K
3kY2JGqOC0q9F7XAksUFwl4sHqjUOcEzMVMHDlTOaeZ1i8WoT9DKM7wvgpizll4N
3Wyqjz06b+K/jF5QH1s3Fo9T5PeK+zpQYKvvzL0it1bvyoX6KhFHF9mLnTUOYUy5
smOuI4PvfQ5fcLrbzVVqQSzcMXNVVdzDsqZbYLuA6SIky2FkuDQbAva/rNNmIhdR
ArA0TaYKYpSRgd4//DWXJk32ggm0/mXxncEHAGrXhv3lq5lwVXOv5OoX3c2X/2d7
NA3kplc/dskFizPZpT87VwrQ+DNsNqnGh3P8spDtngPCKojzNWJZm7G6XNambEa6
63qjgwuuN5ywkR+j+LZx+dxprShRwcAIaYvEUJFhc/ulhwB8j5qyT+G6w3GfhN9f
zOxhe1CnSJU5XIGSmxf4nNIhPmmZJVXwTJbTg/mjvgxQ+7Gl8KDvMWyXoIoFw0le
T4jmME2lyWdIYRvzkSHqjZSB4VYlsK5Z1zZ576/IhZjmioKJYZ6WlIw8HZbE7thm
fm1pf+xwtGBjN5YZyfxd5qb9I5inDDKfiAjuuwaQ8ewXatXG4ci3x05fHxBzZ6ZS
w8mXVQxSQf0s+7nfrEaZN1MbbtWHCiZjLkLqcbUWwA8E0l3Cemez8I3Po5m0yxx9
D/koL8ABfj3jEA7qdtRcNoPiZzmM3llF7+qm6CCTzITh1BpTTs7fmPg42g+qPoXx
3epBEstOv/sP6K+2IIwn7TPG5dOXHxC9jgXU6NHwWlSQChD8zOJUvQwoIT+dXvSB
3Lu1WNjyPG877/PM+dKLcVfiwZS0g6CvTP1f214dfxzN7OzPXXNoqLsOYEfr7WK0
NzIRHbR7K7iGK+cfDo7jgY16BUbt0qw4OoseQhwPGXxZAOBajWZSidqfySukfDHs
7CXFXmwc7MrPxdDKZIfbzKyFf8yu2yeGUoIfdW9CdlNUJdOvRYDtDNYf0AHpox7+
AsqTTO3FO8eQ6TYYL5ny262dIDlX9vuwt3g4x5716YeWQHqLaLmJyh9BYOL0wcyC
iiPoN/OuKTKFqViYIy3y8dS/YOCRVR0t/LySVQ2dpLsJLtsax4zwOJ7v35XHm7Wg
AdoqERInW5QnOs1oc9Ll/JwTzCrLgN8biij9fp2gcY/ZTSpB931x7RzFh8wk+/Yo
dtFBAb8e4/+EJthrpueIVK1mXF7kw1zC7BiLlItd/txYvwwmKt0PmNMhrrco0Ii3
2vmbD5yB+D9Cm77MozHNDKssqYHb2UvKIOX/Zxg659jtvV05W2V4Q26StLufzSQr
Vfthbis2F6zG8jbQqcvis1MRw4M9TCTwM+TVSV/LmSk7hLVI6QmazZIO4APSd0ap
q78dC/lTp57XXoeW6euShR32HOrhg+fmcou9cN6Yvnfy31tpcmQIAQEQwnSI3gxw
spmyk1mgOoA88WUBMsB4T7r7oQWEPN1iFubxnlxRnmY24rUQ780DLgHsmxUBbF4U
ZXuZ2RznVmzDmPUkKkVUjhRjY/9UsuHQ9ABB5huNZPMMIUMAJT4XkfN1MRHLXpIG
KoT7jgg25R8H3DzU/Y5sm4CzvYqKyYG54NRne1WZQb5T8I5yGBVcyYFs4hrWNdqM
aoCoQE5MUhMGS79NNErNHaVSga7LJ7K29fZvMHrdNHST8NTy4axEs7qoebZfxoCn
XrI/ha5X6t38SH1PQoSUQsyrvE37Uojh1ux+MEVHVgl/EmoH2HCQwgzxdBmkrj5x
0HBZTcShCmX0r7NnAy3V3l+AkTSGA4XoC0tSqTXvnehy2kIYZHC/YM3tw502qfZU
q4tq0hNIFOBKupDZnxDDGIKjK/2eQ1xKqOMUvbls6n2Lq0+2GIHJi+wTKDQddLdP
pXSzfPNIZrRyFtZafjCfXSngJnelOeBDFx6A29MWQlOnFkqCid+k2f3YYT2gpCjD
imSLYVWb87VDW2WC45aUiPkOlFdWU3F5P2AagDiZt7LkP+QobNb0Fn/KKY6Ao3L5
At7V7Q4iFBARdHr6lMYjaDiIrwaEptEZ5MNT62nK3uGD3Yagwbtkd+Fg9vcX3Vtc
s66ag8Y+kYf6gdGPphK4Byekk/X6kxKDBrboBpvH/guBGhTH+mvpUzq/C9uwqN8w
SBn9vkj+cFvs6qh7Vt6FELCegEvamcLdUj79w4iv5ooKrDLH6pCCkAmTV/xmsRGB
fuHN2eKsQdwMwaQeWdhODsTc0DPtowVXbbYW7i3X1R0poVx4q1Ehsr3Bf3NH5Qmw
HJGeCGYw+hPWAa9ag73WNi9mHU+gOg0cenwefbmuTdDbhBZ+sdGpsseZLrLUiePL
QRpVWlMK2hXUKJ5N9ino5WW9UMD9I5JUSiSk7UHG6wyqQ8jcNIdKFb0GciLCql/f
pLxJN8nHoukCol1sS8PBBO/lZv9oboIkrYHSvkiw1hkum4hIU9A80g8JHzcrBB6G
eISIT+zJzlMFeYO04x+RlaCRjvgK9Y4RV3WfQwgVic9PbtjH3uGBaQkEqW32yCij
WZMTnksPk8DLMKUb6BN7njTzPlVdm9+4d5gJNNg0Mo/kXzGZImZT2LmGh9ijd48n
e8RcAjOKJBRnm+9xTqNW3GVMhjAJs+Y9YrOckdAlQ0WwdA6KVKPxvxeZlyERtnry
LiIKVjSOarsWOtVgE8DgWdf0erbL1+K2Hbfbrk6kdMRBo4PWN3zF4qPM0wQKvq3K
duN5dnEWa+UthtAvGwU7cWGrX/iILlewqdBjvNkbCzmYTNdl1SqEhI4pRenz7BCp
GZfbjNXNIAyeng4Je2YLi/imwZZYkZ1fkTL1JRETrsntbLZP0fJlnbSgzJBlIj0S
MJABZy37kxam/EOOcj+MtULmMHNNg2ZPV2TsbHRPE6ZsxKizJBS6eYTYFt0AtU2H
bBjgEv3+BT/9/hUEFSTgp5DZnPNVc0emP2VEn8LN6hEaPfytkhXeja9KOkqGQex0
fNxwW2bTwxvgj2UVluyWRNx4RAnIQHVsPPPjuyf5PjfQHaWZqNhv7Yug/1pPWU/M
3Ew02FleXeynsax3AMme3vpXBFRVsrIpbPwc6Y+OXe5lYEPxzrJZF960c2ZqhZ7a
l8CV0NxGLYgcyeHnN1/DWA76j0iGOhCO5KXN6D7KhFml1C6o/30Q45bJgbF1y9ts
bfUsdVndjdaPp4Ufog54JzP86A24t3LNwYLb0dEGiOaLUVQwW4Ie3+7SnRDBYj8t
fSOodRo+yqroewOl/0qATkdIAA2qjiRsz0eydFCFHKpPWYSJkR5Yxw1+l8nPZ5A2
6XBRi1GhbVxG7vrJssgDugUpJM7M7DOu6YaOpDNIwxMBq/FvREXf90BaJEF9tGfn
StikDf9y66hdqWVbt0FAqs1OYLtX6KbACV2ugYsrgG+Rd9wjokTvQJQ6NYJL5qOk
P/zukDmGzMWsfQRnss3WljqILxwkk0WnKcis8wE248CpdKEYHleKhSAFFsXLwNR3
cgDKaNH61fb885qjY7s6L8a4ClArMcgFmQMz/fhts7mDclrbfapUK6Kjx+irvuFS
3tm7oIjWUCOG6CBc4TnSILF8QRsoK0PfkY/akqEW5F8c0aYRE6/idL9p+/PyQ+4x
eBeDFYZiC7zraTm2wiyZDo/1jrwWGFFfXpSTmeLG6IPHIZQTunnnuuxLvz0AS0Jx
POW20BWpayEjKK7rTBMynNMzv/12c32AgGgT3ey/mQAlMMj7gpvN3wuHc9iTccJO
Z3XG/A7PTr0ZcMYUWRAg5fO+eMr7+FHiwcx8BxgWdH6GEY4fo6yWLN9l9ogVZzN4
Pre3yZV/kjdEIn0adIl773rh7QxegSRY1GS5a8IGJ1tyDqIUWkz9tnkKAyINSTde
3WyYTpOq3SCZ2g/f5npsF95oi4sfss0BeJHEMtQSAbB5H0yOZdWVpHsqWncNTQG9
nuiV6+zRQW+iVQdtcx6yt0f3ewqhyP8d80nkdRV813s4UVfgs8LcZ3GhFag6bnMe
bc1uQF8mR5UGU6BtoBBI6wLQvFtQPCZT0W26bUQOtQVys2LwUOdb8hs7aeMDNJHF
/DNOQuBt+25DlH1LE5v9QHy6RMX8vtwA0LRQpsUd/T0LYChlMrb7mJuFLFyVIwNF
kbXjdqWc6k0Fc5Qvuu+EWnwtZZSKlQL2jvgz68Z7ejc+j3PDURRWqyHot5lSACd0
e0Pc1feUdrxjcrIcuAEicBqWrJ2Ym1bWjutUSAFs4MKa7jMp2KiyA/ynr/RPoK/A
WutxRE51mSARQoA3F9NVSCX0GuVUJoB6PK+rkshZRYAPw9uK17+T9vuMzk5sOuDV
ST+CwLO5qRaFzN9Xz/2q/6Ngyu+CSrwC7/L9J1/XzUKHi9TME9rOlmZ8SutycTMO
cr9C14eBwBmhu3+9W2t5zxq0roW4gNZeLuT2YOSzPHu/eoowp6MAQMXTDrsIboOP
4yxMHATZrkbWSO9P/kalTG6L7A601IQD2tE8b6v/Upj8zxpNGTRfNzJqUcfRkrzR
V5N2miBHa9jCIZCfN8k6JCZG0gTzT1r6nUFaF50Xu/nyNdCHPzOOBwa/xTIfgW9y
b/hZRB9IiR9qwKKUtJanv1wcbMnrYDrfGuVeplrNxHRZGRFtocl/3y64YFQkF8aL
xTPfK83UWrtn+DQzCbKQbh3qVWQ6X+E3unuQICl0lGR/eozXRVXWKBOIsiOwr4mX
UDlz8W18XBT+Pkp6kPQ2CRpfbLj+s2E39M0RHK9nwQbpVCZdXYHMGrJmy3HcOUvq
R3Wy0/S9p1Q7uT2AixytOEjwf/pY6P+10V/2stFS0CsiB8Ka0pASuZUlf7i9f1kE
KFP0B5qpTOeqPj8tp1JCSHVbVDlQbP7RTITcJVfnaGNMNPdC92zyGRI5rNaAQrIO
JyNFu5TUCTtBQS4jowewdgWcFPPjwmaJv1G77rQKHvn/Dqus+Z6wTTiZfr9W8EPm
usLWnecIf4fYrwRDFD44nBx8pGIGpMc+uBBqsx9/A+Orz6gjVmguOCE2Z3NtG6hX
SheYO5M+MYhADe1H3AeM7F11DFd4PPU41OKr7Bjf+L0s30Q+vNtiaRHDg4D0vJPv
Nt2+F2L1ZzxcM5d5Q3ZcvbtRan6bC8mX7lUYQ6ey4tBty/A30v1xtXM52SZxCsGa
BJ0jSv/FBL6kv70pl0GMn0xJlSIsAk5dxy8980nb9vq+naCrv8IlA/WCEuT+imNa
bgFUMgiFq/RSS1HnDE6LC0qpSZYLJcWzvkRuYOQIlzC+5Z7g4CXXRczsHaekiqkc
QGqtBFZed6Hk+lrQ5Wi7svEr3joA+3yPhasQ5/GQtLe1NnMfLAPMt+XjAjyh1HjB
kUIx4OaJyO9RN9gK10jKjgW+wUW4hWULoZFDsCwMf3TayvH0k4RCCuo0cByfASb1
itS9dPs+JbOci8r+hUsoKNcF86P1AdW7/XEvbrlV1ZuOqVBLguL/BfxNHdOp3g/Y
TuK9LyQb5nIDptfIfzleVn97w/f8PCVkzDKbmh59FtUgNFkZ+b5ndAtFGgt4dvwb
LfWeHHuM+joA9skhPgOPUORYVnqbe1tsZnGj6RKpSwTF7WRMmRIjIJnP0jS3FztM
sAG72WL5v8pHtI++rTevxKITrv2X4PfTjSDgY+TzZhHp996GPXPCzeNko9swhhpV
QflDTFhouRy+IaYbEoFwiYKbS+QejaJkiqdCr2YZ5enMoy3ZpkhssMEVPZeMAzWC
bPyIvpuoihs3WrOulExtwUFqgs00WB3LyuZM+z/EMszz53IIlEdv7al7bJk4hcU7
4xcN3EM1rQyMW/k1LQAxCIUsrTqsSp0VpqUTfOI/sJ0LzpJY2u3rfI9O6uzD1KFH
b3MMmkIRGqpxW62YmyV7LfT1JE6nRbuEPoCKwgjgJ829hEJlWLxPowinMbhcDGnP
Dzj0DjBIluSOJHAJB+Xhy3NjZhJBFxyJL/vl64DSduKbPJ5y7UABqIh/PrnZI/0P
KvykN9e6S3LkNPS0hooxV9NxEi8EFm2o4G8/0rt57xiiE2BYynqMarZ8WYB7gOnO
bUS0aC4YXd9cn0DlQ6DxTA0dkHC7Wc+wfKVxWk5DJwbk/7QcSrwdTudCRNOkhTiC
veoGWr5gRwBcgqHGaoFI6XQb4X+WvwXBK6K7n+zeUmsoLnqmjZng1DPaqQu/0LZy
b1lvtm+IajEo54Ih7pjpN376pGUyHIZR8TitDreiWiY9mgL7NVK+qKEJwWfCRssp
OSyptjIDju20Pa8Q9kI+RYJD81joCqVR8da817+71zGL6h+ycjyrheb5u6A/XfQ2
1RLWLMm+E+yyTZwuhtPlb/9KO/iS7C/lJdX85tHk6Slr5OwLkcTPaoSdh+fcZ4gZ
Ih40X7klTHBD3MQeUCVajsBCyfLs1RM1XiRsS29n0DFoaWGphYqbtsBx93AKKaMc
Eg6Xh4Zs+63ULlVrsKFZjQxwKOnh5/N9P5FU/vdabxl/AawaSwFXKG7W1Q+u3OX9
FejMPWmoCMI++WY14BJQ4b4Q6I9QZiAcMa4WiqhdrlpvJ90pMPy2hjR1FebWTOhG
qi40nKTK0dXRXhCZJfDamLqN96mMWw/3EHiTc1H5D4HfyaSpPFQPsXMLlmB+7TLy
HghqElZEFz1STRBHCvR9d37VdRITnlFAWN+pRYyK/1AWGbQGw/azBzjuIJ4kkBhV
IOBtlxmEiFGceOr6cKM2q5eUxs4hLuhzP7MunJHaAzGm8rgW3S0adUWD9hgXTmdK
/07U6QM8H0Ir/PFo9cO7V/pYZv5BpQrWLe265yHQUmYIATX9Fc5yrR4GoFB2wfNe
9cRbD0711KcJ8vnIEANz5rQbwCkbUpIi/Th7jB0QKMwx5U0HDWirODOWq9/OuDjm
h6rReo+7h3Pk5qsP4uipaZE9XCLzO/Asz/HTNs+wUvlrNYFEceyz5b/xG2WvpOb/
CV+M39HrPX4KqqIFejWN8RxiSnX4NmxbtUOAzEiUJKTzJKVq8PnP87JgDGS7SMsA
I3LXm7xeC3Ok44o+BxtJDSxBycfLKzsf895/tQDUtrEsHvtktzY2MXHzZ3hRB9Yv
F10LdDllGrgBsvaFYIkncz0lD9pD6I9vFRrr6uFQFABpJWZbDG5ylke6SAqFwLjP
j6M2gVLttw18iN7EFwKAEJpu72C0wEueW/zjlsRgwwPh34ILZ05ru/fOw7g4PmKq
m5DdVuIoxoToykFU0a/JuKkFqO+jNe9fU5f01zEFv8lepLf+fgX/+rF0Hrt12n67
wyv5p59Pq0IlQiAdDXSt2CyINWDpCLB02/3Wl0+tYmmqOrkcLUJHpy3+n1J2mvHD
nG9g5vGoQCbAgPGr+m1lNhe5xiu2rITHLtw58ekGFmr392Nz6xOSMWo10vZTx3CH
ZhU1GTV2IgzUC3j950k1Bqw6cmun8cIMjp2Vs5LGCdcty3Uf9gCvX3ddKJyBy2z+
cBQNh6wP8xdPJTqfM5Cf3HD2Y/OkeSKb0cIdVokSpmCqlxy872xz2sbak5LHU33u
l/fs/4oer3htNs9Daa21C6ng91KyrD/UdzQFLAIIeuZaaKkb6PZa1Dj7Me579KP3
Hb8YqYIRIR3/k8l2AWxgxYbSBoEpP3BYZuNFTEgdu8+5QA1ZyKwGrbuD5GZMGm0i
Dea63LQZOkocvlEZYoUahQzHEobiGZcc/wn2G58tlgopHWxlB+zxUsfgbsfHqaYt
U8WNSCUnlJHa9VXvMlfidClJbO+0ttRuXpk0tHUIwp533BH4MOALyMRyZabguOFa
XqQVUl3BDbUZ88enRNeMwpDCCvhLNYBVUEa2gQ/OLgw1NF4p40qw6opp60dV7OXY
50Y+Iz14SCkwKYh+oZs2zKGcYo/mMnyRy+LtPduWzATXnmxDG5iUx6SP4/xtpPOb
PHK0a+MPkq9XYTv2nGN+DMJFu/U21h1Y1q2J6yhdh+VRvDKrLKk2EzUwu1rcp0vx
yJq63yPfFOL1XPzuKgG0I+fBugf0KczaI02W9uttxKl27E5SjkP0R2FU5tT0Eap3
HlblHcNO1b6Yko50wBKA789huzL1nO9dn6A0TrXN4P0Yeo/DzVMoLYlIIM1nFy59
cLmo724ox+PAo8iakXU46K4JMVovqxEgWjGDpSCxwfINGqyrNoCJVEbx6ijJDR2p
dAxz+OgfwB9i7ZYkCUSeI74S17+mQnnCac6BR1pG8QFMlzvb8gFrCZVxJyUKp0pV
vC7dIopU41PhlBS1BrKjzeV/My0woe103H5PwvZjbx7rbxf7hqyIPp/Z0YExi2LM
wMuOKS9bNJvbkDkU6F+9DQu293cgg8VDPOmwODCW1GbLhOQcr8j8UTRQdV9uvn+x
+y1KOFgFBmDTMBNC2gw+HYsU/ip4sDLSLA3/IBs0BV4srViy7NwaHq6C4N8jePwP
jmmc6NMz4dgfcXEKxCTdFxP+GZlK1RXs6Wk9EsBtrFfVv81DIlY+6LhrRzqAPsH5
Iny6BaoECtoSuHzi37TPIDi31LvsZKFWIt42v6L2wH2FejH3Ef3jTBelkhcu1Kji
QJ8pBeeaZMDmzGb50Tc3fgjufGUAxuikbNrWCS1hr5NfHDfZeLRYFD8qEU5GzvON
XS7UFfMQZwzF+smVrsaJeCwhUbwUNNqgyANvWg3xWJEyqZqsJ3FmcN8xqf31U5tn
kIfwyAPO0XkPbF8iHpjWI45wmtHJD4+QE5x18WYlPNg7bVNZpwSzA+tQZyHCQXAO
GBikdXlzxo0WPrArFl66IPKbGZPysfgeEznZVLP/EL5j7nBEXX2r/yFz6bbmMZLJ
D2xapPPm8U1akLAc4Epoz11ZdPk7KNb68LsIV/9YPlYXYcqdKDSiZKPnQSvVx/SC
wK5uVMr4I22onRmdV87NO+lQUQFmK63uF+ZzX5JDgg4oLR/RWhCoJvPzR4vn8S3M
tGk6kubtpsQs8qGX12FhsoOR2x9gnvL4obkcCgQaNZrkv+Bvy4nYxbZb61ZoTkG4
MXkK3eHJzHjUzJxWpQ7qdJSGk+pQ8n1KH16PCefo9Ub0/Wg/dxlkah1Wz160XNJD
ViZoBRdAwohURSV7bXjoqrF7+Fml5f9pjWQT7mnn89oQZhT9OSYPkq1VZzzM0d3y
TAirnE/Q/FtmTaKw/bt9Zg1pY7qckhv2mYx+7t8/iZPBVqixSnCbkn4cdtASJVB4
w/OFqWxcl/gkzrj3FvNl9JNuhflR3tWfSbeYSpBUUnHubq+bCW8sGB28JLX4l08l
ajBmsqO81zRs8WGRBLn6GD6HnRVFL2E/cEopGW/58XcvdqmwuXymb/WFajeZsnWq
G7Q9doHieJDcHbhGZi3diCYNWwxO++dCZUDyvJxZeY/HH7HgVwaSFcSzfT0nLmJy
fmbQ55sGwoEAXwZmmi2Vd9/sznyg360ZwOnOR652FxBQxgtwdG9bDb1iSgPDnQA9
r24j1gOrYSvdFg68PEC67UNt2gAdXaOeXqr4WWG6JDSpQxI3KauoeTM7cxsS1xGy
by6sjEeWMyvvds1wVsEyAxY9pk365N33AXcYF+GRuwTv5r+i2hk26wxTRiaxksp6
yIDWCp3gBhhyAy1npzLBMaVIiNTRpQmzjyZ4babCMvJicJe3kav1ZGMy/MVwIbKW
ntdTPLzpGzTdLGFoAed3P/yCLBhgeFDUmTj9haOm0j4M7iYQRo5dRzbf3wYYbJPx
7GwOrVQGw2O3D7XJsi2mZLjMDK+Akt6oMR3+vzN9C+9i24bE4WRrd40E+GauD6wH
xQbfI9x6uKb5Gl05AV5WGyb+ih7jrH1z7buDAMv7/N+Kku9GHk5yUU7DKepoM5Dv
O8BshiGFje6f++xJfYL4ion/95UzXcENwKNIiL7IGNzZ0oPwZmEGhuPwQdVuAWLb
MJjXFQtsqsRU12mq6lvb2PoO0XYkciWynrWIPhx2xg1pAPSFk0Jk0fvqUEDyYh/W
ytUQjwRZsRGp6uLzgjod2WQ75EYJLQbJaK9AuWO1e65aQUTHp6wRVUU0VQaTZQb1
nicmOBk+WJMjzcvnC7Ag/BhJIO+mB0BIvDs25bQvA1JS8HiSrD+YZZ3f9A+tfl5+
pPi6G4ZYh6mAKpT8NnNwrwpjbHckBYahbBNcVZr/PDOHey5CltRbLu2d0M+sqKoq
ETOm4or7NNBmwegYimYZjM89DdKltDjKlMltZMxRbnp9k5AliR0bkbSLpv52PgYe
HJDndeSl3dXWVeEWhtpvJnEKp/kMPVy6TUI6GrTzbirjtR4cEeDIwq4WBHqDbC0F
1tZGhx4CMESu0Ds1+RMKs3koHgTqk4M7oGD7e+uqdE5bnNccxhPSELTDWuiquDu/
D4YfG3RvEwK9jehlc84PgopdgbP/0p8Th8CoWzyreRQxWyyRYfjq0GAynXyi9ZVS
CFhGDGYMIx0mNnSA5hs3n5j0SXLw7HWzIXo9q9vMtQNtBHqXttd703KMUIwb1NDT
fO/J1oH+UbuDkBpBO0Tz8tGnMwM2GeHA3rfrqx2+lync16xTtgmhA+ZzXFlnn/Ty
Jx9KMaDW3EOGLnmFjIqVY06FO7EkXEqMOtMdADlgBaQW2b2D7sy1TZ55/E4ytLS2
5UROqKctth3ghjxRSweajumK+LIcCdZFRZD8imV1bEpMi8R7Pi0L5Zx/VRyWo/pw
diJUBFU6ewrqM1yUF4EG+4QU5cudtoPdTVS6n6KrQ47FRMvH1f7ziv/Sl+SBCMx9
Yl0+AuhEk82dm2hpjdZiqyhRG/Q1uNfoEMu0/dpB5mIfPf8nPjvDGxoWEgC0+rXE
GBVaE/BQQUAk8Exbu/MMA5SxnmQzM8qSRk0ex1LOhG2LiZSMAXPpIbY0WKtoLR1B
c1sC+Ul1w62BFPgWhQfMGuCrRIEOBtt5uMNKAimZCb9sHINZAuTYH3ZBatV6BbH/
OS8W0abyLjllycYEP2520nEK+OpsSYkrn5s1rPc8R7QtgNsO1opv2ZAcnFzpilCP
AbGRYyWlu5kWrpv6ouY8KQdQxGW04SsJuRvCXKkd/US90/d4lg+Q6ktQzLHmwfvD
+uaMY1t69jhL8z0VGQ8vmJmYbuf1BzKbJhzt66NEMucxzFcwj05ozEcSr1ENS0s0
JLezXteAxwM6Q/wSCp8P/FuTzfG9Imk90CeI/Z5zyvIOUavdKN/6wtXG4Y+H/hq4
ZTNBWJq+fyCa7p2U0FdKPOteGoeRCgefxODfrTPxNePWtUrvJYGghhmLnd2DLkex
mhz+NtK2kDLrRLmWRz+Dtk528bG7HmJnFJJNQnXr9RTwjwJVQOjna1/1RNQwBnu7
oSb53+50FB51Le2zyZmVmVAGGw2ci4966CGhaGugMZPSQEH/Wxw7BcLn7M9VOmBR
VwJrtqMGPbud8uhqXRR8QjRvsIGKrI3TNFxDxvyIz0caG684wa8BXawWoq2QOJki
h88j9Um6dSjerU39bPn/sZAlQY266W4MhNdCUxDcDgyoELaz89rDElFVwwwZOEU7
lq6mjHdAFD1rMxQcnDvkpiHGJGKzkbGyYeK+H4JVx2lYEVcMZD7lBW2jwxo9oqE/
4GcEj2Ky4R93aUQEdUTqJLzKjCma2WkXMsj94EOu0DVkqyQq51ntt/j+zRXnfZk4
xe31i0MCbO5II3tpEO95S1ssvtqeAoFhAnC11yEiuUhLmcUJhJa06lOjZLehkIC5
sneYt5ByF0JA6L1rSzH6Kc2WU12QBgZKpYVsImEizW4s5HlypwDHtoBLiHri2eY3
rVLKqJzkKMWKDRxSv4Ru0t2ixHXd19NxIV1Khj6NlprAyNqQMYGZERv1xu/MhrAu
TFROHQAAA3fNE6sxqOX6IH+twJGw95KsSrl8OSaJ9L5zkYnp6JIbv0TOn1qunzCf
jzb95NMJnWssvydVu5YyfofGN7MNl0BXiuPr+qXbhizetnnxGjLqA/2vgbTszZOi
G5xvhUca5NjuNvaw/lak/y/pSTISJSDlv1p9g9/j5IfkSX05HWmAGVBSbJqG56Ey
5hz03iKlp6ltvyuT3gfe2bBoO7JHNeSTDvylaOsMnRZcJxhpIH3W7WvlUOEWc1r1
OUUouloFmwcbn16bRGBcTgLdJ4jx5SaRUK1MTe9e0BKFgUGg4KdxkgwWc0u8g2BQ
5/gLLrUrnKU2Weh+XLEwUNYec9CR6/wDU30pFm5k0bdFs3ysAoneJ4LarQDJJ5Vi
x5dLTR3ijEPhAmaCgYVBKb3ZQjJ29KXZ846fSFoXiaL+F0Hm3Ce2QNTyVAINMkZq
kNZ581MpGFeZTEiEyH9QvO2+tV+YIxciqlsvouDxN+ZBWXMEklbomsqoLNU7grT+
bkhrCIsAPbnm6XBQ73U9Eox6T8dTG3hIstW8ig5stuE6uFeiAhqU7jvtxv3dbF0f
QfWo7EQmenyePjuiGgLOZOSClbowAsjhOmcrmMw3WuLRkpstd2osjq3uOkg/hCEu
jMgHWTtXilupI1Cq8f55rWYlSgo6rs1HAKW2/QE1VNjHYZdmyEyNmT7qCfkhGqGT
ahb/hdhUcHp9RrXc6cKJ4C0Ojb/ZUA+/Qn0aBh5aMSWZMEGvxD3luWxY1A2fDBID
4a9OG5bsYS2FqP8Mwr2CGp/AGC1ZLOIdZ6j1Vk1u7ltK6PRGFk8UDeLp8RaC8DFc
+B04p/I8iM/ggadGF+Lt4EpJH5Vydhc8OwvfWzP/X9T4hdS5Bk4D81Uk5jX9t9Js
4dlYf4cY9ROjlZ4GVv5FZBTgke/Xv6v8zqzgyTjTAv8Q+RVzSTI3RxRPuZlzQZu/
Y2uKHlhOToPhOVOTHYXdPdVqjnTbIK3bO7b3pp1DWn2CvdSWguiXX2cC/ohlAEOf
Hkce6raX4pofeOSIcKa7gsejJdVpnqOyg16T9CCFzT3k01napQhfjw6WrdAgTS5K
uD4uzb3+gS+eEaC2Cy6N8sRam8CyaRg+Nr1s7jAbLf/9YVB2CE8hfuSd+XknCwCl
Pn63ZBKT6Pjozst3lXcNFaqvJwLTZz2wFI2TScPEUs4vPK7Tm8Kh3fQI/rk5iwic
D9G10IHO56n8aw+F0fj6esO5RPCRTMW7/lgErneuaRv5bk0wG4W0Fponl32LQ9ok
Qo7ONTSPm65DZxDw1pyHl9GwIhqEfMZllt5fiY8Wpz9BHTTsH1ovA0q8dAKasQtI
yePaVYJWGZagM6yaYHzY0nmEPYR3QKOd1iHR2Oy+u6I8iEQ3uDf/jNaz+pGrmFgU
3nai6wyCJIaOwEde24McxZ+p6TOYUsVpblRsFYurrv/peWZqYMj93LrDrecRZ1UA
aGwVlOL/EsPkcCh5+7qe9fjRg4o3LtogYQKboUCFhGTDi4c+0hMF7Hq41CwZNW8v
RXe0FZZhlPICc1UbLE1GVugdNgMyUQuRVvl9x+ZkqtrEB21g7qDOnNce99rc4qGq
8C9M9lJ4MuBFhbgDjDzYmDh9eaxGw6o12Lxp/RopNmZPw/wPToQikyTj9n0mLHEd
Ka7j3szyzf6mWVVp1l7W5ex+rBsk8AnKQMHCJH8wm05ACO1Lq53IAgZ1BFhpKoN5
q1VzfwZ9OslY6JDE5ft3fC06PnzT0tHLP1igDd6C0oVWQ0NBAFBNu/wPWp57HvAf
epwEgSsDNC3f54LZErYB9+FZi5iRdSUMW5+gI22fTf5zTJbxEThoWTG+HknCqoz8
v3fZUrIqX57+Y3Nxdu8FIR8Z1SsEp3OpwzIRsOedPI75iS29MdRJ+qBo8f2l+vcS
hR74p8xnT9terX3HXGU2qcIkxbkwRhgDV5Kupdc2nCQJ+6OIwWQLoDLBOTET5ux6
SftWddjdSOTqpJVJ7VR3sO7jI891eIy731jrntjaH9WO8spfvMV7v4VW3BADNgIO
QhASI81r9Ahm7peO+hq47PvdiB54pBI2ULSY+5sYTfA6Rmqq+HwMzi9LQrhEP5Wv
SZ9WRQXbz4eGsvcp3n2wFMI5rxptJpSz8LXLg0J9/ixdPokaIJnFvEvmXyqkIWOi
4zvKf0jxOWpe3XCUzJfSNSE++eEmK5RAOuzsD/UjrNiW7myzMAiAQ49qks9cefwv
elHWE0+VF/E4sIriPCf/poPTxCUvwpIF4Xcui0xaWFzxs9SzsggHCkCb5xqEu0MO
pWWfWGDwGM2x9gkc8lK1Lj5fzz1WHUVkLhkz8XZGTxDpv1hPN/3ruUSfIDwAhPJ7
HqYEjmihT3Y0Lui/RbPTrP0vClag03/wd25HiySmHfJVurh5JW/1v3Q2mSQSIwPo
SSmqHn/XNsYXn58vzO06lIUcUMEDCJ/20oHj9tKVN7+SgnBss10cEOgnZbeSWJdb
sJIUwZ9SpwSBfJn8ekJmBVXtQHG9gPOrE496pXnZZPdPl8flMEx3V8GRQjnZouvT
Vl9XYwjTQrDUeQLyuXQV7rzGdNniUu6QubsaA5uwiAvDTefkFuL2etJy1VSywHiD
Q6BaA+2qF9R0kJHHTlzgMolK6R2EgXhMFNmXnsHaPo0ks2WuWhqZt2TYs6Ghim66
5gPfG3KLBcdpbMQrGCSo6j8magP0Y9InEwEQLpKaCRLeUbyiblJycPznLP2jO+di
BKnIihRAXUawSfFEeZhifgY2RrngPyca6s9C1fIWpI5tZel7aWjW4SUiuyZxL+ls
f2dlzVb8rNyfosGF3bF6lXe8xTyaQgOOb8LPoWwOgw2IzWDSMfiWB4hVC8m3Vw5y
XQGbkzVFehhZ2zecThnfgM57Zwf3A0Fkk2PhwhDYlR1OHAZnfkUSHa1DR6WWW1Fm
f77TYsokcbo5enSBFOCd4XSM6VFZCVWLOpg1zNi8oxCH7WwPQbh8xmkvwvPYsANm
5c5RrP+lt/b5DCfwIJIOPtjHA+pGo20rspTd785/TdymGKxRS8/swqtBgICszi37
ypJnJtYwcoXjqDpnVT+KyPHxTowCzJdTJMoHP436dPzRzFccvtlcAYffCnlvQ1Ia
yrkG+jC5v7PTCZaRnG+Dp2V/2OY61qIYgmJXqGHyVKYRy8/8tXqchfIW93I4NSCM
ZU501AB7vPloDHsx9ToRePaIbfqk9fxsfP55fcKVshKPJeIhLt/zcluJzQck6eLV
1EQFzr1CBmVg8a4PFyEr3y1W/VUDYL+b9uxF5zbtPTXywZxj90AQ9aQ2GHWpsLXd
RV2wCbJB4WzUBoHlGYyiDhsHUUr5K5WOpgl097XpeXnJv0kfc7+6sMEYKSKDZmrw
h49p825nmNbQtsxWGh7upMXrruJbUSVqHN9O8mY/b+Xt7Ew5FboMZrE92HScPF9N
8Ib0kolfSvLhoqylZscou8M/ij0N+PmgDQtcT9nonPQT4u4Dfz2IxUUGBRUrQTjY
rZnYbeFEeJML5+kNIbeo9qFOicV8UPtQWEhSGXT06Yq7MEG+TfI5K1iFA4WMXRXm
7h6P4fQkWEC1xC2uS+x+I464NoeQHQnAIJTZ8dU39oSpsK2AP7OpiuuDBgI6jeJh
1uHUaA4szNb02Gl+hh1qek8rfewV8nLUTHueWh9Zv5WMmU520QBPj2NNoh3cJ2U2
A2rwyuE43E0imct26a+jQYAejAWfHCp9gNVoCt8RxbHJ259NrIke1OMKcAiWy4zu
+w/WjTFYsMKBN44GkpPaaQOuwwhShwSZweZ/n54LzO5tO96LK884FjaB84yxiXnU
v2AE9eWt7b5/wDFGuJyNaNt6xm0DExm3t92QbElG4kPLNpFs1wY3qnr5wVjrcmIr
F9kSIKPJAoHdjhdvc56RhVfutKdaCbdjiZ6urJGAXi90F6GQbn/BnYfCCle/x3qz
/j1Eo+NmEG9VKHbmx92mzBGs9gQhnSXTVKmhw+rrAqv8wEWEz3NP/2+ZgZGXt3Cl
syb4Ay2qtJY6jXdkrWkriCFeSf5y4Upd9FagZuA0hKjWAnhzL9cee/H6RV/yI1w2
L1zb7EJJafTa5PE5ivNJA4BCmsEbvlrIXtAOXQcFK4maqMQsKOcljKSIgExwgXLP
3vVj9KnvoOZI0aA9IG5qrTJOKLwsKr2PCgNZdGEbdybnb0j4Jx2T4DYmRH38wLKz
fdxQ3Fu3b1YhvHcq5UOlIx5BXkzbsrhsleOYZj/HA8xp9HAAClb62yrXEdRwER1r
ASpHKG9g5vu//s9Wml/N0KoX7zwtAxae4MAGrDT4dyJfzdz2ZaIRt6/vg4bssFlI
HNMZLymFfd0oBlbs40GIh3y9DAKCmYMLLmlHLVuDxwv+0a+XhQkdXkvUMv33m688
9t/o/T3JdGWGyaydV2Ar6jF5ggZrxa3lkpRQrV3o+a7c4nWMK64Iu8f3VAh8uC0t
TYfC2936ytBJeHVXWaGt/GY8w7BD67066tzmeM/nV2hKh5erdxh3WYSU78338tgF
nimD1nxpx+13QGU1l4W2QPCyCnsVctWpFUOpf7Z/34iwllCr2MuwskkA9xbsoE/F
DtbyaxYatcQcmuQi0Kz7YbOjSaiIPLxdFkyBaPLnzH+wUV4SloqpldXBWZ1jk4al
XtBX+Gxh0EMCrl/MJnQWMAlAnJ/XFQ4vZQd77EE7xjPz6Z9O4puGtkQXOeZgpmPc
1nsDT2Y/DheWhwGhGacIeWcaG8PWdMhq8ITw5buLa8z6ZwQMaobVZf/mr0Ds43pb
QPDAP8jcVJucTUrEE1yXvyhmLf+E7CTQ5fGP3/HrouLhpHHY3rdVaAImjkn4Ycvo
aKlQud2PJCbii9Z/ZZ+OkG3aVixXnx77ScA+IQZqBK9TcMHy4ORausZ/K40s8pBS
cNx+JKLDZmGaTmc8lus5RMtvp1gZH8aroq79xcAopLh11fH+7PndsE1xGvuJSw7L
E8tTVasdDBtVdKAd5NHRqTHYFZaW2lR/UPLoQjXAUICEWGv3mO4wpmuGnlM33IfS
mZWP67QolPGK2HBveueo6YehyPKcjyIgv520NLorrkmY7M1DA283e2BOw6QR+pcA
5n62JbrWSEhvrYdMGipsLM5/nBsImXzC3SAy7q3C3iTlvghi9qe2BynwGAIU5Vud
9WNmSdBG9oZ82GzSOhxPcxayS0P4EMHMaYoT9JANXShUs5yvIApdKTISfpqDQbgD
TCQYKSSkBqSDHqh+fLsw3UH/eZ37DRhx+Hz6P3FWrxOA5+Mq7g+LBY9uFAK33Lih
7NRaE7JE8noGFYnaj9+GB/wi061QYub4fYx5SgCEXVkRW/KNJI6Vt4GPJu7kgtRO
3O753fz7DnXQsvOH3RwOS74I06qjFiNFHDS6x7Cjw3yXQl9qdyHjMkNkDvjy2BqV
8ozkC6PvxPBjA93lDMkIUxUlSB2HJvSvZYX7hbsUI7/NzUdp/J6mJ5TJbnmHRMfK
+YBl+6PkwSfAbMPPApOsLc0RRH48ETxuW49Qi5dM/REmBCTNJBtEoScAPPRea71H
mD0d1NnicV9Bsq/A42ZAyfdjV/bct5aLVb/HFU/g2XTfis9OT4QIm9Y/Gd3IAV3K
Cgnrgfbkk3pT8togYDOySt6Y5vJAFT4TXyFwyPWXBXSCNi6m+FaBistf+TCUH6dI
BZuZdOy+4qvibzO4V/E54icIlZ7GKtstSv6P6s1SuYAC7sI9N8pnnVU3V6vDywDQ
PdzvUAznLl1vtLfL6Ni/33onrlai9G4Dhy6rTIoFv/7cWmavpcafzcSp/ZbzCrCW
++cpXBDrZo/Lwveuc+BbCk7pmYVfngPL3hGpcMY/ZMMLs63zl9nKXCtvEbU1Kebv
lop4QpuDP+3r1MBUid/7z1K1NAn7vXruCoXFPXDlZDvXTS6R8naMLjjoT3RezzEh
iivTZylxxhke5R+/XOnMt6s5/qKezpOBvdKLnDGXDfs/z3ebuwOy3qlpaew7q24A
EGdDekgxfQqjDOZi8YZ7/c4r4kUbVvloBBkufv0yM3/QIxTh/bIs3bdLeAlY9K6d
mOIsxMNbpPrr193+WympWcOs+gVrWIyh+0LdDrUt67yIiazYgLGVc+eFMZc6SWpZ
U0gqC3ZSgBmCCJZhNHS9x4VriSXBYJUZL37nR4QIBw/jqTf5lcinXzcEQqhpd+/7
Ae9Jvx99TewOUhPUmG6RNU+Rr8tGOvWBqP7mmWPO+dt3SVpnp36XKuigyk7Axd/B
nhnW8Oi/0yVF6cqWFqZtM5dQj4NCv6rB7GSXuyQil6x2RL6TRFKB+O0pDcWOfMWW
pJqrVXmByo6R1V/YJqUy9QycMUYhUfq6SvkUXtxeCmKla/vXh73oaKOAUWPLH2H0
Lnu8ul6ytI5s3Wed7tUKmS6zkM04ZSI3zyghOQ8PquVIrQVyVipUzWu2i1whqFQx
/gMbwNFBJ+qZ50uIN8tQlT/mZMrXNp9iMUUNPUR7VwcNVFWNTFquetN4Dac3XJt2
prTlxkDtpLcPxNiOl/lDdLL3dFQEaMU7eOkLpQQ7iWaMAKIS+dfsDZ7w7l8YFJbU
S/jfhBNEkRGhMXLMObh91HB1crnnGwL9G5fklRInc6ZCMBq+qsVjiBQw3Aji2nQE
0VwzRQeFlpoF0TSgHHjxZvplaQLZV2+x4StswmgbVLD7ppDtl0XuKCA2nvsc0Lvf
yw6JFZRCOSTVcVqGydP5u53NPTwo60hOIPLgJulY2NA0Irdqu7f7r66rRz+qcRaD
53Q7KjdcGPDukG0EKUDaB7W3CrDoU9HoAWBJeGs+hfUjvd9dSi/waCz5i9ZMUdNr
FJNA99qg7q2ipoYanC7DZU7p3fxDxNBUe5vEOngKvaoqNlfDmJezl/6dq9c6+qmd
empab9rT14KKBpNZwtdYnmo7ZJwBKl3dPpVz5GJPLlL53DwgGWv9jkkrPMd07CQY
N8U6rRQTYTJOTs7D8jes19B7iO7G9pnxNC+7IQLONxnsg9zD20Gztf0S9cvI9Isi
rfWTkeOx+YAmJr3wQS/FZ50OTpEgFTV7FqdWqrWX1I3gQGTRMzYgG7T5clG1HJWp
JguFZk6Cn1wWnMfxOoZY+uguAShW/EX9AOhKHfkuFAPk/dBEdj4uGr1IGx0z8NtO
siDmC0nXhc4c1CPazlWdvxZ0IGQ+ElV0IgOYwgPsYSJjXXC2gicOKDi94raGtm9A
WRl0wJCU7XsX7tMeVrVoOezJ0j/Suom8tvli+uiFgLqH4TiCsSB06emb+8s5PSek
f41Oe4Dxodv2jkSiqfLzZRzyiPqAYVvL7YSyR2ffx9TJMIN+u24rocWDBCj/kE0I
T7oHj1jVX9GPKbAln6PKYsLuOpEwty29YyvPhAlGEyoecVEXbLwHk7Y9Dpm/sIgP
2nHLEzQu2ANZVD8xjnFtJHpx3GhDo75iYNIM8FisqiajiK5vah5auIw5wH5V1pL8
ohxCzgGlVnnXhctfkiV1QKyFo0p2cHecHiMGNWoeluJU74jWUp7BFDKhdhTXbchg
fhrNBSof7EEIjJ267XPyQmQHSxI6J8Br+DNZiNbtKyCy5efQBPPseJez541K3sKV
xShjTr9k7cyHj0lOt4LDsuPYa/nR8SKyewm+3LkJqjE7RiNvy81QPXKSSotn+Tki
jAp6QK5NpJsgSlO8N+xyQsc8qkqvYwo6YyvUUlXjRHrmH86CxrhVG1NIeel6Hb9q
pKmA8ItGl1lJpjl+C1GsLJNf7pB1lRvCLOz5+ipX2RzMBvTQcTMyMtWr973WqrBH
0mwRa1nj6OZvFkMi0M6ZtT8l0ySFLYxGRBW5efu6rdK0XgQNHCZGzwDPgT0ydX9S
+5OmfI1XWt+rrYlYsM+ZCWVzArnY8VPQHsg0L9BnqcewdXKO70UT68VKKrCeAkE/
CE67xTJjlYVJ5gkBb2GoCagYEwE6wp+BDm9P/lMlc8GIQwJIO++lelbVXUuWOHbm
oxw0ukLr4N4KhsHHzgpafniRt2FSQqB5NK6/g1NhE4j+sGeSK9IWuWcohrgtGJyh
q832UttEeo//QPhLgG2IpeQ9PemMVrROi33vexAwZKllEAbpqolmhU33HoJbwe2T
XTMyGo7XxFA5Zri9UT8anvzDVClUw7glxkfzoy8KYZk96zMWJnMH/71O62nLyF6E
xS/yVfec01NjWOtcGHnB/cJNH76Hpn7UQUYND9xLnPvBsBb0jJtPEG8kLavUPFof
seSCCpqSv/AXPCV9w3nb1yri8uFoi7CBIOB6zdEx+6kJEzcSQK0iG1shYkuBPkM4
M7ZWeQRJTw+SHWSFD2MSmE98wgMRy2nyVfZJReijBzWCIgXxZjn6DnN2IEC+npYI
g8fgsWPw6R5vNcnWW1U+w5yYSMEg1RnkedPZSMmoefFln86BhwOF1vKfhiNztd7Y
TJVkYuLzInJqU2MyI8+o/E2X5tg4KXsXFutAsM8TIP4U3A3yaqtyiZDd8BJccupp
nV4KtSfjvla5N4XMh5PZntUcghn+wIf+KZtCmdeOHYs6dSmOLKqMPJONvqgHAC8V
1BfD1J72LYeR1F1+rY/f6zL1pIpQIbiL3jX/z5V799ZYM4blJvqjMMmsPXEUKogR
7olMlWrEvlzW2QPizKkQsVnElmgEAq5azXUXlT2Jl5ChEuhsXoir9S/IJenBR2Jr
sID0ylc1E+qAEbONHY3935GmJ/8gQzem7WgggwJ2smIV2A7RbaaQ2EOS0FraV1Dp
Sh8gJiBxlyoCX3lSY0GCmfM6AZXsjppE75jYcZMJgWq6/u6osWxQulUu1ZPZzMAM
dzteaxQCGfQI1QCKXyRWESdRd0wq36yDBntIbeITraTmGhQdHpf/S5VQ1TellLcs
RJYu3YZKMt/rxhIyOqZSR/x7aH5QPsjGcD84jYhXPaRcIaV7qb3cXZgJvLVZksh8
c4UXZB8q0EqQflpWtfm0FNxDFAuqxvwCJfNEjoIkvf9dgnyWoqCAOpJP4Sb+So38
iJX3FxZTdZRFMszoyoEQCPW62mfZrCNCWoRPKqgLCCVBLEVVQFAHY+FFmOTdJUkg
2JvI8lpsAE5YbalzvTrl0KPJ0H9hlr5sqmROQtJDAPkDH/xVyifHGnVHSLJ/Pt+s
GFFlHZMdM1du8qy4JFgs93Gv4ck9x92lwgEG2sp8Z2+w0v3eHaSlimNhYIltNlRK
dHbCcxnSFE9McLOnAuQSkI/NTKZo7/nmBbN/5BAqt0UxNQM5QruG/Zwu1aRb4Mxy
Ynx9dmGJDto7FZ4loxlKBzecXrYj76r6l6Y7KqwMMLUDgHQpbDUvN5TRsqqOLya/
Qe8RiHEODrkY0YGxSwgaUk1K7j3GaQdm9Cn3QVU1AUem73Bpt8g9vJcJuMkG9f5S
b9EMTSwQ79rtijEh5dSsG9mcKivFtt8J/jgLJhMfa7NS4On1BXUpUWnCZBUYzPNp
GlBoIbQQrhI+xiu/H2Ec1DxYKGnnG63jnXmI7zcYtcwo5hXq+g59ej+iYB/6Vvj6
v9OMHjPQyTB5jfgaRPpKh/aJR9q9/Z7xUdO+QLIW6dwV/gmP7hy9bo0s9QS6mO7d
0Cm3KZp0CFgoMCijIXqn5S88tvWtW8Xbb4cMsHZ+CaCaE/5Ga7UogUyGhERmAJrq
7EEGo0p1tK7Xnkj8+fcxicn3FniG1OXpPcC+wITqno/EfxDILtuUVi/01OvlFXYZ
CaRAgAZIQGUJs2UDMgplz4pSzeF/uk3YjkF3SVb62CfPhsyyaiW/jJS8gGv5Cepd
mL6N8ASTBFLbV6QJMMf6qicri/W/DdBOUUduXXWINss/o4r5h4LKi2T9TcgLV6FD
IvkKEBc5PIcI5OuqpEdshJWdhL3zqi2N49qQBuSXwSFE0l6sW4JUFTkEv5wHdNgU
bMCw2jOmOJmcDKjmEtNgkERPDwgIZxLjLta8TyUCY9BGPlnFXA1GCVzI+AJy4GUl
bTYLHw1D8yfdFQksWIozXlvaRxdDR0XdXqeM/FHL9WBhkRq3/vQClafCh71DsvEx
sJoAa9U/IACNeMAloOwCgBRtHDxNe8Dar4akubWIPhd75y+xvGjB/mIQmuriEtmk
alIEQGEbbvsM/XTS8eKS/bO5EkTQD6zlc6GVgNbtDIWb2lbTaKbv+fmRWj3kDF2a
MOddvd2uziw35Rqac1LfcKJRXF9FO78xicNVSFCFE7aJ3tTggO71RMoFYXvEullA
LUpe9cMVL5hzF6Yh/8rgHrv+BYJnVqhilm72q1H5MhfRjMTVIZPJdIrfwhnAmJNe
uP18s1CwIIBD99P2wXiMXCljsARhJvANhPZybQc+LDAEMYqjmlzodzd6f3A73n+x
K0Qrbfu6XABXeVwWj8DgKIRx4iWRa3xLrsE11pFttitNTwjiIo4E9BGXccm4iQ7l
UipHnkZHsdjBKkOxHozF+jv6c1DNHAHGxEfD+OR8ygyWGA12kiGPkE4nl22wYud+
VDtPQBCdGbK1raKFio7ouB64Y02Zov8rN5bCMBd08nUV2d6HbGLH1JWG8EI6qw2g
ouzOCBBphS5Idc65ES5G2JZE4TMGfBuHUTc8bpJqcottQhN8Qb6CvNkpQiP2i5Ki
wIXxASnbJwZWKt4IiMwC2s19/8dYHTj5zYDI0qQGeP/5rur3intOI4+FFIHpysu8
69xqk4D5ky1T6BnXapcpPdG3LDtREBc99ISRs2jE0DPonQUDYLpVyrk3zDSH4xR7
tVQesRfd4aXXDTHO4IU0wA8Wg38kn4Ny+3hc+ZKzbSknfSmVqOqiKSrN0oxKeNmS
rtycwFk/XedW0FMWU5OWNnIpAvZ78DpUgOIFKo049chGBOfeYCinSZ2yk7FqCy+6
EFFPn3uX4cCCzMshSeXCfCfsSCOOxJm7y5CKAVB3/6P9sLaeGczAAbPa6rAhTM0N
QB7iE9olEVJKTj8sm/GVGryx/D1m93xq/paniAiEq4JFX/BGlRJBuvq7+OvjIGHz
fka4G5QMAVb5QCuAafMlQNa7mYHAYuZLeD2h3GKK0aOSRLO+YC1LjbdArqqvg2qO
kI5fxSgoeIbV8KNjnJB/eoWyLJSpzsuaT40zpQfCyW1DtERgSUKUhXID1wzLyy2M
VminpHX8jGh2uKBYt6N4/6+G59idIE9nBeYnUCEHN54MggBXJd/9d2E+WPrnF9+i
JQU7LxLr8sEkHjPFVU5PVGWw5aDHJ9DYEjv8aEIwl/H7i7S6XfWu1SZTNOCUMmYw
JugFgoPsGtIJ//3WRM9qNyL8l5X86TyF8va1W2paJGlw+U6kn4ydSlheWEK2g881
RRn0vmfKJqFYS6wsr+KcTm0l9liQV6V2YNUKPHYabtvNU+z3yfQurxp08+u6NQ/6
XA3/VSk3pHYD8qWQjlJGEyvpPUqDTy+QgXg+yIL08qGYjQj0Nnl0CBP+eEpGj/pb
v1nR0wTGwAA5nyVIQacarvbwJBgAMqEe7s4rN6cSGaWC62sypa7OI2sCTlXWhbXK
SPz1bMJSAU8tzmezhkxTFHmyczKZi3oF27qteBcASgAPzf3jXAMxxfBZALeqQgRb
OTipAJMEIaJh0c2ZKo32pGABCjKciHSmveCMz/jWdZ3QBmnZx66j8mfcBqdInSDF
pGd/Spcvrihk//hO+ChK+Mol6FWPyKWhckPSFhs9MJOFhZBDGi/yGvg6jnexNwjJ
TPkH2iYE+je3cDouNxgCj7YbvufLU7sqh7pwQ7SqaNRgpzDllC5ZQDhTCYM4fMZK
7lSCbz1a8pCZwKzj1oOCev+qNxP5KnXV39Ih39BKSPlWReYH+uiLI/Y8PBude0yJ
FyJBJuJS5+Hmp4O9TeaglwaD5ZoLY7IMvS5eiTsu57+LsI81bRBp+sJHurt2YzIg
GRFe7M10XO/UyNKN+jySumI9UlDuxd2q4QLlbQziixpuvSUYcDq4YDk7vZ2uQqW3
6LLebwXgVexQ7Kc9zXSdeMkmw+t1EtqvX3onfy0On0ev+qCz9YDL80tOoWRBuJSd
zL2ozyWPa8k1gQTR2ZkpgeJLzLb9VBI2OqjUe95v9nPIx+Mb9GfiY4IZGZM5r4Eu
aj1YLFuEpN3rARUhuRnLINeG+ZqOpl9oCP98gnEuc8UNwVEWLjnbTc4wBy0eCgGr
H2Sb/7Ptfx1Eo1P1so0ZX8uPnbMX4GJQk0hTtpGFIGmh5NkbJonDZUHD8OAseyfD
+DwRy3bxx+yoNyaru90agIvvOEkHA7IeJc7eAPtx987WmHvnqVPM+IcXTup2ZVXZ
JV3Mlk47wn0Nf0WEkebMuhvs8NEMm9BAvCHx40kAot30ZeHf0HSVk27G6waekKbk
eEHVyMCLUXKs0lrWONyzxniMZR1aGCjkNRGsFLF/tuQ3k5aP41tCktZv+OG3FEqX
o0hoZ+6+C4lOyK5vZYaapeFqvg/QmOzuds9+I/uhN2LGl3MXfa1adr1BO73ptetL
ocZEq8QrKk1fU6ORq4DK89yfNUFwYtqO+YKtW9t4XrdLTS8dE0j3+gOZvin06kie
vFb/gaz2LRmks+HmSc2MgvdOKqq69oF00z5PMDJ1EHiMkU1nG5zWL4LNQv4qBe1X
RoTIQM9JEGr1z828cCQLW3Z9WcTSREj1kiBXtvEqPp9/u9KXVZBnA9nXcF+m5fFy
gKNFpoWPMQkuApXtsK/FKqdfue2AfJDLquQxzE88V2tl2btW9mrGK+avv9yN8mQh
C6rGO9oZFPGUiZbrA1dGlxXgf2p5V1DzR/hAV2huJuCCrB0vGmZ+Y5S6epT1q7Bi
p8zlelumN6htIFgBtNTJJ/t5FotgSrIxY4iDi8+VVILtEYK6grx+GWEH7Cmqpk8d
/b4NcZoWxJjh4MbDu9417qwMiMUC3LvyyTeVwliimbs5E60aRhvUYiDM44uyXN4R
81JYijgtxGmpnw0j907TkhA2G70wbxRrQEtB0TRGOd3JWZg6FHEsSt1CXssZaPQa
nsuITN0dOs/kVvuFHZP4IKm1a41ZJi1/QklxT4aUL+AyVigUZeQ1vbe/hoL+whQp
3FI/7V0INtvPsxmtplB1Gu5FbLGdvV/oKHkbnu1YScj+7kqkxGfynu4e8Ytj5GmB
AyvXlP4TAaIt+dNOZacGPOrHL7qsqYx6eVvzWykmjNs/0DKjzaITcJIez9cSm1mB
hTUHdgqFUTAa6O2Yho8kMpbE5GYQQs9RCY5dbO1Q6kL9LjUXM9lEqAGaipfGYY2f
9LEi6yk5yWFzwvP8+bDmsKZ1Q75aBpimbnYYaD9RA5XV5QLR5nFCnMsFOTZXe6NO
9uo66oMPD30lKpLXCcqwjKVzOJSMFp6Y4OBp8/1pnve/YVT3T+WUyEala25MiCbE
sCcV3zA6qExtkE5hB1iEfJDA45MrcXPaaMzkJYwdS3qNoZknGz4y9kaYDtBhHXDS
NXLfKtktqwwsm+amTPs+QxWw1gh18O3FD1dcXtZhTMPioQfnRkk+uYQrQOwZ+vI/
2xe9TwIkKeZAa3DbL1cB9gkls0nd284GU7UusC80sDiON7G7j7snoFOh3OSRyD7w
kAtpCsUx2Fl8MImG9z26IrhEPqrgT382JV+6RsaPeBFSg9WKBdUcHrefKP3+A/GI
o/kKokDk+0cUNbS7W6WgMQXHXQx8PFgPD9dWwbdZwm4L2O3zree8na/Vv15gqvs9
61vgfXo3j6wzyf1otWucgRW5k/U/6sZeN02digi5Zm0dJsWxlDEwgfA2pX6luEvM
13OJI/OtBsIV67PpWaeZOEsPgNinpcwliM0T4sjBsPOfbyAkvoroeiLAagzN8Hj9
gGoq/YPOciLK0j+eqRrVTLjarawHQWl7+qxmJEmJo0mhl+fKLGd4tZpkBzL8xN5t
TOVejtQNiLR2Doz7SasMkYV2Oe+QYdvKKocbzlYWGeM5uW26QXDN4ywwsPjdNyG/
lI4fvWCOD9DhX4wN/pa667tYuO8qlTkiptCLajftdEs1C9ZhpEceQCWYrf8gZa4a
trshBu0+0iZg3NXHkOsPViV6yNx2NghohILpPlCQXRVwsKUYvaR6aeKzkXY3mBSG
s7QdghVQVNp9tCshzML6LCKrKJ85n0dlynLxHepM8Nwowy/2OVyTm3UM2lecT9hV
ZkauxQcokcPbcYGfJ8FpwfSnMudruafZ7Tp5i4nGqI6V9+HQmnfHgqQMdPPSi58A
h/U0agXES7Vlz6nzXi5TTVO2ZJOEc566xtHyujBwokJ742M82PpW72n4eBtDIjFy
9hfjFg6Yarkz5k5TcAulbXS/evJGwjEcablyZF02+3blxUbJ2EQXzAUbU4PigcFV
loZCYRstry9JM4yu/N5ULIwPl6xaFpWIpZ4Mg1cOHF4IChuRH/mW4wnsvjgRX2CS
PV2XB4gsc04Mk7KSf36xue2jU2i0XRynsyyv58IQbqYQsb+Ugy4CeZeErbb2wm8y
SR2Nzy4OG55pumlvz9464CGwibPKYlf7CSp3V1oqzmVEyouaQFPe9lpgIJyp14mI
Xbom5R/R9iQxUd5jWQciWG9iAklSy+Jt/djvljZYfrmx760JL7p3Ogfj3qAO/c5P
0hE9+LO9BjESN3i9Mtn8npyDV5X3eTpmO6Rh2Htl7D+66YiAJI/o09jlTT82Nxzq
N/+wJjmshA06QB2dcj3KdFFU/yFxRw6L/9mItvgoneglR6v1upoUGFFeigtFL3Y6
KMnY7N0m0a6FrcXM3cVbMhRHzT/DJ8J9n8qBDxWIcyrr1WYMgQzzw3cYdDeiCFZ7
jXQrbJEEHS1vXRG1Z2LU3GupLRF09QLWtdCKfdfCCACaFG/IbmLRE6BM/Map2HSA
Era4R5Y++n/JcNzPiCYclcVoOjMJFFIRA7g/Wfh6eVe4M8Jv/Rc4l1j203lz7RHf
tHIu6kKiNQQC3xKz5q+R21ZSb3s33gq3dG47RMmR+QtAVed/rOeoQaUgmBQgs1jl
yDlAGb1+1i1daCzxw6QhnjTdP7mz6S4sDziNpV5uFUze2sd90URXzeooKQlhdRUw
gghMR/fvBoWKZe1cVCFDMR/1oE7wpWTqE9+usK3NRGjHs8EM/IXsnqMbt30Z9LL6
NvF+Ix5hdxzZBKAPha2LOqU4ds/xFkH/fDCd8ZjoVYW1Z/NWJOK+/75+OTHNqgxI
ykPgN+WO8tHw7doyGYpkTwwajLyIbhCqaugwR1AzSr81VS3OejVVNWvJBQj3v3je
DvquIioHIUGKT6nPXbNKp47K1ETq8YqXGA9ZUL5Q7gmSTuaKEzvVBML51gLx1xdA
6A9oCZjHhcFDywGueUhipmj6iTK+GOVxEFHpH9ZsougNPc53AWkoxNS7+1CL745n
DWRNy3nqhbCiEu+4q0F45FBXAG2PiorXxt82t0xGMah3Uknkd9T45KmbplPhxDsv
u8QQO0Ik1wQlvwGQhWpevvB3Pi6XpvXlTG924aZ0vNsd+jOt9eDh/9FnVh+orAOL
QiU9PVWwGv5MeBa1uu53ZIs/9mLEQAkyFU1E2BD+D1leQ2pt5fDB58rHQMjarbI+
o/8mWSjbsWd336pV37YXV2pHuVXjyBPLgVH/RAxfbH+RNjaWX3fVK1kVXHqXEObu
G2vp4pOaGtTNrFglT7w9yzQaP1lEHAmpodP6ahfXDQLmSXwk/H2EpICWBAwRJNR2
GdYodH/BNFlFiWoy+249gr4nMYGEx/TbBWdWnPBQBOGPMkBAVu8nVBNjkrD6NZxG
60uys/fJiOUIb3Ro3oa+kMr8VqA09IwOCFnzqA7NAvudOVGOieYuL+jmQjEYgKA9
xtsINbXdfMr80So+nmCWlDAmaP2lcQ0+lSJXGeg25TFvmK4snJuq4QR2+Sb/d5Mr
QlgG2ZWlI2lv1nYkLiRDA0MH/Zp6t6MQTTb1zsrB7Wu0NjD6JQVflERcXkA+/jEW
DJztYrYtnT3eZuCNpDS3zSAq4DreqXl4dnMsLZ5dmICHYeH/TZ2RxkmUEKyjCGsg
eETg9HfRG9rs/oZVu5fJ/gBr0rI/fyJ0g2ySfawmdr1qdSQJe4PJf2X3KIE2FQRD
88obigxVtwrvxvgJsrVxea/r6CuJ/dC3RQ9NiPIu8GcGfxQuu3Q547ZAqUAnKZaH
btqTksYoQ6SPC0lhML7ugoxKUP50kkuIqjmCVXJdOUtGj91bCXiQhWX38pyxL55s
ZR3FeU6w/+E1W27sQLhT8OUbDAYqGFWcSp7lrx66KL5Jix06WTIGQaA/AE7cfxaI
l0hlx6H34AIRV72FjNQbN0qNXpNFoXqLLssK/5+L1u+kqbgNBZ9m1t9Qc60T87bh
btEwLvag5kMyVYdWqwb95/IlEFC0MYSJnXQfS5l7dNA2XtrPnt9wmJrhygU2RvvI
qi88df02cdzM2fNt0DjV9sTH/1sl6mWa7GlMvHrzcAWhRz4hxq4G7/sdi6nEvoBt
hkwsJMg6eZIXZZVAGUe75jbQrM9jy6cJRQQYjAcGlnT7hDmcOfeV09CRl2Thsj4Y
mi2wD3WKFQY2JiQDeeYsvwlZtG+8nm1iYcfq3rp7qC4JVaNlUIumUHa1f5Zyq4mg
K0EL/qA4tV9enRI1lnuN2WdpMKPB/j9MKJ0LPzGfXuq3VCBt+OZ1CIyYglxhydGR
nCeVW/zxYibh7jmYPJg6Xes3rXDhrqbWzCaXQ3f0+f+W7fNumEB+cdnPX5oGAy54
nlGL38ruKBZfTyehRTXcHJVmFhLeLAhsHi7tp+3BILUpe6QKn4wg4fgjvzfhVojo
8Oz2j1iecJB1xkhob5rK6gXoh/15QhPzo48nfvGYWegsCQgzrRE6pN8jsTyopIgZ
X9uFCjv3+bNb2pFtdTYlKSRuQiZ8M4HZDWWqgP06R5nPrGuatiVG8FCJBxdT4Xwz
VZw41IvSnE7z8XO184yAHYmPkN1t3i1dTEFu2+eHhRoW7kjEF0l3hMxOgrkpW4eD
/f6MMHoSMEjxx68SdseF/gXFMQqA8evuoYpHGveTYT3tmo3tVJJY6ZQycPktm4EY
2U/v9jqjYj1+F5MrHaIvbEeBWRHoywBV5UTuX8wHUqzZuuhhatiRJPMNe25wRP/A
EMlTsS44VbJz+z62kx/jPHgMNbPoz05zCTADHtll4bT4g9egl+OzPoHbIei7xHtp
6zsep2+5PXFcuycqk6jOez/5Ygklhlgb8AYiW7xJgswVWf/CazYrpVzDb+ffTsB2
vRk1rHG9Oeh96QW0CYtDkZ7pv6MiQJP6Vrzw/ELb99QjP3jkWyYuj+OfXabiFKCt
Ga+JjYnUAPlFTKoClrmg6X75+dXU+2J9P3fb4RxY8iCVq/mUL4tfZasmAWrhBrId
XF+TLiHrjUOM7Lpj8aKGLM1Ii60ysWnnXTvg1unAJjWpWtVpZHutZ3VyfNMOrFqP
FuVqv4HayJKTEYpkU8yg+lO54rYwbRJ5bb+DUqMF02hvii71iciu8iaRAD9eOMpX
3RL1Kv3x4FoN3jQiS9YSyvRP0DB21i2Na6xbrKlafP1+YH8owd/1KDidVHwhZQq6
5JEolBXPbOId2nMzOv+V2DbGbehElGGr2NjBe8MypRVJKb90LbHgYbu4cK1SqUwR
DKLHjgAKuWC66ZLlAiFVSBArHtTUbwjeuLEuB1ZOH4uAQpKX+gA/TnPziHbnVQOF
H8ib0xST6xZKrboZaiuAgW60T6P4GKhq4yuIVkZxV5ww/wjKW44pm1zZ12VEPCV4
kbX8SsO4F1e2L3rbc+F9lcJQsqEJ+c7F0NGJ6aiAhmR79mAKWwo7sdxOlkLFsboA
KC/wZ0qm92xjx3Gu5PVbeS9Wq3FR3kEBxnKzef5/+mRUaV66ZPjjrrD/udYofFXg
KMGZwKL5RhuKvX+La8uU0+UVbeOTMu38cJuVfxsI71ANpcMrFJ91xDPVde1bR3Fb
MH2Od38NNiH5O5/t+bMh0Sru9d6bUnuaPkd3Qc+3NAn50taWtSj7o3fojaiGLGFz
ZRDvzksEqKOFMifLzbGuLuItR4FSjPGsQDReyN7NgQW/5TRvOxWlfbAb+PWBGWsT
9h+KM4InByXx9DA7QMl+CKQSCDEC3ZKc2k3q3tzkp8oiPnff7aBO8FoOYMpih80s
sdX2PS+fU3t2/rSecQhXLWzKQVFyAUuk7dgofH+sfz11HD9Eyq+9/v2J4n666y9Q
QjW+LVS8rKo2SJYBZSp4ZT3b9hN6ZomItYF2cgns5Q3ATUodI+685PVKMNcRpH4x
wpmWF5RC8ISMml21rtIowNV3CXO0RhW7Yl1KEp1o5+NUSmBQRu7rx50ZxYUqKe54
Pj+Nn7cCvwKErFjFohA2GetYuQppCJEGZCe9VUZjhTLgXF2USODkc+YCSdavhFZf
zMYnEZsjKY2TK3JKCjBvzJVcmOhpOgWhcPQ7z4vz+MsukJTvootWfnZN8x573Adl
XBzb6ufB2PxFMgSk+bj48FzO0s3LF/Hw2tsr0Plew3wk0XRW8+EM7OvuBmc8bG+P
IiNl0tfwu/cPRgpUF3NE9xKOiinA2lIcU+4qaV7Ii4a4fiq6vPkbsO6afxGAvAEF
1KXRzq81QQYQ6b4X9P7qaW5ugpKbJ9zZLhvnbXl+UzbTTcOtOmEJUuMyjeSAhi5C
ngQsLWUHbndR6OBfoUcrtKqNCc+1J20VcQdGMe11DoPH9nCvOkiskos8JAe1ua4K
cFy8xGLUathN8PsLvQ9jbdGLwt2XRX4rpqB36mY8EpwNEUeqR16OMJ1tBtMgAUnp
wYf/3jZYbTgi+abRdmEupTwjRL3ipiWT3t8P8ZuJGl5Xf5REZ8slsuUwfXuTc/LR
t67r5ICnSr6DV7YzQmYy3BtWbLSamLQaP4GIGmWzA51cjBrUdpGtNCNRGh4Wq2mC
cRLP76kzidxN6VkpU7saMqXyijeA8/EoBQeaHcKC9gKAg+M2OxY6/G2ToQ55QS9c
P5soKXC0Xe71C2JZRrKc/2Yr5v28hhZHJJaqoxKca7qg9yVVC/fgJ+KDl6pk/NpZ
2uLStDtOSy6qTkKFciDPvez+fhZmtXr6VxxHru3+aDTvNWG/ZPYvZJGeCDmAwgsM
edbFWW6UeShXh6CoCr7RufVG+6qVD3Fmvsi1+LfLErntkC1ua+BiLI/UQyhJpKxs
Fbhyx/1u2D3GHbAemkNR/FjFLmxYmX38XKHRsv7mGBDVd+6d+f5QqdSVLZiDu7pH
JpBMFYcoWQRpDH8C2LNfTGvIHsNxz0MRAIrVv+pSZK02j5Htd6UF+vIX409EeB9Q
TtiVGqaoefsydmvIDuKdSMdA/31H041tDABo+leaSknKqaacLIn3be5VSdUy58YN
xWJUIbs30pLSRmp2Z01A802/Lq83SJKTmaIB+eUNPECt8yhZJ4XRwbuwNGPFP/+9
BTQkX5rdxuCllr6Y8R1ybDvl/6PazPPOtG/Bi8uNZXTWiP8yTLBOxHNwDeVzoiqQ
1UDjBsixarhvf7cRCDp5LwpZpkeqwl3liCSUcqK0X4OC4USYOSKT/YY01B8B2D9I
BgJAZm2R12ZKvwPmf4GJ2iUoM/8w6FEbuxsDlBig05L1KKnzuEza9fRGevYPNJe3
arxjR0CNbZB/YH1/0t31WcNy+Wlwi6/R45f2A6Zawficg3vIOMccAStFVYlila2n
94P4PKqTZBCB0tfFxSfYtPDHEogtNJm8tm2C1A0zRqwU/L7JtfJza+apMhnW8MDw
79FQ/OIXLc/HhtLq2u3LaAwVIgnSuPjBaoPunK/VA8ESYrq6uODk680v4OPhlKqO
wMBBAZoeFvWtL4r/nHGXWQ9BGOENVFtPnxMoOdLu7o0k8e1H16RKVyv/CAWdGTay
DAV5arKL5+AqMVot+TxQOQCzm/r5Ru5LcBkpxP7nhXG+xAI1msvAn9atApSg7iP7
1YKf147+XuqmIUnn3TbJjqEbogPG8LYdqa4VSc3GYSeXW3sxk8ylMHxhFh5UhDbR
6FZNTX8IMXfDgDK+hHROPsbKXtGl120XIzVWqsQxvBPGmYg60Nv6rlK0ZaiT+BQt
rMImWzQiDmnG38M4pC2ekZKfj26Ko9K5zsFmCM50EN7GUMtoXQ0/bqajshNyEV2Q
nHuTsznOz48jorwv+DhVOtBBlTYxJHj4/xGsMAiPYX3rHjMzPRdzfc0X+7GKYqRP
J/k7NeC0xs89fWDs7aCJ+FkYshmKxFjc3KNFzciwQ47yHsI+U00nkp4oCnpvRWW5
8L/G4vee/SRKiMDHCgjza27fBYeiXhBlPoWiK8NdEMK8FygCnW7yEP9h0NjpcWEY
gNWROtDH17ZbC3QDRo1OBfaiYW5Vw+AZ7lfr7Fl+eNnCql+N1cwZH21qaZ5kz2rp
0mxP52bzooUcHb4sa/hOUm6+fPDXd1rMhKzTQNeCv0EMTARNCC5hZWAVfggi5J1C
ab2ewZzIRv1lDtnNuGs3/A6LbjH1T3hFbKBPWvG9TX4XA0PQdAXc0HtTfuxHOOyC
6E5KtLWVmo+FMoypHyUIA58T3UFkQnXzSEr/TmbHLkj7GFBaleRCHnoPLtzsSg9a
N2ykGsI/zQkuEWaYymdyqpoBnd0amL44mJj/cbeFpZiwcyfs+yzt6lC36a/GMON1
M5kCSnPrbF4Pu7ulre+9mKWer3ng9zBXREZjlze/f6MBUtD7wErWxogqXsDKVts3
pkPMuJZPAzobUCP2iLeIRm/8ootG79seJ5aPhRtL+7QLfQHcgSUaPmVCJyRQo/Oq
/eykcz1pQ91n5e3nfL+6Z/3ioX4l1ELmwJl9Hya//vtSp+IFe2M0Cdj25NiulnSR
RYdIANdgTcOO24cBPhfibkv8FwNQdKXbX11iwNxPAYDqjb5CZpKR5M5u6uTiFQLU
nl3fT16ezQ9c9+PFYObCHIM3+OigFZap0/r+Q1/yfo6FlJJrmeiJK0hVgp+jfLZ3
IJad2jTDRRoJUKm2jJ3C1Z6p+PLZkh08zkGGX/6wTPZSfp0mkyf0OGSJxRmiJXPU
Piy3+cZ8q/pqcqAvGtSbXZm6tS8z2TEjDQNjk4qGwffTvHgjzkQgELIUZH17ZUOr
dj8cJ8EKhsRDaZ+sq0SEMNxggGJJur/4r+IQds9ZrPvjcnAM2T5Q8LdrOTX7CoWt
mE77Hbu6cTv/e8y9pT2wGWlDIW0CL3bnjlw5TkIp7q4LPuMJ3S+FRYdscUS9QFXk
r88cHmWhEAh1U5syJftdZeb9i68hqYsthe6BvwuMuelsVb5jREzXSA3todHs0wTf
68vLybhEUCoad3NcZDyblRWfbq335flL7epDrIxCZiSk6+oWCdbDE2LxPRP99nJy
3nzF6cUh348R7rEcTWHFdFkC8yK+pNm50kwC7ciWKII8L7LgHPfkmgYlXt+IeWRT
pi3wsSrlHYfXr6RGOGb5tj01P0rK0tVgGZ112bntIZjSBUe4sA4B54s+5W+e722F
gPwPdn6Mc1hcLWk2INtx2TmLg8bfrhdK71KdCz/FgdEdy/DN6GEZKTf+8rKhFqlR
KrI62xS0hP2TJtH2kW+mZC/Hu8lhFhsM1q/PdTqtWd2EzIXR9iDp6qb8O+jE1Vzw
PBmrgnJO1zxybsJqFdzzlpUKSiZUSMCGgdzn9+JU9hco6yw9AbHCy2ZIHpl08V6l
MIsfFzC7s3P+k2ZKYGFPQQyu8aYoC7+mQ+FZ8Zajp+8iemD7n3WLsfCYl1v0GAmn
JQSi8AlpsbGHfduanhD/g0LgSmbWLvfhDC3U8ln5e6hVnexaZ7pYlP73RET7ZvnW
CeSdTD4uHKf9omrf7Vt0o4QJMZxA09bZtGUaj2EKTByh4Zd9mLUYd/uYSUvmQ2LX
KUi+mIvnkSuyh8d7tyI5XwivKBmduuVFPw476pvTe7MScpWvaUKnwH5tLtya4Y4N
fjG0IdfXcpnpiv1xPq+kAzqu/c8750Nu1E/yaoHtPCRiTHEhKwSMtDOWCMXtEVka
Z4+r4Z0wZSZQDU4b3JY0e2zsNSq6tE0YqQ1T3/qfbk39xryg8VPupRtw0vA5COgT
0YP+G6VbvQO+E63jmDShMbwg71qfydVuoUFjeNd1ZyDUz4h6v3fncyM+NxM00Ae/
hvhg3ctgzSWUCcCwRSchXC+gkHcDCy1IGeWzSeD8CCtAqj1D5G0tuoxrJTiQNKl+
BVRVgAHrsWHRHirv15EYEiMuB2kk8Gaiu1+FhVVl+I+X+l03yj12EZcHSCpqsLE6
avexPSQZbKQzxuWjyp9gL2K4kjnNkxh7UtN4KFPga+sKynpvVq4V1jF2KTAQBR3f
qgBG6f/NZdoazUFOZPIBZiIdOUDTljXAC4hoYDtP44CahThdBSxPpbbdH0AuTGIa
bI1NfEo0taxRYZjwaOEvXt/oNf/XBJVvwmWgCpjUpOw3H6SpDR2sj0aHSwPol+S3
NRKP9weovvbnaMX7/6cowaD2f5YUK7umumgIpU9bO+Fn2BAvzwDTEie8p77DjPxE
ibGC+RV1YK3OM/z77RvUnOmmVebnstkmVv2LbLA6WPGKSomoDIShLl2p+2mT8PDu
RRMTxI1/50E477d8nm7WJVnOoZ1SOEfuy+kmOcuvZMjZzi+hUkefrRPBN0XtrohO
tyUz7RxTt6NSlCgKgBhKeYPUugfQ7QBDJBOeLxu0ZeC5OzPQ8ZKXdSl8EDy5+U2F
IncTPnsmxIueKcFZx39IB7xIa5tyyERr0mZcJe6TmNd8hh59txXzsIWvuLkU2AhT
qFAIVqpMLLrRleC2JpbOKMUruqnPOthlpn+RBqF3eAuDHqNfUB/bBK4UBHrmmjpR
HUxp9TPzwUTCUW9fZwzbVEEOwk1WvchInSCw8t47mLbZGxDeBJ2BAWlNc/zA/KMq
lToaXXth9McJwUzwniKK8FefiTDV3Z1PyPB71ZYz23y+KBqhB4R3BiALqCCQnXZN
ITsQ5GvTQRGup3VqbgB6VS63K2+JjYeepKzO6wf+Oratobo7vSS942WHGdOpmfc4
ZTnWFVzVZ/ru8ERH3ssLB0yyQLI30GLO1bdJEaeoMokNjmZosrgpWQ+5+N1NmNkG
fGYmBs/XvhaWqHBNzua9owiGkxQVolerZXb24rwAb4PtPbYUTwUjvXQK8U9UMc1Q
NX0LoMP7wqhjN0L4GxJspq2W0BnzuaAhXVrOxQZPLetg0vMt7qNDjobGcCVcX+Xi
7cxnpv0H709rapg9Nq1osAbcw6vR36zpQQHDEiT8Qlz3x2Xp59hyf0cd3dX2+UEx
NWm9pp08AwxavdWevIo96BpN3sFIbn8Bm8DAo92i29TtGtlQCVQWKss4jDPYDE4O
m4m0Fu2feRcbAZPGOSFf3Nx0lgNLESizKLDVcyz+L6VDp/VyEf7nzePOEl7CHVw0
L/+3GrlUfSvWeF8Ys9e7trwMojbjIgML36dpH9E334aAMt0193V4jZ7/zK2wj4us
qxUXGS2mmGQcxGXKRmcJQwclHqh6BYuc6Ao0oKN5tHFQRRfKCT7kNPT+ZHECvAJu
etr1SRPZieTJlADtfnXmTW0GPjbfE4WV2aIrAw6dCPmjLZ/FfTD/ffjAeWEFfViM
obgcnz1NBmlH1z9g71EeiJikzgHuF6ia+0y+EMOnPFFfmv0ahUzvfFF8X4CWI4Ht
II5iKd5LqBs8TaREdFIafY8Zh9EUIA6y0lWodF+o9ClkFRibjAfVUppjwz6Qz/2g
+ZK//icDVXZIsmm146ljQa4gbx1V6qvbWKJy3FdGPf9ywKtpVoYb/wdKacDEZTNR
5Ysb+Y7EYa2ffuhe6xER6He3XChkE089x+MBbiOiKaRI+XsZyBDmbK3lv58wzIeS
yjQDj2+C9c5GrWHFLO8rsaUThV2//K6V4vWbPg9Hc6remG4jnluE7aoQD727xqnK
nbAoOx65Snm83IuQBrbDarU3utlP6//GF1BLMhcnig8i5zzkLdJ5WD+og2rqtu6f
Y9KoQ+S3BmwHkrLFcp3txypi9SDmxuE3J9pFJOSt3WvZtpt6vJvWGcN51dPGaZzv
OkyxuMVnofAhzjyQdHtDCjJaEApSfr+CVsoDWgGP75EO/ai+sOutI4iRuvoJ+zyV
1uFUrJgkItXt+4vqWHFffWGJ5fDKxOM44vOJNTag25piDrC6OBFLoM0KaV4RlnJi
BDLlRHN5WQes/r2umTxwnwW9PdWw4b9i/8bw8mJZfhAF5QPxL88vgBAV1jJvISLl
m5vBknCzlzrRQ3fcQxNUMYJbtvMF+c5Tomo6XtYngXA+rtl8ZFMb4OosTq9v9/M8
oBziKnvEmFC3pjxbfP7ho/GBhOmwDxyOCLUdG2M9Bn4+nDiJZ1zA7oMoKcc6cQ2N
py9OvmpPPi3rkJE9qY6WK/qSVx/aySHBnuXcv86irVnzONoWXEQrEkJ/wtI0jBOI
EItI5Hyc9dfL7Dtgc7vkSG/mrGbF/at8ujPhzMtL6nzppyye3qD0Qa/A77Nv2IU4
GrVA6YlmFRqvdcHu1IZNDseoa0i5hyX7Tp/YlLRPUGuVPaOSnSzgCDMkF4do5Vij
PTb16NPzXP7Rkc2Q2pYGC9gB38Be5ArrGmJRNPuLxnOQbw4xGeStGPv4Zi0NhyVM
Q24bruFVjMtCgwi6Dt4eHNdw3mAznNJVYAIw4cdw24WcwXexS9u4eIrtZSFiclNn
tLLrFDa/5Dq52WgRAuyZFGd7HFXwIgxak8QRwFPFXXeVN+R6qIAsX6BvZLQ6YRwi
EuO/nAAEIi4qVd/xCjrUaCBr1ENTIVYjIFi1YLYrvuBOmYKYaJyNerPuA/AZmo6c
EaG2kHZw8dPJA22IJPUe8WNczHBOor7gnZiKneqOOrQtpXSdIVTxj5pPUKOwwY/X
F2JjUW4URQKWVxq52Y/TlS4+emehoxiYtzlK4RZV7ryLVu138prMBE+tIQR69dFC
E3VmSHHfBypeS9ZtLdm/yYpT9DqsyoiloSD/vCnW9orbYZbhqn1uB/VaZmRCPb8Q
8SkcKMRKl3VMdOzfdC98166x0l2hJYP9NY28Q9A5vjRlTH9Qy+8Drcd2uyU3D699
zf/ANiBgNVAondlz3go59ni37QfdbhGEdMSkzkwnMMcl91LjUWqMiIYyFhIiI//A
nwNwHLeTjL/qNOvafVrX8MOtCcwI2MSUNycATjnAfwJ3osaqN5SXltqgn3BQFICb
/aIBuEEOiYS0iWw90or4G9/WR82XRb9KzT26iKRlqTvl88OFp/X03irdzDRermj8
NPw8FB3RSLa497wFuxVJtun8tSToaOvXRdhwsDe5l8C9ZbBcLUz6yGqGKCIBRyJS
Nc9JVBNGFF5QFI2sxe3beF3VjpnnvXYpgTcZobuf3bZkxp9OgxJCML2cXkmz6/A8
qfl3W9yAmcgljtqKBUjKwhU+uoBl/LipqEiR64Bse0UlDIZTD8qnksPtqVKRQtE7
pFSJgzllGSmV9kGl6Zd5ntPyPPDhR1E6hARED2VChkkGzxk3Oc4p+66Q7J/q7xlG
m13HrnI53jPeYJEP8iKS2m8OMCjRz8IUvep96WKT1P/VEDbcCR3A5HNBLLNoKoEm
fw/5K+8GhBene1FsOLjh76Onh7U8NhOgLIExsVLuoR04KV/NaJGnYS3Gko3rAMPI
vIXHlQuA0BI35tSxlHax4CN7kqO5flLeJRFtsLFJPJCp+dtrnXtAyz8lVjLiCYWc
x0OGywg9zelEeJ+0K8SREYJpl4Kxt29m1QNGITNL9TcJ74W58gjOlRsUDvWrcOWH
lQT5emu4nwyMl4NxI68XRX8AtuEF9UXFIKMdIU//tlGiZvWwBYa4nE6t0OznZose
eKsN/vC1xd/sR5MWitdZAqfZgUh13c3fSIjINVN1NNbnlzaly2MgzN4g2l38uSxX
ZlyiXZOkuvscA0LJEqdqg/vINgQh5y/RMo4fVq3evJkhE2yPPGUC6QP7szNcZjVf
+VQI8raAKWMqWWOsqCxSBtJjSYvKWl0xOVzxcWsxWGWqFKFuekvqi8agU9LovDyd
RlhtVbrRHiXgb1HULTB0iN3PYXQCxsm8BSacqMzPh5qTAUhVvXd22LACTXBxS5fT
8CQX7erzaw2RemATqF4+ahPGcBb3oeZrdF7AghTt5wwGEpAjMLRPNdaR00CyPX3Q
tZ2pKTICoRjVw8v9rTBRz2jvedZCFp0QBdJXYT+BOkoOZH2CG0vZ5Jm9/QvV7sC+
5q+c8+4Zcts2XY9HyA4h2wdEuSmZrIXwNGJTJNftF2AfxmdUp17OZkIqS2uAmAGl
i/pSy17I8p/IxQSDYQ/zglaEX36Tg3OCafbf+jh0C6HjrgvZhiLQ743cKYrtVnPS
UPCbGa9p17UsvArqffi5LccPGt+AcOOBT+CsfhhQwPLs5VAfQnODUUpb7kVaevHV
iao+3TVz3XlnrV/dmolrOk+ifWi7etdEuSFkg+z4F5nLmgEllpXtb5DU5gQ7QIyv
yziCZ12xZxo26Vu5g8OBSs5RoLo+ZrKou2twi0alSPoR5mfrjaSabSVT/Wg5SvWv
cy+hIahftfLSs3zNPkacmn9AEGKA4BpxgyeTT9ncxkblPeqji+bhYL8uJtwpo4A4
6l8fMvDvwfaU9kn2qbFfKFm3O1UOfnUFUS5Grm2DYJAit69h+u5OoJ2Z442Qt1T+
vNdmk8FVjEjdiLo2rVqb+R8F3Ax3ALhap75tqNRZk7XZm+WfaIl37gjcoyQeVErB
ux6CpiSCwI9IVIVeDbqwb5We9LRrjSzPIwY/hTr99TxtnRIctUJ6XxuuyuEzkfkq
B/cilkAqSsGE52l229yOr9RB2XmI1rSzukFyVolkno+s6jfiJpRgUaL14GLxpjMr
5zZogZZjxWFiSMpd3GVP8YO3Mve4PtQH6EcwIPiuigV23vvLG+M7KRhdRY4fZQ5T
FRaGDK0mg0jLkKz95AaX5sdYqPTC//j3U+azS7+c6wrRdNmaMozZ3Brgj2Nt2/Lb
fYxqIQXiergd05FCnfUM1JGsQZoriGOG2JkY8ivviOe0w0xkmPGpDj5QrUedGC0B
6CwM0qTSDUZqqzgrV8DSMiIS4u9p7o4yCzeVRA40JYRg+eUNrKv8EUWM++5zDgBd
kR05f4XTwdTTobivpwBhv8Cq+G5eU1I5HA8A2kw9/peI1LxDsqoEKnlhdnX3Yykl
hWIjaI7UYd5qTBiXjfoq2I8Mvczp2wzyGzwIf+JN3gqxVb/mcPkNrJb1qOucfEyy
FIiWBRTA7wNamqbdymn1brDsu4xtPUu/SuOEpwNY/uf4lCf3WCm8znXUE79aAtuq
i77yidM4/IOehDOTkd/IX/S+7LWSt88PXPaiDGeN3jUaWTY9QN2XHmWHN3NTmsJV
YwNExCYxWNC64M8V2733BL9gLH4AFThNtYmxbZ0EIziYlYE3zVWa1cHg8yCsClTD
iLAIpiw3kabFoVZ5DWJmheQy1skHA1V6hIJSuPaD4ar1wgXAJTpuD88TPkK+xxAq
4itWvp6vhKHJCscighDJoSqJKsJM8BKfmb4kIknkTJD5kPv8pB1s92t1OlBFdKAn
MaVj85rqlaJyb2epXsmoNAYHRw2QdoXg6TD69hU4BFwzutfxBFeXdfmBooubfX2A
Ymwjdh2WfvInQLWGeWn+4U8G6vTLwrPzXmxfgEKboAjX5R0EVEnUBaMZdOiCB85I
0nH6c9fCcWqIEIDSC8ZynuzGbfxAXHrS0b/sDVZ0XIKUzpGoW98YcuHnfs6Lz+6V
CZ9UN3IxgX8Il4QxYU2T0SRqiihBaepWvvhnpdLH2OlEMcR4tq/icaOxo0Ms3Am3
IoZI9R6tuWlog3qgREufggd+m7UpXLvsSljTnZX3zxJGzXCV+6hINEGDTx5Iuyjl
GbYdySGw8mUKlJK17PNXk9rV1PKEd9/SzON++pXHBix8JdVwdk8yvNnYc1GqfwLy
gZLo5yvVyedqxDjQV1EnpxMi5mATcGbG2dDe/Izu9+PwN2zssVFnY1pilv4Fkwgn
FTzbJbWWrJj04nzQ3b3Di8ZxvwqtzV6LCXIgVNnKFDrxHxznnP4ABvauTs0tBfQv
frOoW/eSq6cU+/xWirTb1+LA1YtdQAqBzbKEWU9NqyymCLjjkrtFIGMXqNo5rZuU
9esVTfzyoS57SxjvucupSxn01wrBrytVtZPIT2vjeLC+Adxw+eQ/WsJCyT18iJvn
R3RcD4q8H8wWcZ/qnKI6QApV6gTVt+npUWPZOcj/F4MDcWSBBXST1iswkgTqWY1i
PsTqwkJR9ZzH8Pfw7X1k2dTrN9FVnnZ6RjPX9STNNhsAcWtDIfQpj8RroKJHfFY2
K1RBGfUkHtn40wzpFmXQH+DAV/YQFmQn/x1mGs4F7YJyTQm4oaphucEuyO0TqoF0
4NNVmSnOu1UcEAmnFRc8Xq/2Lo/TTqfMi2giNu7npxmnnErkvLn87h1GbJkRtEnH
+VUAuDAEAOqG0VZIxqXfDVPVfIZ6QpBSJ7fCuBxFAiJEf7JRlq7nMVKpvBKh3hGn
OkuKeLArYckC12d+rUJTKitHRo4bpMtQmmRV9bDy+QKMnnkv0+pCu13opp9j48Zv
KfhdorK/aYQZDbUTRZ+WAGR1/1xJ1eGwfOhGATPPI8+T1WVty+ots5qpIV0JYYqX
4LqLrD2RHuYtdFOUGRmVdTnNPWtricpM/D6m3kL6Yx94MFEIQKbN9JKGMTJWc2nj
WRYZkbQUoGs01mWh7idDDNii0UQEikHhjXtyo6rAUzTxcESr5gFOK3x1lJkFZRA7
7Sl3Zid4f2XUd8i6MyTnjUTQ2DbQ630dxEA5+TnZLyAWfqbhvICFAmFaTTn2QTCf
jZ7np3OZJk5c5c25Dt1l9opBKh094TmevGyKPlo1btnawV6wVOgAzYBudHHRPm6m
WzonzCDqFpF1EP+YhkkgDplikcGy4yBF/ZwijA7KhmkOAPsFqlp+yi3u4nuy5dNW
RJ0aXo+rjPBFP451MvfCIBj0C8jOdPo0TWl3tV3JEu214q9SFIIsEOt0/A7nm3+U
hkxmZ97dqrMGPzw0zWkG5WwGjBSu6wTemDu/23awOIvdr7Wn0hmesqpRudf9Ud3a
5P0CrEbGayNAqZHAbYGsUx1YHg7I/EwSBs5xRc60nEmQSl1WLHgp79/uK84g3D44
mxKGk3lPObSIftBtBB2KijunekMKN2j85714g3rqpR4ZdOpFhlMtPwW+i9Lj2VQR
dcNZfOzhaJMeUSIjmJLt4vXrpub1V4WOWnjClKC4QkR5efGn+Y1k5RHPi/tXrksQ
ajaqTljMAV99yLd+NzYdjS742/dn0Db2pg1Xs9srKw/WDhRed8wJXiw/1b8y8ppa
mOE/lxDslymNgRdRVzXc5cOQCE9jt5HmKn3okgbSQNKJR19ijFZarF27mBqugL1b
9WDCpfVI1rnE0H069XxaZf9k9Yjd/ExV/kaGfucjHWTm0YxsR4drWkOBliwfRq5a
bY8ILTKSsNuYCSxHGi/AFYDBEaP/VJ4GPdh7LscipxUL7Yw6j66HrUHWQmFD/Q7/
jErA7xBavjLl5VUHkGPqhJGF4OlMFGRTrUabv4q3AyOm8T7WUdTlSyGxw3wB8stG
M2rl4g1J5EygY1KLfV4G+0t8slmB1RmXiMmlT8ZPCnO3C+qYUpwMnvoGXS2/1T/y
qr2ry6n/pzyNXAo5Al2J8fddxm0TqQwKbPeHhH+SbZ+v1FZtYqFhZ4w9XqvfHlR1
l4FET8lTsEvTjpErEr826z6zcICahn3lP8TGyTLsxUI/vQEj91NdshiyccMiL+4o
WKqA3IDv3AVdFHJKvK/Qomw4codbvugtKHpBfxym5Kr5mvVfnZWEK3Z3JJpVHfa5
aPeHpWg+CqfFeo7LMhMTYRF9mayDkjZDzoiplKviCbXYbNGpb/WnuMjjCIGjm2Zr
zR/spV6Zj4uIk6lr6TjtlGKBgFF3/VdMnfEDmHvkGS2h9Yrn+YOhiwDDKOvu2qdM
8TPFLGoWW1o9ajyjIrZ0bvwXFhhEpGuF8+YTdeg7e/tYLVcMMbuANbkrMiIATyzV
6N735uAGYKbkDxW+XnZm7ggBpbtszE4Qr01v6UoyN5sa4R3Nk/44zOLMhCs+Jp1d
FmWedBbzBEF8x4WkAbZtBJd3BoqJQdKsvo8Tj+ue28hSmPGC0OuEe7wjQskNBsRA
3ow+5Km0UCQUzPD/RSgrSzc/cYE4cyT60sW/zQoraYIOdnWqMM58D9D7H7+d10DF
5/PU8jUkoIA4uC+TiTEUko9t5Uazeqy7SdJeqXju0AV8uvjdRAhbW4uk59l+vn2y
J7Fum0kNu/TLmK+7OT6jMHxFIBojs51qFwbi/nyAkMCtZDVpYXDBYUNZ1oqyDp/W
T/KNlDDoRUhzQ+iYDFgWyjxHgBvw36Tk/v72qgYMRcgeqny9mhrP49MIjk4lrEck
3vRPkMzHrwu1RnSClcbZMi1IyJMPk6HcSrDmLbeEngYdQ1NaPn5O6IpJht74Giiy
1EEm+jbCMln4LADOP3xqjeYlnfQ5WmkS+YTALbZ7Q8uEjCuMwlDwkBCawrJMQbTn
4LjU6slcg/v9HcAsTSoA3XvI81dmJVR+HqaYDz691+mLSPL5tONTyCjuhq+Relcg
m9koeejZDA0MgAc36WZuk9YrbyfOtHd/R/mWSZXwWhXCeWG7jcgo4YfZ2w443mys
bAB37UTKLFedmh3mjt+4LVWz/D2jdi7+6rXjKAj8pnQjOA3xgSe4yQFaAY+w/SE0
fUS43P2ivVSUw3Dih7jAFiF9bqrHdprbktjOzvKgYtLFGJP+QMCqrGnRd3CA/v/d
JCJIPrjKSZCyiS2pDEXwqfUnXQYCZPvhnBS2YudvfN1oLxhr8TksB3fTwBwxV/jM
M2ubZMlujDtU8CwZZA9pxqoeyolkmhIhk/6JAL8FGvsVumXXEF6iiuZrM5h0FcNO
VIyA/Et6lX5kKS1J/BtZrXEVggOXxd/cB0KWJHYE9/sj8nyn89/Drs5EVKwJzvQ5
8+Zjmb2GDX7OLsbSwVP9urf9wPvuS9sg68/ekyppgh8mE7PuaLg4AptwlQAz8UJB
SCxMlJwJjj/J+sJYG/DJK8s6Xy1V+scyDtPS1DY2ZSIR5GEIUJLdP8ejocoIZIqi
JYcwp+Z3p0g85YlOEGzpGOKZqW8GYMwG5exDzIUDTOM3Na/U/Z+1wkYaeNvTXVtc
nqeUUa/wCzge4QnipgBfM+xbC27bQ/l/DOCV33TRtBC8UUnZ1Dpon5a5w94QW9Rh
z3hWDaSqfpR3+ngQcJcDbLlhxuOy4IhT2iieUTPYHce0YEhPjvG78MnCREsBjmRX
FsTfbf5mawcVmFuIPTVJflpiWGlf4QSr4IzxGaXTXNsNv/t8mrimWiwyHoqtQtTX
qrk5QVsjV+8pgk/+rnUdeb1jqro7K2k1XHTCgGfPhAiyrqUrIy6s6IiZpF7421sY
lRMCF8OhOp0pRyfo6VQfFdujH8CuyrTJ/QuRRdkiODHyJ4rfg/qI57alZTOFMvH1
3qZdCVe8Jtw3Rxo5+Gb3Wc0bbo5t8BEzn4dz1eiGTOZNOPyLyYbbbRhZWC4pjIIB
An74vPSt04rtp+gvdQOceFGmLD06REbmemleYn9hCoTWbGbpR2eXNAU4h3Rdyz2Y
tJrFNxlBHsVrLV5Fdj/Poo6zbupbXaY8v5r3qx8zawkzd9qjBDePu/cxEGlVFHGW
3qF8mZM5iwNh8ZKFBT2xVdfzDWmNTM+5UGHvZ5D4jyrB2t306qd6wayd6xoIfn7m
8Fotmr6avGpetNEa91bQP4QBKRu5NfUsruRqCVycFvCaQTGcxH9HbVq+XpyXjtQ8
foiLvAHyC97QccrqwFH/SMHX2E+wq03Q2DSRhVbrvC9Sdbub2AB30iN6oyWm7EFS
TRFbGUv+9VNFCAy/WrhsR/ZfL3dVBdtg5/QrFqadiIA8CXXrgHWmL0lgRUt6pLy8
puVa/rkvasaLcSsZB+HDhW4a+lO/eWrBgqauT8nJ5AxwaWC3JQorTHZ/rFfymOvs
H/3LoSe5tWi0JLoXOtIkh3pumdHgZJhAzx9jznZ0XV6NpxcCbPpmZ6AzsWtVlMPc
irYfw2idxppX/JFTYZpZq0LSYuGI9qVv+iSau5Y3kirRHbjG5rtW+QOZn415sD9a
vP6gEB9QpLgRrjVB2yZT7kcu6r0ESb2gXHkCbsr9EqrUBvvaykxsbNWL7DBPSwpZ
pb/3bZQxKVXGbG/Spc16ZOPYe0O+fQBz6c+DOPPjuLi2ST5zcq38Nw7mbjIV2Ylp
KrH+aAjQfU+jGO9AGnGuqHOmmGS483C4W4iOX+vvDlvLJA1m7f57st3h0ReBUCPr
wkKAkThlYuvxAn8eg94fq6n8EetKWszBwTNFva3zTFN/ijIoYaH84obf9jO0QNyH
qcz19+BbALXDaS17HzZ6CB/MS3XUx7t+m20LY6uuQSXP0cV8OOmrcG6B2u55hyBd
bW1G39PZnmdOAAT3fUFC6J8xeo6njVM+1mhKeL5UHKObQVHpErs6osQSv5NRgIYo
ekMi9uARqofPZrTV0WhDhR3N+79bkcBqY6SWBXTammealhsbk5GznjicfgRJlpY6
LwfhI+XxbsGDEKnnwDkkhadMg9YdPH2iylogUEiCk/26B4MkXK8iYRHlbnymsTxP
VbWKIqJH9/9jQqj8QY5WiFEN/Ej8jm7E52UrjZS0QRHMOdqLbgcLWJC9cp4T/is0
VQOWc+p/ipEOMzaimPlSUflWktj2rfWNscd5MAyeR3sZHw8bftzaT/6jKNkd/Wba
5giNMyx+wWuS3pYunhfymugVZSwb1tfDHUHa9gV4hLJAjasHsLfdPEHu/ZAhdSpn
YU72brmBfA7ZKZCZJv39lKZhFcTcGn2W/8o/D7fAvkrCN+YDesYEXeDU6CYrR8ij
IQ3fFx8oqU2IA3taa3aE4CmoykyUI6AylYkNdYfrCPEtNsdw7GINt3+UO+OIXXx1
yHv+jvSZIsRv8W5AFU08HNr/1eXHkb8X2R0vqffTNZ/pTx4y6ikKcuRQxMI2CZ/a
n4dZxAwjr6XCKJ2jzrloP4tvjG6d8Z946Bn2usqgjQ8OZYyFK++5B/IDuCGImYlo
xHNM5M1JC9eheFHGeP8igqh/FYvh8EMXdJcodwk6jOcIbX0+3cQInMAAUXlAv5sI
qBJI5y3TQJ1BC1dV1OACWtpIDz7tvVjOEpvc0GqJ7vKfJo1d2c1Q3fHn8jy86alP
fikBFzQlN3F35S3Qx/qwlah0LJpz5OEFCFZQBeHXfKm0TIFAMpLqAQ3XBYsw/1Ot
/pLQJkEl3+ZQcrvoYiL4NVFljRhGX4LGOZAev3jI0IZNvWHDhDRbTIxKLjvEh52R
e4csXAtnG1w4hvt1C9PhmFaU5loYMf2+hKpz7B7OwUo0tvjUR5CVPW0O4WVADEO/
IDRxtYPkOcbUqasvasGnqw/xhRQUhtQbyschqAlKwPBJfNbqQU8zMQ8CsrZY/SxM
tneCgRvLO4EF4+dcRZbqIsrRsNMmpusDjyq38B9ytcnEUCNOyjypH5R1l55Xs6Yo
S0MubrNTOY1tTBDR+MoyxyNvC5ATUzEE6kanxgJU/U2UWP++KWw6oZyXN7dxVlqC
kuw6CMwpPA432VUrciJhXziQ6vnW4+UYHx76L+mmFejYF84w5YVPkABypl+a+EuV
ZpawuB4+J58QNcEmyDgItow1mz2Y9nKJTmntpt/a6hAM2N/SXZb0Ji5dAsFszESV
Gr3H/ERp4eRArzykpgFEQ6mFd86Ah8nMLDCLzoYRIvgbbIvzgAQnihpk8vwp8AcN
BfQ+ba4irJ8VIVtAPR91a1whxDN3LEDuKuTrUz0/Nb4anbfsfHH0WITz9SC5ZF+5
8zIgYOXBZCAqJHkq/0geWiM2HArcNmqyg0hvGFp6eKPBO/rbMBkW9b1UAT3X+vxP
Kd0HPiSjOWQuQpRYKTqAUiGrLVZs8EFYvEGIfmG0c/KPMs6p17Cn8PoALMv0uMrG
PxXVnmE38BeHPNL21oInXKpAtjdzDn/OMTHYZzUuCDmoq4G/unLoPXQbrXf64wBa
ZgJU+igIOK/6rChu4MTuEIoZS/QFrf5CkZ18ZZqwMuVT0gD2QDsgMbM0vGkMrY/c
FasvUEcp0kgYyTKlxiDm1lkv3EIsvgIOK1EU2R/PDNbgH/+xVaYPhwwTvGkNq1+/
rlrNmihOl5n7El8jB73i2BiplChOhgxg2dwIPyh5MGd+VNO+g89De4XVGXkXPrR7
dAnyn4/u+7Nw9YriHhs2VsZvR0iiZRYD2mlHdfcx1ve78LBdJt8C5zec6iF4b0Rr
PQ8wZWIma5vPLva7QVu0xp2JuCnUTjaD98oHinUwG8tjIYsyqief+muypPqfIjoh
zz/lLaz6qhUCCAtQDoZT8rqwfG0/viQvn6tiHXtK+Kxhqs6EO7yEUV/fAp71tFO3
8JBSKwdg0bW0ew38X3kY7zrwEMS2DjSv04AGsYmn8fgf3BvMKwCLQYgZLOH8MjHv
zgv5bT+bj4Iq82PBQLZP7ypRnxA5FHDvJ+JJTJsDUFXmyEhfvPp6ZM6LiWXdi2bb
VLU3+EPDa9E54bT1J0y8KkLxM6lbQUOr19t0uLXAYwtFPWBR9kbwVDXV8mzMIKZo
JSbnv3Tzy87GhthGzoHqMGUOTmAvFU3+oENJHwSsrN1BQcxjyRqdrWvW3W8mzA+z
L84cLZmlivgNYse2jfT9F19M0OrdlQEpQzrwJRz32MQhmBNQ7cfByOELq6lQm65p
FMqvyqBWOZvrChhHXvUz5zkuCBBp0vXSr2B5e8VR4oxakwGgE6clGY/twdsulxPc
A3jWxeobzSL/gDjNhu0m1PkdXOPvA9bpLN9PcqtY0T/V6zx+yd58VB95eoH1EHdG
DjwwXDTi53Egrt0ICiJTNLDRAZxjcyIPA6ik/lyPCieCCyq+Vjnwi6vndPcizE1s
M1DF4IjJUKZGZXkrw/0mJyLfmZUfRwQDWhGOYlykpnAaZCvsy9h6cACDcDAyFEJj
Xdp+DsVbM6qMZ8pqxrHa4Mtyx//XBp5la/kT25GO+sH7mEhTDfmxI8wYwT5dYIyd
VS8ycs8OX+7mrzq9mwU+y4Xa1Xr6FOjk541ChSFblSliEuvE9QPilfXalGwdtN0d
wHYBXhdXccC5LRp1uyjugaiKQZPPNWpS8kjANMgZlR/PQ8e/gGLAaspgPb6ZQiI+
EtmVkx+7RiFeglN3ksH83IvNjiUUCvz3U+ceuVNFpInkyW4uSHg47HKlFua8zvKo
9NmyMr/9SVniSSEh2qGTk6Xr6N5PVLlL6dNRe2rfRTV5n31OD8xlFn5JOBn44ZkQ
efbGYftkt/FLl6kC9Aep7MV+vDWCKB5HmhoFboErH2BHbGyB2y0r4h841kHAhqmb
E1ZpPBhHPtlsbMLCzTJdKstRrzEzK4KlnVRtoCQJ1cMOOUaE92Ut3EyJKA9sb6CC
NMF15l+Ptti/4iAgVLZwLn2W13Bb1IgShKeecTH93Dm07DdpvKDbx+n2TSM/3Zmb
Abf0GGZ1Wt1OXv5a8rMPA3qhLWBI4lqWqgEfopjOsSM9UxFkCDkAnkhVDukG5Qcs
xa4KZ/ZLMYg5dM6Z36Mwh4+2tSmvShttokBqkP8TGG9YrHI/VvX+jXcXYMXshzpB
cwtYQJ5GoOaCvGS4v2V4s63TZvu1VgowZtfqDhUVZrr8ma8/m2hdeUeT4ALrx0x/
B9A/8cJCeRDfxM1h+aTdmjyvUAqOgoKvJ+QrG1/4zvv7FSxDGhSNxdyQc4rAfxxm
J/L8gVS2H4LUjPPmFbKwdLRSo/HoBdZcJz18DkRVVvMGAMUD++asELkegUbcsExk
A6pF2y2PkI4PqEpPeQVfkhTxIjAbG0q01Oht6w3AU8iHKhwjCRjPLB5j9LRc/xcJ
7wrSXFKvc1s7PVV+AF4qt5GwdH9KI+Hd42jrwnDasgOuuG+cvoKqCifPmR39ZVmM
OBKSls+3+yBHbcqy3UrUwj/x76FewpQL96+tUtecxu7fcM24ArsLQs97NTUG8h9F
boQLrGRRyNizCI1ySvxT/nW7z2G9aWRe2Ce2KegvFXUa1qLe8tDEwHQ71ieGCmpZ
/HW/OVUluu3qHTAXJ07B8DbVlrfY6lyZyW6tVF1RdWlIegbEVlNFB0VdJpGta/4H
UhwpOHL+PXjYll1nKhXMHq5wLrkaodT3+7SNCd/2E7ijXoo2i5FIyomoMECfxbDR
spPfTgrqUwPIriLQ7Lq6MIpvVullbuwomhCXOt5C2wQszZ+KuoKGBnCVr+imGach
I4pAyTAsyRL4XzoGwu6oDOS5AIo0uSd+zdpFxKmJNNFRXYXtRz/pKzscQJvHbALx
cbbK/vzNvo6gk121zqx470yVS4YVrrHBMa/Z7iKfqJfPqQoxiNPB0wdYg5ZyCNel
JUkiAU+VFjeKkG54WG7CsMVKChs9dRqHbQbIBPjmDihEC6wdr0Zo9aL0zMXtF+nc
H+DcvKu4Y4X+vkmgIF3prfzmn+YJd5IicrGhBbLOhS21tX6L/N/8L18JFKoXw+rS
m+gepXYfa83UFy/Nyupqt+uVWGEBYs85LB8TQ+gwi55boLmBv8bBiCkaoOGAiap+
Xx0w+4eLyoEX00RQd/iE4ENxIYiIY4T6dPTztKUUHSQ9YpjthLXyEL3qZLhfXQyl
oIXTB/699P2L3FmlHfKrLQZQOZLgvgnqcm8ZhZHNvLydC9OsCndGYjliuaLnOgkH
P99JfzD18Mn3Y6u944j4TGpksJXjFnj47IlJv1JJ/S9rO7r/k2a4cZai6cyLQAF9
kojdN+AUKSSa6dIYJHiwQxHN3ylRH9dEly3lRoBEBke4gcvexYAcrlSZ2tmK1S/8
SZMWyeAcJElUD1YSovLzvumQAYtD5rVRwEbjyd7He6plhtUll2rMm9cTeleX47U7
+MlsgluSFMrIqIlXu6KpKFNmGBBtUdeJRecD4H9gdHEFH65ujvmOs7rsbjdiUKYv
cpkYmx6+FcC4fVyAZcNG98B1hR6zWjiv4/ETASa7AYBtvC3ntr6sdBUQtCTdlCos
wRcYGF92G25eD4f2jJM0wH1QLaO2ix3sF35E8zmpds28RYm0nGtqsR9fqYticuz8
ZaYhZkXD6W/hNP/j/fBJh1QH3B6QzPFv+nWPqo8eAfk8b4bt404uavcNps5FVx6g
duoGc8vU9wXoVCco5TlsHB4oWlGOaRpe6yPVf81gDCK8StlHRwcCLMGZ81tJoJx6
sQjRy3ocOFAGCUJOqXttDm7OzHFld+9l30CsSSstW9wfdNuIL5DTuc5raEUlvG8H
ihWCDQxFM/k9jN2s5A/OLKuVWHh4f+9+dz+IuODm4/MiesL/qEnE7RMoIxQB+C/Y
UrDVdfAcJohV8z25PSKGvuRu/Zk3v/Xv+NcAR0r782Yn7/DpSk/tQl+kDajZoIkv
FtFf2qrfWFTmPy6m0rj9IfKQAeui6jAGzQLeZAmYaiVLqagwOZAmCvuqQ6hjT76d
LmMIz98Q5CF0tnp69gHOPxui/3lYNcYF/WjPaed6WBQXg3KN5M5+A6XwqcIvntPw
ghnqEcnCyw8xBAVlVuKy2dtL/s5XnkOCg1vcaqgtJq4OJ6WnWFdrYTcmns09YJIx
7Zq9Icj26aQLwV7WwFhlQvl9FVW6lxO1HoK3agFgjY/Th2DfzKDLZvKThiK1yuS4
BERMDu8Wsd0Gu4u3oAAtskqBxNJJBMnMFGniwdbaIbNXZF0olBoh7i+KyzjjwYx1
Bp2G1XfV4+CeZTPECPSFvyYNM6jYMx3DHOnEQM1FJ4iWmo1GeDTPRcT3ZPZ8J2e0
jMpaYGModhTszEgkAIm+SboOxRxJvv9ouDeaxyfQydutD/ZO8ece8UGamMPDrTXF
5S2mG80fGZyd9zxzspiY28doGzCSMXrAWCOO856KHpDRS/WPMhlXbb7HH50ZYOA2
++ORok8FOKLBBjsJ2qaoVCZj8oka17eceKkUNF+a0XOxI5rM81MLfz1BA7XUrQff
C0Ys2JChrtHH5KYDC0S1gt0uj9Z2QcDtu8XB1qr7mQtH7GokWjGsXNEtMgzAYd+p
uR0nXYsmr8k0X3vBXBXFTfLk4u1Y3gTm6JuHfWAaTVwCmCO+DA97W1dgt9eHWvD+
epSYfJZylOqjYV8LRuIH/9BfLmlRHne6S5zq7vu3dU3nWw//9+Ag+RjOc4xJ/x00
lh+ndnZz7fYSdEstbcR3G+x4nFyFn86VXH8ZJXhfW2AJoNRTWzJ2+fi5C6MV2d0a
KKzXyeMKl1ehnl7J18tLyzaF7QJPBrm+mvaAlxtKzkoVQr3++m2KXRGNC8ErFSnW
J71EI4Sb1OjuGAmOBGrE7ckd3RstHXBLbDSfOlJfKCerfPXjsDTyjNvPY+gNUA3X
lnXnYSk8SQAMp/XTGa30rnGQb6xfH5/g+gAJdsU/lCzOq4dOysFs0WJ0saw+nmur
i3Ltwb+fAQvyALzDB/Evbi9efAj8Xjnlml09pnTFTcrg1xFP3YdgaLTQfifQFPNe
APqR5cJk6sFi7PWVDq0VDO52MBphfmrru1ROGa4jLKsxp0/qMZWDtbjWfwGtSr4f
HDk/liGX+RQNg5e+85ssT3yiwKZOYlAswDtkQ6BFNcY/HWN+J7NHr6PwxYQiLSUf
cCziY0cBx0yWf/NorU5aqAyPDAh+kiY/Y/4wDRtEDP03GXe/97bE4ep0xDTBcRpC
06TYfi2xOVSBMY6p4F/TpPxTt6chUV7hM/WCBESECaTfosSoFHr7P6L4g6C4gavj
6T7ySZBkOTx1vHbFe+B/lPvbCrzBCJrA4k4TgL3yw8SfCh7qlIV34mh3DMhZ5ml/
IFay/rKGI4NhX2baiYTHN68r8i8bVyDhdfY9lzx6PvI9lzeVqNbp1u8KcBfelGqF
KlWJuy7mjQuJLFH/GadX0GgB1xbkjsm5KRdlfhl0klLg3RMBGGIbndzbxSIAtoHp
HemihFigpWQUa4wxkA/g3VQvnwMcLCMvVbtpQK+cJiNEi/Kn82F57rnEU1oWyos/
wsYSEobZT7ht1+zKuPjCRwGwgeIjW//nJ9baidGYKJq3GcyA6a03EvT+yFEjItZk
n3+mn9lXHqof82T/nnFn0HLd1fphQxi15SJYSeLX5EgnnUsckvhO1rOLNwU8Isgx
T79PfZXizZBP/v07bTpFpIsgRv0dYRmb/o06s6ebUbpjThI6OFy6pg5pGFBBY+8j
OsEJGbZOnyIEQwlZ2lSnrIEPguiPBb2s++nzcGyyJds75mwLXn24NWZpNB+ou0Rs
auL4usuu0Q6G0kpsSbyfw9rhyXSdyeMal86Dze/schKFTtRQ1caCuUPUDnJhqSQN
uOGgBS/AS5128mjqpadP4Al+SxA0UTwMVoC5/2J+NLEQt0nE7KWPj3fDtEUzDFDi
H/y5XWnD8RPWVRC5rKANrLmSIPIu8XPlMPYRwqXNWVlW0TIYcS2OtBYthJPjdvIr
1D5bktvyG178uIPqAYAA5j2d6rOT96saXgLNaD2yCvvhRMaop8ezEK7aKo5sphLY
PCBc7EhIwvvkwFRL0KZVsjS/FHi79PvZ/fwBt5dyv2hCYLcOf0YNddaxC4JSQK5c
nfN5kF48fDrXNbvqVW843iGmaQOxP++yiVppDWlBnYCJzdwsaAabXVSrKm+0dfuW
DXuA1vY8reglRRsje7BxCKIFjS4Ruu+TJz3F1UN1JJ2iIFOvr6qMEcNfa15hIyul
B0H8KfhHnQbbCCcGs6T7Rr4NrLno3VUSuMUBmzJV7ONVKYxfFLXmAFNI7lrJszjc
TEMuHKQAZezu/tOxhhKevPsA4Z6WJN60MNEQsVe+E9L6wuoE21I5dUn4c3tHY0jw
oG6PsJXLlQsS49IrCRsV3LI9BDLEpkPWuhvg89nbbYgHmps+gJXLWhPo17GXZ9tb
OOlfbBl9yRhyKD28iWWuZ/V12s+ALp11ppGyoHwybzlfFW+FD/XfrEXMKxRdFpo+
yGRiXxFwuJTGwfjFNSzQhrXHMVGOXQBujAyTh2GfmlhOrg4KHT8ADwTeGzGWs+Fx
Z34BSRpwA0w4R64jCOw1EYwg/xHpa8TJrQkwixGYMXZ2sI8jmiVDxMLaB5RV8+/3
T+NlHILSiJWcxUMyXDyltMBTRjnjL6QK8CS1qKEp+GGpuEyPnkLe22alf3EW/rVS
Sbo4QHsjyN0PYR5xlr9pC/2UqqQ009q6mA6mlnr0Os+aEU6f40IdOyUWTcgUaKij
4p0XAPjpTCkr+aXj2EkQ9oCUvI/eXfU/g2nr4vMcaz21U2ARoCQPr6pdKZGIYOSU
DVvkvG8jIAZzPuIam0R4xprMhOT8/tFrS7wAlPNXKMAnRpdzXMVmhCJ/SgMJEL+5
zZVHwsjDmQXk4dT8VIDvdnXo676UIYmK5kAe7sviO4X4tIG4Q0L+NMNB0lqcPfhJ
hUHAD73hqGqodBMP9rKKp7xFF4d3MEcko017ZA202ncQZk/TTSBzjukqOzr444wi
tG255mpn8YD2r5V4CoANCA8KCP11dPwba4QeIITmvlKjl/m8+YJJ20qw6H0AmUGX
kl/DVaT7cjdj1yR/gdptMJ8rDH11CI4hWlxHjYkiJtwT0tG/rc2h8/bYlpoxA7fO
RdXPllcw+h1ofCm/fOTa9OE19/pPUMLW5ZOOtoXE9aSkN92HtPEcvmrnjXzvxK0R
ekfL2VZPxUU6nGvTutRNnCPMJHV4cdgkRbPeaJA/Swvrae6ZswwdM+xkATTvSjDM
dfv04AfVjzq4+/e7nKuGAb4oFKrE35ehI9R/g98vg8i0fZUa7P7vSplE6MGCN41r
5SzBlyzo0mKBUEAeycZtPjFyvwhn4rk4RZDv6hTDPe6k1Ujq/QJX/hf1+75yxmoQ
GKkCeCFVB2KQ2ccC2pBAVJ4N0w8J8hiye8zZii+b6OUoAdEss7C82sE+1xv6kjU6
DXevpeNi5uW1/DyCpUTeQ9DrPcU2wekCGayrUjyly2mRqFhZYM1YuW9IS9mdEA9b
k1ZVVPXQjNsk49E9Kf8CrQLpMA6UD/gAp+IPGQfFynqF0U/KsKMd9YY28rqM9Dvl
xZT+nNttUPDtzjoiLfPwkEQW3uGyR8BkNITjUoaeqfGsTXpdC687oWLEqAXx69ua
OfT2B/bJOK6yhstfOe+LNq/YBBpn4mikLPITy6duOgGOiGEsPEt8qY38q8xnfvB+
71edjxGBu9+yega7nOA8VDryRN3rCNOB3zGPaFqcR6teIe1CpQjKOH1NMEaSi2GC
IaGp/+8PTTYDR1p8Lqhm95p+oN8r5qDymoJAhi/qqDGcvZ6OU6uz1c6CZVTKWtYb
XvSyXxGD6EJRpE5ncYxUhL24xtvAxsVPopnjKOFQn+x3TKQafsKgQWkAGNuGw6C9
30SW1Vq9VnmRWSxQ8eov/hKS/dq5ad9UVZkwz+VXWqQ9Kye8xLg0G53px8v8XLmu
0K+0Dp9Cd2uv4h+XyZIrG7Rcq/+/2XJTyUCxHdk1Flz4FiSUcScVRVqPPIKrbWhm
cvF8161/sYFLI/r4qTLvpedgarywMXs2gjEE2IdjRoaPDZAKnqqJR2yiIjw3rPqN
bc7+42ptQpZA3XMuVbLc/g+mI9dRPwg57cqexvRpiDkVbzO/2yXYx8qjSGZrDA32
BBIOzBwY0WmUJN8RpFx3EyLy4UJibHw6kQWmn46Ci0QmUSRBXh9p3mCy9irbPrl+
Xc4yS5RpOCz8N8wCzLKyCcCBlCo0ead0cIkAX9G3fXpl4ErSkMxzlUtqqDCVO/0v
FLG+lKhz+5jC5RmYDoGhwIVig97Cj+DCXSVH2v+LS25MXqCYtL6hn31fpi5bx09h
VzLADAgosXl+5KFDDy3Klrfa5ILw6m43l6cAQUZq0eBiaTnz+iXpv4xD/9DbDpWi
vGAURteME6S3gBBbNL/BcFUlYO4r/TL2d+0gVVkQHWz7H3Dj3DinXtsuY080mzzL
bttKuJdpo2aX/AeCmsG28pNRgpGBTZTxZPazO3YPDZNbaOHcoVg8xKAUYAEScYpB
bRdWGwGOmXuhYlU2ghZtrNWDKi3ed6jpHD8YrDKy1w5R5vArYA1f+lTumFE53aHW
FBhw8Rmyi0uXFH+7zj8IcXAyQDHO4fBjw8xwvqwCX+69iMkLIoaJR4UvR+hJVDAc
QfX7FfqQ2VVO//6i3MAtSsFNxQqYILfRsQyUuGFi94kN8fjT51fnKQaA0QdElvDG
A89214zJntGEN/sO4xRDRg4dJ4jxKApEWV59cAMLOolQEOXyCZ6stOeRgGuwuWAV
8i0MOfEJFT8u/k1vlXyHmJRYZEEG3EZLPbqnB59eBKMg/oy1QvpBe71ImJ82boo/
qT5kaZqyfqOTXp7zHYKSl7MwMHEiwUNGX/JaPmlhwb4Yv5njBnzzaVblbHyP2w3y
JV3feCMEdKss7n/eqqjQJ9twHrYr4xkaAiiP/4lL5FlKq5BbGhQJw1OFL77cjXf6
VpLnR6uWCF/7q/N1J4omWRVEx0Jp1bUf3K1wpJVlDYAIE5jy9dDxJmbMXqrm4gLX
d+za04eC7Pl1xo5kxiKhKvyrD+M+yoKMmwplpsOuZ/aDNrEMJttzZYKec0RWIsXr
L5jZSlctRJ/X8tAetLnCc8bU+bSV6/3+H5Pdq0v6JILH3H0VghdVmjgHBQStfYr2
ki0ypmfWMffXw5oyIP/EtXIgDWCfpMm2f8bE/Fww7BdwjcD803z1BIzoEIOCu2Id
B0S3jcV3M9WasDYp1tXr3tfforXeGHvlulg32c9HbS4lAe8qaPoR989+KG2HGtz4
Q24ce/HKPe2D0ng3VY8eZAD0++XuxgXOEmi3pGk2/PFxXCB+iIAJMCfi3wBfoMmC
4SWIS4WFHxttRVFTN1DzIyvyJbrdWV6hD0Dn1V0TvQExDMliDR7RzLA63yv/uJ4m
m9tVx5H6dWdwcl40DxokFiHFnxHO/77Yjc6IGzz3pkbqZYBCDDMECFqu9qWlzIzK
wqXG7IZW0FbCbzRU8wRVOEh9WLggS9eECiOTLs9yPFiDy2ZTXnZJLgLgNUEb/re2
QdNrXg1lg4rPdEeKeS5qoP3nhyrEaesIi8ufKzYx0Rg4tlF7fx9y3a8A03GISkD+
uOPZibwi/yUIrO1G7pB+erhiIEvqV87Ihnm8ec6AzL30sO+EAI0xb/f5CH3MkKjw
C4W+NwM4jXjJMwVqr02cDUcX0g63IFf/sCjStoamNfNiBCuTHPaSF9ID17+zysUt
UTgsPXYuw/l/fTnIVtknxjrdCZafukEQkgN7kQxBqw95DYAqpK5v6P9H0IEArfQk
LQw89WQCFRLXgynlz7VPJL41CzJv3gfbkoXt5jFsj3c6sW4PjRcX2s1BGpITLeK8
XbjfOM8Bxv3HIfSnDC4Yzo9Jw/jmVSErBEhKOtuzK5N3o7ptaZdxyV7cgk74vBsD
ikQmDeSNGQsXLlIhT05ThqNkDPXALEB778ZvGQXmNW0Pz34kNDiqbUfD46sAUSSX
WHLWbPY2Nonv+pbPOZ+UYmbG/kvi7UH4nXdYAvxPrSuTULwiEx6RrSty8iiXq9On
70zhnj5AcgBRc3q1ofM0rHGNuGXQIm9qrnQ4Z4Vrko2ZRUEc/IijWH+zBL7XEcig
aZWlGwqfv2UhqkAhRxBSNFri7OKmR0NB74/vFMUtKboUYQJSAt11gkeCtHMvb3IH
5MpHGF5vP4guAcUq9nKxVMWrGu3g37Ogpd5jDUsXHPJrXIZYPIFthHiv4+82Kn24
rE3bOR9D7CudIgX/I9XeIfImtBiBwda/WkBap9cmCbY98bI34pwYm43UPL5U4Gsd
IBf+eMXnadpx+De7NK1odtYR1WiAnBssCuF/z2Vnl3Y1FteQmZPHqJ6dyPspKW/w
mjFBW8hqahPLPYI3zur2dWW+aF46CYtLtD5Z7UqdVG79xeasVyScxnKmWlbUzwlD
MNp4v6maFbJtb1NKWp03pDRtoXh/q9jD5lbLcZ6EmVmVD+eMOBCeD3nUwBM+w2M8
od5qkRhlBVImizGZNeNxrCNBI3lW8LlHqpQXOmCjJNuKdlsiu6oXRFRWwzUUfT1W
Ts9vNTSgVfbm1jFvfaMWHzIqqfaADyVFLwiE0Wo0EereUY67bHpoX4qhjmOAY/Yg
Lb6AymC9Nv1Tz5VNR+vbRHFPGxPec+e2k2PPVoXIjp0KOBvW9Cw/qFY64tHPmv9S
PDGBhScbEPjhypVCJzGT8OeUZgm+Mx/E75DSm4uSFJpadlj3ygGzVmWxZsUiMMUm
cR0rDyiooGyA8ZpGM+nB87YfNNJlDxay/PCEt92NRFYKODZYF4YaRb21VgnqaBme
smfrGV679BO2rtYkHYzq8EJlETRfg9IR4X1Scy1dTPUsHqdsBwUxQgxVpsfUfd5X
FmMVLF2kqa6qqV3BzKRDtBPyT4oaFeKGA5sktblK4jlg0fOGCHlXuQmyqdUr/YGI
xYbt8x/KuNd+9zOWLbf1+JUnyNeAXkzeBcp587f0FFWw/JCH6YP18uM6HA/5s3xT
tM2O0irCqRdx4oSxePwaayuIGR1HhHRbP91X00GJm/RDsVkddi/zuP5B96wfi5VI
rOHmrnGw4RE4T13ktAF57Oq3m04WzphTeqHK3ORZDAZlBUIjM6il3SOgNQgZ18t2
1DZFkv6fsrZnfJpdwFb8/FStchM/67Zf2B1i6ODr5PuPkGyKGDak3kiEPDlDBZUS
lpyLaS6BkiP1CRnccmJJHsZsTP8LnWogrphxJvsEnSgsNFVNrojF9jm+q7fIrhUR
8YKFpPiZKG1tRLaXz5/wp8DHY3t1+aCkhrDjO4+zcPv2NvXEtIuJVfpsrZWYQRmb
tUPUWWDhWpjpQ5PHu3AP+xyHR6aDsdcCtfEktOuexV4vg6t0pP1Peu1g8PZLeBaj
JDS8SUIu2IWQluD0bqwnREqvAPg9vECYB6McTa/6jQO7AqonhK+DBYv/ePKBwiCN
bMqZjftL1R8iJMX4wLN3hZ/l3mjTdC7dqFrpM5hF6cEnoIPx7v494+LS+jtiE392
PnwamLh/xUKJ20JJQaNUQpPvy5kmJS9t6e6K2gMoacX0plbN7/ixgWKU6frTNFoy
da22nmWLnudCct9tX9vpMlbBmO9nXrblezfpf9zbD/EbKfNdWs7CSltZWu1Fc8qo
tBj4EUfLUXI6L/7MwNsNQu+DAmCdBmJ64bj9YjOLIQMJv82T1Y26ANNqydw8fvmj
GDlFlBFot1iyHSfJN0IPDw5NmAYeiAwfNC6ekZ1xY+7xRSdYEhNGKabj/OMIw44j
DQqzwH4tWHz0byNCgdlL5fWCSu6ect3G49CZ8XS2ABYuq/5Kc5IUVqpZDeEPiQVA
AS6udK0/PWHzb/JhuN7KDfsnR7ijsXmPlYFM+eYy9q6Sfah2xPXDLnLOffPiJwoK
54nKSeKNxeuLluffGHBjOJu987Tbyaeb6w3UgdVNdRhXtnqvhpfKDaLBztsh7yuy
um/0XZaH47gx/rdxjVjGvIYiyntfl9oeu+eSCp4fee91btsffvxeMswIFav+80OK
+JP1iS512AgtolaUGA9AW3Jj/jsfjn0DxAygkTu5kQ0iLTBKWJpfvK8NsXZmvStc
jSUIO0x4f/XMRYn0p8anoyBD4QaB9PzRVKJajgdfaFjn4Oy3pnfjaiylkmbZ9cf/
2SRyHSTbbQDtblGvcGy6BgouFf/bxcp3ghHLA8RgbVOmBDn1ozN0SaHRnvystYTa
4biDZzJxWwqqe755N2JXaUHqx1GLogz3JWqK9C1iEJ9kQj0x48aeJh6k8ssWPXFn
5j1gldKkoWRw17NP2dOEg2fm+209au8OKKcikjIxso16rFkEtizAyq+LK0mo8MLs
O+qRBlh+YhjHqcXRl0I+v1fwR3A+InpJINYp61DTNtWUxKgW7xKPYB+c1yjIEZpo
UZVEQRvgroRK6WCfNdDOAgY5hu26Jj8xMmnmm1tTO1HPQUdu0b9SxSR9A0GBXRUG
KY56P4tidLfjXlK1A87hwPDdzLxTjzhLbLrFYz6RB7MMlIJ39Lqis9/HL1F8gNI1
i6jpcPDScoIE0l/O+Uxcoc1rW7vY/vUF+lxUqEPd/HFGbXNEOjkophn0xoz7Pjf5
sJ5+LMiq9lWsf39webR2vHFH+kEq74dei8h0LKjIMPxtnRcDr0Akot68Cb+oKqdE
IBXV2PYQHGLQg1+a4FlY0abQSpPRSdHVkrP8eUau0BwBC50LedTQX+txslhXK3XN
6et7pTyievBiPot6tg9aOfiDQSNVplRAcxN3gGj7uUp9cpfj8to6pVartZC7jOjo
J6dvqucKBPi6Z7J/C+TXLmRg1NFpBRgMKNOvhJiPtcvA0QX95W7IGMaoUxibS6Rc
wxCk08Jo09Cdo1MRNBebaBYkUnbvzzvCFnuilBJWKIF3YP8AblDzGE+Lpjqiev5G
2d4Q0iLa655HAGqa04HWMUxp/+rsKpfh5oPEHvWqop6DLDTZ0Mw2sfCdhgIlNY2c
2r5cJrIiOGObjRsYyzn82uGFjZ1kRls3KIo/cLxWhHR58W7ndcFop3CeDt0K2wQy
TG2fSKOy+2KRKdDS8+ON3a/HmYFwCavuHGehlvJT5ppJ3KoKeWqjnCM9QBqvm7uR
Ybi8RR97kKAgcMVcjZGpoh9OOpHBD7BbkR8cq9rqL5+CfU30tJ5ugLg+7FtGqSRL
K6TqDAwYuSrhRrs9Q7Ap3k9mLlfg2FU1Qtn4S0Yw/VG4RBLFWMzwOKjTyk/ePDV1
sur/e0f+fcHodQzcVcX4y8S/ZnHX+PqTrh83wGCuMaNOv6XzPl3CYG24nzwODfvY
Qlzr6FBD/vuUXCQ5nLdMuObUJ4ku87NZdGAFj+607nhZPpDpg64RJzAb6Zr6lyZp
mgjICX2H3xyhweuQ6psvPBR9VTB+MGym2rjcGoitj6Wn337OHxNfyG7/ZWehgkoH
lWARWRJlIwL0dIwT+nHfzaT5DwAbhanDcIRsqqpEeW3WYFVh7SXRarEErb0tmd2R
y16ayYqM2DkNyVornRn1fa6tdIN6K/+mq6IDYDKa/xcDrCaFzr229ySvGzmrpUU1
eiLrs1cznbrhc1x1numgGathS5B7V52gSjw7Jn3ITwC285Mx/7AhFGl5QybqhL+z
2AyV+6/IeqI4zD4lSI9gXc2QfUHZb4rp/hoYXfuuYUnb5uWov9v5vpSPcZwVzukc
ohItj6phmCTiF4xExlIhMS7LaeKtYOucQwB4JkMk9mbOKZD2D3Stkg+g6IgQBU8y
AocHriESMP+yfkQmR+kQxZCdIuV4mVMOvixNi4xakPpQXNMypYF2gyZtEfmSgNkB
CTS/BOzfTgOrsfRIiBTQlovyG+nDZO8MfxcjkNlJs+Z5tF9/OL+KJw/sHoK21Cd2
jpxAvP5cJpmre/b9BuETGzcAWcV+XD/Wm4CaqDQ4jVWlBr0kPcGhDrSkMarRIqhi
koh1W6Kzsec308KsiCuNd85SWjQHiWAMASiCmS+SUrQBuGmRYMyDQ/R2knpq5bHB
fmUbVOVpcHEyTezoZdZuQMDlE3fIechP2JuFBNSsIulwgyXxcB7jKCLq94F7+rbp
cnSJ7yVJL4+KO4tSSregMzavTv4UTaqKpT3x1r4/X3eO0vOY1fexTkwEAH8hiX+j
JwlIrnoVk7EcDKjDWCU7wjA4fUKwE3iVBLfUo1Lv9CGNjjfJjRrp9rsPJxdNRIjb
geDjQAlaofBf9ZpKPQzx25qav4MCbxS6SBZQ6Q1tTk6FzMv6+6d9GoSpUFKpSWfD
ln2ufa4DRwmX4AvQ3fG+FBMpbCn0fKUVzKffeBzlcrbv87uNQ+5ONgFhsIALL4Lw
KwhcTbaEV+tejKxenlvZnVFV5V3GnHCxyLn1j+B/nQtk8GsdzJQUHM6koHJAktmI
gQpX9wyGnQQjeoSegCjmVZq4dyi9o98/5fAMexLf9LUSize9AUhgKDtO/uUZju/c
BOeYh5pEgwrXl6KSWMYVbtXJVOsL19yabrKHUnhelOqBZKvSEubuObqdJKnNwZ60
bqSuz2OyGsECT++rsld+DGIJPZckI6Br4W7KpxEDRMfMgHNpbnf96wayHTvHZ3oa
aslIYSSQ9nNtGUVQ5qOTWiUh50Hfbvf/GTBqFCSab21QPEkQEDObxgYlXIoYTp4T
NU9IhWo4RxM967LnTNcgYJr3fL5uAjkiT5gY8+Dh/6HLH1YR/mfeLx1PezajBn4n
hzV3bVFpFe6GjHFeXHVdCwPMwJ8GSbvigoGomZwut06lj56TEdm40/WtLwLhntJP
910/iYD3LmwRfjGzCX9n+rH27GZGXZjNmTttodYi7lYMZYGU3np6GWtcq0KcetRc
/ZofMRUiMnASmvbR7QEFMh6/nxUSMFFhAYYfKIS2uneiB8vlDeKMNJd+NXsuU/kA
tg6ujCtSCARnx5Q+DjbCh0ZEt1nRu7unVK4jiX/xdhdPlu9wHqgVb7Vh7JrlQCQM
YyqjdrSwb7F20JYX7m+b1lCKkiWueK/eU1da4iXdE0eGn8VNzL8H+HbikJaQXs13
YWZC7ugKK8JYfe4h+1y3CPhBvK5nXb3BhagmTjr2pSS56NckjEEHAX//lMr/XyOl
sY2AK8AFTSQ9JV9ThJtmknfx5yyxpd/M0B+XrqAK1/RCpyY1yHY6OpRaB9OeH1rF
xrKdJrN6ve4RTuphLuEMw6mYPo9PnO2bFEIOa8dlw0ICwkOgwLbifIFhYkYc2DH8
pZDM4hms0J09osVFGFphHz+RdKwHN9HY92dMmVD9atUujqOq7HQveVjv99MVP7ao
ydRJp2J8QB7z9QtOkHuJ8jz/Yj2hKhSZDGfhUsysAs50dV0NkuZEd3b1e2ZT49hv
AhXlVpHzSAKQvFvLOyZIgTETDNBL79A6YOr9v2+ThOjHViEYohNsLciPQQ6DbTjk
EgVEd4SLcMddlKiBB+DaJcRPPfN8QUU50FFnR7tmxDZb9qMi7jEAcBPE+4u0R71A
RD6fUkkCxx/rOrrDpGsc/spLOf94nlJI8GUJWl+ZT0JKc1lSet0384l6KgpmLDDm
SJ1wl1Wvjh+vRW8cuUx4i0NUfvsdQ5a1HS8NPADvs1AmeR4ql+76VHbaRq56rys+
7/6+fr7sbkwJ+booBkCAW/5vVwWxCMA8E4sFH5iCiBzEE2LMNkIfxxDFZp+VAR7K
VMjvgNtfAMPzXDS8ZSHQwybkrp1bf68XbsjaEmWBOhLS8qgT62g7WwWFlcbNC18n
h+M3sa5rlYlnzHhqB0p0MbmetoQE1Vd/Jb6qKF4x3IaWhYXv3IA/3luXjFzL77J8
RPnPz5Rgw8kKREYJQF7o/FYRjrO2Gh/U14yKXw4eTaXU7Ee7fDB95lGOlSPiHOgi
+SikywqoRX5jbR0fsW85Oahfvp4OPROlKsGNFq34XdQ4bUtTlZgxQMQi9iyM8YEC
McAGNg5/mzp3NT84i/NA86WHPepuSLpT2okqyQJJF1wiN7++r6n0ra/oFudeVF9B
mZeK6/VDKdOmQpnooKyMLFFlVns32hSzDxll4aXa8ErqCwxGcGw4eJ/26iSdd1+4
xYuWxzXjFeWItqkxbAtXujrcZP26narKI9SZDlvySwF1wGZLQQQrgsMhtM5tRj5g
UV5ZwDJn6S6Nb0bBBGIMIquaP3sXINX7jvIIdwLQMLiqL63mHaGnFNzoDwDS5G6i
uh8cOYLRAvYEk2drEWYJV4qZnvgLHNMNAYmq1iWu6AzRj3atqaX5laEuKTXl8VhV
VqKfgbTuLKoZimL2aX8QyL1zbYXjMvPZ8z9AW3RZxlyFGADRS6IHt5UH4RQ8VicT
G0pK7MF1e60OXduujlLQrelbwSEKm6gARicVWeaw32meK/YVs9GcD6wmOEqaNH9B
NnqSIcxwllyQQC6knnBISPulRg/3F4AXLizB4QEQRWkP3xgNK0/AAClNW1RIbm4v
IL64ZYInl3zFsPU9NT/tOyirPmH33fZvCFw/2SYolwbORi04WHIKzQ7Sz56R3KNF
ZbQWYrOXuhObV8Wq93KgksMqTIL33c0eSpteF4PQGXYdxbJeCJKLpHN0fksVZw4S
5w7HbWAh9JM9FLGC74nvdTAw9cGZiB2OxiyySRCRpKbwolyOEp/VAJHRyysCnGIO
2QYfE+YSug2vqJxV7+VmPSC8F8QWLqNBLEKSFiD4vIRSDwm5d7Zsmrs8cRZKnBGB
5Aixb9jzgRA+04okQAdZDtIQDugk83cmCKBiMDpSyBNK0hhrTn0rb0UB5YaVD0Tj
TO3qa1inzp6X2yc9Qe/liaC30WCoi6CPZYsggJH4RXm2SegkefHYNKbm9zm+s1TI
wr5l/+TSVraF1/Fu4X8MMt7R05Quw71liewsN9OlSnfkRrUgzP6zqeXg00xntPqS
hl2lrqVVIJpIjthB0AQjO0ZQ1xwHIlmYMCUAKLz686Y6knpZEAZUP0BChkhfT9e3
qqYXqAfLdIcLxRfXwsW6IuvN8ceURD/pqQD0QDaVMXUe8UeEpJWNJogIuCtnJDjU
pdOYkNmoxr3b7nf/jXB/9sbXzwv/G5Y0We5U+E3YD8VefL1ixjZ257VHsPKfwBI3
mqIti7h8NNWUo/7ZlOcspqPMUIloWIesyDrLInVB0kw2xBy7mDL8JGftY5hY1EGu
hwBXL3umh2fKWdL6VBKlIlp9ts16CRWe6yxMQ3VwqSmWXMsJEdE8snsnGl1oP7Je
Rwnw7YkJopy++k0zuOUmKEmFtrwztSvEmHPKPYtL9CiHYczExp0WH5mv7WOB92H8
5C89ysredHAuX6eZx+0A9M8BPVSqWnTiYMX0FXLn/NgmWVn8ZpqXJhNISeiNB4oT
kVZlvlg0Irb+n5K//2TFhtqUFv58/JBy7p/ZUaN6UTTM6lw69gBJbgyO0gUW2ntc
QCSqX8M8BvYwVatNQvKkvNvlqoBMlUVmrFkMQXcrXLreRsnpP4w5acMhmiX/hnEx
ki37e42savrniPIXQyXMqpdYGYMzkz3LYYlOl0HmvLeM/ohh+qVAmuUIksq/fEME
vdAV8XzN3bYTxJ4hfugK8o8uPL7AofJR6PBEFdgJDModP7tlYKgWm3jzK0gEPmBr
nDHJwKNeaJS/xt4otwE8X1fEosIhDApIBKF5yRx9yjXJw5oeppRXuFp6elOKAt8V
Rlbl/IYk9Vkalf/64PYmJoSYf8WSvvqcd4y6D4r4sg8S0Xyl0JrZ4+xoEDMbY4Ao
K/xGuU/CDr2/txwWFCkJc8S2zMXV/URqFBR5Oic4bueX6Lww4RTEfpDlwvpV+O+L
xX94YOiDZWo+OZXqfFEYCgrea0R20oSNNi6b93jxBK7qG2vnD8dIlFZjU0JKiGVk
40QwQYGObtcAdYGrSjSeL3VHW0qEc80yucBvRH4kng19me603Mmv+pmmUWTGRvFF
yvtida/I/7m/vpjO1zd+O+EkCqpP23a2jtL9itDoIpWw7/hYzZ1HZujRvDIogW1r
3JFe2cxVNTXhyJJ9LbJzrEnmaD9Flkk1I3Z5pElwRtpklocfg7/Mtqj6qpwDNfiB
c3A95X4e68jECLPlu4r/N7mYiorVUGs7pVImwcpcdXH4L9lStv2r+jQU8juwUWDg
3ZsIikwc/9uzC3xd6b6QDAbKP9FzyqhYEOn0aXJ1ufG5aK60QFwnl0WOtr8Ua7Py
Rcd+P0BNdYhmVYA7gP660VDDNsG3FR1F61jCwNpE8FDt21zzxI4hqqhop+rpKPbL
fhvB7Lm4QKR/Es5IW1StRrnx4UZ4Y8E6D5YBnuazfM/LC+xKof1ZoTg1/8G0JlQd
6omQTMIvJc/9QyDYGHUa8sbnfs8cikPS9gm1QvIptrrnMLEGj3qw1bW/dTFL0eEc
UCbUoX0d32hRarUCpDEeeBoDm8nubaGsEoD+ubhgBxtISg41uPMHDQqD5l8c2u6z
GhnhMB1k+dm3HOalaVXOHNRhE5Qp2jYtBIkUdt5iFFXXX92qvqEnvNYexNQ6A/y0
0Bx3W3E8P1HUUKwJgdQ/CaG1uoDM0G111yqcuvEA7Pa2/RRHkrITOk82lqRDRV3f
fw3zwyjOt1tULy9NcI6RMAneXclwjI5DGqQqZyY8luAQto5vl2cPONQKnknCiQ4v
HXKCKGM/qfsOUmfxcmOjv/4PnxX2c50LAkVNGlxNNJdP3C1I9VyAGJQ57LmsrdGU
xl+9+RDSq7Kdmrraq7Z9i+lbjTYJ0576kQqOVTjM+4ab+rZhvxsDUROZAtaM+zV2
rwzAt4Zkcg8rhR4f7WieA/2v7wCxOguqWboy05OpMJn84Fbfv28XquZLvZap7/8B
HHwMP4DAr4iTsLeFd1AZJ2pyTlIxUy+OMMyNTnBmtUx1vbjToDwi3cBC/b2mldjL
ctiib6LBf9NAg4j58FNnLHYfXATPm2Gd1Wy1fg+vRUadzGbC5CZR+Hsbyp10H7yM
A+rwV4tUteYQ7mizu0O9BjrdT4y5uYHsUnSuGYdCfWOf3LtPLh7YazhAPF4tNZ04
9tZXgBFptPkESh6nFZlm1LllHC0hmP5cYhshNgbHxdoKH6+6ftvosvsjOG/ia2NV
PlMGO22FvMup+TixPgVMQl/M3tvx64US1UuypmSNSqSf/ARgwRhggIf0bezAOz+1
VT/o3k5ZXI9IXL7azuaf2kBUq5L+J9B+jCHvITPe9fQ+jyOLF79OEZbaLrKMw12T
JGRFHvwTvkO1bhNpIgSYZ3jBtrW6QfB3tLlLiULVffMvineGKnemMnu39avdM7Cp
PisslaHj24dNSkFtvmOEf57k9zN1zgBoA4yG10HZ8S7buzZnYeFWLWh/eQITDsRJ
mL2ra9+Jle2hPzh6mkhkpNqL8qO0NJ1mmClzJbOuimD5MtpmL1uon2wcqWLSof3V
nnnf0Of0/mWUs3L49ymXKLX1rcx8CRAExJhHt/uPU9HO+IciQfhpUcWvsiyLDtff
FRaoOtKKW4N7wSrt9jDZc4+2Qn0iVgm/f/kzpdPQ3zgV2spXq9FiX7Fumn/SQDby
Qgj4ot7nuqgNDD8vZjIHaVU44PUGa6S/5fpqvR5m+UruAyjL959nVYMAfnQFNcXO
PLd3VKDliZPHcHqqIoWzX3rKePWuSjTD+bvDVT1QOlHXEdnUHp3J43r5HPiy24nZ
JuZ2navL/BafpsePIgxMMlDHPwLQfBbs9zbJS3KZN8flMdadiXhB0vEZjiwjqbMj
Eaxha119YBH6nzDJWyYN+byO2nqzhwS+AGvus3qMvdxs6DVQqHz4lR2QSDwOrBrI
0T97Ev6tM6MDLQrT90iqnwdDFbGSmznHaoTZ1ME7LuUyX+CpR7VhH/aC4Iljwifa
gA+mDeYX2830RWKlcFhyu/N+MvFY04WAjcejAJFlWM1t2lK2qBppvx3XPic/RNNo
biyGM+yohjvCMh22f9JaGdSelxWqk7jMOGIWUkuFQUl8lKmI8ernvploAmwQpZDH
uUg+fw6uEkKWGxyUpHhKYfgJhGjd4t//Y+VaXA5DnN2kV7zC9d0Fup2zldU5g8Kx
CHDMc+RJcSylWBeeDLxBVkT9s/YKsIypQa7J4dPNTkSTr+d7Z+tkgSVMgvnC+GRV
z6e1TJPgJiUOlfqr3FXCIjApvMAd7ohDgaEUj5Nwh7GZHHxfCKFGn7s0jAOb/4Yg
vvN8GUIr7YBlo+/J5vnsh2oB1XIBtw+mkQJU6Ggy5MxncD0aE18SyQE+s8fh9m4Q
PP76EY0PekHqKLAEo8XaY7nzpIs1HlEv/xgBYHqybql1/kIOcwetBfbTt3XeqIHV
kA6xpWu+kk4ZFnfF53mrvcn+cYdZ+i+sICGhf3LW1xrUJNYk1crJWfKlWJiJ4P3K
0ZN78+Vf57EL1noer4oMWkE44skwrgshMQqk59T+97W67fjpiDcR6OX0XI/Q4Z6R
xOedhj8y0D2Dv7mvPV+ImGv4QYdV/Jf4Yup/bAruMei3WrsW8rE4clVCBEuivHUt
3iS9NqffysSZ/p8G5EasXrAc/i4gay/Znfdc/pQIARDsi+vxU0AVQZpQzM7HBsiO
l4bjgZkxVpoLbSCA/gsyqvBkDqr3ZuKQDbJDYJWhHGfop4QMfDQVbNhmo7yIRPKt
RZ/AuA5FlJ0ig6CjXfjpD4+siU1T8g53S8aDXP5CENmWO5n96ipV88hi9B5ZhaZL
2vJ+pfFcR/vp3ALg/DQgmMLoBu1YUp5abX34JDvWPr2bICtGqEzBYPmcjr83eWFt
gaNmalxgm+QTBLjIHP1ybx8V5YRkQzwmzaol2jhDd60ASqCcXfpF066KkDQM36jv
RnR0f5m4SLQDZ/UNX9SZXLVAlj9jutvu35nNqFmCDlCRZb70g5f5fGqVwOCv8YQ+
baO/F6qXinqZTD54gPpXvpDPRl8WoTtRbhN4fgJzyil9jecFkiY+HxMVMeUb8o8i
4rxihsRZhTfPHXyjEltC+XvIhCSGDjk4faeOKSuD+7MD440h12haNUqv3Hj0NFuI
ixkZQrYa1Pq4xbW0axXa5U/ZBFpYP+4MRBT5Rj+STtpVil0b9DszJBW0Jxhm4eMr
gP86QEYVXOlCeMxSQEtHUhidCjTNpj37ZOw70/UbI5xuGjqQnglRK2TKWE9cfuaR
Ub9doGC4NhQ2TpI3/YeMaiN6uSmv2Ucwgv7//kyK5GJHop8gBcCDl5DmRYj0hdLt
L3cIZifpj4sF1XOsvJMxtcqxeQ2fjL2xojut+6/aRCoLzWYvMaJd4fXkQKK0Ho1s
2zjVWrSaLTR56K91y7JCx1V4Hik88MW6qLaVckp/EhyMR4FznlcS17pqjGAc1lg7
seLjnpLcWncI9CiybIJliEoECYu7LV7Y3UaglBdHaTUS+x+L+fi+kqyEs5A23JSP
twff2vqQ/o30SVHx7UN/vpn/6zY8tmU9q69hfCCMbRYMWFtz5GehWjiJ7+AWrSZW
WWjPjNZAcI7CFRYX5dVutT85WLFLxLXo9DOrlFW9KbRMSTVgovdstkVJJvcw0dZC
5QOrOoKaAV8FO87XrEN7LldPUgZl4HDVmzGdf1BLxXW1et0u+UjlCOss9UMdFRHj
XxEQdTUSHcci4liBsWVZyW+Vpdk6Nx24X8G9wkY948tvOjb5QyGbaL/bH2pPWHmw
11m0PEkuHMQT6dYTmvoDKfhKdBlOJ0tIUdA9/nt5YyxlkXiJCMiV6oUP6dm5OPpC
J51qi/TZooftCfCkixqQbO9kkvX/BtpuRLnSjGP/k5CrViVDqpvCzkYKAw6H1A4h
KRbHEPa4TneFwpxUtYMDlqN6OhOzG/4+2ZBsDT9f9+1QsEFNoKsLcCXcbNQBISAo
1vCalBzsoP18X/T6fOfhhpRSgjRddbjLJuyhlUZ6dMN79ELNs0MXmXtW3yuWEnft
vGCcPDwUu14TwDnuNi9ZgB4/dQA4hyoE3rlIiSXYpNQmAAIP/GSG1ZfD/7SBAQRX
nYvukcWMNkCBFeMLvnwXthPpQXKnwthzuEbhDtfL6rm2aTBJ0BboqNeAtyAJS37D
afrP+72UubIDBcN37/TfNc0KgbZXlLDsbJsAExcc7QP+UBgu603iiL4jfZ4G3Lii
O3xn3YsFX7VPJ9gaY+/glpSiLSARYe3YBmDoaPJoHjghpwtBzImS4Q/QxI46i13w
VtEDhRDdog/0+7k97KhzhmZNoQq6CIeNFThQ5ZdM+ADASjHBFn6zztUIr4CIA9ii
hT2pVZhP+dq5m++DcxozyOTaCc1PvQYDYCiB1ELgt2nTaqytoUdSz7jhj7eDvwkT
G4Pt4F0l6BfZEEhI1XY2z6O3UdiXhJKASG2E4OfzzJ9+mXdGRUdalJ+IQfhdYz/I
KyYBy7l9nSOnoPmqgLUvi/YxjKKpeuf6cWc9w3/rFAEpGWCK4V5od+VkPU+VztdB
z8WbJu0+tUhAgAnaV2wO5Jxnhgz14IQlGkgaMt2mt3C1X+NvvgSIFAA9oDMlV/Re
9gLGtsm5v+4tFi4LwQgk+dyhnpgwtsgjnrnXzBWL8EsbSzZYS6SWhtaVlLelJSbI
6qyVNjF6zPkY6VDZ7rDSAwvq3n9+9+9Q4OuhzAdWH3RmNH2cGqGk0YAJqK04w0IT
PpTozy2Wc9N5aZA/dgINSeVKRHaOZTL5J0PX+QduXLj5RIFGKSRMMRk0EmWTSwOT
5e7YQBNc6RDMpUmpO+umyAQ6BafD8g5MEk+Ixo5qTqD+d7ysLvvLb/NspSerFyBK
aRNUtBfvJHPO6bdF8W4W4XBFJfs5vqXlRjaIx9ZkxWZgnC6ROsca7i2s3eV9WJdp
e+wK7IDVTI78ImTJ1EoxJlXjJbJULFfpDh4Io7bPu2lmj6sbOah5rZKNK8lbplBq
GA4ohfv9brb2kTQhPGB0TSvf057ZZzNVO4Tcs8XXWjg/DqGOqKDsX5LZHKcz0bVv
CUEN+6x5c8/3vN+pE7ojir2juuVLRY0u739PCQTnP2kWY9pYCpGLvuzUNZoF0iSg
/Jk3lh9Re/aHGHEH8rlWNS7BStxnDfHcjup6wLwbiBZG8PHzvmQDKl83PcC8oPsM
qCMxxHR8XTbykXtK/bknwg5SO9Phs8rwBIOo9vMwj/XJ6qfGXs7ShQ4flesjPPWd
TqajAXbVkxOv+RueSggmZXnJBklD3iEzZTSmpXjNEaHEwJeSiBbVeid/zbXHbf2w
G0wgi1909LeqKRZKKrUaEN4StpwmF2nvM0BinDkulhDWNbGKmOGYNhdPwsFY3FsC
UFDe0pjSb1Q6ePreHHyNARRxNvD9Da2rcgi1P9kK2O41Odap8pQI/XCg8a2vXNue
qDG1eA6n+Noy798RKdenL8T4NfLhoq4ES0I/MjQFaxeqEMrNaITA0efeVnl9sJ1L
Eu5VK0X8aeqmQlRbgizPWh2qQJqiDdDtKzPzASXUthjlMMtGfec3qIRKcMhCq7eu
omCyYDWtdm4I7AJUP9K4wyKeHgXSXb0kR9IjZMcVNchyoPtkF6iAxkUO/J9nXTjw
/cabIVrBOCU8znqXokWkDUnO+UBX5CnTj67xFBuaTQxR/qqXzdRul5ed9NxKowsF
6KtIv2wYAtHyPa23RqT9fzOXgc0bMjdA5P/pLVS6HXpI69lQ33rZr/8zgsx3cAg+
1TjAJhNNxzxbVquqQEfdlfMhj6iXaUWJH2kzfAs6BVe4jlpvZ6/Hof6qP27rreWf
NluqYFSdo9nsGzzC2Cy5luLH7uHgeWmjOyzAa+xJ0Waixwpdpm2lCj3gtwniT/G/
XywKZBMW8pGF/36d2VbAqceYpVo2QLOCF357qn0DILmkN+3nPZ7sTTgTNHMh+GZT
XLWyOGZUIh1IkmhknNzf56O5Gq3a8hfLJWoax38xsSHJZY5t8OrIuyP7PpNi7ANW
bVq75C7E9Ct4oKexKDu0bvp7cy+ksRY9kXzXEWUfrTvvm9lzjaEa2SsefNY+gUHN
N2c2b71vrf1O2SZ7ueXV8LhC5YddDsL9XHscn+nvGSfdyiniu2uCMBDGXJo0kigD
8FCbfVzliumVWCSyYMCOYN/KIJ8h+2KQufVt37QhZpp531RVWHgmzizfFAiGa2a0
EL9SRQCDShZQQ4iRMX77j2ZGD/CtHLmj/q9Xnl4c8J2D1S4hnvA3nUazfjVgsSo/
pfXbZuc+2dS4yB2S9LJ30UQxpYYtQIY+tHAIkURuYmtmzatOtVibPINnmfTMAA+1
v2tmctsj2UszuaRL4LfnI2Y2PDb4WhWngIY0UlOroua/0g8/ASTgyMstfCZQV0gw
sRmQ2SLkb1Yv93zKzwutXfqAaEFzBMHU9KsD6LvyIW+GGy3jvJm7tBJFJv58/3z0
XwPLIhHPXPf1E0lCkAcug+SjSKLARvMw6OKs/bFMhkyh0xYSwZTRIdLabYgWkCkF
XD+8x4m9TR4wM64FYvyv/o9XPfRNqZAnJnle7V/GHduVQn6F2nAe5GkFCtYLVFLV
oqn4DzfEs7aEnMQeAryICp9urYgUAnt3KH1ZQB1gHh5U1fiTF/wockLWAT/kjQQr
4p2IDQ4eNY7inW6zCy3igHITmhd9SYCnytRdVAEUo6i80iuoNNYmQAwwC/sZv4oT
hyaWu+jU7cm/urG80Z0hytulggDTxcK1v2C4kaCByLe02mFB8Uy+y/QgQUseD6D3
+n4rgvU07X9RSohjjSIoM81tsyQihkMPvJlEcSV4zUnlzfIkPqxNwWmIviB41csW
YkVdKshLbMXYDgsIn5Whca7ZwHj8/LDiQVybeGlcZoHtHAIMihtcaVJWuZxjqW7B
KwUCG1632a2Ha78esq6+4sTJgbtvLYKQX/YD2j+fUJtBzIQ+YGkOvl4VL7hsv9vE
EGTE1oyC3sEgtAzwIdJ+DwTUoqL0f05fQeS+3nGWOqiMFGaWmQZeBEEkut/qLrga
bMY7Dr5cHcvTyi24XyZmkFyRlcr4vJmuCjb3f+se4Zwm0nx0pECMXphrI3brrw2X
BK01q6UQBQsgkXvxQQIzRm69Ho0q9BJRc5KDs5IZUrp8sOObB9JB6ds6AgY7uSGA
HhaYSlgHWLe1EcjQCkXj7VAnaBPPKAiLcZ0KkDUP4oTuUa+DG+awGa7I3RJX7BQD
R81WO7+2ywXaRSumeYfegB7kQmyz1T5iWxYgd8fHQzBEGUMcOMnIF6jqzE9mhbof
lTZ8TqOd8ND5nOUQVBPoNjWHFHsE5udSnIgEmWX12sHNdXECOY3XvB4lzQHIxa3f
wN+lInAmgtD91L/pPZAtFgxbTGotvrLa1ywp2PyDjA3bJYjnAtbjJ8MElKSLs3iN
JBh8p+RAJJyj/TrGVIzTm8fzY/qg+DzR2qbal89JiwAmD2LtHEz1Rhpb+DK5eY7J
72P62b+f8KNIe/O8BOZPT+B1K7Y2Zz2tDfEgdJyrUmNrEbf+3MsZNJviP7tiFTPp
NTBLYyX/YqHqTKlvzgpHN/0VFErg9U1b8jiU0zCckwI3Bn/P/RQz+hhAVxbZvKT5
vUpYtymsaxDIln5bk8R+RjG5Eao0ALLMyvnULR4ZGsisEKmKQMIJrR9/Ddtr0TfG
mTAQZIWlLeN/OxyGfzCo9nrBkH5mqiisR1MyuUGQ3YYctizrloyW0FrSd5MBPUVs
QU8d6C3xogbV/1Q6XzVK2oJOW8E8mVDxfS8VSzLm/dTAYbZA5+V7aHCzhZJcccRH
uI4V56wcMkQbS5N3pQ3Y35TCl3w7RDiOX73P2wEe3IWdWyjDZHfZgUTMWkx/DoOl
RFJXNOZUuSfUre6mUJsGZTaps8v8cJ0Co1iCfbufMKM+/rK3b9UVAUWn1AV5izuY
A4Bar7M+k8Nes4QVnBE5PQg4SEPS/IBTNuHXGmfCp/hIkc8yXnQmsprLlQlqkmBO
zjKPGDhrlfwQuVAh/5I+stcIRc4cxJH2cx7uSzwgm/Zz12Aa1hoqMG4zn4tjJ5Cp
xShEjl3kgpd+3JuydKvTRDpkXUWIn1wv/TUMpDrEg6nDyFTLG0Dgj7bEXbspfsT4
WEnOL0tTvWmy2OkJhbXsi7FfVa2tC/Gv5fPGyiRGQJYzGCYJEBppmy3jpFvP+Crj
qBZ1XYKOhN9F4TnhFveGs8YoNrlV9u2/tncHcwqA+BfIvHKPVJZbAPS6TTvUtq4S
u4Vs+cO1+JcxZr6sID0g5b79vowDMAtqZ9qULUFbFlPADvTaSL3QhIq8zw6qC+D7
QVMqfP0/egpRU0hJs2AcmYXYMGLZ7qtXZoHRlEl4T0cpAmz1CzSxAUc2MqtLzYt6
rkNPPXlKcqR54W6QpC6L3Xtqv4DMHKoeT9OCgkxqand/A8BFYzoSlaP0iAFc2EVg
k/6yc52ckSb+JGluKeCMJbKkZ57ZL5vPMPDt0HYczbO3dBEycJNEhrh1e3l4qWSW
9S9i0iSMmieMOfyW1kjk8nki+mIgORtT/gL5+BixnmIf+6wNqjnkpgJdhCZtK5At
3xnUhcyyApZ68AwUmaq2gOCxCkAt0myhjFF3EeydysaD9FDMzmZGI9SEtkqQkcv7
Rs6hzsIKAH5B0P0BKFD6w33b748gp0cZmVHcV5ePC1GXrspacfAAy38ccwc35wIq
vU/YsR9mLvI844xf3UmnjYDhwaZtqbhwTrKPPqNDEUq3m64RcBGaziQlgoIFCipr
dfp178jxDiJUf5Ji/bNunzPQfywEsGDom2+ZVLyYJfbn5QqmkJ3J6LnzqyluX0bA
fZvh8J9k7h7jCAPyjST1N+E+kU91cUasL+0PZvXPuoNc0g6CwkpeUPLaex+pKeut
Td268JtCj++TsDhd4SnXuq8Dzw26a37FyZsd5m24UsJe7zKCdbdzx0DJpTSt+/Sb
kKpVntar6qCEsH4ZiKCSPXZt0mmFx0aU1cRipMofIcmFVUC/guN/uLl3UoReEe/6
cxQbOBpIDKpTPdRe2cv8r0t77Tmci8N16dOQfPqVVtViyZ6+ZvqnMNWf/5taGJc6
RXaQwuyUJOTlN38/Nd1BFpdDTMxDtvXGbswK/BfbJJGdNZr0u3vGey5gEzyPdVJH
BbSGLbGSlddmVWbj9NihpLOKbg7FZDIkQuEdGG6i2h97GhAKgffk7239huBgH2iI
US6Bx8l3tnvEMaV7/PSY7XPdPgo21SSJ6Vn1kJNhPMQSlKSxtDA4AGuKY+QvKiPZ
SAwzK+I3esPIb9zcrA4XWhjDHXzF/hc2Pm46IPEjdeRsP2oZ/4XzRR0YOobjPS6d
5uhh0X8IL94OqcxPgM3Hg5+27F8rH/B3ymE/qj+M1wbHih4Xw4QlqM0N09MhEPu+
wcZgfcKor7t97nDwZqkytDzAYDSoMvRWbMsJ4/8Z89SbEe25qFnNXhAmj1fr2uoD
18N89RPXKI5wJlDRyZA7wOKccvHuFe6lobKTS8OxGF4A5hok8143sikXc0uL/qH9
U2SqRVorYis0DipzSY7F2cyHtGkoSpNxWtGcQ0S98/4wbDGRBncWlKVJ/3rXWOnp
fI3GoME0fd78J54L9M2vTgU86vap5lwiTLlgWe6tSRSFqAXOmkHsUL3QYso92PMS
n+5skRMu/qVIoitBCd+V0tQpepXUcN5SzXDdEd6kPDyThIFf024SEgmzoPTJ0XaN
pA5lDDW7LPSPBCSj2YBB65JG2q1VfVxnn6w5Ju+Vvp9f0ptIT242ds0+6MxN13J1
aWF0Ib5m/3NWKrYZWLUNpWdIU6aNJWZQtvw2DaMP3r5u5kbBmK+1KuyL6ubHTW3c
A2kagYSczuD8rPG7ZEiI57sqMAnSw9Sp0XRZ+tbQeE33QRKZay/469pcVhB9SAb6
sNIjShFFteatOrDmEMlrsJ0N35y6WVQIQHwWmG4rrqVpeRQ+LXkNpQZKnglOWuV8
6QcyP8teEz/HE1uhp5jJSMrWjviF2jNOogGJQ46JYPw44EgLH14Pv+NLVgpA0ftV
BY+wvyHRJCON12AAA8LsbxbH8z8a9C76NVdK1WJqpdnJq8USj06VuSTuIDcMpCYb
53uW172aKVU1uCLKOyut+9twQfDI2IwC/E68m85CalqHjfUSltYDF3wyumJpIXKD
WE+1KNfsm4Xu3PKBtO12DqBU9Xc+Zapqhk6I54wX+xfkzaJMunhb61BQg9vvWJ9C
9uXr5T3aQL9eAjjPpA7lfCClMNai9TiZOzNUSnQ52RFQZr0TAmFL++CDThLSEnT+
HOE90t9OdHSmnqCvjv19N1JvG/9DnUUR+G1/eBOkzUKcDs7yjuLhsdLmSlcXWCLL
IQ6edUmZ7Ko6TxSKBQ6DxpZ6taLkUXAX7KYZYal0W30mbaWCp7mbL9qCzk+sk6G4
Fbr1K6dAHgnNGfN08O5Q0ALEy7AKFfdjZXq1xdo7ddTbrDeRfs4yPOyhUQmAnKOd
dpOkAUHWDpY3sVgcXuPuB7dud5/u916cLBU3PSR49vJrqjKTgSiWLNRpyQhFzD/c
yXa/QvTR0UCD3qytYUCWCgYvOORpxZnA3v1EF5/OyZ38n4HOidH0+3gQND/lyI19
FpDa/DfbBELSZijQwaApGfwrGUNwyz69ZY2k8fIygYWX4yY8vl4Ap1lZxTSVeIgk
V6MjrE/nED+PhGr4gQdlNdhlvqtWjbI7SPT/25oHoq1LUtg+b2KIM4+gO9P7j3KV
kfzhmvWBL5ABWb6078oXgFW2ZZQlnB8c59SXQ5hL4BUdycZ4cZNtzZ/ZUq2eoC02
uMdb9LOAK/00Use/RRZDYpnmaNHteTaJZy92ZbxVjfIRS19/awCmHOHi0tV1opRP
KE48QsMvGskqwWteGm/TLRZ9g/MyDrEN7j9Z6MRNK9rqGaLay16EHeeabHlew0z0
1xipwy+BdnnmDa+x47K+bbCT3J/L5M/CI6kPcoFAcsWKzou+qCvDqSRIW4P4B/12
uyuqPocI4ijhEXu6bZ9s4UNjcMH/OdnXM1PmIQII4+wMghHfh0i/tlBMzA2lkzK9
OzxIgVdIiRP/FKloGCG6Ikoxj6t7BzpUo7ML7siICgrPJp1kslVtSXtvybN7XnPL
zFPIPQWGVuvzeEYgJMYPLaX4R1LsNy+WLsRivK5dJ2iwvQ2Zb1xme6i3PsolhKzq
g40Aq2rakymhpKXhA9WoNJAvq8oDFxzSWOBFwSC7nmFOdEWj98aZOTYq3yep5Hg/
PcEoiV2dJa3QO+WxPR+ksQeBkmSVYJVtylAf1FL5Po27Iu4lRU7erEshmAKaeICD
ZvZ0dsBgNd80VGl2J1dS3+OmM6vKOjU8tbTIe6FzwzwWvIFbjNURjt1tHz1Kc9st
vRza3ix+EBaqvX3uQ8LCtdiy/Eiv3wwYdhTV6PExjggz9p12rhZgaXUbekrkUA3U
Dj39SeDZXYG03XZo4joohzbAs9XEVySKktxG79Le23SCrw7DwSk+ChzKpSD5u8AR
LarrRiKstf8nVO1HXi3PVW9jf5uF+6eMOlDEwQyjSWuO/h2yO30MB1WwR0HXbR7h
oyoYiEaU5ZTe6atiI9UeeZNbc44J8NkCbBtXo1BTbi4We/1jm7GSOJbYgE5kFYBC
0MyYPwFGwD1Mgsmcgk01xrbW9N6xtgV0fEiYKjAj7vYeo/JKY7qcmuIY9eeYOfAM
bCtFaHURMyPZQbfROo7bL1jI4qgTEJ+JGYwOduKMKbqn8gHe0ChG2FmRusjNkI74
cZ5cnmMLQHJyvft9FBJ8cPdIpUvb717TZp7FPxNabbBKWER2rdEtL6ueSDVXNBV8
k114LQ/WxTesAWEDXIYLxL527coTBIqroaNwk6c+vknvitvxzYV0anZGfRue2qwA
lkv9j3TosItp4J5HMolojFfXeXDCzz+7RWnJ7EJDFdMEY+tDyw3YrMldM8JaPgMg
/2u6kkTt9yncqaEnGwJv7STSQQPAN0R5gBYe/sYBFB3sPHR9yu1WAV3aqTuPS7Yk
gadtE3jvbUUcd7z3ghZqV0Oml16uxqZxPc9HC/OQpWyI+EKUxvJiKn09PH/9Yfhq
OkFwa68wFd+LldFWJbax28rKRY2yyKMcm4/SVvEuTnSbeig5v8DuVhIuzeHJuDgP
kzr5lI7GG810qdXNrnj/9B3l/b+2JTRHLVmHAOebPuGrItIJVSCxMh6CSf0Z7Cjq
A2ZBUQkcV/wxB3wv4w6Oiy8D2f8z4x+5UKbp16FaTHIFmKBr/UIC58QxWAc5zXGi
KZneTipSOfSFnefmJVnPwSklWR+O3sinDxJO3EsWplni57l5bNTqv4hOclSrZLFa
i89QMA//Ddxt2VGmVPBymStOq8AcPdwVKf1efrVbSKyoGEx6q013o3Z+FPwxn0Qr
ueTOhm+WdmIewtvqs43eLThG3vZtziab90hqvbqWdg43li0guj7GkhT8u1B1A2hn
0hjuwhmCA9bjr7zeyrdYuOehEfAj7SgeZCocyaa14Dylx+ouuyzQj2+euNKKBC7O
ptTexoyn7FEICdR62eWOVejuY8eDVNcrnffjGkuRIelPxqU1cpKXq1Zq8i08uuFp
9Mxhazjerb45uFRCaN0fpmDpXQVcSa31xXHqhflsWU4CndysEDeENeY3wlIhOOG0
LuiXwTwol3i4O6QVt0oN6iMWvzPez6PMPQvvFyXZfBHWk/GJnzPze5LxyfW/p6sQ
lp4g3mHLl+/5VforbSLk//OlHKoyfmiarv+5bVtQqjjhDvkMVLbUIcfpc4GAMCDx
e5TVha0n3mRebLrrhOW8CtzoJCKg5qqV5vjYf0HhxqTriqszibx7YFWrsARCY+eP
CCN2zmVk9n++LQ8AuMcNwMObimMLByTF0oJ4D5r3IQoIRMTkdM/yNjevFOwHV46M
8JosS77BUOHtt4Itz0QPTNQzHp64FWM0Dsoxk5ThlRGG5DLrmUCbe2JHecCbrIPL
3gnO1WAD3OgN7GmLMnW8u7d5hvHgbD52d7PvwvCGfbjepft+D5GHmZqZlSo1r/p2
yD5W46+kGkjpHmiOPpt72sHMS+XXie9548zHgzsKOs2o7f+T/ex/Orwhl2QdoUN/
BfK0FfhpEHsaqXDjHaJUdH3kaYfkUQBrThXFX9IqEkDfyzkuNeAoKyVAiRig4Wnd
+zLTHa9CCvRuqAHvjSqxkn+q8FaQ0m+zoH3l91x38MjoCUpFs/zo9J1vwaR5um5v
Q4vD//E1vEN3dHqonDciFaIhmgDK0zOtCyuoFPTT1RDihZqJ4oAKZ7KEtTwomXfV
f2L65FE3+6TqnukMznyNSG7mCQ1HYP5kZVE6WLhpxw7YRvBhtI58hAaQkNcFEjof
OMT3l/+boGu5v4HP/iaQwHGp62D5HMs3LeGJMAOhqIhG7kP6IKt7orn/lIcHaAuv
4KTrmT6MQcNKAA2LDWuRVOnjC9o8cnmGiwTYeLottZ2yyZGkxq8tOlRe9iMR8V3R
onUdcoU2o/vn5/oOB4GUI1WZEkGWFsEVOwyUOFXNp+ol5UlyZlOG/CDQ9chHX2ud
P94mRU+1uQBue8S+u5ZJ1bD8ojuQR9Im5xEI5V3/0D0GNLP40UmeMEDtYPA8GIXI
Hwx9oIRciLGpaygQel4TvFzvrjclGoTC8QlLzN5ks6j9sxPQFErBrnd8RS65yaTF
FTgEuSTKpxA+QzoViCW57F/cX+cBPn6HFf6HaYNpEFO1Aznp/Sq5OjDaVR5yD6/L
B1FuJ6kOhWOoC7rdrgu8jVHsBRqRpH7+CbPv2fb1xnrnAPCE7nk+GqfTazb3FA7K
+TAg2QHWBeAay7nB92Zb8l7wZ7Fux1fhV0aFAI/EhepvHigvhUJJqvLrdftWis0o
aYrt2F+P5bGW/WslXeciC3fUpxA1sjUKXF4G7/Z4ywEl1DjUMQxquK8H6DQzZCA0
fwBLXVNfdkpoxSUY/PKJK8Lpv5ZX0v/IcaMEyrd4rC4knqsF9SupQobKzm5XZv0O
qN2/7rx6pk/CyrE9BWuMDhnCYKChyJwZ2WrMH2rG8MCPXCAWsXD47mbJAodwCDCS
Xlq7dc2pQ4Gfby0co/QLqMP93lPTvQ6OhPVqTq84j5ZA5NPU78WKUhPsJgaLI/7F
hoA00f/6qacA4L8z2255e4CIboL+mjA48xj4W8tgZTEcaau6xTjhNy6xOabAQRfE
3WVWRIV+cyBDiOU1WTgy/XD/xehUHmMO2MDlF+4+XJ9FQO6GCbOVc5mnuxLcbwR5
t17O9TnOHn1k/pOqxMhz3rzMgQLIyGZI6jA4uXiA98L2vsKYSH2s5J6dYcjhK9dn
ZFNB8Saj8V2X2RJQpq3/GBHJc53YEwSNbZ/bA2KHf12bo+FUItyyEzkJI7yRzGV2
AodofKbWFjng8sG9+arc7U7mHcf2TbWraStriPsR4ibXiBGiu1bZBFVAua0tYqCw
+qfwxbdST4nRVvA2s0A5VKhDjOhiSbRXZf/HYmJ1ifn+Sc/rWWt1DIgVkdToEQCY
eHsxXUkjNTVKnnQEraufD9f+4ZBmjT2DmCHwL8WluSvXXAES8chl/prpe7NaZOLI
f8o7vHRltDBesetJ7OP8Hv3cwLTrXb0S4OaU0ZHoEK/SP5TaxfvXsFbemm1WjaZH
lCzICzdE34PE9oAYHBZRbtTERQH9JqRBIW1NBk7YQvCulUt88Ef+fldMXbbikqvo
0OkPNfZ28fmKhC9RYvvL5eN1sQpDML0IwNPYLwa8yB0LTlDPDQ1BMcId3VgSta+z
3dE8Jd14Au5ledOcyyAC4Ht00X8bI8loc7O2JD9fD6Fgb3OT7GfI8H2RhKZ+NJlc
w9AaTygUDoAyRsguA5mg3sW5d0Ebnjr9/WobX2IWE01+ubAMo/qsl+Y+iM4XApLK
zHhqH+LGhoWM9NOTmlNBZ/ybJX1BdnelrIMo7e2IBEY+thG5qLc5B66PmQlwMv1h
2+T8SDL2tulS/ongoKFQVhWOioSxE/1tS8/c7ExFuKmjzpfEFHP/n61I4rwKh8jc
P9xf8NLxu0l8DcdDidSaeVuni3NQFleKFgHKiG26ZKi3Ha/Iakc58DQQamwI3SPc
3Uhid57GS9BlEU8p4u+POtZbQWLhoXGDXQu3IiXOx5qOU72P585mxG4CTq8+B0xM
YzM2qd6EBfO3oS34y1obauAMgUm/xkBCir4JsVxQZeXivHAA6TFC/6NW5qAA2VLs
b1dmV84i2AobemVxrjf3QJ6mGu8mwxFWOJm9agBxW+zf7qk40vK5nqN3zDy/vQM9
dTXKRjzQr//9aXY445tI1CBX7zP6N8KbDWdbAX6TwGMIpCvGNNtJbPooYwQJSgNB
3tk9iu5Xtnjnv/TT2NO7L6dtvyPY3BXMbOBII/eOF6mT5S8vd/JfdqM/UfwQqor0
zfNZ9phpwnn9kYc0ToTgC4AoMzuHv9eJlDMYgRMT6DLWXE1paQgQdwvuD/fm/lMT
bLHeSvudcIs481c198A+NrJch4Mb2a6zi2+b+99m6Kxfl2GyTbdahvCSWwTBoZjC
bWzluhNwtmwsnVmUgsOUgFiJlziqvPiN+U+oZ6hNgXbn4Irpc2+5V2zaK++A8/RG
IeqwRZZ7EKlZIz9wQeJ1hfbHF6yUzbe8PcyDOzWIFNl1gyusR/I/g/k26ilvlopG
8jBaMJeiHh4+O690hbVqixOkC5GV8Vz1gcDPg5VEOsJItaOZsCyJGuymY8s1rmt1
F+1RWR5Li5OH5CXjI5Hrh/IYT4onQAzUh56ZfuJ5kqZV4L4FWvVouMjB6xo0BEE8
R6snjUhbPEj+JPCWOQ1t4OHjAtnditd2dPw2uXBx5UKZOFwTAio1hubnCb8uCRhI
3T7ge85Y5GzuInl+fqW0rN0QsktsM2xP9tmPq4u1bn6Xkp2Ka38J8u3Nt/M+NYZU
cwZht7YH2JongCOmfCrAqxLSLWENusVRau9uEbM/HWgrYmWrQFjSU1SwB3pYoxRO
MOHwZyVbKU+SfIPDThQSbwbci0AWNQxN4pf737qjCC0dEKpsYyjDVuKjAvBSG1u4
fKirYyM8H9zLnB4cSGOwEO6bJT0YLHXeJ+wvkBCHxSz5coSAmK+LeO8rMkK9EzrG
Y1a/BA4wB+1UZ/STJv5Yfczt+kN3ux0xr6K96oz9YnRTJMos91fyYaRvwaf030gU
LtdtmH9x0v6Y9h4hu4B0bas7GptEUBmFuJ6ByyAOpMsiiahpZvpO0rRZ+sHnz9Ud
XihRhVuxSubLwo3FC48kzQ4p9ZogIDxWMa5BERz66+N9pfyhvG4VRuscX17IkShC
4918dClvGBJj/3h5KmW+KTFnshZvb7TjFOHgmmd4cENKYTzI9YfJ+6PfXWP4Jyqf
pdkuT/C+hAhsDszuykqP2dBXAjp18dm3/X9txNeALcJUICGPycd0Cu8rJQpXY5IE
Bz30Ax7S75NGuQHjclNi2WTdbbGnbMeP1SoNqPAvufnSi5XNT2IuESdIouzjIWCJ
46EAaznufNC4a/YomiqMwax1wIn/kynp6N4nUS0DuHfqb/XJUoZaXitFftHX3iT5
jYLKT2M7rK8spjRoGHnCfGTAoAq4KqdX4rU2lZSGsJ6YgUt9OiMWwaix4t37TuNY
4wB5+ZQMfCwLiSm88klMrFpuGJ3DHQV9xwxWiX7LVijkmnDRlD7kLlSoylijiQaL
S7eOzkM7c2z2VU1xL7wtTwQB9kSj7I0fuwwRBrc8O9jmEn7F5vFdYOBpKWVIi78v
1GLRaBZoiJZlN3ude29Ed5MMfWrLscdOqXx4d012TqLey7LTcpY/yaiFfUuocjGn
PYTdKXG2hQNoR9OUJ+BhM0gsgd887dLEFCefuIaMm7Z5vuDAX3mFOgjlRK5U5CCZ
lWqcZah9DMupybeAG8OgoYUdijEqP5oadOsIyk9jit0qjxiSjz9Y+/Jkk5x+u/T4
vkZKlvTdPzr0lERfPQojwegF2r7AyE2lFcuBtTx8dKGoTB8rgEwtGN6QCAy3oDxM
Vs+unjhmudjjNZ3awhobkqd60ZwAiowkVFQbCveyEbs64Xdov5o+J1Xfy8WBQZiC
huxtgl+tIqL7++RbuGnJgdG2vv3RKeaATmhWLgRlJvefDAYJbCfXOaEVaxtNwQ+Y
/sDST+q8osnJhTldpnvLbYQZsFolB8w6g6yNO94QDPg3rPl7fk5tbFq8ekS81cY9
/DVWDX4+d90Sat+BU48JcjQ1G5GjejsI0HFp49Vd8LNgvEH9aRTsUA7rShvFICm9
6msWyEtgYGmEvzBIuPQwBIJf9PdpK0BRbBa6zPdKUyrjRMSNGFUgXClp+Y/Sb4Ax
ldXCW3XqEyQTMzQhPv3Eg3UXhef9VZ/Lp8LKVQhnopbBsSkC2ijePUwzU/XGhDFW
SEtIcET8jAfkeLLqnQpn47RnZNSHYlR/5iUjYXCOGhf4lXsWuxo539ESc8QKngk4
NNb8JVQrTPh5PmHZO32yjjV8Aj8BzrXGum/mOBAiehRBkuCeAnWmyjAp0aFotEJ9
NkYBhzJgqDtg3L0HYEzc4GUiKT0s2Jz58A6k98tnDG/cdwmexMbt5qiXMMTg4DB+
Mxy1jQ9Yy7Gmqt2BsC8yz5cHiAzg0WQ81nUWGlSz4uaI385bs9i1A3RiKk+TCeLy
Y19H0cMiRoyvmWaxisZei1hnrY50LNIEaxPXylhEkQ9ec1+f571jE7QaJVFHMQpX
QATcYWfr5SnWkFW+ROJxF1YAuqFjrkH4PY8awFCx6t2knhbnAqcbnDQv+1QpRJas
S5B69OaDmbIDnI9vm7pjMaG/epX3qS8oEsKkHmZBKydARz94cBj6JXyMXwHJCM18
1HFTGP4v8cjDaI5eiHxP1o0av/AHbdQYMdlEaPXISt0RZXPpu8wk+vG714aPAUN9
1BS4kvFMW5ehSUy5GqIFMVweGBx3c0fIsT3EpKkJ/1l1d+JelzllF+ZAzoB3YmZF
KpbfifZ2cylwCDoNQ4GbHv4fZWsbMuYzVbeegKlxT6U6ksRa8vp+i+M7S57JqV9C
40OZIVRRQ8H2RCU09Vu3K115It2DgJ+2Rv/qTBzNHL8RG0ekuHvRQL863XqWg/ZQ
/KEziG6AErbzge8mQAupTccb5M0kQTCB0WCg9pWmm8t6wKQE8+fMLMduHxDDVjpN
5xjI2uO+N8zSMrnBMYdF+Dsq9HLYWt1BbOvZ1UXIhQeE0GiLENkKUxKH8R9SGgnU
idhykDpavKiOYrWdgFwGUJ4DfvXEqHPXwjE5xzw0KmzNjKwlY8GEr4Oi+dyWrKaU
y+uZbD1yidFxLFLxaQLuTIfbN+T1RV/sDdiInzid1Ai9+6YZy3sRV42TJ2/1wAth
WBJRax6RGgDs8cPfkH0Ui0iN0kDQiOFpxTZAJnk1VsGGVeoAUaSAtkudAt+zccQ3
tfEsf2Q88/wazHx0aq5tr2bdH/TNWN98OFKrFbwz3ypQ00BLW4BO7UK3HaT/taSo
+xQQoGH20hvfnAJTE8INaiUscGMk1iJFtmh0hnqo2b+ET8CBAb0Zs5tO0yJsMcqW
2eyx900aMMGf51se6yK2rYIbn+gIzXnE0LDeienpvn7vb6Wx5pwQoMwEHG59b1+q
0czu/D4qCKOTeRkzzBN9kfD+70ownF1kKVO1ggvnsglKql2qpPUqS2RqNXFjTti4
2xO6phM5VXlPoILLY2LMnbjIFHxarHc1lIl1bu+2e04CXVwcQxHg2rqrIl/3jN5U
Njebjq7hWVnsKP2hOivaTUoFQXuZ07+iWI5PA3I2KxPBC4FFPG9SwMI37V4Eb6FK
0YbrvCjui3oe8a91OToeSlCu1KYZcNVOlQDIzd3bonm1DghXZiHmHah083udnjLn
Tp4MBiCvGT0KOwqFfj5BhFWLd+vLunazJZHC4YzdV87WqJ+BkcCWLHGexauCup4C
o7cHAtpWe8Wtu3bzfBIdi21in9DQatHJ3o2U3l+c9GELnEmjilxLPhjZhtepu/gO
05WOIt807iajkwVWaY8xInggbXPsnudtOSD0fPO2lgMAQqVOJlINGsdIqL7DrY/C
wlV4/nwEXd0KwK/9F2fFskbM+k5sfImwIyaMNpFG4Hm9dz9mkVTnDBjuCptRbp6v
IFD/uTUkQrCcuvRUQgzQpgcQmAc4Iq5AyarnKLQCJxK4JXEfl1L9BvZeARIjmRob
QZCI2vT64T2o2haj8KeSxcVvB8Yf1HEwFavlYBmz/lITLDyFaWrXVZrUDkVc5gAm
QvcHtaeVFDOPfcyGrR7mA0sKga+8vUfK3fxFbQ+VgHRnjDrSYQ4qap3AqK8cnAeS
hSORBB14xd53kXDq06JiwVPTz1t9uJVv+KHn0YpiIJGeoKldcI/plgPapUnTPbIg
ieIQlIkekAgBVXAZ0YHAKKUNfzeEUTj12m7athEnBxeJU7TQ52sZyQBeDbJGNUW0
DtFy6tTGFm+g3lo2J7FTXL4n32fjjYZUvzbUVY8ev3WzXS/dCuOSjihAqQulYZXo
yJg59JSRTAzoW7lecg60sTZ41isijsVmfPxcFaTIePA47SSpmJ0/lBbxea8Ddjdk
q6a2OqFUqiNxFry8VYOVlwjrdySt6nEYgOnyDky1nwuV2ZmnKdmpb09K9B42VFd9
MoZmdxw+CdKkGT9IJIXjTpf2NA23fiHcAuEUVU4/I1dtjTi1RNZewYlt1W2lyKfj
VRs0dfDjsxQ2eEwMSmaMKuCVHEqTbPRwA7KocYlJl5MpBA/4NWWdXh9aLP8VJwN5
HmnI5V9j3cgP/AOc+u4xCvdsgjF51cJbU3129IviQUz9N6DZan4upt8bdvsccBEY
13PM7tBKtM40hW4uKSE1ZlvXVhe9K4WkBHhWKqUnjrYpdm6jwIhyDqSaVNpiddie
aPcufwWx0MP6QJYdawRA0KDBv76OwUR0tEoe1/RbXYcKv/t21vEqekhyijhU8iAW
Q5wx/5YhzUezNYLXjC5UY/thJkMkQfzZCCwlKnHVJV4DcpKi09flIAimem6k9vq0
hQ7bdUxudcMq68KL+dJDdq18jIb2rTRHmUXTLJQ+gHazL7hUavI4lBCHRwNOmpqy
g35Fl7MIVVuUovcQlHCNM3/NoPNpQz8+kfeWLuxqTGt1gDyeSpLWcLcUxMPu1Uqr
MwKo3rw+Ya/htJAeazK7qSSybOaBycQ7HuwVHtc9rzNH6pUPNlpco01sn5hW661W
70TtV3tCi0QYg6kinB7REoyeE4ZdDHsEpVXSp4dAu5UWVtXPjsmSTF/VNVex2ISc
1TlOLI+2JRanmInJ4p+F8BuK73rrosx1oHsR7qDNTfEoMC4/xS65wQqAs37D6b3O
PGaziCG8NgCPm5Zkta/APYcz3E8X6b/oVZRqssQlV/Ds/jufAb9/s7osvRbTwnus
9Fa9KlqP1rUlay5JwWBj8/1kR2dFk2Hf2aKsY4v+VHx7zxdxxgPN1BfXMMB0dgfv
xTCpTbxqgcWuVHpDEQ563RrjoNcLBrjAXCRwUBb3xUTZo2cVCjwpDCFVqYSdI0MR
ekTYY7eIyCcjZ3jX3quWjP4NwhUbgAwR9hNw9N5vDcZJdtuiyH2UqBxn80siO7r4
PKe12uhGaM6oVQ8JLm2SvbEVAWbUech165c7YNivaQO0KfqOoJtKMeMWPQXZY/cY
H5wir7MZyVeB/bgyW+BKO5HDqFjAYxZJCASDT1QhwPGEagwCJAOGSieF9fT+GxnX
XyvZuak+8kmkPfOYn7LL0zhcWhhxdLHu7rMHoeoDp2csccowCNfTHhks77GFifub
RS/2kJvEph2Qxlxneyj7qdE9e96gmsPX6DMcfMEPrUaqW8Yv5859y8a+IdmEd9S2
pdV1vvXxJT95zHF9Z6xO30J/kdWsoJNrYYaLVRQppKmPb66PWZL7SexpK+K6Pz9U
dFdCnRMcQY14h0sZmDmsIdRgpAAo+2TGqf+p0jAoHlA1VJTvyIqgybh7nvt+TVLi
vc66FA25f83zDOa9yQoNNRar6aaN91++evAyz8JfGCnEktAa2dSjs1Iu+fK/fTO/
MoOsp6vHf1jbox5UiOLJUsPrPkBsSINcWmxYtS1GuZfUyIvdTLy7nZIR5xi9HScE
BH4qX0bLZWfveqDjrDq74gH+6Oz8OPoeh7kx8xri5jiNzPaOY7TsBIyitpZS2siE
uDZYQnnv7UdpNXa4mi/jV7yxSwBMqZp9IJu3qnKse/BbXQsUDxLuqI8tIorudLKw
hQ6zS/aBC7FzBylp0n6IGxnZ/rDAUd+QZO1+gK5/BLQjbwNvMmQlj9iGfLn5cCeP
ohYsiO7O8CudLYFrFJSn8Zkq5+osCK1pg0UgdSAJLE7HFZIskWIXfxc1su02R/vo
Pm2ahaG/h9yWk8RYB6Z6QClwbqB979LQRcKzJIRiVjFr19+z2/0/lTltUWR10+LJ
6Ier3eBKee2FyfMHUztgLhPbruLS48+KOINyPd1+NQSJiT/xw5uTqKkXt9xx+WTX
5NdyD4JyYgbTGEv+asyepLUJIWH333VQv5vDi9/FXY66DLrINKD1c2g9o3wnZaMW
pyQD88dNTMKKONypLRs3qzqvZFvYZ6TAqfP6c60H9R9DK8RYcAOa7p5IJaKMSJPT
jodGhf05dRPhZYkDpgvsitNEP9rUKboFQcjpeDGy8bPUNl6HaVhURqpBQXN8ru0f
emw/pY/SNgE52Phe0UVlyjRkqBdbtvPiAF7pwaSOUdpASZ/wMC/Hh2q5wESM0cQN
u9DZqpC9r9+AS6McAnxtUvYNgTeqoAQbvkutAZMxOWr+J7SY4KPaCFe4dng5OtxC
uLZeTnsNtLnRcWRSx2FVYGAO9F908QT4AsvCwMcCzg4ZkLz37nq6WtDrGXOz536s
+vl1YmE4mdni6b+YdBTasxFGRTduvwJBwhnUx9RkUcWlqBrrXL8GnuP1Qnb/1cnf
gHmSDEBoxtzx3PM+cEssr8NPkFuWOTc2nRO7YY8P5qNtIS2o/T/vRyc8nrpvfjZ/
C9kGDlHCpnsRH+mLnh7b9GRDVve3iDzx/lMM5pdf0nw/Yxiyvct9mTIKXPdGLfEm
8VBjtuTjtigPhU083bWAmRnxLsT4l12/jr0ehfEW6iF1fYa+tn6wCLlWGgFAndeJ
2yyDKSMIQSF5eTp+rE/crTbSmvErkWpCZu0BXynKs6WD7oDDGpBstg4M7CTZFEzk
kcYPuDJc+4Y3crsWegCnhYaMJVJ0kcVVBgtItyJH+WhQRZVd1BftWQZWBk78sRLv
CvM3Ess5LQPkHPMlnncbndbejoiqbSOFkO7xGzlEP6Fd+cPma4lJ2lhIcDlMfjHE
taLVyBrmDNScxOxmxd+PKygrHOainqHBYlhf4taqaKs/3jKAmKkl8dkrVjn41qM6
FwR43TFBneV24M4NyglXF80EkgbfI0awrPbwu1SNyyZVTyn/I5aDbxKzCMVqXGcU
ZIuqs4u+J0lHN3kTVM8MNgwh1PViAZ5H1Pu5Oq2xl3MgejEPpvXMA3hiMqapD0NU
XnP5LnDhH+hrXq+0kqphiNKySFK522faXkNvg7+p/FUQ9Op2fTSuoAnW+GpGJSAY
XAYmPQlRi3h4foktc4hTIsuexW3cHnIlVs3ZK9kK8NtmVLgDCc1VLfPga27ePrZQ
Mll7CVRqtIuxKhl7P1AlNFylRvtC7eGFXkgdV16FlU7IFwrqF3PloPMCkBJACswX
g3HvdxpIMmN2WpOUT9xdMRp0iQpDmKiFidRyT0CECsAGD9dzC+PciWQm2ZV8m6YE
zHaFZOEcQ46euSpF7lTYjbcLohvsx6Tn9Zfw2erpySKb3p8D0Xs+SIPsepsM2q5k
DDPR90M+0kUFwqaydaMgERHmBEv6Y76undawrm2XyjjSxmX8lFnd5lptlLCX6r2J
xBitd3pXc4AwA1gZBPcdd3YUBwjQ/KRxgnMOXiwW5rreYsbosjyzd3oEskEKYvsA
EEOVPMCnroljP3FZDDZDWqPGc78DbAgYtInuMzUe7rvmVkSqLRFKNHnRhg9I1MwU
HX46RWvMAfnX96mdzjKFpaKd3p4+JytDgFgiPsGVEepB9wf0FyOhvdkiB2aZ7eRx
iwLYFPvmfmcoJmK8ScLqRTd7X4R8P8UbOOmoDRKGj00vlMSYZjIhCvM4XRrwECBc
XzdMISJAvWFsftX/2AKGIm/qY+MHk6lL9OphcpmLY0iRQvDBOwvT/bcPukItwm4y
3WwLo6D9cb1RZQsW1FT4AxfZUM1LiHAqDpGSLnM9EczD1bX8A8Zem90ElYsvcSAQ
VodfBGrHupFn/aLLu5QWPqROgwGs4sD3R/+3Aw1G02doc/FOIkWmRx5r/8X9PXqH
Lyddwn+iJAC6Lyb+GmltxJFh8MqsxrvhPkgVUTIemS+urqol84SUqOLLtoNMEV++
XzKVtr4JhmM5x5ACS5GumA5oGsesvXilw/1PX8eYN0bR9v61HjfvS//akTptjf3A
mS7VGZEGbujKBtgEAAUH8n9nyCqrnTwbig6hoc0AwBvekLgFyxO4WBcDo90W5G9K
VYB5Oh5XUDFdfACwFsNpv/TySAaVx4Co0whV2RchmmXVx8gFTdsrPfIBrPW79sJd
KMKF3KW5DgKiQ9rB2mqzZ3MsmdHPO2LAXIZ6FJmA0BOQ+3BtmSyJgzT7wp3uoMmL
kD4nPLHrgOB0Wx5QevhYdrrWD3d3KAcc1zZozQ2XQ0CNCEVc+mVX7NId+Rzwfc/L
/DrZHttKKIa53lyb0j+euW1bJzt4FGkLqafsVeO2Ky9GJC4rKNUNePVaCqsiEnS8
ul8oj/82/cxAL0e7Mps0/EYjaiAqEOlvzrZd3YVXHb4+ePZNHASlY+6psCxaLn3o
dP+G1y1vYJ/Lz7kEkNQ2Lrx5TI7b4/C22hLOxSv6s6Ab/chrUtrUqyZ+zEyOLKYR
H3McE9v3z/cZOsAlHs/nlBAhbQfvT1U7Bu6dwCYnr+8zg/vg+kwXkuC9nF2JW/hD
gVvvsXGickdGKoydKYKW/PsoyDo37WORSkXYeDp/2NnnMUon4bW15pgIzj1e3eHt
MW5WLQoMX1Ajr1vUYdMHHBpOYAQZYYukPe2cJk5v+jz0yGfwhXFa7MFM6rZCRv0E
A+d1daKoauoX8drw+Jw5yfRYpPfI02y+Uy28VChTD5VON+AU55Lo63Y/ic5zYHXA
56A/zgmBaL9z1cGO3Cs5wuMXOgHOmr7uutaE1vHPHerLEJ1HZa26zZnWUUa/wzs4
IvM719muahp2KnFd/8hejGss0k2xBya4VzCaorS+36vQOdvEhv//6QdZDZWgJa5B
XN1FI50PsTkjzYjDXIfKzIDXtNKRKNCSgBzFqszg1DujYiFteVSr67BET7KGIvxN
pGu48gEnLutM+y7/SpRYRWxstfr/EqDFfQ6OMFFT8p2UU1X6pApb2jtld40NIlnI
ezcPTgm7vH+ajexxM8SqDLmCNrngFqO1rPtOUHs8pF4XgqX5tb2iiVIFDbt2OeKp
3aZhPcxO8E4iSGtAHoSpVnLcgGAmaOexuu+oLz+8uf6rfV0Nsx4D0u71YYPhYKZd
zqE0d9XBKlJr9gEdkh5O89AlhmovDlGbfic20PDXrgvxYPJgfglNbBc2rTuPaE0j
xU2dEGLYFT6G9EJA6quSrC624S0y2wJrJ32M+2c1D8QpSPswn/RtcHVsKKJxa2Kn
h37btKsfWPeoqYZoFLhJk8gA/2WFcmV9+oK59iKW30D893Eq0m04SH8r/C+X7Qrm
XfjD6ArGAtoy1dIuocdIqh/sM9HKSQUtGs28BshitSij3aLzSwq7fc6Uwk/5e7PU
vtpsMU3rJwGOBu2UNBqgqnGc2HY34eYCQK3GiJ4WpwP+OdGjvq52F7mxY9T1RTIJ
pD4+xGHotirY4S4UHip5Qh4U6cVpZ4s2mqJs1olqKuRQxBmiDmKsc2+v2FfuBCiq
DGoxS4F/JnZg/cPdz+0mraFn9gCpFf2O9JGrtnr1PtaijWyoCvHKCqjEg44s6nqA
0ETGtd+HYy+1/hlTlhmaB/Rqp9tN5IsNaOGY6vcACjcs4DiP01LRt8Rfj6kYr6Z0
gvpph65YjycY6CyLrvj7gHbQy5SIG5ekb2u7HMkd7E5pE3E1XXoYBfhXnpTKO3u0
Tk6vJD7gbgH1MlOe5ykKnK9Q+1gzM2RnmOx+2sC65w9fwMFHCqvbuflZ0AP7YFbo
ke5Jb+PDExaS9gSVZGc2PWjZBmcJsoTFMlU44NI7dt2v2ruV9wyxL1vea7a55cP/
BaOhkQmnGtmLz24TVbhrQpzR8qfS6FQSQ6o77dqefxTjxayi8TLakbSEGnloh61W
iC2DNcHZjmDjN9kOewK+aDrBCMcl1ZzvrCwF19W1RFzU41jdMNs6iYiyguF3hIxD
/dGh4Rt0cOW6fnZ1+ZkvslfXpiNjSf3bV5Zfk+uHxTSk4tK17h5kHBuu2qHWA9w/
JlTyVoZxY1lf7nUwa2PA4tFgGK7WmXErDv0nfmWkKoHM6scDCVFuqn3SDOOtqhvR
avjT5xGfzahbw6renbN0Camn7mE45ybzsHI+FgCU2TqDB3Yt+0JNKGRTfj38dlRZ
UKvCr7HelO2gwHc+PR52po6dCIqBj6xhbl3Udlk4qEzORVp1OlVbcYkxadJ8WVHh
D5Ncv6UBPMSNfYRMeYL0UdWBsgkqFU7RJCYXHQ6XGtK+HNlgfKudx20vqi4BJXNL
wAzwwO7/yxDwKlQb869x+9LB2mbHjsyBYhvYl4VCequ+yJ2buOySO6WBqI0l67+V
gFtNsuAuGlD0yw+O6W2G9Vcd2lYvKK8mBdz/XcE1lwKKG+HH83cEy/qZKBMBcPbw
LipAwu6nnYBJoZhbD+CP8sk7A9nEQlQlyulTVc+l5Fp2jj29S/PAK+iAUhMEU+nI
pyn5lOhxJssr+IgdeZ5DqKty6IdT6EsBIQdOgpaGb64zEb05StiFK3Eeg51IWobx
5qIrizBDO3K7jiegupEwx11tUTFWSN8u4UcwK+p4MaJ/8B8T5jUc8V+tUO71Jfyw
eHf6PdiyullB9R/Yq8chs5Hw97O1BIlDhPAR4g0+vnzjqPmAlV/fJUUbTUOYB2Zf
gfMhyxVw2PdoI1ed4Rxacq11ejhWB97vVd8olIQ+tKWWyh8f/ZLFLGouGSq5YfjF
Zv06H5zpPX3P0RP0WVOzL9ppsYipwxent1yhyIQVFPc2m5KtNQ/soFdzrtgDnaFi
b+fph0lMOfm4uM4QQgnuKUhBfOWDPfmyJoEfMqZY8tt/+8UyANhyQsUsxolh6Rtb
22PWd8OGjhU/K2vB/DqgOQY3sy2AiFTua4h9IQhMLvMFQFzkC64TsRj4TbFw78yc
kRyGXm+YsKzhIe2s49aGYAdztFZ695FzPBW6Q/euppkXHDeHAoK8Vuyjt3VRp1AU
f7r2FftV0tqsanwn+LVdFFrcLqCLRFAJOU0JE0tE8KjNR88xhhNJwwf6+XFifQ5F
nfPQlNl+jGhcsVifUpFjC1TFd/ZiFl803/EoYpyG+avmQMqELbrW/4JBI8V/56iS
Ng8yV+oIB+pZsBSCdSntd6dg5USgWixFQ6QLa/WN4D2beND7ImPKQkAA3xy9IULR
tJ+ss40tGne+zAoYRVWAtMboudjf09UrAnT0bTfmUZhKkBU/a0TEBlFOwaUUke+H
XNuCfAc9xtWtPYjcS6vslRy/BHLvq7Mxo6O3m/JdTj7KHLjH9xHCYrmC09K1BHnP
uRton3zqok5RDGK7O1LvtXnEm9Nc8TnclVmBm24FKT/RRmN+n8TqESuViGQkCxZ1
n9G+Nt3dgQconib67k8icewz+BhgBWLVnfL2wD7IwOitc8QYI+AJrm49H+XieqXr
doLDeXU20CXJUDgQX4L70QPqoyQGNHIhK/qXS7o+KmqcS6/JyzA3xs/dtxqqFe0D
Ubyd1PY2Sw5IJAZb3Ud2GZkWFTNaGxbJI9wk7qxXiR4X/rEoGMrIXJ8/tMYoAsbr
ip/hJr2M11kj5+bg4oDs0kfFq44xQMMDk6u53Tbe13Qi5c0uBE0v5iL/xnkVTvLO
jwProwxskUHi3zLr6uU3axrZ/buDN0tSrpi/UY0yJ9n6oryionzYF00xRArUzFQr
oLqfstFmrOR1LMiw/fodEhMa6MQYa3l8FGJ9gvgkReraBhEDqallH2b6Q2SkLS02
C3wH3bzHK4pbuzM+6FzOF61AYjLK9CuzZWq6ktRR+v/AKE0GCq+dzIfiStUkC3CU
8NY0ky39/0SaEkeBPvpuRwmrdFOenqLzVE30X++u+Zk5G50BI0unYYtZHgn8Ry2B
5CT21bg1jtgWR+deyWSGbOKxAhKPgMONh1fIZR25jgUKeNWjTx38QAjAmC/ipsnl
1AsCgQD5jF4Ytk+cG0HQf3YguWXzZ6uRcQMk2rdMUPH/fJE4jomxpEtf+mzXjALh
yQzVbToAn01yeRYzzTJOB6FdC1DYeqKxE53vQzP+OTBjbqyZbA9thZh6bQ5qdm7c
YHJRCicYGJBcey7MeIclVwejDIgFTcrEYlHZe4di/24dAjP6Jw52a2pslgKYQfll
9bQk3m6g6hMz9e4Lw+av/HUFvzj7WYoFH3Jsqk0Y8iaHshtIXaF8pc5XPhjQTygW
mjcdHLs/gPOm5OFVkjl2gP41q6+2GiW7DS2MHHb+0IMuMWr16ubO4wSmNkCOiBuA
EZ8xkrfiI6mqus+vWpa9xrHMIXVO5PhqMyaUlV0XMm+2qZGR6EYdt07jn2ysa3T6
zAVv8ufhl/aXb4+6OQwR6kbM7UCVQXaBlhky8i7/0FaLsGkm2a9r9Z9dgFfzXU5l
9C1Kh9ovpSOEZPY2hvMYdWTHg1Myp4/rw6qbU9AoI765iLr2zF2Pm8LLruePi5VT
5qRl9uP/9hGWIHFE4FCiTzAcDJ6S3eCLWSYRBL9+ksfID5k6/fxa/3+OMmDxw77A
JZK43yttnNBT1rJ0brgvuz46RUOfZhA93aVkSv3Mq0s7PN/CG18W0gyz8xVT7vl3
Ytq3eqIxqXzUfvVdS6WcG9WeH7Hi+colee5lzOXRmdsQBk88rtEPclj+jnEoDszD
uHN6QfI3VJyTk5CwIufMcPmu4Kwp3vLMXhtgRcY+mRPV/qwIsv1s+oajkdsBCBjH
ebaNZnU6cjz9PWLa5qcRe8zZ9cxTO6bOL15clM3UNzNM8r7gi2Hw+Z6LojxqM2su
Yc3dijhr+oB1VrS1qIejqLWJfsmE1Ul82sIZ3g2L96A3bjwVapZQ6q1NEKDNk+cU
EeH/Tt/DaawGiJDpR/7IVEQWAOvxiTIQElhokhuz7JNeDx8EDVNFLNuotsyhz9cc
iLxe3317lqpMwDc9jIytdnuZ71NurUNiik1RBpW972poTFJfYmWPLB85CCenwA4a
rkUkQPu4MU/c2Lbg+74rz7tYiuWViFtPWYUWlHLnfNpe841ObBTOHhGr/Sxw2ymf
0J4u9DCx+0uedQFLQvT6oYTrWT82RzaF4Wlogkxh2DKaIwihvjIJSnrNvYwKm6zM
nphOcjcLDV7apFLW2KBC6HHDVnNPBn9FtMa2Yl4VmPcNg28c8Ac80ohEhF4jsSv3
woPCgTtk/jTzcHcukVNgcivhbafnNRNkDq+hl1PZntDPts74+2sl8n7LZWkIIjFs
4fzUUpA1fe2uz8My2Kr1e9488UpizvPOMHCDaihSIF6v/vJ/2Bsmgdm7/Yrknq9T
DzOokvTCBwr1vYscHHrMDfcEk50vh30tdEZ+pNGyJcJRQCyI5/jubmr3ICWeGF8J
cGo3Wr6q0+1lZz56UNzMV3aOLzTak/2hYyil5G0Q/PUddZTFeLVdXPcwHpSUMmMg
pvjLghNeN6rVpRATAUYyIylixqBNxmn8GdsUKNTRJyr2u6iN9+HuoxlXEQIq5aDu
ldCvxb0g2PcKDBFtvypN2Npxr49aB9kb1goT5gfi6HGhQAAocc+nGAEMIooQTnpq
02YM7NC5weM/1a2kIn909vh4jgriGQpCUpzrdyWdxSK2ud1ShOhCW0QGdGzcJcxv
44b1TRt1Xt6cJCQMuRrrZ5aIN1rs/z1KQct5deZjakKOOTvj74yPThpmm1z0o0UZ
Cl4lrP+GdMh6pUH89aelIajjEr0IiA4Xwp2TQOB5JLQSfCaoT2YK8BfkuXAflG+R
FNQrmHaXPT6xMfx+goAn2RGdnAAEci0tvwiogOBRrv9zPyjQhyTYTuEVuOu7bkQ5
qAd0rVp6BCmvLM4muvw44jTP6Wf0fFYNqpgmqGeFuhbGJIKRCJTPBgUhgRtHYSY1
YlruUIFHem+ujU3MQ09AG1+UsCWVAIdwzgirYxGuXk/iNCL7UlWTdrPyyf7ZFryU
lMMOtkZK1JVaPo/FcUmH4OulnjprH8lJPsVjlvOhRf2yznBBWNW/3ING9/LmHXGf
t/Abx4o3e/rw1m0ZW1wCpHedkHPVbCIhsv8l0/UuELj2wyjywRhuTvmP+DC0MCcK
fVlGk0Q1ejb/uaAQV3qNc0SB/CDWHOsz92H4QSue/90+EQdgYIUw6ixcIfv3BAOr
1DbvKo7FX3PKpAu3XhwDUXUgX41zntEhjqRJqjYCPoIhjrYIL9m121+h7WjQCYJ+
OdPJz1dm8nBsF7Wpu80L6VmK/DLkeKj/KFn9p7VwACuGZ+cMrVd2rJJlmlPEtH+P
cXHWfKdkLir4+9wJGg0gjxfaOO/ErMAJ2srbxQvAOaZF6jDWbyynR4Eo65LkxHe/
hH47mQcgwF2c071DNcYeXMyZ6jYrGdt6Prz5iDmGTPJJOK1OOfTf8CCbaihjEAcy
Q3NY5EIOam+imlTdosaqTUp97WY9/Xv7O4vh519ASVaFhax1/5CulvuciOoRiRa0
TNf49iP2Fg9eS8QRV4Ul6kGI1IavkA3dQGeE7oSQOEILMTmQT4Y7Y6oQ3SreyqhJ
OBG7xhM1vorsxoQJ+fhc4seKYPJm99vapOWDgAWo55IDtwRrJJ9Cq83P7pV+e5as
kpeDa26ps1xhdsXbIkklAUW04tgjKPCgx0c4McTc9KZd6Y7tgxVuH9mIi4IaM5rd
NECU31FpizWIxWRYURk6hjQP3fEjLb7FBRlvvu/Ito1/RyA5MkmduYUz6XUmOK8H
Df4JELeAQ1fh7j8rHXUXrYMpjc52PjANm3b54XxPpf+dN9jidV2zPMVPKN49EWoN
o/89X4dd/uF0wA5WaQRnJv/lCKLAZxYVvH2yIiSTOeo6TBAmnbHY58rpih2rpc2V
iHjvz4QKVCtkgwatVrYMoEyuL1nin0nTA9BdelM4c/V1uOtJPSMCwGdPTN6G91Ke
eKt4tn+jqTqnzE5qE1J25haLlgqtOmNnujTLDG1MW/y54BqZ88Irbp0nZTgGOdtX
Fwt4Q7qYCxQbu5nppsozA2qlLS6bPhLWo6EqUoIppVTzCjUkk43WS95l4KK4P2Is
X9Ee/4f3b3UnVltEmU/ehHsRMfleehtvAV+/ObEvqaZ/ZQBdYinw/EtG5YnEvH41
Mh1jvyLEi7cvQBL5JZ9gpAk0QvsJTX/OxHtQzBLOKgaSJohsBiICE5KyGlueQ3mk
Gi15UHrDIsHRACJg2sXIdWvxQ4aFFeSo6TslgVQddQvcgicRsOJGn0WXCHsu1mzo
6yO/MPu3d+b86rXhlugXkAHJ1D0R5l1gzmEN3+5TUqS67EXyzFbkwWkhHzu7KRc/
Cod72XhEiphpkz5cOcVNeITAjngIOUnzOh0VKZV/M599/Rav3S2XoJ1+DU4vnfL9
TBpx5ATJF9WMu1RTMH0wsWvvZpl0IRQ6ovzNm9VGRSYOqDbD7a0Tt+3LTWErwjEW
ip6Dd6xyzwcXbhHbw2BPWEGFsqNKJ0bXHaZauxghrU2brv+wE0S7/Yb4WfZKNgUZ
5uJKxwUZu8ofg3yUXoM6Dbp3M2VmMUYPAcFNCaUxqiidti+JOuSwcUJ7XGKuhJrU
jjOfnb7qaN9xbdXcWFgoRSx2ptzmL+WGOeiJYK2M37bWAFKjb+YE0M3pyKdlOZV6
0Nb+BqhOBqsfaspw70JEw51XiJWyuIjgJ1MLwJWf6WQwEIK37+w8EuSV4png92ac
7ZTcO3PRHd54RvEoEPIF4a/ImjY9T01tOkwZgo4IC49r7HnTNWkBt465r2qI2ztU
WfL7wHt2WJ2aOIwJ5TljHoQdnW1eHihJ2ckWo2We+z6dphE6KX0RINW7heHu5Dk4
nLKmLqkvt9hT+p6wvQjWh4YwqkcPkjUP0vFvlLn5ev6+Qjd7Z4/dyHy5HayF8wqB
tvvuSAbloS+UejmmIEZ7hbw96K+vaZDpUFEfWFOZWG3G72alx8cHb93zdqwhoRbR
gmclW7ccE5m43uQu6F7Aw9ecpJJ7PguoQshiAYhGLjXTDUHYilvfTYfY+rPHIlp0
/+P8Zrcpvw74VqGp4iQ3o7wOsCAZrk2iY2C6xwVhJfl4uSfao6r6nQOYDvAQkiW6
PYnpcxdPtAj5QBjwwTooYOElcEJu/BU2Ux4q7iubwX/kbBpgFbCj/uCA+eXlwBSo
yCCYIRWUBt3WRZCoi4dvBJZJ+Tcb1BqA0hkqKVxldVsrnFodXMcvfHWI4A4OHpCD
VeDN0jS1xbygsc7ZzSD1mEhf+kD0sjxMjxfBVFwqHtcBgM98ddEb1XUltrEZgBDe
kJzypVkShKWGHD/bqHGhrXJxpV9krG/IrnxHj1rv7M8mcYyzWy5HkUON7KVESX0+
m7VVySPq1pvoPbYRP+BIlB+5ooU5bl6ZxF0rCRjkB0kBNHqFr3935ZmXdU3yjWAa
g3ootLtJMNBTCGp/sRpaEAVRTxdNVf8+s20xbkrpT7lnNUJReKEyjF8iyRIBF4Tj
1r9vYHMBmnirl6/9hq2eepk7cTOZXFes07jym2YqrzCuWMq+9d8Y5OxDhz124vVR
xuajOQ0s/EEoQPoPgey6BjmKIubpNQEr6Jp82i0lhYvq/2mdsvirgV2+IqG3r9iv
Du1Bv9cVNROKqerUikDQnUmF8un8KqATq4vFZN9mybZUuDvvGUwtEmUmuwLShbhW
KNOOMQ2xdtuqQ7Esziu8pzJZZKPNc7Py6MMd1LCd6o+F5alEUuk31yp3ZOZv+kmV
1Fa5vYrR9nqMLQQJ2hK/n8CoT1XQLFfazBLI51WXobolaklqnIZFkBrgCGtpjkaa
ndEwo4s02XHOmu5nto+N2DIQaHiDXWLXiuooQmSiy2H2mxaAee/NwcMLfmAv9tTY
nBJ+3Msyl8oWSg+HX7ZhW8hlwsihlkZ8oXzK2xTmWnmxnzE7mvKVzGwYoIcLBgKR
eGgew2p9uN4v8FeT3TDRRSBdhWCKplbqjW4oEKUZ/yxJhaIhVti9yG1pC2LiZM16
B9hRntrlCvP0fBjOFnpI4t34dCXM1qFYls224hutxFlNPmZol8I9rHoYS6gEwpci
jK8tjI4m8aqlJR43/9w8hyiy9Z/Pv82AHvOHL2r6GcYEgl0wqa63hHFP5MacpaeV
lWDAgkA0ZKrMB4YkBSfZqeJL/0GdpIclW+dhi3js6OewYoefqpQKFrsrBYblrerx
zby7yTzcsTA1vONCgiACC4s2J2z1NVATwDKFOW4ahocm9WL/MietXBctQ2k/tS/r
CfFLnsUrFNrmaXISMYJYxgNd645n4pNZYuYQwT8PTjxEY7q/OOg38ZlqHqVIXZrn
GO1NMpOldjIAppi1nEz+ljUFVSccBKq87HoFDhj7NhFR7YXc6t2NSM+u3wQZYMdt
FsyTrKdP/RB6mYGg63eZRecFK7gpxbGzRJtQyXF5c073xxt2VNVcqZFTxWITVNoE
6IGX1nUy5pw6zyDXGu630O51yHF/RciCL603MwSQ5d7M2I5FydtvpcxOLS49/fVY
RoKqW/YQl/VzIbsSLS/rtiox8+Tc974bCeJGz/LRkoBQ4kCUt8zlY4pwZC+l686B
MQwd3W0Dof1zdOGC+oLWhjwyVgLcp6sdApO/Mzf28AcLIWtIm4dxj/rQqZ8c/UPJ
5WqFokjXbyeTs6uoNIyIB54c3vacOqSyZ7GJ3giXmYBsP2VyRqy9Hx3maVEZ6Zik
oxQNTIyetiAOt9pFP59rxtEUWr2/gN7I7ecAkK/TFONjERAdkG9d17h2dYedcjHl
5C0k7ynVWFW8GHbC5AuJcMmGWeOpwKm95kexs9FOZEeg44wiJhFyY/4uzdmuv12f
8atJFggxh4+/Lwt9xEPTvPIKSjZILCL8wi66d831H7uJb4axw2gKN8x+K11i/jtQ
WYFqSdpHMSMoXlsz/Te23lNwITvXQUAkbK6VM+4APZpj5kgUr6zkUo+KlWVmI7q1
rTvme8CGlqulvar+U0yZpFQrJriBuT1HcnKXuYGRkBgq8tT41KNaEZ/bgk4PyqCT
IjM9M9+GGwBZwJdjVQ29HQT1Dif8dyWYdphpYUMWojw5pt+un9ZPdCRFIVnNQI6Q
VEnvyehtmPXGdyngdaEnrmLb4+UwfLeHOkw6A/Ir2Tzx8VgksAybkRy5D6Wgq6pJ
0Jyooaot+EnzRyeDl8oiayaQsO0+ePv7zGot3f4s2dZNlNZnoWcWELR+a8J9UoEJ
tV19aLyfm10myE2RyzmDELRpqucyoWQfx0OPEi1sg6zvYIP2ieaIxJNkose+h2l3
Ogj//UXJzarpadlSMM/iNi0XhnxXw6/OGOsDda+En2xwSydr5aOuXSCSt9Zq60Ak
39NeW1J/n61wJ1JvhZoRi3f1OdSWasi4yJLtQVLYKAkWXBw9O32wbYt+nHKZSukz
xab0lOD95aeVhH+7LKPZj4NUCd4U5PEp092Lc0SQ9sQu/vlmdpKK/Tm0KZ97Z/AJ
gs/a93B9cgRBasMGk4gEZDLKXRjcS/6XoSTbiQlh6/TeoKWFdxrvKkk4o37BEMqg
+xshf/zH/8vJHXl8fNp/QNbUCoF12mKGs8lWEpvm17p7FAlNhQRuYFwa1rF4YPh3
EMY2WiFRPQvQAAWoL1WV+BUujybks8VhOOuXbITAiZoAfbsdiv5wXmfDuduIsNF/
dI+H9KRt5qsbWyt7X7GXDfmoENX8umgmVJ6lRCdbSGQIjJnkhLGoYWLzr0hQvaCq
6rYDSuG2gGMSvfk17wkVGKXp4dEANyKRoOqCcFv41GOcu26RjFDjEKs/IleTFi6H
YX/P+o8B2zGRkpcJchVNUVIkiC+wnchuDhL4f9i8YzHpJSfJSJQ0dxjpRUFMfkXb
FK0OJJ2zyH2I0B9WnXLi4Vf8aNI0jl7R6JlzZkPTAwtRwmR8n22XvvsAxLYzrVT1
PcmrGutj/i908nRDQyWUunOnMJvpXEZBuBc+KRbqJFbQrxlELTFxHq4+vThZrmqv
xEnM/nY36fThcgpaNE8C0cfSNZ+79V7A+CWCkCTSYcJ6VctsHbQXyKjSe/IqGF8V
MG5NzFcua+YdGZeRdZL4jMe53+Y51QujF+kOUf4HaaEN9O6D0ppTDKZNLQpHoOm7
tTilVWIIhT92EgqX+k3VJqMdfqwoQEBf9VgH6S0pKJeXaSqjLgKmLnJdP4MCPBn5
s5IF7zns9kBfmSvU5yCtVLMq0NsHMXygbVORjlZ85Kycc7MEf/SfJZ4pOX9ni6HH
UXZLJZ8kYbzMdg8sBAOdjjz2JxL6DTBIqq6FSdVAzq10JP1JK+5hdhlPhwN6P+MB
WQi8v8A461cGFoAW37Hxk9GEWUb7OGQ9zCaG/h4QI1caH+VMTuvJkljFSBZ6C+SR
MzvtERfBTHVe0DowfSG3mFLbqVC+9ZEa112hWKdMPYEXKcp4VlHDEzi8dpJ96rRJ
7yukHq7y5XcvgKZEV99c01zhvsuO8nQquGojWEJI5rP/0J9kNw4xFy2b/k96Paji
1IdYtWQ/v4BD1Ob8WJnMUO0jVCPbawwjX1FBGlzDUwR3Ns1XbVSyHpkFmLJib8Zw
ihQybmuwtHJdjh2kbaRcIVImBZ2Ylz3UxlKMSpiMALwbsFfh7B7oQwhELuNpUpo0
aBHoEk4vOXE7+oLlNYJNINEqcBSUvuWscN2HOR/cgvhNYftNhwcMWVe/acSQ+1k8
8Zq8C2lc7b4jqFwSGLOddUJ4lBEJW1nwsdv2ac/zx28+5sDnHqi9eCpxCEWKZGBs
NSMUCzfoJW4PLzrWzejXNoNIhsI4+PJqm0v/ox57/AACctNp99+ZIr4ZHuxHaVbo
aQ+8H+logDqGo3en7NlJLvIzeCCp7rDdBtbw+s5Ok9sdAQcq2hArYaiq+s/FzTLy
4HmZHhww0q85npUs1PXA3BRb14+9qWIzyendRpkP4EzLojrBJzIBV8rXQjOmuZ76
cBZLksAo41YryEF0SsIifyl6ofU7X/ZfBXGVssWhmdRyIvNATtroKmzcl14bXZxG
+FXvbU6YS7p7BQumz2OQryV+H0WX0TjQC3ExcuDdTAJFn9RvjsBZwmsmsP79YQ7g
Z660HNSy1z2XvS+CML2XjVrSDyBFCrd/F1yBnbJglwHswvWjfg81c5CVRtIYYCgT
m6+hPODJsitl0M7k4CBU2Taostm6nSIyC+1lYLz6YpZjfGpds4kYgN9brXQXEyUl
4uS+bdJRr8PrkkYH9822kyngOVzjvy//fP22pfCRPRK98pUw2A3cDPgp0tfYNeuF
Qmec9nj68TW/mhMbaTV/2V7rJmNdcagucwEn8HrlUqZMSePoFgC5FjD+K9YykBJP
q4i/sOaJW1Esg8jczqWEGjzKrHmjwuQFNuuiVIUJr06LH6GNr/YZI4L+8uBOVcYO
5RGpgEwLBjMCMvW+rIsClJzu7GsDzOxSGerBdbN59auwT98arNZeoOQTS/HoSS+8
cSnbyqFHcqGMo+4Zo/D363fBeHJDl7vNvaCStYE+6OgpyWujbejkGxNy+1XtIjSA
B8OjX0oPS3RqKE6Uka6Hjw4FrOk7Kf8uPw+C/hXGmZB7VrR1TVqlyPPOfZFe+FNl
YY5zpipWQDl/OIJrCL+pK2SOIpc8hlVgDGIwtNP/ghKxHrwby1lsCIsNCXmqBU/m
lIThqgx+NHpSjDRIso2oO19jJpuvAVjIge6Syord5g5Ggr02nxocOA6/LBtiJOFB
oIYE8bYnC6kp6oGnN1ynbF9OSqbPy6EsWSh6CbAv8VdPq1UsRCGdEJQ+zKQ7Nh8y
Oqp+MlgrpXQDGC+yUrIRQRkceFOmaRKnJeVeCDzd7Zqs9LrrxiMS0/Nbg7ilwj9+
whaXosB8OltSqOJ04D6smnHrU1Om2vm9T4bAUxzQlLXvugGcf9bo9376Wj8ol5sT
2yymENvxrVCNWA8X0oLZ/eVNV5S4J7A27kwc3G05w5mb+CJW+12Bf1fW51n/03MG
SpL7DNQGZQ9OrlLBFO631YN6ztk6Bzzx13rxrtJiZbbNW9qftCmrdzrEMtkBVj3+
alk4sTwgweVQGfA1hU7hQ8NK4iu5UafSPmDxYWCxWz6OENBUMNVrIxxplW07Odhm
lIdOwnt714I7b/RNBz1YP6ZNjIOPJFIlJFWwUTluB15+ddSwL3wep1eACRlujppG
ic6XfJYpgeSFPDJBGDx+Odn+ot2gnvoM/A9KwwXf8hIAteDRr/zuL0j1pWqlLx90
1cwK6gweEJIoMfFZ5fadRP73zKakQcvV2k3DG4F0Nwu4bshPLrxKnc7aN0XUBSr8
o/6DnbUttRBcxhr+eLcVt2HTLMkp8o4wDbqw9vfiw/yTvbLhmM8Mf8rgtJlAoIA3
UIIe5PWD8u5rScQIZW7/ofoYwIJ/aSj5rLroCKn7Duq+eAq8Mlz+QG61XTl6C4GY
75b5nWD4EZpj+POfc/Lxx+4Abf6gULBlug8E4YoLudiODp1FdD3ZsG1s2RBW3LU/
UbnKeZn83YNYGmPJghAB7GcbUpY5OgBRxfgOhAcToY8OkngfXB3gHwhcBvAeMJz2
hiRWrgq0QV9dKXxoKe+Fg4OVuBLf1ZyWgR9AbnjBSZUbuTnnzRDNsXzOFKXTrCXz
OvGkHoU9TA8Lzn53w9p6L1WBGgeS8vhmogPpcGmHsIf7YY26o+TBX0bQMx7Ugbii
wM/rUlL7OjQ5HNAY1bhnSwJ/Ijrc16ZxRI7jwUzhewS7Eg3fkBbIAsUpYrQphCWP
bwgwohpI7BnjNB9wwGKUi1aZuukyI5nXOGmNZbJD6YiC2kB0XQChPapi2V7T8Bi0
VyH7CXEfryKHkBVQoxvzOStjxNaMVt6fGXJYm5SzzhCNFdZDX6nWLWtJ0GU897uA
sgTfKDF0PfCgq7MfHlAxLlhVooBYG4/KTx/uIted24CrMTW1cJr4LazQSX+KEGjy
EMXI9RRjqQsgsavhxk/mv9EE/eD6CWhcVZeWD+tt1dtHnhF/atbHs1JpKnzDA+XB
nvOPAiaGlSc9EjqRKay9TcCexXM+vDvZ0/lSSMig/U6EfswwzwtY9a7k9ZecRF9g
LpNX78bXZnBHxWw1aoGcRikUIypEM+FRMCNgZ7/Pdpp4tenMWKbjoIitsed8cfr2
FHDAaKKwIE5xZYCUbahBBQdZKZEyqb3kaB08j3rmOAyfKkFg+gJ2ocDPNlG21vge
mYLOsGiW6/kt3u0wQ0WGqupaHMOSIlCXxbJBtm4O1uo03U7wHcZYJx6LUL3OGQKM
aKlo5ZDl8Jfm+B06egEWfYVa2r9ADoZ4Wn86VqIjtmF/bUquLFkUrrkqHs4qDko8
DLqL+lJnrnkqaDYhxRSZzAFo2F8c5Zzrk8c/kS3LpbTr7Sevq0Vd22PhLKcY7Pyt
icvA5k1s7kHm9qGJd6eYRgRaDW332yv2XECCFWvAF9BxQci/eObHUeoHXQJDrZPF
V76Kjd5Uh9RZdP+91G2W+cRtjUNAVJhsBeRcw08TXq3Qb3YXZBitalUu2Vp+xwIX
b/Lvws263wBFSVZNk7QgMaGGWcJMpbY9uMtn6X3cZsmthN6G/zsenurRLWKru7rU
//lET/duuJC5HoOo4qtf0rkDLEskfFRiwcxZLhMzLlmcxiDWYzfwSQ3BIu/qyU7u
teBYiLUMqIS+VGDL3ZXoVXRhW5eN3zkaFOLuMEapqBCrDhWk9rmwb3l48qAfDYKk
tqhTxYDNRMnp+yA9VPWCDYfXkxxM4YrGFJrT5QOvK4vTbbrHzhZr/hkQKpYg3T6K
JKP/kIEnSlxNNu8AsnNJnuAIGk/IUsEPXK7OMGZz1OTXaWrLougJ5/e5vz1XcsHR
TA72dAgGbNGwbUSBrDB+IZhaJVRt1vD3gR/+WLd0qSQXtobUNyJDWo4mEj9KNbXE
6q2otbnumMluH0K/BjXm/24Xovi/xiA33/DQtubWbYvuezv1OvwPaCXGPep0c602
tPsFKi5WLBGq/0s7wvIwYSPLLqblgzft46IIbTD7qGnhv+qO0hoXR8+SlBk9RyvJ
OKZ7fe5lFovebPsMdOM2WrZ1vG4L4uUR4mMVaM5ZfMgLbiv7uN9OcZHSE2+AATRX
CJfcFwIq89ZcFhBaIQum5q5wy5FEk1izaUY0YiS5ZHREkUbJntGyeDZ8R6vYttVD
XAfov+b8y+DKHm8wpI4tOuuXo0zN1RgJEkJvorGJy+FT7WCBdOx9et05qIbloFZh
xd7EAlBlVeEZZYAGCDMungqGZadsNjqHHnUxIBxWU86scOpUsJI0Ng+sP0FxZpXw
5Xaf/4Qq8mOi5AQQavRQoOlqwN68I2bmrgDTbX8KWzE7fpwQ89GW1AwBkCWQT9W9
dvlHCFc4TVx1AnLbdKjZZSI96sPYK3ALoDBHAp1mJm9feccfOMgKgSslA3iN1/Qt
jlkB6Wl1ZfnP8wG6oQOVjC55hHTBoSmY6hwtrGIlGGU4IH0cdqa08TuZsOKqMck4
HXpsPFu4MpVSIk/HOxGKdOGTFnm0egzBe3toQNsK+eU5GRTbOX3QnUd/YGhu3oIT
t/88yG1JOsvUnI51JsPCDafKi4VtVTiHhrMciPvIl6EsmVSc/T//cSh6V00HIiiL
lL+LtRCCU9rtyDM+1WHthHugg3ZQ5UL2mrtQm90eHEeMuhN1p1XR8+qex5ml0l5t
5XXRzgmE1ip+URKRHfybnPYnKsKG8vreqizcM128kZbgFpUFt7zbRZMyn9aVxTfC
dUfZUhMkKfcRlutLRAqftqrGoQ7UNIz6C1nv/85M5PiVD5GhLYCnrGsorhlGFhQW
eD0+zmLoJQhAoXtiTVRxXlakZu+8j3gNNAPzsMN/kghE+Z3rqfQlCCKpjUcaEI8q
Gwe0VFGxqQph1hx4oYWZgsNthkdQw6LTUU1Uw5Y/vefAzxyP//1MGCdmF+khEk+x
bjZG9YgmbiotA3m7pO4G58HVtgfvi1RK5TeJIO4YuaLFCyV0DMWM2cunpaCqvzAy
C7WYLKmxjdQfMdHQ7Pxc/LefNVNlgAwfQ4PSOXV74I2ECIno9d/H0i6eQiujw+p+
thretw0zOpUnCItIkaaxBqfIZrluCJJiH3B0p6pmiw2EVgikIub0AJG9Lybb5HxX
01103BblmMWk3hwNIyFjSwHudVWyZyjv3w+8kXrd03LqdjFhiUh/1HfXnXi3Tex4
p5Ps0C2kHgxFrfqB8rMIKsqTP6kTo37/xPGTBlJYorZOgYN2rtM+i6s7hb9jZh3M
LTrJbD8qacEqkE3XY7NdenacYY6DBSOeQfzqh9dmjXVsrGe9UsuGGbd7qS9RSv0+
BqfQbEOJ1IrN6/swPFyacr5tlw3eaUc3PUL7/07XkzkIjEuA8B04tUh25rmRbMjQ
6bF/ylh/i8G4DBqpWUPMZ05vcaibmuL26DPG7M332HzAMSJOV2fVBdE7PeChjyhK
IOnybb6XkrJEXp9rxbDync70RowVA/3PYT5D6+m0QIjTBDLhgdIC+37YmlsCPxf8
3mfcRAvqTCkFYo6vb/EHy9EuSpzj0vSu+HWoDAGPJPZKHQyj+Hk1IdInexKIBWcp
r4U98O3P65t8ifAWhSvQ5m0e9/5UxA3WZlujllGGaBt62pb1Y28Ana7cMAwYaWgf
dz4VQdBixtvcq971nnuAwBUHIC9mrl7raEgosJbtiomaqp0b6dmtSpJdjJ31x0Sr
WNmjRlN1vVTAVYMWe4bj3LN83EbTCk4DJXePjQ1YrAcd1NGdrqSg70Mr5L6QdBKy
jD5hIuKF+xV9QPtuv+cvuzwusi8Olm5S7ZFJYYGHLAvfK8AWrd+awsgeqget7nGQ
HKn6ZZhy52yhWm1IFOqsgL+mm5XEc3clk5JGB88FjRa+M7Xv743t/ecO6p4wbEGg
Q3n4+2U6sHzRpJEb7O5FAFGgUvqkEntWlbrWGDgK47AU3W7SBaoI+PTTCXbxLCrc
aOqTfphVBhRv7PIJRyO15NQHO8NPJwl0yRASpSuTowzyz4kSg/bXVD0MFFPHVFNi
DTnjneDkS68NSvCCLEY81ZR4TLjsMqbFGz9cxQ554pTmX1yyZfPN9SCZ11WMOBAU
z10ARINSwAZbMFYWrtVtFMW33jG6hZTmNqmEg6MR00S3PJ1p0RdSDohRa8zkFeMp
tytHIyFNutoH8QTbfRV/NHIN1Gt5XKj3VArC8gIYc/mHin6eV8J2jZzZwbyb0xAg
jKg4nzdp2jI4099IlLoiV03Nz5Mh75QXikasKNcPMR48U9csNTF1n0HqJzkX8kU+
5DvxvB7w8iLcyxsrW5Hw4MkOgTEsBR0E5gHL7mWWGfWUd2XV58aXylpLTrnK/mr0
KfaXmoHfE3e3JRWHj4MuwLel5USUC3aCl2DYwXFlyiOkYErCZ2+zK5NG9mf7XCws
NkdMaCqABjMtRdjgQBdIeWCGssr8qIqE+Np2n7m5Is9/PxY/bhwQdIIEi75RddpL
Opk+25u+t75J2qjM3JVf+Pt5hoRaWmV6h4e4rcZND5WVcS3Egvb45Auvg5Ax7eBD
S5gyISYlCO7rwxej6JU8PhTxEkrj2+CIyQ3fHhqZhdgIcjT0voqIk3xeuSNwXIxC
Ycva7vVmEyPdgwmeowKEN43C/qKN5Xy5wrGWrbm7CF8elPKDa0VQyIz1DiUtKzMs
PimzPp2avV1Npr/EsBRfFXNB5pAp5HpA67vh6WF9jqR9tqnZhG07dQsA4Ocy1V9s
PJN7KZPf2MdMYVez1FeT+MLk9d+K0+1Iw6qy04N7Ev+AEvjBXSYjQwS0pLJN64pd
DBCj3DRKkdyEbPtw5YSCmo/Vh8GM2YXf7G23bRLAO8sB0NxzuBBeXg5XXhK+dq08
jyG8S1xd5YJ5DrzSHGsFiLQC7kk4f4MAI08Tep6lgiw+ruSPHUwzyyZc7AsP2EJz
oa+xLzWwY8dJiaM6pDhTzkDYM6Cv9v7lymipXbl9YdOZ2+CswwUdC4eGuVGL95Ft
N5gph/mk6RKIEPBhUztjFPcpJTZPhMdncjF0IeK0uzttUTmYrrJlGD829oGDmfS5
oQhJ49HuncJcxwZo6m+6qCr3r5sL5zM2TMiQ3dlXCq0XRIUj0Q7ynm5qHY9cjQpT
zXRUxypk+oppBs4TOuj6/n4db6On771y7Uz72B7onn2J1tyYqcZ/Lba/CLsaUm1N
A/18T17UNFkX7jbgJSf0ysNWpBfYszGti6oSYFA882AuCsNzZHCv80CVIbXVMZ4v
eB/ue4WNlrOrif7z+VSFWIm5T9aPpi0KSHJQjjUvQHEaIhLM9/M96D2FMj20AG/h
j+7ab9jgpp/Vsapd9whZYZGAW4PtUEZoqJNX6VaLIayPMd/+CSHTFo+Yg4jW3TnX
xJg+Pnv7s2xYMjIF3IhewhrS9eKbyff4HNkdf9qJIfka79+qvZqV3cJLmVxIPhP6
aTbymgig4GaJVNGoDg0y+NK9Z5pUG+oIHaZtnHwhPNdNi4U5bhr2nUOjffMNfaaq
IzH6y8Rm4oaAVV7JEVvG0kZ40KZM2D+ak3G6f5QtiZGvLeKuwlmvly9HLVGHlqKz
YpuhQB/bUKVUqOeGuq1OQvzfGMHv55Og5RRD/GY9uwo7xSjV+SoU7ylPCmgoPyYR
CGDwge1O2htnxr4zt/g8nvNAIfhw7A36SMFHkdYfxbl+W9YampjthPckXnjV2IW8
kTsP/g6I4mekj8kD1udtIad/OKWDhYWx80AmiGU7RSYY61aXfenYMPp+4EUFGv80
nmp9wOuuoiANj+7t+EOQ870+SRNwv9hnqw6qsLiFHH7YYkzqMhhzgT5rcE+tdBd/
YyVwwIByD23Md4Lk5uQOCaWOcnq33WPpFHHTnLlFfezeyGsXOUUNXIEfkF3HOUP/
c3yT286hbS4Eyc74i2/aqqKcOXgg0jzZwvAkR4B9ktKj3yCAXav2lY75z9ZOtOv2
F8FUzcQk4MJtZFaLC1Y8qSkB4JQnzy6yyai9p7+PMKhAJN6TWmriber/qFFGgVDO
rqTRCP4d/3kYMSBErSiQK4xz2l1QE+fk1vQkX3ETOE6JotlaoCBxWeQ/oFDNGRyj
p+UtxMm3jGMUdJZ+SS0qBeSG9SKc7BtGRvEk/txoBkBsun2YvXQIyoGM61P2hLQb
9223QKYI9bxN+Z54remI94HDNjbJQ0B9CNTLqBw+ZFgwWW9HZhCySNBAoE1ckKEO
22BX7Z6XHsDDlVTvJnuc0cQODfE6Pae7FWHPY7GusyeyF6U0X8ppDdO8U8l4t410
PwUsjD3b8BI672iNmzjg0l/u5L059Zyfs5dobF27qotXhnHj9Y9+BdNg0GJPtCzl
9Z2DDol3eL24sft/XD2fnklzHWYtAHE4qUEYf2oghUI7QBAn1enegWw4uKUx6s3N
FXaS7ucmpYBlmPOEbvM2AL6Q6Pu633TzoulMXJzVQF9hIFPAasRogLMCprkM/nCv
7P9yggpFp5S/VMjMx7OrZK0JoZ5Hc/ZOuFOhtwe9OI9ckgnTr+aEdUSLrOCbmD74
2HUfJF9Gwgzi90V8NkWLixOR26F2au8fcwRvq3w5TvsNyVK9z1o9aNcPvMySG2Ph
N8eJbGCooUZCook9l/QdmlwAR4WdPYWNRtES7BeBLtghKatsZCCnxEFkKXxRdGYh
d49EEdgjMZTbQneavjvXXEDhuxUjAoEvGfSNobfHCIiT14dHwaXcl1yaiS7sjzHe
JBqNsrLuC8pk9SLq19msCBeDSv00QZ/HzCaRB++VIO7ujI9uU+sZPRldaykNN3F3
PRSrehqZwX5eGB3rr00hZFqqPIaPVWSTSav6WfT8iiiKdnRAVLyybfW45zX3u43s
6vcpeGhA4AKL4ni/rgxfu1RRggyb2Vt/ewekaFyeibGbGLJOFX5T85xSme7cDNRu
8P/Faaa4sJ0Mhdr4eUX+FdvFkXn1fqveB8ltHqpyyCo1fienyScKv6TDqrdHGzWM
01jZF1M3Z3DSSuzi1ddicAXpnNWCWVGZnUDef2Y7kXlzZHxgrtEJVbenbjswmTrY
QlbZxsZvHzg24LigtNHUcTch9ekWJ0LJaq1JScZFwQxNFBzv3ziKx7KA8xykg/hR
3Xmt8uWOUbZeptDU2AUV7TPDCAiGc57Pbd5/MaaU89jdHrb28kCgbv4ooeoKFo1Y
qo1BceZ3pHC96KewHaBKL48OTAVXDYS1WIKExrOnHLECGtksnonis29Y+gIIcWuw
p0vh+Rf9FV1fga2IbyBcZdXyNUebJB9EMDp/VjZcQwL7g4Y9Q+zH9foeKa/cOg4U
ulaql4+uRnb2SJnO0jNwMQ9EWXUqXnHhFMwK2h6fo7ItqtUXWk9jwg2Hjy88pjFR
yo0ijdbrP+dOod0keFErBJtqDVkNn6txXYg/U4DLZn3PoatCTqMP4eabzE8OvVg0
3p1PdB/LxSpgu0t/3XZbmUO5jMR4o4VzHypx80xumHJvfdQKBdkSvRAY1+JMH0cF
zSww51veGipHQGsvFfg90dVXaZqqLL2xQyNAeVPXvKs5WEjgqPkOD81EUDYfE/aw
BBffgw6xfDXsKeMcj8x0fGa9SDDP+cyMu7NrQXHqADB2p2HV9J3133yoSxGH1bzh
qYtfwyBMji7uPYLNOFDuIzSRSLpymWsdFeIk3JNJIokcY8cc/1J0m0aL82acT5cW
c4tOsfeVr50TIIr4MuKH87DpB66D5lQpQqVdJX0h4Won4BsOhDRn1LZXSG2gL8KP
vFbX5NWidLOXyY+6pr2nh+6ZlMvfTbZ/3wwYIEqrApv8+vc+MacjPwt972p0UHZH
54gDJDtQkgzdPouO1Wu/8vqVLXNEtBHwggGMFcLY063noT0UCrE3E4b6mO7+QViD
i+Sv3RoKIyJyJQQi85XC/dl6BuxPL3ydgPgSBUU05A32g5mCr6SkzcNxe3YQdBgM
An435W/0sl0bwrFhYFWgC51Q4DMCzaCtm/Z/pidQBME70VFY0m6z5YJ88y8G03m+
orm5wiVNei8/1JXmrKt1eif9/m1AzsonahVtKpdPeVLYdHYLM0ST1M541b/EA6gf
SC1xlCMIk7gAZau6Zk3gurTzOEfgHNi83x5TSJMIofeLZPbft0QkXeH/uMDTCUiL
ZZ0qJ7FTlikrYiQ7KJ0tOs5O9hkzZZ1MHiUvlue9S6wlOXYpICGlJ6V5MRcDhC4t
KvC+mRBypcvtcD3pJQy+YLSS3SyOAtYhA5pVvOWSi6JZNZxyGnqtcfmvcVLygeYu
fcuffd0BAC2ShBMJGi88KZqRs20ad6ZPz6bTyrEugG24SFUXxfWsmXU8X/RJMIjF
Ya+MsKHHMVMgdUYHYUGL9RH1yhXsyJw9WzumqxaMWRDN/xA/xt2I8Z0jryrIEaP8
R+f8lkjcwhQEsRabpsqEUJfF6/N0+PdWu6OWeZDWNFzW/I8PDHi8CXfwVa/TjJxO
Bz+PSrlBvhmJIJM/xGDh+4u8kOMAsXwCCrefPa3kh+u0E0SZGzMisNrSPRbXO6G4
NevA9Og1tc1bz1uJRO5vJtm/RqbPZih+rKMxwP3yYIBDlbNuF+JUBDycckhA8TIJ
hsrIeJ0E152vDVHUYSNDuKhPIm+gNs+wIJT+3ltHH+fBqUeyARkt/QDFR3/icP5c
qv3E0UMiKpt5U4X5q9St5Lt8rTpF3QlK7ZdmoskHr0LUJLEnbX0bezuUyh3WIofL
gRM4uRdk/oxfHJinQuJ8w7EzkwMndFjfCGxQ2naZJR3gDB85PdHQRrr6QRVVW2xU
eMM2OrVI9dxmVi4EAjjQTDLolKsJiTibcveMLFekSNu5P3Rhpq5zmWfQvjOKGgIA
Va+FNjpnM9sj8N0OulDcq2J5QFbddwANzUUcSoe/uNOABeNnhg6fXAuPyRNLlfl1
JLn3DXwYBdUWlXwTMsQU4AVe8P2NoBrqukRdx4A4Omby8dIbczR/lHNB4psSeNut
W5jBYBrGJRkKpd1cD+j8smey8ne9FpJbA5tZ6qjDIGun9hvl3KwMoikYpzHQWbY3
G99pBii4QY6DGGwglLerfMPGrmsZzaw5X7zqP4bb/LF/K6khh+C3xRdzjxF4z74f
PlBxy8T/yL9zVdsMQU0MSo7Ai8mji4Zfe5NWGJQca/fejNCRZuQ3vZjP791HeksP
E0DPuBjclyEn1K8bch9Pi5i4ovA2tb8d6dgaA9f02PfcIFV5/vq9SL/J2nLnXveW
cXHWt//6oRd4uhC5hmTlowu/GbtYml3RniUj9l9hyrpzcADRPNuQ8w1J8N1Tqi+3
sQ0eRVCN0kRKa656EZBO7Sn2Shej8ZjMSTHSISGZrtCG1XeKVS6rJ2YQqKqb6FVb
o2ydD+tgb1nbP6mjSb/OgcEH/k0zL7nRHe8f8sYViqUqNLkD1Pe4wj974WBWqHZh
XCkr3Tyt+VwblUghoJv58LATOgSCSHA7Ptob3m2br9vS8mlwTXHVI/0SxTMX1Kx6
MQVG630YGQOGzDfj4NTc13GihYilV3nKuDOEwyrfiBQU+KKI+ExKyajYT8AEwb1A
xlK0/zFL0TnuN2ZS1HbYnrK4sfmpJf32Rc+5MvGtURJlp/5Xn9xP8eqkvrFaR7TT
AAqsTn8eHQszO2Z2yJ2ynBGE75uNawp4HSNx8ADnbnDT/gBzNd9i3LKu04KgX24A
XOMTDT0kVDOTecFJrZDFIXi1Oj0hIK+68KBfYlIGaM6G1xQ0a75ntK2hvXEepUR/
hVvCTGjTPm6HgFa3h3BBCRzUY33f8yMml1CbbfD+IhQm+agmgvbv/EWlGVbaIH2P
OaTKO7cU9W6+rswex7+47lFnF1tH+C+jSAyhCLreLTnXm2rmfkoXdhOkMDNWvPzA
bYRp0sBnR9ptHzDqp3xOyGDk9DTOGIdjQklEvRXZ8feCx14htEeEocOL9GOb01an
Vs3A/oQAJ0yjqLCIPDZmbk2vrM3VYyy30OAhTXqsJa7ZCfVrD+QWzbCOcd8bWCWE
qlO/DquTvHjUb2k5IcfOn8mCAB3QqIblEW4MbRtZFV3xHzXmvUSv5EunmVHw4Zm9
CLWhS09ZuFADgwipKY5/Z6ysW0j5jBHESQ+mIfoWP043munlfI8fDQQu4zZ274q/
iOQNqIN3boNECIMl8AAh/M8q+24faeXZexFPjs4AZYR+s0mZgaUONTAU9RqwOyMt
vnXEvrA9k6oGF7xsl65iPSXHl6DohgXIbbOwwpGyqDz7qwL3w2+7k6lzMDaNezyk
Tn1KJa9ZHK78QYgSs8mKkiQsZoh0vrksqbNp/m+FSMLxRUC8tozQOO55uA0NRmBc
+kDOucFzAHW1RDlGnnWldjyI4n/BRO31AskOid0khsWignIAd3mfWnmcTfR3C6pF
upiBgIoKn2rNvQz1CbTJHhUvwK2qvO+q91j+xti6UuolyLME0dWjqFnqPPLvBhd1
cAoBchTEpmKGZMfmXpzzTuPoophzZfldzVKGrq4AwC6KThwhUCR9J2t09RB25xFR
0c4Os8/XYnHXLkxLbcDVZ6QmSsqgsqm5NbbLcuH5XpM6E1vjLnqb1kynoQcx8560
5ncEMSACTvUmYg6Nu74xxmfR1TnqsprjmjMNDz7Llt9jUyT/JZpF+KzW4iCJ7tI+
n7ymNhVnHQZ5r2q6ngDFZ++g8MbpRS6j5LrtZlSfgFJ0aaIST/M3SOhexv0J5T16
mt9RVRcSmzhfINUC/WdYv2Mu1bTduykr/DMVvuhsvsKvgbBpy81kwTaOi9Jqv0Id
xfEK8ppIxSejmFuZtBzLhBb0F8rBJBGuNa7734dISWdCqD+fvf/GlC23cqoCQg0T
ONLeA763V5CXeQJv0BwMjE68w1UKr31YDE+qg50Gd99dnY7FSyqw2BJ32PfeT4qQ
7ukexyPdvH4RnxTBdNXIF50Dd0z3qVFQUC82SWXvDfmxS6FrsE9Bt0qv9GI8T7Gc
A7NbFttzv7dhO0ttOWCjI9ndcwPJF0YylBibE90NPNj+cWpuYOlURV1uRsI/QI6t
xbsIM/q7RySwcKrv63+FwqcWkvQPu+jim1rf63eUfWMR9xY3XtaMB5l7KL0DvOiC
3vCYVuLAQmHkX+aDoZFjHMOdEN1DiyyhiJWOVFzm/kybnPYbVyVJ3wbIn9cZVZaj
vKOgIs91Af8IFsAx1/WD8cZV9R2s/sysCfrYJppe2TNslKk7va+PrkYFxN/eELH7
PNHGmoDXEAeRzDlHMbZpl8RXN9twPua3/CvhpAIoOSmTmFbxTG5Qp0NQhh/xHim3
8eZi88CgVwgUDNo0CMQuq0loANcPjqND+7XSYqHsW94yYSEqYdiqYV44wIZ0sQCW
lbi1ogT488w3au+vrD55caGTki1nRibvetDAuUHN6mGVxmgH5ccB61vY6UbbI6g5
u2z0TDmDFd/60/9fplWEsEDGK3YWfR1RoR4dqMOgsR6ywnSacU88XLlmy5omTLy/
PCKC5Qi63X6Y1F07pnZoPSgiqOpDnl6B4DegX+hPbauqzydzMTcfttoXJ2+xpegc
QS3Xo1bpoM5LtJWeZW7AdauVFb+l9k+3sNtg/lwnPk0C/U5V0+/f0Bw1JhPADKSI
K8c5kcmZD9eiow6SFJCMx0UfFxq2UyU6hQfQVwLR6IgP8TjEPNYcMT0b1OxrkkXw
iytoRVXaPCXf9uhIMz8ZFSpcNjWnqyytOoN+e3FRjcOfMATzIVM+P2wZrhiniOmD
JcjDbfiAtn+vWZ2FRW64YU3q/UxOaLRmWGY+huJ54AtF4v7UyUsIIGveATZirtcJ
gYJyuKGM1HA+mWDW75Uuultba9mB4e4t2CZWjrXB6n5CO98eesdr9uk4Wi8q4pKd
ZWQbAcg9Xbw2E2h+z/GG42fPklK9qJEiFJU9nMM2M78Ereiuju12IS/ytMBqiYiS
5qAq9H0u2miiWzo16ndASvUWKXOGlsjgGFC9h/f2k2yguF3vbqO7iB4/mwAl7EmV
GNbqHw9QqqA/Hu0RfXqaUpeGl9kXk8QyKj+1l++MB25ohDyT9tO7oIblp26muk6z
IkHxO8GsBGN7DMSp20sanlSBZOT4vkM5AhMh5QCitkcevX9kpiZGGN1eqfYZnKNU
PDRS1iG8CFzhzuZbjNy5z2Ci3O5PMXH/j2yl9mUz3eRNjc6B37ysDYQs2rdDEYxr
Ddd0D+Q0x6w8X1kwzZT2URSxQNdUemW8nwkQA2LobgDSGgG+89yyzd/jIHSrAIRH
j/KUv1FOqsHJL8sxJqNoOeJ9w+CXRFKh7/kczAGtp48w+rHkgps6A0+g1Mxt4EjO
QhG7HbRPLXmE2QZQnul34dikZBeJ5K/4s4wl+ObReREL3PBpSS3IdlQb2QH3JgRv
LD2SiKOqDsutLWCmqSxYp5ClX8Ybvu49dpwMIyS7d7xbEQ9rNiimZ4gVvhxa7aw1
AKvKa52viGV60JcpBTE163GGTYY2LF+QiN3CG5l5KR0yn09+gSJG2TbHeEgc3QIn
GP/AWhRD+ysPFKdtHk68umjzc3tVGmQHsE6YcRfwMr2bzx6cqumRhj08HBUEml00
LqeZQcMtah/HhDICfubG6uTqCH7PLJKAjt0LNc7GXW5zzrgDFWgShtYoFVZg15cV
X6S/DSjzwZMPPQZ3oSO9rI7qAreEDwII/44Tni0ij3ULANPqAJ6R9+rkwkoz0PFW
d5KGgNEr+Y9H5mLsCfe3stBgbLBKav5TNG7dRecDRWz3DrJQPAiYdHAtaJwfiRMx
dFvG92xCE/6NQcUGv0WtWiqpHEfDOoS7DahgUI1HI7pVJAdK83VIwA9wb0Ss0OH+
NjJwKovF4UlEh/RRRFNlAP8fv/bXajYnnoo1u7vwcfJ+YXNxx3iC1dULf3ho4Qtr
pCz4yMe4PPG+OKS3VHOvD9V9lF5kgSlXHsvkCrBZks0mAQo3U2gOUJG2FG0+iC5B
z2y+5N9+yEDOqNvwkn0xkckspdG3s2vqqTWifxbVvLumSgv+ikf/cYOPcCDPULEs
rVHt6vQuShr788pzNjo2WeeSZzBmJir0LCGvfLs0EQhrj8DeqDUAdUuqap/KFNes
s/HBJTVkh+uN2jcp4FSxZdIXQ+8V/D8DXz8cFr9/LP0f/NQul1iYzikpPcqWG78x
MremCdJBwcZ8ccPcoHHYjXP1ADwQaw9xtxp7Qf8K3n/fhoq6VbfRC0BOszTfBwjw
AU94oxVbe46t/3rJYRDuqqGbYxb9FbrrVdGKbhBN3tP7lUWdINtRAOFPiUisqJmy
Euqn6dVFr+trCxtdxJHxy2atdPbZFHQDiLLB8rV0kRsDQDQ4eEXqn8Cc2dLIJ3vX
cp485/DDyn/wkbGnreWvlc/s82/0UOgbllFf16RXlidoqbuS2kMpW88dryrZXvx0
VZL0/N/7PNDm0HrefRwpsCWbifr777dTObazow5q96I34Uhfzla2NBMTs2RoghWA
veUZNhVWg9Nz+1JPt4hitSDW2f7rDTvglEBFke7sEN7pwOjzRB8bgf3OUAmgad5A
a2bWpgmZb5PAnNOsCLffA4Y7JBkZPZTvcl6fF2UXqqsfFQB9eWpqMau8WAN3zSRX
UKi3RDI8T6i6+zso/flp9ZOSftSTijfXFbFmFvzVduMxjUF1yWRrbEhccDIM6I2o
RGTTpUueSBvuvf3OdvMZAID/KybP/Ry/GhNWvydvjrYH/f+pKOwu1EHnhmPDFLV0
6QJsHssVu7v1Jlyg9fEMC0C/rsz1LoIn+dvGCX/+QDp0UugBW2HNT0WfK5mopr6H
ZzQUibJU4+FGb9prTzUcLESWxfLWd4Rk4ZTE/gr2PdS1aehprfyq+Zb79DO3/uwg
gKvbOLaChjRSE+v3Kxxt6PnRBsaA8QhmeOylmKweWqo1lYTArFXZjxQJyIEuM7lb
rJu6Pb3BCwEBfwJkXyviYgWuufHtqtC3EVfLFL56UiareajTB8FwPsCpUes9e7u5
vQFqLjktV0SUA2XhY5hltcp1wPfzXn2DrnOG63zliUrS9ZwUMCuxyiToEiyDedGd
CAAYS7UHJrjSVuXNP8GwP8tEpwJehEfO8cF4R2sTxaqPh1l/KcaB+R7yIMcfw4HW
fNp1HrBkOSA+9p4cH/iaUtHWXtFHnW1lF4GIUiNgCu53MJxXfYqqnPcPrW307TGP
r4/lRehikuoVuxN1pnzudS/SNd7l9R+1cAbxYR3k6bEA+OxQtgc1I/pcFKm6MWev
pVTgEZyJa2myRzB19/vhD+rGgq2UiOIDF4/M+uw24kjD/v+JekT6dUYzotiN0Brt
40drIWQiDcWI4rBjIwZPnyRomz+eoYtgCQtB8VjLqIqMXM1v25YRjsPoQjwaG2xo
SFpKda9H+8AggfU4CQw2F76jnvuq3Dv37xgcLiZz6eJsJnEaifM7CGAag7Pt5ha6
zWNyhhV7xmXU9OJt0pgDYagT1B3JBBw9SURzlJHg3pkuvQqQQK6vp7BNHMPhnGdA
zh1ad3D2aCx+3eaK51ee3EgN8aEnHjO2lTOFx+7/wigx4Yo0pfpL6p6+Vnl/qqVx
YYttIn7F0NSEEya4V2XUeyKAEkB05jef40KrjdvILEYgPTWndaxx1pu3qkzt0bCn
suwzlmqxw0VUrHAhGeSsD0Iud4z1Xl1fTavFHsDfGlr5x/fDvWR2867ubmeN/Vck
jCsDYCPa384ehJtFe7xud/SF+lFedXtFPJZ2jquHbbbB/NlzMiBnerUdJEIPF4Ea
ld/DZLPBmcx9klTUoMmzofdVdVs+x6ADmLMdTicSWYfWhwpBXZmLsK0rA42JCt7D
YATRgcsNTU+PhEZ/5qnJt1Du9jeLfkg+SGNFZ2vTamu24e/onc6IAOnwaeYeTloZ
z+Ku5wnCVI7Ugea9ncjKDmbnuIcdb8yMfktXun4kfVY0BJ1waNVFQz6s4wwRjjkJ
YoUDKC/3/PhuZLw+SWMPaaNXkXEQWG1ac/u8MAGm6RqxJEZw2BgMC0QxOB1npnxV
TLspLYm4NM452sOnmYgTfKwuYVmGorJj7fNy1wPXwfHJ4FxCJ6uA2ul4DnWQILpV
7WAfpkh3b7nhvRKG37Je+TncWBdVJlNqrHJa4kODD6wNqDdhtLC+JvWYAeJ0yo1m
pE3w0LLAUOBc30zLmFfqOZv3+4fCok/uKzM3ORVXrpJeFJlYqKZbjMvHUJitsLpQ
ASfYazpIo68QiLhKbh8R9E2B+s9rB3bmW0D9Mc/XuRdF/nWfbTyGyZCPC6jTDbxF
mSfXAaQ6JWNnt3394CPcpSb8uJzx7H8tb0svRMjuzJWO8CARtfyweGZLYY45KJvH
tywh9GH8QZNm761K9kCyKwUWniJzAilChIchKE2vhYeeoxWckeHr3x6c+MROADcE
gVtTpchheDM8n0ol0xOdFpQ8YUEYDga0feRTqiZ/0H6T2uufOVsCnGtHTewjRJY9
gpzsQQzEUmXTt2CNQGLfnW/s05d3jRkLEpmEqpoajEgvXtI+rVOw2Vc+p9Uic7fV
x74jTWLxYwdeMeCX/ffVNbXpX97o+ebybArE88sUh76h+U9m02IQmuOpGepywzub
wiFFFNHUaKuLq7cnwtubXMx5Loh5viTbSR+U6a9s4EAhHrH/z1fEZiHqPuRXQNgs
0wMb3z90VjoyiUid0N0w/URTu4mmeRGeWBaif+I4nW7nOQvqAEdT0U9D3ngGTOwk
EreOUCXwlctLAzRfYzRQszGHrDNtL9AiEKdk68ZGHmVRkYBtcAsGZLV7hcywDE6X
TAXWxsFoNqsFopacEuR1NVJd5Y0TolRICto9VxTwh/jvvBIw6AJLlRw40Bn08cCX
ReufuTNkHZi9NPV+Yk2jZ+aQ1x6sVl16h0GAtf/9trTxzau0lx439zXH2lZhq4mW
iSQh8zQQNQllVFpcHVbJPU4SqGVdNRLqEdUAL2ipkMSL2IzorfROkf42VqjWpeop
ZiuKr1esDlhSUXeJDPRxXpNgd2tY6oYNOgb6kJi6ECZ/07tlGRe8kszD6L4HIjc7
qYE98E+LJ4dJeKI1gGlkp4pkPCXoSj2y8/qHzDNBsTzTNO1Gldy17HSFOA80+cVC
Pa2SANuXEpLZ6CJOkVExDrleM4xj5Ir9qcgq52hErcs5KMqzMPAYdAzAuXcNGMMu
WPwaaQRPAB3AOhRwTwXDj927I167/oXa6w9k720sjRusF2lFRYrTGREzM5yBydpy
fVt26pVgJLKRinBOpRNH7Psc742WJQWn8jqb7jl8UGTi0Tr62OZQlbyXRyLJRe0I
MlYX6AmUNNFlVYf7wZKOUrt2MdIQUOmWumFfVFvQVeX9wxp3zFGtiv7QIjwCgsLr
H1eTpPnRCosppwbxHYblM0MV1xhnZobRD/3jYcRZIVOEz6W0f6SSVVSchkkgbNRF
F2mvZaWd+nsRcDUS3BHPHryxIJ1HdrmiUwC3J+1y5nRAoWlzAhtvBkgskB2zrkea
Mn3r6z6lojUWgTqiUP7pK+xlo3poi+goiuB1BD8xPhjJryep4ne1k3eaG48cn/m0
7ZTSCBpsyiXX2Z7IfCXzbuW+V/2TehQdP9Qz5JPQTsBjogqklA2MLsp1YQJcLQ3m
mIHWYwpC3cr5hgtCo5HutKcUdbEeCzfSseBtBnOleWkfsV6P4zJOdqpwrELNTXlt
E8ih6to3esZ2QzzTHq9F7NJgziaS7D/5QR/xpc9lWYY/okBb0yXFHJcl2svBo/GD
AeQFiK47FQMyz99j2ZKYjnzNyMatSasgpft7q9U55pKL7tFfbFoZGj+VDNWtXm3L
PtA2YRAd5GtH51KvzYN4YGjWCbni0FCjGCuK+mE9W4oI9iH4dqGMf0iKoJ9ZlxcY
AGBna42e/MsdNoRjDonIwIm5JcFFuYlvcNk+bk//BXN46LB4bsyUzSB1REp60O9C
isNah5jB4twT82z8QznCBs/2+UY+VYA4uOdO24lOVf8d+FOWZ9z9AzGSyfpgsphF
g9xl/2SYVTLbR3cepSBqRR/tU0aI3FdXpQHRxsgqbrtnMeMfM9vssUPv3otmriVw
jv6xlxJdBXLW5O74EOYpdjz32pp1X6hFt90oyLe50fCe8A+n1kCMQ1SblKY3SraZ
+5vayTH5qMruvcmrxWwoW3+c45gIALLXRfeccaBcYQkLdENn0aig62GWefa3NmxW
96+ja8H9vQJWIgSmdCY2ExMlk9ekHAwtbxlPyTrGihNxi839l7tZZkI2JZutKrtL
CYDNB42wQJ0ZK3DrCYEatygt3o6fPKi/SA0zIVep3QFU5oW6NXxQmh2cM0AAInX5
ockRXJOZby0e3AVCLQr+l3jCeoaUTLTM4lUE98dqOiNi58kgQtLOHZfOQTgd3XdB
PWOYhQrA33NtFzCoiJDkrK6mO0lbPDwPNv7viYGNjpc53YTrWayfHoVo/RrbPKrw
nBnA5CSRC9O/maX/gsABQWPzmBwv0MUoqpRasuCkR+6/pEdnknwaprKKqFdLyi+L
Ap2qE6ZUdR635ydj3lU5LNh492+tGrm0edXeAnrkB7SQre6FGH+20woaNIEDEhgk
/mOlEi5i7hZHEZ3EheKrIuzcUHeMekSmfjedOVTXaF2HvCkMYEFGq0HSrgQmFV9K
pUoUf3i6xJ1YG5OMB73FfsEkCc1zx1QrwqMjoGZ+J7EMVlSlHg/qJTHI7VIzTKlz
2CVkwzp87vj0wGNagPWvzzl1/0+qUBnWrHsiOFxG+QOcp1QuMPdwhtgEdXmr3y4c
giAWyaHlQ8KjCR9njQsyrW8SoMx9DS2Hv/HLv/AnIhBLx9s95cagAT5uu514JGQ2
PReKJ/mKKYIlnMGp2heziHoYkMSQbpY59aAfR8KBWn20A3XvNuIsrV5WTzyElwi9
nBkygCtQ4dPIL3+h8GmIYqbu7DCGXFazBmHwORsN+Z4b7lKfmJ0YnDobuMMvxC4S
L7CNh+OdxWGZtjiphp1+6h3yo1d2iztwyOY/ci5ktrGtBoXQq3KOeUqBR8ua8SrU
HlRFmshkHhjek9HrLCuE0xORJZ6HKO9rg5F7fVmA1KaaCoKZZQc7uCVuQyWfhtZ1
fMtjGNkUmBGs3Cndby+104oDIXJdFgpekPqLZ7a4RXYu51JHOti2K4pYIociOYHP
bZvRuZajuxTBoO0uIl+HNpprbxOm89cbQS2ez69mbXCfD+gIwNmU7hF0HFHGpPVY
iiPdoQLImCo9u/TmkG2QYSAIfjfofgte9MpNx1O0aZmcf7UDiCcZHqRUrOMaV+jY
xNgZaw45SIjGl0sMDA7jr0gZvAVW/ShVdz2d2VfnwdDhfmSqNWJSxT8bi16Zi5zM
A7cEgV7TIUdRHAeFOCFGhTT0zfowu7J2xUcw73KtzBHjZQEJHg40r/JQ7cfC8HYh
EGAFtRESVVPbU0Wq6OnWbAEm1x4cMQsFxj+HO7sWNgAF4b25RiPakadsTzwpkFdF
rwLHH6kPXnMDpEwrZSZ4HUeymoaXhGR86wkg7HPYDD2jZd/9O2xYPIveyUCzF0zA
KfzVMERmHnhgeQE35f8dG9wNow8HsA0IXKAH67fklOSDY8ZYYTF8mSP22O1ynVjT
Ef61GBwYqpK7Vfw8JPyisF0Bz8TN22C4jYnGtwwkUhRvgr9a242vntAIwYHxQ470
T5l4uxxUMgO0p24SSDktzmIEB8Z0rkxYcIIdRAlWzP/ObkK0mYrekzRM1tHGKQsk
/fLjER68C2E1uq1tqRA8JHHXq80aMJisPf6TNJx42qAzqf3oYafW0071C9CO6b/3
AaHebdRV4220sP88VRbvJIpMEPvo3qnM6T2FuF7UWX9deHEpbwJtlw3Q55B81MPb
844YUkWUSSW0bFK+c4VxJUibHqOAgcq+baFY64zeeFIOXAvayB4pJEH1K9ZmqToP
q5hmADNhoCq/w4418l1UwFvz8Pf/+OaW4CQz9JkQfUMRW2TvztDuO6PPNDJLZKEE
g50RDcRBN+2GrLVToAt6CWinAsjyQIuEtG5VRc5KWSSija58bPcpLoCc5cCMtaHB
F77E7QGKmjH5EoiNdB3bNKocz5Qj5ZyUi15xsa3upOaCzwK8OIm5igjxLOw1ifSy
v8VTppgCuTtEE6gAIhWYd9WX/lussBOpGsuR2ULKNj83V0lFQ5PkTIhAxl0yXU4t
LiCb3BwUYuF8RvZ1tQCr4hwC9/pYj5cqfK/CUYus7DCUEEjfjII1jFpXUlhkRQd/
Zny3IUbwydZsU0nTSORBNZIN3CkRoxdomMm/tybRhmzXlOybFXBTh5zWXm0jZDbb
ksTsZMPezPUQJDV9g81X9J0s9jH2oc/NQdkksHw68TOcWs+S3f7fVDgejjLDV8ea
/t4y2agR+3gIG0JkOTtIKTZYD4RZbcP9pbmbL69wnXTRTnf8waAFwdBiscYFCp+Z
1+6nQMDZWaUyto7esTDEEtugk6yej4ZHaEJzeqEpYEtTRpnOtIinD4epE/gv/cQc
umAFl2skhdFDQFhC3BMQYdHhc5eDsS4spHatYgSzvmgxgbSpuixoLOxt8irntUS0
uuUPrvD89t3TMYu3qQ1Wx+w1yhgC1x6TvB8l7ysYc12WsnKmOhfBGPz86duxlwWA
yFy0fQMejVwdVApWrrYGz8Yy4kKeK1X7ujMz6zYev2J/WdV2hI9LC1u4Cbz8z0f1
hRqPgrJ7vR5RoyCIpw2nZwpyvYwRSU6kZiOyMMOOjyEDj+NFr8SoENBTcP9oTleh
Z4AMzTRJYh0ma7C9po86Ce40binJVY7i/rAUix4Lrax/pX+ULzqzzXWlx+SSeZ5Q
aQF4YdFqNRP08+s5+W6+wmecR+OrTtxkRd58g7M4l6aL0tyxJpTREV9WMiafSz/J
7V+rX3gh8ZIMwi2WxFzWfG2amjbUGLSUJAJYr4UkgXT2mCv4k12I8SMRo3rD/WQJ
pFqVqddc9fT5Rfy7RXr2exFwjMmi8jbGnE4UEQXREkoVVllfvzPyMkCcNADzuQc2
G4Dzkbc7k1sTS51S5GSohL0YTAVvJ0uXhyQbHB2lAkKreg75/tw9pP77MgZfIVug
pNuDz1EVACScje8uk9tFHQZi1Y12cX45ZbatVUhf5sJLuGdkNcrV5fcHp1Kve6Pd
1mFsZ/MPAWANi80/I4dHb2KM+H83qxz8mplyV/lf4AKGCAp2Apno7Zh81MQilnkc
pryxEyRwS6Dg5weoaQBnYhhDz+EueZQzirtr5736a24rv5r4dqbBjzZBjOLS992D
iCQOserv68FbCHqOW8iM2Vt9wVmPfPEzMoPfNHRHsKY8cuSZIctFWFrw1OZpj+2Q
OGJ2GcnPqAq2F0vUO3pRZC6Spi3vkA8+MhoTCDZkh2lhEOvdvexd00BMTbb6Vogl
MYP5iy5vNItOXgcvmb3IUJgxlz2Nt27TdB3bOMZMIeK9xYJ/Yz39oHU4czIYioVg
v/+FK/gXAn/CJ05PVniX8FCTBsCslIYfwLdahALuT9esptdBTumk3cNSYXN6034E
gu+Do/dGiGogbKWj6lHg/yYbdTOSfn4VYPjIrjPtRyUxAcbC7yAP/vCP0hCfUme9
1eqEg8VIv0+Zrg1IWcQSZh3iIM/jPR3LKRMD6TBWYCVg8s9/7LvHSir3cuYcCKtY
SxZw3h4IyURi6LU2Ha0CwVGDPBwkxoUWmIrl1reLw5qDXGGHj1ghjiIPdF8RQoTs
K73NTvLb2JR497ESn6V3KW6YH8iwXQDj4AGsDjBDFZbG++DSCMuCOkIGi7umr5Na
2OO8pEm/LQNLv5PCQGFfEYdG5F4y5eH32NwIorMywt0CykraJOwuCZevjhULs+Cj
9cRq3e35RRXY5y81CybAuZUOLnjTa+l/RnZ/7YRgCusf1PMu+qnc6Gr06PnL9KBO
79pTUgnu2wCEj4c+BSn02stHBbdAaQTH8D9mC3i6jTusohORTgTq7eJRDt0hSgHN
ACTfHet/3dDr5rMf4vO2f1vXxz9KSHxLilOaRekq5P8UKRkYbBSN3pt7QY4ezc/M
NRsrTPOaBv/FxpJAfmivfNtK78AXcEl3pOdrPcIIRraRaLghk9ZxCNLsm0Q4AtOe
9mGqySMVWRB3MEufyu4wVv5jdgNcydjn152BOc6FsfqB/7lkPVMu5NpoCmB7/piU
WP7zyieg45VhHPyKkSZD6ODmWc4tGa5U3EmVybgQ09wt6DJCE+r0O2lSclRxccPo
TNHIwhXwm9xIH/ZLuIObBJjGIFmaCR1D1KpZq/SsJU78IZArng/nXxe2sqE1YZDQ
cpYR3WUS2FUMOx/iTILx74D300d8ITpCA5bnWmj41DbQf9nOHy5WooFAjf3FvPsd
FcTqDwjFj99kJoje8oq9scS4bx2J8hqZRIXD4NQlmQKYlzDUmSpAgz/4sxUMg5HM
2AacQuB0rDXq54EoLhc0YqAABG4ZZTIK4oX3S1p6hFFLA9vBZYUs1U4V9PpdMx5q
5aw6fF808TnSDYl3ChJRZOBWswf0dRpRFEcLw/RVvHPeyX4hYcntfqXjzh4GkPfW
2C8GioxLaWGL/rmsfzggIeBhXbW5I6cHxGfA2t5Ti5SzoApmgXDxhtXG3GPT/P0K
xmy6sgRjy3X/68suUAI9SekT8/QHii5TJEkqudFrO0pBRcbqHY+MNv9cC7ODKT4O
a3VQYHAwjaE2p2gRSKaxbrQaZoZqjl9ZVHbhbI9/XlZGwPPP/0ANChvahHXj33ph
7cIniVdTRfcEGOriFajpdlcS+sEJ1OGZPSkppxSjwrxyMDbYm0gC2JM+fh/PFHP8
m5RCquUO3m+9J7+UJgT/2YvC9PcTUN1Y+CT8c6cOc2r4IHNLg1tmg07oAvXPje9N
xGlhMjHqxKW4HK8Bn2XHr9NnR2nlEKvOH3+SG/XvvGLTk2nJ91gdLMlhH78fIR2G
99vwXTpAUaYFGFJIYv9IAx5nJaSGf9HE4rGt4VS7elnu22IOl32f26BlcAgTevLW
m8+1n27FZQ/Ao/mh9jH9+nz7HRfCVvEPXTA8OXxD8HoWYrZzeyH1n+ajNOoG7nkj
aTYEFD6nQuUsxJrtE/3MSSrz9olxQgnEF5s4xSDR3gCxFb8pJ4StBRP0vi7YPD9v
axPFX90BfCN7C46XAGDRFHS/1NlWaJpPWcrApeIxaSdHsMWTW3m9nAbQF7akOK8H
/DHlVJXkIQEgKnAs2sJeV0105rgWKYgccN7AKf/BGDQRw2XlAjyihSePTm5URY0R
AIrdjiDI1NDEjC2O4/hqxLqrlTx+ecH1RGEjCn0crIEs9CPclwOBRguTc4tIH6cn
dKu0nJPwC6zLhOk/757zBH7muoYuDMzB+qCW/5qoEkDcZODcBSPwgAYLzVJFOrTL
kZtbM2+NyqdEk/2mXrXTN3mlelRGuNYG90MJlSdImb9NCPv7YlBeY4fSF7ylArVb
ZnBxwRF66RJhTU2xh0rK06KXAVqV38LscLQaVvHCpXZSrUzKAkkT8q+jK9CHkGq+
F4jC5eVvzt1tn15lazcNgXwb8wi6V2g0yvpVsbiTs39K5wgzk/7Hj7Vx0qOiEK98
9DnCpkSIdWsZ/xy792jS0fzdP+C2T/6i07OIIwlgwI1B6JkNgBY82uiaqGm8Sr5u
aUoNxTXJdolh0V9swOaY5X3z+6UHuAT4tqB+rvHA4ZSTqHoz2nhjh9ARuRV0BT5R
lwcJMq/VAm2iB0T5Tc/CJ0bN2cvRaBGG9HiuQ9axLWx974ZZaILFvAlOEA5v3FEf
uceHSxat8hSx4JZeBb0hatBTBxA5SFk8e/ugvIhZu1RDLhLDduA2HJC/szLgka7Z
PZ2C5TsWa9hfshaOZs4EFWguaeo+SvyRi/tyA41hjQOcCwi08KafwNFCXKInyNw9
LFVZwUqHPvVEE7qcObCnHmwmASixoX4Ged30vcqHxG9HFPbI8cCTmF0r8A/FvXNP
QNFssnN/kNnBfFD8JtXeiJhit62bC6AFmbaOVKRodLaC6EYQgWLyqWGI0U0Hk5tn
cc0Rf6GqBQZGCP2OEhmppeppjA6yla7Z9PhEa4TcnIVkJ5DftYYe8L9LnfINwg/D
w11N0RwVkgVyCxmEC9J29RnWPX2nxF4VIxXx1F2P6FVsZ+RGhm1nvzIKlIPwi0Rc
B28rInQk2QNUB/5seYiOqKj48YBIxlQb8Q5qnov5dAb8oDCuCDlzEi1T7JATynp6
oTR5/KYHbOcp3J6wMKC8stbXWv2TAp9F6AHC6Wiy+3+CCuKKzYmUn1Y+hM2ZVJOv
UHXN43EJuY2fcMAVn5l8358Zi+vC3hUlc+9/shcAMu5RO8NKEUyOMyxBCCe2kumx
dM5X2w5UbLTz8GF64HkBXppqFQB4p7WXpHrm1kDA1XNb/41Ehigzv88Xu8bJDA2S
/zVUIk+EpAPoSHGwXzfwh0LvcoL/KhHX9WjFjfAsxm2ojqNCwvAScsBHbOtnYWCk
qz1EUXRi9FmY31N4KaYb/GfdBGJjo2m2v1PITQYr4MXQqlQFLj5jT/nGaFSTGT2z
ObFCGt8MVj7jxjDShkHrFfD2C8rnGqObYsxHor5JFgPncqVPVKA6Mfv645CQvhv/
kjez0knWVl0FsPpjy8jbFc9PniUGlnlVw/oqW6O5YYzTTBk88Ej38y/RRiiX67ml
mNemMwUvF3+lQ52Q4Q3lV3hVRqcWFW7rNbKU1GS/h1LBgmUTs1vWozX/N2wJYeoS
wqPkxprgHDVD2sJ4JRC4nbaxJVgs+84Ev4S1QPn5a7mTbNu7O9gF48DhsAym+xog
/V0zuRHovpp+OhF1KbgyYUcTjw1P9vyAic9/0TqEyoPBeNALz5ZkJAF0Y2dyySg2
xF7QCQ1IEEpnR/Gh/ji9i6Ky5s2wQ84yEOYM6K3d79GwUPHwivh/H4WU55wjgvez
XsTzAOw0PjzYIOwE4bReMKSc/K0u3vT8XaYLra+1qKXuQy4jpc1Hh0/AfbT6/hnS
r3DCGJcvyelQh7afoZFR0fpOBgeFheXw9HCVV7dPtGiyvMZB2qnmkGp184ALimfA
eS3y7h+t/7jVEM9vdWuHtZWf7Sri/ogk4xzT85EFsdn+j2nK+RQ2aKof651BdzYk
A1cEQ1zD4G/vNCJB8xwJ9w0qAPy68d88h+ERWeQ01r5T/cf/Nh5ei+ODbnBxPeno
/vXGv/o2rYZR9Q9Ub7e22BNCAOyRHEDed0gYocJamneDXDTRbZ5ngMG55hWSqY9B
U9gC1k4qJmw8fZ0RhLVjPXi2ZRxuWc6rf35QSadX2Q0bxokBWdqjoWUY2MoRZI5M
e6rZ/pDwWS5HyT6ulyQlgEbPS5QXsQwR7qVWbZQEUaww1ESZrJuzD3Ldfn2J3ce4
VysUEnrRWUfgkh8LTG7asmcIrooP0CIQ9TeqIP0UJ/s2gQiJjiEAXA3kRX+4wM8n
vjWw+pqDNaCKTUuR/yzTLNSvxxam4RCbzfCzG6xCi8+lH3nAbc8nELB1AJnanS1o
nSqeE1aYMvGVe/2d6B8AyuW/XPYiGKANWXDM2RZpmOqHrje+X4KdRG/IMxqbJIwj
PZHiUudcbO65R3J2qwD2XJY1Kea4essyHosyHKKvErq6IHpRgjy3KwJ+KfopFlq/
nvEQoakbsCMQf+smwDqj7WcZ/Cf+rn9eRFHf5lC670uASDuEikt/rT2PcD8j7Fe6
i4tDmEF1LhKQp9o6aFWuumQ/ZK5VcCYJOq3wEQFUtZQ1RPrXVpTBKmDInUDzoOQu
BTEGBMUoCYvRHMuCzrOIEAxmTJ431BpjR1K4774JIMjZ1KtGURhKAVR1yL+I2q/w
ANkpGuxL1iufRRxSFIFD9b6oRJCiyyx9OTBnWlRWlXDmrkgGC8qY45eHwUePUNbU
/+CCIzu3/sCvSgQdzVX+cUv2d6g9S9snAm5mi9LoCGH4NowliNI9AOKawmHc+fuF
Oqce3+fmw3yUFUTbbdjFR1tEpp4ZHbHl6KvWzVaN28CQfC343HFAqOJ3/D5y8www
JLiMABnFXY8nZ5ELpKOyitEJYATxzOfBORkpKbPze18dHfGuTthfEPEtG5J4wPIf
iEJKXk1iE43kCz/AL6KSDBWwayGGAocn5fTvo/rJirA8gzIJeIq6Dx2f2N6RuBij
dFtjuqKndMwYDobywPtB0npWYGbN9uTdXtDl1Q7vs7LugckJ30J4TZyuT/PnKbrr
fFts/fD3ULQPzKta/amDZwuaaZhyydfog2hJym5RAejvDZoUeQPl39ZpMigppcBN
HVrwkG2xCtY+SgcY2pKZU+TtKb4UvQa7tYmy25rNizoYS07a3qlK9TLQbehrQV49
vZCqfwYUN4rjLCHXeTMpeZW2sOmYCoumOztcBOtw1FG1YFPV8IxcG971RK/486Ni
SN+ou7v7n5c2XqbctoxH7LdlGbnPPMdYAxu6we21Jhxz4E6DemakCg7A4eaTPw3c
EAytYOemI/UeDYThLlsQCxitLdKTZ6nrZp3hZhGaxb68hwDFpQmoTR+ZNYbj6mGE
72mXcIBlOfUXbM5OpnGvhqiXyP0ptC2+h+2Q0nTSqtJQWHAO7D9CY0AUaKLYINk4
dhPBYM1MEiHAsadydehor6z8pY6F+F0VpB6xpsX6YgWKXhNS0m2eEpT5R5ga8x/e
TdDwMGtSJ5cpDFIb8MQdjagaNjD78u7tAxckw9Kce6QPSpja0GTwNDXvxSjujr4N
l/vcTE0YH45s4WX3fxuIlQTTmVMk6J7Aqzd816A+KQpZWU+4SN3iRKPIy9spb0er
mErSwJh3pERG4FXumT7URxIGuguISjPVoVlF6idr5Y2JuQ1L0qSi0/j/YYS2IvRa
ql7lYIKS9gQAqO19Mtpy56vULzOEHZRmFwxp7MDQdxAGc6NpZqn9mN7xZCNCjq/C
n54Tpr1XBdBxRF/tq5UgJy/dGU2FRxiMeh7Vs2rlujLVEelPubtMxCeNh+/sD2ST
EmpjNXEZqAodyslv9/XEtZyZtJ5rze30Rpv+S0+ariUCh6Jbf7lrl62ecpC/x7Dl
8frAHY1hvbszI43yCvEa0gh+D0DTaks0Jg81mWBGOPQJe3uCL+ONkF0MpOECbM5/
ED1iMQ2DQzyRaGBi2bWeM1Ev/R0TskyisxtEJTVZL4dRABJWIauYHLLx7Fcel9dG
EdZ+q28l3v9yZybPmVclrjnvGm8RVfoX4/EeNMxS+kT2PZRS8SgPwKJeV/GjX61S
T/d76HN5PgeFFipA8AkO9hun4sfBV/Zu7qV97f19/wOjBz7IEjm3Seo0qpb7dZRT
OaWRwB5hezYrb9ZCrX4vcaaxea6US4+/10iCmEj1IwkgXQjBVTfKvEtKgmXjMa5+
MzNZ4S1CHaEBiLNjT9SlBR44gcAtwX1w2NzGjtVH5CN8v5rswAf79sGTYHXiv83G
molGY9S6x0w2g64q9BxSR1yKI3RS+XKJi4YsV0fKivL0LoRMA/ysJ5yl1TgUCRNZ
0WeYc41RsSiuFwxXiIBRZ5O+zDQOUkCNE2ipt5D/d1PqLxg4rose7UpcvM68DL0g
GhDrwSSzyn5l4Cj0Yoes4wzy/mZhTh69k9mwj3S0g+ixbbTo48G6Dav5oBDtoxkA
uQIHeWoAdUF41g8JIcmCLaIocSQAHosJ/74p3iRguM6pu3TlpmN939Pzn/qAPU75
2W78OqcQzwmZfFxJ9oSjq7ux8SYRE47+toY+B0ZiLWi15F3Cgr/JBn+YvKGU5gik
ohbo/U7+/t3bQJr+JeK24KZnsbAil0QaXTEssr2mzBDLhUH5+NspkMZEc5sMABLq
FTDk/vquYqA2wP132/lPC+cy6xtawRme0LiL/Ys+wwVRUI+TKp0SfUO0CkloszHZ
XRQRaOAZafo4Y+mPSL37H3IeLkc1JSUmInaRhxc5OWU/kkOhxATJs+Ty/Zz9WcGK
6N/Zm7lQQ7Btoas/dEdTsgubVIwoD1fltLOv4m53RCq0RkOu9l7wVlF6X0bB7dK2
DZBQzQ62iuNujPGAYt88HKBrt299AiebmctCjVp4BAoh69wbbxI+G/WPn4Tz0qz1
Gd+0P4JPVOf4coeLe2qlt+0DDf0hUJq6KhAIK9yXSNVawctTX056YZn/l6JVDDmu
GpMl7zzyGExy8OPIgvtfPcuHXpEbudI6LV8MrYMwqi4Jy3VqQJ+Tl2EB2eBbrU3i
GDeq0HGhleH4C5V1P59egTAoSslbA621Vo4YWzhryrWWbN2MgcAf3JqZL+T6NALu
mRq9xEyPIj/Jy1RPKhJjcPjzTTxZXOgHXFy5J+9EkujQDkhYX9MLfpNn3V7GkYtM
cVfVXNboKanoO3fgVtmtB6ZoehDjhBXnvngVf2HdrqAGmMy7MUJj4G+dSCKCvUSc
vz5AO318OVpa1G4bcKSWomgemyS58b2Ipmrn7LPuvnKYJPViXBSWSIoXP6rMCTQH
3OTgYG+YROpxx2ZoJx7v313/2n1MXdmbkbAQ9Ig9n2Hgv7ZlcFsUJZJY1NGYdFTB
JLA4xCUCEFwCIp/qwhL5RBqx7Yc9ZS4dow75E53Y0HKuMlD2kfDrhP0LBCoQJZfj
L6BAx1bCYyZWTIAYYa32hLZDI5KxyGzfsk9X6uLuVNHFURUOkz45j7Avq6XjSgxx
eZ7y+i3s/wohsadussBkqupyuNitmgbjwvCCzNfE8NN6R+nBRLHtst30eNkisUPt
YNUOjB63lX3UqK1kgtIf4a0urUEc7vDetKioN1WvYww/wvSe/P7di+Gsm3DbupHZ
vNZH6w9M+Bp3eEB0SZblV6G0eEDfO/M89dxrmIB9ypQJqsbIgZZFfthgpDP+dpiP
nVIbmvIhhd9RdoJvR9yfB1ubkPbeg0DhocVplqJ7QIdPVzLOI7a1fGPMHQdkmZpc
bzdBszC11mx/YbSj5WkiiWobokCjg+QPIEJBti1FCcyFO2UI5u1LwdU7zTSsAIom
LdzPx6nNXDq041saas/FlFwJh4o8Y6OAJdqStYwlvcnaQgGL2gTtgY2DjaD63HhI
6y6glLsFnv4vie5A1wavER0pkp+5tg3fMxoo7VKMJaOVnIrVH0ihA4aYqCIPKUQt
mwqGWpgJnPV82Kk2kMwyygC8zNnbj+2dCJ1SCBSZnGt6fG6idHoRhM+e6+5S8lq0
yylAGVym75al3fqH16f9bZvPhRKRdsnVlJ3a72xaC6fPB/opt3y9jfplOdXJdisZ
dZXbdup7sqqUqLSvTJ9ivRdl4CvObo+JknJmDHiMt1J0BwOdeuEmtdcQJKwyHkxB
F8CA67hSOYviJjB//Otg0uSgPBojD02W3Ht7fev3CijIUQWMc92Go6cLmWo/AJdh
7us13Xe71BJvNCZbuRhapUuLa1/sN4hUWQ7XMkTRTHegXGExSwyBI7u94PbsVV2S
P4vTxpFwaJ3o4vCPwdORAFiABOeOaQNgYdxMvQ9uGv1XXPwx1x9ASReIZhUPPZur
DCcFQfxTu/S162IAkCMwIEuYQyFtssS/Il2ox0ID3i6JCe4IqEUsp+4FsINpPfEu
PZ1b10KA6IAyy1cjwaEFynjfy+sHarVN73VBMP5StK2+568XjhF+AfJ3ePzX5fwX
tv6Fw3i14CN0Pbm4G9lOXGau7cDlHB+nUKN0mgAN1+56ndpOLGIm43gZsbmOGn7v
LmRJV6PH8pXScrK2JxRS8xMmB5fz2orpO90SmhIQ+xe3TrYaLPRdGy0juCXIvhbT
mIsRsWyL/eqRO3HFIF9dfHqSkieRb6anuOoD69nj5ejKnSYNq35H4p+hPeETOaCG
fIBLgVpD3hdWAzqqly53XBqDAc43Cg6bwVgN8xWgO3zG2jMXyeXCodiBjhcAmHnb
OVJtHf5QqtEyMg558oeR5Dq9vFpZt3ifKTHh/Gwts2Itzzl+qHRFRYwjprTiRtEv
N8IxxGpcKCZ008wKnW2AWtNZ9WMBIr9QiV8yg9zjWJSABXYB7EOINtvwY7dVZr58
LY0A7OR3zRjzry55nRBjkLLkNL3wuPegmvBUiTwkcYesI6BHCDEg7WVEAdEsv/Cs
thR2WXjs0FduoUXBgaMb/F0gx92ZbqiEpKCgEHh3zB22DiSZT1xinhnxrJf2HEzY
p/7dlfJZArzaFil/ORTF+mwFSuoLC7HWZHdnEVqgF0BwuNTmwGQq5MgoQTnlGSc9
py9MIqeD28WM3c7M3spMe+JI/Y4KKEClMH6FFHJkIbAcgISstA8rdkcnYWR29zz/
5msPnFJzON4E12nshg80VDTiqgw3Te3lxw6iIhPTEtd3Q4/gfy/AWuNvdFydmKAH
sE2MAHoF0g7tIS0ovt0s4Ngo0lnzja9iUa2PvJKP5kR+M1ws/cUNiofcWXjbh2uV
Pb0ohCNzUyApHrmqmX+ylQCrksUqvOTmbbaQk8PcHm8eVEcHv/6zuQOcv0T+4Weg
3FXEMNWNhU6OL/GF60qeQE6m9KMvlYUN96G/64viMBeG2JuDYdsreMU6QUae3lyz
nMUavfxfCbFOyo+Jd1MUbq2048pAi+FOCTylxQPwmlEC74BiMqLLNvtbh3ChXUkB
nWknfZhl0qsRoSNfYY/nyq5ro7igcdVmEuRZLkBYktnX8MbrK1eTmEaOh3COUgUj
hlEVeTRRHXVGnApgGk+tuYxDL0HpybKNfRC+MJZRDrixi18OBaNtWGWu2XFymcyG
5PI36PlTiywQUVjSdSsif78TNsGaPVbMwrBpvkW2AqXK6l4JM46N1dWExxBhP0v4
2rUbMlEkcQT7dZvEHJJqZXqu3kM9LVSRYyx4uDqRlzVpCunzWC2RNoBdU2BAP3ar
19mygSMK2xnGhOIVsx+B5gagLsBOu2WpwY2KrHpXBi6U6quYmhZE9YeBrfxtgdwv
mlhhXPWAfXZkN+uwxM4WDsv5TlhLji3/6BFjmXGVSKcw8h6DyiJjyYVabtP15u89
J3y2ekKsh9IqXNkfF7LCJL3ls07Dk1mZ+bGVuU7BlP8yLBt2wAc/647NSZ9WCS2O
KDdiCTZ4k2WB/SoI5GA1EgpIuYJYh4gPfwlJ73HuJB+/21MogC+l4tcn72ITQG8+
N6vUhruyO3c28fud0q9ncxRu6ggKdaO16cTay8Ct1J9uO92l+jebifCDJSjemXtx
26KY/1oLE1a/mhz2PKOiOOF7q1HAzGbo5UdYGPF3y9eb/TeVXsXR7PLEPfiUS0hG
4YwydhRq7zASPScA/cNYoTEhERYgOAw6xT4nzL0wfgFpOHuc4j66A0Xbg15dN3gf
zLDcI0+0431gHwVzNCrXuhdCE7R9xk2tW2nwm7i6HfcmFcGdIuk8Uk4ociyPiGuw
gSUzAubit1BJpLPlJSqbXaOwsrfiHgIlxBbArGv/VYKIJ7cyURahkncC4pEpYEla
HoDbYf6FqfDUQ7TDUj5RYBLkc/2yRU0u20fTxsh/UJzWnQBITzCtJczn72iAFl27
PZ/3JQyhHEvLgB2AcQsOxgNkXBVTYmr6+RVsDe5Vz3oaeZH46vAXtzanX0Wchr6C
HnDVEaAfJkzmdwV24DC+6bvSWQd4I0HHbvX+Bk3LPMRDJ9get+3r4q9nz/voLjCa
xli/gyxb2IrShvG8QaaAQLP84EEZnX7Dh77IARrUg8FMk3C+aq7f3cadK6ACgXYy
+bZhJFhIMr/Zufom2qihncHvg10ezvJPLyN+Ch+TMxdh0VBCkkl0kiAXHwCrnHEF
iH10wegOg5uFXDXW+k/BaJSRMjt0LB0AoFTcyKhQ4GTvEWKc5bjA/5C5OyddAdto
yHcH3j5z8YmHmcostalhFxqPlLtPuncO9KmKKG2Lg4y5JPlCXhc7i3Vpe3gSyPFh
pfxG5fk5OZ81sC6vp/h28Mx7quC6UwOYYooL+S7ZxxNCQJBHhTBr+iAWzXWvew0D
dZ+spFSc5dzVobb3EBnphrG+vvnnt0jMIwQ5ixPSBsaHypKJMIzEzlKOr/7MYmGq
qjWVM0mbulsvXj0CYMbb5G27mUIvl7mHeSo9hqrN/SaXB27vHLGwuohma349jI/I
Lbai/Rr7VMq5wKZtZ9WKGzjdPmBWLzVZYPMxTvYrCQiJftp/jkEKEx60znm2W5B0
dUky0Su6UtbOpbGZaytWQkEX/PTxVbaXpfw8IJXFTo9OKpOCFZbAlJxGu2v3Wpln
rAsQKyFd/EhwUP8Uu6ArE8IGFdnxnYXBjwLswgRgvkzzq6PSn/phT8rQUOWbLZo5
vItp7p8wR3K89Wkk4tR+h74ZlnGr4WYMPRZrxUp6BbHKKH5HIAdI7saxiku3ca+/
Vikc3vxuZZsj7lopY3OfQy9KK93CAIRHL0eZmA3Wpowe6tunLLlzllclN+5Wo0wz
+yEre5tijdsq5KgsLddHoS4T2DFyLt6r2Y6ipovrwzVhUlgvVNsuz+b/B5UK6Kv0
TKPLvXW4ckjT455P7qi87KnFRtMa1k5fE0j3xw0hfQCQLQrVrUzTnAktkR0VZPw4
FjDlrKMKAfBvazrJZcy69V9xs5LDWjmeKhJm/AbP+JXDOlBYdQtp5+PHvqQccgBj
d4ana3bfEBwHU8SwOctilLOn8qIHqHtuEDNU7ty6daQztzOMIbFt/1NKtIx1ilYr
n54qX34x2LnmFxNxfRptTyEgtqMH6SlBQjCBlWOmyqktpx3wIqpKBxd4uhpaqpuS
YbezMOGRDHJDmIf1JHijXKghC10+6RamH+IIj6B464jU87T7JI/oztbA9jHKWaQD
ZRHp5475meOSPuoopUvY4h007eROqbLxc3XuPynRwZGaBf7z5bwcuZzbfqPuEk53
uGZwnr824TROOLjILostsX1PupNKXW/MWe4mqLCUDfdQZ4J+WubjeLqPZXWwr6HS
VRE/beBgTZjl/VANQK2z8g7lk3ZFBfpobaJI+QVQcrjYACSEQFzYkymiOmQB5ps7
EP5ajU8hNpiKHwpJMwaJ4xFikKixmf8u3Yg5yoAaEk3zJksZsvuTnPc3JUN52XD8
INo3nm0oIg634LPLW2l9QkkdcCzZJS3vjanNrfBPrWpdIfpKXy09HF6EmQ4rhD0A
KRvfmf49xjByloC3vxpna519f2m8PRVysMctuogrgfzDS+c4NimLUYDE4Q31JnP5
NVjhqJKduaMSQtPIPQnxIMXBmnNWHE1KmXcDpSBQ+sr3MstBV7V9PAqMd3wvI+QW
JwMAyHITFdQobbYvqp12gXqCg9KGx4opd5XJKEdTKY1OTFGQ3/GjbZf4JCaNqwef
akW/baMrdYl9811HmIhnfK9I3HrUw+uJ5WY/To8iOnP/XyR+LcTzpe0s0havbO92
tC8xLt330tQqfoAhRm6y4n4HeI5siTjQIZGgrsKc7gh7B68N/LSTqAC6kA6uhCfu
uHkAxTZ/aJKXXoAlHbks7ygH40vwP4YLM3tNxr4LGAWUbay+O1AD7OiERbezi86y
iyCUnTsdbfMpVBHQZXhB1FZDzi9DfFhOMb2iTAMz+Eve92yHoR/Cdmsnwx119cvT
PfYOb9ThLuH7r7u6po2Dj1hBA0P6rLveOfA4Ge6jsfEBUlYAaTH+XTqLHSD8mW51
RawEPaRD6DL3S9CnSVXi+8LB7crOs1JU8k2Ml7xOO+jtRbkgNcW8hW25g/MYbUml
kcTdziXvU+jDJ8A6C/D9xUyqpLjjpO2ZNRyEKTnRqJozICRbfaTWg6WgBc49u1Fb
fJFI/XwpgCllYze/LOk5aAiaRK2+DCwPBtu++MHEO8XxceaLW11aGNoia0lJXvn3
vojaMRjDKfrG+ZRUDuu41rLeHnXkUutwGJ0FEnS0K0d++9dYQAhQ2n+TGwjvAZer
UqsHTtGBvCLubTPDxIx/r7UR7ViVovyWgCDR6NFYc6GF4agCvWKb1ooWVF81vJUO
QWSeWlNPzV7F9v7wk2M1gvmyos14Rt3AXEMtir8t4zVNiPLB9OwRZthpjWjmPbyf
5rEjfCBPUZ0aSehlG7Dh/Sd0F/ZDA6hT0SGWhxfmPeV39RtP2HFWHrFgWfC+u3n0
E3MGikoivAuTRDmpMkj4+kOUJnrXddCXwSmfdVmMMke3qNM6W5H82UDYqz2HbqO7
riZYPhkj/aiULLrr1nn+GYrLIQeV1Z11VyXO/Ep+w3TuSaV6FmGf6nzIMWk22JXl
gHm8UCD2JcTmMQyb5Ssb87sG4IqDL00M58nevtT+cpYpRQ1qTJSUCCHx0eyJIi7b
j42ZL2CBRK3wlwW6X2ufVg6qQClUR/OcfHwgBitXxrwXwai9+JLlSRc0MXUA9UFY
H7G5Mq4xrB/ctHkdzhlwEitUzweFOEzJDHWKILoCCa9XznHQ7ZmGv/qHHHIUfUXG
g/CANY2BFBhkFN97BL6bGujh5xPRXwFx1in5qXUCAh7bxLw38x+EE0mQtDDyHjM3
IEEYp+iLxtRxrpAe7ISlOht38evBl852LmRlqaWApdhDz/cOUTF4UMeOckEcgmtF
t8chqUz+Dw8iAXOdi1o+0JQfvlQZWDPuYdg2GcKoUgJGsYi7zYuXd02J2fLZrliE
6AAkKeRRmQZ+9srTFefPjD+HFVfdlxbiTQJpMTlFm2nhfCN2y1dnWFW6fVa4+aK8
vnK570M+VGUo6axVLTtXW/Gw1IagYVUHOOR4m4z+odXNxOd3b+a0AQYVzrCKka/L
YGGIhGI3ECXYtSklwGVeKq77rgBjQxyQOKyKeyQydMJCrZXytqadONK7ixWti83L
hEw1+5oiniN2tCmnEHcMFYMfP87hJmqm6VtXeI3Qc6WTR68hdtAZEd/0gdnOt4jL
3HZDvCe0w4zjOXyJOD0E8lV7ICv71CNDIRh1nEzVFCrOFYPyMtYlgGmfKxjlbknr
SGaoXLiTyxsIGAqy9GD++OHTR7zvvMe7Q5wAKTzwCtSdOMSOezGQtFcrbp7+iFdE
0uPzxKKg3OshdsMTYLl9p05oLHmlO5XvrI+b8La+3y7ltK4wWVJlK6KOw6MTPNWI
vwd9mo7tPF1/mOJxN6YsM3HHZ0jJKiUv2mwUS1y+fXyNx96SsqpyWNUFfxMKjJ3Z
O0r/3LHsw11znRRoPdXzWL3iyr4yvndjarQ2Nl/ZcFNNt9uLy+aPbaZflwJR2MeY
A9Up/UcApPxQqYN/W5EvrgOddlk8sn/kShtv7FizCM8oKQNuzt5ty5KoeFmMlvV/
H+fQTbVVukJbr8fY+4QA4eRu6ZGEOZGfJBNJNCS5NJ4tTs0iGSB8CUIlOH6LxQSg
NffXWTNH/PTJsWIJsSpNsgbWNgm8lAyAlOVwdn8xnUfaniUuQhQwm1diV5WjFfjN
bNC/Rgnysq3e+T4UTT7XpBqgXU2G9SJgYupmECERxeMtAiLpON8mf8ajIfS3ZXHk
PIr5ks8j+BMt/0d2W10cViGJ15hDPdFkUR+qY+2w8Vx8UBOaOQUCJq3KLVyX+EDo
7fbnOS4Ki1bve+KyL8AhJMt0HXbto+65AOaYFwEgbqHxxYHMIaOrCpFGbfz98WVQ
iPaJjiRSQbdXTr3qrLU2nO0cHSUI9YGGDZDLvW3Cj/RBwoqOZQRHiQmfjgmDDaY3
IClCXxy2AjWZ0SrgFQFTPPw0kSnJsHK3ZyCjxQrgk5AORsu7jyfAQxFQq5fz6A3p
3Cfa8z7JmNMefiQJUEtFgLQ+zegrIShUb7O2edevEfMk+wQLVJXzIV5pYGPo4udG
E8QvW+5Y3HyLTxX3mXE+dyVp2GuNXxOdoRMQtUv+U3qpmkPpc5olTtXiPuHYxG0k
w1GPpIIjrnvHW1+0E9rlkCSIayQK7SHQlnbVHdncaEuNkcBQ/DBHNHpUN4lJEJLC
B1bcrWnirrbsAm5V8ClXb20qYw6r3IDldRG0yogGP9LHVcgHPvkvUMEgdFoxN8yJ
gUx3VIIxBAq/uruHzKAeWAUl+3Uv/cW1+ygBPVuu+v+3PAC1TMOvKFIIATylYwmZ
u3zNK4ORq6PjKjCJ0IvJTbhot2QQGtfNYIU9D1tmBOzO+abdWum1/ziG5sfj4pwp
ngGNfUvfzxpcCPxYd/rLSr/gcPlzMtcArp7JGyA9RZNktwx7gmQbrkrVourFxOvA
v9Vz06mkEz1VKJr7bjXVfE4Q2P8lzeAjXcrj8MO7MSTlsCd9ZPBh9E6I9IPdvr7r
Knk2+V+0aMNiyeXvx9iO3Qgs9//a9zEixlS/3VmKZ+pDB08c2etxY/oFP8P2yRDE
ZLEAVVRxrfnyTAm7VTJHg8lfNCzBdHOdApSV+VR0CeI9D6ep5kvDCAU65bSDdoyE
Ga9QM8wLckT7DCHZaQ9YE5CpI7wy1QEQfC2LeoP/3pBVcCv8R9JTNBmW/rXnlS4+
M0wOben2+0rlNmH6Bwr8wqW2NpOCpfrZ+VsXigCgo80tDfdYoO8Vw8abeQLsfnPO
8Hquig/HcqH7QgHsW45Y89DDXkkRCXe/kFQyfpcNqHtdbGC5GsQoybkt4J44ZEul
3ENIu8tuw8I6k1G8GdjpmampFuy1ijG8zyCwqpLHAdbL42sr/JhQlYnKnW1OlcB8
3zL+IA+1TbL9bKyBMTtep5l45hKoCakLquYFAQxDsOhYsCyTcUOwta+gCsP8ZcmP
7rB+C3cLzUQvp9HFDr/cOWItNZhl0vz0snfMhgI5e/zNNwe0fAHZ7izAP5YRcQRB
p2uaLUtEHohOrhK9FVTiue/sSFSP+EsrR5uBjhrSrNiaurNCVF2jE4Kof+scQk+c
E4LuUdNlHl5SqjMbdpMrAve8tm9wXRJp0vBFMqNbo+HjKXhWrPGa+6eyfbmOj3Iu
F06pO/2xBAu0HshEncYrVWYR5nRUWmDZ2vBvukyeVNmOr7OOeNs8MGXPtJCJGwp4
WkirFIow4WGDKYeU4k7RPtLtqg/BOslLOXh691yHeeoBjBxhgy07/qTeTKgVYr+c
/AbU7nespr0w7gT9WHFsXld3xhx1WBiB0MGRd5aPMCjmPIvnUzxdnB8EAX37yuzl
ipdDctN8YkKnXYA+fJgW+FtC0kamHqarf392fNN64/xcrYUl+VuealRrgk13Ha5L
OCb6FKScPoSsMNewJXJx8heMRxENvB1c9NAUUDXJ1NRGe+DgmsiIKeSnLwjQwUQ/
9PSkinhm9q0JtX6oUIzUlUu5K1nJr9FUVpCMADJRom17H5FBnkjTqtGae8edXdVV
RK5C383WMNVpbuYsg0bcwm2RQVvtv7PVrjhRCgtiJ2JYg45Rex6qSjE01Ifjbr+F
7OR47r56yc9LTGmQYpeSh2CbhqYMn/s8sCPvFOSnI9VzOPmqLnyw4Sb5PnBbD40Q
JzqCswSV76v2G0I7sRWZLCXHEZS1Mh7CIfqjmTYvObSBGazsIP0qCsXcRrlJTh/N
WWGUU2/u2sKI4aMRjoMZCpXdnz1vmGgrsfPZuB5sAL3fjbuoihGUnlQCuJBOAUrp
tIeGet8tphONkLealp9ftz51POyGdxm8YoZdf2deWpz6l+JWIQZOaQF04sPIbUMh
1WFNEic+asYArAr4rhAHc72ZQNGPSAjqHI+zMCqP61tdhxJvsX2yISTZPW9DLk4A
sKb2YK+AY3NQbg0LptmIaXotPuND8OlCLI07JkVf6jeOFq8vsQqULcFv7qy1Uion
E6aMA1kPfQ6O7hW0XBBZ8ZdCHsINHrC2sZIkyrFa8C9b/WSWZCTFswSEe8BBWjoK
eolvjmwTntNOU7N/X+XZpiX8zUGKuuSVWM0Ky+VD0+l4aEP5UX0ZEZvKOD/zFswi
OGLQQzco/Vn1DjiE0gJu6XXlqGVSe+n3qG6GKKlyvW8lDHuxBBTD59tKZJT2T3dy
vplP8El4gGTqVy9cIUDSatMLiAWWIPNog/4E/MD1z2V/+/0upQe05EySDxOR+HSd
sjdPpUud5xeG3KfogIyLR6go6MYz6yt//Zy29ejKgXBCH9fPJ+CG8q5Bf1XSop4H
sSHlcY4Zph4jW1yrGH34CT2+QHJGY/EIWGqwXik1p9G7QVpUF61o2UknqOOA//rp
WD9nZOuIOlMZ3oOBsCGs5pbnQoDDcUAL6C1bviwamj8Ft/dPOh2uKdKAtUzdl3HP
JjE9QkvlHDwixrPMI1WQiyfdWRy/XI5ZsO+IpWd7z39ihh8TdB6Wgsowedp/indy
gZgpgyupD87u5el/4k+qbwX8SdE6uc/iasrUKWYjWNLKsqmRmEwePyxCgoWw8Nou
3I07mNymyfx91UIZvMG64cfsclrV9K0EWW2k/IHX/IVutsND7x80gC9LvKZCKCfb
6m8gkEVtSc5k4cesFzU5NgJOhEAvthLZvSZ0jFTVQPTWN+5dXa26tXLHN5o11ii6
8uWM+MGGDtWGibBmNiNvYJM1H+y+iLyQaNgQo5halQMP6dINc06lo+RQtCNw632l
vdxlRW38Q8bCmVUo7CL7cJwFQyfDit6b0eRxueYMFzNIeKgiXkzGgcCyj7EPfkGy
GjsYxP3CGRG1k27+7p/9f4px3V0kgscvgjMV3LgL+rZgC06eANBVbH4CUzKQGpID
hE/tQYzEtwTTGlti7ZfBaJ6lgH0LvIKLKmoEx/hmOZ/pu3oLAD2xKaZmTZc1zL8N
op71sgTR90Ze+8Z0mXjokN3Po0pISh/p1WbIsjvVQrUbEOgATek7ELM6luTKGDyg
weFdKGiBJ3UekEpy6qo3YI3yHwC2Vf6+qxr0o9in2ocorcNi83F83LB8zmm1bgjw
iXz8UyZyvN+Q4DWtV9oQLfmEIWJ94v4YScQdsgpwFbFtkAZEzTk3i8/Qx3R4FgQr
643qhxLEAStQcGrs5qGaDZFN8+RXEn+9sZ7HSja737X4tfp1DJK8QekYJFebF52T
BqBlAVUEdQeycWkn4NxiITq2/bPAV+7V4MtkjDWCCW8mwQzu5E3eCWVt6rX+Mg+c
0tN8uEBXMzEhAKJzp55WWO6lqQMvH4pEqH2g94zpe8y8SB/cy+lQVCrlnOn3llS3
LbcB4CTJWRbu2MQxajKNogfgwy/1m7Cjir1KYJwCBiw9l9cu/vMwqBZ23wiW0Gwk
WKpQQFSlTLs8MxuJVzyVDcDp0n/uzGFJJrfj3vSiUvXIAcKKuvbf0+d+LIQv++qF
07IsJqv5FtiRRqfVddmUXrOGVzCg1NJIqD2EzOuRowk1/xIJTJAXATXHXXfImx7Z
TzVi6888MGm6a6/zacI93lhsQs+4RFitk3TDtQek/yWLv7fLqnMbYcHg2xO5nWBk
4p+Sk1GSVV0ct3Uy3Y1xkulun4JqcGXxk3IhlDAF3quVhMDk9mSK2r4I2mYPkfLV
FA+SLYLNJvaf0SqqLiNUTtTRf360oW6zYKTfIpypkqeQV0fkyq3ISCDTm7nCnxwr
bjqGU9Zo/JSEi4VVebsCPRJfdv/5rkRrfKzyfVJEkBt1W74jZR/s7heVL6m6aAF+
dAhkDei4YdG1rNrifLrC9L98R3jjG5leqji+EovPfjOLEkPcpKQ0qyr8eO6A7zh9
vCwe/bqNlqTeaGIid3o/NpnOo1Dq0gLM2CNp+3PJoAL7vrEpFgtpjN29zMXInqJm
IWnj3AT5oNdhtAze1HOVcUlTBP7QTCE6MwdGr1Z3JevgCPb+JJKhk19La/OtP4Gi
wimRR9jFYa1Qyrb/JlL3VL0YEax7LWms7QQ/Dbk3jtlp9mX9Vo7gsIVxp4UCKsRX
1pPe/DCUp/HOwq9Rjda2ZwtqaK5aWKuQDFTHius3eWPTrw+tuwJg/km+bu3RUhtr
7HEJXfky7mwM6ogC1Wbd1ZCqm2bnbuDBRKKMmNb41B+5XtCzym/xF277wXIykSFc
yS2j6otPAhUvAEXXecD7M27qqStaQoC8gyu6yrq0lnyQUJ7FxZ87fbsj2cXZs35Y
OZa5gvtj4YfwPMQm/va3N9x/QR56cV/UAlij80ZmAK/63x++aMQ/tvfSZOyOtgp2
jd9qNzbzhhH1EFEEFphmQlpBHM5E28IRNW8lAOlNWhWEpiDt7jGBXVoXg0nT1TW5
Jc5XkLwDFYKBP9SplQUvVcfIBksMvCBwgFs9TY8+n16HmcPx36BHK7q7EUkBhkbm
/oPEXuNaPy5FJ209WX3RPqg2hggE0D7DVNA6kO/lQY0U2hQoRYX2P2R/25aDEg3a
O9Z/oSqcmoMV4kXOkpeYgK7LIACyK5afAMdf3THEdKu7kz96sGFnZ0n+fnQbjSxE
M8g6Fc/Hq/QmugK7lihTg9CBNmnYJr1J0aKkRnVd8FPPh4b9rdUCd29B2vpP7znL
KU4yGyLUDVEDJm+6QiWjjrQKAeWQNoiTFFz6JUtZfgxmMEkADDjfOspBVSjwwfJU
qoGcWI553gpdemJUamtFvXmG7r7wAbm5cWWEeDaHBRYqM8X3gEnU15wFDkncpvLN
5/7Zi2HY1Nk+iyUiI1mk/zAiz6VCqSuJiHEvvdMF/ZiCIxb1ju8wOwlDN2sPe5ob
LYafccnYY7+GYXFWIFFbGOjUmngpnULlXtRGdWhpf+/dBaxUfJbkv8JpJjKoPwp3
pxIlFL/6f6JJkklFTPucXWpuOJuXEobUMhxQ0+/g9biY4FH/5fe0OSWPJ9bgCFOg
ELUXfO6bVZpOIXEY7Wb5PHoapD8HcAzdOn0k4eZFH69mPBn1186YhUoiQAk3ht2W
3XqvVvmCiDZrUqwZMx/aOUK26cQKA7pN+3Hl7jwkFRrStHjKFw1CdYHkelk7b5E8
a6wcN6IHFAZmz73UC6612mznVTsmSULhveGVp81Gh5Ueg8J92wKkiQJwPNOrbJPb
gErveRQ13ohmOsxiPqQSMVTLY/UF98B6Xj6RAJLF4PV1Q+6fTlPou/jpk8pYmzHJ
+33Emk3Pd2klBXSSNMINwgkHrrlNWpB/7OkX4FNswHr7fIud8dp3eJdDZplAxw+d
e2/U+Dt/XowOh17d7k7yli3PPLcRBY8EY7VEflutVCQNPzRQ3njTnQFPhekz+18g
OjqaUt/meqYLurs7Y+G9BFNTWpRdsftk6WvoKBmlFZBqn/e/oHCYzRePO+dqB+tk
yOOjDdgwy4pMVImrUL72e95CB5ULjtfjmIFwgGWW8V9Ofkt9C3p10ki6BG0GBtfy
Obl0/Hx0wKFGnBeZiy90yDInnjwMj4NUCcyAin200e3TYnzAw+iNW/oRMKYz7GRw
ksgbQ15qNPMIwWQDmXml9rLIHYKardnGsruceO+4VDYd/sLG/pQfjdVW6WcQY2yF
pyrZaQG+sAcNFC+1IGALKgzktlaHVUFb1iV6XyzYCPgV24k7IEQnrZqgiyVolwS1
TppoScVDhJqZRrDcFTuKo4EfEIdXFWG1JrYXp1gVrqiODxV7mpfCGoV9oAX88nhE
soVDkypKrfcobsDPS5qHwAVP1LGDYLuf8kj90j+jAuEfDLC5ILAikJJLE2VqCyEB
b35RdL9deb61alnx5ietUNlrDCDhTdBuXgvhVUhqAnvzDJNNSENm7nCud5WzXJu/
fmwlxdZ4POGCiC4ma3Fz1iedhfuFcZj84f2RWky4/fhc7RRKYwcKYMPME2LWwKeT
D8Jy4vgckp3J6qlhTL2lcLEdOHtFOjNVSKnGw2fAyE+S0fsmoMOGrNV1kQ09Gh7w
EM30eoSlZ5Ahi/+4iDRhq46bMhe1YqUgQ2fGnA6eQOqGE8yeZTPfKHwQwbktzSS0
oI4SSob6ih1YzSBKWRSw1PuL/cBu5OLCslpRdDWKJQd+5hlIuIkUp1ZxyiDDNhSq
rPo1KywGMInXBTdgLnMIktk+VxJN9nann87YY6fZSLvp/BLpUJ6l3/EaVMDf7yvM
Wno6C/EbzadLGoRuSLzRry3NbL7kZNnRSztmPsCHkK91pACip0kcggBdlRuAGsuJ
bw85wI7LO/k23UIt5g85NQaYICfE8l3uG9zFb0NvRhr1l0eY+A9vzRAYRrJ6YjwA
aSINGHkaKKBt64l30GwYCOEfwVClEFepZvOsn8PmkIAg5sJkqgg1peAGrHTBU8z7
e67yXe//E+JQO25Z7dRwGVvxswk0lPEoZYB7YFgLfGw5Y7GzeNvxhNbP/Fai7fkG
/Nw1k88D6YEerCbLmjQrTa7UINhS7UapYRxqmddL7fNSewLLDco/x7FqhMC3cDZ3
+76oy8IVSH1fegcnaeEprjaD1yBVorg6zE8be9/OrBP2p9LSbEwPrKRlth4f61VT
5w7JbWLYvH5AHlVVKW5zoCe4encTDUQMmarAysldM6X3oba+cngjLNzyJxxackBI
GzlNiotac5YjtTa6L3mFqxt2s/hxloicwWm/th44n+eh7iFiQzrm6/JKBkQaVZa2
u1UOGP72rWjRtzeKdgXSQiek5sHsyUxet3nwBKeC9D0dCmgxEy15tJy9VfNjBDwc
1ulchErSOCutnNDtwq3tPaCZln+TWlBOTYTKwThcwQdqmef98WcRR4llvU9tSLWp
UyblE8ZRCPPmvMGIhCdUVKGLydgz64iI6HG43mMu+PE/miKRn812H+XP+Ourmsgi
R9t+JIZ5pAN0Sx78wcMauxiVHTBYZfKXkLf+ySC1hOFl2g58lZiEGUcnxOwv4NcC
dG629IilSFAdlpMkxaZdEGI3bN0lwRhTV6WKQSsrlMnSrpyu8BVP+6qEOiSy6F9I
TzOoA37s/0ELO2LRtSzpiZV10vBah9vmd4I7m3MvuBzrji4/CrYdVqUMqAJuxNvS
Dlm03CNBaLjp1YhhzwV/E/y2r12W7MpeRr4C0l7hx1nPXUbQoJ6ld57ljeu+W3Cl
jrh5LC1u0l8+4mgoqUFg3O9mPC9EBybOdnFacL5gHtmilBHsxJpaxjgM20Gxa/bt
8H9D1BbGlGX3K6CJnNBSYxfzQKV0GlDTHEAwWtV5jv4+dvHmV/kC0BAMDXgEU95H
+aSpUCROpgstT4F9peXFLz80b7y0MUV8gM1dXj4KldBzlaEI8JBM4K7g/6yHdQ/s
PrTPMuw+iCPq4wUN8ZZzT5qqkXjmSUBFHF2JtlADi2KkbLzzuHPHyzKTRxsXL7SX
7/2PXb2Q0qFTGMFOCYC3WiOJjeoN6pREaupKzPAK15Dea2ElKas9M0sVx3t48hTg
tkmskd6s2K+KG0OXp0aku7G0aPaAK32TNfi1BeDBsa7/yqj/gsXg2d8+1q4LK0J7
rcz+XP+fcxN5qSXHCV+03tfizaqnJqM9kf/PjFxglXo8h+UyTTA01rbWW8nrMdO5
hZLs/lIa11SHniStz2EocEi0kI+RhSR47ui0a/ngQcT20ft197Cc/fCuGh+UpVmk
HLHojV9MlJmrsBFyzkqIyExMLyyLry/Ua8OdFGkgC0LCxmqEBOMWcoUuziuar2Ed
H0Iy7XvEej203BF+S4f0l9E8cu41YEwTPrB7YK6K92R+F8yuKIa9fFgDfo4TAXfG
x09T/4D0aZtrSsnaAxB+nOOBDJyKPOUmqzvwkZLPT/BhfzDLgrSw+gPG4yc5sTkb
cJVpdE5fRvnHssOufRyFloDAynHi62nlJndEHP891Dr1p8ccIsPLKUa32pkuLYaF
0eUhFHV6bnNzGm7aqU8fqLTCiWl53hsLL/rBr7aVyULk7WnSTxc+ig9uZKKUW4zO
yDBLI4o/k+IzBDBQYwPWpX6rZoEET8uacsWUz+jbg49iNfdMJz+a99zP7fJogEgS
1EfuVOV6Z6gw1vNtD/J4nBNKGSazPlmoVBafPULnlanK1n55VIMsAWqiHf/VM9Js
wq47qUJK7vJrqxiN1ztwyJwBNOpZjI6hhYRdWQKnFoUo7Z75SSnnZ3evwjwSoLaP
lv3uvt3DCJfhPId6Tt1bgEfQc9Ojz1KzWKKAUFMY7mpuHpWJb3DOnIMX5WEsxEC1
W3kIFqTPt1ogopqEOVT3uLSlXAk1xb1hKu9B5NfrOxVjn0uUjLePjCQXXTfMfwJF
KYqFTttBHtf/zrgnF9aaGDvN7SUQpjrM3oSVkLMmntyUfIhfwCc0JY+SWp7xtdVq
pxWAVoqbslBPsZEd/3AzFaoTC4YKKeo6F3TwuH/PuE3oMff2ImYN1DTW9PEMVFlK
3T6+81f7SJdIDXcLUKUnbTSzJakQWUGg5WjAL1qM7XV5jcSCwgCh1iNoEySfuTFI
+eR7sGe+qgPfhApokY0AWrgm3T31c8sxDDtajkIjqMtRgg55jzzzuH75VNZMBr4t
jMAdjzGlE4qtyTy6GS74F2ceSRYdbwtqTj8XeWV3nOg+WoPlJEQc3BAh5Z6PHUx5
B3KhWsR+bLjeTiMpmS2DA4Nw9nhFJRt1hfaqCU1cm/GIHGBcxPLWhvs7fI4BIPGN
eb6q4tb8vHH1nOVqEfWJggu9ub70K9MBUT/EuwwzIMT3ERwkN69i3CNawMkARvUM
HfPU+HVN4iLNlstLzN884i9Y2l95BjKPkOxVAz2z4k7FsmSnH7oPrQLhpzG2Cse+
zQYzm9PvEgQOcpDvL63a3Mi/4gtg9eT4XMEo7R+KZ5Pr5BoTiuvjIT8hIl+n7Joz
zMzZA8HgCwYjSWEI09CY+iHfyfLkAQl/TZ877AvQKiYpEZZMAX3NHqUwgzWDu0OK
GNR5XhvpS5R2x++E+EZHKgCq9bjDSVitymfudgX5xF6EunZFbLTKRUbY10+FJgvY
23NU2NjqHt00gV8NpKAyxw1a5O2Mv2xqzfHO3QGF2o/x/L22qwyA61zYlA3AM+2P
uvVV13blQskO6P7IDc5PvTGGPepXCy0l96o0NpBs50iyS+NZ8spflItyxeOYtB0Q
DquA6N70iGQ0flkcHo/pFavw/bjusnQLuigPJs5TAUqJ4VYjzNNqGfYMFaSPdruq
Gt0+VOWMvVNIhHIyCk2vB9+N3qG+0xGJ5fJ4zwaVtBlvAvtMP7lYgElriwU+3J75
qL1GxIdkWfG/LZgDLFJ++oEW6YungmCKG98wSkTevdYlCLboKdEN6hy8e4EAs3Jg
+NYQPfi6iO5cY7GRKXG6Zc9NBbpHSzwtYUhy4sIdmIuvlUMOis1v8dxZdNW6+1Pc
GvJGfS4SsShljiHNaKjQeLURVmoTjlupFnk0OBK3Qqcr3XYWj/CCuroiPNqWZzDl
egsZj9XBEMRhMNCieDBG5FEUvWp3MIIyNg6T2VirSMjidBV+RMudTZyG6eny452z
XYIDWuvhbjAcbPKUze7VJi8u24M/FoMttWBMjax8fCLkSPk77A3bL7PwxppdkM9q
2gEy8KzhkEHPMkEJtsAlTiG9dUzQeOi50XyampUCaIEoZo7TFmmNWMDT55eHYXdi
Fr4qzFdvJAfdO9q+AwiANku8oDLPaAVZ2JdKFLiA92REtHRFNRYffrjV48OOuw/t
N3W7tUdRxStVPwtO9AW62oSm1PYlj0IDR6htMhyoRHPnbt7wdL1LIBPO4ZF+mAXo
6h3zV+znlHQ4ybw1Y6O9CWGNQmJNrpwgE7xRaMCpaMsfx5MsgpGBAmWQhi0nZCg9
JRzXNta1KGllAjmBRRDCViuZ27qMOk9EsqBwKuQSHgh5bn2Es+l/vdL1VFGyJpXM
8VQe00E6Nz4rFcFQX73kDNdkz0L/0qhZ6u9y8oDKw53i2h4UW11E/mT1sQ9OZAgm
XtxDzt8paVDUmMcYR25vIvoE+zjvJALPLqbf1/oTQUYdJskcMZdkUIZWLXnbUmix
ENqdmXgjnp4R2YbibfbEo7GRKKrOp/J+g+9PccpppCsWT57fOCLVCHg/dsHGxEGq
23joxJZepdcbg+OOtQCk3HW+eva6oKrQYlzJAe2gr2cxBDNMyXrJxAHEKczZuoK8
bybQz42J0nTVdFYc4WMu+uD7ZOEgnWmdzZL/AJw4Xe2TST/35FoaV93EBxPrnC74
1CGAU5whzD5tm2XMMS/0CHm7r6pMBOBo2xEGwvN1yOk+znhuk1wemkPZCZ1QCCPC
gIQOWuPiZO6kvu32+gkVQsqU1sXL+vaxgydQheTLE+234mnJdriqyB23roPZJCyj
bTlx/XSyH/E3MDo72FpFxKMJAilTDjul9iVcZOTw3KdJyqnqRVowZR5V/8J+d4Mk
uDvuOi4hvOPv5K54mlRQi/u5IRqHwypFjfl8sJi2lrKa51MWohlzOpaTSdLTUl+J
oG3nqsovJKWNIDDDjmLTJZSlr3Y3AGr1pos+5N/TjbjOBv0ZbPWMswdXaa6a84Fu
iczmKmZDD6BbQ4F+B1obEcfFECt3uXoEtagH1xHhZIwVXfP2dUzP7ePjjgxmkS54
L8wOyhuKjllt0T0OQAIj78waaDAOZRIgyMtAwwUknzUcX2D/fa02xyHikHwcwUAW
o+tgqViEpDserHSvNg5gogIlQr/eJOh0irJuCWFceYPKbuWM2G19igjTTQeY3Beg
uXoVv0Kec1nR6VqfDDFXILBNT8SnUOdvxS9s8OJ8cwW/9HfI5PErYP0RKNe6qlgc
y9s7jMbloJZNP1zoo8b7gldlcQI6MPSR69MPqlp8dML1aKbYfr0HiGTG5MASgfW8
JkCokqy5BSnYMAVu3dS5dZttuegGiCgM1dOGY7mt5W7861PQQP4py+fcTKALU6dF
tS/JZwRIyDIad6+CLAHBJgjyPx8R/Z2pFqnpdV2/uKZJ3PyujjogEO3akYCdanO1
rHt9gwoLO8TgCqM/HQaFhRs9Geu+pdiMCczarPu+GvWGVzam9kRiRFzrIzR5ocC7
xq9vd2jc4yM2PMlX6B9bPRyJiFWmF2DuaZaROxso4gZ+E2eTpMDxC4VZkuB8dM0n
Pm/P+/q7b3e/VcvLdIJsuaXmWi6cwetaghx/Cvs3Zjr4Pnqfnw8AKwTe+z3N9g6N
u1iRetkuqum1fkQBgkYqIG9FWj3BK2reqOQFMMSYoZbB+KSFK5v+DupjzJ8qBmFh
xnNT34OqfbYHf/Sos8L6l4bLEOEgWwJdixdJxkxHyxdRZdymt5HqY2jBJQhlRgVq
mOXKyRrZu2/RH7VTNxQLa7RzbtFjORNfWER1eNJBxg59EPtEOoNL4Jq68yO70XwH
+YzTTsa5VFY3d1tviqF3ErTnTFYNQVhaHAmqctGDLTz+DhGdwjLvfsQgcT5ui2zX
1SjOiozs+fjyxWPFIy5FEQ51bGGSvfmATghacttVvi9no03mC47BEsAQJlXzHuvp
Gjo7I1P9Gjgbc8h4w1IG3SVzfxLYEp8zc3Gbkk6Xgy0u/PmCgFYum40zGCkQf39L
AmZkl3iQwxzdBCyp/7ROONM1TFq7zclL9EpV2RdXrQGzttUO0mGDTyE7mg1BFUkp
SB6e8tRLI04BhD6mJEuk7JeT39uewJJi72pRtQfD0iAifm5+OsDtTXJJ/mQ2OLAh
IqVwdosFbjeEazGlOTBqFR3cpSi3HOSQGLUHzFel0APb41W5mR/1SoQ3iXW/e7jW
SKzbFMz3GZN/XHjLykACdaKyWOYeJQpOwP0SkXBgCjJRx6Dn1ZDxerrT0c/8Nd+/
jC/+DluWDUZfEwhleZeD9k+luZQadtAmaBgcshwJ97BsQi2keYzBXjR1qGJ1ReGV
RBRuzYof2TMo7HjwXUnSU+XHeFQe8lJXEF6xOOidH9W97gqXy9aH5EKgA2UHJguh
UvTUlRECLs8AgHEdRhXRFqajU/jzJ5OyX0jhaW2ZTeRWZRaM1qeDMVI258XdXBrw
SST0rH0FOldfMCiMiEj6knQTVJyU0vZR+JBHi+kgy2wbVrKvC3fDvlLa3QgyPDYp
HHg0y/CieDmGMGAzfKhUpfgO0oHfJlfREHI026jiOq0DLj51gQL7ramfTDziFN2s
0K+4YBRyuxCVudg8lLXKxsIKqY665ZOkVQJC0VYmH3eMOlKuLFjW5lB9bTC7HMNj
7vDJzGU02JNaaDPMAmdXBCtMeP9BPSROz6KeQaUnN/F4pl1YZ9IpRlL9+zRf+Kqk
DPJAQTwuYQwgITW5jJLju2ByUGWeDps+E31LjF8ZrqVRaxvJY3/5TSaKHAYzmm69
Q+6mqQMMoxcD9zejKLyXRuNzrG6VnpJO2h0yOs5Eq1hN0hM05IFO9GEa2rXT59Gr
UPzOyH/x7hc9+7mvl+tJq0fdmWoR8QQ5ZyejDrMj1OFwvArlf4uLMtMf3lDalVST
v9LXzXDI5nJoejErtH9lc1yb1GgBwZoJdIxPZAmKXoxvmYwg5rFceHizGyQcT0C/
LnOW5P6X1X94FJthPhxGfanMXKMIlgVrNnfCNeJuGmkTJEbRLJl8z+pApiZkV89F
XVpMj3vai3fVrhaHu6psev7WzY+dcQJAUGMCIXmy8yBPDmOlWBsJBoPfacG4t6sy
8MxgvADQrDIp0s9gZheqvmNxTUoPGj1zxjh8KMxRMdj5tySe0QZEzS/fN+Ztzd+4
PmEQJoAYdHAJV75Pkn5NxReJeUrhDZ7rNBCcoU1KDr8gQna5OC+8kUWhtt9MHygh
PUJqd6O4mpGftj6mlfv4psqqhgOo//0EBUyukEa2RvfINfMvEv0yGoI4IDvbcB4n
/RzSE2A1mndozm2ur/Og7kWm/zyZ5kmZ6AVDghWm3cAlU2s3sd+Os2BpRgB0WgbI
SELyKONh5EdlrROBG0DgNIx4CSj9xQQhujj3Cn8m/Hf1/1mHwTbv82ka0mXll3Zz
/89wucTqKDcuNNnm0gWVgtKn6g7WA1XoW6wJ3V4JZV/gPuYL6SVvigYa89BiFgpk
jL0MhTXXBBB13HUoXSIIn9ubwD9EYhP/uvoodPMHYAZMj1qQauO7i/KMitnaBXpZ
i0U0WouMaODwSuxhVbXuLWsWCYiKjyK8GRzfdvP7eORY1jmwScaHxgl3QjdSfW0x
mmZOrdpChNSE2U2hE7bCuRHu/dNPA8ksVFkNZ/lSHoKHhoQ6L4g7zg59h9wQ4BVW
h4pIddsernv8Q8mg58lDO9l/wUlvuH/JS4J4Ah3mR9GcTad3cM5fasMd3QZm+97b
kgXHh4Cs2kktuL8y5V6NXvg3g0cp6kWOzo9AmOhJ/vAKJjCC99wn5g611D3+cRct
xmHrS1X/4nCpOS7OKRU/ue7dgbzchBdgy78JNoK2DG0+ax9WaL0rgJchhfrWSwIP
wB9i5c+eui3/Ae1X/YeD8Rc2ouEn4RmH9MvAr5192h3D7AySjvdNtevlyygvVGfB
Aoy+GAhWXWjemEII+cTcqdFeBshb6ClfBwM2yRMARKK5mpHjJLdHrDJgZK6AriRb
2PYfmM0DTnfKJCiIzhdcrRHXiMhYQ3IttJobso0ya+HsPgijAUwb3E9IC+iVb4GV
7MUCA7RjfYEW8jt3tDJmRhnhCxHJvwqk4QkupGzaWFAb3shRXWIfl6wh/WGebqLr
k0/IUHZaPXPkW9eI7c9ZR2qP9Q9PKlIOAg6Wi8/rXfXNuEvi2hb5XZLspPgppEgr
kzsWAc+YMH7imlOdbRjTLa7e+2GeYH44HMRgGNqLvR1UGwC5jeEGgTnuejsL2fnA
EzayFMGCKPSW2VhyJ9mUMQlAXhP7Ch0Z6xbZ6J//M0VcxzwM2B8fEV9uVCbYq9s9
owTpuIaLp1IP4yitmU4cfVg9BGgT6aS+qGnP5U8VuWk6H7nxThNg4tZbySgVCTH4
qO6fjgxfWjHyDkDkxUWeX7lAO1YF1/zevHsfKsFXU3F4FWEs45a0lN7Ole/b9muc
wL1oiaY1yQ+TMBLE4bHrHemzP7n+xZO+WRbCWI7Lbas3h8pWJ6ZU9G9IrnBq6lO2
OuG3fKgCdmXmQqPwmbVUAi5Ez44DwYa6kOLX0EQ580a/lSmgvmljqjRToEQQcFvD
Yr87p3wDPoN1c+H4feuCvcqKa4fcLa1kj1NycfJxsee11D3BP9131rAco/yIPbCM
rB+QQ2Zb/M+sBlI5rVbb7PDdbdD4f9U7Bjg/3qVuGMm3+NcccpM8+9WmxyvGhSyU
9cQy0ZX2i/A1ozqo/rwoH9IdfwF2twS9z5xmjh+ataF2dg972ut2scpWanhJzx3f
EVfPNPNbztv6wwJDhWrmynpF9xx5Kz8I6hvHC8SBLlwxX0giboBn6nI8UQsgGNVp
DDksM099Rx8KAx8zysiPbV6bz1S03xsXXupt/zNO7fJxxcnUGK1Ls3vUfWoz9kwx
3a1ogYNjW1Xf9CUalyhqG1czgwR+CZl8xrDpjwgeb5o6jnc9R8jJJj5J2NB/DL3x
6W1fYMe0ig4YhQp7gxjrf8S2LHxD0bc9sG3ORAgwCZoqEqmtr8ELcx/qER8zmkeB
v0ECX7RnLlB1sUo6mpdCrwA4LdWnD+JjsazcXBd5bMey7XHeS/DWj+cXgPoyuw5X
07ADatYZn5NuuP/msJ9gdtZmx7NhpphpcVkyUpI0mo6o75D7RJVTTztLUpEhKDii
Hp0CpnZ0z/OUAlipoDuSUjFw906GgI6mGBjyoPbZ4u2lwMcGPRtWlrMYfnZ0CUub
AXG7eNtturWMe7/ao8lz+eKs6BEcYxh2d2taZ9KuveNOQ+yxNzoWRHv07h+BjMGB
ScBrK7ZQCvqYNmMgmlsnZ0ecll/6KTh/TtxcbRQMAmVNefbewlk2PJrBSe0mVZIF
BREb8Jte+ro4czj6+0PzY8IZ5vJ6dv0AxmgAo30PH2tok//G4Cb9PprZuSOrpFBx
kkb00pzjwflrkK66J4i6NuwY8IT0yaXKK0vf0f5qoDRlFuWj64495Z1cNKnjM8qK
cf4MY8j4d8OrgHZtWDYjNikesXdPM4axN2aNKF3Ib1ST4G3pxpcUOVu56sNLf2PB
IFpYJNuNp6xa7yRVxqcRE2nlmOXaAVFkwTI1o5phIlCQADbXtve/RxFW5EQvOYaZ
vH4nRBsSF4Uot37hvIOTPE08tf7qUrYtwgfGvf/hfea7RD/IW7qHfUqn1/qL48yX
LrjxrycAfiv48QKSOAaQYt8qKZpOCKH3v+QO/4Apay5Qr5BsTb842GE3iLfj6Gie
vx7vkszWNUuEicvX/RUr38JGxK3l8bIxmL73ipI6vpon3DoRDTFmCVpTopuEUAQ4
pUWlZCeIpDBarQzX8EVvpKD0A1D+J10J8jASslPmTfxtxEfvyZE/CczTyEAYmYjb
C8KpM4kxrXRt3vp8c5SpPZalPga+RNxnSRNIZwJBQ7oSPLUA6qwDb0aoUBXpHqdS
BDmoTAC4hMBXlenpLDKQkPQ94HgeGf6t9m/FL1x6wCyw/OwGC90e44NX5WawtAIS
lUSuVpKob0JZWK7jMuPBBKdpInHjS2gGjhsdb+w/gkR8GjLyp8e4wUEqCDe8S+hz
+VXTRqpd4L8b/Cf8PzVx4tc5s77f5lcq9rMo01V6xiBy1R8I2wrDdphh/lgjIFn9
77GhJiMBAvh40yAq14nBdnFJIxPYGbtY6gMcMteJbXGAPZUtenKuIMktgyk4mID4
zdcDxV9paSGond4EdBXRO0lh/0eqv+W0bCnADvWQvR8KybQIWnTWigIQsMCzOdEL
7D1NTys/H71pvoTkv7W27c4gycLU6urjJlDz2ZoxtI+cfKmdVYL8ux8sgwjy9S86
WEl+SpE1MGKjm7MSZ5nUmbRjNdj6l7pIlYMeEPV2n1VyvTIRdsee7d2Yi7oRX2KQ
HjU7/BZ6M9TVDLfGkFX4I9QD5pv+fiEE0Xbyptwlg/kr4x9YT9o586U7jVY+wk0n
YKx1paUbsSoDqPxmQyEFwL0S4inQ5ESQTgkGYC4ot1twsC2NL/5npzdJrp9lpIem
PMb1FbV1Gdz7pzuNwO5qounhlU/+uP3A8lTVBOVqqaoFeWDzk7UyjwTDCW+bvEfY
ruZ7SegMW9UYzKPoqBTtU9bjLChqM5O0le40KRU1tS4J9uVyRmlY6PaKIgvGLj3S
GgtJ4r1uiLeh9FhU1akIXFrCVUqAxOdU056uZeUlWPwELlpqqErYHAIe2G/GuTmM
cevm1kAVo2ScTvjNMH7D1986skAMKlpXfWYy3G3FLHjWDa1khDAVqBGUcR7zbLPT
vI8w8b3Lz6PC/FdYKJm2i6hQH/xpDBmqaU11L1YFDs/SFAaC6LHYFXMevIT5ryC6
LTzecCfjK3aYR6jQtlbIdGIFmzRZDel2ngcehAIg4Atyo2M0bzR8T0TME+Ud445j
ESch3nyhrKcm8+ffL/dNTpBonjg6vSdkOB0YOzFiFbWAMxjd0fGfpKHKaEZr8Uxb
trZrI7fbliHs0FVFnJQOCu4GqXJVsVatlnoOy0BOxbhJHtqcUrmhuyrnVGdK4PKp
rkvw4IbaOvmRXu/okX8zPz1KOcshsXlTzuKnEYSGl+o6HdNUoJilvaNVWyy2T8Kd
7OolHT+R/j5JnHDuNeYUMBQyUfGDBHgUYR9xIzwulEpWhpEOgR2mqowqWhWOoKax
Dm40nMd9y2Sj04SdTHv+46UAIQcfr1JASnCM/+3VEj81Tt+x4UP3SEN171oK5IWP
c2Or/M0C49WkQzt7cJOpFNfKpIWavNGp2kqHaiRUuKX+kfINOazXA01lGfVnpbpI
yFmVG5VcoIOjqB8pnOQ1r2RUep9Z+A3K7yOleT2IyYZMvM3Qvy9rZjUHR/FdxaNE
A3UmQaB7Uj87Ro5Vy0/+KjDZ7334v7NjOn/pjMxGYxWKkU6K2msHyq8QO2FVAGnP
KZ2NL/j5lQHHWixOHuA+FyTu5RpOWK69AVklSck8CsLP5SF3ZD3MYS0S4I+0UHtv
EqNeJtQlfLlQoVXdFvd2ErHchbUzElmKFHuEvXCpLuxisbz34W9xblkRUN6+jKpr
297OcOhvrWkVT684sZgDYy+3INwi2p+n71/6XJUBnsDrIZLOYOlFm4djz6bkcipp
UrNAVRFloy+YkoWF3sBHeXBotG8x26YWl3QEHQbWp8z2XCGBzpdcH90rmFJ0BaMK
LE8OURHjaHIWSZlbV1HZ0Y9C3l281LavvusKDS1YYW5/VA15EJYJxEiGxdB6lk6u
RGEfM3JHBd+yCCi8Fqt3vDXGbggGeLW4/qny5hAgIX/sDcF0NzES20wbiiSsz7PV
dAidw8YE9KPJ6/1iDPbswxo5e685PGBHmL3AgaJtg0RmW8I8GjQltH2SxVI884EG
oG0P9nFurKmFnT6R9ygiGrxwOXhNPeTDEU5UjWDj3fBU/ptA9Dkn8meBAHi7IUPK
JsImtaJxCfRo1mz/VeiEAmdEydF8YtDRHVMUr/0+na3g2RviUuZ0lt9Msu+nKDq/
Ih20YtimcSzXn2H6AL8HJcGfktN41AOjXJ34Q0q1s5lnIU9cPZn14BUvVGaU565t
GS2bcjN4m8X79Nu5RJRwAJUB09KVJY0yaVXS81nF3IEJqMXUCwcl6TJwrsEDz0wF
yy0Lrg+iyg5qR8ItgJNL7BghS8IegtJjHXi2EkdWncDhlx/BE1GhJkjB4MwOuN4D
K51v9bRJCnfsQrf323BYM41X+nucqhfFXluUjq8Q8Xp59c7QiJoaQtibDTNw1HTE
RHcFtg0up/zFo/86sm0DKMQ/dw/j6bNvDrM1X3K4pPaMBfowAkahPRMGYBVYEBLu
TQ6Es5wxKmBSFz3hU/zDsBppCinf07yWWs8brTYT+WoXwhJhTNzlPHFmL826yAZE
+4gyWnhGLMNKz5er+GPqw3Pd7Vtij44Zv5PC29W+9uLuwOw9aJhvIT7QHlrHn3aI
gJQnMY0xW0eW8HEgbPORimoQZfFXfbYSHFSwFQHOJuhp0QPL+wQgVZAAOqsypEpK
ao4WyFCyTYKPw+VCNQpZLahtIt3TCHjtP0rCLqvoo+vJrsfdbEiaGyf+bkDPxZeo
CksUOalXoYyk0jL7QjVqITQCj4RVVNEdt4Xlav2QM9xumL40H7SZvB+/EMr/ZZuL
YUNu4sLVB0BKc5QQ+/T0uAvnEszz7rHdUG3s6w5dFZ0COURpr2Hr/RxPtSdjvhvz
WaFmFmfU8j7uQ8tTxdpHQmLIJkB3fiQz0UjXdMFj+VP3b6eJmvNFwGD3ELK4ZKO5
S9BB1HeSb+rV/dOJXTdAseR47/vOT2hPmKekCYNtwrXegzGyKG35snjjz3DiWSmq
UyIouCy3FLjbmlktc+HGQ4gk+cT9rdkgOE6SyQWa/IA2D73xmv/pHEZZGMkLQFQp
Tntoi3o0k1OoNtj+sDQ2GvYmb1Fjprqq6nNkJXD/f0JoGyxi+8MNIWh5AB2SZWAO
ksuvbahDpAL+hxeNBAKc/01nwTXjgAXnSmTp0C19U+JKQbe/8PD8OX3lk/uhjHVd
2OW7NbmpPezZXRwAihYtD4nS46vApVcS+FujuhwaQ4+Nuec3qQvBe6AiUj2leOHe
KeVh+QuU70IcQw0u/5RP4Ti4B/1XJA48ksETBNmRa3un1y8IMKxsmZzIKP6+ubLS
GuJZXKU+yaI3NUM3KR7ntCk2QTqzBKWi7HX+Jb2bMxCpNbPA10YR2G+nzjgIVwho
wQxC3QuLlZLzj0AM3sGC340kFoeXYJVe5Rvln6GRfPCUF2YPn2gd2DlsN/6iboBJ
uj5nB9Ipd291RogNjSsKEKMb9chZNvAQ/LOmVhvOSTyCaH4okquyKvfI7L/DBmAP
iagV4XetR27YQbeTpZDcq8WU63FPIv3u+JMvOx7BpQF8p2bqeZsQFCsR+bR/iGOd
OH1gW0cp/HV14n/TjksbS/iQbIJi1BSHKz93kLI2+fxa10cWrVODKpOS3p33Xljz
3fucXHvOnk7iOgc1sTHh/OCEhURfHxNwuUm0a/1fD2jQs25DD1ksjWMmyb5hcU8Q
rS0TuA6Alayb9KxsmsWR8MmYQO53Z2H6ZPOrHpQpvN7rvHO7EpWUTEllrd545wsP
VtWLeryDyc+Ma1AMXSbdcGr3dAk1o8SC99DbtoobGifnfaDjaWYhzREH61GIoutX
7y4uXeh76AVIsm3l/zszM7xRpS+k9j2+b4vw5vLuuYUG8mUjM8Nkyj+P9kDkjMvG
mVaeQhGTRlhUyRnrg23XNr1pgjICZ1qx4rLpzINnFRJEzRqPM48CYvKAdh7zNsTP
xoGHJJUB9uT8CtvcB01X59HaD9V2OHZfzQrVG9vYe7CC7tWaiPwq5MI58YVxHi/o
byNyx6B6EYyw3JRZtqdA9UMbmNOMxkNHYb90fDagY0vDerlSaRZyXGE7D4OG/k/H
JSsOo6tg4TonWdVDJhjnorNGwbLeBuNe3wjTsSAYRe0XPkbfp6YDAD2t8fZ9RnWq
j7jZe514HlrCveBWCAOZdKgiteLUczjBoU2oZGPWn9AsL9Sh6FrGb2HT9tdxyeYq
n9vdt2WjOp7JCvVLKN+f3psXnIPzmajPW3MlZ+4fSvHmkAvZJYp1Xs4h6KGhH1S4
zdbIWSKdbH5RWdhY8v6V+oAxYyJ9eX3Yu/G41lsHVhsMdRXDfSAZVCICjnCl1B0+
KXWwaV6f78Ng7gI0xKJNSyXMaljJ/01qZOe2u+yHa5s+dOX4tcDjJoyQL2/XOdRF
jWzjAQBLfO7So8JMX11FX/Ah5HyLLswNW+12z9rsiseXrFWWLPb3+BPSkpAHrxi/
+409mXCjXxgFG1z5kpM6jEs4Lytw2ZWOF3JIFdyCnF4ae9s/gmEsOSd084xZVkF/
zCwG3kGV2LfJI7cMVjvDmHhgR3vgo0val9n0E19yBH8U2KwEADOV25SXcHKCsaCR
EBHie/HHqm0A5ri6IZliPgRRa+A/YXmJ9lh2T+9IgPlvZY0nrIoRYgvpOuex+x+Y
VgCN+oywOvCemtgQhRFPOe8Wh6t63TpRCvx/0YJ3EKH7ixhF9m5Ui0GJpUcoMSdJ
sX1LxuSsuyxXAq03Zf6WTrgqse/lu6FQfvqBsYr6vARiYlyRfosoFblFHrsq5JPh
GVrp32y85c024/Nv+fPgrXgM/NFKZIvYFtHeXGYBsD6ZCRJRuTDbS2iqLmJB2lLV
FjoT8xienyIrGgMxK/by5Ax6U68ouoWELUTEYH1ZenyhZfmCxfc2OghYJh7ogTky
3xJlF+qYWp262UlJRE4VWb2W9/Irqig7HPhS/mRyGw7Q4gvrCSWLwCAa8jn+ii/a
DGREtVJd0om7rwO1Ok0DkUP2J3gkS/xzXmGKx+uCGRe8h5Vv+G/oYYr0vODQMEew
HETSzKeRlCbguzXeit3dOyCePm4x3mbyRC9YHeAXo1mAXSlZXawYqXE1gY4Xq0UI
ZfkeoMAI3kWKmFY9nRGoCCmQbWw3IQmmH8pmoyKfKC3HDvvSStGzc64WGzQQBClw
Lniz3IdqdClK3Geh2W3H34gT17VAZvQrR5qsJH4jB1X28OZNaN1SfizlVByOeXzE
WrEB0DJN7yaf/25U2oH5SkiDTSQgkbbCNi2Mo8skE1r4t9EOiQObTbMhQp2Nk9Y0
ccpetXgp+WlcQ6ZJXxSJdd46DeBbfRLsmSsVth2gl5lU5u1MVFqTmTR7trq4Q7Ua
4H6Rse9vNzED822+h+5MB1SPmedG01pjvAIw4VXDGR3DPcmKWeSYSQ17ifphLhLC
C4K0xZXQImAJ7aAaW+7beL/0JZVZnnc0khItpSsmS3nVATTFBdTNiBG8Wk7e16Qw
pzamywUc5TUW9JoINIqEUs/lP17YX+vP/JkJMW1SZN7KAuHeCSIYMauNfFudMfsB
ntRoWPu+OlwXNjcpPa924NM+W6Jlv6dWrmcUwuXVIK5ggQOY8IVLZQuZzZABYSKX
679B0zceKL9rslD+RRHFKe//EDMNL5AhNgWTcRnEysYtnKF8KRRKzFDR58j+eSAT
iwPUykouaajB5dbTCFyKTm5l/Y6TouCsy8+/AyNEWZjrAqS/7vHFTZD1jZ5gLxmF
XI8xU+OxAv8g5J98VobJCuOAoxnJleaycdxvwByBFnZDqyAYlTU+TtTuMeW+Dihe
YbPyt/NYVlfnW5neSOLhJMeWtCx/03NMHH2uIBtMZ8jCjcxgjdiUl0R4v/MXpxah
mwDcKYgZmam57+jVQe6RfCX2INIWK7ht0i/HVTWEha8s+hkV2h1JfvC557jDQQM8
PnzJ9GR7CFMe945BnXdeZeCjPCS4IomF/LvAsVhGjrWZ1ao+r6HS5NMzTuWYqQ2x
w5XFCHcVhS2lYZu2h2GHSURCWsdv+lasPZ9agNLwVgzcVX320J/+ZzE86t4xkohi
6T7LJjtPizXN0n9UVOMlXOh6LjYuSKjuvo4DsBRfDUYzbLQ++LD57IAlHr0pgf0j
Di3Gro5tPEnrEj6ebMGhRnYy9808J2MdNibmBRWVXhx9fl32eZZRh15AjkiK5UpF
Z8LwF/fx/u4I+8xO6vP4vIOCddx4gEVECfW8kXURCGnGnUK2jEDrOWj2gtdEo5CO
XK6b5jSMXlA+tSfiEKUV0gPnltX5m7+2K9W9h/35b3PAuEXkOXKkJONT1G5miZva
VSTDra3skJd5fkmonGTiOzyyLx+PaWa82zE4GztZVzAFvSi0i9kDMdc6dnFbsMyZ
itmDmq+R0eMd2GGheFfBWI2oM4RyE7IvuGMzQteq64nBHUkP3qs4jilyI1WJ/Cnd
gLLIciqRYOAjPmLhVA2ZSPGnnTsMVFfbYW9tWxETFymMsVQd4h81zp7KAa8LGILy
eBGS+1abkj1+27E0vqL19z7Zl+MF3wB61IhxxvDJfp703EUU+tyCoR4f8VI+Mx6+
xf4j+jEo3Olg0b+y8QiMhrl1z49TpwUT+HNbUaO69YJWyjNxAh3cdSGR8SlR4bEq
P5cDXGH2YpJyvgCmZ/zxpAd+mQl39WWE6nX7kuHodvTzmCyAoxJx9VvyRwlyv4li
3sZziRmD3Cw5xwirkGvggt6dmBO0ScSlGs/nD7rfhsQGuiol1ggkfNQ4/HZZpX6R
MxVCCcfJ2yrrGZtNzdDScmxQCr4J3TmP4RixwCS3boeX3VVLVkG1Jsy45B5df+6P
NiWOapuBO3D7PK65kmBOwnIJtqWkcdZ745G8Nkas3Cad/4BllqDjm2G6WyIaovND
YMcX8i3HEjjEzwiVReuEYwi21+aCVdx2/DCqe82/667IwQrBxny9joA3MJs0JQzt
zcPAsqNQJNAseH+y3hgre80IywVHHjjovynHNTIjVKX3u6H0/G13mEAYTVJyFob1
t51GWDigJaZ0Ss6DKbM2u5K2rp8IrvOtPzrLh65VuN75I8LDURGe8GqNO7q53/VD
P7Cq5mL3/B3rG6i6eD+QXICbl5vgVR7DqbygI8E9UcuMeZdrVb9G8J2cAEJDquVv
9aKyMv8Rsl1YA4R5aSGzVfTfrwIOYzVFtv1vpWD9hKWjZCDGRqbLqY2WOgMefkZ2
DCV91gf0tN3nd4uZlNg3beD/VS+wYi4CWCZms2VPlDLCgJObrTcl676kFDp659Zb
+cH7Gsjl4I1i795JH6oCMe+WSr8h49ctp8uuRtjkRHk+2KwcMAJdSFC8g6mM5fOA
vyNT6nfQhYen42+bU5U8o7R9L9snIGH+oYwWwrfDvCQXfRXU6GMiC2bw6Hl23X2w
yLnQOf/MCyLrMRp+QODzmO+4XwStIWmJfhwALTybYshZ6mmW9RFdeLkxMKxBShYB
5zGq75nsGBp0Qpd421z+uqQGDLOadu488mndh8rPiYIGvvoEHUMXe5hoiBM7LXU2
64texe0t8zoCf1C66MAsM+wbTyE5R2Mc3eOX+IBBI2/9JvZ95EMImrQsMmwYRYzC
fFfCr2sH05t0oq+hQn1TAvUhRZDXsIXkdmUYYC1/QnQsVFx1vRzRfKCytMw2jFKi
n3EuJXvWZitBQP1+PWHjiekfiHCRESpAAVbC684pOTsQFafs6IUo/05LGyTmJLZF
nxmnf/TIML/Zmr4lgrbAhYLoIWrKo5xXFmmj54Umgap4b3+sX1luLXXrOQKCNCAl
/rGxFe8BUKUFIFrQCYXAAT1zX25N+8yR4bOczq/1eziduNrz0FRtcfzKYlFJMnrA
4r0SmBJI0dzpG+XdxpHNo+8ieC4KLzGxop9E6+IVyb1RI4gFEnX85yFKTujzADmg
Y6m+kTZWz4GlH0Xe5YOxJHXKradxtgGnHBfQT0yRA9eS1s/0VohXvqsNA2g32vX0
mWuEVIsJHL6Ab3HRzjSeU3dTe3WvLl+YNtLrw2rF7FLCaC5Y6k4RspnER5emND68
xQ9/mIKNMACxqAWYBeerv895mq4zsGhBbmAxLcJdup1xjFohqoXk2AI2aIg4oDe4
2E/MWXzfDVqoQOhGRSQYm9TgYmdYCGTzFH0ROC1czlGEZ9bUc/1xMQDcaIAabWB4
1EDr2oo3+thrmNZK5Gff3foE8tHEy5f6g0lE3LHCfKqdFuDWD0XoqMPw52R0a7jf
YLJKzwqYPKlFIKUYUzEbb+91rLhziamqxJwicY4XCHiuWTWfWoDATe3l1p+MVKR1
5kVkQiF9Uv9WTz1m6f8LRhsVL7VB/ma72Knv8uvpW2c5ZOvK1y6U6ureA2NbMjF7
nRBODXSf+k2BnKoXWzs59beKyAUerREkFXB0PiP+10U+Rn7l66/dFjsxg+CUKtwz
UQ5h1/0KmCBzZleKvaAn/1u6sTTuKe+TATH+NanhXvqElgjaTieuGf6ZQnVTY96I
b56BahBXsu7SpcOxPMdyDD0O/RWIAh4G2+jjKtRwj9zdwP/2+Ne0guUxGtd7OKph
Tacx/+ftULruI/w/05qYVKXJb0jIzaP7HvT4oeOIazkqqya6TJrO+4YhMHDRNdI+
fWa3xC173Av5Ap/KgjG/uxOxRpcBV3BKnzR2fpsbPyjBj1QPKYhY+9jiW/pbJSg9
CusnR9L7fKfCKTe/V8p2n+MzOIRQqTYQrNhx/WP77pCvB52ZLbT+cDD3Y4zLv9Hk
NEgtmC06ETEPGQZysACVb47/81V6WIws00ehPmNupksrts+6+GMj3htB9mSLyhIT
eGGgmLA9bf/gpSn7CDTBbhhrqfBFefRPR1ImrpmWTstV94XNwifkLU3YSyUr3c0M
1GI2t6yZ5XRORvfIjZQCh51s3Z1W2PbJhwfmP3ZnzmJ2ET3O5LZUYSe4iS1cQw5f
W/HdjQxkPvtZNflKrqzGE59le/nD/QbBppSvKO9+ip6emkPeqB+OdY7aek9ArZHt
rgZU1m8Sc/g2LjPc0jMev7uoTElI77vYX/7s3rcloEeUrIP7iNWZ3auzdCZBUiXh
E8lF0xnb07/uGX8zVgoTRVfWGzMzE0fpBnNT6glokVsyEt5oBslSUllM4zgxFbcN
cTHW63DmcGLB9WMiw+2av3mFRrtmi3e8TSMLsqFqNM57vz4NorXnWWs9qX+ZnVBt
2bK5RHW8N54p4YRZxXPk9Xsyf9SagBPf4YJGrej7/joWAUEWshxU+FX4fKAVS80w
va2Y4WcPY95LENFQ974xuf2MMc5bL9kpt2ceYe6SvdF2YtJ5+a1IQ4W58vPFIYQG
behYlxk/eF8ER3WvUOm1vieHfeb03Y7ies8WVtNvZiJivsXC7PjTvX3OlWNESf2X
krr+raoW3gE8Yb16w1uW2y1RGHiNbChDVR3kdEiV6gtrqRy/Xj/v6sPizpmIikvO
8ueRxmySsHQQ0ihnLZjkiKkdVbCXbn3ErlYiiBPh+DWa0pEeFxcMgubBOjc7CxI5
yGFxuHNXxoq70G0zPTmFvYB7NotANqh4iWFlW7fCyihbahaMWM4hsWvO3VkQ/TtU
HFeU80ZDY0qEb2QbrUaQyNazEjnlbJyxMOKCEZKQ6KpVnr73rLGYEJWsUPqm3veV
8e3etik+qzEhL7mfiSs4NMi5Ts3w9HS2QlL3e40iVhdLcLm9jO4LpIakhHmnl1Lk
IjXKRkOXeD8FH1a7Dg0zayadbD1jlkGR3G92yw36/XgYBYY2yqkPR7uq1U8BN/QL
iBZtEpfmNMxwNkrdbm0Z8FXs2WHlVzMzXXVZLUFsksGT83+Lb+LJkpEHdtBEHgs4
C4i6iliW+1uKyfMZQID2dv/svOTp42Zl9+z7IO5rWl/WPAisl18nnh2N6fr3m2Y8
YnK5ymyHfThF8toHB9drudDv/sjpU+lezoriXXDqH+3oEn+fi0JPTSmdqNFZxSzR
9F+Zj0GOaw+Pb+fzlMM0eyvfvzfDi2Q9gUWwwaxv6r1i6yYDVgfG85xU73P1Gm93
Wr73Lf838hoB/sObt1PUy4c7FeGDOmlTghYbsKPSH1cWEsQH6X7tHiT0VE2VuGp0
eGDlXz3Z8tfwJegdSHFKgkGK8PIvVmmsxsoUc14QouwdmXrQL3m7F3QcAV5t0Mcb
lhpME09IESrRE4wsdxAL/ungNEXUdUjwAq8iq93ismPqqDShT5MBy+l5U5ul3P6u
8xSUMA61ffoVjiOoI0W+wEZzZ4fRjVJmqNCjnfWs8t2RnCCIrjvd907u/D2aTxNL
YwXOm1ELjIJ7ZZEkLf/xE1aAtrRbG8/uPgfL203RgPBshPL2mvmau3NRT6LFe2io
DxVMjHv6eU9olBTmMozvE2Es9wDkBvzDufVJBOVFMSuZqdkhqem0xiIT9pBQX0l3
BCrvbIi/WmrOr9mMav2tX3dw50+Fi1lFjrfj+cwmfTwezSC8BmRRvb9VpSQ7QEfQ
1uUwlraHtDY74MMxgd0TcTnHRpB45WdV0KWeSNKa2ff8IVD59wJi6V+Yoj5Ee62e
6JO0ASJSasMSRE38+KMMGk0n9tnPqQLlzOodVM8i8bphwMJ9N+4u+bYY0AGlN1Aw
IIwj78gM2OVHZygeNKspd97psHEVwpKbkbtkZ9dEmuzGofHVJ0j4ouayTGnpMZp1
jkmtHaYVh9cvtBnODTC2kyOG2N4A7a3wTeko1R8Zil8z/jbj7F0yV4zl+EPmm+FU
RFox0uBNZnJ57kbAuGE+1V7nhS4q7XP+GoYEpY6lZ+TFzr31yiJyUMNbQW0y6sbK
NX2h4YoeNMTT3+ECTk+dJBPYWapkRdqZGR5HEuXStdrC8LwHYx8LDl3l/ZQhLQ11
U9sAXbsFT21u25CpMPHn9NyaKVFh3H5SFnWPTvNI3uWIExuH4Yj7tPlMlfOAh1Ed
LSOGnM+0QmJdNO5dGCyGfqWxJODv215rmtu7yY9bAY79b9emUkdCaL0Y1CqVvvOl
6eLWaRxJmSJouaw6+bbpXu8hs7ZTnZL70QhYBqfb3zptRCj9EMqC0iIKYO5BRBpT
CwcK8uQfpeoHNEdMoMEcu9sTFHJZjklVrfMLEYjK54GwVZpatFOComf272f8zbDt
3+x30Cd5T3bjj7Dyd44YZSTuwVXiepshxc1NmtAQF7G+mVQlJh1deJsPp9DLRFHA
lqJzCpAJwbAgxpDLnLhdEol+HYzngP7YuvtcdTHUlxMooJRmHyEXe6Hp7TXK799j
tbWZJEmvXs0dETdZMfWu1gD0DwnqiP8ijik2pMX2IOGth3/xOBRld2Pmszfrclbc
5j1lpGUHjjAdpqD2eYVkyuYxVmeV0APVNWy0uV3Z7gOen7lveMjL0Vg3qEww2Fxp
mHQ+H1/HiJptcw36/tS/gf2DTuUOAipLu/FSclbXBWhbOfpKFHFAD84hkzAIjAQR
XdIw7Bbj19dzel38PbRs1Yepgm7eKCHzMgObDW/3q9Ir9UJm4gPjeAkBeC0muXce
ahsb2qi7AEe5428XX1NbxeeusdJ8EYPIVoijoekdeBUlzr9lD5MyiPgIFVT0oZZe
LKv9MnvaHc/Z+GoytDttKAcNy4dVdnoWb4TqrzgIPo91DXPvoj8LoadLWJVmAhAC
F3T+mjotdyEIwXsB/GVHkpNVVqNYnPXtr8bKaNrkpcUU2ZuC3GCZoh7zWur0oibb
nxh57ddoBCXAsYdbvbWj4rLXbqDpAERDk6tNTTcw8FCV+EoPJfdQfeHeMv3l8qhj
LHOgY6SlZ2QVZ38qT2wkP08xDW2zvGYRUmon9WOshHEdwWU/UHcUFAOv9jFLUklQ
Uw7MWoux96GXcjIdw6CtewKoUmuVGMJ8cVzCTkf1B9EK0Hjsn6ujM4HJZq6QxdQh
7RZ4JhryPj16Z9Fa9M4i8bJtIAiRLSoUC1m7RhuVxqZGesGVof4Tc2KhqCHci8n/
KW4U+/wopvNXkx1e5vW5aJ9wRIinySU7jT2Fqvj8KoZHNgKJXGSD3CkmCCDxBZQ1
OvhL0nSQTR7v37Kq1JxTCYpKZ6cCLOP30HQkNGi1k7CpvwuGHr4FL9aITskgshlQ
6zkGV5kHHXZoCTIdsf5VVq2FVDc8Hk7fnSwzwo39B66nGtSkzqhwwm6dGxwj4RBq
KYabetjdbql380uSXnBefWFoNR8shxvRyn27pH2LcDm32WBxrVDAvI1LkaGZYPQI
MWEiS2NWPtkeUTl+Cb7844offXu/aQixWSxC2rVfgu8+KSMkpXRVjsmfkDy5QmVB
JKyqwsWOdh3rXAK7DxpoPlKWcM1VXvsQZvxihmbpG8ESMywsovVNl6TjqIvCK+Z8
ckGwi0o5jO6cpxXIHTeo8x69s9f3i+JK4X5+f+dT2LP9t1CqMP5lvUU4l3OX8GT5
QVPYpTZy5ADNxuv07uqSEtcGNgxVjXuUo6uLhs7Dg1o9AHhAxHdn66Vle93jcGy+
D05jKmlq5uOWpDNKV1WfueDEU/RJUDKVsOmx5ChSh4sdzgmQ/VSJtutSKSJXjkSS
pHUBaBAZPb3Smcn6cQZC8rxrBjwZR/Vk/fT+47plDypDEMf5BLPqBVvB5FFnH1mz
HSKwkVBhdH/9xjPFIbgBxpBA9OmTwVOmoam5+P3XddlvC6YNZBBp+SUUwnMgZQ9h
1c1pMDtCFHdBXcvLSBzygxLqpq6gfW0vsoniz4ODN/rgQn3PJTl7Pb5HVBWKkxno
dSWbXz80y4kRRm/ILpxcPjWneUy6JT97cSqo6/LHG7L3yz7ju7anVtzgpyzitW1M
CqilYeaEkdJHzlZQph9/hIFe+Tp3CIA3xHFyaDntC7CVQMVXL5zSm8N7vLp/OszR
erPp2vUTlJWKk4SuGbf/E16coRvak/TE2LziwwZBcUOl9oM67r4ngQyw62GHrlFY
6k0NI+b/eHYpYdPFbAO3WNsQDfXraLyt2fplIZjMCtTEZNhBWS8ddXkLczT1z/t8
yuEHvnK1JZkg3CWwWri5sL3tfYluyE031wCahdohfMZX24+Aw7IjhfJ2WbrXaHYp
BBDxOpPxQEc3xC8Sk79dP7Qt8hPllWydRvlB3DSCYwAgBnUL344Cmy8Z1qU6KYe+
/4zU5QsRf68e3luyllHCB5PdBnVgDyhmjZsQ2cHR5MBeKIUfgajMsAC7Vs8Yo0mc
NPGKHyK9SuH9V3rT++4DU2vy/2FE9FAuXbApwb/c7dM7WlfVve2JulVYeWM9jAia
zHPB9KE8qTwLrsqBrlHRco6XC8rDKdfLu2pTNJvdegwH+0wFGMZpY7Gy5HtAhk7Y
3SkKWkYqBpCrhgdaBYChDW1DfI8ETJ7cHfHdYHy/nGF7GJP6CyD1MkmOVQ1tuTAa
gs8D/Nb1mUEOHbQfwAuF9kBpr2ubjmR9HTKPJCzz4g2gLMkuzTYZxTbdtyM7+VKw
FwqBt5ASJOhwiLoWvmZsqBGGPsL1w3zDoWom/hNRVH9n1ggnZKKCz5Fra4IBX7hF
+PFJsp1OAHpTMIXkFQJHN7hQO/tNfcqFZH1VUIYHwQDKNd4Ja0wGGsHv+tGNLw9c
M5UT8K4Tn1z0XXcDVIoJH55tzATTGtH66qCXnWoym6mPdIlfxA7+11neYtE9vpib
Sn+YydYDO01/B1uUPNI04wNlxItpg3uchyd1ZW/KdUhzyGNBvxLwEozBkVWM5UP+
gNc1vVsAttSxxU30ujzWIHjBDckT2fOkDy4Dl+xlqA73KYTORXXp21+6WWkQdJfU
GsaAECaeYLdMPal/Cc7r/lImI1ATVetGJ/qV+RTofWLiuEcXponqOgfEPZxOxQC9
FMDLRlD4zcwRn7YlWTyk5NZc0Y4cL8eSh4UTlnViypuRfer3nuiGCZW+8Qa10Clj
d/4wrH4T0yn6ZLqcR6bNJxtX7EKMXUg8AX6xlQjwEKfoiYE8Z+namg8YrcquNy/Z
uNtPRI+eJnzEpiyBj3s5BfuOPafO+5HdUfUImJdO0WDKFt8ccCCPz2Xx75js5zos
LKZgZoGh8dcztIRd3IVM+leZ6nXe6mfJ2WcqgQoiv9U4Zct8DB/lEfQSEgoTTaNr
FhEQn0x/rMKKbvxeOCubwwrGv0c53IOzFIbjB39lQSLlaZw1UaUPIWrR3fubWP6d
AckXNm/aDiQLabtq1zUSTjhWW5Utt7VJErUF/0oO+CJaLa5MYcO7/i6gt3JkEnqg
RnTaE7rgFwHiNrJdI4V9Qmz2sZAatfiZUCPijayjDAR55rtIlW7y8IA95P3LFNgO
0C0nH3yzKDyuFwFzo0b4n4dTupfbNhN7Ti6Bjnei8v12ltSF0BNwpWq0zVDqkeyr
vgtLEnEK5s5SDIfkOpjTX7EWlCr0tCSNiWH/JGGfAXAeEWUwPVnl7FqrqgwhdOZ4
VEkaaXCwFWFLcw+psk71CI6ih7qSB82V60BDfAZwkbH7Gqn6h0fcxWh+UbV02sI+
P5OqExsWNWM7ioegYcgP+E4B1dnDiyac4qUG1ZCsWPQIFTZOBosy9i9YTadox8H0
uOXOOchAqOwpuMVSOM+OKYOvufdh/jLlfeuAnyGbJYlfqEcdT9FspTZCYUwAj6qE
vOmXy2Qw+tzLcen+PodbsyyAC1I8/t166kzeHD25sdSjxZqIHCeEMT6ZJIPzmvD0
aGzpGV6BonHcIwTiUgjKGDFJtgt45lhcS4w0y9Zxh+6ubhawDNSVVslTUtR3A0eZ
St2N/cj/94UYyxji1nQYybAC8WbEf2ZdruGvEx5nl0bvkWh3zlg1HzeKVsnayUWW
9jxH1B6qWAz1MUrTlyD6hxxUd3nuIkSv7SxICsSFzkdQD7ZqUqIcrAvelkOCh6WM
fsNTuhMxxMOWisRgRHK6/h0rEGKtmhuzM5/PezKmQgz2IoVe1gxZ986+wmgSLktK
6HyuOjkhcfFSBSaizVHgQdD6syk4ev1U0+BmKebGyjb9I2aiJMso/6J/qyiA7TfJ
Fvk23qDD3MrNBIcAOgANrTaD79hW9Nl5g7kDP9FfK1DL4LXii0SNf5up+rqdT2W2
NGDi59ajKFPHOAC3nHUsmgRQZcOEpdAvf/saBDE7MqnADUQzC86eB32X4neG7DHc
g70SZlGl1Aywxm3CJSsI788JsgALlyD3sN2JsDR/CrGabTIODbuCGPVoTaDAyxhW
3BRn1dUqnVSlYZH2Qgil6k3EAaPwLhb9gZbhCTkE2TE6wFFXGH7OQ/LV4keI25T3
Ccm1WOd0ScgdXoeMPleGa7+yNcuRO/a5gqEScJpRRfTnaU0MXPSLYMFdOIckvOLL
DFVXLYdHKnIyC84CEtlCSF+NQS4lkG0vqz9p5tvHaUX2I2xQ9SudH2jCA6PgPQrG
EGtNTYeKscMsBGKGEv9kVwceoTJDu3ofZ2Hcz58P1e+EPHQQwo9XHbc5djCPh8ID
Kzcv1YOx9by61+CzpH5TXXnhreyyBnT8JcIpFpa4uL9XjwtE68SOsuQQYoXjaDSQ
JkgFIEWPX3nF3raJ028JzeiLyLnKFPvzFMR+vIVViTes80CK7Ky7ocD6NYJ+xeLb
HHyLfAOnekAAbzzYVvubUWCWh/JAj+pm1CTB8Miv7XS8rKKJCwzTzkXAz1YT+ARk
HGHftcbsfPL5m2AMJvpYk0lvmpI4VhuWmCTW6xxHq3A0JTSL19UN5kLZW6ZZ6UPr
e6Tng5gJDTh2JXQOEYtGICXNWgSzr8svUp39fEz3uOkOjW4ocdKI4f58gv1eKRqz
U2YFP3ChjM+kFYh6GJANiWvaTR/K1d+0lrWesAkzeMDSqF8CErc8L/HtUqt8u41i
Z+seC+3v7IftR4hrUiWH1O2TqcuqR9XEylEXNGhNBJWIG6SY0DA3JnhXVOBzuqON
IwAHiSWhtJ7gbANLR+uNI7FNQcEqTmy5Ad81v6rTnU2zBmP4JItlb2Xc989ZEXiM
xCQx8Tgo3lt67AC/X1KJP6UJc1ljcGllQSlUTS8K0zugfCE1IhOggtSXZXX80+8/
yKfRByEpb8MRbmHzI0VDR2nTZGR+uK1i3SEfLjzw3FfwKX1Qwx/ItVHg3/cxa7E4
GH4pMIl2GWfsC+ef1i0+f+wFlyWgRrLBS1YVNzziFkLsuMGKSyQlJfCpeRzkhD1/
GiAXAb9IazX3Nd1VkCk4pvjSxgjG0Hm+2ddXdv9p5wHgTzZ0tpQT3v/ELbOLK/UI
LEySSNXhZP5kb/VJkHUX14sOYU+VAQw8OVCKG180fIeCrvMIqGkrLmL+X1ihUCKf
J+IiWBRdrHdkmjsegz5jzXDW3sRX1ul4JAe/WPHfJVgMeDnaAc3V4MNI+OtJVaKQ
eHC8Zd3J5/j5hqfXzi5Lc0w6GPEdR+JgPiusKcQdkMkNPZ32CwcDr7MaNyp2sQuW
UFx+nQWmwWbVRm48i3IndkJ9nUx2reScLfy4d4jHlJu7YEerl5dF/SGWZcbzRYiR
EN0EUKJsjX2QWbzXxtDADzDR6dDZxv90fP5RmyJ+K2Zc7mfweZYv2bvtnw79p/B4
XDQ0ub90ZzT5W/nRi9ycf4ZO7nqKUE6PIKELj8i/AaShBQoybD7HI2fV5MsJxufE
Yzg0Y3KEmpf18TnjF8ZOtlDPNdnvMUQirD54R0iYSWc4/Gg5OR2+3Ftq0ubMxGjM
4/dKocgEV0Vd7MpF0Ta+KO3HjnmWCm74JYHepdQNuhqMzIh+t9un6G0dKiy9HMk0
xvqxafasK4y708gBr71f8Q9bGP2kD0jb20Ncea72gBh7alHcarnWCa2TCYss7rGs
dBfLGjmLoX/Wp3ic1AQvp7BRLE57YrQ39HScS/BT6muIZFSibD1NXPkrhuKuiMqy
wgmF9co7WPGbrLbJafZeHpFGsiRk2ojTUGbKTvARVocbSm9ED5NYVkka0w1qSwl0
f4UAV7+lfyOwY7BXkvXaWO9ZNY70DZaNdntKHIVp80zCE+vZxkrU4HIaPlb3yiWC
M0nQd5yoBSxuEYQiYnjeDyyt9XbZXE0TNyLTvPZt1ZM3F/L3QDhny+K6o3/M5ET7
qYChfV0L1UfH0WW/2/OKQPWNABSgmLBqWfRVIxAvNDRuXkEaNPqDFl/am3D4ly7m
/UU89UTjKDUWJu3moqq0xsTrkwfS1MC0QBgZ0PxRyXc0daqyby9mTmhK6YNJCfLl
TlF4KcE3obfByRyVAV5elhbcgOZDb5z2MBtfxEg7vEI3o0ijAlRt1xQHJRXvPLt9
m+0HHAuiTli0Sc63RIdCb170/yNqf/Pqv6kvH3+rY3DD8HkxWTTgHNO9EgTcnDos
f+HiAei2PMhv5eo5Rfu8eAozOsMT10VC9whjkED8Cmf49iaeEaaBaaVUEjbL9nNv
6y4NsjzBWNV6WmzNeE6xI1JiXnH8yub81VPJnP3o7slfqpVIMI5LRuERFZIl7w9a
WTmsarV1q0R3zX8Y8dXHajaNt3uDBcc0StHHBWpcx1H0tkra3AqSsyCiIsZMpZaI
c0tkl9rt+EPZbcnCLeShvoYbsTPjXYzG0dCu2RBj+T7nL/QRDtLQcCInJ/edE7P9
8FCGSo+NYuzl2upxy8Gnsikx5Ub+K+HA5g7UWHSYhuVvRcIYlt5m68zgLdLtJOxc
xl4kfWokyrX9kiLg2Nka08zSTzFQK3RlfmvFfsVCn9/YRZug3WEABoUCUHVj8bMB
/oECocCobfpKZPstaWGjYB/kyBSjykwjVPzVFad+ntrM/zC3SfY1mRKXah4MYV//
QVkpZymrMjcBa1xiiN4IgOM2phjuRtukV5iEeXfFBwPY21m30vXxapPe9K+O1u9U
kQD0i+Dx5qxQohY7FJJpsW6etJy0m61fG23oIKowme5YcjCsQ/B+R6fkvM+KirJp
ubxQbZ4GIMWA5sxhc25j2iTGaswHdAyW/LPNwigja9RMDatVs686Wp1qp1jRc6/n
12Uh1A+7Imoe286YfiyfF9Ory9Yxtvm4QUbKwGHeYXdA2d7RS6vki4zawGl2CPAM
15TkXkhzzCObEdXYNWECPZ+UVGyMqisCWY8Di8w5h2fOFOCLGfoGBd4Of5bEQk4L
/g3dVG/29CQ0r5wxp+0rYKxVidD+rPovaESgzbVowIxvv13TMur1IFoWdud4/Qnu
9svk8AbvIRn6dBo1gi/Lth+Zfyvnpx2tkx1UCrWO2I2uhDbDj7dyepf6pu5H2sAj
1CRH5vrEBfiZZUOpgGJMcWfHMibeNqAA4iyuwNGbOHUIFNQO/C5Gx3IkpNf8zpXS
iZEo9X+AcPoZDCg6HgdXB+jKezkCarKRXUSGCYxN4W4igtt3widu33wpewxPbQIM
OcTiyqzcFB+8sXjdOfVRQ6CxKDaZpG/zS7Gke0BVpwPJ/4Ag5ZB/NqijFmDBaQ2U
5KoAndabHl0kIXVFaMMLRv43aqM0Aucd91YEWjH98JU31FOisEvrMxbw9noO4n0x
lJeuciYVvNmG/C2e9jH2pbboMMEJFd2EFKTWwjlWhwW6a67PQbk2QIbUuzof3/8J
W540fpr9ZpXqyzRDKxl58EAICh1RTTejwGuCYFMFCSDNX72UfOKgvcF475KzxdZi
CuiKS85Jn1/TerpccGZlhEGXIXPf5cG1T1S9+60XBfh4ipTafR2OFEl/JBXcyyaW
/gZUIWcC6/0MoR0v6T21iJFXRS45W41WtnjaeZ9O5Gpy2H9VykrEutWkk4cpRssX
53zDEIsen9uMI5kk2UGCN/xpIs6CecsPIaf+tTWrD5wGKwwhjlbyeQvwe/caxMiW
iXHqvvKU9lEnyAwVagmy+m9KmYm8hn1SHsOLBeMFhPVLpcjGsQzH4n016HJIs3gT
2+SebBuvy6L1cLh8GMQG442We5N+OTcMn0AyyBdgPVSsxwUyU/JdeKa9XEs++3s/
KgiOPKFxs5hgyku9s9Ox8fwoRp/Ng+EWzz7G9NNBZ4Y6hsWy99IvTJURUiwdLxfn
KdcAAsvn2mfJp509BYZIRMggvSgOc6qTSXnVFSEhxztuKZ0ljTj1eUslmmwvNnSs
2SUeehc1RnjlQV1iplxD+8T4k9Y74IuuYryn8vHAQGlxCii5k1Bl2DPZQC15+KMN
I2CcLTV6xG+V8uS0yIoL8ncIElANeOuZmjFHLrkTJYpBoqMrq3fU11x2mZwgVo8q
8uXuvDToOP9u2dkn5rGjEIvkj9FuOC9xNI5+zGzz3vOl/Aiu90JhA+tGbwHJ7/YE
MzVoV4d+a40OGaoYAMtyd09q3ToFUUQI+sLdj6jPn83Liox+h9fOxungeuMTeTls
4ZlCl2C/bfNHpNtsZsFN3kHCMpIK0lRfdFm/9XfCthS8uzVIvA5palPM86Xddwtn
BZ86j6Z1UK926p4h3cInImWZ+JkLpvyVYHaqOjtLPdkhHg42fCJ9D/YqZy8/Nmvy
c5AIjcvX212uGfTLOBXv2UGizpiLZ3DEJgGOaSjR0Oth8Y4XXxaRmk16cBkc5T5Z
F2ldXIxgWCz3/yLKA/gf9Jv5Zcd0U4484P74W2cbCIZDgrbrYp43RU6jwLQPPK4Q
E4vnMEBjhgGN5Nh1HjAvef9R8kNTHr5DozMq+6A2lH3pYgLJ1Kn6itRBNCNToX+0
1FOfqvKeP1bpRUJ2b4mmSJTGsqRQN77fp2f2AeMjEyWMgboL1anLD165zQ001Auy
OK05OrmxCGlaJ3IUWxwK/UCDts2u6QgSFz6V0cvcpf1Fc1LLBtrFHNIh8FEH4sA3
0HJcMWnex5MFr2xJimrV78xYheLeNcs4vAombT5a7ULxap8bth8vpCtacM9n6OLR
5amIOm0hk56aelPgLRTPz8JwtqL8GYZxYHvQbewG/QtMJhmCRvhTxAa/YQWkmKdX
kDxjT2MxyhaP6So1WDrl+Y0Ws27fHhAEkcMDzwEwaNp0ZaKFmZ5+pUF2kISvufbC
0sS9Bc2GIP2AnLb7KhIOGZcPgKH3JObaSvoqeVWXXEUhgzGilmknsDNs2ge/n/9v
pHTei/6vXCU44vwtbMPtxVNb4wf6ALj4a4CanSSRlimGV6R6qQMC+cxgphUJvz7a
fG8QDgqDJWCyhsPX/cakYs9TxsolPxjhOZ+BSkhc/sKWwLjUeI3P8UOGSdaCoIB5
WJoa8KyYjvcuTJ7tyslls80h2njOJ3Ifx4WWQAjZ7toPNU7H3wkpPutHM0fbPDrx
GCbPmWN3TPvwmNc4HwBLtLwCnHOSJ9yR427jfx3KQSRdh4adHQdDf1xp4V6YcPAM
vjXErenErup5BjGsIkcCB7oSKpvsR2/FQ4k+ukdC8ZHfDC8z/KTH0deYAU9M4bPG
xG9rX9JbIfCnJeDtOnCyYgoHVxoXOH0WNT794t+wZ7iWPkzgZjKRmgrVSRofe0HG
X4dJm8qY5ZKOS7GuvIhNXQvWghQKIQNHRl/lkDWXo7coTLPT+4Pdn3GGi8bts5dd
g9npLbK1iRN1NO3UTXRLGh1nLS20aJ17hidI7+xj1CXZ2GvThQzS+fSBPY1bvBBR
/7uL6vXS0+2vGzM4Cad1VKxMn7pNz3HcvssRzdGe8W4EFSSTfWWTsLUZ5bCjwuMe
oAtdZpLKqqRf8qukhPZe678Ei0a7Y3F+xAJ97/FcvoxqXO8DwxtDN1GsASO1vuJH
EKou8/bSTb/SpfjZbJwKe5raQ8Y54TORax91bDK3/v5jX0ljG7S6WgcwaVV2oN/2
6SNYgyGFaKSJnaiTMaO+Nk+KOjSYEzlJb/d3Qfm2QuRurhFPjOLKDTQfG7YrxnWE
CttKkDyzSl9Bc57RYAVTonXGYUnkUjaYDvGjWEA2pYcE6T6B6C42/LDhs2zvuucn
irz81doaj9XT/ZsuwwKz/7UuJruNBcJATLdp4C4IsWXvyzqSnpyJ8Y5OP/eqLAtb
VddiwxBSytCljHNzKBBCDOW6GrhjkUn8yL8LN1BRaYm9H1POa03gTyJpE9TKap3S
6sqbCQPPp9nMGnjSWuKoZ95Q+yJGlKalR2dUmtDkJVsJ814CWD/2IZ7oqW0Ho8nU
aFET+aolCE01a7K4eaGQ96hCM2JN2EFrMh2pYDbD0RjbC0D9S4aMjjg+4dRQSaFp
NGYmRQLAtC/2I26AQvl0MDiL9Lx6Z21cBclI7ZlpG1EVL7dWGHnhf6Po6nhauxzJ
8Y1cHhABmLpPo99NX9B/QLZHVhc+MF5QN3V2QMkDU6Crl+IQu9kJEUu+kvUUq9At
L1jedoAdk9ARZAOOaZs+3/u7Yw4aZWG/U7WVckPn9ySl5c4+ru7O94Hx9gLxFH5S
ymIcm1xZhVhA1C+iK6N/BoCxp3ukliezHXr+bGCEjzl8Oj9zBDy9F9o9FNdviMzW
2D1srE7Lvey5OiqAWnuGhtiy7qZaMcO2dFjbX5353/D1trIOSLaU9KetaxMuR3Ie
fCFsf0AbnS5S00krrqZOiaIzHBUYb0FwJa402FEf4+NTo1f/RRLZbnmCFG5EKBZJ
04x5yX3h8uYLAxwqnqv9N8vJwVQlwBH9poiLmoRLbA1pDoE4u7hbH+uxbKXUGZKC
jG2iseVT0bXoQ8mHkpWj4886LJF7t2Y/ob+QJPLD08+P9t9XhSQCnupXF2x/dNxk
PfhfTYiFalxj/yEIXC5fJBCFgCO1lfDFt0faoU1B5RTDWpRNnuZNH/zR7AZffTo2
Ob4og0eBZjQgl57yh1Ld4oQox1MRswrJa5uaP9XtPeAuqOzKZsn9D4z0SbPn+05w
9GCDG1Zl+l6qbtuTgZ2bSCk0oWD3HdNjmeBhyhJoOWPAGzyt3nFug//tF2pGMkQ4
PLjwmazguOFgwGnc156jvrt5YUPZCfq1/1KUYfq4YaL7/lLDO5HaxC9zTyzUUSgc
tcPfy257+djLvVz1WI21/IB2lPkwu0QuS57vU6uubxuDdA0oMRgeDSTOgF2XxpH3
NbFOQ0a9me9LXgwoJJIdLJIRIM20Iyge6zAG3fxPDz9cONmMHJbdR6LfrEDGA34B
zToG9ehoHdfWmpjKtNpjGKteV/Y9mA8dMHav3peNXwGgWL6CP/pOFwatS8bgp8GP
8qE56dJZs6D5YSiqf5T/msiLdGZiJjYjgzhD2HZ9je6Gj3roJA6x+VHPEB0jhlCl
RUIRBLwFl3BicjlUfripX4DP5AIA1MnKAYDRCnWgJuaAA9dYsIFCCcJ3JG9Zvdea
oLn1XG4cX9Z16fxt+Vg5N/E1oZW9EWVtL0gwSFwohCJjh/ykeY83Q79ca8XZeZwG
AVDhxrL4r75zmterDlsfJNpt/A51OJ1NDIF3am1J1L+2K05fTGeumutzVyj/tVol
fXzDys0FN6Wi6RMmU/2ZtKPHMmzVr2xPtWaJBJWQ4ftv1bDqGrQLw/5rV8h0UJUP
nktrdDuT1bXp7WVbxBunT1eia1i5Fp/xJ2Bvv+7ADm5V4IF0J9Fm7LcnnIQdxK6p
egGRpEZFod/jmVifpKPnM+YlDCwD0nhekEsDzuA8elm9Nlzxc60eS3IkakBGpyNC
167knnnaaOW6YBh2SMYHoydyHK7E4/lm3XnN6savYk0d06HzqFKs7KeVaKweAzyE
oIY1P7sZs4fqdOSR1fML/cqFjAjSknCLglm8eJv6WMZ9EkM+R/9rK4cQXyQ02QZi
TNUL4Y8E09lLm28MQShofmKxBGnsVMXlwSI4yU9Uh88TThspbUhEkqxHlgD+8juJ
Zi76wY9hd7wiTFr4tNjUvan8GardkY+T7aOqrr/PTnkWeiprge4TkgW6N//92LtF
upCXIGKlRQuJTyyGwzVKYYpij1pKXdjlmkEZ3rUkAvQnf98eEo0Ce13Jvo6sF+VB
Dfm57mWQfKuXwJGhHYLcfWcSOD6ECvUp7wumQ8EYvKDl30j7ajRlfJ4bbhf9/Z5T
f5uFmetnmJQG25PIJb7vaxZRe3XbMDC2zZJRoYJee5PNLza1+Yobn2sgk8OVdn4F
H6CgzZjTwUtJvycECGc8QWimhtaIHXnP+Zhl22D0pi44HgGJ29tYFtYRYQwU45y9
at233YpwdntzB/io1hBb19vz4uhfIvqbr97s/C1mid6Eqh16lxLw6n0jbW8/r7ig
vGRoAzivjl+6hXhufZMn9npsYSTuHxnBAEp2tuU1WH9EdrvH07bXF4mDPcFWMBiG
Pl/XgI6RRJT8lNZ+ZCC84+7sGtZZDiWFElgKfvw8P4hAjCU9mxkZhK2jlKmK40zV
+YNSC3TakF7byLy4eq9VebqeUevoFtiukdYXRJ6WZxESfLl0E5wdMXAdcEo7605+
jr3w3vnwqn/gAEgtl9E4YSK7QUzSAY0C2bLMdhMRpP38+6bsgXPFhsBSRLj3XP0J
c3iSGigOIOocNUSxzL8d8b6PPPgNxzGhfekdEJePvSjAJxvEmvdER4XD9mn3Cn8Y
8pAgugfoBA0Y1xdgDTN1sjNXUpgGlyG8fr23b7YM/CvHwy+L2m+bNlRL8n2PwHHk
KvllZwRKoIZoWuIISI+aNTwTcDOiim9dYLJiFsG5fO0BHrE0YiWlm9zNh/oD+q/R
C6B41i9AAgvGckx0B166oJ1aWQ9lTuXMNdGwpt2pcGFPAgFnY9GtCGBQ2EcxO4RF
sdYsDNDWXdexX/ws5y7BlT1S8AYB1FBBg2/mT9Cl5Msnq9DvQWQ6MCOCnwkEETdf
ZTRD+bZOHB3PWkazLwSH+5DqfL7oZTtd6Kz18EzfqtR8tExVn0wb+m4Kn58lU0W4
NfUHDNLNLaT3+nTITSgVsy6rq58zQ/vFFQBu3MMdA+8zNER6KvrL59DI9CcJQOMI
pYRRXeCi/IZlO3yej34V7UZhleX95qv3KcFWy9240Zt1gnIV221NC/ZiW/K/Zd57
08bzaasAZ0iqJhdR4sKhaGwd0fuw5Wli/BRfsUH4i9UTLgBSQAY5aiej9xiynyfG
sW/pXXM428QuRcP3gtHyYHIdhCTBiB0OsX47TG2D0m5uzyIkE18lsqRQdjaInGfm
EXaqGjsw9H5QALYEORAxSv560Hhmf6lkXixNXglZf6aj8pRCN1uAJlvSxgJFMf76
PpWamR8LiNbiOqSLLViR23RSfJbxBnXF1hchOOJTXBcO62DApKrUQbQjWDJCbf8s
Zd8jLVb5fRckfWaLvB6FwgS22xzHIxcJLx1IU+pIFcnc7e0/LgSd0LB2KMKWjWzH
OygyCm7TJDpqqQietcd9cGlK1igb7FvdsHZlQ6soQVI9647mtWRcDjju4Z4CaDl6
+N71yVCt+hfoCEvxv3QGYv5ogE42C4Ml979NM0nskvzURzQKKo3QvYwDaDrW/odb
e/P83GEu0qEiDcjMgAzxhEybcFCtThWqGwAlp1xmoBj7lZ70w7SoWUI4AZOiuSkr
9w3uaZMmtaupxR+O2+/p47BX+zmWtsKr//vKQLbLJgdA7VaPC4ZeK51X8tASrdZm
d6bhvNNdqBxNXb0119AujhFPEQYrgEPdqLQ4YoFAv/KsoRVtAGnZBFLva78VJpoI
mPNdNFK3QH3YKHA85kEi6W4oqfpI27VJbYx6BxyoELe2C168qM65I0za1XEX39dO
Rc0KHLQJX20M2/ucCizZ3j1tPIw9wQtVjH67Ktcki8EEBkkrOmYQujVjUIcj2Mzd
NEw+5N63FCHjYIqvwXoLVMCyC7k325h06AeGi8xEk4Hyvoktkt8GP81ueH4Iqy8+
6yyBXR3Mgjkjs7/CjGpvtGhjATWPzNfR+irP9pSWdC+ciOY94ERrJnUjirazw1Kq
OYSM8aTpt4BIX32+6V0SwZR8Yi6uI0rNrOSbaOuf8camaQbpVS2fJuaCcIctSbkP
W/NcUz1eHy2/nvRqdmOsaZkiqDhO9HrURZi8MWSGz+6JQLuD/XQy3jkhiTRm/Vl1
iQYyleIyewpBgnTedmBNodSzcLLLGINWEp87rOCElFo1Xn5vhJj7U8i45aXjTsSi
LNHKctDlsW3hdHcHnnMgdD0fCIohWgMXh21RhUEiYzR0enVTEk06DPSEp2YZdPJ9
Uc+DSsP0ovPEaw8vjODpWJpZ9GrxV02fiCXJu9v55LKW8pNsOcCXj3EoL27Ht7au
UsfPhjHc+f4yOuorgsm5cSfktj49AH3xrzaI/vu7wmYhcz8dDbBSKCBMKGgqcTty
N00tT7ftY/27xKuYQgZvuC2CxuO/n+ozWaczwn7dIoe6U6cmneFdTzTZQ09IZDM/
KmDoygTVh4zEydYWCvzoxIzypRS3GHzURx+99g81jf3Iva8aTexxy0y+593O4Ldm
dp0SdUM61DlVe4N/SqAmRYCeccNfVSkgcE+tpUct+jEZ39Nn1at2dluXMYs9+Gdi
qf0nK+EHlFpEmB4V24Du1iV15BtWRJy8f9ui7vRl15Ta20Ug/Ntvyyk1QC9LQp7D
YNXaj08W+4eKYu+5OTo1DWkHjLZHj27H6GLM/6MFwSig4gVOumr70JhjNgmZvefm
IqjTcsiM3i8UMhjkBhGTcqqS5apKVrbCuzdSbnienu+ffvdQgM4nYM8r/JZqjxqF
YgllVJNkTjhwqypaUCUItP2cEwBxD6+lTyuJ3L0yfkjWot0iiorAlNHaFw3eCt8O
Tv/PjOwRDGH5oslYCl+VA+iXjjwqndoONzLRmV/vuwAUHLXVCH9XUv0g01B+V6GL
bery6U0vSRrL2p+8I+T5umxumpePbsEcIKspQKQi/n3ifGkW6pZg2Ch6PILq8ebr
CfQJLRwuruAINpvi1XOIo45JpZEdud3Tae5IBFoKTw5mG+xWt13zF4IUqHAesQQQ
kHDxcVcsFia43uNiv/8fTXecZ42gsbq1/Dg77QSMtt0/TfGsDv/4n/D/tZC/N29G
1y1lOwVdNij6hA0e8TQvJ3DgahYle8AUpq/Xn/ayUPcUmm1vNDjjkDzBFMNPMdRw
PSmAijGrsLF6nCPUGLa8auhQxPMRN433SCzNzcm9qbddhebIdv4AEAszOhKO6KrF
Bc47g7hK4M8pddb2cXgHfDCuOPBiinsZD/3JdMNls8028EqRgbE4RpHfxlxnhpgM
5UxTDSPDUJ96kPcVJGYRZDS/WE7eEEz7xLEvphVjsGRY2nYIbfxc17PTvgRORG1o
tar39ziTnLBF9Fr7LtBPVfZfMg8ChkO8JPGkS2hZf1NmnLNiub2uQLG7qt9fWE9y
Lvc9bi46TxJfTcItw8oigwUtumSrLZxFIjbvhsLrZr6QH6lF34s8vKl8cW80z9Yc
99RbHhjnu8fgWY4mcZxuFaiRoUg0D9MGnmJsx1P27ckSN0BQdxIuHQWPIGbTOOeg
ZkHnsP1PHgOeDFXy5TTyaz/Ee65KDxX3+44dFZHjpOJZHxuO0RF/7+d3Uup8QoCy
S7EosSdoSTZGDqIbo7dct+jQ3KsdFVW6JcctzN7Gsmxnwlh9qrritIQI8+NVXxS8
pBqUhrkd+whLFs2tZUzKoU+dYghswu02jA7BuaZzhFMBkJdg1SjLbHHqdSR2Kvzw
HMS5gH600FG68RZ4MxzbOQ+alei9cbGUX5n6TNYe7zWSWkLL5eqK6yAJZAaY4DsA
jBK/ysXgLLD7LWdGL8eVewDtntRqjI8+xi5rkqbXDVLnzAIFBa5kuAEmATZY1XfC
ZHMqO3xrQpKi3QPyhpDrEBQeCaA3eMJ+FDShES9BjQN/iClTI/bkXJpz4W5eIoxP
4DEy7yhRDZFbYF06QFkms8sRbZk5JNBCIkpgzXlgOR5vDM6yYmVaraEb+b1kfDai
YwQ6WnBn4PItpG6jEzEG18IGzIZfaQSMJsDm/A1D9ADl554MzuExQ1Vp/WC2Ko2M
AHfto8Lqts5qLjviULnSOOWFaO8g446p3aWCummbJc7uUufOLtIlh0yj43vieq8i
0xqeAXFRy/uyJol9v7bWn5sy2iAEmzO9ZwycGmse/LLfVyxOAAnDVm647fGN9Cio
oe6ZfGuzTBActSjAQLuKQVM+vWjDWLfi46IFyAjPeeNnPmfSB1mj1bbsW5nPk4uJ
WJp1QfXqBGs6yPTq/W/vjd9EUlB38n87zkT+73VY9kLVjAEO6/Su1fnvJPFVcJSi
pi81FiW20T416EY8UgdceK9QPWsgeJxT+PjGbAE07C5GUuGEWCT6xEfX2nZK5JmL
ObBLomPb1hQGeJISLtyQmoPUTcbSugEsFtIPN1mfqYh4HhrXt9MT3dRlLzfljEjv
kCiAmm8yuAyi4ESfLE/cfCyzUlF/x9Yeq5wIMVRVB5C0bMP9pqpYAsCIJc5+oKIb
ZtTeqdf8CKWc1ryxgvHjBCRgTehysn4gVjzv5AaITHMuh6xYxSG0UrbPl5s+Ntar
Cj2Li9LXi6KYhP9F7eWVcxuHW5jJPkjZgTshbrnxGb6YwZzPTdDia7lefjVTpjYK
qNEt5SURfD/8t/MF4WDct27cx5BnNzJeusgWmR1gdy4V1tjrIp2UUImAf/RrA0TA
Vw9rRwLcaiAqVT1mvZeSWNGApeqF57wGDklCK2N8WsnVsrnW7q+L2eJ6J6+b4z1S
tQ2tarVNnwtzArqRpP9gLOeJF5bl2IP484foKW9C+nUefwshB6vPJCJ0DCHh7tw7
Y024X8L6fTOn7EXynPBKKWQaYfmS1RDtbWN5DalDpJq6GVz5fNcNpJ2eI7ikgMp2
PORlLvW7ft3JJ1thhKbku6VB+9WRC4MT6HeHJCiBoCmdwxX+KKbh5gp8pJHVLTVW
vlfmyhiIrVrr6OQ19aKN9RMiX+csBq6XeSpo7YIIULGZC0aeytLFs+jHuan+bXtK
fyhEE7o4jaEOExCowtYdcXR9DZavyOAyI0HBv5GsazLlQf0aghcSw2wr2csGIiXx
0Qug0cspya0bKSVg5CQmcUUMLrjmGCVd47T+7eR44iPCgI8/o6lVp0NqA/WCb+rL
ReTGHXtgYlUagobZsT6+Fo9TEDwWygJUPVe8yG7PzXQb0Stzncrs1zMd6EHTCzo/
Gloq7HRF3t6jFRt+LzovlUGsRYADX8Hc3LGB+OM8CYZNYAJ5p9kpLdXPv9aOe1vv
/vaS65rmZFWPygEvYuSuC73/ZUZdkxnIMF15jyN54HCgPXcREJ2wE7qiFxzPBGVt
EaAYjqqB++nZmCJLS7zScyV4yYJ/L6dCtLGRxCONEId/0gZI5vNAgX1Oud/rZdtQ
TXrkoN92V/+tDZlLPc70IBLT7ma17CPNydg0OpJLl25JCgXigLvzDbbWOqKHsU+O
SDp2zuLLxZIFUTM72/VtMqSD45rQnmESr9/lTUgYp4rPFXX88stnh01iN2+LxiUT
JMrfNJJWKXaXHpPFFNg0lqkfEgMxqnTp/aSk5QaHQGPvHJsnwixs+I1iBDRa5F2j
k6WOF6lSanzDxsc3KMGQJyzoyAsR+bJr1qxAcr0UjUN9uDR8jVqZ7O/3yK1gMly5
nfwdO0/3OnTit2QTba3jxs3teS5/EyIMVOSlYtL5T0YWmcXotToZ7yIz+0juOdIU
pC4w/kGZ3uD9N/jG81tC5iI8dz4X5r4e0TIktKUdYbqQhHITx6KoGvMWURZWjE5W
75fMaNsFrgT91lc1Vg6NwPqwu+tzjEra13x3GoYzmZEsK99fAFrgbqVBFi55xQIr
+PpSpwbNAmDjIXTjaIbBzsQewOWYp7f5belaGNo/hJysFeGD+7pBQm+ramYypIJu
9RkeJ7WCHWUoaKYlEhDRHWRtrhW7/oqdOCQwJGvLrHXhC7F0plCVXVivIbIUbATt
RgScmDP2BgcjKs8rfCB7fNQ8W6bv/DKrXlEdEWQeU12Man4ExKvpugF1jxlC1huD
qKVSun2MggGA/isFWBzxNeOLQfDHg1nj9ATjIWMvcAv6MW6lU6D0Pmu9X9UZoIoJ
Yn2zU+Etq/PpQMPswS8wSC6zG14qyjFrHqTW0ewXulVbKdAnbiMwIynRUFr36Hhe
J8or8ATzhENysx2KzxYwOcAifJaHeAzCAoP+1j1MR0hlrvanlenWJXUQ4GbaYVfp
yTsAGUa/QF3ObVQHfAnce+cQcXJUZ4HxaUTyVlT3W8MTGEZvXGlDzkNwEHaQEGby
h+4NLt2/S402fIiHP5RTcIqW+3hRNx6Ar6TFzpN/AmtpKckPCUsDeVMmhFrdWZCa
yO/SzTMIAKQ19eZyz4LQpPCCOzp8Y/xsnmyMvq1hvLtsaKVu7KrdaCGNtpD3ex+u
yl4qHuy8SwV87WQAzfJMRC5rXjEgfBmOSAxUj+GeaW6paMM0jstMAQ0tOA3ThGAn
6LlBtJpWVBUfdtuK9Yg2UDrDF99JJTFSUa/8JQ1LIZfGM9E2AOLpmewP5umbaqQJ
FmHHo9u6g1CHEXBAtI5pnxDuiPUE2fvmYMWiVOk1STmzlcDrxt3lNdIFJP7eRMRq
CeKE52kteid+SLlph1SFnmDZKFvwjp93gK1bbgyDKDFIjgDAY+HjZPqy0Jl8wS8O
ueSMwtq8/RFHmzRMZULJX72OdOBH+qOmTSW+I3WGfMrVuZEUKHTdxSL45mYtyY+d
`pragma protect end_protected
