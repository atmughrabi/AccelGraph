// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e76WAvaOp2iX1DDjyzbpAnDITL4CG+PrMftK6uuWSlQSmtGFxkCnQDt5h/WJnXh7
ElaQ7gU8eODMULXAn1OwQsrN2Z2GD5CI24yetm7t/pvi6j4X+k6cc8BjVwKYvOpn
eSkuA+LthjkaWC/eEVWOeVi7n0h38xxjhnMsMEr/mE4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 132992)
s6Jk4PA/0+Z4eEoS1jTgsN4xuosy5Tk7aFccDzboXgfFgehAC0GeJfp8SI4OlWN3
9DSCBuZhYtnrGf+B0STCL0p0DhuHVNdh7GwLNbhClZPbTJXRf/ZZJDjfQXuPObH4
BK1AI3ks5jywsscb/xlcXmkscLfdz9VkzfzY4woxROQz+KGZs7feVUsOsq8U24eP
QAscI4cO7SScSj2lekAFd47GgGeIF9Pzfg9ZexFXZBRK1i49GOq5KFALIzi3B1+6
ogaNHw4CJknYYaTYCrAMsi8v9FHp9w4gLvhnsa4nzVP6B5/u7qOrnoLK2YRt7Ieg
Y5/hmSg2wh9KUmHGDv82Q/H5HC53jlYYZ0XHi2oIaSPFcghZwIZxI1ArrsmgbM6S
Ko/PuMM/Tcw8EKS6YeuIJdA9bAUkYCl3wG+S56Aj+l94kachX0B5BVwezOzU0JHK
+TJ10fZpT69bighyS3vgh7s7maP1cgkXAl3uJJwGOEe0X/bW09eziFUt+gRfNloy
6lrKceD9kuJuQer+ktf1jMI0CY8dNRO248qgqtSidDZJ8wouopuRMYejwMGSsTIY
CCF0o6JPtmqAhfQrJe+p4KtgxFbBsH/gHdqjp9lu1+I9LY4yi/cDcq1TRuj5/Wkc
2Ts3v9cDfnQnXX6STdx6yrTA23cHydLbcPZIPFaKLslS/7bJgTmJXjgqIuFpjcjM
x1qGNRdtw1M5cmcaw1ez+rj9jWpLYlxHqfxX4BH7AHY92Gz17uSXIT9ZaVvzo0vZ
kRgKxAdULOTRSxIHOMawWw3JSlGTDrobkNxYsgKplsRzLyBf76wgqYqTep796hJp
ks/1Yw6Q6BsXCXrUSCLe6gmRShoXM0QB67Cmt0VqDzfO8JDmASIBIiw3dz5im42I
sm0nupLIGPi6rsoDTzi8yf84INho2LTEyp0vj/7isrJkQcJ1ojnPtlwqS/JZsqV2
hzp9tJ3q3etKdCeSgG+VB601FMnHKPaIcElYetmBZxnrtWYMRjgVOiduJh6sYMJT
n6Dgl+dZbNwd29ZZ+AH/6XeG3OgH2F4tvc5zaQ7cvo8gguS1gVVaMMylkVMPz4uX
z5famH81yNvNas9WcLWMncNUprqympO/h+WdPG4w+EzKqYL38M2JfbmJHD1IhSK/
hm1T2Xn3LXn5ph8xnfKTtNxY/Wq4AZGXU3couweCtJ9ukB1/z3ntUeZ0pul3ezWd
StmfbZwq6TFmcNWNYB6AbhaiGYJ8ed7+PnO/RmIBdJE9tanNG8VkQl8J+dCWp7Bt
sTeHcHBJQzrbwcRuRyw6+cERMPJurfkFi6061fQjGB6pouKvC7TJVP1aEqBkoaG4
2+bgBmyHo8YQi2WiHD/dDwOW7cL2Ps0BsLTp+ayW3yFOKkjJLCtCeO18BpLiG8Mm
XnlLCP3RsgRM0M20XNpDcLMME9g8VeJin8+KqwiWI915BRwrUgr7+aOv2M1kVWJo
kHuaUumcc8ao/l/wIoy9AOPrIC88BOrLdNDG3j3QA4k0WKDX8ktpZHnyP5bfWzre
qxrSbChRRvasN1oIDCU/GO44TY/DeyFdDUs1U6AXEpDXNses7diXRWbHnLvWJYrj
v5eD0GMV2Hnnkjrzm2NOz4CDXj8Oz5dqQRVOdxI+NT8vNLi7FWTCBsJ1yMpRvT4/
YUn17ffam7pnTmhelHKhL/abY2aT4sQr06Khv5o/r1dINO2k/1PdTy9RLXgj5KkY
dtbBdlrZbJ1DpbA73qvaDU/ZfQ1FY5rtbojU/IT8adbnyjLJn9iRJuH2RyEn0RZr
2u/GZATs0/Jf4z+93ZI0Csqqr7yfEm3v3SobP4KkLq0K2iuE9Ydk596/yT41qaep
ZAM6Dh/n/5ebgTfuyEMdoKW720dVom717svkmP0ZMt2b0vZwQeXHF8lUddZXyV5o
ykAvyBIM4bwBVh76Xq/TjXOWBy9L0GZHt3xXqv8Hg/yAIEWGS1O+i+vBuhdwPlzD
Qd/eIMe+0AODN2ye3tp4GpJG4o2ZCk46XJaEQgnHr6J2fxH+8r4LOUx0zr3PDyP1
TvQCei4pwcdxdsHQT0tlMoEqk8zxF7cX1kFeUUmjPHe8U3sdLZzGtz6PTjxB1Qtc
N1+rvgYIme/ioKs2Ofx0mgiPhd3jV0J/X5uVibf5G+mvjFk6ygq2COF5OK11RGB5
74F9/81IEMxw97OpBOp+SdO2VNHKTjEPhouSAZ3zDb3z8AQtfu6OhJ/te+k66osS
G9vbzgvg6z1kW+ZNYvxPrXQbjP0b8NObhxt4Rh3UjHNjtjeFWTgJxfg6A66D9dbC
B98TEGwOqrE3SMavwN6GW3Tueq1Dq6f8MuQKO81wuJfkE9QmVyyndCd9Tlwh12PB
v1YALSF0HqxE5X5Y7f0twrCXECdkqZGRwWTGN4U18k7/PvBGJdkPCNBus+EqSywv
BSCt8NQxiJ4B0Zt8dYepCib8ZvuQGlf5nSLv3YT0QtQ38X/EtJ3sFLyI2Lap09u6
A/nnz4vUrDoOajHoze6d+upwowOyM9oikP3z5YD4eRL+0H0nNzdbJ182khi4gC8D
7WwJUpl1Nr47MyQAPBsJ6EWeXDA/EgCK/sokKZCjldZfhGfcutfcHxnFRRpC7D2/
oakP+uvwqyOjThiDpNVASJmG/1xY5Luv2gX3Bf1RLmWrSahyzZS0Aaw6PyNNT5jg
ajeVUrOmpIWP+p2YwFJHVGcLcFFeiBxTjiFg1+GEY2VQSyP5AGmxFT+FIPw54lxm
7LnSAxmvSZDeBrcIDjrWaRFA82aC98s3J41cd3bokJG779w+tHM6CYiMrlYcw4zh
zEfxyVB/f+rlsuDs0Zbem5xcS5BU8VAMHkKxkIFt2x/BYlMJ76pqihLqG0yJbR/L
zear5OvLhIXyrfuSPiDnSyj0hwmWgW9NiBHmPjO/xi+fCOZOH0xsAj57l5DrRM5c
YukMpviAtA8nUYGU3RLogY6fhGklGSvhY+3bhuLg5bFaAS7wN5sF4II4f0isGODR
PORtJG626QOvq6DFEGyXy0M67rUT7FRxJaSLxyOiANjf2Epk3K9dIhD2Y3thqYY+
D58msoP4rT5Cr8YqijLZNwswX0TnNGWR3MEXn+gbOxrJr5Y5mWYo7z9q7CsU8iKC
HJaf/A8vdpamvK37iHP3xR+aCrJ/Fb688qhZo+v8dUEO4M4FhjS9eowNkv8ukfX8
Jf/unNlAj687DP44wgqtaQ4sypg83rF4/8daQJdSsa00tmd+t7lUZZrE8NM73++E
Pd9TqBdJAnRc0WeTwLOEpXu8WgPZX8+yZvTGhA5kjqxdVjRNvVNvnxj15Ti1rD6c
9mLvwIUY2c0FnxUvMXjvw4gpbppwzrKBtmfAkTSPBfhklHZYxtONC5R4xNQa065n
rurQPOP7igmV83aclP1z8JtcBD/u+uY4saAlHmkFGzxQkMzLYbYbXGCzE5LUB4qT
ElzBtDAxSqyaXWxznp9HzhBI8mYMs/GILTFdVqA9lkc9U2EHJTFVzJNB/gVnUA8p
9jANP9Ncd3VJUpKyUYW3JSC5StntaPXZPRBM04zedwHb7Tf8FFbTL+5leznmBgeL
3tlLBY0Sto/rWJPW8O9SmG3hF3dCKXMKlaM+s3Kb3aI7D93yMjell++PYmjPHfp0
lnMiTlfLAmEKzzDk9THHAxHwO8y0esBhV/Qjwtxh0v0bTu7LvGEWtBbv0r+ms+hs
XxcZ+CGfyIIwJz/giyUbzk5Z68a9hDztiK8xMm1GGhNsT1+3siaI96TTMWJhu4Wq
bMpQvxSA3UdIcQ+GE27BiGHc9465XcnpOq2EYyv9QyN4IYffztCpTm0KKNytwqHV
DJHGBKAC9VpIEKPplur2t1fD4buGIVN8v2uVkgOSDp20Mlbrgoqc8MW6DiiPwDzD
rvtV6ZasVUcRJT324UCn+GSzjxpYkSDL6sHGo4Pi5ueR/e7omU4uaE0MCWyXqiky
6VWIMqI78/mQu6D47ASYXTj/18dBGhuq8tw0/76Xr/0kWC3XcKs/icOcwaC+FS36
eL2DOg9/bbBp7kFWvUw1f8wJh7wXq2lVqUbuxL3HPVA6pJwpb9eanr/NAh9nJwGq
7hPQ3uKc8OOzaAWi53lZpRlOn2kgoTRloBdEpeNqEZ4ch3zDSO21kuQOZf0JT3VG
1X5rKqOBN9CPD//tdTTpn+3QDkSVeotwzx6DbtczWIfrqYNkUV0V9cPHDbJ7lMLR
DwqTgmQfgeQQDf+6Yu/ujTYaR4LlzSHNOb8R6q5urv7gyhtDR7JMkpDNG+JFPq5E
Yxt2b/ycFqK9nIDWfFCu17HEZGolVAlHQK37YFVZA/GvEeJwhfZGmwfVjnD9moeb
TVI9z+qoDVMuqFjUy+4sFustp5LACq1n7Bj0Q8DPzwfvFt+K5lf9WDuBJiwIG1Mw
lZbXwHTLXmTZUH08LhjFd9QNQtdd8R8s06CTXoBOO8ri3CxsrZKqw5cbyO+6GMue
YMqvGD7HuZsfJBUZ3M8ci717pxJ9CCGX/nFHvvgdV+Litj5u6rDX778tnNV5UZ+5
VrB/49yw2oNzkxzLiYaRsHkARj8eVdYLRW+0FzOCvaF9FUISckW+f9CZY9E+LPCR
eZnwJm4LM8KHDpQBSPf0kJBl1DmGY85mdZym3I7laQgr5mpasNM3SgD+Naq8YNzm
uz55FWQ/H5Nnjz0TBaaEoCDHCjqERR+VcYXYK1Q/p0yP2rY5x+gXCVfHWKkoYvbN
0wWm2aIAwN0WPXhho7klBpONdNIMkVAg4HkUoUYlqBWdWwN86xtf+iczkqcX/E7V
u1/YkvMlHqvmsc7dY6GPAz9rfSso5guAt9vyz8pBheHGwtYdK4KKk0OGn7eHyM6P
IGqob+wFoKnOzIngXIhn39LyBiQpnthiZFKszOaZ5H7kqjcdpifOTJuNZ06zVavF
5UragQxwz97Wy0KaEr02VY0gMQ2q4JsnTFuH2fOKbKH/kQ/uKFZTfklmxjOk7ady
f7RRd18WT2+MS64anEjr3v1AbHvUV4y2yMaQ6yPDOgA5L2MZfWBEqeGB/B6SgRx4
I1TG7W64zU0YyRFBu0kIY+kq9j2+HwT3HaMWzUT1W7erhC5edX+aFU/hnHOtGj21
bOILCAWoo5i4DZkc+4/tdSsoPqoJbBn0ArmcPDzMwFQCcO550SNJvD7QumIsdHh6
lDOmLvAFUDpO97JFGk7CryfWbgD1n7JeBa6TbWxAZXw4AGlLYgJzH8BZsJYvdim5
vxFxRuFmph7KfQLy5vw18kjSUU83xsJXlNmbWaBPf95xsYk4D7+MPNlblGxruf46
RnkQjFY75ox5TLNJYDIunFlD7hw84bQET9UmJ2gBv18HsM+2Y8s3yp098yQzznwc
JFfIgwnVkrMUFDotxHO+CgywGGeqjACZ92pc44vB6ce2Uwg7CRoGZ1+CzyDUc5e1
MiS/iTZ7V+i4UYKhww+CdxVPyEDoVBDJDKHTa9KqgOMTdgwEqOmojlGSwdIh8Rmh
+fpVCOspz8JLvI8GOeqOmLyJI7XSxUv0UvculqDo9hUCEmrOODdjYu/a7NnmvvM5
wuDTUO78/sIfI/mo8uWcWtB1mmMvJhbU86gR0MiODvOF1UtDrHycP7hHrtDCUulF
h0qO65NxiQbfZRsj+SgMUuNWTCxmu+1ze576bW38spVKTKvwugHRUJwcOM8SXQiX
086ZpAFS/eAhyjcdDD6GwWAu4WlYCmKmA9e03D/YIT12He179zWWC7HRUBuc5BYC
+odobgK/SYmg4/3vDNInstOuLwptceH8VeFNfjyJt3Z7+cK55jF4hHRahV2t5sS8
krBEGvCZdfLml/6VwtihZ/GAHyh9ePHCBCuokBjIsgQ2gZwcsR/S/Sd5RXS7/rbC
AujAwE7EOA4QyMP9iQAWMpGJCMSCYl1EtsGmQ31t6AmtGaJD0bhVjRlqC6uLM0BX
gdW1y/EHW7YjG86nzxX9BGgzjmcbug0R1FZH72UU4E2z2Vh2gHF2H2nTyP/oaGdW
Ze+pE13cd1rV1Yb6003J9MHVsegQFc9O9ZiIXZrfGeO18z90FE/fhxHUd/wRI8fO
T8dt7ya9AedTt1OeVDR8FeIBikOSfkn/JYpoE6ge6It+EY/qzljMSRonQMurax+7
/64CQrvUzMjkmQacppWXIra0RrtYuQU5y3gRiIs7vRWVt1Yn57qVgmiRw66zJR9U
LRWZuKSHrq5bTRi8KM89wyWuUaWBiQRs79wv8DdVDPYbh6XLHdZNuE0YEgc+t6nd
uZ4ly4AcECMAqVWoU27B2setjSb8H2PPaIEVDV67SlFU1K0l9UMwG4FnSsaHPRQh
zF0YZyKLoMSinJSh0PoFJaGKe0+epeyGS3nCnB0hlrbvyAgGJixh7AGEC2MlUkBA
Q35hJTirUoGKjlZEsZefoFE+7dNIZFIXdrD/9c9zmS0VDBCDJoJ9xd9d1S8YIQi1
N1mt0N43v8CJjY1IexfUmOyHI78Lr0R2fraB4RHSQ3M92hXbcYBxKFJ2IRYy2lNl
1qDKdFezTRBB395egUz7jOOXRZEClHqrR10Ik3AezFJZ/rkzxweumfmd10EAplE1
u1JnLRZgrlA6sQ0aXrgODOPUDne458YAObT+FXYYqUlEa/90PO+Hw/RyqG0453zP
OmPgJoqlZb5G59wNEOdQuZ86pZ1GMTnu+1z/yp1JVSzWb3vVdj+ZeMI8qC+tmJ1X
DZrf/7x/Yd/8YpRkDs6pkltriS+hEBmf5gdRu9+M7dWMWYQwNfGzC4ZpkMZxG/17
Qj21m5Oi39Nv0Z9mBybyZYcuS5x0hInbxKWR8VfHhEo8KQ9UFpr9EpJbOel+ON8R
2ERvXd8fB45vFFDhpVraM8+clNv1ezuVFyGWsOdIw4o6O+68ZV3DmJy3xBziHjTU
3cckFeWXsLHEHLOzhrTKJw62hkvL4FrtNptMmKra5f1j0YRoHkwCeW7mPbK6ARfy
W0dVCjFntodSXYo/vLRtdZ6+qJvZtAV1MkYNklgLzkou8SHxeVa6dDkDV5h7GnMo
KMouTaqOhovaPSHdvOWJwNAT/+MlSUIkgxb9ZLdlKlN7Zw2JUotWpvH0FjY3f1Pi
mlFR38gcSZh8lapVXyt+1EtcyGvHb57C1SjMfdrhrS1ZBaAwOMzqM4TMe/SvRBWb
zrBeW2vkBBgzGokG4/rQNzarLPEg96VwN3BMZkLHdU1LkN+XPUflZDegmJZ+lThm
wdn0RQINVEwuwcyiZamUXFZrq6RKKW/wN/OiYQ2Qq4KDuAowDCKulIIegUYtUafY
kzblUZMvX+cKom3icllAmp9PdZRRF1h6SUBIXFiCM5AlQZsTC94VRQBfeNMYxKMy
BOQwPMQirWeuziZaQVV3fyb8qPOaIP4BHwkA4zcP/m1SgPUhieUodddR0KkcJrEC
AGULxO0RKHdCl09yq53mGZezDZ9w8yReQMBh0bkUbFC1Hd2u8gj8Gdf3zNu4o1DB
AmzZwypU/C1c2pfkO/vvcYOVOOgDuiMo7zWvdlgFV22mJQnIb2+uiHzVGXcKzJmo
3DnVj6QiDaYTbMcPE1nFrnNKYZuSOP6aen6lOf2B9bx3abu54hjCNUsbn72AQjcS
rgpFZq6cD4A46VajzVqt0/EXKLP+Pzl+DgjhL36oC+O4yiUyK04EMvo3aLBaXoZ+
hwWDb3VZHvML3jViFO4eX0eHD/jHCS9Osq8mRWb3U1OMd1ViJdg0h5lQ+vPq4E8K
bRzHJo8L9QhW23Y1rMIZmqmvhvnMfezW4OmUwedQryRlsrG0o2VNrW5DTPbyceI/
oX3Gc2kFdtnvJh733iOGolkYDG98uiSJETA8+Un22LQ2A3zKJEi094Hw7e6ppK/V
TTK+mlNaDCEq8jwLdfthdA95QYDNP7tPir5jEhCnVb6GV9nay0orSd8yFsLJNP6k
n3O/9x2/SE4NuvZ9QdiftZ99wli5G1T4ohmDofX8T4BeZ8e8WUuNOFUj1NalUYVV
Ubf7IVK9ebPdhzJRnrnS1LG17Ano2M9bfE6eO6ySFEOSfPwFMWg/ks4mFvTk+dgO
scZaijIc8VQWwyJAoX+K8B9sqN8y3DRAItyZNAY5Tje/i/2uQXGwCZLm8CSM2jGg
EePgni8IUwItHa/zkHubU0Iea6g11WPBBEYIOkHm3mEd7tRwY/2X5eeSdnPn7MfK
9EV8fPq9WFpoX0aUwZLAAAEqpj21NBc0/l6oDMYle0IIiIwSMuCGwKAe4NNcxNbs
ekr/2kM8EDySgaqJX8Qcxl6x9UZ0+/Coos4yOLUcc6zIh1hdaksV0WK033Cuzbs9
ApWXfHRgU0dI+dTYdEL91gLn+K/KyuejllosoNyvYLiio9QoceRusvSz8m4HUloJ
wIvuupiCOR9niU/p8N5DEXU9lxB+GMFPdHCtmEI9+GTXTLjxveDKdljZ6VL9buiD
Rqmir8pKnaCI/0zzoxM6r43Gs2qrP3K5zmnJJHF6Po3RRqP2Gp5vkg2FqWEEkrAd
NHTMxvPkPrnGiH5I4B1AFGG4rGk+hbdPryuV51E2k1VuzBBMpys8Al7i78LU8mpT
QAkACayUetg18RrgjjUmyyiUISJu+OjtUeYCVs5knGuGIyAX03pZd7ftwsSKJ0i4
7AbtpA5yHKgGwqzjlor4oAXGmQ+4A3ToPcgi6bAB7EMDFJMTqjdC8gIlQcPxp26l
oBcBV3oNahrL+bVMLFtvR2kt6TgA7kTTQF1e5Vwtb2hQUxExMzxh0Y2lxOrT9LM8
EJR7neP0ONTj/wasmddGFgOaXZUvmtNiOeTqRzlXKSPke8Oc25aPODlEsECtDwmt
9YoLN87B55mdK21GqAdylW6ibpQVyNsSJ6Uuky9EAMZCARM2Q3g/8JmLgu0saO19
qxTRKHw0Tway+jgHczrlPFAdHJhPbYS/EpYj5LHqR9vHRNcn+U5yeEu4C7/1cQQZ
49FKGL6+jcT4E4TTFZOV5XZbsGzRPDeuBOfr2OuZVUKScCZkNyUKK46hAjPo1VnK
DzEvJ7pE3Qb9CJ6/hhV7+b9ouptb6eqcviCBi7o9u4BfwETV95jGEXPqjMKdDD63
j5JxFNqPX96E3qu+k68/2KV2GREIEjNOGTvLnwl65whSHbAcGmOrvg7z0N7tTv6j
+AHW+6rt+AfnNjP6BZycPYFx+BR6B9dADpgODWOJyA+Vy0jDtBU4xxOm3bKgYn4x
c9clKT61oJGYW0i9vBBFsArUuK5jsmdAM8So3O3c3IIDKx6iQSqCUdcTpzvuRrdz
e5AofmwOmwekZNKUZAPs6kozkuRxECMFz+tyAe9qfo3OnDCZqZ3pUMOUXlcc7WiE
5EtxUFNB4xkhA4vUtieZ1cSeNOAumI6USHlsCQDG5bx7GvGOrz6hYISYlXdqAu8+
v9nSWYtcFo9XFb8lx31jjOKjOSDzqTr4e62YhtNllaH/d2W9Fx+Y1mVDFiZfVoRw
i0IsAr1/5GG3vgxL5EUx8aUW7m3449i0KnrBPbku5m9J5wpqCs21J418Y53Ly8Iw
NyGf4S2snsSmQUc3S5tys3lWT5qJnC+l1fP/BiXjbx6v1OsXzZkW2OgcwoSUI9MK
N2js11GKrbL0GfHbkMHjl9KDcPpB7uGuedf75uu0FksxdFFAZSIAyNlkj0kVMUyG
28A4MSvMoAjxX/6UK5Hm2otFULPcc7t5QPQP4m1Cw08o3/qtB66vsscqqzkCyXC6
2/BfxQoFuGzy0e8r5zhpg5ZgieEErSoXU4tnVKRz81k19kofADgwzZeG3+xLyiWl
LWc/YnQUCgDRCJLKXGo1cy8efS5DajhraWK+EVdBHsWejwmQm5317joMLi6yaQg2
1PMSS97gBwBsIS/QetGUWVu2eWn3Ev+IIUJTRvsr4F8Ux4Nfs/JZWPyOAB41m1EF
y6e7Su21RegKgD3bthkG/fo+QxKlpERzuR0fWJ+0/fUcZzPlCkYhEvKGKaGrjpqX
cSg31fnbyyr/mON8OHK+enphKPuu8+ob76+TSYk8Reu+NG9yNvy77kTfgy9F4+Q9
TqzS7o8dojDrBVETb4XpgWNlbu1TmhjXk8xXWHuQ56Q5RPsMAsjJGjGTQDqriwUX
WnHMURzB92L7I+JACtlcRs2G0PAQMNlNzWVknP9qhVZrA2+ALnms/RRTPHIe+q0o
QWtw/TKGuuTpmkctz/wS2ey3ELs/DfhpEBRgkj8DpwNOubE368l4COMlPPgttDku
sz0c3eA9yPnWPBAFsqXdD4Cv97j3nPf75Psn9a6XfhvUudBVtF8qksgXCtMuqFZD
YvZ/G88mPuwoo/36gDlhvKoKhrmJSATVAE0ux2peqiBo8tSCoshhW6g2DoX3Doys
i6Ml3YyuNNh2UyBpC4PaOS7n+/HmUdw6oFdeNwJkME6bsg8EasFqKXrCCPHOeSUy
MPVn52gSSPXmSrxBVivAi/J8g7TXz7Ntivrl6pQuJIH+Cn6RKRSuNc2YBMQybVlA
7NVia5GLS4YPNNJH5jxfEETZc8IFY6cbT4ETwzN7WT2RiJpz/cCKy0CHr1hVAnLe
zxRS+7yDQqIcOORB7pef8zMErjAcw2P+dE2pPPSR/hBdBuXd6joB9ACPSvHHpaf6
5LyrXGv0+rkVNCxmL2X4LWUn3sO1/BAdNI4ExrXJdrZy6OAEIRZkrWXAxuCRJ22k
8dbatBmUkuwTS7THxtic13xjIsR4A44GGTZn6/cL00xFk9P0XpeITmOi5TY/hpKl
wyrFfhyq6VXKzX8ssJPN6SXL/jLxQ26Nr5drrmCgn/WfmAWtFa6NSwneKgZC/j7V
r+6ewUarEtm+8KJnyup2bklZ+P6RDUj/vItY7VITFnDAu7BHyfODlLguXhJItHSf
cc+lOfZsjpfLYlTDC38tJmeWl2lTZetS1E4NT1lc6bVqkGEBCz1LdTZVv1Rd9a4x
Wz7wETVE5qwYGGxpdx1pjlU2yaFqBIbYe0IbCATSfGbBJClCbgi59i8Ah2KukEhj
dukzvMOTEsLAWd+aqJuqu8aNKDUidMcGcfkCUTcuAqLY2hTOwDT3/9eEOd+tOtfY
PKjKgo1l+DMGj43Fdj7lCMklrpprJyJygnwhbK/DA2n2QxYio+ujVj38yVGGJvnI
v2puYfDu3MY0HCbz+uzeW2S+3ikHfXDdhr1JaQiLA5klpJjB52IlKd7qJW34JGWx
G6rR9mxUPo8ipNaTWbgM47fnLmGbOjbgyzJ0IktwWpuH0cp38AfhREHVcrQLG4gS
R0vIBG6k3hhBmrct7BETNClkSliyZygDZKq0eTIt0HRAeAvS+sXcE5N5Dqq0xOfO
B4jimujEszjv5jquHuzVaxZjLDjsKRT4sYtQfYJrdgjxezcOK3U6jfBZ14rg+LAC
R994OrZhRm2KWvWc+YaOGR5q6Xy35QtZRiMD1eYEFm16n+YKUdRGLeHIG1sGW9FA
wVsGSux1z44pi3g0YDElW/sR43ncNhFhB6HGsUo13nbyA6J2DXcF5+NqxFMDK3NX
TeMizL26GHS/HHmZwe1Ud42vMs1TJCMw8d8Trar3jnAc0mZky+47ssvG6I4R1z4P
G9stnVKckq/2STelJUEc6+crzlgxnNKULZYNClBYmWDU27Y1LCcH31NAl7mgE/td
LUqtFwXbnm9Uh3DoCdfu2+PpLy97OAG+mPu9zRCCvj5eCx6K+J72amRzYD4phGWt
qXHDeblrfgfuDlAvuiY71T67Sa5DeR/IACrLLdQbcHIuv90jyR3VPs7yCbEArZxv
XQZ4gD929syHigGtM1LZWXC0XIoU1B4v1LhQtm4EKCmKDXVp5i7CxV/JJ/Bhpwij
ELCqA27mlTa/653weoQ2ymopuY7yAR3BvnvYCppIJ4xPwZ9rqFwp0N+ESKEOd3g+
WjJxzMvVNIoaOA5/cBFCnSc0J5+1v3s/4t6UBDuOjDEA4FMFZO+9raNin7uW+M3h
8NQ8VTPq67lbUz5kGPh3zcPY3495Smb75BkT6WDcsSGF5xDDrzhG2sOpbZDvzHUQ
d5mz3B3P7c6LKycefSRDZgo8XaaXpo9BISRP/HtmXotwrm5BxnRtr2cmRDME3Aa7
R43OT+FfxZuXhfcix0i1OI8KlvDM+Tn2yBMNe85ea+CL7/fAxbR+882KWkrkY5v5
T17iEFxIO1nm5NpsKjiS9WeDHOv1YjB61IP7H2A6ewHu9Uy91Y7qs/oKB8i3SLKn
/WHjVLwa7nVwfdRed8W+HQB9hiqigPa2C/O0jLSHqFU1Bk/xXkDViLsx92PIyLoo
Ka1NZt3UjytccE3WkwRxQZB2VRZJQSqiFTDsJ3SuzSgijyY7QH97s1ksI/fw9lZH
u0MjzqfcEzb8Wd+qpEZH6XvS84sDfGl5DuJldfYIf3BRZQj++5+isskll0dhJZ+X
0NQV/xUuG92ZH1oJeU9wjfZCAyQKlU8FciWvI8ZQWghvumM2GQFMvOmNwhkiDRlA
RJPPV5Tlm3RiOtyLQNTfCqWlBSdG03h5diHtbrkmUc7t4en9MgRShR2h/wuNe8fj
1D/r33+DV1JIjv/lWY451Jp0IKJU+usTlhgdYWspA4MUDsIHYbjOUHPeo9JMa16B
tPK0Rb6aUByZWA+Rsm8EuQ7hLqTnUoYqR9qi0Z2rkYP/h4mvIR4MF41mhIfsc471
JEJGuV5MfQkvnzHVTMh+lB+aHqiYutQuDEBz6ceLkOxOw/dD6xTBSi+2PjaYBNui
I0NPIDNfl5pH/kgZ43pJjQvgcV3onEHjgTp3yEa1t2qcC+vdi4VncMyTi3XWErIg
gtTocvAqBKnsZZiTLLHRTAYe4alXUNQ/S8CCNdV9OzCRq13NJGy6qmuohhbYe1wn
OzLt3T3n+9SzKyqG081DxzvYLbgtBRIIq7aubhw27nOpfIsRjW8hpp2vaInZAnnJ
AhqU/mky1aYJktZDGEhvwMqcO/T3HGFNNHOp7+DrD8tYCeVAtAfxW7+s03AhfOZq
H9lf4Uyku1Zca0ir3xm8R37qduMgx5vDSQth3wt2BUjqjl1U/UNkdoDnWi/6CCCG
FsnQrO287gWRocTY1kKo8PBFB+i7/o5DH2dvP6SaELFLhySIGyvLff8uicYUyeSM
eIwiluD0qStvbHZsby7+wrYjCyaJ3TJ9JMem2atDOurWhsWpcBpG3WqGfwUo4yFt
bynZkOhou5XCVCXB6GQRBpV3UsK6h6VccGvmzUf6SPTHtHpaDN1UGaZN1H4CGkGE
wHz9TYRAMenxBHxIgmnG/C7dhogI/KyoLSRj6ylK1Nq6I+0TyqJ2boLHy+Rlclw6
72vnPuuWcDcaufs6cjF869mOulYc/jJAaFvmZuwqdf8EzJuqypKPLy8BgPUM7uT8
lIwG/OX9jTSy+O6twcG+n9KCA09IVliyJsTggT/Nzc3binUoqhlrwkSKKUXgnp+e
5HDZVzVu+CEu4Guj2lmVmv9EKQ7Q480KBIqlJQSrE8cmtthzQitVW/DniVMDvdU8
NFH6D8OVdasMLDb2ZNFgCFndUcerAard/F5MfZdt6f5y2VBCT2NKDRjyGckkGG0Z
aLArrgHKeSBXZcM/Ny6Ndxi4Bt014zWtIU2ZuEB4A0KaQdW2ITXYR2XjxsYFL7hc
SUo+fxylUJVFild2BfEC1bNj2IN6L0DTsrkYSUcemytQyusqXgMtaXCtD9a5jzPO
PK6FWKfUejlHHSwNfnk23NfOMu0rxPnLG+Jwh5bpJDAVOisywhGVc9fUy7+78hBR
sWMZ0Bo5dx710AmNbuIjSg6gtxIOxG1EjR+noQprWBAWTCSUImZebWVOf8gBCekc
CUQhqZ0SFuPsZEb0tFkB/k+3AjHCq8Y6LHQ/2rIvgslHJrByA8WI0n6UtrwMBj6X
QSVd1rvyAo3mz96aIEdjDPLQgq68VuC6ocT+jp6lqhs3WV2J8PjW0hGr/2Cadogd
CHeFJxi4RQMSM9tRQZ+acBojXGIFvtLhSEW3JCRA5QGBh88N/WIxLTJh+eE8M7+Y
34aNpcd/pcvnAcGlbG7zgw+44IWoSxnKWyNhpQOMnmwDp+o0zy8Pj63d/2Xs9tlo
RqoQgrALoAnay9UHLCJDQafpHBnjm9YrZrSOUwCQaVpCx2P2gG8gQMzI5Uxhaqk3
/QmKMfO90+HNsmH8tXz6UkmTvWF69v2ka9Jeg/dIMeAvljLS0xOaadnvVKF21XGd
lk0sgLn9tFQwVnuwlN5AiSAXfK2bCsRAg8AAWSttNkQhiM0N3NcjH1WGEfJfV0/s
hsWbKH7JCTWKFiTyhZTj11cTmoLMp8D7T7hQqVk5bUTXLH1iLeauAk94GFuZRHl2
RVmlTuYiooP5qGdpWQPqYqyBIqbj9V+wxEcdQGXAfq/TTgg1oTg6LuWMvyHiYoy/
exEIkVdor0TCfpwFVaPUUMWg7m92ehtK1S9J55HUSsQMRqZi83zAFzBJxH9+Kz+4
HaLIWR8LvusX4pLx8niWviifne//AuL0zjtwgjTBDD29Z8XSQm65H4yGut25Nr/O
pYbA+xCN70Pa83gvhGXGwQLFdXW3Q7lncsbkSQGgokPNGh+xdNvubA0cllBwPfsj
xZjGYmAiB2SUfaE30fi5tiD9xaOOmM5BtsPI/dn3AHYNK20dkLww3K/kYKHrs+4l
FWrox+6yID8Zi5vUCa3ogpS4lK1lPYWwykVDOVWPQ055IiCy2bijzhjRMxR8+CuW
xYmpoh5/60Z9Zhpc6qnoX7bniRktlICuuQqFQ+fsc2QQhxrg6/1uG+2TvuG4e0v/
DJX1eCVUcqeeS5eFIpyGlirMt08qAlZAhPV1VcB8uHIyrolxRySLwok2CmqH7+Yo
Uf2PYgjFoiu7lDh03gnpBj5jcUOjxke+XiVLQEIg7oE2jmzg1Ykh2pRLewQcOD9U
VMXr24qUaLDKq/1LLz20pGZ9utvjnEqc8la31Q9Ft7ZoxHzfVx7/iFb3F0m8Ccvf
PcCT+UETefecFcFMpUF5OW0r+9KRW5cGTIDzgIJ0ZPbi82NWYMb9pkFfEEjuMMej
rw5DFqj7q7Q/RHFJsccs1pjMGWZ7Kub+ZH7etr+oXgSruq0meYzbuC3dUKIp4zxy
HYYpu3IPTXbp45EiBc28W0ijtcwjNrCUG+1YogfKGFN+RntAloSHWxXMWxav3t7H
fZmVsYUuUsf6RFsNG1ppNtAdz6peHc3Zdz7aRJ5sgPTFo7bc2kXcAhb4VyGMjOQb
iOLd9VEAuxNGhUmIe1679lWn0xMPR0SKeZrW9KyTyg8MvHyTLTUi2rphflTDortE
duVwOaBijzztf+RWi7eRnvvgOf+DRMQAau208oa/nYRLr6igvw3JD7FnmaJUQAL9
UV4RpCZZbQP37e+5UpDywoGczsDLxwFpOJD6hBoCGxTj7YxCKRMYzZyI9G8UcMit
k/rr1Ix0I+0JzCgKJFjqXeCiJNTXuo0C2W8XJ+Pzkbh+TCVnFj48Zx1Tlm2Wg8ph
TRMTWP/A8XE5+dsbo7FLlXu3c+SMGOc/37IWWa6c8OG+ocDCBS0Ep59GIfJzdibk
roY+isxsIkQubX11KqTISzta7U2xRcoxSwGXcyQuv44U8CXgid2ttvCVmA9zZ0wW
O9nI/bDeqMeM4Y88YUWM84e+DLriKr7+v5SojiZdys10FXOteUhEjzXUPZeXRER/
rWMslqPI+AeLBl7BP7Zd5PGIVLW8uJYm6Cczoo3PpH1GieLFFUmRFg19A1Tc+IZ8
QNXMfib7lhn3i3qjnxxjGsCKrhMjBX1r+lMj66hUo8mf6QOvgj8VphhNly85FO1I
k/wmyJ88NjI24JV4DgcAiw9xW4cqZKwL17rpmwT8OYfNnQDmKh0cIXWjJzBnbsPG
FqV/D9wNXyRdoAmgM1c6G9WoG24j4BOFJpitRTmDPyijoTcrIFB/MbIRF102oKCo
/D5i5MAUERPiO2gzDTZ7qJEXJE6W7E/jqxsYM0HrZGU1iRPUwDmwrS2XtTFs2d1I
5XL6FSygAKr7DGuOI/TjdlAwa/0HZF/N5ZtKSERH31H+wCoxgxkPLDFbl73+nSJa
WUgspJ4BeEA7wApvN3AZx6ZMtpuzBGff3liwq2hlKo3iqI971C4ceG5CKTePaPTQ
dKgK1DIOFut/IzjVdrM4pxJuyZW2eIS4mILYCJwvcOHitBryeF5fWg7/Z6vuWM71
hmcVyRIqN7IXPE7/5QilVonMidf10KUIoWXYEAglaZG9/yrL+C4ffZqvd7I/7bsc
xVNk+fy3Terg0ety5bNViyNd/c+zleqWmfr6yVlKsVtQcz4XRQ088hI05L8n43Lb
WVq1/nZ5sJf/q9H8EY049xkEeSQymG1vlc+ctEAT3PlvmZ6YwzLdNK3sXyeedyuU
oYD475Xt98sokA5OUdAd2FLy46IU5ezxXxl5EHsWC2JJFNVAQKNgOzHshQW2VBU6
6C13Xez9mFesPYE9/FFIWmpWyog1DMzm787jCpnZD/Ayd25RRTEITC1M75NIMaGU
GWO96EygkWIoAJco/qXEKJmeVi9R5ivmXsWO4j7PJLublu2Aet044SUW5dKZlDI1
K/w2/2quSHzbTpuHZd/hPtuMc7GJskTvn8DSf23Dbkccaig99TnhS7rk/7l535+h
aaxUgjoLNjTf/sP38uHmVWuZFc4J/4AAGzBPYLECeAMsbROMS63qIVbrwJhMunqA
xF9AgTyzaTB06zeLxK4ZhRoWbiGCIOKRGVoDyuqHBXHbOwfnCwQrA5Wq/SLBO4L2
F4E2u5WF5Lc+mQ+Z9LUeRcbTKORFjzETYBOgaDBD7pv/Xk5+/wvlQYA58bpT02tl
Xg5kOukXcPB8GQTvvnO76BItzgTI2gALlK/prvxP5HvrPAdAzmeqZHkfP/ViDaGh
ovAv4tu7XMHS6OYKD1IIiccfkVR4JlpLVy2qZ07zeSKkIR6+R/DUhoM7SuzX3+74
ydOVQ7vdDsmSQY1vzoGlK92ClSYv/4Ije3GX+mi1szvR4sowQdpqq2axNxNVSnuo
voW6K5i9QhdGBJxtZrFYPu0whBbhWIeqSLxmjDYfX3OX1mdbEXJLdffapXzrNDnF
dpk33GhCIukSklX4MWJaBLiPwKpkgKOWJMSxOmRhL5kUpOrG6roNbxXe48DG0DEZ
swIHTVfk3BYvVVtvY82bCXIwwfOA0S0jk057SVRYiBYNFl0vA7ZnHifZhSnx3KmR
AVIQePUADvXa42Uathkc+7IAojzf8QghmhGPUhL3USdsoNJREnUGC9h0j58hdVlg
L0UWbjzkACt3qb7v4BDcAP5yQA7WW7nyT3lAkmkAOL62qHSplmpHjXSK6mUF2iiZ
oaI9S1vW5j9T9vpPosVZBEdeDBowyIw7UwQQEVXCsQ1GyQqerMNvI1xBP0h7Y8+U
H07+6iFK17kHmiWKkXE9ISPQ2Ttk1TDEhf8KA9QntK/2gIyCJvejY60ZRzOBAUog
iL2E1xrvMyt/YF+XHnSeCq0D9D5ydRJF+lmNVT47pIsgFYFvKxHmMtQhIRnt/zLv
YD+ffE0VCTSxcYZa+35z6ddWrMtYaGxfk1JoenCWeVa2gVewWzS3UrwizlixXgeq
NsX8XIKhUy02j07DNZojWA8yjn0tbfd/Ku6G7kIwnQfdQcb9tmtAXvBgnV4vHK5N
ozxZK6bmYVRiIr1HS2M9W6mLRnvG7E+fZhIQr198zzoZDj21by3TKAGUNjHMBfLl
vnvUCHeK3choKJJwA5DAe/hl//sOz2Y3a0CNgN4F5LK3XSipiqXqABIaMwUa31yl
/uXX703OpIETQnihs8ZhmKr6lhqjdh0GOU9H5QS9FJ4ccSNM8TRqgdNZRhk3UwgJ
HAE4AOebHIm7O1Nzer82ElNXNWMBkLghuh2F9LL2MOdJ6C2HRGhOYmjAEZIcDU4A
BW20Fpzrrk1z3UXMwL0GMkg++u/u6Ha2GRsIUzm0FJG3VSJWi2wjSKtpdR2q9Ds/
T3OL9PEz1xXMIlwrkcdHUpFjsMhKxRzIc8W3CxKBcAjDG0oxf4Ox6K3eWxQJ0Al/
eDiJYQq7q0RxDAM7mXaA3N1WsIdUQl8rs/dJ4kmuWHp4wR9uj9kGSOiIz1gmw1mz
5nYonznQmbmSkh6R47smYslklvd61OshoNCXwN1a5DO/20g+9gE9G7+7j/s9+JpG
x/+1hWdufPSkbhKiCWspltXgl1JYcFAhatfYHlz8hUt0nXwYrOQtMlmRNuUZnv1d
y/fkylXVQaxRVVL5sXx3RKf+JLZp3Ke22UPVx/wha+fvXD7KjQD+mlqZOsoqkSDM
ZcLHdSCD48BPOp7hE8LxTpww4tNwrywjKcqrjOVd18BGT3P7VjPcv39/uyvnALho
uZBnH9jrp09luMX/fGNoXEUTgrYGzhTDKZLx7u8sa0sRhMTR9zOhkrrf8g4lxpDt
Eqbec0tNazt2xh3xo8+dVGISUokkuP/0u/qYgziGnXR0lmWmvl5kb0crRBXaYeIY
mIYytvXsZFTybd2DpTy9BFPVwF1gUGZa+yysMJrn1r7GkEFzfKJERnyk1K8gSddK
Egp/TcJbwT3e/zdSx7EEzo8zO0qZfXAoihDWU0dPG5KF87NQNrJP2Bz4fMFTBScJ
dmInGgZcR0iyHZPtbsw+zFAD8N/mu8dtPBqwPAHAnNAh+lASmWOMog2d/WbdytAG
DfD/zVVVb9lKRJQmkUjm3a8tPuIjnyhmFyG+DnKMj89LoNwRByRbe0BGYraGCKi7
CEoykvuw+NK0cK646J8p5qZXA7TYl1UNfbe93soZ1mviUH4CIY+QijefmSN4j5pN
FuuhwhXr30csjYlqmxIHauWWsvfLBGGrtMMhZJcOh6dMjcPPxkkCbiaRJHsOJdQh
L86lF7q3SJLFPENNEcM6kWQt4uVkI50F8ItXuhYhOwNqZtlArk+zlT+s/Tgtv+SD
JRko3wjFeurGYVtRhn5Vpl1bC4pQgHNxURvouuXctWf4tbGSMC60xrO1HscurR/A
3GMitpvNH2tCzW5my3UN7NFDFDdAMeGJlO3u2LWyOrBMnYX2n4UszsjqXqZE8z0j
ZuJPuTQDQq8xTlvh1iHFgNfr/9Nx4FetwWoGDBMXOk/QJEN3yR1xQWBtP670+36I
JFMVynxaZsLnAKoWxU7Jf6a7R2KZFAg7lHH3ci/FpyY8aMHXr0JSJV2+tO8kiq7J
MC5HnM/KQ+GEAgMUhxNVb7ZFfi2a3v1e+26sYB8hFtcB3w40X2c5ouv43itJHXXE
09U1sGYQJLH0cUJawi4jAcaEo6jgMQLIKrUiy0VUUbSXedsPNqcKGpS27uqlheZb
LjeTFHb883YBkj2H2x5PQbpioXF0BRPRNd3Tq5ZwXBPnK0IkBqWL0nQ+hJZuGH5d
c+3rSdGBwrYimcCxf/K7vuGhchMugPwAqw9+q1HkSuCi3Eune3SaJKgOninzss04
4W0KDt9o7fvNXSHl68542GB2IaHx2REehARJW2FrPjVvUWrB1bGr4RJMarBjifcp
nu5nH2aWXjHyJ/hO6Qg1ggTVRegrQjm9JJmxpM0Jy3qRyCFSFoIXxooWLurbtQs8
4ScWLItJzf8eccVYaucZLfDxlVici34xzLQ52RJVocMl42cQZxLWYYcqVHd89WGD
VBCaEbCAP9I+USsmK8cio6VRoC6xJmfX/40IBPZvCARlAqKDbvWFMxfGqnxyX0nC
w5AUV4MWNt3PwezRjW0Cm3owz7px5gJY0JXzx8UztZXS1T503bH3sskxudVDOu6H
9ZiJioB3JfyVLPZ4iOuYWiCTd7khmcwnoXVdZGhz9SqbRSUcNsyKmsOanI6R0zXO
UnzeX6ya4/6c/gaO83Q+hixVBOU8M+bolfMuuI/4AHBFXCNwv0BSAACdEIkivDc/
PuOWFUqScHxRXeT5uwYDJAPIzCI3GmpLXyncTV2K3mxLXODDAI/KEOvgflLVDvgj
QLQGfa8eVujOCJVXnjeM6NvcedtadXHewzhGj7h2+Ue6y4hwAMoLTLPKbeUtymqh
9sMbdmN3je8Ptm9Z/aWcSNElRo4ViVaZmkHJWsWkVWeoTiAb+8DgfjwHwa7U0i8y
9cwIntaED29QlAW+yeJGiD17MutirPiTPuqkTQc3DXUTRC4rnadBRYBEXtD+Z1Bb
N60GEFMf02ndAOUohqSK+hcQjOyh+UaLMzceplMZ8NwszA/nxGQ4/BtNOAfwG7bY
oHMBenu9bDmkQU3EBDk8RqUt6VHHZNw6Jk1kncF+PZQPiY0vnAKKWmkmdrvK4Wm/
VkisEpmjali9p2lbfvJuCntjo4WHloKTFIZ5U5dJvMYHZu5nZwLxBkuK6dvyl2lj
Rhp0q/lyxg39XpeSIc0Qz4/wlT7dSSrZFRpMElMOXBMaqCE7zMW2x41Efee5ZPv4
gCr0EF2r80OUOF+exSuYQG94TdI8Bh/tOCdYANcBLYxh8Rz7hVabVZ0/iIFKB8/u
GT6SD08P3oo1ROY+8uMn+cwAUvbR00aOayna87mPIn+1eWWa9X8mKhH5/jiN6Htu
Cu03A5SCKKVn41CJ1UhytdAzJqYqjNjEAT8YAcFpVHUeuWvIfsEtgWq4hNZTQd4F
UftqCZcHNgnvd4bDAT0IaYQYUAji3I4oqAJtqtdgg59aLbfFYIhOjFejKbZn20BE
cQ2eyrRMRcPYSwCwYxggSqZbxKRqm8ivKMxJ7a+BrTE53Hnsa4S3aFg78RC54Tzc
BR3anOwxMw1bnEOXmTGDYm6IWFEoka/UvqonyN1sA73tLtKU/LGTJp4CwZmX8bK6
owin5Xl55tv1J8vkE/k9oZiDmwkyLALsekm6ldgXQ0My0wbccTwQcRvQUIdEbjde
QVBjUlwSMe0j9VzFRiTVKFsgq2YqwMSbsA/ZLfxxI88e7U2NL9ubtk6UpQlHMr9s
f/E+96EKryF4awxaRq+uz5MfomQUY0VP+hu4B6T7ITi7klLiaLst8kn+izeFcfMi
siaE+P0gnlqNlkwHfIQzKpulKhbUBg98fAxarmpC+C5/qFvkq9kNTibIzZbqWYSk
qnRjpeO0lCp5vKQrlSFsuNxroEi73PSOfd5YtZPB5rvwBgDwmyG9IClHIQaM/y9I
XqX2PoQme57rIlpmTKr8MtX3w0eyEhO2x337AHvPyxCITTYEJRkJoTUhIef1AIL5
O/pW67wm1DCPyL1pHXArDlZvEaSrIyD65oKC9+8Vu4pvWqddBDYyVHa7lCNd0Kq4
iR3jFRrQ/hhP9OjSJcn7foslnmaxiGQkkbPImeUQNxIBq81UudZMdLdtelWodBL+
9CNfTbIO/Vt7JLSwkNfDisei5qNDxcRVcvsPfbkPkes8Smmyt4ylCTqAl7MT+dbu
GytrWAeKr0R3M40en2NJ38MhYmRmjJAOHRxwpQfrMZBpcxXEG/yD+ecrzp2c9hEM
iKmBeXjVYP0PfIlDO5dnZ6O5+Z055qF1I2yiTsa9Pwib5m/rpPAU/oWY2sk+t9dI
6x2VVdWqX30dJCWyHFUR3MrLn84XFWRyO5hGkd+ZZzCoqshn9/a8Xs46CmwFF6gM
f69mH6t+/VRpzFTjOwwM/EhmDyaxQfr/imaVeWxfBEcDBW+6PPu8KGDl7JtpJ2JC
XWEH9gdZslwAH1AZUOSgGfNSEMZhguwO4kBlGN3MfrkRXLrPw2MCzh296gjYcNTg
lpUh5JQeMY9mv40OeZolwZB/ik2QS6D/X8ScMGKuVT0snzN6jXYA/S+D4llVVnFI
NVFwxYrfWLDAKkOJ7VGA+KTrq4PkD51LHusR+qPftbHbP7vtiL29kCz1poTFVnwn
xUuBda75k8s7y/93hJfqC6ysc3A8ZoCW+E05VZ2yMlezcLBUWlbyxq3iokT4HyV8
oz7I5UDXpzunNXKIFDAtEkHH+yysknXFkpbCHOFwAPi+slc3p1Ng+WAxfO0DYGaX
SIZUIAYkJzhUlFKcoekvxLuLfgqd2SI9LdH8HuNqGk1DpEBQP7d8TtOXlzo6aDVs
Tc6sek8JNHj11xRPDL6SuZA6xMOAzv/AYN9nNkRyBHOILUUDjlqEtr6jabZCynFt
XKdETSKw5w8QzhRDV6pUlSByzh9Ih9bsAl7fEhcGDa6WGoItu//7bB7fJ8TRVPiL
fWd4sf/t9Bg8wecou0HBpL8UQqeamIMTA7FzwrsVrV1UU2nbB5FjNAX5fhcsD71T
MozBmTWR8iprJr5nU2mQ6bOIzUiq//lpUohkN6mX0EFQbvUJGstRv/Stjrhyx7fo
42j+odKyaTnknYEVvhnzSmZ60ncQ/OA8VA7tqC8IX1ItdjHx1RZPH0y6Q+J2WwgL
IUEogorrASXlGO8nAMiQz5rv9Z9fOnaKD5R3NCtmcZnXxs1UWRfDPCTqdi6arAI3
Riy7I6rb+s9zmb4vbp96oqpCvYBYHwYw3ODZwzIRzMij3gt0aNLQcYohpJY7CL+f
ACdxnEUP5tvtmydvbcq40yk8hl2/5ZuZsZaYYniBTXQEncj3XcJti/9LxMXT4aYS
MmaTImgeEpT4crQIc9yGyD3D3T8hJ1UHJtoIuG9TxOMplNOSAZB5vbMiFyTRFJhc
HzUd4gdW8yDtqbgovd9ubGrNPE50AMKT7ipJlEGw49WXNHRpmB8VhEM2PuLLa7tB
7rz+Xi+y7yDYtCAmfqwWJcwob2LphVINZk8zoR0Q/PHUrKmNE6VrHaYFUR5/jlUv
SetvRu+Xyd2NCTZjBwbr4q0GlANQrp3H75qigtyTCjGO9iniIhWq7u1XLu/n1Hjm
oai30QEzpJ6ErTqtNpgpyxuxoqVHQk0a7CSHJ5ZGyRTRPmVDnTmqjF4uYSwumTr9
MRoEjb49N2Y5HOdF8aTtAM93OTew7MVJYvLqwRlUMPJmRZOuRG1x5dmoSCS9ZkA7
20PWtAQJaaIg8kNtJzMRQaIkQzvzma6ePmLpCbsiwXIgSQq2AXVyfzh78pIsEem0
rPKYgX+1WFnqryStX1TpQruioRlZnFeL2FkkuSAcVbg4PPv+M4AMrUcb1hSNGqr/
mGkmoy3LHoDRrIFg/FdJ1rsK35VboFMiZZkmC1dUVSm4l0ODoCyZ3prVehv05lXv
N4X+xQ4GiQhCkXTqm/8o1M5/KmTIYHK1IDSiK+N8tYN35B/7HCK4fcAMrnOC4qSi
Ml4PS3W6Ud/UDjob5+djg8TywuixQVQlpd2K4NzAh3j1YBb+CRN/6LAYev0ld/or
zzHImMkytm1qBie4tJehvvYtl3MAvm+Y9OWXmnriD8AzdBWey+26RVSzrOcgRUrq
nioj+P3dk7BkDxu6q1jPpiIFh1TUfihCRdrokJDsuNtn6Dbq8KYf8bsO1P9h3nTw
4vLENPAu7ECAYafTlBJmOnFGkjvUfQjQJPsHPwISwrc4v8j63O6uhpdC87Tjaj7C
tWk7YzF7AsRzEBKwBcfeHDmuD6POF6iSdfHgdjQyRAo3rClDHUv0VdNrZH9MJQGw
Nd9NpoxYrUEPZlhiM+KPr5oy1O4LgkRHw+FrPWPMjSBJHIWwJr/I35xD+WDQy5XS
cvUEJjSO2M2O+FmOjO0KnDAFQSHjza9uk+IU/SPg7XMIggQ41oqYgGi2hNRr187q
/c1EZb/QSv1GU0w4MF/V6hzDiIsAmV5UmoYZ0Zv42GIyf6O/Mm9hqQ3KEuz4SDag
uueBc/ALxyGFXx9rzoSBg3WyPixS1FCvEMDIm7kIZQPptvEaSDrhSfpccwNgbO3W
SqszfTFGt697EW2bvNOLIaTgA/YSH640ERqEpBlRfRtUCjT1YMNp8m0tZQ3JFJKo
GnQhajjlUDMrMCbbVQpv8PQIqI2e49/gCGd4bZmLl18tGeIjo4PB3z/RZmTDqTdf
N4PDdmtiKtdp+xhYGUKX8sVeYoVHZHNjWi3qCdGbDKth76NPiOhhowae0LevVFKv
QzjWJE1L2t/fo2UuQ0staWG+Tw1QQyj95inp0uO4EpLXEKxJ3+A9ppug0WrJ3qqV
YlqIitmOTReawL01OGg5nHNO2Uxgsrw88BW89C17IaQEcgU9AZIoGb88/qjsl+fA
vf5atAEEsM55YifEGN7Ce3t0MEZTCM+sdrgtEPAoj4nYinPKBzE+KDsV1fVBhKUQ
+GTWGpTE67ImwQrdkD2W8NzIQRQl+ycQX96EzYDu4aIPHCQb2DONRKvo6/MrA4G6
hbsANj+tGLvMZCJViODY+WFbO4N/9nWYvW5Mkxjhh3J5XzpE4ttZ174XL2iEcDt8
I0qA40WIJWBsErqXSuDrbZ1UCv8TybjnZXZfsEYD2l0fYDZTQV47rRGqBfv2c6uz
iOKsee54yLXTpu8IxFDNwkeqYh7eBN+MkbWzKXuDyfV202WPHqUK4RuIIGzpDlNO
fosd+R7MGI1+dOB/DbBra0oL0VaYit0yx62fl88PFxEkManNOJwfKwBIYHV5AmDl
DdTKf73If7I7xtmeObXyAMXQarJG1tWhUwiNUQLLKRxGKXCoAaeNa+DfQH/J2wW0
7mBVIVPVWC5XcZjqpOdQENBep8VCGZ+X3zP0hK8NKFHgUjoLTld8rCamn5hOdtRQ
n0YV5IbxA+7SBwLGNNFJLg5/sIq3gB84Y5OZCpPEiTjZec2VPHjrrTuwW3qicRJZ
V3mQ7kH6LO5gNdjlWNrf46SNQ4zr0ZxW89mkjPb16+q06T2u4Dy9WcKpS2t0hu3s
vhfOFq9HXMXfOVV4EEBuqz0Xs8EWM/xY8umCNmAW5atJco1jBSG4Y+D5nFuQfLzf
nEgGQBA6Z5YarUzlTrRCBJlzQXSV8ca9UWAIRsxgHtrwSpHYK4s2yqwKPSXEJCoE
WnHJ0dPFdX3zOxpV7HnR2mJ08P0EhuAMoBFXyB/TMyJXheXhKbn3cRYf0QgbXqYH
RYTNxjrwi25DwZ3PlyUe8jj/6b7/FemGgf8NxcahWpJxNQ44XUBBkDtDCHg7b5ud
w21KDnf6EchRlvgN+882JxRYRn5m0pRGh8/d6GbEzIEjYAzYw+deg27aAkkGtAzD
fprdYK9PYIL1rMDNeQs0XN0Qcc1sAlMrp6T9Aw9ty4uM6Dzz0eKLGi3Fx1Bjt53/
NKMOiaw75Ub6BibtupBkUZOV1Ludck14P7lIZmEZDqJoYtXLKX31AnQ1HunemXyi
6Aeceqs8G8R+MwQPXHVqPsAdCY9HC/rbWaEL4hQq0iwxZ2iS74dSHFL+SBMN12hI
rMDs3jJL1H5O2H4Ke/D8uzMa7/FgY5BcvyyiiA7sBRFVU6bJ7a6fTFHy8i7bsK2L
4I/Lcl6qdl3d2fHTWk/+jayJiO98soZKA6309dDU8U/QNHH1vbbbztJHtiTRvEuo
8rLSGmCLqf4u4s11FzBNwjfF014Y1HZh5/RUZPm75M/8YiCaX0WmKiYyw1I3L9Wt
cyAlXFAeRcQ19/CJLskYccHalzHawHagSKouMGnVbx+miwsZbJASokDETLjDTiaD
kmwdBdowYvosnB9JPxeZ1PCvwyCivls14WYd1Xu5r+su2Hy/hf2sdyj8wNoINuPw
8jNss4F88NknNKU64vM1vWnQXqxn6FwXROZAt6KgLEstc0Q80LNv2E/fahZBFx0F
+JuJwxk5Agz+nBJ5TOIbUi3NYCkJwRfeO7Mi7r6C8+jo1dwKxF/ZoNRnZsmfOLHj
3nbR3o9fd6D7czhtChQJ+qb+opkz+fcelYLCLlMgTZT02IpV8UQ3fcYz1NB145UL
I7L3UMp/Q5i/Mz5cAAdg4v5RALT4wNEuSS/N3H3RiYAyvEYiKsgwFLKo9JuwAcHb
DN0hlBuLFW655oRqVG1Y4F5TS5YiPDgJFKtZ726sXrmurjPBmoSi4xOy8+4tgUxD
d0BDKbEuvoJrKlh6KlU6jeT1iZajZDGeWV/4eODasOe/Z1X4SXl+VR91HCE2flhO
8KmR0Nlf/F6bUPfcB9d/arkonP/WaHRoe3lgxFU7rcrlW49OyOKP3nSMlItaiN+v
mKwlqMQsJsb9IRvyKuHCfcCjJ+o5sIZqDuAb5aeZ9oXC6AX+0IuYgdoP9kJps8n3
Eimp05EuYYJw75HmA7v1JsEmWQM83avhWwGBc7lUZb08NxF3UxdvVOSWOLyU39tr
eb29JbX8oShEXL+1TNfXXweg6a5riIsH/wR8hlPs6OU/fAjWbXi+XGSjJ+TWCXRR
qwZ729TuB9TkyFjfdiDxH/nZ4KqLzWUV3564tk33ZvPZOx3wxxCb3x5b4hiX644D
eixHyfybs/YPonFVTl7IdqUZLbKI6zqjRXMBYMzYfbv0gIG3GrHTqHTv8hsNPcqk
jzTorLUHzVgH41U3mLkQwTc55w6fTCtKlU2acviZT4rHEmXbPManxMhIFlUHmMxu
k719IoNxeJHEL5mdrfwjUk94sC7OB6G0WXtkfut/ajiE1IQnWSIoX3Pn3kjE7Vde
jF0sj+eyHmZ4M6Z4mnnU+ccDPkOxT26SwCytFPNvxGo5wdLIcSIS1Iqqe+81ax0O
rZRjqrNNefdgLpSnkq048Uih0Hl5rQlv2FngCTnNFpOhjsBPr9D4CDaj9HMMTdnQ
JHFnruZgGBO0AHJDxQn04OmjDP5rvxoYWj/L0IZZvnSZy/8nxbEk6WboZVNsvhIb
uaHI99uzMRpcGrbOvWrkxWHhm2UgwG2jEkA2vOnd2N2HVfVGoVR/b/dPV3nnm67k
hTmd3Pd9OM8I0zlm4STcqDcFtG9hmQXxsjO6tsHR7pEcViBjPw+V+RK2l4bkM5uj
ljFCbjGoA5t9aTvOA7yNEgeEhF1vuhZtqi02PtRWU1TiI3pFBazHD58180Z7OkxE
ZbmPbm4X4oC+Q4MPJOlktaG5FmWOtiw+15UdEmVPWIxjWzX0IR4E/zh0UFdDTXDa
A2kDe5TZAY8XXkCXNLTq3+EzzdBbKWXBQNYBnOvcM9GBrEdWoi3KnGeMnITJy79x
Ep8UMB1o/QAnoGo0+aSxcWM9FA/wXw8YhL/h/yqpfPUGSdp6wYstZBvKQvgIrfz0
nAnnu3TSCLoRPK2kiUaDGEvXBcAU48ouP42Pnie+EdliY1GQEkzlQTOBLuDWb0w0
LRSx/xz40afq3oAQeXNFbXKiAtKlL7Clqnzb2JOmx3Bg2m5OTr2p88SXb8WlN5aH
Zy0Nx/Onj6bG66qigYNE7bfBZqYg8w1x8/yg3FirW66bkW2uV+QHkhCu1C9oYEjY
R5ZFWdN2x60GQ8mqaRYdgpREyWflpdYVBdzxYlSyvNJdORZB5TwcI2rKVXkwKsQ9
aI3P350VpKvjNx2tsPfim0KLCSqPIZTAXff9JlRMDucaIZC7JlwftIJKgnGE1gXK
7Fj1nEHPd7K5ruZbvPvSbcGBzwQ3X7CDXnnO9wAJ89HWHEBAPJYum4Eo+CWo40Sc
tFIwPuYuH+Q2dcfn8lrWKy6eGp0VtlIqGB4VsYzTDnXBTXVVKrYk+oLo6fV3QVF9
8+OaGOIbpvDQ/dH8pp5e7WGf3OfpZeswXrpPKUqp1JE6O1JMTGn+Sf4i7wpuEj5v
+0J/YxGBf42tWhVW7uRhZlJeoQF/Yo8ewLXDWKqK6NWeVxa0mfoUHfmKWYRylXwp
9BJxTPd/q+KJ5fVZVbSSlRTgO2M0LGFe5x8UZFnl/198arB4sPeecmuNQ5Q1zwON
HRushD6kEM0j8xC1FG2Ptni6RelpW8vyHCEA5vUphHtL4cg4I7wReJAd3XdsoSwy
oBJtHpl6A0O2jXmKduXuzI8TfZp50Z2Ye6ITWr55MoNkAgMlDParHDNqbkFt5YBy
WA/vo7a5zkVwKRuANdxEVaynENXelgLz559ck0jAsjeek/+hnRfuCrlUWXliZ4gr
yk8QSSS6yjBYZEzd3gu1GBpoMTyuYhMs/wScFNzaMQ9/eJ3yGpYa10AQ/6TReW+1
1bJmqNR1O7JXBwFfJIJ+cQK5IN8kDa+Qqkql8s9KXooiTKb9+k0mHKAz0oidzjO5
MevNUKI/Y/Yo/zB4NXO9orK9pHa0k7Yo62ILO8XIZxYcPvhMROUkvjUmZhyma7zf
sZlLgT7+yLdTJ64uh87iiggDvnWKSejkKJheAIBPqAIwNnA1jYB8XHSvJ8xeepDW
G6sdK0OQtacYZ5rdlMpnJu7sdBgheUFfe+5DKA37xgtN77hbWPpULwCNmtDRaV9O
aCkKKi0zERiCGd/3wvcHoL7Pe+YCkOOeBIni56a10yx3/+Zuo6+dTS4au4arYbOP
MVHTZvweW7VwaxR4hyuOPy01Fdwev+YY79hqI0HQJaqUtRD9HrIb2u5t81YPN4lx
tlorA6MUJGS5ZQMvI8aIYn/QIOrRFFhIv9s09fERSpPVslbsqv5tJvEPseLeYn3H
P8kdoW9MIwdyeK9VO7EK9qNXHrE14zWEoPgXlY1T5gshnrLPq8uWz+SeTnKI5DRb
2RhvRUfCy+v/p7i/N0n4M0QiCbOvqvKZeLzsOXXN7JcO7UB2Alw9EwmIRUe0hVwH
85p4MBozRhbLPooB2GAcqhZfqgX3Ej+v8DPgA/Vlmzze3tST97ebWPzVhPpIoSM5
CRi8eydt+YMYoQvi/ZAq9iV7R5tpcoikbMhtF3WMGJCugTQA/gcQdd9vf8w1CtLJ
f7l0/q0p9RYTLl6jW71TPfRplZbsgFzt8g+v2VLr+ENr47zjjNW7zzwUUM3Jt0fp
9m8JChyVewrgcTbkbA//USJanWvhTEHumLOaEd6GBD7YGsJ1AKC/KRIFP8GeHt2E
DNyCQWEUOipwwuu2Y/xDVQvgheSP2tOT14DeaCaBM5LUVlfgFKTH6XCDL3vgwo/J
VVzMfUA819OadhtU9RM2bJAyjPdGE3BLp2m6wbh4qkfPQpmeadv5bcEjsk5oFUr1
y/W5VcI8VKZHc+GvvhzTLjP2R67jIilfxLRlQEdqvZpAUrZ/jp2IwYeOhjvL/Egj
2tx2v2UUGnCWO7dFaU3WPvbnw4TbL90bZcqzBt+FnbpOhnOxuophuCuUkfdXER6y
1u4cXic8Kth4BAPnjrsbqd27CIJ0q0FIge57X5DWNvC0fsTae7pKEqnZoHVsBqwJ
sDMrTx8oVjSa1owHa8D4HcDUFBFe1bbT6UMKjujGDZDcpBpEwJzfZqmoMRwu5Uiu
YE6EkE1UpXOp/obkSdGGYB1Ou2jagvzNOAm2+984Owd9BC3IC3Qp/WX0l2WZFCGw
UmDpd7zGk/jK7QdeejgdXg60vEkqUL3LpotohHkEhOShHN8nwRck7ncHIW+wXQXw
LqODw5FprIfIouVbzbkP3eYa+3DGUzCJPZUE9g7aw4K9hBkZis0tLsvtcc1MJnWQ
qeuVL/0a7FDGWT/JxZc6UIThjCS/weVe2QfKWG4/y2VdrcWh3FJHhTFquetBHW0H
34EtTT/ei9hYjKkYgQ7ROn+NqONi1aBOWRo/K5Qtrmy7JrcWz1b0n+yBPRJeyUBu
MD0FQznAE3SLHywXMUKav79fVLMym9F+TjZ9xmBkNn0JNQroow4vL3Q3oxHPKfJK
OO+rfTlQH4W/6KMU8j+lfEBS8PEKYacwCNx82JTXnEBKTVHjL4Wc0fGhrvgnPo44
gZBPXPp1K4f5HMCh8ifuatuZtGEDPwcehAK4ABa1iS6EmIEZIMFRUMIIAFJPu/6Q
pRSvXoVKDZDRXWgF219BIerVRo/IZBK/CKhcichWtbv2aFBjbkINFRdvfYboTP5s
BXizpI3HjdMC/vD3cCzQ/VDWwipxzt8NrLkL6DYDxqtZRTGX2IIuvDveAKHPsmFm
6OpU8r/ojpOWh4sdaPdJmt8HW9xytHBA+EVYmxGC5DZ5ifznY2mUhQWoXXvUOp+B
ziYRk+vhMo5GKQRX02Rlub95Aep2eufKYs1MVOHQujQzM1DZaXmjMrzIzQTwi42/
OKMOW5vLn7qyeFj8EBlpw4RYUuAiXHzkb4MOD4x3jDvPf9qMmG8NkqGVTv0ycg6D
szxOxZv7QP/gAWj1wjJyNT2Y+MJGB3K9ztqOYbpBshP52l6CwyoeDqK2TiF/dInr
0WRKptQPcSFjMe6JMVghtR0FL1Vx/CAjGzgXp/7Or5B1FVKEbsNDl9S/vET/XvWB
TSsan96RkvlPMdsBcgGYD+yH9b4ZlviO2KSI7J7RqQdqITAlYcf7E8mldxJxNWMF
msA/Zp0r4vZP1leP1WFvzHGohRM0zgTmbmDqJTJWyPkSYuAXfQfQVw5LcRTZyHYt
oZdQ7xd3YoKSlQl+jFhQWNmsdkzz3Ucp++fneHrdTHkGOMbr0luXutpCIIkON4UV
n/TkmM6o19i2uoIq4lxFASIpxnb+VnHr2lsbh3ANgAk/KxqE/ZlwDOs/aKVkIxOv
55ocDd/ZE4QWngk+zOFNvB6G4OU4LFrwnd2hNes1SIIT9O36ABStg/5N9RctvQmu
rNhU4dvd+yA+/CyLOjMIdISrmqLdOrGGTtq02ptgwRiiV4uJypTxRpI+CnQ8Zv9W
PYKJDSPnqH98YLs7G1ksud9LU35VjPLHWULIrJmwUp/lpoFbhnTTdKdURLZh/p+x
EYV20f2cFlybFyTycX6/N6FIp/y2N/tlUHqgJqyoOYf7zs2XG7VrfRtjz6DJfk20
XWlF+DAxFwxEybeMHw0+UKx+629Mz3x5tkm2sRtcorgDz+iG0uSxEvqgcE9QvBAn
gpLdCZz+kEPPlqLM1qXttxij6e4OsK+5J031ba+P6t9p+lSS0UpPCMWOYhysCgsY
XL4S3b5PuVlgcqg/GzJEzHpU+d9Xcj0ErGpUIq5Tzh4mKE2diIZFL4g6aflintWd
jcr90VzSxY3y9/l9LGGbVNV5Q1ebzJg+nRdzQRk7RaUafWojsLtgnn7XxXvNeAYJ
uAOl/nVJ35Lo1kZhnSr5YmRf2s2XEMotTMIJK46qHA0uVgW6zumypTS29cSK3AIF
rAgmPw8bBl60JXC2hiQTUrFyekQ86m7S0P4LOTYY/l5uabE2IRkYC0AnVNpNUsa/
j+NUIJCJQptZi+m+RUKT3tWzwKkrY0ZBDzLmlSaWdu3k1Lu0hJv21PjC/GDmppYl
S78rM0JPr6f5OOltrzbJ7A3+szDDUpHLcz5CCEzOAr5/YanzolHj0MCRJK7j/sTr
GAlT7ZK7oWl4XUDaUhmgdewhmpBr1gQCnXelmgmG7DquhBo44PVj0kDOpd5HYREP
T4U9HNykVgVQZWtYOnPlllDaFAaTNEcxwnqHgG90ddTE5YGFG82q3joeh7Of7cOy
Mb7krJNKt89GSRr2euYXwAmxCFuAyami2+rhf87+EgmXVU+bJslVqfsDhRyuOj3H
Ss0uJ83IbrOzyE2V8LELtMFq6vBRxd6oI2qM9AKWid09c+zjbELj1k7kvOM62nSB
VLht5dHMHuTR1GAspsE3TVWKNYv5GZSIY4Zl8Vm2+KVbNSGSRAw0nPVwK+su3ufH
YQzCj1NM0u6OHkSAUQDzvlQnk4VFSKPbXlJ1lDAQl3VVGKspI6ox6HDG5z679D25
OPjBwJRxelSEx3T6jp8NJG8k6V7Pn6Ntx8B0gk3SftHQNtRE7iyJE48KAMqGuIlT
90CzrfxtyExW3tSGyFgQNcnG7UkOPO2DGJDNtzeyjeTTnsfQa3YzE2eiJFvfo+22
XnF5anI5zcFFM6Iwm+a0JZlxtOkPhJnLdYUQGrUlMZsgpoDOsYLOwd2OnySJJobc
JI37e5JE/yKfPUd3c2MRnGUYQ3KKFWVv5Jlm8Xyed+XcTPqNIqAizykqO9ziNVx4
C9Oje4lGK51XZWsogjjXQomivT3NJxWIDgXq5ElmjKL/CG7Fa4+KP7wDtpvLbgXp
VhIyiJtX28zYCAQxhyzd6qhJ+vNJIR6lGwLU/yGUmhgNqBeEsPvKXwuvySFdbwlC
lq4iuT1O6qGSN2lhhZAcUN3kF2gQGB0HO/EEHf0LL77yQ1JkGb1XChZ9OXWl/HZF
+4gihQpkLvrk4hLqt0DtmTo7A4SWmHBsjAutUYiQTkXGtQvAcxYW5jibFw0pDISY
FqdYS6gdeFRDtahAYlizjdO7ZfAAVcd+R0K5G+YLG60gp2hjh5UMZAFbOMIneyJy
EuL9KYTDp1uksKi3gdEIUw8RbjV++WSi2n0s8Dkrn2oQeklVlP2R/77HRlK3h2Rj
F4Ga8dYBLqQ2702DVrG9/jFqBPRem6oiryY/vPOTd84DZP0kdVwkaSfPLyDWwYSw
048VDDSkxVGBzd1FUfLVzFngzs4/ro+heJvuMrLgbksklqoCWRsUqkFZjVzER0iK
cyw1xeocX0OTj8h4QpJlhkEDi7qJxhe9p7DKlLVYmTgcBUJ/mwBWt3WflvgR/GpJ
dwdv1vLeBUjBxcoVl1BP6d28N57jqNN2GlXDelvifzsUy/nk21nAkA3cKq4Ri7yV
Gnh6SmCZevAozRuLBOPr6Pxbm9d4JjSbzcpiH2r5MBQUW41W75FSKTydAX5pSmb5
QZu52GjwDJl+DMSRs+FYvZnDwtn2AnDIj8unEp6qsirHFCx7pEYy7UF+JHvPMtiJ
71rskpdQjsPmThH/VZJeohTmMIY6/PAfFUViDjuI7ho+TlrHqaQCQ/sEVnT19D67
Zp0s+NncdNI8ca9OO+YtlFrofiNDs0WTU6StaSYqPFYh9Ev0zewImjo2mlR93yfL
0Ft68z7lKhqtTpTHP6uNrFRw7aI2taPGDziV58bkVQJx/JEf6ffp2ci2O9Gi2N+U
7LxndRoO/ltJrV9l9rPM16h4KsU/lZ2bHuaAfb4vyD1UPsRXQQe8HVftwSslN1fC
hPfDlaV1kDt9ZeVsSH5jolc6QSjsqFMrw077+hFEw0RhKGHskJWkn4YKLMiA+jRQ
vzwnHH4q5QbuWHaMbnd7T5NxhjXTEP4A8uVFh0oZXXv+N/70aW7rLLxWM5Y+OAt9
AUcJd1dOjexhpCAN7WHxvarzQvZmO0FBmPtR8wwqfNUy/Oq+9Sgco/ChFENDDdNE
tz8nVbP9+R8IGdV0+++9XxUOs/cBGLVdQi8kLYk464Ey7nQlzubcg2MoKL1LzpuH
uNgKIbeSm/xFzGDBeYwK2HDvMRczmFtbrue/jb36aQO9w0g1/idJoCIWmuTKhSO6
+cskg+6WJ/2vlv/p/+yvh6FaFvGX/sMlYeLf4DpQDycgyPbQefTIzT4MRmMxJVSY
q1tMMbDWiPGkfvHE1ihyBmNt2b6Fy8N10XVezgXJ87AZsBh/SOwgQ4CGkWhKjCA8
0PImnc06frpbar8ob5FcfGqXt50ki0WzI4GdeG9Ay0IffC6WXa9CuMnyWGaxGQlg
fEC5n4nyDhE/A8btfI/mYIWhShqW5q2d24aXP4ioJyEfqNqzflzsti7Jo6qWdheX
2gjrZJf+Artzwv4j+B8OfqTMQXL1vDw9hTIXIUnpKCQWvCZjTMp1RxsRZ6MVyCIU
lWGkkAt7G8N5rQTMnSrfqmdEgFG/ADj+6ASR+J7gkIqmV6LUfJK0BNgRZyREjyE4
ivs/qn1jNbsjKW81o+riJiolQZBAq+21LoRju7ph798f/F22DGc/TAclH1iQmrKK
hwgVCLEoZztbYGa7WskViA5jW31t6Thtly+yz0smrcpuEdAY0L7+9oPI06bbGMKT
drx8wfycO1Si2iBveKG30mQyhEvRsIIjqip6IZvtd2dZ7xKoGlwGos6CL2VmBYoH
G3rLZImAVwlEcLZyKIVaQ+S8P6jJksFP/GM2MU3Va34wl7/b+KEindNp/nvFTF9I
n+oPjIoVGij86+gry3Ddkqq1m9oLqEUd96u7uYp2dl0T/zUD3K5TY3Mh/UdSG25b
+UBZE5OFvL5Tok11mjXvb35AHKC7FyUb8f8UrMDNFa4b/LCHy+kobOdoamAzEFHH
5gWhdLsirQ5c525Ufpl1Rh86d6Nrkh5KPlu0XDxAKZap2Y2RqpHlX+4MDxTOT4Pp
HJjm/aBeUt2g+2faO6N/onIRxPT+vsgmLVWISHPkGXA4vxGYUUtfEh0KQMtTKspF
nM1iwZ+5kZqJXiYdfD9DBr0Xg137pNmLHqOo5C3cZ1TnpSptUqbyRhxL0x3SrcIL
ZWz1RFYTDvh0JtUjZ6w1hR/8slTtKnS7RoYY04OVjDs+m7jpnDZNME90laRW4llJ
DSGTHcy4m+FwbIGKWmY8D4bFRlWx3fPeJ0Tig3z+7XuaNSYV39CrxYMem71I98hT
j8dF3ogKiSEXQKoDKQ32bIC/gqq11d08YikUksSsCjx76ER+8Ti2J+d3zYPyh/KF
Kq/VL+q3nRJyYZ7dePH4/yXb9+w1M6ZoFiQ9CJKrl7mxFj4suwNquFn+v0fEg1Ci
GlE6gvbUQmnwwu30YdwNoNE4T4eQW72JQvfYEcJ0hOTKh02JB9CvdRJLRb1uaKFJ
tbnga2ODb0Qxcjoxy25K/sp9xn7n2x9LmhUqEepwoYkwp/i0gN3xS/lIlb1s4Mfe
L0M8VEz0xfr8axcH6Gz3tAcOjU3YmlE7h+7Hznx6MQd0gULsOejPjGTdCaT1SqmZ
VcqiWHz27gtQ6NcpvJzP66y5dn6DJCZEDVmyXtPDnSXu8TIVqRVnmPwhKWo9l6pD
qFORir+7293sF816iQVn+72bA+MTmik1ZDVpHl+qptWcKZn7sNIRbG7WVaUku/Qy
lIhhScngjHF31HsMSisOKvsc4Z+u/7tTvRMhvO197FGT4JlWlYDKHvGSZ1v5we8V
XRt7A2Ba+ZPMuul7fD9feUzksbaY65J7ID0cXdetbyI0QIUCg4LS5wZQiE3QOcTq
BrTa7AdNRzz/DCxuXbfY3FdWDYMFcFFqdBT8NIa6XVPG7mpDa7Fm/2y6kReFTn4i
dsJChCNSYDiQUr85D96i79dR1Df4ZNzGnyg/OWh1JhfJmj1WoQxieAt1cvBWuTmw
8CDt+qdsGUefi3InRR73npYPV402sYdFxFN8Jg6UroIJVNQAA5dlT0w7XT9XKVV5
powVZGc4fWFD4fKG97Vmy+SjTUYh1bm/xO0IMrr7uG6Fx0GJJVOu2eCCZJXOr9fT
Ykik2gxnyhnXwJT/++/JiwV+U+RSf7XUbKq2evbXm+xXAAAkppy2hTF7ec76ov5u
elcz1sDbCYjfTG1ND1fYJ4ei1haLu+6JrwH/qahOHME2w1+6PDlLfeAQ+Ga8WVTn
u16UeusiLgMBrw+H/jvff0GJv+CbGGWZ5Oe0dnO0N4H2K3bnnpuVZPrSBW6nfRdt
qM+FnKIBT/UGdrvfTwGEj2Z12miYusydiAPerFUsVVFBS7/oMpU9UspxoE4zZ30B
JIae66yes9X5gPPRoD4Tqs7ELv0ofsXFigrNpD7WSDjKXh3tGHESl8HivtDbJ24x
3xK9ktlCiU/mUiE7273UKX+txx1yGNcBJSfwDoGdSrI7TtnrLrNxWjVGpfGsHZBe
UL7JIxWSxSydYye+xmMAejROrfUquTdqeqTwqCDDo7H53FNLu3Rj74X7Arox46ON
bYkNekSJmed67rMETGztVhXpjzKPhBkPaFeOoHtKrnK8lQueCkfRRy+tfZ8Z5gEq
J4g9BtYcDce9nX/GXgEEr/sbIeV+ql0n8QBqK28CjrVXP+EcPjeDYd9hzOxo6XPj
1O37Bjh1ux7sWh/pMgU1hgkxjsHQVabcJl89dGTBQN/j1il3zG8OHsLLNKXXFNk4
Er47DciUiypcK/ZI/ck9ex6kH4NGEMFLYYfpgbbuq/UILZCJTBHEN5Hzy3mPziNA
xSi8NnJNZ96hW0/XP0c33zn+Kzcrb/vtw3hSq2ERn97/nBg7XqSDfyO8WusOH83M
/3FM1CiQDb0odMtiIj0iuTAvSncO3MwsDp188x/Pxzr1KNrGQEMvNwLjGWN0JibZ
JhqDchxe0bELMepdtTUm2wBVZlHT7ecyRokowuIBo4BOofn1bH2CTpvmc1+y/XRd
9SsCWgDGoJ5JWfRv7ahGWLWqGWNY2LZMu0Y6ZOKzAW1fJik0RHlqh9OtSjomDSZ3
MhWBidT7BuUWLrbYtl8Q7QiL/bJmBGvaVY4CKl+Gxn/rIGrvdgrGcLbd/4XinaDA
YyA4w1Z0D/a7DdrqfVw1JWsAs0wyheWRHJn5/rEl5xOnxSvpmw1w1BWhWpAWfNl5
IGqBDfhLNH2DyvIPDjqzxew2vuDUAt4PgkJ0lnSlY6v1pBtP/9V/O/Yfost9Wuje
fi9r9X1F1ctOjJpVK4d3X5RcTPdAViDUQQTe6ji1gQ2XbtdYIBz7zKeIcCzhENQn
NdPjtmEdXktIs2tKlA0xBd0MdJPeTqy7EU9Nq8HYFloBZo+hXrfKyOntlfDj5Ne6
H9h0/iuY4snKZH6J0Ed1GX+wIUMjZSKb7b01BNvlSaPHDrTlrFtHJe+sbF7VTQ6u
HXznkof4vknLZr6tWJ7u5/Obky9OWVU/Ul1VgSvPiYKvh/UpETaBnitn6LdvdiQI
6QhSNeRiL1MkenEK/JWN0qDIOy+aumYjvo08KyWM3rUvd6Jr0AYusASW6TmzQiE6
m5uZret22umFuR72u5ti65f04W8cyHV/STyUxz5Y3DZ8rQjRjs3VCsRHyMjHQ+li
4MM+b0MzwBZdT7zFyPWQAvyxyO+c/b4JG+UZJLFu8bfpgIdNnfgKSQRtZ2Mz0VB7
/QURcLzXeLdv0EqFwJP5AKqnibkq2MxU4RqwR8X/0x0r5wXloIESUuF5OgA4tXEp
cpcW24TYI7qJxfKO9epvvHVL2jTR3QqP18YiQxgjki/Ku3cG4GzYNiZFCfYRIQyY
jknE1/TWp0V1AW+bGTfu+LUaH7TtXNN7aaa5UJoIqJ1lUx0zPbRnoko7rD4CcgWR
/O3/SmGBZOrCkio00JgV0+EfF2BgFt14+omUTe+S4gxqHHdAE8LZvxFvZ7ONeJA0
1qyNq6v/3V+6CqS6zbMX780HkSzkqbK4+pEJHDk4ZboXj7OCpbSdqbU9e56oWb0g
lLXJM+sP+a8ubg+knOKhBKD4aBRETmiHuT0H2u59GcXlCzKdRtsTNNUqsj/TMDV9
WA94gXohFcV1HwJFCF1mxt64B+tAlUOwUddbk9wWOWL59zbhTK6nAEGuO5enS7Sv
lENR6AhzdWukil4PkIUroUBJIzBBgmy8cs0mF1lJufMrOWnSeJPdmZzfMoIRS11e
1skZW6tuoONwENJ35fBNmwHRXc0ehSpt18KZybMmvb9NlX01D1q8AD9LiE7KUBqb
Klb+XDi1qfhGake763ay11U9iDSBqIJJAn2CTJQscFjAkAeLeJns+z/HHkKUpfVe
CiKYmDAmsIJKu45YfbpNWMzykmLndDvnF2h0h4iSTLaq5tFegGnp+8hSnVf4XN8L
uWd7kzH3FUnHlDsRZefSA7JhDowZYFTzoZr4sKPj+1CGDQdkopHVs9O9H/783bqP
fhKjGUlp/9PrpOE2oQyc7AFS4SJRTs+vPljEv3ux9lGnveDlNwNPlaHqDz5H++MD
8SKPg1LEjCIwvhMAd/amx8os/NFwup2jX1vj1hz3fco2uzpuAPGHO0vrqGFZGvcJ
7M4YnSTqTjDcOCKqXyC0/F8K95/xmxtz0YHZnEu0gY4eg2Hjd51BRLM5ODGA7G62
bVncECIj/yz9lNzjHu0qTFz8dFijTtoZVg0N7sdqBgFtPi8ZN2l9SvTGc73q1Qo9
JGvgj+1cgbfdBKeJGXOBI0vws4oRgFHI0HdGQO2HqyrDeqpXk9N0Gt7nQIwk6jlh
9S9TkfdeVcHuzfQmodkzewaAeUcaJapvZ/mjtKtihcKdsB3pcqDMC+L9U7iuwjdK
NscnawLrgFLVucDo/Ficugiv6ct8y/6NZW7mul5jfwj2LFpA7Ey1VGWD/X/U0FOH
E+8fyBxQI0DZpU/D2KnpHg4tT1A97prjtol7nRx7YYKRE7c5O/xnveUra0eb4nD9
N0dxwLi/lLm2QJZpXlJxwQUhqfhabg3+CK+gTYHZ69cy43gV2+f83nxM/CvOR2PI
sKab7eEXPgx1sDrH7byNFn0bdj7T9V15q3A238uJkjwr7Wy5JcyCUkm9aX5eIqdj
PNxFkBObqoWoyK9FltWElycVNtv/rTzYmhlGFUwNi0XNgCy9b+QSoDW2f2tppz5Q
c2c8yrgqGc93HPaGmIGi+l93tmhlmS8UHamxMyioEheeUd88J1jmpC+ha0ylQjR5
rqTWYv95jdZ9nTIrRsVm0LFyURybPk7J09AGFIeMZoQCyfw+pPAdSZNMtqwSHZ/Q
UTnAgyovgy2LoNLHdIVojzdtWQVgR90Ve/MM0QKksqnn5yti3Jfv1liE+UjnHBej
JsRBJw7PITYl1korGNfz28CfFk8r2Xp+37LDxFgEQtrvCPgr0eudT8DqjE090/kj
JPXygUAuJoE32cbav3HRiRYgL8Wnfnm40uyzHSqjp5vyzkteOxLr9fCKc3FWbsWy
Qqid605y2uRBVdfzPFpSCtS20xECFedyoxM3/PR8CXMpjbgSm9ufpibz+Pa3J/6/
6Fr1qRCFpDSu8VtjYQKAOLSNYNlLUXAjtjazfbQmANevLxRoX10BtYw41cZpsDXr
NuxY6QuRIQ9/dSjSDF4tA5/km/s8lvp37oAewnxEfjHRsWdCYXOw3kIXb8Csyerr
LQQpbBvvh5QncmJB7Z1KV/BM70uHhHvxQCeKDaEcqyJlejSpGb10RdzU6o1gvFLQ
pHb46AEpdY1YyEfULtXOKx6zpGavsNd/JRFZh5DzvN8A+sey1lNr7phONbNbAhVl
23deQxMJxoGZ0oz1mqRUgHi7ILL4SIwj7VNxaLizdaBIR+3s7gUx9m6utzDyfW3o
xWD9DnIBkgsEYk2/wyGqIKr5QWJTjgA/I3lV7TjAVss9oSiBD9Anw5FDENwDND7b
caqA44cB9zh5S0Ar93CzfgVmloBvkwXZTQOep1A4l/wwyk8OLWs+ov/XFYdSX9kn
YN3pdWKrtC/SvCjHwnTOOAWe7fsYa/HHNUOXlnd4OEkPf2R/OnXiBkIbi6tkucfQ
yw3x9eWARorYN2XtbIvqAysy9EBmKk3Q70yA4LEYJeUH4tPNl+XLvlMCDfVG9u+I
VngjFRRb9OcXQa/fZI3SfWTxytgTgLAmiqc6WT784ifxcNfQ6aSjk6+m7n7gcAC1
+tf1jCeeJOVqGCrIkwHUDlGv9lAJkRtkgEsVk968Sr2zFaZ/cUXkeu4Vw/P5VatH
FB56/T4k3peldmewZXy9Y5iK14UFQp+4qFyXAu0m/s909Ubjjmmc0eub/ht5VvFu
BRgJRpmDRR1NB6VW+aEymq0BvKO9esEFKGWsBCCAoE+Twr7x0mwA5ntqYLXkcvMs
6wmINtmuuyKs9PAXmEw63wFJwHfnazM0EHGPqIQY6tESQXqmucQSdYe/SAp0Bx6p
zBI6B8sd8cuuwKF4J5f08KcuC2Ga0M2gloeZfT9xuDcUelCx5BNDeipz6XHiKhkw
yaukIb3d9Ft9hpr80fp3tf+vvLLxiAfMn5nb35/kY9HPGygCobM++tN0ixZVkE6D
6T/e54ykYaJweoorBs20W9LUD7nRvUYVE/Q6sVELgJFYV6t+ezIMPzVKf1EW6k9w
tn7g6NSBDfXNSx79Jrsi96k+5XGr+YCne2oBpRxOElQWVTJPviEl/JhUz+I1oTcV
QFg9eZgxd8+Aj/M6caFVEUa20ueO/kBb3xScJXGuCKSbnrLWFjNRhY1vpGcrlZ7R
zT3aD5X05njNpUpWs4NCuG0BjzeIgCh34Jls08I0/IKccpgFgOW2Rd5x3EjyJEOe
rPzn3T8tu6Whj9SOFEQ4XXsaJPUn7sAQBpyLd6SXkneBerEeRYnC4IoF3FENei9i
i7VGvucCx7eJ+rKiNkBEfAph3lkYrTl119P3XxdNFkns0BjNcLlFTsuvvJW1Xj86
T7TY12GogrwDTZwZoYq9/RXsh112Y6yluKJe2wLy1U2BerfcYIdMHzMw2WLhl5PD
yuHLcEjRKj/WGLckNoTaBqDEqVPbrzeTXeaP6TNkYWNIqqxVmZVybOw6uabq1Ty0
qZgdjfafB+jBN5nLK8dksVyaA1YbQLFb3FrygC3Pspl7J7CkhDdzDlY0ixYsQ+uN
xyZ6RT61p/CasqBwMYe6amED/h5KeLl6bDGE2oKLUb4nF3RnfILVrVUJEgLE4+yz
Uo6/AlUBpFwlgdh4wDf4mbp0PsIgHJ3MZV0Fp79hn2X2RNfnPkVZ8C+wdKa5ZHnt
imr38SuBV+VZGQWMX2MdbxjMmHZVgCoeM1i+JJiZrFJ1A0jR6864skmdUNDAy5cK
zbgN85vA+Z4XBD0tRd6aCybPVa3Nig9IiykZNx2i0gpPUx6aewOi5uV1ETXigJon
hMCHCGws17QA59SFUw8cLAeXKzzQwyB6CYWEsBXTr34ZDMZ+CFKI4LanOYXYIAqp
gaP1mJwb+2nf5w6pt2wZTLhQEoAecjtY04CK4Bdd89PKhzEIFfDm613mZXkuGyw4
4ZXQPqpvPDrCAGT3Rp9DN/VJl1275SgAIW4tcrUeRi5hyCWKcNCfDuFV+V9G4/Ht
/9isPEiMHcCj01J6CfFgumZl9jMikAKs1WtmX6xjpL2tavTJL4+WssYpSieEcLh3
Yx8lMx9sWm8y3BDeQTocuxL6VlgKNoFbtBeKx0TLtHluUhau55aqcTlOa9jOCH+e
tts5rjm/Ah0T6qTSs4afv+DH7vctKqYfNWCIOdESyaqrC0ah3X4napRJcFOMNmEC
TtNIuroo0tXKzYiRVHsQ1HL59hQrPrnlGlQfNfZmebu64AF5rHaovNVBOZZY0VHR
6L1FepEZp8DUqe4bhCpIEDvUPOSUlDEtTksZea++Fko1UYecJZ79SX2H9Z4/yU7r
sCDMH2+hU6OhfvfeGXzZdrQC97z6/dnmlRoN0VoyA0lEcjr9ksT1sPpjssAKe1AU
WBuCUXOkenNhLEGl365aNrdwjEoqECSE27SKaVhinT2cP4k9Ghk2yQg6yRZr6BtL
8/F9nEOzzFNvbZ26DpE7pQRdMoNppn3S52Kp2pDsP7P2eiCXz42SP0Vfpoii4to4
M4yihWTaON20bKLcDgSitNgrwbHGEKVruea43xcIiHk3IR7Chp8pBZYzI3iqpcYv
n42jj95aedFnXAltV9O4i8TorAGRQbvN/G1XWAK9C5T+JtSeir5Kp2XC6KzI6DZO
eUzSTuysUqTDGpn3ffpxKI7y9ZgpmH4eGIM0Pv0r1p7ttAK17UXO1OMcj7pdHGpR
FXxQFyrGCqzzMMvtlSNbDyy3KckIgjtI6pswwPCecs11KVx2H9ZVOmk9ZnqODGfX
VcdvALzNQsjEMCqQyqzkaG+sgdPlBiUpAkdHSu0Z4KdCWgmg7t+bHojyuWs8E6Pv
1AKF45HPzQEEkQmBWqzx6r2UY52XC3o35pCGb5gifhKtpaHdULRXwocdTv8aEwSL
lSDLzk37QpN8fgT5R15ybgP/uIkkJpEHc5jRNXXHZmXo0B+lO9+o6YedvC3sqWTb
UEQGyOcGtYqYiboQzGOnAjUW6HvKFXGGoVLvxq3y+jcfbW6uO1sf8qhM97t27bPE
PkWXYIy7Z7pNpWnISWx6Poaa2LYzxwvY/kwudvcjZWDFOxtpSOyWVLzELAVo2jgg
Gh/DCR2/65Md1vxze1HoWq2bPm1KDSW9FmyMqUpCk3A+SCPbMHP0tQFZQ6LL9Ewz
Qs/6qMPeESkC2CVHtUwqPuB+S6RTbv6AG/eS0HRKYmGUY1PC84gA9/zyg5+FLpzv
3gOGjOZQPghF2LW0ovK9lyHT8scxTT2Quy/n2aCAdbn6G+0z50BIS2GW8ulcYEJP
tuOAButK7H6hV6rEsyQoOmexqBh0Ibh/6cT2bLIDXE+FT/mWNIKENf+Wfje+vFrh
TdqGtQVSH8mWWFt4SeZ6D4y/savtHCGpzCGvC+agVJGUcmbjfO5HJ1o6dPACT6xI
+5F+iftyzetQ1cNPfS8xeB8AWboGw9Wgf1uWY0mpgKwbcM0VTzRGzcb9PKZDIqGh
mq1VcTEZx55S++qU119woMWYxU8i4GnrzmWrmzMitO2nj/fHDrAN6LfrTGGCyxUt
2X7c5pzzE6hhxfVL6UbRfs5UUSkSIk8c/2yWx42tSPeCDHBV+psxCA1hdy3OOGQv
WKTFMc+PT7LrAmYIblJbS16dSmZXBtj4SNXX9akxic5APmdupBQLajmDn39pFKFv
sTIjbfo0FgIlmaBsQP0DafVwMj615yZAq+bBOgBWF/W1L3mGPaZFhxFGQh20pMoc
2mMzl6TUjx/EmLsb95kFV4aHXLMqcDPQwfu3cNo4zKMkt8ZbVTVGxrfOtTBgUS5n
1SiUoRURJll2jaWQF25SKBUDFvGRU+Vco1CGIClJrhpIEcA8y9fLsaYiVYH+1b3E
xu7nWvDERBiEwX5f6xZYllqBJhVyoYn2gwBtJ9RlEFWF6PqUJUQ/FbPQxPC2UBPf
UZrkk+6YGAdnf5hp6GGIGE4pEk14WEm3AdTV8wsFlzZw6wKRYMdzs+7itxG2oZQg
3eh3ItOFTcY8kJQFxEWcovNUEJE1CU8DDE/2RS2WqdwpKhdWuLefshX6QH0or1bU
panXw0utLb19APd6yVUDj9Z4bDkT6CzjqQnTaqxQPq+0Iywe3BicMW0XTYbvpta1
UaLRIYa9LUxfpxvwzW2mXkZLGhwu87Q9Mki5tCQnWKaGohYtI4FJfajW0CiZZ1gU
9sS+d/SU97OcfVDGCPX/TZ5J8fXirshr4M+w9TitYb14oDezgmuAdQZIWMfOCEdj
ubfcca9choBb4ptR9UCwexcjgReg8TIJ7B7Z0nAU/78ALDhfe9vMt2TnRIocqN8r
XfHXR+9Sc/GKRxiink6ZIeam2I4VVGxmjv3iCM7/cdtfl1/WwOUnK3IXkHLSolJH
VhWJi2YBgVSuFY4wv6+lYuysqEHh9aNwxS6vWlvGc7WSRiMZyZpRd8+Vu/UCLjGo
hwdx3BRrDUOrcDmmX0yIWFGFTRvT/sIbFsKRBVQz2kMjh8oJvqLCOqENpMNZHUeP
gXmAA/FWRfdwjJ62Jzo9OvHQ2bMm/vMSH9sksYQJ4aAEpfIqhO6LpvTQORcsDPAU
qmGqWs24qo75dp4tY9ywXeYWzfl9Be954hBh86qErrUHVAGvR741cMSveQsqGfSB
qnUz8ZTK8FhvhMk6b09pRXdyM7FUYWuGgSrowWuJXn4ML5ECGClyYbweAh6lpyYp
tsAuQKSPu2JTRkPwjf36CiBd4+mcu7FV12QDpR+yzc+K6OSqIVjAhME+rP2N4iiz
Piha8JmFMb9QGiLwwgA8B1DMYZSn+o3YU8dxbLZBC+DPNAiSCdBc9lgOULka07Xt
PInTTOy0drMyAu/VkudbejE20xxrJMF1Lcw8bKYwK54WdQvrOAGQME7XQ01OeGxd
nV4In6v/WNHLrEjosdFucqzFNQspGM9UZ6QcEhC5CqPJzkeFJcOWEgB9JjFMIMvA
TIESWdi3yvC4OW3P/lzX42lkYsUM6G9Uxu85LeLGSBXGTy+ilteBH+hZNQ2mbX0/
gHv7rLyXtlVE3vSl/KFdIzYUss0VJDRPd2BilAqDHDDoEVcLVFtBeNpHvfoiZ6wB
EsiIFx3YwvhYCqWkILIwfF9mvWBWswoBZnTPMDjH0MTwIZEXly3GXVz9xLovB8h2
gDUOERofSaoAxQ6GSJe3DYRG/5YIuf5WO3A5UXvwbrvY4txMUCmWc16BYdlCOAbu
DYTIa788VTnc/luRFKZIP1Neq1nemcQOOY6gJlZ72acSjLPb5XbTecY/cyFPs0P8
RSw8SA1M3u5PZMYmQJFwVi2vQMiukKOqJeRXvlOtblpV01F5IKW5Q3ucL0OORUMd
uQLpAS50BenNERl935p90zH6P8JN9VHvQhqNnC7Ir2euEPUtZ2FXZRcMJUrXfG2X
BtQv+2OhlB+MAKyuYStVC6cYhjJ17t2bS5Q3QQjPbMZgySt58izwi45VGj5GT9ON
GbpnDrvlshhLHDM5Y3HzeO3RQIcD+v/0DzhT043R8iVl9IqJLR7X/hLEOjBy9SJO
7xLaUhxjAmj/Q+QhOIrTkTtoDky5ndWztuey9BxlNBvNbpJj0mWSJ4+XvbzOU4sR
8QUPIpTnZldoXlWPoUeC4VwLcR4TRam7gwReHq3/d+mW7B6XKdwqX1XplN5LXzfx
ovDgOqevdkZR2u6QfkYU8flRpJJZdXwmFi4tWQSgLd68Ml/6WSzx5vl660hx/mXL
xTDf2i/lUFBdiUgwVOusjhCB96rEgh+NEN0i1+zPypTRKzt25N8fzv150JyrqKkH
JJql3N4WhTBfRTQUpnXoxTu2zpS0DDPtChGVSHUOKX1QOwLWj1uuTAVYW9vKlPXD
YD8hrwlb+Oqfsw2dxq4LH4NoC9umJh5ClxU0aRgefe/jp0vED744RXSoEhH6wIPq
xMEsJQCatVJtN5q1bm4z2kQmGYaGU2Y4knb/A7HZlWnUWQ+qjaSSjvSSJIUf+FA6
b7DWQICVRKcT9Mg7ARvKGQ4DctpH2NDVm1zqox0uNWcrk/s1EX6dKBG4T03pjlt6
ibDIv6s1Av47xyIrQyGsNOcQyXU82fKG04Uf+RKuYiHGIsCW/ag0zfZpxwmp0G98
BMeybxSgyZT+3jxKxHym6kA199XxKAmChuWXLeye2aWs6uahcBurULxhPlVowApM
GsONpSJwzWTpMUPwgLohANnMXrLRapGAGvreoFqJ8RRlysSMqsiBDU0MdE/dd9RF
zs4B59MkAbh7NAM93fe8ua+lKYsGQmywj/G1lMaLTf9zlFx6NQ5lFL8pwx/i3BpD
S1arC7dKVN1iYz2rLlpzdTkJdnlsd2Xk9NFa8NIHmr+wxGm45+pFh+fiyiaPtZTj
1/haPP3RUNJbZAc2mpk/STyEUoBqn/dSuNVVOh2GAk7eHF3fY1WGCtxWUTA2JSvs
+m7a0/oOmy9uyF+eQb9clwp6K8YugzBEHpbhfvEQQs67Hsifemu55WFyZJ8ExCFy
qwNfo+YyHcIrzrxfK8715ol63UduFZwnb6cwiuZOe4mTLKfYp8Es3PXYRtJfL0UO
7DFOkPobLecRg6Yf+1wJc3QTbMbSpVdjk+NjArNPlzfmyMB/u1yOLeTmiWJgujpG
mT+VrcVQkBH1H+iaJZj/bs1tdOe8YVyzAqE9iBkuhJzx3iWUW8iWsIHrYjed6C5r
8XMzRMW+22E0KqRhf97a6foUQe8yHkBlaGvUDJkW2MQt2fjJMB6TcSQ2CWSO+e6F
7TGGh0SVGMsVlIhywBEDJrxp6PyQyXH2P0k9BhfxBiPSN8WedetZAjxRuVZc52jo
W7pLCi587bDblyzo9LLpnkPCusHo79GmF+y53aVAQ2EGTjoHuBxInvX0lfjQWATX
e3E8vl1TDeE+tzvEQH1kIulmHG5bni3RWCOME9nAvZmli8Hs1GWZF0iEkWjGHT2X
XfE8NsnVCyK9Z3fWPyfS3pag0JM8Fa/xbgo2WNJS9MnYeZuP9UVOk7Yq6Q6Rm128
XCr4V8tFTesO6hSV+pX372uLypzXmVFOJe9AsHE2LGvAqWMq4nicmiDdk0NpP4WC
FlSlphVcDm4sOFpmB0hknb2RayTyx75bZ9JCgO8nPPsMNymxWTtTrg1vOoRPNQNu
A+cvPmxEApKsw70UUZHvFZV81dRUahiEpDsf0b6mX85T5+XB53dirAyi7HLBjQ18
Vz2SrEWQfZq2rNKnIwCVeNET4CLxr91nqKTGw+OxZ+wEKTjb3SqI8IKjT2qs+SUZ
0fQ0lpRbdtk388WJ/q7K2Ciq1B+zKrfNMQdESXaDQNqwtMIPOLaFxCm4BW5PaNwR
ecazcngL3GPcsi6dyka8x4my7HcD7Nxr2bzsUP9Rdt6/HsSY+RRSy6cqrnvDjDxw
hVY5Zmmw5CRczV1Fl14ytZqgS3eLPSIub1TJ+rEQBOoeWqIkT4MY1hXZj44u5oaY
wjZ7hIkbRhw4t/C3zC+/jGvh8IxPux0bW4wouT/vzv1VXrU3ynJ53eheMXsk0ynr
Bzb5rlitesnJJu6Ygo1OYU9OppraRTkDsVXzMPppY4eTg6qQsD/fhk4AAYmMirKE
4X6xjkc0vbadDijPthRrHnGv8CJ3UEWjHfncB4KxRRpniZwxKUyYGQmDE+mUDQ+2
fFVvhuSemwc5io8JSiP3TEKP1+U7LsPH4OgP5BpgY+t4a3IGjWgjloai2JRYe6jc
/8/gJFp1w2CCAD9mvs9/wqL8SCvbzCm8L8c2qiXPaYB/7DNxyCJ0AW3RHtlZ1eHZ
sg/iyOy6Yh7jWF0u+h6bVM66BBsClL9cY0r4ozwu9Bon7QCFhUoh7yl4RA70AtYW
5A/vpLxsqtqEllRzX3aPAzG436FRP/oaj65LZRIqJU79vdsXcdmfdVjZZ640gtAC
Yxij55koucac4tpO8unV+1VmAk2aGQ4Vr3c0CoNZzIve5rwuwocb0bzw2usGbRUQ
fxqEbjZqK2+9EY00DYZ8Oc7cmTT2wKXFNZ2WUbHRf9cU1RVfT8x5ATEoM6NtVRVf
67f0oEh+pGL6AREj/x6xmH7kggP1Ofw5dVXUef0GhCmyCxs4UPgxDPlac++KEwPo
RmPvgilp8uBDV0Ub5Ivlh9Tdc5iIoJY6T3MVRvoX8A9DFjg9zJRSU81I+vDZul9J
y/BVwprfy4a24RqtjAMXato2XHGpwaKUs5l8Ddd1L44GteDiJQZv6O85HtSTKbkW
swexORudX3PWSmBkBX0Q/TwDFFKPTWSiou/xjJVeSAzthJ2EIShtw98/Zl5Vm6Ty
K9HCSjzDsNX94Tr/BaWn2HgcGSAxX/FO4jtbSLHH8aw95yBkCQ1e69wO6k0WBggz
Lk7d9mJN86Qsu8Hm/Vwaa0NBi4o4fJnZJQJN4+FhPpGkstdR0iXcYyjA78lXua2j
Lgm3mFtCfX/KzdkmTiHwSyviX0HUJ5JuBjGO/XmChmTL/aKjUtifO9lXkeP3omzY
r8Y/GBx21bKT2uDlxymL5vdzLKIum3j1O0yUpyIULGtZYN8YI/MkbC4C+ScoyvO8
DBrfPzdAzyDy1p7Z8LhvatvWiZkeqkFV5AslTuZqrtoLjRgyEdAK08lVjJiXBVli
YNFwwtRJcFTLgN9IMyd34Ap9xzZoPhseN68x15TSHWj5t3iKjbbMwK41QukoBaI2
2pVQ/2dhufozv9CeoQyhrfaC1s/DF8cc3KYIAUYuXsMZdpJzj6CDwAJovsC+3GTX
dtDzy1YynFIIkI4oAl//+A9aD1MyCqpRbud2Wu9sYbMqZtFF9UcLJsXVtwBKyObA
FuojqGQu6bniMkLbRoaGNx01gzCS9FI6A5vKQRiFzCLAgbXwiF4cELpdn+DYHygx
4X7eipPjKHRsW8/g2l/wjb2U72epK641Z6ThZmBAg4sQGyiAEiLklGZQ+0kAuNCg
Gd5eqOCti1/+vPCW7luPP/h07bSZI2kRdJey87Ta+gPJhdbxbgqUCIGBZi3/1Lox
LGLr9kjTL67PPY03zuLd9McORXxoMK+gjz1c6NtoBuB7DDR8rrePGy+Vxe+9ju7d
pKPr/2ZWeDesX91haD2IbBPm1lW3NOKY4GwaVQqLSWEtS3Hfc0XBI2CHSsYzDSvm
1CoEY19HhIB27PiocL2rZmnqQhUEW8AVi1UN6UVQJOOzaJ0nztrDoqQnbbAFFoSw
YOx42LyYojYVNcQH928bOpw4Z8z3Qn3I40KngqTO7gvNZ3NVoy9aFiiwRnBH8Fg0
HWQCEqxNho/rW7aP6Jlc07u+P+tHOzMJh5ojWDuaN4MkRKRZkPQCX6EUTkX/Uzl1
03jg2XjF2NzcnoaLZ014PvvRveP7ix8YhUQklydQ3anS7qAhzb1dRa8B2n3mkZBG
hVUDgJZx1KzftqigsqtzV7EYsUTt+bOEtHev5iL/Y28Q9fPziX8h2F2ROWimBtsF
ByC0lcbpX8PgBUr18/YqW4Iz0uBDOlWDmQGAAPqLBl+UZC6cey4F7g+O0+xETF06
LOI/pcoJh1uhCRv0M+GNwgFlIBgOlJrGjxhLLKgwEtlvPWcIORo0/JpB7N1RcwX7
SGBzLO5coXiyBGfRFXvQad77JdZuXpqP5WvhGBK/TVEDUzBzTykEyC+y9MPpWjiI
XEA+RpJjtrlnIbfmcOvy6VSXAY2W5isJ9Tc+BsWxeO8w8Cj1CF+hEOe5BHLi/5Lq
rKAKN2SjeA7xUs3vmtP0XYZilYGcCLtqbvZXBjFl7AMt0ITLAP95IPHvUrRmycvW
x7XT88H/N8BK46BRRWyUURoRK3aPgoUJKKbQjO7zV1mqzj5Pj8PS3toRh+SzOl3O
ohKIxIIjDoTVC+G9kJtWv2nYWwovw45PSH+Oua6biBCs8AzojmzfwyNDd0F67mto
ZWwlK06aMStcumIo3lBOyS8GxbD4JJ5V4lIgBaypMg1g5VjvpwgjU5Taf1hd96tH
wbtC7P4FAfMp77s5r//dof88ulT481noLdcLDzVaVD5B+tsZm4fc/JMO8QbCjY5N
Z6/wwbPtdh37Ll9qUJLlqHPgBunS35um7q1m+Se/iW08jYHOiJn5zJWsf679SSen
vShxs7hKFVgp2SOf/V44Fwlk795ix0thc4ic8XfXfIAM+81NK5iFDJzJ+2Np9nUt
s5SlF0VaPfTdQ0auB7JXBDPOEYAtF9kLsTM2GoK8Z7PwzThKqKcWs2cLuIshS4BE
C3ZTtbSYEK9AmhvTyJsi/73zMq+e7BiVh6LWlfDK7Z6aEvE2bFnyAXXvxR7eL5kN
OxPJwtV43DZ+i+Q5QKiJZiTf3TZ6hMlwbC4YHgSBXM9X4T2oQobGVeLm7O3xyEDJ
HRwQTje6MQh8vDmsKcXl7tzup4nyPngOJ226NNhEBJDX9Kenp56og/ERWAN4qy4J
OFgpxPRmY1ucwUnEMjwj+lkdgJ91FjoKXXBNyRfsNHQF+2+gfDRf/Q8PtbAlOhPa
phuw1SEMGysJHWyA1mB7GXdY3clZtAd95XWHpsmeX2YmAcZLaRdILzFt2fNeWcHX
6CRkAqD408BRbseKp2FEO9NweMXS8GEUu01ZH5MlfjKBn1NzkUqpEbtirvG6e4M9
5CF3/t1WfDY/lNiAY4btX/s9Vfp38GExSlAAYg3R3FWGaFyHgToVjNmup7iIAaf8
xEnsFa7Tq0SMKMfMYpl7ActolgvQc5Cb+lBoElTM1DHd7KiQumdVZKjBCLnFY9fD
u6JN8VrsguIDBm/ZwLX1eZE+hSFwUWfQQiCzW3R6XfNrvCmA3jRhaXU48ZAr+bvB
jqmKVflytJg/KTruW6grFBQMlEljZgucsoof3GqzaKqyTgZ4jZKoxtl5WVApnkNw
pZn3rT1HQN/3sLEnjCdCo6/32hUsJS6ghWAo6gvtcuIraPDVTomGBKCUvZnrV6vL
HPmkZEhMS9YAL6aso8vwjjKQJ6Q3IVrw6lgXxIvv0qcZ7xUo6I4sd3vZ43anzUOo
Fe3rxf7FeyDJHL0qhBaMrAd91nCk6Zg3ViYN3YPdJNbbtwAI3/KB0wWfXnDOvOsr
NaK9JtIH9RoPO/zK563KsP7iUlfbvYVv3QlIbph8zvnGtfWaMyIXH/HmK7ch+VGv
7bwu2bMnsu+BO57adJPrn42ydiFAJxt43Mrfyoy0Wa++/UedP2sbGeBKT1vN+hwo
eLh+rHYtGQ3lFMfiJo+7kkHVAiUXv5HL/9DkEtTRT77zwQyAa20SC+oD1aCeiRet
oDvfM7S4T07Fvn9PL1FqZicGChU1T5CmAt2+PGDlVJG7f+pu7HUKTqvaQEyZYddV
l8R16hJsTvPfAb+d2AdK6/AQHgnIQUpwvKdy0uF6jRXCH+NoAlTJU2xhGUVLFugX
SMYjYnb0+P8zoMZU4vMMn5wuVHlPGAdaxMTHuDjnybkfkYZFDYR5GAwgCyl2DxLO
eWL3rkr+cjO1EmQZnEsI6cKAHsFdppVNIV3baghG4WJUzjLEbeDfNzCMQRxF5R7t
Kz7ANOpz1DW2+KwBaJlge32WHVYqiq1NhADsC92R6vhMQ29z9czCHpv1aHsXvg5o
Aq5ze3fvyR7V7yE7AkXccSPviIYcKGPDPl7BSiwEVuYrwZFu307yBJHebo30tv1Y
gRuvN0Cg/4huExy9lF8X4+qQUVIBVOOd3eXN5Gs8CA0W/vStOriwKtzH59S71N4O
+8lp0cSDtl+k3PgMqCk5yyEfhCMXA+wGpuvb4Hg7R8FhzgbLHiksQhdlgt10yTyV
1uEvazV6vfrD6KC6TRTPmVZCNE3j2J0sB11DdUiAmyvNrh9U8Ts26YDHJvF++pCP
HCFKB3A8RgMF5frV5q82/IjAAy1Hznm69EjQcO7Qf2bl044d5RpU9gl+t8DoFpyo
Z3TQJ7qzMkB90JmhVwnTlfz7Bz7s96y6MpsNaTzrZO7TAmBIxmgCgExOdWbRu/M9
t3Yc+LMrD6ht/7N3PKZKy/U6UcN46FAeK0hZH9CgvdZ8WzwBJ5YMWSBaPXfyJDFq
GU0/P47wKXpgG97dmVGnw91dRdK0Xx1lkgGWua0ckfp47P0qXRrhEXZq0KfQdD8T
PgPJTdxVSEKOYPgI+/wMdke+7/ytbnOTYZjoC6hsNVXR4w1JyqSk/qpdCN7AdmT6
tPlOWpg+Rvg0Yy6CA9sfr2SlIJGUMU8kREapTA48mw8wRufU196WxfP09YqlqnkO
Ovm+zU8DRLgmy2LJ8ZmORQYRJe/jq3P5yDniDpD6hX3Bba6EyBl0BHWSyS2mHffV
JijuB8GuCv7N959sjKPVDusvImx7WYpF1Taeoq77Y0lBmZoYkJKVbFYBPNwCZ+iv
p2IXQY3dQWL1Sk7/16XQrQy++N3yu3Hu3FCdCGXikbwyKJWlLew1K6uBMMnWuW6U
boogPAHzE0j8WyVDUA7alo8ETKY/lBnwM372YmK/hGMAXDc6QxGg9ELu4ALOde9v
8mcHTEWFjKfBA3OvpV1YNnRiT9k//nyRF56mYAkXTHEBjJ8fwTMm9FRJa7ifmpPZ
HPzSae4QHwkbuDI/cibAS5d7H9Dop2vTBAUhY2n0sPldflrOmCfI6CpEd/SD6I6b
oFJKbvVvwsDni/iKRPSkzG3tpRG2PpRLZyEeV49UaKL6qt521KRHk9Ece6cXGNsX
FoTFgita+GsA1uu0SEZWb3Z1p0tzW6pzrMQ5N5rl4VJVz8XPHo5zdo7hqC6jjykM
AR39r+DCu/yfsIUPlItahQx5ovCTgZ/HlM8wsFsa5vHrENcl/xwsUvjF9QjnH7LI
0rDz3S6CY9+uAVIfEMoEold529JbhDbIHZY750H8hlDeyBq1eQAfQstZkbPs5Hpb
Mm8RzRQlqvOGAdI+8VsFC38tvIJDpwy1EvRqlTqHS7QmKBM3uqZi2vXu78IoKWOx
pbRmHpgGEnrldmBPcOA17Y7Q7mXk/ceFoZE3yhgYx8rS6jVJ5U4dDy6Gvw5FEH1J
2l6N8Bheqhv0dZRYVNRugCOc8If7ufoZ8FHmulXDswITWRWPdESRfulI+bTLjtzz
tvL+WcQR6Iyga1cJ4H7fEhrfrIZJ2RxnNWERAimOh4zVi9h7vda6eY9vLgY6r4C2
Q6B7JMEyhuf+TuhHAFop795DvxzvG7Y5DVbtvFZ9xCxGD0vaeOC1GXYXVHQ+/uzE
DAnEGeY0D6+RH4cd6S455sKDm8FWOZbBX/T1ld+H8PC4RizNRFlhkf2ngOJwtOnj
Dp6HXGXmIYuXAPpIsWju2KMd/x+RlpdbfeMQso7XBm5vbI9Fa3/LyeJ73Zpbve7G
DD7G6MYYw6F35AlKKpMv7hN8QoACihH1QlqvED96GZ/S/E1E6fV2yQPPzJVDW1ZB
eMbhAm44t1JAnPZrQxbMNuKcrjDVk6G3JgTudOBeNgcAHIDeVEKySdZnVUaLMfR/
WFKqqEY99rEzNvBav+IYS/RDr4T/FaiBJG20sDBB4Ds43+zMwwY2I/FpeORi4SKc
lvi4BNdCW3nqytImS+v7P2V7T4B+FELEf2MVeFGDsh/ZZiEhZ8ge+tmvBFJLMLFX
E4hFLZxTL3OcYZTCQIznLcun9ZgnNQLKaaTcA+APVfsTk+IMOOxfYkP+9dtCPp1U
xghRu8ovV9MjnPcj/UAI2pmUj8/VPCSuBt5o0z0jGzRZIrBlerPGOzSPzWbjc5QU
SivqjBsenuLrZsCTDBV5suOlXdaa3tBuaMIXzs3J11sNZuOC7M8CRChLuUEBYNii
Eq+Mj6fY1+lE08t8Tbf0LRdDEt/aUV5L3/XuwXmuq0Dxc+hSjtgArmw+XRCONV+W
0CdCx/3f1bprenG/ZfdHkC12uUFCbsOaWxAt5Oud3tYssumtPJeBhtCL+KtkNdqJ
trzzPLAPAGvckehA+6xBi7WGEDAj4sRh363OTgt55KB4SHNmuFC+CEhdR1HW9aLF
0OG31TKcoDY4kAw1ImWYaErPtOSJtPzTSqKJ/geL7pkZlomBSgjUhereXnuer9E8
2QiFAN9AKZ9p9bJDDLMkCKTTNp0ASvRDqFpKSxRz0mmmS5gcRve+0lqT535MA/ti
SH7swkrnOPmI223Vt//ZCVu2rskQSGk+QWaqlACKzFaLFDnVwXl3eljQXTyA9Dtf
ooi2NRoPtakXMr6bUV0K5P0M94MhwkHJa9BCWplSp00GTiGW7TVPVfUzmP9vgAHr
LDMLTFIkq7amw4ItnoGxVzfNJNqaxfv6xCRpx/lL5S5+tviRo2nQ/Yqg3rZz/Zse
zRfSLF+sQ92L8tjX8kacHAlkAqhvqSnBOVPON5cpyNS9+UMCyyGef6av7NtF23Ci
8jLAQuCodKr28RV/MY928jHdF6aR2G8Ga3e/MHgZLWMHK/2pnUByAi4U/r5lLWCT
9rTjsBvVVnlSLuTLNQ/ZoCyNo9Hovu1M7J3Y/KZiDmjm/A42cM8n9JG8d2teqWwb
h/9RqUuV7AImdIxqTYzSaawulg4Hx7uROLP9J+HNkvAxY2ehXLfqWIYUD/Pb9LGb
I4uj0AWTfFva40IZhf88njLg3xCH/CIdLM9WLLvFj9IaLh/tsYwY41uqmhe83GdL
1nL17hXjFGLfpLDBZWDScRWNmJdnpIrl28qQ0PzTV5/iDGZr0wbSA6Irc9idUUuk
erYfO/4+IjJGHrRQsaeU7ODkMT9ZFuoBBmYH8D12B+rq51IISlEy38ynA0nnptQg
q0o2I9ALMcaGJ1biRDUNUg3ND2+ZecrJrHyYfAkGoBgTt0+S99CA/QP1fBaApftd
29ETP4HmoOl0fiNJdjliWLGuVznVvC8b6otUFWPIA7Ym7eikTbGPZepGmY24isAD
94IIQZKCDt6RcR3a32pxEiQ8tSozsFrGHqazIZdhLidr2lq5cGgPalwbbQFaD9Bw
tQn0uFZl6+mt1ps5TCQZ5JMoOvwHgRyAuYuSnFa4FOKQg567SzQPQDHM/vDEqiz+
8F604l23HGFC5pxx0c2OgheAxYqoiXehrwJ/OpE6Gvo/ZmO3Jpo76xrxGIlKPqcB
9ecPqoYWKXsdot2uFTu1pWpuTtMng6MBarDuz18HlKzxY5O4KWATnCGMlp3shrD6
UkMrbSswqHNEO4TH0sdxSedsAkoCx2hR9dLgUn4Nr+QII+a3bh5eLeWPy9HadJFj
9kgZF9NgcLfkWgk5B1yqZwqpbQAdmOHx045W8JJaWPGoumeBcQkT2LfyV2TEoiT9
SP8stH+167N5kRSAEVnJdTjRLzneT/6uxevKdHIRwXrjeMtyss1WKQPBogLUHSqF
qWN0954Wa2YXKf9jzwMHmmI6lRhEgcxUdInPM0/RXCnRvNRF4ZOt/5Bp059G6Df9
0ykMjNj0GJpcMizE17ApjbwRtLhsfggy9JfMgJ/pY2ug27aDl724VEmyP1Gzdj5C
VITP9uI9mDas9Yu+ttu5f9cQLsxGzVAFdNO7a1N0qhN3o8QyaeGqQv9z+TYaErqC
1Rp8GZO80bwQ64gakjeA+GwfiB9fjZXEPJKcR9yHP9q7lj3M2Y1sFwsX4xTpEE19
mzxtJSgvs6vaIj/ZBxIRayQg8c0GLmR9SPCiAczZ1e0CmGGiNDfPNRWgZrB6AfVZ
0Re7ZmMmPtaHo0CHHjVQEELYZKK8QyD7mooCfXiBn7+HrtG+PLFfPyf8fWd2XZEs
jaOqslrMstibGJiZE2G9VvXlWusdiG9QZ6I/NDgtZt4nNoacBK8m2ypOoVFhjMc1
0PTtEV4/qXrDlumDJFkW9OJVg0uSUolGwA5qdMjkDogkw6jFAsaFAKhUjQor6Gjf
78CiKaMPudN4M96uOYAE76ROIOsa/pM2apqqZM3tWg4M+T7wJedz4jy00Rs4fc+j
tLC5Cv9oDGUBYEjQ6ZNvyIKBq/JDhAl6nrIISbS3H3A0vL4cq7mXzhbc/rWa2YEp
tb0Q0F1yoq0D1XeTt7lY5R6laH+9O4x8gLuaxm7+d8Tql+c36cCgCC7sY7GjYVmO
oqhD8Or2q6qhO8HylsiHpFBHsHIrkcHqMXX7b/Xagsp0Ugsv1YGW91jpbuJLDu+9
3bztHL+7IrLjn0acq2Jo+MSCeQaxUVj6nWdHBpcH5+ii/QZy9iLhDedwiitEpFFq
SOMG1tU1m1rkl3eh1l94y19DCZ7yKQx5PtcQk340JA5WsvLJJXyWrRRCVz31PlTa
DAcmmKPN1tWMTvGb93zUuuebUgeDYgfXv2W+TOGj8fWfmSYMY+VI/aErUfKn+y10
6PKUZgEma735ifV9EmxG1pgV9yZCGNgNT1eLnvuMetZuHN1Jvz97YjcR+CY2bGHu
QPb6L38L+umeDRi6O5XUAQBmczLWywZdUz5Z7dZrThn5VxA8ORjTIMo80ly4jYRb
1iCE8HpWDrehv0kDMMHzYLFTnfO9AOMT14qXWiIqQi4Kf1nXROyFyqU4Lwnaiy7Y
zSYIH1no1bl5B9uZ23v46KnxBWRU7rf4WKSUuxrNMfzxyQUCfeurhfXGF3JFaRSU
Rd6Dy8SH6ePiNTXdov7XdljUtXaNhyqBDEjBoKO8yWNRDdQnxlmGZimWzLQ14/hn
70r7ho3or7FyEVKFvd3AzK+2PZ9c+JLofNgdnfs/YgfGWu2BhYSDrJKwMzbhHPCB
a3fjQ+ZMxeURvEllCxNJz8Yl79MptuixJtIB9L0VcgX/YCoVeLOcK86In9zgx01R
fiUfByA1oDYaE1chEfNCdfXYaGeED1SaSuQo7gU9EyjQwx/D36lrIIdJvphPasEv
4g2ayoACQ80u+OQN03T76pYaRLeeDNH3etIUQminb4na2KCCAcRo3P7yESITwstT
78VMoz5vsx9SeLxdPKhFqDvvRPB8xEe10vgxcbgic+dE/OtKmmmJ77a+qF0BD/T3
vlyimtLpAh24n89NtrjM6EidKkuyb6vir79nel9WFtfbuyCvlN8e9PFzDP6tYCJg
embYbV2y/GoQQfN28X0Y0AvMeIA7y77ABbGljv7dMGMPF4mu5Olxh60scmThqr0W
Rj69JCq2OTiaplbzCkXSXKAxfeZEHyGCEchuNHJSxQFcfFWmWOeCrCH7vgQMedkC
m9IHH1qQF+e6KJ7M57NeWYNTJW+Rxul0TIxhm5hqHakKQxACQKG7R4Nq68yjZuxR
z+WlMAbFqof4nbjlO85O7t0HWuq8uItgpjJAgp/n+BWk4aaaz1XMv7ypebisAhEn
bsH1gpibVrHCmEtGjTUJiFSDKjKvpPfqIKdmcJYAEZtb0LYvBPozT/SQZ58Xj1Ge
4P0vpbVtjF8a1ZKK3INiOWxW1DKmWIkua30sY0dm5kL44kqhoC0sIO55gtkauvzA
FYlYriniGgQqIjlH3m4YgBEXmbFE1bqzSlHxkErPaFki+PdRc/JIW8Yi8F7MzanP
NRNyN4xSvDt8ZaLV5nITJVw/LDYHcRPUwMcD6vrYoAZxdAzW2pWrcSKY9Qx75tNB
2KG+oeXpQDtYDdfyVudTvMT/xMh9XTn6JqdhySnX07Dyalj2COv4QgFAnYDfaTW0
NuBEfLw1qt4QUbquA4dEA7N50aBqREmDj4oifjCJ95CUzlF2MioBRq59ufOGfkfq
GrWKphzUquBt/8o1e4A04ZvH0u8BwqnwxnA1rZLUu+2hrR5+DDBZ/Lq6HrwzAXZj
vBeW/ZvdcyHx2eqLEx++ersaJgsMIFC3EIOfQRHLGer+sUN3s0TR2e/34EkbzKcM
0jvkAUDItMcRCRajmXmljfYVYgP068lL9MJXQ5E3y26Og5/fJIInrlQxa6GxHK4s
vBEZZCSQJnG3xVKJ35NPTAME83ilIAqU3V+kuXP2y6N+yqbQaKY2m83PNRjnDFUG
sTeNNPFUslFMbeHtWX4s6zETAlEYu9vgpRIqSZAachwNZXoLNPYk8YThDyQq+6cp
Al+K3p+QU4NF2qvA6+5EMyIMcHwdsnXPxpOb/vMZY3I2YF56boTQfQj60CAErt7g
jqz5FfIOAIRi3XG47Axxs0TEhpqbN8kMhe7ruSAPlLfk5Lm684UvpVpxXCTRvjJw
ami7axgukyTymFQxx+7OEFc8WiCgFJaKZ+UUL9hN7sZ8cK8FWxvUCFw86VYzMlQg
Of1Prb6XfZp1yXLTpNXC7KWw4zQybn1yZc9MXJOm4un+x/EGNACGV8NWkEuoPp5V
P/x1i7CGM7+F9on7HjGQiWKPe6ReaRNEHJct/RiABRHqTKfNqlAa2kDAbTIBcTi3
wsQB5/WUsqu7+/5vPkMfcejrBhD+9L8vY5A+MR/JJGSuFjp21fQfwA7KoBTsZPFm
p90RS6FC48bD1EsVuJMWveBktPlRmKk9HCPmfN269VIGoRo45F3dXQ11ibEA9hiX
ZDwT/cTybJUsMSsCuJTrHL4nBQ/gk5nkmpfTx7vedhZHfRuCFtj8QfW4E0eGPGGN
d2j9Sd0EBaW0yFlHj28kRFUK0BWRPT3jF/dRtD3h/Pu/7MyjwjCSTDoUhbkhFcaS
t7W9HMIHzBVp0x810C5ZEfm7ncXz6HIEMpGu0hqDBMx+0qpdmpRL5hz1X8maOnPY
aavRf+VD4j1S9VdajZiphRdQ9MaAlv6H86HeaFj3OCF4tCCRVR53WA13V5m5qiaV
U1Hn1LQbpg5+46yG1DrDKHPBrbOjdFTdPQGZiXr6slCmYZXcmqPjoWqwCAh2BLlx
xacoASerVoivvQqkC3O44GOwmxyde+aAqeM7e8CtkwQsZ3BjP2I1BpiUUg6V2NBj
3BXAbySABETirRbpKIL33Xu0Nm3CgczLz/2r+fpO4ZoWOYi4yW8VnZmDkiWBRkjU
ou5eIBdsJNTzfrMGga+V1m5HuARtjSb4f50UXk/p0pxXzmgV82MfcaxEc/8eYeBJ
2X88ya83jBWguHdbywYdYmNfPO2aNERnztg4fFHeSyUvGkY7Ps38VeekT/S+M7Lg
6Z6BhOAvIxpgdEoaqxywt8kKi9yk4DktIj2x0KIz3fl/c0w2JH+QmsCym4uS6Ubq
TDJ5s0m2JdhSjdG+HVsvPoMnUefDnNhWO2BLo6nw0LDCYX+WMAxTv0eEDGxu8cWz
RRb62vv26YMKdltUq2AiqMT8ZFF+3jVNA/rTLusVfGfmYL9FJyahb2u76oG02mSq
YPrOnOxt4KkoCGduodNVE6psajuCb5owNLbPR2us5uQDlhZl+oThxyyOBvYqAOVX
VbG4tyUG3PnHCk0S9OLIygWk19Z8DIC3I7nylV4tcswixkUVraDYt4B8ZFyjVBIU
kx57tzutxOl5ktUktA7JX29wDZtV9h6lApcXfYqFfCx42K3x28iWkTkbcjLz7Ukk
OLA3qtpJuQ1P3enY2RBzWgMhYjhWyMjssENgSRet3EHvXRu5GB7yD2uKC3koEkI3
DcskKRRS27SW+74nHM2uoylohEwH5IDh2AzvjSCp7LjWfipi0BEQ0Vnsl3LOKJYD
AdUhlbQNHjVJwweL/PRqWcjBgsHnF9V41uqfNysh9VmSet5en25LS6wDnQlcuW27
wWeIAQTlQawQGg87x+AWiz46rfU7klyWnDu0fmvFTYIZr1UhVTkb1QF8AaQ/Vkk7
7bqw6TsTUIDInTa/6hraCZMeh9qkBPCKCQMNoQfQl4w5B8EHk++jESUhWhWo8nnB
h8FCkZ93D78tuso1ZdVehhBbyGfdvJ3Uw4h9AUE8pXlt6SbuH2m1LgppZd06dNka
+WJhh7MgDvaZxwxFEAb6r63RJxiiwk2gixcg/+FZ+uWLIW0WfCX+/yPTOGwlRQ8t
B3yxnjpvp1SoTzfko+aKteQyrHk1MnN7qvGNYv2XYrGI0gXA0CmWXgMl94iYHgaH
jD85zSxkI+j+4w3FHdOctYGliARxpDzqKCuZQBfbqInZxNqKoOZUyQW0aucva8xe
d+jHxI5lhg71jckdPJ2gbX+oIpTVDXELrEI8DkNkgNMIi3EFKu69mSfs/Yy7kTH2
MZZjLS/z1TBcwkN0FdAkV7VYvWl7+2ZSc892aG9lP4z4MqJ1Yz1qqGzc6+6WxIVn
lhhuqQNvbtxfg+E++w/6h8C7CyUEXZSk7fNZzBSk8m4bD4s0JWRlKllB37zsA/4o
icZm3LmgxOjHUdzHVLzz5v2x5HGef9BlAO4/MvS1+Hj2GZs0zWjq8UbqeKB8Hrtk
Q53dd6bWAFe79WmdfQzGyBOI0gHBQ1/E89imEe3j8R+x8ciMVNrV3puW4RsxC48T
OzZzNq1Zsc024zFDU7RJHGMTd3M5PuQXI5NgQX8hu2yrKSp4grjKj+6cJL+bYF8l
wfsEVQy7783yHGdFaitHVZ4cTsjk0a0u1HFllnS0H5EZnJ4tlNge7I3YjDZzAB9I
M2kmnNRDB4uBn7jjFRRG8nBJqt2uRHtb9dMm9U4YAm6HtmfNFbg0BhghWW193lQf
1JAJmNIcUCAdVD12X0dYiwn0baqNEZ7oMMinzB+EpGd3nR80HJK5z4+bEsG6X72Z
m2hUVBw2OOCUwtHabzWV+qZYqbpVm8jF9hiCfXxs1uiEWQFDPOETBMqruILG9zRP
nxf4a7QYBX+H3887xlKP53K9TtxndUNqmF3253JOxkFH7le9Qrhu9+gIpnow0q2L
9GO9OyzC9XuX2yzKblryp6XbGOcb0SFN93TaQ9buN8f230HXLnQAU9sSggHU2UxE
6aWWqG6j6fGq5nMFJXPscKHfXOhrIPkj3xODTmXEWphquVlVg6iYZTYzLtoWtkRx
6GnrNEV9E3kiSpn+CQKKm1wlYwcYtDzErRQCddCf0UekzQT/AYbPUJCdjiS6pRHM
87UuuoXTNcRMCLQPfJx2PPDJdiuXF/RjPcfcVRELa0+PNhtlfae204acOldVSnS0
mqLtZQ6ZiO87QJcYo1ROLHMMywH0cKNFis74E3x0riraECz8O/loPcqboIalJPtx
HHrGWNWqbmhasl6kOSlaHIdVnHFYmr/xur267lAzFaC8kT7OM1sLvq6H39dTqBkD
69BPhgo4++x6Ln/QMVvU1xoGv2As1/gydiySCo5wVdWqkHay0djk2KgN/3QMhwsE
t7l38JWwQdNxbLLQX4cN+t3UeuQKr7zxPnO5gW8CnJdUFSDgE86rwLTkLtys2Blo
BnJKOD9mTnMmiRnqg6j2yqEe0R4qCaGd11NZ6OrDmcvpzC+Qm+ITqs/I3epI1OlV
FuRtsHxC0IIsfZI2uQQuHKChJsxyb6azVQ9YlSpKDsjWYwhsK24RXrvXDiBOjicu
eoRE9n0Eal6WZ+/HjErXApyxYEwUV/24CATR2/pHZ9ANsJGXvyNr80FjTHoeqzkg
x81jiyQ792IO3rLtihbZbaLDvFVWYp8fUG9hZnmbNlDalLdDqqAbtGEO/T0+1H1O
iiBRwNdeTthmlW/evoJEDhvoSaX1200J52vm0dpmGMijXrvWiVTr4nTiN+mmetf/
drAMJNG9DMu7/HTzrsRk7vuZiwgNuPTgQASX6OG+3ktqkB08x4/f3V1usoGBsLVp
rJJ9d4WDXaAZNL9/yyALzCSuE1Xy0nE2a0ABAxErf85RFKLhB/bVDTFmVz52xISY
PQfWxvUUqCBbVqItQSomgN0czppg4QtWj3qLtyNHA+lALRh65JBlSGWyiK9qHRB4
zhpkm4uF74qb5cKLKtHjsCwlDUcdlEqj2nG1lqgNHS0R/XxYeHMuLgKaHOvrA8wV
uKFhrHbOFT8G5kbgTK7vax6gkCqXYGNb36Af5GbVCOM+5Pf9/Vr1TMi662slMgUl
vw+Ek00tVneJaRtMcpeamuq4qf4CSH3b3K5TjC/QndZuvQBRnfxpSfYIo3664PHA
ELL8m1/6ZReAf/JQTu4av3dN+rxSm+zDgX6Wrja/pK74UKMlhb371HpAIqC6ziyc
LV2cSEFcATiTBXQcZEQBvYd0ylLmSknb3pxUPuJrEl6uGhIy52jrItRrFBx+W89g
sTb3TyOS+yC2sffSMdxTtSSxYOyVRDj1pRtrHnG3F5Kpj8Z0ICuR1xKWuaMqSPYy
BIdfNjVzrL88FyUlZTknFA18zm3gRuRfyTHaU2wM2CrLcWr/iJS7G6O/O+pU33xN
yTxA/MIpOmQmVk+/O7rB2VpG/++KESVhf4bojADHTmSThsdAe2mJnLPAzHQ0Xm3P
afQ3ocBx3+gka4WS6b22G7ehb2y2axTsppJMvaZw8CVKMMXKrdpKyQAPEdNaDwpa
XF5H4ygSPkeSyXTIDOMWd48oY72ajv1T0J9ssRJ6SC5P++tySpDlLq39nnygzIN4
L7xwdzmwMmll0PmEMIsATCgRixL5gYvD24CIm2F7NWRiUSbd8cKeZvp7iPDyw/Sw
mhS3vkqK7MLE26RvxY0A+pE5x+IVKhl94tDV7HpLTHvQAg5Yhko7rCFi0rl47irB
mpAp5xfIWWvVer7gVmeOQHi3FZyJ9/u+lm6bABXGUDVgjmn8W4cFbiT90Du8b1EI
ghOWqdIs7lL0gJLRkyoIGaP4CgihVmThg93qG7Qejichc81ePVTk9bVPY+q+OPh3
BMYaDZU7q2r3L5rphIMu1drpJTyWHYHBH4NyU3IjUE4fsM6M4/7iMb3cEmirAxPU
m21B/cHFCM0NEJdEW3Jy/wOXUB0A6SF0y3kRZHfoHw94Rz++5lOkHih2KQoolRSC
Q92Qa4sCwrxxvNNl/mQBSVFAU3TRppP2JzWJA/nBYP/rDWjwxgpTqQ8mDMHoWkl6
sw/rUowQwnkxdnzZ4YHJJU78d915y7cY0WUGIKA4bBONtG6XS2VktDD2arV/6M5c
e0a8xMUL17oLGhpoS5isc7+L8J78AOHO3ItGaEuIqdOju3mXr6vTHhby+upw4G7B
iNFvyBuFTRuk7w9eAErioYuXJ+LXOWdGo6bOhQ+Zya02CGVSehFrVHgP4ZlFqiDT
bRV601Wz7WHxXCQuLCYQMs6m7ZcxcW0t28d7xWVvMWE89OQYCCkqpeyKAW9a2lL7
x6pjDn8DiOu1nUmfwHnj1TVTBp0IxY4OLriGa4HSt1bo58F8wNf0+PzuvGOjPrjo
/eO1PHlESsw2EJ+iQKTvA9xVMwXt9GC3cC5Z7i0AHaKplYd3jyQD7JlylpMxET8d
ZkBXuOm+7O/8l7UUaWppzUA4W1Hxc4eoWQ4pwI3NM7zDFwjqVVlfjRWMQui9FiP1
V5mCTSCT+dFnSvtDv+iIcJGL9UJOIb68N4uA/8N+hZw+eDq7ntqnU3nH1iuF9Nyo
o7I8KSki2tK4RCtmuklEEFv3eW9AtaKP9PSo3E0fvrhLHt+8xnqw0VJip/YWObS/
DjI5rQhQCMRwakSEXfy7iA10TchyD5NB3FGGRRhNg1+VIOEbF3Rmg0B4CURkfssC
NO+xUd1r8hK3/fKkuyg3/TFXre8MSfmfMT1yx3ALHoz2vX5/jj/lpNxeS9qmHdmC
ahaVe6bCnA1zykkWunxR9KfQ5WoQkmH61PQFdtuPHvcR/bjCAvPCpOLai1VLuQQT
HULcD34l0dcwlHgnyQ5QU5yKXgV6vqPzkJ6Tr51Mt49TcKbeWMXlSIZ/pfQI6OmR
cSTFqurUssd82B3l6L3NlCc0/fhBqXNyoc4bGTeMosKQiRAiHvWNZHuBfjQRX7sa
NNXwMsBjVc65BvdEltWgEX72NzIOY/Voczjioy9mJ+GKkhQAEmkGHpcSbS5Qsn7v
OGM1Wro38vVtu4MoKtbMIokud0z5FJ0gLf5pjWdtwsOm/tI9A1gf/oLD1YBt9lF3
qgnJdGsSL239U7z1CUAV64PUZioZBKkUt5CcnVVuiOv4QLMkPaZdoUyQZ3A0ikA1
aQKuWYs76IhhkztiuAWgB9hPPxB3fTLNN6Kj59vtthyZWTZr9dky9ZiUFqXlNc4U
6kNf6k2MQPFVWW6ySj/6F61BM2MnmXXLM5qvVq8ag6oFbJ99tZ8LTupQ4ELw/+nY
kWoe2rOguUsXSrtOm0M3HeI/GjLrwxzEcDBdB3+MJ8mjLPwuLGw8zRzlImje2dMr
1cjYd4QGB8+XRd/wbg3PaeEjTjey/Me30oegAH2DrlNpH9w/uGnYWI3wUXguMJza
s+7GsJRrlZYHZo8FZCwFEIv5djqF303bpM28UKKMmOyedHKMZ+sugDbeouUKeCcM
S0x+W9SeuCXLWOlH5UDB3nkoekWvhFa1vK4HbcoT5XnNOb3gF/Mp4U1TOy8MCb3l
EGYF5kmu0XY18Z20V5Gov9x6DsJ/jsjsfUzF4eELJ3DJORrzTK+aJ8sNbdM9RsKb
OlbZ3o/k2XedoynQLTaFNsnGA8zkfNWaMxLB0fiqShNwjeZh4zbIcVoDumcssjLB
mhnIh6K3YFyHj+tRVQ95GZduF6gBWTKN3b8rRs4/jTrseNVJDCTpzRcsvjoWR76N
gZXgB63+kSTc4rHVyfokd/UJbO8pqUikcSbBzA9Cz8qNxQAaPjXP2klthCVEYoUY
pfV3jA5XRHLnlqxkRriM+KXqZ7mcgm5hdhCqMUO+l1Qy+bzXcUtiV758zmi3NjJU
fRBT0mzcovNGVoXSM3mcg11tTmRwlFiqqlwsSVlVcMePfJDlKb2RRb/iZ6t8JPUF
qRrzjaFXZzzHLaBHkkMZf5gimUPzUYVeaUpx4e63sZEv0KNgtdl4BAeKuC/qavK2
Mwy8WuiVVCsXlespeDrFVKLsevB0Gfsdeo0fwGW9S4oSmGgbKB7W01W1xI5wgq51
ry2m0TtwyzuAkwzinYj+ZKyNm/Xv65xICGgD1eQHVypQ4I9/p8KFUWxI8qzAHTqW
GGQqt3HTxeyWAshKnIgU4COI5sb9gqioYdB7OWSaWd9r4wfMWNNoorrqbyGqp+gF
rRld3oug6psDIZILmJChSKRefev/ig69CHYPzr+CA9ZP/Wx2S1eHx3LGxLKlUT2P
k9Ljr5OJAT2G0jrc1iDKKHMZPSzATSZrn0HrwkK3kQwwS1HeyZIYhXi4KgIgWAcV
qABIxyCRr4BxQXWncgE8Ba4VQ5n/f1U6SIBRmWyw4QLZrUXiqzPJeA7ROzNQZTEN
FJRUOmmVWdeN2DaIsgXmB3SOFbMl5kP931ErQYCK4vGuh7wXXGOdUjpyK80lDjxA
BJjK76DbXxIxusXmMGhEjZckNDD/OoZN+fvB4PiphbCXmBWaszsghAB74XQPMirY
CQjTYOTAjbDo1uCIOFrttt+d0L3g6KcnYg9oQxEmX3GIxrNOuixmenwXuxo3cuyj
SR9RyP3yawhiDTr281suEdl38O9HMBL05qyM07Y2EwWpRSrLh2hpbYlCm3f8ouEh
5PGcdZjM8HDRw7/j5LhpzC2KIGmDoaSVdasVQ3Y6eVFouXq/R13daz0M2jrVqTPP
YFljy04Ay4GLPHaWbphXZ50PASfa7gqyaQckEtc0qFvHA2xkk9tzhMUvM74P8tuK
iGxTQTjOUkELVBGSCFPndfTUfgjfh17hxkd22StNLvbC7i2fSt+48gG7FE4uf6DT
nxShmBB9St06SCURDevHPVNU8UlKRwPlsolkJVaGWLclx671wYPuf0eHSqAdS2jQ
oen+Owm7PR7RsVxTIxtZG2krIk5nrvQmTUUYnWJJ6mBd3tCPuoxZ2pVAakYfN3Jt
euCL/Gn4x419kppcqL44mwfWK9pMtqDMAuSbvkWlVD39S897JavNPt4RPwfdvtMk
BD3AOwYpDwKvL3V+K/GWHcvWugjD68m4UK42oWb6TQkkKx4cwawtyeJ1wkVSj+Gs
U6gQFJ9pX3liQr8UWUi8ZCRhxvy6VH3TnmrwNwjV9s2jQMT1GYgWuzaCpkuRshAI
NhgoSKR+eHhaWd+QufXiuEdYWbfUkdUNK8PAb1nZeoahfRCcKrgpXFdSo3FC/u3S
7Lvpog0rvI+JXbHidlGrl4K0dwBRqd/RkP2Eb/iNfg0Fw+sRYev4WrgxCr0vDZAB
YB8nFPIqjQHR1cqQUIQTOoBgdpSJXrAfB5idE3ablJur0t6SVVyAbBMFk4U+fMjX
ff7/T2XDEjf80MlOSITA/OO5K+QT5ymaydIWyLYV6TYm0MaX+KqVdNIQEVo2thf2
GGhAxI/uyYaQ0xMOJdXp/xGLb7GKkl0m00FQy5mIea3KTmD9V9hG1dcgTpfsTo0J
jPOsRWImNsEhyihi2tOMEJYrr6I9dL9ra05N5VByleTveaeoSXHVv2A98l9/NNje
Sqynd8QHFi+mk7tBao/53B9Q4ea/plbYQtFtIvIJCv4KRxXIQwYLTwUKcRxplGQx
U7MMrPThJ6yQX/mF8bFRktVHa3YkkAN3U/x5GEfZkJQWiiw1znXDYQ5vwqJEPuda
RjUlmorsT3VnvUN+2pujXr3cb7b6Q870QIgRiZaY4nefZRH0xBGcUq+yCfOeyCH4
72e5KTWTu0Zpvq89HHJx4FATbljWOoy6DEp6uA+LoL2I3aDSt8jTkM8aEP4sXMLp
Dj+3Mw+kZ29ChOpXe/EMEBUQ6xH0MZzEMjIlCK58UysVEeCkNW4M52qqji9zkvUF
nhqfRxNwQR5VwN1h39zLOR1bOe9BKMdUGnFK9i3ng0CFwVuuN5mIbDpF2SnbBJob
wVPnyV+KTseYrhoikWAg8b9qbFW5SuE4qKgKZbNGKmqOtkLDMkYtP6goxUylGTQw
TOkYRRxjtYDnmCke83QTtGpawDnPZELzBarPHgdLVuHPkBJHOud+6hypxwqP4MzD
30vewDL1zLsKxBLNh0zEjNzavWCPlxEbeZXO296GlmcpXUUe2hdzOFRyPyKyt3Ep
0IzS5K7who3IvIkc3povkM9ij48xI85hpqgsn2+hyW7QMYtcxrbmEdIGsYsSAMmP
QXws3B+QQdNaHfA69ZyECDE9KtfXbPJhdGySbnKwfRVEmTkMJCbjMdmu9FVw4tqW
8yIS9Rk5wkVetj/dnAW+99lnBrtOuKBgIiQiXLAmv+528D+REW6d7SSo+Qwsf7+F
1DVZMiHbvYs+e/Ur7HKMKkHH/l9o5psqdcKGc6oCwcWbCLwPmZmVuTc3a0KV9L2R
ke7UPDFjZLcc+trpBCmVEsFNNeMSCzV8H67DOsu9ai5u1nSS4Xa/bWnpDdycppfn
Qn1/BVyl0INIJDQu4wiQTKPKu/Jxv8mB3pza713WEwdM4ZHUgnwilHmXalJqR4N4
dbIbAlcmNRpO31EKv57WEbkzlHYmlno76BxX0hLdAvGwOru5veWjJS3fzGmL6gys
WyU6fp/tHkU1bqoZ3nDhzIDE8y+2rulbkJlK0zsmRS9csu8zSn25ZpbMEe4uMsof
htcCP470IZnfs1ru/vT6shDjZRH/95kCXXGRd4ERfw0rAsWwYB6ABbV/Ne3BpfMb
5zjF0LR6QB97dn6exQ78vY/dUXn7+YN/BZn7muJwvbTfjPF4CdW7LLRnOpsXJ8aj
zNszxkLAGIBKRYzXAUJAQxjwm+3H38HudIJPr8AmEzal8Aa3NqEkm+L5swrj8nwf
EPXch1JQ2jUgcZXzu4BSXTBZaRLOvvuw+baZ7Slugw+vzoEOKC8HJa1ThZhL22B3
yljGsCMTvCRz8BGtECAaEM7qir0hSfIGR6hAPgYkU4y/mNG9S6/Zfxfviuf+bKKa
SlDu0twBP0EMp2G9qx2LGFtVGEdfQ1JPylnFr7IGoyuR7dhTwzW41ZFWY89/RSs7
N+DVIM1kxBi/DmQ8e3aEZndW+2hvdGGsw1SynPu7EjimyJZNP3TysoadDsQG37ES
lLiwqKCxckMSQF9T49LsdvjYp+gAP+82H1ya65eH6HdxBpcTXrHP81CFDZZTQHIx
s7b/mGSDxOM+ny+Y2Tr7PSBH8FlrYVLyddQ9nw+zmHqafUJtL0MqjKE2t1CweVcn
8fzh3WAOnEL2APO1N+euRAJGpErhQgWOPqWY5y/246tHarzYPZ3G3zFSmbrqxbHl
M8nIL40XqqgBRcRlr+J0baIjrnIp6YLJKE5z3LkuwD+uYNEehZPIgy7TM9SJ8TFs
8elw2U6jP1xnfs8Q6N+Jy5nRaew3NY2KTGhJqMn81YUTlAr/bfMvtZRLVKvA2aY4
xe4Q/SAoEXxX+9rEOsSVr9giiQNp2vkjdK86vpnq7DGkna02rk6jdEYdHg4Otiv4
tO39x8TGASw1KwE5KOyNvsigm91rGMhk1HVPnEK93g343uE3Su6oBQqZpHANFb+Q
TFRKxgIJAP7EiGz63RVEmYd5lwsnVEC6Q4u230Qr+GiQ6wdpNVxjv4VZV0b2KIQC
r2yoaxgNIVqG9V9CV3XkVstVpHxBHPJLm38IVyHsHooAH0m0TZENk969YUW97krW
jTtfVKrkR0oz9F2bqORFcinJxn/UWnKEwnNnmIJoJ4XrbIv1ILlSOR2Xnkkst/4u
eRxaGeMvthKdqegww1gn6D6WvS3GKzUxvnCe/7IJob6uE9MXJry0QOLLVkLnmXKL
WrQssSG8Bj4gXMrftBlKDgL0r9BJ4Yzt/h4yIgpMhfAf97o1QHd1BzZwG+kEGgI5
w4Pzk/otI4yulEVhcCfadK9Ohvrm/VB93OObal4g7w7Lu1hgeIosq5HaMrEDmUOV
468FG/tgdtVWo8o0aopoodrRaVAnvLU21psOflBhB8IoY3VMP0we7sQ+BfWHF749
IOnZrclSBwUEf9ss80/dWRLyjSsV0+gq0tYuXPYW3l9GJgTMHy3PTL4xj5K1VepF
SF5ul9r1R3cWnujPbNM+UuWpYoQqqZ8lWwNbOPwVvHpMfNoYpeQLjtpYlfvc/0/V
BpD3P/jOmtD2ERgZjpdQ8reVmmFXjB06WlPBtIi6pzZTyHff1NX1lfFwxVmw2tl8
uOgUmURw36SA2O9WPG6mMtK2lpdJB4G9qPURGfKOracu270yqZ6/UDJc94Kb0ETi
ClA2AZpweKqoIZv2YaX0c6OzeqPILGENsZCEa0bMQB338LzqETr/z1oqNzQN1khC
VpvXNkz81f0bNXUYu/EG0zARgIn7KzoUvGjBR91z2utiPF/5ING/Bj7u35KuN1p3
jwoH+TmbpvspT0rqglp3t8yKH8bgjmDLniAJWymBHhJL0spdawHLmnvrb3YPDfCY
1OV6a80NEdQNXLIkzmi6TghpYfx3/VfxcqZ0KeOBKrK3vGNW+2EL504jytTVdAQ3
MdQW4J8Bw5ur8XvfqQb+W2FqFkPItrsND2Tbyv4hCAewLPbviStNf7d7PvaHJWQt
JGk9mo/0bgUGz9NFsCKNe+qWpq0etIsBuZkcFQDvsVtworQfkKZUIHXMav55fUeO
u2YzU/L+3/zDdqwXPYlsYGSUzAGBnTl6nTDeOKTB5w6uE1jEGpJnJXtuDjq6iCYY
VHEX+xiUXmR0g5iba1ZLGPuNPtai49wFOtZSnxM//eusVs72j17t1xfn/eGyz7ZQ
jRDf0vU19S2jnWCeThiiv8GLoeuB9L3R6MHQgcHipngaZ919e8mDu7fdsHQSqJ94
lCNrP2NAN++Oa9k1bJMB8frfSFDsS0MFsgugsijgU4cnDu3yNHuOqydM8rtA5zch
o8UFpulJJC8VI1n2R/dYXjnriBqFTEAH6HVNzgqtbM5heeJeioyPFcJZcXSjhHD9
anNi5WZRqZGhg3nVKFJeXnV6FlKdl86cwKv9ArRbSsgrlsdGwehDkz8kdjpLpngO
qLflXZS1AXu9wyJ9yYoj0dR1zqMLpWsQt3gW9freyAX1QwTuBhi0pTGAb0lXViNh
NpVSePhXbgp56tNMFJxJNIiosEmxARYXzQrFV695IvFCvF/vBhM3A4GAqoiqWFL8
oNB2T9MeBktApP3S19BCoSNL+cdIDZgIKQF9soxbdwit7WVo4J4kDUpmoodUHGGB
fuK+T9/VIosqoD+Wm9rgmtTmHh1U4Q4z9rjxKyVdT7mxZY8NeDimEjYeqAsCDg6h
Rl+6bcYxfeljHESqQa3bvPKBuJKUF2zdrf73QugRWnSi5UMfZz9fJcez2h+emICe
L6Tchpf1ykhI0XdaRfeKiO6cJgo7Ov6uxkW7NQtX4se51ux/u2EqlHb9iNdSiqem
SeWejNiri4Q+sCuTAhQSmXsxpuy6R+e2J0zw7mDhpmY3GrdPX0XmQoodASqN+sNv
es5YdlVNa24FxApafli+9kEMYP/xsf+mMcCkoS2JBp3VxWv26mM9MDZhCucD+HT7
126jf9YM5jRnbmwRndYPGooEyagJDlU2WoiKH2cad44yRLNmY9q6IqJTP+Xjs3Bp
Cg77iUSx7nP0x1KFHovJnfh3qiNzF9kP8aiPkrRsMBkAxDVvGulKzo8BSA9WO9eY
WdNpQIDQiJNhDnhpjY96n8/Buh5OY/DkPD+DUuHvsZ4QNb8jBMu2OjDWIA2gwfRg
t/mbIv0Zc7kjp7hj4UYSt/BKt3Lzxfiok/MNC6/pKEmOain+EilSKOU69ZlQoQM5
RQI6jYc81jevrZ05pttXsKisD2N98PKxFqF75zovbIVvZW2dKylNYpfSvrPGP1H8
X2KuxbYOeB9x2wnxeAOv4oX1uV7nN3ANfiNAbbW2qhj4kdrXULTm48NBKTSzLfpp
Wc6oo+R9llsux7K2Z7XXFRp7E/HGDHuBaKdVxw15XtmJx7ASNrq0hWDLbOURQ9x8
ynzsK6VQig47bxEKbE/7ye0tBHn+PFBaMPNUVZpXTkKv/66mBbdG7syLEy9POg3C
EbyxncY0H0x6E7Zyyff16RijmE8cTxSthFncBXjFSX2MrJbzececVYs0oNl9caZO
OW3suKZz5RKWinllBp7qSaC7l/hwCYzU491VqpLcXdEq0pnrZHQmi3pCrJhoiCaX
4J08kzh/W30D6Twl+01v5Zh58wAwZY5sPBNHC3I6NbUVzZSxu8CYlBJW0lD4xjwc
OMTws3NTyPw8vSj38MryjzryEaQWEWn64fpk2TeLwx+zZCEskP9l9zRcaTNaj83V
pTQ7/oNcKwsBdMRF2jQw8FJvL6HqY17RAMTXVZuKNZq0YDSiULBoz4hG3zarWhze
sMtVj10MyG6DlvZxbHEdDnmFgGT2W09s8IMPChVdHYQ7TV//pB8dQS/VIO7TXelw
re3DvlCQaVYtLX8zuWVY7Ujf9kJxn/gOYQBM54cpwfgafsH6i7xTvMakDZPbulwn
PrFPFwL1eT/COetfUQPpIWIp73x47n5VTUiGgYMNMI0OlnrDeiIccEeyNtLaXoXm
DcJw271FSR/VFpIn+jlpZMog0kfHHxwlkMicVBNcdSFeGNEa8ncSXq1vzX50EKTE
ruYK1JEdPLVw6B/N0X4ZkLz8vzZCuUcweqART70ofCVUMB/flyVBJKmKVLDP7qzm
/jsopkHX/anLyVJcHgNEeJ0FUTipWHM6iTF/giODSXYbdpA9ET5mYvfL9TyyB7uq
08gp4QK41kr96dVByE9T6vd1zhUWVIgkeCkhOJod/n/SNN+FumWttCmNh40j+i5j
4H6fd59tABkC1d635s5xoJ80qDLTK/0fRDEWoq0wrgs40znFLEmlPJlWW+cXooah
cnOsnUbSWe2bfIy1MKQbGQLP/btdOlnxFjnOVmPzGG0roSwvWsR4niC8eFtrpdME
K7OwU1RzuLVNjyxcjPcfr1qEZIV+5ijE56Dq5thhfKtY+YeOiLIRwq1XKb+iMX7M
hmOtNOze2XL9KZRM5wCvgGReV06FUsXz7lgnt173kJNS8YlMhc9CC8tRPCgUfWVE
6dcTZ4l7flX3c/Hs6JV2sH6NmhesD7+VqEMcA72JHU2sQaLn77t1jryqLxf/aPRm
yHLqlr8rIbTCSwg0FIwTI82ikJ4rBRs5ZwqQq0tIg/+XEbGPB4xkfzovmNsc7xxZ
akdcdijdkmXfjZE47rUMIQfpHwwYLpIpzfc+4H//8zXd9ADK/8GYKRnzAax/VWXd
+YZdLhJFyeFCKXzJlDkF8xSSR8XenE6duZxVDKWhTDjSFNwYTqBm5NHU0dZzsDLI
B8ZqBKEyII8lm8jQ6cGkCJZoy9RDuqNwXtF2/vaL9JyZTz+x1H7BsLnJMDF9fv7m
xHXyyHMuxWdy1Mqi7ryEzM61Y0JySdQTZyWnzRiO+GKqfXiIGMWy5QPcI8cfEgvd
JrdR2/9Sv8JU4jmBFkgj8qZlSzb1t6QWSs89tsq4YQgHq/IVTwPj6K5vKenjOsuR
dynwAjpTiwpTTaQZWHosVNAflAj3pSkqKOJdZIlKs29BIwOZRODqvqlwgtHptO4x
E2LIYvWdfm1rzF677r4tOun2MwXfhnHbJXutrQqeY2SrKTtOKxYTnbigtgI0qWLH
wXtMAp3DElKbAnYl1SHYpdyH1p4uU6Fp6Th3FD/MFXxAnXpxOBLlTOEIRslkzybg
3rZ1kEhDs8xCkaK9/A9FxlnVVuw2WGYehMGo/pZac07n59zMZ9Djk1swuvy15AMM
D14dCgpkGHYSOFtgWn31iG1fRlkeKoKxef0p5y5JX/F7d2awfxoHtExOJjq0mguO
n1RZzkuP7MbGhIC38AvTbRLM6cJDm28eazLvlM6o99ab47GBQ1naPGvCdjwxTQQN
ydbacAiySbL3+EqU35YqimaB+sgbPzgfNLW4XKLB50FINjei6kDnVZVn31FJ9HrN
uqnfyy2Ur7+LhmCLhDgqeKph2RyfhhLx3ecm8f2Z6JqLmoIL08RYw3sJlNocaXbm
TefVmknWQp2emEvKpUi+xbKmLw0Iu88oOIcUJCAFRSBjiG3AGXAAK+7jgmze6t46
TH9FPw/H2eIVQhOXdapaph/OpP/TakZgHk51ETOHioAdGYYFeHB+MDvetY+8qf7u
MucSqFfr7z2QkDgZkTZmgQ9DyYd6USbJVbgEjRS/HDMwvpxleKtdJUTeUTS4f+p4
lHPQkSrVIzLzdX4eYlPwa/gI4xyvNyQ5D9zHPiNcL5GEKAL3tHFDzYKW27HuCWA6
ehQ9/4HTHoKHBlTHEE9dSEACRdcBQE0ltvXwvCWpVAaDLktWTdpkUriv9wjQ2VP3
3srZbVQr8REB+b4+GyDcOdaTAQbnoZztcD9YX3v6X5E1S3hBXUEEfcuSBqpwAcMg
MqCQ19L22622XClPkIN0k4rHQAz64Cv/kNbRtDvPaiPYOtr/LyhmsaHP4NIwW6af
k9IUzSX1UjNnhOpB3cbux8Vuekb18fmggQJSZ2LfMoaiN/DbcB9cpq8gHH2ML/FL
T4vi09HHR/P9KvLxRVsmIobpvLhsncKRgycNd/xzsLGcF7RJXNX/RKvU4B8G+owy
0WdITDdIs88UCs3/3cBtlGUTwUEszpFpAgSTK6WBSpC91Q4P/sNNDkzzrTf4x703
2+b3NZ0L27UqxsruyEuIm0Z8xNN7NVH/hjad2v7vx21+4/yY8YP2VxTR9XqGryQP
NRUBIhp43kc85SVZnD7Aq2+iGboviEKG9mRLTjAPTgMl7OSoSXjr2Vt48GPdqcuX
MmRrkXllcqDKZe93Rb8w5pv2Jjj2YcYyt2c/iimwBbi0I5Br3Q5LnA2OVETmWlAs
NxO5x10LSWWm9KhjstkcxxBO6mutXnYWo+bW2liAAbo8lSHUQZNpaMvZwbA9egCx
yNFdYfOya0h0SoqUlV3hqlWy3vT/LTHVCeGYUfNqcsk6r4F3+Neh0E1tMPDn8WE7
smMh+3r8zDf9zicfOHC8Y+L6L1OijkZ6r8Ob6/kGlogggERNye14cfstpF/gEWvM
Qtk6OBxltAgL28PXZOdPE7y9BxtsaVCuWBhQQvl842C8UwYw0xrzPxFZ6L6p+2j/
1nNyDq1d8CVhV4ZJ5cWFp8W2VDmCaX0v2yvaIaM7Ws5HaKK1i1e1YnDY/R1jekxM
jPrmZAeplaXfEMK10BRo8Na275xnX396v9qwZcFveWIVvlsPnk1Tu/0vHU3T6QiJ
jtRqOeCGXhK64KGR8HHHE1WMw9opZImFy9bJ5pwNxg50orEzl7a4oXrGR7tVQ2kn
csOS2hpp7skIXXwpB7FQtOzlhFnYx5yePfhxfnjwY/Bc+jbWTVidr13u0T/UQsWQ
yDKxmOzzzK25Ce4fztqTIs/75XpLeGaGOIW0Z1jZBeaPsoR8csqCfdbMAr2xh035
P2MrvDk6plQJxyfGpmQfRfUELsK8SQqskaza1fuBr0/ntV19Y1+P8kPfWUaIPvk/
/0FMPABApOnJDwi2eYDfRt/h97DL79vO3Vm3nf1JnSy83dQ/T2TCKqUg33hQro7i
5ZGN7EBfSDWXMqrohNgII5gXt7TLfWa8N6LlY3eCogNtbNImh+KqR18B4EZATV+Y
mZtr5//ULe/Ia3pJSMWYcskuRdVWXaMRBAH2kdxE84oitRfp/MnIuhydFzOCCJta
KTHvJtm19rdhEh16CQLCj6Ki8scmK3mCdEp+thSeF0++6zaKeF2KWXuIFKv+cAGv
2Ng3z2Dvd/YTVYAZ++4+9Js2BfmJZ+Yb9t0WI5eg3EbUlrG2Y6ah/ovdfui6yywj
fK6KlgqCKpIkYszvg9fBcmpKnmT2ObcXC/HFM3+S4527YkrzwgzmkGIdvigB9auk
sVDIPP/+FBaRb6QZZXjB5vpHR99FFbxT08QQckubAh0c+H5gVeqqzy6vDth3sdRm
RvUnn5swhI5YmYAAVZa0oMIhsJUAr8O58RZt11zIWFS4G5/u08fJNtNkJ34M/B60
nBPCqB8QG1Sg/FEuMQUK4tPCooZLqbOgcdCOEE6i37t2c7rB+Wj+kxWT8jhs6Y5n
GQivRN7kspxFRtgS3kWdlzUyLmDoDQRX6oCdl9+ovExGWsDOZVYmid24dOs+bEX0
EclcfCrI3W33bIpbhvrarnO7vJ9xlEq1fiQbjFT+biJPaXTS/kJ1tBvrfbgGRpIf
Y3MzUYv+3Wv+h2j4uyFFAxfJ4+7o4dpRRnWk7KGb8qkej7hHXWMbKBRmIKdKbnpx
J5nP/amiZlI2ZWl4c4Z8Z4Msp6pN0dKqgjgtbJeOCDYGA4rbrHcDjUgIPd6HQBXq
UVwkSjcbutzbo5AzgFkbqFMBIjDriXT03+wsPBB0/fUtQbsPkLmHJhK7jD0D81Em
pzdqw4Sk2T1zvnLSweu+pH4sCPSua0PJxr7PK/IGyl+RYYftJgU7sLG0rkJnqGA2
Hn5LjExDyIVPVD2Pd53G0LhOmMqzuRh164Y5KWYbuLHE6H/lzRO5WOU7fRF231N6
mRvWeNQa0RR2sCvXYyFCqbgGjawM6K9UG9+lgdfapJa3XcYz7e84Q+xYEL1a8IXx
qJYoocvF3E1NmChgDeDNoZpnEdmLytCS9ihos/PZRQExdtOWTXMHJSx8rrNBBcKi
MgUDW2QNfFuNX5anoiJ9zFnbmtrLF3KZQiWoMqJhk8mpR3uh3smnru2G1Bqu7+Cw
hQOP6gG8xUXMPkcXBatBmGUh4u0h2Fqd6OuJAq13VplMKo/mP8Qp41YGv8AS+TiV
Rc+jRENdB7txGWt0fLjioXQn9SGTOve+j/oC7a/YLkRJQ4qBEeu/wfwu4qshrnNi
4plse+vQMv+WxqnUX5/mxaDKcg/S/4pgDoQVZ+RnrnVoUkUBH0ImWRhVtHTKYvEZ
VPjXjg+MW23Z2K7kCkrvxnl19PfuwKTE2n2HKnbTgEjFZoMknvUFelxRgdvIRVR6
bkGCyz/ehYW3nvYpXMCv48sAUPI3A5MbCKj9LM0A26cBs/OYDVuu0/JZO0kzXMOG
gOEEPpWu5N0FySnIAGH1cwxID9lWGM2gI5wAhfGurQvv3KM2xu1uQS4JrYbagvmB
fKsnQnHdteMNOmkSDos+Fsj16eCkJuVv1Skwu9fPN4kE76zJ/KdIQf7ls0gZzm3T
kipGFEinDA2DBnIzuw1H6w3EUHw8DGhT6Vr6oZ858g1tIjHbIKh3FQ1LlvzVkyHk
H7+RpsGdnmFR1jmRZM4qBSHdUMhxzkrwa48EWAj2dSEjhDgq5gpHu26TjazBlFwO
cZAzkh3cndbyn81A6ABboBABVZdCngiMp+7NKCVIrnyhs9nPZl8ow4dNpv5hW8cW
wScpIL3jHJvyi9lYX7KWoviyHKxy1YXl/wjEaGSw3cWKQE90Y7a8VFQMKHG9l3jd
aT1weCVkQxcpfFfnZKmAMvPjOsD+G3pfhBsv+8k1QoW7QxBhPxoDHuKyDM72YdJ+
vStLq7USW/QrIESHt5MJlmZJFTx45/LhAMCggGfdtUulDvkTDwFl2KEs4rZ0xbw3
25ASIeKIqAhmviVBqYvrmcdeFHvz673Zk435RPINM2xg+7tFeg93iC5pYjYn+fn/
LDIfr3NYmziwOd1U8hhDl62yrum8oBOHYZ+hKt76lHUfvmkaYezeHXrfRW5mWP4l
kG0YNJFQOgVxnAhOWrpMu50ajhF9QmnVi2GvcOloBg3Ab/yHuw7aXQl4jwO7EMt2
EwJ4BsrcGcgn8p/jEurhtBTs1splMSwHAvK83mcPhjM+TfvSdEpUsm8J6Zza9jMO
fbHIfHMX5zT4D33TUyaPEdAouuXkT/zZRN+VrlRsyY9JcQBsKd5If2ks+7zabXli
97FqLwYUMdDt3cTx/rERMpG/UyrLG9f5IUAGUCXgIe/AID6VYfKIE0ywKIfBSFyD
TeT9hvnjLVAgYDZrIa8hOKe7vGSQ/vugtuwNXM99+xiNiZmtj7BZklVfjfzV+yck
WhTl2ZeDUSiTm3P7Hmzn0iN6gIQZoKQdrS68oKGlMrh+krctWNzsssJGqAGxEFFE
Qr6lUHZE44HXxybVf9l9/QfPpdR0p0Aoeb7h0P3Tcu0xcvZ3yQ6dNI2xMyquMFMi
VvYghe/kW0+2fZd5UH5zEXy6gvUVWhrgw9WlxEvS9UU/3OxIIgT9kQ4mJY6pQR5m
33IBC7w1oXWbYhJSypO74moA+ETr6WTZ+keJe6GZMhWG0xv0wpq6VmzGkxzSkcpP
gi1qJa2MBeHX2soZ22u8AIh8l6oC/2MyyS4JwfBe9VQ5BFtQk1Ikv/5pa8iL02F1
TXyyqJgsXZk2C8U5bdT+5IRdjDAG3qLrtH79oiHBCgBKZ1J3xI3onxBohO93XzVo
+s0TLy5jP11BpIIjY/jsENJvcx6vXpTHxtQQFAC9B2qSzxPVGEgdL7m/FdF5piwE
cwbyrw+SKzy8J87gZ+Cf4r4pXK+sUQE+Nmu0axX/0o0lqYQ1lvJ/xmFA9s9lf54/
kL1eifnOA7u8MnmdmVFPNq3P/u9W+2E52AzHut2xkF5r03p358px7TX3Vhaln5Ox
RCrMOZVI98RbBUVbU9znMjzv8vpOtg7gIMXUUXYHMY2y/4ZopKTXczFzVsZUgkG2
nwtb4Jv8UHWz+1hpHvAbAYqtygkQuRt7GCqXZrk/OOykjDY1YCf/6itpiR83gflY
cUdwqQJLCi1faS1J+7ZsQ9OnX2598h35obpyqFyK3bmRzJyqKqMDe/g7i6LDK7yP
mGc5MFasAjZWhudWlboYRGnqdqXYf6x3Q6fJN0eWceCsff/3zvC4Wl/a5Cgzu9Gv
8uTiFBzthUT3WMPe+kO4OzQ6OFBSgGl3HXbgh+kt9uZcgadGTvkNennWUxVQGbBv
DMvw65GWqYZBG4KJqD5k38E/9CCpHLkogVS3rrLOC9uQ3lSa7J4qK30mvfuECZ0m
xSjlETXILw5rqmZek4SeiXSpCxogYr2m2BALO6ssV12C04oDHGC5+nAhPvZkG87U
4VxZ/7dVpR6lk331mWlGb92lZpgzm+4TCv0liy8enRjfdQqINSlmjJnFZ5drGAOm
YLtM+xY1PrnaXPDAsdGtZp9nqJoJEptZaMEAOtB7tRkOyLcvhIGzk1tprnkGECsc
qLjMbpEO26UtQiYenhpiBsjTkVtU72AqfR40cF00CFEDjHoJrcyFN/7tY8uRLFKV
tSJJrPmZ+TzNhI9xef5y1x3YlT3Kb5FH7tCg6kv0ZfeRdri7D+XC4uEeG342oyNb
wku40BdSU9zusEBWDJBiNzyYUYTFHfbpUKoEgjSSn0BYFcpBUXfvxbC9eQKGPaDQ
rLxReGzxXW30uXHGTnfsJyA66cfTr44Bsr09DKlXHeNaW7jyuc6mfHPSWPMAC17Q
B9gEFUBBqD1Uzopr2eAcGENe3XbTlUwpe94IJhFhstEtqGwYqgghhchk/GkaIVkQ
vMm71IJLRxtcOBAIKqIi6fduSdtKIIxLz59BvkoCbKiTSZpr+y3k9rEzD/EkiRFl
z1rHJ6eVU/oMHeBqP4e+Dea8w/QTH7wbHs7y1SIXCuZC05s4DZhaR1JX2/Mqecry
X86H+Xj/XiBb80p7G0S7KdJiovkIdvz4mL+QEsFtPf6915t4DJCxLohX3dvgk1jb
alLBEOo57eXljXK3NBRJE+QPOrRuD2VOpbrZYWuBGi5qMhX74e8A9xK2zQnn/7oy
IyHIx6Q/t6Ii91vGPWO2TETHkiPVcb93kYXokYoBwoSVxB2fw+PwUjyE/DlRNGA+
1i1h0dCO/TKre/qFozMkDDU7BhdKhsIF0eDMYaf23CQ72/sisSBvJI0YOOMWiyWI
JFPyAedO/OmSslv4xEQtQlxxx0CrKnrVVbuKXosCYyrOBQ5DpabMOVUtx1NjI4Ob
+l8TXz90r6zzygH6MX3LrWeF6o2VZ808nZMpESrQSD873FZW5S3OjiwEqPauklki
SvV/d8XWGruYW2WcXiz0PbDgx/fejN/lP6BTMUV75PNHF2xcqaSn0LCr36rVsuHW
u7Yrqesjuopvk9bkAyRNKn8EqiYKseEBAndSeUP2FGCxLdM+Gldvkayj9g6sZl5N
jda62/iPPBlLdIfORwqQuwk6SEo/KjbCX2/3KuHUp09S0zopNrIdPNH7dkOeb0GF
AwcdYjISe1qbwky2Kevlw56Iq/7/M9r4TYfBocTiTwnH1yJnXGdJroq2Nydf7pB8
MBvesfsaDi66n/lR7k/+Y3CBswxEMP5mlcT1J9TE8HfxlndKqF0cURkr6/AtIJwQ
OKu0WXL/QzzX8TzP/By+A87HiPsi7Ag08eyc4UDu/WCsPkyBlK8BLUxXKvzamyDb
UYMP6oudA16HzVH2V7/kQ8pcIPdFq9Uz/rFvhJ4KhBvRAaKTvM9W9Ol17BJ2P7R0
0t+rD0pyir0c+2YHNKKxkjsCsmooF8FdoN0YGEnioY50WjEHGZ+SYTcBbIffS02s
faPeQGSr3v8XsUF9h/G+pHsf0fvpRpSrrPrRdrMfYdR1oubdEMEu+lsXQ/DesafZ
xlvdQiThVE6vq+Owh+7pMx9WIhrkXOzXuu4kMefjMBs7c6BfeBbo5tuI4601cARA
3aIca758DBG4tTENuoDD2QUbdgCI1Qq0Po2G7KxKN5q5oY3rT3hLqBBnIadHNVCA
mYvA82Xfnt8jJpRZNdYEdvL7r3YE4o3/fsha2psstzAfsBZiNzN3m4Gnp+eJKAVr
7iuiow/xhiJKDCoLilEHv36ZuU16P8DM2DaMvOJoinyUKQ/dkJXSwQq9s9f5Fi6J
MMiPHPfcTaANJpYmUWiTSUQ0AkPTAaIFzONW4y8HvgSngmP2VMCjEFhrJ2h3oCLe
V6tYuqt9lxVsagF4fdEPKK6Zo7OD1YrV4U3aXctgpDuv+gO2aimiJQ0ziVx6G2+K
6eVtNXyOvzoMszVc7gLCBcQssKv7FltM8TVDimoqanIa8hld7gBH9s5sQNCii32B
+njZAaYAZ0APqu1J2ZdFRRuNBuMvavzHcdWK8848gulqGm48HSKon24Xn87dLPSz
ub1qiBU0rrnq6+nQjlUDAxjjZpRm9qVYoCmGzLNwJIkkflkl9Q1MiOcSslgvift2
bzzzxtMCstBNcEEyURo4n7PdpjW/VZSOlPB/3V/LbVR9CmxhMmCO0DkBrLJlg28a
OOl5ujqPHHkPbMzHTuT7i+nVcdT0pGvhJco2VR6iAzmrZ0mEEM8cBRHtOs/i22qx
QSCRGDhr9zFfDm5l/wVCChdDpVpUHsT81WUO/Mw0aqQBZuQn1oQ4FXRgQTXSmXxV
Fm5v/Gi2sTtmpOTk+m1C6GErc26TANsl6PpTaJun3z6TEz4snnhiNdKzj7slydOy
tw/8NkKrSLPV/T+79jVIrinzTYSzcYaRMNA7FTpFr/EmR91r+rC/pHo+AAQsvtz4
ASYpPnkTvC2z+2ed277EhcJhZHb4T485nWQbf996T6Dvhw/4w54RDUO1p3+ipUCn
pNTqEm6HipBwkC2er1FTBhKA1xDo/Fr7d9rX0r/OiWt3fA7OJSPTtaPgk3oBaHIg
sOBIbe0wq9kG5NqAlwp0BAIyKI14+Z6KUutKBKbBntTpVU1Dcw+s6f+8OqCm8vo/
FBffJMltqGFN9o7Wnr2T35s9zFXBmYMpd3E2ozj0acplzoO5+4rrNBnvey6uOQmA
uN+/9+ZLtiMPqivC2LwUcfo20FfV+uiWrDp5h4tlu4LS3FLp3LYgMeWJ1KLeqTxY
fRjfpOPX+xdhBj+qGHK/c9Ve/OvpO2c907yd+5TEcOTNKHQvZErQJTa2d/LLhYBZ
gcDJ9RwdGSGrAPfexkMnkt9AOlLnLP97enb9ruzqi7kPztmd10AdNlVbXEQoJxHS
lpYOZg5yV4l1G9JHKFJasguUmFU+9+ppeSwQzMtdZc3J710IDyDM2AxA42+W/8uL
RZ2RcbsTQGq2NDV5x2LIHco3PcT2m03ZKeBLs++5eZLBIKBPOC368kSIeBGNAyB1
kJSCTJ439AUsc+hH+fFHoTehMeVc0EF7OAMmUG1B2f1rVG32aii/GOPhcaslY7HX
zUMHrRDI3ErdfwYr78jRNPEKf2BAtZylTqZcg74rJGNdkyph2HVHLrf3DizPauCW
YN+pXRY4JgSI/01Mu4FR3HvVX96+qoIRxBe+pRTmYnGTk80DfpBnvr3mLUkLDS2E
BMVeDEcCbhDyUzVq3ynohRv+ff0x6HPWCBmWct/5Hd7XTlXIP4K0GtxU50jBsrBF
kXA1gvBmKBrQsR8WTEqNFgQlmUnl/sevytctKsUQcKW+o1R5r4cJc6+vh7pmNTBa
vCi4hDGbtsfUJNL+h+CcKfvNGwvnpiE3MubogCi4AuZk5jRRKW7fvSNja02/r5bw
FlfS8autCnJFNILaFMoajRU3fsQ9vUGwS80qYQixokJGef8IKLL9DPb1A7jR7bq6
SOegsG5JpQiiUgAaGLTqTutrFnhnIa7EjDz/Qr8F3tLqj4l2e81rUyJcoGRsUr8I
rOXz28nKuPhtO82omk82b1mrb6a3zm5Z7Xbh7NqpxilScQvzT4AUJGpcxEezwPNG
SneHHsEcZV9fiHJN7n0DAMaY774idoBlJ0CcPI04R6//JQihi1FvnWUKDIt9UNai
lkRQVzmNgubUhFQE54KBBU2ehdm3yuxwz8JW5EcGMYa0+DxzryXUpMq9kZ56XQeh
8u2YocPRuZ071t3HXirDOyt1P6WnhsqEzfQ9SZ9snZ3SjtiIxrExivchY8illN6t
DZK87Se1KciDF4KPvY07+G/jhMoF4a/8br2War9NM1TudSB0zUlv3kWcVYXCgXh4
GYPELPOOmMElD4sf4ajhQ2SblMbYnX+1iLOFr+JjYqj/mDDuVXvN/z/TGr/MqZjQ
/K7hYwFfhBiWyWCUYjk7FWHCkwD6KaxfimP7dC1Aq7a02qa5+KeC8IUE/G74nMT4
xu6J2Yzqe7VUrv6wv3LgAu6LGzvioh6ajzUn8JEJCBbv8ncjXtWXoyI9cCJ8qaQO
LiYq8K+Uk3CK8klLsfDvNxIIPKOYvKRKJcm/6smalb9alHGDtf2O1lMxPVdyFbx+
tfLyceTAQZ8UiPpXo54v3Hncfvpi/6r35gjgmlLQ17492h0elVHUc6/VbqpZvIM7
4Yi86R6GCIpfjSQ38s9xmo0Dyx0APlVDHX4E/C3ZDj/VN0lsZmmOXRWCvM0H/RqF
nN0znusd01esQ1dnz6NioPgZmgfFVxIG/I8WBKx62y/WTMSzThzQavlvmMsvtNUV
LnGEVaOyaHe8Yg6QIH/cmqkqmtEitrcM9IWzaiDe5vuQT9l2RipaQiXYkf1ZNmn6
UGRMSJYKgrSWMpJ6WPgkrYbYwb1bope14xrLpYSaB0fcLcs/apVqF3wue2qxxQ7+
ZeJ+a5bIjc+FHXaPnriBca/nNreytW8mZJ1bepZZFNc8ObhPq0V/iOB1W5REZRVa
iZxB1qkvq9Z4Y66MWTYjKdPQ3vNXijieGgC5Ts00jDsshdAzK3Zl2QdjsmCk3rtU
S8VB8QkCWmyY5ZZl2uJ3v+rCiqoMp/Q56GodJtGtbc/Ji03UezAOBrJHcElBBrOJ
GmqiZ2fqukz6IpWUg/kCp9KGwtToOBkA5cbCmQ8x3fp9y1V3vQvBUxtAVR7obJKv
nI0q5ccGZb2oi17P8xMUEPqk/3aAgck+yIzyAyPjh1Nou+z6Q83ha8vEb31ZjObc
NE1Ge5lBWFdBnEQ1NTVUHQNqATAnJ5d87/J9npRl3sVybltHrhlhy7M6HlJ0z0z1
pPnAiNq4QOo+hQJHUKOlMRtRqImVVqN7R3JznmtJ+ubkHqo50R0fhBrEqDa7S8z8
k4qB7VY2chPniFJyCs4zd97wjw/j0o45Yx/6KemrH+YFD9NNobHK/EZ5KWfyDPNO
MwejogiUfZICwxHqOgbbA+p05BtY34y8MXgRO5XUgBLeL/PSj++U2h5HLCUoWe0Y
Wt7bXHGKYmSoVnYkAqinZbyYJq9YouUClRjE1JLwPtwZGXQ5AOPHtCwoZb86ZOm1
QMdou0m+2oPuhZGyJIvDMMVWc1jhk/n3Nu9Pqswrkd+ZSp17Yz8vOa5hAtKgCmXm
3zFSUYEqwgmwUxmXUbscIyLP+gm0y7VFwFYVdx1Tyn0Trrcrtt4toDA261YaDkLP
Lem64a14C/jOEhZFOHpLJtHjfynlUjmP/UpMyy+HOVXhU+o1NljqofPIM9k6+XBQ
QMhXdM4FFVdDaYTSumfPwhaIcrIYvaB0J4X3/BjfSRmQCN98LL2eLLJkPhPqUOri
rVBf8kzbzJKWwUVKXIK/J8A+d8mTkcT3p4NE0SpyeZvlBTWKt5zUwD8yqIRZl0YW
NX7JXNH+/BXyfqECuKwlBTbU2GToPjPrlMY+xjqyiL7ulVCLFgfp+Jeb5bxsxEVx
so4T9KQWbmOL7rNdEUWWcVZ2k9Ck0G76tTpTUi5KgdRNIc+0r41i87qLQANQ4aVp
XEibQ7l4Fu/WxfmUCxKW3EYKgIdclhRMFAAnS+ntY7tYXl9Xn0vEEnIacGKV0lWk
v4rCF058oqaZ+CPIP3p7Lrb8PrUNY7yEXqs6tjKlg6TAFKzU12bvfLgBYyZIucNe
EoFUzfKBwANjKWGxDbNc/PyCvhXm4OLIoY7WhLBr6yg6PrOXavYGDjcEkV/hxkl5
45QzC3LnfgeJl89RTbcL0tgllKl4kMclKj07mk0d4JoZ9JonNPC9XHXu2Jf8Pe9r
7iI6o0i/jrMXKz5wHH1s9aGeilVn4DHRyo8ff5eEAS1EnAMq21u8rwGIUZN4ZD/A
oQOOeUAdihfriXwUpEpORFRQM94Zio+NKnSjsQJilt1u3ljGfOMxvhF8dxzZ520F
bfhQabcOS05kFwmR35i2/naOtFSl1QSfvxATmwE3qkBaA7EZ3hkXIbSUjm4jYrc1
j59xtTQssvqXVe7HviUBLXx/LPvSj32afDU0opTVJL8JmUJ/jye+zwPFJi4uMO+H
eXx+oNDNks9LIT+xs2aEQcZiiZvEvMwQnEdJdUuVY/9oTxK17aBj/FM28M96XuPR
t7vlOMOEMhxQ3zwGhHGbhw1OQsfm+Fh7OuUwLmAKYWUsGDpdBB+cHnZgB4wbM9yJ
KXQtlgeMF+k85Poh/qPrT5GDW9h+iNjMw7n8XfM0T0/qMeuYx5GRvfPu1pC770XJ
W5eqtf05KF9swHbkBvPg9LghLh+Qll3OufipjoDeoDcb0TUO9XHipCKqbpQ6J8K8
Twt0uNDkMA2VDmW9OXsIUhipIOcOuWXfHcSzvlzb2vaKWdc5joqV8/PVgqRzifpb
70zVLVH8COe57cXSxu0RqM3p/5cJOt0VV7cj+kcONvbUYfWy3FzM9V33eAwGt1tw
ZqEUOdi9qKfFe2qy5/61LJwbwVSbaebv74KAL1EjygElye7k5ZATyExeSEjICG1g
/zP87KePFRzNrUOOTNSSnPa0Qbb4fJT8Wv/JxbMEUoY0ZFeOZn7lcacyvAe4XutU
Z2hkiR/+TpNaiPs0CvCI/6aC/lzBuvxswPGuW0uPgdfEhqixS3SlfEpvrREUQrzy
mAeE/SBoUFR6t3QDLOZ0MZVPtJNtJ3u/aJ7hTmP0CBRo1gOTxnFI643wQbv5WVNB
124ADhCx7TEquvp4ABUxg4R9bsLBFhRQMA/oDE3rAmkjhL5qxlPq0FMp04UKod12
bYXxcjyp1tiABNegVYtkxtMWI5aAA3k+r7lXiv9jWrDVp2Nh3T1CyZLk9ljBiCJO
tjjX13pXkYbQUQ4EIUCvYCp2qmO/EapteCz/wxniR/6iszF0MoMqXkTscq6P7Mu5
gcfJHmzefY9eT4iGyNtSJrnNI3Z6USEeDoJt5dwU6erxTimkd1hOMGwJNmR5gj/H
lI0gDrSsHaTJu28YaqcXDFW0Bfh3zeUXh5ywEu9iqSn5GehatMnyKg7VF5k5Ar3Y
UvuTzgh1VEk4yjp6IS/JxaUeZBx0sS1nX++qAsQY8DSi1xBaV9wEUil4szi2z/lb
GZ/R85TValgLyiiZQr7QOvJrPUCJrEX+VdSPl72Py2GDH0CQPLn+w57TbVsdd8DC
nTtV25C3Zu0Cl7dUiuwdx2qpc4+zVThVBmAWHhJwdU2OEZdfLg/hPN243Abxp18f
wAM9hwHS9dd84AHnFCaMRMZ0l14q3TLjkNqlXC/0rKZidL4jHRs2TELqBd6Z/m+w
SQTpuMQzlIIA1kCJdHRpSHt1wvu16xG/MUr8OV1PXllOg4FVgloLOurr6QZ5cUJ/
Y15cFwewW4xYHRdiYsGFH7hMzaVOvseKHANSlIB9UMZN2u7/Nt3qGMRU7M4MwRxG
CxkNOm4vs1Ny8Wqevk+lAlMAEnSWnn2Ce/jNvR+51bzn96Q4L4D3i4CBe7mvChKp
gdxZte/0evfcY2s0DYs7hQJGWnbjATN+8aQJyOBZA9Zz9hcVR8cSKOyiMHsuge4G
mnNeXnYsmzVFG3AqjfY+Luyz7+qcVemC2gYJ1NbH/0waalLEo+u8bDAJ3am63+cA
iw13p0WhEfaQVO/pvNnX9NXuQ+KNOgJEc0cI07jT9tb186IvoKB/RkWh0byrVYL+
liVRKcV2Vv3WdKezoUcJWj2Z0YPPjlTu10P4r1iS51B5WST1F9OqNFAbiiB5eIwm
8YkQ/WnHSlPqkxrdfNVhWA5OEQz5RLeVNYllVSmu/sSBwhjfw8UCoKAxX5EzXy2y
JR62Uik8HfnJQdiCxu4CLJc2hcQ6981ifD/SQ9Tj+TME58KwZ5RelVqL9hjmlMGl
kw3SD4FegVCwLNsFsLLpUcKzqGEqbgUjqq6QwThNVaAPx4vCcOQoGm/Y78Y6yyQL
1zGC3IVjvyVWr25hlyZG5PsgeWHZrlBehO1rz6LOjelLWaAvzY673vQmyAp1+Zs1
i0HrCs+n2sJmy0hRWI3/Xxvx6+NsRiyQl2AvE8aKXk4CU19WPK0WsPpMlsfsWkPF
Wb/96nGj0+Rvj4x2GrxydTrYddF3Hrt4QMKrP9XsjCRF1umE/VceLHNF/MnZYe41
T4pPjxAKopku4N9iisOax0EyCvKpOF77dxxmrdmnMmVbfdF3NDRCk6bvxdCdyB0n
C1ZLGcquasFutjS6QfZ+q9+OstaaJbVGZAZYL8FLIJQc+gtigqL1FrLs3iUhmEgc
GMzDzdfvyNeeHf8Xv6uFTZRMZRvKdvqQoL5nSHyfndogQBU6tBK5gIWLb6nAloO5
WuO3zqtTQ72E7lAk8e3wcFdxnwTrlDEkmjUD0w+T5qPbwrxZb3YnpjM95LPc2WGw
13JYX9t6EgcDQMVpaQOWmmlfTo7yH+SiqiSyY0jaFxZOJLwAt+G5plOCn0+JRgfL
ioz+Qck/dhdFo5gPvciT/rEAAunH1TMBKxc06D+A+8nhxLn0AgpETCPheZfTPaD0
3qQhANyErEmNRqNWyLdq2kcr5eaCcd3mLNsJqh/9q5jft5nxmdbXil5hZLz6w/Fc
oEXf3Jji43lecuiAd88BbPf2jtaHeEQm4Aw855yjsxN7cN3TcLzPo+KsGcm4d2XZ
/Ns0n+kddnBrUthdKVZKo2vTcXrKNKllfo9JCj4uCs8dl1aXNUpoR00WeE77NLFq
AxrGcRTVhUSjXa1Qh95jCn+Z6aHXuY0fpH1vLfWP1URcUXcN9/EZiLghL06zJuOV
zFoga7H9rmpe3eeyh7o0AYPm34Oi9yfFoWOvuTn8Vo+JnP2NkKFHl41T0h+jwAPj
wFeHuU+7x2KuCfeFQShdfLChf6ouIrZ3eYJVgNqlz9Gxp5B1iNl5HhmD0V6G+TNi
0gDV2H6/pq+FBaQAsB+sGnx8nC2E3BSIy5mtTRVFHFa7GzVX9n1yRBOBwCfQzbmK
L6harijc2FdHhpoWZU87M/yM4hxgO+56isLMpCAECig3GaZZwuKvqvHwbkzC2xeu
6Ogr+qvJu65tgWfz1PP0FwTXExvyc06SEEax12ZexglGkw/2jXfCnkpzTjeMAmwt
3Ue49+kN6tCUYmhDoWGM++7V19bfSrZEqEfiGBaowzii7wkIjY+uWuwCvW+Wg3i2
RfdQx/YD2Sd5+DHq6l6Z2P6lfzem5NmJtzeYFNZHU4W7ElY1eQNowRoenz6lu9DM
9Fd2NbypdZrWd1riadMGXpt3dOvWp2O/hvl25HLsTI4L3TN57sVsPjpCifte6MkJ
4wp9kfDV9qCcGXnQri7CqPcLdVR+hy1l/x3MTda5aiLbSe3qVzBUS11ikyCZ7z4Z
EdD1Wnu6KFPcvNj1HqlZguCGtl9vQQlt8GgH2oOq1AlLaOoUOkOlA/mTmgoAAT6H
U8bPMBdG8Cc3Do2VK+bDvQeEfACzzAUVSaggAQIIy57o5bRT+D1dXGBnQkuqVX6r
PrwBJUGC97TVm9BMzjtIQEsyJC1BFxAgkKGdIyZfgK82cWBNYxBv9ruJ7sRVEovH
BuiudQMGqnLPQWwVEm+bIIN1p2YVhHaun8vg41ibn2lpqjios+kv1NTnmNIjcMbK
HdMbXa4XENweNa7SSIz1evXMLIa30JbWSSz3gRMdvzZjMEZWFinfoqTs3CJXHj95
cHzJ3jILC2kCLxv4BRY2YswJ/wXMN1X41pTIzRUdcpZugQicioe8a7vWRCK8U2Pi
h3X+5b7tvwPrXF+KFDH316iBNMXRNskYFb1Fn6t+inBC6OLQGCjdms81bIoRdreu
IG6n/jS/mOfM8RYSvS0swYeULsKWSV1OP8canql8zaUg/OHITUeoQo4MN1Zd7KbI
7l1lwwIL3/2KBreL1f4AIPH3Yv97lFxdz/d0rTdk+KnR0hd5MkZQ+hLgY7+Nc0xV
BDhiEPKQ0uATACKfw0XMZkQzbqs//8ahrUWwH2EWJifaz+smAAm0KRIPK3nqtmcf
pqpvoMPxn8TnskEYEINq1/rW7WIELj2BAzKQHmoR6Qu5EeXTH2Jg4OmyYwGJqzWB
jDBcepAykC8/QTLsVhEAk6fSqe5/F1caBffr8x19X2cbEelbs2sCXHpZ0sykKono
IH6n2g/gcfJVckf7JctjHWqU13SsV+smPHULJf+OwGslHuKak7los2iQJA2tbyH2
ZC5Fl05q6k/EpHfMhW3bF2I52lO5LNwWsoyyxmcl5Y2WVLMh4imPVO5AWCmXkKt7
+VCIm/tFW0hEYk34yXDWeCNMjyN46pL1xJePCdC9hjuc9sfTpbEwt44W3/imKHAu
U0rivk2ur8NDZXLloAb7bjGyq1K0oN8bQR/flK7I+4GBCXpKwLO2CArvELws1aZS
qIMtf4uZlOJEAiXHcQdu76DlOLkyp7GEs7ULwra+zG1o6NR0hHAi9fdKwrqOj4Q3
Xhlf9aipDnxkPuFFJlp84NYOhJDBFbc0VbEQwC0Hl9ECb8KmHw4yThVDY20ZPhvH
gTK01EiP9D3u0MLx+hbaxrNL3g2/uSOcOzozb8l22QoThJqyDhCNtP4BqGz510iF
B+VWCavLHW6ljdyt7WMzTCeyb0JW8zrxAsUBGM7ZWGglpOQAg4keO7s99IzirUa3
R0Dfo/YMKF8EeWULbsrm3uPXmrImjORyRTBhEN3MFS87oyVYTvagdwU3tji5EZn2
drupquhGpmlBCHyh73HMx/BO1FOWf457rA0nAhObl5qSJTAbZTVMe/GWquzssNwE
D1PQC/xy/VW8dJn6mhQQxBO20cofHKYYGZhkskM2zSDxS2tu2/PRy7TruA0/GWHT
IYztHjCFBUc4JpzZlnnCppmltmbcMKBy689HVKdqxPJFA2fdhRLSV/20P8rQ2V2z
6uqOUEsmHcfZ3J3VHgag+GFHLplRyV21VP4mDz+tVITtrceFML82OuG9VvRARSyi
xat5UKpnq7Tg0BECgS246FiUxxfy5QyB0G2hagrDOd63sTIsjLoSm7ZTtkhz15Sx
EBPzxVOvgELKDtmd9PxZZG0HRRESgfhyMbXmBFzZJRXjnld1NH/nxxbH5Lvp6NGm
LwthBnjQFQ8KE0NGcGs6eipEj8Vf2x862ytGfmvhRhuDIwi6w3Kvq60//qDlTHuE
cv3mvNCa4xNwy4Isp+QAKoG50Nlr0NsECgkRu3lW4h8Yt2EonBTSlwRtu6Bx8zQa
F8f2/z42kDxAUM/KtkhhIxTIShSpBTt4oxr8BL7+MFMpQkgTgYZJ1vBT6Lqt5nQB
ErfcGNxjvJt5Di6zfF32oVTbL0h9rekXw9vfwVxLtHwjJE3nxkjzEvdOcWbq+ee/
Y5dUtm5YOHmk65ItYux6k4kzNNB0uZemnfmBhcWdVVpCOPecv6eJseJzp7oXrcFy
ODc//Bb5M2aqHMGKwMbxTWaIl0DaHHKn5T4lWtR/0dzXoyiIhTwLp2rxK0+qqAe4
Aq3UmKJGkoW86ukUR8F1zd14zvZibQV3nCGXMWkKuYCfvsaT9cBOg4yW6e/rxc2C
ZjwYPx9Wi8XhcaFHkZaHt/fijoL/EiH8EASsl9UydYMSemnxUiYK36B1AflI2Eb+
jAs1BVPJCFXduxIxWcLwGsm8NZQTTm3Q3Do/Z45CSEjQKiIqNTkflotaK4Xf6wTj
VeFbM+p8YPRgVwffjS2EJ8f+uJ6ScXwwUQ1he8QMB2/xAuhVDC22SaagmIqDeU03
pvFWCcrjMlFAoiqpRsUQkbJ+9uH9dZM4CfDqf/yRO9BkHiZG7kuCu9V6qpouD+KI
BT4tSel/m36R27HgT2TNn6jhUbSatSQ1jOOwjOZOtktOH+WTBC5aAspaSJnE7/sy
XG0t2/IQAiG5HXW2eV2yneGrN5hhnkSNQ9zPBH696a0NLYBEVKdpxL0e6yV6GQgK
I3+2okNZqGLW8MX/SW+H8+qthwOsAv65ECIrmUYHoZEX8qCRPySd5I70NIIJ/h2I
saLWmbSpTXLeNAJnp2d9f52+aplKDMK5UuSIZOGURlOqnxXuN0kWvqXkfBidZzyE
iLXxkYzPnwO5Ms3dMJwh0tMnkhhqL5cNVgYWE41NF8Edo6fqSzMprnVQK4rbYa2o
7os5GNz9E71onlrWDDYcoNBT6Ds9WU4rK38zplV55Gnp4HPLCHPxS4OvMcGqOU12
v8m3PeIMQbQj6iRCQOKRU3+Sv1/vW96BSHUms5MpCuCbuX7S9bOb/cytiDDl9Oi/
E2YHMu3jqBsGQII3aPlAukKijl06jC+1JiHqjub/wVSua+q4yXdbgpcF1WdjbSXc
wTP0zYdwAryGNt1B8/CIz8brEG5QhbKFsB4YZT34FoelDL0+ExuDZXB9+Kw5dukJ
f6m4MiAHhMdJQrEuW5yxD18h0dvsB+wB0NbmQQLvWLYKmOKkeWu0feZytwmGdDvR
O0wA0A2JK6aBHosq2woC7RRIdg0Ib7eEvgw/gvHRmYQ1wgwo/M+Siu3WErS+4LT3
/wZCIToV7BT/g7lsqDiIiHdLHC/h6N527NZYbXaAzLY47qgHYJWfHR3AcrrRqDW5
uHH2bo3+sBDY0zCBTG5sRHizpXHXtd8NA6rIC1kcIAhLrST5ADbnRE3qaqf9z70U
IO+8dduAMCb9Vhl99Cm7I2rwM2ejC4f5bUcc9t45AmOmojlcqq2mqeHcKIcNxNJT
2jjbPzaN1vC6vLldDAcRfjYGdKDIV+Em2CmP4FQ50LDrPPoRWkqpfk5q/lIPwFDy
HWKjj/VKMVZVEaPeusa2mB9hyBozOQ9aLgDZdQH72mz+l+UPZ0yIghucGyhwvR9T
BcJwhOPVomlXvuZMGjbbuRFgk53UywKLPVsQeiDfZ+EuhreLSm3hzCKB/oW9P1ut
9lmxbPl4CBl7qgKz9/GcTyAeJRHXPP4xGR+7aYDdB1PCAQq1zAnKuqYV2H2pgAVi
KLL7HuiaBwo7uNkHz8UnGxDSaVFmKK0Iq0Tk3As0X20h/p2xJVM4wp/N6Wx3pz9B
DFkJGaNLQM8Wczz0MLtmuiA/1rVcBuXazb/YBhYOmXjrF8PdFpW4jEsXIhIBIJrY
9FB0JOzR8sGJthDfP52MQLdk98zdgp6sqdkXARq1aRES8e8/ZDL8ccw2rdqYOJ6g
5sZ7LQkjiTeUua/C9ojtWeBKCj9aIeU8CA1T6Uv3bCaeIApI5OH05zEerek/FBfi
lsHFYgDz+MCCs4a5h2J6TXjw+l68Cm/CNMU+5FTV4Qb2xAFuGnOeD+QGPm4eRmYz
Pjkdq0D10GYPoYDGFGKWGPsf1ywTbBYMrhPHcEeO4NM1dGUBeEpS0ZYEz2X1r6OK
uV35jth/VRS6d6oSqxDmVxmupsVb9MOQ+k42eaVhLrDfSHZT69fArRKR87MwjzC+
RyKEmbHrGNM1sHpkQbUe+gBip/b5RNn2YcyGenGe6cyI7k1GUJgHv/xLaqNCe7iV
d1H9TqjsMkAggY5z+Jcvys7EqoGuE0mNMa5EQKQcYlp6ljpLDSp66+a8j8REmKqI
T3D8sCbjR7i3EWI+VmMDOyZwocMZOZvVTZI9zr4yzEh3LBg2wiE5HXe4hm60zUEM
xg58GDreQXz/oHY3zjtXcGVYQ/5qQUeg/ZTL0jj5+obUX4oFyY/d9q4WhzVfQg9G
3l5nqie3Oi9mP2jQDyonvAmbeQuQSzw0MM3+qil5ktbI9FTkRZm0wGv9chh9zDjN
fg8ZyVcbpCXQ+qC5paqAPX8/Jw5SI/BY98/8a70ftDUWVSrjubkv9YPnxiTOUpL9
NwQ+ypSM+mWXSvZjai7EemF71/RYey48AHzXBop6VBfTV97+JMKc+HpynHlkToKg
VK0D3eB8gcWyVYZBGJH3lHapa/Chxm0wzY/whR0N10u3xcY+D7oSobyV+y2Y6Q5W
QPYSjUqwoWmc7s/39Svh38+7LJO0d+R1wwXDgkTOo1uecYd7gyKkCWXF0Wdca1Xp
HJNTYNw5CF3IUn4YrrP6Ba1b7jNyD+7hza+BeOUY1o9OC/Lj9CIeq/PLesOXNjrx
FRVVjttmCqLMhZRcQrz0IHaOVNl4kwVp/hJRN15QNVQREC6uhufPUw1S2t/AGlWZ
ENi9h9Qm9Z6o19D6Rl0Q8ynWrSbCr4PCzzidAOJ5u7maOem1LvvVyniZbzyk6hP4
tmymsSP2QEo6+AvS/j/+bnWYytQqqQ8okcVHFitzcVF8JL8JtD+kQL+KMuZ2lzRQ
u7R37bSxcCCnq7pJUdyIADkRTz3uz2a32eIGJaH8S8D8pjiSxd42KN6+jgtsS2l0
m9iUNxUVrCyJg7m+dKlc/JnJ0ScLBXTdlQB/xgoRaYj38fd3tJlF0Mht5yINDKL8
sZ2IdQ1pVMRWjpoh+1EHJ5oK9R6gGFzRPtEHCCFnfojN2X8XMISKrulg8L5lNHj3
a6umXdW6kHta6x5cxsAQFQEyiFSD/k5hP+OhOHN686vt1lZVGGn2NTv2doHvQ1mo
jesxvfMBD9qpjDnfjCmDOnB/3/Lo1BOP1FWkxh7Izvd8X0juIFBWlYCh2Lev1iL0
wN9Yz7AX2kQ2NaVGPQ135eUqaV9ynZvMBvS7Ut0odGuG92B3QvNBMVFf8zNLUZhR
WNWiiYs/SIRWzD9B06FDzVgRRdnoUbikPWif2gsOe0jo6YqIaZCaxqopJRfcb+cM
R3fTlKnlrg3ab/dcADJhwuYUrmpSgbtzIeQHrC3vKj23x+4CObAXmSCGBGVxVsT/
ld1/jHM0jYoNyHX+cYvDyvtP/PgVYfERslIc0iI854Kzh7c15nJVd9iXlFC6K6o2
+pPPRG1O+IQh0dT8Rtra56avohCAvlory8FQjQWZKHV1wuv5E5nqmHe64XxlZ6D6
DQP2f0Cty11YcZZJWcBBAu8kYaXcyXsiKD6FMnYpCsaFvv4LgZdtXaG+gnRBW6MS
bXtQlia3AVIH90HXM/W5Anhm8Tj5TTgyZ1HILt8kfExuiW3BhX+phsHQxuYJd+KE
Sz6ySogKyDjZPLZ8eURlx8T0NbB2ntppNQ1Ych5jXtm3iSYx0DxkAZlXlPViV7Gf
Qnz8THjfxfcW99hqr0ioIzM2vjyESfX2LFxU9bC9z52FzvTmNhdLb7NrVu3uo15F
eBcAmCSzeM5JJZbhavvr5CrfFryUNpLdKwBJxK4cEh3d/RG2okYhYJp430F7bKjK
YkcSk6D9scuXOQtH4LNEY6tQi501YBTlFeFOpmR+uVFoqIiHV/ALR2MISk3RPhKV
+FoaSXJmA/5rQeHGmCgwbhK3v6jcEtpvRvsRrD1xbK116Xcw9Xj7DHy5vtoiygFu
C1k6HwybdJx4pzmU71elHYt7tfIkAgvORr58XaJCAg6ctO6abOH8zIJYuKF8ZYjQ
wbDZ5f3rG2qLuhhcVsekZUp4g+VBHuO1M5Ao5PfyUILb/VPFlOZDFcl3sgKBIoBr
3yvmOI3kMx34mqxyxgJcl8EUyCwAlNY2J/BGbVrTcrw0kxTI7cEPZligSLUVWOSM
z1MJu9IFrVCN4YlWML55403BhBlQ7ofeLYdgXC7LjHeEiJX2KGo7kFCInUWYcsk9
JHD8Ojed5I6NtGbZDE7TdZcfbVdMa/d3zjBop1MKpN3MrcfhUzq0+hF2KYAqTfsT
MJ0ivUmb5+hrcbrV2NKFZ+KmyQr9uXT5RagiPc+vHQO5kd0MlNyUSpTsg42KSacg
LVt5W3jWZQP//t/ZvQoXh1dvFMfeFt4ttgPalcNQKEtiFDAbERC7xpxqUpqwRhuE
wGEghBOryHwzSKKke500sGOizBY9PTDroQjkF+24+rjPNlgdsFBIuwTRHNoOMkpP
Oiz6b6u/mi035Yr4El2YHXmDZE8Nu+9MveXVsRVNZbKS1AMzRAipqDWcF4rEw+gY
pWCCIyY8JcAetnpop/2oOpUh+9MwEPzOlNCZ+bsY+8n1u6MeUS4Xec2mT7TLQMO1
wqSbsEbu/gDzw3lBrdPVNdvOM6iFE9iq8egaPoq/3S/0XS2LMBxE0feHbgoFimO0
nVWnqKQqNVFT7hMj7/PA1OJIccvUcCqXy6EbRr/EvDYAwfpc9WJWlya4X7D9hWBp
2aFZ/KluT3nS059Y9F1c/vYo0d4Yc+6MGefnkZPv1h1c8JhmrPR41Nl0L1FZlSg9
Z8z7Q0Gn0tXsYsf6y5+TFjlE/EgMz5ZF+dZAx4YBdZmtAYOnUvbMiA41pPajn9yP
K7SWqNOfTiQAvWKrMGnP++ubKNSCDcSbOz8XKR+BjWWsSZcfKOVm3KSuMCnPF/tC
4FX2LbFOyI+hK96LRk1/r5tFlTIihKeCicnsJGQYsAm2aaw7TH0lcU6hYejlzDEG
ATV0J/zmY8AVCox9OQR8s+oIZiZnmmp3Mc9dGkWZExz628CrY3nXcgTcYPy5IV/f
u7uNcHMpaAObjoDK86jA+TUERct1MIt293DMwcbb09lZ8KdKYn8RRL1KaDirXFSK
Tz+OwT1CeVrLXUA93r6za4cJUXNBMV9lkXswa/X3Gt6zQhN/vHYXUBOiB7JkDsHh
oM6shm7Vfn3CBkeD8+re09Tpmu4dRt/P+AWlcSvWZAU0Lm156me9oqLIfhHkzCk8
V3Po/aepfnA+7cqSxZoOG2e8ArcO/Bb8UTIgJj7MVVfzB4njn0iWKJTNzgL6T1ub
uXdx88ibrO2M5oJmPTCF9F2JVYqbDy1Zef+Oj7KXASKgCBDLb/yhmlyZfjwKh1i0
aRoK45hYz99+otGgif5BQgdV6OJfHBiR4ySfzoeqk3duDd3o39ZeaTmuKwGMvGHO
Op1fuVi5QXD2wE87/SWkyt2TxfrpW44b1VLnroy+SPnZa19EsNK3GV4nSkdIg/D5
hUgKoUVFTPUeWDZ58K4pAVQ7pcHuvq4+Kibq8cusj+0hFWhyReKWf9TOeb9Z1HfF
1BjyL0U+9dIsaHLluM/fnyHro00ZMpScevmQapRDvrsCX0kAUUQ7/5CFr1ogOT/m
0QHXM7/2Q5N0JURlVmdS0eSH2C0LP0YaZOZ+lz1nZAJDdcLWUzhbh76sFjQz7Hru
qUlCk0gsnvgfJwXTyWkIAXOI9Qj+eOAzJfqoPBJgtRFgxfGtcEtqA6rWGC0Alv63
gfjL+0+4b+ThEdQXaDaU4g9TT8m0S0lc/ut0+xSnBb2jgVv7Sm37CbYBQ87JMCRM
XJeYfPGBFApeVcGT05SCJw5Rr/b4atuMT3qYOdRhwvAsf75mo0pNxpeJF8SfQjwl
EM5X9z4y2VYfwkGCbP9IkC69Bx6phEaxL7l5w/iCFcG9QWlNB8LsDB/loDNA7nBS
t1VIxW27nt9tV4NzaHcjxhtp0ETURuv1VqQ8ossIYy6eorQnileCSN3S/BAdbP77
CtzfDZ2jmTtBCY+g7F+Ust4hHPcx488hzjdVYouXHr2TEpXxSAtzox3cRQu3uRz5
obtDS60gvx4l9e64RfByJHyA1mjH5VCOwRZ+Tn3ebfp2xyY/NU89zpuaGnJlW3TX
XyiN4z9n22KD0FWGZNkSIOmIvliCRXamfXLuf7vVSDr8w8u6N/BORPrEiWtRM/ZL
DyDA3B92ZvEZXTbLMZV8p75VVxgq6aAfA4kKcs0szVIA+21s671hIMU+61xS9EVx
2zuN17UMT5xzudH2XauhOPknQcjWuiZNm8lvxFbXGq4zGAUtsHEwfnX3yncHAaK+
EUXyFcljNFvbQowoUnBADjsHMGTJGGmgaBHVSF6yRZqZjm+iblbNKVIoa+eKhPP9
KDT7GWaniLig6Rweg9lX8cIa7oCfODFhbXw+QiFE4ZYJeGm+KISeFt8wiSAx88iM
yfDBR/LfHfxtkd0J5bXvNlphmKghF5Ea+1/lIeHi649G8+KnMyK4i15utgY22flQ
LGUeSdltoCrOs/TzpC6G9mbxWynKdw9rStehewlfgzKDs7wvsqhZusNwv1EpNk5O
6uEjs2LwNbeivHgk9aJpuxUM9Dur8e0+0pys8pC4DmLkiqu6D8FzywgmEY6ykt7m
eEE1ukwAr+itG4DykOFaASJSqZZtlf3hgBUQGUJIRFnnbiOrnoFSRTUBn2apPR1C
E3bhAqRqle6fEwevTM5dHP4wxb+XVLyG8FFHPWaR3tvBvKXDlFhObKMH5uqY9E4W
MxFnv7KLzary5it2RCDkI8ZoTCofEATABwjrPtSJCTAPvQv4TA2OjG02oEKRQSJk
QdHIv3wMzQKwcC2lfAA595kFzH7kbCOMwQvWS/AUfll5JRQagyCJDFeqGcXxFILg
+WBJ53mHDWoptM4hsW7SxEufJuGmp/NxXeuwf0b9bxnfy8aXc3qHpbAfgczfc9FC
dJKSPW2wKDV40ffOzd3UJ4NyOPhJQHc9BvL0jbpLDMT4uNNXo4jDJ6kUW3vwqJx1
lJaCOe+sRQzdUQgB4BCK2x7IFtThHqYi2NLE1m++pleUDGKah90tHmPAWHDR8HTU
Vy7cAfxzczGd5sssdZSkDvQzciIH+OwP6ZlTIsY8Qdh47TFHvCFc6ygrMLlAQHm4
XB6H/Y6J/rkbJH41vRmObBYixD39TwuztQqwx+S9q3cby/qaDh3TTjtxwKSGvG+5
2nlNUKnOb1+I+6eNZj7gnXC3fmDKsp+0QlVWdimi/53jsrZ/0U/It8/Pam/P/13k
AfBS3nlSXFbpZeaOkN7zd4TdjjC37eZM7zNuiKKBVer63pjKHe8BCY9gSuW0F038
KuyYehoQjFcGtnSSieLftFMWz3/O6wWEsnnCxTv92MGnWghpnuu5x6fjmX+MBqNV
4jc7HOLsNWLr9YIkFlJN6+7jICyhmiN301RsKg0KkTVjexJcziCrOCoWgTbc7HTg
reE/I7pznWi4MoVmsrD8ICdY97v+kdPlLQKaugQuLU/twoILWhWz2AL4SWj7iTyz
/TCVuYdYzrZkz337yuSENP5mauZGERJQNXYquPvo8jmjU/HYuI4A+ySPrT0k064T
FCV4uIogVg3OeFsdWr2NbtyVcFHsA4+gC8DbXvtTQKZWdUxOKkzRsILGqnIC8a4p
XywVefn+kWyKJNbTfDhgknWat3E0jy4o2drzDYeYlpdxAgFS9ndtHMAvvS3zJnEz
7GpbXFnI5qENKIfrRiZFET9Q9fh7xwckHgKpJGNsRd8x1FLZo6/hDEHED9T1twIU
JwYBpPP7y69LopBPv4mgwEenlNlBjSsQrKwlluc5EY4Ge1i+JVNNMQFIS316g95W
AR9T5vc4vERvr3eCpnYOZOch53u7YTqypYJ5oy4lYyQdZyn7NjbCN6PET9qnn7U0
N3m3lYtnOTmRCNTBT6WWfndxKpVuihiOhgRosCVn80uV5fxw9Rmv6sDU5TdJlKJT
xsewIjkV64LGmT1EpXiDH4xCU3j7hw5++rD/3ZFQTFVMyExYOZs+3sTIn535R2WL
OPapAn09RRAG88oEzNhpULNDIGF75NMvajuDdR+lPqalYnB9o2ffoTcYV7ExaSvn
jp2XtfZgWXYSilJudgbWcgIjQWFp8Fe8HPzPmWNk1+MaT+HFj47s2X+vAMc1yB/v
t3Y/wFKBHEj7FHUsphmmMVpTHhpk6NSRHdnylWHz43czglSXFoJxr/UZkZeNusqJ
0HqFSnEUxQFp+01OOEvVVv6j5buoQwXpaFQKAWGlpmt0nx6JAssRShAxa+HbbreB
j2yS/cbymw8gS4kimktuFm7ytfjAAuZlGzAvF2BgUG1lIBMDVyqNR/U5fmSOsWhu
2xWr4VW5crwEMY2UTRdX2JdJNeX3QzKI893gwk0rz6mpoFU9HOkt10EbKWzpRzvP
tEaFyhkizt65DrByXAOvUEkPiRWT5gRugO2s8JXio0MBoTZmVG+k1W0w18qBju84
HgSn8y8BWm9Mk4A3IPYZ1B362hua6VlcegnQ7A6iemN9JW+Pfp7yUQZ5Ml0sojY7
xmXcvfk4X4JT+Ou+ry5lKRulK0PJwROURfXf2o+2/ZAw838Kcn4+Z7EvsIAQCQnd
WCNuY1Fog6VvSPGaXs3MOJlghOOPVdW9Mn3237tPOmzUnRu34sOACM4V0BjbjjOB
OrrtpRS09V2Rl4PLuTykMmHuipaYXBEKu2vF5hK7JZJ+YCO4+fYy8UNuPEkBTa5K
h8taI6l+unSyDfmcwYfpw/qAZFCAPwoc19S96AyC2qR73r60bALqinoKdz1LGtOV
S1nOXKpI+o7zNcKWWqaQQPyc3PxPhdhhtSXFm4RheB25lu0wRALWOyRkSuxfAarw
ARPr+r78ixA4obPqvIRmeaipmdeVvH1LuJipcfMjODIs/MrEpnAy+JI7itPOFA7g
kLuAler4j3g/Z+It3svd6qqS5IR2N7l0LXMEtMoS9V0yt1jRtJGrLHykjOtxZbc4
bxg6nr9Vn+3tOGgpHwjAJ3CS4Qao1pdxyVgM6tfErJ4pfoaXig+GiI/grGnnz/Su
7U6HwO7EYSXtwavy6Z0pczqUcaFJadDmDAcyFBCFvF6HpMsvZpqxrMyTyivFytrL
5EqR1gOeaJ4MOJHxTJVScJehZxT2xZZLOb2s+eN6F0oSNQ77UFhFrmOrkl4Z3oHi
CSSbWU6kpYwvwA6o5X4iJag0mNbNC1xr2SyTu6NN8cK9Fky/pH5wLGelAlvtR+1H
H5tei7gnq6LOsLAS+7HmCFMHHf2Qf0rCeKwAdtB46gTynKSMXurYO7S12ud1GqJv
JuY4aUpryjDv4881QslRdEMBbNYIPGLRnewi+2Y/b2bfhLzqQE7Ygs5ojqLOCQVQ
+5+HIDmIDx3XBBhWXaO04Fj/V19nsl7juoRwoTKg3rVO8atQOCJyh9M0AVt04zxB
8Qr6jHbSirmb3DeR7DmDYnhhFbzYpg0s9t16Md1qo7DIzJ3Ogf796MDvXp/Z/2Ep
rwUkkbZZMY7ZVrounYihk1II3koJusUeKbdYCD6cc5Y9+vGRyphL1Gx0q01oOq+Z
S3tM2ntHDEQZMvyevm3j1WSu803Oj4acRDsjyoNwGCRCEdJsn/MPPpXSEPbOk+nc
4sZFgvxL5yVV0kPjDIl48/ORzcTu3kVtXxNvuxAC0xGo6gU4We7yeNtsUTTyRO3X
144WmCobcOZRSRyoYBQUHDVqfRl2nzNQuvS8j8Him6JimneOeCx+Mw9g3nDzkxHF
QXHOasPlGt/pK4TqZvWYrxP6+mW55wYGcXt/n1dIxjCMz+qaPPulTdmVnSkA8RTj
DMYLmyeOnfIQ4x5bzm0aAeGny8QAeD1XxUOiVYzHSuqpPkS4T4IZUHGRGW7cbbyW
1ubmGVpCfbZdfYl6nX/6GftP4UaeMgA4plTAgLBmxKp5/qqNtt9OVnB9WmhJyC7o
Ckh9cBhUeQwGkiA7/EjacTcIMHz5h4nVh0eu5tSk5ZHaHm/n4rlyQUnFGoulnOUk
YgdRsy7jedqd7k/3o45p6IkJZmgDD+86hmZGJVsoXOLdIwmCEEgp0Yl7qX5wXNBl
CXqEaqFcxXUZ/Px2aHSQi1L1n57nDcdkqQ4TWSP7jLZoiwn0oM39wbngKleLYQab
KP5aporKVUsw/cH1ZRmcU7MAoAaToGjUnrCgte6bkcoUWCeF3px6cvi4GPm/GRH0
lNichvC5x6rO3OuMohqQYzxRwEXbed9oR1/YJVk5Fjtu47co6HVuBMGjT0Y8LyQr
ePUuB9CgieQfDpox8yFJvkCFWN6WEk1BxmvncRYiPCrVZ0f3ByHotd70mqNfASKZ
jgdaWNYEJihQeBFJvHbjNe1UQQ5Yb8D/tzCbDiQKnriqZhtVxyn69pllpRZqyIoO
FTcNxIa5ei1LcO38K4aykteew0Dos9VK0t4iahZ3vbbd9ZyZUvaSrATPIWSHFJcx
MmgELxWcZ3g3ZRmcGrn9ZGPX+YcjYbDR19Ou6eTVcYesZ0xAVc0UbiiyCy2wkvP7
iCd+easR+C33PZtf2LjbqHTcxxRAdAzQidGaqrdvZzxQqONVi/J50emO997x6RQd
nC4XM6HmrLMudIkm4yy8nZ3NSwVU/5vO5PjxRZfsaDDEM68QI91itjnyfBd3lnzS
xdr8fSk8KM7iV5wlQOigHzGCxrBpMtUZEtgpJhpmlWAMY5b4w+69dkk7sd1O7I75
3w8QBMNv5U5hp5x0v4tgPankffe4mBlhiXy1oIeo+rvrk8GhWQM2nKHrx+X4WU+d
y1mYH91vYu8XBvI6zM8mGBP+tz7GxaW3Q7LaP6a/hTRxr4KOmWH2RxRDMoZLUSz9
/dpfxSGlDcbdW0nmQX4b6CJV1obJr1FXABQlm2S34SDhsA6/pD5/AWKj+AW1eVry
clwnpbmH0j9Y2Yj7aH+Y9Ewn9NFT2K/MvTSOF/FC0IP+5jxkn9gvGmGEvuZozygK
H8at9BwEzFi9kkgsI1nq+pBb/Ismr4igbOYecOVtik96TVN+GRudReF7M9xcnXbr
1Ve/HMHBHDKxkS/A7rvXXfBL/fUpKKi6wsmM8unOHM6Grh83HWVoBB7w6TNz1oUq
GLlHDJ/L2KhJQwqB6s17z2B6f7CbwPXgWbHYz8WZ+Noh2NYSLWf89J/RAfJzkPMK
5OJIMkAmXIS5X2t21r8YiY9UWU/nIQOET7zeaFXg6kLTYesjsPIpr7eTliL/pztc
GNDmTk1Tln7PFfCCg1gSEHSsjhOoPlLidTIV6oK9BB0e8zxhXq5J9sGO6pIsP6CM
/6mc1AlZfE+0EfOIk5+Kheb0t850uH+JbkqbLIPxSFQUbleGkKUr45Lgcs+YZQb9
5HNIRJ39MpEU31zSiq1kktbbMEPumkcuj8grcon/3LxU5L2vdq0K23M5O9Zsf9Nr
x8I8XYQUNSDcKYBSosqox09YcKbotNlCsiPMRiqBzvgEgU7RpE9FjA39dTJ17m75
dC5O/pSBVvWrui+fieqMWTDzzaRTERghCFlXFzLlkMHTacwyOnBHxd0PkhRtQ8l3
s9PXBAHNQ1ohWqocC98DcXVygiLTw2smQLScXbiI7Xy7j35MjKOpqFj65lXaeUmM
vU4vZo9KtA8yod0xtTtFQUfI9PWW/aBUeMmFETQCTOEmk2r99KZHi3rlTf+No4bM
e+WWacBo6h/z3FFIJ41pCSMqjoLZdKgIj+gx7F0MIHInrPFVZ82+tFiQX4Nh9iXO
c0cBU1mzAFTr6V/Or9BbRgoPeCmFOo66N4JC639H3OpyXq4FgNG61rxqaNCtQLTK
IzQ1BRaKovLtC0/2lDIzV45aGGtoj7wQ/7ySPXtGVYt5Bclm7HTx5aV8ePCdYevy
5KxOm1f2W7L6ad+u2vGtz4yOw/dhfXZV28A9R9idJjh4kD1gtyNrsmjT3o672YsK
fEs03TgzQwS/dHWPsxxm5EfYPajxUe1nnOEdYTaUX7s+Q/3E14Sv2p5/22MxE1g6
f4erQLdmoriVUbCNX+XaESIrvHTx9KJYZTyZScpsfRjgmOPtJBDkj738wIIs0XjL
QCeYa3v/y9T/2gmXNB/lM2z0nu7uLZbZTBKEHX0MC+RodjoWclvJwlfO3xAt8ETx
eFDxba8PeMzOiV67iQsv63mK3EYA1v+tGIrwavR1vjPMSS965wyRM6Z3UUDgM6tn
10DgoAVp0L992DDbUm7qsf+SbbomSCv9bYN6flYt35e2eKaEnJJe34JZlH09krzj
wrfQjo+uA9eHpYMgRi6MC2GauX6U5C2z585FcNk8Gk79Aw+0rOIJ/jLPmBcklWOS
7W/WNpw3SJifcpx12ZjK7yjK/Rk1+i1RTvemRNAawbHdCRJ1sSbCVDJOP2Vx+uKU
fcbfZYTW0ozck4Q5qMCHB/GFEaC5b3323AeCB1YaFNhLiWxj6D9klfonLNMfPNAg
PEETT9tjfc2+eukqIztqwHKbcN2gRlnb+PU+YuEKaPBXom5Aphxdi91GckWkWNKu
OgdOFqoCLCLNqBujXCnhzErA+f+ICho2F2rCyUYz6evqTYPNHvOzBrpAENbR4ZbJ
r2pr+sMGMGVpxv7NAHcMIbVRkzFJSbW5nG2ZglGGQ+2jsfYCC7CCT8el4bPKwNYn
ITvx/Gj/rQ7co7nG7PnCluhp2CCqfT6yX/YdasSGO/xDsLXSz4Zsy5cS8dF5K7Xx
AwQOiVuYWNLWPU03gPzXSGzPKC88bnB5zbOy4JWkPFxwpfRrCtzS7inax0crzvwi
HfYizoNfpCxWB6iTRRk9SEU0vq/a6z9mKoFUPJX9wuxxrZmEczjXyC5BS97H+e4d
sUgO+vsJNNrgaK1hlQyV5bHk9PeGAZNEkOVxoCSJVqSulSJ1Md0YE0DhwDdVTchh
pL73ZvFMHAh6F33D+3zk8RsXh0i55OerrONz1G1CbYrTIAsijQgObOAkkN4Y/m/N
uT8TRIT0lQ6rpy4OfX1T0qtcMrYWlsJCqQ2Wk/N8ADYhiNywwPwfUDxchhkjWDLT
6uD1tGNlfSuxoRmiSN8Bx1OaW+z4oxxmvEg76osURbDzfJ1a/GnrrTh0CWEgjtPR
HVD0Qo70uNWDBm2IN77bBtDCHq4dqZktDmkYbZA/eata4MEB6fflqrs8t5fT16wz
0DCUbRnVb/IRa7iMcpYkxY6RsqJYVoG3JXNefkm+2/U6VpjgR73/Bgs3Y1oOzNAu
ZDY1E6Onlp/aAxL2g+iXsUEp4PbLylsq8zZIjIr87GB/65C1TSWPyvgnYsTBc0zN
4SgglXqCcwcCC6Kxw1PDZ3/fvgJV5D/utt3aizNmIVAXv+uT4DQN1hhZ4IXefrkE
Q/U7xJg5L9okDVXDkOngXQjiMRmT0OU/UaQG8jua0eshIHUuWJhdoWJATbNA+pY7
FEe5L90RC7b6a7Ynr5NKhh8HIMmHyWuc4PSaq0ynLoluoLEuwPjZSjeV5R37fZ+P
NFoquO5KgKGzphHzz5P7S9mbixrzHs53HPPYxnhl6OWrUaIOrci1pts/3GD+WwRK
qIWO0tjxBgUk7oCYNBLZ3/W1+940GJ/O6GANHxiQVXGUUonLGQ1iy0lHh7oT87T2
fJOGofp3YpvWN7iEQG/p4/ck0enSTl32uhxd75yCamJ4JvzZyX8dxVforubPYh2x
gQ2ZEMNGYF52NOrvwDKmAd4xKmCsSddn0Ig1SSVY8SniR02oeuD28Y5QqKfi9E0U
Cw8zgU1D6a01PgxI3Em5HJTHiKSSbYJwEwAbeMnlFmfVLoIfq8HHffgy4WdbKG36
Oxm0WUxVbW/V33ABSWRefSuOTA8M61boEkO/HSw/g/ll+wBMEZgELgtTNdO51HMQ
9JuyWl2uhJeYLlUZ9utVNomSxfzfvQiCv68tsHVRGT6Y8WgvHbqdqFUK/1G0gYHK
Ox9HXi74FAqtoQzoIq+CZ5s4H6/PC1RDjMP/YbL2Z/wuIOXZUMTVVxtcLE+KigFh
dg/NmBFgdE4COuRCI00xvkiJEnKzWAsNbSmKX1iY0hBJ8X5xhRg8wE9dElPjtvpW
HKgSwR7GJkZRMYcabhZhSiMfrfnL/r1YTsCcG2dzYJRBOILTFWb2LZ0Vhf3BsxP0
fn3UF7NxcgXk9zuYfvzGyO37P+YMbNnFsJ1YesF08u0AuiwzwGqmgzM020Q/OsX6
A59WdDvcEF8RXJJCeHcSSeEUA9r/AewOym/A7FSmbIDajr04JUahkvBKH6bdL1WC
e1S5SA9QqTTU7OQp3GHtwC6utOVaBwwxboXVcn6urkW5ikgDDaxjQYy6jH5dgD1l
+mEc1PcJgB8KioHjf35d1WrR3N0ZvuhT1kXCnosJz7w/TkA0U+rDkmsgHEMeNhSx
2Zekpjdj8mYteN50vFGoubvcIdb2Dayf8FRr59A668b8T0Nc14ce6JviABcyNkog
8KmOvEel3GpVzsUuPDQc2Bf2ar45E9bxyLJOW4NRARV0sjdtLaPSHzIc5oUy+T1n
KcOqgOyk4Rw4hBqylM91CtLcOkXhCWU6Ctxk2q9ajRGmG1Zc5kSY4/BXZsfyJP40
zZaxGN6dmBG8V0UV8FYtAqcvsJJMiU0bvHZtjkwLiXB7U0EfUZlumW7UeBsvzq0A
Z3A+URDrlMQecT/FHee3dyQinzOh84JefCiFlBJBv2XAKyljeZLNHaA+jfXAMrgW
994ovwBnelT9ni/+NYhOL1ha6WiZFnhOmQt23AnTGuGa8jn0ROchxPQW0c9eYgKB
MrSCE7onuHcm7GB9dROYVJwoE4rVVaCUespLJ5yaLfQp8V2Hyi0M9ZTmdlkMbHTE
eATID40LHiyhAFyVHWqngnE366GvQnr7SwaAHBVOs9gXvJdM/x5xT4dX5T4/88TZ
9Q4O/KE320aTMOYNBjD6xWEt8HgzuhrQQG6PwLTptZMTMrzVetzO8Y7i6MQOu7R1
9P/YywphMHhpXmClR4CyBMyk+fXZ1S2RUwm9J2rhF/Va3gLU2FgWjxYyZGCdLHWE
FyDqRA315r7j6pYSv4qCpXnu1UpO+ZwLyGRdQMvl48Xgi8iWLiGnN4TA7y/BQSc2
qBmhZQ9dVAVvKcABk3ZURFq2R8hXupPYLS/kHube8baLQ7OuoWC7348BPU36y0Qq
8/z3/kJxOGZMQqAxlSTQ7idcXko1fKGw0q7Ve+kc5tasQA7iB8Z6/IcNm/vG7yWB
+VIakhO2icDBMwUcxPHVe1k63P6CSBZfA/xJTwUdVVC/Bbm3yTImeNcwe6GInnTq
DlBCJL75VdObfus489AMbHQqfglx7oDlhrN7h5NlyoDzlIz2XN2s2igvDTdrrutx
gElsliktCX3CoPoD0BCDqNOcpMzLS5d1udjxfIItLQEWpuBPB1JDW9VRYlfdIHBy
hi20RyYoKWGiswqQAgvQjG4KHTQJ+Ru1/Prw2pkCLBBnxz6wppRoK4a/wq3ge+Jf
pmtmWmo6Tw74oAlDvlTTJ+wR96ssYPMIQc6hJ5OqBrztL3MY/YVl+IgYO+dsTuGY
VCX2FlXUhGi6hoeHdNYMyIFJp4Jdd3/6eLz9eugnCTE8hL7u6PPdRBBW1B/cIYyq
LbsGm25njHCC0kt3nwrocK0/G7lgSSiDfyzPa2L332BWGJO7/0BSovKbJ71an1GK
FC+RDmD+QSMqbqtfBXKNz3dEunmz7XUXC8ITGuyVvKsMMrXGKwbOWTl/GV+tglpS
ev+fOCDdjn6AwJvP4L6RLDNcK7cp/+yb2do+9IdfvQ0qZr0iUMyDXiFeqVgNoPj1
FhD3+hjI2CZtGLtHT2hj4SJUVkdGFRqQ1Om0yiBdGSNPHd55KtX6F6Ga87CPpetd
vkRgDzJ5j1b8vT4TTofXMVTuMXqWNtglw0bCj/9GMuijNkLw9dLipNznlHrZJlgu
n5SyNB0UKkbALTuC0sSP9ftDjw7NJlf6pRFCee/q8egIOd8SAKHpEinBiig2NSmo
OkolIo4DtvtI76rIOcTkUQ4CAc8xZp/9G8e7HT/lLinD6tsaU18bZZIsMk8KNjz8
icZDe47Ah6xkcz3rYW7S0R8xaxCM4+94t5qlvqcIpENiG5e8ftnD9J8S1MvRCVek
CsQ0JLhzAD4AkG81THOKhpcL8PXBMcjTXt0JtWbsaAgxSSxaDxrXjDKA7mCA9Dyi
HwMYSyV2M/hrqN8+e7H0AeNmBQuLpWFtn8p+g+jAY2KxqChfeY9E3I0HrnijHIAc
Soc4l3+maz8+N4+Gs2tlP2t7pGB3EDE1Zv2thIgkFh3Ea8lXpHGH2GiB7w4KG1C8
DWySC57NRKAnp0/HcGH/rWXH3CV7wOLsh/RWCI0B+98nqVARUBP+wTxf8ULiG430
HPFr1KIZn1T8ZjsTKgL4lpCqAb8uKdz1iiQE4331Vd4zv1CCcJRE1H29leCZd8dl
bXYkhK9QoUCFJl9LZX5YYp6DpRp0lGKJNqGEcqKatm4CPO9dItJqPHgmZCbUt72I
aSQTaNU+EiJYleJBcU8Ht0Qm0HDexdsYmcRGWxzIA+8W/CPYjM96yVXmZ8W2Vaya
1cChfQkd9fw2TTZJK5kP1UkVCF8kUACQPJcS2O7P7csk/XB55+8Rq0XqdpL+qzhz
8aDt+tgf/rF4bqSN4fPRCa0WV4c3e9yjFV8vnObHC6ZCFlpeI+X1F+hz3C2yFu+x
qBz2H5cOvFYLm0iXzCmk67xrWBnu23jtLLocFIgi9y1zKZCu9v2DCGuK4eM4ABtj
FooJHXvKWN4Vu3oRXVQCe7Ha51buyucOCDCa0lDnhaUcvnoGtlAo3kOEjEUilGlI
/MMk7fVU1pS/GR4HRv35VboZalvyL49/f2M58oQ77V9qMRj3jDSLp5YKKDAZs6AW
PfxWp9WDTJ5jtAahDykjTqndzrM1X0FjfTOMJQvS+p4mxEGRx/5XkqenqYmw7DuK
jwECfL5eqdWsAMOOOrlFz12g7PR6/kuTBJRoeNTQZYkUBCJLymtzA46l5LfGNrch
wpzvdu/oK2ajDquQFDSLims/4Mf6/Ng9U5pSzMyBcwpSrCBb4kvitt6M1ojLCTpN
MB1wyxWYV6JhyopnPqeKpCNxWhBJ1UQLOfb0TR3jelZw0Hq3bFbUs+VSN7qEa2qE
zqoxXVoUbNhN8/8ocPAwocO4ohi1v4a59za33jujm3LdU65nPIQMbIOa4dmQWs80
HtYyUPzlmFvC3NwobEBx0MheeAZGOvvDH26SsWTFPvZ3r8m43IFM7+VL+ftIzFjn
uU9R7PWCqFDkgLKDCUP8X0W4Tr/2CcNcqwlsnFSkCwagArixmcViKE5lur/D0tgW
RAk0fIRN1XD3wsPfV/dtKZWSLI9b7NEeQJ+hm0ylnLCLNu20X5yDashQmOd+d4yO
+PzagOknllygHSZ/XUL+Je5MZkQzF566hcpEu1ihHCqNlOov0LlOJEtkjfmL6rSR
isiHkVg+RlhsDgb3wV9LaYhT1e19hT9wNhTFgIMVdYVeL0rzeSZyR8g8++ORgQ0h
jEDOQ6qgTY9vVRgbna9rQOJQdfu1TCj2MFjsbI/kdVwlEXSLPbchHFiuEw05N91I
NF+wkwA+RfdtAJYTsucig8G0g19AhahieGdcDV2pMW7L1IqkBs8EO30VNNbwIJpa
Rl+wYo7q4YsIoIllkCJxEsk4Ny6bOtnlCOo9RyIgQh29puBV1NgvUYvr8ioZKqxa
fsHLAx+O1E/FIaKKZYj3xPvvlojgXXhdHd0adRT2yTJkX/JVYnead4R7KdDZ9te0
CvNLvXQG+r/0RrnPZtzAqc+Xfhv9v4Z/gQPhFUxdbXVYHwlnJaANB2r4bevXh+vH
Ot58IgHIqKgRMxDRNW37rV0G6FtCAsJkXDDXjq2j2aAVWGGA0KKwz/ot0HYvyLtA
K05C9Z7QyzHF5QasNDUU8UCZGN6Pf3xiLpiaHphhA9VeOMvL+QVJvw4/sm3qYciS
8FguEyL6Scsvc4qEF909hc7Jn8ymIj04FKFHPatWk8j3FSG0Z+/gvwY/DeC6C1of
iMBebFK8RzrZJTfgMLxCj7G/z0dSpddbZGgW1xhrPwOo9cmu1wUczuEl6tb0lBBI
RNaXhHA/WLsjXi5h3HT1JEVI6uhM/9XR349HX2/EpxlU4JeS6GwU7R93dIXq91cD
7xNqVGkwJqJsg6nReKVcp7FJL8Stfv2Wd2DR0dgTmuFGMcoJjCJhK+DFwy4XT/5K
QdAtV+OpeMrzKKk8BQK4ds1PY92zlsbqgeaw5gM56JcyfUp98hSJvU7oh1Xu6BZ0
BFXWxmm009fQmOohpGqKI5JeUCBViGAJlBUmQRM7dIVjVwsZvnO0Z/tFfsaFK1ON
W0S+C/qWJ6TgaH1bIi79UbsQ+XYnSk4vLqc35+2nHaROztRuc5TXH+wg0Q9hjGZ4
dQMs2bMRp8rbykhllx6/bGXYURzwBU1Z38rAsjeF1vSn5736sexW3MPTtKUE8Su2
G9l7qaaEOCI1+uCT1ihNZkhqsi56F3StLjhjMr2WXbEtK7PSs0+Kx65nGmpbrAtK
DG+zYYqSdohPOJPAfSW5lfqH04YwjNwrKahpSEoXVEytFv1jmMvreng24iTqt6qM
Mu65yTDDKERBTwPh6cbPuPUYwFJ9GCtFrC8mh82bxqJZAn4vRUlguR9US3ZnPDaV
RzdkjTl6+gwF5dgcSwIyF1ZHGKNgn0qPfIqEegEXRMOHYINEBd6JDSIs4yeOVyzZ
Mu6hPaAtDo3RqzKsplRLV6QcbvoSTVe2UAvnsrFRTnzZRj3OuFWI3E6/hgAoUjRL
jDWlIwPHt4c4ijz/qaXwJ3lKxQP7Z7lMz8A+s71xT/eP0ITvt25Mcr1n8QBT+Ori
RQYjBvERFRudj4WEsK67GLg0A5r1CkGzX10b57e8dQj1ORoI8J9zp68nVpyHbvFT
CHRhoXBn9Fiua6PjeRHS42TbLLQc5PLkT2E3sUVA+6JNoRABbtjKpOwY59b5H5ZG
V2fWafZicGfOezGL52+r4tvqbo8soYT+B+CTbWwHjaePX36rw3wwU/nsRpq9RF6l
mP42xwlYjq8kZ3IT00QVYOEyV0oIQYxp7GwunjFkyynX0XEAZItoCbEnZkEl0XJP
EobKGK18Ij0wnDa5we9iaxQUr5SZGZ+Hrr4SdBu91PSyQXX6QdM+qbKaDNU+V2D1
d1/Lp7oW7pp+YtMpZInHfZmRDKSTFRwSNIyIA+RtZZ2SN/rc6eUDsJwts135T2TL
OWhVhBjf7JJ60SiC/t9VN94ZhXByYRCxTpeINXCjP5RixM+59ioau5Dh+ZWy25Jy
JTbyA+YOzpge3wqP+vhESG2wWsU2JDfXoYYAFUI3H0hRlokevhT6K3zvgfDWreej
PQS9PPkKxxXZiMTSoNuZjsgx/ug0DNzk4evgp3C7DcbY0OgpC9F7lqsGSvhv5vn4
TkcWsuWocJsA9258Eyqub5Q3RR6iFxM+e4h/COlniY1Kqk0P7yIQx11Y+XOh/aUh
ltWHDgcHQMhMpxmX+OYaZumyNgkxO0MCySqaHtHLUiuu4X1KEAS3pNyxJ0BrTpiB
JUQP5xW1Exz0/L8y5KERu1Q12jbFhhCvEdcZnK5czZg8LFDSzXwS4Eph/gFSIvLU
QI88+795eTxJhBv28K2lk6CpAYdj6qULZ6cBlokpw4FPZJfk2ENGWh1xkFpeuc1J
PZ8X0RdG/NCjgeqwibfjIuSx6DNPAfwUuA0QoGhQiqWzsVf7owQh7lVBRAP5gYaR
30V7ulwYwan1+gjvufFwBnksnWwSR6RhPxAOq8vOuRcK43LIcdnD7nfw5KbiBH5W
sGppd/DxvqJ8WVrcuD8xloMmK5XZte1pHfIhdnndp1IxpsShIrtpISFshJK72wER
Ycb93aqFtyzqZKjSEAyJE8WD5dqKIyUrz/TtXf44VEq4knjdeAr171u/esXszfzE
XsEY3QV5Vhy8XYFbE1XjKYd3R73MDBbML7BiOvHWj5QwJCVx8mW52DDHrc5Pnrgk
Y1RnNDpPk99R33810rcJ6Lrcbqolh+lGJAr9pqdFpKPcFmOFLA8MIHnMpkM+RXJK
5QerfqK9NWWHQmYv9jaZirKjFZpFpQ2q1cqHjqE4I1tDRh9zkaAk94R/jryI0BGe
E3uJ3nSx/J2WezgxMXCMRz3MauLtD5Z4rj8gSV0aBXHQd8OXVmim/PnjoshGRkFZ
vy0clvRcpSlychEsBm6Jizk6tZwQplvb1HLb1xtMHJXIYax3YRuN4eny5mOcoYzF
NKEZVF+85pGY7vLLKZ3esZzPktkLv7f6g0fs2s7MHh9nObdtuJScYCMmmbQECnOI
EUGJZBREOB2tT7HmfbUwI5qFLFRyyrVbZgrwYN4e4PxJo1xCL88kl8q6nmuwYHdy
ZhgUv3eYZcSRYbHBJSACS+SUkAPg71okYYyg9CNIaVvjYUt++yo9IscFbXeuvaPB
XXut4DACGAidmUa7EbPm1i4MvRA102JECjy4v+vYCq8bjnZ6Hak654yqT+C7F83f
1wGNSIBGzySvlResrXKRA8J1tzvNU+nh0+zqSmzcqcGT2JkOcwhEs9vLUi7cp3UG
jBJHk4eEBwHKd091CQSXwXnzAol30MMBAfxyVy6jTZNJ8sif+sMsBg3d2DzEkiLG
kQMYl6Kpxt0GPoUJCF51XiuprcDWDCPz5i48oW5QZOm79vV5zpCRviFY4qmIK7mW
wJjyorai9T4ZLN39XZmn6Gqz/b5FLFxjS1jtIi1ZFidfhCNfhYn3ihs0oLQzT5f+
f5TFyNCl5nu3I86BqY0DF7K283ClK64OMaCsSRB95diIUXt7lUut6izu87fyMuyK
93M8jxdHFSVvNl+KsnNHRcdlHXyT3bC7Kh+lpEqP2NnnpH9eWYo2yJTnW7HabZL/
eGXxHK+OCduPVm2DRW+/J3sCgcjwkGxFPYlgTkz3fWYUtVFXq8eEtKgKaTd77R+C
bywm3oEpxBpCgYnO33fYOC098SlXSPCBakCrx48N0eB1Vc9mVnOg2RoJHKphlYYo
UN5Ny+Ry0t5NbW3KN7Q+cMZujZJ/qLZuja5lQ+1Wis9zdE24aGSFleA7plco77k4
rTR/ETdeJJEFbWreV4lOz7FmQ8hCLyWUpqkvTQCzHgoaOukcl0VrBcQX0Kc1790P
EPR4on0B4DPcGsjlSrriItwIHiW7vn6r+oQdKeg7iZG8AbhWyTMnfVjXhH94zilU
T/jszhFYBzxpoXL5kDREj5qSZPlW3aPzBbmmL+ku8PG8/fi9NcVmPiiFb57M2igL
bBCGQVSRQg//qexlCiudDJhrtahriTNeuzVsUkcmflQUu7yNGdtd9NMIKQdco1dj
AKu5FxNHSjllhc00WeTdjXIL3FU6LW7JuXdx2YNL5LAipVcwXZb+hoeB5As3FUOY
27f6Phn0Keq8jdeurjUKl60vbf2cSTu8pqqz1tqHNUXMjLZ0MV4Hl6wVF2xPt0Nh
YBWnB/Hy3bBOFPuh2Zlz8PAe28tVVIuAa6F27RZNGfLOF7B3Zuf8c81wJ6Kudo/D
OK9SrNx677IOQ3BKQt3DhfA2Zef/C5V7WGt4bQKBm5uZjm1h+E9rn7lVqgIRp9Nw
07YzKmPZmw5Hn/fWj41eJmiT3WjNyCOJm0YDo6Mjf1/UczCDiTg2GDWaGFvu+/kn
6V9l6/d/OJytZAPORcTTZH+x8a7WFrekAReiQZYJ8f8vO8tO//2RKdBfS8ky4D91
YCrqzkjKMYkcOqV14i1hqKATiy7XfnyVdMszSuTQzLpM/h+HCzB58pE/GOSMb5FF
xN2Rn73XK9HnHSSO1OSEJtGfvYl8RaRlnXXxsV7hGTEYqxIPAlrH3UhUaaIf67En
nUF3swgnS3EdMhb8DI17pzWx6Ae8W2/PF1F5+KkDSuKenoJe0SBj48OMY5u2sYcw
YsdyEaOR80RZrVBPATRf3sOQqrpy46VWBbNYx2wZvoRP3R10BlWbx2rT+iC1/M9A
UMghi5B1cEHUdhx2Xt0GVsgUoWetFIhoNuNoXZAnHmaRVOK1cKfFfK3K2fjPpWrp
p4UrLUlCZG/IeSFsLGR9MhG1/B9f/s2uYJJrldOZEXnG9kjlCIXG585uRCKkimOM
PTKSn69l54JiZFBW7tAdsfqWU9UXY0H5DJH5XDZ4Zc9spXPkdEhP11g1Zce4jhYs
4B0DSvMAXgHL4FsFnEZ85WzhwMldqT2SYXwiWrDxtRd0PiVuZNAJAuxqwvJAkbY4
lhL/beIbC6ILQMpLGdvbmXqNatR7KfbD4LADYDPdYjTFYFFi5702do6pYkKB7Gx6
Ofe4bZwQZlBNLn+UHffgPAs5rzowogWsLcIBpkkhA0sDdveN2bLA/yj8c7ou6Xww
oBZHz+DHWMF8mrhKdURK3vVD9qi3St6d7azCFrHMz2FlLyLU5OLqtMJKsr3fT26D
l/OLxU5Aj6hCVd/GodR+emuH5jZeHwv7NV49sQCuwSalvDR0ZOXU3rw/YTayfp+v
uOjgooahbD8j8KyeXHxwLuddR9n2Wu8yqy6TRDCLnUxmcVrmWlM306B09VYY4cLp
Yw/7CDWrB46kzlK8KlISeBu+ZcjBh1e7KphpWmHscrkT8ldluQHhJeyviH3s2iP9
lKlcmY5JOD9BpUIab5tDsUP8Cg18kPRa4o4GY5nLtXw2WqwRUCT4W1WWE5i6+BWi
iil5el+gmi+l3Pr+eJNvHTcKvCxZV4eG0jRwqOH7w5LX1JztiCSrT/sF0bEsI0ie
j1P1wr2DONyo3/2qWr1+QVE6L5+fkrAJ2x5w6rWuqZgRe6maDPU4H7UHmmJavOxy
aH+ZnP2KeertzGMjPIeHHISFMx6TGR6KkWH/+ebtJGDPhYwAyd5RTRBTC5JLazPR
VpKTou0RXIJ7g9iWMJ+yHBi9Wuuez1tGW8PuDCuwP9kcUF9v2pHCNzWf1eAO/ll3
YzKys/wXStZEP3Yr2/HYhKlNt4Lp0VnQgtag0XKfYuwMnxfh9ejPMqBPGY56vd7p
MFAKBEElyt8/9C+RLyA2zSwHQ0TqdOTzQiCZgL9ASm3dYMONSvjzqO8zpWTQB4gO
CtQznHNSGI0E2Yuw5f8IK47hSMe1/TryDaA+Bgv1JJa2BQQMQe79CX6opx8xKcGE
TCKH+B+QqGM70/a+BKveRUMGQFpGdDUKXew8kQLjjkbE/KWwV7jBnfoY0192Zxw2
moEIwiY530G/SS1bxrgoz3o7bQPeU3o0qyJRjG8r35qNvdZDu5/Qq+OSekxlL5sL
8PuELLVnbPu+oT8jneNEQeYT1lvczPGotBWk1jQggsfZFmSiDg/fEioP5Xo14fR3
J1Lz6TgCPsKcG9vSKL1hRIA6YqXTl9ImuepQkAd/svYuI9rhoGoLavHntJilaE9U
FFs6zDRGBTqVyvFoZBYTES+gEljMLT2AALe295ugSAE4l3iJGw9WR0jbYjAHKk1R
OOmfzU204ozrADunyV74wWvd0YbQHUq8Pw37ol/nlpzA3LuVSOVpCJSPPJNQp27b
TZRr68SVOWsAZwwuCvRjswV0hsJYYZvJ2avufeYdE7ssghnRSh8lULt0R7nr9Cja
D8pTePQIQn4OOMplMyi/YXIMTznP6zOzoTusUgSgXeAQj83yawFvCSg1sT1FhAfj
HXMc6I5TZh54Ifov8PAKdw/lCRp7cixWaVEAIiZ+Mvz1BtUgoBr9kRJzRR5Z0YdB
Zp/2b/gGvqsZNPeHQDKY85EYCOSAll6V/gbNv4l9k00rguzrF3zmWeVPtueqMHTP
96tfTSiTYPtVkfESBAZk4dt5P0ZFEe2a86AgEyEDmDGOvst6SkKiqoswrFB0KzCn
BICvWQpg3L/7CLZLbGet/VOQLzHLRogJSWbrjHo+ZLF2o5yiOX6OVUKo1NgdPdAz
wbUwjcyOrFEwCXjgLAGmoW1lSNcuUJ9TYuvaKHldZnglT6P4/kV5o6uYrobFGfI8
CCJJ89+Q3rDG//o7HEfTcYFokUlzcaSYCwY4gzwiOWfd09Y4hi1F166P59SvUjY0
RzHqbhujR7kDD2BXFGI74WSDFkEhrcZ78ob2YOAttfNeLERnRPhG5gSFprL/RNDn
CDs5KJffsa/fgMraEAD9RdbKA3mj8Dja4pU+CMH+FXjU6zpdTDVu4nlat4S7PxNw
6MiX0mod613Me/svuc5XX2aQFAX0YBbeHXf03OiYO/wxiSdGqAxB5j1hx5+yM/2w
qJ4OqxJ5GNhJWZYOrSp6pm+OZzDMmSsd1rV7YNyMoMcZ0/07IXwPAWBOhncoFqYd
NC8x0okpqliLfdZEtvi6BcgWoiRVHHxmI+Y6CK2FsJu7YWSlyg2C6i+V2bWDiYav
MONheVYDQQzGW6rROseIQDFB2VXzIM8qqAXg5TOEchqn4qRAtN/mBu+7132YLWaH
ioxBCVd59zjGQdkPBD41GF2pgamfV1SpfXZnG24dVZy9wWTceT8XvJ4mZOLXTKL5
F8gR5njp9HY9izyJ6Tgpo/+wDDMkMoSM0Qm2tENEs/yaL5Fut0mbDV9cKX7fBppT
CkY1KZlFfNNEVvvv8I0HY1OIPS7+FdoCd9nrYNhW0bsZw9DcJL6cFmJ4/y4rtONe
jeMXQ1omMqEBwR8u/VjnGz8vcekiNCgxyWxrWDs4l6GcbOQeqhy6lf9TGalKjxqN
8aE2SqGoV/Y8yQePooP5bsa7pcQ/iR8YXA2x0ok3q2hie2SQR/e3YPCYlC6fBj4c
3xeGYaheIHhGi0W5lOhbUJXXkW1u6Qw+XGAuJIPOdf0D1w7OethSsUrd3uLHdiTP
KLiSNGD/zAgGwiLRNCT1qCcnescKNOCF+8813jQhRGisZoHpiIcwr8O4VzWDzfN/
plHlmrsOAVLD458hzm3NigxYhNr5AJy2tCBjzKUHF1lEEqxQuYM7u70GkbZfkhs9
rIMUObGlD/xoEo/Mkmion2oN3g+zABRyQGnNC/rdAKEiTEQZNmEfDLZI7YIuk+aN
ZABCgeaGcNl5MtWnnoTDzdqaNSnmEWrcTL7kzLMPOSMuLvholNbAH7DIvjqnAQV1
2DEf3kypj3IRbd64OtPUbuldz8ZpA6A1DIEQf70qM1j8x+u+I1YSd1fwSoC4fTr8
F5jHT9XRe9F1h8K+GAhTyuTpfgOb6KAVnj4hiiTsVZnteO4uNZau7g2aZQP/LzHB
mxTOXGxPMhltD4WvdWZUHS69s2h7MNGmqxAnWqZC716qOxfNjiElErC43ZfK9cs5
76y+NqoVC+3Nl01BBlwoANfoXB1DlSIUzd1VoT2QgFalcoUz9TAsfo5sZ8G03Jav
///wEl+Rt25iRl+zQDEL06TaA6ly+GkGyCpNH05H1mHxgNmn5wxICOb7aayK26Hl
bpXGMnDs0Zsi6lC5Jmdc3lzsh3NxrJuh+zIEvIgHnXal5VqT9NjkBgbEjrWkDklD
ZJ+PcPaLeeluYW7wEZrTR7w2NHBjSccjhFdh13ajfAwG+YGzlFyUWDLev2N8Iwzf
pwrxX1VgTEGpAtUpM9NWq7kHcwgLSrDYlVjbNbFL4tAwlHsnwnyHm+VNaSc1Kczh
ChEaMj2d6iwtFX+mqk/3iJPaXpUFus2/Vjk9d5yv9J/v6V7TQ8IZgMGwPIaMvUv7
pcBK+24OMllVWVFZO7zyQajYV2+TjA+WwQTjy4Gfx84UGLaOYK30iQcuT3agKxGx
0c3E5Go3ThBPrxERlBNJwAzhG2DH4SrOGPndNaTz8n/uCgj9znsKAMYHkQLB4Y4h
kpcHfbty83aKC7uAsSjqRfsjJxVjzf6FBQ0fysjC/UPhAR2c7UtDasKQy89voKC8
lpmyMtjgaWq/CkARPK7YJif8ZXGSTKj5JslfNdMvjmQsKep5qPIYQoeGLfTikEQs
tVWs1q6YeuslwcJMGKTi6+V+4J97oTkCTk77Pk2tA4SCtX/4JLwiyPwimRAUOjpq
KXu+tsAl6+4H5OUFuFtkd1KLbPxmChNk/VaEtGfQQyCOcfleKyWKSSZ3N9zemvc9
7naGiWL6UWV3Ei0WZtJd5+zmAtRbekcT5xVRe+trAaUewVpJm4nCbtG2geACRdMs
gMWI4Mj11QZUKqHWL2rnAbnA4vFjzDKT0n+/IGBRSYMKasQSM/xsi1Ln47axSMDy
BkEubzC0usL3P+B1h7mfHBuKCfSBUiHm2uWUWV3suMmP9bHzjoBi3AzVzYW6KDqw
8r7j0fertgp1T7+9A3/+YzYjy1mUV8ALJ4Fh/60mF22D73rNdMuvqhn+PmDPXmrO
yHB7Jt5w1zyzfBbThbhFc4HIJlSKOSeO+C/iO1JiTOf+YGVP+LJxji4VRqGiTjUs
WSAzoI4QFO33HgQ99Fhe389W9cc87qaFyfHshmiRm4evEnjoDYEuOYczmB2fEhnR
lWqrSGdMsRYeZ1NB15IEivSPJPXVyxZhtKcqITYVgpWF7ZbYHyTux9Mm2fpJ1bNu
hdHpBflDz9b3Qh2TVG4RU7UtcWlvnWBpSrL3mcBXLQztl8SVrlTHwmBOUcHfERTM
gt5bel1vUPKjRBiQ0CJKQr4MKJOVoW1WM9tRoByDcxYRM5cs1CmE5xi06DIfiSHq
d5mSZ6xlmcN11HJq2zxV/3atBFUv5sokK6n2R1qpKDcvJxuw7aJKoO5Cx26WLViP
Q3PvlEAJy772Gv9ca8MdJn05yGjmiP2n6hlLkMozZml2NekWPhhLyFIbH4mKtjz7
rhME4Uy4tPSIw+26J36xrk4Y+Un4zOvqo4rm6OiF2vvDg4kF49pwKyP/EjaPcwib
dhZBPGs4VV6vdWSnsT0xCPy9Ujh/DYGCSFSI6zZxAYIPGS6ErxYmTZecsU5U/oty
ZfynmLHgIqBeMU4tR6vRz77kWbMgprfA5yWujY9t7oo3P5j3BbzcGfLOrN1bGF/2
7havzVZAKlYzyiL3PwGkOR9G7jhfmYdtd+zqOtslA1jQzY5xulAZrKqUhi9BY0Oz
E7aMPVeHPH7l87kA1GYTct5ypneUoCFZCzxmHettlZ+yM4Hvv+hSvcVZ8PxlTtpk
Dhjz4RwuoEnkKlUwplZN5OOqqlZv3w4R0WSNXYTi0M0vYk9aeMD4nEsCRsjBi5mO
/u0vL4x/k1c6AtGAzE+7xtJ/QrNww/csAzVw6Wut5gWrEPrHcI5iCGxY3BMF2nKf
Usa7ZWv8/AmS4SEU6IGBFxasw9oVW92i3ZNdr198M4+QF1XF/mnP4VTBqjih/QIx
YTsCztsao07y7UfVh3m1qN5bI3VDd8twc5vcaQIG6ZRvOMHBhWZhI7k8UgFJxbnC
klmULhGQeOE+gBHPI/+h/mTvXzbYsshn+dPpXneO0zV4COGlW9TMsf0DBE/WSgEe
f9v6EUvRJVpz64t78lME7HVbvv7yQI2nTlehgmOmezYJnpxAFNAgCeH3JXpBr06B
n2sPZVK/M1Sdb669Q4ynLxGGr+j1u/pJoOdU3fG1/nMpCiqlCUob6xvVtaLvwWRj
hEGouZWpecmd9KWp0SpGEmtWpXwrzx4uX9AY9ZwZt+zLo9eGH7ZnSUX7fDUY24eV
M9735/ZheCkPtJAEd5z3XB7wv//Eay+0o+Mr7t+P84IJYaTCZcvkmdtYGxDSU5as
4CdCs7hA2LaN/H3vn2E6ndrHzN7VWb9ww3408HbU9UnUf2jHVSdVQ+w8qFS+j/Gy
6uC7bb+fXGEu0Q/Y0x9gwZvSKDYIp0iGvnPXcEB+XHcZ/gZfnpsfyoPAGJJdSYd2
f3G26GGvfmjabtMaAuuWzPWuXjKnRXZ/dD1loxQjbKvx0ur/ehyMeDIPJ5ZeuEJ4
KGOFKZSvhDnVghWDBXrqRzgLo3jmlJAs5/QeLaw+v9cCmjUO0VeWcky9xs1tlmRe
wQSXwSIe2QB9AqiPGbMKfb46Gl5HpfbHu+jUEtZjYvl9gJbqnGOzmHpoLwaehnz0
IlVMczVvvNUdbiwmV75Du9hMytb8Ro5eUE+BdNzhA2zdMyRpNjzMFEBVey1nKW6W
XnCA8MEjOSOxQCncgyYdnU2Py60Ym0dQGdkAugOoC0cfdU/JOpJcRwPVVzYtUPwC
LyXFHaW7KXXzTs0Tku7F+ZZApZwqsWQA1o1WLn+g4H6jz+F8FPVzzJH7Sg8DZMdg
A/Qf1Yxrvvdm9hR/GPazJSomFRf+2lfsPvp600ANFHY/4SH63Gm7tM7jL/q1WDkx
pK2sQ/ehO4Zk+YeUkXfVU9vfwwrHWlYMck/hODrRyIZyyS5tygT/5pirPn6A61Li
3skI00nF3UYJsICxefKgXiUgSaKIyiP0TrvOo89DivI1MFFHsxKH1QLy4fH8niDg
5jKHDRRMb3kxGFUCkd9SAW5v1UmfMSNGctzfCGk61k1QTH6O8kVkNKaHsB2FhojJ
QLzGoBh5gva7/Yijo8HRuCffBmcYWdup0/MrukKzYiDKlDO+qIOuL93WrTq/o9b5
oMPCCL2hBA7dOaXGu24xGs502IHof7gEfX4UYzzgYAvmQ0KFi/11Dtv92FE6IYOl
94JiYRywX/JAlHqZ+aoyqh4HzVdofqQAllX5DLcczw+3fGbUfRz/k/nUzKM6pYl7
Ca8+irnZYHRC7EDBsColf1UgbmvUIko/gV8TmZCZgLL+8UpfAci9GgcKRaWRhON6
lqfgUYS6QvyNTovs2qnVyqsJ+eVAACp+q7Jf+VwgH/4q+OFUtUonhPDjVpf72/6Z
69uUsguWbrRKbAnAPtcpcYow3pyfRbwblBMIr08sGdhBx9RJqNgZF0I3vjhUnQnz
PMUgW3pSXfzNXj2phnpO7qDHbqvZZj8xqvU9JVIRbwF/GllA4iVil2aMgFdyowl9
sO6kIwRA6ZdKY4hOsHdI/RLFSKERXkr8fs0QaAKDe30V3Vv4L6Wxt5ANCeOItguE
jDWDfpVRjhan4JfMtuvqZlCQt+8AdTVGQ9X7bv84P7sqZb4Mr954bvhDIO7SQufU
KdcIIX/2fYDWMdCrEk++pyW6DItFfGpKd5OZxCJjzDWAKUK+4TvWkLF/LV9CERmM
X74ipZjCCe8SKkl6NtSX6CC8/ZIyGuwpgY4dxx8nkxRJL1SbcAP5IDbZMaaSN94T
puhGA0Yb5lviHsVN+z5tBVjFz135+wZoohHGd9T7FrKfGhRBvJK20A8jvz15qRBG
ErHzlk5cFA0+4a3o7YL3lCE1PFHOTl6TkyhM25AlQyDfNKJWr+8P4R/2Ern3YzdB
YTigJ0AslM6rYUBc6ouWHM2ZxfeptJRqqCjz2WaEKtOcbx/nJt19nBgFk1Gy9MPD
PbhoDvzGssYqsBgIc1sxkR930+54qNgi0WBToVPZ+fQBUTWmk1e1qQ1IcrXplMCv
ItnZIrb35Vl9PnBQShe2yXdR2q3sBzvJA/wefBVX7ZMUFfY6oucSnp4bprcofRam
w9oIfIKDYrW1BrO4WEbRHiUkz+I0MzHICl2E34aeQVHwDSmFq//TSgOCYZ3aq1uO
KLIeuYIUqX4qxHuNSa0k2nkgb81xbDRgq/suf5ob8zN0UxNgZRtjROFXxJwtFOVz
/SVcbqPzCJhdqbAQwyDEKAVa6skNriqNtcqWXqjCNXWs1IyXdEcw3ZM+QMx6YgN7
pEwqAX4Wqa8e8YK2UPSPs/4iLA5X4fpEPw16+7j28oBDfvSfjJ9SZ4VudlCOTYp6
prugp24E303rUHwvbNs/IvDUf4tzb8TR9Gmu3Ht3El8Q++3Q7LcFwSK1IFj1kgyf
jMKQ6UoXH+zNwt5c6fUbjZjped14DaLpKZahlXvYYtuGZrxr4Atw2k0OAGOT6m0G
7CuxtC2rBdf8nKyyKLEKRPpZlyDY5H59n8nAyonJ0n940m8V4txXv+MYiY1DucGV
XqdOfWgSsfL6zdDvyxOyCTlM/Fk2fUkfpp0OiEZDH6WsyGkw8ijs2y7Khvxb7GtO
P9lzpWlUXXYPIINMo0oBbKH5HxSvbnfWsVdLpchL64Mc/yhDQq/SHXxgYlh9T32z
SJ79Vo828XH6EuoovbpF3bTAuSnzGx5NKP+yQcrCDQk8CPb9dK8rsIkKr8Zi2MGM
J44oYmqhhLi0FrtntPhioDw4rOpbTrCB+hRZTpF21MieHn8izPfHzuGj3tVofWqE
BkpiTXzouSX1WpSD7WScG7GXfLAHbloK/QF5+D2REfXfxYKeIOLPjaPuwDczUQvL
D38QWPKdSXY68QG27VTWnL6kil97P9wmk5NPTPNKH3npxtT+JZn+FGVxT9icUeJw
qy5TCwTVVK2BxmoMgnDLbl9SBAxO+Fuw/Ct1Dw5RvKxxQQYUObGPa7h4AsVjhMHW
MkWzSZVAqfzr4ayiFeDuIbbHSBGHyVROm6D42pIiA95wUOt6mS22CAzYxGIT3ttx
37KQYiOVON3lbl33/Yqhw+M84YIC3Dg9OegTkyV/fi9TLXoYlFSTOj1LLzKoPXHc
WGEXvpH8LESHO06XTCzihIE2JVocn7rUtborOYrcL12jegXmOgGgqyu2K+wmRUss
uU5PCrovu9qiO6k81kOESME9jyI19435vBHcDYEk7KKXIA+xxw1OEcpzVcLoF8hp
sO6gbrCajdfHUqsbEGMLESzGcUw3lSYLWvFJklwb7/hA4e9gYVsYfv5FTyHAk/6w
HQtVeK0yREc3TtOwOz+TQoz3yaQR2oSU5SBdRhF48XnGbMgYmzMKz5RuKSl6ChB8
1g1Q++QoEIgFMIQBrUvGj3+mSceyKyQvSJ0ltxsDyhTZl2odCegSwZWMK6f9iZMs
9Bi6ir8ajQXeUyu96VST4BBmJOD1r4l42mPuAwZMC9lWA6EJxUkwPCsxfWtPZ11p
l4vW0Ij7AAAqOmg9AdCjL0D850zuSJL2Iu5zg2QROeEeiXSMYZmMRW1LpT6b/2zI
47BC8knlFr73eU3NgXXz8KZnEk4DySAiE+b7S6ZtQZXYi8SY4mJtb591JN7696YB
C5XoQv9WNeD3Wsimzhvbu6vXNWlbIZgfZFJVV689yYq3HxU+SHMIqeC6dpnZY4Q9
laLRLe+U0iHKLiuHAczqPAPRQWSijyr//tS+M7eb4cjvsGvC1unDXRVTxWuYwlBS
N+sA1iDPwEikIXEv5F8vdKu3w6lGJyqIx8h4QmxSLaKZvfLei1aHvV0Es5aJU2sx
SDmp6t+9Ai/YXS3rR3kHAvOoWmMm7P9BJBEZ2radHSmhZIfpdIHiI/LW0nlCjq+c
b8KvYxyMwfqK9Z9pZUNutU8NVWXaVbewPYlWQQf5IWG/f8+Ng2N+PKejWfTLB84P
mnmwdl6gEDLwYU0/BCnEurSeJPtYT/CbDgwos2+3gbqZw0ZRxkMEfP82mldQEaI+
C2Yd2WlD9ccCwINmXZfNhL5/QfQ11oj//6cRkRvVY1LHRx4IP8xHGkY+w2jNHGLz
ude0quBPvoy1aJjkuh3hy+qJ3ajowTAjfZUlSZ22anPGUXV0LPn/bjyL13kv4abN
Fh+c8QushjRRr5JsIx8W/2GjJCzKQCHb9NGvGVTmRr9+NVywGB29+RweMlO802BO
twH8WSEt00w5CCwUPQMc+/P918pkwMRQSTzfGAKhLA3itYlsQHXkCYWkO7g9WJI4
BgLsxCCESmmTd8DqjsnQXorxmOxarthsS8DBa9Yz2D50XySL3QCDHvyCaEdQ08GD
A0BE7igQQKeYKBq6+edurPgHrwIb1W2h5wDAKKfB9KsSsImYGVNNNCSkHHtG2afK
qfEAdLajmBpT7UqcsuoVsrnev4ZsHkd7vAjzntUZYlUt8bRno2OGhx9DdUAJxhPG
ROkuO3iWzjn8x/uojoAr6VdKf7sksi9VjGTyiDXS+LC/HJ0EE5A/eVn6wl7mDO/G
AefSpyghLc4yEjQN7CbXfbcaBAQP/qYtVSYgiQjRUfvslaj4cDHHyfYRvt5+f5Ga
Lkr+pT+AEbeJzXNr3EvX9ugyUIcWFwn5ac0uRlr9Y2qxkU/zQV8Yty5yQZ2rO8/5
96YCNhVe+UXaQADLK8lXnATGvJFuGFKwP7LyOj6+HwJgGME9Qj/GG4F+2DWOsuXU
pG1IBjmIUm6TLD6pAatjnTYd65cNx7AXSK996unzrs6z5Bm1682x3ifzFueDOct9
d8pEPoKzJnLwLwWizqr9G7/RZkXGXRSLiIRjm/tMNuRK7avIABABSM9k2iUwbShe
2tH5tmj+iowqmyacseZ4eNGkh/l+XTVaNMURlMNSW/n/W8PouAa0bQNDT7c+4Sm6
jmNBkPM0Zx2DbNByjjMd4kSJLnVLQtuUhStuUEKbKzCVRM2j+9UWNou0f0HmnGSq
BN/og7xBMwanu0YA9xkonLUImUH4lp1tFCFf7BLa2k0EBOilWCWF/PKAD1lQ3Rk+
Xau9xOf3L9jFmF+nCf6u1AGD2Homf3t1mr2ZoZXmWfijbtPd2A1y6lKitWP11kme
mNB/8J1G4aFAtLlkoW7leQNF56yU9MNDrsyBhjomvViTnD010iqi8tPWDtjWMcZA
ranLw6GQX+XqrhxBjtu7QQX5S4WAShfMXE2ASubykOvC5sp3bhb+3YwNBgjScWlX
o8lxXA+KHy/CglwHJCxqGN5pWFCfPWm/kjdqfgi42Pek7gVNkJri47XmMBbc33QT
pxtcLqWUUNWf5+fYM4EeVt0p4LU9oehmUriDxvhRP8PbfczzMPUufbzf+WUz2WGo
m0g8h8J4XormQTGleXMRiwBUygxabD2cJ8kyoDpDL3x16TQtkaZvaupb1ddAw4gB
ySUi2LdiJXJ3XoIequWppryYgezshy1tRvMmf+MPcnMQt4hXD1JBWgi0Kk+t/xcg
n4f7tSYJTpBsS9XklAIlZTXaT+TiQ3Nd03YMy5DDeP1spmGgI1DSnPiE+BPy8BWI
XjHDSOsqxdkJrx5zwyllQsn37Og6j2F7+1LEF8YpSMw9kwdMIuBTDX28kcSHY2Zd
JcxK4fcawxGwKQF6OLjnemS1ttmccY0jYlFpFz5TvKmEzQ1MBLf43ZFE+ns73KI7
C6Bjeyip43frX0bf+aitR/wTN6j+AIaSHQH/3n8i2ajPX7+WPKEzX/SYGz+uJlTZ
HyY+6O9a4pUhbCL2ZwUonnHWJvdwLyMVcBWNlWEnRfQxVewn+sUNWnxs+2h7wdvV
BlGzpaTc3t1U1+Zs0q1Z7w5RyAGdYaqurroWjIJn8sD1fu9rhmm0KHkrxIo7dMw/
O0Txc6cck04KRj+AsdKGinQ1BM8Fca3tXobtGEiuvGqJMnBTq0D2Zkgl5rIVOg8W
ajXedJG4fcKpvWm1Q7YbgWFgK/lW988B4A/33r/X80uxmb82qgpSxIUdXDMcrnIz
6rZixresP3BY3oetjNr0ohIWw388iA/hprcIC7Cj7r6zSGFi3N4be2HOLFYAdqdg
XT+66cVRrIG8X5e2UJIYn8fBBUspYGQ1UyZEwXDhL6+VobAWuapnU4/t2mG8rolb
Z1D9CIqur6vVihpvaSnep12WB7+L5d0kQ93dJBgYYrU1uFjBh8I0oTSVpkU04EbX
zVDlJPoR0S3jz8mMULAB6E7jKGrYF2J7bRzbo4w4zPVsAC62pv7de7fbKTjNin9Q
Y1d94xP/ZeDsP+bA5nC45qOjiWuEOy19Afu9V79LLnH4yLqjLsOpKFyMBsQxh+7L
qs82l4fmsnOAo558l/MWCBBLAhxudgeEGgzYfQVEg9XXKTSdPiT7fxglQsLkMZhc
IKmfEQ3sNTzNMCZ0vWrijSjqPukF7ffszLOJDsXKcHh/tOUzwfMp12ToJZqaWpt0
BqhKCC5yQieDDe290x2/04Oy1m2o83ah/n3cP9O+2qEs0aK5LMyiPu8ycSELbR/U
3/l6Z/8bQVpgA5Fhu0bc3cc8mxRrhP+N48JQnLhkTBxXQybL6VVEWwAIQMd1vrAT
8apjKlfMj5mDSW4riD7ixXdgfpTWpdF3y7wO/ctMSYph3I3ktWTgPw4PN1aWMyl0
DTX528CQE0QCPp9IGg6YUx5pk6LqUTtquq8BfyGtpzyAccQvxwOPIv+fMtj7qkCP
8aXAS7oIFooy8x3x3vUTiScMADf6EeDi3Rrj1tXZhGJeD77jOX9CQRYxzHz4YhjP
pk6tQ+lIwjEGu7ZAVEEAxC3b5GCHQK7acRjhcvZzbyoPEr3B8QK6tSIeFPl83+hF
kU42leEaPCy4rgZ0oF3OgJmzO/1L89CBcAHb7LB3m+9Fur2rJz70BPQYRPn2MosJ
RNQTbRM9lA+/zDC6mexOwgHq9au5xkAnOZ2Xnv79iyYP1bLSdqKQTmgxNZBLboBx
IzJOBQSLWBJKRnL57BJDZSbofyL3CT7lfCfOtI1VukRUT8V79EMiASGHWlZVJRyw
aJYSg+d2UrIYILdL7rVUuqm4ipph66v6dvItIZ0z9fsZEkQUBfAsHvxAYrbRbQSb
iGFCa3us0ENI+stAL1uOnkUZOnH1k/1FcehNSX6vxnPXLNC858SAQ0Y6/8KlARWW
oA+qfPhqYxPL8OMGKfdrT9JzKELrHASlJB5fZO0W7tiTB2pobDUaOMP5RcCbtweQ
H+t12Jbbxub6fly8lRZQBrpEp+A3DGDxOs2UswUMEKTubBnIhsnqLTbcnUoSNaRI
/sYd32GF+3Dgy1zB6zDZnDSK9rzi0vIgjt5yi8pDQHqHy96Vjxv0iJOesnIqEbRX
Dab6wfuu6mVyALDFUexR2S1KF58+pkiGeGWEj0jAOLKi+yL4bzOixQftTjr0g77o
M92HKYxD3b/XQGu+OZrn5dELQ2o5vSeqCkJ2bs17hQBbrIT0qp8olYTDB4mxb75Z
FZD1ot0JY8zxA4ezvkoanBbxcGuhYnlSv3spUUFXk8S39nXeG/kAJ0OfYM/HVhki
SZz3Mu9K6UmLnSHNsFanxGoxgU+hod6B7n2VlG+VOD7dchpJpcDzLEUauKRvjN/t
Mvtv7jE8VqY4FyaePRxILameDJEi6ceNXC2ReGSgslpm274WVRcL8+NrrnTQKzCt
aDUtjJtJWlRBNXU5HoaoZCHr6E6utBRPTFROY0BlDZNX5p1uw3iSmU6EGkmxU6XC
hr/HR4nt8XC6LfNkIb0ha13CnroB8piTl3rPKryqJ+w9cYyMLcE1HqhMdNRKJnEv
9KKv5qeQGnQdJndF+UdzqNF49UD5m9ohLbiMcS3Yr3CkorJ3ZX64amjuVDI9BlHo
UQ4FfaeOOwoPE0zIm3NDYoVnnqOB/mePrW4+L2wkNcwwSgLZWMddvO9/5aI39cNZ
4Wv7WDKpM8ft4eBXr0DtK6JUwXTVlKNNjujRO0Jbg0DNvLylHitPTSP0tgB6HYph
E2vBdHCGPF50+NI60rvxPFActhpWV8M0qIZYk/AWLo57Hu0FOlsCLyumaqcrkesT
Xsw1YHT5tUUdfseDDvQ46bEPYv50hgyDwaLzLaeY8CbgwWKo4antavJjFhG8gd7r
MokKLE9LjQWuJ/9NNrQmZ0gW7XDxNLvvB7v3M8P7eIalPDD9rjT9lK6BeoWoBzro
WNw+szI9iIF/Ru4wtaZrXO2q6YhbXRjbpVWKO7vg2rPuhOeMemakkZ474CRCbZkU
7ThO0bPXWSlePdZM9EOT7QELmoVknROp4TCEi8EK9GhCKKS5/KbKNCd25WgLbHJP
5gnJqYGb0Ve+cSZXoI4vufYq1g4n8OYQNkD9WkcBH9nTlBTR24q31oPbc0nZ5G56
EEUu3hBqbSsIjLL2axYOuNF0NOUC5mRujKKZ7yVAM8ADkweXealzWegVO1ZSiuFa
KqA/HKFpWplnlxNzkj/39TTB1kVZokxRf7OqaGCjGJrhUB5Rg/c2KIOh82Tiyrqw
jA8Nb3vNlIzpRgHrvXa7QD+AfjsHk0W+TKODhWKL+CLyNxjV0H7zrZ/I3Q2xyHtm
7X7dv9tEhWJSlyB7IvQOmgLR6yae25jRR5hXl2uiDJOWHyGybAzZFVJVlvamgL04
pktVdol7/uE/l+1y1BaPPbooeMciSJNrqnQwt2Oq3eOKkOTVPAotW+uqJTYg2kGc
1H2LNw3dfBKtNKCjAJsPOZNSiyE7nYk2KrxrOZHkH+X/R4ADMQ8W9N9D2WyEg9kL
JoHoZpc6ItKxWTsX0RH6Zwgt6qXLHlERyBqoHDtyHtYc0OPIx6WBsLK62iHvab/D
zqOLhtg2OYA8x1isGmMgh+7GLPj520YXA3Og8BGefuCtA99Za1I3vdEQu0NLjuhu
3Pvc8T+ZmLHD4A63VpYI93KwjeXS51x4VqvcXmGkCxtSf0yFbxDFKXZEz6Q0DLaB
r1YuYTgZSkrs+onD1bG00f/c7FTtpbyGGq/vu8TiAIxB997MK0Gp4tn3LmjFna42
YThMSc7SrK8A+0v3yQtH/IO6XaOpufoMEZvmVhmGyNYAU5arCeTxr8h2UGnJ03Aj
DqZfMawxxwlWHWobkpPOTpkMpb4axrRYiFRIo1yEMz8v4y6ejY1ZE/W7qaB1yUeQ
yk52H22iz2qxPIaHZvTNO+H8S0YRT9geUvNL2l3MoNP8VNIQ83UR/1R3Bt68KkYk
GhWyVT/OvtytR40jSn8cSjHh+WXifx1JVrr35uvS0g/hBTbVYtvXfay6ljYBeF5N
xCN6W0m27lvxMegdURKdOX4NdUsmi4GgIBKYFbjr7HMiQTeBSDF8Eo94khHyGZyk
7wnX4BbCHQ66Txa+qYwxLESTw2UpZZ0JuIWWq+9YEaliBGCzZwwmo7LwSR4Oa88W
BBBdRooU7KtBm1Ruug0rXfbbXtL1B8RCoXJ6OcivAB+ggMtxzQ20NEGlAPiv3df7
yXbkrYSWw0iyCWa2nwjzMBXGHk//Z8aYb9t5RYvyoDxxZYR4llu5zxcPbuRNNmlA
LTVJCRkiinrd/d/xGrh5t2DIjlV8n+iCVLasfUBset3BIBL2Ax5gn6x2PhA/tynA
Y3nukjE54sVjTSgkXABDtXp4SlPFSTRnT44WjBW7qbyQ0l0+qHd/DptEeyyjcQ/2
kvT73ip7HDPXjuto2L1/gUO79wnZ0bASzRagnTD0igSCTZK0GBLT7ANFe93r9ckJ
HlszndN820UCuanzD4eChU2aZ1ZKf7FhMKdrqDruKsQkDDRQBFbh/RW5W/7ayDkP
2FzQ9F7rcY0ivItb+HhUiVUzFjKzcsGwzYYUBjTDNXbts8+pir3KI0gmwkXrkf5n
p9UuMQTi7sZKv7s9QAQ8l2VOKTFhl1ZmMKkiidRLH6jBglcRD2+yh0zwRsvWgt3S
ug3yl8MUtdQJrvVGQf3jPtwOd0Q+OnaNpLQvxJVFYQomByeNim5j5CaZUE0o/3rH
PcCoNVPseeXrn3MxNIPYzquJS1OKCllQAjAdq+b2sVCI5H0OvS7vNbmrFr0qt64y
z7GRzGb5eR5gZayUBHmFqTaTWgxicNyTDssCeKOWsYtJGyWde7hiXEjd3tyY5JbS
MghzcyE70sssBPYGkMnystj7Bf8SZXUtluZrNdGcp76WlBYyviiJTGtEt9xJNKIu
2gvZ1/vJ5WCL6jlK6K1/YWxLBVO09Wem9RxXDdipqrjLw0vH3xvg1Dt+DvDsEkP+
k+qAcqDlopozkTStBja1/ne9U9yP2bG2xa5tJQumjQtUDYBzXikEWh/yTcMRI3tr
SBLjpG/HGcDpTo+rJXAIqFnhcn9npcD8uyPrSfuAIPjGn2MYbepsHS+iBOqIGwel
KHr7bHNvbXZtPqxQ0DcbVxtXhnUSpb04971wjB7R2ZfZv5RK5lhpnL03VQYPw3Bc
r5DcpfjwGS3wl6969WT9V+nvZtuTtI2tJF2vXhSzLyYTqgi9KqpyNrBFbcSU+hyg
OL9sRpb4x1+aJomzdtxkIDu6V7fYR59Bcz2xqHj7FkKCsugvq8o3VmQRp7fKYIrz
t5X98AjgYg7SOyzlk16jRRylZ3+A9UZKrvL4y0LRucz/dHr+S4tvIdbCtN8kJ4q5
vhz2/EZGGexajPTEF0EpT9MOCT1yFQ0YygEh8BEg1iPe7tHp2DzqFR958vPBV4iU
ygq0C/mDO4bFJ7mVrVpxGHx4kbdVVioq/iVBuTh47vXzyg6TVem52B6uxWO/WwjE
29Kv1MhS3mFf+iGvNY/uTZdynbG8AstPl11RplIp7VGa/Jaxu0WweaqE399I5pOl
XAm0lwVOFS2IABYnw42GTkItBPu6Q9cFXSJbcJev+9ToOT2KlpYw+XUhLS3gImyA
I+/rBcZYpPfyhvltpQRyTz/snY9niE4rqabL/gwlxE0zh1dW1FDnNRcdldIcpOAr
GzDyYPo+XBLkf17GVaiey/vlLRkXgciN5VetXZBHT42aXK0QqfV/JJHRX+lqxrhz
InOmjg8QT12lMXdy6TwubGtxeAcw507Egd2HHhzf74K/Hoy9t+lZQIZJ8Ol4E5rV
vkfU95xqufXxSArZMY6a3L2RbgDqGT0jYJ2xHnU91Erto2aLHyMFmpxYIM5gFcV0
N4RCF18SnB8IXGlGuPOrXox5OMMaBApDE/P4n0nUl9M7zvI5Eg/iRqmeSwJkGJ9w
lTYM/HfKwO1PPs/AeiUd9TbaSss7SMTUZYiJWbOuXcKVjIpwSrsu/Oc6ucfnXAOh
/9Tw8kxSek68NJb31JXY9FB/eU+6ILbZQZ84VxJW5Umk3i720+0asZDGGJwdTi8P
sDxJ0YvFNK5O+AvOsicM6RLo6WTeqa/qYQpP2DmzwbWvW0i2LQ0ACPuqmF04dBVH
WM6ZYSS1BpP9NDIJrbALIJzYV4Scf+Fn9NzCP48pXeDPM0AGGxL5YeGcr0LuW7uA
ExF8k5TqV1MVVJb+83BMat033YERvv8RtaE+ySpRUmoBgGSPT4EVAvtJ4KWM916E
qqvWrqKdlMTZcHg5hzg2Wf8fbfstMu372a2eHDZm9yRlrBsPi0is0V5CyF7YT5eT
YAbirTqh8yaV9barbTUiU66Y3Agh4T/lj0bpUKcCLJ3NftROGiWvMKRjrZuOGf3k
8Wq7vapefxjKNVewgVR3c9RcMCx2Srekt4O7UVNvVsgobmg9zDCTc7X5GNHv1jKN
cjPjLpIvozgUQxik9PMAkN7HqhdbmfrezD9NMFxrKve6ukB6gDa6zp49GLuwa5m4
iOIYrLe5bySv4Q2r9Z5G89Nt7vNE9aTZHpRABzfWVRYz2CqRe9UvWpzpFwla6Cbq
CjhE/s1cSHPoMzSbAlak8HLb+G7VGbvLcjjCsLlrXtgDDs5R1IkTUJUvcOd/T8xL
3Km0uKs31dQyaxYJxVtRJ5vqQcDhmXXBIIctI9nHD6ZdHxNHuEuId2ThLk5bq83b
KKYv2Hoy1+8T3HouUxcUvzbd3AMowIAuq/JueZEaR0csQNzaeazz8C2QytFX2JsT
/sqgFu1xgwhuLYRAh3QEdAWjVa3ZgEG8HqycFTTp8urgwyttCyhwcuSjrmMrUgB6
M24dq2HdM+jwQZsg0OmHtLKfEA9KOY63MU5Af0YLxm0Oz8iYMIc30Ox3QUddpMZ2
xrCHKAMN3fpjsuHFPVWDlR1vVztld7g/VI+erqD37O88DKYtbDLBrlpXc9egUl5B
60cLf3mC5TB7ROY+HCX6e5GksoLzr9Lzh5i+Ve8TmcGwOyq58+M1CjyGT49HjDxo
Jrf8pphFDFIGZQyprC9n2RnmrjT4Udmpsed+iv0I992ptXliKscaVRMUtJ1Pinty
O12pg2+2Ddi67c+ja/emes27DAKe7QjgMQ3rtnGn6k4rGM7EYj1tEF/K/+xtwi8r
UtJhn7W6i6w6bLmM52fR4C/M++pZn5Bh34AJIdDsVGJi7MYrniN0dZC3/BxeqP3z
rOiHKy66GiFGI//zeEmrtuYHu4oYP15iimm8Wmdf7U4H+jaLT64WhicCcxZAq0jl
xRyE06zyvRuoRCcxkKP9sWq8b5RQjAnB0NgPlkCLUjvJ4XLrpuz0/SVZGz73b70n
AL+RkTHWBf54sTbFG9Vl/xeQcKCONGvi9tOHfsx8zG9avGSO5ptZ8Xy+0tLmEA7a
WZWCev467DjWY+M67a97mroFNQZbd7spoaYeXy3LACte97QAH1KAIRq+4mEO2Kuh
0tTlTuloJ+MoLHdFXtz07ivFaVz0ohgqalNnLog7DZdizGLJUTogI/hacogZlpTD
T+vO/pV2QYq0Fa4G7ICX1ltXU/cMmz3yWkytVYFbvb/2n4hYma0SFz/iiQ4ZOapw
g9Z/eTYZZrE8gLzWN3BXNgR2PdSq7Lgw1VlcwQ6OgkOUrLferDDLY0diiyMFTTEr
o7aGRgJbPD76VcGvviMyUJjXw70e/3rOSjICLDQ5am9EeM6cR7U/VYDiDo5Ox8tZ
dL1nRcv/GejD7RpoqVyDanaUxXa9moAdCMjA/8KjsKB3C/3KoleQY/dQ2pIwL9z3
AB2I37h7CxvhsKMPIDizxI5+E8ck5LQlsVMprCR7cHDRngkTAn8VNM3rxy8gM+e8
lbjZQCtpDfbnwr7jX+j8zRwwRP3jzcHHgpDCK4bjuZ2FEQnLcYNc0YRF1QD3uIXu
bTzQbL8LrCll56/so5ByLFnxQOm6MRnrJloftXxqg6bqqgerf+Z+yLeOJWUGOGC4
Cgqq2rXfEkIH1cp0V2tY/k8mOK763vr39sdrIMF7WLsIENc+u1yWql9Yk9pur/fw
dKPqQeey00iFIagQpEQLmo3kqOeW9wm+zYyQoGmmYV8djA4qJEKRqU+uwkDKwQr3
2Nfla2rV+R7RW4n0hPpxfPZnoQyKHSsWz8CcoYUTxXyBMpQdCmKLCowg0zjtNYFO
0EZgH2kq7sKGIFFC3sXR1EEu/Zd9L2UQ8JEYcI4E3bX3uIAF2U7GhFkeIs+vm6oX
tnWA542JvXwGLGNPI/nIj5mTsOrt92mbhckd06GMS3jzhxuQA68PFtRJRNoWGcpx
uYBVX6oNcoI2BHepEuSr7xphvX/BpWuSHQUq1w3e0/Nnaff0LH4qxh8QXDIJ7nk8
ZK8Ox+PJOkyCRK0Nxt+zjMp2E+OELnr7keuE1Hyf+0jKwKGK39D7aQH+aHJyCwTr
2KTuV5Sg56AZ3Idh7xcDyQED68v6VN4TzH26th8NrJql13jUGxkpbw9qToz+zkv7
QJaNocZ5wDtSuUBs/WUShvtsbPPLVVxKY3HibCM0lAg0E4SSwURZwcofWPo8C2TU
LG6K8LfMFI+Nlfm/h67QRtDowBGxtDCCmHOXZN7BI+sXIc1Sy/JOmdfUFhnHKm+4
DdsqYSN8jwAEVtIeMeuz8ndBATt7n2SmZ81wPbWTthEnLqKVrDSbPW1eC4sCy9MX
dvz3gzu9fAgT4BettDRPVlFoUrUF/d+mLYO+/M5IneLBXRmb6EnaXhhlCSWN/Oj4
rjIuAP0Lsj/CXGBhDNp+AMmPsWHhJBG0+3MgDVbYuaqsu3zJ1iqCrmmcHeGkOfeP
CYgEPMoVn7JVhN+MQq/jdAOJeRCQJCPtWzKlJ5ZfNnjR0op6UBgv8bo/sepah/Fy
qdZoXkeBapl8lVZHJUW14Kq5L0sp91/qA5u4D2WPsyWOrnsSK10NrtPvmM41oUbn
k3HRGjHO3fbHz4AiohY/uuwplKG/Iev1Jb2nnQhwQj1rsqHWRM1UD8hfFgpSp6k5
sQyBQ28dPhQLJmdjNDJoqQALCzFYWpitUjunvn7u2VCDQ4LOiLLAytDwPnsUePJN
AurMK+VMGdgopdwGlNBIsN8ZUoBoz8MRFTB5k1JdlbKx6M45SZAeCxu4xaQsPIzW
amg6sa7ySTxl2iR3d8A8igd2e/3fLMuyfUAw+qvGwSYkbea151QCSE1NxPMNX5ME
BHpmd94XocqMwQmamhHqK7OupXsGW7gVc4O7xoTLoDhuuA8qengdMGfw4WJqSSGP
ywX5Mh7kF5jItKxni592xSg4FBaAM+LxoDn9URo4E35A/VOpmTDERGAzobS8OzJu
W1DHpw4fsDralLk+D/yJ1Mv/VC9Cc4u63U9HYp/WLjLEkWUf0JOQNquCA31RZzaV
cEmMLxa6hAlAB4XBd2AVyXKWSTlOcMffpLyTEpYvprylnhMOA/JAH/VbJG2FkAgW
fhdreqw/GSfgRdzDIwgdYz8CqWogIxc7zV7RW9mLurkprTUGVUsUGi2vQ0WkYP6/
BLSltOP+UoTk/PdlyItLvjzoeXTUIlZCccaLXSbVp3Vb5Iz9yyj+rMZT0/5iNUf6
PyVBWLDi59V4wi9Yt7GIo9b0O8gdkpxZZSkuoRSUSPBBj5i61E76zNHJHbVYGIHQ
1ZoXevGdaxuOb2VgPzOtggVK0Cc1Oi/ejdwsiZ1Y6uG+1LqG5t2GlflKXF+Jc4ET
GYQsbviBmbY8ateYriWf+sqfsAkgGrznX1Jkf7pWgzpeLKvrfUzS0ERh2fCp9Q86
A6P+eCUNQWAOLJgqYJMNHXHFFRN5jTQkWFfbfD97gguFvrNJdUEIbIRp5ry4nVae
KFKc/xh6uw8b1/BT0osPItzRc3GVnvHyl874/jQ4aRh1EQHMT88MKc4R/whhS2dt
avrUQHls6a3Mvgw9oVQ99n0eggAH1C7MdlY+FvfO8xsiHSV1vQqdfTNox18qy5oh
JrQ98OibRW7W45UvB/UjybFvnN8zdH/PnwQP9mFIruGo89mc55crJ6NmO33Q1uoZ
5AI5lyj/JjSkaiTDtEuhP3fmTX2tNvVSOgkUeTiYiSfpL1qFXWTVP963Fvx7DlZN
FFZz7OaTdTukQaZElI52X0MPR2GVkLFesi6kN21tEKRN0/kHcNBspgfABs2aD8oA
QZ9bCB72uuPu+InZfzLweu4r0kiRwTBe1K9vV5DwTxFdI2RkMFPOwVrGibU7JzRZ
7jBDeLFqDFXvYaA1YYvSnMYRRVDhFQXfTtHfuagGZbY9lxipkIEU673ULiRnOvUs
awD8FRTyYINbFNajHlGTL5SWv8iJjli50DnS80u+piKlE0VgNKqYUK8azJI6KUyr
03klH84o5ZAX6p56Mvaitb+lr4YFuIcXcHD6USDTxJV/IKVfLmiHFypY6woEHIda
7oBNspeKGfk1Hjfxmt3BHx8NN145mTbWxWzh8yGpwPFgmOluYgeNiDUpTPVouZnD
5FcsrTFFma7us/2m35avjDAhdt9zx/cPFtk634TYhVSITGEHZ2tT6S1D1QDxC87e
JC8oebncaDAV7vBWgJU9EKYV7pl2WVJcW6Jv5f2fBEQlslNBnJ1P9WV9TqmJ29vA
PAAOvEaEaVxyKSqw+sXnaH4H9iQl69gpXJpJRnZLSrGaIqdXXCkR80QDuKKgFv0r
K8dAb3WC/3eVnSvw9RAYrAZ663Iu1B6b9Vwy2P7Bv3bEhPttQkb0Cezld8G2erwN
EOJ/NdR+DTRgfWgpvbV+N4ZoYXyUko20m5GWQSgp4/JJ9C83QfKB15191VD22aaD
ikG2VjdwIuSiFu+2bIkgWgkkl0FcJTroJfjnrCkDS3nCv+RwMCoyok11VdySJP08
HUHmTD2zElcLCcIz9Jgv/XIUYiAF9vGzAufCGRIU8t2MkldwYG8hgaZkNlqAzAp/
j63J/5h/8FB+axi9KEjrATNwhdEt6EhEa8sD/Kw5EymI7Te/yNEIqgdbzcHfNVMq
vo5puBXi5k4W23lCWW08u8Wi8ONPIsdclVCRDU26tMDjhpBhCslG9YIt67S385gx
NdB42MapidYsKZojWr4Zry/uj0FlqHT1o+cLvNKWMSr/xiwJE4y59f2fmFpvIq7B
8pbwVtqtRMN720ulhX3NYnYJkjIrZMF07Yhknq7UGQrEYTKhpiW3GGzmuIXYDPXb
LRsSYs2rhQuHS0iFGtQHXVD1M26dSPs9Mki4xVHXkLO5kRuGc/SNrXytSJzAmPqO
9PGwhMjRE+Q0PStvjQdvRrjSg2A1T48+oQuknKWyHyEDdHI4bwSBiyTGrzE4HvWs
okCMF18JHBi+5n1alaTfa4PVRC60S3hSJu87lDiCB7JJ325LMQKFNqNL7s4w4VUA
dj9XUwe0Na1UvrFc38KSYDgzcW4s2lyDY7DsnYeYuFZt34vqxtowEJapv7C2Mxql
WPiDoYImVoOnwBdIRYasNjnQd1DueU0WR3fUJqLMwOLysrJUaL3pFRYAaGC5n2zM
3q0YQt2rz0X/ubfp7GGJwTmLbN6/M4YYtvkSiHHVhZtrMvbtM/f60jAdnms+9f/Z
3/3hAAElYrphFsz3xsQjUCGTYttrcDgOgUl5dUmZlXKX4myhwJvwqtlYcm3ypAif
AF8r6+w7P2Z00b7fEN0QBEbhoHjW9bT4rlhQU+7CseUGzT9gQ1ZMcq8L4ztq2SKt
3cPplK33+k1QXdH82/cOZcrVRorxPnv3AzKpE7zQV+ddnBHDWOiifKXq6VwNlBdR
+0rtNFqlkFR2dC82UrMsaT/KC7s7i52U9uhffUGa/W5pXNkpuw8UFt2W8JQ4fwWA
k2JxY969GO+9eMfjpkwYHNekaa9ur/kAXYfwnuwTLRmlAMcvUGlCqZ3TodR7ODWt
InjvZg7DhkBHk4P9MavQZTKHu9++K0UuHjeMgP4xNl8we5suj8JBWl0GZuUrItzf
t1T39qe/0zgWxigXJq5Ow5UzCvc6zm35gQdG2HzBQa27mdNV9PANnk9tIJF5eTf7
pnN8YccnbnfiQRn+3FTjZ5M8KiE0LxsuUReEkx6MWwmQM1HDzWuVmTH6GTV5ae6W
R5+JMp53VPjHH/Z+p4KjBwDonkEcq+FP5oNoV501D3lKFHWl8yh8vCP609Fh2bHC
jlHgA/hwaunSraWFdnLJKFC67B2dGsAx0AtKoJHdqS9fh4vK7L7+QUnjIsjm1Vyt
N7PqaO8nr8NWKPrF9BQ2hse9RGI50nhgWwqhzR24nM7LCyX1x3L3VaR3JlDqmuJX
L8WaJm0p3sRkiNktmjbjTIkkdfhed2aHIgDeZxQwJYUQua2Kf0C9fE1wAJepRtQ6
jQ/S+veULfgjpItSI4tU6qic+eCF6jfi5vQ3Ny1R2mnlGpYkjPQQrdO3deTQ+2Cv
hJYpEcE6Vi+myQN1JHHG/AUWoO64XYDfU0pG2l8v9FkSkFZuTzLvY1IsHHm5QJOh
WZkoLaGAvLzaiSzsG9LjeuvE3FGWgw7BMZfz936yMTjz9XfbewCLOFoe0cbisl4I
BWGhBKwyXJtUTeo22iUnvPDjDOstioYw6v04ePcKeo1Mk6uXxfwcMUWgGhWdGwFt
IvpZloaZB6sEPvmOVBDp9d90D9jIJshzRpubYcnu9zGJbHD2K6qbfAEmPeQ+BONO
Nd7KAx54aoV0evaVqQdY6MBYjkfU2xZVtKtH54ych9mtWmJTSkkjHkRvc/WNAda6
Sd8nNM5l0CJNSO8/2c7AmVZV0BN0f2YO0CWyJHPiJBvuSe9tgHatWXauQMh6aFmu
R/fnjNcTvXoomijX+AyPbuZxVJbDnUhZ9Y86CPN/8KvpkPEPPqoC0cN1tLjfwbTS
BmjE+G6oeO1xKw5j21x/sV+5Pdi/C1rqanS9a5KAqs1O5+Ex4TPWtlhXRO6axCyP
XG89eDogqUJLEy195QqdYIgSCaGDBl+B2Tws8oi7Ch+1vLvVj507YLfJjKSa0+6D
zX/ZK00X52YB8xPRBPK8HrO+8v9o+7Yyp8wrqNJVVewvZhAgsxUWE+ZDWEBFZ9TS
l4el3pOl6/9/lHTYYeMD71Lj8Jgx0G1+vFUwkHKg3HfN43wZ+gUI8jy5mjc3pM4V
US3yC/23nCP5lTE4mQerJlNob0I6W4bfA9UoyC6ReBEo/XV4DBoUaYrFClIY9LJx
+YaTwA1QHbkCR+bi9Kh+IA8k8s0+Qmi79lqE17VCrH4AWYaSJs50fGlYxOTVeP2J
K0yD1w+OrWSTsJGwNs2dIP8E5qedl7ymg73B9TQ9SWaxEFiZCN+XlH00+wtd4MtS
YRmUBRzGbuFE6SRdB62zbijcF40RbQPKyt1GBfbLnKm6WwqRhTDL2k4szy+Z3rRc
xfp0XSPJwaFRredroLRl0rNI3y4TmvDQnK7fSQp2ro0IbhtnPCjpCUx11hPZbtma
X1WGvU1qB5lWWgH2EwKZOenqAjWEWqn4uisarmLzmrSrHI981SRRkEjBhHh5pQGi
bNI0Y2eSoPY6zJeJ5hQiz80KXNTPI8cvadpygCfVR1nLh0heRhGQYKqmUFtL/yMa
HuClXMdP0HS6uWr+x5E0AML6EOBJxooYB5s9pBi/BP6GJvgtXePfHMOIhwhhV36J
Gg41jAOgsY1gO3l47zOv/qXziIjggY1haSb1gCguLcb2CwQIHLic7XSZRdjIYN3f
vNUlkZyxXos2fbmRMQx2fjkNbwpKYWlNI71lbuXe78H3xyQlecpBMD54i3oIs91Y
03ieF+bKesvCm0KILz281KHI44VC/Fb2dqSQ5ZLzemvAJouX0H+i0gtoiH/63X8z
z842/sGaEk0zuo0G7HtIA6kbJq/pmQZviAEY7kXnBIQNuAmjRGJof5CjogddMgkN
ja+h7qrlvft/Jm3WsP2RaRzLELWmZIy5mqzHc9wGdRAo8A0JLZhYmI3AdcC5T1h5
OQVrIyJP47PdbUvOq6vPIRqze97Q4EniPF5LsrfxyvSr7PztevmsKvfPDDYVMsHm
EAIrrgH47H3A6QIS9l0/POC5wQvUJWjwhUhzfDshb7mJB0+Ly3wx9SNqc6dv6x1p
WjIk36Wp0JeIHSschLvn+dH67Rwa8DRue40HrWwgUdVtxTms+7yqy90iBC47gVNQ
BqSDWLtacj+JtspJA0v1sMRaeLv0tmXGeWvOdxRyUg6dXsx22DfJKmzcGvrhU5WT
wMLGLBe7EmZWSKxOFNqo4PLW8GHXAS163ubWXXnCI010vcNbRoBIOTTKJ4W/ju4w
waGNPNzcoiolFQJQVya98tpMleuKWanWtbwUYW5NpBxEUImwCsO21CyNS908lMKL
/wjbDJFhLxeITOAV+xT4gSWwdv8l/PM4ayHGI1WyGyo2Asx9dwqcduuCZ+B49umB
qpfLxKNJN3Fs5vcAOAaMs9gpONTOTzExjAaEu/uife10dctgkap6MrivtEBUyRCm
jDlpDk7wCTAgmOzKg0OBaZtODw6ty29wHGWqsYnoRnRiGcJ8geZ6FV9qeXwsN6MB
6Hx/ZY+TchxLbi64b7qneLd3hk5mjfzgU1N9/FUiaXkmjvoBhLC3IE1xfqYuoRS3
oaTurpUX8tnSPb0UlUlXauL/ttX25YtuUv2/pTHSwEaIVE2qxExjBxNfYmmC96jg
3BfU7podkk3uv+PJ0m1IikfcJRj+UzWwuhD/m3M0QAuFKd7eKUCwhz9oK27ZYK1w
p3UeSp5Fs1aElnNoOZQCHn5G8ZVxDHScyC2DZicpyrdoRQMfSxhKOUBuVQ/QLjS/
OD5ao2v2kiFLmjkMhWHcjC4+vrJf3OCDPYRMz4XImwHZUsJBVQtfYPIRKqA0ytvh
GThZqczvKxTTF5nS6jkJrCgGShART6rLEZSTU4lND2yS/oYs0WnpQ8jOfEK/AyDG
NMh+FNTAko7+kR3BKpZbm511i0uU4ttHuAZrEAlVWf8YRKFiqUhzG/VAYhSwJAqB
13VMEUZ2lecC1mdFO1rfwqrBgTa6waYUb6Yz6rZR5d1M0avyq/sGogNGb4birq3t
zIbF1mtq+Z8SWMiGXjobpmkxhTIdL9DxsoDvMLWGMGpDz4K+NNLgoOtMXv4Lo8qp
0HPhL6THL93kDQX0Dt9tPQOjzBGE+N6QEYSM9GwJaCN4KxnbKSoHgMsnSFSYRQEm
ylWO8nsekdhatj/bHJSVGBIDfK0j2wJjoinrJF2PROQNzyPRGDpFRQeDpttKG7ys
B8RdxioC8xZpfnTnBHoSBNabSX91mLF+yyCGjr0MCo9yC24VxMOqcQZBCGNDb1Nz
iMnqKWQpUSOkkbVKdDRcRv4JWmVdraJVbVHudReSVUrirB5tnoLKTsUpvd1+6+u6
hiqBV1gu1tjKaIcnfDugXv6+d4qo2NFstsP5zh5GrdxjA/xh1CweV/eqLW0kqaMG
h/fhWPO/3BCAE8GTbSUcCCUgP22dzJR0sJHioLJCjCqiPAOeg0MIA5ba7ZRQKWG5
X8POquGkuhpfma3jQM0FXtaHE1+0+DkTObWzO1VjwS/MHQMWzyWbJrVjoEi3yUw0
/ydfRnCitpr94U/wAocCsV5FN7d8KsY8cEPJXHJrRhF0vMo6EzEEFkfA9P3rv4EA
xDT8XepH1ciOS7ePKxm62E1tePoR9yKFhfsz5IihJ9vfzVQkP3h8vkPrKcntEZpv
CFLa+lHZX/0lkzw9cC+TZJWm4yFp7Z7HFznoXan6xku5+gYpO5Wa3lkF4Ku8nMAe
xgkMgRnb2UA6jlAgYL8TI7DAh8iD6pWSYGNMeuCAcCCYoiPSzJcOkm7EC2Yei4Kr
3SaBScRV+m+r+USeI8dptJmnMpTQf9qErq6e3wbTFQHEmqQPxzWlsDebWyW7r1Ip
XSV+CvPhGoChL/BOWYR85aoLYyKwgmhEbZjt08gsWTHsMARVOR+y1cx3PVmQiwob
0qvnYFGYWiauklMoJVZACSHpQG1A2PCCROeecXiB/BqQTtFDw/RhceoQwgBnjhHA
bvResXtKzA0kjWeLwoV5magafywvEanAWI4PbLbOz9D1eDs68NnElOjcjzgoKTgK
EH4TjgUf80v18Tq8LYbQ/dgxwK+8jI/ACNK6ajtrzzEA70QEfvSoJlVnDLBEkciz
KsTNPxSk2WdxUdgRbX1565h9l7h3zCRHEUfwXPg77DPmU9Wx1yNlCWPTQCnVZO5W
3PtpVY6BuhmS1sjhfAloHtNbEN2tGgQGtxOoS9Q8bZEnEaj7fGbpu0GWfPvLXGQK
4/+4Mf3BN359XUS7ORmMaOuang8s6CVpa+el1osbMCSIPATUkJlqZV0p7Q9i7XIa
SH0dX8a/W5RWJQN4LW5uqD9e6tOyweIqp3CeQ6ml4GvUEmW52OjMp9ARXdvIi4kG
FwrNIxLXNmfAv6xyh5SFRKZB2jslmolQee6VEzN2U5AASE4rPWGg5qBpEA5BE856
jE01xomtS3vRDA5ggvv57l+0D3jdGXeYQMP+PAM8Gbh9Bfk5Vjd3ngcunIIkFlJv
PiDmhlBeiBJiF3IXFMFzDvgD+HyByXZ0r2ex4CUxtFi2zRBpA/0tymZKQN11I9v4
k98Z05Vx5nr4f+gUa2k7g/H0L711ZeniV4Eh9lMxTV8+uij2PuzFGQdFjE7vWppb
M54LZrIm1yRxErnQmNfAINOPzm7wvvVbvVJCRzvor78pgQtFKQXsn/8911zdK7FW
8pw+3r4nUpjEUj8iGMq/tsxZJZVcHNFGLJBp07GmKMOzY102ZEVW7n0BdyK6NeN5
njsnGaW87Fe2i27AUpcwUxkUV3YfaX70rBbfcogRewP2fY3NPWFCj/kZHIS4Vv66
uESOmt82pZud42pmXspa88BvkcLxoEoHrXaMqVHJjIu1KH4Z02uAZPsDPYIY7a5p
q2sb2p8QwI9p2+XtZ4oobFHyVm3m1ucaW6rPAt8w2X8+oA5H8jLi8ef6o7XKxto+
9ywDjl9QKGJSAA7WxJVh6GqIcZtSkL3HgDVzN8UTlVkIPdbS8fh41GXls0IZ/Owz
bhWrLb0EP2EBOT5UFTY9a4SEdrhao27tfvHCy7C57nSE5jOKT2Ex9IOOJbtLNAXf
tL/MnUTERpSjDM0IhUikOAZsDdLeK4tUHCu7FCq1oKMiMjYdZKVsh3uEQ1mfUpH+
ZTkQKpda8ZW1D8L7ChezqE9klVo6teti1KrBBJeYn2g52vlpplvN3Oulyz7yZdSQ
lEQjNH8SXtRCz7bpp7CMFPL2HbLbhcyyAc21Hgc2a8mcKtYHfHtuH0t3ka5kz2LO
xPu2UNqyRP20OIAsWEwMFW59cv18etiHlNFDUNz5bx5SWOJTqBZ+z2R2p/Pa0gnP
Y1t5D8+wflHMRje7csPeOZT9RFX48uNJJyG3QekmF8EgpuWCMwq3L8EHKzJGhUrV
DILCGgXEIgkZSCTO6pgRWhPvt5YGuhQxfx3uVLA4tSAWlQO8On3KdujzyjGw7VSd
535jHIztMM4PAsaMVqIu2v0AODq8egtUMflImGjLVqb7kOMjCoT9YKMd/4lQf6v9
0ZRQTU//nXRbCcLFOTq174lIZ5P8KwJqcNxJ++VBDv14iEh7dmGGffIbu88Q8Sg0
leRK/gnXtcSDdvlOwgH0pKxDf8tRHbzwh5+TqYn2l/nBfhV0ycxUa9VezzhRZOhy
jPrcmTT7mcD0E33v9JgZBWykR90eA0a2o3HfaZB/kHJKJiSEnF2dgEU7BEK/sbOf
uTsybO+H7t8BuBnLr4yRbKdsWUj9XdozKplPipAtcCQKbM5mMV+rhlhsn+N6wk1K
B53hAKMph9a0rry426/iKeY+9MLvsjw56RtOlAqLchJyk5FIwd8JXGhChEZigKQh
Ztoipc3IXO1svpV1bRqAGytSB4xBe7rrSoxUa2f5iZOOLrfgxh8DTqSSyD50Gd6/
v7TLlNfbgPMuJEP1iyoTG8SWYS3aNuA8y8Kt2FqVs3akDCYqD9aM/5aZTvRR/b/9
BM3AyxbDS6r2auWqlbVBSj73s/dVVZSZi2dKiVtajhaHxlqjX9SxUvgXqAsdZprs
6wliRyqYzNosnQ2AH89+M4V/FcqAjdNbj9UnMqdekLkWQRrmhlfXPy2Zyrql8DfL
4c0VxXjlEtliIyJ0eGdBfklYanf0GxS0ogQp8EEY5UWycniki5XpaV9/+sbSQKK+
QyAG3mYhM0RjDeqRHjr/m8X6X4UKYjo0om6tfDKZBgJIdSoJRKg4044hmsoKqrke
YTPaHBrk3aPEEPaQCS98Y8ZMkiQGwCR1Wpy+LyyHqvuAoPkcOWFNYc/YMz5jIi2t
/fbynuTpaGitdSjlLBwSWx5D7Cn6LUrRzCiNw9HT3+YAVpkufkP++dDzicrRvb4Q
ghHbhlyUAXUIjL+M4Qha9xBYixwF1+54qch7tlIGUxeSlRXcdyGcVlzqR0FdBO4H
POJVTspnJmL1uf+mr7+Rqp672egtE5QE+3SREPRkG+eJyg8jg80mDt4TXUiWYmEe
tdrlAYPW7iMG7A1xKKld0Zz2EnHGwnZ+a4cSGDbCA8/8gUnxnWfs7ri+b4u7KqGt
aEFSigObmKKel8fW/9WixCZtohTK2jpmhdZ6ycQGDkRsZN5ex5Wl0OVgwKkELh6C
IBqsSs/KnQEJLqfyodhlqtDePEc8ginKC33r09y0lrqG/C8WvcKDJ52FGtDfK48S
mscG5jxY7h9VcOaG2zHPh676xtb7S3H8uf8c/9XtWvlqH7EJLSyu39q3Knzb53WT
irIwyB8yTfY3YUKrGh+mTXXW4JSVZYwU3U8guO9rOUsT84vw2/m/PiUC/PHDyNqE
RVKrzcnSNyzwht4dhMrUcuby9c1TqFSkzxdOdJZqF13OblUeqDDoAgGDxWB3q1jG
wsxRi85lmDqvhJ450eoKSKRYkUdEBABG1YoUS+C7gB+suTXkA8/gW3b6T9Aemm73
o2TBCD1uc0GmSBO5A0KWQnWfiQ6qrj7NvWQZ7/lHPpig9H1QNEOe7l40+C6U0Spo
1WSoxm45/hOdmHCSq9HuXwvYqR+KcHp83LxEGoUk0kQ2Sz+6rwEZu3uK2mSV22q2
uNWWulUaXqlnv2syP8UY4Itqu/ljtuad9MJJE/Sixh4iC7E2dOavYncPQA7L2pOb
DTXnboRxN1yjGZWS5385FJ7KfXzHwA8VSzA4zcRRtfLj2aQCM/TJb5NjH6j+Mqt2
8Zv2yQS0t7LS+h1e+c3MgHw3DVIDqq0lVeKWp74EG0M1fp1QoAnqG5boQC8SwNY4
LSl3H6wVQuMlHufOQwp3B3QdF3QRU/JWkBCGrOWam1J9OJEej1E2b28/FMWVrHhC
Mbw5wumc1WlJqqoRqXngqymCXk+uPs2DT12zes/1QIbsVAbh7rFSlQOMzs9JAkm9
381dRIB/sQWPDNk/zZoqoNnRazoKroDR78RR73Nd7P0oqdQL4WTmis9P7eP76vO/
wONffKxhyhoYsK2dE9E+ACSlE5o8buaPFlmEGmrWEbdLvvGCMckA3NH7DZU6TWm8
jr+i9k7gtqcymTi2YQWD0uWNE2l0bupVo8yYCZLakA/Vou2o70CAlvGgS/aEgv99
E3iUIIz3EmbaCgw+RUqSNXFXla8RWFehJIe4KEVuyuH84QLT6PBXQZO0nuMW8AUb
U5YHDZ0h/i0Bb9QbidZH39x/3dpppT7vQLcmJNfd2z8EjQjlJtR844wRuTHPeyI8
KhuXUW7l0kKPuYMmySiiSVlJ87++2Wg12mWHouZP1dbt9mqkRal0xnlHYnIdq8/x
4ZoB7ARsYO7TzsdfxXbDZ9DlUtCRUl+yYmTBG+lc1N0CfQ7Wye3Gg1hIMcGLINDV
sVC7bi6YphZTWYhT2GbqTAIhCUrDe/VUsi00pjX8nTvF9n45C2iAdXkeJMwC3YcK
nn5NDntnIj7NieqWalYCJDsBsYs75UXKiSXIHTpbYQhl5+YNd8Dw9WV36ifkQnkH
/rMnwvVJQOhVrT0dLtO/PK/q7lhicPl14GB9VY125e7ZvY3n1cW6x/5UhP0/8rLN
P+WYRnnYsbrtsCkdY2Xvwy5sQ1NKrZ76GPAgUXSI2eGXT2g4vSjHTbmK9RqPeSPD
cXycJ6HxT1Wg7coHRBRJIcJDI7lvolxUIJYbPWxdm42maS4vDh9xllhmxDA98/Xw
Wx1rj51gk9N3bWpUqr2gT6YitLAqSSnpGntOUD6rIkofVo07xvgG/zD/HAHbrhGU
PW7Y1gpcIvI2kXKn9xoh0xzycabgmQ+Lc3e/Q5oO59ocnvboWgXTALekDp2iMec8
pqCDi5m0LZ1fsAJ+T5njvBU+A7ag+P2DYi+oHuaml0qEIGhYlcBaep8FmGlv1HDJ
RSqyG/A9mg723zolE/6hZFotRNXwhvHnROSeX5hNMZXsA52+fuWmVXVa0qcMUkB3
GDMldwZNsTgpuwqr52FJuYIA80VUuKGwIV05TfXO54hdXspioQb/s28xaxupLKXK
H8C4HA+dZoN9qNJxF5n6q0x6OP5Nr4kgHwIqgQM8jz6w+yT/SrkXtJdHZUVcEL7U
5fi5rhg7JZA0Ol4BZfwUc744+clXXei5qyJbXk2U2R3ADb2JS8le+LsDmrD4rBii
m1DPMbJvLnjKF1WHWxoiqbJdGrfJYLoiGilDR/BATkVeaQRnducvKUxeOWM9c7HJ
qHSyNgy6HDitmSZx690EzztqLrRMmUaX45efy0/rThZ7/Ls9h2kHkfskD0x6pOLM
TwT0PvtG09T7oPtBm7gpygpIEBj2wV5QMoP3sCQdtNZrQextSazKSYoHWRUsmgvD
QFe2jT1oPYENMGokhXuLdeJKCElrcADeU5RG2AsoCUwhgrpaHwUJ8EMjcnpjZaGx
OD2F49MdKVpAl6syDeRyvHniRsHeH9yWIJgQQc5yZk6qdhuQfjDaK1pqJchfPnmq
iG8iK+TU0me8O3p76vIpllCbhQBAWqo2PtnSFq4Bxe+on7W+Upa7mb3RGGOBcWd8
e4vBUFkLitCcrTmU8Do5iqdqEbsCsS4c06z5bIwSawTG66kUIAp6ZIWFmj8Ws5ev
kiPhpE3+IqCrPiV2d5veSuPz6KzIPzwisWDyAyunjABjvcgjWlu1Sa/abH8O7YNy
x2KxtF6UQ/3pFx+khZXn3nxrUpmAwMjRfZPIvd6OpinCuQvnUeSg5CVpUnG6PRfX
PWc/4UO230ne0Rs8LAyK3N6tYCuqXoxjhUHoLsgU/Nt0jtzdz4zmGefhDZ9lGhL7
0Dy2oTxdgAvMkRa3TVFsZj6SPwckyRlw86Tkvpyk1tXJNpa8755HpsSjEn0jusGU
yKbPJF5Edoh+KXnQZ2L6DK0AtR8HW5WHIR8SWo8qqlhGJj0QSKvD8MtfRnKOVp7W
48h/n7dPElsinQV1R0Ym1wqhoAFbloKiUpBymaPNcP7W2oi2mJinDaWB2BqvuhyZ
AGdHGaMzOteJyLlPfOUE44Cwm2DJMyYObZUBYLcoLJ5EfsH+8pHDYPAjPNv0ie03
8gjMUUIazgZfi0TeAchbZg/zh0zJCSDWgYT1kFpDx0J8yFUIZKtClBMNtwk3dAFD
baEDnucv3Lc+9ATsx278FPyzXqWmh6vDjq8s/YAVSKAK5Jon/wqYRNHTxPJAoL2p
e/EyQas0NbTKsx0eUd+OBzAP0ZLKfpS4qC35YJ9W4UOArvpxYVy9WczJJoCEW5aI
52m/SkUPRVN8DCfNvAoi5Z4qGkCMNF8HWeTfdD6MfP0Km8ykv4rF0aEbQeGgV06J
E0RovOeCUVo8fQ1vJK+PnFAbbW70Nyuqf0Md2HdKY0M7OM+mUs/hWH2HAB/K+miO
7THJLrfwe9aB8GxsS9x9LLcT9qGNp+A7FiIWShJPwpotaS0xwZzDKjcVxIvkKEiU
4ecThnGXbAUY/kZrxeKia/UZrRxsDi7rWfPczUlAxoLfcy7mbIz0RAtJytA5bPQa
yAEvgdRe658tXYNPReOacKb0jyhrwTwBJlEDsx2VOBYPjUlcSrKj96qa7r1jaR85
kuJrN8L3vkfZomgnaJkqAXsbfSI7Xk7Y8F0Z+nzsCO0onFhvnAF33mNWhgAX1YM7
FXGDqrrWEpRyBawazmK34zLrVuuPZXxetpb7na6ePF9IKfIKwsCB/XjKRHvrpe9Z
u6gLOBJxoG4RmushxSwB9A8gFmiHwAbgIxJWjFmPF6B/XVwLCelRp6L2hOnY4zxU
/NzCf5wPgW1XnF4HAbW9VkUlLmKXy8WGmSbxVFjvGfWlWczTLF39FGQXPpWXT3xe
FKfP0FvxadhAM4hx9kVqnDnLdJLsNN4SIR3zJKP6JC+eyQiB71TjlwaICs11b1E+
pmimiOvyIB0umKyGoPEafOStmwAcFht8WdnyHZSEkBQrcBzPH9z/re6x9alQAnOK
85s91oh+MfUB2qdglrnKMSbvQUsYxdlfoqnzeB7nrCkreMkmsTGmUAuDEZohLtHy
/Dq7Z4Ndo17Ed+ATBseVPiCjpMQkoHR8oPerHb8u4La0HY9LbAtOwCciLwuuJaxb
Tnpn/mu6fZJjlsmHSdcoUQjkZRrNz3YKFfz9+OIJ61qoJlnRiCMj+bwi/mxMgst5
lFRpkLicqYmZtcMFDqAUZYtvXmD86fOAMMws/Qx3wTeioIwvWw1H7tHXQj76RG1E
oBlCBXyOCxLHwOrxnXZ9bf79eLif806Ggnpha+fZdaELPyWE+RfMSQuIo11TFR6+
s0bh2LcqILwFtkesr00tA++bHfjD34LM4ri5NmXWFKbKxyzuAk+GSRB571vQ1NXy
HscM9fDkwjoUk5HpkqLEDxJBWYgk4cHUxTomH27LaspgiN6xAMZb4adhK2uUEiau
wz0397kPi09exhQDZfhN7BjF7vh279UOtU3pETR7CyT6g3YfxoWeGy86kITQRxR2
vAG6Pt5fupkScwvU15W3z6BSl1IhepemICWliAE7k6xzYS/iBQa2p/mdDjoKeYGg
Gh+oyZ9uvvfCi0K2d325bGoX+/9Xqd+Pzc5KcHANnApGfdMLxNCpBf6sPxL1mnGJ
6eU5qMkhGF2lmskEekdyvDQ2hm5HKXmUFsIi28fmTICcifwyW6RgG0yyZ3F9DxU0
bQqzeiULe5a5PLgoaTLHqRSZccMdKeTRrkPd2bT1NgQ7EVuy5QjP6IC5bydxyRtT
cEAqrr1gdLCcz2SR/dGg3RNz99NdkzaP+RwiWvz2Ll+MdTILkNibBWvEkvApL3XH
VClubH9ymGu4fz7/H4X7/nNGtWocoHR3PGAf8MfEi5+Y95Qn7vaC4IaLbAHCtqG6
0bQo5ci72XWmms7LS1wulbuQEkcEJOyGlQinl+jXkKcJShWvwiQPcDiQ2zwVBNv9
PVjSVsyFcTxW+0AacPjxtR98v9WyL/L3Y7AqRHW/Z3E81zEIjs0E7ZrMfBJMHOsH
Ff96fngZBicc9s3AbjAe1yoc2KVzgUQb1hRPArsKxwRWsV4p3BPLeBilJlzb2Zbu
6LCNOWohKntcIDO7Af/c6oe+K5WENoXzoKacSltUmBNTzKaKAYADejF1znB0Yvy/
7x7GYsRfWEJyLoUe23uYRITbbSmyiT1IKLBuXeEYQmbNLTCOcZ4S65YWApBkoOvF
iemqkNVOg52dsbJlJfTYpulrl8L5vq2/TgaISf74CqlYjJ7L8wVYEx9X1OkwswTS
OzL1irk4tp4b9+YgRztut/gDqbOusXXEnPy1YYlNt84jowjTnk7T2lGOIzgH6V+t
xVRRrWDU18P2yMZvTHfbGjWNl6Wb9YDsImHftVrIiNNKEJnW7nGcXKxWJilf7ZzZ
LG78XOjjNKhW9Jbfj3dX4rJPi1Rb3IHqaCN3HhEjia470cX5RchCfZuYvsJtiBIE
slTkalsLngJ9yX39I+TiHIToJ8a+h8KYxJxuTv7TEYWCQryWWOaIT/Pla5LUGdWe
BfWpSRTpIsV0Hf2oGHls3G9Lvf+ZGSEgoTCvkvM0wG1H1NGdJtDl7khAAR2+Q/86
CvTmm0qhvXtyRriyoXUtbvsXed27HtHtGl8JiJpRSt11y61rhymsV5R8oRJYoR1k
lvpdtk6Y9FGeTXpUAY5Qy4bKjUU1kiwJiHfpEPBqrCL88a+eLsrOsdF/yQY+I5a+
Bk8dGbWFWi9eMaERlBNMYqQ1VQOt7OHVx6x4lhdjEe9IwnJW0y4RAAQaywtRZmQC
PV5CX7i0SMhINbO1+i/+WeoMsoN9kHXh/KdKz2O3c20LmE0MzGr5xXU7EoVG068x
mYrO7xU2n5xtNr5qOZJ3s6LDLcX9f9z/5qrguiBz3z4Duxcp2t+4+q3n5hoAKrjD
esKA+6jgPIzFtj41+pBYNNyUkDGf27JcM3qgpaE63Nd1urZsEH5PfAY7TZVN2e/f
Pop/ZobJBnNt5+05AeiRpJraOuxYEbRmIqdhjPoP7pM8eYVxcTeX02+zlO+NhrbO
AazgiaBbABArbDFHc2uMT5ug11zpHnLnQw6TADdPxuK4qy0Qw5MIH6r/cDLFg+JC
Atyt0cRnvit+rv6GNTIXyaZf8ewA5Kbqg7vqQfgdaT4+qnljveMOsRUXkzrdbbBf
qn4kEW0MzL08og46SSUE2V5l65HmP4Btd5p8iaR3Njj77vCEuvkMikmMlylFNevM
fQ5jJJrHlg4rw7/yohbLqeyNGZEpE5VyjMP1FhKqIHM1tMfzsmGCN5hwQXVSsQJy
LGcC66L2YJtFHcdBj3AVfsj4DWnCfFNQnWA0DMaUEeDfQZpC0W6y20QiEj35Tuqi
h4XdCw+elZ5WWmnf6ylJ8Yocd43jXz+R92jmPvMkoDBBSGZu50g8SntGmF8Qk0q6
irUHXUVlxnP743C/pVAvFnkM6r8BVfrtYGU4m7Fh3SvA1D1PWEPtWWAEsj49uj/3
1YQzu3rrYNnAWOOIEgJ0OFMCKtDEQCWpA8KfcDwqyW+MKF6BQKL2Jl487k18/Zuy
+nWTT9LyUaM5nGkd/4NdKkIRG/KCds8O0N5QMAd7X56SUpq4wOyApjnrDXiQvN0R
+hqqhqjIiGabqQrfO0e1VJT8nNESf7mz8zp5li5wOaTaSPWcdUEY3/w8sdwF+6yx
T+mcswq8JP8+AM0CNeS6WBoDDX/YDXhjFumu44tnNm4bXjQby8Vdm19XnzP03KLa
SRiC1nCOIQQJw+ukp/cwQD2hO1dIoEhUBQNOA9zMZl733SuZIuXVo/gDlyXJoLwT
JC9xEfbbE5wMshn6pEmsywC/CznC4NYId6HKBiG6DeEUfbOZKavqu8EOlhI6SRNH
8dPcnYuplsBLLO906O1X7fHqinWjCyfeCHKitl0lfdF1JiuqJ4fNw9ZxRDqDZzRB
SdsxwjZiaXhbHyKTQNeIB+vkKVllJrdPQRtiLJlVqQxSG1UL3T1XL1rbWAmHxJFF
Y5fr7BkUxBdIaYZPjdBvf5Kn/3WNpZX8TxX9jqtmtaizhyA6r4647x8bkIffcxrp
mriNEI/IIi6V2UmjJiYc+TzdckY9DvmhiGJ0DlcLxJ+ZfvBmPWhShjbNehWzvDkf
RyhE+6v/O03hMctMF/506P0dynAPWDAUOz4kBJZlUNn1zKyhYDUu1uaKu6swAxf2
5y5O7iWdN7W55eTMtBn44FFkMkFbbTJvH/yNakcD+CQ7+n5iUMIHSn+NmZ/qTjmA
gYz1oSN/fHjseahyMjp1UYJTr+sUYJat6wPNwMShL8G9hlWbiyBSz6zBHGViJ8mB
oQxqtxySX2mnQmHRAuWtOb+FbuMO/ysxQHJVIfAR9Pglu5+3miaiUP7tfAcfftHu
uuO1J/YHcF4lEDbx/HLNSoLB6BdNkQ0fZNQiera1+UFSZwUPfeI6Xw4/L9EELt7G
FP5JfT2o0oEgDYWMH9kPcldiReJFJHklLpwXMEULZpaLxaW9FL7GUC6DjojF/y38
WuvKHVIlG8+PxDqm4ZUM0aJ2Dd6xe94n5cJN9o6hWykjsbMYuOFdBX3tjSutSS91
kDZdmCmZb7C2gcNIQc5ixxWVpMFtpDDry4++f/yxDVA/HRKqq7SdqOYjlC0Ke/+d
/TbwyEaoqGwGVbQxJbCCqhUG2RKvMOTIjQsEcKGv3VI5oDU7CKBxvpR4CjMuRVYm
29gis+r4wGTYbuLz3T395Twdzg9U31trC3p2UrPi2jgeR1rt+t/uvZk2cyQ0LcyN
dm2X4O9mvopBz+LJEgE6ccSMhhXgCqnCwIsnINviUziy5Py6XQO0SyRMJXo0HDhW
Fpdz9Cq/9e3zjVZj/gbHg3caCbtw6Uwqn5JPXr3ddbBZsWW4akPtiadSiDludJ4P
w2PdbgSKeZsMuv1kQQt8okvD8ggzq1hKJLAQgsZLwNkTCrNsDDeoGQ93yWJ4Zpzc
vZXzQh/BdH/HxQtbfVBTkLeKGWbTK/u6AmevsJlwSEmUCjoQ39InyUPWT1GzJfOL
x0EQTVe5Zk5Uw/RHU4pkr4tTWhmJTh1vUL06BUt8LopCYnf5FJtqSObcXVq6Y2pp
lHrzGthaVLBll9wnezUClGn3JmwHaRpTGLavUCN6S3wnEQnjWrZSpIBxrwDLJf1t
qTHv1Q8tax5x6UFtuJFpAZQLHWvGBOYQ1w8LGwdT1iNqI8zlWxV9ndhs3D8pJz+u
AnzDEa9KvkFjQfGVdkzRdZgOOLK8Kw5SkMGwtKI5BIZXrsbSsYvmeBlxtD4rV29L
lV09JrmfXm3ikYag0rMaLFjqgqlT9e5AQerPD3k/WgSe3sY2PzX9R7Sko30OktnW
7Qi3ISsjrsFvsCG25osGWL0SSoU6vsDW6Vr/p+MUK5Npibxn4jryUkqnl3doqjSK
0LQraMorLgQI1k47+q4iefZx4vS6QA9+pWEPIpjjZqhi7EQt7/wBG9azPEh0yRS6
M6aMs79TLS0gW1sWhL/42arwauNSnRPnvJiENl4tnbhGaqif/mNdcdY6vvkfVjuM
trxK4nWu7KlQjreKEvelPexM+D4/Em1eBKC9aiOYl3PVbL28NQd1F27zFofLhsik
i0zdgO7OrflqIw+X5uucF/LLhREvtCiyM4NCYNS212SPp4yT/7UtnewZZy5zZHOY
fUQafFdcdgJoijhHva4OfneOnku3Zi1/HJgqgrWjRK5+Bayy0DCIkYBM49Z/cjYt
ITVV4Qttltaf4dkQc6JjEz9LUMVYgHLO08AjaqOzRlnLhWA3pFPNrv/N+A3bQHX5
XphGZ1y1H4GdYcCFdLF0IbVKWyKWs9SvFLwx16RZHT+k7bpf+iHIGp3VSKLvYpdB
agJGfCPqRKa1Jh1NA1je7ajmx0I3hrnk2+enreGtxiRSZ1+ChfXVfAorsFIk6jxZ
9oTiNFgoWn5tfK3BgYloA0F6Gq0lrpZibScdiBGD+XHEiz+ORJ9RxfI65ZsYI3bT
TB36kl7IBmEoZK3SaKIKoJ1OlB4IJgeqVmpt89bYgRsK/+mVuOPGOLuGkt5LeOx4
blcLBZhcrx3yyVbZT/EKB0BxIx4/oFo5PNckV1VbQT8d/MzPENpBq2qAQLQ5jXRe
uX0UlEDwn1SodVZWJzXRSQ+/htEvAzfgAaWthMgNf3TscmzfWXcDogwz4mZoZBYV
mNBjVhR6WKilTQG8jcRUcuwcM5ys6xfPmDTHuU7gxjAKSDW4wG1gITQx6zbc+4TF
QkyWMgUHpFa4Y7rdo8BiBns8mFvipFoXRHmSkDKaW9OaI+YSM0T1U3pMkwwnzT5m
AoVTsJlQ6/W2gJtTF1MPLUZ0xc2AGM8DjCAR/Y+RzZFhdgIJ8f2YwXbpQSZQhVWM
s+Q5HndiznqLWmyGOb/0ZHXUKP20oUg76XmYd9W8Xae0e6gg/kVNj/MuLSIiNeaL
5CBEnex+o7WE+FrWVj5jWwBSOVcnW3iQzhLrWkaifCprBqn6mAb4gY4MtjlY0Igl
znWWaWydbI60MkUpjWOnFdfXq+TEQJbUeeVoAlMkXCJzzEAK8y186idPhl1Bq70Q
k2bDibNKGwgJKi77V+zKqJhVZMxzXoTjMFkg40DhOTrJBaPzHzkKLhdY1jduLsu2
zFjVaWP06TVitZJJGk1SQLdyILnpfg+sW2WgiMKttWUswX6x/hbx2gG1pl5nNXvK
qDaJMxbRldV1EGU79uT0F29/ngQ5F32LKMNPxbjBlUkBSQPucJD3W11lT5kpPXYD
79m3GG5QJp6SL/ey0/qgPq6+WP++nZ8Vk0nYYL2+SzNqz3/IZ5JlCgOuBseHMSHi
PC87OITrbsLvbgn3MIRYGaxtj6qrfJEU8D3g6E39KYER4lFiXwzYcdOdfHTyWH9g
RS66q0uDtgJ5RclmjXRtZVrubqv/NgSkr/hfvAXsUW4JZF52qlQnrm50Gu85dyKE
ajwQKtRpAotFXq77ZG4l0FuxbHGgBzpnYqCgp+fYGSnwb9dMgucbyjXkNsNDeNEq
hTZNfrrCKpmbD0Us5DO3CMKg18LqqdUS8DmdGZQPltPIvAAQrcCzd/mb0wp5PEgM
KArLkIEoty3TeTwDozMkr70IAGXGDoKMxsegWKkFGrYjjkd09XY2oEwwc3Y08kZT
ZWKsUY/87U0t3ox6YkeF0tcaJZGaSmI6hw4aK/Uw4iK0UggeKQJ8aRDbErTKJCKb
iATmJD+rUPqr1/MvsdRL+dnnHMlO/2Yf0TojGttxNqK7Pqq2+/J8c4JE+SPkK7wz
dDfN5W+Ub4lnUNL5ZOlX5q6n5D/WYX/71DdqULQT4YVzk9UhQFe0zvTpZR2dmEg3
X3T6ba3GsA/UFhDhDV7zEUAX6cqiOlzzmyd3YWn2co4XRzphbYdcKu5yexlKmasC
/6fZOfygDVB81LlkdY1B8p+C/yPl2YmM0CaXX8luB2FcAza6QwTJiiKfCsE6wicJ
u4L1+tVHADDvuy/9+h2aggRkBqIHlxglADkUFDtXT1vd8qvK7QCYCT+P9tt3ucDY
uPGJEg+YTnsf4odZFT/eQIvLnxI7dYoEIokSjtEIUfAXeTj0/rau1PHXW0M6ox0R
ORNp4NIMJpyjKyppwrfDnj1lVrEfsKfnSTiZL5bMWJWpU2XDxBj10VtWks2ORuwd
92j50Jx6FVROTqXkTkhdIVvmX8U7ftabL5bnkvqCGR/DE3WJBBPDfm/xKL1sNb2B
UCeVCJXc1NxS4vDQ3kRACLQEKvByfalAQbWMkVjlqjqQ1VqaSKMapDLNEa8aD74Y
wBb1QBxKdu2vIUmSHgZfRVwhIBaFEc0WsuunptQmH03Zc897dzVD+Nm0lCoX8qGT
+MTrAori22tB4kuYRuWw+r9mKhwp4jYS0bm7HW/VJ+kB+NJRLoVBvKR+KFRtBcLm
c3c7vNS4jnwpKBkg6/4XJmnYlBfYuRTMdIyF3VaI/O0SrgefSDjfR+S3p0CqzrL8
Mycd13TboWd3Gj6vnA5azC0MxL4868L4cCbtARjLoKwV8weSAyjz2ekMoLpcO9hx
WtJyHO5L7M97HDvDsQhl8dGrtfGjiLh3XTWqyKnaIlV9InnJoQmSwce1lic2H90w
lStFlPVSTWAM73bEyTPD4cysI3QJIEcMlol5x3WZ6nz8DKgarbakArubzuM3axTe
ZopvkxEAb4XYp0oSFTsRIshS9R3BiTFJV1RSVPSGrUM56m0NbS1/Cf6I0a/6Z1YZ
Zga1fbP7Jfbdw52e+CKve4VpHW5tsbuzIZOjBZ8/WmJgKr1mEbKieQFMLQkiRDZC
zKzcbGSuuTlTas/cqOOSnpEaxQhs+1XAHww/6Gv6pqCru8X0CwK/0NySLvJ3ELMj
uIz+I6srHYSeNLT9Vv4OijdTCMcmE5SqaTOtytwUIwYU4QVrMyaFgT7Nk1h7M8gx
MHsRxksJmDOyAJQJ5lpjdjjPC0Z54hZ3zbBS9BQxLmZapgc/sK4kL1ICSPsFsurZ
z7eWpPmLfWKzdPq9xDdO1HtMABOU6AN0QkW4O4OwYT59vRCAu4HNVPwW39ajC6nz
BZFMuk3efv9R7Pq3ZooI9gcVimq1+FvrsjcLqP7+kvr8iSEfcL5pADpbRDesVnrC
2ZMPbRpbPKH8jZZESj6WZwBbVepqfuNxe1B6VSlddmuY+u3KMzMEAQpVTdOwTSTI
B7fTPcnVSYPWlf5Gnfhc/EuMr+rgr5vgWmC/5Hdqfceu5RUe/Sd3ob2d8qPv0Xdd
LKherEf3ZOEHrKVJlDpDJQ2KhkOpqW2f9dDH0lH0q6aM49tKGqrXfrNISTZ9IiVF
VnwMJip6oOhYJyQNu/oSbsDDn+bI2D8rkuiKb/ruWDivMe4P/pFSz/2Zy71+469b
CwkqP6lKsC7b/X21Cjyt29BHJyTiO6ltRCTeP+S13CYroSpv/fA6+G3iUnbD6sQF
305njQPVtRBTkM6u6CSGH2OR1Y35i8fefeeyPybsPLuxjWmAVU0IdhGwmembUZad
/yVvU8LmLBT4guIwS9uTpjQpZF4+6QQn6IMALSkxO9Z8bgkTSzQfpqXxVgVpnnPf
XTxkAGm4nK280Igdp7vg+yfysQfDbVwvnYaZiAbU4CfJ9+sB6MFXapvSlNGc08aZ
WMTG7WBgpRBECdYS/9cAZgcEEDdbI1J1d2Jfpkijt5HTKD+0JtHNG/Wq0XVxyJ5X
4BbdYVWSQRBtRz5Y6UFFKoaLf2SUYBsA1+8lOyXNbunSwtJlleimq2n8XBJIe2/H
mMDMDqXZ4/nqUERmzoStmC5hIl/iEdYTwmjs5KJpjija200ua9+bsexkGFZTgtV4
DeozRbpbUZAte4vk6eTc6thfWkhX76p14mKnGmwr1gIiILM4jqQdAVNYug5Uf3Yz
hvG8pA3FqeDJ/ppxQWcCmvsrA3dBspedWz/Dc3zBec5v3r4Si5dYsLXjADkYEdBO
1+LIB1kaNq/CjML0wYrvK+kIUij7uJef7JN6Pri+CNEFm5cK6o1C0Fvje1m2l2Pa
VYZAFVbzberL5A0wcP6EwOKDa2/jFvyrcLTd8RSTw3OjL0cZzSJJEIPdrPHM7cFN
prXw6XvajVqF/LiiUh23Sf009ksEjnFs8W7WZBvg9i6Ywxxcj+HZl8IaaIuGMC10
kpwWddMI4PT5wb1+TvV3pRW+JyOXUBp/3+E6WaSdX1Kg1jFUjC2HjtxgJvxRbsRx
HXTZaay8LxV/IFCs1nY9WAhZ18R5f+CPTkTY5ZBCWXqz4CK/XYEZBZFW/zYVONOr
N73Je/r95w6SckwEqX1IROk8AdnLme3mlaGvqpXmG+H/ASY6jrWhIBn07TZvbkG6
GPa/jm0i9g5Bpm/DXfImSo3Mb4jDFuLlPx30wQhlTg0agb7pdBZ2+z+Cb2A9cM7z
fW55jxQC8lhrGtzHMR76afBD0cXy1PKaPX8y2aOxswgGalkD7lWhbZ+TZlOu4HHn
YZrnLcFQomqAKihabCOMZBV3klkOv3uzBz/c/Dx/USugx2ZlfZnaW7fKpX2CvT74
M4Rkj1emkAgiWQvWSWP8glqk1BBE8LdT72AqZGzEDglvNphhAYmBO597hnCFmmeZ
1uNNnR4OiN4WO2VpzU6bD2EFpdvVfrZUTNFZcLpmHTs2izc4eimmRrhNFpb46PGE
XGp7O3WCGzDZf+JddzANLzeDftRGcjX2ZJmo+LLjQJMv7+6i91V4IFTBLg/pY9hU
3CIgd/IxalRV0v1KdNaKm1vWAujnPhEemDueJ2PemFnwOOn7x9NAwljsQwOOHVD6
6weE1doS9KWlSNa4KqdXXpBi6QbT3QigunAzqYsHDup7ztD41gau/WsO8IONRX0/
Et9gm5El0lyxtN3S9pVs9dKeIYk01MzXvXkfHujenYj3TJ9sjcclvOonYYOmVpKE
vUPOUnUrjt6L6mQSrdCAt6It6/pz7jkQ5kHCt/DuUIVn8NHizItdTJ29cSnZ1F6g
cDmbJlF0UK8rpeXDnmd+2jqdHc/IKebygYMBoDMHaqkrONBAZ2WFbvCC9Sa8eZ1S
vfKb/FBmjlN+NaxW6iSO/1vDq3w1CyQPbeUT8rVmgsNsE5zT0Av1fQpOBjC0Vp+o
y0KfxoYRAs7MZ2TFZfHjFP7E8m5rhMym470M2/ieIU4NBNoM90zEQgZAuCCLUjbS
7e0nJzPXe/0HdlffCzGj1K1k9ypQTZYL6GfWgu+9Fto4yBpOKu/FeVqTSdgqPMjD
N635UwkPouDQ/uzcX44qwogs6OhvDl2u7dIB6XkWCW37FblmlkrA45OGUD4lv5ov
8CEEDAB3jBHrIDwgbLc9T/+UIu5ztlSGvpvtEF8dUARZAzpq6TnJF7/DLm5t7W6y
Kl7XcVEPEy7smu+5awjo6UVzLuwsGOGWl90+d7CvZmEaVyyov6Q3I+v5D7cwZsHF
MHTYN+DB5R+u3XGhSQefV9/lIlxyMvtiN3sSF46YBaqvsDNGk7Ub3f+PT+ymCVqF
OHuG00Cjyly/La9U43XhF6SKZSmr5vnStqt0tFlJ3Rsb4KEt2O2//CLXt2wS7+95
w3wmo8tFbsTzfHerzqkOuDl8h/wnGw1tvsW1In5ghQ6e1hYswYRB5rAw52aYZnef
jNoP3jVn9s/EFqeZpsqR+5L9bxzJWKzO1fgP1Qn+kgzWuoICOr6Mjz+/hMFi6Kvi
U12Pe7rcmJpCwfGVaf9/XTjb5OAQa95YA5CEY37h8gKKSkzgGRRK0CmuYgjvzVHr
ssgQF7+47MZahIVr9IU1/MvFtl0bE4DOKig9jQFZBXuvhVHtVUiRWSJhI5Ac3srP
OjfABHj+Slf7dwHMNFwYBQ+FuSb1Zr+U2jd0GYWm2c3CfNacBgtpNfhafe1A+lwi
29h+g6yDjAYiRYl9/o1qYM1w/zF0kOVEama8pAtBU/rT99y745828iULV2ex0CQ6
WXKP8j+alZ9Pb4sKHWSBdSnne1G/q2re/Wa8OHiJOxtPRBNExFpLCmn4KxRZyFqS
esTwSawSIH0YfuC8LRJrNSuux2qbT01rmd4eGmLkv54eJqvEglZsveoApqKI3sxb
4wr8A+9/+yMLQbJgiWh6kztJysUEBWCJZZaT1tIb2pos+bb1f0KcT/KW0/QsPh+9
465q+oUkYD/6WoH+Zgm9K7eueLb4WndlMHX0q34nuDLK28e2/0LZCHz8XdhnO9ug
wUhMXs4BvXSp5EvTWll9YY8ng0lfpbAEu2Z81zwbegccY509RtaZm406q1hKY7E2
xj5aLMhuHjaigD1svKRYiQ98CDM7gaPlHLPKMT0WKIGITCiRyfdeJ90jLTjuDh/5
NqjfXAS4SitXobT49VgcgRFpd729zkYjak2h3rU6iQAwj7Goo8TxVWUK4emn15Mc
Q36jN6b01IHGR3b85vRHGxP3Wxny0lXHkpmMp+sopeSI+mNSSmUoyOqKw0ouAQhk
QvSiWmcjLWwxHfxpWccTLdb8KlUjH3spncj0/0iKyfnkskXoBxQV6W47s/BzJthg
a+lnBzSDAQsg21cQTyXS9WVPOmAbWKtdzLz9m1X7IConHAziszBGzw5SsQTwVJAc
mrI4v/dydPIGG8/znLgS3++hP5APzVOoT40f4VXFit3Mzcnr06H1Heu4YCy1ISDv
cQPt8OuGeuZhRPpHLbAw1ro3+t4YIG+gPshR8DwGjGXukGKj8YrOfEvHkVspUKaa
Uxv7FHEKY3uwI3dRPqsat4N1YOISSF9k1OBH3cor6Q+oBWpV2IGnSlltdNu5PcZ8
R408RaNmd7NbKhHkeIBKKh2ebLooYNTUWRvQVwJu4JJ801V7AVpa2UFaNRc+oZDd
WWacHjW7DxchuKnl4YNfZpv57D0xqkq5XLDoo3yoEUi/gacqlsESpekdj+SzA/UM
GojK5HtcH0JjYktCSF3dl2ogt/xdO6uCrY8wg7pOuA3e27/3+VQPfzrwWuTt+QO4
rZc9r4qFKkPYDEBtEFDw/ginajaLUdmrnuNQ6+AIEpMSxH+sKKq+IYOtM23sB8Pm
kuHtkp4g8LAGN4BTeb702NRIA03v61L2EW5QKr8UcXK3BExWQfSKcEuUd5p9VEQt
cSSJIiU5z6faFwpVsdD+UukbePnFPS1MRZ2EZpaHFvkTU085BmsUR5njxJ3yKP5G
qwZtR8sO74n1ctCLwAcCv/cSzmr+ZPkW0Ow8ENzu1Jfw+JnqD+8pxQMGqjov2ghV
W34PYlrjyLsCDkPSu9Q4hEVbYKfA76vOkU9vkiiatPctleWvmINKA17O+yc8on+E
zcfVCMZRrIGEGvkRaVuDV+88auxDwCSUXJY9+jRvIpx633JOowon/4klnWS18Ocy
/k78pXDCDHfWHM00dcTvp0XF7mkC6dVWgyUe+nOG1kAVN4j/mA97wdPtnTim3ior
TqzJKF9LmIH1mk+mEZzf+x8oEmjeoeeZbfeei17EJlMDdn8v7BgZGzk8tW6JnWj0
ipSYOGVqr+/u+lZbvQiAvQrEF72fiqlv5r6S3zcjH4KkWU15ykxbPURwBOcpS3bG
v+2jKbZyMozc9+UaxP00q9FiV8u8H8SSHWLhMOsG60t+J2l+wss74rhazfKt2qPb
UOXcpK4QMQr8fnmpm4yBHGkbf+sYBgC+2nsyPl3cZqzxuLZ58Ce8DnZ2woX2dS3b
TSwAOWdEI/f2UBjFeyQSJ2O9fO0hUEzfMkEdVSymZlsbVJvXD2e57AontdhKOVTW
f7jVEycfD/EFG6FS/jhZHIz86NY5Lax7v8UxYdYEJs16IDPZi/HefH3OgtVo70Pn
3LXZ/a9cubzV9DdhDTyjUYh4h/6DohjEuA2XO4FFQzKDQBK7nRuvu7KfwUzJawCv
B1yFQ+7jnbuqVhDHhDv7rZUxo7z8Dr6ueP8rpN94r+fgQ/FD8WjDDirscRvyomii
S/rKOt6HfnDeSB8CnOei5HMEyiPkgnrrD9KvNCSy1P6atjdnb2JrIk/Uvmd6mWvF
OEa6V58qEDNKgtFK/8WNq5Ka4iu63zvIoRoghACObX0+kScPpxSEvu2YiNrgiU4U
qHTJp5Ub9sDiguO12rahkO9usdpP0J0FepIt8LDyAcwlH2KQ5q2KbVCh5rIYs41R
fkj/xWvXkMawGvnxID5OI7tMMzbbX9T2NB7BK4KNgIDHy9mwW3X2REUcWKKRPc5R
te7pwgIQfSQfEye4GdojYzlbMUCJgGY/d8pH+9oudQlGQJtKCWOcyxLmCdXev0hA
tysmC1UAUp1THPm1ejTEMuy8TAaxdMwe5SAuEVMvVGiudmWQYTRSBsUga34QgQe/
uJ076K7553XyTch4pIfoMzwWA8pMCjJnuFu1x+uBoO3937PYIniLxZwxGKvGKWFL
7C9zDEeFRXBP3NLJJ4+emPIDZwttAaFxgPXlupal7KWxEKUw9/WotIiAgXLHYkFS
l7L0MrZTtetgjqAwhwxFMXHqRY4+1iV7m13nVewuIlAp3U1aAzkbzOUDzj5igJ+v
QiIOpAv1q1kUvGy9gz+j8osI3MhFpgRq6NeuoI+gJqac8uNqOxXmnV72GI6Mpyli
NGKgq0ovr78JIMphqjMKoyBc7LAZtZ+f9s/ahbBlmcWMG7bOSnbL1NYvK4n7Bazi
3SQGQTdPeiH8P7aMallLWczhis7ePZFchZ7bYzyfIuRbi5gowII/c1HqW61ltAJS
BuJuEt6F4uzf4tGrCemhbTUtCuqOCFenooCQB+udgSWiT9r6N/VdeUWKVD6Pe9QB
DOLHhLGRWjdIcfBy3hOeB73tnUnB80gssJcEE9wYodq4uKdSGvqGjpkKvokJtQep
kegdeYM6ywNxcHAcPGiQmWeVmuV98FX/WOavLf8ADgi4I/13k3t/wEWr+x7cAIek
EC0ci2dai2IUdr0TjeRhgXvPOrJOev7sply+ERcX2XV6DZoednIueAJgFr9KwDhq
NK79+yxkQy+vcOraB6DfaKws/5apVZYKHiWRzgP5rWjj7umDYwp9QfdG/kg9xyCS
Q3v772BtVZ3JhmEfIKeOrZr/AU4LKEqtZTF2m/GazySBmHpSM2GzOiCf28u3ExmO
Y0++T5bRS5OroscVh/m7cWDOBRIdmTDYN7BRCn0MbyNSELXOurY2aGxeiutHpU8q
9tkrzZVynbq5rkklw0CRTf9GXTOK+UFi0ngjPLS6oh8Bc2wfuD43y0Zbq94syMI6
1wPTaJNL776c5XTXCoZrd54fZ6uGlRVR1Ogf0KgcH55hIAM7oT6025J0ZBFENAMU
gNPZXg1w0/QzgtMsfGWbsIBM8ozQoGhzWaMCefYYzRFgCKGJLdKatUY2pankPksN
OPBnlMZaq4eGSF+9JZnBhKz7tNBKlvg89ZFd3q8e02GJ3Rq+BLVhrVZ76wANDG9c
9SDR697ZEH6NFVh6qv5dGo1h4GO5yP42JJJelYHlVXQns4y5XWVX4xJEIkOnSeV5
BmkPvAqYMzV/NIinZGwsBxa5JZzKbQrGdEXXbUqud5X7nMHkuSqg6aT4Fw6KcjzG
IS3eA1BXUgnpSOpt9TSfCf4c4Axz/oiaQ162dXagA9AO3LYWz8Ta9ElgWFSvIo1P
W+WTmvB2Wzvj857t/5JwA9nbFSp+cKM9iwemzFMmyuhbyHeEArna4epTt3MgLHw0
MVI1QiHkprlssR+Pnr5NVEq05waOnet2prRenMKEZ66JbcF6/S0bbD9rfS6sGg3o
9rSnd3FM5qD8UKxblNTRibM0vumQwm4hEIPalB5rMy+JzbmEnhZtcvz1WnuFGmwo
vHcDk/HW7lvKT//DSt5PpeIoXm+IaCVDWaNma9D33sC0X308lmOJ7aLi3AP08/eM
KqcAo53hT1gscZQV9DfczDdDF/NhStaCEMHlOxBHd1i/xAx6c1bMAErG6OhbEWn0
aIPoe0eDh9hPKwMjn2jKh3SMvC2CkFMrfKMMANuOrGDat89ZGMsBD0ylvtdqvA/5
syki/3c6XdcihdpqWblw3Gjbok7aaplbd+n0YKnvctlvwoie0FFxzRJcSnNFNZSf
pgEpyDQRFg3x8DS4Sq+TPvIgxYg9LcWTjEw3qi6KXMMBCwV88QiR7V2CuqFpiNCB
tGc4hLG2O8N8I+e5Tjf7MnOmncHN7nJonVEWFzZYhb9DRELeVjVy59POsTNIEKSe
Ohlv+//CMl44lowhH/cfRZCbZtFcHIntGapGNxLdQ38R2RVmnCi/LPWmj30Gz+QQ
/ISc/wqeFmx2egSiqnUU62yfldAmR0q2/PUJaoAnLv9lHeR4Onjm63D5D0NZ7XWR
LM/2BkzUtr0Sfh7hfFiU2GA3YhVTajP/MLbv2OJ3CINnw6dPo+mKxiMv3MWuC3V8
gEgg7CW953zBJlcKD3X9l8iLb7rl8xHNWVOL2sAsSmarXeMWaO/5A46rUlg+4fjh
qrrCXx6IaG41CF1FkRYeJsgag06AB6iB05aHUTIT/pvH9bj+lIh/2JrBQCNFa85+
MdiD0H/2A/25r/LQCZg7IkUxPYsP7bbo8TSh4rgu3YHVNrhcZ3dO6myNaB1FmpS1
4IzP0dv5+Ufr6f9tqDs5JhtpkmVplDh2Dsvka3EZ4gB3CLsumk1VWNtcQL4kwwaX
vepZgdSbacusTSNcpzBl6N+uRvrPwYIdN9ufFohKqOEWHWeDT1F5SWOVqlpL9lcP
R3XLTUf1PQg1bv9nybFprWjsf0PnBKlXmqum4EF/Y1zigaQN4s5g5/3j0/iPz6Nb
k8mBgSsinflHArCvJo07j718RVm6O4z/8kyzMv+g8HJBrKCNb02eKCpc9b2AdEWQ
6QeIAUaOhzl2uEWwagUyFbATeKsKsbambRFvxIqya3jksKJoOk2OOelGXCyl7ENQ
EAtZCKePHFRtm+6Qq//8okhbqNs/ftv/S3dLQQklGQqgcGg9/gpgo9LlLM8DxF0q
y9z36/W9eHnLpcmXx/tBtjmGjWcgG4sVaSmwZDa7rh5PALYQdRqIubej3PtQbUIw
ZumKr+3Bf5oLh1mwa6huWf1mjesVo3uIxVMtDwaN4LAV1rBCHpwtyplrwpul4QN0
LJVO0OPIl8hY4sbeURSsuxceynuaXUA7nxxVxyPH+Ard9+29cp+PJVNjjhm9p48R
/y3c9SzJqrAALwwuYMQldsNls3Tnl09C1qBjBdMa6m8UKhrWmgp0M9lD8wF4UbTV
XwyLL5rcO9+l+xW0aOOl9Oc+OWliELATPD9TqX2i3953cqsd7mh5IzdUV8wgyLTH
tlKVQ1OHJQPEwjMsjOFXvB+RKZ2H3NiJcdrJd8W9A4ZbEmKy4iKLDnCwi+6WBDPi
boxGYyeMdFho3bJNPI/EYcekaDJgBrHyCAcSreHYhBcYO6ldjCjQ1bT9yEvfiHGT
xCJnQm777rU77xYPCURlphGu1jpzdWbmBcIvyLu1km4vcpOOau7Gc+U8GBKGVzwL
JSk0PYoq5qTvgwtug7Idwj0+y3/qHmZT+zdJCoRECVJve4D6xDhKPoDaFLacaMne
5Cuqe5rYLHMhUu1Lyt5OFOcsarPnFH2/hoKe+/T864qfYYybo8zNzTwJaNBtXG9q
NHQBC1NVq8HZ0VrSnFpLDIe5YKZ75DcTAobt7xLgjb0NyKTzuUMjo0uR9aWRfmwp
ITXORxA9hAkb7OzDdVpnGb2aN0DD94lsnKZdzfUM1BxNGXVAwixmhWY8ciZkaQtM
yZQgv00bUGEbB233SEzx2140SNxIvITsiSJ42uNGSs1ClK2YTyHusdy9EQTyfSyi
ZZl+LEG6SDMGf8gOf1zi6EdEp6zd0Y7RKtxawnrDhp4YcCZEurfnnNn6leDmYi9M
9bz0GM2Qo6E8QJssrl8L2AoEebJ9jFaI8Lirml9c3k1MnsPhLbEZmdZrdO6b0VyA
b7ppmalhfCDxsYoo/d7bs2JuWUHrWINbeslM1osCMRSAlMvthdaOEbBSfL4XKD+T
UFi6BkDpMERuGseju/jgVYvzWAMqV5hbWrNeZepP8RFTZI90qaGXzj1lsDIcR2Qg
lNY8q1v7prpEpctCCKCgMBVA4XFiqSTc+1uOyxu3qiC8FedNu5xw7TtM4pmQI7ux
kOGWnfe+MtASQgly9rGn5wktlsZel4Xz6+oNhGpJIQN10Ztdu0PVqzPvCOE4atdg
8nATnNBo6/HD8454eT+78pe3AVeWK0hE9bgqyY2ATF6ofJHI1Lxk8Mlo73SGOMjX
MdwBeFic1yJ56Rwy/q7ZEORNf0jeSBH7y44Vqdpo8HU9XFB7z0BHah2WmhoHUB1m
Div18SzrHkkaEI1qRk42NTW/ikxhfKHWLnQssAEv9D/Z1WteqA2HaIKugdGU7Qds
WYHtc6DbIMeXoRPtGgktmjSBCKi1qvnxuuqnalbewxxFbUbTUNNbIBbmqoj4Qzm4
/RWKi17HJEnx8D+uUtTlDPpc1PI/u/RQknSobLvh3VueTycG6l5UBjODgQQz+UNe
zmk+xV6iSKCZs86LdsR/QFQyw7ySNRIeUsgibO5WEzb5AErbgDSM2b/llQsa4x4X
29iY9HZgXxNGjrDZ/OdsgKOgEZ/5uEyEf3Skljf8q9vdkKVPwFatVCILo3nenIdd
jxgDLNzqNug4ovr91ulRzSyQKmL9vXUJvsVLwR+5mXebbYKnCW9l730sP58B6Mbd
n+Q6YbNqEubBpCmBkK+wyOINo/eDgY3BMXe09OOVSrLsC52zmnudz9y10o7ejkg0
2K++kEDkN9NNtwTiVAoJBzbqWsJqmfFCKWJzWm7praXoWXvlRDgdPQ8gwJj7ahcs
ZEREKuH+Mm8g3SP07BkP3SXwNPLQ5/lNHge+qVdhMSvJ0B3e3rJJ+EfxckwXLJP7
0IlxQNb5/HsTqEghp1koqVewnLGF5RQgy4pJMs351gPLtGcYFqd21NqnDKKr2x/R
EsYDIVFtSTFPPRNARAP/7tiRE6Du/BKb6vVEPJfqtU0cHxJ2yg27m0YuAjsjhvNp
n5aUmSFKzcHIx4rOl8dUXArXicXrBOZZ+c1/YiPmk1xbxiKmVeFsd7A2Toj7v0VF
FKaE022IizAtOkcrb0d6sh8juhbqmMQTrStfyVKEEi7ytsVRzaFcP5Oyy1K4NcHQ
oRu7m1/AbME3HvwE0/PMKOmmpa5bEpO6je1t7e2z0+14CbQju60eRTPDLEWxmPLL
D/iOPvGSnk7Dx3FCqRxm/B+TIuNnDGh+zDs9o6a+dJSDeD999VgDpHnklwV5YI5T
kQDmmMja95nc8DUErXN185Xgi6Y53HUreXg+i58/qiAIjFrXppgzhIs3p42RhXdV
Ja7eu1is7PjUhwFsp2w6FG4hoLaZ+EqdPe5h6O7VfxxHWGxnZV0mZX6tNZb22uGY
UEzwk0+mp1sarv4H32MvNGMS7xgpGin0mwBLqwV3Ft+BBqRq3aWK8SbpQOShXgYx
jBeuPH9CWe29Da/By/1Af2T6+ww2H/tDxsoqcew154xYNotPD+WsOonVio2SQfiL
fEosVIVcTfhwDPLYrjcIFxHC3iUGScXehddbvQumHd1CRFrsNhFOj+6tVBsZNewo
ksCnBWlopLOu1oplhRgc68OIgDP2F4JreXIcTLexEA6yNXNOjOl2mFmqPu12e55A
hHW0Wn5d+ebqYpp1SjUVAX4VRApK8pn4oLHpBxW4GQtdWU6qTLfDeRn5s5ZW1/oX
OG5Gi0IfrjbMGFgw2v9Ic8x2j7JCb4kiNJPgDdqotPn903eqcQOBwLxbzFHHdh2e
5/6L3pePnl8o5k7E5Y4MNuakQ5RAoXVzIPPvrbCPpgzwaH7mlppNixQHFD+pOkAQ
ruogSMTWu2i2qS2v2i/ms61RFSs48u9UeC5F0TzX7xlNsWkphnPzMcnA5Cnm0uMM
crOj8YaFlXzOR7MYsxcmgplSgNhJKWgyLuRMNdZEPtUhArTDYG4RgigaonjMqaAU
pzAd9sf6lQOqAyr28gEN1jwKn7ZofMI57Ua1qHQNKItOQ5ZNGx+vsqfzCrGvCagb
8OrPbBQiGQNmP1TzJoV6v66PVXSYEEawLcRJgqDm7N98NqpuuTBAPVfD5wDR2ZDH
osj2nqArIDBjYpTI9+5m/hBuXCFRHC4ykYTA4tZyZPl1C0rWX+uRnBj3tu6TogZg
Rs1E10XzEAX8spaqIAAinhlyYr7pjCLkzID1KCJ44KauCVDGRdfFf5YEA6KK9dB3
EIQLmcevcPyDeWu5CYVoP9fvc4iRAuIiulFdEzpOjQBurJQkR46kK2PS1ktEpzn6
74ypbW6pFVV7W9fBXcO+lzd2kVoia5d/FMVArsBmZJ4e1FTFbzPiH8SGCLtLYGfK
G1HPjyC6X5rV286oSW02WKBUaTCTIz34GJontgGNL523L0AyWHqL1IbmWyCpQkrc
99o1EefMOpEQk26h9/6Zsq1hFglMxPiDRXv9Xuy7E4HJCO5wC5D1/IVTYSMdxhVf
ZEroUEVaZiMIVuLHvC6lMzjm7WV3hH3uFym+t4AAoQYjyEzMZ/mNIqHcP8wPGjz/
6X3M4b1zWOgYnKeEmLToiNfVWJzAeWpkhEkPD2E/l9uBkpOSGSB6odaX0JtbBwbn
lbMKyM7fvAXcQBgwwoAzKlKD0aHip5Y36l82tPZw2X4kS1IulahXiI9OD6BT3DIU
DC7gHI5GZ87BvsUUxHZ5C/+eCBCbf70zNbzW50+Jn3fDG0rp9w7SZGkfH0UPaEJ3
cNW5SA6RY7Af3Txk+05ZF9KViX1uWcEc7qhmQT1DZlSdx/BAsNKu9ZvltrBOTuDI
r4NXy7h8N8svJTbTbPnOpobSwu0ipQkt42ANXd6wE8qxkfHe47oubSPYe9/zVTmL
b3zsdFqho6OzJ5lp+Yqu6dBnUQatM2ejggpCYvYO0PZD4Gv7MXf9vGfQe362BRLW
5d0i+ZhtqWL/zDeNI7HyymIS6XCCTNKl/82MHk8nAo1ien5dDUZ3pdx7GSRrYXkl
ZHBerc1uV+FwyO/Blv2JxBPscWDCcroZldPpcljWOFDjtlmQZk0f3YPTmTJLyKp7
OLGbpvxOF/cDaX8gDW7Y47AQNp75rBPHrJxzykJHkrxSMD7mCwVZXZnooZpYEnPI
LZi7fiRStSk+ldFZfPG/rmbDxYWRXIJrg5ALvc9pKIzP+CMxB0VJI1euGBdt7Ukn
7fGPpLxKEIEPODEo7g98kh8YS6Ifjyvo1VfgDu9pychEdWgc6M6ZVGL0TOM36997
yYZSlMF3pIvA3/SAVarkxlRwz6rbimbqr/V55F4ZTNDmSlza6A79fLlTnQIbn/K3
uMPTgMPVmAUtj0Oa3RMQOyxR6apIYDitMx0SFbi4jveaGIIDJODGi7sw9jLbL4QH
PjO+jyOBiVQZJtq3gY+CkwtlIQWe7axHTOCTJu6FVOz0Xt3VpqkYeYi+sv091e26
SNxDHfa1L8c3SUxxClMR3JvTT11VXaMWGcQI/ZXXfowcT+SWN+9m/5LrvElPdVTI
lU0ioyFIbLsz1H1Bqzs8m2lHGBjVn06tNqMvXf4luaR4iTQZCzatlj5qNOSyrmVn
Crzou8ZTHHGn1xVkRiD+MJ7NDkqhboqXmF9Yy968BdQn90QemzdYIqJVwB8svUfr
tQ+R85yYKMh0KokLDGlpZB/4yyzom3sjpK0iY29xvP539LehQRtg39S/BLMxzuhT
zPv/q4heID/gKPRX+hZvTr/5Ci9ucj5iBrNAxDxiZPsomFH3kcOGVdgk5eglipWD
sOqAQPcrMF7aMY7GiquXKfYU8RKLP7tcAbWtxEkCy2CiD14jSLvjhCHTTIFvrdhK
eBcMsJm4aus4dIlc8DA4jCylV4CqJ7+SSp4k5bWQAqBGaaqxCcnMdpKd+McXkiF3
ASirWYgvfKShqt7oIyOE8iHsDowQD26CIHYAwAW4Ywhe3Ba72FyNcOhIFpZuL5ao
sUvsjWyGHVgNGbxDvywPezQ3/o14VXRle67TFPLxE73qgJBNX9UzS701ll9J0FP+
yvi4a4wwyXUmBO8EcYuPY7PrDWXPY/p0BkxRxzVXqjtM7xfIAKPrpU7sVL1Qc0QR
PVIdekQ+mmCjqc5p02YwvZ2PcsGUyyXdu8WjXcxyUQx849J7hXCTeoK7dJLJkS4O
++6ll2O4Wz1fBevb2vlRn7dvJseMqhaahTwSlkvWD34fkwrPmsJltzrG5HPatja4
EutGEoOCBZ2TE3w1uuotCnMxSXCxFmPtexNflne0o6Ol6eh5jrZDRc2Vw52fzeor
5QJzEZAX5E/C8UesQiSvxurxoZEYW7LYHE3U9WwDrVPT6Hq1kzbvO0yrnyRqv0ps
FvZ36CYEpSruM4kcMdjQqAytlpJe1lL/LVXLXXqfUPcHVxbczILgEEXuNiYHvqRx
+5kHH/kWEvgcRB78qPQSVUD65J3ksGvqQvLZk6FSuOFfYcWQUGOpgCZZLuJEOKaC
h0DlCEsHCGctYunsy0HFYGxPDwX3I2BQYgpcJJko5A5X7a9xCFRLDnw4Hh4sao95
d83AUTO09akBKceoj4eQLDrniv8yHwR1nfSvlX9q9t25JrUTKN/Tn1vAy/eojt2h
zPX+hmP0K0F1NzSsvtPfT1T+ni24p5IyuQI1i14WLCAn7evJNMXXMWSyHWngMEnB
f2Gam7Gy6vaKpAxH8vSElLioPiPpB5+AjdWRb42KOEg+CnSdsvKd+GoAut89rKJK
APat5kHb0dOKDr/dkr6CQCkMjo7cAU0qiHiCw5QrwhquZwQbS7bIwiDEtU3GEj1/
8ihFssAdaROGyDVm6e4Ic28OKD/eCrJxvXQbStYSTCf31SOle3AgIHifBkvouGJ9
kqXSXSiPXnxgSJnABgdkrUM3XeKMKrdsjgiHdW0TdwkKgGzrKubgXMiD0s6yFpl2
non3gH+rdZSVSw3BgTfRPMyknYBO3QMi7+IXVTsZaVzt3Ivzgep3iRMc+WuEBiff
MR7M2Vllgpq8iV64y7I0Tl0DBeOhKp+AM7NVa69wdAaHwfUuCvZxjRja/2MieLvR
0a5rcUH16zxyfNBr5GEBXr+rfQfZMAZpF/3zHMOnZXrIWSkPCIjg2h6/xBYDiJtJ
UzYA8Gq7E0UwLhtCaLtFJQnoVOlsa87AvCbvqNlGvFaB9yoO+X+WiAEcx7YCJU67
pnnxIklBsPQm8RK1KQqGtwmMcVx+YdaopRx4Zf9EnT9PHl42dSK6eitMc5PtsXbw
H6DmAdZKVaf73aiXkk4OCSkxGtxiCyrObpPd5CTZpjS7Bghtybvoy7XdwwdTQ1WB
kLIRVRL9z3gvbRmvLzXN7fRgH1wC7jI+HgSq33PpDq/osjOalcIOxwZUKQ8eoOA1
Oujz1UI7UgeNA5qk0cpJjQvz7YqmKTflvtkMoedLDjjg/sHMXdDA7R6MXLeXt1Td
8hpijMt0IgIP0tkFs98t+f/LgMOUWkPuRHfbT+qcYS0qLeDEG6pOmlFrYt1IFzkJ
hPnk2XO06hCJB4bRY+R6qv+VGgXjT2e0JOQomLay55wek71Y5wWNIAVKBfmA3U0j
psOdugJH6c7oGV5olaeww0I7HUGf1HPnX6cjMOLX0stMA5MkzNhbldAcJn7NOMSO
rAKgKrjuGfsJzZV8PhLgLu7voF+Ywv4L+maulytLEp2G2PWLq/FAJpMGTqFxB/tJ
QM1/B1pBjcqXSUMa/IIQIZ2VX21NhRmdCUGpyt3mHYnVM46Eu2dY7NBu5HD8R4S2
3oxQF/KvpWdHb04gFmNVQL9L6comD5WjCQnSHeO+v1p8R1LoGTlJgeQRgS+LEEic
jfSO+Pqn1L8eMu7NZWgxVHQnvtLjuSO8qE75FkNxLf9KS9xrDiVCRU7uCrV0ZAnv
q4uQNAdAgfn+5RKg0xZ7CCjhZpMP12kEK6BcaQU4+ve9H4u1e4yY1AQ6365iUZGW
REXqha5DZkfugVv+ZS/b6kT4BkacidIa6TAtkww/BzsExX9fNcW6NpaJ9LmA/nvI
qQ44qMDFObYE36tI47pmkUbMiGI4pP0M7PnIclBtb/G4p5pFE4L3g0D7AU50yUPI
BKneBUgCfnMTdaPsT2JC2fhZlLF+FJTKkhuf4vZHQiJC+bUShwgZdvWz+6rmqzjc
fwIvt26j7JpInZQ+X13lQ0hGGvBWl2ZKoee/U6b/h3UtRjOwr11RbwcCg+/BLgve
IOhPNeAgmkbQmxDJk8+NkgygDvs3ldjrMdTXfSGhCAeEodl1cBwr8Sx7J3xnmlUm
EnaxtpzVVDHuvUDAIM8Alb0G+Q4HbR/mM7nsOZ54LoQBFCBfB+ejZ2xOcmJAxq1d
2/tmVU5kyVCHotMkLUV7sb+lxmiZYrn525/ajYZmyNDvA80yXkPuzPgq+W16P0ZJ
fzgBm+ZFYpqrpT6UL+Df2A0cc1WvGEdHibXRQkTvIHmkmk/QGTfPrtrtKCPaf1O1
cxNy55OpeSsWnJN4kWdaXuoiS62O/yFrsAsDNefyLY/vwwClPUDiNjD28DxnOkmH
OuGbmOVgX8FzHaTl/VBD6US9kB/i5TYDUdFTzJpY/HszWYSmhTy7r9M8JBeTi7Fd
SweJl/Z1vKfS/RMmXSqjtlrzM+3/tnfGKZCwBYYTBVqSPLiBl/8pSybiGvFhHdAy
OVE/37NFybETgyfKrDczxuQg0LrvhoMu4fFUQj3sTHJWFYcEnU4w1//YdZwL25zM
UEVO3ylvu/mBFrnSuqylA7Yt5TxYgB9ukjZElJFieXOX7B//FW8AHe87BvxIMVbk
Ai/Rjf/eqnj/BKxijInt85orcOgJHfk1ccNEbIUFfhy0/uVZBsBnWprDmIS24R+6
+HAlQI/yQXGJzJkg9cbsrCyj+WbRWIX1Mm1v4C/YBsvPy8vEfq0kBfHqeBDmyblR
jF87VZjgOgu3q9/7NyVtF9G9rFtXvc8/Vf5C9raqjZjARPu5KF9S2+gZgz00wde0
BAUir3zEzK3z2cpYtuS0Aum4kvCCliYyIeXnrbFraIRtFSC5HRvQ067Qv//KfSqk
YXxb5l4CU99HhknUnr2qV4587zGT5gR2Ej6nKqmURP1STWMD6nUiiIt6JScYGXOP
MW+XRxBerNLL9Cj7vChVy1J07oiajpW8sKB7l4eD9EgTDFrnNmvSB5tHeszX3yzc
98qrpjLS+G0KV7f0EcnVWhY6UHowmr/rE3RERbaQtnZw1neljcyKS96JtQGYOo3Z
MagOfdfA0MRNvidOCW1y4Vn8+Br7MSUHhTHCeB0Z/cIfhsx+cWtC2Gr1mY7irk+S
9k5QJ8hXhYYeyPxxTwvvTm478oz47Rp9W/i9J7elRRTWG/ZqcAHxt3uQknR5dc93
m4gkx1R8wysxeWGDxbqzTXSSBNjon1Um3EX2o7NSvEqBeuZJUPVMEcE4N6Y5Cb2u
TGZ58x9QFtGtMnmTeYEgDMi0HcJIZCWfbms1/mAUQWzZNEYLyHPbLX35cLFReGSQ
/g7Qub6arxxTkcYI5+S/SkPSFKcBWC5xDNe4JpZLQy3ChoGCH8QUvMX5SNidpaxm
FB5o7sIyJtggdRdwa6M5Pk8SOccJITcbUPU0pB1PJvpQIcPrCo7p0YvVix6NrlLN
xkcF/CxSuVKrIocQjZO9VetLBqSkJXET/2I0wqIK3XLfKJqIdH3JfBNoIqkXHV12
PuhrHyTU5dru8H4/0U6WwJy9GI3Ov7S+Yktoe/o4OMHQG8LmIBkV51n3nTxm8Fko
X30pGDaoqPlDQE45sl1qJNDH+jGrnAPUz0NMth/4lKkeLEFMyaHW45OJ7OCPgUOk
KORkBIwcGTPDBP9wTwjK619SENndPuO+YGn70Och+K7ZBtnl/P2YsVZW1X3X6xDN
9byt0XJzV5GASYNBKrSh/rIHuDSdDeN5oAD6oioKFPdoKiF2OJoOHebq7g4oD6g/
8J9DXZL8PJ1c5gQWXt48W4BWitn0nclv/aVcNhovXbUPjbHhqY+TmFBpEOeJpw4Q
u/UBOKaKZxApf+Fu11eGIXxzVKyWA1/ngu+sCSNkZ41NJzwB/J01WYS9NgBaB/xg
EuG2zp4uGBSsBKlMXo6ZtBJCDNyz3zCYNhIJHgDi5Mq66W5KSEJGKMqtapZsaAeR
JeiIrfznM5NX7rwNM7nFo3kklUaZOHJeAnj+wzCjjp5wwgsezzElvnbzu54H5YnS
g72gRMFh9xDeZ9gb8G1i2KZk4SKgSNfRtNOwVPu3WUviaQGs7ay227xhPxNSYh2m
bgD1aRlmpeurlKw3R2fMgcaFI59aKO6pC3/o5K9lEpa24NpdBTcrEw6MUAidgN/b
fozkyfGcySex7EL0aPDrdlnL3/Bh3/EA87OuH+2X6ssDT/N/wFUD2D3UN7seFwPM
fykCALoLRpjTHxoiZOUH+AFb3Ahc2BEi/wJrGDnTVJpXff6UrxxVexVbVMMd66kh
borTe5z0jU66bewZni0d2fTux2CQBxRA4qNXsMLoiXpXDCQmsPRvs+88gmQ92NrD
jEG8umfBZirEFQ+KhjAfwfXL7ydtcRUE+WRYVPvg2+ABqZ/SzIaVTAv3pzS326Sl
lL0KNyp/20151UpdZuMjnq56vtSlbzcadnrUivO2A8KxNIcOJw0vmFg2qQzGFAg0
AgvhBTsQ3CX4lcsi4eEehwWZYUHFaolcsRZZ/LIZcEmyEtqbSNzudi4cFxPenKXD
XoIIvf/yE54SOn2/3a++HRrfS1eg+wOv5q/bIg2A/mO5kpWPfYWkG5KaqCjHwW+W
yuL+wa57EDMtcy6Yjb8tQkWLb0nSNWH+lY/Dec8ALnhIkW4pS1Iyk8HVW79eT4VY
khn7EXZkYIlGfl3f18jgtwb5z48DI80tSR9z/pPgH4FuwTPj9l8mTDJwVimBmAWw
7k2NQf22nHV/4EKCmFLuDr+odsiRUhDJgUPraOfon4saFfofr6yEMUMSKzXBEWUM
C8HOxula0ospXzyldBr1KAH+Q2YMPrkRqZaLKQAE2Qsoet00OPSASNQCcW0DQbWy
vrgDcG+LR3tye8kqagCMUu4MnwI2hiSNwtLvXK5rVOMx7WjOv41XMnZZu+X9F0+h
5XH7niEOHRWFTaszQTwQG945F1dI7t8mcOTIZRmxLi8fRx05Ayyxe8pNcLa7n9hG
jTcQkCkTOBti983AK0q9OQKyXs+L5GBvTP6mHd8FphdbunGpoLgufT0zgqY4Qpgb
yH1hVxH6y9agAAi4QpUuOzdaggBpDcK5ggizD1Y/Zy3f9dDz6ewsbJbkSHiKZk5l
n0FtP9Fc5kaSLVFIEPpTu1HGSKaiK1RTq3zZDhDmi1Okbksr0HhAEKLVkZJgIyt2
61hAAT/KGxpcKjQVw9AaN4i3/SZEGp+g6E7eoFVYz0YJ5UQq1Qe8rZFe6U/5IxLt
lwg28GYCW+kqpKR+YTAh1gxo/NS/IQx6Xz8Wgt5NvlULcTQIm/sfHUg9P7XBLsL2
B9x3D2JOJSCh4T+XhkQfgzsEtn7Xm4W7FvSAictYI0JpmgjOjiW70txlZQxPonHH
jg1yjv4VA+RB0HmRfz6ItD2xVOlNkSfAuYq/nceTwb3eGOfQYdGVwtkoGf7qRoez
JDAMbZy1R01p6+DWSaBucYP6fw/XQIJtxxtWpt40Kkss0Ha/e1WFY2BILdGmBQEV
b7Rb8tMOGhWHiGdaX4201grpTAutVGJUMafxfpRocXg48Vz3saTPphWiur27h2VG
PFd/FvQHbuvSJnl3kj/PfvPUVfSWft2oHH9f9KnZu0sNqtYOqhbyWvZ/glwXXoX9
jJE4ByOHobjEM33hKixwNZcYoX6cDU4keKUkUnZH6MohUQE2dvG7uMcN5I7lOdTn
XmZP23sR6Kd1ko7hq3XMmK+UI/vrfj6hi578R+H+q8J2dXrIVD21WNtbBB4BXbKX
nuEDNMGrBbGHRY6dSVdaY20mKlSW+LGIZjSquIU1UYe6qlQbrYDX3oBdB5cbBIXK
bFqZBAGbT67Puz6qrtKJ2ypQEjiWSFoacLOKeN2HSITV+gHPVXCxl7oFHWv6/rUd
dmXaKYziKp90UyEqAkzyUjXCejoxi6dUfpK9ad9G0QKUcpusgv8Qdc0kuGaFs1Nk
YMeSslhGyUlgxTK5UgqcMxDcDcz6oVGCdS0WjNTJpvrkJuDbaDA659TRd4Qyg96M
M8XJ9tFN2I9IzpJJH8sYpXpsFPWj68JucZUhe0pH/UFPAErj6OwPfElB+Xjr6n97
FLtYLlPN45402tJOMO7FEyKTW/pPSawGv7BWH9nV7IGl6WzLW7WZ72FgaNuw7NNh
/MC493Z+ZSPkjN4Cyfn9xF2Rn1lIc4bL4i4nThcgkthY2+nWCjF/0WJieHE/0c2B
Jg15tz0U1a/OQ7vzYeX0+BNVKRVC/CqcrPNUUDqwJEJetW2QgxWVLz86pLAlJeuc
NtVh1nLNDy6EaZas6K+03Fa4MyMFf66OPCLP3Ud3h4LD0KlQ+h1UYk0FwZ0ZAhsn
YZUPH4F07t4lMjalSFbaxBfXMOLevR+xBwLt8SOSANmI7pqmZ80y6wQV1Q0ySMoZ
r06U0YyGThu5J49ctDbKF3Rm07cDtjmmH6yQOCtER6RY6m43qox5q9P9u+JUbgci
tLQBT+YtNfd0+03dH/ndy5hHKP0FhvmOXrMnkrOGCGJJinkJCBjdhbcHXZruhH1q
lm32HsxE+KYlj67DpBNh+nTNJYVAC9otrDb+4CVscpBtNfygt84c1cuPsIg9NX+g
AuiG7PEiVUuhY0BLF7a9hYo821UFxSnMnUjmPxWlxIToXaZLYhcxBT1cvZsN/K1N
9ZdLNMl22WYgdDH68tRR4hwJ7qWbk45zzGp0mHWcmeTNcorNCpwg+OIv8LjJgMHf
zVHIMj+HcVyU4IGANUAnlt3DYBNqu0/DnXoqB2P0zGTkHkyLZvPzMNroQuLcSXq/
kb9mhTWHZHneDia20J7JUSc8O8AmERdAoyDzYDPej0GwIl5l2xZUxiZLtigdaRzn
hjR8dFG+v+nIKuLfZFww/ow9kr3EegBQTZwPgD+FXigGiwly2lo9nT+uufiZk2Zt
JhdwaZhQU04TpaVWD+xXSUCnJaw69abvHqY6NVcO4yHLZSQRX1LELbxxZQq6XXdH
5/NlJF3L3WQNZXtLh43EhBexVTmOxdjracTuupQR5NGPjXF6na7dT9dFG9bYx/VL
cu7j01/xgp5z68s5WFUWsTgA4nl6oeWobmb85uCIxL4bBNuv+qAym0Xx/yzaAva3
yZd3nCvu7WJ6rMKHINriQQvJAnLmhmZy7VT4mgMG1UV9AUcW+P+jwdz9ZjbaeG/q
/CWeB2wRC8CGA8Jq6WiV0DpaP28Hkb8IPaOyjbkJ48zOaokhMeZ0Na1kvLyWVKPc
5qaX5rCXgDf80OU2s87/LQtonGFqsNyuaGozY717PZg69Fi0asVpOLUhHWf7kwVt
NsIW16XJFT2OXsY3Mqnabway/VLSUgorUwJPv2VNE1EG3D2QicE+qV/Wk5JP1fW9
zVjx2KlKTOkmiXswKeIYX/FqIVuItsG+GOXxdWPq5dNSzijdTMxzKSv5SC6mgg/X
xxEm+DJG3nk5Rlu5GRrUmWDsuXH+vDNM2ZisNhvgUV/azCdoqIliCaTzTRQJU4ig
uadcnSa6qziP+bDwvFkLBTzB0PlUN0ywSjP3iNWCJnvxdJawEUCc1RPYrzh3C2Yy
gPcOIPtDgQMC2Bm+axJIMZSbk2WgOWbkWiQhIbfEFZ4vYSIco4yUlR1lIWAy36fS
AL5WAiWC45HZbQE4XKDr0hUnL3fzid/xBOOgKLOKzykNamAR0hHTJggt43Fs1RSh
92NSSE63GTlbErKf+lSACng3vZrykUII3sMOI26bQaEUhv29e84d4n2JMwP2b2ZF
rJSQPfLFXRbNk2NxVcWTQjNjZbL1DizEaSbcKZJ6h61sgZlcpOecomAv/i0rpOed
OyF4jHbAMhXymEpwapdeVwJAptAVkefeY7EingkbYJH0mBr4ajjBqVTwgx+Y2fbA
BIrJL9eWY2JO3KH/XekRiCovsFh3vUZrTfPJGxubG5zNu3q8LW4HLqrzI9o7YgPI
sYk3vXsNIsrPI3D12kz+c5/r4rSIhXaqKQ7qn1377x358mNUshyQOijU0onzEOfQ
F889/Y0Fy31r2PrglxvFd/190cwxFj07dkLltptuYYxp5i/t66PiQRn+gpqcfh+d
H718yFUQRulB+yNt5Va4m6FhQq83ZwsYef/K7Zzm/BErp/EMLRtvjHwJNnziwPOI
22jY7Spl5mrVOLPSzuO0rneqjG9XnERKYpmoywEo7cFN6X5tx1thmulfRH0zwTza
VzpFy82JYleicp4e8LU11fjRstrwUDnDaFQYVjdPw2TEvN0E/sXEMBIYjUjtc8YI
Tl3tXfCW+Mm7ZENw0IXSwMKlphRMKpLQF4HhWdQfFQYZjEZIXYwerQEp3lHXiqPk
+45F2fPtWSCc2ZVP3ABuvHQLSK7lyFvpuHrdb7FJ2UGvFtYXkGrCcz3XTS6Dsb+s
Ja6oHqLDWVoNWbwNxuToxJPUef8HAH5jhwiyQp1un5vyMdjo+NQg/N6pgsCRNvRU
8SAOvPt87pURMh88T6+JRdV9IpK6lHycN+Q2CGcC4ZpnXcDD+dPewssxZRObJrMD
T+qFlUAIjNN+pQf2bEpT8ODO9LbxOXzIfHqqxssAalY+hOyoPtd6jeSgbt7mqHhl
mak+G0pI5Oh6gr1H33X3FCuTghqX1SyNWE2KE97cYCXrol92EiY03Xadqzv6gWbI
Bm6p97UsdlIOi2uZJO3wBX88VD8JaAIXkBGXhHXWCZw9mNoWLT71/NQidJP2OVSv
Y2zip2C0kwz+QzeZNs3l5ga8jrf3FzZ3BSMAkfhK6eksm1lbOytXaNOGMcNEtUpA
NObaVpvbonupKeofJ4/mFkItzOKIELJyyKhZw0XV05M/aqMREv4etvprHF7qF3dM
0ynOtEZr2uV8Cqy6XjeSEJF0Sk1o2WTvw6SpzNUbFr073d79/p6Yy8R8nMoRMddF
eIhH8DP1C3fvYXA4ZvBZnvV37/KiikNI3oCEnSlST+chyRs99jW3h2Q5ikc25/kQ
0UUij4SHaHuQur2ERwpXLacT7D/fkqpcf+c8oAt1aB8ntF6usbG1zFRKtFeY8GAZ
Z4qdYcMoo/auE6tNna8wXJSr9mMs8tCHIGXmktAWOTS2wtN8ektA6EG7zfj39B1d
aNFEKgwsE6Fasux5hwzMXIIH6ywyG3Lrt8D52ugpWaPW5KPjAKRjTXgtFXzhexbt
Jlel/Z1QuxD+jl9SMF5x9hTwyGpV1t6Ix8ey9dVdYYHpcl8Hgia24zmqbMbASOcj
yr+iRpx3hStAPpKpyZfw4ji5JnlNKJuzBVDd4nPpMQ2lQBxilZUoe5kdLJmiiBjl
rXUSzj010Fhiz9cf+qAujAnoTWVpKP9otxgG/WlRfMaMM41Cw6Sr89clCFU1Pxcp
a2QJSZUYVzXg6ZFM+2lcs4soeYT29FNKs4UCPfyI/bLBpE7Mf7vKy4eSyayWZKtb
HKPbjVKEAu5mx5WOvHtZNNwUOlzAvw9OFJCpRe/THhM69M0ktHtyBnQYPvACXI0L
aD87NsY7CcGmmXbEsooNONC3Y5l9UxPDXnXxHK8NrOibIibPdPZwWbX157lkflSI
cQV2Fs8I9NUMohnXHd33aetrsoOIoxFS4KMy5afT5batyOA/l2Ha+sf90Mjtju7y
Ax8E6E3KIEGPipQxnxoW7hrvwJbRnV1IjRef9E577xvQYdTWEOjwQIw26npdw8eM
5RWl5GRb+J7zUtSQvGCGGD9It6KB+OPz0utiRsrKghK7wCWnWTkiBAFKdDyeGcDI
lC/pwnR+6tP48x2UMog8OudYBkpC8quthLGyhAmQKaampIOkjEoxhyWxC95AtQBy
SWQ2TzQcQfcMjb0oJuBHxPWSp4L6TrxSf7oVHpHFiTIB043Fy01+GtC/BJgzsn9b
sFtFap4B8hPk5hCU48qWfjSTQDpxak9Ho5aoBPtq4M7/D6hytzpeBrtb0OUoUxcD
Nz6RUQwzD5SZUClIb0grzDzwBtaH5UicfCTlHD5U0g2TjpkePZ3KM6tOcEFJQzDs
/8VquzlfxpHO3OxFqZhUqyQ28FJv3BiVf4yqZRo7sWvSpfsNJfunMmNz/iILRV9W
A2tZZGEgneR2d3eGaKr1kKcW3gV8Y1f/fKYKwIuUhexgSydqfcqIRi40tSADxWPL
9kcPOi2nieSB4/JoNAvDU4LFPOyc6vF5Pj7R5v6p5lITLsb5I3/TLakTamPiumC+
A5kK6LRAYielUIAjQdjHf8Nf8HZOooEcniiuug6gOO/7I0ike9nibEMJhzHnCAk2
Wp4MKwE4cZJvx7j0L/Tk8seWeKvy1sPIfa5vBJn9gzPG/qkytsVrAhGwbfbQIBgg
hwW3t/s/w6hciUAj8wwkDFZhnLiaC0bz9HUgIe/sOZBuX09Lgfa9gQr32mCp8P/d
b9oU5LsiDQBPaoph9oui5LxBjOO3EkUSfr117u8kevbmiWqoVmZir6ureXkF6aRx
yZ5cGPc7G28h0XbsZurgzGO9/TF7RnBSm/BYw4qzyEfJEv2mxwiSdSSAwSc/SWqW
RRL+8l0gCAYMMblLZo8JZ/npwQPfspH/87Ht0V/KXsny+M9m43V8fT/2UZQzE1Jt
X+gRGAor+/28yuROYatV8hPFqYXtw1fxESQeyAuidt2kvyX1gkn9eDSjUnuoFAXh
SasRajHPeSdmA59WEsGPtqqslAD3MFn/c2FmwF9akthiiPBhWYzDBsTuaZ4JOIk8
cLTLSoQJqfElTc4JQVXSDIl8B48w6k5ygwv01/TotMU8AU07hpT0Vs6QzEsrD+E4
o9awGFIbrxaF9viOri/gnMFvNafzRYR8rlIz+hrlNc5Ud5yR2nb1+8KSGtkRWVEB
dPnXwprzOCBlPPtaCj5CsUrSfGKHFu1Efp/DneCd5Thm/xPL2EQtoSIhfCpu4OOa
XaOYDMt61PX0FLIBJrSNuYfHaKOO+vSuEfcyaebsG6wLhlUY7N3/lx2jxCjdbLdJ
g2u7wZbLJ3VqVAu5+uPluSZLQiyv7SvJr283j3+LvyeRKVNeFwWVFvzA/KJvwEDN
0gd5yROVVwAulniHCPqZmCyae5ApWLtfPi92t4YCEyqHSw9dcpAZBAsHUFr2LLaC
7Ip2jDWVOXfxa1sjoX8bV/SZ38a3eYIs60cKGC85LLMmKN509US9fB+KmTSrZylm
OTDrJCjX+nQIKdxtaJyPCoGiSZw+hV3bYvbSBh7saOScEuvDEDvSgupJ0Rjp+sGk
3XoH9dZpbydZnOGF/trd8fJ7qGMOPg6h6gYaP5rigsZwBH0cQHajPN34gl9UvXlK
H9zV474WSWtLY7nlRmzp0B7RPpkF33Jovfro2+OBOeFcHVpY8yCSmaPulqJyLgDQ
tLitbkAKfSYoZFTEUxvuhwYUZonPZYWnStGzPg4lvvHiF1Mj0inzPcoN8eZEndsN
1gDjvAvIT663T9iqigPL9ZkjShrzLn8rYGemIKFJoBz3LK3q+0mhge6lAL9PKEvR
VdjW/giQjpHkdgFhHEym1ZubL0aQPFBbfmX01pG2qDlDsXg1VSpDc58EAY8gxrqR
XQfd+Jrw/NcxC4WnYnJqUlqxhnl5KTAFbKqYA3IngK4h3wK8843TWMiDorLq2buf
TBG7GxxJBNiFwhgnMwaWfdHQmCaUrAqvwcMOOoJnBt1JOiBiiKbnwF0xB02SLmzk
qGCSpvn3PW8pcR0dYRyw5zHiv1ztJCBst/o9OJ/CpI3lfWkju+bJKqmxtlDVzqvI
o2xK3kMTcjxIzUHQGz45JQ4YEGQplsPnVVCGXfKSfetSXj0P+xb4KPmpDE8OLuDk
sDjnieNj4keWa12ZyuSXWD0ErkUmm874Gbq+JgmlEqYKz4Vc8WnfijQMZmRElHRD
w4B9wS5lKPK5iN4B91EKI8xz4dhzNJ9FaFVY/GE04xKR36WvOhO9nKOP1qS7iLl7
cc2TZ6/3OLDwUxCXxaYG2AMoAF4iz2F2JAQ9BaMZd0B4DiqXwGPoJKTtOxApunBu
3LJcR0TSRi5VZfI4Wg9+1NlKimbdfuthEKWoCrhwl8AD+G0Yp8WV8Mq/7qEylkLV
ujB/mWn7Fy3sGF2W4gVi7EEMUkp1oT7PZ+HsYAxF1HNkRdPn3mMX04pAPIFNX9W1
ewSh6rJ3YapbiIwbiXlWHn45B5VN2YF6NGTMFUCIfuQNBir70sH32r1FOc2vDuji
GTH0lEeOYHwztlEy3+U5muSDgl3vgkerZSgCMszKfyoGzkaZDfWAFPvLhoEVtfp/
B643sWZr2rtSVxGn9+YMzqRBbUIGmlypwtknrsPDKs7gU7QLz+Q5ytjZDCFMDxD+
kBQYDYxYr7yyaKnYJtKNFN2nW2tHFsfRNBM00oB1hVHT44eym0uL092h5GsL16cx
p8Uz8psfLfnMZq7+WPTQTUF2/owb0HCFtPg2hLTfXVJdGQDHPRsjJSTFyVk08yGV
kISAngDrwH/z7IM17rKa/RBa0VTq1kFKedQdW/CWOe2/v6ulUxGNILVPTKYQSYB9
eJqOlsqyUWDA/MEuecoG711Dv8+pfJ9M5yr0Uu4xlQBd5RLuCgLaTJ6aKBzOCKFB
Y2axEeAsRYx6ygMiocrRh+xkU0Ze6KPANRhWRvz6yHz3voSRBzPH8PMh3gMUZRAY
KN1YmtKcC8DusYl72mlVy2h0u4qfYj4S0oLzInEGk9vd9Cy7mlHPUGM2TmCGHjD5
Qy1lFoEYwVGlfFt0gzDC9dtl6XoxjM0+JVrc/BbSqEshkP6cdz95+/ZjQEQPIZTf
C1Mgdh7Yoy0BaL3bdfTjbp8wlf+uRyT1BJcfzxSsoceh0z7ELlcek2zxNVJDADED
ECqTZjBXqnTd2/Un2HAcznSxZVdmhRm7D7vRK6gxeVo7HXSagdRWeUM303Wv0mo3
lPTxB2bAVx0Ki6K8sisRWCQuqqqaHk8O8VeREJRWub8Q2NHk2l/pBIepHoueSn0A
CR6majBYuOW0bZQmgLeNzZHO6G3hVJrwjYQsO2NJf/7QH/vHCgez4C431yeN/+OJ
6YzgjzwJZfK6C4RL/Me6eEtHJ5O+ILXPL9EjbrUvuedhMgt6aXRrkwv654pxi0yi
HzOC3+PRx34WbCYDHnJxqgdiJIQVUWgPIePk9Xu/+0J2Fxl7unJakJYjFZ9qr1Nd
4RWKHYa5ZXDYMXGrGB0uZyZlu84hvx0jD2YoMPB+Pi9GxbtZ1XjpBWyqsC0LndFp
wkdzTLORboh72MyMrxYw5/9qDyemf5PrzUwYbhy5NCIX6bXhwuMuOS10AOg25PZW
upjj/4z1ak/TL6QG6xRVmYIkovyUIdq5Jir20YvKS1jWlz0+Y8fGuZWBX4NVNm+6
0ANj/smYXC3E2rZNUepB74eDIVBG0T3+i0Gl92CR8jXYGyCdvC3l/9reoTXhBpKF
FsGfJEboTeO2UtwJaQtaUaPAppuJXb51hkQwc9Z1GGjaz3KZaVAgs5eZ+tPhjjca
PAfg9jP+Y7+2pyZRdaunN+S4jzlRaDMYAXduBdcDqfeGCzDvVkg4AhoCVDMVs08W
Z1ztpz2AA6ovk3qOWMOJnyFt0Tg3diQeLv0IIbL3Os28/1iRaMBEWGpqGnCADkuG
THSBsY/vYSdNXY4VnuRyY4R9mqTFf7q3YFSuB77m3dqp9wNIX/a78IRLPP7s6c3k
2YEidufZl+guIAIJWPfmZz04LqsTMrsjbZ1eYXGaQJPe8GMEw+D45Gb59b44v2Xm
+iBhLNDUdEa/Sng6UN719zecv8Xh5PTGzd8ew4ORlSDwOzlDt2ZX8OTxVNsBR8i5
OxEqd2gcIifZQNLGfRWMeFic1HoXjlChf1Q1qhiKzkvw1vgU8LruMTVnuvSyg1Bc
P9f4n9aUxOwnwxA4r1SiAVg7QJqryHHE/D+GU5GFfNNRuXSCgxAs8GOAn+6HtPcO
LnXxSvIDQ3hkDpRFD//6e6cYTZrBxb2FgmdKamdcIyD0FsYv7tF0bZVrLRAmd6DW
SHbx97yEcYiuURadbU9ayqkfudxS9mhE1w+KCw8mxekhVy7XZytPQu6thku+H9K1
dNfSq4zjoT0FVWm8nmEfXT9H0VUCwjb1slvAJXnUA6JbzC9g1InwCeZ34l55YvHG
MMu8QYG9WkPVQCRAyiEe8ezDTUCNJRLG/PzYNw80Ext+XN6XkIABEmwo5ZBfg+wQ
Dc9uIuYTaeff+lcnH07kpXc/tUpFy3JwDVRddHnIMs6s8lyL9PB31Ik99EU51Wbw
26pVQZFTWbrLPx5KXhpOhVGnAv/XQY9Ov5B09EATnXNA5txDIbfJE8ioiqAWXRsR
HPZOzDwj1Y50t0OUXvOGS/UoN06u3fefWzXKaQoSy24expHAe0Gi8Ox7FQx+oB+2
X4BrmTDRApCDSW44wsAw81WNLCHsEdPbYllemb2wo5Y=
`pragma protect end_protected
