��/  �c�9���M2�ޗN����=�\��X��\�UR[�<������B'��j`-��B�&&W2ȿ�N��cz���Z�~��e)����L�$!.�f�孟��������Y���l���������	�۱��P�#Ӡ���;�b�!Vo����0(�9߀�����5\h�פ�M��bsd�$YhW�c;KodT�f��
���ڢ���Ћ|/�F��@����|僙���_�mE�o�4��d�N�O��ROG|���Q��/�	��t�7z�Au��I\?���zm3��ՔB��u���Z�?��m�&R�ю>���5[��RAr<$Y&�
�7���Ǹb��B>���T��畺�F|�g��N5d�X�h��`b�`�$O�+�d���F8��&KT�L�7\����#J�t>�X�E t�`���� ڢ=�`�	[���p��5�
���$�g1���	�Ƽ2ƨ{�7��td��&���J/?�ĲZ��\�=rP��ܗ�C�tm�li*������C��E����e���tD�O�f@V��[�ʏN*ɢ���#p��}F�NS�6^�\�R��_L؂x�F�м�P:�[5��}�u;�<#Y[����[צ��<7���ׄ�0e��P��-Q1�$C�Tw�&��w�f�T����Yp�+�7�� ؟�fq�	]w��S˛z;�㝁!���]y��y؆ܕQ����y�B7���&`Yo�[{_-�W�VQ�¯E�
���|dR�B=���O�it�X�>��#o��_bmFѐ���T*p~t����8����:}����ٴ�1��0�vު|���[rd��[�����GT}	  Q�	�P���V#l�4�~am�s���Pq�O�|��K�7�p�檬�&�(��in7Iv�k�V��V���|�	�Z��kx�>�T���t
�>b<>f;�ס�yY��8AZj�^��#j8��p��=�3s����;j6L�!�|L6&��Z�0�l�x\��%�T;,*E��\*tf\��a˪$���*���-��̎9�$�)�]N��WCA	���Ttt{\㮳���7���<��M��zw�l�E�b��J�*�^������4�2��<\s+p���P�ENܴ�h�ˈ�����AH8�7��a��TK��{�}a#�+�/����Ir���q�^R(rmס�������%S�Zק{�ڸ2��+�2߰Hfu]�dOi+Vj1���W����*+�N�)��vQ�`��ɌE��-Ͱ�_�\c)���p7����#�O�'g5�*F�nV�����G�R��v����[��R����36{� ��	�q��k^2ĥ`�@�'�$�q,mk����6%��0�h���Z������j�H)�޴6��e턋�6�=�D�;r!;��LƂd����zag�q���s�5)M��\� 3?D?�(���;���%��YK�w�n_�h�L�,��7c`˄��xH)� ΈG.'�@��t�\���r]�͢�ٛ 4O�R:% ��CnS)��$!��M�Sn���U�89�⮵Ⱦ8��x��.[$_�&%��Y7��is��N^KI�]/Q%�N)�t��!��<gPO����Rl(��|�z����.� ;�^^�G�R�j�=����5`����p?��{�������E�Z�#mGӘ�^�E�,���Ul�
���Ġ��_�&�qi�s��/^F1#*"��N�(�ow��	�&�0�$@U砱 �D���9O�<�Rz-�C�,F��V����P$oy|��b�`&{���̚�D�m��o�aМr���6,��"��|5ͩ�yd�^���w����K�s�]r�,��ą���&� ��J�2�N ��!��`c�~/m��?js�<��U��\we���+o' r��������@06_������؂[�m����}w�S�k�]X�����S�j}�{�.$���JI�ÙGO��7@@M X����D�mv�}�\M���C��>]���(�������^�^XB���'�l^K<ʐ`y$y��V�%!��;>0ckV���^#�ћ�U�1x�wn�z�?�L����e�Cr���E���ȯ�p"V*�p.x3V�R�O%Uz9�j�24 |�)Q�>*��M�3��谅�Oi�|�g����F�`�^�7l�����w�.N���L�=EIQ� \���z�Lנ1�H�nU���t���/z~Hzehz��X��r��pf�5p@�C�����b�,$$� �=��o��H�A�)+�#V��"��p6ur�ת����JH��{/ԭb����8���t�37­��2_~��Ap���S0=}���U�ڜ��
1��Z+�xW�e�I�-F;VMaI���&�l��I�(�::��v�'y��Ȁ�9��5d����-� �Nl;;�NTlV|�F��J0���e~���f������`q�S�*�D�0*T=�7��<ˇ�	E��±�c�f~��i���|�#��-���0x�rb(�S��k;D��.�=c=0qة���g���1 ��?�PM�0R��V��	������\<�~���#��{��� Re}3�ə?&�\(��h`��"���#�C�7��0́cUZ0���fL�ӏ:Ԉ+�Ezԋ��V�F�޽�x\+n��!���!��t���
��~�X�� #K��x��:���##In�[�4���S� h�%k˟��1�a-����{�&b�����3@��{[�6I�`��������D.��Nİ�+���ᝇ���c(_��`�띤D�>�f��>*�V�U�t�Ɩ����_��Kkqq�R]�g�|�����MsM6�#�B�T�vz?�7j��cy+[VY+�lq/��dPRp"�x��3�Xl&�Y\����Լ��1�C�C�oj�a{�$CN��Br�(n�)��/\)������!_�b���wk��t@H�ӏk�u���y��s$E��;CZ����p�Z�9Y���rRͬ�S)�xa�tk�	8�Q �r�{0�߯����xY'H�7qv��0�f���@���qg��ù�G�Ò�Q�BCT�NX�z�����v�
���x7����я]���֨�d�{���SVgKdV�A����Mڦ$�6�o] b�!��r��4����L�+��̥(d���=��O-�۰~��SI����'�-��u~���Pot�Q���"
.��q��)����^�w@�C3٩���8k�E��3�O���7�o�-��ԯkA딥�H5~evw��]5���.
�v9��=����P@���?�q,A�o�!LFܱn��ew���l�<����팥,̥��Pa���2�U~������T�y�a����y"�睅ુ��|�k�R����r)(o�d�{�<iS�j�EhkjXy����;<8���R���l�R��r5/��`��7v��D�	�e���k��<�::�^r���x7h3`0�Z+#q{�0Fb>	����U�)��\Q��q7�e:��U�E/��^7��Z��|<$��Y����Vu��-L*�'.��s�t\��e�(1D�·Z�0�ڋP7���x�;���I)��t�K���
	<����
?.�]���g��/�iX?3ݳ���1�I������x��TH)ܖ	Sp9���T���\o���o����aUd����F'8�p�]:}��A0X�CkM��pc�:#���3�5�d�Z������8sX����R�E8ͯ�/i���H�vDm�H}<��kH|�I��a!��}��^En��K	S�'���ȼx���%E�ھS�l��5����Ͽ����9q��$�´$^��`\�@��(˞ZLf��P����" ���S7!t!�[]B�'�)Ha~Ӱ/!6�"�<�q��r�E$�Lb j����a~���5'���;�ܓ.��(�u5Nsq[H����Z.!mpE�_��J�T��٠�[�1�����\"�JQ���	z��<WO�t�K�l����T�ϻŒ�S���K�x�@B�9�޷ɫ��?"C����-�0����hj�$��FTexpӉ\C�q�i���IR̢�g1�`:�� :�r���fn��v^�����P��3����C���0�n����@lo`�M�%�H!"���ܔf:m;��&1�o�/2"˳��Ja�-�"`l_Ν�z�� )a�b��-�S��F`����$����ZJO�j̐o<O�u�P"hx��".����{��r�"H~��݊5�W�����(��>+t��μh�/�;����F�%-|$K����ңp��-��t<����o�1R�ϰ��9�#\�� ���7��i����fP
6�/�U�'�`Q�)j�}V*���aN�V��,9�/ýd*"=��
�2�à�5H����_��C��H4	]-��tʣ�zav� �7�K�URG�� z���܅�����7�\���
aF@M@�\IO}�zم���H�"�7���^�7��1��w����nĝ�*�����tJL;����>N'�,Ŗ�&�/��^�mK�f�y�m�2+�lyM�A�I���Gݶ��ZOC�f�[M\ˊmÕ�b}Jq{�G��b�]�𶘹�Z%��'��S�A졊P�X�ߥ��x�02�;.���
¡��jڔ�*/bxmx��ϓQ��7,c�28��C��9{`��/��Aa�$~Y_�1"���D�����MV����O���AWgQo~�
[�d��Η��w?m�[H�:X�`G�CM[؃� ��̘�_�W[�sEVa�<x:�׾z�R+W!a�7 b�N��t�^��Y��S�^~Ҿ���!.�2�u���|��,�&�~�$qF/�)����Y\�to����1�/���3�bTԽ�v�rU�7<���.���{@&xv�"vA��Ӎ�D���6`���'�
nT��޹�C,�S�~<��A|���^�G�v��zJS|��EP���dW�T����8�`k����y��`�,@G2��y�D���1�rs��=@�M��lq�+L��_���P�ϻE;����|ՠc�%��Ū���x5�56X�!���y��8Q �V�\��?�t��*C�T��.z��i	����Y�-��T4���p��6!qI��5�&���,��;�L$��`�������S>=M^2���2���:2nf,�|FB3Gs
j|��}n�wn��oM���������s��VUƸ9h����������k9q�N^�A�l>a{�6�@�4���h;v��8�LA�0im�dݠK+��D�4Q��]�[�N��1k����d��Aa���[���R�#���k���|�h�'>��5�O��2"�_R�K�!(�W`��&�5m����"Xzjߩi���U>�	�c�ӸΝ؛Z9�t=��l�b '�@�B]� ��>I�ݽ"Co�(�RHF¿6�d�3��&����K�ǔ[�� ���G1�3����|�?&'V��r�H�-��{�-v#�z�������ν�H,�C��$�����	�=]I��}CJ��]S��^���}2sg�Jiq�	~V���6���xF�-��Ln�,�`�	݆�
S��9ӹj�hwU��7ʶ/x��6d֧T�����!By���d� �Z@aR��������.���I֯4!�c|�]����=�~ H���(iZl̟����8(���,��Az+���,��>�����Z�6nƯu1���,o	{V�L̒n�rWQ�:Кب}�K�j����S���^�E�������B�&�q<�]!�_�{W��(�U�usbBH�}[�%�N��b�n�o�k�8���6��#������p�n��:5�۠!U_E8S�l�)k�PnY�S�P�vԆq5p���}�7�VM���!���W6�z�B��2�`Qow�)v���<�@	�wcUL��>W����T��=ȘX�?���f}�7r �>�
+ dg�*�}j�΃HҌ��\=��i�����(��~���a3 �h�k�|�H5�+��i��[	��1-_�sݩd�v`�rщ C�܌����f�͑�b���D���_ڔ��
u� G&#�{���.����^5�=E��#�s2e�q���bi�(�����旆7��u��|vQ��h�5bjf��־{���d%������d)-������!��dlu覫���#.i��g��u�����sU�9�HE$���,�n�82h�؃�����u?d��p�HÇ�s�Cv�ܧl�*�j+B�Q`0�:������0���+W�!�&@��J�-=s'���}�Xr}?�E�ս��i��[`j}��:UȲG����}�v�ؾnQ��2,n�M��7'���@��:��[\w�uL<��|��2D��w��i0?iLr�����tb�8�Cnk��t��G]�y�X���ZO7w���~Z6���ź�g���}�QA��A�R�QW��#�z�������o�A���リ�8+��]{�����*��6��X\Ǒ�m_!��%�r0���]c:q&��q�g ���_qs�ö:T�����8kβZ��'���%�VK��KgW��UQt�R �ÜY���D�}�Y�(Q��%��6��g�V����\`�H�[0�5���,f^��^bWZ����Z�6�w����˼�/�2\H�/or<���'�X�G���\[�x�ݰ��b���M�M*�x���vI���|i�>�#4J�z�\�O� OW�d�G�Т�����0mL����ss�L�u�ͷli�<=��e~��(���S�����~���9>��u2Ihf���1��Ppƫ��m0X�(mCA4��p��
����[��=�Il�p�<z\������|Z?�ė�x�;�i:ڿ��ƅ*�h�	 E]��OlkQã�.d6�r��_z��)��V�y� �����.�X\�q��I��_Y���9����)
�|Ő�����sj��Ϣ�n��|��u�U��,Z��	�B�7&¾&�{�QPځ�.GP��ќJw�e�����EcN�L�.�t��'�Xư�����*�h(����j1T��-ۥM~SBkp$Bs:�K�DqEL�9ʃ����"Kb�*U�AYǙ5Z��x�X�n�$d����m�f9�7�T�X'��J[�7�W⑟1&R�&&�_M���_�X��O����!FԴgܴ��҅ ���p��f�n"�>}`*�_�P�����*l�������ҍ�
��@ܳ�w钅l��e_�
1Ğ����+V��`F�.��CE5��\Fv���t�h��T}���;*����7�qf-:�e���8�T"�m�}K�[�^�IV�9a�o�
7+w=3��|\=�'k�����1������H�m`�@�3<��]|���d��&8U�NC4R�;��[�.ҍ��N��F�{.�A�Ӟ�--��/���j[jS(��(�5�?������N[�st�ia�P	u^�^��ҕ��E��%���v�#��*�N8�P��F��yp~C
������Ǒ#�i@I�=�ɴ��}lÍӆ�?�OV;�|� �IL�.q�/���p��,���*�u�/x�K[�E����>z��7m��**�ӹ,��ɼ:s,��o"��B
*���T��!��+n����Rp�tZR_a�M m�^3,	�܈[�*���IDI�@�D9�-�lJ��"v�̜`j�pU@��J��
F��C�Q���!���$��w#��/� �m!�wp�SJə��8dD����Wu$D�s�����[��f�R�5����ъ��A\w���]
��`j�
����f����<�ή�<� ��X
�Se�#���z��������	f����9��%t�u�y��%����
�)'�u:�o��Ӵ���X���������x&��]A.�#Bd9��6�|kF������N��t1[bME6��!9���QX�)BQvѺ1 �� ���q�%'��o��F�v<�/o�X��"	ո������
0�A���&�DBJ��x`d��B�x�Ư�B􁑩���I�{/|%�礿�A�ᴚ�~����>�PB�'�=���0j05��S����2���sn_Cq�.��'�j��<�&��q�`^���YB~�S�1�X+�S.4fRc	n$%
Vc�� h ��r�&�m�S}L��-��D��2tV�a�9	N�Ck�:�@����hjKGD�4�<��@����0?=���Aq�3�<���e?��q.�N��ǜ����U!������i����ԳO(�D�gs�B�<6G��b��x�Z���^��.��b�_ �>�\>��%/m~�}��ׁCߙ��2�(�6��-���k	�[��J�iI�]`!��Y�=��O��,>Q�h�	/U��e��f�f�iW����	�a�Q�H�[{%H�Ƚ[m����ڐH\���7����.U�6��Z������Ƚ�#XsR�R�`�-;0��폃O<�d��T�N"4	a��A��@E�=�l�Y]iv��#M.����^�� �$d;�J�fZ��2&c�n�[.�6�w7��x�ӝ�zv���N�w��K�r3�y�s�=�g>��1S{/�0fU���S�p1�*�yVA����c�9	���B�bI�}��Zmdio�"GE�_]\���� � =�X/*�9p
�@�]{ղ\T���+;�7����7��$�-��(�ȫ���@�VEDt���׀m�W-^��#9R�<m��M�wC_��
"H
w!��Ho�j�iLF�0��W"u^n�6������nX�i�i��b5§�D`�^_��\O��Z���bZ:�E����(dI�ڤ�1�b��uS�bu��Re���'���}�>�i��[�-_+�x�>+�R�{��ih���A>�	#�ģ�����U�5�Ӵ6|�5��1�"
��	�g��=�e����
�T�kVІ�.�H�x��Վ� �
��W&��|�Q��6��
k�����"�{{�&��d�6~�2��U�!Ч6�4pv�צ�}@��2��9��_�{�t�R�d��y6�-��Q�-$YG4ѝ�o�s]ئU�l�F[Ê(%�'_�q�D|<Y�%f�3���0jE��i8=�����������sJ����N�J���C���Ð
�����5[��v!���"�"�%w�fvo�=�ڷ�!��u�53[�0��֧�V|�MO|2C
ME�K�xg��p�]y3K\h��5�{�@�-ϙ]l��>4�sGy�S��>�B��\�*=����팿C����"KA�L�����4�ɦ���.�<b^ǖ.�����M�������~�k2r�ZV���-�*�x0�F��!e��\{Rl-l�6������)rJ4lCSz,�Hݴj6�
]aL8���E
�m���㷙:q�9+bz�&�zt	z-�ح*m4�2�?9LH$�o'��qe(deڑ��C�����$�����a���v,�5M֝0�4����Z�E��YG6V���5fttV��x�B̘􄽗c�L�����Ջ�X��p��[�A�G��X�d4�i��v�^$ q�����5�{?"�z��=�� ���k�s/�FN�oz$��²�|ڂ��� m�+�)UY��
��5Tr��	:/Ѭ��DZ������)�A債�_�z�;�^ӒWa+jk�����0?&��a�91hL�#{s7��(p��4R�l-��g��:�It%O5Le�Pݍ(���	W�טMFT	 ��#�VKS��c2�0b�N��w^�����p��2fV�����"�E�E�Po��!��V��c2����-�L�&���jq7�E�<q�jWM��DA/����v/��b�~ d0ܙ�1
W�'����U��M���dr�:�Y@�)MNW{[���)�&��%'�����Xu���C6�}���Se^�4"�pR��I,辊�M{�|�z�;�Ր�[w
���O��.o6�����߆�F��P�g��-�����7հKէi~<\m�pm��mT�1]Ff�����	6��XE��A�I����y��M��c�&��<�1�Ff�S����(�D����\ND[�����5��yU���EN��}91"����Ҩ#~�*�Wy�o��e�AM��N�ɝ�i$�G����.��̺��Z���8!K5͗v�Mi�IM;������g^��M<.�40"ELq��a:}@4٠x�cɳ]!�]a^㝘,"0�gEK�4`�3����d�P
�o3�H@��|?LS�YFl_�C$X�t��A�Y��4� c�0��﫤��mݏ��7�A���f��rp��ϛ�%�cz�$� X !��}背�ԁ�y�| ��!�C���4��3$�[ ciKL9�6�M!o�̯/�S���I��p2_ZY��whB#�SqY�Ͼfo�	4�@.PQ�٧`���~np#rH
 �&�q��^���2��X�EN����Vv���m��T�k�"64#�U�o�
&� 30L�@h���h𭇐����a�i��G��4�%"W��#��K�)���Ny�0o����6�mک�3�JL'�z����º��	z
U=���Z
3�yƝ���T����d�oF�t�\xi־RC��Än��`��7й���![��5[�G*���@�F�U��
4"\Z8c8"R��7���a�Q�aA�M�V�#�#�"��&�r$�����m��
YOr/tU�5hp�k"����0	�������[��灐K��a��Lf��A3=�MQ���,�_R5~H�-j����P�x�i��V,��Zyx[��>Pn�*����i���^"N�õqK`�ɫ�Ї���Kv�F�O%[�P�H����}8�Ä�g���#��S1���L!K��ZS��Ґ9��Q8/���i9��r���jЌO���	���	<�#�b�Nn���l@>Ȗ���"ү�чa�������QV�Q�КUH@Y�.��:Q;l��#E�{chb��$i��_=���.2��g����n�ۇ��(b�.������L.�]?��MM��yBmU�5��6��P�)$��1�usUy���%�B��6�3�8��RAV��'[Sa����
k�q�)[�E��xF�SX﴿3�t�N�pY�!{�Y�i�
�
&ggjuEʥh�I�G��&�=d�fA`g�g�x��/6X"d���ߞ`����u�a����o� Ia^�E�y	� ���6����.�4� ����.��r�8���ɯ�4M{�:0
�n�5(�H7*U	�5�b����%�����}d-�(��?��h2�`��X�-�&n7�{fL��WdO|"��*��"oɍG����]��n q�z�a������KI�1E �L|����L"��nk���$����%N�0���ˮ`����jJv"��X�|���TÀ��+��>��(�^g.멻����R3�^�	U��Ջp��������{�s��]I,��iEu�Ixs0�+G6�>�;�o��
�ZR�(�K��4�#s0��L�>|��yK�4k�R�� ��F6�+`CR�L��=�M��Cf6���8�9RF�����5���T���}�F�T�o[J���mrS=	��#c���ρ�j��d�9�	um
�zj��ly�~�oX�\5�5��O:푪��ο������ɹ�����������a�}�0b����x[��8!PEq�Y�h� u7עO�r�R%�E��H槐U��R�G����i��z��t�����wuUW�W��� Ն��x�U�t6=P@�m��h�vs<0#�0�M�-�r���3�KPHT���b�.�Ť��*�Q���e�TQA����}q%:��r����z<`{��zV�&ܲ��^��RoD��|�ߧ��|T���"�<��*p�!��oa|J�w�/�X �TS2B̻+��'�)�-ONԯy�nwqz��83=y�߮vO�CU�wB���Ne��s��r�(�ou���ޓ罥ێ��O!����k�)y	󡝦���$���^5ɥȘ������%�Sk��P.��&MD5�&���)���_t��h�p���*�z�('�̱o唻���ԩ�|���:VWԌ@���_
�ߠ�|+�sɵ�����P�1a������(jw�s�z�����ϸ��;���m:4r[DGZ�� -9��Et�|�y(���� w5�r�M��F����Px*�|(n�S���Ȁ�n��!�F��LU'ǲN�-����Yo.�+����e�XБmˠ�j�t�H�~Ǵ�t1�em�n����9k�:cs�������i"�^F������2�0���~���J�awg�.\<��摍 ��+vZ��3O�NK�-<o�6��b�X7��}���S��"�3�_�y:����kmQuv<c<A� e������%j���X/����L��Vt�OŦtQv�o-��=��r2�$�	$2�7�ںG�����;���/��'�u��ſ|��%�hx��v�6)�Ģ�8�F&B*<D�Ȯ��T,�X17?y�s���"�	6 �(|O����x_,�[8f�ƪ��D|gHn5�I���}�#���-T ���T��\$
-�Ҟ�� �5 �8��fOM�ǟW�.��7�hmxGJ�K
aP�����0R)q7g^�?�9!&"S��+%h��\����6k}���=����������ʆ�l:��V�mZ��K�,:�� ��z����'5�"_{O���>��#�q�52�f�q$� ��e���A@��͂��J��d���I&T��m��䀖�3�|<�'�)���ܢ�~�`u��MO��#8�V\���V����m��)��[�S���by�f�@�!!��j����`�уBiڎ��8�{�K�'6v�����!+o��g1�N���:ui�+I4;����g�����i�˨�7�w��Q���lL�[���ŉ}n�S<�s�"���z:��z�W��#  �d�J���������L?���H|�g[>�HՑ�H���4pA�WF��f�S��K
�  f��G.
��Mܾ��G�tP�qe�zI�����$�jTЖ2q%+�3���@��OVΑ���^�6yn���x�w��uK*/xaU
g�a��<��u͸�l2EJ��}4ė�rfАu:o�j�F�*.]��\?Xd�\фz����1��p�'9�bΟ^�6�M��3FM�Nz���zF<a���<��N'H���V�͌՗�$�v�j�]�~=����;�MK��[pRa���}���
��xs0sr�0��k�7G^2��`&+G�om[=�Ā��qϊ��n��θ��H�$�ҰN{�!���ɽ��}�u�z�+{�ZZB��T4�X����G��	Շtph��F�`���ү]'P�N��o}��m=c�8�M�k��J���॑�(���Տ�fT��Eѧvi�#k�ԢW0���?ѥ��l͘�5�Л�
��ٸ{0g&�58�4a�g�j(2X���'/�����!��Z��B�C��?�krFb񆛆�Ԃ�a�P��۶?�v�V��eg)��q@4�z8��_V�Eb��Ņp������I�UшA.х4�kE�4�\Z6�y��?14M/ �ֆ|W��L��W�GP��)�I�c��}5B�Ϋ��l���|��{�n�pV�W�GBr���~e@MĄ�}
�h���c������	�g<�DEz1�|�,fuPDo� J�A�4�(}?A��2!�jQJ��dy-�����m�_π�ћ��]����Ġ5���b���:*�ϧ����ߓ`&Tw샌h�)�ݺgoށ�V �'�T�8�??��W��冄�C-��y���3$y�˂L:�h	L yn �֯'r3�<Nq.����0��zQ�a�zc�a�&,0��^��P8Q�{@��%��MVg���y%�u��C������zo�3GQ�����D�-x�&�g�=��n*������I��WQ4�2i�����Z�2\�`��K^*�Nu�fZT�)�Ŷ��1���l~f>�"��R�s�AL���3嫥�f�CL���:��KL˾XP�������+����mW0���Dr#����#�Ö�|%g�dx�[),��8L���Bȭ�-�T0O�w ��T}(�4Ld�cWY���]��f|��a�]BX���?*�b�*$�4Q5�����!-I���I�Iܦ�rP�*)wƑ<�Qt���Y�dZm^i��+��F�j��gyzAu��i �MHg�`%�N�c����D�E�R��8l&@�|͇tb&�E�n�ȷo}L��s�`���Z�R<��ix�g����@#"�:x�l�C|���[!˰z�َ��b���fk#��6m��䐯 AY��D.ȯ�2�;����`����2�T�WsQ��3�� C�"b �z+a �%��!�bZ������r<8�rW��`����o�VY|����\ۯ`v	���V��W������+Ю��R�?�3���]	�{��Y�_"3i����ޔ���J]x&=�69#	�~yW��O$��	t$-�\V�̵]���yr7A΂��_����
��)D�Z�5 Q���e!�������iR�A���}X�������r��s�t�Ӝv��mC���vc|�c�����0���p'��i
��;���˧&�9��a��9Q��Gy�8ż	LO/}���{efYA#��`S�ʍ�Å�ށ ���P�m�h��Y��*��l�³Q�{�ZI��iNs}>_.�W�F�3 g\F��I;T�40o��=-rѺh��)f+�Jx�K���Eߓ���/��5M.���7�3JޥM�����E�C��`Ԇ�~q4��~~ͣo~��Fo���x55i?��R�T�;��o��/$������m�A�^��аo̼7��q���+�wݲON�I�������ckV��@?~��3 �"gP��|�f�<�׵s/H��S8��w�����@Jl�OU��'R�+�Hb߃�=�UrX��'������k��lWe�o��Q{4����������F9P6�}@��ڀ�6=ȼ��{�pP�[s�U��Y(�D���uK�z<Þ��v�l����v�N�@��b��R��A�-3�@��L&\�+�pqu�lzd"�J�3��'���8͟0
����!9�65������n�OCZ;�X8�,,�����mbkN�bo�ǘ���mj;'�mF���>|��=q��-�����ы��/ˌ.���.�d+�F��d"R�����*b���g�4�O�K o�)���[i:��:Z�5E���#��_���e��M�p4Y@�Ћ��["���<��ң�-S����A�c���s[�-+ϛ2a2��<�6`��ӨD[�]�0<��g.n.��R"�@�I��k 3�[;5�����Id�PR�x�O�