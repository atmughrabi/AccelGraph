// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CAdXbIX1AGFVE8rRCxmUqS5SFQ9VvdzG291V4pMkmGVbus0n8aSTCVtzZ7AwMX4d
IT0st60SBRWk8VWixK0WXhX9Cy89rwO+6SimIOi/kB/4QJpScde3K6U8gS1FVj+s
fxlUAk8qmNA8xVQ+PzsK8yOO6t/Qv5Yq2FpxGcKef2w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11616)
AiR97OR9kjUknsdtptWM7QE6yuRt2vsZw1stQ/rBjJw2e/nuhCYnCQtDClwnYH9d
zKzESL624IKnR4uAIFx23yfzJW1UKDAlI+rC3QpbeR/LxRbBBLRM/AVPRHZMiVJW
x4RzsmVMjrnsOy2xELPMRIBfvYgJHPn1O7VpgbbeB/RYbojOzKI2rhHFfQc42nih
5XUDqs3ec5szYFmpFL9JH9p9Iy1OM/DQ1+X0jS4QFSWnmqzCelLGM+yF629K9Fgh
yuxitpgQ5tAl0g4Rnd4cGzRI/BqMvSpxPIO5zod5PI+EOQwEHPaxaW4ZJFXf6TN1
VthX29oSfg8W3MaPuD0ZLnElfi/DkYWkGoopL4Fy2ORERFfRP+SqOOkYyiQRtD7I
d7AArp36+SKgL8ZeTTP3usblsDK4JA0tp1VQhp1RSmqc+a20uh/bfoOvT2v3KVwP
pLtSaSB/cN8lq5l8BnDxowVL61gYztIAPaJgCqSsJ5ibjQnOWB/tUd9E56H7GAeY
ZSfqYE6Me97VBXouqHSl2dmn3kXsuG3VZQ12esw25H3yqpBkucwnwZS0/OJip/S6
JR8OG3uAI+fDcleqxWp1G0qifIe9HMess+84TB89Ze1VXTWYQvHAqh8ftj3uUrra
vnNfiPjvn4rV0Ho0KyYM88XY4CLnZ5nD9HdNGbXzDU5ukFtS2BKGkjUY6+CXJe2x
R4PlqsqS9nwlThH+QXEolww8a8ECWQbiz0bhg9jYPtA8+3IpVd+a1XNi2AmKd3Z7
KseUuJeucZkNwp/BqzI+SbAHaeaGgOB/jHvOWfCyZOUhU/hYUj9bc6moegw98FxM
QO076frdqD1aOx0ZIpZ0BgYEE7EeWAUxN68u/IdGw3p76muHYvxe3OgK5sf5q2wr
obTSxqEKr7ifSo0hmYPOsvTIZYXSjqMlIVnWLFc2efxIs+WqbwHSS9qph9s9pQZb
5FctLlpDJU8PM6iFlSbDLxpY3zx72VB3vodArlZLqq4uqX6S99MsiOciUGiSIexV
mh3OD8eelBfdtYSIE/gg7JPktrAcTjmko6WtZ0cmC1oXBlfdo7iWGqIqmj9PdbVf
xMCbbN8lRvTGJfaa+7cotfN2Eoy+GKMp9j9QceOpqUD9Vg+Hk/Hr+PT6r9cdhaOU
JfUb03IvqkaSMqMEI1S6CLdyj9/0W6FyK0oOAs/ApxaoTYeZdQRk8dhD52OfyRhx
n6eWVBGUkL40aE4Ub50TbrEb6suZbrXe6Q/SWwoCo+Cr7XljrnM4FwQ/gug+yhwy
DfyzThfVEZUwMT5RM1I/T9veLr4zx8iQES8aOsr/7ZwjhiTiEsw5HZqGcAkmiuI1
0nLQYw+LrY7dA/106KOk9dq9VQRm6yRaWpT+ArVLpxkujYoxuj77oRDcu2SNhYF6
Zl0xhm1hhTGaRX7XaslxxnZOVMIVCeTnj/K0njteehcJWhY/vCQM1XTw1N+rQMVK
CbBlV1Dz/9Vr0SJcEyI+gRmFpwQoxSTRnzGnK5E9EQmz5cqZ46mkYqzOM55ihbXE
nnIMby+LAWLOJc7/J7U+70IKIrl3HjWNjR4ZKnhKupvHEntlw8s2rX794zhIHw3h
9yNKVUbwtsVF+XK/QBM/w9rc4xrqqgjwV31es0iqZ3RM4HomUmQayZzX+pVcDG3b
X8bB9r28gSEqpjn5nSuvXFO7X2zJO8Dg3wOP9l7eRtR7waSEsPbxfdl3DvmMhX9i
Dsq+Exrlngs9gh0EHfmWezimWNb5qtsYYipyBcFRMdMDg2Obn0NIVUEgB35OHe7l
ohTuRkDiHcoMxjvF2kInXJpxWJW0Yq/GSPyjdvH7iAR4PBqMaoa5bo+uzzBNLcK6
HqJAjtgCD4gxLvLGBCbBwuuTVUu/tVq+uw2ZoQ9U0tvqSIIXMiAqxOQNI8z8whkz
k9NS44IdBedzp+aidAonkKLS4UERf6SbWi7uDC0tmKY4v0/RqLrNLESx8POwylfj
xwwmtzUVpsi9qj9SyDQn1FbliQWTkCB30L4fIej5+RvjWaQIeSbO7PA6Znk0VRMn
M2Eo9/QyQofxD2KF3kZsANn//575ga81iF0C80HD+t/+5/cbx79wNT8QuHgWBR+b
5/KwkWJsMVM9rKXhBi0Ibn9FIaxrZTGFnCMX6lEFHUTpT85PubvuUtc337tKPEW1
lLKBLXGUFdJ7lsg1BTpvwtrs5T2m6GPOUGZhD5ZwakYf4G0LFJO4wM2y6/wMju4P
+r9QoSXi69gy9riubTE9Ev7cLoBxG0EFeCzvwgGeQTVG5uzCjmJlY77RJtXpsT2F
GrSCWrM9fZ19s3NGNe7dhf6I/PJ4ylfweVrikh6+p7FUqx+HznsgA6fFq3d+Tsdk
fSMTkRDfq2lNYbjzj1hu+gjaxr00UHhd6U2xszVzI5ICj2GgUrLZ/PezZiOGt3PQ
75aEywRUn8IyCB3bH2vzSNN2HmjI7sIsBcvz/u7JloaztuqEJYE7ts/H0W5heNTI
Y95VGY+yQdOxiI9+2BhI+okkWwn3D3x2RuglKa00Ttycw0vngbS8ucYB9DpgouS2
q9tDr1e8dyi08GI4MazlYPMCe8eps0p2qg1/vbm6qmt1tmU3TF+B4kLCg1kEjmvL
ipSykCYAZln+Q2UF97qxjCsYz+CfxA0HQtuONrrNDaXRL4hl35GXpAFUiqzQVT/A
awlPHeIyCbYvWVdIvyTwi3x4oNn1mPpiHbanHCwPlUKAwfktl7B4BfJV/mFg6SUD
qNNjXnT/H9QolqYNOQeuS+ri6RLxlXo1TAJTtyZcIfw4VSXz33gutZE9vaO/oPVW
8SrQfwnh64bk4JAMkWJqXrLEq3XpPwwaA+9aGZ1BVhmFLuC0FOdGUcurRamrbZPi
fdXVkFeFRpWxiQeIdZfnvwjYyuPQdL6LRVQ1KZ5qqGvmxYLqlomwZCJwW5MaKWEK
bM9yfa98wxLFsFKLgKv/0iLs8JtybbXRrIdaKGE3HD6KvsXVydcvqxG17MvGXiKA
3BqY+CGrPc8pZnFEMuNCXmm18pn1onALKPy6wndi3wWkUVI8foTAWt02xUmfNSKN
cJKB8gL3gKkTMsVsQ5hBcsU0fP4ajeGm3yI76GhekKHLT8SrqAppgcG3j5/o/g2w
BSQ930cQKzlJ7p3P/hXiYeVG6nQXVxMVFSON0ttM7nHrWrTefQjIm4icO4f6fibE
nXd/bmoq0Vn4o01bQ2ER+SxaJ3biH0FbdhkWC9+mT87vY2XdyyjWQlwoO6R2/+CP
ifh4mrMPH8TUkWDJR9GR7ZYNRADI9rrO2Wvn709N02nNjO0I29M6hafHfZ16imi8
ochfMalrVlSpryBtFs1P2SQ2Zsc+PLHvppl5s7BkKYqnYepgRJ4h2vkOGgDL1s66
vMljxRJww59tEyLHb6PLLEDijFbkUfCmqVw6Cod/zulcaNoB2TVpue7oePOV9+J5
HUtZwFuKI6dorUR49VVbu681q083REcRDAkvs44O5lHqQ1X6cNOe0IGHMfBAYQn+
3x+50cOEvPHOpGyZyXqWn58OfeUy1BGVDFBfE/SASniAuYApR+AhcZuYO+K0pMYI
WAdCLgdDmUxS2AmdC5tXBiQUZ5NZMSzNsZcOesnLXwyQIgeABKsnCO4+TRYKTxDN
sEPTBdwd7SMonSEDr+S+0dJqtgvXOGDSUyYilnF7Py1+jJycvsAeNjJStUeh721b
kT6MV4uBpo9NbDXWUOGjNC98fazouwOEWp5U+8zIzPj5jvxC/IF79qgOXM0SRmsF
E2Pm5EodGI/opzcLzumNWuLwepbvqkvX2Jb1EXHMRfg7RJM815HOEME3q4dEMrdh
Btvtf3u0LCf71z6nX0aEgIdaeN0p/mmYG88GM3Sa3TDHz4/ZPhqzKAyYAHm4Ryp4
loQKPCsdaO5UCT2FB0jNtegVQvJCjwt2EHUoTrGGOULMdMiFvt6r13YQ1P5nZELX
sn9FlRLCrgY6N7KMGUYAkdjHW4YSKi/YM4TVeWhrt3QEjjBqWT4+GUNMh1YXjphL
jQ2/D4PDMXo6PzAyZxgEcsOoTArxFNyLwj95iFochCztH8yzSYkbGfo2lfZtdc7D
dLJbjglz61xV2N5DUgyQLQzXdjrhVtgAfkJ81nfM3j8Qfxa5Bxzigj+dJdZxe6cD
8jKcB0iLG2S95v7XTG4cacv0lv1cnLMZ5nStZ/Fxp8cSz2EU5c8UAnhFNTIKysMS
/7rC5KAWPLHmrA8MbB4vNUaMvUnElKfWyBHDba2CnBCwYgr+JSU/6lWpOAt/QbwU
18HwM553VffGmM7iuL+N3MhjupuPXaqU2hN42U/EF6iG7Lt9x2DYu3sL+IsrgFXO
7fj/zK4HAMQxsAtzsr/rch0HP+HM8cgwYrUFIrg6+WYlI/8GiQEtU+1m0jJ6VKTP
gWb1eolz9yPBTSKP5XsIL/ugvBsxKKA+sTnwtwAPCidLt7D6sjJQqKkKhhr2jxnL
A2jRveFXkJgynoVzrYsaUqs8zfb6HAOPlewbNb+7tsxVR8lKBbCDiPLEskxg5dHT
qcW9jedNrLNkyoUUp4C/zNQ3mNxeGe+6HQ8oWX19XsHZc4wcMigFqpfWgFaZW2Bq
7HVVuRQR/jNS9TyaaleZsxuxPF7++U0UHkRQIWhO/J2VsKq66l5KIvejnoF7casX
kKV4DSl7uY8AjuNWMr7DSe5c3pgnn6nQuYzwDJ6Z3NOmCLzEmTyfQdiRmQyxzGhY
jWHFYkeCgY3iIdJ0hubsAxyoMG4uPwR3sUMXicTnynMGioEYNk/6DEOj86GHUHkP
2v8tup0g/ptcFWdIDJd12UzMcWUwLRyWAFghLYW09O5aQmYHf/nyqyUbrJRgmzBk
q/tB3ifn3SHzUs+7wbG7DPT0QRRGwszq8mC2gr8VSTEnDCnVtWtaSLsxIPCQKbqC
MoRT942w2o8AeJnNojfZXD6dLrJfc2FJ26uftwhkVzaTGHzAHRjWF0ddkxOwDN4E
/DvLoSaOOiv5q/y/zHWjZft7RcuiCCJo2mb+jPah5H0HTpBOVgvXvoxTQcyn37Bb
unF2Acfd1fZK1qIcLK5Lak1yr6HqvPzPd+zm1LXIA1o9B6qeEtNHCFwIJI9yDq8R
GL9ybZFV1LGg5TFlIprfOxFZC90bBOcgOLWnQFhpGy9IoQCEHLHBev5GQ9nPBox9
S2ex+u9x6zdwVuuFfcGl/51MnTsbQIi8hJ0Dz35bl5+3fZdEEbrbsIuFficN0rnK
Dk44+e5PAoqL0S+3GhlW0J3Q+nFORDQHULv4d2FL0y0jfcHzaEUaVkHCECSlmfZ2
A+j1d90JfAJayNMwViQg0Cuhj9OXMjHrdAHbY4kJdLcFtmR8QJNvNJTKxBi+/le4
3+ExBltq1Vb/q9bUwTFr/P47aQJr3ns9msS6tkl5AnKOZsw4UP7oohJHnbZ58glf
nEkiA54jSEA88WYU91y6U83/UVQp8TM7sjGhMOnolpXNZ4Hh4MHOcfJm9S8K0UsH
zy+WmvF+uem3F6J2K7IcZGLX6ESkoNclpEmuL1z8kXdji1Y2bmK79myNlVRajreF
hrAA9mbSdDgIaZMxRBNzvSSFIg7olKpZqOo3dHcSi3gG98q46ODecXigZ5Oi8FGI
FwYvPOvWouELnz0AhWllV/1zCVWN/iXfgoCRi83YJ9KoqOz2aVbB3bIymD+91pw6
TV469tSrjAVq0x+qxdY5X0lWTe8BPfsiWB7Hga4NVuVo24yXCE+ERcC6yeuYb/ET
1WAjW6l7lnxHwmVw0F/bP2ZVdAKcbNutBFPFVa5ofRhNu8qV1vr+SBC1DyRbAkuD
p9sedHc9z/XVTa40bpvNmJ0UffqjalUpDkPUukM1B060TWBz6HyxrjNph5wqyQdy
ADKUFICd8P8140MgOaDlxGSEENT1rfGl0n/WD7IOmEmLUYYsZysSszZIfalYMYBN
OG/2TMX0LBtEyozwDequU5na1UkoyyAQKrTBkBz8HBT9UdK4Wmoi+RyRC7OYLiG+
4gCxvEDF9wtx3+9MNRS3Bb+XM+RpHSy+pchAXEQJgGoriEsRxdU/D7uRejlzWiVY
DCUpnD6BUDSn0Y8LzzXDvYxjSfrJplQ22QDC0WIwK4RPcFf71qVRu4f1u5d5tpfn
tKqUhQsANT56m7zyzvo4u2dm5APL9EVCT7CQnFV/ZuG1//nqiNDRnTD4wG+jH6xG
TV3Dh1/tROPf65Qs2MC+okONicxKaBdfRRlKy3KUnGxxbVfmkXvroDi4talG27jk
zsej5zNHDsQDnjo7bO8oTGZCnhWIcRsYP3Z3vp/R6e6ZLJcmEuNHY1727WxwxtMs
9wdBDTw7nWMmZyaxFJa1bWKGjVzeZLGIogYYVOcNXYNwe/Yt9NlwW0q2StwQizHc
dIrF2MP92UySWKNSJaJWO/4OTc/5cf7ZoIgoBp7Fkus2+B4Q3FvTzNAeXIP2SHoZ
iUFR+NY2UwhgNM5euXnQnuwOxj3U71L82ovhcZ+h1jyJo+vmOjG5QuDGl0sGngD7
g6lrpSP1LT1QBU6ONwrtS0fQ3eKVG3hqzrsTV7T6OU01zjdRrEY3M72WOum/imnP
ycEvT1q6NxLt3ZFA7LW5uQ+eVOz3bhuMJ3uNDaKndA5Ksg2wlppvc762jKYm6Ftk
2ztf5TyqGcL/JfuSps+y0zqz4ePaPdqz1dTu8UIcn8wh5SzURmG2bTnBhwVMVjS4
xXGeRJTfguHE345gSRYxTS4i6vuT5J4POPmHsa3QbFchb3pU2vIhTCO3sAAVhJiv
xwZ5yhKPlEh4CC+yOXG3B9NhK0aEBn67gDz0nSKqz1j9hJ9PHRp0DewS6n8oC7rn
pMbm3hPcsVRObT8ThrYwUod7YXURxuvZpWCUUTLt2RmshG3WznTgkN2/Fc45n/QN
o/M+2Ir0cYLdj1uReQBDtFckVy+JwNeNmi6AUjLxINDGHZaA/7G7UIPkvZGkrasP
QaKCNs4/W3nUlxWQOsaMhSWLoGRbrrW2KHGlJ0Tq5nvc6gfhIBAV894bx8ucA7ca
M0JIW24JU/c6AA+Spk9awwpKkWcJLTGz+Ely68oOXLhk1vPf85G4FTS86WnOvFzE
eUCuUrtD36OVA1JQPj0N2WV7wvnyqdTCQp7jyNEsOdkKLR250fGRKC78aUUki6Y/
Qv+Ho5aH4NTaEcW5KuF8NYjqXu4gFdbmdWX85CCoMq8DFfUNpyItSMJpJz2fU+0H
jm/mdCIjZjacgBsOFkGiBfL5G4rrg0w6EA0HGosniKCwijMGxNdRdm7qD/oubmPn
wkJabC+8ePREHA3HBwJXIquH38m17QD9Np6h82+cM1cWUF6fV1T1D2n4rBiYRpo0
tvSo8TPHbsCtAVYhJliCu3qI+KKmJ0Fiqd+JWvH3je52wgjpTG8A6DRqPg/sNeSo
ZlW+Hbe6eT7H91XNca/Sm4kep/T2dAcdHyfbMFXP4N93IIwMokko7u9mxEjyGibx
fP5npgupfVOO2U0frz5SFIJnfO6vGe/iLTRTAifaLL90z2PdS58SPVTIasCbYpod
R1BydiYeIPjKLTuFRKonrseje5w3ZPZmCutY0qqXE26pMdN+3HssBQ1tR1ruRNyW
HaMaVVv2BlUQ3Sbz5J+uQWip0AsmMFPfNNUluWIphXqqG9vAPtyn3jSxERUQbgGr
DHn9HwYkV008fhmMVbHwJZlxMZ53yAJvY10kUc6r6DUUKnzEdz9fOuUp/OYcU5Tg
DoWW5fCkXfGM5xrsN4tWDHulVYctffIHrAYVr6e0f49b74iSA4hkkG6a/+fUXNqp
RQfJXdre9a2778r536N8R1OxN6SMCevM5UX5845VLxfoyF+oC826zG7tzjRNjASb
GxUgEANs69gB6CT0wDanWX5M3QSDcbdWekECEZaxex1c4hk6V/jUe1dnht1LCpMV
QhWu+39F7mAdZ/lyZhfl/xxvhHERI9jNo+PVCklkTL5vRnspfCuEi8WSsaiMx0HX
GoaF3mHc7uwIoi2OuWAwt5hmCW2QEB7xBX+q+qrbq9Q5eiplfb4RQtwjzRkTgZHE
u7t09kSGkkhnWX5XMGpmL/nM0QTItLxoLJv8t9ldm1wntOYzR3LxjHhu0vcBF+MH
1ot69/PuBhQVkWXfnuzSEyhyf6IcHcFycgrva6VUdjNk5B9TPvjHYY/uL0/sycfL
7DhpT6nYuKkyHbh8Lgirdn4ZJTVUkwoywQTOKnX4LkdbSbUr3607o8MMiCfNEVsR
fJ4u8iw1ap/O26PpeBQiracmUcSssevt2k+8gwZj9iYbgb2Zz7mKUncF7SDtxNQ9
1B9aVo8yLXJhu4vCSEjXn+vmWLybkOD3YTtBNYxOv6FFyTi32Wx7nMtjAOolvPOF
54H5a2AxNZZN4OT0Yx4mJVMzfLZwrk53LNMpxrShKSXJfUResMnlpUMf0Q2ZInqT
HDOjI5yrCF2Pr7aEY3/OEtnNrD2dbF9vC8g3iBlW6OChnonvHxyPchzhYwnfBEy6
8eJ7HDDp3I7ahN7nPJadVF+G2sF3NM5DoFWhq1QVJUnIHb/L3rcPYE03PP8aZlVj
4nVhATUvMfLQDe1oUupOFsQjQa4qE/OOovsOvRwziqYsem2YbebVCvdTFcPAf1K5
lEeSQx9R/2ts+9fOrEBvqgQID7bqjHsJgktty/mZ6SCpqNjQqPEfomM5IcljB1JR
k4zSrJcjh5Sf6JXWnAYx677eeOtVcMj4AcQSTys7wEDZ78DLzJBUHGwutbangN8W
VUEs8hpxsGfMSRDXrO/Z6+C40IPW/93XxJOuuVge/8SwDFDGkth+mkZ7im/Q9zNp
FjdeaDBrs5M2jJQrR3B1DujmlE7K6zCMcAoCpxwmWZosawH1otlybWbhKkdgbbDT
tBNoOGyamjiCKoxxW4aqsIkxbQSWedn5O1t3dIG0KT+vZxm+qeT/86NjTKunwYVC
tAMxvj3j8wW0DtzkGCtofJWuW47eHzxq/g54lJOJEW6eXgYs9B1U1AXrKp8cINiq
PClcdsiUIBRfAoLNs70mQpE7Z/JJxjcwGwF5ToS9IZv4maUvk1ueuHEHMlJ2BQbl
suIAi8d0rKvhK2dTK14kHyLnk9XLbWq/3f07vjUKOpjhFy6Qj8LZ2mW4QxDYNGii
YMM38PdeuqplV9qZJ2fYN96d1jNwLBlV0r3Zfxf9q6lf0AjdxrWsO2dcu5RHEu54
bS3NmIJr+LfhIgYVKIv9aR7ADphU+MRjuA3JNGa7hYTqfdG74RRbR/buRel+OmES
OzdmT9y5qM21e+2N4BIHHb9/D8+q6q/gB1xqVeOZB348vYE7nGJ1HxGPhUZWpETQ
zpQXxL/7g6y/gG8E2528na5kehiVVKsM2LYsEoB0udGIrtp+lPji+qvKeJ63Dq65
KJUUyl+sExRZZDgR4Tl9EmE0nGoyXp6SIbO32U+fvXJomo/54nyGHAjbhNi+TXPc
xn2P+eg3bb0nCcQ4cd/eJhVw+EP6yPkN5SM9LKFl09PrOH1U63CFUVbpOfHIH4Y/
P2GJIClOKbRAn+k6+puS1FNv1wSrlY7CNa73z4aYIXWUgoTXST64YWPx3kVAn3pP
INsN7kDohZDd+2V6A6ywRF4fOR7i7QPY6NmZDOuZQw6ifDrYC5tuzcuQol8gIZDO
QmWD592Qy3voJ5SErgwNmWrjBL9E9ZI//ha4r5pIQUEhAKF8fRIyAXlswtijivLF
6KbKkufbOLCdFLVnCocPVspqeJ120TrLYbnV2EjyOin6dV1Jmn9p51hF2Eo//Vzb
UhXlBydu9VhWzzDLX3u1JqjSXBeDBV2I1/O/v57D2Czuhm8gD+65cmUSDPI2AQBI
GDNqoWNFAV7IAsHujQQleI3m4VxjHvuhaef4KiMGiSNh/lFghYjtN7xFTgfceQZz
saLI/S0fWJJ6V9rTcvHWeYLWOceWFTlQ5B5+OkWlafn+RoCQK5Qitu4qNh5dsIcV
sw9C0RoYzqZyWzYqJvtWBpRa72Bad+s5MgN0Yd0ZXBobcTN6fGmLmmQqbTcFPB+X
+UIY+PIaXIneL1HK1wDsW0674mmUenGJUzRLIAQdAsoH4KkcfQm6z3qB3x9gBz8w
xGgLEpZBQS6xCNfIcaNsVXte3P4ra/YqRvLM5WLp/Mu7Wm/AwYqc8iKaycme8e3N
Xk58JepR+qLZ/mC/mkhtzTmQgu9OzCZexe6GChAjDNoz9ikOfqzUxHCzwTuK0SLk
Wext15ID17rGXScxAF29YNl2uHXi1sulV0bT/BtFLRi5jkZctr2K2i6z8raiU0n7
Y7vGAEktwvcvRMYlT21Np4xaPL5Ho9vVss7k8TY+SIYM53gb3ULzC7GCl2j3wlTi
fzFz8G6UI6/XAljC8j7AVACSh+SP1LrM90tc+uXlbdWNCffSESFuTJfsxidT57w5
68gOphpngo8MDVgX3L0wqnZoVU1xptEG9A/sO9zs2mb74WALX1zf6LEF5akkeits
G1ILH3wnSicKQz5yRYRHVxT4IoQPmNn75RF+MFRgMgYzlyktAL7cSDpKwlqyJ9Wh
iCmpY510uIq8b4I/niLVAINruXgr/ge+6UDckv+yxGXShzhDAg/azOlqrOVnMo3D
lzlNhwxUl4bU/xEy4zWPj9u5I3CTHRSvFJ0mehMk0nTwsRIQhzLbfxyGt7XhhqBq
F3tZ9Tz25awBTJXBhuNhMxs/CX/lHyUeBDDoI+0yFclLfpJj7qeodHFgLFi3H0c8
keAU6+5eIgBKexKWjNVYLG6G/jVdisogfRh7gUC4FH8ggjTroifrc0gye2L6LKbR
LByyt29X0lkd6u9eqxlLijXc2D3q642Wciuey0C7jtfKbVkfaJUFqiaC7i3FJcOA
kc/UQNqN/g1Cz0W4BSuKZ7euW1mW2hbVwEz6Y+Idy4E7w8XnN64MyR8OmY5OisoC
DzULeyY0fZqxdB89VYwfyFKe5b4uQZzNfc7KTEGSefcJ7XKKs7Dre/KFSEXNZWrX
Qh6Drquc+5WT9h6HB2CnleR+qaWcBxkyrBVrCH55JoJdguaUW5Db0BMNj208cyg6
VcN7FFkK13z2UwRVS9PyXlTBMkVMoiYczA+j5aMzRYCe/azQl3YAnCZyQTAWSwcj
alpgA0gAZsnvGfmWbcLxTquA3+AZr9DolLYggoq+ba+g8iVS5qqCTwujvVod4D3H
CQs38jPgZ5ekyNGwQ8TdSd3rPzPoT9sFjtrrGoJRY6wfo4evbSbU9KDbvVYl1box
xIZxJG0LXYV834oCg+8IFBZINbphweNzKnDpCw5AFfMYuh2jEllqWN1yDAcSy9Yx
BdZjQzTxBjmV++1NQQZC7xuIPPab5M1VArIo6ZwhNQfqe4RBuGFPR7v1Inen4XDl
kBOpgBBJ1PUv8MHJHZ8h+3OJvcs/U/QreNHEoBu+/CTmT4K5jarP1xN9aeJMlZvS
ILa2Dx2cfSKzbMlyK2ry8+Lvq3qa/fQ29e18EeCm4S107jPr3tqm5yRbZ/Sj1/XP
fb3ZVnaWZ6eOQ4XuyP7YBPR96lyFEORyaP4tHx37TrCYZc/yLriOxezor4ooG41A
9+lhJpfEvDWSZqPVnqgCPofTSzzNsdnT1IF9wNbMrb+obi7+kX/9JjMmcA0SwBX7
U6Ytat5CDO5TSr0IqHODjE8O5Ziq+1+tA64m0p2blFf9JJchDqUDmif4EA7wK1/x
qYkt3nxnFBf8/tXGyS9vumUMC4akP6/+DcWDfmgvaQ161tHkxqfcltXQEwwaeGsC
5MSYEzunI+UJc3f9o8LfByH1zRgk/N9t7SeMp8oEg3ZGPHp36FP94lPFSkix/1TY
R70kvPv+MtIx4/g8HrZK6QcgRXMlTS+wNzjxsLrbElRhCmftDjfjxCQPCtwXXf6I
uvYiSI1lsal7Y3XrbhKdJARw6lr4DBbyrrvqdoWUxbVwMzjHIr1RVi20IohJHgH0
iOdGoelTfgb/Ho3qKEMJJrANpkplA1SpGv/qvXE/+BNGsbMy0nHWdcwlPEWq2i9s
rLIi9wZxbAqsENVBidpHHuEhbPiONS2PXDujd7/+yK3x/yqoYxPx3eIWJ1Rg1w02
xbGwbdpFu9hOP1SGb6SleJT28Yme98FP4o63nQAKfcCL4ax1zELR3XMAw1Bkw3R5
vzveHqAj78vSj4aslBHpuAtEFNFm+uKVNepoNX1czR3PZ9G+0wpgeZnTDjzygGOh
zA1SY/Aetkc7lrkc3mIWlg+h3qpHvIpVS7tR2aU18FibYAtVEEBmebWOE8CMIv5O
3v2UjHsnTIK0yVwNy3fMJ+kJoRJT4Y3T1iG8/HmCvIyTK9CWhcGcOh0znOFa+EbA
NjlTrh/KFeVBviD8/jKc6tLXdi7v33Fq7HrhDw2wZ3dp0BRjF54zpwopZb6A9LSu
Bv3yZCb0NvtulUEuY8yPL330qrG7oMR/krXoICVuqcAY55JMItpXipP7zpkI/d5/
N9zQq8jDH5HYOEkr6WVDwd77U1cDyfCbuNSiPxNc21iT/xUm5VRE7VKeiimV4szJ
E+mVD5s8nmmKQHiBqHNePRqbE6wS7vnboh9o7k90YXz+E+OjEEpGrDHdcwFaYe4t
3qBLgFgHqEU9wOBoEJVFgJcS163HXOCXdt3+qOHu5jR2iShnXJEpVXk4Dyh13v80
ML0q1PBVQyi5O5LtnnZ8c43lZxb8cMU1sJGEZXBvByC/hmfyPWAmnvsAv6Sfznua
XrC/dMPM1wt8XnUJ4konHTAurCDUrVGdlREG6e3m63Be2PTeaw6KFSNF/xqEuMnt
TkAcygvMeqPaBCh4XmREvihXKBWwhsKJmh10HgBf0o2+P3Gs93H+Hd2Rn8vom9H+
nlY7TH8wgthtaoJngtwnqZtB5Yg5y0dt+N2ePCschzHB+1gJKFxOAo+f74EFogae
Dy+iHixfPSaKk2qR1eTaUHmy/sfBn/T7c2qcUd2pLpg2UW38b4z6fPqBl86d4yFX
VDN0LVwEs8c/As6EqvRRmrtIMLniTJZ8maOssrIOHwpVzoV1E1gex4UJ1AR2HaIx
ZUCj2S8jj4vPzB5/tSDKJG7f+bYXAZTJTpGs/fdzcySGXeqm3W370j81RcLg5zuH
5Xc5uO4w8SZYWmrSB1aUQle61lbdr8LlJKv2iOE6147FsXAYI/tbH4EAVTS2B92b
2zyIclWtFmghN+EtepzZjl/Mxe+3IFA0at+iWXAyH6K0GnuZDy69gbvxmVc07sFK
mQJpo+roN99XrB+jROhVSeai2wkYMhhhaGRV+XaJvv+pAFfVW0zaIDt8yKuN3uq6
TMeZEteXfrln8kAYNNLXm3sJHnQi4DHuUscvd4I+KRsVhtRUrRYbfgTZZn7jAHIl
bNy7zk7vPjFwvSovIJ/B+l6a9HxNzcuOClBMe15TmuxqiDQ10mXV8U48VcENAGDH
RmI84Kyrxg/m1VPcDMTs6Kn4si0TNGiiJ/p6KUcTOICN4X+ubyIGEYjRtEES2+NL
0OX1lLizfRYPNM06QbGQfTDr/UYS3frXMkqMZyVPgJO/4/L+wxIy29cSC+FMPESb
uL/VxuGeqYvsI53RoAA4TwCcs409LFqoZlwkvWVOquPfp/ng22OBPdK3iUgwWFpd
heJgkjKgbhp132huPI0wy/0F8tdLCPfiggq8AMAzuwKjvKPvvl3DprBFZYqTfrKw
ZlcsLs1Wp0kVkW+YUmerS6ETnZRl2bU7csKwJWuuR+ZhAahgH91SocOEsgEt2tZW
Qudff74gTotDpdhUbNbLp1qJy9vWU5N0F/tVrweg2kSXoYoU6Nsqupixs86QQrfR
u6eLBsiNvXx+tnrdFlCxjKiVA0MU4rJR0EDorv673mZOqq+tZDGMTFwj0wZwUJBs
7BJjOXtyEp3eZuEo28s5f1yN8BCBLYqMiBZlT1D3hweaUC7aGtJQoNmvA1c3frHT
g75AwvKNyrSfbLRvBySaPZr+up9aHdUnm+xIuUNOmt4mrXrJ/C/9jQaRYesSTcMP
GE5AkEsgbrCJKeVKR5RI8ccUTFQ3YJ0CeI3CP/IBsfkcVt3/P0oQFXtQTANFLmDT
nywRPvhfaSaBD9PzTeTLSp7RSxpyjY5fHT6V6Mgli/EYEZ+2KfcLR3O3Sb9poZX8
5d4hq4EEWcXDZcRqO9Onk9OfmeaBLpEBghgmV2gu7xVmztCxYQWY/wGw42BuK0Bx
5+mbON3PoANt2aE+vuvHTaKmF2DpolZa/+lRAeeTDQBx73JHItydzSLKCAsTDBjk
dOMZpqzXYXNMNI+lB6abdtmaUp+pYGvP6DeScOlDB+MUWVtWMD/aK+Z+26JwXml4
Jv0CIdk8+6KyUNs185kF85dCElfEXSvaPB5YOP7HcBk7uVGgKcrry+F+/zMswzih
uUQqFuZIo1eLMpiBEu/GKC9h+HWbqnxq7iYkpMbKgnFWCpQRzwLqyZReGJCt7hHa
sFIw9V9YpqP/Nr6UWfnBvp1ZmBVL8xc2mCbIcY/a6ffNnwawyOr17OPPD3Oh6LuN
M5A9amXgtCyzU97tNqIKhedVWiltKFn5NFX5ct0mYMxlvBBMRQ5x37OgaN0bemBd
219XM7t+QEH3fqCOzuEKq9q4lmZkr1ZchTafejLRFI5yEDEvAFZpf1uVKUA+BBXj
OMhzGox/LH2xZGC2JxTzMQwvnWCWjP1QxNPV4pYmvYheOCL3rLg9Wt+yBdx3Ydez
5NEimRFJ7XVrhKxswooT9cHxJspZ9smHUDjVSmyuIdlfBnuq/PyPj0YVJ1mi1TOS
UyYLkwFKEuR+tFQpS3+HtWZzGVPihwj2X0uVFeGkRHdjUzQ+RocRfQ0ujNmxMTGF
gBIa4QcdfNmkv1y/GFQ4DtEms7h1K2zdE1l9bIAgcBOu/SnMv6Rl6IuGxbs5ylVi
bUSAhd5+suBk8S5bwSiFSpNw+50oFdU58B1DszDxxRf+WyZ6ZNXpBCPFNtC06Rt0
GL3SNo0GBtU4zYwtM3FDgE2j6+u60ij+B6Rc8tXyO0PtJjSTXDgGUhAaQkJpDFaN
bNDNyTeoTkIZaHdyRwps36919W2ovU+Ba6vtN7DdboFCWgVL4ZhtvAhg/82suokn
dUBx6EfV+XuHk826Jk974iZhsCmNKG8iIGOM2gFsKo5G9Z5Hvm4+W5Log1I3Q91L
dTM+Uq/PBS20RDSmXG3Rm3bY39Z9dL3In0XDk+0hIpey+CLbNrcfxIiFstbOO9Kk
pQjBimZMGHgEpawKq5D1nVSIr5ozraM1kV023KQcv5Qerp1YoPxTwItrWWwc5B3s
uw6+y24Ml1iDeFj/mVKK/lyXFQN8KntzmZVX0jFVUe83TKePHdrTW9sEiGLWnQIu
+UL4blMvRCCm5MWjSeL6RnuSWJy0XbypqHK8OHV+ExyTIvoPnrXnQSqL0rxMfpQz
yyWsL3Ll1hyv3JAWktYagQPLA/dr129vo6O4woA83R1AXuR2bAHxcphcg8WHFGah
`pragma protect end_protected
