-- megafunction wizard: %ALTIOBUF%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altiobuf_in 

-- ============================================================
-- File Name: psl_vgpi.vhd
-- Megafunction Name(s):
-- 			altiobuf_in
--
-- Simulation Library Files(s):
-- 			stratixv
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.0 Build 156 04/24/2013 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altiobuf_in CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix V" ENABLE_BUS_HOLD="FALSE" NUMBER_OF_CHANNELS=10 USE_DIFFERENTIAL_MODE="FALSE" USE_DYNAMIC_TERMINATION_CONTROL="FALSE" datain dataout
--VERSION_BEGIN 13.0 cbx_altiobuf_in 2013:04:24:18:05:29:SJ cbx_mgl 2013:04:24:18:40:34:SJ cbx_stratixiii 2013:04:24:18:05:30:SJ cbx_stratixv 2013:04:24:18:05:30:SJ  VERSION_END

 LIBRARY stratixv;
 USE stratixv.all;

--synthesis_resources = stratixv_io_ibuf 10 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  psl_vgpi_iobuf_in_h3i IS 
	 PORT 
	 ( 
		 datain	:	IN  STD_LOGIC_VECTOR (9 DOWNTO 0);
		 dataout	:	OUT  STD_LOGIC_VECTOR (9 DOWNTO 0)
	 ); 
 END psl_vgpi_iobuf_in_h3i;

 ARCHITECTURE RTL OF psl_vgpi_iobuf_in_h3i IS

	 SIGNAL  wire_ibufa_i	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_ibufa_o	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 COMPONENT  stratixv_io_ibuf
	 GENERIC 
	 (
		bus_hold	:	STRING := "false";
		differential_mode	:	STRING := "false";
		simulate_z_as	:	STRING := "z";
		lpm_type	:	STRING := "stratixv_io_ibuf"
	 );
	 PORT
	 ( 
		dynamicterminationcontrol	:	IN STD_LOGIC := '0';
		i	:	IN STD_LOGIC := '0';
		ibar	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	dataout <= wire_ibufa_o;
	wire_ibufa_i <= datain;
	loop0 : FOR i IN 0 TO 9 GENERATE 
	  ibufa :  stratixv_io_ibuf
	  GENERIC MAP (
		bus_hold => "false",
		differential_mode => "false"
	  )
	  PORT MAP ( 
		i => wire_ibufa_i(i),
		o => wire_ibufa_o(i)
	  );
	END GENERATE loop0;

 END RTL; --psl_vgpi_iobuf_in_h3i
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY psl_vgpi IS
	PORT
	(
		datain		: IN STD_LOGIC_VECTOR (9 DOWNTO 0);
		dataout		: OUT STD_LOGIC_VECTOR (9 DOWNTO 0)
	);
END psl_vgpi;


ARCHITECTURE RTL OF psl_vgpi IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (9 DOWNTO 0);



	COMPONENT psl_vgpi_iobuf_in_h3i
	PORT (
			datain	: IN STD_LOGIC_VECTOR (9 DOWNTO 0);
			dataout	: OUT STD_LOGIC_VECTOR (9 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	dataout    <= sub_wire0(9 DOWNTO 0);

	psl_vgpi_iobuf_in_h3i_component : psl_vgpi_iobuf_in_h3i
	PORT MAP (
		datain => datain,
		dataout => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix V"
-- Retrieval info: CONSTANT: enable_bus_hold STRING "FALSE"
-- Retrieval info: CONSTANT: number_of_channels NUMERIC "10"
-- Retrieval info: CONSTANT: use_differential_mode STRING "FALSE"
-- Retrieval info: CONSTANT: use_dynamic_termination_control STRING "FALSE"
-- Retrieval info: USED_PORT: datain 0 0 10 0 INPUT NODEFVAL "datain[9..0]"
-- Retrieval info: USED_PORT: dataout 0 0 10 0 OUTPUT NODEFVAL "dataout[9..0]"
-- Retrieval info: CONNECT: @datain 0 0 10 0 datain 0 0 10 0
-- Retrieval info: CONNECT: dataout 0 0 10 0 @dataout 0 0 10 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL psl_vgpi.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL psl_vgpi.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL psl_vgpi.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL psl_vgpi.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL psl_vgpi_inst.vhd TRUE
-- Retrieval info: LIB_FILE: stratixv
