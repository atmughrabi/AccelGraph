��/  �h�s���G�dU<�PK?*�E����rgJ�Db5�y�`���n��p����/��#'�i�F��X���#�u��,,��'n��'�����Dn);nK7'rmGB�}@3Zb{����◀�F~}����&�jx����
n���~d�{m�Xr�u���S���Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9��@���krG��0q����=����U	���\�_$dC�U&-�a1�3#���1\Ez8h�,�'a����i�W+�瑷H������ɧ�R,U�$���A��m�C�-#��ƒ2�r��I}�&B�
ئ���[���>���T/�:�!����R-����:xw�(�Wɯ�|+���p��L@�ly�Bg߾$y�d��"q�B6��H*hnT��(2�'6��GG�W�tإ�A������� �Hgw���X�x�g�s���8�РH��eA�u澿����_]q�e�3B~��O"�i�ޘu���
��Ђ���Z�[Wְ�̇6�(V7�G�q�]�?`3Z�%4��� �A1+u�_*�����C.)#��Ə��+G�|��2�d�GệY�Ҝ�ww�h+��q���蒵���d�k���g
�7� ��1����f,=�������=��x���^�AGf�j�k�-P����L���
#{y?=��,]��d��.W�Uhg�
~p��;�G~�x,�7KԬ�^5� �32C������ӣm5�*o�¾;j��ve�ޡ46�H�hm)��p����r�3��<t�$,��zQ�-��]uZ��o��7ƫV1#��e$A L��^o��t'�P���&�Ak7ݧO���ᾣ���ܪo��[�����D�g�_STY�A�.���2�HgJm$�=�;�����M���/�e=N]�=D�Yv��tC@1�rn�����D0�JaC�OL��ZT
\��^�l~�R��F�/�f뿇�5t�R��"�^����~$��u�}�KŐy'��8��1H��@#���)��&:9w\�Y�Ί'���F{�w�}��a5)��X��L,��̭��g�A>�U��7H$eLCFu䱕�[�{�sg�(6:gU�i�5�炒��Ŵ�(���@��e�6!��3C�^���'�g��K�	/�w��xRYW�j�P:�D�v��V�B[c3��,���y�G4�vu�fx.�mq�_�p�&U�B�֐�֨ēsPB<m���Λ����OV�!��l�D
xPC"����=�����W��o�eW�u�}\E���*\3NP�@af#S#I$ӎ�ρ�A