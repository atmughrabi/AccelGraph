// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:30 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
afq6KSvEn0+nDWkLYplqWAL6b0tCNx0vbdtbYvMXVGSavGDU1+LSwI4VQOvLDm8o
+8aw5cQFamdSatN2E1J3OkiGtbLL/BUMJJlGeuy0awG6mRENhVDN/qlETq3AaQWm
8FaQcsJ2YfDHj/PdAITNzA3fVZOOfdcKmxwtk2vYzno=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46160)
AQHiF8GukCpeaF6iFNjsWNKEJmZfZluQj2qHmYbvIgASHZny26V/Q3LO1Cg+UdQS
C3OH+IENt+7qMmSs1UVy2O2YgFZ9bQGxUV96RMYdEEUBaSUi8T5vMUKrEQtRP/Al
sl2U3SjLNeRfHc57y/Uku2DMkKU52c2Lgr+m1ROS0hg8yTQgUW0OSZ7P/q63LqDp
NlrksGU5JrxFswqiA5iX1bgc09nPZwgH2VIP5o6kr28Gl8mUrf9CXzjknD05DiqY
TlayocF7PJCcJf45t6K0te0o70CTO+/q0LvEZMiK0iGtTosrHH4zzEbug1QEdEHC
T3MnhDTSnceprUzKqJEKS6gc1kQlMXf18IepEv1faJE0QpC4QBkvBtnLGk4wiIr3
Hlyvq7Wuyf2UNOdyAYB45rBvnEyMJ/0qU7CUj4xKwu10dDxQln24Xvx+HO3V5ljY
QBbUbNC+4AAlSO+XdD8GaEVvd2l50o3L9/6DZj5L52++N4y8pXg3sxsNU96P8gGY
IaJaIbqa1comOcemMzhA7Y2dV5eY2414q1t3JZ36IZqDzB6sqPNIjZ3ZUJG4I5Cg
0M7/WHI6v4A4pl6+zQ+u0QEQCqixkRRjO6WjbBehcU81W4oHwn115GHdczXcKyBt
kkwB4cRnj2Vr0ZZ+XXpHWpxz605LKslimQvq4NPf/7UBGw1x1QJKj1DeW9cvgx0T
1Oxtf6JmqG/9CDYpmBNIYG99wWIOSaHqh0MytHrhpMUM9acX3V9ciy3laVH71pxI
OWd37OKV15upGSCvxS16phQcL5eypQs80Ig5Sn1bOx0bAqUDrYjt1v+hKm9NyPzL
nTsLXzuepNRf+RnKp8fdpLGJPnCqYO3k+SH773ml+V30nGis9ZntfAw0vbyC8TOM
BUylZKrs23yVyBdaztTQ6bcpZo6eA8JGMp9wupQizyOCJafqdLO3KglnO5YVOU2Z
tlL2KopsHdiiEiUdWrvG6D4edzNbLgc53K+MVlcaqogo/CHKXyUNb/qf/IMPlfQP
Q+rQIOdDt6HazyrQORE6KZ9Dxsqeqw/Sly8OWym+s+FTLfGT9O+TDMyUyYmiLNHK
THKGxtV5Ji2HQaWxYupQAS4Erf3xbv34ztE7FSxRYcZeFqn4ZENLnbUmTpwgC3Ld
BaO0Bm6FKqFwuEHNKdLTLe3sWmxVOTCObsX1wME55MGRMb0q/dCUr+AFDNdwLmKS
QVRx2VlYnAe6j0s3Yl29d7a25dU+P/Amiu+bmbZmMIpe5EOfhBeVGu7hkZzqAt65
u/PlvRN/kbd4OFvUhhKkEiXOMzIgtK4MumiOHm7wfOu/LUxbdH45P2rnWH0EpByx
cZu1gy9YjVJZGi4p7nHJVq1sPMnPiBVrnrJnAxcDV84erUgbtT09a7F9nz3WCjen
t+WVRpZGZU9iZllZj6EjRcur6I9IdlGYq34tZWRveGKvXkiTX93EF+zZK50j87gt
ydRw6v+GZiagBHqGGZN2lei2Li09pKkwTpHEDb5p5GRdiZICQXAQnatyyFSI2GNW
moxp6ITRIg4XZri/lqo0nY3epQWp1o/7z4HMTAL5d5S+k2geDqmLJb3QiUIfmWzC
YFcvWayqpC+ssbzy1SjFf11DP5SWFYww2DKnh/FAxC8CK02FKTmggmY0M0oVCTGQ
yRArpAswieA0WIvS3Baoq3VQw3dRclqktEKOJKIKKpJLUGo48U0Ui7EsNDlsTxz9
6YNXSD5INxhYFKEXdWKNK/nLnAYOrjxqJf6pyzUxYl8qARFMYXfwIVJ05uRAxQz9
aUcGncYjZzK2IQ53k7n8oQO4ku5qtivMDTwCuNaMEpFxElpA/ZOXrE6ySsuDbEjp
OgXIfmxce1W9H3bHrEXhBWqOFez+Rr4Z+4SM/3SNIQK2EDw9Aukpmmi4jya9xUfO
P4ct+TBTXM8UYGFIv0k9FYCATYsPrVuuh/ClfqVAjlDQ+mm1fYRZ4eTP9B4XEC29
QMnS8VtaMpBCRzNsTv5ckp63zMWzXW7+/8SxK0KaZy3lfgHOzd5DJpJEqyfbRaKc
nHhYfvEpeGaMD8h75DOQRVZnjGOPnYQLsEuk2D7FUeQy0QB2tQm2/wJRVGxhkVh+
nWf1DEHA/himeFMgnZhms/QuRLenPMC0/hp9XW985psr9wfva+QalbyKli9UkMDQ
6qQjVOGCqgD5/8f98buqKgrgoddGRbXQyqS6tTQw5yfTkObGGSEoRzntvukl739N
6PISOjH6+p3jdcgRv0t22YrF8aY+HhfrIWoIa/XdkHvu6Fobo4ZpEnm5SbF7RCfF
aKHJK2rsAgujPKaSNNbIBnTsNB7Fo3SF3/THwFEwrEYsAsK34qlt8S5I1yX132aP
LuuhLiIUH14VO20oI3hL70tq/0+aiPzFkvCL+Tb5H6Lpt2VmKP4mkEKknKErdtH/
0dzwvEdlyP8nVlBT/s1fkUdqvcj5LH8DSkiy2uLuEizlQARddfkNlV/thKsu5orc
CUCwB+IipoeBV8aAL5j3oOPYWA8DCXyW5f/bSRqDPaAWaZdE1catQlV6sSe1iIfA
ANj7S7fibWesfmFLO7PIYaEU60cX0+1tGBXes0+PmNWQvtgD6S9EYs5G1rNB5D47
1c9Ie5TPrToGeXNTXRUSpiP3OdtBK8KbpKmuXojAZ9uOOQtBtt1s8P3mlKi2F5gC
ztmJ2ugFdY2YKiPG3QPD5HFUm7GSUJgo2mCgcG+aJefSG0DAbIsaOgiWL38DjN2c
nL1ZGXxxJ9a0b/iXjR077T0qnFOFQqNsPCYc3yzM/cs/HVh0kkjTfECN1BCuMbTY
1KrvO4/w9XJMqLYWztRmUYdP5cfg9xZM4t9X7s3sgs5QU7Ua7rpNJL5nyghPwJmf
TJYxxfff13DORBA8b8PM68K7y6RQ+sONQ0KRgHM+3KcNX7d2Z2s5V97zR+jKENCz
ZwS0faYTMS217ms5kZq6x/F8jI8ph8NuOPGEpomMfZ1OJ0T6yCG7ViQAGpoVXOoE
mF1/oivk2OpMs7WTJ3yQNxDzWOuPR6mGanF2tRW3nBaZ9HzibpkF6ex3urpo6z1D
UcL+0eIiaI70LJoXFxvKy8gCmWyEV1lF9czCstptkajV8DjoVyXrbm38h886x7E8
ai/T8+dfWiEynyZNLHvYvOXeLph7qCQpKDxW1iUEr/mcXzQh7qhy3ocB7F1oEQUa
NSq0cCLdhc64DCZ1NH8oFXnwHHqWTxoHU7b3FNQRzhfCVnyulRZ+e52GAEsuDWBK
tdTyChOWTCIFQdkrRUnZUhL5nwO40dW6FfVo4aQF7ZOVJaHOtwm9Y3dNwTelIzqZ
eB9X80WAcJlTRPxdXWmTcpB/vgKckUozh0C/7TZGMczoPZS7YYbi4Kde9xwqdEt4
waHHANdS9yG8anTXfslRpuKAFLv+a+ZYKMlStg7yfe8rYfY6EynDP51TRluD4UjJ
xqkqR8zXHSySt8KBW8C5+5glt54yxWkzkCsJq0gx6QmEYemi8W5TNvIMO+/Dy+1x
upbIdM1/4GJaljOfclxLAhhe0u67qyFz273jkn0dPeEjOtwPe10w/Y672w9eYzvQ
a1dxZ72tBRYiLmaTHFw0q6bNpA52VqZLgJvYRwSgldHtb+uSaYVvYTu87pYzvvCw
Yk3v8vLdBrN65R541EZL3uD/YdRa8gNVojRGd76LOxDFo9esyLNmr+gDdZrWm4q2
EmEMdKgay3/Bg5N7z4cTx/NBc5kpz0o1+RAqRW0RFvM02i1+hvS1jSDunf9cmMFN
lLWSScxTtJxmkfDYcGb/KpykuDzRikBmq3c3MC62Hc/ehLHZUnjMV0VrldU8QaKr
ittRMa5O5zk8SHVQ2LJy/qWJNl7+3KMFo8gZ6x4ZIf4issM8HRaFzPGO/ofUqqGs
YvMHImPGpbm+EFSRHOhh+/D6Fjm50fqOD9/vndnNUixyQ/TQ1qnj/r9RcrzUO4x8
6Is+S7SmjuByoQaS6F0gXvGN5+riZqicsVpsB1BQ/19DzTb0StYUra0HE1yqTc45
3xT5a8vNjIvGsmZgX5cA/uEGkw3ZYbqjNRJ8XeTOB8yW5KjXhPI1/pNyRq8CAVIl
fMZDdGGuYwGauFYyWIPaxx6PJ+VWZxwkhWPRF31QSnNyTIzln1NSmUFeNffJcQe7
OCcq/zERzVDdQ5CATs2cuMuBJz9AraaRS4zQqkx776qz87V94hMEGaYYbBPitW66
s40UuVEpE3hNDwBmmf1C8/E/V21oP2jvTAD55ySSFYMD5/gs6LOfD0V0QRlxg0cq
ezHYC0Z89daODc6A9/AbUf06t9V4iRNcuVO9hBnbtNYPinCvYOj+NMPMWlw8AI17
WCvXpTSfa0TsNQ16yRd7x3ZvWL10Qx/eWagYB6kq14DQBS1HwyJzsthJKlJAsSDT
IQSeoJFi64IFV+L4i4CTRw0vsrOO0DzT6vttEnPXiosx7K5AxN0A0+W5J4oK1pe0
KmMRVzF7+ejBf95zOrpyulR1IptYOo9B73aaXWhYRBXva7wnU6LFTWUUK+aPpMDd
BV2vF3hx/Wdt+4sVOLr9Y3VKRIgsP1OCrvCjOxbIX2MCrmnpYm4mG48IDMn3MXuH
nHHk2sNVgF8D8MY17L50shG8GrJpK+QCRnBA8XPyZ7B6lL4S1yxvKTEbgXbLZyBW
nIr71PpWFkzO3UynXva56kI7h2spH9hbwn0uVPJvDButF+eCb5Rri4aG1k+fDAba
k+F0fZszMzJjnqMvo7YY8Gnf8xDUnCxGDO3m1JFihwB44LJ2i/C45u3Fk2PRwAVo
kRBsplQd1vLfrUuFe3NevQY21CKtXeeCLmEkWMglzQaW5YLIDDCNWSVjRVOSti59
wBOvf4ilkUJV0bE5mF4HRpZQM6TxcPlPlBHfXV/xTrPjMkJk1uum5C8CCRqvSH5g
0YYZQGn0avzLGFro7dPFBIQ3YhPcFadkte2uCso8onK1NgeAhia2aufzyyfquuJF
RGoxArgFnoMbdG+kYEWyXnQjLmoEN3QTCp/NfoylggyNb1hc8hioDdLqWfRXpkzs
8fuxruOdxZHuMzU/uSWQfp0FrHCMShqNa6F9cUTBokYDMnhZBExyh6lNMfK6DsDF
Ueo6MAh6LlkdZf4otiuNZl5ko1yFYf/Ogzyrbt9N8OE/wmd1qWLLUtK/KTq6mINP
iwbiJmzSLo0Ht5JcS0OVl7qSjAsdZGq/vOqhIZZlrcxiHntYtS8qIx7aFAzQk0vE
+E1m8OeQvuG2Y4hlUU+z6fIH2SwhdDtMdeI7XZ1K1S6q06Ulk7pOaJMxRgTtlS8h
dpbSjCC49H2kSgXyWdaPB6SAjAYubiry3A83+BuQzsgsgCxGDEom9qk/ZZlG4r2N
2+YkG2FeGfFob8csCK7lG/32ciIfGTZbhQWewrVOPeojBAW4PCi94VLwvifWNJn9
WoPIDsqDfiXATujAvzg+nEcYXI5R//obcaEcr5+/glb1fAbxSpI0MBn+5aY9X3gQ
5FwrUspXf/whiQi/EyyeX7DOxy3/Zs5k4KsEcdxSAOieEPDcHTcKqPKdrSMtmQuK
+YHi1gXM/GatuPHtxgz6BBWLouDw9GWdZslMRbX5RutA9ydrWsdfu8a6W0pvNsBR
k6R7o7/hNnRSQSWb2Fu+kvNepOqpugdZ2F6/ZXLmQgH5007wrKOuN+qQR9I4IKE4
aFcKXtzwnCeMW2+HxgoltcDaWsnmBb0bCWgWrnmLMeyPZP/tT9fkB+3hKLgrwEku
y8MQ1JosBG179FGa8XaGrFDvpqy1NZMMLQvuNeR/DjWfkDJ/YjtS8pkarEKrJlar
ow5HahEwiPJ53ITlc8XYxNcsJ4hxaUzqpl3uw3ki6yCDnE1FXEGDJnQAvyLGhio0
BZCBZNQUd6l68g97pSmZsVJB/S0smsJ76T6V08qvSP8DAmMVpbpMU7ZLDbTAKTHH
CcDrPEtUIjyMcmEhw2eJngpVEV+/SgXbcAufRtdTTOhGxooDHjxcPiM2RNc4NDQx
cPwxWnYzIw/CaC7+/LJu5UR+ejEL547zI5+YR7bPbMlUhy06NdYwmF1ezCoDuhtj
iBem0TXa9vP+ZxD8Jh8+Cjeqb/QcR+sAjGktFqfdnBlheTMVhj3YVZQM41Y4De48
c1XJCWhOKTelemlERw8w7wIVYOzdzusQjAhHu0R5op7e37rbwutwy4zzPm4Ej6MY
ARKR8HtenGKdGXbDX/3uIXWG3fiJmUPBCmX7kCd3AgxE1SuK7f9SjhxR5Q5QlrL5
tOyNwbXw1fdUNYOdlxOwOqdCelCQcgjEq01vqa+fAtq2ILcZRGv+w5p2vdb3clHu
xDhQ2DejabxPyXLv3OxtGCv9ZXF5npcLYGdlSqeUaPAS4fuKEAJB//grYl72cQKE
cQJvnA3RW0Kad1ijwWXZfa2uWGq0gKw3SUDyswdxWbzpa1Xbua1ZV/T5JMwAqEGY
0MFa7MCJkLP7LDc+VxG9DwXcDwrLyCt9Mmf1fP544lCt2S39iUBs363aVTvEYMyL
qoliK7kkATSRt43WZ3Bj7dGp5lLFI31E1r7lUjIonlZQ0PqvMQuVSNDAEFPV97eu
o4xHaRexJVx0bU8DwCKaG2VcivYq9qJ/BzA0gSDY9XYdgLZ0757uVJWZ3tAvTsfD
WyJNYSorldFEjjzYTD3QVm84lu0u4CIOONGMzBljLGSsy2UQhePpCXZkQVcpZ7rl
rfdxwTZkfRvaygnlS1Uda1KSlYpZ865fbEN09kBhNo5tBj4tCCKdJeUTDyhrTypy
RV7xHsIXbMtYu1+bXIzZcfZcX+w0b1lTCMuA0hlAm2pYwUlhclSBwo7LVFa5Knpt
6ljyhMENvE3FmDsREWoOTEkS39YjDNGHx6cqba6ExeQpAva7zh44+FoNH7MtAPo0
qirs5NnSIWI48JiUY2dD0ZnxDppYH7jwQnm3OHW6fD7WzzKXO/O24gN8jcHydj6p
pyv7J2jxikFso3MiaUx1jKonJT5u+ABoA0WbM+eBTSnyzXT0DVuECOjt0/Kn99Ps
o6QBGs6byEjt7bRC8XZhzGBGfkCwE4//dHfkXZIOfXde9CLnBbY7G2rfrrniV+lo
Hph4kiftItiU4lsnAGciaNR5+H2851xtVP837Ecs88SNPiAVzrqVXOhqMNiWzvAU
5wi+hl7NBr1YUksYIZHpy4HOb/A57q9PEYM4kiRQgoqNX3Kr+80LVL3peSy5SWKt
AOmIbBQmtbdXzQmByMXCQzPk+7TjVq9ydveTtPA9arhR+WjIX9+MfrQWmWu9GwZR
UC0nIP9QekBoLqzfRe2txrJM3TnRwjsMfL5517xxxGwQyKXL4EvfeVpctSGFYgZZ
ojHe5klahvt4OOC6s/YHlXtSHMnJBFZN7CNKd4kn4ceYYO6XW+PozHjazE0rmTnq
M0vy1dhlKyWJ00GPXZPryCaqnvVjyqaIOGFy/sPOOWSkvuW43nQYuVzl+ErLq+4r
G7+F1He4cCM5ACp0rolFuU0X/xtqM3AaFYyYORYVNFMTZXVV8hOokvePXz8oWdSh
1p0lXNYHS5DAlTYCAq/0Rn39IHXkdZkf25OP/z9WDCRXYOD37eccFA1FOJ/rCwVd
4Mvm7FgmbUJNveXMqhcKJFbn/T5DzwG/yO56zt3GZYWyNIqn5Sw5Ff2HMpNKVCtC
NgLcJcd1iC85yZyFzlEHaP//rAZ3S/1z6E9ZGHvN1Ea9UxNVshw+cz/qbTTYElhQ
fHW3P6/QKGiE2ZjPGMzGl9cQj1tidBghSCO7828Cl9Fz8WS2N2Pq4EBgLvu9SVIH
guAj6ZifMzseXzfK3W3jiw+xnvx1uWgM01FjuYhh3oTv9bXnQgvNyqdfE+7tSnpd
nS4TBavo0y9ABLAFl1Oquqfy6fxUXdAHRFN4XC9ZhIZTGBgE9xBbM4fHJqMMVGLO
/leNar7kXIcv5d0q9c36NJZoSG1fdt8EnW2Ld7qVHKjM6LADrIsOtna7Q1hT2j0t
5KDYHC+odltExVKZGPok+o6x7M3VwBx78Vt6YrW8lls8wSnLEn5HUVSUCoIuK3zv
bfPjbUPSRZntZB9UotBKdCtSzAEcpwARjrOiOasxQQWXH5qAMdJUSTG2TkJaioUZ
em4M1kKtZ/bb5UNwMr8HQOaUFNyVk6xBaXQPJCnp3DK71z2d169snFniSoz4l+sn
+DHfYDj3V89ahBnc7KIFvarn4HfQLNCmavlsZMBu+dF66riyrdAQv4TzO5tWz5xR
ThWPQWKuQY5JclyVJsK2zkU+IadBrqVtBqMCA3+ksvzFvSRRXKciswDn6bT+fzoT
2Q9R0uHgDUOQ93ZgCaQQGsLTCEIZUM4GVWYdxdfAX7ul4Gn+O2F2n3eEU5SU5pGz
IVIs3sdOG+BBLaoffaM6XRxmWyjj8OTsmQO1J5eJPE8h2VsyvGunaBxk13Z5JXvg
Mt4FWIgD4eWNvPaYI7a7Jr3EPTpy0VDHKoLPJQWp3Ghy3ZBGBtPOQU28A9vs+wit
lXM+E5m4psU5Aj95sreYqv0zgvJyOQm8UHMrBKTCr909ungMXVsL7ak1Jsbde32C
iV6hsUZk4lKv5kb1q9mKRKqwrr/Iw9Djj4qvofKnDdJ/doe830g5LISHJeDF9E3f
BiUdVWsYMQ1UOBLhpf1SKhIV+xbXXYtf8rq/WiHoLLEsAK8ALfpRYstiqwdYjq0+
IMfhN/LYHetAuyP/Qzl4/sQunnCoVVf3XYfRmg6U3BlsHC50F493fG4um65vxDrk
Pd8m3i1znvtQ9w1kFgabcqBJLWF4xnMwFjchRfyLpmFOx6uo5Wyhq62KuqBRJJYL
+2smn+JVIWfExhzHM7GkfOnBCI5hxJxDMoTXP88sRDMIRWzCQ0edQxNKikugGopJ
nsB4KJ+b4u4S9dY6uX8ppAwc8+vLIbHsfPrLB4RmpCAjq8XfUiDrFf0SZfVVpiUa
YNoVoZ4HVCG5sa/lVRVtXcUquU6lncvm/5FQY9rk92pyH1uILtgKJ639G6XWXaoY
7iJvnwyJyUEKweWhSQFp9q52WTAWF0AtUCLwM6gseuswj7L7L19pLEM04zX4zPGn
DfNUQ7zDmkmN6yLbANLeLD9VeeBVGk++JRGJAi7c3ZRMNQFkjvWlo/KpxOiWpzy2
gneRhKWY6AcVfB1dy1dFZUP65aMV7YZJdxfOHZO7jWXGJMiiQMp+nuFWGrBdZiL8
LzQ9mq2aceDGxM03SA8G+xD6x36CVGO5zKR6b6VDUCO4nNN/P84nnHpdFd3vlECO
FAkeIRgbY0PBxbHLtig9asJdSYuO2B7Anpbdkm4iSI1PPz1Ag5kDtSJ9r6xCmL4i
8/UB9UvMGTk/lh9pkNBhnPLnSNCix4eHTTzqQoh6VzP4ZJ3rcS1lhbAeqGXCUlEe
gM5HFU5bIF1aFTlKX2+PsULCgSMHGdgGNUHWSrje3QdUYfStbH0knVNeGpVTbVqH
+C7gt30KRquxAf+NuYpmWzziqlFk0jEpzHcNcTmj5CyeWfJkhBlmgDIUy70pMzP8
LLP8dpoQdmfzRJLSqdgcFFfaIaSygECBGAk/OpgWPFlOURZuWfEsVj9pyb9YdKUJ
lMIjZ/QaSNiuQEzxD9z2Y/6huvBOGo8/DwCit08zvfIoyz922FmgOnWkAzbtmLUN
njJxfnpfu+DWkPMvBxfKzfiCmbw7Jt0aPOdlhLN/Bxjua5rYmDuYPjR2aig75OdR
97xk6CnLTMH0Q2VxHoE7YD4bQybUm6q9X7yzzhnHRDk/EWzyj1YUv8XL3/Zv1FqG
5l3HzkN0KNTRU4SWum4ujknLnZy3dl/u9APPACClcTSGUqoInAQeYmP+17/GT5jd
Wgk+sZH7Te7PxRAEVo98qc9oSsTdpEm7K/m7WdNXKpD/2X72QYpFjEtcMpEBDNG0
qg1iqnrjIkvxS3RB/CcYq7sobMqIITHRihCQZ4ejANfxIaFQc143IqDutL5s2/64
hcWmvCr1E23sMBYS0DVe4ZzwG6yLvVK9ALy6nk4sU7HpD4uk73bJWHCQmDonoSfE
y2BvMk37POS3WFnNACv+qc5R02j9QQR59aUPvUnSdzcXjZ8IFeS/KmS1ABEqofwv
FvOh2p9VmkVqgl7nfX+aqNaDNEo+1LCQX1AOc9fIIa606KWNVbRl2h9RwytlDudS
RJiE6RVyOz3sX4PwB4sYJsyk2DBS71A4W/tedpWaxy5YUv+/aV93V7K0rtU9WgKZ
JWx9Lq2FBFO+dTtgc3OyPK/jT1/AYS+tEf8TSadDOzfaN+y1DXYHla//eXP10n09
wMTXSYaPpAyfWnJ1Qa9ZC3/PIC4BU1WAsRKxlqFyci08GRpYZFyMejTKvq3RyfRr
GJcfQq7i3C4SbHWUiWh68zztdApPgpM3gQHeaAqrQyMajg9c8M5kfz8eHPJuoOgC
KSRv2b+TpHDTNTVEh7SYFGV86vWfEJ7efAFBRC3hvwsjiWDfpMR0+/dBs7DBKQBa
vu5RK7t14zQxHki+4hZcZ1y5X6gCcOUCj0x8ndUSWsWUeTyc4sndzaCez4pkzGum
7Km6qsHedkENujub3oP8v0KQNfYgoTL3oKtRinOzzVbUbsBHZIe2ZN1TN9EpVq2h
IcDfUhPn3W/m3w4Y6aoRpRycHTs74sOWfR6OjSlB4D24fkvstrWnfKyOEXR++kve
Bvj1aXOqAaGDVBXykMsADEjPfuBRMnln73XxSwuaTdIMcIuRMLgGVlFZZNXuKELt
NlhZqhUdfdt7lYLybKie+eFZ+F8dssACvn2TX+WKQDINguW70zAuzSEe2W2jAIJw
R0Je9GbwYhqpM4XQzoFE8+Z6PN5it9nsM7fSImSlbtzHBNXTbHZIdAMi6NqH5p1e
bvVQ5eadZrJT+65plxlel8NNnzyTerJ9dj1bCP89Gc2wt7F10EgC37T2kd/yF45z
6lXCLIbt3xOEeGjdhztIMd49LqMOgaRo+6eXGVXHZ43nK/TFIqeghjM0ESW5wdoY
ep2PUnrnM/mbXrg5DvkKy8OHV73Czssks2/xuvoO7f7V0VB+3QbdzYtyRRAJ+WNH
iFvFn/CmK1bpVQ58B2Buwr499VwWK7fhi5q0v3aw/8Ar2QgkwqJ9XhkwGLttZRXV
m9S/RoOpnS2Ne/Lwunn5bGUg0nDTUtwPg49B7e4eqvdEqQIEvHG6zcZsjF4kLM85
ZubTq/VAMTzUbfpf9AplvlGxhKX8ZWw0cEgGmRgPyWARefSbw+nsoMcFB2IQYVl7
Z3jOT5Yqf6LXiPKGaba6oYUAfeUdnAvjOqZ7VmQStWPqcY0bAHZkCYT0Etql+FLq
qqb3EvzrJps5gTVxA+4PshQTR2sRrWXB3S30iZS4H/kb/lALeL/rvc8ucCaycCoj
7Niot7tL7wCbeGfRRjn1j7mVOD6f9rBlodT9Ycfnd5IygGLFUN3wJBUyLecliEWi
oGIWQgbzFa9TYOKpHx1OQUILtmPiXYH6ggyVhrledwobi/xmoEL702bJ723wqzCn
YHb70m7on8IQM9azDAo7sLHvN7gLxEj/6/iFYkfDeNUj41WSoBYc0jp0mxxD5qRu
euJjfVGD4iHA5dqU7B8iZFI6XeGytxChSZnoSnXjGZmN8lTTpR4JE20Sw+80Elom
Lhy10q/9+THPF43Kv+McjEnp+20ULKCaeTZTA5ithBQPbI5qJYW9cLrP3Lvq9n99
icmCgZp7W23c6lEDrzm3pflMIkv41umiZrF8xTCuhjm5RPBW/Y+rGkgom+AYtA/D
GFdzU4huFIDHU5dwlzmt1sgwodyDbpIkrJH3JwONuMDTBObB4y6rUxTC7E7PURTV
ZP661xWZNpmbON7rTO0vS1oDqlfrYnWUIADDpm6EF3jw4/oGsME2KVwgpve2zlrB
P6tGDT7SHh0KBW6SFHXUOIgIgVhWW2xKPTHB2JVFw9okaodwT1I3IFTwW0hO6cLD
u0BnEHR9zCIkUSEpjIvL1aKdnO3/0Iq+4CxrCUWOq8SvNk42X3eQ+xDKkasiB+WH
W0ecbCAhKckOvfEL21ii0MnLygELiMztsGmS1btfHqnUw1WtSRdVreG7VZFnVPaF
KmL48MU4aztGFVaOrYO/MXGYV0OYBvBftgGgJrik57jahAB9k1pV+il5ICFepuLS
A5AsA22TRWxzgFmL73Z20bF7NN+BxjSknqlHOaKhUJ/blm3eHAoM9Y8CrkOCYhPC
8cDQ3R2qu9B/ijVtFX8eVVRxS02+FScvYDmEdELx7mUZbWey/rxwnHxCI8fngE1Y
ZqspkmOCQmiygtCqRtz1YBSt/FDBbQfNXlS+lDMNp81Dl9TBranypkFtO2I63icb
m4CpPQo789Ny0yP4MZG+YPsa0Vs9C0UiBttRfrUPfna9JZxRJ9F6ugtp6/bEReXx
lxEgMVvib5mVKjLqVg1K+JJq+880hpwTXjtnCGH/AQrtc3bpNDew6EiniYfKeFaV
HRC3AwT1rmuoaEqYcEwubqL3R7ZVshUj2CpVCUJASjStS3bIChgtRd2DB9ORrdV7
d1iE+K3sIcfsJXu5E3XhTUUmj1BavDo1+MWnrswL5h5GtnySxs9FBidxaSpsZrFh
viAEEWvhfwlPsGC/CL/qQ7woIw96oTLpZ+Ba7/jc9GN64w2NW4v6QWMmAoM3hrKU
k4Zh7Ynvj5PDUhpvPSJTcSWEJ3Q1J1eKx/gMLkBvDQDPvk3pB9kp4tR9dIpm40CV
ZTTWzFK/KTrA1fAgt8afrVt5BN6nk91gi1Z8FvlhXUff5NfTvdC9jMv6TFxWfxf9
oKXNHFwTNKsXdLYEqEIphkE8yhAIrDWOExzw0THW8VyATYpMBHLa73OdFtfCeFwV
blD02JfO3MnDK9Ns3nv6MDwtE7bexZ1Wy9iNtHBpnMuqUE0XZGo15yEpZNRayOvJ
VOTsBWOw7aWW45rPTnne/L7xIBpWnaCxA8PfqRx1GzrX+tXvyhwcg61FUnlgPb+A
PQv2ymfbqRatCJHKDpJg+qPhyqkbxmavGjFumNbWnGRCgb6129nA5vY1TzR53zFQ
yG7/R1W4uC+RUyQ2AtCAZEp3gBQmrEJGnLXtmte7vR0xslFitFES1OzOvUpMghXd
8vN50HuMi2zcFKN1so2j4KEUQG1ufwXP95nKjpE7QoKndGVyYPYYB5qKt3gqnFHD
eDinYJi9rBsplrRw7GmqzvNLSZOocPek9nIhamX74TXG0ofF5Rn8AAFUrgmG5PK+
Uc4PGx6dbbGZzY+sDPLdlUUTttFJHi7uCIxVISLIBTaGleqfcCLvcklM727sxFct
cDnqYvhnj1vi/uc+rwk23g71dFOW8+x+Hqz+/CXR2YSN7qhYTZDv5L7fvQAPtHOe
r/SLmOl50bGynwUpFHffkyCsn35PeHbW76ztYtqFc1FoRUd0pC4xnl0kF4CZDyUr
bAs4057St0kCEN0xgDMKhWwkMWhF8f6tZaPo6Tkc5NnHSnYph0h1zy3d+oya8Y9B
kbiZtUi5jCzY5aJnYxpasTvzPi5HjyGFF+rFColCaIRtvtpYgjrvp4a9Qqqr7006
yTTTUksbyt6xPb+VkeXXj3sqbAB0c65X1qUoaJVMipb5qkScc8t9ONUfkESS3sVd
hbRWuNWwI7E/faJk5CyasHQyiSpnPIQQ7v7A9ADdZHWaJEemDOdnQgfyTiDUs0s0
EJPlnacyzH8eONNvdVJK0Fvf7kcALlrvIkjOX3XwgjZR3o2J3xkmhY2g5mOlB/mE
flnF7sL1mqxPMLydt2uWfhxNl1rebKY66WtTTOBlc0C43k6GNPcFKmWk4V87QktW
v5X6FS+73DIGvqmYlgFfaZmWQhJQRBKhgsBZwQyAAexIjufld/9Zvcu7tGT0I6yi
IO5MpB3F4zO+HXkkCp79aCgoPWVgl7rtgdcewOtlzWKCZGz/l8Tsl0CpjLCgmkuL
8/ALT9ATGAjb3OAt+D40KipRGeVDabQ3CxR5mrU8SaEAk1C33pp0s47nhHcwENxm
2X7801H+y0JsNVJIT6PobxjlbB9yuUoSK67CJEDeg5ncOJkSLTNqnMSXIOo8jsZO
6vQ7KNb28/0pR2V7IIPQ9vRa/Ru4wpFHzjsp6PQUg5CIC5PBmqvx/A3lz6wsJTzI
WYbeUNXwgouQIQxh1wGdcXqRxAhkhfCedgJhS2gFx5luKrn5bwGCI+SIpWmjFW17
psJmhssU4gnTwTwgs6l9aSM3hq/b9RfgX8Xaw+ZUbCklBB8eaG3HkDaxgzZqIb2Y
e8QbaLgNJT4pbuAP/chark36ItownVxUrION/ZuA2pIgT8OUDJY0Bq0LilbIc5kJ
+GL808zu+7fdS9256Yl8OB12rP0VExPnLxgRh/mcaVHVEU6q6jAEi3Svg8mxYirA
ZVMDwMVhXUJTPAATpv+XnmGYIa0PRkuU6SMrroRo43ybOVsuDFAp91klvnEiYlYn
YPvADZTSswjAKETJeWXzkSmQGdImFzv5M4D/ilZGmjteAq+B6t/j0/16oFAS5Lz9
dQDJB+M786XWKGmullfqzxkbMyfo08pdv/cgjuIoNYT+pdlGORLxG/dQZx5/EDMp
E6w5E4GF76oC/83Y/5HaqPjDn3nrrblwzrEUydrYRQ5xHazys9PRllUk+JKhLORi
0Pf/jVYmbR5EUeWMpzcBkHKayBXPxkvVSykT4f5LvcXiqjhrZRl8Kkg0cZVDz7ul
bilF98T0/LNL59I5zCh2Ayt3Hw8qdbeUdNIe7oL7q1jkWBgcxwebzONmIJQseBCg
SBw+fed+7TiBOhcxX0GnHyqR69Xhmcm4shG4wPzDTsKmuWLWlXMyxNyo6IwXe5fp
pw/7+cBkPrXAVSXxqTV9CBn0xRbP+3iAMVu0OS+bHyTxlwwejZ4HEFTPSgRPSw9F
DOnJ7jlmOCde1hpa85eoqkVqUMUkuUXhLIxq9yekasGfrTnXaNFUN8EgsLJ2mcGW
JCaHoRaZxLIK2fM7qBDQsKjokrV6ix1JTzEr/rqvGcwm7U5Ws+r7QTkjZ7OFg7HU
vmCPOrHmCtupWrbu0kIWTjePdYvT8/aWbSE6lCMQa4Gj5tDQuPYPfMhB7uGAxz1X
XB1Ta1DFCuTMn8KApPAcZN7/kAtVBfGeDd2ER0SsLS/VQtDfgCoixUiHxahs1wE5
JLdFk1Est1j6xFbc0y/Z/l2KrcFEMzZ89muo8yGoYso0SqtcHEWm16RQWD8tiVTu
Vqf85XCOecx42mvjLRuEtR+c53AYi219QoBpEj4CUdX6YE3v5GjpNtZpxsHJW6rF
LlQ/N99+wZTEMUI14bzGt+tt+OurtUmSxDKBkCcZ/v2//MU1lclwTDb2Iknkwaac
F+TdRFEHz5pNnXNijkqpPV25tqdNkx5o8PjhSm2/txWXSMfw6n5SwdE6zWayfb8n
d3a4CNQGLgUvLBm4a5RcNdmb2l2pJllIq6dLb4oet2mwX91EJDccKCZmGM8jqPRj
3E8oxtWsXSE8O5ryVAA81QcO9H/sNNd+wTreP5W5y2J2+iTY1OqG7OHUTo9tlsXq
dTPsq4i55NW7+CNNXj7tiKYMsvSoXw8jZBXPisMOC1EDfkhEjmXcdRmy+ps7JIP3
EcNbnHO1/kMi8q1LrBMKb3/vx60RnDnkNMISAhwz7QWw6CvRzIBwqzk9cj1tkXc7
VbCIM6hSI2ABN1EgUgHf+kuZ0QzDDl6Mpct6A2awyIh0cOHCYH4DbDR0wpk3NNpi
Plp13/4s7RWjQORkGSujImTbA6/r4u2urPtQQOWRUsXxEtHIhoT4sLDveZ1ApsPH
mFLMaHytinj0k9IhK6hm5EtxDsvnk5Cc7fy3MhDplxpwccvY7nlf+mLUNoqbe2iC
fmJlLVcctPRIKiM48VPd6dYLxLKIfCjL9+ikrw9oQNju/sQDl969Xg4W7SenaCEa
ti6g3M8RBnYU//1Yp1V5d5UlbsKreVUg97uuE2I81x8FXN16+py0YiARGok/gIRK
spli62BPO2o9jGf/dnDQo23xX8pb8JknsZZFyc/ct6s286thaq0uxCZiqEikATuA
9QhL9O4vmCEDnT+IQ8T2lQZjL+5m6F4FZEJhpSt4rqHhicx4PAoOU924T65vBv5H
tQGqD1Wc0HTGR8RI6m2RjtcRRfK5iO2D74EK95a/Ozej8P7TpjbnpAp9vX4x5cnk
910IRUPkPOCdIoQnmiZRnlRfjps1OM72FOPiRD3yombqJgG2Ewtlgyn8JvqI7Dvy
MlQieHyw9Li4ExVBDLU7X2YCGVI8xv2b8ikiFd+koji8v9+AMzD2oHgrzLMv+Iop
4C95B76BzKeoY4NIQ6FpOn4p/v3+z0UipEHRT4+svcBfSComJD4wgee3mGSqNPcq
JjrgKNCT7eBqxwcxU50676eOY1gMw+2sGiUmm1VIOe4w9ijPdsvKJz4kcA/ZZpgB
niLHcSG/gsw1qo0Yz6qL+g6/o1PQu46styCHxdd8d7g1Vjd/S5sAVPN2UtvowNN1
oNGk5YXzx8yAkCAC4GhvFS3V6j7Z9HFU8fDXBH9hSJgT6mPZ6jZxgzRK82jrWHhk
8w8127PKT28Mr+fFfFwOG7H0Uzq36cpt/Hgkxs3ZhDbw04ZgXAew0pNZUMlPugG4
1y405IVrQYZvUmuGGHdSqDRSqLhv51sRHquaf4ba859PXqLtT146QeD6wdz4FqvL
c7GqbktN1jXz+FI5P8tx/Lu8evZuQF9mFVDRwBnnsbqxEChQ2CEwwSGKqiYVbH00
U+N49ZXs6aLkWZpUZ3oNOX8aaO2OH87wMHKHOPqlCXkAuipTy34bRUdtrBrMiLYf
N8xqccoONGfmp/ClnLtXeWG0EoT0k+BUOl2ODm3BmbW42AyzWO50Ir7VyWZbLT8y
kv3fEDEApa9sbuj3Rjf2/iQkJ1tCYI1Teu/53rjGUAjvIc2p4e3JWCU8YwtJDyRm
AnesFqNEV2K0bFDksWKWk3rbRWV9jSZJc+mqRyMV1He/15e2wIhyCiMuqPUCx58N
YY1jvWF4aCAX+ugiftcEqH5KZv/HrcGhyecc/AdvscPjCTojKS09d8/gn8udumMU
zabW5ALYgNRD7YlXeUDO36ZcXXnViSzUf/nrqR5ioYfrF1fk+43KtPip46JIWWgq
El8sjFd4GfNhOnMw9KV9v9ipuZFBy1eoH+QgLb0O7ltIimFPpeMCnvSpVU5nIZuF
RUc/Qqe2L7lMeb3YRgIglyPWZkipgNU6/KlC8f5iHvNeZZ1zyhmsMBJufzzfy/6t
TlibLbB17GxEGqTCdmUQdMroaIEp9mBSGLVdlDL9T7dGwDOhjsDUjThGBbk0Rdn5
GSZPNv9qhQeXTbbbXochReBKktWVZIxHu6hlrsr9zqOiJalLSDk24lAL4V0SPa1P
A4hghAoyf0Rzs8FN8H1cUBEtYDfo16RSqM+3wPqkz7Ts04WPlfdD7nVoGyweqkhJ
2V0tztbn34m8RPV5tB5tq21mfZvsa8jiIvU+p6acSzR4K37Am2I13LJ6eGYgU1v2
KMMDCPlYCrRD9iIZLmiLYjOW48oTonhLg7jvInEWCMhQB5qJsI1QIlArrkXf0xHr
pZxRvaImRPuEFt2HfPezXXZw2TN4dNaDjjtiys6QzkDgya7w9AU0y3yKg4n4f/Z2
Au/prp1pz7N5U393XqYrywvG9DJxsGGtKToEgcWzZjcf4Vab2TFYH4zpDsG750FH
o3SS99gXsazOFMdgbvM6DU5Bty6nklTNSt/8doevZTOSoj6keFUbOAduQzzVwSH5
OAK4+iUsVso52CyNvybP0rSZvZ8Arg0kWcp30zHx8oR1W1Uf3E6lvXqDw86Klzyu
VOn4NyZ02FBtRTozOZ2NUQEdpzpfOcC/MgN54LKGpbgkh5zxqFZklRkNXqhXmV5t
gw21pgAkufHQfPSfzjQxFpIoK+CEHSEH5pf7/6OfXbltYSyo4gV/Jy89ulGI6GZ+
N9LPd5V2ixIU8yKycE8tiRu6lCdUCpc305Vl+IZHv9hC/dQ04mBGbsRmzsSSRBIO
ErYxahCGYJg+cO3u71mw4jUdvMywFw/JXpgawIm9nsv8A52bZ3l5QcZth2dS1LSh
4tT6orsredtJDbDKk6DPHPgDDIixGzPU4XuoKneKybUw9KNLIqF93ezjEkPxyqbu
rdGt5AmGfdVyet3RF+knHRugxiNYmBPPeiisTyqP/IWxb1gJxnA+KZ1kTRHKvVRb
ITTazeoh2iqKrtYeCUdT2zwaBH5EJLFSn03sAjGnJm3bLqBPJpAJEGkJcFqOereA
TUY+0fpZnhIINEu4bHKp55Dwtg/zw8AeEJ8Nl6GyR4hK2rRTLIJ3ZKcaMF0vgrq2
h6XgHuMmy7yzGDEgIED5yQdHwSa63eYv17DBEj63HFm5AO8vSpreompoT1owEVtp
v+1aSdHNd3/M95WrqcPYM7oKvSnozfqU8TpMS7clb40PmEEhiEev6jRg1OnL+yvK
y/YAe6CC0N9RPjbJL4BgyGv+qFVq3uq33fkmE+o5AlB0liJbgK2qqU7KX4Wyen5X
pkRifpqEUfC8PPemkDbL7RLeKaFLHAPlHxzQMNFi3EP/shN6U9JfGzDUp/KXoYy4
Myaoqkrp9/sZIRg046cRQEpii9946nv2SMYjBYGCrYYJDc5jY5RnnMFeOFSnLnpX
nb1ywyrUAwoMrSO3VTkqN+zD0WkSbH0jMElXPDXENV8T0mgFbfgu9MHLwDsIXKfi
XpQAi9/KZIPKEAla47n1z+/BIqDrO0gF2tF9PCYMr7sKNXvi9zViQ598LtIitccJ
TMCqUGFZUXX5IeVoR7lXeiaINP52ujG2xy33xncFNius524GhH6JvtSBs1Wfaq32
T1gb6silpiGN3eTi6iAXoX6HzWih5yhrMe6Rg37QG6ncqhppXD7IoMNQUsx3dIlu
bC1afPgk9RNTj2VGJH2K09pPIsov99Zu1i7KKzXxAC5N5KrtO2QGyztl/QlOL0ok
INpJj9lTJe34ocMQ8BIMKL4EE1jyLYxPlL0KrqNUta/64VXqWyoMM0UAdJYbjoSv
2HaWW3mKtmZSCR1LU/j2YPDKPnUWbQ4plpVWjEUjTnpZpUOGQbvpmyvXbFAMFBrm
9ORG+S4bBZ/4VBMupJYr1Ylp2bJ/iDPHRJ65NVbKgGPhfMZ9zE4OsZjVfzDqbvP8
1F3N8Sfv5Sb0zTV9jHV5oFDcI7V0hJjc5DXPVqsPzMF6F1SsT7cJDNdA9T3uh6QM
meO8l3F+64d/PLB6z7McSiYaMXoEFmwov8xcM7hXOJQ8BkeuuoVIF5WPAQ4E/Ds1
/HdZ7dKG6niwOQiZ0/CsbKRXbO6m0KTNX3bn/snGa/tLQGtkb8cAsmjcIBnV4FtK
sSKM9I3D6qhaemD6xydXIyI8d06gSqtCryx2drgvJGQY1dLyYl63QcmkMNRjYXe0
SbR3jmFSksmkuB/r52WRoqcYkecEZUEaDFRrCg+48ZpicFAdMOtMBXX2HemM0JiB
yQTZWm/UeRAmWCSzKZw2fOjwRyzF2UnIGwT0UL3yLhbQISenwLFiBZIgcv6gbpWN
cc5cWh/Jq9bvrvNkZJ0Mp9GlauSMGOQXOCn7I9BuWubyHQnBvvTMnBTi7lL2FAy+
siVwtPhSWjdhJ7OijO6RXy6g+HxNQyrnJkprAoa74x/oaJ23znxW/A5ZeDDwuLkJ
Pg23aiNyPR5NTsfmyr0ff1wYVj3g+lI+5CJPgrMC0UuZYxwDLGFJqYPT5yZY4kML
DkHjd40pglZ5HWHy2wszPbdcNhy98ImWsy6HxltlRhiaAga24OmDOdNXs0tC1il/
mYCqJHQrgKrE6knBW1i3ml9C07Tks03zCWnmL243JH0ftJ1zp0RAJTTa2g6l04Zj
TWhnlAWag4TXSEqO3fWc51HRhabquhNGUlAoJ7sbzqQtfhkAFPGGb1wlyiAVC6SP
+FOn80FkG5W0UUOHj4nUklrUvghh/63Qn9Xpx9UUT3Urx9LDa52dulcyrn7qZvEu
W1w/RMXbAXt0YYaAF0J881jnxWKVJUsIS1wPUsZkLrEZYdLjlHHXePG7jqTWftrH
ASEza0jl7hRtrM6+O1G3/zHl3l1x5qK5QNarGZygsjlU+FBURrHTFqeWRej5tSv4
dE8duwJMt5klXbygAgYUtlzCIDDkAuBzMxv5XXldfWeTmP1mAobGDD5bAC6wZ5fO
bluYT36xm1Vqbxi9ZNf2DcEj5NvmOt+mx0n+/rIVXTdFC5JIngw+/8iNVrLKZc33
TOecwPKTpM+6WSE9kTSZ5SinYYTsGp+vUHfYt8OqCO94QaG4LoGsHexl7pv4OaW7
vm5ba7dON7qMGx0/KP0LHyvcKiPvXQiZOwHxoCPNM0cP/spr2NSHfCJ9EPYmRP7a
SRdNmojTRBqjJSGcDxiWmyR73p2hxU58TJL9bPlW7tB1JPPqpGPURETpWQf8v8S7
O5kFwEnoVIeDb1dcMOaSjwk/CsyorvF6hJzcEi7e197Qn03YVIClfGlS9ZW8oXrX
OHJjpo0j65A4K/4kEj2Di0Y1epTApdialhQegPJ1PV95kAYpjZByE66WGGKQgI7b
EA9Ibq89nQCujZwR6a9pjDEyar06Xl3FnJgi8zxVYA9/8V5zK6klbNsIYzE6xMKO
wo7boa7AvpCGO3h0WS8yaOGga0NtxLFyYAY2AJdPxASDvAZ3p9tMcWn+bUPUDGnn
rMsbxzdG0wcqh3TBFQVnkYdz4ZDRjsv8RlxhRlUjZgkF7sw82FnmsqzMrPChpDTe
5BJQEdMQ2srySQYeL7z2aQC931rUEqZOwgc5Dgj12BilkpkvQ2Uqcc079r3LndCG
lxo2M0lelbucZ/jWbcrtbTZMMv+QY8iwjhpvWvRcXmqcWGrF6iFkBzo4aPp27G1V
j019AFm64fRXYGv92YNdlBlXN9ng8MVFSDlscxqa8WjJykhHWYnfuXrF/uJKiHrn
dmzNlgfuSxJ2a5zsqYcCxVpNlOOaNDQUBXFpKY9Y7SR+yorXmql1yaf5ZFXj0XZa
aOeD7qTHuzx0i467EhGry9Dx1OyBQynM2YJEZ/DljQ1PWOHkVG3kRgiyljbfcJqI
P4CzRUomyApEPC6AqzXC3AWhyu59TjaJFn3bS0D26WGcCt2Zm7vQEC5ssAC5u0gW
Awg0NdGMSa+wsLiLoGVHdLGD+2/knouxNb5uhBI0EwpnXTc1ivWhW1VrsiuT80zz
NSu0sbnHd4LyGI/oOGHWEbnA8BTxhoMdtq7flMvjlyDanpgQjLcAcfSJ8Ya0Tzia
Dha9l9Jn0CbiJ2ZK/VcjjovlzE/v05G47OAhg9JBsDMZ8XuS28pa3IYk6w+pdyar
UO/bf36CU+5wURH5usUts39Zctk4Btvbed9orKxcqodg0OwTlkJxhkPyEQUdhUBx
zkUEbKJiQb+dyHcKsfUl8cYn/T8+d5sY5UFxd5jP1lcN2gxG4cjTipcXKy16yJKz
PfC6j5ozhcFbZalvfVPrhs+443sOnoXPf7F0UjmiBXuX1JwdNPXmxt26hP4kVnq/
Dj5WB/W/Y1TjNxkuW764prZdFN5RzhU53L8eHPwG1HY3QsQdUi9uIlLlq3lCrjkZ
lbLPC/TCOP81sDyFw0o2eo86kCy2Dw6XzHJVK1BrIa2YMvRqFz2Ps3921x+QZUTN
33waIPePAyPXtu6pyP2xY++REnwdQAnATiyDEf1POLBCHUyHTH7HalSi5ofgQGHc
snaGAeMhNSyI7FlbiRsyUsG3HW5dsQ1naNdCuZHBKxUSgkfPf0zh4bg8gFmuiV7O
eHRlcDErBNaKyb6UJggNCcsrfMuViJtnl/NkaDcsxKZYnafxnjHAsXGeps8gDW0I
tuA8Y12xHPjXTs0qDwjoOps7EMR4OsneW7fxHqV7EM1UWom5UZxoTPGNnAiaXALc
0qYUI4tN++U9147Fu6x6atTuTjxdAQpPGAB32CRoJGxXj5ty0QfsRZLbiNwTtKlg
gxrzK64N8XZT/9sy3WEpOf0e4gCYzVbLUWPofvrxQZvvexMGeLoURATLYrkPCaQe
zgQ58bD+sn/+0z+2JwiOGjyXW4o1exqVJo8pb/bjebOyPEQPYrFBSoxJ1Z28X9h+
OCkf3fOHkOTjeAoJEXpAyIgFSe2WKeR1rr0lU7cADrlsopMwZdLZf8M18ouqdKeR
jArLYmH2XtUf6t8blwLoqP/0+cCXJoGsR8p+dt+/uY4fQLoNLZIRq+FDP5FaGCWO
PgTyXGwfKITRnVqkMxaXPVq/vTJaDXE9OIx0Rayz/M9wfY/dMjCoZPZn8fRt9LYD
YV5xBomhBN0VJ31NHTXSQn9usUk4PoGLh4zyOse0z8dhpZZN5C1IOJaJOAB6JEsz
D2g0QtA2erSnCI2xXgLOtT4o8iBMVXNrqAGtkn64gHJt66YQ5lxeCXubzkfxnG6p
ovd9F00G0XLFYeswW8tXsHdJnD3VL8jBGKfwxRYMqOHZSaO/10RvkmL5jVuRPutu
Y7QEE1J0sYhHn5UaZgFqeSGKzAjETshD6CsVSGUiCn4fUhiZiJozsnQ9cdkwpF8V
WO6lWzFCxFr/P6Cdi09k6eWv0PzuswUXnjsvx9Zj8ZwvTbioGkAQQEcBfUK0pZr/
8ONJaAkYDTO+Z1qQ9itEN28ciRbXhq3S0FrOUheH3gDc6n8On1sonuaLsgEdmaHN
KVlfDT6vPY49Ng2Si7dzL+cKll+W4meTVzwp7uZFxGQIfWxwBbYAhZBbOOSicFvA
yXhaLBm/yBZ+IreLeaRn1rkczdE8cJ/IFbNH40fTVe5wWuzt2NindpXr7xJeIquC
Nq3myi+WDlCXatzy6yj6n1QkO36/fcGTr43T77hCsK35XBCxLmWS/+QYpLSFXuhU
Qx7u+worxkQtIUtzt6BsjQ4jIQuyN9bkGalfaWxq1LUZ4+gZP5HsppWv7vdKCX/q
OQp4n8Ti0I9v5M/VqieK3TOUA8rri7PJswaz1IHSR3t+dveZn2wiFvHXFloVfh8m
/h9MtuHLrilTWVdQFVzGIMC1ZVz7TluGbvzQKlSnEJVXFTLqvlNsh7bQr70ijXrR
80b+B4cjw9d2J7wRlepvT0iLUJ1hWaCzmE/L+38LhlQOD7eP/wNm5ban9AUR9pV5
oTx7pqVuYzny9XldoIM3W1ntTkq67/lxOCKhE6rYHfLFPv1gz/0HoGoqliYX/oci
9GqyNJViIFnrXfragU8lkHV1OBswl9bEsMchCx9xMPBmZd8YW31xJupQRotjb29u
PA6HyfCl2+7S3HxxqCI5k/RAaUNgTHwWzChskhmeqgXQTAZBGG5K/yBJvIlxqGZB
XjzkSvDXov13qCSqa5LAcQ/bhWF0xQ6Gfkk4jyQRuUmUjKrBbAHV6cyr8zoTnqA0
BUi1FVvEVLn5o7vOkFfRDfPyGZJCkT+RipKz3lsjFc2wwZ0wdfDJ0n/ife8R+oLo
vbz/VoEBue6VMRod/OH/FgNi9rTbSvFROuoClwzDwaY1Rx2iEFjOILkVjyOjF+Pq
DyTXaOhEZv/G3kNe+GZjHhBMRqzwUBhGvGtZ0ybd/F7q6T1cqC58YoaVdYg3IwXp
VcHBasWHSXiF5tGJ7KaOliSAJR72VFv5mFngyG/pmnW3tzSBpRMLF8E5FllCr/R+
8xWzI7Xu4sHNsSwaCksTEEbmzQmDh4DusC2i0ckE03wksRUfqfZ/6jg7iaFESDVc
2QnokWQhCL93yDs1ZaejLGuiCsh9R9DWSEjCkwHaUF9P8TPA3O19fJAESk0D4L5V
v7BWTEcJKK29xxtRcT/umPXifpYcYrjt2zq6GqNcU3epKtLG4IsflEYWYkZodqIk
RxvQNVPAE13CBbErDMnIAhMAkLsNzMJtL2xekm6tsHoqxFIt2bokL/woVFXNerLN
Otv1iRzPGjRqpAIFhN91tyGSJJx467Geg+VDorM7UZmHjq+uIZiKO1WDyDN+ufm5
8x77CTH9duaMbdI/JcMdBn5X7Fp9/Wun4cE0dzAh1Dzz3MNvRdFO8QdNCk7GJToj
igX5M6EFVJ8/dDsGYuFJWUVAhG7cOr/Q2BOu1/QDaKsvqnvcQJUyUZJ3L5dbukU5
YHvzk37GDiv/Xr6zYbTgSMfBxT8w18UBkXwO489HDplGkUBzr9QReGgGN6ikj3z9
JihWKBIzcZGB3k2ezM0c1n5s36GNHa9FNP+rK7GZaq0FNy6uhUGcOhExSyJsuX06
aKsd+fLWueKTNsMv+OIj3mTsOyMnWecQWVgouofdp/S9UtNwxryKvT39CzWZXwKe
H4hj2ehxnCI4zy0cYJM8BDC4O7nUUfaQmkCZqzxVULn3NhmuSx0NAlEvhfDUMIAv
g7mT6EVxDMKXAGCM4/n6srXfLBlSEY10gqgJS66qACmYwz1BnwULZsRvsAPbxgMT
2gL9PfAeaeCvff+lJZofZ3StKWBhg1TI1vSxxD245BJ+fh9U/T9NgwhHroALaOkf
q+6lA1u1QTcDN1Gt93yyie1gjLQdGbESMui2gQlOUbR4rHYMUF3Pj8D6jbooNO6s
LifWdHMrs4aii1M8KOKnvbToLNEwsYQ91vTfMe8ZSRjbfreTUGPgv0uEQSHVSESH
UF6kI8z2r7KmsJJxQOZnpV6GM984gBpcnqwdb51OuQWY7yr8O6nzUzKuB3T6F5rH
QkZi/FTRjqTAz+Fv+KvWQ4wOoe3GEn2QIoAVn0cHsg6pr1wTkVuRw0IWBTBia7pA
6QknAiUjMDvFX67v9GD0lvqX/GL0yJ+sWOncGZJ1lOdEE+fiz/eQprFUyTX9zKaR
xYqsSaGpiCjZGAC7+hsMeBIUwiQzYfpAqEU/9eK/DoZkH966s+iUc5FZ+9Bif7z2
wgWXrNAm8P/7T0gjMewpJ5su7D2iNqMCpm4cgepXAAsb6BSN2YB3+BQ4BoGLqn4+
lpCjeQDYkJEycAugatGtGJAOr5AA/gcNP9BzwfXdZHRRoG4HG9docXpUF2BmRI9p
sjjE7jZ24+qIBkKzCMjEhxVcVUuiYfku/vHHmnbHTMvjh1GYDXHYlUsz4tH/JPf9
UFufTE21wVLs0RTciMlCtXS6qjmZO14AQ0o95JPpA9LZXg38bkmee3aZJRpQgHaS
MfydCZbw6/GNTzx2YNebS77IWBc6xijY6JAVf8TLFXflH3uJm7qQaxURD9BY2wpg
buaedm0vO/P5xVluZAAOhjM6N7rJSGaf3gKmosQK2gKUILFVinJE5zsig3bmktq+
hT5ZOW+5lfXhPrmW1UzAnW5iIzom73WMjV11W5s/kv09zowFYz/rXwEM3XR5CG9f
RtAwwHNwUt10U3qp1wuBJC7FDWGuweLZNb6MhVC4liyutPZR28CHyoCG+4xWTPuQ
hEaT9IrGjW+artLxFzfncfkF6aC/ssDnKMULI1AtgUtJ8ChlqxOzCnB9S1vKvW3J
QKC+p4b8ujKQK5eU44XRvqMoX5RE6Ulcn8/kSlXWc1vKF8R7wD0ksYPAp3OgOL0H
jeXFmKzjyP4T0qiung7KTB8fy5ByOEA3DxOH5PfV0UJJP4KQFlhYozOpxyaPI9uu
w1ulJHwAX/yOYQLZWbyJHdUZZYz6rxXEvnsr4iWWKQoxLdgXkEZMX5gRTzgFSEfS
qILikmSM5wWjp0PP7W5HdgfasEqdfLZdh3/nQ+txcWR0DwO5HpjrCBLnm7FFYVAt
FNKmbGCZPXUa0WwHbz0bmmm4fwN0A7OLQRwfCU+C+tpqNQ1xzLVt5pPfJQy3QrFG
FeonpLxlUe0HdzTkQmR6TXXRZ2khjKy79V4L/c5eFK0PGN2mRadxMt+Ug8RfvFyx
akgNRDmeU52vSU2ITuTEaPg9UIs8kNffWXHU+JWOuJf3AtsHOraHILt9gRvuDYa5
Ksr0xsiN5hSjLxzr8g04HL29JGdq0D/3FRmM4JBp7GLN39AGsfQI9JYgY30/xw/t
vvDiNQ7tIlpjKi91sFsNjgEMncCm2Frmk9McfSon47R6BDKJvTBSUVEce6hsy7xt
bd05Ktf1ZMxqU8s8fJrIbknWv039NxwmDORCcrPpCt38X2tOAq6fNPDUx2jse5l3
C5R8cIrGQNOMjBNlCgQZQ27E5A31aqlRWPiJibjosP22mxyJek0wRduCmmL3abzB
9BoYu4nTmHks7FWcjVDzI/+NxXLXL/zPKEKAhvWCbRfQxTavePd4TUHkvdQZee9A
uPgoHcxc6PL3UtKFnKVAHTJ4IJLQX9RZ+6diMpN7/Ba6B4QQfoyCy0d3UpGhdJX0
T45jZx+5KbQ9wwvzj8Au0ngMGzo0TG/jxMktZHsDAnJpmqcoqNpomp8s3PC8ovEQ
Gx6Cm97caa6OTRJa8Jc5ZfDg+37bzp3p7/xLTRrcYlwZLXnurKIvBTFY82sYFEdq
JYDfKXePqp3plmmx1yN0tNK4BkdyCWX7INpHJdYZ4Mc/BVKpMU1m2vI9WYzq9wTk
U9fZaUcEfxqTdsi6AocjVWiNM28+3ZaucUZHQkmk/CzTYkL1NZELH9RFgmXyjAZt
OJN4ev7t46bVAtLw/zQKUsME55obqdNvidNkMOi6fvGpOkciDUSrJXNWtdZ5I0aQ
DEeZsVEb6owvPc6cm9TMiOxFNK525a5kPe8oD7OjnChXgYrAHez5r+jbarkrTXnN
+yERJblw0jhcJ7kqodfobCg3u2hLq5eE16x6ss73tIduyqxkI5VwRJj7dBZBolxs
Mo1+/+nKqp9tro4F8klcEZqnLrEI/Blh/8thq+v9DyqMguGt6DlVnH7HTqu876RF
2yibr8ctixhIaf48aPKQeFiVcb51oNDA+E7yonqcHkqs8yWG6G+kBe6dbKy2qVeP
+NybpuRPj5Mc6nPgF94EzdO/ElsKc/R7rVym7MK5R+KUeFhtoxDmugkuklvyycwA
W5bVFy4I90c5X71+f0ZuUFKBqSi2eRjssM12prsguMopHQnxd1STUDND8WmJCvlv
Jzp67slGeGRY2lcJbvtXnJLp8fwo8AhDiSOAVI0iA4XfOovha5tsodS0A+D/o4eF
+tFf0usYtIrYEleJYnToPJ1of6q0kCe8WFMg+Sr0uhyBLdR0cb+AFoGyWFcK0rsi
luzd+VdJNJW1O7OqZbgHRzer0wwdOZlg92ePUN098iuKAQe/h2XmOztokTljQBDJ
h+J5lLU7fOwgaO01U44GYsoKveevBDqyL5I3CkVbRIafEUMqkKoZO+OJLZyzv6g5
BQSj+ry7C84N19tNAxx12YXE0RvXC1ebqGvQIKOwrsd566Wc3o0mYuYtp5jgqeDL
+3uIK1avjq770FMgU9hxXHpPdciLzAtDhcqRpzjNEIytUG618dkIPpGQeFr+epVu
7L/x79DdHSaHd9OBhPYLJSCqzyOBoqQ7j8H4V5sXBiKF+OWlBK0m1HzKnZ5s5tWw
qHubrx/WmsVcj2bVyS0DZIf/Pe9sNOe+g6w1sGMJKqlkGGyANKti5NEIth895T+x
Br94tWEYMQABXBoODYogthjrR67aR55oO8tWuRomZ3iTmt16/Ypx2/dn3MauY9Cb
evgW+3fwCZmy9POOVh/S+VgHSqhB2530fJzvMKtT5FKuYDOsY3EoQByL10p8oRJd
IHFoYfOlDRvs80TWAfNM8qYoFg2mcdsK3HpBxtggqK2jM76mEYnfn3lw19zMlhld
HjzVISy5DCXBcU6BS2VuZujnqfz7+lQcYf4N00VyzKsp8VDqJM8EqAhhunlqP8N6
EaEf8w4UpYTVGzdbGpu9ZCa9t4zYAEna5T1hOK7C6Y74/PWh6ahjU2k8iOVGRM9+
SpHhMnf6Z4WIimZ2C4e42hcaSeMUt7tYTUvxNBKWpC/9aGnl01HFzdrHPLpqIg+g
HyTM4LrbzhuEqWUkvLI0iHn4NO5S+5c07HvwJPn5sMtelGYqmc0whqRfcVeZ2Zk4
C594u9A2Ikn1X9GA4+RGPOUG5bIrqqh7/PjWzWet3/JHjj7qO3M2o9jCt2i5KdBt
p2X4cnDIlsxuqvXwfLRS/g63N8mMBC3lsVZu2iFc+lPiv2v4OOu+sQtjR/ZO7zon
2laZLRO8JmAhhtP0eYrq6+iMAAkbHGAnkuA3E844AxMntMCTW3ondR2V/JdShD/Q
x+QBRbcJVUi4PIaOlpkwqUMKJUvl4+AmZm3LJH542VF9eiOEFRN6a5GWCrrBuw+l
GKZhSpFLxYyeREaFb+3y6SGwVySpdlVUWViXf5iOKhOvPyRUlgZCGRs/pZlGrqgm
MPmF9m8L+ULIrKVebQ1ym8qzMbeplzpv91eiHeX+K80/DYnfyrQLf5vSPu3wWR2Z
oktJyXPUbHEa7NjvUKmcfozlnL4JHB5M/p1jRKPsGmA1rrPZpaVp8kVOmvDHc4ok
NZeoaia02NdCj8nt6Q+t0ke3k0J1C4HKMmwzIlRYV5lqA+L4UGvsiNR3GRn56gYn
L6siMQb3Eol4Y65j6qJnc4dVZIiOs1uCUybEn67HVMy/+Q4houweSKIdZJKWip10
Yk15i3YjZ8+U9+5Ob1OsO+Tju6AoYZWw6nftoTSCT3pXblXXUnOK1F9j2aM9oBh+
rbVUvhPNMGzjMC4CfaR9TFENMocMkaWG5+dGiqRgPDYQ+6XzTvgiBeNwfedJjkCR
iWGRsRvIhocfXcnWREMfknSNT2Vq5JwfCCc4+xasoUMaOafc6DGBm+DQZOUzA43g
VC8f0hyqKwvGw/wHaoJSiEUZvJ9hpo7cfrn2TitDIWZ8b9GEZDnPxlhm+6R9JLyo
ovnlULRXFoosxW66TPWqv8JhUDEiWA1Jp+tMoV9L8nyOhMuGZHmA30mv0UtpjOWr
3aAFBRyPHM8DMP6GlY7y5Ruzkpa3/drtqcvpDXTZ/idHmZKVC+VOyqoC5piovbdi
u+oQTet29PDaeroFo9eErLYAJOpGTrBJfRqY5MHUnVftPqXO2CICqxoFagb5eEwD
hMlOc0e+iVbNLPivJDVkwlT3zr8vweY2qOWhKp2Qm3brKxs9iuwdEbUzE+c5VC8w
6OPkHK549O0cPFxbbblC3YYl+pPrZpiA7cgv09wcZpVhq1ral0Xui2lsYAib4gJy
vxU/sWererUguCRUzVEMHIqx17fC8sHInoE026YiNYDhmtlxcMQPpVT/FE9EdOCl
hduQpKsqqGJtzGR8y2LPcVA5gtmEcpu1K/GHN83ttLN4ICqZWory287IdrmXjeX9
x5ybQvfVXOQpbq4sYf67v8gCNVAqMk0jA+uIJ0Rweta+1DG4STiNspZjZhx56jxZ
oDKpuPbdqwk9EFMNIcd1mWhkwzJ5ZY8fcgJJXy49docneufBbaeNeUqrb9wuAJsu
Eu/OpUjWHeaOA7ir0q+il1KokrO9vFX9PwbqPlunBFShC+4SFcGkQ7CpX5jqj6QH
Udj3HzlHRkVhzgXNkDHcLQr+fuzmPY8Go/r9S067EAafYnIIzT/PfPwqdbiGZRdm
B7a+CTvYviF88VpqBTkD1pDdriE8LMVFeCugqtW1oslIc1BlfMI4hlzEndZj528+
Gl9RoG55ePu0AxHWQCp+105UK3mOVv8ioI1zkjCFvz4Dbo7NI6XNLrs1btIE+ncK
orkgduVh3NBt32TRnCs1sKAD+YVm3V/6wMoeePp0JELFzMiXfGcVK+XDi6ASD3ku
01kQsE/ePZW7UmRvg/XM6Zg8bxDk3H6Dn3G2NhFUhK/HBgxT92H39gGs+PPttXj6
nombbEYqXV3UBh3a5TIpCgP/nqSD9eopXV47SY8Aut1SiZK4XHc9xaZukBgN03iI
+2OodyEWj0J0msB7mn5OEJjY2CpGDAgMMp7N9aFUcchNHx4gvma2awqYiuXT81vi
smoQd+j9d/SqiIpORxKT7r737uBxvbNXbd1J2YfSXpK7oJGRPknXOD43jp/oPzI1
kJHM/pm4bMD1CxiYazOPcJBSM2dGVGVH1rjHsqYiO/+5yGToieM96Pz8tQY1dl+V
J6syImG4dqUkd6QKWuVALMqzXwgrPr5Uui+fygMtl02cxf6reDMsRQlqfxKRPGjv
VIee1kRmSKQ8Tw2SPAGbxoIVl5dSz0evNoaslsIxUnKjyA16uGK0e5yx+hT0/oki
qZd8nlnW0aNGx2PoybwTQQsKZAJBYLp/6hseZHHQeVTD4Ktf3kYiYRuhstqT3Zg/
VYma+jHaYT/PPXn96hLEDEAALmrz9vdZ9fEjQPFNKomODZjh1cXgllYHKZP12x3d
y+ofd/PlyPppEAx5gsQrCMVgY5UcHOszhOJB2MAqWnKtSE8/UflMPgTTbSa0j7Zz
JYZ4XuRyh/sh9TuzquFkLv5qXcGC7LOqFy02ay7p3U/ck+Ossp9SJTIBQTm747Gt
pguQya6OJ5Sx+5W2dzuPJvR8yh5gwYcizWhJK23KI0RFCHg+CxVrk7Sd3PSfj5RK
I9YAT7E+rbBOdVzAqHUwYypS8VERGdpTGfnIII+FsS+CTXC5FLVOv2+qsYpYGnx8
G6iQfqb6jiBTDK4sYANTY0rWWVdDg4w6tp6eaoFFLEZa4tUwB9mZAjMsXdhKkl1y
kzvybt86bK1f44hBOEMI47BV+yMU+0QY7cItTp5NuJRdf1z/s7c+QC8KTllUiIOV
660oQOdENADZlNy0zJKXqVf31/wZfpb9g4at3EftcpsKFlo0ZYK2RK67of3zMiMk
3JqvfvvU72RmaKmS4ilGRncQsj/OIuRc7MbSIX2abFz+C6pzpYy5xB11o+fAwvAu
vBXGPDRqX5uhwJl6Wg9lMyB2P84xnR9Tn24LBVanXnlYH9A5c8GC7+dylwvYJI82
whtUy9YpS1frjXkKbD4OABR/maW06O7HrJu9ja/+eXn3C2EY2WfmewoPdDLJCHil
p27MLMRCllyC91s0KqBZ9/O55Cd7/e001jeXYfv1tTKlJJ2zh7BdFma88W4c6Q5U
RC0MnlPiBAud4gzyAKqoOYxrGxJO0ent9GsZXn+eYuZzK+QlQICJTU20fXpMtqpy
3M/jiukHzXcosynGY5G/LS2h5rYFfdLt5sC3CWs9PLx+5XPnDPI+LXcSXhYzJWlc
pWVg6ttaHzS7YVvdv7Yc5f2iVoYoX8jnaeN7WqRMRTct9IArSH8RTZ9wZ+mJ5Uqo
5plgye4QMaOaHcChH9k/DybppUradx6eY/pTH/VlT6e8doefnEdQEyDzET/2uQYN
XFKKHHt72wrh8CodqmPyZ5w8LVNTv9YqIEyEd0h8kcDhXnF8CE9y/G3jBIfm7qJ4
7LcST+qoHgjj+zdlcUBrUWAQgjab7MXdfFldeUHBV1KwXnQ1q3CUVmy5eCqXwusa
PSfVOJexLpYCc/Qh/PbRhLhQ6d6Ic9gRDdayhxijJUqFa1PY/9L4sTDZxrcR1t81
CymFvA4mENY13c2aoiHy5IG9IOkH/PYGkX8RdvmAaeZxzlzSQN5nyZv5fLro+YlQ
4+2+OVQlp5OZH+Y1etZqzNj6SHsFVICije2SvQFCaVL8I0VLH9wgVafflg7qsPU3
AS777IGeUbdaAr8cXg1TVaQKfd0/9PuFyHDwa7khJELei/6g8HnA3daRfUcYYFP2
IEuU+4bjNqAU4MR2zzFfdQwZmhNVq5GnDkOj+UmXppFgtXlPIBT/u0M8fXDjvE0c
yKyMXHEgxX+DuYimoAAa5OAoHOgsYQfCcTVmzGHclORun8aWeedCH9zQIpJ1QBnq
ILwc9EiaEipWp6SpDiOt4XTqWIDfPwc7o2ixX3R8HbBVCok9pglj5pLI3xjfySKe
EOEUH6wJHuD5eP4J+tXjXWg7MFFgKc7hyryCPpzhTrAnOnSJLC6QwgHkaLx8BiB4
tOceZvq9NhmdSEwsTGHMqASnoBNJY+C0KZ6eHYVtu+wa4Yc7RB8IS5t9gw2qV8s0
CXfC0ejnRAvMQLDxWK1E5qnuYqGoB9pe9WppZ+ISo38ry6bI+7cgHyW7Taln4k+5
0L5+KXyUKGV1RT2o3tH+ShPPYzuZnvqVK/FNz+i3GznK4IW/TTq71nM6fkgUyN+r
E7vMkmzg4xBeQD57hEctEOZzQios85XtDfFQXRjrLhzCs37KqPnQJWYw48FM4o77
NTKuqKCW+vGofvKgJiVA6yM86gMLorshaCFqQBGz9StkihhDsWIx3FKwHduoTUwD
eOEZSVXyZg1e8VFUbQWRR2YJitRf47p7ktP3CqEEJTatdkxHPOjz2CO8Suf92gYl
5VFr27FHO20+R7EMHWeSQ0/E98pRBB6gBz57u6J4eslHx8z7EhNJdH3PcL8QLfms
uP0wqQSGLm0//4ZPeHJcz6T8cPwkLklH1jQla5jb6kCXG1LMIZkqWBF3SmgUBz1F
UPgPKvKVhmqu+H3TDRKIWJncS5KkcOD09FkY0RzIi54LE/oEWu7sTB7cHEEoPqE+
KmOZv2UgRZy49KVlZVXXZSVTlORbWSCZw2mNpZalaUxG4EEIW3x3G46JbNFlAGn2
iq6MAq8WabSX5c7RfNHPKRUGybG4YBsxmJ1d4DyMlZxPmmDtS4Mf+JpmaBrbd1m2
CM5s3Wc6/YLEoB7oAFli0zhufmmNTJZOMjXfSostgyv4yEUcfq79hADu22+HHFEC
cv2Tz7cDiKzl7rByeZby9tSlqTO5NAjYJi6+KDHrZ2yJbLmpui63VvdwK5Zkie2g
deEgA5WKye5tDGq+cm3PCpCrJ5oBoq/pS9zOxXwuyCh324DPE7XzUg+0uZZKIhQE
j/VWuJ5z/WmXZjDUivRr1zhEgghlT/6cVu4/xtlIps5jx1XAaFKgvehlKCMwx9Wd
+QgaHiwOXL0BGEtMkjHwIhyN/kYDxNIcMv9evPwKbvLfDAyAqn+ibcAop1uRhgvo
qMXU1TX54OPPiTSURjzbHngzFPBkoHeX3gtV/ikrhOOTgVoMMrcSurifRZKSDKIy
dRlzi54C0G/z9V56dkFXy2+bEJbjTwgSUfc2qftEGj43W1FKlNfcNWZJVvwUCCUF
o+UCaDHZQfUhm3VGH7GgdE1ayVZPBre6H9hqIQ4iw7cE2QjVwB0P6tE8G/dgbqsP
e1STOAMWW8ZpTDaKW7vx9xTKmnkNayy6K1QS2En4DfvbqtA4wI7p0Hv2yl1xuwh8
wYExbLm2M8+dbPgpMPhtPbEOi4qjuAPY3th5orjKqVmpc2PjeFbO4ysWZPTjGX+v
jV7NkmIk/+N9sz/Z3ebH8fpVsWbJJg/vQIVD1FoLqn1hx6UHpZNqJxuwVVLH3+QC
MUQjLo0LkUmkI3NbpWhjnosxxSlwttInyCXLGiZQ6xbgAF//Tuw5CZfP5jRfk93M
dsXjQyz6Xaaq+LJDtvIy7nf75/FThsUinndNx4e18R3CLoU5zqIGaDUV+wCMIrVr
b17fbbgsv7JfcGWEXYn+g4E2jWtiDkaPHMzXSpO7QztRAb7ZdMGkFqBvvhIhpyL0
2pfmaq73ciq6eFamR4y7Ju/fIEMVP5RCbIwgJ8dop9w5VYOil+4IFdIg1RjB8dIF
xGKbhtuo9qMd9HOtmAGJXSL7762w4drOdWd0CCm40t5ibQtr3AUkGrJDAp4oSB5b
ebl2vTvtniGy5T3Ccjnuvp4atZZbYDfQwDwET9/Flpx3Eef7afNeW2bKqw/ZsSVY
Hwe1jphGKREWSslWrg7Ad2KfJL0OCuxRhPoeCjeHKOnSulquaKpO9saPuvD0dYTS
TRdnzYDEMNUtVQhVfgh9nMXsWbk50Jr+cWEb46ViW1YZXl3DzWw2+xKqdq+9wsLd
w/DjafcCNcuQ4o8UjhxiKecrpPO7GW34ISzWNcAEfFcvNS397Z+L8vIritBPsaYb
DHLEIQ6WGOQbQS8pr9X7wpQ6LoEk/4EeMYrMGtop7efeR/597qt2DiENi05m/y1H
zWqblD3bMJh2V8AQXh0oaepeGBjvAdeypa4BmDBQJpw+5a1z+tVvBhk+U2N4rh0A
IGpnNqP/6nWoeQf70kggGYd6dAnyLbAafuJnCFMHX9ZrUCWCb/T5U03+dgM9H0mT
/JU6Y/vTRkcBdWIOBj70u4t+Ksg/9Vj9uwFVQm0TldqDV1tv8yI6ZJi4H94hfj9Y
g52xQMMOv6K5Vz+izRUj+HI3jXsTQ1IaXfRcBOPSNhDZDHg0o3ATsY3aLzD0X0sn
bK3KaK/MIbIeYc3Li1vEm0hx1q7Y7wxybLjB82d/mjY8VPGpin/DWJvfW2tM/vs2
n8gZG/t2Ip+EzLIVkaUfOjOvwuowlGzuiTL89oEzVAVv/xLVg3jK9QfUDc0fdV+c
MH/OOVFOKo7nRc1AO7X162G44M4XRl9Z0cNLHgBPJAQjIAmgq2PO4tKeg5lVCAta
N3nclYL5yEHuADPfU0NdAAtCC4OHeNP45fM+0K5mdNxHMj6rUtLjOhg2n0pYcfZF
9LcIXr9dzOcvcggGk0BZL7bLs7Y4qUzNNw9ZIMrWZye9KgmokbQ7BiIvPhv3XNzS
FazWHejxcgFju1Bk9O3laV55dKBvjOdJOjaGXdiBF3rblJUl6kw/x7iIqYmtEHPW
d0zlFNpS2DaR8sf2Ezoi1F8qaiv8MmKe4LwmT3PjQgD3Z86iEmSm3U0PHIPOzPj3
nSIXA9ZJHCmnUMrUTtVVYblMb1i2Gv3zuPk6JYAwGB7isWUNtP4NGMcY3cUpmaWC
GmQpm+37JpuKBnr59locmP78sMy+5cKH/pNHHGMeci/59yW+tnQNqLccBvwrZLPB
5BLHq19FZW8btEvuKdu2aqh72cJAdDUY4ZpYqKrDDXJCwV5ihCZ+xwGyi9O1qI3s
nfDXfoLTxua8FdRN23ILjSKgnVXoEkTWbNoREaxcOOJODYNnagPxuh1Jct2w4e71
iChX3cxOtADLANZV0BLB5L60yIJm6MzH/EenUv01+HoCs8WL1Q/hDNP0r3hB7kbe
Pc8r4WX0PsufjFcevF9bvct6WUVtBxSkD5O3mmKOSlSFjyAHuw9NOozwe8vZrNDW
8NlMF4msGkEWTX+HFQy2rwq+8EFRwcdrlYyFxiWBCBc3w+hpZk1sLHsJ/88vFE3J
BISOvJme+ZuwgYeWDm6IfzSPOEnCdozvfMJsIpo0VEBFEaIFq7r3Bktk9Ukdi6Z0
66zXgEbnb2bLqxA+/OdulJM9iAx5OQEkaiJwUtW7e2ZR5Eqa+EqcHAA5JVN7Uhqj
SrzrdUrCbpwp1xwD5Skx64Mr4v6nwGtvCYB75NPlIwdLurCFrPFD0N02TlF/Fnfz
Y5P+2r/9kjCuMFSDnfGt723/cN5k8uh3AmdeMzH4oaFM7LqsCCy5mlN9Mul2+MFm
pcG/ZFX//oZUEDgfb2Ny42t9Hm023D+/ZjR/Ip6DdkgRTVrGr9Pn5cK73JMyiEQQ
gMGDID9ru0I30g8WOUXpPImv2+/tYhbAQ55h5l6oN4P7GotY/lvNLI6EXV06nx5/
zMbrNokjyG7wTsI3CKZUxRMRCP7bHod+FsyB5StetgfWLo4UnQMPVJhyJifdtwPD
lQqdkT8yRBT+KF08j0eSkeqUHSpxkt84k2K605J9Gt3pIUgdZawsgpHPX+YfbzXF
VnLSVgwXPSTcuZoa/Xv86H5TdIt+tpyr8E/uCNUZnng12b9DRATfp5TOp/txIK2V
fuGbd2dbZeR6afKvXZuQwX+7GEJJuyKtPOtxEtSq2R+5Kap84A+96dKP9ne1PSUE
ufvFt0JryNixqNaGXiTTROiolj7BrCDc3n8oKv8KtZPTXD8Zfhvfr8se6dOrqwlX
CNg86kNkrOz/Er/Y0T8IyvByqn9XpwLyGlWCGHujjLGq1jPXYBPc+0xIOPUUQWhx
idwlgxRDj0rsgnMyE6mhtDLAChcnAM9fskOITKIYPx1yXtuuwAwu8CSE27IezYyB
CzoUvEresU89U3QIoB/xQwIWVStpvvVe/ca2zWExF4kChWbFPzqs9LDQAV1e/u3+
v8KESS3Wfkn0ln+q4bR6v/AarqvbxkMNJ+g6WYkq9DKjbLdW/3DC1u7o3pTMZng7
TjsMG51z/CaqxGQWdaEWN758gZW8zOALYP+kUlE9ZK4JRaLDsjo1/6pnfIrTOZF3
gSIt79MAApLk9DwTKuCMN1FOAyp6uobDMVr6eEYDURqrVewzgwVzM32ApZTwo8ov
RhwZ95q0VGX94uStLstxGlo4XpcMPZfzjnuIG4aMqJ3EVzt/QyJByOmnay/7+bTR
YHg9T9fGSRSEi6vM7lldEsTWfw5pbi7rHaOVKf0bs6MZ+XfvSYKvi0HaYDvQfKf6
yHKkFc39MJMnR6OPEEzhqvDx/MEgNHzUXPLkO1wAbm8e4dTH6Wky9bugUEv2ooKr
LbCTzOlG5QxLfZIfRuWvXfPxnNwwCaXIG5oZw8BiS9PJ9tgo38323DIK4F3S/0F3
mXFoPXfl7qKBkxBlN/wkpI+Tyfwk43yCIx9E0fK0u4KcAorwA1Kvo+lu5vwecJST
PytY2Im44bfXsruSw/BxZHEmMGJSpcRWDnldovDxm8Xq8hE/aH/1d16smjurR2id
synaaONPQmJvxqL1lFum5os/pjKWanr3NEUlm9UMwQ8J4+uyyatSKaf4Jd4joTQL
436K+PbFHesXv5rBV/bmKQf/N4SpS6KeKpmymhKUMOffnHZqOeXeGafVU8QXmAeH
171P6H43ureOkOFhJ23BCFWn/v2pIhBIblGtsQmeMXl58zHe+YD+aWHVJ+/EF6En
IsNFT8s5DbICCbnXbbLF4j5bTDBdzuL2dFKOzEtqMVaoC/Mxr3p1W3R0SjC5iLbb
IdEehfQzSrqweraD5dZ3mllu5ldpwzNcWrGa9ExPan2cOGTbXQlLuwHK0Z+bt4Y5
1zMvNFZr4BW1ntoYhCcI4dn0Tv7PsYaa0P8yUM3Jw098PEs8lqyFOmVoX9KMiQlq
9fnr2yH7nx3OuT2AeS0PbXNH8uarrVrkPWgWzyQj6xtPpK5hmoiwGjsbewueQU+Q
f615E5JoEPkJxOCa/MiA0dXj/fGvDDRO6FSx0PSIEvG14tIqSL51evOnkp2EUlfc
7QyTcfjObVXLEcn2frQK4DYFAXV2BO1MIkAh4UqKhAXuMVhfVtzgaSM4j+TvDPPz
J9tC1nEFSUHo/9ZENF7pmPvTyrjpJDG87UY/bRR4YPNNFmFs8GeLNj7DEmbWVJpo
0Q4q1yY+n5SlHK3PtjXgpgUBYRjDekHtK2iAn/saEUJAlwO9bmxaSw5niNUtZ6OX
wZ4c98V+yHSR1jLMH9llMMcXXr3KEKQTRi4zvuyaUj68p7ktVaWlNzvBTs2P+H1Z
xttvEQqALOX7aVsI/wRkp9ovidzWSxWu6ijlflALNKM8Phq+s0aQUC8heft8Zk5U
Fq4QVVb6xjDfx+Mc3q2eMfSNkgVXNn/bYnvvpTWynrCZu11ofhudVVb7M2qR0XGG
DeEDz+5U2LoZqHw5HyvEwBrz6/KVV/vcESUC5mnHGLdQayvv1oMaspnabyTiftKG
du+6XjRYmhhVoXBU7vXsisnLRyA7XZFpEMLck1fcoWCyBdcJ6JyfTX2cEGYXmISF
HVhJyQTwwmImEzqDZbp4RszK/sogPOQufV007x/HwjBJiCgpqclB5Kk4YVKFDEfs
S1Nvkgr8tRh4XTbz3a59JthkU1DomjbWHmNJhG2EMnXpm3EAGIOIkoEr2WHFenh3
x6mHdkGckOwnYF+KZq/uC9F/pwiQPC2YXczRgzp7D+rmEGKU7Nm9jjHrkqzkKPEO
pST2wI9sVCAuiFyi30rlsCnUupS05Yh4f4q+XZ1rlyhAPZVrc+WZXjncPrnjqoTN
6eX9c2/Wq8ax1mDJN5lt38JY2dw7MFaBXuFtwuy3DNWAvS0izLGdxvS7ZcsAQrCy
J1kBQzzYuJx8lwCd/z9BerOp5PN3HbRB+3+QsJ0eWYKu4llasX3MnODtRgI5HOwv
llC9RvySY892ixxc3qxjcUjMHUKNd/ieMbJoj9ZhUS8E4RAp7q/QNhF1RJgWCbx9
qjjrraGrkaoUPUX2cNH4JAqGP2cFMCTa7QtLL+sVn7c1YXwReg9Gd+HxJbfk9Cw8
D53XMww46JFYY8FD64JYZmlVRZtUGqCOxaYTcNAfLIUapOUPzl5+NmFo+21HiyHZ
OUtdxakQ7/6hE6JW+lRhTkrkEI88+07MBHzaTdEXQawjuJ2/3dd0mPZvY9XN7yLz
Sv4Js2BlsqbdxIqgeaR+m4VTnhmbDkk4In/lTvQmkrUFBJQS/8iewARgm6sDeu4s
oDBZdfn6uVRB9p5m9DKoWUScTZNSOWQON3yLD31XicMmeR5OvwzG1awFr70FbrcO
PHA6JT1aCT1QluUJ4GmEdZKEPrqmX1NhC+5lfQwJ+bIaLQncsa+ojPuqlGbZwu09
XAlFV6M5qifyRV7Rz+vnZsHff8meIkrrut+Rls+2qsFoOSdoFtjtaxscFwUy1YcX
gOgyCHinwtQ1ZKtKUkP17dTEOxUVeTWEYpmb84yujPRRQz/Idq2tWJNeIwoeJEhQ
A03nprfxZ7byFlHxMIssndTmKYzSHoRJCAhSpVcyVdacanEDg8kBdz0PLwmb5BdR
80xvpomF3hp4WQdNbw4vm/bBBiApoNfEtdWkFQMat3LIkQY8fZJgERW+DW7N90gt
4TxpHrANmF/eoIdBClrjpIIwK4bOEDBuAKiT5AmpoyBYzxendyfD9f1R2PO59V4/
TpSnKVqqUfP/5IRBKUZCWafOZXiyLcsHD1uS8lJojnHRyaWNfWP1Wez+IUSVv91O
FOvLMOmfzpNeh9YZyQMBjKpd42NzPhqD6W0akw3zP77t7GkH8l7vOwJI7DXkO/0Y
YrhmMqUX9ze77/Et/UfeqVBr2DnvMWatBw6tbjoNUR4JKVQZRkGuBGqg17i6F8vD
w/IW/QqfqAiSq2HwdP9Dmc/KeVjrDbKj0490ReYj5EREq0Pjwge0HoAvDqcyLBoF
QqhcQMM1TtRqKcj4YPfqzgJUMG/yffeP54tHbRu5CcFNJcGt+gTwPZWT87Y71vCh
kgPVFU7SYmlFxynRioXd2T2v1kqq+TmytaxaZhd/sk/+oXMK7/tvWLno/yBZhS5M
J+F/FF0IrVl5Wlh7/nQ7/i0p3fRRw9gZC2tzp5r5sSEYN/4zVHuKZEksZZqKOYmv
07UaFWVV4/DOwrnpXK0hGSxdVArrOEgpaJeaqtqVeFC/8RsejW14FFJKADJ8hHYU
y+JXP4WxQP6YJTlev3mxJY3O+clREGfDaqIj0LTfdLC+NlpT9VpCjZuLRp6uW93N
4sRGdHRm6Zr4+l9/MdmZY4vEv0C+Xx6hpqtS3OyhYGhJfaUuOCy3+0JlLewctGgH
G66uVFWNRxjdYE+TupcnuTPgZO+QbIk8/OqUIbALZDVtwqhuZu0U4TtYQP00BIRL
BgAPT0JuKxjzvVAqkZfPC72419KY6JNmjMRpNJT6hdH+c+NMKx3QGh4OshX/4jWL
dROZgX1wy+aCZtqxOIaa5kBjheVlLWPSyEiFuusUJWGIM/kegU7hfERVbdvdftaY
ne0xWM5Hi5wuUyxqfSeR1/weceHNCf2HNRy+yH0U816hOx59fZYl4jjmBZHBazEB
EXiDtexVoompTFK9kTnolqEMDnJaEF0fe4vY7oUETerRbWhvFW13d3PpYhLyGOKe
H8xUJFhPNejwKNfK/h6+e2/PwHbFWvTeaq7Q8iA9P6DRaWB/fmsK458Wi8J4rsur
3Mo+DqLL+kFzNnPFXBxvxqaai4mFOeEB9HS7Xplukcub6gAWjZ8gH6y29IgjaCsb
B2NnHUZMsezZ3YwYg+4BXUsMZ1eDWumyHpWi5Hj7RgraTDV8UQsiGAqaV9JMB+6F
BM1MOmb3L5Rdy0dOJYWCTaxLVM3+4Dspovw6BI+lHgqDnPJG7GuYno9fdWNQT3As
fnyMxXbhJ8EabzP7fK0kw0m98CRBaDM98SFs5m4k9w+w9DKxSWuOWSoZJe84qi7V
ETimP2DI170IBKWucGXze68tN3/b2M9RMbZ9KZisZepOGIAlvgPiHM6UPxiGQI7C
XCL5usH1oRiucHSoLr3iyNRKIRx7U3KtGSkgpJNpLBt+VQhHYJYTyJXkj+rxntcZ
YGIINiyigkN3jkai9H99WfPEoSqLdTh8X7J1xPlySmP3t1IDLrI8RqqvVy2jZ72g
cm3p9JDobQFTSefOn9KXdRukWekCzPBWfbOvuRQefW5vgAl+J6LMduwc/YUpXq+c
/UYbvniyLtYsd1YEUYlk/f2LLKrulRvtnQ3kjSHSlVB+/P+9RdRZchnS01oFrlGP
kE3eUgDCOrYOW9yvUJaKCapWN1jr5rqHutrTd21mQXCD9xASb21TPZZCzoqobRyq
dl3kf9vZPRAaEkgKmwoGQAWUFRF7sZsnwxF5rdAGPJKMTTi0no+YWNIuSNhd0Dsw
Ewje2wZzNWxu9JNZKnj5qz2hkfpqVATzsEqFZD4/uxCcGg5c1YmXz+VweWClGquC
dtPxdjPFTV25oXWe67HeDkWVM2OLsJ2gBX7DgJIfkPqr2YeGK7GDTrcSftaGvt64
+1e9g8NyMBw3FbTzapCjJxIaoJwVp3RB9LohwJhYqyc8BRBT6vKQSim11MVZePjt
vdLNKdeH5uBIK4cQcQzbP8Cb/h8oO8sx+CsyBh+NPZ2lT9rrSQaRGvRwsWsPFGZt
G4ez+uLa4mPBGcfDezqF+LnEXm1uDHaXWdnOIERuqPn/W8gMHF7bJmUZDM+F5pVa
8QpxbWJgS0iLPKn+Ih4HUe1VomZT/lNuclNOCKUB6OEuI63RbdqcdOM1fm07FIfO
lVQ0li8QRHp3Jr0yAPzyUAdEnqfh5ESE8gKJD/LPAZh+COloedkMUX4Dj+xDXqeU
Z6nq3xppeCW9tS35zr8Qmem3tWRch3OqQ4eeKVfl2yB7KccRpzHZxX46PlTlx4Fd
dxZPOVGw7Vj/DpkamupazG9TKw+qrY0C40S2fprSwZV+H7erBS0sGhrWKNuWwQhu
fmv3GMy8HqEpfaAVYW2mlJCz1+XYONEiSPGRdKjvMjdDbmOY+L5exgNQJ+leZCyZ
LOZ30NkmPLqRFrSjE+0m24+G8SX23DK9A1Vz6242zq68IswdTuniEA9L3enCotxY
fnGIFCFQqB1TJ5v33wQcaPcpimZIRGy/afRmPr0UDtNlS1SHwP0y8dLVG3Qbu4f0
ZgdjpXpBDl/J9AT7h+wSADutupQNo3PvOqXWXHjMiWY2EbqbUbVwLDw/EbPKdYH4
zcSjubFyI4HVNTzV5AmG4jc+d5X/LfhLaYgIKxTqhXocVkPcegVKPNlOYxs8aT7/
lC0K7Dw1Zt4lRxsQgg2cLEsJ3pDse3qIBBZl56w3FW2Fsy/9tb9tjQb85jyGKifG
JSPCJayXLVjFfhZqJgq1s3VSav59+sMyLfjPo5/t5ejbJSnQ/5e5ySHwOtumBsfH
EKqckvsV2lsRKPgs2b3XLLfcQ3uPI9l4r/JU7l59L3feZiQ4io1kvOkKScMxRAk9
vXrGWNFpzs+vH5/+OTMN13pMXKpemBkCXfiKBKW/8XogmPokjdu23Oo0ZCi1URKb
CSCr502VF4J6jLAhXjzcCw/5MSsuEFT3PaxQ9keLEgFAxs/bAZ2skvyXNggf0as8
pJ1mWOZldvmJrJfXGTKz8W7s/6eyPrNywvG4sFtgPSuyw8b6azyPUSw1Pj8rEOqn
xLLgbcDMNlcKYFop3jLFyyNn+zvpO0wj39BaI6TT0yJSA3hOTb+xY8shU6s6neiW
/uSBLPBmpxaY3BAD4uAVDE1b+wVZQXts8OivccjoAmSKZH4J55zU+oKWLA9gOksh
BA0GvjNfdCinHkkl7YFQpbnxD/67YYKX1iJTAdjCVcyVtE9eh/v5yqiFqL/iOTJt
DsB4UEKymZHNcQK0YyQ+aU1B4d81hSgly51kSBvLyTLwnf1YVnxAL3T1RndTYBgY
73nNkp3FjjHp85YJp0Y5KLueahtDqQIbYPzitVHvmYFWgH7HiQ31D9LvIc6ur6OM
DaxaeKF7d67rWgZuLciTPYE04Scirc8/n3LinTd+1xK8RO241RVKs2lfUEFlkPx+
pE0O1wGUyv1ZVaJUv2uB40bCzEq7UQyHfE2BOBZHHeOpwCXwwUM4wH0cBjTMinh/
Imx4K+XijZF4vsQ2Mg/z1uymM4BUct6v8vwK/Ln6+awGmXeQLx8ZlAVj88JF61HE
KwkiBqpCna5D1COuH5vd4K8iiWKngPuZeE4X4G41732qjW4cAa3bIHpGNEe2WlGa
DJDBXMIfSgNIQSqiWSeaukDjsqr11AngIP4Kt1nt7xNZ6p6dA4+Z1Xlq+EjQ5oO3
QeCIL25TYUTjbP0etlF+8SfyMJAEpOxjVR1j/96tW6Bc12Xl5E/8ITEQ5omYVQHt
X73tsIURFQUt2M3JvCNyGSLGzLFWQEpHrS+NQFxlB3HyWNdTVDlp66IrJUCdLXy9
yIcPpRJhHO1LokykAOpr9Shc+jHyVIh7PYkZNAcSsjNz1cCvlnGjdm9cwtT89TyX
Isb3GzLQrk30dNBtt7haLJ9vcFdAVoTwvJ/8BKUEaaI4Rs11e1v+mWVQHu7ISia5
RrodJyo2Qg6yDaQbBSplwTplOc/BDI8CL5SkuqnU3gPQx3tGjPFhe0d3Fmdj8qVb
7Y2quwyJAfBxtlxWy3DRFCUDLsqly3RKln1sruouQgpVOFIZJepoVflOy+W1hJyo
Z2atHu7NxYutpLhJuTqZVRaVzEq0OGaYfQdMl5wWqo8y/PxzRWSNmt+LjWtSAjqQ
a7whuVxQGjfX8rI+0snI34I99aJoZXIJmDCoHZtoUEybbmN7KZrh9s57CblcigP7
8iykc8EVDqusZaVsqSBA0FRjQ71KcvS/jO4mKl2ZROYs7QH5OVjL9AP1UDnrcn4g
TeDXpDm4uQAcsYW5EOZkwcQwvPpr7DAIEce5Rltj4xBUvOqVBEV9Lv6wxFZ3LLMm
8IulZyWgfg9zuDvUst8aevKTvgJ2GxRinm2ugn0kpvkp7bAv+CoP8cg2siCUK3m9
SYvySprkWLfInNVy1aJjJIVEVfBAtjefpKIrsB8BGZYB0uDoqaXCp5RuEXjAprn5
KstO7VgVPcdBSeruCN+Sb8QKieGH6GRy9t6nx+SP0uarHu2OJE53qjI+1d58WmOK
Fee8lh8twRTqhvkVUe0Ajs1Sx9qW3q6Mw2LwgXpNx3U+hkjKGywaBFNxASxoc9II
teBKBYExGRYPAIFQ5FI2Mck86P/V8WHPKRxJwoRWyExXfKb/qy1Ju8dfFQywRv1r
HI5Whgq7V4hatchOWgeq+coT0dZWq5NW86TDOA+k05kfzI+UjCtjzNcKMST02s+R
+jotg7+47Z8Eywl9JAcbFie6PTrKFcNGQsotus+dtp6Qn3M6GpxfHMtBf0ars4ax
cPTDn5Rru2PGLxn8YzsziBfeLlS9gV9Bcdqu7KqxnLzaEqVI/CLt/6xn8sUfKEN6
Y+XwE6Nj/99mDtI7IjPJQsfdYpLj4bdj+zHRPWsS5qdvi2if1A1Y0H+LGrFgMXII
5RJKdGS6EYXXSJESspd7TjIxlwH4iWypB4foEonvpBGQz7g2XF4g10Ntwr2WkTxU
ttcMnNN1Yt8x+bVGqO041RmMUHGf9aqZRxVIm7aYy1adlkRFiaoAjnO6tu2L16Ac
wjoNdSXfLfygpRVAnIlRXetNOybuyxzkHNn0krXu5xNph9WeN7QOx37ir67OXB+G
T1OI+VBqSbbZYhZtAwEQO1LKdOE+YeJqZZvu48OHyyw4wsf3wLJnphEVUWyK+JjJ
pgb0bqkeSjgRWeIn+eHFit1CPfUGFrIyOA28z85zsxaVKFIQBDXoR5Jc0RULXGuj
CamePFl+Ylaq3HyoUefqbs3PUExcD10NuT4bIUqqQMTwqHfPbTY6bbIA7Q6ZEmEu
FAAMgdlT/d0vm6ggG/8UnfzD/GKXiIUtSW2OOBgv0HEyJR+ufyLfwIYWQAJjVcPx
H/ReCjwKgwX1jIJITHACzHjyNpYJsEG9QKMYs+ryhOAOQu2out11AvBrwk0WCmWs
NoY1B1HAYIQO/SdaIAZF7ndjMiHIn1+/yH//lY9dl2JbtDs5GbEy1vw3YeZqOsHT
heGrul2pO/LA2RPhEtcPgMPzkphc+cCO0/J1gt27ECX6oyHZmPVruxLLsuu0oibZ
gu6NzCRfgHmMm70XXFF1kB2JExqMGT18l+MNbQlvW9bC5EnTV2cnhIMLWzlbYAXU
sscd8+koDNFbH2+2G0F0Cahh+8TH7Lvv+QoaqQGuSPF03HcmDoneEEyz6yHWDeql
Vk4YYWp00MGGcPss5a/GyCcq8AbGE1wqFqJgmhmdCqKFS7v18MxJVob4etZJwo+S
HaWHXv/s7GSlJN/aFXVt3onFzYmfN26JP+jihuw0vC5gSNb89o/+DF02IFzmaVmJ
2nzud38bhAJaF9MbHP3OJwfAdCw++I1J+fVVZ6m8nWHKrUQSjBpPNNAsQ7+FQIG/
gohIfpmFBUH/sJ5NNzBuB2G/BbaNtYEZZ50PhrrcVr59EJOEQuA4LMmXsJD0+HfF
BLklX06zdN6o2fNCcRs0vvGXjPcI2sgdKmzlq17H3zGRrrFWyKxXd5VC3ByuzGo1
loHpuEqlmi8r1eBc5u56gBlCACUr41tPvfsIW19fRA00wV6Lm8CHxvrO5gJ0JHVv
NrCOJNFs4xIvo582hH5xuNzhkeSSe1qH1joxR5uQhfhCN2DM/A/K6Kfd4jlSGKYF
j/4jE0vCZUURKI69ZbaWXiY5MMh3khzCY544NZAKwoBHK6avSeg2PrBn6M9WWHyP
BCihnOXVeBDf/22Qvj0zVEcuSwXHdDNtUJy36TqiFFpEq+TjVlS6Ps/6zSIkBN69
bkd9SqLcPURvfFg/dGwtcRCBfUwTl1CZf+chUR5J6jh+Efcxd+qviReuHQ8dNNF3
fWQhen7sM2ongh61WQWsQ/SrlyYdNS9v+h76aNXr4qtNLOT/SP4JZc2zcvrTDhOo
axVquNBESc42G1DLA/wpDFGX4MFGPJXbvhwEClRW2BlsqjqnQ1z5sFQqv9bjAFcr
GDShrCm3hh6tJJSVqqYy0OHlgeF5ma13EToMQedphz2FsJZi3K988EI3W0EpODyy
shNkaIbjUcjqwOxwLoINOqNNKBWAikbwn1xM9MG37d4voV+PGw9gfMyoTypXQCFh
dKF2hpyXWTfeaSrMl5Weu3HwtDgu0EszJVawqhvVWqkIgbERqSuvV6F18NDR5gQD
yws40NxEJe38JHqp4k6AVvLwj1eNZcrXC2qWmWNfr4cFS+YyBdH4SPwMr1i7zrKy
Ris7J9I/euRioag1CYL1DgQA0HmToHlXHpmwW+bTS8aiyhhCh469UsTFh7ToqudI
Pc6fnEFkY/kb+61A1H14u/uUao11t2vfffA0VQzLZrY0y1im+x7wqK2N2nR2OGMa
ukqsb9rkssB//91rf/92idBtK9DQLIPTsDovtHOgpGcCwueSTF0X+EpN7KF/Qt3a
Vtlu33lskXSjMSMobimoAiO7KEWO7QqIRojawJYPviEgIgrMnxPQGZQqWNhtvwmp
jJcS9t8OU8W4mDrAOy7cstNm0y+bqbT53cAS4YauTWEiIo9XZPmUUBNWALYjfBwA
xYFincYU1A8VRuZDqf7YYOMY50z/F91Ea4BRhDfrefbX+BVeGJrjbT8dpn41nXpY
6aDCdgS+bUfNzm6KwkyDkol99D70q3aaKB/ql/o0Kqtn4RkESbOyho4278etKr71
NzBMa1ZwUTgm1573v2kqYlnOU7jtM4Ocw3MHAjNrcPxRG7d7smP+s7lENFyQYYXS
cvZWIaD9tYKnfXJRy45yH4TtFCGiwGtkhv/YftqnNOKnr3Qf1qb9COlluoLrmwc4
DcQJszs+GoIsHismQNFkb3LB1jIR2CoEXiZJ27uGoiPqNzjARD3RkgUOYcn7zkyn
V2I9yR7ZKHLQDMm5JUIP89vBBjopvzqWMIWU+AxKoJUYQw+UuBCnj2PAqDSzbC64
SZhgswa9+792kW1qSGuoSNfEQE38F3Bn/J2uOAcAYgDumXf57qjEiSadta0p4qqE
1a8sWyr1s8dxyCEZOnRuiQ5TQ688rpA5pPOvwF7kNgg7+k/VKmCwDE+LfcmaUUvi
ZWMFgFLOBf5sApBXANA5QXth1ePmIN298Dhb36FvZ2y0hgUbmw8UnaXxdSGsksoF
JhRUo7BCcqbMC5ja3/rm05OjeFW5xlw4mqtUX06Hc6aRPjHdkB7FiHGkv+F5HG0d
3J/pgRcdBxyqaNUvg3p9/TqrYDhSPelljz8Vs2LxozC9kuk6Rfpm9Kjz/9BQiYJh
DJHGpY/CRO9WsUVJgF3PRXMkHFG/6wzuqJDBtTSRmn0WX8SzthDzmVffa8idHf/p
uPVyOSwu8R35d2h8v/C7+jlTMigdr/DhOLn8ZD4OlD6E5W1FD+SshJAW0yl7oWCJ
DAd/1+CrjOVAI/q1fb4ix9v9l7w9PLGI7gpuDjIGyYKFzqrH5NHYOvY8IOcN3T5o
bw0v4Br5zSuqLBRCPdz6X9kd/iBsuMLmd/TX8BG4VVIuEWNxovPxv/lgsxsQQ/aw
1zpMkJKIWHlAxRHS89d0uguezbOaha+H+PxT/d1IGlhc+/J+z4XWQrtnbndPpDf5
I9PRvq5e/BfIQog+X0GWBlrkl07CcIwouMTle2fpWZiQgeIpPyoiaCEtYt+9R4z3
vMXwh7A20bs365gaP1u+ZvdbdWPeQ7+yoNiLspYr7MU5kcmOHRTzxpANcC4/2gjE
7hFK2zHgrQ9B8zWoHSW4ZCZzUNMt6K2l4KCqX+F67TReiCdsKq0GNQGQL5dOP6ZH
zMzHfmu4CUHMSBlQ/hgPTqUl26F/qaODfhuVAhWbkViIJVPBqJ6uIgx3NHgFTcE1
GXQQYHBW1j/Fwg/tseKkh/IWPT7Fz3jr5TZgPryA/IFy9T+zAmmpF5Hh0rw/V0jP
X0v/emWgzE8BC1Rv9VwPL+EEgJvcijNs7fuVx50xcocWk5L1FGhLb2ntz70Tdq7+
V0VdlAPBvE5i7nqcphry8CGVwX+VP5Xjtkw5EA0em12+u1BgNXj2s7PZ7wkXaviN
4Ugrq48ZtJpEsZ1ONai5X/ltSZKesiQkS3uWSd8JEPYbrOzpKFZjpxFIobIs6yE0
tRZXQ+XjNtNrGfFJzma6bLJUNyfFLC1Z7j9v9L/iDyF6UnwOJBrWyG1UgDVatuoL
6/Fd/W8Db2O3uSbCfinO0jGb6zx/Cb3iH/4ggQ3d2KbHNLjj+ez2qOz5UnGmhTZK
u0hd2WjICzbA/3kjCn7vD+X6yV1g14/xBLqcqpWmNmqtXoSj2Sk5K2QyHRBR7K8m
N+iPwjJFvFEEfV4Dg+yuJUxAITxjBQa/h8IqqvrF3NvzdhcPwmpR5hSyTVzqlGW8
Jbmzyg/9TXHwaeuWWs1xpIVl2D2LwxYtIpBRxKM2BdZG0Ek1J1YH7iKjuMtPdqci
OThaP2Itd0V8qmdhBEW73M2hhQzgjgwVIuPlQ8hzryDzchnAKhQdDyIj3xmEFRUl
QfGmaA8Kv/stL2/0ahSQ/kX4BMBMb03fLLqg7GVMofqoOSJT5fSq9EjFCn5VFLpO
ymuRT+mVPtORVq1G4rj4+KfTPgBW5u7bdVC+EzWLboIsPAhLeCp1GzgFpq69rvCN
essg9k7p3DkXEA6zKlDaKsdFlHGfd8IJpE0jTd455C8z0cWJkBGqjJDx01O6Hqgv
EOiemP7BDs0Wfg99Ytm7SVWyNcXHOCpjcPEBGsmO+IBeR8+ifXi+GwMH5VDCbOAx
pbnqJWYVnvCwhWa83oT0TnRLTLmcjoY/gvkbx4BQH0hmDVqraFu/uiGXeu8RyP77
8f1JUiHQeaoRHbzpxZygFvbUBBpDngq8xYYRo/hB7fdN/jmGWydICHPE8IXs0ykE
Fa6bTKuZfd4O1OKyqR6NPvOBwZoJUTb+Oj3ZSN4AHD338EH+cpQl39CsDqTC6YqU
01DDkbwiSeORKReI/nuop/75cdtoRiWI0jZubYwDjQWjLhXEzCeAILNvce+vdynw
mWJLpUReK//SCo6usqWgQuGSOU2jW4FnmtqapRYur4uEm4tYzIavKTGPQdTJflxF
czHEc2/V5cNCihSItjjHwcYO++0sz4r3nkU1e/UMHdjYFYiBYfK/2uxX5UWoJo7A
pVun40rrI0hX6PMhuQlieD1lTiJCy5TRXs0YhUyQbQVIQPZoiR9PxSwWGAa65CXU
o7mfWhlPK/WoXUHcihZKwrrZC6v1dd+gl/q73onwsvfH1MPBcdl5uMvDkQpTTpGB
eP/waZVO+JUwn56Unyosw5SF1XuJK53SdLznsnSpy/9QnhBhRYTfSIn25cp57OsU
wfpJoD2HTATemx7zNosAXC3yaP1J3hTqxF9K9j/cwOtuV+v+UhMGRjXY01NaF9fT
U0f/6y3wGPIdGd7Ixk++n7j0SOsd08Qfaf7hjJ/EUnBkC7e5k7zZKeYb5FJD0tan
NjyrZpS6WUaN/TPGwUdFrWEO8nJRuklXTeMnWxzhkBISYLECV1vxUSBnam2Q47jK
uGjrwAQ7rtYC6J7BAgEC+mZHuHLzKZpa4QzN0etvDpKjLezFKfiTdAfrdx2drcMc
ys70PQeyd2njzWhGrp26r989ajp335xRh8egFxZz+4a4aITyjQcXb03bAtNeaFr2
ZAPkZCxiY5Yc5A/kwQhAeFxX3abuSKG3OS83l58elQ3j/BOreW5hwDhsUn3Vimzt
M7PCIOuc/4EYyhxGVQ3/Zrz4vMPusKDR88Uhu/Jv1eWOnxfGb9070bknhBb0By1v
MaDVbzkOmxx/Tp8zL1+yPDfwud9OSX8cP/oTiOKIsq5PRBxwSRFXljnFqzuAdkkB
7iXACqw4UeWZfDMbcjXNs1tUGCYhR6tp2FwPJI6AnIZeWwOoCmIfIoPLX8HwRJum
+vug5SUCajV+5dO5Cjl8A7pJVxjB1ZMNZhRYmf4ePqWT9hg0SUJbLVJEFojVesBA
+IRCWbwjKGNYipnNdTbmxWno2I703plUTrOHXrWar4l6tOCt7DzuY/otSsdIYDNF
lHJcMeshC3mWwsiXWfMSB6UOSUBUObgP2IoF5sU+inpvhFac2BXpRndBzukYFj5B
isfNFH97ERwdTlg8pktGaTinte8V2zTYjpc6zuDMGRST4MbYXIvF0EJtFfVGs/lB
mHio/25ByZV9F+iltt4zDNdf6g3XgkYGjk6g7P2vyYhPdNVHstEq0Av3jFv0ma1u
Gc/qPnc2Wg6WPyGQgypGozRLySQIyUswML3B7ZR0Lt88fQNhmjGYhmAjTPN9CFXD
uCtcLwMeryFZaXhOkzgW1S3s04I2gHxGtyMmxZNp1rtxTUUBiHD3LpaUoGEGCvT/
Ueyy+qlZHdshzWAjHqO2FxkJh0HWAGVRLB36fAtjKhqG2h3c82KiYDWfIvgDYR52
/j9OEk05bvUgrbFZ5iBjV3IrXvSoa3po/15PMHXsPedqqWKnebACkdRG7Vq0URDO
GTWRoxPEyvHSVejv0AxB4Mgtv3h++iZVNR4JXkde9SZKKw3eoW0c/DRDuRQHgjFy
cBnYxAZ6DZysWDWYqnDjZY/sWr9R9lX9eUMwTp1WXJZ31WBlFof9eY5pjGiH8zDK
db0b5bWMEZGsWanr7FbqgcO8K3QAnlR4+x7AwEVPCi1+zZ0gs1PjSwaXhNTc/MkD
x0F8LY2o9rWM+4a3SiYqPaiQp7lgBwffxfD54PD1NBywQ8ZLNYwBjBUpT7RpeVmG
XaRzlx+fj4+lR1prRbO896fPO8VIZiNIoQlDE0jkN/zSFqwUYLDV4RSnTzmQ25HJ
YblXk0aLs15unuAKukB2TkRLNQTRguUP5rVlkL4qhPrD+bU1IdZlnkI0qlWgLMWA
Cj7W1NOfahuPeGKnUFN5BliTHHtrwGdJPBzKr++r4oDEqrG72sDFl7c6O6hlJsuI
kPELTMNC54aVrvAxxTpyIWswEcDxh/Lv99+U6vOQYNJjaYkVAFi6nnRWZT5onhma
sUJDgd3+NgDf8MpzpQMXA9Uyxw+XeQtjbalJUEqTCiaEQew1PNq6QRl4MGFzPZXc
5OxPG7LaezD53Nbou/Xnrau2aNBwc+HaLinV0y6g41wY7oAsAkcKlAaeuxEtmrEL
7Cltrsgm2YK8rKD5xOG5Elz+aq5hBHAFI1DEkPydkWnK04qX5G/xdbtUCPZA0s+0
6JIIvognveA3vxc0EMFvWHbZWFsEJvFMkcHWO81OIHyWTKpHOet2b9wThTuWfa/l
Geafj4KvlkjydAI/1moS/zxbW52OUf7tWaAUeob2eaUln6bUHBBXdi1/HUsWuTiK
0CuDJgOYIn7nspGPXhWwdOBLE+KXLfK5ek/OLKkS5y6RnNWET9HaNjH6v1YjBDkU
Q2hGedtnHMOzYhxm03o82YHKRwhXX7ZyF6eWYra437i0OdV5mJO8+eMisy4zVp65
pKkdg+M4YHvRnZ8eYnCbQYPk2yyznG37pS7Eo3P6oOePR7hv6/jgAfxl91FyKxXM
8OXfMx6Tysctu8ZjU+ZuaRLitnHzOzIdGRS4mrsiDBAsXfkVeVnW2IdBaXnZuUzp
MZvwOa4aFFaBQpsvg7dO+DSz9ziZtnGPsPQXRNtbzoFBA37FYfWXAmPTUA3XmBVa
/h98ESoUMRENkyssc/+pBg/wmSlNFOXMdtPW6aVTzeyvuz3gw8jg4xo7YDZJ3z2m
x07iU4EFZvFRByqOPUqcLb79K2Zg5W5KWyngQxLE+cePoD+7aNsGE+4zPTM5aLAq
JeJ5332i8HELNpDg0r3nLxWzgSX9xCW5TiJyqazS6mtFi+XCiNgxAMk0uY9shJR3
PD6endE2xTJjytr3DnJNA/GyqCvOnWJ3ayhi1bN4WbMV5RPWtnjJA4w2gV35QAge
gwNlj0HBLL/WflJasXAIxQdvevU4u5BC1Ogx5F6PaoFeQqqlMJvZCnbR3yAZiFiq
GF8b8A/RFHnlArjjZ1DQhHLDkt1OuxOB8hLr4Zr3+jZ2BYHqRoMLy0g1Wj0LHDqc
rAncvojU+AvWDylBvjvnyA2ySI3MAzUWLPF9UYQUUhHq2VfFabmaT9FVBHgOmlCw
heEcWTmBcUgo/couIeL2umi1iwAT3MLbUOL5Nbiuc2i86GI1jrYw+h20hc0Od1UP
YOMc3I4lIZqRII/hmGDRxGrxr+c77mR6FSNDTRrRyD+Qx5/MOxPVdthRVMs8b7lB
R/068iQG4dweqgfZinBCC60yoMkqAZQCYBf5xf9PW5qptVPMFgNJVNTYpptF/00V
jLppajhOcOdSNZ2YfFD0sK2iL5resgB1tK91YJXKbsttXk3L/+sdeREb7dVaflc3
+ayAFHMhmylCzdXrSwhsw7jdlE2ZQV2aEqJlxVF5TDAyNOpOZUU6X9M/YRoj9/sY
LYWAbxEI1PlEZ/+Q1vbB3l5ZA17K2dl89lwlj+8X2gR827aLjIranrZsJQiycoig
B0xCdKS76YjUlPH/MopcXOtbFWbBDMYIQ6T/KwacmKK95vAXb0+pNhESW7ptQmVZ
MEbHYbReCHRkpTAb1oN86LLNYejv6zFjtH8uY1ezVq5QNMdP383pZbPBfTEmXb2O
hlwSUy9IvwxFwBlPut5huQ9DEGe54o/mTKSKrzXjcXBLsETcQJSlY9YiCQpS4ZWg
mSk5stWE+sT2u7B1SdvcKA9QiEh0vNK/nHTjEew0D4n4bDlH5v91eNLN52D1zYu/
fy1xkzYbEy+/pxETLXP5pJ3A4AGN5mE9gsMi+dXYfHOY7zPZ2AWvP7UxWdYGR6vt
QB3Zcgn0kFg0csbAfXreDv+qDzecAkUdXQ41QFpsRrFQcwlJRDFHLA+rWPEzFlJS
5uHRQ6rJ1s1UtHIMQT07zpnJdxj21iFnU4oV8Fy0i0VNaA5lREB+e6/muqfiW8TB
oQvVfA2N2x3WqNhnLi2tmY7TJTFbjDhOeNpS/o+LOjgQoKAqwPA9vssO2Y7ERBvD
NSrKkHeMXrg4emkCi+srcKD8iHSdXWVwn7T0V9A26p9DpgOitZGg3Nh+5VM4tqqw
8y8nzx4W0Lrtgp/cucj3xEuSkuVYScUDZtpjrU01dj/47Jq0td09FXS1Rm5B5Pzm
4QIxpPIK/v+B78v0o3mRlJGWav80cuZWAuSqXetmXPkSVIBIvohKrZoyTAmuoxrK
2D1NDWBMdADkoFzfizBuLHLbPeOf3skFE1u43UzaDYabAzPcaAoRIKzo6QPodV8e
Shbe7UvFTfMr3elpJd7lDcjuk/Xx+w6yChcv4jgpZfd50z9ORb/MVnBhD2SDsERI
nKU1Vim7umgk+MI2T2nojLxxbBzrq69NntP8zneD92d6eutQBDWbG3qz1JxkW+4Y
UsRKlxan6W2aahvPobgEamoAn6H+l94gUA7z9fkj4p+kjHtlyY5N9NXxaeNzkBsP
e96j1m85g6wlf5zByIOypnZ4WmFc+kfhQkcpz5vAx4aJAmik1ImlotkbB3kPhvea
vZoKR0rbj4vDE0Jy7u3+RoOlT5Ue6N9488sQYWifnrSzOZ2QKMb1MU+eIGNz8RVw
D1yluCnHOpaEy6To3QIJYHl+a8zbpE4gmTo22pHBPezl4dvNgR3fGMicdGB9VMGA
iFVmvPyJ8dE/14JRnn2ZQHbP1I31JVQ2hqJ9XTwoNH01hT3/40cVj98yf8HXcebx
sqGFpGWLaoVZetTGhdnILpCsZ10m4vdWfrzUUfnEgZ1f52rl4dgkRSDRc6JWEyAg
A3EX7pqOtRmnX3H7n51pPWHTwTt5MadgZ4Nmi0U5YJd8P/YA0/zEeK64dQ3rPB/b
9tdPGKyGC00u1iCosb9lRCrbURhxgmXkw3xcOqunYS5qwh/HUd2ftUuDLllR/KIb
lX8r6/KVAT6JqxZVqjAM9ddrHktyWvpeAKltrNrXH2F4K/kOo5Lfh6MKuAOShdFK
BmcPsNXdRDwIuJEnlArU3hDeMwZU+amndu8GtROW3ZKU/a8mH8KSKwtAOKaePxp7
KZyiuH4OGdjbfeZwAWvxCDAGfFZcoiF2TmXnYcqFLEsJrfB74vaQYzs6BLzrhlHG
Uu0UcewrLUxSGI2Jmw4BFCXpXLHLYdwYoIX0ZnjSchmkMOyvPmNW5EtiD59rUglr
AMLy9AUgOsPa6wkD9OO8iZNWw+zO5qKDM4fvY2na+9QCyPFYWihhuGS1491y9y5W
H+0MZORMEueQgZA/Hyg0gukoeNOuhakK/Pix8XcU//38dfpxToX09BnJVyIZ2n+4
YaLegkp+wUCnVnrZchAKZ1v0lzewHodjVOAnx+RUKqywFGblRnzQpTMCUgoKGZ3x
CIiM+AeeZWed+XbUd3yTZQUsKU0OHoZfXOrMK9edrnsWtkAQIrqag6pQdB5Z9MdW
jC64k0SI4uZZ+3nNFWHBza8Tc8vKx/b3fomvrlTl0oo6e5TuQdgzXqLi/Czfw2FT
mlYs1HDvjUiCVb95Yqe5OAXNmUwxrzmH4UljYidjuIv47mKKZQPzpQbbOXNLEukE
FFt5Ws3XhY9OYRX+C6s/B8RGreXXy0clNi9sG0p8PrbXOEQKwgajdC32p+VjnKkS
D5q1aX1Ph+o6bHtErzauwYQ22Q14p4i1L8WeRSSwIr43NHyZsJ9yFoTdlTYOulIz
l132ve5ikK0a5CeAgh1aqUDIbgaqkU4nYJQYzM1WwB+TefJot4tNpkr95G0zOyCd
zvBhAuvD2HUDHqrP74kRgr9v669rpQ25YKNUNRkGNTuJGcNJNhxhqw0sawbnfwSl
LTqBSKIy5jMY+87FNm1TbShR8uvlbN+8v2+5ubjvgCQfZntJkI7A2eT48UOwSQNL
IxJ9yC2KiUSVxDpeStQM3jipAmxK1eP/+j/s0ZwmYsXbmkEY7cUG2e8qy9a0hKUW
l4JPnCRd3tRD5MTutkP2H/3dyAYlaNAQpy7uYMbJ0f/l9yh1iuw9uEso4IEaJusf
ASolZEvZ9xgLr9EjM+u9ESY47K5FPQbQqokda5mXW0XLr8elKDbI7Ubs+3LeTVnM
B/mZDQR5BNEGZHpFVuRiNGPbnvBIEJeevhIRbkc/LgUccz8c/gAsitDUQGtwVQK+
yhMCOw2nQo29qvmOIkROY67J3JMwWi/lhe3aVosBFfR7yS3BPJcNB+KmAJheuhj4
HT08CUqnFK7aqCAU1PTxlxhBNgUR+aO/Gi7PchtMqJSx3x0rajcjzaDRUwGVewNv
hRdGwvqIFCW+hzthPF+fYvfn5NG1udYY7tJrx4+GpzeJZsiBUjAYuqKwwuXNaKc4
ZfjgO61dzXtGCGMvy7rANBLuqQFiNLPR9orWlbN9GjlJOECettOf54tHOs5LVH/n
HwfLFNKLqqe0tq/AxEog4tIgneWs4h22hYt14C4yh7qkQIvUAiv1H/oWrc+El/7E
F2jQn9xu7X9l7Hxo0Ned3nduIds5KjLtSWqQ1GVaktZoNIkP7hXsbXCta+eKYpfx
zD6wuBR2U16x8kfRqSRhXQFS2mY7KnXVu7TsPhM4IeTpbP9RIMIuiSs7teC00iYM
kYTAHlACt9WetCxvAk2jI22dmu+Ttqv7rS8QXbe4U2Ls4BRkVlFbhxGcTUqNOOxX
pGwQ8irTYtv+ExkfUBYSsBhHKqJL8+l4nuzQ1tj2qdIHzlX85SAgK+1yZ5EkyUCd
rb3aEXkBWTQN3AJwohgWEWNoy4P5NgvHcnLOGlhAW7ArfPPBoTPHdGu9Tbi3K7uV
xb33eMVK9wGH5Z/PNJ3woCiva5F8DP17JIbaGaVjGHGPX+JlT3Z0fQEmYOy6hY1w
9ury/cBJPGcb7ZRcW7NIH/dF6jLJimjwkMCPTgbK5QYKw5Q6QA3vJHHdV5ZUzHXz
KUh7yv4sAwhqC80m6R9SCPMSzlBzSgT4e5/Z9O2E4dhv5JLB642+vSXPv/8HKxbV
vx6kWtzlUNyEr6bBWrKtRA00CCH2vnLhcT+F1VRZvh7i5Mp1/LBb7s46MO/OHWNF
BU7a7zjWneHIlBQnQrXDrW8xBLmqSVeAILUcU1G2Xgtlmm6AfxSAN2GP4Rc2Mh8s
L9ep1R0VgsGG4zccUs0o72RPKOWNxHyOTQC0IjH8FgH6ybLNASo5vRIKn+haDKfK
KX9Qlg53HPl3gl7maAQYeUS6xmuZTCOKjgnVYfszr7DxWpGtj/Ap4e3Quq4CKMyf
ULy8rQnCeHnblYhYRCkbb6KJuoheZKnvHhjkKR4xxC18uHuOcarDvXMqZN7/UFC8
hVVSTBWnNFNrY316ytw3PsBxXdFy2fU3je6ph+LZUCmrI5WN53roYZfMhMBfbL4J
rxOEIsdmb3aFLM+9ZziDWsQ2nSifgt/DdGycXmreVZRFU0V6KQbJ9wxXcEw4k36+
md9F3sagBL8V7bOkHbOYsx2Vp3U9S7C4gk4m/sEgiyRpdSB9bkfRtSunALd26pKf
4tHm4q/olDlJvHv9xXtwF+ssG4PiGoFeJnImYWoTPTieea3tZyAwfFDbJxuyCyE3
bO5HTWBuitfHh4HsSiWDi41qjxKdyvR+RJmZwh8bu+xiRRnP+XynNvrzIoWx9esV
TeiNIMYmRlYc6nTzfLDWmPrDvIw17tJQOPJXC333WZ8Juibz0Dbs1HMxnh3YCY4F
IdJ4zAwyZh8wuGsHhpPwAOpDgrp8cEj8eCRW9cepnPJg5jy3WnXJPU8gfSE1quTy
efBHQfu06Y85Lic3KrBJoVKk8Jk9vnVS73+96v/828N0m9WOGuHr3ISiTL/e91zx
quUAyFreFk69cXChIiQCcPOA2PoyVs+HLwJVoMUy2no8FDviG9edEMjQUnhI4kvX
AjLUynpGrmjDRDPz/l5qLyvniDnOryVgA+AuJUAJ4bv6afAoPod8IdEQgT3RPKbk
taqRu/1W7EvIXiXYftfh6wqvruwwK5ddN75XvfBGaRNg3PlWOn6rK3DdqYftUi1I
rs9ziavSfAw7bRMksNqA6m6mEBR8SP+mBL4aBAdqLOzeB4Et4Rrai7Lg4Fd5BAE5
GZFebD9jOaYQNuL2xYSy1XgEBwDjQkGwXDvzdr8a4xDJKAVC7WBrUbJPCN+cCp+p
9E5LFgDJ/gjrIx5WuAtNHquPTWvI9da/4inq76Fpc/aOPNoDQZioauE/JKymjBv2
MEKmwc/mHyX8ekjz9FiY8M8OxAhpvWovSy2/oeKtU4fLk1/xyY9OlxTWMRFvnsL/
6PAgk75JWUDYehGljYKcE0LDkafBO2Erb1BK3v4CsZrmzAfiTnHSQRDsb5w42q7J
Y9Ju1vHdNfKCAPxUpqQqEcWG1FNaP8zn0r4PEoAG7eBf7iXHNglS+J8Hw4GnjN+B
B/GxlZ34m+Q8RK0mFA3bc4rx/+iM3hTC919shUP7clgivU+GMMmwL5bI4/7HSUlo
0OQqbcwvjzmMK1YExTxRWzcuJYr38tampQwCWYmf0z0fJQOpFso9uc0Cl81zkI34
VMKet6SKjH7IKbU0enhB/O23iZ8qggWV+/oE8kA8VyG07D99977t076sDkmqhabo
mUVaqYWYCtRuCwdvVw5SNhER4wk/no4lz64Qyw6CpPE4Vi0Ko0070wKWnOkYwDUj
YLsqcWDjQpewoMnDzFLMfgZBMiUshVm7FotJl8SguYN7lQb5PrxfsxlCansXoYRM
dW0UJnSeBCeLCFvChTQxmMqJJWywpI1iFNrayuTKZZznS1J87E0jpJzUCu58Wwhl
M2FDG3bAOydR6wkLa4ppdS7E2pZcvNP4DkDDMvhJP0IAJngw8IP5tb308g8VHHNp
/d8z1DFJuJYU7Xf59M5BLmPdRqa6z/6L7Nx4CJ7BiZfayCGAWeqEgOABdjru4ZwE
S/c7FLaY8nrVQOJggyWrB9yYPVWI586InSbZtkECJ+dp32DUfv0/sBpUwV4SMhX5
piHL20AWQJ7SUR6qzrqRK61kj1ghD5dMuQjovEjvLZQQbYwrIMAeVBm/n7+SCDiu
vCdyFHGMJfeLIaV5+EnN6XWn3y3xFoOoWiftrbgMraHH+z7nnIFfo1nm3/CJTR0w
bzxkJQrXt4Pu9vj2QWBqJJ6m4AuKOec12mxQL9XsNKIigUkydI0Ovw5prxILAHsE
5Wxxl8UZCsQG6JmkwnVKzgbd3BafDnBHLbSLtQAqcLKrUU+4EMJloXQRpyc9kGJq
xeBbAJabzkGPiskkYBf2bup7JStmS1cjxNzK9Nmm39JySBHNeZQEtZNZm8wZ+cA8
vWShJvjAHdFya6T1fimdWcEUzl5s69x/UeVqXPCLpcNEf2bv3OoqembXeWtNqXQX
E3MsuWGxxGxP0TkpA4Dm0Lts2w8Bv5X9TEdlkqIIY3/5u85D3rhb+FrMrK9PpgGg
eV8RO7FQFF1ufMquhb4u8qceDnnSpAzkqVaifzI12UKPo5DlcTLeWT7a2WVYXwTA
mtQOHnFdDbUQo0v/2AgLHGE7V6ml+V2jeKapdFhjKC7l5JMEm1265bUOYe7jMOzd
E2Mw99XOzA2ODoHO1kWf1iPo+VMIiUQIx7DX+TwUXA/YHZaRGVCO84RehkZVmuYm
1qXDlAMr1sh8NRRwYzG2o61T36CVXs3NZa/VZIIKiRCrsxSGIq4NPJkpPVrHLT+0
6JnSfeRNfN5mH9i6PLwL3gu9CINbistdM9KSTKiV+UTa/2p3tRDpo1+oFjPMj5VW
CZGryRtdO5Qv2BIOxA7PrQTDe9ZocXmI7awglASqh6xqlp5tPCDnroKwBfH6EZEQ
Uuj1uWoX1Xl/EtlrJ/8giEtMVE1bnNgTiuYlLJ5EfzZ2YD1/8LHyo2sHo/RQn9W+
P/pARZDGXnUH1+903Q7EUYYllHiUlHEKa1pkGEj1+qLwNHahfAztzCwILgoEM+Ht
kGmKoUycNiNM/D85e/EEudVcjd7vz3YO25WyWkFksWs05nAa1d8x5C1UPKD7/Lwe
0J2GnhKJMUM0dDg0BJy+0iIfL+xJLKCqHZawi3Gh0UvOIRjNjvNKN3b3I7pXW38B
5KVcPF/dItzVVw4qWujMzu/JBnS2EMtqCWrLjxEHZYrtqnEU1SIMUsW9+HzOmAdV
5+SBeoEmckXQkOAAtdYcxZVIbrwQXnoj9fVX03P7GUk/yMUvj0CIKvgAR9edC7zR
9spwChCricRxBGssTQln3eec7LAw7lShLhKvrY4k9Uf4Hecmw8dA+yn/BgeUVWOx
x90854VRdPEPkC12AcUbTo05BS8l7E0J1R0/gZQJ3iDAN+CydbNqP1ee0VHeDGTA
xvk1/oealsWmPHrcytcEqx8fu/MRfL2Qe4oOM7r99qBXrx++XRj+vNbSKktzqZkS
PVrlm7MpT09htov9qn4uE/A0ZdbjD7tycj88D8nQ1ZCwqigK74tfPdgEbcF8wEuD
rE66NV3bVr86njpqgfwg+MldXOD47kGSfrTeVYRfdCW84nUUlAuktGEJkeKWl/Zl
q5mkT3lcaOcmMLTgKaw08nc1LHRbp9j8hWoIGh97Kt7J6vish4SGTmH/C07WDU3e
lCg7vof2MkvMv1NDALYqIZYepOeXsrpK4hfO01+4aIyZkca71bWwfTHSw1esS81X
CicpaE64//xaECe1wd6AFrYnc8X235Rl6WYO2o8dI0AtXFAIoryA0cYfeSz/fZcY
1159Ns4y/iI+BAIfUtfdd4OtQXuk7EAFrYXXLdcEAIzLSUR0o4k7liQOTLTOPEig
pKqbj2lCY7iAP3zIIoulnt8lxJQyKym6ax+rNnhHwDecHrSJM4cZlwOKK7jZtZxq
VV73qE2qTfOe3vsZbnNwiSCeELnirt0nWRc6FAXKjlvickMUVFMu5ZZNgK/nL0zM
BIlv1a+n1V4U5rjGvScHSkGnMo0IriBTFk7qr4E5SALk9KDb340smjaFlsiZJYCC
xx7oTAe+/eYllzQZ6UFlLMqBsDrwyB7ItwERgl0mWUHvBS4W+u/60a7ucynWBWDV
5g62Wqo9iBZc2sZeVxFZRR2ITa+IVkAq61IWSW6bpQe6FofbENirbwMFmTjaHynK
u38GInegLFncruy1/KJB36Yd45liXu8D0BZ6rPzw+YpV/cYZ/oaa8wuJRv6GpfmY
/Zker4cF1ommWwXJbC8PtmU9EiETDNhTieVBdD8GiSqo2eR646L1i6ssmPwSZ1hq
gXBqZSf0ddUU/vGmFmy2WBDvY6SyyzGZcynQiq4Io5V1nq6JDT+z+hOkwg9etAK7
7YzZoRXDGPsYBtdivm6KT+nSvo8dv4J2FeEuYwJ20bFDRe9qYetFeI2pCci3aHnz
zbMxVK5/r/3gUt7ZmDn1Gud0bmuP14Bg9qy6NGqSS4sBsnFksIE66UNvaXQcz8qB
W94ejQggADr6Nhdawt3nx/PYQgBHVUYPtJHKHJuBSE7ucrgwp+oo/v5QOW7myYVO
b9t6aCQxrBW6tqHXFIv5W1qtBjZkalTswT3o1EE0i9pd1uZIRva7NdYmJzIgCfmf
nLDE6Ipiox0ozkvcnUTsZZyS6FNfiHRHyTyHQZObQHYGOHmlWVF/XdZV1CStR8Fh
mu1tClS2ufsstJiLdSieJuEOnnvltjEBS9RMoLOpuHz+T3Tdrhgltmol8cvzZQZT
fHyy5a3afdMS7IRFqs5HSIYo+zjiFNwMYpTdGm9jG9anTTx4rXshUZFdKwcYnz6z
TEKlRslNO/zI2tbSf/e32O0wkXbVQ46yWb4z6OoLf0GgESxDXYJQxF6iZI3r7e+k
XSz5QYK3uNgTnWTlNe6Iey8PFhMgCNRosZl2V891gSQpQAx/Z4sFiyQA5Bors2PP
BWr8Z1re+sOttB2CAxuu9kdbKcxEfG61xwlJ60E79/ZjROc9jaGc9RHHTYTnjpeN
tJpC775KSUFu5WjL2+Ng5/r0RalVii3L1ayyDbzoB9nEg/DY0WB4waqL1hBG9TDS
FA4QHvd61rOlxteOuy9kw1zuITnChFykRkgCRkO7ZkVsphXfPYabvR8PbjL6oD7g
z7I2v0BYZbXsoWtB/ATNSY335MhSSnNXHEDiNYFchNAlygWoWZLX7uduQOmGa5ih
sEpaoKVhNitWWtnFa4gMA9QrHRUcbevBvwz3/DWm87o4HclcqrEeHLZtzROFFDiQ
8egXHXJsyS4r990PMFf4L1GnyquHt5G+O2kAQqQ0j1uGLov0Rk89g4Stb9f4PuCB
xJyEr3+saJDBzRvhUqzT+mR2ppYjckiMAOf5Z6QANpunk68A4ZMJj0EvKb6SDF8I
tb6qkgvEo8mj4Dw/1wLETcnk5+cQwlxJrGvtWYXeL6eo51vHvLYJ8PrcRtSLTQpu
TWJ6Li8X6vCcuV1AVQNDaQxXGqrFc7pU3sARb/Zi98w4cdlWhXWEQT6lyC0YtTXb
ul5AINMrJgfmYZqN+yWWlC7m1qTwmuDu80zTqgN+OLATAdnfPos/FyBj1mQqfVGU
v/7+zrmu0+PVzkpbyqSInYjj1SgYgkbJwXUiP/5A9I1W0h23Zxy6sJIPa+ecyC+3
g1qU+2sbqSKPILGSXwA3W4lJCsdzdJGRrBdBz7T7/xZWyHOEQ8Bz3AsE8VsGn8aL
b0Pr/o2qgduZmENnJKSIsN24Srs/gL6tMM4lTLh0kQ1dBC8mRCILcFp+IIPMc8kK
NpL4PTl4KD5iC2iDwbbhXJ2nsqWRASp8im5KbP2dz1/DNzLHIhOMpJ5OfY6h6K0T
g2HjMU4JMKmDOaFPWQHME9i8dIP1n27Qpcj1BvzrOsoCAw2p2sMpMSz2JAZhKJ1H
mUnhMEk7nSLtVfMl4mjMoircVFik7aHd0krPEtsppIBvYqNHSwO4kz7ycKLjbVra
kMOpwuSeDY3putOqcJH/rLPRSkvdMVkGfAp16EL74LVArPFysR/mjxCeIh9bkzkb
B49KpykSSjWW60x+S+g421cUnxz56h27duZI51R6+OEZeP8j8Km+lB2KHZL8k8p1
brpTbvRHt5FAVekg2X4i4tpQu8NLRXVyxTeuhrjOo7gkd77mUuBYUwg1RG8hjQph
tTx3r909uKja79WAvFc1L5S6BsmW3cKi4eP3WYVnpbI9Y4sAy9+HSybvvMh3A/Pr
FWKkaJx1A0L4a8Kiw3rVIVDkDTg7DymCCzNIaAMCOrToMi+mqpw0VHw94ybJo3pz
6RsH77qdQTqtjFHbHTs4XgiKkkvHAuxdRM+9cM5IkCN+God4rQY/oxMsQpQns+Fx
gH2FRruJ268TCGiHU4WAWHHKMI/tDQe4a2D5phmULjY6tvTGPZv9AfQxa7yxXQuP
pn45TmYgWUpiS3oe4cBsVepBqYabckmoRu9ArDckqDb+vRRnD6KvgDQOKgjHKfmL
OAeoQfUTGOM963ADGMNiKvxOxc6fiZv+Dafple3DIeeZYp0OyGnY3ZdBxujPdb3i
Btak2+7/p843a5/5uKIeVFMEh08ldeyGif0vzw3/0w0=
`pragma protect end_protected
