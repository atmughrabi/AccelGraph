// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FcmcYU7ILdNV5hdPWLfhbh0tMPagvFdAFkL641LXRQ5AgqxI2gEiet9jXN1N9lGn
k0LO4wjjbfFfHAz4JYnwovGXVxXi92pL+5wLIKLk0B0/soMrG2b8ppXbb2vaGwNy
kKxICPat9g+0O8HhGiuWULT6uYNujmAd0jJhiILklV0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5328)
6FtXZoK8unBrBr9w8/d+1cXp7Bl8WSHJBSF3rN31NeMHvPo6AxboAaxJ+iymjZCw
zVtmPy01EHXqTiHYq3cNSixUby9GZYL5DqlppYI+XCdp16blYhhisByT2tUp7xOY
pqn9Hqz6wk9sf8jlCwHffd3a2/X0g1uJbNb8l8u06r8Tq4yAvIHPAuHsWTWXZpxS
SHlHJaNr2uiYvNqPMHoDat0h88l9wzVBjKC1y2CIZNijrDYne2i5JXc1sQxlt3ER
Rh74O6+0bUwy1SJ+r/91nVKcjvmV2R2972mhoGC0nltsBFp2esm+XkkIV+CA1wrd
MoE+8jeFU7A6d+Q2xrLkSLDFYy3B5GQjP0UCjeDe0G4gws6hD0TyvKFBDIfV67X/
fCbhIGkif+TKWa4M6cGorrnTVcQZp56VQqQ7NC5BTdks/Kk8PzdG2tLm5tEMw5Gt
rDNCd2S2LpMRqJ08rTwN35oBuJwSo7aGN7CIpQ9MIEATZCsGQdhKeeOO5PEBj6nx
t1q5CPZdkarLrjCeikHZs5ZFhbCTNtvpXwQzxMq0g6TKqPa13l39mq0E7Cvj+vu1
hojYT42LEC7A1kgkfb5Dbx8BZyvEU0oYUXXtPHcMYTENlLEEVflxPIeHE/H+Zs3D
6O/CAeM52Mntpqw6lDhZs2xYvIpL8lLvLZDf5euC++HGG+7IyGhWE9EgK1THwno0
JyJjKlVOxrTr9Bha2xchbnD/vVR7Cn4yv1dSoqgOrrlw4ESwqTsQ7xKbGmeK8yE/
7nW+V8WzQo/QAdNVIEt0pj2Uh+HDyoq/B6d7qmEgbSgULf8ynRNa1RFrikG+pt23
twb+yzmU/fdexOEQ1Q/LQrJ/NFUQ6Plfkzkss3SPSP3PawNVqKnzsByRTVaBascB
It0ftosCBb84K6XdPO3YFEFzbkJxYeIFFCk/DV87tuaRaJ3MQVOJJXUM2n2EiQDT
zPBxerXXDgMuilpGKSo/AjoBzlJ7qX7ofGdQQJDmA617R3dbQa69BGMly2DGCwyz
WmlhlF9OLtBNN+0hlAu+syaDXwIZgo/sL2tRvNGh9YAmpcAKGkop119drBjDG4C5
Gq64t1a+YStemKg4//CfroqmYQ3eMhxaQ4Dif0VTFJrDKJ9No9tLeEJ4bnRjXfCl
H1FWc862O9XAwMn6XYw9pteiqm+bhO/cIUguo/7ZgNo5XERmF2pY17vkzXh/3py8
kphvxV2Svo+upBdADLqeu5o37ApJaIlIwzBLPY5uqT+XO/Jy+vnwCMJVBwFbX8Is
i/lGj7b8uNiRX7m/l4CDvxVIA9vs/RDzeQ4PdEEtMDCRAQAJb/ReqhMA3H8ZnfgI
2bQYltrzcGgx4fiHFz+2pKMPxDUHTbl8OBwwtwmeZwD9/Q0FR1qmXFwxs8UkBhnb
stxgzAaRXXJUFKL+zMXmocqEDyDTwpQuLIu17o1WvASgRbqN+tR5pGIiFxNmKKaD
+iiO4ld5xQ4CW+JOMEBSQWaZk6xsHvuk6NiVerUqerwvHS0Du/Wwsk2+R/A0TN8+
NlFhuty9gVsVoffO340VPe37BVAs7kTGCeqdD93AGdJRZDEYpwRceGw8Vq+yhtC6
GahUEVrowf9UrbXdxOFPKcErGqMKSK0cCezOp9d1GFViNu4ANXj1LZ7rQxdmSO2G
ykPfAYW1r5P997VwbcRznn9w8s/8GhL2xUhdD19S2ILDzq2MM7FMg3Wgw9YIjD2q
H/lIHKd1HRkQO6nkO8c5Z5LGCOS+FHLSPqOuiMsMUTuVjJfaVqy1LY+QKb+sVPnE
ATnH5YH4mS8K/7Nz+ucTX94q7fvUpDIk5+EGxi/E5PtjdC9AvmGvZyyGcb09HtHT
nzGbJH2SjCYQpl8RiPcsbJcWyxwpS5hPKKNfAH7grHcJOa6wLG8G6vG5QF7gl96C
2odG4mV5qA1OxiecUpIdD1G7vRfk+6EnIXJXCtDx3Xi4EfX6foVzLGf5at4AHHu8
kZ9wm7jCf1sxT/h5f0xLyveeRFl9GjV3TCdImvRvPUkG2plk9OKpdTdTZmDI3XMl
3+e+5U93FEVTxhL4t6YHQQtonU0HtgsEdKFkyYKn0eg1rCcMNMJJTI7yIbivhi9r
jiCGn5DfQcfrngIYX+q3FVETMcOc0PwsJxgdIm7aNPRtgkUBhxw49uZY95hA7SqI
x8M+Z/gxgeSxpkQVhLXWwVSvqGPmXN5JDL1dG7YoFjlwViIje2In38YQ/UGO9pI6
hUADbePfRmHDWf7o+5wccjUgaRQAnqqkHWW0gUQgGuWccyLDlRd1ypm9WQISbaS5
aO8bilH8buxYcBYedpwxf7BgOT/GwglIG0gcWbbvQxgwH9h28t8VNLfFvEA1V1Z6
A2dQpoTbiSInP2w8JV3BI7yiqd+0NG6/f5/APEOnxN3ivPXHYi/MISLslo8DCdkE
V6hssYMsPKJogSkuZdUS5rvTebFE5lCsz28q71QCFfg9JGpFDJai4rMsLxXaGErc
7I+jCTIlmvjC6QONEd4wfhO2nRK2xG6UK1jobxjPQgFnN5UIshJn3W8r4lKfkM/F
51Ey3IdOWamuKGZx6mUbQezJfuB1gOg4xTU4R/MfdtoTh1HhuvwwQyFFBXixvBYp
166xPfim/8eNEauqbMkNuOC7aJzQx6vhAWgBT15mtEhdGDyJSGFIC5bS1J6RmIli
dJUKxSsEJj1iqKi43fAZhPbDKqEV7W3Jmci68i7GfOu1fblFsftug2CcDH6iYVTc
mH7FLXosCEU+PaCiECPhPf9nyYO406USDKAROpvhqgb77vTc6Nt4o891BC0khEfg
GVAsI2+5A9KwlyCELf3pBIdqNm8732vXfVV++UZNOej6pNrVhve9e8buNAGYz8rR
Hhqshjuzy1vlmzxEQm9dsoOLLhu5WGomQpdUtpmdwLoScQR3e/4543Pc6RgoZ/LW
TAqKhas5OMdzalTYc1l0i/YJyJU5C0wZl+nb6toUZFJ53KNoUZHmkgFs4x6ABxlC
4rtw0bRnXO2zzSdNRpTbjsomahiDEUN5fwIEY7gl2FTHtmzO6VxW/j9+D43b9VSC
v1OlpAcrdkZw92K4E1/rnrud4e2dHSYxn42Z7GxYm53+FOMXtOzf4pYkZAIyr9Nm
tLjRDxD3U3zduR2oDNautteKqWa90Db3TsOPoybWUnt/lhs6rFAS6OUi3eN+twQy
RZxUSG7god59E2hTL9II6kZWNXV3lZJhohKJXIay5WkcDRdpX+K4q1wrPjegbPjA
Us1tzTzWQlJABBZUVVlu/VpvadMS773c/XQwIoyHfEXia3QlfTv5w34XxZ/ffVG1
HTHsQui+FMNcGQqyKOVbi/Ij6SB9UsOuhHDRiOPjC9n9jvAqF5R4/V8HlsEuRapP
euTGu5h3e/pTMIGpBOA3rf8vER0lXLxn7xuTCFAvRR+nK9AdWPVPO73HBTq7JCXy
cfe4/4+iddOpSZu8j6LH5BWAofgagq1Z21H+aX8AVFLjpIWtCzmbYkal/OQOH9Tz
nMESqwofTMbiZOLS2+MwlVKAMpQBC5iXKfkFosjG3tfnc6w4ZH2dOztyY4sHGHJi
oQwtXGsl3av2IpJhuO6C3MbzjHXP625CmxRasqWYoDHuHMPGOO2XArqtbeHEw/PF
v1zeiJ5iV5WVCq+1rRxzJRXBhmSl7E2o2XqnZK+mIAv/PHLWfy0z+DGE3Oisi/m7
l5ihr+SYNBvsAxgHmgtQQsWd60va9kku4HfAccT6bhuXBjApIC/V5ziFqcjlXiOO
3lkqDS7OBJFStX8WH884Wtdx1CxhHI2MERoEBkB0qziF3HTzznNynaWc69f6lXX+
IhZrnKDDWtutZicmrAE7btEr7+rHb7OMoM+WdQz1gKDgpigPdWOgM3VCGjGJnnt9
gdp6fCVV9o8WJxPDYq8Ks/rUkqejrsv7PHhXOsQVM5vyfjD2NkZ4tWqqPI8ajCjC
Ntz2YCTCWpiggUIuDMZ2riOlGaL3Bh7NYfrcfJePlHlZGFlkVttU9kmCtW5YVWiF
oSn+tzmTPHjQkDeUgLkFatRij9bfOLXhQEJYgBhh0vWIMo4dbxn76ZFIsriY/T8c
rtwrX6joT7oyzAXIhNNOp6Hs4VaQ2n8mS9+/U4b/+uGm8C5s8R6W0w7gtdxmw2kY
fM+GV1h2opqfZ6S04sKpk6rC1khe630M34z4HZcGVzd3PyhLWsVURMwj+f/wH/Tu
Xs3i5zr6fGlNH7hCQX5gHWPrvYjCGtKUQMNLVQZ5lPdnBf/V4Ql1yeea+h7t8FPV
C3eZEkxPrPiO/wNKjsR292Kxk6LTjDuK/bCDrmHvL+WjjV6dcoIRFZgYR7vndp84
hPN1PzdHhKlaYN06Qwp3NNGpB7dMWPa/UnbeCkMl7hIF38b4CUxPL24hUH9SyeC2
BMszppaIM6VPOIHMJfl/EeVggVbRiqtx0/zVlvNof1NnI0hK0hinfkQMO+Peus42
20rwDRBlaAPoJErQQH0SlwqUpWjmDx3bT9mtEbOIXX0OF2pxlVn59atga5FF8Am4
L3rTK6OVJzEYREWfsLImgEO1otPzMNa1qLIL+1DTuCm7ZV09eBDfgmBvzPaf+ztP
HWxcV9egdoOVV33AAvw3mNe0wb1IuoXGe7NKmyE60VR2ufvp5gVcc/hen8qNwY11
qZ8kfBnpLkLsaRwdpc5VMNwbgdxpR70x+kYUmXGwmpYF9vVYXnsdLg/J3xQ6giUU
9rfVqFBI8NV2q0MLQsYoHAElMCSKum7ND3JNv201EW2W75jo8oEmW9qcNUGhB7yy
Jr9cMyq15Eiy/bz9tbLz4B9EQgJjvmqFmFp1xHAuxKbBZKUsQAAKsNWVOlCSf8lb
W5SR4zD/3Uuq/XYxXV8uxzOlHd6O80MWRigLOnsfFk8zPF+IExa5kcK7TKSKm3by
aTV+1kM29nx5kwO1yKkuZoPe9zQ5JPvdubWhlommGfrvJCfSY3EwUB+6hOPxUFoJ
RF5lX4l5B/fYjjc8BoehCuoub6uPGUWpZOrYpOmekcVoTfShWdXu5+p0ZUxKY6MU
opnMFJzmHRDxS8TQnbu8o1mMoR8q30ftGtpWhpj48uMmPMN6CmdQoUjSDg7UVhco
ANRrbtRA73J+0mHU5XF2jy+z4IksHKT9GmbimQDzajiPJ3Xo9//NT76SWPtW0Fvr
u8lpoH19blwZYrd+8AkeawsSLmOPOYhg9uQUD5hsGfmVhD6b3k+wF1JgWENN00uC
vcCFKODpoBVzkdWcbtu95Fyoh21IanJslpSs1oK793w9PhLN6yjhQsG73qK1iqOI
ou657y521MOX9uKAChtlVTedNRogrDn6ci1m/rw2H+Psh1PKjILO2Fq45Wu4jR/a
GfDEghYJKg1zQb0rBMrRFxbuNKi6QjeEYy1NsafblWOucThCRx29ejx4TxB9fLiL
qhcFWgmoVhw01seENqcHlq7fo1DVbLj7YtiNAC7xJZLahKZ3lbZZoIam+ytHtudI
ooyYmLUyNYrv5tILSSDjbse5re1sQDyxs/sKn3vXXyncNKolAJCtYpfmbRCersmy
GeiLX6///bfl1Zfkh0IsSibavdrCcxf6IcS9HtP39pO/UBiJ2Fc3TISuvmkxxyk3
NJLGa850GYBUHVi7wSBvDzOy92jHDKG7d+CWZQPuAatAe5OjWjiK7Y9TYqDLMMXh
dbdTux3NPpBEazOjWl+lvD//ZfTiu0S9Fq/3TDb1IC3z4sFI6lB38mvBXj+15w6F
6e/42kzfK7kiwGdqooEkI9141E2OYZwiohnN2fGBwPgD0FJVrzdp+st+Zo4qSf4B
reFz8va3LrKKyozIMHzODtZZEGTFcvzmnb1axT3wixNsWzUUkuQ5/tkseV4NlYPT
XQaR6UKGPoBAj4zU55BG1WWwj+J2Ahs6vdAM22Z7HSHUuKpIjXIr6FX6rnY0UDKg
cEn2BedFGV2kHKMaP5LyBkE9uEIWkGCh0jpB1zkyzAYkCKid0C+xbZguSmaT/c7/
sBty8QbCmfWx/u/oL13/UNm15R0JjVZKGAp7gxkkXdCW634ePQEM3HDkepUM3onS
Tro0yMQUjWwlcBQS9xI7PvO7nbjOk9y7qclczNClotgZu5SFVyVG7vcN4iAhyr7D
+zn17Hm2/yT/UPY1EmxPk+wv7TqvTQ6WkT18D9VHJJtoWaHXdZibgzDqhp85dBgw
EzaiRxw0iffVBbxULgr8VQSLMQ40geykn1c/YVu/6UVAQoikQPYY9AK6tmr0apJF
3zlWo0UCW42V/IV4Nsln5A2zT4NiT3mTaAaiKHdo90h8kSvxslBmdYavOoe3+iY2
AxQNNiImlI1CYzY7vSjKHOcRXOq4LaF6GLfLCRqXGI/zozPVqt6honeN8PM5KhyO
2rvy5msaTmlr0IgT50bjpQS1R4u0EARXC/9iOxOEYUEDBVduBKsdouAdFHRNsrF8
wUonuTgJVNTWKK5kqTq92beeRQcuhyfNQuclMEXGJOiqNRfr8MJvgyhfEGQGDnxj
UGlGDY36vEtxZ9IZHPgv1xxse0e5DijPHUYn4sEq9MYNy/nPPWqMYUz+QS7qlDCz
tgbrD0i4xXVR9eFFQWfQizS8IufdJcfXYhy+Tvfqows9FjSaBksQ9Pk0YrwkrKP0
dFQf7X0HBDPi35SgFC6c8O2GZICEDJFFhZDr8IeS+tfe882nJB4UacUKaMKi4yYu
V1QWXLbs+JJTyxOz4oByAuOP38ZOEVXSmPxr48nPZ2dpPzMAyd2IWkl6oHujMtu/
tCuJmjWzBGLC63bX0L7YDzO1NH4KVafsquqp64K8y4Klm4RRh3F7tn90Xeutuu7R
fAEd5gBjaH42koCUTrqwHpwfpaJMR/Hzw9pO87OVHnXsMATXiAbizHLdsfN2hixf
lgCqXzn0g0rb0NhTHTADYDAiZxDBzYBohFqzO4SWB/tX7GB3syWmBu3lFZB3sOac
GQ1lWZ6akHBpKcizq/9GJEmm2sx9VkaKMKaYrlYHmPuZD1gmcGJ5xdomd+UzGbXw
p2J93SCFre5aqhWy5n53JtQMjLAY4xR5PvwYU60CK58aeSq7gvWxKyBySFashzdd
`pragma protect end_protected
