// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QTNBCd5Cql1Sa4LErxzEFm6gV8eTTFVpgW058lSsDJ8TbDB/Xkdg9MuKx+vCEq/o
2I0+LgtWR5EwzOkg2CZxZAvoY021rdKOHZPt3KRUu3qXGzIiZrTfUy4qmX5b2i0X
QPxmXhL12iEDU2zS0qQxeJ2oI1CG6sHfRIaAmdeW6Ck=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8304)
n0Kh02M8J7MchwEGlSxADp8QUOjEO83u4jz5SYMAcQ3Xj8785pBPWJPy7aTW1LqE
aEHPBzCZP6LclB/cNsPkL7k1kZMw+ptm0P/UpfjQcM0fPoFhzqHElk0y0zHe4wXl
PZWzAK3ER0oElqVne/5CQRns6A+IyM071aiNz74vYXZgK6u9y9Pe2xah5RB9yJ8q
mMSTRdVvnqYIhbQB2EkU1umn7PRtkRdQgjInNnO0Y+ags7VJDN9cDIFifVNq6ood
lOucGqsRXTbgnS4lfDQsFk4AfmKrXYNM1jfyU1L4ahaRHcPPNoOEvLNd/rd1j8lI
7OjefiqFlSJF9sNSGbHbvfnmum1xB18RjB4X/A85kuUyC5zxLCqGX6U0wkcy4cMQ
sP0xyfbcvJmtWheGHtTCAcfLDQaF+fo/fTvwUSHyRFkTr4+CWbLWSpSIgVssfQeS
bOmfsdigFnwOYyfQowWrNpred2bhp1r4jgL6QAAlkPMu1b4u2TQEkJn0d//QWAZr
T5ZX2Cb2j3AYACy1+rkge8+P50aKfDPCn06SP4DE07oqLnInES5sIrCFyuOaNqUh
OfCfKdD47MRUBYAtOts8hWNlV1wyjUiv/MUP8rZeUTibXIxsvsn9+/XPR42xaDz8
StxoS2bCVio3tfUxDd9ub/9r0vxdUYkT09BQbArGuK1yZZL7q/glm48YsxJ4HlJ/
DHGDy7+H8forJbqyKUgCHiURgfO2nTb5ZV+95suaBDboS8os9KNVBUeUGS3DVw9m
po6HWzIdMOSTO0f/FtokvQiDdULDSUXOmMuqM9DW8Bk/skHU+pUfRgzEtjDq51XY
Z3zm5kwsRmAYjOVhmh0JT6emtcQQ/BpALQop5aw/Rcz0MOiIoIuXid1U117BFrER
DzUT/+cTqn+bY6j2Ybky22Sl1UfOIWc/7EVm4uh0HoVW01wy3y5NrMQ5siMM+RRP
yE3ynvIke03cgKL+bdljpfmyhbV0jpoEQRA7xbpehfpWgwpkIq2HFtPwvi7beLg6
WmuccQk/Jd/sU351aU67+7aoTIL8vgeXIEi+693TmXwsDuy7WF8RwDQp0Fekdk8w
5Xi1Gt1OJ9CMVB5hviySPWuGh7b5Z+47y6sekNM0Ft+y+7YtiQA623zvhuMdUdsu
uLWX7CF2BAH1cq5f/s5HFiesq6T4EbW/fYolXsoEbRSMrNJ4mV8EWq5kGE3LCWPV
90Ol7Z+Fx/I+t3kMYE4p2mOfHi2/BsFqvpEMVmGWdSwHho0Ah3ys4Er3EGNH/fqt
hbPvGqkz5uTSi0sR50C0yufLil57IEFf2gksbOm6JntVcz8HpHjqgrEWTC9Miu1Q
LNS59DA7BcDdDTh4pnqS5xOt5MhU4OhfItyOQ4wrhi+s1mQ10YrmPDYYh10sud3s
lPeAlaOlcEvzVXUuRt/Z7yjKuruhrOeQYj4smiPYDFBUu2jSMh7U0Xpyz9b+fSbl
3LoW7e44bNh1vkdtOsKW7rJMhCqiASHMsQYrqzbyWdtUbMmGJIyiIFyHQDKR2kgy
IDAILe0KYi9kJVdiu3CKuu+mQr8fpFH5Lcjs28dE0E90pOKODlPFSFjYqL5/sekO
541GTSWQV3SVnaBUnLLOC394wY0wRNkHqrJRzZYb9V9AHdqZKYHzkvWcxVXeWlAW
IEUL11Eim1nWWTwmRx3SCooTE4Ll3hlYXEtk/xWRBFtHcFjkO6rjZ3ACKZtAj2O/
xbajIqGub+iktIcx50ds9P3y2jd5bq2bgqdx9HiPWIhZIChkvIYQu9b8ukvcTrj9
ItZ6LM+zJIzZavDCdTZWRSHKWn/y2T7ggt4E/67Y5vJRwatjyWf3Z0tAO/t4mM0q
55WWAcYM2xABFE59mc7H1yWAE5UW9HUzJ8W6iJ98wg/+QHhVPj+uiTCdbhF6X4fY
/EgNE50oOagT3lAVQF/B4WvwYqoCk6WOpkJgem4sAThoaAqCHHvIQFwErhTF+d8s
w7H/ej7z1AySgAZDz4nW2U2W+ijeHcZFx1amooZPHlYHUbFyFh0UKNddtsjnFwjo
YK87/NpylMbkMDEEZnseuJ5H3b7ivJct/RcKM6bX4uE6hfkHA/+Zxl1YvUDaJtec
jcKGYvkY/T3by1AGMGxf/G1o4toguo6mH3sDhdRIBbHGaYe+GbdU/UkJc9xVU/po
FNO/MKAQ+DoJgKZ0iCRODiLMBfg0yRP/cxaMsPyd5ECvA5OlTMF8U9qhxBtMyeXF
0nrT28zEG/NgnwY3I1r1pNDAyDZ2yFtmTkZH2Icjx0ReDEZN9oKDDFM2A8A/tcYD
3LY+DExJ75lOSgKp7TFaYHBj4WpYbREvQBxWz43OrrCDn3CeTuJgKiZMx+KCZswa
WMhoy0fPYqWEs4lPaXpeT3bviwXtwA44aXo0gxObEAhnYTy0XdRjVzsgAGxvyE1F
WI+9MHXyilaxY/6BIWsDsUnEGt8BzPjf+MNBEGxC+Aos/oq2KqtSRFqx4DkkUGzo
5/INpJyFdUiu4ihGiY5p7OT9+sIvSeMzWjgOAuOdQo3dMuaDzYahpewgU6gVJO7R
f1B6ErRVgmoM1zN1NccuvZbyIVmf8E8Hl14GREWZVrpVrdc0+2VSk8aeDdVgaqRW
aZozxBR/zODYeqZLbfueGZmTBdJusvpjbrOugallkQ+zIXp4YQAhh4UUk4b4Mtty
EjhDhwy22rXbf5n9iLfxJhJ0jK+5cq4Mno6xFBTTXy8c8Q4ImnUpAwxxbktLKn+R
IEJrv09KX8pxJ71UYiLOoEz15FG6nDFQAcjJSeg5nN4RubKecUoNVFaYExckhV9J
HQhmREJ5W6oB38d6N3G6akGrOSroUGqOg1dezUrPRBP/7N9ISDTIuTsimdFLmAFp
87wGUQWMygADfzBL/Nh1IeBYN+8uL5PftyejgCgUqb8dDdZRuPV+mfIqHkt6AcL5
p47kepgNuOyBMhmtA2EP6sEFi2IdEcJSJ+bRwv51XyUFK8NGX9e2HGR9Kj2UZpJc
WEGOM3sgF6yt/fCYxvLN5nKGTZrJOTLlGSHDuJCtJyowKQucPONTZEXbcjFwvsHr
N7Tg8h6KJ0KLvxBB+AihubfuPseUEc57pXcQ4QOJg1htEoJ7KQl35LYVYT+9s0gZ
LlQLgwiUz/IvlugU4ISQz71Rlnt5XECvgpU52T/J5IkMD4JSm+EHWICFhXvuEuVG
nPnWu+Vn9QRNzCEIAgHVSwN6Oga5WU9u+0L0uh70mvUxFukwH0vx+KARiSbnUjdG
nyrOS7U3XRkEqIvJU2YFlxsVTzBsFLf+qw1uPMMakx/rF/OI0mHGon4Pqy6NYMzp
fF7S+xC0ioNqbSZQkCe2w4+OK80yBm6jlI46r92PH7fGxn2/rBBfnZdzgnw+AlPn
rzq+FqK4gjemRbMOn6YuRYnFN99i3AKZ3ioM7+UMNLtF7HWA7youpYmWgPJYsW8O
mM/Qze6iIpUiG+BZr0fsS0R/BQOqvShh8lL1wcc4z1tmLdJiARa3t0wzhLce8IsF
ZwBMMfR/3F81bFg3zsbIS8abnEhITAHNTdOrdTGEdWTR8HU7s2S7ZKgGodnsHDP4
IFfawnDuSqhGVRQC/nM0TFdDgNVVrQH4HCcO7F4nQZpSYgfT+BneCpeOt7nn+jql
4Wth3cTI0O2j31bQl71opGuph/zWqndhfR9SmDke1eFMQIzHZI2mGC6qVgPyEWzW
Px4Itu+F7CAFGRFzVaLPX19cTXzf9HrpjjJN1GgqbIaJd+saJYQiesSPW53Q55zH
dcDUeKT4kMvv4CplTE1ZjrY9++pf3OSCz48zKPNkHHmd6dMNPMfJ+CfYbHdEzZns
uFMrVisfB8Oy78RL8ERNVyA0gE/CgR5WDb4ap3sISmHSMCC99/6XwNsT8PsS0/VV
48o4e9t0usfU8yEddWTmcoYDITyraVSlMuc8Ak0n3xsErVd1XLX8icjpf/3GFasM
3SRH/UKnrsbJeJqVwtNC7hvzPB9W1mrM5a8e7QVsmk/NNTQigcH02YKMJETcmWjT
GPU0ZRmbAWyT9DI8O3Aav6DGGtNnGQhXJ/yBPe3a5CRRNsRcl2qa676vCmDsokUG
EGmfhv8d1XHPz/jOgWG0PHsPJKJtgbraZXoNqMrdJGMaS+L8cyeFlD7DHUnhbL/Z
5DHJjytJY7hkTbkF41vWaB71Hv+fYpMpxd0mHSR000pa2Z/Ri2TKLU2sCLoCNEK3
9rVt4vdNuOXWEK6cDDruTN9wtI1dQpVAy3QJ9pu7WPGa+6ts7ouwhEuObLoNdxnM
GVHWY3XKOf3VsgD/CVNu9iQkgcC2acDH4pwraiSuS2UHn8aUZwtsO5oBKALHGRMC
9yzHFwL94rtXBozbvTCxC8qEwoUSQkaOv4m3nvtXhWm1eUIHFbVqEfc+cxuQOhKW
heqVlhJ4rO1BuAqaibD11HEqXCXp8EEDvO0RjgqJwCce3JDWY2ezGjsDcHeb8xn4
OBeZjlFcxXvRdvGBDSYny3gdoKJycRllYvnOOX/YvX6UTYyWZi4tY350OoYwffgQ
ecmrFKBonezEHMJ4hyaSrqnMRMahFLx2sYZ7aO4IMC1yM3ykjPsZR4b/JOAjwTAb
4l8LfQ2jCN4493uyi0CmD28NyK/b6QzT8O57ZMVy2ZcX5Iy0BtqZXoMTKyuT6DzX
0iIBuwwkn3TKACDMF13ULnMz/K9N8D+3jN/+4dOrAuxIVsgD5fyJ2QB4EySbCtVE
fAlehrWywPZ7Sq0jDlJCxYTIxQpS3ClGkjjYMIKc8d7Qaq+PamGTIFbtv+G43ga4
hwwVaC6dDHhgR2e6WcpWn7JcnhXqVmB8ODL4TMdifoqAmtQePrIKTymzmA+kXjjg
T4slfECcEU9M3XjkYeFuR4EWB01RVO7YZE54oz9o6BVm5PX/C7dNwiyxMbwqKv9T
3SSsuNZz3U96AtI+Eb8aUeYIujhn8f/tplG1HD4BqSza7kZIrff2isbP3o63SNw8
VlMQ91lcLvpBucswmwo1xzuHNhEBi7/GQJF7kml3Qr7acL/EI1vCzCQb1xHst8XZ
YJya+ioQ2+Jl9KG4aGtUUf8pcfTDmgLvER54vsJgVvesyPvEeaIbDAW2KpfvyaQl
FW1RrtO3t5x7kte92A/0dwQJbeSQqAu4h9My1QqEGHsA9Gfqw51egSZnYhCWOmM2
vPHbumKFYzqxKAo2sgndPekmERa6QQJ/SSGgYH9nwvSCI8k0ujyZgZ6yJXbgAKtp
TL2qJQZ1kDVtzKR5QHlBRFpIhfWWuurBKqu2ZK/n4p9oKIpiFoKdeTZhRb/dr1kv
2R+U67XP+tcWm1eGMsYOhRBqhVwBJ4K3iupJomU+UYw45XxX6uKMr5XmZpZwrLle
b+yu+CPhXbpPn/Lbk4bel5rMtdCDwa7KFNWatk82QmLKXf9R/LNa+nKbf/2yQdMy
nz9yJ9YRfvHkM/t4Ud2Rt3GPRTNyJ39poVg1luQWetHgM1M6MflCUyaeenMAGI59
bUt+lwFayWs5AlzrZ4V+mRNI4nTX0Si13KzFTUD5DOXvE+lG4dmd+CpD5wt4oKUB
qta44agpFwL97t3mUt4KjcXp6R05fgJB1EIvSxoi9oHUHQT/hQUOaEs+XlypiqOu
GvKr70XqMdTALKI1KEYMsh+i/e8+fXm1scU82MRbr9il5J6DRiNYv4CZY9PI6aef
six7dCCNf7n8dDKhgIO/k1WaGEA8haUgYJopmFBACCouFR9GNNexsqznkkzLsaZy
oF/bVJdqMjSwC0b0O2tS3SiOVWSIX7CvOfDV5o2Yzdstp/n/ftA2UYFsUyIrstHC
aV1/7fuV9pHq7j/OzwIFgxu3+bfVApbZ6Q0eL9rlF/yYepry2/hvhsz5npsUgNbt
kHlSWnsWhCpjFW+pNDEn4R3+27XkCWsNvX5KODKUyqT46ioTzgKMil/ZjuJazg1K
p0rOaeGLMoQLjnCyc23BziltVYLQ27WSZTUUKO2J24w2AjGcvlLmIVk3mdY6/m33
ASZaF/BHRJKneZ5gOpjlXal71sH26y32ul7eo/hIfGGAmlxjsHx/8stgUdon1wyP
mXB6BgQSsxETh40sRq2ENTwqsvXxWRebiPADt2J37beVnhrxXZSXUiRscOda4oKN
gm3pnruXMeNbV61d+yCspAFhOIASG52v70zjHrEz4dLuIbi+OJG6l/7cXcp55CFK
RMn1TGn6mXZvCoVXCfXEkYz2lV9eapcemK+khqnxm0ctIjUgUO1byJh2Zbu94fRX
w7HX3PdueBCdwg8q9XI2CpcDKqbHC48kUPCNNFMqplllIDjLqHAJd4FkJOluFikE
03As+oucdIs1pXuZNIhFkfPAAa1xhdV0px8Bh/mGmfgKBS3YvsIYhYSLcbm304Nc
OyKYq5xnqEAau+yYjqLE9+y//wvCSuAF6MeHaxJchmK4TTU+HvIZ35ad3OAXF5Wf
Hft0enbxl81N65QO05Z7aXuHpnCuYAGWqkaI50FkH5FUeeCWly+wyXwocOdMJwiq
Dj3oj4Z6Z1ZvqEEPdf1+tdq/icLQrqzRyeNteM8ORnFaiYol+EYpQoBljsqhyJO+
oN32LdqMiWYIm4NGwEM84Th5p80LL672nI/vn7H8X3EQPWAowVCi3ecz+Cws+K2z
t4dyfcaVhcZEzTm3E0jR22omRX68IZEVOUTq/43AE2NsmgOD+oExHCvrIpERU+GW
A7zQcfesqXzvYhMGop3bZ7SebCbYr6/b8gCiRH7Shp26eEAu53vrT4ePeRCyu/mw
LsukLpBs4OcJkRSIS0ia5Q7XWvRtff7G07TVzfhEFU44H5otuIFuQ933QNHd7A2G
mAgKI5rwHPVpbAyMR3q5HlzHdACH//Cd756RKq+RHY+TmtV0oBrjwkBFUYo5lnXw
+kzWuhrsiS6VQQTLO0ILwsfalYIVB0nt/ZtkKuDQEduPbWia+tqY/gLmiTIMeALL
0l6UGZmsn7yRKOPeH047+kbqwfElb8lnlHi2Oz887hdX8wWClJMXlUCavcLqT98L
+wrKPB0JRhCatDAdHsenMeKQ8EgOWOu9xhMQiGuIPRhP8uaVFUquG0nb+EDetar3
9OXcJKByqkxpx2qeypJFBXMymPgTyXGD0QypfRqWuujrPSZkEGaQHcTB2vtv53wW
zx8P4PtSQcK8Eb3tDWEcu8bt55Fe/bWI9JkgYfcolgfX9M4yck7J57/IrFx16usC
vDwntqnTlak9CQRLxVLgJLJE9zIvLoZx3hCXH4fjh3OXhwPkHT4YduJRlxtBR/c2
WOln3qM9IhGY2mVzs5uToD3yCStlgZt8o0RHHkja3U+jqMHBP0rxaIAnmPS/553d
K7kymoaPyEPNcLL5UBjwMke3vnGIv5CbL2QXoOp+Y6p/ekZRpqCoZMhdGF/FBECz
fd8IfBrHGTBjjtQFoL3GFp7zFJtrIGsgb6J1jRKyonJUo8sAdmokrNi6SHd2ryHx
+FdHo0R3kqZy8nhZiTArhuovpJEEWba4ww8C8+hO0UkchkcHpAHQ6SWPz8+5yeu1
pZDeV7qDxGi5y5+LUeERWRuaDi2rAJu1adCzTW1v85uXwL0Skq9oSaxMPm8Da0nn
hp91bvDY6j8QGnDZRStt24MuWBUoxNI62tsIui89xk4BcgGb8na/sRsjq0ICQHRz
hb81Bllag6a8vq+HjYueIHP5jIwqDt512QOt/n3sAwfMDUKJ0n3kIyoGacXtFniJ
JXFzAH1eSwIJebpUKPR7AiymO75IQPGYyMF4+4myIjrLqJ/b2DlljYctGBchg3Ap
XETxSiRgwl3209VTGutXc4ONJyeSw1u4eExFmtMFE6swD/9yUjHyjUSIs2lYBJxQ
mpnAh8Z2EQv0GOnL3RoiUn4JfO3rktv2fA83cN2k2LX3ywWRU0k4xU3fQm1YpWIQ
Ax881PAGf47orgrFzhPikSBb0MzEoWqqcfpfQmf9o3ojt9fBg8Tmhd5a+dODo6+L
ZCbHxXPqUZZeuo4HxThjfsi7Dl19E/bea4REJLlRXHnCmEmy9mgMrCsQWs1svHTb
3cr8aTriqnCopXgIiD7YOzp9/4fUi3/1zSjSsD9TPz3fAvf/MEyA2UpH9p0AuTEn
eR4N0lOusptSU4FAgWq6IM+EZkODD1z2YOYcRKHKcub3Pj5khky2KMLdYbqHHtSD
8gN6Y9ZDUvQEM4/Txaf4BzwXiQYQi0szH+21Usg7vx/38CEeoE7bBAbJkAWCp3ng
56Tf1/bi4ksIJAY0qT4UtmxO1sVJ0wZVxPb71t9UlEyvtPNwn9fvg1XpU9xjjqoG
6C09AhHVd+RQtHGrLJg8MSdBJftp/Yb1dRzB7YURa4CuFL8Oot5nBiJaOxK5Z55r
uO2qVGP/ZGTmkzgXJO5aQybMIviR93r6qTx/NuXiWjAtaRR39xAONlop2zOQmCTV
fdImtmSO5zBJmNGmo26G2VF3R1tSWKUGmM1CC7Fmael/3TNx1NLnJoMPdl/U9yJv
zvHJjJrpUywgUrEzQnVOZzlbiCouOqsSFvR7wjWKBS2YIsc29oHojFyKKl+c/B70
VJj4boNhhvpMpKeoVy+gRGnuruBTtKp0TS9W/wOL1META+RW3TrbvwcMeGe6PnwG
EiBkpl5XTI4xRHx9Wnr60BzlpJK2ucEPGAriM8KXCmRIMeM0bNp/3Cg9n7sjAI0Y
z85zMTZ8+tza8XT3vgoAuIyP8sPe41ri1cLEC3dpDbwySdZWH9ayQvuh+aBksag4
/VeZoiEibLtJ9NcY6+TdMmMDo0Gw+UcHQ+QkPiA9w49Cid05EoTQAgRe8ZGVQvDV
EAmM6aIQqS++OVqlYQNpOK5ggaORGsho8900epxvuHXGAOsb4daQLPgYUagnal7t
h7dg2X13/zmJzUfEaTKT299ZPrVO5l33bdYzWICluqjpaO7la+gSna+MgpTTr90F
dsP9kwFl8ojUYPta+Pj+ors1t+jHJRYcuSkNVtdKot76hJRI1WoNaVk33ocVqUUz
/nQZXYeUQt6qMJEmj2gyLjjRdEQEMpNB4eZH4t1IhMUdz8jL2PoYW+hwrxQYTr0q
tfmk8HEgHjlnt8t9pAKCKlOt13ifcnv7qVp92GORRkhZMLTsViXoqgLzgfXU0GrP
UpXQGlMyTRLjZpzDtLm/Gonh6EQmQJFnVtL8MiWYkfvDnsDcH1CgkMFWUf7l/E9k
bKPNebcheClNpZfX7eTYFl6Xh2kEAMei+RBWb3T4jCqC1+j2aEhjEDi2scbnE1ks
PdFl5UkV6nOo90itC1AWm2felRymzZtPwDM284FiNs3CyVj8kWQHwR7MqzVmlcF0
uZcyY1E5boc57ylnvF9T+qVlulCw9Wr9s4kqATXCoQQ05fCGWuY/NiQ1hT2UJCIx
ICi6zkNle2iM90ArxSQZF50GKO0k3+UUrXyDQqwNEdi0vJhFSvpn68sYV1rMHiJN
5sxcbEwMbymZ4shvO8KICKNLhIGq5Hhe4CDnAcys0lEnxZuO7+wYvUBj7I5oNvfg
lB/9CzFCftkccucWQUbRXQlUvHJdQTq2SPKh73dG90JHtifLwX5GPv3ZckwoHo7W
jFwJRDT3wwzSUuP6kxb2sLBQTkMpBZnDZXh4pafOcAdpS/Fvk8ee5pxlt/Rh+Zgj
xcdFnuEI0WWcMB34NQ/T9+e+q26mgBCc/rDDDZS5EeGLG/YcPfVgtqOGop6iIWRA
szD+JEvOPvqNhpztVbenbRMbg41CBkbhXluf3T7nziKqgh6GytBN/OMTeCSR2EKr
RLXNPJtsf0KvP4aer13m8NT+Kkhs0slY3HKkandJDKaCzxUIdad0rWiPqeIlvFPI
6GZ9ujZo3h3ETzQabjZ8WC6LA/+fV64T1kF5z5n2Bnvv6AdUfQD3cI9/+vEyGU97
wqdWspN+GR2GwCXaO1CzmGRoDdsHWnfEYyu2qPe89coLfyHPfBqVtWnq0fX5M6CH
YL+qoMzMHGYG8eIPoiVDwhzGq8ajgI9dNE9k3OJTVvCgfO6aPBN+DzdBu3fsglj8
LlTK/f3SQQPQJdKbxlWDNdkjdKZZyeKq7ai+tFpZQcq50ezNtrY005OABcjCbHzN
Qt+8rEtmzdyR+UxlQE2pzMezYF5xyVEKs8JAksEmXBvv9U+AF7TLNf/r/msxaeZh
3U2u7MM8bekNruJxukqULY2EWwg2+EZi1sAUoeKVJyP8S6j8gB1RlhAArwPvhU3u
QCRHYpksMIHcjf4xDvrYuYtNTWVclI2gM6lcOoUvKIB06ihVNa8ub6WX5LOweEvH
a5cYDJiOW53Was5fqkzgp7cI3dP1vFXvQxheD4N0PHIgmiP9VUvRyP/ioCvA8S2w
vC8TVcgYYLjsHGcDCTX6VQAwSTMob+CVB99eiVdfzXuFQ8OY2a6oEWrG/POyWkB4
oxNZJkchCi2ykP0JTlq90b+xr/iI3P7FQIsG1PLn0upW0GWxhV/OYWDwWDYrHy6q
zpFIy9lrsM6Y9HQ9UDgCn2LuaHH9e+g7TKw8eLXTevs7KU1pAoozvzNVGejuxH60
X4TlR+EZ3lCo3Of2O+yBhlqWaQuhrg4XIzta1mSJAi/Ab90ZdJYnTHeqjOUPHlBo
8OBD3gFuryfAC0rdgqLOPe2teU8UOQOUTZjieYJn5RKuaHYYZPahn/g6OhvsR1Hh
Pu/Q6N4alqdiEc2yMB1JM+fPET0rnj+Qb1idVbOL0YQMyUf79gBjy43P0/55skAx
EFvUZlDdBcopO+vjW1Y5Yekh4IcoF4c2d9QipgUXw9yvFE7sU49YZNMO6oP+WlnE
Ga8MEC5wQg9zWGE/vWLOdz5d1T0FrNyRNOORcwGKWk+wGeAEFDcE+iZ1Ugh0tWmU
MPtHck8hsMfZEwQYqoYdbwiUiv2UtYpy6kKMsxAPGLd5ZyqefUvcZjAltUfKoLk/
+Y4MPK8ua1IjYeMEXzVO266r3StWVaFwY0gE1IMCx7dpDwSCZ01aOXobYvG8JyGa
kFXyrjpwH2pvC9ql/x5xu9iaivFP/vrTkd1swb42ful4PjkMN2cEleqPo/8+edHX
`pragma protect end_protected
