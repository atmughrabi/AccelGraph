// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
UQkr7Qk3ZRtJZRJ//q18orPzm5W3zfKSDHiFubQQGgavD5Lb/mqXafh5zJ/Z8h19
a1EmLWQg/NiDrWSUBwMTnwIaJgX8l4nGiWZOiyvPLM3EQpRdZut4Z00IpFc6xXKn
MIAhzRylge6T/cg1bhgeQUAoSrVKUSoRPgDTChtLcOzkdTJiaNqg6w==
//pragma protect end_key_block
//pragma protect digest_block
qnD9SmhG0HtuIIRKUH6LDEOEntI=
//pragma protect end_digest_block
//pragma protect data_block
vHPafStLHdPHVhj1A3L0gab6jh+lA5bNUHhm4uya5p7QmWjkPTjuswFjrTgm0v6h
sKgzg3hMtzG/4u20AWDZhl57Q0RPe8xRBQgGKSfshXHdde9kuT0ynn2S2fwpp9wS
Vzvi+1b7YITEmr1nunfNe3pY9k41zafEPXKyHphcNpIrA01HRdQlWHNeAS5+EE82
XNwycEdkKq2jUfraI+kfuRYdmUxaqLcUY147+c52hN/nJ6DfzRgeDb7+XpvvYarT
xWHpdSxWF4C4BMw49c8/Ovy+XcBhKp7fFoMRwHhKfUNWu0Cb8140nKdyU1SpDz9k
eGeFoTdixBeLMkbl5XX0Qo3Hz66/E0TIZd5uSUwN50S7V6SE6fsR4SBgljQ5JRkJ
p9bH3CLJEbKNOfT9iDCjBPt1eZa08igPLybrE1Vkm8dc0W1OBBigcT/5oR0ZVx9b
KmC6coQUd3HXJgozp6Ws/h1qiNpMCZTqBJrBawWwGixKeKyBEAAsV4jiAIsISDT4
pOfcqauHDthc5VRyvPnsi3NgopHfhXiZlSFIz/ovacm0zbQAyLXVdLk+kj0buUEB
eGCoVBQG0MDTuvaSj0m0h1Oz0ak9zSOkDK5QkL/K6oD9Vc2WrFmvlPsFE18e6h0h
HJwe7xTWz6JKURfaxT+Iu+sSOpzryql7XAraiC8n0GtY688cl7MvMOhVdNrRHG/w
zAMn3HseIlNNumowfcyX8W3GwLKveNYq+G5yM4q26ASZBvleHVOG606Li85fLpI0
R/RaaxQGC3YHXJ94KJroFxVUKTsROSm5B/ezRUWRZwyT6CWmDCf4j2ZzqD3mslcH
Gw/9YPwmDEuAWTSGaPTjRIOtimEEyglwu2SNC1vc/n92Mv1Uwm6vKDUNYO9bgvkP
GVpxxhoOA9E0BwwYKC5LNKL0AtV/YHHrR80kiJi72Tdo1xGebK5kR1/VIIGll1F2
xPLj/Tvg6zFaVxZ2EKiwh2pJkmb23+1KKN/c9qYQjWgBRYA9t+Oc5khVfBHVSy6B
jXueZR8jjpXPTge1bg+WPkURKJRQrl9RPqHEGFufOYxYrFKIeIYIyjIVx0YFOmGa
M8VtJi0MnD+VcCkqJWM1luaSO3UTDlPC1MTUhCN0rOB+2v8EYqdu16UUtjicwsGg
uZEfalaO9d58ACed0ECvYRuZx/HkoHyD1d4XrDDYxwctbAzGOAJ8lPSmF0Lq5ZXP
MvxzwUZxmBad1D36bO2uhaXBbQDBnVQqpOZ7WjuyFO0CSj+b5MMaBaWE4elkhJBL
xksTj86KGIhHRpoVA7yPuczG+Aw/H9ikr2ArQ6h++oM1uQoLnRhrulC/Oim28bQd
k7H/R0T8TUaOkkQm2aOQ5ySNOiqDUZZYc5XAGlBncPmhOlMysTsSjEG/alLzZ8tr
AUP66qPzxgKIO9z9kD0onbme2oe6Myj+oGvaqCLiwkaFMK6lpbmsm7AxE9xc4B/O
jGPlAUcNSIXe6/0KepgTZe/r8s/s37SpBM58yJicoNIijjg6L65DJLYDyVAs4hRR
OGNbxhmdeOoFVVYrcgW9q+4bh5qJLkww879aikBUJfK40bxHzs5YsW/eAPPwIc5L
BvZOkWBwA7ymkUX1Z74mNqMPaK8K2bmzRod1ZFgUoeDuC/BHeX775d4+/1v8UdZ3
889la5WbTjtPJA732dY0GoZTQuKMNQFpDyDWF5/XWfPlLBUfwUAzIQ9ykVOQ3eql
8RG4O/BuY6GmW8c/1qlsjV8+7k5w9Fva6yZgE9vwR+lXlYtJxBA1WjcRCapmzKr2
Nq++IrpZ4phveCl98qp3DotYnj82nmQ2HrxrTE76rzYoGIoXD3qHqK5FRvlCCAPW
k0s5HhU4D0GzFl3rdEgbH0XhoQSfdUg9yVCJNLs6HuUTQXZ5luBTi7b2xMkXPlnT
BgQWcbqETt5NGkdj6uXnVVyDsl6IhmY014vVBCoq+YKYenj2p7/ZSjH8n2FxJDb7
hfvADJdvgnZfVkAaP0tp6kzfRUv6Bt2LO4KFg9JE5TXztjPHDX6DD72u9Pn2mQLq
C4M15Sil5/58QUE2Yw0o1PtKV1ophahpHI/K6HqMHdhYaI+MmzjZ0Zj5LjYrnG6F
uGZZkwJuBctLUpXVExlmn/h2YOjN0jug34BcZmNCUw3cf85Tf9GmA9oE6jWYNUy4
QbcXNbBFTHkR5TxgKnhDcCRnmDYS1RKSzcUlcO+NofZaRUQ544TMfY3VNFclXJLh
DtSu5GKPVYzbZih+xt1Oz3FDa6OQt/1PY9y3r4zlYgJOLC7iUBw1q10MYadWTHQs
DWAVpfYaElreG+BoVjJV41bB935NYs0n+NQApnGPfASiNYuxV1L3wxs5fmnJA/Zj
6k45/ZX4LRz0Gs7jIaEoi9hHhmJlpE2oc872iM+vPyiIfB5UPKwxhqWVKk6JUWXU
jQnaqST2mm8bflT0E551vwARbNcxa89Lv1oSpWasP1OVraZyGsmXGD0XEBuEunYf
kW5HLtuJul5I0IoynBso2xN4bU25yydfb0FxYGW5R3/F4QoKqKMMGd3lBILR1Tjd
TgKmnWuTbrVClA1BzGk/OMWXVvOE0baBCQ5xt2hvRz7s1fVqplE7I9MGPdMSJDU3
lGirVb4b343tA5uunFe+mj/PCWh5y+2+UwYDTk5lI4hMRGwgdLZCxLStANSHWi7h
Vm3etKKEQONYgIeaqN2qQe/md0BAH/4LroGYkL0tRkicA0Hnv5zGjUk2Yt2xhzVH
HqvsK7n36P+aH508ju+96kNCTSck5vJBLBAI2L+LU8V8xDeVHbUWn/2NDoHJ20d2
S0ivTvH+WryUrmvY7ny0g13HV8GS0Fq3RFg7AtZpgz0Bh2Jr/q8MAThq/LhtwUfK
A1ZE9DKumrBcrAalDAiyyx8A7j8+hI3bPYX+7beDySnDLr6lcuydX/I3uk3WpAzq
RUQSFudrXEd35NUPPX5QdhERDgIeibLHqJ+z7EP4HfgshmIMDB6XGWxQE2HSUgTD
BUmRq8MRlntDhoP82T/t4KJHYCMbZxahyxniYDIuh/ujuwEIxIRRH6Kns/SOmAMj
3mFwxcV/67PKJwJpSCc/P2P+N6JrR97DVWXYgqvux1rAQzWZ42M1NMCMQSog2Ojq
i43MZrKXFvGgMbnPPBbmiRbaHyPyNWFSihAnsrvqzigwYvDEDA6tNg2J/NMJA47v
eZlcR5IBi8vZBC/Do0OtmvXOl5/HOzb2EK/7xAilOV+Fc1E+oIzwzGb4fV58y5/r
ejxGioqZEu9eoSN1hQ8evnJpmviz3XrS6HUUk9R79TeRgk03HC80+OnJ/0R8nZTM
8HcrYDTVxTgzSSB/Ut1W/xqmc5v0SmX7lcGZovxcapIZF+FVqyS9UeEO19V8DYI7
IxcAkZUNMqm6C8nTxrArmvVg3dLnHk6Eyx/gceTPEG+nx9ZaNzTT1J5eXIlPxeDW
N79w13Lmr/IjXhOCynqyLfQaylDiV2Ws1okSrVGYR36l460QafPeMcog3ur3pbZv
kLITblFhYJ4nu1UFEn7ALMngVYBo1isIu5rAKQPBmsE4rSbjIiQfJXcWgHwUkn25
4G5P3tmCvKeihsrMirU1KIrKRxmZ1trKtajce5V7BeVVVz5cgy/f8bZ/YjgVn332
A3qkmjQFzGKK6kqOD62Ti0oP3PfN0ZmBrrcfriXs4Mw42Zs9d56mIFyn7Jq3ha3F
Exi66NYJFSwG9yU4rXQGSQsew+38mWrTJnxG0FZ5FzkRjeqLXrOkgK0ZtpmdmVNf
cv7qLS85047RBBzZqkn/gtKXwnXUFuiawzQcvrKFXrcmZMk7NL52Sw8TJx8zdc6j
hw8Ni0mx1o40ex93UPCONWKxbkvQLAlnJxY6UQU4x4q1eneW8Gbwm2bOqNBNb3ES
WSqA9aGZbvF6Vi8XYukrC0Id1/dNrH+yubuTvfUOfx9WJOh+zCkjhnv3cAH3NTr3
f8dVQYL8UuTQQwyDIGbHkhK0dgq9HY6n18pvaIoBS7GUUos4PRYZa+aTWyrhBnRP
kNdI1RnRtFPqrClqdaUyqCLjiAuCbu9+ds4mc/eSFmTXpOgMD8KW4yrQAnAnqG1+
xIqt0TCII8mRCmwmCGzVi0A5C3JkBy0nhfSO/c73Cox17wqLLLZ7CRM4h/dwegIH
1En1n8zbOtbbz3YmBK5V8UYfpqBIfHSQl3+b+Fnc3V+Km6Ow2BJ9VTkIUufd/CSX
IyzjbO28bdaVFdAFRx8ol8oZyuGUB9mMz0t48GuJkYMKVw04qBm+OMHzP1R2CaAo
svrxHINRZxT+HDDyHmbtr9+bhmXy+I7Olud9SOpKO1JayA0u2q/E4QVABt5DI591
bVIG1e9CPU/xU3Ic+XWbA7COMe1QIIxroi3onjnBbsuLaiURoCypM5KkbFcLfh89
EKhp0SJZuzG3W0rtbgNzh3ozbIpn2FWLapLjFKu6u3vOZjcv4C02MpPJTm5INpwu
TGi/079wTocCJS5nZOWOIdYzMkEmUWOoBW4cCcqpPxyMJ18jhKWgFNcHKSXdyPEQ
d5vh6zyUkmjvecnnmW+7yETb5+Vmjh8ip5VjHgOmyzg6bY3YTrnZWzPuTlqEv7Og
OjG/RAtVGGOZRjyvXJzLLemifwHBbQgtgsVBpvcgIkJs2Z/Pc0k6uWcmICZsfiIl
Qkxds8z4RCoekZgBN8BDEaWl+q5fOivgo8CvyBkVomsbb1a9FAgeG2Dbg9j6VsAb
+goHqiDdC2iFb9evYkixvhzY0GUqGoBxW3D1SDXWsU9kBPifiryzRhyOLrwI1lzJ
5xRP8I4uTFWOtgMO13OGrLccW36wc6poQ0wYR7al6QYP9KK0tYslcmiD1W5zcmPv
K7ZbbtMAANvoiIvsgFRRr2NxlAvUW42VHUtKkO7CSkE9Zmw4NYKljK1qNRh1hBvo
gLKQ6GatPccac7BqafHPNI64l5W4FlVeorljsfJUU8wrqrFHIt4ZrqKG+L3QiMeR
HgD0DsVx3zlrsSoDtAmanJrX52dxrTf99j4OPrhFuaN8avXFQ6Y6B926bqEaKm+X
Uw1iQTCizkvcagT5hWscgnG7tYlhDVBea4lDq/H2gKX64HivzIAqgwfJayQ5IpmI
sadfksYp2WcIVrYpdgd8l/kGtJYimCNdE1kVT8S5FWkqK8KVp3mt56KcbSV8byVW
W7kMeObcXU34OLLUP3mgrg1dOSJybhjALD3I90Hpu2HEsU/BBrYvpFQ9ecUpYpzk
RNOtj7XsxZcMGX0TV8hZ3c5sYEm6EwJIFWC8H3zVRApf3AS/ITFEZgPpaDgN5F2z
PTTnJ6RA4kIEzOXIqTnjGB4UtF3XeiewPF2wWkRH/+zoOTPMRmfwnzUhix6Jbpoh
biGNwyYjnH7+WIcuZoh/l6jNPEUskcmQVsLd7k+5c5uC6fNil3Cczn2vdeNSOJZg
7nhY0n+AhfSEHzEiJKzVJ87BTuzaeQbP8AetCns3eE1FMuS1t8WYqdXO2xf2yetv
RzDucwBXV/+J0cTnWqTTVllfPpyE54wxfYdnviXFbtKCjOtzR2k3o2at++bpYirc
qEAZMYgRtKvkl+9h/cdeTJG0ARUdcdfKahUOq1N7RvPiQhfU+kLKqTC5TiU0pmL/
D8qVBxmjM2iA4Q7X4GhQtOhGxSTHvK2y7ecnAvTE3ZOccjM2NGJqoZz1DC/FnVJu
ENhnBi3EKW1OF41ZOE83QMDqSY3K4Us2JqSqTdh0M99v8hjrbfiBs8Ys2yWhJn/G
X3kSwUDATt2VWo6SLrl7HhX2qjJYgX3gEozTbJwRcBhRQNigy2zXZrdVOAQFvxxq
uFw88UvwrbbAcR8gxRxMTSzeT1hRTShG+Ym67F2Xc5W5RGhL6J7bSiIMGhwIuikQ
iBJ2q31A+oiHiR4cYBys7qTSGA7gPAWskAbOGDEgkvDOI9j+Zc89kw0wy5Ij3o1f
sgABgfjKx9isBNw5oCCgTgLXdo4wF69sKlrOF0gh2WuDZRdAjY93EKaTVuUDTBlk
PGT1Pg+HfhN3kRI5ZWrYDnHnALgDMb0B6Ptegx4/KDfmjKU59o5GdYyB7hj6CHyF
h1/HOmcKVV/tpDrKiaMaMEYB1oYhzhm+gryDGNRSx3oYr3KqL2OXsFOOWTtk8CeV
WBVHih75mhL0Emh5xaNASW6JSY2gYpz4Z9nDimV3ODdMGWbB+Kveq/XzCWHvxfut
jLJMQJqrZ/Rs1qLgIBHMOz+3N1/khPYrkDaqsOvgtb8GgFBJRlgzRRPIZaSsIsjJ
OP4dMSa16Ke4/8/0vFFSvc7RcDUEJkspLt6HnMTobQVjNJMy4RbpvI6JCxzp0Fzl
JKHpNJjjApQqF8rUyW331aPEDMrbnR86SDw0AKiTHDzmyzf5XLXpG5B9fGzng9uM
akXt9ZxUinRxeFQ/naqpfrcpQ3p4fMHGOrk+Gmu/lDzrXOVXhU1Hv1pHt0PdZxFW
71sYpH7ipKHQyT8XodvX/91q2EeiRnjq8oKdD6XZqYDOTCcxeg8OJRps797RLxl/
K9EUP16nvwUatmqRTszxxs/3soZZZbsWxPYWo6DO/5r7FrFTtQipI+mrV3kMDkNa
VgjhPLGwwq8O6nx/PX78uSAKKU1I65jqpOBS1qm9zcD9dhrcnRWIu3ZsHhovDcgq
Q+UOrlX7El40q5GWIX3xQT4hVdxZnJa6bIPSexbrpoXrD1V1PmnoIRKH84uohO/O
qo++To+nwBPT/0F96qPvRQ2yW2l3tlHojK6HRDxQiniLftipN7fNShar+XEMUzzK
bcvGMKJqp53P0AVAaeEa+knqnwz2VRnE2dUVS4IURHUh7cOzfV7g2JQfW99l2zzT
j2iijlnrpSb0FRjBF/iM8Gxb1/cTZXxXM0ft6iG5va1b2vDoWge6Lqnlxusy7fwX
BUo6TXWGLsRvRFzDzRXQamshSHDt7gAScukIma7B/PshHAkTPC+r2AtXRn7N/OPN
sIlckzlmE5mX4O+7iKZDhAJ/77VBr1ZKjQ2oLXaGCowhcK0HEGZEJQ1WDhBlizHu
A0T09FRXd1TM2f/UjQrKYsr0xBtYbBHw7hjI52Qw/xjnmphngkuK6OtjyGJxYkMW
o0spuj1dModxRPBIM33CYjDO4pObdGUUKhVRBwCZNnujJDgXLS/Cv5yyBBXB9wSp
RVznVTzjT40ANxpyCXgk9bYcYhGbU2eyKrqXIJKgcpimiwic99IFmUnxrTaHeFZz
ScalI2TbhfhkN8/JKTA355GPqnxJqJSvO0Bkj51vaah0InnVvOYVrfuLeFYUfstF
UMHX440/fy5g6OUsroe5mR3JxMD9qzMLxSOiYnwk+JEwCEFhhFGq/exuLeOfmZqi
zRphecNJyYQPCpI6ZcplKIgn/Tw4hq9/c4TgCf24BZbnvoTnEdQFFOxWp+kqHV9a
Iql7c6X849XiI71eI1+33orxFG7kPqAe6/ABxrMI7pwz8KdXLvSq5lqCudYXFaPp
pU1CZCoz/o+9qJrQ96VInkZ6xA1G5sl1m1GM6Q2vbflWqXZSHchXBUp1M3ftnyOS
dnqj687r0JDfauHbUoqAeLHVL6qy1GlLddocT7U5ojzn5tCdgLvPdeCco5/9NNgf
thG0SHua667fJ+E5srpNmXmJHigcUUFYCtLBfHHKIIKcjAgS4AwoMuwBVTMOEq+v
aBHWHCHOl620iXdZ7xt3Pzp7ZPnw7S4LHDfVy56BUIFEdARiz24NMQfhyGW9u958
XtJw5ZaKbsvrGJpjSPbS7j4PbRiBh9jARCD51/hiZvMfmewvdJFf8h50jreKuLzi
gHAkmTCiBhe2sHZGcNW15nlf4wORYJpmr3lAxIEmnAULtCm2T1yx9Kx1lbTElJaI
sv2WoCAWeTrHcQKNC4ItdaJN+AbYqtMpsPHPOR+yxWX/vFMmvhGfharzICMzpwqc
i35Gf+lyYKeNJt1LOtMLX1n7OKIXIDwoxlWe3C/xUrLWC7Wtvj5PRFgJYUjnfJq3
wKcQna3zokb47nXtIgofQqMojcR0gHtv/PgDnyIn3fhaYozM9cGjqMw0v12FvA1i
QDEhjWpEMyWX4Pr6XPKOszZ0QHsxDlvUPDXFvRYIrC8Lq4+JfDRH8VCZzO/CacYK
HixASS7rzog5ouaqJbLid6gMYLeft6rbdmMS1AWLMxMbeJ6+0BSQfD0bo323+/4G
rmI+RIfPDQ8NDfMo//XtxVxrgm0JvynAgLrzwOyfrmOX7jBiL/66PejWWVDEIiDY
vZYXz3BFp2fuiZP7fj1ZPNpmXH4R3EL/EWjgrh2iDj/iAQv1i6Ar8ag6O2pDqkaf
G7uFQPXw69W0lPEuazFll3uMRFweRk+pgRMJSc/exk9NGTC8ERW//VAocVjgVcPl
zwaX+wOW0kkd2BnNJjPNf28+vys/S3XvpDQO3uZEaJZdfqCJVnzYu/yvXIhBXxan
Q/g3GxiqCx7yolOXCqWXJyF+W7Gpvuskm3PTZVwBRyYs7X+SYp32IkR/ClocZwj7
AsZCKd/vco768dNEkz6yhEIdNdlqP3Ak4LfxWfDpNV7GyhqdoKRes0JGsHdMSP+l
7+efvKKx0lPbeXIxHO97CGCm2Qh6oMLuJRMjJbrBk1K+R2yJUGBikscRQtv9GWlt
xZ1YArSPArrFZc55/E81YtZwkgw/Cg1Y3mdle4+A5B7lrlvjNR8E2Prpkup+lsF/
N22OKJadS0Cr/CXdK0tito8BwUn+NbC09z1ufZQThq3uo9kbjw/T+ssWItELlH+f
E/zSAMk5TJnAADbsXAfnlrfuMl0amhTix55PQbiC7G+wlQa/6Cavb7cCNTWtWIc9
JvE/yT1mfWUYIbda82NV6kPFSjvePMgcvYfrM1OYJ9jOYCzql7s6eS8slBGWEMBV
DwmLnepqD40mWGR4kr71bF6QVaIINFgX3QGqsDXfJ2rKUWlBSbQSCPLth1B0MsYq
w7X76uoimt9XdgSjjtZL2BUTLVKJd2pSuz2O+VxQaxnMTqVwkiVobEVM6jto56SG
wlPETH1BFbyMrOGvcuIDnctI+C3vK79EVda/X0pW9zs8LewW228SA3ldL3Wo0lxv
p5t/BW+6Yb91jcZpi2KB5girQ/nDt+MPSbr04ENRVs7TrPp52/23O+QLiYkjq0Un
kouSEChS82ou3XQY52R4J8YcaHA89NxIOoZmOkmxs7juMOVH3mn1qd9JG40KlNE3
DDl5kbr3uqP6sHZPqrSU7TZsUHivQM5kF7NPEqzrc59TtK7N/xggFNOPzD8F7Sly
cwjfBDtIQD5p6oWGqp/z1tnhVONbvSIKIKR6Fbb9ZlaCpouwEg4C6XwVWS++W/7g
Crksi+Z4Rx2zV8+pmnYvbeZ7ulwkm65GAlnHiPWI8ojUtMJUkj2hfi1HbUHD2rUF
ZR9DqpAryr/4unNST6ohzZQRouPDFRteu9GYk6Qy8e8jUIm4jy05Aa0FuHQlHIjv
a5FutHAwQHbZLdClJXfFS8cGwXj7ZgCLd8GscUz8tCzbxOc1ckRoa5YfZmWbsiLz
PCGEy4jTZfCLy2atRli/7ZaMyTxFD8zKZLNWgs9CmBF7gMc4Hsn3phDQtIBGoCyJ
w7R215/nfhkcjbA2L5KegwBtHOKilqHLdoY39HMafWZBhJOSzHydkhV1uvEWeasK
6ce7qCdzh8Zyv197tfjSlcOMuz7TTn1+TuJqB9BYdGLN7yZoIbJuo8eO26wtXIkD
A4e+w9W8suiAJVIgglzxi4EXBmXPhr21sgAT99xb85BTp1ugoBnSvtAZgJ3oLguz
TKD6/wD3Be+gr7SlBgel/tbXBym2vmJv4o2hK6ja8EVi3gcV/EuiNB/1YeNQyMur
qYr8WwPgWEBl+U8b6qwut8gb0/32AxNH2FVoAZvTNW72HVAuiziMh/giNQDGvixd
ufzOp2ZHWyTUE9Dlm9vo5aH2/PIn0kJkNinWRQDb6aI9jK0+Q+wVHOSyqVCsJM9B
4BHH+SEhdn3JPjIdKrbt/ZmdVfM2QD/+Eym2s2X54kEECtuvTL2nrky6ZDw2xPnP
kCEKnmkVlfCuMa5NSN37nVgY1IWC03D1KzX4yQZJuTNKFhTb4g2g2hbgCfFa92Ub
YFUq+MOVh+9fzNny8gYpwAEkV8ozfikdYYG2UCGBZ4RoFJWqnf2BoQ1ow3JmLdNa
QU6K9RLSK0ntsWoBm+WtnU2vJ5nz7dqLkbXLLhknQhgLbM0Bj6Yg/0Zu7GA2+YDd
uVOEIvfB2/19/8PFTd1T9W+bQXdsuxBpGLabJAMUJMY2Bvf2SKlQI/+6cPPE6/Gr
3k6kMKCHaFPFqDWO0fdNBdMso35Xn6BjWHqz8u4cUeTBY68nz4OsRt0WmJKp9q3r
80jCTlVCrnyvX3okOdkH64DHxiBSRLE6fXo7/lHCt8JX9Gbftt2jzS2I1YJ1/WDW
l1J+xG8nC9iXfpXjxK4G/Umf9hgiYkw/WT8bPltGJvbxKCaVDJ7qVtzphz0JZ6W4
zTyyG35g2jrt7mDL6A/MtUHHSDteubIaXkTfMKtjEaejH5ZzWfSaVVv4kva8o9Tu
iDfLHTMWjLVRxzP6DAPyk5FziqHGUrhS3CDpXfc4J348sgkgrpa9EQFsngdRAdHU
zb6A6vNbgWJpF95dSvFWIgs+rxTQIWvN1pMRROknzhS1Bkmze5Q1+7GbNPnrO2XD
lA6/bzuM4bzmsexF6MvHD+G/M8nltmt1og2ldzqh5ldt6J7IIz23tzb2SkkkuAgZ
e+qcFPdBVen4ixJ+9rbK67B5dwlJvoOiVphlVP9dg16unz6EtnZ7qUr1n1Nri6+J
RLHNt4HMkYLshj7wiByBRvGWUEsbSqbRnRKGlx6K0p7JhlYvkiNA6NUWn39EOXnl
4xZkjcYcIj7pdqVV1pBTgrrCht0ieb/eTFnCi7IaBf3+dcWO5W/YOLWPm+Anuf+U
54XhY9sEJgnyGHKm1cAIkslOdaLFFN0seHvFl112VvSaYDLvn+55FlrMBxd3BudG
Ya+oGFj2VK5wBzsphQddEz/m/BXqWWGRNt3Ww+fJtV3q/QUhG1LwIRJvVWzp0oOy
zlufa+xC7G5d1Uj2kHELuo5xR3gPTxBmw2HcvarlZPOouzU0hKPUJnquBKpQzYL/
0KA88JcwxgIGLXqEkV6+eVlMmJRkWu43PvQWNIzXXu7d1Suyse6cEl/L9Z3FY9Np
rzgzvDRc5EKki7kUl9FDK/2cP0otoxwZ12T9G8jVVfSnXAd6oV5dWHiHE2Nou71h
ij28JebCjvtKz8WN1pGjt/SLvI0PHtNES0Zo8rGACvBaxeQSdss8gwq7TSTduqaz
d5lYp3fk59eNtMoPMBLUPLSVrKpQsGM9pUoGZ9XnhF1QXsNetopfrMpuwl+Ez+98
x+tcD1m6vwIKjEvte4NmJtcGhb1SXpaQgHQQ98xDkI5LPidjw9aJmwhGj7zi9/Zp
SQO7IUfPdP5w+pJzUkuZhKQKPxohIHleOTB8fpOSu/rKahNDDduYE6p4fTggGvXy
XNmIxYZ8R15sPJ9z9PB3CBFPUhPoD9TYR4nSeBamXJIC1Ls/j9SSSklAg5LHIJtc
WfnouJfvVkK2Cmy1egYTFHpFIhBJRGJJIVMC/LDur+B5dTK4zl+W5whIrUZGqnMc
0Lpe+pAfLuDeyd/opvat+eyz5fbCuAUQoSJAKDOOXG10geoFA7qOUeTSrNvi3ZHC
NQzeK5Xs9+NTN0sgBCnoBk6ekqMZeHiJw5PQ3wC4XLtD61PMdb53jEcuITbMzoJr
SYNSjWQ+HFkS2QiZbQ227sN7zND1pcIEpPaOmbJFUv/yrmjchILtgNcCZOK4xUOI
pjOE5lZ2ECVWzG81kcetP0vtVM2rFRx2R0Pk+tXpxAtkrECAxMEWZeVbgAZpap8x
KtoX9HChb2Q+yrY9u8Q+f0NWi3CIBLJBuaQUsBTo/sksP3hZAyags/bBaD/D9c9c
Gy0zKDXHJbGQqP5S6dun+GQB/O/jpX8Wsw1Hyr71CeWr6ZRVP8hoM7YqEuN9SN/m
XUVvyMKryTG+0R6aN91zYoHYgWTtxoOkyF/NluiwRCfwCAOVSeUt5IslzcLtCy2Z
OQCaTbyzODelcR8cokDTgCviLCjnbXjZs0jOrpJikknKaQgqJaA353STzo3YYGNh
n8kw+5uM5n7wGUUAd4L7zJwKJBCrdoe+bsl/cG22T+ZdwF9lKOaua2sYJUJ6434Z
k5tksWdSiECrs8MWiWI4R+lPuxzImQeyb/nNYx9BObq3H5awWzr/Ld2TBpIPVGMK
dy0Va1R1SuhWUvP7m0wZVKoDtBLBxp/4T9BdBMqSjy3zxmyOHbiZOD/HayYeq2Rd
/6f0wDq+3Ka5TzG1ioUVh21UoWHcst2D8FSP8ELHFHtit8kqYWDVQc5WLC041M0v
o2WOOL6yPOODo7k5umBT7hoHrJksNv5gqSsG+TTY5P+R1QqsdfA48fuqnoqEJp2x
tHKdwus8zKz1qIBqBDCla5CxBamPA/FKzkVi+bRV502jvGkhFNRtbY7u5EAbQ0nj
+8XwocOH2SR5bOaniou+YIxu9he1TpebAb9IZtF9ccnWVe0JP8NrOufJl/P3NgQW
PURtEIvH2jtbr9anN3Iyf2qAFjRA0+p+6dm7uetgVC2fhCR9dk0wcqLnOnSUHQom
0bnEacOu2FDp8tjfZ/IWcS6FkJJ9etcsOM85hbl5n4cVVFtDg+MHgbeHkWhANftK
yStFacpdCc/3On6cpg8Z1/HobU2AkV5N7D3HCvyqgVzj8MDYrevQP4ccWN0+ttOM
GOlNyCnQeSq+mjgHfpu+wVlBcaKd8E33OMSegBnhgTHEazLXKBy+1HhuE4S5RApe
9+fV4HLSiTUDuyEbbJikyGKGQbpK8Op2RjJWNVhaZtmO6oZuul1NBsq56TP6SRzQ
Q8Wr092FsWtrx9UO2ewFSV/RqtX3LSP55fIN1oWs8Jci8Z5PM1atXtHwBUR3srGW
8/aEH36DskCK/63BIEnDb38PPPqy9NyIK3ooaQODuRAH2/QWtREB3RqRX10jG0jT
/Jd7klj/O0e/emWuAVJPb3FdYLg/Vy3gCNUtBwKpUTqPh4lMHr4x7tifZxsTLaW6
wakIlCavR9/Ntrmc/K9ugmXCsWd9l1ygVXrQAQy7N0U64SJVWRGVTB8Bj4CZtDTK
sdnUMKNzVICz6C6HTKOYD0bg8049Lby00aa9ZB+sfyuVvqFrOUcbhOhDoKlBQx6f
UU2fcqGpA/UF7ihbdLPvlxjcPNs6MVIf94oe8xsTNwCmA9LOOr9Z7VgckmtW7kgj
b+stGY/21ct2MkwkB/OAr0IteYbPBUl70ZlNrog6mTR6BwLkuzZf5lq9EKujs6PN
mTP/RUBrNTIZ1hztr0unAZX1ntgvdy7kfBkeKyfUxMKIyS52FTyFCQNiW4pmEcq4
uVvObiFuUcAFTj5JIRP5i0YoKXoABJHGPNV9cVvEegU51NtQz5gWrc5glwTKsFiz
xNshpmgfeTCHjRufOsTSDWha+4Q/X/UK1gXVexuzGzv6LltvsyL6bUsI83ocuKhL
gtD0TFnt1ah5AyTsn7SygauISJPgqjsdwOiM7irgKVDpxm6krqbvs7EPZoirXy4E
Y/w4mrUXxF43khDlHFgqoewLy/FtIlm4cwI3ZJKzcvVwevpOx2Y+sXeu9mNbhnb3
ph3sxrW1Y99nxAq0lJAc3EcBAR0jFyKHmxfxyyvvMdGbbQ9R4EkfiDNQBOOlI4lt
vS8WE0WAAODww0D9UkQABK5prVaj/bUL+yVg3TGcikcJ/pJb7Ct0RlNUY5aeYa5X
Fa/hvoex1Qe6e3HFwf8T2JrXwwxL6WkMn78/Hvj8iIjdQ/0uGEvOr7Ab+WRjgmZZ
Y4lMhamU9yYr+U1PXlSqCwbqeppRoevZa5m9npqlG8YH39coz/HWehdQwnuVsWvC
oTxpnCJT9Fb9h//5xuPQp0tXqozY1iz7Wwh1uw4gqv8rncCy/UdeTaKume/RbWRq
urZWDzcd5jTcsy6SsuVWXQ6E8FRnBduqWAo1fs4AFh414VR/1Kcvz1wuY+/JlHld
1/TBrHsjh/XU/yyc82YwDuD+EVm5uw3luBWYCi34YtRi47L9mp0O5NyO3kDTuWqt
qJjpaLdFhqmKOpQuYATR56risF/BsiP7UHIqMRxaINGsyUUj5dKtlmFPhVH7AO8P
X85sxl2LTPygp+v4nD7M6z1upFffnA/OHfsPdlK4XCNoffgoTK0nsRIy48aNQpzx
pGf2JZa4/1LOnB9FRh3QqN+s2kJ+Tl98frbWXvTujprbOuc0u8V8cK99nTswanuB
f8Y7KoOLqMmgdA5b/4FcpnXy5oFqnq1+bNxiZHiBD4ki+wulG99o5nmvpi10wcjm
7zJMVs5Vkr1BCJnBMJNPXUVBM7gIWrahcYfRgBvgjPLNI1nrItnxr2XsxXvfX1AD
nHBPNRCUUhsXb81zv/OdBz6GKEch39qTilkZEDYdmteS/E5ho2ciZT/egKqbxAFf
p+85yWEPmssFYZ02+ExFvJcyZ4Etfnen6VCr+NIwX9aAAMwDJrFKU2eg6tQerfXt
2vC+U/Z/ZX+B9HFvLXdMnh9WKOG65GeLUpL3U3ugJlv4uD/gaMavVPV6nSFvA42x
Ac86uWGBy7uUiN5zI8yc7D074gdA1+P7n6X2EsX/b1OeYr3LJR1g19uKtaS15l9H
DeOknbNgHDD0vxDm5ArOFgJRXsTU4wZRABqE03gSiS4+pkXsMQm7y3u0L9y3l1D4
8QNbSL0HVkZvNeRg4c5LTLVXP6SU7ysvB6N3tOh6+4GvbVEBVehMvoNYXDlZvGZS
Y9TiVOeK+1Gawn0Tyagj+W+21INNnVTKZ234Xz3R5AvUHUQ9PxqWjNc8q49HAwv1
ewbv66Po7GfQnNTeH8gKAjFvkfDmcJAMRq6lnogh+pHTsRgQpBmCPLRLdWTVkUzb
u3GGV08Sj2n+FU9c5WZQZcTp6ElGMqIayGXeDPfQaLKlM9qU8oRSHJFfrNGYW7nj
Khomb0L9aLSBbCofLzsJ18EXUQTH88dAFwIoo7B5Syfh3XclBwzsY44g6ho2LcTi
FrHEXH5RsPNgcYUkq7xhLFu5Gvqe2TGZFLOCsbY0CoH2ty5WUgDL0HQn8t2Q+60o
aPaDKG2o41RZadYcHnd1vsz0AKUuZsGuNAldx7G+JsAjO5mVRZUyZRQb2DNs6tyq
D4sThKeQlWO2PyEgXI43AwvEnhjHTtGiW11V4yM1mytU/Z8nRTroAyuWVAnaAebw
7MvURSh7qsZpdFi2Aslf64e6gwpM3/L3AXdIWlJY0AtWKAOPyUbpx4TjhoZIiLA5
R8hqdsBFmLfZ3bZ6EXUIAHguH1DPby3xEIzqRiE0A0tq/Cuo25nmDM2MvauvQJAi
9kSNi5aspdTpLj0Ep/+k/8i7iiFasNWUMr9mQmzm3Klu7WX0EMiJe7G6a9VByCvy
8vN3MA6LN77zAzTbIIT7mUUwi2zrUZhwBwpgdECxdNsM23z1WFd40j+3Y8MDvh1M
UyLeviGPEJH/1DQpkWXgg+8Uz4bvRiFXNTSposYMGLtSXhbRQZfk1cjYUuhlty0w
Tqybz2IW2Q9A1iUu2pdUujFIOEBd6arWQbGYTwdIbKqwsMO0LxfQ53ut3HNxeOud
tZ67zz3BtRtP4l9W1NHbLEJzYu1qHlkw11mhCJqeG9uYELBqn/X+9vyrReVsfBEM
Ekd8AoIUTrzzjngRJZITXmU5JTJClY2yUq4prIf/heSiEevtxCNd1qLgp2BJ78wk
4RCOqI7fLg855Rk/4FbJntw1K4BQFcuNVvnSInkPTPMgBkCTMKVFwzdQFqep67cm
YRHFXGWanRGTE2l8VogKW89HKDXxGDe+AjrN25CpCpO/JXzrQZyIq27qpjdwnExa
NpCbF3nuL+LYI/4AZDttB7jiRVjss6hGgjYV88KEGI70mEESZGG9kBwJkcaNd0DA
G3kw6l+IRUSGkjzvG8H+y2LR+rh6lwz0aL8ymQRPUIy0i5uxDeAR2MwGn9DMFCMM
p3yJosvPS5g1ZvjsU5XNrAl8R4t1GCMdKThFI4QOGgq5/GqEqcgjgZ8X05FYIRWo
quMZT0GKDj42vZMhg12NaTQHEMflEJCvr+2CMqiDfB3yWMxazXIMZzVYkDTG0n4M
0CgQ+3KTDT78jPvy/ASa48yLd8NzA2S1Rih7uXxNP2AZj2mYaqPMsXKfmf2i6Mig
Z8ieoxUm4X6xejFMhK/bNRo8SmCO3OYy3I83vEDI7g4ppH4uFVBx/OFGr+96WE4O
54NyzkTP61L+arjBkmJ3Ag8+gANx75tMRD+xZ0T70YD6zg9dCs+ZFjRQaej/iNJy
KrRxiWDD83wgRK40dxH4s1aB5b40r+aRSAEtVJV9CfGcV4eVWUe9oZhWfXwRUlEU
7CNuc3giPZJ83rHd/cPhlyxh7WlVAntINvwYulC1p1V2wvYQaGGfwrzLVPE8rfeb
Vo6a4I6hFISkkzdQZBk6eWdjMl7FIpYjSr29T9aVBWtbE2m5cHHjYmXcjMwLBDlh
9LJSgljYh1QoS7OoHprja6nl0VEp1xSsgb4l9DnBQFiBo8mew5RkEQy//tfnIgsQ
j9wttqpM2Zkqza8gKP3cUEdkHJRvC6FRplqpDHJov9/dVcRGdmGUWiLDF4V7DskZ
Oaq/NhKmJ7YNPJquWy0vzY+8b4X+Cy/Th7r0tcTVNgt8bTZl+WFlupa8Oa01UZJ0
xYTS4LD26kIy5BvOhiN2LOmWY94LZXuqaQLWPL8w3/GT6mVipOxyImFGhC5iufvR
1hjQBfl1PWCg+wKBmmg1UH9YasXy0VO27N4NvfVmL/Uxi02JSc0UGY4lpJRYVRQ9
HDzHBeZe062JkgpwU9uWR5RxcVihaavsfAinBk2M11LJA1g2wsDRGn6JNh5G165+
7nhrhWuG032DkSl5TA0JkbyGDSG/HynrJtdBbaS7HeI0b16r2kYqYMIHkIByDSro
oMPD8NA4YMC/Sa9vjvHy7OwqYkU0y0TTeW4GtbPmlY2XWjP+twiNJA0RiQApBHw4
6yD6WNd4axWL8P76GEf9IL95Mr+hBGFuYKUym2zmh0PXJeQnJ7hV34o1dsHFkCWP
CaawL9UdTwhQ1daPOrZxyQ5LrNyNIE1YsDjRhj+dADqTA0HQa7uJ2yZ94Pu3sz4l
FWZpew/Htb9daec9XrXbPjqmuyYrlFnVddJUJE35e+2SCujmj/q3dqBosgBYLaJv
Bx2BS8aXB2kCkzp4AYtZowSr42ZjsYyPow/UTC+sCgxjS4Mp23ld/Hy3YNvwJ/il
Lhy3971tfebK30mwqflKYsIF2ZMFNZ90Cug4MtwYCJgZdQaZjx5T/tWfXqPoLID+
Mu5u/i8AX0qbqPKEAPLLU95hInnh4uNORR90uaM29/VMEYTZKxfoP+GvlwbU/hTW
VFLcBLcxjVqd3we4/eqCCAcVlzxxkdDxUXbaaRYwjl6qbcx5RHEGyfDN+AcVRGSA
9TusavLbTFRC7GPuk/98fd7/KsrEXRaYvu00MOiXJMC1UDc2PJz0nDBmHJJdMyGp
4mz2fpwKCqnkwwSUKvJ7tB48Vm5rS7SNgANUReWqdpiuQnZFsthzFM0UnA8xAKNv
w3R8XaDTWM1gFRK5QfPJh7F823FmsTaAvV2rJ+m2VTTYEGbB9s/pvJkhlH5f/Pm1
K+MN6qZ8mUMqMnBCqweVghOeUuE74LqobEf4SQJo2jk7sAJnZ0hSfHtBFN9D9Eo1
8jYrskwo2SiBvSl0PKgS+VRci1yq+LYNtCwsKOiaeKqdfJsVEidIBU3tYyD8YNHd
09s8JR0D1x+pW4bXROkSxZcfh1thlMFIaSjoYLDrjk9TPuqdrHA3Rcz8qR+/SBG/
Ou75POZWYEUo50QPHDrRsN8ZgHC7l/BNaYL/ULg2NzdW82afQ+U7TqV53+OVL97d
+HUW0tKGPE5CG4/tREHfCh+mF7ZOqdbXkpoT/DCuephWq6+va6q/h3uIzeYXViUp
i2F2RytisJ4+gTZU2AZycnBDPi93IIari5fghfFAtxrWWSeKxBrH18oi8tWyehU2
+bgCa+go5iFSreBwwn3BJZAOIZP1LzxV+0qIrAz2ANXCEtVRFNDxZF3HuJg3Y2q6
UDiHuQoNSxqL2vL4xAJHmmPGjSP6ABnVQy1EzRw07q3VVpUMA35OjM4ll6dl1xv5
0eMbpJoycJZ3y3U0oB+oQczqscjfvLsmIrrtwMC1FXsFixlt89EpjV1nVI6gccaV
8Xy8sCpic60Vh9mDnNh20uhNFtR8cZSTm2Z0e9Utp6slWmisFePdSYxG7kPRF4xx
rXuGiDdgt96P1aS9S1e8f8TViZb2uY9YSuRus+fvRSjCsw+GqBICKxD3jBqVrp8U
7/43k61YCKdMcDf4NU/aCkbNOl2fiVCRo+Ise99WSje/VUz9vHe7qAPUswiqcME8
B67jH0xPjjxnlMI2ox+v2DMoywzKrV5L2SsQaUuz6XpcoLH69PP8jlBgV8eSQ/1t
z4p9s5ZguvWJvdBFhKT0UK0uj6Y/2XKMKiqlst3uBclWnSnnpsvNnHwBYqUuXBY+
DE1K11hXaSbtzgDs/jzYghk8vr/KW9nmpk2SuCFVyqKr5tetoLJFpJu4vrvZuWN6
aA3Cj7u9HMO/PZGBdyV4B76K7QPszuLyUF5u7AkYw4jT6uaBZwFZ2uHZ0q3ErAKU
0m5WE9Ot0FOLazMFsZa2QtLEzmJ/ZHkH7+iJ2qCE7Mx07lMAdZXezNzWFZYAtStc
74phEY9Lng1AA/NUn8uCUXFlxQsBjKC3jKF+jeqNX4Sq6JbP7yCdvi7QF8IZNr5Q
LB2ho/eYtKrHP5Srs6xliP/Vmtsa8HGRtYKfL/SzBiO6fOCAHZIY1ZiiBiWrXPfw
7R3t4R78xyhwlrkNmUKN/FhqnefrE46J9YWKx7dzrCsd+aTp0ohercxaE2dLZFK9
YjKxIXuGZg0J3gAXERzg/JBO+9zbmfoVXI1lPiW9iOmIRd6Vwdc6McEc4aBRaGyh
OYKB2/vwImaA+WkoMk0AAFIlDsHdWKcHHDhO7kYCiN41nfx5RfuQSxWwuVNzRYD+
PzLb1xkVf4doIOxym+ZSZkZxIHYMfHLDGwZsQk71l0eyE5thQzqpFzGfKJyJGkQL
mm5o9ALJdBJCKxxN4hFEyVNG6uZYxkdHJ571KmXVgnJvKNRIV+CiuDM0e5Ve/wKo
qstQtJBd+9b7AhkQtJKZheKgmIPx5vKh1wquilmEOErlgZduRmunddo+iGQ9fNiN
sHs6UiDzrzClLJzB/57p8Y5MyAP4W14wWAoqTwu755O/Qyy1q/9y1ztbFn/GWvsV
7NfjlCxLt23msvLTRKCrRfunjUfJXktQD3h1PDmM2xmXkbQy8B2l7ne3eH4dG6H4
4EEFfMk1Wi/kKHI/G1MFYqlQpYcc5sYZwJ8MbQyFy4K5OsJgBVszKiljcpwwW+2Q
pYShlERn90kNIja4je9sejXpPczXLNuZF7EoXrZCnE8deOXyWviV9VxQzO8WUEKc
9nKdyTdKOIJK2e7v9RFHknCmEq8eO2xpm6tLhwm41v2CKefqWQg9R1m0mw4JZqdh
cWhAKwZq7zZHyJOC1dHq40Fyn3D8Xdffzo3Km1GhhC4zM7TmGcFTfSccjIj4us+P
IFayehjEdSKC3CHLfxZGlxoefLZRakT5CVyAsMStw69OQxX9KVcanVojiIZStp+b
4g3LyVhgXmxwWcobY4EoBArrDM88MTHoa2XI+iIRpjLp1dJzuj7Edh7E8aICJTu8
oLD0BYQoR4IePaa8vSzjRV07YFA8RTHkQRseacfdDoQIMgegXFzZn2osA1IArUMa
Y3uFLetUpndIDzxYeWqCC+FEL92wbAB0AvNkAFmuUVnlag1O9tpYHqMhqELN8WPQ
vPHnncAfPOkoYk7f85EH9qMhElwAGsT+8fCIZHJ4v5jYSXashWZ9WwwR/stBVYlc
/1QTFepC/GmlIlyNVLV6KTHzKrtCjE+E8d/+24IvamhEsbEmKbZpigkiPUA9igZo
UK4c6fx/OsEhj3vRCtGUAyUk8rBbLTVoLeliIVyLFWHrFZEtMEbEecOWi+GkJ3sP
QPn5C26Ea9weVv4DS+SZamwvZ+S9V2P5Te/7GXShK9xb7zgxC9UmwSj79+M6rLUg
xzoPZxd+0E1BXxrWg9d5itAg/LLlfOdZXqslCNzMIPFRvIu5JQDiqQsZVV/QY64/
W5519GVq/IQGHpCoEomCTNIrem8J4t1UxJnSBag2QWPDp/kwe+EO0ozAA8KLvuT0
bfRjDHJxrYXwO5/VCucaj/XEL33BoiyKqY5ua5toNvLsZ6+YSDOpar7BJBzNSnzB
Ej9PZ92zV6faMghjlPJAU2su/F2DUl6TOWf9AqG9GuweWTf+d+pdxcsMpg4xUMm4
nL7NYZldPVUkc96xmTDCD+zRDZyJff6hI/YWEmQe0rXWqUSNOssIUA5tPd6hFDXS
SO2efKtyBQtrg0RlArT5QWhLb+7vKXDwkhqCPj58gA5FS16a/rcy0Te7IPX2qMBR
E5JxM8OWKeND4KcHarp2UQDwOC9qouG4E4yE0RP7QxEGN9DRAa9kVGPXLeoZXnZp
5pW/dqfCOdnd8AyftzQdzDKhvj/PnLtVX4DcXxJIxPdH2/y3KtrQEHYqBK3a4otB
SWCVhYLiPUtIsg1j+6wKotl/1y0bNPOYvZVDjYyXEsqCo+E1EY2pp6vdw6iL+5Wi
5y1cMIF5MBwzTrJ8bUt8NXX90kHMNZ3YWkkWZQI3ct4KK4Vb3lKr/RvknLjd7+zg
IM24XB5IZ6vC7C+RqeExKzNTPtcSm4DuiWVHPg7VzqtY0/JYhXtRFyabcQEmUKOA
w4kwEKAQJdDrQqnOj1IYySSK9M8exr0yD5jQeVd/u4tU61kRUBisdG/XHeTQBqx5
Pzk7mPJG4WcAAfhGUMfiVYlY2LOCAlUX5uUFd4nOj0PGLkBQatDYWvf84iSkoqKL
gas6D2dPHa69/NtdcvrZPg4svIgbWRiTBUdHSeNtCHZr1wp6s8YJOnXkrqJxjzSh
4bXdJPK2BpLe+EWyaikMVpUmbxetM2F1zJqtkGeIydkGjuZzjNkE2z06BEUpDfhq
cHB6C3zc6KAL9sI7lulI7ldyYizZ6dnF0bj2wATVUHNOy5+bgs0wZQLp03BKgvSM
EsXn3MxVZIZ+KCRzJFi1bZkef6uX872o0XYfZU1LbXex3j/xcq+gURzn3FcapSQe
1Cf5esq5yfpTtagKTb+kNIssRFarpNUTPoUSlyduQiSLxzXq9D94mldQfzeACS/a
LeN6ELatwCfbd3C0PdW97/gTmw/PenJ9iM0fCIMs021NZkbNBNug+SNGR9t+Hbyv
kkdL7WaCWhfEysEBGk5lajhH2v+JCyaQVHeWa7x9r7m//E/6qln2pSWsoit+lBJ6
eiyISbW9BkLGebSwdqQLHmSUDcuXZ+GVUpRpNiP9WM7GdN+N/smSBQQPgyFnswwz
w73JF9RExDpSjewFMfITAGfTON0cDM6e+xD1D4jmGmMynLaAoB0sdz/Jy6WJHjIg
LGPy2ePhS5EXbl2aXMagOxT5C0yJ9JDv1565L8CLSEhbNl0lthnXBxt13HiurUwW
EHisXxpR404P7Dz1U9WGqzW3IBkJxiSTtk1RCaGmCcqYgioB9a9j6HLCQWf97ki7
Wj5SNJ8HCf2cZtgdfGdPdADIIub/Vz3operf2vqSj6ndi/QbaeHdHFOGBK2osZv0
T46tbTtuIA3ouuEM4bae4RAO1bdeC9upz7L7uzzJ1WZ5Rw9pk0KMPLTWDj5EYtpH
RJZuKHjpukkOBAqlAfIiN7Z20MhIs/4M4/2SytbDIm7h51q450AuzwE83s88Z3Bb
11dg0LbUQtEznsPoV//5zdnmkz+IyOFUJF0rMOvWqgX3WEUzSuieUlTw/NvBd3I3
JC97rbvs/zC2ujGQ6D46HKPh2Xbo1gO63WM20dkamIpzjqxzbhUiPKcyI+JvH65R
2kYRxpzCV9I+1D7PLzrgh2XJnt08sfrJPWPZaImtAHstYFHbHYUcSV2MZrrlzzfO
9aSUm052X1fo7DshhF53a+J4DkoVPCMFhae59F9QMMxhdagAN7GHvmYr54tAtWQl
u+Hqjl+Ee4+JfbpZlAAzRdUjWLyA1BGi+jTMxgel1hZo3KCWPNNsY/4de74WXI0c
DAJvEkKBhJzwdezClGC94k8U+jaslL0cC6G5QB6Zn5MntWEEzCn0aZl9V6rM1G5X
8deKmMCG+cwYBHcPhl8XhThbWMRg3by/iY8JhXAlXmUxGtOU5FEUc+k6nnUJc6G/
+fkCMzV0vLydPJcVCsDCy2gYFZyo47KwK/qCx0UBH1tPDWonhJy3CPo460EhdL7F
otG58eJ65o3QlFW/kl13mp6x4Pf+oWJfyWD1pOIWdrdCCD/6JLFLs/HFhPknvK6O
6OouFRswnUz/q7dspH4SFBIjeiYo2pKb3U6iPaIRwqfUOYqDcyaA2EgTTKEGRn9b
whEfxlqWvbnMKsqOPM6i9i/tphjSq4FaLqJ6gr1cCkk0G+OJuF27O03OzdVoaJaG
uHJqCaWZkBz0gPmmFkq6hSR5H84ZOvFi8eOhNbRtpkPV/wZrIxEsRBbDgaKdTab5
VggBGV1lBsmt9nhiM87PajXOTX9eIHBJlLMOiUWNdwVcmU3LUDk+3kZiNfk02as/
FUG2ZSXp+lueEC6ZlvPj77029G4CtoNFWg1vzVOJthSpv2eVTUPvRXCaz43rb7lZ
JuQXs8D93e70RHsF7u9D/e58vbtPyLtNMUAOBkuy0y7usbV1CVzY53DPrxEjj1KE
RDlNvwt604A2WpPEhEiMGAsvXwuxHUTBWpVzb6t65tHpqdzEEbXfxIQkk3yJAypD
OUGN0/uxe5J+oZ5H4Sy4RHwCNf0T9l5UFa5PYwRVRc4CwWI3vY/xrojc+adwu4qB
C9GBIW2Z7io0aQDuwpGXldpqeqyvy5nW0cys8TjLKAQj9ev/SAic0tMHfCJO+oBA
in28iWzvJ8Y/ndCkAA1a5e723Xet5E/nU/xgIk/1qPADIdCwCEfUTuwENWCelkGn
KMQrVjWg3EncAoczTj5glVXcgetnuXPvnwovExje8oAPMVgk+Y4E4DUpFJApSzDo
KMi4xBRO1qNKYIKMUNfUIOP207tUFxY8w8cE7ZgMhx+LM30s7ONaM4DsEaW8M4+O
cAUy2kVrAMJK9Nx3IargOS/0sq244OViAzVEA6/bRv8mEGnujrf+C11XGm0hbVak
3Z3oakTk4kKCaJHfaoP8C0b8a7JXTUFbED/KnAp3ECmBYOvP4bwLhltI0vS4ORqJ
4KtivbFFb3Gq+FfcvH577Kt3fSRzJrXEaicjVvsd+2T7pxzd75aoRQUy9DNc6T3P
aPY6sqTcsPcVE9QeYKtDEKMXB4MHp/HruyhCKKJXVKGgh2kyBx2SWaY38KshAHfZ
lmE2kR+9cpBJIATFuHUaiW18F33asmhO/eDzln8jVvu3CEcqouMtNNDaMFLCY0MA
2TxXIo0Z9pTPpf10CZ4PkG7OnHHKG5RaELbPBcBD7dMaedYXZHZ08ijY5uxjRZjN
eRJv7j52/Oti2MHlo0mfuOVzvpolZQE1e6l69Z1i8QxqACgDlA8no6yuuMpiXcj+
+8KNmOx6hYenntFnjJmzSa5xxB3d3WIEQcf39aH0rI47m/qXnZXvR++6bdh0S1KC
8HX/DpRboP4glXHxGobpOACksm15KDVhTKs2d9FJHGmB1BduwBXmm8xBoImog1cI
TFjnkRY6Bsb/AyM3e8+t5qD73+dqRpOvU5dUzFDa2EM4QV2BDqK7VTuAni487rrC
JqG28zjTF8ywqjvl1poMe4Thmm7sIRwxd77cIBPO70JZxzqkcMqaIee7oc2qU3+k
FJ59mBQol4UdKEhUgfdfhzcwLWSQuzELyQAOG6WcYwW9ctvI66wL3v1hj1CINd8O
tiRWmRgIsOXcxiOF0eMBrZs4MdyepTuhWhyJAC0Pg1N00JqR4gEkGFCq20hfJYDv
Zt7IH/3K6qR8gfLFp2PNlFbWEIi73reE19Hdm8v06PQvHCza26p+5kobP1GUQzYp
zkMZC0FvhIdqw8nnkRyzMEh1RsPl1/Yz9op7Uq9/QNtzhoS0PEBFcDMTWiOpFUka
I1A5MgQ3aHcVkdIP8c6IvKCJGEXqGFSPaWKT8kIsFdnT7qPT6jwzbSHCDz5gT4r9
qFahSpaiMrzjHgawhQWMvqWoWu8N7YUccGr+uJPhiCoA9aK0K65hv34QpSbGnTvz
hfKcDGBbRvCy6yGiG/WDVwseQgLUb5yos0TymX5lHSut87Nh+gozTCkLzD9MH/m8
pq237JhB8P+VuOeWKT4v+BgB0Lj72lVOBWdXgr3n+/z+40s4JIOq2ic6N9Jhc0N7
bYEU2xSo+2+z4dRK8gMRfnRrLXJhf7zwBifN7j9axVW/vW5CA4A24/OKo7fk/BZP
Uip570/dZSJj9O4SUpAI3lf77UY9L12u28LGlklGIbzEvakMLe347nsXZa5DP78k
e8GT6E4Nm1uV2oW9TJTKB+nlbPpMeSeVNod3JVxq+yOfDFUtHEY4iiy0BZQwpcf2
gaqIQmyjMlbPYLnqDsFVPOg0o7UR5LhIwMsqZ+3fOPAv1i9Ak8AmNjpaAm1h5P9G
bn1rG3IeqDS4IvWf/ALZ/MZI+/LzPw5OjYSKyGXnVSsF6l4Jptspxgc7L1I5UDTO
Cu0NkxD2XDMcN7eE2yddsiLZJ99N8n2UWFACVNex/9soVlfvq2hDCA77SEYAoaM0
q0eGPJyZeuayApGYtgyXPYOS05kNNPjBfCteh0bm2bT/FexTdXFnlaTxNmLNnbA9
qcc+J1v8xgl+RLEXPgtSGvF8/6AIg08RzrBFRf21/37PIoopp2VZ73d4tsl0NdNV
MsGH9RSdT+iMJsWZ5PsXP/4euLT6IR6x5SZtjXXOAh32Dv1+hRQIQADDnlu9cYaC
zVBU9En0e+7RvtuSrXG9jCEy7y+QlSqOetVH1iSys1LqL8i4+wceDBxvmnWVSEGr
Ybt3xD3z/tCi9crUL5coCWvy8D2iiCHgZxwEt9CIW7wolZeobpCBXc50j5YHiA/O
CqV+neOYgVzTVrcaZkvh+rGL+E0SgTMUOrGsvNr+2iHZGP8Sqdj0aX++CoezwxWa
TQPzRCaZBpu9OsEMxhcy6s+3KXgX9HJEa/zHt2UG8ATOh7SV1PgxeO3tDa3Xrmgz
GQE0pWlxnzBZ9ZyhpQ08bHYN9JjFvfgW1y8pUy5+qGF3D7pluCsyMdHvdFGrDKpu
Ku5fs0GEkKKPjxKFPtdrp2DgbX5tPSN1WCt2Ma7sfgOTIIFKTA/W6/YpQojbb84p
t85xkXgN3a95VosOEo03T4Qf6c2xMtUXTk6A9BVN6p4PWlLO8/QzRZVeEb8IApDt
G/L3VYpYZbE+/H0YGcpvdRfH8WfK6J+4EI1LR52HbJq4wVyxHxzr7p/IKahDLckN
ie3jT1EO4aANosGAUc30vbVevSUDlsIzEtBoDs0cHVJ62CdTCaYe7m3c5KGzI/lH
djDUH5jCA1KwKwKcZY5zYf2yMuq3mG6JjNUcrNeLywUHbr9EwA+pnLH67Fo5X4yw
pEGkjStHzHw1xaR4DjPAs4GRnyVtnMLRlgonCPcu2IfZLoUkSHbtoFL1o4kkmqJ1
6ZdVAIzgM/1o+c9zBG6OViYRdpnJIgBZHd9p+5krFK1N9doM6oUqn4MKRW0n/vXT
b1as8KZWM/UUm7T80P914llH3umS78ujF7fHUtucbu2nctNQ0+bG2WX0bzXMUQjb
RmIXujV+esHEKMUnJh3B9EruA0JQaI4qcPDVnMkvqdoW2Jpqd+ubLYevL+OBbNyV
RMjIg1bT3axumkoOXqQcbfy50rCBYTglXRkBuWKJhmVaHeNmPl6Un8/VLx7pCFdk
RsaEtYYUkxPMzDgZT4rcwNNAkX+O+S60AI04/hH7nV/Pyu0r0xNy6Tt3940lLtx/
1QqfXLKYKVNca+aQg8nOb3eRJS++9c3CbXBzVavB6svRVpWYTFz1xjduLRLyEBda
qeRR0wyI924bvm9QCLJb7uI+ViyZvPyTM3PUM4Q0xnB74cMba0xQFzvJIR6wgxjK
40ZmzYdK/rYs9tg93LkI0KbUsZ+Qo1kJpOt4c5DvzoXXAffmemqOW9lHnIRtYZP8
JAmCiS/cBpOujmKWS8nj+YKhqQCBbvPurbjCdQQFydAAYzPyndRJ9XoIXrrh208e
beMX9goXhGfbe03rfSZoAowB81MHNKE0O31sJPjdEqsjtv/WMBfIVnIb0Cdkd4NJ
SdT5MXHvgXagCTEy0GNh7hPnbbz4mY7in5lp1d8pV4ykRe+trzAytNKs9AirIYUm
Hk/6tDxFOqm3VcNGdRvgPrUxWYlyfsG8td5fjkZG3ao1jyQb0ID+cEkbSiKBksgE
naqjSpv0r0TB59ySG1yvRtW/35QuKDiKB3TuCiKY79rZaVHjgFUO/CyitpUge8/y
GfJkCv9L9xG38WIXaqFCdrRWF0KjmCB6jUr1aYULldDMH1z0ukY9ruQJ/yzmfALu
eiJ/uJQwo16TzspV1uh617x8bAp0kqsO8LGIK1vkXvgF7tf/7HzqssD4l2KYEb82
GyBN0iPBKORA9YxMcK42csrMvFt+3KzfUyP5YLCHnYb2HRNnPoFj9ZN4v218XByO
rhwLFbSs+H345CrrMdSPlHjG5KoMOawPZVlNY5b4wkM2WAEp0nHIuiRQgj7e78Z7
2lwKA+0HXqD4BLVQq499ggp1nIdUZjzK1JlOKVhOfYX2qJ+zFE4vIW9IyTW7xN0i
cDOx1u8JmDlFvLgrWaT0ogXaghU0gphDvxCH03bKpyVWT2q/+sghUgLga8Ie+HUT
uVzspF7kMlizb48LkMrA353jCL5JtdVwBR903eJr4v+D1XhfLysal5tU/ZyDx0uY
Bjtvrz2soYaCey4EQHez7qu8SekUZihyJv6yWWF9fj2+Enllu3UbEepRzLNLNQkS
xBV7lAjWEU+ewZgThhT2MTD194OOf2Kq27109EYZL3mM/9IUCZjYAy6llkwaNgWI
DeKbcbQVF57xTfXoaaSC89yyPQzKzURBjsltXJsONKgUpphsd0mukiYInaswsZo8
Ay6NIPseuEFBoDxJKePo8xul+XY06xBWx2/DxrVd67U+2jYaxH2n44hspHcpSPM6
Uy08CyppniUxTQj8bz/ME/g6RpVGNlP7VBnFj7AUtgckSWArRopgLmwS8dJFEkiK
wKik+CmMJRtC+yMub1iIj0lvdU7z8//am26ao5yXOHKe568FEdnx7KstKNm7ubQR
KqbdJOAY5LCG5T9+IODRqYNhXlYza8ZAzlvp6FONPU5sn+4BRkAqTclq00poi+QO
UeTU5L2Ji7hgo7eGOyEbFqcHPzjz8m8SOovYfejjZ62om60XkzkK+0xz1TEB5N5B
3hkHYiXvDhodAuEKAJfOv50k9xEj1tXJEMQxPQkiv3ZT0liQd8O5hUy24Obbd4RT
jXDglNwGYKQWYDWREJKxvu60eOWmDumNjDBj2sTLJtq2jycM3Ghncd14bkBTeYTT
pH4VGa3wR+vSddJpH5ezhJfA9GzziPhyWf0q4f3lW01KB1e6Z04uKTo2Gr2j1c/N
aSEIB31JRNxq3c618+KcgVN6nj8H39pQQ62rlczFROla02yV6ksL3M5puak/GzT4
MjpzpdwwXz6nSOlOs4vdnztq7lhQXAur3xA/LsRKVNhxaqMbACwDdcuQHJJ7plAi
wSEMZAhuRHJktTXHb/fohK8Orwra5Lqa3b8yIdMlLiPmU+f+JA1EqnMcORXAoHtt
pUmhPTQrS6lLaia3j2S2flkQfanyGGf0tCaKKf/hLa4te/kEi4TwZTOpWs4jVA33
otQPGbgveA+DzQagiNG0B22/f/wbA32n5Dt3itC65R1Z7aJdn2EVgxSUDMihcDMK
hbHPzvvAQ+QENNWW1lw1SOYZF0zjKZRIkOWCbrKJA9gtzF/UW9nIRgoPve7oCNE8
rsuwth7B0oC2rlWxz/2VewhTrB/n33kAErrcVzzawAgs9sRC8lraX4l8jzA577lJ
Pef7D89tWxkeb20qjLDm59t6hQC8Ei36N/s7NBIPm191bPgGfn9zH8gfsOE8BK5p
ApQbLe+lLTp8n5ZbMKdVecnU9HpgdzaqrHu7wGXzB3tKPmOOig01HJHLcKgqX6M3
zhRO8L73slgwyqSVLsBPeoJ+AoE0cqCNi6muBILFDBnkRdx2sLGNBQqwqMWgc+C4
6Msh6VtqV8CWIjTcjyqI+C3uv8noTpcZyoO4KUsOYz7UuPb0JAz9BT/2exBlytE3
JLkMKgfkt0CrYwDfcs+U+39FX441dlc5hHlcFDKnReOQ3TIWulF4LwS6tMRhYboS
lVH3+H8Javysw2+ybmnPqaief7LTngTM97D5uY/W0G3BpsOVoZfqKwPNi96G01jX
e7roKzekYMAAvXProCXhqPogR5iogP0caVf+v8qmRQeH7vD37uuxymVx9NaSAk1L
tYPDkCxohu2pMPb7TeCRY9/pguGclHDTsKQ50BxDPr16Qk1jWYdYVV5c6714WOXs
k+OYOKElzh3Hv4+JuNYDpd/WnrFhmzzG4AAmn05zVe7CQoVWvZcJz+37+gG9/c68
FJUWdQjmXsx0Bx/pjsyuajpAtWSVRW/wLJjYOjWKCgcUaLrXt/dSVtKJqakuxxDo
Y0MdFwDXBmmCLaWNc3ABjmOFAZhZd07LZBijOxi9f9z/sqjlAMyE+a79PGcXIfpn
+HwZyEQ6Yol198ln89uRNkKbSscgqFHJzj/eRRXNOkDB3wsfkYzxNrHsFwJzWzut
c1K4Z4nybS+36QA6zJRQgbiTalEwm1+9kTWHpFu/LJGsyUNLIn5yKU+rbpI1EQ4U
UytLCQDI+hLA6VPKmbp8nWdeIzcyDdh3Mh4KdM+V70VrbfQ4MIynZXMIUL7rjTR7
y5fJG2We9E9QdodGyGMVm/TiFMZSctEf5KSYlvNacALBM3kSvqP9NySDZFRl52f/
hEqCvLo7N2rOoH3b9Rdf4FUnxuZRYW1dART40qiP/06CdNUv4V8TmSHL6xV1UQKb
caGgtkPbW4oOIuI6fi3/AVJqiYfFBF4rB9c6ELeKuU9SMj4iy6RT3EUJFc9AZdqb
gAxlk29AeP43Jl5W2r+/zz6rz0dlGb67MuBoLAuPh62MR1Uebl/BKtB3Z1gbBwuy
1Mky4z1Hg5NABsyvi4P/awcHWcUsRHN+K1nQn2bzcmFxKSHa97RnVo+hxsiXuS9g
rClzh0XrQRTfDCtiJDYdpL5C+TX/RkgaRrQ0rJ3aeR51/hlwvoXJhtEWhFuIzj37
R8CQeUd7IBeeN7OqErj0prGAUGEdzNmzgopeFZHfCHPNEgP+lHpd/2GYP65etWhe
j66DhVP9nULHKLNMVyFaPSjH1bEubXCqEKXtNep07HLo3IkxKYYzXojLirbaCbI3
uZAWpEvjiGyflQh3AP233OvzSD2rvIX5GK2JiIyTuEaXATQ6UP+ir4rSvMqi3mZY
dh2jdeJIkMA+/dlC4r5O63qNilACMr2UU9WV/I/VE/Vd1fgpT+B7JebtNNJ0v6Ij
f7iqMBuWVMkVL2OxSz/I3JgrVEp5R+AEzDOWPkmKFgsn6IXFQ0Q39rZJFMRsn0rY
9jyZSWQ4D+pf2Gk8zPTjtIicB0WqofGFcaujpjMaK1Z09LVk2qCDAS4tcdSJz4pu
NMasVraDKCIgT6staPttGUyHE23Cy8ytpkdL370+fglUf0K1rvy49aJhtsKrFxFW
ZuyeIadbCB/sNjEIp0QcrvF+T8ju88Lui6zjKqvGSoknvKtdFxloSQivHqC+ZDgs
9ULHMdwpX4hViX9iE173daM2JVQKBgIQBvg3sEtnT/fa4D7l8ZFtGBykaGfxKWa/
hz9wWcTpOEftlnTwqLsByOBaiAlLsLpng4D8k2GFtnEwrc5DXGs3gUO8cp/4REYF
LO0m3WthysDPfAlieix8lsesZwKiR/SGk2fmryloGeD2uktDVKlL9hcB22lUTneE
CA2W3VRYVMnhfxTBdMKI1v1zstswb8g0Y75CSoYB4d3yNUw7W5sKM/IoOsjVY1cC
5lle6kfB1+T+cTTkN7szAusFRQ6q+w4E4RTO4HEau0sLoGwfpPZFuX6q8GVdtEJ0
M9RVda2GX8Fp3xeZRZK00ytiRFmuPsvCxG12UM6SpftgMl+5CRxIiRAuLUqLoe93
+k2mJn2Jk+pZ/aOZVY8in0X/ie307U7+0fzZgVPYA+dOnS6x2nCJxhRw+V/Dvweq
kxF6aRsa+htx5nOdPDQhbgQacWrdDe7ZKhGMMzIpAOEKPG5kFl28RBf9W6i8N8DT
foaM67af3mxR74axC8v4JhtVISCKTWVlyoJJSnL98As0hgl9eszpwruMfWvflKHI
X0P+zo3IZiD11eG7/P/7ajz5nJgctgwT+VuoegDqKKe+G0WbxzcNKW2cdupOdr4x
v4+C6U54S9c5Z7SPbF7c7jyt+NkwgnIbrK2QF3NER02pnnRJJObZ1C2lPhQeSc+i
fwRz+uKL+d9SZ+Z67Dz+Hw7cBF+DGHxzoSCzvLVpcpGBEGzumGAeb291/qYibYTb
XOSya0uP/1P+ngZeD0I+/Xzpcr6GnrjuGIDMpUYw8egrPQJFfWxy/M58Pw+Tt+bJ
WQMuEJmy1BQiYCH73pAj7ok+TdsoAWYNJmyIgIdlgqVeVVwEzZIXx5daWbL2uY3V
w2B1HR7wWOa73QN024SIEQjAXCS+PTNwvmuH5K8/YLGtLkFx/QNtRnj/6+G2w0N/
SwJLaKaPZDBYTIWPZSqtJ0qEX9JFwCmwX/xChSDRboQ/9XqIYYt8jv6Ks2nHR418
EA821Lzz1MYqBc+Guf+STNVo6I43y6Q+5oc4jgkSocFpz+ZFBw94JuwfwBR32b4i
Mvs1ygNBXbeYbgIG+C03F1rjVINBUBOoYF1/2egRZ6HvWDBt3IfVYkE6s2drUsJ5
BXD3Omr8y0fsUR8khtYwIYfiKqPb1ZS489lhYYyBcY3vGXuXnR9IqU3MEvX0S7rv
4PLvx/zI0ZbS8UBJCxFWeg7wInfP8hy3DSSgyVKFCzA2M/WvIemRWFJznGTEixxD
mnEov/FWB7W/kw/ZIHCYAmwB02FunalKyMk9KrQPHCfOIzxtFaJmhHU+c5wqlowp
QZ/szsPNn13UJIDFCiWltJgn6fcHEmi/iXXr3u/e8V+wlifMC3qzJiHyDKH5tHas
nKfJPmIdvhfHdzCU/tqR/3doalSEdhsa/UDhQ2c/1j4dQAQbHtFxJzt2gm3SzFuz
yBfTiMMlVN0rdrn4ujPv4mN7iyRjPVtNnNMMJGJOuMp6zx9XqzlUzOSuloERw423
tjL0+Fubje/EiJvKlc35cCZPRWKMhw4JWocdRXIEi6rZJNTeFMPjOGoWL0JXuxCl
Oc3A5KhiGawd4XcGwJPInMmb7CcxFE4ANVj4XwzAS9XfAMahr2XHnVDWeKFMHbpX
PBmDt/hD+9AYRM/QszQ94gs5RWjKetMmFXWQ7vIcgVsd2b/7gu1BRltNarL1vpl2
bNJ6Z197dWfNl14n42WvQdUSw/tAvso2oK9AEUOiC1C+UWs/At2WpwlxOjXtZxch
kcX4oAaV6MK8T+aPU2bmbxuGNFHJbB1brKYtykj+Ce6jDzbFqOkPH8+zhR+oll5u
ANPAk+kB6gwR6Fmc8jnOUfcFxUBiMWELxQpPnjNMJqyOdGdMJyNd1Ku1jaMdzZGe
1tIQ+sffZIDUIl9ToHIQ4Ee/0LyrxoULmdJHNrYXox8FqcGtaYDcFqTAPtOQ+s6m
XyoRPKjcLbLlYw3bY7lp/CsE5dLpy5R2/MUbWcLCVlP/w1++4mX73GKQN3a5qz5t
gKVDkuJfPTvqNl75DGuOGcinDqgY4axhx7KHGm7YISBowy4uutqgVxHuIYjFl0bp
+5hJdkA9UybTOaFW/e/dY6L2cOklc1rW1z0qhStqKxbR8vef1IRTqXuufWC4nxWw
MbMGOX+F4bT5XMQMtHlI1Gx0HM6aZK6eaU58sMjQEDJp1HZyIOQW53mihdhI/yxU
f1nsagcf9R3FB4IR8kPkIQFKDIC7pd9hVh3AQPWfl5FtJZV7SWBX72fQOB8b3JXe
9ebb1qbPtl2JvyHlca/9vC15uEPKYfPCek7nj2xya0wuXb5rZHoDFivF6HnNpLjK
lrWKn13+A2qasZGaLSdil3gM9oPtUp9JdNlJyEVhvd+0yj/o4xNz061X9Xeuv5lw
Ykm1etDCWC3o5zuJIxtMRZqsdnUBg0M1wsQY8gfeUI0UFVRMLfai8aFn1akCB3LE
m4kZT0xEih/d861J8MnZzPSRWvtfdpjf/JB3Mhdey/Z/1AEV6yE8JGIWF7bQc0w7
idan1OV59EWwxEPTtcSES/KIvjcM5L7hZD0Jhn8JBd+V5+dshp0wqn1c2BlMXLiL
Cv3f2VWrv3h2PH3oVnoX5GJYhiny6rbq3zbkmfPlfO+Att/cN0OQgX5QRhhJT2ep
5WkVChI1CMvq4aUl8CBSPAyCCQDXHPJsxFRx0/9uOZfWggPA2NQiqt4WZiw6ZbyZ
laqtdWlSwmjksH5XEpyTAi09x3SxwJbZz3qLrBUGbJ1YHCFU6tOxymfeN2/3Lnwb
Sz1bmHRiNTXvhz6danqJH+wIdV1/8h0hBay3DYc6dVCtSoP/T7dWDCJxSmHVKY99
9i43G6nolYOpKFalnTn4lXKdXQHLjndqMY334La5sk6bLnfPyTIV9YRKEBSgrdVW
tGBxZD59QNNFmYCNlXDmIzn/vcFuWszx5t/tKreKjy2C/vdtAluUK/+EDX7MuCoB
xYHfyThtB7DYNjASQXV48MdmgTKF6A9H/k8uxbqK3sv8AGVLYy/XR86/jDLv7Faj
ajrYgraAypdtb3GWJ2boh9MOnsB5Y4+OGSXg7JPZv6+7/qQJtzUOwKxzq1xSeRqa
g/KsmPqzjH/L6a07sPUNJrJlZ9HZEWgHM7pnL1fZmK76ivqMiHywNvaXL57Y7AjS
yPHC+jdK4CdRr+aMnENqFwcvJHy1XfAXv0llyV+yy3GekggWdqyYI2vYe3caBAKm
GWjAlBp6VBbdH6DxIHwFc9zC1+rvrb6cIL9dlUQ/V/11RPaDsINPm34PliuOd2GI
csIPhejrrMsSVPqqjtvqACdeYJQJmgxZt/IA3P8oFH2GBr60FOw07Jol58igcTLr
OuYC+1y3mRw9tOir2dVhytD7A97eM5K/BkO8N7lZZImBGwEWBgSvstCv6JH+R8Hg
GFUGhLOkeDPFoNb49byNYQgmypvx0e1Vmq0gB7mku0o0H49u8dtfxMKpU5rPye9T
WarhbtJzxcvvAJdxAHzqAkFvvsob4c6cj8/rwiGYpr4vOwfAwVEF4qQSg94m/v9e
7j3RA9xrGmzOwjGilWyId8/0rTDtXPP1Tko7DdXHaq4il6a07Mt9Mjmp63pTciXh
cHwk6ZZ41PIcqtJDLclVHAjAx79RXlbkAVhzGoAJ7y+NgzHSYTHkp9EuD6j8hVjo
f2OKp46S1b+rfygs87uPhcJsbbSkiHh32e+YPUErOXP/N03lM/dvpD5AnIqO5rrR
+Enex2TaRHqQd7vRkIi+uMMZPbybSk+MGmrAwmRpqa2BrszRuuQCc7mrwcMOBRbV
d7riMm4GE4Dw9QMCbZwv8M6vyImewCejUdTEUaHXvFyKOCi3XpWEcio4pxz/fgi7
InryNrqOoiNrqnrzDbdd9cRfwmhX4/dM6aWQEXSQleVX7wCiRqil3dDq+nTUNXUO
tGD7o+98zu4t2AJh1ZV6anQ6ykhhTUvXZJ0NFO96DarOziEbvNuLkby40acyoLog
C5NNv6nn7Rch1AHJXQVOPJDgZV4/YG3NiJ1DXi971a9NXJOiTeF6lhmOWAr15EnD
RiAqQ1/Ld4DwKzxam+vQdEz/xHKaT71GKz/UYaBHLB/Y/fKxbw5fP7DYKVMQzyS5
cAfVTYBVDayAIb45Cxw0jtIpC68rk6eq2nn3Nu9/LvuTWmjAdeu7Nu6pg8vYbh/9
VwaLwgdWFJ1g3KGdjkIUlkmYnjab3LlNVtwys4wA05j+bm53xVh9Xrj0z1J+V+C9
Z1djk51JcaNAn4VGBWvdGrbyU+AR4zHThAxJ++jX71rh8Sxt94/2ZYyxjoP0PciT
8ptPZuczQPru1ukw+y/GAkrcYPg8i3n0asryJzno4duDUi2FAzYmL+ltWnO2piP3
gdNr54KVd3ODEmihVurb0gvozT4ED9VqF6jTtMjjxeVwd/DqSdONxikmwslFrM+l
oovu5TXAru6QfjzLJ596CZrn5IIay7zmCJAEWO8qO1ktlqv7l6QAoxIowjI88qOf
/w3zrlHJtBmwpBv4fxgdCR15vNBRljoPaES9F8Kba3+bJ5xafNsAZ3yxkQh2fWfR
eufLzP8VRezRo9plDjdq4nRNmiMSupBCd+y5yMEIoUMaSKcD8V/kfg1pmwtNRqoG
4RvCTHPOPfNUw/fjuaBmbsYMd5DNWkWQgr/j8osdpKFzaYxRYaQWNvpSOQimWsQM
v8C1R76A/SSg67+eoi9DQ3VG8UJ22HYCaEHfYeF6hDLwKcZBwGJXXP+tCHOdgKkR
WEOs+pauILLZKlyQ9xVA8kBYxwhAQvo9SxitQgmRqogfwXhd4sL/rhA8zjhcM3cC
N2l9M8FUFu2SS0VrptIJGCtqqJRfh3gxsliX9BXPKEmUKsqldFL947QTYxIbe/Jf
ZgVzeclFULeoyuHyNK3Bcvu6idNYTTvDiPCwhXhAympF1AnrzFPXLEwUqKrOgwkR
Vyp6u8G0KlCJxwXV3NKK/8CzBpFcRpNkrkAgIY+C96eIBMDVwSYtLW33PdXLygbn
znV3Sjfc12mWXCpYh/C7/86cPxisNeBbMoJJkBtDFjsLvlNcukQTL9w6haI9rkyF
v7Z9yRORn4u0OmPOQDJ3sFGIhVFkz+LdtJVxefeSh8wsXgU3jTOhihmIRTLl5+cU
mN3EpVdH6uT+m6qSWv+ULGQlcTL3PN1CEno9G3kkBgHYfyLDnFfJWCuhjEkDcG5s
c/VRm4XmakBWJ6UYPC2ptwf71rJjimKYMpcZn3yFojfquQbvkIrvszmbewjj/uuk
EoDJzlpfd8pO+E3tQ98DVlFnHqupSJBYpRKi7WbfuQkSPTTWKrMIQlfdTAmceFly
mwaNG5wcVc4xdE76tGcjJul/3Wk7A+8awYEeDRdYw3MRZ4BYD+sOozR/dMFCAPm2
DSvk0IrIeQDtdve42UZbHWyWsbM7CemxrACwMu6qC+JqkAV3ENFGr5b/PtzrHDXE
Gz+VnRG0iqIVk88WJ9OVbvMeAprRFrLBp6i3824ixVWAOrxn99r4kS7ukSTV6j6o
UYKZpfOACzG/xb9j4iFAuNOJj6K3McG7klYoP/XgNPitJ0aB8DGrbtZVRCAVBy+4
4Mdn+7TJF0iBXtf4A/RlI2r341+kWZy92kjS1zuoN967sghnvvXff4P+GAMI9Iyl
AFfufZmorxN9YN56qMk0EcQVk2pp+Q6S+Tk/K9ifiuyTac+drU+6EvH3I66S1N8C
AK649OXCgIYlRQp9rylbfbTBE2o/uAzb/ReuOvVOjOZL8ZGMd+RyremiRXy3yim2
QXSRqT203t1Qq7Lh4pnpUOWqvMALMX3+lClehEB4gDVGD4LrHRXryK2StL55p9aL
VyNjXe1rJoKYVks7eYJHGAm+BHdtOHvhWH2aaBrdSmC/pOMHJmsbOJZHpiBiEyHZ
NLZKDo+yVQRisBMJCXllOKTfa4ovdOw2qNzrAWt5Y10cfXx3RWH8mDnyA5Euj1UE
nuMPbDhwzjeGxrup5+Bq22dy9FFARHvXrAIfnqZKGXpEY5WsQAPZjiQCchFEcxRg
vevjli1m+fkUuZgpv3OirWkS1o04Ign2z+N+64JmkkYmduicOLrY41hA8/HgvqUR
ljaYNR8WPHC16Y4yfieoHvVEydeNC5MDywnuF7dak6IGQ47HN9lmXF5dbK2H6PCD
d7qwx4G4Yj8APhbBYQCOD8GHCX3pGcr/54gUszx1adIUmeJt55P0iboK5cqMYIme
whcE1rDaNrMEuI101SuSVqAEDFJ57PuLyl6FvxFdr/C+GlIX/nRI/0umpphss/vB
VMlMmxkp9p3J29gWqP8/JI6UqtTO1wEh5osAjguu9WlMl+1Qq4WVCI+FgIe1iwKF
wxcvHSfPeXvAxIuTnQTjcxNfCGsBHaybCEfyy27pRyg7ZuT9udj56Tv80XXWIF0g
CM6XDi/XfBEAj8eQ2ArZurdk/0mx6QzvlLMj8h/hgS3W1qQsaxugqkEdWY4Tet03
ehIGoX5Dm49zpUEiqoWtX2PsLRiu/tu6r6FliCve1Iz+P0oWqvQWo06Xa1gbKMgO
GjHgvXr+BAkxC0sjNmjxqrqGbCUbsITcgb+0Cvk6fpgtc4UFY6YxjkxQb2+dFjc+
ne6QQ+AuXvKUHjZzBLxqQSC7FvLWyk1mJOLVItlayYXyIxZlTdgxTkAxF1PS+Z+2
9KnbzgdAuQjI5A6FL5XF9fZzsTfn5n16t6L2ZsRKPiJI/bKsAVaHnuxQ4rmPtdgp
o30Daz5jhcQtwaI50wadOkNri/nSIKHJEB3kO42TvEH9SGAIWvSbYhZu4lBaSMTG
REwbxNHj8GBXHOBXteWxQjCQ8dA23P4i5E/QxLRt3GPATTD1Jss+ZNHjhu9JUuMC
fhiSoarsB7r70VcnpZso2Xc8RXsUNjy00XPHlLiVdW507DNNFbMXP46nd4YyApiC
hiOEApcoMf4Zq3OqYhtb1glQPq++jeHic4YUbiATQjE1fFJTGychFNVHvLqIT7UY
hBml56rAbjGid3zQ8ov7KUoz2dWxfaH31+Ag/qfL9L3P01158KScrvceEAJP+2gd
JTMSyxuBjgJLV+LseF4So1DdRYK3abHqWu0AJ1j1YJLPyQ3JnGUMmuNdC3RFa78A
0CNFhphLPSSK9GpWmTZrgbkVcQgaDgTEVbiaj7KVERwNSpMDl+WJlbfNtpkzQhXN
jmeqf2lWqmKbpsraRFgoI/yPvSdHM2gTFGNV+zCRVo50G2Bz3vubabIxjz7D1M1O
9FdJhGhIinllkWXQ3+sf6ShQxQOl1eyREHNwpfZgoWtoxlezRfmvJhbzXZhYA2Rw
dqvLl6qwkTaXkyS0TDYZqfNj7LeUW2W0WzGd+xajlBQtYkKRh6thEWXLJEoD5Eww
S/bK+W0RuOer8cxN9Ecb241hye92+ui9MblZkRxLAzcx/wkYxCo137+0ATbQO0rT
VMwNFVJGupxhVQtvD6WWXUUZT4PyntQTijXNv0DPgVzWaqMHtFDP73rXAwnlRPJl
BA8eq6TrsRjXn4IIEs5rp9YMQT0tRyTQ5u/ckoFMINqGHObK+OsqYibI3SAcBSdr
PUQxrHv1Q3E64IDI67wh0zutZ35+74cAew+U7InHgmv8sZJ77cbj5uu7MJOU2cAs
5fFQFQpu7xMdQZIGv6cQUoxSf7Clp99Kv1exy6N/jz0Zd1MzVC6fi2GO8OyP6KbX
vUINo8uNvGES93g7REOyIeqFwbjJpRqrXjXk2IdJjsX7Je/fT4PHDFGhg0OvsLU5
S2d4lcGH4xobgPBXkt3drmlWHLJ/S379j33tMUKJ/uE5EoFKOSEmbF3ZNU3/5KL3
3jfN7+lyTrGwjfJj1qJPKkZbaBlDJd0oQ6HQ2nr7iecjC/ljrPQSpJD9JTJrxQ2r
CEeCAC38GB83T6GdgKKVVseg9Vz7VZ0zQjGgrmQ+ERNUFwFD8x1eW47ZH1n5GPd1
K6ulg9IxodTOWbtnaxAtvmPtjUvwNT7/0yyrwQYo9AQwgUG85mZWgzgP8rdaG0CK
d1tCcD8DnIK6V7WZpkUpiYEWm1NEW5T955MIhuTMqOiOO14O2gxu8T1bIw5Fo2f0
BMJ65Ee4Ia2D+jlMw8W4/TAH0TigBC/57TwEOK6pCMLBdD9Xwe08VVkihrVyzPwx
AtPoNKeT46a1ElVYzMYIxgsvOxREHkVrM+1lOyslsgcqmt4JCZcFEvwNPxylvARw
WTlx/X7Wsh4z5xFIp5Qb6VvuaAFIrJngzznVPmHJivfSz8kxpweXyKkiQpKHNFtf
YnxgUrBUL4F+CeDMWke4IiRlmTc+Q/CXw/VvuFV86/I3KCj9/bh2jxm4xe+WFHrw
dvC/4qOLZuo9kTJ/NThqJ2QH9Dd6vkXHUr/DgVa1nkkb7aDkhdyNENwh1eEDwXAL
bqS+n0I+TOpqOzOzOMYPNFmnSeV5TJBMUBK8ZPu25AYZXb0/e6s/euCb99d4G/SQ
f89AMTF/4hfgYondzVriINaaFqNhpMWj5iUFKaMAZSyRzdv5SLdKP7TvUMoE+zYU
SV09Mp3qqMn1+7Z1RiLByIeOH6hiQLT+FEzEZoDROG1DqIs9qQnjAb8Jm0OC78Hg
cwuo4cmZFXxgdjpyRQtAVjh/xoEs2T9uReX7OaOe07t7ojFj165tLHcbo4U7MnCN
vH6NLDMjhPZVNlnPB/Gap7744ZCzK4e8AzyUWUPVpS3mIMK8hWxVXDlU5WNLXkDO
3p/WpWx+kiA/s4tyeweNl1vxRS7KXsYiP/EHxV7umOUvAxsfHBtvP/fpPgcAIYZf
MSYY78uaaDRbeccKkXAx0f+e9wtnpvR8U4lnZBBHHkSt9Dex891YFB7hei/gcEk4
Jji5loLKjQg3s7vngUNG2q/kxrvP+QLpVCyTOURzOJthkZbYdSKZCXhr8SI75iYG
Q7axLgbk2dg8HRDrAoc/vNY6ronlEq+Rr7RZi5MeJn1C182oh47r7N7ccdQedQe4
39SuS9KZXYoaaToQWqsZaT2h3Xc67kIUArK1dbFdDr2rFYDQXdbPtBCf4iLkDthu
cQEP2PdiKxg1CpxiTg+ZguI5sqbyRE5w1KR8oE2jNrH70XtcJKcjwK+/O33V7dyi
W1M+fGPQ7Z1/YyqqEtZd675niqhrmiboqZx5v6kuo0seyWOgzFlIXJBBEeF8o0n/
6jKDrK2ShDuyWhRVaHS5Cc2uVP5u6El6rl5kcltroUeesYKWLRvlAEe10P8zokwz
lQATtDI1XaYsJHRbgGxXAeaCe02fyWWK4Lxus/OysyvCvL1IeawfNHKHvfChH8/t
X707voTEaBjmQL1p8Tg7H5CqOQjKowYboQvnwuPpNOiCL+fJVDLKNNPRTr2tRyVk
g/kcJsdXfN9RwhHZrosCvrulsGBanL3Yci/1lOuYbO9CNGEEc+PX5/6Bct8uOd3s
iye019IPYamOFyhDbN2lUFC3EEuCf9QLC5AwwP7qE7t1m9c6te6j3c2Re+C3rkiY
1Q1cKb1MwvOfXJDWozm8jDnM3/afiVbQMfvrRpjqwLv0jq+K7rBpLIDa3ElY43LL
cBs/TYl/R6qAML5A1WpzfDb23J+cscs2/lQn7vX1tLsspclRsa6tw9eYKGhZCbJN
fV7SbbhPylYT/It/HhXyim/mfSxnv2fYRiQ2Ma9mgjAwAd4cWFkuiGjbtKBvrF5I
QPZW9Glfw2haEQ57h3cG40dR6dMHc8Kr40QDZF9FargwV9uZQlp2khzooo504RJv
Gbj6nf0ggj0BnZZdS3ecwuA/oM1OYWHr1UsX/fOwdBuOVQg+Aasz6Lb786UmG0ki
vsfLkpT9hNvEsu/6aK/TSuHkVhdahyFAVfDitHiWFjDSpvASkzLG3PmKctyWcXeZ
7HNzAMP8z5Xak+6yC3kbrDfc/9a+KVBkZ2Qjf1JM7jlPN2H34cBJURXfAdUmUPsQ
Fr3p5n4/odQFccKiE+l3JKAbutbvYd9VXmxqaVzhVw7I2A6p+9qhqd6daBP6Vykh
YwcL0YYD/6jRRoxbZz10E99udtsEeqKzQdL4qzs6OXjAInFJ54/XqHAwGDaFQOCL
mC8pRjxF2KeGYJCjv3HSuGmYjII7htwPWsJtnc/MeuOSBzoVGUhXYhYfMedqH4yd
OSWuz3TvS21Gb0l52KYUESBpRgSe3dofcLR+925CCUmmC64zWewy+y0etJJGjQn8
xBEcgTmhNxCm2TTsiyMsDhMQALSqnnJyVu1wciBcQOapH9grSsvDqtW5/jk09vOc
hyIQPJ2BcwjjEBacDpfqwLtRuJ/2r2aNRnexHBZPtvtAq2n62qBD0IOrFIulfRCE
P/zjj72vs1Rz8xRNdG2qGUa+19tFGWcXgGB5GePJ4bIGFgdR19lsc625NfBZk2Jt
ijM6i5jVMqUJSeQheagmwj4iFyiPEDSopeODxj0GQbjXY6dqJOGLz3RvzuI8Tq7Z
EHIhilMq2Csb6WKZ6mXG0Tfx8AWEMCIsPM5uh7M5qa4Czvi0dwEW5HxU7yMxPEac
bIKCs3EyjpX2ymyDvf/fL1X+ncJrkP9u6Bd9p6J2obXZxCHWo6/T9H1NDw7u9mQZ
KGo7RrRPh2pTNxQ1Z+Bw9pnM0Y3G7aJ090eEYwVwqEBvaN9sLV6qJSVStB3VXsOQ
U/izZP5zz37we0TAm/qQiTZLDMwNgDWWynaUwXK/Zk2lzfCG6MeXsxlL3Lfy2Uwi
UCF9LOqRZbtkt+lzDFtkO3/Kv0CjeR7G8RN7NiKjddwHHwrLOGhAMkX4tMH+2Z2f
xj5E9RnRqsEyBeJ1jIh8V6D3aaLJ0t0cd1W+Dor4xUlgScBf4UaKOV7OPYD+CWfS
m4cp8PcVFhdyfcmB+ioN+FaA5sM+4f5o+WhVAU4HetPfr/DL7r5BbIV79JGTnJV2
oyMnTllLLCZJwofZzJW2ZrREG+pOR0nE8b/tJcqZPwTC6oZSfkFSofSdvLjYMyTf
ASMos/djuCgN4EHx+EEeM2wRglbidjDevi9WyeRprIM8JCHvuYIYjyV3Bc957W5k
LC8rzjwilEBLERx2DSXerIo4qZnyvBVYgPbS1wKZoVJen5xa0OpiKfxXWI5JfaFm
J0ixCS+9qaGLdbx+Z7J2Z0MH92Y3UyFY02mC0tyXp3Zzn4eC9+uhWFKwQ6KkuXUH
TpgLShSPp/srsiNycOAg0lzMbpn9XKM4FZRi7GMeeDN8yh6EZx47wlEx5DUPk3Op
6qjbueGpKC5UtiHrgE4gOC3IyOlLLpLb//ADWRBBcTdj4Kczt4MXSU+KFXM3gS/M
w9jIQ9A5nIvSfcBKK5Idk8XsJCf5EeeczOcZ1RTuWhY22SLaleQEx3L7ElRFO0A9
StKulyg3f1BvqPd8R+zVBZnc5zL/+5VyYDfN46FZ4wk2af4jp8emRXpDw49E9gGh
Xa44qW3a1rRbGZI80oHeZg5ILB2AhGTRxmZDqzVlQcJDq8OVkjt90EcwYxeBrS59
/VEZti5puB3cdLqDZB/fnzpTDGTSIBXucIH89YlqiAEuQeVx08WycsO+EW1HpMV8
XO7ZSrkNYK4s4XRlLqJsq/6OvmFsQM07Cr4z1XrSNs09kbagih63ko5hjMRXEo8D
Cd9RJgnWOys8EZDjj4DxminUhLbh95zmOJLwxI1tPC8qkxJ2kZkFdKcm+3qrmpEv
SXjAhtgdZOjeMRFaaQyaE7OVPTuK000akx/4toCPmL/O2DrZu8nP4Oy/bPGxKCn0
qC2dfBs2lTdFOr+V3eN2tymbap9Kszs4FSL5sENXk0EORavPAWGHALU9SUk/6Aor
gmXflKFwrzuxMnMDoneimESF/L2cc4D0Ti02Zc7QlUab72rk1j/93Na0TCXczPrF
rVBH/Gq9ilZiVJiJpd6WYqUEkf5/u5yD9tDlK1JrlzAXEx8Q/GYZi5Oqp38Tz1ra
9t+V5KZhTvBygIlJT2odJ5YBVAmwhCsEA3gHla8sOuPpnp3AsEJu+g1benNhOURC
aGs6snXUPldBNSDgazkX5jJ/JGQMjIGMJJzN5MUMLOQM/iiYm03vO5Zpu84cK3CM
eyHb9NQk1hck7Zy8XO/TjdG9uCDcOaoaHNCvvRx/OArE2hKaJh16zRJumfS+uBFY
Dj61DauEsJJT2tsBHHQ6OZXYtU0ZUYPh1F1qiMuAKfuR+oel7FkM/dL1bRRmiX7u
CB8Ds1NmbgZdLaiwDhI8N+kINyTvB1L7V14NtaR++5AHWYBB/YUR3TmJ1fr1sYW0
NEs+7lFnNcUQDfKtk6cbRat0+5Qrkrln4L7bbAAkvfpoKh6tU+Mk63K4kmMWlE3F
oD6p5rWdyGDyMAJoKZkIUmt5na6XVPIEqdmaj79Em4pjsrsHAiqcDfrBOsNRreDu
PN5J+bX81vRNaGLn0kX+WrDv9jb3JrMLuiY9zCzJFs0e8PShc4HQcEh2lmlRa2EN
qHOxDbPBdqf0lL4BHHGXIAsMQQQHvXmj08+fE3K4Jp1A0NuoF12Yy1caMt3UAPax
k4JnGVq6Cm+ZAOMM1tOWkd0iInlp5vLsaMAX92oE13cPu4qTEinn2kRnLUuwmiRm
Nj2OVC9QE+949XrKuVaJOAn5J7UQ20AO3osCTaxd3TeYaMersAQ/9PT4ZnrqEcnR
jjWmsVwzomXj3ZwAfjHnH9J3U1JR9oURJlC8gdv4TmBmx+uGEXvGXnAMmzlzZ1aw
a6anyZh9CP2CMVqAJqw11clMLhf1cWEdMC9pMzbP1QLl/tp0OVRcqzMPeTTA7DUS
jaKKQNKyjn3iRT0n8Vf8I8N66ERhy/I4CjmYOH46qyfjHT0r/l4L4Uhrr/HXveEM
JnGONLVsMMVRNBL44PYwQ/XoGMMXSHO3aSDnPEurgRowE8FoAfxkGejnBC7k36yn
06Git9GSQn4HtqN3BO/tzdziNa37LipHTTDMQfp7d3kzagFE9fvwezWMBKh0xJHm
LPELI4bjW5PwujimbHHg3RUebyew8ejoOWlMUSL3SbzGK1ECCkVLZ/fZQ3GLRVBA
uGLBCcK6dZO6x3pE9cphJeCBeTp2TY1i0LyYR3eliSZ9+aR31TQa87S1cqD0KjX/
yi0N5UyXfne6qQ7J8lIqwEPuyCjRSZEc7WlC5YspLbas5yrR7U86613b8Piri/33
+gSVEQN8e1aykrFHVqZ9x6a3p+7zDswrLdP5bgA3FRX7jfSq26euYOsju0I03I7Z
W3NZVetyMYz96wI0GOktJXIyb8DozRuuFKcH6eLDnn1yNraqILAZmnOa2ENkOopX
Kc7pH3MXuh2XtVCZzazWqIVCOnuzJ/rg9RCLjeuN6HDKr/i4MQXDGT1ILz8JXWzA
E0xNL7fXeIQycd28u1bQOTw0u4ibzKTFb0OOs2xeycAwSPiHhs3IRiYQOMMs9rY5
0kS8CTrKlr0Xzu5KAgR9TQh0mZ8O1VMRRdXHkhb1uSwQgTtxhDCwckZ2k31fhbaN
CrmZi6DV+pCnRHcT7qNoQuGpq5BEASiApsi8bap13rA/TZazMrzGZ+yVpkZgWNGA
mPsZ+by9SqNOBclFwaizjSkdC0cYvVPrGH6bfAZHotSpx6YGPHvHZYIola190Xje
PJa/l7qmNQTTBX8d9VLGnY4pFzlWZQU5TJvDo3x1rHuhlZDTqIwGpIXYYSjrezoX
OlbxDVTSHXvyDH1TIdq+1+pCX0cRj/S6XQM3h6f9H0eB4DiiMCDXATldFALC14QX
csOaY82om5T1o/o9TBNOwrM1SwZt00w9rdcZjfIMANIFgfU4rpMLV1S7Cvq0M88q
42rf/01ddEGBGH0PS/fEZJY1B0A5nPfsK39jbq4MU+fTuj+cVHwyorUJi6gr355T
BPlxoV8WyXfLzJrZ4906D9+IJypUMyyDrBQ7/LagYVVXHYRVZ7RllG0kW92/TqI1
5r7m/yqgG9DvsEoAlSCnphekoAzUDA3UoZvEwdi/IzHDlGNyAYe/mVxAHsW4DbHu
P7czztt99p66X84s+pPWL2UTbPrRr+Z6X+Sh+tftG7REBifOx6eikWuEVskOe6Ja
ZsHVRWva9QKTFX6LYdhkklzsU5v4ZgGwnRfXYzC5K3OYXcp+ZrE5Wv9jG2uNpyJ0
mWBwQjqgLG17uJ7ned4YG80a8U1yXPn2rbifPoYKCb0XW1FFufdo0Pp2LbNDj7M3
5Ifqa9kOY5t92/PgXR5Ubq+C/nfoUFd1eAeP0BMYHPdKDklsjIEEsDXS0Fw/CM25
gMN6nXlfIXbvhD6lXv7r+eeCydMS/NTBob2S9tDMXuw5MOQ9AqAWmUoetc7beBgU
u9mZuvkxEtpZUe9/sV4lEpkMLVDb6A+s8qacu0ReZA47Gc0sq+HAcBQ2GskpI3ZK
124SltGuxUKWMiYBf6i/xmLnuZlJQQ1kwGVFCAW5d7sUnNlorQGFVYhomqFR1g7D
7pPs6VXe6pVcvD1COzmw1H2D4A21/DHAXrlAltOZIhs1SGutjmud+tpsLNN/v+Td
5FoleFZlTgxIwxJ2pbG+gJaKwu0EnV8xk6Saj58tDW+WwYKTkylAF7as7pnCbr24
QXazoI1jg7ydm0BlS4Mi5oYLBHgepVvXlsQ0HesWaVuQSHTHJG5u6XQsmxMa09h5
85xeYAgh73v0WKSkHu4ZVrxLTkjwz90LSRk4E9CRiEsm7cwlETs4u55a8v5CHnNa
59lGQo5PTP08ux2P68x7uPjfsYsFC7zpWGz2AwzdKTEsnnY5Cdl6eyFudp5CieSL
3ctCWRAN4KSEr1VFhQLGiLOX9jmbw+JjS0veCIQeD83oTNKcCLSZvWAtx4u9vAB8
TsVm1omfAFYW2c3N1yjdBYLWYgwERulL0wjGwh+/NNfWAxAcee5c4J8epkiWlulK
g+nrd23RW+s8MVyRFxq/gdqai9/oNRbrDTPV2pxf44NgWL6t2kDQMG4h1D23XT5j
MEQ3GivTBLhPxbYMYD4QmVgc5Ut+Z7tGPmpFiuvYR7Bbc5xZP2CU9kepJFVcBAJf
kb7eRUvy0SUjvrS0AdBeJE7YrlBntow1ldwSegfRsLg3/H9s0aX3gHogrlBcG/m+
l8pyYoWiqV0ToetmKwV/JLancT5YHFYZcIRhGGaqelkVQfF704lEkcW/wiQ7+ztG
vp6aa3efeVaIYctAy6pzto+vVcOUxpBPMtq5UfA+k03Re0CU869MkaQgXHsi+x3I
/I+7iE+GVreRuYnuLO3jkKj+KcAHSpEuD30T72/TSxUKE67tpOPM8ZaACym1deVg
3T5nc+sUfp04YTKewk8raJ88RwIbwHAmAX9Ipf+kGufeYOdZow5LlAFf/GntVH6y
mOfnbmvtM9O2qKJTJIlabWT3gImqITKNVxFSHYtBQOElxtkxZSyd5Cy+/sywwXnH
llWZTeqZc9aIc1b8QFjD1/DBx1yZK2Xr1UekEJRjSIKoiniDjX1DPirgVMFkQSO0
BbQ7PZrifpvIgFca+R4ovF3KCy7zoMC5aJSmDKPrPcWiRjTawnOGRIk++zWi45xD
y0oy4SkHjNFSb08pqcGHWPzNKw5cmfN+XDn3a2EqU4M0CcwoHIHB8nBg96bCVMs/
A/TYodrea+SXkI7ae33n1QHFFXqthcHxkI8ic025y9kztBsmd2mSnHy/xtGYiYKd
0jRDVIFo65kA0PNDn7S+GMkDRMU7msaHOtZxA02jnAnILmBAM7qq4jAoSH3SZPKn
Z5MX1pXW7Z9TwwHtSkpbZG+lB0lhQnxz8ChRJ6X/FrjFqrYL2F9DGf0p3oWkbws4
8rTcrpfqR9CxwXHe6xRJUfQ/O5vfmJJ2XRp6gqdgmyIXn1MR4ghXzuTztxMc0J3A
sEUxlGoEuv9U0oDLgM1VM7xQMc3a1y2OxD3S+XycgmCWeusuAiZDVghhlbMtUY3M
fkMcmGljozbQ0GgEAXVMKhhBnXeXUJTJoGv9pYakhimSLsAaeABfmh1lWM8hTJAW
9XPRMWffoNMdzy3h8gDQOXcRyPvtBBfZMHFxcfZxz4ZOZXD2ir4TRVXUak/2adqc
lI38qjzGjV7X+OX78joaSl5+XJC4Prl3bbL19tZ+L9RjST8TSqaMTQ/eqbUVlcr8
zGUcjNQvt03eWhtJBO1mKAFNHxxMbnpIKkSbWZQGbAA8SCeI8MfnQhb9OhshxRse
yKZCkEiURcxh19Lo4C4yv5XHcmdAHL1Us9MGmwkcH7czZPHABhNH8yMz1F2DVLP4
vuAFWIlJyOBk16FV71XqqxSTIcpQs15eXAyMoH8P4t6oLxxzt3hbOJoZlPpLxjfq
JIX9pE3mGvdneTFgG9aLJYaNKeotbf4RLGf1Aj+QasNstE1gJjBMreJ0CXOzobeU
LdoRCtVADNpe3smteVCixzXbEaIgynhft9SCf2ghuhXajsM79qSPvf9QIwgktffs
2lvtTCnTILVjpX8ILi2Cb5M63oizeV05dBV9xzkqIUyW2ItHWeKPVt9OHXq/x4sC
YA+Kf9ValTOK8M4mmm/cHWD/fypFnqQpV3mJW1KNTArTt0EUPbQcLgR+sAfqmaFc
PT1nAAAO0YkjaJzinWsNztDbkLbGZrccuBr49EnueICR20wDdP/BSkLeIxQnkqb4
ZCR7ZnKU0z6k+Q1FuM7zaPB0H35ueJUu7efvKwD+wwCpitJdpvI7GDUeBUYlHo3V
V6HsrWLrRXH1mblISsbwpqrCXtEi34q85Px40+/ARG15+s8ExZ0JA2qX5Y+2WOUY
KKzHscFilZRulXAT94Wb/xiugL/KWQej/X7Wc+HdsfJY2v6pJeNqtQhBlWvtYS9V
s9lhKC9OokzmxSoW1XdcWYfqqMWzi79wh0FbgEllOn8oOv/55+GRqlfnEX0KxEo2
4WPKMwRmHmDZi//iLrVRadJj0otGMFYQ+MQUTnosrnh5saBPkxpe2o0o33Xh3Ktt
uULO3LL4bqCsPXZXiABppo8PHTPWL1CkQrPRor0PmkeSh/g5z8xdOU1P5vO9EqCy
qgFH0PhwcELFhSoF0YeZQmM2XBHNqXVBQ50Y32F8BKGMrKQtyktEX8NQydULoWRx
Z6fOJy6kisu6wDHRiabwyRPphy14u0wTHEYcSg+3LeRzYfJCtyCTsppqPEbrfpQF
MLUHzMlxJX5CCpPFprsuasUgzUDECEtz546aT2anffmiuGeDA377GSXTAQuUXoej
Zg1ioCE0eJXoTfB7aIzZ9rDZkUFe5CDHEsn6fan5svT87utF6nGOTIAG/NMuGL1J
NFsyyJLyE93liEdr/hqWSCquoN9KTCdwecGMObAaSEy5Ina0mSEk+wV2bDKqq8tD
YbbF5MdadEVDUkNKBsReQAWAt5sE5Jp54l7Q452PdsYWOZk/GOiQvuiFFOVie+8t
oiWyZXlM/S/xGg/Bw2bJlc7YNvT05Bb5muBNNHdwEwi4MtlQrsDk7DssIhspPuTo
cnjpD72rgnOu0oDxCBiep4EvPfAWkVJgp2a3TrtuHydiBKbl+KJZXg+tcZXRZ79H
kmr1KRM1lq9bzjT/1JhC53EHlyHWfcPSmInMvWaF3/gBnptTaNbyKgoWj5JWOEQU
+prqzb9IT/MM6xqUa+N3zfY/SAjj6gc13C/skpHT+QmVe4c2ne9RwIpb8CWBt9ga
CGOAlokjh5GYjksbT0uYG4HM/xrxqy/BsR1Hs20tQSiBaLcUEuTCfZGWjlppxy2P
IFCgH4TrpXrjfJoAdMvZFI6qd8ZqcYMzcsoU8ajaX3rWv2zjLL6rtLTmwJVe0UpN
bkDNFAGvcDdEx4TiG1HwWWvAa1MFG0g62DptRb3T2PtjdQiQsmLPmjX/ZnT05uBf
mQIfej71gSKkTtXntqlF1sfw7dCJjd1bGlc35hY8cqVSDoecoRdbZ0kGOTFtX9zC
uPAM8mAEupM4aArFZBa+NCeqgPCULtKISGMLd84cT52DPzxxdPBu/qrbwkCuwvoR
GODBGfUfZXKFgq1LIHKH+okQUaVvnD6oWoCxKUNYyvdHFWuQ7yG2cd0XxhtrNKUY
078EWXiL2BCeBX6US7Cytz6ddAr78iMsiMtkjSEyomqPY2ftIBfYXzhWyFrCXnOu
SlM3U7JPeVWxf480VQsY54xEpu4Gs5DpF0nOH7RYdxMJKnk4qK/wKg2CLeCitwiC
kE3NFtftep3OzBfWICkWmjQWrPQ6oYAHAbQdyBUm7s9kx4V6TEnTQacSmeQph6eK
wibaFVOejQzZgZIm6EIaSiYFaeod3qeIzt4SCrpmNYDbiiF8RnsPbwnL1x4+uClA
MsvkOR8o987Y/Ereyp/a6XrTuqMSxZ3H5KnAvmPD13vPjYEz/JI9KbdTfV7JFHtX
WUwbsfLeXEe1329ePfxl4PV1FPd70R9Tq5fAauVxipp1AZSZQoA9Jlf3qcgGNhSt
3xyzDLKkZwFJuA8DaXIDpTyNSXuAMpTmTI2USVaxzoemS4W2+I1uE4pJ/hyPQKS6
HH3vuw++osp5ofjY4f6MYMfFeN2XfowOb3wCgplGGlJl/Sc1+CUa0Mwap1r2NVSB
4tW+yWljHChjaSSWibIv+gPAEgQDjLF+tBuJCKp5sZ8aRLRXzgLrsvx/NbF1Odc3
jo4yIsU678HkwXtVK1nSMnQJHbNm7C9x56eqDuE1geY98xYFFM1o5JUPnBp+OoDD
vGPCDtjWg7K6ys7iwHGjzt0b4+mmaVa6JeSyrxsi1l6rnoQl70ve9lBx+JeB7tln
VP2nQS+XbO7hOZwXYBkYK7w9I34M878mGsKB4HUsO+gPoyA8UMI8DCeuX+OsXwc6
yTPO+PlRNORPNwMy0QiSJGRnZRO+yJoHLT0jbviRoiRYqsnnJ1BNhdieCUH3cntg
R27kN8O0TX6LUzRQpoVQG8xkZOsYsn0YhaCw7mGVlKlBFnPNh8+QAFcxoH+vcagH
fuf/cw+3CITgBQySjn85xuY7Toq+ooqng8j2JUDyJST8jBEjjZS0fAMORJunaSoP
pmSYrqK2fdBNH+qZv/kGNSB0wI+sKdC/u72SBM+bA2c5rVW8dmBzgH+F+JWpvA76
JJlxQFUGGh07/DSoBliDoPI5AbDzDRDy1zCdMIggG0cOLv3UiIKr7KheH6d4v97j
MmuVggZbr0eDJX9N6dd/hYItj6Gwy8uM/jN94VlKe4lsq+2S5qBmdvyK/AbkQSzR
tbzma8aLSvHqp2VITtYuZkIzVU/mBALEN5KI0ZFUP/oavKET5pOnDrOOUR2NA4rh
zD0+XvhK1Tw7Tu51SQOL+7nInhRTUXA4KvsABHbQZus1y+lWsOi9UtBaMOah94pK
R69obmOEQiFu4JIKE/clbF6za4INU+BnRXSy1VClaOmh1md7Ouuwo2pQEc0ig41R
EqxPqQVzcsUZtGAj5w0/1+VhasU3Y8iHB/o/SbQq5CLexEkLfbiyn50+cupfCkec
PYeMRd4iJ3DPOFUYmK65W8nx42YB+qinxngtFZow6+Z27OjIuWRVvLpAyjq8ofpe
XTt7wEBDNET4VOBO+xD7XiT7xW9LsFdwgjISQnUyt1SRrYTdwAHs6mKVJtASeMxD
S6VHq888jPZo0BTZVY4ymeLrej98FHb1AsAP963AeU9C0l1nGR3lI3zuq8jUmuom
XtppG+nrVKozsCroEZRzkFvpclwinQg4gTuxGXsURFak4TbO3dDukS3jSdoKuQZB
r4Wx+hiTYSM8a4Y8Qvf/wck8MnwJs9E4Uwzv6o4L+s4tEWhXLo+C6IlgVAkMkJ9H
2fPjZWqPfZAE3LeQogH3e/fLBC10KHXg7wXHznaS8SEiM1B2ejBR/iauXOkufpq1
DNFo6GW3tJKimWUKWPA+0wVSRHNogtUhY74ZIqaPUoxuVt3muHNeID3a7IM8yjLN
BI4pS9tKumU5byj+AB25dy9Gv/6bwqA0LZNN4tI15BJ6m7GSqPhIPkKixGKQ3U8B
kmyHNrBPGi0xiMyXRGNp6lrNifjrCUIfCT+znCfm/wIsqsEuZwk4mJXhpm/JzITR
uyobYClcmvMMjEMf4Chq/YZ34dAC6N431CFFkTN0bDWTgQRrrMcKTk8AqKdjHIKp
UEc0gv46KqvNrxLMUivXrMnS72rsPUlUImimg7CAjuSPAwMkgB6TPZBmJ+2QVHLN
sw0GcGRQCA46WsY9icrYBAXq+ujO3OErG8GOAti1lKR5/SAfeY0LHTbehXqsLODb
UIeWS4O7R8GXlXgLIaVTJkcVj3ZO7kBWXssiiMQenJwr0v6CIQGMl5rfa85itBs6
PCHEXqVsSwyZXZnLfosBSS+HJxaLqrnEv8T9JtkVCCbpTUMNCcy/bjAuzFmJld1Q
XPAnTrLdVu6ZwNSTbN2nUWHSsA45S88ylvHWPuPk1cE8rphwhL05BPv0ybKWeCc/
IQHpEudfSgYS6GJM66T93dM3bqwNChYP9YDBwBBZz8FlIvFP9fFrf6ApRskUBmgk
4lJJByAwMa2dULa13YfqbvhRlqdT+Qh/557qHc5KOgyCakEQp5ae/D0PPvTEYdC6
mwsXYh//FyW015Gbu2Bs3Bag6QdYJSTQlrVoT3x61iBrix/t075mbK45htDEGOM+
uWm+qbD695Xm3pFHD5sxHE2LOtobO/tfqoWTvD8bkHu+op7Y3X1XmGgNOEQelnrg
bvNhCfoGSncOKphg6mf14pV4TncM4yfqgrDxGs2hf65RJNbUnsB72FxIziabcnyg
DCjJNcsOFvT6TR5WBl5niz6BL5a4lVHoU18Y7A/kprC+Gs/VWwuoeB0k2XSTL0uh
B2kxx+sYD7DF2KwJu0whLHosLNYz4DUY+cg4xNDLL2BsPTlBf6KEr5jimWDX844W
lcgSVKo29Rpfw8ai+P7ouIuA342MoLtw+ZuV4tFjVZzwnVgDBAYB41hSH3JpgByS
GAhUaphOdU1nCK/q9j1L0xw+HRVK9uDIXlrizu/S9GekML+MK079xJO8Hwf13GLa
EPkHlfYzYaILwzZMIztw0WN9G2qWRpbgWqKy0WU/gWbCJLbx4s3jtB1V6jhb6flw
Vcx5zsJ7dVGlO9uTq3neV0bC/birL/GX+rfWg7axtfM4pSqnhkitSEPdrAlSjvmc
nQR+FUJFj48XL8Bmt9YtRnfIdnp3EZ1oXvoGb5Vs9GSSBNR0fgUY8UQO1r8HLIHc
dnHZ5B8vYwEyOutbhKpbSY0Wxjr0audazvNuumWoyTjI20Ftul7RcsCPzNZYJn8E
k/hMud97GFcGisvEIQVBS1Z9EmKlGze9+LLJwMys4SkgNhnB1903EQtJD4excDJ/
CWXwFHlh3290iCIJ7giBoNPPbZsTwBVMmbYBMcgV11FFz68GzxmkeRLh6HZJ/hvq
iutokQwWJb1NTgXdOviPP/2TyLFH2cZvlCC9xU3m6XrrcRHECCrVIOyg2Nl3eNSX
EzhIlFcn8/hV0qYK9Cr5vHWc1rnV+5H1SPlMXzx+QGNtEacRxSLmwcCo25FKIfyy
wdqHYU7c/3XJYe5PZBFWPPuq/NfmGAUFpy1jKdBf3k5hx0BDPBLFSrnmwOnirpSF
O0fqW93Cqq7eRgP3/eyDnQaZoCbqIyycIzjDPpGt+yRuh5pPEZV8n4vpMnRumkm4
sXOA0+o+MUUCUHb4WArWZpcO4LQfGAMjlAdlpXMBFrzN0sT9aVcK9BB691ibiRn7
CynwLWpqYgQee3Cg0mN90c8HGKUmNYr4tvWsgUGd5fvradFGOFF7mOyKkrOTvomd
l/uu++26Z3WqiDUGI1sklRxCwc7Zb3ogehvgzWNjNPnghmHOuxmN+v0TQs35V029
MpU8wXt8UaQRRoYDBl7L1+tt4l1OAP2THBF0shI7SPt/DwTGDvxkdaOEZXe9v64x
lj1bIMcWqkVAsQqYiDTNv4+o9HbiN/C1GbZklaiAGgKLzwnK3aSh8KxpUydsTMKD
PtPjui40wVaGTNghiXZOGzW+IYk/hhQmrJ33vGvjwgVfMc0hY2dhbnLyGapdAZtC
YqJMwXCSIwPbS0GL7bpvC7if3pdVUetj6YIfEpZNGD6Nj6aJ6Z0B7yaWwfTlRsns
CP09bjxR+Q7i3TAd4v83lHIlhmUup2huouxWDK2alEMrq2L1ATo974EVnW1tZDkT
G/XfJ5LaPaRkc1HtUaGdEb4DViAiwx8fb+Qh3nnT8J1dhSVShtbj9xsEk+hK4L5q
l/uQwEp9ex0FvSKQjr1C68mB/kGE2UP/gY73IeNCJ541iU95vyyWmr2WpX6UEV5Q
UBMB4mcXF/MsMzkz0dMtnzSgmwq+GO2gcCh/Hyz6s5/o3Aq190/IAanlWfJ6caGQ
mbZEozOXnZ/5OrkWp4H4Z8M56N5bxHNgD5dr3b+DpbZanGN6DjD06/+WUT6nnL/G
twyZfQG+ABRjwnR+9bVkCqK8ARtasKw5T/yZXPDMKLpje8EF/J6O5MRmIe5rIfi7
tGesLa0WnIai7IScD2jk7GKhxF/7Y9uWcbvunhOmpPkvje3ND0M3yNTNxQ8BMaZ6
EmydhJwtEpK2DCkaIgM/s2Cl8Pmweiq9VUUEm2j49HEcqk3NTuQJ7QdkeduIbxMA
2EWMdU1LCUG9PdkbAZCjvPHCV60t+LYVixreo3Lr6pjeyia3RUEhGeuMkKKqXEek
qpwO3VyNAXJT50lFKNBHbBYKM7wbdChdy5uAwRpsTVpKrDQRtUwdK61nWAUojxPx
LozZhhOxzTCPzn9kEI+qUwZtBqbrnifLmYX9N/7XWDHp6MyrqUKZTTXAqdX022QQ
b7g2bWjoOIz/DDFhzamu07rXZFJZPHtGw85xpRc8+0ljYUfdAE2Lf32Za81Xozz8
vp4d3kKSgf9brMXdOH+C/kQE2ofno+h6GHT9yGMwFYubOW3NRcnDmwB6FP+sqNni
pnOn8WW1cbBUcdgewdpMft5OMsj/jiZQ/7nxLtjIzWPko0gP9FNcrRo82jm1HShG
2Mo5uV86r8bcS/eFlUTXdbCMPZREtncWUd8VCK/t4ngyrztgM4gRGZEKL4yFUWNc
JqjmWR1KQyDEaCzLbHbFMYVfKfjA2n65ZJqUcVfK1ud1C2pKApd6DCFAIWvtH0Lm
PNRApfPthl/XES0jm1yvvX3bYkgqyIQVm7b/qJMODdasUxmGHEptf69FZKmXTpNA
YB5XRezmPFcW9oT3Qm7av07VmZVoyRGJqpjOqLAfGjpdEawQBB6p+feg9inXrEU/
xH7ALALCvJwX6eBMKLhhQmhiPOseKxEPR1BvmZCGoesLaTkFoyfbR0oaOQU4iGHT
Mhgkqgyf3mimflQqPLH5FDCHzdP6p3hEatG/+1ztC0J9Wj2vDgsEBVWLb6HME4gr
OCFPex8JSghQ3CUz1BRTpsBPUxviH93lZzWNo1PYiB4Q9w8Cdk8p2hpPZZ/DvIgp
o636xqP8wwUEGSSLBR1rqHMrrycdE/g6Diu29IgIyroUoB+ibCXx9G8fvjncUByw
fhDGYMVsCyZYVDhX7VpQPTZr72yscsBIdUGNJmg3YnCjnY7/j2Ma3FTYUyU2SbFf
sVJJYI42Tv5eUNFVxG9AV6bjn8B6nFXA4Z/w84McCElKbXAKryfZ7Q/u9eHJYzoT
odqMH2BNies4gnPS/z3AcLK6NOnum78iCY9QXv7QEu334Jb8t1yV7OPBhwUSYS/N
YhLDdbZEUoL2PH/24gKmmiRGQkeT9i/UzNMaCZWvAdKf8L2T8Uwghe70nKtbP7BD
Vauj+052GXWFtuhuEKlmW1R5RqPsmWIawflFRl3M0zRVEcUg9MhPhLTRLnlLzdyz
WPmHSXj9yeMq5+CocXy1kyubIgp0QHVxnZFr+bQz9s0sc2UUT0ZmX95/rCzrE7DS
KPYehWI0xvIj7J+4PwF80aqWX6/6OlJSoH48JSPSq6PP7BN3qpxTwgcFcg/6vvBL
y+0i4sNg57SSgRO4AKyiaxhgRQvr9x5WWsJ2StbDjLWcvGMmQHeA99EciDVsb6Tj
/www5RWUeMEOpftLbM+VdDJeMoCpO57qtet5FGhC9X7D595QS2RWXTQI7m8cYqyV
FHxDxQ1KeQRDSGp18iwoyxXiW0BgFjiFov5F4ON9diwX/vGhSYF3O9y5JO+83qfG
oQWWOxHh2BuiVSSWZmTORWbKv0TleFQ78gbzUMk53vo8G7YiTnWeRNh17sp+C2yH
FQ9F2H0riLw9DALxctpti413uETOYuE/WbdDA+X+rZ6dOPYFmmsVTFiZTjGKJmeX
UoiRtv3mkb2CZ74C8oeE6iVZOy951qHrxxrQjaVbfYV4Pof7HL+L+DqlIt2i6WIb
O5a+yIK+YHZ7LTnJvkwTctAtUGCPDgksa82nr9xLru6r8z53qEGHIeihu/pRVJz2
Y2cinOp0xxcTyiTezaX1/e+h3P69p7V/aLjb9ztel0N9NNG4tvJjGlQCHJtNsd3l
PGSJlidtfi3xNFhiShlLkNVD4IfvrP6KFkacRSFzGt+puBgE1T08Sc4ZKIvu0HEp
GGVyRT0pdERjfgZj+pJVkIndaB5asqkFZh3QIl1i6qTBnMfHN0jt+VU5KKBn6jtO
oiCimDFVC0rHwaA72XDz9UiIjpSKAA+XSbPgd3X+8nuRmsUaaVMNQGIh0ixyHZGa
QfCncyuHp8+xZJt+4qgQFdQ/K/M5CF/iXaHa3hjjPqiRgvJPOkz/gnHqeO8PdQFX
RhB4EjrFBiB+PbJKom8faz9PfiJ9krys80Oji4K5FRNHd803vj0NR6vjMH5cLfTc
UUvvZD60kVPhbw4A4fQzy4BvcqPtngQGxQADcBCgMLfz+KR8dUEJc9deWl875ozJ
sFMy7tq1c6FpJ3CfohVAsLN4NWa2h7R0o5zgsYvUw50+zgd7GNCw/eXgRueKl7Xa
SD9Su+vdPZcHze6xlq1d8tr1EqIo0J9nEFaQJeYiOeya7XaCAFuPPTqEEG+pWU6r
4uMxq6/8CqGSjIijxI4aKpCadNjqNfZST3ocs9nuIkExRkA/hymP1ECrs4SbxxTv
vJ44Is16w/pmfvLItsKKN4RfOgiUWJ22YaHUm9BPPKEXAAakWEWokH4nxkQyDQo+
sMpQgNRxwGAqjdkpQxjqroB6l8Sa2del4LtRZdHuj43tLk27ZdT+HQ8r/ekYMOVb
DvbZxwdnGDxLueUi1musJm/TT3sv2U0nCNXhNK2S0d7Yvc/GXbsuRGQS+upoxqNo
P9r6qozWGzxRD7IkrFC8jb6mr87Jo3X2QFAZeDlx4bNhrCgQ92gL0j/ylW5JTzgr
K+Zak05DG0xn7FwS+JZ8+YY08/Ph5J3fCxaoLoZ4TSOb0GUhRLAj7eXpQ/WY9Aia
wrOzGm/Qd4KUnssB2UzUmx9wiqSkbV8Uz8V15OWmBsp51bMSTPP7+EZpmwZZsAPe
oi3bgXo7h/9gSYDzgZCMKsjC7pTEm61eH2ltkbV3n3AGu6K7sfTlGlx59E6XPjOL
rfuoQoxx+dTNctM9ScVfCktXNtN+hRiITfm88Hcz2s/XXLQYzz31dJydxJn9G1qt
VVXUQUnhhrrP4w1S64FI/cLaK53+EVgtn84o5FcuXi1kVE7n/475zTb8kE1zEuTv
YG5pSYtYF6kjiTUqctSr4zP4bLKSCoS63wsu8HnRqOyMhAnwW+dA32Llq4UYMfzj
fxvwBYBpryUQOeJykPIimw5M0OX/av0grA/X5dn9xzzibim0Z2+shbHJL5yU0I4Q
lPfU6A3RHm1O9cldbl1eO1hjfGjTGy9+ZrpxiwlyaeRwdBXLN6LsV3f2t8pKUZXD
GJzpTh3VEhjJQh4e3DrUnDFeuVSfM75suvAMey8meuf7LUJuQEaPrmtES4n08qmf
p7cA2zejqd/mvteO636iAMVOT3HumT9tzDik6kRMsbeb8Qafbx6ys/9lwPLKXkss
+l9BV29O9iYoGKo7o9zkInX6s55JCPPttpXtpYJuS+s45A0tpgK9vwXc00aUvler
0fmzlw0uuQwB4vApIXg6e+fnGVy6N5Qsbr0v4KSRe8/GruqwRhmIm34Yax6cGO/D
8V1727LrQZoGy8gFp0W4DavEAEbAoXI3cLVxcRDry6x58mMu3wy4IWMOxOnslNgV
QN/hqonnmoUBZivtTcYpvsIzw/uH3fr/LovZ99os6jCqOom1wfHH3/6vAWF5CNcg
b5T9pxbTwH/lCdzzwjmUx2xhOiAAwqgG3SV/WF4GFkbZj7GP5iRu8Lt8jqQFjiMk
J9EzTQZloAkUGDXjr6oShjcXjiggE2wKa76ohvo0rF69sXzUz/0HUMqPtJf4l/Kn
uEOO7xjLDazafJMpIL//zGY4hWhX4ZP9E7wsTpw71tSI/FjGnsbPSXDVdvnI8L4K
tuMWh5oNfxuw3b1zYGptQUTJdPDfPiLagNJSoNPetwKvl+1L1kQGXbi4wyodN/B7
PFA3CkbZLZHSX+8+ZSVmcVBBa0jYQN3U8CRDi9N8T95xNP0+9tYB2ng77Mn/FQZ1
fRTLMe38scAIRqwFWqclzo/hLiuKJHogLWlXE0B/6OfeDwKQY+75yHqreOtwnUd2
2Q6aeXSkllf9gUNm8qR+hSDU+vaUsHgUfCM5UeZCEm1blrDFLli9bwbX584h2ZJs
2hiduFru5tzhdCByrAMi4FyHZTbbJ3prcUQXjPbBvhW3mir4p3jKh5rZYcj20Pk3
ts9WknLhx7F5z9oMzBFMu9HIKWQfz/Az8tBhThdoJ+5AqApA0JydFxYBmB2K0OuO
Yexxukgn+4UOqaWQh2eaEx6954KDvbyvO3rcQI5QUFq1xAOYCuMSBgne1dJawvP0
AnNwRfFa/KMPOVQYVgO+myLcJjB1lWiM01fRz9MF6A5f70haJcCAtlMXbrc6Qv6o
Da7F02xmMURGaeERtBC5wyyJptRsa/GdiOmhZliaP7KS+IGHg3VnkCaTIqiAhLHc
7TI8EQg5LTLviqdSREqXQoabVU7GZItHjk9f/jcVpl+Rx6iA9jALSi/6bnQuOdlq
AihDuIUfERGoCx+mocIHjlK3BIaf+Sx5W4+wrUBCYFWB4V2Z7SzziajntIOLFsNq
+IfuVPVSADn5d0iK65eAbdcH2fVwhCim3KRwuHRGm/h3Kl/1P7uCMqa9ky/9ObFJ
hJKW6qQcr8tgvvXXLkj74fW4Qm/fBo6XE/CoTf4yAVv1wXHlLepApJP8l7JJ2F92
j3h3iPgz1GQ3hE5b33vzL8rBCE8OsW1oV2s8FYMPSv5SQdvwnYY+JX6J4M8w+9tQ
/R1qYqS9rLdek2r54upR4/J9dpHJkpl79lXYOTJnmdKkynkj6O8yUX7zsEOMIuYj
02okpoBBsTqDr7cR184tBU5002xJ+fLEGtwjvfncs9OhUnsbahAAMLfKJ2REKdgT
aaoq0LEYR3Pgm1EPcUGtupX0hl38rCNvWLds5pY3+ZUMlXAr5fMNlfB4MWYOjM+n
5E70EgmlrJCmRkPXxH5CVSZ3yaqrQzO4j2v+RarvNjv0/WSCJn+pabnL2tY9ja/H
TlJcv8OwjZr/XOos/lbGXzDKve4vHXeEawvZjwzt7FDCc865jm68gww6Jsol22dT
M6BgAh3Pi4RKB6U8xVRFNoYtxK3bdClPVYc4KdpRjuHiRctzmpjkVCWDp4Xf/XF8
DPd3ia5dc9ahzChC57VK4Mx3Rpx+ukgbEQs74sHvo9EXHOZ+re5V8B4/u5oMZcCy
N72epmEGspJnjwQ+TcqIuLEJOlApNMejDGh7+kLECE2OndcXQp/hChAr6/Hc4R6e
d5AxhcxE90aVM+7cL9xiPdxvaSou8hP954z8adICC41JlOT2zdNnCo6dO7V7Qudo
RXIKGtsN2coaIfwEeawdWI/tfBM6iHSnRXOB8czwWYmc8xhc5LsB/fWvUxkqg5Ul
se4ORg/QRl5Eu/Kud09lO7BmExumhApm+dZTZPx+OWg4AnKGdbHvg0LPBgaiV66K
PDnSHNV5YglJRvKufhaY4lUUYW7kkmK3EIlgHTFVUXDGXt1g3sgGAyALN5VrL5uO
kqRuOD3DwXg4ynrusW7dWnTGalcL10rSY6kSJvDFFPjt0kXX653V/ry3RErwwi5g
qgw9BmWAffA4AENm4fCf1KzAjNAZTOVA2kGgSNoKWEoFQeg63PQDI7Oh7a9j3blZ
Y2glggJkb2mZpkowAAydWdNBj2i2PE1jnahbqjkNmdyt2HxFTHEY49D+EsipLby/
vmrf3Mb8azclVh9TL3OwEP+8SPa/PQxHsmrEAaH3HbUFQeTSpF8AUB8in8o1XyN/
DmnyiQBAbwc21f+B5KkLfTj9OZ7bLdvV6jJHoP5GzGhjgiQibAYW9qKBX0D1rqfn
HwzLOqdPLqAIlcNs0Jc9Sq2xEbsSZcpWopl6CPjJ8QmTRxrH4MsY3neNiHZs1tQc
sxe6AE77yOboi8lRTjTjtmzuMxagVzOHpqEBxERHutwvyQg+iBJx7bUJgsazneCB
CZ5HMC0T3j2asiWA2DlLeL/4rKDM4KwiR4xVudc3fgzTTzWRFt937YprQqENImFM
C3B5thUW9NQVNF/s6aIgOSraq2BAVxEf/CT/3Ml2YkzKmuxHBP1/Ki1jGA8PwUO+
wvnMxzaW4uvahbbUBbDSlczl4nJts4GKR+RMx9qp3qLV3Yu3DDKVLbhZA6g/7sbU
4IXS0xAq/j8AZGjfmsot8MO/ZAZwMsbSC37dt3UjgjrE9WCNbCk1QF5v21bH7ajR
sR09SLrMCBPYIjwffKaSBPI1rVgjWXJLDDNHVchkJPe3YKXFmISC2H72itNaHl8A
UYNl3HhlTdNrU5Tt7p3mVO6msVE7EXzvGluZQopuYKLa4ScnALtD9iGVOfetwArs
9d6BxBp6y/KAa4bwWffDGZuxP9W5ecQRCrmMTfpUflSmWN5+YZju98hNZI69/huM
59M/KLvkgkgWjWwAeojoTCnrEEMuiyTV2yHQvDCH0p8ZAkeHNWG2zuY4SCXHTjuS
cyKzptLncbYcXy6Eyws+2TL76yyOV0i8BjrSNqVjheEG0DAoAIG9DBg85fL1r+Mh
zwmSh+YWNQjrCbPDk92TswEUJd3BQuaUUOxJ7o8ivb+ZEO0+RgOXraxWEm1t87zy
ZlxOxh4fFKOu4ChM/sJh175KM4o352a0iMAWtZ3WnNHIEzcUJ7Sv36CkjzGFNKUG
MFzMKHLvZsPCbpFPsv+ukpfn9HVNQITbYekvXDgH+VWxI6apT4OZJZ1hACgzjQPH
Djrtn0vwmqm0J/PI604oFXqgTvWcAmMOq7X3m0xybOnClLP0vFaaWjoRJijYpFNb
4K1ugHu4WfGB8Nkm8pjy8dub9KqPk70NfH/LHCu7EvNVBMfFsZ4Go9oZN47mL+nG
9Pgl6NmErg4qJCrwEeGiiMJwcfsazFEH1kI3UjrTzzMLr+czhnyzaIG3iYQSL2zE
TcdwVfsaIrykiscg7ahCWVBHmRC3hZeGs1ia9QAzAIcfPt3Ys/NVajlc4OXkk+lJ
4oGUZk01Me5lJ82CKKWFuYKf5Kv/l7mk84MIsezrmylTHQXg5TFsyyHDv/nuxxP8
xIZof4/CuQVaZe1D/mNbUdACBUbc5zrtNtAKPs1YgZ0hIaRrI0Mo1M6yuCJKNt9X
wzcqUUW3VVOIe8jhmkOpRXOwStiwgDcRlS8IvPmZEmUE85B3CZrikzzGR6erYLyo
jsqDnqZxVco3Jl+TWF+bAw9WdBAC4QKwtcAug3glw3+jvHEe0hoQn1Ie4vqELcL+
wOsdr9YdS31lJtmGJhJCj0LlejABHrDi3S1uUUCBISCEwgPgreGGglnVXvoeV4oB
GG/fiJJHsPqT7YcNDC6/Z3+1KiA/TRcQ34Hr86p3JGaTTXzFUJ2zkLUdbUUwrWg+
qhJZujz9zJ+NKIzGzX0bNphhYzvblxNzPI3Tjdy26iQ6OdM5tcJQmoaB/xFnr3IO
Kq9OWdocsLLbiWg8VEAmHlSlh4zf2dYlmR7n+Gryudlt973sXxAZIQOayl5N/1ZP
gkn6je95NDsgKpCmty1sJ5zHREmwDZwEftZSpkwbatExPEO0PghCPgrxsXBeWS8Z
gUmuzXtVMaRAU9GiL3NdcP/3QOY33SvbPOA2URjVyDVATHAW3o0e7MDYqPeU3S/y
7yW12X27+PPsk4RCfTV6Hv1GucWwk8MEdxHtXZBKa9S4cCTQJCg7kmYfO9Hlc/QQ
WfDljmhe35WrPC1DNmCrNk7G8DO2Fw3EThvgwBkZeizZ32q35630bHHQxDqnjF1d
qQLQuxnOQCHNOzOVgi2c7A==
//pragma protect end_data_block
//pragma protect digest_block
gdygOpTJ1ux73lLlJolP30e1+jE=
//pragma protect end_digest_block
//pragma protect end_protected
