// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
v0uX1eD/MOsuaHwhc4td0i004V3czP4+BT91VEylGlJne61eE74hXJFVhy38Kb+iF1+jIRadQ4id
N3OZTpPh5A/1cAjuUYHsbGuIkLtwqiFYJfqfUTuYZaA7rbRVqgZFGCULeuokqO4BJIhkhX3X+p3y
waQcIzr1SEBrx6auyodSqmhb1cQaRLBTuktIq7b/SHZLHGkQUezjtdve4LhQxZHuEqasIZ63mJg1
FLR20Ut+9NfA2kKrRggOWUANPpnDBMAt/25uhbdOhWNfUpc9jM09y3pJI6vhgkPEaHvUjKTD9d+n
PUHk+jePKH8v6F2jNgbQxctueXGtN9tZIcNNHA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 16896)
GsWzJXotBLSZoJSHmOd8jZNeqW54h9YjhTnGEnqxI9KW9ZLm4IakSVjHj9zjraXWHcM5RAdd52dd
0PGtsJOYle1WJaxFPDtttj1z+Ws1j9RQlkNpyGhxIYsxIDPDCfFdb/1OrDU2Dr31KpyMKtfZxrmB
azoD5wMx7JwLHZ3Wmu+jEXZvJKFkqn7wKyKNP3/vTgP5m/RSagB2cl6+tvBEYFUOL76AC5ec0ajs
Ew6e8P3K/RHxmBjKId16Nj2OXM4xq4Ii7k0areauqagt5CHHGUspyQovzbS4uQF0ZNoDWSYRwoMO
Yu4kFHnr+mH3pnW+f9JEa1XUzeZ42hfmUpA5O1eErURLYWzEiiAaPuTO3eMqLiWy9v4Ls9SoC/Ic
4kAE7fGuiLRkexa8ECQFadVMhZ4nZS/BEQ4XAcB6cAwnpcjBlOizU9OlzjPGIpO7qmA/uvfv5yX4
IcOKCFWUTfgZ0P5WDftBRvuv8UXg/s5sDK0pn3ilPbudelq+nnzvQJv56SOssaGVwWMH35sLNyAO
kM2aTSzZKeypoHBz7ASjyG7/GYw0y197/kEcrpHJYUOkk6S9QLcgisXF5nr4UMKgpD6fTRNQWMIU
dj77crVtRYc7fwVohb8O+vKYONiJeB4BbDFefkA0EkBn6p9++3UajORBUEci+ZD4ZaafQsCKKUoC
OOqTHatU/dfPk6N4AeukvqEqiC5P3FSR4KLUB/fpRaJLhS2oMzTZiwHjCSEgnTyvjaDPfv7T5tP6
thMAEX/KckBZdIFYy7i5cTUHbIzgavLNi+wljlpPD/CTdwbjcqoHu0OUxixGCyUKG8n2kfCj8/wE
blc/j9JYfABiVhDoRLvA45+tBmFfJsdQp6wdtYV78HvyyjZYThrZWr4fJfqrF4/ooy9FWEYX8xEq
B2XFXNjoTRUafgUHGr0ybMHp3JBO/hxXbr2FaFe6Amg7gm2WWxZ4fjoTeukRnGeq4kNNufyJRO0g
uZYYVWHK52k07fpINublCIOf/E0x2FQyL1LPsaMiQnxxrOtR0w5TxRFrsCMeDKdWy3jFsk6MmU3J
ZA8Q8RE0DfEuxw1RRHV8SW2Ef02bClDk/1nK42WC38GKgE2TXVp/dMRxW6HDysSlYRABGNRJg49X
CV7iMV+dNp6ghvsYxS7O2OiO56ekoLdW3x9MfB9jxA7R/JGQZTEdB+2Kvof0EViDVsChtSE3NVlq
jEBCo2wBf3odT6g7QiYSRxT1WoHlImqPItNJDIB9viVu01H3yBaMucCAO5cRt75DdJVJC8fFbuwr
dl1NgIa5mUk97oyigFyxWlTroGbqp68LqcFS/8Hv1lHB2TfuDxp8gMsi9FyVq5baZj5ehJigfOMH
khAo0hUXqCYu1cCOU/w3B/idFbU05oDLptMSEZ8/FtoZA/DRW6UnthN+6+DxNpFI2v/+Guzsah1m
YjUZ0u62cMxXIFKzLB50UiJGCOcZ7a5//wus7GwtCzV37SA/vU2ZNQl+g6hl7gR6F3Fo1wbFUKKj
uFrZUA5YG/5ZS0hi8IGbSJUmzSna9PtSyk3mC4HcI2qz4LIMIAOy/v1XWKl0J8auZLbnm27JtIfn
nYi0+e3ZobmSFXJnp638vvjAPkTURVSR0IUyehW2EEXNrQWhVPep1it+SdJbnJQJtWzVvE277qZH
hVHRtv7JqQjyoKLN8vjy17hwS5WfWAdi2MPEUOe3ghnEJPiyYhhRh4oiSVa9BBnCHewvcdfGqRwr
jt840YOaHXjt14uCrRkRY2mTgxxm2/1vMjoNpTWt/TnJz6dCkpYxRaricPv66KFuNrjDmqtVeuP1
NrET3LmZ8pdtLcFIt3m1/YDj+O7/mtDZvYFbpPnOLCsVwsmGoLx3rbOcfaTVHdEDGKJTTsEsCA35
TX8aYo5tOAMsJHUZd5Xp8FKEyXZdGFWj/Pjp+WpoNem+N3hnzflOAjeHqaxm16bdNs2y4T6Qt0W8
0pPKviKAOcusXXsWJE+uRf97bhBbWyRVfznyJHr0J7o1NcC3S4e7+A9yvDR3AtR0S4NKFZM9wyl/
Ch6I5nHglyLx/uFGaMlfAQABCTt6fjlDf4Wth3efXFkKONZpui2nQdOaqbjzUEKH3T/aeqmO4R3t
cKefJdNWsNiRWEvgkilygw6XjL5j6lPZW4m8HxKIZbk1mgJvaN0utpojJdBGvItCRTcCM99YLVBY
1KAAVlriKnoZEWKF9VBeDWi/JbYiCxqdnEFM1Gj5CHBxP6frhdgiSrw66eno8gMQQFQBzCl1wZCh
9UbtxyJgheS/s6YkXwCn3TEoi6k0oGY3gVt6XIloDvTTA65h7Zq/hRwcFUEFhDcdcvjrBkCRxMPz
1DzuOQfSZpGHwTULY96NwUzXs5KeAzbZOEKPKzb0cP92kgfT3kOy8yFoze0qGH4JtojQhtGXHyKj
lb+mkuMOddGMicjChAp5N/x01MBPikYR6JSqQrwTfQxppZ6iH8+u1+5zw9dpzDkZhIXFXIZ9qiFJ
z5GUj/Omw2oFgsSURvqX3EJG88/NM6mYBBL9xW/7D6ugMO4ulYpy1wZi7dp2TsMjIjpbA50VvG+q
nQAXBGHgXSbsBWH0VvIZHprxIdtwKuCq+bjClhcQFrqgOR0RFmD49A1szDwE3bIXFxlopUL0K7Oq
zUu3WNmwAzkb6VL1vLOPR0M5kzIIXIQfvJUdYWCLJM5UzJCsRKpkWkkmtWEb8WHIaxfL9dnERfC0
52O6tdmk5I3KRnh5da33UGX3NRiwu+FXaMhdVyOPPRY0qfAcsLMHHuZgf8vwi/R+ZJN0XUTFT+FO
Rd24apt3+bp5Mo/ih/9/bXkptkE+2+bz+nBsM5C+x415PsAT9+BxmMzYAUhISPdrRQct1wa3zIBf
V6F+3UIcJ4bBTLIHIdPQ4aEOj5o5I1FtAyk/rZ5CnOgXKdTHn7D3RE5C3+NfF0VeBEFOr/qW0UEP
8q6CBkO5mZuBsJM0SuNn9Co5qBEx64ATA5mjOe2l2nZFAnbpleRKGkWYJHaVNFhZimTRhiG26qwI
RKIIN0Mu8owjXhfc3lp+OUO4ahW1PvJGudzUALcMCh9hxXcjaN9LdZwqj6wlacmJ/mIinJS3ptd6
KKw00Do+JpUfDC66660mu161F9fT31G4c5fKQZzfZK5zpX/6uO9H2PB0PS9WFQDBfw8FDP0qv/sU
4gMiWkkD+Ip/WuzHLh6sA2M37VSSlqGsEGNeDAhIM0SAuRd+qJkVznAl6qDcqnYvAIecwgjdw6Pu
HR+L/SD7fILbcxUBZFJiElldVDjnSdxnj84rzgGtBa+AFAaRoFuewwKxk2KjKz9fza+8/ufdRNX7
8pkbbPiKwCY7BMCu1NKq3RNu+Jj1VpEt40P/rtB0XcVZPcVYdccb2flrxFZxIZtZ1kMFwquPYjd8
QXSrQghOyo9QXQqLgmK9BTSXax7usgqs/CKbhtVsFAi7xbGg50XJqBl27FWdpsd0Q8zWB60O1G4X
RRgW5yoyQnbPIxuxdx33WsGRFFrt5ZehkD6wivxg4Gdb/e943o2aFbla7wJeSFGkcyqoHfIZy5cR
nRdCGCc4H4VH8dVSq3LrQU7YI7hpM54Tfef5rotUePc6BDD06iNWiw4seS4KDEUKHsMqDmCg3Vox
ssRL0WfzSHF2rAxUDD+I1hC6YosAR6SS6NMbHJtkymygjCDy+K/ENhZ9gCMKih9dBdWbiu7xDDIj
sKj1X0oMhpWto0pbpg7Hn/nSWnT8j/oAX1HdnnEdGOtGBpyHnK/95lCRUXvNBgWFLyI+n0w60VUL
eMXHo3w0E2prtATrPUrYsneAi0Z9oprG3Qop9rZCQ3Jqri/iVmuy5vkBR7i3I5ugtaSq1ZHllUA1
B3AdJ/jvxuiJJkbToDP7pDWxR+1Q7v6Fspjgc7oeE5bT6n9zDkwTWKptB76Ygd8n+zEZ9i1MGXQS
tS8mTE46IvKiZtTYx4bIDEj4qC2zAIx5MHf36mHk9gLRb9chYFHDXPUZrBKvSizSfX3lIWEul+Q5
ekfGb06+qD877CIijLfQ+flKXgB+a5CjnLco1I64lBE6w2B6+ILPbQBi8wQYoWWpDm4eSdvg/3rZ
PiZYUS7HuHf0OYKiSCXBRXFhEZzXJ15YuhJ90rZhymLzBQnvMK4TWVDTCdImKkSjJmyrtVw5r/Zj
m7rIKJb44XsFNU7Uqilwd95d2NSeNwawV94KlubKAEirZ6SCM+te2JRRaHMjLsUw4JX83TPbuY86
Gpw8lQlTbQmtRyMd37BiTLwQYa0/thpbc0LvttBTWkK1Zsk+CDTYTC22wSXGOqmkR12jc59QrUAr
2owEXdpaloHvn68pEaHm+Ro074P91XtSK5rFAhfkvz/VffLYHN2vzPYno/UVwW8ixMI8Uuly3kvt
2D8Mz5zRnABAdHklYPQrR/vZHLNwMUDvE8B2L+3Lq4DnECSYy++T0h9IYNJt+dTu1vSONY4FmJbT
/Z/UbMNC0EXNt0+9i7zykCNCMWDPu1kQb9kxifFVyVDXiOucxcoReKHmng8ko7kIFGqY6FJDnRwL
SZXMlc8QdrV0iTTnOWTDNHsNDQMMzO92PvjM0/awvxmVraexgnZTrkhnS4F1TCHa0Z1S3ByJvA16
ZckBGb0Gb/cnbw/be7TQujxg0duWdAA2FktD6zACSizMpDIPUPyNo2+NUBohSZc6ceH3OvZtGHi9
cp8vPFVq1s5m4G/sRRt3LhO7PYWC+xiD+ZOBn3Lqd3e3S0uFp0f3dIUNmHjdLLJYRCQobtGMX81g
+tZyDKUn4h9VVtXFzc715OQ/Jlsp6PaaFBuAUY2/fVvgdPVnw+XucFl0Sx6Oc2LJnLg+QzwDk58S
TBOuV4HpWMhcOejRKPd/OW8o+heedItnyDFf4us9L15OPH4yNxEPSDN+kuk2xm1ADzINGpioJ3Pz
XXjBzEQQQeayO/Tx4+aoqTq1YLtLNDjWEyAj1dsaTmvyaUDBJIA4igIAFYNJ7eYxGwPHzRfYTz1E
oKKqKNzBTW8PNQcOikHBfUHKjDYcY6JSsaBtHHRdO4TdDu0kw22cYrNiHZK7E2N01TJZvQ0yQj5f
zu5GJ7hbsTZRfxxymZwRmDYlBRn6QRrREQZHzDMcyipA3k+5qMjxpLMFkL0OkVN6jeG7fdw6BzZH
wNlU3zvTdcz2wIWMKPvPSosWf0A/JMN+uhJvjZKnNSYckX+NGrH4OJ9IGEvfwcMtqKU+cQ8aHlRz
qOw618vXb8UXZWrP2bdYO3UN/T71PX/ILGVE3chxWCYFaXifcPqT9OrmA21UjmIHNUgtgONJfFbl
Jk1J+oHa+n5A1tHEbTFve+MV5WyMAZ29FT+sjUT2zml6Rg/R5BRVRApjyUqIohEKhH0IYvDYHmlU
MiHf/IQrJDqGbamxYIEgwiXQ3S0YV7rs6iH7D8XRoOTX+MY5xjN8iVX7sTEk6v4976CqT284tdZS
gBQDYbidrBDlawFoQniiZ85rsH91eXrtE/I8F0Q8OuGRrjMkMCbrEpA7AggKFuVMGTGzR5m5CWYc
mdxbMfocxp1XYeT4iGvqBmwL28PL3ZfuiYaDoXOXdHMMcZg6bBGWIAukqPBSo9dhDRGO5y6Sbc6F
ZWS/FqpYx3YjXHwnZnpO21CunJxyFqmVs1CZ8wS8/4hBJ8q0OjXUQhqVwIAxWmHAtPd3vSdUoi37
2Htfr7s0Us/ne3wuQ7CC4XSYSW/1ymQw7TXPuZ9GHXzMjUkFDlCNYZoFwuvKqjza6A/4u2xs3I/k
5o76iaJ5YoE5rBXDkbrXiVV+LsN5iwIcAS+Lb2EdcqWv3HMuewTX7VgZFmr5mqeppC9LV+eOGNgH
03p79IS1BY2ZxvIg7ifdq0n0pJzcpUR8J2a69EUZGDm0fyz+d731mAOHbpuVu6G+JX3Vm55jWb2+
vXJInKn1KDfCFcviI3qMuU7fObmr9Mly/+0mBYAInn8JDHe73NG925TBrqLT8X7oxFtGFAXWVNHI
C/C/7saKC0r3Z624pDCvm9tSlaa6VFmsMct/wg/vAZD4Rz7Y0DZdIoWJqgREw57UplSDP2NK4uzZ
yRgB5RpWlq+fXytCvyCERuF+lvq035137xhKOwRF0luNWsdg2zQ0YDzVxGtHp9qoufrUOC5cZxPl
GxZDQUNVvKgT/AU4E6FD182v7cF3AWwI6/5njmROEF36kfwHnW4GpRlVXjG+uHuJtQEnIJYqNBpC
dRybiA/wpwicdl0ZYpQ5sb119c+DpMnjcQizeJxQ4hAhMOWhKynRZz8zDZIPvbpVM5vxvnkNY4UV
BMdUSp7nhtWqiDee91fXxQ0oTGsBfF4a6eSRjUdxemQ7fSySc7QaM4TRWN8F6E1ZIdYSmvcBnwr9
7J3a/OMqW5XUV0l3n7dIBIWH3aYD82hbzGxbP/MMr1Z74iaruLLDm3tk00G8ylXxFJ/O1MzOPFSu
0AXkQ31xeC6Wd7tpdRMCp6u95Pt2hed4h4taN6C1COxwhcgVj8c5VMlW8OyLe6s1ID7Chi8EHxEo
l9+ybmTx/uAAZ5+Jw8Bf1MGF4MvpagLTBQoZJWH0+cX/YZfKkuinO+AbmK+/eh8CwL+S9TkDv9Dd
bVif/g4wspYVQexQZgjZjCmUe2EA42An+iEpGmjkNa5sTIs2lvIj6ZHH2yaP81gJOKj/5vs/Qf6b
A8+bYr1mk057zp8/Nu+mkYwyd2A3CGFHT87GFbWmfHOTgMeVlGeAIPVjI5y9ZHRJXQQs09ahd1ZK
l6Oc7nhGhrsgfPZ0D4DYWKXtir8M17o/SpITKDVem3J2dYvp8/Y1xadOJmQThnrq66J6IYfQNzPK
BAqfwDB6EZ0Ymdlp7tTItSiGjXoZTfuP9oPt3IkYiuce9pLt80FdXke9w0Yu5y1N6WkdEzmJBJ1Z
0/e+3AxO+q/YF3vG4Qa+F8oioasRv/DJIkwWEQBAIF9hca3YpyXaHixkfsuHgm1ne/miMP8bfNxB
ceDYkv4Zz85kJhrIAjvrqORvLd1idd/kJXwSt3PXdgT6OobjDi2RZNP6lMWlAQtt06m/ETUbAzVL
XJN5ke/5GUJ5VdMrXVLOqnJjGCFahOHC5L1F9/ZG2DVqMqd3WBFEzSklznkIqni21IeOdWsuoeb/
0KbzBVefnSyS2XzDnVBJ2jYTGOIJgdrKmOA+yseNvclP6+1VJlj96E7QodOF7jvANQ9RSa3zHn3g
cmMq+8+zCpSR8FwTMSEs/23vM0vxhTBPFiPa8QqoqeMp3wJaXgdXKKqccNH3HHGsp9ZT3G1QVYnc
zFprnR5c9TejHq1x9nRZrMhM7TMQ3YLweHEE2FRzur/aY+8BHqruNec8ywvSDZHaAlduDFnsAIkw
ctkKFunEC2aeOnjO8HnYkMop/YOWpkTVrClAyNXvFtriixISX8n+X/6PCrGZAcq6wUFu4x2wiqSd
+SL1BICqJFBEagqsPdOFiq7d4R1OqlgSuYpgbS7HSPpHV/qqhZdbvbbya9IH5Rco5gJXQtiBZJG3
C8L5tSX+AYmyyQuTf4jMA30gwViZPNu6gwkZocKpgvCebGto74MU263ACyT/+TeV1iz07PZ+Da+F
zOKJaSrjwOQ6itoOrPHXHnRVTcd2tcmXaxYXiASLfmvRwpF8/LFscnNVntCwmyNiIKFFqFfW9CYW
v4K2Rvo6Q4ehKNMQaQe67k4XB3ucOvGLk5G4GRcE0DbJJ+brYDO09vY/eF50eDL0CuNekxk+rTYu
/pCSIhbSjwTU2CDcYD6KebeOk35A8Llfy6qfrH3yYG9Texalk1Y8QwQLnx3XNXGBbK63zgDHo4W/
fI2jqBTwuqNLl1cIk5dSVXiIQEOg/CZ0wY+wzs1+Hg2JB7qYkMf6V4qWPNXnJHZqd+AUHXSYB1qT
/bbUdNupDXYHy1WXSslNzW7IODWJozXXsr3MFOvjIqb2lxgQkoFKoSCB63YsY3ji+ymg/yUTXAaT
5ijCI2LX8UJ86t6oSSmpC9H4mDde6V+J7OMuV0AWCdmnT254QLFMdYykbmK1uomRMTiGACos82Mm
6zkfpeEaso0s0Kw9msLX8/wLeq8F8qS7SDPzi8jDJqcKhhWiDW6lduOMLxnaTWyNN0Yz8x1x0zUi
6a44wds0thbv4GjFPdNoPJjc34KX4lUsMjWkUuUAkEczf2higwQtonTliJ5u0PxFR3iFftk6tQs2
LvqBjM2i4FEilOpEfroCNUPX+FNMaZlY8lm5wv0UIP/2R1LFZ2mDSeoqR62DmANCXaN6zhqgz9fT
a0gqO4dO7eDNQ+YNWqSgj0qO8xIzr9RsAX5gzcl6dWu5sgPQ7pvbV72mu8Bv0tr0/YHytcjjtV3z
EmM3JmhvZ+3V9UJTZymJy5aipaV+8cabtrnxTArGcGfeP4v5PAsetbbgsqOm0woXq/0NOn1rQCSZ
QSHBBm1aYFH9eu1g5pxcpSQnuJ3BCBnaYoCUvkH5T79Z77OapZsqm1SKtVbfM8aaghUkqdIZ6GUM
4e3nNK7kvDlf81K0Lm31lKs9JSRvKakqkD9WIrjVyVyz3eEJO3DIr9gWfHgDRyqLtawXNGkJD0j2
OQuF1A46uw+ZPT2twjYDiPzhTUvmMgNobmmvuDiAQHdJZL0voXhQPmJ5CxGoxUOTlXiCoe56/5Gc
M37AWyMFlqRywZZJMKbaGrAPfWboVh+uW7nxqSvtSVFJjte4iyD+niLQkT48CYleKURRah71bVs+
+HsD4VucUWgRAnsbNRrmcJaOEhc3neXy+Izhav1rYwYvF2yCdi3NvnW/s2B9YDdY7fZ3kXl86cFd
DIIUxilaC06xyJGEt6p2YuvbMCuEzNu/AbGneU3OlwFvEmjpJzmyPPHJyQX6naonzxE8pk5DiV1J
fP7RoQE+2FZGkyGiJ+YjcnoGlRLlF6j49rO+UDrih337Ke9WqpscA88QAiVLXcK7TGBJp1EoiVwJ
3IUcvpYZwJWm49acRUutyPsib+dQJcz0chIJjka8NwC2gyHuMfHTz52+Za0/44X8ApAph2db1wQ0
NGyoGCe2C2HZPrzynBpQcxmwAxHrjiOy+fQH6dS3r/l9gquQLzCHyTDXSJg1p5+o6rCARD2I5nVY
zIamUg1h+lVPKM4TvOyCK6IgxlujLYJDGaboF5GJD/3z/rCNikm9Iy7dQBbBDd5HJYsH6foI/Lbp
qsGNXoJh7ui/Bn88hOxN7VZ45lN2SjLp0IabvorI0GYtEU3LVCIxQJSIErLEL/DJzHl9CNWxX1ZT
lsEeUgM6hhqrTDhqimfyF5QLPM/6QN2/X3Erxkbw75oRasetyQAIr57tbPY5kw5NhfIZwrfJj7b0
CSphus6QxdSPhSmZjKodyWLwM7qzzVLx+52+73Oxa9wExbjKvVxOCZF+D7Cj4IMjGfaw+znqxFoa
Msg710Qjq5589YTWXyePxo9k9oqhQF6V1HRcffpr/tiBlhHKb6NAVieiydS8r6yFHTg/F4KcKpSO
3ZL4nlO3JOI8dWYLytamJJcIjATbwVYq/SgZTHafqZM5GAgxzWu51CfgMdeyxc4pLkmoJjAqcF/8
fIAAYbw1PhSffI1Cd/SURM7ZBNmO1kaQv6iCucwELF3Xg1XVm69taktaJDpxVMJbemu5/rhjYnoR
cSJgI4JcblAkFqXWw31xJqoqRJYq4XJjdVqhvPbicRYrzDURHx2kguW58Br8f45hPAEUEaVEZfwv
hKzQvp3iRnkw23FZqO+mS7dQioxZKFbCEGGXPu1AJ/qUa3wLTkbLEWHwcigADeAgBp60wPZ/rVnG
YaJN5fFAnK6NPSQoxsdCPFFiFb/OeY3ll4iCRVl79JgVvws32MHZqfj2wCrnmZGOiEgYq+i5k/ug
wfaSREepnOq3L4q1O1FlxnvlRt7Q469nH4+que26RB5tys2hggmQwU+yiiQy0bkPNMex2uGPnWXQ
U8JmOLakTg7ZVKzqQnquy2zadICvVMzDXV++iQePtAGj6rdE/MFrwYVPyyHxWRvap2tSbUSQcPrq
fuouv6tOahAqUztiBgfhHc8qqq7ULd6OToCMIs0FnZzZZ/ZsBs8vrZdAEufnGughK5U5GkdK6i9Y
CgifTwBmIuio94+kdAoEQBShCDG9Po0ceCpuC7vur38FpGb74TB30g8pKD3dOof0lixk2DWTEIZb
a/e+10BhJ16dbgrhMmxlCuq6DpfR8Zd2fiRYkLm5eN7uFbweF0R1Jlu3KrJM4isLilR5+BaTEpPp
KQpwOxtcJZrN3ng4PoVlzzAa5dU+pyRddd1f8c1okMcMHRThSErGJSnu8chyk73yMIWNrQO5Xezl
lGDN7wxxvezmjoCFnAyPrJI3CXOH+sukTlKXKhH5XqVXtmHGrrN4oHiHV7EC16YEwMCs59dwCILl
eU/RcDUjUsCwpLoqoRR2Lk/962Y/yx2usMHaFPEiQshyeer+TgovhFwU3LiReWqs+JGBrDsnKol9
NcSxTWSH7R0OgqtpxYfGTgEldTewVZBQfsrY0ceBStqRRK95Dxp2Aj/IN1ns7dCMI4/5yndavkO/
9q0aeW8v9jbrDyQf44WJd8t0ZUXdQqLDOXXiXbvX13w/r4Bx3V2xKw1D5mMs+MgK+xpuX0BYL4xk
4cEIWfj2ObzTCF8VTU9rPJUquyl5r9feZ6BYy6STkmkPTWZ87cjUvvJ94qXiMsA75JdP555zGOmv
s0mcibdfMUKXRnvqFgdFAKs6ODkA9UJj6ro9DfabxQlCyg08dcCMbxdu93b3PZWtbx15eGOUSr+/
2WGlr9jnJ+KU3tkXnFLbHBDYJ/6vbPQ8djDn2c9RHv/ZSth9btFHwZTS2azhVtMjpJjiFNkWVNKj
EJ/Q262+mMeIqmif9Y8w8GbIhU89NtJEC/Ngx571/7MJN4QG0uWD8VtUxhq4xyuIKjsrC5Y79J5O
TmR4ROFjLPnlh0HI9sPN8krCeQIkY5KlL2wI88ovB5dStB61kmvBe5K6GMw9uqqX/gs+kiDgG5AP
h+CyZR3RNTe91NbMe/uS+4inxCigN4idKMnRTpmYK1WpyAVyqdbkMRzlOrZUKgqdCT4DW5+TkmLP
oTLq8THzIJlokREN2bodh8oo0w0WtJsBwaKTgNlXxj7p8nnAtSrzMyGLFrx7o5216nu+j4pEnOmX
V4SQV5Rj691NLTChL9ehrJv4A16zV7SE11ZsQO//Cr2C+BVv2HYnyCj+vp234BRUpnAtUT2YF5Te
NFEgyl3vvMmnTU4fvBHRAb5EiLt2/5F6ArL+3mhiXkouLxBY6mexzUgKiyjczuXvYVwbQ66YM1Fd
UJWUEOwwCeiYSeBbtnMSs6JPMquLsAjMAJsjtOrUa64GNPiOvhdf9owYZjIdDOH9fvm7wHsvEDci
MNYMCW06+SQVtajGCOioVrjZfm7kyPbauZ3LnLPaX7Q1EQfftFDRLGNz8wckACdCoT6k0CyFSgpP
CMmEndwQkH9Ourb41uQsroGtx8aK1HYtuYcA3kwREvwMdQHQ2MQki9CdTOewv6W75RldhmAXcReH
P2NIh8ujConYbT4aB21h45RXUHvcdqBEs0Cub5XtQjMA3wh9KYCUsMVYkhnEG3StJ3qQAnS5JTti
dSWDDkLVKO1ub7zBzDMY5ekYtXQ4dp7HqSjNoPtsL3Q1OqaM8XEAkqIP5GUHsIsytX6W9/iUPiML
aESFJKH5DPbOv+86JmthUK4jMTp1+v+RXPVySz6viLMneXLuuwdpZQts8iVj4Wk1WmCoP9eptkot
2hkef7vpbJKRhhlno7lprS2EZ5NaDsU7QEev9gkpAy9zY1Iso9z4nuBtLkEt3RejPyHej86OKF/o
HsW5HhLvUlvvDfVgxp3dag8TP7fqMEh673P7fTTgDFa7sQ/XAW1bO5hbl6JtBmdq8VfUmv8+gELR
Sy2FVQHHYL5q8qmKSCdjTyGKfYfyU5+GgQwU/y4jc89aQm37hzq2GYo9/64K5/HwrvC9MdiULXJo
bAQk7dSbQRUtW0C3Yjmq5ddwFrOCtrJdhuwwvlDbDw3krXSMLNCgFeX2odsZ/XO0iBB+xagraZpE
qog9dnQqzok7yu5G3OfFzP4im+a8xN0/SIdGI4toSIjIxSeVf8oklXnKlsILtiE35iUtrmLNmaCg
PCMoCir/UQPIfGRREWG8qG7Bq9ITcfVJemS7PQW0rVCwz/e/Gcn9dh73gDStakj57eJEDtJSA2Hw
VjB5H+HRJj0qtezQu7DuGMttwwLAwTFpEW+M/CcRc2K5NfPPR2SHmk7RftpvyHTuSjlD7ndRxIyu
5OuQvSb+LjrmG/1vwS2yAvF0yhfaJk7DsfXl4cO3mKKxMCB8//mzgXHZg/x98OlbLjsP2mfKsNgO
5ZZNeVuJNo4lNO7whgdhgfrjm3v2qNs+MgCljGEb3bGHr2yPtrl3G9YSXY397M3L0ZnZZ8ZAy6i9
qlYEPP4LqyeY8pDLmBKONkMYhoX5MeydlGyd0qBcdCnOtyJGzfczmJpeASH9dTNIYEjZe9iGPFJd
Dgyc6i6X7vcbOiV8NqXVRm7qHho8psAjRiFh/OVOEqAbiADlkvvwI0uZu83fRpJeFwRt6PsdhhTZ
O+R67X/BbYJVB0zqtYJRypgOpDhVc7I7kkIOMVb5o7x0BdAX/Okfu+MpKfWrpZ9/f8BaFL2FKt3k
w4Y6DSCfVbvdSiq/IMnsiFcC1ac49s4ebNYcRU0WkATID+evND+oGvR2wWtIvoTPe5XrJRpS0RQW
7kEduYejKw5G/fYj74uBIZNL1GC5jJohbFn4Zqm1s6S4ztXZkGf5x3f0yE9IttjJoT1kwsmS7CRd
Gk5AC9Ade2toagZzJrlGr4xthrBwP2Mw6SWW41jNc9L+eZivSB3gLN2+hz2no6CyEQ7rAdIqaaff
K1BMVzWzrtKiY04pKcFbIbkw3qwdGXq6K2nrfKku6M4Ug88NzEEmUIKsppoCtj0Zy0mOATQ/4EfS
HWB+92SzRx7W6L6CgBLODxx2ZHvotSK5ubQ/oqBTjHQqije79bgAQ9S8YFxaJAr9MdPZdaJlOlfX
Fuj54ZtfFrItlDWa2wSmbclUFHGKc/gVrGq6yBSSuok7NN4QjRMyDclaU+UAaLvPkMjYghE/5pCP
PmsX9F6OKbFgtdF4ViAo8TzkqFO2kzBmbx62/yuVY4sGngA2FIQrb9wOsEP+sF+PfRJ6pPVMxC8d
p2ZtnUuIljFWW6PEJsSCs3MmCwWuTkwXsctaRq/4qFwmtiuqWHfBCidLRb0FcthRGoo9LuMFLBJR
ZO/3XinSJPbRwZR5dczNmCkYa9Aphzn/mxpIWYs7pgAYmgjaCfPl2VZznSd8ULERJsrC18iwoixG
3FxbZyUiY4hw2AP7aV5BjKXrRpLVhGyGtTVs3WIMWGlooLZ+ti+WAyopVeqjq9HNPhtT9+AeHG7d
579kOcAW08np3t/qiCDKyrHq/pkQD8mM2ypuiFOYEXvYMJeowQefd199wL2H1uRL70DvPBu51hGZ
Ggum9IEKJmBflfdpogAsGEqMNuFZ+hHqcg+VfvBnFnuMBAi3QI/59cMf8S1SUzVXGS7kcElZqRPX
lq8mcbPiebUEn7lBXztDTXeM7vut8Z9k4wi8nIwU5FjJuwqscj3z9iZ6JC6ierMAetiGArWYCRyr
Pr8iduQuOTJsCnzQiEhJop5QkvmJu5K1wUEuS9msrAfh3srv50M6ij13qB7vpYPBzf9pkvPbZn6+
gf/ndrGAM00wupd8GyYD1aE3QQv21y9PXXBh3DD1knJWX9tXCmMY1Y5y90iFGXlMb4R8/ar/FB8f
kkf9n7d4ydjYYKXSF3xwWwjtQkfpsKvfBxU3p8lNiG2ahTWCsgrtJhyeH32WP8JWNY0aTlszZfef
JHJ3K+pUORigtYCPTKYTZzJBRC7e/nahE3wVW65TgnuzxMA2oBdczb3SIxHjL5leoang4Si9kVcx
IY5pI6EKZXw5WPX8B6CnERIpXX6N0wphg2FUX1JmQYbROKFbntJjX6PiauRepU5TPcUBliju+CsL
Vh+5QJWLHfBrT2OMKoUppjTezTEELUavsYMZu8waj+U0s8XoFq+/vFmBwoEyGkhjtA8ErXcG7ATO
KJNCLQyThYO+GiEEi/1Vj0Rb00389FDyHSLHG1x3sYG7PaxCwfyiTE3s61QJWWRA0kTt6JJngmPG
UIKNfPhyu7stKldUWdH9M3B0DZTR8+gNRVqTD62b41qvqcd+qfqKs8x2vpqn1A+yUJTjHodB+i9y
nDzh8pDjP5ipnnfyqYouQFHS/Vg8uFTRM6TGK1gXUYij2ZGu64vuTBxWCiPHEPWQIOUuJdpjljkZ
hPtO0w+Da5X4yIWk4HKGgRkUlbM0yinuXBkTYYBSI1+O7Wh/52ENLbEQrEJYXIfjd1zDIiS/VtfU
HExv0NG6E/WfYJ7SjkJ4XxX9RdLTYrvjJ8vGbnutSW+Xxx+L4WgjjXBcPGlVEwgRiO/azgiEBK4T
0ia5m7jx0hh1KVZWguD8KlxoFNmBj2TtiayDtU0VVHIPyQAXAY9ojJzeU8Xs+6FhVId0yJj8kpxa
/eBEIYupcfLjoQYsWGLVnpDut9+RHNQ+K0WtfnWRqr+2qCQl+BwQZ8kVW3+2Kxu7TvdrUawczshd
LhqgwaT5khcY/m8kB1RYX1+EpVc9YEMvBiQUH0yFey9/gLL1x9W4FW+G0YN+X+6Ex1uUvebboTp+
38T2dCy68SrnuQ52+3nyHLTJX8yMKT1MrnnBv92kqwvnI/V/oMLCcpdGQqygifvKoGU9kFG4Bniq
0luaCUcvV2Y+4KnPiCXHJZzp2Hfn1NaWFHRkU2Gxnv7SwNxad3B6GTt1Ho9KdawABo23l2IEpwN2
X1lARzQae0N42lnIasNxlYY5JbhT0/U8DbrWL/P+n0Zyi5jRJ3j/yLSnPHIOdk2AYAW9gPZpPrrT
gyeyjKln83deJLeSLjdyXqWxh9qgJzojEdJXD2DGzt/gJHquOGb3wUMXnLmiswCHa0PYH05hkB7/
Nae8RMrEn6KK9zmTtPqCqQgwkQpu3rJQ5y0xpQSpnO4CzHyC2T7/HhvkHXLmEo2tc7cb3yyWl/eC
GxoOUC4TXWyI6aPm9py69qdydRvRVhkgR7DwpMCAVnh6fHnJH7lEe5aukWt1+0jxJELG5NWaeka5
caxt3VcpGX6rcLIl4czVe0oxaAolBYKLStBWzhRtNvYUZYXbrpe4376uGzcELD/YanlWgAOM2SGj
YVV+jaHlPd2F2d+mGCsFZqVZ8nwU/PoAWQmQ4qOc34eksFShXwSVR8xMp2UTtVSWaefqyo81L4v6
7mukp8GMaOF+nX9nvwi4pIS/E9xT9AzkoTu7FVgOYmErnYGQQ1hSgDKrX1ltwnbQ6kBMIl+HUkwG
M55l+kNQ4ycaUThMsqeQD7MQ+7p6ga72pvd+LpePUA1Aa5t7cdVSaWViE4gkWWHXAyrpO794OdaQ
Vkq+2D2Vz4SiAgazPpj/4gPeuhO80uQlJfr1ziEL6JDXbro8x9ZbP2SrqxmKfuwF4gjnWCEtRNsS
0dQYlPRZCtm7Y+78ib4xFOIo8hJaX4hLB4Qnq9Biq76XyusoN1OuVJQdFFU+CwJ1l7qXtC2iJUIi
wJmUQS8qXUOgaA4626xaigQ8gIMFE4vuBuVvQ5YdL7AKNmaBDZlB3dCVFqKBtX/PxTgqV3fP6mDR
YhsWvPTdKoiBym2iR7/U+c8CDZm7QYNk1Ex9H+LSHKQH4A/sr5qMvmQF+Q8UMdvCy5Y77iXmY95w
atYs0/xCWdA2YOEIsTzzmMuJ8SPteWb18pI15mLh8fsdlbowKfI6TsguhGPd/hCsPzRTpFo5eSSS
ATCkGWxgUMJDAt564ArpHNiqBPH1IxegsuK9L2O40j1ZJSTFCrg6Fxg5OUDwPio3EF8+yMMk4K0Q
xYBxRUzXEfbG2FkxYJVTiI0FKe9pgwOkdTx0ZlNfYnRm3mZp5lMnvpTwk1ipNeEo4MKBTjTrqqCS
fi8bZxLZmjoWiz0QWI1IAALLrrU+TdZ3H+A5m9FPsi/J++b/N5JOP66sgjR5G+GV1ixcVAdcJ1Fa
HzAcwx+3GhV26qsJVtrL7XN0WglHT/QGH6xUEymE9wTfcgESh5XWB5OzbHJ/rZEiPoesF2uKGcNy
Ykgf5ncig30Fx1s2R906+yxrZ9wFDmPQcrbCTv04DggPAd9b654BDimac/OI3TgPrrONrtkvHQ0C
cQf0yvyABHtFlqmOQXfkgBu5ULXFfUSOkEE/GsDLM3RkFzp7laQUp+egEEwSglbEvLKl0miA3G27
JH540lyQG3Y4VOTwQk/GuHr2kD9p056Gpu/5Oku86NtuGxTgJOjHa9RSagQdiEi3AYdu6xGhN1Hi
Oe3HDdDDyG1+NiDTtjP/5sC+Pt80BIINklrPk3BkwjDOliznsC9vnr4Qzz6oehvGQbePKB69DUb+
BTvMnyt1WSmXk+4AfX5kKTcKrc5NbkAso+1OsG00kX9Pj9BekiRCD9C+HRttrdMxWG/s331FOjyw
3MkxCyoiDJS5OYIY9ns3u0NKBW+w+R4e1ZhZEvcdF+1/+a9ZiuC250+cs39BldJIcK0pJOuSIfDI
dHjeiVOiBqKyJE2jur9WPTwv69LmQsBxzb9rCNrncefNTPSu/G4MzWVLyCMzIxOFBE2bVIoi5pgU
zOrkKKQW7zCbIdpaEHXT1RaNm3RvYn+GR1VLiuBOc/VBfmnFew200FomcOrvLSqlCb2cNM8MMB7j
QPIIJ72uXV7x8urKYyvSbuPJy9eadP8ftiatx/5dgsb3RdVrGObq87rfb0RH+OQF0AJYHm3cgDal
Lj1SQ2nT6nYifGeOQKb2mZIKBeXJay3ZD8ehO9BgBRsmeROmQgvHva/LdBK8H1AIGGT5/+EnVWtS
6QTvDNb0Dsno9eqBdzkcMNiZiXgD1FaJjFATNDOzgc5LGWupMc1LLkSfAu5jy06isMjxuRMrKjFb
NJ9LNenEavNpwtEy6M87n3KpfNBWGwESYaeK/gfR//98Xc9XB7hNcEHsq7SKhAHoNt6flKjNQBd0
ZjrZJ+fkenjmhp3i1ptDBSBWWQmx4Pzbx1EZ22cbBVeEb6YOuaSnQglYocu2LJuf6rZNuvgvwGY7
x/GvIZHZgerGBdYaUNGIkBgOkTm0hfIeqXDee12RMB8hNhGwzyppC2LPWoKKrfsf9oIHeTmf2/F1
pBq7EMlO3oJbYYa/OuW7/8DqqDHIWj/v98yxc5eb19GPsnNtT2MpVMffdoQBmvxdjNw19Fb439ba
nBDSsSmmt0Uni3BYlNnEbSqNJkDQKujlgKCjqYYJGRv3HvQOXkCB95/xiE1KUakMWNe4Je5ZLOke
xGYfvgi7NwEnB8UOX7/luPdhq+SNzSQStybeM6TTn8BRM2UJyHi4A2QZBhFCrYQIQp0j+YKKnJll
O4u1GEzTwmtp1Gc3q2XQhBlA/iiLBD74Vd1a796IpLPM3h0ZfoHNBOa0l9XjyL9xofiFiq4Axjjo
PtFyE+HLk+Eq8TEv/58JuteV1oqFZiNgK0jOBdb0dIx/pJedRFj0GE+/UzveNdtjMJgt5ciw6FkU
/zWpwU7X34uC+BzVCBawysN/a4mvm9Sv2v1hptCM13wwoUqqT4tGCky0Fb4gfFxDfnH4L37C2LcS
koIRNjeWgEll7TkE7S+xepC+c4hSpGW+zy+bA73TFLXnSEdBlrp4QrAh7mgbcqnvCDwe2m9Ed5rS
bEdr1pUjjwE7M6U2M32fFuz+XEJMCAU6TNG7uix1ifF/S+HZTGvbN8vnQsr1AMcOk1UedXgZ9Id3
r4Xjdf7QUGms4kQLLptkbeX7ZFWWVnq1+xQMVPABeEbqLJUvOON4Lm9+zj0OBIiShLNpvF2OBkhi
4gWLSV2MUttVclg1Rbxj0izH+1z/A/TdIDhQtS0tLS+2k31ciuQElEA6ILYTZvJqXVmQOC7Vhb5x
3PI2Xj7yXbd3RuM2UXheZ6e0hrRWZmHT+JoajHee42Ihtb1mLQuBdq7F/E7HAs9APUSig9okqPAA
snRhrxc7y10LY41iEvALLgr3YSzGBC7hxpi4xqoCAWOqpIBpDzFnpjolZqq6OWexR1hY8wtEO/hq
OITmaFOk1emB0eHniZxefbEeS+U1xOurG6SHk1OForIlFHzeGVch98h7wA5nbtgsmw+j+MxCRFDZ
gdeiZohl6po5WpczS90tD/0y5+MHrDN77xwQ1Qx951BBTtTcMkRXmzjol7en+O7qXmDPdIvlGa0Y
VxjxEF1TZNx7HN5LTLdtqr08x/WBLiPgtXh/hX0kor0PBjmRDeEbPYH4KYLNvQniRjRxZ5KcQ+d1
O/kfcnvYRQS934PR7gZNrNA9sfG6p4Exw9ZpFBKg6ho1Lb1aVux21bub9UGN0JmgbolzeQHoh4uK
Kxg/OjOBO5cFBY5JBBZdc8fut2efx54s0+6uC6b5d6ghnBdEKVzJDBEtm9Q37Z+OccEKUL+F3Se2
AdrMy5Wa80FKqwMg3MgAsUnKj/xbjS3fT3EQ0/npNga1HoA5L9KNQx66FRKjvUoyImzN9Yp9FKGR
RLQmp+x+4W/EKYaIa83T4uzb2W296qz40w9HAD4DmqdgVpiPi7es6sxAS8BNYQMb7fwXbZIh06iN
lsPW3qtCBewxTm2aVYCVKe0e4Azi9AVH5Wu4p2aQw+OS/Mcsr0WTrrjPn0tXEY1+L2Z50aWDzfnG
hXa0+XuFDsL/+Jz1FakhxXz7sHha2IeQUCu4qxPo9MwhPRk6Hu9MUx8Y+OZtB1ivYRe8B5ZhTAzv
44FPj8No+U04UqJ6PwDS3UZR35fqZBZn/a8QAsJsndGoQ+yqvP0EJO28GMlPMHpxC3MZXS3zfSqP
Lvs+JksOYZu9f67PAVwUe60yQzjtNh3RhHr4FiB1KEqp+3hjGO4Q8xsVrDwL1sq1HaqN7vxrjwIx
Rc+XFOI/6v5SAoOb3CTXgJuNZx9W/d00h9LQ5ISet5I5Im4Ta8pUguqDW3t++SIxuy5xIZ+OyMPW
HEWi1Nj37BSF1RZ33gkiu0Tm0lCeKVOZFMamY3fzt2wTrWJgR29EOOfODV85S1ThoO4nBCJJPyvD
ppuczol4zTjwOHGmgbBTI4UxCDKkJ9CG5bJtYIMXFBepXyaZ3WhTvNy4fbbyl7TQ5+s5CihTvlJT
gRvw+HlmmfMtXIpca3dAvMWYjv1JQhPdLKudmtTwpxAFHyHzmNDgGCCJDKocF88SSa1inUrseQnw
Db6XGSBJBGFBW59E/55VXLzdsTsJnS1TVfxWbgrIN8uv64KY658N9mH6te9ii99edL07c4QA79iM
59JBO+htJ/vTIyQDY9foytN9pc2wPCYey9pOgVf7CUGNd6fyN7M7XB95b5sQhcjJQOdPBmsYFzqi
m7OkL7wjnZG0tuAfYT5gHm3DqvsooJbqV74PUrFlBswWA3r2pYilB1m0bWjDr4NFG1592Hq7R36W
/wyvfQ8NuaDbiOxCnidtnIrvhox8ENbErNqDKYCLxqt+h38cXW4gOcglC7l+ue9PdYRZLEvOt7nb
I9iF5YQ407UqJFYDSBPakujfFSwMBAfYty9dx8cHbOBcDAwAcrl3Yu1hZi3TKj6BPxVMgzHjqxZG
3Ia8EiKeitMEn5kXCUMJDPO40jqmtxovsunN4p9I2ABxXNki+US03V36so/P9X3WLv/byi4n9RrY
KbSo0E3DO7+aakVi7eyVVBK1hpcmWt7ocPEyusjuhRrisiGQ/hRgG1C7CDqN7bH9U6b1VZUvEQDq
xgeNCXoouGLR81kaRtUSnY7MSFwpz7nG9dvfCKylU7sNgFOuuW4XGE5Cgt7OPlTD731zhQXNTZiO
1LoruMnwLrYN0q6gaQoMvXvw5PBd6JSHa2EycegNDB2taDiSYYQ2R27jnk1MjY/dXCplk3DDxiC0
o89J7lHHEDNZkKug0eTXeovvUvjFTPPlLM92BpbityxuOvneYGRv9i3LGIeu3DHCe6DyFF29P5wO
YSWATudBu12e3X/V7O/v0paCdVahbS9UFlmZfArtNkq6UiISCHXl8dZcs6XP1N2nQsF+3NifklCc
XoiJ2GYLiZ0YxAhLSMTSiUQYVFUEHU47nN7j+NDiS7nwYteE+5fF1l6vbmw4nWQ05nsis54MTIqC
CO2Ibv+c5n6p1870HdSg/oKH3d9WKptY6agQYEOpNPEcAUo1gmg1Hi0hRqVoNefwuy8EKnZ78mu7
IyO+sEtshjysrW8tap2nwm7Hk5nk+MJlY6Lt2d5LnAP7WgsX51xhscxbGWDJBJgikqtbCNtRFtrj
C17mXZCUXDsRBvJ2NypzR73Rbk1N3+7kPXw0GW3wmmMKYU6lTilhlehttjCVV59OKiFu7PZ40V7n
f2HxUKx2kXtS95v4cbf3dVcDey+vm2DA35jdE9HL7uxpz6ZXjNHOx+LWl0I0LnM3LMsKEJdoaYbQ
xHPV1njn57nAljYn8ZPF3alelGi32vUQP7y7PgstmSNZK3tNyHosZDHIUYvGiDp9MVrnxlSHgG0t
Y2/VGpgnvpzE+t60OOW60YzKk7Nobjxi3fiWFsPDcIBw2mQfitoZKtgXw8yj8cwd5CMGydPMVlp+
VhU4RVI4cl6UMGdN2iGe3a02nmIO0vYRhtUhGUq14/gYwfjy01ogEE/sDY76P42Rauc7p/aP7bYz
k57Q36cXUYmTlO1LOXiuVRRZVU6TMMKwvKAi0bYdzmu+j8EUh3d+634fjZmAa+HhfHGZSK/EPoAR
X7ODbmpNKd8lfCWJSND0dTQddEzKC1LziGIoQLU1lj+J27ySlzlnZX626DshE3A2NEoPbPMKr22+
vLzWG5ius2wnM9J+4Oyh+1QA82wKfEj/nXXVrFBFeRU1dKI4oNb36+9oIx9bHFpF3AEEqaQLhWHc
+7J8Pzm2uY6fUFpVv2Xa1VzoKKrFA2kd7IKRHPFUUDiytkMJknYavSBJkuNcOAAR7UIefEjXpTMU
2tu77MR51JSR02Yi0YdGIZbC2jmeHr30ZHb7R+9VLKP0AKA8hQSDaacx6gSeALXiQ7I4G6QJnlv7
FrRx3AON5tJVQP4MClkhrMXPHJWS0iAh3oC9h7K4jcwYTKFFuGYWXmNG5wA73mujz4uRlDEFxZPL
Y6sahrrG3nrjKqvq8Mh+p7ntclgBHkqmrOGiBDBijvi+YTzPY7h6O8Zv2Hj7tqVI6HeevaN0rxHs
x/E32QJOpakOc02otsSH2xm5DEAagS2gbUR6k/FlvBE6HVi1yCqqp7mDj4WCMiAzp37+yhtLm4Kx
tHPAwLMqRmW7T+/TGH5mJGxoCfg5bUJ+6gUC54VBhyh/Jo0wRLXaY02RmoI+yaluiTDkGuetijsP
Y11AfX/OmIc5TH+3+9HNDk3UHUvk+jydb/vRE2fbcAPXDQU9F2Ni0nrxNGikX5CCkQ77CgGMMJzY
I1FxTuv3ls7CFMCEAxQ19JTKee6Fgg0Q1n4d4XAkBppWMTFUnqKFhh2EjX6kYAe6xj+i8QAt3X8v
Uo41OzIyPeTgzTm7GkQS13QLK/Nt0Sa7ji/VYo8XxjAUqMVpFfi0X5XwYP59eird0TjivD7y1Us1
S1QWF/JcV4fBTXh9bIrVROvFLNhi++pIAWlafBCIR1XrRZo+Y9PegMYV182kbskjAT/kdt2+SMfB
Q6HN7jMy+3cR46tNY0fLNK7qUsab3OmJt1XCyKhJv0U9UgT9m1ShSjitjW3Xwe8jncnZJwkUqAIX
vJ2yWspgD0eH7s303WgwURJrZ9nClqEO5hIpNPxAkmW5imcVitSm6gWMKc9gjSYbys4bzhA3xgAb
ehFiJpzNjp+8MXvgeoSAFUE4DhpjfSPn8WO5X2S/5j8HLwHNZW5xV/7TvtetJ20riNVWNQBwI/WP
hQJVwg8hu+DRAfeI8LpEMnDxS+E1dFxkfZScAVYL30lVDlzt62rkAmWkmIfqpNw03MhwezQiSlsS
uJ8fMOsynO8JYD2Ul8+QYML/MilJzSFpJZydyLbBCfNPGsidIhzW55TND8gTsytAt39PCF2kdlF2
PW4Y7opD4LE6kqNvY5Y88lBxkaPnz7Mq74aAv1R0FUjyJnQzs8DV+mvJ91smPnlMs89Uc20gI/ue
GUNn3oZs0qoa+7sXVt/CI7+d540Bwd1002wzP9vhZhCYU0NXGS2mmDB8wunGWUg8+7ARBFQtwIib
+zfptCbw4Zh61yg4P6p65jN1znJPxxqXvBkEqk5jIJykVrN49w78QGD7NdRDyn4/EekyOfGAJhqU
CyIJCcjh/QS7FR1gWI30lY8DXHjdwg3sko6Us6gqeXRLgXoQtRe1JM1M3UpCpPxV0FrzFr16Fwxa
CI6Y6h+ocVUT5VeuYcAUr+g1lvlZz9S3use/36SM3dHcpoVNO1KBUF3OYLkfjEfPy9Qgz3AR3hkv
PyfGUAEGMDqYbJRp2+cHmgX6okDOOQ2U
`pragma protect end_protected
