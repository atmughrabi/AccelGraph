��/  ـ���ѵ�CEwS��B��s$��b/ާn�k��Z8�t:��8�Zs���%	�&g�P�
�|�l�V�<��Ry!�c��} H��d�.Z��b�2;!�u����ۻ'���j��/�lP_ba���x�8=�F߇�:�(n���8�T*����:�nP������Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9�㑜��8pB��ho��k�	k�ף��N�k��jL�5*����>�}"����6��$1��I{$ٳ�yqmo����4BC.+���}�+ �����mu�]� ui*>�I���q�	]�J|�����{���c�,&B'��;�G��3QL��>������X�W��ҕ��?�J��n�6Q�?X.f�ĥo�ݔu���n�����Q�f10R��N�S�K{�ˢ@h�5-���/��ʒ������_�~QE	2U����ט����u�<3����)·��$�?M$K�@��ć~UG��e�ޗ�+j�/	)C����|w��~J�X�^Z�(_4*H)�
��A�'�+-�=&k2׃����U���Q�N��'/2Qܧ?e�!��T��`l[�KD�����8�$�v��m��T�$�	{��D5�����{������"�_���r	���L�� sz,$v�'��c�(��8�4Cn���N�,x�ݜ��G�wl�����P�H�zgR�:�)۝��x�>/)�gs"���]�P�Y���!�6�<�]���[;�}͸¶�X`I>�f�}�o W�KRQC���AZ<���@j���m8��f�!6���
{�û�g���j�ed���>�p}���q��d��*S`1�}ώ4rm'���jtmw(���?�h"V���]��9PQ��|n��հvf<�̠����QN�d�n��o��G�D���6L�W����c������Ve�g)�"����q�p����E��3���jTy딮�