// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cY17Eg4Lhf6C8yMPTjeWB8/TIUpg77Gn5GG1bXFca/SLoIVDkRtZhFtN7A6OILcu
vuApk13UmS/VZsMmSoBqD1kxlGnlhDGZ9z5nSesuNe7BBACX/HMCgG99/WbIsslP
TtFjCD7p33dG7Xk68mRTu2xECyDbqWTjBrn8Ia+mbeM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1728)
/LoQBqRzX6rqsC+tlh9ZtJ1GG19MNyoG/Vu1DHeyfhxwY0pXK6UzxqS1AbA8HUgR
B4aDreFz8aluNYgSw2b9C2ukISCYyYUY6uyjOHYJ+nqFukSv4QcUfpaEpc8HcH6H
ERuMhXRHk3X1TUjLN2WpGjIlMdSnkCmsshpuR4/q2Xk+bMs1hzewc/1rekUGwAhC
LweWc1PDBbvWMxtIhudJ7hIbxDn3WxAO4t4GWrTiddaT13/yoVqCX6ZWuIfmX+yC
XGcoJk7wviUI3or4fr314FctsGDonQZPu0kK1L7yx1zz8x6f4VVTvf7KioTi9xhi
TPRelm13mcMhne0BI5u4d2OhkE2Pk8GQKavlr7xoc78H+lPmN4yNR67Q12fbD3yj
lLkYuFV0i5HSIBcwg8BXPgTcjzUtENTyyqSp2AIxdMs6J7sFhQk7pqjqsuxYSGJ1
Z7/xJBWfy7BMvGYCHY/HQpkVvjfXWEJkyCRLWZIAIv4GUaX7K+XZ0yMexQ3HO45v
/yzdC/MIOoiLAPTxP+TMOvpO6l1QbFSXyQPfKyesroyhryaBGDmw5jZZlgathuI/
pc27zirNCWItVjU0k9ixVKMh3h58ORkkiaIEZk4h+MuRGkoMLjT/EX7wGK5bEeqi
Xh7ggPhDCkJHMDLXiiNHR5sSJOcOik6d5mWqiQKZvYFvrjZ6Wh9voheWYXZ1RZMZ
lp3s9H06ojCQDPc15Ev5T2BylkGX+Dr1LaUnefzvxYd4J4noX5JAsvt6PLdBrLM7
a2hJe2h1iFeeLNAHZRm0cZZqzEY1ZD2o+73zXRUd7cvuEVJXXoYGahi3gYNz/Kc8
ri0AUyCYosT4hO7jXaW9wl5wIckzepxubx/btvnbNLBuD8xn9aM3YdxpUtU5HBFS
l8owbFnR54TKHais5JiUgYcID0z3vR5T9gv9XFTsFPJtjadEqrkJwNpltOOShC7H
qvzcLjvw5uXl2Z7dHP30J2wv96iFcv2iF+53oqYAY8KiH5zb7VfzDeZ3hDNwR4DB
eKtlP/9exRhxFa6M9ll+9KoJuZpQiS2vfu3IT8t8y8eiVKkmk1I3rZhgLDEnEMxb
xgo7I/rjDP9KmZafcc8Cw9go5G+N9M0e+pwUPYJ033PT866kuQsD73zCpbaL9TEw
8L5jXySdet3zBPIWuCmdbINN37v1dBOiOCTVERRlHDBKSYH7mYUGKv+VeG9FeQI9
cqPDi9KinPbHvGE+aHVSoqZ93psUT011xSjN6SoG6PnSd1ITIONeCam9L1uEBciE
4XfGnIucHpjkDMyVOOcTO/39HvdsOeLcjptpk2A2S5QAPMGgqb8uBp+RSAGFmVH1
645lFuY+sALD6G45bZn8W4zjpN5KlLMyLtb2zUL/d1RP/hQMl3fRuYjMSpDX2FHO
RinxFktRaLLs3WggJ0gKv5wkSyKWBEbDUNxqh2VHvftZ4lZz86ApESyzICeOYEag
L+6ExAAbQArLTs5kWkTvMOBcaHQINHt3nYE003HIzVJM3eJBS//CrThBkkWpEZA0
Tf+mIGX2r3M+JOb+rmM1B3Gm1HMDyqNk4iwaZjlFwqxoCQ+faeG4w8yr3TqdO/ts
15VH+lQ5O8zCDPbyvQ/hq1u3qfV/xTL0faEqHSET+2G+SahUm23AiqvAcu8JYj8Q
szyRDrbNxTYU+RTm5UcvynRNQvVkcugTqBfgo3by/E2ciDHfCQ4vHMlieEgxaKoJ
X0fOpq6v8Vi0nS/53WWzlZYrpEmXk14D+lBIJSJ+enFLYMCuS1TM0Vw8XJwrNBxR
0PlxD3xjrR8IrUFciv9LMUrgTIf7LXoaZYSienaYNw+gWCdh043PeGu4ZF0qClNf
3iiHCwLbz7DTJ1EUKVf6WO4/LpsxX68jK97sDfKqbM+5hWcovi7ROrDWzJKm0u7m
v5CWn5FlJLs2marO0UnVmeIN6sgpRWOSypL31tIEAd8XfM5TfDNf8KAIhTI0Lg5C
8+ST+r4yDIOjLC7PJFHPHHz8Eqzwpcm66XTuwpYjSDX6yWI5fx155H/XiQuAxizL
+UTDgqAf1gD3nXw7dBM4JpG2My3LNDaLO7F97h7msv0h0Gdd1KWFcA543tyvpELS
p+jlvgfgcl7/+X1GEBu/r//6qrrvzIgsNo41ZifAENBsB0uujTcOi3K+i8LPJDcE
BimlaLGkR8xDYRoM0YDqso3YT+vCDh1UJpeX1QYmXH3HWJmV6vM2n8kwy5CQx06b
QVK8M/oC3d8Rxv7B/C2/1Hs46dFhZHZy96QEhhQjj4k28BSq4KPFtGYdk5UoUIcN
`pragma protect end_protected
