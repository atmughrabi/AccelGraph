// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H@7FN'6?D%?%N8#3JL(M':O0?\_?6/4QEC]RX>^+^0C2TO'Z-@F>L6   
HSU*^=$WB)"(VEPS/[Q]1I1 ]3L-F_$#QO0G1*A).Z>0"89JN 9H-K@  
H@I0# 'ECX7!?OV>LOBJ@A*&33!EGI.M7"'Q?.):*)]XLP#!.V<*O.0  
HT'P2OWZMK30?#,TN">"U9-,1OUWQM>8<D+]58<O\67AA2 "'*677EP  
H'^$E@2_?37 A/DIE(C*KF_TPTTQV[;!(?I',<\8(QRTT$4]WKEB13@  
`pragma protect encoding=(enctype="uuencode",bytes=19648       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@-,!.I#P@)3E\7J-'3VQG#K\E<C/MA_CFEO!;?4]%Q X 
@#P]:[4OI(0/%1R0*G59&7OD.6*.*B5B2;4EZ"P/NOX0 
@RZJ+@;E2C<>S<8KW2$;W?4H5/#UX\+0_)H_&5!23IJT 
@4^[6?[.M\H@H0JXEJ^82T\M8&H>6O!6+9](<A<5T>&X 
@P*'@0&-*TQ@I2Q2U\^X:I-?8H%UHOFNI=O*T%?WB,UX 
@F+RX-M07L#GV)1;GU?Z:Y0.1\CPR[B=T6)JL!J3;93D 
@VF]BYE]_:@(YJ,/WNO#1EGLPDB12#(92 LZGP\7%3R@ 
@'J _'#QWHWXT+XI%ZP%CLL+ D82)S?8V#2$?)_<['KH 
@R4<A\0?\=B#K<P+6,D/-MP6M/,S'YY7&9[K"C,B2)X\ 
@"8'&M!$Q_;[V&\VV)2 WC(L;7^F-T?<&Y2EQE<EXNRX 
@5M3 -"A34/5"[9M+4"("\/O^Q#N^I]Y[M;#B_B%@MH8 
@G]5IGS74@V7$]6B$O]FZF9O'K?66 S/WX2O5BH$T.KD 
@'K\G%N<)N#B-%(F,@D3FV]Y[:Z7.%/\!388X2@D.^OH 
@OG/B# 3P481,>Q'+Y0^Q!F_WZ=TA>:/<QO7A;&FKRDD 
@?\U[ W-S@FJ^$LKJ WF$*I68[#%.76,K[*KD-(;Q'H  
@\OWPUY/N+ _6BHWFIZ-'F)\!KK;=2G/?EU"\G7,-0.@ 
@T].> D(80RZ\4B/]_66ZB&!O=^U>$#=@C4R3 'FKDUT 
@59BA\U_Y$X1U?O32V&%18W-'6V#U$S.BU;NVIY&?6S  
@Z%%TR 0IIPMI5&)86F;<+,R^CR!2X0_X(R9>*]D\S3\ 
@16EKO?/^6 /1BU;9;0"S8PG+,.;1[AJ1J!&R/!+$+)0 
@R]I(>>R65E;/A@EF!F^_@A\DK\>:_^@DA3O=<7%M1_8 
@[]#Q^G(;*KHY9LAXZ,W2]V0]')\?W 1PCD=M />Q=B  
@>JX>;LCL82*8RC(WM=)M%"]S@J]Y_J*VO(BK!'.]0SP 
@F5W(T054'PFI5K?3_7B0PEGF6%-L'2#XF(O,RZCXYCD 
@_%0PTIHKG8-'?<F_#Q4XB 6Q%4D:=7(SR _P.$\1*68 
@/4CUT*H9KW>XUEO8EA_EYZ(#+;,?K^0CB<K:CB9,^'8 
@HJ/VP1'^0R0HZN#W"I,5$8.!9MA&7E9/XI!4E/X00#L 
@J&@JW7>6>U^5L''TTB=-Q4ZS$I&^( C*,N;O9S,&,"8 
@^64.?UMWI-.0(!;T"O X/%]Z]P56?/'*]P!N*'[#NUL 
@B*M:N#)TU(+8(AY##"DCTPBJ3T(".GB5*BH-6C/,S'  
@/V6DUE"'!$QA*.]YZ9"K;Q51#Z8%#-;[6?K---3<!+X 
@^4^^7C,[J^ Z "]'SWTM4&IO;I+E36"57:-$:U?8GD@ 
@OE"%F(;BFF.,643ZA;7MD\0N M%4#A@Y>A".BH5:'@4 
@GHG0UN\6_B2<_>#&\F5&&K3POS4JBB<#D4YY\&V?&MD 
@NL..9+AM[WDT?7BGN*QONV%]HEC$RH"85UM)TVD1D:@ 
@VX6!BPCBI1P [W6"@@^R']<_3IQM]]TYS/*>@VMXH.T 
@?Y5TOG>9%E,3=-"2Y?$;G_4RR6H60GGM =(]OVZB\=, 
@R@,?18=&8.Q7 ,]O_R,.[*CV?)1@.8)(?7QKS.X7];  
@K!^W[29H*L.?*Q:3;AKI;K.8:#NQ?5>X$;CW:Q 6":4 
@ !7FY?=W1,V$W@1<.?,'L4X3E1V?=Q%JQC--U.@M*C0 
@$K9(4SUGW<=5",05-2K#J?!W49_K%F.RRF??CD >U[L 
@L%KJKH-*740%5+Q;N8L"J==LQE+RH_XI/J1CS^^ANG( 
@@N9K+S'MV5<(BI63E\C_IIW^\R*G[>:B@P[6JS;=!:X 
@@EA+&E +TS 7$$C(:R/4WPT/(<K;@E<1MY7%_ ^(US( 
@+74+,*/3![S?X,SQ1!V0@9W:CCY/&*.<)Q1N:,H"[P$ 
@])DH1.X3&$)0*6"8RTL[%M,=4YNPI9RW\V//,.'8\\P 
@I=E.'.KNPB4[[=C-Y?FZIW06PYA?(M?Z@/-H*!9;V]\ 
@> RD5VU90X79\M'#,^B7_511F5Q"*0I?-->Z5' N3<P 
@KXNWR11RBD$[5W,P22*%OK<>G0N55-Q3]^,8]8CA8:T 
@\V'Y[7FSYEDO4.;_ZP@,L!?3X%\.H4IGK;LQA?XY-H, 
@UE!Y9#;@A*\B*)N@_)B[>VHXQ,M5K&_?S*8^G-M=!M\ 
@6S).%)YJL1;M]"H$5T3$7P;%K2SS6_*H)2K"D@,>H2P 
@31F^/>WPS@4[5!MG1+D=D?P6A@F;QGB)$*INC,Y_^TH 
@?GP;T79_3%OIS]S:T-"X@">*E,VH)9A3,W:GE3GE2Q$ 
@T3^XNP5V4?<V=R2P2A&=IC@&>+S#*5#+<2@KZ*I/\M@ 
@;.<MV2B M 333% L@R%U>^LZ%J8_W7'GE6/UWO4?@,@ 
@@"(6Z#=9\6LBSN)-?BN"?1%U&""[D)_)A.S!7G@;B=@ 
@?9BJIB*@Q/6N-DBAJ&=@WS[4KZ2"AJ6+G/LN,FV2 "8 
@3 %\&NN*<G*^GK7YGURKB6L]J(0X7V8=OL.DK@Z1L&T 
@5T^2&[.ZVZ=6JNT!.1)Y@0C^(I\-GMR-/%)3;KYQ 8L 
@07O*X=K-9?WM4W5I1E=L\(><!])17/XC 8X?Q"?J@Y0 
@9%G5(I0C@3$@^&"[_B/^S1E";UX-CNTS!RQ[J\,STY4 
@%M);F_<QZF#13?.D-SM TLFTW=9C/ C779+"VWW$.=P 
@4=_*_'Q>.>21P4T]>02E$0G4M/46_<UX*1L%^%G"O^$ 
@>Y@$!VM1]MHCNERGE%*8A$<_HGEOY#$Q_LZIJV6GE"$ 
@#_ CK.LN&UD$)N'62WV;L.]$-\SP-KMIF3%!6@RN;,D 
@N4!@!$AULK$W?WV*NU5*8/V<[RI_W44106T@E@FQ_=P 
@=[,_RE'M!71WZ#^?F1RSQ^T*[.U=+4NK>/MC'X!%7?L 
@=>VG9-_ .C/L4<HARR5]9Y2;ZJW^;!ZP%RZ/F_'KZ_X 
@R(RG@#W.K!&T[AG\AF)3;]@@%9#BZ*/),6+ %?RXRU0 
@BTT0, K5$_UOTE<"5NB#K/IG<[='[G<[2,&ZT#;02JD 
@P6U0>2TC4/)';R'P93VV"V-OZ.)^AY)L^I<]F:QBAK< 
@KR6\_0_VX^W,[H1 5]B(]20@E!FA.2^5\@J/>IWR6N@ 
@I\R/H8[)LS:L$7S> +QR^2@*VGI+(Y[W)HRJE#@N''4 
@EMGHZ]2@\7ZD(_X$,_KY'V@,X2#)RC]G9HL(M.$^M.T 
@6>GO+B$.D[P0KO[8@W.-?2'4^&!]?^Y3'&F3_@1E;.T 
@Q7U=3J[B4@%#TMEYDH5\;9/>.#^E00.MD2@6DU=#5VX 
@F:AEJA<!$*?3%-N(Y#%^>D<3SPRU,UXE$A2;T(# "=@ 
@%-.7TZSOW(GM9G5;8A 8,/9^A#J@S;)#[K_#IHEK370 
@+IP8@VO]''J"3,5!J9I'D)A"[P/L$"Z76$S_7BMZUB$ 
@AW4?S,_P+B "#GOGYAY39P<\YQ"3+D"C^+M8VG. RY\ 
@<ZB-E/E.3V:7 N=,UY;"=V?VQPW]=7*JX3A!+9'"[3L 
@(LB)#S2*.60& +? .2!\/.\BKR[PE1!WJ5TY0W&6B/$ 
@TY;ENLT?ZX%T44=?^494&?TG51S#8HSPUD!57,'3]TT 
@?B^_\K5EZ5DD_#B>_2!0D9@V*HIA'J$;Z._0&;"$BC, 
@?0I&!P5V3:8X=U+TV70>14"/H40TDV";O$QKE6N1-9H 
@HU+:IJH8U-%HJMV3P0EU+M#-HQPW'[?$FH,IN0Y000L 
@]X_Z\F"]*&XT6U&;.66+7?<6/"_^FBYG?89W&U1ZCAD 
@CAUJ3ZBB62G]AR\9;]*]^!/Q)K&\;?L&[GW0P3(#?!X 
@O:*C)X ]FKWXONEWU.U1S^@"ZNZ;=_[,4)1'=T T[(D 
@Z57HC6[":=DE4=MOUJPT/?D'WP]4L'4<9G$*\+]._:L 
@/=N?2;*TCEL?D,FPXD%9>M60X<,&(KC],_\2,Z7[YIT 
@H@+Y2[>I?[2L:UFU'86Y)4O4+D$@L*R 7N8]:OA[;2H 
@*K\<D0GUH#5H?+5>G!DGJQM[LN KF#H!16DV@"73#44 
@[H8V@(-D]M>NI9@@CPND&X<1V?3;7<0FV$.3MB_:4SX 
@#9B-G*?GOQ61%[DW6#.P=^=P:O6QYN118!GU3+&Q",$ 
@  M;WVV=(-QZ ECW<B&-$#NY[,8],T%%."LV)4 A4L@ 
@3ZBGJWW@YW)9/ GV=]DXE6(/>MFVN@I1$*V6H.'ZH9D 
@47:O)4\4=2#(1,X-!SHA,WP"23N)QGI88+.K(HBXR5H 
@ZTH#:^M=-D;VJQPR9;SEI$F33TFCN=;N>'Z+%+F^S)4 
@TX^>)188, OG]%3*A2FD_=/I4#(0^ HLQ;Y,VOZK_@\ 
@^JT%^0V=^DUOA;Z&'&_@@ RCF=&9N>\MVVB\RFPRT2  
@W*W4Y)LP'V#6.XEL,J5%";>''<J A)=Z#/SZC$ND3LD 
@U["U86=_H$$8\=7Z901U.ITJ!U+XD$>ZRBFP]'U?MT\ 
@>EQW"D>SQS3)'&F+A-_D.)%;QA/J1?_00R/EZ1_(*1$ 
@-*&>!DY$G/#FNFS2-1C^F%LX'6S*G^8AGMX?V:&\Z5( 
@]*G 4DV:U4/RJ5D ;8@3@"]WRE$=D[/O[$N^NVBY"0\ 
@A2PW<B%\9(9Q>7/T;\!<^7-F 0G>18L/:M05IBI7!=\ 
@D0E=,22&[_M;"@7>2B[4/V/Z%<PW)?5/:/IK...L^)< 
@9CRJX+(C;0+D"DF4JCK@LO5PL;#O7B8/;Z!RD7@W@*L 
@K.TWQ<3WPBL6ZK.T$#Z(S?Y4+A*&NNU*ZK!#V3(:G84 
@_H&YF$46;/(F:Z&HB-Y*!S,Y/K_GL_N&6C40M)$^.L< 
@8U0C+_7D #4GFQRYU(##'_A+I-B .?5O(2,X+"BRO?@ 
@Y7!&;/ SPG4S_BFIG290,:A-J**.](&!Z6!Z0DY_&^  
@#V]_/ZX9%4M9Z%0\T:)5'MJT- :.HHCA#R>P!GCNB7X 
@#KP:&Y!O2TUQF-O1O-BFFL54VC@Y5+7\5?,YGC/[8T$ 
@WPN>7B@7<^ 5!QP?-[MF 0;<R@!=3 Q?9^H+2S)TO]@ 
@V,*4CV)DMXH9KC?9NV8!8(Y).4^ONV'ID@"VLA[6QP8 
@G.4+2I@H4*R4<P=[W +I:EU$53DZ=XAT5-N'I>]D @8 
@+5[S:AF(<8=K4LSE5OXJJYL%9>"E]%6$=9$<6AIF5%T 
@.X?S_T\X?6*\Y(U=I_9^R_OD8Q]0-'\%KD:@)GQ_-*@ 
@*HV\)ZD<+9< '>].:&NG9KK)@9QWK]?=<]M0,K)B$A0 
@I2FK(E=D<WE,*JH>#R6*0_X5P>_B[Q9HL$T#?QH6H+( 
@U# C$#X!6!%'%@/.85I?#<AO/1)(D4M*R+.HFXI6R=@ 
@G9'3?<'@_ZJ*9L>Q7;GQ=U*+891T?*0<+Q./HF$@RN  
@SF-$.JH\C*>E(GK]]6R=)Q_?]4X;5-]RS.<3E#YRN7$ 
@4L[AK"J@5?7 1L%!A E08D#!A!_@7-9W3E7Q1R2!TXX 
@'C8B$20]?QO6[$P50ZUFF"],I,(/5M%45:FEW@:\^[D 
@97^E6V]\]BD6$Q@B$.*_+61"S)W"I57W=9UYW%5%3JP 
@[#$GV9OE1HG.OUUQHN(/#)JVSV&ID^S_7I,<3V9 #.P 
@<5+K$'G)0=(W"GB\%_^2*7ZLE###I')2I)&?=/D=F%4 
@/WV6EV6KF_]\.M1X%3>OVV*PH"_N/5_I% -FC'6N'1T 
@A8D:1W\2="12A96?1'!ZDR?>9$7F2Y@#!:P$EUHSA\H 
@D#RUE#J_EB52#:UD&7E-I6LK9Q<".&J:J:^7I&3,150 
@?&3:NIE.[SR?Y^XVOOFL1[8":QRJQ<)W?/^!Q66DIID 
@'MNFN=8%.WAU?@#:$P9Q6O\8*W+C[:H0W2J,U4\3W/@ 
@*Z&V<'C2(O;JPNY2Y"'S^>)+THL-TLS;?I7@.%##6_< 
@G]48H@=GB7(9RYLI;NTGH46>K>+OQ)?7QU5E]V?B\)4 
@9+7#+-SNK9M#[/TD"-^ZAUQ5K74K0#==,4;<'5-)USH 
@$AF?H 5=-MN0"K)L^IGL?+@BNZ&U];*(<(.@(!N%@B\ 
@S+.VUE:OFSS*E'4O7$ SHC;6/M-&KZB0S[DBZ44"YTD 
@21/PKEQ^:_R-1$WK1C7P>,]R]I7EK3YS)OH,F D>&%L 
@(8;\ WU&_?2SREC-949^=E6OZW.$,M(ED;Z,9RJ/V2< 
@^S6\GP6^#-[&B*#HBT\$#@+84:& = AKD2L.('KM;4  
@J^3TA>OZ3:/M_$^6R'S%+U<P;IH@U:?Q5PUKAH7$L7\ 
@*!.YM4?G0QHM5 G'"TX!918J/#E:$ZCQ*-/%+*_8S1\ 
@7/$BR<VH8_/F-'LA45_;G[OV@&]:641PM? X7VRZR?$ 
@5@7RK-N4*88OV5<I"P=\<U6U==,,<%X)0MLF8XNRC$T 
@SFK\PG/7ER21+'#67="O@L[W3N.X2]'>WP@=9?84 +T 
@<?G;M>FG)H:=(8*,"8) 33ZV]>)GY-SE!L7-4)O"Z$0 
@"/:E6R'O#"G*'$X$9BC$'0!!!MV*+ -[)E%Q%>=SAJ$ 
@^ [;<B8#H#(4XG&_ZRJ"REW*B@V@Q [L38C,!W9A<LH 
@X =N?;6UOJE:=/%3.>F%.E/8ULWBEJL-.<5A"503X5P 
@OT2\M"&(/8!>N82_/^8R*6Z\;I#R0HBC3(+:4_-B!U@ 
@HSX9J!>N9V7-B%UQ5*F'%\I9BS'#T/7+ET\?;UFGNO4 
@(.T4A S(IV(KC\J.18<>#MG4Z),PA;%,C#8L@")7//\ 
@W2(L_N0B;LXD%%_PL-HE8YA5S$ L?4+9<9;#/4$L$WL 
@\'PZX :Y;3&TQ&J2)NIAL_(%;P").$#*=V&EOHW;DK\ 
@$Z/ZR15;QNQFI#31;5!($UZU5K.36!>-2+S8X6?&C#  
@%M4*\+UOP\$#>S9C+C=P5ZT% Z_*.F<6Q74M=J6H-$, 
@XB0])WQVTTV 7JVXY@_A8_.)G'GX'=68,6XYW%#5F-, 
@[1%SP1R*C8P>E9 G.P3(.N>J"KLTV7IOH",$#(\;1EL 
@$_<@&0X= J^ \5SPASA\@*@'X< X\C!=JO3]AL*VSU( 
@Z;J?B>KRLA@-UK&4_1^E*+1=LPWPE<,^[<A6YN&S 2\ 
@\<3S%Q020%989\J0Y0*1DB;"QIS)A1<&U2V@&&/W*Q( 
@/=7T\NY1X79ZHH9BA!]B/"=>VF;Y8W<D("= $MV-WQ$ 
@<&3O@>;9S)*X)(A,/'<4^Z1"!FU]EKX2+PUY0M.77G\ 
@I2<9V1= DPU]6F/>)]R2X\H&8@Q"#7 !Q"GWIXFR;O0 
@[W<<;E[BW7\3YPM=42+7RI1*TY=$^ 21;P8A!#<LKHP 
@.0E1,"[@U=:P]6T_:>^S]?1O62I>D)$$@X* ^RE<I'X 
@L0O]L<IG8HY<';6Y]E7>G9NT$,PJU"!:)+Z57^@4?%( 
@,W= +(M=U W(9-=VY-2KB1P+Q[W6@^>*83(KE<FM&&\ 
@0!0U/LA\A/ < JBRS%14XPL94TE2JKN/L.N*RKJ+[>  
@KV$_F^M34KUE['>WX+M\5S59$TKW^KPAWYQWB<%7&XD 
@D>)GLH:D?_^<KHD!PHV*4]T;3WRV$P4V FCDB,[L5/4 
@S1*]'HH]S)NQF^0^766/L0%[IB?A1"O5ZQ@I2U)5"Z< 
@XUD*!_&]S,BQ@;@XBLV,1"9S7]?O0?%;AGVNM>V2IOD 
@JGZ40F9< B6JRHE02H&'QPS[N$ V8 YABK^3_+^9U,L 
@JJ842KKZQ%EB)61'>')9B2"D7KI/']G3YE&Q!*!SFD8 
@'2TB?VQ3DJ]BW-N/^_3B3DD'&M,YWE0CYKI#:8]7P/  
@*IO4"F9U0F#8H%O@1\;8EU%XOW=*:?O^JA.S.I,>+E\ 
@YD7N_D&JP-2LGEMJ\Y=7<LEK6#B@N-,%NT1C=@0$P($ 
@W#>7PDS=PWJ#2BZN0'<[UD/,F<X*]SE5+,;&71=VH0, 
@>?US%'Q(B=52%)?&5H+:6_T$,UHO(X,882F0[*%&HUP 
@:G9J>Z<&("+N:,I_6PAJAD.2T_X][PLHYM5 PZXWO3\ 
@9[T;$=_X5!AQ>0SJ-ATDT9J4D.DNUPLH@.#07"?!0F, 
@9DF'S;,?^Z:U7I/\.)?_#YR!)[[!@TY>.]%JT7*KQ[T 
@.E0,5(?23F0_7J+1,"CT&B=TSCG[2IX^NSV=I$9"@3, 
@Z'7'KU1G),$?Q")$N:5Y2@[4R*")F 6!\,!)$GQ_7TD 
@)]%4G,4]8SX6@V:1H(V'4,'P@]EOP&R)XW)A%$/VL)@ 
@]!@%X-C&64/"J(YA@@E]IN1P0^0WKVYN09#+1"M)8FP 
@,5)$E3+28@]P>2XL =/^UVP_YD .$.B8/-BK)@/A>K\ 
@%-5Q=4[;1?L8RC[G;:/3-&8\CD07;<.&\UVZXR;<B:0 
@'R(<",AE[]5+JS[^E*Y)]AH$\+\YAC;D!X$[5L8 I(P 
@3/T;*9J2X)$KBM;, $1XJ4R"LB6ZS3A@'6#_S_0M'LL 
@Q0Z(/;!RN\'A<X?"37:\P_-/!\LWJV#9*1TD3, "UXP 
@E'IXIH*TS5<O&:D&S^2%*W!Y?G\LMHOAD-6$\16O0E, 
@#S%LS*=PL,#OK;SF3O]:'6LH"Z:N6!C%.NW0/DZQSD8 
@*7?[Z+8J['T<RV0]!A+1X^N2%Q>9&#>%YINA3;T/IPX 
@!%GABU2@ZC)?A& HO3, P?(<5UR6:F;BV%U1K(+ZQ?\ 
@Y2[&CY;NX3X+KG.SHP>_/E2T:S<T'^D")JK=*ZEM,,D 
@N^9<&?T#41#[JW&PO]3Q#M.9F4-S[R4+Z>7]MT*/6HH 
@WPD7TZNUA76+&ZG5<'EVLF]_ ')6?0N/\&;E<R80!8D 
@E=G]">-V4'NX.$WBY#>N-:;,R6=[!KT9<(27F2O?$?T 
@*=4W!@,(1V $H^32*]O1"A71B]>D)3'-J$'TP*TQ<V( 
@2K4M&'K%RN!&%C5E[ AT;Q'QJ,LP"[@5RLBR!W-":Y  
@204AU,D YS:PCLXMYW&46+6YKT-5J>7*OK67L'5-T=T 
@6N]=D*W0G]%=?SX!RSWO[UJA1D :.V61H=6)"6%=Z9H 
@0'0'(D7:HMZ(SH5-OOWPL?;@@WSOV?2WHV]7&E38B9H 
@O$/R]$X$4?G6]\#2TNU1*;]#WLS53W7,R POK(A36\P 
@OV'^X+>CXP<**)>1@Y9>B_5VD>3E+-2^A)NX25/NX$< 
@H:H%X$-EWT<5"*.1@A\$\[_(:13Z(XM1N@I!-<CJ@#8 
@MQ0",DSZM#)*"^L, H-!1\>$UU6U0 Q#\=I$=B'"'Y0 
@EP@>2.OD4#,F3H.#F#8N(WSZO275(^51N]HX5Q<-7VD 
@:C"*;U K"^J)RY3BH(>)>S@R"*$E&TU+5C_2OM(7*C  
@^\&Y9^7=+OK22(90$9I6L=-:PY."#X/\<^!I#>PO*B  
@\E6IUV1XF)@^>"K^03:R8JI\U:/H"ZUDQHJ]]S2'KR$ 
@^,M!$*>HIK6@[R,=O!QQ&&NA-"G7M9VWMZ-DJ^?/ T( 
@79:P^J7S&AG_5O#I81)UFU!6[/V-AI[KA8GJ9R^)Y6\ 
@*;T?1!GA7J]-AB-A?,= $#E[0RK0# ;-V(ZXDQ!^%$4 
@OU +<5.'$FS4[DXN0MW[C>MLIY/F(<.!:K?3?M82]@( 
@IE"A%JX>@45+:JM50MOI9^66O[#E-2GLXA,+J,QDG]T 
@&E%GD*O,44%LMPFQD\E3&3LOB$D/G52"]@2%!JF_G^0 
@E8!71,TU\4CFE73;@78JGP\>78A0\$B=>JRVNV]UC7< 
@V-3  C._S)WVV(NNC]$V"2Z;2Y)N<4D13-[L"Z_NWUP 
@+CEUGKQ.^1'1^:"3U.<4-L-:&GRFXNF42ZS1RH]I.+8 
@C;&K(S%.[WX\PJ#1:--5BL37QR<YWJX&$OH8$0S5R(8 
@(#0IU\8/OKR68Q-8D J1+-F!&T[^(,R1@SIU/A"*HC( 
@+SX#KAM-@(B< !DAYHA1B$->](-R"2 EGY?'8K,0!IP 
@G2JC%J5T=>?)%/="6;D9M!P>E'/AJF2ER*VB4,K/)(( 
@KZO_?BJM;PE]^#\ -N(6OT)/">\TWYXLNB:@H9'RR6P 
@K^0,VD*BW30G9/J43['=OZU@<"6]RYZ"G]R(IH6:^/H 
@FU%.Y!OJZ?M4C?$YG@H%]^P92P>)6I6\UNX$5PVH%[  
@'0F#3&69"0#0#^"$M8C5>6'N5!M"+_P>'.?@W/83UZ, 
@%:@*C11?7(R0IQXC-%)3G!3R*Y:5G+JLNG9-^V8PAL8 
@#VC]S4NF$AQC,GL>O5BNF()W(I,-YWR1ERF*P#,GN=4 
@+Y9Z_G:_+#V56!4:_3!$)OO!='!@JXY?!V,%V^]'2[\ 
@\+Y9:4#C$BN'A.[9 M:K"U9^+>;^M- \D6%O/'9V0QD 
@4$P4$3@%@03/B5,9>>I39D;:CKPL4P$#B\4XKY'M4!P 
@- &"04-9L=EI>2S,O CY6(Q.NV+(35V/NCX(F^EI-"T 
@%P>6N)Z*@M8G#2VT]_3/,]FUFO52%N)4]?9HL3!,&]D 
@).]/[&IQRB@' /J0%D,><O*@7C(!!36#FW332C1>2-, 
@X2T3]#B@-F)7FKC#=R"SVFN=9_8PR=-ZM,W#=9X%@J< 
@J:1Y>QD?AK\HZ'!Y%G>;)35TF<.Y BUI0C).[^?LAQ  
@P7"/@36EYMDT.6.R/CM&)L*LB3;Q"Z[G"_,X]!".3H, 
@N7&UK7T)2"80*WYD.^^J^W*$/SJ;7=J :2+#JJ$S=JD 
@)H3AC/D5=I5SLMX<LKBM$'B*04@"S3L'3/&'!#4AR-X 
@J'P&RY*HJ/NZN\HD!=3!7&W,9"27K:R$H"#G((N),!@ 
@HH3+W=<1IF]SK^8^G<)8+=#Z10>M)A%0HYA)&29:LHX 
@\)9,<JK6N0%8ST;C9_*'VH("(X.*MX#[_)'<\' P.PL 
@R5\[889F=0"&''&).!ZC&1%QFA6" .(_N3MEH&)LDQ, 
@H^IHZ/+A+TY1RKIR8C*=V00:Y8HXG:\>R!G@6]4KI7L 
@VRPD+-Q!W\H#?2[/Z$5P)K\Q.N0(6P=)O2(!A6:83)@ 
@.9C?;LJ^91CQO+XRHN9\XV=K3NASG#[D]2@O&-HW,0\ 
@KJ'8Y'MO4/&2[:HP(ZU1>2YY.3ABI71K3.-J@< G"7\ 
@'=OCXH#K6$8Y<:^PK.0?DB19-XEZ9DBDV\S=)1\["4$ 
@NI_,AO2>.:7\;\HO[,E"6N:8D.6:!.);.<S=1EL$3D  
@6+5$NJM=K#SCB"/\8%3 _3O(#-':I:K2(&4*'+>+/-L 
@V-IS270754]F%68#SYJD-V?+-16#$@RTC(N:/^01/CT 
@/37NK(BT$X8 G^-R_'=FYLIM%59VH2D,) 04G'37P.0 
@5M:K]03&9[+P)BD#APS1KC$6G4+GM)J5:^'E+B(=C5X 
@"V37G&D6.\F@/=G0]++4>DE*NN,JP 20JFL?Z1KKA'\ 
@*'O$7U7(;GO^![8R5XAX72$X,9 J(2T@33]E+M"OBH0 
@M:)"F.H3V/\18 A77^.;^?4%7B%#KUQI^B,-&/)I*!, 
@GK%=WJ:XP;4+-;>*?() H>KO@WL4$E:AF7#/ :Q)V]P 
@SOE0</+$!]DSEUF<XL];B$K:E?5)^&XC Q#ZZS:)DF\ 
@.@P./5"E10\C'-GJ#[.HKVG''.9OIA>R9:IN\)'.,:\ 
@12&Q"9[U:ILL+A9^1Q1I3)(XPDG</7W+;8Z8TPRC#8T 
@J0;2A3).VJ8JK:&JDLS =$L&=QF@J\3P#U?VXTT35?H 
@U2>U3#=6,*V.P[*C5QQK3#8O,US$;A.>84"P?0$O&,T 
@JD!B XIA)V)9X[SXY+0%\SM38U</I#5XG< W6]T34,H 
@W$ HUZ/L@JCUP(#<K%B(<GA/$1CHU5DB?36E@:41G;\ 
@<X..O#@4Q\(3+2 KKL]E/*AC#/4F^]5?X-S7^8\T']  
@N:-D=/YW@%P"N, 7$H#4G;53EQA0MQX5.KM#?5'+DFX 
@#8R1Z%)NWA>3OG@<R\_8V@(XM9WV=$V3D!9^10!L!N8 
@SZ&/I."]S\LEGE0#!XGST1B5O(FP&'@WQ_W-)SW#SOX 
@]//8,^KTKW2\SZ]-<D!4"'S:O\?5OAULI!R08O[KABX 
@/'E#'KWE950AK?MR;]D2,-CR*R=P"/.)&O]BS,&,J9( 
@-;.SDWGR#2],OG'71RTD7'7<[UZ<G5B[--6\NFO6L<  
@A(-N3$JPE&RY'&FGV<RLFG,S=6VA&41D1K8G*&QA"#$ 
@[,V[_;G'"Z[_VFU+4C$UQ)_FS#1]L,G0+;Z^?^BB(TX 
@NW3:QM4XU$#1G2+_=,EC&*A]YXBV7*.MG%H[.015?5\ 
@FF-WJ'2OHCG^"3R0?%3ME>:H(,I;ULAI%P\N9<YQ> L 
@Q7M)*I\&R >NF=?2[ KAP 0\:E\D1(5U/H 0G6; ;S, 
@7Y=7T?*EMZQHA\.0QS@[$ !YHRR[4]GU"*IH[59J7JT 
@:P:<TEUB<S9N\F<N=8+R,EI)L8.=5R>1Z$.^AXO!V;P 
@59_8+XJI2__]I8:VB&7A*W5*KLKM #<JI38K81+".N  
@T; 2P<]UUXO;1[MH\$U]E>>V8S^%)F91KJK5T,JF)^( 
@ "ZS*+F'B14&CTP6"?VC;9K.0Z*?P$/8U<#Q8:_4S7< 
@TC>;1GAK]&<9%K+42?^BD"D'0!]253*[XEL(_ M(&,8 
@VY,ME+N&TR8W1/1>2DQD[8]B^'X1/>>[1;Q(P]>9Q4< 
@]&(?0E.97(#]1O5RKQXF?'4UE$?(('D$!;)]+0CF1"  
@=$W=P%@F74C<.O0>*VH0 5X1&KS3V .&M'(,7#%Q748 
@!T?>>\#S2KA$Z<SN\,>2H# $O)??-'AI6JR:D(U=]RH 
@DKWD<D.&20[&)X=#C?BK2"%2O=&1B'_/"S(^?6/EE_H 
@(04$7%=>/?%9H1QG#6?4K;QO[<50#>J] R,Q)"Q:"4, 
@S7"M4V#DEN@))UX2![Q:5CH/.B!A,@/(<,?B"LW@89P 
@&@XGCVCT35IK6'IDH$H$4S;)=YZ\.KI(5A(,<R4WW98 
@SRE3W@/_ WWEO>N1K[/HEK8IBSW/><8GM!5AKO*0E1$ 
@Q9&LWX*[PQ8(E<V5,,J?+0#2?ZQ$;A3.YY7^GQZSL2X 
@T>WT1R$6=<U'N!8-QU/@IB1D&K_[-9R(6B82F\OBG), 
@DFG61[TP=.&;FU_HV;_-6";K ;7N=&2@" Q;T.N1]/( 
@3)[E59I\],D2XXO!9'4 MR.C82B,JZP,SV-+K,YV!7X 
@G?)4_@])V;L !IYYUW%HK=*E "H-[6< JU^G/&Z+05  
@@@!CU"T77Z?",_DDQ9 C+V?6\&Q^@(1P*X^>TOT'C;H 
@T6PUTD,O[>3<8FG!)<D6T*]T8SR99 ZZ1[$8;[?6FSP 
@PP:Z\'E@Z[L'$7M8*>T2-EX;<9&ZS^*YZFPU+S$V3BP 
@@*$H7:5(Y:KCAK3IFKR4X>X#T-8:H)ND-^=S+J\=X($ 
@<OJ<$BYOJJQ$Q)J2_*Q@!I2>\D]99-M4=5=<N;'[_!L 
@_[T9D!."2L+'_[Q(]9937#,Z,2"-FK@AE8;V-/V_LE@ 
@QU6SBNG_4.$7PC!()1:BR%*I@\;&A,%'59P1)&R(1A@ 
@2,YOTV[Y^?0!12^-F)B=*#NNV@JCG[[.>J)N$\H_9Q, 
@K!=R%<+XX>OP1'-K8R(U[=/#&\VUL@O-'RY-5-W./'0 
@O+&I=\C4[?-LI-%RH]N9_U8>'O=:=6YFUTR,&ZG"@\@ 
@SG071F-E#[V()>DDMCHD*2(*A$#& !>+Z5OEQ5%AQ3$ 
@#>%)+]H[T*,6 K-U\%'I!*B=FR)Z_0- X# -PF)F1#@ 
@U\X=6>P.3GB(V;;Q :E_DYKA.C-9['C%APMDK_P[0V< 
@W?(IV9)C:NZ9>R 5I(?Z*<(J6-Y<<D1S_.S)2EJ[SZL 
@4SD:WK4V^3/79=H5.)$&L1PKF]NO*H+"G9T4BU_!<OD 
@<F!E68!-'^F.'H3SD2[JZVTK9#\BM!ZYG1!J3ZT^+7H 
@^[^0Z'O84,(#U%)G=_]9W<2%QZ47V,ULB'%K(@M@X9P 
@,^8K X=S4\R?Z \N\^!=,^KRB6PO(,73?T$!BJ!T3W, 
@J7>#DI=SRA!_T!O:_0910J3S((130D?,G+Y HD,[9B8 
@9/UFC:6LJY6I)]XI=J=8=3J,_YX@'D$>=.\2$Z:>2?0 
@W>:?R,4:-UFH--V@&P&VC1!N,"/)7CVJ3C!Y[1NF4M< 
@[]F[C*B#*" 7#M2@YBY9M+E:GM6P2<:FP2/ZYK?*#;T 
@,#0FNE'7QR(L_X')"U]AE (Q0+D4OCM2@\95:3%<W]T 
@H-PM4@ '1@^7_9I?.W1/?&5MLF1S;:XG;UBQ1RG_+O, 
@:/F7CR?#KT'=GB9;80/)01K&050.'%!(/(?>6K^GE>, 
@\-[@*JQ@;!!TG=1HAN,;46,:>A;]!Y <C*?*?0V /_4 
@8%G)<)5HJ*L*2-HJT<.#[DD<S[K\P#G3Z-LW\L;'/_P 
@08*H:V91:-_8 81=\I97#&- :!JH.EYJW>;"&#08ZCX 
@W[AJFK>DRKCJY#[70\"7H"@W@22J3?94FF41NDRN3^$ 
@,)F[^(6&!'XS_8T3PI02*J)N']M=9PZ'87*7D-#DM6H 
@1NBX 8T%_XD=SGJU!A@;K*[8K\<$E\^G+C'O(N;^[', 
@((=\_],8!R!_YE$_'13UM[7 0LCX"<@*:;+<PVI(@%L 
@;<0E[I/F%L)>!13038P[<*A,M! B@1M7*+_7(\)=)@$ 
@?52 .'\>F<%9-R!Z=<O@=2<M32M/?W<8N;!L6.+E(R8 
@1Q5J7_<O30VJF7^%_,FKFX#56]SC<=ZAAT]$<%>K]($ 
@]7(=A!VP7'5,P64U-JLL@>K-R\W1%9UQ)J,(8V\>_.X 
@=6E O5=^J:$.YXLE2<(MHLT]X>#IG&5@QD2IR456\$D 
@&)CAAT=5PB2.!QN1'D/V6M6C4BCI(M*0V^^2_:RH=*\ 
@!,)-4(^H'MIZ5 Y6S",^:;:2LWB6>#N9L:\ >K[#\#P 
@MB0??,7MV8WV>6V>2K='6VZB73/ZJ!9(,[7[R!O\HP\ 
@V.7\,N&_#=;YL4B:P7UO&.1?;&[%ODL("6_YM<4W"8\ 
@'_FR5Y)&0+F%!T/G,9((C ]5+C!N:X:_>!+IE?Q(8A  
@SBJJY?WT47;1S-G0X<QW\M73_]#V]1^;;MFLX484WI$ 
@U31!. _R0;G9M8H5D;35?@2GD8:QWB&3+X;12/Z\Y!\ 
@WDX-%.:?@<9^6#>,X%(2]!-C+<DIK[A@#?0TU:YP!'4 
@"ZL*>_SG<<YE'?:QU6-$'MCLGC0K SA@:ID0;5R:3&X 
@M_(R39'P/#/EW^TAF O.@_#MN'<0B.>"#V?!?80V?I< 
@)DN/N/W3 *I8JAWIJ6G\J?.%*"X$D898JLF!>4A>S@H 
@5^C>7#P2Q+;O<_?5\*3CI:'X&%DIJ8.C"U1F1LFI&:P 
@PZ"G,4 %SKJ>,[?@'VX'+$MMQ@9_E!)">P<1$EQ<FV, 
@EHAJ^RJ4GJJ:]CXB<F'2LI?T4S)$SPZGN_:OKA5<$W\ 
@9!:;"^XQ2"]Q1@Y]-H(?ZB%NGWW] _LY5'\6:*^7@U8 
@:8;[3IG5?C%=^5AH,3)&2]Z6V;A2_^X.NZ-.V)ZX^CP 
@.UP@)-]CMO2G<,*NJG9U:O4^YH#F%"@E0+UL""KC(!@ 
@FB\H"DOJV>U,1TXZ:95+_=M[NS:LU]PNNMR2"_YCU.L 
@7F,Y(W*FK1OY$?]#.VAYU*\8Z6O'*Q-"S=+<9XPLMP@ 
@()2,4&>A*2O?N6+I79*\7'W(5B::G@WXU6B;JMO^T*( 
@1G1U*F&\<G%5P8MZ4OJ'@8%-<'_!O3SV^MB>+1('LG@ 
@ENQ&:87\#?S3T7YDP.PU!QW[5)";Y^-935"6!6NR.5T 
@0?"_BZ?0'8LNS7)XJPIH4=%3(S::DV\W$^;>\,H-"6P 
@KFL^/_^COAE>B$N7\[/O^P^)U#2RM'"J;K@_L;;5KN  
@X02!VR\]1"RY@":D0EV =@/_P5;HT_N(<VYTFC_/V=@ 
@;PU=:HPJGEMP+4>U<A]N'CDS.^P@9HBU\WP@Y+]C;PT 
@)V62ES2L3?"J&.AO%4S83TS+F7O@UG/)&>0\Z>WSB;P 
@5 :V/""#ZZ6^Q#0_*]^-G/.MV>ZCFP%B$.-W]-N.G@H 
@BGIIN59%HQ"PZW>-H]K]QLP 1]R\U;1CX^?8@(F[D-@ 
@3>S2^> ?T44MEKJESGT4S7Y-R\9H_4?U1*#X7;,5Z!L 
@'TI-Y/:[N1GS$3&%;&G[;+'%5<#'WE GVRY>]\N\4+8 
@98JV"1:;2VP5=0/)DY>(:"/.(J"@EZ^[1@1D*]G+#[4 
@)1.4'B:.!T] /Q[A"YU/PM;4-\PMI6WC&RF*FH%9\D  
@/)8'\[T4LNT3ES",NP+_*0V6[.XWPUP@9Z=,\89)H-@ 
@S)H6NWI9]4=7CY^$+/"_M&W:,H*92<N6;\!9TO)-;V0 
@Z;0]['HO2-[53VFCLPIMI(K?!''L[MS:8A<\%S&7)@0 
@.?RO+^8NC&=R:&) +-613IW>)H#(L8_8>$$?W2,%S$( 
@FO&HE:L(KK:J^AFUA84S WXY1_/;J*P24J\"PB\(L3P 
@)+99G5K1F"8@TB:D=^9K"IL=*1/?GOP'4[MK0P;_E3@ 
@;KD!2>^,S;\?-VT4WP[GS4%Z#\L"LI*^?[_HA2J^)/L 
@4W$5 8OM?U*38E7=A@G>2*3_I%8"G<K@7QXU>T0[O5< 
@_\&8]:VT@NB"HW#V]'[2ZF[&^&K!_>9JQXU/2SGT)X  
@*]$+3SQ^DV=KPD(TBFI\G3)89D?**OI5*6@3;;_#:N4 
@I>4,9W -X)T))B2S7%)*F#@)EUN%OC>*5?]4" ]G/SD 
@!VH9AW^^-EBCKR9&6["UUOEGDW@#!MER[)VVVYQ-. @ 
@:SEU^?QGI'&U!L[-Y8.Q^]7VWIT1L[RX0G<J]&40$$P 
@ %%1-&+Z3+(WJSM6DT5M8[)H @?4;7H*(D%,5B7=9%  
@QVK "@Q?Z6'DO[BWN.MOI/%97^-%B ,+"ENW!A(/2RH 
@.K0;&:7VC_;(_O1'FIKRG'VH&KJ9#SS1A3#]#EG9BDH 
@K#M@A.Z/?SQ22:L7)1IQSVF42$*T_&%X$I:IQ9\9K80 
@1>27%:SDI75*M+/VBQB9OW0D2$[@Q=+DQ6G5YP6;U$< 
@>[>([0RS4J\H;&-LR2CDC?RXC=>)3(PXRC88TM$Q$\  
@U2;]+;_^4F@/B 0#6HR*MFO/*USB0E!\3HL-^J@AL=H 
@*J5\\YQE3\&L0,;IH'WT8;^X]I/WK$\GN)G);CB(U>$ 
@ZS?X>PK[HPBQ5'6H;T(!MS5*(OUC_Y29*WBQD6Y>K*( 
@T85WMJM3H-EP\Y_TL0Y6]2,)+G.&J_=>+7/:*N\4##H 
@60VI:R=&HB1!XFQS]N7X.V+[Z#R*@<<^V=+E8QQ)GF  
@)%#.#R6?/<P[-WW"N17O/3+D>"+7##F+?1-:87]K45X 
@2'C@4@6X;F1 +09)G E[[Z$CSN>)+3<3S,&F%'QETR4 
@X0;)MM?]B_O"#F_RJ=9ZGT5YAI)DZ:0S<L'.('W5ITL 
@SA_G5;4B3OWIB;<9M=C&IL>*#D^DRW(0IR,<Q77XN40 
@=0\>NT8*7N9O7L#1_9V3N"G^+D>1&)\8 _ZF&(W6V1@ 
@R'0O_F)_O,R][N=XJ%\E H8GD#_MN$P)FQ7EE=RATT\ 
@E<'NKT+( M>1-JJDP\6&[.;=L#,4/,J/]668^K<O+ZX 
@2M*PN40_8]0[O^8OL&[3K?=>D[>P&G0X!H.B8M8]J>D 
@%',<#FSE\F'=F 9E)N3$FE75@:5 A@@UF4:DE=."1@D 
@"0/0Y'*JB[%LA;.WF-!)K@E%SY16'!S0DOM<I:3%[G$ 
@6S5+M/]!I8,PX"80W]8;Y2<=ID"L'G)G]Z5)_VZ7M+L 
@]!'[7B4M$AYQ,%!&!N3'-)HJHGZ9!.(-NQ7+*3>+<(  
@DB ]L9 \/NECGB& V:6S[[E_D?Y^K+36$\:A<,0!22X 
@*U^SUJ3$U%"B5]=E420L9*\6#5I/PC=".< MNE?WB6X 
@3:H[UC#$.E9M:L#]V^ Q>_C41M PJ#[:J?1KY,A;QUT 
@J0UA2/8J^ZPS9KVT[%-1@PU1S7&R 5^6Z_W:34.7JAL 
@I/:G]VXF51HON*SV?!E))$EC>]1:HH,!'E"50B*(!'8 
@M#Q08B39EBS(BN;@5;%V<7S?4>1W^&?P[O^X(B4]:_@ 
@?GLN@"M- (2(0='+>2DHL3NUSL<B6:34^-57BG9;Y2T 
@IA"AP@E"#%T6 VF:-N-8=YVCQV2B;]6<''=10<9<!KD 
@C5VM(850;A<]<S1]2=G)EI7"JQ+.'X-/!F8(D&M[150 
@Z*[_D/^\IS#MI&'A*X+HJ/ UQSNBH$&BV]5EPPEQ1LD 
@BZ5)#!;QJ9+\=\H1P>IGCG-,TS7HRX#0R#EM<Q^3:=, 
@%=G;I*VR 7:CM&")#7Z#>\(3Y.(O% ^?L%%A" @\(AX 
@I.KV4,W"/P+:93[K-2'*,]8Y3.)LJZDX^5E#LAH ^U4 
@^)U-L1G=A7ZL42Z&>AAO?JB/B+PST5+YTB)W65^/L,L 
@FN1!:C>XA/<X5L!;D=6.K48$VA[93M6W QNYQ9MP<VD 
@75S\O,M9W;$']")D!D/,\5PJ;__!6U!1E4J0,\ZCD:X 
@D9V+>I7005^Y<J,K\[)&W%[SAHJ\/[@/];PV,IZ4-)8 
@7NA3EHA2 _L8=6!Z&)BV-RX*#1U#/,@-Y<@4_]F<F?X 
@,P>",SQU%M\D)44 L+#.,9_&'&MG S !U4^ZWE3]R   
@ZU4[9I" :!)L&TA/Y,Z _U)^)(C)KMH*G4AP ,:"8S@ 
@OW>I(RS3+$2(13T0G+7!]C^$H>S'5P?<27O$+R1IU6H 
@C8]#C/T9:[P/B/"B:$-9]R )2#O$(5N"Z#3#MTZDN]@ 
@44?IZ8\6AG&+TYU.Q0&#BUB8)7^=MV5%VS8GZ3S;+], 
@J>V=EIN4>^0M';ZBH-S9"O7MM/'+JT.?O ^71SVV?CL 
@A3/5>(?(=/5?Q83M@I$_.5TXW[:HX&$.2--],OWVPOL 
@HD1D?D]U$L*6]4Y//Q;Y2$\NEX37A+):TFQ6C=F@='$ 
@C%/R*1J8Y3_O@8MZ>T\2TLARLMZ7MQ5+\^. OA;>9Y@ 
@Q?W2U$M[*PF*"Z[QG76=_]54GM(L9Y:+_;_'!'VW5R, 
@KN&/!F?1HR@X?OXU^I2X"1[G**?I-<I=<F+I5(E'D"$ 
@9<3*2124_.-#4D6/66>!@X^*>XMY-58^0O!!\C@U<\T 
@'_,*^_ 3D??/Y"3AV>M)'+V$_!T]FQ;4%0,-/3C!M]@ 
@S5TYWA4>\ESIO?8D3333V7),[_K A?>&X0D*)>\"-B0 
@3&W$C=[AGYZ[*D-L Z/BF61=8K_40[,E2S&;G%]K9C< 
@!V0Y=])\ZS)N"2-ARYB_L'38Y3ZC4H6U_%CIMGJANR8 
@?:]Q?L U_3<:W&(0681+BR_'W^]WN%TB$>(\LJHFRVH 
@:$TN=B:2&>?_#FAB =24_3+8SFPF83GV*UL\Y+XR'LH 
@-8 FHZ$(NE!G; I,B.;J"?5E0R_7%+L?--NFH7IY?F, 
@E\BK+!2VVQ3\V:)WB"2^X;YD0,<;0+R^*+=Y\,I1W=0 
@^"H=H;(,_VW4J7\*\?,2-B[,&J&2=O#=OXA*JTA1X!T 
@ON[:SJMTR1"Y++H7]^F9MIJ)8<#Z7R>AO[1LPJ>9,M8 
@+$E1HH89$1^!F=^][0[!>@M%PV^HPG<VY@IBI ]EM^T 
@="W&W/'8AR&^'TAM]DR"<WK>?:P-GU\*F"*OJ)-%AU\ 
@AI%)[73C=+SI5B;()Z%D$QTRP.:=7D49SY5'EN"PT@T 
@QOBU-II8^O]='>'8D!.3EAV,X3_GES%<,]E2Y$&9M<\ 
@.?K2.)##R9Q\G9^S%NQF%+..:HA&)/ O0C"GA)<NVST 
@\T"PC&X=ZV36N,^5K:@J-FOM!#7H?'QR,+/1Q5+*,B  
@DX>FE4^@9,O"XVCD.MT]KRM7J^T$'QEE$\8&!413MK@ 
@&T&G_/JAN]Z+3:7QGLPC7USGV_!""WFZH/W7+Y?3M@P 
@2?O%0]2_>RRD?",9K=0"WI?%WSE#ZCV_!P7E)+YI(;D 
@.E66;VR5%5PYE_/.O'Y70+<J#9P9!=?_'R--@W;);.\ 
@-Q&1'1:E9$AN3W,!C6^H@"JO%MRLLW[7])4F!(\O4ED 
@F^EMD#WYXNT^YV=G$A!Q3L%VM .XC?B+QN#,FK+'A%X 
@SYG'LQ J'(2\-,ED<QO-HY@0CS"[FW,='$.%^V1S&(T 
@MR93FO;%E"#-]N,9DAQ!-]_IO/&^F<&^_C,J)Z7):>< 
@EXG[%9/61'3U(C!'"NFT][">APZ"#AO32[\ODENA-)X 
@P:$>V)C8O]>L;=&<'V?5"A9 &3]S5Z' N?4>#]DNA+  
@__N7<LT+(WU]Y2!-Y:<#N<(:0'2P)V .-O<3XV2)G[0 
@@-E#<ML^]YREEB3[=.ZRYN8S"R7=)K4 LG5G)QL)\%, 
@$CFV"IFG10T'VKV!"%MJDPH"!S,^-U1+J +INNOXTW, 
@E2J[%IIM*]L-*NF,^,!:W7#1>/5L!O7^BB'5 C %I,4 
@4Q)4[W-/_2BC;;LHG@TLY'Y=@@IA.HDN 1CSU_$FY%8 
@"P/"08U_UF><S;2EU5F>A<FZ\])(KIR_6&WRE689+:P 
@/8K73%/G!%2-/J8_8]@FV8R,,GN2^HUZ:I*'Y'YPBJ8 
@T/)FWHY*FD'@'QHT&/' UN9.U#XF+9Z,U1QC4=B#>M@ 
@66J8!W5(YZ8]D2D5:!1%PA 3X[0Z2C:A2DK%:Q[F3#P 
@YLN4<1K:;X@ZR+)4C7JWTE9LQ^08GI&S5%\, =PA;HX 
@N-*:K!<208Z>N+(;F>*Z?I_G>VSG9"[Y=P4RR9Z<2]0 
@""=$,1&E+I *'3-',I!$%<[\.([CZ,_M>Y!Q2YG=8W( 
@Z%#7[E#QA+H!$C?8.%M&6J7RQM^1,LFL^7X<1<VC[A8 
@<37;7.N6O/>/E\ 6_V%X)-+KUB+Q;[#K9G.J>8XY<[P 
@O2=SKF!\[-FD7N..0!82RRZ-\XGFP?2\$=FW<-ROM0@ 
@N!K6'%TJ:-M$C@F.;CZ#K-U4:L02^FK)-T1CRK=DQ)D 
@ =I1X&[$?2(@,M3T"(MB5K>S38'=70]\(#?%%9EB*YL 
@%P-H6$1Z:KB/4OOM$<LM'SG8"0BXJ=_+&FQ7DWS0\8\ 
@7%7!=F62T#Q5L,3P7#X;1.HZR4S8FI.!__(&PS4)AKH 
@0/JH);<)$"J_;HU)C"4_/#RLK(6"3 9WEDU;NU8>*/< 
@"\399K"%L;FBT*Q9)DP+;J2O"9MX3TO;E5([^2,2O20 
@N5RK3+_L#?![0,S2:@1+OAG&X>ATCN.1;*EXLMD<GFD 
@)1P5QOUR[_^\M&TY$6PYU3]]-_0@T B8R)^C:*;3/OX 
@>F,0O>T?'8'%PYR1.IL6!6O&=6?HM 3Z+DG<J4.@'W$ 
@J5D#;#>,!*H4.KX.B>%K'2=>#K=FC;VI[VLM,&N,_SL 
@,[4O])( Q?O/:9:#-9LI42K;%T!I2Y * M'SJ9@DY0\ 
@J3#0>3R".^5DY>.SV_M'P<'J+)&/7OXRF7!+__&*,P4 
@K1M6DU(CQ2$>\NOAN4X09%:J_A/8XE) Y3RMMN&#2F4 
@\FL&I#V%"*3_G_;FQ&FXH E6SWTEB-;G:HP0%74,4KL 
@<R)P,$%%P!<-CRJ02:D_,JJ^_"ZQP.A^)!^W_RE!4S0 
@$FGNAK.@NJA[EV_)QJ??+%^Y 5"W?L&\N3)IP9U'# L 
@(';5I:49?TK(,C45?0R'=Z_1"#1-2B-8B Q*6II./;T 
@#T!(PM@=":06?X#55PA^IG)POD8OF6:_16$[]!*Q9/@ 
@1NY>+4AJ)*B?4YRA!)B@^J WGAWU%4]ZW9@#YV0SL.D 
@3.B:&?$#&44Q?LQ!2%*JF'< .7E^X@8>*H;&C L0.H, 
@5I:HHW6KN"<)&T+%[YF-)?C'2]6/MN5UCY4S=XP'7+< 
@X=S)CY>V,]IW4(+4E =1/2J-N5GU]B$-R-4"T# (?\4 
@87MZK,UIFU6/CTMHB^4_@13(++EVEJ%)KF;\C^.GJ,$ 
@^(F\T^,/PL(LSI%G=)3OK#AJ]B[/PAX:P0;[!VO,KJP 
@ _S-'*CI^31??Y=Z*:7*6[S/7VX:"TB\%@?5S@-H4*D 
@L'DPR20%;>(0RB%QJ0;>QUI2QF;?7"^ RR+4]6@/G,$ 
@"26U5@(_6W_%'7 :?CBX;-AX<@F!(']F9U^@NH"^J   
@8@>86;0)@!5!="+& Q--B(/]1K?7UVQ*S&#4@'AA^\L 
@N!0W7FO=(AC-I@KTL@WC!YKTT=NHOC@,'%A0$:M1T^( 
@*PE86B!)B@D>YV21E\\V3I]LYO/L^!\1ZCE_.##:2<0 
@\T4ZVY_-@'8\,PGE^V32_T^\",!-'6G]LL=3_OQHH^L 
@#DOMC]=JV==-RLAI$S-?4]6D(>J08+U,828@F(S-8OX 
@9 N$..1(6J9F^+'502=?;V8EI\:( ;V\]7/D>0UJA#T 
@Z&9#--R+[XD-C'FSL/>,IKY+7I/R,&F#Q%2VLM-ANHD 
@=L*,4HS,HQ %E0(.L!;.H^Z(@C].G7JJSV+;C/1"F^4 
@.?_R=R-'YA?.S3[^LKC,'MEAV[[&[&E"OE8ECMRG#1( 
@"\0\/PUD[; $E:YLT.30X.E([I=;M3GWJQ9*DL$'?[8 
@P<[EL]0K]O)(%&[GSWG86,.]PY[[YVS\@:%X:DF #(  
@$IS(,:"8Y,X&2_JUJ"ICK;1'F!SP7;!/N EYO,:3,08 
@YN*/_@I^6E?9\ ,1U]"JO& $T=<X&MHB*0.=]+!=;\\ 
@%"1N%6P6N\HLJ/&L OP/4FKUJB6B;*\CH1HUHG\@R@< 
@'=*+?V@Z2+/G18GRM6<IM*?T_?7^9RU<.:D/YM]35TD 
@9X(^U7I[=_5"#-8',JJFD)>!<[?%K@JC44ZKN[>=(B0 
@E2:F<G!&5PEIV5N#3@*U[FYQ=N"SX#D%B3)G_?6".'@ 
@2*(T7%@Y^)Z<!Z1?<<RA>@R='9\GZQ.9KN9'&N=I)<8 
@1]YQSBFCH'[;Y$.<TF]X_J%BQ2]IIPENO1:KE8/,_8X 
@X9)]P'!S*1T4__T-/*MHM9.I.O;% 2MG!@(9<6X24#@ 
@ O<R'ILX)[J>7 O="18T41)O$Z*?[\]Y5-(<ARR6?CP 
@)G1M"J33FY_!JL'F1I6M.?Y@Y-)&J'D_?8Y>?OGDS0T 
@ *1YE*<S;EQ5W;_P@5ZD Y(Q5$$;;?B4,V77\0@GCF\ 
@+&EB<\R",5N+;GW]3X^/CK'GQ^A$Z5:21T23.!J7R[8 
@285I$?T&< !Z;?QFY,M-3]!BBN_-;Z]SXK=9/RU&GD@ 
@W*$FT92!<']H=%KZ@?\S<G"0+ON@XFM.@*4!O/ONF>0 
@4R,.1?G7Q#UH$=<#@4&?ZS'QTDI0JU+(29AL+/H%'E@ 
@\*E(VD5#Z=1T2!?_FZ2*I=NBVXX.HR<IS^SU!C@RH9< 
@^KA2Y,999A[:=JF#E&=!)7_F@7C7H8H%%M/J*=NWN\D 
@UAH&;'2D-CBV%X!6V^"[R'6F:%(5,;%&CX]_KM,QFFL 
@\PX=EL0I<(=/"Q[B>D9GRA,(._^ TJU> V7DI %.[>T 
@^1$_,$?;:#3T9E3>U$R_?5COC*]$A:_!\?'A;E55S+4 
@P"F'GP&)H7*9,;N!<H)%C,Y.5U@''Q"F:OH=A67.>), 
@#LS0?*E2P!U\B.(@]Z/;R2+DR;#M,&D'OD4S)\16!:, 
@U50 8Y?[1;QKWE73UHX7S F;&3(R!1W9/&<>@_Z5\!P 
@$;1?Z'?QPY"Y7!_)^<80F>D6XL9 8Z-:A65DOIF!2(8 
@3RX6[R O+2K*9'0A[<-Q+8D:'FPC"?-OZI0[ QT7^N8 
@H%UW7 Z$C8J[RNG-XW9JP%9E!F6(@E\N'EO3-#]=E7( 
@8^W[,+NDRZ7?.LM>_-LT^DK]JS\6K;U,%T3GMQ5QAG@ 
@MQ *I"K(;*2C3)AQV\]8;*B>%7:CNQ!A1-M84C5?&*( 
@!=3S) +]IP=FLQ.K<@N?)T"[?9=P\K9O1J?\3H,BV7D 
@,1R*&B/;_+6\T)-R-JTJ*3[TG.<[L^L.M^@IKOO3&\( 
@M-,3Q-&4 RG/QP8SY&13JROL1>VZ;9!(J]#3%*-9T*\ 
@^3N#FX(UW]"B_WZY K01V>(F.S1*%'5COROY'UQ4 7H 
@CVAW(;Y+MT6R=!>08J$;EO)&'XOY9/<&X *?:[,Z=.D 
@Z[^R*<7 $*(%A70,$]_3/UAD&B%P-0KLEP3?D$ C784 
@QLYTJ$<PK"VC25G=T+TA D=+I);\J?8HQ3H:48.4>S8 
@^@U]1E.WXUH,#,+*Z.45(>/(XZ0#)VL$%VN,LS[R(/< 
@BHERH*L^.TV>A#=R2YLFL;_GFYA=5G/QBNXM*>![6+T 
@H-NK3,/%#<R\,2HGLQU"_LK!K?*<LL=KQR)]4,:<T_T 
@\X<.MAS\-9R3X$-I037 ;H8$'LC&=@):5$+4@([.%Z0 
@1L0RQ+E7R %I/X8:/AHXU75=<FB"OY F_@^%FO\OC@H 
@ORY=Z*CFA1\NVA8?V59=V0J='4AP/II+/GN=ZXR]K_  
@)I-N-@!:A1M_DG4G>WW*7XU+BOCJ"EA.1I1W/06)Y4D 
@%PL(\0G*JC%G!.I'NHGC2+!EJ2V/+LC?NA/85HYT[^H 
@=R*,.$J^!LY/E%2ELY<K.W\C?9S[2HJJ@A5\MTU[/*4 
@9T%@@E^LF8#%/M4)E;2R@U97P7IX-F68QK2]T1Z1Z4\ 
@%/5,]@O>]7;&J6"1*F [2OQ&5\:!6+0U0BJ<Y74P.T, 
@#F\P^5^XZ4!S;]%KGP3?B#J AR\ C_+-,Z=*<V2 ;FP 
@0UI-29,57E2X%)&+&/O$XG_W'8RAMKR0WBQU"[*W4QH 
@$&-\O$W#S6<.K4OS6CN@2@^8%<C/+#KY+KX?DOQU2A$ 
@D>&9E&OWH7;_<!N3JXA!#7E-2J%<#&[7FXQ3<<3J;UH 
@[]$S\JY"1KUU202D78@]"?V2Q'"O9%/''!R2A:2,FXD 
@Y5=[VI5E@$1,E/$^ .=7(8(3;?$*+=ROXS/6N&"[JF  
@,VU*CR;@79S>KQ#OO27 Y4 #5:V!VY5QPMBBV//YHTL 
@VB?0,.P31Y21'UF0RZ8\W"9+E)"%C]C??8=NP1<_?LH 
@?W;^:%K0K24,*=DNW.#K>Y%A3H@%^CMKAM#A(,W7!6  
@CT%QM EI:4?,1$]M[ 3R5*>.E->?VBI(Y^NBM]5%FB\ 
@08_[!L.BD<$,>?E\XZR\PBLEI%-?] 2<\'YNBI U#_$ 
@?O;I0P6AI63C%M9SJSUS70Y3D]N"+#)BSM]PX5,";"P 
@BY26UW>CX1Y6I;ZZRWHV4%[K!LG<6C&RZ'4@'.]4_[L 
@D:A)F"&4]<"$-O8F:O,O.GGG_MP1UR>=;S(_@$M,6Y  
@;=#\W5)M[X'[.Q88((@FKO\#[H)[',!I9UM>3!]%M/@ 
@/X&I<E/GBUL;@,U8,IDW)J4H'9[.!/@!'&7]247\KHT 
@QD!&[.DREZFTP[5\I[!;"8S[MDY3@U =W!?K%N$F'<$ 
@Y4Q)F]LG*+",.P]-OGKRZ+N+8H\O#Y4C%=16;@UJ*B0 
@-6FBX2E5%J: P]O@&:V RB]88FF_4&P.?QL%*$C7*1T 
@%[&!0FQ&0@M;92G@0323@U^$XZN?R511]]WD%<OFW&$ 
@8Y8IFJAOVK-L%QNX2J85]&9*C]LQFL(+V$/3G.U Z,< 
@:P[-J.+UTHA7IZ<[@M)=:P9<+D5CBL=0]]ZX"#^;/&L 
@Q;^N'Y'PQ]C6_VI6RH>7W-5P+/I\DOAN&K(H,12.DWX 
@A<]SR3@6K6MJV+/Z[)X0K57<.OI573X90N?.B\M!'!, 
@Q3!&KJNB&F9P)E^HJ?1C;Q]*<0K!<)WPT RRIH9"A%L 
@N^W-C:_5C>J_R%>M6PM)3ULMF%PNDD5H2#DITC1O.7  
@ZS#FV1;C09[_[K&WU4]C6E)Z4K=8>.CS$7/#4$(D;"$ 
@,%\9,'F!'M?S!;7SRENXRWB3GO>_4N7E#W1/\[:BKNH 
@AN=S]AM-^F>I#EG'YE V\=9<BO+V0],XTT31K*(P&+\ 
@EF  ;'1M2=\%S#:T@&I[RTCO?7C6OPY/QCX2#5D5@[P 
@5]D11@)]T&8'-^)H([26+[.>_YZN3FDEWR:M8HM>1Y< 
@Y<8!T*(>P7 .PAP40Q;/[*#X4Y(>RSN_RR;^9MG_HF0 
@6JXF!]?A!' <R,?":&77Z2+ERK%#S@Q*13/F)))U'*L 
@89/#;/<[SB.:G1W.3C_LS$__R2GG-X6>4YW8D$\_NWT 
@,R#>O0Y[=>P]J.6J:C"X&0A?#)8IPQ=Q4(15%33SMZL 
@YMO01N"GU5<!AQE1Q$]>F&H\ZM'0.C?VVHNG31*:J&\ 
@D,R^F%X>6DI=X+=0'KDF\V#5:"@8,%9<\ZN<R5=,#N< 
@K16^#1/G0L4X1^@%.7(V<%-<?4SE^@]H^6.L !)/5<@ 
@ME%6TI88E$P SM^A36U;EFW)$/*.IEK73=(@Z)#;M&H 
@:("8.PQ(WS)7I(+"+&'JZ+TI34&1D)E*=I6T*;0S(H0 
@MJ%\'8[F'+5?IW\.'\WJ9A16AEJ==8[B<M"LLW6#)X\ 
@:&'A:8&SHO_J7OBAG,:2XLV6(J5QGVC2LF\OG23-$^8 
@*&%H0TH4Q5VNR)GSG-"CDGP_!!A%3.6GG5F*CMNOI,4 
@L'!PNN+;9%1"SQBOOQ9M?:YXS*&-Y+BJ8;E>?5LO#HH 
@R12@.+#Y/+GK'?%X3<M$XH%XL(#H&M^\7PDBJG\.!]D 
@4(F)=]E[0K$FK&8[.LO+#M,1#67A,]SB& "R@;.Z_%( 
@?58VKM7>%_MX;"-!/WA.;XMVB2KY5V[/OXX7$4TV$R0 
0HKF;J('MOU-J6;$$@*=._   
0S^RC%_/]+K2RMLZ?H8:ISP  
`pragma protect end_protected
