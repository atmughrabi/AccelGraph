// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PYw2U0ls0kw04Cn2KA5K7uM3xXRuO2KNkQeER+D28l0UUcfmXDfJfj47DTBSRQP/
KLR8mwgh5kQwVbVOWMtIMnLqsCTWm4AtHWCmb6mJC5DVM6oPHPJwG/1hzdpYdX3b
b6X1DdcNl9mR2EEeCrwa7p9ZomFs06Rp4YeAxTA4xEI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42752)
tIO4KGwQTUk4hrhp+f1xmNCFZoL/v74v8c7YqkrBRdAoeAPQERWQXQFUL89VJY94
1jJTEjWf+v/ezMBQYNRPPmsC5PbzMexUAW/cS/xSrpG/o2Xzoq6s3DZ3fOhEQwXs
4HuqbKH+N65QR45F+2UzOv9ZKpWTnST3rMNWaZis99EserPw7HzYBK/VOYB9zqks
xPdFMkzQ1E/Z1KvA/Z3KAKn2mAvfFV23zy9FS9eyqDlK0UbzLt/EAr7IZx99PNL8
mSd58sNwR+PAD9+6aezLHM0NV+/2fiCLm0a3KzPNb1M13bgRQzch3/UjDrhTrRAe
kP4HcRM4qeu+V7xxXXzZ0Ej0BiuVtJWHN3LfS4UsdvHM3jS2FLFSGst756ks7cLZ
qlZ0VscqBvuHxI8nRdbZ2oK0YiQqvLx/wUAMaPJX5vPHX4rqvHUSp3Vi6P3j0b6j
xDx16P5vAaddSHwJuPXqVLcMYbSTJHerCDUFTfjmMSEoT5e0Yd8KZHwkDWSmTdDg
l+lRa8ylZNYPB3wLi9Kp9J7FJ1rI41YIOYd1B9zRFIeNikKaAT3AlCNsuTbdAkFk
JJA8HN29Sf++UqcAWHf3KG60Ivz7Jj05MuorwMTj7U6Ma4JoLoSYrfsmJL8CLmoY
zA1LXcnaPhk7ofIL5Q0P5UbJ4bSLGFDNH0taJPkxjWlRWHh/3YJXmCg0lY6b+wwb
mXkR1MqFZhCLCEYK2p54ucyosFLfZOYqA77k6kjvojjeOmLHOKEJ7GFW9d6PrWTy
1hELELHyo74H1ipzYyLXCdEJyhKOnFxn5QufqKglu79oUu/g3CcYfZn4dwJamlm7
qb6nr2vMn8WB87Gt0nwt4HdgJdjlv/+bey/HCcVA9KfD26Qmy1ywwL2K0UZZDe7k
Idfzo9ThSFyfSTGEqURNp8B9l/29eY/eoPKCjEyi+3SR5FRbHNN8AZczYb6HyFXb
ng9srpkevV6gIEJ5XovyrnhwV12ue4L0/ZIL/iC9mCgBZD+MPr7Qfsln9XUbL/JB
TIVPZm6K7v0hRF2QQN4MH4p/wgE1HN3iULHjU1q4WPKLPdHNRR90g32A2P+Qt8hZ
uUoyaq0Jl8BoMaai4kIhfrpJsssqryufgI8PCQU2bizNpSnZYRBivSfRIfZuQlWS
VJiO0P/l95P9LbKwjnjoHGWVNL+ocHT4m0FIG4UMGhcjsBVxd2vW5UHv+jwaSyaY
lKH1aVqEYvZooS5zNi3u2Q2fMNXkBVe+C5jZcjT5KxWDwPDDzhyj1zKfuPJMDoss
lR7+xijuknC8LqqFy4kqUId1yr9oQu9zBYvGg2lkiRsWX/nTlQWt5Vz91MoS8Meo
90I5z3usGzmQnJSGYU8rqfsJRdGtj8OVUM5+6oGjrGEMDrdZUZHYIhsnXT9DpAei
If9zqrlSnEKRuel7kNIeUf+yDrJjBkqhvRKqUgS3RYPmCCt4vwSa4dW19oJZmhqU
RzWrDUpeStuC124A7oLWiO0cZzToWLPW/GkY3ckB/gRbOdUf948ff+iZ7s3ijl6Y
z1kphCXErjWc0akvIY5h+bVrwBND+1l0Z6TyTC+YuVuoA9ThAyqD3mx46g4jsc9Y
vP1QEJub8imhQUQ3eBkr0EFTab5h2x9vDTY9kExDj6TpptAKFnNglx7Pt4O7OEEL
mRf2s6LoclQPn51z+tkrt910AvYKWWbxJ7QznzwPzzVfgdgX8a99u/LmxOPuvcwF
azG4wNMpJTazZDZYNB4Irz8gTk59549X0gy3mu6WoRmq2rQLnkmyAWtJZw2nNcXW
SGm/3j0iEsGGg0MsuD+J753QaE1SZbeJT+zjRPXosPVfPsLQPEn+8o/PsL5wSSQL
mBsKOapFVbWu3nVj8bwy5mbAidpKVsrlcw04EVTYh9A+MF19Cx/WR8TqQe5Q16Ob
z7ISM716s7HKgfVB3uh93IgwvIX47tQ5+OlszLxjyFxmmbSHRG0HtQul4w4zMMTr
o8EuUZue5GUL4ToConJBtWszge1CJiBLJUaCGVmKn3BRg+7GnJ/el2HC4qIP5cHC
vZ4nonvyNBcakHafoSo0pS1wJkpL05aOomQcvT1KKbdv24Z5qARoMlMHt3LPBLkC
1PjWAGuD8tDN4pWsoVcP+BY0v/2T0VHk6wFQpYTfRQxBkuwoqBSlfRqQqrx77Eml
ihjfaVPRFxD2LE9Dz+vqglaZBB4EqIyWjEvdX5TzkMDYomwpFRWjuplDWjLntSjp
UsfCbgN700SbTO9vXwHwOuam3GLtcziQMANKBFp9ZegqU9hURaQ7bJeeatRgduOB
SgkyTKd5YpNs73IsH5LPezx4M4/1hTwg9XXr8NNs0hhPvpsydsvIJ9h9J4Zc+S9l
SHaqrptvg7MgBMPt4oGMyR1bESy0DHv6BbSRqXBJXx21lV8RjSjXRmqm5kBRnAQO
tiNtDiO9uHryomd/Dohw9xBSYGGlAoeS+NQE04tsaqWO/8jhp1XgOH9iHgcY55Qs
8Gze1Y7+Q1Y2g9IuqMZLLnMgsHcULD5GHVuTZ06VlHFQ8HVpRmsybxaKPQ10AGA3
nrowpegg0QGZKpBo5a/RcWfxUf1DqQSXVTqxnLd8ZMgTKwHPO/7JoYRZTkj0dGXn
4szZOReTn3LfORn21JR/iJ/tnoDXpmViiM/ozMP1yMANQpEz2wy76U08HUIZMu+S
yn9rVIlaUhJIlJfc/nqroQQ76e79rtdhS3vDj/WvTVDJvn3zg60QSqhalFyOP0IZ
w3t3JEZHhxx/vDP8hAGDXTyLXVGkokosDAJ3jnKGLOxQ+Gfc1tBbt6ZmyRT9J0J9
RIWj286YezebdCZ2t4qFlRQdAI3yxx2RYOHncI/09U5p0Xh8+36zp7oLopvhDbLg
IX5/+HDLgtsEPHj2oWZQSGgtXP7hBG4TyGG2hIKgOLZTD+CC1hTzmEjz7k8BDyju
MECLO/2j6SFwO2EjiK3qUDckzlCQfJe28IGC1sgO5P19s3gc5HUGnKFUr5OTzBBj
Amzvx+1qDuRYxbarLDuIA7ek9Ind9OtFA34GNJKZ2Azedmm5zsVxfe7JKDOrBCDb
d1GCVUjGqBpHvacMETPj8mwF64R13d9MmUsKjxXhMIHDtnEHsAhEa9wNFn22rzCb
7hH6QJ1Y6SAP5TVy41UEBtTYq6U5Eat/40OaIiP0ickEZmGQfqlZ5ITVUZg2Y3Iz
UWlSsozDFd2VSMnAHLV8qBiZ2RcyQf28UpjPlF/PUzdoE1/dF9mYHe8FX5qH4gSj
ZtAtJWvb9xPQgRgPlJ75mFcmXd+0bZPPFAac6lFMxssIeJJZJPZw5YzHFyJEXbhr
PqL4iAadDQEidk/ioq3ORaF6rfntFrO5Q2s2uQ1IGa7oAmIgjYx7YmJuVoVO09qZ
sKwDzwuwn8co1ve3vsEgVx3MZLuyhMuUyePqmF/QXfek8FbCfgo2FGuO9WnSKSQg
QIZmM1piJ/AEICJ9vqo79tv0R5/wgVXkm1fom6SL6VLFhcAwRAPqbggxY9vo1D44
zzG7Joxfktejzsr7n/JFGi0ESvqZlW1uAO00HwHUsb+ChxNMjZEL82cZvyOeanXK
+3WBCuGA5Iy7W6FHjvXgQX4YGjXfZBVCSLe8GWxo8x2AdzdPGUNAIU2ulumo6Vqz
/u6EkqKqt6Tbt4kWDPqRaxkyUL4BGppwcKnY884fZ0fED+qhxelFCi/Sn1yELf6o
NecfWQl3S2bSh59Xuwee6kSerlda2Ifw76G0UGMLA0OAK1fS6whdhbg7dCVWcmaP
NaicHs5SlOOw8uT2ORKWxeuRUJaAXF/5ZynhK/RwtrAlYSejH33nJo5aRNHWEMR1
23yqRCys2sb4FOphW4pklFx9BOZcZMqKIHnMQDMnQMyr4/VMeVlooJ+TVtkZ6NNK
yMYJmjUiVNBknlWOWcSwTbPXONut0WEfhMk+sonsmoTf+nEm6URgKZURESY4st/Y
NrVBZ40fsu27YEMEPn/yQLxUTjHbiZt+bQVkkNxzlv/7/a0f2i8IEggns+2y5kZ3
XGA0VywuXEFd+jpV+2/Uoa5PmNbtxrWjpFJcDCY3KSTPnqeXrsc/Qa47lbGQ38bJ
M9l51WQF7U3USnckhZaJ4BcKKsSgdx6ojBjZdCp6LJagr75KDcwN2LVW9MicTA/q
eKssJvEbTLQR3mS0rslsK2HwJNSOPa6O2Gr6Hph2o0xS05yqhVRikl6CbVzeplqE
XCLjKtmwR6LKhtQuCPGPjOfFrU96BgmN8RYBK82yTCeuXJujghrc0I8b38yAdBVB
OiQDsYQf7nzp4b5Sy9ZVQ29Wu2r2P1XXuO5EJo4EQCbJHqsCWke2HZT3LgcIG3l5
OYLuTMVakZeG5+PeaWwPoUp7M6CT8Q0dKIzNkXSfp9YPG0xNlF5JLrxCLcHJ2GCK
JGowLp4wibwawOZ3ay3Jkj6WTfRLMLMxNTtzxhiAEouu+GXmXOYy8QBmPPGh2MOD
GYlEUo7lxj/mVSaWiIKOKnU9gDSf0kjksfaxK+n2ner+OPl1Pwnr1n+HyNyu87N3
A/DN1ud3i96nwnnYx8tfNb+3SQdpbmHiFPRwK1KvwigOS4fMqpIykNX5k15zxhtL
RfhJ33yE6FFwnh3o84qBrENaC7+DmKGyKvBVCoT+lKlLhWRPHJ7oIWhXdWo5nHle
wqkLTOq4wxlTnyg17eRksyf/MLMASyJL984uUh608WhloIUVYfUeKf4kWYp/fSuh
tige2eu4CJrIs0RJnYDgqqP+IN4aHoP3rgYOLvUN949uc86mD4hlSOZreQ7n2Ooo
8/2+bNNpD3awD3QTjqZEzVg2NaFefzLjMtmHypzEwz74vyMEzVRTHIWP9mVmt61B
SwPf4hopOrB0h3k/Fin64oa/WaXISqqEwxeJXf/hX3TLzZBnQMOcWuHpaTE0/E0i
TmBv8ciEn/Bh9Fe1awhC853+nn/a1aGFbZkuYQ4n/sugzFbW2LfaK7H0yFpnIzxT
SAa8c5o+CcQu/a2YusDzwYbkGP0mk09MGYnDhXn+sjDcQfgyAbFOAkXsX7NA+jFh
x13UBWpZq+hgFcAbi9mymrd3PGFSlwyteuz2p1IdUvYeNcRQgpXoEv/WfHi/hyyK
A7YU9FhI7CmHO7KyUn+XhoMbSIKEI8f+Dhxwik7/t6m0oyrJ6pIolWdJ1ZnVjvcd
OYKvX5uR1Vy9C1FWtwgF/Uv4UQs0TJZks7mRWA8xx/wnx4FWmAQ1Ow3RlQTILMZx
w3OUgWAh0RTDvPDvhUc+MbwHkjS1JUvAeF19io3uKC+4y+p/hPySttzrexcHzt4I
0oMecJaqDrsnm8TsID4u3li8c3VfhAiIzWoxJydFfasyrtzjnMMzSqQSCOe6aj5p
Gt1nQiAXHmf0He2cVBTLfzxY1WvEMjmj2ILJc09+Lcdnoj5/9kVcPNKISiB/htq4
RIL/Ee9Hm71biMi6XAmEP//2+o/10zzhBODUlDzdwLs0yAhUUd4IVpltytp/bvnQ
nVDbLoHagZm1F6fRniFPHnXPbBat6XiLtEKvWbV1mqRpxGCkArGeW+AEjHSO/iTI
sedN9aIp+hr/jkpWmbs8wcXoJDrkly5o9aYX57YZBalaEyy1UiusMpAgB/Q90ffx
3XzhsHhOHI4mFN6QAHzhmizdIIZkyTCymo2CegxW5AP/XoOyhB63+S3ygiPOj2en
1BcFWnXFAF3ivmiAyAnamqZ989xaVVfg2PVF2jwxlYKQYnezY4kkN7TdkHOr8648
S9Uycgk+KfLZLmQZSv2AHAsSG19h7/WYPKr8g2LazRsIY8cGS1TTIfOjmQBqz6Vp
vYgIFqB/hdLSDDJ9OczqbJSBxv9lJygTI3cSUFDPaxUbbXIGJRjJ/ydinybPkNXk
xQUWSE5NfzyTwm1kxm+/JKxP+GyqxU5EdNuzi9Y+Jbjfd83O0AuYzb9DCn6g5KaF
r/QUbSEp/edoQpe87MSG063xWySrcCGkURlrLXdIJ8A/rCgH1B6ZdnomGCCgBfWa
V101lnx+yjjhbekBdoclFmFlGhIJDIFDyKeDYKSXnEhLkj8ebqD9ynzHZ2WCbjpj
XYxoQrMBcizpjjYohwVyAcjzRoojbnFgzPzjHUURsXtU9BUyubtYR8WPs6r7WmY1
gfzhPg7LRHV9kly3IqaoBvJtRZxy7ksFPmRahU4gYzmIYjyi1oys1iekCuo7+xDo
DeNwBNLlxAsJXDhf+WG1Ch7b42cI/JoDjO1t32SCCg1RGpRhPgS5PPXv+ZOro2/t
/Siccpl5OJibMO8s/vXjqGeTWG5efSlr7EhbyH/Dm9YzEA13ZW90vSkNb8BXCNtc
xMh+coZ3Ru3BB23fxX4SD4zhdUDTHDagHKEpFBXuQZTmAp+QBSRG2B/e+qGk7Uow
4uMx2FXTIHGYgxU6fnMWjhy2JheVTPjrvYLc0820rsr97I53Dq28AUNzVn9adnJ6
T/k5fsA5Dch4pFdrISByIAPxtxCyqGXCFGXEl9j7B4/Yr9aGaAh/mHS3i9JrAGwM
2CycwhOloXc18a1LkchT7KloUOIy+IImXiqY/d0RCRzMDlPA19gfTrVUMeVDpwV0
2zRHnoYh2WIX5FUpPX2bTdkULmqQz7j4wDhsPRWgyHbE+fAenm/rFHwAPcH+7CR9
l+7tsmNEKcIDTqUBCbv1MN2eWOgLWPVlBBAj1uvfGnLi0945R5A46UA0cUkM/swN
I2zQPti1RsPMzh4TuvunUUYEuOAnWBXG9/t5zeVaYftj6f/5H1KFT1juFFQWl6QA
DavI1CZ5X2kqkBL40jCToCHnJ0UBrNTNdosXmewaFnZaDpJ/9pPydbatd6XruKZU
mKmeryhEIEiQeRfju19P7izgd6/c2+4XikOAmS3wVN9fyVmUh+MPw+lsql8l0waq
Xfr6girgHK7toOpoMsJIhanziXxCYNwT/MRZ4o+0J5oHDla+gQr/aaSneHt2pwqV
TSRZoX2SlqwZYXoWjdl1ijXNZPkj8S4XPu8d/0MrbDl0bNu5NSRWayQLMLbhlob+
Uf7uO5O0z69LxWvqrlX8TR8C2ybzCyR+JeQ4Ee3fVaFfORpCvgPgWv1bIXp7gO2b
6ApYRnpyQU+s368UB842R1ZzDaeSgE2bU08li251oszv+ayx1tBMq0Wdn5Iedn06
9/DhBXZy7huzQ9g/tFt0WNZl8n5oHNjEEldESYear813uOAMjFA8WnrO30660tIC
sbudH2Ne6o1UAp4tXx1X38DaIJAXmLNLkIbPhEN2bzi2nAg0IvQz6F1b4HL3NRNH
eTEtkARoCV9bwQBWPbepJ2PxUW1zj+c6O7rdyJkqpUZ3pA11M2PON44hID+rAkxJ
Ee+8XUiJq+XLDeTZUi4sUVXO3tAL9wN0p6ERe0LS/9DzCZkly0xVVs5qSXpgrESa
jectzulzyC9B1QPlvUdNdxl1sYTk2GSbspo2XY3pFRvuHi4IrjP1wlf1TNCDinsU
f47Gqw8NFYa5qy7uJU/QNpTUApC5mwV1drciANheZkSOZ5FsFTj5JwEM+ZuRFPVJ
QYFVVFucth1Z8zgqY4euedWVxpWFAPjhFqGpuLtHR6t7IRyOSvMz2g3IeQCVtclg
wbaY/8QW23Kjye/nKRje6t4tKpcaZhF3McdAN8/3itnfx1F/vt9waO8TYEgWawZU
I3rgOBy5irXgxUFVi7XSNAwS/nC6OIV48W7HXiHxiUt0pwr2Er1XR5/RXD3c7/Qe
GESPb651gw4i36L2Df+4FEe6CdhMXiS1zMqLKR7IPLwZDlIJ2+C53GLQ+LRCEf/k
7x82IePttbNSLJOGDbVC83pVQt8Ah+twcbvpTHHwGCrJ2Wyg/PyvSWP0gOA8ou8o
hlAI6rh53AB81vw9vI2NyW5ZINGbK9TCrAnj62jXepdOEDM/a5evVAuatqnQQA3b
fjQaYKEBRFi5fSkcGh9mvHGimkBin4nPHTsaG+RZiPwnmi6Zt2+pCA+ncg4+uNyg
TifwdBxdPQbncBHMdSRyahF+jICKq2tvG3znWe7iEptigZMn2DcJFkikz+HH9cn4
kDg+QH3qGatcH0raUlWMukF/Afr7GaUqsNm5aUx9wO/j9DGSTB2HOgkdIf/nZMdZ
S/43AquExiB6M3VGIAsayK8Yl2mFeOqI7Nxpb6HpwUGfcJJDD6SjwAchH+kJA95h
kp0YjnFX9I3iotzKduUGbNhbticicHUZ/YM2C0Egcqi1TsDPa0oQqDp4TjZ2NS6X
Rzqul09WMHUzvIakldcEfPHkS1IZdf7rKV3X8oNMm4/TgkJtdgPtbE88K40vOh56
z1SjDjKhZsbNvK47+J14YCn79UqyI4++4ynU/X9Z64kehb9RojhbRf7FRL89aPHD
V9eLN2D+614egjblCslJx+oZZlpPYQWgtY32JgjvGr7hVirQSDvpVOFcES1h3f3f
mXMvHiRw4HNAmmGdUH6BMvJX+0YfAklQiD4+ZI6hn8iWxM9t3gI0j6Zw5ZvdlzSi
RcZmT1G+BEZSlSHT8B9GfcYg404vdGVWOJcmkIphevIw+NZZhPJqyu1hnXuv/JTX
qalrvAFww/l7P9aeEp5x3MHtcbIBDdAYYkbjDiOdmii2qH6wz7Kll7oA5YNedbux
Y+Vbqv/psv3nzWErTM2mY4TCiEiV10ROhhQoNJARzFDZN2oDc0Fnmfc+hDGGNCoG
bEFi4CIFe8WOgHgszeLK2FC2Csa6BzLxSLMkwAMj1N/wBL0IVyoyRpoDgZas1kS1
jshABBymdiK4fmi5nJubc7NrAXfijL/zAjoeB5JpY75W/yA04oiiVq7+cJojfzL/
S5mzLypuHuiqsMHnD5m0taUjVcmsBP5YygMlU0pyPYPBLcbLAx/DkCZdPtkq1ebW
//6ThYmZarubvBSLFXN7tbaXUk31A8amI5F2sfm4aKjyqanS3RJ1fGCAQzMBp4hZ
VOn01vy+8cLhOUp/WCQXIYheWOdXr+VRTXl/iXhtYLBE/sTcz8cXZiSdALeiS38v
zvem1FMMNEyDLAQh9gMitJM4VHAORUJvUqPFfVbe3zoLyXMFHt6OCppxGfscQ7ZH
q4pyQ2VWNoJpQu7OBS7Hags8KhhLwo/SyhdKEk9zD8IMXWMDJ1RDyM5QFXQzVUex
gcHPnzcrnUUX9apAVXGAp2dXxLu+W9VQ7yLRvpEeXuIaD8L25qWtirQk4HLOjqFf
+aA+J9NrlpxfFmFMlwudxWZCc8Wr4Zv4WqYoLviSokOYIKu+4hOMiXPkOjzREaxt
zv4hpdCWYZttzP07jTD8T/5UTx7asH3DbNcA2/1nRbWEZFQuMGcCFRj9Pn3zgxTh
zvMEM+D8XxTz3Y0RJ64+q4FWVbWCb+HAlfAHcAZFUvIZa3GGlkdx7fxMSc+KquQe
NJ+0t6OtkCiy/CD8E1Rdqwfso/VN0Wg3tUrhRk0M9xOiS5OvgyBdkUTT/6esNcbM
u24m/veZWrhvSN8J2OHocvNWmMnCDI21zN1CRIcUpVes+QkzBv1qMg8LIKlhzPVU
EqEfuyb7TcbEd0jZ5nzWcKag/ZzAhosmDf2SXLnzVZ4jOVu0gRzXL6tYh7muEpmB
XQ2XsuyzlzMw0BPrGIYndxI7YO+xwvA/tny4L7mIzNjmj/hLQoHNzi6maRQj82oA
+r+ZA9XMcubSqJWMWOoXYTcDsavckF/Ztdc+WcVHgPbjbRQ6swJ8YC257vRz54WL
UkglTzfxYnuku/3l1mBkOIYH80R5tx99FbQcx9x9aCEWim2NmXwHkcfMNd93pNZ3
0f6YuxjFUr+yXfp34Xv1dQEUXbjzt19V69Vn25XPDGV8BkaIfN1lheaFNs53j+EV
E+J3+JNlxW2jEree/4G/535t7Gzuq4XuLkb2L8+uyfWe3a6TJF6r9KivutF3eIC4
rs/yYSWHCK7N1yVQncWmTfLNldWd66UEDg8qAY8Tz9u7jcRMqE8YJueBMOGrs+0g
EHzzyqrwE/m8jqNXEX2JSdPRZKN9yfEsuv7KdpHVIDacdbKtchRq08h3iM8lCxvV
vCJyUjUAP6mK0Ltk1c15Vas7llLZQmVGJo1/cN2aW5off3paAwwOlRqf9lUzOBOC
61k4FhXDXBa/5TVFP7Itqh+rGcm/Bu6Hws1Bcif2ox2n8/eyo7g7/oglLG3eKey/
a/N6fPZ9etltAzeYQEL8Uat+O5yuHDc9MYwH5Tno5dJgo8nYx0a1Omjba89xNEg8
VSKSfv4hHyVB8aSRnMlHOfvsiHko5mfjVnlsFVoxiusnfjMOidpB0bZs2MoSFrLQ
CqnHVfphi9NA8Sjjs+OTQTfqNIXpfM72ZSs1BqUorVcnPRwHpJibf374pIxFePIx
zLje3Odc7zJyOQAOxCie/2NMZubzSxiP1gWcuTQ62jpFa06pGznO1cRP0uZkxxv8
6dNi7ivqbbJt9sWUGvMGzYZa0izj14Ci8yoGRdYMYfHpSQPtV+iik087rhviR1jI
Z4zt9kCBgDub2FufBizMwb6SezLj+OB0Qlx0yjiV83jnNVgnBln6gwnPgb1phJMn
PBRvKR7PMUzxNL8Ypv+nCzX81Sw+AQEejViB6KRu7/q6kdvL4VqyQBKFyfVQ9SOD
ht940LuPDG4FK2vvYEIon5lleKFySXiTJDG6ZvU3Hi2PBrH/0vr+CzvqHSqxR5/Z
Y5edViIjaT0pS3R3a5FA48S9IbwBXbAMmqFekRAALxjz6F4oi2cRXX7V2f1P37RV
rfYAwOCY/ZRPjIQS1CBNNQVbMkRSw8+HSJCcTxpp6k3nFhOIxBx0dZFbfLjF6YEJ
Ewe0ug1EmujtTNBMEwvmhX/OuBXxykt9VJvToFpT7Fi06xb/CH8gVQAZziir5i0a
OEPJN8RDPx+43gfjEWPmGy39jU6Ch4GC44vRlzuZsydz2N7cmvv5zL6+trDJdExL
9RTIOu850CFKs7DZ5m6Cd/ovXYWPSBDZejtkWvFIxFzvSgx6h35cw7bJD+QSO7pu
vihfhSwVWJq4xOCDrLaa/J2Z+LLfi9PaMlvVV1bowh7+oWgvzNkD2DqN/oAE5aIx
8sM0viDS9S22ZhSHEwY3I8YGgG05Vg4ZHTVGm9ErCscb2EJZx5rgd4843V2EM8NI
cYUyNJ9UvOYyNIGq58MdoBGwTfQPl9Wm1jhiEK+eAMH/cYCBL9CYsR+wZMWENsgn
29lmLMl0BPP5Rb1baJjISMHwqzO7nyNpH/k4Yn8EZNJFa0WVW/GtmciKW2gApDB2
kOzl6gr677obvNKBlNt/S9tyCHlHo0GsCeLmhI77aACA+R0t17v12ZywoYE1B0Df
5IWg/xYjz5814+Hk0y6w95n419vZFBqgXaB2z6QSHdtScFVI7LBfawti3C+kUks9
2B5UqDEzsfOtJzJauRIz7XHNTmaIoVPG3dxjqPd408MX+r1b45cL8K/4GKF1UZAJ
Ev18/ZBCJpMnkxz0NoVPLyBiAjnN1CwXfkUv9fApD9m+uJpYWBcxHArOE9rA/R6T
Yd3PFkYUt20EArqbVQ4fKR7HQlohlwnj5I2C9+3QoKHYcUnFeOg0wem1FnSS+E/7
FDeiEgJa7bEJG+wat5gR/PGbGNRQyzK9B0reKJ49JcImh0S3zDv2db2IOor32xoK
uSF9ntX0FKvBLkCKs4IfQJ1DyeZBqyG/xx1Xq7+lmkTphJHlbb7h75b3qd40j9tV
dVt832u23QwUK8osW26XQA1ttk7u5uR/kkksxxW+koc8PclbdJn9vFBZ6Vk6GaXp
maxxaV+zT1jdu8o7wOf39xVavIRXs57Px4zr47WwUHXvWwHZG2VlxqdHjpDXUOfj
+PL5v6BS2cu20/OYTCNzyLxIoylnal3OkpitrT1u2aU8mhiGCmNvBrb9ldUQfvdq
fYZlboRJIcDZ/0UslbNA2Cr4mf11bt7mymqB2kZjnY69yNgGCKirleuLbzYLnFjY
GdtaOjUCOgZWsFO1lgwy7OHpCZjlZfRPCojPl8g9L8sZQsrQyNEHZ72dlZ14r2yc
lOaGQ2YROD49obRu6NE21b/eDS869uoQ1l4tlbfxu/7z7A9Y9tJVqnsY75t0W1fD
A8GVYtWYvjVzIT+hJ2yrVU0ykwo2lZlRsiim3LymhE6YU/oluRDPLHaAOPx8gCs6
itOSJBIrMn43Bn9UIh1Uccl3Y1vUoC2EMjjRz7Zr20stnYqOIPXssrN9nVjGGHK1
aslldEDDXkLLgvKvW524fHI7XEfSgc8eclBEbTyk0GTNBAg4KEYtmL2saBmCgkIb
z8TzLB+S8qIPN79Hjm69yc8cwFVAGbCkN6TUCefsZs2DvG39yVM5pV1ayabBx/Q1
1u1IIoKpvIV7gpopA3Ta3djmNGLgyVYOQkSp42gAlzzuyhpFtGKlVmfBfVgnx9Vp
iUNrJ7T+mLF3WKvd2qO3HWYy/hlaCkWgJ1uIDR++6WSjFGIkXMOX8BDMbHNQOrD3
eJ5K9zWqYWSs0FAnTcuJV5t6f8d9+uM54+ncI6W1/GZwbTX08hSKttF+wRl7La6o
MEjRwdjTzfkD79cGDLEG8q1mzgT56zBXbBClE3bfrrWqo+Row5wqKNRRd+ipR7U4
BqPPUQklj9rAltgHZlAzxKrxf1fOfJFRP4mBwGCJPt2ty4wd30N97IZvcxb27chu
Pwf6qnY3vd3UTvwxu/yISRRI9RtnlEGeJSqUugB38qB7VtjS35j+CC7kFnVCEz7w
NbPxvmb5wjyCT7VTGcYMBWYt1VjCv6SpHhyu7MyK7mOmcjKTrN5PiC9Jt4ZQbQ+E
QglK9qc7LDT98dNApbmo/rwUbYU6MRT+4050+FDljY+cPy7E1HDvklJGWvTAiegV
BUhsILI0Bvy1ABpmxzzR66i6phlF7kmJJLCdhnTpv2+PhtcAoy2qdXq/IfLsHSAy
XpdR8e4Fdglv66Uqhhclgf1Ja0bowGNF3AmwpfmqL3mdaxNn5Gn2jvTTlYEGejss
NbFz7SCutWNF+DHHOT65OX5EEOhqyKTiwKNzrnWIHPdKclQ5Sq+zIuM4vnU6wRnl
fWYvG//kksNQ6dgCusOf7uNCcYgM9+k/QF3JNb51gwTO+P3M69ef4dC/bQcelxaA
JDo+tFw0a1NRYoRKzb1FNvagjHcXDdnJXgvlhgyGqpsb8xqm00bzbUoIu2enyiF+
E1ttxyjNzj4IAgPJCoTyIHyJAU1tK0Pa+SPLhhSzk1oyiZBwbeW+gM+g8emfjtFr
7iFBymTVX4tGZHgn2i8nGJv69qiE5oah5aZVqHrJMUhOKrt5CfIhAnniSWD6vyAh
LQwgv3WNbxFx6RFXtpyZT8wtt3MWy7aINe9V8NONBu/p0X3MAHRBI1P3qFhg81hG
gIrP1hl14LE3ffSwVDnvWi0ZlmiKksxsabkTdg8lL0UAwREO0PV8gN29SGtVVu+r
cb0tgr8KBEN3WhAK17LaSwK4a5P0IlwoCrlV25Dtg+lw05jz5EmVM7rW547PEvNf
eG53WUnhxJPaLYGBy3NR8YO+WCwt4oZX11QeOMHk1AoHfy6aXfHGagiVUhn694wr
SZOCrOUN2sc7B7Gvqe/6sTebcaue5U6KQAma2WiOeqx0gkQDxypz4S4IQQUfkLX7
1Dgc7UdUVkKYqk77+eliOH7wypfgLvX3UzRvC+rzkwycxWrQveBauZrtzOCl9r5Q
BsBnmKz4tLJQcT3mGnS0AyAG4VZfZBdTOotEZBT8MA+0+zMKm/640u4ZQ1wryKMo
vJ6RiIbA4XtfX+5D+8Td5M/2QS11U3NBkogmSP8RPgOCM3MzEIb86p/LTfdgZkG1
6jAUdFTXTbQiqzNdbUYRyaOcOqqCh+xci9RQKSQ97kUGpqMhhBX7kdU9XiQaEgH3
WaGquM27dbZKMyqWDartx0BzgzuVBNmGT9IZgM0KME08X9m6+0yNvCGhueS/MJUG
5Qx75qG5d/g/TNC4OYeQcBOR+NHogs0HhRHEV1TvtZTBWQstYD2wtlJHgUlTsoQJ
7ieNERAx0osQIp/5abDY3DrY8ZNzXn9pWLVpyRuN4RiItuVvZVnn4fRfjXgJMmaj
auRH2Kz7BJsYY+Yjq8EVNTVb7nWLft+4CKCIChq+/lulwDgtEw7W/otz0FTBT8Rm
FwkD9bvK7QOyDpt84lVYLTi8dmoXLEtqMeQX7b/1hoDlpCB9MVmeH3R1jmwlSUHo
HJiyzcSvGMmprkZRECc1LToXeQ+mK8Y9EEqDwtd6E6j40i2HvxBgQnovejRYgq9k
Vjbhmx62dJcc0RNd49gPiqt9Kpu06p+/ouXAGm5e8/eKwtfGw/Ll54KmD+sn6c4o
U+Kk7ccf1ppTjaUBdpDySzyVxSRYXMasYL9GYJxvth8XRnNoJn0ecmS0oIqKRqlC
8ad0+S7ZsnhgVVlCouzStGsDbYCXTCEL06i1jxQABdSYu+FI4yjMnTxbgQ8g791M
aClbwyb62kyVItEZ4KUB+pSgj3X10DHijvnysXq72UE0cU9b4mEu2OC6JPbzpFyG
hBirLzJArwyAXh6yK9pCN2MMJ5sS8DyCCCi3UC1J5cnbaDW20J/1tudS/4g98Gpr
dCjjFpFe5MC8hLFKmw6zjdIajNgVdbF/7gvaspegIjx+7RUkpwOujsaMe03BN0HR
/q1IiKZb5CZ8Y+6Iom72G0H5YVghNKKoJNaDgAWwwq8qaY97ijwYwbIlSN/B2oHH
nHBKxgWoG5YeZuxClQvDkJJzxZgHGT72MhWCe58etgsxKPnapQ9pjKzFiqWwPB4P
9v3STnzrc/ziNn+cNbksJ4nzJjdcDxDd0MDEWp/PrqQK2zY41MbiIyNw+LMh0j+s
7Sbtk3QBKT7ZHPUNBChkmzP+rkr6bZN5vEbtjbDc/+my6H6ffe9pBGwZ00Z4y/Uo
f48fqQYKtcZVbajIFJBhWRTH0/1dPCP21JO5xbA7Laydyc2fWIJUb22BOIJdLM56
VfQWWrmngr/f/hNRk46CanM9gx8Bgyk8pS5BufTldS4LucG0y01dXx4PHFtcAmpL
VaULZywfIF2h6k+N91MUiilnJjuFHkU+ZBP+PrkNkpOLbECzWdORceGIDuD8dqV3
jroyS1RwjUhzN+szN+9L38gfDd52E/1z4nxt4exbODOZ+rXtVQ9arKSmAobowTsy
qu082FIw1cYW3agUCDZYpdyfsVB0CuHE/R3fXNUbHueSrRQoWXUdUvtlhdA5E0SV
03PKlwNaYDKEgscMpr14vwnELltaYhcSeaM2lbTso4Nw5+o/nE74PvOcgDE6C+Uq
5eBntSlVQ6xoaDjwKHCjv4f6FRJJmWChZf/FqvwNecijVP1BH6eNJpNBaQa2pdq6
aZRMFMJugwR10Ejy5mn8x3hhyA/KkYrcIOfkF9UTro7BgVO0aNICrQGrVzAKe1zT
ULMmv5m+CW9Q3ewCDieB+cBY2DNR+sW4wYtabGgBJQVD4ZkzH62rA+pln6pmxKM0
1mmcMfMLOsj1DdRNCOPJKyBPv9CuoJ+NIqw4WEum0GQxZe8GjABpUZnP7y2mzwyf
uTLaX9LNASCxLnn4U4c6+AU/2PCFszJ67ymAikVOmVCEP15TiAtLi7cZD/29y+Uy
993lBZPEkX0YBSx4oIFYEiGGPWZpUOXPTpz9TnUB7iI3MdtvxR4waawY4p/E/Ii7
1UqgDHAnjuDw9X/M5c2AV9EAWQwgd6sAZj2yeEbigBGBKiqI/LBRtYlinxsAK0xd
Ih0l6rQPhZF6ZUQbFb6Mt/v4J4rNlhAKY+0o1M9e4JDNqbnT/q9+zwtvBNU0xCH2
MMTPmrGoIvhgeRvebQdUttXz8lRubMvOTRJZixi/nkh9ryvtnc6iu6dvvn9PAmI2
P3SY9i8s3Y/E6HJprl3/Hz4cAXsnBiHUY7QH0TNCQTvTLwSeFtZi4pA7LdsreXgo
Fg7rpca8ho2URd4OVwotky0fgI5xa/yKnubi1mI6z1aAKX080voeNO7ucY1teSZi
DlCYU6nr7MueHfSCsbgBHUXYHUe0lx7OJeN4AnBkPF/aHJpU2+4QbiYr2z1o2SyD
zLr0jv+HqNxmVvpcxb1HE3cXSFb9JlDHoil4avhg6gJj9FRhcuSls5ZXa78WOckB
Iz39ez8jx6VBEc6PH4j+IVUM2PRRQ6wbYfW72ndEMBZRoPdtg+Ti1bmwISei6Na6
dpE7E31TISzDffyZFZk6l/6BviMeQqS5j30J7d9g5h15E+WEd+tT9a8Lo1UznsRY
TRVLTuvnifqlh62SCr4MQn+aozPU4D+exO4BjAcoaMqsUNUwYNYjL3JwPVyk5qC3
Vpe2K7thvddiSG4BJoLw0aJ6jN8tPF1A5g69oYm+yyR+p55vm68hZpOXcH7YUSPA
cU48FRJdaebfSXIkWw6LxKpyVFDFw+b2qLjK9AJUADfVy6CS5nkZiUdc9MQ18d5k
MpBHtxAF4cRXIrkZVfWw8rDQF4WntPjngmv2jgdp01GyWnadtF1RFmEt8Rfjptks
tMT7Lil3clmCPg9gN8KF6OwQwFfWO+aljr/sJOLFh7UAZkO4fKt5yvfVd/nShLbo
U8jMFT3H41OJXj7ExRd/BQ6WqWMw0LfLDEJY1nH35tcA0npL+fdKt99wIcIog2p5
P9S15eXWxRU+lzEntkn/3L1QS2yagkdJ7YPq72Uxd3MVMhOYKFpP+R/vzvmwPqBw
SIURce8WoyGqUuizepEbuC7TrGytySLgrC5nlCb4Z9TaUaiswrW0rj38FYqX5Q4+
o/4sfCqIw0l3KXDQN+I2dvnfis15A3Z6Mag6Bghi/KcjXapyvX3Yk8EvAmLRTBXE
pmdVsAEFqbUBHVn00u8Aldl+X7/836RryesD7o/yQtListahtB6sY2OODu03+IK3
/4zjFCSCUJEwdUZuP2fFnrhFTySmcAeIStI4qY/DV6Fp1pwNlca9zzepS+SO15F1
yAocL2y1enfX1APylgEpC3yOZcwrdqUT3qABHyR3vpcOktlkvoOB07PvfLZrmMJ1
mK250bv1Hqx3stNqyBJaOaRM2VYseCW5RgZYCifk2G6MHM0SxtErrHLOSbnoPNFx
NK6WpedXTZgoav4iWJDnt+Pfi8b3+rk9T+6rgm32b6yJV8mB9IT4XgAU1R/CV3mt
JbB7GcFHoio30HIyVLzp775Stup4x0jJ8peGgJ4JxG/2eWgcR56Z87ddKzcuencm
55VV2UiIh6fJKE2P9LeIdu/1ffhLwlNBM73P9ibWRL1cn6iKaUPEfGIU5dpJ89Dh
2ccGjULtb0657Pm+fEoYly7uVjy/7fi2ns1QdHY/6vUz2lQXzLiauEZnjv0+vwKR
mbNgjs2ASzPhC5PGdpF1fadzaeulIRIjN61qfT7RdOg+5DDg7uHuqqkUdH0/rt3m
LAiRKApSNqELY6NjJ3zx6l9IRrf9dCNBRI5cwR0CSKYivfy/P4SKwWO5aWmDUEwI
ajuQb95ylqKm6anjf6S7TB1+ddPawA8G6LTd0TlS3u8TDivg3XnCduj9HTrrpCoi
Rw9NqfhMU0Iha69ezMAR+qYnq2vyoGNs821T2HcOTHQSmz5zxUiw+OtHr4dXgS/r
I+BqpilF54MRWbNrq3gFiXp5aymDG+wWnAAtPnOPN0RC8GpWNMqKlWnUfNBpRxDN
J2rOQ10Soge8/7WDvANecfeRMXPevlrtDab0qpLfzMEwG29RiKLxdYkanglElZfj
TUXgae5Xu3vTs3RyOdPzpTSfi3GhFzbEppjgOAF+cqgK1ngviPD9jkhROKVJ0oJ7
e99GKm6pM4rsG4EE7JxpSUhjLDPi7WIWcerQhdttiC1F8n40pJWZqD9AuiAB16vA
l8HzfT7m31lYKrrAVwZpp1JfiwfamRmJTncQJhavpmim8wrHJNH+q0kx3w5RLzgc
+7Os5KZfgaOSrIMRx6vXT8cvtWFXIMP4jnZQqh0yoyNET+u8JoyF1n66pW/+xS3Q
gi9eTIA042txorZibpoDKYs7p4UkLcOzkVnaXOXnGiwA/D6AktDjkCiirD8DvzR6
LW/6IYfn7PLO5wVEa8bFjkGy9Rh5O132Cg4XG8mSjPtz1I+M+QcukILRkF8cPfP1
odBBILyqFARPZhne96PUtppMzO2BgX0dOwdlOrsp+BNqjMWUUrBfQe8K9nYQD8Lx
6dqfz3nGLE2+GjDrEvrnm47PnqTW48iRJ43ZpOkGjMkS2qNAuN1fqpw7l+8kWgVL
TrCatXRUAowIyE3GsX8lzjnxutxqsJ07OsvPvDPY073rJ20UPbD6dtpL0Pv51qO1
bwP61OUG9h1hBHYEih3+BuS4dmUc6kOh0/T5Ur+466Qq1QyXEXCcvENDyEomKQ2z
8eL+LwtqDOic0z860wcYhejkdU2uzTJWTJH3SMqsFosH9Q1P2uNNTJEEAF5mFLJL
tIZoxk/4d24Bm6Asm2IdivTOfngY/UkwOIcC5CwrRnwC+cx2GyW2OVJhCINopgyr
QGR3zJmXRl2ufBGvkc0q7F7rQYn+4C9QNlzltTuxm/0F8J01IrUycmLSaTa4CuGN
CCjzHWkyUTbY2xfbXIuMLCfsIdr1cT9Qyz+W0ISaFB5y3HySeleP0TOJpVFrAxli
G6sosJ+89s5wxXk3E982kIJsnSqk7RW9wnoM3GcZp15rG4eM9O0JfgpurB2oB1bT
sZhl2RPAq/QY2dPM1poJpB9LNR2DMge7sk9M6RqzhG3Q2AMUvdBHzH7sp5UquOk1
R95yJWsPSSPCc7Ae45SmR+/5wFo80eOQ+iV4QNRGN2zok6SXiCYwBpf7ZZZqIrF6
dtq1GBqf18/OyOKRGVzsVEV/gh2lt4kjJ+u5c2/UlnY+phqg6ozp5o4de2kBYY69
1cPPViPFPMHDJDfT7bPA8kXPWCsatqck71hYJKjHvfAPR/qNCc5TtGQ523WLvHCc
Nyt4IbILlR+CSdLBXSul4vImld94i86ntc16hC8X5JtD7AwFhKmJDSmePjZtN2sW
vEhFIEsPMLXU77/76woqzkcPbvuSah733F2epVF9KrGcqbiJh1obsJt74qG+T1QW
+LniHSwpIiuh+6wSfq+xr9BmfspAa1F0NYtdgoVwvAtiJyBEoOfPujHtAqzqvXJi
3b83IZbOUid9+MXZCBp0NSmFWdC3uM/EUwlmvwQwfiOsmqizW2pJLKEwpTbjOP3D
gINdK6Chjil3kZZvpYtRM7lodMzSpq/cSLf8o6DhNX4ynhNGahaQztGV72aUnzCe
l1dJU8qIRxptQswaOtiXcN6RbJbhd49xLoQ7A+1RvMqlCZpA3EFnf/6WT6iFmD1q
DPLgf6/Mp9vznHqoZwSNkCcqADAup8/uA000y26WUAU0Js1zLjvJ+o9fPD1bDo8B
ZPd4lzMz6WKPx9x8Pn58fKsZvf3m0pWX+bU3eLZPpebiWyjQkKLRYWffTyIv3omz
a7pADE/2tIagj03Q+pj4ZktpgNx3EUdjPYpMYRCzEKuash1ccIJAzB2au9O3ElCF
CGEZ+fRZtNXG3czvDuHy9zAluogSA1mFalLfn/LyFrxzl8X/HKGJwM/hlLhJS51L
hJ4Q83gJvFSr2XwwtrZeULS6NfU/5TAjLduiChjqHBuPw3irJdZAvEOOOQXL1GcW
FNbaLkRdXytPVHfLeY5NMbahCbv+6VIsNCKfQ07eYX6jGzPkbXgewMOubcPDEfxd
mOHAT3k5ojk6jjsSCR/fU6kkGYGbNz1MTQufcpElPBM+8hc5MuENMIZk7Q8WGiKX
6koxaQc6Ywli7iw68o7WPJhS/yd4SoQyDYah4xfDiO9pLXKqBaXsQefLziy5PJwW
P/twafurFB0x/M6cyTSFrmkGd8IiGzwqmBmcnu7ppTY5LwAW7HGTX1po+Vh/2Bmb
Hlhj59TutdFAjxzDELQIY2hAdepMlV2CYzFG0zOJT3nY8QgA9eg022a+N/GWT+BG
Iq3qdQ8xEHJ2hy2VTweGiLYtz6C8bxl/P+QlNEvgLNaoiuT8FQWKTWeRzy4iwKAk
ZWfkA1iNMSEaZcRPlLRTLzxTyfwsrmfM+oJkk+YyYc9uaMrl5sAErxWWYkT/jmp+
M4QxXhZopk7QXcouOooNjCRUZpVhntHlMQmke+W/5EUwXfOUCY15TkLLJf4PwZZC
exd2eo+3V89qJsEyhwrjx9TmYyg6SDDS4ePsz6JYjl4IwWW5v7ejXAhEL5lxES2h
FBKUNw7aIxJAXXbbIY973v+3xlEz7Nc4ENZZAJh2OPbUxW+OGDp8jlbI9FZbBe7B
DWZlEsBegkJHZerwXpqTFdVguM4SVvmmtqm9I9Am1oCo7p0a7BVZOAikvpreNkm6
ZITC4ZMHCZq1Umr6+X82wToI7wiGcQHddHMFRnHCZHsElgvwgYhCOPmZp+7MhrnH
UQHZD7ZIKBgLC6PAE8vF9hZybuDEBOkrWawEfBHW5j7ylayTzJ9A4sBoN28cx6ep
nKTIBZfPCWaqyUHijLDnlrwO4IEJSYfRy/D9ppDDozeLSzMe9Ko8jIrNBE7lI8RB
RjBPyXwdjVIL7Po6xjTKVqdVszYK8TrgqlDshBnySNSgIPjWDnQSkL6Ykss6qKfg
wl10+UT0p3VRZKZxHRGwpsmKzsS1z19Ab6nUOLQEoly/I8iemg4Ir32UZZE/4xaA
aiwO9do6oFYftCVHCCQhlJLi9cZREOSgYrVpY3EWfWfbuGGAFoEoGKBNADkc4YSo
dLwGXewv5EZ9cdwXcRQfjXDMt4GRmRsXGwxxIfzowIWLnjOIwos+/GDTSSpTyhCV
M05hWR1EMS92OwyWr7ZgyJJG7hdboK8g4tP5i/M5TBrfIfLM0aXGdG5jWb0g0wJB
smRFDYxKTk+CLzRNo+vYqS5r1JDqfDeTMyGgAMlOzE3ulEoTKwoHrRBaGK7KB8yJ
N24MAQ7x5n17vVax/CgbnHuqZWYOCJ6zkhX6PETPhM7Mybcbw/L0XOJzOGB85us6
jcayIIxb6bvG+/xgJgAa5pMsRopcXZ9bkzy01FEA7tj2YtrW9XvC2tLapRpSz8pb
r1kFM0Y/Wtc/NMn5on1wjG8THsw/dyK1R+dsv/GRZo13x2EoTUZHL+SkxP5ix08l
z4kEzYwfXVf4LFDMWoQS1suMLex0DE9FdZ1ayLarehAKZ+4nEhNQfivL92aFF1B3
zaGAU5RfAckZdskzYKdGo3/4st5SvNK/tm9+g/UGV68PH23vwACwlH499hQdsAKd
GnDX9ZrT7B3czZrqoXp3F4yIMzys7NJBgL4iwnBWQRADjjArW25laq8PC7PzijnD
0gXTtoc7sbeAT5yxf/duklMldBk44LCKMJHD1NF7g4+1eZ/Ar/QH2UgsUHPAVv3n
c/BcWrtQboxtHduiVqtBWV8AMiccgJPlA/XeTG7LMCy1yX2vADRp02k67N6Edqk7
CBB7d+SBsVxZ3YnriRpjEY5DDtk5AoZvQtcbiF6aeinUQh9UOsCURYn8f+4JNEIr
/BwdzR3/nDl2Yd8kjIMdOrQ2CnPL3JM7vGbNUZp5OsLOvP6xAsFBqk1yv3iJdoQu
Kamywh5nPnhPOH5x5/pCrvTpbJP9raPl5RU464+KaeGH3WlK1ZV47HBABF40NDpN
DQlApaQpY3AQhQyKmOd43V89dOwc7tyCWl66aGKJUvmYoOeMdZaMM0FofAq3cmXV
tW09ukMQTwFxgCLhRDBys4IerBgAV9WqxWkZf3DPUD90KNFyrWR0YjK+VBVt3X0C
tLCD+jlD3TK/LPYPbyA2z+LQm4ll5H4jEDO+JJ/Jf0drZYjYTrG3kvUhVDjBXcfh
ZW1DfIWVEbOh3y92r2rnrZY97dWGDiwjGvCGeLqy7miP9Xy04NcVna0FQNqC+vaA
G7CqpK5Y1oLBzzqxxEuNszQ8Dk/SSmndt3z5pmnt6Hxnc8xN7bqiXTL6s/EjOM6n
nVCcsUNHqFsKHKiW/zrYc9Q/pBI2ovsKL9bW3kuBZGUNrLSoiSu06/SvO8zMSD0g
7Sa1oOYDmqO2O4X3WEIxbXBOdJaiZMR4XE83z/0cfrrvjUGC/53sfE+xKgu42JnJ
sKUXdr/3/FzbWc2hK91Xc4RQB7B3HcxAReC9DbR18dgWkaw20wGtQ1+JvngT3Bgj
lcPws0Re/rQ13pO1l8FpsZKeGE+nPRAeTm2vxQqm51YMRwvAVWfqC5wBH0wUMVzu
U//Vwumm6Xsi2bwXKhpn4bEp9Eho/3++v4t2BqXIXOKd5CoHXG5hfcmA5pMo2vPe
RvABCG+3/xNlayyhX0y5U81wkqw9yzZz9jEGIwdqSi6bPtVtBT7JQ2UfY2fqULCt
XMacy4n2uGf+sQm0NImto7pXkjmhtRPvWjlf+2IRzyidd0BIIm6LNiZQUyVIeLPL
fjdNRZQhJwxivKGZcu13DGdiXf+VEXH1dBO5KixgIlN+mtA6CpH2fHjYRK9yeVoP
sbvskXlWyrngAh99O9DpvpgI2NCIJVoU5QDG2ItSpX/SlOOj5ywW3iEhJLK5QkUy
IwUV7GXdX+S31wROisk9HvHyvlZ5ltU7igHXwP7f3O/7b1shNpKczWNaNkvtw4Fy
Mo4Vbi8zxMul5FISWcNtfNR2gZKXsNAC55EHtdUsc6omHumNrTZUr4Har+vj9zg0
z28r0e4kTaKKsIVBRqAqBl7Q/WGCjDoVT+AjPw+aKAOJnLKe8vOxV+5m+YPCvSRO
1dsd4G80tLrvB1Hr47Ki5GSVZIPO7+moY18mdziLoD6xr4Qhm5/mXO4LvljoOOwj
K/ksleEPwXsG36/n06eZgnX60Kh6nKldUHLi9ciCQo+uTn+X6QpiwhF3s2BvOjYT
bDfJpQ+/YyguDWVyw9VdHJ/4LJWXnC9e+I+n5bLuYy6UXUKbzBmhHW1ZQdaJ+dZq
KpW6vuQ91YWnsDzzjPMxX3nWDX9QSNnTRgHtjzVYIxce6gfV7bHjUPPY383r1/5U
oH7FLF1EizZeg9PfakSoG+eQur3n+JnOQTYdG29OnoPt2pKQv93qH8MNH2W+5hMj
pTL05f37rf3tF0JOwIS/K4+lXyOflYjZHanTz0vLlAGlwL6cJE/0z1agg6k/7xYK
SCp8ZVeBDYxWGBJLrLPJw4TUmbfgfkUYdtciu5bJA3oC2PwRpoUJm/Ig3FIv9LW3
dMP2daALqpJ5Pq1IEyooUZ0UgSYe8+JmjwiSAz7CGDRLWqDQ6U7bGtioKCwBmKs2
WYNZ95p6BLt0Goih1XzA9OqlSYfFdM/wnxP7BJ96n2kRUFUm0LcuRQYg4vtgB6Xe
uO3uSG8BbCArRYqhI8YDBhZwCnSXjtHrhiGLXebyLJHB3b2It6ovD6PGXAfWoPdP
bNEQIRKItqn7UQRSk5Qr7DyRrpzPAARLbGHdNF5J7VTpgZ4tYDuxRWDSxorwAA0c
5fXzpuiwfsVxi8GGnHG3dIwBBQ9r44f3/a6+CFuACVHO1BP6tQOwslLNocwCgZ3Z
DoI35m4KqHeQ9/LTx9BMvRbtNnphYbWTqhKx0abDAc0Nm4zG6KYD5AzSAQL+vYs5
GRNo0jjsFb1qwrniplm7SAQvtmlEdRDEczigre0Xng51lgpeofSVYRNRafes3Z/Y
Wb3QPBzVSAt+l/sUw8cPKpzb8zKDonryxEa4c+ptQWeKMs7WesV8Qu+1pgyH7Vsn
f9mqWzFN3ISvMvq5LxUyE5wl87z9//cibevx1ssF/3DO2dfDeuXy4tCx4ci7f7kA
faZKVTo42hznDg8oTUgMcsPwRITN6/ATDhwaSQIreAId9FbGlQqSrgYPv+CrXIP3
XW/ioyXrQEHBlJ4p9yb+sIML9tQsFKHblLQHt7jFxQrnGBhhhLkkargzKiimMFdi
zsChnS3aJl22Hn2VWO2VH523OzDgCQZmgVkH6Tg7UYRpzj/0VzApqQsUiAY4IcxN
339LgQkXEUzYXtyybP/2ggTZe1YjIkC24b7krcIo3jFtBUnB9iAh+j+9FIjZCZIJ
A1bQTPHKYG8YX2qMLmuTnrvsVfWXXGvE8//F7HXovTU+N5FxToKkm3PvhviRSz/a
vHEqK/q4YFk8mSdQxNvB1MBA7yXHpYvF5fTu3i76WkM+SsSCzTPvtShHnEdc5VfB
SOeTwOX1fz4ogZMvi1J1E9BfAN/yQlvwGJxtziTE6DiZBrd/MJG3rh3ZPGTEBywy
MsS5bF5XBBGtKFhy0YY7x+hdG+Bh+NVHtOcSktJP93C8dUDEJ5zNCKNeGY6tbTTE
/xhMXFxV5f0yOPdFMIdqbjK5u7mQQCKxLwB6d1LjBqlZu2N4u8e/DPhGoGIy892Q
3Xa4AnVstAiMBo+barVGZmetEqdYWDXC8v6B+7R7GEL0igitadd9egAEfqXck0KE
J1EnxtaMNiAHpqqsKHvD8SMdZESEh+QdNIak9yet4xwO8OVRWwY2sPlB018p8a8v
KmFfIUgHbjgNgosuHCxjbGbWYsjYdJhrwqD/ihvPZBw4TbfVX03qifU7lK2Q/zzD
nht0wFndorh2QqpNqzax3g+rLtcskM/quYMD3tFseeH/935vmv4XvqU0GcrMK4pU
xn5fkpKllNMKw0IgqHDcCRj/qxE7NxX9ErskAEz1ByEfl7jH2U9riEN+0LIRXrkr
lYgD1vPjJMbaiMEIDaSyvxq6Cdy/CDC7FsMw10aOxh1VagulLTcX1CUWe6UGARSW
HnSuez/WDo+jDRnGPoDdlRmg2LnbtntRh/5CBE7fRAYYboxjXEYD4AtdMal4d5DQ
CHco+PvJ7Il8dSu/8Jssl+NFwH7L8dZHikPZcGBbgONBiqG++1RSavNIrg9/q42c
woyVBwaCbyi82i/cZkc/PCCRJAOGKpzolwB/FLsoY7iYXelE+3HKNrcBTRxme6LQ
2Nz5xcASqZHEEzuSTFgbYn5fhSVFXDy7yQNFRTEZs2Q8Uzgwsg6znXlMikaBFSBG
iArANACvdr9k+UGHIMdihbfPCcijZoXzuRpj+f8hnj2FRzh9DS91c00hzt1a4bVy
d5OafRkW8mQM5VknZrltL4g8izhC15+cew6tlM0WP73RvvriCcx9ynBYoQpYTB+4
Y0n1/pvHL0aq7Fl3PpOtnXrljVFjPHn6+CsjXqGL0pTb7KGd8JNy4acPRawwH3dk
3PsTK3jIq75QRv/NoS0HTdOIXVf3e0wycrPJdEDJ+NwVxeeqHZMtKFg1Sy6Yoc1T
tXZVdDsGuwH0LP9c9EgNA1kJSmoIKRF63Lg/JbafNSYNf8dTGLVTksl3tuzhJM3X
Qhf4yRo7Fs8GKThMFCsVAhLueTCVe9zZDo50WQjFU93Skz2fa5YDFQfkpu+QG95r
ly4c5sPuh/b7V8mgqT+SMWEonyxyfx1cc/qKO7CKk4OAr0rNfm+BU+Llj4AGlzlr
pdOXGh8st8+EoJZKFIOgmYHSg9qBWDkxwBqira5sOPYSad0UuBEmZOwy11vRv5uj
5GliUUMjbrZ6YN0/snczGds5kDGV56MVILqnWqFkx/423r3T1vRwGCcer6ofx5Om
7YhTURF7GsodOXEL5c08qDMVwhaVvcGUQ1L5v9LHD+vn+pEkxNT/NFtpuCjqZE9r
1cE/WF3G0mtlwZG7tmvAx0ofym9nWBOJajVrpGB13fOp+PYu/iEiw7wm5r4iqu0U
WezxH4RpbfQXG0OvvhZZHUL40+A4DBVeN0ENofs4K82vV31zGNqoxZJq2dWM2nRa
qxUYdVQEzoOH3JEea5gLeoI1pt+85mdNMCXW6howVG7tQIi3pmATjtMKW3PuYRJO
JIF1WX6DQ5mbB8IvX2bZnbXFDuABCkiR69rejWAgGKi3pDoBVgkLFBYhvFhzYVg4
Fi8CAiDlAlOBte/tGXSRvB3sovJY5RHlYdqmfq8035WI8owfl26v9E23BxAP3eTH
VjOAUED9WdYkW4QdtrYUyXMskA8a8sjynqG+TpehkXFC+Ys4xEehBJTR6BDqYG7R
Erjnr2W6bzvaE6thNd4C60Clyu7B8VdRvfRSgb5vmfjvSTYu6KZ0XwfLFRLybI3d
73irCpK6jocO8lD2YrALLVctjU4a4Sc18LolcVOTiUgCy7SW6DPJMH3yWGjIRlWk
avoh+rNcUI1CffEj0qx5ziQv4UQUoeSpSVoScMrM44CrSpOzFckt6GBaK8U96Kbl
puZvd4qZChqEi9owsr8OfvAeDSOVQZKH9Un0vzPbeUddn3xjQl6bRc15L8JF7Ni+
umPFL42R1fKZORRAHorCybdn16FASLJ+jKf32E3kyxVChgnzb2SfD0q1GTGKgrji
ddpwEmOOOrx+sxgpS2+TDXOF/r2ya88N6KgX4ScQjqspcqDGjmG8u/biuBROdi+u
NnWb8TgWoyOf7MHNU1iapprI+JM48K49lkqC2N+cxuv1BSjb37tNj2F3BBNJIGYP
fvksJeOSptkCdYVEzgkknA4eB+/eKtPRzaGLbwOq45nF2WmkXOnXetZ58NLvAik+
3itkt11SuWPGCLFP4Gmh85MXuxlnPWv91KVgAeRBoeiShxgKTvfOVOJm9jPImdF5
d87JNe6giQdVBWSH7IduEE6OKcpCO3ekKIA1NDh9wmgjo52mc8uNpXYFe47PM/A0
Fo7iHSQ40vPyt6HelI1NIjpYue3ooCXHXhviJqNBmQSKs5N2Q1cE7p+5F6DjH4/l
wwWGf77ERw7dJXkTP6BVau9MZHPauamqvpstZFfDQRk/lSH9e9NbjOO9Old8koeB
J2DBn0YmQu2RO9CNJ9E20OAKMTDj5uwDgC9no/pfa28lx2yq2RUaTBLIvUeCwvTI
3i2AMETzHThuPPWRojnoi5bBgJbgY5GZeHtveOevaxU7isQoGh3DW7YLo1xt2Awi
UPJSsq23bLiHCajDguAGgXcS44msZijejgWVSfhQ6BdBv5Vp/CVM6Wmo5MsHtxJp
dPz/G1euyGHXe6n0sB+HHJiDC7TRCoR1XTnS6SZipeKtM/uEsARVFROpc3fMF8NV
7ESxlBMPfA15IClCmsoWlGi8UNobt6DC3d8hFR9Q/9Xc63miqgnHTFtj2vrsR+M+
M4WVi7fC5eckZz8oNv8yz9CXjImloJfhvcwyAem1xPK6fisTc1wmhMdlVF+1roZm
pwmuuZn0zag8tCfCQKcgzNWcyKDy7HAmapE6h2DYRMzRXUejk23/sv2JFzX3dcGv
wWnSubw1ZL5PBM/wG8rqNzTsXcTb5+MGUpBG8zC9lvfDhJfIThGMFc3g8vI7B/hD
tHyPbxDO26ubCZO/w6LV40Z7euD+udGh1j75ddG1gQy+JPdRnt2K2n7dgfls0hlW
oYj4PuWgzVvh3YIwkXQWh6sKIFeU2+lMr2zvklOSz4SzL19Hl0aFqZGoSQQ+W3XA
E/ujwwuTMtEJQnF3RB+pIab3nlovTdT/LnNLwHtLow0K/9fJa0dMBUmKM0UClqyu
lRsdqkSUZQnQ+yDvFnExa+wolGN1BX1xHFoJ40YBA/Jwr583/p9MXvYUEC6wVbSc
GrNI4n3ZByAgoFNiM0YWECBbuof5tjlG0n9T5U90E1obmlNncrvQ9FVVLEEeTTjf
mOmeZ6YRNUk23y0DHFlmxm9oeymbZzjdnlyKqVQuciDGmBQaOrtcKYGhpASuUb/J
2ZIn/E8Io7nT5nQGelmWSBllneuhlPALYAwOd6KQk4YahKaX/EKcR7qpqveCB9pa
NZsjSIfRFl22N2jZgKa27AdsdGC1D6lAmpa3iQWO9o6+h+8xg9Di4wGo5Is6INXm
xy1S5A+dCb7jXqTZRJSBgvzDNSPzgeePY+iCgDe2zFGaoIP8wSPHFW7/abuzTg8c
RtBjBwzKRenMCaRz2IHn+giLbqQJIKlp3JyLZhl5twaaZ/hZ/RLOhttB1sD5eBFx
rJ6qf/lT7d1tBWPXis8hzVRQOYPvk8nPaE7DdnEX67Q3+R70gpHA/Abz5FOWwxLt
+HSDreVwLoaB1MBZtmUjUZqKLoBexssUAmd2vn5iTakjPruOm5Y6Dfelj5By7wKB
7NNZfKQs20PFn//sviZR4w7sNwbyAa8aPY5DXdRNhm2fy56e07cg0REAW/LSL+Fj
ALiuvStaiypNomQR5XL5LPjNhn6L7j+zPtDTmlym8h9LD63dg1ORd9jjYdkSTMiA
Mh/schUTwEdkdKAT+tZOkJWduZB5wxbUftEWjMUIflIAjathDuJyqEe+jQnoJqB/
y4otJsn9u/u+Ys8vLQjlpOEKErKNj7mg87mkYeP8L5nCGIrnls6WCf+E4ej8sgCG
haf9wndZz9e6bamO462CtDuCTFun+M1RE9BuG6hqA1XaTr3aPbG/0HL92Fzx/0Im
ZZcf/EHQCLfdOuZ5DyfP6O0WdB8tzGVqNwqK4FP0XM35MCiKgkMH8b2VhzZvzjam
U6w8/oCmBSuHcnKzwg0mQcatLHSYU99ovHqRkBydh8O40bi8zuFQUtHC+tU0prWN
LqJl/1F/gmmkUkQyELRADmJRmiDWw3SxDe8Zvhegoj7L5YKUYVqZ1HIK2LiMhO2M
3GP4ShrrI+NPCqsMfFcODNwiO+bgGSbnZDh1xPM98OVeYXUiq7jLwg2mfpgmu83b
3GT64RwEWmW7NPV2DuvlCZGlA81q5wfDdHm8tkM2n0wf1/eqDP/GCgZs4SeoiUe7
F5bOPwEMnkdwo6EEfKCHa6azfG5MVhgvAv0hu8LY4UZ53/EdrrbmG7u3cQV8DI9W
oRhDplFZRXXxlWBBo//jM9XBgyxeajzmQ8BbRG0k+xiUil/BuBwesbZGhRSmQzQo
jJIbVkhRZoyPpweVNhvnlUrJnjhL/nh/6XSeCHm0fXjmuPOF6QKThQNTMzB78RNI
oE/C59IZJu1fuiIussm84LBZJAKiljRUj8+N+E5iJOyiBcIJsJncU7+EuJyqxP5c
b1Rhknm8ArJltSlTVDX9JxojHI/J/J8+15Q0D7CYQXTldtnRJIwYReKd+dH9e4xB
7Tw0Zm5jzD+YzEzsy1AuggqkQlr5uInopLgdiWH2JkEK/ZO/N3cQOFG6BpYhmwjS
Ig5dnyN0CjdaiOKpbT8rTLkR2ERCu9qellYv/G4q3oZBBewffS9ZgX4c/CrSxRnD
UL+m0d7/e06VXeiG7Xv4UImE6mOvSUE2qPGNMXf3O0FB+WPo2+OLB8cv0jRxJtqn
amJtNsFOZFcEs2lYOuAtxa+YX0hPjFBCdmed1OC3NzcbaWk9/GBcDAsWpfoEIgTr
P6krwhnOenq0d+F8q5/thI2fG2h7++K3wviLcp1cTu06h/aSTXW2q/PFcmHjKeQi
/OV+L2G5CwZaAnLHy1iJ8SZEv4FLA5NZg0uf3nK7On0BidaGIUtOJKKdW1ScXOaY
om8feqPjpSgmFnxixp4LqtcsNVUbv8tu6ASauye4oACrmhFDeghlIQWznMb3VPJF
omKe8rhjivNYF6iOroz0MuUJkh7kuIo9yumcoEKIWRZ2+ngOtXxA9xZhZaoxJezY
kqPBgNFU3pN2RMG7KDf+udjFsxVcOAeTmn5jZyU4pW2XQWf/cWx8hBjhTYIfl9sj
QD3hesdOZU5vgH6KgHxLcI0IVbEFWFVZWkps5rBom5vzxCeJAZ1MPewmxuf4vU3S
+uMWrZtrRH2B99c6bWfqbqAAHdXKQUmvf3Jdp4RHDC5y/kaw8b1VM2Teouu4YwG2
/S7swpMQyvRKUk0G3w80cyb2ouU5G+n6DvYEkHyY1APWn9M0k5/Fy+AcM/B9exvq
2lyecCdJm0W1/pb/jl1BbHo81Tx2ZKPjBtko9LNy0VBda69QK6XHJcdOnV4k48F9
Tk1dyLNxdQJJKKED05P3jrwVVIVuhiwHBVnm08Lq1xz61Ye27AyK8OW0uwuwWf/f
7Ds1fpZXO1/GAZZxqvyefpGdyyAKzhjEuELjXPH+LWg4X2jnge3pmMdajs1WY+i/
P+NqWOU+spDE4frKuI+ZK0SzZz9qlVJXCl6uyjWO/QexbmZRr1nqC8mtAvpxCd+c
iJsLFwlDuVNd0jVk4RN3+lZIN0ETQQ7XU9XxFINqhxM2bmGwkU6LQ22TsYZjYXka
RhD89IR3r9UX58m6vk6h5T2q/KXhVk1VLkoHUmn3JZy3volfBbPOIv1W+G2m2/um
0YWsGKuuVHVbsuvL4wSMS2ejQWkLDAIu023sAeHHFIxkg5uItl4vCZCxNGZvQeXA
qKY6TebLFkal1qyulUov9cSNaSBIU5acNNfEAs8bmq1zoXpQ0ykllDtlyQQzkzsa
2Pzz6BWZy9jtcMptcUhOKXJIPdE2FZrYbjy5xEoa5m+7RI5DgdJv4KazciDXt6Cr
r3BsUH8yNdr9PVQCPqjoUqmmUQvhueHCjB8xX1nC03HWpOOY0ELCiU3JyY6J2TFA
ieN79strCb41BY0z8Plr7jHDgyz3AE6gqrVQuuG0i6rhR0TciEQVHeG6wXd2qWVP
N6sH8Oy8jr8Qy3CkthxQDHs2qnNj1QqOsEdODpxtjxq3/u3U8o4fjo7sZZZrFUqn
3J3dMTOpMEkStyh3e9ikI22gvkD9GBIDFdALtgumY5wUOfd/bODo1CJZIvPV+NNP
b+PH9g321cmk3M2vdSbWHt/IMAhp67OeY3FIeuNtwQLepZdHNZ4mt+lGXOatefwY
qLyP5seNdXoN5wKySUgl9TQG9sZ0NSHElWohxoSqcZFFTfDAW4wTV5N8VOn0TjHH
MX3QyM+lk1RTa7Npf4ntKHUy8MDqwfCSTt4m+MQqiFaahRxB/lOIrkEou2emcKw5
To1mlXegL9AGOOuRVzuZSjR9Wk0kEOdwTBK/i0arUGmnq/aRYz6VStB5/tlu/keE
nGJmXsY752QaRiZRKDZ5k1BOjud+UrkDBgHyQHeKEn01Q7xcxLEic0QwGKnIvN7u
X2vHXS0VPLkkVFyrhhHTbYxZdH7ZFuv/POJD7K+RASZI/RydxqLowq4MAQw4DbUv
yEhwKwyOlwAbrVFelDkj4dPcCJoNvYx+YvR1UP1QzZ/PP1RnAeDD8UIUpPxzzojh
9XrqWts5GiIzAWkcrSIYitVtfj1fn1WAEpr4jwOBedAWEPkPkzYh/eDvqVb5smKP
1VThEwBJLxDotau44rZUjxaMPxiSlL/AxLsqaizCromXissZwxm7UT3rOyKFlaQl
BGiIf1okTHgirfUlQne1dkwKNG2k7YJqSaA4tuPIFp8ay7HrVhcR22YaxLCiwkoc
SMm2RGl95bXEj60BPbW+6joNaWNltN6eX2vpKhsSz6PoY5XYc7FNFrRpQN8A5NzV
S0WKU2YxqqyafEE1fPmuz4KkE8JGd6tt3hGWPeRpT08DXEeLv6qhmZ3vSundJECg
Gr7g18jP9fcuo/d0EqnLUnUZ6CaKt7uCR4vyUDdleOR4n4E0Bfsbsei5hmvMZmF0
Z53WpZ+rJeoMsyrlQch80ZhyAFdPMefB9eO85lYyVv9DWy/yNoiwSgZ8d5zbx4iq
17i2xj3kR79zV+UDhEhuBl9JNN/u8QmVCmwgul1HEPcc0416+vY69bIBvbTgpnTC
13Sb4UUiwQLmpkvCp8cbRP3kJtfEDVl1Q+LR/hEAJJSUjJL4G1Rho/WY4HsNlgSi
K8VqWklbnXWsAfhEpJe/45Mr/WGdL/P1ZVN0KXDQK0UWxuiSZiiOcYMt/F/8yQSz
NfmOiBVNs70lCRNbIBY+BOgYw/IAFPT5vetvEnJjEwhVWTLkoqB+30fiw/uoUbSi
06UK+nYSrKZHpfLfDxMk2KPF7VnOwkV3yNf9pwVowoQa4cBdQ8yzVW/YIvUEhezk
mCviRVMs0QcNASrGxwNqAPk+C4MxEZlaZLVuvaZUx88mqQUlgeJ+Q6ijH3Cy7bzd
cav0sozW9DRmj7SBv3AmLrypa2R95C16cefX3S3z8lc0RCXosTZLBvalHeoshgIq
5p12NU+Lap7iTapGGMP6uY+pDcAFddsg8sNDrYgtuRux7mDQK1mkUxf9XHpUMjnr
eudeQI/fKawu4jAjyrqv2SWTc9QRQvmH6U3GZcRvxb3N+BEG1ildPZ15LgSLTH4V
+ulc6ZIbKFlUk3zbueUDMdPjsMN02qnzQTyDebHkN2KC0DyhlvywcT8dPympa431
gsQIj9fM7VgO8mAQrQB2GIJQS0I9t8xbUlY5MORK2xVGS/WtJx4ml/QwdlAP2Xb1
LIepWnS+tvDANkQ54jVpDeGoF74CNSJ1ZqPhldp5x1Gt65oBPPoLC5d5kLhte9Gs
dIxHJDcpwTnbllHr7ZjvMlTeDUfKANR/2HuJ3+75jVXlkRsmFlzwjkHXiENYFMZ6
wtG9v6pRH9/fIkYmlANbmF2G9JPBpx9QlVVbcI5UqX6UMGk6eG67HrQs1Q+VaR6E
I5LwCHvVnNGY6nLNGyE/Ws2e/xWugatvW3yEhNc3vN3gEwfxOJ5YwklCENFBU9S7
N/S2GtLlS2pn+8Fd/Wbnu9hM6RLKf5WQ//39nRzZQHecBWwcLwDhakdf++CBhUZ0
RsH1Dv7gJSEi5YXIXeZcBUd5+tvpzviUWW1Bzj8eRYm4tG44EktmqImookXsGmZM
ktawXoK/hnuh8F7zby7F6Tg+Co5bLzfIQYtdvV0AIzQrg8RzHlPjItuVvT862gdz
llwpt9fVPfbCXV7TFYdBPBAbHyPlhX2LX1afEAIPK/k15OqlIkbXSr3d7ENWOR2A
XbSExxY1KnFfUb7skHB2aYyyPbVeEqAtXhGpCGgBlEk4zlnzGDz2R/Y0qRXhhPib
RMwBCWzpqj3/xFmWW9iRqYpeulhqq3I2CwHlmz6BIVEHXEQ81XdsAa/RkoVL3mNU
0Sb3/llMOXpJiM9jKnHjvWqyPuqjLnrQgQvDtn8JVtpClRNOhAPXrFCzF3QcJGYt
QYmWNKn+XOCbsd55MXOPmdsVzoYLDtFGAR+ajWn0HZOQhFal8qXJpAkse9CkVbVS
U7z8VOUPcQv/XfDQU0vnbWucr6aoZukzIi3PJ7CrTkblGFN+9hm6NdwwHyt3y1RP
3uyZcHJ0yQ4jUgN7nGz1sEkYVNK9Pm72xJ02wTs/eLFe9ndBjvmFGuvG95ljxHGk
4zG966znSjy3yON01C2yE/ezt2yT1U2rTcF8ljpYyXySxk/nXABDR8pWX7RtHstl
5hvvcfKa0s0JtGEdXsV8/i4R3Km6+Z4azXcrmcJzxcngKzEEDJATnbnAk1UiIIt9
/M5boFK93AuBoEtq4gClDwYQWAlLZzQTflZhKgAItK1S7T4o1LQFGbFijidzr5j3
ByxT5nLaKIxBGMSMwLkdiMgps04k1iApCDLpZlmgGENNLKYx5bcG1bahRjKiVG4o
dbq/DGXaIEnMB6mhc/H0h7HpzmFzMVjh8D3EGceIZS7jU3B6dPYdLzxU7tWUjtmz
zbaVUYQbJYRxXxd/XJNEkgD9fS3h5Ky/yVYFxwkLBMDU31+O7BqANLP8AMuiqE0n
h2EmUfiiIkCLgE++x6imh+HWII6nf+Xi7/W+0q4x6w+IX5ABCxMwXa0k+A3e0+oD
mcOB/rQnrd1GW1gJNOpalg4FQqHYSE2GIua7W5yM3eTNsy4Idqh779HsrWe0Z8lT
YUdX/dFNQc29aJ6jtTtdYqQe7LBmZNrsr+hVyLlb5RY9M9jk/fzf4dVY3MqoGnP+
D7SNqBlo/+Wqj+vnwOwpgc9cnSOq53SMqdjcsScQC8iMAca2hmNpfq4fKTJ/iUqE
d1X52OlNw2IlvahvCA+rLTw1sPd/+2rvWG+9MzPWNI0ymAC+AmsvN9uji2RFjYbM
/6gTp6yift3C+n5scT2M8tWzp+TMDEgdlqoY7IrCo2tiXWaEezG0NHVtbAoRTiTw
U2fFGtjoE/sh/sGfK0u7k0WvC6xJWQPJdTABaOc1RLo4+xxHHNr1aROItFrqdVfh
QpjO//BGTQs1nMb0/PoEYP6Xy9f2zW8Vp17vXVG7gvqkzgbSpcuIfSEzcUdWdbWU
iW+Be83gDYYfE+j0OPIKaFGdjnpWw0p1LFUOScRh9WNtY0HyiJrp5h6HB/BqnSQI
/DpkyVRobcEATz7vcztoiHSn4giVmOG51a8hUt7qcCnxjI5qUGSBStUnfT92FEvL
UppY8b/SjFss2VE9GekwY0wsrA2TazmU1f1LQIzSy8KsBJExSM0cyIaitqbkdoNe
4Fga29gGpGwWc+V6YJTH77szfwdA2tLrElAIRKM19czqsBX5M/b51Go1eII6KoVk
lj4m5XDzNmSV/bYuMGAeoWbzTlyNAuXVB9eGC2nmFZiRGda3AohZd1xiBV+TOgse
mOGsFqv/tQz38ABLG1k3dOLIr+nHzgRM1/hptvYvcvoA905LOhbL6p1pIYvFDAu8
yZD/Yg7Lp5iD/r4zJFzwZpDyMnxpVVhKDc7DpKMrGUFkiwHVv8xl+4CYarRhlIsj
6j6A3kCnupaQhpP+m6TmYRkTQx0NEdDIOBLWSQ/gd7cfwmGwPUL4iPb65piTBjL1
oPetiTn2UedJl6LWU6iruVqRKw40fRspHtn7p3XTZcC+90NHT9QjdVe7qnPXh10/
/xd9m8h9mmCjndiiPA7911La317m06pqpMJaw9SuLP4toMwkxrY/iDX/3jLwUFFY
DN0CWDAZjMGfMmQEyBSmTKVhEkJ7CE4DUDuSZa2bJmAvUTYyq740jsc6BlfJudZh
SPgH/La6E9SJzT5ac9HuHjKoixc66HmZDRiZdUXnNmZdi1vJxhZ3aCWUIh6QarBH
+o4Y9vBpDU2wZLsgMKvL5vqGUuucmuYIQNIeiHP8GQ8Pz1qN4cEjKZjMMvyUs/r5
PDmFOAHzvsWuucKVCf6Hvrou/suSxams1qn7O4aEubzmT7x+zAlEeK82gG0RpINb
Xgx+btOa4HB8UXTIeVlIimU5MreB8rMN7Cr7xGzPwqh0Ym6bfx3RBTMasHOfNfRD
RNduE09DHqwgkhN4jeXoVN9a5V7tBhxj9XKhaKZ/KqE5kab5pIsqOqqvvY7q1ZUX
lHkv/Z6mmLSHPK1Ebx88iYX3yT5HyYu883avz1KHqZHsanlP3ccLofnCTRNnwLGg
HuR99WOlRRounXLvszU3UHDmOz4Sf/+T/3YuegKt4yco8Azt9hguxNW0DK00u4B6
fSQv83f/pjP5kadmDJIlszw5IbUhrTgkuVKxqwYpvgqLEjqpW4FqUs5Z7+yA2qLm
j9+ffJpGfSiaw0LDXVIY+6f648Q7gfzZUxtoRgthmJ1WBAOjp9fiJVmu0acaJZLy
LyixzzoAfi5tQpgQYEKFNrJt/3RhoNV0WUIxdfrdnI8J4jOlcI8oigv7YkEwtAzt
ZYNPRiSQaImhde2NXQ/l2ttuiVI7D70dpaFVdUjWXebhUGOtOrgRIkp0ho2EeCuX
bzT8JEpub003jRq+XxKOf5BvmIbOBYMqzcl+T1B9Ja7i7tAPqoMxUeFufUHOJkDH
5GvkB+m5/bK0EEAQnsTe2P7gs4tMpL8ers5PncB3suYSRCJ1zGuQRwJkHvoXRhsZ
4QBS1n6U59URyVHiEVJgfAohNHd+fXZhG4ZRFUA7g8yJBrs0kQoILVCBFtp/S+BQ
9bG4UTSR6EkurbicjLIcBWvblwmSOa9qsfHpQgwgDb7Xqeb5hqKpHd1BKXX4yRNZ
ZIXZzs/4ypLZMm+am/WmTMa1c+sBFZn3yiU72Qk+r4S5KYnsGAU45yZQTyXtY/Ks
h1zwZag/65NG9m1EEXJFJPxiukpAuzrKjwXx+DfzJQc5Fqy8w7rEtTQHmte7rZUH
Rv03CvK57McHWCVfUl7NN+WvDMiX9nIvyRgfaNT3Sj/DSfMB24ezoEB/L1hq9G+h
krGAuNnZ/6ay6GknH7PFLTrZANPCmOmELDADbNDarZHcT3/u8ZpJMRIu5tAJ5rOu
31W8dPGKftSCIL9RbQaKM8TH3Yy6kxy3exB1d6FwebmP9N7xpqwOxm/zCodUvRY0
SdrRdce4I7pb52jjUPNl+yeVTxnQMT4yxrZwqkwXOKQ9JwUYVfvC6SC4E7wkF1vA
xWwN62pSB7gAbGAENLQl7LzzzgAg/BpIzro0i28rkpARlG8K9WUvxuuhf3wISshO
KtiKtCRMG6Y+QqsbazJTnHX+b7rpvg1ZOd2dpVY8iV4PlOKi6Aa1etzMnMReJ9x8
YyRXoBDf9kplqRgYbZy7UJ25ST0hYd5kC/9YccAGUjwLafhqrSrWKzGexROOcUZ8
r4mwAGn35tG26IMMJ571ys5ommAIe/VSaoSobqv6loOif4lTZSMfL6AAJW08+50v
n+zMNJ85wXwBAyhO8qSu00Mndr50IkJRV+uyVKR59MfFisuXmVUzJy27lPzAGfPN
4t2H3XEjSNCMU0StrSWgJoF/RpbnkyoRNInqlqyOMaJ+i0V1jDVn661qGfEjGpA5
+TFpTzxx3GMbzI5QIbr7rMyUTKFiaIuRhP8+le7RtA52DtU+wusacnRVlNcys8lp
LuV+z3DkmjaakJudYdrPGAhb3YDpbxOcsqDv2ixPDJWDgDYKTS3b1zwQxzzghStm
vnB4j14uLS5O6JAxRJsXKoPlTawjjesCUwj9hR5mzldELBPrL91dr/Y8+jrJINzB
XTNGTBV95sHxMEEWmz46gFw+cmYfjQrtG3DqnluB1bhVUZUhrQGmiFFSsphA9ocF
bVRNq6YbZoKbYtIywPfBcsntLY2mavzlESu95FgskGDPKHpd0L19HlidzIxONALn
XAHCJUizfAvy+fIHhEYm0dWTgFfMk4qEmTA6kCG6DZ6T78v80uodfxJf8Cr/t1xy
iStOS0D0mypfwroClbsFzczn92PZB0zxlYfNe2gx1o6XjfethBE7MzHxkEIGGtPE
dV85qyLy5ihZVFzkY3P9pU2ffAtxseLe6+6TtkE7z0YTfIpMkxmHI31eFfazNqlg
ClCHpROnymIvwV4tQc903QFJbT9uuLjz5I1IKYizu0nJU3DmfJzvhwEXxn9yFGeo
xvVfVD0CVd2Mz9Rexr+vauqmuAtjcIxn2EJGCNHZnjRfEth2/LkZ14TcugGQlWW4
VSt6QpgGRBKECPUaSRL99+rUVQsX98BscwokIxV09bnBxe2Jh1FYMGhTFbNKxyv0
XIrWsL7HJDst0Zhr4QqVHt0nWnRhQPzAtordWuzPmRX0MVaj04BryDPbgDiCPvFV
VSadMIVUjNcdoNCL/Sn2xUZ7ITjd7gjtgzNrRWaDCqyv7W5dM5/RBrYv9/aZ1MfT
PfrFPzXxdqllrusc4I+/DR76ulk+hXu343JCAF14W5x2l9g8aWLpaiUKej/PgMq5
jIJfWC6sbXlfj5JP8ZpuV/nuyKBz3VTBiyupZQv41EKp6faoU5uAEtqJv14ULK/j
OnSQ/Q2rUkcbm/oUCKJHk1ClAs4QgJK8bXMjsdxcddosqLL9PWfVl6FNnpLOzZxo
MMYcPT6VQ8djQ144Z7PjmkmyCzphUgL+pVEhOOsvY7Ds6U8LLQmXUL3qyZ/bK7LV
Be8YdDCvWessRF+BuR95m4Ht4WwYPoJtIRhzLWb0UWuiQmUIbPVqOR3p7HbFFOJH
bNXUJIAcnrfIeKGN4C0aHvg8t+jSQTO+Y8qplPvTyvA+Hqqm/Ktp1R28tsDuvvFL
NAbvA0RHnU3FnReyX2G3csUZA9YoVrgCpCo9uGPqK6uy+tWdTu0qyUHdfOfsIqHG
7UMkNjiOvbsvbh4gxj6/TQl8O8bnhq9Cp72iuoshzWF65dd8qnch4xtpyaPMkqIY
xtzcScsnGLzBq1ULpfIbfqEVbvICypkE1yi+VPOxPUNJ8v05SsCszLvJx7HNU38S
+dtpQVsFdsndww0/UG/8bs51wk2A+Ftsj08G/sKucJrVLOHlkPpqXAYZyb6ASj2S
Trne06hvvcOpW4HezLBtiIw21VPRB1QA5IeEgJ4tqw737yCxqhBg+V1PPxDMsQC5
5qnSKgg4bfvfl5oK/zoPkojC3H164OyiLEX74PsBY7S7j7iNa/oSV4X0GHpspWbv
hwCH2rr5ko0X3NlU+qB5vANX/1R5+R4gqvOdvQFEjZ851KrX3/wQSX/i6e0ixA94
I2bI3u6lOqKa2l53S7O9NcgSs+iN9sr4suddE8aOCEVVz3MJ3F9um/l7twP7mHnW
WRivx9sF8Cx6lOirnubvzQEqXiZhwMpNGgH2Nb7pHsHiDb7HiLN5MWdYSJqT3Mf7
2m/zBSIylSRlP7tYB9uZ3bkrZHUN/yA3J5Xk+zvUpC5OnegnNGppIYsxv/A+hdjO
x1Q55/MZyu90yqp6OncGhNKDSanw3TtlRF6Qg0Bihvlz5wR9R1/Sx1fkOGfywTQ8
/+Ue+mOB9Sglwvf3pfevQxqyFApnyzAm9Z6aHiX4G1crdOzlMPf48VuxN+Ib079K
7W172IEYaiy55lLG25q9VUxMUeRBFxxzdREUdyI+mx99vuWudGib4o5fBjwscLrB
wHe8cMqDd6sJQk2x7HwajVwGw1sdpMKJmXGuepcQValLgRX/urcu6OLnJBF5Shcf
FPV3j7gsrpd1t/sxnHE5SAiOpZADXrFeChRF1NRTN4bBuywtpy5PS/T/wmDWXT8m
AUro1GFeUpK/1StUHtAw5pgx2EindakUMFU/KyWcwj575G88/9x0Oo7vcoBDQadf
+U3MAtn7446oGYtW9yLrV8HV4tKJP7amOkTli7TUsTMbfpY/fnoOG2Az13bS8sL1
T6ejDQo7kpef9RAs9XgDuDCDKKBU+LYHpvseySKKsefGzgy4nQ/rXDNMXezXsYO4
rAO3VCyfQC90lh0YgGgJfp103zxpjOTQ7gCRdQYisWlsOf5Y601YpmGCXdl99L6m
gbhT+tLIy6fdFc4UeD+OWB9KZ7nV4QVTLdEk0fgISsGEthorbiuYumOP6j2bT350
X23EQeA7wAJ7NTg3GXWNH1JbfZU1MzNBy6NUMEZHU2dPp22hTxhlnuVWwDJuP/m/
c1P90N06oIJDVWJx5zd7iBREjLqDoXvjo7Ae6I0evXaF53zqgkY07K4QiCpBqkLQ
VLFlCnHYxf46b9ivOzKBEpZc3BIWdietfNwSwvTJgK8Odrmi85WLBARfh6aEb/I9
OUIJ0l5CY8y6QS0t8MW0cKCc5aGfnNBMDudyHFXROSJW5I/nDmtGgq5bpyUm9a7u
jgtzoCThAJvdSI9rkVDg2XFbx/9WgLtfbMqmIsvcEDy0owSvrXb7/3k58+EsPjrh
9B/v1xG7rFf/w5p2sCvbbX4/EGFC1s4uytcwpTW0pjI0I/+Snqonvnl7VZ7xPCGK
ZdhyOtePET/kVMx7dBm5ssP49f3u7ow9KbH1VbpiRW7IW5ZeEXhafjDFGnAQwg09
/TgNRCN4WDNRIyaUdfzbVbNzxIZ8SbgB1K3LX0DoY3P9uTgPzHIZnjSak1XUdH7+
TupybsXY7GMuR0ddOGsrRdS22SjEaJ4207gGAJdngcgdLWiw9vfBAv3XlV6h2DFG
QP4wXjvihM9eGa5Crz/Rr9cumrSoMyCjjI2AvZGzijfjEWHOWaBZitxE+rAGKvar
jf5iDkMIJHwJN3HjJhWRFfrbP0qbmLaqCQc7GHPR2t9+y+k0KtmBSrgbG7Li5Rag
IJjVK/qh4I8pgeK3ZT284fc0S1VeLk7uJSNiirWUdBGP7JszI9HX8r68LNt+y0oG
y+BKE2vnMhNXphG5nq241FRLjRH4/dshGweD3P9X/7a3nUujqeUBOwlG6m8liEbj
5JwF5cu7d+74vQoepKb9hZMSUIj2V7rzV9QgEUL+nuRU66gqwQZ7UOoOwWw4Xbiz
bGnMIYiHy9nYRG4ViVtnSAhjHCizj9E0V71GkpBI1JX1/PKb8Y2ZtxCmga50lq+u
ZXlOiCw9vvxpd5p5ZGFYTg4W2g/ONFdrBIAvmnxXRzqxnk5aixpkfo3H28X0BrTB
qzhlUGAt6ofKNWmUbpwhygIat7B50CXSd4Oh67As56hENgSTPcwPsi1eu8aNdMd9
X0NeLvXH3luwiU0jILsAe0IuiaArkT60JLTnsLArovkK9Xu0OypBCcMFlfpUczpA
XDh2Lu+gjS3x62nDtmx40DtdJNW1gnMt/5MfYghVDLLLkLtfXeMx/Fx8Z37uNIcT
yLLBHhXh/HiHTSrutvpqGHhwi+8I4QlEEKXjKBi6ouxwk76dBZLegYvbTSSFXXLO
Hr5VHWmEJXdUjBH+01h8YJlilURhpbh0pLlceUV48p0+izNB0oja154qDzYQaNmJ
H87lFuz5g/3HQqWMVja/r9A6BkxxDBR3Zas4trfn9emUOwe2q22eLxGOV9Jj8vwM
LuIFDyN8HO5P/H9/05WrqYPTUgBHy6OjS+NzDIOn3uWUIh6OZthozCyxIXoVBhJc
Z+QUwVuhTjI+SOcu316VxDPif65Vup/2ZmE7+ziybWbNwkd01EXyuGrmLIPbB1Yx
i+Dt/PzqbvFGpOQ/FcE47G538G/nbSC672UxZrMNw6sBC5uEVUUgmrDgVqiRnaJc
QfvYbZuoyUnCaE+MK38vH9c8IMYMqgjPxwnD6u35bs8nARs1NblsH9PjJcZ4PZL0
b+ak8Ar/L4vuKlnX5WJR1zf4fuqwYEO9z7BrLa+9tPl/YInsJnOZB1z+8nAgkhwC
OobSBmHaV84FGfcbtBbAzM0a+mBLbsMJbX07X3y1JtWDcDk/YyiU5WMjrUoA45rF
1OWbTzflfpxepn7LDg7HkmnJtSWnl69oDxvmeUIrJE7FPUdaU45+EUBS5a9qRb0q
93d5RPfooePIpeAI6GZ/pclwSVFvk5ed6ElAxEzjNk6vdl4hKNEKOWNUPsKD5L/U
UvV+ENmD48yNlnP5I1S8Z/IGMH9wGAdTsEjLx07jFtX4T2XLUsuCFxeyB4S/Gh6V
y0c+dNorDQLJ8qxoz98qiRWRm6Dg3Inv5cLAQGXFEnmG4gLcvIZTvbVj4OFcLlPw
hAKqxIsnIiiEmAPSB5z+xTx78/nHPtpDES3ocmwC5iX4GWfBkWj5vXnxPdTGRzOb
AOd3NdiXPKvTpSxQ5l4cwE6wk+3+Vu5Q2PugPuuYXMLStTsuzyJNsXSLXFklgbN5
8Z8LchAnC/K/WN0Fi/FyI0xK3w1IoSoLJ5xLZ4fUFLEUwo83VKnn29q0+mZMtFDo
fl+6LOF0Zc1J9gwgjo1TOivEBOusD6CZ1ZZzTS140p55RBvO8T8ew8Pdy9NFcE93
mDsabS459mTdltOwNGAllM2pRsqg8go3Pl9GgIUJg2+tH6R75c2HRCH6rA3OPQXu
suudHOvQohWSh6bQgbWNHROCogauaPaOk+FkZNNRXXYZJcpGMlhKmrYn9GggjfzM
ckQy32gbCBZYwm0talainRKASIVXrsNpBmbTAAtO0aL7QRX+HpTdwTraoj12C68O
ARuXTTv5M3auVZ6yBr7f5TPOsnJfi2K3CEQ9Y/yll6C1fOBHM5+GeItklSZC9fcq
+iZl3wPRTb3lYRxhvKG7Og88Tq3Zz8WFyD1zZuEMx5VEv7RmWWQDPoUG8u+F0TGi
ojWu6hbBQhZZwOk6eLwNYifyIe0ueyHvr5X971R/m7zsmdJORoorzjEQIbKEz96p
aydAHQdsN2xAmAoudP5tLyMQnoChchuogH479NgyPAQmwf9yMmhVMdb3HLaK5Qi4
uMqVUB2ELQAWBKQdxmX8u7927Fa79JflnP/lS8ufCykNWcZU0TxA2zLHLpO2aHoc
D4nBOQKhFkk/KgjD0KHUBP3/7Zs6GgEI5ZbK0uWlng3Tk5av5L5fvi8rv8CrHv9P
p3bpWKMQKRneoNlwzpaqWTT0OZypikupUMEasR2ttPLZZSEqUlbjWi/+QvmDpRxC
sYdLFQKwc4Bp/7DGzc8NElCad5KvC+4w0JlAbY0KeYy7yMdfoe+DX3MIamscTQYG
LVkLDMOh8PggilSB6m9XiR4XN20n6Pf9JFbR760AJVyYQYGL/YGy2amisy502DSj
F8UAU3RxwgMZE0Vh61vWZg45Si9VEYosOXUElhRnLFobxm1W+D7HWI3gRj2nrbYr
KeTinXmWNGmyr7v0lkqjtWibABNG/LQfOs1LReL4ckefz18MkLNC7hM/x5hUI009
enKUh8HSv7Q/ngHOr9kby60rVHgm9bF+xZfnOx+w6Zuop/sLAOPiuH2zngVvVubO
0kfjZV1z1YHBIaVUbz0i7BpfRD4K04U4nB5L5QpKPwCQ6Z+UsJ6pfKMlNI0jlXRw
FHMOb6fKmvoi6gqqCo7E2xoZ9DD8CLbQ71espYIMPj0vaJDsnbg4DxdiJ/ZDfo9T
4/B1isGd1ZaAW6d5CabSosFDq3oTqZu8nKsqedTnoQ8LWJ7z8mg7mm+R3IdWrSXM
NV+XZWBsrCi7vZazbtdHIGufm5D9x/cHUEP64Eu4Az+OHFKA+kj1pYogqs4MuQyr
VNf4vbY3rIdjIFTSgpXArM62zBRYXXiGBsvagzIl6tK/CLHTMtv9t+BsijNNsUoa
ODwitntCiFoK2jDT0gCClHJKhejj0bY+XU8KsHHMSEH+rKqAypF9fnO70kXNyGwa
aUAGCxa7RRZo8/iuWcrBJQ5Y8EM/cQCKHvmqaKvz8wuBpTQcSXni/WrC6OfximXr
g/0zPU8fniR+Zju/OcWeq+EYTOFgJ/QPjmMviSJ/3PkThfNasBgDTzrIuAYGa5lC
OZtSbrXSwqMD0FlWIMALbWtbqVw0dwYuW3qUPHfzEzO2pUripltMXScaIHb7wutY
QNXHvfUBNe0TFrpvq27mF0VdXZufdw21dOmWpynIATEk3QpBF97xF39t4N9IU0hq
ryRihIs9FpWuQDg+HvRrCDo8ZGJc7zMNT5t7XRa5ETDuBSCYu0g7kb4MH4srmLQk
ChVe2zcdHwnGaZ0q6ckqL0ZUMMBzaVq8Vf2qnQKR9jv26p4LdV+uJ3ot7PG66mBD
QCrPrtUcY0IK2YSLdoDe/bcQJkDR0rlz3mhirdfC1a7IZJAalhYoK5VmAXr2wRdx
croJPKUrguy9BsohhoSQvf0FxkXcTLnoeTutTLA2V4P0cDT0w4/Wi6oBdNxVSWPM
daydTqlJHiufSwd1LH+rG69+WBqZiQYGje5RjYoE3z9MiT/s9u3II3UkOtWjCARL
3HDJkB2UTE58B85urNdpvc1yn7oxHoGVDFm9uNSS2si3ipN7VH2n7wcmDAaYEDP9
E79JpkNiMx/n3NBIOouiryu1YY3RrI0AMFiINf9Oz4osfn3ut8sDp3P7wtHDzA1/
1aOIRQ5/doLYp887l5oKDGEeFWOhJdPTdwhPbHeljNtmeRCx3Vbj4SSY/J9Lu12U
A7eJPVYK73JqA1MFQkjGvIZv5BQR7nUY/HKqtm4gJqf6EEbrC7F7tyZnlRANNIVA
iFTyJonzMpvHrkNUXCdUBRKcD30V6Brh9tShbFSDxgbMkdnmVKfSJm8Yy4KMVBEL
iXJ606IvrewE/u3w00eK1T34XFo+ECGfK/911dGssiPKp10GYNPYPD3K4YBZpokN
weEjihV7qKwgqSqtjkxjEcKmVWBwsu/4Qlpx8kyXy3fxr+WIid6QcggzDNiKATO1
in3H3JH059MOhOs2jGZdZf9ReLbbAjpRx8wXhYxYPCtj/j2h8gxSeTZIxfZJUoan
7AexAMj3NxBJT+tSBnpH/glydR7clnaChbxS92wbTFoGQTHR/C+hPcurpCuwRgjX
TuAjcxlVk3cPrvPmVYVooS8OnWx1JGym+NLaxlGgTFP8ojmoIS/5vOE7aNObKQGg
9GLJqh5eoCyn1O4yC/3m5RY7DsPsvosc2VX270e3uIU+yWaFrSei4ZA+z/b9IH+z
jrxVeH5MwQ9P9TrhCdHHMRMMyGzokTmlFQ1eAt7baGXmTjTeVksGIFkwbSlCn5yG
pt1OllPlr/uFXd5GvCA/k+ry1REZBYyj4FNSMa61r5jEIfoIUwerb5PaSDTXwjm8
+txsWDlk7JKquE+BgRly0GE1BPJfLOkaNdso4uMJ/jHG4YPrUlGgdcNrbSHLxJiB
iDtN/R9OrpoCCuOcNGTPMbq6f0U7rch5EZahKyzazqFPbq+I1qaunCbRpaLiqxNG
uFlcFMeIVzFQjneWs2OCUhWAQ9moPSKZOt/KTMTLs8LMTjW0Nkv+ygYxy0+M97dF
FqkbY/PVJro2d/vbww0+10gFRBeWtYrvXmkzmzqYlr/CTqjrYV9S5+yqIo2SKk65
T9RB7kW4D4qBbT/Z6yluiYDZFp2geTyrCjXQxOider/aWvGaoevL0gGfei6ZiR0W
LPu6b5zhbW6V4py6vvzdJiEnv4eVuKsofYTIZ/tazudrCyZAvDWwv+GWt8J1iPHH
VuhaeEaqOwKBNGhcA4WFfNBVXZNQz4JXroBJRi9u8R8VizuvGVr0DYzG2pM5unHs
NyccXaehpcWg4gLWARbLmvU86SVB4pwIBMrYJFCShU6oLy5g1MER6Mp5gr3MgVON
fSAgOoZbf79kjGx70TEF8VoYS7DqgDw8xuiP/vJloQUyeMYVZDLDFF7BJ+Hjx3e8
8dCDYMaOTi123DxNw51WXN5r2mcan6szLggbkc/DAWeO2MZ1XPnUOWIbIP6wSaTt
MvnTfb2Zd5rvphD6tkWD4s+2XBbl/PJ8gADJRRWcdIqO8lGw4rP2Jsg9M/y+eU9h
5WVrYC0jFuYnUAeDzfc9Z70LcjyMZnTMaXmIr9LG6X9OaWVRaMGL4OZa4t42wonX
8yEh7zzqRO3z/cmOH9KHimKylNqRFwvgOZUODc9lFGLvutZyz1Kv0/NBbi+SajjB
eOPCWVeBsTIK4dVLv78KP/MT93S/zxhM+EL/aBXJxLUHxkEnq7TczacwRu1dFSui
Z9wnfelffOUo3CWXvFfIymRGE20dOvJycuWj7Xn4A7ZsSMmxBu2vAHDRHDsGeJMQ
5RufjK3wgvetRSI4t3EGLBwwI9j4doOLeb17vcMaAeb4JMCBgHeunQg7ntAjTxct
ULPwAcD39WwpUb7H1Cw0x7AdvGXzxmXHooFHccjI+ZogI1/QlIHgGKk/Z088hOaa
Wdve/euBzoF+EXdDhVf72AID5gVVxgVIYm3hTkHQkQgGuVinIabnR3ELw31V42xu
yCvJOpJg0YkchyEb+0gbtbNLeNzeVHQCpqiYnLm5SVT3toTeOZOumj7tQR57Deby
/51R2w+BA08SnqvxZDogbdsP6DRxbene86zPGNi79hF82GiVmWQnREi6YL8Pa4M0
bJh5CjpJ/Znq56yMv3Rvw2x7fUPvtFtMykAqCXMzhlo5Y1utOG5jAsttQxGzRFs2
QyRG7g8/qB5O8599TRH2IyzeMmJGgZjn/t3SwVC7D1NCP86mYIRNF4o6GpGsLJHJ
z7UYi5FC1cEpGyCEGsfy8GJn4DGRcdVEyg47SQ6koGI/L1w98GBsqx68xJPBzxdC
5iWcUyBa/HqTANjcldc43klekf1F5OM3Vx9A6Jtqtz/xmIdmwRipjKDWkhucAj9+
bVXrVUrclB5T/nh8uiU96t0P0Qbmxa5jxJ/s1+tJWEjSxUnrqNd04c19/ZT4exs+
KgsyDQ35Dqvy6c/ejP6xMITYdvCU6KpAY3ZCLHJ/ItObUkznpEHzjr5jWcpTWK1J
lk/5J8HtzLSfyPwZYt1Cd93VYUtZt7ymMCEnAu9gQv+nsNQ4Z6csLqmYwKiBt4Sx
oNjBY82qKes2fB+tPExUnBjMXoMun0gstXNU+VVmjfEa0MXdHi/OqHapxBy0ytLh
7f1lRMN5X3wZqkp5AvRpjbUZlin3UfJknnXDOSvuWHVOe96O1WwmZXQ9VXmxMQTH
yRpxfs71k4wgnhFskho+IG2TVRprgbH4NiOw5Kq73Y7DFxt3gmpCKaUOhPQ1lag9
toRhSup8/d8qT5TSdD1/4ixwS9XozGvN7zT0Ig7JO0MYoACOf3dz0UZ6IAlOEZXN
0jVUVpuu+nFj8gEl0En4v1xtOZ8sTXY6Nzz08MzWqKGymcZAwSP3/8I091MhdeJV
Zdb6Xumii+lsmPU+Mk+YGpZoz+92dzjVNDmlRaRwpupSgjOJlP3NtxnPRQ7lmlLO
2J9xXd7XagB6SaxsQDXl+c8j9WPHcTM+d/oGyHDQ60JbFFwvhyCM17sEhGQX8Hjp
3tJfDpYJ+PGrWNxk4jf8/UhtKgYBXrWpggc8LcsxIuQvyxSclaIVYlEWyo07qnlw
3THobyKaNyIMhOjPnp0Yc4gvvdKR0B22EIjMiSeowW0DnM3LbGlJke2cvrhxfaY6
W4AM46atSR1jO6E5Ui9/2296wozuWs6WYfDqMtBIdYKKY7yqN/2zNljt/JqvHusF
ZcRe4LHEDopKXOMeXgk4/qg40wbuws0ccMs9Srhf5zDjkrL0AfmpM+uS75huYebs
QSPvzIhzWXRU7ESdVrssvO3Up1UfJQs8iLQnFdCzoJmqwc52n5SmdGmCL7gdpSG/
2q9FHrVtxTHqIzn3kPCUQGlBvSV49aBmLrxnWR8up9ox6Cgs6rZMidPYRgOo6ivP
mpOQbhwio2QUm6b+oPJ8g+0lBlSfpzfMIcrasGB1/qp53d3vCHMBqfO9kccsWSBc
w3j28+47CGPbgdcBKH9ivdE9+cIi5E5ry0Y8BAa3ms/EljwYbsn8xs/BTFQJYY+v
QsPCwPl2zNZ5Jg7t5oYK/y6Vx3D2t6yfZ+D8rshPi15+u4C9w8rL23/Aq+dZDWt0
QTY3Tkz3ZGE1NHkw6hyI542MuUguR0jT+SG2YUnfHM6oZtOPv97hxSYdG0ds72Fo
+E3XFODCnXn/kXJvXR8Ov2eDjA72bhooW/ycksPYu5X6Ql1qu4mgoVjMh74u+rj6
Q565Ehk6UkprMcIbyYJ60rbcFf8lzl8eLweUVgW9PBLJL9AZmH+5mMPZ+ORTOR0s
5Gfuz7dtyyGHMnLXwY6D6GNIR3HPLNFUV3n2jj7CYH/byqV/uentY49GDhOPUkdv
FGIkb8fWJsxLWN409MfGDkgh992cScYAKPwedNBXEDjLjqGv0t+8fLhtYGgL3Erw
V5ahaQocsnNrOn5767/mp5N09BE7FKIK/T/896aezspxJg2JqaKGbO9zhX1dye8U
g37/OW47bdqZL/gnJQrg4o3KcGPdX+gz4BTLyXDK1rIxGBQ/hUH3fw067rbkXi3K
2UTSmtEAxUFKlwHEiZlPFdu86DEf0F8GT698s98co8oHV6ClvzVDNDdLER1TV2M8
SvsP72ZP+esS9SvYk3P/SJGr/cRS0KBDO0DHFA5Fo7BvvorpQEYNXeA6B0mnmIff
/lLenLyAgp1KpouOpM0YsfKraYT6M1m4QOO3QQnU64LAg+9BNzPLE/VPzYmoa8Jd
hKxJ8leGR/WzpvhkWlYR27DJV7NpArsIwPBtd7P682r6u10EQTltU8RJvSs/2SFR
zhBSuQzz2XDtSsGlvE0Y9kd7TEkYGXnDv+ObxBOyDSU31sIJCk3Yrwj5lzBZ/syN
g1fStpxPyY2XT9j5DtXYIcluJ0GtXiYh+MR6gMxpqIPxRRDXx+/yYB0paKzMXMAn
6FmzK4ZVobXp83T7ouNuGXL+y1XZp34xwXG0/rCGe5b8FSMF3vnA7JWONzMpyMK4
/yxC6qNPxyuaP3zs3F1TGNGhqIoRWcU/wln5m8bt7DAw66Id7uawqndc1Fo8bPiP
qUYZFI906WEFcI2EGj+KIsQyHH1BCvWmpFmzs+htEEuMy2pyc2eD4q/QLDiKUblw
ljZZGtssp8nMAZB6AkblwYsgde24i5/nev73PAT+UQfDLUtK1jgnQj0au2kCjZ48
jlUr4Vng3sVnBAcovkZqAwKYZg5HxkbUoCcsCa/5Wi2uI+GHbXObWW4/MgXPdE8B
+pPV41tHI9yFMLGJWsZYuKW3H5JpOFDVsmhK8zRqGeVdHN4a4qNIGAG3/iAz0/9v
TqSU8qFpAcU6j2W+JreFFeH9PHYi5T8jhIR6+kWPLaXU0u0/MgqLfdSDfzZ8B+6I
Wq1++Pi13j1L6u36WaNKqwQOY+IYTzt4tBHbxbyoMYWP50jCX/Jer/wtVA5Lk9ZZ
nkWmShogDURYAINcpbUCjHBdrXgTNWl7fCMzLwwFBiXPOjf2qW3XO9o0ZD5+BoGW
5PFdDcxTx5AiQTc3RmD4ejMrDVBdL3kGvqRK54hym7N2PO+i+3WS9iQbzTh/wbh8
FHBeMnqb/+HHIJ4gZf0vHR8ZLtqpXfZUEeR6WFbIqEDEu2046NtQStwjJUdy1FeG
HOACqCml2TxX6nbfmfcm2QsSPUtHNqVgh1rIsWb6OBk8uaAYCHqn4QlBD/8qyztv
1i67WfVL88vx7hfzdJitDcrIBzwQtVzFN0M3fffaAGijG6wwCaHfE1TATgLFenM4
ZerK0QDuoee6CsBZg1OfBouZ1l1auOFAOqx2SXkjMfCtd3o5HUyb/APv5GuLQMhZ
XDyOBDHw2nxMeSToHRCeMDWUZhwsHuLPImuQB124Q8IDIELVlOVAopP7TKzJ7xXS
du4LuH46cP86iSFeQR63F3m7zLZK/Wr8k53UZpS4ESRZBAKzI+FdjwXQAUXMJXN6
6Ffd6w6I0sJTvpGfpB54kPC85eUo5FNlks5SQwbfPYJwBmzl7LeXOc9bz81J147O
igDZM/hJJRE0iD5hfuQ4rU31X+VnCHJ+zSJK0KNY8iJb8fVp/s7j7gtkqj3xPn4b
tJhszgAO60M3OX7ZzhBzkOyzemagMGp9UrvC4Htep4n4sSahxWbaS3iXmT7g4CsY
Z5fp7qphC1Cm4N4K1R9Ki/8006BNHR+jkuZmtMl12p/HOsh2J4/L+kUAhyHabFjv
H3pT3SOIwVTCaX/6OCr/1j1ChqOLWXo44gAa+hiocpnfyti6CUuZXCv7X8dO8Zxe
WFjxK4mrg7aPchjLwkB2vb5RcF2+AKxczadSduQjUZL9x+XA5Z+K0t0+b2NPVSGc
CQfA6t09FXRiJv4C5bdk0oHEd8nbL79CEvGoIjfaz9+fanQ856zZsWUVien+L0zz
ni/txYGBer3bbkI3TCHeBDjoDW6PzwSRcszekVENTa9benfQUs3R6p3Rkka6cH9y
gNpV5jztCS42OOdeh/PCGWSUjndSVGRN6mE9Ykt9/UcJZNuMu4SxwpVsy1sW3CTZ
HhC/G0sFCvhdKpr/ltIeTzEbWeAn1YVwfdZ9+t+m+6DlmQPniP1A/6b7ophi+Eep
T/MzTsCO6cTe0fp+B63L5c9mWDoXL1xZqxzMk8AoT86yrBV5d52GpGiDwtQbu6+J
vXy39+fApbhwT4K2hwes74I+em1dWfqceLhWzlnjnp69ov71ZD0foyzZZvfDMw+t
/5sLdoJTyJ+8L3gcco70DpLuk3VILGSL98+KP/kPA3enLxY0UCOx4QwXaE68JBv8
Ug7tCF/0bU4z6Li2OXrwtF1ErwPHyOJl9kBd23rZ8rckKw6+XGSD9S//EVV9JrN0
qk79mqiMeaDoKMp6x+xvcTa2QApQZmTrJEUlX79WisiWLzgaynY/RIfFF8PJtiAL
KFeEjI3JA6nrwqcGfg+sI6Hd7tSwDRshonop9nuGLqidkWNEZ37HdXXR/uUWbgyg
WCicL2WKGYzOqF+uc+/2/VZOXr+Zn8T684UfyJyvu5ETo6b+B8quT7LrnZUWk/VN
BsraH3hM9rTnpTJtM8HodhGaa2NHP824xyKFk6rzruDvHTkgcC1ONnhS6UUw7MKr
4qJZLM1mb7Rws7Xj487MohxH17Ax9XWfvngVnmhJcegjfhE3mv11IAYtXw+txOO3
cw1vmezx67IjH2XOV0Lx6ZUBF09kcGxUc4GjHa6JNbG58JKFeCTznwuqh+Z1ABMN
BijUxk7DrRlgDBemCpAF7kl0NgOBLHdYCCWfJgPPnNrb5pMMls92ByCMnhOruMSV
LwVh1mT3W2/fbzp+AS35yXTVuSprgwoDecVvlRWPZBcAmabsQNl5SqDkPGjIYolb
o6aY2bdLRoCJV9pmv/+tz3R/tbcTaNdGBa6/sckWu4gT8sClMXAmexeGJN0hgkZp
FVvNX2MBkJbhhnpvLVtVP9KD0TpXHMj8On23cZALVagPp7gI19BDE+eUqpmHlyxy
lN9dwIsWs/mIqVkokcUth/l/gHZ9EzQyRA/wIM4zu91pfCqJzCHIlLNqiq2/qkt2
ReUhhQ3E9z4hWFqGB9D80M5G+ojbXgqpmCinZDKZYXYFrtKmrWX2yVNnpcICGoKc
rYo1OLSHO9PtTOeWNFQv7NsJuOLOvZCqvKh90jzxf4/SsThl6X2/uBD1Mj/Gu4m5
aF4rrPAb+VHiVgC9d4BdS9fU1m774PGu8vJs0f2wxboGEQccJWup42wUU0yS2HMJ
dL/D7nEajVFyRmxjdSygVcHO0R3C9DAd4tDDTFUheM7Wqi0dgcgIA+uGCfEtEeDz
lvCdIinunE72WjEdNusrM/ikztLUfh0fI+T45pviaH0Abjuh86XD13v7alR7C7Dd
UuQ5POp8bKnsccGu9vwAiA9aMCBb54kedGv0+81HuakUdVNVLdFy+vuupJ26+fyH
HlFovEg9t55TJg9gYMzDkfbKxjmpFQkHoXI/jxKxc4sTyDh3xQQRdt2a4895rQ5e
+04DPtcoU+7l3fFBX5hGZ/TCBCAwnhLX5ZNVnDWlWf+WaRj3PTm1jNEffc8X+bmE
/BYTVMbA4CQ6gyh7HmoY74IQsyXzNW8kTbSn/vX+IoFVztL4Cnqhfi/IUVoqNIUh
7EBOGTOtclEBvtEd7jSpirDEDMidANaEARZe2u+RhqJH9fA3SPbFBR6lsJAbOuZ8
4A/pE8Llq+Jv8Win3YsdJZ53zAmxZ1B8p1J6eiYnEdYnGL5TLvZxQq6Vi+SWRAoe
vd/7BnqGeLsq0AQA7Nen02/iZY5fwwPBmJMhaW9NCOQ9r2WgOlNqIYAwl+yeRdCN
US1nrjqJOh2lazEXkRjpWfhlyYeB9HeiL1FgM0/nN6kXmezjAxw0/dmFEt0manIA
35dlD5TwIRoY6/NtN2+ATpV2hn4n5s3GaoyywUGxodHl1D79SSnI2mlW0g5Mly/6
UTEuCdfZHPl/302qp32Vl6pmKDh0UghJgI4vQp5FS63xGv9yAz12k9vVVAheX/CN
FJDfdAmyAw5oKcKu9yN4RVjtTTjZANhI3QgalwbvKQ//K/xvNg0VodpWNiU9wUPr
LudG+Pz+7DpNVLc9Q2vdtILEKNhm1RmJJNOx5LJ8irMZxH1XwCXVHf29IALv5lAn
uETKFJMQzhvnil/Hh0w6xiZjfMp71B28rjcfjGHYklw5gNDTiDXOfibjFcyQL4U7
Dp9OrEOY8zmdx+FnGOzumrrs18Ju8ff3yNK0T8tCRnT5N5XdMwmOkLoM2xm5OBCn
8FBEyPqGT45nqZEGrQ89ZVU7Mmg/x5AZpvwKg1sb2KPFxtuT7iDL3mIat5ZW+AIf
Se+20+/s+CTNZB3Zj7CRk9IcHqsxBwIsXWFHkCtRj9K08jZAO+71z4lZ36z+u2vX
xM2eiNuF7yfdnh5FqMPS4fGgXzCtz9DxR+pZlNNWdZ8VSZ9oKKymTcOPvddrtLcv
v3sNHACinFmCA4HMsvvG9vdIw38JKUwAfw6xtCk6Gf2uH51NZDP0pix9HA+twVh2
84gVJaDzCKhZowScmgxLL9qwi7A7yK6CvnPuhvvRzpwgv3XsDhCxlZsLLf+9iwdK
jDAiG4i9Jbk5AF9fkeLJpMI8G7+vkUwvI9Evpqe23QZhuNkit31Na0qWDWHOUznf
v5mq5vb+OmSWEGBwGs/7zR49LRYmPmYKGJcwX13WspwtEi3DG7eNx5RXJVeLFY2d
7OaDIsZl7OhO0xkYhfxU7e7vaD2UgeNC+H/cqGzM7jh1T6E4sDCtXVur29Z4eT5Y
9v6eyWNEfFZa7ilp+6RtwrodbT+oEIHg72ey45NCtzPorO7lLgWNCPnyjyA3hFQ+
L/HWkhZjDc4/NY/f26nPGxyWSGUmtbjJ+7E1Wfo0Q4bETslkzwf3bM3qmRi+XCKi
kTrpjfTzyL82p4hzZ8XgL61gw66nJXtQrT79jZU1olfyxz1zhIYcCZVVj5BcKnPL
Z13HoRJAhbSFsPyIU9oXspSHBHiXBHye1eWsEuUT0lHGjYk41FSh+HnyVCXNtQsj
FTy08il0LjzBUIvOE3UTC3UB+8zti/b5yCWR+2prrWHahM1hXUkBhQAocXsoP/ek
mOUUz+AqXZpV33mM/0xRDrrjj2np/mpsFbCXDCByIyaaOxDqxgC+WDdop5TrNHG1
0EfKYy5T5xmL4ful7ABRu9YbG3rH6Ref5usHc22xcnd6aguUu7ckCVbFrerXiGqM
AhJqbMR0Q1oNKRARDQDUzxJmoUJaAQ9O22p8wcyWp3m1M1rI0rqaaeJJW5iMVgaN
edaQiuKK9fmBT9Cx/hW1DGPi2kV/GUmAoRI+frhKXL5TLzod0OLeXW1Om4iY7IVl
y+DC2/bl/opEgSIm6dnEgzL2U8lGavFdcL2HHgq2KkLn5ZKtOFtqu1D9R4qZHzqV
hwsD/j0lJATjaojBwPM4z52xyRB7yubRWthVnCfHfclXOnOVQzEtbxRTtkEvEIOJ
ypqFrdbL1MaLwydXOqJMkvj6ejBdiH31aIHE7YRooLc9F/GDnPhKOzOQAE2dQHZ1
B0CqRCh1PZf2StywK5IEjyRLyq4o2LTGBKiT+QsFeBz29cDX/j0RH5XccCIQHUYW
ZS2tpC1rGwSIyJvqjiS8xV7uTpfUyK6Lg13WILGLguMkVprc6X1PxJTRMYqP2E8h
lduAVdEFIfEZKSHjhSYZoecaPsyOm7IrMNe19AfVuwIO5Q7YwOARdyHk2DoxklaF
u73j9LtXmO2h7wVDDmrf1L0wTJb0mlOO+5JA6x9MKNrBmjOeGr1yi2THH09nMYNG
hwYWvgl/4vW1Ra+1Jx1GlhqJENlgSmmrHSkr0ZZw18XuzQ7DdG2ztagkHItbfGI3
6v9VGXVIaeJuqyR/4Sla7KyK2ye/IZD9RlclB966S/br34At+w4yVXfxBg80bR+D
bYoegdJ/hYEOIT1ue7T9u/gGXea3gBl1rgFFjrJbWI9JZ7H2aVJ7N5mO2R7BQpKc
zLjrRiVUbfjFi2vToaMiNm6Pq0nsAhjr/PVM8R5xHUxZV1VYM8bk7v4kH2/U8V1f
ZPCKHfhVLXvTlZgSKu0AxKx+vLghpvCmEJiG/0j47nnOIxY2qHkeHChgggFuSs9i
Gp1CuvO6JNL1+dY64F0HXpduqXEOhKJluneLsqiBJ7dE39Tzj/rsf+YsHwu7RPQH
MXC/hmD9HhKFXjpU5T39It66Lgb+9crw2mtFssDMuFr/QrxI30unvHfcewWnbSbb
nWNjNCmeCmc/5AvRIDGZsFK9iOtIzPt5zUUv+c01V5YUmO1TrnBIfFn61z27qfCS
TKiTlw7lAWcWfaBMYQvJvNVc+zRFwLViCov9JrlGC1FmyNnFsmS8uEx5YHcaG+np
UGFB98GOigo1xufoaisg7Sj9SH2oGy86wz/IpmRBj4cflG6ioZSyHxbDKmdWIdk8
nK+7RhjU5S6bbt2tZ6cAkJzc/bwuJfNgEjbb/N8UWF3Nk73OAHReidpCClrsfxg3
On5Zvf9ParoCpp9HtUnetKvnLtpXBACamqxnS4s58j4zToyKJRrsI0fA33M5d5So
nZQetWXUHMiYJEfKMKGu6IzYzY2MAAr1XgKmz0W/7WY8PmULXX1RT2l3BfM6OmVn
+2VH5bwHsUjGq8olpLq6M1Kc/M4ghANMwSz/ApmqAgOJl4hzmbk96aAN7i3NwHkU
pzmGwiVdF16KIPOIVNg4lYSljk2zGhrSbBDehljTpR8nOIKEiaRjIAjkfAl1Om+p
tEssfTzW6HwSvSd1Do8ZKHAv73g9MBMBD3tT9XqYzA7CZZPaTFfh4IkQoNZliLma
WHFhJkCcArgLgh22+xKo4iIpgn9/Ap+5BiUbCkx79u01SaiEIqc2KiTpUxkCQhSF
iAG4H4i0MK2wVnfYTc+Ele20fA9SrceJW+aGzS/X6H+PYk5qCnl7YjIJe852cqPy
MXObUG0CqGhmIUa8GalrB/UOgvqqrn97qCkmIadEYAs1+H1fcNqLk9wDiIpHI0Wy
uk6vuw50I3CIavC/v0f+GVUPVVVdcTVX1RJRWt2VdqnLRltEWs3eDZGnG+gxpmNk
x/t70JwQt+SvJw8A63a0G+7JDAyBioKXGqlK/BQiBat1d/b4oAkCxRafwMlk6RzP
zSsvqmxylLqoZSkLPJPYZD/cOXMTTw+Eb0fYIogRUbIo+M1vHtelzxMGUyU99BhS
qoJjR3Kxpk5wntRpoN0jy1ggp4A+zEa6CvbRQDzG/DmFGTd0WdO18J6FjaiApilm
S62AtFYoA28oLKFBjosV8JWeS1UiVXLx8V1GFT1UsxpBQ1n5H+HM8ppD1z/8fFyF
Kl32YZY2J4mQ94klchl+LxFO4cqkOQmJEENoM83nHkvYAtOj6AYjG9nVK4WUhGCK
cQc/nSJAuuQGVmLnXzkeJHxMI4/6qJcovrQQNoDAr5NbBG3Pg6+WXyEPVlwO526T
oElptT5PrCK8pPeak/ESY5DcI0J8oy85C5uaetZJXbZUY2rsTUbjmGddkc4UXb5O
9euAx47IgOgfD22yn1Jx5+Y1jrN3JvnfD36qKLUc4ItaXkWLDuVxoJZfDeuMhZBX
uhRITiIrWhDjXBGoC+MdZi7PJ3dLWu6a459/NVnrn7yl3A1excAJQTs5HvowhE9G
qNWqo97DMY4muoX+2qrSrgOayjIisIsU8JzpAAkp1Un0MtuZ5EVrrMxigxmGbOYB
a77+Bqhi16NJhckL+TUNGh+/XwUrdZ2/Vxow71d87zZrmcgLedjBH2EqdpRvO2me
GkWuYNd5sub+8bHiWa5z/p1pZGaVnvCDI9MmzA7mO56BRs96H7rBq805Lz8mtdgG
f+s1YPkiaBLZRAHEO7ArrHpzjjT8PSpYLqM8XIXevAAkTjeubz8BfwBRFbGh5q4q
H7xO5vdKJ1kocDdZnmNagxfsLv+TeNAIV+sm5kkTcilG8RJe1WGWxIhv9NGun9UR
EoPvDGqP4/vQg7LXPKhnaK+R3farOElHfDK+2neiDQzE9tmU85wZdEdMxukX76a8
TRLPsTy5dYlt+xql4WVBk+PAXMtXanxqdywK71qKxd/DMhE77/Fnol5WhrXG7w4Y
CYFBb0B5xaxtu1CSwkQpzvutcRjQh6Jzvz53c5vmuNSluuonA5udxqUi3nD8XHIx
PgIM7cYZ2mjC1d160ZHukglS8OXyMAkqNxe95S3K1NVhAgIiNCwMNr1xrjfj9x9k
SLGmaua8x/d5NldtWK0NQtmXlPt7G/+HYUGZbMOJPUh/yXL15K537We8Taj0go7v
SEwF7Cnqz7wcCi4rX/SvnbNTnb2k3Ng4Es6yla6FVxh5eEfHmxu+e8UE0VsQAz7F
uYUEOU8uZ+WSJv69jcbNEe/ajdBB73VNVy3NL0cfnF8lsBYgx6Eryup3asMQU1Nz
v8t4u6WiVznA/ExRPPo6Oix3wgS4VH1rYM/IaP3y3h1DzC6rxAnxH6h0O3Y02Nrf
nGfKrHaUldzUr9skHuFxiKAQuZs9Y58VEn2XWeimteGBv1QzbyLJdQ5wTS36q7MZ
PnyVZklkGdIzYP2NOrhYisBGp2rtGCZ4Voch/s/9Zkc+822QeWEkvoaTxhiR6yy0
daISsiqJ4qI2QgD1eDlQWfpNepMRKB45OjhOS/Q1DuIqynDuiRsIG1lBplP3D/+F
yfGy9KV9Ph3ZvvIrVZmGK/QbPBg8eXWY6wqGOOSgQiI/72QH9wjsJuDKvYbzODl/
zduEJWQhCD8ITOH/6CAlTun8+qwxR9DAtRF1ZOrsYmneW6GbGuLHdCZ5NwtnAel/
WdzCLCuQusVWW5AYQZ9WXw+9jnzmo0QLn6ZteXc7dy/271lqL322I/gHAGWRcCmn
xRU2eKcgTaNb1FpTgpqYt9mC/sh0qpkzU7wATm/DIMyzrDae+iFKB0XJiKZhd2vn
yI6oh//kkE37JUun94ZvF/jVIzpnfgqSDNbABdpjDLzW/Toe3Q9eDA1zqYE/pwyM
0Ip4PU/fsJ/5HWKfFWYroefg8wd+LiJeF1u0zE+oNweEnfeMkf1qllnAwukgySaY
YP3GvGaNuM71rdInhOV2bGST2aIxewwDTGLYUEWqQqFSMDlt57OppW2wdldelFq8
EkYCJhSKvN4AFiTnJDqE+lFE4JPALG9gkWU0rlhcYsxXK5LdemjDglb5i4pmHF/O
SAj5CBQxoiL2PlVGStKRB91Iq9OWHp8JHdwRGyTusThPmnnnMjQzsgzVpjt/cZuz
R8gI2Cy9d/Pb3nMOOXoIp8A0L1rRB+XCLbwk4cm0E2y8R1M4FiXvu9BdS6LNnNpr
WMvx3Xr4Ctah3G6bD/8Z/N8ARvTAmE3A6o/GruYfTKpUwXq9yXKQaB35bY0OceXw
4JkTS1VFf8DBddAFpnk1Ryj7dfPMVHwObjx9Um+2CrIWQ+acFoIFKVuFzCew0Crf
kh6g820IeYHpdnkWDdBZxk0MwTk2Q/GgzjhliCNuGaIvrRG8gT7ZWy0U1uVllkad
NzIj7v8FzourVe5LRkn4KdNm7c7F8ThgfNKSfW25gBSargZfac8mtjV1mbr8tDcU
sRYRX0FFjd5Zh2Cb5Yoxu/UOJxW+OaTQX+K+IM94/oUhcx0NxnwL7N6/Bi/qwZHn
BVbPFA2l/dXW+loWh8wu1UCKtLI42EErvA31Q95K5EOF+Lp9SvNBYNiq116U4BI0
i1RvuYy/1hDTg1MfFSHHfxEmKpRonedIap7mJCO2k/gNkmw7GIRQYyrlnomL4QtJ
NzyEHWWrW4WVRWOFbxVm2EeRIPhESYii2gplOTfCozsCjcdz6FRaq2MnKstjM9SW
0yJzxYd1GXAQ+gOahO7USafwO4QavnKnPOm13S9SEj8=
`pragma protect end_protected
