// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
dVlWNfAMdmGWLpm/YLdAp9AZEcDOCUzCrBWHLo7PuqgV8GeIvZefqDSxvAkFgloMzV9KGgHFA9fK
ssBzT3EI5zuHEfyreaIHqXuXB2avuUUMK8x/gEg+tUOgIU25trVg2967nB/sdusy04XiGtUgDsHo
5WoYVn7wwRW+SUMgN60M5Uq/xH/K11KDiLM1clq85Lgkkzuky7+6doBDwjJGBThswsWTzhT9SMOv
3AjeqvSM8o8jp5ISPwf3vfQAAks5ePOc2djCwZjVfdk5lLUmN2QHjQemmzBP9P7CbgwPc+pv1p2I
ICojbffaUtQ+vny4b23jz1yb/+lpVq6ivg1iaA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 45008)
J9CiQsXXIAplc2huV5Cj7PGToFmd0iXq9HbuNIrx4N/W4gdhoxXW/owqLcCtuQ+wUi4WzPfNmdDS
6STAKP7I9TGjSuZWUoyQtn4adFFC/Mb+zzy2afoE4Gh+TIJgF/1a386K78qpynkzVX6flJQn3ZzE
IDSNv7uFREkcXNrdpkoxTX10mXCeArsINvjo5Q5Mnd+VHNiIzLYoGv53SFwkJRMuvNyLiKhu4P4l
P1SKZpEhT/1fCufLM/WggC+FIohTKgZpGZUhfBlGUBQelURTAlx5zKSE+22Jjsk0Lkz7XGPi7xcW
lBhDzbWbtZsQM6nKfvIVVX7xbp018lEFmLmc91Dyh9BHljgL38yQDTyug/xk4GNYeAyJ9ctj8oJF
oRDWykdGpnkokkVazgoPghH2HVOIkYj5JlkDB6v1yQ9y2S69JAJ4pOgRM2gOrkEcjAu63iinveRk
FtXUxSpAS/dG3aeg+D8jZFN/DX5onHejcaVoIk5lk6CJzYzc4ZGgsBlFEr+q8Pc4eTspJxh/gY00
me+/3fEyBRYTMJsf5sDA5IvzzljZFBb9upI0+PpOoy88XoeMXNTP0pQAD1qdPL7nOkyM5MDoR+OK
gtsBsKMW6gKhlOBwo0PuyYSlCuLp3weRERm1GCg5sLtnOR3qZnqz1AFO4bzKDd8qH0yl5vWKUpAY
MkhmMwS+A7r7ZTAA6GtW25uph9JsWFECgvT+0eA13GnhLp/sBvDvxpB+uj076pCCgoTdM629hEdn
jduFZx2YgeiJtW07ruK3xLlBpJ8arRJtQL0dTvRAVdotAIvLcPDj9yas85clRHV4Wx58tCUQxA3c
Y87EOQK430zBo6TGnHvuhatBIiAqt5cWKwJXJvDM/QaG0IIWcEwweLNsOs9mjQjhn81C0NjYIxU+
ynt+fGzjJ4JVwIgQ+EJcE2SfzCDP4KHU4jRgr1hj0frNmij3OC56q7cAmkKFu7Qaq+sZw7za6QUu
Nx1W4XQQpYO7OBliTvGM/7snH3qkvJxrpGaznPX+lNxNaxPlnMpAfxiWh74TIsE33f9T3VBKKhI2
kyHI4SwkW760ShbBsH3hMIGT1lWtNejyMtzJ5pUdhqxse0V7xniYANIU5TdWLzwQukbMNV9PCuLa
5sdmZhEu/KVwg5ouwrbga7dVhLU8S31fpO/fNpgIrGPwlDUf9Xlcco2pyiMP+EsLJ1t/UmsrKyCq
xFfavNb/d3wj5M6BntDIJyhaDDMigz0hXbXvCi7wsg1GGwEE8O3RgBDmucbX751hilu4MZo5z/So
m5lB/LuOh/fyRhtExGx/iUr+TQTtfjD88Xviln0lsUta08tIVaEhEczGfCZ30UfQSqbuS7jApZiN
rJZM7RKrH3etlqixWs2Kk+UnJD9o77eh1Gg4GWfQ36ywk/T/wAzMfxoRLuAz6Y28KLRJ+J6fd5Qv
9DiQo9f0DVYl0Zf1EzErzT6fM/ncW9ONO51SVZTe/kemzJOnKOFb2dAs833hGc70lt1x20y1hzkY
TxQMfwEoGelQV3jJYr30X3jjxhBBWZ6QJaxukSZHQ5k+G9SYc44Uk+kLiDo3EFdCO2ryUrzyXwqo
RmdSoahnvPZ43KP4UEOPmS2PolBxRzh9wGGLpCyCYHt21grbThG3F4B0chJtotJNykzQCteIH1hY
RHViNQ0AdN1W/pgygfFzXf23FenaVkbfO6scuAXU5xoPx7fwoed9TS89+KAVYWBM0Gx/UDqrLsNE
l5yKANU37rBqYC//uNPtKhTmZx9Rrh/y62dI1i57YHHmUSUR7U0844Cb1IHq6uaqpt+JJeAAJ3GY
JjFy6kWQpP9RnrIKksdI62uwXpdprTHCdvkZuIvGuE8rOICF0tKgH0YDxNYW///Hv1K+T2Swo4Gb
FrCcgC54o17Zp/nD3H0bWNnQ1Jlh+ERf4ot9NH93PN5L703GwcigQPWWT1+dxIg3UPf9dUHvUALS
R7z02QhTktXoOw7pZ7kSMwaSBp8YvXeu81r5bG7t4XWJErG3jL+OW2hf4J9eCN19rO5Ifo6Q1zjM
EfaSJKzsFu9s0L1C1qfaHbAb7abKjnHFjU2QD6+v0+Gv2uitq27D2sKNaRvSSyhkq5Gu0bHFSY6R
z3fFPuqm+2yQOa54F1q43jecjsojYZgiV2F5PJsMxbk29FWXy1qxt/QasSh+TC5zSh4JuSBZ12qd
t34ZgshqFWx5e2HjwAK7FJ0N9ryftBJvzGlwCgkRGsKapDMDjr70nj4tdceiHJ8+wZlcxrjc+ikg
BftKiG453B+HKOAjHngCgn0gYgl1MjvgtOxt1xEBTlGEx5BLDv6jdYcb0KJUqZ2SE3RQE7IUk+gT
vm9tWHhIt4MrCQyOA4I3Wr+vy591Dm4Qjl34+bKb8/uTMaIYNku8Fe5ufWlEq5rePpVNFb2yFBrw
LFLZmfovoCNw6ifHCWiO0CCuxEwIL1UMahUJpLhIOHhju5/rDKtovWc7+j3/QL5aEJzgrbekWt3C
ZpS53siVXcHRxYHTLJojFcitXPPgFr8BbELziNIMI6kHYyeRbiaK4ZNl57b4muMGpvlpEc29yMV3
0J1bvt5zsEI8J4JlwWV02OOJQpe3ep29NtWqzcRscUsqysxy5P4Zinv4qneEtGM+DdFPm+FHjd4N
1SIu1dXGcx0X9LcYSp4cKaugk9ottJDJPa/VZTLaBvbNXA99w7emlrtlwh8CHwNpJIU78206e/9A
aHqVTKcis3nEs29EAebqpsOKgCQyDnmMpNWh+bAg64OqqprScKiZ+KiU2NzagYVd75/g0TLodpai
mwKTLL7eyonukrFzKh63mPFO2/4DQteUVr5r7wjPl6oxL2k8K6kQQDp2nRAGeTYlHSshnuplY9X5
qqQ+Z1hJeunbtt2dHVoci0o15Ug2nnhFV9RUwNTjwdBemTu+KO7qv8JL3qWZyxS8uTD0HYCbGf+5
W3xtu4fFa15UYvivfvu19M78vOT/3B31np4Y6DVzzhWGtLvzdr9NNtz97TuV4Q9b0G0I4bYZgJYk
Nq/zYlpBg8HsjZDUmUoIBVjSxjWGEIt58vEX9b7g0HHBzp+MrETg8rlTxZ5IRf9cRvhPgGPpkbOs
jhn3QLFLCf7pJ01tPQmh78an3HmuAKtbPukpQa3Nbxwc9Yea82UGnM5wOorB7ZlMd1qNzepA/lI3
hF2WxuZ/u8HGJe6I15lRmdQEB/+1N3sMPug2megsgQUVMvo+hNplY9gT69mw5r1fntQOOJ+pkcMG
EUUauSw3YLB2uNXcjr9msIXCNn2CwiTTJIVaskokAY+lC4fWnHf4oV0t0E3GJZ2Y46ZFnd+OWgXX
le2xx1aNXW9dCuANVB3WGiJS5Cpib9kSebBXZ2c/gfGmgkMkzcBQOqgiabKm4MNPGTaM9JKW3GOl
B8Q/9rIK13eIzi4GaIEoFbRfA8jdXp+xE8g0hlbSj3zZUHErLCAdFssLl3RJPxwbalo6yVGHhPrk
AHy/UOCVC8oE0bpXYwnluElykjv6+DR8npfprsKaSXDUFtVPlkziRGHie9ng1ZfaikRCbRaKkUWN
oN6o+Jd8O8iiipyNrBKnikORD7l6W2mSnTleG+lZvKeklxV2EcON0368qojHwZiv2VpcJhGjpa73
WTXp1arz28Dv1onUsMVO2uExcTFJ7ZNEcBaUSFfeS1ynFnpjAArfX9Tbo+TO9ty59xIGG0HmGLKQ
enx0pd8SqDTffNi0pKG2zeomlOgflm9BTEofpVSQdbN9p7DbkL5hNIDvz0gNyDfqolE+Ai4EFCvb
JMsVGk1rqRW48KdF+DXuepoqMJVwQhNcKiZ0J+pbwjfqTbQx+9Zt2LlqC8Bhtjm/hCD08+JXJGcN
rq18zoCkIktpvmwEVsHYoCmUrEq/2b+xBPGYP+CFCiY0FhMfaz4XUWD1zXLuAUzXIPvbcD69NzSk
sM+0CUrnrp2kxqU0S5U0ZGITVvEl9GzXs0YiVQ8SNo8YSL960qdrpxt9yytnuF5cqwvY5aQOcecz
E/tQGtd9k923bJAZ0M8OM2S32DTqrvkZbAhnkaZLePZKVabSyoTKjFwT1i8KHDl2gTxlpey939R1
FCbJX3rUUfB+pkuSm84e+gKEol1+iG8GgO05840gSPGIgx8/kPc82rwrhbzPj+a3EngjMcL0Hcip
R4SjsFqPFlaCUZBR9vXI+D9jGZzki88pMUv5m+e53SNpHYYuGy542lSULHA+iQ0CsbKVTg6v5fbd
XSVEjP28bNGcxeM/CunUjVpurf/qfYvzrSdAtkOf1j7C/31KjOwvwxQz9c1NDttQ25Wk4FvsP2tn
05YMtErGw3pQKmCGXtE3v6Dezrr3NSLcvkHbfY7zuupL4xe7Q3X9Y6GBbgMuR5z5tRtpMiGw5ktp
iXQUVeoT3Zws4MBhbMWwm733w9EGaE81mpow0kPmNSzvUlhJnwrf/YAD7L4UK1wUPG91h69xPKu2
PidRvOzDA5JkGwmFCSU+yp/LxF9l03WM5eLQp0GfmuswULIIfADhgaKQQ0WqT33NtBgw36DkBS+p
DmGZeu0yd47RniNU9+btcSAAZh2SO64zfgj8eZ6q+wqiwcuJVJsb77w5w9Z3Nm/dEuPLyOyOzlVe
KO+LDuva1UDZwPj9EaOA4uaMZyIrKFsnmAhtRoKa7VXWvL/PJI5y8ZJA/sde61mijZ4qGM3l/9Ji
rD7tco2T3Ub81myFAyeyLqEfphyf556CjNlyZ1B1W6izCc4grEoVF3ZgDTjKvv7mOGWhimUWdVSK
Afha+K9J0kqBlcXmZN8p4jQOZ2rpv+8dZHB2cAegYs8wmjn8eaRNUiIBZWPGGXg5zUDKmqxX6vBJ
qhwNvvC4y8pAu3dzIHibRpnagiitEgnnQeK9Q3B3nTKqPJHPsp1tljngT5TZbHUnTzb74y0lA3z4
SE2AbYH1n8Ly7pfouf8wqmPsx902I8JYOrH/Wa1ab2m08EQy1h/waBJZCno9yWSAnUiE43lCRgVr
Ja+wTWnNcXRpz1EiMdg5cwQy0M82HyV+36f8zLHhUVePfDb+IcSibUFqxG/YbbWqWnXcKsWWw1Md
lkSDytxC29OP/yhgPNkRR7Cr0vZ8Hyjf8G2uNHYZbZHKuiMfAgS/6EERrTTZRbHeeDEYBsL4z6Ap
EQ48JHnD7gYmjGlqWQQLwPej4VghucGscShLF3P5ke1Ajp4hE8pECpBFO43F1ZIASlq+RCUZBneX
ZulA9yKdP0u8FYLrqvasvD/67R9y1NRm+Hp1Worgxr7Q4s0OUIZjtJgJnnPZJPFbxVv/fTCB2JLl
DAA+JgbzFsUZn7RnlGHcxXZRzTkaIKdaRrM9H5yYAIcH/L/87RgQUkGR3IFXRB0XfIeNAshPZxCv
Fei873i43I8FIORmPRmGkjLQ6rJOpkMPu3Rje8nfrhkqRSEHBNXw05zDjezYBwTV+ss1JA4o/roW
/HS0Gvm5tEnQxxHaYYHx/09w8BYgTLJBPebhYKnWQBSfGAxnbD5utNduZOJ4pAbhFHyLv3egNJVI
nmkw6cCdlFcVb3ZDzLMyhTvjusnJh9pya9MhtvBAk5jqcwToJ+q9RqgvDjUKmEukBhxg9ntTudsn
OlAWmyij3BaUSdQ8z1EjaSryi+ddXdCxGUZ1mp8QnnO3OhphBkjOCOqFq7UpSNJUIQmV7Gd604zD
Xc6nkmHlQf8wRNzZ9BrLQ16h0POIhDssm9Ifizdcb8sw7z0uuRZciSUviLwfYrTR9/h1O57CP30U
LbmB4ns52zVF8maR9Y5dPRa6T4wpDLLqVOCnYWG94kCHAoQ7e3CbmFAq4aPhL3scpVmGKMdY/zZq
kjEFPeyBqAgXFvw4xAVOxFPoVOu7uhdGVyKX4y7yduRdiR7xQIISuppNzwWWUzwI1TXAV1mcsGPt
2Zf1snhLtZzRAyTt5XRFeIe5YqtWXflH99PK14/FCx5wHXnC15SBbCNm9BCR0uPZRmaBtVvlcklw
5Tc3651oJ9fBGCaqSzugiUvZNtEldJ+bM3HOmks6E0XY0MzDQxg+0kefC/ukLsHYt8wvJ8QcWd7t
dxL0O0i59oINcQQmI7UjNbsYvy8O9roCglRMd9i1mILQRWe32uCUa1qE8mDPznJ1Fp8eNwjL1Hmz
gRRORTABNUvCR2A1swEFfhaoISfO9F50mPKQHNDb5sPX045EKAbfOR/xzxJfbH3Zyb7auyQ2rQeQ
xJ59XVU6G2J960sFt2jSh+O+EK9DqzfCOE5ieBk0Wu6B33mQC+yEmSuqzMFYliVvGEvIMdCfoZCM
qV0+mAS1emgbHTQUvFaf0jUTeCxAUwjyusV/OshzCnyHQTDCFbhFcAWuy2CbTuPtdx70E9+uqYV+
zqA1Ty3dy1NgKrDbPGWTR5f53wj9jA2JDFyfVALD9i5tsp/LIf+dKNgS32PiAcDg1LScthezh2Kj
w3oLkosChIBZmFOQZqwCP7lbxnw5GLyVCUGR0TlsciFK5VazJ6xYBhqleJsShXQ9tyx5EVeEBdtE
Aq+UPEpNr8HH5W5SMGI1lSv/6lfiRbsw06Z650Cq6BBCvjNfZhy7qyX089KIBuJMNywKhiIrFOON
JtuSYlqas55dPDsLEFEO3vIDq6LXXZ/OJKaZDPf0HWt6id8qQmqNIQjkdQleUkWgWe0qwNcFGNCH
k2OLj3IY/6x/tLqWdNFmf0mhGhmUtZNWjmqR0ms7Tw3lXKWwD+xvOeNoJzd7/BEUwJHRIgY2j4IO
WVXOqZhhGCwCXJRKEM2Wzel+gxntduikavJ/AFZjr+9ECTwRdSoaFPKDNxnhLi6S3W2RzM5XkUbe
KolxqCKNq1xfXMjpWB2R4Y+aCb71NVNlsjR82fidVCHjy6PhlKjVg+HK+/r5TB+gskWpRRpmcdNy
mMIJlmCc9me11u/jnpic1Fxt1fiwHqyufsrJhvPnyk8mOP/Mpt3dvBXf7WQXAt/uBQ4l2OAO++Ae
XKQXgOjS69RyBMhRLVSBCVyZLFrWyK8uhNhMin1TUmNkLQR8oC7sXqAZD2KezVsKSMZ1CynTwbkH
I8eMNXlkkp+BtKbX1WXsi7fHQLsWlF+jQwwIkgysWP6n3UOj8biOlcK9aVn5aa2HBbcQD74wbJsC
RkMJA/ZP9M0TrjAkXR8oEPrGOcJxLbPKR3IOEPft1Jz31tkAzR1uUl5nZ0F8JTs473Ua/Sv1Al9Q
HrhMHCc8dIK/cfTNRw+JW46lha6onO1cvgObqjN2KDVZ1OurYLcN36Yj0tdVIpwAjAe5+aDQc4tY
QKJhfIvmVKOmISlPDjNPsHnRa/bTqUrysyN7kcuuBPyTbotlRqcOKb1d+iYS/D8cix9zWmAeRlzM
e2I1du0WYrl39RsOhm66+BZCfxqeul5x5TkYo6LrdFdySv1vE8AsL6lWxI3CbOveygTi9G4BwSM/
MMyZWJ0XXHnWAkPWUCZvGr3XVl5phRaL2e7+8no0wIXvqFiEmCCkQyZxF6ceohf59cxJCVV7DXtT
u6Gy6wWj3vkvAg4F2esr5Ju2IlU/sRkJYQAnyJ3G8zx2EqFbkSBVAZTqWSUz3UzzjxZg4ZMAH2ZJ
qHBZrk3+aboky2cMPf1S+Ed4DSqN+KV7Q8aFtuoxd6Fj2TUS5OBMwmotMdEsHPrJcVHuvD8bv29u
rTCN/Io+uHm/a0eHSYlKklUWqYqGCx2+W7uTh2nenrHkypCSp2ET9qeS2OAB2m4yHPKfnDEmMiQ9
ms4KuJWPoaK+BvFcYtuPqlKLN1IPcGCHs3UR6uYHtkOatn8MjwFrRtV1WPob7ueBWQ4djD8Lb2k9
V/xQ1Nd/Y8I+XVcWsur03K1EV9qkeNj4mutBqxDkKu5by4jy2l3Id1+USm1ymzTXOMCbyXrLI0N9
h0fxfhKMpEcY8tr/gdbtavNIoSDNH8ysP+NdCO4LbMPHfi/xzQZ9iuopFuymZHZ1eJtJuvukXGvH
ENTsiuM8KDaOxDfBnEzj0xDRTmo/9WwQUrGOnhWlUS08MhUmGc0Z/yPQTXHuRiPjZy6Fip46Kmrw
7KRZuG3jKNTqj8jw+0rUf2gThQiy7EFySNvbcFykP4GL3gqSHxc+xttJryimwofSZJYJDc/WbAwe
ldwOkioV32af3g1FWe9eRiVwxITxlpreShpk4JCDKu5B6xSaP6G0Lo9p6g5q6ICKFDmSpNMNuGsp
d1yBmMdyu0JLH+uSeXR/hk85NP1qRdQuBlffJGRGHXVb4wlIOw527lsIiUYpj0SIIB4Oeg5WxVlj
Ttj20G3QlZDx3UHvXXUe1frdZD2DCpPmIMcz8fPnnxe3jVNSlYREIpY8O8h2srLLXv/gbrgUvA5k
nQQswwINE0ZCkUvR1bkoubf1nEMHna1ipHc0Miydw4TxoGC+NnHQUlt0v2ZWnCi8QR7G6o3dX1nz
ALDONLKqcB26QksAs0cKDvub2GzeYoOfMA7jwLgv4pPF64NeyxPIRXY3tSj2bl2itJWwQuQ2CBQ1
04x1yUVlotzL2C+PBWJzSuiRluLLkkxmglftraIcey4RqbRpcKb1wTEFOsmoYxLJJBb0SEh7chLS
w46xdqroT/HgzFbrFpaulYpa+Q/C4M2UByO8KjsZ3G6gBdeXPCrNV31FmpFT/RytmP24TW1yM/Q7
+G8TJe8RInfZcLaES8iERBZr1LesOQ3gMt0tAzoR9gMwB126voQFa3+br2pd7Zuq+WPxoSlBdUNo
ERG0ka3TSz+YB16dFJE5dNzq1TqfDvOSIFMCg9nkybhmR3BY/+XDItC1n5lf4Rctw/Ch7wDBG2Du
HEj+kd1vbGOJ1+mM4FSLfWbwNJNEEpK9gkp5RvweaqXImexcI+k33zlw1Y8c6ruShCmILYxaqyvs
5N1kz9jvMTkyEA77AeRgMT8xMC2QzM8O3PbJ6ig0n7Ie/ZVlWCFlLK+UBTg6gHCYYYbxrhBdB6d5
GbXJoRcgmz0rrV1mMiwLelOZR+DIGTIqiHfr2Cm1yvbZZd08ABvlKglueTMf2yEZ3BRtDrt5YgTb
0mpCYL50xJvoxbGlgpitgtVSXl5IANfXwlfs+borXLbiB9+mYLUclbkEqOtnGe8LJW4jryJDxZoQ
eH7XyoQaFcTDw4Cxlxsjs0p+HxYOXx0vLu1G/Bd3YFd+aFloobLG9rl1n91iSNAx2oqG45eh+N3O
SFhOvILKuJWtt5BUcxIu7CSHbnwLU2i6hkMtRVorECSDWrQaFqFDIAUs7WocHqJGo2qmXK1X5UHp
ziosv9l0zjNJXz0HzzYSwQLVF6BsFzB/33gRhiGsZuQKlIiPw6St0p23aKBcJL2E2udj14Vic1vQ
KHLL8Ya171AtorWYaYar+bQtMtvvGYyYdK8iLLYJrRTKEhSbK6xfZ2ylrlyrnUx1P5lrDbhSf8Zn
HesZbL+qZfibwzfSD/x9Hlr9uyvLPTi2hhTkL+QyJqnsm4V4OQyvWoR8R5vyrOEUiJKVtHtW2a0w
9zEKWLmPeEhg2SaKbSrSnVXFLceoL4Kykfj/H/mWZd4OlLVJTzwoDT+ayfNlk4xxzPCCFXsBisNx
rmsYf6Q2Mq/D25JyGKE4z8Mt5qTQ32rBQW81cVgoMwEptpnQ0D0DrzNxSJceBv0STlO1zjWjQ5de
2csvFvEefaogQWV7hvAjm9AT/PL63JjQqalGIXhmSUW9E5Om0rVzi0+/LAs4PT+4tz63lusenHrS
Jy+4KDRh2Iw/uI04GQ/JlONprw4gEGN994UwcPuHXCk2Z2lht+0kdSxbRJR/GPj2B8Mb/uSG6ykm
dVyn1Dcs4yemhC8lNuJv7wlghxPtFr+6Tpi6YPYy2VKd1ccBkqsMeUM0RvNuIvAcet8U9cDtek5+
clAMmjNfL+jSda57AHNDzb1BdUL8Zo3VHGrLrGFaV35odxJ6YUH45e65Strjr1uX6XAnv2Lpt80l
dkbpEuoeTUfl7D0BzIVPRNYebtRZIF0Cno/7Dg7HJkn9OxkxuvjK4ixNHITWXcg1GJs1ir01iNBw
O7ehvQlSRnxawMG+/QODcVBGhJM2GZtnwBPiXKVl6mWmNQd1szQGnFfiqGwEDXPd7mWCE3leOauF
fmphO04crOAY+BuFeOK3YeTMOEqyn2qMgb96iDCvJZp9WiCVBsyjgFPu9A7gQFeT11zOmMJhlaOk
No+TdGBS6a6nHemtKnKoIj1FrMRZrQaxrvRr3ZZGxspsyTHvLQQiQ+6Y+VShEJBj9541Kq8ruMro
py81uFUqYtDtpWR7txU7C/VtKT/ko657CF6em3eFxKdCr8Pg1fX+Mgaj8aB7wHKIWbnJCoiK2crh
bCG8Y1B+yGZshGGn7jm0iO361w7q3dALmAJvKpBxVCgLMEBl4NsyAjOna+CdB08Rdxp8jlfuaigv
Ohu+9fhjDgUOOgTXCjW61kDOxnhLfeqiZClV0G3g+QygVM2A97E4ZLtKPdhi/4s3VZZDqy/ypu3T
igfqkzAneL9b64wCk+BdefFyz3QcGKplVraB9BU21Uu2mfDGomyYk6eERcmQCcfVCZSEf/M2zYhK
uS3jDHJfyLxDrjVtKlN4qmwCAv+5g44rIsaGlmhtIbYcZ2OfeC1I0i7rgo7cLP/Np7DHKQsM4Hv1
8X21eaofQmKftgLaEykhjvSq82pPVIgrzQqfrWwP7OAfEZ1j+wUkKdgHkB0TLa5+kCH/YDp3aCT5
boZENiiS+PqGTBp/mFrxI634haLduXoL2opTjx4Xv+6qG+C/sp5lwoxe3gyYC2nEw3vOB66M5VPa
tRN+sxKA4CY2dm4yxY3c/pTih1oKtcd4zu0of3ZaZZ5qNEXvnjEO92krh5i8hit3OMIH7InvLhVq
XoaG/3gZZ8/HO6ONk7FrlhtmycyhjxdYnAXR/Pf9LmrDiuhangbbldlJFGFAuYeEhESGUwytO2Fn
S7ohZpm/WROFTcm7bLvYT/k/PfbbquFZ9ibxcstYYvxTLDsW2JZ3u9m+2mUV2kPWauCtQNWmlLfL
h7E1j/Bn80qIMGqzTrZ5Ri2YACZj4CqWwSX9DOH0ksj/Ssomcg0+ZC7b5DOKwZPQqmQAdYm4opUP
S6Fjcw1H1sM2oWx7pgYIOV+sdaareGQVNNPLUKfiedB2/QvZOVxWYS5msYaYNO54zZFL5PQnj+YM
Di57Fw3L3fjcq/7TlfUUL8aTN8GWj7yY89XMrmgXPYnn04ITOjMwGKsZYAPZ00wFVHdi8z6WKw+i
SxXpuhoT7vwiF8O4e35Dwi24/6YXdLc9bsEEf5TaFsXlGPoVIt2wWV1QonN8Uvicn4zO2AF07xOV
PzoxVOGQuTyonRcOAeWfuG+WNfmpbkbPPr6EVaIJVOzveFW2tOLehLK98iHQQzbJdsHbf6bbKCx+
BIQPZMd2BY+/cnB0CV5HQvhYG2rMYnPoW2Gpe0tEHQkKNmOMnxqtu4yy0gSZUoPxmwSzPNQSMqSq
hZ7QPK/wegzsEiFKgY18NR7+awSbVUDrNLAvzK9sPu5qwPOZQq6GB8lUatwxJtJ1JdGnW6hL9a3e
5N8EntXSNbSCJ1cSunYd5Vy4KHyTsjQpvOBe7iU0rxpBLnedA3D0jaRJV+oWEv2VTo/BCVYeNH62
83MqjzCCxBmie4M+Zv2A1/TTzpEOXBm6bkIDxn9YoTdI0MObRPrHjHr4P5DCxBcFi0KHw/bdt2J0
Qtm1G/FLrYHwXpShs2g3r6ln8pWxwHv5jHfkqMWQlcJ6tO/f9NZ+ofFrxSWr/d4jding0wxPNPwb
fmvGA50LVEQ7pHk3ZiY2vgFE4Gun+MYEOv2dyrsrPCosZ4z8dmVZm00uzX00KYl35lGbTOrWV06B
kNdU2LiHdMLFwT8yHWsDyv7O4Lf0JShg0akY1tr5Fvg9JUS++Wttkqog66tWiD6Tm6q86TZdSVLB
icrPPRcAFYkOUurvc7VB55xgruuORHYkZIqRVoxuIcXnxfbqYc5g+YhvY7XoCukEOiuKjWmeW3qi
n7PQRO583mPaJHmGkx7gyn6DtOH4P1ZQuzB1HPV/GOSaTR21sG21tVAfzWMg8nRBrHKjUQYoB0Up
D0Py5eW8G8OBrs4nL7BOBOOlTgMwTNUy+o3L4GFjLqrBJ2eDF6YclUBjbdl8xeCHloK4MASUJhPv
8BYNFEy+YeUMZZtfkLBoujUkpIRGuYjhaifbOGA/AyL35M0+dJanPPWQ91LLsVD1XsiAJkfAl0EC
21+6v8z7HpV8KQZCObiNxKK+LQgKiT306y1ukZugjZf6dQXGK3eJOAsK7uKa2vEmFDu1WiSVAPRm
AmgaxRj8XFrAD2ucpD+N7X5T3LkiwRGEJ9u3ePWtTmtH+Uwoj53SxqcwOxEkeJ2NxVrTr/h65rnq
QFn76PZkKOsjRpsXgt+mbAP95cZa01fm4XBxVn7gJm55ZVPVdr+KYRCgsBNoXtUrVu6pGA4BNl4Z
Z7rVTImwt2j9ZpzHIGS1fT0R1KdeA/sXnshWxZw1AH7jtbJ20KX0dbdNLCRCCwmw3qDcVBY3+Y8A
2a3fiOlggJaEUfCCIjeLd6R82yi5p7GhtdqbCw7jeU8HfA7uXE4gllWXz3YCmlrnl7uH8LvYQ0/P
+rnouueqIs8w+r0dvYyG0bo4JvpInwH+3HDF5djBnSc3UtXDqdhI5fLOpqKCSh3wVEvW5Vd0yaTJ
aom69dUpf/vEMiN6QHsNaCTcmGEEUYpjZCPumlPh6N2nKHZnZBR4zC50C2AIZoOI5CywG8ZC/5IK
0bDmSezmY+Z5tq435SvC3vMjPM0VB3TN8NN1gYbLiY4pk1L/zAvKTe7xtS7d1NfUZ1nFxKPuNjai
xu7zY9qSbh1RJ1tqoqvToyGC7rhZGaU0Pch7hVcAyaz40SiM19VjHIg8xqhgExMQ3yW0CZ8dFlb5
t24fTwa2ZSD4+RMENVQtClX6pljKfevnN9rjGFrH1cLCPsFPR1Sgd1gvpJdsyA3b42J4JuU3B9DK
BKTusVIDplg50QPsn+A/p3YD+YMKMuv/Ip8Kfrs+8Fq/CyhHIJdx/XHdQ238PV7oCDNFrcb0ZzC1
U23ghPuTUFkNvjqI8t/jDtugk0+aIYYzzVvrtSLt7+6kfRaiz3uTeUO0bWhvGD7P+62jjO1wciJ1
sVW0lDZIqKG2t8qGP8qG0slGsiz+aeYrpr5ryUB0NsY76UBP3SCZ3TfoQYqbMzTdYVxinqHHGarP
v4Xek9Q8xIGn70D9yuEpQlAeSQFgFWj+Q5trzG9cqha4F/KTdkRxpVaY3KiNkL9zUGggwqvGoayX
6hUXThh0uG5KAFNhWSCOmjn9lqQu54NBPsn/cNxmLriapy76LABZCBPjGRrr8b9tq2w77HTYk4ZX
LVSbHyfwofqq3VwFqtRw2AiT+gTSVcAF7KfK5kZ9tZrgFG2erCypn00B8ps82aE4SQwdoA0jpd2y
xkLImG/7Owy1HEeZizeGGG2bO1Y+AiWvJkb99pCd395jaQquCDETucYaYXhOhTYA/W8v6HQGGCyB
ZCiKijIox+shluCsKkorHydDsN4FtthNwcfEmDiX1IOpM8P6CWJapUknaxNLk3CkU5BuGYQ7gGuG
z3LyVB3HR8MGAXf0HN/oRBMIw4Xx/Ye6dVOd0h6zusoxDX+AdSVdWSpnG0saQDZgPv7A2FRJvKHW
LfaROnd6Zvdc0M03KiNZOVthwZBgo102TNDCJ9ppALFOUGJSv/j5ks1nrnUuO2NwJsqRfNGXYLPG
ISzDyU3X/kvKYFuflbRTJsZ5axYqxaTpLWuEQODK2qgTbbp7NE/djYnfjrd1zTcNeIjeZL/CxkA7
+G7gNGBbQ83u8ZsxYICLRwrd5O7Z10v8c6Gy78JlGWbUGSi7D1GO7d+Dq5zetSc8ea473/fOLaE8
rduuw4tOxckR4PxtjpuEkXB+cxE3ocd5PO9bwQNgmEWRVTA05cRyD08JR6gk4+/mH8kH0x3loiYv
AcPu5QBzN7cW/GzOqZ/hSYtiDepn3bHuJi1uX7KxvUygGIS/TAWZfrxtBBgT+kkp7M7WSogOy2rM
reZoh6ZYLsSDSF/NLZrUVP7BXCTp6fjiJwjYxU+dS83uMGR5+KnsUNy4pzr/ZpKjS55NKPpZr44T
5Gi9hF3W2q4RPucgMKmCznTGJeWO/O8V8+AD9na0U2LfvuWeliNJlzigIf2Ic2+FTmgOxQHhFbWD
0Zl6MeT56rmBKu4vGMjD7DL2b91ILSP7h72FNzbIkelTK61YfVd0fqdtNXl6ZL1GLqOPOeQLG1l0
k1HyU4iYc5+kPa4eVwl3G0sbM5c9jawvWX5yyNsA1LZ7859nJ0i4D3+ncPlTZZsHsytn7UnSMMU1
WppbmhRPSwxsaJxxti2p8TVrnrbvmKuJH+Zr5nKCoaMUQWA2Cn+ipcd4HVz0gz9sfkfAl5aZt8cK
wvkM8c1DS6oGp3c7iZ3eQ01wwzeCWWZ0fqnE1JDPJnNH2uUrhQtUwthIhlONPB9YCrXCZXeqmBT/
lHBgjQ56fmRLZhX+4qlDmntA5J6woY9ZmRA4YTxpoMqafK2yzKrbEBNbT24tX1fOuO8nsu0Dc6Ua
kzqq29tEc4ki/Fr0EtzHt8K/s8Tvc+hQLZkAJFnghgnlfwGWk+XhhxQy9VG2EL0ZKCYKAdIbZukl
GVaQ4MISKuoB6x9Ha6EOdrBH7e1GfgoYTUkMBxb8IIaKKSDP//Fr6alwAmDVWuHZwP5pwi8TCDdN
JkESt7PT+sUQuzYqxABfwDWBr8OG6oq6xm2HhR0erO4POy5GKWW6/yskVWp1PPM0ofTeaCXNDM7d
sjyGcAfV4ALoudgwnvORMMHQjOM6B2O++mMJ7X3ht4+/2NmkU5PoRAerJdF9YTxNIrtBS/TncmT/
VLrw9QXh7YkZv/lE8GgrUB8wagZ+ABWqrg3ril4yiyIiIDX4BddqJvDiy7v19cZsKI0KAZwJRnJq
3VsPG9K8lrfPvnvUm4oKPynqq2UPukdRISio2iUi26R+WaN/eKCtER+ZkRLidhrOCl8FbR/70tuc
3qHjd+b+AC9rUtlhvPKPdyPcUdecIAUw/ch6OI50mi8Jgf581la9tYUPLR9nVik4/UWTZ4NdG0zP
0Sl+fhrXx1sxXtqS8pbUIxAHDOxvEA8TtyGpoLqAvz/ke77elzZnIc2tfUG41T4GJK9K/BRwQqWE
JQ4viNeUOwujglD38r0VPlgZ9Riz4lPMwxLIvSWVGeYHm1BkQsjW0xQdfITd2stG3ggXFDTeBY99
NOAjKB/W+Jm6SRKvT4nXc2cObaTQ2sYMpzZ9EtCMRkuol2GC4xIP9Jz3B7Qo/7K3xwq5X5TO6nxR
+qCirvFA3c80RiMNx9zX5O6nAZBk7WgHCBr8ZId7fLh/wspTtU0st8QWaMJ4loVGs7hvsLkQ34L3
J0dETI0Y0USwd2nnL3bxI1DsYgS/syPraC+jibY4T9nnZDqtlVk09De2yOSzsEjDji76tp8nXiTV
fG4IosoC7uIFqg+FBvnglmGay+HyvGjXaShBHiMiMtEhmNNvs23bPgPty1HO+TzKFAz2Bah4HaW2
/kV3DzCUJv0y5F7CLOJM4ieOIzLRmv7+MRnwmpoEkvCcIVu7qxEUsFs1fyIYc05BJNdozcHwUV1p
+hQ7u/zGnEFGVoq8VOCsVhOJuNan//B6AHT87yBRJWlGi+QfBK1YF3VruLOjNGGNHj5NO8vn6Ubu
RwsxocL0iHn8VJLGODXUl3/UKe2w8/Vrx3q2pOWfrDmXXm+ydlzm7vTWnrZ5tVCpUWsWP2VtbSTf
ZGl39BI5dLahBrd1xKnLUJI+rV+wLMWd3S3jJZ0mU6Ff+Exl62cTuSGvj9N3ch6UrbezOSj7fDm2
TT9Jhy0cBfuGcjROdgRL3m+JC+qZ37kKl1JxvY+atQ+stZY8vRAdhbS36RFUI2p+DvbjYPWfAJ7Y
ldILCdqsUgPaWwGspd7YReqyZAwGouSbhrhhDjdza68tR03D1sfSnTv8Cz/RTdljN2QYrO+f6nMH
ApKOdnC+jmqD0c8MH1Pn52qNA/082VG7/yLcP69mneK0peAtaoPc8tJPjUYGJHxPAVqNeDgizS4X
2xk6QJ0+3Xtih4ZjFkAouQmgaYppVSn4ZaCi64fcsLem9v6nYya0vjPL3GvVbFJ9L491d+LMvjDa
uJyj+XOSGdt78y5qv/iS1Nz/8F+lvsaMtvNcQg7L8TmQL+exdohELlTFdcrDQlhTcgcWQ/3bSSY0
uJVJYnLpuuLMg/644wCsrMpc8q5GdkzKz0T0i3WLKj3btp4ZgsU9uXTqSGPHahE1hjYKL65wmFWg
JEtkM2MKeLIUBA/7a+0X3lWWWm6SaEJgUsoSNqFfpmEU+YHk5usl/WCj6EPAVQcXVR8BpGgtoffs
dL+mqqlaQqfj7CH8fMiNiTKAN8tep7hZtKQ8yKUOBLOsPH8ZQUQ2a1PsKZC69OyoHxgzPs/Mgg1Z
250R1OMR9XGGd641+8WfThYmN+5kfdcWB1oCNB7iV1trN9KPsDeySwEzqbIPw4SlsRhotJeQHpbP
fC/85roYLtJdDY6HSXFCrChm6QJT2z7QA9UHoUD4BHGlv33ABeP/cCnaF54jy7VTMqJ6sWNleasu
EsFtEu2q+Nw/NuBTZHyrWtVpWx48WMZwn0Ex6Fqj0bVDaLsKaXJDBPwg5kW9hWgNorW5yWte22Au
oRvkZUqzwfCKkmtfI7hUJ6NoPCn7aAp9YrJmB3+Dm8svrhkMadvWSkrqPBvW9v5v9pPTL/lu+sCx
U/7r7uxFqrUnRtrp14D0MCc+GfFdTNXa9pkSyIbtMJm7kcM0NxjrV83DMr+ihCMvrPKDEIaOvD/n
xS2U0nioLqv6L7X0NME5P5jk+RJ9de8/30GqW/YHI0WD7vk3mND6euh/bueMaEuO5G4+znIO+fqd
+JqPThgxG0zLmfetTMCiByicC5CNtQ4QG/pX+Jl7qegc0ZbFlvC0At0nDZJE9KnJiEqn8qEs5zRi
aatJiJOKCaulyp4Wf1xbiLM3IUoMOib3D4yojZ/mW7xcfSUlLH9smXOE8FnX4UYEdA4IscRf1K+z
a0jomVCpkA+dNxPvdiIAAqyTyGVcyYAQXeFke8W54dnwiCKxCi9YxiWQNElNRXOHv87Hh6dLUm2q
5pFk3fpEfW/8ciws2nF/QmZb1Pc7olRJp5ge5wN2OADfh0jqnQv0Amgqg0i+yKPlmeItjZI1UWls
k+Wayu0Uqp392iXRzkrd4u0hIHXBKskPPUf3eqH0UUydnniu9ixCf11FMcjnL7yStDhFSzg0xFpQ
yS1yjXEbi/V74OK1xCqJ2gM3a5FJL1H5R3zl5PTiXJQQ8upT+0H4u+6lZVGcf2v+r2x5LWTJG86L
PmiSftXWnYSwPyVhoTcLgfuNDiiGadquf20fIDWP0QE8GvGCtxywWZKqLqsanCfboBYc4XkpHB/f
OiKBdkN3LqpwS/WWkE28TRUf3islNkQ5aWuqFysJBuujI21f+lpS6ppCBlOsJeK8OebWCNoZbHLs
L0HvG1gJtu9kNU1H/Vly00TObDpn5Nhs/SvJCXFOzRtq7270U6LzK/5arXnPFDayAfcGodLLkPr1
h78ppfvID0n+Tfj21Hu+vTspO5eos3A0oZa1pIWPvikTwFkqthGMRXT8G9MY9K0h2Dc7ZKEDDPmI
l0JGsPXvXk+hON5+CuTgSaCrQ6ozwnIiVvtBoAwGtaZrkmqt2m9ho9zUGWFxiOCNieoI2H4yPAZJ
l2698uPvzu5E7W/Q9xialqpXrxNsPKQkiCk+q7wsxVs4mBtRKKN3XZ70K2rCmz7t/5CkbjYrw9ZX
4SnUNt2voNKq9/FqtaAJtYd/tUF6HxvaQ/3Xv2fhzb8luSoA222sJft3OBDoyOhGnj3HRuPIN796
NttwqYVDNGIIvGUBM+BDyHuZBTPLWRiv6DZzktkSiqEg0RUsEaOKfS63mJndS8uePNVy3qks9+AQ
VWbeht/rBpzbZDmQamq3lXN5uc7Sy+TCOdS5qECWOJPNIbGsphdPgYr2qyhmYO8d9N9mQnR2ODJh
StI66qBIsZqopQYAY92SYR6JKvWvbV1Wg5+ud//Eh3D1bXRNF3fdvUhvIpSc6i4s4e9abVQagAnK
DyaH6EizvuMMhFc/kqbv0ZfCzAq01pobQZOOsnW1fk3QmJi4Eg1rfx4ubwYAkl45VivxTrA8r2rg
n7iSfvMMSyviTRcpTHp+y8DbDyGRfbuBb/dVq570IjkAbyFfEFmQs1/CHyFLxgCo85UTkpdWa7qq
Nd8YKallA75jeAXWblFMEvS3BXLMm6IBtOH+aRoybC00a5WMELu1knxcPeH5VFk+40JuFy2mvn81
opuXBBaJbzRwUSEsnskS7zHLu004R4MdT4fi5v1+ZSCnwWhMXwVcr7G3DyXiGH2CBdGUgvb3MfJA
wdCSac5elg3pT8f8ib9BslobYE9SCy5C3Y7FhTj6Wns8riSoTL231Mo7sg0I0J1ZIcSBnZ+J0q9C
bezLOMbRYCQif+qjwKclMqDLgWlruB4c+RPAlZvc5nHTHp4Fp9mbDpoSW0I+P1e3MgKA3G3XfDEA
SG4Xlz3hZSvUe3GMFUxtEmQ5Es0cEZs7bMGg9QX4kNkR+gxKSqg7Ap4oGYbc5GMl6PHrGKFqzRIq
OnHpCdgDi1lp/h3uYJaisM5tBjjjdsWGVfCDLQB8kOIxepoZXpV2uw6Ta3oymi42c/JodlntN3mj
SBEY0VHfYT27YTIZkRdpE3aL66VnnQZaJ3kN85sYGNzcF5k+G2WJAJ+j6rvf0GtJSOv8vXnUmqm4
bMAEX4mDKFtkJx1/06IX1WTMVyNbfZYtskANV3FL/RvyZte8LCkoK9fcFnKZ3EtGsOupD/LBQpmY
nAs5KAeZ7bk0N0VbBVCZXqLSUk4BQAyUzdmrUGpWKwLsBQuYQ0eeOe2rvAIcW5K+PgI26jwHuCYz
mb7hv0ifcxTsulg4f7y/MhvZCPZu8lxzAxybZZ92oaosR7UbB+1H7/bdMhPEafIhqQotIqXAcuJO
PL9Kzt87miXv+KgIm1dDa1nDn+BbsDo/0wCctRG7q8fdJi+zksghks9mDhxbc6NBIBZR1+KRhvku
7LjjQjj0hNW/hMdGI6ulBrXxw7NmwaYv5mhYeVcD7P1H2QyrAxLxwnEA0fBCMf8PD/UgbayrwypK
uQ66gbPazWiDglo556JYl19NpHXVgQ/7oFcwMAANKB4jYk04cl8BBwLwVyQl6MNaubXkdKg5oOwG
/Ei5g4DEWANIO065dCwQg7TBlLH3x+mjoiuaoMLp6J75Qw1exrfYx+o6Atl7L85XL32IR5C2Hl8A
hDIWyAGaprx6OEqyfFVeShOrV5FO/9v2wNJcsECi56COB0h3Klb5PNagJ3L1ojb6zxl21qlPVzAT
PCyGuZBZjDB2s1w9Fp3hSUp8+fFNiEjvE6khL7SCHmlbkLXugDsyeTJ0QkSAy8Ykrh0zQHOFj4uq
5Kmzq4k5UWOLgw6mHqm9dMUArGyMrFR9/nBR7T4mTgfWcjcgtk8+WRUIGbkmGrRCBf9XHja1EhYL
4N+Hv2oT0xbffbVfyPRFlRpm0pD8xOdqRKSiUBdFvD/mLG/1pU/MdJ9LHKetc7vf54kRAGZfJSUL
tBxQfs2f7o5x2EfGM7gRtu3i0J4BShQpnJLtvHuvEV3JnQsSJHTImGFLCEwD32SgNAWCEmDPSbIc
H3YHGujp9yepNzYr6dAJg3CeR+8PRIFyzSejia1FHFG1JXYUpjRT+LqzmV4bZvZ3M5rN68MUxoqJ
sb69+4P17UFsaHfDCq8z3bAwUPR09YlvRcxtO+TXWJLFc02OA5L+WVUs4e3H4BM/B1pKr3yzXgJF
FXxh/CcC2X7uqiiRWMlectdVOd4Fj29VujbJ0NxayYdbNGjQbaDruxxVUwmRdVgMWhgi1QhlC2fg
PL1Aexa9VjvJn+v1mzbHRpn8eEN2zxUMZeSPchD8y6vVU0BiF4nFEOMzUt0+bOyyBJiNvbKotacV
hindlfuE8aIP4GTWxhHjTT0+d9IRkFgu5v0qPNejtK77G4qsyy44dsSN2M3zdtaRDEQlZlJCLmO/
l45iRNmQv19ycldAm3NH4oO29KOWh/Kmlmobe2ZfMSYNxq7gskL3FHL7XcxXCcQI86eWYQWixPN5
UDVZ8Uj83Q0ra8HhU2mAq4yu4DoYVcz2RVmfgTKv/r9a7fFd9AyuDU0xpuy1luIBDs9X1zdmhK/0
0gh5z3e777VSxrmtZYAdUSegZHRNfz5OkDVJTYPl6UqkGyUcYDKURg9/GZ3z3PM9YT37jUKFfG89
+LkymCHr8/TVNA5LuSh5yc9diHrxWoQPEwDZV35+dwyAmS4SmlCSR1Cd87g9EWNJQxI2oSa0SnEv
uFDxxRw8Wdl5apWs5E46yPIrAslsnwA88P1bmTq3WR9YvtbspOCT4JRXqWO/XHxA/P5+7SXwgmlo
e+T+ypM/ryCnHbHWtUBjZ9dgauG0+vxEqlC1s94MsukzCK/sL2328uNuS0iK9FX7KuFBqTf+Bm5J
5urLTWodRsdU3IueWnLeBNeT4o5voG3bxpTQXIZvRRxmsUgsEJhFziy6B8LLQgd+QCXBjN8N5JG6
vItalN2iOUPYkh+CoLpT6sSOzJ8yFdu7nfGwRyKU/tQznPZpeBHeG3W0gQ0Zx8P2WNCL2L5Svflo
Ut+9ntNJymV9WaZI4UI+oWPbVCEwkcev2kX9sKyPOB5tu/9DevnwR6cTQNNfpXdXQy7TfzWz9yXc
m97f05vQeA1LLmTeg5XsHzweWnumtGGvc/v82U72eGE8YMScCb3TvOU2AciDYmoFcgIW7kyrIQUA
rnc01BNRzYpN4e1X8kZCqJqdg2SwFKZI6VaMIZItOYaST/TAgv+pXOA1d2Du5b+DcOvfxXGHNVBM
aMWSajKbAAHtWQhJDgp6bfAiZHDmuv9BeT1aKk1GaF0vJZImZiJSGjOKOxvbQzclje45kgq39F/z
HolNPNKl4vi/7igf5vcGNY5YeitcTgkFDaaP2e9T4f9ir2l+OIwQpGkisarH1J5E4P+AgnMGtKas
hufMY64/gST1fy4Ll8cn/W2H/Q1Dn6sp3PVRgdkIim6XlEjy+/dBaALqpLRBbeZr+rEK+Qri0Ucr
q7sqW+sHWBN7CynT99nic7T060JpLK68g3uVu7iEp6el1TvvhapMhTALMfV+fTgomOeawpoR2nb1
Nh7Yz6bLfhVvI7pX9rivGMP8SK26jUF0aY/NX9iEOKsbA5BtHZPlc0qa9l1ryjzac3hcmqt556qG
kPoEECZLBTVZDqwe0GPoYPh8U9xQAzUqD2ZLE1G5Ag6CPQM2pCJ6HuWxH9PmK9FKcS1dm/5EYnXx
h2Tz+Bd0vsRDTyDYKPmmCKg7CL1z/1kMZG9N5LBIfwGZtPc3AoQFo64Zj+3/yo6CvUC3H+/Vwoa9
k/qhPD4LJFpVjaiw9vPx7LlK6AVn4XSGQBwN9d2edEngOQkY+Yt161yvLstbffsN2BOIENJg03Cd
XAFMuRE4/fZZpYTEnEYkVzKNcBytWOwSlxxp/4nsEvcMp8c1FRLHCKFNJtjJNUw70b97vJcRd37P
SoG/j7NpLV4B7sXKGw02BcRBQgSZwcN13GmGjKlwwH9Ao27QR9fTEzaylLzfSi8hBrc3GcgjtJEJ
Sxa0snbeo28AeCmLL5YrYOj9+vLTsgigj3qCFKiq9ZXzzJPLgyozeXs0HmHmD7wey5KIVMHL77CZ
81Oakrhqz6EHOPD1MT+ZeSRFu4SPJA+zLDPskI3qnFzS4QHYJoQX0AtTzAVQf4OTFfZ903qsfgbE
Jm39X6VNoDT/D6qRK/xRGDwgj6orzeyTB0FmCAe/uPFNHctk/EnnMjP3bh7rLwCAlSc6zUDytY88
PKK7tHIlG39L5JcGdTLpa4bVy26/bdgCQVKx9Hg5zQWl+WL0ItneSED9TrwOle/ZI5yZSaYbUqs1
NKOwP+ex2Gb6H0gP98MVrSr1fWRKUhzLZ9ssN0udvxfeVPb8Bkam3/5sQO5zMrZA8/3PdWlAixKu
yQMuCMmjGMxDWKlfiigMvqZR47zVBVjDEC1g4qeANvnWr86VAU+W8zYbicRJ+cxrf/l94gMEFxrr
WFr7Tja6JgG4tjYFMZM3gEU6mIp4+j+yC3AULaP3B8Y6kANy5HL8Y/6AwLtFeotqzgJZusnmCIqt
blxuKZBmBI7Dcrbrl9hu3zaqHDkZl3Dilh3MeRUfQaBaacvCby+q7cMMNcl52o5SklpW515sBPPt
ecXwmHYqi0rm6SP3FZpusDyUKpxt9zNkHJDWEvdO0paEuYj22hzQM5Ap87C+7WB8i+Thn8kIxkAz
/CyjwYHge2wIVKxXrIBG3hv2oM/HJen5OIaAntsjnEGC3KCb3NIcVjEQdg9ZdiTlihXAUj6UWS2W
0lqWhesxgEKEYqKbYAg1DtQGfgJ9gtEtcspfKWxDoFQeabMS3FUf1oMvxYbrPPBmMQr5kyGg4gIp
jebwiGuWSxf8I3ddRMBeSMUzZs6HaW/4jTiANxgphSpTvT3Zu6i0vi9C5wsnCJ50Z7ADeIzXNzM/
iNwFHBvYo/5KFAARIZzfxCszEfjZQEvR3qlli8AzduOtmBrZp486s0nctisDxeg5KOwAWDWoys1r
YmjqR6ln7I2SBGnI83bpu/Fv6gC7+gBCRBhUPgH8fx1Yl1Zg3QhiWUyjKUaMeGOiRD7RcYXXSypD
lZvfurJZOHo5/pM4G3LyMxpwFa3v2sAZiVLKJHlk5RkeSkcVFpRo3/L+ECV82UBnv7in7D6Dt1XP
Z0izyN9IcgKXlUPWvNo4pbjhgCGvaBW96CmSCOjxkzHwWYhBi7+ooaVG1P4BjT2cYYfDXC2BdFZa
VFl6JJ54jpAvF/JVnq+R6UJrPrajLBqOImIt9nap4IjtgddkgisMgJR3ZaZaBcERz73rjkMGjdWD
wIRX3+pxCghZDxT3hE9xJQ+xTnWmAEjpeAqdVedeFc8vTWR8mYwfRa1ZGJen02yuDtkbflBBy+mY
9W41+5rOPrI/3qBHlJAz5nzhFX5V09STVMja8t9Y51nXElnX/kb8vv4EKMAIdQMUjTarHXpEbEzP
smsM9alKXuOUU1AHznGiB5ffEYqn2Hrc0gTwKhmWkgjbNLsBJJ5+DtIaq6PGpfNaL/EFKEiB/7tI
+aSvKfhsy8UcX9puQYPYupudxBcWtuiLoJoxTNBQx1yu6BzZxDKZ0odCuixGv7NDiXrYGg+NTgT5
JFvKJU27LeGU9SSaQvvHnL+dXg0yylLkn2ZVTL++KN3heRbb3muL/96az5xP0Z+HkP2qaPD3T6M9
YalIR8jziIKkkl5Fk7o9l/uJsxtQwWZW+Sd+TSCPWsm2TXYPr+0uTjN/rxYdV/AGYqk1nwg6xrF0
DyeY09aeIefVhgnMJ3qdeM7UiZxDEK8MvGmAA/uuey/Kyj2iF/2wqWFTMkDU8mvU94MMRO+SCdS8
+WBJgVhKe+n/Ba5m81EK1711v+r1PyTPwS+zw8mLMZkJDoYSuQy12sRE9/XJaTkWAfpHQgRhtMcp
hnfH32AIArP3zWCVsE44Qin7/fh6uHItHeshweo4Jvj5PJR+WCZ3EZEmlA4ueFP7i6RjNgBHK4/V
H+fxtEAF/7SKrM4Op5VznLGM91epFi1RiK90U+zn+2ovFAgAmVjml98STZBEo+vR6G2U+67Dqhh6
vtqee8uS0EdKqagRxLYhG+Rl6YWmmnlYVK/gYKAVADMwQ6OdG7iGH3vZNpWHN0Aql5psIVwi+Hzi
gZekC3Bj8ej3pno4v4Kku2EbYB1HrJ4ucX21U3om1+0ArxVA/fhAHMwZwO319Ct3Xdj/2WYs8De1
vLiLJXpRDAAwC1fSqY++CehjhoDpuNvlThKKmyX+AdUW9r+EZw6lJxO1wOxRdaXX2sr1RE33REu0
raNo9nxhj410WyOfpQiyKqSz5EWK6sLwpAJq0pDIGxiTfrCY4i1tz4rHprFaZMP+cFfGNgarmCXe
lnsqNT2eDpUqE5S9juJWKhlHYbj8crOcefW9hTY4s3i+w6xhTwlPWiH/Av0NTqMO1Kchbfh1dHIy
4uIEO5QVzuL0PEQJXZzQUEdEHwKEhaz3uuG02k1/PBnjeGChbPhfKoLc8eBYnV3BYCBWB+AxswV8
iyh8f7l94/+fcoj577eZ1QUIw+UazB/bXaX/KFpw0eKo1oNKUXdJWH+byMVBWRXq6CIKUG1yO7Ns
6MrlOelybq4buKugp7UIWq5haGBjEc6BEeSdh2jEBdjsXDCKWmT6de5fktmQB4YxYboRlB6CV4wC
Lt/DccuLhE8nWyjj1EfnQwgXuYpteFcBRm0fNoM8StfJZL1mZlI/86T3aN35qpuxthgQA9uLyr8A
uTqndLUH0x7R+AOoK3Fc+PO/KcIzX5vEVfzixgtMS87x2KUrpwXXXmjeCxez3PavoNzX5vWKpvoG
4lQSiZbrl0N5h6i+H0MfLZWTV8Q1DJ1Tjyj0CynbOQCFPOrE3JDHCKa1lo5bgSme/zO0H7Zr7dUr
EOpyeoHa0o0LkDqOjHZKY7Cj6nZtK2BnZ7liG/m+VpiVpzY3v/ss5boBmFKUE1F3VDHGdO4ChbfL
KLlsVvPZVCBHgT8bBnSgQV67Hn2j2tuYctYe/QxFbWHkk3aWRKlALhis4gdPnyLi4k2AtAbhdj5P
a6AS+s+DvrrCVaexQMXOY59JfdXzYh08f9lZmDW35z9u+1zbNOD3nQYsVkCxpyl00Iwsxa64stBt
EJqB95Ax65CujpdNfXVI9cKCPMsqX6Yl60wVUPExGBKawN8Xwp30JjmRxAUI39Tn1y/aiNP+6sFW
pMJYG6GfoRx4PY8Iz3zh4QD0r65pXYJAKPz8McySitSwWjF1Ym8FeY3xJNBUum0UN5Qd7rrnid4I
bnWkLWbH4nn9z8N50YML4ZqcKYmKYYFVpcAue+IoVlL2tQKTWPvy4N57tO28RajNoJYsuKRqdETB
2dduP/cW929NzlR0ApXI5Suizn3zBHzQV9ge80w2UyZe3t1U4ycB0wY/8YixhRKPZI4oj1YvxnQy
Duq/k/Gnrs2MsHsI+SllpXpzVDjPHzdhSVasa3M7kuISZCbuwYcUTFEVq1k9s6X1/+E78OJI8D4W
FDiziBgcgkg4u6FfVVccdq2By5cBAW/BT3wFYw0npxiHj7svqyWOjjiNCUbOo26/GlXkg4E7f4Fb
i6jg09KvrAW41R3RTro7n0OGIP8w0KZUYwCv/JTi2NtfhnOHDFyA6Xwx/L6MoObCJLcums2aG6Rp
u6pPoNXqIoACpuuk6uvLsngcX1cclvcLfcTcit47IafZtZZDgoyxcnwtUPoXfifytBj12mpMEAwV
v1cXIzjjTXJdSuugug+vAtvPxcasJmFrnDUTh+8ukF0h0ixMsaY4yCqZHfc6wAcc+h9vZxMUV41A
T3YDiLBR3SLe2l0eVFn5KekSFx7bqzfoSnDrcqVB3B3+eU/1Iq9WlME9JIgdXWZ1PiVfInW0+azp
w01Lj0jpDjZaK9RqHALWuHIr5X889/z9HhEBLV54f2lADWTIRi8GhkAKT6CgfrXz9W5bg8xe0JFp
8V8+VaTEFHbQbOooFvK94eNE6dWxjgFHZf2aEOkFgitg1jV3g2ucg90kVjJXBDgiAHINlGn2gZht
YHkYHA2FS9EMofWPgOHBhv34hN5o4QEUw4cnFZFOX6dl/yki+1T6OG0+d3u7lRjI4jOjaq8bk9zA
v4IxOtbFB5y9qTa9fC8RXO+0fEz9Kdl4YYXKGbxZHN+DqxYxkK1AW6E+J7MLQNtNoKO0rpjzntXI
bDKF6c3iaOPdyshtk+rlrdDLdWRYzM76NBkxXrD3jaD99BC3TeB4eV3uovYJOSE/eWfX7jxpX5X/
U9GMWB/uH9/QOdhQ92uXPc1MOBaM/UYOW7/d3UBQDSlkcRwb3QpnLXVS0LExWERlS2MVgSlTHDqT
qAOdTtil6ZMdqBkTFnB6UkU9S7a4nn21gKvd21T2kyRzynuNp7R1t9aySWDxeJS9Qwo3iqcLTjBW
zpMZApeQrx9X/isReb3r/QRb1kBrtTH6sd+sQRbHa40UoYXRG3KTtynFFGjmELUtwwcyf7++qNeS
3wchnNqQrovmyynN0MwSkiXh11pTjf7pKbirMKvItNmHll+a5n+PCNkWMcoVBfvDCVXboID7kQhk
HWJMFSVzB2hsM68eSuDs6O79QFFE9Q3WA39ks+Ize6Cl55NmIB6QQfzY7RG53qcF8sXL9UuSCeSO
PEiTyUiRv5G5YwESft0LqA9XmEpAAFQ0/SKkA45YaKoVOi8YDJ7HlMo2UZeYENIXxfYQybSTv7TU
GU4zNUO24BrWI6J/LeoMXGtn9AX/pWDXeCkDYDRlaadtbqiAqj1Bn8wZ+/wSHA/p8/gFKCEP/Qp9
vE7YoFr6/EqP3urpTBtw76NzENHi566BcwZIPVsIDueBCxgBk3ajrNOYHbJn7ItTtFrCQBIsnQly
z2nS8nUEe9qFJUE37PIWVRlR9WMwqcwTFzAurwAvasp2AwEmRDPR8NHV31RrKTB7vd+kINEWv5hu
4mNYILipO/pkKEQRcNvC8Hcf4uzgayGbFV2RIcbmNT9aog5JSnmut7k3jfdrYhbPyHqoIbi52SYw
8z/8qrenWCq1+85VmUGbGoS7ZZtRyIWc8/IyaPcUHEuBTLwcRuU7JNVkEUxCK899xyOKUbH/lg9p
6Y6aKV0wHGTW5kOv8yXU9ieOBgv6O8+wlrSzR/Q2Wg7TARVA7yec/t7+VS5Ssu8DMGKDOhoUcTs2
85EtT2glJ99KmqOLYEMqOtelNUJMoQ1ubKBca7DZwSZ5f0eZ0QNwxZsCJsYiGv/AJ1E0zjluCdGJ
Ec6r5OEQlRGs263Hwy/MV0mDuqvrWOrXYiHUbIOHR8HEGDRcxRjxgcIiBFMl+aGiKyFnAuQzpcit
YIW9UI42M9R9vxknkqhc2X1eURLPMZfnmtS5/P/R8MvHv2j+KZO5Wis03YCq1hoKJ4RBeWQ532th
yqBfTf1BoGAYN373LRcyyplqvWDdS/TQaB6cBnPxtbJDUH1HqeFfzzof7ykzbtHEKdqk1qwNhcVw
E7qxT+10Cu6prYxyaYRkM6AJONWLU4dOtRVhVpHZLr02Vpj9ibzYhoXEJKaaInE5hSdF8zGIe8ID
THNhtmmKv27ZYLLLCl3mOWSde+O8k8Ct20OQ8YCI7Ymco2bC3PCLp4ER2E2DfTsvGSh4hVvHDfKR
VHq5aeMTrSGlvNSX4CWKQNU3ZYWAlr0rg8suI1ei4k6IDl++BdWgkmAfYVrwKYOLTqPZCm9Dpu3Y
PycSeKHgh4Lxdk9j0x9neP4tiDpgk4V+dTdfaweEDpuROg22afvWq1d+MCx/z4Bw6G/aoQ7S4YM+
08HWQMbUDVTASYhtOdIb9MI7XuPPM8szBnfhDMbwHgmSgZ8+b9i0yCUmt1SWwpGqQ/3cW6CFvquv
PY/nOPlkf/nV3qBRkih8Q5Z9lWBAY63AGMXS0xesyPEv06HBVbXYg2g+cZqL4rnQUwr0/ugAbfi9
y0WVk1ocGSWkSbVuHOYy00iPUyBJfCwWYa0RAVrNymEomVE6YeUbiMXHTyIPq/wAVibKm1kJJr8k
RIoMTZ/GARWVZf/ll5zSyeeHR0KNyrpZMdq34SXuAySbSAfnfs3n7eq9gSIB99/jSw8PAODp3cAe
1ArAQv3oh94oixuVcHwE5joEAg0+y8ExTadSZfMfH4PiP1Cnu72xrc5+IlYvShJrOK5i0J3eWnEH
cB4XEE0pxIXqbOmZkHzpivGpB/VeEi+rVIJndcLMLsKyq/xf75P3JvRlgUY5xm8wbdMZMcecgC/9
PQLvkqpmwOGcPhTaT1t7lgf9y0HdZM0W/GqY3YUYbVBSHOEDVocnabqEb/YLBafTpebSdu6J6qQ+
M4iTyyrSTptllJFZADZkY0/vnV1FFEdKx7HlaIwA9T/8ke56bDFgP1XttvcqhnrJizSY/lxaqB+3
GcekXhR88aGoBqjXGuZuO2H1f+38UpseWN/7vAUseO/cKlB83v1WVBb0xTa8Gqyu3H0SNZPR0wtZ
0EkSrrKd1C6sCDhuYbZC2cCRuoIocSPXEGReh2BrziQiCBSl5Z1wot36WxHjRLtd1F7gzy9lbQH1
Jeg9PS2Bjw/fguUOPsA+se3Zej/pTipW3nNQZeb0ongn4kA+fZRMk5cytIRTOns7qvuECEwnkNod
KZd09yvhcSqjnTzaTpSHRlhcXxcFGPJYF7tVG0j56eVkU36EsiktjCkRb+wqjal50ocswvHEJhRy
hj7noDm9zltyx4kfUpisEU7kn/FmwUIIrKRsDgeZXIPVMZXl5yufAaWW5IdRf8UTACP/h6NKnDCB
Go18jKSAwGbjWEinZfv0WIKx7JijEGqqzyPVPOrwhY9mjHwIiNxm/uuk6hFYUvSxYZo3W7UFyaS4
SN0s4simFXR+lgEdUt4B636TSPF+CdZrL74WCTk22Fl7WRcRg5nO7P+bL/htAYT2AfxwB7oXvS5Z
KAyysfCMBBnk0A6biKLo5ndy2pYqpTk9Ab5RBDvdEt4PVpP1XQPLatXr1cXmY5S7/cHaVB3eNkmy
XdAzBzYO0GZ/lDtKtdboG/5BN1PwQooBjIMRY53c4TbtXad0Aeya/2/ffGF1JNPllwtHREgMoyez
CpMBIew6bTi5dTDuOBYZ6cFyIcaRz238w3fWdhh3IJI0rXIM9cZQ5xt36RBcM+qPXRl6OsV/IobJ
o8MHPVEManIPGZmKZniyZ3/72I7jQQaMFeapSeItdOquocx3dvgijXrTSQh4yl0tN1ZrlQpUC+S8
J8UVegjSb5iNhGZ3ehEa/Mexwp4Q/Op/DWiVXa9xt5ueo2B1E0CMb0k535p7y/1zIJMMVlHkRSt+
RsQU2WhPlBwDh3gwPQBik6fQy1NDyFpEkXnfTNrwongztXL3t7opGAFvL1IBkTh8i8eoRJzhnC5I
fgCD/iBXhr9kHAT3eush9/DSq5paETgWKWJBDamnf4oXLUyK3c+P85/AF+Fz0dN2uGWKQYmBJpMv
UipBjfKdHAGhXuCZQh7TEcukTlxPJdZdzxmnwr8bm9T/526G+tPHSZzBPo4caMFOv1iipIv53bnO
rro87IDh1xTo9wCSNOciU58GA/eGIJNbj+BMoJ+CQj0+ej7a933n0miyUvaHwGnqd4QAz7YioXYb
HyEZ0SXH4fUG7fvCFRAhDIYb34T3vg4qa7dNmieZMUakT6gE/TKRpJ91aI0bmC+MxJyEw3bYqKeY
8uucs20p/RkYH4aNGOai1nbHYOFviVttfxWe2oTOxAC+RI08syVTeSk5jUxTM9UXnVZI6IzNG9Sk
YCC5LTGmk0441aDzoNeTua6hnp+caEwYUFvJNyrTu065qVv3F8bNJLwHspGiF9s4MVor71JuTxPG
ynBzil3h0vZ80kPausa1xy+HmiG3xVmruWwqWNX4AmTPda95l8wMcLhT80OCSmFxGD17USDrpoV0
Ohi8mKhHShNB5138yM6x/qqoPx/AiRke2lbhJ2uK2BhgeHABrhYD4pCJXMBcZ7bOY2a3+AgYqSiw
LI0y6bWrqzg+bMvn0ixah0tNfuGcsC97v/+5ZL3IoXW+pnZPOFGR2oqHFtnucD1sVPAtdekD0udS
1fHzcVYF1f70oKghi69VSu+3cWpdA+TxT/aiwre3MBrTnme+acWE07V8TkqO9XWR+Z6/XtubUpUj
dT3zROGRyvAEXQQciCU7y1M2/bSBfafWTaWjjPbOLCwrZc1y70U3Q+aMuFT9r8XhWCPbGYzzvfSN
8ezzZGG3N6408YupfvMlCVwbxa+DrAtaENzfQ83tEFJwoC50HZGz5Ckk8P8e8vY+OOS/ekJKBZd1
5Bu15WdQGHoS2/Tfx/nLS859j0g74QM/ByTT5giFBG1lF+a3BdEixj+rVPW87qXCBco6iDeWgwoN
oBymXw3UDZPUC+E2sl58RBKeReBMi5Y/nUgbgj3YvzdT7jwTJUYOUFsIH3rux35qDwy6Rso6NAT6
XVoGNkbfpsFD8v46lg3wb/z62cDAk1o4xFLnpEyHcgCRsbcLs2v+prX/m45zWQzBh8is1/+HB7Sb
jMjncTS/TaYA4kkt2a/ZlKx3VMei6N71vWWdafgsqBmoxj5aNvRO2sVTXxmaxyyj2lcG4O/y49iQ
wYusv++G4TbflfJi/xxMW/5m9V8DAcojhYv4ervvMVQvcRBM7TnrPl1dy2jPqaER4tXcHykSxhSV
asN2pD3ciKbmbid74ZPwiI9yTjQ4cDDLvSS0oyLx414CJbhHlTOeUfBt1S1X2VJADMCJtpw3B4eM
U5dPtatVcAZASNIAQBJLKevhCPYt601FcxApO8wNTdFieqqM69qWjTpWglLESc+2jtRDdNaZtAnj
V5qjdo7Ow6CwxAvLRzK+v9bSFKoKniTwG2cMYdgxTT9wn2ztOGyM9+k5z8fuhtUxutQI/TbXNJKD
rOnZ+zzLpLU6XOtO7UtML1YYmNR1E4Xp/67z9g9WkAfKKbKbPxCJK0p5eXmqRRgKGwVmVu+crdaT
Kv52rl7hhbx+hC860ayoOveRkZBVkJkcb3aNIvQ8L3aMGec+7XLyxqK1JS2lIUcqoZ7lxTy559zm
EzxyoV4FiSty22nrKq6xsmlleP3ZiQ2gQm/SwborRXWJI/wkR2CtTsGybi4c0IQ0W3sTjtXu0kx/
dE3RJBS1FLDVBzNPlXqr4GVpeAmqJfgGvnsqD2ll/FuFrqhiL5O5bMgtspclgsaM981C6wWaSz3y
14fFuhvAPCEyvcathGHG01UYqqaX4e4FlAfbtbILm3NKsyJ1Ha131TxzxiT3zlNKIL7lO094XfHn
4x/LxewPhQGxvjewVBcObIVgU076naXEHOlPTNoEvaL3nw3/zJ8WuchscNPZaCoaAWAbEQzVCQPU
uxx61KDOD95dFDx+WAl7q8gyFDkRc2OY3sG+A5zMbmwHbXT9GyTqy1VWJsEItP0L0eBd6ysDp+pM
XqwR9D3NdOL7O4G2rhdtPqZy0WxmLeRYeEA+81ocFrvHrzLdvHOf95h2svS1ne/+IPvCG81N2Ls+
2viqA15K0My48waPRWq29rJYv49lj8pRco2ke4Fm9+ENRgILPSnkn1u5ry37Eb7VyA4RNzQnq48a
Ap2AxRJk9ldv7tprAl9OpWua0kOQYbG4SZvt+/VIfFldOSbjXFluPseSw/8D80x/V3JqTqne7IDo
49edU84Gsme84ag/F5K+adzN+chHPE7FTSeSvyucNPnz0wI4U3Y2M5Cg4R17fea66SdV7ppcmGQF
YBYRXU6sWrbE5ZfVEzli6+HsakuEm2b+blZZ1yaU/EiVj0tZEEMkMST8lRzHnOQHiEd5+qwIfzUA
5mTeM/Lu5STHWWMdR/K/msa02iSRAS7LYGapW7XeigG5f83aFc5u33AX1CP45JrQeDdNjp1vetuB
BMQjFfrz6EkWy5F1UB17HSBUc2cjmN03SgRpxewIilyYySkykWhQiNS46MGlzIz+MG+nNp++9/ch
0dZtm9ysSo6pMZTw4hKm+QixzwVqhQ7V47LHua2Nl+yL86zEJ46Jy1lyTa6VgT2VbPRJJQsBD9V4
QxUGQLv1gAv2XdYP4j7dStKUnL46AM5QeQTKLm++WiqM348XamSKKlPNqi2uXAtWTy7LieVHF0QW
eLF9gpTiGwR1tZxXMLjq6Pe/k8/jDZboK9WFi/oev+/bO+maXKTZn7T4JEJskdgQr0SPe5NDDiYr
3Q+mQYIflxWdbwIULEMHhW+NNNYQRv5sdqfCM1Yjq/jGN9izANJ9VhAl+o8Ls/5Ll8+PLty45pOR
d3Z4Cv8Np/1Rt5lhdZquOgh9Z5KGvQss00o8QXiubQHQCEKb0QCm8ygxVlPS4CVFZPaDaLTUtZFX
PnRyPZKitJSOLTLyK6JQhPm/EDRLVp+4iBpuInCJo3OTc5mS5sGZXvGOHvbqzNLALFTlQjiKka9i
QdTC74uG3C7hQcd8TAB7u2izTbhmBergTAmqCM3WFOFg5eyWhpek3o+HT9n/VBherv92rTzEih8r
B74v3tJCj4W9/hQLi5ZPDIc78M2l242WHPS6FkWHuvIFAOlR4WI1siWDgcrOlwk10ooRWDIxpVhF
Dl6ZIXwYBf9dZCnq2RUCOGgbHegy9Eq1/8RYReH3X1ApM0aa37vV6D3z19H7JtgsgaXqy3QZkyDE
+WEzT09B4+dvL2gwSRxlY8Panx5waaZ2JlRBILuJWLpa/vp2zM71R7H4UE67dBD4Lyys+khA2ByM
dr40O3CoTF88kdMfI32gQME2uYSKeb5OlbTOAvzheXsTcFF9tpEGgggOflABCD7+SxbzR7Y8J+/w
S+5+2BRft0ah4yLPBNBuqvGIlHjNuViqENuaQlotWqldK+aYyFJJQzdULZQRwQUtp1+tTqgNlGhr
vVXnPKQ1/df2b8fd8Y6hfTmY2bK/hOQsfhymWITvVcY+x7nm3GMxviTIs/+OM9d2LyvY/ByWKAKI
LfC0ZQTL1HONyIYW//5P5aqN7jKAuV+mSYnONMbh6kmGOHYDeLXlfWK3tFY/UXZMsjBzFc8CcYr8
li0XfAqeMQkaTcDhPSG0DCixJTzR6sTQ8LjIxH6my256zkScVjHKDHxv04w2S4MWGwSdfnCPbum2
4QxBV5yvQMFNt2612jInNMvFnyIPwSpcwf4WRRYmwSWeSjPEYLGv0yBsu7wKYYAd4x36L3Kng6E3
Jx1DlolltU/KFxBi8Oty5z+ee/y+YyP86NP+vaBcqcgEN7xJZT7Tdsw4QCX+DuIvO6aXrL9Wq7sF
+whrat8Fnwy3YARC937vFI8wSVEGn1o1zj1QjkhBmrZLOdbkkK4MIYkmn9TwuJpwoR2BRVqA3T5w
SCSBHM+BiRLc2UfM2/K2UE0A68ziWCQYmqANTI6LC6spYV2v+wvxOi5yZCzjM3ZkKB4O8t4ZcHIl
WIESVDtfKZh98OoFvsvHtGxja3DnhF+oN7y8ppiX6Pyf5Tczxjd18fMxgUau6Ap1Hjs/Y4Rhbcqd
izxzx4ubUUWJNsGu/IEn1iuQ7o2v3W2dF+I8JBHEldltG1Hu4oIjzoN/BFqzPiIDY7U2NXGqgez5
8VfnO2YFWTwKOtfYmt/r8zE7rm+ZLoomVid8a7diRooiu07bCURzH+U3aImx9W3D2BmD97xmTHOK
3KUro8ecNhmBu+cfhO74kn5rlA16lWtq+uxlrb14HF9lx5axIqdVJ1S4USKtk4sjDnmAEFsWr0l9
XY/X7yZLXBxLOUmwrIcDS3U3sKzq0e40QEp4yQ/7crnuDnc7QIDTsnECOXowuZ/JZaR36aGspgXY
iWrQb/2HjED4efAqvkMfqJ+jFCFzHldMzaFuAzghV7A8PqaAZBGeEVAYIPu+nlmbFVS3T5JMYazs
bUQXtjptj9tBpSUD3i8FWaJY8YJGeMSkWSFulABSt5QN2RHBdSwNdMIbasaB6EcZHDd3+sFqbpXM
Y8SvNnPWEM29FxiC3rBauaWOtGYtWiCy/JDv94OOoxBdMMyoNYgTO96liMKPw+Ad0KDiZECo1lYQ
dT3EfhAXvrbixN4i26jI05t5EtfXipdBUo2nhywhgED2K+39iIfAb5CukvZzFqDPk7ujtoW02zej
vbKhK6zCtWJmy2fFH+VrGFpiqKIiboyBsZd7F1UzGVQ31drzVw5/BMTqDeIPf16u3aiJL/LwyVw7
Ruz1XYdFuPwRbhOWc/ZmxSGrghJT66XZYJPBniAyCtPAV9W/KbJltwx13p6tQs2kpBF/LcEcQL9t
/lBhdvERSLlSYWPSK2Msz2qyKoVYn+iZY0VWC1Brd9otSQG66P9SoLWdjCFRzesECSgeizWdpNL9
qAqYFvfcm5juM1QEUpBjH7QRFjaCYTfWpB4PkT1zGKrKJkJ23SvL2SVY+ner+Xz8MphJcXb++4uY
ddWPHYLtnE7toPIvDkGQ46spGNy8celhxssFNnUNg/EN/pQC5wfKtPfJCH+FW5pby8w1xOTbWM8f
eB9+WnkFx2jkQJX8ekVFzXAPwkWQQyw4vTmkPyzVnZ8N3upL76+DRg5NK7txbSPmNjlLjRXGmtya
cLm9ysBKRFB1veqfpvvB7lbMnNv17lM8jJTbk5R+mWDNDsytOJBAQcvxZY+9meyctW//6MipHlsK
jKpgmDKJsfk8T2GAQOUim2gmdJg4v2xx4iuKvFy5MPPRXdWH8vNmi7B9Tq6HNpfrnIIa5YIunfnl
zr0xfFKEbXyJt1BB7KZBSqr51LAWB3r/NBKDWepDbBLty7SUG73rIDajgrvl8yzkjp+mI77fjtpk
mnCy8GLfrxEjjxVhC068DyCUI3JsD4KGW+u8pjgETMKyQ3ojXiZm46cPBnLH5X7KmqswHJxIST5J
qIV4vavHDNmbx0kf1hkI6GMLjN31ccIzgo1ZKJfgoPvkteICR6gC9valXliOMVPcJbNSEsUGGF10
phZDrzkuaoYWbEapf8njsKFniSPEGXEK/m5zHwy1IapAz72fRm0IRIOq3RLV3n5mk0FJamL117yg
dYIHSrt0hc79HNnUUx2ueb+/tuzcLxP0nfSuRbYpzCslGqomAR3oe4+2eOsEnuIkZRwctf1tnAci
HCqPe6nIFLJLUfhdsMUm/jcYzJkAYlGmth1puGcxyZDxr1JerkhDfm+RO3Qstixfwq6wDmaeE7xT
cwwBgGYMCNLPwRQOm/Ndei1PgJvmlofeFC2v8Ap6ohQxpigTRy0iNcIR1RBB5g96L819PT8XEtHy
a3SdfUeshQ4yacwW255Io2AN6sB8121X3RTbbW0u1qBT33rLxk+Z2rmyfyEw0FbtZgtUG9eQQgwC
qs0UP3ACtuKCm5yGbt8EyvSAbV4Y0NIOTQNZMeLGuwpnnEF1+mXeMeSeoMa0T4yJ/WwNZclnofbi
1x7FeH5kK5omtI0u3oe+lvbh3WSTJSR+maovkn4GXZZDPzsA+nrARB5U3E+jXaJFXhZdgKv87tYG
Ov7bJONbFLy0S2LCuRIfs8lwvio/KqXXb8CH9VutwDC9pyv9B2pY/dwWyABjdg9Pu2jeiYWJQF6x
ZYi9ZnuzGYa77xRVNk9BpfpBwrWYXX+fW/cdjiyJ9fPLwLMkBUHF88Y3UAgjOLpHRZj1Bdxl2kUH
rh+xp5BnNYPod0IaXnsWyxs35v9aWoXJ1vuCmdGpzlLuw4zuTInpMwMeLdg69Ne4g38Rr+pxoNsR
BRAds0SxY3rUww+aCQ7wPlDx0Gh/m/CtMoip7y6yORtJgmlZHZwSGkIkbQAdBDA3qzYmwtr0e0/f
+7XJ3R6I7nzNYXi3Poiu8gsA0GtR+vl2cYfGQHXrvkZhG1SQMJMX2O1C+zGdBezRIJfU8n0z0+dI
Gol6rPSJI0NpKhw3LMDBTa3csaZKO9KldfM2ecCOR2iY2sX0APvZGVpVjUoAByosNCFFiJoMLrgR
Zv+PKXlL2yTpV/w2jreIQ+AOIB0/by/lZE+IHB/Ekowo4xdVogECL5FIPf9IOvsY/QQtoZ/ebZNg
UKhzBeBZILXsg0FP9vHv1XojU2tYOZXlgFCLbxdur2jzABJdbq9/Z8HF1VJgs2RawBWuUKZtZO50
5IJpPvDOF4zqWxaP/RWZgrR04jtiTrnPuAd13ETgIU5mTe1DL8grA8AQjbU4AEX4TLEWaEBdh91i
Ltg0UTF1oocFv9pXyiAvYxG57zU578nmmxU5ememaKtqNiRLKR3lUL+tfllYfe/KzbWp71JVu1uX
yVLi9+sknqFxnz4gQsh9GR3P2JH0XWBUqIaCQyss//RmgGWOHElx7CywU/ptj5fGL+zhEOo/WB6S
s5XXQxDs69FvATuRP8ie3rMESnK1azxjYp2GiUTGhqJSrqw3PfIeJWepnZAnztTuM9GtbtRNuzaK
b6C6aZaIRNJtDJxKOPztVaOsbOuClBetjJP14A23Z9ul/vJDN+Ds0VSDOVWBCblQ2H9QOKSIQX+v
a3Ue5F3T9kwLiCGjfIiE2c+lNFndSOvBPAd6/LtqPsrl0WzttU/S1UDPGhlYS51XGuTTIX/sDQs8
ZerU7Lvp2Ib31gNpaXdDzeqFS53O30Z/lIwj0OLuB4kiLpTrdyNcVAmrM8BrVzYtAZh7uU+0mgCq
KNpkiSYomoJo4FodOhzZQXACBrAx4nDg/21vhAm8BZ8o+nFZQGbS18l6zvDIlBBkZaa+/TYdwX0R
eBsCElIeReyg6PQUk34L2AChQHJX8sVVZlkzHL198Orlk+tBXOkS5GajcIqpvcAKzrgWmAC0WWZo
tOJOiPIYNDAXFjvw+p3hyKosKtGLqudP6xu9XF2yurh4bu27lmJU76QVdpELQ5Na/OJKJzNd3EGZ
9bve2oAOZLPKjc6tXbJBs8XCrm3vBD2pATdhRxyWtht10j3Xsi5R4Ej3in6GI2wvhrlIyo6VZQyj
dpYyo5Igc3rPTGdEkTRfFAE9k8LLyqxHs0Nhj98+HbtuGq6L3vL/n2AyQCBFk6HIoij4T1aEWhRU
IBq55kk3pP4OtRNDwvRDKFNePANb38j5S/9BpiStzSMfduZXbnrg5uepZ0HytLsl2t4voa0x+pMQ
Zg9/+I08MWMfckwvkTPJ5IQgHRRhVkt0hBjHx3YO8etiWKyEsY9nTzbIGUOSPBTmGuoOEqW0SsnH
Vs5UvZVRzHhxi0p5LVBzNeUj5FLIF8K7xLjobqVf/OLkTg5oeJUeICsuhiEVi7k5gJrz5p/qIQEv
x3GrUEzBmUEy+7DstRJdhYeQHiw1K5uzzuThnGszO/BOc+e2oM0goVBYqWwv3WOG0wPAX+b7Hr4+
xcgSMARKRXFhTIYmw9SwTBuqgR6znfPQHsNE+kwjErMDp11unXS8BnAjEdOR4jLmWzO9PhePgZWY
4oGSu0GeZBvGpxlx0jexamMPtinTT5c2s2NjUCDYBnggqrPpYm+DhmVe4qQZVww7DAPBthiURDPu
D9+mzVlqKCftphSrw4I6KF4ivfofVRbzFOdv+uXWjUtIwnH5y7qLcXqb11sk/LWs42+LgwXbKBTn
kDRR6om0j3K7iqWjpl89ngex5xELcCxu+Tn6pLx28s01kdeO+zUJ6qCXFQ21zIPbGJ/kE3g1e8Dy
1gSDWU2RHNX/A+E5l8FxX7avtxKgvon2lOsyTZk1UXfV8WgA5SYeeuAHGNamPAZRcepfxieXPgyf
gdE3UWJUtlHcoTEviGMSh64oRJl5lk4ZKslfOffj8hPd55tbEfS9tFb/1N5oOz7/xiWgNIvpeY1O
3DaMbdWAgmy5RNq16lpV33g+8SZpjcHB6cN92ENtLvXj4mf1leYTDCovAhhZHWBUgfxsDCJ6UrEF
TVhROcpIMrN0H+rdrDekvsxNuAohzNkyHPsQGoqHlZrj5lmSwsFNBqW5VoDX38naAZTvkk/kOjml
jjvL3tURHb/2FKffdRu/WPvy86B2SOqjEEXNsJWJaIY3KibXUKSAjW5OloXGBumMHoz2Hak2Dn/f
0pfsTJAiTPFF++Nqs7fwjE1cbVS8jHBHV5RXyWFTxRbg4pU5paClxluk8qHJHzY0+OGct4Ztg8Io
HCg3JCmSJCZMDCqJ8JDSDBT++k7rdJGKsURQKJlCJSPKB1OnylZuPszsB4qamQxgqFlnwjgq4z8a
4dyUoxS4V7lVqZhIVUiouT2gezvoV45ZLb7fEGVyNAw3yUOCSnW9qI7fKOPjSrGU8DwDLwb9jRuz
Qe9xwaGyINP0HLVgrKqXw0tU4XAiNYl87/pJA0//2qrD4dzuV7+owQaf/D3+4xztLKmc4fu7ehnf
3qZW+lw/g5PhVc75AGyPskLoF30HIW9zu91vBcCtrv10d2A6UC4UxvXL4rADA2G4MLHJOmYalgYk
amwzNfnZqwu7HEPKRWavNDBXfExYvcgB2RT+lkJ3YeSB772NZi/zr5y8Z/IPRM8VZosAczDveY7y
telj0RqQ3N3OMyQE7UI+frwrX/PrpLCq9B16EPYmlVQp+KxO6K9TbV/eup4r9h37jQpEnYS4b6SJ
HxDFVEqi25Y5Oo9tGIFMfXYGhMnamI3c0VOcLX3lrfEpjCtKUfs9ciHps1swSl6LykAjfgFPWWO9
119v6QIgGrHQZaygJtV3JI9BaOJNrOkIl2Xn+sPbCH4Cwr7opkPuRPQd6nb3+l6aJhVWiS23QLx/
bUnWaCV+S+oDAqS6K6l3NphnrIRnwFWIIBymcQ016rstm9P5UnY7u0a1NLpeWfEW1V5imaaezVpw
xmJ7INpmvI3G6p5WfZ5UnS3P5Ao/VDAz+QJuHgb/F69WYrNHwNQQ4ZwS0jIJos7tN4q1zderxZZY
feVl00TQcWNmmIjzv5YSGADnNiwrkqQB6ExDBnjaTPTaZyo3HGd3wI2/Jf+p3kCuqzRVYwl2juIu
hX822AUzOvk7HLlvuiazlcpUIH3kGrvETgrBPvXFWw0SJMwRFxtOQOxGfUZ3mU6V1lTMh50dGXlR
8rB+/JU67WTbGffl6va9dAZM6I5LiqAU2iLG8BSMpqCZPbPjiifp/x+TCYWPjIYik1O9s0MKHL8K
mGsLOC6Y/qmyBaCNOS7GOl8VHaBRnvXSBZMy9QvCtlltoi2iraPgBuDKYHASgODXwjYm8h/kYFMA
1ATgdb7awDiZfOelKHvto6Ag5/kDE5svnJlhaZy680P5EdpUuuEPHQ9HzzZYBiio3NSURF5ghFQi
DrMfHi00wgbxrEKgoW7SeUP5pLA8BT+6jYVlmjGcMRkOufqYFyWzhzX9Coo2egPXHz2PAa+0orqJ
ESq78kRaVjJubxKTvtgYAzjuiF7AbE5Al+AzjsWmzgn0EotBAxRl7vTj528heI+QOddz/X37UBAO
JsPdfsbKr2n6br6NC9dI4HsTpIstjJrBPrknILvx2m9D4qQLmc7cxfRH9wCXNVbbbn1oI7F5NltV
AIQ2Wy517Jac58tRonjepn3A21oclhyLaVQKdargAUxxJ5++jN/yBw199EJH7swzXOcnTvClwxhB
+JaR8SFqCW61TPRfDKCKCsj+V8AZENETpDHMLrdL8MB0sNLOpM/M7nJkyv7iJTFy+1Hy2LoJeq1d
f92v3LVGWg2GCKtmwnBvLVzDAUOwu1RFr3UGtj8gjP910W7mQ1h/raf/3rgrU+oatqg6a5PMFPRw
XumckVpze7gin+v8p8aX+DbgaPRUedB1mNYuTON5ytmd6leXdE125kwwAk1yD3QvQROluLSAob5j
+YpLtyfJZVsraFBoiea0yDNSBsijGAVfnTa2SJPBkVEjtvYBRJudaHkhjTugRezzk7hZG5RtfD8A
ZvxzMOm5sphXtTTpdMdFaEK0oneI3H/Dxb+fI5XOlwGqqgXrBpr0E9QnmnlcchxWG3R3PVLipuJY
W13TIxmNyXuz/ecbjJZ8SjJE8THXU9gNQ1WUTTz0Y1TcFSlCjs9JK6CTFBHWgH8UKPQ1691EZq0a
n76/bDNnvBq+RIWBh6ec1q9Fv6dFpjM70xcFoA8ryba27DCxa0IOoX2N/gZhJgKpNxQlThutf3+M
kCp13q+LQmQJpfnaX0WR9ys/POBIFy0UD16UWFwhUcvzd7v0++sehzL2GG+txMQCbdRX5iEU8lJl
E0nDrCagE21/GIEQHXeL/aa8dMTgk4ZMblkR4vceH02loE+aYn5E+0DllkhdjPNrjHKELf5qgkmo
TANGcrrvvr5fA+g1wI/cDfqxPTooCwKZddnFmEahXP4a4Ne7sexj+iBeVowvejjuUID1q/V85TeA
2CuyIE1FpZ+LqlMfjM8K8Lwds7jRJXEM9dWgvskdHirkBFdmwCwR7sGa3fupcmQ7FNXMIk4SlI+e
X5KGx7Nm+Re/dMkotNsovxQgF+I7o88YGl/VNs3CcSuYPkzynJYneXWWiNZOrL4fyTkz6HoJnFra
y5oFtnFeIV0dTfXldSC5eA0cLyPazGu9FVM0bzN9U22ddzALlMvlCqfTpns0xKRkgz+EAH//9Bxf
FMRMhPbW8tieFmz6F4ytD69ilAmPrthMvHOb1nUnH/1nok5Z5aicSAkWOtkbCBEY0qXDxKrtpdXH
VVVRcw4BuG9sSWyhTkO50w/j38b8X6jOL51JjzuHblptYfWA2ANFAbPyrv39aSUE/4HMKgrwE+mH
EXh13fpFtkBAkJYUofpYt2saBgqpn2VqccGYsW7lqjeCC/WSbt8NbqJxA4fx6XWzXCgEawA+/vz1
4vBOPbMudF2Exg+gKQUN/kp74syuMxNCYroNmASewK4weqhfmOdTaLJJljNdbG6rLAZezlBzQ22H
fWDA6Nmf/60YYakAvNvgXEw8m7hMUkjFHMkFLFn1HCi4NmPoA8x+nV9OI3D9H5NdFKgUwFS66Emh
iWw7UcpYjFNg9rLfhQSue1V0W3XrF493NjrcczRSDf2db6LTMF5dbRjbg/aIM8Xje6au153rTa3k
xlxNpJir42EnENjF093Ni8Wp/WoomR81qKssHb19wKt2wnO+owzq1DeOmNP/5bGT7rHpRM73k7yl
58hwu7APaIkuToxEHmQsXrNUULMwV/nHKFCd+tCWfdRwkSGJUUmo0FPGBUlRsZ29EO1rMUs+76X/
9GV5Glhrn8DMMH9liWksGyoqb4Edd6Dp1fe0ATEzw7d571jtOVGKFHk8yQrtOhJkHQMGPadI9ONh
LzPhaGbpTV0cLOPX6UNN1kwoft1agYg650tqkpxWbpHIZjMiodmHZ20aY9YVvbO30XBqtriQ3rvJ
Vj6vTA/r8uqtKuKVmFIFXj+E1/KE8Zj3ncUWYumVaJIi09+4pOdhI2BmOXmqI/5wrcOhb8ZPJn+p
DHAPbzpPdFQJcnFKfkwkH6Gz6fi0OjotE+PBUl45gn7NFnQ+de5UqS+KfZ015hfp1l4GNQHEJSD5
EJnZbrtHJKxScql7chq9qU1nZ4usbW+HrjiTYhCbI/i2aLMEthg8WMLphlULV4wFP3pGBKhM0KtR
lCF5KLAFerFGYSQ9QmE1lOksWyJStuNI3kv0laLrm7mBFVkgix3KjEzbb8kQpZZNfmizFx00KLVV
hqBVxRIFAvQllQQlQnVYa50okdLFsCcmWKIH+xhLXVRgFBEQ87pgi4JuJR0tmma/waYQOdGCBKLY
SpCt3vAZtH7r3+rrOEM0boiRTXdaInLHtNWRsoBxff3NaqV6ZszHyopwa3ko07h1LjVb6Keo8tyc
b3RD/7BNKJ+idTvoteXlRljZYTI3QLHcvREIlIfj6hmp1NWhD/rRWleJ3BMgflTx0E0gT/gLncpA
JW8OYWm3assfaKOaloJQalLZZW2v7hzdcRunkXwtEtvi8VoAuBaMQmgjG8eoYpVGnOwa+gX7TAGy
KAkZzB3m/IN/TzTli8quT24EsFYUvLtecWvQaJnIwiXFFNzFid+ifnsV9bV5FX81Yu4001hIXnqM
ZOcbs2uKSxkvx6N0Og3GLTe4XiqwMwx7az+Tl8MQ9btORaHdNgRQ3+AQuSfz/K88sFmY0iK6RINa
Hth0siwVedDZCs6DQNjKco/F2Kmm+sD88uRmJsePXhH8u2clA7Zx6ErUiaqgJ5eJ51NQIg07KQDr
ay0gj1KH393YlFHxrrdilfk0w3LefufxgbpvOUKtspZfE+NYtALFJ4XTUQLjx+xBhBYPjjxOglT8
+Bh2QCy4tDOZJqDzbX6MAMUKmdJVwCaGH9d/3/ZcmNY2pW3l3UOxjahCR/IJxeb4KQoZf+tphH0X
61QbPSHf7QfdMzQIIssilfQ2lF4VkAw6nJnLURYst4lCvSZO1MgzV37fdJ1ejxY73pLC/voADqMg
EcYfN1Pnps2+VgIAe3znjqoCAzWTl4XmDYCe8gZI+M63yHuUC17QjfXvF4qjDeT10JFah/BjmP0e
owpmzqNgE4mZhPSj2IyC1y6GHfsU1qsGWnDtyd7eM+mdXEpMOMCS4Kf7riHg6RlwHeRknn6A+dE0
hdd978KkPtYseLhk11bTyPQ5ePYxHLqL9b1MJrHwEN5jSVg5zXiXmRGnSnTjDLpRxymoJjplZ8MQ
nPJQZaKtNWWWySHAMX6EXTBH1ovgdlz2Yy4WXuH8lr4fFK9bdpnpWM5gk/5VN0lXFuoY6rvanD0E
mpMr2XBIIGIYCHmaGLEqSSM3mI59mBh8ntZAKMtjawA6HkdyQI0ra8utNzJe38ysW19wcG6Nfb4H
kwgxrjJYkYNK4tkyKYb0cawW9x2ho/VMFw+DTgyILjXtSLjR19SK91Dk0ZM4uuDxeFWBwR6zhOuF
5l3CfEvVNAnoZWoQXn+9g0CqQL9NubOMkg95cQ6i4CCkAor66214J0dcZlMCHNokY5wMyFfSF3ZG
43ij5aRK/bqjyRqpERf7dOW9VPZ3mBBQD8SCjhnPxtqqAupxKhFb5F+d/mHduq5l78M9CHroqSPH
0ud8gmZ8uSCy9gQXMcdNcGr5kwOTHmbltOJAAgpcodHvsNn5nmHu41SaqkM0Br+4Zs6dzM0Ekoe9
xm55M+aDteXxTeHEo3JFrg4ranFrTWl2Tj7YZm6IbG+huZjgeC6ZCj3reFZZVTh4U98lxxm5jSYK
mkGvzrgFJnFREZtsbelsSluhTDNJ+QfR5u4/T5pggwSXgo0VdbF7OfzOwYJZ86we1OhaxHlTX/iZ
lI/lfjy7dLReIIzl5FQ/6NLw2XgemICy7ewI04xJN8ffP0K6PHwg69HT4w/nJCwWuzax++96ky+r
Cce2oCAIHlzgoNK8Z2YM9Y1CmYkpIkjTe0SjA7TxwVzCHm8oe3Ky3RiIgER/d9lKBbglxAuU5dcj
sJaNPkOURDks3wjunMIXCOxp2NiBxERqvzOKzX6BUUcwIrPAhECfFfA8BHkS38U6J1S07P/AUc5F
HNXLX1sKVCrnTkFXBVSaiGQejWdz17v9cbD+yDvgjhVQV5FkNzan+BkOHc6TDkfeB+XADETQ1Skq
OIYB4uA07dBbv2czTgpl7SgwzbN+HVVAYgGaUHW/PUENHG12ZLKZnerJAgq8h1tJYqsVrvEr+ioD
gcdbzCVwHHBQnZ5GrJ8G0+WZ1LrPkafEpMtl+kse1TDaBRK4A5OJri8Knduj7WQNtowxmfkmIT7O
HayuLcan5vAH4dFEgFL8YSugJhWqo0QL6FvpMg0QTCwoTLmpLHHjsvp1mLvFOGhrCd852Vb+t5JB
lfZpXKi+R0cagqLgms0BGn4+uAs3FiU6e0K3oXwyUqEFGn8hDfKGnmTTQsLvKxj7DJaYPmUa72lq
izMz4eh6uYv9fNST5wyQbJMXdQFtYL8n6lEAeFKUXZHnVeL0B6oMj5U0+GAgxzu4GI9CrLri+mEl
s1f3/qZkxt2g6Q1hroUXSVnnHuhwGn6X2+ZW+8+S8uyspXFmzDW0wWI/jURHccN+Xb4/xtguvye8
KlydQWaYUqKD4BCK7aDgzkBdfpmV+fvbga69iUuUv7jCLg8k5wisvmz0rZca8pJJ2EOJTi8+2C+b
MFEliPimEKS9yxgnxxWKjmLBADdZYvRpdNTk8n8a5gZBnLQJz52N3At0JUDKXnAl2WrJqmpKG7XZ
7z7FVsxmSK8jkmxQmOcittRkQdcpZgRvJrhAjXdXcyKKmGEpSIzxAdd73BINba680wjE5BNSN31W
XWkzarmv5W2ZY3a5rW8vWA1KxAr/Rlzn65Avu8iQc4GYYc+GfqXQdrswilPkE+DRI/5vN/iZCpDM
pax9I3+AeQp+2edaL8O+ev+/vW/DupnoMy5RIYWuFgW72a2egbVu0FAuYpT4EKX8x95nbCjj6HXZ
WT+/eRYF8qG4CyPjiLJ5j1v0rWJxl5s2hzx2bSebCZHnVKXnTlbVIqO6dwwBKdN9FdvhLlAnFxz2
kgGqdJ6V8FAX4xZbPGq7Q9C7xDZiF4zzaeeeoAXjysM8JoGy8wWdgw7CP90ywPo32gMlh7ST6c9p
K7qk05bNQkFAwio7eaRfnlrUufa031e1fO3a+E2u+WFCUb2F2u5INq98oM0a6aBRxuIv377CyhmC
opK5aVm2P0JKcciSgRRh3ZqT5iTsWx3yqRjg/14LgUUe+ZOibqRUFrxCLKEvE79j1ohTbms05VP7
iCvrg8muZyx+g/JdoBZGVRr8WtMw6b9JKttpXjF1uTn8PGKwFCBj0N961Np7cwIt4flzYJ4ZDQWw
a03UwDorunqu6pbF7RWhcAV0NCKFbEWrfLpw4md2LpIe7Ay0tG16iN/EWZwoCob3P/lc1eEAd83V
1bIFAXENQNDXrF0KBML7kFF1+BnF+wVCumjPZ/cibLq9y9/pyLaXeT5JijDybuOXUrbweL7n+GqH
wV8OTarB6KzxZf2nmVJsJFu/NdgSNbDTJEQP32XtBHWah3NZh1maoatw+WgOX6gKst5gAcoekQs5
Q08vTbQ65dDOJy0/IX72kVE3zhuXStaiktX8YnB072qv1oakKtYEnRS07jcNygWg+Nu2FBI85Uux
ih5cmDxgSG/BGvnuoGEBX9K0qYM293CQr5V1DHf8Tch+HXxOj1NNRDCKxWajzhDnyRuNaQNkMwaF
vn6ex6QWJW4G7nolQ6DRbC9PcsYZUEsT5Ube+d+k0LOOcdky6A8o/2rjk7aXfd2NkmUrEbwtfZ9V
uDIYTS6J+rie6Hm5Xx2bW9C6AKNa/JAp/dVfZ3Wlg4V+oU6gYZss1W01UR/iiHBV0toLpLcx3x8L
z7zmFmr+4q0MmEXtrf1Vv0G63LXqC18RVaSTjpujjl5ZB8emMYF+vLQwBainNItHNtszo60Obie1
pxTYbzORoKo3VJub5RUKs8ioDHbXyKrToEV7fSzSqWhYeulY2HC0zatmiOvBRDOBeoo5D8rhKRCm
tnvSxL/LvihnSbairt8mgHD9CaW3HOsjm1TuBz+fcM9prOWUTq40NdsOx19sh+amv0Phm6tBNVVH
7C6N5yqAx60T46tyRR6ajzWnoj9aCUqgn7TfG6ENlmM14jwOsQWxo9nl2UigIWM7nWhcCLgm9KxG
1TnWPZs8Uak2iiw7EM5EUpQC7GOl4orGU0lnr1nvXPHDxDLQpmXKHtytkljzwvQgjd7rs/HPLaVK
y3Bt+RcZ0gypO2duheyX8ImSfOJYGysTi4yu+DjIW2OlhDDjGqnw6K9A1jNxkV50+dqdPntE6lHS
McJQuevW6mMEIv5LVgtIDyJrRgn3y1N6opKVj1JF38Zu7uU+BSW8X9qDYzTKHk+8mqc4SlKLwS2k
awoK3lBVs6wAOqGjyZEBIljsrJ9UDDj0sRWNO8DmUHmBffjMev+igDbVEEjDY5LNGYWRU9PylDYB
U7Eytta+F4UpB3oTY0mHfJO4JVqRuD1qhc+DcjEAqVr5DwrGJHacP910sqTKtES/2sPxbIBwyrFB
tsY104JCQg1R77flJKGdrzzo7qXCh3Q0Q4jnVCzaxbKmmEuuRO1LpqdAKKOVz+3yw3hGSFzeKBIk
A70WsMdoGQdfuvSJvlA4/3HEMuEMYopc2LQEa7iIQKjTsT6EzDOH7NU0E18/HWNe6I4t7UrfI54j
M8Auepi8CqalWg3cA2WhWdxQDucmrhSC7v7TxrxCxDj06lfKzpkA9ydcYtv+CEcumNAqWiiH8hgq
y3I0Vnxw/AKpeMhkPZ7ZgdrCt9JmlR7oPEYbD+VB39NsiA83eZKNkzZVEEbhpxGBmjLjExE15vbI
VgOOXBtvUmn+NrVXi/d4aRedURl3P5a0MdwhpXPveU0AqlCG1HgGkI71+uzRGUYJYrwtAOeg7RkE
r03gDrkOjFCvop1jDZs2mHKDMAx3vB/d35m0khQlFvpuwv+K+IsGGp10AdHgnkX7+UzoZaYoidSx
aIx4YcnBut9jm8YMA9asXoqKZAP5ruYsgeSlTd/nfx6jLOFduMZHTDWerMIOqDbM3D/vf5u3M7um
F6Mj+U+Bo7mHXJOy0DPVZ/BQVy4FWIb7UFbna0bASBh+BgbHjBiSqxyEy29a/pGCmgJT5ZbgpvQu
Xcvax3qat8knUMy997LO7RA2ieUki8/Rg/7cF1jk4SzQ5+M9Ff19a5ILlTMyB+k/esoHHu1Pa80+
zBUrFV8cCRa7GyTpBhe0PpsF2Vu3R79RMDP0yT0tqXxwiBjy5HI9CnpaxZR4LvOx02Gt+GJMK4b/
VcvRWXFIzZR0eLk3m35sdOQk0SoosBM9UXgjVKsfvW5jaq8e3QXgkPt022WZxvc9Xa35z64wqPT0
dAKLsJHOckygRgtTJYXM8qwzAW6OqIHlbxqQXcrJG39PiFXQq1FIfzBBJxOd5xsaRhSLsSN5C0EA
lgXy9xlSwlNCTEUW3xsXJ+DTWJiHW1kwZXfufnTSSwDXFG96t198fMgPirQOPcGN6P/y4/vGJ5cy
rUbrCYfO2yv0WYhcHbUUKs2sHtpma5HOjoC+d74LtQuVaDiAq/qAsMmNOvg+QJG3OLP40yhHH7Ru
VR163oqLZ+NZmRT6gQzbzxeoB91My/wYqmPV48iibSuPCPFBL6m/MlMpH+xgDbHTBIIJntbJMAXl
4j2PlwK9GphYuoWk7yHzZgxUYGVawbUxV8RuTV3FwJcPkpMBetJ9PhreA470YxgIoZ1XNH/XioHV
8pkPXLlOudT1MhHPAj5XpZFErdblyx5V4Jdll3Jo/mqeOK0Nnx6vciuSsAcS84tkdu1+tRrPSdV+
XoPhpVCPku1+M1jqQ/PxODxKUmMYZr+FK3ta95D7KCyA9dIegoyC22jEaIYourZRW9kWKABKPERK
Bdj4fXuTkjm43RFM5tNZCQflOeyzoX8ZJH6alwVltJCnQU5GYjVrHOxCa1LY9h9XlJaw0j51zc0f
pSbH+sy8wtOZKWqln6sxW+pZ7eBwqyoqcaHnzZuUqUMggJ4GIh6HPW7Xzd8jrFbYo1rZPVKhu8q3
QPnKnXCuzZoAPQgaRMNVHFAqqN6v14Cjh7geUXMwc/GIsT/ByKam2nvNRgKRQiC1nFf7+flDTU/X
ErPfR/2qPm6nng1HPTrnyw4zIcUUW+Tw9aKqaKIMtrZwK+GXwp84k1EDxNZjZfZrLV95Qx+XSKXx
X1HafEOIQILtCVYRtI9iXpC0ANSliDkW6/2bOYIKWg1ChQ2WJpSzS+ARN9IQ6ZfvB7Y2RP9j4RJT
lwENyLozYQkTLqGBS0IwOwqbYjG25Hjrtp60yOe7WYQkMXLyu1RzQBxtPhIrpCKmQ0Gxkl+J04ay
d7ni5LmJsX1XJWfOkA5j5HuSfPPGF5SatbJBzXhFZp56RJAcG8o/sqgDt5A9woDHTzFXlQCmKVM0
qfUpOd8wGBUBg07W+dZd72SNIYfGBlANdPRQrx0WNZrVvzvgTdJxqDKnLTM+BsXI77egBQ/sk1or
uHa0XYLuQt4Q8eDZob9Lpk75C3bEdpKWT8sI1GVqQcE44t+TRJvQOX1m+HrZkDrsZdIXjQnt6ZhC
JglN2BeiS9a6nP6d+QP8kyR13HrP9RbCucYGWgANc7d6q3MpEviAAaTlF7YL94foAWGOjM1/6A12
G3zV6JBSe7mQUoQ1wGTWb+8JB8B2gen8ZSFlDHXdE76XSS10jZ1kGZGd1PECeK5lme05XWwgTh9S
xcQMiEd6pCKc1K3MQBy+SsdXyG7unmQ+E7rhxrsZEWz9izwPnbgtziz52TzhDLG0nJeE6obV8WJI
ZIjPfzl6rVsPoEwYGVOviNfDlF2Nbgvs/P7Z5Nm6I3+59THKPYoS2cTU4tdpt/cqUSWZyR4VPi3s
kgNnh/3yr33TvBWr6bQoZQ/d8MjqogwZuSn/lGDhBI5ScreRXunajCh4urkFR2c9Rl5GaXNlP8Oo
VPEK4sYsNrydWES4Skxi6pgIjC8qh2ACj4/SsQzXheibrkjjsN+EpgYvhLM4ihPJKwms6BJSwTwV
Z3X1FHizanA1FwGnb235YGJdpUnG8A/J0H/FT5eXQOHO3gaYPQ38VVYc5kVNUu+pqR1UDgvTEA2G
ImEIw9gHzUP7ooazaxqJwoCzqSz2D2JeOkgqQSwijsAZ5KS4hY+6eLt8YG0CbCowMZ1rYAmSUyjE
a5Q0zQTmcU2Dr+2oGOCWLdyCg2/DY+xnUqYob0PzAW+7FxkHu3F1YUXzi3W93kfb9xd5msNZdSKz
XtM5ag4jasEw/nwqMlggHqUDUd2izMcT6n9yOYtBix/CEa2FWzsCnWSgWYU+5SfMpuvu/EUi0Sfi
lOrYdnbbZeNfpCq1vTeqnK4PP080ZFqdSr5PSksmui9JBvGzrkN+0iwDoVahZXxXQrF1fUFmadNe
LCCm07PRsq9bB7mMuedwVQgwX0KYo2/Zp4Jbq8S93JskJ75QP5stUt1NkmexI6K8zdRN/X0VoZeR
RHfl51hI83gpnzXIo2DpspCszWg2Rz5r/damzBr/Q/mmLcexhdle5lR408dcqF6OXanWXrYwzTnc
CXAMCSkrJNR766D5V84/4tqArf5fi6/ZNcNBuicZo8HkubRu4K9Q1P1KOpc0vxNZ+aYr7NYsV/r/
eKPwZlWehHLGHeuxpBGMattP4uPH/K+UFFL/unNNrXwA7SkdXtY7usbueu6Nx4KxfRV6aYK3wLFo
KjA59JtjK5OlyT0sCAQ51TBA86Q8NSypV+p5PNWbYoyYKGGDaKDsT2cRFBSP7NfMyMRK8HRwFrJ4
g7fwckaV4mbceDDWgN3z+Zx+GEEH8kPj2i5BHXO6BLtCT9jXweXxoi3jHrTLiTfBAcTbuoRX84mD
CdfwYBZDLLK7UtVBmYgYgoIncvgztXI04ol3ktEdJPksrAHh55nDp4Usqt8YNi/7AuLJMG+3VGcT
scF5X3S7kRY59qMwfaMG56M0o7sEx72cAfaMAzyqKA/jloD7CXKUzd1vbLLVE1zKC2cONkW9umio
rBUj64Gg3MF9tY5zcwWpUQK7OM45wfdaifTFXHmcFTMPVxlAlc3JI4F7wD7C3o/YU5Jn5k2YOHgT
EMLwKGkFwvftTmBX1jzReuYv+FHeMgXZOPmgzyhEIPzWDqSOUsjnZTwWFZH9tNOHX6VMtmJ0I0JY
BK3/QEC1cZnXXsVr6wPRClAib65PRrViilxNFF4k25IDmzY9lceJ+BiWoxxhBsRTt2Oqc9iwIkKZ
uilmdJBQBhuORmsz5CZ9M1GqE/kdyAJY2JfSA/e/iDJ7rGYokFDBklmIcp3XUlnyL9T/xcB+pK3g
itUP4PcRmNsPdxTpOUWB+Bfe9GFMZKwBnQ2zep++ulylD36iX3NpJ1bKtRVdIM/NwozxHA1qI1YN
6u/GBJ1X+fps00OvJBe3nKbMPIU8OEvBQyjG8kg0SAJluSV5BjPtzTTtinKJw/msLLoHw+4e84zv
4wuZ51/ercJAeRw6oM1RyXkuJJaRn6hAtmz7lcZw+b1RnDc066kKC8SHT62TXPox1/n8WUHIjZ/T
dAvlrWQY2s2DJr4XGMdg92Xp/bQjkPKkZJSUHxgyOSHctcZpEw1N7NIwn5gXkJ4QOPUrCAqETGkx
qjjC8SkjdGuzOK94PQchto37iaoyrfhXDJGxgdb+c/CJBdv6xbo9C+1hqC51f/NoBvSf0+9kJvAr
wnWcvi7U8/LkQTNZKj7Cr7s5qvOSv7hndce/H7/LZkfhY925YZu48z/P8zg++p/IkoobjhHWKWba
aj2A2lAtJ+ks8ltYVHoHJiWYvPG9nHeJLNWBV4UXRTX5LGpIrAOJmDNjq33xTRdWMZOYb4yGWa+s
ujFkLsebZaqqKl7zLla7t89YwzV9FirLqqUB/TZoxoWGgn4nmNx/iRTDDI5tyHOql6tmWhhIV9c2
I6tpmF61woNhDmalYsK6z8n9kF9JO8XiHI+4tjLmOtXvlF1Xo1232nYqGlb6HichBAETEUfHcgVF
ChO09XlGhXOmzHWdf8MkB9NPc4qOtY0t7zOg7bQSG2PcoG+paC1KPGLjniiYB5n7smSFSDQtls8R
D+iqm/lB8FHC3Abi+BM3TdSGQq8rEupi9hQnmtJcBPUaPW0fKh/ln17ZuqnMt+svIKDK+x33V3S0
zb92bPck3mMFArqVf8xdK/7kvkKC8UWwDHEbz1A8r9/6DoCV4Yf78GuQUYh0QoyF2iczcGlEAF3w
a0Bf4W1pLH6BQsM+gXOydT9vlO3aAr9J52R7rqftCiyZOOyJbcoWxjJhNIJzD0uHBxv6TpLlBzXK
qFRzXUAwbRHGSV3jVrfk299GjLT6fZ4HtGlCU745EOW3W1qTntLSWohg8scIHBBzJL4cXCETBkem
sQ5k0MMDwmlcCHybt/PrapB1+p40tRYcsmY4gYTkbdfU8S9E72LvE7HJfoojrVNYO4hVA8yJSlaX
nuI1A1HC7O39MMFzENF4Rd4pOLs+/dUudivRDN99F8Y+t7mkf68Jyx6+eUp9MAlumjW23JwTcyow
FpIpLWZ+QkjMyEaPphKbCJMXvWVTjrgrPNrnHicSDDfcLZSnKFZ/FoFQGOs4i0Wj5bsxRkvR36zH
bPtH2eTChtHiv85QzPPhh2Sh/5kl5l3H5DEBx10jM7C7FLN5j2zZTGxdosMNZG+mnT1r3Ej3+GJv
4oy++P9Q24i5Q9gsMKqSms5CuH0I0fOag01HZ94PnDNFBmQibkEuOrrI3YycqNAmFu0DjxCEU66R
NZmK45CLrk/qfMQmhirWveI2ozDbZenQRQOxdaDSnYPLZ046uGhMwlNRNmV2eYRr8nUEtOhfQtEt
6DOzl+X4p8HcX6+yJDFojTvyx2WoNSX+OHosAP9l/nQBU8ZJjE7lVM44CxQJtYThhiF0gANZmno1
9wNqOMDXyfTLxy2hjV9DNAe2xRPJ3zrR8YN34L80iW1lqeI4J1YCol3dUBJfr1ySxsyx+vxDk514
eCQdBarYUEnOA1QhDIg4DLiWELAzsL93k5UxzSnisYI2UORpDMtzvgiNywuL2E6gsuWn6C/uLA0G
Uehl+KHT1yS+9GEEmZrws+qP64VHVGmlTpEWuGtozihuCotZ0VYR4AN9auPVXAQ1xZWme1UDtPEQ
syKT2inhc8ErxfAZhdYVjIeqv4aJA1rkuCTm2Uq1ETRD/CzlKUHifdJ55uRH9LORxRvG3363xU2L
fXoyP3M3t+XGvlFAXGGlsKjH6nwDZk8/h/cooGMEvOC+lLfdyi0fZZOKqglFrqxpON+RX74ruCQH
Vu3VwFO7JGOjQJDKBYSmNzInYLNyCNGd+NNS1CxwQ6jX8s0s+CL5mDlhvHI1XuezpnCOxA2kYkOX
8oFddkdSjEpeYw//ziJUe5eVcFZqb/Li7ub5b+rC20Pv6CUsst0gMcpbSaL3sAiPHo2Yp0IREv+q
PWFaeWQKqsHRTKjA4n1FFGcW9IDNI8u2FLQFWNE6RdsPxxKV9h3rRcoECwk/puyzVUHaVhXiOq7a
36RXK05JgR+ACCHc25oLJal+K4b9lJUCgbX66Fa4Xlk0Db/tQDYhTfNJpHbw/+SEE6IwUTTC2MA0
BPI/t8pTLOVMoVs8I17ARzmslhcex1rGbWsOugg7UXq2bcdR+fXsP0f/vxL0YI4y9nzMMyG680yd
T6YA7AM9weB14GFCEm4fjN2fGli3mohZHUKeKoRPRBOkAAzjsT9O7LVEVQ8GzEHivFd9ldXmi1Bc
jlFTTQYuSbH92aAob5NJOtFTosRaL/VwVsJzVheZJM9ug+i4lWYb2IpvyPrZuKpvgugh2j23O0PF
FX/Y1cKhusH1AyuiOHEk3Jji7hA/y7fiZss4MO9jQwyVNJp7GA6qHS7hCOXQWwWgNwZQAs1MOhwM
AYZiJeDu65mzfabDU6WpEQJ+JEtpCMOPl8rMKQLzNcifuHHqWaWKvKTjohSSCyG0bgzGZUijeFOs
C/vStf0gZQ1T6CTRf4OiqSjb9DPCduE4X9meoO2C7jBwOYDTsX95u/Hgw19odKTsr1z6O8QExmM+
yaONB6Bj8LOJbm7MC4FvZxkCQKxU8lmEIpdzfdK/35dcW0I0OT7489dwGztWEJpXuSYfqmeK+3jb
ypmuf3Qu3dgSFhAK79DYljkgQ9o3tIszHVQ8Ok39DT/pPpiejYAjXZzca0dMqIUazw3b5xmm0MJX
rxwRyMH3x1uifVgbHMQ4lyHJeFNr1zA3tFgEsoYR6nQMeXFyKUvQF+quLcQ4zF15uCCSVwpEgVQq
HIfQme0bYGua5ZHmId7Q5JKdnGFriQVMKNCZ+DlnyawWOip0J2/xgougxcf4qLJ26q9knNZkcbqp
VSnYJD1EbQwTvWNiWKRU5TgEjpPTxrVGksLEsR9N/E4+EIHsRsIQeVIYW9ICmgh+8Vg5Spg17/e2
qPk3s7QESCehXBumDUlqz3rCZIkDXBFB5IfOY/0NcZ7Vy9IxQkoNR6io1Bl1Ykb6QgY1t8zWBekW
KjATJU/hnQPfo0YVUUGqfGQNC2DFR+vNWxPvOnmbBlmE+IWEW8AirOrI8z9IeTOnqmpHwtArpuI1
cj/P4h4edWl83E/tBoXbQyNXm3ymquvSNmE8sfm+6WXDuIvT0MwUqGJ2iKZAwbcbVth7g5N0JmtN
0Y73FwvFEXDkCQ1ItQWqckAaljtsY3+pjXssdeTwGRrHQykoVaSkCTS4hNfAJfGx31g2f8DupacF
u8pVvlygX6QhpVHByMhZ6ipalkI2GwFYdy4kGWQ8/3jdhpCLpue7yN+28xV+J47ixIuk0MfU1s+k
xupeV7i2yYe6zWUifThIhZKEeyBw/Z0PJ0pBv6uo/Lp0zKTFTTzJkWhmxbGb5ByRpy6x0NgricMw
IEatY8Ri5VGGwz7VyXVCHM7TY5h1rRkMkUvJn5ndQka3/ElWVBtCATYBYPqcijLWpEpx8Jn/X6uf
lXOM+zOjX6Ufi/AaXTbGrcOuEmTpcr/dTqbb+G7q2GlUI6ioAFhG0B/ecQDI9Xt9L9WMPolpATdk
XrXWgF8aUWrJme3OQ+3Z59dgiJ3O5FbYVFkg0lUbJA8fhdWPUFm2A7vIOQPklXPIxPU6UnhG89vU
gCCh/l7h3nwCrtpWSyRazpA9/MfkXDdjlbHFFxWMLfeOKNHw7jtnUjqPAuZaDgBBB1DzaNA+uM9z
4RB9QlLj+hQUNOJFI70UvlY7dPVFr6y9zLQ9KmYQWpq/1dJTDKBNCSQxnzOxiNthZ/q7QCIPwtnW
Ib+fGvhzX+8HPvXBkkWHuqbbsNUDtZgoWFp/vfAB1l4RFJ/oGTeP5mGRGObKYnokc0QCAsQBWOEr
hu6+GnmEs3VoIdn1+yawe9ieXpzCVDuYGzGmuqSuJ4tovVJ7nNtPvAguZKz7MSQE3GIg2rpYBUU1
p6LcH9tRo6R/EidydgMDIPe1T6JA03LpDYKJUVVAGVURtI04CbSnIjewS53Mt/skz3LbZm1N5dSX
F4QSuqFeETSFaolC05/7pofx6/6cmDUhJsVqBWvU+DcCHA2nzo5Zs6MPMudA/Uvu+9R0w1SEh4sn
0soP+OzHHJkNhjd89WU6/6kpDgE8xnt+KTxDMRZSqK9GFgfYUQ/Umde/XqUiKYEJNI0+LqldVWby
aLvaOauXn7uWHyx5VOosersmGgQ8Kd4Y2MmmSczG9vEnVMuyROCcsT4GDAE94uhWX3yB5oogZPWB
dMj02xjgEQySsiId6T+urcBhrF+kot75E0KrK1gulAsrzqPf+h0X98wT9yEJDQt4eZI7PQlY1JJO
hjHwGFt+mcb4o25LCwtDRPdB4iYp6ZVYDxpvsvZaeHHNucTEMncv6kMt7Y4Obin4t/ciSa6UX615
XTUzq7OFigb84Bxt1kvg/Y6aXK8mMT1eScR6qiY2LIBQB2b+G9b6MNgzvNYnSi7A7NXHAk/wn0k1
HZebT04mPH9hZDYgYv00FvGw9w9gcmESUtuY2943pPw5+npI0Zj9bKcEs1KqgZ4uZh9/HEA0CVzm
fQr9xF+y0AAXFXLWoEuhhs78X85zVg5l0SUal8Ykd7kUMYjWOhxKKVyp0IAnog37dXbQGNowWl+q
YWiRV5gJ47MFRuA54dt9/Czl1MEAzod7H5ERcY7giWEeOmHe9prJOra2iCrkqwkCV7RgB9CSJONC
mNm2FHC45ATMP3GbarII6nj0ekmXpvkU8Tgl1zVHOXOXvphMqkyhqT0Uyu0lhNNxWpYkqfpezaEn
mzDGSTBN0u9wfFJm7qPAoctkKfM9t6W/HOwMcYw5q9IgJkDQfya6OQjmaHO7hOlD4ZpdYZuD7LE/
2XUfjkpjYMGAXa3gBZ1HJauxYYNJCpHVoQ/2vvsKrx2hEVJdVzBRsvMeCP2Nf4zK33NXETw501XN
gLW47pWkcpfd0apyyKvB19ojLjgQF3HL4iJchSqlfq9JD3rNgMDlttfr7MilYzPnNvKcj7Ruhq+A
mrM/t2mOqu6UUHFBjeflPH8CmmCgrbgUVma8z9JiLftXUyQ9TgpRKg5pWvFmGsLiz0RwRZiADRzF
h/b+xZTcgp6Lt3H7rUAASiQjOccek1yAE+ebuNsvXHUogINT8K8MWvfEO8zToVfhfi9P6fL/eUSA
HD63EYNvJbpDazVA2KmI5rT52qSsRjCVR5tb01XNToIfL8iwKXcqB5RDKG7XPXuBcM7VcBuU708G
1cExR0gjVRsPXlBMhimHAxbj6A6pwoH4RtfxE6PqO5laRhMcDBjPyKGsD0UY8l18A6+7oVDQbvzc
D9MuFzHcqyMjMs/03e+kzg5hLJSljfSVkfg/22PrZ9YVMP0lzgGod3sXX9OYu5cdYeUhoVFZpMg+
aUK30KOltcUfLkZJFVqAazK3II3NduHhwubMpyzjfqDoMRrEdvRDi2fNVA93SQv3P5zVkbct7cZR
L5u5BgI7niuUnhd2GhB5QTYNvUnbufrqQpvsBcorFBEALIXmyegZ+JMQBdJ0XDqmTEnTh0OGXbSi
fBfMBupeOMPilqC30hijDpvTTN2fk2biS8sqx0eQC+bhfBFcfM0AqgF+XurhY3F8fW88dCi+mpzp
orBAWzrKnItipfyRH5pajFrZJR9VOYS6ZnZPlJkUFlzfYiBqcOa7bEh5fn3cqJ6ks92Y8Od3Ju0U
3rBaJd9C2v/KQx/471vGu4RKcAQS1zMh4HDhFZAPpo+WbjqCGcFZO7WCc+OKbGsCZDxlmfUQ5+8f
rU/u4q/Vn20WaHNABAEL2SCfKbvFeYfCyHYXU23b4Lh/3+7/vDpY6ihhX/tCRiURSZXcaq7LnvNO
Y622xDLq6ZcSsWbU0vLv7Z9T2oIJ1qnlBBLMKLbCnH7oM8vxtCWjHgAEzsbiAF+V9EdzVXovrnTU
5xmKTCUE6VefSBbbNSes281uBrWUaQ2rXLW7QLB3lv5RH4XMi86L1XypfuhrwQQ7aUvld2srNBaN
ok5icHImen8hApgI66Pcw+pSd7ZU2j1Sh0j3tcN2tQ1dI2goS3iBV+KcweT61/giRtd/PwfA0cHe
0CSvS8zWbMJxtefP7AsJGi4TyFxr53s+ow630xbhwsik94EBaqsGDE49m5igg1nOGm8u2HOaDo5P
2ppyQ+9axt9qpeE0sB7X4tHOVyCtDfolUg0UVaeYyZDvFHQjlaG7f1zrbJ6XF1vWC+oYEbDRydZm
JMiDtAKffZ2bUJJza9Rr+ObE8zFVSJxuzRVDuD0ttXLBn8aZHSsIdVC8NawgUlZeQU+FSJjmaszk
HfY69b5MelTi10aMcLH4dk4Cu7qmspXKxxXSARW+SGeg7pvQlhJdReKEQf+BhuHSVgtZKFG1UXjc
L1T2ag6Ug117VU+dpr+VsCGp3GAIOTGWuf47O/akzTCexPZNEUMUGV7dxMJxBq3GdPh/JHPj6q+g
80QfbjEh7lvM2w9HHSjWUfa73DshyI7+ynZPLaLYLLgrqVqCw8onkkMdfZt2yJplLxANIoFcuUhz
1P7dD9JQP8kEy8hDa3OX3aQ1LJdWSIEpQtzGeh5+/7Xk7rvdoMTnqzLNdugVreXrsVmcf1z/ya4V
xzPPpnLIv0U7zPAv8ByfVqpbmIvSLurlOBuyML9rKEFGGQwit85bquKqwvfCtfOMV+3O2UmDa+q4
IpV3gCDmpE+GtgSI43aqlqvSTaDQjJzcdnS17ci3o9xFa8LLoxY6QhPTtHIyM5hus3uUiabIbTq1
NAB+Zm3B0w6Fhtq6qvZ6ZyBLPWhQPBcSmC90maGqLfuraz/81HTwPV/iBfN1jOzGJvZY+JcElw50
khgxAxps/opxfDH1dby4/eoaeLBXzZq3qPuZTqIIowib1Zv7ZTrHc8LFbKPpRYYFdJackoY1bUtJ
P/QCsLocJXrJOosHrl+OGE1tz6NpP9ALUZTNpLrSe2MoAEIvb/k29kkpGBdTFVhRUJLgPe7AJGRF
ccjdYEK9fdxpUnOS9wCNrix3kHpLR8yeK5mCHaLctOBXrBDyJCF3KLCEiiX+3Wa6fFFT20WTivCB
MDlQEpMBvq2aB+Z/7nMbGPZL6mhwR/pSiHzBfejaf6j+IKjZcXhTmSNDU7aeE4HW5scOl8MkF72g
HRuuhcyUjXUHBzz00Y1L0MBwJ1i2PCbzz9OhWoGo12CGDiW84kiFRAZPbFbhLhEa/8ovyVteqbmz
ELTlfNC/0pskNmbIUoRAn3YiM3V+q5MoqDbMroK897KttvxlnAvT2/xLvh2Lu68Ed01peT2JhcRW
ob+PkM3mK3QK2ngSuehJKW7r/Xijby45jY50oj3B3cUV6fjoTAUlG7/3IVmSRXpLxV5POBhnUFGf
ioo91XsFm2ITPgCwvma2tcuphAuZZNr+1KIUJ1R71ikyclmNzc4RWMdLn8St4p8OWqo0dVBwPjcN
Q3XA7+ibo7ddDdGm1H9xNujnJgcDxgX/0ihLM61tH1LqqDYkrfJzVPNWmQ5aEWj4+1dCZtP+BajC
bC5eIAOnrOuf0w6DvV+hM/lV/62A/+AkCHyw1HQOtsvqlD0y7bJv3nnKY+fmEZLwa4mSp58hGSCW
yVCNBZilJuswJDQdBmTb1MRrSQYiNKPVoE5BYOeE6c3kbsWzX8kmBjhBtPurEzRXPwRfEkwNy4O3
VSuRYkBb8RrYbc1RO36bK6+lFjCLLmYsgQYqLCopQ9btHdvgybWv+AMuNQeBTw4oZsWdolfy0swK
VG/VZdXMSQaID/CqUPG5mJAOFf8dJhLQfzgKCrO2U0iqjFNyGMxsMYxo8ZyJ0KBzZIM5mdL8sj0h
hYpDKGfGaHBXXV9icwvzJjggyXgPMId0wxyiSkxPCxKt5dnSlu5xWTlyD3wWKkjnvNSgr5rvV0Jv
MbEzsmzIsOOAXVQHSBZ+DFH0rAUxeGFWrLSQ3bJIV1Vg5JfRZlgF8zcofd1MyzaTtJ7LyGjKb0fN
BEC4p0L56YPX9Z85MLKi320WKhuHZpb+2+NyFEqKoC2iRi95yAPF1o1m6MASXl/qKsHf27qiv6hm
n/OI2gkY9g7pfj+zIi+nn82PCnnMzn1X7QgVVnMFaNPWubFny8vIEVXmoJ07xODGwryljIzHvv4c
K8X6gh2vkK2UkmaX4/Ou0blIVXt89ppS/fXSEexwDk7tOyrKxT4QZrugkWc5EX7bUGNqK76gCBgj
As5cAU335bEw6qIfoBkCjlwbrOV/pnxIcbbW+mg1hGFzCQHob6rHLkcFgsvmdurjVX3Z5T7JQUk9
zc5FXTMaflMDiHwXFC1q+w2DC4eOMHMLTDyCtErxF1PLE7f++wj8sgHZp2Xmw0Fgz3WQHGMhh95c
+AqzEdA/K5Kpb/sJsLWMpe7CA/WpHH3rKcAIZFF8Qy83dtkxp5YYZVFMxrcFHqVRL3g42eHm+ijX
o89hRz6Rgi4OuA6xFMgXetgbPvYjwJjKp05VDmPS8wJ8rUM93/uhbUW0fAKE3LWdoWJHd/QiNSBo
UWKKozQXc+7APcJ++kRDkCUQe7zW+LskpF5cCeLZU7bh++KP5x2H6EiqIHlEPRkTSjzEvhtafMUG
P23V7jOB7KuyApGFol+f+tgr8PCd5wuXXXgFHErNK1oerogu7lqq8TknQbkrsvh/noHlFaVH0+Cf
+QikJ4A3Y0/7s5pdRytFwvdj3wRdeN9YU7Y8sIIozLTji7mD8QSZpb5mC7tWLGrirfiLZ4b/bfoE
NK5tixVf3kxCjAfEYSkqchXcUFZnzOI8R0eeOEQ9YZPyD+GeS3y/FZghjfhtKgDNH5JXjSAh+uSN
KNiUoL8GZKixd3w2DRCjw2R+WvoRVd+So42ChspZiPd9WpT+e2f//9zFGyQuCPLfEqaSemzYrkYE
oH+K7l9OOUsYZBSTxVuK7UT+qLbkS26wETA9H5qVYm9HV7SmVMHlkszGWI5FvGEdjuPuG2P2hqSq
rheM31gHlueOVFAZLAYspQQf2GJmtGsfti2VaRVPLbUrOUlKPTbsXIz6krOBFsk+wI4ehdRVie3m
Y8a1U4kHpJpVOBr8k8Ep8d6QplltHxBk+HmuetDeez4FdyhNnhL4gaC99XOnMlvTbR4UyXyCpHU4
v35+1lPWMEDVemWo4Bb0DXccftc2xSRGH4MUF6M2zibs/N7KXqokcgrnh8K9TUFjZhVL+/lru9Gt
zJNxSNNwcrdeCWTpE9CkowkZg4hKv3bAC4nPQSJjCZmozf+/Yv51nDb/9l/HCaPLqf/NBRawdINN
82n3kF3DViUn8YKcS76oFJhDJ6+LwSllydeVOuQYs99fLFohejDL0m+YtVZeTIsZ/qrRp0FNCrAB
uuVgFrdTqz0MtBWAkciH4Ix9Qyz5Kxi+a/jMoIdCd/xXxkTQ8ZeNtFr7s6HyHUSM7UVXGETU1M+d
M6/28/25QQ04bhRfuapMRnNRva58J7cJNCorAAPrknsiRypp0olV6uSEWrT4umRarz/8BXQeFrJl
5VOAGoEThVjJY/xtq22ns6PE21mWBVjl2nEB48o+MzcleVX4TpdMd0XS0N0GxlZoYcgkBmf1tuG9
cX0zLFjPYdsBJw9qt3t3R0blWdoOMscS3CnekB2yhgb0Ky2r+mPo0D/Fvl8FwWQIrEvMlGw6hooc
mJtwRqERfR2SIVV4EdzJ7cReSroX5OP+djiri3K+wrt22qpdV1jjTdCkGbJGSlH82vZFQVzsRcJK
/zIzVMBNhskJ+IKiWBTnMLntfnYfTvO7g0A9j1wXk3eVFvhcBFpP46oU5evCZdB1nH84qvL1Vxn4
/es5j5TK9IUfmiBhXmSdovC8NA4IMZ2VK3/oP1wvbraqazui+hxgjOU2rpcZ9TjTfH3fGlDSy8ZJ
QzQydKoZnSejIAQdJ85R2R3G51dVb87fxGhP6Xh26I3kOv0S6l7Xj5K+THgMBASQZ4cHp5wIoo2+
eps/i9e1Zlf50eIc1GrwHv/yx9EPuy52SiXlPft/zd6tItzkZJ6D2iUqda4FxaGkIC0JOvcNU5UH
hx9XYhWmijQHAh8Phr/mJKiiU4wgmLNnGXwIN/4xHEMQqisHIjdPbII7AJfGwPVPv1gMWziKFNzw
v3ih9yV8FKQ2LSyBPDLgBhWlKM9uGeZuk+ywx7qVmlJeGl980g/WaW4PJkE3ivItl7U6/iD6tT46
RtMZ2fFATeAcMf5KB6S0GyHEN2gf3yLHR3JvhO4DKLoNUtHK/2siWYjkSjCxkWdl+sjPtrzX3Q3F
Uifnf+OoPDN+Nad/rKSdelkyl8JyZKdlU+Zmak4aXvN1m8EN1ocdV0FLjdbH1UPuKUHshEpL244q
KRtWEvqmSYaN7+kfw8VFQ/QXrWHyn4pDeaVL7O8mQkf3tzXypT7Gj7ss1DjpVW67HtZcE9PzqpP/
NWk76Iv9DuH8qMH8buKZVWbzoIKqsIc/LqrJxQj7tX3n2L4=
`pragma protect end_protected
