// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kNniRXT59xJloPCHNUOm4T9DTn6NzGfOWMrY1knn/EAmaGpNTKxMjnb6RqZXw4u7
dhJfSeU5XBNEH2W5h6GCKJMu/ITQdnNkAz+vdpeNURq2d1nE3wTkpDSl0sKv+YgN
x7cUlo3M00KO1GXOzvvAb9OQ/Y/1n79Hc8z1nzr4qYI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12064)
b2bojIC7z7IXn8RFZQVYYRmU79/kpWSAW72lxQ5T3qtWSbGSFHIutc/hC312IY2u
SycgOMNHbMUV+Tq8wA+uzzNNwMEyIe0NP+CTTgSoxO403VPOFcLye5CZSrbg242w
FH7wCOHTywlk8XvrfQv15H/g/eB10+wzYT22B+19QLf3OFPSGxHc0+zp+kC8jxlu
z156cXJyIG2gtD1E1sHaK1nnzFOOCl1ZpO67kGJNhwG1n/FfA82/M3FCXGq3fUB5
RD8xpReUgnkVFrs9zgk+ELG5gCDjCxqn2cYUoHcfkcFDdPM16ueR7jGOVambj4s0
EyGMOjBoiUVw5bFgEwliGIww5jve/iUg+DWaVOCd6G9i7BWqTjvBmyiDq76+jBo3
8LOyydKp646OPps6BgO6x2+NTwnKcGnrrUJ9/89+a94b163E0c5cU04JUHrDwPBJ
XcZWnl7Z2Txbdxcx1uJnGNeA4keEjPBGi61sF3NLkPlAtA86+5bQcaeUTG3OCxdU
v1t7N3sOjSJeIbCfRmjQ1RphK4F/Z/HRD4g6ZcoYX2tga3N/w13jn65jkuUnGwhc
+S9vWRvGdojftxepwRzuJcm3YBn2qWpiCj4PZbbXDR2P7tM7rhB7FbFrrPlyeoSF
Nur5mP2E2Ixy8cmGniEZHvh0tpqUQJpxRxR2QTM8BaCZUHug+nG0f/n0cxl6QttT
BVxklxES9OcoopaVWzxJ387qAvJ4Mp3+DG2fSeTJUIS72t8W/IoAL1HyCZxmia9o
Lmzq7+YXly3maLaguCIhyTP6xetXc6aPlboO8d6ZIf5hPqsMc+/sktKftCjptBxf
MbTnmROgY1mXuL1WxtHg1BZDe9ZVKGxEbEnqdSnD9O608H6hzKQa54Y20EAvF6Lv
ZamIoCbz+c/W5D7bzCdsnqCeiljXLqOQvc4J/Fx2vTOppn9k8c+HkrDBiVB9ebVl
E2+r48c7QZi/GbXLV+lK1zqgFxSZR5lwhJgKb05pTNrO3fGZ+RsV1TFElOcRDFXx
BvwA7Zr62FvyTub4/JG5HDiaP+lV6/XjiQ7Hq95ZBujwkYgv9y+sSWI8IL0CcR+Q
UrpTkVudADylYgvq3EGCXDfgfdFZRCIhmnqcUT/kmOutVnpTaXQkXaGsCTD4MCsg
ayU/EiSbm9kF3nObLzZh6ieVC9dIlhdwGnyH3Jv/aEmVklZZbDU1kiBbZnAOZJeY
JGffLFbHNN//YADwKe6HPQ+JjzPKP1k7A0GIc88Td+T3iA0DzjurDMvOCgwv6c3d
hLrAGRUKbf5gjcSYbHtY4EF8HEXS/hsIJYsR25jRvvguy9u5mTGhF31j7C9OzyUd
RU7WT1wfs52wf1EL9dX1Ouz0d2lY4C83CUSDne2Wd2RsbCc22Wuz7TBbBxubtSKJ
O6YSUKZhfVq8L2o9tuOXFZDvkCaaWR+MRv6FJtxj++cEnSX7UqKx2g+UsDBACXFc
24Cgaf7cbAqIR7KY7jT/cBqTBe0j8+c+0y56yRlkDG2zJhtYuSzJ4Elf8PoEgmIc
PHCLg4qqvChaxR3UYBYe+C3FF3X3wNDM22SiCyxctQDVaJxNKDLOINZk9CSf8Gnb
d4UHef2k78tFB6ZoWdcmWiGjZMN8nlylbRCSX1QHvDjnAcSBFe8mjGeXdVAH24sL
7GnDdnqqVrf3Fi2NvaEvMSsugYF7phY6mGArM0q7L+4MVvw+RK2gbLKKfNfN6WNt
dFNYh0pXyD4FJ5dZAa9hMgVMdoO7nhiubZuXa1NDWv2dQF5VMHEfJ5bOb70jvhO/
tYJUrMo6wtdi4/rCe76u5mX+Mii+UskHweQOI7Gqu6LB88aLW9KWBCj4JtX9UnL8
tQcpQe7Ebk+qVfAM66jL2h6Fh5bpghAJ18d+D897nRwhveOwUB5DTCBS4wVp8El7
3Xjv/lyToU4b/jUHdf9tnA+r4d201Mqpy9IByEv8L70bT1sQY4DYrg4O+mLvgNYQ
dm/wAtsuJ3N1LCt8Wb2x9a9wjdRcvchD318Qe8u2Dy/O7xhvlH04i26ZHMKJ0Lyy
JOx+SnEiG4CFt5jyTOEynveJ7sEMWUUVXW//rKfR/JktbQnLrHYT4pWR5QCfbQ09
6sAKgwFXVcMnRGZw8eC9+Qp85ICz9MU9epoVFD5AkmE1OknxvYNCGr779RgvVGjl
FZHuEMniL00fE4ITavviX9JkIY08rnpFzCkz2P2E4XMvoyLEwDl58tcV0G/LiyCb
pcsXWXPr6UA8jkljBEr0lu3mXvY+D1aLOI2b9gfSMuKdLgj33IQpeaJzSLIGBjwO
QDMJFs8qdbQ1NZDSVicjdhxt7s2Dty81d+qdR98e95T/vvYc9My2NdG0iRZGhw5I
pfWptG5nVp8KK4AhP1B+T9wiVw7UPaXfvIR+O5gxk3scpvuex05CRsrdPrZSIDaH
OpS+mmUBZRd8cLACnR7NCXI1ljgYcrOReYe5uRxZolD3Fnb4FjKDM0Cu1l/6YZhv
8VvlAPDUP71UTqsE3CAHz+IJFbZwOByYm9NCCFS3MlCh884exQn0cJPzd3rL1Aj7
IgapcTBM00J3lGg5g5PenAXw7hyJBM5JPHKVMSqxNo9zLndzSk8tgESep4/D6cBW
rKhWV1Fnhj11iwi1M0/lsEGPzpgAqtKUM1hhxyxnCJi1E/8tXD1v20B3ud0maWSP
KISGfegv/yoPO3IpqSfUz/ix3HmUTrzGf9D2FNVdHfTIXBueIjHs+mpkoz/q0p5k
FaeGgswkprI6CMq/PYsTMUvVIz9J1MyJsJ0zP60pFNGAuSk0+v4ee0KSM6/5EgQ4
HNNpJq5vciyTM59Tob+oY7D3Wi5rOFwF2ov39oYBkvoZOesy28RnEn5wHBlWB1Fa
emAY51RFVp2tI8+9+ZPuguy2YZzCi/ygEhUDghbpNShyQOyDRVOOgcQzmFoEPfBZ
SKukU0QHUf8Q0g5UsiCI4ZbXKeyovATH3hZEofgQgKpy9JogRjzULxts19lkjz84
a2a58keVFRUAP5JYeKRw2lT/St5LzrWBwt97v1UbsL1Kv8TyA1OO6+/lEEFClx65
BVPwt8zB7UPJJvCpViehCfeGB03NCKhtVQiHlDBLHm5dTB/LNq7EX6NteL8kHPhO
3jAGHIaIZsGBak5yyon244OUZxsmH4KQgIyr9IPlRuwkQeeSDYFg2uAmg+G11IZE
NyiGQI2KfiroxrlQw5iZpxJvBv9dOfQJaWhqaczGS3xe1vVGCrYEPOA1vdD49LOM
Akr1GSFrmOnzv0yVu/gLOU6yohQVqts2qWbKD+5N63waI+PueS/8Ux3S0uv23fjj
nZjhQuD6Oh64sa6FQVFBNVy5QpEjZGww4jPhCjMy/GXfwfhwLKMSonk4UDcMzjZp
A+bKKyEwu+vWIQYimfrzyTTn21cHbwu8OxNKAvczMrsP8NYRXqA4ZA1c+VWtUjwE
wDt33jd2e2/rtJjrnvPNXEXgm9lFMkVl4e2oOJ8ceWjsZvIqIP+z9VPil6s/EiZw
GlyvqieQ7vgAGqBeihT90Ec1f1MFsJXp0bN9TL8xzcLq7GfE3zjA02zyWdyMy6mW
SKoOqn3rf1FTN6vT6xxqvXjkPNpFyqVfvdOI1pdleWzfux1pN00sDtfvHjFRz+mO
u2X97vEM3M1hSvoaVMwKV8x61HdcrIOC1FrGGCNIll4alLdim6hlMZP4d9dqpwJq
bFtvE2iqCABDpb79xg98lDaMXo0ZFlQ+QiDILHbd9rVpNRIsL42m+y4R5xFrhTIx
GEWxWDVmnsY9EB5qQyeq6jnlz2SZR1v+naZg328gXRxWfJYeQXqtj0FOpG/3XwDQ
TdyUv5vvYmSB5k5ue/KVFUayX+rB6QEXgLTxe0jyzrOlbedHmga2uzXL2BCYQ76b
mYR20FabE7FsBzrAesN7x2pPLI21DRSZZpiyCmeAbT/ZnrSNZEDN1aRBkWsofKRy
FKJ16UnwwrGL0lgP+1amSuFHE+hKkGxN7kdN194xpUqKeeIf8wwelbymhLwyDyZt
mAKHQNCe1SYmUOOfyTeD+13fL03bqSqGo66gdPAHl/9Lhq7gI46f8P+utJ1OJ1px
LmOgZIcYQ8JqCzWuk7PHt9NB4TPZzLh8GC3NGto95Wal4QaKRHaIMqYqtJCN5AAf
hKIRIGPq+mfAJnAmDtwxpUMQNix7pHPNkN6GuKaEsxjAyBm1C8gwVuWkL7Hgqhov
Bj/wcluigyMo+0d2JJujPGBI0cX1qe6fTLo7bEVLmibq7RmrjJPl/KEQY97IZujf
2t6VgdrVgQpXH0B1W1JwbTGtuWFA4PaGadOBVKw7Ltd+Wm4R2OmsG9o/27ggYIYi
VI0KmYg3uQYu7gYsFoG4kwyKhkYpeMwTHOPE32pTbLtRCrevFjRIsoC+Ew0Kge7C
iQHUx6Yw9U8CtySPbPTWc3/1vrwMBFRVkwiUfCqzURC3Y1UxmRAZWvD52nuGr0GB
LwcVcarkpCoKnun/2SplGlPQmOCSRLZBVhFDqI1g+1fDXwU034ZRElB0Kux2occz
wsGNxL033/O3gEEbr6t2F/SCwyCri030Xgp1GxFMfVkBW8hfpMg1rpZ0u27ifAbK
rTORoxWnDVF/Xa/ssZA1sDp/VNGukmOdqZPA/ahDw7Vao+QdgAx0456xkizQqSLo
frjjE7ae+TEX62iwyON6lv6ziInUGJOxBTxXYdSajr7qpIe3yMtEy3Dss30lDpZC
BcD2RM171l7HR5fMaM8CVsolNIohQKUhAZglFbyN1yoKUnG+ImBhjNyzDwbUG91l
2zxCtkBIcHlDQBZEU6mzIVy/5QD9Id/2O+n5FrQDzIfeWQkxvUQG7ypYVabmlgWU
oTLGP/Ii7Gns4MwCR+4sHm6WJ20NGneAMZ11WGFLv9ZphrneyzhfdKJgswo8Fbyw
zTQhExF21RzWEL2vzn4yJojS/1hfZUOp9OuJK60u/v1Znlab7kr3mK334koe3hs3
3fZpIvzuEAeBNHHVCaxNUbcGx5yzp0VQx1aNe8QpQ9/ma2WExdsyie+7mCv+IWUP
68o9gWhoS7k6tGCUK0aLVG7PRfTYKN/F6Tg/Qw/GU1xstYgluEBttPU3B9V/Yq3s
bG+i1J6DjR0D+PtRgn+xA1HitTTZE9d0NZO+gJIBorMd3QNKGV/nu1HytCs1XsRU
E4+4Z2rmeb9aJBWSUHY+VMAVbjaaTxb7ePqyw7+kYtQYUX2nPrWo2sPHGZ6fiqKu
kSDM1QEaUdzWcvXwpsWNq+EDZv+LnT88Zkd3KkupEPQps+Bl5dp1zpsQ0ByPL3Vd
d4mPmmyaQg0Uue4TE6Vn0/bdvhzqmEiXE5ewSvOWWweaFHzsFh/W7EkqK8nF4HN+
VXYLx3XhJYKGBXrRpeJn/aHEVrKBYNBfRVSQDNF2c7YHeoZN+Z5tuvx9+v8juMHU
Dq0fcwDVoWsSiAxg98rVlrMOvjRkpFGWHazzPPi/I1BVJ50srTmHviuILl4yttQm
66QFViTNeiihXVfZ9PoScajHsMFsQJnOlUkAUwTLaTVZPpg6Vkt76Jlg2S405woE
sDtzhKv4EjMwbDiquMVO4VPox2dktFYAdYqmpKmjYfjeLK/LGH0SVLskP2Vs0di4
XRGhU8xBzorRAQDj9nlBL5tWlX0bbhJFwdNIY4tiueiU1osYQsDMOXtNRVWIEK8R
G/wjBEgq2HtiEgDXi6Q4TU8drGkETAx9VqYMUhwboDZcsD+SYVMwQjdWOO5//PHe
lmP30lNNGaZvYTN316JXN0ud5M0WJK9m/TQRLO2gPjQk9pMdEt6gBMX6fXF+K2V+
RjVPZ3EWDusOJU96VTbrOLo4HY31GgxSm/eOTMqp9gpxJiOC5Ibj3boPUAGCH+pk
7SvNtZYlcf57bYpYm5GfKD+n0bTP6e1RyVLG8IkBllKiiLG2mloHMNpPfszWc1Jl
ZXtc2B7CkW4/PdXQt8QcI1ecvFdnAGbNsi32E4mV+qX+k54I+KLzjj/g9NAPiqsW
3hmH//GNy0OLVmn4u/3kagUG0FGA5TOr04s09ct0e7it5QfrDQOx5hbDS4yCZaUr
9Ye2sYxzGZg4YNwCRdglEFn1JJvP/AM0SozLh0xIRIlKZECyqhF2r5nG+NwcvNDA
AUNtpKtAmT2p4xSXYopeyU1msJVfYUhhY3hGPNzstG3DmQZJt8L5i/9teluThXcX
sAjMyvfxrxBLTw/LJAy9R3Q9uwCNjnOn1+uOvia4Mngi+eWHDqUGhOil8kGFwHzF
Dfu6UtinCPUBGkbuGgd1XI1RU6CH7cqF8fmIquXpbKeHeVD+IMNVmTV2Utj7JDFZ
SUffnZWE2dNrS6AKQ+8ct0zl/eGBHEwVo3EBSY4EDwgdq7eNY+G34e0o0gwE5b3o
7KbfJzcYEV2CO/k3b8V6pK8jgivLvH5jMR6P1Hl66UzxPB+IGDpQBPTiz57LREfF
afY3TDHWMktjXu4mDXJviCxZGeKWsES0dFgEvOd06zQ8ijg0l8zxM6TFpRyR1pbZ
PjjaMMh+8q4kV0sOiEJzhRqTMqws0jgcPtuJTRxIKtKrd1J8j2/91zI0J10OkRaB
u2C2HBE2+9a8eNRHRo+EQo10dH+r8LnsaqnOeB18MYg5yPrkVxBt3YUjOM8WszB7
KSJom80JMZZYDvDzqhBZDyxpPbfIrcWAQv9wZ2Wk/4pOvDuGG7/G2pgq2G2W2Xjq
/oBsJIcxHnuNCXZ8fZ2kSKxw82nQ5qb5Tj2K/UpXG4P3zwH28UXmt2TZs3Lyyl6y
/O9ccRo7WIMjI2fodtKlb2iryogFRJjp+K1/Vri+3rW3zku/rcYl7iAexUylm5hf
noVh8Lam2vPzNtQrAXIW8ctFXqYMHVKufWiXEtWxqwju5DsNK8Iom8g23zThKShZ
08WzIESihXhrWJ2ziTWpu7J6QRUxlWvSkVVUao/Wri/+24KCT3kk6qBGo9OuvNQV
G7Z4NyUidjJZk0akAH2AmUf43sFxTl0xLOysNLo42+q+gKV9XrVjMKA+voYNEqrj
wFbYD/fzDkxlgoLQ5KOSzq6Oooa9SXyXz0Z2dKXXjMUtrOHWFgq6YJCfJ4R8BLNQ
KQIXIKAHV1QXmIBueXOAx69yNpukuPhJUgaQG0QxN+jDeDMM36yLe/OoNI+HaRmq
EJg/VWbFA71aRj1aC5Qx+6iAE0dtsPenZiUm4/qSBScB6qE9b6x4sJhYIAS46mcm
h/ajsiKz1LnUWWsbFDB130FZBzHWPBgD1v6Z2hCuRqev5aXNvyU6sxC7Qt7Ul2t2
8QVJPJsBQ+bIIZjEIqF1nRyiJt7EU1mx3vZPAv+9+uO/EP7dehyhoqqwcPqfu8a5
Zfm6GzNjhWDjoDXP2r/aJ7L7cwr/lyBFBPRoDR/Fw7BqIecwFEYCnQ2pGVvQ0i2L
jr40HLvOSE0kPQlsO51OgNtC22vZ6/WI0sMtv3yU2I8eILs6LqZSc1Euv4mQxTS4
LTLToZR7bTuUudvqt7+DhxyAOckCmrrdDUbJqgAwg8QnRoDMKETY8Mr9hV1sVbcE
4lXI0Cs9XNHYOlfPqDlckODZP6OIkFoeXbsf/0q+65ibG1t/sMZZcVMoL40RMai5
Oe3ntxlziqJKJ5oQhYT3F8CTAVQIIFPx9/dI2laU2DNaHRYlF1QjeTJP3hVk0Ba/
2HOTXDrEmQf4Qj6fURPANM0b+kE+HfT9Irs3G/1XZuP4Pgbo3SGnEz/Sr324yAZf
0esy2aUr2NF5u1+2h1hvohZFnIeTlLV17nfIwF9q279owSQXN5lejjZQ3OA58Xyu
syjMBDnU5q2J1SwLnfUVJ+7ZN6owbgKgAaJRQL/Ovo9IKGR9sLfM5DfnVT+dxwWg
jI2bS2Rq8hoHvkFiEH69pdZGqrsTx6XzdniXf5mEdXsLc9+D93PVU2Hl6AX9Jhzt
5sax70CwVOzzWQoLnS4dqaCPTvVwZk9y5MflZUwaKGffMc+a6N+KgFQjUeEwBF7n
Wp7610kloBahhrYywSaNU0XNo/fcPMty1+ZbK03CgQvEob05YLlciKMqXdzIAgSF
KsJXMag9GhNxo1IXVJ+gKuIFosQeyPEEVHmtx3XleFh8/oEPKnXGSfcFAwqVeGtr
xuzXNh/l2gBthkeiwqwT190EekjYQed8Nq61lIQXqyRjqd+RgUlWT/Vn7rFSLIba
WzIamJKIm0XMblqHv+G7PNYDpWQMyx3/zrxSLBU2NkWIZqJN7po0PaZfwMEhqJRJ
dtl7WAaF+PnpJsGBaMBMv8b7FC9BStcSHLLIwVLU9bkH+PBCw2VuU9oZMNIIy2yF
U9Qoo3y+4N0GuLHIsW09dpMAdWH8RuqI033N0J5hDXApE1m7NXs8TgEtYqeCtrKc
scgVUIwwVzOWHFaE/ZHMqgQtNGJbYehCu1JU70HeDUwDaSh9wa3lNC5kDvuytiXb
Fj+lqKcmYa3NFRIQwmxtx1fjV3knkNXMDFn9PDt7RvZza5bMwPJhlq7l85+yCIhz
qN6yQ0QXRz8MWlaV6QG699wzQupg7BuBLMzrTjSjml3kYBv8xrgcKSGAJ28AVMNA
bhn6bJwHJvk62CcoGFb6xOiW7ABzGxZfmxDY2aoLQ3+N49TGMz11cB6XNpiCQrl/
cHpirGk+8gvMGAASQ6aCuZgTnuSaQTBIpnY4TSlBv/q4jf7iNknB6zT9u8jflqMv
yHJm2QUcHyuBlJ4eufZyOh81aOOorxyvo5Vw6CBuzt/cuRfZ7R0U1mR0inMqc4Ug
pmKFezc/zABOyGPCsOuKsMr9Njs4mPUVkYwUj9qCzN3D3s0ehW4KgEm8JaG2RzNH
IsCshFsz6cOZg+OUV3GskOKQmyCq4Yqq7dDVxpV5zSas8mf4r3T0MIAA8hUFICXD
EAadPq2se1eYnC+it+LEpb6t0hOCGOiHRYFVMbFsHnIzSRxiM+ergUb62dlvA2LP
h/xf0S2cQd61iss2j0bzydfOQasAOWUC6OK5UqQro4Ukyd6J3ySW4TLlP6fOefkf
/iUVnogpbshyDxLRKAK7iD1NZ5BuPmbDpFjfu/eEUMtP47QoVpjsNzFKNlzbNaNn
yuSSDmQQCesfvHmo1HP6E3VIBD4DF6uogaEAwG6tNJ2uSqmvobt58Lcah2sb+akG
wNkDEETe9gEOSRXGTom/Y5PtO/JNG3Iz2j/Cn2f/mLO4zxbgO297Iz60Ll+P0AjN
gZe5cTcM3cBSfJE/ZL0lmug4gYf0uKNE7/XP+QncRkX/EJuf7S6W5F21L5Qh8rrq
Wnh+S9rUMUXH1GqqYw0dl/ZdqiegbMVfJCuqxmzoUPKA02r2ntmVc1W4wHbXdXKJ
iJIvCxlgWu85kNqAHJroSu3xNkXVxq+mKKWYqk+KxxsUBxJ5rOIHNQIdurNmmGgg
W76PFqxF8r5LmSlEEJPxUgWfxxysTd/98b8+Wiv6d2IyNd5t4wTW3hOEDCOdEfv8
zLD3YX0VXfa67uNQ2+QH/DumkOOlszY9mClR/wcYoBtcU2ry7aVKYqGt/OEeEu2m
xTYvNdQkpu7wvfkbfqWKCDrsq/59jaA3l4Y4wQnGRrYIEKgvXGxfL6yazkXr9DGK
paznCnyqo5zQsardhFO2Wb4MXpqDdrJHoeMO5sHP4GDwVSPx8Bd5R6yAt2G+dk8z
gaXlcNzgN1gh/FiXhaCxPkda69nO5i60tgoe/9XPX7KSnbEWFhgKrSz3Njwr6HrU
RZEOKlqWg76GHWjJsICLLsjOPk6DpvvnrW+x5hMtvq3KfD2hnDrEXqRbpd+wCARk
pHdsu3iAbEcI+exfTuRBSXbrI8AShNpv5L+GYhc1CtjCD4niljUnE0qeSomEo56F
W0vP5e0lfKukELUSFdXhgNlDsOEvqb5oXqZ9UTee9+jEmXZC761u2J6Q+EJZqSsN
5NEXJsL4DIbOqHSZdBmmOZ92jouoctDib8Sn29qwduIRFIEwMNCGBhRYJk3Xbzss
uIQkJpCmYzQgufCF/9ITsPGuaY9coWlB/dRFKdaCSP+t9AcUX7O28yH+PvL16Jpt
QNd7IjUSdstDlSljiKx0Jd2v/V2JCv1MSYjXsAK8izJ+7mLQJDfpApB5ZMWT/iAk
XnuB+40U/bY7k9qdD70VXsWgIzTpAiwI2FXKLioAv17g5RGXyv/XrVk9I40O2N+0
vj7oH0p1K8rl2eLRi9GGaRW0JrDI5lsUL8EU+sZjxaGfRyweLDuMzwpSg78ATB2Z
ns5N8CB8F+EQZgkXwbiQfi2NKiXFAzg5Z0mJTiSgCSHWWdEWyMMt/92TemNfVYip
RLdDnNtKvn/VS1DGW5VzUqDRVQpMwdsZszwms8ZmYOkHJZmyBCT1LO9ZbMxpKnvn
LhTsgCWvOsJYxc9pHALuUYotoQLsY3GoHQ/unLBKn8fzugT7p9N/1yoqQANrcWbQ
fU6gKB0Go1k0zJz06Q/XdB0GvYrpel6V4kf0rUEn1Z2G7IXB4XoRoOvlN6q+A9iH
kKi1ioYA+GU+pS9hF3XaoLPaj4ZAmynjtmpjDvn1V6IIRPXgQaxLKQwmqLvhSnok
SiMF4QRZaW9AmBS2qmpJxlzeKL1GccTBoPI2kd+eBYOhkxqvMt3CwvbWKeS0LkgX
TO37obJs48+i0m/AcppCcLJLLuEJE8Y1j9OHSbFNwO7U8qv3fXyk+cVSRo7M78h+
leXGxpl75fhf2cCCI8xFrc+683FjAaY6Sf5kdoXgXRa7TPg3+GpaEAfWMQhw4qbM
z3l9SDJK+OFDsCyC/t3qLDCZZw9WT62S5CQ4wls+ebqvH4BwpfqjZk2WMAnOjghe
HTvx/ougbotM1wKysHZWrM0i/RkLdXr6e1DBki8VYlu+i6ckuvQtls9T0R3ORxRn
9qwkUxoJNU1ZiuOsB1Vj+pL2/5CZ3XTVcf5yvJ5jVl+d/tUfzggJOKwdZ+ujYLPQ
+4Obn+O0fTFbmUCSdBzT2f9FOzp9H2mymXoebdu+mRuL1u3EV05m3LaOorz3jLww
oeXYPZ5AuVPcAAykUb5/Es62CFUNrQln63eqZjG4U8SoTqXwqjlIJmld0lvgtC0X
ftciaLGaEp8ChjtEfGBADrXBHr4aLz9YkEmb7MnSQLOwBbcYiUSvWzq1rxg0oZZP
7Q3if2t9naUo59zgz8nA9QqRwMVr1pf5VEAs9w0tsRHUB5BVXurl2SdKoh7TeRgz
JX6LEGkRyrPxZmfO9KH80t0uN19CMtMFl2rbuvr9DKzDT1ltXpZv9U83ilWIjZl/
VFe9XeqTYIY2b1IGzbOJBInDEqPx9LaooKneXdCfrS5x5vE7UCCwPFHN5lo8ipo8
3KiYwMATMuP0yCkjsM1IdO10WDPJgAuV8jL2FlxUKzZtCxe+7aLqemRy6FULRUPb
APgKvrHzC8Wal+8C9kfh4LkT3HIQ2uyE/45KDWYU396QFZCuMTZt2g0raBCwYuVq
Ryx4JAlBadAxtmSwsCyyovPV2yLbiC3OuGj2JKuBNYVUFY0+C4NQ0/co175jK42o
l/IVZM/sqlwX3kOCZDuWqVIwnmz2I0UzMfHUNaHNDSywjXXraHhyeLect+UIrb25
lBfV0MFf1P4m8EizaEfR60HaQCffkoGzA81GxHZaTN3VGDNanjLWmNCUqpoCaD1F
W6LuLZmid/V5jwGmTQbpvjc674QsWTHEAhrAP2xMTaUQLn/d5HxQQ5LMe9modAhc
L8jKqaLWQbdOxnETm2GPdYyfwAGFQcw1F5pWF3bf/mfqQgIQ88IOHSCmSSi2LJ9U
kD9FkQqOCzpbPCVmzbhSgO1aysB6n8VbMWepjXV2eO4HLkfJmcAhLCm+niMpPdp5
zTQjqZMk7+BrJssUHENS02Uz6GQKpnp0RwhF8Irh0FKQHDxNltAAvSzwp8nXxNLW
f5JZjjJVQIrhHlZlWWYCI2Gt0gOpaoN909uwBysFytZ47vdVK3eYNbKTI2GWDQTa
VeKq0F9nLJPy7ZDZR6wazs9C6UJVE5e3Dl8nx9KubFbyd2+DbyZ1B5M8mEstvNzn
phtKoW7IefVGjTH+FGZWxPsaWNlJJj3EYa0tn+lPUHwjl1ssSRphxqhsDZuYhTfv
zCQyRTC5ZQ4S/xqaZynQY6GPER5JS2VcUf+Gy1AV+C5uoZp4J5kuZH6otbFCp7dz
YiwN3VwHwO1Z89dwMYr7ZZcj9ff0mvKt93KfFeZUxwi5vEZpFrDIlDz0M6u6KSL2
pO29UxGUxC0yPLKX3Iz/i035feGh25CFFXfYgIgnc1RCgo5IY6qaitLpLZSzEHsA
porNphYwfMUIQK+VuhV60bEl/6HU9RViRNFdC64owPf+9PRQLQZfw84tZdL/NGmY
mZAn51bftVj9qmt2ivvksEohbE5Ubme88dsfkF8lbhSWOUd6Pl1UnCnbiWMxPIvP
F6JFFbGeHnQIpFy6zfsMAM7VcaeT5BtQIjy2o9WlXSHvY0Ts2M71zqL95B1XXgQ+
L+T2mCrMGDKKZy55U5v3MyGcj0RxOjUeeQAuxb1ddQUbM5IKzlcQ2rptOsz0bTsZ
AuxS/PWfvEHzHf6LsJx0SvWiOGvBo20fWsiYBNdiNpWfBYCdBEGuyPaSA92x3qq8
w268Am1S0YmtETefiKWb5x8P9EM+1S9wMhHXkt0+QW1TLBvOfQ6HtGWpBkFybiZm
TyEV/vNFAiQ8CnSweJiE5jeOVWmY6RZL2b6Vi0qXy90ui6FxNsEUIXHRgaBd7DDT
B0LTSRRskVk6ycmB5XUmXvgJ+8Wh/sgj8se9V1u9hCjIiCDU3LculmLW7rmHCFKJ
9PiwipYkHZaJBiWByCr2LF6ucVSV+08Wiyuaqr9x19L/Cl61vghD9KVDCTFgq0X7
d3KdWAZPRBY3IaVCOGnoFs1Bo+G3GJEtVcxmmwNVlIhRE7NdCmNstSPhz50Oe09j
ae8iUzMWegi/RQ/ShyVziVzbKBL2vD6BquaNU9BSdfNTm8wh0nSoK906QAYqvwQd
iPnlcHd6G7ENmr149TRwR9Fq+8WcmdZ82v8xU1RyNq//PBwHNbfTQsfztpYqfAUQ
9fsnBjkd7AyjdlrU76yeq4fYMUIU+hBNya/7qtcImG6PjOBTmvs3uSN5jG1goloF
nLDMfttrxwQ0clITu2QuFYOjnsZqlg9huYC3Nw9Ns34GvSyZQVNv9w5B1YOh0x/D
HohXs6k6HPhftzBRb9kSRKlDj1m7ePWiyMkDcqUw44G73pbLLgVakpF/kvejRJ2U
DCO+UQk52JfM4rVDe3lwn9Q6ZcV5gfm1NQlJjChHITOH2ywmy32zQDwz1GZGt57R
8b1Mmg1pzGJrVRrjxj6YKheDcHP8DDrQ/+2XAzENH3KWCCuSVgP5iyRzU3iXM7SR
icXxtR42QJCBuhHZazkyJTdgqLJWr8zaPkKQN1iqDlhHsww2ARZPUfJJl2IOJdN/
tbbrlNiGetVibCOfARY502WJ6YVZUTKeTh+U+fyvwrI8feuQcAR1eeEjveoKEKqw
BZqW1/3yZht9ClN0yR8pf00oPnul2QV/txyreGqVwPJVR3mvbLcv5MGK+ZX4Lwfe
lXy5wt//89lvZI0Mr3diG6fG2QxM4vvglbbsUYBMKtfdE3yw8HUQ302epcbX9cWU
GZhM9mJUGSePd/cowTrZf1P7QUzTNZf+kCdNJwd452hRuw6tkJtOJEZPz+yRnW1L
lTBL4mKFa0NX/0Ubp5dWp+a7rd2QqtIm+a0+Q99T/RQwEOiaI5Qj+Gb6keDu1d4r
ncMxLQ7GSBrsgbnlY+2Q2M1MazoHXnroqgu5mvLK0BzY38+U9ikZtOiFSBAzmJII
vZkeSRnjjkz+/xfm7clX1W44V/RSlkgxLhFy2QFgHE1YzLd4+L6CQjatPEsFPfwr
giWLAlxWXUhedDhhXi1dZP2RTAMjU8cZTqpdYIBEu6AS9WpC6dCp8s/M/Qj6GYDV
leMKL04HsGhPAhtM4o6OoUo13qFL5UxiR/kTLodpE9SHLGwKlwRLYsZIr8HtIUuN
aOKYo2DMvjIJc452MnHmhi5mav6G28UbVw+Wj2kByilkl+KB891LsrjwlmtGMIyQ
qyJ3v4pEUlMBKbxToEzxgEnGSPCukYQiet6h4g9xNgFxbancZ+CG8ggnO+tXOWoM
YmV2wTK0g92U5mFrPZ3fB0PDxUmqIlFQyrYXdIFmw5z+evMDIFBXZ77S2vdAqKiZ
ntREkPALjT2ifDxkW2ykIGuEfNEPtv68JvHO2kpacLDVKHRstg9ekCDEpgz34NMw
amHWAsedjbOobRAwHFmxYzB+5unbNYABu2Evvd8MIJU9l90X1ScTG5Wa4octvXp4
3myIlTGe1ClAZi1diObP20zco3Q8VkVqb/UykaP2/cy9f6neniOgKStDYi1WVCfl
JxxPPILYhzYa7DESyo85EAeFPeNpuBukRLPXWTd7WQfj2jX+lcYjRJcF99c0XayU
O6DIGVGkqEWKlDCSYWwNWeY9kgbhOY7+6iHN6bX4nb6PHeFmdl8+auf/aKGjwMsj
GuGoSKQkWnmxwRDO7KTEKohN7s9RwmJXxvmi1cEghcHQQgX5Gmu7gSy8bdaJGNRY
csWhbhJHBvGBmUEQSb+8RiIiosX/xW5IAnh2Jryhz8qQaeWUJ48+2UJgvakeAvwc
HKeVuocUqTkN6nuIVRHbTttojLdh/HKmeDC1i0EFf+ouJoyHVl4nMkX81CXwdCz/
pgSfiT5U8s+fDX6ogYWqoaark3Bz0PJhaxjGEO/fSDHsyqVXgobY8SjGJAfFKVLO
tzHpVDxxpk2BZThgJvHLaFXpIk+c1p6k97eFhBP2STWwA5ptvCx9XL1SWnMPIERC
rW1BwX1+yoDLqXHVxQIbiYZf+HyhHvqV9jJ9HQtG6hOO7mCEKv6E0lUYB8Ye5C7Z
xQLj/l9+3yOwBre6DynyfCuTjZsmEKO4Xf+4trzZEcBEnsVdJCyATTUJ0mbiMkdg
LxAYOqe9clyHoo72hTV6HcTJdG2KHLxiJ4FOXiRtL4fcegAQaGGWhBjuRJIv1bEm
kPZYPvZuBee5XQdvBY/hy7UEoyW4aWc8LsrUZl+nPWC8SB6PwQIRRTDiJPYre575
dV7i0QGPIqRkvZwSQ6ctzJXadrcJdaq0RJwiY7w8BiaDEufamQCmyPeIWo+n7P9m
tlEI1BUKte7RFMgN0qzyNgvmXfayneEqjkT7JZP+IHL6lm/DW3/YAQep1r8wPpff
3fYWk6By7X2KQ/SFsUAV3zUkoKxg71jpukGiTAS5Gx+rXcyCtN3nqleH0YuQ6Gw6
XXyHpikAX/SyqXhB5CGTsr/vXLzmWC5G3W44cEzwihvtNigV5jYUWrR9pRMX7sVv
sWWFXpTffZs7YZ+BS4ZyYxAFLonCsiyTwVqMHJAQ5J1aXqMnZ/z5Gi0t7wAmhbxK
S0lz4jl9yCtC1aEiyqOYVQ4eV4bvfbTfp8H7aniHb9r3/KLzAgpqyHSvsoxFwNu/
uG3VJ8PhAzKPFqZ4HtIG3ELHg6yYGURbjMl5iLNwYpPJCmLPF8jSw+nirsdUaGpl
AVGEKjW+rQjbbU33Ud/jmAuQaoyteRo14Cnf0PueUVO/DdrGAtN7SYf/GiuIr5uF
g4sXEXbWQNH5RYv/JTb8S2kiaH2L3efOYxgxG5woLC/2DD/Pk+RqOIzqP6UvANAq
ZBAYV71LO8+zUTsthO85OML1g6xr1eSbEP/d2ZqjCB/To71Jew/mr8FsaQ5PvKgN
TVPZf0Id8MzyAWzh/cRZS7f2PeLJEagDcLkIckrCYR+8Bs88uyby5nFjlWwYZNJC
KxeBAN+T2K2R0iK+Bi/+DaIQei0dY2Ryp9Vo0Vz0KssFJwwv3GBWhQh4wzM63A9B
T2qtYxp2xiAOFMuTL/NfGazH7J3vJdomZlgDnoSv14cnYXSd6RdAzSjslfy/eSDF
OBUdGB/NGD5QKtTVCGfxnclJMe5wkt1/qPofdBJ+RcRn/RC88TiYahupTI/7ZJX4
Fsa/nX5jSHmU/z3Bxb1jl6QWOaL7GwA+3NIh2eOvmDMleMtna5ZH9uHeVfPoEnAm
WESA4zpZ98euuF+1zIgZlQ==
`pragma protect end_protected
