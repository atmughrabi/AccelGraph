// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iEgMOcPgJ4lOxIShwqRB9BOQfITjSMywP/6+dcsY+7lqCwztkma4JnjS+xj9/lYi
TEBmjVAwLQOAbMA9Q3zrIYoy66wPOerKHXB0zZNmV+NY6tdrM4pjHpeFdDG18REF
8j1+2wfLb5snuBxzKoaJsMMKnLDNlt5VtRAD6n3OoMg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2672)
A7MRYHxMa+CziQd4wwRgf986d1kKRq954I5s3THJysIrWrTtUAtGP0nPY/QEJcIk
sP3k8Yq8FGwRIYBN4/JlWNJcCW92lS21AV8pXF7sBn6bNMPeUBoae6MLouFmjF6/
TqEZzSEkq43cNGZv3/1OcarfKPq3KYZEys5tAjL4fj0c/1Tg6F7xVg50TxMmMBiC
Kw3on64PRYUOukc068pK/5a+OaTkckGIAbpyiJW29IWfG4iTU+kMWADYssnIPgkz
mru5mPMK35qVaYJ3VIYGT2Esm6AgSB2/oFPbyzu2esd75W7cFehfX+mwFkms5zc0
vZ/j+XAFcXlYRHw411j46AFSi0jgGaSEE63rJwIU2wVA9AETskFSvD9Ipq6rhz4J
rchffFbxw6czjg5SkJ2Z5fu2y7kzULpUWGwlBu4vnfZiPfY/gQk2h4SQQYgQXQQG
k6i4X1mEwvooyBPTDBjtZ7CMdbjYpeWTYIRsgfjUDfjVX1XLXE126asPH2YwziCW
87S6Vu3w4edzazTYH54yxF0EVTKoMI+c8UJzEHmDj7pe3eQgLq8g1n6p2RiJ1ivD
OWtNZ4dxl7R6LCShTfdL5HzrkVyXIs5u1/qcB1QA3Z0PBWP3vWkEcP6dPdGeMMkx
TrsOAwS8LDFGKch+5sCAobKsFvYIYuxLnW5+rQvw+tdQ3BigAwhlcA7st5yfu5Hz
N/yrRec5/BHcawRyLQkUCdCL0PV+MpgA001aE3ANcZbPZ08faBez6QSreJtgy0vO
clFOF+JwG8RF5vbR3SxeCw9zH8GLs9AiQtxeZAwn6KqHuhE4NwzYRQUSLmGcOYYV
fGWaMjR9RXu0lYANDkxkuHbGcbu1a6UkZ9tvQNVyhOsCpbvb43gwM5QBBzXfFiaL
1b2hQMELZiW/XEaOwk9wvOAwdDA2Hht7huH87Yg3IVJfcA4CVfdYGStIhbnlmEWR
fBjg8HSZ4Dt377g5xu32zNSBXkL0gjbpcDZN8fWVOj+OPwUwYWrG+YTSZ1tmLJQQ
JF9sIxwbp2XPwgPz2Fd0c2RlpmLOBXNhZAnke/oo4/k1uYWsAmcEjh6WNnFDiaaK
9lf4CmbHRK0l/aow/qCeoXQmYP1bNtG5thM4URaDnz2M+VEllLFuDgU4RzZ64gHI
qM+M25LNWunJAKjixGLOjKiiPMHPycH5tKJwSiomvRpYIfK9M7TmLbjYVBNGjViE
2OH4kTXiqJgzySj7irHKay2E7oF2FiIzuNkAk87r8G/dx1VzUprlasqMxmTnQllX
XMgZ95y4I4aZ2imCkmkyThamERFEsH/yvdR5o5qtzKHU0/MkHMvVGtpRKqE2RIvp
/ahrPf92RJiGOzJASoIzFE1H+Wr7DDmg2Olo6u6ZJhKImE1pxuMPU5LpVz3qJ5l1
vHpHh5FDzqmwd3k+Z24to0dnDb9jEa7O7AW6ChfjuNQeEooXvucbu9TaQcaKzckS
zOQCrqly4H0AlItmHx0bllVddHY9cmbHJT6Yaoi3s4XAr5yh4Le43AFWCdgRHCvS
TiIT1Jc4lU9/IjifAuOPcgoKEO6hSUEUi1wvNswlcbetWvkEXme+J6/PB2nMkEmd
SFlTu8ukZ7cmbKZhaQ98cNbz/qXiEsg178l9bKGrgRwmX8vmGh4OxlhdtxyRFEZR
leMi9RhVzBLkjjxg1IG5yQrl9yFu3Ubf/1gvVsFRZSuGNbUOa9DViawQTxqnaCum
trtohVs5jSbKvfSxu4w61+KH5xsvQGP5MBqJhRfwgFpGkQpSsTD7ML0gxSNKo+0J
ybL12ZikX9T+5AZrsn2itIG/JxdwQMgux/dBG1DyXyU+T8jXjKgYzNCTzXVUfQCj
C5/ekTRtHZ0rQJ8l0mVrg6mXjpO+E2WBLZutDj8W/XQIYlEZ3baUy7FH0n/WHv2w
oujQkCmNcOA9W97XfuT/zfyKSdRABX9NABjPxxSqOX+tORG109od0V02L9gmM7dD
pNTbGpQ4yb9IOTDB97DrRm3Q3uL7T7lWXtMdPVFxDMT2COzY6ARAIUZcpgImqcHS
l6xdVkjPdNcuakJDGeRAby5KBu1wGaxV5YTTTPxafT/hS5uGX6PCvHpw1aGsB9ru
V4xSjoLcj+0C5BHuqwdxUBUOOZRUruCyqguulukd6omFYLEr1M0k6aSi3x/GzFx4
oSgQEv6F2nelYlDXp7BWzosxi8xvxdnglh/hYv7f1FqJkncDjg2Jy9nMkAUkshiK
BFDt007JjPUXTp6cptFLyQOJBj+r4DLjVsdQChGwfzR5kdZqhq87oEab27EeFH9n
A9LHd3v77GqDyNsoZnsH8Bw2MpRiZSP6MRjXSHIJDQ9xcFK9JR+/yZmmh7qxkH5G
m3fTwPuVtruc3F9TZ95xxVu0R8Fn2CcnPppJfeIPKhmcW8muHuJ2tmLfLD6q9UPR
Q1ytZb8nfOpFO/9gwy52KtB2fdp487vhpNg+Iquk/cXXvGD1avn9AQWHYvwN17tT
NeuzVtEedTJh/PP4BoIuHsGKioeCaRUINW+2Ggw2uYFIizUmJKJ59fMAbP2a9ksZ
7NVZIeR1hAcvMDOgYG6W4JnGGuszkXBKo8dim9H7rbcSAIWPWCpdkUTug/98/G4N
JpuJk/iRVuZv/9N3T3rgeUeUfmr8Qq7cRwUr7AG71ihuCMdkIORUDunaruVvW3cZ
3QcBwKHaFdBywTz1+5O31KTolR80fRlFjDYyt9g9t+FSh/sAbcPhiy1dUXRod79x
LPmxfoffY6bt4wJDIWpEHuRmiTDtoP4Lme3HWZxdHcCA9kKnghDu5/TzpPFNUSBo
mQodJZJyp9vd0poYrWI3LVnBbaWjWYb4Yp3DFkxxXs6ic+AFzrXYWnmei3DL49Wj
NxRW0wPO5eKlfH/mXKc03ceaINyire1Cfr+5la9EGy8hKg5gHW2it+jikf4GeLhl
JBtzuV93cm47n1gEmDIvupAruoKaMVrgpgxxGz/hV/ZVZnmoTYMZk3Ein0IU8WDs
xlkE5HQoz2Bi3HvE0Sj/PR4EQF/ddcYebPYvYtXofHAZ0Vjg3BsAoJEvvG7VJflh
jJNK3gAfzR/QbYknjsqbnCy7KeTEFJGKQbrBiAv3wA0/WPiLB2UpM/At4nUxHkz4
GANg94hGTFpEG0uRf1NfnTpw02r0vg9tEj4vYFJpiTDde4knWM5j8TzJZk/gpOCY
uLJc8oBbey5uW9J72THHlbYikmGTvm1uj6R6DW9dk00qQEmFNOGnkocRqxJvNnk8
MCsRPp9YYJB0MKqq8g++nSBznlRJDOjXz0oBSIjlLjmTkEOI1wMzq6UTRE2p5ZaS
fcRI03/+m/UnEYvBS+trQT2+IlJCjrlpDVtypxLOix0I49oCLMYewc1gD98Rwkl6
dE1/gTE+UX103MFU4K+DFXSRWrxy+x/YlY5RW5SRijksEbBq88FbzoWWcqppyRFr
dMfGmcPEKtI4omIexcxHRXP98FxAvCQ4U/x2v8npiLdbVyzREogWakftPUxZgY2I
pzlwXdfVdW0/9PN/2HqMTEeeNHcc8tBcZRMkI7JdKTg=
`pragma protect end_protected
