// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GS5X5j6Kq/QnQc8/pBUpOp2ILCDPu8O5uTKaoY1ZBv8tORP0JuRc1LFditEOHKA1
x96AK0E4UEHHvXBZ264a+NWtSAu2yBTtE+4wO4myftRZil9WGFnEJNnuaVqPJqP9
1ppMtw/rjJ0VPqlew/jDyLtWLm5dmpiuquYmodPVecE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
5g0fz7Rl5EXxbxb7Z6jAMA67tL+Kg+7QpdBUXI9HNLDV4BNT7pYgY6Fex1QBiTZE
AKOLhXoVfZnENUsazJyrT/QolgdMAcWVqViI4nCkDKGiJ0j7Tz9g5Ld2KwYcxk2A
9aGs2rBR8Z+rElveuwdkkBjDZ7g6X0jIeYYCHKRfDDV0hPi3vSXz5Ho5stSWsooX
wpVQKI9g5DhCNFmrOGzL8F7EkouSxXtKqnds0llcO3PTK+y6mp6eVZhP+lU+mIFX
TqA1LNzDJ9+9L16GgKT3GGULYTf65L3/2Pp7ygjn5QSWzvy3rSkV5knoxc4W5y6i
2O5sCzTHLdcXylW1ZwErgEtdjmVcLDV+1QyUJ96YFO1K0mjJS3mXi6o8xX6+6VTW
WyPeynh/0YXyyf80hqmRmWm1d0RiyX5w1bPr+h+bNn52y1t/Tnl//i7CwzeDZAUd
IwgTz3ZlS7lqZW4RHRWR58GAQDR8hKYCZIgExiB+fI4lFQjKiHhsjQ+J9TPLuSr4
lf4I9GdT9ufcUe5HZzoBQEvVslLwqi0VY+vwRxqFfxFfJVoTZkAPCCCXnN2PUkV/
dGOxbZy+MSGqQhteiMN+YdEF8jp8ROHaaUdbmMHsuRQD68u+zmOMVEpPhw+m9lJd
KZkEh+aHrpW3n11ZKXW8o0CjGRG+N2bWGK0a4LHHuz2TH41w2Yfj8Kxos9ajTdYY
XkDUxrO7rCKv6gkCc3f9R2Mfr7BWSqzt9mr0oJVff8c0VLrMtpvRVV0xUnXBYAXu
HGsunlFK7+2DMReaSyl0h5mlNYClTDJPEe4lYow+yFDQFtIqg/dRwjjiowPAVQ3M
ZwFm3KVBl8znNkNFrgf6VVLd21/eashLAcwual/Jr8I/scH3cIUf+yCmiEE2iBKg
XfrGw3db2sfOvaNjTX7k0k8zXokj+3zVFOpziR2CNgOxYTPfIBUHfQFGpIZ6lu/T
pFpegFoQbmDBTUTvm++CDtnBHcUdCLvlZWk/w8s/5FCUhi/lRajjwp2qlP9DzutU
9G4RQABYj2e19T2JjfJeNFTXjczXpW8wSRQUkkzUHNqpu6QC/ZsyLuFLyKKzrYlA
HKYn/MGOmLSpP5rsmwrtNzRTU423nfqGjgsnI94R100Cb+mzANEFRXKWlUG3XXbg
G0bfBb9qOQQ2PXa4L8V5L1MibeZlut3ntsrvGQvAWBzi/UET7CDDvw3LyIusi7oA
6HT3zEe1zSfu4vYBgmUUBKwMXJ5ZZM+uLsIftyQ7mrg48dxfmbb/eTLk/8tFSLr9
am5ZTMhPA+y5bOhnYgROJEHMYUZidgytFhAvX9vd9LOM7OqFr1KXJKJgj+lAwt6Y
hJBdWGWUJ093V+kka8JGUQ6q41dNbZEuvi91ZroS/2ySD/d6T6raEz8ScFglhM4f
OXNUR/gE6AFSu+cWlUlwOzpi1Ge0VUf2736zDn7gkF8rRHxF6nnLDHEtOAJk4khm
PzTJFvCE32dYQ0K+Hrn9xIXuDmMsOiG6/bjm6JgnSbl8LRI7qBzxWwLJ0Yc06UDu
+lBUSS2aWgUL66Wz+nkno/vV0XM+1MxktyAXD8YqZ2m8Fuj5nmE6QaNXwau+SO84
vp+tArcPM3mFkk64H5e/A+vlEjcsDCfQ5mWxjB6K8F8l9CPNw34TNcS88y99GGRG
jdEj/aQ48z9O3LVJVupHFNkZXaOLaciLsq2umA8As8oZdOb32lKaroefBz7oCHWA
54Gg1Z0Q/qYEKS4PTlA9KANdYlEIe4MTuYejDEWOgxQfxsuK2G6/Zpsr8KK6VJmy
DCJgE20FNQGYEGwMRkt/e7SXf3ZoOf19D4c17tOG8NR+ckE8wrKbJJM7S2jA/mCR
p9CQPEdl+7nOk9W9MDi+lSPNlg+wlobNCxFk5q46hZuLcl2w9fd9PMYTal7kdKOx
49b+NIk+pY3ELUKEn7V+SZgtJUpoZRRVfQdCw0E36pJxAInDUVvP0qiDr8i6j1Lr
BYj2Emc21EwvwKudcyNdsfP10K7clLlS6fibP3mFQ0X92I6h7HJArxTiacLTf5xq
sJwOeOxzKVEabxNk1ZL65+HE0oNud1qzjCbexrTH/qSWn/QlWQQvIlZA5szwX4R8
QSx9KxBKfhbfK6DtJqslfRBfVgfyII/VnQdxu7y98oLmUtMWKS4EOwylDPeGWHg/
pVXnEQbT2Yn6rvUMFJ7mjiL9CTInFuVmhcUStdXJG86QqCY6I+sdMQWXzUYLBSDA
q6nMAeMTSGdwuAKAWTH23oKkKSdT7GzXNfKRMU7WHTA2B470zbJf2xSCsnQcL6N7
Y+SWCdxYlWRe/GiUZTWEHN3OPnTotXj+65yGSvbaSY9QNvltLU/+aEiUp91Y6cYt
oJpNnyu96/8TTrNGjQ1+B0RvIUhRr/ckGqu4q1R/i9+CYabWvxaqWCuUnB9MOxZ8
RQk5uGvpe0lW4EQqrr6OVfAwUE3ZReMJwesFzIP52s2h7VHZsQJG/GlheM4Zubgi
JgIzVYLwUVbWT/EFwQW/gGD7IHNydEMIWoRGlhrqZPzWGtPipWjIibr4SERjZbKl
Yx0ycARk7ePsfvdxV3gpoR5vtEryOLu0s8rn/2hF39N/gyhvmCCBVC+9uDF8sDNQ
RL1l5RxR01+roRsHaR7hTCsodZVPW963knaDlK9BscHdpN/DpuPuWJt85/7UVSDk
eMVa6WOYLR4LKpzxQAVb8Be2gydpE001djzifWKrpCVJVSLBuwXzgHz/3V8mO48P
g0PhOb5YJAJA6GpY05DFOsXIj3q2Yl9vr1ZhBb4lIF0Gne8wd5kUYW7HP6Axufo2
g9SpI7CvaZWVsaVprrbchxZ3Fx7IK8N1u9xXKGf2jAjYQHQdEpSeLLf1Wth6RAUu
4FGcv6F5RwDe5PQocbUDJtz/L4OQjVMh48CBWH8VSGFmVH+1UJ8e+967nJf/SVOx
0teO+S4Og5MF9v/UhFs2czvC4iVTICe7Fvxc2cR8Dpx4+f3FRNIoqgdGG+tQ+HIF
wpLM82i+gxqKDuNVuSHzm25f0s/NLEOtksJGDPL5xpaauwGVled/rQJKRMkulH6H
lUjalBgbo48jwlZSnf/JcWnw1wG3JDBbn50ijZ3TY4VUucKChOPwStMx/507CgGK
5upBbEwKdmfxg5QO3O2LmwK9RRGx04b0CNpTHVRIHCROfDWZz7qf7ZQbnGX3Z9G1
zGC20uVmZ7QYuuiA6X0WGHQwvEQvt3qiy0EuIisBzWFB50tqsfxRFs3f8VttRXIi
40GHPeqoNYjjHDCX1LqQCLLrGBRnWcJDNHVALwxH3rH7+KjSInf7azRqUrCmMRGe
R0pTzeNu0VRsMO+wKMI1SGXi7G1A2un/Ddn16bsioVQ+y+KuwpZjqoG9pZ7wHrl+
0Oo84zzbY4nPmLEzUJdohkvCXuScWX0beeN664kzvcrwQhpawMNzkMwvw3IdvoHo
yS3DlbQxNIDjog2VNuf9qb5aXg4gTTTIk1t+/1Hts1zn0PO21zvrdMUbiR0gX98V
RXxjHXzFBEsfBUv4HMV93+gZjFKwHEeCeD3vD5MEKfYYku9TWekrSxIJbFcQ6Gnr
WD5vdaMQL5UNUoPNIw1QS0cMtPYh1xCqQERNxJtK83ztfiyG8HSGzp2CHSxrWyOX
3fJCyjvqWRkERAVu6tROxnqCER0rUFFrhh42Y3b8eH/5q8ohX06dDj8WuKQtF5vB
2UAmcM/QfcSS6pk2lEzbR50fUnQlxNRVcUBXDLaF/mAcVZuvwcaJLyY2ska9Cv5S
5YBwsXevez6YQ0UohD/twvvxyE1x/5mK9MZJI9lF3pWYCnnfHpN/wq3uYcJDKMQF
3UrcyasgqLpYKHY4VR8Hu8UQXI3vRUqeMIZLsT6BcUqQH1ZkqZ9WjOMD3jq5iLRL
6AqJdr7be0ezuxl4dKJhW+Y2iFBoDhWu5ZVtW1GR9Z5oSo8BSAoPlU5ilpLlibm2
4O/nfPsY+qHeTgvzF+DvvR1MXpmM+LG6scUkv5sJbds2rUDTPw3vV2EtVgM2PopB
irKvOyzKeyQseGIzHSpk9ez5XptmuWxehxNYuVVz+doZU7nusvgocWYnybUyochW
gAcU07+lpTmSGl7uzRrvaBFo36YY/GbhIt3Ph9XQUjArWAyXXJSCMVYkTYxd3J8z
89A9a7uwnCffRMn8IHHGw4T/nLGf7sy/Sk7Of5hKBhmX8cemQqaHRnYXVB/t++PT
3lkUDLsTObryF/ueqxB1Sj82u2Wv3pmi3pAFTAOFcUxp0uMAA1MoVZazjwI4S0LS
tAK7C9WvJFtfq8oMYX8ZMNcZgaWRay/L5Uu+0IH8gEIPYPbbIS71Sw50lii7TVTF
Aiftew6CW0Xj2rupTuaAbk40FZz0drBKt04VAD6cQ28QcsWtp3BewVegT9PNO9bZ
QcC9yjQlxfsz9/gCuK/kzE68mG4Brqxt64gixM+k/OCArOMKEeVjv2pydY5oQaPw
wNfpmDYsNGglrHzMkTp8IIWwqW4AoExr5Nx0FEDWYJgW4O8ya7Z0aRsFqj5K4jqN
qP3X9w+pV3YzHO1KJ2RcXa/u/JHSbhogUQVWZnDmGgNn1RznZRAmShGdNtoRvZkU
/S2NGRncPF+7ptuG4HmtTPTFZPj81a9SLVpgpPjtzcacolpil5YhTus57MtqiLqq
mtFIyLYRwsOqqUtfnJcf4/o+rHN6Z/R+5ZVDhRlDijAHSHza/i5gK10UxZUy/OOd
aphJ5fv+AURdRASeiWuKeaURNjiYhlVHmG+a5/6LbQBeCWoLUaWS67uUmNEqyTmu
vbeqJT2Sr0i8I+B454RNqCRApzsGPBH0OLZdxRlVfHv6fYu17vURFthIPp0IyYAh
8eQMYpnUh5bSsHDcrs/XdlPXb8WQaebtqHX27M4q5V3GqeXdBfbUSR1DveW14fME
hsGyP2wE28lN/3dneTD7DvTxuRMmeMmb9zne/pKVFYyXVaHusQfg6p1njNSoQzHs
Zk4308BX70OQcJpgom9vElDtmV9zxq0P+yEVEpxoc6qlXDfbF/gfgDsnXJI3kGDe
HL/0Qo+XlYGZNKDKNzpb7Hb+SCEzwIuJrJYTdEQSXAL/iglHe+JFbdJNtkLfESxU
18ozkGeMqkFLIRZcA/M9zfK0UYUYNN14RrSRVYCLoaDWjRJlFseHpKc4JrGmQf0i
oyQaBb8MdAexF1bRSOVr3p12na1V2ball0/6TUTEobphsWZ279rK9utwYauXXUeq
eXsl6AAx79nQKHiSPc8916oTRU3joCsUdNmq7SqESUIPLJLGwEwnlXKuYe1LwYsL
LFgcoSSdWUPu7UY88Kx+AbFRpLWqRQmk8QBb+a5PQX2LQDVoY7YcYKX3vO6sUAfY
h3KfA1rnXm+yDPiOQYu29l2/d3m75ZYhcQAUtM2T+RGW+mrCxfsaPTwvPIZDHDOG
C/3kcHEAF1uLggdi02JYUmDpdGZo/jhQ8AJ2W0ei4khJug+CJjvNyuV2XCpJtwzb
EaXeYzWZZn2EeQlvcdy64soYXuiYujcQJvandJixwrvfLG7iOri0AAuDooq6jMUF
c1M02QN9l0m8W6go0u6KiRNWIFNMvAYM5BOlzzQKnhRXHPgRpzVQU5c+E5MVj/Jz
nojb8A49S9bZ7Nn42Nr6gQ2x0IHYbR9lz0y52zQe61fS7gxzBCurxolGjpIYK5gY
kBQMK8qPhDAf1zShXeFwqs/I0khs61qrwn6OOJqp6wzo0l5gxsnYoGdKK7GP3JOo
OJJPNdpSXWwp147598H2p8eoqC/LgrEkFp6RwsNax6kgvQPxjc4F+B/gw16a3z1x
wMQpDnc2aUfwJZ5EoiYGVFJte3bErfjSMO/YYTXJnpeLAHOUaGZkr5n3hRolpORZ
PbRz/WhHgzefXsigf4IjLXrXrGWgqAsgFSI7HJfm2mgP9/zbe6fLSiNumHKiyArE
2B6tS054rvwevSnpmpOH1DaTR8uS530T7gSPO9vtaB/QIFb8e5FHLmb6x5tdoPzb
Tj8JBZY94ke9xqquodcYgdt4GZFGjy5iu7at27cufmucJ9AsBYjIpw1hdoUF66AP
dUN97t4hTZpvaIwy3zNsArUME/6pRQboHXqEFiVZj7RfZhBh+Yzyi2AjVl97g4Ev
xtGojGvP3BjVeUfbz47xlFY4AUjXnC7cjRBXShdzBCqIN6dh4ambKix/QmEFcu6y
LdTvVDtTNhx6qR1GuW2Ay76l3caYXa+GcIPv7ZM2ROxF/VI7+PRFaYSShz2XXBC7
Xohal9qyEwL5V3fmYbVb9wPVaBjbvuNDf4NHzKHP70xDT38bhgdPGKU3+eAWq6dH
o+r6kGDgvTSabtyDG/ljJLu2yoVhTgkNFPR1gbe+6sN2tTWG8GqTO8Nug4nh+Fup
l0Yh9OOIM1Y40x1Tkm6COmb4zI3c6j4ImXtxLox8weRStE1ZzJHeypNNQjJ8iVtS
wRgLLvfw1Q0J9nTEMps1sLiiHum3rNaLICZyISEPPpJSPpg53MKNA9AOjLdEPAc9
jFXhEM2B2RHMtGqDb9wPyKpvrh1uuyjZ9CEprCyaop2ceOceXlyMJrf1vfiCzYik
M8VBpo/lRtmfeset7iPLy4mhDchQSVNwqUPprTMd8M/RWGL0pRGDkr4rznt84wlc
VHIl5d3ZnKHQDOIglUS4qoD6uvz/bIx7RQEzsSPkcck0sIivT8qJBjgsyjxE4P53
rCwD8CY2Xir5ikBLXxwkuqLKDPiZhV+Abk5C4D3vMbIH9NDqpdKfboaM6Db4vznT
ar9hULPS2IkG40kYlzUARIbYPJ2qoj5Rs7xkk7J7RPTp+VS86fySnzeYTWXwrXP5
l3ETJOMboo0YjXpjkhJyDYlU4PAYoA1wtUmd+6LzYXVmipqO3sLLSG/TA8d0PI8T
fSrgD+bReOINV0KuuaTVa4opctbrR+R/TStpB/wYIce8I/L2uiHU0knumG/Y2ONZ
6aXDaqbYgmU+Nj78OxUAZZ0nl4fadYIf+tKV7Jt/uNza3ipKBOFmNRoeuLFwftl/
gaeCHWSBpu0EKrfxvcd+ZCTdeXrwX0Pkn5lY/BzyklV+VjGDi0oTQQLzRBBuKYxs
eJRYLWn1kUAs4DapIOdAiYABWdiHz0NLQajiJtBzFV12S9Kd5oHddKgX9WOSPndy
N9yMmpBqBnKJFanR7zNzRbHUpkPJIQslMw53X2l3ftYkJkJAzaecfv1JD1GhMUyr
V6n8TQze6eR7upnt4XyABMAj3QVpfKYypxUs0rGrASAdom6cQ/Ev83opO3VHN5DM
xmhKgR8tmXzIMRbT6GE2w4V3s0r+yai/A5k1N1eqyfJLYFVg56pAxfWyp3AURPeC
55fF2/MS3YCy9s/8GfLvtjQ4iNArqsmfc20YOKzRMauhfDLSnj1ZDGqy//9yckZ5
yGnnxI5XivOxfXk2AnfUulEvpjf3h2ojrDGQtbGkuX0n9xocQb+dNMR8pDtke4q4
avreEVSPi4FBBm2NC0n/NVCk91uAhSK0kCiJL6CN/UxSO+8NzkJIN6fBPb6A4lm1
zUXw3i1/5Sbv6UpagW3P6Pnw5TTl5fM9SuvZZ/q+rxP0Xw8rThHzQvwxJ2bkmzSI
1Dvmsbwi/0zw0fC+FqXMZttXMgsKhP/9WUHcw7lgOtGPt6UMk+oalu2Tfag4kF2a
lXF8eU1M52sbVi8B7MmJm7y1r0K+G15tL9wsODB54f4=
`pragma protect end_protected
