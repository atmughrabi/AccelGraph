psl_gpi_inst : psl_gpi PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig
	);
