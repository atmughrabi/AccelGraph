// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lvZrMzK1isUoE8zpq7Fowi2bh0BYbRB6TC01y/2T/pOlhk8UXJUiPOxH1Onxw3J4
JJREf1uM90xo92QeoJccaFINmgHQMk+dHNWpMT+4uihYBEgkLVaMq5GPmbrY7cbd
Xe0TFfz8nTe4O1EUYUzRs8WQAz0otVQUfGeLnJf2734=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2976)
hyQJDZzm6v+T4VIJdhmUyHoqH+5O0euiYhHOM/Yfqol3jaKO7QVkG3Ni3VF2WsGZ
vUuzUkKkMFM9zITzKNKY3afxAxRk3t7Vu3bBJzJt7SjDQ3hpci26m7GUW7mQfWOD
jNrBJVX57NIxMNTQxPLzhZxwJejNfSzlMMkDeCFl4VBZm7QZxg1lAzpjq7GodjBC
Zf8P/GQkoiR/R7X8iYgLJ8okqET9Q00fOmmjV/Pe7xJE7GO4MeU6wBia4C/a9vAH
vYwrPPzWRIJjY8hc0zVXr3+aWKNC9P/4wWU7xW2laFS25Q0bsPz+0+MtbZBo3bSD
Bmp17aOQk2fCYYwrtlBy9iRnpwzZEp61tZOMikHH4wCddNhditu4MqeMIucsnBBm
4Jj92tm9HKdhuVure5CA4m5xcVNGV5G8U3tY4Emi2stl8QxHq+pXJPJo63ECzzbT
SayO3lbYov6YCsbT3aqVKszyalZc20ezwnk8i83dSrleYcrosKmWplpWHg1d0at5
+yiS6xsDho6mP4trHk2ntufYm2LnRxchhSJVABiUfgDxTzDuFfs8TJPWsNKdA1Sy
3HzD34u/cRkfI0Rovt2CUfit2FEVYn5krqHCHvNeiXiHf+N3qOjiAU2US1830n1I
cp3hiirmNzdbMG6dao/rYLFMWDUBz+I+T5Q/vRhrvczH2b3GFOfKZIqv6GyGIz1g
ZOpP/Lb8wxaz0NhuJVSZKbAJ/umycgdGN3+18g+APNO80YpGYNBB7Qw88H/YMifD
qXUNWBsBvxOdSHexEmiomRJYVHJTwnNKOTmrTTPi6E39Dh7eA5ExItwOxD4uxdYV
PKTM1a3uEO3qKH82mGl9LWHWZw33X80tdh6MrVCCUjlzQtXk6aTnoQCp/Kk1DQ/N
TyfXSCjQS2Xw51bpSw+eOOI/ak8ETQlbmKOiI1q/hprJTTeJkF/1J/zNAkCy8PdC
4cORCyC/2VFoD69XHhRek40Pysb5VwbtXBuQkctlRmPNLJ+unDEBnBNuyRiaylJi
40Hg1Lo8obIFgkzdS11U2DzLZaqTjT8vyh9cJCvrmxLA2bIxL58Ksj3DDirrjzDd
qxQO23Z1CG19f9GwsauV8yDHSHr7c+GBLrVRzN5AOzz9s6fAmKwlrEjghx7Y91kO
VBhPmcmuVcuoIJ2vVfpqXU3USgQGgBoVueF3/NJl6+qhat/YhiwnVPB7tbgE04kn
85MRO2zOBe0eFEEDw9HdY0AH46D24Oi2hfAm9lDPIYqx0NDOylzu/uKbYs/823VV
r9dUyBtXcmyDK13RblSjibbLMlxPcKYs0qLawpOTvxEOjOT472XDBTRJwSmCq/GK
LpFAoBexw9f/qlpEAQeDkSeEi78GqPN8rrKin8KJNCmcF3aCKn0oCk6OCSft4RRW
aC01lgErwMsfm/p1fiYINAHf+rz3bW0uoll4/lZVsrUNhrkm4ZG0oY4bMAfymMfZ
6Q7mMDIpRPlGxQ4ytEIR5kq93yvPMFL7tsxX7kR7XIsLD2KIt9VrK6GfqiFazmHw
IPs4Z71vy48t3HeIxquM+Ixnd+Ip9gNfXnIAD6lG+p3gVMD38khXPfrNSlEcH9Sh
pIrFBOxlDneDwyWTLSJ792d6AFSk6za8YaMWF5xgbWkoan1LNagzrtAs82AK0bFa
xN8W4oBrBwAiJDLgCeLHswW/5nbPY8/m5APVnVKnXSGVB7N0jmkod9s2XuumLknV
4hg6LSo379cEse6pPPsKihlnylIQOFNoL5yxWAK0jS2gM7nxtrZwzxYqqHZErmWk
eTjfqaerGl6fC4zhNJFGTU/jQZBUGxWdUI9F436AbcH6onRhBq7Wh33CHt32pjG1
wFsv9pe9rvt62Se3baKQE+pgh2mOdG2gNUOcUq4K60NvAR3VM9cAj39yoAByUQxR
Cf0Mg3jMIh9sMLlJiJhXk6v62m662yZ/gvU1UdpHzs4Gf+nSH6HW1opJmJzYWi0j
b7cRKlvCq4fDEzr8hlvoRTbH2g2LK7kwBNNMBezo7g2VKCkgISdZSXjecUU1rqNG
eFmF8miaePai6mKikXrBWhLzjf4bC5bkJVg9dRQLAllecu53NmW7EaThu98hsMVE
aMMUCbdkrxqKpy+twg7DkoolLXN3woNUp2VKL1hOROcChiWY5+THfPrxQ6px5EGI
uAm8xN16BIL/bahawcNY/J3ldSOv+NWMQ0tuBLGo08QC3UX13Z9ggivxvoUtaDF8
jEnbFI0oP9n/CymGK4egQEc/4CKlCAcN2dMeB0VSUl47MNYIrENg68BFQrFO/7oG
fhY6z3kl/SU8qQZzySolzLE3+WVKJhhYvJsdB40te5/ypirF4va5i9RBjKouf/TH
fNUeOfYbhy9uauzKJBZbqXNLB2zQDifJ2f2S+Dusdthe94wVTRHSULTIe54ibgZc
hny3qDkBKu6sk0a8RQoM94CU6BEz8iBf7I1MgFniiUe5MaBriaFYG8CdHk+Tl4DQ
p0LIlF2DaHZYhFNGyC8E2Sx6ubRv4Gk8t5sP9iykbphmXlyckGyqiR2ieuDFIvxH
rrrUq4LEFZNeBORhxL2/4/tRCPEL9S7JrrWbgyX2QTCwLFg6OS/dH84stpMNyUoe
++74Aq+IL6pOj/vLnDJfn7JgRcn4r2vS9nGTxCVDadx2iVt0/m0rVwpgv2J+gnnM
FvlLk//Jd0/BM90SlESK/LvYLnuf0cQo+Z0dNv5Pp4EoJZhHqyVNzssb2VVSAcz1
41nS7wTrTcj9ZyvAL7pNrtTF8YpVngO/gUe82/6aubUMmok7xLvWPbPojHZ2F7LI
BpmEVyO52Z/JH8W2ezHRPP+qclUNB7J1qlim9pwpOFbRTaYAw/BDYpTeaXyBApBG
v4mNeQRQ4Hyojt5SoD90Wquvw3Pb4UvEO17pdswVjkPUrqS6DbTZIsNfChFLKRdj
Mf53hD4qsDHhOnAfqD1gDOu8FAspstmW4+4g7vIHFawK65u/qb62JE3t9811IDwe
K4LQEB5BHJ0RmiOaR9UP7aMGsJULgUk3NCjtSRpZ9w5mW8ZFgZdsXGsvMPe/ZI2Y
xC8lLhzQZSFf1MOUT8nq2O9Y4mpNsb07x/Za+ouYla7y70VHLzOuQ2i1soK3ZoyY
zTGWr+33QKAYNSDwxa7+pTtl9J5expUPzEjC89ta91ZW91img7OyQ21F5KHYe+6e
eLDHUuhFbkt7tmdtTbgdATzIxjzNq2sSZpzewe6fDEJw/v457w4WG0QMYAAdt6Sw
jtz7ssx4tj/hKLoZvx4NAPqGBUEoBTn16hKtoSiSV+pBRb6DdiOxZr1tBw3iu4OU
ae4/inaS7sK6GK1SanOeZ1kT7QsqOHgsQlnWtjnF7vCBaOMhnaMgxcxcDst2/nCU
FUbK2dE5DnyFMfiEsp8NpfmgSxpB+CczWPELuqWcehhsjUac3UcYgdrhoyGhg2FF
GPI0aw9tAubMX01GUaOiOked1FGmuGArAsl7Rf0aGj84Ta7u5raAAMZWVRTWbjYj
rhY9aGTc3Spa+YiwZr0/tSaGSYY1OT5Hutbtn4SfB6rALk66uUuYarrOIBBaKmyE
dx+yL+py+O7iMVsHMCaKIPwtFb3HKnSY4fEnbndM8YHopGiOqTQXn9oJ/Uuci704
W7XqhDYIu9CaKcSydeQGI58uSqD2Gh/yn7pXsIaFPMRLkWy22Kom4LJCmAp1lgdB
exBxP3rqgeiZM8h91lo8DWQbdlw8LszZq75CS5amYhznpKJDy6AIis/31tDDi2xU
NF7WO5Ghedw8R/ySTKWVQkztKY919EQqLODy16UAbP11/7NMyXHtjs235yDOuTWj
fkhExJVHYP6tfI2lBRiKH93l+BARNqQ1f/X9bI/BsHwTBOhCNYl6f/VbNBQo2SHv
kIUOQRGz8d4oVpdxvQnQITufMkjTmP4yZtvxzPQF7vN82ZFWDaIgfSWw+i+7S7fO
`pragma protect end_protected
