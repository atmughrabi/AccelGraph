// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hqJcCy4kJEBJB/q3f/n5N5RhIiYk/7gN3MyohrUafcklJrd+t02jrFsOz5G2OO5f
iDbjCnlA2HuxUxFpHlALbTMBbSbCvPcIWCfn3OdWgrIGSCTo59rTeZyi01yPLjVE
ApkAn6dtEUKdX2qFtSZjAmOTXsGINillHosCh/5R2TM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 319824)
CzwuOyF5Y5kH6WrHVQMERyFn2GXkilyOsa6TnqcsSkFqQ+q32+kG9m/YSLc28kqq
ITD/XiKpGg0b0s6aExA3X7K8/lt+O/hoVwHNtBlD+IWlGgbappFrb3IgPdjIBxLt
w+FoU3UGw65fql0VuE2Q18vAl4ig4Wc4NfzK5SdxR8SAF0gMKlOhr7gOGuVS3/C7
lZ7TxBOOYR0Tns4eu4HVpBP/aaToEQTqFJdaYriGzkOWI98ZuUkk+kcoY1k0bmvo
0tmxLtcGlzj69GOiP9aTjR6ssO01CkF+dnKMU19XW5Vrt3cIHfEgBoKb1X4uvABo
35tlW6TCdyT2BLvd+WRMwSaWzMH7s0dgMEniN2ba1n1DbibZZRbym8kcouIzsui4
5GczjeN5zOBkBarwQXYxNgm7HKoeZoirEUV3Um+I3jqU4BlxZzrTPvq1I7TwMjUT
hFDVSqZXuagnBuv7HCJYYoK6apowg2RKauI1aGQKExfip+bw732IhpW4na5tpprO
FTE0yz6zKkbSxxDJtWO5Coh9Y92J1ZIoQZY44tg2Cgl/Lgi0lj1rgvjm6QfFBFkF
xaels4NYA7HG0T8cbe0hE5zLuRTubmri0uluepvbO2gJbBh9XRCVsor6WDTdRA9/
JWWYsKEX0eQVRLAcn0M//p/o6GVHifGTaZikLKqOI8hkn84kbsMB4xSr3u04rlnN
MroZJQ/RfMwTTUhTvWAHFrsEdhbHRH9cvuPGa4p708kklqSelsmicVbKqx8C3z4J
7yLj8j33Eap0oBWndW/jqYalyULtges0X1Hy3tVptGgE0TGuaDmnmPpjVbeiHXBh
KoriB4YO+lJs2HQL6ANveAHMpSuR5Yq08IwEtst0LbxKNpj1OnZl121B4X8aPKTZ
cc6v8Ewws/k/RFTJTe36NLBP9JhckuIYCsqcykdHJBAC1/6qZ3Wg+VHfY3yVEx2y
sntUahHnNUeTztqhie/iiPYhwWTXoHuK/mY2ljU/GfzAEvXV1Hoj1CqDxycd2RB4
BCIMS9BKcAK/OXUu8aBQIXrmg9o7Mromc0TUDhrOLNA8gd87vLhbcqm5l/gJ0L98
ekgBOyF9IL1Yk8zJ2KsvynVDSI5VeTKbp/j2szYDuhlF/WkABthoF/bKHeKmjPWl
WTx2Xwuz6ElNMORaYcHR0Ii3dmw8fN94d1pA5jaPPrrGPejQk3WawlNae9nHUKPG
RIKmvHIUfeW7rIxsERKdVP1Zl4VRnV7YTLtup+Zpeoa7oUk1jmhUeTjmD6Ub3q5e
qSp9a8zJ22kYq36CzI6TuoTIP3LzP3dHXJhF8CY3K3QtoH6+bHJGdzsLmsrK9AcX
NbH4ofLn4zPHDYtW67UvAsuvLQcbqJhRdJk11kb48nJbqmsCCOkiI+ddY+nLBSYP
/l77Dm0FP6N239kAJkKY3qSEnhfyP7A4ULaqNKTv0vqHyl9Cpkhe1Ias6nuw2Frx
RDxOUsoAlhgDrKas4WLJ1BFjdvpGkcSaOE3QWLg3OrsPBAXEDXD1sas+WatV6RwP
k/hOxT/PNRv6o/Rbcx7gRZAL8QdH1+1rtxsW8TYpFwRWEFW+0ksPmUeo7Cd9Th04
iw/njNgjalM8eOSF3NoyaTj7xgwTnb2SBxA/hrUvy6cdPBvJKnuF+XZIjMNuyBkE
v4p3GN92fEDwTWLisQFIsd3M8xa0p4g7Cgq7I83gFD9X4VT7R6Xe4CMq+dmcBaBK
Wf5ehE3nwIMFoWKZZoi3O8l+g2SgQj342IYt62gK7IyOkhh900CAoNERSugHbaqn
0X8Q0zjdbbWxXMae3e2XA42qqms5LcYAyIPwU/d4PZfkHickbKoFm9Q9bHFVr0Li
jf75VQgBQhwk44mPBCaazSqkBgN4uW8sbNZ3jo+GQVCVKXhVbaTyCy6e+hPimU8y
uOHZb68SIsiLYV5+3gA3vhcTsVdN/knMUCyB1iwvdxIegsdPeqpYFUCNmNVGajGp
Yo+yeX36ydkKVmdfH70vTr6JyNyFJM2/PhRu4YZ/018TaBfEmA14uLukvFSpAlkb
6Jw7rgQ95PKMVE0B1KHKVTFgrnneggR/m3cD1aTLLL3UN0jYCeiIQJyctyld/X/0
T1UiYwacMXkUyhWHhFXyC+8JdfEC/++nlHQ13zhB2bQcMIcMzfeFvmbIZUNadMUV
X7Wo0R4AZ5ImNqgcUwNVL+7PAu7v7LwdwhKrCVAXNWLnNUSvUIgQ0pjX0kPFa+9D
oM6fq3rIbAD2vHmyBcUNrpYkoXSMlKNauMAq7/b+4/MPOJuqbwU+d5m4qEE0QoHo
4kuL735E/Ev+6gp9UP7urnNnz5y+jYoiV71DXt6vwnEMpkBMO0a9R4TjYjTXk9/y
F68hHvE7KyZZrn3bcN3pWrBTOuG5QodVUmZboBHLRUG8XHI4gfPb0Qw42eg01pcv
FPWjaleuhttdSMJ0mnDF2ubUyyAO6k85hCBJACp3qRNjRqBUZmYcJ6XtGqIqxoQa
5Psrr8Yjqsu8ibj9MCIRyhrk/i2t1T11Rup/N1EGLAJ1B/aMzCMy9sOS66uFu3ua
xDoibd7VvecOv1l5+bwDX9nZnWbT7VRWeWqu6w3jza00As0ram8EyevyxiHNN4h+
E2N7WeMQ/DmM4JvwDtGeZSDXuu6XDuGDTBoCuK9Tp+OzIp/2/A3Gk35osPyZeki9
qj/b4Yn0ekWDRIY4nX3DTdqAbbsFxXpHv/tVzizb8tQwSuCFGR3WV2loIA/AvdnX
f0w1F3FFU7DlfBXJ7KDAJ5fPooHzzm1Fo5tOrLMooByKnM19ceypLhTXlmIO7Aat
xN+d61TzB+6CuBb1yBYu7mwt+m/AL3KAeq4g/iMmJMJ78gAQFnCHouxiZ65WrMCK
HP9QoM3p65i/fBnK2IxEPmFn1UsG9UudEeOR9eKUMPTon1ComCCi1l1jyci2mTlj
O2vAaktpyrx0VkLHVlZhw42f+shGFSFiB3Hd9LHLyhrW1aXj22LPPbk+ko1bxVrq
mH+bz81q8I2eZBwYeNK6GUs8vb/79Syns3RMrzMD7AOQWmJb/vl5bZJw9kjXQ20m
pPBkgyYF7i8mhoelFf6SxWQeBOukAeC4DhzlnGfLwvAm3xSyrj5Og3k8ZKJPv2yY
vxaMPfpt+Qr3vVKywkbYK96mJsH/385iGzdBYvBuEYjipverT43z3eDvLRCp5e13
K6UG4fwjv5+ACbA7cwXSx3z0zSjSrnOo2SLpZdPMuZBQxwywkZbDlrSoah0YIcYE
inNTs/VPVCVo9iCVOAjhQYmSI2k2qVO+NNB80txlEFB5qJMzIy2Z0ciccNCBeMiJ
D4a5MlHkAWCWdyrpycmVA2eSfYPCbtH7Mpm+3nqFWSH6iSF3MVOLROHpewm3JwPs
OOFtssMfHN8YUKO22JbBeeDhMRMX6gL6OSQ0/rUdhdkVPen3EG3OedBFslOCjV4l
SAMgSPyiZTZT9OSQ5STM0HsViV6DcAtdfbJ5mikYq62fsDxVlsjn4k3SKiNIIzth
DfZq6h/J0ExcEbPaSvnevan4/VNnu8+HAEhwUX+Dd31x4BOkhJySKm6YWxHiIQj2
XGr4lacmHsyUfw2nf3B9TOIglTBTlGu+12VPyDr2twPf1CrD1xP5bJhqttOh3xBe
Uv/XFV2xv0T2soWqa3AzF3zXzJL6B+TGB4mGsMaMB+5L/WvgF5+MMFqkbWObgiMO
m8/LTIQz3SKnid+6XEXVUXisSiqEmGgKdq8tnJ7KeF478qHec7UNNrPUOiTu7ydE
7kFOWStPk/OPjIL1pcrZXq2SgTULajAXrHvownqYZ8ogLbUcrIkNZJyD9IM9fsF4
7uTOCU3U0IzYSSg3IvBVzyTx88lBg4syuNlgFdHbA0t8nd7urymdydhmugDXcvwz
nM5ReoffQg2H04yOqJlGWZzjDploZ6wBjxzjeYkjhrAbUgm6sGrSG6gkhjZa5oIy
wxEaqUVZGzs9/WEPXHAZw/GbNlNI2yNpY4HxxcXqygLOVF12pDjff2ytoEGyDwJT
wyWBKVHrIccpr0ymBhv87zF+6HFLnR1kodYOGaDDnI5FZG0DtWO3lzx1iNbtiKbb
FyXFmbyHIPFIoIH36greuC42eGurGNLrLyC7q20LOeYRh5S7sfD+hUDNYrYeJb2D
Los6IqJz/DLANjvQY3rRRzAbOm9rEkLt1S3aEfdXRwlOAVo241hVb7Np7MYj04ZA
OoZFMuuBvQgncjyR5FBIKFeMO/yuYss8PFS8tqG4KP/dVykjLv5Op6CFZWhZHaMF
oPLOak3mAtQs5B6a2PmsJOWwng7Ui9wcoo5wcwIBxpVYiNyXgQz7YoYV72RRDpag
qnxN3to00URZuJZKrH6dQip3AK8swV5WlOtLH1+gT9pY1UtPI1+MERqe5MfI7/sG
3VkM1flaSMrpfMLhwRs+sfStlA6JLSXMVkMK6cqY4HgxqQ2uqXWXR+eRdb4nnVBS
+QR/jhUmypcu0WVOBmXOZwTxzLYjkvJ5hEUbu9EvqlLP6BQn6ETFV4DSW0DA1gfB
yavWHyrW8Tl3L/YL9qMOcZ6p+S0HWSaChajWEAGs4zKuh3eVO2T+6Ppu/yNcRhX+
6VqBIRWp+Km5UNeYVJo9GvICcnR0P7XA0xNX459kfd+xC/bwZ4AjtNTBmDPaF8qy
FaLuZ44idKl5lm+Yjb0u1HyUjxmCzyUxWzK87yB0uQeItLJeW7FPbc6AYyoPhYOa
lEPMTJ75A0FN4OCNnNfAnblxG3FFXmQ6pV8w20CmfKPgjOGL9d0qxbQOI3I9NNzS
oZX5PAi1gWGBBv+2UaYk+C5fNzqlK5sZCcGCl8Wp97sBLUGPlQiA2IZhNx5Rb8Y0
1ZLsp8VzglZSgtd//B3QtVJEcWhNNBekWe9TCjzlQlP3kVn+LXI05R6wPpS63HhB
SUnOejGA48eHDSr/1r1BaE7LoALQbX55jF5isVvKTgtmwxmUUKpU6g5vrcQN4HTb
AFLm37kRRdw348W1X8tWenllMgT0zxgEhJ3tw+1BkzPJQK/isB2DnrQQWhVI2/w5
g0mk8u/aR3Xtjpi/zahHl4AodhJXFuWrdA3zY4Z9aR/1ZN1rCADvP7QmiMGEehb9
SjF6n5IaKyxFETeZzjT8GsLj6jPK7yspeEpTcYZaupsRQ3n9SNlmO++ONIU8Xryt
ug63yua0RzuUKPvvtzqEjLyAhsSIasCXAooBTEPcFC++ac1wgBybLN+GDPOrKA2M
+T0T8EeO/+PD17rGnK0Z6qYe18JOvZ3R2tVqIuQZ4JJtWze1Y2OlSpXCxwOVwxix
O7t/wwRxn34vsjr14ONMwDl/KYtT19N4oETyQAPAd/VVWP09H6EAQhqUn9lWibjo
Z7jf5UUqD4tDDxIM0fSB0DJtYq4EIQA09vStdMAFYIE5YhFGE7al7U8gXLWScgvp
c3j0yWivnl5BYNWEDyQLG9/OeHIVDgP6ToHpbQw7ciq6pn6GCs95ZTt7RhO6enKj
+hEroFqg2cg8k67xs7TLzoNRT6tSlfMMEo/vTHp3Tv9/t99A9n3nQibxQyKdEkgH
iChmGx60cAEFXIF0VT00V/TlrPSkaV4Jy+J9PsJziDULTczzT3fuKFse2GjEHvwd
lzlw8CJyvifdteW106xlfncaMAslyXDhVA7NCCruGhrodSWS6UVRQRON9ZkXUvJk
IQo6lRLgkEIiGCO8eS67tngQWwXGSF+JFCWIj+9gjKJTQwgZmSuzNL3BYorUMhEZ
jckpbIDdsTS0jP6940d5myAd2+YVUSKDOU+Jk6nGbvO3v8vMROYfZKB5wQFSoar/
OwQdGmdCSGt50j/l3yT30InUNsdBz8tyHJbyJGrBD50Yd/V55Jb7UgEmZXCkOC8Q
7WFa5SnIA9c4j7NQr8Ul4a/tqAzJK1uYWs4/kRi0qgmPldkq5bAt8wTEIFSuzevJ
xMnGU+UiQ/BT46NQGJ1rPfKgv1zGl8XRym/PnEYGvsG5CVr0DdUYWMJJq/9+GdQ1
lrWJDENF5ilPK15Ux+rtl52/CqDUntI3eCDBwODJyfvvZpi0WZIZvFEpNCZL4l2F
QOHqQ4Wmb88y9hqUSRiueyyVLWUfyueK1cZgKTs8L7BoP4BJnoQ2NHkIQV2syphh
r85N/zxMinH/eDZHL/TEpSzOOpExdIcpNBHXQqg1FzO5GdrH0k0U9R3reZXRNJny
X+dSUPK8njN/2/9sRJVCv6H+FqinjxMLAJ3ZZtlYZ2BUB4xXjezuIQn4gBIo2Pyl
YmmSG7qJhcKi0Rb7/8kyCsXEByu+rYm6lyBy3MZ9iQ6DLI18j1GeRDGTyDmEqrJO
33g6Wn0bAwsrOtkzTFTqovnh66JUzfKqH9JfRRoISOxc8O0BGSQSE4aLBFS+l1Ra
Fw9TgtiAHOcSiuEW7aawycEm6rLnk2mPMqgVVvniJvh4jbk9NZvB+92Xq76StO0P
Vmb4DnfGvFWSVVAy9yTnbnH0fD0CiNlaZDvZTQM5edgXSiskzf0gPPHKuXjQgLGZ
oHDwZiEO6EItoDfqycqPE/xaAaTIaY1u5ks+UsG1TYrbjwxel4ObbSI4jxqTjagF
11LGPDGo+LDqFJhL/ZzxDyLD8HCs5FcvzeRbF1WM5naiZTJfsF2LbLPAMTg5tFfe
siquoW4Yt2SebrN2DKcVi6BT4dBKo2Dy1BLIvH6tSDeSLJ2baMsrNVuJiHy+pwHF
hQLqeqz4pgWw+GQ3ZqovelR/ofsT0EDLbVdCBErow9/nQfzWvadCP8DGjIpUZBLI
NbdQ5zFozV35BfbY3f4oAp++nrpm9LXzJUo4VB0IOL4MdWGEer6ImruC6egwhfo/
7VTfEg1WX8evixBRsYTPSjJqxHwO8Qwta2dmwvUgIVswOnaxHkqsmo+Fjm7SZc2N
IiuNSp+WZMxEOT1coM3E0WcdS5pkzCVnYEnWXGEFJfPGjQt6c6P4tcpiGlB6fSkH
kYUn94QDuqP4RbqGRAXmxcrtYdsxw2RPoBWwyvhQBxrE8QKutYVkwdiZFiR6oR0p
QHmL8xbxr/1WR4C81t3MZ8Q7GkaRv647dp+1Jr830lJ46GywHw/6jmCq0obsi+p3
lVaU9RsotT0DuBWxkeL59qIlIqcZo6sQkxXFhVvjThoM/uwQh1tgKhgLX4HMT2TJ
Gt7qHOpMcfwMfvoucj9vdY6CWX68uVczUDcHfWs9n+TTDCO6CJE4RXNMs+8I/OXN
368q7f0RwO0dooNA2231GEEdJU0LfC6pcZ80zBGPrc9b79fN+e6AuTczeRlw4FzX
G4KPv+CYZqP6DoOBqIkjKymgjwXN7WQUb8ViFG2Bmvl8zMDyXm34kbrtkhQvzXHC
9pQCE3oHqlpO2nqQrQPR5B5WeTKRJRL4IcNWrMiBvOcOF4sN+OwxhoZwTi1zulqk
T2h1pFjJskBKVrNmMQsqNDkPEn+OUaua9lPwPIF6D+qhkbbDr+7SiU9cDUrUIBE4
/7givJXVLO51/RptBez/CMxrAst0GUMvvuCCre2kNNczTHwc+l7zBjMkNVBzvjn1
GzaxOz4J0do3lW9yP/s2/h4gUO4Hh1bfi+gA3IOlz8vQX7ZsgNJoALw6acnn+VOk
kldOt1reROXWa/RAqZqpztwPd0OqwnlsdJs6FZbf+MfmxuU/ySQkIRbdS8Pem1OB
2CoosPl9AG2JuWF/GwG7TxvvbneNCHWgfFpM7Uwj3TBlwe2+2iub0g5X8/37vjct
D7rDTJYy4cd9NwPEt5JVkW5FVVlMFloHaE09DgX8DU/X8E6LrlWWqvXBQDwcg1xg
VgXTbqWGE/X0Vwaep1IvTVe53q7VrNFUNEwtjqi0pZyH3S8jBIApkWdETYSbIQ+8
tvWoDrqtNioRj5Gk89UqkWOHsc2MIMCB69KdLDbbRz0+G9PparVzvaS+Wb2iIo7I
wc6GXFJDTjdLuDS0tSATQ+lTNUKyuODhwMjYBS6vNZluWhQMIvbR6BCS9nME3nO7
btjjHBcsBDbu5BpyVOWkLRbQ+4NFuHY/sLEU3KY59z6TPp4jIEAnjrEM7ghgRcP5
TUjj7jgyBf72hGjSeKJKH45xPfWNxeMGpg9eCuKuC7vYzuQL3yNlcmcH24zTk1VI
d4WWJ2tPBytui8Gn2bf83hbUP1poUkZ/HeqSVFZROAjqEWxbtCMo5PEVbjuK3aDR
IHyvd0dButMoeGQJHyzq+/x7uXnEh7G2fBq5jbNvg4g3U/SiQZwGAEwrkTb3IJtd
VzFSIp2/Hlg7HkHwA6Z8MBJv2t3oT+GGFXNZ7VUpKVYBo/JPXq/rd65d252rHHZp
r3/R3B/vUVjtlxFnaKEPGDhI5YftdeUqn6jLvlJ/xgwQR97tWos7b2YmVvkGuJLq
fo2x+MDYsweoMA8wv9pgQHfdlolLxBbyz1q8E/+yr4sAZqjp+YFcrHxXbHub3USS
kBcYjQ84aEjRhkgKj7+bbnYLK9KaNaw57Uhj77KWh7ukOr0Wgv67B7rbHwY+/feB
0zeQfjTgDr7VokscTQuXhEi464Vi55EPDlHngxwvcDJ+qV7Pteay1+K0I38hakyu
7QTmlPpe/tscv3j7AGj3sf4i07QqN7rg1Stx0n7TMxQq0Moht7TJL2sr/DFmxD78
WfaS/5cZYpAg7gFx4tNwkOp7VmbphxmpP3JEYHO2SSsuf3LylpR6rkkar4YkdN39
z/br1nGsUtwbUOmGXdb7LaopLwRc1wy9k9qYpJkx2asCjxryu3wnZU4y5mUDJRdV
pKH7dQPFhNCS0zzfbyudgEo91hI7bsfmiOaDBjJ0Q2vSWg0t6steDGJ8nEHFai/7
QQCKElB3cX90i0hVpTZjbkZzAL+DHLuTsHLreoPILZwYs6kmCOEHN8H8R5vCXO9/
owPKISJwiVqYVFjSheGu4lcpIOtgY/9DVdqB/0+udad1L+RCYE+GIyye8Xr64dET
fQbRM3aei/CSyLlPtVHKvUCkmVba0rLL+UkE55cBbU5B4ZcnCMsNTRrQ77J9jaQU
/3aHGxgkBS3rMKz4yX3VA+wI68lb/vRj5sEC42rlmdawSFF2O+i0zNywOlSznpFX
EzkAoNH/WI0opYbcGbllCse83dvDWXGNcyp+kUkC64HUYKPkGhCBVgriAkHYUs33
QOebsDs37AE0YplzzyPYnvb9A0MDvgGnSlG0vogQepeZCbgxFRfIVFzR9SbhEcMM
m6DJ4bjhzsF1oeCb2CVYRbMK+ok7rwNiTGUhW1S5E1NCjTkmGaaozP3EOF22wa6c
Js/wKKB6CrQCetmNtukHNhXlK76++e6bFO8hr/hr32O/RNk7r+hdXKpT381D/WPt
ZaF9oBeWv+YmME18BiMJ1yhGz1oaVTUctYZJahcihvois0qQ834CCltWoVMRYdxq
CLcEFhlwg89m9C5vTYvn3Zahtnje/co58YCSwNxS1V2bMr7RkJuIisX9PcUj6D7R
8hEAFlPCUp/OZoFhWTYGaUZ5atSBUzt/p5OIiVVy5L4Sw3Ln2/FUCFBpewtewX4A
y7W9qkk3w6O1rxK+nb/dSFSqteW2t0QGT2Q20wrFI9S7ajWvclTZ9za0fVvMOuPL
V7Ne3+n2xZhYDMhDtsOE/8DFceCM7gLtEjOdq3NxcEZ1FgnUuMHmjRQurBTHXK9D
7UQbvKY0SejKC/ub0L9sHI2fj92vDQ1M1OnioQplpVhKc5mJq6ZboXEpKGhtFxOf
aMGj86f7AdfTarODyuFY0oH6cbM1gp+ZyU5xW+OjNix/n+Ac93bJVcufc9Pf+rkq
W3W0XqtKaiqv6uj63Z82Inq329TuG+qDfZl6PH72jlbpcr78Es4yciWGRLJAyLg7
M2TzVvHJB8D58Q8yii08aHQYKauHcDB54AgKS4ooeKr2sF8pn7Q1SbXxc95RjI0z
QSgVFroaCa5MwT4azJi+aPj8kdWrmVK6MfBj9wUpS5qqMmVYPCcSwt1Qgy5dnk/C
kOZobr8EDjVLxa+KgHVdoosFhmXEip3j5Tqql7xe0Nqk2LpramBXqiPqdmOLPVY8
9jTUrLtIpxmMqu33bRjbc+YnjNhCn6ObQO21n+YiEJSnUvOz6dRZYXDs5B0J+xhq
FPWMA6mA1lTVKIlYD9CeVsSTZwhjlJ2s8qNKhxqOk3b9pjKtOkxoLAa6gpWWO6XF
wusz0GKzx9Zmd+049NgPwU54M0Tw0OCtifrxfeY0dMed3bSTM6MVLZfWu42iQDSj
OyC52UR9c6Mypbh14/pr6IbiZm91PhEtMS8BFY5h/lX72teD/renBacjmRTZpQjT
d/av3xJBV8aFU4uKuTBkcoGlGnmuHBnI8k7HY2aY3mhenQ2sdw4WJy+j4zn4pufG
npldtPNcrIpVESbQ9MEpf52+r0xprjE+gkr5NQ9+EcwF1F6xFv4niM3w4NtHif2C
UZXjPrNaiNJ8X0I9GtMNWvKRv2/2bQckZiaxpTCgVR9lqDcGrY9UoEok+kWflYir
YbVvZJ8GtbATpYjl/1N6Y6eatiEKaNkzMIko8ghn3P7HvtsRcuBNQA5xiqA+BdZo
50aU5PPsrKjJACsa6l+fUbXP42u1hBF6JFw43+aJhSz1itmLO2JfC0KZzi0wMZL0
29jJGy8pZHk3x/6qPKrm8NqiawlGLKp4baM1FPk5MirT4LY3TdC9F7ZjseQTZnXO
7yHxRKZdp39ow39PuuYkt2miz5vl9k/kiQVcIrAyJgbIHFYdhhRJwTWJS7IYTZDn
iOxmWR8PySvNvKJRsu8CQ2L5UJ0ILlgSjBwsSG3dBXgQXhqfTeN20jyzQYYKk607
nXCxkiPhPYXM1k0TcCb6Ktej2ht4wVFbYRAnh/7XkF4j3Sm8DOxIODxjuFDWa0D8
2/lBGOvyXwlBaUQvJaMFUGnC/gTd8tXYl7d5X4KFtI7ollUPAUq03BD0wJLGzXOv
gj+0rL7ymnTE92sf5RP7tdzOqkhgO6J48nWcnMXIS70aAXiQT9u2z/gUFNIKDelr
YWymgmewiNk87ZUuxW31mLtYfvD3Xhw7vvavSOt/mvj6ok+L1rH0CcI3UhXA8008
dq+mY7doEO/ZUsA+2gmiTydEqLlkHdmVnTUlANrEjSk+pf6ixxVoP5L2AwLMLW/3
Yortk3IDLAI0VY65ZKBvw4R5n5x58CHHxwkqibJXOwxQrWRzOtZQojuvmI+givq0
XQ9Hwh94D49xfZhsBbSwg6oKjT8ZMioydqo16pirZqB+FhvNR5N7v0bj6/1DAw/X
jxl23qlwcrzSZAgAc3rdrM38CpxuJKwUDp0tW+DM1As7SFW4DqwJ9ipjaUIUfSCk
ReIfkGno1u3xVNqjFlqa9AhHGRD66FC+X2e7majQ96chgf6i0LI0Lbo6TnrvS44y
+okXLhA7XIFJlSS3XpsVrSzfzCtQYe7P2Q6IkHdyk5SJgl2iAIHxV1f4vyvgGh1j
qDK/mGHpeIEV638YYHM4cS46nKexgRhkC3Zuy2G3l8DYqYCWD3kcWHZYKEs2H6Le
NuEbT1E6MxVnFDmTAzTS1g3NNxCheyWvw8wNcygK0+tH1+n04+AGlfEgktYNiQPB
Qfp6+YE0SppvkX3Ot58LreCIDg8al2JSvcJwsWnCdHmmX57s4XMI8pz9N/jwU7qJ
y+xz2Ps4Xg23g5GxND/cONfV7ymCbnOcjq+f9TUkVrnUYAb2Mvo6birkftqLH5J3
mhIxLLXHJDoUAVNASiru4UvZv/hHfQ/58T2gy3Imrv0dIwInHO1rack58FvIM4Ug
NEuVCiM4M3sfnuTUjaEEmbAMInau0vrL5QiI40hKMFGik/9WsxD0pgfYP9hOkjHO
rGbgblBt/evQ/+9uHsuDWaoYUdSVYl4+kBukgidgzwoLSN5brAElgIt/WgKXNQVu
f1ex92s1WMlYGsGEZlnFdW5m0kku4HJoGIuWAQi8xv9FPFpM+6rEiC9kHhv0CZ3v
xs/VSrbiSvHaO+P5B8BomqAHKhpHjUVZAyeEKoXvw/foiarQAOEgXYE9dLojzKwa
10ZoQyR+LaFGUnh+iOIqdPeI3cDrf8jlpBadjahgxV04EYiSWfz/O5CdEkxHlmJ/
m9iNONP8RQV5bEhu4U04BHdyPvTXJoxffUBHB3uvYwwBpbEBQHV4Yj8ICOwt1E+p
gSPdInafiZR6Cl6ddfrLrgZCvJ0rn6JrWgGL/fKOCxR7KdcwMwjFuuNje4/v0rbc
UWICzeuk3r0QcJGGvx/xBdxS+g3ryYFOLCgOVXnRC/tqJRf7XaBe8SQQIgr9GURB
0k45562+bZSa/nkzghbPpenukh/cGHkknSwnH/EUgUoAb21ypKsHua6MBWwz0t2V
r+MkxPrCgn2VPr58snlCeK5UGtrPytO+FZ7cI6ewsIi3e9lN5CuCo0t49XuI+D/3
RG9KWf+7YlEbXNO7lhL/Idd/w33ev0Q8HvhR+A+m3fo0XX65F+EIjZF3pEloMVUJ
O/cVEZQsRMUlmp7fDsY9gnPrcggeiYhp5lbLGMsEMxnHsEQexPgCHZsDJw3U0Tvm
svd7qUEMGYeiT4/d2GgLbLD7hQjyIdm3ik5Tjg5pqoe7UQMXlAuBq3LB+OmiYkfm
ecLKi1vgbI6eo1dVUAmILL0kTTfHesgbxY7gAM12rhS1dNXHOXNgUkVSGytRM69U
VSTVXl9bN5YkaUbyjE4MOBAvU5AZfOtN3cNQSpHKdg5CoPqUHFfeUcaXsrAau/Sf
nxqMyodiySlYaDOuHDMG3p8v0ZuHraGgCjZgvMfnmCdUU4sagNMRWSM9B6FdQsKN
/DRcw+edWulLa7KwgAgmovg4WCUxioVcH+zLi8xEskBAsrEnK6+r4HNNEzedcpF2
Etv29KxXqHGu5POR41joalfg6YMIjPegyTgoXqWxb4Cj+Gpj+RqDlVcBy4c0ms06
T6058cCu8S2pD1yrDQmUOV+VmvxVKuyM3v8+KqRJqpxtgwBVNCBzX7SwqMiEL+nT
LbQNmBFbdpGmts881assoWUz4CqXqmeh1i4wf2O8Pueq0jeNj3h2a2qml30pnfal
zLzLXVlqHMhqwonMFLpQZ+gl0dm7QaSAdSpHmK1xE1E8i2O05eKn7Zx8wwbU7zri
FCC8dA6AVa1vw4H0Czvh5wVPLtWOgadkmdw3q2bRxG2Bx/Xhda1quFTFiJXsaGdU
lrZOPfN9DQqjJSLzDlvOV98u0U+GZyoqCbJLqhCnppb4UcLADtA8S/FhI92lasSU
Ei7AiF9XvTQ4xmOAdfVCWjphY6WtADEQMiZ3V/uqbgxsmUot4zzp/i/FV/arfLYC
W7544kzZXNh0Pan0mb0csptHQuOZ2HlYnkOLQ+ZUvlqYI+SizjZnCTR7itr7Tb+u
R7DTlOoPJmJMxCaMRlPXERfX4LkJg91RM+ddqzMoaOCnJZWUJ/EoT+K6aYNFl/Zi
kai+z17VIU+aYdr5FeSUH/isEnrMQAWjdRNtVd03lhkGlW8hVq8EyVV4QhpfmjR7
m+5p46fwQhPDA/2SY8259aKKyVAcF1/MIIvNJvG+QidcSrnoBY0rVEhmAzUwKs4O
DoTxDSlSIF5+7VvTz3ANBX/JnGKA/p9F6qwp0NSkJiiZ9z4jEcYRSPfToarm/bNo
13etnGcryHgKJrEoWXKCxTDDtU2fz3G6b68PEr53pRqbTP5Dd3vs14eLx3eFt8Uq
xUiFYzPFq04/e9xNGc79Nl5HZHbrtNxYISkgQYInvES/oKSxcfiR0JqWzjoCyFIt
KKdtx/JR+vyCTuHRv1sfmXIGaEolW+OjtFqXnk7de81DbxfpZAgLvArAB49tojh/
kyBImkftKFH1rVFzyjzO1HYwTRLlrfoZAFtFt7Ukg0rzgABkaeokzZmQ7vgIZtPn
NLvyo8mupAjXTk/s+lKOtpFju9jrv9yx3PyO1ZrYTylCBOZVpLU4NAZOHb1ahqLn
+l3LeHXh8+UEB64XrRt/1zPmZbLueeH3wBeusnxEBIJAD02Qb0Mil8e94i5gqcXG
E1ksdhVrBdMMnOgzWxb1bTbpodpwOoctfVXmibjl7PpWaJPEyo4wbzhqcW89LZCC
xDNxE6QO4ccc7j7GAiMMz2XPTS2SUFzu9kDG550DZXUmrzQnsL2bEnvzkmYqMHHG
7moIxVAPzz8CufG0ZerCxLrOVF99zxgyWotW3JSx3eYc87mcEBG6M2YrGMZ+cu+o
DCTTZYtylquu1Skbxi6045NujUWQIR7/6stqFPIiQLU0FYoRcyaHKh9H/XGFVa0u
KT6bqjyixLlMPbm7+oo5TtYmKgCWv157+QuAQ/6w6bUd8qI4/yMGuqStgj4f7OHK
5KLkBUz7baDimzGStp9Kp48PF3uE7ilou4lBdrafMCd+/1tIMG7EW2HS3H4PA9uQ
8B3mIOwviZbaO79ShpevPNaupBUnJQbLoqKWlvKGXWfXZ7ieCDy+Ne3CTnZhqapO
ND2sXac9TX26+f6NHfNovBMPekJmas2Ai5Zb+7ymTSQije9gJH9Hb4E7Q+mBqKZE
em/yV7Uc023CtfvnI6xFhpTjFwLhOOeEkp+fM2ir3iZzPcdd1AcVQE/L4BdgqT5q
Igp42FpGOzkh9bjWsVzCQa9/E5CGSDplFZBsdd5Ai4UivwdX07T/RsbYOCQAbKLp
mFYJannFQGdkcO1n9d0omfuP942eFpe0XT0anCNjUQLHHosC8dN6hU6CxmYUTsOs
YmMznpFI/aJaEkqzeFdsmql7E20PZl9Wowy3U4RiHKRFjt6Rsft/Q0XjBICd2iYw
buR/ohcTdm1s539H70cYaBlyCWuFlxl8OoCP8sc+vDsNJEnb/Y73bmxGqjrfzzQK
+4ge/uBRotgiyJD2DwEnSegpPMCqTZvgaQ3uNNL5zHJaUewqgEmqWHEutimAOsFX
JRQZyZ2xQ/Ccu1STdx9cG7493Agqp9AsxWexW2i7wZKYyCLARUcEwBKedFjagXws
lCp7ubxagpMBQ/QT9Me9s76E5hTc8QIZ//T0NPU+8yiDj7DIfIfijYOQ5TAT7qVV
QT5uGMBGTF9k8QDMLeDpmKTvTU21jj9BdcZz9MQvNmEvIfAx1+0qy0CvwcSPWQyY
qCtv1zbws/pNwMF2UsWbtDlRCeHr1mhDfUY9XEhb1EzXmt0c/eO1svEBmw6EEL3i
8bJyu7okwgCiQm4GXv7elA/gUtFlLlrpxPtgRFsBpwP8ec3qtwuitJgU9yFJ5PEu
ld0HnN8d4J3fitfmvnFohPclrNxosy0gotXwGGpqNy8hvxeJCMTLBy5hBq/dFjij
vvJWxYUcLp2pRa1c+6CSLK4BMrGINbdtkFCMTwMz/IBjyT/QhHibvPPOxj/5o0a0
qY7VvvnWHnF+tCT2DacjAlcyZAj4ysp3ftUw/RDkc6GDs5j0hzkNLZyTmrQawKLu
QtzLrSRJ5W9YCDb+8C+ZBLQKPmxDraksc0OQs+s5mHO0Np8VcI6/iuKL3kxFKBk3
P45pbObgw+J3VdGF1qKRnRAECtW4JkeHvyhuhMil8NuDID2VuIvjQPxABxNyvO/+
MlL5JsgRFHl9horMR57SM1UuOBZf42liCKvA3imF11J9vwmxQ1lkxt0ES1Vl5FWu
3+2L9r1dDPxhoM6I8lmEuzvO+SmYCjEz5POw++oJpHgoWg3O8xD4tpP5fJrPYG3+
mCa8c1N47d1+eat2Fsy56jwJFCe+XwgV2HoPcjybuyXmlsTO0cYbdrL8LYF60sRw
fSstrOKVPNnPJQaQsR5ErMlm2dmhn9sUhbf0HoJ0BZ7Qr9G5/7humrPJdisrsGJ/
Sz0LL3I46Pvdc2ePxQ/RIK0id7ELuUWBxIUFNKPbbVhu4ZcNE7HPyWf+adFDROBj
q1O78Nqop0yMGCB+FF18pFH22ytCsHgLEJbfnG96Um1JBDR6By8pgWfxj9cNeM3g
isb1FT+Hv5ncrbst8jAkmkgd3zdG5gzaL9kJ2A2k4ffvbkKNYXGICRHG+eewdbDF
omxKs5UtPpc0MIysXrbYC/KAjyjQD1bv2QtPwLSUhVgWhNAGalT2RSNTT3lqnYfy
cKhO/ROYDc+e6gxIqvizOvcOu4TRMYGXBP9qeYF9sCkxwcSu6C4DwGsagxIuSPhx
Ojzml5hlGUX5sUVMFmyFODNER/oxkIsQDV5T8PB2Py5vw2lYJZMGUG1aFT18aNU/
ZWJaU4AJyptqsL5vKRD3crgMGrwFFHsXbIEqme+hLbSYUuOrGgwOhY8MJrapU3ZM
2or0CSi76hS8Y01aXWUNlXx8c6+8nNIfvL3R+sev1+HzeCD+LoYADdL50RsiMVJs
mRZCClvecybOVpnR0xFrsQer1KHPrWjp3xwhvkLhOjylnAf/926kzdNtSzZT6b16
R74xIFSC1T0kbdXlTgoaHAEXMTObrxjSU7qCiqDj9mV7j+2dS73hOsYpzrJ6XdFg
lwv+2IGtvDgeZTcyomXNy7J1/s2q5MLr3ixDBq+nvIMq4eu5L1XidfYTbVb4bc4I
1sI+kKNEqOAGYyQLBcvCu9D8MepMii9TY12qd2IOVa2qf1BjaMnMr1ZkAM9pdW4J
0ffz+pDiaak2piyag6XIzB+ekT9+B0LW7v6qHhWtqu0IWXyAv5bWs3tq5B5JATFd
eSYpAm6TrhAW/9l0Qg3MpbOvm65KOrISPcU8+cwwK3H5lSMeKzqyjOd2RcCB6hRS
HbFNrht3TtzZsMZ6Lk79IKqbyK64NVhyEDL+xpXMY/NXsVuPwG+QZluLY/4a5y6I
4Cb5DVAH1g2kD3mMRIXiD4VHfiqW7M1pyv7jA+2FmGtGa/EgXIyyFelA3/eN23V3
6ydKYGtXDrxjmAD1eAqTH311JvxnJCrYUA6Mpup7OGnat8FcUwuCrBW8Yh3VQKhP
xT8jqMOiIki31a6eCIeym2V0AsQVOOJ/ythdYOefZ+Xtvmmd3/vTE1vYWYVe5CNZ
R/3+zpIJgIsOprkZvX6IoQfAEiYFS6ennhr6kG8FutNNk5OHcinir07xa0CfBSBh
y+cfWGbsd0sE9aCj/DczRU5+5fkuHP/C/SlAXBVyMS99V9mVjngetUjU3PL4vbnv
h9iyfj2hMwJceb7S7IALTiMSgKGU/Nthy6LQ2Nhi8YjrIn8qnRJCWEH+szMN/5bi
XzEa9iiu+WAQhZO2IzKFXDzwGw/ICcqHL5/vYFMM+6oKm0Q9wP967pqv0M6nX/VM
SwosjqZhdtxQK3nZxsMUgNsP7nvbiGxXfJTxIF7B6YKg6BIKnpcvLqepDRUf6zdB
Da1NuRWS5zrlv2ADvtQHz7bHM6kNlt0YNHPw4jEI66xcKghuF0mFyaUouACQRwHd
U22NJUVR8rFPn+KAAorcvQ/YXI02q8H2sLUE8mR2Q1k+8VlkJyoEp8U8JGndTyDD
ROX4zHb44zoDdEUYm+qB07mRgkYKp9e+N1i11TM1x+VUT6qT/THBKI15fWteYm3z
lxN9NqjjRbBzkmyeq06BK8JbFDGRyhvfU2qy15WUjucuPmrsEg8cpUym4Rk2glkM
yj6ie/EqYIMDNDA6ZHzHZIPW+/RsNAQyBblCNv3aWT/ShJLXwkgqt3g4ZaMnq5Sz
/r8OlvvluMKqhzyHWUkW9B7pT2ZZXYPZlqAdTY+9YZGtMrajqvYqrNE3hkLT7YcO
q5s+IR5a9+TKLjqGom0bsZjYKmLxdQ0Rqmtb6j8oSIxHvYyImBtSjWCvx3Qs52YE
iY+6pcJlB0ZTTcvyY4FcCDCSJrDBTiW9mpwNMjPC94W75h13nNqpcBDd2ujnb87E
aZC40KXa5RuPz3b5scaJyvDeBYHefwcs/6y1e0MAmn/tvsMBjmuhNgMXnw8jPLOS
l4+2MHRhbqJ7IdUKW9OB5L3vjumqBIpMH21aF4htAi58yKRCbjTY5++FCU5sbSQD
/Wo+qZKtkNVXiBxJRg6CHQd6I76JfMVAVh0He1WaqwQ2xf1K987avQecuKmRvLyz
Ns1ajkwAv4oxraP9o39vzFZwBmNJ2YU5GBHCvo0VHhjh6mgjG+EQPBgKzCtyVwPC
JLMFgjtQPHhqPumkcS6E+RoN9iW7uk3B+EWYCcnYAU69L2QiGKRpyaGmtlv0F2lN
HkeXOv1CPFwi6DMLvdv5D9Lxwajj9zmkipBTMhXWxKKnbpx3QF9SvBaTPUZ/QvEf
unjSNZZDWG0KsO2s6/t7fnpF/qJ4ALs/uTH6sqW7Hzx1c6VTFuuQMAiDhxobgZ3k
SKw13zMR90pJiFf4xx7XW4tVxgOr3O/0WoD5bDVlOwQagOI2BqnQ+3b9oM8wqSk1
wbMYuC9kk77UwNUA2kyHhBcmVjBcZFi2ghVDAjidtW8yS6A8OhQyvLA2uxUVZzuh
aX2oJtmVM3MU4kiaYmnBq9uFutMVSdwBmYhBIXDBNSaxZNM4SHitnhtFOaKkUG/J
isaUqoHKlLjt5mGgud5QZwWkB7OlUzFl0ss9i3nq8suJPUPZzd4rPqAqB1S/oFWX
r5AwhXeRZbsvR9LGH9dscgryXxndLOUbum2MXz/xyNAlgsRU/6QpDhAo0GeNATcg
OOA2O9DTHCDF0tz2+JmzT/ahgZiuSSVi3u6bm8CeOc9+Lq0pyd7oKda2pqIedbEx
2Q4eof+mTNcJGOMw9PDmNE+cZBM86FPzKu0NDVrBcEVtAGlQsiWKFXUX85/fJVmd
8K1RgCwh7GqNFsA0Vs10CKrKDtDlDUNq3/RE8Z9sRRhsgnlJ9wgjIpbUA1ZTNgcR
8e6y8qMjihwFw+ljfDkENsOBnqFTCq+vWwiiL6VhrwoVe0YctK88z3mZX3Nm2My6
LbW7wWUbsUWrQkcifWqrEaFIfj299RHcGiOaRqiSPshosLa6O0zWyVqVjdGk0Uwj
IhGrjN+j5dX1oLCcqGpg7XvgxyZ0U1NRZk+oMmeDlB8MgruCPkLMDDZlhJgUwNwQ
t8TCIuyF2jb4xOLzqkHeRow34unJtb7ydFKZxE70Q2pUWstn+GK7zlR5A7N999gw
X9kV6fqsqOPfDttf/v9RqFIRZIh7vA2IVFDovoJYYzt/dE8vYD26dEtQjCY80Z2s
8lu7S+W1ezWstho21ECWh3+gPNUOyRvr7PSathqgoa5ETiwqu9hw50ISlQoRwrXe
fHcq6uNahWPDMsZ6Z5S43bMHyWsqwGqB+AHDxpxYZWYz5b+mRCQvW5V/eUk8pAxn
ElL5T1//rKQyE3PkIHxRem8tR0UyFUMIZ4k2zzwu0zc9g+SpgooWqE4hz6TA6L2J
5r0P+KokkKhjiApwdg+Z4K6fwJHIpdLr6sBCA2VROdCv3+pSvKAuM4UjZxkik6J3
OonkUHbsTRYuOx7ySqaMthWR9o8eeEqklVvIj9BejV3bhEwamzZnCxPI54VsJf3N
qoTnvwVGsncIXsqpkR3KbtU6M9ChxDrwWey7E8xesMlCUdVPzSh2L2xsDfjWp/OU
JNhqmuUSYAqVZmHnS+mg15EeG/Umv4DXbJZWIIElwWTTwbvKofAFlQ8qVe/4sWf3
fFqAIiEycHNswdhHo30ZFpJEp/IeuoorOJDg7aHIK0Hr3Xt1IYHjRsLCkENXtXQm
pv4NlV6LHZY9tTA7vQsNDmJSpPE9apokqN6bVKZ/nDijfQR4IobIs7De4RAZqGiE
Jyqjc3kFvXszQxpArFAEezpwX/N8NBxwS48jrZA3QnlXVNFF9YpTaWvjjd6v+lCf
QFXM/j6YDjBGvAjfW8GIR5GeZPlBnbrSn3+m9kmAHENUmrykab43RFoY18Q/sdyu
OyIuzmQemNVk16+Y8/DcCMLEhtPTNWRynPeQvbWyCXANiO24gzfR2NS5ONP5oNoZ
UflF41kHnZ/aMODbyBbiLV4YNYAle3W8LqAixlGJ8gnJoCx1smQD+e23JbmuHKIu
JxnHwDCdcImLG1fCVQ43Ekigq+KgWYhBbPvqXvs+4xTIUG4nEn5DS6o0lA0TTdOM
WcVeCIioqgQpgaahP1T/AYH9EVDo61rvg/QQPUixxInIixIGwsKNZridFmHn4q6c
LjzlY80kyC0l/q9xKBtByRepsAWWkyKWQ8schre/1KqlvhKNEtcNbIeAasJ3SbcK
2Ub8EEQQDIQNfo+mJcqtII/d3ris820EKlrFPE0Z/7+wvePXgItIyJFPjrs6b/5I
16Nr7AqEOuucnVoWr5xtRZ0lgwP+bN/2OpadObxTYdvkugw0niDmw/DHsRjQAHbt
yssrmg/YMs8XM+gUP5R9tEWb5972slgVeQGe1RpiKMZmYOM8DSzbuIzeotuen2Gy
Ez8rf0YygG5rFIqRTdJGK83wWkQz/kPToxDPtKhjSwJRKlPgcPGZ3dHj9aMsICi7
lCfWiM5xTD8hasPmF/1EtMtUBkcsokkc/V2Prp0pB9frXyPZKrYsb2xJ79oksJ5Y
YXCKt6jm/4AFADHuNOgVhEoU8oMIbZC8ABkPGN6u/MrLrMtmND+CnSUaih3iGoQv
R8VK09nqsXCuShMVU4PdwiraJ8QuTggaCTJbdWaP/VEzdYg5YkooJ9qLaaU0kY/i
xF/dAUCUees+nJk/0jDUfKp09yvTUuctEvWCqsPzET9DmJ2qnQzxZr3l/wO2skrU
Emvwss/OVFw29nPtNHt5N7UPLBoaPdoJ+kqJzePXhp3KIlRH13UxM4gEm4xEjxwG
rly4Huzc8r+hVF9Hl1ygFgkb9CByjD+bhXkN/FURALYhFxnNNiMstjNRcbTBI4q4
QmMnot12jvGi72OTmN5bR0T66H87WgwWdr77bPVGsg8tJVcswms+UcLSduYJ/+f8
tT/6qsDCdiSU1NjM4MGnAmQbq3PlFg4v9Y/FyRJcMQ3WPjKPtiyxngd41VrfzXuR
oDPmt9ykQTYmBWUGvktvXA/w2U2cHhCgNgUyaiCndsv4J7IBoOnKfvqzd2WCvEcS
63usW3OseWUKPYvKnnUSXWoNT0yHT9ePqwZkn46ISw574SaFCbg++oHMpsO8pnwu
LyxDvxVT/CagfNoQfXrThVd6UsK6gnGq8bM+gLEdcFrDKsquJsF3BSUkLz8Ph1X0
taznkMtQG/oA7gUZXuRY+j7+vb2lzzde34E2sslqWQ0oy61c5aoAhZPZvFiRdSw4
+SfuV/v+bC57A6btw/1A/gedRMNPoeDhp0HLyV0nY4U5YnuooneTY93tzCPHJBfu
ETN4q1BJ/PE545yAKsVBi4xP7ozWGXZUc+OjTm82iHvPnrv4t5cpnJlnQp9S5HXQ
5hzfJvKuXM7XNo9nRkz6R1fmeoJWiDi6oqXQPlgfxbnML6WEmtparBEPcqdO3lBt
4ELbg7ffy1Sx7gSvPZZKAlguCWOjB3JmdPAq2asw6tNWaawsbiUQBvOitOungpS7
QQmCjsyJC8sUgnNM1BmabmdVAKNzQ0ohR/HWCf3HSdtttE2Rwe1cEJw2Fm0P5B4I
5Nr7wtrW4LM2yGMsTDoM+VifH0w7uKrzJjQyyt5t/X+4xe0SaHbg3i/1tOjZEO8l
pS93xnlQBp6WotofbRNb3Tfdj33jJAGizEVNUp154MV3On1G/vH2L79sDaGnEScB
vX2TUEWmQNxBHGR5dwtHV6YfSCrRAI7IJpykTqXSw05KI/YjASvQLQMzxImFBer2
ywwWn+YXWgKy/DbTpBftqMp2uGXRCKYulDGQ6RpMSoMeBPVqqM2X22m4PO89DmE3
LVPyKzyaRszWtXRmvsZRdqEQxLdMfcRvx3Ly5Sz0C4j8wGgLiVfroYLW1PJiDRpH
hEuzdPVqF2PTC/0Aurd7d8Xw+S33nkJAGDmX0RN12abHq6rLdnk078qnQk6jiXYO
9Fy7cJinzopSF1eNVu9Y408kQbsJ30TIlEmRIABzzwSy5Izp95oqSbC9f4eeleYV
vHWn/8puvSGvXW3M70umEPqjNyShbMtXvt3Tgvc3sY1lupHv6InD/IkOrwN9Syb9
KFG8Ne2GFbRbx+DDMV3aStkTjVsXqVTNMcvG/2BqRDlWLIV2/8WqSL8d4zyga/o3
Riqw30PV/H/kOR+VAApOT9hR9EOTNUpC+t+2Tky7r8r/IyicXBRGV7KNTn9LJwai
1pGeEd2eGQhHlY5bPap5NLTCZE7TJ/noPH726iR1o1xqluqA0S7vYxUQT+K2h96y
Brc6hj3eqwUQbpbIe8/uPt/lO9lkKE/wdg47/iQknmqNeM/FUJ2JW4regqnN+Hwg
cpb368t3J4G4HCTrfYhhKQI93cD+yJtoKsx5ZNAY3+SkV69lyT7UD8z82sMbiXkt
q695FPB2pCfesU3AHI5ioLkGbjy2ms4qi/F3B9XnePNftVI6yhE62wL7oFE2RcLb
NNyRac+30wSG9jo/wA+sthRrmkb7jdCVFbZKNHWOWFil6Yu53Do7mhNtKLXSRZQe
gwOunvIK3K0c+2DQWJOkr9ZKwRUJU3dNBI3ZjxXi71BAlRbtqR4tz75rtZz7GGLD
khBS0J+dZx/kADdTzcgeCMpZ6eNF5H2qXcy8nInTx70zt8ilFGJHpAmYq4wLdW7W
2GHdoVzy5JbWC2lawo52eEQ0xWe1lz9LiTMgBbfNK1/jPTvVLRN34C6DQPMZbdjU
3ovcql1SYiBjUXQUFChNdMd/ql8+s3ch+RW0Y+TWKNIgcSUgWOwMVEz7NiCvw8Ov
GSI4biiEBpNVEQTQYdcAQKkhJkuzP6zESSzEvr6s7eIQ6i9vTnZDLn9Cx1KeEz9a
1Dh3Kogj2sQGgCWvekAbSbB0iX5OZh6QcPgIvr36Pmz8vyVH9h+XLBN6FXy5k9u6
XwSrNmhyjYtr1pTAkBs2enKskEw19T8WeWO4YLr7f0BKxmMvVcFv+bxn/2QKtowT
UmR82tCmIewGw19EdzHgnzkYWDchUtDD3rtIXfY1kckmc53s5/5ZC/fdiXKETS7L
/UNtk6QTl/QTHpk+tA1fhsHyH0zOG213h+JnjjcmTXHoGAA+85OuN3/Bh/GGgnMs
9LhqrOg69wPP1qehVUjD9YZIp+bi4NuQUbQC1MmSNLS83pHbaAwgmjLcLH8b99J+
smaf8yaJnDtF4PlPnBbHNwf0sY3BxYgZA9kLavm7uZfW7Z3pyPZg6bcDG3bLYx9I
QfrK9+M+/dN4P7NoDT8/s/giDchksVk/gmGvSrtx7G+4gkyseepGQCXOmozz56o3
S65YMBnswYZy/NaguRUiMgej9D/XoLYFGTuyRlPafe+Fdfdo2dTxNxkzicJYnB66
6sUuOB9+9CwfdJYpWFvWlTZmcfmpEQT+BXIQFdh1XjOyvXr0Pi+M8UzqqASsPZLE
J/BQhqjL2ix8GMR0X7a68/zBjLmxMdXg3iuotnrjmN2wUujPgf/lmf2koL4c/V2h
I0t407/xwdR4izW+Otg4lW0I0b/nUkJuSLdISa9A/5Jyt40RrYnr0RDR0wQIE1CO
8l+2gO/6+oLXOYD1LlX2ZiGXqlleEnftGFTLIuNzSO4xyZm+BuBxsM498T+68a47
nsQYs9DjicdExdrRJeckr97C2woz2zFNR4KlopyXFr8oVDhPzfSTFAB/o0JV7fyi
J0oZmiS6AqsOCUfh9RJNJk95pYQAjo+IAMyAGE1f/LIYOg/9Wgz3K2ga0NFqqlPp
dF8C/0dkhZ5akpSenSd1AVZSnSyNpPjw+J32pLZLEmwVxHn4mg4Fu9cdx5g1/4dR
B4USPDyIzE9L8XcWFsq1Kv8GI7VdfMt4X81ep6e4dFVaRK6IRsdHywcTSJUJ3WiW
sOo07xybyVvRQcD3Url7PKsZGnCBw7hxC35SRLKJs1LRKIohVsC9Ez6y/yz0tFi5
QIhk7JBBMRjxyd202S2sm/5bLw9Qa36VF3vrIqDohXLyvhO4PJJADhD86FFHKoar
Z08LBQ/krbuAjfWWQv4nkjuSePWza6RLAhBKwcLsQSFSoDYeynJ4g/Jn1KCJBIAc
knQYfvQuQvudajWpn65VQTHKhbaG7Tl0vuBp0mJ1kAbobnWLRctNNTkDztrWXgzJ
+YZ+84ktwRxYXmanezEzM34I7zQo0IF+0XAU6ADN8uiZ7iARSJODQaalWytMfkJG
8hKdNUPjbJeM6nUw7KmfCossrUOf5WkpKuytv//Nr9hO886LBDAHyWHxBoZ+xmF2
MVxmR34Ez4UJSEYfu7P39m4vssXi0bskNU4GsjemqylrMQ/AoJ+lkfAgSZGtqYZk
DaoxL8Ibw4xRodifQdXjoSLHCqc1aBDQPTAi2cmo/BKjI4RoomQ26X81hig1Svrl
6iq1KetDvnh35OuBOrY6PG2hxtonoZxTs0Hn5qMe6AB09DNVZj7OWXoGdT189xkV
KGCH6QXNjgv8MkcCtUZtCt79wJs8npYW49f5no8Z4aHmXX5Huq6qFvExslshmu6L
t+PgFjOtGqaWY1d3QALHI89HRChXe5H0vxMmeoxCUWM/EDjFm2Yr4rk56fPsOArz
Dy4pzATj7c6Tc33tUiZxYmkLVgduJvPGVwU0b9h/c8B8v1nzGfbDQCRufVpCv3iZ
3hKhaj4662p7jaZWGGMb7RR9rlixOiAdueHsAXV/YQaSjl0X0/nDl+lNE7CFHU4j
/cvjmtI+dQZYkHIGXG275g5LFMty+2GzQxd2BXWUP71Vo0qOosO0pgXR6z3c4W3z
4ROsapDqPLh7t/Yf1BWom1L3B/tKX5nmVU6vG8x84aMIjx3tkHC6+/MUi+0Xn+NM
Z+SnH6kCdGpC6uzEriH7PNHOuZLS1oJC/q9UZ+uX2INQeh3JbyY6aAyS3iV8vWa4
BwvosYw+9pLBkuZ1JPLf1UpKohB6BNfUWE68M1g8UmKMFviVPF9V3zSInu9R2Ssb
BIVXx5JbYDz0cYa1/umHKleQyZMCSwr5MOO6WvKksi9wUSODe2tL4vvMoSFAQ+oY
7O1DFkio0RBRZ6G6022Ks2iFVyzloL7e0rbcW058GVVSeBx9N/1aouEiC18R/p3a
Ls0OT7mOpIuHnNRHVvBpd0TkqazziPRU9xsEOaCqqOXPy3wUg2V9QbW7t5u9r7d4
OH0riz/olZCvfKj4zLDotrANHkTH8ww6034241bgxCnG2Y0/RyLo6o80jz+pxSbX
mHrhyXm0bRLSRs7c8rxfUR6r6iU+B5RosANE3xRMWX4CrCZZKQZqlBMEAAfxpYJQ
As0D3lU3Q6/2hR7tMR+USGt0kMJM0WDDKDmV/PHNm7ut0pgyVkbFMnp0CuiQ5whq
ORFOy5UjjaPjzYLv/KDgG4imXrGvIP/2oCZoEJBcI8c+oHuNEELoqrntGlkKAxYf
xxB8sEnwlyV6BW0ezx1xB06PVdnHkQXS8paN2YYleag+CvzSMSbg5udVEg3Ki7mv
Sm1N5mCeROJjGAFf5k3JZ3my910wkux+nPBXbKwWOaYhAcu1SEjY50yDkhglH8NF
lTJx9syTOJQOVv2s23UMtf5oNqR+pqHhKWul0nz93OGq9TeRqNYRrEb+jc1jpCQk
KAU+VvsFPEEwwOPMqf0scShzmHmbowHaaOkGmuXyVRnqAJUGJT3tR2EpgZMlaklK
FVfujzqXaHuJ+/PFK+WE8fOnlP6sisEZiOyordrChFP83SZf3pKSZ+JkmBn9sP9i
ELV3eUKYDCuT4G8f+lFRRXHzfaCvBVNyqX6WrsMy1gjClGiqHBS0r4kxPQkj5bW8
i0p0OeFLbmteiunqjRICd1vOcRK3K/wcjfilGVPSJs+hvdFjfOeMNjKbWnpZ2tgT
SwKZTcQxRuKfHCKxXJ8IYQADexan6FKeXxosib7Yxw52wWcRX5IYsdRXVknEiSOe
0EpF9gZ9Qy0SySCx9A01oU7AjmuvC2KucKQ5PPpTch2k/KIi5N32G8TBx9PE8Ss7
XDeur0TXQsKeQoJyvYdV8P81xu5uf3TktBIPEUm2zQIP7WVRypMeSJMRNYm9DWoU
j4nIgBkURYiCNRNLFw1k/R1/r2FlcCwgV3DdtKMiJ+GL8dRsU6reTFVlrwuFt/Vj
ijUyyb04NszTWTYJd5ZPlLcsxBCs3o/vD5bpwGDZn2EvQRWSEKBuesuamr1Na58t
J/l6QB1uDifV1b5JdJkSziLdQSBG6aVqiOzWJR4Ps7W1KcRp8uT0q+VY1+h1GNDJ
hWx3z85cctbYc+dR/kobkdQzhRflYn1v/opljw90tZ4F5WgShE+wHsNXfSrvYqVq
PCarGSKvWNpGhbTsfirAhEL8m2tcqvoxf19rt/Pl3U01pU7YwlTxeWmSLglGtD5Y
1guKf5GCy5OJ8qX59IdxTxd5oW7sUJ1WnJC/BcKAM3k0/CTXZHkYjb1VnasT1to/
eVzKmxhvXTMYtyWBhxuO8uz5MpXXg+0Xc2vr4fA866x/iSKskugiemO/q0eJ1Yfw
sxNRPreo4o1X2TQIaCyNSUXs6CipSCclukNNgJanG1fdLDazQwkbA3tLMxBht88q
fWhksWxajigM0RgCe8kRquqrT0lCr+0hVnlpWpuX37HNCMz98iqpubbRJ7ALGMOV
qPwUE4Lks9q7vlp+Lxjrv3ugV8wdfaATFF1p05y23X9n+B+qw8DVWswwI0PJLOs+
andNCTMtl09qB2tJm34QoHm861zCW6yh8DkBwOnc22UnVPlMSTYPeiUhKrBbP82+
ZMCZZ7WF4kWrlFFwNYyygZoyONW/6n9WCkFQ+YywakQJiUTGO46oHRleyG1FS+wW
ELKyXqZkgukFNqJwxmYdkRgefyR/4vLrnplbmmQj03RUEEXtEU+XYpo2UE0KA5gV
YVegE8ZjnlY7LpMd8AgHHjxSMmuvTPelDuL5GwePmTQ2hC0FVGz9Wu1DPx8ihnr2
HGTFSeb/zG5OErCujhOtnixjPYfubVlvlEuz3vpyi4UVDcFweCYqGUxopFEzQP2H
wR8sDZhR07tnJxSq3WAttkDXeZ/S3++DMZVzGlTN0PvwpEFf+J+25zigt0NSwOeS
VvXH2CuxQK4Uf8JNIlbleFo50DDv2leKFDIkBNquCYzMdqDAwrjMnG4ZC/SqGYMc
9RURz9tDGKtY/UK1a8LWK5DWxANvAOJ/RxGt/62efx5WXczXFHfccyz9GgTeqGO8
qboHFPBLLcKIowiETsh5IGKbxMgy48ZGZ6fg7SgHcq5eXxRSMCqKggr8njsu5Pxx
uaiaDoTbGl0z/Yl4dCfwJWzMMj4m5OYCBuCwW2wJdABHHYkwJ1FOMIHcN2GA9i2m
zE9E+mmf7n4gWN4uvQDyND12ZcWBPuVbSmiG92ulHLfC7EK7dOk21tV8BXVVjmeS
qydc9q+LRd/kk0LtSx5A59HV4cUVADQY7cpDghLH8ijpR6PT+KZBS3OAIpsu92oS
XkfVfvCHLYL79Bxldq5A3xi/56MDBucB41sFYVJWgU/pkbVqIu02aeercI665gzO
ZotL/YflyaQcP5mUTukGhbwDJpshC8D9bIXtIonh3N/6kNMvi4i/bC41lg/Wofyc
/FSQiRfmbf1ad1nPNS9An0zaMQItT2Aah0lvY7yW4j8ff6jO+cYYIS6cmChVlWqi
ejlTIppiT2mVievmn+2B7IEQTmH0qaGt8UnKDows1b3ncdv/PMySUp7oa7RP0AMd
7dxCX/GupSm34K0iDKgYlAeXUQMClOOqEKZPIjUvw6Ws1B3h0FnhZWpQ7tJuw2d4
Kb7l7MeTmhnatCxeVDtAs9olpF1Dgit5dKnkHqh+o53zRK08cBuahnXwB9LIq6OQ
H5z+6SYG2DkfaY5l+DeRNTfhndY6Od8jonAhK+RkXzcu+Na6Wf0BZdg5Ne3wVhAp
zqWOQJwHyegmopyhTlF0paIg3qYKokEWTxiDCxtW9hOshxnESyR60j6+/V+hKkT+
mc9g4z7ZWHoU4ZN1R9WbXpwYFouet5WDFEMptbJz1u71hYaL+vT1KlW9vsTeWaLd
fhQwn3KXJe1OxYLUdNQ1O4k7Tuec4cSCydJR4i3XeCxOLb7Q0PyHf+JT5/Qvuxnh
qbFcUe22aTFE38VSKlNeIxr3/cliY+jgOyDlJ32WCNnydKdvAJGrkPfhwDUR8xJ1
nsOEDpfx2Rm+iOqOHdlPe3hyHTk39HjsdHq1lcQ1uyPOiXZqPgWemFJEIUJKvDxI
6Vi7W/aLSPB60XJ8/LMEorrtbLXrN4pYLJZmW4r04JwMblP/mNHM0wvT1/E0b6tv
K95S/2NRXdulTZgIBlQu0jcKaUB+tM5rBmRy+ARcaw4XeNtn+ZagKL0B9vITwjKC
bOAvp4N+c7SXIOtL0m+zi/g7hUuXkdQ+45t2R2D5KRiyCwZI/E0Wsz52i3Okc+Pk
AVtVQHvqTfp2IvlkwFN8irt8WG6KfWZ/XkUt2reYjd08kAGx3K5aBLgLnjAPE2Lj
SsUISxUa9xZLzQTv36B6LeR2U9a3TtNwoXIQiROCq4w1UW1GCqmhaCqZm6sMUb7z
Ss7PMZuXweYP+wAPwYVWgR/A8I2Tc0GjoV/FfSOCV7aCUWq0HTsLOL/dEd2yGQpu
JzUpbc04eUsu+6azKPUTgfXq8M9N92Dl5qng2AVP62GfyxXMXXSsMNclNYmjRfCM
IGB1Hyuq27slC8+CAg7Wvpad9WvpVHKu7xV40/8/NkATraF6QsFSGM+iFfTcY9OC
enUd0DVX9icDyGNOkEr1zJN2X85HKZIzG04gVNbmZ3VRFpp4cuHMoNY/OQz0NeyI
3Lx5r+I1f1WPNfclybl0cJ8s465XOoRw7/yKE1J+1Ar6PfgGBC4R2OWJai3uSYaC
F4eQK5l15BDogoWVuiKgS+6blzrJKD5njjQpFtuEZfTBFcvlBbw+qiPhON4JoZ/N
6I8yK+30QetcYQEAXOENs+DHdMS8+lSJd1gEstSHdrt1QeKX5hCyTivvDHJBRa1g
Fg6U2haKW2X2PJaNhMrqFPG4tvVDcLBk6oy1ZGTQ+Lf7z7H2XK6wdCCfxdabxsPF
yEA+6nBte+xGRI0+WXIfzAmfkP4PG8ahDVYWjwEenLBmJntCwX/G0gzutZ+B1emT
TRbzQUt7/3LuWkVQrGPiElyjH+/3ZZ07r1YaIMJD662fTAH9Bxvcb4ElTKMQZ/af
FbOl1ycYYWdmr/Y95dvxhk1yh/+5KTjiIXmUdfaiOlwDOI/xL36dHxnA0GV2pQEd
UC3mZNnMuzkDA7jquIHc4yNYshyrzP76/mk8MtCZNFEZBG5IkTvMwlE2vzJjfcNo
ZQ8y7wjDKz1h4cnU80cRM3ZdC+wrDzotVE1EXAA1eiF5XCwq8dw72hz0w0Syah/b
7lZXI8G9aHB6dg0jdNhwkuWvk6qLr4yMON7brwNpipyE4JBgAPcRC0+abl9qLgep
oARypXkJGPKWyXIIN+OXrljx/KigC+Ld9r5EJ+ZLcpyN9HlIRsUkBGvr+9dlMIgL
mTCip/o9HcPMw7wBIhh4pmXMm5vUrkDYzvhVmElt2wnsmy0Is6InblArzloeNb00
puoRvXv9eOd98Nphozu6ZBZd13XJndfEuBJXDFkfriREXqNDFVQpPZVzDS5bCpac
TK6Aatj/3HoCQ3kzArE8V9V0lcbr3ehOapV/tuyVfgGJK5Xgpgh2TNWux7veLqSf
6j/NGC8JE+8Y0iiSNSOi61S9qJiQ9bKiL7JWmt+5Ho+mFlFkQJ/qvTS1GBjiE+Vq
vSTU5xWceXMNARrsaj+SIzAfBWg6oLMPjuNMRLYNy08U6uZ7OR6FRHGErL5RM8X2
/wHFUekO/+QQiqsslRWaags14Pb6ub2SxOw6X5MbBgJ9CYfL2smLVp19BBpBWVLg
xTlV3etss+XkLaH3Vh/vTLvTAiF8gs074hFUfTo+SeumPHQgdGllV976HikOnoGu
H5uY3cepJbv5qf7BaMdKydaagCmzFFSMk9USB2YC3R9eE7+PHkaLF+NQxU/q2WbQ
sGm/By7L5cCMYAFQDWl4S/6fayJWSIj4tVAny69Zhgs6489e9qjXt4qQgK1xW46C
GMIv3dmfaMXUeI0Nt4uJMzANhh5MIv04sWS1vUQkd8BaCjOQHhIwfNWvVLAFYb//
KwH4Eas5JCa/PssZ2jGhHY0wiDAf6C7d12D2jpXBUu531bTPZB5usqmW1pvUBeg6
obFEU2/lTQFPNnSkJaK4ijh3UIP5/ghZckEU92VoOcHXIUICxeUokw1IFek2gbbG
NyFDtHhw+j5DrrH2CDPGknlP7f03q4BtmvGHrYF3Dv0sThN7B7xOVhGgCjGpEukT
HLOmke92fTreoFogToxz/dbcu7X+64O16J5sJt/pJJ7mG1pjelQf0YuA2P70bk4M
zfbpS+HeIICYXFhi6isHcSBzLydLXQyTECbprQkTqgkE5PPkaewtl5xjrLG2crCc
es0GZahVt7NJvQCeK05Td/WrVkEppsgfQL0OM2esoBZyLhZMDNWQQqP8Jznc3Mpb
FZRa1MvDpmpw6d/iIX0rPkRwlMk0l88iw7kxhnNs7oEBaO0zU5HvyUJGjXZG8075
e+McMfZv6HcKefGzx5lXBqzlDPT4Zwl0bR6LhPxsjynKEAGkNIqPeW73ZUy7hH1e
JXYGCWFKLeFq+JyyR+/uFqJUOZMSHO9XHZQhCmiOTDtwPNvHhEyJv9Tz+/+nnlIV
ekfjdrGQ0OACZomlVXFf+wEGBFMpQnOzSa7wNQhWiGukh5Gc47kRZLdHNM6NB26U
cwKVOjLoYzYnwfkhO4IHvYS2VdAqoMW/4LQhiHvAssY7oNaiIJmL6yLeg+dU0CN1
IUGvMASs9y1HB53oXvgLA8kAD+PKkrIJ5gM9ooMNp7tCo0IaJgTsTz5/9h3i62b8
R0SJ71y9pvgUKQFJ+LxRiX+mlDzV85s0vYMb6Hgr3js8FCjYI+byKQ6QOCjLD7aU
jokR7230862JqkCc1DKUcB2K2ZHJ+I7EG1y8hqeuYuh//h4jF3VpKFFAbHhvPWuv
lODt5OEfQyJ0L3Sgheb9ddt7IQHAHPw0YDFNEj2JMZDHOKoQR/NMXOd1c/7OkbLe
MmpgzFgPNWOIXB5s4OcI9t0/QLPQ1eRp/4iJjcaD8xC5Ita9FS4PA6C0GS4AP3VM
QnQV0xBmMqJYZ+AWvujrNW2hUTT9TygJZy/lgCYQPpUXM5RXRN0C8eYyxZlVPtQW
x4CZswQ+2jN1kirSLl+T5AvOCjZ+Ng8eieU/qfvxAsTSfT7tDNJvysof8kzkCqTk
BmWiBqwH2p4OPNvEqiLftIEluMZZIdiZrtVpYc7G97v8Z4VqmWi/O9tbiwUpQYBa
kBSQu6xWsAV5yE4KK9FCnc4WZPMi0nuiG+YTD6Wy6Hi2Jfnb2L2H22O68vLxPRZf
QbUlQS+qgZK3XDXtMwWtPNlTyZoRo3ChU0n7jDuOyG4wwS5TJlqeiF5joc71jUpM
w8aechIkNCNnnsnF8TKwvPyHbQLvmsIXq/ZLM/K6MS6/cbI7raEi9cQX5jUA6LPa
6ZlHQx1Wy5u3ftJ+W7ZJRhq6pLBXDs2hK8FeyIAbhG3h8O5pQMWJkv5lobw+DLNC
ESU4bqeSfzqatt7Qy74V4ikYZmzs9VPbWcAVatUN1sorFqoXryKRoioTkaq4PmPy
A1j84mbPLKX6BhIBz4Nw5+gQSjKVh9dFgtniQzCxZaC6clY65yHfhMiFhDHEjESE
/HdwkN2yah7Rb6btPLMwUa77ONOhDXrXGJy0FVWjAXWA+CCVeDZVUm+okSPLZhW2
+vyuexbjojZYB3teQY3sBQmGOl+9Qx6ZN4An8K7Q8BF5fbQOG0cu+Z36Swc7DTjG
cTOk6jgcPA0u3SYoJdGESWC9dXXE565z3ZnYUFMWLmEJgir35Orgx87nui2zFHco
XLcGN6q0oTtYLXW+sPFxg11IW2k8dVBnKvOC/w3/1KHukg2R1Na44DQ1JRnwZXFG
glyqLy+wPQT7XlihLK3ZCBsbtOGmUiJpSe88uxjsp3fgUtB3QoJDlEqSTRDedJfN
2u0WU0yGa9KsJXQLurTMBKD1tMt/xz8eGDjvydKM3glKsz0ZknDNqrJK3RCu5Ze6
bhfNuGlQVoycLkhi0TND1+6AfC3OWEuVkLflqpTOowAKOOxNwSbZd37/3zqyM1t5
PtYLoLkM53ZlVMn53DwftwuStEN8APlBZOpsmoEP07HbohMNKeq9c+XTn7YI1Zue
K7stVyaEjwzZXCbQ4YXvBA7gV+mnAjrjJIh+nqre3CNbkx8YJd2dRh9ZKPJw0z2/
nbIoO5tv62orqqFRmRrxKdkCx3RNra2APlREhdsTD83EAvVRJ47ht2j196PKWsc0
j4S7AKOpRHpxOIEWcuoRNwpIbRO/E5B0AlEuEwgH8EZ/wdvP5kd064iKhN8s9+TV
jMywIX8u0vOVEjKmeibUuv8qNZylY3mMHsbZlSWg/LZbaa6Z2xkdssdIjGadm/sY
UBzbATyV4tKc2pxzlqI5hqdYJeGMiOv+iWocE7x2D5DW2eo2BEqpQPn37x/cRZwo
ot2QAnP2vLeioLcMNXHnoKUouIyN862huD8qRxGPUUi1sGuWVlzVI5gGRUkPY94Z
LdptvWApjYNET/mu/X29fwUglFsLGoLeQF39zhY6IbOd30rt+ZylIw8z3KFBIW5S
el9HC6Ou0ChxDioCukUF2ChHN1LKU5SBJpovZHNXVU+hihGGUNE47GQUfC646N+M
HkhELUVVF59ZB2ztUUKu1NvIznyZNwBSJA7xPUZGELSzl/24V9vxZiXJv6Po+Dvf
a3JWi1pZROjdBJF7XCxyOkJqH0iRUzkjdjvlCLzNjHehiv4XyWHs87+Ot2VllC6T
fkuibwd4xr/HWzDiq404CfZiRRGs8yS1/6xruF//3Mx99ktBq6wUkF7cuqJKFNSA
9NTZtcdYTE4e/rLjpWleClhvZvr4ACzj95axRyVvCNSmVihjNU8hlxc7h2h3Mope
ttNdrAhyqpqeQUVyK73esfjP1G03MY+PO25ACwjlYK448g5h+vxg3ExX5hATinxE
vthKZb/puwtTHTwwWCajB3weEgH6NWo3qcexMYNQR9VFhDJ0Cj9GpfOBTEGDWqtY
alqzSSsyMMLS4vyYaBlJ7T+1TuDBV/FHA9Ep4AcLj8DULYgos82acDLwJc5/kzSA
SqAgyHp8WZXMofjYYGK3A+nnlUeLmwez4sJqXsJLGC5AB1Am/2KcBROw3d7suJdI
w55xdNMO8YFYJITLV3x1j0Nv4q4OZp3LeyXuxTkzkAb/MhWCcNWmThQd8ZB1Sh8E
fXOTPyWCP7CmBtffpIp63xpPgvIuJ6NLrcs9+PUfYwIrKnWnqLu2f/ylUuQbJdfk
ZnpIv1Qng0ckX5jyylqZfsySpgOgZeuOfFxk5zJd+esL6Zu/Lr/SsB8ANVJUdRQK
Z7lJNYDvO1/Ucx96ex+FR8cnHOM1Zq/U1rACvUrl2J4SMUM8ZFbyu3b7UnOwv5mU
eSsJombcOszpHCbHSQVl5ZQViiEPt/Tc6VunXCJSef1pgYxXvHDtbn9zfnRmuY9Y
/5kjhHaTi8oh4tf3CMNDL1YhwCfsIg/fkyMgk5GaC+DS4jKnqA4xAStGxmnXXjF6
ETup+kcVLLV3VBlLXTlSTdjFovy7AIqLc671iLWR7jn1AkEWlNq1Eu9r/2vLRnc/
PsxlvZbGXRB0xxNY5et68eaBr7onK/hGLv5MD0pw5PweFBuHwbm1SppwDmAKd+P7
nA7ioQlJX7/kI5IM+xzhjdj670oAkqmjJ8e1OEir+7XMRiIkLl2I8oOfOfHOwZz7
SdFptTbfa7kkfcVjbw1U4ZKSkdrCiDQkbUwJojmz6ZMo2ZcDRrso2LINGr/fKOaE
M3uu3963ZnfAaoaMI3IcBMjn582lS9R2HnF1rALO+9yRNB9EU35d7Y0J9g+9Pcon
9cNe8VkT981G8aKSJAslSsZ83XX7PfJAMYha+EubeNtHfIbFfqv/QM2596FXQACL
Q/Gmsnbr16DlKM6uxjCVsCL48OmlzAs88YtOjzoE8p4GC+Fuo5fNLczFJX7UXHDn
UHBLJb0rWV39Jvp7hbhanmo9Z6Pz1XX/qQRZc6i1VMxIbCwUK5FF+J4iOrCUrlT9
hDHenrpMo0D9WQnTbXQrY/F5mV/rU/9bnjlxJd2Oy2gzk7zuFGVnuz7X489Qb7qz
6lrXYEcnKX7cN22NUFer5ov0lTiXcfuePvPaXO25uU1ViWdV9LxneMhLruOZ0jXS
UF00asqozKHJ3u5L+zmCdRSa5j7y7uyodldUhAYXYMGnEqjQdbddt9SWU2sf6baS
gUQ9JGvF4PiD+rgeGxOYFoG3xUQMVk6zB5zxvLPPeW4ie975PmgG+H8dsdSfKv3t
ciUMzNuJZAn7Hfl2D/zJzHghjUKt+LVWxWVEVG7gfTFltR9TrM07R+5SCtOc/LcQ
SKaChqrnVdHvvHu2DaYQ8Uke9TKMoIOXQrycB7enE9AVzWiyxEscIBmcaXTIDkd4
em2EApqu1Ya9pIaXnzFxw25/66pg9zemU6v2X5r3bBe1iIwVuiW6/bC1Gs0nzBJo
WfFRE7qunzLXPAsXgmpJoQIcP9d0IuqZkh7aoCHtsd4uhNuD2lDvY6fgpq/HzTrI
doIbM8xFFOvT7Cy4rUcGjLzzc2Hv0ccKQqy2pZ9wxwdTLomNI8geGGPcywsoYLUR
ASuJLEoMrs4mMroevHbLwacUxDsh/RMWg7anzRN+dmYOqEBvjdPbVNedvRjGMRx6
Z/aDkNiiuT2OnQcmwLSw00JJo1L8iiAXiNEKRPQ/Zd3SMSWSo4mzRAjUN8pTV8NC
odBFu25T6bzo+vj4Bnx657+zy574FwvKgn54Td7zMqiGq5btlEaIa0m61l1MZRsa
462lN92+rg99UHzdtx0Z7LBjRnjjW8rlpSDu6MYdzM+PCUkzZ8cNlAI+j3oGscoA
tB6HMDO6XGbz7TZNKGZMk46c4B9dV1+RhT3IOvVUHS2Tb7nCjY2Erb/O22/y58TF
LTn3UA59te66lwMsV4TLXEfMPoxIOMV2Lh5PwkEPvcpTj0pVDcwxuyMwiAZm40/t
UjIvkvavb+GWbGoD/5Q/SCL8lSARvuR/vrzS7ssnl66Q+EaXwKd98RMU2BrU6s5o
/o5Qx+25gUlEhZQB4VeNuFT4DeYhqnOKbdgpL4n6LzjAis7WtKVSDIBtNngint8z
GkIn+BK7TIx4XNI3VlGRLVPzgNS2yesoznszAH9uKPjiGdbBXPiy8x2YKNRfeEV8
GRo548/4YdlFOqAujlm6CYru4J6g6ljGTbve4+wGUr7wVxjTcDOwo4/ExVRVeXnq
k5BvGz0NMyyEMVmHRp71JNLiBZ/E04aayhf4avXBFzdvq/nRFjrNtS5b0Jp7cBDJ
rf09TBfK3fA23FZa88k2IcxJHM601JtdE+dQxU2cRN9xaQQ8IYiJnWLwqtJ7RTS5
RgGaK/cH2fTce3yI/92iU25DdPgfweWDFfWDslIgceefkQvHxQPuDMOrppHTm9n3
naEjh8kgBkj+PkERes7ku3oCCqO8in+5FZcHCNKCTu37yjVtr9vV5vM/vlEg4knd
+WkeV4a51A1Y0F7WO8LkhdsswVXnwT7XbxH6rIuk6BUFQOoL+dmpH7wVw1efWtcv
Dti29JEpv+qF/43JetCZ3jCuHRd/mPfoAfXglknMOXcIPF2IwGhfWI/KQhhOvHWA
At8e6ozFuxFnEGvu11iLAn6hJ/Iuw+UrXCGNcmne91LpCIkxIH6xLrhX+CQicpYm
uhE2/Ik+gnoVjL+Zyb8xZh/bM703mq+dXOio+BEZ7M1Kf6BZrjIjawZmM/SLDQmr
3zpORIJ/ZKsnGRJlKXQzbAE2UgUYBhZY/CFX5lSRXHQuI+M7LofuGfMVTcf5BGqM
18O1fojBjzZmXeazL2/L86JMq58ZoHUhq6VB5Be2vxlkdzSJUJ5JV8wt6bRNkG22
zWBb8Rmb0+EmHlpjNc00Zp5LYikyuPzjJWNr2LH55V9pKheRt1kGo4T3J1n68cT1
v7NKKFDkBfvMft9NHUXIff1bGP3VOb7OOK7KhsUhbusMULC3/KUBQ4ILEh3IwqP2
mb1ke8nIPd7ejGmf35EL0UImXTDGfjiqjaci6fTTNrgHHz25obq/M60AcnXd2wOH
l+HiWrZxaB6kIbMjPkshnBqmHLFZD6uU+EntFwVrklJD5maEp3zMGKMJkaZTqz4o
3N3A1DchLuONtdhsBuWo55845ruCtjZURU8T3EV+Duum0iHZ5/Kc7b+XtwTcXl6Y
8VaI4rZjCLveMcHJp4nhaOyKH4KNIQJu2orQvtCuSCx0Iu/st028dBI6QidZXVoN
R0XM1p5o5PmJXOgL+CKgvFrpjR5aqfRtIQJsm1+yhVWbzHKpdY9vrCJ1mqX25wHI
Kec5ozW8eh71Pu1aUdHOWXUN82XVxlsOCGMZoaYXJf849RVyBvJOFGGvFDPN3drb
l+J1nBtT6AYYGkwDrcmMuX/5aPhMQcqL938PI0ZOsEUGc9iJ6HbfWqvOyMCtJxns
svp+nZWl8spKGJ5r9Vd9QJyocPeG0sl8ovN0U7y8wKgQI/l8Fe0KPDZYxDzKkBCQ
Mn2aHRCxDf0V5K4muUE9aUv1JKU7/nGHagKzpu31Z2Gt7P36q76qI642LcB368vb
Rdz2vibZTVBrPuU6f6PWHuDpMaLuEwaKA7G9yP5QyzPh0T3VScEwjte0zuKyCMLg
+5xuQKbLJsr+V095+SlDqsQIcgGM/37AisFTGHA/T43PfjDfgEccCJ2G4JqLlHHQ
gdsPaOCmx1xYPeTIxgXTjMm/FnskFU04Vy4+fiitX4QzpkGgrcBHtvkMc/iZ7Szc
YanlD1gRoV83fmaLJETTmQ18ekM9SxN1942nHNTf2Bgwq8ErhQSJa8hEP0trLKti
BzWa35XWC2bH6oYyWdo09srw4CuSATELCjemxZHOCwBz0JFjZ96eHPkXqWMfRT3A
V/nt2/jlD9TZe4JqnAvv+nQuoL8kJo6CVoehYVojUFht7LU3NLgdV9ven32Ln+9u
ooIRCV+Fb3wYOioNH0v8opkOkQOMTWd0RuS1itmMZ6iRCypFOY2mDuflTNmTi2UY
4flnE4Wm2Q8fQEZiC+0u7+bYnvOAYzKAdPfaqnJUK0raMQZh2xNvHfKEe3iRYtqw
uDKMWUKn+rQdyiiYjtolWUVhkGfIEnZLZQZyhpnoe7tVPIByolHYmQG9YYM+E0Cj
/EptoYnIxRCJuJBALcqPvuIz8DrZSrdop5UBUCtN2YkknatA0RuFfTT8r8mch9cp
axmVaXSKA9RTp2Xzv0x0lePpvDSfpG0WVmtcbGWAJv8kdAFBerQvIwE0rzIdZRdw
/8dXX+Uc99d5Q9PAoFkVIKlHhHVgco33iu0HBDt2Mgp0MoW8aqVEDUXp1ROvRItI
TykeFCyYqrQzrGTmVS5pEa2+A1mE/LJexc8Li5RRu82dSaK8tBIXXjLLuryekKEV
7V9zZ2x0DcQwg8G3sf9eLFm2sqa6xn5mSfx/ovm5kg3JwiKNU0bfi0XGze0VHm4Y
MqRUiN6eK2axEcHuMdw9KmjSPeTNyuW7SxZEC54JU6QoLYxr/gsxJ52QzQg17h4n
3y/KXTYhO6R1kLQdD1asddWM/KnyHyEpvUOAjPBzQv0Ym65fLzoR9xo+Qsf9IaeW
b7LLO8LnpevedkQbbrtV8kSiYx50wPzHhuRFg5gq4indQ72NWUf4lLAP+mu4P+vt
ROlIU4gt9ta0qLpZSiaCB0KzMVwvdVjhgl9u6cpCVXgitJtwq8ddYZyWvSGAXRiK
+K8wiwVWaqgzfU9vnv2ruQ7ANfFzSm32AyO0ry2KMWkEDz8iAK21falgz6Pn+CFk
M5N+GW1DFJ69qdCc4QFN2UQjUV0rV7HDH2dhbD+e9fnGgwjyXo18xK3cP/OcNZmL
bPcLL2GJxCNHvLDuWiN/RlcBgpi70RQ63doyE0Ehrk018M4V94po86j5idQv3b5W
r0efyMI7JS/74VR2dvUJ5DBEih+xzJ+AvcYw2W8m/bDuoJ1nlzligDwoZToLeIgH
oaFKX7oM7g59bwnWWysqsjr6Dpbymx+Mzoz/65fTKdcsE5j3ASVqZ1lUzzYCWQXT
TW3L7CUz5xgALP+XTsNsr6oHNwd76u5hmvMPRbjNWo2/RcLH/PnJb3YSYLf5SW8Q
ojCLxxUVvDHu9RHGB/M0XP3ywHv8lOQR4svpqrCXKRVCnlKvVGt7Q9/pPtv1kacz
CxZR3Z+m7U6g6s2I4Pk3Kbuo9slNYj87idEuSz2Ecdd6S1P4sP6zvFPSBJyhJa1I
3IUHP2wgnyd7ZonFiMO/AlG7/HziAJjQktSMDmx2kGkvQ3GFnZL8L/RycM7yETZN
PTSSKcDDMopMK5U7C4fJ0jBrTJAWTIld/QACkZMHewFg7J/z7Hw//2ZU2sF+HjWw
sC0ks8NXD9d/itRqOQ9oILq2kNFUw0lEsapl8BO5HEQ7+NEDlmQ7i962I9Z/ouOz
e3vBM8St634DhAZLayLSkK+W5OVB9Vf5spkM2WXYiwOzufKyubJK5cG7fzU/j2yY
mM7o2CSzZxCPLYulg2NET1rkYhHf6WHqPgw3+n07txzvBlsFNhYrP/d+Yja1mjKk
lE8xqYPvlk8JtMrumd5lUCYP3grvLUY29aOadsvwmou8KKr3LExSE5PiaQ89Fsag
jzVacrEqWz9PjNNS9hqR8DGwVIqAVP+vdiNX0iRRplJxLKBz46+xCcnHf+eB0zOl
3yfYVw1qfhYm38fg8YdskHLsbo6IXWfqLgNPLAgXlysHDM/uoV7z8hpos1QZsgj3
vofEBXSBael9Ms9AGTEi56eg6wG0jJkrJa6yyGabICwpFIRtPHSpN97nqmTlaYHD
RgrfoJ9nLcTBvmouRRL50g6hJwvnB1whLMqZfyR+bi3MrtJiLs9vKRxNUDbIw+Tb
GvRjFc14b2iaukRAITtqDj1ZTNuGb8vW7KpBW4oyFhSgox/96hdE3JCEURIotJAg
REkNBqoq0LUreNMmjNNmLvVn85dg032F+HMdhHqIB9ZerjxAGjsQJfhZiFuTh80U
KyEzdAalwGhDhOexkcD0RkHx+86jS7N2VmX7Tjc42MRZxHH+eQvDBfwD9HyOP41M
DA+31stBEA9euhq6Yw52c7FJD2pyZcx62RJBxlqxZ4Io5UMhXS5NHdHZT8s/DCN4
eqdTI5ms1yVvLhTTfvtqGRNXrWDGJ1bqpujsWbXeNK3HXyJvJGprVIeisfSZh5lS
oIqYjbWD13JUueR42wiZl2IfiFzmDYXiF+PWIcAueCavKfThEmxTO86ONvlysoa5
QrSceh+or6Df4FbkNluKtBMPaOl3THuXaqllmwICTXh5XH3LXfT+iFV7oWAi3PHc
LysTo1mt40gR/2ZTy8y+8+L8j4vGNfo9agse/htwiyuToarv+miChN7WRIj8rAOb
BPIH0/yBBbsRc1+SDGLEHPehxY81iVdEalQWL+vbUIH90F0ewKwVTOsyzC+XA0GZ
PaepY+9PfGP+rCV+aZ/JsxIEQtSUn+4t/VcE7cHzdO4oPsb75eCL4sXihgabDNBK
NZIdlHb2sMdGWDsiocqNCfPeyIbGhYqsr9fVCC9uvLWESNvLShuJVUENDfLgjnhz
u+2aG9Tc8dzqZhM3wFJ+7/uM0uoPk2Lniy9LlnzxhvotFIo+SrnzOY4JxmLoc8V+
0CVaj8RekYiwvl7zOkmBvFTR12pPBjkcfpCj+6FwO36PuIyYszhj4q+v3VeyFZAS
7+gHjl4g3hsjxC9tH0LfngfQoHNMYUPLZRBBHVHMucCC6Anb7XH9IILu7wM0ntbJ
2PkbNXshjFEiYMROmC0uzGQ8g7sjE0Z7jGU3Yvp+hxVhX6OjOZMj/5F+eNMnkQSw
elYNl3xPCndjngmO2cULr9sxmh2+EQr5nNH2ptB+sJjmKp+3r4tZE7LoG8YAVX0i
p+nqif70pS5Y8tzxWzKX1LK2q65zLNVqDp4WjbPdMUj7o6tS1bm35vSObteC1LSx
1LbgnJYU7EJqrDEbLPM8aRakS8SK8hWOJuvTaOSoexniOZlCtwPe/ROVSDyvhjin
t52S9xTpN4ZZtlFy+K0i2c+3jR8Jbp8Wnj7beFut4UgMTZaYMR8ZPw1BrubAjAST
MsNvN33UebLBDfwgknj1N38N65MM+3uSNyxhPiBBnDYGZwkRDgWz98k521ezD2Iz
oA4H9jfgiNoeyViTs2vRHqMYwBSyfiGEUADp49LU4z4JT2BmaeCT9hxn3iEfjyJ6
52xCVdluhq4K5X6yhZnUwrOZa8d58KqeiI9PTTZ6Dz4VyOYsT3FM2ZlBSw5ZycaG
X2nuzZ/ZHs4gCSV6Kl3J+saEoO00Ksut/zgcnNXMEhwjs2E7kxlrIRt+umy3IRtV
EPfEmuG6fDgNrYT9rw4sWpTuYskpIcAz1T2c+mtEjyOsOGBsffTpoe1M4e0tYOzx
CJk2rxyJmsGobdyN237odUO917iNclOv6pFC0SLq124eCjSUWM5FEJCmMEdiFsBu
hbcZdtnXPQlQzcsWq54N2rfoTXhM8Jccb9qHkWQNWmgD4ZGrQrAmNYwGa8GXxCZH
dcTJKzU5tuJ/HQiQKfwCxPhMDAyvYVx9Y+emo+rlWbYFCk09Ephiw83elhfawRAU
ve7j+I5jf29aARipe3ktohpdQcyKPJPq95vRoHybfIPo3VvXT/orZZvUjCtkYHLX
RbJsEXrE1YAz73Ii/TaG+RuoBtb6yiyaFc0aApjwiT7yyhscOJtfTjlifKhQCA+3
tnz8wjWvWqpmqV14yf/nCNZCLK6ahxpsh3ggyJxocVxGRuGyzHoUWyyli74GLORR
RQ909OSfTHUJMqQ880lHEPbD09vIsH8VwYs1HmTWdx3/z7EPalnm/hQFnQFx6+NG
8KJ9cwwrqXoNaqMyjq6aQSTKiDnyts/QP9uQutrYS8q9UBGy1L6Zpbf0WO06fRc0
zJXCUdRIkBKWudi720UUyxRz3wtBC8DKj9t6VjbPZlmjOc/Q+p8TK2B3p3xZfG8n
gTBpcdGOfLdMzhUtsOd5JMBmIcfQJR3kVOKy8pZmp3AYaBeIlOWNHCOt8VcwLhoA
8lIkI44TONwyVYLlfmWfT/XL1j/MS+znyUyZolX4ZI9aPVaTxbfixcehno8AGtFt
365T2hfZOaPu16O6Pj1N7P4KBmESAI8rd9fIJxpTYzaBQZKtkJyW+KHkq8syreMu
Gv7f14JvGLR2QfG+b/SqXN3WR7hP10zYePtr4p2K25y5DoMbpuYhecsuA7wCilw/
vbcUurSXZfZ2qxd4n/g+6JxCes2fXLf101AoC4L0GvlVKmMGEx6XC35amBelvwJz
j24fcyMvSS36IpqjUmPPSBYqShioQqnOIThl4tfZ8rUEZAIGYx1qlNQXsGA8g3FM
1EZGbLgMyFPBYA2DLCYqCWjZ5meSNUEJy7WrwuMheHYJBQ27kMAW/Yjpq1g+vPLH
LZEFiOryOsx/RvT6S5aW1gowfaEbvBy/XvNv5ijGXVs/cSK3ZxE/rtYuh3ObhT8T
82kxn5xMCr4eDPsG5hlsVXb0GrYhaabYR8LGNPxIBXhHRLMFRWvutfZx7l9tYGpz
AzJEfzb5thAJj0ZGrEoW+dhv7zqpl6i4jngI8ne9n4I2ya4SmkK92nGE+E2KV4l8
PwbpQSWaJ6OIOlzyJkQwgaWhZlbnfR7VNKuotCFmc0VqHzmTcJqgs4qCqxc0cDeK
93JG3zQaOhaek/YH6Ony0bFvQ1TywKA+Pg5fQzJk31fDRkicGpnfSZJYbB9fiYEl
yx1fj1xt3FkjolzlmNpNnwTcMyU0wkFe0aljvHW82t/UsogYF3+DG0NTN7gE4C+m
8bzcsQs26LB7AikMrRXXv4jUAAgs9nhLIT78XDHdMocnuHZ522QTFpNbaz2Lrjwf
AYI9Vl7tU0A+itVezeW6yFkQjnm12Lk58NEAd97h28URs5l+aCfwa2zOQtk1yx12
3OasxO0Hj7eG1HPK9XoTW7fzVO/bl3qenpuqUSx04D0SMF/VzjU9gQj3hDsWPN8i
BiQHnQdTgG0SgkWXpho1DBaznLeSiI41IbJjPTXHMQhGVyJPvqcH21pPUiEJBDQQ
HuoR2KFT3RJ6cmJWT3W1pBRRVtckAYs+DqtutHhScEbfJt++EUP7Mzq0V6nINACE
QXGykwlSXL94im4du30svUz/f1AobB1YXe4RwM6aCbaoGXpO2bybwKgYd38EO6fO
CeBelfk4B6Db7Hnp4UsPIvfHuDB/jSnrWwlA5Z/Z2t29YwfoLY2uWaObJpYPc0YC
DQOI0joLGZ25vJdt0wFvuAvvYdLDb/ioXyEvJ1VImv+IUeLm1KaZwrFl2W0slF+u
QH/xW9CktVmpGQyjLgnAQC8iGECEOCZTOMFa800FpYOdukPo0e2FEdGSwFSe4lfU
jVEMg3f6m16RY74BJ2cjoVfyaZ8XQWATxzdEeSl+ay9hROWFLk01CoDS5aK/zM8G
11oBe10WOw9seXNLIZApltEORCSYE1hfYRlkl0mcfce6ODgAPxxrIQnjnaeiIE3i
bR8TQcTIOcf1ej6crLuf94t6j7T13lF5WF/QQFxbfLA7c3gbd5dxb8tnHyKxXHfk
bdupy5yLlRMr+Ze+Fin1TBm/ycNWOWlgeGnqMx7vKX8R1rPGPBqYkRKL9zA66JfS
ISeCcMebnaBaUmb0k6XND+CIdeckYXIKykaCezS9e98Vk//SbZgqKPUSTyyDKxvx
150M4Bdx9G81w/nRETCwbULnSQoJgMMWkv1x54aaehuEK6UShhvX5TtFL8LQSdE0
GjGDuk0WB+S935xnB8AOp1SSpNJLqdkTxnw9hOXwHsympD+Gej+esQ/azjYuZji4
sHesLKmrT6qu9QRUD9zwPx7iUQ7Y14VkuBGjDgWPfUi8UgKFEyhdBr5K7ikWpeBX
zuXV2d1s3nhoLH9u5enfEpZVgFek+nbeg+c7Tu7fT3Ftk0/C+Ry42FVtNmG5kdLR
+7YjiajDXEADB02lL+Mv1n8cEFPot6ZI1fgggUtSLjXXsdX1esYBTiCd/96t/bbV
O1l3xyknYBmuZxCSXFDS6NfhIsRZWGX0z/EJ6+9mC+e1h2ozlyyuckd0EHY7FprA
vM5CMbBjhyCK7dObrv8rZFbBcpO5LpRiDD2+9CU8HKRYm0eTlCoAj0PHhjVf8MR7
JAUpCh2TgiTO7GFfPAkwf6FPhlWaz/EaLr6ppxYuydh8FZroHYWa8+NTGQFkzX3F
3BYK0E7W2MqekSFPEMnuM7S9Enj0ISnAvolXfNxCRZlBd5ztThepviXQFjBb47Mo
QbQ14frwMae2vaa7rCv9617eWW37ohw4/ZWo2tDVTanIoBdO1dON3CXx5fjx2ND6
ByRwf2KPgWXyM9XrC1BvwIYRVdBjTSEAHsFJCD1YyQJH1kt1hvEH5J/qjzq6dmC9
emJ7oO1ei6C23CaafrLqrUuGGYEwFbSKP8IgFKJUnUABd1GgMsyBz0n63px7KQDY
mYaOZKvMHrGA9zZa9MAD7ts3JhCziDSL8QklPauyYy6J8bPK327kNlo7CwW7+rW3
uavigqitmEVFPad1uxi1+TiNrK4vqp104FjXCHJhl/ZNSFRKC7NAKXr/6xE37ENO
SgWZfZ6atLh2kC9zDkLWnwTEoCU2/W0rCDlnT+EPcSOy3VWc6azEJh95r+IustdD
iEZI2hqWM1Fg3Rc0BozJxlZXU1aIvMVNop8WUsYg6dRShawv18J1nPE6G7LvnnE/
0ff2cA9WaCfx1DIXvcB0MvHFA6xMpW70TLzQLYNuPWIx+rK6MZ7wwzrCD34xpv3C
i3d9oBjrQrldjF7d+2xsYheJ0eUWPw3gEsPv1hr9bmVdZfrdrcMRxfJ6oXyzm+oD
2yDzHI+WyRYN0Ewl4vRa6mTMWbTH5/ruxVQc+Aqd6ueOjAwTrw/Vmq3IAaSSwjXO
PKa/m6A7k0w77YMG6KAQBS9RmOtVpZyrOLCpywPYDKbwWSNk/FZPgL6OnqwSLCg6
ZcsbNEziyTv2iSQz9Fbdd1YsfIb5j9UMN63u2XBGK8Fg5e21gR5AIq5oToAAz1v7
np8Pn/EE2f/TMij7Oo+oYJ+ZpQF4oc/ohwq4w1BfWI8tZKOkzVWfUPVsNxWfUA+/
HBJSVWJHQcLG2ixlFhnn8Hs2/nRzR+HAhU6XtAapGS5zlWfTixKgCImkccyJ9T5h
LRHeJTtoxsjTqJynrNexZ3jQbvjY55BPrAeSTv74o9I7nvsid+rFNXF1Wmd+2j3o
WRkvrPxb+wcVTrBakpNB/N8iCniRG0S1VoSEL0xakSGPx/Z8xITeXYuF6i9ygCFD
5RXc0UiGHDxX+++7T1a2gXCKdhVgFlFkJ7Q69ScjNOvdty9iHM3k2hfdhpXDi7Q3
7Xm1aiBPUpfqwsMyWonjg37aa8BnyaXqGDsqA38NkAl/vpJ8JqVCzmStKssJjKs9
N75TShlClku0h7yYGe+CAB/gvaqdyQc/e4qf0BmbfaQP8oYhtWdGFgI2+xxW/3Iq
WXAXRzjLhCQFx6rJ1qBUGcn4SqhNa4v51WZEMjThKqHQ+9dZvcHFu+3/M0PBCawF
2Pd5OzhWGYK9yf43fhucD9IuusRvmiah5zkWNzfZ3V44rB0b3HXX99IsIYPZ8NfE
pu2iOLD/TU4t12au109NbMnuvS1/aNuiU+CSnNTGP4IRaYUS8lQdhvobE88q/ZRP
gjFuux5lWohU8prKK6TYmVtYh+z3XscKsHhwi5Ue/HdHWPFh7yIQI+j5M7bYZvBc
jCmFnmqnGfc+h2iMJyCZvnFsF6Q42aCb1JRVlJAlRODhnJSUjpF9mQ/zRO+BpPsm
/gt/Kb42RIyBR233tFjW5ccs7rTXY/g/Y5egJ3R5QW/+d+WsRa4h0pwCttV6059t
XQBK1DA/Z81UcDQn/l2raLgwVts+vVAQc5ltoo/EHrdo/X0PDvN19NCg3U3oZ72C
4Wi6BiCPUZVVTF/+hOT3bF3GTjlXU87LZE5Z7bINg11bEA6jw4p3WOM2nS0wbQHk
eOjmCNyvg4avQo8ARB/sxDbkccPLyHLgrtb+s2XuH3EAt1S9RDTSS4rbY9Yz+2yV
5an+iRm0TKzMifq/TQ0MVHk3AT6rybnVG9mNHkkVvd/Rq2c4bQ9TLKqH9hMgvAC0
gQ0MCw2QMerfZO27YRFNL6IgHqSwJTqWcSkYHG2cUKKrTwCGgs7nm3zfQa8fxDFI
bW/1+cBPfq6mkibtiwd6ggKyFfknQxNIv9hID8FDt3ABNfKds0blmHDLPbwG/ISP
TLSXaKzBtdp+RdZxfdOdTupTjsC60jJnoIavKBpOtACD3vehPdH33vzx4wKizH3f
zm3SZ50BjmM2maN4X9ckO9FLSp3583jFe/zSVmYBfTIUEKLoa9CnhhEWX3tWQ/ME
IpuAqZRb8tTWkBInK2IvrwEbayuEAnWuIb25jhMmLjo/+theORMVLrZYgor26jGC
wMWqg6sv/LVIEXJ2Dp+0FiXtuDNy7Dnii51tQzeaKL5U2/DfCXPuDT5EnMVaomml
oHE030oPYeYveKnBUTScnx7aLnVeXyKnE6EAIpnOt5fJINGpo7LxTzbXYfO+EC2a
SqY7ErS8SJnaDR86hISOvZpnl+fC+9+/Neqp3Ie7l/0/nNOrf1RSzUK5RA0rwCC6
KIekbgDBYoowDrPDfc7z2k20Y4LJz65zgZRa87j9Zrp8e62EKIG9M7FwKk4JItUt
CFf0879lEX1w+I72/2HRCmWiY4YiyPNj+q3OJ298BRCVzjxE4Rq4k2RuUPZj8sSg
IrrOuS15nB+lBRFtZRCE1E91CNijfUZVLAFikrjdn4ZY9V6yQTNwKe2RBWcpcMqJ
J8XXlcM/HQddjDwOYsojYHOT1a/gPCw37yhPuS37NRkBG7QE23/Qxql9LF+4KdHi
mVd5GLh4qh4pfQJMhoJ3JpkmiR45Fvd2FkR/rzjxmYXdChxfiL4A61KxcgrD3gF7
V4cmvJ0xe3mIe1MqW1W688HGPM3ML9W8ZCNAQFemTMylgovaYtIUs424094g71cv
5qb7H0J5TbI08SNTGrVjeJsExBFaWFNhZFA77EUPKcdCcVUvSOSReD8tscqzmF4d
ZgU0cLj+F94ZJMGn7u1Og5631w4tqZ0UZI5gbxpJb/DDJInWExN9laYWSY6Rap2m
r86eJ9c+WxROJpugLxTixeTVj2mUO98Z+NsvzO7sH53GR6yGjwvyg9CZ7m0uv2Wd
KqnxxGiwRJATc/of2RTzzVUKabqYYCWW5bojotY9ULmLG71CPs1YH/HBUyulifsn
riYIPG74kviXTCYt8pF4d9LRd5UoKzllXGn7+UPQB7lUUS/W3DDcpZxleGLdq6nc
daa9XDxhKlih8qkS/ggb/7xGXnHe3cOAByKQ3LTY8KvhQTXS9VPASRLhipkz2/ZR
0RIHaBQYKa6fXxn5W5NhMiiRPPYVnQ8GCZDW4Ik+QCWo6bvJ1yJ4XA39SulfWAZM
cut88+19QnSGrOcQ8dIW104jKcj0cE9XAYhVl02VRG2b11IVT1NDNfEBIjnD001Q
A1mKjByt86o6SLAngC31zCksZJzhGq/IypS6Vq+sovjf0QjnIcFRKrkW+yL20q8i
pbSqm9JOTycKFI6cYB2vfsOfTsFf8R5MF6sn1kkVzincyKGQ/FG1uPib274aJt6v
chbaWMmqw2icpnyM12Q6X12KUkcQ8nD2zEQpLhjzgqwIIRAWp0gltkBOa7j82daw
fXtGdmpp9pcsyQAOy0VoLWA+dJ/NSAibbN5MwjkSBwn6ROHKp0EhiTTOLKGRI5LY
Zkn4vVL3ERanJttP4SNaWqrPsPZ+d4J9riJPjPZTijF/B8XzOT+HUe+D7NpFC1pL
9SsR3hFU6X89rSd6QvquLdKezkiJtdC2BjQIax+kh23QvvycfjmhdGwsY3mQNqsT
hvtgz9RNPPBNbwNMYAA9yuNTWhDlxql5+sQ96GGUtdl+w1bKw2zsH5M1f1sFzz33
fmDbACOdD5UUtu7WCay1YREnOBvVU45Aj1MSzHxQ+EzwcvbqT99SVget2UuCG7YH
Q2vMJ4Mz5gduXmUb2HW8MZvEov0e9Pvmgi/Zch8vcg030lV0ntjQ+jWml43g+F/j
wqcBOA60POUckFnrtOwOrBMCYmx52gaZNhmdbXIIreemwWyqQQMHbauL0nXBHipi
UMljxwcp/8fffQ0KL22BED7oukuleuvKN6RfJH/F8l5WJMQBUf3dU5H7cwfUqAPD
ycVxeS8bJJ+SsBDjYrAdBt3Pvlp5n1xyvsR2oh6ZMSB5KIvDrrUkw6qdwi1/1xju
yvtFAjQ8IcDoAxs/3fB56QDcVzWGy7ClNTX/E4FkSBBbgCTvzyY835fm0rDAqmC8
rjPGhlekxPPjCiQj2nYysPzhnDya2yAOFyS5WcYkFbHKD9y+6qYCBzpMNkfW/XVj
ykyvwbz7HFCHHBOtANhEZ9SZUqEz9Ukgvq4z+RParinz38wsIYuCWqmxe0RmH3xk
32gVF0GqMnqO/8zxn4uVS4GC7XvtaE/13v5R04Jj/59T1vdJP6xVKbuObNHtXRzY
hIOIcW/9x8xMx/s84gizCOqTPEFdY7EMAZvoNdI6HZvPuvihunvJIhfpZOEbql2p
m3hGnkJhsQbdpf9Q0ZGaLpGz65hiSek6BW4D6PPdAJ5lRbGmGfx00RYFqudEEWwt
UmPMxggueSZDVF6Zp8CPpyKbN16xE/Nm8PwOswmR3cduLYiFHSALibADyju0TN6w
tbxaIRQX8oicjgtuMpYkmNGro/GtcdmjFGPPObKvNg0IOOwK7/GcU+k7IgMR5q2P
V0l8oE3bH8f18EHSlUMvgd1dSBMOzAXNBkTzQ/x3cHn/OQg03bHYrVxZPmArXTzz
K+jepPWQlihSsG+vFrpcWh2e/hDjOjsWP8jiUBVYJGuYv+9ffgOzlUUBHxA4DZtc
UWaCESOAqbxWch+7WP/qh0xubGpBtH+VD+ci9q4E5+6bfqGVgm6iowWrnV38ZSAA
1o4YJFSKEXfAVubDTFvbhgdHnyikUlu/OH9lV/5Is5uI3zBXbnbK0GMDeOB98knm
Ybnv2jRe1KBELiYNX686sULMai3B5AYfjHmpCncgzDC8HDSvk24+3Ha1u18Gx5Zb
oo0x03riK//NbCtnJrrYuKg9tzhTChzphKBiExStJsk6ahje3WfFlqbpFw+rdHLK
zk8O3glGbyfVqjbyZgexDkrOc2LUFFZr6nEqC8//A3r1Wx2LgpB8zRO6Y7NJO6/e
5uLfK57bPsakKPaYJN/A+NlhaqEbPQbS2b/LQZUspItc7ADh2epmHT2kI9O4LbYh
7t0sGQnT8P7HhIfyN4aY5PWfz0JctpHUibZd1nrUjuJfTIc2I6KF9FXLM/Fu6xzR
xPSzlc9gsWeyhTSnM+ZCym0E4k3i8+l1nrjZOvf5FROtMUwUgRMZw2CkM1253Vev
NByBHU6XhwUIAhQIuXknPlbz8ohLp8M0LEolf88pU1zM56wxbKDTBUufZa2c5Oe1
9dmRcEUUsBpOibd9RbnQr000gPucgd9wJf2oMlj2lGgeeXMKdtyBqpUj8amw1wo3
4kTaCvRceIEwlMM6MvnypmNQt/zjJtS4u8Uim0mu00kubOrJoWsF7HDfa8sMZLcP
BkeHtDZs2Q9l0mA3gLGGHBW+YAo3W0JG//WoWGaz0VmOgCPR5dhmULOJ23siBmi7
m7h7EIoZg/ZgoXu8tHkuOU7ZUrns/ZyJx+13pxzSXlvA/xZrB46BP9vNPgHclzvq
JHfFn4Xp260oeEtFKsvlQ1RvWPEocVVi4dMKY84SCze5pb1ZQv16UTlN0/P+o9Ym
Kf6W/n3o/M0UEoUABTJquAJsIl0xRJ385y2vVU0f/GTO3YVy/uZ5S/PmDc1HAPrf
PXbQ4g7vFO+Ht92b28ORGwqwbKlY7k/eq7eYfrDoTYQK+OK1FBXp/EujpELfhMJM
kh5BdEfO2KRmjFqNLI3hyGIKiotgkxiBFJyPnJ9zYOKHHhQrSpOVxZC+GDe7owep
ZeYlNuYNblqOtqgbqbHH389Whn9lqzFudGeAKvgqlrM8ytBANmDfdYRkuQJHpGQx
gyeIIrcq/Bbw/GXEyYQSgG6OFHz5ayKNMo4LVNHtBXSGO10Nmgp4Uu5v/qfWm1dN
0Eg8EonLbBMNtDeIQrntrWuuv9foGaDHGqowjt4tzBq4XuZNRYnDTBMS/v1FaQUr
V2UwkECmL43QRC4p5oTqJIUojwYGspaTIzHm031nTHXTOy0jHvoh59O2AbLvjjJg
9pqJIsKApoovggaLPZ6RjXl9aJ5rwc9oolafiKtN/DUm2V5DWEGQZQa9AStWuGpq
Y0f5ystT7/UbJdTQVMlQuNa1DOz574MERNwu7pllek0Cy+NP6fyiy9+3hE3dgoqn
j1JGYaINcWGSHJtbI12tIxK9SQWyBU6IujBmdOw+MYKoNlK2xrhmjZ632GRpecQd
yKnovXci+WgldKNCo3JPJvpedbQVomKSMSbfXOs++vaNx8zRKjdeEWSsc5SQyMM2
IfHbgXaQpiLH2N9ry4woWfEFreywSEaXp3tHo6S6/35RNde4JcO/VbYN1/paK7Z4
j/08FdmZFT1heW3rKC9t+vP7YCw3dfC5uhWBYPDzuF8DpxHLVhk8Hv9/z8/YX4qj
X+oNZ4trGIdBvA5hrRIuEyLRL1bF6RThjEsNSHcoh7HOi3S0fN4RroPdxAW3boTp
wCX/CRw+BoQBNk73VR5sxsUHsox8C7qRxEoFH28DTlEyd0HTV3GlMVEnlSk43s1/
y1epSEzwJadrUjOLSvx+AfW/h8VeXO/vvS14EaRGY4BjLxM2TRjJyJ/fq389tArf
xtiwYTgweN0uh8R7jrYksECUO+BDcmFj//XB42omCQ9g6BimPWPAJiNk5i6Vba8s
OkAahViJmDvImzr7TwGaXnGa4pjtopID7mqkTpVlszRjJf4bLgUsEKEoDA495Szn
SBnRKj6i3RUAGqmz2JCYooZF+o2UkwP8OKChMggTYZsEw5ke2DbIb9ZVCOhI1L7j
isCvOciHsxBLRCj26IWCuK+YfUzWViRXqjG4U28ku7L7YkWBS3Fi/VRS/fAq6UaP
F5m65Y4kRZBdoXUH3RlxOBeZF4ivSiPLZgwOwQ/j6RevWnsNk7sJE7NElbHuQ+2u
NvX1/bnoj3ioUhXoJzqYsgk9lZVJM11EBRqa4a9eCFslk9rqvqxhCuxWi/AJIGVQ
Qe76KMVVLZZHdoG7mjx7ZifHjnvASfciOWxWK1Ry4KMKPFcKj17GjjcCm5yLAU/1
2cQcBXSFGwEx2sYeI+zzMjZ4DHhSGtWFnTIXW57YF0DVnWzI5qc2x709T63JbLOM
GIuUH5+Yo2LMOKUUSCjY5cymhpLjGPrWTDnOBSiZX3ODDqoce50cb7WbDl+kaGJK
DH6eneqxtpzDRF9HzrcaqhpheaXBFxNz4gpIDRT8CG8HSsz+h5VMtzX7YcpoCtWo
o7mQWx14G+7gi/xKlsaMzXYzn+yv7afu9j1lkwyMeY5bMKKHC8AfFOfxZkZt+Bau
kW39qZ80BdceW349PL/3POXEdkmYcBnENvZoE1XmMtKM1LlqOvUYcbEuAxUsFPAb
HKQOZ3ChkNQRnNnEQ1HLKdfw/4ffgPOC1eK6k4bIWJ1Zy3+VMO8CE+Pn3g1/Cbbk
mVl+N3479dw0z6IUfpsQC43Ckr0dAZQFjn6UJumj2r31fiFD8WpRxi9gnofTWPBV
vLjl/kxZHbj5T1tPlq1fgbqI+lCSS2LbzLWpo8xHcns/qMJgMx74SWdjpWfI6pYU
WYv0xGUv136esRkiaPm5wVrqEB5Z0IcHg1e//yYI2f1juMnIrF2flPXrn5htrb2R
ZosaqLdVVfMBsVla8j9eV2Av7oufTOFVRi2TcGnlU8iwmaZAJynBYXGxBNlOqQt8
zTWfQap7hyi16Xln8QdlT65WGpuwSOyqQGlke7j223hToNgxFleFAyUibtnI9unL
+mXaYNrhA2hdPsno/jEeRmQmUZ8z6PI8rozKyVHjDrStd03pmwVBm3SC8T/HUqlu
hehG2hW9veAM2LjHMDXrv2XQj2h580CbAIfJUbm6WAQabdLREAn9RG42DaGit4WV
XkLf1DrUPgf0c8H+uAEEqEvf2197aRJk/qU23ysQQLwsuXBnQvkDY+db3KDIH7g4
8eMzda/b215UFx5EEnWxiJw4QF4WalYAVjl+v18W1Tzy+wDeYOkqrMJafC7xUkd3
HLYDGZjvnW1PxPKkOpKEFzNpbH3WmHGfuFhNcFqm3piE0lQjiOW5rgyjeLUlxMAo
qvf7zyRCxHjOJqClxsDmjzlSo3mb4Eiqh0qC/VYVSgBJSWMljzi38FjZyDZGBJ9j
zj4fcEZmzOVWn33W7FnljjaYkNoaGhnxYZxOXrNYQ+6pz3qSTw2aNcQuZnWxONq2
IdSzzlNjNV4cvMjITSNt9vFCFj0R/BUsco7Y223WmTty0sAEAkllcqjfXyZmjECn
fIThmKWpXEZAmLUBg6PihvG7Inwv/qwCmwis6K4WKYvjwsVRG2JqihfN05dplaa3
r+XBEGB7qy3RYK3pU88PvFuncgVpI5A//PPGLQTUQLZSPxWtRsKwxJ/guCcS0Qx/
1zKQcIEFMecjvHvfj7bFy8XDqfNDsebgdOuCTx15xZgwgQBl8SPECmgrQ+6Aq1wt
FvzR4gmGXmCpkx7uRJEsLqTny/j2vH4vIR5CGRAs5jHE5xZGBY1Q7ol5D2bchbfa
m+SnafBYkzyzDgen/fquMqYtVAx05pd+0Kx0uamG55p4y0uBgdVLJ3D0GFJyMJIA
SSWY1/GCWxwzKkhY2Q09Szfh37Z2XGIQcmw1XUsksgEL7gYnEmFz1Lq3rArCUgZh
1HtdSsG1/tnqPmsFhMOSJSH29kWQ9j5ulR6Tx6WOSkpGjWwRnXOp4dvx6vbfGQBM
pskUCbnrHZRMufUOKR3Po24KXBXQeEc3lK4jrsDWtSJbgiYEs0/wKryu9g+iF9n7
p4akDczML2GXuPr+cKc8hAQ7vdR+aOlEK0GflXiwnQJXTfqqnOvZoaI+xrISyarq
AXvxUdPz+oNPSk7Se5n8ZBzzuZrVGvy83dphqJKmMkgvQebRaRit3j1zrNKRf6VB
EAD1g4mrnBiBsikGndPFJCay4Y1sZeBfXcf2wZixzORE9mUfcE3KmZr79aTvz00F
nwXvsMFNglxMsa+QxK+Z37O7PLKA2alDXNzGrgOjBTRuRChlKCr6J4Lkma2ImoCE
uGIIl5uaAckdY5r3xmbUiKdxiNydFhhclWIfcvs7dQVKkNn4i+W74VPVjUMNZ63B
x+1XrKNUSfbxXYgsSk6bwXq5eMYW8Z2MvbhB0fuvPA3UMv8G0u7WzwoBi0UDZ/Rq
39IbpQf4P8jhwhphGedKS6DN0Q9aU7XIkHJlapEAs/5xsYXYIE0xRY8wJmyPsCXk
23gvLi6Jhq0RH3HueKl7Rh7mxqNkFaxCmBJO0Iz7wnUdexQ7ztPyI+2LuvuYSeix
Du/uCgmzRqPzVqTN7k8rbxRpIv9aX2pbI/d8Qu72tVmfHO4GMnRS49CdDSqd29qx
EhYWVbN69prbc1yUvSFFpjCDvARKDskCphq8MHuDUrWMPrRDOVy6e03oBBrQ3obk
KoTQ37InakX09hJF9xDtyRYtVM4nUigMYCcRmAVQrINuYnorJXn0Uqd3CZz+Y72n
0UpdqCEhySkEQoTWygoIWGIBlm0I8CClXT0wL7bpOnPopZ9BXSINB2Zg5Zp5lZQU
E/db/3SYEuguB3v50WzAB8dQgHqrJ8covpR4q2ON5YfhKFOQ10TJOY/bEpyKSYXt
1Phu/YIPYK2IMjECXX26zSMBMTCMCDRWukG20shV/n+RPP+/l642IWARbltXAtz4
8Sr7SADpFlRL0ylOIDO8HfAciY40+3R94fidU4jAJOpnfv0GjxBH+umHNepxDV7j
rJPqK91fr6yxrBSlt620p8AdCmQrnqNzUgBOMzD3OfevYvmUjj9F4CMyZfslavBZ
J0nVeOsT7SfkGULKaAln+tGOg9/l6s6Cbv3iV1smg58sQQWodSR48ls0iOUsbCfg
PY8dJwKuwlSEltkvnsaVFTkfKugad1MEOYSDC6unwWtVqIrQp9r0q0iFKO2mV+60
Ytc1sNJSeIw76wxvdxiU1n+qAj/ta8lvKfaSGTM9Y4A36Fnmbg1SN4kaDjc6LSsO
5wu6MYMKzJ8LjgGT0IGsZy+yglp659HuqCKI5NH0kg/T52OCDV5i/WKnzRJxcLmW
f/YFRGcOUpgSPjb4zj1rBBI3LPnBhj/CmAqOjlyW6SIZBouktw2NhogzkJWk4YnG
7FzqxkhxYo9oikhSIoUzTqR7i38jpP81s173UuaBuhiNWFPEEmV6pgiKG3fYHQAh
yjmUPLHCk/wKMC+tnXOgCtowN6M0szU1TZC1O9bZ6B5f7dWPVF3XXkklrlVgKnxM
limj6KZXoeBIU7amcFKAQl2qIt3ZRJh5MD1xSVKfc9A5qts/WjBoQZqq+ewlhAk6
VODOqM6gtujHt97Aenzdv2RDx/0xw6SPFLi2Qa2Ro6bKVva76bsvP8rZzrG1UzC9
36x7AlVTfelL7jPlZmGiPWVbhrZ6Slq41mwZJF9vMBCPcTitw90Js4mbxffMQVnW
IA++AUGOmkwyhc5IsbgfN2BSFgG+JSrpE0+OjGMNAjqnJaeNLDkQss0Qq8FyKuLC
BEQ2WKAB9yQtOVgGXICv8eT8tv6UD7HzfVPLC33XdRJU8dCwYIH5jRzrBVOfiwpb
h1duRhnAfzoP3yvidp8gqpgTUsuZyDHchRLWyXYCZrHznpkWQg5cR0wNBmed9fEo
Oe4w4PgA+FMqQ2WFNm8q/6Tcm3l4qA1zxYOVE0+pR3oRWHf5tP0oA0OuKrAJN3/n
0gkCEPB1qf+9AqCNH3zoDmdgpvWsUb0SwxE9Gw5XZrgLKr8KjKXZ5bf0ao8sdJbj
yvqryu91fy5vzAzwyfnuBxaEij0ysv1Q5Y713yijdyaqCAG9AgZ6jvzjbGH7G1k7
ZhGAG09GQNUbtdLAE8Kchnm00wo0ZTSCQN6/AefK7Ext25+Vm6nrniDJipIgb4kg
Sz53AzRHo44GuzehO2Y/vfbjJYij2eyYBOLbHOLKUXDtz3UCYdK0T5sMiXXnp2lp
FwNMsN4Gbp6TUzAMgp5sqctIs+ULMVMEQlE2I8jKd/LPLqRKgHxdcIzq5Fg8s4+w
Lta03zUTG+kg01wJuTewlw2Ndi6NlVY5WRn28SzdA4U574GUrx+hIaC+7YHEYGEn
jBN1n5j+aU8ZT/G2hmYwKngIpNdjO2oaAKCTZVLZAIdoCzHzKRwSsUfTpgsYUaAH
fk+yCCl9SjOHqD79dJpZQras2mQ89TnXxlaeVcAUBNcW3sGLtR7g53UEq9JiPGC0
0aoRFAPUy3+B/Ao2seyMZu/ECTRyf+oEgiFDEM9Rk0pEcwFd6YV2hqKi6xzXzixg
XdtRNMxBe4YQWccP/LL/dZyUs/nDYvEyei4+20DiaW+Ry3GDt+ezEmc8WXluwr1U
BPclvqmy04YPGu6IwLiyDKLn0o9BJnVJrgYwEQ9gIbYDA5vUEU30DV1UJNV8MX7+
tyRHdLbWF76S9muewG1Y/NO81nSZpo/uHgdBAg9LA1Mh1KyvxKrwtgPnDRc7ZkMv
eonav4cPcrA27mpdh00rlxB34yonqJIR0zen5w7/k10AWsbqj85WYMrlMTkwNDgW
h5MDmCC8cqXNwNx2zfMByAJc+NMo+HR2Q+Psqx386pr8DgZDjQZ9wg0IJhmQusVf
PB36a0CpBsrAEUwC5feyMMSh6yWs0H08oGCAKYRV73y5a9U/8my6cXLEOoMmqvrN
7l9ILeI1bG33cuu5VLJzBayQ/R5/EjhHr97ub5FvyMELvtliyiFDyPWYcrvzmU69
ygYsOWgnrSwjaJ/S3hURlbCVVlnT6bX4hUjesxBGNEZB7CbxG6PjivT8QkH2acvq
SwJoqIk8jd8NBjbU0ZwcwPGWMM+qE8goBxKbHJv25Dgx3a0NgvQl6smcNByvDTw2
Fmm3pgdcSobRntDXMcRFo7ORwajfVzPlvy/n5hL/KNCDhOEHy4j+MjK9XEmKip3U
UxnIMdw4zzJJJOiCEnvs1Sb5z0UAu/JjAoTGLlUpNTeNk1wn9Aqn8vU0oH4fig6R
/1ZarkrCFvqcrT1KP0/GqyOmYy7JC5X/mQtuEcNzS43gXliVUmUEEaf49ZSH2Z9T
fNwBIJTXHA9ABb43IGNpMjWlpqItkHVjMmHqQZge6lQ9wzhjOL4xwlA2kjvuPTJB
o5XdcemzL50xW2JNBa100Ha54WxcVKdGCCtWzVPIpxa6zwk77UTTnUlnWaDsqont
EnXilJB1Ec7q+0VBx5gWT6cyrCCvfFQKJ4nySO9yrVvc6sWE30Wm8h11+fPhXt1s
LdSGgfyVJ5C/g4EGOl0dtIza744oTfgVZuwdUZioW7YCxj2boM1xjAiLB2qxGhSQ
KYIS+vkgQlI4ScwCS8Ij10InEkE+Nsx3lrEmgQfWE6ZrksddbSDM12zwn4RRfU8n
V42IxQ9vpX8jU2bZCwA0Bx2wxgCWFvecEfjt7fO0hArZnJ4JYn/9iK95mUNbexFf
NcMFuTWyZ1jmeNmB59n2pFEA2HEOY1zeao0pjcogu9NiDtF4mwIVa008kiHWMWvq
iIQYYWB7HidqSPYgKN98ozNkbhh+vVu06DLSRyUzju6xtE0/cLkocSq1OfS8bRxL
QujXlLJ4tA7CY9I59qbpVi9EVae6T3heO2+WQmwTI2l5ZqnFveDlX934Iy1Vq86h
m9c0R8j1DLaIQUgMmqY3j1vBWtfsP4xQWq06VIuJ1sZN4BVQeXMS0KGjFkMe+XU8
tabE5yQZxGacCP2bMMJT0bNoHnxzgX3CqoYfT9zKaOCAGxhXDublQg733MDG0aV9
5cARIll8WLN/lI9oFHPvTmnn+geLOGP7TQLmU1RsE30xZf6OB+VKrgUGy4c8O9dU
xfPLZY5I0Ek+mANLlnczq6C7nWZESPdiVzv7oJxglY3PLgJyHAoEcD2KWChwAmHi
iwve/MvY7bygK1LKRTETGmUVQeY4fQY0yWQWc6h4XcvBXFI7b2WYj1+fQO/OINsC
6jh4vVIHNUzo211cN3WF5JHEw1AuMYHAJZLhZe9dMS7m5iFjVEnHj0Rxnv0AaawV
4HqldveI4w7aWuxvWYtDd8UsupceqffysEFiLE3HmF7fOEkyUabQSIV8E+K0RRek
4PJrvce7X9g/kESwbD6Wy5eavPxwNCxR7n2Mk7c6+xrdkbzkUmbxc3oJfRERaKJY
r9yp5zd3fFhoq4BYugDUVDdbGNd5l/FXYi/UU53yMU6Ny4SNtyPybH9z9tTfn+st
rdXR6g8aCVm/t775Gb8+f7JbkeuyIrEXRv48Vj29KwB5zz0ke09BtCAy8E0fZnTm
flsU1Dr32dXTzOITiaIP4Q3U9vFZCzZFpiZ7o8qDGr2YOLRf0526hhIUyNjffDxc
r6baqT+0pghC6RpbZeAnsPCZ2L2yHwKtkrIKr6CD5pPpD08rA9Zpoh5LOzykVLmR
P6g3T9kVAoOojSUHBI1ViVxoO9NYkcm81mm5JXjNI59A5oKa6ToXtGHsTFceX2Wh
qO0kfe7/FCRLLdxQQr5ICcGrjCTxP8/11R8olZWODmTp8DsZvwDEFrpN6occF4RC
sa2RqkO5AOaCKUBYjlETSVskrRuBZqE8TIrUrAhJ3HE2s8eQzS1pP+uRv95C2rKI
ye0HY5SBfD9BdiFPpzlzz/TYbdE0CiEILQU+34F3GMdkg6deKGjIoyvTVRIJEv0l
255WKsb7kbQ1O1dGDiGy+ONfslaaH9l6sEtKzlM744Qt7q60g9z9BMxIUw/Xl+Ey
Juugkaqzj14NOwvfYWg6LIOxa3KG4dwbcTf8h1DwH0QCh/PODeIRwoqCUenmdowV
YgjTO2TyN7nxbtp0UNCwsDd0NC2cemBlQLOklVm3HNCxwnbNBUYZygB8Oj9jyx5A
FZ5rBPnpAlpZMma9wKgb/VR7iufbAOsSCrLXkiJsWVn1GCfr33kljlf70vYME09I
6DjYCN4C1mbSKRlHyH2DLS1ZWAe5UG5fosf1rJt5R+WGGUK7vwgYt/L68ll2QTfD
17JikrM7Cha+wpZbSZm8OF4h1Zi1YxiVU+ukEbEhNCyjUs6evO7CXELJCR6n3owN
qRiYJ4n+bvE1pUtTuCo+Z9GCXS3N985Sx5UZcRZ6+OaxHGyv9RNIZ8eDQa0jxA0W
WBugcmkpGkWzu1TitrWgi7HrdRU2I1HMJ/1a70KVZfnKdIjGD5eldcgvhkP6SAbb
V3j34KKVE02y9pqss8suyYtBDaDRQ2OqlHi8kQqu09b3ozuSFxWVdJ3+p103vlmy
kJER8UzqEL9TQ5blArTuJzJhjAG6E5uZnNSyvr7J86rzf69Ey5zuWxyRc6zV8BBJ
dFJM6iFnhGI+vPsG+OI7OD9zQ7SDpcIln5Gk7TC8l1+jNDVyGqyZqyhvEn1VighH
qnGzsP4s2yIycuObQr8+CwpHIaItH6Zyty++3LjKq0pfsqzjEhvXXTSt+iIu1O+2
uRRAE0Y5JiWwyoPtPaNRQ6/wjJNaLG6xmmGKMcsydCYwvaxIfyoIMVP5hHV7khMp
ocyYmSck3Zl14jEg7R9LlmDJNsQ7RMuPb9EJnbeMU9xzvZ5rrVHfQmxqrGZk5cxK
xNn+CYSC6dmLBVvX8iCUvN500OKW1wx1QQDNus1M9aSlpgxQXzS5Bn4oX78ScV9+
Nu/0qZ41FlnTwXPpnnurIVtJwU38bqDokO47wA3h5LBtS/phfQnYnjMXeaj5+kou
AlOEBf962L8KStx6PBudMvH7MN1ppsS5D7OCURaAy5GrmyyHaBsNyu8if4zK4eIq
9adf+PC+IpC5KlnkgueMn2xf0q0fAZHeywHPTSVHL7v2cGlGxG46XlSqPWlNsl5Y
B/JjhtiQhtpAcPk2Kb1cYfAvcbAQpSxurRTHgC/+M2NGzclwb8l9YrwH1TXVT+g1
mtS4OW9c8vDvG7B/TQV2mK9g03X0IJ72JHdWPpJ2e1rk3RzZNL1nsUFawL1m4MCA
n3/+6iX/mccy5xOZMv+YNMp863iWsV5aCZ9z1nCDbHUjwVI3uTQWQsNrpkgh/Hfv
1R9U3qpaumTFnDL92vjSu88cTHG1R1BO2JLq/RTfT+fSYFKe6uFXPy9xaeiP4TB1
GJ6mBQmvJaJavo8CqpUnaSh13oDCU1H5mEuJQ4wOLKDCcod7JeUTHXIDK2AHvs7+
H6bXA9+5/8NIXYF4QvHuYbrIKp4gZi2BhNA6YANtGjWHkLbTBfyiBpBjGukcBzvV
7YK9Jmw+Ao9QJINqQArFzWNfsjWbhHusp727VWPPvLyCTCv92LyuB0hJZbDI6SY3
oTNbU95dSwr9bNGYQpB2rNcOAl+NuFC0TAEJ2DOQlMznKImBtxwEwSNaJdHPNfKd
ZD6y6ACpGfuBlEnnly1uxoAX0E+6Irf/FbKXqI2me4qsvDHaXsk5oJOrYy7JGsXR
tIrV8HAj+EFaaVeJ/HSjZPRnEr6Mdn3kt3sstj8ikRzNxoev3a2ezB/bVkA5W1SQ
9/dl9MV+dESvAlqlUxA8h7m4zWyv+dg0Rm3+r8GWuWks2wTpwwn3lbVBxK05iD2N
vkVhziPERxXTkHMCxBaNCVGyBvMoCr2oW6oWsGvQtQsBuM0tlfZMMcHK1c7jM1Tl
MsJMYh66CfTJ/8DSmYT+ItnJ8MYznK0j9kJI1BVVBPAMSOv9ozQE+vwyqlq4GRpD
ap0H3jYdQyMACOWZ/ClhgwzxaKqoR9ygFnhHgxfjdR2BHIByG9kl6+mX3e/tvNFm
vtolPosOegmf4d+pl9Yai1iMPjAumL8I0SMvI7wn1tUvnonzaO3lzgaxXniNeRFC
/0hB/PmSo+Oaw7s+MxtbonDorsY1gyoSWGLcP+SqDTd+uwct+u1GvSKxbdzGnTlV
zTHtiiPeylOgZIAIkXp9uzVwpFge3TF+W4PTEBFk9zYSq1RUYiBPgtUpOWQ/itaq
qdb+qWSfQdIxXBDIQcInP5CK2fZsQKAvLTo1+VFbChy8Jbxyl1BmF/2WaBFFr0o2
q85EVVmXWDTeEKnGLAi8y6cIuvfNH0l/4eLq4UKM71IO1m7ikjCvhmN8+ginvGI/
XX09R9GjAbVRqOhvRKOl0+zZyMhat/9kv3UqEr7cVCRAoyMJEOb4Mh3wqTsfqmap
x8Nr4dZr1p2HApZY3kI9HbptUNLCPnwVJozqh5+l2fbbw7bzBH/Yg6zZKCeMJq+p
bJPGkDcJDIPS8Y4Kb4YcD9grH20Z0fSolWtyh2dVuP6kWhEjUmhjPluvm8EGlgD/
Q80g8ehFe6r1EKanCxr2CAXbRlyd5VIXjgXmS4BamLBIAMfQAZ9lhBdZUAb7D2vO
9exDl3xoifOCuxjexIfG/Bfnh81w3+bIQ6J2L3cyUVHkFxaupwSS5EgmlpDJx4st
5MEMUmYLV5xU2yvYAmcZPc9YA/GOqdwySyolV+uMEm6pr030W/aYa+Yzn+bHK/23
/eihyMfikIixbdtb0jEyoqDF4PCAie6M4RLRDd93unWBcRogDm+ogLkdnFBwvnE5
EGzy/7ZGGXWz0J62/ZsXFsDvvzICgXWj5enFm9x1Qzs1gtXqQJAHDrDCtLjSrz46
t7R28SRnT00UvD+e96YBXJp5zpspp6W0hRTAmfEgzFf+FiqzZzVMiGziyXDr6EhU
k1KnB+bK1ixJecYVGg+nUKG/pQvgVsVvpsdbfJ/asZ7z6gze3hijxdpQHBf0Eo1D
JjIG6uAm6MJLUaWkil7IBvBT0IqviyCOKcDgMSLEEqa1WfwQKH633rkBjLo38NKF
AW1tzJBkgdWhIEQucTLQT/Rax9h/h55scLJFHR2NEIcFuZWl4mKjdFF69vSWgQy0
F0lD/q/R27cDxXktJl8u5T0jebvFMtzY7q3O5I6CyHqpFSCu99AHIhcV8rxXFXii
hldAsLGYJWjjAknutZqrL33lwdyf4tnlR2uHSk3DhNNLGkz3xnN+3SyzZpryPCWh
CAc1g1ZE+j7qmAwbPEUDS7bljcOF1SDYmlo7oFf43J7cfNhfAdcfqZk6ehe0M9q4
8s1goE/l+4wuDXXnz/ReCczpEWIpXZpn2e3qTVQy+M8FggEgdFvkjNGSFaFYGEgd
ABzZRC+FdmSLqIVIixYSrRwe1nILBm5OJmdKiwuVJgjcLSE5n6EMHlgknohohcRK
0tFmqgJToL14QpQEsCwrphpAM0koQaO8CZP1MLobenFoDYMYoJ3vpDgcXSIrwjsI
vAxXERCbdz7TQ9c6hX+PQbgnlVfvzSFzuhAsMLHwLLF5T0TPVxYBhCuPk9/dKU4Y
RpkTWm+68xCib2uX3eKes4P5RplGY+plvLSNFV611o4rXB8ZkOVFxmVsE4fIyn4j
w5psgdne1PyjZ5lx3F/wUZjP6Pl2ZGWLphE0wMohN5LCw13cgIsIhLT5HtWsO46f
g95YfOmF7l1AU+PZ5NlBWz57ZBoShJuwqBmeA11Yy8Bo05F9qVWZqNKG0rOUpqVq
N6f2RVsLsmvjM3/95pz872qDFW20t36Apeseq1JLLLVRzBnpmoRpgTpcgeGYD/vB
ktyVlXjCk+cIEeTVWsfXwYA3lMNYEW/+ZQ1PIWttw4o9NrhxXMavkPp0Ds42ra47
/CANt3ZN6souvgTTIE9IdD8DEjAA9npNA+tGXXHFwYQtMFZXSUV/PuOMmWvWLBWQ
hnBjQgojzEJalZxl0m/CFfGQKRaQKcJvhQXS1+q49Ll/oG5423cMVk7bmTml+hPR
LmBiHh6mbpX5Zq+ot2cUlI4dq++aYFDRJVZLjlWm0NhM7ob5NE0XBzCfzJqcKmvq
Np1P43PQd0xF+FzHIjsZULCOpgWxRni/qzPLPfT5GcsD3lniCdYs8nJUUfdg1q1i
QMbkw9MhEJnh3npLIZI7uN9h6wBndLAiZVNFNYCla7uqm/zRXiE3Uypa4JKfEsYs
0zRn0TAGKCPlqZOtQWwUzCKBne2oMymaKB8zepbyxjI65bGtKj/VZ+vpMxVCvfxU
bDF8Ze+0RIMRQMMwA/eUshenast1DR1ylXl0n6Iy902eRxXUshcDfIh+HvfhaeMv
h0zcIcb+wA2SiaIGtB3435vsturpZGGdrSGPKHaOizZSULRs+HM+OXu2E8VYQ713
F2TOlJrzdFq0O7Z845DxHgd6NVcjEXoDmFDuourWfW7q50C4nj9j4h+4mwr+BZJQ
xxbpTv6cxB3zXgIXkguIqc3DB++fDDDUqST0AJbp3BMdttRQH69718fbapzsw6ZZ
FEzzduTutiupZhqYGzJIwNE5CLLaZdsbeE5f+mrkHOrcy9k9xqNZRUhMo+83QzV5
UAzYpO9s+twSSounR1mmfcOL+l5n8nWAV73hFrLLjbFatdZnDRGWbKzaFm8aqBX+
WADQAwEtDUCCT9HKGKYzu2Xmp3h1OOWB81+l+Okbb+dYJKFDH3YioRJzaF+9mR1L
WymgEtVBCw5iDvxwHEls1qAG0IIUacQiVU7RcQvPSpqg/wXhebgiFdj6cKLjEu07
DbaV6fTDpKJAqgvnoF8YLt4HOfCDIA55h6U0dzx4igxDJhVQ3/0cJQZ0jimLH5F2
deaS/bbtg7+vUQ6bI6tt0qWia5LoiKfaCTIDuptVRjOZV8TZzbJg423yykBezUPA
VgRLQnR/pQeTEgwPTA/FRYXVoLlQf/fzq0Z4geOty52hJ2enqz93BdQ5/Bd1h0oH
cvP1Qd10suGYZrRFxFgg1+JLDvi3qM6gJPkLJr+Zg1TK7aM/LZANX5C/lmMn8nt5
02Q/ZUuhlzjdD2nZOqNlPT5KOEf9hFIAV1BrkrNZ9LdITgeckLm4b4Y32sUp/Rom
kb/H24GUsCnSh5U+Q395/JrZCVS6aCTKq9cpZKxyixbGxWvEno/wPw/kYh56JiUr
8kj041mQF8q3UjCXEv7N6z5T2i3W9TqH4zcucpqPErOjXPItcVJtZlCq8lFnDNXh
l/nVpdJCCGLhFDk5w1OYA09UgCaJjwqEUGUQ4IOUxDOErIabhtqDSnDKnh41XZbP
yPv7Y0Ne2uR1iVwIQmQFj9K7iV2PuQ1Zt+mMpY+8Tvrp4XUkoa4PnwNnPBweEMEg
AVcf2+CFiEbCKknIizPOj15esHp/pKdnHotewNoVOhTGD9Asb4kGxhGHmZlQQJw7
tFYioPsd4+aoL63N/VTNO24q3IFU9exPrVMLM2YhbTHOaI9hIoYtPV9hGUrASEFn
GgC/xGo272V6BiJHIJvnIS9odxa5acY83mAlD5zgWajy6B4taeVckSxCwhFaN73K
EvqNQxweBJfjjgdpuroRXfG133pr4ABV6Uy1pXDHszPap08eg+cF+YR5r+8fASIN
X7VTNi/9YGOxk/SSkaTCcBOftoRmua9JDv/MggKPA6QT9MgTUcHH3xof6sOTZUeI
FlDoB/1XMb7gdVzqluq1XgvV8FFRNqQbfwGaqMuKe3rPvaGlnx7+hBujBXpgkqKo
Jvsd0mTArgsZf0RRUMbaf5L/ckG+vlfLJ3e7ZW/QUZWrfGp8/U9QM4sEep7wLasK
AG11pjCwChV+aRXCpRPWRbpfs5ceYscGtr6PQve0/J3Oy0uBsbecygulix2yOC27
SApt2NrJ+JbSUQ8opoKhjLCLnWQB8LZ+uEwXE/mf1WSHbu8G0YCL2e95sFwFjV9y
5Yvucqz6L+sq8UNmwVjVMQnYtXURVPaWfj0sx21iHY4G3ArMqKeX4nXS1GyRoY83
c8B2OyxHe83RSC4wuuXquzQQodLSx1VQ3CE0qgUr1GpweCuN63g18h/71JjgbZY7
zNlZ2HLcyzRyVpS87bq1XxXgKO80ChidxvEilTweeYLejpjbpfSIUGIMmruAk0SF
bCJxipe6ZQ6Sif1cWbtxOUFLzZgdJYBzdDM89Q3HgugSwgOrtFwSZjxNujFOt0ok
SB1Tag+b45x8LSnGUftZHqtlbW8N5HbfN/a6FEzJ6sAN4dRP+UX9uRQhIuyh9udz
Y9loZVPW/AWETENrwpuOBSFhk3VB5M8b1+phF/N2RK9EnnYcmDwkBnx+psR/9OH1
SJ5DYtf20p/eILYG5B3jvgnY1fTU4wwVzwxsOqEiwhlMDrNXxnimjZodxmvh0qcd
vVSAUclIR2hFI0nNTjD3jVy8lvd09o1tRGy0GenTnBNGPlkbMtyV1L17LchGUZaq
7DARWgQWg4MGViNaqrXen59KnbgAt0rX72AoZ0Z8Fyf0j/Mvtg4eN0Ovjgwb+qOs
Z3WOTTeAnzj8ERdz2QW9apOghvQBXmvLpGibv/Z9/jTndcgSlhrZJhotJom74zUZ
mXQxgYjx72TAnkz3+uJIudEQpYH9gkrvmGsUkWPXnv4snNtGGc0WTg007Ho+eeC5
1PEoE71NdV+jI13XOXzN9G/RSo58ZUSyVaykf1PnWU9I8FlKH4wwipD9Xh8mEWBk
s9tfgKQwTbzilxGSPQdIlRqGdxcnuCLevxoMaj0aFKXe3par7ZYz3kIDyP/wZhy5
SfPhH1YZLD0EkyyUgjnjDkHAcHX9u+0ffCrSuosRo629hm6ux4iz7R15tU40eHOl
XytR+xTSodbMdXSI5NQsIThfIAK3lmEoS1FnfXomOhd42gRNWiLUjsT9AdJpoNXR
hP731f5HOcVkXDwkDNu2JYMS1q2w1scQmi3jdrduNbGihokh33CtzfMoaGypqTtx
lpLcGX2oFAebimYY561xfRDllDxuKPzA+C6NYx6AxOQ2ByP1M2qV1QPf90nm9z7m
p1vhbNID93NqhmTlwfZs61zEQzzVI+PCb7p664HbffultkRMcklSFNDkrSO6kVeV
NArKAc1y/LJi9KmOxbuhNAjDb2vAwgt6dwLQwJd4qIRUZVZcJRTFesa6Yn4KU8wy
BLVsrClFl8vXt89pZMBVUugQV01bDMpkO2RdCEOStnKeCiMnQdZhv9Bh2GbpSIbS
HdZct/06FvWnnkTEgL1MVj4W/E4H9G3Bgacvz6giPjIIhaO+xWPy8rfT9U9F1gUC
DWElg/s1ekb8rL7KCUaJ8dZO955DTzlP/RSJcgah9qrG6qPjobkHzO6p+ZcHNwgR
qf1M9po1qBie96FxXjpzIS3sZxrXW/Ib2mkMp4KWrEH1Y51KxVi4TZRU9zyp1HMM
KVKuVE3jjUBGQ1Q3z40PwLZZY/Dqh7eUkvPH8u8NxECq0KBxmpOMiH2mUJ9XdF5+
JFRMULZVIAmTN8iL1jA+zYPYgwerNM2PGwXocTKNMy1ovfJgnv91dHzYXgdysyOI
FsXVpztU0J6hqv08pqDMT+4SVThnslJaHZbclVe0STqK7Ax810VUvg38hQW3zxYk
spwd9dQ3gL7n/Gegh3u5M7TTU+27QeO1fO5JEOIkXsW/h8szGgOBLAJUX9h0lqMx
Rf/wj6MekgBEJvFMj36oQ2KyXmVM6rxYSXa7xGcREVAbyUdeNUWZYZ1cfjXsWoJD
PlMshc/Xf5rviP5NJ/PpFBwV7h86noRNN9pp06lQcLba0f62RVPeuJAHhgQ/VDqC
a0u5vXgZuf5bYrjZDFojMUkM0gzmvVm8wCKxPp6EbaDDE/vwSwJmQL6Ppnqq6MH1
x79qmttqIu4htYQwX/TXEWndaOOOwggwTUA8pFNzMnpCrfqSrQkYVe2S2I5CNvln
CaBGoF81DZBGWX7gtBww3ODBdgLxSyTnPb2YGoaw9bIoT1AuR4XeL9YuDmzMk2nA
PY/SrRGpl2fkvXywv7NyRH+izea3udl1nfnLpfNFuZtj7em+34s7uC0L8RBjrN+/
Yk1YIMFV+NPOSHhJ5xjcSBn0RK3TICJmv4WkgDp3yrgsAdVq7FJT5MEnhPR7mJGY
wARlNYUE6Rn9sUH3bEtR4OkL75qVJ64tgCxeU0VzX/7sZuAYqHJIeKwqZIyMoptH
GquWWR2nZUpA8GjrygQrzIo/xGH9kTHeuVlLFxVdzm2xm0GL2QsKDk/q2lMbDdnG
Zkzh5ydgpd/jsACA/Dl1DFpk4pwLmRBXulAbl2AsSDlajGuRvan6Wadp0IjFgEWZ
n017CYoaPAqHFv9vDMYpic0JciABWKTF6bQFJz0FFIS7Yww+R89VL0CU8aYz9P05
qrjCiVFqvgNKH0VfZGg2R1stuGsCT806HIKk3g0NDEEZCpFPg5upr6hEOorV6CU/
mdtcfLSadKYliqHFOuWl0tORzAlGCf+H4jOTdy3Fxv2dBHO45uTwHU28CughXuvP
D8WR9ZchSeNx7DZEw4ChvfuhasOHP3s7lKibYZYAFc4oFVb46i9jZqU/peTp4s5y
z+40gG2tr1IrA/yIa2ySyyb9h59ErMDJyMQ3TX2xi3w17NQIIOB4B8B0yQf03Vhr
xDOIsAqmoCOFOPYS5mac8pDjvnMLr7Nuesb76YnwMHQedTngMpiPVBTgHo5CNeqH
91FTwfuBX7rGUWiZi9lhjSv0Dfy+Pi5g8xu/8wmY5W0pfPTcGB8pyRUThQhUJnQE
C+V4aZrKnhPOaxHNhJNoIlqIN0A+qyEAaFHZ1Z08GpeM38SrASx91PPPQUk/XqJX
haQA559u4HxLeen8pd2itQV+23fWUT3FPmR6YXesn0nnTWKVROh3aIdVY+c8XuoW
XahAd5sy1Vz4s3wSwdLb6yMPx/JckbOHxdSOKYktB2sS8xYWeFsGSwYEbLjlFcpV
pjsrJBFf4CuXIFs/c0QX1hT/55OyAqJPwdB5oYlYDs7mO0OL0k6KvNe0MgnF9/F7
u1kDW5rV2QOufWaHCR07hJHh6WnEe9qhyb7KI/LT2wXBCD0NjZ/TsfM4fzIavF2E
M2qqNlIEA194pUAH1bT0A0CxClI86+sWu5kKDkRt9icWHm6SqRyYPtZuYmDjIvW6
yQIzAzQARwIwbwjGd4RQ+6L3uF3Xcr4RTGDrMGNLxjF1LbJoP7X/js3jDmXQIdb4
zg20ndEgs4YjYVF2MjFdefCG65FpEEhd6YS9kIOGTAtef+IqtIQn9aQSga7YcTCK
5Nq6Vgtu6tL/DCVt0D6XDVCQ8EC3r+veYv+Be26rWYQ6P/p/+G3t98DS/kFwZ0id
yCM3Jl3JqRZuYGbMyoXkHuDMvR8Q4nwV7ipancHzUUVvK0xMtCp63YVnyz76ucf2
cc7cFW0bGRFMtQjxrbwLWUI1DBLIIlujs3e/zAg85Sua+KCwxTjchyK7MBBap542
roJWTpI9ofoRpWHpsVWOqJG1gXgkTWyHZ87qQ5GBFB12cEwIMH64zGVz3+Hbwnw/
TEbX10zdatUa0rJKrnk5FcO8HvluUaOY3xyYAitruOheGXTid/nes1eiUkDZdcAK
eYoir5RzDppE3DsQrXQGDMhR6mnB1QCNCkc1mXK2gMzCMAnReo+AO+wTfDsJ/pyj
ZhAMpG/toinM2n9Mk0j+YmrYZKr1xPFFu2e4G74D67FBn7v2ywRTCec/V20tWszo
459yoiQVhV3oJB9G75s5r2Sga6nuv8vjkAUlKxrQ6qqtG++NsykO6Q9WeBbu8vp+
Id8G3wwcj6XyekxvYRcvNvHxgY33boI7gAwOOYl4V0hvmKQl05PHBN5+a5eyKW9v
5Df+QaRdcWqxiBQWzDWFv3MM8JDpPScl1JiHW+VV8J81GGEGpC+N5aXQKtP7suPA
ChC/vLa2o8NpmvQk0QmK2NggDD8rOGtZZ3axahP/xuuU4XqiHi0enUGbWWrQlqiS
EDNHLvfBejym3oYRxilaCxqgGI4EwGpUX9M1136CMzIcLtdc3gInjjspyPR7DAcy
TPZ5Nxm0K5xhsRVzleXRV2adpC4yAGMHhPWB3ene7yN+8+SchSEV3TVD8Flln+ls
qO980xVY4tHP16zoVKqGD1Ch5KPpyEPZVcKRjnmu+R2q8rTp2fw6PvkEp6K0VEk5
vdtgsg2d6P4E3ZBSNLckWsJnVRQXHBqkmG6Q4ZgQ7aOogcgtxYtCUf2eqT71L9tC
YMm8sUNoBW+L1vR6B5ETo+T1x3sPu7z1hA47zG0XeANSBNZLNTb35fuYH+YsullS
gTCpcQJyAU0EMmOSzcHdmuCstHMh92Od1jhBDTCip38bMT0HU5H1+69RiwXY4WBs
d7G0m9hRq0zBLL6mMpGVNQCuAj4OGFgpJlvUWUrqBhOEnoTmAvp5az89PDWqTqzN
f1E+RAcmA2VeVCuwr+tIdoJIukdomnKqEV1nNX6AYfxBN1T3MP9QxZUuth5iUike
ynV3vuagLG/GxlRbYP1jOKugiXSPBE/3l+VVSL6zuJ2B4yDzX7AVbWiV9tQljom3
yrcwJwq0p5dc9Eri2KKVj7Nsf2S1NhlPYjc9aCjYmdq/gjaJXd0aJNVJkCoQogIt
pa775Lh9G9BuX7BU5ptkkkoF80xZ6ju4w6pbf7r2KCv+NWk3llqKw5LxA0VldOPX
M/BNS+y2gQdLckmwLFd/ZTU7NqhHvhA0aB94LdcBsYeOhI0LEfm3XeFHA0JXin/y
9WaM04IUFkJLx55o2wU3TeXkYEeKuhxQ8FPWGqc8mN6CHTgqcSIFt5dNGBGnn3Xu
JeBbWnOR2KsQqIHVqq+uFe2dpiTqyF19+zucwAfuSpwFcvDLtv+n+wr++i0GPoFU
xCnfnceRR7J1StxYtBsb6IOL6NgGNY23JR5gux8/jDyWEAhlQ2KMwjChwa6L6KNR
97RRpi5orh3nsGGnTlv2OQFFkARADl6IKsslWajFLMBM8anKYPgKbKDOkyqazpB6
39bPRiwrZVRzkfgjF09xPjxdrLWCEOc3MyhtQJwEkANnmnvwe72J3I89LLzCAyYL
pGpQflWudQ8N1R3KQTBJ5YEyEG4I/6+7HJBOcQ8HeuVy2tGRRMQRb6zL0fD8auop
+CBI6Sq05Djt4a6NNyOxMEZPiH+YkVwNtnonaUHr2tXotq6YVegeGVDOF30wPvtB
sDGumYwKHUccO7++05rFbGJg7RaP2GF4gbexnnzh+BTDOYYrGOcXuhBWIl0bG+Zb
r7wuRj5SmzVEAP4NHnRPOtgARIPXPV1V479PQKLQldo8O5P8Adwu/EXb1S9/+hYI
yziWJ2J81q96sIMwmUW6TY8inhGQXab3/qwvU2t98dtvI4kRLXxzZVsvF1vqdLzr
laEDAGWb//d9BLR0hsyqhvLL1HqtheenJwWTqR/fXSKxGdMITNPfXVce/5M25nlV
esK/aBA9gBKKLCGk2l95nsgb/wSxf3Wnhfg8m6jgqKEpmTiKoDlKK1e+GNxY8EcO
fmm/gdFcm/wK+/nCuwD9sRtHVPedRCj/bZoTEOygCPw7G167s529Jl5kLSqRtiuq
EMhvDx2tKBantKa6IW1kG4GfCCAJf1+0G5riXlAKEr5Qq6QjTU7zLvWoOdK6Y3ht
Ylz8GBPaTzmIeP/jy2HTKS0vQjLEHlNPjhdiTuL8gqG6OcfgR1w8BItDr4yOr8ef
qP/uKu50Y1EqNcgV34uc1SZF643v7vQsWlhEcNCPnvR7VgUAkzvK0dddv5Xdi4on
FdjKp4XFg/l4SJVI9ujVMWo4Qh0+po9Ing6C3ivY9//RXpUTsVOXWV8UOphlqZYi
ge8LFrXKk6E66luHa2yhRaXfNVMFwVJCfFXCSr/qejgyKjDufVZ7cftCXdaNFr7L
tpjpjy5+PqoeQCVis0ztV+mKXN0VbZ7tHijat1YA5zN31fO1pyh3jNLhwpxvBcbZ
XIuK9I4vjQH9QiG1kYc1mfcS61PXWkLjgrRRfBTf0qipwbFRbBH4yYXc+YZq3ZDS
IIiJcjGTHUv2b9MXV3OG9CA5Bi4JOkH4M4t0ZmAu5ycFWfpdXg9UIjQyM58tMSYr
0lOjg/CcUyPC3iJrB30GG/7j4U98WgjmTBZ/t+wVh00HDh4Uy9U7BIv9vm/I0888
izD/5iOrDuhCTyDcuPPyV1RNhI2RCf7WuFz4wf3lQtQ4Y4lLqQqGRvtvpWg0TmNa
t0qEBEInPIQeud07OQoX2EY73xZLTXR9P4TU9/fSB31gkoTz0O58JmfXScf1LNEj
JLkNKbLaKCQKmVxwFnQ/W9I3R3qOVyL/Pl3NvlDNut5mFg8R3vW9Un5HENkeMpWX
ddS9ML9lfOTQyl9zWOXwVlv0DP35KfR9/ieo/XuELKMQ2D/THv/Hd4cLK+zKsDCe
eYRi2ojxRo6OqeFppwb+A2iukmaHkBMoo4kRnHVUXnWtGRV/0Jgxyabj2heAhNw7
VcHlAcir8TyzjJ+z0LOZaleFe3nGiIa+obdTdxlOp83JM6xbtRTiksfaiRAwxYU/
2FGl9h0vnQGavawoBwxVt8yyqlpkNDb6xxiyIl9zEWHS32Qpn10PfJL/zU3aNf7A
pDSS1QWQJq/Vwph52FCJhhINU/JpKWpwqugu96dACYVE8q0HROcs1cccjvrMhmxU
Umbuydp9zlVg1JcvD6KqAj0AbpoIvFY7ES1jL89TSwMpegPViOaJ85xxnv2T9qgb
p8uWkJk87UccibZGNjUsI2yaPrmmJmyJ7TO2A3yC/J+Wu0mWZkz9wGpKgdy8qyuo
98aculhV1mIxf9/qDzitHt+osoujI58eFO6ifnUWIzeqej2MGpnDDT0JWU7BqBjo
Uhh4x2G5HgG19ajt1tLu8iIeWmv0FKnu5te+5sixSJQWDqABXzhM58bT1AxCpafw
vlfUUIZBRwqgZGiZUP4lI+gUnYgpM5MRstoCSnypHY/aF2avoDKsc6RNaTxWe5PQ
G8IVtYytYh+rVTzJsrxlur4a5t8T1U99uIGOWVZFmCyP+UGbEQm94rH9vfNCJm3u
KDt+4OGbIXSpwDhOOYhWQeaAa0fMk+g5RP/Dn4OKwRVqy3qz0ihII5wI9QBJV4a4
J/Tf27qwr6gY+yAAeCT5dKeidIfRdahOBBWOFrac8jtM9y9qg3edBiHYuDV1z5ds
a0wOetIE4/ggICvaRY2kXogVJTNUNlucd7uX87A694UWRm8spQNqswhyWLiAQci+
HkoObl5XNPsEJCFi+IvzlMVBS6lSkU5mfyPKgvFvo/m/77jVEnIIDRaLzzsSsEcR
EoECeL/GL7vthwAlKwMCC40gMZzSuns+qD8Hfu3mBkdJhp570GpbqpMP/c6m0WmJ
2gSGbyzDX37UMsg0U5DEds2KsmWXKzJWoR5FU386EcH5KovYsBcu1jQ4LmC7rpnu
Rh40Hr+IE7F4YJ1+bDLk1PZQ3lleopg2DgEggg79a8GLdO/ykmiuNbt0Zg8OjEdu
U6f8tiCFXGlbknIc0vO0t8V9BIddoyIuRDCmzJK2QVkRsZYRTyyEYs8g45TJd/fI
w5QAGo8e4I0A1rz/jfmbAEyhePz/dSvHQ0jLZU8V2GsiPwWwsUWp9H2/j6mcvgrZ
tj6BgDHWBAmVKi5JtnIeExOvyuySoTLBM0gyznM+XdhsBP6vi0tTZTYHCnE2a73Y
8zODrJiTGMcCG8bZqWRyUVYg9lJbD65AJ73NsRxRWFcsVbgvwas93UIQPUmuJe7A
sHNsL83L6YF7YVmXkEw9u3ndFYF29wpqldgdwvLeVPZ4YC1XKpDa1rjcFyjMMi9+
FejVRUvR4t7X9WwbWF005MNlAHaYB8ful99XkMDT75/SqvQ4SVac0wGXqeoNfkp8
IHG8Fs3bTM3ul3JvDLjXMMypuugIpFD0oLK1IIC1PGqCeR92lfaSiP7AlNZ9MBcb
vWgzhM5XY7cpfPgDlcSrSoulQ0rnNfuzWoaEsdIK/ikiXDqrdT4xvVEuPS0RpJ1z
u6kStig30QchwO6ykCvTppnEyAqM025WyWLRCy4XkvaalYkmqC28HaSt5KkK5XPj
y3Wz409uJc98gXloPxGhVQwCAoKeEwySDUehUyDdn8dqO3S+syQ18i8BU7KVcC+8
A3K72IGhpwIKrYoItxqS1DXUIq6hYiyhUIa2yPa6qsiimNL1pDUSwCnWLaW/poUW
XwoGS+jvzMwZz5SPYG3uZcDECe3G/dmzrkmMRPyPSjW8YPJ2feSDXmlpajbtQaxx
Nw5UdHcv6hUABQecktsHDlynNW1jL2fy/l6xKyTR11tFv9FhMpHgPzEsW9yeH1Lf
bsWq6ztnxzHdHcFoy3J4PoS6B/3RmBqEobKohFHwpw/gzPMiHBTbE5RS2ZywMUhM
vLpeR/nOTUg3UZ4OCV0Qp47mMbQxZtB+RGV/GcqzNg2EhUhdFsvsr2obs9jJGa3i
OIT1IjnRFLOh8f3Z2cN+AjozBrcCXmqCQBlaT+IyhbRI3ey7whwlch2YC85pFPov
6HzlvXULf91Raaqw1h+2u389bUxnPdvVH+/DZGwitZAf+2/1slWp5einFDctx6J6
1WSnu4unq1xQc8HUxBAx84JhTNGJux8Yqq+Mj8j1UEm+Acb19M7BRwJmteFUfSWd
HcfjIt7Wcui3EYKGVogVImZr3xudjL1wMRF42sbyOON1Ox8DY4EYoeqYXb/w3pid
Ityw6DXB6p3BQEmxUlO4A46P05lsCU92rrD1cxD6bsml2x6mPFS0McuMafqp8mby
+MWyRHh/rCXIuzOIWWYe0uFsI2aW9TlU+7dlNYkWXVA8BA2JH1reIpBW9jizKmqe
JPa4iAbnIBjtnR2T0bna8ZJe3tvqeAdGfo5h2BxeiCjyA7N1eqLW63TCdahdvK2T
Vc0exKTWGE/3Xmj0WAM2R+Yzly+1+FarrfZdHs2KEpJ2pm8LwbYv7rktvrLtb0s7
bbSIyszvfSbHwGdyKp2526d0q8/Z+YsR/yM6qxQxH0MnuTNXcK7AcMz9J6eydXj7
TX+OlRXjAKOpXAXPt2mz9EjVQwrS5FXSj/GQ82Ak9he54pJRuzNkrxo0Z9Ugl9zj
+f+WjyfVfrPCYLFSZVZJ6byvsABUZJdbSqM78M/P/8g0Fxe1mO6RraXSD0xOUtU/
0N8duZeJAcIf2KOnIlNjgD9wbK+ZPKuxL0TlvXrjFzH6bR7gvLnCYW3X3Zic4cug
HhXjW3r3WRxnt9+tQolMc6crTJVjdbQbUng3c+oCUUpY/KryXiA95DlUER19E9gn
6Lhfuw1iGxqp7mSjdon+M6+KH2IVd0N4hheYlE3YHboF+RI8Jzq0q/drmMvk3AaJ
RQyRgtYnRoGD1rJW7VGcnxpJ25Yq9ZNRsN2P+97iPiv/Fd1Fh0eH5kRSb+It8zbk
G6yZ1J7CLtqPHV2hJV+Adqs6f6YKpCWO7Yn2gjqxFqJucbQG0TXZ6uz/4pBc3ZW5
ZThJnk5oJY5vOjduTk4NyN6WPXthI1vGpGR9gQvKq04AmVMXLb7FNWVpFIJglq37
LjePWFLfYDCQZMz6rqvP6AHwRP9YIW8oMvA6TVAI9B0bC8Q0T3FDaCCbtxm2gXIT
dQcsRZUdjEnK97s6TydHz1t6cERZJ4g+8Ql7nVkZlVBjuc+Ejow9FjcBRQkmBUms
AvcFJrRZmKfLdtsZEB93YfaJjm6bLXkO4A6IKeRJ1ITtuaUX5rgu/IhsZ2386nAO
8/78/Xlxwye9xQ8j2wfjIEwqlk8g4Ulo+cPLweti77Ntn+S0CPM6qABdh6oOXXc6
ngD0eylOANWgLFqlsXXHIRp2jewUmVVhtNUnSY6bEjXmUQcZtGZefNxekvbSsKPw
ITjI+nLw3Bn3dlqdHdGXbApFLnHyayjPchuk0jayk5zk37nq/3fwwUYpjxewtaax
W3S6fGod8lv6EJF4RtlEUn8myL6gzomDoBFsEzs4sk5kJFK2gtEJ40VbTrd9Lzke
Gyq1mIHB4fsnjV0SvKXfes2Ij12lbd5V2N9mo7bhc9HQ472EuHqnZLKd43J0vPfC
OvW7q7B2orLEQB0LaTMfjt3oCYkIWb7bfLpPJWbP2pD/x6qdFZESAmqLuOGiLJVL
aqtlmu/6khw/eGhezOpNXvdBc26HPzMDZE9VVFemYxgTK+N73L/U3MOCJdG5y2w+
EKYeC386eO+vLg7BaOWBn5e65qxLP9BCjsnt77ucfDor9dRlSzyWEjBfgV1YqMrg
+EcqxvlDPqR1fVFUIr9jdQt4zqtuFWwIiUHpRdO93epE+txXsoIhLq8ph7efM59x
d1RUTEHThm57lCRNwoauRPqvS8oRxUcs7RHHbo2oK40lsNGEDerFcdxGoGbsmuBi
erYFmT/Q4sbsRD3oqSKZL/xsdod10dy8nWe4o8cAsmHBFnzzSHH7Ona6sPGpNO/W
fWODpqLvKXUbF/AogGq++rYkZxwvUbry/1RgF+zAH9lYX7uAM01B3mDxJjzvXETo
A1oTRCLSsVvNhhYnLXfhUbxafGAchpXfNtRXDF6AD+CaKz+BL9stmpJ5pxRO4q9B
9jEAWtT6ouMN909mxB9snIi0o9KJ7ZHvGLNOCD4ikfCSBYvsqWZdlQ6CM/6kq9li
KVQ/nfPDcHBpsjk9J9lQHSQAioVJMtcXjhjNUERuzCm8Hyz76M6jdFRTphnX3xwG
WItZEl7vlok/0J9Hwh6jMuScIS5UlXmyoCBqQybKnwG0I9WWT75TghcZcoH4QrlM
iB6XH/FgSCS2Lmd65T0v4UWtsEcn+dvjc13uIVz/7Q1DK7jJ24gmlT0Fa9B2zREr
GUKnnFkfmIzlinugiRS6pmlHATvRwJ/y2lk7llsmTbIJAl0hFlL8P6AOGLBFGuJK
rKcmB34c8w4S732LtpspZV4JBKg6KhV/k+sj2mpZWlb/q4Wr9nWUW5mxzb8cy06e
tk3LybK36nBfnAwLYOEdP2OJUgQ5UygCiLH8Y5TIQkw85s/o2QORTFduX6VqF+l2
+Na4mVePyJWICv7YzYw0XMG0BZRVsju14OA1NX77KsuCHsJ3YdIYYPLBRsaXB6+8
P7DWIMRNiyskjfeG4kYy3X7eJQiQlKpwt2Ok/FaQvww9OTXKWnPGutme4V8FvYpM
waldFW0tqhdRrUI9enPgEHSi5Uhhhlxv2ywDTpT0Cg6URF8IW2YtE+OePxrxpuD3
RIdOkNbE+9HIRMntNHLowEhPHCTgypNf0l6LOgZuaQW/eajE7PQ4ZJ4fbhfaFMUD
ToMXweO3FRuCtmUmQJxiSB8yDP87m6ifyVwjgce7jMCjcpWKPDYvPvYUlnQIXziC
KiE5GzVbBfVmgOCTV0WIPCAK/qdERPsTxQX7F0smCzyF14a9b4V1gEnEhU4tqQWM
DPbVhN178RSnjC728UIEZ6wtxLOJAii/15xV1d6+GClDyS8a79ehppG4iCK8y60I
Bc8OYJvncvYFeXdHgLmfGw1OfDQzLw0LUkO/HYsTEpOO2tTB058ZSDnat8/4ZAX/
HTTDH/zchLwYuo/5NzvT6d0ItxhdaTeYMLMhCeBMN6ZmhPehzPx2wWcYF0kEacgV
ucRxOCYNhG6reufuHGIfdcVJpIbYHA4IcaLWxJM6D9HLDBC2OUXESFkpBMmCs6eY
q4V4xFr7ZldkSiC8VrZl0cJgjuCMWZ5ifL/LkUVgM3hToIJL9kKP56QiO/UnIz2p
nqbyoGTtGAB5hxzIJ+wYra9FyH/aR09oo0s6Ex8sqGJ4QO3eOkmNemmd15kZ76cW
XhdlQFLSIZm5zXrdTW7eC+TzxAUoBGfCIhVZ73rjmzpPygnR00SrmLiguX1lUike
RIUC9ALypTVeVTQD7PRcVuZ2Enk3vWyvTM7LLusnvrQKsALsD+l9NpqoOq/ttGr5
ac33zIxBK1eLQKzT7/MRL0dFzv9it96aPOxyoGs4+toFPJsM1T83YZG6E2sYXbrL
0OMH1laLRg9pet2KbrisjK2lLi8YMbiw3+CfmW6Et10+M7eTcnyPlZdeqGnfU9b3
qnXRKjKiVL/dkl61q7dBzT6cyQTCOgB1ET3Idz+7gA12Noo244wqK5mY0HZU20cx
zDSrtYqrY6CEl9vy9W5H5rcJ4XIqly9ty4oK4rPw0iw2yxA3l1wUY40rdI53CnBf
0CRxVd9kSYkq+bGkcZjQxx82UAjfoG4fjOABhF9JHLDMsOORpZV7EXCzrb8wKCcb
/nmXs9MVxSIh7gu/3UUA2sbLtc0M80e6GATdrEHgC/TVWZBujnzlbhvniQVCSRsE
TszdHSefGHBsXL9097sNYZJkfRAEoWHjq2e+yzKeG7JZ5mwJCMlJZ0YR0XPoe5SJ
5ez2pi+ENiTIj5PN3tkHGJlqeCIwYxvv2+gCCYuCOTD+mrwfXNtS5T1ZT3IdrxwN
FCLE71IpUEeCt0YrqZn1fdJIR/HwbQEk7vW3phVM5zFRjPoKncfGo3kwLHWAS0d8
LhWxQJjoQeZrhlIB37CsLrsKfh7grAVN8o8I5hHH7JTvVwT0hvH7tIY7BJASLLA5
NHaG1YfGy/mWAaP+53ey6dCuI0Ej/jxHPAC2ThBY2a8Ewq4TCRMeNafo5QTVD/HW
gNdQ/Gz/2SWyeBxrxVbpq5oXV0CcMVymWbyynNpdBWkVwHN2XPmCzNvyJ3YLEqT1
wWfjNKTpSVD1pmSIRshlxTZ8qXwLkEEsB/smRk9VlFi7sa4umcl23nHgo3SgUaUL
09G2eJCXcQsRtiyL22CZfJVNHMXgcte44JjwyyQBCKkKDqzomHG+EnXTWyjex4Gf
DgOW5voo02frftWxTEiFbdV4G/FaeinCmJuOBcyqdw62MqsZZUqO1YORQW6D+O6g
ObnjHFZdbx8aDB4JoHlhdN8SqHXwe/vXqQQjWnhb5XFnEnjNjdQFMJlh5rvJYQMp
uCh1WGtQbYqEx5vxa8+gtII2Zpbe9ANZqGhUqge8nadSF1m9GCVe8Zon1Lez2egS
X7Je+QDeYBfa44ggwssUC0ifx0l58z8OU00/djlwtpAD+OkaTBEX43Nl9swrhUr9
JvadvBsfDgKLMrFGNbce+cDVaFTdVGjzaQTr9YfwO0p6CJHiknnmhWaaNgvwn/RJ
NVyaJeu3+qMYDB4EZ1V7MXc6fH7u50LFUg5GmHi81h+nKJW8O+TV81aZPJobU7eN
ngpC6B/+c3oeehyFVZwbWSot8tBrvMsqAy+Tf9A6foEi8sAN8AHnG/gARspYRfIV
dCceKNr/GKfFeaVgtbQfV9Kb4Q6cEJjherlHbNMxLfCAykiLqiSBhMDv6qDFs8uV
U3OXwCj/ydVE/gueBWaP2J0kghEkw6Q0B2qZErjT9vakbuMPrAD34P87LZLcpD2G
bMlqkxzWiN1Prq5SImNcLHGH84AEvHXwvmpbKf/YDq+/dwM+sc3lwV95qeQCpRtt
cntD2t8UaXwfa/Qsr3oV8YfgDR0u/5FYE7KnFwX9i64tDApFN2m8bvEYXi67dHp9
bYObo2cWMKOqwReqgtLfoO/6w27MlP93ApsCvdhDsbdZFJbn5zC7FhKYbpGcsgBH
1hzo6JB4vByLt7CwOi2L44j2PHfxVQoVw88agSN7RQk4GeeK39dYnY+bn7RC5vIk
5N850l4o2hvOLm9//5HmhfqBeEH+P0HZeXcTKytZWF/mEqsx9JDEzdSHJ4tgOlM4
jmxmKDANXkrbrGUP9cP1kBkjbb8GUgolAlPcOONvtAOfRUKQwpivmVCYGFEL0R1E
lK3hujECiH8IC1JAw8B6orcsOlU0xVugBSeKYCJTxfEAxWXDi5z7EHzTnvpxLzwI
eu6NszKipvdsaLMQFGUtiiudrMBPLNiCQj/YuguPXuHsepj+WiwLzbYZhNqdujOa
FPRiv09Jy8Arp7rq3Yhlmu4vuGdxK9IO8NjLXjKDi9ixeS34z5fTFYg2a7zllMw7
6XpT7jfce9xjYMR8mfX33s2dQB+2J+YC0sV2CrEHvyIoTY+8cJjrFk0U44DlM8ib
4PQxTmMnCovhRJGdLqVgB+wGPeCJjA5H8ywm5b19MhpASNTPl2ROa5QCIzGU0WQT
+jWt1hVYeaRhxEUVspOjiIRHjfscGn3NCxe5kF+sqPt+nS51Mf2EkqQuf/CRRIGv
5HZIurQhvNKmW/k9Nxy50X7cyj8DjFbMFCApUj3EoTpM6slu59FOoVqw5r1NXXyS
JAOivhqb1Za7SwnXFHOdfns+0Dgjnjwr8fGx/MJX26BE8sTq1Oe1PA5BIGqh61bL
KLs0TReHjK7AHwQIsomCEu771K6NJDHdhpmAyDm1n58fPkYsANwY3dc87oXycjDA
yEbWHWZNm1vwE40wySmMNHKkvrAGavJW21L4lgFnMnhF/Zg9l6XQl+HUenyAKw3X
Cjigb3u9le5cDNWkxU8WfJn59YNR1hvbyznY3m4nNI3JK4mS51plIBkD6gMMHwwF
ZMPDxmr3lgFqk55D9gmJoKcsQxa1TU0Ts/9JVCgHC8kVIc+auvp6gSy6ApZHuBrp
154tg2gsPPHjIu61NwPL3jB/qwfD3FwERTw1Q94MNSkwef+7nwKeFpVAbA0wIaMy
kUNajw1+YL1izK90xNCv9VqISQWHeBN8SBCbnVkIXAF7iqbeXS0ir2ELzGOK0Bvg
Xkx1jXIlou606LPGAQG52nkrWTDPKvNmq0zJF9zGPdqRKHzfk+eOPAUgilwXsFCJ
BBcr+QTDzFN5bI2xjQqD08KZRQiCYU5K7qtohI+QeHEg8xjGQjgi0aYxjHTqjMTQ
Cd4teQWLwFTDeENV2k/h0kseQl8e0sxVRc0fAmwADu4zn/Tg6+ftCr8mZQXPQCkJ
Hrossh7K1FtLqq5GYggW9yqjxQdfjAtYIiAm/00vxDUhRUsmFtJiF8QVp27NLcE1
G+nVCEp2nlVSx6QNq5+f4RX/LDRNOmaVjigLuA7J2y9EBuhgN2kjtnraJoxj2+4Z
hn7rBqHZhrs233QrI9nxgkWLJMzebXhO2AMbv8Q2u4TerqzLfLZRkSk2/Lsmhc8p
z50BUvlyHrSulJTdv9psCoe/txkeS9/ZMD2SHOVYIxTr3WZLAAdal2KWliALN1Ml
9msmMZfyMbQMjdODLV55Zd5TudXMy1jfqj9gNAKC5dgBs1gKZi+hXWG6T/FYkxzE
WUq/YBfOQzzUiP43QGFBA5UMz/og+lO1W+huxhgzhz+jNtFOoHIl43aUxsIOWzvS
IuNd0DOL5MTuoVuw03amt7aAHqqX6yDX84xMio7tUB17e1No5xNMpXPC9qdnhm6x
W/GegguLiNMGHbZgfZaM4CUeL5k+ictmz4t/KvaGG9vYUYjIj1I2OBXIjaPe1IWj
z+zBdyiacSUO5ysrj+MeyiARL4r2KIjK9VycrPPp3tmasRe5rTigtqVEeN3l91JJ
LbykUY2+2Ih7zMqV5qAwaB6teH5Ul8uYO0aBk1EkwgrZeEWjwpMiCgwY8DRSN6N1
UuFfmZmVs2aRTUQ9u4aDQrfwEwnRsm9+JReDo2HK5gCCihZ8RARmMHwodAromOmy
cCCtiWErFwPZJRzPMXB40UeutKrSsfsycmvQ+1kfAkJkTNXI7C0XR4fs1+M7xe7D
5PYOVT+pHAPRvpdZgDtTURZt15sg/eBlhQT2Qbdkk3CDViFPO+W6yT3Ns5LqZZAY
1bJ1+9HHM3xRiTfPieo+mkpeLAPnS+3iNwr8mQgp1CeDSoBL/YesCnhNkszRIu1c
VuK0kjzSESqWs8tg+1ReeU5z0mQJsQ459aWMZt6ZceJCDpkG4PCyt3yYn6dQrwB9
DkQX3h+PaE3xG9ROHsAY3EQU+Uh8+R79Wl7xlNWynQ1Yxy7NDa93cuBiqMZkAfqi
4r00vJ1bpH3UAwG9agOh34HmFLe5GhDxJMXaqkA3se618QS7EJ8hxvNOwWkeGVzI
YpbplILdYozFLyl2fPH2SkwDtOcgVeNvy864qQKyGwHsR9ZfAfyKSIEW+oxfZ1ja
Z7KIuHWWIXRiyVgxEN3NFIeM/1q2EwLYK/+8qk1dL8Nt1QwUJPvcGNI5U90yVfzB
WLinvFAPyZw4Y8T8/xCgm3S8DFsKZIGO2lYKnBaZYHJ+KTQ2txNwYg9XhAZbBjMw
mxIdBeO+fg4Lict2epJ5SrHSbEKnAQ09rtuS2DQTLQgGEwfIEhCEaObYVXtzZFNo
TRI0YiQ3KC+qstkR/4Ns8UNa+M+9fKUxY3rZ00/IfWR7+QYRqlxxDYNXFx3i+vxZ
66s+7OVeNt0vc+I7PNF7B9fLXo5vwdlzOVFNDDdhSX+Ww6YRnhFoaVxkoXKie2wh
BQzf24rHoGZoq242S9J4AHA5Og9PKiHucNdTO/89LlyLUCczp8ya2hTSckHLacDc
2SFVZ7N0b5KYVLGdJ9L7KIZFgI/NOOaXWCkGTi9w6AZQ7HE0TBayCwnfNVx8hEOf
PQXyJpLDiIw2ZXajilenuEmuTD83ATW5CwfezLvpbhtdbU0yxCPb9tJUWBYhY4Le
shE5VF0lI+Ilxyj1p6AI0lplqZdR0d6Kw+MRdsFMA5t5gIlu38BVEOM7Mbog9D8w
xKlu/67pFO6EzG71YYISiaQcliyLuNgfFObsLhricr4s9YkYbQfJjLTfONQogrSN
7XHTeQUBo3EqogswG9hE3Xdo/bTrxWzDq1oc6oGAY3FyZtHhsar63zFm1atFirGP
vKlD0yppq+vzJIbHq3Q8IgwBfpTcu8JyXpmIABnMmYBYHak/lY+ITjgKDYCQeNZV
vfjKLsIaAqggT14W0MSeTlueyI7QHa1yPywA3x3waGR7OrcFewbRLE2AgAXYm05a
H1hb3akhlz+5uSY7Qq/as46mrMRF/BJNV2xmBMt82o6pT3ARO1VuYjjYn02RUgL6
XyLYZkODdE8VsenA4bo2G1gof//3pWURaGVD6bA1wNvkBW9CJlXOG4zCX1CStFLY
LPg9z6bh8bxY4N750+fPRzzyg19nWMpVspA3yJlZXwyImSDeHLSrkLS9cWKVcyoZ
tkoGU5aoxXsUMK0jIBGBREBkmwt2Pb4gwcNCpeUKwcPN12StEhIvn0sQbahI7scA
2G9PGJ7G/cVyWDa4Uop8LQIzsvb26G8pr8qB7I4aNlB5x17eHkzp+ahutle1SC8t
oI2EThKArIz+GzhAV4VX6uXGyGrP5fE5TECNuAfhegtDtygsdnW2WsYWUzfC9+9l
Jg63g/6iNm2ZEhs+7yH8SpD8KS5d3aKU9huMqe0MgkeRbfPIADf44pmQ3wE8xpRQ
59PpHtgUUxIcFmpzxLPK1XPiE2zhkdCJ1epso99B1jIsJF51Mk/RnJADFOd0rBN2
bokFe12swg2Fq1Mvu3lpgdYI5Zx4r/XMID2lj0C55tbX5Bg6pO2oGsjazMEwg7g6
Hc09fU0V7RJFDoH5GGce5mFuCCn8ecdYCGbplrVrFLGjE9gsmlHJc9Of5Ita/k65
v9cBF4hnTUX9Rx24UUM/G5nNRa651V20mIAddK+d9cKozTsWhrAwP0ZzWR7p1Lre
nsw0Czo0+vNuzFICup5JJluaBpTtNVl9UNdJuKBg30eYE5neGj9kgjZtRIR9MVXq
atGlDLyhny9grkuiWUG4wQvZJSvufldtaaTHW8Erbkf+0ymxFSsf/dfNGOXUSwas
//tC35xy/OoZkk8nBRTR+NYJGZYRtrUzXoNDfUcpTyd7NO2StUUZflXaA3iY8If4
7pBF4xRScasonA1uGr5+5k+awK3cMmPw9RJqLZLLHPcrZ8GZAZuIEhua5i8mZ5ec
Dzwu7jX8eELQB164pElXBwSQOE4alSABazACxSeL+iNrfyljsIVJu3gRgjkSYnmh
Msgf5uZYR5/X45q87GpX4HpUfUF3f+ACOnpbs9Epr+QUDwa/Fc+2dZ4ioFDgjYjv
MrAnxaMr5iHUbngJ3AbyFN4EptElfEuzey6gj55o8mo0eTx/d0iE6Cwke2Pp4gYY
Faa8gxrgCvYfhHRunCJoTW5yMzMEL7+q1aD9ysBBOF/LxZpOnXS8rcFg5xvAKVUA
4zMtvL2L+9QTKjaVniXGxAy+s30VRw1fXvb8jylCzz+ySp9+uvnGDG3Wjn8ZCrxL
9q/U8Lz73LTIXzbtIOJrjVzLb5V0UCGWdyBhAwUHRTbBhVLink0VkvljxEprZaB9
DDrjnUjdaYOv0T30zOk1Vx80AowQckRqupkrbMBuZG2YJXQEdHf2gidfR4MVFOsQ
AJHdlU1JgdYq/1rVj9hrveRLScTogbV6kenmO7hh0GZh+tspO0WO4y+jg3hqU9am
rH5Ap5heYw8kzKO5AW4dw43tANpOTyBlghBT9aL5wwM8WBL1mprms9I4tGYqNq/+
p6jWMeUGlL/8rsrtJ85g7ex79LJI+QYR79pLvMa5EyqXr04UPNuK7AvaYSLPl8++
W92IrQBJJxbq8Ah9DO+mNO8WqHCI7G6b0T4u46xhlRkkYZcXBP231YDQJf3th96G
VHdPYOGD7L/xVMEfstZbvixo4ll/K1W4F/lEv9utw3ynv0SrJ4QrMDnD4tjMmOpv
zCKZjgE/4vXLfV41dL2lzs1TN+GpyvrBgsMshbjoIcyBCc0C66X6kRDPlU4NP6im
O0db+LCAfpYr5Lt0YFF4H54aKJfmtZVHv0GP7sydBv2Dm5E6P7TQMWejY/MitEFc
RRjjPoQGNJ+o8ixwiL+Ggo7Nn7KcM/WpK/jCP31lAic6juCPkF6I5zuanmCijx1T
QcoAcTibR7u8ieqnlBrMYsI0Yrf5CJSB6n0qVxigM7xnr3k5YZzK+ZnXK+5DBb9r
0+YBIMYvu7INowf+hQJ4uZoMcuI1koLkzJpsEDGmQzh/vrCz+6jnp3WZWuRRAcWj
yvto2Q0QaCaKrTqYBXvwP9WriXbhUEHLoujIWTRHTKFhTm8R80Wsm1RIv6Nr8qYq
xOb91KryClBq/qwSpOfZyS6ekDJ8dmeGE6xbxdku0+bhro7PnI16VDMMdDGeTR+E
CjQlwL/K0g3jA0lr1oKsAA/uS4wwkt7xG2752wPKJzlTUBe49ypOdIRYM2ZRDlJc
kGexSf2uOhkIo/PfuAkAkBt2f0SRQp3KnRo80zSAzPNOQRsqlzXqQE7fH8zFiZN9
21aCLpxFm2GiMQzECCdaYMjDNcYhr4ykeV152DVxOqnDyida9yzt0wuIDeI87AH8
NOXDX9kCOkGo+gwKKKBejq0tYNOiyzpB150/jkfMjpij4R8OixVNrfgFutFW1T1M
wI54anZXLzRh0y6thH6vIkMwQ6v7/ANeb/Tqpx3RLq3SJQ28VHQPxL1SjTAegBy1
Be7910RbeZMZ2+6FnVw8PbYh/OBfUwjqShoT2CcObAER5m/av6kZ/zcNaySaBoyD
4nG76mW1CMzq0tO79Qpz1PUjrypwOBF6QteoVQsNDT3e3OqJ5ljIgYMoNwARFlRl
uAW8eyOylQSVVUwsKLNwtYcdfSz+VgC/NA0PzvpS5vvP5vqPPzcP1yHJrjldmDCy
EGvEbnfvhxuN5l7QkW2Y63trH/+MpXUNVM6TS5M2ZnODlz70J/QPxJSLpspHsEzS
vTkHt8LP+c9VuPeK3zU695vGfsoCdEBAVgR3Vkz4KiiznRi4oxZXseCs1CcQppkA
SriKFSWDPC3UlThdFFgGz2Ok4DKrbQTR/q/pTbYzW3fv1yiBAZnDa1eUh/PURmDE
zeGgNyFcB2YMFwei3W0Ld4zny5BGa0rB2EUr/19tLFqITje3jcB4hzER/Yg7sv3s
8IQBRQipr3mQ8KxMtQeFanravikjJkve3XFH1qzZgC0c76y3MG6+9eq8G4eqwZTz
pZ65/0alEdeXwRC7XEd1b08IsKxfbkmz+KjFU6+ttAFZR5cCBsgxUXszcppdVjY/
LEUJAqce/E2dT8bP6jV407OJGWs1kUZWB3fALzVFmS+7qBeGI3hc0Z230ZmsHOP+
GptNztZzKJ8cwHALxCRV6W1pjAiHRFhyxwSF5ysjp+3UY2frWesyqOka4dB3GXXi
h0tjD4xTcAzSWplJawGzSVqQE9RLCdEZaZ69fmiFQWJ7I9e/xc/0Cvefmyo+R36q
vUusb814d5Ifa5jUmYMm1+JHApvyaSH972kicD71TYfE0jltFwQ3kznRjSVZOXgL
p77LrChmTbTY6XZ4zpQGeqgcI3ln86UazMXXBgy1IoOxBvvhUCUHt9kzzu/P15nR
p5xvfVOCaNs3rHcwY0wL9/aWRDs2SAEfHv/5z049KuqwpkD1BiwHRbfhxXv7WGdM
HKZ1mGKqrVqTOWaj5hXXbfZ/qzaFO0y/zoF0sM3gYhjyWpujcoJ4LX6YebkJSFA/
+UXyiuoAat5eNm9gH4R2fIdDRDvj27Y3u2u64CJnO3+qaFgClBITqHAI4Wkgt+ax
cqppbuckYGkEi1ktQFD+Mjw02lqzI+pLiMnThOQh2WZ23MlnbcuZhjnsE1hY7MUL
IlZ+DsQ1NUIB/IEzk0g7Jv4yR4woeoZDlZPb1NxWSzG5fEUi39Hy7ENiqMRMx2+0
uxHqq/Fitl0gPyUhVZoHvrYKnv15VB5wSoaKy6kamqosVGc+n+amlMxsxsLPOs1W
Xeo00Q1+jW1bGDOUAWrnA2g2mWDRNwZkeejYE7cynATc+ProFwdclWr9zryrNjj8
q4JmWZGTchGrqrA5CYIGuTOfSfKCH4z0jSmNoLCeVOT0p4SeY3rXIY5Hn9WfILmp
rq01fbnJDQ3rG/5mgk0UUXGlfo3x7RDf1BvYpPCXyW+zcm+WIAwKU7SZr8Rg6cRk
t2YidedmzH3beOYPVQaRL5EpT53ekrLTs40HygHKTn9uhZjK+K8hKV7b2KwsRZzL
NHenwzKoBigFse1bDz/q+04b8Rvdfm0PQlUbYR7lS92ruEWNgkEwax0DQQ5cRbtv
Tk5OQNW/MU8fpQXR7eTYDqAj1jAtdl2l1Jltqcrmc5VG8zfnRXb/gQavrHAB6Ib7
dWzLAyQ26YdRzp1P5mxn/Z2nBBqv/OZDwfJMjbjbNnfVGrEjUGLze7sjMxEVbRU4
rtPr08w+wD0pSNNIErAJMGByl9+00lllzNkVd1IEMcH1sw79RE0y+TU3WhCi0XMM
7wVxSYroQu37qJUrcHUWBql3lEldSbfapnvUQZ3mlXfN0cflH0T7oaLUcmI4bBVZ
euCkZMbCHCMBfYicp8835bD1sVFIFoUbWAQUnLAlbYV//fxazgmZHMzgrt2fh4yZ
VoSOOORyUSWHRdhcdhHqIgQc5Hg8ccZBWNuzGPVhxclt/fgOzOe3XdUU324C1dHV
pOQ0mop59jk4WANDVp4a/zJWz69PpEQXDLAzQwRLZs3aCzSFmblrfBmg8PM45JvV
9DfzS4fo5jyN71TMYJAMlJxgX52ZNnPKNjPxHvHk3meENOuJTWclFtnIuUwzJ33w
Us1Cy9PMlRxpLfS5Yj1X75qq+moce3bgbqbiKqqM8ui8gQVNxtebqlaI8OxfzQjY
xsCpFyrwd7wV6HYEdI6DQD7hSsdGPOiRsdhLA1hnlhNYUPT/ctOsYCPhg+rcee4R
bCXhdsHt02Isgm4sRQ4ntlb3G8wc0V0bXz70i7v0Y37QdI/rdfgnR6jcqtBUeGxL
c0FzY238i5RV33VO+JiAoZgEhiI9orXuKw2MKiobMvVcDWBbddVH7WEvX9X34Jfq
Zo5nVR3EZAudvGJE7X6SUZDeOg0HJbKCoMp5gn9mPN6kSDkrTxqRxBPE+ew1NIR/
KKdnIJFo+VULPrtvgggIT5xuGXOUqxqHiYIoquF7eFBOrFpV/lE/L/YIJD1BkRmM
JZAJgv/2rnoJOSQBpVlGJaCN4TL9U14y9sBRNmGWHcNwNwplpzfdYOrbN7qEIqhk
aYlIVNuL8PqMfDTamFPCakS+NRQY7uj/CmfPIB2eOmeVHrH/8llVNIdcwjAGW7PU
2OuiS6EAREXRd0ApxbaxxwnUaa0O1vjmmGAOTHdo+Q0PierCpNTawlC1BqBPmOcb
ALpWp2XlIk/y2PgNyV+L8qbAzvN7GILbGlfqAJgkOPwPbzymGp7/yU0mjt/dsfqu
ZJli6hsU4CvTIDB0AbM8CUJBuf5LczFobAsn2XcRBJWqtMswhaAxBH81EHR3DI8s
KQkTJtLpUBn2H7DkCU4ydXaXYIFMxdBIfzG6QMiITi9cpFMCYs4/U/wSBDW+XJA0
7ahJGoXreue8y12C8rCM7XTxpFmgz3a5fVWu/RkvqZjpbVetHCoRPJyusGEJVRvE
PPEqxk6nJUdGKZt9M6XQUhd+1OYnhlqOGYXsYqRXBsqXLS+SPG3mBOHm5nMVCg7d
VtG7F2TEBuhwoallhI8CbYgGSLsB37IlUBvxynGoVowBLgXnwOVN3nNvTg4KUU24
iH1Hde05kWeVey9H5w0svv0w0Pi/61K0gf5jJ3qHa4FPMdZgOepEkHGC43aGYIbL
EDXaehFwRqyFocdb5uhXg48daNTa9FV5GaCeQUQiwjCI9sKzARV8zvutFUs8dO6Y
MNuS33ui/rJpyidCA/W9Ou/gTOixz/A2tHg85HKDO9eGjCzWAXN6lSRmVv6r8d+m
H97KxhO8GjDiBbu8aXr4ZcnjjpvCRfOmOmNd2bSKOlK4wH4lhPdU2CEQfvgBMNPH
60BUWJL+H+HUh27vwvMEb0oKrR/+BN0TTX21STh8dF0kpbs/WpV+GqBhQ74XC/MH
AlBvzYmPmTVt+YWulxPolFsVaUv2bH7DaXHNWF/Z5jPsX8aGNS0VmGSS0hESjb3O
9t7pA9CAAQW5Kl9/ehlP/4L+OGGdXHR3oBANhZAemub8PCtISiqmQnCtxGj27o6t
SwGC7G4d1FdPtBdWTRt8CFBKI4mREsHTTh7XRxFjRYqDS3gkEem4WlwxC6NALuXX
mEf1iOT+b8TGMgl8bXlcQLfMiSodQJ1gbNgGVQWWXxbEPrfrTxKoGt1WPsg2eB4N
zpRCwzbx8wQoZABnDCluRJ5MaPLUQGkZoaxinkC89CnsXDN7oYUbFAALoCPyKiiK
vhUbYdNvKTqVSrvra+YH3jJFDBBhjR0wi4IQuprBhcUkIWde9UAVtzl9D1a9gp2A
Ph13LTfa+pGApLLBszAcMu7mae0zVk2r8e9rmoomO/D0Yi8S2WYR2hUqC19AcCGU
yAmyMmgcHFclErL4OlEGfsam7SRChKVU32s54Xx5qasEq3pJKUWoKL9W019Qc0XK
B+WOFmFZpgSwtMRKFN7Jb/qyHtCjeok0/VMPR3TgwpZXICDgLLVlSrcjQUGhXPGt
2ePWsmDtSw6oFv9hoYN1hCdvDYCG0Hc+xpT1bbS0TpeIADlt5ShUNzegqWaFEAMq
F8Ick7aVts5EdnqxNaSTIypnS84QrabnD7Kpl80kSN1Nrei0CMP/htqRX6bZmufe
mtDJZiNnbljTUxcYXUPEgl1ZNZ9RpPGPmGztUOcRXjcp2owhdlprrtqA9NJjo7gm
X2gRs2m/58R/1mu1MMkhbNsY+kkD2sSr29bZeFBTZMyqbirDyAWJaUqdW6ZUb0fW
auqLmVHJGO/wuBeAUtn5kRp/uKgVYBqQjbbTlbNu9opNT6UBRY/0l8WdrIXdahLC
XGzxhjuix0d3Ofd0lvMNWONxxsW58VDKmjFoRHKybK3l17YnarWZDU1iLI9GCNPa
FZOUsT+acLAgUj9N47CMl+IYX7G0DeY0by8TT6jYohGSLu9BOHzksQwAnyX6QtEo
/wHtPTLfEbu8ddwSfWA/qrBGB8BE4S0iiAEUUHOifP8iz+SEfe6Og25nKvZuvkFh
Gr6GoKaDFONm4a5EJtRSIOmV91qEWAkMZaJAIsaNtUt6v5EslGBsWOrvIo+AwPs4
6jxeVBL4sTvchElXAcGz2pnqjEcrn8EIUu0d4/9YTdkzcgVi6cGDUPBpAIzZagdF
5P5aZO+T5TgVGQ5ALItan26xVljqN3f6fqm5BV1mDCThsdX0hcM22OiIF4NMrAGB
JkJYpTi7JFN/564GhkFvl3Hhmis8NUvJ2Nq5l/byBIo0R1lqc6M/lZmxLiaf2JSu
jQlzxrj1UCe8UqZFEPXWdSovh1IhTQK23625c9MYu9E738XnWjGrVP+PAILGGQg/
ahdpvXo89862aG45Lmy36CWWr8DYsoYcc8rIQrIKB60c9na+9CAbG97OPTdAeOgf
10jb0YmsGHgBY1G8uKReSjd13toufdWp81BOGc78qTnWQvhceSxY7DGu/in+9Gat
nieu5p1sclU5Mz+R/edI7aNbyS2kbCTW/NZOEqGT+uk2SC751jlv1VoOpe0jDjfb
3923mWmbykqknfv/6pMZHFq/pgaNpZBjYYtnUonL8ITp4SwycOBgU4xYQKXG6AS/
JcEK41YhrpuPdKAulDoGYy5z6xP1PomSmSL0yfgginuLXd8Z+82QUU/DUktLTUi/
OoCsCjdKtZUt7w6RhWYtgWLdaauTRtxIxa4+dwxlSp50y2l+/vd4OqwS49EuPnfh
CbJvY3+08H9iCVGlDVI1pgBqpVAZiTY/fkkB2LYS3CW3Ma3Ye1e1o3zihntjh+n+
F30QL1txczyKaEzQjTAYrz8VQEbZDPFpVQvtyq6LC8xeeoUsJt3qYA8hIHocxmpl
mafzgyRF8NWDlKs3pOqso7fOOOOMWJkUObHMX308XSyZA2Jh/ujk3j5Ilf1U2dn8
TYO2N3pwYBQkpOhsR2wuRtmwENBtPB1rjbDxT8pQ5BdAt21mbgZbnzSg1Ya7uaTm
fRxzQPSqmL637FnwuGR1qLuFEr8D5XwNwcPYdDDqG0Q4gCsF01LILj9fxTJAHLyZ
eFt1gFMtPidMtcvhfBLFp/vT5Iikh33Wktx03bWAiSuEIpxei5uX1/lYSO+/MFIe
LawgRPPWWo+35a9bJj2V5x0saerfmEnGUd2Olu0ROwFLAjB6R5w9rRTtX9AAkmCG
GnAunN/ioq/uRQ0COPBJKVK9GCwtSmAFblQQzNVTxysaapuUIt8G1G2g36e7GqYf
NuJflUhF2rJpV1NmxscGcafvD3nfZqU2m7sqkxefNiIIVEYglRB0coWHXV86mTAw
dd4CsQu+kZnIQxv9Rw+AoaGs8wYwaTWVuN2Kj3qUNZHByk+0fRvj6BMEpYcALVAW
9tva7Q8y4K/e+mY0f6qSQ+OQd1XIBS0Fvglnt9AqdiglnUvlMWxtxgqln2MigRBX
15Zy3Hx3qLg87r1la8SzdrMFy7s7Ys6lJr9NIphmHekpA+qrjMF8XiPMaMJX7YHp
RJ5MEzoZoFRtHqy9gqnUxksq/TxMozWvwxzCypFFvuO9qDs4JX8QgdQ/79+QFiQr
nM+acgi/ZkN8AdQUjZYxi/ToLYhcCjPELSkER67A4e/VyOcYOa4cX0jj2WBP8H2w
A9uPZrJhTl1FN1Wd81s7esANK337nEuSJWE7OeL2y33eOETgN+LOO9ayz/rloDru
/LU7E3uA/Tx9JEplneHzM8eaa8KWRf7pn+V4TOoKycPFXH9faxhIozeSpmeUIc33
1dM89N5SeOkH7Nqh+tyC3OVU9kVH+ZbxjCuNYtsaRtF1K2ydFpd/nGcdsdtpOEQD
Vn5rKHNrwaNBQHLLiYjNRhYgIC309U8ss2Cw9/z1w2I31beleosGoYeA3BR1pi93
J+GsuFYGnRwgKdpbE8OAy6lTraJ+ocBNXhxO5RWsFnXAdNxOf/XPIKu7EwWQ9ctB
6fmZtcquA50621E3/LZX7vVHcThkAZrfYPN0yHcFjoDjIjWBt/hgejmewxf9fdei
NUPLfVWJnnj5MCybZMBI4/XYcxJMEFe3WYHIy7iuGsLxUNiwNItGlil95IysPNXk
Tq3gWkise/TrYYcJKzx30KUoJEzvcMAtBbxWEcTTfy2VlayrGnCpaDjO6+mgNJrj
Gg9+eMm4EWR+xp2JEfz00IKgjA9ULlgmvay/v/fGZ2OLsbnvQcQrNc5otyQAKu5h
xImhh4L7FxFk2vxiPVS0UFxqhS2LjlDgGpaOxhXEO0nIx0cYOMHudDm34NJg3anS
DRn4w1f+eYZBRBIzRLuI8EwcoVLoy0A9PeRoCaniAMd2on/ZIeKSRH45ZJ/QjBAU
JWc99MaoMDdACQjjZs+zv//BQMEWhjlOzLVEdNZVvfevV4Hpy9YczyJ50Ldnccl1
QY33UVw33diS9U5j3mT+3inUDGjp/s62gMYHYtVjwnVCgPLZJGxJyiZnIzIcOCvk
m55FYERsKc9aTchbQMipBey0baqjmOs1Tc7Ykk7i29UiZ2kAmoEip1uNDsbn6zIu
4c+g0hMHHbcZ0MNn1t18IQkSpwcjvcOilEBfiBci3HUsin9JcaeL460EWgXtn0pV
Ek1t3zCnAaP54+pqGEbO8MzYCOaC39vinPL4W6Yq4CzjnirObgJAFrTBlsWWx8x6
PEyEXCQsi3avYp5dlOipXq4HEVLNyffU0yVy9BX+MSqvzR4htvCuNqcm3yMEJEF7
T/IDevreUxFsfDmtMJIyGIclhHjlIVSztyqIyQCYnWaGhVhf5TL0URuI5SHgxLze
AYo+NqCXPi2HNcnyin7TLB2EFBn4aR3QuQOnfBPacgIWFnmD/6/35MPMpomrVitI
3q+YXMNES3KkLQ4sWfCa39rySxZSB5Z+7hP54ZVjHA7g2bcqeTYdIMGfre3DLdoc
gbFdakgrYRCt/otc2ULVxwIvgc+Spuy4hPiYrBzQmBT2lMJrzq5mpuztKimhcGsI
PSyvX2GJELuUPWuArEX4hLqzD/VCwRfKKlGIfnUi7agNACDkf9XDUa/Rf/Z7ScTm
6zes/z2oRqHVcdOi4c38fLst9NcoxOuCpl+1b9i/vZVjWvJBTO6Nya3OzTDk1MnY
5TB51V1xtU3Ac7aejE0FthXdXyy1xeqRplPnd59ZGls2GO6VmCrtEtMHzgME4aMG
AU46FUcE22ywfWpY9eXrEag1fIfCU+WsJshlfGMI8Ri0hx43iZ10oYWcySlpVJjk
r2H0HjjQD5M6QzMhlWk0ZwAWvQLcngpqSC7BzkuYaae2DlUZQDaAdeyLnmJHsh+S
3tLK4DB+0mNV+Ja+IkK4oT68onvFbDKg//BGoJE7I6tdFUMiV/BHIHp5zii+9DQa
HOhVSTP/sOJbA7ZHGgHT0JNvReymUODz68T2RSYVczH7vHVerr5qN8q/4Cx2Om5H
39Z1BK9CSdpJC5Be8NNMDwQe6nX/p+fHHYlL3E+7ycbrx4+r48FAH21vbqbzkoNZ
VVnqHF3IlxlptMlkQ4Q9D/ZEASexiZLBHrDnfYe3yPRNvQiHfBIqHgM2QBWf08gM
c7EoAIwCjMkhMl5aWj5OzDYQxn3TGxVupTl5B46g3JehvdXjeWI9Tq71IudTo5YF
iL66DzjHqiV6g888SMA6urBapn6OiEnCcFRjih8gHlCbSkSvzc2vaA9Gus9Tn2Xy
IJvxgtlEn5Ucs/Hc40dMPI4lbOTINWYmgpj07Ivp2deVZb0RE/oLKwViK6PA0OvN
CxgiuFXnCaslCKhJitTrIxFf20g+u1sTrNZuMox5Ku6e+qlaj6x2+RT9lgixWwWh
87CdtIyN5SBquSPXcqIkiorfNFLRbqXk6NLIkrCF7CXr1FU5H189tINrFJljBibZ
r2EzER6TNueA3xbrjCBlPglk1ccDXEZS8woYnIxNXikzEacvdbLvrN0SAQmBfAVy
enmxs42m6UeYe/9DGXFfZ6g56BfHfstCAhKTSQDqNTa3Tfj9ORaZwnsjkNwhUwN9
D+Qjq7YaVRcRaW9fc23O3BP/BBkFA5Kl6Rg2A+My2HrLxnHE9E4+G+z1l4FZ2/9w
rLApbuFmZTfu4YL3hwqCWh7/MjqIhpQXwodg9SCpZ/1Ur9TnrxVo0ywWeP+V0pId
vP5D9Qjge9vsW38p2Te6UVZBrPSG001LURzeLQAxuJNFhC2ZalPJy364K0eq141f
HA8gSt6DL9wnsQaMfGIak7R6TZt7oHE3GjYOtQiLeU/obfsAQqrh0Kf9erVQCl/9
8eHTSGQRErL31AhyB+vVKTh/zjxiovr0aWqyuJoU6CUscDOKvH04+nbaH/bfebCO
bEFxBkhmkQ5LPliD0OcciS4/76CErNXr17POQAyDPCCyukJMoqTeRLcBHuGob2R1
yPilCwyVsQPewkxkwxGduNn1/LTjWHSK5hvvOL7ygXrIWsp/f56Krws+oiEXyzhi
AORNHMeUyBZyUWkvRDw/jyjykZF+8M7zwubCrzQggp/Uwwz3mzb7VE1dJlti4eyQ
NwGRSOVSRFJfk625XkozDBD49xbT83eR2gdAUv00mmMnEl6faAn6EPrJW7w1+Zz/
YQGxb20SpQF4oHZgnMBVCjujnylHpqM3MUQ21KgkKlZMEJRE8cDiQsph8at2Jivp
/6dWNm1fyJvODmhWZobS2MJ3qLYMQW1iC6Jhsw561BSDzwqBk/jyrRnnMhFguUFp
fBS8M/1/ZjkdX0VgQL8CC7hdJGigQOzc4O9WVg8/DXR6nsINlXHn5u4YebzCjY1V
9ToS7RK22w+dpzBvIke9Th8kgD3RFrP3XBE6WT2okO51n2kr6pXrfiin5O9aLypU
aReRzgNvvnsOWHMoq3dZ7D0ET79CwGQdYgFUpiLIcbTif/sY8UkRfsm+/CWwrsVm
uwhfAe2DnQHtS+MdYoRWMC0HzcXx2RdxbNlzPu6Kukpk6bAIiH91r4CAEXkIxm+j
GOr4mJSsa7YWA+KiqtOWp8W/pkQlutz3tv0zsrCiyUyrkRdByjBYlct68JBdGKOr
sertN1Ceq/+aCmOlbdaxyomDQmuY37z70Dfes0G4hn9nuoH7W9/CZs4cc56dTW2p
AHocD5QSbLnzcfv8892Xba2vD7Aq6bov64gMsT88fI67JIGwajaoff2L6404TCvk
a5nMr8PXq8qQfb2QFXX/r7YBNjUx9D1QSMw3r8e8YDDiXpwboxFTRxGAofNVk8K4
h8e2Xsa/fCeuo0ROMxZ5/6XTWwsoT/Y87qH8anihkBXlaGmYCALCyftXhMhJa8B9
2JT51C3vra8EpcFzVpNWY7cbKyAqDWXeCXj4UY2dwg0BsxEl1OMzXAI818+Jw5Ac
3KiNCbEFEVnDAwwNN7+gOLr6bIZFMTZMVrQUGmsEqBezO78md7G8dK2HtL8VWk03
suUWOJlP/WPUWPwX/F3vTRn2eDa7b0SV369dFpD68UO10YA7fcL8/Mvd8IW+Mbwg
CqoMpiym7bOzmIiJ9wklC2CKdU+6dC5BZA0HVl/tDzi8MlZutXEFzjwmFc3luW6E
ivWQqyAe0dBiT1x3xHgFhLBTpT8S2OsCVs4iWau0q1T0iN0X2ifMeMATFqJak3FC
bO6rTt2jnqqeJqdOTz+fyceVp0pAXowoRhwHOiTEq7mnjZO9aDCQm53lgnoh+B2K
ITiXigGibhqkqBD5Df5ZdbfHyKEznilq3iZouc8FKTzxWA1JVdfjTe3Qkn71O+pG
GoO7OPiCgi+b8l3mBb08/URZdqllk2IORkxdayXW80tUhz//tIjSxdLZ/tAvW332
0w47Pc1+sItaqVdF90UIS7vCmSMGAq3+fChI4X8X1/995PkXZpAd0uddt+XHEYTS
QVLEHFCGbdhRzohcfzGvKTlaakvt8lyoinFEn2y2Dsz8XWIGx4bGxz96YU3GJ8A8
t5JRB4Lv0MZPv3IxlYliGNrG9PCJsiBPsmtE4jYgcs5qGZ8PIpH7kYuFfLk4OBb/
oZI2WDFTvCUKgBpoPbYONvoJYb0U6XUhA38l3yDEpv4jCXUDPD/Rd0BRe6Xm/WZ8
gICP7PuInnfu31iDvHKwBQ33QP3AIDc2ZTF/ve9i2o2Sq+eT2tdB7XMl0s+21RIO
i6b7Hsan3hS28TRa9c/98tBmHX3aJwGChFdpWX5/NWd/+5RKYLqHf7rJI/F+Bu92
+gqrJhN76ZrctWMJDMABCGiM5ozqhpJRkFqVHXjzhZkyxP5+efKb7MXwpBEnAdjv
o6zLQ2QD8PtaOdS4iddAnCWgyzfjPa2vNeEhkP5BooSo1UAAkZhe1i3x2/NnQHas
YS89BB/ciiyZtLwHGYvhWkDseCx/MLbM6YaDlv+fC0zcKRQIW8moEtq2C2pcmXeL
vdaeEdhF1HGd1TYkGizlKoyfW9kaaFL2uFOrOByODN3+ncDpV7mpXDVzdYvDVNFG
WmBJ+raZitce/De1vJfiWk1TqlepTxealLvV+DxKB8Q0kYPg08f9rSqsauUhQEPd
Ir+QW0kOe4OekDgChjJG0AwZ+e49wjDdAxFDU06PdEqQzAuYt+T6592D3oM20qrX
epA4IynCKQd7IvwxC+Rz3zV7rk6O2XWqmU7QG8DKZS9ysa3SIpZU7fBmMqwV3gOJ
zgTr2CHaPg2RukTfskXxfzR/PXzCStAJvRkCquA74G8HLImmNKku7eDdj7k03SiI
u2jJz1JPL5JFLVwnDH+Y9sVSwpnlVzmIijJlGtw2ofWwipQW212LHSrP0txhGEBn
HdpZIto2lK0/LjXWX8Ymkl4E5KLrvy52gC3Y1FF5Fc/5RKAEGnyl+1TR4rrqMU1o
K1WGwiRxB2LL3VrFDegpdVdSVfOTXbPPJvSkHPV7cMGTwB5KQTKwj5E83Q+Yywrv
MxUm9KDUiXqgWLqAE2V6hxjM4qpHO0JXqu9JFwVExRf83afV6LkgCNMpZ8a3BQIR
Iw2tVhF0U0/fkHxBvox8JeekykdYyGuXnnFzwvZKrf2ZQQarCoxj9lBxAk+Iv4Sm
qSw5Xuwr/ZDLb/jSGNgZst/gNEjXhY3yeTyLtjd3YEmFUVFQbbhCVwW6tAV1X0ZO
1GW/5Fooz26MEexiMeR0F/M72oqJYjQrtXh+fPlEWDerA67lAb/HtpHuAIcOodnt
lI+XFtjbFUw8pPgv2KSrShGpvqoDv6/o7qJWPkLKHig6xmhLeTr35gF3dD8Hu/0X
xxmFqvsWmRESWAr5+nMd4nn5m87+/UoavnP7vwQ9QCsUXK7PHSErTKbetOwmxi8o
zCimQVb7Pwvtpit73F3qo1fsi/KMnLPWHS4nepiv69/x6RI0w7YfDZu2A2OqxzsM
wvuMtTcQclmqlbb3v7+UqPpYdwZ7OOAzRuKmlviUpC925OLznCAgifwc5cQDs1wn
WHsIZ1udh6sNVKqvbOzFwlQdA29Vhjmu+KqTa12h6ClyNuyrGm+H1YQsGsbR6scn
LMUfchFWnLo6+4Ex3ZUaPrLj0x8htbRAAzkqk8kBaCpns3x4u2Bo3THfZ1HfXgzI
99N55mF/UISZ0Jua2/wGawWxFqUSCGE+ujEV1NJ0Fg+viq4KQn6hATl/jYiM2vqe
RP4EepcWi9pLVzZAElJ2N+KiWeJRrpC9qeynTj/d/w0LXhsqTvAf/JzFkKDscgHo
BGL+2gzpAp01/5UACBnaKFSaij/ZNo3zg4ntWrYFvlso87UXIICBli/1nS77fcBk
jCvoA/t44a0RYrypqpWBe2rhuuNt4pPB2Mvjn/qMl2YlBE3v/tI+yJzWjIAI6t+5
ZXFxO30ww4jcmccB4c/dg+Hus5l9yXAqKr1BWMpNTpEX41a9t201T3pGfOL75+9Z
g4D522lDfwbX7zjXpXKuG5nMi8qLwWk4N31gFqLvNQCFSKdoUnDs8AVwFx0N4hj0
mKYTY1coEzUh09zXw0wyYbLNpm+wIcUY0V6DHghIis2Fd5g3N68vFoSXlymVnn+p
5/1UqO1DxCWozIOHHuxnYVTFV3Tt/EHh7GWh8gctIJao1VqZyeHgYQG2JxASYxo2
XE/W1OEcU9T4Aft+XCr8/9xsKuxZJQnHOh+iRoFd4sZhQJW6422bucvCNrkkcYjF
O7cKZfwhNAUCkXXBIrjsPKcI+LIQI9I6T2bQIPswH55u7Rw0k5NNxHYnY00kuWHB
/gNMXS5qVpdaFiOPG4VXPaToiNX7Ok5G05ybvFCAqKMdoGAtiFGuQA1TxCme9nd4
D1oWql1j/WRvE302RHIXGrSXYrtYgoFxinFOthL1dh1Z9iTnmo9W7T0fxj4pxHpp
CDs094xJ8+iBSu6PXHRA7qOZI/ZUDQjfEreiDFcHpAfPjk2PIbafvr173FolllMv
i+d0s1tdKHIIe/Gw2HCbTi9kinrWU8m4fvgIyZxFeAtfW29ZQ/jEYFkxLjdzI/ni
7j6BSOk9SoeAhKgiHi4SRm3QZXWxX6aeWAklQZsRCZeFoE1O9KwEtaBM1SEly4AO
q6YDm7F340M8wokg86IJ6Gq4qp99qveTzv8LXm7KBtmD24FrYxeju6DTmzak2NP2
89+7ncUVVUTO3CZdNZnKLdC02PbVumi1oZdjfnMSU8ZQMRvERGR9E5AXLnU6m/5l
mPulcPJ4IhF64S3/qbX+HfaPUbIURmp39y0pyfurqLrlblD9q403bmJyC8Pq1Cdp
RGrK67nBc+a/FCKlIT6V+w9XwlbYSHvqSLJoSPYQ5njPyWm2mTY3ffeNvp5TE+8n
z0Iug5OOk3u1n7XQ3F6dq8YKXH2TXeQGob8XmqzOlUdtFmdRoytyQzNx/+Hq0yxp
ElkC3eeQPQlD+ym+1nZIzpaCz63eGSfhK5B5kdZwA+rQ9YBQmYSWCAHXuRrcRgR3
fcivBAAEGGe3Fa6IBoJ4Sug4g88Wy3F2n1CYByCtleS3hqwIu/vYHhs+7W4cVzmp
j15up7OAJGqdQ2o/f1TNrle/yWbajkYThkb/0szuXGCIBCFyXLDwHszgqWWGgHVa
0SxZXE5ZdSjDmrucC/A+VzW1/39cBnzb+45xzrXBubWk2UK2ziG00bquIx3s7WU8
AlhFvna6Zg3I1NY5OcoE/B3FL2xvUUHJy5yWAN+opgr8PLJsAY6uuTUFrxEtjtwz
ymQ1hSG1GmAGDLKrW57dfh37ZQZky4HVM/7HAwRiOWDdSTnljeErxV8rjiTNZwRd
otMn2jWlgOh1IKgvH1Sgx+XmX6LF6vc+kZeU3uOO7WDRXf+sx09a4eE8dCdYmR9s
QeoZusIc/ZuIHlslKTxG16nWdrv7jf8dbcElfXobn8ak3rTG0nWZZsE0G1hzh/4H
jRUlXfojA4TXBmo5H6PM1+5t7G0xXcAAEbXcE/6f3BV9zhlisOLmt1XbtSNkFJkt
1kkzBstA38Xi6iav5c+aLlKg666HWS/AS4zNjieijB8lKOsmJ9/MwU94t5x3gahd
q4sFUJ6KwxQzDh7gXOCRfAvBhNhSsD67dh/Q4ivhaNPjHqz88qOqIjKSByh+ofVZ
twnKHD1miHPe4UkFuaaurCZKJhd2SxbdyMd+pXyb3EOMsMCdn6VYyo3XGzgmxiQB
0FF430C1ZlnL6OAYijN9RhhEoi1NbJOP7FoG5wH/VJvFb9ezDZadtjNv0YfYt7nU
SjvMMIDzi4LGHFAuFPaunEwz1lqIPbfnl0IhaXOLox3Lu+EmcuAASCb/Q1AtPQAq
8ifizYENeivFmbdOb1AgqXmHAJEmH26uR+avMZkJFFgUQxD8gOZscq4eXXpqp0Bk
vmasBYyHi9nGtjuKKtZUbEdgLuGPuNQBLeSwfz/41BfZvYueCza/9s1xp1dwLFku
zd58wREtjlQe9oKGls7k92m3RZ5DDnj54Sg/W7BUmyGBPgE91h5ine/JN/3o5r9a
7QQsLnIqCQ7jyOdLc/BW8f+d8F59XQcZrJe+1raUtJuhmrIduL3XAgWaQRSBvvo+
U7ldkEFN86Gz+D6CEITQ85mDwcvs9RJ/2N2AE79mZ1/yb54OZHA1mApgLNXRuuQ9
uDfo8yy8aRzpVU0Qd92naUWa4uXo+hekjtwGN01Gy7SiQhJ51s1ZnjRQ3+M8RDK2
JPB7cEW9nyoCSKmtXULaFSnlYQ1b1m1K2jfww/6S4YEwajaPcVbnlLaPzjsCpAG6
ahIywX6E+r203rwWGjfPm/iBdaeJCd7lMgdTqUbIahQhf+yYdYBbv+eYy3PTYhDw
z3ClNtLG9gFB/Wv8TUIsI2Tm5D4fEGn7Vf8ThOfZAOzxurzWwqFQbRL+I7XIHrpp
Wbx85xt/29sEiQR0D3J25f/675EPmEtQZdHdou8oLylP4MOu9gZEGSCPWpcdxIWr
JJJ2UTOSnmbA+i+00uIq+/imzeygZPUS3xQ+4He53A6W5/mHgAsQztSBwaComdqg
/LPAK+fuilqQpvFE5mTOW2SS3kGT3H2md3nVSW6b08bi8BDciqvJ9SzKCu/5kyTe
rprtP+TvDLVLhTsOOlpKNoFN+VK7HRPgy6A1bmp/Ba8FnQCu/hYdwWP5At2p78PJ
wnhfdYDhQ1Sk1OWgjVXGsz86q3R+IdyROjrjmMHkbXO2It4WGawaeIj0LM8zMVUU
dFQdoHAxvgTnR2siKDXuWexNruqFOJaZ8PjbKqrruQJTgcSrthVVA7YdBe0yEXue
dw8joiBRnjHyzHQts260SYzuDW62jNU+pY+xYpWhEP98vLv6lSIvxEt0fHVrf+4w
1TIzBcPfBR17YUbF1VPq8vOlI2lBUmBGgMfxAz99m5i5SZJdmF1nmqBReQLlgb44
+BEP00XQIy49rPBtn858IBZHDSr7ZOkGNV/mHx2nlyajyLa/cjEwocpthy+2EN/1
+tWw+8SYwkwPXT3XjnhIe9np1TKy2YIeyKl7ToKMxLdkjVu/oAq100DNxV9aNjCp
5kQIzU7b2TIohzqJsqQnJV65fIh9UvsxLkRRQScZIAHAfyDgl+oYlwejOkRLBIos
6HJpv73dLgAV7O5frt5hjuzbpS4Z0QaBF+cVfT0yn76+XCQwwA3UsR0P+X7/i9Ap
xWW3q2qhIdJsql9doBR7N8zkBnjOv4sG2R/dusUMDoKB/Z25QaT4hhkWcQ+jOv5+
FjpPfAy6Wmj/v2qjcJy+xtTHl08bFL3e8P9ir/19EvVIBF4/k1sNflnsegPbwg7G
2TzuU2bGaKyPotOae6i46DfkCS6GHNanJeWxXa/pm6obHdyhTUVoO+sHHT9SN6Kd
8PMpGOm5j8/s8a/5AgMHQ8DZAievD+FQQmHB3WCTqUr9SomGgc3dIncD6v42wwyW
7R8L9MHt/GUC63lz5CphC4Vg/9qdIeo9ihKP4FsQfOCapCBdTqkY9k85R0/IvpGV
u7un8Tif82AfjQg3w8FsaVNj9PD1JtWBM+0xwwqe2YqsGtziQtQs13PLIMUaprKD
FHJ7QNfXT78c4tqOZBgaPNAHSvLKGxI6+Hp4JU5gz9ENHRi9dLG2+hq0THGBZpM7
c8HAMLTw3NQyNm3Aqc5yEJcswvpyO00ke6b25Ti5jE+gOCq0z7aOBOZJA89q3NP1
OmE1+5gnLwcNZLXa1iETubb6ktvf9VYeQ/UxNrWg6uOCDBg4ApHIIjIZMBY90/aO
athmRZG1+XRLVpZJoXsP+pJnP+Q73WIR49TSm0B3RDQ3s8npewzDe9B6R43/6FW6
246js9rhWUcDPFjK0TQnLZ6zyH4MCrzVHCevkJDy6Lah8Y+AoqsrhgG65BCGfkFr
TT3C1yzr03/Lxqe7/7Hswq8jbbplz3/DKwcmRKaGZW06MFnMS+Zq68jSNx/kNFbh
lvemdyr3koX1Y+OLZB3su3j6WU/yoFgdwr6eQ00oqYqrLixNLViYig2VZMXJohNO
yEIeHR6xvmp41uX+zEAvcideJ3+qz6nO+4BW9GodFNi4/zWTsEoW21FENLJqdNAC
2n12jcrlRVE/Xi07/lDJG/+dFgnYbDfOKCQCSu2GB7Wmcli7NbTDfvUet4t7zOmD
71juR2L0/Joh1CYl8evut4LbNAncH8yu1w7LX/jEqKKwgIXHF/fM4myUzL3jf2rH
tCdJTRq54PVu1pxlO38v8JiEfsZkCeQLzFQoEP9W4PzcrkkhzHBY0XPyfZ+1WE/L
qSvN5NXJgJQ9M3nFJ0GI3Aw+sWB9ZVIBzLZRzEkqGPfXQ/ZUDlJELQelWZLOM2e0
YYS41DGy7A1SM+ZcEzFDx9uno0mtTdmsmCnM832va4S3o4TSJY31RlRqXiV9lSbR
FfOOt2q4MJaMMIknFxJfHAK9gogHVrmfatdDrJpq9p2UNnAWUWoHHPv+5jTUODIm
+9DdswrUc8bk+shw0FHX/tmuRazsBB/NGshJTdTT1fBvt2ziajYGzbEGNW2YwKAC
wostj1IkzK1PgfyBIm6foPecrV4QU1oaqn3uaGjDZfbdfKS6KOMku2ZoTRU/S5qI
Q/FLgeH6yZT7iAdKEIlE+exyGgdB6MUr0xCNU8TZ/Yge5SK8s5F5BuQwm/sBoSx0
UcC8i6xvboSRPe1REs73y+4agjvQp2eX9f93vq07xxOpumn28SWAdVelka07qaa4
3jt7RUQnLLXbmtgyswgrz0wHEoC9dJnXtmHI89FZ5ehOnxaFpkqO0Rp0GOtBgq6h
CPD+TLFuHKNX43hsblcqYatZMhV2E1Qan9D2HbzcouGZiGa2jNU0lfBbcYeKNsmC
Lnjg1LhHlZx1hEAayg1HCnFzxZ6U92oLgMn+H+Ny7uJ0yc6yryzY+kgn5Ut8rJy9
Yx3z38fkQtIOJMpTqyItBjPOf9RqhjcBU/tSngIk4ShA2PfeTrZJZRiz3BEBFc3t
dxkigxM+cOURlst+WOLbmBBSQIQgRcoaN54A+ylsQfVPh40ohiTxDmOykFLXhKj2
1NUtOOhorJek4BeQc5PQoid32CI6sR7UNCjAcvzuCSMy6bkfXPzTb/0PYjvBOlW3
EQt3P31rigWdtoibZAAzo6vFyVHsh5/ydCdt4OnOklmj/aKZXkmnVmuH8gg5I95p
wqM17p+aAjMZQo7nb+RqBWi65z2obtJjL1V5FNdsMCawBgXvHmiOzWWUPdhwbXJq
D/tHSCSfoWwwxCbQTmnXEcri3KAHtGXB93L+cALeMS5V9xn+YThHkjQs/36/WmpR
VWk/ppi/pezyIGTR3Rg3masBSYshL1/QauyqgWzHmatTOyehfCM7h8mzltf4cT7x
LYWJ7b81zyWtX5v4eRL3BVjYNyeYpgfcNNGJ/xP+Gc975mzP14bHisVCdphHh4Sw
cUsLKpJK3eKguehKoOWCy1SsSECi45/m+grFkLHcH8zNvQPduKBRmz3QYPXq1biG
XDBciAaUYnJnioyCVbRqAOudDKdYqQ3nkCHnxnW8ipGqRndAEJWZSv8sAIoiYWjG
6b9+r6Zi2d2lHe9/KoeeGGQ9aSkCn6MWM2En8r9C/yWh7MTokdEapm28JAMxM+gY
KxW2MC8iWUUnucHi/yqIaRY6ggaSkdox/2nAb1BN14aKcQ7+TUgTAB0JQatOngj1
HuxnOwwPx4qRLSUOGP/DZMB5yHzmqskwjrUe6fkkg5tm27QgYJuMNxUCXWeJt0Fv
d3xQrHCEGZOBQO+ell9DSsJtxPXJqbJ5uVS7oiUOMFPNnN2wYs1NKVHSiYmw+Pwu
VF/MOxxkeONu7dFyT/HnOrrgBHQ+UW37PBFAjIpYWAS0ejxTRhps+eRFOdCsooiA
Yptpuz3xLSHGefnXpj1S3JHqCxMbDoLCbNyMCBQQ5CSXeBfbts/rBIi78Pw0tDpn
6PZshGe4JaAzORGAFFw30F01jHJrOX0/po6Gepb6U+RVNUl6G9QAQ8Qwe2FKPJK5
5oC3pTgQkiUK6rmbKl6Qi4RSf7nIOw4Eyli3iafg2B9SrlZysXF2ybC6GA+wWlU3
pmEYDDGyVOipXu7zWWmugbiQ7W+yd5HAhbBv0aPUXn7bO0jd40wxHjkf5/hl4cHp
MgZa+v1oCBbvdAz5nXbnSb6s4ZvRhB4axhGR9aVjuN9V2mG1yb7V0lZTxNwtZ05v
NLv5vsYOM6pwTW/N8XhLq/SGgW5JvOicaBooE3ghxq/tCHyzvCI79617C4810SGB
CrJfVbRvL1uAVdvbeEKCuyszqsmn3ibEdhBWjSEK1oReWv973bYi9WnJfiobxJOd
s/hjbzLE/7EWWAD1UpYVa2rGMwweOxnq0c7tvMBVE2n/J5sFDsBTPOLaTCa+gVhd
KTEVGRXeuJQTocTzyHiQ6dAt9QyUTIiXjpwg9KpKlj9oKG3YjfmyoUM1ueGizVfu
vsUqT14sDkB9fD6OVwbCviI2M1NGR1O6vaKRTXWtCq9IoR5ibJsOkZ5zT+ivy8W9
7mRVolac5Lr8Zmviglr8T7XMDebb1B+nsGn3aiWsTrbRfu5kLyyvQZ0TUX14LR9j
6THsShrALkXiGewARgZZHT7Llp0d0NYlkynX/p/1kdURnoY6v6tjAK5QzIbjcLkB
Rl31r271jjgNlTwNDr5m9Kx6xnfUba3lPeslOaAhL3lAxIyNmiFR0it+tz1HgdsA
pcZJb4zphDtne7cli0hYvF1MQXa6F2KedIpGAPpuBeZc53+/54fV8qfFOSHn4CIx
iimbv0cXopiXzDF3whFXT+dOe4kx73Jj8LnptoJ1jJVqd32n13ADY3j6KL8rRzg6
yr2+oRSkKDkb7n1jRNfXOvA7SRDoR8PmWdA1UIzEXgAGw+aOfNppMKfrSaAXDt85
OzO5KyBbqgyTXdeZFleajQqTYdJV3bx3xmUckt6ZdaB2XbLSDqqcNihjJHCSKCsf
ETbAwZGKjuyKIqFnr6bpJL85OfdAPy5pgCHBavuO8wRSQijzi3u2gD8U9OGF6uKL
WHmPMhx5VRRcY2XwQ8kqTMLk5s9Ta8DMoeM41X2CDK5a+xRbckfdK9aKXcH5BHvn
U+jTfmDIFAV6Esr5SHhDXRvJYkm0DH4xs9ET67bZmgdoaWJG5dY+nIDdUO4IqNC/
RFK4cF2t+96AS/VPbVya7EDI11HUqOVYG21Ay2STcFyA/FTdzppKBxJo28vWfPXX
nML3mHDAHIViYzCGRNoouhR/oDF0P3z1ho0dB81AqqIhlPh/FFMfqLJGYcXX+Mng
OH0OgeukRzqou5Y0Lk3pg5uCsLc+yhzoxTtaiU6VsfxRt4/j/CeKCZVn1W3qNKGx
8yLJOA+DZ+AUHOwS2T60xR0wveblOwFWW3pMLbltgCnW7TIdLzNsrgoPkCdskHFm
HutKIHtrTwib7k4ItrPCJI9B8qi7imkjMD3ozTIjH3whluAOsuv6fsBAvWiDIHIe
HrTlyGDXKFsHSeK0OEg2Ras5u/JNQt5EJB/973xIf8MnsPtgHy64YpCC60IGYkQD
javvgtoZQqHqnG16cgMO0lAP0rad8Sos1SfGnFmKclKOwR9AtncZSBMY28iG5BIa
ZB/uBmQIcZ51qFyqUWF5u2MyzkinosOEpARDdma5AMrXNZOrlqpOkHCjVnXymAhO
/8Y2tiXkjqWO5BJZfAS3VBzL9clmm0DjbcRAMJNAArtgn1/Q+jK09Sgkz+iXrQwI
zNcOwe9Lp/Rfru7ZCE6tEc+3Lnh5XpS7234LT5lJ0neUqybvvSV55IPIYdeG8Ca+
BG11V/Tndd81IzXd8WXChnAZYmB9E+2G+bwuinFJ3YqYzgKM9xFWP4YTN1YtXgZi
rAfeazXbVewEAbe6k+wu00n36iL4VKitHTkv+chliLIlTr0sMFf+e5sSRggidmLv
LaPCEG/KXndBScYl2gjl3M58dLFfDqRpfAq0/BeUa5NBxlR2Agbf9Cq93ebGCPE+
SkpsW7MJQyinQeEeV+53XHWKXf++2P7x8x6JidCygF8wXsBH/hv2I0wHBHzizGqC
/0SewkZV/WnbVi/aw+XsRpfMKAKcbFmIrMXuAD2gVpiWZSFhOVvM3C4Hlyi1nGXL
1O+bW98/ZsEZZFAdOTC/g3Tb49pF0gyeRK9T4zkxaVyBo1+5++XSOYzeOcCkP3tF
Mm7cyrXIjHqSF5VtCpTsbkxw9NWzBsINu7Kc0FtFiFLgKtUO6YsCyXjtYpr4V+KM
dmO41RbylrqbdwBQjRDYgVgX0gGesEh+s3lqUvS5yq9Lh+RzwZZgcBUv1flRb03X
6sb4dFWcxzqRg8C9Fty+LJhlUEtZO2qwnglf1z0I3+BEGjUODSI7VJg4OFe0ySy+
YbmQfSCqP7VdakFmutQNThhKHWKnJYL08BgbxVcCpCorEa8gxLO4MV1OtMkISB9d
oNy10USQcqCfME/CBnGgRPM3wDz4xJ7RVC1MDYDIcpLZwzOOe7FG4MORRkYMpBXN
gxHLiz4xrZ+EzdyWigqJsDfaVEAD+ayjch0JPmI1Kkim693rJpwZc919hFW5X8ZJ
WNt0TpMOXP7E72Icv1B4d6Xp5tipXNGX7TmJeFFBA9bDVTIhCgV7jdShHSbU8KN2
JM89Nj1dLdb9uTZfihPlUv3SewveMKjRnxA7h6FyBmDi5KFzDx3Js/EYnQw+9jXX
wTXWcALd/KItaUyU3okpTjDNpJXeE8IISGbqu/kMAU4DcDXRn1ZOzBwDCbyNCOwv
6rVgs3aKzJdu0HMrToY1MQdqpZQ4gLaDRsa8MONQybbkClniOwODR7UdMu1PP2Fs
+jXyMz8JwdU96QrvT+AHOb+MKa7qIvDbZFl+1WlplEjzXCYBAJEMLM8nDQTotsnm
G1b5STdqn0vBvz9mfvB1elaE1OSs9MHfOJ0ZlI5pK+1aa6L/X+unUva2zlB6omYm
kDJp94hSQBFjw5pq4nrPsH3ZeAMl1IDSeiHKKOFOYmQtQfzTfU9yZexOUysgG8Jc
ayg4ml5JzGXI8DShyJvJ434eLfVFddwWqH5y8iD4ZTeZ1EBaoroQZXsoD4u3+orr
nnSn6JUhi68zIh5nG6WJJrNt6CImoY7OK2rfoGFvndFO22YyC4Q4iQi8aL48PMeP
f22smoJzp9CBg5Ke6RNYvuXQJAP9Nj/QYUwHkXYH9CaqIRbmoC/FJ3Of8sfhDxj5
h/3SLs8SjuXVQrx21kEhNFHYsISo5aaxqbgDMLpuO+L/JdfoDS52tZdsK7xIr3yP
nDV/zzdw4Csmm5GvVf/KUP/ZqIH402+GZV3daNc4AqBbHn78QQAojZK3ZK63aL8d
+D/90balVQOBtVBGisjZVpJb8EbF9iqqNuug27GdXAcKIiuFNrtw+yG3v/V+VMZf
IkezCp6bViPA6EZU8aPDzrB0sV8CvGBibdFzaosuQh+hHpt3xIBpbT6PeTW7cIVt
NerE6rTGLBB10ovV6H8jqkLpXXXdAvRq10iVHD4Lh3syHqt2Y9mzIZKAfO0g3FZI
sv4yUQYpxa0zgrBwq9y01/eofgRYNcywFc3/lnMqXjIAPCUUAuXTSgBAwhF49g4O
HIE6LguWlPwD/PY26wLLvtuG/xHemOjmd/saXkML6B8SxGCmJ2IOLjtqPrBUmk4O
KQ1Rbi1ZM46qCEZQB4PBZjTM3dLi5X6sPGwfSy8QK4qavVHbj7yNIoVdGuWMwXco
ifwxTKt7NrWPw0Qzma/M5Hd1OR9sbZW/WXkcbjq+1pQkqlhDRwKEDqdqIpajw4S1
gvOqzW/USrSukGCAUtZiFBZc2vR+F3H5dJRXR7x6r/lEj8HH698Nt64JJldL0qrx
5/EgmHpPpuu8p/BzScMGc0/NX8YG4dTaSXUbnqht0jmfS9yc3pLmhiJRG9a0+GDc
oFI9d1TqEyBiY15RW5haBFHozPHHpjZE3ko/Yv7GGmKuz8ZTJISFJwP1wU3bgBzh
7g13iks+VtYOzioCA4cXBUsN83h4mVgoAMaP216Lz00m567yRWuSG/rFoxbq5/og
no0R7jHbLHaGnda98BDTWGAv64F0+s47wnKMcV8JCyUMSudDXlZMojoI7i6gTiwN
nW2YWBqx1ZrgF00UML1ljT4orsEcD+64pfMc4ri6bM/UYohssHygKvqLHhyI4w1p
eQHumSE6++Y5d/hE/A7hdPVjuQ8+EQDzDYjuKCr29gzy7k5b97p9AlsWCnkHMWy9
vjtzJjRB2KaqLvGi2BC3flCM1yO/p98PztjRzZyJVI/DJNqTe/7AFFKLgjp58+Uj
LBbnZPZYf7jh8zhE8KGrdkjJzfq4DVYoCkQIlLW5zyKaeiHpMLdIH13HTXbsZj5F
gAcldbOpavl5jvUWy5HV13oTWdzr0HGGHIbvR4r+nCg7XjoGhRDMZ2RTu7P7G1O0
C4EoFPm9yIvYDbP1UNI3vK5LmskdiDz5py//gwggUn+8fCDOFXSINADJNDNBik8l
3X5oIH0Hltkm46CBeaDzMKAq6tLaDGK1PWsJqRJ/dZ5MI4wR2Sf8KLpRcJy5fY/U
sNzVVUgLvJ9i/r+zbatGvgaqpjcRfyEFrCxjDv1cjEyGhQnak9z4gz7JOj8AOwUn
PV9fZgtWZV8/hwhAFA2DZTlhkZKrWHOuc9r91XsUsJPnao50HdlzcKHPGgGGapZ7
EUjX/wQbu9+l2GO0sDmi/UK54gPxE0eu3jb5O7r5Xfy3GDVy00dykMzCr1dGJR4/
c6V/lOTR/2xz0k1+/z+ZeTS+oRxlbZw6vjcePGCmmTucp7W/tJlxi2XFSovoA1MR
CCogbJEQYtwnkGN6OqdQ4P7ym3CNZjtzs/NvUeeOy3MX7n949Idnx5p+AZARReBJ
WP2mreleV/LYJurd0JtbrnDBKfLSb9jrhUSUrekxSUNAh/V3rhzw1iR0Kn45vQ6H
MjCYL4h11CPzdB41tOdOTIA2i3L3ZUHDy3pkVP67mrvyizGQFFgCDPJDpHRViYlz
VDJeVhuW3OMIyaKfmyisHZZTClURA81y8oH9YzWDSp5L7WEY8Hp+Ys5zx9bZL1mE
2VtJN94KV5eITk8HYzHbpVIM7c61mviS6OqTCsADVYw4X9TRdsINHvAgLlic074j
nkOEV6Bmi/eUVaSgWTwLSsdSzIPlEvrmEQIdMJGjGtLQUFak8F6kpK1pMdDh/1W+
eJhXDWSeDOZ9HZCBV/uSGaftAODMk04PL0OoiosWs4F872/AALdjhnJWUx2SzpfW
vr4wEem5yPv5mc/Dil0+tHmx1oLDetDigyB7KcjKbj26wBOtcz8tQlkdVvSxDTeu
yfjOPK2rwdLfn9V//Y9hHRNmlZnKKnByeUer+65eaeW56kVWNg1tuzyu7CTDZYuD
w5SL9QiNU9DfopguAnRsb5FSa/duJTNHsfANx0mG3T6JCvyK7vV/5oBdrgnMUejA
DLkzS3DzzAUc69mGwoxx6ftWZaanBCcSCB9PC/5EmoGCblZwkRoVpRODAL55dA+E
Fm5gQNvhOBBzPZZyib+y/je6mEIUU66uVIiKY5nhItRLAQAVprZVwPGSOF8sDTBZ
LYuGVUAEE7Kx9hnrqdYrBLDoY+owqpQrIv1QEHxgTEBguVC6FGW++JHcDV+Y+WHo
8VsISD02QQBknKJkO5u1SBsetun9wi33Hg6wM00B+rQa5FJKAlDnjakIGq2Gznaz
kvRClgdBr/nzN5mpGEGLTgK8sF0/aZZubCAQg6TVeqlXt/UQRvJBDcOMBoUdUOdD
YSbIHkxcDKqYG7gMcLoj5Oc6RRf6+oxCsXQJJNwaP8YjhaQHYOsMiJ+HavU8QX0D
nAEYhF4loivPcc8abj00efBBm5LfDviaVevJyYNPdwLB57mbgrTeppVPhJ2wGAv7
7EOlbjJLtTRbrN3SMgOrZ/C3GWZ3rdMcQI/RHI2XEaMwGAv2vPwH0EFUqJY04gfR
52TSKSs5OL9MoY1XEkoEFfLar+PFHg/zKU0Y7uTkDXfZVURqwVSUTT5tLScoDYO5
+uQidlAk48YcRvY4JBXG81ikUnUBLCKYd+WjPrHpQokyw9dHvk1eH6GarFNe8PxN
ptwvOxz9B38L9cyKFdNwO576OMrZXV05hbxzlJU4mRDV0PFnIlKLhas3IZZU6tzY
EPYbzuDTk7F1cZduBBhmYz1aa5znvpRKAE7Snl9ztiln05Dwv6GkZ0e+YQ2uYamx
rlf8OML5yFTJKTr2quYLipkWhRRwvhGZtA7czVQICPAJKivhLjKLZjrCOiHrVYhF
4Gc1M5/ZYa6/tonoKIKPxg9srOVi7Wa6kQ8CufAaJDoax+xfkIytRH+r4suob5yM
EHSrC2EtXWRsVOA8K849LaY5+ZH531ewx60EtwvAoyDGtBpR2fIJaLAGUNlQzO1N
u9SqOE6DxMyb3HKYR1gudCTVSZ2BYQInvoRsFS/1VWbrijXtqmBEiEOfQ9tuJcoC
X3BtSyOhWkYHb23UJSlr4ph1aWdKZIdVr1s37vVhhthtB2v9Fw3ytre7mUZ2ub0d
ijKesQ3jz4DPfu6zDKHy+vWbBKhXnMxWhOc1BM1d33LJ5ueR76cZsB+W2dqo8cK0
1aSiigeuVOdAR75SDYdH6fDTCc6NIq2vQyxYt0mL7bZWlotTvtBt6wZdkP7H92ES
LpLFeWDsF3AJB32vRjh9qoZNqYmLfT2palfPp5b+UgeSk02Zc3zWhHbG+/3Dq6AC
TLCCAnAB8lHUZMAGFH1dxaqvjQ9tonGPFHvaGTzCoLr6bv1SDQloDeDWVdpKDEiy
7tmT10Ku3yUKenaFylwA2enOYR5nUVKEl43UzuRUWFYpwwJDFaKr4APW4IOmNQ5/
gO/EUTYLZkiPbRwVfqz3ihoVeAxwbbOGF4CILZLzSvlqqYFTHlYSFspXboA7d2Nx
cMO1lxlLPwhqUAKnFy60F+6A8aDP1KZTqfQRQ2uy4b2Y7HCGxOsG7BAsyrvkOKsP
KPb1qgDh8THAoI0x/8NWPy3a8OrlNp9Sl7heB0efdbJNIqrEDbWfyIPKdBSICxRK
+47dqfssk2KaqNgYGJibX9WT7iYHJmUlY76NCu5j+Ml7Q4vFwHwnXV2poLs+WUuT
UOv+U4PHhXTZffdFo6rFc8ouqyEguYQ8LySaLkPAnMkR4JZMtA2f9Y04DVi8tOwJ
9c38Ux59KjAgbIjHYchLE5Sj4bPqRBmyJQ1UDoUfyyonlNv6Uac4xEjniHc/P9uB
c8ic98E1Ksa+OJwM07KBL0Q2b+ekZpoTAhmni6RyPS87uYKmopE14Bbh36SjSAdW
WLD8F+FcTO50RgEDbYHt25NmZugWKjk3Mv8QGvE7dbvxeSzmzxCpPI7Rb+he8U47
+c78L0LOgiW6IWMivcJ/ZFBfCIpSK1IcKtY1OzfAcdhTYYD6ZlHKVSwprDWBMX79
2dRM5B7W3vxKoy4/I8hFvcEauiqLUPEZ05NYofZf84MDuPSh/qFMMdziBx+a3Syl
8Sc7L2yhtB2QjZNVxZUaelG2qPzEF8eAs9855DMGgv2HttPFkx1mgxj1EpRYvNEB
cqIOD1+KrLX6R6E5DBrN4X5qZZpoApJe9Lrty7kXdKbZWs4FvhN3/ORzDx1k39+J
VLKziVcGJ9R9YqKssLJTQJ2lQbUyg65PZ6imhrJtdZPbFeSWq+QNOBGujvZS9tsM
MjSk+3orK6zzhNji9meoBcfD0EapEfos/fPZ0wYb7x2ThL9IDGZBVUeSyH7z2600
NLjq5BUKxPzWCinygdT9sY7kSN6QQYJwgoWo0fTi3fbH86q+ccGFTSn6CEysSElV
WphfHiZ54g8AsxE2A2Bwu1j3gxtYzkwsNihtnDNuKTXpDKg4RE0fIqs2p/tDuhYA
/k3ikPUoB8VYxR312JnQ0S0SEZHycJ/oZlbDY8zeOBi3ffeUfeYieu64jzt5P2ei
WkL3ZZ4n7cI7+KbLqXK/R7XCrADZcsPm3otciL5Ef1bhr0nMZUsdA1XvTJcA1GL5
pEQjSCWkMmXfdaAnxDdGbgEFZJFQ6i851PgJgypkKz1tyIYKN1iFHqaNZ+KZGeGJ
eusb9vD44KrFv5cXvkl0oYJkCB3q/6wKVRCy8gtYNVaLFelDB+zRJl86Lxr6D2JW
sNF5ojCgbO0T6a5W/CF+0DgPt75Qc6ei8NTnOC91adUkyRxbfWev+eelnuimsKOu
SB38VWLX758tqAlAClLQDT6GxxcoE+4Kj0bpu3By9qXTKjU+H6JJL4CDQ/YP8/eo
1ZUV964u3P7m0H8gRh/wOMkp36FMlgrAbzbKXkZRKtgHO6vhF8v5OnW42qFI8nKN
QToKh9bT6mSIXe+MaOM1Q/OBuZvu4u+ipEj+jmS7nZ4ZtQfhpckD11fvIGUjCGsq
RtTf60odABfHOZmN8SkOnKzNq19LXU+Y/FEpLoPI4PM6R9JzfGry97GZSiX2UouH
cqrPJDl2WUbFCoftNsSIPKsrxAb21eGhCLYz/g5JZiv7VbfvThTOGT8zju9e5Fih
afB8kquXaE6QlZNUEhsvkywUcRUZgn3yrj9Ha1LmqZZDXDk3z+ul6LkQ65VFXpNL
6q95924YyoLPs28ku3rR8Gzw2i4hbjFMCVKpE5GrE8NA1uM0ioVQgG8dEkr6vnlD
CUCCHTja0m1SdLj1mi+jwKX/tDhVmPbv3egY1aWNx8SYIU1vjHdomtYCVJosWYXN
WV/QflgvySqEq8vZjgydNtYgJChI6fwdwb6F4Vysz80UYc2Q5xixFos6RgbtLN9A
Mki6rUHLEimYwrtKdEuMYST4aUjKllXCRws6FupwYxpX2K8LloRbAh1/0J9crsIA
JGO0qV5AzwClBqbw1lUVQ14/+fvHofzvgmiTwjQuR6dagOvERt1w0O3m9Pph1ZlB
sm49iMrlB019v/2emaGbAXag9S8Cc2uruZVKBObkz5m+x2Z5qS4CAfb1aZReav22
GNykP5w3aHfhpqnoA4MCkJ+Avaqt7/5qFETnf3Qv970Y9KNPfdubjf8WoBeq6P+Q
KhAtpLgype9ae5saTSfCmtfsZrfs+OnMXdenEyQyUCITB+VdOE2sWX8MRdKI2SOu
L2Bv5M/DEZcetAk4qu/B6FeZV/Hrm1lwnMt3hrKelSN5LIeftNBB7APMBeZ+Mzei
jz5ELDF4c9W2XTH552GAr3z+Uh45WqCvj6C22iVk0KbO8PhS68VWCU0yqQ8AuTLO
c6LmKsq89A9orpXNDbWUVa8p9QfTDym9V9JV0lvHXOU2X+dJ3T2VrKDf62t4I79+
4ueVo0KXIfycXnkvKeGOGS4wc3YN+nRAjyaAz3CW7IKOZC4TVozN7WpRpcC0vEco
Ocbuv06zObre2PaYgiYfSivgOrRRV8Q44WNC5WaB0/m/1c0AQnG3S3wTVfqHXJO0
59YoW6dO02ghCiCz6k0/Gw0B7TJDjHBT4U9k0ojScViQwT1A1MQBkKriCxgn5nc3
xcFKMUkXu4B1RBqDuQLIIpcJp5JoRBRFYi77B8tcA2ZEKUmrqLJiLbcqLx/XYW2c
rkGUUt4NYakBSHmkDQOj5SUU7Y/ZlcnJYCjGfztumvBKR6t1GlzAqlGdMgxlPFED
+4mV9Cjvczp/5brNNZ0uPMwYUvIgxvknJhq09COfT4T7S/lvStjPfgm4j6N5ZIiZ
cS49vZtGH+ZNp8rRIW5Mdusrcde6iYCCS99rcEpeQOXPAr38ceBTs+7ZoL9hkuY2
2RSgJNoPgG0RMPqrZhZ9O006ExZPvKYUl+NWfbZQ1IV5q0dRCi3xImjXRaKgvzRi
+L3UcaekPu3BGRbq+QWcU9vwk7oGv+ASp1YZGbE6N0B/5kYY726R964mllmYXx0a
nupdkBhGdNvq2HF8QMokggUGFuThO8bVb0a9tT1Jf6iZNch0eqaFL053ONHdamXx
QCgFPmvQk+6uZoOFRwzzuDbjwPWAE6uePohSZyuzjL4AaWnaXFlAF3VghTZ8ujUv
/4ZUAjUxYR6otx0Yrlj2bnWyTQwObEUYgDp7rfamLJ8F9yr94d+dYLK9QlxDz+Cj
BMdhBnBiPZUuAexsYV3ylS3xaPXzVKJpj0rZMiaLf4/N087LcfsWNm3H/wr6gr8E
QPKtXM+Kl2QlFke8bCJRZ8rZpC0MAy4MEcc6eMqdx7Yxh2g+Wzpq7q2ff5KW+5v3
cP50p8t8aIrlNU81dlYUXTTQqhuliBoy+ndFqvvb0Ss2MhiCon/C2cXGyb7DAHt3
my9EA9IBal+nSrYyKzEg5I0SSgRmv46T+4CX/0fytplTArO3CzIJ5GX5QozRQhee
BK7+KthCVDAiiJOJXu4BstI9YF0ewDaFS02dHLcBj3k05XIk+4CGPDfoqJ6UAvct
VK1aREUsrylXa05PybV2lJtnWTbyOwcuIyLqbjFDd8Zl8L4mtdEb3J8aOZoSuYqh
u0IuCn9Byghin8+nfdNAQrVVf+wTW5Rbo2uZt0jV6R2KGX+9oaJmbhqhpix16O01
O71k8dIoQL5Y8fLSbF1wsqhmLYJQbmE3BiVmRfQ1sEyq1IibxYu4WYn+cKEkTE87
SFdDmFxBdRLJ3XEkFL7liGBhbtK81/MqLXDLAhV7nziNkEc03yrBggSpUe8CaHih
bRQ6XUlijM8Tr4m6/89UheJ2CEwUOD8K8RekSvSVxPobargjohZQAw6TozH8THAJ
/jEYRHlfAXFd9RXCstwPwMzsTOkxkO/u/T0yeiq5kGZdF9nmFv+DCRsZoQEa0pFU
6zVP90VQKNll++aL3uIMljTnwSEUIXASpJRbFipYWyY41ZLgMf3x+ie96K/j+JHv
aosTtEQD9urt+Jop/5JprkOpDogWfsB30e6tJekJevpkN5727oa+NiURwc+Z5MqO
PNd5PlH0AO7Sowsfwc24PbTQoBRsSfgSSZ16nj4KcyW5OA00VidaSX4EiFRMr70s
IguKsqtL49S67gIxWsVk6jnq9bWOzQvSdLijbqItdztaL3J+NpTr+Ro1s9BsYpEB
977HOW0W8mqNP0VevdfOY6nbuSDzFuu3BJ/IeHaxq8aCxuxO2YBu1lVO9IveAviX
cAKfgd/GypTJlLMK3jZVIDLFP6EZHKK9sYivVpKrV2laQLPmmHY9kgUToulbRGVI
+VpCmvEsaVXkxOpFjNRr75ySS2E1QylwQt1GkeH31iFZRoamSTKOro08DCVwm3px
vjA0FFcbAsAxczMrDbyT93LQ/SBishnE6A/l0I4sVzoy/84l6C92frWgqgG32njw
JkzLEVnK8oXYPwspqBXBEuthpSAIBrmmxxcJA9PECIfvpmnU5G1yU5rWnerR9zG+
nL/dM+byR0QNDDeuNmEHsKXgX7BKPM9XFEYhzmMRNusL9qSNEES2cBpf9xVqZp+l
eWcPWFAKroylCW9pX7Y+CRXTr+g1zx8gf+E//dvU+KJZvviLjT7xDUgO43F3nLrP
1ZA2VrP/a2SuFsavvXsZyJS4hRu++4VLG4NgJZ9q8nu4d6a6se1yOjyPWwynmumm
eM0BS3slSEeJlVV/+KbftpX9jjSkW3Ox9m+kuwUXzpDONRrGqR7tDGn7fJkluzuJ
zM7zNJxCEWlgmvOHRZWQ6lEq4vPWSooXxiMLZmGxVEeEdT40mVphuE5E/Vx3ezT1
ikNi9pqQX0jYPEPZCKPrajnz4BwVFiduC+DCXh0Dhr9+4CmDDwc32UDQIHI+/3ms
dLMPN+Ql9x3o3zA+cw6lluWIYTzx6SDmvTSUYmG47PWbtOI8nMHC7LCrj/ZJUdzQ
EcYtoXXitK/cgZNXrQVVZ2Ek41Q7368ul8I2+8V3XRAUiIVUlsevv1ybkjVm3P57
0Y7aU26qm6PmGs/rrIehP/s4AXnCz/1XbVEYehu3EUNzRTeA4pg/gHoLOb7YQ3/7
dfdabXpp9DQLIImwMDwM6umjl0sA8S8E+pJJhOEPM8jXs1nKwOK9qoGqObWrUVAH
Tzf6pzjTd6jX+8J+W6Qde4/dMcHvz6SJWsPjkbywBiHL2FuXBqy5vlgc3yPD119X
xBs8RPHr63cJXskW8PZjQwalO2s1T9vHX0Jp1FeZUp3Vukd2aq+QH7IWfHoWMHsy
RQzzwmdBUrkuGruAZIpVpGv3rP4TfLsetFeyCnxON3+KVBdXn3QON9bX6b1Hg8gG
bcvhypotZwlfy289V6b61nIqlJ+gNjX2AYV3Wd2S0b6ysh6sfyqzi/fOgglBcI8u
jSUVX0Lb5SldOWZ+5ztpp2PlY5Vtia4euwWzwnx2WRy8/gOVq81IJRTH4wMXeytr
gt6lUq37Ga+CsO8Dm3ku2jUxHXeTnqyyfUEn3di6DskrIE6U0N4MZgTBQ/UEEsxp
KM1gxPFu+rVvYCq2ECirMnna2UTepFLxrATDTSum+JPbem+iGrBqMvFr2VEnaG2A
vDL3YDAh5s4rPGkXv3rpzNVtrle9TdBTMEt2G0b1tsYl95simIM2fyQ6HtK0H+O2
uOEgqjK6H1raJbkPKPFoeTa1rMavoa0jAf/xkVMq+kP5CPp0PBT0RLc7tVw0fKsC
L2rraqp3xgvPKWIF1c81nh21xjJBfJ6Br7el4A98o8bQ0jhk6pm37gOmyKr/JIPs
JAeDr/ra64WOZnAw4ywYBh9H7Fso9Ig9vU0s20RNhlasgFuzOxFFQkk7qMNJZG+R
zCLkGJn1OOJHU+2VizrwkltemFdPvCC9PLgGSO/0VIQ8uwIukadXM/ZIZAHER08U
Ain3WMotLBpHH3LqEoB2EUz33jM/K5BvaNjK5r053xytGyBpCM+c+mYgosNn463V
r/yK9XDc2qjumk8hzNsAC5TqmJbu7ZRGhvKd6rWJx8VkRihVMUaC0UraQtNg/8/4
Ws7X1imprXOfgefmtmElag5OJ6B1HOpYp22G7EagayYVBEu8MuRGcD453pNcHoIo
9GI0fwtV5xYvJd9cuXv5ixt+bMQVEOSAo1uGB964DCl/Iqz5QGl7T9lAvzjxkppN
CU9ZzqBw17YN5zUGr0QO7eaWUI59jGylPcSkeb67aTFAD3NPPlgHTe1idXcRZIPq
X3ENkRaLnVsRz4aS6BlWiw5a/CjlnXbooLs/19+n5GFemoXCZU/Jnru23y+7iS+B
wxt9aM09IfF8bWqIU6GWOftLEDqXUYFyiXgtG1d0M81JyOXZqmxSg0d0Gx9JutE7
KdwOmcFreFO1mEGZhn2nHd1DKxkEK/d2Af5RNSj0mVgOJRBZ90adNTHmPTPat4gp
jrVgw4SjMYuoItV/JgLwhua2ZIa5tYGjWCmSTNWmQI/6nAPZwyHdB62ZaLoJqIgq
bwCtGwvKfiGnEUwgll6CBXj5E0/ZxqreECStFgVxoVnKkbmtt2KpRARdKKq6jDlj
LcmjYLqRbBJjGuJCqqBcsdWTMM/9gMb5dLb533mYMIreJIaPjnXc2av0xISV5dE+
2sJHvPsiCJ3x8EFFcb05io9Ilpq6eLM+5H5u3cBjgaDWlZjxa+58pE2UoR7U0zX0
+JVPtFvDf1D8mK0dz/CcyrbTBdWOmAQ2C+Okurt2KBgnmLJoWiPpqlYAGGqiah0b
B7FNxmjZ5A4MF5rWgo6yB654o4gsT/THSI9T5xaIxqXITbSe+M03T0KEN0bgGKpg
6aoBoV2X5t3pvsUghyR/i9QhNg+5MtDt9V65kOlSNyW0QwZa3KMY0K06VNbelyGY
IaD+jZnbUc4Lkf/1QbF2y0apnjlq2fTOEvjciYUIwVSArAAyNzDzEyN6lOJ7sTxV
MlInebx1QbeRotFHmXGOQippCr7Wa30M8yo6c11SfIEh3xc6ECbRvHjDhsQGmI5J
qWad4J0RpYaUxV4CZVqmJYaNIKfg+3mVyLJxSl0SH/d92z7sizIoa6LpoCBG4D5R
BsTVunZDqWke0BkPJ2pyf15yHhlXWbCF+d+AZ0zHkHAz0wHN6CB8xyaM2t8YBoDz
N7n1QYK6M5HmDihpXKQnLGVWPCKiZtZlkBn4PXpCwfoaG4vBXR/nTCU3zBvo67Xj
65rtIe6yznFcu54py51YMntQrSoFUQbSg30OJ/1uDFRRV3hV2lyRgWCEmmCC5oxD
Krym3aUWjY88NiQe2/kPS1yNHfiFw5LIXVDMOY3lCVQUXa6PqpPKmXDwKSrDBZY4
FWaPhRueBIn8hR1t5Cw0n92MS/r62z+16CFS5/fMogwiDljtCpQHH8MXY5a8SX6k
3zTTVIDuNHWQDuoR9d9SUgW5KGhsrf0BRAndxqzt35d/vBl9mB/PvM1LXZK+k0Je
D2PUUw4BYTZHvCtuG4+2QJuax52YYkFxrpDJJj3C0zo2+cLznRrs4ycTiPQGjUjr
79s4fXYXq2tjoUpB7+a5iVhlzXCNqy3+dSmI1aGzHDY4kZocyeEBZYAwUIunjEnh
26yz/aqYIIJlOanjaJ1Y4CiT+Jygh0i9M5swCocIEJzIfxUrNhb+fc0LGPV/vdHX
W3UkcsBP1Od+AjEt0jM8HXHFow+n9C85ot/zEIMDqlV++qUt8k9TIzxLEAFSTliF
32YxsfmU/FIrCpQzDIbXA6SWdbLkiMtKjLhQMxKP5tADXLUJ2ihE1lTrLWR2JVmp
wL2ldpb8T9cHaE+ZuXi0t7jR18tqMc4fOUltc5fOQ4JR+yB6wOBEpmDKRViUhJKF
SwMufxcLOD+pZLa6okcL8gplyYgC79lyucdg6QfKPF2NBdD4cDitW0rgPbjHeqVR
1B+i0YNA6U8JQbZG1e/bDNxp+8/6ov8YYY5n65ojD4Ko3B296chI04thkqch67f9
Ug4g1xIjqfevuwGXCT7jEi6K4Vb2aYOzKiv2vNBGTxtzQ56JuSnRcnVbWNJhEn0+
r8vgD6LnFUjTgXQk4QYANC0sFwZae/hZRNZprFuQpzR1C4ERHbARMrRfasrEhlNM
nKkzCjSt5cB8HIOF4Vpi7+/OnEIdZLlEoUqjXGfrZt817pUJJt7iofp/wiFUDLJR
OUXhvtUppq40ur/R5zG5w6UZMkG5I7EL3PDb21CUFEyQG6LPhH4M0dlYHk1WKgrq
Ji9us2Ty1cueE/BURx/30+5FMHSfmnGZfMFOSGaG4qdQFAc5i4uynX8c/kbtycCD
mfR54C2ClmDTZV2RsAMuLlkEuQumprml7DDZjHRNSGFlYduu6GDIgpKDInquawvC
EN2ouKax/xaO5Gx8NsVHc2U1cxFZsiW5h5ermNiBFx3SEzHVoHhU5yCHKjkEhoYG
jLopxDSqe40hDnMfQWmdvfOzqaekiDboopMq+2LaoFJAEZHcraH1YNfT/nEChYox
lKHr/X0DkvC89783KooDcC5rCIJnpPC0b0ttd4RXqoAVeeeVGVfTOVAxNt9q+UJm
487woeNE0/lGeHXWmGakfP8NbGqmPbtF/AjvPjg9PDtosUW7c7p4oU8qRB+8iKWB
6demI04vNdLgtwXVNP2GI/bzecEr/hm0J3ETO8h+Z0WtfkGIg688QE/DPNq/vGT2
q3O9wtCfWf0pUAl/UAr9y8rat6SI7H09WHvvLc5kw+u+P9CIj3iWyxWEGBui+Jad
01NK2n+CnXE253BD8rv3YxmasLemmtlf6zJ4qoleC29JcWUj+nhvgbKu4eQBIoBO
8ERpJKwO34BouuBzTMAZJt9jG+Z0wTq5Bl73wxT3g+bJ2nTKqsbNWM/7T1BpbrZK
UJ7ypHUlm+t4+LJhfdxuvWObMV2TLk2/f06GnEhtkd5ZZA7UQMAOLZLEbz2RXM/t
0QoNk7REP9MwxpIOIzv1y9VN0zqbB5TsHeLq+N1AQscmJGUg5S+kVbtJRrpBL2mx
E1nSm6Z4ccMZBIJDd7/CuChFFv4v4bQZYYJEqrWu7Vbc6xYCmX9p8kkK1GCOhsPS
ZpDgf44iuTn7CyyW9QxUuJvBCJEA7C0EofyCIYAXj00PWzUuBgI8MlPALj23AGas
GBbUaK/+b2ZZ+5QQ6YN5kM4i0iJimTsA160SuGfnvtEioDuIX6hotKhKayCwrtkM
DfjrvRK5j2tfMddcnCvLBMmk7WaM8wz4ljpgrVci0abpwq9gaOhyfnu0SynHiWd0
hYp2vWStSp6VbO4N7SRv/i906iMonF0x16STsdQtYSkFJOl1VwsHTJxkoGuH9AGh
0SUqO7TCBpbWsggBjLhKknR2c3T64oceAs3vJrdmIu/kT9EyrKgSc2k4awo6BO+Q
ZlcM1h0nMXBMn1jUoXdMcShjYl6wB/sYq0A4/NiWMgrK3urEEfsURiOx5AWPDqQh
D/p2YcEtTi1Flxbr5pVEJaIAY4+4koiyEdC9vylpgM9jdQx/HdYZMBfYLF7jTHF0
g0VDIOiBjkB8HdMakDYFT+B19cr6rtjvPGxKxjU9eBIfa2DWbdoywoqkzlW6i20K
oe2+Nw/PbwwSoB1M526ZZNti5TkleEbdY1qu5c4xEyC+Buloqkj7gntdGR0Jgfz2
eZYtU/boZIyB1uJuvt/Vtq95g0uD9GHW7GeCX9RxgXFicZwqM0d4jBeaPFbpjOWA
z57T6Zxt4pN/xtumf6LJyCuFH31ZYyenHFz7CRdEEuRab516NzY4ELu+nD/VC38G
YIOiCAzPdVmJNRSHfEOH1h/TWBQqfqhXedbThU4Zl5NX2nk7+OAtnSZRHK7EflKK
b0gJ9g/Eix4EncZRTSlCaCnr0LhWOz46pPNwgIRCNdnRTmLSp4jqpOEuf383OIAS
vqZpnCNgMqYNZ0DSwbnsyaDV9vcLHydlnBX0oX7E3yNNEfs7FdFNtbOe+EbqW0TY
h0wRsKtGtf2WWeFemv1AbxfGveiDiclBzdM2O00sPMhC/NNo0ciWF9s74eH5nlpO
QCg1at9HoG2Z4JgDn8W6jKv9rFtH1CuRhwFMXoM0YzS/+bCq20HtJ98GLuFkI4Mk
QJZifCaQKsPu58CZ+JvNZl6KY3V1oI6Cf+OFvoIZDE1tTrbX6Fn9j4opLraqQC27
byhszLyWRaRdNXlh8PtnCzlejc4RSJbCX5MJ6vd4hTDSkht4GErswQkYhtIgmkzL
iRswlbe+clmB8DMuWm7tFCeIihYyJjg9tUKHzwE+VPE7ZdHOhqzBY91s3JJmCTeb
ReAc6wm8/x3jlOZW3nzQ8OfsIvuhsK6qo/DZ4TA4FsdSpcpRJdgAQlCCvlvN+V9T
IwBCqsq7gBNTQNv8LBxT8j8GCFUzlMUPuCgaar7NfC2Euv1nvvo4v8cWLTL4BWbT
xsizFL4QLvJIVpzf17efXA30klqtwwxKgwx2bJiA1dEwlWh8E3RnhHyOizZMR254
1mliJNjTCqdTsjssYm9mDE6yrs/Ew+FZuhp9VyqOkKssu+JCD34Q1Nifqw+CvoCI
9JsKdZIucYDSHt/5cXzRLqcndZbRquXDgPSklXYHFWdPN0nyUyNqEGPG3ujxqHn6
ORXec0oxaW6/0dHQwxct2w2SBC+3NittpntQgQ57KJ+EeD7rbxDwCK66851Op0vS
RyoHhflLxfPvZCnuzLt+eXGAexqlcw7PoFJbItNi/k0Mcxu6ANlwy9ECfbVumckr
VBt21GhQz9TcTMP5LwJPfK+ju0WSFEE/1NpV8ZzZdyDii6yY+qkLN2rRjSoSvwi3
VXYvTarvKYh3Ed8PCSNLjb2ZLy3vndg+nCcoKe4hu0+eYo1EXiTf94vXYvpVUfqH
aDMFqkcUv6V6FY4DEvB/BxOfnD63OAzAF645IQIHKkqDsbmZVieJZY3eO3xs3KqA
WgNqnss0W/0Gz89Wj6WosZJUvocWnQhcTl+XZ1iZeV9hnO1T5fMmHH95/biVFpt4
x8FkoN4cNu1307LO1vCEjZmAb3bSRvepkCMWTtNSkRupombRFO0t6FZVWi3zANuN
85sv1F8blea+19738Tb24P4XrpUEBszUOHLECbIRfqFH6gUOPzH3m/H2L8urEyER
XXvdl9PBAs++fH3gv6X+Qi2o2ZkZCgImT+25bcXKz6mVU45CJNyfzNfG208qNGlW
o6rfAqxz0xqHLNqnFoCxN7xPv/L3NaR1sVqy/ZyVxnWkpHr2SXW5tKj+GA5BCiUl
liCIHMtlymyhfffGC3fD3v3ftwbU60aFsafCvuQ9lT1VKJUD33OVYQ/XVrmgus6q
JaxOrXoZxVHU/YKY9rL7f3UxclTNNJEbkZQ71KBznhIPD7g65Zw0mn/dS5V2T/1J
WGKMOwpXgVMhhwhPFzDqFHGdfv0C7AHvsv9LTlHt2L8kuSKPgRHjynnyKVv+Q2bm
v3BJ+5R+gJ4CAVHhLaDTO5xBUFPdxmQk8glvbsSIJFpO+vUPAmH1H8qc4r+rxtp/
EH2LPZ/uziRKSIVsqw2EAGZuviBhHSQXQ78gtZof014tn6BB8+l4CblftQm3U62J
hQcurmPPTEMmZx8wKPYKQ88bdaq/PjtcLDQcJrAazqlGAUREjaHwsIt5nZweUG20
Ve08Sa36SV6lItxHbTP7lmBkDfalRg1nNzWV0392L8PZEOqm5KhORu+CDb31A5nD
HoPsn6LdHwkLQZZkXgj1/dubMGPvNpniszp5wyHhTnRnOnX8vOcjDADdPxHTIvSL
DHzFfzOOdmkHRJGEuAaCsrh9suIKdQvw7ui+//h5aW67+NYpAcB0343Ljg3wULIG
R44xFCXgHXwbQk6UY+C+9nwLu11IWR+OILmD/Xdy7PohW5fs1G0TYdEImXenk23S
ug4+sT8B6y45fsKkM99ZoEuALys9pregPDexklkzzYIF+jk4zyq+Ob+ibcU6c+eR
tcYcJsdpl6Ca9K5E8z0GNWQs0j0vy9wgW3NV+28bae2TvxxodhUvrc0elfiZjLaq
k0raJ43Hu3AFxmlKsfZiEpn8rMeyBw0ROpjjq0mvQOG1Eq1+64iDsvZP/xjw77E4
mYHHidxIFvoY5kvxFCFrT3Nb7bOA71C9ryJSIND+yhyQurWaOwR7e0GyUNig5sgq
aUOkvuuwJlEKdai5F2CdbE5Vo+JmLd0DEX2eU/MkNBDqsm3MNHFxpejsQBr3H3GS
qXy48E6g67uvtL6tcKiaCebpcNBtxip7vCwc5HIuLqgArmJQqWK1q2JFeoPjYZrl
9Wlrffw3d8uuuDMGPF4HA9oQZZKds7+tN/tnlFZHGBm8qMesxBvViu8oCFrUxyuC
UFMaAqkMQoBRMy6DVxmeDw2by4LShdAPDxpl12gSAzMiSS8tS30QfZChmFlEM3o/
WBusPApW4R37Ea+R++3i78HlMCHoAn2QRVXELy+OADFjAr0SRiOeJy9pGr+oc0P1
wtyj8UduNPIQdNX0FmMMEXDii8/XvYDsuGOW4tnGAXR0rYPNXnuQBnYtGYXO1FO7
VrzuXrWj9VDGEh8T0SafWStwjMC3hLltKlBsELcRa09l8XS104+dHkeNXUrX+Uue
2/uEOKZdpGGecAYkFJgK+fttbUQDSAR4U+sm0Hw4iW4qtth0mbTzU4z9UWZojshp
bk8EDrajaGqqywC/2D3/zMFYYv/tWbK/4BPpE5z9dTJ2u68cwmVgBTR2t7psIuzy
huR/f87of79bbdHsbfbUMS1qmhxyV8TIkyokIiAwrO82S93NitcIOBViodURKjGV
scAAGYLKVgC3TMMJJkUEmGyRlEpgiMdrmmEALn96wx1ARO9PPZXHcH/CeJ2DGvfp
d6mLkGE7lrXWsr8ST+Xnseqc+0z07c5XYsq/Z1v5oM6OyZyWF+PFmnp0Cb0nNcv2
+CcrxRS8qtdFk5gMMpk27CW1PE85b+zHY9tmA2rxjyqphxjnZbiaEm8j/X9YF5rS
KAYvtOhOXAyed7tT1+AAb081vWzPNxiF1wdA6gHJAr4E43s88JX7QUUvsIDvLwqd
RyPMFibQYkEscznRb57iZhhYxEM2DVueGZUaZQNQdmWJNYrlIdpKH5fzEnyL54aS
NEPmSRwDVJAuDH/5W8UmWInuuiH2tG0n5+x2UKoAIb1Wm9uiHwmqcJPsENHy01U3
Y9wdvVWJyG6hVg48T7HI2zCpF71c6cGp0L0ssRsHEPzCZpqdUQ0OJ/8my0IbQ0Y7
+Pdn4Hd86Wtc5wuRMo6NjZOXGGYSFW+pXYqy/L7JEp1x524ExS374QpSWMaibkEd
CNrYhdJcUWlBzTz3tud7wwEGubAMrWdDqOSPXvzPvC9CdOOfBOOgxvup8/jnIJd4
bh96UO2IwD7CtgJNLwVE4tUM5FDgUGqPTp16W4/FfYWoVmVsUILiaMCE3nBRtCoQ
9nambJruPwjol6slWnrZduoD6K2O5CllSjSkc2p4MAdV/+RGhCn7irPveM9OVKcW
khOKT0iGKDwCxRq2HY8HBBIRzLjgHU4E/sMAnZLlGYTjG8ZkxVlCvelnLbt6EHRN
06JEjaPerYD1Hiwk8XoXrQrL1KQuiT16t1PAjZUZkXp4gSjGXS8wAbvOr9oEKsvn
x71HzYu/mfusbQXIL0ZhpJBsgqIU3znayEXLegJFwL0yDacfx7sFbaO8W/+IxAYB
awAlwoFYW61zILOvegu4qnH0iiM1Mvx38pxjmF4/pymVHFN2pbogPnWRk7SBT0h1
oY2kgB/VA2+uOClKZ97JLlTJl1R+Oc6W+9bpPQ4qRq+PeJBbsYegVvmT8zXemc50
ngrURC4BCmQOuz1ujQBN6H4Nqn9kfg+uLvuhkyW6WNzP26RDBnjncx0dTOnsZnmN
TeOfPBkT6rKg+HgbO32V6Au2BbIQsxsJMS8SPCQldjA1LggQBhqZlmpHdJhUCdJ9
D/C+FK+PSQOe0HhAmXOGVPLb5JCHc9tuqFyfrpXjlXETNFH6C3fmo8UECW9pOjBP
GVJJLKfQ5l7vMM6BDG0oydTKMnGvxzk4mwMlOtQY8hAKUTesBAT7uAdXLs3ME5DJ
BycfB0uPfZGCipEIIpC7aivDReCe8DggOsr+419CjS9ozY/c4TTzkNuBXMFcV4xt
CZgNCC6FUCbxnsPUTpabZY7Fpm80wMz2imkOsmvQUb3Ob3O9V2KjiM9aX2rsJpIB
IXV5dKA4PB7IFJAa6rH2TmVQv1LYrPGMZKFf5g8QdKKI5rHpDq+2P206Po2JqeZi
bflFe7SG/1kMp7YmsQwu3+x0lf6I8+oBWBhVE1PkI2pzn2javNnM/9spt+KdvO/f
VmQjn+j2Etz4NSu4+0TTKwGfI3agEobRG77Q7MoKZI9Z8QVmxHS7g3MWIOpkqcTL
48FA4jlbxvUy9hmfHJG7Kqr0wmldbAkp7Zi4UsZYVnWYvovaKbnsKzZzL4ZxkoDu
GEPwgQNH7oplI4r3wt/BQ+elVqhV5PvltMUA5a/yoLkihzUu5Y4iA3eK2i113wSh
DWXYuYbcR4qOd05dRAGfDmoGPiIj4eyHiXV5mY5sOoNSpiMgdZhXkWz3m+WTWh5o
2u89SVuAwgsR3Kgn9QxVMWUS0Gq+iXsZIheDN1lQO2sIWYlAxrExgMH+yv9H58oi
qFq93ED/vDUch2kf1nFIvmbpCBKd9JWTNUYkioqMoPH2ksuWTBYSjFm3lX0BViA0
RXx4kyE2C7MuL9Yq+yrB/cx5CEbEi5YfBLWQLNMFMIeRmg0Wx6rcUvFtDLy/TtL+
Uf9K5Ifs8KzjTWv6cOmorxhjo9nuz/n/CqSE7jNsO4M7gXV6hoAzjR/0Hg6AR6dg
d4q/z0t2ZjphY6EdGXPVXtIpY7tclf2jT3g/gDbrZKszV/Q7M2ehCk+SUxN4Fyq2
Rdp466heufLiR4Rd4abnNTUEq8vZvdG4lj7n2f4LW5dTEKlwsuLhff+7HIwaX7QA
SAyXvrNOe0qjZvZ4c8x6xLKtBFwDCTzvaLgHSVI9cIF/kGuouW6PWyeM1rwjI3UX
PKAk1w0CjULJNF8OlLIHW/iJiFMirDEi/we5GTOa/CEnHVQge1zdTMHsx74V4D/I
2PTIkTuvOwu7Thki5/ZN8JngT4jETz9t09ahy+cfG+S4pjaAW1aDlKuNUuSo9clT
bygEzpwtMyJWN2o1o/zJbBLcT7y69qwR8riOZKjdwN51aP0TLq0q58dWBaPYPd2Q
lJJl3CWoirKuZtnwLGTBwXxVgdjAc3WDflcCaWDMrHy7tOIavFoqZuQW38oMslnQ
3rWTzyouJvT4iRP0NWyQ+6O44tmDzGi3F3SJ1irOUMdezxX+TvHUHMGhACijvWX/
NlTYsm0iLN8YUF7V894/vxYog9B/+BRSnPB0RAyklztEz8bObrNp4ChMuPvH8QAF
fPho7A9LiyP5Yr1+QluGW07rv35uA8UZaZ4EYEEVrXqOKplIQoS7QXkCvpHgb9FD
Y4914ISuJQJYdhX1VzVO5W5ckVeQF82EfJH8aQtmmX3GaJ/nEod+kLcEo6WkWgDi
LAKsuekhSSjRaol4TzdRCQdcQhiGPw6JmgB2r5pURkqy3LegdgbJdJfl/Qpmdlux
VvQdpnupe7usIbHVm2GtHUZ3bNMc7VzM9W0kZjycK/u9ZYF6OMzdW1KZnsov0uZf
HG7aZ39f1qOe3N1A2ORx2NCuO3S8RCEBu74LJFFO8nDW6zAgSaqdOW5ZBBEjW4dZ
ppcyzArX+Y5IqiAOmT4Lj8IGEuHrdxe8V+SxuPsWSBooz+TT0nG1l7O5XSIKC9uq
OuYGxGxJjO8YcuihVd5r+an+I6HFq+aKtU/EhB53T2GirJSVCUwkuStLX8QD3xku
VkROmeB0wZZaZnTibs/yRRCBB7ffo0zcZnE4oz7GiB6LFq7KnicK+9ntpl9qz7KD
lb9Hed84p4HGFmVlW+ceUatN0nkgHXitzDgVTEILcV/CyM/yM9VrTJ59S+2i3BhS
D64cls3vw9DO2vYHyd6FOI3n1yt5n2xl2ZLmroMmxHRtzFk+5PBbhjIH3RjWI4kw
ySzbVXTtFVsNT6p8iPdbyZ7+IM8LquZ/+AfeAiPYFDCsN8mCSpAu9MzKI5qOOYfG
a4jbtPgj9iU6JkQpn8lKeNzgsEWx5zqW43kaHD1hHgDpWhzE+gPot62TMBAhBrJH
aoAnPZekaxtbIgTq5k4Jms1+Wh6hwkJe40L84MgPG6/6z1bw8vrgqO9NUq8C5GXn
U7d+m8A/TDDC4t0kNzaYteeBtwl+DAejvoaMcF9D+e7xA7gLCpF11qtyaCXM4Ga8
w4HtdOyndQzZ6PsH2qrXMavKDUVpfglDXZqohbt0cUWMSW8REelHaW0S+QQNJ2Mu
yHngFTha0nYnUadDCg1mGVb+k9JrAjDlzNWtvzeF6W0sd2rl0kYblSfG4uayuPdI
17ClgDq6gj5qz2kO8mJ9nT5f2+FdltroEJyd75pZ8PngXFYMpZpNfxE8o73K2Nwy
pa+hzIoXXkPTu2c8Xbh2agQHXLNY9530Xla3YPqn5UD/tcQk0IPmPOsSIxxJZsub
ftYj+UYZiPYLrGucPNlYM9MuDDeBgjBFiFV1hSgdyMjEACtNgkZj2R9kpPLnHoA1
He5OaKanjiJAwzHxnegcWbo783GqR4liqGjZ87aboTy+geQgqxW5WpUSGXMkfwOw
Wi1zHur7UfiCY9YNuA48cpuY1Ot9HAgT0cYswGhRMiEkkEMb2+abYESFLGq9bPJh
k9E4kHacop5J7dxf6ihCCl5RpcRLIBWu1VngIwWsYcgy0ZBOjYHbaioHSzm1JvMV
o/tryrpiGKEQBADsIwpft7uziv8oMW8tHK3nT8bQE897cbasaqSfCgmU7s1qlXi2
+fQBnDrnZ4x114pTf52gRXjceep528w+PqlSZqHf+f/+pRrVkuGusLL84VSh6hjD
pmGfzjbZFRxXABFser3rqsyWqHoyddqH2mBqFr5Wd4yIxjEvk84doavr4ChMtIiY
q4CpY+1Pdo3aehDz4zIJWWL/z9hLVGN7Sa1KBduHeRpqTEWEqscgA7NJwikb9Y7p
2hUHFneYaq/G/ZXjxIau9egYN/23XzMmLtZmrZoaT0Mie7j/5MHFIBI3MX8NP4z6
GiF9OlL7Su8cW+R0K1Jpr2XhUF/QnV43An1+d0diatjA5p/qqsCF4Ju4hSTHKnC1
ntKpdIcwRGoLYlZCPS3P4VzCVpnkeTIddD7rQ/QNf7WuSJ6ehmHYI2MeCXYrOhVs
bCdQR/C+psC99w5W5x7E484xtT/5OfrwgACfVwzVBja45aivD0MTapvLpQNNLya2
FcyOheIUgAM+pWkb1A6Gn7kGxr3isG6wr/xNoWj2Z30jxHjkEP72c/psbq6OaIBg
LXvCqYX2amRc8jpj5gsfgs/ZipV/LNsd41NkNJ0m157d+1ZAwJpxXW9e3LgcjBHx
b8blolYuutdv77gWBr1/73XLCCSdpIB8nHzvas4LR9lrRX2FoVetxbg1TkbTb7/h
yhjQgyUNXOW1N1KhJGjdvE0T0EKFHgI5MMA3MBF7LLF/gh514/fLhr0BJQ5ej6Lk
K3RtfzvecRzB+v/6pH+47uebR4bbKIz4KMeLlRPBboApL7dKg2Yiq7nb40/GeAww
+OCSSXPc6YlgVbKOLMaLYMI6N6Va2sn4rrDOey29Xe9C/AXtCyb6Rt4NgOb5s7Q9
tIv5qX9CqWfmR2KCLLf4WgZUG2VpJyZPs6BwYnSDoLIPyWinP7e/xH7nF6qfkjBe
JMKl4TuLqWRemzbbiznbQj2PT9XWts0tDjj+N7TtCCfAvWOStzOU9q7LxIOOOOTp
f3RUJFJLXZ4aNha4HpvFvrttMPfVLyqmGS5CDtIizxO1djh8H2KpyjrD/RohydkC
NgEVjunzzybsmphdy3vqUgB8kt1i5gDRHtgmH1MTc0fro6r1OYw030aL9z5og6le
7dup+RX3i9XUMVkQhI8c+ogmMldVCG1Jb1wWK2t1JFBr2JLZ3L7JUFV3ldKZJFTP
dvAsugw0a76aBnYosaisiYMqy5AoZoNS7/tbE2Y9jVqLVlWpeoKgUTk973mLcTnQ
/1Q5BzO/TccQixiJFKNjRWrsbHI4OyFgroVKqI8X2pXT0vqGj+5yrC+eFt5pcbZh
ugU8mf4TjrTqXqXlcuAfbQ/nWYpG2qbafP7yzkvUstVvI7yg8/lX59cyxTPFiyEV
znp463hOgTM3XEtUabpQ1Z9eBJcrNF3cPwFBmxGTmSXiohG0xRlp5NX+3NqlLWZt
H7CvabD5gJgKGBV84PrG0tVRVgkD/zNipzvJzfXMS9tGQ2Arx0F29LCKRSpLN7kQ
PXIbR73iDcNaMNtmpBVxFC6t9Gdp5uj93Zgi0YbRk4gDhFEnSqnBIvbEU0ubvk78
WVDVQXmTg+l+LbfZLDUJyY2CVhmQHd2VllMbXyqbHDxEixPKacMGdpocRNVB9mw1
yq1Pe1uZ/SfSXA4G4tfPiWOi1LrjB97FnUk+3MINgTFhQqugdPN+QNdCRTESOLLt
1fUsxVJEztKZJezI55p2PfqbmB1NMl3C72DRJBdK+CsWFYNSXn7xq1YVoiXbGU0L
CRaZsvd63wvJtVODfDasxOYMKUvemDaPKrIuArv+Ippm9yIIo05symmRaqh5P6aE
1d9oAyIqFovsTMiSDHpdfUcaQYu1OsfSgns1npIRhIOsC/8wMH/J/W0Miz79Bp0i
d30/1iVB1HZ5t1JshkOl3qNZiu1wyX0e6DrAcyc6NUxhvHPYqW5pf09y/+E9tWGQ
+vz8aCl+nOLBRz3zfZJwvTwhjx2WrgXwbUUcOrDUlXSSiaAaUvEuv+q/fg+l4sGS
0eIHAU0WqUoIQglz9JNqdiriGuiPu0mq3AQhCVrceNralYoVDicJMr4x2X8mp273
XSLCFuZQENT0hQGXE/Qk+mzA9homtKtaYYPV1I/oBKVgDFzrgsJwtzHRyUng+lfo
lIiJkmWahBkyKww2i5xtGJEhfM/w108VJh3bD80VWlL6a0s6Ew3FCvndzG9LG3/n
uE2483680PujoocoI8LPPw/Ajg2qNr3lu+APvuIX+yybBV1sBPEKXSL+pZwfwIOs
/OfiXSZOQ+Mf1j0JeuxjjMz1koKDHh2NUuc+/EZjhN8ijqVJKwQJ2ocf+TSYxr29
h2NSmfqYglNNmPL4axFAKkYWB5GE8hx2G4CzWrruAbkK/EvY9Dp/Pxi3JWjLYdfZ
2K1dCnUIQmQ0j+G7L2GbAnCdHyPAPoxbT3mp7hYcN833lKqpDMGv+oppJ5/xpCkZ
lOCIi8hF9uAQpMnqGshoc2k3+etdP4b5XmsDBRV5sus2U9q0uyDp+LhiMMmO9OdY
Q8FYhWQr0NnNPuSBNqa6ep4L//mnPcjAk5nKIIspQy3MXj+DAbhnnLelxMjz0pgw
Sy/l0DMgwYZcJtQLi/Uc1Npwmwc4pZeDoNAD0Wckjvq2/fZyGzfIm738oLD4y1DL
wl6ciqwnxTbVZx84EcSeKTcAv1LMirH8zlLy75EaI7hdGP8ymYAtxZ1lxPNPUGpR
q9zrVZuHIAFkR/qwV4dcYay8uyr5c2cVEjqjC9tmmI4TdQf2INqGJQn7UntLeo03
h0575w88cfAFsVrzd0EA5jx/e4q6BY2I2P3KjmF7k1jIWo5P43z479xHHqp+gd99
IP04BmqbNrbDRLcJQhUAY9vcQ6jKUd925nW+qAQEQ6lI7kOZLjeR6Z/fwL8jxs3y
5IUk2H+ocL3OZuppvv7q07WikrsogbCaF+w7FEeOpCGvW7ikHk3T7X8HM2tUjlTJ
TFGdiIdBmdboC4kEfmuBoNY8td5bPTWeR38vQzjjkkY8Wu2xMAV4qSqMjWIBhcJn
z+2tzTcIS/BknXg93xXbnP7zFOBgy33RCyE4EybOB4o1biFqAWPbRRDYnlqwJqn1
HDVCpU6nTFefgPleItgJQCg4F1upC0mMc0dGLUwSK86ffxu0eTRWWXy/lesS68WC
wYXWoamOlv0LYLCQEWVUNFdV0v+FGqenAI62vseDdXTjo8LTrMc1gxyy0UN7VD6o
b9aTEB2UU2vDc41DhLxOQwRrOFi5IdziG8VJcakgzgi5FV7Idnjsa0nC1tPjJVhj
UNZpiTxX4r2Lpfdx0F3J/H3KfMMUD+yUtfBfb8K0x6RZSd7TMx5FgZPufAu+wEsE
XzuQELizdivf7oBZz6voHhqgEEkjdvcdxh5OJWN2ZfoMI/ljZ4PDUfnlIr3lTV3v
7VRmZD3gAv6UH8RzbEV9k9/fY99mCAx4VBOAT6DtCOeMbRh1qREMakR4YyPWeIQ2
kzdKjMETxpt9zFDYlFHqftHmr8x+q6oH4F+sp+/IhRXfqMSxvk4RVVpbMMEN0Ant
yTL6M93zVT8n9S67OSzotFcVL2q/zvMWUuXkqzG0kpbKPfyl6nVhQkdME5mlThq6
n+k+NbLVbbQsjdtggQuaSRwT0oCiE6pi1ZgDLpgMWbviL02uXvIXpJAlpOMy34T5
t/AyxhoHJ0+GZVayknZXvlDtdAjQQ1Q8XwnamOGrl0OmXoiHBZAaKoIZQhtnYhqj
Uk5qI4HM+LoyOwEbvdaSlwnykHALvU5jzrkNB9QutjHJWkAtBTt1oTVxJmJ5TmNB
jkSAl8VQf/T4ngQX3byd5tYXgGOJHqw+ZvJ9HA6G6S7n5Vtw7j74lFu8S0KT4xEA
Qt9ySwIipFYt2oPSeOwCkfKBv1ycTwa2ZjiLUkC6Le2o039AEDYFYFWCEq4mvyfm
nNMDc+/wHhe9IEpYS/3Bk3/KiyeOymLOSAQfUPXXD/IgWqx15kSJmNLyrH1qC6ig
4V3pC8/rNhjqw4nroXz3q1PKHVQFY7nhNrTwc8+kKKucdvn8FCSRv+nCNI/ZmXy9
6VBMPymIYOK6xDpRBHP6X/5JnK4vavBz01AU/EnNcU8LMv6VQWtNpb1UUVglgmIQ
/Wu6kjDzw0rrpqCd2V7b7QslS3kDuZKV+TpHv5AB6Su9mJV0Hv2/aKhMIsIW8MCR
1rPYYC6G/Uf4P2JqGa3y28M3hF2m5BQoPEYZggYuqjXqm+nOqMhTlXJhx5VJybpM
WKiGt+mbD/MWjODm6u3I568S1Y1sOPD4y2p45DNoYkdAcyQgPHbeF7b9WpoAf5LV
sJrLs6EhN2aKvDOynO26RtFKtV4Y5xYQn0q+cTubuZG6es6Up2/mIoB3mibqZDF0
5FEg40g4WPRi9KvDFz+40R1G6d1d9AgvQSVlwbW69aGmOqoqJAw2gjBaha3WD/L2
OIZuWGuVgr1o/9lkUkawSIjybEypyPaJjbtavMqasCSq/lhOExflJScJQ+ZocZtm
p2PJ7BpJTxNap0mymoPjk7QtBnlCtOyMSyKyLmHZC/A8oVD9v+JPW8uRxYqSB2WJ
NeJvhKy11PiklbLtmjFJ24r3dSma5AoKpZJ38/kvVnNU07QBiy4OUdcrqranJ9xT
2avXWWdzbGMifHzKBVp2EGSL52vlxB/trE++Tf579UP1WXiOmzUL8pd3G2x+Xou5
Jh26uBWAFLiwew8N0ESjVT90zbS+GPScYb0kGHRDyU2BIJwmALFPwTnWYg365MG1
WwSSmG1OHkDzmqwmhXEdqYpW3Fytsca79QFPWRE8uRY0X7yNW/xU/Y/K0NeENRlW
zsJohjvGqo5jHE/Q+GYKwAW+Mttio842PLaKa6O6Ib7CDlo72rft7LMZsS1PvSLQ
ov4Tt3ArkR4JnXBe6fJ/GQnoVzTiaAmCFu+9ZobiHPsl1wHvzwb/WigjyYLUERd3
uanGk0OpO4IC2Mxg/DqhH0ovrsyhLDBtPDiuXg47bp4GjenY6kqxJwb85oy/Vsmg
QlHZTB5Hn+tH11M+eNt6D9xUbYAeYVZTzMq/VwfKrDffYCh00TiMkpFfRXlIdGwQ
Ggl98UWhgqbDTIO8k8R7JUUXy6ihohYyJYknK9fKRZqXZzkDtAnMkgvyjuE5KrUK
x1/6WiMOG7BOQWMN+XtEQYaUJ3EL781c/bMKPOT2B5kctimTKq1e6eHhTTrgHt9g
8QhJ+Cy/BFt3BMRUHBV37Gp9S2cMeKN8sfKASN7++F0qryUEc4Eg08Xcxr4obcGC
sqgx6ydH0OUZk2XOX/FZ9IlixaMIFyX4rSXY3rvM35gxkBht+Hn2/VN/Gv/cGkra
J9SOxgN31h8jZFEiG42htBSpmHAWbQfMPWbdJsLxg11ZInryAV31EyhRT7oFDr/k
QaAC1hTXlUXqd3sRpBvHjylw7NnrWOjnbjEYsm6b8/Z5eFGrdNKrrmg9Y/4/sw4o
89qoQNqPq5h+QaMY+am8jW7Hg/yBq6Sq5niJMk5p/yytBVQvrmnxvrKbt7IGhlu0
cOWxoKmB0TIxno6V6T6vKKGvpEIbaQC8VvP/RLdx8XTsYlZC2OC4Kqo5+VB4UAlu
9dm6lUCmdnwsoYwYYXeuSZAknT7HZ/Hg93qP1CFHQLunNXXrZE/XmI+rIx6RkQCc
b1/lJyHvdmlXOmkwHNieklpUTKapX29OSWUcWXQsw81t4huhSLsNO3bwx9OjMwBw
ZysqLMeMdWlD83btocr9va4aEgkOYIF9IlIPfJCMm0sYViTmwtgctRQNmohaNhbd
A8Tj039+/Rb7/Ily4HXJqEAAUHjdFC5IzTYzQ3DbXJEdNtjhaPCdUibp6AR336gT
NCI1Hk1rG0PNUcQ6+ueHRwKws9imHpu2PeQk13kzubxzkJ+IfukjOWmAxF7yI/j3
xE7dVU/UHKsfLl32iSiUoUjksx7h6WR+1qguTOuDnKlC3hFEgXoxtsS8tEVeprQw
w2lOfQ1hIYnDj1fh5iCpnZAJs5pT5mvNKTIyGKYWK9oSkmyUGaSBJCXmZQQpSGoH
M6HcghTAg/4oK2+8L4b4jEmn5J8Bqx/KYB5uEIk06KjExp1RYp/aGiIwLrzIxMC2
Rxi8XnDKHgTVitJYapogBG2cqC93/XllOcseNhaaaBdWPqNXxlObSu0vdyXdevKT
1GCYccz2f6Obb7zIepkafQzgG4jjgBvCb6aRDljhH9hxFPNKvB7phMHRfFhI6RYs
EEWbXnzRiyPtZFpG8eGtgxm9wIwhfJ9k+zIGJ9ErAho9DPuNFSGvZR9iOAdDNbAE
m1sL/PUDmmo89xERc3XbVORW2Zkcb6y7oj5ywxUua9aYER9WATSNbAWwxhdden5t
eEuuuJvehYU8M0r0cKccoxXkdJLWHea7otN1UmpCHzyjY6ybtqk3LdmV8+oWl9pr
bQc8GVNXTPyNy9MtYREXafnetS1GrFmtUbuPFvcDymJbd3E8RR++7byEUFIhcOgT
legcFslnZKrVxx/oNQgO7+MJAN9nqR4Uw/y0exBUjsBzb5PA2zYUDWbfTmMlwQ2f
RJNO6M7uU0KTL82WvsVaYB0jrlwN0ZCJZA9+109rMel5jOuSZFrrZoApB0g6LpJx
c6U5N4cLSUJRO8BNbruLKmGUS0wRdrXpJlsoCkXeQDhgXAJpPfMvntNVKNrmY7sQ
OSOt7ifqYSQtAJpalRqG6kFhytgB3JoR814bZD2nfsSLQHkrM4Ev+sUbMq7OkDWo
66irvWXfvvP9RtPcYfNLAz31i6ynGWzXhsaJj+2fkM/VxUYOBn6IB6tUsxBaPb/r
mq1GTr9mNhDc+S2mHqKmyyuPaI0MkuX2aIJv7/t2VcwqYrL40GUD9mXK2xPU5eJK
tK4EwbrLkIRVwZ0iO7J5zSWVOIHL9JIwGPI4RJzbCrqVbEJ4WJEC9HO16lW6H8CY
sYH2WkOqYdbKK5LJaIC5S71ooISxw6ct7Hs34tm37KgWm+ZTiYXIMU8OS6g0Mtog
BSuFNxOc8UJLGephb2LoNw0iUtFaI/r2arWIc+uys6611gAkiOahTVDB1/mrA0c9
Uiv7kLUCV9fi8OIU2g1YOotUxIuyIzKY46i7Fn1GMyOMvA0KhNRr6VhFTysb46hZ
uqYeV8vmYAGS6QcSsQcOgnpSXyz1ozyg0g9FIBNYE9UuhkpB45ERNEGtzSssfHnn
Yk8zS+dKYoVc8UgmJouj+sE68whq0QUH4BkPk4F6vkHRlT8cR0e6Bxs+JxS2JLww
u1IXYGs3/J+0uQhEtzveuV9Szp79BZ/xlR8UcvSoFyHApL4AKTfY1z1jLr9N2/DH
A7IqE+X/LX6AHZv/saSHe3DTUiEg0Kzh81pWk5tBNJZ4+EdJKNK91zcgxzw3kBGP
0mxU36oYrquNyQwc6HLvWcnYWoXv+t0o/gCJ09DDH9nR7NbRY1gVpQm955ZrPiqU
9T4I8lwQ/ODXXEvoritGYTJkC1CyGNTpezdPNZKlSr1azCBjSlGUDnd+tKZ1RueF
+YHkvgKsVyJCGkFVdrFAqiEwvaV2zkFBM7PB6m1KnrAQeSFKPBnzkA4m7UlSWftj
RjOqTKYeO/ZMqUI81scUL/pXMmv/8vfYI4X2Rqfrx3Y1Z/5aZUf09eZxnYiG3TMt
yiT8Rjo62GKruNOPDUgkfHX0y+0z2BHK6Rqi7k/ziZgRawtbkFqn2nJ8OfRH9qFL
H2d4km4b1FNsK4arP4u7C0K3lPicW4NQonDkzLk1d0LInvQg3Cy9Xto9VYm45rxM
AoBZsobIxhgAFRIUAJFNV8ozoFY/pitQCcEZoRjoBRSW/AXyaZmxJfEOitVXLHsK
T9N1xD9lnpu5KgUe7e7SIitvNfJODSnYmr2rodMDYkD3h/lllakfrAzYFgIOKzaQ
XoG6/BZg7qx4KFwZmf47INFgAaNX+brnL9raQhjAixQf3W3PW8xIzoERAsGMTViq
4HHXPvuOjXLkW00iM6q4oddZ7SChOJWLOCPMOozg+mxcCcfClxYNL+qI8co26sFe
4M05WZkmXRAeT2SFZS1B9COamAYCjBTEcwYH4LiEZ/pgkRFUvqg2DgxAT2ome0K5
wkgfMNDmOA+26dqam7WXrhA25GyE0k3VQRH97bRBSg51gKT0AgejWCyxjX0NWmXQ
Eb4qbUA12J4Qd+ATAiQ20chcpudUe0TNm+/4jRgBhDs1Jb6xkzA8na5KdwkKUpMB
3u/f1pnnqWF3XpRq75buzuNW2G7m76HrgWQJFvUrapphw47RewhwOQ+zwmU4WfuX
iNbrD3luTQGAyc7A3gtW05+1FVczgErEE0heojDtySog0WRRGVQj1OoxkTmArQdG
OCRyfkDrL0WQektCoYjy9Jk6zqJLOE5QCbz0pw4Ur3pUCmSeHlsVdAyLEcvCp4pL
69w/VB72T7dWObpBp/acuwiXoM07wHtbhH7xjY0PnsLtycDiS2t06cVvc1G4xOE9
1HuMbJj1rDSRgXsoks6Ecmic2UUpgpG3txYADPfP86lxP5lf651DBts/OJgRTZMW
JIHuA72m1Y2UaUiruHLuJSyqK31VFpknM9nc9tMD7WQ3mjWPjL9ht1V2+wytn77d
3Lm3dn3SDGJ0aF4AAPUaoMzstZ89BZN114gw8NXBdVxlUbSjpqJA7LlBy/RlZhnB
0gPA65HwWTGBDpAouD1GZ27x5lu0XXyxhydtEc70MZ+dkAUPS+TdLDThYllkZqz9
j9g7a1EaoDlYwKQDIvfk6oTsG7ZEIxyQdB7birm+/yNZW8Q82QQkbbRh3VX3iJWQ
fAZ5CHFvMpemT3tILT419PAQwy0+UT41k5rFqY0MYwzEYf+9JPuh4jsG+AHv5lbq
+yKG1qSZIVk0BNGlE1FVonKRP+3jqm2KvNpgyXv1OIxcHL/NRb17XVM9jcRopW3R
L/GM0e7RFkKiW7MNwezof0vBSiw475BnGfKmBjrs0iBu5dMhrXstdo0KWUhvo2vT
CiS1g8ibOJ/kkGwiFMqNH7ThyXt+XWRfEKQqlJVKRIgwM7fm8a0dFVvkn60Guckj
HyGTrBU0oEMo33sxaiSmT/au1CajzOQY2/T8QR9AKizipIjMSKRtO1XV1skHF9Zr
NS38QQNa8B/O5zrBh5ZBxmk+PiwrrJv1iyQz/SziiJp6kQt+8zXt2qJ1APnpm/7Y
I+DTECDbL+gDEsq5eaNm1CUCuCnkGP5j65XwwZ2Qgclcis6qZFwhjT24lviA4bTU
YFEai9cPTptlP11Nvlj5QQmeF4TUgtv5kzBZJM4Eh4ZCQcAFJQdxhRGc8VhXX3EG
jcWHyXDnKRzzXWVrOfCIneMrK3LpfWhCKHRiPPFi0FbDB51SNtMwslYKtgeKep6U
e3WklrA+ocErBvj5f0D3ipcNgK2CsmyhVaM540D/ViqX6J9pmkPs4UOmjqpMi9WF
blCnEwR6/R+UKimIhnNPNEospcEknqdobOyfVN2nj5GOcdZjQo+uxqJYZgxkHsU4
s9N8xq/CuzeVIZ3Gkpjmk7X6d7eN2mx0LWCjAVPWmwur9TlNW9zQ1c/CWioRhAqF
fOiI4HSXzAa8xulRusAf+XsLJTvd7ew0xzR1Jyyf5HiVIKtkh/Af/L00cHNJh62z
EPKMQ+FxedeMUji43pmDD7QCZUrS18jVc1YVZ6xwOdLYf3sF6KtB4aHnJRr4cjIT
FAEoH+NDTrblE7hyzllvW54DLMHO6l7aAb6RH/BRmZ/xiSQooexjCbU8jC7Is7Ci
Y7uzrt5qF1MI9tKzE2sHkD/Z6SrWy4iX6+EcArRnBZJkdtEJLTnrKE3OAJaxa6v2
AxT9pqpJpmb/1IiaYqX0UMAU5kh6es7nDpv330I1U22NIw72Se7l+daZ7AtTk/NO
W66i2YRWvLnIXMcv3+alNsOgN9ubYyV/1mMMQ2wgYsf4I52hMvmetSmthnRWVAYh
HCJ0VIegP/YcpmgnIli7CKN9Bw49cZFvwj9y1vpMnwaiasKkBESZYZXV7qGqvVfY
aIwmOaQuq+5CJGa6YR7YuFB9C/5T6iW7lja37GwSbTYhrn+8wW25CTQqJRZF2ngj
7kEkVb2t7SuO14K+oXW28lUB3kWXHvKKQ/8201otr9Dm+AMwvSspTS/AhFzSHeHm
UVeqnED7g/xEeAC+ZLN93OSkXs7osHE3rYu3NyrKAZsM9vfThxojBtJP2p4eMDJb
OcVcc6B04+NATXBwsj7PC0I1SzS3aNaIUQxlEtZKN6CJDF3a29UFg9ft3xUOoA/1
xHiLdrQ7jINmwNAQ0sSvrBsL8gyNcojdZvdNxF70A+sYZZbqCIT4qiyhuEVucS2R
uhrloBOdAc1/vf9QgV6tbwqfD0FKT/h5iN82gJaM8193W+XYpsxYH7YH6Rp08cgT
3loO+EKg9tn4Y3+cb7AOZEXmd0AYpqpnabCrizDJe8zIP+IVkfo9Hp5MsoLSY59x
+Kz+yhUDu7ZOvqBM5p1wET+j/7w2JnCT7TiMBNVJpxQmr+V7TWUzPsdqz9jgg/Hn
5oRrprhrpCF7zc6ktJcpWjwpamaMBKprk+XUwUlI2oM58UvIA/HRpm08ux94U/hH
HyJ2O/S1xyDesItTPWTkti8uLFy6wBviRUkN0bmYqTDcgq6zrhhjAzI9BRBiiIsc
14lHIMy7emx/Ec+QzX6wj0461JBNT3+bLE3hu/sHv73V8aECMfxPHVz9HofUfhrx
b7vFvwV89ZweDYWb4QVCffsi7+o/N6iYNSK7EVcaTreZHHPBILh6tyYYtvVeK7XX
/hlrEgq9ZXaElNGaAoo7yqbLM+KGAm409dshlGEhNkm66M2DHNbMxYem35mHLi7K
DEyzUHcOZhFUQNtCpfl1EqySDfrOruwtZ0W99QfIOglMBDMMn0ur1wCzTY4HIaBZ
/Cbg9sqdJGwuPetdHHqtoRGbSrTHWQ3/ejKiYjRzR8l971o/rGUjWGEPdp05aR8f
j8iodDu+oFBbmiUzRQ9328GHRlAfkFB3nNxdiH4FkXpRqemy1Rm4yWLEUw3AX0gQ
WbqsM7m33mkdUTAHoTN90VbfwCfU76zT3SJreXyOlm0XgyCw0edfryAatUWnlMbM
6/OvwUA0b2VC70kYTKgaBr9uIdt0s2M1rYRKf3/BvwHGIGCnl+03pUD1v0HGNP3I
3c2G2GLXrWhtGnPTO6B09dVu9BdK3K2P1Yemvtpq9e/LSCFz8IQ4TcUE0+oIQ7wS
Md6BMd7sdHShORF+DH06VAENQimtPqI+64Y2HWaiFwvBbQz5svFq3f81ZpqdoHVN
kMeBBLSL4IhXLdMu0gLDsDexPa54ozo60ZhmzC/kuxWK9Bee2nz4QXKuf0hTmsao
6LNEZfmpOdwPhyLuex+NRfyHqECTG/InlsZTvAruUBSxZjX9p3eZxIIcqhlXJM/X
xdLI/0c7UDrGktda6+j2P7pJz7Cdkt8x+v4nq4Ql9Uba2ooeQCUEp1uhfb5Lj8KM
W6Qr45uLhkRsrpecRJ03dDV86bhzKIH4Sw1JXKcJuWwEeSjFa5AbasYeZdJTUVrJ
Njo5PYUdt7t1qXYRl/q+RnLOGpNaJjdCvncrRlJg+vB8kqvWYx3IbKChQwPBHlxN
VOER34XdXPvbSzv7POQN54RtOjPTJbWG/np2+zACRPHAe4CJHBrxHysV5uo50r/9
2T/ImB1ot2Q8Vn4hRdT3GLZmsBjJRHC3S6uAnldUeNxwo30noSl2CYWwhURVgdog
CdkE+yTd0jyTdT1D8g8KAMYW3Yq44tzgNQJXi+HwVyB6BJYmlVc4W7mEwOHt73Pv
sOL8OqwGccdzmsChrVKhW0IJyaTK4LZ6E9wgv/PVAWFkxgbp51eNe1bw5UBI2f+z
xgp7KJWBLpcw0sXJN33BwaC3VycD4aHXr8HxZuLojcCe5IPKb39MxeWZC6Qvo1wb
+zvql8rdzqP6ux0k3Wd30kryP+EmyFVe1jllvHVDWO0EO/TiOq5zd4b+WWn16j8h
dR7NMgQADaajJbaF+a/o3pZXVtfvnr/BcBAGhIytjr3WSQKNC3PmnvXxCDEkpjZn
5W0Gm9ZR/GR6ogE5l8dvFzO81Gbf8fHnQOP8EHKBtcVxa+xPq+eSONXIs1DYEPxw
gFaVCrhhs5WkMjH1itaeVxmDAemvjkWCoU9IcUZ5bSmrPzpGDXXElA9uZZMsUuMb
3gcu6oOzNbeXvl1zaMZ39AQRgKrqd0+xOfmwmJr6ERQ7iKOVHKqlYyvYA6PSIYq+
UQSdBCnDl1Dsx6Y6rBZR6W8LMozg3wv4ywVHmumTn9qP+IyV+TD9N03QaCC0ez0Y
X0XioDlP27+TQnKbmD3VT5XkzhqHWSa+8ecBR7NU/FcY7BXzlt9D1N9VBAUE74kk
oB+V6tOIQLyZMB6DF6JpdEI+7qdcs+wdVwLJE/ge6h3mp7u/ZgyFuxUEftO/fwXZ
QRcvIXDnLt9qK7D4PZFq43KbD4D45LxtZsjtv6TBQy45/1VpwQYts0c9RIXb9Gav
dyDoMZFTxYG8+UfJ4fgv3HJgJmq7UHIW0K5h/bekMv0Wv84rpMoG+Y6ETclexPLV
+iFzYqjuRgnhH9UOtV7gsF9YDgznMKUzlLmQ525f1nG4gxOFPQ7Is6JBPB88tlxM
/PYAWlVu1/j2dE170AEHFouQBi3QDzD8CHxnEF/QM4/ENFdKMohi3Fxb/3M6SQg+
qyCq5EsiSfLYhPL4onHS7QS8nqXVP7ZMVikhi63zMr8M1+YGLeC+YErRyVqWX+3R
2yMECryISAwDvb1HjhYeq/sS1IcHHvyEemR6rS3cwGyrerW9EiYoLCHsm2XgxM5+
lq8kGZo7xmNNDJa668xF2RACuBDhmtdQ6KfWgtqpWXeexCuKbRr1tmKlKlmHCzQ6
SSrkNSIAFMxujfk6dkr95zgTJv1yZITCw3x0SW+W3ZX4vb+Zz5NcS3kzieNLXkTT
YiQ1lJN0UZVgUOkAMa9ZYlcWD/i7rA+AMWBjg+i9nN5F8dWa936q6Z3AwbjNgB5j
5JAEHydT636qpzX3uMLZ3B+sh0fTgVdVX7fgDhPlIbvx3Ka1qjmMs+6dyg1byDLh
oWOEaipuw039qK5Loesa/t+L+M8old0nxRJ/q52OaEn8JBGYBmAiPEA4uBcSdqXJ
nxW5YBymrj3KMtIhAx/cxLD91R3z4dp1C4BRWsEnHeo959VMiC4FUxqhrl8bPkAG
8qtxtVigOjtsLkCFBZewbwoEJXGwiBZ8hfIumm74URPoudgAgQq5MPZmXlWwtXu6
Tr925IY0NCmNdYnxT5KYUh6ZRDzHxcpBi8uBKmiAXJeqs1BwevUYba8cU5ezukD8
qN5J0InFb9WelsUUUw/BCmrZ0HgQWlRg5liPZhTRdHJR7r4kDhRTL9tliqL5LKn+
eo2MNqrp03oN9aS+3m7iIfWWDFVdsnqBWXPX8xVUrHuUU7CTmnVn9QEB2Z+QL8SH
EO0+3yd97YWKxiah1Pv2THbPm1e4U6NLQce9h28kdY8fYPCgAsTm7dsKpm/6sB1n
P/EaYdygPRMijtqTmEf1gGdmfobY3uCLF5HllfslLZ85GfmOABOGbLNZWipST4M3
i1jVSwIDoQ9GNhHMp9P7sfHmEsJiHLry1wFUVCA0ry0zR04uX4Bkc+r9PRgvvBiJ
YFuXNYZpdEb6KTqm8ShyPlC2xZNbuxucIxGZH38nn9dbzWnupXKtEmk3yVlJ75lT
oFK4vRJVxya0Gyrsx0voY1WbzZ4MzcrGcFEPjkvRNO9VxHiMJes8yZ26mekxyGHT
I4UjHnrK3KHu3Fjowxys0Wa75OH63CoDC8/5oixVFqSYxcVnvycG++myLu2T8QsA
nAR/kBTKP0WWWyzHNJvew7tks9o9KyE1SA/2EK3uIU3PUMGZyfWv08Zr9XXOUBZZ
f+W7zsrZVE1yPpJnVek5qppKcT2yX6xkwyoZowM8WQBNaxzdiUqSMeDqLlhY8626
SCseA351trbwibuNzrB2xTu5A59UBgM9Ea1atRRXjzSODpWD9WOOeKadSYJOWfza
/8Phqd3NqzP6EXzJdYhFcv6EE2oc/r3oDZfYTczr40AxdSFdQte2i4yXxP/9Rd1W
N4TjmAWpigo8ihc8XBewL52oBq/qMsxJtLwECFKNQFvZQyHKlOYKNCIFr0lgFz8k
GSfhZzERRDIOzh5cytcMuipMXaeQugijyAx0OZrVo7pGR4L1UmKY4rn3Xu+eKfMo
VAM3j+qL12hN8HblxIptQLkmoftrcx1HwKFBniWyIRoo2K7OiIX3ByGQPbZzOyVL
zwZ9/Zf4D9vKRUFbkFeag5sRU4WhmnLsvWuiyI00X+lBCIej7bTneHLWnDnVXB5Y
LVnepZ1DMaD8X7H/c7gILuaplEyVkOKxSvoqD+hpN2xpuhwKZF7KfzqzPoS/A3Dg
oPsYW5CNmLjekql7ID9mmO/4l1d4JLeGGL1Ofex3sGDuS6IFLiGRszr+khq9oddJ
2KzPPimtpK6xZ34mp4RJdEiZ7V2B1NBWPP9PkoInLXeKM+S1D16eCgWCOHN1onbO
Zizn77xKBUwBzvB/6B75h4W6PF2kd1VxF5/ALzZy/+PMdLTtho0SMngLcdjCC2AU
/cuad3j/3Jk49BM7CBU++6Ni1otksL9rVWoAxW60gsCvT0+P7NsKCUO0YX7iS5FF
vVMeTjWdxWo/S65qj0DzO8cEDzTi073+MIPkDtnBiEBtvwPlRsNLGZASjMMV51SK
yrK44rBumPjw1YbaANoWNfPaz8FyoLSqWPJ5XDGStgH7653zPCScdUUM5cCcwWRP
CQMNfjJsbVAs2jR5WO3lA1GDTWIzvqihA38jso78niCt1KqLCedKI3VKPrKTvqV3
+SrfzmpKhV2MNvqq4eXH/rM0H3jkXPkzUOn6k9BcljO+bsluHXkNWv2yi61bgn3x
1GgGmAh3bXETq2XiSj9gtyeCgGmZaWv/yoOD9pSLk7qmejaK8FgKQYF27Q4c9uMM
u/4U00nWqrR708aqZUZ/7CJm/Gd2+idMmmMmzpFUJShzn5f10bOIxcV2Eg7YMY9O
rtvefTDT5j1nH4Sf981vsteRWWBH83gz1HTp1dJR6cUrMUjwYyQIpIl1xo1ifYBT
IASJlQjjBKkhiQrr7zGlDZXryExJFDnW2WV5p6Yd/7GwG7jeT/ogwYYz+uRPUh6Y
x0JG3/A1K/ERNtiObeWqvWmZIde1ILeUvun/tm2ddhsN+neTWw7q+HvmBABbVvou
H6rb9AJ4adWrAJHWY0tVKp3oFgAC51yqRHUBHhI1cABxDVqxvzGnnhtVuuYPcZwD
lA+jU8vtmqkkTQ8wwnCzO+rszJ7tjoyRuO++5uX5QnswhcfuXmDF4c/KCbe3GHkh
T0jr2HakBd4WpYicbmNVsb52mt4Q9GUBrNIwdppZjIVUYkTPYmtGzCBDf+jar8t0
fuu8PxQIow7YdJ3PuzpSl2ohp2g8M03iUsuuWR5i4IpPzFCikK2RS33w99e5DeNy
dqVjBSMRbIHfO62fu2VAl5vIokTkafCP5mUKS6VxR2eJy9E5ms4QOlaq5uD1TC8f
zrJ15YuMQ6c3QFBz/a8FTlUpxcdQx4ctok2sW+cLV82rUtsRR4KcPZE4szB/jmy5
gZBr7lp6qlZTvqu/+TrNBoZaJdPgeWw+l43+qJX6MZuNRPHuLkGT4Ne3X1UfbQGt
NyCSMoFHwXjzj8Sw2XDs2XTH5F1z/XQ+lacS3/tpHWzDCulhX0oVxcq4KZYTvpoR
W3DhA+QdZkEkLItiiWZpsaVhAXjkRXgM5IpHJlICZXXTny6NtoBr/MU+Ni+6IVa5
mFVOlmlOhRUzqYSzOpZsGpDZ4eSjX8CAEH052+A4C003LKeaK+4dYXoCa1uzQ2EX
5yaNTvFFow2EGQAVWL57eNThreSS8GP6jn5AROsI8/35puSdKccm05ufh1iIPrtw
+ILU4A4aOXtWmvW7h7HBU8sxnDfXo1YNi/ck/5t3lzMi7Pv8Kx5uCtfPlVABc/Gk
EvfOfKYmL6w++zA2adFwvCiqma+vkqudak4k10djF3sh/DHRuOYvSTQbyrx7zxsa
ISpbEwdYscTm1MIKPgnI7HQbkJfdZ3gjBx0p//y9ghL6mnwNIHlKBdei6qCLjSza
vdJkkjh7eX8locAhzD1hRIRCGElcmSh58BpxwVg4i2gLKofmmjwfGqOpfuZo97+G
Jeq98yDYDcWqjRikYkHkX+m53/Wt44LOSu1cl08tIL/AqaoCpw0vjlTrSOuL998/
QuNmfU8rntYlQnjCL1kAb4NHNUgnFg9rGKUggVKK8h1jp6zGiPuqkyAUUAdyGypK
dcb3KlfrvVnNPjrU7k+BgsnINBlUGLUn7trgveR6d9zftuAZd/th2AkOKbQPSFob
Q+KccQociNLMalaxkIz8CaT3zjQ4tHsRsV9pUZoHm4nffZqi1aHjWxT0sIiDI2Wu
BOUPkFEWJJ8hMPGDn3PqmBF7xmNyCP3C+kFPE2ZQvS+vNJSdBr51rVxo79GxQ3qn
fEVmLX7l2ud9fW2/ggMupdqqVE3RS3NGX9hKhfacqU/qjU4tNAmj0lLwqIEUuikr
Y88YCniR9TXYRef8q+sU3Po9mVqrOwlJBcbSrtPX9cbbFuib8r2f3GpuwqsqZ6vJ
naC26i9rQSaaY4ynZYSYnDzl5A5fbPjtPsjxlA4bAce0tEV85Tt+Rgh7EzBOiZua
BCzEMVPdiJBf45dlaCvgOIzL8RZcIt4XFDH5pDwwXBpufR1VWYU0XL+iRDs1HqSZ
I3FdTJNeT6IDWZ+2N41CXwn5lDEGHO5V+bBujhf+Su9i1V+VaTcw1uYGvFT05SJD
pMyyOjXeRtXv+DlljzX14mYOrWMgpX4MYiY+IdFehXldqeVIykURoMe9z7JcLrdW
sX2mf4dGnvUo9SmS0cfudQtH7Ov2+qyNeIjJLe4co9X/AIwxwit6N524ZjN+Wy2y
9xemN/JtW8yvhaTrNNyzkm12fMJcNqXEfK9HSR3qIHtHVLPYfGMHCM+HrE9bIPRZ
+dA7g/WPGC3T6VcVDatNuHCRESeHiwjCwaG9ixeYH7YmywlVtSbaILveLhE1Jsod
B7uJBxCv7Avn3VBJt5phgiVFV9EI+NK/eMR3SXF1+/Z/FqvdJ1ywyikDQm0CW0vt
LfeY30/IJbbj8YnbkA6aL3RoqDjPP9nObwoPN70zn71CvpWD1gwSbKNPAtEPtfCD
zrJFpBYMMLeDUkAsAWc/7DqgLS+ZZbeBcea2Kunnlq38XYfb1ospXqAjs831BFwy
Qx97OvdrL8L+0zqsKQeZ7mL9y+2lq3Yf9sJP4grnANYsWfFTD1OP/5r/DAPyW9WL
xSMGd1MTwqkdi1GLzTjNPJ5qgzQ5VDKv2xfNCY3xpkQWcAvUr9xjy8Evs3MaMM1s
d0wezcKx1u3xDiT7gbY9l5TdkyVlZTUhmfmyuyVEgbXZ5QgogHl96b472ibhMJRG
jF1WR0OeTrZ12Co2attbPl/hF+ghC7gyL+v7jRf+iP5/3LOR3S2vsD2/XK6WxWLP
jF0tljGFGS4wkSe3V6uZ5vknUCT8UMUD5hbU37wZt3OBcsk4N7vvIm7HW4tYQjs9
FhAN2sthke2L3oNqZXUinrA3C2CZF5kmzkYVDWsM7oXn4I85EKby9pMe+j1Joh5E
3IOMsiElnG+zMzzr7pDu7DFrbkISJjN9k7FZIZLUrX2Ha5fH7XeaN+rUVhLBnN57
vZNHDmtBKwwgYyN4SkxURz7iVHdaTNGkxLWWzX8TZnVW5gv9axbNtm9HeB5m4cy+
z5TXOaznGDAOonGf1QDFx9A+ifkMfj6OpR/82D27pjAkQiyVjGlGezJpnBfQ4gZK
x1heDzVvUfOeVGc+jmYd9UWSJaJELP8PbVSsJEBCUVG55qc/snhCGepQB6auQ5vG
00fWDILHo/8VvjpLZ9QBNzH+MBR66VGfylco1iEUV/87yc2QHFtc9O6AIk4g7HW+
uS7v1V+6TZSAsigqlr5KsYCscUoNjxuMND1du17TMoJ1uTH869YR0CD+7juAhtKw
47I1JiKrMaKOxVFzFkA+9Np5VwrsotycANDnT8mXHQAiEcOzynfch1e7YK07TN7W
zgpyn0i9SxxotX1h18K9y9Dmg0Ii/OtFEjiscUaw/YtGiORQjHFbnOc4ux+TacTd
cmh7tmPgYOdeoZ1swN5pXCkNvgtylgTpbOmzOG8lTJyTSJP6OAK1+hcBJ1D89EEs
dd9PgJENch/zEjHkR3l+1Y1x3v/eohSiRl3GVp4gMCoHXelqQ1MVkWcn0cOh9fvd
/lysEHdmczLVeIhd40f1iNiLIi4YPk2Bkb8kqfEpslq+kaO6o0m7QfeZO7oPso8j
iF2AxaGhHW7I72CA3f0ykYG3QGBAmu03PyiXX62roaffyqoMy55ODa3YqGzs+cpF
hiFl8GyfxYfLYdGjVWh2nq3l2peXh2xzZNJomZ1Vag1sxm4C/uQIdKVqqhEABpO/
ewD+83hiSc4eTt/xGWqpazZLdCKsE/LQ7NFuhzPPvsZYtyBSQww4HhSLpq4Hc+JH
7uVF/NQwSpLw+XNOGGPFEc1onz+WuEMGzE/5hDVoyFUH/zJhXD5lcDxpJ75S+v6k
54CX+uhr1mmyvluM66xhKHdBu+sH1vL/1riMUGJnge0fY9jKA/RNA/BShvcUp47p
QZ4TpjdJnf+WDa6nNxeSHEbcvpbzi1wauPpcSEeKXz2ZfC/n9sBuHbVBWsSxREJM
an58qw9ab+YnEUMU73L4uwAzusj2ES3GvxyYEP+JIMMWn0KMZRzkZJ9+3FkdlXpg
dDi0t3gLy+Xw/eb7hKGcSM2BbrjbO25Z84aovEA69lzPmGh5pSWBAePCx/LwDbdA
/vldHJT9L4UufdvCpGhZaINQAvEMNsfbhtgx9xnxroHnmiiQEffNx1W1CLlB85Zq
l6rq6CNNGnnz+InWb0TNNh3xFxux3G71FCjx495O4egIdBThbEv2YCalL5Fegrp+
nPiiwSZC9FVnB2Ses6jymFJGrpL70+H4M3+qtagpbhgF2zxmmS6+cJKyslG3rIdv
pYphejrAl47no6ZPIJdp283NVI4cLB2OE/RQVNgdTbXe8U/MtGB/iyjLX8U4k7OA
sPgv5MygMqLMF25gqEcJaLggR7LTvXGcUF43Zafmbrn334uNev/yGBUMQ4GyxZXq
G02+Ds+nmkziwhQ6iID3SsVcmtnaERT0jFewmWegzh1/gGBefFZvdoIpD0lazeor
Fdf8Kz8pCQeHFeKKfpmXIku2SnSTuc0lnwYxdr1NxidiBg5TkLDFhVi0bF3v09Z1
fcm32GTsq3+73KbHT1GN2Wbi7DKXHggYBxG4n5J7KE5bRJQ8No/9rVJj6Jc+hy31
LBBGg+OBWtZXBy7YlNWq/9znFJsyIJYRHAAMwSgkOPqFx0GeIukx8aNJ2vQcgl4+
cXo8v5QPLlaJTEdYCalFAe5hnwU2OKX3fFkO9/0NZ3w6Fa2ZLftUFjQrM42cRftR
EHk+tRGRIVz4yGOAo82OCZetYzHLRUL3Yv1ygJAiztqBgi62L8UZTYkMZIJva3di
VgAeG/1C2iqORphBd12LYCz1tzomv+MccFj1uiYvGMa67NLIxxqP/45GBy6ffkb3
X4in01pEfwgUBKtB0Cjewq5ofB+np/ghD93ijow1ZsY3o0b0xWBkKXNUZH8VpNyb
LOExfEBExmZIZ2QxZvsDhEpMCECvhaqbQF5nax5Rk08zqthPn49vWi5djcifJHa9
3iTC2/PbgLYk//dFw4dXHmPQSF8KkrBp4xQZ/dA/ECdo+AYyl0T+aarfZk1k/s7Z
06lpHe5wv85wKn4LRVQUlN/aBAhukBhIJHkyz7IuBHHrQmnOe4p7tlCioe+iOSbq
H5THrT8aX7Rci3y4tK0KEIJlL9VCM22d3LoBRMmoiPJTaX2WB54r3a6Viks98hgS
J35C1afg+EV6B1vABb3M14yyZ4j6613kPFLpuVDzG1HNJmBi+U/ayQaINFjJTW0q
SyBIBXAGF+YTJI3g7CIgUkhnZz/06hYHopQGp8fkxbMZ+0eKTKD4v248rvYL9IsW
ph0D+6ZRSXXqAB4lGeoK9ox12ZY9c97ffpBRga4kBErUt0Yf0BJl4sd/0qHxty3h
MgF8zGJMM8Gf4eqrp2p4+XIldSHMMmBQkb0QlY3n3I1MDZ0/R42D0fYUZyuhtkGG
NVCxO5TT9Y3aS5DakL/W1IKO6IJZOJ+E9yC5tARzbLXrn/U1wduDLWRpRddjCD4r
hJIL3oALJHzc8NoPzaWJhSRvHVykZxWhGEN1q4I31ziNwqXfV+ITLJbcxtj93SxZ
IfFZXRnanLA28SPw900IEKUsidWIDjuMtTzw++/zZhrllXs/DZd6PXY9aWtY/1rj
y/6WDSYSBSRC/yyTUaBC8NsAd0nYC5Ri4V5ETSD07rUMJcRSHT3/nRhy/jgMSdnZ
FOzYMWTIDS4YsjfnKSGLN0owVk6KN3vzZD42Y1NIKhvaH36oHw9GQ9OY38x1leu9
669zvzIzXSAZWLZzIp92bEIGWdk6JiA51NhfRgJKBHL8lP+2jiBhNx9Gt8bOzDM6
TqY+drqDMQ7lULrWkxgc9qcCVaTNuVCVXbB3Z2vp86feYQhl2KySkf1nSISPaoZd
rukrQri8v/jOa7Lga2qG809CFhE71FziBwsa0EBMVfqFd0iZw05jL6pqTAvCBJrE
/Qa86hjKO0LHohkNLlVYJkbyaCLJJDSa587kbNRdtcdlOFo1I7NhT3Xx98cGvRki
Skp19PKQCILEQOqEtaIX3JRWF+C6QA/Hk07YCQDORakHsWSm27a0fhzTXJb3w9se
sPj1AILN3YQyOI+daqMoaRSPq50sr2letBNcR8e92/cjxGsnocsp+ItszWcnif5D
B6j9jCsZpUYUb/ya5nYQvhTuRU9AQ6nUQJDs3VrG50Dv3m/0xMEw9N8ENtZSJSwa
KXroB0KprsaQ9eGsQuyhZEoLBBxMcxr2nPUwAnxX8nrX6D0Bbp03wvNncKT1LYPH
KE7vltXE+uWIzuN1a5qcGyKQf7M7cK7n813Kk7FXbhz910+bD9jwZ6MEE37IhevH
isHKlyDR37ul/IsZfbOQ2y136qtFD48lO+GCotGLujZG/umKDvJadG41C3xHzDIg
xg7jSTc1y5brlVDtoVERbMpCCRSDW4bGxP+gag8fgx4Cum9oASDChPvCFxgyUJ4L
2Z9NP3A1n3oGqW6NuqvwjDnNK+FVQDF4sZIEJblKPKXT/TKwkYdPcaWGfu51s+wJ
Jx7L2R/NPPXxh/Tgi/FSjREa0Dvpb87m5AAW32XbluILFH8c6ooMyNF10lf976Xu
ChdLFlMlE2WqbCMFI4RfOjBs1EvQULxFTL4zkmgtJ3hU8FwXHrqFGjDRCC9AErDK
u2qUm4xJVYxlBgRZ4GFzDq34aQq0awfQvMKy56Pjjpw0rt+fmkuSPgu55W6c9ent
r5O24s/84S0Q6HgldMN5CSAke7dEW4B8iQPv8txHQOhxa+Z7OApGyt965eUYGqXI
ZDwn0sMdjEdMbTPE1XI39WA0JLYkyyh7HOx+YjDjRdwwUHiJYOpW32E282lm6cw2
aQczdRqeIEZL0a080Gdp7uAU11vkTjJOwJQyg/6BMaVOzynj7y2wv9QwVOMKDbgS
FfudkYA4CtBX6F4wxrmbRP0AQYcMa5RWSvLwvty6pDPKT5MWojuyaYYOHDWEIes8
sSqqlN2it7mpRcMEY7/On0rY1Xx1czqqzfVL0dVs/Ljftx30I2ylOYXjoZdXDLar
eMbMOYyuKsc22LR/O0G8utAIbcXIVcigzq+UciuFyEee5Y+V4Sg6SBRn5H/6QkF0
IrkrftP4V6oJ9kTX35wVyNxLUQIQc3MgklEYaA0D1n9ikHsIb8MLqXHZU3qMQp+K
rr4S1c5xj8S4uK6dES7Adq7MiXM7QmjQPWkOuYa/9DRf+RckPg5xOsEkblWD5E7o
0QxOI1dEELSsGV3kAWiihfQ9csOfpYUnZD9fAw/Fcczu/VqREjV5PlSc4Fl2NzdZ
3XpkV3Lrs8uEyGREm/IXY/1NuPsnxlFmzhBSaStCn8no8Gf3rLM/qCXor4p8w/Wi
9XLyEVy5vsyKd9J8dk98XalbD2BIc7Y12bXs6G8lSquVlM51uraos0L05yf5Ol40
03eUuH2dpaEeKTg2e9QLh3l4341Ab8oiZWwWY7j825sKWw37uv/tmekp8p0+bNe9
dqEyFl0zboSxkxB4WOyry+F9GoqmKpETEuAX9Fyqh7Vcr2EX3c2QCFiLL9hlolBX
+NhcuwaR4LifZQyRIFC1PbKt/ezap0P49LE6B2coifmhbLHDbnGhzUOalaJoezW5
FAQKNssvWNGmuAvW0cLntRZ5hKfU1igdKYGFsZmakOAfyxn5/Ke76xFFOZPxfh6w
zyPafHuPk43c++yqlgINIK2PvhLM3bIprnh7/HtTLPQrQH2pr8ibmd/E20ErLF0E
xtsGLxvUU41zEAMGIC+dA4rReb9j9iRFbTRf+DH7pp+VtmITbN9qvMAVoLkPaKh6
pDD4UB/77Mw92loGXBvKOte2eLxAeCoDfuZZxUffsd6weq2G8SEkpL3gUVXBnnMQ
Q07BSOAszaGW08HaD8kDBy1RntNYE7qZcShy6j63VwanKfDgbneNZCXowmWFKjP3
HhW7hh1tcU8eIx0CbOfMuzB/mwQLFeZoun/+dCQe1aL4RqSwOmvDJv89iyIe2kUa
rHxCEBMpiNc6VQCdZbdHq7eZSoiNvmaOp3zCjVj2bdeYEanMW/BJsCrHfbpTzLu+
XPvsq83JhosF7cdQGyct+r6/Jf8NFu8U4eOLF6a+hPKT+5dI8eohnIn0S37Gldif
L+LOCq3VWz9ikclycdYegBWEZRJ3XbMyk8iitNB4yh0F3xypS+gn6CpsqY/0WrwG
KkjG69lbYUN4gg/kxftsDbO5ycQEWspf+ilLNRu2s8k5/yFEoVGtY42rDYVwscbZ
V/g+FhjhmcTWNbRqzl+LhIG+bCFQBREvc6JYIoD0+fELWAYIzv6KNqnFyyWg0rKC
pKprrqfk79J8efEmcA9GNztQm4OnqUOQdz8e3aNma6HjyohO5nFOyX/iPCiKPzjF
9Nqm5Yo8JKUemsKdlCCwnQzIG5kx7aiobBkwWtaR1ylm40cLbXYkDQEcK3374snI
GouUTSeiJOXED4z046k6o5XHVlIv56Sh7G8Og74nq9V/gjXMt5Rl8Bh+rtUQtcIM
p/WnvSzr0T41xBPt8ewu0dnSZ+4Xitoe/HKd47zcpvWY343EftmuL9j9ZzA0xaRh
tWpFcF+tOkmTDHPzwmcGVGvxASyaSifL2pJ/uQXr0Fr34a7luWejQAqvu4ZY+jzh
DlW7j+pgblo5LRndfu8mmM6h0/4aGcuKNLcIzW5MIGcLQdABif+a/+j8wPzXwhbd
pSw6P5Yg1jRAEFzOOo9iGHYxg4DpeRNGc3kGrYdqlmofbfb7wU+H3xVYCfvj7DDA
KKlSahTo/fhA6fN4dJIbTH81pkQ0zwKUjWvNQrKk97jaE7T20muoKbMp+Ut7KFVn
Z+NUxWaSI9365yFZb7gbNY5cCOEQgRlolY2VCeStEpl+xJDivihW1ia4dfnGRIGC
jl1yt1G8cJ7/u6b1D9pa46lgOhB2+86N3xtfG0k7RX6Vo3A/bUL3HWY+zTdgyHjA
ufuFOz4Frisw4smAziboAxuBlYw5aK72bAKikvwktkz8Rj6asjWCarCR6913C/HT
G16Sc1plWrH3iH/xYf/uGsKrowP8NDOeTjlk6H2X0Y/PKUTxLIxQSekPMn5MElT0
bBAvH4UaoyHgUDFw8EGFSV7VA5tSy8E0NB+0hEbYbBjAmMjJv9MNd508Z0t3PEYg
05zZvi5Azo1fuKa+/iZs+35doy3U9rxjyYv17mlk7Us4Mg3u+A9j9jvYT5FvSyJk
wqN3elKAyc+hSmrjCksdtSiuqrkiQv/dgBB/HvxMfyCIdhOQQUfnN/vbgkYg2EDt
8hP8NRq1rmBnqdZ4n/1BtpLSvVX7xiZ+x1jJ8RxMlI6fJwShMYlIgq2/BoiYZw/R
o6JzLJX8+P1NIOV8Of0w7PdajtIJfeOBqIgmS14DO3q1VAuxVwi3gN3MCz2rgQwj
IigUnikg5qHBDKRZmxFrAaKHr7fLfxCQS93JaQwsFfwbGKlITs4CkpPwzfURvD5M
8IXtCX60MpvEqsbvzqyxj2j3gG+B+ADweyVW0wzL9mE0svB5UXmNMskHa0+MJuJ0
qiNj9VCkc7exp+HXphgYG4P9phGNPLEFnsmqYUQcR/lwBQqRgjP3gkoyI1snMS3c
2Y6sm8emjBiX0PRMMl5e5azb7u4SVx7mqd6jp+sP7NDCnEmJJubPkj5DcKKWM6Xu
mSXOslQwU35rsD6Cmp2mVNVaP2Ey+a+g17mh+apGSed+voMpw5BNP4bl2FFRAimZ
wh7clpDKzRf4lIESE5X+c3L3XOiD8D+cHuM64dWeTrvQvJq84m1cN6vImX4FyTIP
6li9F+euS3whmJFQGes4H7ankBseuypyyY8Z9YXSOgPOKZeXWaF0/5Oxfdb6c+21
xO2luDC/8A+jENUxVlCXThNeIhQf+8uWNFotlWOYSk//R1w+WrP4MuEOurRlLGSN
DqhVihJ8lgHMJ+V+f7hno73ljZG5bWk8feCKKCCzL1Pw+HULaDx/I3wDu+0goMWm
T6ja0BhlPds573GitAaMRSXzNXAC3pzNl+0tn+D+0WvAyT66vBg9K1BrCIpv5TT0
B8hDKupGXoCM0VMdOzR1EjN6OE0vPYlgKbaHCW1ONMQKlBLLmjmyEtiteHIzXUQy
VUW0ZmAroD5QF8Ke3IsDPRuj/hNYWVLKX5P4Rd6nBrWTu8ijA6dIX9VHbM6yFD0W
O3YgOvee99dQ9aDVBk8B4/woiA0H4U8aEWFh1PKFEcdNVep22yX0B1V9zIJEzOZl
i6cxmFHp4R7GIs1SdqXE+vOJkV2nHHWMZaK2xfaE6BCTgnKbUutR+yA99rqb+b55
4RIryQqw9WlJSogbK8uEQ2ufIKvid+IBL5i+SXUNR4gwZGY99M7R6WpQTHByKPii
Le27xmLtGFw6hjZ8TbqpV8JGATt6dAaesa1k9IYzwLY5KqAH76Rp+wT5XFdkR2MM
4DYgKnktD/rPfU46pR6yglX2aF2eg55bfzelADWxozivMP4YC+sgS1oVH9G1RDRP
U9oWy+tW4JDiopngBdZ/kQPzrebLx7YPfvcbbVQe788uha2G7cBvDqfOKUQctx16
M1CzHZDvjnA7hO5/xp/SGVi29GGXfn6sNczaWo0LQFrU4hOwa5pwzVcGlk5eRB47
5aCyePWX3PEEoaEdMX7oy0THEvUue8xvmmyqSOhBPz0DiRUUNMg1rTGqaTYZQKXa
ZV3qr6PzBsLC/DOPmAtQToMmNqcCeTsiCf3rPmc/RJUz7/MkJ2nCv45S7l/qdrdL
TLM1GCK/1hT3yimFwE9CrnUWjMJE4JNuxUxAAWXlqtNhh4xTbbrWwoL3V/Q3PhKv
B0YtetUlgD+C7yqn8DEmrbvo7DtkC+U/9kFEmhnuTCybfhYIqhb4Br0oXGkoYyLf
pzVCmzOuMsP83eLQ8leV1PfdEpMQXEqtSRlCzax8O1ovIZRFYAKy1QQ2OgQPcUmB
5d/T9vrCoWpREycnWBTy00lnBT40Bvb/RrdCTA/V4ro7CLQ3o3a7utxz3Djye78h
IHTfaTn2UlqqOLaP3NRzPQctDZvrxUfyXZasBcUG5B44FD46Hh68za/qXd/vZDhm
p4dipZHN3kJojYEPakr8zBmC8yoHRm6qpLDXtC/hXs79RaONO8liSYyNxdaLO5oB
kNVHChn2YX5AlSQHe97uM4F08MylO/4vxXzPCZCkyxULyX+J2j3SQktNdXayO/o5
ykwtv2oemccRnQCFl1WOiliIBcTlfqwN+EZ1uM1dUKko/mVIIyyoRInlJRY1R2P5
s0P7Wp9pcCfg5QeVeKfJB5dwRJkbLBw9PzqW0hFFMoSUR8HFGaD6PsXoUq8rUCHN
d4FBuyVC153rHzItpTnS+RhGKr0kQD6srMkpOxw4jvz9uo3GVlwK89BRcyuCm6pT
JaFLmQrh7TGratB37qT0tcJ1MGkYfCuUFpilG34CLapiLphaKdUGF19DOxlbnLcY
mllsKScVljmEI2B1hszNaTvYknsEXWFXlnn5IQhAXQtxCz1b9NtvId0Jbb5gRlYo
i9UwETQ0b0XDwzkm1wiRypk0P1SGBau42jLFT5jV7jmb9/CophaZAdKAh+DKteFV
BKU/5iwABn1TP/dA32V/HdSArGBTc0elbjFbVEr5co6WWlNRghc1I0uAawyTzZEA
l+jMhfgmQtJq7chddU5mhabGTFd121G+HPywMFbWU6bWK2bW/t+zA22Cnz4ZTti8
EHsDgHQP4Wad0t5eY4Bz8sgyym6Z/wBEwItNpvA7nTMUqW0I1T4U7v4UCbR/pXmG
Nmd6RIaJwolc3FXEN8FRhd1tDAPhbqdZpEIa7kTRNoDhq8ezEyJ7Tz12vtGQBG9K
ICfZvOIzV6cPdhI80pdcusX0AkzipgvFLwE5wmtRJt3DqTHiiU2zYmK2wFb0i82c
TaxPQYKYQlgzAbfLUFotdcsfgfNIrjajNvNDtmMF8h5OoaNnn19OuaMTK1I3ZpIA
xsUC97SbnBKcCdqgO0EgH95BSV+ZLmCkgO2AACjjW32qvQtIk5QDSkJ88kIQrKZ5
H9xeqgMTSCyv2/6fJ7yU4EbcpTxolkvogeFe4dH4Qmhu4iUk3lfvJW0W5yM9zMCR
6vEDX2DQVbMwvDkzHjNzvidVjE5F8oM5s7xb4hCMjbvoBpb3Fyof+W+jRGAUJrPv
MKkSpHUkhVhiqjbtOo2JBDpkzQ6dtw67kInJf2wqZ0VSfJXmk3SQYjzlHwTeBJh/
H5ybHdO8YkEP2yM3KrBeii46m+GRZtsW1N70Q3tVI+39DHZZ0PRzEUxUF0K//juM
R9leFQsS70XYlGf1eoYPUuQj7JGmGPs65ZLAh21ql6oKcFpXK3eeQPLKJJw8sgNR
QFXiwzC3M5aizSLld02ZakIxwqSHrzFGtC+xiQ7vefb6w8LXiLG6Gny8OMdhIAbS
a7Abp65i+rqm0JkJXQDGL057QxwMjU9dYWn1yedxw19qdhfKWDnxGJ7E96GVweNl
frwv5uNKilFGfkaLYDF3htSCPJ1HBOVO54ieiW0lB2kxYBnzc269WxqYM3ljMQp8
ZCg8U1nyh8HOiKlhEAwhUeel1Qm3MRuU26k/L2mKzvv0fcvz9B+JE0noTRRs+iMI
Il+uymlkMjumlsFO64eUHiOgbNhMKML6HqnfOKmYHHvWncDbw1i9lvPCRpq5oLPn
rtY+rGhtdV60loZYcNmkacyVvaXUzHRvE2iN3zcv+1Abt9RP6EOIKNFd0zVzL5jW
ywB2olwv7jWyIM6HlnDRM0PC+f8dYMOXpOf2ZDq190EYWYlX7de+z7ZYvF3/09zr
cnc6X04mkL6hH8ghVNrvgBax6TObuqWn5ldqujSqxapj49pmc3REzatP4fivphUD
U2tPrZgHnyrjDsEQlAV0PprNlr3Lx9q3G4FlF0zxjAULtO/GmE+q5X/pOG/e8LT2
5zjI7jfK/YJ12dgnAtFVAQ5nHyKPFaq2+kwpxdPwlfQCfEv5FCY64MR5UAZeCq+b
tUTcGMOk3FKb1PglNGAK1MyW5OY+CzL5os4+g4sAW77JNRNtIFl6HU9MY0rhVAci
R5IL0lAPjrgInvb5/x78k42d30+VjqNr6oIiUxsCYt/TXR249/9wWqcKisEqEYji
EmMxoluw67l0mYMi3SKNLVLm96x04OGqHuI1crWKndiQnPlWM6mWN7UvJv+Zu7Zr
XWkfzpDTeFY6EohZQoP7VsYt8GfNveTeMeXisJGj565rabcwsShw073eZuUZQHBX
ags9CQB4DGzsSZSL1ToyoeLzMtFW0FDx8P7fKyomr/fD6jYBkz5xGCmhN1LyN3BQ
25wUvLU88Yo6/DTNBUDZFTkAHq8iU2rVvmaOnpL2jAL7mlDDI8K1GWHKQVIWVVZE
it3dAXAhdUA359rMaCRw7qk/L/tx2HDZ832nVUOTTJtvOuYmufcMfmoeTGRoGQ6Q
bG4wPA3jByQwQmtlhdlevJP6KnLswTjQ2ynsxxx5stXbOqC19U0sPs3O7TRmghyh
N1kF7MaxCtYTOU5p+lssiqOR5x9NwsBRgqENd04f3haHGcxKwqrU7XHiLJohhZt1
vhYpi79ys9W7Aw4EH828vwtIxBCMcVPhVQCqlbW5c4JKSQBbxij4TUAd4aosKl1D
WvSKzRtcvJfuBbj5fz5Dhnn9dSDUu7sp2elDuFtxQ+tgRtasVflrAzXC1tLHAGom
k1cY9T/Vwf08+smoFEVHoyN0JDV1ZlVRB1+sR9HkYncgCUjDBSHfB4ejrA0Beuik
+ofeCeJUkkbiNY1LUkabLd9yBQCiJcRKN2PhOcNQpBfKTc7iP3/z2vKhVwLt4IYs
BcQ1y7fh90zT2rHfvbgULEDlw4n9ajREWw/5Y0QuPkFdvY0sUHIb9/el7sph6x1S
j8f2bMkeGymsHEkAP7ydFWhDHSbMNHPwGGOgS8XffuFQWp0wxGrXorVtme8BLhXf
4hV7wd9ljIc8ycJI39SfjHYKxT3gj7eqlZVzjX5osRIRwwzwY3LM1QmkNlA6Yjl5
WHn8CwBBtdgTpgE08lXWdNkeBaIWjIP6k/nxkvBek18O45XZCGPCS8JqJQXyt7Zb
9+gKOCeig2NJ3hCZo+fPzabV5jsKQM3oVl/Vy6LyGQ1t+CIDsB9WYSIWnDnyyFnP
3yXRjTByhYS1rro0ltqtpp3li8q0wacTO96BjlFe7BRmx1AeG5O9H3K8JVt7V0BA
Pfs82tWewZQ+S0pDvAz1DJx4tk5N0ViOrfb1oSOzASipaDK/6BOr4FikNCQk8m1y
U6of7TigqwuHDSSQesVt0S8acVQ43HFcoBrtCcYOB4eJj6pBWw+/9rM5rQb83Cmd
ZWr6eo1kgsQl7oYIhJKleT0xxlOtE7M0ZakRKaS3JiaHIMkFdTsmD1q5Byj4NDFH
rJxzjflS9sl6zD6+vzL85zm9spwYMcxvaCaG9pGokKYHd23zsEe0mcrlvIn1ik1q
6tzvQKIUcSAvB93lSxqDuWXG1lakCB2yxqwQbjeWoAjaLZtBtn5XHwbljF0VaQjW
hMMl08L9UPSJ41Xp8Fv5crqh3n0AZ+GQNXS6UAA2ZptrKDfYicTCiYL2pUixWmjw
Iw93frpr3yoJzW0I/7kU82qCrqmNlm914wmKYpn4iCCF3R1skzyVKhe1sxd3QQO+
Fkj9zqUFZOdZL4fKIyRSLC0x+Y5M78gTzDsZD9ugGUAInrcz7H+2oqbXruyLZiqG
V2BpLGyX0ASpf7NMRjQWY0+okwVdn14bHnYJtnLFtixocj/g0I4Gx8qo7eZeK2sl
FnoqEb/G6Av4H3TU46Zba3xilo6MoYrOF+tSGMLhE9ymb6sWKu+hdjaiY0RUrh4/
Q1RPS3SBMENihkHjq2z8Jduk7olqNlddSOxSYF8S6JVXfZgo8HzpMXWT/OU7CwXA
miOxnyWZClfMVEBe671nDAkOfjeLgdh3FjYvLgoR6Kt0C6+qxrrtzFd2nj5mIBIv
/pWLe6ptwLK662acAekxD5OPPtzrA7aKZ8NLEwsSXE3u17DKHGXTNHaktZxkbKqD
JxCJdu4U0Qu1TBaRW4wYNX0JuqAbtOltC+tlsYHj0BKoXQmuDlVxVHACpeTPAbed
RC+HL+68O9bABGJcQrEcLpU1HBbuetnrjkQsCpphHE4ob7HklFwyvKCdsT7CyVpg
+4lZW2ttw8trTg1PZutc2ckUArMNv9c47itWFlDRrtYWM6mx+UN86erJE9GNsI2Y
qDJmnBgbKev+tHrLLRKR2Xj2rxC7p0mr54DMPsU8fiqwrvyGncpNhtxlddaD8NNz
XMk2KQplg2/Hj6K5aCNmAhCNGSKrWKvFX5wqlqgc28D7aXr+rWhsBrJmV5Ny2j/4
oBguwxQ9lpDjOp9JkybeQ2YRGwJPc1+N4kKo3fEm3Iyy9hBelzqWhrP+reW054ey
Ho/fWS1wkXtLkQ92GtxNThe/jfc5RYkHHXnetDV0P1IEka5OFzKvFD2f0z3me4/q
J9LpTp1hMvLJj7a7OolN2KeEHvlXdWY0tU/r4GSPFvw55ODMaEP9GUipgEswIE2x
8rx7wjuZQYr6GkqMCW0c011X6XQYnM73dv67Ty6he/Ie5MfZH5LtUwmyskT9FQ7X
kctzuaLHu1xCcdxTjfECvdgoWgzAbcGpfhB07ZBB1W8PeWeMFEgiHOHIExeWUwjT
Shjrm6cVRZbf6qziiUMT2qUOj7YJFqbaN/bEnQ80aJDyWVXHtJ7ZZcIFJMDSmyaN
FLnl2Ona8wsOmhtVsuvTQnjnZDm4e1bNPB02SstgIv7enrXqAKF9R7BTJPFE0zif
ildjbmrUar1WA5ZRd3MMiyd/pjI2Sv2bn095Ag9jxsAuaJ8nZJjieMvOnOy58qio
ZPv3aYQIegPexGDETV8ovLJwKEB1btQ3pF7qjRa32FQBrEH52gnCaaDqIw7VURXd
OBGD3XFLOiVDiA0uF8IGCAZemIRmYUhusXRiW7NGqRh7gHjZCc61YxUbZoaFJNJM
mYFCoJQIEdfZ5FJ2veusv/m5Cf67o7wXQ898cmOHOAO8q5YV9nTNVfHV65voNVqR
cIB+pxccCAIpcXO6s0idJa5CEyoF2DaAnsUJrGseAZU74cxlCwsl4mTrK4wLxboG
72+C9P8Hcl88x3Vc6hRYXGVot767qedIufTILccEhf1SsUxwS9x9SGNE/ufZrz7k
2Bm5fKspePRa70ljJWFvMFXR1c5lWdCKm68ulDRGiwDWBA8ZOy0wRD4m7J6oUmHC
u1eDVe4enzLSNCePVLOz8fPkOFpM/MNvIXTsca0w/rREZe27/bozZ14AR7Y7WHDx
r8uKSNQqauwxU79ZLjQ+yfrJdbN7phKLPPjmiYigKm1xAt36J77TIsizf7PQh5zj
XyMeNvrtjrV5sHDkoxinwPJdIt89wEqIgn1gxROS3004QBRQYiE5lSHkEYnaPhR9
b7NE2KxYxgasTEZWlPaHuM3pqOlxb/J8z/m8nTHM9zVyoUGFKGQ5GCRYQ/SCTmCE
HQJ/llxVk7aQwOM0Q8utE8dfPR0pP1TYo28hAa9P4xjjpI5IGzwa9HCZoYJ244df
MXRO6jMrvrPFZcZPYDM04ksSSadhQGA8FfdcqjGw1qtonrOirJgBoCQV0Ah20bvR
S/V1t9DjHrmYab5mQz1tAytUc5cMFocIwGVDfkXDHFvGDvYqqZy1xrYXFSxAn8IA
nT90MAnFBelnpc7V0IUsLijWEXwU7xhU2DXNT4xSfJI1hnSi58WtKW0HrVMez4s1
SDbqDaknWZg/yi2vnrnzcr3gqTSJ3HQ7Wjh64XutpA5PIMju4LxKeuw4RTO99LQj
6LWfgw3P4ONuqCT+7WAknvhmp3cUT9mqPc6w4OTfab7f1/IwDmb2tj2a6a6VRCxt
jnL2lx1MAWx0OWq0CkT+nkfRdDV+8Y1Jn/WaR95FlqyPvaDO98Ypo84zPq5+a6HB
7AcjmOBAEmruLM/UcHvhq1/0mmGHolsuE/J1+lER/2W+jo3/p1ZGjmDnV/o3Wgxq
r1x2ZmF2Mw6flUsQ61dJmw7LkAWCwRBO7uVumB28qGruc+wRa60SxNzFlbMkMm8s
Ec3NQLKt57qRyjKlknBic71qCLSDeT4P4B+5z0IDZLNNjlVJbroHthpCoTZf3XH+
Ddd59pDtQAnTCcNvT5juWsr3cKE3xZRdXw1lTcykdgBd9zKZU57XtuWqBndxGpla
W6AkITEeDhqYX6AIyTy2hdGDBooRaKmh17OvzBtCcVNkBY97s0hBoCGpytRu5+dh
nC1RoHtL+vIMabHnZQA8x7+sfF1QJo4i7QIUNSuxmlIqRtyqhQUM4oMAMAkza6Iu
XVVdVr78mcnIWkkJ5xgfUZfhy0svZjWIZseqvJsfEh5tJm8/EovCNwWh1z9r/1bB
pqx3THhcCCQjpgFUCqqSfqhEOMJQAG8bu5JZnHTMQjuCfbUhJBCbWO3ZwKQp0/wZ
J6n/PomhsS0KNJJ5bMYpEPLY7rrfVqtYs1ZqjfycXasNL4DBsE2Bmhzzv6sBsxOw
cT9jfnrFJ7fOTSaw8s+J42AZqNqbpAWpZLvWSQDzafrAmVqia5HgdCaDPDTQv5PU
dDz5Hyhu8fQLLl2HwrwlsIbrZVgEs9A3f+rh4yKrrDH19xVUiZVOtWeOc02SV2LC
ASpmjUkil5yb+aNmS4s5CqVbINNrThlpWGbQNdJ4kzCthmlf7uXRtsyH60AZM7tU
2KdIldhMyHLGgm2NUEnqhzfRmeSyOAxV283GGMeZGIxUMgsfZIOhn/B4qJzjWPKi
vBI/Eu7gOdm+d/Vs5Vs0jww5J09Np4XWFe8D3YB5xHXnbRBW2CUuSa6MwfvLVoql
ufwS9FwX5Soay5bZ/zy2/GNOHvQd/bF1QSyZuRXHj6vMXfKoIEYnYPL+JNk+bERt
eySqU3oHRANUanBZ5iws/XJ11qaeYqYb7LcXzLLSw89scsT9tSYpyoykLGfVhsjm
HuaN8i4MFVx5DfBttMmc7DsDdDslSgE2mEQBMfDH4RYYCbwopABwNOtE5Eh1fYf5
6fCowlZSyJv6sHvjf8Upw2vtn1t7lgGrHm7RV0vV6Vc0jx+Y9yQne+LQx6kw434B
kOS5M+uMydTjaOUPHk+fjAw2bB24p/1DjUoeCsUIMCahh3+6OcmNLXFG9DNTcg31
Jx/eJkl0KNcP46jzfuPGDZN4GqwQFBQVsycCY0KYWeVndcFxO1K/CQc/BHpIuNpV
pxaOEFgH9wbPiVuxXuQpIaTt1EHZ64bG9t+C7mieZmb8sovmtTt9kJn6exuPaGLU
S1aU3HA5c0L8Pv+YTQIi5F/ZBlv1KJbNRV8W2AagTGb42QJuzMTfAvBEmMhfoIXK
mFb4adtLpjVyKgO8wxoQwF5mCiz8ijRGsoCrdzMlwYhcFNkvRNduPbp7T5Yv/ziP
8hxjTK4Q2A/9PvzPzU4zwsCLhikjWVr5Z1IIevlDE1esc9vl+SAehfls19Ehot88
yEMqvW1D94Sjv1TCoX8yDzWx2jVay81AoNJOO0rir1/NC2cxZQbCiFtpmGa/aPXU
QwWLQ840it60QitlXGTL9aiqkGG19sGy1Pn4FEBCn9BsFSS/UZMYh8vx0cpjr56T
lMYGM6y7gAm8VGNVUevp2E+McYQ2H3PmDsPfL9b2vDJdmWunPohWACa6dmFutsUx
bvJ7prd7Ys94PPPicZFeknbtFttaB80ry8mF6hj9uKcEpE/Sba2+JpoNdZDPh0yT
rbi+/dBZuIZNzsao9bqlXw78CU2i8C1vzZ6dCklM2sr/WXGVWYHZ2OoNKAvihVCc
xTf50ICy2MxtTUa8vb99OLNQIO0YVbsEMMiW+fJRQwkb7vZFSFFwLebthTOocTiY
7+S5eUKLHRIWQDJaGdx3ZYeU1tqjUKJlw/Qbs58wIt8waNx/ovykbg+O2t6Pg5GW
MboVfbeET56b+nanDNqroboAFlsO3BIz+Usz73teszuJEeTUHahG8icGrxi2HR+1
nooDtzsr2+Js1l7G7EgEVFEia75Sc4ANCYawAJF+0HCH+dIVr+cXGzDZiC1ch0dO
c/bBvkS6EVbzeK2lmBaO3PCHy/cd0BQ9dASaFhOvK26AVqfLFX05hhu7+FxzMBj/
FjwEe8XzM/juLldiFk9+ciQZbA8MTZGLG0oTAA3vWe35Y7UcUuX3HJxo9eP4DReu
xwdN7+iKm4qYligKfp50/vEQz0hdQDxWt/nCAv5Z5MVtOLBqZ2Jffg0KVceHkSxK
YgMJ5ndzMqIzoRu66CBlu7AY90GkdrI//swinauQHbPhEgxBAz9/EnBuqfx5kOPu
sLTF9DMNmJnfu8j2kQMYcGzurtfI85pvemxRg5N95S1rrGH7Lk5Zrp2gmCMPs9RT
jA3VFqG7AnCzmF3ozJo6qsBZ1P4wxHQOOCqY3D0j0T4DgbStgOWhhjoEuUbxvwM5
QNqjtJy9zuCtimw3lxMKDbKvotT0niJHXxHS4Wn3JvPwfsNXj/NZwgjaswcNoUcv
f4FDdH8EHfV4IouSESLVGL41OgZ/CybQSIOxoRStCKmV/7C3IdOX7BygwK/ESCam
Uii43JncvqfTajF6yw5RwpwmIT6FDajltLRMVcgUNzkA+/aqqeQ486zyKyh86Nfz
S88k2P1Cet8vv1kk26/Y1h3TTR8Wk+BcMDEVujem81bGS5ud5UYAoHYq5dUgaLFk
mLnUNwwrZevhVxH6rUO4vSXgy5fM9Y1C3zLjgJOqYWNuJgZU1Hs6qZc2dr9T5HIO
26yeWwbexVPnnL4mwK+GIrsJ+QSe64Zq/Yqik2L60dEfDBy2blN+mXfLmIFznxXU
ycR+59SghybE+7wI+e9C0ARHy5MQ8qRVVx2L9dJnVyMaba5AjTsCZWhdID3t+Hj5
7fU03wsyqxafLwPKLXD38lSdVFf1Hg7yf3A12iWhWXnunldynJ4whf//HGzwJWwC
cPFdPGmwvoGuwMsitx1mngC+yTuytrMeNGAyqlrWdvoj/eKQqJP3COG7r0YjkfT2
OkzN80WrBmxt5wHifqs93LHNC9i2Yq7d0pJyfpE0KwDbDWO9wJcDm47RHvASxwzc
WBXql4ufNav3n24k0Xnftov765qC19r3pylziiW/AlAa6QR0/o8BnWlkDPBNPD+H
fFIAsDtK1pDQX7iqvrW6NEL44rMmob8Y4IpgT+xixfYe8H2W3WVdHUI8lNE0NFeV
UlhxPQnMpiTcndPpYaOU9Q4etjm7d+nQfOhKd/PdzKuaoGT73TWYobApTpZpIYEo
Bu3Z1NFUF9xkq3hSS/iTbJFFOURW1knC/LSZAmL6Q/P4ztmDyqj/faiQY7WUD8hi
6MQvEe6/UQ/vOGwcvq5ZawHrVtcMVlziaPI1F8sZEWiTn0GnXosQia0plDWMNyjx
MYv/3+OgKEOv73rM+WxftA2PJgKjbV9g+PYMFhhq6/9CwlqKjEKKhkFNsgqSeIEI
BoL0o5o2UkrJR/iW+PIDo1Nd4ZwiFaxsxwZUdEb6jFgDrFTVfw2t4VQzV0Lf+VYS
TAdMShHnZfT6PD6yRpaVEtNKCmCac2K+23y/GiwoGOQioK4+yZxp6cK83AOKXODb
9Ue8SjYzh3ZjZs86i3uL/ZU8HL2RhlAiNUQ073lsNTsGWZxsubFLFiXR5MV6iwZo
pUQ4ZrSWoJHrWQJEE7B0Hw8+8qXZpMNQnPLGs1wxSHht6KNmLIsK+lC36Fm3GvxA
TZaOLrYM+bycwL14T9I7wJPQUajAdtahFVnWs2vycmsUZ3aUe0x5e3HwtOLZiW5m
tZ9oygFkHWHEoHPScog5lqI8vKgOtCpgPuUVWMY/gB9P8zZmFqohTqTZCenmfUo0
o/0fZOibUH/DJYSM3lbXEPozQxXXuiv9krNbkewZsj6GBOd80hL5sW4EA1GSP8+G
5QyfVcm2r4w7YSdvxj5hS5lWG7+mLLPK0FNuu6jK2WrX1LwIgg928QXpUdf9hBCG
S+Q73VWob69jNUWJdn2hmilJSRzwqT0wXF+dqLQJN1sOqNpbmSuLN76WzE8Z+7N6
n2UXt9OKVMSEXEDukVT9lwdKmWo8kuLF3QgUrX3/xXpQIi4Vu8FY6nf59hq7miF/
ZKs5g/qN8iKs+mDrDsQ4/5xkvV2oHNXyfHssUL+1xQqJsxZP1uD/UFX2tc3EoHrT
yHlVVOeid3lPYXqtnXSTEdsT5pJtDHq517GIOsdhknaowzqh+CaNryeIlGgAdNnN
hXICVJ0B+ceLy9pMONKNsqFJ+OR8ESu7qd2wibEOqlBmGNCPP5roIOf/OTXF80p3
S4q06mcqtvd0GW17tf8R9Ei2f299S1fjc0eEx/CR2/GnsJSeVMgh6c3OF0QBLDqw
l7nsBwWcaW9RNDjDub1YtkOTlXp4dE59lpFSj3PV2F5nyylBudHwAjbWar5liry1
JuPtVcRQIgU2cpdkTtEyb/L5wjDG9W8GgA8AmHT1MffX1zNoJW9CNf7tFmRSzosU
26pKh6YGQU0OH91UJ0Wi1qJQqxUAu6ZBjPjheuwbPwY8Iy0yD76JRr2kf2CJnIh9
6uNogYJWxhzcaMlBqDVYxb+j/xo+sckmAyvx5Adl6RJfpD1sSqduVuhgLDCUoaji
AIAvKeG8YS/ybOax2BLE8qLy6X5W/IZBigaDSilq85Qn+zBIk54qHqMSRHAJGiV5
ksuDf4MlaRO0E3yv1EQ4HONO8qPrVgF97zlzxdSuu4tQfR3/iib/ufHSzbBKljsG
3qKHJKRrq4tsU6Lma3NtdW/O9New3GBnvzbLGpo99zgMooHDD/HUDYRSXl430KyT
E6Slwsy48SjTtEgwTcu5blD58ylDmQWvpnXftdtprW77rOVglkKiOmXvZ9DAxo/2
K6bRgHH9jIvJQZZk5Z1Lq1lkkXj2Bj2pC5bLWR/eigWZnG5ielrPAzoTd6hEuDgJ
alIdSFhWeIhjQDsCimkalFJnGfq8IVSlA4piMNW62S5VkO8wV4ytKKBNsLiE0RDN
L9/pWiHMWA9w5w13vty7cJx6Flw+L6/7Nf4eC9WwbdMeMLcxBnNoAy8tmbgD+cW1
m5hzZjivJvZ7dvLvzP87+s5g9OJwEkZEx3rOklLEfPOTin+w+VomHxxwrkz7GlmQ
z1iISWsh9MJH9XNOeVQyNThY3NUBwghA8B/JIwjUYD3WoxJ2oJuKTqEgCuJ155ml
MuI8hUu0N6J9PokoMskRXXzKiZDuO9C48mOuCf1gcZFf2qs3tZrko4IztoyzzicP
mxKcnagWbwcakrKY/EkaB0T5qtImqCxIn3fN3pc3hj1aS4bGUYsX557zVBy9xChK
nuw2CKtnQkk7Hn6SyjVaYlKtnkZ93B2DJFhEKhvkwfr65c7G8qQajUXfJ/xGwAll
oth2oILhcLQ/dnpbHB0TEMhVXUKoVDYotoH9SsxuSM1c9aa60M0y9T95KC7pIAMd
c/8BBR8QNvTxBP+pXmpIRHmRZIKOIWE3Sx5I9D53KzsEPD00ez39TrQ2KSqazKLy
GD91S8ejQu+5y+dAlRjO8qU5ZgJty22ae+0N3vWkfKMlZ7fuSDJWXJCIrn1RvbJG
Rz4b/r6zniztSJ3Z+bsDMGDruBNVU40ry0QO43DLO2tCDBeYrJwNxPOzPJJoT5zL
fHVofZ9WMUoRZp9Ke2l5qv+88i7S9Kl086mGvFHB4o05DmhAVNbzeCqEu2PaE56X
ttptij/TWDSyna3voXXy5owbW/61R4qj6qtCSTgdEqTJjsO8Hi3+FK3zgXYDLTgI
9SLJB6N544fIj64NPdnhksDHT7MGqez6VRUt+tJFiV/zmJfqYL8zWHjhiki9Vepb
YF5RFYdDDB/6F943xTVrzlTdZrbEjRbzqKxsH8dR6/Y1gCA1YkJwgWNOLQC86kOJ
NCDvYTjS8ltivL017qsZ54/MvBLWfI6vQTZ0wOgj1ct+0YCnfonBsZBn28TF/4dq
VejmKk1LAiCg0UqxgS/MB2Uktwf8+njDe6eImQF9f4KzoQ6uyLLNeFjpEXBlg+5G
VZg048j5PZYYJ+EiDdLLfWH01223WYxwqlJosBveqDEbDnNHXlX+RSotp33Wv/FR
uNZOmH11Nrzb1Uh1wpHfMv0jjutWkCzOg04dM5qrR6CZtvnHD32DNsl2LTRdges+
go7U2SwXy5z8lmwE1wrtM9ebomtKmHyydFhx7GyPDMT8mlwaKgzVEhF28uF8i+jD
mkfEtTp9ss13aruh7PVokp0FzXz9UXlpyj7CGHkn+xO8lzLiO/9arMkm0M5widDe
07Q+dpkLng3JyW6YyHNie0BoOCry+kyv8PDlPenskziYR4wUg2DpU+nnSR6EbXRe
B0NjEIMbDw/FFs+cSN6/nESWufX4WkcA8vbQLGBnuTnH9rUSm6gcq92KFpqutuHC
TTennAEsvRmYcaP9gbavW2VSLZsGD2PTI9IctLGBnQ+wa9IgR1WVDuo4CjOrE+Z9
qYd0VFFeeMHqNvgwNbdmEhFYzmikR45kZYR6iFUMyNzCRVirUBThSJEzLjFQGwoY
E3r8vD8w1LREYO/vvHJo7fw9P481VrHFIuJE887yrpQB5b1GjCBbXG/c1u5hjC1A
sujRGKcnTzHj4QH6NhaM9MBaoLvylyTAl2wvIKih2sAImOzBftGA0T1Ov+mNRPe1
eZabMQaKIVfjcA6IqK9Ex1R0dT6dmQsGTx67ZeJtsixy47zwC9J8zstu/7sT3Eds
fnPD/ogpKag6j7rk9UCDuYKY3Lgf0SrorZpnp+gvTL9DFqRFx2ZJx9gynm7Yr0Ht
AjaswtfPKzDTC9YDp/x7BW7ADQnOnSaSWqn6emy1cDv7vSl6TxUeOpg09CafzJli
Ydl03pfW2HHwHjr32qhN2r6CVx5bngEIueM0JmhQSaX6mYSjUWzBA69kt1PDnT1Z
Xvl85UjpTtFSeH0/eDovkvApHrDXUINRepoVqplMc2cqETKflaQcgH5eM4/RlIr/
o3JFO98p2PtcJKmQQ2mKcy64ZLw7Ec7aY7JxJ5IMAGX5+5ZS4l9z+9ea3FU+l2YC
+squtc0B3BXfTOJwhCdi3X525FT7wWULScIloFjo5r6krAeOE3QMXT2MDwHv+Hyh
WJpWX55svIH3GUZ2Z50rKvD434X3rgqfri3A5X1oyRe7laRRpuL+6rnRQk5AssMK
2qM+xYHmfaH37tfd6KtEZZmQAWLpIwNorY0Wn7U8OE6+yDDp/cx5IfcTg1xjddF/
TX8I1kxr58Tvcj2++LmNsV6vnMfV9kS2FAfzY1hnFbPcdexxcfEwpZ5bGmOn2B5A
TeajjCJpo49X/KP4H/VkKfg97qG4Z9RrYAojntu+iIaN7oaKt/MSk4xW76hlgghH
CQK3eUdSqY2UgdXWdAmp2ay81xnDf/C839GzhTimkwZnDa0sqZEvCaQ8xYYnRCA/
/EbrcmPHgJr23KbSJ4aPLh5BJqmg/LHfZPDi1ajmM7TJ2J+kAEXImOJKFydxYZZk
G7qhEJSe/t5tdfpeJZhrd+yMDN62VexC/t0UKbz7hNiKG4DdUwHRAUDuLWqodj5f
h6LbeWdxfRKZUNZFGbePR0SANS38KW6zWy5DR+Nh9EdhgQCZPfXkLEJKuBM9pr+x
rPGsEgCmWBVlKHCy+8Frkqg+RFUDNe7fJ19y9A6KROZ1z0bzfFdq223lEDk21IpO
iqUv61o/kqj1cm6EP2/QcpKi9DwR8u1I5Yorozr0Sr15+F8xfSSWsFqCY1QCAr2a
I6NgE9HEqbybEmK6U3MPO33f6kgMR1jVW4KcCp0DJj7Gr2WXE4/AS2Q0h/OlGFUq
gbwli9SjqAOXmRWVavlO52s1eGZMdebsNp026ebhb0Xk9HwsDrc/KziI7DU1eMHS
1Iyel+wn/KxnBjN/fjupskHH1uv+MEKkMj00WM7JEEl9CfoArJE2WiLADxPhsYXE
H1Sx/ZRq3CwNOq+xFvOuf0u2W6qm7/bh+rJA0OIsos2afgYhn1/lV7Bn7IYaUzDW
p9IgoKu3uegprcOO+lg9/PrsEGNpqXtQGQ7rtRmu0pGvCERpdDMQ5Lxk6uySx9NB
t2Tn/vENg3O/avUzQKNkcaCwadrc5zmLWo0HFZ2fPrEEU88OBFD2Xr8UFgtE5gsW
fy2QKecknq8yYzryWGRNR3F2JlRJKpzt5Q66CNYFIa9xN8a/bV2GifEA8IKGrdUq
3mW5wSw+KMPnmOOh9D2GqJ89xjRT1I7HVfckCLiWt9Uou4AcHckSgqZgLXysrMHh
0MlHp5SPj7L6g/MtbS1zPU40TJkvj+k1S1d8k0T3SqgTwcXrA34Q9RLLqVLJ58mP
KyZOBXxSSVI1nWXueoslPxeDjVLrF20VI5soiHxXyDb4qLF3ntmdwsKu+CVJquYS
WtYwLgGMVPv9gTgtxRBDwpS5dpjQhlllg35B4RQzxA0IsVtw8lrtl4erOS8kXZzJ
VS+EK3WSL7CD6As8aNB30AHZtrYjJIqMZQxQmPBTTUHCULdjWdYsN8zTUV43PQN1
Pyzgv2P4XZTdGO2B2Y5wDL+qUmaYOpYAPY9b5qncW6wN2Uf56GsQN8TcyG41bg8W
NoMNow5dIwgqKQdgh/FCQ8FzsOlb8V93nXUv7oaRbe9RTALSDPV/Alb8FMOawcR1
uyEz2RA7UV8ykcLIGcK1f4eZaN4sKHH52UiZHd11dArOeeuZjNzmbU5OlPRJE8zN
dWbqxvs9XuGF/SjDCb93ugczt2KyVcKW/fc61YuFiSjufMlHlLPBopliBDrll9b5
rzXXlW/I24Sii3jEEWCOzIQkB5ukun9zv8soaxOCG5U7y2EQhQ43khlUvqE2ghJp
WItUm4WvKzB4eEIjaHkC80nvj8mRk7J35EZyAyolQrrGYT0L8lbMjfyd5r6qyiV2
hdQwEUaYWGtr2DygHahtWaEgwCac9Fq/VDIspg2vFq/qBotzk0mRg04kFc+M1tnD
8AVOCU3m/o2XnUgo61nJ7L+SF9ukTgQgpYzvz7Ndr92pIRInTEVyej2o2fwQ8WuA
2DnHtBvzReWnhrRUH8Hc+tfqOMRI7/zIoR3axJFKzP4/ar3bvPghsizlNPqL3cDN
0qdNavL59US7gtMvS/t8f9t6MZroxXRdRhwhQv76g/UgpSwJl/RYwPAH5OxbEzYd
d4ZKfGTH54g07vDOZoZC6wGCme6V7CXeapPezotBV+kmqsEZS5IQ1BfnUPwbRbVa
Hasn/OzKaShI8yYiSpaB9yPGsL9zs0TdlwYU0JP96V2ObOI6QzJWX7Z4vqZYrdit
gkjs1NNJNPUhQVjT75nCOniliRd8NAQvekHwVOLsao2JSTOpVfwgIG2tW+koth29
hTbe8r8VzDl1Tok6lbiZMdgKpUzymwBwN13BcsVLQ47S42Esj0M5dHgZmwll5CW8
AVvxolwSpIogDpEFfWzeCf5NpUWfOkuNQuz2joSLbwsNII6NgmNPbRTfWWEcN6rf
NTjHduz9CveG56iO/WT6cXD+ppUCFGAZm028i48oeggHkPq6CkqF85ZSt3NgW2Jn
S7y+M3JDt3tHI6rne6JEZqhdnrLorRRHk4C/4ZxE92MWnGrth6Q4OnNjURP8OCZm
Xr24zMyGY829eMxo0HnOOG1RL54PmTdm4a/crrZeLCbhin/bvk5Mi/5lE/JMlmdw
JOhs7D9N8oXgZZT5zBbeGN/zSxbHR5rpuGnCVM5tilslfnc6P0gTV5fkZxy2i+43
+47/4NJeV9G7WF8ZOa5440fBjiSji1+qsuVT6hEeLZy7TN2k8G6ARlPXoUWKw/DM
0kmB9AF6Ue7VOuiBEAFIyQKiDXNoC3SVHRYt/kXHzVZU9UHeEy9v89bwGAF/iQkV
HLKIuUk8Kxcp4XoeDyQ5s3oDm7VglEeTVRcw7FYI0kNSbt0K3mDW1buP9MmO4wMX
g0NWG6S82xAMQNLNTOnMOURZAq/TmTsJ5BpW9mJI1vExPQQXyuVfMkmZcF1QA/Gc
Tbmv8uP4YkqEko46AMZRYU5vT+nIfMlrhEy+zazFDS1WzYvw/2zwJ3HXWATJF2dD
+SXjnSfJuSe7nvzJfd/aaZ9PXrwinCoT13QJIhFqxgOSBjvkl73Hg+qNP47j8gA1
rzHCYJwJ2GAHRD5puNPfHUQb4FbIJWieWEOfUVLjON9U2x5z6p7yF2fv5FkuLajV
yI7R0PhsmRAbF60uknER4uO/n93CdDQlYeeA+7rJTCMkFIz4WG1A6Vcwlk4u7YL+
8C9azU/NfGWOuzxw/ginoabgYzxUYEp+Zy5BbrhjNtjhG0k7uuJwCTWInuuU5eZP
+xVq9RUpuEYT/COoSrzMyTHdHmgwLeYoyeyk9Fv6eJGOpJAqY4thC2ZJcTgU95Jt
8RS/whp1WjZIsh/GFDovQh9TXPSN3duuP2TeU7+HvVjrDoodYJ5HBTJzwKTnRtXk
vUmwcvSALZn2MCwvWrWpJHCOQi3JntocyD5i30aCnxhbYpCrx1/DSN1SSXYQHJb6
rlgL4/Xu67TaTPC651VWwPCdvWr1klhUBBhyJPA0ZYdCsWeVy4z+VQfsNtS8rH+d
ffx/RdBUgQa6mFrO5WMH/HiofLanGiM6UOlJBDZr5PPqSg32WVzsxM2aw/GVgviy
xILp/OKHuSu9bhnfmHE/ZZcQuCTzBHGnveIE0H9B9diNVTNcGYbJDadkk0vbV5Nw
f7mWnCoTvjSXU8MwyUFJekjJf+oLj6Zi2Eq6dzFEvFyfaJq4/WmQzyTQaj5WJ426
CBwYVOCy/eVTF7wAvTADkqUIJxRc7Y2FzBWJZdb5NQic0+aq1/Gd043ojVpIWfHQ
LhO8oGAsXbsb5JbYAAPbZAof0cIfKHsSYdZIG3mw3jMQ97fDyG0P+rwIaez2yJgQ
IGyo3gyGPpl0KjAosYRwd/c1ggLWeWeCdDE4V4xRlkZaHDBcu4OTIatxIFb6nwvl
4EngJ6vkWo07zKlmABFiOTzKsYduqvbHVPXIwAPD3qB3VsHGO9QkRdN7gaNY9etl
bjmQMaDoI3eX9kKYzz0yYqwFldUtbpBe0xNSnUWmwdoZBIwIrWMaK81nOpJMMUH+
y3DX8kKKDj2c2E3/waqi2K3+hWTKslhN8GqBZ1cNPfd6Eu+mQ5tcFMcDr7uzZ1uz
vfONW4oXA+Mdvo1/284UBPfvJl5tkm3ylSNxLMekUQgw1z2D1VraCIdITJP8pw9T
JsaJ/P78nr5mN5dzo0BbpvGzxrFoy1N3NLspaqFnqcL6d3XfRlDTTIZVNrdyAGVG
JTQsWNN+BuT8EIdf165GUMplnqbnAnViK/Ro9bjej/N0/IUR2703/o8lZzOGtLHo
ECqCLLeWmsKnWJUIAamLwZFNCMhoDVcct10NWJBExhgnyzuJFSI/B1wYjXf6Zc8/
QoVLHpaTZk45jQ7JKtf6YPi1z4RVeTf78OSR2YY7AGhZCNA83Mm/OkOOtdNqCJer
cK7qyToYNCK4CuYyx9NuVio86vjWaci06ec4kKnqRN71K1gjL44QrdofefSw4g2u
8jhmeev24tSFBhw5UVonRxSREidxAZoc1SudcRPzN8Ih5huUNgGdCubQzUd5fJPR
tA+os2Z/87TNN5PcyYA1BVu3eO7Uk86LUVtpouRudm8qtXXUqNjtMnIMm7YH51AE
cfTSKLsb5EFQ9m+yy2bIZRBmW1/AzpbCGhSHH9gOYEZ9WLhM5Vtb6m7fcFU9LMi4
qlP2Gb6X9YW2XMGIXHEYLpKrXn3/AD8OWKjpf5XT6rOETxnRsdAtvHnsRBSVhuE2
q6eQiMFKhsSIIX10ma0SqD5Any9UlthmcunPUrA5k/orfIiCUb9m9L7l0OFBdbMl
qsk++mb/uzCXgMHZdgVrZzJlfZTxr3Z6cYnoOnINFxY1lnvnkiwPME36XaBTmnze
8R/5qZED6sXcvXnq7gUYuoCMYiL0h7CCaFRVHNY7OYupEMmw+7f6JUco1vKeDq9D
3fArbHhTWwim03IfMvfHvmxcpkqt3k6MmZuK3oxSziqZ2yD1Df1lcr6X0ihb4h1B
tsDt7bzfasJZid14jB/LDU7hkqU32h9vsVeSylW0+OuqG7pRGndCZUKSbByFxKXW
XeQNwBM4pdyY6ujwNaqRumTDa1szEGMFmnB07GT+ofCLaUPf7I1Mk4BCg7cq1MhZ
g1z79F/CzFoernmWwoZ5LfH1ma5yM8Kmfz4KBihY0CnUAh29s3KoWPbBvB7UJnm7
RjpSEeyz+CQJbQ2H1suEOtv1b4DlJN8u4YpTG3d7w0bCvqdjU6zyGP+mTU2WCIko
EfRDUmtT21FebhxDK0nBlAIwyLOc5aVPEfdLcvYHSiuPxVwB3KkG6wVVXbJuLxGE
sEo93M6ZaXJKOnp4xbMvM3AI7KLrd+gbfyfG38qHZVnjNCshrgLH9B34n+v7MHX0
j0mQqVOwnDisxPm51skLkTTXY4GgaCCr2xthlL22T9UEhjUKHnvaJpV95x/pH9zy
YHoAQVucI+cuDKDhleK3er5DdONFpo9zbZlV6VOqiFRM/HiwGn39JBJbnHbdJ1n9
Wfz9fMt4+rgqYI8haYzgB4OVZzuirR2FAsIveTw6gH18Zrck+0FuJ4CKu1JxEpQ8
Cg/p0TV8DyiJ1GVjlA+M9etPyOlJewhpnt0fh5zfI3agIkr6kKgfVIHf0AV6KROe
+YVVu+qHMObHcnsVeJ35p/ZX0nqP+ei7FlLyKlpjQ7pbvGlP3ZdZURB+AiPG5qZy
nQ+d4X9wNoQl8AV5zg2HcG6sHpwTpUR/S8VSpKVYftIriXcF9VTXhfp5ivV6DVNR
hvwg6CIfobLLmaZW8rgDZhDLmGPH9wtF3EEfeSjBPeeIE4dwOoQX/udO+hxbdlUz
8b7Rh43Uqaub2HnZwunichmKFhzJAAF323eJLia9IL1MDvK47CcVf4xHNJ3PuWH9
FZzCYQgnqI+YaLPXAEV7dJE9ydMpuSV5k8YyZuNJG5bl6fPFPfx7AwwscPSnijPq
uLOE+RIU4rtVhGaUVlHVc5EFzPXEwpD8AKSZUwverIj7TciKpD5HYhyHvByoLUjz
8AuYB405kjxfsWHY06MZLaX8MSzY+CahjPzYumADcAEdZF4Se6D33MQBSpI2XswM
a4zzy14scQF/ZKxwwk0IgdXO6qYMrv07nykR0vzVpwWovZDjmvjhZogJo2dxHyWX
kl6AJNUFNort1/Qi9NTHnn+onZ+Mcmz1qxKPq0w4prNU2RJXCRfY2X5UN8v69zMo
J3ppC9/9DvEuTAjGOK1I7dsNE62I8jGDOwuixYHsYCmCTWMbDklayNdc3yAz2Ex7
vIGmXDbf0echOM+ZNSOni4daNd7FS+C0jfXi9/8usFfSDxgPYnb/4h5DlLUNvWuL
3NNQ9ATr4+nUXRJTTe3f5XOslXfz3+bUqbyJ9E9c/Qrb9e7vRxRuOBmQMMN8fIC/
DuuU8sy2BAo76WMiAU5iehpDbgvgYDDb8dDuv6XFvMVuCOhbvDNgdk0Ikxfn64sE
L74YrrtIALT5bL8fP3PhNWRfSgrYqDU06WstO0oS+6fWzgELYg/FMVnazlNgbX3S
O0B/b31cittOcy1WjkleJevJ1YivPEF+TVdNI/eQTpUVJuFwV2rIjUKd4fQhoQT3
YVbE5/Md1jDAiwXAFdKNVS0KSGIkH1r/ODaSrMqXd6qy6TS6Ryimf0EIG1nXITSo
lFIIKpqT2LgOPwc8/dz/bFP0F+uox+mJB/m4VTZVwelhP5HNNpItlDECAw2YcfBI
ON/+mckhr4Usj4WCO2y29b/7f5k1CudEsd+1NJCQ+Wdhawn4FmH8IZ8s29aPHQl6
ORJWKTbHli1I0d+rRvcYDJAtXZ3JGfZIThpO4P98sRdxppeWD8067NN4lndIbDsy
nWS/k+kqlFFwbX6TDPQAb9kWP61lI+RrdeXfuBSXFCPjZSbSzMvbRlrvqY8e8uor
vqUqtVVo41nM+DQRZAuhIxftuWS72SNdq5j5MYosUCS6eFUhhCKk3N+LhXHIQncs
FHAM4nby6tSbfUgJGbyWJsaQB0ZFqUWbzP47ZrOTpcJeNkAE2PiI1piD5ZsD5dAG
4gshWuuYDnv2/Lqq5a3BU2sYnJOEltG9kbnI9o0OZ2ECm2pcGKUjydv46uHs8pAS
ft29D2JAE4oipfm19zYIDyeBmoushdON+CZKYlaLgeoNvFoe64fl4epE2wsF6Q4d
pFtwZqh7ph+WjlTvU0pTk26KKUDv9A+VoBAKTPUADvdepCuLVdBntmaddwewVWKc
BVlOyU/LflikQ81TXBTxm+ZRCzfL0QoyHDjL9GT/C41vmKt8+weE0Bjhk5/0PEhT
uqSfqkCO7+JvDkDKujN4HpJ8icZ/Qk8shFTHhyAgLaRaE+XkabkwelP6DrBxXbVk
5e4cIA+S6Q8VGYeBtRGTqrjQDotS1/BMYXoayTM6PKxWYEBv1yzQevvqUkQAvQHH
L2i5elqt1kQhwKQX5Gt6zUVVTkFtNtyLQ34SH5XBzB5nrEWrErJkP8xmmPq5Zkaq
wHiTa/0t16cRrYCvW+8D3tMazjJesYDFfJY9LdMbIsV5UqQpGxq4sDDFh4S8lmgZ
xW2zpNzfpRHgY5FGLuGVDKeP/xB6tnQ0KCehiHlBgMbl01Z6WId6Pei7ifT3kQ1L
OaUuxKg23Q/2zy5kU3oy2wttFrQRyJgEYtgu7cHkesnQX37CRC1ZiNLyBnp90nil
tSnYnWAXkYElm7FdwnCMsdnxxxPPMjaycu89+L9JabrmIeZ0KyvGmYUrYQCNVCtx
dPXHOFqQpo+fM0MpTHVs5mVt4upT0z29upPmoDSraDmE+Wud573Fb6wTXgWzdP7R
3OmNdHmYFZfHz88ovAPSq2uSASz0vvrVRNWILDSl8GlKUB4bmv2YXrxcjTrRTNfl
Tp9Bq1psKOcC8HXcuGVOQ54+8GMPoVaynR1xim/saLJ0y3wXuUbCfCbJmVcidu+m
Xk60/UXL2O0Iw+/CcZslFyTUGhuxlWO+OSVl97JqRMexK9nJq8bc4BP/JLAde6xr
YHspG3iYUBhBm0R1eDW3IS8WzuSkd7jEaoXaUzS6EoyPNzpxB/R3GjKcqxXuT2Wa
vDBuZuGI5nEo4izHRZL/blG6IkcP177l2VgaCDyfBUH0S/EeKbx7mX/7zMmp+kAY
M+xiUd9icyS5hG3IrJx9V7Inrfx5wL+k/tnMnLMP+XLB1bXZc1nHFd8Tyx6Q3/U4
0zv/DhbKE/rPX8q2yTuy4MXE4iAp+nfAPIwuAkxQrr0+OrqAfjGrtjwTSIrwFkPp
WBikD4XJ4Fawp0eTX6q7hHhS7PJBeBGmcOSFvAJrgKKNKp+KMkPlokuWGxGHwl3k
1h7t/wvfPO7a6JFLvYa59T45CKE2OcvaWbfxh6nBeAb8Ww7gpAHBjkLop+02Vlfq
RdRIB7dhtpVYA9uVX+eaEcE1pyKS0BRC3fvAW3kIJ6tdepKc++4k0+fQj0gT2ER8
52N99nSxuhYJFpRy6HQX7pk0wCQxrOFdLQtjK40k+vAL/jHUZknC4zkYEuzrQzTw
syhEk6TYC20nS4/Y1UHy62oGuPgsbB3GBNUQxlh3KrSlmtB77D4K6x9J4nZMz8cI
oH2rOnG6krER8h7GSAFDNjrm/9dMtpaMuGM/aXvdB/GJJBeWHvL3I4BnFEJahuIs
75jmBsBmFBgJ0h5+glpn82r4gmIMgfeV76q0EqUZOl7eWxcqJ4MzHEBsc7ppJQdi
8uDpSpaVSE6HpubSU7sG2jM2HgIC9/tT4HgCEzYpabU8PG7jmkziusK925mR+/yi
my/BpwEIstUe7EcrmQLbprxNi/xVjGTrduRax8Bgl9wrhojRpItPQrXOrB9m50Nr
Rx4UtgAFtW1G9j8479AfODzydQEFyLcBaZk4EM2YDATblLJGWPjhCmRdvz67n224
w3EIgArKBhfyA6LQFG+ATmTXqOMaT1RL1ovvfaEeXzED2LvJyTaBR+xZJXnkLvZB
/O2TzTw5dWJVphLL75BR2vwmEF0v08boPyt8SEZoPVep/jKUOybMG6RuQOLCCyrY
bRkWFi5zMoG55rUt8/GOkEKgSTr/kUarqedvcXKj3/QX7LAymJQ32hhwIPl256A7
j7U9kJbeeXD23hrD6d9wRRVxi7eKpv2mld5rAbGEFjeQhtrFM1lDZ8oRdNUpLszz
QLWMlyHXYSw6gl4k7Ni9TdXUtvDqA1w1BuuJGeiSq2RGFLOkUyrOyCQxEZ89QfKI
IVyQCmLvNU31VqQ8W37lGj2iH9DVjRECiymzjgpM4cJVc0nLlGTewl/Lrq7LCUUJ
5J4v3DIwx0PNDQTUF9QkaRMpcEgoGI7l6bpbbaSe5hvUA5W2TDjQX7HgGqmbDnB2
+ZcR2IgZvzoBrHa76vQrEfNnfs4MRkG+58ohy3IjclBwLAiA2VfQU/gFpag++FU/
FWiiyIXMvuqHZzyTodeVZ6fWSbEQ/ksZoQBVpjI/NlMZoOtEQVw6zVwKfQG3wdkA
j8ZWJn36jOdU+DcejgtYmJKO3B7Wj7tgENHlobUL1ggx/8o1ugxZAiN5gPYFmv+s
IctrYSklC+jx1ubzcYQMy12YT6BM+vA8fzvsf/RRapPSw7Be3CyFPzg5vZCcv1Ra
NzDXUGZ9MTUrMwV9U98zPz7l8D7nsLaoAwTYA6T0yJ2DiVou3q3cRw292KMwMPcQ
Z4usn4vp8YnpwoqLR41TGtnO5ijYLdJ0ebiS3lznbG+V1Csh+V1QSxLub30DrDMy
gj7+F7Xj6WUDBaF3t7s7xOya5HQCSmsLOagxxbTKzbUF8J7QhJc+Zjnb3jnHFAeX
dNbqjH6+DkZDbkL3QdSAvAb/oajZhSx2Xt3VCCzo9Rt4VLp1xZagybq1NmcFRlRd
IFI0rqXCAAbmVyLubGny/VdqmiEGLW3bxXwA4jqW8kBnr7EnMD+2vNj9BWhoWlOW
Sk56jW47rhljV2P13W5EnuujPN15E/1LfeKj/X9TLpvNgRo6ssHeHkgKtT9+UR6W
xmpVk0N1c71a3U9G4NWQKB/afEI8a9SK97u8t0vu5w6d4FTd0HQlgnrohq7pAwB0
ZQ3bYcG3ic2WmHBv0hu9qMmfnQ4/ryvPjOLJyCtL0wEbK4yVYBza1L5dmNaKc6uI
xxvT69AC+L/j7TIxnCbraOqGDhRSwE/LCFYhJbAKzfo93lvbVFeYv3BWNX3/YfjV
A+bLtZ07M8gi0G1hq07iueCdf3X2eDlN41DyYUbfuN0T3w4p08XZ7yHLpuZrOjQc
NK3EcqZs3xAPqgATNXlxktfBnN66WFdf0RfoOYWdDT8ksM7Xw+NVFyPpE7CGxjEV
0MhOEaN08sNOG7am46aQKRmUyIcArpGeUAxucXDbUkxcvULWPXZIYOcGQd4QxgsO
UnjO2FQ5FiJ9yCcWBacusPE3si/APyAXkBQ9IXWkDFtRu1uARygW+iIhvMbUhsJU
UHVVmymUEmO2vc3vSDohZQQr5hxMpcsLvucQBscGVRDr8h7K+uso6h6k7vjcnXnE
Lg2S/4JUFgrnRzDic4X26F/7PKFpQFyazu3uwKezJQ0PBv67vU0f8b+6WtrWzjUo
zbdUdFlvKfZ17jGJzgjCdzxzeSQerML4TPlUGs5u9KZNg+cHYbQ2sjk+Apy0qI/q
7GSzd0lPU2zX/yfnJYSzId9TD9lTMuh6bMsWeygFAaEk/irz2yA8i3GgeT6vhAxI
lBXaPh7bOk6ISId9cKiTEOuodGOIskBxdk5091uas4qIlrJP+w3HSpVpP6+R0IBu
GWverS2SLv/PTZPQkqPLL/2ARU8fAfZFVsVKeknXEetR06a5iR7DTZTGkdQ09fcN
Np/OT4Qz+LMewtEwiBOH9iX+XF4OblcpZV175mUSneUCbahK0doQLtEisNPOnIBQ
lieyc5affMKlCr9CL47/7MY0VbfJIYItgOlQSKZLydo8Ne9Sg6i4LpAoYexiNzMZ
KVCeW87Q18bPZqwzOxBEtJqCsPisJEfP+BcJNrA+Q1Y/FqtXjqEpGSaciuRtY2PE
wWk59q8dsHCcdo3q5Xrq656QCUrtKO8Pcg2VcOTE53FEMqL6HIgjDBm1fz3PRpfa
hB42R5/bMvFyWdU5IdBPFnqR5wmsmBmlPxsPhc8zGrWaVVo1o8Cl2E2neVndyole
+fqYBsuUPyzRmYrfGw6VAtqwfBHrIqsaSvSqY/IPo7bzmAj9duQS0LSdTk9/oI6j
5+WX1cHmwF6hnrZuOZ+qktFW7J9yE0B3gwvHVi0B5zvyhDBwbClfURqUVbN71T8u
Hq+B6gOAPjajimoUEmKLpXYbLIk/+6ADoEgDtCG/DZVLLHUwCjoi9cmRj0CT9S7B
xd3w3fi/8l7a99SYJAP9XYidLTB84GVdl/qLsAbDVobrI0U7UHjGUX12fcbZuxlx
rVvW1REBIbsusE2wwcGLgzyjZnvTqWqSkUV0n7dW1EfqrvrFcyhSvoKiPjbVfBC8
C4/cbPt1R3z0MdwPwwMrV9emISW9P4XgSJE4IzBZTCnDC6D2XUYd42Y1QfWMr+ab
NrV401BN3/7Yw7jWdYYOpdvl1/2qAm2WxHc3lSNSX/EAslWFxm2lC3fnfB/qALd1
03yle7weUV2MRqnTnciZIX5VnmA/lqVsihw8sl9GJgU5lwC1iuS5R9EruPpd+Qt1
o1xInSizPg96h70jZ2wM/U32GGskuaknikfhNinsrpnptOnEBIsHQlHSsinLXYuR
2nrZBHOvqpNl/Kd1X+0OKnuxHMsGCG7FZFksUKqgvqMKwzvakeXLb65iqYtfIUYg
zzbAphfP757l0SjDASPg+U8/i5wkOmAv5hZ0QEqIA+CyeVW01cfaWlMRIg9BsNLI
rlrj9s6pcNbAPdSgHWORK38N0cXcFHBu41HoQ15MJIpallXfJERsEXjVALbS8hMZ
AoDb3KqfwV4M5QzlU5a+M5/rkxjPF8BvuVAp6615aUZcdxb1rx36FRNEKw5KjkoQ
POqyianlKw5xpvTsIYGmn2R1H20FcpK4aZhEp7ODLTzEmSLvxactSjcuSJC3kYA5
8NnR8PMPxR/JpAEpDu6C7Y64LLjLJWepGt0RAXjVEpBl+X7/PoV8/1iwOK/kmYWd
7g2D6roqBmxukERp1xJTmRpmtcfS7B9ihvNjA7Q5JuBwL3jP0S4Unp7h7J9Ybg5B
x7d2yQovKOWQpNtULSewH4r8K6+x+WWiEPD6roIL57AU+oWJhlchQhgWKkqzsS0H
UD7/YK/exgKEE+lrvAPoiF5qBoEK9akruRR7KRncfnKfmov7LQEjVAEpbQSfs29t
5+7yWdGjlXIipKWpYgoiGGnJvQn/RWxSiQnLhvpK1/3rSjrsluaW1NEikiPY/1HQ
6OB1QD2ZLmJPg8GQYqyDffEfti+IFCFbjiIUdUeL2uVb5ljhtmqzbZquKtXyzex5
ujLz42126XtU6PKLw6PAZFpSI7PDQDOzafF7zEab/4yNBc9tEQj9UPO3hjUa0AVQ
NJSNOCNB0OdDzbUIsIFkdx4LnBM0mzas+t9XmoUCwc+Oung/5x2iW2tZQcE5vuqP
sSL8A8Ah/wDZlz+Ig2BohKgnUdN3Hu3qpBIYXmLCoSnlfRXXnlga0U2knXa9xEhz
ce1ddwJfzM9DDJL2upNuw9mB/U/X55Cli0QKhoBkhV+ZwKIstaIJmtkwfizmd68t
X1/c8LsY2scevHw4z4bbhoLFlwnW9pAqCUQJCKg8ZkUVv+XVEQeZadcG9log+J3z
/23dupgBuOGV8rQHRWHfVqP8etZBiwa0nMjCTQlpyVnvXMJUnzkjtiyiYcydaSVl
B4at+5/VuvUTixLs91WvsJ7z8SrFr5XEnkEPsvKlKRA7ewbHIVTXWikskoGKhD/1
Hn2E9xNxdGUohsV9Dv8z5i4gFg6GlX/B7Ot5/PxeJ1FB01Wl79LJ3nVElfTxIZj8
Sg5UDzrTr627XSyMt0xZD4K3SmHyGP4/j1+tGvQwvUKG+EKQpfQ2gCWSd9Izf7jM
PbePHMO5bT6q1K7KCybGFlxGbD+yWjpPAe1CUo0cBwm35FXvzdEK2KJdR6FiFguy
KEGWC0riWQUNkddKjCFP9Ankn4uFca3LBpnVNY7QtOQTOxQQya7pNp+nfE126nFK
6pByrjkhZCiEbHsyuYLBmAUncoSh/Ya3v0Or3Ql4K4yA21nif7w8UTZdX60ZRs4G
WKgVG9uHHrFejCS7FAvwGEcNmypaasPoluVM4G3e83HOeqsMjzcRX5D1iz0P2B25
J614P7bgeVoPIOHE+Ulz7Qk291/eIabhEa5T901xTuvstlqU48E8BG5dHrCCslxf
9/6F6eOEsKZqRcyHPZ+0yj5VW1zkBfGyWVn0rnNVhFULFCaicWbsllaOS0CxzuXo
/GHe3shkrOmdHTGIUnfH9FgEwk0YLK5UBvHfcGsSzbCG3UUy+LoLZsNgtqXepYWM
ys7M5Jm7DpmTExPhSBm1okV/aRcIREXn6SVgXIvQMabi+M8zZGJ56LzdYYSk3g9o
BFIZ1iFi03uFIyyymHbH7YBkCWMo1wr/hWeD9dkkj8KcweuovcY7qtEGFyaLKjrg
hn/minVLUXpNCj/jwr+LSKkPxG0EPguXi+nbclDx2Oab/iQZ2iEho2Fnd610Ca+/
yV+3HLGQ4ReKTVyDqjTi+GSlKtWiCaylgtMcY/wH/aV7dhHSaGFwBaVMep/yJQvp
vDWSVMY18T5POR65ziII3FHfEJjvTZbUZkBe4K6veOjRDGhzdDFMPvvptD09pnJ5
kQFMEtXbrk90813iDrH+OfF7wqEuF5gzYl0uPh6/vZCgn3WbcXlgkwZC9KooGope
TIczun/xMkxZojIFJ0jva5hk/hyaIINpaDhMO5sRyrSualDLmWV7ZbSoOLslPazC
wUJsgbXsCUsRhD5J7QDrZqKkPz77TJ9xg+6rpr28IvBxbEfQaWd6bCC+syYQQnjf
mF84dIJTvsFGEeUSO8QgQjnCoyRFiqYnjo3cyWGUTHxT6+ZhNX8FQ44m8jdC4SLu
3dmTKVRXbOh9InmNF319R/Fh34LjHCoQF4KbeQVvctckKxFGuXRUdRrLI4YP7vlM
kKcTP+mUG8wXUMXFwYwa9vSHcTNS5VB+4m9RwRzKYWb/sAcxeEcJ07ARtirZmdlH
uTwAF620qH3i19QMDuR/f2mjVxEgtcP23TtM+iZ8RWiMPJ25/DfIotGETURo+CCF
6f2o/hgVeqZ2Aw4Maq+bnabrqsDnh2l30dZztSfmxnAlQAQ8tDbck2hE4Z/0Eoog
d8FJuRD1dJ46Q4fPfXToEh3dRuU1sh9+HpFz/AxUUAXE6n0b6HVlpd2gGqH7v58m
YgvZnHetI7vzwk7Y6vKtXouDSKOm1TNM8PR1nw6s4qRCjArbASRMgziHVQYGjjH6
41mk8IkcfrO+8yn3I0ytdRSs5mt+/jtQkHwAB6X/YI/xbS8vic+mCAtCKoTFglbV
aB/3gT5a46aniH7zFk9stu6ACm/q0xf2N92z+ALYheEkvr7sL53rFAb1dnd7UcJ+
1OwDOPEmahQVpll936ys7bIIBHujFw8ONQe8tl8qmec3QD5PHC9NCaeV3Iseg65G
uP0gVo5rF6uKtkV9WLQ829tH+goRzI2Glu4DBCLwUd/w9EOUQAYeYb6gms+GWQLp
W+le7uvLs/pcguSh0B7itRpD1CkP9b1a7QuMAxcal+KJRv1Vx6aGwq90T9Lnogp4
fXBdhvlNUufvGbCeQAlzvHwwWAN3O9wHCU6JLbN0l+pfpxALb0B2ByPyJ6nsGC/d
mn+TFLVpSPwhIj3NKdNtXOOT+pHJ24kafpHD+GhC1P1GBopZUtRtpTqaDy0RuhQp
2fVZGTVrthxV0Z+A5enXeDmNyIxLGJktNMe7PUxMamRbr17iIpanBzvEd/c+UTNS
u9rJzSAnmdKvLVwt20JxxVtS12uR6VvTkatHGQzwOcgo09CCGcfBPuRBWLwCa5rP
NZfPChadjq6tJNZjWatdYzLMSXn97SC53EVXfcT/41qMLoFOzPvv/RS1rVNQfcdl
WOl8/vWwj9xXjPkU7u2Ik3dn79L4oNtRU2Gh23os6e7VYB3Qk7zO4APfDSYuAamA
fm2QwC7xkVX3IG1kHd9YJLAFJNq/NygAYcSKbyjtxfJwPOjmP1IFfrqzC8XGEXYW
ReewKXWlHVdrgBKnoHzykUprVk31IdtKBGxHx/aB7Lag9PY7MAfm0kn7B72uqIqJ
KisEzCS2e8iwZ9gGPZnUz7wzMMLFA4q9yCCxgbmjpPD0wjnyLyyVeqNd+e5E1v9I
2dBoPMCLGMR8o1mAqML1MXMYuXcq3DXzC9x5KmfeRPMTzDD9knED1yhd9fKe874r
DSuQ1vINPI4YZJe4tI6O3LaWaJAWveKzcOsGgZl3W/WKM106fjyWLKQ0gphwm+hF
Kwdxr/lSukUH2i68XQFMJdMogY+VSUzezVmCvljFX51D71jZBFu3IolFaEaVGyVf
TckAuEwR3UrR0/iwm294UEnch3dO/dhuTkLx7DN1ZCGWhvjHH8AKKra/1ydDH3Qt
hVlBayM+j22UIwjdIALGNNakKmLN0tisknB9hv7fiHz5Rqj5PandKsERvJEJFjys
9TvXNAaR5UfwovCW8wGN+P64mkkvB2tQIX7ItmgcQvdc4jLhfMNPcSgIC8MmqWO7
+89g176zi+YoyrJPtd96mxe9lhbUGTgne+2gvWpeLKk/7xYhZIiMF1W1mpDX1EgS
yG9K7Dpqn4lxOLXwyOCVaZHPXvVmKja73PJBfsiys7KIxyYv3m2JDhnYw8WZpv2F
9XvTVq83ZUm5xzNj27OJ/dXVosdXITp8JkL2MdRHNFKX/7KKQ2rWF9Jnf/D4raZY
+dtWuRFveOFYpxfcxvX3Xgn4NBnfHTfQn42ZaozxsXq8MyOr6j++nuVpVGQBiY24
Cz1vbhY96TJ+IPCjRByRVnen1sXGhH8iL8i1b3n32sc+usbXgm4GcqsmUDItmDoj
Wm8P5XpabtxW5RQnAE7HoFdr6NFqjgAstrxzzwZUX9fzkcUuPQcfpWzz1SJIifOH
4Wo12Sy8t+olSO3c8SykVZ6kAsZU1N+zMBjucsp+xjXpJfPc9CKLUPlfj3XVvJEt
/iaN1RlRraKP1QcdKC99cXkIrh7kKHxUXAayy2AxqW6QyWiSu0F30U0zInKFWGev
vhNCry45cjdOPkSCVc3L30k/cp7N6rggukoDvhyU9uj8P2Fu3ZABRa3AQ/9Jnq7I
m8Pa0k6RJCQ7HUpUON9Lh0e/GNgzrLlQ3maWnHWj8QakIyovxvs+Ej4TjHI2VS0I
9p1kBzaB4JOwZUOsEuGQpXtVgk6w1/Dyz9L0Ku2xaxddVpru+kEkdB7vLJS0L9Yg
+g8Yv9F4te8dSuH3mmzMqWlm2D8vTsV27Tjs3QKOAqGmKmVVPswBBmgOXqm4rQ/4
mdMv9pgurSEa3F3QSJ81mI23eqUYofks19RYYAnIyASsp9FZ5lqsaH2DM5/w++9h
beDq/v6Xhwn19jshwyzd/CDVSDM42m+z9KC+Yb7EZ7od/vzKu1+hUUaLR/SROzTM
1a+cnjxSI/aHxd64ugOFgyrJOs/bHuQODnlqC5G5X7QLCjvJuXeY/23e9AA4Wusp
RHo3EWRfbY1UL4sMrYqEE141M66WKUkOIIg2HAHWieQ+4Sg7RwCBfXnW7db/Ip1y
+Jr8D2xU8l+9l1dU7+F8i9FNBzoWRnMQ5ZJDFLhA7A5A5ZQYi70ML81O2hs6qd9T
3AMZ3hIR4vJwFFR5ERs5LuoRwCUePRYPjfrVlDNzi1nyGbR/bQyz7VX26b9mjWpZ
G9/k7exaM683JAT5qaL3sVGRIzaGvjCpEjF8UBzkNvp0dQo3IRvkvCaAE40zBFnP
9JAQZTwb9OyDyx9Q1SBNmhD4ig6sTQjXL4QqCtsK8QsoASOgaeVrztwYZJsMn3tf
vA8xO6ByNzxzeD8oo8B8SiETdaswZEHzZ5ASNitQXolsAWbPyWVd9nugQM7PKnsf
QEFhkqDK4aysCsPvPQfFnxZFCOAJKKuJ+mhqH9CLx+i9UYTtLizCLE1hBqAJd+PM
8A1iB54fvHZGBTzicAeG/6coNKvYX8oajSHQ6F6OsiF25QaQCmVLmhVl11R6QA0L
27IWBZhNCn+PbrIK9NcPz1//0c8/LPevzUUgg7tjbou6be4rE2a+UnGSQMJcyg11
buMuCO5aClhyGCM6+ip8tEvlzWr01a80zq9K9X89ZoItf9ISaSfzXEuycwpjG/Xs
InbPDkJm0P4GB92WRfQ9K+OSQdKW0wzTAOme/QGCGzaDpOulHAhdveeikdktRAID
aJ6iKQ2XqQ9rzZxgkApJf2MBy8OMgf0pbSrysaq64daCcVXNNC17TnEqmgIrY//Z
grF61W9bBMVD1QSp1TbZ7Oet54wSY+S23SEc7S/mibTEXpM0EveRWw2D+E/nq/Zq
sBEM0/3AhyWVsH9OOahV43yRouTB91WkkY5uSJEBxtzrMqnVLv65che7SFionMxh
I79Ja9GNra8/tEHeyY9YZgL+rnU6ABrKsPQiROUYW8LMlLZXsZNA1TQzczq2yOci
eDRbLlYIirFyR9dyN5xMGZWPH8F5fyO4FyAVya7HA+6KUEMuBrs1jYtSSTko2TpJ
Roy8pPH4D+dDF/iuxNtfkr2c8TuugeL5WmnXpilIwStm3xipMaCrRx0MwR1tavVd
1XxcTTB1LHo1Cgr7kWf6BWyi0CHaxkBV9bH9IzGUF5OXFmXowAwxeMWJqkBcfhSE
PeXPa/MI4A2Bz91u8u600kS/0B1FjXqzgSEyjcFDjFymbOdlzOlVygXXIC97DWFl
ThwIPvhibFiEGf7ne6CVanRjHIdwnM7ZxUbm9oehg03Jvl+r3WdrlnA+6eJIc655
W1cWhkBNOqHOSn96MdLDCUIYS0yvt1us8uu+W3REQefLsb5LW3PjYnhDYXDJMFEX
J7Yp/Ed+A+5Bq24tYZVu8Y9XfqIMQ4alKh8GB4aVGFbSw0tmNtYNSeoIyecB+Oyq
PHAblAW7RZ0ISCykcDGg/4JXgfRBj5RDUDtvMnMxKrMiJHfONnHFcmMMWEViWO7y
9gv62xvCUZx3/4pAIcnX95MN57cWeQzpI+JQKJngYwcjXrax291gBFrF4PVpYZUV
hnSPc8yna08sV9u4JJEfsn5N/A4WFhyfUgW0QEMWgRVzmAZ0xV4Jgt79f5OTpEtN
jp9qPC76D4Kjnu4UIxG0MtePARlG8NAB5ks/EqNFIHDk7tGmSJ6ClAQHqEs3T5d0
hhhZuAUOo+ujdEHqCZO1M2gcZImO1hpyDrpvJyBPxueI3YtgzC++DNnlaQS6DqLI
9/N/15wzF4cSQfALtPXb/gkLWDaDNaWxUcJ6DKmdypRhfdC9/JIA8g+UoZqU1r0u
QziAAxf7H/I0G011jESnGJJ4nvx3p+/e+K/6XJRtKZVNO1xMB8YZ/S/OTs37UtoS
l4iryn2i8ntTWvVB7hVCGrFGUBg0gcaFRQMm8AaWAYmU5gF9rL48UJTXoNlKJEXu
9jV6wlVAhlxIAc+AAKgUBCdHPRSuHMme7mKAzyWh3e8ckjk1LI6lZTkER0chzXRm
jScnfnY6ZThrmI2edxleKv5iOewYF6Kp+wWTCe90ZizVFCuig4wPBOvz6hZ2NxNG
dyW1Hv4XY4Ft1GaUDC8g6z0nflFKQ44p6xDQhN2cOnvqDKuRDeUDwuZoltoW6Ujm
F0kn3vJWtrSqsHHVFjH/C1kiVWtPvUk0+nDkHJUUyz8Jgxy0sddY+eTWqUXTG1aI
fs4r9/SLYRqhrAgI0NZ5ngOWytukeFZeNJw1xpYpox7yRg1ZgFE1n2k0DpDh0T4a
YmfktXg2vxY/0nGPJwm6TgcS10j14hJtEjunGVZoU0A07Voh1qH6mEPhmwHTafM4
zBvJoYHRAHKTLk5M3XVJV7YmlVTJjdC8DV0JK82J1jDv55VSicMOz4fwEbh3O0ZW
Hvxgb94xtXVokd7MSLWB0BGjYs1xPJ0NUnRLOQxd1r2dTPGtRRCdWGlZzNZ/3uSw
rjyLuUm2yfv8CXND+VEZS1wd/9O5M7liEMKITroqnPKIqV4qxfOTlp2AanrJBim3
giwk6t94KzIhhphM2xZOSE2Am7YruHkWp1+D8BwwPPFA9AUldOlExcfekx1tQaOC
/qcaO+9IaBOX7BkqYPm66D+SYsNuJXPC8iIyX/eq9XGHTzLAmSIVe1mrylYKQqQV
lhjY+eamH1KIzCm+ciZNqvuCvYdUfKAoVXPzcYTod96XaQxxfI0ry1E0pkBuUcFb
GkvG+BtgI8jTtxh//Y8676EqU8b7HXPEF9nbDDuvwdZXL9Gc5EvosEoCiBSZItF4
6NFw7PiN9gZNXg/PPmu6AOQX/1zN8GaUsy/dUxx0j2cNoSMuqW6kIlevpNhc7Xvw
kGMOlH9oHRvjuhn90ddtmWxoJh7ToocH2SzRptz89OM71JXu4WCc2M+DJXD1wnqd
Dfds8FzYeIsyDhIeszAkhfFgGA6nx4A0L6Uq5F7HJUvMzZevv52nvJiHpG+MQ0BH
qUrd42cKKWmUpXJcRDfGcZJa3fKUNTrpw4QNCLeAYNfiHaWDI7C7vuezG9pNlwo2
69tsB79vSTWzlSmp3OUQ3KOzMMNP/GntgyLzBQHZaK8p+eeGbzA+02/eVpWEAjJ1
Q+4TYMFpilA1yqwBR0/zggUI2uduqTzZsl6ajW7zz9P8yOwZZxnpIoQKY/Y2ZKJW
r/f/XOBYlw78aVcr9F+0DiLblR/0c4UeaLi8AtX1IwvDQ8T/G07ls/5GEIyyIPGl
nc8L5fjxgFI7wAkzaYgDyY3cPdbI01QKpIOLwzqDP7ui98tUcqPW8k/ydSSvVnkO
E6cAn5lAKN017zh+NEngptcLyUhFDEkVYigFNhFFZtxxATGBPS/IQB52hiA0zXLH
z+dsB+AO00a8UlRlTk+YXSmUEfTJy6qzO2JOwMNPt5IWhgQy5uyM4Vo7Ti7lorHg
WLZrrkBqmQyjeModhcFgBQZdu2GOLqsje3wKuIiGkNkMcsKXIDtJQhDRqxXC3ihs
fnHE4UD03nXvQ/AyQ+sCqAoNN+eMPO5oCu87/C7sCzGkBkFDoJUS2TV5wG9QYZNj
SZrW4/hEfvB3Dcufpq/RYbywegdApyrguY3Q7Z4lKKjUgayHADPb0hMnHSGUbWZs
cQW9z5serTlnJ1ud9ZUwhPluiS7he0wsj5jRzYFWG05helL/WfyKBzYUm90w8oRV
rdspcZGXhvgtCywuR7WwCUva2j2dgjfChUJbDl+nBEUfpQ4cYQc8QCR0ITtuUIX+
/J50wqoO7RjxNFS76OJHoJ7Bx2R+FJNLLucYXajcZ6X/I7j03JaYfouyqjcvSlqB
jlRmcWFG5sNds6KE0vDM683BDIysJDz7Dshb3aApzVKEyx49e2Sfssg88yLZddZW
6u8oJxqTyW3sFcNjF+FYL1Yqs0dgdYmbbVCR3p6qudDTOM50JrzEaaxqj3OIKojS
JVp/6B3r4+ezFpKvKUGQdOsOels2jRfkiUrpo1TwRMotUlz+qpq8nM/aXKIBbsCN
4ZZryQLgiQdreWWCPKX5jyhWAkeDHYJyszf/9QjGKfF9X06LpevSqkXAoTt3/vyW
tYoZc03Q+hIbkDSjum46hqclX8uQ9IKGCk/ztD2Wu2hCSrxl8FLhmgykIdT/OWtV
1KfRTtl9MGaW+YISuO1gItJs08xTwPnYQPPA7w+6/M2yQkR3wmUZr0FkwjW3ofFk
bDrR1UIzB0zQWvBSq/DyRoPZMjTAysZX1oPOMJWIuU5vfWYFKoUBDG1VWmZBMdeI
GftHuNogXU4h8NxnaO+DLGWN2wXA49upp3lj2fTb0Ghc5JS7rZEAfngxufxXfvX8
rqAllv/YfGxH0Doe+otq9Z6kDPCNfScDG99xE8J4szoodaTICb7xbJLq6qm8VdY0
KAzUztHwC61bsBs4WYmOvwrG0oTWqVuIA1w/jibNWelLKLIG7tylZQP2LMzsnRik
8AKw/wOgjNtqsp8RWR5aYUyKRExXEwxoPc+YebMUS44TKqPSe33eeG+ST2qvmNiR
c6QseQzff7dVrQFnorZ1wO7Pjazsx5y6QYvKualQ/XJaciQML/DiahqdYLKvwhjj
j+uKDiXdeqznJYe1qktr1pMh/n3cPXdLjlATX9DtIG8yBdmnJz9WlLnwnGu38VUd
CLF9UwhRD7kfz2UAIM1+iBN2hbhtb5S9rNW68+Omd5T1tTsp/JxomY6CC2U2HjQ9
SSnasarYL4QAeLkrTXypNqSb5ey5Or66WrkdtEQJfCmEky2K9G8n/R+HVjsdl58I
KWjbQyUh4A/FZHPdw8wI97V6l3DJgEIFRXkmnuaj1TpNVl7/XGrG7Vr9HhNucscj
rS729JSRvJ0QcFmOMsjl1nbNDXatLBhqWQTF9lbyRDmhtqoFr3EuHEEkKJJ1kHqt
JGr4uA8vTDFMOh66ox1Ve+Y0ycrGS+L2idLBc3NnLMBe0vIbAmvo3gIdNAFpf4wH
3PMjQ56Wh6QuyvSbAlaxG3tByHeXKL4O0T/VX9sNumhup0gPNOC0e4qoN1WhHwHy
tyiD3mLZc5WuUd7qdG4nhluULSY/PVzL+Wt8PSwsMIKd5s7o8aW5C7n7p9LWskyX
9F6lRs4aqa5cUOqu9wULI+KM0pKL3gTC0tJXrbOYHBr+KXuP4Zbo0soJ/X8ZGWGH
BDrgGAcFe6ajT4T/C4BuMQZ1vdcj7q9dbFSef17KYD8Lmzi8hbktNqnjhbJ8MSWm
S/45L9UtAgMG4mI0Pg6IsZhCVd6EP0aYm/pIm4n5lp0CbbneGc5VRkjByK7vbQ8p
kRFOAAHsm2E19Ek9E4ureOC5hWs5ZyhxZMMPVSMcrGuLmADR0cc1zprhaTSyfBHp
42XVNFj8P4ixV85drQL58ruFcytedfcSRpUPvzQS1zx1wJIFKYak9VFmx1xuWKvN
1Qot0568UieP7X6iAmXrwSG3K7+BSagcKrxY6r8yQDHQSavGVadebnwxaghrSPPa
OH5c8ESqYqQ7IPmUDnTp5YZL0EiMpQANf2OtUnpaXbh5odF9sXnrLp8enuOO3lpY
JSSBUF1Yb4s21LqCqoBXGPTIeMkDWPY4qJoiBgi3Gvhb6oJlAQ6Big70+VtNAS04
k1bq4JPjZ97NAdDJDGgqHgliArAlnaYMc44aMumCkTDHWOvLXvwGVN1/+dJkTqPh
ZUsVc1fFbrRnX4rmCMlVV80WW/LRZTl3USWTUtqDEjSbfzD8gashwo7d4IZyQObT
1wtRZkArC8jPC48Xf6laf7Vi1tsrNbq8GsHUdARid2G1dZwXLg241S6Stm2vSLTd
r1SzoJOGfJL7Ot5MhnKqbpD7imZnApHnFOf4Knn5itVXDQC8UBDLktqIcVhGceVX
/gkV0q8ZI7tKgY5oc7ASzmuoGjr4YvqS65OMdrdWwObodjFGyGlw0/KSfdFKW8my
hLLm6tkF/ZoH8CBo1blPYEFfzW2I4OaIIXT5UeVd79aY5INByV/U2wfccL+BvfCA
k6Vaw5BFp2F6DUk4lcENqwbXX7JnisT4ztzZIplp7bkVX4lsiMSuD0N7gUd6hn2R
ReFsH6kncbFkmL78kMqu1qt42kf/qXpd7FgCNgjQCu94DS8Adzbkdy6nYMux+7D4
tbk3fNAFKirmnfpsa0IexBjZHVhVrnPqn8QvkRnfOELD9iih2W0CHTyzcTijavoU
2SirAyuvmdnUp2iVVoLAUs9YeTWEGPzExT+a7s2Na7kr/eJ0o4bQhMC+rAWVc1mq
oA/KXBQ7so3XKofcDrrTEntzVx8o3pIYtsYp0xYe7yBu308i/+PTouFm63wGVe3U
bLIDYTQkYXg3Yp+xn6R+KMTrvApr7v11yB4zhuVReaGrjPbVn3c3Do2FA2CrcRq4
vGJxr4cpmq9fweoNvVbxwb8YJ2Skl5qF/5fH0kEoAFvo4YymZ8d48YYJZv/bEESk
DaomYX/rGhG0PVDTvTg+zdJObonKAlhWdPJZ0YDl/FO2lOU2HUT03G+t9dSK8rhe
fsL2oDYt5IGG+eF8KqjfgUgmWSRw/C1F1xXXgmjMA31quKCjojLMcOm3OauMLKK6
DEhYx6dH4Tkaqx2jIRXlYpYH0jBeYiisiViusnsf7I9k+XVr50YXkC4FPWZJZ5T4
GG2d/Sr2z3+CBroE8pl2KV7iqkCPaix5yAoAIuY59d6GbrSsxR9PNWeJYH7n7/eD
Gq00LmwIpG8syRn39Tpgjv3KiSfBGUX5gKCmOhpWi6aMZn0WbQ9Dme6KgUVMW69c
wrk0R9wgevWZ9EgWrXHIS7q4jdhcvjSBcP+nHr/2f7d8J3moxx8O12/VNd2vOl0n
HATjE1FPO0OXpV6faaJspSDk0fmf2WtEsIW69Aa0DSSzci4mpZACE0w9MehvZWA2
DyvbMg89QT9MkIjAb4n40qL2qAUaxwT92OYhCbzMP5QtOSfSWiwKb326J/bG7jKn
0XwniJ5MgLLxk50aw2f0uEdPCh5MQgpPZ4Lj9mA+5bTo7a0udnVRpYhoWNvpdnH4
1ai9G4GgOAV1ZskWeN8QrmmAdIcW8gXfAQKdf6kesE3860NS4ul1AVMYoAA3IlZZ
NzNB2ZfFcXN5U7Z56OYVOsjPBY072jHxJbwxM28M2nCRrmz9XJKjYqK4EXt7UI25
V2XaqpU0Q4Id1YXXZAM3GPCh/CTzCRE3v/N85DHiihQMMRzjWJn+FarQuXD4B0O3
I8VHRL/oAOFNw+iPHUgO9QN8Vybq3M8eNUQqX3K4clMbfNyHeyEACXMF2rdtDGej
LZXwJfF3NCVsMa2bhIq6/kdRDWIsTvawrIT/uHp9gt+htBvy3Z8cn7xGKQEaL9GG
PbsmeTMsyqeGZ6ihPyNGrCEWTbm4zZzKqHLsd4ECCgOGI6N86Gya0cUvR/SA+GWy
+WscvaYoOtgcfG/QsluS/OeC7e1oJVqRm2dPvZf7vxK+t1Z5w0qwfrPOz2xGRNhu
BAEELlugO4Y85E0lnvELOptNLvus3mDN5qGu6fvom0kJ09ULeK0ouwFjm0L/uBqt
1I40LdhyG/oiw40sYUYHE6tvxndME+m9deG9x0kcL6Rs2lfluGT3HQu/RckJuXM6
loxVyflnP581PilRA2WaTMhpMqvEHIEPvfF4wdKzq7eY/OQmHRJH/3fIGhPOkPEo
awPprEIfEANrdukgu4g9UYxxKSnz/TZut5IcUrjsUom9A3yoDaQ414mfh40Ho31Q
kvEIN6CtxoMHAcyDTA1xECZr0Mb1wFazcZyU4LXjC1htcPDoQu9WUHKL85+xbmUk
s9h8hMF+uk8913Z/12fxI92qkbeGCOTS4MVQGnJ2Lbfgy8E+pZKnRGVvN0pUzpHU
LHLPWIOdpoF8eH1NNBcE0KDnAmrF+1TXBCg5FoZdsfL9IfW04EP/t3Som0JPVgf0
XoFBNXqZMI0nQXm9vc1W0CVPh/yAv1spW1bz9MYHnatkXB0bu4AwO8N71fdQBgL/
uQeD/kbIFdaJUHbLlkfVXZlLUlpw3nUh+DaUQU34n/OQzWKXRn6Nt213uVvxzdfA
wFa0KgV3Q0w8ZUgBs5zRh65il4UoP8/WAENcBqlkmyDw2odAP1n6FU6gy7fyydQn
l234QwK0uVp3ET1AFs/B/blah/eiaBIL62eFqbYZhnJtCO+S1eV0elDqNrm5XXhN
9lzwe/HbT5N4u/Efgc+QuAqW1MB6k5+g/shN+GGlwxrUBnmMDX8qrHXCx3mumzIs
3HgH68XkZ0a/If5s8WCYar5D5N3E7V7FiIOjIeQwWjQf4qFYHyKqfspYdoCh1nMo
WGUsXsDeOqHvOiYOSETIyI+6lbKuY0nws3NWqlV/LSXDIcFiwEhU5UqCB/LK64Hu
D3ij/zDCGJlMcgUUbivmvHjw345Fdd7IxYDJJ4n9O+Ebvb+6KnDvCsiQBx6gMZeg
kjjxLgfNiRtIv0o04FPDpJUoZYLO7QmHdBeJ0j6N5M9lyAf260do+fkzOnJLdQ8Q
hNb/yxWGA+W+XX4i4aPhydrNL7NY19BgkcYzvDJkO7jYDe3/fPgxv1F/CLf1D6yP
trPG6r5fVRNQbPkO/IZGG/J1GZ3zlMMecCfGthYV5jdu6LiE55jIjgyFNHNAgjwY
3VAPaluwBvdtHL079m4mVGadPqjJ957wFBsaZQP7CLzTlopgRsRq63RVReCQhOIH
H+S6bJcPL/deyot1kfv0UC/3QGKBcF7/m0+XBSLhNJmNR+KcCwLNf3KHAGToTbdR
8blmWnQRL9wZR7tQoE7suNiYebzcVRtDFI+uZX8Ua1RB7PyhxmW+3xVc96MgnYfq
ZLO76cjCrgvMn7j6inazub5XdkVdg3GZwqX9EdlRwK5fvaEec+TBpdQ+XomCskyM
EmlK5IhaUcmqHKccIa9iSNHxk/LqqyJK5fia0H0NwKDCfiKlaK/5qkmGp2WNiQQ0
8URlSnaAv3IW1xXqwEoBWmcRUkXKN40AbX/Df83ytH6C/AJHGcKvJ7LPRzuZrOBp
NOFYwtir0aMgnMuzuffNnqbpyoJ6Pi0IuowkOXn4QnuibsP4gZPfqy9ygJehBwx3
ixQb5nFthdtqDI5KF1ECUCHFixB5XhATZotVr8ilC8/gwjBn7ZAhOXRc43pZyjxj
OJ2PeAriL7GcHq5W8ZfbhPalV7DxBdVL7OeWz4/ZGaoj81wtdbIZfKkP4iAidB4S
XNC8t5XNpA2LEAZNT6uHQTj8MBrZUASZfPk5WqZkAH6gj/qIytPDHoceg/s0WhRE
FZWIO4KZe+NjpMCcgeThUx9xMX/+/DXjIAYd/55tT+SlbAgVuCTM56N3+FfYQuzo
efVuiDcoiak8mQKt+V4/hQfcng9w4s/waGBqaEQCtlKa2CLLXudcHSoh1ka4oWwr
o4lJn4iZtT+U0XMHqlFEmN/4CLMndZxYV3GhXzfOdKiay4abXksjDZ4FXpYs6wDq
MZqewJW+NHDdK75bk4olFcTgWsn8Be+BdcqlUlQRswHf7AzWaO1i7iER1F5DJiV1
moSqjwtD6yfp7rofu5hIX97ZSdcOSuslK6VirhQBPiUzQjvsztdjrljwLg/7NrTt
mzz1/ZTjCqfClea9EfiCB/w4gkFP4zLnMc0VXcyXjMC6309qyA88fGoJ5CX+UCUl
xbmjuRzeF/zXeusW2B252rRwTxXVx9mSs5vAvoZPFHrs3GXoq5txXRCfMWEci/jc
6ioP/ysknDZCs5LjJwv+nz58STKIF2Q3wDVmL6a+RovR8B6WBc4U7Qk+k9vKCSGO
pagjpm185Bj0jUMrDCxRo1OOQ4Qyel73sZkPiNeat2252eYRAVCtv7RFWpbmzUwW
OtYq3HooZ6q2gH+H2qqiz742eb9rtTPfB69KnbbLHeOT06gDjZfJBXNlJFFtGI3+
+4t+yLTgO1utX4qBdkqzfGUkQjisF1QeRVZaI3BnA3eMualFL4XtegPU77DMHsv6
YWuuq85GwTtlnAj72KG3s0grUY27H5CwOaGM49r8ygsTqfUJuTqac7TFV6NEIXp7
2PSMJgLtk/sS6t1vRixH+4+/eKSPsx2OWaA+OnF1afOyJK/xAZy6v7YRYeKrQPu3
YGLg++oWf2dUc0oOXXdFUvZcTN19cMatrPw0idFM/HAPlIjeQKNfBdwi0uGm3MnB
wkaKBqVNIjoJGORBVkO7cxHkhA0FzQl9osHwQFdm0k8R84aHDo0LS5BeznQrcm7k
qQzcljqqxbH2Why+3O1iZ2831fUQSWY0C0RtOQmQX43Gtx4XB4zs0BCZ+iXG5rvC
SlRVW2FG+naTuoID8zkC8GkWQOsJ9mMwVeheY7nDvhETkoeSpI1odEV8qFI+vI+P
59U6l1Q4sT7Y9GALlkARB7eHCNilQRofFT1EeS71LHAFwgqJl7buzTFCDM51ydIb
KDavlkk0daabJOLo8z5lM+6NxCu5w11HxtEx8636Skgex/0rqP5B20OTLfTPgvop
VqMhm7cjBipUWIaLXbaGZEAc9ntWpgbW6M5lPiFoMpLDSblUeuInsy8DxBxNp7K4
0+54m+WK+4TL18IWv9HZDJqGcIFkBz7wtnmvPEBT8IAijRij6uFv8843imjv0fyN
wnUup5+oOE9pf7D7reigHoMsmQtwlhr2MBrVLTROaBLZkfBHHs1IJGbbX3GqWRQA
Qu0hCM8TFvbUc00/BA8zSRHpcWbuDRsNajBGI0+nKvDk4u1P/WiN0tRos3B15fi/
hujUDwa/oN2YxoOxfMdIVAYDrCrK4hnOya5/KrrQjs0l+hQYn1W9p5j5UCL6R3BI
nL0hIDSlmk8AxPk9fwVwOPCsXfRULJHUUWj9ujFloL/mq0GPZ6HS4IRDOMkxTqYM
wPI7PpN05AxAEvrIdnbRTnJ1mhYDijjgZE+0sPZYGweiFgzcpWJ3Jw5MHc/sHJdL
a1ubL6zlyg0peTrmJebieIIiKMkEw4v0AQKADt4pZIvVgsrkxB3Q9nUrVVMK2tjY
CGk8xPCwkLlpbfsN/eBOE8Bx6hBT8D0D5MjoPRxbbJyzVsQc4L4gJG/rQ86V5ldE
aUTIPJbYwT1F84e7hq0Li+CQpihCLIkkRuRQtp3jbH+VtV1mIVcqPDdi5CBBsSU0
zIJlNMSj3GAG9yWmy72hlkwu9xQLPnS6NR45mQXUblCwkTuds0ThyNFve4vYzcBu
nECJs2K2/+r/pIHXeF+lnv+cqiyhdK5OmYDD4pHosgkP/CacpoYFp7g4rgRQa0ro
86D+IJebXs7rUX0+yG2ZpVW76orgOlyxeJh0J/QwwnpqAZ7tYiAfPD12fhnSTm8l
Gy2Gov3Rf3+2NQq3e5wA0cf0IjX9Kq0p8YAcZ4DKCbn/CLdDT7ZPG+hKMZ2PQnEo
cr04QGFKPfQJwVG1n1/yeA7VpeIZtObIhVl8UxRTvEYxKeyPXnCYu7NJuc6dAN4E
FOXDaz+Lj92NFWEojBfVwJqvYU+yCkJ8ESco3JkEreha4XBiHhpsx0uvocoBsSr+
KcQyCEvIZH+hHnM1Yic24Y8/zm9DGkP29fNw9tz6OPV4i6wpmpGGv4H7heBUJZei
2G8++kKJ7flUSREZ4eXuMssHfJaLbHQ1ULp1hzfNe+QyHHJvavcFiSAMZouZ3Jk5
zJQIfGKiKP/n5iuYNKMeat9Wumd2tiwe4ADH9T4ciEgiTJL2S4OKotaTVNw569Bu
BeAB4Cslu/eij4bYBoUbJQkJKyUrgnmiId9bn+KlfBDwOUvGHXku56+0RsIazr1A
2+5oZxA12e8rHW8+stxqGH6t0mvpZUdmy57HIPcvSffanKwdFbh/jUFlT4VI6yJU
MXUmbhT8kSie98x9SZtqKGdnq4YXDKsQuape+QDXlwDuL6YFA/qswTIoip6jVbao
odzmYJJ/1w6F91nFDdiq8Y+56aD+vxrKrt5cqcN6S91MLCZ20VYvS/Wy+QStNzEe
y/NIckhG4ErHqOwfxsCboTvIsJd+f9aRtSx3wMj9pYzZUFWUL6coH31+SyyQf7TR
IpVvVFE+sYh472D7xjRbbs8t7/rfKw4nIPiJ9W/CBB2WvLmY2tMNcOz2DR3DOmtV
ugR/VKHTBgCY523w1wc0ThE8jjteukenQ5mhPb+ux4Qfda6WXokR3O0mBIIeFIXE
qj0NH9cCCsWEwFdFMJmlXLoQnVab/37/d/Y8pMsDNNfEQk8J3SFCTi/nzHakEXWi
5WxTWmcTTrGklynMHOOC+JWZFLZzy06WVOsw309abeejD3spgHjj8rD1L91Yqvuz
mLdvp0jycl+Y/PA+UxUhvVhf0vLr0tZ/tCwom3vJQiQ1d7SChZMeGI5QX42jwl5G
+OaYHw7++ktfUvtpNL6TF7Tg/LvtQBWZb668qHTVyOg0m0vvOLO092FdEYboysc/
hknOwueUALlOJMVOQg/L1TLkWIhCXl0PoFpMnpXnz3/ilvL4roDQrY56wlfbG4XP
wrE4WWvYzmTiiHE4ifbY9KSmjd4s3BG3DyKig2bJO0o7GBS+P5SlDaDnKs3alFiP
0N51YIJfn6DdBWUEbHF2WrMYzJxVuXFeer+vARHzNLRkA0btiHF5V7C+9vXw0ejx
NwudMmSqQA+24csKvqjgPtSpgee5LpvKbd8rh7B6D40jlguTNE44kfhC0Kx9Bo7f
JhjOKAkCklEEkEAL3Rwt1RKt7/Ll51pjG1K/cy2QPZZoLZMdmoeBcOva40XNoyGe
vXYbVmPzaZ+2HvWeiX8llUyT4qHWVkuY1zzQqI27vBGYSy908y3oCglaK93jlsUb
v1/i+kfp00V1r00zkFJiMG/by2hOomVEV5ZTJKSu1dyuQjlZGiw5GGnV9aSiL8Sc
szh4GD/RMgG04/2MmryVMyC5hkZfn4Q/o9J+/D8+I2G449gVjat2LNW6QyDAO//e
YhklzeJyotflBqNvM5hGQhbHZydml7pmli8dQvZJfcuvOMorbtBlVjlM51cuMFH9
daY6waXi+D8U6+9H2b9JOqYnnmlx0kdlzzXB7g/176+JQCZ03VrHPy3l3YsCRMM6
mds2FDZbPc12SvldoTriqvg4Evhqzw+Oxef1RxJZS8Vy5CFvSOwpWhSKhHGu8UzN
3cJCfWKaFvTrw/i4hiZKgm4awlAQk2MCmTHPdA1OriYuiupZLqFG0jE7SL/jPjol
kxB+YVkZV/0OvYwWuBq9uzr2xwv+IEBh7UKMNL9ctVTaqKYBaA2Ncyx0hY9ZAsM8
lMpxwaXWb5QKxURQxakHMmgkv/ovsPcn/V9BVovKqJ3jjDu1SFMhpdo+n0ImHl4W
Z3gijaPtQ4m4CnnCL699DAFqe8TIDyX15jgU4RSLGdsHP2hxg6OvLPpJtjHe/wD3
BVqL35ci52utk0i2lucHQAqyPiQ4OFafVAWWz22e578QLiRK+Yu4NjV/iZe6Q7Fg
S87OB3p1/U6DjVF9RHmLBmnpb/4M1y4hKsjXD9ZlO9OYEV+zZSyxYTy5gy8BMbZp
xvdeJ+Hsmb/asgkM9egrlwee+oFwawZImDEMl+N9wR3FgzuBsVxU4m5gNNpX4QtY
sUoBouWI7o9sD2eGpibs49S5YDFlmdK3do05ZWZvU/RmMVy2wZvgeuuy0vA9AhfD
ZG8/8hFI59mp8rFfAEaWcPBJ3BJxtbq10BWxPUweBQTN1EeVNI+IUrLNLbeqwvYc
UkvhLtN7YHGIpJo6njxbaCu5WlY/xf5m25P1Lhub6HhtmG9r6Y0L7AW4gthaf/PB
2vkKMIGdCrVCK9nf9BKtwRgR66wYIwgqk/UlS7r6KsxAJ2bwb6LNWL5nFPMIjyIu
8y+IbwvrKTmm6GuQ5MRZEq0SliDlxw9UVM6QHvzlCChEuO7HvptblwsCPZArPwl/
zt2sDZ+Kh7Iuy35a6aBAMC9k5ahfQ+IbxbYlLW9vIoRbtmuPwGGId+rKu+HfKBj5
oS7/yLHH9HsoNe2sMVA31tJNu2xEpoiD4n74s4Q5d7HMB5voTMiJcakbcuovTaZ9
/KC6AxvpzGJ9wUujB19aOOgeTa1v7EYiy+RAXZyEDC4uCGWhxfOowsOAu30oYWjO
w5ZNotHvas+J/TPHCeRexIcjcJLQOWG/E+5OER7mAEskJd6ZSEqO9zH6Hg8j2KJr
kzp3gpl9LNQf1Dkr0PxbcqWszxchKpZksvF7IZ5GoymZ7LU2ttBu6EWTxnu4YZQ4
Octl6uGhwYJnTwZaREimges/olLyAIfQVm2upzJBBpEMEIT5scOOOhZYUXvjYuC7
XUZgO3J619WxwyTDJG1BioDyHf96XtRxUW6uOzLlkDSXOcL+NHp4Z5KZ7JbFO0NA
uBtTIAvqS90V3D/Uri3eZvAXZCZnUYhBFt22WuR8kG+QQ6osA3GjrkfmkQbZK2W4
pCsH92/Ek0euWK4t45N92vpFRGjck72mscX5mpovNXax7ScmxJUGpx209WqUwX6T
myJGUmihSezOAdFr1bcivNhJUU28j5q1q8SeW9OUA71Ml78tTjEZB8ffKHyDd1S9
wM3xgGmQ8MlovenfRBpUrctmQjlpMmRG2gLgCdJsUmLPpeG50Yr+RJO/tzLNMP1n
CueNGj5WPLckhX0+DVHkn1ND0H4bG6q8cgK+mqHt7SIgMPJupy4abqgm2lQSZ7h6
IXrwMeOGIilik1dleikS09sLrCeF4c1Tnfcq9u4Fvm0rL0WF7EPi+5JvP59Qa/+T
jHoooitBMmV53Lloq2JgUH6YoSAycjm5V2a7CmUUkSGeMUYa+5eYiQTpBi2iyapW
uG0hX3F+zyyRbcBu8SzDm3XnHnDiRDEOORG284IkwEflgb1c7oqtz61ruXMI8QUg
UA1EDl/02ECWn75PYbI78p+6AtLKufZktXn/4sI2Ligq4CYxLmyVjtv0Q/i+ZQGR
lNVFb0Se5foMu69JfdvgOngUANlk+HbmYOchgl8ActRJM+wauYIkPJiAHGrnCBfp
LrGHeS0QyET+E5ZHke9JJ8Y9z6PpOX3rL2FKCndlLzLkjMcHhl6Xz6I4j8PvqWZT
GJUXKq96/AukONbximfdFjfs3jCGfHDgGXl3bgHnfVtOqqL1VyomIrkvBlTOude1
djwZwAtp3M30Ib2vUKMvnL9M1vs6c7ZtGXolud2YlPhuTouCumm1eXBL8ftGFpO9
QMNBlbapHl9Rro5IpwGszU8Y9AAyFY9KQwEVCDn1bi8q7TJoAo9jL7/iOylym1ah
Kz8ugCg9DCdSXOghVztFIl1Y+L3yC/jXn4Xl4t1fn/zX/4nikeDcDlUvpmbcUbVO
UNDeh2Ny/i0+FD0nX5qga6YGnLw6BMi1Wu0ToE3S1z1K7OVtRNJoe6idFzK94G9M
v5xMUzduTHsJeqV6HssHqc6RGgWa5KqfjRvkx4R85bByr/mfN5xCh4BFnZ/zlwhY
imzrA2/CEpjZ+z5I1rv//XWJEA3RW5zi+T3g6Xo//IVUydMSWtZlRyNUvJS1pj/O
NeB44AMet3CQM3Xnv99w1hfpVCZ7TPx9YlIkH8J0RNtV1GoRCtkFpPEaKirrN97T
IH/kmPQgstB2knLLAPKgQW0puWIIKHmndeKGiMdFYuMEqzPC5IM5Ja8JRJBGJLQw
f9KXNXbuPQc6zNw1jhKbz9NGSYJkMf0sOkPCQpUsRTsq0vL07zVmsvBQJ/KGCrVn
eyctysIsn4fSRNPF2uHL0D/MvuyhLyWmZA05cpyAWwXEz/EeUKNEvYWkwgzmp0i2
goYuTZMdt3E8Mwc1gucORgt/OAlu4Yz94uOs84Qu8GUl8yxo21ZgopOELK8PdRk8
mm8SS1sEDBXhWHcZcMqqAz6Hdz/p66EHGZMGd7C+CWQF0XMChZLTwociizlveD52
kyztMJkKm7UvZxG+xem5ZVm+LdoesGLh9+2S2TTyrXhhIENmuXlYSQx44r7lE3tc
3lcgIuIgNLTIWlUDlDwYTh3SEd6rYxa3+QLXxM65Gwh+hSz8Ic4tOVDIj2MHbwTj
6sbmPIV3i6cHO/HO5gDT21ZDRP8Qw5l8X44UbVNnnFbnQp8P/15tkAc1yG9qZsa8
RZB/nwPM2bU0/nFQlB4ySeen0oRGqlwViJKdzWXLnG85zaj1EYbMWugGzi1T7+Jl
Tf0HFMP7EJt5jBLNc6Bez0WOaHiNe2RouOaRylF0tJXcd1JVK4ZZ3QfM/g5IbVTg
PonsEpUdNWqhUwzoahs/rwNPdRisNjdfEm24kMgainHMyoPZig4pueTZjmEgwj4V
jieZysWHed60yyyMtOtEPCD00y/ZML7c2uINBXVDnup3bQ2AifqFqTHaffflyCdt
xPM6ptRevdU5ZJ1C++AZxTA3ERR1zXEms2AOFdGG+KG2HD77QwFHut9OAdp3w55l
SnIpCIznzouj3iVXHzM4n8GAL89tDygwDk1yom9k1zNt2cOwc6UlME4AcgevI4xc
QWq32x4k7JQ/ZJtx3VRq3AqnSLsQ1mBLqJ6GqD/eoNNefSmEUEGT1oNoJOxksBmU
d8f0O2RyoxaIRRpfMlayUzUe27Jv1IrSFCRD2bRmgP667xho8ivSICzsHle6+kA0
zlxlg/V8oCir8fa75jeSLfR50R+atSQAnQbxTRylgaj8oprbGOMqLg3N8diO1ERG
E8yKuF2nzeS3P97Ddub0tIxBWleVXQ6Y3l4HLOCbPi8BYI8h/UP6K1mJvJ8ASvUb
jqoDqamYqYeS+rFnfd41xH3/QhXLEDOV9snn7WAm6l0++itsVjzer5Cp1HrqBI6Q
AW4ZrebzHcSClLbGXAG2QHACSBlN7trXgO5SywhO5YJqOJa9CthLq9An/5JTIgqD
ljXukkqb7CED8uarm+R0Zt3wA6VA6f6h+Ar2j5jjxOZTnOKsRglghMfNHh5urSvF
Q4+wddk64aH1Gq+DJAkB+Tz905xIAbww2gH+juwJetKForoid2+QJc42U0sLAEiy
QULNhJJR3ayNwIzJLb1lkYWh3WzQz9mto5B7dzBPHsX5SbIqLeW09hjR5FnInN9w
19dKZcytypq9IDuTi3d6g9S5tKXhCpKTnKiTw7ItVGqhj5CMi4+CkdoL4G+G7xpW
B8mzvEb6Qi3ppnBVk/t+8EHzJ51o6mvERZ/QPfFXwwAkkwPleDXDdyyYyRFb76CM
3qlTtK0PDvEVnjNQwyU7kQuxaE53YU6AahKAdut2yrhAlwRD8DZmjiJtOTNiPPy9
g6uKIJ7jGqj/2/BRZpVH4bPH56s5meiXHfnfuw5DXM6LTGsSODtnjUOTOmrjnrXT
esTYUNUb09OYH4ukchvPJ9Ln27nUAtO1i3xZG6KRK+UchNuENipkIkP0/piSlFqV
89APoJjwHIuoOnClfBU2/NKQoJA4Ej/C4duDi1u94ByI5YgvSYirPyjspLgNY3Wv
v+Aav8KQJepQ5LUvEqdc0iUP1ZFTlBPmohadsI0kVLRPVLP2VsZc9G6OnOi64PPy
0gpej4vPN5OLztbuKr0aV4nPqsvVH4bV++Ao+k0hZv10DfyL/Ci0Kz2N6JbAe7av
6zczUhl5LkcPEK9MBUksnFReUBqX3jTfTPXSqWRxqkEFGHjpPpJjeVa4vFHcFunn
dEOsSLTisGgIGVnQpMVWl6cKpcvf0OJm8Gv55HsxFGfUMN4jNX9appnsqGhyKcP7
k18pAFEw2Jtxn19vdEE2Lp/YiOCnCeY7cU2V4iIXA8eUbIkl4QadKjQk3Var2/n1
9wJIsgZt/HAr6hKwyHpbJJ+57dnMPrICi0trKuLTUuflP6PADJybTZqVP71kDQeU
Dupj/2xlOyY3XHgWv/JMEDfQgXionhULJESEh4hOqyMyS5iYzA28a8WoS0+1gtcy
kK1GyVVBf+7wPldTikLF9ZazbkH2WLku624DrFYeUwu6HVnYZR8jXwMhxMMK6suc
m6eZ26BBH6Q8Z92TvhDfzDLkZ5DM4tjtEOiION8kDu3Sq5K1Th2YsnWyxNxGbkyi
dZts1EiB88eNQcnaokZamSPIWZ8gNnmd837J58YlUilHjB1Wmkfi3C74b686Z8pz
uOhUUzAAH33jK3GfkDw/zexAC+WNmErBIjVTVzz4NzU47nN/7DlcL+At6RFSR7SF
btQAo63eHVGkLtVw7TjSohwSwUhX8+YYGW6LrCWnECytLfb7LGKnfj7z7gDXGhqP
qlxsRCHXbYBkyIAKF2a1uTiUgsgJDp/RoY2h+cX2yT7a8YNYXOSK7vms7FqFiy+/
/MqGFEGelNk42Dq/1C3SIf5wKEynQ9NHRbL5ZUjTKRn7cGf2OhP6c1mmrRGIqZoj
/RG5sHmbEejNgrpSWZBC/SdKQFryIjrO/ChLN7/sgQMREmGZk7918iQGs43Do+be
F71PhRw8uzuorY7Jdr3vrOlqdavGOTXlr7Q+rGTdQxajJVf66Rwptc7EzVnbKgvN
QCh/OJoAbzWKu1DzYwBR14OYtgDjWmMun5aM54D0SlN4jppPcFwfw+39WXXQkyAe
QN2ruwSPLbixK+cM8oVg2wW3e2qU08ig8IQbDdApFbxb6dpQwjrfzYeEaKDxi8Yf
4Sb6/sUkYRkqSgPG8V3VY6Jc01+Oef7GuhSn9xRhZxPt9hnxNvJVsvofSHFbKr3W
fsFLoTC/DWSRPtXHt27cokwVdswmvqWKYDzsoC4hhUO8DqyvgnAiMxGZ756Ki6ig
Hz9KPVd+95W38byBsCP1N8E48RKckrpHiHzxADsFVeEYJ4R6n893fyaYoog1U+2E
9hk1l+dTmslOOSgS1+duSanFgwcQXwXFq+V5mS7jjX7RrCzMd00nS9lBoDzTl1yD
XXOo0cm2Oq0P6ZokRjCbJhA1dl5s2OqVGqwY5NOWr4+n8frMOc3cpN1IIMN7AwTk
0WXikiUYmCvhsipPCE4gxDkNtfIBBG+T/7ZvbsgIFg+6qIM6SAmELvCieKCAoVHQ
gIr1G842JUBjvLhhyeWcz63gT9slmXz5HySyO91gNh27jwXNd4EH35rAUVBQipUE
4VNhyZJuJj7I5kmYIwRiMk/VBkuPiqWOyQvfN+L4wjbRqQFTL2zQQo6AqJtCBRpd
pcaNY+LD0mcPv4Lw/bj318XKl5fXy1lfeGfEnI5gn+Pf6Q1qMqvfJL4lpwAemlvy
KIX+u0m9cRLsz+AGCBUVEf8r7zr5NIW0+LS/gifLYr33jUxflNxFTq1DEyVT1Ern
7AorqYhwUOuKyomFlVeLaFEE3x5MongHq0L8dNKddunromMYMJqstR86t96Daajc
WZsMhSH1RteONLKH8cm+l0/Jw1FNsXsV0SsvjQfs0O42nSqvAvaL2/voq9KzbPmf
aBSXkdF32JYwOZJA9+pEHzDhI+D09YWcszGAm3pHgrO0Zw6luBzTLQ/6oXeGsu8/
wZS29gFJFqE8IqFSfcXMykJ8I7BD6j/3JFCcU+uzu+k4WRGNcO0lqs4lyCeQwJve
RtTHHEHuZtq3YubpzHG8aFzCYMZCwRegS9nIuwhdN+b3DuFKaM0h8axzsrkE7Sxn
sjfDoxTk3024gSR9TGvAYtUMcA3YUtBVMihV2SRG7wn93ooZ6FaZW2h/L7hLw4UB
a8xmGN8GW82H/Pg/ThPCVBp/BMzX3PiLaGinXJ6CYik4b0KGctPcGxFO4Mv2Faxd
jLP7zdNEmKdj30yUh49jrbJ7zIg2/5ZqtvT6TL8ihy9UZWDA6+rt3wW1qpJ5pYbd
czJr9Q11/YBuwuKlyNk1rZrytP+06qOGo8rgTVCizpQfkp2AiP/vu2VVYytJB+Qy
3b5w4bIUeM/4Pumv8HO6x+H8aE5NpSEW308+umthPVMKEvMedQEjOEgd9HZ9DagJ
gJGjgFkIAfrO45htIlZB5lFtoglECebUw9ONDT85SAhtgKHuV3AV7VCpS3xUm7RL
nxaadPBZk2ro9OBmWiLw+kjr8imV0C/Rw5ZgeTuAvH4/0tpnO6sxPBbvs0xwZT/w
5wVVtM8X69TPn1/2S9LC9g6KFKCpqVLZtkb1OBE82QuXh/fOEW2GEqOS3WPYI0Vr
N39+ivuC1bVaVKJUi/5WR7+tDEgua/kiLp72rY/hWoGKGf+jnhkJ2QaF80Qd61Kf
hACnILaLlVHBsEESz8ugF+b4bGIbKoKRbWnkQJ2P8PMoqL8QUJ9EMqPApY6H5/ph
PBLFZiN/2iOF6F40YroO13ndfI4YUxiD7iwF4swSSuKpvo6tfeBMbf1CnmCZpXR4
/t438iVWs8dHXNIx04YEehRST/gW589b6DSaMFTNUPeLGhzPB+tO79lyWz/EnejC
wf+TeWU+3JJeNozZt4fEIdYfoOAbsAIZs9vLrfJ4vxyCwJjr3/+/IBYVyRepMVvM
lOYxbLvhWgCL/kKTWkbgyex2O3Qq41YWBMlZRhsttpA2GEFTzfi32NPlVT5oaCBY
4zasKudLz+RWEbbEl2FvKu3CNzIMciHNUp3jycbG16DwoM00DTls4ZEWloA53h2v
nyGYRnmAxgePW3cJD0jW0S2maue4WHOor2ZbvG5nwaS8tSy+/vbUSouzd/7AdI33
FJkqPFoozUJZBSOKQVXwh9K3Bj36cdgICN6EAUEvJ0wL6k479LCANSNMA1fgDesg
IC9+BaUwRlfisMMNw8AYZ6rKdZHQom5z0gH7P4xnRumX3HHPNgbmraA+c27GIRYO
fxBEwrsh97lvPnyPa0qaAExXL3RYNZA/F3+ToHvBQ/LUJWdFO4+ume8Is5SLhI5O
jN+n87/QsvXLGpI5HW1m5p8AcOKxmQr2mcXAIKr9Ylbe8AT26dNimZ+9miG84fs8
3l/Wqtmn8exv21AOqAiQlsmXHGP8JxRAC6EVaCTHDk0xO9aRB+zCYMbu1t83dDwj
RNAJPJJtxPPYznxco1nr1JvPykHvCkWlayBeOu1U2uWlSmL9ejU7GcfdXVKYqVyf
eOXN3Qyxqm18cm2yZcs85UpjxsshUceHmIZuUBJFW3XKpdZGBA6L1zsOR0Gbn6em
3rLPLAeeZgCS7s+ifir6bL4QeBStcX9bB82omRcIl1eN7dBR3UGOq4YpumQM3FRC
tq+9jQ8fjlgCTV+OjszcHVNVNwwyIdwIzEp9BYgpOrsjkG5YqjPw++pGQWo8Fg8h
tlHgCCgHkciHwdL/hZr5pJgzVnvGE3b9V9v+Tkhk+YfGRB70Z2svHwHS+NnjAZbL
zIvVS8uSyJBAe/QDojQNKPD3x3AiiE43aGSEQa4oXlPBFt39QRvOhfWOY+PhGznY
Fm/8dhmtxb4HRfG6utFbCU12kdN8PK76QZcyDkABercaFFFpkbDssqkbHVAWDG1P
q+iOcUMSZQUYwvsDzf8p4Bh0loEDSGP0taNEN86+Fcx59WGcgAoL2muXKMt35i/E
SJ6KiacrG4Q1XmjBKozbMN/gHbzXcSwqrAg021jeIitXU75gOMSurwyHsyTa1pdg
R/LaqlekpVWY+8p5OITmS6xg9m14/luoT7EZ9ua/uMksPh2afNSMLnoRa2SV+Cya
blXdIrOj4Bdmjzg24nBA6k8tTCpYnE6YFH3KEIHq7p5hi3+bL7Cf2P2oXumrUjHz
uvdkqfLThjgeeDsnN2zAawciSnR+HHvtv2A54ZVhsj0DOUzJ1zb6ysLpyTrMR7Nu
cqBkQLviXMZ8d1sMpufp3c1myrBwPLoJVpW+ZCE+SkaqYRq1VdnrMMrDG3zdMBCp
ibJhNmvPw1sQM3CU89/g6qRLAM9CL+3n+mfZ7Dl668VLkM4vJeVdBRRm8SwNfiOw
OEacMV9YoMhnWkfR8R8CCJO89+MY5JciU1gY8fsQ2Fp/ANXHvJVpqFPiHZ0PraZo
zYDhrrPv1FCls3xvXKwkIeeLZApVjwD/N9km6tGiTNKCcakaWjj2k/OSkeSrwZKw
tGh+SlSSgKC8BfEiAJO0lBtXJCQbOL/34rnBQRFyOQmUgVtdiQYSy2mhYO2jnelq
YKNxbS/SFFSwL2pyOvoH+WxidHXUDNDzXIsI3qIwwyTRYpp7Sa7TqnDeUhH9VVjr
WTRwfa2MHg/Lc9ThaMgl1UCbEz62xMFkGkNcnF8isFhF8oSp2d/M/fq2lFrjv4bj
XTZuzasAht8A5BXzH80mAaCxPR+zrd9UqyDSK/AGz8l4Bi+PQPA+kw4a2C+BEKUZ
ImdtkvGfySLBIdnyy4n/jdsRkdAPDZ8tp1SUjsyKHcJzKkrMBDzoPglJDo0m8obm
H/SxfvrYYYXZSPMbFrqWZ45E/nDtoycMZA/JC5fvbtFU8oCckp6V9Aem8rBsOumP
VYvhcfuekFDOwdauQ5c0xDkPY+6fyL+fbPz0ShjIv4mRUjlKBKYUE2DrZTrbrbqb
7tTF/PRX9iEVdopsvY3lIUnrq0LR+UJJPhxNqkV9Ph9IpZi4jkAqpKy3aAyR9xfZ
2yifn/1TkGoaqgJI0XF9jsahpee9XVSSXOKxwipmyQxOhSud3rTwWnkFoehjBvAX
obwD4uXBsgjzQFaYoF/SYUlJVstTGZTarGxZwXTyIWHv2qB4s5VKqi9krP4d/J8Y
iudho26zXwwpv4g46fQTmW0uMCOJyMiFVD14TjNF5CvW0FpS33IPqWz66iFD3hwG
yhsLnwxyA+S1M5uBhYMrEFzj6n6Ld1XPTUFN5HPNjMXXE73x1YogSB4tqzZW/MPS
9Sf4CQJlG2PVkIr7oaCfUFJ3/f0ch3eZeYo8cIUHePPYIBcNXv81R7DOm1Ir9hCu
YH3u8hjbPtw9Zl6bQsWXIuWcD2rBM7OLD9RxiyrSPFWsqXYX/SYyVt+MDBSJ4lpW
GRH0IT7qmNfPO2VlavJiPu8zd8Ov1jF9aonx5whRac+9Ky/E1bu75SC1x7iUhNOH
hAHc9Ps7BEieb103JUmTl3+UCGQaBxxXvcmCE0v/q4cDnOXq40GhmaHYT7obisbW
5i1bBccM2TBBNWxRDswi2eZCyS8XEDArU7o1Rc7t2RaUILsq+LdZ0GOCtCoi5pNt
kdSn9wuvlobyjLP7UcvYRG3+kDe/YlQbV8iYvTQp3BH+l3+V7hMq2JNpoBcPaC/f
Q4x3Wsvbeia6uZVNYTLkhrCfLZ7qUICjXs/glhn5rYFnHtKOaHrb6FIWxfnkk2FA
dlsU33EnEl8xixZiro7TLSJugAvxFkY7dchN+eC7aIUQgeTq8c04IG0DLREE9BgU
isZSaUOE/zoYXF6CJCzEnVbbF+oc8TqZnq7LI2uhZtJ/gKPeltZwaQGYzUDoYFyy
BTjWEAKEsTaZxr6SA5LZ8hw1oL0AgP1YG7IKrVqy4IvJdR5kvJFX9s5obNI7BFu9
uz4UqLcvppKsNt32Wcj+vXPZySr2RcwxnRz5QqeBqSGLf3cQhqvr3C3SGuNATrY8
25mZALQBfOEodaRHgJ88J5Cv7HRwOiJ0dZsa5d8HFsVYmTY9q57Q7LBJtprYzUQm
5TBx9nu1+HKqceU8saok0mgIINRY6ZGfL6ARfRbyIKSvNEamWuI1djsgO4KeKOgA
VGQf+DPe/88dS6j2Umd1X6gElBKRYWEDTHzRJBbwYPkf1oHDvB1nyfinpEiZ/ubN
eDNClJ8iVNlvoC3vGM6J/MnsLMah+Fvf6lPfRyAA2p0wXupfS5c+SNfEG36P2iJX
ZydY2uBh7LMTW2/73pcoPZkLu6dcSoWGXOasCxZbrZO7KZVwwa7Z9u6lIxhRQdEh
CcuVkwGqcsmbUv8+SanM9nLgYnYWDlu1omfy5tjSi4oNInshSvGuiwtzikfTUUEc
7gMN1vbF2UBAf6VmBXxSoZDOW7Lo2dmwh/cC7p6LqO9HjPl9NRApH1wphTwL7zXp
e1ZVB7Sj0FSOot7vycmp0D2AieTxB/gYwtTRX86o8zTMwnodDx7Y9LwwnZTd3RNf
SNaQSBKk+FJk8+2fn6hBjaln1sf4GiNy+PH9gyWs3s/iOHQy0+7SQPcWusMD3cXy
ObkGhlhtjxhAelG3XYnwCumLaXJfNfsPJzOdRZMYGl7npXktVpHzVd6Ip19QBPib
Ni+5GU21J00TSRyMIImA4PhgaZEFnGXlNYL5yKGgtUv+gwTlaiBo1bunHvP1Oa1j
V16JAN1F92h3b7F6WoNIz/SVszQjxKj+nv7oS6SYg6S53wUCXc3gTwz/BYgtQOaA
HbRabhE2kc7yKk/zQAimlQUStXBV/VeP8n06uY34iMEjPiC4e0343R3Hu0YzKwNs
eQHPxesB7O/xxXxbgV7jkIFrI4a8D63tjh1GG626rDq63wc7aExkzVCTl8TMmiPL
8x/wg/1YFFP8hztWYN4B44IERA5WWgkXOQDB8ZxWViDQHgwuWSLhoaRYvAZNpQ82
GuGD201MPt+BzPOp8nEU7Gb0RWod1vZc3u6m11I8xxrndEwZrSYPFuvJp5RnXaI8
x23zqJALgz5gFPTL2n74AtSUB6U0+z/D5X05/bZch8LbmiQMpVUzQ9PRQcL4Fsge
SFT5f7BwKnIK+XC13q4TCUq/Yjg6vV3K3vMnUo9AX+1X6xiUhMYuJN8epglsr/Mx
XbfIKkFmDztKnjCzp6MOzuSLXQiZ6w3h8NXszj35rG1RwXRPYDLdiYVXNk0HBWVw
TEZ7MnW+xbT1wKXRKMF7mfspq+4IlGxeNJ8J7btr/3EuL/iIOISQjR7uLyh1xp/3
u3tYT3PQblxx9ZGN6IxaKJimdrqO29WWIkw3A6zaff/K2g2WWWws1YICAH0/yJu3
vRMv1ASKW4iGlH+PrLWbGogcvH4KHIcVidgO+YGuSS694yR6SpRdTzDCYrJ+9bAa
iJhsDG8DLyEZWzNdMCccbUnkqF6+EZSCcdP1nYQT6EFuibTswfPF8P3OwXAcgO1S
V+i4d0YG6NDsIGZT3a98mFvF0T9VKpUJwA6BcCyyVaXhxWzbCqfWAFmhf4F3noyi
hn3ktY3E64RtmSe2wayb/TX4HEcnjv6IsdGCbWMyKOPtuRyIgu8eoGgzEuxFsrUa
VzeIL7mqIZkXMC4y5mJwJmK7+zvK8UbtAT01r7KXBYjI9+IWz0YAfJHQ2WzeyENh
cvfJiMdce8y9kWzcH+QO5wjJwNEOOFAg7c4K30AlMMOJAffoflIP5pl22yWh1/PA
r2tzPkq9E4mX+g35BmlYdRIkHFcyiIDqeMU5HzSSUIuu+9GTKK88yoHb+Wugs7oA
SsLfuuwL7Z94Zfeh7M9mZ9muRZTekD2ZDzFPHHD57lsk69ZffKHbVGPXwdHIGEG0
UIDxw24raFUJK7XG6Wx0/q0NkQ3TAnmankilDIgY2j0MPpkwFS2iKP28wlNynR2n
sjOwf40JYM1QhZAHXqIyhLFQrL8kXVhElTMlCu1qHD0a0uuT0gRKwk6NWrkopJ3e
XErRcy/eAzYKPs4uooogdEKT7LjAuMbQ+42VZ+ei7xM+TiKMYbImmUy2YTlDSd9l
rFV1cp9Bx0oVD+1VOVfyDDZ4RN7xurGHMVpAdj1JopnDtYah8Bbm+My5RPsyfy/z
zu0RNbFavXQ1cZecUkXDMJ4U0YBBq/smJRoF5uAjkppqnxHd0/EGw+sEZ6InbaAr
nfD9GhZo3q772VUt0dv3F/33cjhmJE6H7s2tPQO6WflHrx1KFgsQi4/U0eUYuSkn
tOG5wCZvcBFNuSDsLwOTskgR/rp4MgvlbDogbBme7ZBBzyMXh3+4hVCunekxkqQ2
yGqL1W0jECc6Y4EfcfhlCas3w69p8EHiGIWY6iRCwsabpvCvKQ1xTt1D+CQCNfxB
4uHLELNtek/+fXWiuj87XUDtlwhLB8/Y565xD8LaShmIzLLJyRl7aEp2pdUsieZ8
ToxaOitTfPdoGMVJ6Lh3jrqG4Z2IA0zkAvif1WxYHA187D+H/DaKXng/V2mnilq6
JBxcm8QlXoLXyX8BTcq7q5xbM2ZpqwETmDQnEbKyxLuXzV0E7iJfqRyxPxW5OASE
S4A9dc86Hcfy6XxuvuDtT/fQwF+U+QOFLRtzv1jsY40v0zX/wA9yGq7mMQWUKiOv
fjUyv5AQvT2n537tHO74zeNJEc8z8yzp0AsSgB2jth3g1OqngXpcRwv/5oVLONWm
j8DlQFyuXn28ekpMGh0xPTtHBye1g0fze70eQ7mK1Z2VAus/zSMIwj3Sh28gkwDt
fWLYzGPEjGCdP5q8jk4pslmpZl8OELDbDNm/AVEZrAXjQOhbRDOPWx+6JEeZjhV/
z0qJVDv+DCoB7ytge4Nq5QVxbvLyuDcP44uY3OKNJCrl7CKkoJBOc7t0r0wL3zxd
UfBEc0kSOhB27zR4CmtquCC10bI3RH2ZUuHHacCq3cqDjDeqHw9S1W5EHTUnDLVB
YeuoMwsKQvaKIoV3F1cq2ievHAPDPLQAW5Jf6tf0uF5R8GvMan/8qj+H1Dnvv/GH
UNhp3XPNjWJHiRruJfnCMUcD1hsJ4HiPmbZPP45WjEpzDdruim3Lb+6jQ9TjJ5MC
Px1i6/RBDv+lmzhGpvGXbWcrFrAbULfvwfclnojturzpIZ5xgiVx7muIccRK0qM8
qATewKIZMofQewrleFALeFLetDxun3SZqc065ZaiAHeEk754FUZNDHiB4xZVQrKM
LuZ2mNr3GKy60MaMuy9SslnbidRvdcqJ49ESZjk7hmWYEkHs9jz1q2EUrXJbzgf+
HEV2YziRrsf4vPBzsNpcGFuUCbTMjhcAEoObNvVDwbQb0METAQVejRkvJtDwgFqF
9zF/cCLlVIilJZFpjnLVN1k0m183faAvtH1EXWUmQZal9PAOCsOvoLRN6gei99t0
ym49N1PIvr9/vgPVLesnjGm0kMC32hFpOhZqNIIAa/H7zHDJ2xrbK+o024E3COht
i7LnozE5PYI++MYzOYQDnB1lpXTCqqYD3JRNkXN4pu6//cz6iU+EextvuBYvuEaa
p+A36u6h0rKbl8OarLsG6n+SPoRw1j7kRNozhQq7AhrRnD99c5eZ2K81iHocx9TW
klXNjazPQpFyF3eOnutn/2dGA7b6ubZOLbGd+BtwnThbp3zwq14HZ+qhAqzDWKu4
HbA4E8pW7KHlO8JgrxvrGA+Cr+WzUoCcvUepYB+yeAmVFN50SlJll8uQOrHph6PJ
M7YBLEdpO6bJBhwAXLwJojiiRxZfQJa9OPKx5HACrC2gaZrEaCElMskZwkOKwXg5
bOaeyRirVwC5l74UZp2Vgn72Y2Hcx0AdE8m526jCOAyStSrC4H16t4uWFKENdKgj
tBT5iCOkcRM5RH52mKgIhWtXVDvXPV41YilwV43aR/u5FWF+HRitnYuXKzUTAb9i
1+HeafrQKkEc7jHXCFL1Xv8xV2u2UXJSlnMTeDttTy/PlJZ57T7XHZ3GTgNSjsCR
/5iT99mnioj1lThDxE/3Wa5ErsYf2qZ+NCaQgRVgGjhJ00nlYQiyV57ABVe++gev
0DoiYdblRf/xOY6ttspBrghrLtvW8LqeY3kEPr5AE5Fk8/CPleSItm01fXW02Ers
vDgZvrFvpNP2XWWjYssucpY9qlJngfw8zxda8xqE+zSdx9xoZW7rplf0qtN2A82u
Ty/VJw5LveXxxALfvK3mY/l5WJsW4vD4tUeNXsX4s/h54ovgRDneslEkjL+4l7G6
mHujkxlUeE/TS96TROHUgNmBfRED0WL8wqAE6ymuc9UlCcmaY93z1ksDQk68mQFU
iQs0vEt8HTHEPJ82fDqwgEBGxYN9yr3bxjvK60lta1Z38bAogSwQroN5BZam7BjY
DHipb0nZRx9MQJsSUkMh547JxSHRFDYQxZ26icgVgB9+zUSV8JaFF1UgQ+++vwEu
EJgH8gzM8ejeGkjSoh/t/q7j6Te9r9eyyKPR3k4/WFZFhqgZMDY/oD4AJkzmd1VH
yhz3H6RVwlOO8D2X3cw7ZXpvBNLU4P6Sq7ZivyipRXojp4WvTNwhwElj6G6fZ5xF
XAXuErdp9Nn9PLIAq3OO3873Kl6kOK+RVCic0isaUu71nYTPKoB2tictu4wB1AQP
M5CsmV1XqrtbNgESaTZnQqTaHqM2jmxNGMfyHmpeeV1TfXRGjxw6An3PftBjjjXd
zNH+0qxgzIQpBhVHYaS2OST3Xqj4P95fCJkimI/Va7CtDYXBaTL0aKt8y3KFT7xq
jFsmKibGSB34NPAXbM7B+FgTXlsXfbRYQJR7fcInAp/B6NvjvNkM+wKhlzXbr9Dy
1VXXP3PReGoOkBpPnIMF98TXw6L4y308NRYTf+fzeyRO5Sh8aa0m+Fh6S3J12cTr
m+ubjOh3tRZBJV372mQGGYCbKpzgk5iruQ7w/bskQaSaIQy+ReQDuu8PUFlMpdt9
K9C7HP0JDDgh2iXMq+oqlY9bc0+pieV+EmalVkNkRfL/6nl16V43uY7SV1hscbDr
Q16+KbI/AnE2p/+pxuMM0s4pzsocSr9HRJYfxkDsAPKt6MD6rcBBbk7To1lPnNe3
oqir01CwDvnoF4oR3qBVi78s0GJ2s9ukVg6YK7/9eIvPAivc6lk5+Mi65fYq/g/b
vIkhaqWLzLXyh3YS5HsWn3TyurI+PU5jKpIWyFnuPYP3XSq586xQ20rxqSkt9q89
FZqK3Q9MEJ9iD9/dmHP3o6U8bACxvE6fSgp4jJOUQt65GlgrtRg5itrSA+N5wSiX
o4M8oXozn4z8zaIvCY31g4sxf8X8525BAPoSWDr6Y/PmvYkd0YDuqNwhrKmyjxNX
j1TxWoDjTLvpPXqIQ1qpJgbTFWZ7Ld16habFXJzSWVt+zmTH3uWlYDI6Sc0N23c4
ZE17SpnmCGnVczKGwfKAPRGEJXwuFvMe3x35NY8idoUtvWkii/6ghYjRqIHVwLsk
nEeOukrSd6kZa9CfeaO4dTHIP2roXBxdICHplLdtxOqoYSkXpVEJ8QYGMgn37MWd
gv6je7Uy5rKzSkylDyDj2InZpDYFhKyQ/oaY0s+KUDYB3yXVptkPA1aNBCPVOl0A
6RZeUC4oZYMnCuSGQ2WJAxfUg/voxjd0rqN2kwhP9fTP0u0OTJAsAeSX6X6PRVwm
Wo71E2iEKXek8j+g+zXPUPv5Ep4dYevNAKCEX0AUnp9ceBzvqi9R0qTNWVmyz9hh
zC8LHd0FkUu3M3p+V2OsqlwVepvUCxkE+zGMWx+J2rZq5FAVvMHceVrKV7cmlTd+
A/2El7nV5S3VciSj1DG+97zAtVuc2R+j+tFcw4wvB29UH0mzBs476xOBsZ0YfY4U
RKVWpcOYiE8JFffalYr/8zRbK4OSfUJZx50RqAFjgrvnsHq+mM5jxaZNYjSroWgm
DEbtbbv2cibmMn1CMhNeS/Cy32nxSxoohGc2FcrMZ0E4DzcfqlcSDiY26wMHD619
iwR3rBVMFTNAPDThdz9wLbqQhHlaOMxWzFvOHExBLeQ4PSMu0b/UpzL48VrjKc75
jk0nMWofRC4Erc3DFG8fQLb8zxDXD1aFPs4QvCO1v319aKnfhhhP3z6UqIMbHnbq
6iFt+yqAzKGrBW6NoxqshWPB5yC80LDK/zY/74bspGeGnr+6M2KHhbtgTTSp27yM
RbAvtTzbs2RBrxWeZe2m/w6I1/mfxq8pwvsoXKrhmrnQh3/bdYkT1gEE+gSyocQ2
4wC597aFyS6ovv9w41hg+yG7Vs9S63pndOcUrlEGgtLY0Ir3jfo6kk/E3A9pYcBM
/ibAONg44K8elb38otf1Du4i0+FOr/GF+Cs4hGC/9qQyj1POYQey0H3YWb2Yp3AY
K3aIoYVw8cQkEbcxe0CmAYidf9lUSMISfHp/WbCI2Y3W1Zlx+hat8SM1D9xO3Y3+
/ObL1KCrhRUvoZm2/hPKlkktwCA97WA/9lHSugxUvL2iEVEQ/lsO3SI0Mb+anpCp
HrsqY3OozTXhW/yQOxuvnJmJSsBjCQrzvvk9ZM8duZNRoUwNVTwS4VY559HA2CrC
nwECatAXdC3BtcmBvH4EGI4C+lZPSRF8C22l1Tcwm83NbRLmiUxW09HXGNOp7ugH
gHybsCNgZNG3xuq5vWIooG/FKmYSnLN0s8PEXyY4tw9Ea5K45fNwDnfcve4jwk37
kgSLScWNNpdqDOVlZQpu1hpY3pnt45OhaY9s86/A4ijCXv6d5dIOl5ohzP7OxyNC
rl/OIs/CgxFYYGwE5X6QDxTGWOfclgUPoe5IgRuL3nlV/IGXCpaIIYqwd6TlZL50
1JCtzTFGq/wvjro0z8StEVjerDJuRm6+CZoNUkJzrffiTk2TdSMD9GyVE6Zb442R
CwXyLfrYaACs48qzMaE58qhct3p+MtYEPNbEZSA2WsIHqwQ9EfAF1ap/6OHVRqe+
ypDaLBbhLDE1bGjFoFWl4mRMpMaiLegvqy2PcxlOqBXaAIvKOk1lELY07t5HY1Di
SQ+mXH4zH/q8WYsuebKSzduL4qmGNTgdOVO5Bzg6ElCic+EczijSHcHZ3qp+wYWN
1iEKTdHU2Nqr0iFpmblVIv3a9NX0Mk501F95oiu1L4s5GLD5uB/hh5QrsweIN97m
6do7HN2rblz3bgV8O/G6IXkowKjbdn+QeMFYrO2D5lKtTZ3pob0wXZFXa+xaNDsm
l6nxLWmrPwDCxK0rNZieVvkJ87t+qmLKN7k7dwGPQgmYvkccl9c2u/szYWIjmLBn
qoPnOInS9MnbzN2Els10aup3Rk0kSbbEqDHBNmnN5qrHUokByCYCluZ9Pwfpfr+d
kFythzttLy/TzcBLyjTOQ+u1FrJpZkyHGIaMcA3X2bau3jmV1+ut2xAyHtqATisF
KgDWv/JuDVfhErp0xCjIpEWwOMzcrVdo10+sJseSmtKfAftXC27Y6kuDqh0pCMyN
XHYvIJHXNDfrU8Bxi/rApQtshoM4BqWHjuHmJQCsLvk78yOldSNcVV8hoT8ZED+M
u8uxE5NJjW6KSpA5y2c3vLtYIJKfOcuYqufrDykxdHT42iJrGwhHVXKHOP8UBG9X
jaBGapYonHXuNW4PJY4l6RX4WubmEyXYkKF3NqN6txRsskUvTarzDs93coGypbgo
Qyb/F68NpgTJf5A6XRctpxUR9sh2qk0PRWbYXWwmrf4RfbxdDkFT1fwVgKx6f8ha
AXOJSw7VESNF5v2mx2HHXsxVeNs/VCmVs/Nk7VpqfOXmg7nkp6ADWlU5IdKqe86U
hx8RRW3l+mOHKSoDq0I0HembS63nRXuSVpt+8B8IeTaxN1KJiCGstFgVCe1Z4K1q
sY6KcppS4pBvMnOhOv9qxDU/U9xij6bqAyHLA2nheKffI3WuxhZGVuFS1XewQySu
a2b0pMld6APHzmuCWjxX0tAsYNfj1+7IXVgWWWiO7/rX6lRpnIhKrINxRj95KkWc
E81YfQL6/ylODJg4UY11NF5zJBK/Abbp+RiM6XGKNWwnSVTUUvxxH7FMS4Bj4RRF
m0eIOZiVwRIYirXvIFLh/k6zeJxk3ufwXRucVhJCh1S4ZvEuJkdnAUD7g1e2XVj2
5sbBlt0LB59pqBHykiNidABcytCUfQ6a6+66kgAnNzPzHszIIwy2GGzcOYm2EJ8b
10sjWQsVa9y78Eb5EOV0oa9k/tEeS4HMsAbZPPt2EF/HBxBOq+naUqc8x7ttI02A
ZKlu7Uvz7p+LZWNL44HBTAcFnObIMkYq4JP1mW0rUMlysNTyw2GDYVPMX2xm96oq
IiGWRAgPSaAVvJN499qzjfejCyyqt0NZa3zXPUxqtCg9xO8ESfgHqloMkjxPi7RX
/BU0vp7zgULllG1/9Apj+y5MtytaMsksQRh8XshTEYiKABXxUAnH/bebHEKILERa
VUv9sSpopSlmw9xIVKtxi0cCajqsKFv42cnDWSB3RjxahJNP/C2YtKIONMNU761B
9zostsba2QX0BZAF+kixruDoOwnKPajmOqlFGnpJtcH2oX4WgJfrfl++BoGH/Shi
GjoOkAhyoXNGE1qbI32vgBRujq3nxj7Z7xGmwvzQ4R6UTiio5+gj2OO+fwW44YAa
fewjwmDLIpzG0fSO8Lcv13ylNOxGUez0mw+KaP1Hi9MCZHQG/vnhwTV48gHor3lc
w2CO2/VuGBVMqc+X0XrpqVVnTKe2DtFED4ZlPzHz1r04IRoNFzMBCXlvbKMS/HL7
K5syi1VYjj594aTx7kmXD/Ws4hfCzTLmX05aMr8+pUm/J4qoQAbofVvdugc+h3i1
SRFIJJvbCM0biWNt2q8Mq6NCzMqtaeoEiJtzS2aRpNPz9Hd7Mj/4E+3tt8rtUT3x
zkaPxpaVaxJ7Eyrp+T0fvTwl6YxU1rFF32xK1K4nGkR9UYWOtTdpuBsrjNrR9jTk
w0e4pHpfkGS4f8nPfbiaTkiTR3oi+0pvZxYcW6ZKN4/wWSzvj56pE4GJfijcQ2QP
c8BcDYIrSEwUmF9o20tMQZrK03cMn514gNGJ4Bot1zbLknuGwcVPrBcfa3a4kSoB
6rs0DdeXWupv9CapCqvKikcscT1VPYSz9SJOkunSHgtRtmWqtap+JFByHVjI+IAI
OzgP+42OtDtZBgScQaNE0EK6wQ1Difb+9FIdLmVpenunjM+gainMe/CRzRTSAlhg
07D3HqOoP/C/2AnbrkO+wkFS1ZeBrNb7z++CXqFJdQVULMFATGoQvS9SIVA87cKn
3ltbOxnb/LKNgRWZ4WaXNA4pXC7wydynvcDw4/FlSLxThzol1r/nnsbtei19W4Kj
M2aJyJrdOuuryIn4WeSG1dk+3vgsifOaRlqzOeLJmlcrwqhLBjtLqH4S300VLvOD
eF1Ukjaz3UpI0Sv8/UsNIHMQiTc5S5qe91siJeE9SWLgsa8+VvqmsbuEQGBbRaoS
zMfRL3rbc2+87CIcJsZgEo/e7pTdWqMSypsZ32yjwwNxMvQ39SdrnAiFFH1gJan0
xLDYOT/AyUu07aa6/UPRqDihzswCb7hjnhsLCfG14xJ1t3JyiCb+EcigmytnpmQY
NpsgkxSJgHX9wAj7qIl3A0mp6C3AVajlZMWmODQ5bQMJxzFFfer6LMG3jeJcRAKm
WAbu00DiA4g5yJh7SGvlRBv85BMjD/Dovm3r5jkoas4LP76lySnNsVsooR7wXp4R
zmdCE7aDE/UdbGWD4k3BAS9hIiBYSaV1sWv8latcEcqh4xDpVEIvzCjivuDHtmab
fLYTjnS15sBMB9Bdv+nlIn89VlQkHN3JxafG9AeGlPr/YieD475O8JibBt5FayIg
ydovPBv5R2RwmoI/TPsIIysxsiEczDy5O+SQ8Zk1vO3/f4jaXUtR+5TAa4rvTyzW
bml7Gvd8N4KAtTtLfSQ8HfyQ1hbQAAd4772eSYweZDoz9etq0T36eDJhb7mvQIN7
gvVal6w8JiFA7qrIjYvFi3ecwTzHPC9lIVRIupnE8XWpr0Gc1Fu35WpkSGCRY9Aw
g/iLY/x7c83r7NC375ZbNvyzwqouUdK5QWh4ZhqGQaRCFyisJDAuGujnDYFmm08J
m5LZtfhemd//GADeGzBDaMQVgookuL8hm64lvAQ3s12L3oWphVWEVrpBQ9Ji6AXQ
AGa9WUVyecQkOEe7iqYwYYvZXbght5fWTOhw9Is1o0IJdeA/5DKYMsJMFefq30iR
7kOhR/Fr5ZeCEExYDhUGwh8nFbW9cAFH9ISjgdh85/f8qbwQgQX9T7qfr3Yd/t1V
PzhTte6B0TxwM6B0HVdE0NKpCrqeAQy5V3+1MmytqeC+St15cdMQfGCLrv6PQ3r7
7beshxJJhKYHWorgtXARFYMfhX+0qAVj8an/22AkmmxxB+iyHqhrawgy5fpJ1mhk
yJZ5mohH4Hi4CFSFqaWbJ4573FojcOyKtiks8+1i5ymg+hFposRJCRhLcLyyCHND
shcj/o4YkrhdArqHAjATPe9lsHRBHGU7a+gJ/lVovrNl86REarx44BYe4Sure3No
FgRMojw5uTDgx1qZSV7cSehA4AfKJBG7Mn95NJ0BWltdCBoMUVd8XTqlknGwwirC
x+8G1ElxKoOarP8WQYIuKAOEbgxcOBUHd88dy0UHvPrvJsZrnVbleYALWL/RQkuA
J7MQizcTPSop+7ASsPWeaqUUbdUiFs70vpWpT9erUS9kIvbFkecVpyNylnJHoHyZ
B3wQFMH0RDy5+RfI5qghRLE46H2laXNJ2EQnjLR9ib203ekG2zrHw4UnGR1/VqhR
1minWov6RsPkhcR2N2A6ck+mLin6f0x2dxmspgTGcTHqfr4oh5c4Mt8vQSXHcaeU
jNIRcMEElUU4KMxo8OLxWL3WNyQgSFEExys/eji+JeWVnpOxRr0wYeRrlGuq0naA
LJvuODnTTsxoqAMxicJa8rXwdd9+vZNpkR8NeR8DJnvR2Nu9vfVy5aZlFS+85NQc
wlSCkZDtaWBcoRsmAEkhLvjq7HEH/3DEGS0tvF1xZ7AUVNthkn2D8t7LR3n14oFG
bVSALRs+cFO4c+jpQIrUHwHq96j6zjuaU2eIwnrmnDuLj18UfH49/CuPTQ8ykump
x1UXFseL69nQ7+vJgPR25jBMsV8Hs86DLRK6Z0QnPDOT17eGdbaVsUCYNVDqT1ZA
SNphklvK0RBZFkq7cCuBAVv7VjFz/4LQKGgmjx+oboSFJ5bonLVgc8MXMKjUDA61
EdfAYWiaZ//k2ZpwoW2J5kn7BYKsEGxzn33z4i1w3nzV+QSuO0G95y1L4iivN2Cz
YnyoNsTuB9E8yqV0rj5s/fh1r9cZt9xQJ+hPEroSIvgdd7pFtCUs4B6ysoqBMMlN
QyV42RmqEfb5db+FhsIndXhOncweZw5CBRfrKtu8/txVl6nG3f22nhokUBrdLawT
cl2Naow5Ozj2F0baC65C07Guh3ax7vBEkH3Ks1/m8uP73nmVrL2HVBZXXNTiR3As
AQeh1n3s0jgBth6dpenzgoKkDlbSTQ8qG5WRyv1QLY1PGB4si1aEJJHPuf94tH14
0CYxiVfZU/CnKhq08z4KxjBo01SmYGdPV97Hb1lN2qF9WfXzwiL51mBNSVOtKlrt
otU2zMwyKErDkyJ3PesvYGi/L3BQInJFiWRmZnGGtUjZLWpRV42AbQoF8tzX2fMh
q3wwDewtpVjkGK/Hm7sag9pcG6vo6Og+EwywUWV3ygM5Rif2jaKHDYiXH5Dlv14s
Y4QHf6QfJKYofnPf/A3wycf3hwMHSGkB01/ORfBqO3lIJOYRP+/VSz3Ax0+EfVTP
+2VM9+A9FHr4SVgu8qzsI3KLWSQG6qOo23fkXXuYcsqML/dl2pEvH4kP2o6YPE+5
qX75CzGM6pdsAAtbyVPPfbqyrrmjqHVC0mLn/1/YLLaIxvstNyBEVe5jmPFvTMyg
nOuEG9RvBuwZ5V8E2/pb20IOT0jA2fG2A+SGzIP1pzaoPwhJAaxZTSw79enG/a6k
LQ/Wn4SwexFD4sS83fks4GXnC6X83ejMUf19MthTyImaY3eyeHhmAVOeL+toRHHd
GgU45XWNDXwB9FkAn7PK8NM6bGN6mbE1wfMry+uN+RXVDlMrUzc1GtX0OrlIU3GF
MyHWjN6KhdMfQkpJg0rSjR3IT+/uAr0dyW+JkQE1QCI1bs97i+izrunYVZnjLMZ8
E1dPJgDBSUmHtbzF3czouIC39BUUSSHAavpzxDcmOfDmgaa7jOvcgOP91Dyn7ZBZ
UyU+qvmeMVg0gHvEIzcIEuhgy5nfjkvYI7z4Kz2hUCg63xnXmyv934GO4J32ytmE
THeNKj3Yog69zYsfXT3kB6VBYXPwIHh5GnfYT/c+toKDBzAVEtld+MXIamDylN38
E4PvSa/NCpO84nW+wMhrP/1P7o3dUHaUFf0xY1fe6l+W1IEPW5tN1+qvIldO9h7r
BK989SHbnSdFVqQBPyOVpg4pbhfu4O/Jb0uvvDTY7+sw3V8s9NbyyR4XBBobbrDR
saU9VdhdU9RvQX0OYJh4FzO70QeDhq618dpNNWwQL+1+5Xn4HqLEJHBFzJLQHAjO
EO+hn5rs2hpNInOwdeqqq/PveD1WOKXh9zmiQ+1j5jYo2drcgdqLdFDYjvoQi0WL
WzH7siLjo3keSkpSrr5+0o1l6DZ5H6f0vfxhaoIniBk24u0QIWnhWD1xU5tLjoHl
EvEHDZkoMqWCkAOUX65y0t7+aywlZ2WOAN8UHrSnXiNQBSXPMzk+F3dvP651c6L/
m9trQoLzXVNpkrgDw8bh8mj+0El1AVxEQApRkEZXM0l09Qw1q/2C3faR7DlNlK4S
Hdy8H9/aMcgzo+5FpgYdp4pIA/qgA5A4CoRxvl2AjWMf20G6IPuVORREz56r1cgl
A6X5Q5/94KYhP4ZdNDDpc6nTljCTacxopVmxMwq1G1M5TxfLyXWP4V9SrHdoQDRu
TBx0DTIuxS2VJB2vIS80kHBTqYDy6imSpKt/RjCr/dUpCOhbwMAAjPk5NBottSPH
rDQ6L+cvq7gz4BFCr+0AUEbmL78LzexF88eNZV1HXHSf3ZKRgVJmXlrgGvaaLx+I
0uhICdqPvGx0mq8DzoUyIP+uQBZb1sn730eqTBsmb/J9ObOxtA6sgj8RpxGqt7z9
55cq9hln1/xyMLKcceQq2B4dXVtMXKQgGbeFyIGF9Z6q3W/umE3Z9HDyS1rJpPRn
zJwF6ojmpRbZ82v43ZxRcDGoLfvJ3WkhRKrH5jgc/oNhGgBaNkw47rrhabkZ5dsj
bilzvBxFvX5cdswyQbxgERRkZWPWjD2UGmqWH8ZyXkLIvSewER2iqG74Q3tRhoHG
e6xeXVsxcZxr+IXAFVERtSJYCCZQYaSssWHgbMjlBKiEABJ9GeBZttwe3gpwjYhL
Zsq+ME1tbJX8Xegb8JPz5s5YnX1CBPxFX8pxqA14bUzoTq3RKmvwns3Y0ZoLB6dx
Cz235OLRnqBcvzZ3hu0vWaJi//U3fjifvabsp1Y/Kgo1UVPaszPz4+v1UwDi9zes
7rmUT/bD2cJg/0HZj3wCzHZANDcnQMm7sqZ5X8BLdlKmxogKe6GyxH/RucAg+eu6
5NDoIQTDHaBOUjFUh6xijpurk8JaeRn6GFj6Tgn2PYDWgJQARDijZRSU4QdFs9qo
qHZQx7DMgEKtu4mzJ1JjWQ7zq8UpqewkqYgInhbixSuBaZVY6FNDxU+m3GxAc+Tt
YELo3RFrcAC4ecvbRTXF9t0BJic8C6YA2Yk/HYUjns9i+Y3+Fsi6u0LtBpmu/Tr8
+STYjS/aJJX3HQfKjWBbcABLSD3nzyCCCJE5XquGxEdURRNmjss0URJVCfj+SXuD
CtB3Y8oOVVcegrx8QN7K8px10E8JLECNz8i6BeaE97adec1He5o0PVSXv5yyqPFj
YkgYQNFQtDabHPKLcaERPbMqYD275SIQw4V6Hdv40MJqxYUsL48PjcyITbUIbH2z
OuJLbj7fOJMRYXr1+xxukxAb2a+znKIjbPd4I2nqFmAgWqVs8/LgiZqcNxd/mmAj
57GrgmyxxQeJFy4G2ET+SAP4BcmlXqK3LzDl2IgKOI4G/d9RsKiX2KM4OHLDxy3i
WsHJChjADe9E5a3/tnFv3sfUH/0pey2pbuhcMc+A99xm/jav8mlp1VF2o6lppJcg
MFw5CHPp40xOi99JiPWddzGs+Rof8xS/DXPcV4nS7EaZ0vPTwcEfAPviIzFv3oUs
7UFyiQi/Mi+FUK9hikYN+YflSrorT2Zwk9IjCMS1bXNNMKwSrav/Q26N7C7mDXLT
EjkbFyJmb1M1ZB23e2GG8Mco1MI50R7Bb83SEH/A3fWb3skB7UPNRA15rPiRaftt
U4/QLcyUd0ets7JE/xNJw+8Q49IxC4PlJCstLjCV7q+pdwJMRzOsropHEuk7IZGA
yo5vebbqdaqVoxjdVK6Gb3A3zOfHEiI1/5uax+dgc21f/p/+jRR/j2GuWzWGSnrn
NSVFHNpdZWcwkfS/MAk9M9LjrEmqLAMFSAQiXB5Pq+lQFK2GQaC5pwuJxhADoOiw
6LDaVXJ8YycTsFwIZzJyXb+P6Qou67yyIRrldlzNLW1Vn/dKl3V20VeTjXW5wPEW
clyleyDwMyHCvGgg+vw72ZGR1lkpJ8qgtaDlIWOQyG+GhLrhGCi0kYriGgGFMgum
sOp9bpuWU/QeuIx5fM+Y2+WsJq//0mk8SkenhwqPx+78zShsp6djFFB7/zNoeXBa
M7BK5zpqnbcZY0mK/sl3WKDBpum/NtiSXYxfwtLNiWt/lJCy1PLDCVpUcx6C1SuI
dQjjWtN7xSMBgw3iDRfkjl+vN7Q3jOBcMMR56BMgDRnViqO0HcpRQDCJDTjBTf84
KU55UIeSTVc7NsIPeSqIYnybbY+S4040lNK4xp7oRQLZ7ekjxpOxURcc4KmPCCpl
e4hR9In6ouldo6IpoQorW9j7Tq0ZMJF3bgOxiHKOMI+0wMf/5oFlQoZFkGmxLExf
aeRrEGQRikz+m82Nikiy0tMw/0H/ur5SwjuDbb4YG2JP5NGmyTdPzR8qMLdsijzg
unp4WDhdPaJlbF75N6/fMx8M/0g01rLtU0ajYaATBc3nRjoGtLlpD5jnv2JIz8J2
vldjc1sNUQ2H8wMAhUIRIdCSmzkMNRmXAHU88GUuRCE6Cafb2WCvb3tBdNUbLodJ
vWTAwrx5imisueDsHF4kGGON563dMp/LUX/H5dCJvClozMIgEcN1RP6NbIQUCzXq
w3gOECkK7j2HeM7AV6253SdhBNViA5Br1w9fC6sBNrmcbfndl1JBgzJkPzzN88k4
WtxpZDXKflsIiT2KDgVQYAVzUxE2T3nZ9TV82w/AToCZaoZoIqy38mhhHv0omO1u
IZ9zsQJlwpX0dFK3+JqbNtSAUbV4Ys4LbgQOLxjD+EN3SXRLvL+5K2GRRmSzFpAx
+36oEz417lhx/rC+3V0FxO6MT8fGCbbmXme8uFkjRqNSj1OfgXR6+ky1PTWk4wh4
htxWnM9QEl71wxEI48rmlswG5lhzYm+6D7/mSgm6aNJjbH4Ox1n7uLTma3gQcnMl
U8avP0Qegd2MTww5r+/1O4JCF+df0r/maB5HPpfGqXQtb64qBuH2Fpcmp35uzsbs
Ox08rWWTLnN6Jst6ba2xOYAplivbp1P9fwG8oF4jpvpAhl0L6gUAh0ESndcSJtuf
Z/k48adPGusqsU6NKt8TC3tureoY6nq8t/RBsHku3sAJ3skaC56UAEnah9IKfki9
52PB4YShgFls6rQqfjvQAysEQksWUNGwKMHGabDmdfyQWx7SHJBPu0K7nw3orBZe
ab8+OgU0sPrBhB52QO1gWpYAsgDSZtj1pVT3oRiGOMYZtwUklv9rKjMLqB+FTdCI
iOcwlIx/EQCAFi+Amf7hWKpIpwM86JdMhBJ0/Nz0UcNxLG8gy5h9v89sK/SET3rC
pFNl5ev5Kw7GQ7N1jc3SFZhlR20v+g/9wJYodwphNVMd8rRegWx6714AIT+qG4Qf
eK7ctj/TD8MFtbEleIWXM3JoqBj7dVVolSl4tVyrOGpjo/Jp+SbGmsUhIuUBCOQz
Ckr3usqDyM9HsJzutQfa8qGvQE3yfENt/CgV13GTXCjNQKlY0g2LKNMdHq9dESwh
m4lRJo+0BNvXnka2HbehHxHB4DbeyMpr8csVJpe9rcmaAR6nHhSfI2AMUrKCPWuv
r3E9qLo5N0E6rGkWSXhZpXUzWH+iwG8xHMtUG1CMAbpbHyCoNblFslqsNhuig3P8
AFUmQEsnCZPbC4uBeaKWub6TO+hiwtFUt099gnFNI3QaLifXtB/qMcsE2r4D4rw8
EAPQyODoSI0vthDFzaruM08HX/OQje4aUQgu35Cj2MXdZPg5NBD8we7qx42SkVtJ
O1uXbcGmkgK4RgW3dtfP/uJuFM1AxyvZImJ58VH+RdQXQaJgqO8i5VPOPe0sFtKh
oRFKSgf+aRuR4IxnXH5+OCyawYNuYGvs8SToLuST8k8NecG6MH4ogjy2MQCZ9UKM
MNXkEGDeXi87mPM/Wa0rBhNGf8ctNXot3ZoI0p6B4K9O2BR87BEi60fnFAK91doN
THAL+QxHME7ZZgjFgS9iFdFBp7u1lNd24g78l8MlL/qDv1mJjZV4GMQzePk8UXFX
6TgdZmpy8TvCqU2TzlSX5FHu0o5HJawNmZJ7EKGipNalKq3FdDI38DtVf/X6Hi37
Zrq4u1EOkPXhWz3LIe9payB2DTW+XcZpjXPPHBCgH2QaBaKl0deNNRsNz/fGNPPK
fl4DXG3Qi9fv7iTSheZd5KtTAI9XaA9Z1w08pXmCfBvX5LXHkTjZLM255+vR9hD9
4cp7xI88BO8rNnoa5xBNlUJWXPgFORUGDzHvcTaI/eQflAVr2AnWCUzGkhXHU1k6
CyS9/dq6lDgqMMLCqv9sTXLa6fPCFwq/2oIAQdzF43L/xHcO4iI4FFb5LbCqd92G
OIw3Nzb4n5VwTsTOVRr60EWhtGRMOiVq4Dhre2xEQO7aVvmn7T/LtWe0AXUmEMR4
yEjLnNwN4RlnPeoPpt/GhGuv2SQTPAy7EgiyloHefQ5z0H/AWQ/VV3y+tsWjLl1q
VR0xUibMAoSWz/U0gzQn05LT9leh2chI/oeAiyK1gaknJk4MLbi6AqpY0E4m1+Z5
gN781EsVQD1dgV4ScUmD3VkTAaExR+hIDmSPAe+LFMusvOvKna+KgmIbkCk2QXkT
Bh5TC0sxhudZ7zDzjs7O3fU7Ws6uggtk3QNtMrVKFtX4ltUuzZXbt/SGg7NGQqDQ
CKzbeupBq5DJKT+OCiUgRUGp//rOPKd2ynG9jPrOFDVMKOKFss75Iik3qpnpgJY5
RnrJZOvg3BU1I+J876bIjjAHiaCEaWnmo6vbbfHcoT7kwDAknUmzP9mabqmrW6Dl
7dfgXBIcD5h4p331owoTlaNJaNluODPJCv0OhAqqbffjOAf49J42r5brhv4esjdf
Q6UGUAnIFRk6zrBUTVfpB6gTeSbYohEs7eLm+ypN+/lDJ7be7/KBadVllMyKIhYW
bBZMTW3iMmWHahMKTxyymomAwVz+JDOdcErX0Ri4hu+UIFT3XKDNzVHJ5sUEOK5q
CUJk490b1LIM6OgtMSoaPv7Naw/7dJRg2JCvGMrc7/xYOJjwA/4+dO70QQuUvDyu
3PaEjgMnVY5uyM7DyudlDgwxvT+RVd6hbrzJ1LluPVVURd4y2HimkRq8XMcleQeM
GM9QR1Zwoo43WG33UaaxiBPiCY3aV3FcuAr2zp8SqCNVGTPwHyJZbfmRvmQxe00n
ACoPEbLgZMAZ6ZPstm/laEGF3FoStRvRrUqcZgv7fpKKLvsnkFY/uJ2bvRqXg4QZ
hEXaZyi8jUs5ZJ7GOZ2ICRZOm6dFIdT8kaa+ndpGhKw7X430q062rV7v89W7e98r
Ac+1JwjSVPDlZKHaxicobvKNHxwNzg71lPI8huKeBBeUp/2Vvv/g6urxL8qj8fp3
WxSDsqdHKbJqNDwxbVx6n+UyuH/m51jsZu18inOFNeq23Wef0G1PMvL9NLeFpcW/
Y7C3HpHO7FBjuP1S4TsfGX49ZUzxnxqZKsWmNit4uoOwqs+71f56ti9XkmZJkPLT
J5Cg9Hl97ThDYBBXFkEzEsfNehs+T2CkqAQYbLjN3RMF2N6QtE210hlQSyazKmhz
1+X+3MxGF1QIpAOL6EvOoRPN5U0qS/DwHJCf/40w2KkfsfAKZWXeU/QSoLYkE4Hz
wRAy7XV0Ek2L3+7LUmJvEQXOKAwK/PmxCYTTUsOHLfU/gbR/elrylFsSDPYiZm3G
bRahzYuC+b3PdtCZpx6zDwDbVkxileqzfD/6Bkj/PVf/e3bP4Aa+rRSqLQG8qbL0
4NC4s78YYF7iae+sBroqFlNI1IjkbKrdXbFbKqYhIMIe7nciuxfDgABnOUS8nYVk
crYmdSlx5TiftImL65AGtFlR9XeVvUBEuUg1nPf2ATxRP0kzc8KNrL+umsW2l+TU
21vvdO6RLBugQnsbYouOBMIWP/FZUjVOjgwoLksP407SJoyjEThLz7/sLtNRvmOl
rFbRCqM5ddNVzQUsIJ5uBbZ/8+l3MG8p7yx9P0SItkUrI0QwYagvqkm1l0LpYl85
xxdw6btW0wFyJpfDOc0Bu8WgSu74ivLVnm9x1aJtqhHpDJfMgRUldbrbOYfutCTz
RvGZoNhhaNy6tlUC/nTjBC11jsj1gCJvRM7gsn2krQLPmFKL0g22i6ffAE/OO8Vb
wN0Tr2yNVoVbgFvWmd8j1xoly7fStmt9j25njeor26lGQRF91ET6uVtPo17C5/PL
eFOszvJNu0DAN7pAsRL3jIK835nvKJelOxba9yA2W8RZBRXy80uTvwq3f8cZMotI
MPG2CpNlgiNnTAjJP8RJ0R/nDS0Wf2ydu19X/9Nm0HUhU1Rq7gl2nIV/hLPWcaxs
UqauHcVqgQf5gapFtQP7gcg4/tZtjHZQueXOIaLP1cBEnRcmmCUZYc5WZVXME4F7
jGPcT2Vuo2tedn3+W47WzkOmrp6NEVWeo7aSsubAbqx4OPL6NRmMpQwxmUcteZja
94957bzGPviqj/NITVPpNKpp5E3khNPRRuSy5xDY+1UzARJHgjG27ea/ARJZku7H
d/a7eHcli9O9LVlt0VCDzpo2GBzzuTMe1PMulnJjvciliKtRtEGI4YGNNDGlQh2D
zKJIdnkD3ltO6aHyQHtp4tSFesmDxhkE+9XtZEOZ1beTpHIwGbss5ihCVlMNdFqB
eoZfr52bChpyblB51TxB/nlPU5bwenoyqjscdE9UE38yo4G6r9Mibvb+I7s6g/tO
hVBNLJFwaNSFlgkTQXkXzU1LlaXy99A6csIjLffiE+kEjvMQskkCiGHv4cpNJwwF
aezjxEkVI8F/PHR1DdHAC2bzz7i36roXh9hOlB/Zhyae171/iv77n5JU+04Ifld0
UfpPpXWBKzNsgHiPZA/uRSEBMv5zLO82nyZXDW6KU3IlncyfdZkWIVryv/8OED89
AIcXwCf2T5QkaUH9aOi7FhMbJKFeGCj8zD/JrxO/fvYAFieYQtGdFEvV8tg1cIfH
EBY1YzeTahO1P0Za1nWbiMF4xB+/KHbADgIGbq4vMPsOEO/JZfG3FSNyd3R1Vsds
ijOLhFmN+klLbH8p77R9rk1GdRJoF7NUFtcrWWMdNTnhxKX9UK1n+M6l5oZ3fr53
qkeY5kld8b1AaWeUDsQnuUqU3qxo3UaQy1JwzkKsz4luM8Trd3ZVsL5j5y9goUUc
zCpQOnQoDwJ2E+DcCOrSqgXaD88nWKJNXXNMCCvUfFca1hEVbkCggocJsczZru+i
QI552uB33h3QmJqLW0PSTdeo9YbEcGxLeSSgZb2ILX3Oda2tap+XcyZ52UhxVFLQ
Ex2KFOPRR2lKJCM+oHyl3EHMT0SMM8vr7nz6dwwz9LIw3zOSJqSKJMKcDgakMIVp
k19pvuLwjPWC0dEst6OLP3oqC+8qVooSoDi+YR3RB65VHfWeKJUd+4qhh/mxr+zs
k3Iv9iMAs4rG0wFfecR1H4z+euokeAOqVQJh+i/vMqslbpjMO6U3O63thpAd1NfF
vQJ3bNwwPTXg11bZk2bhz+XAMf0TuOTE3p/iWdUMgoPQ7Op8IH/1AcydsERMZ7VP
qvftuHkiMzSaZFJhXY+eQsdoE+DEJhIJj8oLDQWjXbf7OLbHBvG17dsZIuSz2oXE
YM3xoWaAXf6IStw1oXxFkftm41P47wV71OY4W/nw2YrHjDnYIzw5OeE5WjOIZwuh
MsAG1kv2dCiqTbfy0Hr7/JxndIFKeqqcHckYxDj3ve4H5FBTd8KJtf4Lx0sHS4TS
7rcEWLUu4o5xsGu5G9aMCeVm9aY3BTi6KgUEnzzFtiT8zOMrvPQI8nQ3nW0rTh/5
K321ax0QhGmVdlxv78CGO/3SbAtPuklLcGr+zZWVOynPV14j2mRfs5IDhcvDP53f
HyXkzIFBwzW1CCzxdwzgMw5FeeNGWHQegNFhc34mnDjNxLvFL0B5I+1it2G/vAQq
TbpOPiGHrp+bOpaiyP8FaF6x3h1CE0YD7KLG0MTrRe08tOVP5jss6W9I1xgwuBLO
+fKTBHeJk88BozEskqDj+Acx/2ZCRvLVn1Gh9MQiGoYWuMsIu/0eez1k25mgof5D
rO+KfZnx7mFyTz53gOz/VLUsGgd00QZkOXQn9SsRsQMrxPw4gDJNZm6pj8GIFSbD
qmBV6byYt51OUp0VL1eXnUOfAmM8gAP3ttuN6P0qVxXBRUyNZc5mndzQkS7B52U1
CVw+WCeHYD+4VA5uggtsDx0/xoDNYbXPoKcwidy7Scg40bbAd6aK6vcFPogicuix
g+/X6y+ywCz7cGBrWt7gWb/ccJYP2aKW2irGhCHwwIQZUblL2QWAwGK9rRkQj4sq
QSr6738jt1f/AwuQ9lNO0kmv/sEbQsyb9Q2sWpslRA7o73bJOLLcGtvvIJRM8mAP
FrkvKcsiqcJ+/FAGugFMZRaEUm0tTPxAP4R/dhojtOa8RwD0vSJ4j/66tsbHJlv2
eGfLm0+KJsfvjaJNiqiU8ZenIG/PzHDHXLAF/RIBUB2jGzsguRUtxXo5si9j0LnS
DA5bL8/1q2gorOKDbNKalrglZ0bYXh1BQWL7HxJrzzqdgnyEBbP8P4n/RPFmIUID
9eHX/nVvQYAlnephSZ5s8gUqPd0uvKXaZqbJJAxjGBLi8CKWmQIVCaqDWs+3Ctg5
9RdE0qpHURyO9H/p+zmF0rbrWGTUg91hf0WuKI83jf8M03ZAetcIQ+lqAI6vPUjD
d9yDulYZgk9/jFkp9+5hDPjNlmj6H4LuGVjnWjN9evMtIjBsZqYnNas/cs8dc3Aq
CIrJw9ELBn5sRhn7mfQdK9nEWE4jIBl3keh3cmuFZUb0NzfPgDuyKsEd/a3acqpl
X4Dahq8GFPaq7zjVgXAMc6j5jGQj3bYGyQVWaNrCE7+AxoiYmafjv0KH+BvXHITP
aFuhpO5WEloyK4FaPO/l2rS2irFgy93guZtn5p+TuvGqaDTdpXlUutQqksqjcgwo
YD8L93MyB5kxyxlW7oBXuWmpL0S1NnTXkCmsbDuNOKUe4VT9Qvhzq5j7lk7W9MHy
kqLGM05GcDKy8FoVu2x/IyyRkMScBLFm8zl+rHqnwp7qvfonfThccjXfgiN7peBf
XxD8Mcb/VHAlxAHlQOSmeZDALj5X9jV++D/Ek1ozFQ6aeiu+9lbjQwBxS9ciVzoe
s4fy5pOUgFWoe1sg/uDlXtI5GzpNnFjRBUHaEHBqVLjv2615MP/V4fDXKHtSN6hd
ZTsUlZOziVe9rV1RJAFun3zk0cqCPUJqQvEuoDv2/3EQOdHEUnBEyQkS4UHKACpx
aNmQQvGfy9FnyBDeioWdaR/6PvxxPtvMTBwsK5up9GaPbSwCujg7ZeVmHaeSI+7J
lDO2UuoTyJA4NY517UoSb1dT15v0F7DFAK0QExzfzEUDRdb2Sn45DyNg94Sika7x
kCrCBwFDBtg11ppn8pYALDwzmgWy8EEoDYp7s/tXym5mgIPuZSsu/qyOQffGQfcN
+KjQWSqxQDBmSNge3exvaVPUx6plyqheheT84MI/e2bjK6OoukWPIBvZ0ozcxomg
NN643W/6s0Kruyd4XDT9Zi7ZDtTLlGEuHFClbfP1Np6d0xexGcQqthkJirdf7Uu+
LY8+KGzjJgF8MZgmh1LNR99MOTJhicWGA3qE0yRDB0GLWBuv5nSz0F9n8p8nSR/i
DfuPbNy2Mc/5zZ//eIXBefzpDECwyu203iNc2TcmdimVg2iAScgBHmDks1ydS0pg
y8i/vOBvUSGRae0WmtGRE0R8/AaBojs7rlh6uSaz2Gf9fOJ/qKuoat35AhvoVPRT
GchPUOuZqjziNyhl9cu3HaVFXHipSBV9LQGt7K+273UH7xo+5h2DbERPKAL0f7EI
CKTnJ+nGTj/vg+F6M6VKO/VLcGdAvrWmHXqH4wSgMs48gC35F8p5aeUlcFSqVZ+n
Zhti07eSCO0937/rw+Wdl3FEgvYUPncUiGfKbH7pdJZq92s1olE9644grSYrP2rQ
EvwL4+I1bORd4QOqtYkqiO3RGy+mrwGJQZeq7tDO3hz7DXLRkgWZfHV1Ns4ip4zy
le5hVnQlgJXPI95y9YnFRTgpRhqrhXVMEUzw1p9g1v4TG4En57OFlml1V/3ZndQQ
fdQANyf0AHIshpBwWznpVSY/9gciSgA9OWdUw4oHxbmAWl5sy0vE74tVG6GADNZ4
ChDii9kRI1xDFheC6v0z4gwTtzBe+3yh0FNRR7If47kD0iNbVHosOvZxN5v1vXoE
HkkQrPK0ecEj7uVXlOt/xnKECVJhFrrX/SMJzTzDBKniZfdtVLwuVG0X43zi1eDO
EFZmk4Is5Y609Yaj559FOqkGveMKVs3t2nh1mVCdu3az9jR8v3WaLpMMy3PKApnM
9DrX7b19tCSJSE7OQlnjtaucM5UiM7c78aL8BY7xpwJ7KDc1Od6sdb1TtFHF91wL
itdCVhhQk96X0Rw/NrIybN8cTc7HAoISyQVjiWUq+Gj2MI6hFZKg6xgkjLa+L7yD
nLrAMNjOsWRZCkux1n/o2/LIcToUEWI00dkWb6IcqGZUrkn9EOvLEiFVrL7mWjSm
/PDN0WokgyUgnvpBtAW67qMdQy7NLC8Wcwp/hHIzUmBb3wSB7uNlaiBIqKetI3um
uUeZj3P2n4i/rmqgM3ZwSv5ibfysPkxFW9IjMg6US6nOlTexjBA8iWS56cnU76T2
TpSJJ9ofSVTd6NuTG+nXL5coCjLznl/u+y5f/UrFtRnWqx+7mccKr3bqnrc4tsS9
vEzmUYYyKIlnZHBnK2guihUxh3CnFHxzviSG4Ef+0p9h2NesaLkyLymfJ0YQjyc6
HYyCJz98PpwVX7xB/b6o9RtJM2DqcI83iBi33YqeagK4KP4gXjd2eYXPiKFzdCs8
Q64vc9cPjRzRFMras+wF9tm4gMXsPRu3fA87q/hh63LYDcsyp/qXmV7cAAPCw2aU
CZms8xJXaZj5Xl1/MN7YdRwUubLzNC23LdxC4bTY6xf7iSb9rlJkZnDbLtfphpZE
jpv0+CsRXAOnWHlF77W8DuUlWZdDp2B+j8wp6hpccDGkds2a1IUbHCVfmHsf7Z9t
6ZLVtw8WJUsbO/zcLJiXrglHWqmdmzKPjg/W+pRpk/4mwzEkPWMcjp/IeNlxrPKL
pN8Hr0rzsxHL+lfrivCB/UcS+NBcdJzIjZt3Qejx+2mLL0u0OSuVGuC+6ncRwdMe
x1Ng74tpjCZTZrhgKDowLJ5Ve6JSZYm6hljBvbJg43DECADM0IGSwqLKVf33H1P9
/VXVEwOGFYHHkj46g0OE/Hcz4QW1Q2CLDV+v83Xe3vhgggQZ4SNMCmt4nE2usmAg
1+6lZLD39Nt5sk3cXcUUeTdyrqgbgpX/G5SI1It35gQRdZK8b4U/2WnDTls2BBD6
JibLU6Pqlk2mwlwBdx9J7UE+3LkyScrTqkR1z7HYETfc8UxqbTVxKgU8cOgKcZ9C
H7W6+WvIQMVD8lwCYQdCKkQjlj7OpcvnjZCO3LLtcqcNjJQ5aKRic/cYIlYp9YWg
UrTdJHThVkgSXSNh+trOqb3cMaoq4ZQUaJDjuw/wg5AP9aCLR5UpItVAxSX0X2e7
6kK8ESR9QnWFBvrD9GhvSQd/uDqbMSilYViQoNPQjGkeThoeQvvrNL7dBcbFUeDR
Tcwf/atXtKtYOqSzzZbbXW5j5u/SqRKiPCcfk2Myo13jArdxuBki9Avy0OVihDCc
d5ndGYWtKaJ4royKnBQBbDJP2+G4bwZEeza25H4IzXGyabAubcRrETolZ8oavmMQ
RUNE+Ypt/L87rqYGDPWPX7zsbdbIBPmB5uifRizPUQ3wWXrDh43L7BPKByO0tIuV
419fBbSYzAGKrE/RlO8ed8wYf7+dLE4QOsnKo1T4KuFB834ceohr26oE3bTeEdJE
TnV2eOjNIrDr/HH37CHsY7C/gbL7GDtR6KN4s0QPcb7W6XGqrG/r7u4SQLDfFXXn
CyILj/QIu/+oubBqczFipvvkLA3tGBTofjAnBqEFtHrclXY1/cwOTKGF/9SG6SxK
Rr9UhpM+44iOUSVmLGSHJB1YY6rsz9Kz/QSTQqrrmjxyQ4mhDhw+NTsmdIzvv6JQ
nHR27ug3Ap+fYh0S5d/jOtuC1akpo3uJSbQXVNqagr8VsjQzn0JtQIsPT22ptV3g
DvHHDOwWnLuEKlmi2dKFVRDAkydCG3DM4I9CcdptPooq+IX6MYPaD0+5qjKaY2Ps
9YL81UzUL5mpvmUnoMVbaFcP3Fnq9OAhO/ekoyjMKn1lVr3MdFPgjjtIR60Vkqz+
PqaqM+l8QS9mx9ala9tNa5siO3YZNMm77EkF4aLKC3Ywz+Jx55InOADppHHZQ40Z
xpcr/owywLimSQEeg6/Ggte8yr16WvAGbM9WS8QDHJs3T4j+HQh4dbht+0/BChX7
mrvirvtkquRkJU/kRY88J4AGCSkP7rnVMTTpYPuOqROUl2KVNl+gWYFe6TLgjddG
g4hX1/rM/gTchHORkh4v0eeFpqjkKZ0XIfPRBipFPu/rxcDZxqeEseAd7niF732q
OtBQGscZovNiLjRtOBYjz/ni/Iu0sJbPIO38iLoYjprER0iCQwLOw+H9M46WaOyI
56HMpru14rNo9qttKfz2LqEqZiNzTab/D5gOgHC4Wi/j9jRlzlfrrphCIpLwmHcD
U9SksYiLBDVDAzgSNhfKLlYqXnAyG1Ith3/FOASR8M5wFCT7qBPXnBU0t90UGjvl
U79q7F8rHJW/up3nXO888ikj7MppCDJLi+rLfvCqUDE2MvN/QMe2T3X5KM8VOz3c
uWec5X0A5HDFJ3AVxSHODUpyuG3mNX/PFkyTUVsnIFI0K+piGdBqQXOetMK2uJ/v
l/gcpRr2L1sGGDbT1fsdL681McVqyplfyLpLxyApJZQhja3voaUeA19s2w/J/Hzt
CCoKOjrcSGzpfhslYQpf5FatzFILG0hXkQg79uMXdtnYX+dRFj9RALZtAmKv/mC1
IgylU93oTLIv3v332qUzAKxWvCXl+9mmlFMPlKWU9nRVXDSlSswxFdh/hdBfDKRM
jJcdYvTndVq+jFWwO67Xt+8W8DdQgVBKH5f3V8PUHyc5qil0l8hBF5F40cY82ku/
WNd4pjnowNlMKe2KdP1LPiTIDcDJCnrFYcvV+iq3YVkMgMg2AxPTa0rAsa5/R73K
mxAjozPa7x2JvqEg4lhXVISvDXQVLovdxOT4F+E8Zc9pMuF1Ykm/7PZAbbUYTigy
UsoJQx96ozwGD1voyZecW0Y8UHAJpu8Fr6srlLw8TK7H8TFynXuUxypg4NpaRVL6
KSm6jcBXmc2xFBpYvRiBZiHRsueuij3JnNLuB8354GT0TE1dO4DFSEo7LVuJAcIP
vNUhyM3P2m/Bf5Q0SLa7HSENsw8sv7qfspJCoGbNGd2BsireoBiWOFa+Qt0GIrvv
2A5lkR6a0wFr8u0gd7OuzjvLXx9VEcQkecVpJ0JAP3JXc2VUja+R5jtC/gowJB8J
B32oHpp1A3WyDIQaA/I1kNIV1lLCZTNB+57W/cih4Tu0jSF8TJILbQG+SmlRm9iS
BndmpknPlj8UzaKyaaCcqXJVNF2d0Z5DbRdbut2q3wcvXt64ybFJTSpPkEISgUHO
53eHiHQZHakMBk4NM62rt8wZh5rMHc1Iw7sgRF+bDFvulKRqLQMP00LWpGNfl82I
ZNVTk0c5bt8PVZKVrZMoUyQ8GR4yVu8aM8wXfNApQTv3Ge9bRNDWXz7CCx6hKK5e
dr3kHRfKtbfZ4gIKYcO715YVFJit6vwZzQprQzTsR76k0HcJTO/W1dpO7V4ttd8G
34gebevVK9LPy8BaSzWolAkNA3tCE2KXX2RzMQTyRNspjIKb3etq3A/9ciC0YGYj
+Kg/5yZSHld3iM2eipKoyhc1DVi4YT0UM94varWgusGtsy8SgkYBVmkKI7Mamphz
Vjfjsg/PETzb6vLr9jZTtR4GTBZvsrbtM0A49bU69srJoOzdzc16Plh7LJ1gFtM9
MFluJurvwMVK8bsH/3ZIAsPpAvm3vBuufLGk1cRJurwNNdQ8feC53itX1zieL9A6
qzd3XKRcuWZhvd64I5+WhrgjTJfG8MXAXnREygFKI87U/UV5PFD98LfMishGe2KJ
fic2ar7KPVtKM3nqTg8/tjXKGYuozaa02Ahh0U9Ftw1dFXc8dbPQ8weknSPzdYVC
8HQXXeMm8pNTRUK5r0qC3Y488VaUNX+18nHuKuy/niSUNYEL7Jg23BDf6qRCx1Je
ECvPXFoAjafR+f34F9FfdmX7c8qNWk4LH3nf8yB5Ry8zWr3krMeWEtNkedktySRW
u/AFnv+RpMRXtZVyCPQKmOhIQab4sGoy0HBrE+BArJpZojjQATZWtxH0IthNNucw
4fTDu+HUvy5mJx9f4aaiamKT1aoCTPSGKB++DfONXeyv2e4n959oZmKETpQu6c1G
V0s35gLq3mWefxpxRnmjIA3CJB15kv8Uy1lV3UGdvD9ev2ZviG0LXhR+pguYsHko
7bY4+IVHJJsXI1P3MaBSaSWX7NLphl8/fkWYw6NMKD2X6lHBvaFWkAjXytJxDNfE
mWzVLZqcWH7Wyy3CavbZDIC50xaNBbqQhwoYhKDSlKiHIX8EfAvLqiuWvDM2w+BH
ckUv2lbUBY/4kmEKvNDK8RaUFKZGhynwq8RN3dkmdKDwBJuPjZm8dfgOyV2ieSVa
2al236mekScAuIzlowBjHY2rGwYrlcXyNQgxVf+SlBVZIGOIwPn/93j14BeXDI4H
bKrYxJahIsZIDVyjkfByhAJuUGZ7kkle7REmqjTHBV5dsjeIzEcMC1K2tB9bY1lu
m9uN4kOxufOmIJY5zP2Hcg43uxHSTAacg5N22zDfNnR1MArB/tnXY88iUOPL+mUH
+q6zw1vjPp7COB7LboFOScHlK9SW11JLYxvUMtt6lAXxjRn1jx7lI0+qbvOEtCaO
SY2+jJb5f2TcPHBNa8Zlg1PnKpebQFcbtfR931EMNAxtB7L+jbQzLh6xZWLkXTgK
CWFmP8YuqCJoxriqzNcrNPpXlcnDjg2VTLOlCv74e29+FNp3rszX1OR992fQyxv8
iBUwQBXd3bglzWkNOECaypqvOG1lsCHKeGr+jhThGsY0Q6TVvokzFpBQS4iomjQW
7ANf7SiAbM2ilCqtH4FmS/1z/pUmnLU+rLVGYbBu+JVEUoonmZ3nz59TL52GpAWP
Ilh2+eCSj+ge1cFbegdHS37OiyaHGHWBBGKQfSfLYaTQB5hhg50Wsjf99Lb0pQu+
myh8F4uOBacD2M4lI89+4S5hhejmnJSb69BljD34Uzb1vAhnPjB/F/3G74Ugzc5p
9aMYYyOP2XrZ9wYp1uCfe45jtCvpb3rLu1Us3w7jQW3DZE+/bBrjUYvM0vHjYmLZ
QkSsjjkl8wjY1Jox0PSgKAqut8wCTljnXayMlfgmpIRbUGnI2ZVybkGQzHbSdJwx
zS0QylKrAtB9kh99da4CxeWyDORnDketmGFc2+qx2cAPzMeNo1ohCxpzBmipPJQ2
dxuD5mjS4ymI5SmjeRLZmljQg7K5pqdHuZjwYqCk13MI6vfY/T6ge4wbJQaqAcMC
HPdyjvafyABoyvlw6jgtwQ7RA6a0u0IoBokFUlGl0pYQt2DkTCxCFvmnhiKm0KO9
qzVkjydJZoRZRbVVisbk7wEglTLNlSDFeIphsKkhpLN5nW0fdnSQOSjc5Y0ZqFlD
z1jNz3xM+buqPGB9bFOAPMnOGvpt7CJRBbAQfbUttgTkkx0mcCdLXySDi6ujxKHM
agePgOOrDWmkIkTA9a1kuq177LxRuBEJnQFyi4zWbyDrpMGr07KxBr+7HNl790CB
gQYu5yLHa1ssB6Jr7nRg4TylmQsnNY8fkWo1HzzoyyD3qClm/9PgxKlYhuIsHfdH
6hdnGAgs7+7yALUhFpelcBw5YMIdMPwbyGmkt99R+1sCC1i52jT14i+mrOeAFDQ3
VONr0nj4kunRCv7nMiZxXFUzYYW9SmQamMWUKvrprKc0onUypMkypUGFfnKTQc9K
o9+ImF72ze3fMOa8PjHgpZhr06CBPgHFyhQSHwOOf+kgXPzKH2wOyS62IweIZmgD
EIIDWpvPfd98cU6iiDvZRerV8LA91s56PvhLxiV+b3Di1UmU+ZuiQX3H7+ApCAtG
QUtUEbnAmyh1kM9k8cvYWjdya/bVyGHN6dvdHN75I9wiDQ7xEmjoVIFx0cquksV/
gKXlNwDnx1vrDiGge8lpjQMPZjZtlSA8w64lK+j2fDZhL6B4mTdukgE7iVXmj5uT
4Ff1DJCQsCr9XIe8GJqRZgjYVYH5RywAxy6lJ9V64SfaZDnEHCrhYeqcGeuXTz3a
csRTmshHclSAY+35le1+FXaUzQ4JxkSKlJhOt6/28FwcK3hLSFXZGk4IzxVq1nh1
RCXwt2q6TyEya+T4zDoVTGx0zqODpHw5w48/e5TMfDeuwLcxNdDrJXcxfZT4zuxt
Mqn9ZXaaowliE+HJ8Qm1IS80XeC9r7cEy04iZVwmVz2h7RIahnlOUDJG8ZC4CPA1
tiJlpA5bnC3xPrKvUYa/U1Vwe7qFjDJHpMBR+yJYCZHg7RxzDBtO7PANY539q8he
nR2pxzvOHWzRgiZegzA97ksYT49MNMzx3vr/XBcGJJRK7Xzt4zHiQsYpN0AqAdzU
dGn7Dx2K/D1jt3xk5R6kJgSnpMIbCyAiSMye9mu8FvqGmm/AmbAXBDfCAThTOXE6
3n/QdjEUy4F8lHwkIESNoa1hyLXcCv3ZsqcjBBBLha9n2EaQcoeU3fgkTUEeJk0+
BeV311b5kIleV+geoByKto0gS8Ttb591g/lGl5Nx+rD4x+/jV1VyRGFGOtSuNiqA
lXGEzGDgEqBrPoRy9IQs0Wo8+Jj1F2v85mI/3kpZDRb/9/ApRDhUwnpG/kdy9qz2
/X0VCNoCZuim2kElvvj9kwmmiPGblchw1ZxPHWnFhvguBheR80Pl4CYh33AKYSFs
0V42Q63MBXeO7sk2qaXnVPrDjTgQAVNpbNZcu9rvzJLCyn+wKBF1hhPxCsgsFkyE
IQu++cUvh6xquDuIctdENvbqs04wB4yidWttCRdVJU7ibB+0HutfppiDDx62OzLz
F2Hzd/NPidoydvUrfYXqwwkFXR8EwmZoGG+eOBdta9zY3vqDCtAxP/dWH7W1WRZo
y8aSyIzuQzFuOepdqtmw9lV83xwCayv3OSaabrpC9aDAlR5neUJMXOctdJqRY/qk
aV8DFpR/z/IaRmYrTvTdsTK0+MzdNHSfZsvuRbMXGDNnh3eqT3lS7+xr/5hjppYc
w5ctE4LU3TLXgnr7O84c/gKHR4qpHzy38SDFT1kJVyiQDL1NnV3zpFtUCZGQL1Tg
iUfDUfc37m0GHiKzAaghUO06s2Fdt0UVT3WAHpZokUp8tpsAJqfrpkzPhpkgJDo7
Pjnc97K26aKZhoTKl01ucQ98Ts38jILGsacNGsjCEC4J7wug+FQCJN9OQt0Fum/I
A2yiSHuBKyWTmqafW1//kkH+is5vFM+Ivl+hzLZOyf1xWqRB1Vp8FubqWbpAPGNd
v7W+uS3P8hGNkWqnVsNsTgK5tYuBmvnJpgPFzJ+61WdcDn3f+85VtWAur46O2lMW
Vw+G+yrXmCh5L+3p20NU5JLUDN58PFNPaJ2bsC/6IxRCWyoWsaGoj/3iqGiMB4QR
7cO91F67VU+jw133MSwPs9YhzHemDtN+uTsHEAPHlpWPFX8+cBWOZqwRwKxd0LPJ
FynDDevJKrv3U9pcqxKHO0TYF5Wcdjcusppr9iaw3y+R46OWDJLcVIThZ78Mvyxo
PTbt+a7wzCg8+nn9MTvTqcv9gNp9QAhGLs0nWZWeT1IM1B5mk3q4SLmBOWRUBdY5
9ifsSw/n2jzHGnjiRSMhgrJiICxelw7NDdvBEdsZIA9O3s900M62Dn/yNdpHd59r
6gT6td2YDVLH244NKgAnMMOpI47n7k5OIfFqF1V/druR6aQ6tc7ABXq1uQz0qcOb
IucAg77xcfEoM0zFa5BlySgWgtAewo0hso1zD52uvjpDc8dkkJ+X1/rTl5v6tW7e
9ynfw2sBbjUN1iWfkYB4rnVfO7bVxZuVYwtL//d/XcL9ZjsCKPYE4yedA5z5LoPO
MFBb7DNF+xWauVZJNsBQGsLvZQD9xHqx+w+7dS+useo4SXPndw12W0VQ9KaKNz3P
E6ZZMhK+UyUspE28WNhK7JcyoqRGyEY+183Kz2PPHSVllVtnmRAregeSsg5JknP5
Ix7uaLFpuZHMFPwhEVNa4LR33br/yCOWwWRY8WzPTnv9NGqFWW9TBmBMupQzX2Im
0hiSS4CZ46t9Fqz/dTiqfxLKgHesN1gSRyZtM9+U50EG08p/JMI6nDCXmR6NjYo+
5vgGXSyHbjXB+rmrU1keYxoc016ovHXG7Wg7bdoSfJC7sXzMFW8rMnTo+wDPKTb2
2WMrLHdGc3HTrrw6Zia96MCdjSkoc+moPHRl1XPi9tG3OnUv/NsW81ikimcxD5hs
JgkC7AkDBkXcaub6CovrMEV+EDG19ix5UEOFdQmT1ISxZS7T1HuewfLf2T18IiwC
JCvwm3iJIV57wGt/f1wIvco7JAdyEP+XFuwwK53vfSXLGxuPGAEACoNy4Bunps79
hr4PoDF9UYcgWp6cjCb6vwc6SIwrRiOeZ4vCUtrpHWILbF5asOsG46Pg9xc4xmJj
rBcZd9JhqzAVpS6aD5E2FzleeWdTvfSD1kDy3B7yoRVYOFm2uF+Zs9YQlBN6tcAW
uZGA4xGCGtEG7OVRPXQzHgLh6GMYdocUggGwgZPcioAq3XLYNEOWJsHxhB8bJKv2
5Sqf+g2IpofQwKOUygWegphQqej9rSY/JFt1bYNwAJNjaiuzrP45mKGhT+A6nXSC
+QpcdRFKFVcqi6022FfaJ0Npnr9DtydjSJL0GSpvToJLoJLVJuFDsbmxXkU2OJZF
W318VWVEZk1YZS2wnIMQce0PPtLSjhpdFd11dxQI/WqcPHFGxOlGeb7+0U3gOSCl
cAR2Eo78QtMLsUlhLSeRP2BCpbL1TcWZBPa9ywxIWNfueGfrnEF1Khi9sebNefou
5M0VfQajGEOQ8ozLYJmHG3kb9Nhpx1Yw/0XX/mG2XcPfCJVIo4BdSMWwrVcJW9Ma
WY7ql8+roItXISbZFmlLDjIFa6AXj0GEH1SBK5dqG0sN152sry0i/ZTSbID4kZFx
1WTOyH7es3cIrD2OKIt8GAfqjl4RoETeq/y/gRAFbdNI60nfFXdQUxGbJctZYTxq
Y/KIEVqPb7UmAjVuEwajOZMPtgeGEcdZ7dz5qa0Ga/LFNAztT7uaRHT1LK+R/rW9
WHSyQJjes7JcclUJNaRdNT/JLkhqzoG9N5FxeUjYVCrJCijF9j2t7llEgO3NG5FO
PLNMP9MKzxXuRbw+6OE3DS0BgpGE14Sg7sljTdbApNe43gru0tPYJv1kpdv5vxCG
S/eIklg5FyCTi5OiXy+vwkxpvJMC5LIpsm3mfDHpMIZO39c07zT4d+pwhLIiMXYh
BuVHqvdwxrxeU7eK+80iVG4m+nm4HAQ1BsqgRPU+AUdVjevSIBOMyldpKDc9Yxmn
BHl9BXsuoGDZpshwNg8KpgcCbdP7ziO8RIzBnmA1Kph+HnEeTDRwCj3vz2FoNK/d
7pzkDaLPo0AEmGcGfolX3KbAs4zWukWIec703+P71ls5sJCCVjP3iJp7mKfFeOfI
YmdFe5OqEdu4Tc7uQKBz0/TRaJ+WAaBxEGPlcAklBljDItGmJrJLEFhQj8NwVs89
Si6OtQ0is4FVFpW3oZpCm5MBa+94DqmDWidKK6jiyLHP9Gnd7OJ6gjCEXsVLlf75
sg576p+gJbS3D68Q3W+WhwQWypEPl8VGAkdKjmsF1IBMx7lP3ecT/U+QgQ9fdhzo
gL4ZAjzQlSX1QoCeK5FpWUfnmpAmmiNHoQizjAHO9vi3eoWlju1D85MIdVR+SDU1
lOYNzcN0NTScdg2KgCbnlHwlXAxxfJ1sErjOJbCbxroecrdq+ZZjdWW97ICNFDuI
dHI8E/NY0I1Mh4hM37LNxMCiQ4kkRTz1aCTyDLoa/3sKoNpCsmg0o4z1mLsSPSNV
gMyPaQXAx9sKKYmAfRM9FDfGjig9gnuHkGnYEpHYch0ImvqP9rllIoxPgEhOGxtR
1HOTmgKml5BdmSdnBxEM64rUGyzD0oJqn2VH3cBMxsBmH7R/9OO3U3sApVhJk47g
BHymOk6u07oFSqDIsLvjfERxEIosls5MWZENfw7m29g5wDBswy4jpWzGKVl7k6xE
zQkCIZskvfpCizU6q6UETvUhHApvlqYyqX7suvCl5meKX0MSb8xwPFgtxsHw01fs
6dY34emFwmZY6HEqhO6DoqJMg9xASI/Fiei3L5Np56lbPmEVkBGfPGnlliH36a/i
Z3ygHcGFt5vpxPuuOPK0rMLSOk+ql15x8ADetjz4d4jnqaI/WnWbaNVPGkazQhtF
zWDnONEK/IlUVpTzpyEuLCde13P7JAiw1rxMZqnmiXvLTU+/M06lgdirjc0203er
6YVHIPr46ZbdlUSKYUAK6PX4zuTdY1RWjoUQWewRkhQSuXimCKdU1jb4GgJwlZGr
bzGKq6dqevBuvgH/Yyxg7oQ09tgPcWgoH66LGx2Ea5my9LJIHw34Lfmg56cHToro
UsLLZKQi3FJXbkog+JFZh9aVmLklaKz+FnTKQOG2dcBG1zVOFFcK0KjgCW/Qjt5K
Yol/IDzzYcfhKZVBGw6jPI2KkggLEv5z8idL78HrvO4sKj5RXOGKwqBUs4uY+4nJ
pli1PKh3hTkfJg4WfZQ1AqLXYPY/1IC0byO6HKc/4sjU871Cj2U8xHBP92DfKSA3
rF6VMxnojGKJmWSjElrIiKEG46j6Rx/wmPqX3wxqmwpn3MwR5o4W4QM3hqyoUUaC
0SnGoj+GK6mWwVfj2q9vc6rJmzF5dHYJvqZaOCWYhojsduia+uTaTbMYKrBhWQhp
hL5GgIH+xafe1+lzAJbIsd8V0HQ35NW7+96uzPyb5y7MMB8y9BI0lf1FvhEpzkhy
mMOujm8ZPcVpX2zCpuKBFcIf8vSGoMio9tWJJNBjeEXG1ZihR1mTSEEoP/CVgYQM
0T9uHTCMW+PxrqvyLzZIsD8gcIOOKKSYjPnG0zwSsAhwnl01IDRo8Rm7DAJnc5e2
M5c687IoXGk/daqoZiCdPl3J0N+GiHbjXG9C/EldxgMtLHgSS0zLTOAhabqLZQ5a
d9vxCHCM/V4MF/C2n1bstoNRRSC1YYayhkx0qYEWKfEq0g4H9Doznm/RajgX6oFT
g2wZxZRCN0k3NrbWbIWgTZdPMWECeOeupwgcMwsaChn8zPRCkvml49EEQel959Xo
esd4ft1xLjudjr+Qyx0FHp68O57hvQMPtWd9bAvAltdxtNEvekPq8+inkoe3SOxt
lOLedG2s0vUR3msShD/O10fTkKK1jDJGEwb+kDWXoyQnwy7cyzgJELJw4+YrVxNe
dthPWhGm6DSJwvsqIxd8Wsj/X+dnntH5KYWx28r61kTKcEFFgledpQm78eCdbCLF
PKUJIgNEsdH6ywHY55qY6XupOC609m0N3I9WBGsbmYGnlXa2lb2/nMGCy3tU59VZ
GZgsAdtgiDG6cIm0/LXZWgl6qr5CqqOujeJWC1XcfI2viBfau5Ng+z0iZjQdB/lB
ym9v7FyZergjGnC0+CNXsqRTbVl4b1hjx2/nY81K8Ttd6k8YSbi4Lg3NLcqFabeL
lfE0PyZW1WPlIcWGDDdofPsgG+ApR3diWm0GXEWzYlkOTF6r6mukI7xd0US+BlrV
irz1Fkhb+YSBcli0FatEibb5P/4VLGi9ctY6jyihjuLCBtEcT4ssx5z4NsVVCYGc
0DvNiqFnk5O8Ue2YBhguSYj3G5mL+RbwRxZfFkvynveITnmkmeK7K1hEzYy4v6oI
9D3GJ768ZWghMDGsKyYJ+UACzzzv37HvRz49fI7xLAW/sA+HZVM2vXBkRqwpyYfx
Kc/7Pmey7HKDkOak6Q2pcGn2PXAGR0EZCNqzKJgJBqCxzDZ9gm0vV3iibrtCCMYO
1z0LCZCQDOKFJgXxUi90FDEIcVumW2VWqH6nEJJnAdcjfTMkYcQDamLVT/3oVHH0
xTYWmZK13hB5xgX5lzzpD85I1RrYYfeMOPVe/l0PTvUMgOEgOy0hsv0Z+wUnaqqE
e+Y8Q/HgKoJ+q5HY8EDXkkbL997v3Gtw1F/WmxGAuP/JP8iEGuvpViPD6QVganOM
Yd30hBoC0m/uVQ8Da7Z564AKq97+mV/JmeIxl74SnAne+dtvDCjwC5bqgy+UO/vF
23X/DJj5KD9XGeE4iKEnVYJsYAsNQPjwy1TOTCjrnXSLfpUEOr9oV6x2TOOzPXNp
3uUBDUakenYKL84Sp0lnlnshkh2oW+zrp/SX0AZDWvHzmComuK5kMaXizU0rk4th
38YrMyyIDOEa6TrrDepkPr13h2JMBBS6OZM2aFIy2V/GwAa656nu6EZnHdKwKfiV
iGyJ9maymUg0dvzShA0wLdhX+e1nljJVy3MXzYA7ZSE7sCFUuhNueLS6lxCazPQu
yK8U82P70ZTsrUP6bqWu/HxXKCO4fF7/lIz4/7vOWTfmpdKMzMuRYR8QNPlnvRvF
XjedtGaQVuz/25VHFcSg+yGEcMCQ96CQP7MV3LO7kgm1j6j3RyEfl4rjNbTHwmcv
YKEWUJP2Q66pV7AXgz3qjcNyUpGy+QrI+Mmyo47m0Wit9Jq8XXq0iN8JAY3QMP5B
ZIwguBJZ9lpLNv7tuyaO+HK4oVBmm9nzbZwpPMj2DIm5C5RWlgfrQjmdTijvDCHp
7BexjnA9ZKWHUmGXL4lydyOgJVUlkLyn+enxRz91RB0BEvDD/HAyLOU7BOknpt4B
k061CM6BXtMuHcwrWpQJ0xeW3ndpAkyt3qN+fdLTsCAG7ucQ69jJyQk4FQDrlIuJ
yS8bhU+sdZ1HQ6eeejAQKXZ3HGpp1+MwW6qDeaNVdz0Xg31SOKd6I99ubs3hpNsl
Ic1AOR9b2zewSz6rBEH4ugpPGJZ5UcqxDl4M3MDgwA2UXiyAWfcJ41eRPj9Q48GE
QvxmlG4cBTR+HY5woE/EUzWZfRbxflpGPDWLkxBQurdqY5V56+c833VHar8ZBVwG
rBo4zLDawuUa08wnrkkFPsm5eVRYzBbd3dmGU1BFpPSA88qseOdbTSL81HsaM5GA
TMXgY5UyXs92UyWSItxVVpYkbjD6qSkhGRJ/xx0YDGJhEN+j4JdQgRSo6RY3GDzG
ppWxx33ssGWh9dIbrTWn8w60pLIw8Vi2UowgciOOaxh0IhIWmq1rStXm5hhpTZYy
xobQW81GSvl7SQpCNYXDFuSKQo6gFjUUatRJVsRtmL2BOdHTuPgK/vRUBnyJhX1G
X9rZq0dRyUcW89cNqvlIs+10nQeXzCe/GfsuFV0SMgFzmYZ9KrrYoKDhRC5vhruv
iRceZXo8j+zFUnD4DZ6XJ4MjtxDSiC9/YZY/9+VZqCU1sR0jcAQY4nE4PS3OxmpS
r1JgsiiIPIdZ/zncX2M8HhR0lYuOWSp5UsrzovzyD3S4datqiLOXJnh6FTPWyJEs
6YDn6C1BA20zPp5kzugyy4PxUx9KHrbTR0o9DXO7vNpbxLAkzc3s2Nv/6mPLCHs/
ICI+lwrxIqpeL4BsoG4ggA96vKMLbsJHwsiQ1LX8xT+p3u4nQpLZrLKOpYHUxUsp
NbrEwxVzhlesTD0RdpHCaY4qYfJnrmYJ6DYJ9ZgH3gfid1Ih2NjZ+RKzc529Om6N
3gYSk67x0IK7Rw4IP/GYf+Yz3Il+BU2gubqz7/dr78e5/GAJIN8QGAaqc8+lyhYO
27a0gXhm38Mnj/8Zygudzv7YJR14PwL6oB4fK7Z1m0W5KvjEcqSDiSaOgS0gNLlJ
uCeuKtlcMk9X/RnMOaxkQhnPnYAB2RVJE+dHdmLn+hxZzRjEEia10uh3Zc5FcWRl
tj5RdKa+tthxWHJRC7St1u6mgqSUqcT8p3MuT0FSemznvXft504q8vPQQXf4vn/Y
+oUh9m43zd+a3FMcgvj7wQt85LEkODylr7IZ751WItiVWJ6z+Ktg3Z7eF22GzbXl
d4KfTCTzU7WbcJk5XDG43NyYcJXsdH5oUsJaFV6uZILQmmaU7PYLefbvZr4bt1le
H+RT7iBtlMFBTxEjkjPaLuibZlhKX8CExDnskciQhV3qDQv3wYpiG1cNODTBZeP+
Ig+ylp42HKo5RQahtSluD86gYhPyr3EyoEWn+IKHyAGh2VUDoZfDrjdqusrIMWYp
UDUsZ1qGMPFVhsjPXF7XGiedqs5X4qU6r6k1ebwUjWAZzWTOvSCUG4Kq+S8rHj4a
n7yd+Biw6Xnxc9JvFWFR/c9aq7Ue8vJ5u896sdmLvLIuSnyj6nEoNn48LLWieyw/
v2pe8em/ZR5WT/2HqrYv9kPeEyGNKxdwdUKLqA7h7xMB1/pvOEo8RrQFmyD89aXp
3AsJYFFeQeNQ5ortjj/NF8V4/j8IpZIManb7odXQFozOpuqWg60jWJhsM/nmMWdX
zvE111Nx675JKuVjC6kYF5oQ3DF9xeZ416CZ2MSStd2jhTglzWM/QAeWW8/huuJi
YjSRqWhsjU0+Z7oS6OROgi4Segc9dC7l+erHSIz8PEN4JjDHqFhXBOZDX7TbsPev
ZzFcDBijTnYVjB6UHmOdMf8IJl68LDID5SyfnUDNZUiSn169+tFN60BuoJl+W4Id
zl2PsNyS/mtWupFlUS7Ad4e4erUzIMKEZ3V6DD8SFOiGSnc5g9w4GhSHQwFvrCXs
NaoAfLHiGbQEHVpGXfj2Pb0V0lVT+UPyMS+xAXUJTcInYY7Y9iryrongREjL+tLO
KdGQuS2SKkL9UkSOYvx88ZR9qV7yGLTTX3xfVYL4KrVkR0NX3NQ+gG7aRtFYA/Nj
P17d548Tg2joZkVVACMZuH/g2DDoYNz0E5fS35RAj20XZJlL8zOW3mQYHVTxC3ks
soNBPuJRQ6GfS6YGNX0VgcbEiT7sKTqA3UlX9lBeMtx6AN49GODR2hAyur0f1M8e
KEN1r5U7UB/cHl55amXC/dj7Xa9ej/x8EDkgVxQS8O/tgu8OzrNUbLttnietMMN7
eVAc7AKifjR2gr0URuACeS3w3acEbV3DQ/clR9yKU+hhJ62inPH53xywkwEW3IZu
yDbX8324KNzMoEwFsadhb1O8zwqA8X+l0izU8Qh9NLEu1SnUxoXIeWv+ftYdI68M
ubIqAhyEDeNKfPvyaXQqLeeaAScvae44XR5IVMDKUboHwrh/BTMAqMcS2yRci59Y
VKD2yxmDqLfTOR2ojGr9F3HK/mny6KZPmc5DBt+SA0wKrG7PEJGvWMSNFMc/L1ec
d9ca2vAFp3x9WGWKhyoO3Zw/+Oj28O0iXlNxQpw0gnSjJZDNqfHvmy+n8495dTHK
1W677yQyct7Od6t4zT7NNuGjKY/LONudEXfLzrc6R6/O/zwUCesg3RsDy+sRqUnY
TxhHKEjYfGTJ6Tps9Cd5bPQC2QLUaUG8R6Sid/hMMSP3grvZ+kiSUGAp/oK8jrmw
FMTKKsIxj12caYSMcYAz8Fi8yYdZeXqhflRiyboeqqVP992jhHaUWjB34Z9ghsB7
x6st3nZj9i+EZjFniKFbo99kKevlUhGza6y/aON0WxY4E1GWf4LUsbCn1CYMuiSm
HOXA3zyuNv9oP4lCeFgC0hDmclE2FLxmnOxEzrZSNIlhZ6juAHhyRT5dsnO3YhAz
vi0rwjNa75LGLeUtXIpRu97Evs4QPAmBoS9B1RaJnIZqeXmIJMREE9dQBc4QkQrN
xDACSHQcR7o3bsOrhJ3lcm4Xp8nrvDB0NszK1pFMkkIJo4Y1iWMa5wx8jya2mkPW
fOu3QlPe3SjS5QqfjZ+CKa6K9l/0ww8L9yrFV43saZz/7n2CIHiNZbr2Mo0Iu+/M
pu0L5xKC4rA5807zDGEHIBOwdysuXmw33gFVzF9zDEjtESZz0cLrlA2lJ5Q/fFGE
oXMvXjtYIVgCIJM/TBBeRG3o9SQAHL+Gu4F+KlXcbxF737gToEOaEBiSzm75mXSQ
v0ZaRHwLisWlfse577DGi4eUSErm5ILJJzfaQ5expYtWD4rp/Olx21a/zGXlZmGy
mlCau58WtbaiwUrypef61FzobGu9SN5TVIXyjklkBO7wDDl4lEtlTfYGn5591T6r
qqGMb4VPfgUKxurVRXl3TRPgX40Q11aHOtXKIQrJIjdd3KSxN4g8p2eHWoteoVKR
7j6wUBijsGvuIqlBbyhzIzEh5fhs/MCS3wu3xUk1GbBYne1GV6EOVuAjcCNbN28b
TfcPkQW+SnJNhbuZdotIUKTWhXonJDPVVxl8SWGeQ/X/OX/O4S3RC1QtbTPpIacg
yW4mE7SJU9z9w/YGTCvHWAExVLMTKOu95OqwZKqHCNDFu8GIcJY8zdEoa2HqgFNi
ITHvE0KePDXows/AyEnPCZsFyzCVITz9xBibDlzU2TNt4DGjyXL3vXrmELETLOzi
6ldAeQ4JRsW/IY4g7RbYSpGuQ0BRlvNwnv6j/3rXY8aEv2ReZ4zScMb/7nuZHS1T
QnrvUe0ty0/qO5HZ9AgAjxzh4aEorrmBPpmKT8SPdpEvur3wP+a2anczQvwz3FQJ
Eyr3QMdXkCjPBWsl8H4wk+/+y5Jij0kLF3XBSer0da8w3h7Ak4EanwEHey8TDYn+
tKsa6342WwLkczxbbb6NIJHvXVuT9CYwrU1PIx/6Ei/80Pf9JHUrAYY4GPjRltxH
P3TgmS11uICdYH09gdOot96nRZyHNTWhhQlHuGRGE5rUsuPt/qPPcZ9dYv13Udqm
t3Z5W/KCmxyIgJ+3tlS8/3A7OnVFHr/RbWwAmVm8IkqZ1V0xnuy5I4xOzeyzZguf
HqyWN97otp148EDkB6Vmewu5dsmuGGlI9zPCECwrklSfbt+T9dfRGR3BNW0mxbLt
TylyOlDLfGpj13wHudN54CRk7BdB/hDuxa4hknh8bD6TW/Kd8wTqW43zk2a3My7M
EBWkNAGzPQ9Gzm+9zq5YLwXShrrDCdPWe719e0JZkjVgSIN7Ruf08I+1OoidBdv9
4PcnfNHY8qo11ae1G1JIgX1lBYgBk1TfBk3R+HoR9I85L1JhhruJyFHyVLDFq+74
/+FBtlI0LqX48Si1f1nbFyBfKnrySo7eEOSGMxqmNxF2co2zvTGVZ1wURSfZ+uXG
gBity98hjRf2k9DYQ6balmI4W27Z6VoO74I0YrrSne5suDM+XoDvWt78AE4nds2p
ocnlLVA/CQSAqElLYtweQqG1jVHrhPm2X1AXRSq9mrS9JRaMduwZT4p/Q5YlDaDW
hwcPAmY9BVCiCnF4b6BhPTI0u1dq/wPFWwcF9B4kY6z9He6/tTYRQmVngIPjYTA+
yP/QR9ULSMkefBmetta1qoSfpJY7n41SYVJZMqxKQ+8MLBwX3rv+3QeYMYU+ivsi
pdQUu6H10zP3BuxLNBrtfTPAJCddplZiVQkaSJ7U0uuAcohAWhhN53uAtqtVA/WC
PpdS3U2+GEFYN5qHN4Qbv65OWzmXjCAl0SocUKfoI1tpSlxgJns4kkKwebHH5+9/
LSXV4HUYJhve4BBtSmuhQZawwJHUoqlz1PKBJ755/PxGvD6jdZ564dFDna3gFylM
e4wC5jmttTp7RM4e+ojD9QS53IdZFQdXlWC3RdB87pCythfOxfKVy8jZ6YQ4mwqN
JhWgkYroOPtjnoqr1jXv9olC0PisJnadoCxOSNpxSLqKjKzOvsFOCNcBGX39dEA+
B640YLaKNbjF2Q7L7VdFZOf+Nhrb1p6bPUdVOG3vNrLiNHYDL/OnhSyw0osr8L6W
DvFufY46GDMC23PssTQSWeO1X0N7hG2I17ThHldh/NxxUJjZkLxRVR9hSHYtlX4m
vDYIPoyeZ3BdqTSBx81OnZ2ZCRZJexw5E0lntjs1bOMt31Dzv54op/kPBkKKe7qE
3ru0eukXrTPtii20HJmg1EfXOOXDiCIP6AB3g9CZb2pkGmqgFVFXOjncx4QFgjRL
ZXyZdyQZr5k1tvi+4AKd00Z2+VFAVSka3dhCl5dNSzzxOPjwjZtMZpQlY1o3Fklc
nu8cznfDhLbiVNLOM3NAVGZx9kZ9P++u4SQPlY6pNSUmpdKWWYdEAQQd2IS7znSj
n3+ablhaanUMUb91w4YAjMsAauCJWwp5s7ntW1byU24W/bYXaIYGxwjZvIaMqGhr
YXXjVHztK++t/8JcCiMvHhuwdnNLRqhUNRRAh9HAdk5fUnjeqiN9mSWioo5q7kVx
zBU4SCiOK27s7EANnjh5/A3ycEQlVxVXVBAHidmkNhzAvc6Ax4qs7looslKoLdDg
DuwNt8iNV6bmSeKnT8OUwT6+2dq8r7XgiKpf/VXVlB+t+weRziy2TOvOXInLVngM
9kEPZ2N0Say8tYtfa+4pj43YdkGjmKw7JshDyyKavYWqYu3Bn6ECn7JjQH+tdHYl
tTGy1TZ/m3aoLdJu30AG7T/Q5GczjHz6ESs32K/yb98DIvplsk/RNmQ7u0CPFcaC
7I27rC4IdhcvSz+l5rC5+kF8j2rvsFLSdcS6cSrTJ/WmfskURwSG/LX6yHXXrwOI
L9wR01mk9b7kc0gXbkWq/4rfKndh4EUR/SGvncFWpFqSKSWM/PKJPHLR3J16v7pk
OpxKuP2sio583h1MEDCZsQkb9+DB6J31ArKFrdcdUx2naFi8Isc9OqFqSz8q7Js9
PS1bM/T+u/BSldFizT1xuuCpVEUrwDFcT8ickRrlcE+Lz75fSZ+fsWmZVR1/JskA
Qp7EnBIvuG7Kcc9jz4x2g1Pz24O3dBOyBUQSh3d6uetYQXJQQ/cBZ4NR+cZsnfVb
ydxoXGt9P1jFDJ5eDcJ4znmH7b2tUWDoo+JHq5G9BHDgLtst6w92lZF3DkG/Zz07
qOIZE6SZTYE5JkCq0CnHcibCC/DbHmN+L/+AbzjfgVYOpNbTSIdMMRMiFCiXoifx
4g84WV2AR7zNLr5J/YRS3OPDj+sVvIVLaUCPmZ2lFG49Q2QNRBU17qLFDGxaMT5a
7ojLDZ/OCs0ds0kaLb+g3iW3uWDy2/K57VosRpE22yDF+67nJapPSNThvBYSJZal
TXKlJp4WOtWPZ5NiBx2Vtwz+2mQ3OM0REudC2IgdskWooqemQu2YE0H8+tWRhhJ1
jVslGfHTOMAVndJWlCifpkCVu73XO0vq7vrvVs7mDGTOFLT0LqTx5j1pMT/ff+aN
K+Krh5IiXkAldaUTuGxO0RSvYeGE2OmFzR5NCy3aviuiI+dA3zSdMDvOQFHkeGrA
oGa0VFCdmzlnMsRH8Rs6xKhGbawT6aXz7J4xHXUPQYJ/2BFjSKNtxjybgzP4/IMx
bvaECTl5i02FOC7z6iR2+iC7lGXumfm+nqOTi5v1yLZ3xmT9BWbo6/+bQrs3kJDO
tmsKNgV1QQDPrkkfAUTILFK9Zn2BuvZI5KYXgR9JDGPoUihvQfZ91y0FZ1oHJFwG
/0cZ5GJYJOo8EKIrgJCWNExG4tT7FDMcMw6+o52uxBY48ADpeNbSCPTWOl93Pcwx
CD4MjzynYpJoXeQqx0O9Pa/HJnmKZAb0voVpLC6lN9cYHqcnhQFU03KrsTGcxTkj
P4mqEbzKftPFxZhpvP9C2VAijTWqjvlfmy+WQ2796pupD3DUBp/RRQPTKwsyD45P
kRPWI5L9/NGMntM5ClX4YXCLlMLS4ww2kzxDYxUohGeJEkhbJUAWITfZxECbz2GU
68NwkrF6zm+2BmWcUp8mV+WLI1gj7q/YOvDyrLAK7XL7afpRDhVnS3UAd1o+5DX3
1xWhzwH4KaZ6TNsbB5yJS0/D2tG7StiQsECxvH5gkdTSDZFHHLkr9zabz/hxq4ZB
fkoe4UrCE64dLQ1lKIg0GwgD8cn0l5HIRVmMIZ3yq8EK9J7+lHCU+0ZE5h6Cwuu/
rxhDU3Scu7+vyQYzeNiZceVqLLk9TnrhBXB8UkhEGkHOlEId3eRXp0aAGFN8s7fH
c/CIbaucH3ITwOe0bS09vCDoRCtactj7YZRv14R47yhHBs1u6J2NLM+gnaF1Pvh3
WOGWE0iqx8CivPBBqqQTH529tEVtkXw6+mcnweBUAZIUAtSzkTyIpY3rEzXKConD
P56l34xy7bAR7wFddloQRsFznpmluV0rrEgsapZbg7V+0cL74kB+9sQBnR5AAsmQ
xQS1oPFY5K3mVYqMxwpEPgUZWYqzXSX0nQH0+mtQ0uf7wivMbOCkBMUWr/lF3adh
ggtx+FM2RW+BgKCnfMwwruD8RPQBH4BEJwMLtSNA0iM6UWVeGWN1/eUGuU7aqcj0
lhJECwkn2z4Xzqx8Rqh1cEElWyDHigutXd9GqjQOUlMiMSZpRD1xrF4Rw0vcaPHi
fZIiRzEIRd1qB2iRYWcm5SwevdzZmqhP9NZ9xR02CDCwfdHaYT+edIZzjnrBm4L7
1op+fp2bctDUyqRSBLGDlg3EqEBr+t5GBSVmW0nGCcUH2RK0zol4yq9LA06zVBNG
S7t1xkeoAnhn4IKxM9EE4wAXDjoXYaWgqYJScPX+xnxRZXtJ9rHZxLfNL1jo2Zl/
NS+P1kyIlC375KqZMypDRouxMFrSu13FkdWV6R3wo3nGCEpuqDpMMxRyl7rgE8xj
jLBoXjXtIHcf5pDto3HjzRPeFSTlOefApls0p+kPdym/H3iWPC/6hIqZVSq7ramy
4R5V5orMYCQqmXnz7P88C5MxNsvoux5fEKL3tq8GMn1C9ZJ3ZiBy0lKxKOI1llop
5Oiv6GU4woWTaQoiOghFwT5G115iOmnKzoaUDMR+9r9iYOyHHmhjN92ofUDx48VH
oR7iyp68fIgBRk3ZWO1QaoEq7DEcSHZFspK75i33aPIr2/Bh47Sa4ef8W9ox98IT
jT8eby0g6NpfHKYcho6KLOnAG+qDs5azu7Y3FAf7aaroTSgFvbkeSv7RnYhWfn73
eQFbXw0s0m/tnvHg1jYw9C+XxGQlNuygD73EQ5Q1NJxI1IpHhIUL62VCMksjwcyt
KQ+9hBfshujz/8KDDZcvjQr6RzxnYBAblb/UsYOoPLItNtcecXUL3PKW7FRSt3E6
RZXE2cUrIBXRgnZkPgUVYZNPPmDD93BMddUzB0NVV2NHuKm5Xa6x6Q/83kvJRGcK
v3UGiNEtUx2Xcvl+8ISAmpzdJ1zyJ4wXk3HLhNDDZJZko19k7G+xu6zMRGmOjPvN
IXrWmgyh88IpeSjINNLN/gJAyNj9NWWizAJf0xz62D4qg0JGWCcvB9omkaADClmw
fsyCpYP/eRlaRIsZS2g89xzuM0C78jJ406ycxS7ufHAN8yprkhfCFEorxGtI3E3k
5zjT7q/Tn0W/R+uzv3EaX8nXfv/kHv/VbNcgLwKDrGRlaJu4QnDXsagS0M87Tv0e
wjAHqGIJXsSCaO+68tj8PAAp/ymU9lV8e9E7zNVsYd02h1QPU5OgDShEM6HXnpyV
TTqUD50m/ewXI5IXSRxzVok+e1lGzGv+r1X6cOX5T123CKqyri2WPEJA+3I/xDW/
4EIraymSuBL+L6/P0CWX7/WpaWpL5Lidg1RxexOxlZObMYm+8caWDfu0H7JkIdoP
oWZbNxAnkUbn/gb0iPwcQdsDA2qFom42bNWDqaXfLJPrKIgsPzMH3oqYwtMt0jqz
V7MtJO2p4DupbhrHhLfgVkjB0nJIKfHcMD89Lgw4i4kU7Al1p67mUsy96s3Xc/OO
TPoV1DE4FretNOPLnb0XoQt0nHl5tmDJ0f7890rw0On+iRczqI5ajc3QUOZerX6F
Zexq0M//qUYq9G0GPyS8k8mXV28DQB5QsZ/H+h1Jvx20F6YuEFzOSlM1IqH8Qgf9
N9V0rGCkk2l3jdl47DkDR83fwekTBtfDrN7KzVs7s31NRHaJ9OUj6mciF3rnG4mM
NA2bcb0UJGEJUQtrTqSCqV5FBwPSElKjI0ynHPG75gGfPnjdi220YGEyNvkDg8uB
6SCNYKG7jGnjLkAoRkf+E2z25Uf9WOtYtdVROZGQBW5IUmnVzkjX9fLI5EAI//21
s2Npqk2/tdn3mAut4YmJ4leqqdf8EwlEkVSR3g0Rh7kW0CXi3ZeAMmz5RZz0kQ0E
JUewppXJJ4BZ7oegff2gtQK6Yq55Yfe4/kwZbOx8nJxTOi9PJdG5HQZrLFAnK4E/
zZ5Y0U0lkE9AXLGbDCSjP/OjFpr3c8IGDDioX2OVkkGVV6x6u02myVCz8NJcy90m
/XRCGFfdzyib6CeNydrYGEAntkbQSuv5J6sRe6c/uNTOTnb+mPl2Eio89qA6fZvV
VFx/pWbpB7YlDp/M+9Pi1H6u3lw+ZtUFaLRVV1i72F+2AH8OPN3cTGNE3io6ZywP
F14oWsqgcl2+8lCYtuPmzmfT0nTNqh67wyJe3wMjvDL1gBkBvLZpviZp1rtpApqe
VLQSZ420yEqxSY7QrotQxtj186sw5vLDDwQZHPiyho4hgzOcjtdmwtGpdU3bpKTY
PxFND9wJLINqPyBVkiM5/5gVjs14Hj4DB6ySfhDm530E6WwcKkhPjZlsqSsXRFNg
aDcBgygCAlIfNYok4lwe45ZYjh+s6aGSGEEQBAhvh9NyUA6wCCEbQbwepCW20cYC
4VmExjEOXz+VNueni76L8jGmaBe46IyheExuDHTkoXECwBYv4+cNswy0wGoSi05L
7hQlJJYIgcMdpkAPyWk2XGp3mQj6UT22aJG3eHJbHFBvHOpsWrZRgpGqSZMRzj8K
mwESQfXR7iwvG3MlOVyqxIYNOg3IbXCtXK/zjCEItXJCkIVgZi2qJtd32V7NY2qd
ftZ5sHqgSoqj3BIyu6YowRO7wuNf77hjKbeGkQP/GOT/tM+reC3jjeEs7hupFxnE
JhLBaWxWnAfpgC0R5HinfyEtls0lzbzB9reONNR6FlSZI9imbd6qO3qS2q9NB6/Y
TX/pnGjH7nyvQ4zIQ5tMfIL0Wj14MoXptF1zLpNnIJQxy2btpt7qlknz0FNycdTy
omo//RzouKjyh33vO59+fEiWdwVG3Y2J19ET84MZkndP+FGRBmkBphdVw14vU2rR
4csbe0jYL5SQnQuQrEU6aH3UKLd+8h8e1m9sDjl08Wk3IqkC7Ni/Xniy08cjmeFJ
vPraYA70LBh7fndrDRF/BbgE6kpt59OlcO6M9ecgyLIKuL2Ef8Yv+V8dVLCm/yIG
GDQ5TObEh/Vryi67dQ/613nY6PHyQOSYCaQaVbRST0Q8unbOlii9skxpM2qGb95C
yLyEb2venly+kXizb/plLfQCnuRCqltpeszluj3bQ/Y//i8UfXfU5azp1hkX8dWJ
FflBxGp7Mpcl3btFcM7hMesdUl5/yaTOCm0HAFqcE5SMh680A6deC138rHoB/p3g
+z8Bsct6sVdqkTKNE3R0Xw8TjT8E76DWxrspjgssAc2oGipdiaFKlFflRBfgTee1
htvE0RAmEGq2KRpdY4VwxxzM65ve295LPn2CoEXklcZbM8y+qgfakU9qQUoXgPNs
hdVwRJk8cOSkrrFcG6RwMAnfyhA/Oq3F/J+IhUjmAaFCvPr/loj110L+aFLDmSmv
awVm8+h8GWpoeTy5AgjoRyaU9OIyjw+OSFl6ZIfkFPEXWKtm9Pmo8Fkq0lx0bD0f
VQl9KyhOWlfzT18efIVQvqon4wH1ZAQv/r2OjH51HP032OWxO4nncq5w7Z8xJwAS
tafyG3IOwUu85PzJhecuTFQTYrzbdsiN3gPBzA1Lo0mN6quMVf1QjGSncBRjwrKt
mariW/ulMx209AAYWCXMoIiL6wH83DC2RhpohUtA/7K/XpRW4xgcZdiALry1lQpU
qaN9qIGSU9BMAcE83vKeVdFiZ/yeS+QSlwxLk050zs8hjWYrXRZB+Ls3g2Kdweva
tcOrNcEsk4gMyu4lyv4RtsKDvONUfcMRz9zQ4jIsZwW9cRUeJr3/K2it53v+ensk
+xkJOMPx22C2D8D0wEn4h5xhGhvhNa5cY2f6yF8tat81oyQiGMMZNl1j3c1mX9sV
BOyJJtCAui7U3kHtX7GPm1/KjfP6Ql4AtK4esTczWmVIMLPj2qnFiXk7fPujia1z
WJu5UsUqprsWZ0/UqnSO83/5o7V+uBox0nexEt65FgEmIqyZJXZZH3XIVGwTC89y
U8AFpI0JTlUA5sSjiDr/fo1q/tNT287PxR+ZlSFWUwa0WKaSqJWVUBICOsDAi+MB
FzQUFl28F9AMcWiTai87jtGbcUu3hCqlWEgGCW2atOG2f+G2iPIPdz2t0BCm4wWv
OVyeFF5uvQ2Wir0ekg2BV2yDXImiLUx5YhchdiOfJ+lWzbM5j1lNhW9Wpw+B9JHz
yNZNy6/aAvFNLHMU/78Go8vGzGsF9jCyczdGAezt8Sr9S8vPZUjTbxqdd0sGB+jg
8xZCclk8ieYdkBDOARvLOnACljLzMGEdeR7/eBtY1dD/2VOFmDHXriNN3NI+sgDp
h8THOtCrUQ0+qDUYmjpOZRs5HBK4/I8YKVaiLYM/Q+KpxHca3DjMbkJl5YKdYsEw
aElJlaPn3ouXEiHtZnBskpMXQM4vmPEUY9Tx8mFqk5AhRZqOSFnrr/rvJ9TdkrIT
FmasxLDwUJeZq0VzVgLF4+ml8DutMrNGq79myP/wpZusINTrrM/z0mYj49uMfV2E
EKn14/sI8MRZMoydz/Gr/vc51zljbIZlQBESZISdsKDdSRyWXcQlz2aEQvWz+wAp
IZuDQE2uiR3L00xWzyxOHcRDUfij51p+tBtvrxfV52XwZEvTLrtlYCykHzVnoDYu
KDKayA49H6K3H8WZjfiHfB7zBF9/2QP2Tsanv8B57o/jNV4A1357pM0NI0uY91MU
Aa0PPEPuIgnMYrQZ3R+mjAZrCJKTVXplzrMRkwZlf+geSAmAgB15497rQbGLr+jS
jiVJbXuLgHkKnOnfxbOrvGDpxm/4KEaQkeUyZ3hrVHwYBKZoDShDZXGvPSGCy4Wb
NqW+eNTJ6EoTIN6LDWHaOzhapqVDuIbx7c6iuOI7AIKjeq7fZTP9o48okzdtaRkD
2EzDWK/37XOmAEdYt096nlBBJeyQNZvFzRvnPd6MCwUXmU+8fSqInQ3OieDqvfr2
8EdMGALv6nTBGA+U/OpngWbXuA5Cl/Vgdj7ieGQ0QNvZ6Dtrsa0cCJ5W7y4wWUSi
/2tN2i21tna8eyg5YxSpcP+5xiq4Ldqsf6p1wASa59RWiV6oRwPh7qoVMHu2mhLe
BFCp+Oea/AHY0LKoMj5ugE2B3vJIAc3HIQaBDde60CR2VM8iTecmGFGdCUSghpTM
rtaUcLHVtcvtL/tvJ39f05LR0ao43SNxkMekOfDD6i9wgFsQ6YANB0FjZRgDw35U
wBVnF8YcnI+1q47COYxaWreRJYOP4s6NYbKI8awthj0VxKYa59ngXCsxm3xAqH9E
YGB0oq5moB963t45DErfd2HCA9ui9FUrcpjZly7UbdFJ91xSlYTrxOEB4CxSdvTv
YenQIxVDkxMfr7hA1PmBfoMba/Hj1cDPl5hm6WU7iJxSUuF4khpg0dDwJCXHV0NT
60FHopV4Uz15h/vbzj/iDJUDE2iIEiaZjkWdtrrjq9FlhRSqgSj/32hVFTj+9Xab
Um9FOR5eoDDIoEyfrmL4I5DTwCvCADOtW4dMV2zl/l5/grZ6zWm9S3iRNvE/BRfG
XARUJvRpV+Ore50dkxg7Gu8JMeJlPhc1xJhLsx3rf18uTBn6U8IpzogBkbF5oqZ1
SagbNyDzilZgrctJqaYlfSVQEX/Z0UX5nxrJ0ODJ31fT7N7sWpyKXhC5xqphKgZZ
uOTplo9mrZb3C0lG3m//hDQP338PNHptBESbLCLj1lF2J4i35tk2Lr1hb4HECQlF
rebJVaDgea0PxY2zqqPdeEnnH+FLHYI4FvEMqLMHW/e8Yv2lB2t4AfA4zpRYYjv8
TX4trdpx+JYgtUoOv1qS1vMIdhtIFu2741tUHHduUTYZfOhedxpbOTW5MO/EXmZy
48a920iPoGfUOBSqejEl6861A3S7YrhyhcBqHcg6xtJydi1p+U9cqzR7UHnoCHiC
K6iS1xBIJKyrJO06pBEy6H9ENkmAB7SfUoz9JOyhanalpLVW8VPW+D57SgNQrJlf
vmdW5BgAwgqaF/Q2MLYcJbX8t63hHQ47vA1261IuvySnOSTkZGJ7BRBjEtjLiq5D
vDdi9HnN/cXBu4V6RD0eiT3pIiX4sPt4HB62gXjPu0Ejkm6h9V1kfbzM16gOq5Uy
YDb/FJDmCj78MumRnmk0Q7/5kUWx3u7Twv7EiCAkcJgyveqA3RnmbjgVZZzGC0/g
DEtXw8ZKME8zAycup92AOqyCs7j6oqSpLmZ/L3V16C4zRjYSQRdotPlOTxl+qBsN
M2Lo3BdndiUsUM58miJyiy7bKspBtaRu6pScOsGaWx5v+VWRgKTfLJOSqsLVErPN
5oWN3PTAqbTKh2/Cah4CygdsB7C3vHRYQHIWjHBrTDz+MGSHvmqYU3biGlKfD8x+
X6HfkLoRFKZ//fY8o6s4eZvCo/0LnzoQimygmq0sMlR/5Y7nFSi3HPG1tpXTr0ou
1WzcRZm4nOHAyW581DRsxm7zuVhHRMHDuB4O62EndCisyUc3J/VmJbHlKe6QxzWi
fJj1SrgPTd2Ar7XfoZiCHFpfmVbuHNnknE8A7g/+HCLSjds/DMY5mLUiY2pVm5oK
vaEDuppg6R9cBTJA1LcgQubLlMI3AZitbFglEnCkUTu35x1RI3Ap84LfEGf+ipgx
+GUy9URa1YSeH5MGdgNVL+QRO0bylCyDD1RuPDrSuSl4igbkJZMCS+TF4EyBUzX/
HPmjZRfmDiyAMLADybknuFKFAxvs63iXDDodscLulRilKd10ofvIvmu0d1dT8f26
osTNrE4MvsTUNeI0UHZK+u3pZBx9jaku35jUdek8aaka+GHG6exd9udUgwsicA2O
csCshte9M7O9MTKicDUGMEyeWgII6R8Slt7ah6WaHzlN1o2voEHzykYzq9jHpB0D
Vcu3gzEnHLv/oSqcmY2VW1ovMlXUuzi9dDqpg1BNGtFHpCIuqfXhO4tlZKcJjF+q
3WvbdzU856dKIpF1QVAtPJ5P1B7OPyKgjJvbjnOk3bvpjho07ffB2yGAYSzJdIUG
vjBMLcQKIhhVgbDeocBzM8fySI+n2Mm9l3nJwQHYlNls0r4pEXL3x1rpkW7p8dTA
GWgsWXraQQ2xI/OsYhAnARhQhOGWvZ64yjUuJvRD03VB8aqq3eyNJmwWHnNwRWIt
VNhyhidby5U900bY6AzN4q+bgDt5SlOjzgYw2KyZsCY45ssYt3/9UJVsOlq1y31O
kR615ISf5EsRNQMqkK2N0PIYKcFtU02KuK2mmDx5w42BvkRrypHB9fsB2swjcqZs
1KIsggROdKz0DpB3SDMib8KY3RBDJ8G8zCIvqUqTMV5g5hTX+i6sMdaz3VxNjcMd
Uy+UuvtJCMAhbUv8yKgPka+R6TMAHLJwHyaE51EpLUXtOtxxzZEtxHD9XIt0vgTq
AQTO1X9SorHhy/9xPk27SKe9EJIiB/3jNrY56JI15TKJ8WX2lQRGt24MIgRSngpq
PXJHfT2/eWHNU7aROjVJ8OBeZ1asaAutiGvMftL5xRvir2hXT+UEI5uscxt1jY6i
S0CGSVxVGAJtRHGQAuf+KcpAW8mH4kKuWiqCxsQyFXaW8ywITP7j2pjAs9RE8+Yk
O0n1OJ0h4OZ/wbn5a7cBVBGnt34g2Gkakpu7aOEzpNYyo9l5Utt3+kihZux8wE/X
DEHdHiUBv/Losbt1K7PQcc+vhAOkJENywoSIPfR4TuFZUVKACkbhuoB3hiDOkiyX
yUs7KCgfw8ITk4znStQhs9ipCTOZGYWIg896G4NQa237O3qlzSDSTrD+e3ABGR2C
LCh5piFnjWuiHXRRtx8DNQZeqA7lNoqGrr+lbhfgUjxGF985M0V7C1rB/IGI/8OQ
4rGdtvnxf9wcaw2NqBO95NrGZZHTFCDfdjijGl0ajwcwSoZo+HoCZJMI+M66pf1i
h1oYCviTnMG/uLp/kJDRHwIS8p9q5IlL3Tpw9LdoNNZWGbhfEC6pZnPjr+Jkdm0j
++uWCwkJDr9wcjITgpUjmneqxDJVpKasABncecJ85IYt/IVKvmdT2wkYwg9COYaK
7TADUyv+QnV55foq55V7BFlv8y7grGwPxX6kLjNEm7k/6OPj9C6qhS0qQj+FJIgj
p1Ku3ny3UyO+JgjQLpIPbbeyaR0wO9GEfeBAONELyK/ucYyXgRXC1/GlWoskgMYA
/iNtAB+kCxgb5Qp4jtHtit6XmcXoy20i2O5DnFhy+oTs/ZdIYQjOujkkVQLUhuRh
FBsoWKGCNLCDzFoYclKn3Jh5+26ToEHuwnr7YJgiejBQUDxxl0lPUd95yKTXrm6P
4Y+3GBtZwlQABHx9emtlTLI9xKdap1XhDZbQB+nHGvt+VrO/GWM3pCfE0ksKp21F
jHyvMcPH1IDRY6D6adQQle3o5I7NVUYYg16yULRgbmjF31vvJsgvNZthJI8f0HXH
sOR9VK6ghC2de4LG+v/DhsbkOIx4wIJc75FlCjChaUZXtSx3cG63KQzBqZ4TWDLj
Q9GROHgVN1SxAEnZ9nZLfX1Jw4k7Okmayb7U0YRmrsrhFDK/CARlJZ/PUEC6SFUF
01dkPfU4RuGI2USuuvficvmAXvWg4p6ZyJ6zfKARYAXivShifCGQxLz3oNIHajkU
c8dtyp2rdWoA6x0P1rGNDUSuJtrPmEo0G/peiJZefo8aaSz22xgamhz/f5rLtxkQ
a+C7ril3azjm8yrX4moBHZ0fueJSyS5F/v+MBc1tccHc0uzj664ntyI+qVfeViCP
7cWtd1Paf3F6sbhX+ZFt1oyZe6L91dYsdVi9MfZK3CbhwVOGQUtC1x1SluUmLSBH
aVjMs68Xmk+9R4TyZNo4L89lla9ecLukmP944evZPpfnmJcNHPnL7agkDBVxdiA0
5wi+2zxCyZfiNm9xGyVjn7TdTWBoCa1SIajQqpk/91la5l2ATx2Vlr346PjjGEP9
8Pl4/ls7toUt/HqWhPdIYZJWLYIJge2nhQAomGNNNRQz6JnAx8kk8xz7Ct7F5F9R
J/AmzHB4Z+GgGT3eWk3jJaoWWE+WNjDBu0QBn9Q3lfanmW7g2RJpedt9Agka3du4
3q3MQCxa+CslbH+MTO8kwD/nNBt6ZYTtgsOlnL6UMmTIGlXEhvWHUxoHSb+Y6DA6
ikJUj5h5ArZIk1WVDroEYCp3fQhq4/3SR4OV+BHapeb0MQp9Jw0If4ZZhZR/JNXC
Tw3hyMlEL7btaU8uh5rXIINZ7/MAmaLFuqdHPqinMgQhkj1g4U5l2+CuMIcVJRVC
6ua5hHShqmQjnij6f6WknZxsiRAl/m8MvsrzdZD4zg8fyRuKww6TPAM/hEjXL2L3
I7PHxX2Ap3uwSHeEN+VELHIrZLaxseBNSgPJM8iicLIPaxWU70OAxJakc47UkfsL
Md/YQQkQ0KO30TNmI6035VsdfSqhMQ+HSkCVd81AleMgV0qiSHslyLOhYgiyqUsY
gL9+8DPeFRa6hXgdUIAxYYjzKxpVzlEdZFjAjXpjRxIRq75sRbpepoZVena+Fp0k
p2tpskjFkFNKi+8LuYdGKapsTZ/2XAJkYzHr7n06eL4deUcVu84p5Q/z/W9Ya9fo
K3D5PKt8drHfTvuEmKrG4hcIBEcRdDiWMWlFI9ruzqsaTM4cjg/cvqXOPKzu6ndn
0phgazApmu5rtI5wgv6R9kIUnBsYQnwffutCAuinK6WmDRT275SQRg0EECpXQnJ5
PTLk3pPhiTJCbRGUJNOAbbsg3oDzsUn7c1aHsEVs9MDrNPF3aMaZ9aq2rbjctuj6
e/D59MDKFg/yb9GUq9FL4+Oih6S0gm+8ltHvJO2TrT3W1wZ/WvKiiICPOFwk0NwM
ZiEFgGxksdk1MEbuEYVzAcKvdgACDUNMPY3NH5nC+xlR6PSp+S1Cx9PvDPsXBa5p
q3VcDoFUHP0XP5PtiE+wm7OlucUJYOcANArtPk0uaiD7zvTgbKg9yrQbonxNffUb
lc1G0Cu4PabpwKLzDlOIAqunEA8X1VFBWT8yB2GK/NnZaj8KSBsNSG+o1dUbiubr
DqwDDva9cjkOOtgunD4mAz6tClgpJTzhui5UN5qg8Y1q9JwstaGaeVMyUVvR0yT/
m2fyzyteLcyBj+vfhDOw2iqIoEjyHb/O4pqQdw5ohHE9KxNMP6tuGQK8moKDezST
+ZNw0cVaDKheaswqqhNF9vclRYtji2aKz4+msKL3n9yiIFZUC8vBMpUs8aj1k28h
tFQ2nWQooAkjLEchEcIL+MNN8oHkV8AOAefT7z6XiwEJ11m7BGbpw1x4v5wsIqPt
pruPJJCPu8Sl0K/zBEp50fVAN6uQLCN3gc1juDsvboMDnWNzpP21VIxw56xyIKsP
LiEK0YX18vo1i3N4NuFaw3kWZlbf6De4YMFKpcy5YZJ1XyxDkB2dklx79yVfyfLJ
CYFAZok7j2GIEiK3T7Sw3G1doJqLr7DSB2o1SlScRZx90cBcNujjm50dA09DWLG8
ZHwPyk+e2qnnTqn+mMt81rjHASD9mKV0JBFJmuo1FdxDvKW6i9mtoyex3Srzl0gq
8fmOArjoMyiaRhcdUXxrJxahsgEp+xZVmt0flRg3boKPa6fPd4uq/iO2GfpaFfkl
/B22oQv861GSYzNBa9Zpvzt8zsbOHhls/rzUjuB/yPwoNAMRUQqPZLfb+r6lGV6F
Pji92466DBWV4FlIAj6MkArN+VntxPblEjJy3CIYWo6kc6tqY0GPunH2tzqi/PwX
QqJ9hK/R+ubwQoqhMtAqhG/Xgu02bd6JEVwhzhOSDN7CANOpW+4f6m3pcOwRQ7ux
A8f3xhyHzoW3TEAXjQTjxPxozH7Tk+ytv3yMbACAuTq93VKzxrNyfTmuQKngrkNS
LpNCB3NkEoPyWHqkA4RRXY+U9hcdh0SD6SIICrSmyyarC/lkUZMQGRTWDV3pOEX8
sJ47zOkKdrCslkPH+0mvq6QTfCVzcDFS3QBhsbuUue7yGIjDqkPiXMKrZX+rAgZ3
ERVdsGQol4vKtkj+CaEtWS/8b6TfelQSa5/oPw6ECrV+p0pVlJBB43eLcrSemnwb
c+zKhPphkbLaS/y1ETdA9q1zELR330z1oXAK7/a+iD7d2Ztw3xta0PRkIG6eawTr
mnC/pwFPp942GWpICRSaMWNsFvHJPP9jiJI/K4pFsa7IwsxIYlrFDxmzpdfGIgat
S/54yfTXkshYxMoxEfTMQYNkJ9gxE4QvvHXZZ8hUzckBk2h3ZWH0GkalnqIJ6DIL
2QkumebNCJTF+VEgYKGfBUDJEoL6KYiyeetKRFje2vwpX7qujnAEjSvodzlK8MjT
xPPthJuZpzDHAQKGxyZJJsCwGbLtK6MUpFqvCwZ2Nxmy78yMhzGy2BKYyetWBrac
iyzq3HUG/RO2aP3TtV9O3IaFecd6dAOBbBueh9x5RdifXbcOEUT8ESQvGhbU/N5z
9whiC4me4/8mXuOOJ+rDGOwbMNJAGQtj+szjYj8WqSbN/GCDs3i8VMJknNLHRlfE
5tD+WtlAWOWi7UNjyGUPOHsnzxYiiDu3XXodsGASZUmjXyinuCRGk1U8WoYyVphU
Jyu7qh+se2izxqJ/OcfJMe1jQje2+AEuP9UZEQa7pm1FdqIaiiqB0RrhuH0s2wXw
ggvBFiml8FUkj7ekuG7yySeLBS3ZHMPmtitzciewgq3Zr3Xc9uVkqZjwLXaAgYzw
uWRg2H24ytNOB0s3vMnvjQFg8JlMcif8YH73jyvIR6RvEBMAIAc83MGWiayoDpXC
BzUFNDGMF7BTlf81wxmM3Z9RPyruSbD4sewqpa1K4JJ5kIzz40jxKax6tfyLUK40
M7AFA2WWpJAQW5hgjZxrOJBmAIFAif+UAfqNLhqNNh2pK/4CfKMuQNED1KVWA0LZ
LSyFtZYiT7VwyenxhibJgKZJM7DvYroxGnFROv7xykA6qVBkGKGGz4ZCisNmOu9X
Wo7vbVVNokdELQl7toHL6ryxrdrcd32/aX1i58S28vJD5Ap2FUzTZza6T1FZLien
nnkahg+sxua41zkYLTnNKOSbxrNfLh9encKFOsRH1YyxipTLx5OOirQPbzN3qegf
66NLfaFqQ47CnsH/80oCr3zuoXWVXVq3Atf2bOrl+GjnjlOhYmB5TTbPqlX2ddCH
NOCk4+b6DS/B/66RoB8qVZdeBf9ATUKPcmd6ASThcjf0ORewNFpwr+N0dpRM4u4Y
JO6+lqp5QB4USTpoQFMU0Jp4J//3ebpqI541/fLU8ob32un054DoPpi+Af74gkCo
V/f5isIfnhJf+lEWWLVcr+7+1sQlSqKhIj2vv4/lHbCe3fhl2vevPdja4a8dvlmV
6PuBIJbTktfzrJCbh78/hZ0liddMsEb1/Pbe86LiPUXFEimYnBdlB/Cg3g3M5BiL
YY4e9DftC2EsUevbNpj2hQt++4nUoyCaJp7902dk2nabCPAfvfd9XdPVIDZPtnzA
MWkIjrTZ16eLDi1yax6FZ+oT7eebct3EwJuJHhxhRsk6G2Tgh0uNGxWD22DY9GtG
+MC5+Xif6hiriHQ5rK3vnmiRIBKYsZH+RC5YQE85RD8S/BOCCeSfIymPZGJmL8Fh
K4A+mhC6lOeCtGjKYvODfM6DqwP2Lg88vOk0mGn95m59LEkfCFrYvH0Yz6z620lV
HMU7L3vEAJ4jRlmimLJmrDcxH5/y8P27cN1EQyjUBuUmurtlzTJMOU/NqS0TBv4k
a5BKxiQQuDZwd8vBOAA/ayrF2IQO8rk1oF0A9Fu10nYOQEUT+ucEyio//HCXDWQo
mcj55jHK2e6FChsfyC2C2qLkJo2x1F22kUyPnVJIFCt0IAFTRXT/J9M3HJJeAh9a
ZbCIAfEke1ebDRWmbBpRj7MjzGX2/kBrauno2WWZ7Lu5WgVVpCuboyfLQsWoaGuL
+YmnjYO635R+IrCEXAO0S9MyyybLvTVgGv5yiEI+WGwsFJNIuz2LKA8oZAxZZuk2
HvbyBDGYLHeXPlQ1XBOrdjPbDCMayTW7sQJZ4JsAiYalALZnnkVL1Ot2khsSOFEp
FGneXJR46r5QM0RXIBuLrnwjRAdIynT9ZJ7EN/4M7067qYTtVuEt8ESTC6A1Zxqh
us+0p9eLDKW0bU8+uzSl8L2VE/HB9mlKPPIqMLmJUh+97KPUZ9MEMv5ZlrbqgyW2
zpv9h53gCeeu/nasIUgxkOh3TEJTT228y5rYiS9LUIsXrDVZWqQ9KrYJm/ppclgn
ZU6Jja86I2HTbaleGgzH/FVSpPIMqZIAZFsDFjVmz/nJ+dypRH29fpsGrPHi27dH
bpqunnMgSIyW++sG9SxG5yas/MIetIWrGrtd+6ksA94VDc01EFIst2RbRNdoeDla
SmIqhTpH7ClYiVuG/FZGsiB4vjqVrHnzeZeR01c1nOBSPE3zcgfv4tr2GFPyxbvu
DdwHTfKyvU5FbcCX8hawpTa5BcCViOcLvi1HBWoQmaevF+9nacNUZ+cimPBHwipM
OrGvBdrIKPJbnSk1lFpn6kjx1RrRaukfhb67KW+GWtQhJOASGWCHrNX15L2iTict
soxxkEJ45hAWhRL1dltJE5ex5eCl7rwfEuu69u6mA4dhbyn+7dKdfdA7UTJoS9Sy
3HF2Jor4Y6O4195b4N2C1m2VojBGL17isbfAek8Cp6Kuh39pgt5gbHsJ8nFs1OGz
p2guOIPn8zmfVioudg/LdJ1ag+sRwaLdpdVuN3MZtD55aiY9N5DyXv7CBr4eTne1
FSkLQxE8qXzOhHqSNvgHg5+C38lFXZc26CE3M0R7m/TSxqFSHHVsBZ1TfNHl1lWj
sVC85jA/kR0nQ1MQf4Xj5G4AdKv1XHLVM4TVpR+42gZLFtb2gO6UxFEVScUnj00l
wHrntj4NZFObka5bcInlfb18bpZAMIIMs5HJAbWTFQvHxTPkam8SSWTOPdgTmSwo
8n3dqmjVn05sf6Rki3h4NbpybCDN9SYq51kP25Qiqcz1k+h2sRtNOszFpEmgGxXX
vPVt0UOtEpKPbVGwsk06t92tf4i4Yl19GYEYl0/nPsPQxIABNAWVLB+FhTGtO+QK
IUoW/3Fedt/kD82GEPdtE4C6Q2FRpR7yK5PgUz6YzEcLRR9XsUDc2k/BRgkLU2Kc
A5eUw4vHCuLCgfBPIfgObc1rDKfCBmv3vWbItx4OaJLgbqe6xgnRHPF4EauPsAfk
+/uNvrP60RGw6pyqu7nPiGjHFMgL3hWJY/RpDmUJxvRBfLCgE9/BFlwolpVnGFcV
v9hYOGCN/9RJ9sCZPOfvLftOOuSygrqYnZOHK4wHHtAmYCy1cZLAzmNTqOtn4Kw4
9+QiLT9IXJo+Sp6NNAJYKuLXQGhZ77LCLOLGoEKK57dZBS25b6DcEFq+4177Wf2r
2Xu0pNfVAq4Dobc3Pc24KU8JZURXgzR3yEsv4N7MargsvoZxLLooHrd6CndYaDd2
8K8t9tRItXAlj2yiD2c53L2bGIffgNlgWnbUEKrCBabwl6ZBssS/8KYmCiGGpWXJ
1ITro0sv9sH75JEMmtFKVxnBIN0q1nqLmz3T/J7KImK+6R1pN/gcCH2eiR9aVf2X
uI39XcXqEI4i6kD0uduhpt4k18vGlt2Sr7mNDZeBtKLKXdQldvtg8S2AHQYDgHS0
xcifWCQF3RROid9tFjN742lxVWsvNuGVkkp12qF2slVFNEU+kQOmSfwgBMm3k4XO
2fECDrnNQveulJYxJAqVZARidIGINL3nxcIQihnm0OfonJFJGMNoPy5fRdueaIv/
+/NsA0HPuIebcNLJ1sNuAP8Q5mr3QIx9Z+v5CYpxNsyD2Jfu87/+75AablXSe+HE
8+PeOYiypgOyKEQBt5X5vZasiALxM8nhRGSvZgBB6px6o86HAIwaWveV7aAzZ5jp
HWXJayAB0piaqyIDNzb63+PVwwVdNHInO5WR2BHBSbWvpnW6SCvC4Im5DH0NRIWE
AEWKTRqxfeoXr4Pfubr4JFon8ALj2TrPFcb3s/NmUk3xgkp2LhGTcc6M3tJxsNqV
tN2e1NqTGbasUPYCsmB0MQJCyem9IOv8fk0gCWcHZJ2JA/xkzXvFWcyWR1dX1/v1
okWngCfW0oFtGhQNALJT7olt2Y4qylz3lFrrJfZBIlb5HYF90QQwsj/5bzWbGKfE
t2FjDXk6UakyS2Dcux4e2GQNfNsoa9XOMH2BAJQk8iO7iwqx8sJiT5DVfaytnJbb
YH5B6LZrC+uFVXCCIaUiQfZXVcXxImd6zZ9sA4l0/X5eBoNifR+rWwzxHSEJ9vi5
8FJN8PFfFbCuWf3vRlFa8RJb0OWJOCT/cj3nhILtn96J/Vk7YfDbIYMMjrMVGVSC
os0H4zNMQIlnDKRGOXh+aWF+JNYTUKI9Ygc23s76WQlzNW+uWYuXsxQAx0+OCIrb
UtEfQpEAqn3vqYWf8S8r8jGsag+5gIdB+ND1Ss6MbG8egpTbXfID5V36T8y4IBb7
WmHWTE0vtT261foXSYmHAlxHY4uv+4xamq0swjiZvCcB0adBxALPHMk38Im7NFHW
adGhhEhCJb69u7lpItpFs0jQp4Y9Wu5RPkMLmxFgzNa9XDWWs6AkYYl36RevZWAo
L0D475WKe61/3czJEexmvtgJcrh/J/HFekx0H5gc0MVOg5p9vhNVzw/GdBBnBs0Q
rw/nLw4N1afqjvOBy9NKmBCCDbsGO2/1W+MGIIcB7YqJP/SGNcx0UmnIRffgsVZ1
/bZsJLYa6p7eQpQzeLBsXi46yTG2o1/Zj5zDRLN+P6kAZnakxrq6DKneVwgGwzdZ
n0Ly/ZAUzUbRPXacJpIguTaZMUkD8Xq11jVE7MBzKsZ+pWDFHc9GbyKzpymPISbQ
f4McVsTeFninedW7lk8kU10qQb/v/pkF3ym9JWJldjH5oVbSuI1wI+sM2YrgaLU2
ti9BMV2EYkgdRlRO6lUeRWeBr8SJvp7QENzFUW8utQgO1FANFNaNj1gzKnu/MMlB
OC/PGmWzXbGKki9dkaNy1zipEgGzIaX5pHudEeF8SRuR1Sx26cl9erQluCnLPUdC
8SmZgZMzuAfW/y+Vb+uoJjXNHCtafmpNutx01ZG75SmjvEMP8+80AVQEX885SOB8
6EkBtXu9VN/hd7315V8bXkAC/Pt4E0ceOP9K2QAzH6cRXnfakH4mgeakc4ARHLaD
aMTIQKV+uGemauaxQrSjS4X3W8DXVU4h3sP9j+eq1BK7/UNLZkpbNZyp3WvNNZ6J
zxl4kBJeGMW1+42JJqmWO7mppwqbxbpaQTCEuYpsailuTnanCZ4JaDWwjJKeoxhA
5jQsCnOW2OUJ2ZMnTFkDaJspYZXbJ2gDtdUheMOkk/+igE0ojRfg6cglZs763b4a
32a7Kr3S/J+ODnmrZr5t7mg6fxPzh5fkSxGBQQHm7iKfK51tFk37QZV4ZV70uGED
mb4FPfYfhkEtCsS0p2U8v7WHLCjJ8Xxfr91FE7axwn1HcBqzswLwq+vvxFK+cE1R
8rpntq5LyRghEuucDONA7xdiSaS9mX9W7mrD6JriO099VfiiHaYVdFSaznhtOdSz
1S1u8/16axIh1SGNyaTkFHN58GLdYaO8+9YZo12Ap8WWz2zFxXNq8vQe2o0o+32m
wrr+iCue1TgULqndgazjGBf59EfzsZzp9Iol9irFPt96Qu2KBn2eSOYRlxMPZnz6
0tZf0masaAjpKYKsov19e2YfaVPzZnEAtayNhs2tgjPPoODIb852qGIWeyqZu0LL
zEuk4afhJ4EiDcZsVActh2MUJeNPDNCw4pgV/9AkHa4M8EBuQM+WPn1J6qPY6yIX
awHeZneQ8RF8+wB3KPx5bFv3vl8uSZ31N80Gv4cA4kIqb/990UKWCfXagq8JYhfL
qNGNWF5fqKXLya0U1nrDMpYS5ZKtJfNoi3QRkfZgLtynYCaPDUbeYiPSBL5Q+6qQ
EZUJ6yzCGe8RvbBKAJX+1EhdrHenYnGkwtgtkwBSh2kMYZpTqLP0SQ0tGY7v7tJl
rzJX4NEuz0+XL2zlDOlzfiBTZrsG1GTKjlM+yi6SHguEZ3G/w6X4it2P4n9hbE1U
yV9zNKOFxjTwICOn7UZliy7qoVd5n7N7V9620xZYZX0zYMcuwyA6+CBcXyh9CqeK
6ACpdlWQVvX89hJu7fz6f7zoS13CTXC22SkbLKJCEFY6pCs2tyby9sIwJ49xBd+n
rV1+boQP/ErKW3GiXMlufN9FGqBgPJP6469jJI/7TUynYwahCi4hCJxoJk0jNuQr
96MhfjSS9258ooJu7VGgahUWGMBDUp+SFhsNHnoob7EPjwMaF06JAgQdY3vjrPGV
D3u/k87t06hLZ17LTI7Y7c4j9g05eO9Yl+ODUG54L6qC9vFE1+E0t0UWPsCBCojN
79VXAen4ZPgzOPSiYQhpVGQKAei46AA40mYhYevBUMSknFaaA5H69cTypGCjfkN6
YoAy6RXDmvXmt8Kn3VGl0MIlD95WxB0khhi6R0QX8DUs5ktT/QRx935TCuE10xYv
BnOTVDNsU4nPDAkkaMTsozk9ggUJIu6mp2ERbCir8bSmtQw7Dn0uyT4KasKHjRSt
Rd+KAVTxmpjL3Mtg3/5BOJnqtLkD0UiASGgfGLSSrkKZLXeY2X27LH4i8FA7MfNj
yXdIlobwFjF5jaKnoiDVtCdPL6L+oh3grWjH3PHP/Vw/Zs1Ypi+kf9tupNi4gQYX
Sef4+iRcfIVGZB4S9Y/YY5S+aDFJDBfTSEghVbpuTVnzEQAWV1iEHnyuvEOpgphV
5A6mYe4mTYtjCeAr+TlLzkxzl96+dcdazPH0VQMs4QqqZfQXs79Rcmj/kDSmUIyu
FMy3V6vwqegxDWS23HohcW5rxDz01BCNy37agBRmLn0zW/YRkuQqokx1X/cvoI7r
Do+Vw9RwNbcVV+jwhAaLDy/pbeCqv7BiHhrnFPwuFz/RAqIw5kg9cm33KNSuL/W/
YgE9vZR1/8f00x2+HRr7Ze+0dC9TUQBH9oqx7Of3NOYvfmMcXz7GAca8286z1rTA
Z6wqMnMwfrM1D4LAa7vPZa4d96rlOvQDSdNAPYoB7OrcOItQS3ePeHwDxB0EVAp7
29KvywXoEW5anBol/lIbO9FN0QAZ7sxuTdjjSf639zmNEb6rz8zIwMxKC13rOE5z
m09XkAzawaT9qWHW205C7SGQhCn7igtSmTJJysXvVyykLsnkVUBEdBvCTr3zXGau
FGy8cCbi8A7uXb1JtgbUtcVSlUvMgrvcxS0AtrWa9UyIt/7Y9k9h3k3FpzC9+hh5
Do0sdGEfwNqnIFNY+L3V5cgeE6jLaKPdarAyQCuRSbhYsYuLbnBy23M7tAL/uAeg
5Fn/oxGP82tS7i0/b6StxXheyiMCO59SAVOwbOTEvxAqtbVk3OvOoImp0qbdSjcI
2k+gj+39aqBJ788Yojcn9RofM3EhS0Ycbd1qTM93n/aZiA7MQ0xoIb3o0+9kjgOw
gX78dskN8R6uYp9fbMU811/2ityxXBkoMfN4RgBWTx27lO5DjEYzUgmC+NIsMjYK
8wGUJhtK0HEGkl/0sUECSpq1RDmWv9NWBl5+hZdgmrwP1rsXwaBd5SJbC9u5rk1u
NmpOdi/TMlV6o18OqZ41Jp83u4XP0nngQIiHFq2Gu773c/uEaGIZvbuiRsUGR/UL
TQPu+r2gkQXB/YNDb9bUA4iZJbrVNh1WvGAD7cb+IQJOtSJA4VWmiRf38jOZGY3s
XdhD1XXbpkNj+I74KS3h4WfednY4PTXnqbtrKIDAdsUFNMifC37lKBTxMWrKtC7E
7zpn8eYPx8xSQeC1kzCl4IubWNug6QWfJaG9pws58gGQsWzY9+qA083lKcKl3YY+
FHK3OYwUI7gGFOWsjQQ7aq/7XDJlDfCV1KMdR+Lnyvy3x7zFA5En6nPqTAGg6QFK
TUt8hTAV60dh4FUnBq7O4ems9pDmhHqbsJiUNM4/RlXHlLxYvQ/6NHPH74euyt1Q
yUFWAveZcmNnPmlHtyYktc9ZzbJHkizhCfXiXScmu6uqkqscZpdnVnGJieVssFY4
O2f2vp8dWedYjJJinMBpYtUrhvqSrWUsvCh8cufja/mKQTXOCBobgzzvnfzb+ScF
EX++U2WPpvRpdO2SYSx9fRGG6JPqAxdbbKXBWMmbJdhI5l2H4iHdlRS0zsUDumAj
fZCdFyVEeN4f8IiSSf3648F0vqT12Hi4T31VtMvYFbGOxnzVkVchSQPi0GTcFUfL
vZ46sxON4uDlsKh1imp9RabM6dG4sfyHzEgFhj8NpagrCALKd0biv20bgmWj9fJt
YTPxcdUSXl+WuD0oUriyHWzGRCGQxvdtn/p9K1KFJAJcV2c4A6xNRQIpzUWgnFZP
I857TjScXOObjVlYlKWMwrwkXQqw4xSa+5JhTZ0y2ewXvZaQ/cMhz+6HUQgpfm92
5OsvOO6vBPj4ignHk7/oMhvsBXI35C6PlHY4e7VSmQ8oz7fP4KLPUMytPWuK6SSp
9xf5Vi85Hy21KZ0KER3bLUXyWdkUu46rI7TZmWk6COP2bpYOVDcRPjGmfDDpay0j
6ZqZVj7oObxhwqCy3sI2IIMhroBWMW4Qtzlg58u+HzVUEMbpCJLgyYMlpZi20vNe
ntnsrhERyE1zNz4ShNtO35ZVDh4msg4iYlesGzzg9322PH1dsUa2OqiW/Nmnkm+9
n2IuhwKIuQtYgcdQ06M4buwBi+vIsl++n+L2p621fo4uFkX4jnhMHtDUJ/T3uwLo
ugkxCAECO/Wjtqf6TAaBeXg+9JYU3L+31pCo+CHcgxBl9HzRCRRlLkN90+CUUK0O
b2oauBFQ2kCTNNlHoh3FyXYwBqsG3DhpB6zhjciIrnwcidLon4mC2FD5UKvukMhF
ShWt81pB19L7dgpIGcohl0eghsLq6EucsDIIvdPi1i1jx4YdrmFj9RXD1nmqSPGa
CuzFPihsS1TVZIfVv3blaJ54PJCbbbMdSlUyzHTC1NpRMLqpXl5+laQcuTUclnGM
6QXHW0Otxv+kU8YtEQDcEYnMB3Qq7stDRNhyC1hcO+KDLTaeaa9aHBQd3VkmEmt9
gTifJvohRvWXPB+sFBmomBxTbCd4CNTkF0xRIDtAK7c72KhgVM7g7JMF1VfHPBvI
FmmF5QkHqlAW65OzHMtUi2t9Qq27wqtiHYDdxV//+BRgbzouTpIeFfb6RKysoQmD
TZdoCEZUdxGCRMjGi3mPnyXIdSyb1b8QfAZnfqR9K194UhSXDvs/8iSr9TaN3SF7
vqZ1vCsYhpuEKaEKpJLnKLunFxyGFSSbz1niF+vY5aH1IOe6D6Xl4A+8oiwVlPVk
m4M/BtH5teMGFWqo3I2G9lyEWiO0TXHl/u48Hw7K7zaospUgety1G/jfbGLkXb+g
MctPaJJZBAIDnI/Kz4IWuoRvei1fUBomGsWkSl4bPegriWWfGO6F87F+zDs37Gdi
70XFmhgiL4+Umf1ERcHIkRSa7pFHU/lASV7EsFkz9M0+CqJxj7PmvXYcOhvPiZah
ZNsxIHF3wzJoaO0CJlMrRKNhnCw+vrhrjVVD7l+J01BhnlUIrru21Q3kC8BMG8bH
h53AjtT0O1AvrZ2TbFjPjdgBEDG3+QQZ/6AkzRhXONFGGaOvFmRDzoAR0mWrzjlW
JyrTTlFDWBT5Nfwes65Ht7ILHDP3ZE/m2W3TG+//AOFOZivr6ySoUTp3NfOJTPCN
tLz9pNYGEspbysgY0Qpd/WXuKPCMf6oWsTGYGiL0scxz3VYJHULgHb6m2rESRiwi
7rlacGH3QISI/4eDZ4V37CnMqvo1/LXm7CvOyrhyaWsBdGYc2DhWwkH+ywjpxJ1B
TGz9DzYyIeuFSFewU5Ysx4yagOonVOKP20ZxPW8v3hXd8CvIC7enWJzoug0A3S9y
Pnk1DvLFLshEoHIcz8Y58h8J781GoPEAGM+8d1oRF0EL85qK/7fsK4H0rBbJTHa7
9JniIwtl3cPw+y2OSzizFCRKEFqiQTOD9NO81xvnNSXbV5HAu5z6BYYEDdLzJk2U
7Q9K2YCMVMohOh6AZIE2tutK+zQKJYu7BcUOg9o5nUcJTkyIrHidhJ4blHmOkEdg
/wjXQbbMXpS+xGo9eFs1KpP/ANb3qEyDdorYjb3ZwiEFI1Br/TWWsLjDClJ++1+5
lU9ABvcUYVoP5vQftUZ8iub8SxWQ75LAS8HD0slyjls25kljqCZg77hKL6GVet4h
BZVtkpWZj7jlydNoVaUVB2GIDl4SzrRb2dGUcTO8Vu/lb1Z3OriUg+CKei3pX95F
ViMYS0BswnMpGPcFoWAGPVkhRN+p18q2FC4K4ZR/vhGfZFBuE84bu3tpr4EsWMJL
cgnZtDX4FYi5dUtnAlQr5Qynh5bQHkIJum7KZDZoZWYUQQfszV7eklDaYxZ9cZQR
D3UhXpZY+I0jNddn4Dcon6+QOrgnYXDSrT5hITtZY6rKNn7FMwQJftslog2lrbaB
n3WOnL6ahEXDwKA9ffqg5UcB6O7/gyv8JHN7LwECjqCIUFgT31rlRRiXnIfavxeF
idUy3GeUfhOI3weJTVr1i5Hs58mz2Ohc2io6JL9RDGENF3vajldKCBKDkIwy0ve5
9BCURfVPkQk4dfyQ17/W6sJHfG9XRlBvvrnXCoTMcLNYq2QslLS3GJT7aaOWGWnw
jqx2z2+hR0FUkOPsBGuS3rYBNj5VM3Fqn6Z2tvTh6YCF0A/wU0fGqnOtioXqx/Pv
IuBEC4VbCMYSjzxSgmFJKomRBR4/5D0eAITEax0VPXiu1gi0/Rzj/Lmc0IY078/n
XQG3RFClPg2b5Ly/SUrw3D8vtT7c4njzfewxzwuljv6sNSF5vPvcfxjcjS32mPkm
3XXRajQG6FYzWGXhMKYAE9rti+wCgSBHQhnTAEVDycGsi0mi9QsFXO67y1Id4RGg
hbAqsrT04rvU8umN3NOPE33Rw5MnuMQzjO0tTa0dpGKsky+qEwN/CCUk/necIR04
YIP8vktqLv6RBiZYA4zPjGxrv5rNR807uu9ys1aXZBAFG6Fd9AxsxumCxV26fHv2
9ccjO0cGWuTcanJ7J1M0IBnkQEPyU8ZqCiSahLbFlf9Nk3mWgEy7g8PVMP4gFRJA
ODx+3uZXxNzCukX85ASxDoWOaZSOM8sUozoTneNZbzn9XaMVwPYUQJVCBHuaDCf0
7/7HWdCaxbEdj6EEgJurITOmjDJr099vBIwoFBrxnpzQCFuZJVlbKYtJ234oYFaE
N2Qi4qXRTA9GuDemq3j9qvRm1an05RP+N641mzKDnHQfGqSIDPEDahx1d4U0ausy
MP36eKjT5IcCGekBgb6itwyPDDMQE90y/SIdmr/NiDE0PRRCH738KLTTLZqM46So
nihKi1aKwPFxx1eSvcL/Xl7KtgbrWBTbMhLIMwhXerYqWi8P1V3R9TSzGNd7VtQy
+xAMD5UW//TtrfQoqOQAXM9tStIYQ/XZJAOVs+T7FCtdZV0eCkhl5hCp2KVtmxak
brXhS94bT3UhqpToLzcqgzRFhs+yZpHOQ13qcpz3uGMa2n/yRjSXK83BbmtaqXct
nzprnIG2M4TfFZ6Anod6RX+ziQOU3j2EZ/cOZmep6WHhIhdjf4cgQh+A8UgYuFRg
1pzLumPKootGfneIxkFUXY+2yOPhzSIXmGfbpYBc80f63//Lafue4QilrE3hDy1E
tzSCnGXNhW6FcKxzq1WQKOz5QWmnvp7TZ9ItyOUDzWOgh4tfA8/Qkpmu8YaZaKRE
d/gfBaVjV6rTE/uFR5J+57g1TUqs1MR2AFegqWUYwo6TuBwCtG3QcQSvXoesq0RW
DDjeio7tNPa8gBgRGdRnk5pnlqN9Jo9z5lgrFfgVSD+4BmM/7pPFm0acBIujYVuI
utl8ePeNeC03ajBDeDiV2xtxrZI6S7mbV4RqqsV4UIChNhzNAfYd+UUw75xK/aZE
toRnFFEzvSQjNkz3q6yM9eY4pVZJ+X8NxYN1oJjuAXFX2/yJrgVDnCkH4YpBOwuK
I1MQLBwmdArXla5Q4s2ReBdJcxGwFcZzwi/ou5HSIu8f5dBHz+xnoIiFavyx8QPj
kxYhNT/RG0B024LsGgq61zJWGqKeQDuzv/Oq+MxT0hjW+LG/ivTe1Af4n65yepeW
/vvUwyH2YoHykuTBIQESDNHPoMKYgXcAemXSlu7a+Z6yunfUuF/frYC0KxOih3Rk
T1tcVQYd9k3Def7FRCLqmk89kQcYdatu37ZejXN/KtEJctzJgSByxc2VBmNrgYoZ
aS6fbNeOVCy+UNYx92Fj1a1riYEuIp3LgJURDFz4sZCgrL+QfqVHShRouNf1nNfl
dCqZtiuCvIFVnwUdh5FbNwHUVBl7cH8rF5zyskJOqx7t6JQgX5i66uMveJslsQXN
JKuRLb/NdCwgK8rljEpF7Hog6iHLBVDiyuqWe7FYOEZ510wAKUR/HE5U7lUkgV9p
mm8RmHZxqhRi2e7r8s7n0FyKuduqRXbnJ87oIhTwPViZ8U0rcgOZ65HMQUfxK5XV
wudMnd6FHz6uZTwmVEw5kombXNqk5k9I/ID5R7VijfW98/YBT8tVs9nuv8mbi6IA
rG18/gYtj2Pjqyym+Kzr2XXp10NIfBSGw+FbgHhmaYbmUIA0lJhvZDwUB/M3usCK
uFSAk69gPd63jS8S0VesSxYxmWgDyFQ3GILi6qT+HrpGGL11KXtTwISrJ2uyq6KX
mZ/N42VT93lxcv7CYU0kuEFT3klSBcPyPBRKsJH4jEEksmiFqBhIfiVzvEBj8GjX
+zEG8W11QCm2hAXOQLAxHznfnOP9WNjNWuEGxENEGPvmR9rkkKfUx6nDfl726H+n
VUZIYdTrIpFOwgiVX2ql4SBEPxUMWGhICBx8o25LDsPfvwfz+WEhYGWIOfEstWsZ
sL/UKKnIXpI2pGhsZEa+fnFoMhqUufJDoS5ydzCZP+KOchL1ipgL8GurQYfAwcce
XNo0mhEPkWFIxolrQOP1eUQPq1hYbNgAK/ZPe/rdldgBqfT8FF5wzyyNQIqI2QIc
WUvvvbuNOgYMuMbK7JqKwyNhaJxVBZR0HDGZv079o2a/ycvTJ3gh9wdA7cAFoYzT
fB1B92NYgpqcVG16CNndUBmDpcmT90Z8aeT/JQFUVQL+jMtMfpcMtHB5Ge2sIXUq
y5b9VGEyOEB0gWHtygK950kaxhsJi+5CDQr+0POEbFcJ6tGSxNrxCgOCCbDv1pW7
eeQtR54V6FxHQ+xPtprQOiUx3kDPDOXuD+bPOGl5mWauCqUCcRr7tYB5NufbvGz/
nAuwplYB6KY/exwIUo2rkKtWGsBd/wZgHaveavxhH78/KZzwLqiv/+7AATsqCc85
1NgdVPFQXh8cfZXNxIXQY6dgJkCg8EmNTLNzkjXfmLAt7416dQNKXfYdP78rRzhr
JEiCHmKFtacf2xZZz7rkalWB7xv7v7LPJiv5+hGwOI7MoC9vhhsOUMkvVSqlsFKP
JDsI73MeGSbVvF/mIBD87DebU8THKWvmdQGfxJg0UDjQ5eYnGMVys0qi5SQ2ePZW
FClTzvWddGXVcgN320VMnVvXLKGBRWbV7ekVaj4jR6EacjnPp3SDRRpj+3ykIgw0
Ogx/lyfwDdDrIyCcGMZ1uGbwqVyqtWaYrQh9XuqwNqJkilvcaJnlq+fDq0yUu+Cq
3DyHPxK4WjIPDf5si4urzGIQ4MWuWl4V2jZ/PcKXcU6tNUNiT2ObWMrdbfMusacF
JmhWUT9Yu1Fo45y4R23f36sA6A828xmkpm6ocNDHZXV97vUXRzFHy+zw50diE/1n
mGen8Wp83TiFNHroifk/ZjznnSdOfo0raiTtSIM9MWp4VLFmAV7vRecACFDCKWl9
I/oqu/oieZPv18uBJo7eNG9/SB2C0mfm4KIpdYQEMRs3/23zahdugg0ft5akNpRP
d/k+p7dQSytSlmNy2joiyCYEwiNR7DhPmT6scadYRJTarT3wyoSQdZPCxFIE8SDM
ffbwfEtwU/dZuoBhtEvAaNaJGXstJiUKXwwMqqeXdQYHKppXPkg6dIKhAsX4EhKa
3Ra4oCnEpHfxkWEIc4KzHl4ZvJL/5gF39MDVy4qbw/bfAnNijGTaDW+kDvgwphw0
s4K/9JL2haJKSBQyAiOeiwyYQ4R8c0zOiRlZIhe5ll2agj6gJkJXnfwrNtSDHigA
VrvnU4CiGuL1rG/dx9HVIUINDYograbi+4HglQolxNUctGx0mqQFvMKj55YP/m35
4dsgQXLJT3eAQ61gQpvsTGhGW/KvTc8j3sOn+oSf58Dp3qzCciHbl2qCN/B736kw
2CmLJfNFHL8u8i5lwikm2X+RZaJmai1YbGhYO/ojhsxe00lu2RFWFnVCQhhZDDeq
kk5bz1s4SwPcR/Jy/kQ/dVtd7OG4v12brjJDkGlVOP7WK4aSrKJqCNDXioqRDiKB
wvUaALzl1SchmZSIJjw1aVWIBFvbYCLkySW3yWUXn+oUQKBoHl07bo+4/T+C6rwB
eDQrOYRWVZCbCTYfQ3A1t+JzkkjqjgcaQ9N0y4n1Tqvn5CR0pEehRPTk/DdAkk+C
ijVRv1g3R0ax+W4lHAwhD4fhoX7JV9khFaH30373cElkAcBWJ5DqHrKGT6J19kIt
cOFpdWbQO5FtaAtFa6b3Q2pFzxdNUx+d99oBNHRRblsaPLmCq2XTMvC91yurDdsz
wU+oL/sI7qXLSb6MGnQEByIg7wFtDL3N4/rEpzSuqdVvG1k2Q7NDUjoMDMXyXxly
Lp4POyUW6GZ7RBlK3GwuWYxvmVUceaifAiujR0FGFHCwmzaOTU30m56+uMkiziFI
8PzuygFwhj5jVepKdtFPkvFFo2A3LOVZJdGBqAD90+Go+LgPApPtR5j+Uqegoev9
MGuMd5Yb4ZgGv0YZk/kmAibbbNBU0Pek1ciFrPZJxmFNlU3JSf71cjVwxZlMyzq1
ia/mERuPuPX5zM2VE2/eP/mdMKsc7uFE2QAlJZNoISdNtEBBTjA09CXr2OOxgOX8
WjhYfP0GlXa1k9PKgn3i/xTa0AcHQO7Yr/PBJ7FKiR0pM74ADVUhhx2oDH+0IoRY
s/TQ92sqXbA5d4OjvcTtC9FK4QumWfEUhmWpOtCNhSdCZ8/l4AWkigvbx9BJaVQ8
fikkKq2eN/x1FGWeariS2IKehoo4H+377G9UjKJ1UmlO1nWf2bxrc3onzEflmlgt
R+QEzcCT/DyPVhM3YAciwfhOOMa+fUJxc6PtjMoPUR82dxVwnY3hIUrZby/bGwXf
WCWTCtpfFyCx1yckhAtaEDLPYOo3XvCI5vNhWxuC402HkJ9uuJFGEJJOkLgzu7Ze
m4zKXt67zF7vWDqjNO1hyKBgeWC3S3lU2si3yXwj7HofSBU6egcdIM6FVo04L8EL
nU2WYJdNwM7mpEts30SROE+ZK8cYvB7cwkKXYYs5yVPagAXS5cN9fhqx3ISPoBsf
eDTKFgRaj8BlEbHzPybDIz281eneEB/LWRD6IhkyUO7StaiEhfWkS8X8qgiVhPzq
8v/0DpD1uHdWHKBKc8pQv3QX6AvZaQMfmock6F+i6pjl8nxx98PFWyQ/L0pNBnOA
Yov4uTl1EDe3rRj8W7nXK2S33uI0f7rRPmIBrYZOQTJ6zDgPDMG16finGibAfIGg
TBqKIu1Y1g0CUydVz4p6pzsz7Nff+p/7ur1jP6bEDSfsbQ/+CgYP+swJTJrbswLk
D+nUhzplSCwpNYsR9jvGLJW5T2WoX9Y2S+DdLiDF2pazOzjdE+gL5A+B4HtLHPGX
65MFkzsJkoEI9qm35xDge3T2MH/LqOzssrLeQX67VzCH9kRyfeErsQg9wkrdrz7D
SqJFFfjvMdmG64ZMf5FAfCpXd2PKPefTZ1n3ULwn2c9fc0XQ65iHy1MzH0pnuMYs
zLRGxO7W/vTWodMqeLyP6ZryjyBH2oi7+m/kkML0J6uaYI/xjEp4AJcuEqvb9o6v
y/oJxjgglMSry2jcUfCebarxc6rPuBOzu0DEF1SPvd6OKWgqhZgMEhzAZB4igNGT
l1LoswLSdEZau089H288xwKvUehyG+IppAqJHp5iH1uvmml+tf70/jzJ5dG+IHHt
hkGgBdqWgjxX24Je0sMS61ZSC76SRsu69Nc78wKmGs1Ia5RRAMudIgarU3DAOdoI
eqDiTLA7cjoru7CRB22UoC9nviJnmtmmRfWykifMquVtK53OIkBJI5sq3UbNjDSt
IgZ76BkgKYw+s+p+12gyVB8H1RbQsgKHCj+IHQSyiT9jQpSDMP0wcArmTCBPOZtO
hDtkhm+LAqhadUBUllZz6d/8teZ/oRbKHsr7Hf8UILPkPiKZCoKE7pLWJ6h6c5PL
qZK5jVjZnHlfhMHdmrJ5MQLffHb9QFjwYSshN9v1zkAZeZlgrRU5wPU5yj5j88jO
4kpFCYrEyr8FhkaK5803AxH/fFQMbmH6iY84M488fbwuMCzTF3gCSmE1ZinEiQej
hn7iGW8LTI8E2mwzFqOvxpAKM4n6icKqNOVk+lzaC7RLUETkv8YKUxh+J2+zmKMp
riMg53v6dJ+nsxdjyv44Mgoodeu20zGKt43uDY104iIQdgN/ZNVrY7RA1u2AM+8v
8jedjwbR430KnDt4EJKZMbtYuQqfT00MB53G295gK6le6216oAlbPU1nhqFsPdaQ
iNtzdcE2KNhBF//raMaLL8iBDYZZb+i8RILfdRl9pww5gH6D2LPOa+faPi67zJ6Q
qzyBnpbQ+xCOvVZIGYbF05KGLFn2mXTEVgfdTm8wPMWTjhhbJk6zOz0XguC02NXl
4WhoYtOudo7rRCNUGxOsK/5838W1T0Cgxp3hOrVLzuvlnuE34+A5QvMloe+m+0DH
3FoRmTzsjKL+S7dtwjPxpdudAFny5bcIG/Kw4MuWWkxP2BTjdAi9SbipyuiA08G6
99inm8x4iusXlhM3uTZzTaJffJa70jRRf7nVHk5gT2H41nIglVaq7+rNJrQdbClL
OMC/qXVukPewfb5Egt4kNFErq0Aq/B/Y1ik855/7py/28VZRZg/Ldk5w6ieWtjDz
6TjqGj4ESdTGnDS93n6xM8quU2DfY+TGlpqy1Ew5gv2WNtLanbWp3gDir8maITDZ
WzqfOoW6Q/+JEXgrcIyM441G1fpF0+vqO6/NLXbRADbhl5/o+0REyL6M9vtEF/Ym
Rn+MSK46Y/0BbUp+n20r6DC/X3S81ZOPDMGgaWXBMNlgrjOJtD7XNqnu6adp3otL
vp5C4tLzB5pjl2EfluP6u0QXhrmE8X8MsHAmKN/TIMxJKAjBVGZ44c0wG5S1pNvZ
hDD4L9oa0lDGZL1DtW06ugksKzMV0M5B9/u5swaI/R60Ta1KeZelasOWLU6YWk1l
pvAjNFz8zETL6TzJYSJ2FcnVIq5lhUQ21RjYWWa4Jcf8n3eZFlXKX9JtJon0jpEn
ncO5plghHVlKG7HoXUZWlC8nRutPF1xaPUBM8N3dekc8NIRj1cXOxtl0y7HGfjLa
1J+nXEQ6+DsT1DVzXUJjuBWOP6ISybEW0ZQIU/h6xY2u2h2JgBgQ5B2HqCD/TRdQ
LglZ6YOSJbtjQ9SdlRxFq0mszQhrnj63UhoewisPZnMFgs/B4o8yB3eWoJNWK9D7
Xz343ZdwwK0xKAb3pyT/KkIJPuO1iYRAg6wlqGbg9xvCQrkmj38BN/xh/qcDn9pi
Xy8Vje+nGAXNBSIQFEJ036A4Qj6ePW+P/locHFGcc7Je9583Iaeq/Qmh8j1x2Glt
6QCt8WKZIMvVJwioGDOSCRkngOidB/oH0EOs2UnFOsLKny1Q5qaUq3FyrUR/403b
djDIELNnY+gUhioB3W/J5vxgc8oOrNiXq/nfRM3sZaNQr8kZnxYIMcyH7eTKUWFo
6ouMgmX/ISF5oqxPH7fZ9bq3OfrJRUsylawb0j8tx06RAcUogAWhJFFLCshg/h0p
aQD+fKne5bo6tkG3Ioy0ckvpmjU+GbpHRbZ//zubU9MvkH0eUy4TmEel50bGSOMf
8Mwkthr21oF5J5Zw2t6KOCd8ICEz6VV40jdxLyTsSW3Cjfnd2qw3wXyalOXmWXqj
Ib1+IzHdiEvyjr9N339jPHCZ4iJZdNbGCgCk6+znOC0kbVK/o1gUyKnzi86H5wWH
Vh27/OeuSTDrUQHRZ25jiMOAE6bhyW6IDx72X13jlHeGaREWIkzOBuC8w/ec6zr9
6E1zokut8YnbQYUsweuI9QyGJNXkQPm5S1WsSCaoqsrltswFBnqpG36qj0cEOfvT
1+LUUJShDIurN6GIT6drJIfzJ38e7GMqLNPFcTAz3INOZmZyBvQOpPfsvbfY3TYU
Ew4O0Cf0t/VP9Tk6BnRu9xtRJjNqOHCOH4805dL8DasijSPha0I++RikLG1aOpCB
gem9qzOJ0zbVjq2HGFCwsX7X7GHLHeURAgrVZurXgHssLpcvZ3KONCMONUBBvgv0
qh/682ODZikFSEhqO/iZ7O+SB0vpZr47oml4b3PB64ZzBTY+6R6SvN5FuXbtksSp
vZSdTH9HkDSs0wJA3wjhwvVZfKdn8upFsdxEznDYKijOCnyL2eW3EQuiQ+66eIIB
93pYOWd0kjFN+dn9x9NcnvBHuWWDfsoOgD/iB8VG8b2IQh7zyELNxvjZ6tiX/eL8
0mD1KDMm5mYUl6DFCq0bA2ARetW9ujOgB/4FTcNIzCOckbIy4CwsZK9LqO0YFuHX
WGcD3CiDVEX+EZzItACKDIXzk8ldCe9Qv+qPxE1oE8YRNRz0MMTtwTcw4NWbXzO2
ivU11tyqcgX7uGGsZRT5t8yXA27SY6CW5W9etweeiJU+gyZp66NlpSA/VbHsgUea
JveC5UzPSe/EQQ5WAnLr+3WiAI0XJdAf0Xj8NphEVUMEv21aL/FcXtPGS6wLn4i5
OrVLpW6ildmZAqenRUmk45QhxQCaoEmjrqXIXkrwIeWadMk34Z2tCKKmb0sKss4W
eduOKrTx1CDWBns5FpRRV0cCM4l17cRH79PYk4xGyJd329sN5stnffegseMiJQ8C
vepTfSktdClc++cV+rEfhd359x+MuVma+4Mna+fP88oFadv8Eixpajd17Bezmslr
S2pb2uzvcKX5d8EFFowIqmkl5WlwAZ9GNsQajLFqzevj7zFk8JS8yTFaeuxNGHPJ
cGXpwdZoMyVX1u5oEdfQnzuWjYTbrunYkyUEgP4uZRIed41FQpvGNICfPHYapBdq
SbiVYFypnrwWmC6lwLL8KXVFhxxd78UPGcHAwCUDXNIxPzWwRcT6velFmQkCzOfv
WUi2tsFDoKP1M84u4PFmnATPDHlM5X+2jhrs/mWomaID8HygXx0acpw0kIqinge1
dA2ODc8f7E37NYCwxDB2sKR3gqC7aRgB/RSDb11BocIgFDdA6635hdrOUcP8t7a6
tWKNr7DRL4toIx7ukup8w9KT23qjtIDW+QSznzrb88ni5CNOxe1GgbIZ/PuSRnlR
0NCp/CY/1kF94YAFCzyhC4cwwZAF3IMCGQpofngJwBuRp/YpBh13JFFI79Nh7/kC
wXgMnkkI9qSoQ8rjcV0CNKjX3UAk4s5Z4i9gStjfv1daeTiS12pBaGiSylA9OOB5
AviESCmrvm7yHT7ROtETd5oNqbKHrcPyysWuariKrtr0vf9khHsDeydBZ1VAfohz
1OX2Bk3EXXnZTxupLyJesY7Wu9Lr/s5kqzXIG5XgL2wf8GA+oRFH/YY7Rv4wop/S
JTizi/WU8x59/z2axvsDXQjT3xUFbxCTgeUsOWPE6Cr/QOkrOYjjIWDPXWe8tbtR
WwL1gUyfW9Ic8k3bMwTNLnabYv/RBwjiAd8aOKo9FT/qRcEA9chWCjaJvmJHvIUk
Jw2qgdv+jkzrjdOk7J3k7nGpNdOtwVs5UfpLaBkzUNDcrsq4AfPsm4vDRP3Rdm6t
6R1pkxG7Ms3MBvVRuv+uMwQKjTOdChnK8CfrjHrIgZmf9+0uBQtIipOXYcz4LBLv
Q1ir9W4aBO9ufRaezZ8mBHB1NN+YxvGW293HBk0/C+GKjGdXVNhlWmSPwj2JqTI0
lm9TeJCdT4lOTYqHnpLpwpT4BYpzoZKXePsBWtR2Vqm+IubZLrwIfSgcLZa+3fui
fzAyUCHTtpvpRIlRdlwCAzY34qPjGy2K2VI4yWBxlJhaRA9LaKgb+RvXQWHFp0o/
VcJBqcYXH2UWHcCtpIQLVvNocFDvWgh1RQv6MVwZ8Yf6AIRunu1aWXFvRd8zBkKQ
Al5sUIa2unOMOlgMZsk8nQ1Drf6W6Iurn7aZ8V8DFF3o7TzyBbMqZRrpn/iLdLFN
NYMJ27raws1hKEgnjd0FT040eb0SiuDF/3xyxLj1sHc/bsRmsF9wAxL32bT9aMJg
wvxyEvw7mR/N0aA3x3Bv/eJqQJjjx2czOLgIhpM6R/P1mQZ6XKJH6qOLED8V0ogx
ImvwRfBctaJTGuTjJXZZ6Jx5LNc7iY7tWP5R+UszH3ED86LPgjzGXN6hPlwlwb84
qs+QRrwQ0D8UyqaC1kehRkj9foKEnRviDZCbebPRhpDHpVpnrhpzCOnHrXXAoUtm
Y9lq8sE9AmaW51CRSwxf+8gFQGtWR3Mp8l9ZIqp4rprOJ/2BQB1u0t5YIcfKPTYW
5retywtZDOplhXlBHcREvKMgIb4zB+GEUH6hpvgaLDO20uOMZB4D1DLf/FkA99t7
syjkiieI/cm+3Jc1o/rSVqQyNWIR1r6hbbVlrbS9p1XZ2Ol0kSxbjbLSmJMRKyis
j57GtFMC1CoIwx165ZuiG16rCEgDM/j92d78U8K18/2HYKPVbOwgd1bpma14xjzi
sV8A8Ok+l0Stn8Vg0RAlGxMV9AqEBCHn5bo0t2Cv9piBv37Xnyjp6MdmfHK9UZZc
fE4g9P/QuuXgKnYlpe5DfaFNT8/kSDtRPiwMGJAgoSVsv2+4dZhBLBzZXdUqwgAT
iC4d7xaj6xPXl3ULjDbTZW9I7sXH2ZaMPEctvdgZqW2860aKLcJ1RVzDAL8/8/U1
cL0T5+TYM+9zUquiXfXHDtRYZcEQsmUJ+25ZN9srUaR//meS0L3EdFSF5XmOdvL9
QlwL8PweBrTiWAT4L6j9YZAKPbqc/emYC+WbGimbzoRXLeo58ikBH6OgmIyJT2n5
rqlXZ6IDByNH/gohwAPRAHrMtaosEi02tHWRGibmFpJSsBafR7FgZ+pOmbWXrEwh
AYJQwIhqa5+3oUqn1DMucMERjUsXesLFhLMChl86U4i9wbJAMpduI9bHfkRWfrAd
5vnEnIHIZ8R03SQGYlaFmA3u5w5scDotYO9N1hcaaFKPhNCScNty5YQAl+P7F316
IU9zCQAISIwL34Vlf/TZs2/ezb8M+ewXnKaHg0EUJFuWUBi9qRIWTdYQMxZFI9in
Z0dPPE0shPnyq4jozvbmpa4u4dW78L5K+m7sd20GftcToD/OozPSf/fJbdYFodPN
zyGzDmtKsbxXLxV3lmWhqL5J41+SFV73Tjd1p/2fL7fsimB1Nz22RtN/uvrKhaOR
zDG7eMqq7+Y4z+ACX70j+Exy5jk3p+Abi/fRCacWpy5r5I1eGDMvoQlvdItCjEnF
GJDhusKmEaJ65e1iBuu7yfCzRbzRQjhiZoezk1MyIXafQTjSEtNkPqzxj7N6F5Dq
UbzyyehzyrM9hNZXtPozx/XZ7aJsZMIf6xqGgLdwKcqpE7FkefBDAGPAerXnJE3u
CvAED3z94p/CECvtyEz0a/ifWjydiYJEIEAU8Jmx8cze5D24nYe8hpYFFoBOUqNi
leXtAmHQGtDUFL4OrDTJvb6HD1V60OqEezTQ0EEoxqDYHit5GqYKJ3zEKbGaoNhE
Ql8aItCr/5wA/1Wgo6dbDiXIYqIblpnEt+v955vbyNRozcD+G0+3kC5p9Lj+T453
pKbPtx7mOe9HGY9hNvLzsrjOhdXfEFj1dAB0jcUJCWTbz3LMu//BZ27k9FJW2nPs
qG8PW1bbnlAuYYsKrgmkjVclQkZBTjAsZGPD4nExeSgcEMp0Rwya41nf2FMzpGBt
e/rDHj3zEAPwggnkjmd+fKAH0T27PniCENJUHtzX9zZlccNgB+17k3bq9lJL7WKP
kRY21v5N91RbhcoyR2tqFV+O0qk4C8oF4tNULTA/S/nkTaF9eq59YMKxKKlSLLNt
7qzyFLNQicY+/ulwmaruRSUwwDOKGsKKdF1AtlcK73WTORsmyYYfpoMLkhFHlQ1h
TjqSP2Qn6r32X29JvFVlkWLgfhu2s1KTaxc2kMcuYM4auB2hiHije/vEDahIvQFf
aZYp89FeGWkteyD8WxUlcrMz2dZFXPofPr7TEaL4fof6jVm1lz0A6e6MnHmoIOvy
oNKqjyYfPHcaqGW7mFlYEY5R20FVpB2wcxtYQLFv6CI3AvTKgbqVtUBYe8ihcQne
VO3xnR49o2yBlooSQAdppLml8+9VrCTCcaVeqcZCWxWTQN1iDUh8x3DvXswn+uHH
l61hdNuasfr/E7at/mOqG7mGH/xRwd74+FXABv0qrgcGiEN0OOhq7nOLvO5Ib+zm
6EtPKPxihiF49at02C1STcAxOsEhbTUCtPx5NWhyCHgg4PnNP6c9/4rhd/I48ldX
Eom7v6KTxYtTT8a6zkVbFwg4wsLOj5a2KiPc2tRSTAyOmI5k6YQQqc79d8sIP+Ed
5JSqqWjOxPlxYI1kejQ7YfKUVuCMXwiSpz1emthk2fd/lIOIYzydLAYL5Hgs0FXO
BuXrdHT8DAIIBAVNl/2aK7Eh2R64L5cNIPLcnOe22yl+Jd1dBgQtl+j3YsX7ErIT
C74vTHJf1QCNdprGZ9QTWqca8Y9XSE6KPBr1O8lb5yx2gaHp13nnk+4ilquVaTe4
x9FhOFtcMZcGqyoMUWsPzQnEJ7tqJWUP4mEjogkTujQJv4nuAHuT/6ZdiAIFaaP6
Ry/ahGN9S8CvWZC8I8KBc4lUZh7f4B5UTN0WtZufymFa4Ntqjoc0iYk6t3jlVXC2
ptjJv3gAKmGzObYh9zhgeA/hCQsOKSE6LTHN0OKDlChkfTN92Q6hhS9c6M4WMeJo
/LEbSKfVldsAHPwpymZuwpSYHn16oaqaPnAjH9q5MiPLExh1ZVgCwfapaYfYndu1
o3Bwd9VI37cP0/DtGUNuI9SxZ+3z8lEYokfR+0Iccps+RQScthiwMP6+EhgGgpvL
roAAJ5ClTCqsPynaSl8DBUZTAnf6rfFhBQ0/fbaR/0nd4m0BMYQRUNiNauzJxwmE
vQP3c/jSWlipMOQF9hEVU3q2W1oL+8f6cNKdlhpQ1I8hXttKx/3LeGbwWo8Yhfha
KJ5NllpEnORKHx6sc7kWJXYTsGqTJdfzIQDvFg2Ty5bCoj6/ktWIzqwf51LzL+g1
bFI73uYCwce2jz6LIJwCgP+pEFn7Hwn9DlX77qSVMynADYT+fAAPqje2S8QXq4lA
lIXP8KsMPT5S6b46vY653x/2E8OZpIgQ6AQjkY7ZHZAAJMTGF/PHUBi9pe9X341v
cGtoHI52+FWmYGzj78G8Tns4Tm2mg1kqNl3d26vnYo7UV8kAuq1xFIW8+hxIBUB5
ErOwgBPr2ZRY9GFMaiKc/jdCux0RuBn1UzcN5o216sFg9142T/kFbOMeMIM9L2rh
KfqFo0hcYGb68oVBAk7udjuZerrVASNrSdojWFauo621SB24D/JXg0ZcWEYtsJgg
wLjvqRTXLCYHHkowuKGK+wp3Zq/7/BBD4hE7R9DX/4hT+s3VjOQ5LxRjVy9TwrrF
NZIC5LuHwgsWDbY2XvHRaDU8y8lA7WEQyKpxvA6WB1MqVwoDKu7LOYkQV/Ll6qKj
swVYHJ5z1tI3NyOR0hK+yMoeo5mI9+qxKbGlqRgnQwcoZ1FCxcXQ9sLKr99Hcgcp
u28QsCfD0t85xIGNT4G9zzWM3WY0+dCZHxxhkAJzViheN+eyQJpCNVEVELFHRLvK
+zqL4PB56aEDDp1vydv9UBgFHoG75kfnPZwrxa2KpNfSnt+AuyhXxpldPDBGstRn
kq92Cz2D81Q175sKMVxTlYCBpfLSe7nP20/JYcXfHYLCkfhs61nq9KtDujBx5rLt
GjyWvOeekk4MwBDpn26IEAvzbGKUNiNbPnI0Nt/yuv77GrB0zlLz50txNZoinUK+
LUnwG2n7GbQqyemrHoS9R4iVXyaQyCvzi5qsfBGDZnScVW7QVNL2KpKIerJKqx8U
wLBlKV05ic5xvfPp+CBs4ZcZ6lPOX5R4sZVU7nXI9WpFY0MM/rnklY1/LMVTes4h
YE0Q8V1yWdWXkPQDZhAx5NrnY3uHevGD3y6vO1BI836mSbvbYk865ne1DJeHovLE
c5fvlXiMV1v4jGTOMtY2LsTYNIvStA+mpizlEOd1ozcFudsA94gdpLruIUTp5aSL
TY/K3xqEDJxOKywbs3wdECFEIMdY6C3RP7vYJbtbtQ1tnp7+vQWGqpOCLP2jwYV/
q40L4Y5L16gL9IZvqLaUvpf+oBOTbqrX4UmG+gFNxZ/E9RTGLKuGNKaniuDSkRDR
zXxV7QmADTYl/uaqhNhss2fbi6mZ1jqJNLx4oBgwjs/12Zo+C6EkeTox5NYPpWEw
EEXEzYBRQpmZD8+z6By0lEM39AOKalJNvRXap4fKkgAXEW7Hk2uGKmtgzwpstJ6E
MegQBO8MZ3WIz+ovgsuIs09fpV030iGblEIqPbwi4goQAGkOj2ZS5iaqhMJ2EyU1
zUtSBcDkGOxELTB7zC+nlxKEyAFLwVaYau1LTjiOpMKd+IrCnfelshzpbMuKeYLs
Y6Dy6L89h2Zxs7+/y6AHVCM9i488s+axxlW1gxzDL6JTn2zLuuOeq4fdFEJWOCUN
GsscMSR8vfGwAm0eqdb1uwpgiMTH0nW4SsZQRApt7aWBzweWAZhPsE6VZTZPjhVh
wq75n2mBGteysdB1TaFcH5v5k5etQm8QguMVvA1sbXHO6cWD73aDQ6NZxjAz2Hpq
jNsyyh21/Jq7c9N44eIxskPYPG4rrRmI0vKk9qUV8FZFfpaJv7TzmM9OhWsSN4Sm
cLPqfhltHHlLmGnnA/0+RbjU7osPvt4I3x5ThiM7I0RVmOS1Q7PJXEFhbL4Al5x3
DHCgWKsV+ryR0/Y/ZyUEErZXVvG4WUkWq5WDR4qF1bjJwRspjwUxqSpjHo2ruASd
4j6/+76hrk1QspgLf1HcrLlRZCV5tYmEhyl1MQp+LL1ytreoZxdNOtHY8SF3nqBj
U/FB6HTLzHYAOqoWucffSlTWZkJIeZAmuPeYpGETznYE/t0Ql/E7E4IX4K0iRtB2
4lHjvikztvrzJArFoTyRmXxd9tygiufSUIYAGqK6wTz8YazLbiGPtDSXyIfaVBo7
SbBqgCSrmHkDEyZftww1Tp6kpcWqvi/srzg7uN6QQBHuRMAcnEUTM+UpSDsMdZT5
wQQZx3bkYi4h4mZxSPZCRYpltnjvxPtdGOh7g17sH2uH9FCBHiYk9+qPDSNL7Nit
akaqkkZq/Ff0T8WYv7SKgTtRjNqZMKITotQhwVY133rRc/86T50Q8tOmK7eIZfvS
wuMSwMlkiQP4wcB1jcWLQdlpIHeWy1Q/D/Zd0yDGs9ir/mFfwptSRHmPQOFZIcAI
vW7Ul419UFYAULXHMkRRUm9F9ADiiBZddhKwKj08kJ1YM1n5fAMCsGjZl5BUh6Wz
n1ywy33vojf/7fHCvvDdfxLalQ5oVFwICO51w86NhRdHRoG/ajGuwKLFjLR2waZc
IFaiy7PCkjr8DScsf6lIQw8bCIP8qRSqeMoLFKxtrfkcBlT49qTF6pNY7dJYeruN
05k7fFCO2xZrZJoGvlALLB6sSKu6UC1v4DRh4QNgLWmk42YodoKZXFc59l2G+PCh
oK8oyPpIs9GeWgdp/I4IhAKtXV2CJjuxqKz2KTxnS6DBKwop/Z8bAmIxz7bpS3cV
YBiKg//XyEgJyaNSP2MqeMJO2tXZTkfXm/cAku/Ud5nlauaNhyPVvKnpF0TgpPAS
bX8XdMSSW8Je9lZDJ9n8DlBJQ2afRz+un+gSnmkAGKLKvoY2hoVzV/nSv7gp8K4t
RXm72wbF2TwWt/wE8I1E+oDEz0VWwRMu72empMdOEV5SK2laWLADOaARxsfcwwla
dsbp6oHvnYUJrpmm759qMZTVjuNKfMwU5OQUiI4j9KSAe6PCuZ+Rd5jROXDfpYS+
Pdb8GemfGHXF7YMDfPMUb67yFqq3/XIID7JqXiJTFWKWH8TSK5BSVr4oVFoOmmuC
iRo2BJeLliqH9LjJzzOo63SPa+VprlEFq2aX0/LwTd5jxc4QpWE30HFUW+5dyBUf
ZE/avMgP1frSnGS1yI9Vi3iRNvB9Pml/rYu4XeN0Th2ayHaPQywxf+o7pbrQ2EPn
s9M9Y4NPwMLogsdG3qu2jPKP3HrAjO9jCjXeY6aDvKUtLoAo7j0UGVzAOcKSi/Wd
0eO8FtZFQoJMGOPmlPvy0ZIynQWTLC4dMN15SqUnxCIDflp5eIT3nwIhgMhbYTYY
917qjZBKqW7y6Qxo7Ipi7dgV5u3jxVEEwuzQ9m2dijXXFb5QAvZkEYLPctvEKmre
EGvXNVoaf3fSb2TW/H0AaAwmu5o4tSm2uE59av5RxC24jlzL+ilWsD64GxQd1ol5
PUurbfSkSZDAdxjog8afBmMART4Lv8Atk7DZOcUdgT30JA2W40eMKBMnT7ENvv3j
tgN5K6lgnFXcl97b/aej4Mgpc8EtcdPSAVsDFJHbxXxGpTB0vyYIjFIey4ZTOvLt
ILIVo7xV/cT4ar4KvIPhf4VM5ATFzcdCEtzRBxRsvX3wjteIpSnh2oUJcx0qLfem
lySz54HjlYFkN0KJBAM9ptArDS22RbCb6Z/hEkgP+fi5wSt/ByI5QJOZY8GKBRhk
Wy6Lh2y9a8uZzFMTO7fcayzl8Mh0/DXRILti6F4M6lbnmgdrmvs7mlhGbm1IU9Ri
VXWtz92VI2PSqfp0u03GvbwCISFR5v5/a5oAGRnPGuBXf17vJjy+hDXjt3tkhGyM
yEhTKTALsg4CUWD7WnnqEEZUjs+W6bJ5aIB1vgf0VRzNN5JQXdkhXE0VDJa+sIgT
afev+1fFQVfVcljWAuVuMAWOFHEULM224jgczfip/L7Nm7JYQcEkS4UKdp5WT+NL
tv9WG4ON/0Wo/cX0BVgaQEo5h+Cz4L4Qqo8+xJRg5w6ucbt6iQ79PLUN2uXud7ZQ
SSgEvakKTL2poAQhsDHvQ4xa80k0AZBKoaWQ82uE9w/T1jgIJXUvjCJo77mvR7hF
XJ3wJjWMX+hK9X2IrSq88I30K4r5+9Dlv86v+tc4Hy/CMOevPG1SzWcI6IxRJsaO
xdw9LQjstMj0a+A7IGVU0vPP6PLxA8WYNrW9UtNbzGWUO8VKWC0WkAPgXkBVzu+R
H9o5iULdPLJ3iZ7TEJQT4hETdnlJOumIrV46k/g/6xe2vpCM5hXT5umIYtZY4f9D
3kt+tROm95JWLCFEJ3UFlGTj1qhWgEuSPJ/iE3logOBf2OjISnmenNxqKVKWY+0k
l9nHe/ocAjAmB+8dwWOcUCCfQ4lAhIjWHIDGe4QgfNERPmCeehr3aQ9nMkQkEZEg
NPAeH6557PcvKai0D1rJelFrfyJlJp7AgVKfhwxUp8357xrRdyw50SFCB3tc1Y01
PulxIz00gV3dh8htu80lkWkxG/8oDpEYc4/1MU9+ZVQg+aRYbYIwOOh5tPW4zuph
+ijjAgnmRoVyXqGn+Stk/krlIV+g2QN6QDV7Eaywh8qD/PJieBcDRSa+OZeustFt
jAd6xRSyQqMIgmFNaoMVAejginiUCStoC9Be/6oCn3+uGe5uTjHa6NO/eKzwvT0U
UPA8DrTk5hvT8zrctqKNgzs0/CANb7Wx3SJkFixmfmo3ZpWKYFV8sdTQAivM6V0E
ZqkQShnKCaLcIB3kJrInR6kxPv8qABzlnbgHQy3sBv+YocOgMuSG+xj3113lS9qx
G3OC1PfAtC7HpFoTLcH4Ab6Yb6sY8FcSy/g+jWnZxlp4A+ZYpEZFkNmgqXbeEsKD
J56mJuf742mcFpKvIMGkrqC0RCTfQ1SmlnM+V6XtXeO69HCeFAaSGx/Mgrurbqad
lf0DsZSedldmXPzCffLXAbX0Qq/AvC/nSvlp9uX4FLY1PK01BFFB6Wu+vNOae1Ez
Ht3hMQU1t1RTBjscGZ9u0FmVhuyKMnd/UlPqJOW9keLfYQYLDmUjoyoE5i4F/yZi
rXZuKKgsUdlecNuP+A+lt2r6+HglyN2Hn4m6u2Q6XxXehJYirzU9mIh/j7lClc7l
jF68isdiQV5L4FoFxCte+P+n8STfz8vcvalhK1JeEF1urcL/NPtWJSyleftte5X9
bZKN/OujP8qRzm2dcGwC+AVIjVsnPDUhRes5PJyWGHFetTZIvKgJYdvbSUk+l+JB
sQ9evXDV8/823MIy7spaz+tOFnRZSVXCdX84//METdx53biqXibYBrA+DX5VPnZO
2M/E6eUkWVAWriScYygbazxHPD586E4Oq4AWNHHulFTMoYmYPR/tInXL9MzClY8V
/K+18qIhfFBqmMOBRenyDqNAFFZ53taPjgJNrFRkZs+kDIGnFSC2ftzfaM6UU19P
pJYCoAcO6FyQCk5sM6ZpQmqAWvfmwGUmr1DrZT1HEEaP04/aN8jf2Q4vIFTKMB4I
1t6NQPyhx79F6k600uXyp9juOGQX2cele7O77gXg5gBxV0PbVI4OWwBLE3KT6EbZ
ZbW0q7VNAc8XrTccROxvXb+3InvFGv6zmfKhL+cyEApTv7BRZ5oU2lRu9XtClM4L
7STBYcANBVZ+aOzfint8XQVRXm5FG1JWBSV5/qjNcVPaBvYOv+cFc3M2l4Exb33y
OKuLX+BJV4h4ax+ec3+lHJpZPnAiFa56Z1rzoIAyqqtGlo9R3Bf1ciBtQyZRLz0Y
t6Ssmo3ZvFdTLGRKQgpjRErcAtjx0pIGgTAT/DeWA6PSzz0SPpRjIpliqgH5iVPs
HsZ7Fh8WfAC0UAJFUyHjQWBtD+rOfVIOklaCckIFe9C249+op4kg2Jk0K74dKLSb
n4ibCEBivDUgFZ8l/vVONXy0LGvT8SV6zllNkzMJvxTtCh4IXviYFhvGpv+knSzx
wFpJuw5/vr+vtwxzRdDvy4Vutfoc7/0bOc4OYHYes4YQY9/T1lPZYdzaTs6dcWi9
Pdfd+kmfqqk2fcU7MzOi7Ct8hf6Kvb7HSJOqg74dcCzq6MqsCJAYp80yHXey5zOz
C+9ViYz9U370JFNHRkApAIy+xkNRhvufKyRAqAmdOQS3kNSaqjhmQCPRRMoUEwXt
YoipMADT9f772/oafvDSROkM+GgNOsFDDCETtOc6mo/lmcDsJCSx0aa8Zb+LTcg2
AOn5W/Kck7UxiMA8/N/ZUUbuFaLuqYqgAbWd7lbNci4/wrMdMcUY5g+rjX2PJpOD
pQ+e6rbrHxdkZrReYhyETBCuLgMGCOWCm6tYFuQWOFelC9lrIFl/uaMf+e2rRWpS
rbQrTKSGbpGYHcwnGx+smOrqExuwaJGSXf5VHsRphjn3OUqlzaZgY9q6SWS5PAww
P8Aw8vtmr4tWIDVFzTuLwKXR5mvnjDrxzQ6nCS2VdEObksCwDxVh0daJjK1KZh0u
Bb3hsQhbOZuviYOKNCD4hfwIM7dPNUJTaSeCVX/7Gw6Ve3d/3uiZxPFWK34/YSOQ
RxgG3R8qK4lbi2dwhCj9Bcqhp8XtXAzb3w3VQZ85+TCzfGsp3c6H2xCAdidO3WGT
q+HsDyZveoflZqJ0xrTMr+frP9BA9twnmTWihFqWFMpZQ1IuZcjO8bxNzZsUiqVH
zycm9mCnBOlz/f7e97Kdsj6mDLM1ljoH2zdtM2DjoG13MLH2qoIWf3o+YQw+aP8U
mEgpB9LyKeGFB77+yPqBJ5GCyMruNV4TAFRBNqX1+tU74/F3UgigJ9xlE1dGRc7E
h8J8j97rPeSBynYurWES6orrhn7jg9ljd1rUruqGmL6cPbWdngwDqJfE8PG0ivJZ
s0YbLRunxOr5er1j9lRTrzEpfxlmmunjZH3P/njZxPY+z9sAg3PJ+ghjU2DHHVZj
vi9Qk9FtjyGsP+CM0ylWII7iQc+0PCENTUjsfsHs0+Y02TCmujHTb1Cgp0+amFTy
y73on6c+a/gAMtia7+ic389aR6CxEtvnKGneF5KcGe5/8RWKmAxh8chLwQCVPdxx
nd9V0c2OBzVgY9Vcx7qfh13HcrXegqayW4As9FkSrFJv/4FlACzHrQE5FAUPRIko
tbVh+eGZhXsz6+wZ96hBOlW+LGoF/HpbXythloIsZnlUdyEThdNXMDjUkRaPeb2M
fkIkqP+Ni+FQcbC6ZjUZMv7mfppzGYyk7P1I/+zsUQ7Xho/KHr12cMSZ+YrdjYFL
dXnQFicIAfnXLD/zqqZU3aLRSiY3DS6QbM40/WN9FOWpL/YQJKNx+r4kcqF7yD7c
VERX7GoNTrUvec3VTZZlQs4G8j8WoHvO71vtez4bZif1esZcnoYCMxG81Jnk0v7B
Q412IgpV0pGXntL0tEH9EvraomoSEl3X1XuvsBeDSwoLzImuX3FUPu9Xnznei2W/
KrcFLZ9Obeafay6otvxTtVW3k2pUajnC5jZyRPPqZfK/H753VM3JU7vg7FT7zS+U
MCaj8Ae+DagHAJQoj3w/rqYq/4kAvBCta6GvZHyD//1nwbqFjlPwJJjEFK2NgKF6
tOrMp8aleiZLYta8SFst4uQn8gL9aX21o751dW8FbBf/OgcLdi6NhKcr3mEt7CWj
JuBhIeJSM7gBjedCyKf8lC8zkBssv4rqKVhNYyVjr6tgfkKmEDW1MVx7oshZ/DwH
S9wgVmL4b/C1UfLag9wXSEcyfrJWkMdW2ZaA7vZf2pY1/AZu9MBWEHtapZMtY/C4
HCC1XS1TsQ/vw9yYNq5thGy6REi2X/UE/9mxgI5ppareqwqR1MryLeRLBVu4Rizf
oA9KzS584WlIgdqpSpAhXnKPLbwG906WeObwuq26y5Cy90SWZ0449ecJuN5KlD2W
Th3Lo7vU/YXujIH03NU0kuOj3mhOwvUPRhPCQIc3OzEEQ8hGJX2MJQoWMyjs/zF4
Vn7SrXJeaAQT6DVWtQLXTgTTHQoSf2xp79v38+APEpp+xygOfDLOY/D3iUGvzj32
1uFDzO2hy/f2T/JixYXstguX/f0dFa/kzcmhWJ0MpLt8bgAMhyUm8B69z/oZ7vuP
zBwsMCA1tem6wVdIMp9n9Bx8oSAwrWtdG6pn3dQMOgbHDLUDZinjdDJ08bAykNht
mlJucUYCw+7EdIKqm9zLcKG4R3TO+hJatA1qDVwI7wDeZAyNGeWOX+iOF11cM9fL
UFJWsXDUQtmUP3kcbrpnKyB1mj+QfDUyxjslaBRXZXWJQcAAtSsUPEnromY9bkZs
SYkdikmbKy6suXbbjqyQYV5tPIBY6mu2VNadhggXvBRHfmm5R42hSKPYlXwf7Tub
jFIWKBzCiOeRAnOldEYb9l+S3lwaflDb3lXv+zrvmvuryYvE1hu9egwjwBBrADfw
6QgXxA8UXxApMbsRfTBwBm51OHBgYbxi3omNihWzwEitP2atqJbXc8XfjB+7UjuP
6fDP4/jUvwH2K/ZCm6b1bh8B+duGImKUbZYHnvQSKWrbDGFk9RLPVj4Z8Ac9ZbKs
7nkWPk+Fi3PQY5dydXB+zWgT4DNfKZrFBz4Zn3n9yfH23WIoyuPyy53QnhMLYoCT
arDng91frHGCw57vb7qZIYcD35V0POv7rNFPCG3/uZCyE4Ef9hs3SaqPhWyjuiwF
83ZJBw3hpuPmcnGP+1e1+iODyQrowuHS5YyGr9WyAvdapqb6tjk0U+iu0YHlS6zg
/FnsO+0xivS/K6o0Wyd0EWf5EKaunr4Z3gfHEQVJbcxNOGoaGF50Pqmcid6OQKZ4
BLv6POvJUXgb8jlEMmacVxnb/iVaXdzzuVe12AZUj+ujp7mEbuw4v1BYl4EWyWIZ
dnj5Qx12d1UvRRMmHHObODzUq1FrJVXqAUh54KqGLABY0121FQYsu12d/hRGDvxZ
iscesTB5KMyZfVhCziVnM0p5IJrAYKtdCupIE2dsep/6lY2Vz6UoEzSWikwm2E2C
Px5PGMj4k4vPRct+ZuIOC1QE247qJGY+4LXPYhUnxvuJctybWxVsJBeGfVAMmOYV
iiMxCBGmd1v1DQ9+avyptthQdaKPBM7HQoFgOw0akKmOBRd/FmLEy2FGqFskJQVm
nLwp4w+r/m1i6BAIgBj8JsnAGAdzkAsFSZx5FmPbmCYekCiHDWeBrxXbYm4w0XgA
QYT7f1zP2q+yTu1xMPy8N1r77PqoZYskD1XJgkD0dI+ZbtmgnKJG5qM7VapQ6KsX
zYdDf6fO0lWqqYUvz6OxygQuBN/JuW9PZ2aXHayfLPf70cn+0SuxrISBfd2oP7Ib
6aatHtbEIEMC3qni27KwgOdHFZV9t8jcpfNpXcvgP15CTKAyAw4YGQ7UQZV4KEkO
qWR6DJ0Y+gvhtP2UsJ70OxCOvDMfYumU4F1X/+vFa7tVlJW9NcyQuchQpNjmDL1A
WoLkgyfdFOrKBv/cLdyJh4KhjPZYwhT1zwGqBTYmS3E7cVXw+VbZMWt/4mnSr+FE
sEOj7Dk4cVaWbrE+p8Bz/fCWnibqd4aFtVFda4sjzh1fMm+FM+aukShLsNMc03yE
Qqw9QVuvl43QwnTWtYaDaYvV446K0xlq0032Ng5UQr1dwW14/osUiyhPktEoE6RI
YVH+TJBWTjqXOlk+OFmMdhKcqa9ztayJzT1uzDvuoILae6FgPuYnY8RqgoWuFXRo
gcUtt4nAHREEetl0R3QFdFfJEiT2wOe/x79u6geaQebT0UB5st7pFclbyO0Mn68c
2UTBW0HoiGhIcJ0UZ3msOCeL7Gp2Rvl74ztrxqif7/SZYbXoahFNw2oU4u2xhFEO
ve377tLSY6kHHara7TBLVvprNL9Of4+TYkZUw4t63iYyL2y3VXcjBn2G4C3OLEEk
a0QJlaaDUTq1DbDL4R3/8+znc5VSCz5r1+RhY86feEzx4OIhv1GgX/I9M/0UpWdV
ZRQCdYnHF5AqFAgklpV5p7D6ytBQkM7GRTp9vE9ZyEMu/rLrUpYQuOhdgHRhR9S2
+K6k130T9ROnP1o/DcNeoanJGm67AEKG8+DUuCHqSk4ZnnPhEQcGo5ahnEO9Tay6
ude1l6Toeg6+58FbLNpQAv19EfZfOMHp2SuG7RCfywCnhYQtV5W/EoTk6D4u+uLf
2tVOYwNuGPdzJwqpHpRNhmrpvT11m9/riVNe5y6nVU+F+j64aTLQP32kOPynlFDV
nWH4xTjthFLQXA0NdUPmS9AODV+zKXYrq4/2UKzfc3jrHcNjL2VrAqMW2CxFsi00
NuaqjEpMhm6tKVQSenJ5TzGKtKbfbs2FtZGvepUIIS9ZNL8ArGQJJjuVxdrkVj3Y
nU+tI6ZbPKuDecnDqLe0oQh5EhxIfOQi/r+L+bwUTqDNXTMmgI73v1XE225yW3rr
7Jaf/zmx1EiWS1ZDkZeZosWFKQQ2ByehWnt7ag4UPbq0wFm1jmK52nSxDhuofdFG
UH69jzD3goGjK94b1OHVZnsIID0l1RGSqVnbOoxx56+4Yah/Gnx8cEPCeF5MPmDO
Z10CL4bTzehBdjn1pRCdI9fadcbxT+uTEEttg6/opf7PcxtZYjnvOVQITLb8CD1g
2asvMNmC9PnzNT3xs4yoBMXmGIZvGLeauRW55k935CjObLlnHHxZbN3WVIVpEBFw
RL/DgZ7xEU17ZY6IXdpvl3ideTxrBZ8dOWbDOF8YgxnGfilSD+0bGLzcLvpFV7gM
ltxK1+2n64O0HdtTZGDphGLfXcQv3jY8NW/APtn7vtcIUkPEq7GlOOyU7jCws7an
oNhLg5SFfdvaMzr5P7hBrEydJfQE639hwf+JIJXlj4vGR7l5W+MhBYNW99RQmTBX
Z+iRNvX/pOrjQ+I3f8b5DetmYOhnwDT5sBrGhBt9hVXMovWk8hWJy8lNaoVJzfSj
9FhnEmg0TJogtjvgO3PgS8OlHeIqWWeiYnl5LTC8h1AxmZEp02G8H3b2lH5bCPM2
tUVTGLcN0O9ke7m/OhaPDfdIAM3pvtF+Q5CjsAL6yLH1ZK1+CtcfKv3UDGBoDR/f
zOlgnLeRTzaFurL+L3ekCnlcve0n8d+U0tTXsFRnjLAQjTgIb/OM7yy8dbtJF33k
jPmzj0kuoV9RIP00g5UPri/1jYqg4hOUz0gsfQfcGMY+jWaTkU1tsh1AfRTzWb/F
5e0so08fAZfRvvbmB3ft9DjZbvDznpdHFfxmWFtvuR41mmahKb2hH2Ps7VgR0jZ/
wB7kaCEGkdzhDcMuRfYQBCusYurUfPNmVVdePPndZreT9WviLwPRGADEQlHCAKOV
tByuwgNAgtSsQq8qXdehEGw0A9Pf+vtJW9MkWinAKFM9NBzO4bgc4rwxVoKaZ1W/
mFK3toYAyfPggu/uazae0/cZ/KC6C13KT7pqH+eZUAEe34eNJfAI3VPCmC5iipxE
TCKtTxxsU/NRvMHF8UmXZhjjL8wrboY8wXxM/yPUG0hhae1WMcqErLOoN1DWLJLz
kE3U1QFENDIC1ZAWEpBFnY8vEq8+q4gKe3sh/bewkECaBRCycZXgZz4ljJDyX1/6
ltx8puNiX79diEtCDFPRmZ4CIVdKxfdU5ObedgNV181rsLeCDSZUTteZQenWEUU6
S9VMWMv/w4ebi1gdfWth8sGDB07dE1ibukOHXUWu//+kusEbGqWjIu7p6hY62KOQ
A0nccjjpx30UVv+4MCwwQX+mLMcpqUAoKmnF14ADzt1jWUFY5LakQDuQ+kbYkdvH
SPHA5U7vCsvEBqY68JIT6xUNH8EWqLFyKdXXuunTqoEVjQeJlsGm1e4uUs1MDRC+
9XLsVr/++xKGce3A7aSN6fJu02zlsQuddESJU5d01LYVKHXj5IZRvAs+bRiQ5sNz
N5jsICsKd2R4Ijo8jwUaqr2GFGC2boaO3VxikPZBepudLoWFEOtJ/TGOv+9Hfe2/
mg1iwX6TZVoORmkSvcZrbwQ2OylPuoZ3Ky3JfcnnIKpE7QxI5nL86X21FLjWkkA5
vMg26rPiP/x+BSsydEhb8Hew/XZw3wRmJCyGlAGQhBwC2pTM4reD2NiO3ZjflqTC
EXJ9NKalozxR5jhYEVA6jT54lHQ8mquSWGz+icktNkJCfFbVDxYG11fCuUjrsjvZ
nwf+EQO1o8hmkJZNdRT3xtpZlmw7RDqK9yZR7IlTH2xjtQj4YOrBdXszdpU6uUZL
CAmI+73HC3WwCLJuVG3JNO/zU28RSJB7a/K7tY9hyg0TxzjlA/bF1ivAr2ARujyh
bBf5IDxEwgHXWOA53BYjGejRRj4ufJHhGIG7/ybKucavopqeLTXd6yW2S8pRyWpD
Zg25UGDUpmvlVCcA3xADawWphPGCKD1SIFgdWBilt83Z04H9N2zq2Dl6sP8MJsXI
nikDZLkK8uvhh1NSbNbYksa/btScR5iwN9dykxZWhcHPw13VgBbXDXzFHIM5SYFY
TfQIbgQgr6SkUScJ4gKt28ODbPXKLjwZkEVs4LWK+zzdZwt06XEpiMumhkw1aDgy
RCXlRJlNW3A/Xi5cHF5NHnRA3HoXSSQUwQKPBX4RXfaFpj3A0fQgcjtHTJXXKUqk
Huz2Z+m2h+RHqhmIDF+yXur2Wsn2imipb+cu4y9lg+RpzL/+NGNfFwKntgMk9si/
VEBIS7v0Lb11LXN52kxOtJSjOg8fSsIiH29xEqmeoyKW1S46X5endzRziSZ90qPY
bQnENCl/NQ8sEhEDytYGnyaXUQu4tiLZLqDl1AHXafpZcIfMuqRCqHeAFRq5Xo+d
xfHNobG/zCJrAUhW1UW5GPILc/+JZWX7MAdYE8IqFwlHwSBq3BAYf1PUSfjdLIxE
/OM6q4bAVxpVv5HduyQsRTqc+T1vN6acn7Rdv+ipntqsOw/nK/DLlKbJ3geQRLmz
qSrXomtbX9hh+3QkMWIon6v1vs0IT5KgKyKWdOZHOAXWbnnm28Roi5pwJYRi4dP+
uQwHwmzaEfNmbMC5jdKwUaiMlC4NbMccEypD/b1a/XXenjuNnH8iG2lSaEwwYFZL
mhPAq1c1nyKfOyt8yUCTM8vMZJk32/fbBfDLUtWhBSPub+PKbnmv8Zz05t45pfHh
vQKd4+vTmuSiXHXXa9bxr4Ow0xdZCH6zrD16axHsbtlFJOrbBlKgbdiJOQhzzzUl
3i9yfj6Q3cKr1/MYcIOXSvPKpfTPxZUK3SN22xLkmy1QBkakT5Mn6qhoakWVtPw8
v4mMAGbMMqsgj08kDVZ/Xt37/VPsW2kn8Wrrs0w7zSYHww0fu+4Uzc+7zrR0bUqZ
568jWJadNK0ACJQdW+wv92w8cbFZTTy59EHD1LFFsSO/0b9ulVxIXTmEMiOBqyAI
wiMnxq+vtd169DbVb0zK/4Wv6KeU5uQT+KvvY6L4SGpKvpcGz+gUj9j3Iwd8GgLs
JjSb3DWWf+J0qE467kmD6t/LkGU3rRDNuAnVWvu+VHHe1HkBx6Uz6sd+XBq5VxwI
tPn6iO0gQR8xTZtElFu2cLGHDpXHkkegwX2k5scfYmxpoxv0OILmQy5shMNSya7T
U+C7Cy/LngmE5pmICAO5eM9WO8qaqEC4znEJn9PgTNoctmr1NBj34D02PGeIg5jX
U7dbk6dcL9yryU4khLk+AqwqavOlWG9swWocHl06ZLbAPmyaCJoQjYt201srMKL6
wJFu5c7fyAQy3pFvkJH7EWYIDj3xOy/Eem4kLUdORqDC/4gWwym7QP6N6gZjQZvD
xTs91VXF7y2s6j3PpqBnzlZKkN5r2DF3tNKgc9MEVCRJ9ZNCk+gBd4FL1kHEtRQY
qESrp8yzfa+NDzyCZBm5tzrbPvPiLdQZQ7Uo7BD9ScNNdLXdgsRR+uDzwYBz5WYP
jgKnSYE1J+C74hDBicwpBs4fZKMO+BYrNzofjEtn4RdKvlknlc1qoy/jwpRwr26E
6q6PO9UDIzFe1yp+mQkqM7Tjtnp09g9tWGUwGYj1MZL+H1QJqZVG0fhiS2fYaztx
/6e44KhyY1lxHugp2v/MfaGfc5s/DThXSxk72WsEzkT5tVozj3u9giAfVC55zpYs
EkQRGzzkcV5jY7Qqf2oey9JWNYV97QA+ZDdS09suHAsPoCv6R753yoheiGWa4pN/
CuLar7v8HQZ2/WeCiSsEr20HTy930vFQRwU/R6m2DHyQTaD7Jsd/onMVemQGJnzW
JRrQ9go2EEjKHTkjw8wHCP9XAtRA0WNUVwnANjDhZ3Q1Grpvfv7gk9mOysTllaB9
PG1jyLHi5HFief3kTCdkmguhTc8IvlNmPZ60/ARLyVlXedSlV38mvAIrFwDV5LFX
XKcrW65aiHax/kCjaGhGMwjcUUhGf1fAirSq8RaRJXbGUeHySzwenOg5ABB5Q7aE
1it1MaZewT12BP7vT5XOoYW8Wg183xxT+p17AL0c/6ZAbodGY98G4s36czuYYO50
vBzQ+zg4BeMAhnH1wI5RkAeLRDCwgv537ngVHgsoUdM28MXCa6t+FRPOc/FeRDe7
yLFWDXUjhrrPnjC5l2R2BA3rAPEOvKGQ4AkqODljLQQXQNV4TKCPWTu41diXrNXx
YccpZb/s3rLoVrua3QBWWODFHvO+RwjIAmK508SobzX0G80jkniS1AEYA1y5B00t
erdpLT3va9n83eDW8UqOyTPG7kkdT+pJP1LsYuhAkkXuSTk8naphF56sKW9UtuOJ
6fJRGu2pgPmem1Ogzz2nOjIw23FNjpTlQjnZh75noD0nrCM1qmVDNV/jn4TDyRU1
RZASirC7xnpuUqP0OuiKQkAqACkvh16MtU67h+IkmXXfmWP4R83OCf1K+oicAxz1
SUBW0qL1eOQzPXnBMFN23grWCB9suiRkYYxRpWClf3cdYQL7cot5TjeVKXPi3ipz
yMVH4S14T5qW4FoWUPRrxfP8OXrbp/tYAZpWz9LqzGQoe8wpSi7Ar+moi+bmDAx1
9VxTE0GQKNzthwUYgFXolIZHzRcHmp3zPW0EgqtMAfsXkwRPpoP9l/g4DEHiPflk
/ZBmUkguYvOqlzkaVVPU/PNc12V1BRi43QpePc/davAiP/0NbXUpZzgpIpOF7j6Z
Ld0JU5+nbGd5QpyIkhIGyk6up+7Dw2i6yxlPVtdUW6NgLBBH4RNh/v9igMMHbjIL
YS2iOqifkp42Fn7RuJmEsJTXkCQZcBxgE1vGEJTugYd7zMz8dIqBc3CuSW4RGder
OYKlYcBAVQkWTFvtwRAxynCiGifiu46BxwQyJwDsXaFdDv+uAWC3fIRrY45KaIXq
Ct0aEXX2sGTiqekHL3BprrqT6t1GjCrrEnYCqJkY7PpzADyHbH8SKrDCYF8DLYsx
extFP2Cfp/8OP/YcaXeJiaCQy++3KgAdr6Fxlxf7Nezya38tPJr0RvQdh0QXR2nT
9qKd9y1QcB6a9VvUxWmSKMhRSEHf5Su0hMEewdqkAIRu6WeRzo+YJlwgVzkicVAv
C+E5kygLHC7bTRNiNsiYLEQYKjjpiIyp3qD9xPXPkZzUDT36C9+8LjaHuOjz6WuN
Xz7+32raVi5x0dfWC2dyP86tKgClv/uZHbp1E83zeMcuACpftkHeEkN1hhAhoA09
UpNbv91A7O1QDTNXi7NlkJxwdNDfjOdbeUT0g5H2ZiRpknUcNOVD9DDY6bHhtjIe
GOyM6mBzExZKWGxM+80Gdy0KvSjKajPZx9rAkmEdxl/t8MFIbi6ky5byquwDHCvu
W70C6DynZpKvVfvd8hfLFwAxlCS0J8D7dSypiSVaYtJhQCzvlk0tyCbLhbXDxVvl
JXVzbIdaV6U7sZI8ZcwmcpcBDqW1WG4YTCQIhqxkd91o0IRKdAzOCwtyroHt4b8k
PzRoSeCMxBVmp9q6Y4M8Bww3qBhKhspk9eye8Z3ej8NGl6l0rd3xFKtzVBWvDJrw
O/YxnS9EbgLCas/3tVwIVZmVe+vH1xBqor07FK8zhC1uG28ouNxzS6AYjWHE/uYE
d7KuwbYk7Z0fW/MB9EcgRmE4v0zFwzv23oIpqx6yQoqkjXLpjmE0ZLXrHd+rGnJy
XDPsNjLoJJaDTx32rl2ZnSQ4d6P0/6+YT6NEveaTfEvIvO+HwdQaAW+xkkIDSRxC
qeII696uaTVgnahBC4U6F1Z/0dTEqfalpR3K/BnX1KnqaeCk4Tu7jXa72cb5OKtW
w1794pGDb84WKWNGy4KQrcBKnVVIvYOm1qm7KG3EfWWtd0HIIlVO6k4C7azQ4BOx
qoLWgW/PJukLT5pfow9pqtJi3Bl2CDPqLO8AJf2H2VoXTbIfZpBF5DZ+7klsLeEK
QzKhbgfVDyt3ZkaWiNJ5aH1Gbqn6YEr3hrAwR6pKc5OPGycof33JGViq+k4IiiFd
Qn76G1xYhfzAFNHq1HRVzXOoSwaFnBa6j9YIbBlduQPw6xHTwVGLvAmw3o+mbtTd
iMkhjzIedsgJkZuyCTdGshZEFTU9iLd1ATlS0lID/MS4N3VgFH2/4iVA6fyNXeYk
C2XgQTj1fNzLL6jLNCEmoZmpY75+ZwDJz/t8e5H/30etPyqls/AK3pHT5TTkLgc2
an7vQGpa2j5GqKqngGY86hrxPCrLKxTyFMRHH5zNTmlGU10WMJkna7frR7ooPF7V
GTIm3YOo43ByT2jpOfDB3BqyLUuL47Ode5zkwecZfylkINlb6HTunMN9Q4pVOCUe
WB5CyPxR6irpJmLjGqL2oBT0XIYqELMICdiVXNfqouHJv5yvaarI/mWRocATjj5t
FCaX50M+sB6wvugLMVcwDrMVI3tdMPCYdGmGfWJtN0fU9d3OmptWa6AnA0eMlOHB
EbHMtdBIQsrYULih8BnkKwIbxuJC38JW6OX6tYGLV8XmrhIfRW/0kCtRBRn8VTt9
S1RH/jGqt0BJ1Dr/Txt15c67vZ3dF64hog60G+c5s9yNN7xUkoMVP/1ThmfYKNn3
ftZzNNZZZ0WAGKt37O4u7oKVmmAT+hzJSLZtUAbY6FdtqGHibvwoTayIfiquEWYK
RHVB/rAFn0kDvXr+V11Nc/Wsx/4sIha5c8SeeOa5Gj8kjev0qYuUjiJ448/fEomX
C4U+N1OXJv3MtqW5q1m/kMzl7uBQCHQJuWsgghs5A3bdV/jjbJHfK1u9XOG7u9fY
qlGLABcINLlDSoz/lwi0mOPYSqpPFLL2/DsonUgKS+cwk6u+yiteaZXv6Qz033N6
ZEAqHMIZXV+d8TziLAQINgiuy1qjBLjYBuyHbAdqmx6emcs2y+D/mFnYqUNFc9FX
Qgt4aQW3yzlbRbIC2prukc9FuDRJlWyUYJNKTb/fynAVfWMewIMNLFCVuiOuqdsG
p7w4RkVuXfYlVY16YfRX3hwTgFlTJJkhv02Jze+z3HuZYjvWZ8ZBXJfphG5Cs8G/
fk0T72fc3axXvXJCFn1lxfR/szH+WKxU4DwE4EcQMIBeymhzh8hf5FRIUTk0H8HM
kXGeKOoiK8ZgGvidHCfiF3Qfa1mfiZlRscax4phohWdWbybRIdHU5RPybIlu2lqM
0UWG/JjYS6SEOe2wiIk2tonTUYCBo5HWQT6+74Vn5zxnP0g5xs6AR42xQBVpqB+j
2mCz/XT2m7Xj7VM3nl5SchRkILiC4+zs0DCKZi8shXtpWwO/+1auE2gTvfKvOoLD
tEpdndgfD0agr6AzHPMqnhOovuFlNWxXF9S1fOVUpKw0OkvE0C7cPeDQsMrqpwjB
MW8E8BB8DA6o4Mfj4ABwYLj83TiLZWqAMEuxLLqwowbGZYBX+UdITvoLFVG9aVsY
CjaXmSdRsinbUP1IjhgOdCostJV1F3yMbQqRZRlCGNQkrB9YkB5udS6udeKGWWNj
VS+JuSVcbDQO3z5mOq5iBOxmtpX2dkP30bpAeiNKkujcFZMBMRfMRGuKq3dqAemH
wVOuFb7kU9EYVuqhlW5oQ0N45+Qmz9I6+EA/yLR/xbm5MGvU9cPb1RHK4LzUpFlT
frzKzLB4eJ3vkrUwjuj57FASX6ayB5Ib2zRkngq3oT6ygHR5AS5cTlSbn50/ThK8
oLhPVD/PtI5AEnFS9+t3aO4IuqaiFgIZuOHcIMgLe22ttHhgK/Yed5tvOw99XLo+
cyV4QRyjjqiQo/zqrW53sPeNTkdm0GLTiKUQcklXyvaGWVgCFsczsq2LJBcptD60
OwKi9+hscGI/Mf1UISNykQsJ3+fFhkRshyVjvSpWYk/0fWcfW29smg25CeocenTm
/fEDhBYlGYnENCmS/ODTTPUTTBa75Y8gWKxEQSOEZb+cvd9vyfatOKvuR+1bbwBJ
nrRSj8X8958KBcZDOSEZsrhwYQOT8lr/C+2LJRhc2eQWF7e5TEC4QLuOXQn0lfoa
aWiepMZYysFYO67rwNLdzS8SJGCVwnHmZmp18wd0Kydxk5M3dRgnrojiYSOJJX6i
befcAckMg2zm6T4DC2cY1f876hldxBrJfZj1uVFF3pOb1g2ZvilE0pA8eOb3F3HX
fAceTPdinkgaHDOLiG/lIyT77AMykOmPGIgXySJ57l9b6vVio11vvTYpcxDDqVlp
v/37auzRWEkhTNm2SBndWWnNipJJqlkbpCRsyoPT/lWyWyCuyTvExHwYmnZNfJBS
hbTz//xE0Z4TV3suHyKnypN5RooJC525/+h1+AHrjc1BwcWoHK4RgGqitOGxdSlp
4bF4S3Tg158hz1gf3jjihMKMzXKEfgWvCDhUZ3MB+4QpobFWQcekDH5owlQ+rlwV
cJImeaaSsORCJaGZS+i6dcZTAaWtdMeBJuigO+WFiG9636s3wSGGEvanmCebe9D2
qFUxedU8A0bbiTwQmhEzjchUR6TQEuOyF45+65ifjeUIC2lruf4D7eXlCCRcnsm2
015YwCCoQgxOzZDc0N7aM//5EH6SEBVgBaMWr/YON4Mz/faYGxQE/zPjOWVrGES8
uOkSogpxcEGEw9Bxj0kQK/OF/urr8/GpxuBSUhQP5pB9YAuo15kXNG1MqxXHH3Br
51Linxn6D7NGeh5s7ymV+is1WE2MioPh94mDCiIz4B3jU1SCS4o3pt15/vIBW7ar
83CXy1VK9izmEWchwtRqs8jOaL/URsznVQFz9wQcmQeGCYOfljfupHp97popKQkL
ET64vPa51dsMGmrj3jvcjmcRgL21bCEu1v82hnn/3s6svAWOtIaG+xtgwO7F+Wxx
PBqK5Hnw3fpHmY6PygaqCOhxxKkouzPpjwXZxLgKaPV+bR95aZXC+a/lAfmtwNtk
5hJsBgByCkIoaHE4yFmMiLXilqWLujsKeoHIoKEkUnJ3F7Vpd9n9QfVyJYaCrLf+
FhZK8ihFlabdFFsNddb6wYviReEvlliycTb1/SmlaVysEwbE61dtX9cbQULGq0WE
x0phB03dHS83u8ky5KXJX01jsxYtwhMWcmknCZfBhxI0Y65FWHIbt9+8jRlYoSz9
9UVJPBROqIdiXoE44scHPfG5Z54k6Kq+A4vCeme/LLQqP3e5CcuE990HPflrnrba
bT5Gnwv9Hnze3wtpiQ4K1phBGxwyluvvW3WfEC2tzX8m4WiFZo7O47vM1LRDTj2x
aUSE0IPBp0xTrfdXNW2AO+yHAfv1VZYP0dnH6IS7AgmtFc+8B+R78qjLaKAQRGdr
EAvZY93FC0C8wSDQgxgW/VLPU1DoqCvoGxs+Rkw8O8fb3jz00nBXWzPC7FVXrhZQ
CrcKosU9r4Mb74Q51baOE4sdu+32HxZJEj/qBjNsOwN2Dii5eQD2drxnk8XAfoKe
GQpOBNqGJMlolFyrRKcdfpM+4g5nbTALkoFN66/g8Sruq3OoSVXvkr7deIUAxa0j
LVkesqo1KBmkNmmy//xt98tmGNqyyXMrRNOtGp/fo2PgZQY1Mb9KAKERGtIVGA4A
BKgor5DgUE4Mp19q+rF3pLLjaJPKPsGfMx1zA/+frAAtVk5rp+eboP3O+Qx90F6O
RrspDGbWeDpXifHIe3gKePQU/oeeeBJJ0sfL1domQVeexUvrb3rwaKPPzpuwr9+U
CJ/3E+VhKHRxWMHNFLdvMt7Wp7bFLE+oGNxWPfnMXgXapSH2VIRyVFvlCMRat7b+
kA4AbgwX4hQYCtAuQgwJ+I1hrY/2EAyKCUd/8miTfXvkOveuRiMUmYce/nIquzw9
QVoA2hKbCejcs9R02M2VuWlKBJNfD5LxrdUwEJC7PzTxtq054RvoieuduUiP0MNS
ArHE7oRGtw6hf2Uo1z1VDzNXGg+PLR3QdxIg6a62ICrl+/tELsuSc42wJrFLYz0R
/DDPU5Oi1AT9XjG1elVBvp+IunxzWtNtLCWwv2pWfoO6ggwYJgIKmIjZ/NihzE5r
nL0vhBB+zkYqsmRQeV0v/Nzv5KJL+x1L4HYTqOZQwo0T+/WKpOF6Yuub8GSrAj7p
HN4PDKlxBrZgGuGiIz3XeGbCxxSpkXBJz+PDyciX650HcTPxm4pTRdIsXHNq120O
eVPlV+aiAhGrL/zI2nLRpjrtfaPeJJxYKABAh2njjGULmN5qhFP7iu8/+lfkUQbA
IKYcZ5459cWPN1+bQgsw/z1c8Hk8Dikve+E/Z4OWm4hbpJWB+iewF8Q/tabyoJjg
Dy9Qo9t7W0ZgRLW/o9R2JywrjvyYJ1axSbFf4O8a0puH3hmXY7tMl+pDMWHiFUNf
9e5Ut6imHFEViAmhW7wkCEQHiKr/1Znntmg3e9mcy3f/MbTSkxtM1ZIKxzGpczwS
U/CgFeLQmIsm+GCB0JIGPRdT6LqktsTIrwzpTTAUnGlHzWOZX4Y8XEv7+OD2uMPF
YFC/3pU+QvnPpUPCuWCTsN8SgcMWgoVsWqrdW+RUUPmPguSFGNrv/d/F2USGwxWz
bwD74blcqfXq4xLctEb3U00GsJQHMpL4iRA57KqBYxBVfz2GNYDCZ63NA7+HCxuF
1ZBYW02ykiKzLc1HSfR0WgMRqVTi9wn+ek5/o6ySGP91ofpa1HfaQKOpvYEWehhA
a5ATAuuhPXc1rg4hLgmm4jWyZP5VyiE+stPRd9JAJJjrqUKqmT0Jvpj5o+YQiaFY
rUxucYWDh2Ur5IgmjFODs2pqQWf9VMQG9S5yeHN1Uutviqr709bk1YFu3fhLREDY
yPrMBRkNTxMdkuz+d8xnd2/z5TD06R0RP58Os/wm1ANDMLjV30IuezGjLqlMcTXA
tX/f0bN+hrrkUIJBMiQdbCEsUOwhNU2SOk/bRQMb2O67K+sbV3A9c6Jr3KlTSVPn
vt2fp/cc7Kej1sDNiUsvDB6eJp7XpLC1+P+fzdpVObjImg/cLDTj94bhnVch14lZ
3lsBlxpFZWs9QqNjtZEi8DRQipkFaff2D7utyCDEoax3Elg+rIfJ4zDlHF1Vb770
lIiozWVdhUa+Xkk6eUJkzbgYwxWQxemS8snJzdpH/mvVWZ3y08ZKPDspOHjfQklt
X9Slp5yOD6IDKRNogGHi6MjH1e2x97HMiHu+XKKdrYhjl0lNDsjzT9KZXQh8b8iR
RnnqZ1gnEN4drwDSMggiTqIxXGs0A9VxjPFf6aqGC7L29MaFDJ/jNSeXZ3+p37or
j+VrdnfdKSMee7tqrALoMNWVBdsOEKjR7yODavC7hRd1W3dLGbcJkDwL3QmTYcVG
hHSvCQjD0MWIy0lB520Bwnk8S0TDjCeNr0mzskaUpsG4elYs3N0HG2tb2tzvHQRC
RynnLrIGVo5OO3yUBey+pErN2IsfH45vzKAqm7TFpHD8hjO+fMiOxbprIxgar04K
W+z8t4Yu6lX50iEKbNFYq2Ln6iLPxtCBiRGcVOn6PltCzMJoAMDGxRdW7hRM+rdk
OkGXcz0HnNX8wGs52vria6ynGBv/a7hMByWdoU3HH/bef0aXMklxeYyj+HnxDVG9
D9V2juEoc1vHO4Djoq7oSgn/gdqqiXES3+zjWfQOD+8qxm1M2GdxWKOyTJnd0VYY
2/El0veAg5OTNtSoZSHuG/ztX6koMXOYF3GlL/FXvtfIT83mTdcKsnHMDMlcb7+w
jCPssSnky2O4d0pRcYu68afoW9b9M4qAt2I/4Y085O2W61h/1bMdGhHdWoGW0mH/
eQDornSGhWlv/07v8OAxR2Bj5rCxRNXjmgpj0Hj9ax67zVkW/MHCmP3ZK+G898bW
K5IuPYzmT0lzxIta227MksxrAaeJ5H26GGV5SwLoDlcxykSPuKXWKGylGqk3rveJ
ozFXSKeV5x9qLsS2Uz/DNpR/5iqTsuuxhCjo2VgpOBrHtDjN2397bpJyzBddx1Hs
CCAW4W68kN9bYRllT5xUINrkAXyGdsERLRhbD9Dc4srEJcNABLTFN1+EvlnU7aMH
2eHrM8Q0MJptGpPa18N9DJ265aaIeaxCv1zGuwfJhvmEzgH/DdhJ/TfR1NPmNn2s
JSfAs4Bkr0EF5aM+CGhgFmcRrOA3p2UIrAVMYTnMbsi8f0vVkEpvYo4RpPdOUtD4
d2OkNhQJCR3clgml+8swM3ASO/gQyixLCRRBscpNRNnQiPBhQ/bcVV7malPOW0IW
IZ2xQxjHdfRcjb3NTKaa43fEX9eruRFWRI2GBsMyVNDXsW+GcXcWVo9fitezQrmj
SEA88tTqDaSD9gqXXGkskAWI8NcJ8RH1v0nf5AfmdFc6Uk+3yFfIpqmtf8mQlyuO
TmcFlecXgF9RZ/UFXj/vDsKYlzYz9V3UEx40zFrDxI8KBddCTCI9oZ8Jno5623Gp
0ooYOWqV7PZHazJ7AwiiiyjKhISqkZriNJUa7tPBm+2XUyWIvGrD1yb9QCvD0p/S
i2chx8pRsmaLWOaRMU1MmqhU+Suw6D8L69M1mh8vyrjfz1VfQJRTAk8ZlkhKV2EC
0jXP7kn5A/LfK+A/xhMS1e/r77d8nbIAccAPL+MEDkB6LQQei8FhTo4y7dW+WtOu
HIJ20FZ6ExWYO9b47evEKqg9pSQwD6mk8zULYdIq4c6SU0qDm8yxX/dckhbR9Ymy
+XFL2xh4crqPEO2rYao/3P+lrTh4HTznN3Rhik6CK9YRWqFnMe8U2W5GOnLzI3Fg
+tl5d7PjeFCqGBQK5DUg1jgYuKCa2MPfQ/Z4M6Okea8dhXaxaqVXqaVasj2Sh2eG
P2YGVYlJtlqTlIiPMpAghKqKSxflxea+nsVmOMcjEbePzsciAg2zjtcXg6gMA1N+
sQBYVtZGtefZ1F7AI6+wBDvoGV2bICeZdQNwuPyd6TNNDwy9/v+cKXKDC9iga6ti
M51OX4+J9r2jqewOaGcClYrq0Q1qTWuyV+i2tGT7QS6Ktp6DGH/f+kCQqdABTjFf
4PSU1npWWrkpOHI2qXVqqjnDc1iLQRRcHgJXAANG9IKmJLXykgZmuLSACwzKumaA
IUp52I5yXVKOgJxuDKdbybI1bN85X9OjHPtgIL4yNe4E2udwkCoPYPSgsRwRoOFH
amlvMKdAap8DX9GKUFsZ0ERifBlKAmrBYm/nbHvG3VRCyH4IFKr1dEEuwAMANBtI
uVtqWpLP05w3WCz/zV1WPdhpiove03zLVPYmflDFNguwdqhCSjqnhys6TYgu+Kae
0Pd00VE1uVAuM1Konw5P5myK5yIEZzG/lRpcU8MvwXmCiW4r3zIpjfdPW68o72B0
VNuaowY9GBlxxxQvwmsaeDCMP7oYNZdDcgCo5w3uGFcnt6a5+ZlaA/EQ1iFPtZpm
eC3Aa1+YPsoZLJTL+L3iywL2tE6cS9I2Oq3uqX9fl/G0l4Z0jJCrhoQf+NxfGV6C
K523v8Lmguvru6zdQtPuBKth+bK8pOnJ1P6mXuJt6Vs9HrtPlVveEl8bbZP+FQ3X
k5Lbthbief2Chf9obRa5zMGPFWgVy6jkjiP3PA9IBvHNcrU1ykqN8WWlfJ5nYwHM
6KsecsXpgV/xxHGLx5J1nHjtWJFjI0yUYrufNWJ6yGiAIpQNQPaJdRgJFJC3SXFw
piKkZUhWj1ay4vp/F28RSUZh8YgpLCGQoRNcj02WKChq8p/aQ9QayCzMXX3HYeNZ
pjkswDp378D0lyJDitCu3u5nBUBxb/RdnUWwvdsDIy6qIZVcRAYEWSd59qVTcmEP
+gj1Nd9ukVUn9oCKyLdw3Ad/7Kvrd0MAAj7X4YjYmKfUoz3ck58UKj1J3gWW1td8
HsUcbDeqfrAFu0BWCQ6g39hz939e+icPpz6yVa7PlmNEQ88pmfYg4C7qzeYwgsxa
q5+qhCBIZSbm7XqcYJbRWEkUxZWJOSKFekPeSwb4qO1SOJIk/DsvEYT4AIg5uhPJ
7trJhJhNq6v3L4lIvWixYuccmZQqRHj5evERS1OZR4ILw8C6iGa/Vm7DPj6wq2z6
xSEUMgzmHyS3bit2gs11qAto8f0iahtJNokuuh3LhwadSitOdba5yrm1ObYTJFDR
pbggE7xJ3Tq7NjlvuNmGhOYLon7WuBIYq6UF41EEuJ07+fZ2D+WCh/KkjK1dqhlU
zmH5jy8TaQ5a3+MiXKhhEr29Dq7uc7IWbIxnQyGg7PTmtEKPdDtha8MbEil/BWDC
2uHuOgzvHlj8TZNpbbPxJq/ErqSa0E9/7N/AJiqjzcEJUh/n4UQjh4FL5ZfasdAH
tSUeQsQPjP0dYzb7mt36unkG7/yBs/eMAqRDegFbeCbku8mKGtrc/25xhJKuMOzW
GOn7oskEAzy8aY0609qxp9qLySXbJAC57/RAIxWcJlXqwlUzkHX1wzsjnSxfcE/D
ifTXfyfawl9+vVKWsO5XNKW+GeaWplaCFy42cEyiA+5BtJbC3DhI4BCtuoDFvnNY
rp2cI4SOm5OEnE424gEW30QTbNxIotipr+mRTee09h0vEAt/puvXDnIhV4OWJBxq
ACcfjVljB7PCto/GHxZYO22apNGT/+4tf83X7G+9FU9Op70zYwww1i3WnqcvURw2
Qdxi+vPnc5HgGP1X1pmG1pSWD5I5CGSeEN4KbethOWbxhLQRCsAc2ohfyS1+MfBp
jBNP6zW3sHW1LM5Z8dJW0ub9VfBHaac4bgOe+PYaWg57mn46rmc99B+dndtRfoOf
yWmLbS0Iks0QpQuYw0mUtAm19/z7QSPJfCDD4dYTa6B3waP1SV9dv9tO3eKntMLp
UYji0tvjhid5o8rQ94OkLiz/WfWWRv0QVaWhbENqmTpZ6KEzk64qq2fKyiiFelsI
KasobDrK4T0Pal0NzOZLOQ4cv/tTMAwa5OGMln8VB3mSMazN+fhaUNvekIrLqvEy
/pBxUsvN6VkCPmY3QKInnMkJePBApmsjk2Ti/wwHXPhVE6URHO9pu6/smLdaVF/j
mNFSyy/IOAcCM9BkFOVKvJ1YxcDlpxNiH5IGiSW15S6VaTXFh1wEWQi1+hY3IZX/
xDQHVxndnwWXjU6lB0rx0KMwY2c6OgAQNq87FQUVkLExJFiz5+RVXq9518fLECEA
kiDZYp6Gv2KAhxf4F7fQ0GtcXZb6BCNg+40pGn/C0malRQsaAnZ2/AABJTIlMljh
Zg+TZzbaie6L1MJ7h2KLp3c2d2V7fHvVxwC+6g+18hyhjkja01lKYnltDiuzU2fy
BQbWPM1uScrkvr2wqhRs39vfxpAZERTDWBMHVYUqW4DRqmvkx7hmKcvr05EYcBUw
+Atbaf/AoZ+YWP+g1A0CzS6YoQahAcKg+XkEvBA/00JdMc7g4YDhE8lqIirdi+KJ
2ocND5BvwoJPlhPT0O/AzEojh6YwmerLah5Xxtkg7wbxg8D7faSsnwtttK9fhMb7
QpZdFx7+B0T0NH4oHak7bj7x2XFcTBh1JhAZGBOoL0MvuUvTsbx+ZJpzxUiG9e/M
3vRnYtw3SIKO8+ehPW8PSp6GYlY81PkerwuW5YNPAR68mR3UlLR+m4zWXWGaR3Uw
WLMTDLofl26aFBbCZEUo6mnpS9OZazZOoViR96TCj6xnoXSAoWWI/sBfgdltFlW/
bafnuXcS+IROxCWCXDPDO4Z2W9rG8BmtLG6XgFvyw1b7UmySmLBccUjVDMxyUVsL
KM80+j4Es5Ri8e+LV8GTulIb2SgU1YLuKZrTXyGP4G6j2dLhsiHpOx389EpdTvIb
meQZUjEsMvfh0nrg04BAtOgSUUN22vI5R1smnod/hvABHV0qN1SZechKU3tVxRDf
kIAsQqkxQQwAS4Sc9sa4OeZjcUb4H+gRdS+Gs966VsgiF6rDuqLjO+6JqU2tuH1G
bcvZCzVNVy/H5xQUlUFZSY6cGifLY9DQKoDwgyxYx7p9tIpo+WqeEyjJ3K4ayItj
E+HotSKQnIVxGAbqDZB/0zs7KGrbvYWWW3ERJk6qDyn7Bbjy35L6RwO9k1UHsqFe
ifz8DI9Syhz4UVZdWLZ1OdQOtl4MlRV/krbxA4fk3Mu/Vg28iQ/WZJmKxCjkkSFN
QpWPL79P4dy4uGdAEwIHcfH4yNXf5ENuJ1RmKW4ANKAtS9UDfTwcJPBBo25U54WQ
m7HMn3/FwAACMX9Q/hjWVdnE/KQIt68Sycr4kFzCTvTd9Austi/3V8gphWOW9fJi
+HQR+SIkAv3hGDNmI0k+QtMTYyzEg+Um/abG3nwHtK15x07HwynGBbV7Vf2BKj6G
RvPhzgX7mXwsEE+4CDG0cJAPex6YCEua7K5cfm4JKhqSmYHF6M1thK7bsNqJ01Te
I1znNEopfIFYxLMnIweW43npKvmSceOjQ66Gf/Krcwce8jzQM0KMx7NMfQBj7tpQ
nbPt5qUZnUbx1y3jbPks8FtK+Du/hEs/SIxYG5VARwHAQpoYlKS7zOkxWcOJ9AJ4
8FWWdFyxSmAEysgnXwGGNs4a3VwnZqpMPwqSre7zJ7zCUachpElQRMnzRUAc3rmZ
g6kPgdPlDmKSA/ix0F8tTrbP+QQUG56bb+IeUuGtR2C0arFl8SoeO82dwCuFmm7b
ok38/1zlnb7RPfv+P4lIO+CSTb8mGgTSpBe7sdsrnqQzP5/hS0Vy2XXDto6+s2qT
7l6t8I1mPvQ614d/kGDD/Ax7ao93iA3YUSzAAJfLBz6WVdPFeYZloT7eipk4Zw6U
LDmdWeQ6vN0o7amYp0g6BsNnUS4nt+BydOOuAksIkwpRyLCzDFqSbWCW53N+8sKp
cswP0F5ia47CUuuJWJI8girxsGiFMymj2nVnXyoDLJNI5QRCExOp+Ir+tL8/ho1i
cqb1yqhZpcEp9rNB3aMQxT8cO636J8Ug66dz+nRwG7vxjDMhefV3Ka9WU1KSznqW
T7k9CZfK/lgolKUIptK43BJfWoY6u8Z3IODqM7oVKi4kN81sWtqZg17FMwX+jOz1
QJ18T7FW6pNhU+9WwC8wotiLM3MXjT1KHcgLH7fArXe5TxAl2Y3Hsn/jgl0yrKPw
L7MerX7k9aisglaRDiqQ/Kl7IlUgTdOvwyC60wJJp3OlO7dwVzJvvxSzGwmzLNBi
/D4zJ8VWwSfe1u4xWY5T14LT2QOxDborA5My78/g9NAhIeKWtQush5Th68noB4bh
Fohqi0YDLAGL52RXZrA1jpsyFR/yxUYbXIgJWmpc0A2KlZn8HoCH8QhZAA4SpWtt
PTYNJ9wdADQYhX7oqa6TtIr793pQHwKPEQJP8RwySS8winNuWfUUkttk4OQD2/xH
53VvUVTULdMMkcL1vcRh8yS1/WA6YNfVWcP4PD/fvAtSGw2tCN1RqtwRp+UsgiMU
gNuttVDedjtnN5jWq5U/8pHPD30Ad5Cxr1h3QsGgQkoXcBFAwITLzNLrq2tRhDo8
9NZoHjFaWqtdFPHrODJGDAGddYOFpd/ZTJMIT2cRqs+gtEij54aVYWTBkgpFAoGv
hoKuX/kxeewDba6Mj1oM4KooSPLvhXuJc9IuN5VThyzSX4PA4PLwYN92xklkceop
LYwO8YatqIb73+xPPm8roy4wcxnhJxhcetqgYkUhyEb/GpTELVTJHzbneymRgaCu
8sRAFQiWIhV3YNYa4JvjAVUIQJXzYfLqPaSb7LKrWyXA3E/hH+YJXwaPPXvv/x0a
tk7tI3gUVbSIAgpUYWUsZuaRKBsA7boGnKPZTR0QnfNsoAz3vmEepK0SlFXKotOr
MUthL4ePoitNX7Fkzd/Pb/CaYxs7c5s/QG2dDUBZLc3kQCI8prDkMRCRWBwGVqdw
+bCTa4+wK27s/rbctLdd3xBGYMGp8qf3qVqWF0vWj/+r7T5hsQ9f2PjQn3l6nm7M
EqED6oihw3tDnlLtUdnAUofqxOoD0v+Xdwk6WucXVULt7I67Wzr0Qph4nLkGMLDl
slEQ9oEXDjVu73k6JsnA8v5cJOa4lSH5TKJ073FIl3WVN1ixjC1yNX31f7H6lnn5
J5PPEH1vALYMTk/w401S2CPo92VBse+HDSbHV0qaVW/rX1wREcgNLhq+ywRa3t3y
PuajYhnpr3E6rI3rXYHttN//UqexR9mlkzy6hgMbxF2cz4Do7FDbHuU9cuR5lUzD
gpELTvNMAEkhPJdqLCaLR0EPvnvhNKGSCbgKI12O8+PqCrJybmwgsA28lGDtTn1p
CdJB9morbzm8f+/Zv7PwuKmKms7Fn0Dj//RpcLOhAg3s8dbeO5mwZM4+n57sK+dH
OxDhfweplNsAe+ZumFom2lMOC0uHNUbBoI73g85HFbGV1KdSfxDFxSuBOUfy4lcU
e9zL8wjS9xlu10+S3ICvDGiBZxT/u9bAQNpEzYLrCukvTtXShm0Dl68JP+g0aoXz
XV01vjoGvwIM8DNj4OlNfJfNSUH0gmkE0nJ9OIPJoNqywqfVx9uaY5iZRm02BQMs
CVgf/Nl0W/uEYkiGOPq/EUVqURmGXMHmnh3vi0QIeuQUe42mJ1wFU097g3+/TvUY
qgK/mV/1cWIhXKqhrAA6oSPsKg+y2fLC++xexm55yJWaBU8E9nZFMwdXopvzkQdm
ALzdprQ4mZMcrpkSpAmlyETMbteRnj6O6oQNKPSyuCcV/FPVN63/LAuk/EtI4TgG
OzjaGp8RrcGjvn4UVksnH7lh9LzYmen03MndD/DwUEgCO0zQ4K3avg6YVspsB0jw
zZy5vTryBUImmHHt0SGUvIWnITyVAdTgw4zMeLrwMknVz/MIfCeWOQ6z+Ed/M7Vf
TBXe/nc+jWAJwJSNuz+8OYKEZOqSVyMB8kv+BOfT/RKyv71IxyyaAV65feOli4Av
Mjx359bi0FYuiiRe0UYF/SIdcdoCGyG1CYdgR6tQQz4OncVTnLdD31+xwUHpNfxN
8UBrhO+D0fpbi1r9vLN6Ou1Ahd3d/V7c2613/AVYk3uldbEwZLLqLVYTtEx0nqkZ
+l2CwMQz/GJzY2DaaakS11ebZ2JNGiJCPRtqUTUHTKgyBFHca/2+ZkExIP1gGBy+
mIEkGaLlY7+oSbNdteD6ICeji6KOP5/G2Ah3j9lGwqoWcRrefP+lfOVpMrvu68Rk
qyLqxr84NrpNYhTAj5j6JwOfjqxwweYMDnTh5YYCWB2c49dhicS/hivkzei/s6L9
Jbz1W0Nh3RpUdDWl5IDhUuF8y67Zn7CiSJejGbSt0Pb4cAXYrhdx1i72hoL3fA4R
dR7hA+LMRqmhusucoIPEC+q3He8bOQ3/7vBOAo6pmfjUJ33RRiN5o9asZ+4+HUP6
Itrjnevb6juGvPphinqvkwfhTbZ+l6rcX6XvWhJVRdK29ZyvviRG+VrCXqRYzrnQ
1MdxoE5S8eMVNZAzELrI+SHnlKbVbLRRU2uIcBYvVd03Hq87mDWa7fgoBbiwMVsU
NISXSenSu0DPpe3JLH71/+IxjCtqtBICG7ltnBxDjOOx6HBUgiQEfyrm7Q+AzKfH
6GUxCvayh6vdUSfU3VWsBLkXtDO5fHQDSwIN0ezL0nMZ+KiXrRs8sN4j/DrsomES
1slCgr1ikn0dkPpA8qhjxFruTsSUHhK2faICX9jgpGOsVB0CB3tk4nrIgh30NLMj
tpPd6DUPp2pxoJp+eOe2V2zfhAyHU+CPmlogVpvyf9PKAHL9sdkerT1tVF6qrU8z
eL3krK/EM2C5/iXNxtgoVjkg9f+Gzk9MXVTr75lCVCDHxC5SusB4K7l7aA3J60y+
3ZYiQpNYVUpGKWqxjFGjsIeK1lYm1A9LNY5wbZZz/pDuMmrrj7Ml2F/YvpE8Yz1D
f1kW8npBNDX5+weliJiaCU9Yo2KeiGW2urDPZ44DQD7ykNI2nrQDwJyZa2nLRYkm
bd15W63Wdy9t5hkfgZ4gYt6LRQVlE/LiewM/LqOwTFJVK5mzf2xu7+kjtP9lSEhq
uvG+W5nKSc9bUtsSD8BZ4iOhZqXfhFvKtA7vpBRzoZp+6sxiheBNpdqsBv3i331w
zNN3kQeVTGVThzL586YonUJInwYSsnYe4bMO2ZPIzJCszos9UAiLpiDv42q24z/R
7KmMK969aX3rF037EncF0U618meobFeUz/eKFY+0jt9PIkX/sPI1TolE7zGFPlOs
KsWcUT73SUnL4D7/t1lPSksKpr38bftr9gsg3gQyKCggSHFe/Qg+e6yfwr782WZT
98+90cM3412KOYTJclBKA5dIc6SmvvqpsYp9BRbKicKKN4mE0ImP5UevfMwZsajQ
FP1IFncDsL7JvsRc7QgKrmWU3+sbpTALCXh6eoQPFM6kNjo4IluLjywgl75AExf7
254Cwl3Dc4lLZhaAsQT5obvlC539shmagHzLrqNfFx5JEeAFzOQcWbxR7L4lfX6n
URWkPB0ozUyTKarHeRUkNgUUWBErxVZ9d8q2XKHxhnllBTmD7g0w90nySGvkeg9w
5jf2lcxwrJI4i1iQxTHfnfRHgmAmVd8DP/TJv96EsPc8y5bu2HKjN5wnQuT2CAqR
JDf4jXtxnR710m/gM33sqxeNh99dXRs1sI+vbr06jCeF2KNVINqalQEeu5crLK6D
8yGPsDbcXgbIicjJIzceK72kD4cTBg31BR3gtH0R6sCk8nbKgZ3BXXcGw+f4VPkU
7MUY9aN04toO/kaBCjzJgpgnpElUIRTxwPeMgeS4GW8mgtkR1S0j99kncSaVd0qW
WZ1C0C7FvNxGFVuBMPBsYNlu3JXfpHQSdES8/GH3eQsNA051hn+gWRYufycoYGBX
b4grn7yZYXjGH7aC694POOf+PJFZUTgOoeS7VNuCUPgxrME2BdLlhfeA+iuCRoUj
PwVT4R09Cq3Q/+I28IOkUggkLd9nxUXwtATztdx2nFcHVOIc9qOy2+C25Jw9y5Wz
XVHDzqlIqZLSi53mx+gTB0I1v6/kyaV2iO+N9RuOqYjihkXPjqipqQ0XW3TerX9x
OLdb9QiXTUsTio7ENIi9nsgE4X5umKIuH1TxzRDjOhvH7mb+4GpfEgAGXOPkGh7P
eIwoxz+NammxCAg+gkhlHc9y3cOV9joSeAGTLlGAfr8l9FhUbBJK33g3rfelRjBZ
hdULU7CzWQ5hJDMbWlX6c3CXXtPW/viBnkKyLEr+4ztGooP4o4qdeKqhGuj3779N
yn5jL6NVK6RiOhsaMDBlxKh2mF6t6FHtDRmznbhZpgntfJrWhsjFNbFj6ICarZIG
xUKeAU5j4brUfHUFmy54DNCWDPYMefLEdVbkniN3tOxlJpBjqBsud4ji7i3Gr0Ej
1LmJDDgDqCh590XYXHvZnO4uhMLN7WnavEkc5GV5FXyzAx+7Syu0DqmtRSLUJf99
Wghx0f5Th6n3qCFdx4mFPnrc8ED0SmEXiA0w3ZDcgT7tPlc/5Uq1nKBAf0YQQLS9
FPpMzRnd2mvpzr950HecOBOA32CrDuJTI+uNhLrOkDHAwGFMV6rLFA7rOnW3WZMR
CRlWUdPrd49S4FzBNOc/PHVQ8AR/ZZtWT1wO719Y+6wPIZ5MFynZ05/W5czDrd0o
/SjGBbEonoI7rbUTSbykk2fo7YfGUtB8rOmyD2rku8O01cmy9+VRoW6B/L4AeaMU
f8HKV8CmvN1R4xIGZJPWEnfJeM7G4JosktsetlJJYGsax39hcHNP7EPo98eF59sy
0SBPQwNqeywEoqZ7iMWCPT9ywKTrNTJ9lOaj20cssvR9RoaEvb+mrtRE2ko+sKNF
zUDyhDi6DFjLKk/K3VUZ1ky0oV6/aCGIBlxqT+fJWLfrUEPrvo9mHkAn7NCURKMK
ntFe2k6EJi4jsFRA6ZA/Dcs8HR1jhZO0ilS0OJMkDO+Dhy86QraqJilpq0yo8XIm
MnEkBMVUatOk2e+wNJGFmukKmgt3LRt2ef5UR9flZ0OcCR5Qwnk3X3tQWxx+94ur
1ER6tFskVxXIOyIfBXmmM+lJzrHrqTf5JTAzGnDsqiUozw+ZErsfgKRxwudVv5A7
iVw/7jzbPjPhdLxJmHzf2M3f6ui4lm4ZL8xRL4SHzEO55jQeElAa5uiJcG7YzWXM
O1CIjBgGnMPK8aE6ecPrqR3hTxATSQIZ5864Ob+7BiDtBTsH5w+slp2KN9FY4H1B
n9HCwJzQ8HaozFVXoFjFgfcQejGl8CRgWMWPR0n/nShR37eS/f5smCtfoNX/i/pP
UnNrc6No6nmbS/7Wprr7KbCErE+a6OxHf4pIDIsBeRgJKf+rgZRt2FGytureKHzh
tn6hrLo5NBECxRGJqdT9COnZXUgBEzSDwvRNrcrm9oGdBua/Wet4FCd4rbEPocQR
xbwNJ3p/Q5yL0wuMabWtKEG4JN0O3COlZ/eNwZLo9/TdY7r21Zpm0+sJ1mgvvr5I
ht7MEiNZdcMelrQolQt+LVzQkWycbxC1D4ep03PfG/an6x8U69zeeVWfoBsQC6Wv
Z4CCKor4Mx2/9G/XCCk+BMwbEextroEw3zsjomkkt/8P06EVBcfOyKv2UEqOkh6B
y9CM+X06OorGy624bu+dPQa7rTG109GWwHOwp21BbkmZ5nIkkKxWVeMUYPag7tvO
xQS3P4pCY2KnVzEeElbRE3uIefObPqxt4TaabfcdYECDUupdwzQ1I2V2ez3kX3zv
BSQEQka0gdqW7evHFlw4jBPayeIYPWu1bK2cum1N8Qo92013RBS2TFAHq6eaD2D+
PSm+g27Paa9TBtw9DJ5QiYjQqYjVgfMCrfDeWDFWRaOLKV+iU/YmxyqH2HUDlKfd
XnUA8QgwIQPnpUHj+btDihwU//IyerowHxEewz+JEXalttXp+p33W1b/M5QE7emQ
LQ2IgV9yvEZ1Ql8N5J/800SEPdE6jKJGTzb7oWCPB9vN80YOHrD76qXMyvu5aybp
iYOxWfI3zwHhs2f48h7Ogu5NV8GavLScUDpJU9EFXDJ4xG/vgf6qE3U1pCPnYwkJ
SwisA2Rdrvrhn1FoOzgrIlULyvYKfQhzjTTuEQsAv8LxwAfHdd1vWWL4G0LnQQRs
JRflFNvLnY4GnAyaDrTB2Ax6DB6XDiz4FQSa9W9xS1m4sZYEUsNgzmRYMe16m1TH
mpwUG2MIqBnMzkynKUG8Qy9b6/aPjRJcyaxW+8xuT2xGJA+9vMwyQ7DuBIaVC4fe
CtnK5SGg2ruvgd3mirpNAh3dueR5BDw3rrO+iYmUAFWtaXeFgtaK0Wz6Pf+P1R2A
tBwq5f+s417bRlIIwZQXwJWNRrxopETK+G5XSS2xSd0itU9QszbHv+t6AQXYylhv
Str37ZxsxLYBy2ehoDkUidc86N/Sff+nqg1+V5iH1HOWA6B6xX9XXlAkDs52n8fd
N2ZGH5XEJA6vwDRagYNz1J9YikCaKBr8rQlkGX3J4bmvm57PnGy3jdyvR40gl5b0
6xrsDRcPgr42lup7O5l+acDXsU1uEQWTbKInnkeH5TuudkOX0oX2/ksVKWfKg9xw
5bKjhRaP7ecigiq4z615wITZOoNhNU8F5DtdQMsdl0CODFPlmVDlpffeplmJkA5B
2WNUR/avOZcIIhqAaJELDDexkNFu/acpIorqtiOSeMpaIqRBQw4tWzxO/tt810w/
VKeCsWQ1RQu5EASLMiGI1ngzt6nbRL+z+UG26ddCoqgAwRVlol/do3JbWlg5PeL0
mzDRgkh8MXEkkyIvydySJj7ORQZh/ROa7vQmDXcvlBVjwa1KvOniQAClbKuGZSYX
n9nImRvqjuxaXyyzFFXV5SWlIYE9SKCqOrreXGrDCsvkxT1TI6iHplrcghUrKweh
1IbLnR6nJRlT564nNEPNRP0WRcuuupn4qONH8gOkLDl5j1O7tJx6alaBE7K+gYPm
Nf+DHJBZ6RtoTGtp5fGrV+ZnZ6VlwkeTCE9iJEZRDrRpxwRdhs9sCVc0czLBJ09m
gQQbyowGHfwjrVmWh2Ng5cje+QQuYSPi6VQiKqrvswxn5XvNh4ADpGaCb55XqEaf
MdjglbKaC+fO2CwelzR4qPQ6GxVc1s5jii0h0fbxHS7wfeo4I4vOLcf932KmAlE0
Byc92rae8FmfUiEZIsy94obu6yQGVg20UV2OKUHtG3UL0ktGYJfatLCSOFPVP43H
8YU1l4YoBpK7r48xihlGKmeTBIgeVRTejTbiRrNpockS94ZdGwwa7OC40eesDqhM
Dlmc3Fmv9svADV8Mjy72HUDi+/YVgl54dXp0mz8ToEcJ7/Vfrp1FkPJt61sEIkVG
Lp6ywsQIAYIoHPFgT/f1NOz1bvKn8MS1ukAgQmAay8jWPLxRzyJAHG0qDUYsd1Gq
6H/Ljak7J/qpGUPDFxCWhBkyT5VD7U2WoMYWJLLHCrSjdkmJ5HjcJ6rc3XFWqi0J
TsUfm4bm/iPeHb0itDe2uHYEKfsPZRnAq5JSYKw+1UCs2sZ0jYAT7lLmHjw2eTpm
g1BF11HxUfVOKyZSjMBplbykT+X3hQP6T10nwvtEW/Cz5P3bI9GvEwpwMnU4AwRT
Zb9Gx4EbKxmlwUyXApPofEoyV78z6LpOQ2MPT/CTy1ztOYXlow6XW/uRXhaW+zXo
abJRrc/uaMPaWq4cF3rzT58Uzg1FQZFODyZCbz6njnYWnttrD9jKlkMoiXlYyKl2
9IFJlqFhtf8siUbA7XJBv4MWAmKtI7Y+QKY44pY3IjXK3ACJpCdwpY5DUToPyLMK
5Qcfs4nyCzhXfGCuwpE0wMXWDNnGj5CNiLXfQlD34ZKHhHxAJXz4XJj3aLKgNopL
OqSMK9DQ31vWl7Bk4Rfb44lfwKOutd6COeC37mKFd7iIhLsnvfm0n2CguRtuK8h6
r0Z6sHQOJ8OlwcxVjQtkU70QxB2Bi9J5RExkxK+HB/OIlOcKf/UEdAo+n5xlnxS2
tKt8oXV9mAqKNw6Of6+Voo03R+FcsXc9znCV8eo4bSjpZtRjBIZhhUsMm8ZNQyjk
b1dD0vtmkiaizfVU8qc6Ew0WDv4r/bO8afLIcTSyRZrF1m4OP8+/U/lICpotKOJi
SHmSgtPXLggtnNtZyK6mWn7bnEWsGjONiMP4/1OjP5qagrbvggwdyKy6WvSpXhMV
wKugtoYJDLr5KKOmjA0i+tyaQafwfOi5Z8QnZ3DXIZsdYxeaSKgUz0I40vwh17VW
yfwi5g2TFY2cav/L44Bx6gLnWfOttEvBpPhhwdc9LV0YFGS4AWMkm9jxLCqTCFrf
K0aFeQ9F0fORFnd0dZDrH9/o0joDimBkbozQrLvv4H79trZlbT26iPw988xclhdq
+OtXg/Wg1BB22g7LDgCW+W3vnqW7yGanEXw1CrSCz/ros5vv+aBW5yfMYFe2Cju0
WdZwGdTcf/LMKaVlDTpWepb8BuMg/+CK39dh3GHGFg+OCRysT25npw71yWCNMP/Q
iw3aK+ZZL6seiiPCucp+9wI3X2duKYaEBpBDgYeGbMF/YqsewA6XpEhv7gPach7t
wkTA1tpHddEaJlQvNMz3wrCCBW3122Ok1Gd+HqhQ9SCBTVrNiIO2a5V8NnETqQXs
wxGNNYzDeRVc/O7N+wWj/InVHb5OHLIqhyfSQrFLONcYOaeEqHXsHWBd+NsLloEd
L1Z9p+VV2o1FM+t7yVQZk1p4X3TGpSfJoyCL8Pre/tuuA+6hISghB1zPiHNPiiQz
lVICUR1Il62TG/HfiyoNOL75Hv+VvDRnEO9nEM+m37i6KlbzV2HbJI1eZ7uIYtGK
3IjkeyX9Yd16Hzs/Ght+mogzuxO0kDKN4A99cyouFEW7QxGYp66wUtqBxLhx51Kd
+Sm+TKpiXHRGwpTWyijepNvK8eMCUov4WtM2aaI5m69rII/g8cJvGTcsbxXrcSbS
sGK++p6ejbNNyo0pkZdoTMzLYwAm3mervZ+6aApra/ZRUA2Vcbe0I76uNK9lWhdb
yKGWiMMOCXXxW7KaM98Tnmz7vsn6nsyrmBePQg3TaPuO4J2jfF/DyVn0ev9pyr/K
UdXVasBIJsD3fW1YWmrKEdCMAMUF5N8y1BBlJeGqiP/6KJ1tL3n6ccBmc5Hnb9Tl
InGIB8scRb7l6HqusvQoOp8ZRx7tW21CaGeq5vo+J2StvC8qkfjYkEhbj3GkqQqm
/XhjdYWDSoG6EYOgnQ9WeH4W9xVB9Y3ezTc5QDcEQdVJilIf0AXqKk9mwwHO9uYD
ofAQ1cU6LmcXeMcOH1Snn6ZisYNKvd7O5BkC9/YYYkBeZXf40vvGvghwPEeAwOPP
9EXH24BYjHwSf3Y/C8G9KL6kCX5YFSvIw0xOsVI/yt4gFXEaj0HO6NUK9WpcUT/r
j1lCUNR8bhVmEwpYWbnFvAok44/7PXahzrJgu4TA1zNLhxozbkQI93BTaeySiEyc
VNYuQnNuGlBPmJOLPveQcl2wFqnVgxcUeTb5lN5au4+Gcfu2s1YZkXn/ofrXBGxJ
lNATKhWOF6/gOfr/bX9KerNKFEm9AT9Kz0aKMmBBg6GJxAQ1KcuY1Hs8ZaFFGTCm
XWU9JN4rP71nuZXnDiGjO0R/3sk1gXSh4vqBY3sSYLWddD3M4EXCJkqNHrl24ZEC
Yv2bpIzFTOizJ/pV4I6ARil9Zm1qgRqou2rSI1a/EoHSYttz3NNEnPOfwHcn5RNx
H3p5L0IQux2J3obJNGdIFdrorj7HQjJNXANZMyW38QXlLaa6hOVkI73jfdrEJ0zZ
q4ku2KcWymz5m2kANl1JXk6VEuy5l//GySDtXqCo6r9Nvr6Z42vkDHGoT/WGzqHs
q+zG3WzUFPEtP0LXLP9SE5yi+0L99S7+Lwzln5EAsYm4qadi6J7HhLfWZHFZVjde
eU7ZuDHG/6c5qUZrPG4c3H+yfEazlcTfKfa6IHm/xFxrRqkqv3TqCRenOeKcRmUk
gGZqIUnnUvvBdFkEO1KkxzZrsT5u4U9aqaQogCYnrQU2UBjr/eA2LdvJZBbkN+Se
xJM3p9QetXlVf56xK/2amflyhKMiCQi5XW4gpWg4imgA0FW7bXrkxY0si6/QOVM/
si1OLgtOHaXINyR6UcH3L1pMqXNcsA3RvFQk1ijk/zw8bF5kDzTVEbPj0d9f1irW
wm4Fbm462Gv+qz1EXW0J7C85vHHLSADdljDcsX2yo3uU6h9Dbiw41onTuNtpA1mI
6d+rmE0JTmTHwtpSiV1uYndlBB4hNscdCMASUYp2+NogmCPheIYtay+5eDmQzSgR
/RdJqVh+E5cQWCQF0UtQwab5MJsRYupGXsypgf67rucvni08W7i1X4qENC/mYqt/
A6DrbX4GiAi0gs3PykpSip5OPQ0aX2DCEEBxZSA5Qq/2lbIMGF4Ugn6mNatGDqMM
9J4M8eBaADA+khGyUFTt2cZMCyWe+8SVMnnBUJojFbWQyk8Esv2LNhrNkVwTnNZD
kHTHcNTsSBliTt9ouPi1PoUYKvVsM7uuQbnv6hfSX6tDAXf4zRLeirL+Df6qPnGp
V3mYOsBHY+W/HQUEhEaGlRI75+9bZ9MYCC3XirXcmm51oIBLYqvFDxzZc8X671Fx
mpfmR8iiAcYVBMNgpePxiC91FaLp/dK6RBQbNeGV0f+FTH/iySvfuPAgikG0BFbw
EOL35gicYpuXl3R9Lu94kJQjhzH/bf9jnXRKkW/0WUJEywJQtyrirWAkbeg/jZ9k
zgb3x70H7zFLy5I+e3OfHYGsvOFwKYjWf5IJ6HPTYaF9IgUVz/GtSwt/Q2l3uDhI
WHUeq/epuvsA/rHP1CwPOF9tj2CG759VLBUcjo0UHBZcTuFQSJVVt2s8PbmFx2GW
XxOJ8d21n1Jgl3tgTVBTRiMm8FlTqKRtQA6l5vYAfryONFjTILZS54wBNTKmC+K+
ShXOnU9ho0x+JtHPUpIQPlNHB/gcwPPpJZIY3KX9BORlYSFYiIw1QRuSPqGqUFl9
BYuDNwkv2ZO9XlQOuRNgBQq897KOxsgDrh8H9VmXPdXJwks5hNgK1B8Pa2rQL9+W
nde49lupiwqELRnnJqfxTFoqlxuF5GyKAEfMHBhxNWnxWFLVR4JmemIwMmpN5s8t
6sXd20KwJDn44tC5cVmbCuSzOjJO4G7hu4oClfkugRwW0wsxe7axC1rN9fwS+IyO
RYXBX6HhDR87WCSL+ymTtjoS/3weT2DQmRJDdpJ4Pm1OZnfJvSywuN5BYTIeVyS6
Qj8WrjiN+hgflGGXU8xRheJS9CY+WJmY5BfUWTkOTjzeHplPro1nAmWLqoA0rXxs
nQblb1L3c9+0DF5GkIFOj/JTsDn9C+VuM8dLlXKjGB3TJCwTxZ8MPli5gRv6n1Bg
kIM0P6z6pQfDLylf5kog/Gwx/aPNw/o+452sFqS2vGDb13OlmKGrNQZrIcHeY3xy
ofSmtpJtcLQ8bMKc2KeJs4XZpdpVx2sha9YBqizw5z/3a24wE0NAL0r8+10bItEK
UeLcnhaLc29MwdnP579QDfjMXsjsZ3mo7bw8WugE2+XI4xDu585zLZm6d+XJTTNu
xkp9EZX1SCz4By0OFtRK9Sq++uCFZ1AryTFofm84JS6JfHu3fKuknfsFJPbu011U
LyczL/HWPnLc0tJ4ed31QaTGPphyhjf6IkIPw4ZhhPgDeHCrg2shTIj94uf7pliZ
BPno0mZeRQPBH2883xyjgdcSU+ZfM2BtmwrPddX8gSMPVJolm8rF53ykyMDloYjW
KIAMwLciGL76DqoNTeBfEbty+Ma5pmZVSZpzyI5FNDwBlw5E2m/Evv7ohqJbfGCN
2G30SBAr6m3DvgrPGHnsmhhwg284PxiilqUd7eNv8P0gsah6FxmgkJq8Vfl3DC0F
XNH4mVG2AydAw89+DYQvKkalzoIVSBodla9QCGQyHdFqCOxtI2T5CLePAQyNNFUI
W9fxgEenzcLZtxces9YaeNtrst2MExue6/84TxlJzcMTkNGhh5S5cdX7WUvbp3jd
J0zQVuoZOXRGmGCi9SiZQf0snmIHyCbpNgka3HAOfwu1K2yKzPyWmow3Az0EStTW
5BnTZtFODvADXmgEFTqW1zuaObC5PxVKYtvGcegTTfqSJclKU6vwQ4uQYScvgvAE
xunRr6TZKwIoonFJ8LI+3rW5XXFAuoLayCowXQdkQGN/rbi1bEkwHQybzSHKXJzl
IleckVOdGc6MPZi0ycNwpu54ucY5JCQKIY6Gs53qQyuPF39WctzNCN0pZlcIIBtx
qliZ9b2XRXPPvBxxMjHSucI0eH6VI23qJr2yU5H2/vnMyimcG/suvCwDXjpSw2x3
eX6RMXRL6tWpeS0tjADoq9ViTyzOQWmzrligMjcwkl5DC60VgUy2UnPQokN2uiNY
dYUn+rGutCCqUUEw/0h7S7nmH3ynfoIgZGwW98m/58KexHlV1m6np6xKbmxQ2uTg
T/jwMr/memqZlwQ/EBx1bShjiTGF24JF49XCXxe7EliZ+/JXjAqym36WsAZT8TlG
JA4R4GqY4gblk0hmA5rR9ciiRTiVQS7UgIXKykfBgxvebJlcK1dUm1b4kIrHG0cY
f3gAsNKOu5mtPkK3beQaovVzL0lEs0uIKgOPhdqrTUC+UQnAhOWviWB42EOCZwJ1
FRx7XOZzoLj/g61YcBOIDLoHyBoPu/tEhAlC5+t2tRyvmEfNFxlOR+aZKVOWpfEt
bCDuc6stWZKj7VDSjjnDieLvhrje3RzTFvAnPG+uvqMGIv5KFoRe35KEZgM6LZvf
G5+rNemYAxM3C7+tAxGTcXqD4v1tQQUaOci92QVnsBtWURB8WQg/D88ZqLLZJuq1
Fs/eQESKftGfCTaIjd3NkbIWo/iJrGcOITl3FAXPeZvQotfRiwKpTzhpsYJtcSSa
tadM2zoA2rAbIMJyvZvR+cY3Bhd8Pz8psFTXDNMTfkZUiffK4qPpD8BExr6njR2j
ppLCnMaVzM/qdRvyQeVRAKB5cWRso9B6NCMvKK0++vE+qhLMIOkxe6RXUXUhVk16
O2lFMY3TGKoUTB+CK+MIoukOqlyv1Crc0KAoYzyBHNC9cZM6c/3Lu0TxhSIVpsMz
4JMZcU26n4bbTFGeQtrNKCEI9nm017Ih6Qz+yynCcq6BXRsD8I7yL0Bve2dZes9t
4sk8MFITPZsCc13J50+yQTMwZJZC+jcEBDpGT5LYD2dImNdWsuvP+B7xTxPRHQI0
XssmxR4vcPL7QDYEyLI1yH9NgMtj0yhzpmjgzAt/JQfpIRSeWHhMm6XH2YOeAeqN
cnrf7kQXODBGnXt0mw4OcaxpS4683VeUmKx1SkO8+heviBi1Ced+rbPc7X8ILQFN
kOYbkgcF8Xivfu2eN4/WTRFk0aianwXPKQGu8fhePQORFzoTDP71YN5+NctFyGVn
QATH4j5+1dwRI7iXKolZGxzrqxYZAJx7xIc/fbcWVnFvT9Dz+79EmeCzF6rZI8X2
crmh4rVy5Q2tS8RwkBXrdTOnDnr7nGqC7SWN2nO3bwuxcV7sHHh0Zr6Ln4DhQFUv
SArkSnMzp3+t/L3VtTl5KcWkJtN95sR8ej1/pwpNG34UizO0dWx2jjc44ElcNhJb
MHoQq+q5MsFNizU7TtBVdFDyn7vg2ZOzKJ1nUWq/0AGFoJfLxvaOXoCrac12uNRr
m63m+q8d/5P/g42tYv2XzQvRbRyYx9VvK1ePGN36zeMRLpcpgEJZeiGFuIahIPw4
EJSVVpKVNbCBKojXEMhrMAht8gUMOl50HfFDS9EsRygvJc4Xjhj2aWyVQ3FfPrjm
nLZDowJwGYERePQ2TGQ5+I/lnKocKT1ZhtxOx7QcdaULs9C4Nlu+5fQo8maf5YIE
ZClMBvP/oiqxzGVpP8w2XOWpb04cseQc6wwdFhW1f0dSkgVTCd3OhgyNmkdBIzli
kj8owG4m0IyUnLPPUK1oN6OLK1gLRvX3TzHQ5WUqyZHJKnY3FYqd39Qbc7T2030u
JlqZ0Oh26FmxHa1WpeGg1/cioQIIqUwkXpmTFVLzUeJrE5llLI1R99Z3Zw83GIqm
11oN3wB9iybsKpmE5nfO7LC9Yl3mPPjt3jwPV+MW4ls6kyZTXon7BZ92nw6aKnEY
5CTWVmYWve2vRisus0QXhBuRSv3Bdzbry4hXe9+8FtAHAJ9dVYOPymRVIMDh+bzC
jWD7qy767iMOenn+sNHPR7+IZPfYNX/kU5STgnpFbTO5FeR7L/e1xeWS7leJBTBQ
oBVbzHG7B1iLwbouJzgOhmgHGqDGKleozlhk6aAyfl6OggAzAHDGywBpIh87gUrj
LZoszwR/oOn5rkD1HqBQF3F1gm7kvJeOM5Td4Wn9e+ucSeanuhZcyPCgUi3iJ0lz
fCvCsfbd0qY3Sfz96KumOv9Hco0v96RdW4ihJmZ3QGyHL8awNuxkqbUcC/1GZfbn
thfRIsDJ+Rolnqvs+mNpvH72I3IclHrPk+FJowUmYW1qhIRsRPmysWlRMtkiuCwG
W/rIpw6pndRuapaFEG59zn0kDFh/5yMIezo/VFsGlzJCeHediKUjAJUeA0ebhMDi
erY6lWKkMGzR2k8w2v2QM3rvdBXpd+G3r6c+5AYJX/NaTl7ZSeg/aCkuSU0Qdk9o
bb7CHKdV6egTaD5BvDCkT3B7Ez2KZ5C9gixt1mI0qvMkUJAUKpEBWhsKdQbKj04H
hicAuVoT7OoylniNk+NT69Eys0LgrXFWqAys6dxmTKZyffHqQ7ftTMTRZmWqDNuE
esyyPW/PfI3074Ea9FXPadEY6BsELiRmuVaG98+riQxwiD4kZrkh1sl6cmIRkkjc
TJuuUFQtaIrNPafvqw0T28X3D9Z+qgleyTp6TjBPXswaVwBBuCiApbn3eFZ2tWIF
ypDBcLp1D9QTC+PDTpdmE0ppCxHI3Tf28oztV0uziAf1Gw14oqqcKFgQzf3dRASa
C4DYomZUqNDaDWdtuez0KBPsmv/KZ/X0lQ7PJECGZ2TMcztKjw8p2L1raWRQrzEW
ZYNxIrrPRxA5WhlzH/wpEoEr/P9OjB6GejM3Zxo3B/dUyN3tK5SKptgTRUyfz6SA
+yvYTrtxHKFnpTAJ1iJVzvAIFp8F4hrPHK0xGokt+eqRSfbFkbgVwrxnFvxGjrOE
ssSrSWJ0VZAw0rGyIqCIwDpB9eUBOg0RrDrmJj1To8+NEeWQ1BzmksOsawWN6N+Y
JUFP61mg7JrTVIsUPOw1CQJOeUnNHmMvQ1drJHR9yIO28y3l/OpCO2A8D/RI/nR7
EoqkQt1y8nG0VvuHxlLaPacEP2eKScaWwEmhlSFW7X7uTfDBwl/nTZ8aHJu5sShC
5ACLryp+UWsgrA3x8nBahpkY5q45HNay4b1yCY3Fxk5L5Zc/nI6ygAUv+w5c6vQm
Y/6LV4RXNTPjXu5XiV2x2uEcGpww9JVqZHPTV3xcA1n5C/qITwg/BVrEMgw6H+0D
lHm5AkyYm3Jjrxa1el+uRZwF3JMa1s0RPUzFfv9OABLc4dMtNU1B0Mzu/+0w5H3s
2z10FCJ48De/5Et3YpK38V08hBZqdB//3gewKCTFzD9zkB+PpOVayEra7geTDEa7
yRtJ2FRLhimH6tLVpvGzmb3uiIREXxGwV3gz00xIobtPIGGtwGXPXxkJywpjz0YX
uMaQW2/ZI4GsFmbjxPxGPTwc5lUpAUGXi0td4pvUPwtnKcUuJ0z40wjOz0xkBF8U
eingpPXWe1O+zfPfiUHT2Zi3iuO2YUSfS+NL4ZMrFNk3dLKJy/lkskcDU7/9zVEN
gDgG2glHWPEVGKRovd1XWfikq7gw96TvJspt9hI47RHo0EDeK9lXBqWzUO7Krfc2
Bh0wvUKS2mktaQrMnvLG5ktV3RNfwA5Bxkpn3IcyYsoixC/kwLtCQsPjBvSn9b3U
v+jb8p1DquG5k4cgnICDMP70jZMJB8Wqgwqq26jyaB5wOKNHJ+xAn0SAjt13zvn4
HAE/54L5wC81eWxwG1/H7a5PNwsmmk7fFMJuw2r1XDMX54f9egzh84WTKIGg1DFx
vwg5i2kV2PogUFHlhSaNH+ByszC7fyXrKdyYAGno9AWrehkhUAiNAxuNIoQJNjZk
00iSIeraWzLlYbBtWbT/EUHp4fgbli5MUmglNDS/umulWySpDNUWqnW3CfAqWv+n
9blgn59LlEan20ZxBqxSHsLXXLRHAfSMDLXIn2u5AIYoTNiwl8FbkaIAtZVa9y7W
LnTZvok0qyb3xRG7Hw2R6Zq3drL+4PW/L4qLbnepZC2rJPkYC+j9kBfQF8BqmBnL
xEMfgGS7RbV8aEBNXHEoxetm3cMe4m7LuoUrNY8PSczbCh/GxT0AYucZyyb3rB5Q
YWHpTHuMwsLV+k92uqFCGiQQkOubhvKDbPPiravoqkk76YFt9i2Jv+6/+7AnPToI
LI6w4kyf36sqK8L4qd6aKuWsGm83F4rCTmWN7oCjvLaxWGvdYD5rrsmbmtIrSK7J
IIGJE+aBdQZIitobdRAtKIYq0LBIQJ24KV6D4tjnC6c3RuvDFYZ9VFjuloUKZwcs
MlEH38Z0kTFVBqRBAKgv02+VrEal6bGY26AhBcEPLPqDvnUHHL4lZwPSixvf3L+F
quEf/G5lavcPkRjdmxF0SXmAfW3NdVrcMkaty1Xv/MBuwwDsIOqdIZtbFZ5ewGv9
gCw9lL5iBK4os1SO7ZTi9kYlkzZt5Krwms1d0xhsEniDBZoFXPtZcJmbdwg2U/O3
Ss4wNrTxRv7gCDTNkkQbFtP6pugMLBIOrjfCzrHquE/gGp4qIcelq/P8P4/DwCGK
YQnxQIewwVkxJdWvuSSmtjoTPGfORqYIlf2+dlbHdapkxGuGhmdwCjgIkKIMv0ZZ
bNnAFD/gtq+lx7/vdPUsdeRL2vditGUnS3r06mBetqwxm5/PoLkO3Tw6wv8Bi9N7
IbJ99S4VjtA7UnnLbJo1ykz0EKrwozk6yJZpE0s/9L41/+RJnWpQeni7u2yna+Ce
0W3QhnN66w/XPcxGjTcG+Thjs5jUWXKyB7KPpmhIBeqyJeNxvstAilg6Ha+EPp25
xcyoq2ahdtKHNpGuA6AGCik6tYu/tFe+Ocs3m3R42zfaq6Y27MRwfczBwSfCWhBr
WHSYl9HYX3QhoVAnzb4Xe/CRJ0PMzv/OiSylBa0U7F54KcpWtZEBa/ppLufQUJ/Q
/EsNadMZ48uitz4/pQNWfyzCtVL1czfzM/sXK4SWc61CPS+04zOgeS1YaK/v6Pr8
NH9scZt+n6Ob4w/xNV2sK9WMGzBoPdCMVH9Wz369n2o3c3p8G5Hmw4nJhHigkFqR
/tWFv7ZMFWt16lb2TfYNdlFjjOJH0u1YAMP8EpcWIb3h3InTfECV00rxoMKAK+rI
YazY76k4wxNerht6YmXlGSBZ6auvcGK6rV1TcwUxph8AEqsn+exovwfpfwxDiwrg
obTEI27P1ir2nNFUqhu/FoZzFrFta3iMqoSpdrLNV5uFd0EPzNMiPPNvad6JnZgx
Ze1N4lGlkNafU7u5E3xdcZGjc7+BMGBxLaNmzJY8NMUhwHCaLDGQm8G2hnJ4w+8p
rLtyleozrOQsD31HtRJCrG5OjqqaMc1uSzAd6kBV5MdDkJLQ+rvGTukeLijT1SPg
iUu9RbxoH72HW+H86cs+tmkHGoUuLIcMLelLJoJkCaPkNsrd+7vi793OqsW1vNSh
UVpHiqDBqS5NYof14XhHHV/RpKgFa8RoYkTfkihal/sa9g9x1+eFelifwm6u7A48
zxCjdclQgp/L6c33CJbwy4I/fCuENVG2pCkz3/ASh/yvX8abw9MGGmXx7Xlw8Rqo
ElDBBmDI8TA2zb0BBo0F0Zl2aQwAdgEdwpQcRnop6uTCzsSibCiupYN57ABTQ9ay
m8wDPMoOhaI5j49QUD/gw7oZbVYCm6Yxbs0afeo+GAs5Ojg7KPMFVGeLu2aT0MgD
YzcVj7B+DU46h7NCPrBvkZn4WkA1ArHhS5P4eFEJxsM9KFALpHAIGbsycqn/R16p
I+lu8rrwdyp+VoOf8PSgpeBtEjF3LGLPum/SM/BmgqBFOpELL8robtrbB9A0lDLS
r/WC5DewkD4xt6TThghGXodpjxbPHaEEFtBuvAfre3n8PIpfCr7m6OK6QXr4ZALd
wT+PLA16jj6j9g7EmZWNOoSmtcALIonEccapkEylBxma06oRU2IuxX6vBzAg1DAJ
EToYiFYd/BDphxLdOdi3Vkm1Be1uOsVOTOcTwQoDps17dYiYUTh9jqCMh9Sjv7f0
XnHn5nMgB4Df7vUQmmhFaXdOHgeodrW/g0K+mLwXVngibsD0H+X0BEYEAH/9yn/4
uxNlBdijze8k4JZ8p6liyuKYZJozVC1Ei+NqnD6eBM6wmzAbRV48I+N+o3yzW789
V6/QDZogpf7lKzq3ZjkgzM8kuHn4lkHiMwQKU2icX1r4meRKeP2D7YtBoQ6VH1N/
yjBXdyRkQBSKghPWqBmyNs5yozjob3rYF5ik+rN0gbz9seF3RQBVnQjkpczkZUvH
E5X42f2nG3Bjd2tq9pK1W27PiLTeoipGNs14uK0fh9zQ2z3swC64jI5cpUag82ny
33bo2JGTR9kqgkXnk9R/iqGT+gmGbdsEL2toESA1/8/8P1TrCHp9rSPpYNvy4trz
ssov3LRpq3FNFqwyxYQBRwAClk2DfUm5GOweIQs4cX8OSuUQGSChSvdx8hCnBdtQ
phhPcpbF17Z1aup0T6wCjmWVy/nyqDBM+kG7ojOONY8i52GNo/fKRmkrailS7c9J
gBr1QBJCzNMLbrX7ARSO0DZEvGcKfysRxuu49OemdpRosVgfa4ap3fc5vE9aNa2G
0/PXO/lAqrndoMc2b0rQAXI5nhoGHq9L8J1V5azpmPB1cdkjQ9ZPdoEC5prPSAV0
VVX60zw5rxYSIFLwjJ4eyXwnvKVG9fetMlXAK7NU/2QjYVZhWbaNCaYK8/MlZaV/
EQf4GSjPtMUbzQ9+6ohuBOiSMYNGQfi26IfYpVsjQgNcpEv/vXD0EIShw9zDLqb4
9TO2XaNopqqORi66PxpGheP+klV8aNzfuPZU/CcByGJnrNgYJ5+c1KNB9Xt8HkrQ
MBVR0MG1K+qYXUd7Xz/mVwxR1/0nJxqAF3a0P4e2C6eCS0tLTUWPJ5nkddNod+a3
+hOppOiOJ6v/jtr5V9EPGXDft3IbItzOX3JbpO56J5BlUOTV3ExDUrIHCxHMPUAk
H+7lDdAEab5K1kWNxWWhtd+l9a/4t4CBcni5F8ItyaI7idhVUMZmqS2fEaPwMCeS
m6GWZEXZKkSej8J6uhymzIUoc5auba9t8kGuTmte5fyNtdCUrLZt+DWItjjkSrTV
/rjsRgf+6rGEWGuTcsROKBtnB58Db9sdN4Oy7CdCeALXMayy5aNKycTiYEThI7X7
JeBczwPARYxjYBPhpSVYWo2lcdhBIKFxuBhpngcIzVQsaY3OzcLmhczrHZxTqX0g
c2p1uTsP2ie1op9NCAlNetRMBwKuqXyIr8pJhPpPQdp7n2hQRgqzexNt5Gyw62XL
/yJUHdjUNjR292GA2rX6LFvuPbmfAWwBBrz6IOW/JBF28vX0DPJae0xpJtigEtot
Hv6xRT/G9/CSJj3avrGMzO2UprwrhLs2mQ4MNIQgtTLeccEKNewS5STeaQCLMiqU
FX9b6RmPAgwycHarIx2yq7wIch46UGAdNwCGWNNLQMOwiMSjAq6TBHDl6AsSkRW1
vgDpqoqLfXKY1cJ9W9SDnGie7vaaLRDA1JHTa5tp8RXw7hilN7Kc/asGlcWnVgX5
ptSntAdu2jvJ/3+9/ViKnsnfnRovd+msKX5AgLdJFZfCQFhXFhkgt5aXgFjcsTuy
a/dasdVeqhjPQsa4Jq5PrdE590Q3d+zEM9i6wZqpHVb4R1Hc3NBrVriAY46eNYTK
OoF/x5ShOVDP22msxLHOXckHnZnmhrsHVBHfWWwJO05ouFG8sLeSD1xy6LVdQ0/j
dHL1B36bMtUvSiFYYjqoeqCrS1hbvfGgA+ixjRsEyKqbKOLo1qTzyfTpwoxXlK12
aSWIS7/KFrIbQVjtQRMUNRelhOIOJy8d48Q3eKJy4aiwSvRUGnS7dqCZxa/ziG7o
AHpOCY+B29/L2ZnGxn563PuVwEBsRHwVa0UrQ06L7DnQtaRKbbD2LUxtWgNLvlTe
wk55rF6dyymakMzzBankqteWHDRYhRz01eSLCf6j+3KafbUk8F217Ga3NC5D+Ty9
zrE342Zg2sA+GtGk8Sfxrt2sW03ygyjWnHpIcrLe/9w1hn0wpy7i2Zj5AAX0izrc
t7qnIFUfnZZ1vv320sUvlt76RCFfmf+k4WSg89B39rtsjU3sD3p88ZbHEZiVkVVD
aM+Xw7hIgrOKl4M7b2FUCs4QSqgx7wo43u7YspGJMW08FFCZWH3W/iN4BVj8NkSS
rnrNKDn8wkOI9MIXrszcETerDkxNILnq0yeOj6DVua3vwksAKz6z0QPjCpd4/B5f
kGZFJwvWXJlwr/FuJDDIhSK555AS2JQ4JPkUHVDPk3yaYkUQrgVmDv701NAOU9DE
eTn0LDmxkuLoYCIp04qkTVf6IBLRw68P3vis1ptxwRIR8CgMAcudCT46yqL8i1Af
iWp6lmudo+hrvxtdpCRxlpGNT1RFnLKu3Z3wz0mMp02mPGB6a1myFKFLslbl4s9X
JTuBexPv+GlA4Us2fGLPG4er44Aqew95U0x9H0l6zRbXhUsWZ6ZmQJmiHf7ua1TM
iTfCxrqs5A+c+na5dYY3LjT+tgcdy0ueB+6kYw1QSjIQXxyU2RDfKg4zQPIQgSx5
nMEgOXqlCETj3yvz8AhgVd7Dy/r5nG8m/miTQZgjgXe4xlvokK3vmLE4RVGLgm9z
02bJG8dy7raYuO9lrdbZSIbtx8JmYGt4qXeWgMd4XA18j6UosxaqUst9e4GcHHYM
S41/14M1pnz9bE7tc/IX2dX+Fl348RSTapGqwO6DmXAR2Qt5P0owDfgkXbGdhM2K
RUgw3ntLrxNYq6ecZIJXrGEygxRpIm68ZxQWmQ5m8TYHkskpxBrkFfgHw+tTwPqJ
DtQYDM7bJnbjNjUwCstvxKaSOZ0gZ2b/OZLVWLuWohZcP3jouIJwszCAZ+0cvi1Z
8mhWnemixpcn0Tvsz99dN5XOYwXrqyzkpMRP7kkTUmVRSKmtsBY650gCDD8IvKRG
PgwjQ9WAbdGb3RlFOIAsD9HdGVnzPMTPaKa811onFWv50NfzBGL790qXz2nrvDHi
k4FLrDK1jBVF/+It0eh3GNxdzOwskBj9LfxXv19BlZyqhHW4beR+aGhPmbncG9z8
JRzRPi0kWjgI5EkE9A7Zi0YXqgTdOLz+AxYGe7Q2T7rG1pkZk670ikxmXS2CMFBv
cZgTZ0/nhI5xJTnMbjA2EBGecEYTRNHunLxvGqoO7/Q4SkD36Tn3mz/tc3V0zKQY
adwj5/TMzncoo1Yk/9MZ/ZeEHldkSf6WZA+64/13eeamqjT59JewMRTKgZeJaBoL
6hBFGaePW7UPbiH6uLHd8QspFmahbhJUX1OVuDWe1TcEQoyhr8vBznJTDh6WtedW
aslC+vrtbYvgj+7w1ip6z+2VFFLwRY1n9NrdZz4Vgb2+N6zLtjT4UW8xbkE8Xmsm
J3Li9LSqMmkP0wYSZr7oC3xLlZdSUH6QtO0kRoP0YXceG7lpugTeKz77Wd2K0OqK
lEkL2gYm3MHGIpAGEKslU6lZl/EY9t1+q+tWAt1FAP6dZwtXUzAtH+KMXZevQyuE
Iv9fnNTUakRk/1x7bekYRQIyjkTggZkRrfzM2OyIenzkyusTYLwWakiJoGGnsSuT
NpaQ+SJhSS8Q9WzKRaBzCkiknhYYIbkS2Z73KqLT3fig1LdTPRughCLOKAN2n/xQ
kzIRY4bL7pMEpkgdoimYdHEES4ql4N5HO01yNeYLuOuaxkKsB4HlGyEIdz0fEIwt
3R7kIIpliFPwbLLl9C1ZIu2vwEbJl6T/2O7OIKNTztUoLYh0G8wkpTXaz+yYA7BC
wpWemPfEuSSywFodtE2jNyNbNyQcf5ztWEs8RP1jnYZkPrCP2kTWy0iQb1agH0Ya
XpLlI5DS6x0dmXgnPVJIbvEVFlp4x7svyP3KohbF4rpupwbbluQanPbiAH02bk8s
SkbqjlvayQGaBYeITPPlZ7vKPBaWNZKS3t9g+2i1Go/B8dD0EjUcfYAt81J8nfli
b9E/QZwpNKOQn/VxTQmsuNWyNZLLkh3NEi9e7c0iZ/6tP5swWOtGoG7pQGzNkgvR
FLtOzZmaNhiArza1zeDpMUAGwrKFVG1pof0S8B6iInFA6cwkT1Xj7csGHHijxGmt
YWdvUWFRSK7uKaejEc9ATCwWeM4orF/Tp4NtpUjfLH+cjRebwxqcZ2/6fFAieDTJ
Bpuyd54twUd0DO4DUdqWVXjAvP+kSltm4OkwRcR2k0joXat9AzYhd1CtPLMTh55W
cJkTigpWY0UrTIVd+mH4S+C1FoBVT/fSyZFg4kKchNgyf8QJndQgvE3Uc6XsA2mQ
hPpmzHc7A5LyFmIL3W3u8/eY3Zwcjc2gOad8BhRnigvXJcSbOL3/oRSrh82DXKk7
Me1zNK8LUau4WRK5Cv+QGhi/bGFY/n1pldX4UxynynINT6wUxQd9ORJwL4o6t+1w
1PL2au7sgFFcg6GKYlHYm4qU4JusVK9c5R+7WfGWvwzHgUhnBptbypj5h5sZGyII
d7gBNU5Ed+ZqB+ysg9lED0+N6I25iwgG58SYM/CPsxT70tx2o5wWEINZz5a4Bei8
5bMfem3+5UuCPCjlwLds799Q0NuQ4OO2EUuPTI96Eu93oWreoEdM0nrWF+45I7o8
crNEqqT8hBiaLVhIKdUQYEzjQmn1BOvxDWPl2JGq/Z7K5FRpaYU/oW4r8HwAinHX
pWarrwYIm85bYB/yIhBEHKQAbuQFZ5eX5OmdWn6l64Yl99hG1X2uCZu37qGgfJWi
el9qpL81h8LaGlZI5QrhvjP6lZxqB2ItssflDtojfWF9UwWatOSG+bEL92ICI+mU
2j2iklf8Xb6yYWjiRJyfVmMo8kggNH5aRQqcZdqNWx1urxRnZBma0eAmGrzMoPeL
wz7LmYdJRAkhH11zyA/oA975eDXoaVDl+y3DaoCM1QEaNQ/ywVcRaUQVHhAuZ94z
5htdhy7bHk7g+6u7SaUPwhM19EwkJJoch2d4g2IR7ZmCRo5zW0bteDSOYlUs86yN
BGS0rXDMh2mLNlfUJDErhfgo5xh5d2mhXzoXVs2kTfwa7kD9tjMiZXNzVKXkple7
BwKDQ5hrsQaHAbQew9KpX8cHO+2wqKFWatFsh9SN5+Q0XdDHPfH4Rxno7gdFaiqw
JTzQIpo52OyY7dFhz5bbiVZameNOCxFlzHtfxzFOt8vfKUwO6ktlL3uCHJWz4pu0
r0FnvtEjOeSOkqF7Bhz4hZCw8lRLgLiZXezjvHxhFGs36hVsACIPsIyWS5wn2ivy
bsGxO1t6pYVQvwz4aLD/rrcL1sUEQKI/Zove+M/LbxW6ESDjUB1kfMZGSpq7sRE8
XFZ0cOu9xVWas0M499vgwVfV799yZlRAaybwLEy5OYb5/ZfpHDJtlCCPQDfjQ8YC
YFjBluSb5e8XObMu2+6FdRU48Nct34T+4x+IRnUXui/TD7uCperZNjRuNEiFt8t4
87jNB3oKfXyx34b/pDEDwP3dv1NllwXDkes3bZKxsoFrS++AGowyg40W4IzQ3PYY
kyHnM5XFnenxn3NeQBJHKD07u8rgIJPn1tcBU6O+DTZQqtGrGCdgiDxsnn3Je0xS
LkKwKRAHVZF+uR1cePOhydIHySuwy1JcwhfttT6VlCU/+U8a0kw4d0HPeXa2dUM5
GbVZbd7w9YBcmH+yrbs7MPueYUyh0U+js6wf0tDYRdbkxJHSFo+XFWHwnNlKLrhw
eB3+1Ov3WwRHUmVdOtGZ+vZq/+LUn/5JiYVCAsERsH8lKJBwkCBLNxubI/slC/YI
XaHR1PBK5SpmyWS9UPJPfxHXwuLiVO8aKg838lKjSdzD4ZYa7RdA4ig9EYt38GsF
kUcDZq/8oSuaLvtyjJD0x1b6E3hHjAcPiTWLAy7ZP/Gpp1XlfaY/RJjEYa7MSC6H
MzqWZHN6kWBtmeSqBhCD3eFrKjwEq8TtaZzVWRr8/Js/qLARfWkxllq30VjBpm0J
H9RZKPNkeYqmoYeTnDdILeuzSOv8NyGAnirFFI43opKh3Li6F6viNypuC8xidDJN
3fDBl13GNWkHasIJ/U50cf1IrAz0eHmZKd35lKCg3bB8VqJmQXj43iNfmeAzHbWv
Vi4hunuT406BXmRFOim1gSyDnM76lYzevrFFOsX6vctZUIVS1M37RPNM3ItPLskc
McdPDUExYbg5o8NFCTQnfw2hyhqtGHki67gTCgkr+rdF+VWZ+zOckFtGZXfB+qcH
z7/TNypNMz8kDZ3SsE3q/zMEbI571/98FzcoKqQTr4dfKjLCm0yPn4sOO6Titwcm
2pc4kX56DkgAD7i4dmHQnEqdpFhMFQYmqZXL03rb8oSfBgtz99DXTCWz8i8sGNzh
3I/ob0Uhkd06I1dCKz7DgtV4XYaxVOtrCldwztn0EIjCIYXk+OYnQzW2FeH0aJH3
GvijQCcVMzWagpJgmIWsme9GtddkbzqyGkoJD4FNrqstrWxSdZPul3jYp7d91AX5
wLlvZS20BIjfYbiwvGc/0H8mq9gccOCyvtKoTBr6BXljexjoARMDj6YHIFDPM+3r
7F6rHovrk2rgKRIt9HRzUsH2DhwnvGhXsl46Vip90pUME/Qmn18a70ijS9bc+F6W
1GpVnIQqFJxosOSIUJQ8CZSPki4C6t4Cy/uXS4pgkCkSx+5o7Jdf/R1Zzp6EwtjD
a3rGE1qy4y2MiIxWmwMW3yisY5vx7sqpGKdFC0RxK8UZOVE9B+Uwtlj4LkbLYxQv
C8Z4x7WWhEs1u0Z8Jx4lqgjL99bEvYXQVUUn+eXB5XAsijxhjhwAUabhu2a1z3te
Vk1quK3TAtnAKrBkDFYIiYVwa6ZkRn+/A9b9n/VZ9rkI0fYrDkmJc1wfSPYzYacC
fP9HqKGnSiaUsuZjeGk4imYhmffbJ4TUzjlEf646mZBFI8lC9Xl+gZjb7VhE88/s
eGlIqoVbA0m/+ImBhDQbhcmHyiDoCLInVkJqQ8SbMDu1R6nDDoyQSi5O1QXE2NsL
3uxlfyPFKHloo5L/TKsJFfcrwUjyjGICyHBrY8mB0RvhX2zEZDdSKPFL/YyAgNr1
xSklY/+3LOpENuKlHMLjnK+SBhuUJ9sWGoSEphC83YQEk5dHdvf8ZddZ8JTeW/Oe
WECi+Dft6U2ngp1Fu6ZFH5S1R4AC47QpVm0jPSxjnIfv2BokD5AanyzMJWdEdsuI
9vuJwlvQpYNS62IRHNa+lFAEPxrOOfVg3r8Il19UGQmqoK0k015rpkdT4DIxirsa
KYOSi9r+z0KWPshKsDmILi1pNvD404Rwp6jF+axSxZrZ3jvZWNjjiKyr8AdR8Tc7
CVObY41S+aZBJ12yai2C1wxyvXs4Y3JO51WjackMHtFQXfRDlmnBc64AVaR/qLTU
VUXgf9+kI27Ix5I9S93Yne/s+wlY17QHqnzd6FoWde0H88joGTJisQwTNwAMZNBP
MrvBrKyRpT+yTlSGUAEVLmC1iIRTrVNEYvuOPBZ2fCT4738XLYCpzs/62Z9P3JEB
wZt1wiOtUFyFKZSr8mi6GNuxh5Zew2VRWXionMF9kiairk5+64bYSqUi4eu6lDRv
iFng/QecW1Lhrd22k7cSQv0vMQNu5XvSumqjnkomVxVEDJi2Addjd7blBehH1hIb
e+AqybmSdEvXeTudcDpTgU0zEorF/ykvSuY1IaHq8g+CNi6315uJ+b7GflemWMst
r0qkH2WyU40aSm/Q9+ODkGOQ1qdAdls3Jo6Npqqyrrxebo0QJmqF1cW3OMLsvXVX
s3ejem2at5mJ27t2w2GFuusxvq//ALB/A7FJBEBPc5k/V0HNzbXNE2YIJKsYrmO8
FO29iNoYMQbeEAQlp65wDZqFIEFjjHXY2qBjQtoJuyHaFk56e0oq3wHqBOnFh21S
gx4xZj10Bp2NfnO3ced1WG5g97Q92xPkjaN8Kusp5d+5D05cxIOy9dl93Mt+hafo
P1cHOpgWdQEG7QN7izTXQvm9Q1b33wbTNUYGv/4NCQMUsSNp5awZ7IoYEos0HpbR
BNflSP5v+554A6RhS6934Ptr+aDmCwLX335BdO7VBFP0XqJ+hbXRB1WjnCBzA42O
ffFeT6+ETLMNelvoaRuOrfG4CSc03U1BKetKaDpcGOZMp/ODeBK8djIPAE0gz7/Q
tqULvcVYPfFoWhqJJMkZQAinfbWnmQuwb08CNNGXfl+pbhLNlPmsfHhb/Fx2y5ae
n2ffs0NWsNgJO1X2usLx8Hl26JRa3ZLXrEzrfUS3BcPyUlimqj2mjftBuY+p/dsR
LlqQLU3INiiRhsdN5Vm8mteo14hYwfsubs8IkIZHiKvEQxu4HuJyECNKuhJU06+2
zep9SJZZNozmwV/gIhJmQR9joTerJx1hgHUKS1XgBhK1orKHUjAb5xYRTSLvux4m
1ED36QXmqAVXbZ9Z/RMCZ3Qui4jHwU/Ijd5wHGhmjIhlcEZ+YeE34DgEsb+DACAM
nBW/2gcdTSwxWQX13gm9IbVcCwOztJ4Zc2A1uswGgwH8L1vwKMIMk1+M7+g589nW
UrA9Z9EPRjDxeLBeMvyXQ6bgaLKm5AyyFjBe9WQlSP512dPeoSb1Oo3Fg9MpgKhR
iTs8SY5lmQPIo+7F+Vigijo72p67MKJTgwGM33d7TBwEVHI0EYnzmFURmohE1qKm
VO4soDo6ku7LEpqtRXWy3Wo0O7xTfGfGCAOkcwlUUUwCU/IOh8WI47O3JO0C6+c/
Eh0JghduDY61n4Iuaa+bzpiI54EcEAXD8zIhcd7AV5XERsikTxTN18ibFHAtRUaN
RQz47UjuvuZ/EnrYjJLG9n63E97xpvAA7YPGGAgvDp9gEgXbDMTWjF5XHow/dPZ+
3zpMyiQpAQeq7T/x+h82ncvPDGmQuTONHLgZQeUbXzVGvghLH65ejEJR0ORc9Qlj
IbfX6Tbx+y2el7ywzAmXr6lHSIY7BWfFm7pYjRe2BZn4/iiL56aN6xgytJQKr4wu
SXYP2HP6Zvmu2eAu6WTBGQVsHnGV35A/Mn3RdPgiZy802jDMVl8PpIPvZ9cgDiYE
gb5j8YsddXPYdcqGLmiLtRpsdgXnBxiwSplPiokc3pelr4lwCLnD+y6YxgwfSxsn
2YV9hSJT1cZ2hQijqIsNyBixvXhCyLsJNcDm26WVZbNIvBLKXGiyddLTw34FON+m
5eSq0aLibfs3nEPHiFn1JaSEcM9Nwfu10eRYG5dX/XOwL1hiBOhOBeQwyqXnLEld
lky8NdJYOJ2a/6eopC5Eon8IC4M1y9TYpQjMyrvSm7Q2SrdyYNIe3ka5lVHBVqDw
/6y4xZkVb8mvpPiaSdhI51i6cCdf+PKDTexKHn8quBwIJuzAXhalQ5vlFGzLsLiR
0a7Z074UD6iKldYAuWQ5cjeFZiamnSxnHuTeIF4t1L7dlQKrFD289cS7Ix1zUwmd
vF1KG/6p6SEYl77IQEmtsEns0AsQk4wW+R67sM/roYQejCwTFCIJa9v/UqRejDbL
bNtUVDWd2+j8Zg9n94o2QgZIUc50Lo02DzJnm46oDxEVQVnF8fkhrSeDHv5mu+fV
JovV1tHRbdpYriBTgpLgnHJv8MA8bin0UhQOf7QcDSOJ0Tro06+vIcL94MJ9DImv
FO+UWz2SjN72b5Jke6+vS4x0jT+KIk4JR43Hzs30bUpQN+/hcWYz7ajjP5vZ2i4Z
9O0GlIcPgqfRe6J/zNbi5nfm9FWcrFmC0ePNpphrjacHVsngvnOI+5blqB+Y2ATU
E5GQWMSelOSgpeB+elTCUQd8c6r8HF2DXf4I5LdTdW3+I/CeskOz00E8beJaUlfk
3u6MGLr68kXl3PyMr2MB8PvLEZyvIquXuA548YoS61cgI/D2vYY7PK5RRQn2eim/
I+Ha2jVoH/CozkHV8DMASZJlcyNeFTMrRrdS1W0lIKGRHgjS+QsyWLcCiF0fh11l
INi009mMkGG89LyAIxBGopUv3Tt63geKFlR/SueGOjj3FY3ZM5tUTbPG/ZD3pp9N
YkU/Ff5IcI0rP2uhu15kawH8GoCIyteaN4muvMQ3aMnjtHVacZlGkTtcftK7d5fJ
KcU0l3b6OhMjtuIKH7XzMC4FdPM6xfV3IpiyX29UpHYxB8J5ZOUbJhYlX8hbOBRt
dSz2r/0W+M8fS1byPj6SluemlotS1VHZKpyAqSU5FQZXqu9tvcDweObWNZ0lJMXj
C4TrqUK7Ff0ZqleZpk5aZi7wFLeM2NhQ9SqkolUwOaAaqGDpIuxKrXY1w7RqfxNz
oKZZKqzyxxYgJnp9CU7vtGbNJD+UBODb2CW7Dq+TI092bhCX9fDOX5+0a++S3HHX
eAEZA+Yt1Np3g84HSOYd6pRXiDE7F6VDj91dwKDFq3grebU3ktSxPxfjgLWy32JL
pYaiCUVSl6OZKAPuRiHGAPTJ73t0WKMTBQqMQBn6BS3Saf/U0TmGXmWLyanq0jGJ
J6uHT1QTB7j1WbcEUZ+I48f8aq9nLmkJIBUWBRnC2yiS3NyNwKZBHhI6MmmCUeHm
J8MCgEMPKqHWSsgmkwEbDtV65+oVTRP62GLDlQBJszwOoSgj3uKwAHs9zzCyUheW
yYym54Rqtzab4F0sQSTfhVsjzvmAF4gZKoi9MazuFMDGHrej1isgI0pDju3INy12
ftl6AANQTflTGL3Jb4/6RGhxlmDQIzpYjuIHWYxkOWYIUU/3xB6wg3sQOb1iAdJP
9nKdfu0K2zRAsu3Th9jn1gEXjKrr2UEFApxPskobP6Jtg7lTkhpPNwtcdWZ0rQFj
PhO+kFIxvvjUJUiE5lD9tJofGAozZ9zZzTYljOq2/uStz6gcDKSFbNRXMGwtOhgY
38yJJI/dL1qPGTq67m1aEp3uv30U2YTThn41PQeYqyRsfO47L4u/k1sjhQZxwz6/
5vTbCR208zu/hBH/YaPeHxRlG7DdPKMVNkkcDCG+cXXwaYURk6NokE23FvZwUmZW
hIJObLd4OvhN57dhyXWboQ2kqjtxWhAmyID3V8STJGTzf+3ko4vtGlh2RLR+pk6B
GyAHIfery0pGYKF0KBX6kZ27l+c8aCFLSUxeR2y7rXnqtRVJEyUENflQLGgk+G5b
MuHSy6IoBZ5PQkyl8tPvW36dzh2tH6zg26QXbfBWz0ZsDIqRMGDZbHbTCjs2oqsQ
Ezi/+HZriqG1PDfWUEM716m7VUruiSzyROZ0egkUxwwdeiEY0iRYqo/sAZE4hMxA
/AS4O6ldiEADPTGbj8vPdtQMJ5PaVFOmOqmMqhOxp22IORolFZuFl7eW3i4S/hgs
BZh0WlmnxMLNd1qikgywTuzAlqkwyFNm19T0jJ6/37LMv6ZdezkPOglBiLlLUU6r
ifmx1AWKtb+VIlFbY6pxuoRL4+yc9sfpj9Ya/acNjkv90PNh7453UQQLto3NbMYI
hAhKksJp10tZXDdZdEHbi95Xt3+RwLcUlZNn1Ub8GAxFQR4SqGp2phNaPbDaB2o2
QpOPcaJmxBB6mA/X3HJe1Mr6CSLPMsRP03EeYPQg2MD5LwEBeGyJlJ2qf5S6tdat
hZnRfVL07rGyjEy7s5zMocwaCHDS74SvYBr+ailYIA3Mh7qYmsL2E1c4Hx4lnQE3
cUGvRE3XSB5LHXF/+OK22M5UjObV5jKMsnWcjeu7AsvhOFZnDiKbhAImFFLhfeZL
i4hVQrWXo0w7te5RcscNqFTPUALmDzmoqDpcghyZUjIjCW1oekD4R9BiEHWJkspc
7OfIl0wV4Zs8hocfQSyu/BjJNorq2aw6jYyvwwTKKU6f7Zme+XiKJZBPpVhLoI+2
oosBuFQmst8z44RqwcQI0H5WkrRoazK0kYq6OfMBWb6FmYuIOTMJDwBUcylVBm56
5iszFATQv2Dh+5/r8jtSqVjE8EEL0H1gUpqEvzsuf6FNDhVAZPwO3AttCYDqCR5O
QSviJrGZ4XOpgihyFKPNbjRKG9/G6peuVMreD1jd+Oy0BsLceu4z/2JtLEYWIJb/
x+/fXA/kJvfI9z898a7gmn0pkqduHJ4ZEMq3Gd8bdHMikSiXeo7FhbUH106banm1
nl7RjIhC41dj/DY2K7asV1qoQglk7tuXKeXkm7OSAzX2dEqjIAyhwv6DoFEe1g1V
lBhTivATmSMTCbDHTzfDhFf7zwW/2si4kzrXmZb8MW84booixIrBwnYdFuXPQjk+
3pJJOEKe4DpHZZHMQkG2QPJaYoOCunUMEl24Nzwo/yOSTYfd24Oo/nj/CEjHXQrM
JVLkPb01UcCFO8vQzZVCUM2YuzZ5bVDHln2Ig4VJMINYxldv3XUGx10JFRUGo3qS
2XpH4Tvc7rufqL2FyjwrwSiXG9EBIkQ6byVwAy8nIK3WG08wfB9gy63tWwxM3qF+
Fp4Nm/I3JKt/J2ruitVYjbLIQjQJ5I3Kvn3ySpsxAaX3+DD6gpq+Bu7/12mHIQ3E
WHD3jiQ71r0/1iC0CpkZa8Ltl41xx/85/vE6MKW+73VPbSuf+pPF91r8hSHQTWAz
jcDvfPXFzt96FegyYAmuIjq0AqJHcy9FA7qJ1PVMWf1YhZ4IZbpi27o4XSj21y+E
9tvdkjaiaceM+LbFlnvfWdqMKa1mtV+tHPJS+hZXk1k9an7HSfjPMs7M+JSoL9OO
4ORcb5JxpKxv5IbMXfyNRXfe7a/Sctyxb1P8awWE9Ye7WBK4l9tw+UTz/pMNruVJ
/b0kLKJvDOwnRB9Pb3I5A8cGV+4z+kduQcdpAj1D2yjT4gbCxBXva3YVxO8YXO2q
43XbpcDxSQcTdFOOn0uYrSW+my9vE4gsRJfy6k8w+6s+LsAP3v2i1eAyFTKCBXWB
TOjqN44JASNbqNsUEl4vrZxayuoTKPzXyRzAOKu8rOd9VmU6fe6mSbsZQQgGfFZv
oGg6F3i5FvW1ZLgC3NkzbzRGHZKAbRqaeOkrJjKkAsFG78xfv/bpApMn8aVb4FRw
u8YjEXspnrluo92CY77pTPbBgC/ynJweoO4y/MdjE5GeZDROl3pajL+7pIvikXet
z2Tz4XWqt5kldjQMJJJzA4PugDQ9Fqe35TkbwJngnCp8Fotv2UKm/1U1h+Sio8vh
g8ezIWLZki/0hFZu3CaPlZX/vbR3x8NN9STO0FmfZhYjO0HzKHDHUFpxdlwCqbnQ
V8PV6oJ2npQJyNwYteirfrqLMLHMwl+Nn7CUSB0eyGDY3XID7wRnduMb+f3UqNsd
l7dComTNYk6saCpMEIXJaRuUM1fISLvRTBqTNyzGuWqKScqZ6vmGwbYZPLRi36+s
jL9MHE7L1yF6FSeER9MMneE29C+D9oo9ch8cKfBHkqG1jiPJQeMcSGFoVvA1XVQ8
SIkQhAqDe7ISThGTx1cln9mVBcjVHD0PRyPaZNZgdtrRj87hJcPu8vnmByc0Bh3W
kA2UIeovOIql0xs8zzP7Ta4mZnTmnkCz5FsZd3g4HUQjofF3tXnAueh/ZhwR+R7i
pScEmFlrdQ7+Q64O9Rar7OCyKfE0n0EELLIJ8+FuFUJsJivjn6+Hpo/xlYIpjN85
zxspph9C2dmthIXQKPFAld2/dfCREFSyQrzLxLXO6ITkWFBfl9q3LRsCdhsUuZ1L
XhpJuuTSoYiqconYgOEPjEPs99N20D1/+gtw6O75Atm/g3doV4zaMWY0jhD3YrlR
Ns/7uALXNvxerR18VCrUG5pMsQzeAcOFFKIoMo9IJKqBw8t1WsYblAQdqKd/wU5A
7U7TiZK7VZV2oFpaHGuBQzZjIX2XHI5nFFtS2wg8NCy4LCi22m+xqaCaTwuOTTQj
mKIBeYrSEvNlKIdYe6mM4E8ChJ2h8MaqM3IwU46gXbosSgBIKRytjUWonGEw5ftv
LjxxsNZkdsJiR04Mr0sPgCs784apgMq6LPNP0NEKxtV184wv3o0hP1R18ivER6bq
SDI99s36foUBiNJd3JYXaYbQe7bUbnRhXmAnzKBKvhpJ+2q+7MGfbBquZOEhhGCA
T2XRMEMlsN9L7GFpUS2g8z0gl0X8jNIiyllWnoECGFaV4T3z3s3uEjE9SIotiEtS
DnYZ61LQemjuapxhgiPnqdJsrIZHNA7TEuR2NwArBthpXFxzoTHPGk/BabzDQmJK
YZ7OMvpEeEN4JZmEPlQR3OPR5MK6nUYEBRFWFbke2+DjHzfnByuR14axgxf2QT9g
ctsnXiozi1rirMKLnCuj23dgKYSO/tnOV+r+/afG4hobhp6F/FLkrXegRZizW9cW
jFGxqUno/TU3IJYErANkGV0CMR/hW2DImjL4KI0hDtMjWxmc1KHfLL6ZWuYOH3s0
jgkAW2V/wciUphcCCKxGFD+/W+wkPA5UHdxs6LOCydm/3B7KaSKb/nbRsN2kPKPF
L/jXbgnT98RerbbhZhaaRBSE1GaFCHSzBDo467H5Im+grTKDmCfnbWdHXMmljVOn
99x9E5ylUV08qddUHmMjurPZCQTiWXWPMNFt6mJMqC1dUyGagWMSRs1KCxRIsWSI
+SEz3TMnyZwzg3rFSV5jpx+Mk0rdCNP+Gt+N0oHmWKLLW+0d54Gjj19M1vili5cq
aHOfz1AqR1q54ZrObVLyJsU2s18BhbQEdWPuRUgbFeymWjDRRSp6PvLwcNSb6+t4
XS8qpUgx8e+xdfYvTnec2FQ1zVqMKCggj3sdljp33f1dk5dPvLYT8t7QPFip/GAN
huNXi7WTzimKfAeo5k39l/Zp1alZ0NCu3jyJ4l+wQZQ1wyTJIFRfNwTOjBuUbZ/w
bYixBZyfAvZxfyH0jPlvRCeg8mf4UOstBIcODl6Ob21R1BYQXEgJZSzk7AklgIwJ
/owWtTwljAOhHW9uamIFnxuPlwd7EtIwaRpUAscKbYHNEiUaTwhHqPuQ7LbnWxdl
WhulTVhzp7iehCfaxO+3UKu06J7CrfSM7YbJCm33Ja50kLJheVysGGDT7BLFKyPr
UchRiiP+TlVmADgo1IE9Q4uEBMan5MTA37BOtaHpOuKVKD0th+uynvWtpRRYutJ4
OaqkTirQ74u4CF02jyYG4WSozouhJQqgSWXK0i0i19YnBLWWx45vCNaMvSJvPR/J
IRX40QAaOYdNK9nvEyirrxuyLPs8uZFesQXYToJt0wRDb5/CeZ6hqXzuiCcQZg3t
oHkuSKX8ANLlv7ZMUYHsSCJMgj9DkQZ8zznIhjfHonWnR0LSVd8YqYu5xG7rfxUZ
Py+/iF8lDHvEWwhfA2YvowZf84OrkzReSXsIgQAxi83OPiqoWc0VHqAOBsZ5j1qZ
KynVY21PXu7ei0FgykmtjRI6R2lWTUGOHeRhNViPHwA1gqVOL0EZ0DyWHkbZzBHb
AUh5PxvRuGXZI3Sof+XQ6YcEgIzjo2HI8LPj6iBCAYUeGWeqahy+Yj8CaRqJAKZs
s7RlyTIE46X/HFy1rj4x5OWjqcb9SJAfLuc5tDYr95aDhGam4+eSFvKkOXyTP1gv
YFon4C4e2aRu17lIs74eHCJgBJlMUSKD3tAshnYDFs0RlbmDzEUHEXpOfwu/AMKE
e9ZKW7sJymbUuHuKaRMZ0xm/wunalM41D6VYFQ7ehiPIS6TcJv65a0Y85TWXcUJS
bfavb+hw2JFUfBNhXrfRDj+mo0TTHOKQXhWxBcJK3F2f+kIDz+qm0yX7JiMlqjfn
zIrSHq0G1Eb9IURDKKMVodNL8p57r6G9dG1Rv9WAbHm1FNpSBK0N7C1YgeLQ8rEh
ZGWnHgtHvIsNQW+1RU+ryaaAo3GJ+321j9R901jg50LKJ06PLM51nEXLAuPs//JF
OjmkhexPUKJGHGhcn9/8F0ZF8jOSynMdu7Da2hts1GvKrKG3j7RVUe0ZrZhavdFu
7AXHYjutydnR6uX+p56nPZ1fZWWGC6zB0IEV1xBGDIJ4yyWSzlBT2u1QfHm1cTo9
uTrkmwyLHNdA+9sJCBOXAU6/t83xZ8hcajzg20CBrJzxLGWytCnJHWh46s4i3nz9
mBGFUFwhZne2cjK4uPT6mY9C4VALCw77MM0W22t54QpI3ON4vSCiv9XZlIZk3nth
LFL/0kZlTZ6gcPRHXfDhVIdSEvYJwVD8sXhnurnCKLIKJc57JXv7398rjFS8eFy3
2nEPrATaz0AMzypeOleod+tXCtUzWNCJtgYp++PTL3OK0ZXa0ycZ5Xpym0eFdrgZ
eNQcpTEQj1M5xp+fzEidyDhvY2Pf9SeX61OkKVHdZ/70kvygUAInh4JEf0TLuk7e
xtSrb7CxX44ER2PG9ZCoRIFhEv8v/f0XIq5IMLwY/p5iC3gbloymQ/AXhcswcqNX
ST78FcJwAD8S8T300MbxQhjutDc8+YIdaZmLUBc6ZOikf2qQYRm5z3ENSK1Olq8K
GhbL26vnA+Omo8P3F/tSS+2mcriM96eE27QxPtNgnuY9Whd9tAnSk15YWagNfyZi
EvLbsGNFNGDBo2G1b0HgiOZUrqxGgHzGyNXiqrLZT5krv692A9KPfuRHCpoUp5Jm
RDOgJCUMeKCGPn+Uj5N32XyUE3G3yJO6Hgtsxo9wlH6SzVMwBLDBK4XkPa7FyPkW
1dH9GRtYa5EfkRxNOi7iAIZuWOtR4aNb704Cozj/wktx6BAnVdxs+o++WoIOJfBO
iOFrNMiCOIbCJbWTKRZ2ZZ6ARgJZnSbqTy9dZa0abBrEUdR1AA31otOI8VIW46yH
NGJwcWWE1MobUheN7XCift0TUVsnceMrDrycrVOHvabxnAcX+rKiJoSOtzBJBjVb
k6SisN6qmU26v9TFFxfCxWSLSz7jCV1awPs/fQXqRZZjWDBi9ZIm+87MossttWMV
rDu7M2BaKMcRftNyAkqjni2i/Ms4UHHp6Xxa0edeTGnainZUHocIMNzYby0Te+5U
8+B4lw28m55wAHUhtXY3AS3luxeKnxo7nO6rQZx5Y4LK4MavxDvXePDKf/S80LSX
2SvMDWodROIr9hd9oSOs3zZ3Nl4eEwXFbp7Ohfb3+Pvm/5DOhKvuXmTG5QVyoAsq
Z4ETdLFgeuRQgbhsXW32zroWAYYGnwmZKykWCK15S8eaZ9BfkYA3OfPS4QNgAoTs
bpJBbVgKGYHu3jYFbfUiKp7PBOGVaFOAVDA0Uk/aLn3uxyTgMwsHhNeK6woXkj4r
0VoTDKmVj/hOMeDy1lp/6DDB2Xv0aaK176Fb/puRSH2mjhH5izYY/pArZZ3Yhvs9
A7jSz4nyKaljAzLio94LwBjPSPfjS0kpq4jPj4kYACOdSrzllc5YMNBtpNrXmkBC
GyEUQNGiFGZblp0cb4HwmH/8EhPDJBt4LS9QoRE09F2dYTx4jzmoV+7+8XZLXv01
rC6BuOuw70VufEqGvGvOvcwWzt4C0QTYdQR+PjYFlGv5OBwfLBVTzroP+2MPWRPI
oOoCovt382NULVPjYko4gC4mi2B/QYUO9A2IhdvxFCakTcIt53n0pjEyqeQvTmct
Jy/JDlaUUEC8+aMlHMczmpdauD25r3w/poJs1VYefCX6mM1AZ+Tf72QG6L9X75Ny
kPR66EAPKpRJFyM8GdvSVEEaVZpf5V2BNcR0eVer/UnW7HlBadnnnkE9syme3RZP
8q1aMPzM02UKZeIVMZILYsV+SqLNZMxOKjqYsy/z8DO404azGg2A0rVUnbP/uXLh
4YaO54WSs7ZHKPdQ/YGaZHQrwFXvd59KdFn2Hnnid/h1dG7pHuDShVI4SKUImJzB
1bUNzagvhDal1Tv6Ryy0g3AdGuwxCLG+Ad//tISFpYp2I3B6HyW4v8K+bxS8l7vt
0Nlzr57XSkucXXJeV7uHRJVsXAcNzA4H3zNVDA2MtNQQrzQHl2/au5mFnopsUiqe
v37GyjEMqwYcSg630x3CAOZXRCmh3VdweqsGtPpCeJI8tWLyvrsRoASaf+zU8gQn
mNOnTANptosZCbHFXwM5+hft8cukmjN8FWUVTNZ0QlC4oJLp7kF4GGPU6ELX34qa
KOWXsVm+sDZgAP6xwmUpXr4BxxiD77gyWMYZ31Sfu8OcIPHPuPlmwe0V4yeFylex
qpgekS/VDqGCSQI9mtz+THtHxdBnM0RSK6iD3p+GqVs7/R3wFN4/6s2yGTV28ik4
WTFb7yBKHC0ItnrYAKc9TVMbT2QG8fUhT7Simj7wYPd1JDHZ8GzTJ9UdNWC+hfmw
5/sU05Ey7h1j9i4Va+2+aBTP11pz4qMXbuvt+jdbQS19YOXJjt2CrfWJTg+eACUP
se5jS36vRhgr/Qu3oVPVBRNCrojEU5wutxyyJ+Q8yXxshlYcUzrnN4ixplGqxyIm
C4YglhYUVmLM+l9O52ajE2mj+MJDDX1TEaR+RXMD6drreJjClnm05J8AuJy1fhRp
dn8OXqPuLN2njtgvq3Si3i51WqVi1+4I5tNxIyqCzt2hPF+su0hj3kOUSblqJkPj
77M7noU0aGAKYcdpLR0uEuZUnKwey99v5m768oPm11+XxjKmIxauEYnfrO/Hedxp
HU3eClPfU2SRPosKdX8rPLK+xFbKdaJ3DGN+SonVta6HahfL2wvSYloJoFlsGVHQ
iTcS97pnUZiKwyM24bJpbo8d0J4tzJduAbKw1dzrx0OHrncR9ERfri4JfH7SqPDy
pOsqjmKCIMZ5+L67DlYTLjbqiz63oSdEeJ8Hnb07TorXkcoGb7sXOjflNHu3ivvI
1sAO3HhdIBT+7VMd09uS15aEqnJdmOU3wKdKGIGNMcQ17dgwaSjbgRC8jWM9wywe
vH+Lt0LB7rWk1ENZ6YeRtPCPajuMXPY9i62eabjvmmeipmb/XbX3xKU4i+4erVME
OIXhHOeK8Xv8SIyXm/SLc/W/41fVcNgPv+wCH3x/GZYbXYYjsTGd2+DGZWCjvu8k
MYm94t2qIz0z7qB6yjuTC8DQtZNmpAazpy9+VrcRkD4hmOmAotEiO+BIE+smVDwG
dLNysp2ZDe0XmWdWmZ48OdXnK4tBc38tXO3ey2Sv8p42LwicxgdAlpTVT/8vGieT
w+nq3HLpOjiHhR5CetZNGcmVbmFAQw/Ivepx6CCg16R6RPd5nTKmTcqcTSDSTN5s
rKKmn8BVgGkPDMBGQ+KOgCGSvMrxlhmYQ9pbey7vvdA9n3pbk2K2RfpqKkEao518
/1SiTsiCuFKlyWnIh7oXPAPj9FV3paZcdmDIIr0DLVQpe6PgQ8loqYlZYO9CPUm2
DSCpbURiyjBsrS416k+WenjAh0T3GQcte9v83gzIlakIrw+C6gEKBTpRED0tm0tE
x2EB1kV3GH5Y4pm3O019lZH9tsscd70Z/yqE77wynQG7mwOlZagWs3lWSC+CHrAP
Tg3CfZiR/VlrnrJus1zVzVydstr6SIu20ma+DYzO3YodIoP63JDxVge+ow+2IJge
Mkh+fxZ6gVoz0CC61iI8f2vTclXcxJwiJOiYGy41eSeim+XqVeUrZqX9ztXi4dh6
1Jzy6tS1+JjMMeYD4Zm5wie0K37qaQLBeeJvs+F0ESoHoGutvh2mKw4mPonqLPOm
P1trZKrwBpwCxtG/+MaUonB+Br4ey4e468CyHqTex12zODFLuKTiuwj0U9BxMcN/
cUAbKif7NHGSRpHegqgKYZmDVtKdDexgOUyY+wZJccRan6J8eu05M2+VAxgPfjdF
/F3tBSO+/EENOlltF2ZitIo+eZZ0T8vonTt9v5Iis+buhuK/8gk25rfVpq0XGXFu
F+gF9dMZgGU4f/K3oOZ2pw4vf4vPhS7QPF9azsUkOIAY07vcFt4WY/dJEYajSCZe
MbR5SY0WPaW5jRkU4rbjd7KehfiffMBaOLe8i4sPx/qG2vCkHFFHXgcMg57Fbkqa
hediUdJNgrfDGAfYQ5KOxOxjziaXhQvuHx4VKNdR8e2ZvkeCQzoCa4/1DLK9DWQQ
GlPq5BMq/th/zL2oP/1bYGJ87xxfd+I5BLdq2FRK/z/hck5F3BVdJE/di2Tovhza
5F7kFVcR0fLIHnsIjbvVdk1c5iS/asMo3NJWvcdNTGDIP6nH68saaQH5pLl2vOpc
Sc2z8HreykPxUw0hseKNXIgP/19zFiIS+wTT5GDga8CYChJN3kjLfmxGeQWPlKhn
pXNzX9lcL24g+KSrK6HO9tU8l5tXNrviHdUumX3WUe5MKRExmQ7gZSDhYCZM2oao
md+47zbsur+CN+LWQgJgO1QdPJiKIWuqkjdQe2KINXKpWytsYpywBdo5wkSZfFv6
tNkGSPiq3H4MNxa9C5P73gRM4c+DGOqSHCr80KoYPbkooQxpgBMJ1Sv649C9EuIk
41ObaCbPOkc2BDshEyP9TeMaaaQHbNVv/4hYBFRcKL7H9UezhyWZZIMtLGw4Cq6u
TpsovBeLodDi8Zj83/zlk+ANlikTlhLDjKDRV0Z3sYfa2XsuQdF5FxmZVC1y7MGU
bobH8iSL9DSr1z2RAA1+HSjKNk0dLlI9qBjo3YY1SC4sScaJ7HLNrBO3RmNrJk9d
2Adz1L7XSbohhkAGjPiAnwzL51vg/YNgQmDJz5fmKXcUTTVc3bLfey4BMUpwZQ+0
Edv6tiYzvL2aKjB7WoIQJzV1anWkshCWJxnnNGqNXxnAXCdWrRlCpKkQAekh+bJc
dUpb655AXGCTSAunMhDitSml1jbBXMKfvbHZ1iV7Jpj0YRl1wRGgHT95I562vT00
HR/8rf2JK09eRMVyQa7CO4URVGn90K6cOAPLcRDq6DmoRsWgovJUAgvo0lcMFXzh
nGDgWM9rw7Qvn6AV72dn/6kqGXO3VJrpUJDZENn6mJIsCa7VpcKn64eyu7V1CDzi
+GlVmYqvy1LOt/KsLQ6VAIJCTPMl/HdDmzaZnlw9mgvVB2b/Uaucb7IrSWhUSokS
v3A6uAyBSX6GD0Jjrktuuh3uBzL3DDtvZ4zZimWrIRZAtfk2gApjUOjro1QzLUPA
il+xdG0bBu1rp9B5pbEsFR4Znvm5bngB1IC6+7QCgofqW8sQnx7CNdw3puTWn17+
16mK4McJwK+ou+JZkkzEQt0VRv6muEF5fliRwnDq2QDgjXOLTf9L+UJ/1M0yOl2G
lUonyv1RPaUDybTGvxtve55ywdUXlc1C9p1rCQ8/l82K93DRNAX3afnk3xCsAa1a
Dn3IjXZCElDP2TX3SWoVUpdC+839VQRRZ8Tm2vovw17npbR2AkyX6EIZcCMtyLuS
G4s8Uy3qr1ZagoA63xoPdOl0JSeMpEa/Kn++Yufz9VGexU4+/SSvYb3tQRnuOGD2
QeiJjrLcUUewunOXfsrfet3SAi69ddIMtYjWMljrKfQ57DIRA9ui8BK2h1MxlANQ
m2ef8RPIY3Z2TLypsdIGBqduF7TUvkXGcUjIbQL4ltY8lUsxKEuWVFKsfQ99GSho
Zpw5ypitRpZdUYQ6Szf5uY5fkVe9E/HIeDOLOWh4SixWd02XSxh9vUOLuD7McHNf
3PbG4y0gcZkojFQh6zuiyBqxGTCNuJZHAAY0rx7MQOvwWfp55BuLpknI3Khk2RTp
XDD0oXFfijPnZ/nT2IpCFdXsjELodYB4sCVb+8WD6F/K89yBtDKOvsJOr3QSHSNL
By0n/4kPfNkMP74SR1eN/BTKYBjqEBMcv8gYRMMhgBAhT0XtZTC2x42ZJGhMWxNM
VaZ7r7EeaOE6UteNbWa7XpghfJXAjSzQc5bwCaJUZS5yejQaq3JS2pqAKrt7NsYY
+YIXdKp4GMtBCrmAElo78kK8ouMNcz9+Hk1yJK2KQ3lTL279hzTd2a13iio9AxRd
N9O3Oj30xUF52Wy7FpbyiY4VR/0AoI2Ih7wxvYXlAPRPVeNJkJgy6vNv009ICpp7
WuHp9JPJZFmIAjxRnNsdeKZXBcHBNLjSQjO1HgIinCgpIn7Gwi0BXb2DATQulkAZ
LHFmu3oSEDvEK7tGL++ZBHlnmF7p2aBqx+98NB8xgc63VkNkH2M70CIAQRNBKdex
/kosIy+MaFHOo1BCfn3L5sePyCGTA2/dvfIU8DkqVM19zggrkSTxX9qVZHUfEYuh
G+xiW2oHoL9iq8WyTsfLgCATJkml3uonsdXIVlxo719nKRPQ2mTLVw2BFmVcbjxv
r1KCs4E/b9ZhKqIk9SzUMZEOtKjwvgFjwUPL18fU/0n7xdNowX760wF9GAiUkIXw
0N8KxMRU4vgk1oVEu5IS0Z1sPIDnhxTxYVdTGGGom9pe/xQqzMEmRkegk8rPN304
se3e9L3ciTc26mF05gfn9c2odXqR9O6MRC+yWmr3XUcqAO5AbO9w2yGrzNcp6oWk
DDhGhhNjG9jQdG7R8oe12l9KmLwi/I9M139lSgyujAHSZi7p1BjaoIHIpLKwYfU5
XvvzUCzntZz+z2GfKX64UXEBIkyUI6yzqR5WRdoJtOvLsoCru7Wf9hGmXuQmkyy5
9NM3KmUPLmDaPKcBA6BeErhClgck+eJHuUrD1Bkw/A1A/VjUvz5CTE/j3BsRCFrQ
2+/rTz/ZcI9a8MSlSawdpzIUSjlhIfxsu/wfFW+ohpgb5JYwRhsss+tWVnOk0Dng
Haikxo2k3Orynv06HukvBpEQohfKZQ6leJqRKUbdOZvoc+opoMOXCpDxijYoq3sA
SsZV1qg1n8hKIeg5ylRp5KqDeT988dC4ZaTX6OdnFIJ5DuwE2ejREj8AojG8W3dk
0KaSYUDY1SA1QYMR0ljbv2s3zErqQEsPJavKSs3uSzma2k1YFWGrLHKwur+1nNNu
kz97LD/TOw5Oo7QPgoIi1uZDnVUF1zdkZtLmsCO2h/fURin0bolLwl7cze5lHOIm
72WWwC89lN0y6A8nlc1wBU5uBfQ+PU6SD6wNShkDyiqjRuz+X5gDAIqzKsiJTyOj
KoVHPZysv77SkS9rvbEyI9T7zaYkidstHuXt+W0QA1YXymHrwHmCirgi8bNYcT/a
tjvd3ngaiEDgWxF+PxwFZVGDkDa0VEooewdOe1CB0XQrbvhW2BTbV+Ud0NYwCnFL
8Hw7Ud0mlJMkaq9xHCN5KjjojWUNogyD/IRgIF2F3RorO/Je9qAYq+ULClmSyCRa
5GnGDjgqSDxugYFaFPsz8JYjzaRoKBiLh+E8dBYdI5gen8kMvqg2dZQPoPZ2ty+w
x5V8eh/a6J5Dl77yyhkK9F78OiZVgrV4jXOspWIuWPrD/WeBXDwqMyCCp+cIBb5V
N2I7+8foUPXyU5MUbyNq6iEDIptJ3blRlISz8nEoHdCyCUCJdR0jniKD71xRF/zp
HE4v9HvYGrD8S1MyoRjRsZLjY/X/W3XNBlyjMTO7AEwaEajwUWcdhvrGQYOY84dj
2vV3aWlzLjcBuvfUEVfNKoZ4zUFh1LlIq0AwApsTh4HALwC9/JQ4K4b6LtdeqKC7
MpbXshO6P+CzW1G9S2knR6Vj/uzRk9epgcgFx0NCHAclheJcvSmRF6K9Lklp4kn3
Wi/EOcCa8/092jrwx6bfe1G8jUPClv6aT/Ke3qARVCn1y751I8BFT+4ChPHIXGrF
4Q2Q6k+nM3LjqySt2ICvC7Vbk0O4EGVBHPBkEamKikr81BOOgczQR63W456Gmk2o
3HIQQgveo7pGZ9SPMGkQcPyA4iUpAcrIijL4AUcjYAJ+apl6G7/fPt9gXh73Fc58
6F2kC6F0gdzh4U1sSXn3FALsCHDjrgvcIxx/Wd0L+8B6hmoHdFLjqAqaDgw0Ubba
UGNNGHhuEF3BuVUoA4RX7gcnT3glEL+DjO4fvXA2I+sDsuMwhkNeYMUK39tx91A9
Z7iivMp3JqDVJmVsgZxieNXdcLHzB0l27DI3GpM9TS/iIkSgSdoN5d14fLqf9IPa
PbykcC7A/77Wd/3gbj6YSrJMvHiz7pHuau/SFC3lkfRtR4gC5YJCCdNCD3RRqDaz
53zs+7OkqArGbuSimL2T4epo/G6pCZloqgYMDIXIgzawC37cjcsmqFv+W3gVcqgJ
Q1Y8Vmhn9AabmMQ8HXbsgi8rPtTR7YwT3+BmfOOSZ38zCBvZunp3ZIvYXXAUC30O
bjfjF6OoqXf4lpOaR89wQJGtL7nj4kr2sWorPfGvvVP70JW8xC7z5cHO44J36HpW
Tm9A8IpNsVN8kp64+l0Oic1YN9i01LneoHo44zQzi6HaVmWj5qG0AfPxy81IARJt
fWIcM9yzZWVm0BjdcYDh6TrlJcp1zlVPfsXCtagku8UEdbd3hK/kE8oeBN7uSSJq
5+LF18kUFI7mldaqd9FkkYGSyoaitsEPJxtxcqYsJZmlyG4OUgfRZMHB3HYiPQvB
BiGDPtXASj3NOzySyJUm7W3na0eK132pw46JpLrH+mLqO3HJQXIaKDJPJ/rVYqU+
HKCtNbrweF9Y4KBeY3kwgLVp9zfLDBdvogfOuF5M5UyvqDMP3fSv1iqhIa06+U3D
Sydpcbsm9oUAcWsYnpilvxSMVwa5gFxVLDLPUi67D+XFHTxs2W7oyRMe5YV9jET2
S0KbM2TvrNBaXZ8Fx7e1k4EwtbJtkqhGR8WRzRREHIdI6Msz4R2epkmuyiuKnlEY
PggJaiZI832bMsFqfcw6YH4kYtxBM2ssH8A9lMtWZ+IDNJQ81wz6BijW3ZSsk1p0
FMHthnOCwsrQvqI4vy0Ev9MetnCE5Bak5FukZNuWiWthhUw7Q90FRjg+GMkkFo7x
/cQG6Apl1oVtK1Ph5N2a6nI0NlvhIuRg7LaZdTmSz92fjXLD/uK7twvwF4JSCFDx
1f3xczJjRPf0YEE0QxqvI+U9CmIhjHTPp6joNJXMiHUw6j8HR60kk0682qhWTbfX
6W/VkPCHK4XE9ym+0mfqGK94UXAjJk246rPeRMcBhP0KAGV5Y48/0Tr5miQLcDyx
ivS31smkr9xUfua4LKXayGrKk/OUxXQNIFcV9wyJI55j1h6Tubhnu4mQTSlZR9V3
TwicTO+N2Golx0vwldsGtpzEW+ydJj3RWlQvtSh3+GyDkwPk6XN1gXXzvI2A/Afd
+gwjuYOYaD1Ecoz/q6Lz4ninbBNag9q4JtFl+BcTOMmuCxNtkWHBDlbunpH8mlNg
HCBR8YexxjfgFqvg1SLtSXlQNw47Vdd3a/8JTgPgqY7fimm2NhW731gJhxXE+xB8
wnAPSOP4xITChRsl/WX9upcmYycxQx4DWchBKGBXPuj7Vuq0LLxCHVpw+DSh02i/
SWiD9NeI6Enbh4DK/TRCprb4jAKHAy65GMmbXPtF0fwSKySOnvLg0Gb74Xfmm0AZ
+D7QLWcpAtE8AWJqK7a2GSrZYITP9Dx/eGi8JTWQq8jEE5s5s2wcMN6js3ZtvB7y
B5UQV3vrI/O2wzM1+XiVBaUlNjERsmYdi4iaF5LrQTmCWszNGA7EnUbkmH1+b3GX
Q1K6r13ehjeNLDTIpMDsQXpbNXqvMVFoVJTX/J9GjU3rdDoj+p3n7cPnGy5XshYo
B5+ybNVnzEDoAUAno9pZOce+7vUHXjy2MVa2rGFmmmDORyTZZu/hM0e8WJLpRm55
QBPsC+xEzKUVUPVL7l8ae4e4BQm1rqalRd8jy3uGeIZJMtk7QHB9meMmDKQnou6F
77h0FJ39kdsrSGKB1OzXkmmfA/4H22qLzcuSOY1T6EHF3oXngmTIjs+zFk2wysel
H0RUwQvk2EVeXwNYGkYVQSDp31/NIQ5n8URbSp6puzxBiH2gOVHChxZaVghX/Bea
DH/0dT/oXPGOTsjTZYO2jI6a2wYwPzdfI0BsFOHO+jm4IwLOIPrafBagfqIVhOzq
riOMV3LfViEbOhYw5RWddjcLTfuW/9uPOl2rHU6nSXVSGBOm4r7NDInmaPy3bLzo
HvAPTvOIsC+pY1xucfRXoxYdcdZbcBW/DBPCnJqFm1WTEhl/CoSBgiXm+y00gg88
ucrO/VPFKVbGHT9d8X+t94l3Me1Mkau784/pAgN7nX4pXoTRJYVYpHkKzNwUPWN8
YVwLnvEZ8q0oMykHSZtxwmFzDoXjvKX9ij/bNpAm5k5kPXcQASyVwn4JZ7wZ/v9S
1i+GnYHxqJeC9cbkXSGbVSWJpgPwCF/1824m5F+zqQdS2J6wlwf/WpvIjseHzvBI
u+1tnH4SSgg6Pe39dtFYRHJiX/DF5LTA2/liM+1zX5tMlQc3i6SH3GCwNl/H9m4T
2kuPX+1ODBntrfRzUNgI7704UJktQbaWnd1ngz/IZN0epeeSFnDTgjv0DVxuFMkL
whNkR6SrOuayBiTMTfu8UCPstewmgcVcl9Goobf1VEXPygdvEl0ZRRDCaEx1NAxu
3ht5yvLFJT0xoeR+G+0HDDZFcwVabl3/p6LTN7iNnZDiASuypJMJGXv7HtsKegXc
iVTQfoVCNJtQt3FlDPmUjWub9hbfEsdfRW+rtPQNYF8qwLoSMrRTCe5AyivRiXb0
hbz2odb5C4ACW5h4XAoIbwPzJbqSrUp/eJ/rGSe+2bnrlFDhRAvIxvg2OZsZ9Zq/
TH/IUJr7VWAvCX+r1h9V9slalK3QtBHNSAYILzokHOIh9hjaUNjxi47Zb1FwiM/T
jmemkYDbeUMEF0ij3eTJwnpPXu7mfzoCVH5L9/LHqbXVCMTNVCjYuf9E8yRbvNW9
CeHkLRd1NEQ40H43q84i+9lnZUYiHX2drYJgcvm0ErlfmvaXbjGpxBkSHpEyG7Ir
5EMRLiEJiJz9KpgIV0fQ+g0Z1FA0hBJ6qw+FjJitCdw3DZMpGQrAUitpWr8SWnC/
xnoi4DbsIDJ6Hb1BSpPw/7Mt1hbNpUnBcP61CTBfdHV86CgA1EXXoLsy+Uj3lRt9
StPOqZhIcFboTYFSTnhd3/G9uTIEElsfQJ/m97FlS1r4EAcftkjl3Uy4w0UsyBfS
SrXjpJLFxoywEvKwbc44lm5bMpeY6i7gJHFFPLJoldDuZmGFSgfOfsjOoBtCIEfT
SE1Ulb87r9IvA6/nbY6Za5yIh7whwgx9ZlbrUcuu+GlPS0nG/17kuAQhKzQF4yL2
gHgtiF87kOtkZaBBGU1CAUhKMnsKjE0NzCSturLhyoWPnINlhYnPq+ZyodpdUXkO
CKzgAMk/lYi1Gh5Ht+Ds6WqeTU12YahlKhNdV7uAHXafnhb26Ml1ezb/GiOkJnv0
mbAi0kiygJw1TtwTXuQWh3+8NwrxIQxrE7uvOt4LaZJe6Q2ssh4mbKjkruE1Umop
kY838LPRb4Rs8jJASCfbmFRRY8VyNgdsri57k7p7BRm6mLAqQzf2/kDYv3QOOHtS
ZQfwCYMQQM6AVfbWsijejx+6MKjm8f0YseuGiwp6bhfHgzw7ZjLj3zz46yRoHZCO
Wefx4Gi1JkHNevYD4Wv+O00AVRnY31JN/P7y1WBAzyxEMfF1K6GO112bKcoGi4zr
yUMArBEcVfkWpaeojfeCp7aQvz9Evu3puKbrJw91P4BRkfXrQWdOb50dBPsgYF8M
X4RmllODzJ0YPP9M9Q89aakoxNU4Gvi73fRG/DbZAw/xHSsVI/pGbtte+Q3Pij/K
yAAkhxMMS98xAoq25BnkK/YPg0yhNCkMHW1A1aIj+n0Aexshwvpj38oReQv6Mhur
tEvBFIGRKWj0WWAOqfkLR97903dgL7ZT5Krex23yPaMQTlAeqJmoeVlYC8wkFBA9
aZdFQDL9WcAHf3sGswrYYalb1CbRTYP6Jb3rwUU2Zr49/x5XfnTwpYogwaglcrcc
c0QfDct1KHrMux88oMhIeIkHvMM2UM7JxlZFelMmd7Kd0dhkvWMqXDHh33MWBjiN
P/1+VnHD9S2likAdT3k0lhDNoo0PleyT8b8IS8BqvNzI+aK3rancZXzt+1jS1KoI
etUIOqPePyDgmd8+QupdFiwF3q9cyGI50FXx6ud1OZTQBQGETuDRFjpWc3zs3FKG
FMCt19Cio/fRYeiLhTHRTsLNZ6ceERs+DWCx9IWqrbSx0MHtkR/K1Ne8wiqjPI2M
IWiu6HQcPge/4VR5wktJj2nkd0Z0spst486bF6Cu6b7/Hl8zmhqm/bOvPt8m/46o
OT5vu56IU8Yx66LCiPYyq6jhDEOPS2sDihfRKAYle3SnKfOIuUGf/5aYJDcxrOu6
KnIY73GhIsTNHIPpRoIYbpdBsWi0SrRSTs8m7paU35nRm0DHc3meQYbwyOIaKEGb
1j1Ea+mjlnhRDCJnSYpn76OflhTtXeCgFFme79UZtksFkPmTH2YY6cJYz/sD1a5h
oLvsisROKSu2OrpFMAvHt8GBroMJq2bZ7fDx1yZZxIwalOk9kYGn23Sn8aXh+n3J
NcEQh+FGMYUaWY0E2ypA7nK3x/0Q7/LEThAE3Z7KclBSaDhcwRf10ecdUxFzBew6
VOEjThim/QoEIhF7INORoc+SkvUiZmhQb9zmpXqWL9CKayg+fhZjmoi+32FAozkk
a9yqZDlFAAaEHd6G6s9EnodeJcgaf3rs4dHTb7NRijbk2kmzWTvBej0+ELUdnv/9
get7iM8Gr12LXmpN+G0jamptm6IC6jh8FKU6H/nUATUdbCOXEXM9v3sSKMGhOg+f
AvbZgo7lc+7Bk1iQLRKObPXFRGbDefwNpI9v8grV9yoxISbORRPLl3xTBh0vrFy4
0wDWLKzROKlVxs/sTFeYz5Fx0QJwgPouymHdfRO6pGKDBLYa3hVm8J9x0VgvqzVk
1A+vw86ThggO1LT/c+CM3+w7v3/YpIQAD/YRfD69CiC3KwxOzMeQIF0vGTYDuy3e
UWFAT5FN/8n/HPP+e1gbs+N1HJjThFS8f1IEBo1E2Kf9sDLYhQIT2RA1U5gAuL6S
xCMeLZPpu3+Vfopt/mPajgiP0NKap7pDjTYx6FxCwBqj3XVY8H6Pe9AHv1vywQDj
taypJ8w4Q8vM/C4WQxohC20PDwj+5IBullBX2As2Gz1jn1TJf3hpdnMCSZmYSUui
W5AwuS3y1ww/oXd9XwqvhkQRy/b1g1SumMkGVcdu0k+PoPNX2kRGDIK6r+27+FrX
8D2vcHKpCfhF4XO09hOFKGYkwmCidF+gq3Wby14Ns7ByiADxSBca4a22jdx1LP0x
mRv4aAywpGr8ZJVGWaOzqeePetHy3nGROQVmLGzsoWf4z2XJfEi8/KlEPhJjrSwi
5mIiJ1i2OPNYvvR7XBrUfP8QPEnBiORExuCPKVqG5iwgP5Sh6zu/UEcY2x9coDH4
K1Lv6UM/1AiWLhQH1RVpehH7cwdbRrZNYscqxRscG+arUfx11o/pTwbj+6YB1/VY
rxwfHGKGQFjaEOfXDAwQZBAi+6q++2uNcQKsWl4ZnYJ44vnXvRmhIW1aKU+FH+K/
GJVokYr+571BeGKZV+SxTxRTKMiIRKkQptqBIoW5XtC2TuX4OlMP3WmRu1kr/m6r
UQJ7hZlPI4ypJ3uV7EQI5IJ/aU90cz6PDdxFQmZCsF2VN6pTp40GZ9JPb+622F0c
rH7aehP+xhDWG/MBPtTHpj4GEJzGASA9CirNkbo8L1L0ZKQuJyzTXheQ5CFVI6vq
/G8nT7YEHy9j3zMkyZa4fgpFrfcjimLl8rQlaN1ookoE41WI2HLu1zhOTmIOf2kr
ym1Nxj9uEwj+P8o/elUSyPBV0dbohJLoMMZr1MU9fTO3GPORXaKouD4cGUo8Sum/
Qk6IHtmbMlKphd28LW98N4oPTcgbtTDS8llkQHr582kvUnzxwyj27MgqTFQj2kSm
56kfx3UUvrK2q0FcekyfjD54nf2ZHgny/cdRmAhBKq57Jl2JArGaiKen3uEh4xtV
eWfyKG4E2WX9bVV51lfdBhOZGPgdsFH7KeBRSSAfS8XcqD+2vIHoR0f3Ar/wgivI
1NN2yfkJ5k9sHzowfhReav+fDW9JQ6bgC1t0h4pipSX7sD2a1ecWGIGxLfYv+H9Y
cALk2veghiAv/UvabqO6AAQUYWvuRpQqjf7FOkliHmb2g2l9sx3y9QLxom8naZRd
/Zc7ZapQN80XGA92Y2YBaXRpoYpHVvn1zFyNmpOZO+wt8u6wAoSAtMKc3JKQmz0v
KzfJ7feuYDlUmWYCXDbqYK7p1ocopzpLv6xyQ17m9gh/8/9M3VFhU95L4ISml5GR
fziJECcJCMFc4539TwuXLfGfoSfpbZE/vn4ytmtEgrLecX5MdKLIv5jzY8OYQUeM
ERdt7Pd7zbIER38JRzY4hl9b1AbD76eb5zwSUwsLkRcl8ilV1Il2a92599x5bUjG
E+bVSzaWsA/4FlT1HeIKH0PUhSATA/zMX3x3xpbaW7S5Y1e9uwiygkYF/R1hHxqW
nLl62nKfC4vQbvydHt15jsJ0Ys/6/qpplOZ9lUx/mi2GYmAAN9pm9RxJwmo5uLmx
wYBgsDkwgTu4qiLq1B2YqUFw7Vkbw1ayUCg3G4WFKvKI1G4K5es951Y9Bw36DkXs
qFjvjTOximJIWhEvj7iVnZ8gxA7MEwCC06ANVDcj+KcTIrxIpWgAjKm0B0eGfAKw
AnOQ9f8sy+xW6nFBz1RdjkfFvQotHy4k14kF8AeTtg5QIRKPjZEiFWKmstphrkAF
8GAaNXDturO0+Qy8Skgv+dpLnRQ5Ezk+Mt4pQLdr9j8K5R4L+DTwt0kKAQAHPkLw
Y0ncHn9x0SOT2cIndr6TGgBV1/DZTZqTZeK52/Qr/tAdQ1L+r95pYWwIIr72tJFd
btyYJPQcz3qHFQ2dHJGp1pysEaJ+TsfzS7oMjSZEtfKl4S3+FBgOTJIgDkJhOE+z
Wlran4/EW8LytnRajw1LGChJE3k8ZHHl49MwgkewbYocGYVBtZTlXqUprOXDiThN
oZSGZE3ReIuiNZ2x0UKpHIJ5nfOcIFNqAinJnrNNBV3uJtJUxLn9zPLpCMoapHBX
SlLF2kjDTZWppJHczB5mEAMnmRewM8OOUxbs0+V4wf9PDE4LZ4DYKmHzEVATVtLR
Vf0WAeMrbGbMeKO5UJUI532WsyKW4US2Khf8m5L7KHeqrgXUCaVwSLtJw6hAvI4b
YCDlLlboJvbAapBCK+uq6R2f0bD7GGxO+zovjCC7tmnq1w9RWADku6NHqGR4VBD7
QpQ7xDE+/nLIUa2twHuKiMPZtDoZx2SWl0bhgk1J2GBG3O2zssCsJ1rvBDNKvCEg
tKbBevjmqKrnaMWtDq3VEms7O7+vUZrRtjtN8XtKUUvb+8ykPNxWnMeGGjM+sllA
yd9RzVCydtVMB3DSZ8J4xEMNtZi+QtC0vMF8x9P+UVanAEZYs9PKk1GDtyGjtown
MW6pv8AM4BbpaoWLh5weu1OgaOD1ws7jF69JU3fU2s3OJaDaGqaXbLlXrmuYL/GP
+YNbExrwE5MvCo3sh2L0YdovPSXejXECo/YvEXLJ+xL4ziUhmK98Kx1z3n6v0TAc
ex1YvGa0u3rEiViNYwFOwhiJQ7rXccUiYnu7UwatNMyBciKRCDD1NESkGhdczfDH
1McCGU16tkaMmnpSGdhlG+L/5J1oYD6Ohhw+Dj9tHynaXmOjuOpK/xPEaFcIvbtR
DliqxJiGWaPecmM7a10SQuB1ezdzsP7BNKbX33xUYfhZ1ALK6cxLWZzodd5KyoMI
4ikY4KniEaQjcuDh4khvXHAiJqTeGz67BrV16nGigefnLrcPmkpkNqqTVHqY/gSn
p8HWpIQFmIfINY5p/uUTc7l32XG5eKgfsOBUEUR9AR0Lk8bzjNVE9Sp3cGbSAexu
qG/7DXQp/eplDXju/9SJ4Cip4pm0hFUJycNcP6CfsmvzH0vdj3ClKSxVIm47Jyxr
vtLVaoOUdCxZJUjaswyU0mvPeLfdhK7Pl+nuEWbidTiJIUbFGp+yn1zVR+SfXb7Q
jr6S77/F9oMH86FSAD+zfqhYutryd1Qlq/ogUJuCd+MGs46fqufmcpnofB/FEEKs
2pfdKpVf14yFQfGcrp/IJtLR59I2R446LJY0q6efvNuaQ6Rn0oO1pNJj7rYiEzl1
o/f5vTgrb4aUqbi/dgzFVhesRS56w2iTEJnE658iUw9JVHaaORwA5KNjOn3dkeb8
QHe5nWWUzyflf5z49tNeGum/SjrafXqSxSAhzEnzNugkBtId/GscxAjUh7UXeLHj
pbDthJJvWd/QN2ueHWrVIvHT4CGr0Od7OrajJFTXVH+MbQtCeZfJANV7YB+bDrZh
8a1/k7r3XiwSLRFvoTD817cURhgNUawo8e42vwqfEVfi6S6CAqZdsK76TPGtNFgz
G2CG1Q3rGW+phsSiWT2i1bJRCr38I441s1GZHOFiwOjuXyjjleBncq27d+tt/7cv
pwMkpqNwpLoSVv4io0OpYizdNoBnModaeYayrM8qa1F5Sw+QJduS7eY0blQj9iHi
aNRNQASwwlvlNQGEsg9kxAShdEswrVbpvCSCQ3twsga0ZcFIzZO6GGnTqqSZCmqM
TdncM9h8syoXfP21K3KGxqt3eponMfqJVmCO0cnpvbbPLsnL6mlICCv3tph3rny/
KguFw5qLir3jtLTSx8Pcrc3dknXDDEMP0yQ0S6Suextm461Ee3+EQVYkkK1unFfM
uTd7+n0rOYocCeBzONR0VFO8WBYY4uUDxbW1CoFw+UXup1/TAw4d1W9zuPpN34h7
gOyhr7rFFguJUYYAdJSua5MAEEBuraK92xbVvDFbcBsLtOHRWV2GIcnfCoLXrJ5M
OMzxHJLQtqxMAXjYeal/gDW8zdFTXITirdEpnHG4gkTXENerHjUhS9EIJo7i2fFT
SJiVED1XdJDWWJDatIar6K+35XapY47q09y0rX7E8OmM1n6A83EAad2DKtnQi5Ur
/3sHBufSwPYbFsrIWY9gzu7/BYQSf37bWSpXnJBjh6r8muuVJVplcllLE27CQjQD
2dGEYs+IvsMEabSxon7Gl3yQfN1As7qcRbUEgjCHgxWIWuosaM8YUVnhqc9pTnUJ
+ciM2wcW6qBK2IPvZm/VR3UTdcs9H90H4wwIWm88fXzwtRqNzOhK0CCzVz/F2Vmk
vjio/XPdquphsODgEADkygswNquewHRnqRzn/3cqIliKpGNBFjtvO55vNcMHc3AT
lsbveMroQNhpzMpnOQkWXmEuwcokm6EwYD8aM1HF5hzWc22OhSUjnrOWEwyvgaHZ
TuISED6uJnD1dzYik7Y094rtEaxyQbv/FYoylbqDBxeraNUJdLtjDph1usIwcgbU
WsDY9zLtbjPGo5w1Yo0RQeLvCVWQ2VWKsuYzMZr8mhINVFKhWLAo2F7PAvma3LeY
ziIsUjNWsIpKLUeGzyUCOGFOKrBe9Zs7WikNyhvbA2w5HETjKn3AcWF4CvcJDBOM
mcCrR8Uf3MlPTbS5nCMjQ/Jq0KPjX41zbJWnH3Tj88BuO0NuEKaathkD5Xd/O0hN
L93QRXZsgxUwp6idsJbM24a9RT+N6HBFXXdwEmdLbfho1OzVOPvbuY4Dm9GQamMn
jGjExVnDpI+18A5WJiyZs+VtVuZc8ACTRBVeOelsmfUDjkjwan08TAtrR0qqxr11
sd38qRE4M6HiCircrK7IPOFCUGzeDUQuMgT4m0VDQe1T9qfP6iQCRJngJJQ0uzzc
p5mwCUCqxkqaItrOc+ovg3v4+L6WPoIUXYAhAQPrg0ddW+z4/V6LXkqnVMOGICfK
QYg8LgLZoyEi0oYEj3fFIx6L9zELROCnev2A4q5TTFrzVJA/7qkiaQgLUKMHWWdV
XvAuhYGNZ91hwnB3kFbMcoOgFRoCltCWr6rkn7HVmODgGf9F+ag7/rMkZcZEU6Qe
B9DYaaG9X1T72DxZjlPRqUl/8y4eQ7MQL7AQXP5jnWZ9AKEXplMGyQ5BDfE7QPJH
BNMLce6xVjEDhg48J6oJsSkggyr0FVMpEyXcJKydZQf2iYQ5PxzrcBKvAZhTkHl3
EKJ+Znv6VcnF3TLtYI25WEuFSyABvDamxa8JeLLOOyB3V7xqbXSDbU64CkFSLwzQ
hm6c8Htx13SLsggf8jjXyOFAtjwZsPwhMZXu/U7qtR86BHHGtkSaQU2nDqDWvgGm
GrtgsrzokhlYvDvX+GP/3yQGEL6EHo2oRxT3ZqLe8y/Ef0JT01Pn4SZWzREPgsi1
xB4C7oZ3puWQ+ZduwDFoxj/7EeDqbQQkwx22m2WCk06+xulPLMqaz0IA61ZR6xBw
w4cjmtWDwGj7sL8P7ZH9SBqizIFv2pV5EbKTXpRPvKguYWcMkBr90ZeRzKJzjtSZ
Cs/elagscxM21DicDIS3ybR5TRh9xIZnG0LpOenECNHodpVyRsXbiVNx+DZ3YQji
sFsr/uwbnEx64dKCG4BG3gkpL3slNE+bMSBsU83k/ddB6QQ0H3jND8PZxq82MT7f
XVyLv9ER91AoRw1f9vLz1/SK5LoHiIYstjJVKCA3Ij3RCViERsoTa5yGwJQ9ZNL9
Bl6N5BIAlPm2JUsYMPHtMMP/Qm9BKdUd1m9Pae6SoNAivyK0PxOiiNOwgavnOZ1U
4KMba2paY2ysaC4THVyZjTBciRF7gVYGOMlTnm45vx051HB+0stn+9TnGPfOSfgM
kMmGtgmQVsobgh1uezw6DruUif4ikxUOZJ7sIIvuszLTfxNdggtz6F2oDKf5K/oB
f7ezVK6zTI9CSKfWWzsMEJOP91GgPub5n1+vR4BbXTRbRFIkbqB3DxKlQUwm3mbV
x/2I3SmIKtKFcehMz3bMQAq8gQc/85jAPWTLm/IqPXwJmyMr0C+LUcS1x36wgSdg
VPhqCNLMzLq6/VuVPYqfab0JqfvwsHkF8KstHfkmK2SwiP1dv68Mupqfkzlzb1/V
NzdCMh3GwHp6qtCTteh7T6ju8/FGpDN4CIlMQEuwHTF+t6IHgvPGilJh+lNKrl2f
4oQBVO5fQDzQoXhkowPhd2CVuC3dQktKtaDlE3fKf5WDiWm/8RtOyIkQlYl/jNwY
tWxT1QJpheY6i5wGT/pf8Pz8fjvThMZcLlzlkZyrCAjgG8C5pP+O1m5AX22as2Pt
yH34bkAslTD7idZwhjpCmYRamB2CunM0l2ojK+ACIUQVpxlZTOAsyKGMhbBvBtJt
C9OaAb+SXC0BXCyCucuierLp+0JdF/BZ7GAmFYuBAxltJbzcFye6V1FFE4czdwgp
W1Xwh0iITiMfPuGMADpwtW7lILClFezhpygFa7dWajXAfphCakWUPvY1+Ib6jWwI
UiAqWjRyomjY9I5shuB8rGwxbagYEi2tw94ctzw1IXfTrq+prSPfOMqLiEHI8GyM
xwK8zrqKx43Zi+oqcPkmfuHqdIo2niVPRr1R+MtlPS5Q+NG1BcgauvA3oqwIJpDR
H7uRbh4LulmXwqs6ffpFs31FSn4PgqWeLGThGvasqtCIGwE9UapOMSm+jOUzrR0Z
C3iQnYnYKSigLllxkD9KR3sWeAm4rqE0elJp06EvQQJzdl8kCvKLCM/L+lCsE5d+
v6busqSVIlB8XuWjc3jhApmBO+eznFE/BLr5IpRSHGIHBl+NvE9GJmMsIMmWZzzu
Lvenwt18G4Sq2yANjBKeqBNtt7/x1R+zxIwVG9r3h44cyTDeCJIXoyKLEA4OEUzn
jVjX9xhzbaqURbAGdnxHYrIffeO32THf3D8WqKoy+nKlzqdWBpfjpT6RjLRTBQEo
54e4BC1b8t0dILYOgsl4LSQ8tzITJeWLRjdfwuIT2tgl4cRUQI4xd2J94z9PwCc6
KMoYD+zELSf4gH+sz7WB5j2ezbgTLwhRJEZ+TvvVNCmKRr7ZdOl0xOCwMcQ37DDI
RAS4f7m1dD1sNRgc91YNo3pwqfSPXpzRWQUshhqmilDJk7dZ++XdniT6e9X6O/Rq
J3daRduQlZocr07tVwC9F9ZsUB/+9Syhgrp3YtOWNga1IO52Lz54V8qa8sTLOkX9
VjyJnpOuoOFoBTtXMPJdMUeF+cbtiugV9LNb1vMnhiRUGJvEmxe5rQAmuQtPUdzC
C8RBFo6YE9Rsz7Saw1wuH/FLzraItuYkwysWKXFfdKnskvtOeW1n2DIIpy1b8JKO
wVb/4c0w9TPzH9SCZyl1JCBMNqnNvlxjCzKTuJ3D0vBxTU+qbvJdeoE+ioPxYCsh
NHFnnYYRoFPJGNNr7b0EOs2amUkJo16RutFhHJSxrhkdkHDzg2yGpDN6WdgwGaxI
PobBTr9BNn3UObJbtN0FF8Uajwesy8a1QEEB5zlm6MMzwEHVzJztyqO2jEg2dAUg
BGuitatabkSgmoHvxQsanReudZ//h/4tsxrGWc8VioorTOlpOMagQZqwmeSjIfX+
WKPHdn8XtTwE8Q75+zsLe3UeLyyMkvZH7w8BshH4eErVkcfKl469coT9krTdrKZK
LY5MtRTh8rS81YF8ZAhS1cOGbz0LAYwVsDNxAcSMMk8KicZNbp3pefbJTPAnYKBW
9qXGCrxaXZ20KHGf4u9uFV+ZVpIjataVaF8SqGl9M1qm3jX7r6PyeYPUFccpffLT
eEj5ys/6EhH+s8RJfqau2eSMotGeVgwEEcujoCvtlmMcOOvrixZTovxBfNxlKLtG
TG5JS6ElzOQVAcnqb7pe9b2mbcz6VirWa84q3gIFfxrCZ6cuGRHUwtDnxZB+kvOp
m13uMwjj3cjFSoHSytGG76/I9hv3zUNbZycccw+CtkFCeZmpIvdvLPZ5zmXDTVHW
lp2PRUrmlgbpoRrg8EIDW82S1qJN+hQxC1+IhuHLs1rmTpjk+XLT51OuzT/s1CaL
81GWqdKqNbM1g/qtsOSY7MBMs4yQ0X9Rykg82tWVEmEcb/dR1LlhDkKTTRzZFmip
58cDvUESMD32+FUrCbZmHCK5PckSvSvB9tDdBg3Cerj5NAIy8iuSXZfTHJ9K+IVa
Hsr8U7cH1lqqivreHaRZhqeXwmi+GkE0rP6OwVU2bcUdRA/Zq/EnlP3ASJ6ueRu+
alS2o6HUOcq0LPCOUtnWzKAAWgY8RwhOwFlaOAecLhtFKtU1uvKRF7QDSNnWY/69
+ihtH2vqrxNJPGWyuqAXtRXPbJRPXaUapZoP7AboZgvL7hHPTK2w0tJKTzH07XKU
Nk64h+TI9cImeXmLGEuKa/7OKCoKEK57lNGoRw+WDsL0QePRTcZAwvz7LA70atcE
WRPSdzrEKrYMF8TmGWZQayFtx14Vg31mZ5E2SdtwRwFVcteiT8ge+4EQve3TMgSP
OZyFbctn6HcWZsf17tfnaI4acLc/F8p8lQialkN8wGUGq1tR8ZPe6Vlho7zQAOuq
MefEEv7aoISxW/YYn6Rv2CVfm9Y/PHyP0QReSsFm5LGHJ2n88t1PjkRGM7gMtihV
o45UpbjUJ+gPRTgz8wpmfhMovkldp3I4XyAO1eJizo0/pEIO0pao8f+mO2jxlAgM
ZBI+4UDggGsATeF77fa0DQpURaH0fPwpS1AqshcKN29X3Okv0v0cSAYg6cad1K13
ni0IvQswQOlHlByuXnRk1g1RmdBhLrATjxtoaQBrmsFNyHW7XKzVtzYIeXa75BCj
xqvAyRgysWA1zTTEQygv7nukMV19WbdQZcijgsDPHxZrpN0NBOYZ7AalKzoOKoGo
FIdqYB64+jRE21qr4sINVdcBndMBxPYle9Tsg8qpsc3lbXQhpw4zaLwjipCv8L0C
6lAdgRU4iFw8TbiwYmAuW07TprKENHqxpuC7bC7DJCKC7haWp4OE9bgbgC3G1+2I
iXowmRbdBRMFnyXHyFMfUR8sjptIdt2+3mXnurSdCD+b0B9bkm5XLCI7E2n4UAwY
GBXqk0al1ELdQj6PNi9dUO/aQ9PZjmywK7flO6thzRrMzTIOE2Wgz3fCwaze2EU4
7Mt97uQucPKfSMPRYbTUdY0FvBxRlQ0i7vbgvFE+3T42mgRwhn0WdXIvhML5L9ey
cILYSghAQ5IbZHMjJmTNu7eYThCj4031nEcLKXLA14fxx7IyHW2ZuAmDjc1DlMss
2jG7DE+GyuTo5U/pXmfTuHVPCduKGjceQmC/IaD7b/34U46Urg3/14EGO3v3QloC
jucK9RO93EyhdIDGYpZM+UdZmBrtAZyG/ckItwnVdXU7R34TgCX1QQ2FjWmC3b4O
gQG2GUz4Pgd+ZsFkPvHfCGmCJniYw9qmOu7u7qTilkmtuQDn5qeax5rMprrcTUiT
ot0SqsXBurzFrW24z+GlAgXBUxjyJpWV+Phy9B3VNFrKKolebkdeNKwd5nONa/mr
NKVFY94Ux0N/dTV3GgQvqL7YYGlV2eelXLgw7C7ZwH+WjZy2nevx07YPkUiDwBxp
syT8jcw1KAbuz2xkJARvXNiQuXx40PdH9fpqIhDb1/caGP74R3xrJlZf5ZzqUPia
YqjMWJFOGyqpb9qhu2JAEOhfdiDIF+RY/BRy8GhFQ1qcSAWJItk4bIblLdwBO3ir
uLfjOOKe60775LMnBvFELPFU7CS8qm2qWXbGOG8DZakD8lyzy1eqraY4MwAPF9GH
y/CFxREBodIi4geiB0gqsAk1ica4R43b4/8rj4jadr0fFSxua1VRZIPgrvDCBOns
CFqYne/4HADfnSm4ZVoqsZHRv1Bdkggbum5YSeUYBIKg2EDiWfD77kJcCy+Kbyk2
ux01CUc4l49X+UED42jaqx3bcUsIJjtjAKAEZ6aCfjNgIlV8PV4goQWxXqs9uwGJ
iWEJ2317TD+j4UHleWDm51RnjWnShVX7hNVQ0PIILT7wXbMgieOwgLAsMuJ4VQz1
shWLv9SM/T3l6J5COHr378/BW5VAcYSJIH8rugYLdlLzRjnmthyis5PhJ9vBg11s
Ii0tP4h6QBHwT61AAwc+wyPWY22icgtyniKkcukKXXt+zyObMgUF+z7PtZTZVXSy
kcxt9/F8q/D4+9DYTtLQf+n11kXlKMKEqM53oPTGZGEHuWVSAXSyP2nJQX5aW342
ET6IgW8WH4JBZ8ohPprx+MRkMtHRFxhlCzpBE4lzWGwfDQwuzeWRoWe2H3E/6+G2
MaHNfq3hr4Tnbvy3JJcjl/BqBNA1C9IDtnNHANHWJxRFvaMeZgOHk9p/62NB13S3
VJZs22bR4jX6uVgPjABjJhQ52Kqehb2c+KIm+BWuBSaVwhCy42PCCBCOOK9PWEXV
1l7J3bgMZmXAHp/Eo9XiJeWFVJObEklgTv+Xnv3eXoQ9yv+9EyocQBwCTx+LVeAI
jQMu2RiVcZf7Rnb1eFBqVeQiwViMAS2EMgLNd5SEE4iqkOhuORXgVqzocRreJnza
OZ8XodlCwcKzDKcQUt22j4tZpGf8sXcED+ozFevI0O3VNaAGA0KKtsr9Doe1ku/A
0rX2hFRtkmyM/WV4ZcW04P8D65zBlLlEVl4aQ7cBXyoQgprGzExaeLiwSEnVIQt/
8lS28FwvWL0NSJJmv59/fU0AXY6l0t05Zwx3HIFcM1iUueS+3Cd3ps3MZUyesex8
X5uAEzkktAY1Xz+EtG1Ta9aY3pdxpUGyJ/cGpGRRDP6s6kCjg8aqM2R6E5Tti9np
sXBSlcWiGDR5K/E3BAcyciHVCCMrY82jGDI5KowtgSTOuUAJ1GpXncpGpx5duDzu
D/7cCJUb9neb/FXvUCDS68LCaFQuRAQ6ULnvmnltAtR45Dz4lxXHvtTqoClr13D5
dDn+crwMWcyZDi4/m5qGO+kc4cuMRxcw3ciwAil0DmYDMbfMTdXQzHYs8kZI2i92
KwDFJ/nJTZN/pWU4XPhZTJUKNRlKwbF//qL91Idjnh+GOJ2DilKL8kjj0QCm15eT
vMO43EksH5EQ6Eil8IrnAViMXAQaHmv0d/oTgP6Ui83uqICNlA3JvZnrPU427t61
56Gd1TCEZVISsxgLCkISyA8L/Wft1Dyq9/04UWMo11/vGn883rSdQgVUSXbRxa6f
jqP8xlk5ZS8Eu0fmO2/Bv6/Emc5qrEfk40FeKwZI+98C6mwMP6T1JADdr486ZLG5
PJlUEq52t/vzrf+x/fjYe0R7iXOcni/AQIobnQTk6fF1o9y9KwtaXtD4WQKbFNPJ
MKSzYgtYGtVyiHnVeGJv1wB43YLn2dazXhz4qtuRNdvf2E1HePuauuzfti4pVR6c
hdkPjasOi+q9RLfCWj9ndIKPG7zqY9x8LvmEzNSXKIhPwIbfCdzxqoJt+NJjFMe2
8vlIKXq4IdtGQ/pV32wiLL9TEYBE9h+tv/Ud8F7RafYw6A/1Zp8zI84qcicwtrbE
OLCRrbyXYbA8Y6oSJxb+vmlYdM+BNvFoTBJQLAuH4QQeXeCGt9xL3WrzWNfhRqTu
V3HmKyPxIHRg1YE1oJLoInJKfr3qRr5Tf+y5AGkZa+20/O0qAGFpg12O1WmPp/8G
nQRxtzuCFwU1NCZkZeVjH3EoW+783ZyaQDfI6n3+U1tSBKiRlucGrcFw+0fNpoFF
c4Ep9CM+wjlQBcKZYFR5bLWCF4Nh8OmbZqwVAckgI0XmVulZUh0XJLmy41SzdCZY
WXRuhxGXPEGvzntidOskd9rHBTifVSKeEtkiSy1DHld3/oemd7xFqY1xFxe8EYht
6pbc7HRKXNVvtnXTIXkIYqGq9YU27yMd9OpYS3eiMDQ3qxXi+Gn/izWI16ZmozpJ
FYzNzgtMBD2hGeyP1y3t7PPMdas/+dCnLR7aa8TaK5ehrZJHT4T4qyYEal0hUM+c
5qDRNJDEXhQkfe3QC0lVdaZulvwRShpRxBl1WoIRuqPEUWiSQwmrxFNaY8h73Xix
+I/z2r4I9eQcRfojvz7kkCpxwsWSkhphPOty6j3Tmd/mOA/KUlcfH+UPvZ/ddTad
TX8auM6FdJEgi3ePEAJVOZOlUJRajTgNNjyXfHf2nxUcw2f9wtfzCnB2UzIlWWbO
c+JBOwFShflfkGL3hwnb5nJIQpXUzSMSMvKSFueHjYjH11tmjSpv1Rurh+kFDwb7
1pGSRljrkY1i4XCXgFkiESZ/lnnFe9wKSEo4bPjvNa5P7mMFY4SiVpYqIpVJOuju
Kfohu6IW2nG/ge7jfMRSCmHID0pMvC3XRxw/e8KczFxNcxOFm7Hi3sGdKolDP9c/
TetCtggXw+NwThifc+IsvEdhBYNMSc0vgiEpo7bHuBloJOadLpcPZDIfAZNiaysj
CEbdYGlDVjMrjAlrdjRZtBtqhDte+WFmQCd0v02pGQCHpnQKk3n7/Mj90XJXiaaR
LUbYZrSO8q48Ni3UOBRTht01X71+F384leAhBa4GaMBYCcGvVeCyU1w8dwFppDSH
shSsWYFsKWPMBJ7eqwulKTBcVfCo7f0GOXgqOJAS71b2HswgDhijGGAVD6EU8ZwP
3tqmrSmD5BXj9lba3eokiccPZ1a1w61KfW2IfxcRPkSdPTY8D7uUUBuc6G+YCjoc
WtkLRFq2Qbawj9LKyCXhLJr1ng3J3Tjy1bod31x80PADgWJVblOzNfyYJhSfrffq
sTgPXHDRvfmQSEPXZ5KJki0GP9VqSZyZ1cLNoNzXjwkUFqdvvaqINk5YZtuczKdA
EUCEqPGQa3BoTmco1fcSeyAo1gCXClAaEYh89cH5XCREGc8ww2yOxknPT05H7VSY
rUhiIbEtlggxx+WIDYl2chpI/GlzmCGI4fX6CpN3QUwo6T2TY6qs1t7f+NqweHCL
SXZrC7z9fxw4HLvuuZw34gciKVzEO9CI3GYXwBFjCUtGAnrYez62lLkzaaONrcsT
a4K+e3yRlrHLb+Gs+7z8dKzpgDmI429EQZKFSM1emoc+P+PaAuk2N4w1ZNE9WFfS
RNfsxVHajmLw3ddey2mRdYUUAzSqto5ML73BMHIcx94nfIppfOecHtW0w2Ls50wk
L0RKJS38UN3TJvCDrg8OdctTpCGpJ2gsb1DD3tyhYchtg6cWCAGmZpu0ThAQvbyY
s6eXsDxhN3te6BS2yCFd+dZ5q0TngFhY551UiUzZodaawn3c/JZU7uFJi9h8lRGA
re0Fo6K7L+KEZyoKsszdddHw7kKkPZIc1Z2zpFgMQiQOq/5goFk6IqvatZhgAbyM
f8l6Vr+mroqhSEG62Eez2Px0doXW5daY0nZblJeaRE3cZfRJN/fN6NbOaYoQKfh0
mlwEE0WM5/ZZLjBdG9tqABae3KH/4EgIQfR4/nWxT4juLEetZYnZmX80c4Sjvru/
JXFe7Yvglrp8j+P6WVEy7bI/2IDEaR7acGkpa+Y/EmTpXi/ecJ7GiMCJW3LRzBH7
+gI7sCXGRaddPQqax64MvhuYNdt93edUD1cjOEVPUj1LVyOlcVAQupKltQqkGUeO
/3/nQAwV8T3aivuivrrNBpVv/ZoGQvKKrTXyQf1vo2A8v0je6MY4qKLSwkupxykn
s2f0okMmkmx01qaWW95zfgSBwxnhXng0G8ZGHrCpaDPgNdOjiZNujz2ZQTz6greL
CKhspSoTEo2ng9miT7O4OlR0pw16dCvRB6P6KwJ51rmrVN5PPsxCPueBQh7Is7PE
2RZNfhRls5+UM8fxuXn10DXHzy0Lfxd7dEahwWuNbKTeET4rQdT086ilbL+7OxOn
XovlFoS6I0/Jj/Rpis32hsmlQbcXneg6ElPCuwLqlYsHdAvs1uu2W13vb7ccrgfn
XOQZccI0/eCNFJL5apyYYCLQ5i9mzQ3MUG8S4Wcdnsi93RjehGGOf22bC6ceXwfW
3l96DYwBLV5jvZ8lOsp/8aMvUiUNVEGZKA7msqJjOD0TPC9LvxXdSzSwdKWg9buJ
5pvL3vZbMLguKMXLM0sNDSq08rD3yphUzC9OMX/l9Djk+AJAUTjf8mK1m1MxZfF5
Qp+xsurfWFeOb5q2/qoqaGe7uheOOCuJ9qU53ezx0EoVIQUO8ikwUlrq6VvunCTv
DQwt+0aL1vU4bBwA7cVvvn2bHoy4VJWhM8kTUiutmvzimzw/0YwG6P/LxGULppjJ
7R3atXbhKaoJXrobcJ0G1oFHf/yCpplsvoTGfiwiMfTN5rhrnjWurUlQ4xXybz3B
2h9j0goTiwOhtfa/Y5A5IfGmDW0I8pqjZAf6ORNhd6/wbIbj/QAFX+tPEn2pfaHm
4FsnMuNEF1dz2K1IBG7ryz0jDolK9R5dPzGuDT2dAuSNrPuILKbqr6+m4apOI+Ym
WHsST9kAxWEjbm2+PD6zVxlMA+TfI6GpSrR3EwAfs5C35l1rK5FSyhBIzJ32u6rH
A/UcXd9OC4rwWQ7jxjuIbOTZJnsho8iLgambg5VHtcIyj/lUYr1yQbEVj1UyzOD/
3PqTwP/RPJXYS91MjpFqxEpx/bTtK+ftCZpcp7X71EGL4as+xGW8yBNcF2gQ5wwR
p+ngvJQYD5lSaHlGz6AFJDzYfWlAR97ICKoyVGVsy4aaQMQU6Wo3t0jbPWJCcK6X
gIAWRk31JcpqFOzfrv0IunLXnaU739i1cqQ5ue6FCk1XEmit6jNtf0Ns+NmdwHWo
J/M1Mem0lSr0JHkXcH+8PxlObu097r1YAgRBbM4OfUlr74LLnx5mLPdoDvaVeEV5
J5sk9IvfkvcXGNXvpn9BnwyxDzG5Ko3mdoBichADaZWJ/FePL8Vcy/pbtgVT+DSo
FxOGDO558gszVEG2CBW8ZiBbEB9ujxgVkK7h6JKzb3Dyj3gB91Qy8zZ4tf/Lvn3q
YZAubHoHOA8URHqIBUCz18GZYfHkB4yCGSKIefu45luymegqyCoKclW124cT/AN+
nzJSy8Qvr1+ntlR9Lo2YqffaAgpna6myvZC3G50dkh6bQOukmyqCe0SFkraDRW02
VxkOakg/crmvQ0re2pqShaRq6v3jDnWMriModC9ba4Iqwt1t1tuBkZ+OU7u14TPz
pT9iPdrQFwe3Ozyx4DxefDld9YWxtPOchAJVinOSy7S4FmbzqwVQNZLZ9FOEVREd
f+p+R8FS69AShVahvd+lRY8nVE88zlsuyZKEH3ym9QcupWp4Ayp2u5rC2qit8+hH
DjGea4/NMPz2l38Zh9LlJ3EsNQ7j3nKaidH75vh6EiU6JJx1ZfcmLICw/hblxCt8
BugCUQOfVqut1PDr6TqtZkyGWke52nny0ioB76WqfwpuGLukn+1iZmXCRv3jJdAX
fbTLOJh2O7oxyjqH7oxAz68h5w8y9v08w66YpYDOLSwBghbehOKhq8IgNYF8N8zQ
SC9bb6faiEd0XYGh3diIEBAUzZQB/KAsPpxCGmGRzswyM4850iAAKUH16RlRExX8
nW8Dq4Mck3ukasII8UKXnHlZLiH2acmWZNrifYpp8wOCc2mb1jy3NBd5sxqwEERT
Gfw2LHVFi5lRVY+Cfa6ObcIYupmFV0/Sp29gc+30gET/t0aHHcSrUzZUtu8oGam6
m5ORtwSaOTgJq/0jn67b8LSqjpIwTwyaO2P+DNlDH1IFjY634qNkRSSOSg4GaNQh
QDsNXfzw7a02U3aoqHyMqoGT4g9keWIO7576p+LUvAgVL8QFZIRRWfez8sFlz04Y
fV99FlLwvUNPkpur2q0tOMAPLxx7EEaSdo2pQTQfN9xLIs7BsDIds788t3P5TRd5
bhyxrmA4f+CCXwgynOUy1wqlKYfyClZ0hxqfUys64ue+i+DkW+RecJFyqEyvTQjy
WTCYCaNnDOtD2ZoDmIt9wEmHdUPkXE7jqV249NtsTInnf9Clh3T4dGCW8QgTO3Ls
FQDADaGA5UliO5iXoue97kJvcZIPL2UYLE2jRzSBSzaEHj/mo1zFMnJVO02R5ePy
8yaumY2O1R0aXq0rlQivi/Q1Mp5g81IfP/rLNGubefFcNbst4k6kWt0t1zIj2VUG
jP1Yk1bzab8Cr04Q8kx7TlqdIzV+LulZCPu9piF7P53KuDw5nTqpt4PQks9/QMF9
GjtpDnJc2cVQprBBXU4UTwlvpAjzeuIKQ6BNj7O8c84lDAwRDypaPphbyFoDs3hw
/3Qan5147aLLR09llfMxnRCSko72xcJ/X+BYClGLqAgb1Wh+UlLXtVdbmFXENFaw
CDPZBPoW0nngO3ssuKyiL0MK2pS2+7t3J6cAGT9S6gkpqtnHeMcbQt9FDtFnsgZo
R1j2c7qRCSNEaouLxJYL7Dmzw8eIql7aPZHyKJ1vV2dO3FRzsjDkDDGcnlI4bC9R
MKxNk2KHcHcCpLi67l1gu/oaUgeTG9J0k0Hiu/B3ktACXNrRNfjDJRnFljRdOaYo
fb6O8A8ue39kCbc01MtwDvgejTDZwCauaUFJK/FG3EclCcDxjFmkoT5dDnyAOo54
qc4lsWitvnFwXSVr+bgzcoeG1UXllIIKW/63lXecNMeONdnNPnJJdW4YxFVqrRyj
wJXMAvX1MmcDt69P9HHt2AIkK3f6uTtNz0ne6aAxP4QYHOYsoAXJhQgZQjdNkd+i
is8dMGtYEwlcbj6TQSzN0g7hgE/BlUhpJZTGOPf/lg9Kr9D1fpOWUrungzB6vDtn
CVHeRMFSy0nCpz/p2JL9TwW/qKYcoR/rr/FwVAotx9Ec/YZfvwtRrl0td+Yjvteg
BNBaQaffjfICZHNDOnv2bHJvUL8UwcY8pRCEC6cAd5C9s8/oJv94JzVUUgRRtqIv
/+JcPssXApLIy2kIf8hPv0oDepy54SAle6mMbgEm0FBntEk1Y4ORRFSVPb/WFK3p
N7P8vA1nUPyrwYwk7kMLIfkPtDywpGQZsiHmVVhSS5HqzVR8m2Yb4t0Wspd/OP4M
J08rXeVt3GCtE3egZCxkIYw4UPEUWnSAJH8GKVw/iRwv4ezVsLqseNT9bKDBDdAS
AuHJU1fOLWCLNX6TemT9hFzqm5/j/8QvX4jFRFX6MqFhwdZadBAbNDNaPdhg2TaD
Qk9lCYoUvAXKQacW+JrRmPJODty8njA6j45OdnxYMwyhEoLDIh3SljFW3piaMCsc
j2Y2SaWasz5L4ngbpkfjBZHibE6Qer/bx33ZzmYfqXumJSZYeZ8o9ybm34U3dnWW
y9g1C5rIQ73Mwdf9iXC7qHl4x9u/lT1iBA4KXRxNKsZsNxofdM1DL2i9DaSKj88k
xcoL4vm1rgTAyo2e4xhAq6Vp1VvpXh0PZBrVAHAvE3IdzpL5ccArVnhpWOHAZmoH
eWbTcR6bo/2UYAkmeDvWaagWj4TXj4MoKOeHuFXcderglhX9T62GwszFIxq64rVc
sK34uoM7eq3uC/4r9zPuBZ4FpCji4qpyFF2WikgKmJujE6YAERHmn0QR1GVAn1eg
6i8Hj1blEIYQ0VlWud/afWSlSV8uXdcqbpAACpL3fWGwr+hyTx6ydQ3lZ6Lws7qv
Rs93yqakpWFTO02tHXOhj6CF66Sndn98k0VaxMmV79EsDABZ5EGpc74TSHiX4XoD
aZ9OBw8gTXvXkw2du170S+3HO/owH6bcmmy0RlhXyp1qfZKktMBgyDfOtCU9BInT
V97lHH5YUZksaaI9x/kBvvFRigRzjjl2TR/KkmoM3rnlBGeR1ivBLawDYFTHGClr
aOWbP2bARU5RLt+XwRKRQDIYLW8otpo/GofE6MUIdXnKsBXttF0YZuug/zUsDAwf
YuY7djBM2k8KJYIrCZvoPdpZ9NdExVbE1+PWSkEBLw3gx5MnAVcbaBudVQc3jHGZ
HvhAm9UnbwOjr5Zifglwbl9rwIpWCSoFoyt/8QMVTW2Ojo57E/r8ImRN2ICaW8XK
4Ba2JYj3gRiqtWroi4jjDv6iKoX1ggryAfS63Ud/RuXm7yrAW8BwkdPjKs8N0gbV
PRHKDixJ9fB/qEJ/p9Lt0WfVr24Cp9PRIr16g+zU/qpbd9KIdu0qTPGDVDhERXLm
5A5Qnes2Yl8J7CvcFN+v1xS1kTkxX2E9OEVC3NERQZDdAQMPhJA/XK65L1iYe3RE
CxWdz2F1RedhnHMt8LkUpYadhivf2jgrBgewamMydaobBJk+DcD6UB3V0GsXLGh6
lrDDa8lZ4QZaO+juDUYiGFSKYuwAsR5Aa+EY3Q2PthVYAobZO0swPeiCwn5+lYNW
x4glHIAXhFbxlgtgpghgI7k2svwCB+/23dGzmy3IrxKzw30doxAR8X+TC3c93Asd
4gH1n9eeBlNLUvlv7EE/fTgiJo90FjUvifdnF9J+ChgZVNcF+aAp0dSOPAwNPpNZ
Dy4tpR7jjIZG+YsBk+Ru/WEBluO7q5ZwOiOBf7dcvtWCSrniOL5pvQgeJZULOfPf
4bVSkfczvTrDuxJr3mZ54PxCVaHdH7jMLhIC3S/J9ur+ZFqkryUqmtEr4FbKr787
9Rs26FyM5WTmCWpSGaMA+onu4U7dbY2+VAXj2032mnYYUXDGfrqx1WY1b3iBUade
svR8P17iZYMFMq0pxqrKHR3wtutJZaOrXq4CfJ9HTZD/rKHjemipNm9vXTa/X5e1
BHNliLv3XcJsn/V6q51IwUTEfA79XRwXkADrCr1r9DEyWQkUHIk1bmz9BnyaHMgQ
35rS3XVGKPTT6i1G11TIBI8Bt9dhdhv0Gjy1FNwkHAHp4Q7DpovM340tMfDd1/FX
M9q5Glo3kxJwRhpXVBdrWoimGdZrfXm+VNaWip8jtHz1AqNYY4PuIAoStg5wrl+N
6EcJ4K+6fnCkpJzYm+AqIzBFG1w5SsaYCbJuaqvVmSo1C5DsJZkR2CRAkTS/uAmO
TtHuC2qeiYilALNyFCiJyoTsSRf3Xupsz08ejC6y7cC+AbeQbGqqTq7LEoI9f1FB
73LUEMT1NuyFJDGkjSO3Mtu93RW6+1aSB2tvpyPbjdmGSlWbkeM1olzJR0aUkLAB
tj0oj51wRD4dYgZPUsFwvETsN7ixuZ7N3YSPGmxhUWY3tUqJRmaY3TaJCgY6ZR6i
6AwW+isGLszbd2qeS/obtklVGTQKMEwyT1fsmthr532bcFO3/7jvLW9W2TJs9A94
MY+/AIEj9HoKoIoSkxTxFxmOs/8T2TjWQxojIMn8xOEDRruMCnFZSnUTuehRGemJ
m+DeMXvsBDHEReDLb5MgynymI3WJPG9/+Z5VtRW/4rljx/COJ7Qlqur6XoP/X11x
AJVVlDWIbxYURMyNSJhAqDzpM7OlKpZsFMbmy4NU1QqnkSLNm8bGqFcQAOfqZp9J
kW5FhJsBRt9zmZqK5NRWFnyM94AsxwhB1Q75sT+vy5VfQtRVPTVy9kuS4kffTDDO
DD3w3XNjeWbMZA8hpyrwF53Z54ahytH6DVyjBoFHTn8+FIwkFavqW/dZfPae29XL
nV8LO89ZG5JIPUziB7A+RahDOvxJpLqZEuoJkrqwMJmGxSytS/Jpyvg9GVYwaLL/
nMedimeOd2vlOg8OZREWqGFKPIVZkRcwAfy22WbvcWzN/hDFmBxh7GC18gB2UOYZ
oWoUs4LXMe4V4TVmJE7qyEuNEqrvikTh9L/KSI/Hsv2hePjCWeiebD2F3ENyaldT
czlaQMlTCALyfCUDB0p9iFJEFKw8M3fAwqg8cun6tH9/xMJZ3BL2IXh9K5d2KELr
FxQ04yZVW/x8hP9y3XEbklyZQycEjr9HbSJtWertqD95FbG7qkEPTz+5QJcTh0Gs
sLBlCRiRiE/H6teZpOeLQ9xZzWo0FwpH/BPSKSo7iXxdAcsIKpfKMvPBjJEFz2rw
VRp3MPSRkGE16e/op0ubyV+Sy7rvea3DKtNJq+n9MunBk8FkR8hJhEOc6oaCzSv1
Q/2zHYmgPrTGWNpUncLMNldsOC6zlSyx+0j8+HfSXnmgIrZW3OfBdG/2FTbF0aX2
5Y/yIsmx0hbotx5jZcVGrt+5FyOvnh5w3qi0fgJWWQQHYHrXUdTKgq940HFv8k1U
FHvm/RSwPTYbpUAidraWuIddexFCEaaOEUNzbBZy9y8BXt52h7JKhEj9lEdYPCqu
IUlFSvym5axr2fbDd4Cmm8N+z9NkRlnOwjFGT7NCXGBiegoiHumzMQpkAv5mAtuT
xn7tkMGU9aJX4iZpkct9DdPhauPWidUe5KJ8YJ/D186xDie2APC1jmveDRC7Th7+
V2AMGWSiwLGXVc+1e+e/llMjQzjSkiPftrt3ET30Fj8FaDmprpJC/Odtt2VDNr32
8MGp8kl9LxTG9gcgwNb/HZ4yDRnu3U1RrGR4L3gxaiNzWxde9LsqmfleIEtfMs65
eOAqljgTwC+TQGtmYyRFr06EcZFJ3LGWa06Axrv4PId4ldueNjQ0K+DvDVBsYk60
3329d1Tqt80mAXasnFxvgFz1Q3DGgTX7vQhSIPgxoQlHUCQZGcXMaJjH2YleiWb+
WSvPX6SK/nQfDUU0bKxuZhLzv1TKaTaXNkTgES7qzuAOZhbwWHkEYKJkJ0D/xngY
DFXFtsQi8IiKoehOKCDOIRjh034LgbNs2Ew7FFDT/ipohZzNbTcfdJTM30iz/Fwl
sJygPuvbZturEzlKP0OX7pBtMmAZns/XBZfqIH7IimBjqS+u2Cvphpk5yAKTTtlM
hnTDIldlMPKcSHsAZwjOyIqpkPvp9AyZERyWwI+TCrpiz2CPlOLLgqql6WtF+Bq8
Sq1nO8cVENQ0RxSKbpiTca7TVSkIPlVst66GpS9aH+OrwKpjqj7bmI1dF6Rm8TWo
aXvRY1lu1jmf1NnbVZAY9ZxRnyOQK35fd7DWXJj8d5ukPRvvQzVFZam8A5H4HIxe
gSCOoq4U1NCBsHI15+6h+qfcwklaHN+W6pCf+Ccnx2y7uNUGGqfP+e9QfI/9PR1D
jSGgGrMySK33Jxh8eICYQJ/yJ2bWzIsEAnv4FQImv/QaUpsxUuIUeZmvkTFLExYp
Ds0iu6LbGgvA7WWtYR8Vb5HIQvI44cCuUTd5qftW92VaA5GcpabQ43tis/iAlkJI
4etLDvWFCg7JKl4CFj5eh2yAnoUO9+SU1rnXeKsRi4G2d/CkaIcuL/yfpkUY1DUT
bADEP+4aQk0FYD2Eq6ZP4TnfHXL+4HgfgVX7KzApTSgeir/TIjydcvq9GPBXG4PJ
byuso8zOcPU5rZKO6gK6nj8Y/d4icXaELEmiU0zLwMIwvrnP1TPl1DpLQNBmfZMo
rOlvCYWMMJpCSwwutWWlixpENfCTHcdmThbvnPsxBsPrL9w2avrNyOrVIxCH/to3
5oi0vG+DkGziIWiCpLsPk3zTEwI0tkhLYZTzOTh9NymqJONpNpXXZ5swdI7CfXLw
cBU2X7MKWEiCdxHzRNncxKcf/V09JZE820t1zfzzidb99DQ3+pJPiQ5gwFG3lNoz
o2c/ZMfakCxh5pfYBUzr86xinhxFggibL/QNKVipIMvTPnNywiiwE3PJR9sIh+ef
lWwCbJGPGfoTnNHYRrge7YUc47E1Q3cxOP40d3Ij2GbGG+a3DXMiHtD2HoIl/Be3
od9ZuNFW9UZ23uO1hxQEC/9Y8DZD+2kDAEE/TIHzbUXe3T5S5JIVhHzWi+nMAWbH
MRljzNfBuEWcmBBzbjuwc1s/fM+jDwl8vnicbhS83br7wG0Nys9yl80i409AqDr+
NGzfIT1UgbTBBDE2n2TkEDZ+NjrOL9PywAapEBfh4qiOixqNfHCXGDBjxp/E5C8k
98N1Sx3y9ReuYpiDczKfChtM7Yu87bZRJQvmF2LeCgbofZkpbQLYcgb0fo62tqKf
wMiq1pZx15K6Ct5mfY5cE0J3xVADjumXSWcGwvCuTrZAUBbzF/Ms6PK/+NT6VoMD
JpBlPLJFDC5eBUuozGQtQs/FGqo4+cHmEsJoidDfR5thyZ2JNxOi8L10keY5ViJF
9pP++2f4KdgJqRfwPdctjUAvjZ4VaOlu9SL3KBIu7EnZxFPfK9s5uM2SDZgGKEu9
Zb+73GH0HlmyBB/16HrQsmrRh9Qg8E0ymYShfFvO+MHPyM3tv1V+ttVwmfYZNrw+
CDDZknRDeKwF+Qr5gtj8cTvjsoQTTtksgxtl/eLHvlewtXON7HWmGoC3PZMjfA5y
ydDmbXrewadJBqR93CEGYB/pXFAZX+hdBIubiL4VM/0f5/o1No0xNHlBXgqs0RfN
HDOPvLj3kvBjNb5P8Fbmz47CnZVk15b1II12b5nGDxqUGcMsdvp8lBsSwWkbqzkK
E3w+b8epHq4lakfD9kYpjjyTvAWUGL2pDYXaWjxaHRzB6E40LXvtGBEeSH2UycOq
n6ijPeEH/17Fdc4Uq15L8sTJPr9u74ewHINd566jq+lm1N3EeZ1q5N8dgkoHU7IA
pb9WH+gqODwFrLUYM6FZ/kxajbiazbPaKaCXvCW6WeUWEERk7MdI40D9eMazXDAv
v9L0DP6KiMAziXVXS5mMVMjI7v7xKKud7f/9VidLMazhzNArZxP27vc/cK6tPvdF
ok9yNQHnUiVOuzF8S+A+7P582AQDhfuJS64CV/s+ncsPH3RSzWz5w+XR4l8bzxMZ
h3NVZ4NODl6TWYKf4ChSBun6UJkBXIAegvg21gzRTxBgQ38yAJ4OGhzshr4nDaiN
qTojp45LZDv2rDzgVOXOHwD2Iv7Ab43aQevXNbSe8VHWNKW3ffuI7qIue4VxBPfj
yWxOhGus7uNxbN35q54D7aIG73YW2X59XmfgTCzjrt/1Ag7MlqAGNTR1iECOuuVz
nvftE1zFJT9529LKr9jIGiON2at0ZclPL4ncswhitQL71SAZ7sGQQgJ72f5W5mcC
1TzEXTqxNL29NTrK9Z+Ejzkr+Hn0fMA+c84MI0tBkQfF34cadLlQZusDzuPMyL1E
OSLEGDAwoM/bVgqhg4fAztPsUjSkcgA2qbxcm9dVeXzJou5froCSMAkM1QGwKhzV
daeqz9P+lBAesAnhRmJjqJpjVNoFW71krLhKI+fjCEc1xSOCYHA0G6f8u1O1SLXo
c4ya+YcPqY/7VgHKaxxZVFCwmBdLVW8+uv/MrDjBOmkM0TFGOASD4LYlOs7ZGH/P
6Y6TbRKcOjzFlYQqQTpf/UMVlxbcYbZ3WMfemYIK/ixShjrMscZthH0WFGd3imkx
NK+k+wSFoiZnGGKjBjS01Dp6zAIQmomrDLbuduUB45mw5v5qg7UgihpzoEm/BU+q
KNLtt13K26uQ6XaA6OHpqLqMz+QeyFmW1kmnDRRMGB1NccYPQmFU7vlnN3gtT+jA
2Jf/KpUB+r+ALbj+4z7VCyUZqtg/hvqhZrmG/L+SUpLyMnduyGxQaud4v/9NXT4n
GxLoU56ROF5CCYFf5rnkY96Aalx2a2ST01zPTSpzmFos9saqciOroIuYJdGWRjlX
FvpPioy7FjGgyDa1tch7B96h5za8YxlsrWhCKvNOPHDyS5nFINWli8APzeuZAoi6
CgNldYikaDGgEC+f4AsZQgEQ8gzJ+f3O1CmZr7bsTQ3IQ49P9zyXEH99IvHRYTDd
b1XBEWOuPs9GsDcM/OXjpVII7M0qG5sq1uMT4+Ea0v5ac5oHiROhiJLCaW8kePuK
/nsaLCe4ugXheaxFipbbWIOQCss5wlagMzVJDj2ZSjWn0obrbOyiRMU+AfOpUp1h
QFVmgEjen0Q3SeeYiVuWLiigYGwDsIr7obvm9RtIhUYDZ6Oq7puVgcRkHp7tvSnT
TGS7BH2H8cFg2YTiyqgOa+UzMY+zD05FAMvISiuLXp3Hrr6miG8EzttGjDrEAmxU
e8QCnqql8I84a4VTDGY+h3j9v7wNwTqa9FiEzHSAEKgdkoTD4avPVS1bXkAo6tTL
fuEqzVIyWG4tunV8X7g6suaU8LAhwm6NhRPZ64cVuDcVHeqWfbs3DlhdHR4pRe6Q
n0w+VK+R62POlf+iUWw+LFYSKj47cxxm4rB5n5vGftpEUim80voNquNMGv4WbnnE
sjGKEBZ+kvMDqi3+mwcND+HEPaYvLeV9JXlAMheOY0vsaWD1hS/PGCOtoQ0A8dsX
VQ1c4mSDsRb2fFxJZNjcoEweD8DTCsM2ejbOODpVmAco28dvTXHYpHeL5hOxFePY
wg1ZZRQgQKv5Rs6PrdJczyFY4+mTxucbupsnSROnoq8N87tzx9iCV5tTNnSu1Xrh
5FkD0uXDlDM4nR2sIUuNxiiRjR2gc5xeAYSv7qQYC4HiaCMn/wmc+ucTdou51ryi
WK2OX506UCOiyMQKuCSQ6GyONso283zsmtwuZeY/qMHdqv2MUg62DCNHCama1UgB
Dp2+QTAXSAitAxf25OLRFH0e2xgiNS182ucUOoLkU5EDp2VO+F2TTM8Y+J2abK3E
TEc6PIwkCPn/S+XHOnuroXBok7en1521OA0xC8N3PbWy+0zJ9sRFwMujyILrCD8K
oAS8W+gXPtT+ibOV+JPDxr+yhNv0dd7oOYVeeICSBKmhEji/a/22xL7QWRWORUp4
YGeiVWUhaTyFTZJG1pSW+K+HdxBqC9TkANdSzbH0CYLpc41R02ydgDuhaK60ENdd
aQzu/5nzK3Gq4xRjMym1rMpCXKwCJiUsTakFYfhiJumC3LRGkYzyyJvgsKO4umr4
TrE/52N1GTqbWSi0gdSyGOWgHncNWJKM5Rt+qkrMGcrvXNeLvgcObvvOwPOya8zc
A5YNPjFtbEQE+KbIgR5mZ9lS7D3LP80+Flkzvbx/YFEg2ogSpFoJP1mO5lklrx2H
Q09X70/wU013xlWekEzd0sAbowDrbyob946AtBmH7myUCbTZScU3ZJ/t27e3EZFs
wzSKMfz6Z0u2L8ZJBAw4ek1CHEgLQaluVwgRQm4Ez+ePvJugjmusbBvq3jcLD9+M
/G5/IhnXZVHAGWT7oNkigeUU+VRGZSSrFzOlRnYhc0si4Ou4uoUbOhR56PxM7raD
6xBxTfwflewiycobwcDuLJF+87zfAUAKO+N3dfe88wUwz1Q9WsfT3m2d/cNjpb15
GL+RwAc8HyCCe+sYTTdg4Yq5prL/jxROwxfda7qug1q44m3dLbqOCrYN47WgxdU3
y8UuJa8K3PBVfdVc2gLDDl3Bc8Zyp0CO7K9ct/IREtoPCc0gLbBIeC8t3izEDMsH
9f09W6XRnUEYPif39aGvS2AgkNNiZyhzY/PEGgjRd8IZBaWcbhXG1XvvLq20nEyj
BewHJDgKah/gK0OulPtEJPFq+XK8K170omvfJ8tK7z/v/ZPxzj+w41Lkqi/5xnaK
rfJqmbNwStmRQrfQvo/UsCw5rTrq0qhJQnfUbs0EZL4DXz90w1GBWWI1r6UyqR3g
rVXe9s9tYhS36PFKU0ll4OTXbgyDgnLZRhKPtO+2wU71aCfq1ibR1x+LjJT9P9xX
HieYbD5ERJiDGnG0bHIumooQN6zdQ2FWxtPC97mp6vEA3j02oDS6CwJMQ88zNPwy
eHeC15al2EOyzzpZFMCuiwchWAF5lhtsd7BhNyywCqH0BaD6BpM4Q27IMok3kjKA
N2Utzo/DQVtOUX5XUzWp/Ux/CMK2UtLA2hqD4Q107bIPKgi389Dg3P5kMnC4NbFa
TAd0Fcb9lpkgIzjUtf1fS12B5xl49c9+zJXumBZccKwHZj+yTVJLv+JB/0psU3U6
hXTaX9lkP2NWPSIK3rksfkcsDB5kD0+SkNSgLc3akdQKDd1NXbKP03R8rZgSVCva
0JRhbiZgERMHZh/SBQj0zp46Y6HFpjOSYhE5PzwaZJ8kwl16MU+8R1qKR8nZGQbX
oulpc14U00i7jFkps+v4LeC7ajyz+LQGf8NMNTJuWpfWPtmuhXVpJcQTV/kT+CTS
n1f/8la84msfwvmKjNbzbhM82xW6B7ahhFhPe0tV3C3JEgBDPURlWOOf4K4S0pVh
uW/BfgtzUmEKlvzTXudgPPKHQSQAQxEzrhb/MECFqNR0c3hpoB7GVa6gsMdK1wCX
ZkrdHJ/cSwmV4ubqMjnCGMqH1fAC67yrFEA0dbJQTA60m4wGQ+sUxne94UR3LI6z
vBpPxsvkIJJ3dpdf7kMrRBI9s4diVIYgSY41mk+YO4lstd32j+jjrvR57rUomkj0
OkW+lKudAvGaRRrwzgPQaARQYDC6d+Ch+zd+XivUfs327uWUxHaXR83HyWFjzEVZ
YroHsLKVD2gz0+ZVHPhf1RK6yLF4rGXboCgfUMrOS1I0JSXmdF36fAcpbn/4Eiqp
Ay/3XmqfxkDTWwGvw7BbRRJhtTeUFWnYyQNvKPwDRvKj9oV3iPDZoGlP8t0fXiDL
POxagZrTz+uHSTB2LevsrYcOR6T09fEtQ/B6EgOIX/176gp9AJE3t8bHoA8OGUY2
1UpDbIom2lxVkmJbw1ajekLUNXDZHptWFCGbEVNSmgMVdLPB2G/1gadPrwKx9TaT
r5b6F3rSD4PlF2gRm1R6dS82ajWDaBohy8wdQjKagDJ/y4LMivBlgxdcmnFzPs7N
HeXIFT0ivY4V+jCsRloLqwALVrSIdbBNz83/NQDz9q17H26hsdA1R7BefRdm/Hua
I5ayywpZCeSsEMa41T3PoX8MpI/i5UbL1K5f7yPf39ExVXaVltMBuMUdLnZbD1Iw
3S+WS6WU+T2JekhiHJTsf8Lvf0hIPsgTDmYzehkgOqqxc75WZAyzh4QrtlrMyKnu
zqnSHJmrC+KG6cI3FEPNf5Z0TR9eeaLeB07233qsuX08hpayrTa8s4J9PtJCVyXu
7MCMnCboRWzGDHLfFkqMEUKf/pxwn3Ikd4Hu5nYb6tc2/PfYy42Gdx9cp65tusNQ
46Ytn3rnlrKRItZoJ6tojwJwqIaBOxAlbxejyyrJTyTky1bl4GSomoctPy4+9enV
eIk3OfGFcYkPViG7tBKR4FCo/iiFvPY43tIWiEmFonGZ3yzLHNAEvhaMZmkMjDZd
uPsjPIWWTyRWSXpPZnDCIl5AkU3kyoeNJ097+HHOHA/j3aI+tTGmjJWKdZd1ig30
IfBI1hE0SRdR2BDoWIumHJypS2R+CpJ06bB5Xkbv0M36rL6FH4R7DVwJMR2P4cV5
ZWr3qSRxlDJ1rRbzXP1wNttNosyg8m5cDyX5A/nqCzD61MMlv5+jNIg+hITYR+6L
ZR0Snmamj+ofxfaQm7s4awdbV+syvI69Z0mxtYnFHQ3XlJ+4LWOpjhA3Sum9SvK5
60/2AOEvqJc304iPGgGenFsxkcfaQ1E9kngrKSNWvP6F4VnD6L+an0wUUAgaHSDJ
Q6+wTw/9X52Ht8amWRX1vEAr0XA1wOqvsf+qtX9Eq08HbCWVompzF29Q92G2I0cp
BbNI6yRoN4gpK6JPzzrhBn5mycmt4+nDVYvCm0v0CJ/HNuyTMZyuV6QBoCsQtyL3
nMCuQBMuEyzrCGxbwh7hrQ+uaCGHyI1FSHg9cOABI8Dk7GkKR2IKKZnMd9N9ilRB
wSu25lzZpnL9BZuOrQAYBCA2t2Wqmmvs/oWackgb4btilWUulMg/MZAwhmi4oPPM
6B7kp7YYTwdJwiPJuXVHcrrr3vtxLMkp2ZAJiUAJoMei59byctOdgjV0l2DipPp8
c1mdec5s9Vj5cNCFRrnmW0oNsZguSN/NOpigAuww1BwHKA8xzea+cm7q9bhhRzid
FuWmM+4sikS5ApbN//RfTuf2flIrncdU8uhZXL2WeSt+ShH41cJ9fwyvzSFh69R7
DrHhoIR63LyMMcHNvIrx8RYvtXdCyAOhUp2GV3BkIH8jVz+0kaod8fsZxUYL0Eg+
FUA3fcMYIZdyuJo7qIva55JgfDgebKZ7yZUagBLIkrLbaAMZBJK5T6xkRHRktuiT
WoFVW84WXNu4pNFTR6bHyxogNFd7HMBw2JFXqDaKfmhoEE/xNsb8DKtXnuXprv7S
lanU5J1qNYQNlCzaMvyv9rXJma8FRM2E0xYU0G2BgAsHAeQv/WJa3ULdmE7ivBYk
tO4I3QWhCppPv63IURxsHwXwVV8xhYiT3ng1243wz3Q2syu8N60DlfCTWcIj9m9E
b43mm4Ka+fKyFbcsGN+GDjqkQKFtJGCre1689+z7HUbdPy1kHW0NiSqxR+G+CJ/2
AUvcFNPSLBGIgE0U9l4pmEtG30Qp1xhpJ+m2hlcmbPU65bVT1+b9tMPlkfjiZG1i
HoCknMD2KW6j+AiTzrdb/dNrvel8nOxwLtMxXu9A84L1OSNpVA7ag7zelGUg6tTt
6R2DOoq0F5xs3NjXZE5sq8VAz9SmG3AAeItjCOHvnUKYtF2D/zDOt7bYb4ObDmFO
aKcVW5+nwnMR62qwmyf7s459cVnzicA6TYCmtcXGu7BycUn+CeU4DzWYUhACRTdX
1qmak5CQ7wJgu+05i6QmV48+8d5wDVxXtM/oqDUxI2HBv1fY+a5vxH3mzTIVV4vG
LsN5OoQx7MsHOwtDkKZNuEgKkT4GE3/u1/MrAxw/Ril6aVJMp7cnGUMCOJLpU6es
f5Jae0xORgl9RyBiqXIJapm0ktfTxFcmYAHybFQxhpWuWBqsyRd6u3fWosTMaCMv
YPlsZF8QwZxv96htGI391uHKQQDyCfg7CbXNKcIm0OzbxTowOpdY379/wWzz/uG0
wHtPJs511+2jMhde/QogMQqIqMJA0tGBKJNVq/5ea/kYyY5B7U27avDw9ABCbxlg
mU9idDq92Mat9KjTuPu1RE3VNi1x8yaY6kuOrjwUpWoQWFelHNrazGAL8ixI9N2t
GIMGtzsMD+Ab8d5EJG4+yFnhp78Xh4hG0/JUDYBkmZ+LqUXmKqGV38w+NkCX2iX/
gxaQYtLNslBkFlCyO/+IJhUhymBpLjo+93cnzNVQ5kivPjQ+OMaF/Vm6nF89MpSC
/uBjT8kklZG0Vvb4cvOcl8wOyEqwl2e/aNW2R6u1514JTRTvxZf6LBCnVpX6CG7r
yZI1SScD+vzXS93b9lS/iSId5VICTWZR/N+a81CljY9dD77YekKTt04HSHn5IBrF
UHEMeIFJedstBdHQMBzpYMxFzyt84l2zYWe0eto+pC8x+F+T/rqza0L7PM1pvVHG
MBxxqKfb6Sk9n+85cQvu+H96F27YdFj1aBSZPaX2gKRjyFzXzBwuD/TQ5iDVQ0Df
ZntUTl5TRaDogytrLFlNUGoIv7WTSZ/FeQ/I2zw7H8nKgJYfXY7KsFRWPWO8ulOD
J+xwShu9TNaNnOiyo1esHjsYtYRTJ5ThMVsld0pUhBE5bpWbmDR5vRcmsuqSMxnz
k9UuUciRe2wojgS+ON7H+504M2XIrxF7obDqR2rbg/FANXdSL76sVZ5ee8+Pk1bP
vAEATNETUFMx2XlpRxF51rsNcnAddMbJCgbty/N5tMKQm/k1xiva540GrT8XCTmF
96B5ypu9c5iU4nr8cp9HGjxyMf93gHDS9XEYg1MUHgRUivpUMo6hy/qEXxO9o8DA
4l/KuAZLRz0rRTDgAiQVBiIeemvAdlV6iGo4XVnd4HBqqI0lh21B54mjhr6wzBnr
bCRQHHY8/q6oFqtqHuCKZ8+UkFSodwgjTqveT7InEo7BpB6axrpjTubFAk1qOJky
QCfkfiuYufOuGOgJgEl6przVZ086N3Oew65E4YWkQlLbd0tnz3aq9yWxxe9fmOnr
Jtj9irMjyJRttJNEsRDSi5XtQXGjv0z4yTO7eGTgJPn2v0LnIZPo44BPdEPDlG1n
e+DboXzRvNADF6OlaTZR6ya6uxAtWBetL1EsrfhGRyQ6nqOqDT6A3WFtDNCHKEsk
VOXHKG2ld3n9LslR6JRhgROJIjvUDcbPq5pCmA6n7gq/lBE1iOflHNTaZQLFzci9
ko01qBEfEmEi3vxtqjzv/dlx/kdthq6AZoW8D6fQMgetstKe4zsRRgP/xBHdvc1K
V3CVV17HxlmCDP4gJp78Dsk3UKZo+9zcekNrDhFScaG7lFI1Y+Dx7X3WwJFHBqau
Kts8wV82WZgsc21d8IshiQuAS7b5vuRe71euBaMdIN5TMnNYfBGvKnL2l0rsDSGh
QbdhT0lndGhCsV2hVC5Xk1ZZnNnTMKpJ7T2DAmUwmg00fobmi87Els8z9SM6p1dU
c/LtS56auVGnePAIGgaw8vl2vdhaLI7SUjX5IDiZ8McKrT4Y5iF0dg9WV16H5kAm
Cv8rhhpvfpUHVQugNwWpu9++kjUoQroXjJXDMnQcbwUREK4QQJN4Vc7Nr/HSvCmv
ZByBEFkfTxAg3myGjlKvgY1dG1g+KYONIpFxzSr3sNYAQJMEyr2DO3WiXPjufvPE
Go03iuTETKKorArNWyzQu8/a2xXEb+YABLaZWVoTEUilL6TyMUitptea42NJQYCU
uM31nrR4+cFK+DC3PMA3KL1SY42fKscW37oD9OLWefCYLXF1oprhpiMEUHK610kW
dkjYJa2tDqUPWBQJ9HboG32owMSeF5J3hydRigKjsrOOeeE9AKgiWg1aBmd18Uwr
sFC0jQfpDAOa+2DJvzTAd91rugmVlxa2QDTr26ypUnSLb0DldM2KvSwbDzSSkQ63
LGU1TAagE+6OOc9tdTMeebtZk6X8WNJF7TqTDjV5+BbBtf75wkQvEj9Iw2Nzz2EN
KU1RST0SgNxKDA4f0KZi7VOEr2FoJHnLba0zuK/UP2tALXlKc3HsmjOFZtZSUBvh
JAG1RTu0dGhwYwjRiQ5JoraYawXl5uXrDXIiRlIBy08HZvw6e58Lo27L3dJoUs1i
JQAqAeUa/YyPli6OvIw0LjNK0HS61EBuR4ttHKZv4ytbncSAupKAwBz7Zw9NF2/x
tgLEbYBrL65znGmqOypzOAwCwg7tLmNvZjKv5iKX/aRU5Y1hrjMpOLAYY03Herdz
Cev3V6Y2CTxDiwbDPgDAMBgdMCAbbPAya7Qb9/uH2C8qFPjUKOYwnE7AKZNBKwz1
XR7o24H1l8u+sgQs1acPY0DWbk/+XrWL/Vd/ciiLkPlhuSQk8k6R40Ci92STKiZj
BLT3JdAqBQafbQ/QqkMfe18zb/NSl7CjdENdmezBhUX07SZC4KJSa/3t7tkDZGc2
lVLowlM6W/NZFj+iitpndlCViikmJDanOfhm2+9x895AmZQ8tMG2i03X9dc5tKaL
7ah3iZv2XNOq1IHW5vAyYGQskPxpxMepu2uzE3REH8+GxgRHUVSl8uUthLQgf3cg
0yY0PSHw80IGXgsDHZVHaocV/9JTknmoSk2fLXlh98Ket0FUpSJPXXUVbF7EaYLK
1xb5Kb7RfG49J+OJ3hiyOhJXDxJ0QWCuLmC/eHJslFlwT7J8qHE3YEmUc9oKtWhf
iLDcuddgsmlBD17puDDinq3DS+Ik1KqdbQ0VtlJ6Klk7vt/dR4fkbgyWZdijsrKf
MLrtlwL2WkdpeDxPTHkLgxiJlanjqaKagKENET0dtMdCsRQPYTgBCDZU34SaxD4E
7AfAyC24TLzu9qYnsdHchoUdHlCmlBqoq6TGRooTYjSMqCbHz9vhDBsyeK/HG0vK
GCMiu+S880Matmbae7ST9AfciOPBpjvX2nWhk+EvXBb49+0Vhv6bFpdygEIIm3Cz
xGKsJnjUxh7dEQdXvRVhSQwDXMjLsPMMRPqD000q6H38ZsbiE7MTGHVBS7tL6pIX
210G6Ae5vUFsM1Dti5OmvQHkgBCgmXqIP9XezRNyCzs9xemVz2FBsFpxL7Fe8JFI
qEk4yH8kJtVHyo6DeFuP2aptca4ch7dN08rrKV7Z8QrHD/oKc4F1um2nw/jYVPqy
gIMmhoiTIBrOPcMpKUUBOWl835l0x+tYyBhp1Azb12AxZcqbFVbPLqdojthcSjoH
K58bql3FI8oUju5OLo077YTFG+NskwbRH2R5Bi592q1LDHu1QRi+jbbY0YYIN+Zx
KvYsrlgutoGVUzpfbpaHQIQeEHKoM3UvW+Ik3PULxa064t39Qj7iLLSlHa1q9CmC
F4VJsbl5hlS2qDw7Xys3Ofuwkt6xYtoIHMRtgJHvnvehXcI0ban/xk7OQ5RWj5uq
3uy1g7SaOijhfyoNaxSsvu/Sg9uAO49gB4DUT3bQaKsO5kPIcH2wQf7qmbWgqSFd
CvkLnrGc1J8PomD1+wlxVEIf4JKOCxsQ7Bx2dZxeOIuvuKyYVgm4BR9UH7OhqG1p
/Jx1F8MhHtQn1cHuXgdDNfUs81m9oPv0gorIjZiLzHzSRvztFZUMFYd4tciWhD86
b5djzpESBnzE2ZlpDZCdv872B5DdP55uZImlIUxOD5968q6gC68ixfSzfVZE8AgI
TC5JDCrvrN5QnmydhQziz7vQRdB5NaGxpJtZrvo8MWPqUaM7aaW2Ui203/bu3lyF
DQhDsLrZXKQJt2uNcpt5Lf+JRe3utPLJ9qdPtUlEqQCTfsP0UJdF1y/JDXGKJgv9
nwmwXah4fQ45DTFOoYE79nEOdFm/ZkQZE7/7lMYNcJ9D0g6WhYnNUmJSItliIGhI
lTk6jzdentvElEb8h979CWT+2ToitNihNziCTV8NYSCc5WzMlj9+Vboo4A1XD7gK
zvTWD/DJaqRLpHJ/oMpKSDzIrLNfdlSRXLXargmIQlrWRTNkHQE4wxh76J15Fa8Q
1wo2tl/ZIt37QHmTxoAY5YjJB07CuFi1SjtQp0LpWs0HQyWlkCkoCKDlF5gVVWJU
ftLxqzSDnzDHcO472P54BV90w6PeNMnqbcWU2fwHG8FiFYpiyQUzxclSlAn0Ltyw
EYVeTgsIlnFuV8lWwd3f9RNL6dGOumhktjyGCcdrGnPQAIw/pIp4zfa7RpSaefw8
cR2smYlTmV5mNjxM81SqfY3p5wXvmFa4p/XIAqwBy+V/NvjR3DRXeetRksUs8vlw
7TGdMMkx6JrCp3uealq8mQ186vlL7MjwIE6YBdS4qf9LOPAGc/cGUZbVSx1ASX3m
bQpuMGyg+/t6GFn4OaWSu6+DCNDB4POPo9Ze5JaIOInvquJ6ZbDJ4g3GKjpGQVeO
TYK2/Gw0suY83l2+LCgtSnk5zBiGFu8m6M3Es37RsAcnyvUTDgqXiqEWtGv+TGoQ
tHK4U9jyOktHscl5OFNV8h4iygmG6qt2p1YIiqGAppN2eHOmKIygXh0syq2UVIFn
QAWSQISRfeRWGBaEzDJPgJRCDCKBZ8OOgTVq9Z5eOym8JAdWgOa46EGb7VO/5Ia4
xoZ6MnKeycYJ5sDyByGgGD7sLLiNxx5SjeMe2rUpkEQYZCF4UkvoZpvWveNs3ouj
q/o7L7MNiCignWCz8jdI6Yts6Q+qYQ6wK8EukDKtxoYpG3ScJh/PslgZLeTS10bP
cPvZL3i6VvvwLQIPd1ZE7l467/du3LcMRFBwjDpPFBn1c8QVkrIFVG6yJLamCSmX
yrlZgEK4Hg4LkDtTZxmJD+AwgAUDUfy1AHpcCvILQ6+vDQpqAtN6zE4Vmn3yl9cC
xOH3l8WKCuYhlJxa0u/0Q0HWRBIOCiRzO5QRWJk/PEmnTd7f+bQ5pCGISwC89wM6
lrXjv4dny/aZRHGiZR5IYOg6xZ5zBw5c+YJsBKgtFIRFlonAnxRmWFClKq2L6tqh
vN7jzUNMnb/V49h0z1y6q4OhFzsK3j7+OriEA00QDFGE34qWYI3QLmxDdfDiKXVP
P2NDEliUkjK98yfDh24H8kwcMqlZ5dQkyXeVmkMbON7dDwTU50/TQWnksZp5vnQ/
s1IugvL7bnyeTtpsVc6tLukiBK9WmnnJQzYHyPWF/0h1NcyT3Ne54pyAlYNkp4qz
JNEpn2XS/x4A3nCJWd2nxATRdlUg+FPsvVEsfgYfNxarCkP77MpedE9zaqChAVCL
xug8IvAssVnBZ2UCOuDTZiHjPnpJNVi7ioqrPLjl2s90kZ9t0DuQ+U4dFP8T289k
dDltt7l1/aAqYcW5GqoRGZeBY34Fb4Z2Fp8q7ICuSvR3kWSx9g3ZzQsLh/nDi9Lg
bfCI13BXncvSAnnO1+UEXtmkJpZQYPHD68QVxqMwdyMX/2jpkRtS1fRxHNl1fK/4
Am6yDQ1EiuJLsrVfccQ3haCY5OeTTSmg/p+Cn1anmV4XYAHw7hCy+LOjoQnW6JqD
bm7AstOiOHb1QeO77e8krul43No/IAE1X59iTzZLqbKf7vGWRD5kl2C07UAS4ccS
LiiexKOi6795y9MFEb4ioDsOZg0lslBZu6dbLtS8I2XlKXUgoQ8nhgQz8/kyn5CB
MPyLJjPYfrLkLyz0sgn7/bk0Ch6vc7XiAoM8tsEsPVBBGqJK9ud3A3DnDAi+gQ9r
m/+udZ/WL0hPC1mfp0xfaS15Rj/wosWGVXiC6eWwTRbvEzVA9PmwhYAtTGxKZ0Kc
IgT1DNdhEvQeg1Wy9ePqtDFaWGiwsKA+sfxMVLJqxMFzoX8kgaFFqEX9/Iw87u/I
h0DJGf+4UFC1h2Q4ztPLsEll5fk5GOJVorqoohwRXB6esGgrQAg38NolI6GEg07H
Pz34iRtNorlMGX7hNThffSgyppubR4bcBmzglLds3aN7Z9Lj25yM/Lcl/f4ai3D/
cgxNRNK7A/0c92i9VbzQPxn9ADYKnAqhsfTz9PbiCtqAgob6xE8O/a+skraPJqKd
lQpsNO8rLJqmNaWWYbcdQIBGB+760E2+gC2WytRvzAOffOC+CpK/EiPfxCueqhHb
81wjzvL/lSD6FetK2OaMc40efpE7mKEKVeB/PLa5OwTAs9v0v+9iWmyZRZWgSX0S
VzUqcGuMsrbsYFuahcuRuYl96zkVebWn5MIfn+QtstJnMQe/Od/wgQGnrQB95rwt
bemaLnDaGaVu4YDWR3lwc/X5HcGPNKxnhAM7R6G53+Ib+P7rj1YQKxT8wJvSCFzv
yml0aoTJshViCeNa8GqQqJs2tb2JxWqwpXVY1zzg1bzyMJLXm6DepwWfRwKLoHYQ
T3z/KRFhepzXDuIMcbdiNKY6Bdj/3wZyOOveVTGY3doJ5z88poZMB2WT+ttQ30a6
WoCts4F8PJ3DQr7bQsXQYE497qQ9EycQ9H14GLDSwrn+QsKYaZSiCvUUME5UlAiZ
uCJUZq8clOg93NJDKjwEIG5j0hAlMbMMPFS4K30tSNMT4XxBH5cZF/uwgZ1nCM5R
atqjmXo/RUJTdq/yp4+B3p7TIanL8FjCA+F5Ctj+I8TqLWma56CiaSuo2IfrQVcG
BVy6rqdcP54xgivQ+EX3O1GgPBp41OU0GzjJSLkLGMS9oFla4+BoNAbAVBHz3aI9
7R78NU2MEmL0DdmKkxe/EXK7NhSEm1xCG+P5bFrNCe1H7+Z9kJrUv93+86bQZuPp
B76cZdC7ksZyZ++7koYJKn2jscIWUzayDoSKOhMjvzOn/Mq0Lyn49oboqcW6AMuV
FyKjdNEi+CFkko/qVsiSg+iwW3qYmU11f9dqFlClDoVGANCWkE2gN7D7bFWZqkZ9
ZU1VDooCQTJQBEKnQvVJagWb3IuWq2533OrH1MqKolcJXVWRf/0ry+Nw7rayOmES
nVcSC41ifm21lDIl/Rl0AReRDANikEjI/Qw0S59uNicPg52T7iCjAqKHHk8rBDY9
iY00otaJMDihBE2m8OlJXMUc6ee8liApHd7T0LACWQpdDCdqDNMKsso1mA0fXuyG
umTyb7WQYT6YIoUwOnNRZJQ4XTatRzwH8e307WmfIxaTQww7oPXgE4dw2e+cDG0T
CWDMh8DVi5HXx9C95APBFoZBrUyxwLqukBKc4wFLNsmZUqh+z9VrInnyXSeiotSv
DCe7nLO48g8tXWxUP0MvGtkb01LhJN0kRAYbgomVR2TirxWS1rHJKxQIIsUMy6AD
m79qkG/PQg4JEXPSnnxUVeeLwJni4omuWKXxIb7Q4IZUL2q04f82xguJvMWmPMKc
zkR7v930PpjoNOz2Fc6NKtYB8P4R8WYcY/miPGJxwkexs5S5iVOFzT2s6NXszQuT
sLrQO2fVzkMM5bgIDTpHz2I+alH7S+x6LZt8gAf5BH7zQSzOzkWAS7kfxh9G4ZPL
l3CInWb0YAHlDAKZ6rfpqApAJkrj4Ge5FMxWRxjL13NneyneZq5GPxg5juOc4T/R
tDJiE+fZxpZY8sYMOTjaRDL38PJ8ZjtCF0mHqpiOySo0ww7TNL4ThQ0Kw/8P4M5Q
9Ps6dNEaI6xMXOMG4XvyNEA1ZeLtE7AwHI6cAbDFFWIPhNf3umRTpkne+ORcTWAD
72FNRzgVCoj4V/aqeHuFLGfGZYfmvGpXlI0BRUXKPOyiEoqNyVLEwI1LgS7RepqF
7TBOgGYEkJ3bmTtkndCGh87AExATAK0Kiqd7+LpSG1FS/GXoQML3qlEQYFEa0efl
AVZtHakDJeRtMkRSDDCzNUGIFEcgO7hkaKvojJdVgDcW+Yu9NGVPy5o/iN4yCw0h
aqmB6bSWuEqWavjUN2uP7HcLhZFILhPBcRr2R63Q3ENOAMVPmhmWjdT5tdRThMlS
nwHwUsrs8OaID/mobBCZro77b5IuvB7WF08emgzWs0fSRJt0HG9ZUJaptNRzkO7V
nIgkUSbghjhyP7rNVkyUOmE/6JVgGZAu8YkJbdUQPk5S0essyc/2R0xbKKp61OVu
JymTVjnBFpPq7fGLqCygiuHIPTNkQ1d4hmfg4sT6hiHfzAuY4acNHs2F/3pkWRLh
Ca1AacvJoWkSfgD8uqtndKkzMPyNPuEyhSQpaTogxVsjvNwWThO2Ab8JZNT+NVmL
6UJA8jcueGlWANvcCBj2Tr3j7DkqjrfUvQxWi0ZD0HnRkBqt8mB7OE//cnTBX0AR
ttCBlcQIaeZ34DWMKccHih/RMhYBfVncom2A8Da6oyvhpArQ+FaHd+xdgRUBSkUW
7ThfCGMSdUkcGTQOscZbP6kdQUUm4XgnVFkwOA23tv6WhkUJzKpwTh1PMmR70CA9
lapsANYfe0Lfp5vEiucNVU2bc8mVFIqQPx4mM3+qdDzRjh2Xe3IvWNJdZ8AMov7o
ZCSOB+TIWmlgEMrEHHHqvQqPT6gMJDXqxj52yRgdf4PTB6xNbfMFpnkEwm2bbUAr
qGH2+rr14mPBqjm1ejpE3PyfwgR5zEDwFJQ8laH6n+WhTjzClSsJWlUheRDfsrTV
rY2F2ZIK6zkrvjemRjP9EydfzD2iDEmafYz0l5has7JIK4QILRrAHv5ow+/ZfIO9
aVe+5Gta0pEZoxEn7RlerftBTvdlVfnj+cQkk1zQqovpujWP9XBRvsPmI119v32k
z71ex4dTG7pOUyIEIIba4V8AxMlNPCnILN8DGOA2aLofRfnH4jI4t3lXhEyw6kd3
Xx3gMNUP6l4VJHbutqh8BzbuXdsss3OtB4mr/nPO0ghH9riweK0CKarnXfhBW95V
OpIoNJOL5GwY1v5ErvYDNFHEhmqx1xl4bb4E89o9gJzNSpYPm+9o7ZJIjaDBHsJD
r/jA1jQrjKnnS8++pUPhEPQ/plcCMnsEBSrnNbNNeJPKVQLmn3GAcibdQG/bTfh2
LnJ5FY2hACikdCidriO2M06xDUOtzGzUTRqNpP2FEDS+nxzxOZ5Z55wBvm4jFXt+
doVo4FrjH6x3EA9+zXvW2rxVcJ5V3QlAC4BTLQge+KJl0GGGiwvxOfnB+fZF3aHX
xjIURhTVT94rqTwu8t1kh7RffkWZYzCqRLjg9O1/PjrREQjhY7th8jAojSw+JO35
T2OWnhpaBsnhCllp9cTlE16j67g+A778YX3JD7/Ya3jA9sKKEuBjx3VxSYL5E0ax
KpufB63e6UEc+pWk+4D7m7sJRewIOSjHNRjeUq/VDzcNv1rUD1lvwJEYeJqVJIBd
Ufs+oRpvBhnbzuEW7fusIQmppLZ53RCpiTWgTlZCMW5NoscAoicugiUMCHIl3CMW
+uBj8UofafQznWpdBJ9A2OW73RePtOx6QuyZDgAwE+Kd+YcKiZEeP96ou+hdwRXS
pRQO9S7/QXoSXO3BHwdpnFBLYCG3eHbzW/PoFmn/KMT94EwS5j8mF5yvTbbsYbDP
JP2tslly1Pdl04lsETpXZYRqIiyJK4TJTE8/Y/FTvRrh+s6sdwLFX1WBvtwLBZaf
yRjPBENUoSB3E1/TXgF3WZG1qst6lJYNT/Iqsz4RNlcj4aSNh9Z12axdWoazJiUX
tfcqXffrZi9BemKnIzAPdG40IAyYkkR5P5z5O3kwz4B5S58JPEpqbM3V+T2b3cND
mZONe0rjqFMlpYRvH4LQfHWrtMD6R9rwhg2i0x80qvcyYOEWyrcytaXnlIGObYl5
ZeqTsdDzRRtR5Ic68Bixefn3oi2kUDuBDHoVimTLyAJ5Iw1ZCErVyL5POO4FmuHg
kOFgwVMHW0EqQxdrhC+vHMhxuT2SEPgbppxujRiQiBh8/yunHeV4jv/Ybh8Btany
FmZ1znCMzyfo135iB8AG14XGhtTcfjuf3GbSUryJWBMrbJ6FA6loPMuUt2Dawgdm
cxuRScyaNp+hiNJZoRuxkp7gae9IkthlJihdZs6AyXZGbT7LwIUbPaMZX/zyg4QQ
gqKUMS+Vszy9WejdVQIUfk3Fq32+hHfErUYmlYxZkRAqDIkUYlK37oWrjfxEquf2
V2fIaTBicFxyD6hIlnBGIKGia5ppq2wV1BrV4Y0hsi2VftX/bk7/+EmF1MP7RQf0
gG0FbxWs2Pzks+tK2SC+NhrQ9hpzWYdYbkw2OlXvQbRVhbExzZ/rYvtzlApOyDpY
eXbTiJ9JlK17+CMs6yrwzoEf9NapPVeZkyTGQ5lQTPsv/+LU2W3Gm15F3f5KrEnR
R6XuQS/sBoY5VVu8Iohz1RshRAgsqiZQApw5u/u9rw3de35L3/qdv9T4eBN2Lzrj
GbssaOpzT7xvlYM0lNAMwW91GSjKsSDZ1Wo0zqJZ9jit25mB3mI/zPXtC/IfsCX9
wFKYbN0kzFf7t4o1omFQrwup5OsWl14qLwDEuLAuLh9quoIzZMgOXD54fu4dMox6
/1PZa+3GnhTiScyuh9yRPpRMBItpa5pz9VTVQ2gqTR+2SjgI24m5Mee8ofdV30sl
Tf+xRlPX4uhTb9y9nsRZrHDm7QS+3V2Ksn2lLctGYYVHmvAQOCQqTp6qx6Vlm23t
E8gC3FKa9/B35dRM3YT4eKxyH0Gb8wAqMO6ILsksnkI42w5X1dsQhfx9G+3lk850
xPIW3yUVjB0Psl4LD8MEm5/Ge2vSntz9TR0t9wiSTPoGa/w424tFA+OIvsjwmrqP
jtVG/T2RdcBoCUgO93Bxx1IValvfTlIrEmUsgrkXN0dIJC27sTp8ewc3x5NYmU7R
C2IyvQTd75BTnzitTEaVcyqTNrdIN9dFral6JbA3lJVPTp2LxAxj1Pd7FM/X7B/4
cnNxrCLvufLSPv9WwvoLz3VYOT+taGwD7+bEUmV8TjEbEEIi+IWkTPd23YGNvqcM
svusGh74SXJkM+damHGc6+9tKbKratgSUtWS1iJIoEOXB5eWpTF69BFGvd95Kz2t
JB+L+9x0sxHPqIzRkfTvvdlDxLy4iYG0ZgYbffA0W2njoPfQr4xi2wyPolUe8o/4
a0jFhV0eL2YcMq37Xf4bsirjd8NX5uRBB/mvXkm1V7IvsF5rTDnxD02LnaGpJ6l8
eeVl1CwU0S+F0dp9TiAtxTjeaYn8frlnN09W2bSxzo0H0/mGgeYPngSWwpg9z+yQ
YImm0OjEnJo0nHBoGxr+3AR0XpZ12CASDz5qk4f+llx8cuUC3nu6u2T7NHg6T5vu
Q6uPQ01V26YOdI+V/LOx3bQfKzhowF7WNEcLG7mlblwbykCssdHm0GagmwnYwjbl
eYr7JEJfj9QrAt90nuRZijDNKiue4zjcE8telBZKA9tHvtLDCAKDU4wQ4tI95LJw
Yw/X93rz+p0Nu/6kZnZQjGQcv2OlINHkwXLsqL9/44Lel+CTBiK2I9hdeKlGJAJG
TimnR59jOoCmKEyCQqT1Ep2CObZj51Sx7Uup/SnrepRe4Vznacaej4unG98vf5+Q
iKnf7G4fAQ1cFbx1k+sayX7u/ovfJZCZnJFCRmZbvwZcl/Fe3dXl34Q+txT8BNjp
Ti09hIdScLGc801H2VaXcy0+1UiLtSyKE+Ac15V90eEXKaEY1H14eoGRTtA7alv7
q5st+mbaBmVTOrp32IPgg+BEt4qdi9yGl27Gxzoeo6jPtAqi1V6nkCPaEFiAQtej
JMEKA0X+5uZDPWJM8msrKy3RiZLeDU6t+xkgKXZjqvLab4QzH9NutAXxAM/YSN/i
p/8D+HqjrMsn18Vs18F9oRdR/cN7zPGj1OS/gc51Y1YpMtEB9P+pgo0+VeobSuk0
Atlj+peuCe0/qS0qTuZ6fo0k+b8VMmxqbzph7C8u2/pE45CJ6HDuX8OWuigL7UBJ
KHITFbMMwE2kISxpyByS1l8iCzAJxzTRyfg7eFnqRhWZV8VIJok9msVc2412h/yD
xtwLfKu7tbc+YBcToXSMdtqjq8HVD2qKSGsxGjqiCW/erAiR4SIDk1OJKHcQZm76
n8xzxVA5DOEWk0ZlWmnMlmOwk60yt4NDuskaQOA6fk0g+Wev0rC8UvBmzJIdBq0H
uOxhs/jxudGxw5Dx8M5F7/+LU5H72XTG92RPgdrLwCYT/AmRJMo5iNqAIsqAQA3K
7K+PSzaOJ3gmjcu0WxdSgyEboPmPGzRuj5BYl81p0DRqm5yKan4g4D4eB1VddYXx
50ZKLRyGjKpTRNN/IzOMyCu4ETOzNUFkIeimLrQcWjMk8XYzrplvZXW4Zr4dU9wi
G0pjFBDzMez6CbbuUnIwLX2vfF/4UzxFH9i9nAYMHm8CNjqO8rTu1gcM6JknZeSv
Mk385nhpQsrTg2K/MM8bKe2NN5uWpA1e/KZBYbhX9tmKh1sljOYGCtPulH42I8tG
1zxl1WcibENrBTK8jSf+n+LbAwrJGKukyhd4OyNc/hos+vRtzaznI3qWojDOIlK+
wbJ+3i9MBglOmN1C1PI55RcGtPdNfqHrBXA9sUldoWR6Dn+Pi30kXFwlGMHM50kF
oCnas8+utDo0xsvvfwQAGs0qUY/hg93x5oDfUDR1LdC0xwR2YnF6Cb3E4OLS4bvg
BchNTY5R8IVfwgZ9HW5xLKOuM6MHqHywdr19ste2Fq3VFI6ZagVWOE/jeiQfSRIE
SJM7AahAUrmHey/ZzNPzS+OyF8kSRVjCZtPEWs4gjBLLegF2FvamnUrhXhyk32FK
y6850gKu9sZ2n3bEb3EEQKbIImBcBshCIXqVUCQWr7Gqn7M9pSTuNjnLoUyoBQQE
SZ5ymZY93PvpSvnG7LNIZ2AYHqP1kvMGwRrk8tSv+gBWrop8z68vsFHEvp+DNC9b
MwUYAJiQGQtFOWhpVwFAIt86YTdZ0DimaLN/qI6itrmFovt+kBARuGdW7JeRFcao
qG0JHulmvxbwdFilCM6UCfdkWcic6bZENqmBN4YWoSBGHE1aEBWw80Bx/8EJ0GJe
AxQEX+j0cVvq9Nhcz92pBC3+iXqaCVbmN30MKDvUHpLnPYx9ht6gQ5LeO+gMhqZ+
AJS3Mm+5uhZh3yLWuN5gwgd6J2IDbLGhdgau7aCMLerv4fnzYcQD+LwYpUDQCGvT
+DaDlj5+AWoz8sUP+ZEhd7aKjvu1F0BZsYn9GoRMfyYDIBS6yFOxNLi/qVAI48Cz
JFcMf1Ezdx8fO8N3voSjIC/rlAhhBzdTs1dIAcMmJ/lsbKv2eANRmijQ32Xp+VJq
xcRYKRWtAytKOEK61OjzLJzoLnpQo9pPs1BYHNAjcR9kF1G0eYYR/gIm9HPCuS9G
0nHBciVM+AoaZ07wnn+Qm4SE1u2FCoSQPrSDM0kXaTQ5/LHTb7BJ+XIzVvt+NEpQ
JbHk0ZoHBXQ+eB4yb8ZhogRCTp+WFS91vxjiw19sNruafNG3fWr+fGdAg6ZPFqbs
F77Vq5+0ZkCMDyRQVUbEH5yWG5LJqniLXaFMaeHiDERZaKXBZZvC3NZ+jZCW1r39
gPd47r8298DmJA86q9Fwib/YFrUK0X8MLeJZelOUBJo8mRwQUpKR5ZExn22X3ec2
e4MHiDKVYhQE4KoGzCptIpAnUA+d5/PLGb5ZbF5n8ckvvmNJyhkVLeHhynjP1QCJ
VbQ83MnJi2TzZM0489SwD+Pfy6V9CegZVBiqZlLGx+CtjZ0HH8bphs9LGyI8HdBX
7O7ItK4p5fQoaJp0Ry/+wExxolBPEo7Abnh7HF0uw+YFPif6Oqivwey9+KbHGojG
sHCKOs68FcfKrcGT7GvnOOQas6E2r/WLQAfLZpaqHwil06jYgLmgzEvwkSxn3/6r
6Bn474j/hnNO/VZb0+iRiW3ZVxQSZrwt2/EdKTj9Ky45TB3issZ+rGXt9+ZTqvxV
2sYGBhTvOXzU6GgI3e6gjgN1lI9VXNNF2HN3jHlYwJFAwxgxBxJjwNUPVkl7CpEv
i3ForzVl4E/6D1mCfv4KH1buyb3msvwSrCKsfUVfwwaPoHFBhPaZDmsRgP4RrlPl
90ED1knNP/1dbSfpkTcHgmhJzoeV/txW31J1A0X7FY/HB/eATVn/+7tV5/PwOWii
oUrBuvJOv9S4miTeTEOKlmjIaKc8Ttk1cY2a6hLH/RchmDyaM/0Lud+eAEHpJqXA
w795SnEcC/wiL/DWpCKqgD+pYtNJ+aqKYW0ZPkq4cUPdV8Q9UFgOKwWpGTSAXJWC
+xU1Ge8QH7G56cedsxpjnMRxUbhQHjRkkicDIikfk3gqaxYoI6RJK7lZ3ykXUGxD
SqCRi1JLfm8AM2BJfN/+MXKSiuS8JdOIImdLGb3bGPuuk3w8jiFto3DL8wVUAKcy
dSBasFcTCPi41wS6Uy0eKhnToCzxTgaaKijaVTtqNDWQhGvk+WpC1bjm/20Wlj9o
jHMOsuk2KYnLPBwqbHxHoWACb9OS0gz+f+J4FC4SMTXdYal6+CtpvBgLy1SNgCDD
p1uNwj5zpOdPQpOG9tIboqI7WHZrm5aw5ORuAsO4lRf4FeSsMjv1uGqucRqhgAQs
graLCcG/FLwtwC3S5mUPG3zgTDq0GCH7kcglsuul1yz1aGx7IZ5cPvqxYriN67nd
33CLCA7lZjNvRoVGn8fssNjcAvITihwppvDc14H3c8aBU50nCCbTXIgH0scVZCqJ
vkoS2mruh5qZPabAqhTQYde7wNY7ZE4TH0iq+FGrBUXCJNwZarnp+pKwGDPkqkfL
0o9denJul+rBM8x47w2RD0Xktx6MRd2+2JULWn3HRLXXrKSdldZqlgkD+mHQFarT
h2i5IokucbGo+6r3rWwsOJDz7yAw+OvneNA2pDqnLU/yGy6WNdyj2Mwc+q/BKFlH
ZeYT6XcNqWaWCxTMLLQ8bYuK+AYw1vaqCD6Px8QyFnt0mQI+fHgrT1Z88PiaXN+V
zYwd7BEAgs9gPIIDU4yIdt+socuZ+DMONmShUakdbZIHgREACRHKhp1QF20uTYAT
eIWep5O7cTX5a4oPk9VSIk5eonjpDagSHatD1dHYq3zxcRNe53wG6Yx1YUiy89vJ
9paVisjWk3aS9f0E7Kb7eO+uHseTnY4PVIsiBTxTEvAJ3aAGVXt1tTkz27pYAJOn
UvmHK3pIug2KVJhtPhnE/R4CgpqMzx5mtj6vNqdTbgON8RawuKA5gWnXhAUqT3Mq
Yl/HDkyRqpP9KUQAptG4DfBO7hNnLjREfQIhUv//fhjNW8UHdbX7BvG7K+Rca4oj
GvtO+AA/CpZlSI9VIuedv8FDbYmXuBCZ+ML7sGTV61a5FJkvZQGpdidMo6ibtAxE
eOO4sN9wULkMypVuf5WNU3yJr8JVBbhApc5GOrVWbbUo/F9JqL+wsbGXe1d6tXe1
6k6s3xeaktmB/LH70ihyDxIOb1ObfeVYlrzv2H2CFNMy5cEeoOWxysj5p8K7qr0F
970H5wprzeVmXMKQoZeKtm5o4rNn5VmNNJWt5qxuYmKO96/ehT2BPu7P8mCxcnaq
EjB5CPw0DSqzJF2C7T4fKU945Q+eA6643iE0UZdQu0jp+QufCQVPTI33mIqCTYoJ
QR3fjBuXm2apU/d+duIt+a0NFX3htBIn6oN+0tIuAoM0SIdj8TxJRiGaNLo26UUy
T8xFM0vOSjKgjCwxY94A29Zm/xQRAAROrNGlZPoyydFR+m3r8C87BPQuDJ5e7ZiB
tqwCqjyAriWyn28ZY1SLd4YGxq/aJHaAf7/QIpckeokE+ygqI3xPSS6U80SGutiD
WALSM37YyXGCypOTNiXWuXWLmh8L+/m41qmbCO2SKGZBIa1meqVE7ZBaBcFGoBoL
hjb/PgOMR1QA3pb+4JHEAngfZA4OyXn9SlTdwnq3RDsvrams3lMXsZAXrM8zniTm
QwbArxbm3Lnt9hug9tecKihlKfsIbIMafsDHnHN+cOJ/OZAbYAeh2v8umbNVNReC
zcWwvmH0tZBtFdvku5lNEARVSrukIHrKUmf9OlxyVqmrAqfNUc/ztoNFzfzmNAy2
GQkUUIsaEMg42B+tyIgNTKbwM6lvBZbT/tgkHUay4uKtjz9rXKsXQWn2n1hafJ6N
VA8rw38aLXc/hz53zulbtXUOEq6x49XypKwI2uKic6WaY3ME6rfbskyFyXU5Nfjb
mH9qjANm8WywvZWqmqeVIxDp/LH/52l+oBYqmqXOGSPQ2/7xOIkSzO6YHDktju+p
M5mBFDjpBRWpr15lOv5UoMsX47OE6tzAGw8DDxlODSLWR/gSfAxNBs44NpfyxVyy
99QG2CuxFLxYCYRopBN4vwHyj5vE8U2IB/PVzv4hbA2NYmZw8fcYH91+SraFv+/C
LC5hWW15QSBRqkFENc/VZ+oJW9IoCo2V/5wFmPixwdQboBX8F/RYrQojLJC5oT/n
XRkRZZXsX/ZhCVVBrkoGWJkulFZmBiQ6bwEzJupVGZcjnpsfU+XDbcH+C1ZpIKUO
kEo0Nhu3Lulk0S1wRgyiaTqJWOBox/P5nk0rj+L/vcFxnIgbLyOos5ZQaI+UqRx6
7GAvk/eOI3KnOI/S8AXBUZh3wM0uRGatGUOdE7B+svSDrFPY5X0Mp3w6ZoahToGr
th2yB8RRoQpoGEcfdIgX52QfD61SO4yDmxI/y9YO/klS7BTazON7ZUSHFz8LOmq0
ut4v2/rqmzrTOzZzOXWTJxdh5u/9ZsImOK0Ox7dIn40MhfTNTQdv5dqx5G5+oGBQ
PF1oYKzasiypxpi8DB//j5ikuscaU8vFMs224Y0jWINpY921VoOEpVbWjd3v41QP
zV7YX/HwCkcfWkJZ0cuJj0xYsRK52im3Tb0eX9eia1ElYBjrAFp6hd2Uas7yCg+h
Ax4Varg5PMj/0JZajMWktNUC6C5/NE+0d7hndCBSWxikCtnC08aNPbniCUIv4naM
02E/NE8B35uRTOcKB2z4Rk1+63kvSmvtS3Fc1tZKYIXW/bCOYV+I3kJDoTMfPL3c
qtb82wnNoazhQIXkWqnYo7QsmmRty/TR/9ByLZ2SIEUjWUZg4lQzC6f70ZW2AmPK
IRHJpTpQ6nKZ9cfLFQQvOwGOAb1PfeoM0iAEfAwBtiRTmn66dpVnBY+YBjZQHhdn
V/B7+7J3wBU+4vf9xOUgjur1cWfyQq9h+aAWEnOfxlHxVH92PC+CHNFE7B6WhxAR
dGn42YDxCY5wLwwvhTradoryCU07M9mu9AivJbz6z4lKoZyl18BCcDNr3fGzi4Lf
f0ciJp6ATfrcgkvTh5JeYPq+sw86CIGh4dcQc8zLniYQzirbEwRCZ4Z5NflyfHXf
J56YeQSXHMvMHQHOMhnlTnjhWYtmksZdHVhgo3QgYU7UMNc159FqQQzWHWBpPJo6
6oOBILnfmmrnkL8BM4/2HPgqPn7c13USlYI6CvMtHX3XKzeYaJusWj2935oOr106
ha6p3hMKJd1j/PZafSnaNuFofOKduKsSk9ZmaIpoDI8yV0zHRxDYb9TFrzoUJ1fx
gMmH1GBJVqshVWyIk8VGBCAyUhTud+uW44DiKJ8mPBo+e6v7TTSCTYa3JS2rWnhc
xRzMl4bO5JEYabJ7Oc7zHcN0suyTVTjf0z+VxMcwQCiL8nIWCfT7DF8IER8JiSWY
JrrZDejGzP8/qpg+4R0YJM/lY4J1WOQ24g/EfWu0QDJixIZ2EV1CCLIENmr1BF6x
QBdpVPB0M9aLgp6cLDhsJ/UrcLBrns2ydumsvVtUcWwEisyJ/deBZHlCwSvPENnE
KqDrLovYhDTAfPHynO9l82P/kScLtcOSwf00iYJxhlyknbIwoc6L0k5LMpBy7q+G
4LdoiPSuWLZzvAsVU5W3Li9cQ6hOx0QLT1UCJe29Q6yst1AQ5CDzuldxgG6dfhW5
9pUpd1Aoh1LifVxE2rKu8dbwYyNQW+j4S3awOyayak4QyUco4br7lWnTk0Ck3Ntq
7Vcjfq/0CZETUEjm9N1AY8LfD0t/oMFKp8wTuoogLTCskANWSw/6aUjA0TtaICnK
mf9OImTyG+jiFVzdNwlqGslQANtshvCSh5kyCPx9jNRrfESc2EdwSuVgqLLmVpip
BcC202SsMWYlIhlp9kMEA3wEn+oj8RxkNsAYb5U2ID1bu+CEnCpcZfdO/BBvOhjG
E6g4LsFGstQd+ulTDVM2fjWpkhrEzcuWW9Xa2r66+W1abwSIM7L1sgZcrHirkkL9
CjCmjPoOpIko6LJf/o4ER/C+//oPP3JZgpJ0kifxiOJYhVSIlqTsGe6yqP5oO63V
8Koz/MGgddqtuB+xXLt0ESvDd8N6GxFo0zQz3cRZysFqGl+1Hl9j0Pl2H9wVKThy
d6ryGbtc3lQeGQXBDipUIIPugphE6Xwz0uK0pTV6WKP2khVteTZHfezeL8YFCLLj
Jr29/vfECSRD9sugd9xfDcdPbY/jjApTwbtP5XqUp8JcgMOWF3Gw+83LdqnFksWl
KcQQ3lwB8FzBS2ORrRciHnH+tnRVxjgJh/IoH71b3jy3SUsqE5CnKzYXuOBJPw90
epUdTaDlKlSUHMOpC5WhXCXR9vVlnKXm9Ad9jNC7PF5IUPAj8ghUF/H3q2IutJdA
7kbV/kYjhQ9vyH7EyMtTk7eOY+0rr4eKtHpBEZEHTMSiNYSNTLqdIKobI50hH1SM
OYnmjlIgbihJDCw4CbUnuE4QBTIR6sPPuPGO9K24JVJJ+zP73d2iZjsWDvAWWth5
/zHgUEp9a9NtPM97NdwMkqqZfsHM2uNjHHiSrZk8rcjK0qbJBd8N1kG4khGXMvDh
zIYFbroN3yZ2/bhI9M666jH/myHHJsfWcsE1I2Zicz9FnbiPFIqX3kCGtF4awMke
4HS0+PhkE8aOAgTsdLo54iIxpof+4luhTjhXBTWpHx3OBSwxYbvvp+1BkNbJwBfn
eMxYpp27HOGUQ8dGbKLoyt3pvRz+oQE6E5/ljhRnLmUOqtPp5WkGoD7F+jFBzToT
Y4rWh7uj0Ty1r2rgv2pgy/lsAPnFMUxjLgiWk0twy8ZJRRAZJkyaiP4ZamFhnHje
3BGIAUuAU9PJNtyfXLQ9pFNH2w7HowRkeK6YK7of9qobMt6Epi6UoLBuFB3jmZ1j
tsN3DITn0sCeo/mVZvrTZZgTAE8DBjxTNs0JXFXIy7RQbx1nNTUe8IuucqQG5S2Z
Y92mo9T3DB1OZWF7VVzLGkInhHdowuM4uDEvjYGypyPyGlWN8HnkpQIj+CyIf9uq
zTg0Ujf+zLEiloD3cq/lb+xHKXAHRgzrBq3db1TaFbYQWvQdjuHXoYcXFpGnX4QH
KlYUGP7eu63dK6cA/vrJxrySmhjxC8YhtxVtkxj6sh3FO4acKXxXeGxsS00U8vqM
l/MfHCOgU7QAcL5vGeS4Yu4hWjUw07D0XYqwQZyIGNnnTb+Hck/bVP94JoSIyFc4
tFm93dX4v89gmrlP75CRJiUFVrEjBiIdx2c2XBCuKxXXS1UUKhZPayleqQgb5AvR
HFHRlJzLAwcLoP1kFnQsJGI3o7yid7Q16U4hfvqWAAqsmElRD4WyaP4S5KWOsvoA
4TUXReJxm7qNPdxt9E/IqOMX0SAYPB47y0qTLme0DmEtGlC4h+hMab8+rh0Z3KfU
saHCzZI0m0NyROcPVuR9Bn8V+KloaO1TA+NluRW5T3qKdKtS0I8nkPIOCaovBREi
xgTpBn+Z/Qd/LnK14SJc9zjxra+UJ8dogmfshJt1g6KnVpHRpG02GIXt3kpXw3Xq
bbF0RbYZNOjhW35CZ58UymddFafW6ADW9WX3pKJw3D+/+ccXhyPBrm+BQODkbjRS
fAEXoVl6OZqy8lZEioq4DCCUYr+JISZUDCjza6EWDZ8+ZQVEZEicepES9rJnpzrQ
5zGrH9jPJX6/nfD/77vDRoVX7DcSui38iNhsX9BWhohH1WDdApr/jHod1ZRs8Txc
FIC+jnU28vQf2gtseTEv1dWzO0kdXFYkKtpuecVz0PjkvSntPV9yLUA8qSKeIbog
A6pizdJQ+77xykqc0v1TJC4LMcHTNEIG5F0RE5WoNxOV7D4AfqHLuVwjC46A91PY
0Yzea+2lCfWBRFQxhuglxz7wklU+FSZMaTTvVxhUwkf8nws0UCZ1qYlxpW9yyq8K
BJdMF+kYCzPxYZgcahWMR+VV4250kyjHhWMC1G/V0LEIdwvSU5KDXyIVXlyMjYHt
8PXAALiRtkrKXk5rMoEXLX20wj0CGJha+6a5jVJKhsP45JD6uyTpH2G4FlVqimTo
wZ5mTcFrCl1EC6hGPEu2qjKUmxdj/RuDt3K2d8dy0vsoFSbcOAMEuNTjx7uZewrS
nhDp7lcqIXI+z/lvDnjSEXvxoHo04nKl2VASySvTO7wD8/aTGcaS8HxPBFoVksSn
ZFOV2a68cwSbhVHYk4MFcSMgR2Znxx9HTwatUXIwTnZEzfoYioiTvff5Gz9+6UUF
n5HPiVdsHYSrRaoDogz38rBeg9+DVu92LXtLwvAQaxQHAU9paoZhBEWRgxQr5J2u
M5x0AsrSCOj0HroCQZqDGngEQzo8yMouUa0D+jTknsy+EOT3yPmQBGEjlCDQKqgw
h9E40weMch1/KUDcy7MuCF+RH9Os985ORg3xQozKocO7yLb9OpoSSfuUQNk5oQIO
OZFtcWadQJ7O6028BoxZEvNqyg0YdlM2QAnyq2r+TKu4LpHPSIa4Jk5HFZZKVmHA
7290n9Rblpw2fQiS+HJ+y0VxC+bzgIEcIBwtjBxmcSz/jJDRV1m9ZUqwpg9btq8Q
KT0qu7QezQqrjZPJ9mv4jGlpjWcd7EhiYErXn3DLaMEX2FJ1RtPuwB+k9B2JmkbL
XmyyKkzh+Tcb0lNIlmXnrfkImqvQumNhSs9h9MB3tsjxQ+YOWYhIicvAYb0odKaf
WMropMoZQIMB73UmmlquGwfZPkEjY94Y4lAlHXglWVEEPFdEG4FFikqoymqj92ZL
PAEjA4h1ckrbWccyNUDCv6HgU7OCgv2auET4euqSokyMGxZKymPgtw5AIhaLN0aM
TMxeWBzCuKEeoQVZa17wXdnnFs5FvY1muG45DJ3AHBxssOrSqEko2B29W+aonw1P
yKwMSoSw4dlH9zoO9HcmZBYcaYKhmB4DXBw8OTo5kQ9z7s24gOsxiNOR4XnqYo+Y
RdVWatI+KgsbER31KLkExoByjFL2UbUlPkwxcl3bmfB+h7LRJSmL/YVJU1AkLovF
2JxAWIbAOe1D4xzNZ/zBMF6nybzODLrIcEVuC07dS5vHDLlZAhM20LNHaFmZ6dMz
hjIrsrTBPlfQ78MpMtklqaeu5yDitdpszKhk+MlPF8uvJKtf65ogx19ZbI1zWYbb
izbBByQKQaZIaPleRiTQE6edkQp7oFgJoltaaSK2jqfhnkFZggIv68y5I59ksyhU
dyyYwg72/G5takmRTqS/KfElWqQVAO0uBc5FthjGnyS+XFDV0cubqaQYmvQC8o8H
6UjantAULjH/acZl8dA5fG0PjY4Z1c8uYrLMF722OdSbwBDmhYFjVyZSbZoJ2zvv
pDOTYjwx3ez37p0YLsvot8gzEIghnsPZKWDDoe2y6/Et6wGsPQ4HLEaytaEgTj4m
F4QRPZqWQIz7koU85K1ZXmFbWLO3hnopGy5LAbXeSuztLEoR9UfTWwP0swBBiROA
h5gPdACV5/p1gzsyl5nTRXLj38p+okyQoM7InBDeqfk7Lmi4YCaI2dz7d8UHd0JB
SYLwF7ypq5KdW0ZS1iX3QTTaPy3hqJKA22/4marSZ4IRHlrpqsRcb4fLZpOxW2rU
/FmYlepDbStND488LJbty/H7FUUJfpITVyE1rjOMf9LE1Md5Dfn5684x1DoZGcXy
c74v0R61bb6G6M//m3IJ18y3yl25QKjgcCL6GAl5pIvP+GEACc8gn1KUpyMXOL4Y
gOTsp3bTHZPDUihthSLL6QE98qh1zKjjMbVYrqiD17/p74XAT4/8wHlHzI887FoC
TzxsMwrYs871qEGD+OdsdlwhytuvUlQmP46fh6OJxRCZh7HfhAAudkPgog7Ml3Tb
vMau0ova1Vf4uwoNL9hnejwkLtGvnxpK6Lbs+T69In0rFINDw/wU/QI0md5SaPzG
KtJOw27WJoTuZGZk/MF0W8yDoPZJ3WCeGvs3G7BF2UnExOfyktfOeK2rd9fS0JRP
M/KPFrWqlzzw4h1XIqnCJeNykIviHeH1vAy+O8fWY3E/qC/fpaAjnbKCNnuE9kfJ
qbjtu0HMPcgA/xu5exTm8Lho584LdbSfpzB6D1pnOOCZJxgc1ipkIfA3yEJ+y5iR
7B+2a61/y+JKDxma5Xa/R9H7Mgrw1tuvndhhm4+bk9DlvEj3AmgeqPhVDWyEU5iX
DGUMggBR3ZNAQvOTB1LpE8GXovlVDEGn1z4ZiU41WuFjbkEqAuX4012pE1SaQUV+
BGRUbNfT4ofCNR2X6Z5YRwDzmmpRjiKOeDjocJYaifzbzODslV2l//f0z/YMPAwV
Y0XxAQ2WzvLTa7oL+la8fesZzDCZzYgKrUY4N7I+DjkNSodcZqs+01G1gNZWuCiI
VbKFIfKQUr4XC5fAqLsQLaKTM8VVA1uQL1+Q37cwbrwbZALMRyzFa5zrT7dvzUMP
CLVXBlP1tRy2MJI6u7LbAHBr/bB5jOb9SebY6zM5jGOOCf2nsDDDlmqCqxF/mquf
tZVjhNYmNpnapdSFuBrjtuYdibRd+4fHpLUN5vIt7dSW6dKev2m+oJ8/WrbRG2g0
bYBrCabHGosF/6A74tudeHjNUd5TiU+guqQYU3oDOk39y4oUV563spsTgg9NCdgN
GpkiqePF3+KnqLtWcVqtNKxREax0L6yvY9wsbqOHhixddeAIu3eJuWRQP6ynWz/q
CS8uP5Eg0QYUEORNkpGHGYamYVN//Kw3bYrPRA982qk0nExNrjEyfvLrAtVGrr80
I3KUwZXp2Aivew1Nz4AL5FWsUAXqvFWTXiTjEU/I4d4swZRy47fpIQLrL0PkFIw7
W0BCMaoEdz/WqGPKSmZ15n9vHcH/sxcoe482meAhKGAmDG8QxAaEwu4Ty2JEtdWm
if+ams8aTSo+N4cAljJG31VLalTobFF8d6enAWpSJNHdIhVYLKgOEU8rDZZ4xoDP
P082bRo4zZC7/aC3FTP8kxfMFqAzxdWqUbcUE/g8a67rO0b7He3RTgt98YU3XE5u
lRc4MD5N7b3BE12hk7GB6pZzQqaRecO+b/nakAJAtEtH6KhQD466wo2BbPUEFzLa
jchhwthx9LJ1YXLo7Gr0PnnjgJeY6CMtjKJFYdsTDrIQfm92uu1BS+duz3wLEKS/
1sK/JDdgcAn6+k8IAYBRt2qdqta5C8LiuSQnowgrzJMbGGw5upHq6nKbkOOVwqGn
kFICNrcQzAeLG8br7KafDImdQt9+nwdyz3/LFrOST4PJkZ14cHNul6GtVjCZdxAs
85Tb2N6rSszlyDIMVwwKxldFTJ/WFugMkCt/5qwYiaxUEsiDm1vPxSWeBnifrbum
elv5oPCjX7D7EspyMfbNH/jrD/ZD8aaoP3iB9S01BMOMVDHMN9mFPSK/zZPeVD1r
nYi/E6DzVBfZF+acfZdlv5Aej6HY251qz+ceR0ndoUctf6SdoAR7hQgFhkVZDE/0
J45uXIscZfVsKs8vtnwj1KGjXtZyFfbNK6zkpgiV0ypJOFiSEaFUVIbELeGOMQKe
L9IJFhPj884BBC1+2QlTP5Beguvi/h7L/u+CQ3V1wDH282GkQjL1hT8NUTlSjoQc
RLmqp4iJuOO7Srz/jfd6iQx7H4+9l/nuNEUBZ9fS0OemTJJ7GcnuWpfxKF51hibB
LlAONzXDVZRFe2t1pOfk6hJn3UtS9+xKBcHAIsBKExLnQAjpyMV7WaGlfI8gYSe9
C6+9BsIaQ9tZVJJD7LUvSs0TtPi6yTo8zYMqPvcEemfNnaBLdchxKyYq37VXh0Cx
CR3v1hSbqcL/gCRXBwbNlgSBFZneoQOYp51dDuQ01C5m3nFegI3UKemz6SRXjbQT
Cs7S5GpNwKaeHkqKpRgSt2YL8w/JCBvFfUSOmhAqdRGxX5SSW8Axlo+0zHgzFDRj
FfdB4sTqdnEPCVH4U+1K6u8yYDUryO8uZzm9VlCyaAHQCZCSnEFyvxo5k34lh1MP
NI9GW6Ouzwrctash+E6sOIzQFJu5NCX1LATO7A6B/BsbHJkJWKH5g7ISaaa81VrM
ekrwbOARgiou0smb4nbW4EKP8T53dP8aiWclDUqmKmL7xVGwFS0EMnqVpzfrzumI
02HXWPrKtz300HLJOLNPF07AcJ6ho4T6T6jaPSjT4UDMUE/jZ/pmzZ+XYQ1hws5R
oiJ5SmE0yHoV9JM4Zkm8I+GMM54NApEiIF04bvdeCitOFJmE/Gu2cfvZHyg+Ti0G
e/w+Q23X1YGAe+8DLw5nWx07AgwHa2HIVKYgTwvslsA+qCWXexwCCTfjdj7tGF0n
9enn/DnEAMxbTCkJtJV1yMmyczWuX45if2GnCRWFpepPJNXPGg/RTwdGRzfmF835
nXzQFqGhZ5/KdKae9JsAi+b+UF6Mu4YCICem0g1QtJm9DlxZ16rSUJvzdKizN1jJ
MQJeiHOVumlXykTFnLKH92FqLM6k11123/ajBggsdnVfh3u0P5TVedaY8tqhQmUP
YG7I1GZAj8JMSwViRw67bnsLIT3CT2y4/AfEJzHpkQ8EX+WcwVQDpj/r/2v2Zhm9
AfeWjPSz2ELvbhgUQt8ay/EKBEkwKrWD3W/tKrYrUpI/rm04NTs5xosGEA6Sud0q
Vkek8nwTm/UYQS6z5Wn1Uc1ogCDTm+LSlYsSOwTXZwF7anQZIwt4P1ikaaoUVIaV
IcV3Uky8iD+hAO8JLpw6vIhuWRBaYH9+NSa/lrc9EzSvfqknqDMX1Di4FRJwnr+g
6+csHWaYqaKRPLOdkv9ulsNrAmX/Vek86S4u1KJhkeF9C54Ub/b0jhAH5cNV7+/l
hi65KZQ3GoBb//HOY7dfR4NlbmvBnkGhmVAtua076zo2hiKl48pCLUp3COOHnUcY
4MD5QEuic5RR9UGkMPkI0R63vum3j2Q0cm0Q1aj7vrWqdrkixQerlTvPfOqg4cPF
qZg+UeCy01NbZT8h7qtWgKUu4Jv62++uGcdcqJXTZlvjZAu+Me/O42xw4SmLjxLp
PrBo9XXgllrasNQKqtA0Hmm5hj22gHC/EVGJ5TC9f4Fi9kUimqFfQcKEewmxJrSC
Az+pOxhR42ltvvGt06O2nuI7tuLw5BZXljCn6wztaqgJKJ9am9S3H+l1Q0tEvifA
brqxaBl6wYjZ4tlBFAqa99YNiBMfPUyfJKBzpubAcQU2cantsTDy7YCSbN/OATMz
QKdj7HdZakTlKtwuXJ9VtqKLYr7DlAJ4zK6T1liwO10du7A4l9xjBBzSinN2aMdx
s0snMPuG6VnAxSiqmY6Qd3OhJCCmU6dO4N5Yc/M0tqm3w7KRXrhtZ6UihRZH0hS2
tbD3PL2MDUDoMshCRkoMuFNGpZqx3fKxv79KQbvPCofO2icDp/sweVgWbBZn8D4o
NzqgZAMSt+xPvyzb1g26v0JrIJeEomj0JwAYC0teJ8OyfmiP6wyFrIEYWHpGhSot
EoqH0+ljKTo2q2EiXuI01A+P2js76VJhztBfbtEvvMCGw22ONSfZ3rKlwN01aA3C
PmvQlsCr51PB/Qspa36HAC+fJlahiFPVd/xX6oyyhDgT1Zgljl+tgkVeMaoQXDCg
P0WYdIN5CroJGVAIbopj/S49lYIazO3neMu9rxYEtgo5qScVTWJB1cxUJ2rSL33v
PehBI3kx0AbQ1CgD6Rhepsapc39N6xi/YDj+XU0D2VXUd8Qmxx/MK5yBN5zWjO/9
UK277G9D55OqRgiEK+ufqAFtTx8gQOVY0eCdBkr/ToO3EWaxgvpZ1OA/yHPyps9i
DiSlmgmXpRp+Grpr8FxDaZKt48+7e8L4ZeiFU4JtHG6gwHJWufT3+69lvF6mq1/a
lb441g+cGas2OWK4px7b30mL4rK0vwh7lDlxymSS1w3lokS1hmuCe9EaShowO5Hc
LOsKXmC3dwfimJksT65UIPcSpkTp+Nk7MmL0yRDayKw/9q4snWPd8DnghDPJmCJg
W816EWMTcJkXlSkMACp6An6+SW10oFHzoQlaclBEi+dXrlnEFi3e+l2vL0LyaNT5
VZfBol9MOO/qpVhiIO5J6X2NM5e6RXAP7bOo4+02/7ARtaaSyFRJqK+GkEQQfU6k
uIeF7thLEv78rvnJoH13pVKkxJuEA3JWSFmYWzHvj6KhVXdq1nO5b8W0qPtjKTN2
T3jvZ7rHqXjkLn+erpFExALfFKkBBmrvImZNll83Z/FvIZ7dda997k4JqrTASQym
JyCFhWoczk8JLPJS0YUT5hqvbmBrNG+qCDNOcPD0bg142RiMN0+mzxoKjujP2M4y
A7+fJGZCd+knJFhkpbNYfJEVC1GxFD1fawv95pkXpMlrklBBtuL1InUMTEVAAAv9
2SwV3xSEUtPTcnhvlDaMmn7nPUZk/ll9EeMqxaNSwWT2RmcYu2g44cxN3UR/cV48
oTPLgGkWwmz8FLpz5nd/PTrcGxyK2MdG+ow7NtiNxgNjiE5iYQtErX+bgWFj8dTy
KAkSK09egGpb2v0KPWqzf9U47WoxgFPHWZuDbg2WOs/xgp54ADuiMVpiL/3E4LAK
91rJkJvgYVIuo2jWN0H6CYZilO2Ch3CyPJDQQ2Dkv+Rr1glLfb04cFKIerKJibaQ
NgSd7SBfX+DCpnVbTN1025+9HN/jEs3PHMqN2P7cYAjOzaH+Kvlk7IHEC/t2jAqe
RJ8VY7LNm2JCMmmr88JGm+SIwk4jT0nHdl7FQYUCt2lwjp4ATRShStNUe+dOLnKu
j9a2aqSzjucJKgkhBsIuwCbXdy+sq6Ksur7QZ9lx7IzO5PFkWDU+q+27MfpQNKfY
ZFK9VdhTlfhsnOV2zoiP2iHDYP/s7NtyiWJwLPGdE4O82YayZLdR9D1zs+chg23z
WOxHeGJOWWTF19CYzCNCnXhiT4+KJCosqrdClkKWdvKsdOEohiOSXKsL64P014Cl
R3qxbprC4nFMX1Pjvghc2OtTGeaeNj9DIRvRWLEvGlMRkaf37I87Oh0PRBZsmXdk
HO/R/Te6b+raZV/iGnNYjNNAJHJzRZyiNhkH3BlHHglxv0T8adyzXp0KA/vWWOfA
JGAIUs3gKp7nxqEima14TThSzIFY01hhOGttrPOg+8UASseXPdYy6DAsSZeTHDZA
h35DpY/n6EdNW4mkPPC8i3H2JCh1ZLu/PqJJiAl19QNLeddE1A8mss2B6XSYZW0B
DUhP9aPcSXC0j76sPN9JMgsBR9xn4gGxC+1AX3EXl6DdELU6+LIG9yU9ZcfpifxO
Ta7RepAeuzfkT/sDttN6k12YgMBHD//tK4xctWDuLpCe3h/qucfttlvtnebyu1t0
JHuHkdcg8Y0235qjb1rmnJXx9y8JtObapaoCeYiQULXYqzYzofT7mW0TsmpHoMA+
daGpd98Lqp44MwlkSIT4mRCfJfp5zGeRXyfwtQjaZaZkcLbNEMKLSNavlIU1+49g
Bt7zmitEjYhHduGWMHukWayZJPpENwFnvW/ZPFDztUJB+BRJI7hy0M9fxapdMZ6X
D66pw3Cc870bnsN2MWvNbBu1Z4BJfsTJfGd7XE5TA6LiJTGKMTSQ5cNg8+4y3hDm
VhlERxjSiVOaua8aU5ObcTom28ebhOhzTaKL8Db1pEEUeF+pu2vSUZ0pvrKmuj/G
FT3J0YGlnDGo/3UIBRdm+VRe7whSDdAyxjItqwK3fFHXokemKXD5M+ZBDqtC+oRw
6U0LhdPiQ4BzeO8nxECFAoSgq6LWxK+Lfxf4gc9XQpKIsgjhmKZUTXoSCfK4R3/C
SX6/aUJuZXTOj2d0KBdgWE8Odv3Oey72cMNZ4J6HdgWBZoXsbwxHAPpXtnMHcqv5
y37Zs+uzUtoZruYBs7o8Y2Q6zbrSaYH6JojLUIZPvKQQ/SqNQsqQ8NYKbULs5Psu
zVB5sW/2hn9JpFozpsK8t/sCIlEfAgREFZgnHyeiOV5Lx1hXFxrbmt6hy4cSt5qt
5EKO98mgyUGOZTIMvjxPM6cFhoHNv3fZJ0HwxOXD0VWyiJpZ5Sl6kiAjjonW35wZ
TbJ+8vQxQUdm89Lk/fFY5a9ucsPghoMrBSmrsd3fkXdqcpguJ8H4DJnAcYhSAujT
iGFZJ8d4Ekdp7niAdBaDb4KqR6RP0/LLX2Y51j1bPTh2EgHHEnBaBROz5vjrcnb/
63coXe7RiAfAZ+JWV9eaTP7aGl8R5YgXFLGFFhS6xy+jGl4yXwkHa9oUlsO6mg/8
sy0xSBCK4qxzrWWgySqxbzJt2rqf98NigAmF27PH/3xHCg7dbfJQGGICjKdWGEjr
8ZJuQ6kdc5losVJ5C5UcJrQyz09+3D1GeqxYS4OC3NhqqnO+EcU9pqf9vFL5qieO
S8YRUkrr9WLe3aFaUZdNtYBzn23140HLV0jJ8yTJAOhhwgWvRvJpYJFKUT+Df8Re
vM0+Pp9pW59v69cbwXZmkXVSPlsLH5KMPJp1gOzRrok3nDdIXpylAc+qMn62op+/
SaRIRAZTnqQ3hgfrgl8xBp4pcZuZooXfLAlEFMtmSkxMb5dqrjA7SUF18T/hgypA
U8LNNZ5qhg5cGyookbf/0ZdY4PQx9eonEgYPCQ2d+5eju/5SwnwonJzlIyMWYxLi
2G5GuS5ZLmrBVbaWEw0V7LZxi9D8MmbPKbFvlB7z+msfnuJKt01BmP2pL8TJtw9S
6Of8gEFgrvYD5LEXm7idOjQ7eipopRBKd3ypHeLFJcezd+7oI9W9NNTsn8J7seMD
jLG6ty8AitS5y+jZVrehurxtAwTXgEk9tA/VxaURSvcPwPJO7V24nsr826JXQysl
gHpQ8YIoKtbuzALWitY+zHsPH9QnN3xG1ZTACM2N8ddSiCrhxKNl43tJjQoLW57c
rvZ+dAa+kh1Pa08UzQLZj+RlHWnaEXX314zdGFJidXrPfgDpjM19RUPtGxysPjWM
mpIwbVX3jq4A7zP/vPrny5dBxarwkLiAyTOJElHIVwfXsSJA20eaeyCIcQHMfC/m
J8SluO9uCk+dN18dm6zXvzXY8tAIElkmnRxo59dAsdVJ6E+v8PJWiu6CYoLP+1P3
aPPfNmFOglzZHe68YVfhxcoQSKWGJ9fbIXk0tkex/GHQkyjkefebUZPu8ez3OR3O
K7qmfzoZqEhuMm2zv9zn5CAY/YFRNcxkDUPTkg6T7AMRTS/kPQaWeiPh1lrK6WYY
XfCauNBVz+vyCt8iVIB6QwjWglbs5rgT+zKWXykadLggKg+RHhY/yJ8h1b0mjlsb
sJFDc3Hj34eo3XcTvUoJgoyP/77TgZFtRpkNheOqKvShRPG6NiIoNzSJZtVnKlIx
/uSqeTaJCEQk8W5WY+O3dCkfjmlHJ9v6dEAO8eXcGJEIJfAcyz/pkbl6O88/joKe
uD7nbLjSBCXCA1tAMZxIwSkv6WOwE5GWylfFvONBjL+SNjWbQkb4tMY+/as+67tC
/43rKwlmaLY+Gne2I2KNtXXKrLYDeCSGMnulobVtt2Xoe6NnwofJL8ieQ04H6qcX
GtWrs4GGm/ksC6/HnO393ZIYs7Td7KQKQMy1k2mFfGEIqDdYelzynHQNYFu9+tL3
bxLsOdylNBGgm2tBqMZfBTht0pwdNCXiCdQlXJNn6NTOWeSEYqgbeXS6WYVWdpQp
1bDCH4de19j5uzBesM9/3FvxKcCDmCwU+DBeW8q6tURRQA8RcaKqNi663A/4UntP
AdpPY5rypQxUcn2UbaEWJFqNcP6tmlPyQGGdH41dBIOSlrzTTaiRfgeafILIZiDr
XBKYctmkmxzF3WyJ3lKZeWvvPfikcOGuqphxJM/2nIUyXnYDH9a7UEN6Vqr6VfdL
TTExprrZrEAgETW9lu0DMt9lTvUliLQsZTGS0TNV82Jy1JYDOn+mlcpiSNHu+oQV
I4H4ykOHLW4KLRBvDx1X/YDSILE0VAsdhOTkjdOVva0Y2H+BVQ2kLpZB/iN/ijfW
ueOs22INOiRMsNANJ1reFGTm1z4BxGpU3IEGwiHpZmrh4nwFVohG7tflaNcDPl6v
PV0sQ3Pq4flPEvWEm3I7SN59Q4+1uyWuszG6WVISyIO11uxcqZniAfTr7LhKPY3t
DfTbenbQIlQzBJHJa3eDRWYjtitbN9uOyM0f9pvnJeUTFIjkgY9gSjfsod78cU3w
mNmNm9cAO89yfqXdZGSWtgk7nt+i+KT8IjGRSOEQ1+sgAZ/mDSQwkO4x5qgA4OeE
IBPB5N/aAYse1e7QedHQjcPUEQe5L6CXB8S2DIGIkGAXIT3BSknreQd+Pbmuqbtl
WQ8vwKT4k+Iz2kYtm4hYWZlniJu08eTPF3V3X63yJqUMClp6tOF6AMm74nmlia1z
5IqlQYz3F5X8mOnL2EZAy0byW4tfSRoZGOw57XcrCCnHB7tBs8BPVH5zzWeo0OwK
chmu5xv+OxmfhC6Bg6MaRpqoe2lpx6YukUlyr7IG2hqjjCqMOlzG0jTVFYp19zs2
wZbzshQ9q1u1wWtpuLbJQdILGGQEVxeaOxWtVP1TT24Qa6zER8g1UC5J0+x98l9L
mvWyXK5MmrlcntTFiv3pkBjkYYFjUhlBKQdo97qPJExnn0ORP+t9naNPvqV+iGLG
RoUO3oBIPM6kYzyHmEVbfLR/FmC49HMQuEEkGV0KHX6gEQlA6HbWI4o9pVnQQZs7
/P4ft4vav8XrpJSwFaBryUFUneRFdmx6h/+CdNnsfvf0ZCBX4J6GluHgzrHWaSHf
bG1htHg8WrAeoc4zhwTRYaOm/7sC1weIgV/vp3Xp7RgcJsC92bbjYT9rTR8GfycX
Ic9j1NJMoOMt4tlRFYWezq1oPZeUZM5uNS5l0bC4eQ6KzZV1jqKJRl34/tRo9+LB
xlh3EwMzZLg787k9RFEyxfT1H8cLfVgcFSv9FofYwhW4bChPNwfpomTiZNasA85n
HFJ0pB26mMRFiPNqsTeGGFEw0POKEQlFe0xjX+tLKd5WeWBpM4I4VT8227Q3iVjT
Iy+mvoMLR+grFObJ8gtr6M6XEi7qhe8fQo7dZVK+6HYUZN6KLB6qG+IVyOWeocLi
f9F4JYmgw+xZREVEu/2PLk5UGsworK9eyWafmBIjxdVkTjZyiqZbiEQQf1xdG2+E
TrikuEE+NbWH7P+259sVnKoTIzOS7uX9aT4y14iWdN8cjZWpGbkYxhWyvbJAKxsg
9V+kvBYF66SZUmYqyRHRpuM7SJTkKCyRgGZPBGYYKBKpMMcoZnZtlSB+NAM4gRPe
Y8qeOxvdbSzpiw3Ojxhdy92rilDyQPq2Rj67Y15pos1BqTPsN8NupeCmQjqcAzxK
7OLIEO82ljVMxC7eQCJrRhtNATcNXJ6U/RrcSfVWU1SDqu+jp6K6CYYXHrlrh9DX
ZPpjoZ5//WU8w8odWGoYzyq5oe9SBU1VUu/pgh1F+c/UL63T36PPXeNHS6M6mTPa
IFQKsZPw4US5dyfu4OAsmYFX07V89G3WXwsEld/t8pxK7zyFM7n3QqEHry60eWVk
1fS7GgNMZDsT8WE9VGPEiLZz3W9NIeg9MfmKzWt5q3qBoaxp3i+cRZ48cRr/Agt+
9n5LiMoEAlmfyXgT6zSbWrx3zfHG4PBI3rnS8/yc6XE7FVYEptOuHaKDkdLH430a
XULeo4BRs29ia5DykFR3+pDRvw4LtOQd/nka3q4mZp1znK8NPnVmmu9aldMQmTpK
+jZ5r8I69b4rRCB6XNmAUQWgF837SRssxY3jqQAluDJuGpISs/w3Sz54v9WF7CRY
3dhap/T4jPdZuQWw3uw63rzDHK636OfleVRafPivhm7wobr/yhrO4KcGfdBqwTjU
cVkTMyAO2uRdZaz5udxOJ7/BEMgA/gA0QtVoUNvYfhL0DXfwrD+AUhBsGnqS/ocC
j5nPSWJDxoDprNB8anVN4TAUjJ88iM+bzMQVObwSwoi71/RlYLC3sv98aSuJZwMG
gracbujsjjbImpCgEe5G+z71la5of34OcUuQ2ExzeEwG7ixCdsfumfhYSkBEKq8J
C/buRVlwnJYFXcyhtQDLHaObsxg9eofWbk37PtcaQe3GMfN104B/yRwyCLHDtUsv
3ON49S826V8dlmixvvzaLlhRQvR+U0SgedjfyElLhscnFwhbjZwJsxe5uVLXZUHX
J/5oitpqMRqCo4cDkaNNInhxuBIcsD9F7P2opIxWKkFDd0yykq6xQ3VL11mEFyz+
T+6qtmQe8pYdaWxUnZ3AMzF6H/zfqvUwHmoz4H0iOouM9gqSNrrtqoIE9zueNt/Z
PDPwHwcmsB7hBjkkDz+3Fh7Yku0kw0GgPuS/XP0wsCnLcQKM58SK6FTkFV2XyUz/
pJxRi4D+47pQwdJJ3t9joBSwfYUz74E24Dd14S9DcL57ftf5P3IpChPCBVxuwq6h
/Jzi+iGFbAhGz/+Me9V08tjBC3rSgmsFzroNEYokZWMvAhHkptoPEgnr3z09r01g
TugMrbPXQBLC3e5D4KshCqA/7wjbgC3BOV1SocOmnkoeD4YsO13mV+0gwhTua9oZ
3g94Ca2TntiWprOH2Wx41HTm/6C/jadZ6F6CG+5tJdA/hSUuuk1VmeTAPjwuQQOF
7wZpF+rV7F3aXf3EQryZUtohz6Yw7XEftPoHU6yfYIZe4QDnKEWWlbx0AJU+cpqM
Uf6Fg0Bs34EIN9fmos4cmXYwZGN2/I9EChTFw8hNfw1rYEw0Qd9i6O2J58m35B1D
tZbxfMtoalqJ0mns6u0UhZ0RvIB0lczXrf4VRAVAn7fizy+wdq4JfY+9L52U5KIm
EbfafTGznNUveK2c5bYE2Olty91XclcPlS8A8QwWYJLuKBki3HCbJP/Qv5Pgv68Y
5+vCiGRZ5jQEoWXYOY3ZSUcUdIM/HOwaR+SneyRp8h4KkCyl37MVFQLbH5WXpmk9
o9Q0t+tRzl9G1UZlce09wMjBQFjU/u9hDPvNN5IY+7IzIWbrJ6/cHY5UxHCl8wmJ
00UZBSU+f3yR3jbWtkVGh4jYNVFAQTtaVfaCv8LxfZfZR6MZ6ATOePR7L02rZKAc
Pb9QjXvKbDfhIIH4h2VvSazbv+7yOSp/sfSGOJ+DhhPZYsy+Y50qoiriC2JgAKXV
FynvfPS/+dl6SqfcbVBeped72s9EP6F9SlH5XVuUq+0n6o6bCA4OhMc4l5SR886t
jMJysP22wr+tllS6qL8FoRBrPTy5Csg361xFUQwHXLupuL4VJJCmVZ1cRzbSWCyv
BgkAkg0E0Hv7MkVuK4aKiGT8KYYFespX95VWGqOAx+KAF3lXaOf4IUkkrx6uxvZs
7aZwojiepRpodZBR5DJbzZ3NeCFsciZhZNQM/cRNFapbtfJqLi0M3oe3FXd4+LQM
yZB7DLNb/uH21OX51+8G65R22tHRfMAJHxfg1frGVw7kpiHRvbK7E5efywcN+67Q
WNn4e0LsXMT1olKS/gK4bK/SGlAF9WjssnPpsaB9dqjbFIPiEq+FuMmYZlMbnRLr
EyFAZs1RtxDEdC7mWlDHNErRtBlxJ++1+YUbGJsAjYmjpLQTXVh5nroQs4QE3U4X
WIlhGnwhVBXjvG7mBp7JFGmNrrK2nE6IYIfG0y5+dF13+J3SCb/x+eNCbXGX7L8x
NYBiwnGnO5xy6blkuDe00Sa5QObSvbifp0g/+3uivh1+9mfATMLh+7rcNG1noEVb
Vh2VvybI+RwxgtQJelZ1Xe7mb3HDSu6w9qubaIwWMiGvVMVCF2Eic8ufCh67X1iT
AGypbKwPpFUMMLE4N3RCfjZWz8dslvQNSN1zHGoHDujN/UXRurd8ZG1B0/q/VInH
YeGUw0hxzQ1/niJWkwEO9ZM593uSp7zWt83GCPny3UBOBtwXjOb0HgqeQBsohlqD
s3Gsoz067SmujyaK0dCMYTxLMP7LClmkJFiuAIKAIGH6AmL5F6vBJGE7RyZFI1mq
4xRESjo8ikmVJksK1aYqQFQ8Umf66E9RauefXaVvZMnfToq5INgIx23pXVi6HGZa
LPntGMQFLWZH3V0SY8oKqYmPvKuBiTRkb1vw6QMwE0clzjcNoBtkROeil75PwQa+
fl//J5k4OC3zuJgyDqxvFGc1Dz2uY7Uq77nj11EGlAO9CBMQL8YKQUR724+oZbUX
S4jGclXwToYhfU/qKf9vH+dvn/Sp/kzQNJ7bBXFW03tf2iQPbFnfwX1mZcX2iB3e
1FrCds6TnB1aGDM7z2ODnmnW1GDAPfrk3GDnul8IANW29ba+XVuThRfQbJOEa880
Oybzg9pui0EKz0HD9saeaFoiAn1ZZJHabDy66JrDlUDieJUx8kpWLG1Mo6NY0zI8
mE9XKkNe5V/VGRbMGsm97WmYb50vCwBfRgNcwqWgAc1o+eqbu1PJukDu27RM82v5
9dCUbpoUCDTvlIOf3TNGK6iH48g2zdqwnLtjgLF9tR/teF95Gq9hEiJDm5bJXpCh
mA0XnuOFFn7w26SAWIaLgwbliycK9F0SujjbUNQWOb9PZ3uh0G5GpAHUo0wCGFDM
Jh96QfRhPdWZbTVRXOtukXsFzqkWnF6Mv+ixkeaIyt2JNLBVazmbcBdoVKmYNP+F
RSzsru9ib61IzaNR9W2S+WgHS5o3xic3/D1iNWMYmQIaxHkQswIruGIjhCAEjQyR
YDgIgoHgPF2yXvoKEspb/gkqmt1TWkq/u5w/2hIB6pb8RKZgIt9cgvQ3xyZAauNs
peKQ9vnGieVZEdcQ5qmiL6j3CtW1bkeKrnSyJzn/kKj5RiDopsvU3GoPVd0vNjO5
DbedfkwClTTRXqemrfqoYchDxyCfVzWA+f2rnmYfvDc2+zq61ydpykVG3/tpbjBy
eaXP+ZPgJvfXOuRGkg/pugsdXF3v1TIiM06HgSl4LK1Pxs4ee+4yF9wsQiixoyR0
CSrjlldpze1uUtRCJY8o36qbPLUtoiY3HLyeK3TZypmyMjsqbDnAgVz7hUuJvi+5
f2a3aePEFFp/UDzC1eo5jna0KJiamjmsS/IvMLDEWO2AMhIaroGqzWt17wzNifIp
qmyte16crZdONbnJtcpe1zfHPX7XCzcK8RH94DPzBl+/CgueOSMIcaibTj6kAeS8
DwAYBgFekL98YPDFYVZfDkvs4h3sOV0MQJJClW1WKWU7KQan99vhSJHRAw/t2691
ML7HOBwjeRU6y0uJKjLQnLjKucyFuqcUx+AupLXm8nbqq193qR8KerNjPMYFzSNb
1pAStiaMFt2e8QFUrn9PenaBcEkYYUW0I7//jV+TKMzxaM5QpliSdFiFZ0bnRPoh
HfSUngGMOgi2Dq0EWe3JcHcLNaghOR327PZNYx4NH0UcsSNyJaWsfl/UibKCc/Tl
CyuPiRSVGhIU3UGd5J438AYGaAcF6fwu5+BZrue5xecMcG9vZUBjjShnT3d6hl8i
ez7JwSlGlK0hEkvK4gdJTVxuhJ8zyUmN7j8YzmQo2tYnIM0mwiIKYNrSuVzuzJB+
2t/JpdPqmVFB7u5WHCNXsjB0nATCi7EbywuLKmpvvgCil90YOCRoZ/ccLF0JUnP2
y3P9+LVveU3T+TlBcw6/UyHdU10z7c4OhxhNHdRzMlkf++CiCMyO77RpFOUaGOh6
FnJhg5kXOTJy8TynMqEBnmF3WIbXgr25Zy3qctflAq+QX3lEDznArYj2MdSatXGc
K1xeT6YHv87iaexNhz41kgkdmf3PxAri/rTmnTByDNc1bMk/PQ954Tv2IFMXR3w1
nL1mOB6t0zIG+hr15nPkOL+Tqeq9r/p+LMKT+Zq4e5cNoXDLkrK6Q+8g6BfPMSfg
xZ6iEmslOGzTPjZ50VLElSc7F7LjBj3nVeQDdYNfUHXRUClBsa56y3zxkA93zNt1
4JBSxwdLhcVlKnYn7deJKEbMBIrQxlPJkYnjSv3ZxpNom/KgkV5Y2bIB0dp3k6mf
VIT3sIBWoTXcrbLfbwYoG2RHzGNm9Ea3P6piecHfl9eIrcG02VJ15EwfoKzML2Pk
RDcJtKLaR42LLMdoa+1O/mknwU3dpA4gNcq0Cc9hIeXOR3x9ugLeBvSLPIn2xyRv
DGiwFZNnUnF4oDfKzMLkP1B+W6eUP/Al6Zyk9nEdEKWMrRj7rqZjTN5UZTBsYM9A
RhCYwgVv5BrbX33uOyimxmKke7BWSFY1oGSjT68hVpL+4RavLPhu7KLtB2t5q4Ai
Ay0dYhui1AGkQWdjHsHfJwCdzK7wP7jWNfRqEEm3fwHNrJI/u4dCRoBT22RtQLo+
AtDHe9hfFYbd109UOaYPWfwRY/uHPjK4CvLmtk7Xz9f52eKpf41i/MuQRbbvLeRz
8jNlvnecdKdjff6w3UMvm2CBMB4zNhrv4OOmuHswKbwGqk7CXCRd4Lw2/v89gP16
g62r3l7aSjYocC6jjjpe6rbLYmvMgJzpvytZWC/TLFBURuW5Dll1wEWUW9gotTZl
2nC/zh5tUVouIpjssAcEYyn6UlkQhht5cXkagH9p9alpIsn4NxS8rLMmTY5NnknY
xsAsf2R1IfZIIBTTbzpHdi2u0xmAlX3U4YTA3DBPWJmFdWM6Q82StOmq/SE6mjUW
WSH764nq0d2rc7Xi4FCKJ71QYlkWCPlxaFDu8ZBexhCVM0NmY13j05eh4S/vs3xP
WpbYLWdY6sYxSbcQ30sI/lMHBPcOgtnPkAiK/o4PUNOLxm00mrIQIEHATo1XoCi3
6wpFxRz3swygV1Y+fzEmY6zuQVBDxD1SbhI3fKnU6GgnYFf776PQS9KX+EVjKO1b
se+CfI+CvfnRkxS1JIeWao5OrZMREgpg/1dCGE4noRhB3m/XnI6LbJ3xw/qJCOnr
cz6bx7nGwpGCsBxWYUW5RKO8G5QsYL6iY38x7mmxDveLckMrxGWtUyZrJ+A/KHWw
lHJvcJbHjMcDnFa1oJA4bPb5IQYbr6Fka+yrxU/nh2DX26G/jgdQqjv/SKJ28xvW
2l5gRYSthhcRe4QlkAIwu3wGb7mz6oP1VllWEZNZvIbHQeoRIX41aG1iA6B9w1y6
fKQlCn2fpGAnNL8Dt7Zr6IK4yCXUDfvUEAtjkqw89jwtS5JCcxnmHSdmVLEkJD3X
iU4PcH0z6AdD8jnfqiFefkhbhZmgym0MSdW9vHaOJKJ3oicIdi2WH0CYIKB9dtqZ
fDoMUNM6eUSPj1iaUlrE5q8K+C8Mosv2t3oSXK6QkNQ6FMkKUo2eQn3S4SgQ8unT
8uTCEDZ+Q5KALUcjg4TYnvO3o4NrZQtvsBlm3EHRFAOtayPC5+50zCLeZJupBd5C
X84vjT+wqxlAUIwoZSJomsyywnKJVEeHUSMn9LimX5F54L7F/B35PCt+4Hvw2qbQ
O1e3mTHqgzPzLRS+PZX5COTMBzDWeEMUonZzgqksD2klFb6pEOQ3E+ZAyC7wtaer
9ow85jmAjnRTZyX3jFEYjIOZaA1ItAYJOl8mDKM4Z9SDoK+jAJkt9IlwHLTxqVEk
bPrOodlQf93/o5fSgQLyvOl2H/RbeWvj9mdO6LKQMY6ShdLf78lcK8oGOVbJNBJp
ZEqtXDijxKd9kdSXDjf5mjnbKYnpHka5ljeVsq1c5Agg6SC1GBAthoHs28R26/53
5g2MMnW2iEtLT7hvI8dQO9jSP2sBFu/MI6ZSnJq8DpnqjOOsmhNJJ4nG+agk4SM+
0VopJ6hX1iBKTunyPWfaNdFHch1+T0bMbeDvGZVMal/2DCg/MpdxdjbzC46ExYmz
LvLyEHki9VW+gO+TKyT1nSHZEE3jFL9emFYUJBXthiQ1SFjrfAUr8huz0C7YTnhD
F/BXGKbhjU5almM+TZ6tx+uoLZPca1Ptq8kfAM0Yy9wvQ/2f85z2zMA5O2340LUy
LP2W5kWDhVs8EZkFX/8hS892AViGzNSINSw9AL3IVezkPpR14/K6hzJz199FnE1q
eayYmWxAwvziOy6JrZI6TKKkVSDD/YkihfCLR7lCchD+/5i9Qd1ZMfnHJ/5Rdey4
9BZEIVhmvu99FS2VRP7wTsMZ2zWGjOwpkLZUFEg/Yry2QixOVSGCddZaRsHmeIF0
SV78+9lTXkSolaOuctmnezS4evT+mvoVtliERH0mdMEP9mkfsXwYVtiIiMe9Ua80
fQNBYMz5jC3PO1Yuw9f7y+XZwN4cW3gtCqV2JIIRw1h9CuKtE+qMW3N0cwf7TsBW
O4f9Td4t4p3f7Z3qnZUbeRLtOlymL4EZQY2+Fx8JE6KgXqrJXxGJ0TWl7yx3wP2H
F2scexojIopt93acfxrk7s490q5RPw/9ZWqPwJCdD4BydissnS+I46jpvrUhNtBT
d+Wko4fbRat4g1pmlf8J2h8/aHKDFMP2fC2Y6lnEVA4jKRUU1x6u+a+4kHZWIv1/
FIaA54I7robmZ5eZvV7epNJoAkaJU3R7i84euwB9L/2ydgsapNApROuNs3C9dgiL
zcu6Dj3WRHwJG8/IcNbQRIczodmcEAV1uUlFCO8srAcjJgcgs+m3WWQkcu6gb+S5
6Tobus4RhnQYyppzElDydFWSRkmpmnwWl14+AdgJh9ylc9/TI9xUAa7KqR1PPAkt
HayBGvwEXnbfcRPBAkdlTwoJkD1gV6SoE2FAOgmk/Po9JJMw+JQS5qEVfwxlomJK
13XrX5SZ+D9bnzYt+oDvsvGEyMi2c21jzylUYAWrtSLABNOsemRvkobPJ9DgSvlF
T+6mDdBNNWBgPdj4TNKNF0XNlMXJcUaG4Ipc23uoy85zDJJmhnwkBQ+5mEMaeQIt
xvSc2yvqjRW69bKolzIH+ZV/lynCx8PYpx57R7iz5IFvtMfNv1MLK9H4finXdrfl
OrYbkcIp0p1uL5tgDCd1cfBU0BDRsNUDn1lpgbVSeKG2kCPkYYW5t5Eoc769PalN
Gs1s1QBDul40gASclNJ9DPfRBqOVP/SRZPenFvYvNuYie4svgUD3RYN7PoE6wnDu
7tdeM7TtcoebpkwfGWoiqH1ApfHGYjUlMpiXmbN4zbe9tAWST3BnamO93n2wUgG6
VUtNcuTPcDn6g+23Bd5LpUO9nG9c5ynPihHAwWv6uBE4Ws/Od8MJccFc3UdqcK2N
MsxeeuK/RP7EADsrx3sgpE6O2wBgU2Jxk77t1/agAI6p8bVTgOeIiBBpnfMwvZCv
OEgf8edkrHtQSM4qBll3fIcj8RW7AqzfkHbjH0AY+gZMa8FTl1KfzQ2v755nq/Nm
tu5sRyn5TCFed8fSwfQufzsRpssn5JPsTjt+eFYC3nO1GZzyguAD2K/Ur4lsczt3
MH9NOTT+ggr1R58Jr1X4m/Y64FdEkFRtw6+WbhnhujZnIjX2gg2AWo4WrkbFzNvb
XED4gtMhbJMeM+I7n3EV09hsQ+mCyw65qFcVrrnTvsJzuqGP+rLzVeweVKt42tH2
hwh3vV7qSCOPlHJMPpaE/Oe97Kc+sJlCTu7zb9MZzvH5RyFDQv0PxNv1XpCf9PhF
V6pgky4HaOo6U+OjlNvEKP8I1Am0p0ESxihjWJAZHJmb3kAKWkZrF9daRb+CgvHC
PMpBoocaalfPxiEB0Y9+5vuiDfWYwQ5+2iUXfdCNczhv1b/9oVAQiV6kUjzj/8BV
5hyZhja/WbGMI62TqJ0PjYduv714HCDHeMEqUr/NVLX/4WWeg7dKifleGvNRuYP8
rSdy3I9KvwrU4gcc7W77S7TtIqhTwSsI3LNXaY5926kaTUyRGKciR1CK7v2d6mOW
5d6wZX7W5nB/i96UQjFGCAYtuOLuO5HRQGfb24Y3DpeifNWjRoFnuTgf9Di301QG
QK6ZV/He+K3dWioscYS44aHbXhzBmOgEdg8fiqDWKS3WM4VJoXmQBhiFBbm22Dfl
p1SeJW1eaYGG2qbBdciDJhJs6+RayA/T58xqprDj2r4+z34B+E7bVH4pMYMVByXI
yll0Ve5FV0dHUaP3XFOy7DfUGPMQGW63UoS4fsylgoCr9a45Vd13iH0YaFkpneIc
RgJa8zKbC4Mc9FaE1JlQ7q2xEs1GkfkPttmFY7anF1eazza58yT6zMvjyS5PW6+I
BYHHXesys+qW33NkqRwJNZ9DcR3t1biVknJ906fH5ytfw94lgMTZLx14ypPuGVnT
/Cb87W33DJDFE5NjFfm/+EroM6kHrJXAVYX7o6QUFpY59BOhGNVEuEda6IKU9prZ
vZfjtnpsxUBbt2Tw+f+twL4Yr4Ig7d+XnLf8WcUluRXlMlJe+80Rl8oIWY5yJERh
OVh8DjDJ7hebevAxuatRs4gnijgbRa2bDxZD3Abkca9HmDX7l8E4K7nMtNZMeO3c
wn7+Su5dYVUPRFZ/zbyR08cqVF/g9ZcgqtFkdFj0vW70yTwo7oi0qzoejWMzTSic
SX/lgUBIVdMZ7sbQFoZN/p/t9NwNnOof2bmUj8ByBihk9XhVmoPDe0jtyA0pzPVm
P1ghdiXfWMcf+0bzIXEquOXpMLAJ9FCAUJM/9M/+I5mAfLAnRPdBzO8F26N3YvOx
ZJe3U0XpBtQ7QEHvl4g3xZN3e4kY008bUgjjFuflVcY1Xv92KSUg43IB29YnO1w6
qcUz2+ffCeS0mrM1Cg8YbOetGxvvZRf5aYAX1mbS8AWhRgdmk9P6Dt214fzQm8cA
gAzvYRYr6n0KTiGbY7RFiEqX7ThDq9S0NUWiZvVg4fExMRCxrnm8LsxQRY5uaTKm
DMkeF0MIuLV4vy3YoFUWkUJcnGFiSUe/jbZ4KCtCOV8Jufe74J2KBVCcdNe/v8Y7
HtY+Q3MyvOKUVpO8/oYjkZETjV44jhtVDbdu/9fP9kvQ5XIoDV3Os4xbueVqKKPG
qwymLroHy+59Zm3DVVks1Xe2gSmzBxvJqZV6GMTVu2110Sx290iESJJAfeO5UvN5
y7gKMcBNeQS5hKKb6aksfK2du6f6KvTxEDuSuuJDWMFC9OEyykUjYgRmwljTH5IJ
Vk16okKvhCqkc/amrcuHRWq9PmB5Iovciq5Dy/cQOSdFJF0TIszPscqK14sB6EEy
jqT32VLukSZf1ahYNFK18q6OYyVP3p4VGTjRYvCRUGZ6+mX2N03CHEPsy89UJT8j
nM5tdtTGFuWbMkcB3B7jhhKsjw+ATTIQdKXeOIxT/8jwfqQzGRjXKbOpMN5xoItA
FlqzjflSYdxDg+4umXjcRZAuoRMwhjNsvQi9XR3hMBWghp+K7fwOEtupOGccjzgy
w2Fg4+ht7LeadGGvhyHjphewK3i4HMcQhUnTEsbbFY/Dvli4e+Xot90XqD6kib0/
U0FSSxAYbCAdQAeBwh7u32+A6MIRci8JERotfACP8fCVomTQnHBV29ndQ8Ux4D4Y
A6Pfi8/J/hj7YE8mBwo2wTSVippMHxBb6sDVXguKyRa2i2gRHGkBDjHpKRyleRtC
jcaqXN7tpjOwNaHGwoYpsmqIwv/DxTucz/mViMjP1JfCjVWWF6LEMGpvpqj1eJiI
DLFMYarHubPEvKRFUmw2BgOCD/aU3mSfUvaFAiUB6fBczIYSG31wOgQcb7m6vO6q
CI5udvKyRcN3Hxk8CD5BCk4p6idEb5ARMfyM+WLFAAiPN7oKY/v1J5kxy7FKOZ+/
e10o/UW3ONMA1d+m3LWV0Xw5b9k1rJxNJ1k2ppWOvTT8TlfGURdmzhUyheQD7hrX
xAbC2xJjkBPNXDFnStxSN60UkkFP3H4LBybir0xxImH3PoNjADvlXR2pjcA4aVhB
MheIeFmFuBLXVMSKKUlUOrj/ljSzxNPGzdk75TlqY4DJ9X5ZOIcbxWXJmQYjK8pi
hGLYMXSzkgYml/4Q6k1NxOXly9WTVIIcaauE8VKpoa9I1pno56++e80L2z8R3npv
ASobaTaoN/6+5+DR4C454LBbzf/06ohzvixCT6ZXiFBX0ADrciXxHuwdwSML4hti
KyQk0Ysp3GPbjNrWNloRJzng3CjdzVaGJ43HlCJD4mWGr5iFHgO20s97vQbxru/o
frlf/TLu5QRTcu0sdclzsOwrn9kWosv73t3/etFFdPO9JkIDay0OClaRsfZJIr4l
eC0Kn8XyjzqqaTwv4mCWPf2CFDHlgE2emdUdmlIsSOXCwM+/10KmMaot6Blq1YT+
NqYlqECqwjJV2ZuXBPOj7+guMOGNCwCuLiHSv8UO2rzLnRFzBB4adD9AyA5uSIgw
phVkEjq/LMK9l/vfeD8CH7B9CfW1D2akvJJ6p0EIlf3Mvx8ZCwPEvAvk/qku/1eE
4GvxeqFEkhSuxj+EbyPg5War6YHEXAUdd3uvBBI+t+7NHncLxBAm8fe9CkRmx38R
bYVFhXEGn4vi/dyWl5NzU1mG9sVqEgMJYzP2XAjjN98Ve/cT3XA6g7EAlV1QeJim
G39jj21Bd9DfB09Diu1nGc+GtTjq69xH8fGZGKml1PFJTPR0vyMFh9a9QA7l6IBX
j9a6vsxZbLrvkwSIIW/40zHkN7pLn5OMjnShkEQzOzOkq9Wk6yVYOkm2nNDP01Fu
s1/RZ8/B5uOhxn/twQ2ZC9GRZAxI83HGevXZLs82X22+ZgdzC3oOvhCrV2g24Vm/
+k1jYCjouss+Rm+wu9u+2TB3CP/5qARnMrcutzMKmEPfIJ/1xNGe30o7Ko1HziQl
Dnv2F+3KmDivqPAcR2RsoUi7sAh65abkxuh6LIOUFuU929MamQVUUaUuUuQIeqzy
6IKhku1Jui4k4tbKuFbcNqr66TuIf+IdWToqD0rAGbPcQWYPIZrYPJ29rylLpDbD
tRyfbrpGAXJnmPWDEWtT1k+SRFIJhyD42q0NIU5GQbAzgq7cXOk064eAlPMq0UKp
vtZlUGLoD6xA9aDN2jz14jclbjdKe7AcOPjoYq/9Kf1rRugVCn1awTRumLHk7j8m
1GCu86CHvuWgsLhHnCZ2kKbU4Eodoxa/lT3cPBfquvUjjbYhHqEGsoNP97ieCix1
wj0pF7KATPM6GtAojUL5VfGpVazmCmKBNn/TDnIFv6KZka2AcE8AvH0dVQAIqB9Y
SiQhUBMFzPLnK9p3hsZqGBBXHwfVfSoBdFKVXA6asWUZlyWcA2AZmpE0xoMYHAA2
F8znUk0J04PHlUfEc5gcLtbIXso7c00un9CVGlR6pLGSYBSTbyBQsvk9TXBva5SI
D5jedLxxqa0Sik0O+Ulwy8CiaACcjtg5wD6UeOOjYvoan0aDBy9APY/4L+7hvfMJ
zwRl8P44mI9TpIJu7RlehWx+EzT4QspLdMmZn1ze9CZVefAE39r3IFyNW49Y9vLJ
pRSiJthe8P+t6R+LefUEmxtj8N/JUtJP6A1GXgIvFsVUderJMLwKZUDPNB1TslFX
qnq8V0n0bZITjhxmjgT7NUXL5OyMn+EdO6ab7QEIe5pM0c44LgSst5exNCW/KO5l
Iv/KNEfsMa547shiIXMeJaEWAdxpmM7JYAo+Qay0Wxv/+joHltZuVfWInM39P0O5
swB8ObPlwenE5Kl3kb3fEOfz3S0Ik8c2VVArJg7t6YqI+aHD/5Gk2wjcovM7TCNj
amM8pX3dSZBRZDnmJbC/YZCpMrhhs9QF/WeFAYvp+LZ43h2osz6WTfBwHhWd779J
io1jSyTLz5Cmtw59hZCkFbxdIpDwGxNCwOTxWTv+jiX1MiDcyxITrUM32NVbUXUn
zZXIMZlk8aNE44jkc0rU2jf1uM1uiSYxCLfbvw/gtdfYH6nDHeNNKv6LH97nWBiQ
yncanyvngrsU6u3Hc++cgpkxiFpAv7TKfS1mwwRRqac702LGeTEMdO6akzI4lUw5
QNvL33lz+Gw95oqIJXHKyXSGF1Myd18zVq5vgIx/VCx1XWd99Todlkxr1oOQbAVf
oya3Mk4q15HzpVYQ1YtCI5l+IYrIW43gTMod3Gua+Y3orsUM6KuOtkWUJ91JzLqx
`pragma protect end_protected
