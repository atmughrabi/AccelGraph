// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hEaP/FqCdnF505PXlWunVnKz56+7IKgqW99hG1zGvAa1o+rDYwV4t6OF4FY6fMdv
ISHPC+HQC6G4B9X/1GtFhlxtiIOMBgW1Ru71ZyqjIJkVeerkAj+upltN5Aa8Z+Eb
SvqOViLepnYO0DsreoRY3CpB+951QuCDYoJxGzoZThI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8560)
zOwWaKyF3xWYhclI3uCXJ1c4AMXTvMpS3Uv1Y4n0E6aKX8LGk+JeuK4G3xlU61cw
obYYLV1yc9T8AESjMrW1FUnXfZikyug3/csraWTfzI9u4xAJdsZEX2AHHtpnpxcB
NuGvY+IDAGHuBYo5H0dsHXM28pc80UxvpH3CWSBj43LVvf1hEIIyqCY5Ez1WQAVW
eRmwa8/TOpkJYgkdomN29hbG/IGyTFSxCTxrTMKT3jlwSMrgWClYc3sJ7mAyEk+R
esTKyukinSG1pICB2I27hLgaGPlMto+RDCDIzerdafWnbIhaWEWawhQj/qxHCBYZ
h5OZOKVi4c7Pn839RyE8gCoJWgbxnfhICUF/NJ1A1ZWP3et8lopLwCj1dGQIBZPX
tJSFqEhkTQK0zO1063FKLc6zksSYJhXrn4DIPWAveTnpwb6R/FiRosTXp4BwOe1t
IsUu8TjPGVJZDK0urQGrA25bOekM97RQIX2W0Vkf3WxgxSUaXhnVONhPh4TGoxw+
82JbjHFUTEzQHAcALUIQxVtpnNhR9qBegX9riI0wdRQAAyIrJAzowgKmh6WtcIBh
51uu0tGzLiYvIOfTs6+Z9RMIEeIdOFXK3nar62MdrO7hr4NjvYUEOfutM5dW8wBI
eEwKtodKv8X6Jd9Et65FccLV1eWGI6tVerymNyhvgw/ASUTmFaSyaL3Ar6kCy/Lp
GEWubT/9Zd8ZSwuZSPWuZDPrB7GZ5kmNEpMkAhQbgYVelBnj3lXADQTFZKVguThX
yIzO+3sVNvmLFC48nlmFHlny88HIObITRsfJ1w6IimOdSBypcrnVWqNax/0sZKd3
bGRYegV/XFGc6L2grr3IQbWTbeqBtAcItCOLsz+JWbWwzFsYRWzBvTB5H5p6z4+L
6uoFPXsVlbjt6MbbwVTOd0jiMl0Y4OawfizXuV1eTq4DK3qFsIVQA1FQvgPwiMsL
/Hw+prcHBWqpXj38jNCNLxFN47Ocn9LYS4RPdO3wAI+QpwJAb34OJLE2o9XlI5ki
CVSXvHpFVfpmmgvf1keHbLsXeGO4XwIEvWWk+86aZcRSF6Bux2BRSpACs77rCEuY
3AQ/X+1gw5bpDQMweZWTQc+S5oIepzMpsARSdR3/D/Mrow6CTTefMzghXeeqXlPh
rQc3Gxwy/Z91yso0GsIXWhrS5C0kVukXAFJZeQB2wgB3yYKDBJqjChiJ7g+JSkPC
1Ai4kvbm95B+v+PijujfnMnhPAnSRykGKImPPI1udVucjhYB9qCddB3p+o8mJXWC
othplbW1O0E01BNRPnArpKui7VzPd0bsJE7RSQEmuTg7uOhaI2+nAuvE2TbtLnad
QQlDXf4inPLqKqmtI05VUjLZeCb+qhVzf6cFhygMTE1JfrnhaSK+xo7h7UmnF+oF
v9G32caZIuUglxR221kfgJSfuVfOaCcqoy6aghjK/SBfF0lRW6yVheYdaLeiMw4P
4fg/tPB+4JDz/eKSTthWQ6vnzb7T2chI1k4Xs871lkjQY6E08biJ1db1ar/5BAgP
mUBSzIw/Ath0yjAJ+nJSvLt+FXbQRGCpxq9GZqtZmxZLTA94I9DLZSUys6dFGoIH
IKOUIzMi2NYuDjiocHmze8juz45F5pZNiSy42zvJCRVXyO/uQ2Ww64Qmk3TNOPLq
nwnbhhHIiWdYxTZX0Sj4j/ph2M7xKU5ItPgoS2NmrtHmzMZiKcH3ZobMZlrK0gm+
2jy3+bh3wNO4+xRUH+qabhI3wT94rCUfsreuABNs/uXn09j87a6XPrgbuZhYpVSk
nL6AkwFJpX592+UU17ySHeiD9GaB5YTAnViaZJ+Bcz89LnDZP6RyGL3cxt7xUA95
rBoYqgUzwLNY8X0Phd/pqsmRnveLDb2+3ABnBfn+tMQrluMtcmOWNAs8sAAfLlQd
cVx6IhSP2io0SlTxPbu/gkAAJK6KDBWwMVb1wgu+oINmllXnVRpHqxfEf5soWD/d
9CvhAPUYbmsECKS/erVpgXJ1DMcveVXaY/s7VISB/mg0Zdrd/KELNF+U4IOttzj4
xH+rRLCnH68wiSqTp472sexP7DhQhRPOR4Rd9iqh3bkmXKlgcdEpjJRSiih01awt
yifsy6WRcJFFungTy/h3KmrMYpGhY8My3bNpV2bDrGlYcjCLCdGJdBsxYXdrnXBl
6dcwvfwtRPECNssmw6kvd3XiBUvEGsisRnkbvzAS7A6srpqdbW/WVGXqs02j5ri5
YoXI81Q8rCdobVJhgzfqevL/35XsKzqhukx9Zl0aOcR1VdkFUr6RR4Mbu6zN32GG
SV9jEMucEKH8d944/d0C1/WJGCaG3rpigKaz0bGyfHBUk21G0HxxtOomzXxKZlPK
MI+t1aC/XD2/Y0doupEoodwL9iaK6sm9jPYkCHc1nJfROVscJG8gRg/rRtBk3Yh8
fskRS8/yGlYpTZ2xMclVd9oHyiigU1usedlSqq8lawkP8koyQJgizZ5l2lIUwdqZ
tesR5+J9BZfYd/m6NCNaFYpKSvrNDZ7czjp3SXVB+yOVwFoztSoqWL3HOI89hLjF
XjwKIaHdaM5z1mS8MGW1HC1oLXsaWYt0SWzM+plVkJMwNtjBZVk1ShVB3r+o7buV
pui56j+dz5HFDbyO2PahAHyN1Zs4pJjeJeperLqm6O4GJqkzqw1DRIDkd/y8nFiN
Xgoczg9ehClaWyXAu5GA4wUU0WX+A8oe9XOmpEey/RV7vAX+S+hlcrSIlKlVAEV1
KDC+k/RC45Q7vLJ8nyc+gzxZLEbE3L28uXfWqcy97XSNWIBca0xbrS7MGPZFsV4R
cQqUHeE8OcA0l8XGb70QQEzgKdoramKK5q+trg130yKM9sxuSz19VUasPhdLmRqo
eEXXQupISQ+rGDnNBrvk1K2r14/RyTERQDnDzPeUNGRGMRFCVZISB//qa3UtjiZQ
eKRQdPiajNm44ikxfIRgtuztP55NKdHPb43jKjRSrZG1cQn0SrVtfdYE/QnzDx8t
BmwENC80YHKoZiexaQsPvmbc/144yuG9CBqvfIrvSYfTSnec6xWtJKgXbfaTYV/c
RxBPUyZozemGBAD+cnnoJjSFbw4DtEJvjKQFnFiz0YGAI4YYB89P+UWNDBo492aE
YQPvbIPsRJGoOEACLN/oeBxS0xqvNRF3oc8oiX+jDKxj2cpkxsV8cc1X+/cifN/H
E7csNzEbO0A/0U/1xvICHh8ppsqw1Wy2XT1wS/heK+1q18tXVrbc+fRfhCLnDg16
dkxnTZaAEGmtc/t+3NKZrz6lNnnR5zAJuuPhHXJqRRsJwwg8/DInC8u9mx92Ejfo
OqX9+7L8LDiOgw34LDnYh/e1i/O1/L1ZASpk+h1m03GgWad06uMck8NEDuXMOlEG
PalBgmUt70DnMqPWS6upgsLPfsgF/Glvul3fM14XAsKLqOAQ/fEx4GALATr45tqf
gTJOUZ55hTqHbU+7Ic94V/YY8SEKPv/J7eqbGXedXgdwvN6h72iX6fjKLrVua84/
hw2Zjn++m3gt8Sn9RiE5DBIIkJSIjfPpP3Isn4Ys2iCCMSaTMOG8JtJyOy1yMfAV
GCfabSMAidqEo/9pzG87C29J55FdVyy5jTklDS1BxI6Y1CrDu54rm1aBxO22CD3C
a9jnOdmTUHUM0gH/CcFNQ2E6ooz6sNs+rB9gogjuCexEZrPf36s1J5SkTb/liAsF
ccbVlgiNhoHdpFywS5H9LBXazFwLY+68PRmaHkdVVcwHs+zErd5aDyAhkFJbTS/X
VTSGw0/GEEtZ3nvDj0aH8JnPpomXhxpmiksN+iJ2Nh8PM7XeF19QnktHjq9E5Jtk
pehVwjWpz7G1sWq4zmVyL8zJDNq4WU6sv0ALfaJo/PPZgU8VFw1kv6Yq/X+a5J7N
o+vpuTpBBAfiYT0gb+wJuEzlEWxWlULzxIBJDhEPkQA/EH2yHIZutNcJtxEjO+CZ
YfzUzcjGaLakh2dK/O70hEU6/Rj84nH4QpDmWjTq+EOGjCfu1f+Ey1dGP21bC5VM
zx28UCQW+EkVuEeMAJ0asqXs3rQOsevZNMYCAca6khQNl7CSnc/cV3ZNHJxKgHXM
YAGrGR6VowF034EVEmWVJDSodagCJdtefqMire2WhrHUp3e+bjDLxMeZZBZVieiw
hfJbkNOQLeUayMMaMu1KhkShVS5JqDTfaq1ADrcdIbsnRnXYvXuiRIaYjKUYyzvL
xMn1poJ/PN+XC2SATJfZAhZKtyKgPemPEM6lQNdb42jijk/71+tl4Strv74xjhi2
775JYcMU2ZfIA64eMXyLtJ2isPmlbbOfxtiHkAYhffoRwRlaOBOEWu4NvkWOZy0o
ETIM7z7aAfkCHdAOePYkAUUJ6HbI/jpcWmqIiCsMNY2grJ7b7nZ21BG3h6ItnUwW
7qy+c9y1aax4EdrKBWHBmA84VW6J5Az6+vcFQsLh2Iq/ftHGLqRgkKLxxThd9AKi
mPHSLjwKB1xfpuIrFLfI+tL0Ku71vZ/Fjk7eR9AP31QipW7DhHoGfVlrGt+IgZdZ
sYto/HpG12JkEfQ3yp5CmenJtfcgR2Z2RBthWd94sjm4nvuCyijLnaTtJXiEimRS
w9ElltIa/e3UogbpbMdIM3dUmYQ1o+lDc9q2gO8ZytcAwE2UmUzyRXAyLWIRALV/
E/DUGiK5MJB8hD+vwF39qzdrvkwFgBRkKcf6kkjmCodrzhrwOkfKxn0Tfc075ava
mgS4OB0w0fZqREaITBhYNHRuW1NeKOGvTSm/05duDKiJJ92nqdP6nmxRKA1dRwoB
8ZBnUbdZ7Sl/s5GdWP4iVB9wATyTbOX4WW0QlrTKXsMksWQv6DHQU5+DZ1G7FlUd
mZN0pZXeIRLIW+6FhKdaj+62A6eJl2bQ5g+TXBplZ0Vfqas8TmSgBo1wDEQx/OIP
7suJEw0w0seAH6hBZQfqQwd97ficKBpf/OFPfUvpBXWuHyXzReWyUD4//LzDL8fP
RwrZvk3woeqmdG01HshuFR5UGzV4w9iKDWdpOhAnati+6MDXiQ11TNgb+zVSGpW8
EopjXaQWNKxtAxDv91c3uNLYGju2NqfXrl1KVHHF6BbXIS3ByctkhJUqNqG298kt
PzpRAMHuRYospN28HL0vP8WQCakFPWG9WzFU72GChyLReC3k1jAiwaDDMO6M8m9S
fyUgQ6YxdLhS4jRYiTNfH5I7Fjm/H4zs1UIiJi2UzcrB5TSczVZalYs0e+iOFjUp
3nCPDAx39qG+q25XMi/qZInrV9ShLUOVsIAGMOV4qzASpR3/hXXMxaC7BC58FVg0
Sy6NNPD7Z9cmKbSfIaGEXqHcjDwatRdKVDL09oArRS5z5ORpsbUMYO1s9SxgqMFw
JyNTnH3BwdClqNTgchZeSOyAvL3hfZCm/8MvVUFJYXaUT3f8Ov5zvCvzeFqSqqel
eFbYznD0TXYBmmvHEJg3H5DITl+TPygUCHOu8TlzgmdgkndhLmOmq614Mw8p+GK1
1aBUx8j5kVROTGwskspmW9kkTXABKkQCLumCxsNiuzObUOPfsXe8SJa2Nu6dFaqO
xxdu5K4eSeSD8K7tusHarezFJz5k57DX1ExA0WqVWiq+o5NZyHDMDuGxaLN7vuX/
SE5eAY8eC1iAAXH62c1f0lf6Ef75oFELARp93DO4wzN9Ks4Ew6jOUQO/ud7hQjG/
jr4NOiM7XdaAKV376zRwyV3QWQ+H5HlPvKDn5H5CtR5mVFDXqBXJboCYxaF8ozGd
CaUIsfLEZWH++bHApbINbuMFZA6yuT9cYmocCBINQd97WbkFhjvN3yIqwINIOfz+
8EcBRdWXApB4m92xc5DOndisTlbZhDp6XVykMiO2ruoGJYvWBcp9OWlPpW7MD9ET
KMmhotvByVxsfnJrLo14o+igvY6qWLf3AbGwx72TnHaDTAF22HCm2YGwgB/o0ROJ
oWsEiY3p/+IkJ1UkWSpVIkXf2CMcD5TJpjy1LMPhKPVqrgpBwFP0z2Gtg4ya2xQN
+gqBEdLOl1IIdycmZJge0JIhs+jx+BuCt5rsY+X/kbJgSfGbMz3+licLAMRAROOn
IlePO2/z934NDQoX4xuwpE6g0KjhOEOKLOb5I2+YyHdmxX25qHz9WzfEPIHtEMm7
76ERlzHyrvZpE1yTu446hS89+ko7LwFX7WdbrRAxlq4Mo1uaSEQsZc05iA7LEY9Z
rBv47jrFoEXMULLOVU5ekM4v0pcscuhHpQax+WvKAtjIqzEBil7ijBdg1a5iy5Qa
KdpO9xiyNQQ4CNgAwBH53vm4v6l74YU8qZqbN3aX5LfDjYbXz18OxmlXMqriYzGT
aaidm6jajpAJTgabCj3eiY7SMAaXXMA7xCwIp7hcTY9wVYikNyXfxJ41ODV9ucK8
uIF84U5d6rBYv5zAivWLPLR21OCZM0OMJoNN0MLQNPZBPqnCMnpvO23r8C3QFO6P
ngMEuD9+aM7ruHXG9ybMO2GOfA3oJ2DgmgbnVDH19FE2ksrGEszJK/A0NeXwaUdN
hhKVemOnxI5Ozj+Nk/JHefBVqQCfJn1+Sdp5k0ilMmBqIpaAUVZOx4o47MtkAi21
Bj6dECDitdwIFGCV129T/UcXNMxve0On1QQjvB5tGRktzHXtbZzP6rGEEgRq6FKT
GRhc848YZ47RgPPtC69Mc0mKTftZ0BwLwMqrpWnuNLSAe9bXdmDT52pX34az3DwF
3GB4mB7nc70bO/srqN4SM9LG+rZOcDWNVe6qNL5wSk4g4qRzKr0exEKKWEfxOAvA
O6yqeAyWKHvkli8z77+FZNT9eGAi+bxA3SD6bM6Vs47A/r3ozB7a8FopyynPIu1j
itMdbDKSv1Gv3tjQOtlDMa0jYrBVsYBdvELJgIjxq0pVC7OZcph/tw6PaomH08ne
DPFMd8sBe+h/gaRJcd+N6c4m8O47u7QNVoYi83gibZYGp29FE8+R/6wRvpSdI0f3
6XIw+z4ZVn0xApLuoRNyA6qb3Lfdq0xbRppLCyjenj2w4SMQrBcV/XQKEBwcmYb+
Q1dwlgDIDgPDpg7SFuWd/TFvzGZwqnTG9/0p6s5AbtGKaN7bQn7XKae7gYkVRbbL
OyZ2YyLhO8l3Gn4eDJIGWb8P8EzUE0xlajlMzHXZhOW5VbxfeDFF+NOhkcMlze/S
uCuWYWaM/cmTZGsoThtYaynUIqS16RoOKgVmJQdjKpmllC2Vk0+Cnueu9Q4otJ5j
pr+wv2X9VYDbBnP7NIQTp62MzwNs4+sh6Fklf2IYZ5VF8fq6vbQcANRXXi4AUKjS
fgav9aViKMbOtizI2CCwGEgM9+7GpKbzVcWwcZyD/otFQay6J/n6Cqbf6BMxhPcn
Bj4CnIbMO6JFb1O641RSbwqER4QIcLdPWt46iP3wly0JEbFFAtQe9sTulGzJw1g9
Wpz7so7iPjPeHDt2Th2/r4MCbU5nDQcPqVOrpqbT1YwnATvDtENiUHtpKQOg8mOK
Fk6dVrFRkM83ZoVPJdp5ojIhNFhL/V84T1yFaZpGxeWF4taQQkqbxPcxqnqpe62f
LLhlVBGjNs2eM3wGNcmqZSilBZrhgaubVUimwQYUyE/KfWUsE/pykBu9EHVeUHAb
0zGqDpe64UK+r7jlKixpxCmzcxSQnq48nfgM8/FJHXjs5J7lQW3CJPaKGqsyhGWK
8Zor8nVyWhyk6dWmK4j9heheQt1b6X7Yc1RTuiwJwz7nOKFsvex4+eS11qlbvK3v
fRO2GmJJHzQdwTM0zS37fxzdwhyRAWw0jKJvVR2cVKx1h96qPCoWeE3VOi+80Jl4
tNDVukX2kpZuWdnSlTGng3I2bRKJ+a7DJivasUQPq9NuV+EvjTTnsnfup76Juc1v
lDayyfsevJSgJoaau+mwXylaKwIrtmf5hHzMaSvKRNNEZ/pJGspJwgBGB1SQ3jIw
aD8ovL4X9/gVtH0BHTaxcyPudEIAqikW9ctvwF5TMXrYuV5/veQOMux+mgF9/A7P
Yh85TnrqrIHPLL05OMFi44dtqwYB+fIHumlhUEo7EP/Riuh0DCEaGObDSXczJtcD
RbkcNQheJ1Y4CLLfXRQbZ6gsyjBp7hpYYwD3x85mvkbx1nppF97zzo+vqsRzaE2x
t4b8FhFLqDXkB1K+l7ZfNreULoXCtfoSdPcNOlk2SiFYXKVtlVpMt1Z0VeMs0n51
saSPyxuQB/X85Akra1yS8rRu0Z3gvj9zn5+NgC0ZDx4PcZiUR70091S9T9Gxfylt
MInIPjlbdGYf1mWysaPdj3I8MN21T85IbhrUutBGgkMDm/jS6EkajkD9P+hbQ30V
paM1Nojru+lwQjNjq3IALeKGHwbg7Y2AkesCPjCxtK0NfvixsAM6Hv9wSsu3s/he
9SmlsmQGS6NVhni0aIXPvUyb+kx3WtOCgJJCq5Ji9gcd2UzenQXWE6d9OhUmmOge
ExGEkmhWaLgxib8u9kFXcQgETzVM86kBKK0lpofn0I5yFSHzU+sdqlnkIE5XH2lx
5NQw3ev17pG2OQeUr/nCHGmMALSVp5MGZ/uTknKodArkOSu712Ou2c02TyYAG8RI
dTeuIR9+VmFnJWtvxbvE5zOfYVHUorCz5pzce1B1KNQwe3WWtYru/bslpzkrsJvC
ee8S/D/sSlBiJA/RU721Z8myH5/x5RrhwSpU2kz2+BGufdTWtxZudHtsSXFf9sRn
JG6uHYCXrLo8xrgkgpsGqAldUqStsBJRaSFGK7J11VSymuj5DELTJNpbiCM+e7CV
XC0k/FCn+oqSiDsNKdAv3R3hcYoAcxKUME3iAUxEId+Zi+kDqgxQ6JRfGAZJr8aY
XHbnQwEMM0fU7kA0u2XrRqb/bk8zxCvfcNmnF1I8LmIRfpYQMVz8z+796+zKaX1g
9b1zSCXL3Ulb9QAAL5d5onp0IuEzO78JeMrm5g8Hw1ZyoLGrS1t3GhgVY1I8nmto
a5ePbFq6xT8re0mRMDnqnMgeNE0QwyFDtPRzC7c6TV3Wiiwfq/XS3Jrn69CnumYp
urlwMwgGQss87DEjyDbThyHTPUq7sa9rgYGvQXvgqJsKfMYMsgBy46vZRCbCanWt
UxFtvLI2ry6T9GYUN9urqldXAMQVIZ8gCH0WHAAtdNK2CJJ+J613QM07HT2cYaKy
exu0JYeG9AfC5kf2JZBxdcg+epLDQ01Sgc+XNDluAMepFSB1QotmJv9klosrzMUw
3BXvs+ULk3t3YmifOBpPhbAfywbecguZHijhRGXP3vxSsdhlJ+Pym4IwxKNXavXM
+O+x8athI+v3RHnk2PtQogWz0XOZEpU8g1r+vt4Q88p0WChuKofPaZqdv/JwWl+2
nQGzOCsc+eJjmS1VG/3ZsOzC8x+y1ED4a1k4biemD1eGx9CmdVIrGd14I6wGdpX0
qc/cuiF0Uh4uVgGjxepVSIYZFcbM7KfHFpDENr26nUPEwgo1svrDyl9/hC/i4Znf
MDTjmiK3bETzyKfKanNjK0Ul8XZHpr5BJCA2sRicTQTdEUGn+95C27F4VSo8ahj9
xLEwjS2gBWmEMIX/rQLhVyBYW8yPe3os3vkKnkaGGETvRrEXreU86TOpsm5nKPni
kaVrl6PBImnNr/t9u7Ab6tKTZAgkO7HiNcpbk+Y7ZFEr/juHYBCTRBtQ06S/md/5
yVxYbnhRw26X9e6aR71KY361r6Ht4eQfXDDmWuHLmZ8KTwO/hd4x4QDxQw4+x+W9
1RMg9rX7SX6IKoHWMzNBX0w2PUJT/TQaW9VBjalizDTw4xVB1NKH33uwakth2cN6
TmDX2RAIYxDyynUHfysv9JMYhQATpyT7sGpfz4Wx2gJTW9sxwOWB7gsi3/3f2IB6
5OTvjRBQxPTzsZ0oqSx3xz27yjcEZhLSUfe5IuFA70xzlwIuI1yLwMZghgaNAXBc
y+yBZit9nEjuEs/p1R+ftQAoB8rUjI2bp7euoKOOqLhBDOYRPOdjwtuUhad9n2+B
nr4hIrLhjb9+IKr1AxYmp5dn0s4lTOFVoHxC64kfbDqGvPoWgFO5529wJrVD6uQM
ggqGjCpQUUtFUmsbQDpCNBNjQJsNOnDHJdaxL2HHoSTTnabieaxfbenqx9SCQyfK
Jw16qqf/IusWymDjhTL4l0byqyg4lcQNeznhUdffjQhUy+nm5scUvJluHzd84b5L
DYMxG5Kih+O0Icw0cpwe+oHIb9ZzFiakCsxg4fOHHG2NwkJYDeJONYr7d8MKSYty
oA7dZtbv4/2EYEAeMyS+WQ/G78MElUmTBskqnJXaAYdGRA6WeATKYH8eyYswYljg
5j/RPd68WotbtScxAPN8LpX1cHawMNK3qO5+iuyL/go99oj+hIeD7Au87ibCbW2f
blO16pdbSi0yxRIT6My41UqsV5eghB90cU/sJo8qfH43+LkErc0w3+lpOvIxy1L5
IuZmVIuZBvVjJC2WWda4UbVPtzN9sycoek8STr0tad9XMkoRZvgy77XsOZ6wtFrX
EN0jeEArAeCckKhwoa/6bozar816/ewUUwtXDLIimhbYXfdstCs5xRum7tDejD0I
fw/grivKVcngaWt85+yF11OCib6QJfrAEBtCpY+qaftTQH2QCfrS+rNPHbHqvx3G
seFeGf+cbLNuARARnpFzwuPOSidkvmT8YPW6rSt8zP9Rrmhc3Y8AZo8TAjX5TmFf
hRZ3CevcUaPEI/dGl/HYrmYvYwatt8eTQCI873GUcZNWHY35ShNCSMh4RrkZUjSc
voalOZZFWyYmgVVF0oObyT7Bv3f8qqlBdnfb4R2oQmNwB4bNTMOCCWIXf1SBhQk8
ezyreD1nP0kVBJhv8072yDM57grZYgoi0E7qZ81EzO1PKwyFcPB+GVrquL8hJfFh
wsYO0P67P/Qi+/mnrk1S3/a+ywtPqbFgcCuAEVxvaRWKdp5VCz67B7XYW35bw0j4
a4o0HATTtKNZ0d8z19/gufrnf6a9xn9TNjjYDS1+xmrJn9ONLzRWiN0Vw3XzSYsl
1ZHjsxMV61ha1xBUeLgKeK8E98YnPNpfqCUVFSMIWPg4lM/rvD37CzQ/i1YmQpGL
iH8nhTHIq9KJ+10TEQgzYlY2biQAfKBurBE0kfMhxGx+mNJa6A9CWhs/Dwyzt3X5
LFV/LkhC/8Iw3bUis159tsIAUKLdGh2oLjm+Pd78D4cW3db7sbFtoqpCnd2fWdcW
dUIG1vubAZY63zhZjF7NBcyfToUS82LVm8T3/jYgYMCcaKTe5WwvSyQFw1jreRzE
Dv6epPhVMssTfI8g6dNvQIGcy226ZEUgwiOUeKdrkdX9xBEExi10xo3kcdIFsbEw
s72BZtXViqESQa0IHRN9zL6od8q8k/Y90R1xG9NczO2Q3aPu9dS6Q9C2P+pcqyGB
0FZ3s6mUB+GU7RPp38fEOQ==
`pragma protect end_protected
