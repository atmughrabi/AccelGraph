// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Qe0aXfq6oX3Q3GAK2pvVhiDWjc1nJN1RrU0w7DPaNY7AMa784Ele3HoG9MWxEbla
HI4PJppJdDTFfob+aTo2mo2xboH6o/JUKl05JwHB5eHeDpg9U1/pCLs4qD+sZtQW
aFwUhOM0mnZ7XH4viePRZwd6rHdp3m+4ZiLDXqEvIV8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 178432)
T3tQswWqtm5MZT2u/XxH1QnJIYu8fX4bf+a0DRntlDYN/ftDvBNKnHMcUN8c/oob
kUmyg5zcwyULu8bLFV9ACVpsLhmdXMBUYrxCph3fA0kLQa4fpIcLCzKtB6iPY+BP
E+1zEO6aJNDovtl+jKsUi0RNj+qVxGk78CoXOv3/rPbxCmxOfvbbcbXJgEMjcucK
3UN3u5ZRRjnartFd6Vr6GK8VmXoggObDPCF0OvmvJNYVP5nAOCG8VOFRs70JXgoK
8oMbo6DONGWaCRLuKk4DZ3j1QNOP6Dsvy7HrDqK8iFu8RE0QUUd7byckMBbSGtoa
QZOItgG8TgI5igAAEM61eD1xn/F/zf7HW67mt+IVIrw0T1mkZSBv4C5nYpH53JNW
Ez5cJotJY9qUE9LzLonAR8Y2Ow40g9i9ZDMSiWUbYaSUSY0OqoEMrh2a5wpzrrZj
3UR5sYJtGeEW5i7z5UjiTeGUz6+95Yy7+1CkVmPFXrO5RuTZQE2SPFe9nEsFGoeB
qx3AZkRCLe4lI9KEVmhStz0+JnrFxSZi1QnYdwMJhAa9eOFk6SokeQTvi/35OxZo
kU18+8e5Yp+WSaU1M9Ekwq6n5w4qHYoh6Iju8iOm4bAwj8YAurq4AnZoHDCzpaVs
5iIxRvcpl5LRiOn4Y5PhKp2khBuFz5T1VQ4aK4AUoh8iQN1YDpvLzOKNNAUcb2WK
muRyC+DRNg8NCd5mT2/XjbsLXvJbZ3wi0K+UsIjns/Ifvxc0GYD/LU1vAMAFwpVo
yx8Na+nDLPvNF4/73e9R86T6zV0Bz2F98syd6l1qjKgvTw8+YX3MzVm/+CFO5Vtl
h3GvEUIW4+ge/7Ye0vM/FlgpeauF7CWIPFdfNtOouYzNhOhYwU+MWAsnY8G7HjaN
olubuS3tkeuhDUHNp9VBTXFe1fE6kbT0xTtL+8tOOW8sFwnK/t/1C3/pve6MU62q
MuYxFWOqKssJOLqWpMvd+0y9EHyXbxs5ZZ584uioFsYC0a+hYbLDvQ0qXjGvg+KH
u8zJIFeQjrmDgy9rLNWRK9vkrlrHCYZfgfYi8brLLrKGrgS9mmLeqoF+1xFn4elI
GgJGGpxcUPjzGErQdtF5U2dhs+UG5cMHyES93/V920rLIWjIL8S3wWHOYBL/2KBs
dF2TQXoD7iuQyUwZ4Ky+t8qXAUHXxAqhRDzY8RnnU+wrsaM+2Dju9QpjHRaEAmmP
+ErZjcUGFfWmYUFqAO8dlrP5u2/+dmjQCwP6IK05ywgtE0l25pQaJbXL7eGGuLYo
ZRrWMLQpDDkWnSQwtk8m3zABb+BxcKwvE1BSk7UfyEu7o4na3fvAJKY5zzMwecQU
AEE3y8IK/qoiKUTpHDGnJZYkRs1PkG0XORKii/yuNKtsR2EWRTZjtVT8foGs2LZm
x2a5JqE9qISIEMhAOIPkW14GWw3BPfmZQ3irqc5ZGkQUSvWa1y2evAY30Oi6oziJ
uCCEX7UGt+ClP9V5FtBmTIip0cvqa8rvbr5tQm7FG9+vviX10b+s3XFKtgJjHlOQ
4vUpm3TP4ApZt2ePULySI5e2AWEzuz9Spvl08PNNIkpCk/N09rLv1xPZgtMztcSj
6jlIdAfIZe7I9k/U2MCsxaeMn51D9nHefFdWwYgieur/LXxvMvJDFnWTog602Pi+
VS6Zxxn9XmLaclP2oO40UT6nHH3sMKmE+qJ/ecRkHU8aYjdAuMMdYSiQsCKF8QIK
Wzi+XEFHtK86E9VTy7Ed1ETGYOrwzy6lWHQpXU8VDsGowqrfx3Kl/9g9CIbbRCWk
AN31053ZY1JLSkdwGvzzM69LnmxMfoAgE/vBEBH4pB6Yf0mf61zrZuGmIZYY62bU
r9FwzYOBhH1cUEfOXPr0EH2Y5F64wUvAxifWDFe00UCrnBFPomjE8RODlzNnRGd3
3cJ3qDbDhkLWEyokUSGjT6YxVu7CGo/JQA5Agv4RB7K98dGBkwrSocp8hnMWnY4e
T6H2WoOwzd7Gj2iEybDoZgXPVbtXJMVtNjk944RoLBvf/+vo2EN9e9cncdh1VJ7n
UAnYE2f6mJcBj2okXCWFsXrHfeBe9sArDgLjbuKj3lOtLzF8WMg6ZSEN1dVhTZ02
eF/9/ezktvZ0YIY0/gNkTUWQLPOpBWWsj+qiJYn0YVXJaF2lVric1mzQwbI149jh
E6qpVVXVvAAc6fXhTGn/9OumPyYS03E7/7/gl4JF3irhwCR2NRA2HQU5GOjohV3t
SMajhBXUrT5NrAah1YbWjJSTmPXYgZ1cSnK8qgfVI9BBtOrD/LzymiO9/dYjnRHX
uiDyuYQDAF5pC0SeuUUu7j7GHQkDwnBfYUsoIR6yHQzSBo/WeW3YBMletowSFAi9
Pic/MqKHsiBeaLLD7cn9AnmhLHh24P4oYnz14ZY6Gfo0IK+4bQCGEADEuJ5o1eRy
V13odG1AFrsUYFpwIOpqSqEWh8jmp+9ZfdAIgv5LL1buLvDGVlnIgesyUqEbLJoU
XYwV+ncgO6Cqb75H6MWuJK8dNbehS6gr0ECMN7tk7w3Myo1rIFqYYG6gEJO5fODY
vklA1EyI6tTG1E/lPFYIeAFQJpldGBSI04/jm6F7tcVAX9vyuOvX7LdvLS4sGCa2
ws6z1dXVLZ+26DqMWB33CK5dIpSnKOuhiD3CpZHKt7NWYsTmzVGrejj89SIiLptj
Se/+cmdiSoOkhWVOJR12y1azhWZPXHhOZoTCC2h25uHzOmPwBVHSBN8lxWxj0dQB
DKsOeW/2SgRsnU2Cvc9aH6KoOmcAkIYwMEsvfGHdZ1v6A5O3aVIXf6IZ5XycKyjS
R/BkCXLuj12taI1gqPz1diwbGoUcR9QAA3y7pWVNTXQUDhUaEl9m+MLW9wt/36if
fP2XGv2MASimiXtJm1OywAXlgKJyluUkAo7z/uGG19UN1af2AlTi8Lrl7WtH2n1i
BuVGPjOzmjuUT58RLrEInxb4j5a2DIZ/xREam3jqdfcgSE7NEvBwSvE5lpMgNHwW
gQDslVSSRbyYUE5YW60/iktQWYeePAI4x1hYU+Lp/kUBRGasMZYX4hGETiVzor3T
05YYNiw8NboEeFZq4pMjxU0UomiW8lSVYw11c2kqGQAEVDXTphav/h5EWt4ah2/R
F7MY0F7teRElkmDKIJY8ZVRH9QxbdcN4hIiU4ZCIIFZYwFw8t7A+vdTKEYz600mw
Wb66KBc2QyiXWgC/vgQB06GlbXotxlIV4cRqI2JOvIYX9y7+Izwzs09pI+PyUtI6
cn+hFsfIauLiRizU8zE9KLDUOvWaEV2hYF9rnazqH3B5ZNk2NTKq7IWqbwW99YSb
TaaNejwjz5JKWVeIwgZqLb6GadDIP+gB4KaaElsHDRdHO9RZCzLl3aE1KHwhzXjc
3eZMBOi/UrRClsDBHInmPXzTzjKt5UbWv5Jjh11x4HulBzkkG7e1a2OUaAVgMNQ0
9SDWIh7pzrDzvTRXioTc4HyFRRSa9i53OLbRvwAZYn78OvpxLySUXO5vP5DMLLan
7R873IW6QyUOA0RlkIXUdNOzqjMIP8U9AJdeTQ52hkeQ2EXnvFr5umi52cIIJ1tj
HGBfE0TXfPxj+GZ0E3cHaKnwrOC9h3fKjPNlKAGQZR9g95BNBFbk3tsTsz85/QXp
JEXP1HgIZ/SgydrsTI4O1D9alSjNq6TXvRvrxp3sraNBlcqxsgC8oEy2wLJjraWR
yUcWnU4OxvuWBAxcBgr8sT0U5VtF/LBx444J8F2lOk9PKpQvc8U6OU8F8mzWHbfq
jPZhivdt349Gi5kR6lNSCvc1z+jc2Q/upB603dPY3H5CbOT9xF2Pkr+nnLFG8c3m
NJRqTN7P02hhMc16ELXnrP1bURu7rIkY6buZa+otcg3KCL6qBjHC4Kga5Ef/AoAb
d7AK1cTytg4ncX1BZb98KJBfBsBUX8FTjXmdhE43yx4yTwfH5EKWoJAY8COXvxQN
Th+eTKl4PKF6jaCqVtpW9i4BLFIITxUbEcDjFfU+GNK1zRukGw0t6OdE40qhW+E9
0Yjrp1R4lOMESMlN+LcxkJt26MTFC89ipel8CY46qupvdnRC9oZN9QYIpGruDKkm
uAo3K5K4ScmFn4RVYZDcX+9wPYMpRaiwn9D3cChCYr0d885niUBPA44rxNI+w4Hn
i2o3HPOWdwzvRSZZ/Pm5Qm7aRph+7rDvajy6D7ceQjnsGy1hs4CixMcOhzgfPEQJ
aaVGNsrKfj9P+OHy7qnV+SRAkHpHBNrHeCM8HVcIVLtTuq7D+xo8/c9X0w1/XoZH
0frkQjDAGg98tlMUnycin8sxkXDEYISYOsEAGLhr3rBkqJXvVMH3WsQ458NHRfDU
8DZR7XA/cOVA/I0Vq+7RaW2Az1IvbVLtiIfPTMYtwYnQXd2TR+t+HoJYn8DVmOEV
EIKukCpHsB+KmI8uaT0+ak5yD+wRCRDnZjRBtRyhpGrSu9ewaVw6jylRhi5TUaac
jjLxN3f3OPsiMGYBuuGHdgY0ERNovPfg0q5h1ydaasoxpAMaAMyOwZVIJ9TC4lku
ib7l7LKa7yq0DA88L7hUTcCNC8Ta1Tzvp6VG61A8Kdt+XO0qvF2xGphw02DIJl/U
ndIM825xccwfNjgO6XmuDAHZu6zvUc9a+vUG68nk0DvTmVCzKEGOs3joYKzPdq0C
DbAA89tPrPf8Jd47xzPYa/nAXWNrROWs/6u70BAeffBoqTTqVNdetE2o6AeceByh
7pWED6d+Rq0GjUBYO23GmTmwI+CK8otgfodSiHsjcxNDURXSDykHWARNCPxWYeF4
bqeoV30xDhFtuL3JkuKnuicr7jvQStsN3126bmuL/AibRPcypLYaFlGYbeEQ2yC0
GrW6uxFX8Gy6BN2UwJOKAAp/AgRbEaVr7dC83QpVGOfowLbURckUmA1NcUQdl6CI
0EoTyPYOHt9HMIqU0W81RM3U0iE8ErVlKuzgjNn/4ArJfqnJl5tIMYej5P2wpXdX
kvrTzICjL5kCaT3i3nQ+3/S4c3A8dtepFyehqLi+nquGvf0quqDbUdZhSzdMRWYf
RwAsAViijSkuDwFTxHThWsUFCdJv8dEzkMV2OAuLPX46ID4tUBap0gl6SW1HjOzT
0Ci6BsQ4p3uspLnD7svsoPn1CQvC4Ex0ddCAbD2YNWdSUeiBS0i8kg1AOKHdiGQO
fJ5yGISLUeXHyRfDL4NDQqDAY6/DqoKunq7KbIKI5zPjiSICmq5DAdT8ECnK/bwa
kE2n9ERANm4jQmZ0TSVbemQq6sZdyIs3JwGCwwwMA+hFULCyU9lCbAohJpX06X+s
/NS1G0lMbfoN6ewL0bNeyGkEEiOkNqu7qQWMnKBM7skgdHtmPeG5b64PsLcTlzmn
S5/2rWJXii8929JB/HMzBlADd+KEx6q0p/LIVkZ7IInp+jI1arOP/RMiuTuLqc1o
AwJCbe4dIs3nH5LfqrG5isENxUv4ogj2Jbe/lv2EoyfhJwTm1zaXTGzTvTwqlID2
jLFl7DjRwzyi44HAZa+JWPYUQYkAd7DmLBFeiSC7Q4ZGatlT/cF6LIopfYsqlUda
SLQEf/lAAZSILcnP3ECd6ntJm8txm9KzYTx51AZBSysNZC6jJySSxyFuV8Os32/F
WkUClYvQxPxeU12ycnwtgofXSOAAuC6VgBIj3cFuPpaygnPbzFF+B6ehul5i5u8I
kCN/FPeLEizUtF5Zzm85faUzqLzM4zckByWXz2NNAxarMRpwMYcP17R/RFP6fBvK
0FwVry2xn4Qc37X3Co67l6xR8Uof9+KGe2TxPVIwiFtQ3OaeVphQv3JQJbY9Ez7k
hoi3Mkj0aSBR1mfsE7z28hH6uQq5iCZKCNtKN9zXrIqzoJs7rEJWlLGnnotQH5GW
MxowKUj6VqMi89PZA8LPgnCmIL0/icBk/8f5D7yn63gDdTjTnkpOofxQH+25nA8g
2yj7goTUkYKKJwQJ4CMwqiDRcMgbqKtRsjOGtoG7oFMiMlllorwTQxjksx4Cv6Jv
dMc0EjJwrFw6Gz5mgGpBuCGqfr4C4X9hc3qjlO89olEimvnEUdkQ/a2aWOOd5hKa
iSOZevnyl2ndUwtoZUW680XVco04Jg0rO4Y4H/Kv2lDEOXmFE3T9A2mWctS4hSNS
LBgrwvIwnKykZpcHmv9wu+7Hh9bBsL/DKn0YGVXw1VI8H+BV9kWXFtChZVAJB30s
4f40E4b6VdbJf3cvBUP2sG7j4XlFTyeOTLGHKRKSISz9F5tMaBoxQO/MuuWZ3UX3
n6xAjtTLd/cfOINRapBnprJotxyJ7phF9yY1eao8OowAsemvpCeY/3iSnAdN8xDW
9QMxy5BGDoAWHmZleGwupRD62790pQI9FQVxUsq9Y22pi1bbVMLDXKYgMgqBab59
Z6BMpZB9ZLQD2ndmtPeu5WaZ4Q+u7DktziwsQcpECIo9ZBmdQF8i0ZtPETYvjKby
mmtfyY689DimG/b229ThOUAfRtbt4lzvZ8XJXIvSbIQ9Na7xcsaB12AD6yMHdywz
Rpkalp7ZfybzpsABeO5DF1zrU3NXRAhKduI76cm1CmU5Mfq4yAI0HAvUvOtw070e
FSQ+CXM+sGKcrR7qxws1MuuRVGlcjEPDMNsG0Brlg792dB3Z6jh8QwwMmiZzcmuB
XK8yiehIibG9NlBonuU0hJ0ixhklgYCaASEmHo0lIOoAFgVq5cM8k/j4dd7NVSVc
+sDzxvJUGBCtrV8ErNIeYT5kM6KY6zX8jQIdt8yZPdJy0mDAVNJ6DaPaxsDxavbr
idtQpfhNOzTrePic+/b4ER1BoNgGIEw59fotUkB49CoHYvvnpEJyWEjbSi0L4BrI
xVYbNY6fR6LDl0cnNOdHlj8+cdce6zdGDYZNhNBMa36A5zXr+CEoTn3x9nMbN8xd
z5FLRljHiSRPHHv6Vy0wuzrdyfHMhHTA5VRbyeTgrVc10lAfR0ugUkry7SK6lyuy
du6jgi+RZeF2YUbRP9UyABuJnoGhXMkONwKap6gwYYDXjfFXi+mDGKrTssYqeddX
vr+EOh6ftHVtQ4UiSSAsbDO/fD9QRq9VkALEXZEa86dZ8qi7EFx2re3ygOVpx6D/
nnDL4iBoc97mnZRfpzohwVVdOuuxRbQ8qe/4BENqxqh6/M4xGME7ZL0r77rgv5TD
90KIOHqYqLTJL/C7KdRqSbGV2Om6W3oLiRD/SQdJD6vSQsd4Y9yHUm4BvwCBH3ko
tMKKGk9VFhO3fgsfLGBPz/OD1Mf12X1+i1sM6KOZ5M8jICAXSFm1+TO0GAhWlxfm
pKwk0SQC6tnQ3oDE5d/6r2xR3M3BmqGj+sKs4qMGP3Lz6JZCEJCrI7ev47g+dSv8
uo2fISXJF161tWbPSnQcH2SQI6RbJTZq9Mf1AqcjMc4tXFEYzGFFN704+07dkOMm
ldAdVphklic1Kv85opW6i82MXudHKFSXzyOLdXaUoBymqNtm5qBfaCSMUZ6ZXJWp
kHnSPnP+TXVnvhu1ktCKX6XYMzPieOdxPKAPK5o2FREmLYI3As5ZduxD7MyrmW/J
pjWQZwpcPm38p1y2TLL+V/IVUcP9Cej9OQNJdsNbpKbthvDB15p5ec4Efth25v1M
Amf5/iOsyeBBYPh4JdcXiNIj7vynouryjnUkfldvoJGBnwYoRQU4ZEk0pQEeedpG
NUM79nlGeijPAnjYxp4tWTVAgWQFK83BWULw9vqtz6Ru5U0RSeUxgHxT3pD38FT4
YB9DzkzIkaemWXBt70rtVTucsGKmrzoHu01WJj6r73FBjKLBgkqgGF0EaVVlsQrl
U/HkIUMdScbMfclJU0kT7prMKs109FV+HNoZMC7YKQNRxAgBHIlZTW2m4GJUZvex
kpciVkCCY1R8LTNOUussWpB5K4EuGJwGf6QfPsge4GtxIDabFcrVF+ene//VeX0S
pfziekX2DC2n1J+O8WZdn3SIKSQHnYNFzvp9uNS1VTwerO4QZ49x+V3y5dMWkdGg
IIs/veDD7pZvqIo32rGY0MAg6ZWJQmmXJOkkGPzoWf3FfmQ6GuQF/h2ZG1yib9Ep
3FA18Vlqd4V5LjuZAbqu0ZoKvq8hVbRYlnxN3lqAXk6NeVUp9k+vHDBaHhu363XY
hUWTXtDOd5bzNaHQCsnaGarbdW9Q0M7NY9BACrSmdwaSDdse1uMa52AGJzLd0Cuq
YgEr2FhcdflpCG0NkVXaj7J8TkYtPDEel+pe7NPMJrb0l3A6/8rizRlurmlfEppm
DqXyEwZrhZlXgzTZ79p3/EeIg8eTrnJMrCOlIHqPSj9pXsu7c9VU5TS5KZEPYuD3
NQs9wmWhqpy29QUJVHURMGK99RK5YzPMvCljE0O/vs3pu0WycvAYS+8EFgSR1sLq
rc/plR7WaXidizdOBxHclhbdBogxPLrVvgKiNIooqrg+Hma2Z1iQ2dnDVXRSb6AH
TtX339lEzd0m/bnWsIOi1r/1t85xIeN3pf+2HuLgmbQcEWE08fjUTjYkfEkuCtCW
pxWzW9CRMNjQ5aXdNiCnIqVFJbuNEfNZm50H2bhNAtlM/d9dQKaiyicNH0QMD73D
f9y2Rv636/74Mlrenen3/Gx464yOENxyWzYvoOhDdtb3j+tpCuciHi5rHCqvGEym
hExMiTwFVVo9uEPWbpB47ugjocaeS5L0roIrbG0JPn0cjXT5NSJdDPs7jw7ObNTP
LDdb4DKLXnUqRCBEcwN4TH10ch0m2iVN678t+IBlmIbq3M7BUL/j2ExpPnREiJft
+UvtOYiXOyuFZW8nv6AdQFcZij5Jlex+nyx9QhMeoA6g2xhiglc6WMSBru7Jqud/
xxNPPhxo1RCJ6SmyPQtdCPzpK9d5XLuhRHJEXJPVxOD0xXGXkSfHEFvzV1Vv8y0g
SKb1AKNmLvEAf2NaBEglTf7XpDJ6FiTpXMi98fMFpmu0hB1UPVBsGpHRHbgGauFZ
gsL9/WHeR1b/b2fUDUOQtD07JimhBYicPhwWzxKqBIMRjP1ja/LC0pXCTbcOg7jF
0mFhYhCatmiSpuKPb6MX47Yv0pCn8QJnvyQZwehCCCP2qBq4aFsBOq9UDbICdqnk
qebQqiF1BDM/4MGVOVRAkxR2m8sKjRygyIvrs0WcunvoZkqHbd3i1bB7S3I7RQX3
4iOYbvO+u6j4zoqwB+yHKtawu8ZL0F0bSHVIzCVsgZVh9Us2CJXKcrS5VjfKkLDs
eBl3ob8IvFidzLzEMK1BLZZQna4VuHyELxIuq5RmXMn3n3jnJw4QYVXHa1jx9hD3
FU0ahQ6UsWEasrHqfPcZvxaOLpB+MKkaEODK3q6dVKvvL8Y9BeiZxjklHMO9QVvw
SadoG9WM5WHUvT4dUP+z0K5KPzBv6fXuWDK2wrP/gXIUifGxWYxsG6KKXi2gvCSW
2bHTVKjLeoKyfKVbE8tbq86ZyTg+9Rrfj0v0e5K3J6Lm5pRCLm8+eso09WUkP+1Y
bdQGeTxNHg7e/9qpBUBLxunifPtrc7GQIwPyHcuqdsXieQ4lXowDJB9/298tpsGw
jzBu1klY63awF1UsgzGiQb+3OG12iywKUVCj12QtUMVe7cMxUW1U248MZIJ/9eT+
P1KgLQcQgXV5CQ1sdLkt8lWBiXPkzEe1fIHYYuIa+2/SjIb3q8SlM1NeoBX7hh0i
NOmmVHsq4SJzZH1ZRd/cNt2ukhVjkBK+kGwJZg04GiEiA/y1T6KbpZ7P9cuuZ0XI
rRC4tw8iV7zuShWcG063T6LT3vK3r2CZKpPrfKFBll69fBeSUmkR5/fnsdckdTLR
JtmdttN8dOCLw58LnhxL1iEvvZXrAD/PaWkCcbWgNRyvSKtehXFLOXzqniytS/Vc
GpGCwnvwoJvZyUbl8hhDFLgezLYmk2oOr6rG8+8zTRyhfnXuDXODuVkcO0MuXLig
0svglZFOctnXtaRbHnc3O1mpGEllDYC1lSPAx5gojqFWiEwq0cGSd4K/vu4euTkI
w9cDJTUaQ18f0ka7/ZV0xep1a9gfQhuxwgWw6Pvi2XPGXGnXisMlpw7LWR6veYhL
CfyFzfBkBc2nMVLHP9C2/PnhykC5Pnn2pQijTHK6pbl/Ww4tFyGqLrWVCzKbaHmX
yUuuAXDZKufTBqh8MnPK6naqLpQ4is/uilsI42VLcK+U9FkfE7t1jrSNtPvjvHi2
KAuUj5fK5N3D6iBWqa974MhNSATPgXfdJNM33AmU4P7jLzFvNt9Hn0/PkIZyiTEL
ypvEGJxSzR5+x4nqpr9mWq0gQXZMLHRCx6vCHgkUK8k9zdRFe2vuXxwDzuqiaSBg
eHzhK3BSUizDDlYUYBQcarvdwyweK90Gv0lFzogtCVf/SLKwdUW6i4OBCy9JO4IH
Q4RtEPrHRn6pK0/myxPlk4kMB3gGLtxsZZCeFfwP/SJsGKyttNgXzL3OkA9AEwnJ
Vk1Bv0/ay31WGX9wx6DZ44NiXoCx1mABcnYQVwK9lmXBAf5YRlgF1tu2SoXHelX0
DlZb//2W1h3xdrtazPjtcPfI1sWrcXz8ALf5Od7lh8gKUp4qWCZ2b37k3WdXCZiA
8S+5MsBbplrQ4ptQ0F09qpSFqyDfbhpMEqXe1OOvOW5ahEyDz7QnMYDX+t/3egSt
5iW5hAJWANcx3XmrocRV2N/fgBT+DaZUxC2yYlzvDIpgrUNVpAhqpAjMBJLv9CCK
1EflLmJ9+XSnyLatEPI7vA1VqgG0JmpSUF509yTyuLsFZ8PcFKvEywx3LmWKRORe
w1AMe2t4e0XIZ4AIIBNJ4Ki+bSxnpzz0XNCenWxWAgNP3zmDgen+7jIA7Dgmg+Kw
cUpJMxG8cTBm55DUTRj9CUCmH8MYC31jJnfuLkqrW9SSBBpHViyIvkC7v3OV74B6
m9AN/zw7k7LluoDIPf/23t+UzWzDLztwdqiKvktyVzshwFP/iUDnF7ds6T20L2ix
0dEcLY7Vi90pAZ/gcamDZnjoZiN6xWbJ11Ap4RFObofQFc3s4lHhXqyRaDxYoHjn
Knys9Bbx7Lg140k86sVrV1p2etUWZaHo3cHxDXs2Om5SrOsmxpNiFUpS/I5R3u+E
Ez7UeGAWn//FoUrDe3IYzCb2TUNKFHmvO5wQ7/1jk7NK/UGF+l4fejVhkiz4FGj2
C/NDPiYQRlYeYt8tCnbxCuP+7KkCEHL2PnC+8Tautn5CRxxlKYsO77L4f7tcZGIl
g4TsDrad4uFdjzYh5yEZVgOYYit4wM5Gj5oaDQh9/J5nThJXNhOLQme9j/CiRnRP
b+1irciBO3Z8aT5Z6gIG7Th+NEwbdjs/bzybJz/KAqowP7Od0gQGMha2GVdH7JZN
podN7m7Ba6kyKBrsCFRHFcoOI1584YcY89oORFfO4KLvSFx7YYJeb1ZCAd7vkUW1
m83ak+/mLHmgA9qjnhc3rlqpdhM0Pz4cpwHVwokUlyMQvvLiixJPeBLYYxLP8R/X
9wcxwpcu5JiRb2Uq+Kgi6BXiCYKPyjntSRhFSBMFBxnqWZ40r0nSscdiuwPS/TVQ
tEuLXZ0JIAGOkIDzGCVzHwgOrmtskSfx/taJbYVZozbW6BLX2szMatIoAM0JbHCK
wnNUvQH036KsheInAtW6LBRQ5L9IIANOdedy4h012d3gBVwF0RdsVk5PwO8hp+bI
84s2/5lQKiaOJCo++mxkw26J6RJTbbfNR1FHoqWUq2HHa1tkZfurkRx8slo1C3Iz
JEAAbIItDzCJkudxzWhKfWqFpsWITgra2WoHy6z/sN28njljVunSo15dPx+LgY83
OHdzN8lDMz5+Xlv+hy0jtPuX01GCkW8KqQV5TNihuaOq274sfTf0dvKkUp9w8Qz5
VIr3DpoPKEpR9M1NWoFLLiKV8u3ocLSWN/dcFMphgU4e/6OJNO/rldhHhs5AcSOL
x8H7dEpsF3qWFhJKl5RgjXjmSAM0usIw4Rl+q61hNAsJoEGeVSRYvxuB/nhv9Gem
NmrezjG9EEqIMYv1RROut33paOLtV5kDrFKq/GqYL8SiuQ6JhBpt1+s5bl3K5E4T
hyW/M1yhlJXWmN3KoyHFen50dqfzTeZhxJBy0bDWpQf5nlz96ModUOkqS+0LiGDb
NMoOUQRpp/r0XnjVai1b1ujUM5VyiE99lveBXEJAlkN03QNRjncqI90iaU8Um2BR
NfzFdp2GzgfhOwnAWJaK6if6ESW9g7A+uj3KA4W7KWDE7SmDuOmdHU9DfS7d359V
rX6Czuq1Hu7y13qABq3SxKTJLzAehJcbNYn6+/Ls41MRgL1978yreOAU0dmXj+iR
fsjdk0GD/f75vD1CUy23KskEjX9CNLXfcbzU84DXGtJfM6A2+8snWlzxkKEtoWpC
r7/q3aOFqnsY6NhUvh3kncqjAfJynfna27vpGcKG1lf9CPkKngsi7/ZCrS4yg8Lz
33YFPG63+a/Im1cY1CuRUlQX+tar710TvPdeUTvVphpPj2NMcKdro3ogepRN2SXg
k0x2vNnQL3R46CcWyzfeOywDyJnveLu5YTM8MhPrrfPoQbSQJVq0cXATtCGNSQ74
W0whs7vyrRvDiTGbD1jeDGlai327Ds985ChKeCVIKZTCqjSbBfvczl5AidsI4yoX
gcWT41HN5WwkE1+cYJzSh5xgG/FDWesU4cdokTkR2JSn86cAScXYlNs0D3m8Axe/
BUe04w4zKoaBu5p5FmPnMMBraVwg2ueZC7U7R1W+ii8NsXPYENABG6VxbxL8Nn8p
REhIuQCc5si9+8XT1G1pGWbsPUelkleHKBDehBFmrgRqpeLAqzkY+XaVHfKpaZ49
XyTdkwGB3hXMsUYrvJ1muvGbarAXnGzg4fUYArkI7XOgawP3BRUspkTTp6b4EpqF
dnOGuoQhcDlXV+kuTPHlsMRT1j1bCHyh+R9gs/pPP4AbFAdQmCMX89NryUfe6Yik
BxLlfOxxnYR0paWJT9RG1CjJucrm76uINn4bOS6ITof+wTNmH0WES7TyQox7vUPP
vAnBbkHx7ZMQYYENBu88u7bMG+zfJudDNwMEbWSDDqpIHR/a8QgKZ46gLTkNiD37
bo6nRZF0Yrs50jv+6CnsG7KZ2g2/CaB5eM3Ec5nQ0hOCOOPkRzWVRkZnhtYTY0eD
wxHvykOBd4AtGlsj+PHI89Amlqcd2QOUFeME4rml51veBEIAnBq24PZfQNnVu96V
AAda8b8YWOaT7dxjDarxMCXmeQ5GIP2tnEte+AnLFREuY/YPOWiSU7PIlqrpwvk6
DKXp0NoIWk3HpzjfsaCfBTHd4IMbFmcmfirGJDgPvZRVK7V8rBdbNgL03JqqeibB
34teB6vlHInTj3LHEW8XlvTJcb0xztRxvOsDpzROR6RnPgPkSqIrB7eHR62UN4sF
GDpzUC7OefuzlMpLD+2Ve2y6pYDTa1RsULN7y3C4u6+WIMuK8d1qy2SCUDeyii5x
fNEDbs8G0ybzYtKyCiNLvlQFu9lwj//1MeOAPhukm+neYE0o51O8jqEACepBYKur
OfOL0b5KiFy+7o8kWhC4uPBZmaBMGW6012zmYgi7pyCRRkf7Q9e/lp0hxYUpliIb
kqwMFOAbM2LLMvi+ANnqhtrNMMK51UKFBo+zlVF4fz3kjRXdYzGk8AJfMPNIjkg7
6SpZ4S2sGweg60yKOQe5eXXTMKUcM9KYr6QupSvtRXIuvSS6WeBnzxF9e9uRa1yx
EMzSfvyH7OHFOzviIUne9vgZ6Pdo6Pi8ockaKibmp/P3rF7vg+OX8woy1ylTqtls
0wjhu7TyYLeTQqesIZb00bpIRMzNdflrwpKHa74aDBxZO+McIkTGMTHpFu287gn4
ZqbdzanBdh1Q868ENjScQ/Q3QHA3W4XPr3gboN5/nDa2vTQ+VRhsbgnxFq61C8KO
83l5hmMxkIYHOCNV4MNjwtq/5MPymerAxnt38fSP+kGZuSEvL4+eGpEe1DGzOhgh
hIiyqMriKVSlGP/Sg4F5+zQJ5I6YP2L5T/ZkE/SozYuqPxCHf/sJe8BzPZ8rLRIh
E46wDbMIkaTBowgQg2itdI3Kd82TjJW+xrXYIg26UhNpJeNadBkwygS9mjrn+C8E
ZujfirybN/XifPVFDK82DuM6H6NIFtE89k3ZX54NAzS+o1wYnjAIRaBLYpEgZYvW
YVg8YqCw5M6GnAPtBrCuQeMLYgUc4YAJAueXPoMjRubIUs5/qZzPLXRooy0TKIqU
ScaSaprLEDfl+Dcc+Z+mAVjxWZAeiumiUgXblTqLHQT4BQHejvOIaAxX5jOjy/Xh
LEJNXzvSUn7nUQBogW54dZJY9tWh/pCagXwMXWa/OD0WJZYxK0uVFvfG9Azn4K3z
tQH/dzn4kx4kJAfpKp0o9KExqn3+ibeJknMd+tAG+xkYIBAI1El/CKb8qPS6dfEc
CyPIiuelAbAbrYCkMlA8ngYjxyRwoOLqlXMwDQP6oNTegT9HKTdfCYXrYYaDxtVC
whUL0vVhQdFIF8ePZObVRvH16AHv+cHEzqDC/qbJ85bCHmcVo/bwFpVh9HAHaZM8
+npwJ9+e3XIf692TE0ipSliIbY/B2hubpLDKDI96yzdrIi3o4QwHztI+PV6XYnCN
yCF5bqinj74LV6J0EqaHGs/yiQxsvPfAGkwNEGM8mRk7pz0+JVX5nmW+X3C13IZC
K8stbQc4mH0zvm1XTU9eJ6mtUcVP5zVaGw4RxGM6p8LLaf/JxnU4jBcwV0TfGoca
7BiaRJEpc9vJb2Mc7VrgqekHBn5yEKVxLDRcfiLMsV/tfAv5B9Tfv/v8jaxrBOOr
lQWVg/68AOo/rhR0Lj0hLWeJBJUkOi45V7NDPk/5S/jtAAple3UvaBhUJgyU1lad
YFo6zJ7zy948EwjhPYPHbqbRlsIB9vldhQmSlZsRn8ms4WrOldOc21NZvDZWPjfI
7k4Zhd+Nt5s6xdtyJbFwqbMWi2NJRUBz3+oK2tnuyKHOwVgA0+Ux3k7iJLKHyYOT
qVVne/FZg8b1c3uiGRB5rq9QQv+Z66rT9uz/Wu1asoliwgNmfRmovUt9mZiLtNF4
p4BUg6DVrqcPFzttvE0BK/B6A1vJlCVQZTLsxBe//dx7knWRVEXplrzOOx1oY52X
BqYaIeprazJUT7GaLJSUM/JXUFzajYeYDJHcq33NwncBPSL43QvBnM/85/Rr1lBZ
dSxMLAnbSNMOXvAgiBHqojEqF8HIvoYxFEjgMJ5vqBLqaTn09Cmnwe6uHeTuNwfR
v2PgfydpMmGApz1eFVB05hI96iax8usn4nBm6kz4GTvLM6D7f91vBTEWLq8VFig0
M4JOnoeKBOfjtGhIuOEBWkWpoLZRy3IoQYliumFa8qVLc4V6FVwW5A8tYDiq25DN
kHRT9uB28oZz9YsgfVf4ZrZgM6qa0TanxV5gIrD4UYDlFtdIZBBO6gMJJ7BBDoGx
jWyNprqF1kLgA1X52RExKAdw5B9IeYLPunw8sG/mghYuWAbwCORJL98E92gTW/c3
r0tev3V/W8n2jbZrEaPJT6bEh3kMlz4hhf5DZpcTufcSimvs49Z8m4Jfp2LevufE
xuwGdGcmkVcFxR2BfPezEr8LUUVLzfVDFyflQhBT/0Zd5Tydxzx//J17x+DFyHtJ
cfSS6EI3SnAmLxRnRXGb6n1mC21SCkn5ZvfcNrlGqI9GR2XoNtX7FnRrgmGfEXgf
cs1p5jGMl93cSXHwPFUWhSQBtlUWh60jCpy25P3kSTVK0/on4dbhpy3vnzdagPa8
GhhRhzN8gblTEbfIp+0BniHxeTTz4o6TNuFLyhVvvFc5Fggq7qfAsJj6IAaVLFek
5xjjB+nqhKfQCMRKcSGirYeU2Jt/BXrw6VxM6JC4sO/AajqVkIFRopdeaYv8HFkB
xVlh3cxu2Jt1k5sRfydfw4f4j4aqpUVsq5mm/bHeruGvq2ihV37qP70+hWhl+iCf
odnycuKOaXnwWYJ67u0smvkN4vEBSHUZRiWRSiNoZugQDrJusjnlnfk/e4ifAYet
2d3iurv5sUJJufYxl+snzVuSgtzuGAxIRfFvM+a5eVLksAZtHCxILiaaJqHvtw/T
6kEUTOuYgcpPpThn5eubRQPQK7dYgV+ccce7HbCZXgxjGgrQNmpbyuQY2u73jkDi
oGvsXSNnbTO58oH59RJU0xGBDvLOG9EV8B6dQnQiSkKc5OMWkrztvxsN1pWus2dh
tQ2a+oNXK9kPVAcjSl3bYKZQIBOPIqc76Xpd7tcFb6pRlOeq7tzu7u0RkzG/SkwH
mwduXCE5s6Blwj2BzSOHv5hksb3z3f8UN58RGPOfVN6++508nv6FEASY9FxPcEmn
fuUxM8vWHqO9OspIL6plo8V7XexsMv6uYGHQEiZTry24lxAEISQoI5JxLDuW/NpD
IR4fCbKiTOUUnSCYXz1UHh3/4Rs8v4Fe9bYeedh+yO9eRIsmSpA+JtlJUZOXA1J4
RCtqAOHnZWWJE8KGFQ6wei/7WQMlYjS7W+3hqcP4E/6MmjEPL21juxtJYtiSemwu
hoz93GlMXAIGma8n8M6xDreaPve8p0HpBOTP2/nHCSX8N9LUE7e9L1tdQHP2Ji3U
GYRUbp3HQGjchmUL7lYpx2NqwIp23ndKD//gjLT2eB3OHuWS4ShkJ1ZMVN9yp5r0
FVp1WvBJd8B3OLF3+8oBVfT2j78EM5PFlapaJoXL8nyInXmQL86/6WFOdP1dLK1b
w1/M7kvRHXNsxm3qwy9wPH+/g18kQxnkuahzr+mUNkvG0jet84a+LkcBhBOhrVol
I9U/qWvybjDVTyIpH22bMSo7UEgtpWX1zoQ8ZmqyvpToijEs3gyZCITDUL4FNI8I
waYqonGZB3gyPGX1YbT8YRioIvYjPyKfFLDR9e2skq8fkY5E2Qh0YvUNn2UKYy7/
HafEt+6pYdywDHKrBDddhvjVC5i0Yj5whQgclGMgX7QHQ6jpLkw+zb0Anvr8KPyq
GW/pRNWuNf9If6G+cgPI1XqbTLdTuAPcQFr4DcLx9MsTrPMl+HaFIXTK5tNZqK48
+RD+OCVypUGykMkAJUzHiFuaJZ7RPeIdhQEI6ocz+GCLpyonJEu1e9VMsVyNbo3q
5JTjTJ56Fp+oG4RykHKdHgj9TqbWEuH6ir7vBfE4qSRu2tRr5gBCstn23i5cfhPZ
i3TYYOP1d85WMZjwPODSL09/YOAL5jwzlu/3U+ONWVEaUmDwzk1XwOTnyhlOpNGY
L3XS6bdrlAvXBkkf1OiRNdD0q+tg39HE+zf2mVe11efgfwbR8gJ+3cuGDlTUWmcD
GKW21Wq/i/cMCIKadZ6dAhnyVcWBwxBsrYQL3e/iS5ni/G1WBqqOgQBtb6IolrUj
QYPHCNg2V7Y8AEEJgYrG+ay+jEZ7D1VkLkLXsKd4YNkGsnBq/CAMEc2ch4aNsTHe
bVZB6Rfei+ub+8Xi8SVoSkUVy6pzGvMg0xecvHklZaJRRVUJ0clsn1L8prpjaD7A
NiNg8+lJMJC78pzRA9lAS55nQsEQnXFbrU11Ou8fwVpWxRzPEZgPC91QrGoircJ4
mXCXozEc1umkuXTlrAsBJgQBdD5vSbToIHOHhnSZM8zVhA43xbijnq0UwyxCq1WP
BEcDX54X3DyHj2PuFhfGYI2PmLhObVSjhLNKMj2GfXSfH3j4shY1U12Mvigf9cbA
e5xdEA4wRkY3l0KfDgwgkBztP4fk3gnDAVBZrJO53OsBqkDFI7zqJt4mdZB/j7uc
JPCpO6+iEGEUOQxysCGlP0eIBpfl6BhuuenKB+QUqk/4R3lTCbcH86ATwHWb6/2W
/E9QImlVrtUvm++hH7PqLhZOv+bBQvCA7gbeuju4gDF4zT3isZbvwmsLT9xm0KsN
xEzRHgHrxpBZvCHd0+HgMLgoImLghe0c/tEexG7hIo0xJYenzSv5GZfDMDR7YiK9
1cyd56N03TZ5seAOKJMgltkQNy24L3pqkV1qlHIRrfLyELc3YZiHF5GkVx3uJYfo
xhgpSQF0A1Cy9DiDl9ql/sGVYcDSOFxNT7S6sQBbFKqZvd5wE+wOBMYHVXCVaGc8
s1OLN03vZ3jkhIssdTxFF2Ip58AlRjVPMdeMtHVs6OIc42Kx6MzxDVUm/ciuSioC
qrBhR7U/jJ2/PpEecysWPoCPAeT2ZS8PylJm2I9T7uZ0VgrCzyT3ENegfpklyOkB
gqXfRhnFCObljx8CYSzQE/BKJDbUdV6Cm8oI4eHQSRFNWPaZ6I+8AjSVkRj15SKA
TiS28YjgUfIbPpZUsFTqf/ZtXmQziNQ0XBVIe7DbS0BuDE01Rqzkv6ALvvUyF5/D
Tk3Brhsy4cn44RatciBvRgM1+8qEpqVqD4Yh0fpQK+pgkAdNfm9w8Tcz1Yq46q/f
WaBQzvanRUx2EQGGYsyXb1mW06urWAQzt7b3AUJ0VHoIyaRcVxgEg5/B/oJZodr1
AxhXF43InIElMdWklUqydSwR8IblFl7gElrMWibEovneWb/AK6xzkFI76pwfhmaI
VPOTPWLq+mAS6InmbIaPC7uXduqbj5nicH/Sz7tG4bOrhr8uICGzwHglre8mf3uw
t11fPX3gGTAeXoYeZcLois9VqkBm9zI/n4F/gYt6yDEBFYIlFgcywzq/6QXwxFY1
PsgIrfHVlEo047YcDSWt06jbCdYGz3owwby1VOykIeZ1WPDeLyXwcJ1pzPzhKFJ1
+zGcLOivy3svD0XhQoUj4jE07BUD3vO3Gb214C3oazScYBQ788TAy5lxODVMTxnR
WqIIxg7LT/NRvNkmhM6/qvjl3S03ZGbVbXXO1dUSVw6YSvK5kAuZ4xdR7BB51Z91
b/YVD+FjSi3rrSHVgUetn3b1RFApjrc7ZHNbMBnZyk+TLfi7fCl8KN6MyM6lO6rA
R7bYJvg2FCVRpJsiu9zxVQxHX4l4sEnde5P/5SdEcsDTJuTUDQLrsT+xtK0g2/IF
JZe2WELCmVPn3Nx/Oo0imvef9ReIOS1r+8hcPcXzBU09Acnk2+TtJLs3Uv3GMd2Z
3IW+pHSAYbYlfX7HL7hPGqRD2hO8sndmybbpvZLSukwUeDkiEDyyq+oJAsttO5ZO
KunubD6JZSVuwWz5UpjpGnBNlpuxJbgx/BBQBNR1g1AcWM5iWmz27U/1j8OHsAFa
O4aeA5PTET+jRMps42u/QG/MsO7wDQpwyEua1+Ea9r9hhuaO6FXW4tFHRpULRF9T
qs+R7sgz0ljtl/QvUGq+9hUQk7j8MIh5P/bzdHaRE4N7JyQzCV3gYcawQgFXvBJO
D/z5MxSOAmmjGWprAcBqVGvhLW+Nj2RIbuQNF34wPlNX3D0ZoTH3zil5xrSrkrlK
BHBrWSmV6K0tHZNgKVZI8JpzvAuHILm/vhNMUnwR+5lsjJi1H05+efovK3rTYrsp
lXyWnZC5gx1UexaJ7G9D1dP0Arp9UDrXAE0oK2gK+0yN3FonGyVeWA9rdUTi1TeA
fHVRFBDvEpK/ksIa/ygF7TI4+IyDRV4cdDJds7WxYwJU11MOVRML7FVz8qDi+Lpm
1zuEvJcAlgYNgjWE16bSv44qvJ7KZ6qHlEk7wMiEUoCCyaqgWWkTP68Rcj7d7+t7
6Nh2gImtGCNRjlYTRYeXqF70TAGkfBoRAHaB/0e3aZv5F85WfXJqJW0dOZfC2eJN
dltA3FYNlPp5gQUzEIb8vDZuJOTYIO6txLSVjG+zF2HCzHU06MM2EsOhnJnMNhIC
HyzujmM0WNsos0qzGEL0vWF7qa04cUk7DQj50FMC9+df8uCgtfdli9RlcETMHi1N
OF/KMANhH2tmKRJho5WRk4ZEiIZQE1/kRbf2rAaHAjTyho02LVzRA1AnPZFg0pHV
qy6UCYeCecHvL9vU2KRbFqb7XUJMR4Wfj11rm/SbnYkN1ItqFQOTPy3j9rv8Z494
T2NHUaRnge3PxbRyuqWqyZ+oDZ8V0Q8nZWgL6pBFEZSr/u+3a8efkfKBBySSTEjL
7NIhoVEhSC2DfCxTQ2FvwDx5yJsAGqElfA8bGR1Tt11GJpXGyZX9w5E3ciiO64hY
ejTq4+UsC3lZ6Vtov2tmXxv9R9nCpDVFf1KeDSyRAY1HK26rtByie8pEFPxxYjwe
D42Y8bjlKEqLP1mMVzlKcCk7qOCuK7anPEDTNkp58LU71IGAzYl/iqNgN2Q+fuLo
v0Zbi/gSFGch8eg1tUZ1rBDkWQpcE9N/3gtrGmw30Xvy42b6KTpsFD2GTpGsOI7x
CcNedF2AqO/RRureU8Y3A4my04/nSVr9ci/dVDBpbvrH/zi6nz306idXaEn9ZREF
vQDv+jfzjrZjX1McswtqSlcfPsRpWMNi7S8M8BPcLMUIOI27ZYdmEGAoXnItBZFI
im6zD3bFErtMba0ZbJvLd7XV3rNY3gDg0JFTCISpsoNmN4pe7LyPgoMMiPBtZw5v
pIxkUB+JGK6nAoSNM0/t5QCgPsPga+MFMVUyxzKmv6pOjppre/FgoxLn3QHmoH+5
GGvkJCEFYx6tu0SeaJQy/L0TCJdlMx7BjvCZWaKstXmRddM6ZKZQYTFRRLjNH+G+
3pwhgyxxCBTiltoOzgaL/RddakcFDkY+CRR3TkIz2mKm4zHZ8UBatrUjmjrP/zL6
BQboQYzF0Z/c+o8a0fbVloPmk8TkNcJYd25IW/f4N5O5SrABId9EQaOoDK6B7+Ty
U97X1Z27t5iOsjtpIzImacQ5snH9x7CHzlVs2uM/eiGfQAAPDAgAF40ZESszmNsj
wPqpEIPEVdsdWGXZ03aoyaNRIyvcMJ6FP5F+CcplNMhvFK4O3Gk5IsTgwEEIdevL
P1Rtu6r5ttxgBFrx8cEc5ksbvKtjjRCX5FSrW1gzp+POoja6isQqMUl59A2L328G
vZVgyvR2gen1G1PjzU3kJpBBIP6YQ6zzNOc9zL1wIlTJ1z6VGOoTCLKJWSKX9iRc
hzZyna9qml6b+ZTkMFMT184BUC9hBUE0+3LuIfKszuIq7FUSE8VyC4KRmAWNuYZY
z0NTP9LeAIhaZ63qDcgtkoabXVYyEpUjyMYONHVZZglcSr/jx0ak47VRabA0loP5
vzDiQpufHkuuliEB1eGlq7PeREWoX2QDRCCUS233dkeFk4W/b28ZviRhiW8TtGDg
YiZ9xkIRUEwD7YY4wWc9GzzMctyAYOFe5mqpx42KqZNqoRWyUDMIJwj5uEUsdavt
yoiDwsJKe8iMS5b5CCLPqwUwDDr715DviQ2xAx2ETq9r0s5NOZ0mlwTyIqz8exCm
723/9N/krHX+M58tpnVmJx86HL3sHmNGkY+sGTMXr5ZkziHMxvy3DdfDJ8DoPGFD
q2LlNIl/Oz9aHvibb8RPwnK1O+uYOQKDLebf4S4scU05vQnP3OZhilBMDipr/Kjx
6nL28ftwqTxcWGAQnfxywxyiJyaFl+OzH1POdVw+cqFzdFXu/zAFVHjiNvXs6vfj
4kq48OuY0HObeooEKqz96/yrjfd9SHcLa2W1Iz9QXP5oFKy1VMD+qpd31ZuFZzCx
pJFTAfcqIqFkeTClbbKGIV0k3VwS/bYm/HfcpNBCIxpY3ZAsvB3WsBXo8mmIUAVt
STuFp2vdn9BoHPUow+dpVGtR4Ud8rlakZ+pSpQdn9fVfJ/oUAeYlmGmpdBO7D2zM
CKL99SzlMcG4RpAOFQ/blS7zDHtQHAsVkPz5HXjzDAjv2sELpxgWxgG4WgNd10FO
AEJ4atH1p5NWsOZOhB88KWlGDfz0M44+PoTcjRb7ifX04KSn9aCsGSPnPWZXCDfx
Cy04cF9FwjQYXvI4lV2z26RTBR4yXlA+gumAMAcELotpMEyz15F/Ofl7VnM17Kcp
NprIpMuNIq6yJxpXveJAw2LdtHsfjoxQfubkGMFGC43aLLjsCSDvsCWYISCN0LEb
rK8H3/8CL/ALBdjsbZxu6KUgf7Y6dH0tInOASaz9lZksPXvxWdo+NVlmcigG6481
SSzw9c3pREyUuu8iQB2SabtzOACn73g+qeZVkEfPSoDWtEjGX+WMuXf+O3ufhSmx
P8u5775ypBhDtgFdIJpfnGR9s9HWvWMh8dlU2MQNaa7xluUlb9aOAJJy+YhAdMOM
qbsPln/ksxySSClJ48pjPnNCMCJx21noKoQsUw6blvVFpvp0as488G8bKAGw1LRV
1JCekq1gL1+DP9dE12DkUdYpDiApScEPuApivauxo+YV28OaQRKncjq0u9/V0a9o
nonNMpoW4UMZCUKF8LYJlENF1S6cIoJv0/sXobnjNce5kikXIiEnhcunOIhcnb4S
KmL7OSg/KngKMS1l7mMJDAEwNMlkRFD5SsnszBGWTl3lAJF4FB2ns+zdte5Iq5qU
t0GNWnVdDBnud2taymClX4zqhrWsXp+PBnCOTqs78315eNNB3d3MmoONNbo7HPd1
x7Rq5qilm4FDHWmudSdxtOAR5bz0M61z0z65uyCWdhVNVpQ6DO8PRPOlSj2LjXTf
2qgDgs/jB/1OoZEuraBT494QQN3QiOxi/GDeym4yMkU4CAVtga/7xJhy+FXJKM4U
f9WeGKe8Z0XF3ywZXzxCoMUmv/VU357ii17i9oWhSnEf6GPF7MFHLLjHAxpwDewJ
LOknD5edDTyoP5cxp5VD32o1vf+hk5s1dD4LlTxQTob/cd08H4p8tM+eJiE4WkFS
hqQTo4F2VCTMCUU6/KmemmgATIZk1pPmC961tSP4kA0/V4NPkZQ45P0QQj84SnNE
//vpnCkyJvxRCdGvctv23B9rVWK1ec/VuWcQLjfEhR9BZKvMm/gd7Dzckqzjqdz4
F3109gsLhcjE5xxcmt8DyWCmIBkt93m7sVxyEJAopIqCOCm19+d5qpsagiOPXc4a
DKijLCXcYT47fwNfNH8EHnpNZDb4WWhhM6iQGEx6AgMivo0xZRaUeP4wWWiQqEnC
Reww3TVbYIPEtGyGd4UNStUx06KMm0qemN71CfoB9EQ4i+uiIyH9qfQqRl6hA924
CwyI2a661zYk173PT3JqGmviA8oY+un/IHbXPyXrgUeaODHn3SOD+ohjy+z9pDW/
Tl9QgKt8vNqo1Z9kn/3OMXEuwJYB+dBiE48t6MojfFMM+TQ6DM7fsOQ/8VGfSeQr
++DFDfmmR7JLXZy799ueDO4m8A9KI8mccZ6WtwCvEttGM8ozxDrf5jPEI7N/g7ON
Ae4AP6u4umNyVnW2NTLQWdOvlH9lQkzzPA7gHe7K9BWQMgeXn8AdXNrTRFNAiBIA
/6OUGYFmpgBrbcnsnBnE67GbTjsXL/Ty7wNWW3UxThUOg0G2Fq8kM7h6KfESqdN6
kvpj8ugcRcmH5hyZJLpx4BR3cxKenDLZKUPWqRatRVMfyfOzD0PyHIzC2Zoi9Hr/
C9iB3SQWN+rlki15qmBJaV+yQJIUqQ4/Rsyv8zgPUtPNxGhAMU3jV4KHV/J2cGHL
Vx1MGhKURDfzmjQXJTRlF4TjBVJpIMgDTK7vgJ5JOQJczVyPlkaNqLxUCOFhpVuo
0DKH0KCSzhg1GEfBxCEWUvLH8AuIv9EZl1vnM7DWeTFUgFZ8mMCjYQtg0QsrrQf5
qP1Q712a2B+Tw2BVuzMi6cqkkyOJFmw4l+YzxG1Yo4iR7gsax+gteiym+bl4JH07
Intoea1Oi1bbxom1dtHXhP8gfXv8ec6DEuzbZin1+tGXjD6frmu9/QIPPTR3WNeT
5VAr0jfbPaESTnEhYwwqI15mmJrMmAxVyDc7gnbpcQUwUuN8phKuArtUTS504GbQ
wDT9YD/tJ6WvK7MGiOka1Aw84VFWvYXBxjJiflzUH946bEV899fnhA9pWa5+KDgW
eJi24BBmYtxyubpN3tD/bdorPqNg1W07leQl7OKuD+A1ZVMzB7vho6W52j6nk44n
09edZd3+nmUHQEeE5UOIm3uMU7mWkTFq+FS8gzFnozrKiocdM4hSBOe+2uhUytoX
W/ywYbbL+Xd3pAwFp5VsLw3wlSElZkizmfyMcr3jIpkwF0dSjdS+zsRAwbVFn9U4
pjfOzJAG4dn1NF8E93PT9c/FgRDtRm8i+VgYXziivX3EPtLWSn1mSEbMi8mGsVl/
cX951xAZRRjM6F/nHEeW9xnNhERy54AzWvECr+2yQ8lQCbGppwjv8eAfGcJL1T6T
DEc5fqUDxr/QslWfAENJ6diel5jyaVwbjga0vKh441QnIng5gQvxb6Ckt66EWwOp
Noc2Ntl9hBjidcAXd4WAybsPpqYqIz8egH1t2d4fI8SpWBq4x5pTAewk3H2UsmwZ
k56BkZC95gL81KBj3AO5wFghg0l91Dwx/olj5QXt1tLLG03m4OuYx0pRDyefzhQx
3Kpu1OM2LpPV9vLWZQuu4Zp8GzJvNF8lDVqe5ieqwADZQqmCt4VZfcmYBP1tS4rO
i1d0F6ngGJeax9zKlxFcZuz1dxGgFx5NVKfra9pmhuUFza9EE+NJE0KW6MzltAF7
9CndY4A9T2obUb6OIwq1fhgtbM/IEIfFWJjJxJZ9x1kKzpuzmeXy8+PoyQvcKKzK
vbr3tY3OUgekhsXixrDDk6hkQQELLduPm6wWGWY065kr/vWAARLefgWufneuS90T
VtQTqW1bNm1htdDEAOPVqbBG/mDH7yTpFi7gZ5ZvYDMOCs3pV5Wa4t8gpywIivEC
xrnqXF1AkwPx9lWGth61PWKSLVGK3M3Q1FMxrBpz/PLsXKKQSXjBGlydupnpdduT
++q1uhsKiFNjlUJRenALujyFnvMeFvLwamGjyZZJg6dhsB4gtEdBU2BBZeBpRYUP
nBW43sNbBY4QLqmMvUupDtFptX+Zu+Nd1yBm3lpzrWRYIEm9xrdMW39PbO8GDkYl
aIY+DaDC55gEtGNMsReqMeyT4Ik7FAKSAJ9aY95GA4yIulfd5R+x2cmf6PH3JPgb
LqP1TwPFDLQzmAxZh2xW9Wg+3FYK3tphlTwP5hEN4MhUXdaWMg9XydAdyJzf+KRe
A771ci67KifVkGgGdwL+nk1t5aRtGx+NnPBRKl4oEeIcgG6ot66VoHZWI7L3r30M
oloNyM09T3Ah82L3LEhTraBoOGK/ggSFPKwVPnh+PJCoIO1/KIKWww6Gi5apB8Wl
7hAlh2JqdJaij/0BlMtISsEGbLbiVT9CYSPKBbD5tJr5fS9v5WLe5blox6O9pEgZ
9OEv866hv7fHEd7FzrYnai926Hmc5sVrnjC9R3t+nxu4hJBd3Zfzfm3KRkKZu8cP
fYeDLnYCxVr+llZzvUmem6FnKmfR10LHDurUnru/kXxNylfSD6/nEvci641lOMZw
OA/H9HDR8HwqAU8oAH0Tw2JwXNA/sMAz/vrOubHQxpJ0HD+meC5lWxis57mjHf9b
pVNEKuZQd9KJWHxYN9eqN3pib8+ZMSvvO0VLl6KL48zh1qcctxVTYBaIVeUOGJFx
vSDbqTIHw98iLsDLmOThzWAXk+VW6Awc73Kqd+YXb9IHGDwI6oT4HKUkQ2vRHsAc
hCSVUeCTMWY8Hr0rj5/m/rXmTcSXSHxODpC6UZ6tkEdPoXuPYRLniDOvCR+sfCNs
4kAoXBs6QJ7Qwe7BzkW1RyjpEhKxOxOvXkXbY2GnQV7F04DnxtrZZ3pbuLkpK0M7
CKAiC6/3BhThoLMr7paSZKuXmAZO/dH5yxWkIoHxbpnlHSXTIdIpYqQfS7JeOx/P
+V8H/iTZfCoXVTtsVZ1dUk3NeuOvB26Z/WRPRCkerosTlD26gSDjEDcIslNvLZTc
XPNsP7Gqr8pqijQBnTDhSj0DX6yMcz5aPJ03SJqI97e1HoAUJ1ofpw1xEKZbgC9k
X73cfCJpJD2xr4edHx9hM4P6S9WBfSvPMFcbxUa2BpSACVfKf3dW/IUV+WuCJcv3
qpM34yZNCL1nW5a2aYXEyrrj9lhvSFzhRvQr1a5Y1XnuxopLRivyQ2+XUkhJuGGY
Gmf4V4JhOcgwIPXfz5lAkW6j3i2jXgIqpWUIrHsWwyx43DqFGWYu91IY2VWo6HwF
doRZk+/WqdEhD97CF7Vqhe03KAd0SqFXqpX3GwYwDq6TxZEOmnevNp07u6dpxAcN
O5e7uK7Yae0oky+EkFH5gj5uHHNYJb5LXrXBOg5OTnNnCrmQRV/0ZstuAd3lkJAE
giJuSOz1ZdbkmpcL3mwIhcEFPqaJ5goKTX68ucC4tuFogl7whS/UWyXw0n/hNgKZ
CpdtaJFimgqgPVbqu1PaJR/OWqO6nhx9zOO5H7CMhO2a5tsVzcLhcAep3A30gG5Z
Cl1PZ9r+nIrY3G3IHI6iIBQeedEASnY6mFkT3cYuJ9jKsQa9ZbxzXLSNIOaByS3C
ypYXe7qNX6JOjJJMy9CGuzp4xbDGp9YcPZ43MUqeZ1vIu7dT3WXPO1I7AX+LsM1R
utgTMk0RP5D3btN+0e13fLAXzbRn5DPPwxIRbeeTEyWOENUkoOxbtu6nA/95IZ7I
OpgkH2VJ1AenZYJGzZiptwAYuZ1YfTBFHiPSPo9++6Glc8H7aCvVkefAFWwHiTky
C/oc5D5Nm4q54Adko36tHrlFRYlSYxgeJ2wfcH2e4M794TMGQX5I00NerZSDJW45
rIFJOt2GJ9j5XoFRax3QRp5Wc+ki31VoJPwRN2bj8REVYEpA1ORwcW6MoqPbJamb
cdfxbmtIvKm4x6gTX3kXfLEdW5VSZQdFBJ+ANPdQf5vpXfYyimdhlkXoj0OB4ir7
f878RQiiK2p4wtTg+BL1FtYo07uIHPhroxYL7hWqM1Lu5VoemSoQKO/Cn4/roOA8
JDdsXT1YdA2z36tjrNQS7oS7pi/PmW60/WwBioplBPp4rO1Sgx4/jFe20nCZ/8U3
LSSf1Vc5Gn6fjGai4RFDWitsc1NnIc9xc75JMXXApF47fDru/zTymLYc+yGJQ7go
ezLA/1WnkhUKCaqzHh5c1ZNlOgLwZIYoto4pS7tb4r46hOty3tzhGbjLLHdrHA6v
wTE3S7+G+QzYhd13VqeFPx3q5P5yw6fyfP/zVvfW5cehX3oN0LOuX86kpV5LdDms
EMilF/0N3/qxNp7QJhJRT6ohfE8p91cNlZIDkrYDsXIqaQfokZDN3fpiLeehYX9v
2IHAln0JadtrtgLlTXqn4W1I4zQBrR+jZFmGFjaMO442CGfhg0HNJuLgVJoDSbx8
OZLjFqzd11KRWnM+TwWk45o71OazOEIRVyBj1FHaeN++qv7nBpoJChPWsrCFaC4q
5/dK7PcHWXYGfc8AIDf1sQOIiTVBNlIdSsLDJiSm02YNhCYL86GZ0s9QKioR6x4h
Y8aSE2YwA05nouyiORgiDgHOHMlVjBjnATZYvPbcnXeGjk+sba5RK9bW5n+xe5JD
Y6N7JhjMqtiNO/SLyepbRhFPwpCO9QpQMXKx4d4HYlnStpFOvEgfZJssNBgEkNCO
Lduyid/wP+RP0DbxvBe6Bs136RE1J74MPE3t594jYK8RZAtDG0xH63zT5eByS+BZ
ghh4uRPCd0reuHaMvp0SqBcxxRG58tjaaIGIpLv7gVMbgcWXPipwTX2EwQJBBok6
0Yfrh6eVeaOT3kATDKNr3Nxtms8rVpedhF2l+TiecLGv7VE22DtVdQkBnEMZrmt8
wXA+mwx+WtuZVzuVrTpSDlREnV/scX5syY3N6TKrNpF6fAPQvYWlry5yDLcw9cRQ
4CQZHbK2U53Ok8qt54zDFWWG65HfD0uGhkwKZ6wi788daKvm4wOxuKAxw9m/QUnp
PecmVuRcNasDcWYSATeGgrI2/u4adccbMvL0AkS1wIyzxWoz5HMB484X3zTXCmoC
5ys5u7yhVg6J1nxnkch5sht9kvGLNsbCFCCicNvvI8m27WMNmZqzGfoBMgzXCJku
MZackIIM+jo2qadAMGhlZmJcxNbGsw4MwsR1EoMj5LHEiVHoBov7yXXyzdgaSrSh
e29RxwPE+4weE7kIWGGk3luR/jF3ru54oI9tlUqG9C8mxJxqn5CCiGwGjHDCQrdK
o9OTJEuvXRwAonNV6b9OhupNqL+z8KgX/7pDGDbJPRb143CmsAHLyCLcMuQjeqcE
BGaMmwf6gfUCMqJQH+4GnYxe5f7K1uSd+AAaGBspgoKNK2HRvV0tgrf9df++CWRJ
HMJcg1zCJGKjsI3O6S2ZTC7sYfuYPB0mSYPPoIbGlrLTJ2J+aLe9E81+aUWJhBG2
GOQMtVVhb3i/YVEgZ7EP/PK/xk3j+ag2sBhYTRjv6UK4ObrwTK/TGcgVCGoo6n14
+Ft5gd/sabDPIbt2Hq8wPdAk1WT9CO/qRgU53D1kdtCDNqsP/kgP2i23yRoLWvLh
u4LAq+NrMWdd3QOOhcZNef9rbo00nDdp2ZyBbcpL8qr0TX+KRd0skUANo8VpBmnW
I3KaAtZlxWUyQ+Yk+hvU/AUGF2KWTFjRuXcLurYQJg+2/IrbBJVpOefPlXfzDnZK
nQFK+dmMmqMj03ZeGCUxAcCMbw/8K3yfr0ZX2XMzBqZYBxoVmn3LYOEcrPEOBxTR
vFLdQvFyK3IDit7/GbTPYm0Blwr6lEkceYtPwNoF2/IClw4QSP68SWH1gGCsu7Lg
RYC76ti/LB1ZiE43iRsfghLyo2Af79sO5qEDB35Uhxydr9MNilRRH0eG0iJS7ow6
pS699hlVSdqZBojeOH5S6RCKB4jpFunFe0DQxsKACUfWz4ld43j6uSJ9h3eGq2yP
EDFJhpfDj+Dd0N5g4rGlBIFCG+BzzdH6ownZ9dAROcmwOO+7j98kGAJYCWA7LfTb
F0P+QO0jBJr28ZFZeFz9Y9GQE1kKmL/Zbn3k0cGV1+YEZxg4KRupCCw978bySmMn
n118QARKVCQQ0sUNpshS4oWaCFvUHO+BIFtv7htEQ4/Rm2i8/1DpXTUHM7dsyZxl
XDxlOHVZfhZH+bEye85X8e0fEavfX8TuaGwwpqUpYzlOQWvkzY3mVCnxS4judScN
/jCPV9CpMLliCHrlGDwNdDjuORuLd38IswxgEogmCPwIzFoZFuTb0vv0C6O+WMgD
xKWRgWlt/FycxiPJLrG99//aegJTNdWvZQyRTZrwVRbtApXZQmBf9m2gzt6UFOHO
B51dEN7EtqOo74FtjvcB5HPU+T3PSuuVUifPOIHCszowwGhqHi3zC/wOf4CLrkOI
rYqNwJLPi1OPoRfyceqMlGk5zeRA508YIpLXSsvP+lFQsieJFI4z+XA2xMKJvlck
S3o+76grrulO+UAd2urxNklg/THs5wp213dUATX984JjIAzMPcR0i/0NyP3qevCN
yFo27k1Ow1gOdeE8MGeKjVfB5bO63Pw0BYioNiicIvGxjqHuZfoB6BB3xecbkLxT
f5GtVZ3jHbGE5r6b/RdyiDGT6ozJOckYZt4iBBs0rxAEGhtLpRHHtElbZvQokpjH
uZgUP+BRnp9aXnP0L9c7f+Y5i9ooIoLJCuoFgBY1WuZ4cqXwsnIE3QUgzBIucBQd
Oyf74/hB0x+47LV4kbUEGXKyNtMEGQaMOq/b/THX2af5f4ltHOkjKbirFRooCBF8
FFEh7UOf9/pS7gEyYA8lphQoXnj3qhGLTvf/8K8dtMEOmHIG5JfrhQ0CU0r9I7+7
b47od+AyBpO8W8ePlI9TsyBddk3lWvF2h9n+1cyFPPyiAS1oIZ+73dlAZAt8HoWD
fULk/gpVb2rvkYR9GuIXFE/pDox8Qz10Io6wYT6WSiXH2mxEL1fRHG/6GeN7ZIO5
SNTVM/KestoizWql+pF0tApFRKPhvcIaN4nYnIiDAErF/11w7ZMX6ZTeeDXAALw2
QE7Tp9sqRB2El2QRNsmF/CYfJ9w/OPE5gkPv2ihO/R1JF91kUGwL2CKaEr1JDpSL
h5HQpW9vMeYQ8BRJUfQrs8FcFEe1HF4FqeWXOX3QBvLAovIE19u7fxODOK2BhDkn
+odzVWQKn/uFXfw5LS3muKbBXXZWJVRE4S/FOp4TtNpux83cXahFKThMjXN0imcJ
JJS/htVv9qqBOWpZrrlPKAUOlnNOBzuG9MRJfb514lrKJ4rnL8r7yxt3sm0ZwwKD
u2K8xHISPu4nbNYKryMvVRG8sSFZe9J7fwEJIT8nANYhadi8dNVZljy8I8AZiqs6
Elep5ThjuBUDQ6YqyXVqBxNLvDd3LXD23gUDrd5pot8/q7m1GRd/0g/Y2pObdtlQ
7ah/aQU0QGTKhRc9ksgmSmpXUP7eww57bkqtxQ58P4J428ha5+w0bkll49wdhQ96
AxK8T9ZDGkSz4AeW7MQ+cUaMdKezIxcC1NcTVeFBCQfWeoxTLpu9xBZIX4gsZNNQ
weS3DMx9sKI8+p0AzhY5aAl/cSlHDOm4F9HXmE0h9W4Mxr4Rswf+drMIuerBls1M
twqKPTKD/1tNCbs/j21nPv9xapMisThSyaSDMyTy5j5cWxbgxwK0wYQmSLxSSm+d
GqZhVtnpo1egEFt8cIT94S0sxB7H4ebQ7zb9k6Bca7TqyK0eSqy0XrybLy3CNV5F
VR5UKHAsYsZytasPt2c8FoE2hhQfAj+V28z7Vf1tnSv+/11Pu8Z+9sGKmhEH2j8g
SmEI/WqIaL9fLN+/+7NzAYnQQi7puqWeDej9TrtDviAiCWud9bkNFjSroE/66XLB
bVieAnD5LHIaXUrC4ofXDvAw2PqY8Aqa30jgywilWHt/uw9HNQfIS6a5Lvb89/v/
I0EhQw2Ni+BPGcCoHBXs6GsiyjXbAgJ5Vm/ede/wkfvHH9fM3qMQ7rzg4if1MVBN
m2d/jp/Yb+9nkkUZ93ZCJbca0czfPaCAN5+i6Qvz+5fOYeuo023dB5nRH3paUH/W
nHvd85R8zvhCnP41S3mpvUHTAdGAyERgAuHSRcBR56vraY4JUhG0Jy65XWyqkCUq
IV86dGPqAXWIlYACztFAET8sJ8iCALTivM8/dKny/d/JT3wFxTFylfnnoF/ESZZi
L1e471NHThrupmwUwlTKrnK+gulYqKD8/v4K7Tq5C/ZYyTL0b6JamzCX//cav5lm
VP6kEOjas6vp3+/4gXC6CzQw2Ns3Tgj53/rITu0wHqCLcCSmUnmPIsHgkIk7drLE
jGME7/+7GeGb5EECHMcAE/q1mDYSyhIG2W4NhQlGHn87IYt4PyjQ1BTZ60vtZfMA
dvcDvCHdgnYPBPBf3Pgp0ewHr5SpCyS8bELDFNuz4sc9FrsBrvn9pPFXwVyEgHNd
LnWWdW0rU76mXAuicIoVNuMPeTb3IIk+HybDxuxBMXyeBWYdGcljPM9EQwvT/hFL
ONI4fzalgyVkUuBjPe5YKF3qhc6gH2uu8Mek/RyMHD72+2bmOYC1vIW3jY9hCUwD
ltAayIFuTItyDU/Wj5BMfPJ5vaOSVtCETorSTimdnu1Vqwhg6qojcaH4PbBVk+21
rIgU+0Hard3vbzSsjHzDrntRHy+5RgOeb12F0tpaK0a8Z8j0myzZTVuqnk897k7S
7mZJ1f5rjEl1SYiHapZt95m30ARQ9p3bRJO2Dr/GBrLIU5hyjkPKGHA5kpmNR1Xk
uXY+PIWH5SeCcVmsAR3DTcRuFAVbK91xq+w5pnmi4vdkoCsA2Q9Vm04FV/uACKb5
/jOjAWZkEqLaN5F6OMCaWPTqPcZO7nusCLd4NOBnXFp49LIkDRJCB3VqegyVAX+f
4B0DCxAQEamr4U7cBS4p6CuPBwWmVe/338YnWrzrXHPM5bQR+PNhYt/Hg85S4Rpd
GHKhzPj0rU0lCTFPZ+kdL3B67zc8gaz78J1aZMr2cxsm1UmOQwPgaa5CD2YSwPoF
BlMiNVPuwc7L4z29VYLouyEGfDjjn8faGMPT6qzRGTEByALBzGB3Xz18rOWKSbKa
2c4hlor960W56HN7FOYGbx7rgambHOcEwgakxUYChS/NMADIYVdZitCNCS0r0hpp
TQJRUS/Du6r+8wJ/sLT7rM/UAGeagRCA/wsue+bzOf9b++ObXaSRuw87W6ynnkEL
+sIBn0VKWLTz5/SIe7DEdi7/4pTul6S9bYhMGXEOERJGiiiMRRDkRjavOzlEtT6Y
/gsTwoPdR+bskwmnVyH7SGRgOI14sjLEaxEn0mJS22IkYhYJCubLKfRtckYEIxwJ
82HBfrUhsTL9thdPpBj11wYh7/GQNKJMuAd4I7c4NDpbYeTbM8oNx+SY3EV5Vjlb
NJJCfLUjS3geOelv0fvaQcQblTmtqu951R1P2DQRcWbAnE8j931ZsnGEMK7xqs8z
WB8LXb5ZCttAF1C1JB9zNySZ1owXAp/Pwrts6sefptDQ4eHI45NYOVdanvSRw6oU
P/FaIlrhYUBKWp23CBXGCIGkVJK2Yu2IxFWafs8JuKKejkB266BXsB7WrJzmnarv
BO631lLYqBLek1XFh4soCryLo+juxm/FWX4eSsW2Iu6+t+uFdUtay7VnYo6cp2Yj
ZeI6NaxlhOBqq+SWwtZgvi1x6QUAL/1cJy/E/BW8fmE5dGn5/TI+7ZkkvO9/tIhQ
tuIW+bl6qKNtWhaH4+dUA9pmmd2G+mO6JaWI3MAEjrlEVQu/4pQQOvOXxU5L8d8j
rt/u1hJoZZPSWu4ptT/z8H35xHUnW8SjgaYDrVqvGnrDh4g97f5mQcyJkhoI4xpS
aJzeO9M9oU5+cpUuYh289lqWvuHt3d+Y2OlZwKik/H0SE4RQmbAIlqmB9zRKM4R6
oozHk6V8hWey3xPIbjPKoJFg/nttXcqwIBubrmBOKyRVLs6aM296fXHVUWLopk3i
I8KC/64PBnp+RY4QIzcTa0Yu0tC8WvncZxdFztpbaqLwv2U1R9OuFzMRuUXCS41v
7JM/2FMqW7K7FJ6Y1DJCG1wlj49Mj0irwduoY0xBYutWOi/TZyC8C8csgI1c/Uzz
F4A1tSqeMYtVb0PbbQs2BF75+HesJKyEkVjzW2BxL+FHB+37UYGvAHpf+eyukgwq
LRpvrLK+PalgAiWPtGVzgkWb5Z3SWbdOsA+ot32cDeTGkzQiVKbJR3ilI144xvXB
cAkEGjONGvoTW+p90oM3tqpXUINBq8zKBB18m/a3K2JjP5Spcr/BVAJqmBbRe0dL
KdE7QPsLiaPjyUmIIDE1WqxSLY0Q+z+hFMmo1KjnpJ3GnKLAjCZPmjhLNfPailF5
ySbO+Ageot9MZVr2APyXZ2IrdyPW3bZDYubqfIxD2hVIvhoafuJ00V1235Edsvrh
st5z1J262I2bZDokdfKxApzWE95AdR0hyY/2VkA+tfkCxcT+Fkg1FQM80vXZajuv
SYW52UQi1OWKvvf0I1MGJ/6w6eSfypRu0S6pR3ZimVf6v+U0B1qBWTdqxJdIhGtq
dKTpV0lQqHzjDOAN5sEdhTASM2Fmmvr5jO14ibfNBf1koJnlmGRhIV9dV51Taf0S
HWxsrXrnTftKcskMUn5MijjmSrwekfonposAODZ3jrFU+zGP1jWKeqrV1GzvePp+
D3WRqW+6qLHaSyjrh2rPD24RXCOn8PxE1nhgjqIMsZ0vY8SgHOaJB/X8wAdSRcDF
BGakzp9cdGqStYfWIFuzbFFgnj6dqxbzjfZ8zrH+zRd6cuYA+2F01mWkysk64pCn
A4gOwvoOzKMHXHdd9F1dkYJCVGEfX465iFyGarUzNiPYka5wKcVpHMZTLsxoQleB
jl5+mgXdQEByaP3A8FbB17qgxAJO2dpK+X4UNpNUbLpj3DHEulQGLNamQ0dB+ABP
8i0d4HBXwsMVxHA1D327mMAsZ2x3ntSGp7468mAGPF9o36b31QCzpu8Wh89Kujtr
lNP4/JglSkQdMNpslKjDHWhdI0nATr0OnLRgSfEPq9mOot+fl/YPuLSHoilorHge
ClfdEr5HWsTqJalTQALRchg70EFE7l7WzAL6+EF+1wKHMM/7ra7eUBhZ3p5ibP12
bzJuqGU3zvCms7s9wuSPQ9jCHMxuBl24lG9EU2WIcrz/e119CdKb2gFULRl14gGg
GOYbGuCeJeXD1OYL6BsnAIolEjkK6dOspvxpupTNc8w8Pd4ELM/M1RrV+6bhFsyF
OfLZrPwcm81orbvFc/IE2Za57E56SYg9ZEBSQSYhoExe7G1pHqfn8MIzyGMLjps8
VTfyAPm3EuSdAumytmAygV2tyZGk9DwKIm34mBVFW2P1mVnb8s1oYg8auj+Mmtf0
clXILcFGJuY/dEvAROpnbMRcdqa+rhtaaDKijCW+B5iEU/ADyaWYs3cU6ofZcX+U
spGlybICunUViTMJWdx4Uv9ujSM2FJk/lBHBmsJuzdNoHcZPczr4RfLgnFQsBk9c
sfU1Wk5bXmz9XQWv2DGw+BsVl73H4DKQ31BoSiEt/BBIuONga0wnAEpy2nLUsovx
64L75TV1y+jknx7nhlNbNJFEn9yIMbbf9TDTeAxr0GazWjHJpSbMAS/1XIGL5/G+
zKyA0cj3e8cSYBP156q0yjoesDw8pNjRv+MVrU9DkoM/obVqLtxt+YLcixDq+XCn
uxuCrTPso4+ismf3TJvIOf9IxcfNvil/Dt3HgUjtq9XzUKeHh1Zho7v8Wcn27PIy
tiEOtoqkA/Zhlzr2hnf/WwCihHANrZQ/O12tLd+hTVB8rKOltXMSnBS6U29kvI3/
nR/A4zLRrPKMIM7wzI1SOxFZOz/cmJFNDXlU7oOK+2qsPVRRWdx31EYHH4km2tl7
vRAHY28odWkQgXbeh3VgnkTHC0iTYfNHPcg3nFV8xWvVtyMEFnhy3P1ZRgU3/yoe
VuZfkf23juFpv5TA/0DJ2A+zBpu8k9FiB6aAMAueokdGzY5Kn3bEned0g+5J+L1E
Q1dPpuTDcYJSrK5ntuLmOSLnNntYHeJnJKYhyIwM3hvY+FBLkkTrCtGRxjtXYrKu
XHT0nQxlbsK7XJ0c1xS4JPYmdzeTeD6JxDzkefPYAEIc8oM9LrOTBbx0s7xj/HBb
B1ZP/m5QnGssfMzhe40TH86ubeWiEcEa6KsM9bA46Yw56JoYm+zLj3d07kFF8ZpW
NF/Wcm/vd6SU8lFB90MnRd+SoOHb7OtrMJifjcru3jgFe5P50MEBu8xmkVHEU46C
BJ33NWermlD4Dgbc4BG2cMiEcqEoEEwRJYR3YWP9D/acyAaYSE9blx7VVXTDEQFf
ler5cakmJOj1AO3z3ZP6J+H6XzXcoT419UPqFBil/do4SqMp5leUgmPAb+3E5KB0
YjFZU1qN+jRVVqU6i7aUG0L0dnpX8Y0wSsxurQOcwDLV0f6UPg1rF856R3P3PZ8W
4rZL3QbGu+gLCRwTDPY7P5LjKkVVVQmd9THXaOAW7R13HtSS1c0f9W8LpLZFH+Sb
svgx0mA7PonL9cVDdRVXIWVqPlBwWjiemy0i71M82NJ3rzRyOe54P/+oPR6Zz9SR
pyYXaiS4iyLmow7KOqCJkwPoD60toCenrjiQ6BVM8Yftw1i0svGi7KUi4D08K+S6
zI/K2sGB9ynmUhfD/EbB2HWK2JD8SCmoMYVLgI38TKBgzMorKpWLYBxLmg/qMKPe
xNY9PyUhqGmNoeQ3Q7we5gQN9C+k4zopsevicNHfBJY6yZSHnoWE6k80YyBqS5W4
yFuje88wk3nokIwMxr5zDCOG/M3lhYeXnEbwzVmof1XTYegMCbyNLRZdYT3upgUD
hPAEgbst9ly2+KTKRRQQOHtAkyLsyYKbrbt7k1c5ShNoqTnDKad9EJDviTs5zJ3r
9hA+MVKZ2DdeCKXEdFHXGzQ/bWGA4Pb4Uj/xPeDe/Qp7nmcLidVAXRWTdPA9a6Wa
2kA8b/DkWKrU5TMwH7y7Wu29JnlB39VcFF1jf4AFIQrUcWyY49BgQ7ZOAXnYklzF
0lX73pFzB50xdAHIh4vtFP5KiIdh/LyDcxdkHvTHlcw/WZ1kjrhfF5HJdFYYZPNp
wZeKk41fz2YF9PPiHwVR/VD2HdtoqiksrHdQBbtMx+8pD8Umt0VcEiV24ND6is5B
gDcAuSI0W5edf1jZF4cpAjVDWkgsxlRuKdxNUTeyRpPIMqv06cEUwK9V7DaLHswp
6Bh095DCU7vqh04K5AOSwyN5iOENE1tJ+spEOEzfwIYI7Ur9p1731gHmQknXCI4u
IqzieV7I1vFaLmRuNplNDKcgBSvoKv8ncpQ7IbTCIAXU/L31xxoCnaPPwg59vmt4
8iMEHAjp9QLub00cyakD72TqFgROPwnHgmzmDISCRSrTkUU5W5cUYnmUxiFAKSIu
Q/04H1UvVqwda1DkXnx1tnCZQ4gJ/SrKLp7I2lKRLfImkRBPEg5IBPqa4PA0/Gst
H3JDaQ5XFNwqynOx1ZTcxihvdrpM9AIIAAPRcgqQu9ec67ugPyoCl8jxBlO5RwkX
JYWxlfvezGHFqX5vT+2pC+OGnaUAFmsWcIazTrq+k8We/2ZNCSW93vF+DPgurUQX
tJFFc72j2wgnni2P8/nLHAzZ7hoZsuWuuA5TNC8aokHLWjW0sWJsYj0qYwk8R3KJ
zXOvnCKEwLQLKQAkcUShRhSAZw/DBP1fYvHSdDRLlPYcET4sg7rjFO09movfioNw
7tlQbvngfPStWcU3VQJU65qT6r7rMrh0dq9WlWGatPvQQ/moNFgwVYDvI+chN0EF
eZALlZwgmuvGD3lCLRhwA8a4eiVa5pBbDma187dY8ImPz92vsjZpFrtT3Uv+2Qro
0boU8SGAzKYxyoy4Mfh3a04/cR/uwpLq+7/JEyL+rAVZSWD51+KupfyT4yqn/ozH
CxtDHSqA1WLXR3Pvvhk5bwo4KW+MvqpGdwOnI2cME7IbPURMeq582PMU8LpMFo6U
6SFXh2YGTerYO/YmJp1+e8dSd9ZacOIutc5KMPnl//fxywXys+mLuCuCG+cAxCm0
7iFppovDO4hxUOaMf5XfQc89TwmlDGQ6CSvxYx39kLXNJCkCpvU4X2b1YuybL6AL
VLjYiD0QbYxs2RLaUFWEA00efYLEy2crQwsHWR/cXmI3SZjtrdzw1VggPLf3apKt
5xPr4mi+luqzbw3fVVLiymCG1/9xuI5da8FpbXOw3kOfXXhN+d2RO8EHgxR2Cb5Y
9/V6Xcx8EQPgN4+/X3zQ8m+M31wlVfurXYuyMLDJJvxuot+OXqCCk1/F0+gH2/x7
oqe+Et+LL2OHuhWdlqkAi8UmEki6BLykM/QzqIEr603sA9DbPgd8/yQMG53jxCZr
kTbNErsm5PYN7sMWCaOfdZrm33S45A7mtyjQ8e0Y/d/nLCKzXgwj8ir4u9uTyu0k
IgT0Sk4YojSN9WQYOc+Tp63jPVcijZztOaughLYRLm7ptLFw4kqMwgoXUtWpOrSJ
h2pGUqT2g2wQqP/jFQgf4c0OciLFK0cysQu1uOZXWmSMkl+JRtiZOrnjUxcVLmUi
2jVA5XosCv2spApC6IT8TdNH6YBqp7zItCIWtfBtwWTS4UezpuaKBbA1GBWfg8gP
f5eZadBxCWT8jiHZpazngX2Mmz71oVeJ1HlTkcnvUmmLGEOgWelL0pB2/tS0AzVk
B6dxIj/8layyOwEhNaIDGJKHgGmI/79CPZgptcdawO1mKXyecuoUfDHMHr3rNvq1
tLzAuV7yKhuF/N1YfF3MJXB093GzbZ1LERYKCGpS3wOlygk6Bf1pmvtSYuLUi7lF
85usWUziNj9e05s66+7tKycGC0qcOwSudAGlLOTSLPz81seivuU4AUPAjGuDdpwR
x9gsawwkxqftS0CpWBW1gCTekjHvrVLx3sbFdotBPJ5PPHKcaCFv/RCBZi6H26OL
dpbtCrYu+kC5+B6bQ9TAOVMTEkV3bG+A3JNQN6x9wxKBC5uC4IAgnbiykHgpeWvl
vdxrgZTGYgTn1hMH2z8TTbLSIIWt/BZxqaJuutTLbVjuL8NTc1IFZnG1GU4BstKh
KYWLPpZEBe4Or34doT+28Xd8eaw+YNv9u+rWSAwVxUQVXcEjuCZwNEM+2UuO4QZ2
RcFUIHAn779VR0XDFTb/r1+WZQLPuUdKtHM56FCPxqf4xUSgrZ3+aFylScRdnNEV
ME3BJ9KxgM0zkZBTruewY049ouZkcrOvo5GRLBKCJJ0VxL5DtoRDhO/ejQo/blnc
EGjf5LklEW0JHR+tfMbc0uzxqdXZXdnKurwYijkrMeBTXvesO/EsKw5oxQXr78BN
kwHn/c/KpT5Rt0LRmW84+ehoiV4EtCoC8aZs/9FolsSRJ+tf5WbIx0q8trlAMzEM
F9o8fw0gZ2dsdi5w46txaa0VPd5jmZA1Tfs1oivj/5cZliQkhgtxRW+V3Yo/KA7K
ju2hZOJSRIfASdkWOnhfy7CuzBEzLaK+wsJLOyejgie5NsK131arCRTEVF9l47AL
Thm3/jBqkD/34wP6pLWR0//Vxrnp3YaeD1YaOLMPYBaql6kazfIrVFTvETAOeL9m
BbdEJa/20d6fyVmIJsIRHE6DkaosMeqBBF8i28wqb36yjBAxg2zRPs9BGcXUWQ8G
urL+bQByS8QBXvPSWYXVX70T0rSp1NkFlJlo0o5ZjYmwTfM4Ds1vDYXGt+jlGmEr
MRFNLEq1iLEqulJGPBYFLyqs60MPLj9oKwb3oLaeO4T9wBHx8148v2KZ+tYKK4TQ
Wig6t0WnXAvcuki9MANeNuJ/6Z90TXiQW+M5aPVwIWwpbnlhbxJZugYgqJ+e/8xX
QN60A5yHdw4rhM0UoaBw2xYlLd/qxCsepxUyy0KNekB2Z+6SKQEMKUUNmDiojHqK
LY2fbnH6Yla1mMWZMD3/CbMHCzxcHJ094bcOyQ7lqCaeKzDm52A1Yu2LX+11vbJY
+7hZ/o6FuZ6Co49ZfJz+oL1W2bwWzLIRoj2+UtkqbuDo8vba7cKgDzBQcYukH24H
zztIXu60966xk0fu9QsYS6ruilcpp++8NoB6B3HGYSKnupqcS5shWnSlxrGFW/eW
QALoWRun2ZU3QXdo2hrWJqAnrra79ximuDMHxIjIKOzSJxfYshdzZJ3I4Qr9c0+v
JhcrDZP6caWIWQofKXUaaKNfRMjBJJKAjnIGi/wQo1wNzwM3binQSe0SWKo1JGT4
Qkqp1IwoP3X1LY+wFMypwd7zZpcpF0QOmOUTXdcmbOF5+1slh30nbh+i2FX+JLXZ
TiW/MenpivhgCYrf1jDmavkxuH+jA7E0g+gYN9sb5s2w7HKBQRii7SoxI1SeEqR/
EPDDzIb7PaSpYZ56PRAEL0MaxJI5VIwN3seqP6Qr6fkohQ1pojISswq6WuS1nOXG
IjlKUk1wXGCFvqub877Jynlt60OU4PZw04TSpUrMr5lfm/Al0Wk8Xk2pctwvQucZ
MNbr0YiROoxc4yq18+cKqEoltmTykBBbJ0OKj+TrT+a/7G/47YBelERWIZupI41u
MHlEnm37DeUlCZZccXBn7rKswG7k1vsO+q8h5d5N6Ycfg4qPvnJp/MSV8rlSMHQ4
1OfoXnhI7VN74L0n4cWQHhLiQfy9xDVL6eAK1W5Z5h8cDuAv6Yrn+MdPNhzLXbAI
K71L8lE3KsQkPGbnoWMUPQZ5UgQ4kO88kSL0LPXs+5JRGEWx82LQL/5HGicOEPZs
9NvJXEr4YWcjbBLoj+WOoobkCyYXJ+AxrH/UjrU43SWTMzN0c1moA0+yVmfNqnAQ
z68MI6u7o2hGTpTYOsj//EIw2UVkKcMHXRaZINzoTEJ1WNfOEtWxCeu4CXUgXt+W
vW1PgfdpuzPcju7Mn0Xy98ogrlEEmBTUgAzXNygINURmumt2btKbasQyu58WJt3Q
P1oG/tcEvGDoFo8O2ds3j20pk6v/8czEGLscyZx+FINGJPbF+eKjRFgOvUgRy76i
UZh0E6aABmTheWg8rK3OZCwu8pN3gM9Vr8x6xkEANfdPAHDUOk0GMHnLheLAM40G
n1U2SbI6WKa/qmDxGUTljLuO9VSdHViMTF6zX4AWTjGnfGY2sm7Q0WbKoUcyJCKf
NZ3HVE1Dn/7y0XHh37GHSQqAyWmiIUSz2qI35eQe9teNrtCE32MFmM7QNRtUPB/e
KGqLrfdJb9RWL8UF0JqbE28dhPZJmGxdWUEQyklu5obHrvx14R3pRTdhDc7zOpwO
hDEAlQMdb7QHlw1iXmNbfR2kV5v6vF1YIV6ei6sItuKbivOnTF7cjq0RYS7JL+Zl
AhP6HT29Nf3xhHfiGqv8HMmvrCCgy6N0YpIRG8oETauqoyRaU1B+3By7dOJ27nl5
feRzjHZBy9GvsdjMNXzvahUasMohtSbJg0Y/+tSqP9rj0PuF79sf//fY/Tq+oaNc
8E7Ks9oXZCdeXmKhiV+XXVA+Hka9OwpIHcB7XMcyjk62oPWtlwSr3c99jgo3PhT5
6+2NsPJ2Ifh8Q4XOAtrS+gG7KzusS8g3hQLzZ/RFL0IYsx97Zkb4YDfrwWQh8qwM
a61Zg7AxdCPSJcrHGqT5H2FVCA9m5fZjD7o30fMmkUJ8zAHr0sXd780gHR9WOHpI
iyLX4R1OnZ3Rf3MWCTJGlC1mOediihsOMe9cBQRPfFyYVzf5M2W4sPVpz9T1YQx3
ye0qtdHBAZbf3SE1dBchWc/RmD6USLVXxYUwatmY3jPN4WATDF7+2vIMHLrj7fTX
6sg9pYrv+8KLGHOiJ/5Z0PsepWVEE//MQT0Z+FK/u19TaJdepc5aYpWIBtmbnNdo
Pz+qklBnSwyyEN6mCcKp/gdcxu5GT0BupeRJaSmelgueTgoSvjHjkFhdvq+kdPMz
RF3iHKVToiY/IB1N1cRQV84tMK0sftXXP9sWWSShRWaddpITuGHUQ4tpVctwGyNd
TmBKtKlbpzvXjqq8J/HXPfTO7awyoI7N3NfVPkvtl2gT01zhmLEp1228J3B7tJhk
VZ2BXe/2cMUZyvef27uTdRD5Gg5sW7k9SXrsyPm4Bj+hWe7kGytYF9a/68KFmV4F
Sek6ECLU8zdmcjpMnlj4Nf4GaYdthr5PwxSGYDGyliC52qkCPHr9A4BECE7N5qcC
CszHD+fLgbCnun4/WWB+YJkfoqCj4glBNgCsAhL49m8Dt5ncqWI/2OnArJgFsfxE
PKAqe01cVkqbJG+7jkvdw3V7vpt1lUu8916lBFAauB77NPJlkcpHzGS+GS72v0/K
MRqF3wT9UPRPUh2IcMEf/R7dS4O96EyAMp0jR1fH92kkXpFhk6LFzbJq/ZCfd+Ib
nG7GRo/KEBRPFI2eJj/TUz/YpdXsMH5sQFVBZ6crwe2Ys3mVBmpqP/OfmE3mMFmb
4gnzOzS6jjPLYP5nMjzb+ALCG0Hbg/t/QEjMJ/GNNrNr1ySVJDGQG27wRIHwZ9+y
/59UqIR3KpWTH5mStuZ9Qw0qWh29RDSPUxwfi4lHaNA4JEntPmDKp6H9qWJPfovm
kSKVIBe5QuO3rg9F5s89Cy7E/h+gEJ+6SJjskuzezVKFUOD++LwQG9jB8GnTT6ob
nWZ25MHWdyUu/nR4LZX2dga2QWnnlshQjLRofZ0bTLDi5PCNAfCwa2bGZXN9qo79
2kIyJ4sEzk5eRJFc7Yl7xCXCHSmFIs/OO/qyw63EtAmRaQqQbqeKp+o/kPWmIDKy
BzJ0/kzBPv42Cx979+XtNrWt0HeRC0LdoCMYzxdByISGluLbRsta5VFPG/zkZ8no
9IleJfPzfeyMuxx2ZpZxwzhmOAEC4hjPoc4E2+/A5ioW/8z+QIJp1Lopjpa72mIc
tBHQl118weCEOOV9hpSG3T1jB15C2SaGX9fqquDimTSPByLZxuTwCDoU0OIALx3M
O4f0nFZrgKlN51/MszIs2soKn+JUE5WjBfwJJARfYKdojePURNislITTrVX+M8nN
3yhahH5Yp9SgtOh/vRDlq/BTAnwFuno02aQEYb7r8YkkV2Rb5IckvHEED6FVlC+P
EcAAwf5MUwu9vvo1JqK9umyVykuGQTUWLUafK9MKUMzjg6WY7qmRHfbb/qYZY0Lu
Oo3r4xoLHsh7qJpab8M8qPxffzNAkl2f8OGisBisKvJmmcIGeLq+wGJGK1sZfBmg
jugWyz/vpRmDGsg6kHCST5aNdu85QoXmj8yxN44SX2c4nUrUvI0vRkpXcNEfv9Wf
DHzHAi9RMNanc63OOeIClVoO3kJBZv6jLf76RRQaMvuLD0htvu//vU/n80T9Iear
/Ak/5Z051lBu3aBlptPAjVMHzW+q2qQjBHadaQZGzgwkS82db5bd6oOInIIKaw9A
4GDiwVgQ3tC7T79cV/k8AqQU7pdceFFAY9gRuh/1CL8Bo7+p6AHo31nvICNEW3hA
5PIpqTj47rhiK2W75ETLsaTuW7DHrOqx8WF6jwMRa2Duc2laBNNBOlFu2ayf7A2m
47muo6O2v3YUruELdSG4NvUxP5cX3DfFFaIWCFbR8zr4yfMuOup4fSsY0Pcp1kx4
OMrgVV3EIb6gCp7Aiq9Puw7LaAb0ghUBO3dKvlPFRbThqH7PVTUJginUKtabjP2t
AFrOxJ0SWc2O5kgJTn2M0gmJ0ItVCFg2CWsCtuEPR/sGYkhhCTSjduRLVzZkQs1U
JpX0ULs4MIuVysaZ3jEFREAWly7QuvIOPh3qj/zRtFAxcou1uMF/IZN4f1r+36RD
tTpXhbYNDY7E8VL2LFyU5NG7uew2u3scLlsJ/IrRdSkde5QeFKe6/J5hGB1FydOM
0roIeuKNrAx+NR3SMQoHlRP++tHewCH8qoefoin6gx5aLkP9vE+dmejUnecOqSmq
01fBj6tLs/cIKpEiY+rAzEG62sWoaNIWTOmhc7/UUTpp+ooFvbwEcKRf+sIlgy0a
1yM8EiRIGF5hvBRGOPO2P5LT6Eq/0iqyXOq2INye+jNb/m+YssT1nD1pvzWwIZFL
mlIn/7JYXnjT/E/XQmMrWZWoKDvwz5MU9ZZ3sWitZVQeeF24KzvuDUyGhbymgat7
8qFGugvRTZPb5rYyzzMFTVDtedYZlZ6Zb+3ZHWDvcQrmYoO8OR5pxfJk8Jy+7K2X
oMglJa4NGWAabui39u1OMURsQtk9Z05+DyGTSFV3uLbs6XS2EXlcXGaQ/N0EXmmH
eqzRimiwx8uqh7KyexE3j8Rj+V7yibU/KI36Jtp3hkWTrZ4hjBXGrUoufjJKJLqW
tisSOnLI55SndL0Cgl59nyxOjOA42OFJdJZNAIDplmYYd9gmV26MaiHJ626OLeIp
vxZIUv+xNnovvdalWD5NnMlWAYWAY++Oib4lj6bN+J75eZcBt7Lg2u3+4cOhbDEP
zG6XS9Qed6/7wyaEY5oUP5I73P8wsl7Y+bIbK+R0a8w7yJKdXRW89IuIXJIg1I+W
3+dAX2JBe5pPSpwaEr/Yp+/SOusSmhPBQlJH/IQTkFifST02FFz+Uzy7lxrErktn
rW/k347xKh2lplG02jBH1XmHHI6XjZ3BSRxQ5lyrATh+zey4emQwWaB5y+OmPCkq
E+57KZWlgZpq8294ua+JWmhU+N5TK5czBsLjNsfsRpaulYWVPeLGqDVhpAwFN3V5
YJjHdR+W9Rrphtm1JLvKqU1rTuqXqBjfGoapFNT4y04/9RLEcqlVnXRJaRRL9sJ7
1E/YRs6Iw7yDTbyw8k4+VVSEHcm9ITX39tvnX1IZZ3v8A8BPTCufMNQVT1znKgKV
jC1YwSfVstrCxOwgMh4/+1ibuIqwy0PEhHuAG+NXL7NHCE98VvsHJwxQxsRy5BQT
/xXViM4TevO7JgIsvOs/eqagK+Pclde/LThTY0N79wGxkeSlevnSu63yl5Uocskc
bfD21h2B7cn3oSKniynXHJsse3L9NJmQs9yVQotsuWeLMvXOXFf7qMdZqJYMUijs
S0kXLbGniSMHi8owZTZR43HnlWQrYVHzP7W6w4tsfFQf3Zelia/yywt6dL3bKbWA
pSSCcdX0Htal8EQm34Kokf5x8zQhqPQGFgoZ+10Vkn69miM53WCY1CrLhMhMxuEQ
9vIL5ZE4iKA2T0aCmQWx6MbYfQeJwlzS8OgZshwHOQH8ZA9DUzFEv2k/Ros3UlF9
mDpwoY2qeMN8GoFO5eWFd1wYF7IFUmjlYwUjTm0dFOnmy7ysKU26F5YGhywGaFcK
tmbe2UwHQl+PP1OLDQXxluoYXccaLiqZcytI6lwertZDyr8YFxgOwtB4uUzHO8fq
RX9si/J5ehGPH5WF/fcNykakqJIKrcFOnntWh4vwd+7kChHBC/uOqlCOYqQ/Y7CP
HuDLzYhF3RUuTvBDFor1MwJoYXFBF9g/l9mYtc0/cU1uMD6trOb1FlZOnVhWwD1i
OETOS+9eJOLvD3zTdd8bDzc/CTcz36WYpmpv8e2iX8XYiXF4HeAY135bymv9K6zy
EUuFHgLyY+XJzPkbQi2FdKC60n9jfFUNQa/2yeEqCfYwwRDXL4Ka7Irtf8CnW+0k
agsx4lrAhmbexwPg8uQixLpCeyO6KXsCnuVPHihhmaleN6CME99V8vYkqxOg8lN9
UC6flyQ2AxWdgnLqf4qo1ZnM/I0Le7df9t9Z1gLBtBfGwF60UpbR8Ivxhl4+KeqA
uRXOlzXAjlHBM40I7V6blJ+i+8F89rx4g6R45Upg704lzjm9qRGLqkz77lyt5bG+
Hv/eAmNEMbKlmuphzj/o4nWkuhbNPu7p0JUou5TRQ8RDXbP/NAawu9bj7rqzOgKE
NjfO0aFmgZCDODNbtR1kSZeUNHVZFC7pvg+p1seZA2V8dZw8TKuyIhT8voWrIboc
Yb40uT2q0qjENMtDiZDRdeO68wu3y9N6Y5xGzEtiWbpY+dn/3ACkC2sbOcc/brv8
sSffDX6eKTDP0xnze5WO1uhkztHRwXL9rkWL/Pl/gu8phaaobUDXIsZtbHcpg1Wq
GAkMhcQpZY7kIiZQu4g7wB2DQTH5tc1Oaj/3l5jkr3sW9Jj6h6RE9YDwI7k67fgU
IsPNQg2V4egTguFKOsVmtSEUhrZvv+nNKg9fPYqdH0H/z04b7Dy/dRIRqBQ3mSI7
LKFJGJOqC2P56pPOf7bXQRJy7+PmrWqspAKFUw0klUba5LrseQsa5Z/rMXQfgRLR
gWB3+970nrCAgrJ4HWOwXCefma8HcpEza52fldJCFx0BmJDYHLzOnEvgz4or4K2m
QHPN3sA5EvPJAac4EFyD6hEBWGxCXEACTbWtozxMC5P6XPuA5CZeivsJoZFFZCnu
c4Ncds3izZWpXI0qmuSXKXkSbg8wvc/y9hjTqsD0x9NTpxUk1wHvdVUtWB0jtjvk
BcbfgC4pEaY6jA8AcwqxGt+dLnzaC3LFtdUmg/xy+TDzt5XAYLucz2WQi2fBopkJ
fmUU1FjND03ISRi0s/BjTJ2zJefu/NMtCtbCyrkuq1f2I2obDmolgBoE+FGP5iUH
sHtNu3RXCBkVU156jZg7gPjvq0Pdp9zctJ03AXTKLnkqG1hWPQiCGtIUpNNgURj4
U2CqEjoL2Z+WFejhOxrgLSwanl7w60Jl4NqXCb7C6aYooIOGqFxt2LCNIDFSImet
qqXbKQU5Dil6tyrLiZxdx5mCVzNGoHbkPuBDr9lwN+aYn8Ee2EFQogmhBnAvP78O
4tMlUr3hUjm/YG2WxSg9uTKKYEIM7SaEfK5t+/w9rFoqzgwbKvOnOR6LAQAAbFjO
7sZouDpvywhoG42ffLSLkeAfCZW3Bir/WHZniIQPaAguWUe5vKdKGwJJ9wu1DII9
Lb3zXUPe+ykXkS6gv5Qd4ifRL8EHuT5KtCGYdUfPxpKKXoSi3inTgQ5rXEq5hIdY
qZDucU5BfTgm8nr7S8lc9OP4H9uUs46VMlvBPqu7GLioVMlcwzAnbO0BsrwxoeSs
xnuFxAaOk+ORFLySgouXViFKK6M6MxLe+5OPqbx7uInGa6n0IYieHiisXe1xm2Ad
bmkw90mcww8AcBRxE3qE0ee6iGqjPPzKQO+6XA6rKR4Mn9LFPBSor6c36eUnBOYB
uZhTiykYWMWIaubmfFcAQ1qSB/wMPOweTuFFX2uen/uDLkVSv/E3dMi5Xuu959Sj
9JpYv8px8fZbuBt+cA8fQK7w2CK5iLa2PDfK3WEbDZ1iQxBL4UuhhzTOiW2e7/zL
6g/Ovcw6G2xOjHC6jk4QTyHclkGYf/yqMW6mWhZ5FuVzNNvuUIysAfJbXWwONqXg
yTB158Lqsw54u2+cwiTmTAc1DxBOKjJqxWEFcDZjZFTcZJeCM2jVy/a0e5v74aMy
Se2plZgNO8dsdR+13Ttc5DKvjXjv6rwfW1Rg8eH851r2gwj87fK4I8RfVrqADvAn
S01srm4B03a9fwsO0A07TB8PjSUDMV6tn4xHEZ6edMj1s3Y33aR0kQkB0iQ0TWkB
U/89XqZmhSzvu7+V134APTY2UzIfsb9zcrOTKBghq2bAANRk4QNE5zXfIUO4juj/
KLshO6GxECTbaI76Ftkfc0UmZKfTSPGU6jWVgaCdGgAet8mjn1smsJ6GHgxoYy5D
D364WNtJ0PoYHaBS2EAdnesgJN+MuzTuJCVJMaFIZ+K4Oo+ycHWzjo5rt7QzFdtg
PYqZPc9P7P7iycAmhYOSZVNPWn63Cav0BATGrff0OmFVa1vzTjq8GfDayZjyK7/5
oIW89UGHPnnfgduNt/uHUfdxwqIF/14bXlqd0z0OxIw+8A/9pMIYfsPoK6Zn2Blc
QvKsRGTOKd69WztLET+15DHvLTnB5Q+sJTmPOl4SfxHy/RS5jF6Ga6soHoEMlWl3
8YX1rufSUBayS3kVFsZj6bN5gvhTH1ZgB0g67vTUnjhUzhCXur0S+wH7fZECfOP4
MukYGYHneucrQ2B2oE4o+j83VQJ1BHQSIHs/WLsd9h0WAUTfhLSj/Fr2nVXrjkSg
i6qmJhsI4HD1khzjf52dqv5qQo8cy7UNPo/g/oTQjEnhlaGH/Aixidl4SUKGsBa9
5JlbEwDZYyW8oC43tTYsKUXkZID2ZgDodE04UTgvX6O7cO5pXy5kO1RV6L+ypnm+
N76pLjL8JVLIcop+a13WBmYseZt3SCGVst6f61cMcr22936wlnPkXd21sfSB3R6U
ZoI88iX9RTJib8b6NixO5oSAH+Z6iq/0nF9WzArkB2suTn1qRP8BWkxD+MXr3q70
Q3rMltGIwp/tHHPESpYNuJYyQB+dR2lZP2iuMq9djWVp5+YaV7RcFyvzYYANw6fK
UxGlSuOmfO7duih1I3D4YeSMkpyaOqPHDhkgItOyXqGBRW2n2g7PTV9Sc8QKuvgV
ZmS/cAxk51Pe+ZS2xAyy1YsQzUetphQtPUzGqiT/JSB5yj9zqasrfnkAQKGpIHef
QhXuj3JiFTRGa1fLCsnsrGvO62lNmlBEsqSGKRt2J30cnzXGcmP0WPdRpYqqFhKg
S3sNkST1d3tIsg2a7Ps9gfhTiukmu91my6PUYZysXDG3JCxPJ1Kf5cqy+KuJPKOH
B0c7bVNj8Sc5Y0K47x+tZ6LZmmggCPlJRRomsCOjD5S77psrvFYrJxgxYj3QuLvC
/BKg/q1SXWlq3yTEajArMvNBTVyhsVpfI4NxdKtunkmLORdIn+vMeFFgk2p9c8B8
zqQ2izfiD0mpQJr29fSst6zdgEbp/y8+0nmHfT5JvAdMavvxxqEaSM4fJk6em4xL
8l5XmdI2qYgzZE6jMQ0kR+cZnprSf0IyVU2kXWs/QtumF1q0lgH1N0jbnSaSCAvV
LgTnUVKEsxp/p5SpAs6RYIdtae43AMEBzt7F/Z4vuhUVzVCiiQU1l7GikOEc9PxE
tzX8NfJIRLqDte30VNuwDL9T+cBnKzo6f0moJn6eGLcSSX0eOJBz+/Qfpvu+A6BF
lCflc7cmC/IE/isJVHFq/gM2ufgxvBCUUqvpcFd6613y1H5bZCHWw7+FbgVUE72a
eqqz8hTPrcOfTZOyGyBGmqm88tLCKdvsmTwW4Jilg9tAAEmPWgmjf6acrJI06/+R
dADy2aH9f1vCbBr8k1AFVxvGh0u9xBaYiupowb6GFC0uKdFfmxGTkd2TCX7zif4Y
K3JRUJ0rdHeAy+nShd5zAcElm7M1ELDpm6aUzQI3DobbSgNZiSew93aJr9fdLWWG
y1jsMxkDzuN9J6if7RzUxlzsPwOwKUy46Tsfe5ZJja7Apj8OChhvlQFygCwEoQ+0
2bFos7jrX2AJOxdssJ9UAqWJuWHAsN/Le6GV+BcrD45RbzZXNi2NVvJAx6a1aFDx
dgse76PbAklvE4VgoZcffOfbbj/Ul41oY8F15nS+Gk9enS0FhNgQByXFTMzn1XgT
sF5CtWWFPPHBTxp9/I6Xf924pISmlpo63C+49c/o1GRHOcidYx5EeXZkteJkvFJn
rHShLt27WqxdNik+KGnje7+Sb/AtOefsLIxO+ztF2rj1N00ipCvwwXkknMj9sydQ
xqmI/3dtFlk0GffKJbCQEzCXD0hj4H5Til7FhrwKkVF0M3tyEdOPqbOzHDSctNQF
+ZCbZZgKQgk7IZ4efNd3PU8AQlVVZt15vheC5NHq28CY8QPIok82GHhC6ErroTKb
EPkjnRFoX2Gmf+MUQZWIQ7ydJXB2mM72DDvDICn9TARlwaaQLa4CxdLpTo5DylaR
/E+glrOYRq+VL3YjySs7GCxpEJJMhScor8M8P51jboPTnynaXd/DXV2PrU7lSNlF
GbrrFMzQJYzbMHI7n2G02dSCSIE+gnIO5oY75psaGBnP8ulwyQpVvmjeMts7Deav
lcPaW0RlCAdjaHD1UA9PYD0rqp6wdPoTDy/Ne6YsLPdaxaXCQPG0Xp72CNJwohZ1
MIltnWo+ll4G5/jRDkJlAhC5uUyDCyOdncjqgqGV/hy92J+DBq8KQ3neR2P9hcFI
rWh12w9H8QkZY5K0Gz5SbLw89dfTU07AL+tuBV2YH2x8FeW2CqPfGsk1ugNPN5jO
QJxGqZZAjWAMvWcTHYNztB1P+Zr3KL1H2S6kqAC3/AqFOTqGGl6GAnZfHbx0C/dP
zv9xacZ+wXfMVyykUfSQIWp3bha3BM3hXYVXtMGltFTh24aMuzc4HkPhSK1COr/W
l+KrrxtWP1HtQ3TUTAqlgIrV0AGixexexSZmeTBmHTT6uvRDwRbta4L79MdmmFlW
kKTT//X3dGD8CfL3O6d2WTFw/vyR1oalw8pu7Cq1VkU/P1ZBgaP7RKXcUHO5Rztl
kGupV7WJ2CFmaAQplKfJeudHpftyIEEgMLMkKTLbXYFa4XgS2LArZnOv/xgtDWmn
XGLJN/obbe99Yt370HjwDKxL0VaNXPc53BmSRdW38P3S6AS8wm7fW6tg4MVSrNzB
vIbt/VM8nVxZ3/1ZlxHaUfIiSKT4EWBUq7kZexx5vioOc3PJ7Ae+xtpaKUn3iqVT
T9EHPrnUFxupA+AetArfkX+I8h+zTT6Ob6fJDwAp7XzCuybVREPKlTKDuh89pD/k
6XpGx2jTQ9WgMN34YaAeYIGVnptc666/zRM3R3/rsW+ZiDaSHN8ZRJsbbOpIoQUa
9Wa1S1zMHXDhrh6h1qZeo0PqKMeU4VsFNMZ4zPYdGPUYwjk064a6AgBEdNFXtFPL
j8KQ3lQGA3s6KMDCid98ZB3QVMNejaZVH70zijNo/vLsotKFpdfdzZXf0bKGKDn2
rbuUtsYr3eFnF9OULNz/VRPhNVU9qvKYxysG8ykGSelRDdZy49pPsyJGrQjjtEie
0tF6tuh+nKPWF73whmRE1KjXbBC+QLy7RHzUHF9wNpYuvvrahjm6nBi2g+zBtRa7
m5ZJ5q4VnwhZCXNuZMvlbwgzVxfGxrj+XXj4PCwDi+5OZCQlCSJZDjhEgVYtKz74
QglN96HKZlrm+HCQKOyBei22aiMidfF/NSDdMyb7w0U5+LRz19JwgEycLpy2NKZQ
uufbhC6eI3HAOCt/TmpYfByGapmpDe+Yo6ITv3p9UQo614Kx4O3+xvOUj5oynhYA
sz3dDg7Shvd9RDWv7kBlAtGJEKO4/QL7iN6wwZfcRrDRf9l9IHBJuVey2gYjrpSm
UiDpwb76duwSNZLFAVhAXn3kYxlnhjKw/D0YJZZQxVw8mAYeayGHEgYlNcbrUY7Y
TLAzqXcs93qorsD919WP9Df1FrOxHFx54CEMl/p5lu1+I++HaNVwGMeNcRzlffhe
j69gzAZkwbZdFWN/5A6KpHm261T/7PTCtA1uQNGxhLydHUUZqFpMg3B+kYNPRZhi
7t4fStoeFAtm7lW3mSCPiROPK3UnWEh/kOSYCa1O1rV5kaJbOnIkzaB9P13Khk5b
0rhqF+lP9NATnNx3fgDP65rht2/Q+ZjenmUGNyajwxMfuUJUGgAdIMiIEY5o8WRS
qotzTfXqJ4TcQDdTZ4V6JlVeiIe+qv2abTOrRHHXNc4d+bwbNxTtCby0UoGTvw03
nDDDHyYc4YvniPoo+jaOYuzDXaQgiQiaopeDIEc/77mWTVSoQf4qjAJUrlJw05Wn
vSkrfdn9pXk3cNpexEjsfLgkX0VeWfC8l+WtynewshyMGw58aEilYTT9oG2FDOgI
ADGBfDReQuMrJ+Y/qbIYnmc2ChLGNfdOphCTAYrar01vo6pypwb3S14Api3gTuxE
gvZ0WjldV+hn/tkljbQh1NdQfONAT9UjTWxMERD7Pg9OuhQqxDVQPlmIRt733mGM
Y/hqaz/xzdA0EMCtuzI5ekNZo1kQNpwoT8xGbeFEfLSQnO0Wcno6wyxIbg6L+x0B
AQi+94ccPvL4qRc93IWUc8DCkqh2/oHX7bgp9qHe0As2mKPjrFvmS8p2ncqIMZuo
eceTgzYLn9qwTRTJZZ+mtWFJjSKJ6JpUnuJe8S1xR4aSRlJcTWHJmfkq5zavbYGD
JM2tCqjZTGOioeug0qiyErijakB45RVmiuzSUtjAoELjc+CdEP3HlaPCNI5B/OhN
uw+CMQV5zwFNHoiS/1McJytZUrxAaLA5A5LsRxO7ghXIpULcgc1Nfgm1K3sWlNmU
vVIs64hT7PVDyPdfUjrzoKiYiL6Ax4Tr6bFQYgpnUXW9eM7P3+jyYvWI1F3wSZyA
fb0uhqg4/v2lxb0VKsga7yL7wk/QNPxF+Uf3z/AGGZzRDbr4cB/lXAFBG2jBs/dE
HNlj/cJ/lB8pXaW7cG1Bg89VqPFMOmkSu0EDUPYVDB1j7yDQ9l2OyrXHb73IViUR
z+YCBOMu/q16RO9IPl/UGZRf6Wk2qzwMs30l2vWye7EXWFTuceEgkwY4yRJTM9DE
MbgZ1BmbTkH39ad3q+qaDdDm4qrbHsfoRLNPSJfgYyr1/ZVGUpwAGImaaHwo2obQ
Kn/nBMj0lllHmgMDc+UTrkh/eEChgolfQze9YLHSIdNSnyBuVYEqB6gjj6ppCHpF
DCPtn1ua6drX17JBFYivrUh/qgef7NFs/UzT5a/kZyJ9LpJXJvRvba7Y0SYL64yA
OKRLD7x/PMDNozN5H0lL/BqGsbThrtUOLQQu53oOb4k68ybI+k613fi9RsU1W9aD
rkt5+dtaakGocr2VfIArWhUMPkjfipwROnvEWhAtOm0KDCashUuClzAM8PHUQIrd
c1GY99RDj28d/xUz0xU1GNfzPx598aLTXs25WuP+15zhDZYgch3yn8U+fl0FoAi7
OolAQEcn/H80I2+hts2aVF1mCOJnWjm+RX2YirpP8dRNhxn3dXWLg2U2Hth89lUF
GPIyM5h5mx/TDM1vAoQb3TcrcIyns7ZTcvo+bPMuXqKZOOqdcT7FPo+5mq1/BvPP
eEwBmP1vpljhanGz6B0AWPygFu/TLjq+JeLI/BuZJwCbV5U42wSq1d3qJDIDE97r
lfrXmZctR9uM45VltE24limdp2E8m9pDFpvUkK8lxl3g3ZrB4q0MaQLS0SKvojq8
TedfUw0XOV6TTyboc0xl9QTTRzNubviQ9yvys8i1gHmu15YURS9S1JPfWVSRlBek
oajLwqorju2wQFKSZ8ofNi2FprKzr37Y0QQ6UDMi2eBswlI7BPk8F/KMX1qXrbE5
z4E4wE5YG3a+nCMW6xyqpa9wPF5nskfqQDktFyFqbvL3byQqso6hWmOfTK9Z2Ky/
unOnpR+rDbqb63NB944dIoDgk7AxVitYI3ufOCXcvyTlVvzp6ND03I4dq8aLgUtA
t5+n6aWaY5S7Duo1tRV1xrLDUDmXW8N0ehJk6F8GhiDIQD8Zdfk+3LCV/yBCy71H
vkQRYSv4qomNxPUtsafD8aDDcApRgqgcXCbE8Y2TQkHWnAGjr6z3M/HLlzy5K7xn
/GuS7qpNeUm80uqQS8mPdpfXBNKtXeK+KZbcoWp4k57MFpzJAhTTx6wXWg+KEkjC
BUZyMeoTsntHlxOHXL3s58W26QQqJvghFqkNQQd2UED2dccxY8jrM33vxERuWXgO
gB+pVbXf0hZB0lWaI5nShMIHmNv/P9cQFYFAquGDqSM9LUM0Cebk0WsNdnz3ics8
yVsTfb3ml5GXPJojNQbrS6IMR8KBVZ6wADYFhhuGW/J3vlJguGILgZm5qyGgLUEo
HjSBs8osAOmvUhMXduNaBlO0qVI1R+r5+EpdbwF5eHoheJX29ihlKpHE4qMt9e1g
MSgc4MqvnynxvVs6kXQY16KWgUSlCJczuYsXRxMyHrzU/4oK/YWUN+JcIM+WPm7k
2AJgZ+jZRq7OtCJvF49FzbK+lr5RD298E1Nqd8JoUhNDRyXHBPmibgJcedF6TOWj
e9MF/mD/vTFZX+aUTJYK2YBB/4hp61YESdaFxLIWmOqRIKh4ptJICVdkir6rpHTb
WmZ52gS2wvtki/qtjxCMQNlMYHjaKIfT8BJ40JmtsoFlmSAoYmmGz2+Kv/t54RHZ
DMH/IszTQS3OqJwgDEfKF2x1X2HN/tyXlEl1y4YcKD1oLIDdmqieQpLl9/5ulIcf
8+nDBlZt5yLjYJ2S4j6eYS6x+oY5xh9q7BoY8B2CO1SaO1xMJLAOma2tvdCRQY6X
FhMV/cb0iIiLjXfrhHYvi2aWfgDHLFBCAoBES70AcA9r4WeLwtSbsObpsn2ehMHf
IQLYqByNshbjYlfO3Kzv46EAspnsawGZIf+MAnBQHmkHZ4Th6k9NMhykI1R24dha
nher8ypT8nQk5P8GZMrEu9jCyI8/At9Mm8T9I+gsfS/hvKVp12xgB34hMdXHa2Xb
32UQNwtRkCaGxtvQjiXoxUdtCJIB0Rm/aRXgkNQUvmMZh0VtmkNeiUxxH+jP/Idh
KswJqgVH2MoMKKowte6l1gWmonpfzKvT/4NIiZ/BHQ0mlY7LBlrguSvrxroZb3nP
c0rsit8QWpRO+ByrtZbtBs5QP5AZwya7NQWToyGfKv+Hvfa3fpnxCcUtTCImhKiU
XM1PpVPqnfuUVINDpRiQ6LHOmtR7GSRFdEIDKdOxhF6KqkZkzr5HgCTLLdJf05Ab
RlSVDA1BVYEyL+IlUp02buo4p4uthzzx9vlD+kAucd4EiOiTpZhLm3t4caJsyCao
DSAiKqL/Xrd0nfbCVKs0gWkzb5v1VNOBNpXE/QmMzAw0qzJBk2Nz+XGEgkVPwOp3
U/6htRIVJ6/0LzT3YQOODXZGl/HLWFNTBs6EAPEBALq+TNlzt6F0YLqCx89gt5H9
svUFPjoNXKxBMkWKJiYazED/TCg6ofSTDLlY7jBT9OA5xV6lAXNAFSmP6APOCams
I0cEQPaQrbJSmjMlJm/pNCJta3jiZMlVbFtLKSnSedB9V+iqxIYvEXw9xdkhP0ZS
uwYu0o7n5mZYNuQi+9RLDGEIcsJarBWOMBYyPP0F+D2nPYWHoir+u49chi2yeIHI
bgFELEqgDw4e75exR2m3vI+Ohu2FzoG8zbt3rR+6sB03XOoLu5tl4cAXKlzlHXt5
KOGazyIsG7EgbW7/0+LelN+fn5XkYIR/C+AiHr5YV48bdC5DQeV8JVDwaG8jDXhY
TDU1TsRXePbrVcLSBpDekYkgLz7r0mO7H827Ji6bOYdN0cATu1GkxZsWxa/k3rAf
tEuj7d2kBJAFsxisdu4H6d2Vgnf52AlPl+jiy3FyAWXkglKvH3SXBA8AsGnzkkPf
p1lC7uIJpcswn6E9ZBv9s+vEsjZw7+y4E/hnMR/rOGBowCywJCvslClVlxFQ4KZN
Pu6q7UaUddqXgYHR660n6CDaIrYG1xJCkLDKQYmP68IIv4ND6pPlk+CbPCsHm2yF
ClKvDocc5ndu7G+35i1HAM4lG1ycX2LwubZGv0f7B0+cLX8jjrGFqq+uQB8YgcRe
QyUHpB9cKhjzXJ1z2C6AXZRvcT6bB5jzL/ItxSOTAJyI/yQxH4k8yb9zG1mhoLGs
H647otRKITH34Yn01HAwYoH6UdRzdLLllDcqOj/2pNECB7DLU4wCEooxCJWx0Fvy
RJT7UZeobhjK0ihUcQ1HE+T3GAol+B0sbB79jJFNdJ5iYQvACp99xQpJ5hSU+J9h
+DLIS0JdqKmWm87shD9OJdVjRLMpyBYiQN3tpbuBs2gRw+TRylowTr2C6W39W3zL
bz7mTFNXzsqETCxrQFdBuKskM4HUzRqTcx/4SMeEBTOPXtSnlCS+9lYFDt02vvjM
AWs/4smH2iWzD83Z9xxkFw33HqbcuSxGmyKHXhyhFf+lQZyJ9uW5/xeBN4IaXVwg
enZ/+rcCaYgZSQV+LDkhIwCbvEsRBhCSopsBQ+kLw28Gj+SfwvLQlv/kTzak+Qeb
PJUp8s6rJEhIs116niv1xhepmOlYGI8CIPQZFbcGjT0roVXPrLMkY8gKh1h9EbEZ
7nuMxrZbfUmjbgV3DJFCmagwxK/TUT/tHSTByUfJDfQXSQl9DMJDsc0ajJqSj//n
BIPZnVAugZM2/njzzzgmAglODdAL+IzNud7G50ppdOpdErKn/3BgK0ZymkLwE5dy
cmiaFORIyoUddLQLto4mMFXx2RY4l+fkmcqsl7dtTchU979CoQjdP2LR1jugcr66
MB9KRGuQQvgXIwc5F9KWo481nZ1K6d9ANqWYdBwkgkz03K/RA4EJtIovilOCtY+Z
VvGO4pzAJwUp3k83ZpxoPdDGelectojP2ZDpAlsACVVssoqsxL+aZ0Q997fUeMcL
lulT2dSlmvFnCWjcBtsoGhFAthqCc4oxc0IV548/ZrI7aVrg2XGD+4Q7U7YIhEVr
K0zXZ9sWfWX3sBlOcagZA+nUoY/DK4TKQLnAk+zWd1OmKrFottOqFRF0KIK73JWS
25ZExqgR4R2bgV68Yjxp/2l3cMYpsLrzCAK/oRWiWWZ8vhBwVUWpmR6ZPe3PDVwF
K7qBw5eaaATsW97ulq8XmB0taTKZW3qjjud4mVE1BuMNUVen9lxpXB0sfBykGVlq
icYKfyYnvyTKzkCCaUK4YmWX59ILVQG6chwvmPQcdt0EA9PtNwbj+tkkY0uY1+bb
0g1M9bW8BxiP+h/joRwfiakeqFLBTSWmf0f8U9gQUYOWkli3VqimdaX4s7FO+UHo
eNkRwr9J3mvygmxGcag+LWl22IEdl3F/XLfbXkkspNxis3L5BTes9ldV/3oRQL9H
ZS30VRsms+G2bFjmgHGAIVq+O47OBEe4TH30zT5iYS/0xe/wOeEzXJDYxC/x19JZ
z8cEqtkMRu+ZkmZGAoA+yoPsKw+dhLh9fJHbi6WBiMqZz4pALNX7JBRMzDUBVS4N
wsLryIQiO2njq86cH2Aed8wsv8uNVRbpp/J1IQzEAHg1pDnux4ycMBt7sA6DBU1W
JgKUK1rQd8+hsN5OlOBM90zjo0hg0eSYU8BFXNNadu1ArLuG7MJVlOeMdPZQGtFo
XhjdkLpNiN/co7LqWWyrObpnw3ovN/4iyDvapxG30tuUru5aFR/vMRZ04yAq8vG7
na55pJmQNi+B6SPEraSqQmxZrdNZJhCIxTaHPWeXV1VUseG0Ph1qM3u/nRFvBEpW
Q2lzQid7SBZA5giWwjUB2T2Pi2C+jEpICGBafeMpnesePZeZWB0W/dseCVf1eqH1
/nUFqSuCUOwZj7qw5ROFS+zE/5egkSGfd+HnS6IyQgztlCuh0JpRvVDDc4giNpR6
l/r9XP3TWhkXa1cbG4ewM+7mCoDqn05Dl9IxXkjBHBYfogUpmpS4aVbKV0EiENrb
DpuwwJS7nmUh3y1AqWWLVIVNZzcvVkaUEXawTyyBwKcTVUHoo4kAkzEjrhou7lPU
Rb7nPXclj0QFcr7LH/1EaKR9wOXytQl8L94ka4lxmibC4nu3SwC9+jpk6sF1Uq0H
EKc2odl9cS33UsPQQS29v0IbOGXhwVPnx+BZnxXxHzfX6b7nw7moN9tDLAxbzkmc
y1trvAP+sVh7r6WrXQExG25nPqOUWtX+eBtRXxozy2n8/s9qmAPdymVzIbFyw5yU
nwsu4jzfWv5lLT5/UfmrSjaCi7FyJEmsZYOnmMN0ahEcFjPEM5zkwRQHy53sdF2I
3Q+2ni1J+Rj3EgpayepECWlQrDkoLjBVzJ7Qt2zf0k7mzMqCD+jyXUC6WM8e1TgR
2JlEHI2AhN4+oghdElyjVsXIKgbRvLDkqGnLMNhfq/8nXJoGfvoEh6ErZRoX6X8a
pJu8rwLBYmzPVGfMbAZDjYNNUWWXuZt4ZJEUx1N/qwsGnrgpwOph+WBJx6abkWhU
mvRQjOSeO0/n4zVnh3N6AjDroVVFD+ORP7uItgUcPm4L4LvOOby4huhQKEuvBenT
2rEQ/m+fi6Eg1lzc6Jz9ZuGykBw06i1shaVSHm32/WVu9Y9u4Zgh+2g44yMX/2jO
2eTU1ZCc9SUQk9WDzNE0hpBtHNW8hMc546o/84M4yOKmyBMHqdvZvQEsFhXtdycm
cSTwBND22aMScOHCMKIJoHk6rEASr3R/xKwQb0pc0jJJoNoarEzlucEPuXjiM5Rc
8JxNhPFJSyGDuIb6CmXDpXaLD0toG9E79TmBaolopF2HRLtgQ72FwMoPvov6OcoA
nBa9piARkJGJFwvEdp8zWUztWWWDLaWSpk3tQdxhiQg0JfND5zbSFqP4Hbpe+tNi
JZnV70n9HKIzVjDV2+5mQ5sJQu0YEZw3l5S9uRe94N3nbLGN28BEzv5sRYZBJZa9
Q6t8Rn3sOpT/NEqh/zFIl1NWIWSv41lnMsn/vuofDfSDTF+r3IqSU38KpTq3cTbu
LjgWujUTP0Mm85ASPvG6gBp6ieNLLhiD6DPP3c4NXWZ81yBvMSd4JqesvqDCGiGw
utr3PwkpjjReEBFoPCYkQqPmr4xIqPC0wcoGJyaQz469HuG/yI2S+5MtzNq696Ss
oyifppl33LhlyOfmawGDyXrflKbfoqFgoSjf0sAPAWQotGobSuzqtHAXmjFa2sFh
4pqCBdAORfhP9/B+ea85pFSAsG5wll/xsvjGtdd6toZhurP2ApC/QuK5/vqLs1cC
GcKzoCJhjOBZOBdsE4Y1L7Ot72VXcRKQqLzKuPlboDMMIXiR0ffZEZKjhS7vFZTU
xw1nzZrgFGP/lzm9jA40NkrHoq4mJgXVIuyZZAjYANUSDHI0vdD8zUjSFnN+ygq0
EDkfZu30ltMOHEcYFVEY3GxpzVVBB1ngxuDgDIT/LlEGphKl3ylrvouLCQR8mnAT
Oel3OxW1vYITuf/9otWgfT8OTsKzRWyI94tE5qa1g+HIjGVYgRsJYdCTzqssJmkU
Btb2W7mdatZLR/ifBDEl+WDNbBicrXpguAgtpNcYKbEhUF0+HmTeYppo0yhYyXS8
FyV3KGtPNMqP9029fbbcZGF+dh9yqTMX8d9rPvX8qmqGCl5o9o+t9ZqpKUEKStNr
BrelVXMozKRsAj2S6srbh2jZExgrPBbjJNPrJlPr0m0n161y5Iycz9MhDhir/iZ7
t+5CgxgEW4z4e+hcDBomYiVw8L3Ki+JJzDhX31i+PU5/YoZLsj+QwICBUXbPkbT3
/pDAY40ZV6hlFEjYnxwLMRMA5jouvcTwZjnE5Pcw+8OfqxB18P0nW2lQjR4RvjBJ
YETahl40Otx0r1VVian/B23PmhpcUcusuPXM4BxDHvQTNvWsJYWpGDRI2051wc9x
XxgFR5eP8AZcECaTzlYJAaAlkN37V71exzdRUhiw+5OWin4e2MHzEG1hzJN8z9lN
Rq/q3XLRb2iS4GUlcWUeruOwHq2yzH5bl1XOTkxC+Z0uteEk7/ke2PhZ8H1eZHyN
+AS7xK0ma4sOvtVX6fgr4DcX1JkwM5WbuN8Y/+o5qK3z+GQtY/Om58PdFPT2fbA8
tTY93ctwK2yzfk6lWcy4NTslI8+InKL3se7S0eOOkwsoqY692+pDxQ97TmnVvcFh
kcjDIDQ/E1a94obz15fQSEZWa5rnAlHOjUetrCxu6NlLRLcbgY6Tp39PpsclEVdr
IJ2Rm/Plm/4aMdGRKd0zQT7JBGoiTnpc8dere/cc0VbCbiLFRLoySsrt+xJ4tQdi
91BtTA3ePE+AQjyvQvfQBOqBsfu6jyR8Loxk5VtBc552wTdZvUfMiqd/gmNI1WWz
kvFkxri/R1rZzASuupnP6BpVeruWDtnkRT/YQkVayOEVhOLDS/mXzk+LWf6iwADj
3JvVrnfEa70ck61+aLKnD3ZNiFZ0RMlV56N+tPI8sww6gH+ygz1ZhY71kq8MI8yH
bMFG9z7my5NERI5G595DmavFqAVA/pY8RDkqYXV5c+3Fp5/+AIj1jo/uw9lmN+Xs
SVuf8HSERuIEzNHt+Cd0T+6gg2fwUDzy8ykKD76vNB5nX6XcmDgiC+ycEAjp4ru/
+yfLAytuYVDqza1meZL4NX/wzn/eftoTCBEJjUrOyyZjmskAkGTrJqBIqLnm/mjH
JdhStg12h1p5y9Wimx8ZSTrBdvYG/7Ij1ji0qnTcP7rPGc+y7AFoMmtsMVLSGG+T
OwfWGb+GAKENaVPDWGfVrVC9f+2IsavJkuvzfZg7TfHJiNBHBzy9IxB8FxBNJFcb
aSOte3mV3Y41GK4pKxUI7AcZ+ikr85tWQWmOi4kKdTnwKTWhEb6nvW+IAfD/PDI4
yS5ZtQyJaYl4MID65TQ+uu7EYuY+PqVVkPnI81kZePpU15VeYbi0xGKSmlcgin2F
6t1RAdAoXXBIH9ENXt/W0im3moeQvovj6Y5pYBq8t4N3y2CVKckwrZurBpHX9I8K
ErcXSb+VgbXb6Ain0FfMgdXRf8Piygdn9B2ipbOCFgJFvIr+4YDFoxIVccr6NwdV
xku5iw+lf5G6cGZ0InYWgU6TEJjnDYYXI/rStvYUJqdlm5COlenGcMIwy2p9SLTw
SJhlXhOOUq4+M7BFssJPnh6J09LKb5woEI6HZuuC4xtpaMJiYtP1IxjnOb/QTZPB
GLVL6bwUvG4sLno4DmIrFy7BXbJmjGhTKITTAzOwoLOBPoG5HkEvXahbRXSjyaaR
uvT1PfKtz0a4jY5h/vSyslP7eOTa+7MBW7FElsldsxvbA0Tfiy6GOdjiz+mjskJv
liXHTRyszemW2EyaltBSa6ny7z9Y7jtRbAmk47oDLIXF69JuyDYmhYCBBgXtRInZ
7NgqsvEsxbqTL0R86k+PS1/sgckOaaOaMoyYlNDwF+c+AYd+PYCna56Vug52FYTT
x+mK8e6vY6WbNOyg3CezxL6Fw2N2uHszYrsY477J9I4+RKru1J1X0pEkzuGFjFu5
3yNczm42pC73pCliHjy2EpHQbmEL+CAGssdmTGrMGkYZ0NXq8oxx3lqxC3fk4XIT
7GXyFejPihQYmJ5wfnal04yoK/wO/NImCUuXfptAicQXqDgELexatLoXUUksYkzi
EEERq84fqvGQZsow+U1TTrU7ehrZC8I0oDBC6YAqNKyd7UlJv/82PeWXXn354PXA
l2nMdlKUdztHGcOa/9pzGEm8mvZv359jo1SDbKOSzu5D+L8851bjeWoCs2up/glj
Z+OFPBZjX0T0OqOqYuDfta/R2mv5aNN4EVR7+W0CEQk5BIU+GecCStSicOY5GGMc
miWubXPsBwnOZSsV6SIljSZHres+d04tPKWbdD1c/Ekv4LxnlQYwODsiYDVczbEQ
KCT2Zj7gnoiBXRBod9Xz5ryGaE6Y3XXLFpvZeeghazLInPv5MSl0tLIcK0akYz0Y
pL9rJMRrMpMwnuWTiBCTVCx2d2GXmAn7TfBE/StDZtEVMuw0P6e2uURkbPtNQS9V
5NcBELaDLkJovFdHTmsJ0sUTJQk4YE9wjr+4nS1uymgOZk+VgiXbzNYibh5qpP7y
i74A23WznXui6KLRjXf6OUxUwNiOiLqsOtZ85Q1exwRn8FYz+LhgkuqheWe2jpsh
6BU+ztg/P9FRvJPe076tKfUXFSB0RJSY+q8TeA8erR0XxQHWqr0fzF30nKBFE9id
FJYtWauj9j5i8AN9vPVaEQ2blX4CfyCv24OHhTCDEt/x50flYe4KVtK0AGP8c8H6
EcjyJRgl9N2rjD+FPH0ru02SoTpdvWozDp5XabJTnQq3i5faJI2dQcTMxQurSjiE
DfnFeFkgT0NtWKpharAQQWW3ioJq2ASKyVli5frMTBx9MQ775Ot/gd9qRTMIZUf5
5eDj6ps3k4uFJQBLwM9eWfF4wPc2aLAsuvT2tZXgN/j61tKJ4w2o3tV9rtPL36RM
s27D6GMf3wcZKgVJE2xFGLgygNK6cVVIMtkW7aPRox06lEdR6WaCRKbbvJSH6sR4
ievjYG+w9EZy8FWT3eUvdjISfHbKZknry0D0SHCcTWQCyvON0TstT1TlSdoxZxGW
O3bjl2L27ervLS9nymsLChtJroj2HQlMALJs65/WQRZd4PfJF+NNUusJjdut0X0+
onRpfGVI7fgZl1NcvTrYZGicssBU0Nzjqt9XOQqLDofyDPlDjpPCCFWPaG/E2JNh
uWmnePJpUyJiaStWq2BbGlFpDV1Hdih6l/5FtqXl8OsPUuFf2pbAqREqiJ3Zfurc
jeDaWldqS80P7nN5h66Hlctx+JnFz5Wn7Kzrcw8VUsEy3j8O7Xt/ubGX7FCjyUDY
hQiFwZ9LXsJM1xLSKBenmPN3R3DXDRzEKgC3HmXivHhv06/G2soD8K6b3eKWAjGA
nCS0sho8jt/uqVCHHS6yr9ivr58CJZHIEbBA+k4SY1ffH1dyyWdw4ix7rDEZiRc3
wMRrnY1N9erTJO8hJSAC1KtgmmkIHr57tCfXsEYGRMqaqDQslx35ykdnmtx2+tRc
/vSMGM9rLC6F4W3hfqaWOfK+RXGr/HE73Z0d6JuvpnZj27c8RKLBS9iIAxwYtKL3
SU9o0Muqxk0TS4LhMr9v8w2UEOX574t9SaKazPJLRMbQe7SddPJ6AqVmD77QK5DP
qmtjM5+3baJbsgeXDx0p6SwP2N6xoQ6gGPvSzPd0SbOnn3VcFBXQeK7cZ+2ZrFco
bJ3GXJKt2uQhM90vpcPrJg4TdVkBvQnZBnVBaHLY9mdV5C1DS9aQjTCUBhZrOq0w
A/GscnkZ122blgCUSJpLYBPf4DP2xRJM7nHhGiPJIsrGzbi9CSFcD++DWt/epmRk
Whqh6xZcmhZ0UNNNM/APJBJNo+P26kpTBdnWv3nPbMFMNGYP8YEE5AS7oah2FpdT
PshhOXjkV+O6WVTjai6JG0LxIQBwFY450Q8ng7SalI+vUSh2NzV4R5+3R12O2cUT
s64yVY6LpO6ZdIpbnG+QOaKkjGDjuCqLgfsM2c/MJg2VaoLW2/uuBATjlpo3kRwx
2PhQcOa/FM5HnCHxmBc95EB4fgAAlhsSHlgkWOT0MAPU+uwA7MWyFL0EnMI11+Ui
WnY7gD6e0B8YI+phvtJio7OtYPSrX4zwfwOg1+fDd9MybglZp0J5TuYdnKzkAC8p
TiffMXw9qo9M0ykbJH3mo5HCfGYMm/sJIh6h7KVlDeko3BrTo8biChdg9JOK9X4B
i5qSyTK//y7O5Iu08x4Kf5j42GMiikLOfcevy53iLcyLOO4yFLlxKEFr0fXyYbTb
vICpA56aZquHHALLYfsIwdoPo8rhu0nXL+uAmqxLBSaLv8O3m0a8C84T1D45Ec1M
NbkpkJ/NgVuHL8H49SvJKQ2E/iZ32BwgsKn51E4Xo5462TPWCnjzC+IhmrAF2kWO
N/3BdZKuB/AFKFI0iCzGEVTgu4e7R87hDO2jreTD0U1PoLZPTo3ZF2Rx4lqgxycV
vI6cnOb18/W6V09dxtzeQQwZhWG1Geq12vaGnLBVjhfP8xrDj+/6pruFUCyO+ssf
v0GBAFdcz7vj8cNr+ABrCXaBCNYiwj0oqEd5cMEewXzQB8Qt2YfTbS5+RMbszaH3
V+gWCO8w8wdLgHKP87sBvJABRqbMJG/0klUkXjmZ3HOKu2rAVDezv3BA3Ge5RP3l
zamIXNlgcC7utT6jOAOpHNIC2IjpurV9++vatNhIs6lN2vmcsfYdjb23Phbw71ac
hYeveP0BS46Mx+vKTbwJyFxYZ3uDIyCsTnTUAg4GzOxN0Jao+jHhRBxxa81S7Pvx
TKRO2xGC9SfF5jjunT1mHg183Y5nx26oe3mk8yt3b0T42meBVIq3oUQoK1O63V23
ziuw6LSWTqeUKn9d9rz1NA3/9UySbPnqM05w3USCddnjtoIJactvOWjfQxMvm3ad
z1oWX4E/iPq6XLVDBNDijfrS+I3kKDGORCEsyVViwxmSjberOtwAe8YNPPOuTCQ1
B8RG7QMHkqJ5Zh5hdx4ZS7zjM2aMNuI77HdUhQalE3Ns+ZLLfDXnntsl04FOEaNE
YZy7dU1wbMbpaEvodNxvL0CWBnOabxlvbVp8RorBAabYTdetNl73eAONiIwqaQDP
1bYkjrFEbo0dbLk0e1dSyl7H9NO9MZmaClkkpaQSdSrUb4qe3hI6Y22l8QtX2qzY
wM3PxzTdQeVfpFFnT4TqQC7FO6AbPwah5fgeTdOpB4DFFmKfeEq2KSx/U/WqjNXv
vyIS9Ws2RmQk/djNiYs0KEOUgyx0veynJegPEGzjYcjy68AjYImDH2Y7NFhLMxul
nEkwXdalyM6iBMtdN/STOytPUihVm+hxh96i2VLk8OkP00tHS9XZQ9d1CKcXFzVz
jXefNb+I0HODzozjS8zbndkGuNR7DDeHtRkzx3b3pTm4DXimAURnWqJho2PUfC/B
YhaN0gRGOssRzJ+bznmg0k9SGpHr2A//C8ZjlEPz4DVT/yykuVMeinsULPClab0s
opsQSg7h2tyiI7zWjXwMveM4emkXsWlo0Uaz45zrkR0qDqUwyKXp9wAPmE9jnNyZ
s4W/orZKVm0VYwI2QmNo/CTCxh9XKeb9mJ51u+lkXNvFvhBX8OdT59Ms32PKp9gM
opS/lZaTxVx0zVyUbdpWZz3hgLzucU2sSs1OBqIxcI1MCK/N9cQYswkbyqmJQxyh
4T2/5GmCOalPRYk5LjGv2WnRsqHI0x8zPc9HEUX3cOX+k95LyxSKu1jmSmlECg/I
ElZgrThgQwgImAW3mvi7GsmvQMOgzqRkQz1yUc19KrKU5jElqKPNwu98YPGA6ZrS
UhMKQ3cCPsYGeYFlc6Z3Bz8mXRfhiaMCkHu44X8GZYCBGYJ2ovpPke4opKRioXPX
1VN63TFl5ZjROX7lJYeL/ItB0qJ575J/7poNbHwgWDmb2OArEAwc9cXFnjYYUHNq
0xxZdymcQl1SSr/Lc6vlRIAnLwQCtHA2RQ3EvE6RPADZt9GijTmLuCTMPSxg3G+Y
+v6N/QfZDLKVNOLB0mUJ+ncN/sihdC5E0Noq9FUXXIYQJHBp7qy/HoUjan2/igG5
LeOzdUVS1iEN7bKYgCtzwvD4XM3FmOkrC8FGKvtbyWaiW3h+5xeIzJq99MtIquZr
e4IQ61NuZlNjj6GxVjvk0XvlyGTI56k8wXSDKYpS1Ct5J/0JHi72Uh1YW0vs43Am
z2Om4v6R7BfN3Pe6HzCCwk/e6bNc4qDG4k6gSmX0wX4FwW+a4dQhRcWQH1phjqy7
146Eby03wrbaXgBr/X0ngRYMkLttBxsKbgTqYByaz5W4XsWgOf2kgH6aOtBytXCc
PVLt2mA2s+kG2yca142rsDF0L28EcqpFImM5QLnl257nfR+zA8bTCcHJRyK6dkkc
LldyIVa+5coKBtcqWGvsfotQTIV6Ia2IY1uVJDfnUWTrWWDg8tmPlw3sbgyCK2Ux
SN/FAC7ETHuD03SGYx8exSVBo29+yl+eQ8JgXFeOuHTUAUm1zHXrzJhggB+4LaQT
WuTM+o1cyattjEfAFKT6X07Yi/9NlxuMAmq/fZ/1LL9Uz9Ha8q9DozlZGpzKJcQH
ojSRpIFJHX2BrJbZj/tb/Y6rjIAL+hyn/DRs8gQ7pHO0XBy+tjyCZKW65FYTexvi
k1AolUsZEik9jgmHKQzTzDUcQHWW74b4pq39Jywr4GfVHfcVNquPDs8Hi+dTE8Oo
/6DlsVLNpcRBNGmuvp8YyZ+wng7bEwRpyOYjXWYu4262sRwkyqaKZYDrl17ed6Dc
//qtuX5s96mCGkmhcFV8r+ucWQ9FZM7CQCLOzHLTiH5gc7Ram0ad+Ds/+MFhwmY6
JjH1aTC9pqjyO/Qt2/GJD6U7y7CSOSlT6uQ+SKVorbCMx8eSjCHm+zrvyMn3KfTa
TjHfejiLmrFfLnSpzIfTvm/2TGBw3UeAzMo84jfBdpFisuH4OBb/8QHf3qGH/IUq
MS4TnDZn1j6W07u0fNifE2KCMyOczzAchzTEFMUeVN5v6Ia/efqKzdUDGE4jzslg
ZwwSQyT92t8JX6z17vHiesLZLurUImvr5NsqzWUHmW8v5LQM3Na8yFT3VagThpRN
eIwcw7pPwKSW622e5NmSlOrtiHrWlDHwoGwxag+620WiOk8SiUm/oYwZAdAGXyxl
EZHtE+1MK4vGPfmI7QK+XGci7LE2Yn9azU4pG/WZOBLLNiHl6IgkGxwgPQg3/N69
w8N8yZ/vT0cYQ9yIKrR/GaFFp/VCSRlFb2BxjJ8FwsdwoYGy3o4OzOrwY1Yqvxbl
NdDXQAhoy9Fri85uX/XkpNzEP80ulrqTlS6PqzPbyOFCM4dSMgmy/RjHL3pGOIa1
rbbXSd7TcTg6cT1Fofo7nEKIYD6QxvhB6L5+SSMhvs2OhY3wVFNan1HejBTpr0sC
xr22JC+AVq7cIFKbTDi3J6GzxmCEKwNJPQxBM7EN7mwOO0oDQCjo7K2LEsiSBhSH
oxWOZtnl9wguKnZyU6UXcJ4zBlPHyoznjfXJg8A1IAj9QS7498q5lCQZzuzDtznU
4Nld1anEyNG6vwZ86Ie/Ti9OGfuLqneGOTyrGYHz3ZXtXlwAKW9Tnzsv5qUh5qCH
yA0jhyoySbXhET6RpyTrJ4i+kanSDDNiC1bNn/rzJdU/WcYz2BV3/Ak3U+4TZBEm
6RgEI4yGLmK3YfRJQdIb9Mv2wgbv6n2ajOgBa9m/aXpGik8YrDfct6xX9pVAEf1q
L3hLm8rLAVAYq0zqG8QHazTOoZYvvQ4itSJhOSE57+93mL1bbhepJFfgQyKYaPfi
CA8KeVFIlBljIbbFdBC19hVwTh0y3+Rh6jcjc6PDALRpDHDNztlQicA9A4psWLit
RHS2BQmTSlX2QAuBP/LqlGhfqz/k7zwnhrMXDX8ffZY3JAvBrQNqwf908pXM+lW3
XFDqNmCvKoxTdSRg9Nvf8hsSSopIIgmHNiQtjZSCaPS9T6KTfxSp9WioDIkYwdUD
Jz/uQ6m+bOwGlUzYM2SDppoGaqcsBH15Vr8P93muNRzl9jAqO7Fg5LbKE0eXDOax
HuXVuskDL9zFritO8skxg62NdAYp0J9ghMahdzKvNtR+FkBQnhf8Uk9SLFhMbZvq
u2c/sxRlIV1D6ZQR/wb/tFUFtJLaig+8a7kOanl8Vjih0wNeBuX9PNye0pidV5jb
j+ecTvhkU5LuEOxzUhM6vKg0QrxxAzJgaWSwLKElEfdSgKuL+jvszcfgRzj+rJ72
faJqM340BoEfurMXUcf+OxPdCeq/roYSIU3X4/x64vStkl1+fKtVAuHaV/vRyAC2
0rz3rZhO4Ry5eAwRKUs5P1ysVpoUug40b70fxTUCzs6ZnnSgXDXvOP0swRPq1ozT
01epxSgwveWDsLjiOmoUFlH+iyhsq1bC90mGnK22K2zeHGRH03id0GgO3RDy4MHD
wNDuUx9GDQx43mc/qiorqx2fV814FKTBnmS/68JXiTPX7SL/qgDKFWsZ2k1E67tY
yMicF6jWovV/YtComkdHt0baovAuBjZnZabcCl+iMvBys14WmnGkZ04OnKXrSTAb
s0rNIkSbmiSZ/+NreQ2bwtK+OvtgeFFZPCx+duLzqa8vFqwZumnArl6hyA2Y7hYu
wPkINWyj+BRk1/2BdY8f0gq0B8Fi59OonXeDE3TJ3VkaqLHPo8qjIjmeX5hpOkse
JqdWf4eZv135s+PUmMgsJonSWGYUGp8XkXnv2O18JKUXYixb2NSVXg2SfgU9Lw7D
5WosRmGBWolbJEcB+WxshWy84H54O6Ay6zU2lvflbC8KkeLxCOSYe/veEqFwDquV
Wr1zgI4SLZrgjbSX/I1ILd0Iq85GIOUkq8z+LJoCAOpSqkYT0rkOcXwMf7zb7Xx7
PJ/el+UpdWDTb3Ark/uDCoFR6G3VTJNhO3RHNCyuVWrI84m5JdsiALo/p992u95H
w4cz9a3kO+FAcw7qP+2OQ+VvbbnZNT7fotJ8RcKUr7hutMSQlczqrcQp/60UrWA6
5Ruh9jDwKeDbHnZpAiS48fDM6CXvK6DOjZbbOOmW2lE5etF5SHSVcTTmbxE8bTm9
vhRrdMoCI42SZXaQf7DqyBROIJxblmHldsWe1NT6zgLDsfVzXssd0hX2BA5ZiW33
+99E2unZKWyqbcW2WQNtQheRt5x7Z7J1rDLbJZjVpUnDfFUyClODLz7QKBQb5Du2
jr7xyKVA8wpWKJ16YNFJfWKTfkVajW3NNwemh8zdQUUJglQ7+SpXfLNoYRXzddTN
oKFRTbgQBWhyU4cmm9gxXMU88sBpUFaTacD58TDQerah0NUiUCSAuPbae3Khl7Ka
P/ZIAnXI4ExTuZUj+pvgw8Ubm37sXnxzuVOPp+wTn3pCDhylPss/izrC4fejTUYg
qwa5gtUMLO++jhQRmAJYY+a/LUR1DCZG4C80bo838pRPA9zUnPLR8NZ8VtYz7EsN
oPpBfYnPhLPYZ9HMyFqh8ldEQynelVuh8Hvl8wA4yPUvUBJg9Rd0zSzi+QrsMujj
BVnFoBnB01VaITAn4wKwbkblLMLeKm4mi/lYy9QjLl9eAjSkVzaqPj1E+perme9f
oxaaBe1AMbFcbOQMlYRHmevhkyjitmr5916Dm73g0W+bCCZW9Q7jfzT/g6xZQ70Z
KBDRru4PcOdDvZRo9D0QxTqaM3FH2kCG+AIM6+CrCBkoU04TECX4RagmkxT+MCUI
9wlhLso6NKhq6zYB3lshBUJ/bM7ZjGKL4z2y0GARfR/8BwjaziR1gO5lYM0pgmbv
ZtPPtFQDRjbMyLjst8kL158Ilo2GlV1tr/FzYQW/HBySAf3PKDGGLt99ViEgIt7R
XKDzVGFeWyLMRLJVLf2UHvXtLoQ5fU2CDGIKp8y6Yg3q3XJorIqo17ecChbpZfmK
e9xqx5OpyCAQE69EelzjaECJsU9g39Cw25m5gAifBlWFOUuRMLIjxokjySq4XCqA
b+ck/KlK1G1sTR97ACUJLI43NnyyUYXxXq+EQPN5DYaxFp0wW+z6KH739amATOjq
8thrX2f/PZ3X0ebxKwuCfctuosyqx123LzfIHv1DD120cYbZsz8wXeJNvKIYWJVE
E/dt5F7qCkOV/pIgyReZG8lCdlBH1ZmeaH/aRjwDLiAp0LqitiQgibZ86AWtY28z
UTyDGD4M021g/tvwHAzYWbNJ5CZCxIHIPRTYrtpG580fQRjOiTginRh9nAPXSCXC
C0zV6ov+5Gv+b2Ww+gFXxrrxOeMqXzf7WhbneWOq8PW3BjolLlk3ahubhZsIv+8Q
e4AAYiQX7Iep3AjkXumHc+hh+g+UqbWSeG1Kwe6boBIJCiENcZZiUrocG7pCBgE8
QhPEnoj/PLw4dLyfJtYY54Zc8CV6TW0YzPcJWjAAD2ezkYU45norCvNljgfrDHOo
VurI08ip9azF/9IPqGzCLcff8/16OkyzhjM2FLIZP8YcIdcTgTGaw6gbBljhkw5F
ckknf8sYq+AcEXrRmXR29ZlG2kpBCuewpVlEdEr4IxMTGvoQSYBBDuEldwJmTtIc
ybFgaQxQEXbkixPF0MSOJiH6wxpq7XPZWrTYUXNIZUqVp9F5/LGRXkRosGw2ZuFU
YXDPza5igAdv1+pAzf9/QqDQe8bkVzc0YNhVVoVMjIcSukeCaGs1fSqpHxscPmJz
o9yZZRDM7aGhYdoTI1GfEhe2Z3gFRSFbvVKOPoeDR8J/W2FakK3MGFAi0zrnTKtt
IaE2otF8K5b7fDUV7xGTxLyXZoyVxnVg4yX+NkmCtx4fJCXQCOxN/5R4pT0DEL/a
sTrWGB/JN4PrUm7oKVfLCEwUMhjXGD+0zmOsdEVx+ifoXZo6Yj+UsqcgkP0h1out
Oq8m7Y+utE7jRgYf+HmDqJRIVNFTgf8Sv5cZ7JtHxUl2T81AI1VB/LXA39aMuWgN
cDu6xL5+/6mIygOE+7FShbyWogXlkybMVikkABLzYMiFZc/hww7BEFEsT+Q/YS48
qckW9sctdujnRbwkokg5QNW00bXHjNhVQWb2iZeusUxet5DlTFUtzIOaxfi/iOJe
o47pWq6/SF6xR7aAk1KPqxogq7777jxqPWUo6NBWC2bjSVV2cjpetz+jWdw5s9Xf
U24cr4SBRdXdvco0383mHZbHyKzV9cPgmme/Nau4/xfwTPvRl8sUCEZUGfcN3e/b
sGw6jXVBWH7boyCid6WoX4VDPgGXKxhkaLh+uA/fpdYg7MbHnljBv/pVdsl8eJEQ
2uqAC2zMl1IgEOXGLVC+tX167TGgZJtoOnSQ9eCt1ZDN9Y/HRaUKBTjEe4cnRHi4
b24YIK15XPSwU4xUOvbPcJp99AvXooOeMunmaLWnELO6aRu9BldiW8gNXuott/IK
StVZzAFacDiu4hBabKRDeuTZFFCpRoeN5UKIrY/s7X/r8vGhzwD12OL/vQbtCa8v
PmlZf2d9TWbGoL9uaSdg4YC1zN5Jvd8V8HQf5d9ZmVDrZTrLQ88JoaIJ/h3V1tFY
UQGIVP2GQ+ZS8g6JGBW6FuWL0iM7WW4RBoAC46uGAbMKK4Sd5BqKp2VHwE+E9evj
0jEriRfm9fZbVgRi3BRO8QoH+rGGgPkEalQFcEHpLQRgmdDpTwmr9Gta0Am/RFmh
13HgsRpBwCSMLPbqvSVcfAmZddGUPaTUwv2OTCSrOAS56xhGawgMDYQHEM9uI0UR
yusYRM2ucVPTW/G6Bv1Nv7teKsDGPzk2WmxgKUStb+RqSOz7hzYlyWjKRwuSG9gz
V95xJ16BD8N81zYtekeVSu1NmadKYZr7+IeC/LC42NL8JeAqZ/uy3MRaLhNr/c3u
VUQ/f3it/8Bbtkt+EmJhCVTwf94UDUdYrlRtwN076+OHlckSiGeFnVQIbXRddYFf
51VZ0zCoyXKFXdw+eMu4PKjqtp1rJRiKbkvR+4Rye38L4BdVk8YSkS83it3jPRYN
gOlMPlRs+qjocLM3uF23j9csOM5d1++UbL+XoX8/jmyTLal1E7xrk8hZ6bTMtb60
ox2JHHwAWdTPJA83Eafalz1P3JFgTK4eFlUW6SlpesJwEn4SZWpq6k03jY7n2z+3
5aFLjtisw4D4g9ezn0Y1zXkL7PC3RSqE+QGB8Kq63eMXutjj7CCWsBT4EXZ2Gsjo
wugLxT+HulyU8Ht5EhRYc5CLQK3Hy15LuuHfSzHjtpeWGWY4CPyFtGzt4P4xa1Rk
jySRx1RhiGtl/jg+1ledMvG+ZO/EDCx43EKG4ILhxA7Gpf8LVq/j1ySJh1RAWfSZ
lJsdwmIPIqqVkkfGlFn33heuGFp9o9I/zPhVqW92Q+teE+mWxxoE3CW/QgUChkcM
jYtwprqIB/Kv9fcasbgnF/0+hdoGMObhVDI9etk0TGj9GKtXFOOxkmyMyUtPNuMb
rumD0/Xa7rle6WBzIStjK0id4VR98cHUG1/IL/tnPH8KgMqHq4GlSm4+ayEtPWN8
uH6r/zxFb5hnyHN++6lewSUpu5rIZ73OofxzeSxjID6+IieewfdYPDHbYQDt3KCZ
0SBPDUPH95mFuITr2xpmCCyJf18uPgUVu+yY5W0ohMh+Wi5vJdo3b0pK0r/cJKRR
nCpd1emJJLd5bll5zgwB8mlqCvlGOY1HmXeoCnz9X21fMEK5YuaTwKMUVPK8uvGW
pqmX6TbdBiHvL234mmc+JV2Nocu3JGktOS38G5uo+7ZyjITLgImu/XGiozqODRmC
3goLplPs/vKabRlj9synPookA+1xGGc4vNHqNjjnW/T5yeEf5N47oHpcswFiH+RO
phHHex7J9PYD4bHVFkNX23CfBSZP0NmlPvgIVlPuMh2qLe452+z8yS5yNCJTeHE3
QJDSTkTPRy8fZO+49u93uT6HSk13RdSvOGlT9fu9BsZm2UdoWoIsOsyovNitR55q
uR6a62LylGYk2zlMhKAnKxSdIjpB9Dkkb3pZDMN+cKnl6mq06WV5R3dFPO9vDnf5
uDXTCiPiaU/57RPTOnGRfw6cEhAdBfUssg4ReOAqNemvKbIycihEmmZ72IY5tD2G
3+IEwjyqUz5vn9b1lVjcEXeFWQNSsR2thI0gVynylTIayqrwqYuEkCkkozFxd5Y5
AYGHVfr6PKVsROdFiL5RJ/SueId0Ne6S2ygdymY+IpLMQFA4TPjul6lUsOqyNKH0
VOok0+AMkrYFLvZhj9xiIpw+uOKDXH+TludkqOLu282IFPYI1wyo72/4X4XNZ5Y4
REyYIFTyqNh6doC+q2FD/SCwCs5wkkLLP8/dzdK/LK+bvm5UPMo3E7AN2GR92TgQ
vxMUC/CmLmqDEvIYVFJPH11vb5OtkFf5mAhaCkFJoOSZA+Nr2GypvrSZ5Adq/r8b
5+oOtjJYU//UdQiT5RmsF28vCxd91I6GGMd0+icHhTymSWmZAFTS3mSy3A02OzHs
SCo9MNZVMvWa15gUWJEDDd471FlRH/K07VPFfmSAWTDfJx3oeVGzL0A2BWbkYxTL
1Q2YC82uxXbl9SkK9gBL5/xN4CqgKgB/jbuBhPyojb+3CknRDmMBzUICmzIXfUiY
BY76D2xtOfAw5Cn4DUACQAwWOvDNeVesFQ7Nm8aDb58f4Tp52uh0xBVhNxjNaLEg
mX9KIrN16WwzgyiPP0x28nyS2POecceV3Zrsc4p1uoTfyyeE/66wW2GTAvxNsbKK
LfHwudvZr7vU+bGzHX1iG+gcUPXj8x80qwji7BUyQnNXx8ACxKk3nfQPbfMX0bAP
JSYidyqqz0KrLpEWjYgQyIVjOaR1uOfd30OsWg+/3F62hDCGtGR/C3UN+mpBHwro
uBiCWf6Y9BvzhErqjNW11aGiKvzQNENAwG253suvEn3BBbZwjxkpgmdH1pxaCDxC
U2VL3XMzcLrw4CdNKdKWfFthvrwLsv5GQu04VLBmM1xjbXB5SRDFxR2fr89smxao
hRPcQS70N/kM+Z646LgVHDN2ZSohB0mKeumBsV/+ZaijLewikddvIjjA1YpwoOwP
B5gc4VzwNnPZxq3ZVoUP/CLskWjh6hUTVna33xj/UfNirzch1t1XpRq1IUKFIJPO
t4rSlqGKbOtVlDZwfEC32srV8KRjR2NQZMxbyyv4xoDECbDRUrW2U7C1uFfJ7Cja
XPyZyg8XcOcywjgPvI48vEmKms5vVMz6CmGiBmaqqcP90fAY6IZw/0nDjjUiykpp
c8RkDgjD6YVWZT7OQmgzuFtXvdWOS/L3C4WAz3ZPxETkHEsqmYD1+/+qVdCn8AHE
+KdWrOauEuGkewPsi5gEHzdk+HTonm3GY8VIYRlLBdFf8mEo0n2D9YuIZA61yBBy
INzSExK+dXxis5HTNcPKATAprHeLl1Sei3hyFtVt7OB8jAoNC0QMg6E9GBd/RLR5
E/sHyqsL9P+4uodJoeXyY4IiaMyPsLknmNyz5CZocuVYAFm8Dy+B46UfUfEceLh3
AZAc2sO9fPRJ95fGpWMVfwuxSjxS2QphD+OiFOb0iazViaKKyv16Yl/n0Wh8GD/a
samrts5g66lRIkQtDDXbmf0n97YXACqY0JBDqY0qoCQ1/XPt5ZNxYHlQBNvZFR5e
nCyKpioOKyeGdQOEBearbEeMCi2o+jLtw99DntZ+bGD+vKwrBRAH7Mzn/1E3FpWi
dhvpAp+eV1vzqv3mIPtfj8edyxYY9V7Vg6V9GjEOwfLCtort6QMl5+zASFDI/bsq
7zXn4wGs70wfuUBBKjIe7bViWYLONjgPYo8c6JNfFkyjaBy5AvC9TQiufVXUHUdp
NuU68dlsaXQSiI1izqHx3jW4NLDBOky6nLL3XTTLgKKmTw4GcCL1RisLplQ9Vfa9
dD96dQoxg92c/OESYxQumgLX6s+8dN27tWk3l+y25BC5j7jE2LrcNDRBxqrY3Fq4
q8J2ju2LxZ3uRDhH6hOcNix8A/ewNkonJr4dk6rOPyR2dqySLtkztO3TnqcMrrZA
IQPsgbOO3CcZ6fXwd3g3D2Qz93x0csiQfzwbs4GtDRlkz4fDfAwxT3M8PgX2+Ghe
ABt/0bEB4nZEgX9+R1SqDgSX788M7dGXCihNo+sHAjwd+ti9CUxU25gLpxraZcGM
FonR6DtCfuPc+6FKbvuHaMZXQaJ9hGFj5hpABWLm8bKpXNI/BcKk3xJQjb3s6LCB
YZbMYJOQMJJe8d7/uXuTWWN271aEVdovQQSqFXlbDwP0ct06OKuDXXYA7C3WRr9X
p/+PRnuOm2naDEEbUtxbzlevgZVvv5BqHAKxqNC3WHqc4704qO++n8FBac+XOcFd
Q2j66HWhdjd2aZpNpnzx2nMR1lUPUnIGwuYoZFHVd6MFncoyAKPJjH/BS8p28vqL
2uM4kUYyNuGzQfK/DNlz75wdCf1j4QRmm+IEp1eRBk/QxKHjkZfIX2TeEdSjDFfv
jXIz7VrRfRYKHs7RT0CyZn3xubGAG5VbmcAxBmp+Mdf6L904aNi8e/H9Id7Fj2R2
xRWRdnR1QjOo120zosUtjzL+cIqPLgUJCgi05mjH0DR1/EFE+PDk4IGQw4vIkzQe
4P/OxlR15ilJoMAr9bVPP0bxCpRTuVRuW6FCxFeIL/EFwcluTmaKmCUUGN6j45Ql
QAJvGOIxrNn8tHnfmNL7Q9wns8TbL/0cgS9uXDp4tA/k0oZP9clZOAGJKIiCvqDx
PMd5WWE6jMKjiz2EiAIxXTX1KPMN0jSQjSoTJRqzEXN4j4ip013fvykOvf7y+fPL
E/4bVa/+vEKBng/FrV3YfM/mRuTzZtdcE7yAiIWVwJM7hOJ2F3eF9osxKHqJJhb5
XDLOZ9mMfXe0RYDQGjGZrXr4YIadTsNBzhD66uGhj+p0tRiTnci+G8/17lcZzNJK
s+USCSS9X1oZtOjWNSXuajPBfeT7amdwgHiGmJFo21D1HqZSin4/Tm0JgjGK71Bp
zuPH6ldOTRGRD/04hhHF2LuZONlt9WuChRV6YmSx7+0ZBXdztO5aY0VRYwrGUNaP
D3Lj6sfn5eZhFEHXzEMn4EGc59OR43hd14ZjR/CXbM4Jm4ncIQA+ARBjGV9CkrJT
G4E9Q8q5bEQ7St5ys9e04LRtPf6R7KyKdFwYpo11eyZRufM9ufWSiidE7ZKOvoxF
wySuNPxG3uQAiPrCHSSiGl1JIbCRcezLxQLwUqPPWjocKRUQ4urmw2/P3H6/BqyJ
E41ljnQv4LW3febS+SBIs8kyoDVdZPJCT8oXW8rqa9c3W+qZPKv+GnLZU4uyXiHZ
ihQUdwJ3AehKjNm5GpenJdge9/SJRJS1MJWXfJR7RZsrdv6dUFlNw1S3bd+6pUll
NAeS+RCIGhzzF4Yy9yVQVhlhbyzzT9/39DTCLcuzUmNf900/UTavohTB0vZ4NdLT
XnM5vwB2NEnmEU+GM7ArpOT6YsiyN4LiPHdeMrioiTEm/fyeJXIMbUoAIA1pTlD2
yJyexMbu9kPpzyQccqV2Kb7/AOM+4QYFlq6fENqIYQO75MLfRV12zOiIh8P/9mL+
RcXlCJb3LtKymVOz8WDX+/Wl+axVp/snCuQdqzbmXi/VH57lY/2YMP3Oz6GNvrSX
wlo4+1Lbt9nDCmEa7sMcy3OFV8MB7paANvZonu/vq9cE6y5GgH40QAEhYR0swcpi
2+hz8cXsrc0fe8scgEKU9xQ6gzqZ/SyiNXCbLAVa9qBbcGu9z7TEvXYXf2LK+oVD
tLtWfe4qxIqHqagdWrAQwZ4ZLCoargCIuT2tNPQ0oOoog/bmnWyEEjzhj+ni4ggR
cOtNbJD+K2hXP44uFWpNxN6ETe7QOtodADX1AezPDWfx3snz3hS3X9W7CWiYMwi1
+ffScRYwcn+8ox5aqkkPEHBONXednfRK/z4QJzsJPZpkvKk0DmPHuM6+L4OsyB5W
W9f9qUsxJD2RtfiPefXntC6xAv47NHl7hWol8cF01O54mC40kv3n4CElyZEYPgDB
4ccFZxSZW1ww3u+U7mbUR47LFfMA9dRtBcBJqtUdf1t1ReRBuZyRcvX51Ea+Yg5a
ED41xU+Hl2r8B+Uojq4OSkKg2/AHuC8Wi6RdGHZ7WzdPtgklLI5uQ6acBAOkgzuU
5o0OPunB7feqSm9BEiU1wHapML+Z5EFGvlnCgsxmSJANKIv3mlY4TPv3Qp2GpQ3h
nUirJPZw3jkadSESjUQbdIQKXOu+/sjP3OcuhJfitP7QUjf+AdrMjr0bI9LdtflK
+8eg6e23I70Uli74iQKINrT+z9ga2jNeSoqNpZV/HFBdtjPRxRyfHv3+Eul56b7V
Tpz09zq9DHC5mcI4pPW89WdpucHc7oxXFEjbZH8nu2M5XkdfulKhyZEwiOTPlNOj
mW73Hce2ws3cju1OLvGNKLbFqeVaKbczhz5+ePFM6VPlq1pkECzPRfGmCbMhT4uW
h5YmdOxvVirS1yTDMdkKtK6mDcxDGFMsxU+oQ615t5eGv7tS8a4UHXOWHUefyiNT
df2nkRqcQ4xeU08xCdT90Wt+H9jW0CRqmcaWtQLPFWmya/Hpb0VrX9aZCqAqEpSZ
lG4efG+JbnEob6ESHaVZWFkAel7jMXvhA8z1z5V3jJafeIhsnUSBVHkg5BsK5zZH
yN/7r3n52svyk0P9IfeJSUzYGVyurIelAqqyITmOo5POPeW3qYjO6wv5n/wzaNLA
4/Y+VmVtrP7uhD/PYkCWx6HM59tRQm6nssHA0mBKyTIEfz+4d5GgvPsgFwAqQNHs
Ay666qv+sB1xFH00mkfZvCjfid6M5652R20BjxesNKMuTQ+zDoardsjd2a8LFy7Y
F40iMMMsrM2VIQYNZmrefrGp2UueEOBGDwmVLXIKFuRI4sD7+PNVtdB6R9Afv6kr
9y0oO+kySJW+u4K3e9jAkSdjFeKK7KcBI7m/QnBOyspEZ7Z1XVcd0rAZrdaACGq0
o05iXnSBEr6dHV9Dm5gbzWexLGhj2yDeaQTqdzDGa9xu0mwQ+6oI6Gq2C6qXpDgD
0DP2VcQGE4rFDWhToQXSJk4Q7f7BV5NOdeeB6HuqiFGADQ0ytESwSb47sUspHTsO
n0Esw/EDfgsAYgty7Ghv6HRfK3BqhQ2m9by53H9/zBATYqBJZ508RKscmYlrBetI
cAXcWB8tWLFszukiOvmiu6K9yK5SP/pqkEaB/WAZQ0+tEAbXx7NIlKPStiL/St1Z
7Wi8XrB6TkEcY0UgAmzXqR3PJTGPgA1uEJ76C19b4M/uCtqIT76dyxmOr0kUTP+f
33tiQBwBS+M3kbPDzqOdauyA791XnD0LAZg1EZPUejE3N+Yt6i+0613rYNRVRaAk
9TxQ4Pj4NeByMDbz0dIr542G8OhRLAz4CJFXlSuvIavw6RmrJZ/B8Ufo0FHBqn8z
S+J07r7LOms2T4/BTlxfEd+9wsO6JlnFV713sDidgWiid70afMrty9Ynf+0foYse
YIsUE7NoTzhqLjrtAa+d6LTKK3R22dbGBHzNAyG5YnpCMU0+c87djAQTMNi1FDGc
+YNOCJ3Hgc9Beq3v2UrvkbM4YPj5UdnkPCPR9k87A31RQq+efoX3YmX6/06Ft2MK
IUL8/Sx2TTUhTiWFKHYT13jBetRgGudxQS42S4tgaVc2vUXnqh8TO5KwBHhhKzyY
6Aj4B2yu8EkJqb0/S842nhKmEBl/c6rgbClROUwgEvfZXV0qVRlIwOrYKJeYvzfK
f5AmVQtGwAwbrX8NsdtfYZeROU+rM/CtdLuGqv5ReboH7ZLUfAz4eeGHPRdkjpAC
hW2czAhbF8Ojfw6sy4FeY59gz8L93KoqjAWR2HaTntZf3Rqflal0ACVlnd/i5YN5
uJ3V9v/Xzlfbf3QZmEb8WK5wBwuSBkO0JnHo+MWUW3htEhmHucT47IUtCGG6qwOa
HcQ2C/Fks6cSq+3BfG7TB1dtf9QVLz8U1uwWqfCSTmwfaeVlHL1d5YL/gV1XmZFN
3NnCVmfvyDIT/zCCNruYKpxfnnicMP4AmJ4NvlYOIQPklEv7RBCeVNNG0iWovYuf
SWgGVc88ToRJDOyrSCcZbZH2OvVl6w3UoE+JgEsc00Kw8gU5wrfAZST0hVPpB+Be
wbuKl/f4r06ToAVjmeGlIvlxTKdlxXmgfJz1sheOh2hW7Ma3zwu098WUIYVmFQDO
fM3GmLasKePFy/fWH4lNqpxJcLzJu7d1HNptQDmu+l0D5uVCKJY8oF497vCAcMLn
gEyuDK73mTAMgQZF0negUsLMYdjjFILqQ4Tt62XMGDtiiVu2XFwv4FJBKdwPwYP6
/UCWO79YXcBULDGODYp5dju5nG/mcF31DDq/8XSGgM/4S9grc/ew4SqWVQsfANk5
6wH3mQvWrfWPKU2cZ3+4x1NxJ66OdM/XsdbcSZrr49BbyvAbgWdvWmO+w/RNev12
xMMqsz6tPDT1UIn65FLA33tc5uNGgI9QRFKgtMc9n3mgyw4tnle3ALpgXZehtlL2
Nb/jerozmveVyiDxcCnvqt1vGQbVrSdcSE921Ys0b79KCvyCA8rHag7mjdYM8Q/e
kUvHPgQNtpmNEShAYKK/D9TKmFeEPOnmSrIxfk2yJwLwdlwMQpCQqxQct8gm84C9
2/5rvVr4uSsXP80kETZQLa9pA1H4c3ZW9AvxHfiJgkzRaaAFdqdHvECDfm3NxAR9
EXug4gV7ZQbP1lFSlvzLKvXL1gb05Z876+WbW6bdOaQT/+jrL842hS7VasGtq5WW
5k8t7aeVVux4N1oo9HQzQ4oGUp4+2rIf9j7otzsVdJdzaT2Vm3Kmw85Y9HQPjcW9
gvOs1TF7aS0BtuhRuPteuKtgBTXBFp5ncKtZKfd57iwjzfB8yZduksrUMtaEtuPz
POCgOK5SX2E1pfXr/M/IVE9z0508nUtYZL+m+dW03hJPtA3l2J4oozfw0H4Tl6is
pwBFVS4U12Z0pVnZhTy9SiSMGmhVztghXa+j6a5MEEY0mLdIl2kwzXApvpNuixw/
6eJfJa56RhLTyMeNBVrPeA19261nc5vkpPI2p05GCwB519jnj0PLZ1NEUxX/4kZR
s7VnZkduG1s0VVsRUL0NeI/ZuOiebQ9P9ssoH4egBpujzpcGUp9LFdoZSETyBS8U
y+MLsT6RlpiQRPjOpnWuUD+tawpwZc78I8aN5WmjAtbxWZgF49UULkZndgqzloff
wd5vrpLsiGdmCw5Jr60mfjk5+3LCyf0vJQqXPBJ1lonOIiGS1nq0dbAQJ+qD9oGb
kF7u4y+nhS9mNiXLfyJzSFPMHbUoFcPQgcRvW90+3oA+GDlIFZlkKI461mHKG+sf
xml4b18jl+X2efurJlnmx8321efg3eKuP0cDTzh+ssXtaf2hUsbvboDDD3Fk34JO
nu1dhTJruCVnQn19+zavLQxbubKPQ2A8TV7wVl3CoK/kLNhG+KJeYL/tsnAma7dV
hbBMknAPAdYCEzX6Jbj5/Fo1FJvWPwbbFag2OAHZyDfI8mjPHYtLivOWp95AIW2R
iDS/n+NnKzWY9+5ac34cPXaC9SApC+szFrWo/hSHHomP1rKBoHsotuit+Ywr1EIj
5YGiomdNg9JtVf4ofggpu+TC//gtHpRbSZ806fGMmlsOYrxNhajbE3xYsPMuwrFY
IF2TNEYBkpZfB18y8EYG65bqJsY+hSIJk1nF6T3QbbS8Mm5I5VIXhV5Amn9C1Dkg
yR7UqjWyjStEH85/GslmpL03rGwkwWdxhNC2D2prqM0OEtyyVlXdGuWtCDuixgzH
27fqLb94mJNvIn3nWCxD9gu3tkX0uhRUZrSI78A804N/xsGBn2DnUcGLX/qa5Yc7
6EReUWm7r5P37jjHbvG7U9Zwzt8pNRYLXovWey8x8+EO7QajhgS2WvWB775l9tiY
URWz9VdDFE1X6UID9aGqagLQgqZLXzpQeqIO5AopZhh+BmEyNzS+bLEqxlY7Kfw2
eqZLXncyRlHmEozDiVQP6MpUCKMnzK2m8AFXJtEFriPd+d71ERd0esEQiGgTUKYJ
DCFmrHKrvAljQUlnHF2sIhhlx2mIL6FwvaJCamxOClWeYGILKIsvKAr0zesK80pQ
G13hIsEKU+53rEvs9V+s7cd5kte0BDYw4YVr9qPn6LEyx+dD8gUpIN3cnpNxVbH4
llqmsjCi7lHhv2T8yHgR+7QwZROj3RvWLWWEH4AMCO48vrMk72cNOHsXUyrNGcE4
d8xanzGdNsmDqgr9AqGqtb+sidNd01/IEO+6MLt9CM6mLzObYFILSMS+kh5E3BuG
vGmK/pp+L1ItZdAXIyOl8eK8AdOCzmyAcBGNVxH6JzBrpujY4nHrpjt6HvFdK++d
tLV5/ZjxiAP+gNUHWrl2ZpshUH8Zc9YPsLSW127dsFUCneT1nfyV+qehLg9VaWgU
M+sWmnBmnCptjy4c5p0zcPUVwnXm8K5EyB0Q9/pUzhdkgu+tqhrP77z9eT60GTKn
X3VgUGFnfFjZCjIyO2rX8Z3yBp+fixYus13wXpCezDCOA4I/L1d4kRFvknmuWfvX
g+NNVt47p98kxzRFezEbtlb9FqTEaT/0ucytN6EWX+aSzFHsxf5WYQllNv+9a1LT
FKshrbhUBK7waRMji8xaQgfqYtsXZ+DpTip/2VeI4yRxf4q+1WIsCga/LZzrpovO
unz+NdrMk2yr8omftOmVGmfWdVwzdcG4VVTWqkeZ7JwcPeL+zKD6ytVfNceSDWVD
nDKw6swaXR09OPfq9kFmfCnRz7fqv8w/MPF6YYZd1Wwab6qWkl3F2++SI87CK2sz
wFm1I3lwTDL8yBs6mCeopEyu58sJvV1LlEBLBeKzl69RJXB9N81v5BBSMk8GY/mu
SCUZfP1cNmTGXJCmNL96z24kq2SCZEaJnL0U+ki0KS5f/sEHbvmgevqjsv8LknYZ
rcdfytwcc64AE7gpxLM4hvaz9kp+uqVDyzkt3Mbciwq3SMpOi3y07TWWtf1Bjryc
+54gKAqPurnetiLBQRHjqUjfdAxK1VqldJELvLOoXVEAv2YzAi3DZPhP+nsp+CzO
doGgvsGQDhPm2OChYc/3OQGFL4XLOm0fLKomJbDqLyDsMFh+emhEtGxP14h5qNBe
IwP2E+//4ky9ho0iTVVkuCca06jRuVtDtUUYq1h7g3AhWBmSt+Kq2kNnKjIs5AxY
nJ1pkE1DbV2oxMTHS4Rpj77rVSbQY4aKNcv++KzP7XKz/gsZancHPWJwXf9HiYDd
km8C9DLy2UfKn93iXkkmoW1ICD1M+cM+hcVh6ZOf6li1ZAkioZp9pDH1FY2XgJVA
d1Y5Kt6xvP0qgeQAyDhGouNOWlWhIoYK51Ub6SRQ+dL4lodj5mY/c2ddY/0KiAcN
iXDVhV9BiiqioNYIYAfCwQm6jmvUE0sLy/Ia/H3/J1Sk6DkJhwvIs8/pXzQdRKxX
EtyTRI652tgzeMdlXiVgr5u4XzCDzhpibpDidO7HJHtFdi/gVOdrGNc7fB8HjIHz
T6nbdNbvfS/dmqIOut0kghHBPrc+eIVEGFX/XySuzXRjfXjUGjDWW/OI2wEIzRjf
mQ6gf5meW3GXpy49UQkZTfA+fWTxbOyC6DTsXO+HN5y8zZAN6/K6KZ1quBeN/PDS
nnLck+rSk8JiELscazEl2Ytco2YU+J7P2ACpWZ1QFSPHY5M0m4lAXO1qcBQgdTQ0
T7tDn8qtn+D7l11PR9CtvQukVX8PUXBYYUut5nqzArpZ7oj4vRv0ZpPJrY2VOWhV
SdUAZUkyPbXYo31aTaqTcJrRKn+EnS61+Q0j408I8E2TxD6iCHQSW9EuTk1G2tIS
v/RmnWEM8diNHO3CvwZCfmr/LMYRvU/aXMGZjSX7yFsvCcSWJT7B9hQYqkNM6zaa
dgNmmIWLDFe43MdNnf5D2R2+cRfLELaTnOw1Vdl3hz1BmcTqoqpYWFeRg7ayNKNz
Log3wT+kCM/z4WRhBuhCeKUGOg8LMMKJiKdvgjtzF9ofhETq5oPRnlGSsLBIFAQ+
Q4dTe2SWTt50HvErOTUp6vNz6N0Wz7DJrk9tQT0QsFi86yNyOKFx/ZLHWWaZUj4A
a//qGYwFknsXaBkav5HHvHM0eEaXSkVYEtzJ0Vo7Ui4k5Hgc+wqpncXH4xYc7ntp
vtSWHji/jn/QS970bRogt5FkbVP+kwtRel0hXSjy25/3Ht1Mf8nepMSiqrA9ayBS
4eg2+xq9ASaKyI5qUKYlByK7MufJAbKf3JuA/exieztr2QODxYNB9/JDP58SPuvt
saQUjUPoKdJdajA7VSOam5wUZWYYZfWlZPqNpQ0ZX2GtZUGlLDuH2lhpe8kNYkSD
ZxsLY+xF931tlhHWM2gRutrQg+CbF171/mWPoRcu0L0f87aJ9ddXguU6gqBMN/ef
OHAEKZwuLWi048jMXUpr7mB+tJbW1CxFJ+jDr4vwVv537YWQyjktP12O9bH8uo+2
mhNiY2xa/EFroPnjKDtuA6Ttu00poIm1VFryOUXTLu/MOD5Ps/jwdyGCEc1T2auV
/zoNCU83xz/WUwF3ZsMLaCsX1BHeD6KCivycMQon40rudgmEa/2RnCzq1ciNjqur
GO3jkzZM0s95Y52gHyf3Sbh7OqIsY9s1fQUy476+STmE2j8pBwGhB2KjkQbbHZkn
YD/h+Krg990+oeZviQnd7Rby1Jr1YOU7ciUY72q1mBD54KTp3kJR8PB+PwxC+GCR
uXfTS+5az+lW6Bx7OttHDf2ygwfEFB+f3u2RLnfNl4JEBKpxLw6SBsV8EId8CUjm
RwDJlObBBtCd0NVnoVahje6qzrkBDdmjeRD+6X75fux4lABjJ6FVVw/5Jxb/urgY
rgqZy2/EBBk+70G/I5Je+OXXCI6TGgve4FZRXpXh3Gu9ZII6VBjlh2SbhaIGmFLg
mMkIvUHRpNlHW5/D1YSu12sLdx8hzbhQk1NVzjTiC95zT0oCqGNNZfBIYBvV/GqX
P52qN7t18p8BHRDLtuOUEjA0cS/g4lfAvy9O39EvEH4HSb5YSaEclHmYiYGEoegD
bPuYUoPfCdF+HgLC+2M8X8HuY34KzYLWIQaw3IkANQLRfH8YUGYqbj2dR0QSBE1y
0fYq+OP9qwfCmH7aWWBuzU+yHIHMuaon+A2pBWyRGNz6T0eAAo2u/nNMCKLi6MCu
ZuprYf6K4ziuMxUxWo0/5rWfeika0SEIKSA+LO8GhwKoaLdorLoUE4Ogwai+M1MU
sc3iegXtu5BYPAjFjpfdyn5WT+WajY4raPkB5y64/1a6xGVo83//eG59vCOAkJta
5v6UHL5uTeZEQMIVordqZ9zT4c86RF6H/kwaWJLit4VdxIEFy5YYSGxo5fcu6Rv9
EKmaIG+d7wSwHn1SW3ylrdghWYVVDJS3w22fUPvoXqOZl1l3iVYOeXwVD8pj8mkD
ibNzsHPBIuE+gLHs6xvn1MgWgXD5hXbnmbyAFQ2Sg3AB5HDYtouzXXJfKUeB7Hi6
iF0slhYgAJzq2m4/WkWplMkhO+K8j6mze28/xW4Aoz9Hixjj1q6dxT5pKVtWX+lc
YFI+MPQJFlyEPDAdXKHeTUG+QEn2I1Xo4CpB4uM5nFWNFOe3eQmPWHrVv5WIBOa2
LFd8j9tTIvPBm8Lxr4sC3Yrtpp4pOruZS/Yv2zPBv6PAHpC/ZCrGcLWbbG6Ai5G/
bRZa9aiSFxz+5YP9cxRIrw/A+y6QTbTGfUXx5C6hG0zmebs/ueIlQVewTIwK3/q+
/rkgtiN3ffPlj1HNM23AiZbLU+OXgXQgJKssZ3MNEUhprJuoJhID6lPE5RzCiiDa
TqDcWN6qlAm/BJAo3/3z+yxZOhhFyFX2fgjXdDpUrfBX890KB/XFbi9lA4/hhkLu
U2ihd4QjYIoYhwuumo/7xkWfDg3kpKrJoJhuOauEulSD2rc0R0KPflDEPjtEbEVG
KJYMIAWKteeRLkwyo6Rk9jQURukSF4LDIqKg2bxVIbSGb9r0SHyFBexlNWszoDG3
Yv1mIus1qlLMdDCthejn4OuMI/Z+wD4q0ZWF+SkzcwMZgo1YWDLXaKZ3yIZ2TJVI
0F8xmcURGomUiULeFftn83Alxu8PdG0K7O4Zz5PgUBSWpv5ZHNPkMcszY/DDn25y
soARJqnnFUzQN4wHntAvNXLXRs/M7eBhlvY9y9yDdFtp6NwW0PZOcZxUviXjwfPt
shnuZNYhVZAXFoanxOHJqjDDztlhdb12up0F57agjGyvyNbjEtYmeBfjHAMdG0AV
DKtetc/6ZbqQ2VG49EEC3gODCYgiEvy1jrP8OjdflJsLDwvMWgzBSjtqIXOy4tNP
IAgY7tz+gWo1fTW5RmAnLDk4nLgWhoHvwyBXLsvTJJ3HToHjlQFdVOd30QJ8XTH/
h69AjVOh4WAzleAJY1IAr/WFv14s8bkrRucvRwXff7nUrlOHfui2iV1Iu/lC4N3h
Ecy2OByk81N+bWCrUhdQRxQR63lRbwneqT2zFAAUQO4AiGvTQxK7eX+tTozT9uJJ
5uEMBlAIsT6W1cpdTjqWiXqxB5AAZ6LJJSYsjpGJKEADNbHiYPuUKrq1h0LUSi5l
fsysKi1+jwjJ84dxgADMIil21ZJLESHeTlcHUyj5jeCzxKH5QSJilArLyC0S4cXD
o4u7dYO0YZ8NfLgYOCbZ/vtnJnuse9qFKgbAexAuA7Bj76roVsHDwrkgPSOov0XG
8XyLxnpenaTGSGeyZJqSHpMfFGm6YomEo5ykdnGO4qWg3znfl9tIVlDy2RTU3Cro
XwteCyWAk41LbyCcf3ijD6ZeVZZnzfnLgPm5CPEAlbZLD+jXZ80DxGRMbzi6vVn8
vZMRFx4zQUDjyOiqgWjK+zvmv4udp1z3W+JxDbpKdL2o5SAh3iV6pTLrpK2zgkri
2Nio4T3fyTINeKnijzEAKWxB+bUIvvwf5pDikwE6gySPn60jyIgRb/oPTytcGddh
k2Z0E94fCsuAoVllDu5fML/UOnHXA6eYCvTv26t5Jcaefe/KkEEaZi0DpPsoXaOa
ShZ6mrU5+l5NjTwQ3V2r54iY84SRy3hJsQCHaVtNlxrum9QvmklOIitnoA1uwioa
MLoXhjnI08niEqbx52vwX3ckQQs2Cf/HJ03hmdNAN4R/MvqpAwixlmMbEOeXY7UX
ciSd4C4kcMCL++499kGL1bQ6WOlefw744aFwItyhh+Ix8nDPrGqGpI3hegAHL4QC
0QAcB/JqPwEzTTgAA4obJE8R9uY2rS5HP4vr8WILD0yvUM/twI80GsATKasLRPnv
m0PvDOQ/0310/vovzaVxyKX/h8QUnNhUdYYMDu+RN4cd8zizqXHDSzxwX5PE87+C
5yYq7Vri44+TXmdFhZJ13enHl+LEXVYcCcmCRgvuIVHycGhH4FgEZToIOuk7sijC
jVh3tXPvPbJlCcl6+nFvuBpZd/VxS+e9T2Q2T9Jb0sbFQR3XySqk6UGf4U8nnveM
45lHNTMF+tdVzzYR0zSqH/KCMwTjmSjxo+QBi0sr6O9+BlAE1u4ZjeEUpCH+jBa6
59BpikVaJ/gMHOm5u0sv7y+jNAS4un6ORKS/r8so6FpoRDmtvWOXoQOBv3dK1pOf
GcQNxRJzLaRIq1XNsBqHO/yMGFZah0RFuctwZddbV3cHxHlAESboBTJue1YIfitk
vItYN2nqxoFrHHU1zTnF+MhDtvhemjHtYhGOMKtToatMQfEi0MuIvCIYwes45+a6
YhjfQTaztOsqufX6SbOUkM2L+t0FPnIGbtcxlq/9vH7YPqKW3MIVFgtzT58RTOGF
4bdzt2sROrYVc7Qtay2C21AUyMRTC0H0lGhxcSBXCkGb/t2SAPsqMi9ecpW9dtJ4
D8IUOx1FjT8b4LHaZf1xFBFE3jEbFXw+WrbxM/nZ1uxie6OUi18vAucLGhQY2UvR
of+3rmSIZ9ktegjyY7sVkxwfxMfh1vC2gBGYbkWHYMriR05LwTp6+lJZTtQiCh3S
8sl0pBhF62Gbq7s4mFXr40LyAuBlzvYXa804+OhQ3Y/Bp0lL/8rd5W0wqXalIgf3
X0Qa0cAFSeYTrEC4wqOzvC1+l5podPkJEKXJ/NR5V2WNhXV8iErexYQTylhKxp+K
ErrhS6hbgzrqgjTIzECWTRhaJuG3ijPKhC0Am3tLnBzZakhVUM3Ns5l02NDWdVME
7IKlPXD+QAvwfno+ysjQUTzb0uA8h9G0pR+UtUZjl2RPvHQ4yh2XZSSlLVSyq4xB
AtS1KhMS7Z2EmKXpzM6iFfGO2zmdTDJCcdjYStjs695baSYnRw1+RJpY7rZz8oTC
3UqtSNGncxSKr3clJyk/jCfBTSWSOhs3/YOBvepRcUVLjaK2/SZbt/BAdvtPSsh8
AYOtFx+wHcdkXG2Zuf5ihWLspIdQbTy9Qg6zeS2yISuf8g9w0ueXNG2X1nLU6Djm
LDnInTrCLAxY6oxz5VGi6ycGCKKYnlZ/7cM0SX4pB2/X/ARJArIe6Scl7iZRUqus
6lXTU/Zw1XYoVlds1c5j9NAs9dDn0bIjXqZb3GBmaqQ5vDrf9dk8YEKHVfycLqn9
VNAS6CwV87NKVvHyJFeLORxNN/CxU+yCIVZzyvanTMN4oXruGMJngPEdU6zyA0XL
+r481zBUd1mAlgA27NfBP4XEP+Y9bL+EuGkcQNmWYkArf9oEuGl5Ef4H3ikKhy+o
YA1DXHXBLbygdxwx2zykCKcnWkQYFPn+iZSvAoorWFvi00Ipk+0ixE4yaWoW30Kl
aQ7AXUbvyUp6h1qHnmHIzykqzc8Ei5KVG9KquP5Mi1PWT9aOawtghKibq3YCvV8Q
cgVkR+4n74a2/nGgNjz2RQa0t48Gg5id5XCqPpcCiQZ4UQWQ3MLeyPMtJrF9sr9t
ewPNaJojXl5K2HZsmHSdG21CozaQN9AvykxYw37zuefkQDvDPLoDddysHGf+UgeS
Gvg7CFTwfOoueB8Lx9v7EB7ZgY5RBRo0HJTgR0XeXIavbgWVdQBX0J+sTuECkK40
JA91bEX1syitIa9rd2O+9uq+2OLpOrc0c2iskfLAFbsPvbA8CccDAkqzWFWkx8nW
Gd8F7pz82TGptLx4exTVUAVd18qDPwUuCn2Z3twe5HlRwiqresxY/fHSJIGQJNuo
n+VznT2mzVcaxDgTqJ0Ov/7ddVIyonO7j9+dnc592iBcXSzri4cuMNEvBaHAr0JC
nh8l5xz6dAP60NT9APd/uoDcl2DtsLNwT9ayUHhos8DkdlMZDR4wSD5Nb+psaY0T
seZ9PupgcBzXQkDeMZA62W5J+S6BxcjBWAdTWRq/ST/0cB16wGMZYTjN35Mm6B9h
QdC6jBqLOb+84QIFFo6UpE7YGMk32yKOvYA0vzBLhgShnuqkqdG5YM21GwEsvG/G
dvu+gRmAnkBMH9a4R0TpJPM72MFeS4GnoSjes9/HGq8EmaFwfaK3JPlMRaR96ZBZ
h72oVEa0YePp89ISMFZPnSwrFsS3xyHGQdiwvp8ZnCGqi9/YcZm9wWHpv5TqxJRj
k8wfEDr24Xzv/jvHg2VbW1SB6VuXXwdegTuz933A2KhV37Ejba9qUkR9Tvee6D56
XOEn3g9uxvqUJaBb/DT8kCp7xLlTTheFdW4iDuGwlFM/U3RrJiDyFDhVhb0gVfzl
W9M6xEg81slIMUU1qxJeAdRd+dtxv01pG/AaqTF1/zstrILyWav3FgHtcxtHPXtW
7OzvfdW0tkhv7Hfc/Yn4mA0qNrxYbj+8c7m1AT12LPLMCBm/BBgIlDDVg+Bspb6S
f7I93roq5DAsK3ZrjxRpp+fQNd0iRXB3AQ16t/9V/i0AH6bK6m6qq+9CU/2TCitX
IpHiY5T11ffwa2Zsx15b5bo4QYv/dHPZp2rdI/IKtqzTZ2FV9PCUvh54l9CrTxkA
empkZ6sZrv007JbG7+42CKl43mOeuKqrtD4jUqxFTSwaouZuJ8a8AJvzl4S//XHi
QtXPP7b4Wo7XhpO1zDJO9vYL0jc/Ge9we5tANMAGYjYsyIkpP/Z0FkPqPKwUvVmj
e19TPtaYVUCdQIeXfkVEVxIXd9mORJ+UfjbzvsoIJG07K3BsD89+R8s0EeHPsLe2
nZCPtLeKcTnn3Yok9zqrOsBM8DB2r6QwZkE8Yn5QPnc+pqwaDHcd8UsPuOaaJ7aR
gO40U2K52tCAKsyMoJAyp9KSGwArNiFbxmY1JY7syNSPgnBxFDccOO3eAjjj6hDR
64xRqTozU4aZldVOX3mBas3p9zqVTnAgRIPuWpQZFmL2myA1GGcUvagxXl9E8RRu
eUgo4DAfUUsUOX1kCuaTV3wLjcKGbwaV9LYM4UXzYnsvtf+3bL0dB8xRNi5mJBI/
CUQ2+LjmCZ3Yhk9Jl/pINs26TOpFp1s6hgW9uSivwtZr6O4A0oe+bRRI0+aG8W+c
kExFqgb8IPsQeP7rZIPntCMMpAHC/e8PGSQro8hkUkw0e+QxFvf9f9sujNA1kRu6
4HG/69Imh39uLHANBDvj0pK/XbPNYSN3f/htiSZvxodFOpcBDrZH1TDOnaDEjfhG
OJEAAmfGfwbuUnMZn05WOr+n5zHf3zIZYaTkjjLedVzfWON5lUSGG7tcrz7q0VT4
k3hU02kdQ/8/G39DdPmejdQTJBAQvyhLLBsEBNuD21yWHTMETEw6e/eSdiTjJ3Dd
FPFj/Bzu9pwtXbseCkErQZ1gNk8Y1xqLghUiQsAADABvTgtmtUpzc0r2ivSr2Jcg
x27A6ojk31vP9IVa+HJavE2ykvB+LaQDRDfHr60a59lYthe8861q4AVMZRMd/v9C
StHKYYz73fyoH/fR8QPBbUnklYxj8IJKNQif3wwc2/BHeS6VuTqS5H6n3+51hbti
YgcR4uxTPv5JQn5ha7PNK7Qbu6Ba9zOWoTuYrv1T7Op4DwwsOFRnofrR1XGgr4XZ
xx+EthRQMcR6Yj0mXcCuuvOLSaSk8wZEqUPvunjbIaiMZ29BEscPdSOiyLpRZJ9W
4NawXffAj9kN5C5BXslhDuy1D1YymmcrJTsUTUpJqRS9A8VyuLKDW27Gj5jd/8u4
p6ui80WGroct5h/GhRHKJpU0whtwp0cxnFb0164GvWw83a3dBMSBwR2vwCIqAHwI
kotNM2Yon1QaeIFyXPKD0lUQi5GzjYLYl0QRXPRKJFGfWSgU7LbE+vORtD2T3gM2
XxjB/rcNp9Kp2ZTEGMZqj7EXUA7jtWSuYfuLClLt+I5RVnG+JM7uWfHuOLGbgCLT
qvrwg4xdWykmQ1Rnok5TgfKHDBfVNjvxlrpGwUew4nJGJkzW/vCf6/E2RLLShClO
+vrFMX8dLVCcaYf2OEQ2bdjsw7Rru6/HBntWnvVfbHbVyn4+TQ1QexE9vzbH6oqG
cDKa5Dbjfa16FbW3Plo+9femxSlPqeNuqjrxS//ufKvMj/4dFjJO//vXi1kjVzoP
q/gJsyIDGU/i7mtpK5Jiu0pm5tcx7f5oxbMWzJJcq861Wr09m47NFMl1BIu6x9wU
SQyM0x8sSCQH8xw9yro8qlhhQrv+RaY64ENJI4PbBcww22nw1mmKHnZvmufyQa3G
SL4lz6LkxG4c3rhU+7m4f7MJmI7sDdabBPHdi20FdqYe2iYPQTHznVesDrROLckc
bbnL+5slCxuiD+CRajz20YjqbEncPhxm0F+sc0nrzEhnm57cpM9m0ZBhdHPaPVp3
EFf8yBnj6lV95uLX1PX9s0EKfvv2mdOl7ncYTdgjCnAcM9/tVrbU7JLtV9iE79fK
M5j2Kd4Djx8dngdefRs7wjyjiOX+Ux8HTD830yoVKhojwqU17nOuAjl4oIIxhRhK
E2Uk6lrSOOFYk6cXWtHNMDxQYCMkVQcnrQNwyZRxNCESco75VdEgb9U7WfqnepKG
UYB+iXx8ptWHEjeREQQ1HT80jciuyNTfaDFDRyYmnjhsv52CzjkqlRmza+dzacYd
t0snYgE7pe0qg+TxBQPoEauMYqo5DghXtNv3giKoSbAPiOiLLU/SfxFQZYCXqxsW
pyU/egizfdZnxMFUJIxmDAh7npCqr7sgTb4QzeJZnuEzFjgkRDIxAiBTMSyZz9oB
Sh7kBu5KfKqbb0w58KMcWuzs3b4n/sz3kXYTH6OyGb5aXm1XVSyHp8+IyfpLp3cA
wwzKYVlxzenMqs0uiqmJmAC9WRlECF+1sDnn8Qsd+2KZaPS8hwDwsqH0R13gsVxX
XphHogGj+XFI4OIvIovo2iCFIDYTla+B+3CFc09egHQty+RZOlI+spdIxXDABl4F
MXMaSQyNtKbbDcuh94aXIMEOYtnZQbcoHvqicozb83f6NwHYMKuvW48gAgz23qYF
gO/SUqy9BI9ruJKiRBnCCQDHZ+y9CRO+cPUuIduIK6lIGzRZLGmA9HH2+rgDQvNy
WFyB/YT1Hc/EWVf+0ni2z7e5RpIGGZekm2sjdH5uU6G3D2m/sa5JZ0BG39/s7cco
p3juupvztJv3tqu9kl/tHmweBcQ1rlO9dLYxAF/oa9GveGOv+HEk1ZeN/wFr/mRi
aIX2D6AmBJ28Zi+tMtnRjYsicR+5ZHIDOIM2dAPda2Omnp0LEItPEmIuo8EwgvIN
0vt0MtjoCAwQdsQ7amK652uSjb1ZdtoR42beomHZ5Yb8jy4RcuzRZxRgG1HYmHuF
ZNovET9BNgQAIdOJS8qE8rUSC7XHs7Tlmz8lTYW/w6m6G471spkP2ejr93HxWlpR
P4PxmrdxDbqrMgnKo1Pe66rXj38ylncVpdND+D3zvZm9lqI1mFikwRn6tl2g7DtM
q5IfTkSv+wkJVHe2Khqrc6xEi12Pr6mISQ3RvZDzgHbWWxgzsNLuUBpAA+4uwxiP
Cb3ey9F5Tyu1IZH2YWi4AGZfRptkYWpyHT2fmKEGHI6DmDrVxfGe2Zc0AnIfBZhO
HgtIVnDRVaL+I3LQUj9JoMv4IBC9fdNqNY4XxxqpYI5JiCIx87zA5tASJlz+/j1+
XLV/qQP8oSMX2tp9SbmAFz8v43tRiGzSYp2cKjQ9qwgX+bRpizmR7E6hGKP1KqOO
hGbWlUwFGTdp8TqYhuUGaSZflEjF3BeAcOeARF/xw83qWlPxFAOUfNHGsAIEHK1p
rN7bBzrh3g+BPYKiaT/C1g1+UNwY6s/sYx0Q9GbM0SyFR8xwxHJuc2fhNuyET1Y1
+AdHKkUWc+jMqPJjd95xoKRNukeEOHb+n067+aQIRergR5M8AL11Qb0+ego7/aZK
cH3yV4d8DNpHw+9XSlFhFI5UkopBgB+8oTBBx+U0Y4tfrnLHi8Jiw/BvxS322GqQ
7MMFN0iL7Pl0ZMQichm7yEfkyKnTaCQOKrt8tlfMwz1pNFFozAFyszvCb4NZG5SE
imBPSQNpVxK/u8uCX+JAD6kSzmIZA2P8I3AtdnJFTad7m1wKYCrTcm7NKc/wJ7ke
bO4ME4LZL96iUiltj+UTRpBxkBoI3piL8RqMo+2TGPX4ov6hK1aGdoiFH8j7kg3s
Kte+Qfl+0/I144iDEkQteFKrraWgpbQdwIEaJXf7+rCmHB5PNA/UNs95iY8sD3J4
8R13NFhHjcrO8nWQJpRo1uaGebGtr1V8tMe2Lqn449yhM0JMjiEALqbjtoUFO9Ui
FZC3mJrgTtlp/gtZdPx3Zz2+292YhUkMyDzbR/sf7J/KMa2zbrTWbqODe+DLlu7p
sATC4PX+OmTBlqNi54JBKnlAlsBOsq2STBACcvqJbiackuHHwEnstOsbnVT9nC7F
Hj44RBbtxnWrOH4vJ6D27r+VYqaJEnjLGTrdo7zwi74/I4Wsbl1a4PvEYpkjabfs
lwcK1Ms8NmdoIvSnFkYy4zwcatkC2vzvI/tTrImPJ6jvU3Ba+ikvHE6CT27FitsX
SRB9smNKT0V/XveNQ2A4PbuL9kn+JFU8gbtpql3vrvFLR1pQnvuq+QvDeCnugEkK
f4BvodNHvWCpec5NVxeDAuuMg9v6Cz8rzCOM44hNK6LX+pBxImqM0R+DvOI26DHd
WYNACSYKatGWg8PUOMeVaRzxWQTweK1zuvEgnR+ogxC2nbedbeNuKNkVYgKhatep
iyokpJz5x9QzUXqbTgpl86fjRCrdawVg8q9zZdtR5RVZZiuRAYHjUH2Z2+gbURwC
1RU+zGpFSz9lbBRC1KyLkRcUB2TkIw77z52vTDkPnsSrOMdY3usjqLr6ssVcBYjl
uIz9smPLzCnPfgtSRoQaaxogbHsMzxgLCrP0pT4JTuXktNCg1rxCHpq7zMu54uzD
qM9EJJTBcdNSW7fouR2H2hdrGiN3qoauyPuoh+MXvQjIxGMB+IP7LsUX9qjFHIQd
GepId7mARCd5A85K1su6Eo4Qx0ko6WkVR6iSAkq6lS3nl/vGnupvYUowXJ6LfCqd
08QakoarVsg5AqEjAMdCo2S4FTFAjseF+PK2SAUbn0qendMGa8pnJkWd50xMcYej
7D2xxI8F7Ibt4FPugS7+yjY3uLiFL3Uny8Vp77x8G8XOpbyZTpP61Ug62Yxd3RE7
LcaV/b+E1kXnHcFv3nqn1OCz1pIrFouaAyNo8RLO9IWHaDua5im4jcN51LyfpTLx
N8Mv9maMs0UCu4e4EOLfxDx+r8/MJpeMX1eq1RY65rFoi0AWeJiC1JtU3DwYnf8M
qHi8p+XIavNxn5rUUkYMHN74iueRBNyCEGwA+JPxFFGMmCUsRYgkTVSvhoIGfPN4
LkC3n6zlzwxPYJ1tIIInDk62A8R7d9G8mL4SCod0d2dzr1f3v0GUaFqnuCLO5eoY
1ipBAKff0pVuqDfmIGtkYk3jw6cC2EOMo3svoH3u4KNMNtRwoPwqe/AcnthD+IDh
Lk6eqVCFaZLBHazeWhNzfq21iapLmHGK7NFSGGsBNUPeKvPDSkH5dsYl1sQC0EUv
s05Hr+lQTmoVcmjEVgYOSLjKKBZ2iq8gg65vW/bKATCrCqeMILIFehqjHbiSE/hb
9PbHrnfEzD1Sz/11ws2q+ZOQKaxV8O3LiqjBg1L2gb0Z7FXHLYVzUskxj5wExknu
r/V2RkRdGamSve+VzUtakPBNy3Gp9reeOFE0SAJYVbZ6wXyxiY5wquYkTRUbdxdJ
NPP4c+ulJk4uERnqCZrCt9+g0Xiy6hD0lZaToEWQXi7z+FI1hSr1ydm2qyWiwkuz
/0e3W7b3qsdol3XrAKTa3OBbbOA14fNlvCafTDfHHvp5XXTNYhkdFHX3E6z+BhwJ
eGuyM5EGl/dZGvpP7+DESARnNd44cEDaCDFtuWnPtuqLDK7gvdzdyALdPEpSlzDA
wwub9rKwkPvbc5N+m0Zi2FKS/wMUcQNjLyHFi6gc1rNpkU/DYJM1OJLB9ga08sp/
oIYf3SgRnx1kY6bl7TGzLTO2lpOyaW/KIuPtuRtlyfQYqSzsPKiUFLQ1kBDeOoKV
Y4AR5bk0EX7To3y+vHJv9+0tSVip5/iGCQSBPPzoFd8Hxzb35hnFE0rRYYFjZox3
VVTNEbGEdPWA3s6b6x1adsk5DSkmhUdxCIygujnMaO77ffFZxY5ANmUQpruuA9/9
QsSv6F78pI1o9v4y8GvSRiz/hpA6MldHGCV2gG1jGei1sL+syzbq3bfcMiwReY/m
4rd/oFvhDjEoj1V/D2Q0QmsOwWf06zoT0SP4fWcPem50gGnXD/mIwnMBifN6JErg
6dRZCnolyjD233ntq81Le0Twl9Cyj9MHSlQ5r8U1YFrPtimTp0uVCtllfCxTWJ4j
1wi444EM7cdaQi3vQ+U8xhNeIpTgrYCBBdNfpPUTD+6hLftREAlLt01Vut5XXE31
dSe48DV6j/Zd4KjrvhfKgiUZ4gqHYzFcgDEYEjKSchoI9UNVhBLNxgX90t3qjD4A
vVrGIfnsAw3pcGce8+H8lJD8Om2exW6syIvP56vpX4vA1jo+GRrNZusdzwzHa/ZN
Jurt/PJhcztb3Paq9meDUbimzMRJQeC9RuzJd+QhozexYaG1sQcbR5KdQIp4fNSZ
wG9u7MbDElr6GqV3hoF0rLW0xU5Kx2WYEODMa7qJUTTlifptiKSQFabraICjbQls
5lf2PKd8YtbNf3FWIneWmVdg19D4ZBktowQg7x0vqT6C1rws0WD1w6FIGUkTqQQy
a11CHHKLoKsV1RmOLS/4yFUgz96MZLG5ApFvRhZely/yBYyIG/14k0muJePfbwaj
jasFGI/ctGnZNCwywD2iB2YCwVU+T1VWidgRTX/vKT1Mjju49+SpKvZKubwy46Sc
93HCa5SgLeVMCqa3UDh3kBS+G5YPrQaQDZpBtCRwzxJkbjo/cr4kq6iuBa8oOS6+
nunpvb8MJEJlhTuwucpf8d6jnpH90B7tk3nufyZlTuk+OTllbkPEVxH8Y3dJsNKJ
PFHJ15vfJhkavmM3J7sqQDB9RPg7d0ZXhkzOFKyoXWhGg0rTfUTFZkO54m/Hn+fd
8+c2KUsTlTRL2l1drvKmBh5tjwFlKszX0M4N8lrsM6MBjKqqRNHBzsaQx3pvM+QB
3WoxskCoHfWBSPqdz3oHz61L8bTVJj0ChIuzWCAGJkm+hHmTsR4wNc+mqD9swlDO
I8njMNKRsMWPjKt1mOG3l6Ycy3Zywnzf03QIDESqFa3MB6ZRyngv12n7sUsTyhh8
lr44ZcKf5bCaRJll9q1nEQ7irff/R1aZfj8wDTqZCK7JRf8Gm7M0XJQH84YqmkwZ
tWzGNnns3/AJmMqczadeqQ92jeu5hl1Vo0faW/Rf4KlpoReOBqGibx+LhJMXduRT
HNZZIQHpNm9w9zaWG/5f5slUGWVBPHprf9EEyv1wvMHLkhJ5WhhdaRVexm/6HW42
KLOCJo5kD/3jvNlwbzy58bap7hN/BjLhUIkqh5/DBQDaz9h8XYhhE1bOlUQmDJsV
RxgIb+RynyTeN/FPr5+aPOo6tf2/Pc3fbIYFDMeLzjWJV2xt11RoBlhCK4uUG0aF
YTIGwr7f5fup9ClRwQChp6e0MGad/zKvO5ogYPFadPDJODBehavazoI52LqLf+St
ZKhaGZKcKvXZjwepqLtu1rycRNbVPmgC+einvYZq+xg9ftxomVTzLT+Zz/sjvFEE
RAjeJxIaRARtfvQ1+HjjwDjEDEYZHW7kTuzL48LFdVBDvXBA6JfEkdqaD6lapP6y
n4oo0QkybpPmYiMBeacZvgUmzc8TNdxEHOdcdpdGK9wKsn/R/vtkAM+SALJcAsqx
4RNrepIVqDKzky3yW2TbXP6Cxi1YOaTGEWpDDmS7VNSwkQuXDQ3Do4rH3l46Dh4C
ShhzyLLiWXiBHqYz6Dr7egeXpZ7m1cgai/cM9uw9oSU9dFTUqo2JfgbFn91v61n3
I05zC68SOREkLu0QvqJ5KwUYcyYZKgEL7/3Oi4/i9Z1tW16Wrq3LKCET4AAnqhXa
j/I65aj0vM8T6BzuAt2tZUBhGU8WIJ1MYEqgx/pLMYQ1jTsZv04hWzteY042WtRj
Iw7qjJC9+RVBvhm5NJEbvEdm5be+zuDt4eWjX4BnVllmFE/F8i/MAfoe5L20yyVf
5eS5qCEgg9NBZ6Btfz1TVBZRPTkVSOCKAWZFmuMA2CS2pD9ILFKxSjYavX+wuEbY
LJyxCtwIYRh+jtDmpapL831MGVb7+e9o4wMJRl2zJ/gKxUbZz5fLpzCj79gVHWGf
xdVYP2fvE1LwOtPMWvhDvWEEu+voPUT3JsKEu+2j+QSPVNMEfCK4P548JlO2RPLX
xQnOJ3G5GrydQG7EL6QjcpYKJyuQ7m3c1xm9+j2LETmKPUHpRoNl0GJjlA+NiTfC
OmRjuncIHUk+GfuNmpfP/q31gAUeLwDSFwAmvm7Geu9akZHjXzHC6QQFc/vA1LYW
Ho36jPln6IqX/tiHgs9LLSOxmhJ71tf+t+x79kp+S1lJQDQjrTnQWy68SuT5dqzs
UVwkq4nCU03n1cU5RtS+K39eGbALq9GV3nOO35MahyekC2CKTOOBCEN4eIjyBiDy
oYeR3LLXsOys/H9+ua5FcR1UqdQNaaaKLOfFLPQW/T2wdunZp7HSTJS+EuuCpnT6
eEY5TjvBpL71xVr+gQRrhxV7ABEx1X68ZHj7MmoJx4e6fxFAEvpw59oASMon2nZv
ROiYAcc/7LimEI4/Y4QDfIWJ91dNkU+eIU8GbXcKpz8iG/MXxId+9fQlUKPv/MOV
MHNkXvEAYsXa/lcJRkT9xCjYHIl1cKnfR7VYItIX3Kn0pyTKj2jrxS4TDEr4vNW8
jowIKM5sH+zmuqyW6PmYcxkhulMmPrer4/zN0Qr0xOf1JnBgHTzh0qNG+sy4hH1b
n2wMUhzq0hBb7LnF0jYYwfdWmgh7n8QrPjhCyfoS1a+I6bGZvGg6TRtVzOAHewxI
3p5AxW4TKOiraDcuwsShOxovjDvf8IvitXYfIJuAhuqzD6K5B53qJMmhekuh3553
SN//HHkKz5qerpHUQ8sovuDhXbENmJ7skFB4Ktx5dOaIJtx725oUf1VUZjyufDXo
WzhYaO8e6FtZPv2jQxnphQ81yQWi2s1YGJ03OQLkwTUcGL9S1sMXP6NXa9X0t1cw
YB3emAvLhqrxc3WZ6DIOJ2WQHS04rQy3/B9hkLGHZ6yK1MtRVq11hgKMwwEPTCkv
FXBl6pOsHZhkcwoUXi6F76kVvVmwitcoJen9qGRv7F/LpOUg58uQVjJoYw7QLquj
ctSh1/ZHLxp3KcgjTCyQCDiKnE88XKTOTqC9N4GR4qhRX6ol01H5Ximv/wphJIRb
VLiBN7edx6GhrGHTCp8nFEd1ZIIYPqdFTWjFn3K1IjBXs4SVZNfsxM1R41v+w2Sq
g9bucaKhKsKqg+j2YAIGkpMlPG5nYMxJnr5vsp4zeDwmzjan/IeSBKRDnsi1Kdwq
W1l88EMzsUgq2GXjDOR4x19/xbfoTRLafGvk6sJ0GAiaP8WEJ9qRpIbTgmNKsrws
Vd4PKAgalg4J/l3iahrsg06mvZdrMWXFaJys7M4oDQUtQfpCdrDnKZWTBDjySLLh
Aa6RKymYP7iyI2dn2eodWIBs2S9tsF+hIRbM8l+aH5N+Y+e/e3QbFoXj/vVpkU5S
VPWxQsix43cyOH0+3YHqdy9PJfs5FD1xJflpqhO/V79ceN7TlU99FepOpzuIjLUY
PX5SBg7deP3UqKCgXoaaqxh7MrFFj5zb6JO0c0cPCX90kcW9GbmHYjNfqtUaoRqS
vn09JFWt3d4uLQKIqGY0MeALuoNjHE9MiEwR2hg4qFE/ZD/6FHMVLrfHA+deyP4X
sjMO5qLuLivJVIBATdYpuS2BaJuv9yMaFfUqk6z/UUVimTswUdYR8jEOPwm6B+H1
NmeNE05dEjZ8dcIg7zEXtoAwWAt2MpbTXEpF9012KR3jAd85m+HFGoD+Nu9rs5U0
as0wWBLIdtqeZIfZyy01CtMbAJOU4drr62sa6BYmjxdUrAFF3DOfilDx98GUlGw7
9mXu4xrriJQSvQzXgXlkwdfRfmKz0fBljNPgVgxbu8EQT25oP7dnKhSh/dDCIKE/
pPVtC8hCPxNiQ3VnQgh5/i3LFDEjW6sE901poM56p9rxmHosu283/I5EAplkqXne
DP08gaquEzn1wu+luBtghgqLaK2u0Fmg7Tkcbwv9D8DyYc2hNybvI6aVL3pr1Xoz
JXIUkvMxZz3AHVdTvS1rX2eI42oZCvDLWd+N1nz9ofGcggQ59SpitwaeirU5+ulA
MhlvcqJLMWiy/xRpDY9HKGUQWJ02ZohI6dwqrneb8i9O6yk1A4McdndWWV8zsrAs
u+8UpqQsq/hJgAHcJG/8fQcvV0wdHsaBP8Am8fibb5Ev7NIr2WHGrTFCUFiBi8lT
nIju7lL55sWzDYhS9Bq/gkWRTllaLmJKP//gZaKKLz0LUp2HJbv9RXOCCZdWJZQl
OsHDXCcUpjdF7ZbKd7tZNBa0jQGKFZWGBA4iiuiEyPQ8lT5xFywywV5iDOG+SzLn
U7tzaBsl45bgez1DNXl1BiIgADR4YmikScsBPffwAOfOC+UGqK0qe6y+45+7If1t
0JMCtuRbZQh9lpLqsO3HWXy0jHDRcKKj05xtMyApQ45NHnu/nwqT46IOkIeYjFYW
vZ25w9R7Ob4CfJTAAu6g0lEbyvLauNWlDs27rYY9ZhIi2dVrPDWsu6InHheKu1YC
R7eJxee2btd6bsUh5dcnPwlWyODMrA+8lnK+AJGCuZy11yBVAhzpybw3iYz6R1fz
0ZtbhcaV+6LaJkw0DG+5Nwv9RTx1wxlJ0UQpl6M8h/33+EK8N8phKOQGChTqdrFW
s2QDfQHx758DZtGvwizXt1dPubsU+M7dgZazsJQgDydCqPvylA8jG+kTpczVEo2n
S1W0rVzFKRVebKtTysg1eXdjNn0WdU0KLR6bYCrEDGRCw3I7802G6S7XovRTDCK3
Ab5aGmabnGmB9MybQx15NAc610sN/1SXTo72FA+W3GeCGqDmuLT1wUdGoX6NX/N0
wlrkJVJXD2inx0RMKORZvYwC3Yqw4rNCPGDKMbshD5FRNcXeJdp/U2v5CoEowpki
LnCFdLWBkbPgxBSnIITHUvpzrGq7tq6gRIYjMYXwgUVX9vaLTJ8DnkpoMjbgaWPD
PUqkb9rSsvF72ZjgwhOJQ7PbIeR7+3SqJpNKaPRTWt8fEGW8tGufhlIyrYG6mbu5
A+ESlIVqSFKYKEy7TFQ449tnr+EwfaFOfmpQfbqsSlL5kGZLdvbvLLp0Gvv/vkO1
ejt+NZZX5f2SDnaNNQqEaAFn+1TzBIIuPVLaSC/4R7RTrsJD4V3Onpiqz2Rm74Od
fO2/zfT7kutnXTSdCIjXX8xVIlKCx/0N2KjpsfYju/+/zigS1awurnsGOSTelpve
FLBaFylSgBL1WNZiCG4LslKbdYYN2yHzX9fZG7jBSFk9Dsv4mPQsUprpFlHl2TmL
rL4kTQgAwyhBKEofrxk7GhcwpHCJKHLg3H/kmgF1oQvnebwYEFxZh41V/mGdIWN3
G8LzTnR+xIi4k4SQtqjj/VSx++bdSDneOmCuKh/4ZkXAiXVbTtzVac8T5l4Ibo2C
nvzXn5lftFGOpUU3ZW7AST2rxcUVkJfKr3hyb+amCfxbTi+KJMZf3Jrg367c3f+N
vmooAjTQK3dWA+cHL8WvFgNuEcLZTl9efCqRFHgIu/LebDsGM/avRgXS7/0TJfoD
E1CRWaL6zm8IXvE4U1eznLyZyYHbkOKXKz9xDEwI/ISy+OZEaj+NSnPJq/NN/m8M
jpz9pNXRZhr6lMfqN3ADUM8ncQYCokygm40Nmm9BL9n7BOLQNgmSeCGuoQyo+H3E
7/VqwU9pVyW+IrLn6flcPSVyk9cczHTGbBiQ4N1lcXRecJtzr1B5wVu8jPhDSkin
xWvUi/W5fvs5iFWjJdDDUykc+zE9t2mtkp+UJ4Y7hTwFtXtNl7CyqbSj/e9JgGbV
CAxrWG5OqoSEiPcIDHlSif+olss4XkWRy9s256uMkbCg4el0IRarrnKay8vIsdwf
fnV7fJkB4FjetA7yv6vabsUTAIyYld6IE6Ye0aSWEthDMPl7yNFeziWqvTwXyrzK
B7dmP9UFlUDKG2Miq1UBVCUqTaQUG5Cq6WNy6PfzC0rozul5uRVMV57GNSItGSxY
Gs0lSUuK6GlOlqQdHaZ65rkuKPuNdPJQYrfS/uXW7uOTR2IZlqQvjeGXzLctwsdT
rcf3qBvKnXu+NzTyqyDVVVFe/SS40K1miuRIs++YGx53fJK8jMz0DSdbed8apRoW
0BRQ368Z6iCBVk3zm0nE+xyR/hWZTDlyaR4r2rFhmtsujmdoiNVByEa3nQ5uwNZH
vwJ6/C9SO+gWplYzw+IeZxliczv+wx750/f1nTXIpd1nYdfPBY0q2PyEQan741A+
uJS6SB7GnELx3FeAF0FJJQ5YkuqGe7ysd5Wz2tzse1EXB0hrcukj/F7D5ot8fWVb
XBb0zFLT9TcAjhKtUrcGDQ48FN1Oz9vtpEXF90/ccODxwXMCMCnlLucNU2JdiRmp
2ug693U0H/6BD+uBCssqSrq2aZUrJWaxXPsz4SRR4dRZLWTYa8fg47F3lbggbeWx
WCdCVqVDqCg8ibwyxGpU6gUq7dzq4NWaw0nFgsMDgplQudvNfGGtG756sHx9w9xM
UYZnOs8mq6fOM+t6SM959xxR0DjFhHRSa4RvZACwuFQegztibe/S3roy16nhYzHQ
49Yh51mshobgUpzu3w0GLxniz7Br3fGjKdlavCJN/P4Uwo0fwjViwZrT7e81pzJd
8QXKQ1PYN7r9W2M8+ADnP5dk50CJ/vjMS2vF9fTmyO0SufuSftyuDdY1S6PH0l4T
LSATts6Hh2uwcUTPX1L0nDeb4HC6HdNtBLsBQOu12DhREFxRorO0jg/4K+Mtek+O
SwmNulNkBHtve3RqayWghhkKj0ztZt0v0q+4zN0VCMwmCpiwMTDLogzFcLtYsDK7
ofnvKkfHFRqJkDk3vUh/V+vLd0Cot66xtn50z6xjbrhiHWcmiPrUsoPpZ75zzVj5
Sfjs7b+kDyWg7Fb6TXTgHoRTZH/ORtx36v31GXG3zBAAfaYL7kLqLgG4IyWqyPFe
y06EV2yO1Np8IuBPesWLfBewtL4Ccejj2LLVjINpGjMM87jsw6xQpMy5g9SJf1M+
mmwg3V/cJWKTZr4kQlwtoHJFTz8nIrnrjSUJgOaF+N8cOLc6UHMuiQgc7/+Z//5B
rn4Ad1QbS7FUherBqwmIBUL7SZimPnWsuGjFhWISdLFtkZ2Y0US053A3X29+hPK/
+MKw/934huRgwpFTYxLkDl/Ep7zEQnIUEMm2wEU5NgwXc0+G+EmExbgARoTrRwP4
w9WbPKLgY5rEPbxckNvbkVSMsVaye5GWTQ4JWixOSMP3iila6Y5m79cTy7SwWz36
4cCadPkOV6oqIwIkOUV0B248uZr7Tfkm7sWmjGDTpaK6924awGC7aHfwoMgsBTWo
lrPwP3Ny2rCshHhmwbdSKL+wEU14HC6fHcIlu4Qgx2MNFYJMrdvNkLh19DYA0Vr8
PwjSsMt2ZOwxffgZfOfCAhPcB/7NqFno1KfjJXVBiDggj5VsGZuzS0EIRuWKn00z
z0ltAn+2jPQwyq3HODXDjD7DgPhRhlp8VXyHKk69e55bzD3vB5RoOmmh1P0p1QGq
H8w0WJ5YhWZ2jJf+tDgArMjrdqghccnMYBKDA11yskvYvVugf4fWkEe0+w3x7hlw
pN/x9W0JCQF4TcggOTl1Byri2xDetz1dsI7YFMomDqq0CdK8sjjn1qgkxGlRq29y
LqRSDAC3xEZ4xrUzBMGk/rv4u3mGiDhdgDYRN+uMNNxK628L14VyzfiD8XO7JWZz
x7lqUA8N7ZsDF6hA/sLEE3Suuo2Fntkvcx94HuBLxDggW9wgk36w49Y7j+dzpgZI
RdbN6LPVAFUzbd6TzeiJfrxwdehA+rgrC8nRwGcAwTzsNpqElOOggSTNvW7JpAbP
hNOURJytWSUVooSea9v09x9mN285ysJ5UkTSmakzuJoQ5WzPXl8WZbaO8bKI2G2a
vMMMzogsQAb+iTmP8SdZ4YhjGooovN8QXU7EU6SpYXInjWvfWzo7lic3qO/o5oMV
Fc/+4DQItlcuJRfUw5i0Y/nf4hTGmsn/qzVNJvVgQYOQHtOfh4MFsQ7B7h6nqnAX
ajM0baZkpqQ8G32RkyHl6W5w2WUtTVSBPZFo7+/blLMlmDD2UYVEyVhyPvHuuPTx
GFcg44dVEzP9Wr3IjvWaT3IPaxKySI9eUPbmCtwhcaxBfxSlhqYleyXJKORmE+v6
n7HxyIR4M/ZubJlBkQMcY1X4qQ7cbqwmr+aI0ywtYz09brBMaZPGxVt1BSNI6CqW
LajLr6OB6ikkbgqFw44MzRLJJqMm3QRv4gbhLNQ/AqtTptesbO+JGh1Gg7nhn5sR
2zStF+6BViazpBMy7rj75HnfX8sQHLB1JsmkfZ+arIcIqxrmcaNfgyN3G1/rr3/M
Cqv2kyaO4juh5LU1sCTgSkZPtBgRLrnhymL2ttpukO9WTCzT/pD8FdioIZYZCHjg
yI0kqQKMkE1utZhmhrH7ZI/pij0+vK+bh2TBypzmcEekaQch+pTnon8IJbBZASyz
+My4BrIOiZ215aZTaMrLeX58gNaeSL2nNkd0s0DdFSjO453nZNP4kZjMs5y6RnVe
NEOrn5Qlgds7VPgXU6UK5Mq0sYfhojIXMD+aePeAX8PI+V1veZPk0gAWLTMQe+ql
ZbnIAKyp3qIdqYILR631w05/kJCRVB3jOZTEk+qqodQBzKCRjpQlyMnzdYXicbRP
VnLvx2lk/6JnOXKxFpGsY7TX9FjQAxqVkca6fWQkQtyWnHtVT19E7n7RIoLLCbhE
xtTaiG4bKc+6U0E1XJMjuKmDFtgEIJ2KJ5GcOuHBjpHcpfSaS/hfhBuNNCS02gy/
DH5laNUj9PFsCYmcwodMMiSMgqljBQX2PvR3PqjWACHRXk6hdvuVbwsWApKvpQyC
TgBEAa/xuOgB4lZeWSAuRJbORcktVBVp7k+SujXIMyQuQn9k3pixjZ16J07lIBQN
XjKIeHmYJ9Fvay+J5m8Og+WwZGqNvdqrWSil8sFh16+u5hkYAn5iiSeCk+4Ymruz
XhYAtD+dO4vH9S9wrMNkSHFFJbkiE6ye3Z/Vf5LZOKUlEabe18FibuVgRVY2cAKA
8GwWcX6ByUWyLlPq1LNd6rnf0fgKIOjdz1a08TVUbYQBAfLOXd+XbU0aKHpkZRDC
V21gymcRvzjOw1I01zGB3XnPS2bpY34wW5pkiehH9owlXxxMaTJ1R6+3A73pDPzY
LJxvh5hOoKsfckEdYz0MLTGDB5R85teSgFL50mYNMTjQ79HrLPShC0GAPH2TY2uu
bMZq2jysNkkZkgnaUVbS063XJKBTuVvOGsDfCjqAp1hT0zbLhZFbOWHxyaJLOpmM
0FArISLzO25wsLHBirFU2lWbCfnIolOu3oSCishq6aAcSF6SUAIdTy5eZRAus2Fq
/3YJTvHrVa7/Rxk4AilP7CNwz31yjERQh/4FXNbBsvnn80uOVHN7dPvNlZ/4I9tP
1Gp5sfFxWz7hz9mtlBKPUjXfJXJfiWYMQHmoJ8DQOGN7uHoooTRHCiJVnJz4QAyf
gGa5bUAAqUHbkruiFWKEC30vWCK4FaFt6qClaj56SweqteeIY/6/5KHNCqRh6FmM
ld3e6YXvfKJ8Mn9uOc4AvoMTDXu06ZPPS7tBJ9va22JruaIzyAHH1UBUfXtjFOsa
RJ3XjHM2g5RS5hvucrQ79kdsdCvKAejPDPZvp1L9sZiDOjwUkIS5uuoezXbMuC6a
egNVWnSRrG4ho2aU913o67yqAnRZIP7olRoSGmU1q+p0eKYbAPWPoY41Ofd8Mcsx
6KVb1XNiebpSjLEHyl/t92Gt8XcIj6HXyLOxFyXlV+p3/u9P/TMzXLBoA8CtYKU6
jvugPSybp4QQ6EWtKtnt91Ke/CK/J2mY3U1Vvx7Jr3HmVkxPZbNuikLmkBtlZJ7w
ZQELsHLSRfVW748Vtlt7WoEFYhtVeC1Nty2sgLEEdwed+IMPpEldTEeB9JzwatlL
W3HZTX2244eRzkYLc8FzKpQwxMiVYwlFawuRciSGI8ydYnNjaE9rzeAu58vftQe+
HdJN4Iqsk3GjdH269c4GBLqz54EOazwbJsK7uWKymx0uDxf26ow7sL+1NfHNDEqS
Rae4Tpd0feZB2pzGvoUz3aWphKkdX747R+FOG8PTFinHuNgBaQIJk7ZUbA7IhCus
7vAPDrFXD8NGXL0Ys2bbQNGtJcGkyx1sSgW3bJgLpBW7sZOKP3Ti7znQ9u1ygYfH
QtFcIBG0DYJzgomJTlzkNNKtFtVSxY2l0r1HOsffeoFuNJ+ABMDBOhVUkwmFnZ2R
/IWYqdPNXgrSjltcIGvSwqmrZ9UWibMdXVFoJGnG/y5QDPiPXq0BojcBwcz1ButD
QXAAomGbXoOF0r+YERj2zoYnfNgcMbwYnBUddpx0AXAezc1gKJtrOn8adMVLMfEr
vtS44EZSWWlhEjDdo/voz77HHYTKLT4S+nlgJpZ8cp1ktsPspRzR9zNwe4lGccvc
pe+zjQHgVRoW9OsF9q+z4xogS1Q2oDYpebH9HsLBHpx9iJWd6B9W5R8w28iruLcj
yxTrVVcMkmK/OukA2CT0hgNcDfbCJREL/oA7F6pYzHrIyiwT3eq4vY2914iDgaz6
0vKCsz1W95SwFaoq/MUHNPTYsAvZ4+pNsGztrpkqGnugf25X8ysKpmm9tm8vwD6k
H5DKMI9gIDIn6M53E19GlajUmN4dBfWfkuknHVtQImzWNWkC5O//emRswSKkLTO3
YTp3hJ3kAVuhNgUK+bKNGByr8NRQu8ICVf72afWlIROZwqlJHRcLo61k3Rsvqmdq
fs2LBycRcpfeImKx84QMoLufBJAXVcGRzSvV0GkRHx8/Jg5nCXmZrxM+oDGoYc+K
ZWrjZ8cC/Khda2tk9/x6MiARYpgAwA5LfONjX5kOFCMd2r+0L15oObjNSgXkvuoh
rbgob/EEWFuatW2pMC4K/ZMfkL5deM7wPPue8HGElnJa5mgdcuAvkIPq1GAjRLOj
nxEAxVfWZA0QnfJJWRdPSyFrqMBy+V6sqbcYE553Z9WS5tbRkD1kqWYCnB3f7/dI
sZWfd6j/wAw0zHEDZw0rU73zxqVHxDjYgGVFiIuSE3okzCrdY2w8jzxnu9B9OPsk
JJJ1oDkZGsy+sH6zm5EsYyTejsJRd8kmQlZUT+/zz2/UhjqQzRu1e78XEKU2hM8K
CyrFoB8p9iTJO0q6a849MSaJM0HB9qeepWopvmikm6BNx6a8PW2nJucVib+BDraS
mFY9cWdyrXewMlfNjHK1Oa/6CH45M5BIBdhm5G6wTzeuiEyscB6RL8Qg0UM/Wf6X
ljSfoKZABL2lGUcAT8KZRqyqYHQuyFWCvlow49a11NJTtwCUQ6UI8zztg4MF6PwR
ruYzLPpvQcN4PHMACYFbcQfRv9C97gPMfCLn7gGTwvVXhG/IdwaGcKRHUygJyd+9
DTS8axiShpVpfg6ZFxczwi2Z3D8tn7jL/NJtjl9ZgfpenEWzZM1ZBybmIPvraLal
4+jzKsCVyHpwRGeglnA7qlqWtAmRlZIjt09ie+jKOjoyebd+LR7FjhEMxKB8/Y4P
MSZy1sj/yTTp7najrTxRNUc11ouHlUbYn74eomD7NRB9tRglwOsuupebo5ewJlx7
EJ5rGq/V7yaN3JjvUTDLBKPkpG11FG+2e7kMySawtEEd5HVPGKXSvB5esjLUVVe6
j0Iz7zPns+YlUrmIJ2E5wp15zI+SGcm4QpHWP88bPlc10IbHgd2d11VGMQV2IePr
waVoJRloTroFeJ7TcwBnVnRRrvzrnb9pRH0aE/m9sg0BRTVCDx5eq42C4QZyh/Kx
MwMkzkDJIbjt2+aMxkfKEL8v4pt6a4jDEhSegvdn02QO7JGngaPt5k1evtas+6lv
mmq9dqLGSi+jRsvVVAUjmtNhfTmbjeqcMhHJhqrvHQtcY4k2NQpdejcfmeSssmtf
eVFi/LtiwerX0yK2rVvvVRooYEUysTuG0EPRu6dQKE5b0LyIU40+pbNDUK5kwb11
DgMlKvuflCEk/zqupJjzId+3oadKXE6Rso3n2zGKFfmGKkASu9LH7Ki7yTAbJc5j
SWP1Agk0TgmYM2xGDRub2m3VXgjtqwEuPkYdzeNzCYPof1w0DQjOLfA+Sz+j/o0p
UeTLb6jMqpdkYfWNpGAaxnvY+AyBKyVp3ljZhDqKHdUMIVAoDF8kFZ8qMwc+DjbX
2sxN8Gp+c5nXVug770eHNJheum4SRcjsk/m8551mHxBbyXnjDM1UZJOk6K54u2Kz
R0FizVMfwJAwHfy9LK7vg5igQwoYNHT4DSIehWPGNvWBWKZ5nInarjiHZbvkISqW
mqtY7DoccRHp/S5UuIYoqL5XVaPOJreWV7kUHgrrq5dIhkS0SOfHhnWypdoMmFVZ
Q+558v/pJgTohBwdqMVPyHFbZyHDSqUAHmQ5F+wOUhHlai0xcyFvB898FmBNOlDZ
cUqRux5CS1eD0X/EX6dWOVxfSIEybRbhnVfAzxbo/3NffeckI9TncoW4rFSck6Th
X1WlbYE3IljvkgcWWDL3ZmEYiSUZMUut//aofg0WyIRvB+ddJ3omom+CvhMuAZvF
ElDJckXbp3IC9HMjPMMEkCfpmkr0E3rZrSe3ZMCQP7Qk7OXm7uM1TkyLRDfHfX3s
5mJx8HEAlfvuCztTmEvvnhXX2tfQf5pYGwTljAOhXREmn25Wwrjd0XY1Csb9jlLY
/xUoD/r2r+cadOBBHaF8+K/aXezKMkviAvk154YuTHosBXkpOFBwycns91pOmgc+
cGwe4w0fJQT+3gJLukgIJU/IcPJkHPc4jf54aE2/q9ZBaEMFuH9KsBcFEC1izViB
rOWSeOUhCaHSfRhhDJqhsRP/sP9g+JVtldS6W0Jqjh+NQTooKty4Vn3xoPDAiyHw
3PdUTHi2r05S5+kxPlbeDD0dbu8piLpFShBr9uiWrpWzQdN4IaimZIyRYtEkFgDm
Kg2e+j2Kr8HhxvrMx9oNMRAZSzfXOpqe+Gd52QAwRLYJ2/8/ImAikRrvABDsYyaz
AyBUg+D+uDrKDurX1NAKpdXl9LQKWswie4fHwN+Y1D24nHc5+6NKldZST88CZgbw
dp8kM2QYUKkLL+WxEC5ZXaMm+3Teow+mSC9WH+fyNBbDpLUVfLJzcsUMne8oE8S8
PsGCPhvqIIyvUuK/Wehw0PTn4RGVaMnz+UorjpQyeQ1mTPBawpykWB5K2oYMl/uW
63DouRCJb6RGVSfiwdfSn2pn7uKyYtSpF+bCZaRRwmh94aupE/cQ4BNjlMcZ/BZU
r25S15/SfsrORKb5B/PNkW9S8QclyapghPT7Xb8t+N8bVGG/zL8NavKAKqN+D81V
TFy2rqIlfZ05nHI51Vv0TSzJUpAut1nTcFO1C/BvrLZ1ZoWJ6iJzLutv40cKkAoU
9hlhWxvtRyhVEYiruGPY8eYvlicBvt2u4Uze2uUbbBy0MNiy3yPDsyI3ANCSGfGl
6lM3nesYeQKbldQk39hhVuGhvbViC4Ws8GUsMmLMuwq7zZhZCvMP/d3cEqS7jhwe
m5REQQjXZxqv5loAZyEW50o4tK5Yfiq+gE6rcNWOEqJYLT4FgNcceATrPF2KrzRl
NaRNwzb1jFpBATKo5gi6yoHPIjY4gDPsP3xiVR5iXp2XtzxD1RdHclDl5aDtJ1LT
/qmtu3krEvfZU+TihFB9ttTgc4B0C0gIwLTl3QYgw+NLRVFsU5SwxfKM9MnifUca
no6xoKptwN3qJBL98MU1w8cD43jphsbIffO//icqUrI8L+XtNDCP1KFAQ8S1s2ZN
RhFu0aG12NGkkGU6UBhFoixTzxTZ3GL97lsQMz74bLyEF/ZgHjMHtTYL50uWerCX
cgx3vZXQJWR5Y3dnZQcJFweirtwFWhZtdp5RDe4VutXX+l6Hca95wLaKHvq2HEiz
C7bUZOyA7lm3GceERivYP42k3u1r5oR0PEb0O0tFbK5iib6jf3sruf+QMZw8itWP
FXFbYAjhApgfbC4L+KSeP1cn/OggRwresawT6bSShdeXzlXFYf+pYexdYu3t36gr
7SrnzfCXKoWQG47uEBeWKuxfF6tCoBWZN3hUVdzqnneVEtsozSzFnlp//x6hjFqe
hVqYR1XYrIfHb0XLX7llkmFBWkORI4p6wramGDlPcQku8aTxPthcPyvaKrsaUhdT
wWofBBxz0Qdt4MRND6Vl6qd5YFogEJDJoAKQe7jN7fJa6PVG2+w5Ms4WGWlP2mlH
E/BEizIt0F+r2Otsfr2yUNO0n0VGjGJoqQ79C0QxUS0ETjmHT63GmJYBY/M6peDh
MVzwmLDCTehwrlN7x1Writ282vRneMyLoC7lic5vDbYw2wTaUwlyNVYZjiVQv1/7
yqkIfo7R9Oj2wfB/X7ow7b3UpRgLJ8g297I8XGIDrdyhB9awCnAcB8hHxG4MqYaE
G3nV3QS7DoSWd32LVd4Mr8nsnEOqwEep5ZoHToYUcJ78R2BoHHbkBom0WSzNGtcV
YQlQrjSm9wJmk3ofq9iZPe1pBc1exqjOQ83pxkrabsjEJZeywEVUY514/2NyA6yy
KSpZ/leIcagmYCgG2tNsFVasR9orASzLvham94mD3gkzy4en6Y8jNHzEfXiNX+p/
x6jJEDa1WyuKtNS1Iw8b8/xHTnMdZnbGltO3TZ6nloXqSx4cNb9z02pWLaoxyECc
aA7up73F5/PYjRN/ga3Vdkkt5ccPqx/1is1y/6POXqMpQS0BW7VmzgRu8mntfkGk
5I91w3eehybKe4zVu5UbhuVyH08WEuXy2XwnVfIn7Ni7S0uyOpsMFgcNwtcfGGEU
bkFRAw8xjKtX+1kSJRGFzQkAMOME0iHgMRwZl8aIN8qqsjmvYwvebF0eDfNTcdMl
5OMyhsWOV8TrAgC2vIdFtluDpFEX5V4Kc8oNb75F7m5IJ1cDiEPDLzq49iMCtMbH
+7DoJyiLkpsRhpwLUBblhx/OtO7S4Q97+FWLA8RYlfQCC6cmZg2OY1RJnROaGeGn
ZyEf5aSsKzTTnV12ZAwxj9x+Fp//fTbN347r9Sslxg9+KA/LifiEYxfY6TUMi+j5
gD71uWzpDHauGihWqQ3KEW8nXiuzsOMjH5WE6ICheBEmOZiLnWd+1sIw4DD0a+iy
do/iI6011kiWVDAXnaM5D/SK6eHnI/Y48aMCBdscSnItFfeitkD22I4WK9PyNSGy
h9WKXCAJw7zyUMF4MuWYxhX9/JJqSwWAs/pQ3cQ8lree6J8DhcsD+ZdO0jD1E8Dy
K9yyBgO1zWc8sMmFvbU5hh55iS578TkR/hVYhmDM0fLg1MQm49XO9CdwDilnenvp
QDqHsLacMbUI5IFv4x1z5MX4UhX5bUoDI2giVIUDgxPt9afHarGj4S6KPYD2T4TY
5YU7AaSppWxlkc2/IVbgYQ2WPV6RDqzcLaGzxvFvx8nSgsaosJKqkto0iB3iAkbg
wjcAp//cAmSiUemSWjFpd4qhk5SNWfQbgiv5WLi7pQfZIhiOshbuDdt9yTxtG8Un
6C0suXXVTzfFz+cxrPGvMtzE9bQ436bwzHL6QO7Twr0SjrEC0Vmeu+yBpFW09Trx
EvMjdL/GYAJk+TEePwShT6BdqW3buKoWR3th7SLYcPgUYS3kZG47NUCh2vtGe0O1
jEdHBzL4NFkolxqpN2E8qByAPFIXbk3pCPpWriNwgrd9zlDX6tG+gG3+ZEASfvJX
C6WdMHC6qtYILgoUyYVXMH0IPR0cLKBM2bWYmaNzpcaIJCmI+vZ8UGWkBNL38esF
SgCCjV0iH9P61OzD/O2TpsUOxF0m0pjbp9RrInYgSv2quHZM/gGoRIudgHjc027F
tvaIEsIZ/KYtMlDXayiwLZEblehL4DpGawfI0eExz6sIoThDCYtSqPgAkUK6wcB/
r9GEb5vxyBLgAdwq2O9EWFnn1ZvXmld7EiPB7NHsTpxs5l3qXj0XsspA4LmNxuGs
UdXQmHdxnTDBb4Lgg+QX1IeBrKvA9WWFfsCfEx94IDOYnnrWX8tLg2bNnXIR3ST6
tRa5pxSnLFdEtmVOeTwOtIrYdqfSlAozU9Mb95/UErLYF+N4XYqupuMU5tL4FREz
EmWqMA3tDamEbWVB21JV2XquXHRYWiCJi9IDi7vKBAIOlQj1yBSk/DNnbNWX7Uom
iVBaFX4C10y9a/YO7RdnQlk7DH14tKwy0uF1COWuGQAuKYpxWDLavjmTUUxxPDn9
dctZqTU0ULOC2Kv06WbaKgA8QxR7ROccJ7a22Y91nzrPwZXFLHl+rt75WDDCDWLy
a+NoE/VFyYTXCiccu2jlwNpEyPJKg0qbopdo0xuOrKqMS4PelF8qezttDn9m6WID
cVYTP3vM1lBLDrIE/VSRLrsmrZja/RVbZGezgNXdUgd/NqqEPfv8jb2A505if0IV
9jW29AYuemWe1rMmrqt8QYH5NU5CBwcixhVDS1yU1EGxjCpclEiUYMP/9MekBCmd
e+y6BjETK/IhGavNO+prWJOB9MAKlgrJgLA6a0whHrrnX0HfiYGAlWnrJhQozpc9
ijNfciNxky2fEB6zT1GugrG9m2FqHAPLjgIz2/trnKWUQeMEfHvGe1n+E26Lco+I
hBRIZj+/4fBlEpEDnHe852rDi//xivJr5REsV0XJtG2M0IzBZ9BHH0P5AmTytag0
JRl5ENL+LKTN+lziGxfLvSi9PHHAH7BoxOft/ySf0FhV4nuGEH0hppSExdzduTvs
vvxhz6ikYlJULA1HFLpSA3sHZu9jxld97+gZkhIXxdERKUBxyEvosjkx9nJr1eQx
DNRLwL8MFDx1PUllM4DfCaBRbVSPuwxospIkfO2Fb4WNmYIoEiw3kCmoy1/Fa54e
2HyqfWCzGnwUOXVIpo5+70D7oG/ONffflHBa6upUQ7NpUEHs54wZbQAI/VqFsEOV
2p9Zxcy7Zx0VHwSaOUtQXl+YaLUa8lCqlHuRS9owbyIwIN1QJ5oa34lxhdf/dZnu
qY/Ww2XAKMM0nAuXLzhJq6E7wEPdiiVgiwDm4To5ZWefxd9+qjIYjWRUBpvYeUQ+
2+xea5JCdV12PVmB5jyie4SX/ELq5lJclSsFntDBomuAErV3Wuiqbb2C4vi1vuWN
OShWE/E58FWqUKwWsj4Rv27gRLg8KuAns3m5iazsTVOP8ODkBYM4HPf4GezXf7h6
rlsdhxWlcO9t0fAn5tsTjHcxY1dERTPA3VdUaMitDG4ePsWPVXi6MObHl6odeEEe
SIs/aIQ7cydPsjgJmUzUqbk0NqnFAsXSC1vLKTW6R+eGX/f8gHUZ+PGtMYyFxJEJ
lItSYwAe9YR/pJHmwPuMa6wdNErmMeGB9vmjjj3WIDTzeuJffnJHGWaTudUVbujJ
/j3HkdXrXLVX828Q2ygNKxDl9Zq/vwAU0Gj3X4jwJvGtAr8Vmo9M/Wx8c7Al69Da
cErbtO4cURmmo/fsj0Hw3uYoeeJYqGLFUyeeYozhGZ6ic8VqYi+MIlRqQ5q1sk7A
Us+vh67tKJynl4AI87pXbtQtfhpExsanA7q8BviqhxhXT7fz7R39nzWzjUDZkEQA
QqiH+U8WTkfbyyTRPc6QrXjtbigfO/LXikngRqqInQdcRn2PwxhXSU60CGe3P9J/
z1OZi7wOeZkeRtnoa1faiDsvrzfzoyfw+//ZoetjGXh8aew0+Vy1cO86bnD+/7Rq
c2yuoDfF2jghF+ulYNOTIWMPUC8Hhe0Y9D01GWLsZBVjoIh2zOrTeUCYQfk0zSEQ
0U4ED1X0CTh+BCitpKA0y8gLMaPzuRyrokS4UsEjKJGVyDDwxuejuowTyCCdWuOE
4KPXFGeArEe6retjdzykI1Qn56Qt6NzsZYNgMfUqHfPQ7jZkWWwvXzFiufZiNLgv
9PykSVncvi+f4it4I/vD8fubAuc0HZGF2/TRz1V/ON2FDrW94nGyxg7Ukii7xoYn
jvwF3JCMZN9M5IubNUouygXcn+UfpudTtQTUQ3cETEarMrTx7/QPRlsyQmLaCzjy
aWAI0YHYq2uTrGU0kqm9cDwaMR2SN9A2mOZZwYO/Z0KqxSccWmP3vC22Pgg7vxqy
1U1kBzNYt8DrFSk6beQy2m51FLqUlopYzMz9QjROg8afpubDxkIg+P+C6OG/lzXv
bV1eiTCVysJ46yFzhulUI9OKa3r4qvDB7/7wjNjug/XBI7VXE16NEFWGckzobv/y
oNg0j++DBZUI6KkNby+xuwLm8F7xzXEPFnT6nYrzvz4qz0V9rjuJNQePftlVvQqd
T/W61jESjVX1ldMre9zgRLZKddZSi87aYlVAuk8fr2qUGz9pD8AilZn2c2xS+9G9
yPOqbupzr/3xOB5nwteEnIZp4PeDqsoeY4Hcra2peFr283d2hptzYOoeEhRU48fJ
Sq8socO772BZ1ye3h4u/BckRaLeZHgFhFhcrD7P/r8ix9Vz5Tl5pzSWJhanVQVZk
VXjQLH7M1EspoEc/t7D0vjv/LmSTvljb5WKzHxLhb8uU+FR4pwRNgpn1GCtHJEiY
CW5A6lbCcBoLoRDfSQvKRmTobGSGpFcHop4GMvaGjCDtRoxrJtaKUF6f04mK2dcP
MSmZ7cGVRC1w9D0CI8gprtCu3CT61gokLMTidcbtfiHJEsbF6r6dU8wZU289WJF+
fEskExY1x74pVttUU6Q2yCmWxJHbXj3T6frLwwpYisfmIoa4ZwCV7woFXCrqYmdN
l4w3DLFR5TmJZI8hlQUgwnXVnYmlMVImQxU9+PbGosSHWsnY/BrJZV5TiVyIn829
YQS6SO/mObtG6vTWi65wxIE8Q0aZNJH3TSC5wrQX9zLvTfJdr9wHBajGHeqZRpqG
LE+K2wU+eVKPOvft/DHir0jKQ1RqW+4D3AIAp9OWuJC/Jkf4+yxM0TTRLp+3PXCg
njLYNhQQSVV1qZwaEnRKR02Juq5bLVHb77kVcq1CkiiedsUVXFoIIbelhzB8ppWJ
MrHR93IpQWk2D1Gg2zcoWthSeJdmlhhmP4DDgLiUkZ0wT/2dyvuHpYHUxc+sRDEC
odkV0ZAP7RN1m4Cc2tahLGr3C4GCPaagzvOH2iE7ppPRUw0zQRbyV54WRSIiXr7A
yXphZFbp84tNBfDZA722nzdQeCyMPu/mDmu4yCNtC6pMrIl1q43fTWZKHbiJH6vd
2b71RwznH2svQhz/+Gi+a2Nz2NbfpI0RKZ+IyefymiER0ln2JNv7yUS8sXe7cEiS
zvADDdPcwvVOwM1m7LrJqNSpepVHLzhQYLV9K7VGrxDfHtb7098ibwgZc5jN7S6U
j2dTBcb2YWg+FsoHfZAw2HV+0YGOtkLDlKR+MtFM04aDO0zKvo7WmtrJawjHPzQw
7+hfJKyOLH9lCJHHBp6jRtbNIWw0pGk1ryyCAK+fNkE47FBBab4o1uzMsFo7la/d
cTjUFo0yVhalzAWyXpBcFMdSJZn6FbaK++vx527FJdpZ0JcFJLkhghcZVV9aDWky
yAvddn2MJUplmXfkVeQf9BrkcwAqQvSPc0BN/VwK96eBpiDmP3msPXtv07mFWvHG
WA9gqJ3W+LQShUAlmirMy9ryGzzskcVEGFUVgpGZ9UuGoxQw1YyeKKKqA8JOzasz
0T3Wg38U3JNBTve4tyW35H8gjplDu0e0lm4KWj0UC0gLz4CEGdP4KOmYSIqe6kqt
vFj+h2T3ovW/X0lxI12VhY1LEwyNbq5RkNf2sq8pdG2xLcf01EGGIOsV7PLw2JFu
+hVZgGr4RcNOMOW1/YXHt933q7p7QIo5fz47xD5ntMjR2LFWdtZuLWd9BAaYQ+Ja
sXRiUX6PVyx7IhdfA9ytX3DkmjoS+YKQO+EhqGHFRJiMhBsSFlij3gCmrfNw3zSF
DXLZlAx5foE3CS+LzQXq3W+rGE2qSAjV+r/wuckP+NMvzafiy16q5uGVPtpUMSBA
eA6lLjMMszcOjk0oZiqsHDpaAX/YDxrmfTaFZSIvu5QhAb1lHiCZL5DjS5+RhL6R
cWAId+8PWr8fcCbdgRAgbfacpYv8Yq9Cihw31UU7O/tolJ2xpKZXUO7p2xZFZ0cI
G7zsMbF0+TWnRx3KtEhIfLzCGbYySKYJU31o8HArEXNUDk3Ihpf9WRK67CLfmawk
BhLdIlK2FEeYTFiebQoyeSeb8Gm08lzIExenHazxOtM21aGTE4lnztHz/WXHgCbA
6lLY3plP1Yor3M7Md7MWP2JaIdCUZe42BZ1ucEsI02o8ZDgW2JyEvJaSk2htwfku
eHoQidZ4EO+AHbIeXsLSPDGhu3VgpS+9d3RmU8dCsuaprOOahkeWhWunELPPMopI
iXHk+FRqO+M7IuO0O9I46xB4TWbqfIJux2QXmsgzLNAdPy64DmzhuloUKlGeS8Qd
pcXEu/IXWItcc1/12Cgh93AbH+UM1+qOdM37yHnWt2e2Dyj+Tb2uL4xuyoJPqCot
UM4G+t0tpj3hD1Ghzcc/zPCO4CUDRb+Nwnr4xgfK+ukzemzn5gjmzNNIn5R9tdWo
8nUZR3i80TI9J8/yzGtRxFvY7DTNCLQaKv4QbFOn9g1iBVUeeAx8kWuZ9KXhO/7u
hgVKzFCqCLOVTCP8aBAzOZq1FwI5jPl/vOPCzXk1M/NW9eHKARuIg4/2W9go9RoT
bSLWIY3KMJFOLX3o+EHjTZQuimuCvEYLyq7NR8gZELliF1nsFzkDQu7OaNfakOmr
ExtP9NlKPo9dih7NwqI3NucUvviBxpuTMS8a5Lp89eY5AMAwomPXMzF/5FuM/C2F
jDpYOmCCVsINeY8eA60ONKfigYYhy7UaYqkr3IoPYchYDvMVM/vaPt4dJIFwgOws
1ypvaZAjwSqLxxzpQIY56vQ3cToVueaK+DCXU9t4DbQaii11IqVy6HeONEYDETGs
Z6xBfE6athQnhyk1xAxcWmClKBGIuLyRh67+JAO/Ovq4OQxbCJ7l9jLC/6/dYXac
HMGqSK4bXHDiKgL8YLiUxc/UC0jSR58avTdLDJfqgJCAzcIIwGh4BxXCsvN9c1dM
3VWPQWuPrUCOzni/4XSh/K6ZvQzYKDovKhsv7N5qYubWVvDI4oVBOIjTyKb9vY63
wWspIfyHqwKTkk/3tiqaboASFvYqIaJQmoI3tspBRaX4jfE1IpVEQyDmxbLe18/d
HVhByImaQcFtNNwyxQPAOYotuohOLdCDUWIGMzTeutz6zQqe854Zx6Z3aj8DD02G
jCquWXMVFAKESdI/Txg72toL3Xg8RdfzuLaNsOG9vI7Omorl7+lJYO9ixJxBqpZ7
G6pEQXAhTLE35MDr7fZNpKGHIzk3Ya87MM2lKC8oqFovA4ymPz7KpcUlj3kKWtpy
qjnEEz32Pkj+hHzLndcDkxhBWXUzcph5JRZvtoHPOyXuIve0k/eP9exob+AImuCl
zLvIJ8KQjKwqt6SBrnB11zoaedRUQ0Qjvba5YInWEJ83/C+0dr5zzvmTEWnqjvxW
ZHms+u9AtkogMVQc+SVqxu6FhcXQxUWUbi7ruHRY+l8mOhGmAgPINodX4JbqhRSu
iJMEONJcRDqvhjwX9Qo7T7yztUdZMDIhHBaTEgjXLs+BG3pE/quOwV7ffwFeR1L4
cVh+oTMvafsGhzLLJXK/PlVMu9r9es6I5ZPcj2HFPpaD0Nf/DeG5yK0JXWQML+4t
8otIlNXirv3bzlhkQmHYbzDkG4rAZQElCD0vQTuyGG7MECcm2/yTii0Dv60x7yE1
jRXTDAw788cnsjeVW05kfhioDA6qICCw04PaiDaeE//X+aACcwh+F8Z4Sm9sywFp
hh3bzb/61xxhUrNHYamJIpSHx1Dom35EShw6f8r6PM4NTlg2XTFNGhAE2ILMUO5o
NmDyzqEhqQ5Plcol+BZKBTcjRyaslhKK1d/Uk1r0jKusgY+dD/v2LDcnl2mugvFB
lpe87ZiTWat4eMksfYh9BxQsr1/m+WAb/hSwGmeqCdfy/RwffuEyvzzOJz/mtZhI
AZkryzqbHtvEu2aFLMOObEKXq14xY8Ez3QLcsHMdBVwD1Sj+AbMaCfRcPNfWhmsV
lMT35k9qBns2JwL5ImaifnczkiRrsA5JLdvzsSX/TD0TVh82dpSXFq8uemprGWli
lxVhYDg5uV3ijm342xsHlqIJkBEN819mX1z+ZRKLXyxk1tsNx5aMNxaYuI+mtL+L
mCOPMvVzaiOvMhZQyaPjciU00pGIRasguffdGW9XiftfySfnYZsFZ3sCwBGfac9b
6SBaQa0VhjYfUsYNiQ3w79pZRohMfqJlBCUYDNbtAgGhlJDUfjlovseIGFzMHtXH
fvb9U+M2FaUQrEhKeU+GvLzD+GvfF9/jjSF+5ND+IWzKp+Ra6h9yCfNa+rPOmwh1
d/5Vm8Sf3gV3jnRmmcsnlHPsqBg+BSsESbaxQ7/o/AI6pOcxMc+hT3jsPk9riFMF
GSWK5KN9cwol6xptkOTBSY0v7ZFsSeYS7bmJewa08dPGlOJWrZ3Ijiy/XQ86Txi/
FnGwe53kLeuZJaDXKI4XaCfBLcUoGhYsVt0C8WSckO2h05GbK9AaUjn6jAW+rHB9
qkRt49L9jp21al0uoyOMbrw4H1PE3uOWnKSRe9YSaOJchxSBhQlHbR1PuaM/g9Cb
s0O6fqqidqnbIdqm5o2wYII6FoJtHKhcyltXJCOS/C18P/tPzGV4SPsECQCrtAJn
5mKwwmzrmQzTSygCNnAY8sKjl5nokio1I71uO7JZ0Z2oBa571gZkNThgXRKLCh+9
W02Orb7mvWb/khR6pSI/d5uIZ0cOqY0IyfwSRVaaPJm28wQTIjcT6LtaemjX8owy
E6NvYVf+lOgFbTjutT8i+FMQDocKOOYqH79x9P51N7Pf4R674AKL2DdzGqXCD8kX
GbUMVIYMth8WhNZ9JcCNuKkZH45H82Z+cxnM3UTC5aRWaGP3IAHt/wT2oZrlreuT
fzjaeKcEu82qVzznRC8xTmBlzt+Oq/Goi3NwXoM+B/2uTMSq/n4GzFUn7LE0lxxK
fmfMUHHZw+JLDisAD7zxKjvm0tV0K/m7z3sJYEcpejH+T7Olmuo/E8nvpLcsjAPk
JhUDb6bXdrSD9nBtTaUbfCeFhFSoJ3k/H/CqIjTJt2c3338ZUePX41TutdrOoIzF
p665vAL8f97a8+hW3P6nGKGQafixVFtKLS5B4QetRKin0gBap3DNMDguPWxqJ/yL
5kaXhJlF8c8Mx51zLcbYbi9RA9U+STJOWHgDGmTWPuabKC+j+G8FeucMymsJq2OY
vojpRHDq4bSQqiY0kovrAwWQDP2PmUr7rEW52aDa1vmfA2g3xw1tgbiVQlDfcdII
HIRjY0ZlcuIbieQnRIPbzxSduB2fIo5gegL5DyTlWiK0z6/L6QutXuHihSt0xfj5
5aV2dAXDGYeGE0pTEjOF1gQ/GaQRbkrjSnbOZHtAucncVa4Fy+T1HR/ovw8mYbPs
BY5VnYUGGe9shbaBZL/7dPssBH6JGmz6JktgaYr8AKB9eO39IWdw701JhPjYo3WK
pWlCd8XSjLLNXrUrk9FCGsHK9uwuKSnAikX0BMabfuej84n+k3XMr8jYRdG6cCvH
SPCPIkdMsjaajtvKTPJ5EEo+ErEbfpwqxmIxQXDQHD4007vtLi5pUQ59x4zx0oqE
gYJ4X8a/m/drY570YpPU1KOPM7C8EuOqiScoCFihFBsaEfzq6HmPIq+q65YPqfMt
trutG36Omn3pfqB26wvYdnEOdTs317KMRSizWlCb+bYEntC8GExHXg7a+4JIi4jI
X/yCB9Mnh0UfWJcgF3gWonjycixwftd+tjWF+Fhk2zqSQqsKczNk9PROPUIw1kBz
Ib5PiKOA8X2GqWwiJV6Ebi1sscWp1Dcehm2bJ5vLe/sN8qP/6mx0qDD6Ljr7FvqL
fUFcX/bwfPi+WeofCKsyooEY5+pr6DFAsVbNe+NOnAEjFuttyLqHReorWv4WhMJ3
jCpnPbU15IGNlhPf93teXEfr5Jke4hfuh1cEg32xmNXBQrQtEJ28Q58AHgHu/bi2
OPwiNhRxaExtd59rD0tSUVRzcVVvz/JBNlEa8HZdhUQstI4GX97kU4pWOLFM/pDu
GI1HW+mUJKMTNv4YK3BFa/db8LW0RZ67eW2DVPkKC7WfsV5Gj/DMDOEX2ev0CicE
Xjob4kxVp1gY9eV4EN/4qYfamOo35fFbSTXIY8WBL6vO9MICmA+KoMM+rDtrwVN/
TQfWkqiB3W5Rg59yVyH4jo8jTjHtFalNZivhKC2HPhZT6dvCN/oUSnAsLc4Q7NT/
cCxpLkgkj07ZpV8AFHNha8ZUnZMe9f4T7Z2/1fvrqU1I0jq+MFDquS8CZMq8Br1V
dGLRPuKqhiLPhbek0cKYZ8eP04rSv4lI0vzAxXDhJzrJrzcOYydZZXONMZq8+Xxx
6tT+bwjGSPOVWzIecyKOFT3wLT3BgOI+H52sEAowf+eRZWQtRiLLnfUKQ/1WHCfv
+xPo9D5lSkhhymTXmskSrPlKmmoyTwScuR0D6Z5utHcbU2W26IGvlBbP6DkGTmYC
mKstELhtV+m98x1PDFgWx3qX1vl4TmOhpdFZGp7M9mcOaU9V1ThTk+cl0uULFo8A
dOOM+IcUZUMq6me6Xmt9coNmcna8zKaQvepCd2u+iMv/4aZIc5De4xcp2dPEashm
PROXcThowE5pCgPL/jrhdT5LDrSRpWmKDDS07IFcgCipXiCaT7JjJyPzcOE32rDK
unbkidtS/IHC4uSw6m+PJiCk2OvUJp2S42rXaEAKOv5rURoK5PYLkEVLqv5OZHK0
ioEJpqWDvxJ/s/99UmSJdoxwNHc5TsmK1EMT6im8UKUQFJ7FRP2wRP9EOD7iUuJa
jWLUlg/gPx3OaiurfeI3IWnYtUaeWKjeGsQ5tq5yvNSaRQRUmRftwnQfG6spfT0R
4xFbgWFQeWpvzsVw6dojAF4/agzmkhDoGJ3iB8u18Ot8M3t0r+IK6XrJBd8WncXV
ineXj0/Hbd6U/RL5pfHQbAQai1OQztua6xAyZCnE5mPPIbd8SPA+l9PgLi/DiCc+
2ZK/D9EaqJu5nkv359As0M+U2XTW1/NDyIkgau0EVAX5aSIGFQixSXTfMgluphsn
WqFyXGmPRwT2OKp5/kcVsKg/lJjt4KPKHA9ezIP+3kCEN9QDQ09yKSpp1/lN4TaN
5rAlbfRqslt2AlbFgSLepoRkNcggS8AJDSWVcrSxVlJRGrQQ47XxZytnw347vZQE
qMJZ9M3h2ngQXZ+Qb5590w641nfXl6UUg2AgkTsPynSR91DTFQL/EXm3aIIM+1qa
FzY5VqooL/e6lGJcxyX9ZNqBbqfy1I+9p1ivFmGIvZSrxPAf2UbbC16R+uFLPVKr
XmXc2ntH+a0z4/KDObfCSjKEckBkumKIKcDjQElsYrtPI6ie+PgCcrI+gEGOJmSV
EJkQ4s+/1y8SsQ0SjT8cjzoGNYIiuRnhwnuMoWLePrZUUdyXY1J/h+CyFmOVpjnP
3KHhve8Vl0zElbC4HZZBJwSwxOWzuoU3TD42lYnpoEgbwGsTwkATRgPRXwT4kaO6
/t0BwnmUF9uV7tBvWJ3bSPMN45nKBaMWCBvfOBtmlcpnxGPfEWUCOMhSlQgg7qI8
lEmMj8sQwI0YTUedAxfeOE+BevR6Qyk5GXXFBBgLkyRF75AaxVLsWeeFIde6XQrH
JXSZ7OMDEmi4sFCc2kzgkRrXK1Wpb+bY704k4X2HXA67EW0ZZi/ERC7C3B6+X4Tp
Q/8LsgxpxxpykW/kroG54nLvtUmhYMzQRQw6K6gKzc2NoNEUewEzXCyvAUoekqz5
9TUWVsolpyXV65URB3Dn7JyqSvQEwZc86LTYD8a/uJvNaVaGB2QpQdrY0LWrgyGn
ScBiVrVvsWa27WQAzM2w2jI1H0EHECe+cp235gcleXO4tTv+xf4gAm3yZKay12xb
8lUuXm7Y7FHWSYpGph2ApYlNcnKklao1+p//fiANRq3XX4LS4luh5nxQIWC2DwzI
kXmF3tYqEZo2y/0xQJi4jHeBtxybk0iUmyAlFZd9VQThvsgAF9NY3B1C99WJXywC
nImOLxuBARS86iO6gbKHEpWHT6UugvhkltBHvVBfnUu5YGJ+a/k5IBIOibZPiA0A
EUzdvUmWTm87N+HnELMor3Xzv5lDGJEis2XV2SBH0mITdd94xVlGExvbOrEHj3Nn
36y1IO7HAAA9niBi6HYmoqYecU2VMrBgEou2r8mJy/t7GKgJA1jzbjJeuHqAM06/
iAbgs4XD3Kx9SE0z1eBY5QdeXR0gOnC/iv0ehWC62EfNuQbBWby/P+ZtweRjoOEm
T2tRBlAhL6x3D/saoNfDoNWbWI53lW10DW8X3J3p6Wc4nAj4z1u2nvaMQpYrUZAT
ct/A42rSZtzPus+po5cZaKbbPKM8MMHRl48MSNbHG/rZRtN/CKf8mQiEMnQoLGwP
fGamZpXGWKYpEhmJFNuQ8GLZUAUBsp0LM8EkxGd4bd8uUrLpTRLa9nPIUPKXARw/
zPamntPdgYstVDx34CLFAf1TpvEZkhKt8Y3CYhaWnFrfAkxSvXpy7av/sJFYlmEI
riUDz/KmfClJg+tz3D58DCdG9bV71ide0Dye8HoNRyTPN4OFHrdxyvehm5IuQtgj
stjExyb+enAJR3cqEZ5q6yuvgKHkd4xHyJgklhBuQRwZrdVNRJV+MkIm/Im7Rrad
e6MMtJ1VvFzZsTAtD59QjujfDlxmx7gV3BHUWhy1IVmVcYmLC1zUhmfLDFQMdzO/
aJ9XKu4do+y2gae//lSOcUn2da+ZmAXL1TFBxtj1hgIsLTqROnUpbKHf/pUVlIV3
bhML6jNbxvWTk1g0P/P+4OJTITpzr/LxxiwOBnmVPEVpgbrLYXK7WJYEgwNxXp3d
KxhESL8wa/3fTrDNGigOsURKJwnIysxglhhq5vwcSJysyMTimPcj1HVxXTr8TY64
saf0hTV+YHOtQIZwXOBCSpitgil8m1UnUZqTqgvIbeSjfvGyrWVLgLc8Z6Yf/Hft
P5Q65Tc1Bpio1YSsOYOvVn5lDxQqqQeBVf3NhALjwHMrS6+WHlIukiBfZDARXO5Q
i6QLIP2kW6vCWUL/FlZZsbIyyQfJkepsY91yzI2t5rJbo/EmvK4nZyjjvwtJXttt
ZCybmXkRpKjTdj4rmd/RwKny/+qtvhXkC7gGUrq3IVFMqm0woWd91Yf0mS73hRYw
UiJb9TItggzKaFJ+a7+KQvqOjpCuX7KUSGo/3EUqeAYnLxNBAjPlXdz4gAeXD7VV
ewAtvaTrpPdVs1+osydN1pkG55I4iUEmRgb/rb1al+H1gVOC4WnAynBzbrIIbCJI
3pp+w1Y84MSmN3AZT/DVoexFeFbY3sx72f1wrOnUO2xDQ8v0XeREFICZub8mgI0q
u8Ap1xBz3CTMglkZPYdz3A49MyJ2WixvXw2SKiK/e/aLz4uTmJz7trsfNUJIsmda
11ZF3E4ZdEeVLs9AqoYkBXceNqthRFnu5yWnkGe3+ybOXWW9ZXhdS0EhlB5UF3wR
8MoUTw5HvHc74EPEqG9snpy017Wx5Q7V3GQmZvzCx4K2JtKnPNoA7sac578cTLFp
ncttejcAXzsDf4xt3be7C8B+P+Tx59PcS3yA3zAntFUCV+SpM9qeyBCtFYxuLXrN
hvdDN3+Esf4UQKoJjGuySsmzi84rMLFi92RfMRKo2FKDmGvn9mk6lOd+1iswkDDQ
oKyxFZZN96qu5+HkZY+nTH+htSTFD60mk4hm7LM4rwXWtgH639m4ImYkCHPrxljR
+3IrjbXA5jfEx/elC2OL1y5utt1DSq+YVBaOCyRiiadT4PyC2KApGsZLhh8o94vP
fmByGQ6UCybFo4mR9zi6mD6yW6Sgp7ex4vlqJjR0TkCS6JoV1Hctucfb/AG6+O6U
YT0UcHmlzjZlS4NiUcKaBVlr+BYYeSQYAHi5tpQ2kglgrw66B2H4tLDIVpU0Ly5I
nvzI3Ktsg7HTlSnaR77xaUuAOk3d9mpKHSWp3wtFkRWQbu7I7kmow4pTkG4uYhYX
/RnEjnbNSmJYuUJK3e0eJasBBktrr+cGKb9J5EEwvQBWDHtI0TIEhwmCx17vIFjt
FbagOolzW+igja/mk4m2VI7ke7eH1nE7Vw58rB7WjngkmvTbXktKrPzgfkMbdshU
k4MH9SNPGaHvlJT6tAkGwZLwGY1abluFw2gTFs4nX0UTxqo+bpLGyw/xt7jE5cna
rwZr2ZFyQwEvSapyeiA96WV7Yix/O2p5I4QThugm7DNkIoM0VMjMUu+yAZCmB5nk
UvmlT9dOroZM2zexC2cH5y7CeMpIK4dpgq2NatkSE4NPw1P5vXV0UyT34BWtdd6W
O3BDZ7jIlmY+aOiyeiH/OMY+btQo+Wg3VQrfkEbNBCJdVbGq5ObXMSKXgQZRqZwK
vuHrvp+p4lyZWTmKDSs+SEH5Yv+p74rxod6/nX6xJO/g3aaH+NDYPkf8q3iR4ose
zhVPl9lpG7XgLY97sNPJbVW06Pa3hYGQwSAqBLEDwIxRoJjg3XlhkG3B5VFXETYp
5ddTCplrlL5CEZrT8HWPXe/J87pimQ/Wp8U0T28eVrawolO3YLYNrzwOJ9GuRm5B
PreuQVdKmRD98eSqrHcDKoVjNZj3gAD1wA/md+4BoqFD7M/mK6pRKn+kCAYcvhxL
xhiEPmL/+9e8RpPVPEjZs3TyusOEpA/G8leeSNPJEHOg+hoRFks2Ua90Xd51fRDt
vNCXGlwl0Izau935zsCPa1GZTBzfwzN4nq/ledTpXCRBEFdBX+lHojaFccsYsozg
NPLR+AAVBvy4zIv8IIsjCmInd2s4igPXeNfIhIqBRb/ck2Gt2hMQFBAOHk20nPw6
rKcVfOmFU30axihUXQyqoABP7kMMlAq4Xqs7ueI8L7ErBVqXBfQcclIELHuP/ONM
7Zn5hxb5NBnIFguf+XidLMPopwb7LeR5cpV04cQwDdVGDhDSYfKmg/kGVGDT11W6
IZzQIAu/WMkSyJ6Ko+dNswLqaYaswzfq4UamuYn7yb3BueUFkf4rFk8BLlpauwqX
fk7+tVIrRCAJN5/GdgT8NZlOzRpiYk4kUakWWRdgcrmhuJgdr48LZc6xlH+VSZla
angY84K+YeKxAwcahDtl3ZQkRKn0ANh0NqCfd/7fosTqBdQ3YGJUP8/T8uyqwqky
1ae5ntKK07upLV6H0n+k3JVjRYoWe2n3RexkMFZUSMMh/EziN5XUbTVNyejO1uTL
nclVbktb788/bDOgSubDRBN2YEVmHwhFZcVvAwnFD2JEAih92h5Sg7NhtLiIxYr+
1RJluW/4uDpXZPNc4nkBilXJWJRK0oaEDonT2Qgy7+5k7z8xqkaouISlITaukDWU
P6iMG7doEL1tvbK2AhoAVFG63LVX6f5XHRo/57u5Cj/O+cA9uj4tv9MtXWQhGDyB
JnzROOjYtiErRfenZuWBZRcyvdaNB4wOLprNjm6njAkKoVECTTn0t3M5K2trA9On
5FeUuS27oqgdl8ZntPz79ox/XMMJLwDoUtgXARQckBJDxM+PN8Z+CjmFwDtxqBKa
MmU3xsOQ4sf3IhND9WZ5Jo5VA6hRb+fwEXxQCvWTJ2cSFMl03dM677GNtOnS4rRG
1W8YXyG+omrZw/I/nAdkgQXeeuEwIRGULa5XQIJv0CUKH3iZXgRLo9346JMRz/jq
FsQyzM97QyaBTlG4DX4ZkAfyNCZczLuhAGOMpX0xTc56nqDgIq4oUq0hJhbx1PtI
Ft5adVBlMboUQQUDND0esNxQiDnHVmHiGzGkFKzWFtFVuVyIvQ3sJEnzXstINAuk
vNR6blbry8eSfWE+CD+XjLRdWCxqxV4YxhlijYoo10+oA5di2A0w37tYUGD5MtBo
ZinllFC2MCKo9tYm6mrtu1BVdi2GN0MkrFF8QSLv6jADusYqFiAWIwB130Ojlw+f
rj8dCz7RezdDfo8Z6rOrXxf0G0xvhKtnL5uMjEIDyrhXmhlW20gMh/YadISxYZMo
Tq2W0NUJfXSH3+byWI9dUkMx9aOgBmdUljVDomFVMXhy3mgvRk1OCB3+llAyLrJu
fkxYFKh4kU7eYtgQLmyDGni9HJiEgQqWe4XF+8OrD+t44KgZpLDwlsFqJ9AyOJrm
6cBfeHIEpsWYs0aYoQdWfM+FjDQk6h0/dcT9FTURNZ6ArSer+JeEfvaDJ0Oifz9b
9g1bscvpGCXj7O9u0x7OzRjOA4MAzqLq+uVQVRk8FgKLq6lZ2rRJOrbqHiwhf1HJ
9C1sFeSanFCGrb6T4EXnpXZzz0wDuts1ArzQuZXFalHwBGIdA/YV6TX9NVeR7dS4
b6jl6NPd7b3UdgYmPoGuHBspdCm7XbKu9kx1d3OXdKKSQN/ogp4Jk3GYKOcLzqmi
EpzIeVF/DFd/cCOI1mLEGmfrDEy3Jjh3tu90VrK2NFk8L2M62gG5aDKdFGYdmZ3F
BeJa6ikQLMkqoTh5YxoM9r3VI9pX3UfR80ebKiY+kz+9csocKIAGh9/JZ4+pywV4
+xXDSdW724yeghqJgSFw48oaxEwKv0ku+4hMzDN2+Tbep/yP1pxDbLnA26xqDFeX
ueqrZN5PI98Ggm0mQzmOydTp4p9UzJxiq2LEnreDfleg4hrbwaaR5YOkQbodNWJU
NDE9lU7iw2O8Z9M6VqThvrBxOwo3KrmqM1o13KbshLn8TxAOwCkgcFatoJEXHLdG
G+c2yK7SPB7e0S/lrWaLNg9Ic1Pm0IB0cJGd7EC1MFoBxqzMpp2QF/luH5e+XjhL
AFVVtC42TDqgB70saGtxsIoW6dBQaVrGJSdB+3ysaX0xSXnYO49UDw3vMf0jhZYd
vLv1uMh11Paowiba9wS6pTTjmY4JcfkpvNdgqgcq873heXVfHG+c23t6G7FtycJ7
91xgmbSnLYxS9j9NydmBTvPpfH5TFAXIdeKwULOk7Hz2TZCduCVHPnRtxkhIkx30
JFe2Cph6SrRYs4C1rwHH9eHlc/khXvR+Q/ZMzqTNo/wazSsq6/UGhPmQ/g7KMUgL
4Z+IoTEOESVWRO+HQjeRZfYKJ/KLbMDxTixGhqQoKN/06LUmDy9N1h7dBvY/d1BA
Gr53s0mFR25QejKXwkEHNFQ+eTUfIytyb2gr6lqfxe1FENkOJn2xbSPvL/jJ0i9f
uTF/KKfjRgqfdy6dwTW5y3fyr6/Y1hLVg9/UIr0LB40K0LGi6j7OaP4ipw+vYACu
HHeZ7rzcOsO30nrbncZFVhJPVPyCu+kEm+R59vnG4Bykmu1KVMZ2uAGkYIkJT1G/
Aw8iaNBziZeB7cK1ao79Unu14O7XrN/LKSEoOEwkW72VGDf79KfX3qHY14Mfbd4y
eLEcoSkjwYOfvRdam0Oc6bNsBGCzqSp/NJybZTVl0+UyHSPb3d5vV5goD4e2ZH7P
tUc3QwJZBfXKKuFViQ58e5u/kFDTuEV0v1lJafDm7+5cO3HPyMSezRsjf4JhDQem
Huy8Mj2oqrKcvu2o8ADM+toX9UnR4da7bOZBazjyUd5zcFVbL6sn37rXRqDqZ4Tc
CQ+1459mMtg667HSJ6t1Q1Fm/woyWzZgCMEhOOVfVKXpRYMSB4HaF7JSSlJ7JX+m
ysUh3BDpPkia5o7Svz8zTeL1iG5TvW6woIIg9YZPs676g5ivxswAfWFmrwa1vf0L
azs+VaWhY7925IcM9LkqX/Fgs26p6H9Sw10u2WpgjzolRQtAGF8vKq5xayhbBAK7
693nKDT7jBXQIG3SZk/eE552Uq2UOEfrZr1xFWrwzou4AG1Ko7uuYPAtFVaQD9Hj
bF/eU5xl1ImQcVbiAuzP3Coorahu8lPdv6T+i9TYbdYDyFUMZTXqpFKtg+LJ+sIf
6oGNOsef785Rfl3+ywSVrmKRzB9LX6CGXuMVy87433usY4wEFgQSYlrhA1Rp/tqC
gWNhBq85TpWZRa+s8XZJItfuigOEswjW449bOwWsMUEysRH0apOF2dVXPMDlzxTr
fy8XKs4+sT/9xUuWR+JdMiK5OBLu/yuDKixA81z1BV//fGxklB4fthmwojhF6m0f
hVT3t8ETrOL+1vhbdbQGbW98VQckLT+iEccqcja59Bi4txODIP0GGxZStTRVN7gO
Vze9M2D8TzvuRIGHHOqR92jCzhg/pDLnywyGm4I+CDAGyRvRACRsFEMu2BV401by
av+KKfmrhXz4I16+0IEXmdAmJjOjT8B/yESZKr1Y47N0kcbXQwe4GkjwW4myicRH
M2tZ9FAxP7+41uj19/kKEN3Wc7JGl58ZT3W55iDYX0xYiZImD9Jypz+ABFgoX50F
W3W+FlKWFvEHKsDLE8U9v99JJwDRwtNNzBncYJwNzhIB/r0YNoOxnsgrmb1WH99I
0pXdczEk8X9YdnMwy3UmhP8IN21d7/Erv+eVMuzXf3BDeLNFVk+H22MujRcHqaz3
wsK+rb5XXRct62q/j5b0u6Ylu8mPEoz+HkTtw2lETYOPmANxUmNE6//8uQ+VRHQw
0lwQYM912UuPhfQ+lmu+U/vNnuTBhmXZfsnMnVEPeye0VvhynNqqi2ZZrI5o9FfG
AZUOhCtqRNrMsGNXZqIQceKH5tVdpQUO1ss4RRsazhpCAN9SK49c0wK4ru8b4xyj
vluJQYbfBEEsHX7v4I7YCGp7jY6vHGvsgoQxqPycP/yCticWpYbIsXYcu0kP34PC
icDBxl2RUegBfA6pGZOWVqS5Gc4MxCIU0u9dCNCLxl+8L54y54VvUWu/7+mHl/k7
9YL79yaMjdAPcu9hkQuSIXM/bbdv53lL18CRzNP29m+jIg7J8uEeA8QC7Zv6PTPR
jLqmbVVT+a5gh9AOcI90GnaR7VFUAu2YEzwVIFEX8AGqbloQ/5VWj48pKtzcMUQ5
Z8POlCSTxFUBIt9RKk7rf0ipLJ5Q377x6LsFowWojlyNVz5YhmiBBClnGNprDslN
T7t+OgJitsoZnZUr4DdsriPytKTnM7me74SMokdkpch8YT4bnvDiH0MCTPATF6tm
ULF9cBtuG4k9VFv6JPMyeF3K3ouNTk5IvfvHEsbwmy5b6X9YmOgtbSXMMcLFJdGn
QZ70U3bK3ZTL7lux89RwVtdy/eXTq8icXXduqBWK4T6+Lqj3YUg/tM8Cfqdynotk
ND/y2V2soVkLpWnqEBzl5JcC9NFQLA9dU250VFzZRgby4y5kbuXVxtGIpqEZGvHp
P5pjdqXo/ufyfDmL8Ij3IO/6llc0O6sZMMWmMzbsYzJAPBapVdicsCZCZn8V3AjO
TEzlYHdQ46s+NJGwCf6RXGG4eDTZbQ39MRY2d0YSIAduxH87Q2pkyTk8SMXj03SU
hsCq70Vy4MWsvflSpr37UufQ7nKyt8y9cI5xRfDQtVow1wBxh615i9vlLsrl6tLS
0lx3iKDfhbvaFKOUTiy4IBufHzqnjj7VfnAowM7acbpy5MOF78fy61UYQJkhLJwI
sZnUenmQ8RqKOzmj0Uyqjsknd2cvEFn7/+6OTIkGGgZ8dYgLfyAFayM9s0pnbpPX
zuIiXZ+Zr5fYeLLsaDxnDKEKn4rkN2jK8UffJwsVu7D5eSHfJkZ/UC5sHMa2+00I
xO8SBGqS8K7xygwvCkBvfLlcY5PMZ4x+pKcgQImtryHs5e8lqwky/ojaEjzNpd1J
FQctrTKVfOp12UXxbAZVwBIj34qKFUou9giifjiPBymlDpCEeZBTucCZNnGMl4XC
yIS1kS1kuxbKTP9WnW4mSvXh20xkq5AXWQcYn9K8NPAtXC45vTSh2KHSL2J2Rewa
v+U9Uqd0BVEP/Jw7pTqqVknpLpkb19JJTaywuxUrijJ5lL/hU6ya6no6IUyiejSC
qd6uxEv0zIVahqtvFN9Mc6K4017IPdxt2kDJAvDBOT9aYHwvfYmqpY4wElXde/WQ
CEdZ6O1lc6nvDS11Lv6G2umryhFpHy6YT0hI1N+agblf6LWgdodSdQWMSQH5ELgU
dbIH4ojEIAeB40Kd6RzHZYse6uxU0NCo8rUynJTCyaSVgLn06CdhQ4ZOZXyJb+VO
+ctg84E2yNhZEZtdA/d2f3/IPHyYVkMnx6lu99tInNpPqSv1H7O9rskrWjxnLb8W
qL0eIkYq7inJId3HMgadFuHm714EdoOVDtvHRQvWdxGlsZPHxNfbaABN1h8M8WPw
p/YNmCPNHAu12c5Lx4JfoqmrontfwjtHh2gQ4mvO7/Tzk+5LJrPZZ/7DasO6Qo80
Bnf6wc1X+yrd9s/s8Zh03XdHZ5LZZrBu+K2Y3lIaR3Xh4gyYPvhjHHv7eFIKUGgf
UkjA/bnTj9HprR8uQl6aw5xVJzOfrpQvRFS35xVEPcA/oq7HuGIFZro7ptaxCvOW
c9aDmBRmxVBuBQkFkrGMoE2NGDw6ru2MGKs7Ay7zbKKAed99P1Rk1Z92GW8kCdOQ
o9OHKMKK0ywge0kW/7bDstIx9A/Umryor/JtapniifqHZ+MlAvkQweZiwHP8eH1T
KxlKA6KnxNE0eW0nbtD4tMDFQOGQ8wfg5WlQOy1zCyg21qXWOZITVGVVD/5tO1LG
UkR1oXJaFlGGhk02wcNzJX72m+PnfJzoOhzu13fK92/r0tKJeN9yQGkQgsG5dMaz
pvU9Uc9NFc7Jka8IhgBUPidUuRSYtn+MXz80A91Fg7kjLUnMv7hFgUC1DYN7eMkI
S01iMgDfzhCyjllAqJ0olL2g72p8JdQXu3gJDlUvm3klmCbcRFPAO7Ue6dB7NS2W
YkAv+aHw1KnlQKn5xTLWzGp9sebTS2UNZEG8Dl4u7xE1nk2y95hIcndr2+ssgizO
Hj3FSpnezUBA5W1hsvYYGAMUHSZlzYL4t1TZIiWxx/QYoJq+V2zroyY6QtiXPAZD
ChkyMKuIIMEzkTQmjBdfmqIhEQD1qLNRks3bPvhyrGeIWrBOo9EuOkSDUSezFmTf
IAvSymVIQbKvbYZjON7nXHE2GjBarSweo1B4mYV4Ds0LrTEuQfnQm9kamULeg72z
FoDvn26HYy5MUwM3hURudqkVPrPVmya0f5NrKoGeOtik9SYbr/dXUFtTNJfFDXzu
ZQsaBLx5wEjAaTak1Xtyz7K8ZlcmqtKWCFDtjXg0TgCuWVOQOFvmm6usXG2kVWfj
ClcVhFgVoHb4w9y9J59fHqZCw8+KYRKcQGslXjgB1AVLQSZtxCQ8re4NuzfjGluy
2iLIagWlW87XLHBl5lgd0H/yztXG6kznNXzDho+SdFfdGUGpmhHQd8PW8UzVSczA
Bk0b96So4nx00NcXsjh6M/RohAp/G0VgKjJZ8sfmYUqI/wDk63CPxwK9ZSjJervE
FguHjHez4Q5ZgFVTCpy9Er8ay2RMDihQICQ6k8G+i+wX2cFCDc8YMPhKR/CH+K5k
glnd9ezuqXwSqRWpZzTVfMasns9KxTxL1Xm1fsupiNTJGZt3su0bHwjdL9uqH/58
nXa2e5T5PJAL1IIHGj9CEkfC6iiYP/QpOJUX1QTxbnD4+UWgl8+G+GNTheF/rMWC
4abeJ2mX+SLdk/1uVqqNgGWkvCirlBHii8lPqyfasKOIpRK2NDjOmzx1y9RvWn+x
27iMC0XyUgycEKX+J7S2ZO7wPEnJeCzCv+mJEv/Rd+qFywGTbgaISGhwdcjs1/VW
qpj3SZiBfUt/xgml86uSX83we6JnmhkdgC1Fmoj3Q+B5wEVX/D9bHhRnzWqN3bWX
WUD/YPxcsHPBqR8CE2pLI/hNnsoCwtOXCsy2/diEkV+sBknY8Oq46rEV6Wq6mj/6
lmiQ5949G44s6krLDqP/y8WM2hSkKUEQeLndoYRTGOmgVIaYgquG8jug9abrZxaC
+6MHNK03ZmoxlTB7CiDbZ4N86w/wc66hPNLwmhm3/P2hjnguy+M20GLudcpiSS3k
fmDk08biajSxONlagCF9rfPulba4v7UFIfJY4TiKPYM8SGKoAzGtlBtcA0rc+DmL
SydAkxVTBK5YhbW1ambNH57rZDZ2oy6Lh9F2GSL/zRODom3dssi964W+aF6p23sj
n0S+cB6V72dXSZbPi/b+waBQrcdIW0UkCa7mXicvwmc4DPaw3dxVRQYOTZDscoow
LdrZLblyGd6uRb0D8i6sBWpPu27ZeX6v4sVsX4+VfmGjTn5fm4OONPcG46ZIY1kR
25yOtWeqrO/b0XQ0I8OGhxCvFNw8MyI+eu9cWL0vIqRYB2D8aggeotJ0yAXCHnxP
luRbKS91LRgvgBSVVwh91kzdhM4OLGCRWAMmFae53sgjptFeAFhbOWQxAt1UmyCx
XHZ4Alp8vHpIDsCtmV2tdEJpwYepGE9p42pLdgxYwjVUItlMtoHeX4Pg7H3pxOCW
8QbEhsemxCdRs5G2OvfXpsRGfN2vT4BDob5uGWIghYTHdra+atahE23V/SeUOTLm
3eYc4MjdP6fZv0pcqFAR/iZEBjcJxoB9uJ3qXDH9tCYmnvYL34iSREVVTM0rTUkg
5TgwWMRcFQY9sZpBwHqjSW0NJDGZaL5Yfq/2eVy5ziUgK5lcp/suPz5jKHS6ElIU
xKmy8LDXiglKI5boBVGkCtHN5lgVqoHi8Khx2iXbL6XqrKzDwx+u+2E6qf/INtMO
cWhLmxhqCk5Fc7ly+2VKccfnemB6r9qbcBcK3chO3K8/zKmlbCjvrHpg8zW1iamO
5z9mOTgGyXuqZvryanhLTyDS+PRMZ9jLDe00kOgo3apMCvhRCJXNTU8Dg51TyCfA
sN407gNLshGiw+5QJCymoCBt0P1ynqCge2uXpiM3F+v+e5cGRpFQkvzMPzw+yGBj
5dkrMaHu/QZS/oqSoD3v+qr6sDLTqnJ75sBDXL2ywrxqx0Ft3Khgz8ccCzsHekJL
Bn8DMAtzL63nbw8A4wQR6YpOY5R2kFXmhaRggpoS/jjU8DahZY3Ad3RC6uX5ieAT
48j3DNadOCxw8FOsXsLNxIpce/FG20oTYrSi1581fUeaebl5hPGsBcyn8wExJ/oU
VXjlB6cquJIVlmE/5Cvr/NKMasnFstwtc9sASPx+UXA5bCyyb8Zxa6GGCbTW+Zyw
Wn+OlKUPSXgGW48u6hlCYpNqjMt0+PthaquJLov7VXNF1+i/syWRpbPCwyQ8Jup6
uesJ09VC5zww5pgxjeM0lWv+XGjYKavnjDBaQOy0YOuiDyAApGhTnM7yN4zZRRkk
oTwAkpEzr9Uh1YkAqjpwBAjASRlHyHDvonSjCx7u/c2aefehAd+yVrGb54rJaEsc
fUviVflxYbYIAgG+5/iwmLNO5CZ+V+xNKOY6L/ZbKRBGHeSqBB6M1i1qM/iczKV3
SPAKr/zU3ikkO1MLHhNxnuXmJaxUcjElMnjmwmWoN+DA501p2nVjOi0j1+KynYPf
irCVOdxxh9/v9TPQWtQigpPCCsaK62fip5KcN6ov3hKEAcnMd0xxK9ITD6sPhmNb
vMb+BcKB7oJLdfwFX7W5wlZ+udanp+234fBfPpWEqG2ANiHvJzzDWuruM6vjQCfF
pb5yz1dOv48JqqBZtj2WCG1kCLyqODG/i6UtcAdqfd8pKPzLxACME3TJnhMO2YNp
z9NpnXwWnxD/vuxp73H0/gkPuHD4X7bg0u/MlHo0kUH6h+y4IViBhDwc/CvmWQIe
iWfRN8l6xQiw/8LxuvBmFvIgx2AMSwV/qDLrz3tov29nfm+fVHNxn+pJQV34kD/e
foYfA42n2VIIMv6A1KbQ8RSoZsh9kcgxcsCcjt4QRGSRgczHje6S4iAP+YIgqPm5
Z7oU3Gu4nUcJIkHy/MFHBUJQCz0S+BVAulwq4cB49scefXlyZD8wHcggR2urN8l5
o8pwJ49AkYi9in5+XdjgSeJtNIqa+0+uKgVlD4LReu7HNbFIRqbRw++EOos9aHqF
Z/TikNYSk9Kn1QC7nINR+UvlGNHeC4wp7TIVz9l7DFHo2Tn4lWFjDTzKyluQ8VVH
moDXpNuuoBA3Cg8QnscxurBfjyQ0AIOXv4tfJko3aMKU98EPgjltXL4hlZXLb5Fm
wKEE/bVXi1nm9o5a5eDREY9TgFWkENL/c7vbtqUt+0bvfK1jN8Dl0FGDSBuuk8/R
hIQ+SBwcwUaqyYlKYElaEFitp5wDbjCNn5PjjnqywteTFJ0jA+eFzawXluSW3eGA
M6G5xo6bEz+/Y2NZSOOzaN6pKiC8lHMnrKQ378DlLzkmAHNoRlU2qs32z25Ej2w2
0J8maDDO23Rr/m1zX105F7XEw6Lo/2brWxINeoBb+ijmsxoulEblh1jNJ0CduRHh
57qVW0KqLxNO3WKHdMNjTeq6sqSnumlc56/GAkrgq9ywaUCi8TetvfVH9/aU/Lz1
B7qqXX092gYdOE1YSgF6HAQfQnezCKPvXR7/cEpjRNuWU4ZtPMbatDNZ1JbtnqGk
ILQwIU+4vBuhCt/ZGdqGPRxbZlg8cx33obhB1Q6TkDoO5R218g2we+l1Ix/SAucw
rCy7Ei6un46s/Zb/hfBuxVkkzYstuGEta7FmwZuKoIf6tA4+Vb4ze6SJuD/7kCfT
p5VCrowzuld3daIpr8qh3AzBlW0EqMUOB9XycQs2cBcRW34hzf6WFWjkmy1d1F8j
klIRMFPwSikyxCGr94yRDwCM61ggyWylGiVbgQQnTRY0fDS0jvj3ZoRtawXKcoVZ
qcQedp+AFdzCiJE5vSDSJd2r265eOjdNu3W9TfsQkUNYYH5shyq2U+s5onndga0U
EEvLWITwYarD/SB1vdsoTWwiL9CfJfN9f81NIFbJBAg7rJdhJuIeQzHXf2utLSln
RiAamX0Vrv3qR7coEvvx0GzByJ+0ZnOLixljjLz2FfczdUNCcAPHZXydZk06Ro4y
Eyn1c17BwXc8/b2sXB9JwneEpXzVq21B3ExAKw6ezy6G9CpEtAJI5rweTAUASfgo
nxPNnr02yUrQpmhbMD3YuBPaFGIDDyBb6BWcSeoFwgX3N7zISnGKuPIjy3+UKgSA
bQ7nBO7qKBL14xaOtbHr2sMq26yRoQdCfBbnIHBx1uyc6E9Cnw31NhgEDQrOsx8w
pahf/h3xS6ZQTwojyO57dVp4finoPNu+aTVyPc3M0Gb7BcNVdHtUO8mHTvgzyDML
gq+We7/cTIZC1tCRbDzv8Pu+cKcLL6ynjKAZuIvjMdtDI+CgSomqNXt/GZTDPniz
CnOTXNXpIETzAW2TigbdOty7ifPSu2IXJdQ8Uoi1IiDUUlo2yPX2csaXKwFUlX41
CYekmRMSYg66tY15ACQUazjzIM6OTqZiVd8nrjwlXQ6VBpeWbrbZyKLANoaWAffl
B1zyfnzKC8ErXT/UZJsxFsPO40XJCabqt9lVO+Zir6Oxc0RPwwhVHiiYDbRXzN3D
hVyP7fSRj9BkSQ+71kB0EfSXFbs638ELLxvM+pPsNa29UnlSDyhzhtBzu9nPUIe/
IzFfv8VUzT26uPGGkpViAQ0RESGNlr2gbGRuDV60jW++gqWvU8c6ZZh0VfUfMHpP
mR1qlyrlisB4po34OP/C3vX0Da2QWk4gIRi/CToJoOgNSn/Ee37wJ22AvUkzWGdp
muYEktS/SY8aWSJV9TzhuIaa8XrDyJ2PXUMNKAHK1NZJpKOezYgAFFA+hG4tPXR/
iqcGNVBgwWad2olz+gG/ValQR7uCeJerH8z+xy3c8B9AJagHlcnaKvZxmsEp7I2L
8l0Ho6EAmGGIBgx12I6UeLjdKPLhGKmBOVS4BEK+am32B3fCPclAYQXSyjRFFWRG
DBeODgp+QbVFgGWo41Hbp43fNGOcDUIvCLhjZeBxcE5tu1nXZWONWPIxqtmvGY6+
1uDrAcvpBxJKtvvffGH5wwxKFAZ/97i2Ku8YJbgpoXwqVZnYe9wFFCR6Gyh1ap2z
caGWZcXrRPnSQ3rJ2RVQfMutIChH3vpjtmEjZRrD+e2Qfe1/17FVb29N0t0tpQM3
k26sNChuELwei2FPyMlEQkSXkBVuFTy5w6Vc18z8XSOyNM3dj81gmLv9xNn8mPqP
Y843lrgvYviNnZgUela7zl+Z+2ibA2sDd0ZT4wJI8ud9ew28l3JyZyCkIYmmEc5u
toZsVxwAbo6o+5t2NuMvbP90XqmjWiW+kKLZ4S40KWcirvNyXn+Swe5kweFHz/TI
lQ+SyTp/2k+zo/nWaoeZZo7XWEcXCoSQGOEwjMj41gKFwHDd9jqLJKrPokfqHzYk
fwrtF8lYbkbUPYEv5JRvsW0c+ZuCU10NxgxQfVjqhwek21VfxID+WlznLBstVwuL
vZw0j2UObttOID337kPIkn7BxPUZaqS82U12rGDd2ApZzOTkiqqyBMKIyeto8YKv
FOAwe7u5Yc/AJ2XIPy645xIKCkYEXm9Vkx1d2is4MzCpx+5InJSbNIsR45TAfi8b
F/G/zKzJlsXYUdykZIGaQMPqSd2hK0N4+MqY65i78mu38oA4yJC3JmV2pP4KTk1R
YKro5+qGqUjdFtYF9TOYoN791w+opfNXh6x6WfTJGadAr2up1l1COFmk1fyTb9+U
gPG/lwhncnmIYO0oRn8fWS89P2crwlP66JHwW8PA1vL/rJHyEIYpJbz7rhni3QKj
6dKh3pJ3OczhJ8GOW1N5L5hj5KsIBr6kK4stQLSHwVLr8/fLVWbuc0PBry8Lz13Z
HvuYw0jDDpSA9s8fFfvGWhxifpQDMFHvCqkeBGIeDp7CIey08FysydEfQMCK5CgM
k842Quh/wgxt8Et9e3j66KozgfhOltOA7Vn4XQtIOy7Og9jW/8IRHtaT5mH52EjV
JPvGgc5SbXMqHZPrSzJVgNy5rzctjmLGhCjPCGEfL+kSOFHHJePgkZr15o84DR0E
2O0EYOt2kC4zWBb/NJ/1JBOQnpQCfSo3N6WwS8aVaewhlFsy2B1TqdDuYQhxZ2xk
WvgSGa5I8AopDcgPHbvoBnV2IHu8s84e4dOeUqPP5vLtcffSilXzVp8n+0RE2I9e
9JyQPyzuUEOzsvM8VvFIytG/fLShp2ROff5XJYgB+t3cAq5x0NL66Rtz9vAmaQA/
sqPeIrUj7sLGeTgiXw+syD2ECbuvV2CiXAJyZiJM+tZB7H6FSK+W7nadknoQn4uF
XZDIFV+3NtiOICPsOghAL8JQ9YTXoA0bkjMM7WmdYnMSuGJA3nWJTOlj+PB8y9w2
2snYOZ6cHccs4QGdRv3SPudNiQw9FRzJir9X54MGPzp49lBnp+c9ECrfByG9QsSJ
6aLAy5c0Ze6CKzNAP/fot/bFOYqNZscCicP4bTZiwJn2RyGWF4uZzd3yZayRhntN
7AEx0t4gFIEfGmdBAapU28Yajr2lx1/sOTi6H7ZJ2hCnP8oqitFwtKvE9ZuYyRnh
eJ/0lMrZr9Bz/5qqMGEzsWsTr20ecPCfVZjBSATpr80E0p7WLJFrnkdQXwWDxAsK
szaR31cRPdg9r58LtaFJhZUDxjqqyhovxHQDRnMXrAHkfw9BSPG2iRfdHLgOkxbb
1ywgUI4eZcyUoOHE+pcQNk23TTLl0Wo6l3whFfwCzjE2kvXnzEWQD10gR0cE9234
1E6eIlB7CfJ8mS1DwD4MNANgYbximPJPo1v61RHNDoAoZRGPJ8Htt9Ej9UsPkPAO
tnXsvbAe92mqbZYJ1DyibdiPlGxxVA74VTzffZywErczSOFYDoWQyx4TRzywVl/9
0mzStqYzRQx7SLdG064pvtwz228zZAZHT9c2Sb6P3SOz5k2WIro5B5OTet+mrRsC
2M+gxlsOqcxJxN7ftpT0hFD3H+4fTVpg/2ctGIntQTnu2V30lCq4aL7cbtRVjPUx
3oLtrWUW4ZooeP5eREFOWyC6sE8fVxM5DjxS1Yh5WQMWPbXtFaEnVO4wSWjgO9I+
BBW59NVrn9RnHa6qb8Sz5KuNUblufJAFC/jwviUjsHgFmgvHRy74wtkqxFT9a3Q+
swFG+BR32cKqTQxQ6sC6VOO4FDfHV60utH2LrNeftbhQt8PZ8rpK4CmsDEceS7cf
LDwy4mexlPkf/IWJCFeLL9fmDNv48dxQYYvTc4bse4eNqZiAuEPjpoGSjUmE3lm0
ruHlyuSLj2XE0p/8EFX5ndmQ6wukI/YXzhDYXxDG0rYCBOjEKJ+xfMBtRxW+hbgz
0x3Kzi/Gi/NsdYb5TQYsNsXP5UH9AnBnlDIX55YMSmtFae6ubxCsT1flH/UKF6g6
C170mR7zm3qnXTkRWvRoPysRVAlPhelHM2Swe8ppUmW8cE8RRN/EqBZZB4YE57SX
8kpt6h9QWksFqO7NJ6CZ7fOgaNwqZ3scByV7kjh3xbpcsERyipfPkNi0IuTPCBmY
Qa9hZ2lUmxUcKSCf6usAbTGcKMvQNGkYwEI8KWBAIs7pnC7tt0NXfJ4xWFyGJkbE
eQ3PTs/H7oc2e+00esVjohgj0o1e2Up8NKSCPGzSz/LQaNCokd7WMk92QzJ/9TXq
U+oq0T+PPpiZjO71YnK+IsqOHPRkyIq0qo5vL9diHHwFZnHjA57M92HuYuGzryxd
/5odWJv/Dk/ij8zQwAK9yX5F7aXxd+cNsm8VxzI51HWrxpTsLVZAzU/I5QZuX1t4
YJVpVOZebwggkmnR59rBu008ckWn/FPyeLk5NG5HCaXi6M4feepkJDyT6PqTy1ot
oyAi0IiBvfCDgeaicF0KozxsdWEzVLIAgbsCybpKclhiYuEnwVyoX2USKAs+r6fA
th2J+6lcHnKEIHBwC8dQV9Y8WoqB9gFX1EP3TWo8ecB4tUoeKiNOnaA65ML0Xc+c
v3k2juOXwdABMNhBSD9GcHfl4dXQKU7DFgf83tv9KdWRBCccU/UHxnFlG0PCqSF3
JIkhq3fGcOZdQK/crSzZypZUee85Xksqd22vD5K6W/sCcOHqYf1olGtnNsEQShft
nDdQ6q+emtYYTwDdF3uVkWbCMHVzklLpaMKiUoiuYkvuaPw5doLFbkDcX3hz81E1
zQhU2Og9VEBHk3MHo5STdAe7zoa2GR2H9jXyO6TWEWHHf/R3DtbYedc1mlr2FpiY
mvRWoJvpR9uZxAbhAE/Lz5POcScRhmQxUi1LcxhmglnoqxmkgmGrco5X0QTCO8EH
d60I16tbgAiwBri7cVOYhT1TgFdBHx5+Fm0a+lq2M889Fjbc/osgCfSsX2drElLL
LfM5ewlYMYBOoxKnBLzckZ/twDhArh21EvEngAkQjb7RQmqvfNsfp4gvFBxC+OFi
LGj7vwSi3jBe0rMUYkCnO7mZqQK+XY6TxjwrV4TGdzyXNRHFgn0u9Bplv+6odJEo
q1OD4iygWzRRDas3xXVUtSsH71a/mI4lcArqrNv6kXh4TWZNf7iTnOd1dajGFJj8
ubMbYp25/srdNmD9cMqdg6lQ0ZabXmt+Bcio7pt08BIQQOHNoEmcUB7M22VWf7FY
6KpxIv+Da5fPWLjelXxHQ4kyPnQi3r5N4vzYQfwbgvgveRTvY7jeH+1nLf5cExrQ
Da1R3xWzx8IGK/CyijFrBdE7E7jVE2ar0DPblQJc4SD1jymzLmOqQev9TYXsJPfn
rHTgSDHeurzgHQWe9bF8wFQM7AsYE9SrPvi4eZEYIESRBQzch474C33RNpCxpWKx
raV7/N0B8QJFLttmqm7MMhfDafGlenWtsOWlV5fzme4miV7h3TCIgD+/SAwB9vRJ
5AzJ1YdDZM2Sgh7C1cEzi4/eyofIKAzlszD4Wiuhd4YhTZimF7tiyIxKH3FcFBsJ
feEtzTdBvqdTtzGne0h92VzmKP2PJaqD5ObAJnrR8hjYynyIPESYLAJ0uFoZS4Rx
gxrTqh6Qokw2JEMkjTlzQPSFVQUPq8xQmM6hBLbVrjLRib8NetD7MgOA04TjB0w5
a5kTmGV+oNBjmK6nmCRd2tL/Ae6fQQJf+paRA0zPtzBbnzitvIk+rBHQZSjhjG4g
B/w2ON0gUKiIE8jsq3kZfjHKIcLnQ6ty1hBM2mggMEBVrJET45BnGA2s3vH/ZwXi
xknnp6HjbgccST6iwULbsksgWXUYq3NOsHDBk1+Czm7jE2f8wK7+NbezZyZTrOYW
Os7RQaw4PMCcA7h95uzhvrVRQKglcjYvxNyMchfWmTv2iE/cy6YzqFeSLGE5XKDU
yvqCRvSfBnOWCIcbdnbXKAP6idD1gr5B0+/rZ/8psB+/nwiilQqenjMqOCzOQ9vE
PZCRRsuNlsI/cjImNp3us1K3rgXG1vdRVzL8BmqMtbQEDbKcN3lhWI0Ys4vbEOID
4GhCk7XZfGSKcyKJ4kffT3kwQ4sEzKbMlp3wEVuE8VOw13RAAdxRji15dTbslrlb
KaNY4miafYC7oSiZyo5QYkEt3OngUpbL2hZ5o6TExxSkub1QSeqg5ENvkc3O5tfx
5ywv8TQ520Fv140OHL2F3de11IpWs8P/oknbKda0yvq00mEpg3qBk837OChaZhM/
QDoRiEHcQHxZEYQvi/xwh2bub67ft1B8gtS6u2yKLHtC5gzkjsQ+nVvfFMzfDbT8
ruqDkKnPj+kBDQg3jie7ozj58Z7lckAuGlnzIQeTFp/cY0/FAVgn8w5YTlbidDN7
EuppI4XzWIxNRWulmGz0mYCgsms0Uemw1uW6GYIRPrxAGhZAI/KgZfCjpsm4r3F4
/U1yI2mSBinfaguD/MTz96TIjqozPE6B15EnEgpblh/cz/+m1srMQqoEmpNDRfmz
dFcAPy4fkakoKLtzUgCEV5w/nPIXtmfjtNPKhPoiL6eC+snYFH4NxwWsSCDN27yB
v86lqRkmeWh3RYF72JDdA2p5puBRwIoA81bbYYAor1uP+ZxdBlxSM4e9pRrNTg1R
ZisuWoYJKdlmtc4utFsD3Wd25v9OnGhfTkW/XAe4rN/iBbQLyB0rH7BWtkcq+AFx
zfsJsGBZz1sI1zSBoE6uN9itGUA6nkS78bykoWGS0bqZN/BA4ojQNlvWJp4EOgm/
aZ7wI06VZhqQLiQKAQvclTPo1hO9d9/4rH7W2lhKx0RvatFRmx8R6Y6dRP1+JTDV
/GERhKC/x4MNDEGW8EZDvEt7Jhr4kuUWpNK+h5GpOcL5RgK5usNrZ66deiFskAYD
0nEvtW7kMCLJOkCsot3s2CJevg7QgXKchgekwvrgUQC1O0g+kdiUbcs1mmZQ/6OX
1cu7DLLfa3A33gCIjALOkgDHe+9C8Lf34EIovG7NihrO1f6dQiCe+YyWfMchNEej
mhruwjyqjQY1gk7RIeHo5Vbqk1ch9V9+0XukVwZODXI23AvlVwV5HBazyS3N51cO
0G7457VwqVXAcz5Yp6DLwcLQ3xjPqMB/Ju9Qzt2ZvcC2qKelZ1KXcNznPfCd55bW
gYm5jQf2p2ZJh4ZC2y05CxrNTGVeXwSahPXGxQeapWlES2df9LZImqqnZCKxDLCG
8BWLAB8yjRnnuHI3svWFvySGQius+NAi2EPAo9TCmN75AvPoh1AmozyJsZGDw8pe
geAjA5k7Cdt/qLvdNvinI1+Wsr9vVYkvUCmq+dGXWpjAkEnl0/hL9v00n3AOyT+e
ZnLGz3+Tzcw7G2CUhrom5zxqoR0edLoyTetZ6T6xNyOBH8A/qIYozoKTjHoUrNSB
2l03Z1H5/rtV4dQq0iuIOCeHRMKgX9kVZLEBs9PFmNe9DuQ8UooyPkvF9ohfwWJF
6Sdg/6oonMm9jeiHr9TC677hT49Pm4XjbXh2+cC6dyhA1ZzDP/EyURonCCkSMiAV
cANxm2c4uW8Bv3/NSybOSgTyMlBiIGvXQKi1oNqoYQCm+UjX9cCd1t7EZmQgRZ+B
mEBmhdN9KXpWFVLTZa8keVsyykQ0TkoNzj5J7PedQc0A4B+W8+2Wngmha7zT3rFx
XscKVO5JVtMOUi/smcoW4OPODRgBOaQYXExPcgM5EzEsQ9KT+dGJPUsVJBMRAGt/
TQZk4YlVMaHbeDnVolZwsOVpBRYjrs2jrZrHkAQ60e/aWeUXsiaQ8bT9mKH8pjwk
2jEkucM2rfOth7eHmsN7WynypUWJzEYOJ/V3tfF0qWzoVj0LipitEoNTPLkuAKJ9
+O/49oibDMMybEKZFCxpMD5ZRRzRrw39FodOTC081pOejc8kCvtv6YuCoa5wubBz
PVOIurF9yXJT0kJ7PVlsdH70KGsGu+22iCJGaJFGmh71xsBZYQP7/N4P6zQU+vbG
VqC53+lSF64vYdy+gcn6diIJgnBt/dp0uRD/3flYGqeStogdc2EdnjLYAgcWRdLL
x2gxap11p5CpIB+muTTRkAC3n3nf9kLC2RZt5Jy9F2dXn0Yfhlv2erUEEku56St9
12ogvnOCKSGJcK1sLiPxrBn88Erjytuj/oHZgWbvjrrc1oyesZTbE7tE2eVOyuei
mA4yqM97+mLaiHlvvOhPIoLxBLam9zqZIBVzfb3g4NEoI+0SpxZXAAWaw+2uQEzF
Xh4YcNXSNfVEEyH8KpJsbzA4PikPZoFoktZiipkhyb9qE/onzMqfCQcNsileHVi1
uwRpDe2Xq7cx5wbvtEGcTh1T8gb/Z2Zso1ZEOhAFuj1ZOsD98+uAlory1/JkY367
/45lVmrm5fqSP+TqK+t5xq3pYkO2WmxEZYsBQZ3Adem7S9BJhcVFHrVfvFFnMlH+
zYX6WoaMNCmcOUgOVM4rIFgIxGSCQTvzEHDM46Vmc0QrSCt09QljWVeqIjk8RTv+
VVi7lQ3Ip0dLOczQkvJmBDZ2hZ0Hm3lT/xEw+p9ZWukdx9MUbuwbwwc5IPJd72+B
h09RcbdVcpA6M5/t/buyThUKjJ8FfiaEmBxRN7VV55OAW3nMEVeW9HjkYuhIXTVH
dk3rGi2aOPX0E3J5vWQb8PkJoEJmr1UdJvLlxjGNchnDPrBBU+xqg5shTK1ll7Mt
zZfOgyUG9TDEOQb1uUxc0u2IVyYfs8Mm+uLNQuZq/JPBnMdIY3ij1kniLj+JlPRx
e6AyoPkza2SFh0pi/tXIJThtmk4j2DJ0/b1LmDxG7KO4LND5Geh7xeUpj2WrJ3Ua
D25xRu8wG2mdsh6C92VcFQS9oQ82XTMsPPQ0I7bX9Yn9JFL887JiBZr/refNAAqA
uKsSNS24WZht0QH0MeZuPedc5Aifrz5CYaHgko+DEwLdiL8AXdydqm8vGfAXuewQ
UKaTgmv6X40ro8rBLaWZ4Y6sb0hdBaTVgDDK8JHMJI+y89cnEKKM1Oc6fAWoFvW2
SRg0ZR9oSBU6/A9QdHzBkRtgY66xH4qVzDPH9/KzfRTQeX7UMOrwwmW5ExmpmI/t
ZkMjcEGXYZP2GENmw2vn8d1R4fhjrbv4cjWnT5VNveIm8aT9h9vDWMNR37bJOEpU
0qGn1b1JpngC3318kVFlULX3cXF/jxnmfPlFcJ6RpTgoEe0LHnoNIAnEfN3zPeUP
Q7Q0JE3TKCYQQRXLrZBp33pof0qVRMLtlmL+nxmX0KSTBcQinQHP2N20Xv/q60KC
qOt3n9P0v6E6XMVO/J64q8LK/C4QasSa3LHgJkyYMcawkSGWbLNqUheZ1em96zju
bj6XpJZUDWhLoI+AprHrsbiHDRYgiXMa6haLGcMxHWU9aqAwRliECN7ey/BkGAAj
rFAN43P48gag4dWoLhWP+z8TE2nep76Ets+O/A/L7v/AP+37wPzdMdr8M6Qexb3W
UbbPxed6vSu359140zHdNVuqmKXLz+ybJjBjWXYjbroFzky2kJYI8iKQI+rx0Q+d
EF45jMrJQgDSM+wb+2CvYFlnwecZql63Dl1MQHxaOhtiJR0bnZtos7A3vopRgGOz
cvIDzCSo/yJy3ptM4bacBbJPUrcx5A37DWTTY60g3A/W/qbNw8ru9yJu0p76kL7p
KAG0tBtmF3JMUn8Rn42vmjVZys+KytM5IKmSaQWjGnMb/070CzpoHeoQbiP9zQYz
s6diAOEoOZzajDDoc0rZp4fSDoE3GYITpkRol5YINcMXE8iQGQv6epqDpNq9Rhsz
TJzxtoBWwxgXItgzPhsaVhX79bwtyKgRlWo+p2cCwHW/S63O1ptk+VJg9tl+U/UU
rDhshV6x6NC+MKvzD4qCTuI/pilehoV8GRuHBlTyY31ZNUjGwGKEzaUkU+R5wJbg
DHx+cgkhalPtcL/JXAVFIGn5Kr6a+qu8zmDm8mEddFrcAObB1xOTn3RR57nPFFq5
FeWjhfslCW9t/vOHKhiwefs7+h+nPJOutbukfnBwyKXP+BRyVKFrHjGjXcJCw76N
LyMQsr6ZpPgkDhe3TSQSB5TvTa4dEPCLXtiWTL1vFZBzx9W/xNDqiex+ah73iNSz
EbTh5ZFTbVWooZUzkhuMB339u8eIEEYDxJGfvzoxFApzeZDuCUfBkPq2Jwl+VW3x
73gqUOBJuONJZaqax9NcCe+tsLaEOIvBwMFIeAQUVBhZF6V94E0LcyI5efDBqmJP
qdnu6v2RiGWq67vDz95tLUEEUjDSh5vt8cICoQQyFcKE0fAMHR0NDno6JydKVKw1
c41Ve90dwNYLmkXD3VhoTw82T1KjqjnPg0N9v6BQSLw7kVo3RJeuYrpr6gPDvV6z
N1d6FX9Cmrwl4Qg7EI0Gnjiykr4YUCk3We5qQEv+eDViusa1nlEKNOs1FYjbbZLw
Jcvam/eZ36xl8IGOHwxMcp7e3eJTyaHlF5IM9u7kb5PExwwx0SJBaajuv0rYzWph
NYAt6/xyn7sBdVepthMnLAa0AFIkRLMqqmjU6BiZp7sJ/5TffyY6lwMyiE+5jUgw
JiXhuKRH6E+B8dP0cnE18UwwRZem2kP+wq7q/l1PvvMsZnFOHePgSSUlKSRFGQQV
yaWoTRgERAVX8NIyMMdyxtgum/fImYipax1f9pUaJI4sUxHCzxkK4LG+DzE1/TU7
CJc942rexsjqge9BugPq7r7nkXPJ110OV3meX+jTFDH6VZsQ1SdNXMos0weXZAup
nBOTfhVgelxL7nofrYSndn8Wq3oN6LmZo6FdWrD8WQC7XNOztDzBPakrzMNgNcjo
DooBN3zqwK7rUII28e1FY5ocdNefj/O5ixOTeYd1qS9EzYfL7pUzwenzftgNN8vl
+51N6IboCPErbRknEI25Jx4YpSGgnlCH60+BxJ+EQN3UZ/TLy9t7xLEubXcjqtYU
Bm7Fre0Gswc2CIHEZUdtvIzO+/EaClJRdh9pZhNLBro2Ui0cTZgBvQY6R9uZL/3W
G9gEWcPuZZ+4ngx9Oj9O9tNsE3M+f36TZRR0LHIbEtcbBqWMz7m2snX0HPZ7JIDT
JTeaaKgerrX3CKemuYOm9IlsGe+V0pQzrXLSyDb0rANGvwxYXAPAOP47C8ND1BKN
VwXLSF2Mj4XmNbzy2vRmVY1hPt634igXjlSaWrp3E6QlrG9dqxQy7FNk9vsLwcIq
pvGu1Kzb3C/gX7kDQzMovq55W4sCTONCydbporp61DzF550g0jJMu6qY2nD01U9t
xgDS4LVna0yIINN8wy9S+uYN7vG5Pro4RHCTTEh3BWpHd4T7O7r6TW/SBiBMW22c
VnmSQ7YeL704MBOjyNmGnFh/RGgr0IL4Le3f26mQdcsQv2SgCnqSAY2nNEBsHG4H
8gEpRfmXeLaYzUOIU2sZoRThHxiYVsPT2iKj25gdEOyhs1VShTQj+LHBr/C/jj4b
hZFk+0gSxXlgLmyHrFCk/IehxDyXLOaZup441fSxg62mQIBzylcYAQ8Quxq0k/ub
vppWU8CkfWgJHDzsUBW7OBoeo8DnxaRzbIjNzilbWwI4bFqpropAIgOZ4wYSjS5L
yNAXqDYoAGbzf5T6RWeOtpVMJaMCEzsuMI154D9zh6v3mjwT67XnvNfFU2eJPBWW
nMVXEiE+Dz2F3lYBH5qkV3W/as42GS7h2xeKodtflckqBcsstE7mdRWyl5J0ff91
3mwvoepz+96HHFFgfTblIabawpBr57Qfjkp6M2yCTBnfuoS6AEWTdAR45ce874kJ
bHqARm23U/Kc8uxT1Pv3jo1QxPU3FttpIMIFTe7Q0fDQ4Uj/J7q4b77CV9/5zCKj
8a6MCuzGJe5jWQcrCHqQf+lwdSXACMp3DoTjtI4C/IknAYEtciDTZg6XixxfOeVF
h06mcmRHIuX0dAMhG0+s8mOyI9s5bP6kLOf8PUzwLvoSP7VnvGBs0Y4isEWZ+QBy
esuP8zkxlgAtqxL2OzExkEOgylUsrPwgDO6ALNi2t5sX00iQR/As0FmcjH/TvM0v
qVQN8T/XtxWLRD4/I/852R1H9qJD4THj/EKRinSPsEQSvH0svFSkUa0Zjx3TWrEs
8DY4GrYyLhz8krKxuXBTtNmxfDQCJTI/7Cpm/M5EvX1ZRnArgtTXIY+qjvz+1icH
1lh5EyEky8Y2gWmiiHIVEn6XjL7piOqJsxbx3vmuubF28u4IMgr4puNnGecNDK6j
DEoXOW27Uh3u5QLbGLpKKuK4IT6QuH1OtWG2eFwHAIcoRW9Yd6ft4zQeYa6BeKZp
R9SrqAEsrXlf0G1HsE9Og2QbdD6XvvGceiSXrXW9Fhm59RoYAOMzDc5uZlS2wLin
Pd5HQRgILQJ/Yr5bID0dBv81RpaN5m0T4ecbxfpFTZfNQD1xwmTCbY6nx//jgrC1
tRwgnRjsmiLRRgahrgfQ0J+Zn6BajzHn1bQK8Dqd829D66axTmEBeIfv4lv1qiRS
kITHbqFpPQOu9AZ75oJnxACigRCPQzR/xmGKrN5p/n6U55SxD28jztttL/ProJMk
mRjSAOtlWnHtCgpy6m5JZXw+SmNdapx2gQp+wMRAwiResNIWSuOdUBENw/pHsPU5
mQspzSs1DxPvXiroHgaJIOn/T6yP2zOH9WCKb5IhrPrGyW2Po2j1loyFXoh1oifA
8gRdJG8jcneF9sZaQUjN8n7ZIuGV/2xnERXItTZhEnB7bysa6OaRjaAlRkcVe2Ju
nZvFQlpmzsBNc/AGX7lIVMj1gkIN9PydWEmXBRoPDx8LCOIZ27F4vabvooIHFS9c
G8Keg9yFd9ZKDclDYkSnHwWLzJHZ5abDkMDWKNfrrmBLLY28UbcVOxGiqxijm/He
ILpgAeZDBFsJDrG0UF6FXCRkVjJ4/1+rfUTRAelN2Q8C+wLEwmvZiXK5qSe2MlHd
c8vLlVv6AfXQtO+BDUsjjBS6x+URv9mLzFbB79noqp1VgeT6OBCSptUIYfkXMNNU
m1KJSEUDQaW/+Z8ggAgKI6XXidJ1goy48VCyMfw4AP2/3Hl0Iwy69g6CeZGnVr9s
5/PSZ5tcwS2l/RaUt8fvYRExfWEGwT6gZHvByKjqf9cE2RRHwUbLWsSWhKSB66wi
LnL/Hlorj3Eme/mdQRZjoDjMM3zkbyKiSmNigqpeu9+m3cAhXVwn5/JZhhAjNF0q
2lR2amMMLDMlg5PJw4V1h4VyqP6bueY6K5d3MOON2WVjN2fCkL9QXPQkmhc47ihX
u9x9yTWyJKmCFJ3KF5RPvenDjuWEYUXXxKlkqiUeEuYs+PXNUakOCkPl9RAgzccP
Fep2mHoXVbzudXDeXinnL1bq3Mt4okg0yO7StKvChID/uNdxj0QaSca/Rxe86yCz
GE9GG4bQSkJdq2dvs24JvZUpGzJ8I+ftW8sGr8LOTLiIM+aMkdzGTJeAiysQN/T/
aCcfGnLqGGkqLZtUFmuLYveG1SghB+kNqEXTPs6D/M2RentNUOUZ5e1qIZpD5okQ
WM0DiIbAcLvvvq4GujGB6yD2J1w3ML2PlnW/a/Aw1OH8QS2NTQBFa8IgMo0kvJUQ
lr6nAPNiQVgPqzZkt4LWGn8eGLaznkrI8sq9ZpcyJmvnsjeCL9Nno5M7lAjAu0s9
cUqFYAZjhBuJQZ++ncnpmkPlUfeHWfYRZysNg63y2+9wKJAflxEmwMgHc4odhL6Z
oxSZnJ9k45uMjmLBA9u80B/NPhu8N6EhiB8WX+TesZMOOqOY1jFfvzg7kG4P0Wpk
sux/EDIH4jWlZZtcv8AtSAW79qVZ8ZRWRt5TNsRLsKzL9fCNTlPPqFAr7nvGGtrs
H3qhocP5loeva0VNScz1H8pUfTvdSBJGevOfkeVFUZBrlRH1aeaGdXDOD1BK1Krj
/G7yFOmkFh19HORVRjvn+P8itB1IbHEtaNhvQucZENRfFjwoETExZiBxzf6kv2bd
K8zWAuCxipaPBFI36m006IN52YKUKzmCZpbTIFtMrqW9hq6l07zoKlYOlFNckyVA
j2DVM2j2Aa4bz++SM8Y59wG9yrGlrsb5YDLGFbxO2WxgQIj2bcyoyrbn3bZ6Rl5x
4A7ozPHquedlbGaBpzoavfZFIe1AQAgO7vnSlgqhw+/Em4NlYySgpyIdLb1inxCX
b+flpoybDttG6WbiXQb2wiF934c0m8lwTepZzen0B3qKq4bP/8ReKgJGXVGU4xsH
AmK6QNxOhBoEGFh+IIzSlshm8Rz77gK6H75L90XgS3T4nT6hCuVL1oyvjqfKXELA
YbUjM5j9jLtXKTugRp6lxaLrL7zzBXrkuayzPIn7xQ6/z3LUgDo5oWIbj5QA0stK
HXCL4SkAyojYITZNqhEFOow+1Pxy+AOp88EdBvjBHEU6YZOc2veYpB0P+SEbwSqG
g0nNAVdr9zyF9G8BowlWA4eyBpK6B9V3GVSMlfxlw8bMMsKk5s8iQfW8RGny0kQL
b43qY1WvXKaSM8Kzn+sClkqQKYRLQhgAhHt9k4jze/WPeDEw4ScJwF80T1/vv3YJ
vRGgXDs7sdQzStkaRhJu/rLbfSFJ5OKj6EXbblUcjcFGj8BqPxXqWI3N9WoeRA+O
WHad4JnGQRmskSbopQAZ4pMvt5i6FAeaE+3et9C/NJmTAYGcKaxCwWzpHiGyV/nd
j2SnGicNxoHGU12jZy/8KxRkn+mkA9oS2D2adD70T18PqetEEUMjmYejIcQ8Z9Gi
gYONT8yaMV+9jhpLY6fclduTcXYBCDc0UvlBC4p+OW8Na0F2DJm4m6ltPi2C+SJT
fPD7clVCwQryd3n7bDaNQ2ZA8iHyPOL4E6hNRLN9Ddd0jsAdBy38hL2Sx5CtZ2iN
I8b5klUezQhgOMYJCIOhm4gd6alkdRrZ5k1mh/CLxYQL2fGC+HHjM1g9eMc47qmT
xiY0Bvij03zaF35gEi+LQP0MElITttCY/8bYYsUCKFTYO+7YyMDjeviVt1Fpb2EN
1SIERaEFAparPxmi3alIPGYAItRXFBLFyGJkyWca9OPT0kHQozqaAnquA+piRi74
+GDHh96LFlEoSTJiNZg5dczgdWhGgHD2wqVf32EuLApaFNOzfiF5SojJv0Qh3f50
OZdytaDNztESwTNJ/KodKwAG5JuPSJW3M5a3twA8wqqQS2fBVjthRzjfGPwfo9Is
YVNew7Elkupn6OxASCLb5tukl1WhFdVan8B7h2s9gcixXYOG5CD4mMdC1+07hvVR
yZLQ9kPCxo8wXGFPIg+ESbLVOrO6GztaZqIcd8FyIlEijEdpzg5NhIITKbcu2lFu
KqfadBq3pd3V/YXqb97GHXLQyThF+2oOoXlFaPSBD4Bla2Q+BMEA9D3oz5NOLLEy
bme4qv4vdNNqgC8VDMf0u540XBEYelj1gSuKlyuDtReIwgaZTgGYjKhfnAuZFA6m
NopqAUr2J+9fVZjJURyEyxNU30XtjcdR/qAh5EzBx9W1Vy1gkC6RrjaRhRmpxJSV
hjfksqFBlFgYnKOoAAYcR8/wC72TEMMe0AT4I3Mc46m5R5nWyVqgEE41d53PDFYP
3QbxC+rHGej4Uv78ufPCDLAvdQxKa0yLz4V4LOo9GFdSgQEktQh0Kd3TOkedaevf
602vKDFawriJ7jb3UMI+T0J6xJhmx9ikoD9y0UKLFWdRCZ5watlqidlqpfmRPxXq
TFY4aYSB08L906jNkc8Thljty066cQFtWEg7eYVlBIHaIl8KuruzdH7JTcEwOYeZ
SVPhdpQT6QZFbxExPJS0KJkkWSZjCeXO0hHN/94CNJGu2OrxZJfbGUSWt/DYzKUM
DD0hkHmXLoyzxppWd5TRs+BtjXFZcxnTkq2cnOERG5Zgt3AT44iHalxICQghQZXu
tRp3GoO68rnOfalUI9ibbQK+QVKR1jl28kJkj6/YJYu48TSaw+07Lmcep7CFl3NR
JIReSxrmh/T6woShuHn01WyKDin3c1RQ4ytQsp7i7bmVOK3AlaMvOBeRMGJdUSWl
D0AnIRwzjhuJkuCn8G3JTe/9tpnn0EGsSkuVM8d4ZaaN3s38+OeiJP6U4hUa0n7t
SfMdcUxeKVfdyvdQtLtnZ05qmaLLoQDUnSBE2Rpgw3L5CWsiXbPiIFIT2TK1tHEI
Z0rVhzYkuicwent77gcO4iMxN0qDjWVt7Dk+HHpkhmGus10s3QbQj6ULPKvWLZ2W
7xGpTyZ8W/x15yWY0kSTFGOkHj+74V8tfiux8cow7NELDhWqdrFBitHfiCjYH6rB
KlK2fTGcf11y/zjy7fm93Rxxat6x7O0LuJ1GuCz1AH+OZXbRBC2DGH8LmMCLBunN
AIZTnKtw3tshHO9EMajMBG+AinWlmseKcK46C5FbnbsAXdhRe4ez8QcP4nVZkyP1
Decc1QinbPAKIImdo52wMLyUC7Ifmj/8Rupi3KfcDou6Ejx0cTS98kRYJUf35jIt
lqsLpsXw3HRK01D8VhERuzoqqOHmlCZ6gNCv0wZfCTHnbi+5i6yqmimSJ5PQW/1Q
M3Bdl0F+5ano0gyLFsNYWntB2MkkXDE8gjMnctc5UbdiSFO36lQ0Mc972/YoEnb5
iuDtP5XFjXVEZfewkLPUOZbYfySLinSWqCdHrQZDPr0rv8xmYo+9Rm/tSPctreP4
99GbJPovljV8EqI3slYleVAT49WqUZZ6QAS0LGn++/8VZ3rSQKeHeouZ6GWci5Rw
eSiUtTQJBusyh5kGFzpQdTh+UlwuqgwcuAbCXFiXEtgjAxpp1QIhmoIq0rCtd60+
ybGfrRIEd3DWBHnoLCyFQZhMd6FcamnT6JTS3wXH3yrwGARqmd3NOzGXCVqpW/4L
kF/GnBMkT8yhHM0Gipk3GVismEBXnsKtvnVmdWzeXr6P/HWZ053AhDBWTweaVcCw
c9g+vmxF3NsYtg3I5vSiYTh9fhlbJGTbub65DGkVBRTMECIxhWG/N6/202EpLd2U
xT1nWsLjBGXi6HG40f00OcwE3NdbE59aTTxWl2W1dZie9gXHbQVnunsutNGI74Bt
b6l76G4OJMphHOt9XcsidhXtNY/YBIT+hciCx1hoUNHG1ELlbHPwK6Z5HECps0Rq
YBbfTisTOCXgqeay+VULdCUgVtBJ3z/lyndsxdpBmZ0QujqZbWkFd+3w9TkDWnRm
wQ3rCtIP7MSgMieixu218p49FhV6U6jv5VnBYib8Os0hiLrpV5TAZDmu1kuGJNvi
rV7s+E0BoyTMIG/m3MD6klHqu9puy0vFqdaMsfuGYbBpYG9aJTPC1+6a6klKvYzo
2Cr9+HqnTIMciPI3OSIZY9Ks5H98HTTzP1SVgfPYQjYoB5j0cVpfjYvnAJiJluA8
xWK0fNwiMLN0TltzcAooZD6VejkXPfZuLX2RFovWHjGNJE4gULF4pz7OgksCpEkD
CRFZH00/XIRgKKUEWMMy/b9EsORMLSSabhj409ENimxI6Gsrh6abgoMDB7RO09/w
cE+LX8aECqUWRBuFUfmii+HfMDfb9bgVOKP7lHV1gW+tTrqpOx/XpfdDUS6roHqs
KuGK5fr3d/Fm+O0iN5rASdy50j2V9T6zigvPoBkhv8NakIRbIvh+tbm0UJRAK19t
5hr9DLO0VVXOoupD0FKYE1jVIhTBtG5zdhUuo2mpiIjtliUMaf4SsfgadF0V0y9/
94Qap1a3SvOi2uOOXHze7r1mdQXgx8mfQgcJXE/ozhteiTZ1C0ffX9S/NZbqakNc
PPYbphEoyNAJxZff7cARGXRnHv8VFJftb2wynNJad1Kyj3tGWobNc3CQCLO/EFsT
6WEQWDLlcw/SlbrdkbZU+rwnW1IQfxNEYsWQz4eytoYb7BPe2UmFckRnbz5FIGQT
Yksain79s80y/uMvWHzKovfUqrESjveEZe0nNM2sfzBbPhMjT0k6cBbIAarMREKs
zF+CBQRqZMa3f1Cy+o90Bp0zvMlGqryGtoz7wfMjhdAIO36vQ++KQv93m2322xfC
MM/P4xky3V6ApGDH/Gmq+jg7+onQysEcRQ+3dPXZtYzxHN74wJRpA3LbhePjevke
CK4FjzmqSHQ9rms1QOUSDlVuU6qHYQY3fRgp+9Z1jQx8lcferfhjUWrfL1Wp8NCa
Hr6YW/pjwQwEQ6Ka02PqTpPW+CG9FuOQqqab9HovllHfFw2dsoARb75nOPVMLMkc
3Myy7uJCqFF6KUh67NKMzRBay01dGb3Fo1MLKW+sKUyPMw/8xzYwBpdFskvxr8At
rYL1OjkNIjLFoaAk5E9Oh6Cou+ASku4Ash30LYP+likF8tIHPGjAhLPndeDOB5q0
zhJyFatJvHHpzSzgP/IEUSgfRzrW1Vv31sMaeiIVWq/WQ5ITwwii9vRXfXcAdKXd
xx5aAMGn4QknothuNfwnHHSc/l0DJzDWPwtNxZ7A1rnfAgr8gLyQWpXqiXnZ2id7
AH+tBs7vfMAZw8y2aQ/5qDPSPuIYTKmgaym/NqKP9bQlDqjRgP4l6p2cvxPrdKm0
qcCq74pCJi+GFDYv1WNXiTrlTElulcDzG3cZjTCXhPlQHEaUhD5GXUxDtBlGTD+q
kguacbD8wy/Rkzr0YFvFGzGXAsrKTYUXWWpBitq0g7lWgukgf3Q1S3rC4tHAhaIE
7TYyIQ5DlB3shFgncGCkZG/uOJ27yosoMrOayZ165/wv3ZK6UfN6WXmYaEpt8UHZ
U2PrT11JNshEuuqpXBmaWrPyRe5aHq2mZdEt35wOHiVFYgP3vfh96NIesxZ8G/QX
N/jbxSw0tRJ77xA6REUcodCeBlpZpqJxXdNWCN9S8ZCHuzbv8FYnVXRycuikfshR
KDJ7ZgUZYIcQ5bkiZnMEm1hB6h56ZKH4Wrn/rS7fcdYuIXRpUTydTJjpRAVpoK8O
eYehM5x0LvCIZt9nPrE7A21tXvNsYtYccwL/9Ooyn+ykCQLbCVzprjUl9il/5bQ6
NfgLF6Wk8piORP7poc13Rw9MWi+PbXIaWmLKbRXh0KVIc0LTvpQCt1rVhK+dvlnT
GB+FAqgjw2uxkjVFuGuVfLh12pGue6I25dRdVaKlJDfAGJAD+7a1WhVhQtjdrMl8
uaXluSzSqi4/LYGbNJ6K8ysna6P+qwMVrp2hrh8B1q8JuuEghoaP+rcc2vUjvoCR
c5yVOPxfxUyhqDFwEQ1lDHaQpdHDxsk8y3FSj/QyuOOHGGyUMQ1Y2RuVU7hz9Khi
Gn2Z7pHsh4c3YPDYTNvLp31M17irYxQiHzoz1aakBKELLs07tXiqGNGmOSZ14U4s
ljo0nyVZC0JpnL370TZvsQfxy3s/yoi9hNtlfL5bhuJbhIcvTlbEQJWFS6aZmHPF
g3gRZPDIfH4gkRTjY065ZGP31ref+jkbZWl+7KUa6SbhoHRpmaCsYp5RVjve1gq9
hPf/r85iYA0vGjJo5j8a7oGprT/IX4hle0JlYqg6WTtjbzim0cgsRk3rypSs0CYE
m5gkF1RcpRLoQqsK8l8zw/PXXbuWYnYGm3g/9qeWVHMfGhc1ASo8be9WTurI7THD
F8E9AO/Z8hxS33AxTMAeUsclCL8ztLh69kZ3grEGyhEAMR0xPTzqfkjgiTFmkskP
c3WpnphAekFivwaW4h0fo/QayIJdcsvIlyZZ0/1OPz/4acpFFdmHbR6JNnZY2xH1
OKSskEMc4sXmy0XhDPz4c0RzfhViqmzTn4erd59SaxGS/SWS5KJTT0mpGNeozKu/
wFpXq3vXFJ0Gnr90Jx9Wo1/cB075av3Ddt3JEOO7wFcPyDocAVD6tQ4jF8fmDvQz
YTYA6FISApXLqKJH0BAuWCK5uem2kyJbKNFbCdiuCpzKIBAUM6R7W/Xsgb8Lx/g8
LLjp7lqXIC0BHcg/nzserKJHn9vbC6AnThNYuc8t3qe91+SSQNzWu0L93SoIlSSx
/cqmFSBg1HLN9iB/gFsrmqdmAEy9u7+a6E8o2TG5okPzNRdduJAROF9o7RP4jbo/
NTXP0Q2XGq1A6t1Ypmb+f3CaQUvDW4TmFVCeU/DDz32IvMvEFTK5oL0/t4LFmvED
My4rzppSPwcgEGNtkHh8/DVXmXKglv0T12tVRHisL0kRv3A4pMkW8PgCtpUyD003
5X2cEwB3ZOg+iU+a8llGFAalwvleyrE9yhxi3WibMbHXX9PSSdWsoEu7ZQzvatlC
BWXT5q7FB6/kDCokwyUcA4GoeraHpW7H+l6D2zNekBVzZI7MI67e5KHQkvpHciwo
OcVRimT205AblD6Qsjk1pxu0q/HYpOrw89tZ7yBpSbHkic5XhwJTiXckL4hOu9O4
F3ovqiEDtdge/NafUc3cT5gQozt6Z0qQ/BBhPQ3te96LR9SRd+rtxPv/QZjf6GCu
FvwDZlDcGaThMzDc9O6FAgN1k8aHWYiX7pTVBJGnC4j5QUsQRRewjANEIMvvdxL8
ecziq6LforzesY3fNcdsrFwkGSWww+INYEL05qc6fd+M+VIEBLux3IrxBxpT6aq5
BHteVu6Wd40DVqiNUPO9VMb4hOG64nz9WLW/6Ooz+FSVsYx7U1bt1PmJIWolXqB4
m1rqfOMKxyHG3pMYOl/xcoKQWC0+f75zu6tnijKOvLpczzhw23SsQ+b5CzDXwa7C
y+hunV1/Wz12v39QJwxxAZvHKRki9Dd4R7Vy0xnbvsPOUQZ6L0Nuwe/LHCygZU4e
0vLSy3dc8oXH6WOlNb7u2oJ0Z+pr+yts867uC3+tsWTeUvTVbDRIcdX3+HEVM2Ti
XG7Tepy5zcsOPjDLaZl75+C1oacrLxcFZdbx/p/DfyqXl7pzkGG0cnbGfRnejVoJ
Y2dLODAMm5ePx+4OitHXVOwQSoYhG9ou+8haFurNqhxZDCaKxSX7qdTGEBk9LTfN
O1Mnax6zyC57CSLsRzCzWRRSk+1K+eTnQF3JkvqoPiIP/849pjedVUDASDJyrABQ
p9EuYPuDRUuaoUeWEWilACGB0Mk6w914piOTvs01tLP7EhWLVUUYe50iWCTHjXzf
yQgqoT/wT0BzpBoZRWEo7Z08cW5sai14Rfi6Y4/uCXwXxKtPTr4gY5NqbRJhE5nq
VdXfH+133RAwb7Q8TKfxN3rMheo/gPvbarYWo7ngd+Nw7dQLPqioz7S21hAUPpHh
mF+wu0Ig1tHKkS1nUfxTfr532Qrb/1Y6qUNYpSWV3s7xOL2s4q/2ukbjv8/2ytMT
DrSf2L0Wr0R2FUsIEvYX9G+qK2MezJ4fzr0btMZK5G7fO7s1xTu3lPivQM126YA2
zRCn+lRYQPPHNDqrFArseeBv/i4ByF9j3O1N/YCFDzw4V2f0qiorE3PgsTrxSKF2
R1Qiao5S7DuwaJG6qqha9WCu0uWfZYMfSJe8bwCUaxnUlBd3g9UnGt25Q2knwyZh
AusyVrOdT2h3hfuba5IcPfei+YmyxUafjLLtF+/gq8JxthK6DYTuq1mixfSZuy3g
ngXidE/AgI/z/SXP9Ir7/zaZnbKNmLyt+T03u7LLln5Jz3OqQlenSzsHLu+v/BdG
c50MMbXF8KM4HFIVms7gycjcbq2AlkxK9wuYDfkE2qBkASkxj1L+ZpmsO3XTCtkQ
RsKAEYXw+dDBZ/Rm7O5tpPR0rDBG6zh5UUBke+4FrW38CSBXtjb1dC/qFJnp67UR
lWOnO5x+j9nSCXZWo5dAbemUIurVdctr1IX0wRuoRxXHELcOrjK9cq7/81mXv4lw
qUpNhaBC5W6nMXe9mWPWYl308blg6LAet8H5HF7zpeIjvEAcgl/6FptgLgE1/7wt
iVEX0hMUJvuT7zidKPndXaKsVdN4LTJjsikHBIbkoFnuaRphnrTtsYdyykFgvqbL
+EPBdb9irm2+Qa3TUE0kmuc/570n10mYeg4+kyDrZ5EMxHJB29FzzPVnYqpJ4WU+
FqC7KjHOuQlp379JxDzM8MbD0ehfGGpZAASfpcttxd9oYJUaxzMEpC5LIYEUGHn+
VBnxJv7H19/gKFWXWaIMYUXw6NHwC49e3mX6PADu6oVkGE8NFkjaajDWW6pCxEJ1
0o4xLxEavi1zaChsvcnCWNgm57fQgE3EWXm6WpEHI1ILPFRhiH+Ovpxuk8O2T88a
nInCagYurrYlyA5vjj4a5lOX4786KClDSXhaVdTN6VjH1lSdWPwAmXZ6bgs0Z4BL
COBlsp+Xquclq3EaBZp2dxuDF3HMJWmrPjTh58ysbdR1b2k2UhhP3MDYZ7t+m2Zt
vadNKcXk+Ofq+9hnFStEN58swIs7CJ38z3VkSoHlSkOCpsnduVxW7sJM2GUz+dHx
1nHINBbFRGf/iQ+q6nXEq/RXn07ODEm8fV72LAFmrXCV/I9560AVu8Q6eUnSZyRI
Bq88TVzB79jfJONPi8YN0K+HzpI0BHMuVHdxeQYU1uF5ZvRJEOrXCHGZXCgo6lYP
Mj4MbvGICfBfK7/Lvq0sIglyRYcVQR5R8RmVTmO8iMxWerWx4k8GdqaCcXVZ2O6I
7JaLMiM8qCVJKqoboftOwGaELCwynQout9FR9ft0yg01lcrvGRqJYd3rUWMuwJih
TeSo1Nk77YLL2E8CwnX8/yvmT8T01hXQffzMSruUQGdIfxQZIMbEC06zVaDtS7Sg
Upo7BDBOQKauK7ksZWa9hD3TQkRNHSjSb3QpEQrJgsCnWAzbX0Xoj1KbCvjmL8UV
T0VzGlUYBmTOPAL6wODYUw1TmfSbijC5bf0yDEO00hF4IjQjhq+2XQK46rzPAiPf
Ld2qgKIMtYPA86+I91kvWjrHay8SYSUS2iV/YKhw9HkG6bXlU0R6XI8zoZHxccCS
w/zZ8rltaErr5GrVMSltFpZPsVIRfrH72Zmb1g81lDn+XEHTE/HKOVe46djgMJqD
yQLTNecLylVq+8yMIZyPwaSQv9pUXXGsVjyBxJCceaHM6vkFJHRO7AA44sPSHhDl
HiaZykI6zZucMvyVEQ/zb7oFj9gKYlrzX+p00UaUgFRN1mm7WkANNAZ3d1YgXn2G
TLQ3z+ZLC9cUkeozLLRgZUVfVZ8tL/KK8PRxD0xRIsbzxMvQJ4nf1ihw4gY3frCC
+hInXOIuF9XayLYSzqPLe3QulmJAQJGj050L75ZhLCPH7TWO9JpzC8hFe9wZbr4x
x72cLiaKxb402CI2YGLjQhhBqC5rV6uqYiNSWpcZNr7isklNhIk+LwnvWOWyj0jd
GWsAPwFvYWEkZGdCmu/tIOg0LUQIAvDwYcYKPMnzVcuC6ERHCG7FM9HxPeG7u9no
Ujn2XwyItcN9XjyyRUuPwivS1xLqq5PaGbmIxlIm71ntlWlWniR9LS75pyjyTaQS
uxPdIET3Uft53qzoSaUTyUyL5ZnCu1Dkv3SzISqzI40xK8OLu1LWQOV4qvJexhVC
L0EDl6gKyzKFzi2AlHTabM6xvjLxtYf1TxScp6yn04k9cV5M9Jhybi7WAo1VQO1G
Fdsg3C5BxYn4+ugPORpF+gQ2OtqzuF+UlNCahpOKW+tvL5S96A9RH/G/MagGR/7u
dfuPBCS6FN1h4ckxL3ojSus6Qeg1nkL+/JjY316dwE2CMpIH1aqEOtHrt95jj1X3
OCybPdpWqvY+tAFn1ZXU3sqHjRImHMmW3y4bAZx4gGcJNasDtO8WPATxJ6PIoxzj
ZewYi8u/G1tWQqLYBZtmAsHnNsunBleUs/38KDWLiCrNrJI3GckxirMRx5toWiEi
tv7Xy99hzN6KJ0VwXS6YY9HkW8uqor/q5J8lP9cGkMd3yGUsjaUGfUn0R53DRysP
EoFturRYnGUusQUSGb3cM2V8fdGVu9U+TzvWhMZo2Y8mS5yV1eS5jaJ/h7Q9DOOt
gVJYHtHjgOu0mIxXr5ZajQbIQaHaQPiUp2QRW2JpOPrfDCCRxp+ha3Ic6evnvkvj
xhjEHrSeB/REhXtOhl+CYEfH/BdKczzb67PMP+RkyxriagYcjGKsao4LCYsTV8FX
ooAhBD0vqbr1CUsBGm6IVsMzPb+Ah2bqxe7TaHxHwiABu4zTZvb5KUd3p1mMmSop
Mnnpv3sFECQSiOnShHZ4kCnistv00mLCB3zaLffyIA2QsJe7067IOwbvEweMXrz/
3KOVEDDUqx4WGjRpbE2NNDDSdWG9HRX4lV59NdQpHeICgHHe1WESFZHoTuq4KlbZ
rqQPE7cFLLCC67JRBieQ+GtBLAPCMBFRVFWV54WQzgLcfrVyOs3kQ7Luo+0ynVo/
ixTTeo/5j5LIbxOEYmpGpsJvjC97VxRGLRFwYs/BaE+0AzShbCBY3cZ/r7Z8P1B2
EdYtwLnxXX7kfOOsiNqe2MzM6DSwRJOVUvAt/zsvcQ/PpxyQ/dlgFqrohtdx13F6
yhELvdu4JI9BqSq3hpaXCb5tpXImy3ZMEBgIoVAa3+wqCDxN40mpt4zcQZvcxYW4
1Ja6wjRrxnxS+PdxVoJV2BMIDSubS3LAXdroDYEkFJfQtFVqpID3ye019U5zQ2G/
hoJERJCpSZKVuDEYrhdYMuhu0x6W9sJ+CAHEwMoo7FmRzv0cGqwFnhNUOMdSSgb2
izkCS4pqt7T7ChHzOOtGTmKujI2c1DH8n7fG8YuUMC+mcHtg6BwrQGBqfZRR5FkY
fkBnSgJGpxufd5j4jZRoF9h88mUhQINIiXX9a+J36T57i3B5vUmlzMpLjVXxZVZF
9FragW7PEBrTOTOXeGvKZrQKhnjynEL1D+ZgQB0KO8UD0hV6SnokMwn0pL5o6cZO
a3yEC+H/3WmbYurkfcSJ79HhPBYaHb/mkpcqcArjz6DDHUPXtYUzV49P3Mu2cb/f
7NlEn0cWiIoaEFe8ZpQ/BVbXhdC62RsmfHnqe1dvG9BtoV9c5BJMUMZJnwMB/23P
wG+LBR9fMfYUNIZbZBetFO1x8BMfwxSiaACwSRefG4g/sEE5DHWCMjQYNTDLDtWH
FGF5vxjiElM4YI/ZB0Rohxk6tsSaMnTgAECev3+U83SOUmNoU8Cru2yI32GkDyFF
WqPhZRx2m4sExkj04qwE41bXI/JIuwZjexTUBO9UxolM5XuIglK7OQ8EheUAzA/E
kmxV4TEEli/KKdyoy243Q24TZy6JWkISY48LzmKmqTYWgy+W05MSQ91oDcpHqBOR
5ZaYqGMyq0eRohA+CeNTSqbvORUyCTwQC+AW2Ve4tqSa/VSILDRVf/OZHd/nCJMf
0XXPrWhYJXZ35MWxjk7b/gBfcmQPMIZf39Tpy0vukAslNauhoDbsJAkojEzWtaOB
IUxXy95bfdMSEew9iyfRYkLMwYsNpWUuAhywno8UsF2NOFyHPVpB5X/3NnH9Mi4Y
JTZRfL/hBNcdHQPodMz2jyRt5xV3tgRFzl2qmLnsXQ9indrFenFr0VpCESJAfR0C
fFLuyou61cdXpL+jKZIV+bWCWpDdzM3t1OkkNeddBzvd3R5zEEpRI5eqS+rSiBWd
TpD7Qs13HArCSvJY6Mv6Y5RI1K+UWLeRp5Ej8RPHBsuRtmy0xGFJBRfX8jt5V7hM
2KwR9QN+c4ByaKRKSia0RzEHd8wqCCG8vpEQkMNnkyygrDYPui8IfqKgDQoJwyVL
5fQc/1PtXDiVq2OFwGx9DmrIn+gZ/jPF94ZVZW3aMdQS8l7ezwKpMR68w2KZVhwJ
pPpCnaBNxqX5JGsnMqWeshxyYwBDm1RDHjTprUdcCGteXlMr5zy5uKGqhprGCq6p
47o2IruCmmTACUHfK3eJkBgIglT7ZafETj/sWV7HSNvLVRHIkG26WuEXTbM959HI
u7mOi014mxSulamfxuB73X9AkojPVIU0+hsKVeDqoejkTjpKwqFD9Ct0YKdbSQAb
2sSl0rLFwQPpA9c29K/KpUARp9ZjtuJ+KUxLC0PtVI+i5P5/CfE3hd1ZqlJUUW70
RmDiBmkfxSy4UCmlt/ZcWOe7KqG/o2Yb3nrf1avrUpPafi0c/BtB2w2GIa8ek3XW
bjdmddEnzqcA5d0WlWvwMPhcgNQDVbcqJ3U5jBGMGBdOQs//YejKtB1HRqdkNiV6
o7u8vhvT/6kOKhkyoM7SZav/4nS0oivlAyssofhq4kCgIYBdxm496QT2N5HVCenV
2YC8zjt+bCFC8NqciHd9tVyJ+bCnl7IEkR6FyGk8lDm52eF14KAvrRoWMXNsWfDg
0eIDnLyDtS6Ze5R2/0A4FPcGZiyeNeBguQGzPOKWEYPCquM2lm8crP6smXAav3do
QQCUyDTk5igOLAcqdBCKVuiyDlBcIZcLzwgHkNi+eSM4ad4EbDZd7znJkehhVjw3
FMTaQHnrUotijhMsGo68L7S+Ddg9UKttSvNPmdzmjaRV/y15AKjrSQFyy0O9007L
JWXztRQYDjfad6m8pLwRxTVmxxij5/RO8YN7EOmrNjUHSd/w9PI27VArCvW4mWMV
14iDjhRTdEHTym9+NWfVITD4EJCpjAltTlaj146FRZBCKzI8blnxKxu0/iMpVrz5
PyrSc4zKiqAiRNK6+bha6AJ1E5F9zyDgzDJYdop5IwW4QCBCxRX5cXXTX434l4CV
UWklkPF9QMt3j7QWFug8j0rSX/zXUfAwYdjIdNMw8O85at2XKM0lyzG8eE/nK5nQ
Ow0EoB0dC1UHcEQsiZ1IysZi8qX1LBhxUS61GZ/QxGA+e58IuQVCqe7lo+qOUEPZ
NY1PxFCN7N/v2coMVOkOcZbMcC608gcyoh0XJrWvykintod/kp+MxBsbWfyGOxDb
7pfedHaHgNLyrLwezt8UmuQH0fifHwpzEJhnZyW0ZpcYEaluYkioJNR1lgZDVH05
tGvhGoNXlPpcFzgc9xSORu+a4bdcM7CUojbtgBVTl7Yicb+HYQFoDbAZ3rQFzl4L
M+nxZQyWo65ZTraFeXn3CBV1anq45UYTHQ27RkgBGqX1y5Etj1tty5gZ4WCnsgzf
Iz3wICHI1SbhIzUGWV0fExd25+N1ZZ/Ov8DsZqWp3Hp3jfNG57WrsVKWuoPgQAx+
8e8PcKE1znkiEFFPjumOtWFR8NuExgnIJh/O0Yw2WdO1Ehp9QrOmWCCbExRhP4BL
rk4/Ojag7FYNqgWf/Ph+U6Ekhv4mghlXEmZvPoqpS/wmrY5Hj2KiqGK6SJp6lann
B/EiGHcawDv1UFVxkRVwmK78LAATwZHjWXk4UPwidI3vEm/nf82les/o3BrXL9R1
hsxZepFA6zGY8wj8WXANH67oO7QEKcTJ6D2Zr0yckC6dlp53SzOmEPA5qdnIkoSY
wL9gMvkY7MJ2L149CXH6UFmlRNmU4gQfzc0a51L/IoU7PrFAFneeEr0j0+nPFwrU
YP7HKJP+4Su7CBPTdcnbpmBW3ubBAGtp6ugWUSDAT+xY3xwYNqfJmQBPROGanxVL
P9PVImU8kLhZRE8JQMRGsxu8ap+Rh8DrlRkxg96TJek/gCKCrnH6PG1sMCRfj6c0
a6UMyv0oKXwRG9qhJ5fEGdeD+cccd+Xs5xRNW6mr5vbGDLzH9QU/bmLXzAdywZSU
Sc4HSr5Pe6cEzGVzV+9SwPLjbhTIKNSwCjabitGcZK9qHf16iydpWb3491GlYhvT
6ToU/3PFl9TTOyxFnW+TmWrmpmmN9JgP0FEHGBPyOio4f3H7SZMF8OGsW1wIzv+z
+yR5T0Vdw6DO5dpMAYrZYOlAUZgYLvSbP6F7lu56uIsVGF0Ku+v4Cm7o8hctoQuP
kCZZO/ywsosyquB4UkqMBRRbVNyjjIlPkGppa/bLa7wOvXxYnipo5fL7to4I6XCb
lF40hx07KF5gQsv8G75gPk4QD31iHyHmJeAUvrgWE67rePWZlnEz6vsSlccjeOpg
RWfZ9W0HIHhQWDET/kGIwpobj1fJo8Xxl79dPsjA6mnFyUiFhSYLpz6DFldpibzW
SZ+UFJtnpK+E8EzHbfYqr7azfZT21pnKMTf3APCtWxrP9aXIHltuPo7s7Fd03bGw
IYw5iVhYwNDaRJxe3Y/KaV1ZA1SQvTPpNHZZ8ne0eJLNUCE2uOlkQiFMkgbzj+g2
vHZmM7h6gAyYtwlfNxgg+BFjuxKjjZgiYDaxmI+fIx/bWcZvFQcHIkQf+mLkXcyq
rEAqueT7mmz5WgOUV8pCsEGAzL8wasudck4KX2N02cSTkFnRsAf8T6PjYcgdMSQe
iSRQjEpPWyMzt8aNMSMcEWBcOgOlZI8DLKWw3u2eOXopP++M+S3kSxEh6wlTTtHf
uSMfWjUUL+GMoO6x9V6RaCXtTSK5YjCfciIzrTN+DA8AzpSzqs+om9riz3bGI9Ro
mCpX1W9Wxlqni7YFY039O2Fhxtmq9gXCXYsiW5QLPg6N6ACmwKVbPZRmTA7AteDr
j4efoWnJJdqEwvnoXwdUE2bqEtjicbi+GL2WF9VqdzNf+Ap5XCOaPU+JPKDZlmSx
E0SmvcBrllVXynUKRGVY7QaymKdVec8RIPke1yeSKCWyddXFBAOYPlG1ar/b0hXh
xM3gDN3qdsjav2UVmm9Lm4BTfRfHCxy/GKB8O49ylkARXWygOd2HSpunLxszYjdp
/KncmDo3x3eoV3Fj6jwSipZhHTHBynRKDdHkZ70Tjo4NZZgS5zpK6QopoItDmKB5
Kkk2OJLg47f1AhhwXOyAOQu9bJ7q07kw0SjV+yKSTAoN4Uw+xjLCzcTOy7NjUlbn
awoMN7KNb7Ez7RNyrym2FrSPXjPolUNtz8YKBi7d7C8PsreO2mjJkDUk5cL+/7zY
/Afztbg+VVjXH7FapTGxSDQZClx+a4p0ciJ2TZvMSgrMq5jxR8we0jHO7/O85XHX
6B10FhO1KZivvJMaZI/EaKtuH137X/xrHXBGV7B957k0qhbYzX/E6nhaYNnlYr+a
eI1ap1w9b3ODr2BChuBejzDcQRgADfgEYU2W4asHJEVnqU+aGQFrOgeOp4cGpdsQ
cLRXVBnmMs+Jfq/Ucp6HFe1Qfp46j+Cuf1h73viWiKs2DVjuMoLc6KFaGw+BOf/E
Wg23hSt1Z0q/6jl5mjkzvyVN6ewIKvW7iJtZduqTgmyY39bl9fdDsxY7vzOcsCtN
nWJVa9kNGKHssvbNVH1YJ5TVrlUq96Fm+85y1GX+Dz5FtRFPGgDjQgtw+LnJCJQP
R5dAs1YV9x9DtXP5aLW+N7LbMK244UhYzNFAgpvtsLzVJu3nAJ+jAiuB69hW6i8E
vCz1sqYsrhyOGAfxPuAe76kisdsWCLT23EvZ+Lu08VxiCyhZnuj3MRmmk9tK9mxC
R1R1bJPXWYUlVfaVTh2zQyhS/hTFogLQlLmRs9eRF/zOHsPV9IMD1W9PXLI2AcV4
veSElqqmwkBWeO5pKghv8zvnFjjpQIeyj+vXkuPPfcUnErQoZn7/o9tR3poPM3y+
J02wc4X8K9Cbl/vE3auo6fSF06TvUrsSjzov1uJPcUnRdPQk+yH2o3Vj+IKThjMZ
zFTpQfwUM80BplJ1IkL8ITTg7u240ym7vSgrMFs8xCD0LjyDnAKz2m1D4PSiQI1Z
WBcjq2TKtQH/DEq/dTmoZBu3JvodjWzRQn1pGtcc4OAncbpvdEaqypwr32wwEPaY
U0znbZlquy08tpWXvg+YhPPiXksuu+iopT3mEflLqTvVDh1i7S5hsZdoj7NYoavH
yC8MYfFesbhn8E446cf8fvZGiWXGENf8DTvJCTsB0sxQ5bv9dsc35rSc2qu0HHpQ
lvZRn/7sdtPT3aoqT+Xav1msiDBILZ201sy7YHvu1Wt7DNLSYsBlo1Qn5WeAFlAf
9vcoYbk7KonbQYRFZHMl2TPtjNsGtlRHiZhq949d6YNPs2huG2nUiLbBhm/oSlAC
awe91mi2fkCmU+Cea2u8wtfRKgSQ16FiXC7YlEPizBlPy5YzciWZpFIBCM3vtZHs
FbW4uisecih1i9LXSrpfpahQo/SLcXXZyKsk6rn3mkwgnBu/5dB8etWgt55N9xLr
zO7DnT25EGOeAtK1zA+/i9sktKcXEFoquT1xf2DMyJ0FqJaRLin1j5sXbU3Zvug1
3b8jY3cMdldOj1/X+VyBhmljGjckJ1w1Hbq2Li0d9k/3rVitq+jhqj++uZ9MomM0
EBjDB1/f6HOUJDcxpQXhr7Q+8r2UG9RUwxNoJ91VXSCaN9m6pU+yuanIeQhIbs/0
fMUvRHQCZaUDechV9qZQl27WGmr6N05LDaL/XSw1rPTnyOu8paDE0VdK9CPRGVlu
nH4CSDueTYLiMw3MyGDjE1mTA3qTleEH/+a3XfTMl39R1aohM+lT0Of53aFKquDC
JgzYpTy1pe8tk0/8U24Hq66rX/pgVhm+0YCWUUmv+gfuKxAA6H3QtAOUU0skSBbZ
0L2GJiNGm79SHERxVH1sloHMnVED7YQmbgSaHUXhTAbGDZuuyJnVD4NGIPzGtMSh
PCtkwp+hFSRXUsU5T+cq5aMLXLWmLyQNzWmFzwVq7v/bfqsBwq+ugF0Irc47eAoH
JobqPW9mG21Q8Nf2xeYcpbXAY8MBn1XKQYegv6YAdPYNoGyZM1wtb3i2ALJPWahK
QAdzpR0DpUt4/I21OVzQ7k59i09cmav1bKDMb5t/BupXBFsYJ8+5699/hD1273QZ
KWEX9w+OVOw1XoA1U+wHk9rIPdEVq0lMOGPazUGLIDldrZwyjyLg1Y5IshZmEWHF
DaM86Wzc6N+FZ4+kEC2uh2xV2eAq9OEW+thEvrbeK9wB6SvNrjNyRCe7iefaVsf7
brri3NfA2inF56RXwHJ0k3jS7DFTLXqVmvUnuAAa6GaVkwYKzO3YKAX1b2kGpqCJ
apsmxPquA7A/eCF3QSob66sskUX+DauAx5d8fzKiXOoITkHJihume8irpWS1HsMg
dgWf++c9te1XvTMuZQtxYMxQEcM3jiHOORYByj/0RO1kM+OY0RQo+rqPVujOkZgg
64ICw8X80gUKIK3EHq44VT1Op0wEhNeMRhtYRDsNC5BxpHF8KWlZNMc3Ohwr9X2P
adSLzRhi4dGT3VN101gLUvYwa9plAK8278jwnC5aPpt9UOWLbIbm3DPh9oysomOv
UYU/cs7RhFyc7M+OqmrQmA7+mmJPME8j6DnkFsZhcoTbV1AenCiPcHj3LnbgmjEv
pLtk6+iC/mCXpo7k6YJKAfmLYSde25iZSbhaRkn7RN/UCWV/8Ot/hq/A0W9wfr1J
/cTxESsBbteOmzVs0l74iawGHMwSsDD5rEh0t4BKsEH+SX5RFFFOxAmTBLapaVam
XBIMB0Du7ycaY7TtL2yCpVKsBbaf+3dyEfp67KyIftdWVM1uNGYnc5AChk/HLBrR
XmnHgNyISRNLQ7WJTFgAE5rG6t1Jq75i6mpVVZQNW/t0S30ejQhaOYFWWMCM6Vj4
t5/obHZXmEbLx9lKuHCqkwp1JViZUMSSiddfbKerCDzvcTYLe5wtvh+yilScxobZ
LdTD9fCEZXe7LdgCE1na/qjxNZfuuchEBbbjRpA7ZRGnzyaGEYTJ0zsQ02WstNbS
9HDd/WK6pPJii+ifzAy8rD383z30k3HjZ36xBg62k2DftRhdkrrtR9Fx0Hflisdg
xrieMufxlNmLg5FnKm27CkpVuQTrX9VOSdFEm5OAY/UfrlsM9f2dgOQwoBUCZsMm
AIVrcfo7u3wbCljBp2oGQIguWJ7B1lNP5EVSRNjz1RgmuH9YQMG/v4T85KW6KJHv
atzRb82917ffOqwU8+VwYbIjzo8PVD2LAXVTPQztzjZgi4zc7Gedwe7ufJVbuevv
z9ATQV5fKATa3vnHpbtNA/fNMWBGMnSQz2ZHPjpHCSafpNxa0Dj6d8+i+HVr9Qzh
4HGf3Hncyglv0EQpsQFjkOvo+DlmMBKHt70oNjt4hh9j6x0MA4xkL9Lb8H92Bqqr
WdvUNA+dIgmH8nc6+q4kRweLVUw1zs/rpum2aycB8N2lxBhLUrwdmxusWqXcZ6Bj
jr6SobK2Lp7LDtmPXrJCbayD1qJZQPu3m5dt082FyTkaD71SFT1u8YKFMTywSZf5
KYwbEbb8DQjJsO8H5E9tZgl6guQHxdpTChOLsDZVcoQZDQtI1kDV9Nmi0Gu3x36n
n7EiVSFFj0dFTKXiu0Qi8JIjzKvy1PVDjXfMs4nfg4v8rzGYMtGtkhPOcRpTkeb8
I1PR9JDf5atWy8YOIao6Iv6p8ph7U5OlSgBz4wgjJRyLJRdUvPJUVMaOHpxzUits
iS19Y3lF8OSj0q8O8KHUFhcI3MulZVDVwWYlXSz3d54+urURH/eq2nUBL1FfH+70
VruhyfYkEpAbRCfOYL3uWl6jnghHKovgzaImmzrw2CqToq2dX3jhmTHtEpyzDmQa
vfzA/6FTJD/2IOuTBKrI8ED9GjjxcuRAZmqhNLLAMIL9P5SIiF572U/RzUsltMs8
uGQ3MyRi9Md3v9DFd8C1WCW1FDdLyQnWbnBhyXem6HBGRhQLYGI827n+pc2Hf6VR
CgmmFxFwZK+FLqeCHlKWKOzfRJf72zBC7PTYc2qWrK46gOl9KDMybLCRPDllsKsS
75j/yXEL0zAE5jhgbYZOVi2kHz18wvjRFdTAMgye0Uq4Z2/U13V0AqJDfxEqqH9u
sd6p6K5wmU0F6OTXrj2VDZDfBGk1eSX7ElRr4QOXPXYsepoXq6R3+ynXq8pWlS4T
WcmoWZ2N7AyG2iMl+oyagoWwRA2lHeyxFUDeU59sxRGmZ1F5Ff0hemxExZYId2KF
8RvquKvkgzzrBYZup2A7pa7HB0ReVBSsmpFm1Oei29/zivkU3kZX+a3CzBRBwyaS
+dpowFAaCaCVvv3s4iBexYAJWwlKp8gJZJWetNB2glOWh0PnIKnRRAahGqx5zgKz
JLMgTJDBkl7BEl7GHit0dHxoyB5A1EbVPBh+yzLOUJgBzlalbHTM0s05OyC+Eqg1
t75XgbdpINpwK0j80ReaJzbosIYosdl7dlsF+v3TH3oq5I+x3spaOSZ4Ve9lcqO5
f7AM8YD5hEvp/SCi4bZa57vFWEzy+sMfIzbV4aPd36mqDUXS1DCClv1V9+5cJqaA
rrHx/yuMEMX7zkyF3i9JYlMlvHoSbh2sB9vIoGUuLmenXXOLfXQ34fDR39QpkzyB
n+98jxF8CdLJp+I4ghVY3lUDaOn5defdKQlapVeeAN/y3zKPaR3l2UCPiV1EeVBY
trcufLaRwKTos+2UFYSuw+KNQkh841bYL9F8YytawGW4UpcvfbqC6QsvO9/Y3Aab
T+aOCDgacNWs4uqKCa4Xwwzn5Cuc/6u0VhV0Ph1U4SkF1RUbunT1yUyKDl5NtjbX
tBrDkG7wnVrtCrK3OcTB27X7PpOKI874wFdlc90sTMr1mAekmnDp/AK4ndLk0Nq+
nwymFQertVFc+gZiZLCeroIx8o8vo6ji1ejscCiJDhXYiinV7eBXI7TYOeISlmai
c8Jd7sWlOD+CZbI+xwGeI/kwD3n5uYaBD1Y1vf2S06kqGWMsXyvRLiDbflgei6dk
tXkFS/N1xMf0cE7cSIUaf2Q4OrKE/93yv1I5U7TflKbxlleIV68yHMG9NvHZylig
Y+B6LB5ScemcRaIbGX1M4yGHRw611zgkqhy/KunesXnxxGrL2B9GbNH3gLSt9zWO
4A0Nfnbqbj2m6HHJym1tYsZYDVMtTr7z1jg5uOeBZDOh57RQZNLM6cJb40XlmBlk
p4JSYxGwgjMcnP9G+9udRkLiAMCgPD+fzjcRNUtH3ltdvCpDTSQVuzUavKDbn60K
V+Eugbgo/R0jZV8lyKj8wOSAkV7uUk0bRkqor2ob6W2bmEd7NKMGt2veIGgTC+V0
LbLjeMtsm/GLU25oUG7fdptQEptLqkWg0enZ117G6bRvgcGGz9Slz5Dptff0hg6X
84AdrQFKtyT6IL6m273Uw1QYN6+HG2urXvzZLvRrPTUQ6ziMSXms5cioOk06krbp
4xEKUuT6m2iaxDtfJxAUTJyXVeb5UwGEHAWCZkHZh3MIExzJuRl7ia2c1IlbOQ2D
G5UGWXbR7h+d2hKF2FXqNo6Mi+5s5K8eCvff94Am5xlPv2NwIASQRM2Y1jGGwIs8
qG2SPYFcZahAqenPT08+1VipI/fhx8k3fJ/0+wEc+WC8nyAi+3AniDrnH9eMkCey
W76RYDxdiY/umn/Y5APVkMbcFxxc6phjYcD0VlgEpWYkU8f02qkoT3RdJpcZEa01
fWDfNtBxDilOPauohIw6ALddnYvA2YZqhROCleN3LXykcU+eaw5PeHfEfxlsY664
UssCo8dLArpepGAiMGFSUkTfRqo+BZK+JISgdGUGCLKFsnBFTn8KETCmP/2/gOWj
Or3CaECIKKKMvShJLl2pw83JIM3RS7iJI+19TTM8B9/SQ2JEPQJHYrlVlhlSXj62
kLAVtpGZZiP8ZCIW3/8pP4X7R1z9ZgZLKS72YrXjCAf9nv0ZfntH/kdI4OCbC7Bg
ZCSNKXzlhAyS/WzdUh+5gDNqosmGvl0gpKxM9dYUBU1Ll1tS7+7ZclNqsIekPOSI
+vY5vUDrCTRxbktttxmcxwdObhVUEVgRwsVA5MTQDIZ5+mUGkcO+ozslahqDYbO5
UsqabfzxRc+GVSKhw4GyQboKmk21QGXW+2HxqnCPi0fVOVa8oo+nkLugNLeSi8aD
nw7YIbBhnQAebsqTi3pMA/NckvuCH4G76YV+SIwhiCSMtA/JDenPj/996mE+ruW3
iodqK0EHreSP/YaGfzxGK2n3rA2g+8jCqW3ybfl79Ig43aV1yd8lGEg1wXjEqeSu
VxTraOyElzUI8w1CdEjWx5yAPEHnQtNgkL8x+d4cs+WD3A0KKSwCc4xzTX9KJ4hT
8v2t2VXGKYzc/egd1AHKHJhfb/z6UXJMWmAnMU2H0ZRzGOPWDkTF2Su6lU3P/DCQ
ZN6dW5Zx17VdbjvAjthC/8kaPX3TDMfHNqn6nKfY7wyBOC9U7iY0ucwyi7eFRAFE
hVIXVDIVVSYSlv6pFio68vNJ6u1ypZbyPgiL4EIR4stjpnxCqTgAL9yFMNY5MhW3
myjeYCpiQjcz6E1AKo7Qy4R5bpQ8EI6+Rz8ghDMk3TUPyhtH8Hlb19W+Hw4NEoLz
PfaIbCq7Htd/JRZpE20mucRNIjQqGXIgHie/jwCf3f7Foo70fQEdMX86XJ9YGdtg
zMr+hTl+6LM0XNs3iAd6FjIZIQW0v1bE7bWlHwqfTGQC5P24rP4sQZXxEV3qjEmv
wltLb/oV5pklRXp0N94TrKSC/4+ARuS31iCPhe0p2FH1MgguBMTvCwyMbsK5EX6r
6tvTwauzeD237pqf/x5XcPPG2SX8xUXkEX3z5hu6fMSSChz7Z2ZIy5maa76pp8bZ
NMu56EjsIHw2xgI1H87mJl0MqqDbaTd/5LAVe7bH22Rk5xEvMKZ5vHA6/c8F51AX
20iPk8NwlP5s7E1K8HKxtzepbSyBnRycgxS/J5o2n1y+TPSf8MyubBIjLU9UUxKM
EZOxou1fyItKSQRBnLo86XKLuMRuKLFnYDTZQcKtTviJ8Lc269luB6s8WgvF/p8F
LkLGW1XS3sMoIG6rA/ktET8tYgDsCRagaqHJzlNEY2PkTK+Gxa19bZih7dMDp/cS
ci22ni3qgy+XeXFdgrtOB52pRsNzIbeMaGaWHUoZvhfaP7yuX3hDsyzwWRQ4mtrt
8zpQdznDK7m/t+8vSfsfzw8WQav+amIFW23NvudaGIhXUkJMdkK9ne6Jt66SPWSA
6GOw/R77nVcL6vhuG5BDF9UnUGFbgj07qRZTj+huLwyYEYkWQgPSyn11oY7nJI5c
lsJKkxuN7SLAFQJqOHStvu9N3ySEz0R4emVa0Ksz25tn8MBdE0Lo5nXNehL/21tO
OHN2OwIpRBsNjNktGjSDJXXX/WAVZMF0WF4GB33t7ub1/PQqDOs7MtypfBgokPxN
JqKX0uxeKKJOm+QwxVWvOqtZ7QX1cwFboEKvA4XwIMwy7DxCDKNQeUd1Enh7kJxI
Cl1tHS0Q65mDcE0yWy7akZXVpNeKzBCuuem8ypz5dXlVxULuxx4WlH0f82+q8ieF
K6DUi2m9jwWrOXApTRzTB2YZartNw9bn8/SAxxIsdichRxsYNn8XwUhdWjwkHCcY
b8AA07ZUlXTFYvZT9LXe+k0B1z9rUMB48EvGgW+DuZTmRNJ1Io7StPkyq1DQbw37
ZtKIw+1CGxx+lzpEaqVudxvk34j8ID2DV+OY17xG5aSFG32+ilOxVm2mj/t1PUZ6
yZZjOxF4r3FA/gdaLvsGpXDptny964qzp/NNKYMSQ4WI08TInKmeTiuLatwRxqYJ
T1UwbKLQ+MYxFJsZggqpRJ4IqnJTgtyJ6dTtUr9y9UD865pelsh8akhmgVdmaywg
SX0NonUf/HlWP5jlqugGe0lA4amSJIjOqjsWuEx0GN/5M4arObc1uJyxIUJmTSZw
Lz+2b+4KcNFtH5lUbFrBF6puBKz7nMxmg+VHGz/H7D3WQ7h5dowO+moQGYHnZf2p
vJABhjkNoZvKTBR4HSecdERLNdOLPVOqIRBJCqZftc9L9X8ron1UAhlR2tn9qQbq
HX+5+vTeDyVcuhEO0ltuYDKKGZ3PsPQ4UpXPF6e+VZhpxxD+l80It29cKV0sz8/J
jbLjALkqQpZnGm8wL6dOS4Qs4W5CO5gul+yE7FQCDQklCsHIn9hpkzJqG1ENoNEL
LmBPK4Lb6/1+9pl3iE940Z4JiRYmqix1/A0CV++6N+EkAbymag/xZIx1S55KENVb
SeRHbN6NWKPXDOCtX54ck7n9/SX9FRI5mztjR6RLdTc5B4YHyeeT99yJxOXaHC+K
RTOw7NTz90kRxmFd8FKkMHC59tjHZK9btfbk7GrtMuhT5xWA1ER8EFlAPRNZDiMF
12fRncifKL/hjuGho2coBxL/IKMHt0QWvoOErhPXY07UB43yU+3+nLctKcrq5tqT
QJWuJB6r9C8qEbTQVIP601G2OooRM2HWuwEYGYxW8TeHZ5K1zmVxfmCR55/aPAjX
6LDhQr0C8OV4loAxp3BMz2GYYNnA6g+nkiuzNmtPGiwuamgo7XCgZ/Lc2qDs7PRy
131gA5F8mIlomVVEk0quLR82ISQ6Qby6VPc09t6LT5kG1m3iB6X4NUYXmc68qg2z
jpP4VX6Bvy4O97kwyzQAY7dfilypeLjvp+NVi2/mGE1DEjpYzLcartNhmDL2oSSq
legd5VDXqtFM7aCGtvL56g8jaRVNuW8u9Clvwzs+dfGFctGnzDoedeUrsHqB02Nh
CB+p9MgW+qCCY19FDQ2yJlpTLQ7Kttb0Z6qivFeuIZXlI9gh2jX/8dJ+cuygS4ct
U8Z34+yJfizOj+sWYLp6OwpHqUkkvbJSUFJoQzC0tAL+4fQM6XyRr28YjRdbY5IG
L5Vu5+DqLJvpjBW4EdOUKxLN9Qx9LS7/SattIZoslabs1sdbnX+UcRdIbi7nXKZM
G4fpibXReCmmHut5aKa1m8Odrdu8bLrpeoTLYKvrwpDAIFkEVzLCFFrWWOo+psnA
qI/MxqSnYTWD8qWxCL7czz+FhkIKkZphzeGl5IuysXyHZaNYuz1B1eer0bftoxzt
FSBDSG7rhfnT09rrMB5GOQsRJm066ye9t2CuEeNXn6ptO6+wUpsaV79bab0j1n7z
7YK9nM2kgT1ADQM8sNnVBuJ7+Vuc9gAuy5wAhcmz9lv2Ldh55qmrMsrxjMpss3S8
ri8cED9OvNmQj/t58mSY+f0ocYmpWfQ5YJ8uApOOvdbZIuTdm+c05GDAnMuJgi4M
5WVDjqz0nf2+XlUGfoIonP3gnRPtpCsqq25ZWCxu0DFn1R5kFP67CKPl0AwdeyHX
3xxMCfiPRWsAf8kLt5ARxb/mxAeN3aX8DFd83GpRvTbR5f5Yanfg4AMH8zVpNPdi
vd9wK93w0D7HASQEYOOFzNQlOKgybhIZ2I76VEX4ukjXIx6zjOo4XGH2ql8MKbMG
tt5WEARbViJwORO2YN1tfhLVWkIGvWej3BDVCrah00108gBdsGLl954SNk7meMQY
AdN3QWk1moCPwMGCfEDxJatHwL4LP/PxlVy/QDT8tflKsu/Kj9O/RDAyf07M9hUT
veEvlwqw+NLjIZnU8MsodxC2aHsH93A32khHyNdP+ciYJM6X/A1Fl1pFFN7tOgIS
Iizuh4JXEN2dpG6L5YiKeA2u6PRgZqbyz0HyYl4yPZbSL+zNN5A9lBXIM2JxxSet
56pHi9efEZOKAu4XDaQi9I+PkemKPnOQus+B7OeNoK3BEl9ciH1ymeryQMpEtnbY
I/H5PlDdPuyVU1aqsReGJGGb/wnhxXUIA1R/aoMef+qGEjXDU95Nifx5Aqk36Quh
0WY8FhQiId3k5lrG+sWw1s5qYG7R3ARi7b58hjrCN0EHfLs/vkeXmQYptQIywzs4
jEHexZw3B4RhMfbn+kOY8pUzSICHOVSHuzVeoTIBzBmbeSpB8cYbJo4iau8IzZib
YKfJ/6eujcb3E8NpwreVTf7SCcr6H8Hc5vZ0rqwL/KAzc4xUON97N5Hwcn8E6XOB
qJnLCOmBK1hnwPNM/ncd/zaC646tnwh3DvEF7M+QOQXo0Lz4/Vbn5v9w5DDw7vBl
fp9qfWYsY+ByWpURBBUO94dqeao9RcZKJ4sBjFGz6478GgxyBCZ8saQ/gi2PiiTN
7GsvFSQaJjIjKmG4JRjqzlEvG826Qq28/AdV7O4jHJrHOEYt1e2L1OTKH3egWxwP
rAMPwDWUADWJSmg70OkdUPDOOsvwbClS7hvgbITndTiKKJxH0zCnfDeHvR4Pu7S1
q1JPqJ/8VapsBeKn3NfbstCu0tfTeaWV5Ga1HNlFyP2QgO6XEcJ3wC25GpSeAW/l
O0syjcEeNZS6QK7zJGnk+J1ZI1GHUun3KXqt9iTG5XGJQ4qNXWdqv6weA7d6/rqp
WQgv7daECHoz8VoG98W3M4Qzvzr1QvzOwKrBJVEoyrPxT1s67wLAOkalHX29Maof
/e5pnI14pWz5x6GXwDaUXlJ+PTsalt1bbdalzkbMkn0PQAKdGc4vGLOmdHwgLR1z
3ZsLWg/q7RtIu5m3UkAXeewf9Dd21HpuGoE7E9wi/DFAdd2qqSfhX1izQWQMkKS+
p/JLQGHPIdSx7BlDSVS+yddL8dn0iIUzMKopkcCAztkjd2/td9+oCgBEGJdGnp4r
x5scx9dhgugI0lq6hj/TBNPkHvmCIBLao2tgSkZ/3knuulJ2PobYyJnFRhFvXJoL
HwqORT/xfFmyGov7SF9wi+3vCQoMx4acxNisRoBoPm0/BN122gyukiiXD5BZAt3h
OZ8Ek7bII/4+ARrdafJE05r+ynaSOEDB9/81j07yZvzVWCmYw/wQTrMpPmfqwOLu
bUJVdOs+xZQqK8A+38WQ/WcqrJCrVre2Dd7qPODNNMNembindtqdw++USt4TiN6w
hwsyGeUYuws5XdVFSFw88wcRC3PGoaeb6CFj2NlWQZoHvIaq50ttB8Lglt8X2NzG
/JDpsO4CRGdcro8+5fILhsF/OV2MqoCwp1lUcIwgBYVjKt9CB2SyXmf4x3st952O
eZObMHE8QkS7hVH4O33KKNGeXmsaFt/fIrWI4Eq90l+nHRmHTbXxB2XjPhWaGJq7
D3DyeVpxuqRByU+rk4/Je9dAqE/LxJyTwZLVCYN5hzG2vHcyA6ScTGWxlVog9DAW
0U/mdx8+y2iKCYV5CAaa71WS3rG9+2M6PJn37l5GtLHUTLWCfxKeHsAPrlX8EfMb
JEKfMoHpVOaTNeLe1iSr+8os+CPjhmOgmrECZwNbwvJ6cFAr9Zm8kWAALiN57mqg
lSe4fcf2sJYJ434QGNtnbuUQoC1jirxAxghYNOv3gEio5ktzdpOenR4nu7ht/jVk
I/xQdVM26q7WssOB6LiUriGqGYTrqTPMyA1Yx4udolJmk/Pg5yhjnwSe6+R3iTL4
OL4Q5GNohhoUvRGMVHNeeQKdGIopevL7e/MlJjdJCpqfAKSpbjB9YUp68o7StgX0
44/97t2fafBIUu6bIprHWmBORi+W6JIHyapMwc1oFzvzuAX4evk/uD/ardL7Wn8E
CYMPfD3QRO7OCVTYNQMjIsyCsJSRFYxTZDyEyLeTY0z0SxZrA7n5G8LJxXJWqFW+
sFDdtev0PPOF9yvfXmVyf5t7Vf5e5eTI559/SEz8umVFKxgJKEGF4xR33/mWzpSQ
ZcecAzJXoBC3SsEPHyFEUkFZ82FE6jh8HR6m/vmZ3sUgvyGuNt+rXDfTuMHvSSgn
kCFPAVSmpudsAo2z0rOvK2PN4l47eL5Ak3HJ7rdfWTL+Ge2Y1ifW3cuDi+mBtzOb
aUix3G93L7lzw+57ttgEPnFAH1ozmU0UKcDpVn2SDF+mA3e8de5fIDx4aaQb/UfD
UNvbKccbiKIvtaqBKZ9AKh0epJVcb3W1z3lD0qOWIKpB2DCOT7/gZe4FXPnngIIt
AoGrEYeNHw9zzFuSrqUBknNWaGYSjZkp6E9Q+UtCqGkUzRwUfYqI1vNHSVXqjH8t
tNDXfqmzYQeI5AvPluTzHE8EzSkgTWpQ+GV69y3E8yjdWufayyOz2QX+w2p9Ph/P
5EKApOaE2Egm/LBkPDY8Muy3ncZjP10Dfq0bkKxcg1LbFsJ6aLLPIEi/H2+LwLsS
GoTNdYW12ExM+uJwYou5x5jQesgjpF2jpgHJt9hg2NDCNf+vFniTOjUHvNYj3MpW
kqneRHayCG6McNPSAX+azEtYGD86wlRANbgo6nvX4K9omztCcyhBFOn3GFj32zoh
qRrzx8QZmGM0z+cdKWTkIuMIVOobtShyCA2OqA7mrYh51xfi4idri52W+hQLLAfa
wAUw6rSavXsvqbv+cmsG1mDnNRHbdJcWpZXK/WzdZfWO1T3H2vYAvYUqRGsw7XPn
CX7FPLxN/yqmKvokWOLP0CGsxvZJg0YAbvy6y8cYQjx6Nzg0YTShqyufI11gkh7R
IkF+qeRmPh2KGSExsu9fQj195hTeHeEG6w9JP7S0tYwjINkvVVI6KRfITRzCeHV5
/RZV2H0KKz+CkBYntRRrjq2NgL+musRJZ6yrfqj9hHxmXfO+WieEdgCMEYxTpcXm
cqLjqJbsimrMwjLTd52z/brTqFENEkbY1dARfUBmFUKmzGLHY/GnVdPc4aqgSR/8
HoCOZcuGjbBUI6oI8hKmqjtrvIDW2hjXItnrw7WQDMMiYofDTYYZnWZeURnBlNC9
U4MwFyvZJmTvCLqgsVWg+xNLyrCpANIr7G+Bd5d/RzWHZ0UQ0O8IONwx1yzK897W
Rtzvw33f8gut9+xZPgC41a+Gl3suxsUeZmmAyYs2Q/KaoEWmTZVHEV087FQ/RAAW
5HUJZxtY7VmISWeZ19W2or/pU+Der8SMUROW+0J0F+N5wnFtcWsOzmBeWjKyS6Ge
PqOdjI/V1MUTmzOwVWSPCQmQS/C6wRGKTczE7z2Wv7plGzVio/443MKL91Yri9q8
L3J4kv9HEz3RfGckY1jlzA7/lwzEJ+dqhn9zJdG91Yo7VTxjX5FHKadwcBFb0JOl
QNiOcT7mjxcXQSL5Y75Svc3fO3MqK+nc1b874sv74pe3X1srzhq32dv2UaPmjzSg
7NCfUXSpQnR9lf3x349T1O8cx+vxzGHgFlUl257T/ADhVGKlB79eJs3g9szc7GwL
fyPIX8MGi7lB2mrDqC0V7xsKMI0w9uIodrWMu4cUyaLUXMFmVQYrzO8EJMrN33J4
nRBokAAfZRP/tuBNWJPhtPZaoZKhkj4V2vWZI3IO+ZQspxPn9aivBtmIkDekBTbI
pAWzr2yalRybmcdmiHD4u1DJE+FIGUNzG4GGA3vrzUkLCeOTUWN01rCnSV74ZV6J
Ik4KU1j6QTzuVJT2WWMiFyhvE5Qa5bKBoDCLrXNMakIIHe1z7a0h1KY9vU2llnp0
oCkyrgGGLdg+iHnX1lwRjY04uhxQ96MENfnu7VK4NL2Uavc4Nh8w5Ap85w71BJaV
HlYHPJqzd3vbN4uAhan1H8qGZoisYNaP2oWbZ0/s4iAKZcKfE3giTXCajLoZRpBj
hLcZljOabyAcIzRJTlc/GZDoX2TQnGE/PHlAUFBA1qdifZMLLbVU2WRAYzJYLJr4
pAUcwxhuEN4lvd4fdNxV6WQRnyxrni8ZxdJvIBKcWWpdLgy/+X6eJAO9Z+DKmfEE
g+li2LLfq/Hiw0MMPiBP+HZ9c/fryonOyXM2Y1foppzO0UsTleeVE10rJsjoEIEe
comEBjJcL5Sh8VDPiVZY9si11Mq3UZy4A1IXYBl0K/6kdJtgdMA80azM7Vrrby0j
cIqfdzhZewjRyMneSQ+grWluYo0nAaSoPTiaGOmZC3RUuyXMAFi7+ecAxWpiJebb
/oaHxYLtGRkbLz0GjYGvSqHugA3pE2ekwMngnqqyMTmaq8g9utuwxdQgH2jIISbx
PM+YOsmOahISxHTE8hAAkJbTbmFpmhr4IoPkVCJ9FJdIw9TIk7JvfVfw4pz2GRBo
yjpRTr35zTNtJ7zqX/qy8tZkn6RoC8V7G60euyNJoCFWbHrtTHa1FaCWdgimrphU
tTZxVtW+qB6UxuTG+AkJTZ3RkmccX1fSCt5AcBV3/vMcOTqKMZ6RT0gI3KLXGKqK
Pl8wa6LZr8sk8pBnu7cJX0YcFFW9NqJMU2Qo6vOwY2KYHEfqz2l8XbgGOUJvbXbt
/CK+B6TS9BgKtPjEA5CNYr786vGRakUmgiaLA/UIXo1jMboLfHJUd8KQGHu3AAE/
bna/Oeo1ZXpiFaJsnMKiJZ5JFZ/QwdpJa5hhNc0Ye8IpANZ9pOnDMBu5GIu6pVmV
oGFUvL0Yw303lJcjbjLjCY9ITtZmxPKPTdjZjtw47AnOifN5qAC3zy8QByQhKL4Q
4doewZbVWTyqnQUhrIsp71sLAqSZKeWSwtbNQl50Ggwkn5ds+y2RO7GS7itb1j0w
p0tFH87x6egYaZESjYxukby1mCQhonvZn6qc8RLliqPkmfC+zMVNXOKplCQ2GZKe
zA6TXDnF4tHZzYWxXUKAWAb/xq7qiPjT1WdJCZQFXTD85bq8lAkMtNjnJOgc2Z39
tBCrgoV162rudnRuYQjkQmfOriVgeCBXXhKHiFTkKEE3wNWJRwoQVy1s0L+gFIOd
ZkVzSJ64PW7ytd/0LRg9V6oM05ACJaPSciDHHuJl4/xxTLWTnm42xm+KB2Mlx+2a
vsop4OQmTRXxjxmWAW56b2cmE2rlUV1MK0Uiz3sdzZl93fax8kUO2VAeIcxWY4VR
rjaP86L6Qb+JErkzSBoHU/Phtsbze0IDQDE0JYDaG5kDI5p+pQMeKXFvjJ9qgm9K
dmqkrA1jJu/F6fPWA8DCdEaVCEwBiiQQ7kuVloHPpBjbf6hw0up7+pcYDvLdgxuC
e5tsgGosa7JOdNmsGmgAzT/TGqk7vNcSdcWS73oyg8HhUxBNtg8ZobuUvtmOZw8X
6ZGhjXxv4Z7Olr/o07ue4yA0TZMIRV6oD9SfHFLrLpTM4WeFxl/9NNegImb9vfWf
a61EbofOC3dI9Iny1DvkpYKzFJP6GgXcSs8k785d+djzK1kQtKzj9F67Qkh406c+
e8t10DyF5plx5IRjOObqzm0trH9b7M1ZUqoR1FfGZ2E8vgFYxJhkWjGUlueGTM3Q
nzuHnyzKzo1an6qdMpGn5RXofUAysTz0EImD2IxtKZwh3fGNipr1zMaVPwVFGEJP
1zHCUx80ng2FsHN0fCnuP6C65tdUULfPjdVP0X7g6CEPfiN5+fspdTTrAHrzVwnu
p4dPfOMNt7EQP7AMD4KIZnooYvpCnoxhlQhZxAsyRF6D3YO2Ho03/D6P8nmZfQg2
PxioIuj6zbMWhVLSjHXHcfBSYm/BzAjbxMyu+FZhinwGsFzl6g9JJjzFKtn22N7N
0CFK1sRkF6760Ws0xwAwgN5Kc61/KB30mQoNznjQVOjFfs7dKfw83HKUShj/RE+q
hG74eJDKGU6GXAltG4Skc9OqoGGfCFqMp2/2pKmDWZXVfFt/3FXtw6MHrRTSsmQR
Uu6NIdaK6V1WLeEy5lThMUpg/I4zj5cP7fGrQ7C5eqUy8yt8jGp4sPpxGri2C6ZG
gMK7rdPagyZIHeUhqjOnpJzYDPNxRr9fdLw2lB4LDQsHCMwIHNDVTAQXGuxRT5qL
oSrrfnw4fyi6rR0kVRI78XiH2dhbxUZnsdnmmrOZLinwgy6USnNa32EQ6wE/+hpW
CngNiA30DZratAbeQzaXtdJTYrQIMpk6+RXlsrPSQEvcWlFErB+RS4GPAbC2e/ag
j9b+j0bz+I2uv3838KH76d42v1/FVJY9/EDhZyhq3AiiquPL/fAHthvietPkV2QV
kkCa3u98IYEG++lHrFlE83iMouJx2c3/tGZtHuYKCN94VGYu5MJPu9cewpvJ1VuX
DW8u5DGWB0/WWxCA3PVtMH9OmgfIlmWaMD8q1Jooqtk/OFeINvTbjbTDpvqewQDl
V5+evbjUi6/g9S1QQuFzjyetX00rprSe+F8UOTOf3JUTLq0TW9uMzvLAWjDhG4cA
lO/8/QZaxk7HjN42HE4D1LUXLPR94C+aYal+vbD9qpeGt8QQxVZ7Wu4C8Vc1J6zW
/hw4+r/wRDcYI+z26lz0iCjTYwgx3cgPVPoQIglvJBJUeoUnYrYa+MZUnxahAyYk
0q8C+lkw25HGPaeDwnqGRdo6UvS4pEI+7kMfAMrVzL6rlTCGDa6qkNgJX9nNnh23
JQQv+D77AJ803TXMQgbWADO2t9CMqEGED1zZsMqLv15zF9Wy4MH7VtJYk+CIw7MO
bA6uk0lYzWQN6Esaa6nKmnkoHLwrwQe+R9LRmZ+N4madezw+21CNYIpfACowYAgE
ffWnsucEMJLoeeczlDWpAmoH8/Qt0XcSjywdYKwlv3MDxNo99Fy1vIxj+BcFEAXp
MlxPIlHgGZuQT9Z27wUBxl64NkHKZ0lqMspBmVYl167Wxgn03PFnKrdgEkthEJ5/
E3jbRQypGHrqedt1wrDelH+cGxppCj1nxEr7Xj9S2lie5pTERwScyf9J2d/bo4jB
HvFho5y9pgOOUV2QThx12UZcmNQxjAn961l1EOPLY9e5ksywyNuu8pWSbLhGO1jI
/xVPxt9yGYFNjpN1I90pISCCdqBkLJig2LRtuZv1mB9gpn+5fxkTGJgZs48m3gI/
umyWd2IKWIBL0YfGMXvAdWsrRdYeSt9SjeMjTIsyKPefpqt0ofbbmr42V7qSrOYg
Ep8oaBgsajSHzMz/kh3FOehlckH3t1B8Vi3eaCM5sHqbdZKzbs0ktxpWseOVmdcm
cBHFGDH2lpK7tqu/RRp+51wfhc994lqemdDU0vLw6q2iuVvip9jC6S0AC7031jOE
XNrkhqE4ktcs4pbbuFJJY5AHDNmFHXVtOfh7uZwiG7XKOL8vGVCTd4a7R69Uhwpz
l8cszb9GKkrsi45sEnVM34N/HbJdtq+KstApDkKuJLbnzlbOo752TP4qx5kBF0tE
iutLCxOMnHJtF5b6HNn18FzI6k+O+OVAAXLk8H90KRbHP6Pvxt1wZ1KJbo/A4lzN
rBT21jX1Ecr2sa1yK9hFu1Zu9+L5nC9TeDfWgkcSPGt2nDQqcg8lQDLos5g18T7c
ObxwEkV8f5tHXNIzqkxjFBNknJ/RpTL9jzg9iMZKkvHNxpDv9g/lden8KJdcAtwQ
g/elApRnswyjFwgcxQNWPmQetiYsOAp43UB8ly4HpmvZO8b7EKKnOujazQhrrWk+
DKC3+S7HKAU9eBo8KJYHWqdoJoiPU0iC4+TSAzq7Y407oesoKuVvJ51lc/X49sPe
3on+KdVfrVhOFOjmRsjs5XNudSJ2H56EpYeAX580819v7icNDpoUsAnYQYl3a96g
Q2ZAI0OSbtQLtppC74GjivVKJ1nxFgrayqDU0vtoCReNcsjFoYv6WcRWLgsyhCHM
GSl9F7ziWSkSyLN3uhjj2QfVaoy/LXG9ePcwIdSlxMB1sPqEwXaGcbMA8NEY9O3O
n5Y6WcCeuIVovKbGQE35/kmWq08g7F5YAxQdL4WbEY1zip5+LyUMSl1zu0/DhrPt
cfKMRcByv8lIf87gqJC5xeKL2YeOkU4sILnkrh2OWLmf2iwMnMOLcRTyDGK4dx83
/xgLbD3fQP4Nrfqh2D/Zm6coiuwi3UOeSVD7VD1yZEv3F0UKI25zIKNVk9o2Emjo
pWopkavC0HM9Ea8ONMaWiC62m3Papf/GyoP3+kDtdrnrXE1Mzwu4XaIvQx7MrtE5
+0YB669MonhWAyBtAePEA/IjPk5h9uDtmDNeDBzcRGHl3zB9PmjbcJ3hwqL0p87c
ojx/BV15HCUYss8yh4uvPUfulovVKuhfW3ebmdpDzhGoooGbZq4+aQBlB+cXRGbL
oB3z710MAnEJyge/BZE5r6s2g+homym5j5FtRCDg2cd9ficFyadE1P4UK5b0f1yc
7cQLYW2qxlaP/xDs0Hf9ZsfPwlgnHNgxQRUUdZWbv/1KqqS/DPu98X9xvSsQqfsC
HhGiQ79eF0haxqf+KjL3pkOPEUliSZpKi5NTP4Xg/viK4AauHaWFOUX6eLifVPt5
y7QyxK5EzRB1zx3SWivOQ6eVfwabjCAFScLOYufCctUErST7171BVU2dGcL73x0w
WKb31b6ImD3bWgx+6HZtCo8Lyn/4g+4W7f99icIt6JUadVGhekhhm5/PLMpmr0Hw
C8ThRpCO8RPq2PNcMYTce8FikIUCoRV2on7RE/cv4EdSqurfAjvkk7nysvFJtroL
YKcuY4IlvFygr2Xji3cbIQnSWAWJDT+I92/PLKSxehB1SbXNE1+xfq0xfdHjma1+
h1bjhDRyTdYe2e8u3u2UNId6kacnk/CXpeF4aYUQ6tfuvuMhk/tFO8+s3zBN4vAx
vSbCJSRCI34mh6AKiJbtWuTOa0mqWrcWUDir5cnYyRr61591ReX0zXe6TApswoms
+xQSbj1YKm1z1ZDg4c6/Eh8mf/jAkHp72NkvHOOuSdP5SwSFlBOxu1DGV1zbq6kV
4/6kY6D/hI8x8zOjQ+dT+0jj59+3RtzuuEhiNFbOzukq9WJnLh2q6WQyA7b0DF2E
ikR7eaYGur7hBp4ca2vYcIiJAzf5B3W7piObzZdTxoODfJFaE/pu2aQ2vD+u3b/t
BCZepLzNEG9M2JMtMEGLQvlDO6XscCf+c1OMQ7UYJKOQjIBerLgj5tkSSRK1cs2D
Zm77+SiMdF5zfTj2ykB5grdujz2nB+xYdyyqNa7OQSWo1BoWkaRjcSZhB15qrIIu
N2VQs5/JKFtH6+tp7Jm7eNQpSpDelteyY/9YkqC62kpln9akEpcewTB8nkMkBt1r
f/FyU4WRcR1N9nZD+FAjp0mR0h2cajZWEW8xSm6byxgtzRIO0Ix6z7nWfW2j1Puq
mYqxMr+kbRBbizUHv6ZrjjkNRD/VODQQCa96K70CeaTRZMau0M/VdvrDuiViA8ty
DZo7TGxEB3Mvl3QHGqyhAKWm/x2sYLPObH+QLukjWeHwDe6WRxOqVLCLS7TeKHlL
Vr9SHdfmin2FYRSpd15e0MSyLbboy1q9eeEUNtWR4lOpz4nRV8BV+wBqyP2FnpEM
UsWC5xiY/0LbRLDyH20O0ddJqjDUehj/Qvz82jX/75ljoP39tlpqoiIG+7FAvZ7Z
I/rivzBF2RK8+wseGUzt95rajDZe2COOKtl9Q/qtW+rkX5Fq6QrUwMnzwyeYRCwk
S5z0AxjVo3mBET+UIJ3qvrpEUR4HUE87LN8/AxCui0YKQgbedymRR8UrYiv0ujAA
t/OEj/aiUn5uCXN4IQ8o/PzhAfbMfizfU49VhaViLWZgfeQabeuXmiwK97cLh+4R
ntG7JIWdawf9+E24WFzvKXl188wxjD3yQeE19QBIlPu5vanHO55tNcMZ5CsNB+Ax
wunsnfuI/sA14LGYTfTm++k4REl4NoKbfaoWJnEs/WJ0PIygpdiEI50wDyjLacnr
OHtIGtdd5VxDx4pupXC4VrXqrdFpJzvc0V04JH1XAoJ1uMQ/DsVxeOO7w1NYFlL3
XZQzCvBL7zwuCmZ+H/rnx3a+izjSvfAcQfN55tjRu/yt/0TS/5bJpvuhVb9I949B
Q4xd+Ci5PelgVkTmiJLzDoq/b5wd1e1iVj19o0+6wEQ9/6lpckprK905eDWtt+Fb
PoBPJNC1FV9ani5sPIsKlVRbBo5uZBEscUa0zxO+KGxvYi708p8McLnVKx8wNbUi
iaCsSOi3MfE/HaOAMuiCpuELQJohCf9+c6XwOdaOlVkl5NBip3j4gOKsuAwrp8xY
8hPSa7gLN16Om8WN/rUG+1JimVcCy32ZnYXckZHw+9KiqIxcAZa38dzFaoTM28Wi
Jj8/ycmMhr1nQC+Ixvw4MGf08Aj3fKQZ82uJvkXlMwsOEfmlzWDkYNimva0rBXZ+
xN2Mh/s5Km3z9Nt2yftpHn+Pc7XitlTRezr2NDxNySXzC2/tzfatLDvfOO/JRV7y
7dvFZwudyqSEktzIKdziaZIDlh8lT2MtQLbsEgRP4jPCdPb2X96ncApUtlF7oaLB
thhDNmQobkhqhWAhAUpM6J5QhpULMkjH9OX/6SRRTRO3mrijZAOUzTU1dwM6A1ER
CzobjThdp6ZxohwtE9CCPUcws+TTeew9i9o/BMVx7TljuKn661PbdVKo0jWqeFrw
Yp0rdcg0o9TFwRbMGeQKeDOvS7iA/SiZ22omggGiHj1pGlVuuk9eVZE9Revd+Zv+
Dg5sf/w8Tdop0JNwDez4xDs7jKiEJBsxcSlbhDMa0MJiLOz2QiZF/TEetcDjNccG
pJm98rNGrR6izmKMW976OlArdfQSu7ZU/HNy0qRhmjkfwsLUNmCjBtf9F258O5Zm
TUCWzqa/LRn+fg5Owol6c+5fFcOVVYrJ8ZC/7luqYCO/d2F6ssW3clLsuGemV9Pj
noFR221C8mEC2xBeol0Jl9bH2vmydl71m+eWLQ+JijWlKic9ClqmLJTLMJ7pfVEw
nDHIVm8veTx2MqDFvr0fLiV+7/H1tAIdnU6A+Bn9nzD0jkq3VyFGXmBb501rKbqi
vNRPv5BrWxwxSDg7R63Jb1GfXkf9UqhiyE6KxBRFuzNMMLkhj9BjaSje4zs4MXZf
1dqQwwziUKuUOJ+areTF0ISPYHgKYWeHW0g/Rpgz3B7qi8q43EPsrq2Q41zEeBih
aCU7oUdImON5oQV2nc3qXCxfB1So+v2GTzN/t/hm37MlI9Nekywf71Y6HxCZIBL8
AdnwwL6Y70RiUMgAMz2zMWWN2IudFHg0w7zUhng70JDWz2udujorxd0s6QSk+u90
x5Dvd3wtgGmBBX5SXO8BpT2tudX8Q2W1cc1UIHernVDmfhEzvEA7GYXhhOsVM4ZH
tfQ9gin+wJxqc0VDCg/i2SU/38nwSbNSsuk6ohAbQeo6eXqT52J1JkGDDhDPFbh3
WygXHVQ04V8KMZslqR+M75usbhi4Zu3pV7l7Qe/yjnLNH0pvWaA46iUVzpREvOyY
HiFDeD+bTREuZRTKszN0MSRvcE2FOhWxhNIX4ZdZqe0ZZZy1KsI+7Trf6Irh19BF
lrWF1KnvPLfYVw4Y+rmyajdzh5BDPI+vnp3dRQY+I+a0vd3J7skwiH0zCwQ9AxJw
9+6a879OF2pjqYi9fLmYrI3HNUDaEqmnG4FPjgVoYykuo7LnsDj2BrRl+2s8pxtj
V877F47uBKOYUWyZ3vlz+8A9rM1tU1EQp9BvoJGNyYV0+AvjQAQbXkZgIneiCUMO
H8Roe3qsH1mR1AqRtWYQbNjz27FJ6upx4I0kVmCwY8O/LB7mmf4ilAVKXegEdgAV
8Muo3UPWrKRs5El11u2+ac2X+BSjMD/diPAe6X0eMG79xMp6idZxbUhpDoNqUTig
Ywj9ZnzocC7s4t8B8TzFT3ik6tSi/K22F9AsRZmiCE44GeCTiWa44ToXX+OaOrq2
q80GyQ7Fia26DE2HTlaHwMSuaNagYjWh9U0pX9Jsa6BvNcp6WC6oMMM0yvhQeLrb
x24jsYqL1BOKG9Ben4vjN5Gmv/nECfcih8JD2QGV17EuE/0EnJjXeaTdBDC1nFyl
RgaVC8M/wYnk3qtCkp20So7qXE1iGM6P0mjmgypm2GdXzMbgGGbl/rztmAauv+M8
bDw512SJ+uYSKI3J7d0NBKVdvcVvM2pEe3xdSlHBSJ1l6s7SQE4PBDU5zOqPTxie
MXDCKkGUt+cF2rwh3URV+njup7Akz9rSvpkUSVJVghoYTA+iaisdqo41aHJPnc49
WxV5OMgpmmu1bz9jkJeoVaZuFGZtZY+OYGG1DY1iZUe3cErUABb8VZkc+3YMyslv
dpxwMMuqr3A/+muaWVNpMuk34p7WN0l+7dP+2NSRCdBPHg2pVIcZJi3+Uih5SBnK
lAN39k6IKlukgW8rWF9EGksCR/8AzeYNV7o/Ak4ZOdw7Nz7uqnWQ0jAkE6rjRM0w
CYUtkxWCiLIIx1riW8rbyNfuB7S8yIqZxXzUTd2l68snKOl3bdw+aNLp2WW19sEN
R2wFD6vLRpJl9rqDwrS2K6W4+LLGLyDjp3d11yHCmhw4EGTFmbMJf9jAKLk+S2Qa
CHThGjhFeq2pkJkG3V5HIcRY9aUrri4qrWvn4RbbzSeCb/uU6AWxOHq4lyTrsrj0
Pn1jWf0USj/eKMB/c2rF1Ncyys3wEThmEHXgG/h17ZOqPNsRchdiBC4e6BYZTw3k
RQrPsIPeMhjknBCZeXDYAZItiQyN7gVAmWmkO/H9rmhKJeWq5iPhhJOLvtfxXDAm
i3MpUZI0gPzjn3vdVunSiKhKlL6QdR5vP+jmX0Y01KGvLGYJNLAIE2FGvukiEikw
0uptZEEeWLR1VNzxJWGrtuEHgnjCqbKWXWQ+M65CYifIlNwk1K7tt0KlDPha7Fy7
XW1hLbI2DUo28UEtIeMn34UV4UeH2l5f3WkaK90ivw2JbmzAMwdeCPz/WZrr+feM
35g4GgbWvIomzSXbSjG7ujCbjJJketvgo2AZcYpM7XvnNSrJS2U9j1JT21PXwjBI
IeuenyNcXTTCHcbbSgu/gaNQPM8OaUrhXtu1NqPLjNNbXacxKv9JNuAJJXvLvGHr
K3ZlCkSF889XwMiuR6m4OSnvi2Mw3DgDwSYaxNM9L2ajMT1ME1D65Izri96lkFrX
Un9+6wUqGlZeADudEow4kKUVZWnhW4PdPjeDYhUAOFcfk0ncdr9f63tlXmxSEdk1
hGUNFUWUSCjwBkbhmaqKuFh1BmA45xFB10EZM20WA8UGqfFoOf1+AFAf4uWkfOtx
Xj4NvH5MiNc0YZ05fFW3LOAvHbV3zOuSr1t1DjGeuNQdu1w9C1QP2e6EtaYFQ9y5
KJ/uozyYZbLxT+gfoxWJp2B2OtbudmmzQzi6VoVeK1Zak6cC1icP6f/qJH39EWWz
rxWQztymcSpCeUc6zBHGF7QEhswERmL5EYWNjYb9ba2mUhvF+4ehhAWlYHJdE52w
kaRaMlRPgbA7q9QqueKGN45D/IBTYhTu71Mojn9HwGaHYVT1UacPMrek0YnutsAI
4HrOEF4tnIzCqhTFYp5EW5ViKGosb/vYUi23ZJv1LxIWd6Pu9Bdcop73XMZVhQq0
unlJgsWWMlzTBc98O8/MhzKapefCIZPDgkWkuniID/qnAZ8pslIWz6YDvP919Lsp
5gP8dO/lqBaCitVHJM7M+n+O4CMzT/mTiFgN8XbVtGPxNxvlxOAb5c8MtOLa1tg+
NMGdtY25x19xMMiF6oOVNio91WQdGlJmY9jVpiqOzQQIzBumwji1qyfGZwczjOZr
wtH77YJDE8DrNp/dJMuiSgt2jq1lbA8oRD6GL3Yh5RdN82PLlMcMWlAb88vJD71W
ZRoz03OkZa1Ajc7F6UkYbNYjx58aNlMvCFH/wC9DKLVQFVYdpfTJpukDjnEmUzxk
qtyhhIMtDOfeSYcefaV/4zaj/bpIHhC9MMg4OibI4LTwWdoYHEMMGrp9H+R77wLA
IwckWzRO1LtzAYv6z8HBLr2s5WBYM05+zRHxRfeNBvivibG2YZSnFGjYPGkwQFMb
qaXlbnTYanaLfcaVauFgPhk/hv91P0EqXwmmzj3p19T82sWHOaY2rdTjmZU6NEAm
uLa8ma3J2tFc9ERVlazta0XpnWd1tH75V6uEguq77Mkmbq6b8P3tYUPe4OJ78MOi
1bkrZQ/YrtfcRS3gyUtCW2qMNt+dXfdZArHY46+ycqzBj3UeM4LFuxrrD9tHU3L/
cvkCAB/mar9txSR0cj5NSODIAXrYD30MiQ7WSMzxO7gSqTTa+FiDBEouYcOgJ+0+
IrQx63ibfBImD/HyiKdr+iERGi7FiQia6v9t3ivMqE9YzUJ5QpBU+exvbDjTFOti
3kexHVVOLDSMN7XRy7AH1lMa1ExBfQ17t6E1Of5ek0GoD1Ebgg9LotxGooLCfSyr
ygwdKJrG6Nlh8gX32qYegjz0kMz496FFh+ZzbgpWKGc0ZoVXlYsHstQJG5uUgkBe
AOvK+ZuFSqLmxPViS2fAqg7+I7xGFA/jLCkZIo7re/tU6oEAfsGKAVMdrMtCRYDO
0GEaTrqPkUA9a787d0V7bz3i8n9YWTm8sACXKTH2OMQFVq/HzNCZKIIFt3ObAzNN
OVfpKsUhB6dJyDdM112YoD9k4dMuO55FIgBrSJxTfjRHzyFIgOlKMQl6tc2+ExyE
TGTm+Egnk3IBKg74n4vGC+7fKFri2ugh3ZRL8Blz/seCmR6Eip9kitGCz3099epd
SSZghZaqS1i/hKXSz+e4PDmmcNwBY4fn3dhKRJtY8Ctrk0mQGWUTr3X9qraHAtbc
LvlKyqZIoq2Kd5fWM0wTgy3t2FLbvnDTCDk0FvKeww7aT+XK+jeBPjpPynQe5OhG
tfU2BzJSwretPncYCr+zOZbzOEOTIVozYNqrVomgBduh5n07e0fiG8qzArXSGIxU
Ac7Pa3Uce2tRBLW78/AaW0ElZbZiwVnDbBVEMmEP0fnTh+Mbfye1Gm2qnAhA3j8l
vz6HjWZ6yMEAbVB7Yz00R4IOt5BrbroxqeURuhTdo0uBTBV/AbGw2gITYYtRs6BU
ByDKHg1xVFYy3euv+Zx3U5bywz954UNMa34wSy5fl4BbEgUjhoGSB++0CXlPDo96
+4vpEM6vUKfUeC9/mtuMtxY3W1JGOP9rLTw7YnTmNPWNLJB8GH++bcVv+Oa8p8+9
9ssEbw0Mnxc0OtLLieXMcyRUYmksddoqFjGlnKvepFwLzqDGAzpnY8GUazUY2k9v
gpgHk+ThpOe119g9Y5QslczVKK5q27fvYQT9yAxN5afsL4zlZiJA+Ul7ZkwcpbxB
GB6nFCdj4x6v4EXTC/oYZ1lmQrHYVCIu3QgLEtZmIflZju2RKhY0GD0SUiXJY9ik
2QNUzpPIvdI4rFccaHGnLRZChu4mACIrbxmrQljGt2ij3tnjf8xQGd23D1ojiuWo
GKqF9VzxahJmw419gSqEG7R0BYtcHx76W7lMnLd46yifeqsxUTAYQKr9ngivu3yf
1BYyM/dYnz1swD8n+wxNCC56P5xR90KKDgc7XKWGkk5G9vNw4EEhnflQzzgrOuXA
DAmJQeFD3j2jHBUWG++Nxb6VRBBip/xA3FTClrPzBt708E2QC/7VSBS9FxrFSEIl
tvQIq8fGBOAibRlsUkVNOBlOhHFwNkKuLyriB8PVRWYOWqeB+aBoYZwwZ9yvIdpf
KYfsf8HjJgrXeVuMMiQo3zf8cDew7PKubWVUZETkAK2vgR6zGYNG8S+Acmixd2uX
JYMrUwKsyC3WiNgvNkYNLIG7bBF86scgh5PHxRg/NSnk/lkRMG5Mouc8Gwb5Oh3A
s1ZLNljB/uEehZlqNWmPDxUIaFaYKF1YeoeQbv2tGzGYipEcEPlm3ty+0dJB7Ttb
EeLtZucDUKANh8mrhqXbeYIBUhxOal5RVSTDhTUwqtUH0Zraq7gsCNcKh2GX8mgb
128kYcN0RuxTS+nquY5MVQJWk0RgRZ/0V8D6soXbursMR2vDFyR1stQqCWf01lrl
YooYdtE436uDGywOS9mvza37+WapLHTYMztmBsk03odScC8oOJrl3/pkj47BHgh/
D1lkmX/zkhjLGOLreBUkh+n1TC3RIPaUV6Kkw1bAGjpeoYeDBAMn/V9m/JcviGL1
/nbxG9QXRPA3d/9R3BTb0eq3uy8CwpxQX44gEmhAEe3QZr0x7bbtsuvQzUn8eLY/
Mee6gjXw35R1E+qm/f9YHFpckPN6mnm5WXUpdJF+4bacsHctbVYanlzhJWOlCGnE
t1TjesT8V7yUVnhFAGt5qKh3w4Y/PfvFFW7umWiUUCTe1lKVZnTs/OCnFj0nKVTU
3TlOrVucWJnRbdOrSu8eTRRokmAEpU7kZaxP6/0aJRWuGmxuQAhMyWTEoSt7BEXn
N/APcJWXMFsaJvnuR9ZOsiE0g1gT0yqR2q2oUNBGne3y7lZCQn3LmEdlDvktL1KO
+DAW/UKnZp3wJAtVYEPXs7T2iIfG/Gs4gYnFJo34pHJk5XKLqbZ6K7/jT6jUZXxn
5cDfKlZ33vYyenyNm0BbnbbERIe14v6N1YaFiKLtrqsa5wwUmXJn5aMu/3JwCzo6
Zm1Fft0ROVUNxZqXbi1z2ZLXQBYbnZp8cTf13RZVJeDqZlqmSpPf9njeFl4gBJKd
ZVFrqJPkq7eA3Rg22oMgTgf/bYsbol0GdEooolp4efqq8cTe/LrKd64Lic2YAsS2
l7Sd20V1VhGoyG2EUt4qahEjYzk1y7xoiprrii0V4N4jwXqqntl+s/8gXuM+HMWp
IXgzn52POjYxB7c/B9ezwF9s5voEQzHAcYpfZjs8GVAa+VCkt2F9Q6Pe8LF2sNWo
nTnkfgOKYHWsB+Ax5jdPCh/pG79beK+vuFw/7z6Co3RX/o+jGhM8U/uMljMMcpv1
DNiVhVtxV7lSbdoeWF8UBDAtfYvgNQL980qL4CqAnEYAW7IrPDC9CpWpGfl+CEgV
DnntXKgyInCFGDvg1zSnq6TxgaeMMLZdFLaS2J/w7uq76DoQmQHFuoTBi4qq7cm7
t4cNkpxwJeXbj1lctD/IpXnHy9/F/hDdhRyrW0HGC3Xvr1uowI6yaDCOEgJmy5FN
9Qp5yUZR7EXCJvuvSDuhB3TfeoGGq+WSgAHcPq+UEaDbSjvwLc2bmEsjnu6ByXjt
w1uOuRAYEKJZVisg7DkM/WAptZ1XoYArpvEDoq0ooQCPr9DSXH/uVZgEfNNeNKqD
pzLIPWuF9R8Myjsr7HtzF/YguBTo92M/nWtoJWVe7KAqBf4nJJ+KuHdj/RJCePAF
TvtJV7t4wzEm6MPZhNwAa5f/E6j3Ga0iD5ku1XuYSlBKLZtfry0hA9EsVJwpU7sl
ZdmYVQz7nh5Cs60BuYDnW5qFzy0TEq/wvqZzevOQ/+faf5cHetP/hzdfaz8SKUG1
JMMELCs1YEnfJ9ua6NjBUclzUxAt1TS9os4Mr6u7kcGFaOZYUGzpmROLqIosUKzw
C8eNSf31q4pmgrINEoGRD++3pzOAUgsWuWFTSeneaYx+m3AhqFSJ8EoPYfZJLGs3
xwjGTenxju6UgDMYJWUGODXn/AXiu3AP3c1z4ZrvF2MwVoguOM3+uMDv6jXK6k0y
opXM2Ulx4nM6rYCLXvRqgnYszr9bKIdGc9WEdKo0p44oYKp5mF4PB7wgS50gKs/G
FBGxIILSrAPM1vPTaBlMt5Pe8QZFZiOuNU3veOLNjdUp+Ebl0l8HYqaeuo/ad1Qv
iUf57g1bYb3dfF4x1a40lFw7xieYm/ku2w4Agjfjf7i3QR0xbe+YQPqz3xYAGln2
q6L5otzBgaswBs50giMYd7x6pOehMJnAVUQfi1FXRC3H+6KAokifbtFmRJDYtt0A
6OMD8cfuAAOsbI+Kfo2gQRSKhohtr8HOBtdIRON0CL7ZFWnvx1lgO/bkUzaBPOe3
kqvCe8RrrxgQSo9ITjrhoXf0CYKg+VrvX6NsMJVgOPFxgBZQqROD+fjoq/i2AsQI
c5rbRwLtf5iNc5m++Jie38mhooYsKyaXCnHCpJYnzQgjYNXijE2d29QO+dz9OoZh
cmxOl6AidxoY/2H6ns4bJFxXPvZ5G27cM+c0uiT8jMT4wuJU9mMPeiCCzYMlvz8C
G7RugNcsC0Y5kkG5WGo9EloXmIqXOAmLkvC8dtT8vqk5lyUhZjiYtQbN3Tw9LJa5
pbkKW7TZZK08pWBNUS7f0dJvJbQyZ4ips4OJPa+PnGj3Vj6Xz2CE+tH3lzPkwzoE
ZRLp8y+zNfWT4mAaLFaxu1WcH+mjQD78sa7dpNbaXHpgEQutR650e8Pu7N1rB84M
gLHOrdXZRa66od0EtgIvxuFVpoJsutjUZew6HrymXzGW6lM81vCBGXYIy+WbvYeT
Hb/Di6BHvUAFV2nbqumXmFO3Rt9T36yaPKG2pjq6Qh14FLQOT8mcGdabGOsI/yu9
Mlk2zPgqeQAmNMcl3zgwjA7Op9KrASsmRiG5dGQPBRG0LLwdFWwL7St9/PHA5mu+
t0n2+QbPbHvwlrTaWGU+BSCUNNA+8nvipp6kb46/KvYwFLeUcaQK6pZEkx0BXl1x
5xVrWtWvSNPW0uyt1PL14JF+IroXrR7EG49OfRmEckIG6BbixGhQn00HbKua5hYI
X63qL8UK8dOZ9W7N4bkaVkCtprukJJRZH1Y8StWNd6bisUuL57xcsTyMHNHgX5c3
YdcATq0gwDSz0qG2a5M2znx0PcAU1W0V5pVSjcQcY+fga+ruuuRDEhgt61wjVTbw
+hEDLl17g8EhAEEKALe2KAvlCBT+4Q58150OW0xF0wFdP1dW4+rbDbq0cGlDCjFx
JbT3RD6su6Ztzf8LufOyUhcsi48mNQL0zdbVdkHtmkRjyr0mKItY/paf4pou1CMO
xPIutHFigjV4K4OXlWhLZBh1Bj1CyObUBYoosGoDhnu4KB3V6vyH88Y+5HLhn3ZZ
iCXsFflXwkmNm6WHyVKux1qHTv26BPz/SJDezN/W5GTvl+r6AK/9Z36FDlMa/xJB
TXxUTCpMSd+QQyD3S8xkEexDyA4RPLye2u/E5HAlZ5eM264r1/BC9JMjnaiF1EYd
dfQ75zizprzQgyZBkKCTI3/dJ2INhUstLnOG/+M6uuGnohK7sY1ZalgWrzMqb6Xk
aHBj47hj5oIOtWGuyVds3g1rlpDidBMNd2HyeD6O+f6ell90il03y/8rgob+7oji
wf44ZK+Eu/Mw4VRtPnzTAyTRw3TeYYt99HKAy5/4QcyGrH3PXoo/41SdqcOXttIt
G61FDUE/FHOGThqx8UFw8akF8vxMaBMy4sDkU1js4lWYCfFFfj2LOwFF/UNYORYW
0z3oerpxJyT0s0uZWgEXSWH5P13U7Vk+ZRi300QPR4ysani/1ArWKvkJF0FX4YXa
l6KTywbb0i7IqFGozP+PWg6gNDztWpow80FHP5bBdfBXd688EOAu1DQDMC/VSrUA
l8XonYWMNTPxYwLhbIO5i8OVXuNnbXyBQ2s8ZsrXi8zuThUWsoYY+viwUy6YzsPg
fDj/Bj9kndB8Fcd8QsGOSbkc8FrGarakiIlaVI+pXWrlc95yVdRoB35xyba1AHTp
km3c+5+xQnLINGZr0PpVQE1H8Z6AbDbaqIm79XR6Urc7YJkS7BED9GOTusNY+SFw
E2XAFBwjeH9pudYbo6UoZ1X/DRwh+iNJode1Rf45vKARtbR+6PoSRurY7T0fYeOV
Mr1ajPZSNxm+OMFv2UNx+ntohN+lnX1Opm4PWKErXTIZQS2IOZODXV4jKTX103gL
v43OOtin8fWzszOTg7AoWPlPSYp59Rzs7CkpFtqX49TTgQ9xUYGimKbOHpaiUKbh
8oYNIEoobIWRtvH2ziY55Rw/g3mxFDbuZplfLhYzv9iB4qGQN5/BRmnRlAAa7y8K
2811IIMmzpvesqsE3twwZR8njOyO9/8vkeSQisDgs5h7j9oE7Z8Dr9YRQf574fmU
c3K5yxtqdY1C6KRR1eRvrzL0tFyQsJK0id25ZDG0826w8PpGWZx4Xqoq0fK1MX1B
Qo//Emnxjb5+reSmFhiC5KQZYXVp9a5mhvY+PzLQsxE5fMalkO5q2ahFXLIPyCER
2dQv6Hifqo2G5asECv4tED4WMStTPzz0WiaUfnFiFBlwXOJqilBPCgvUNFrc6hSy
wO9CgYCZS83HBvo+/WwmK7CcKPwwgVKGpCko/5JBVwamc3X8EK0LDdAmiRVIcFIQ
PWsWEPtgLrmLZK0inkgiFTkAFldUPfdJkwiS9MwXv/kfuNoJwQTlP6uy8Y6YLLcp
o2TYF/H3q+3W8iZmx3lfbN6qlR1Cq9ghhSDF1JJJICibSmn0w8HPitVcoZO7PdnW
qBHFVg9pZc+xKIS8LBJgAEQgwCZ6XVLoDX4u6WUOS97j9TaTjNDIIFLvdjRN++IQ
Ci7/0yWL7r2ATja+m1y/aPi0cd/ywRzFBiRG0W5RKrWmZGCdBXvTNt2MPfIwEad/
EvcrR5ZiAHgizUGS0wTHURHv2RjDhnNnltis0foY79cSY4dbx+xCNPppXSH2zRuJ
Wfp4pgyPs5+UerXAHAxFgMp6t6REIw/c1KH2zPiHzNkMzWCssnQoSzTA+NnXKIBx
4DWMaF0OxSFU/VFXb0GQo1AR2hhJt0rjkASl3xbJegph6aogxXV/ksnLu2Gimwua
znb1q6/m1Z0zMNBWkw9ap8phNkJSfj4yxHzRjoz5Mn/C/U8Z5cS0DSwOjmhptdJ+
MzLX+dcGDvEjzZUlb5z5BMbIPVlj52aSOdgNZxuFtuqhpRZLLCzqhdsgS9zs5rBC
sySomF76Qoco1D1tZ/UJ6J85WY3r1vbk3WfGV0gUmk3Ejb5DzUMPGUnpxvuiiQFE
5XrMwJXWQiQHFhx3zAHdyIDf0BMCXLIerjP6ElZd1GRlWLQE7TeuE3gD1nL6GD2J
paJH+zZkYAlyxq6FbxHaij38iwJwIGK8RTKOXeDL8fpyUfPJylEiCbs3X5QhzMFp
dz9t7IwvU3PPGhh5wp4XHjShwbuuQ7MnTYgX/zEA6gJyCY+kt5q3DOe9Dr6Kyyd9
OTU4TDxbXCKuvW3DyHUKV55gelpIp5lR/BrDzAlQ+YcC1c1r93i91/gAZ69Jygas
2+ZlKmnVQ0FOo6gnzMSikBQvCKhizcTCeuf9EuhA4kR48uezaM19ZfoZK99e5bgg
1rz28JuuDvV31OifvtLUtYgtHaZ1yX1kv4TH74pl2QaLZRvZV+6Ix0w6aRS7tQ29
LNAmkDMzzwWCWJP1ZSrHtGrBjVP24szX2rKqhOF1OvZ7AsUrtsm+FVYXiHtzDxGx
F1ghwIpRw2bJl8VLhsPdBkea+YqFWVUfbOe3dAuq7DrisMtTpUhxqI79sSFIdryI
DzdOKEzMTf/L7J35gP8oN3TqBwofc0HCuwme2WwzTniOCWitwgWZm4dr2gQNi6of
bCOOFWfTpmz9njYYGKnjlr6hxkl4lcbT1CrAmXFqGZY2a0a2itWKYPTrSOsEKp52
fGhilPikXXlaNYAQc8OcV6gkKq0nn/iOP4jPgdjUi+lVD4RxcULg8ah3BK7lxMJ7
PI43tdr2T8+QLw6vKAg6a8+fKiHkGBcNgzJHARAYVEPmOMwv5CGrCpKVbUZ5bOIG
AenREm41d5sleetYT648hc67ESHZcrjMG3TrQbGZme/ARNqSQwgyhDsmpcc3ubgp
C7WPelNvdrYIKVgP6RaX8xr9n2+3k1HP3ko+BD2MX8pfYfXPQfI6UN/a+LIw13rD
FxfRdoWBq5k2FMvg9pqTzkdlU1BQOVQBmH1RIEF0ok30Rn0NOqZEDNK7l0HeUqKj
xHv2IYzwqkKKJEwYdfgedi7DiL3fNsq6Rjtq8oOPlF3p1/bExMQ2mUvwRL4lghR9
qrDovHLYpoCw62fZKNd4UwSLoPgAbltPAceyfjOP73fYKn4emAC5Mz/xIq3lMEUF
l5M1mz6LIET0J0RGJccAYJ3ZOUZnVVLhXTe4J/5a0veTGO2nKhZLdfpuKlxbUz6U
4BLGVpIVFp5viWjgibR0ATQuk7lzrmNj/RLSdQwG9DWtGMX+a8JXn4Xobe3+9WB8
UedyG9sADYR2cpg8cFm+tlHKqRtC0GQtKGMjRdP3ops2o5PA9ejlB3G6viiT8w3P
qb4ieBzwD4oyJh3AkKop5EBp4+s/z15JbZ/Fki2oBzpZJAuXZy3GqakF00+lRlwy
VtStTbbhVtyUUa1KPoaP5eh2IKLXToymErpv4VEMusFV52tb0dcZxF7PjczFIpoX
TCIoyFx2lqCvIzWDqtNMhhj+qaZgUOjPryGHFyz21/Pvuc1nwT/st4Fro8Nh2/Sl
D2I52pATPqVh4YWRzoSzaC//3whG05xdmNVwNENl42zIFyPpt181J0lmmRwLU3nA
Wz4miVYMoiwmV9ld+7CORTmTq9iWPG39OsrCj60BcplRQmpR/Ii5nEmtY28KzDcL
Lo7YiZRpAjSXfWKpVWr0/PuVXc/8oxgSHSZVJvT7V8WcQwGFPyM2M2xH8vlM3sj8
S63eqUBTzNdBGDmxUbqxRWdraAjPSuag3eMQbBZIQq4q8onJtWD16f5jtmSxgkN2
wtLtpj9b3Pu+vR5tgWUHKHGoKQaNFXw9Cwgts0lFdSz+XihkgmCpNeM5pdYSRcX0
pTGGr/cQQzfmH+8ZPtdVmlEmI3qmB25+b4m+GRMgULxcvJxv5XjGK435adPNYiBw
Fc1/YddkR2FypiRRoH3Ki751m0Tt+pQnbo9VlVLBpb2O/hHGT44JfFi1ZvOyeR+w
gk7Aq0Q5aZyCEx4V3h5foOYA75L5CqxVPCEFUtk+9pikrQhT/hMhFOy2MwfgaPE4
2ucz5N4j0DHOl/vFu38rm9WmcgRtFpVk5R4Iw0ieBzMlioCBxmRbisgEyUV+HKpr
3rAIEprUPcpV22uHHzlKQP/S7sim5pOrtCJ9q7YZRXUAJYJqzcaCGD6YFS+Yzdbg
XRvSFSieOjHczqagS1HwBA+o00EDx54CUGJTNV8vu01e02V7Pv+gJkBRGCuwibzD
sAbevrk+WEEJIvQQUyPZTDQ9rJvxwVy4aRRiElF/2CA36/H3jvQGw0/2N8UlGtPi
PF0TNgZZ/14d/2QC92b3squ9brC9V85nirDpymcQrxU9Cr8fx3Ee1TKjgRyybpZ1
jYVvkXE/URJtthcYUsvBlPvSGJw2iiKXiwqJfTXBmmUxevwOKfl3gnNpxwc5D3Mm
fOS3ohUfV95OhQf7quUq7mjSj4qOo6SDt+7laSn4Syn6H25q+K7LVRWtUVkKYxS4
2XbgoFJuwYBfmRR8PCstYdbOE3Tnlmx+ioSVjWqaFp6dEnmMKZRGtjWCbzGNOYdP
xGcz0NQU0I0U7s2Y86TYAv7KCVvEnf/OuhqaM+B+dFk7O7GUsgVvl5+z+jD1gA80
+YSR4dMOskfgt3gQlYY2HSIiGcK/T60MpFnXgk5nSRBhK9bvOSUf9/U1MzvqP4Br
LzdvT4aOmjJbuv89eJaO9+jKmZopJ48kY8dIwN+f61ZvRVzVQoR9VmYUOI+uc0sT
zcZ7NO9SOF5LRJ9Ej9w3pYZzpIZIQ3wCYThZNZYJtqDeGAG4APTCqcWWGXo9Ft9H
wUO9W471V+oenrPCkv7LHNd2vTRPYRlWo6KcMVoCUDxmI1WsMrdtP+Yke2hQiJXm
Sb6uAUbrYtP1hvVM2KbNLQOe3UQaFMk8i33vo6dAcnPBbT/QAld4nZ9rn+REzxas
fWGO/mg0MtnK3lTiGZm5fBzw9ubZrpHed3XwZq/kWDH+vTYVfVRYXgDGiF9bN3HD
S7asaz5W3SL215iC4R5TDmtVa3tcY43jpcVDvUlDvWh+T8S8lvw3druJuO6GRNpO
x3AdhRCKbtGlBuGuhb5PbAnGORmIVRtT/C9DB75/tk3Ybm4ox5nd0/nPxj5R3dPH
jN7OBZsWoifC7gsoYBdhEA5LuBGdi6hws6VN2/lqAmw1AOjBgzlScPxHR1H4Kh3V
EpZqScCTVWy7aGsCzs1S6+OXBzOg12reXZ+jiJcwnxopGewBtSBz4J9mfmv9DI2m
ChIc1Kvl/6zmVwdfkFxFInNqNzbNdgvAS2fYXyxr/cQxzTWXHC6/jbauNPO0sqnW
mfgWHdG3pVE//LIffaQG4akXjkL6Qmgh0JkgsdwaH228y6788YaEW/Ox5cmpN3w6
v4gGXxv1836GY3dVtecnZ7p20Nrgs7q9LCnbTSydOSdlU1XLlOU+tgtYm1IAaWKk
Kjyz7VxQimmLOzpYNhhnzONyPl+FqsQTtte3oNhj0p1kZWp3OgyXzo3w40dpboaY
kEVVhgzMW05g+6k+Zqw1mCYLOx61XpVQN1PmQHesgVlpxEK6OgWIXt38A7aOQ8x8
dgqQUMEV9NuKe+rVt2tkVsX43Saz2KGFqe6LgR/KbPCGhrcLP9D9YIU9jatWh7Lk
OJ045a46Marecr9l586dmCxpcSsBamvLT9/jbBmYIlLDJB0x9TFSzM3yQQvgS4A8
tqgoV3QokSdpcTGnwb4UAbtKRzKnB6C8XQ1VG8RZqhaJI6hqaSgmBLa4EqG64sjJ
VoJ4L6Cbw/6UEFyIi76bmrtbya9weoJ6PUyR3vGoQm9qRgxM1uRHc8IimOyRoo/S
TphqJsRylib4Hu4Er5PGURlMlEtlb4kiawoAAs6bBNrF5QGf3/3LKusrnWnvJmIp
aXgFIXVNUDSAOvCooCGpqfHkpzqwBHLKsndZ8dLGdK8zk7dNgel6RZ5TBLzdp63l
vkCbjf/In7lnt0uorC1vjTHCwH/CVLosuBVBmDeFQrEd2C832w36vgG+oVnYDPst
st62Gio4uhBqH9KdsFEwUhwmGdU9wgY9B7TIIDa0y6658DktJKDw7qIDfyM9iM2n
JeFbAAQteMbiyiARnsuIRTSGZSuMSEObYT4psN3BhEOW4rIybnuy5Zstc8nEgaqE
ys9eLIkDgJTWrGfP2iBa5B+supeCjcQu0lBfp4AthbcXpS8VJ0AUAlfJkyuuLs5Z
+9Oa6clvnSxleRLCXAh/ZOYnnA3W1ePFVakizaCzyjS2WJ9+HQcuS1FKoXhgM9nv
yE4VnNCEip/Abc8UlvZF4mLBsuXrGaau7wWfRC2l0qQipex4rJbfxYycMXhy6ZNl
rmBBPERqOllhFGNfgl1erivvHCNzi4EU0CZzJ8c1Luvj1Xh2V0xNSBGZRzIDYWY6
gWGLHw5DwLC9nF+NrOfUT15UqoWAxY8D+3Afo9kbK/c4JTidaJO4A2sIOiRdK3qB
ZTBGPRRUGo0I+1NnaGn7AozdqEiMF+FdZgAfkehohgxZgvhGsV0JQE2whLGDxsPq
sNvAEIPWaaPnKczpRejD3A6lTriODDi2Xgno2T7iLH3ocQrh4jUgfSxXfugUINQ4
ZEHiTG37SVBo17317fAUOWzirUuRIO2nKAvaHu+eX+TEQ4nJh973fPb8J+EmMSgA
+Ze4d+yhpEgW9QXlL7fKX1VtGe4eQ14PJnfgI4s/stW2fdRH6NcQLs8m32VL3TNu
U1wm0buDJJu57RuWIRaXaBdHQiNWvi+LCqnZ2XNe3xCQGEXUgkUBVNsZPNH8cVD5
OpIDcXn1ZdwfIp6oG5SCf82noQAhmhzdhPxvUgj5uhb5HmV4sdzNP3w2LUvS5sej
mQEHPsinaGfdyXewyRlnzILHqQ0fvccalQF1DJgwE0pX6YBDlxb+7qFkXvyVmjJf
kY7Duixz73Di12tkCG8sjLNlODrdLFow3WPx8lZg+vaIMnz9mFZa0rRn5C03EfeS
uFFIScCM/3ZC819DON1kPap5nxh0EnQl1Fe/idFkpQ1kmuK6Z8MpE8GZP9MPzowF
327cL6mZ1GXpVFusx2/cZKvibYLSJ3s2FLx/IrrU+peNRg5Z/LY62AuYduWubNYh
712PqoR2sac2HZwMbTu4Cr4d39vLrGL8ERcyKoQtQsrqAOp1fRk5bJ8cTbqP5qvp
WooESj9XHKwDwEpoOrfylz98XYtpbg7ZVQh2nJiA6QVrq2hltNkBZIVfSTEwU3bT
XLkkJ0bh0LYCFE40BQxMCmHwgi4bCuxDvsR8kn3ECcRfG5HtvWk2qH5EPYkWfROO
FIPirfm8ARiHebC6aKS32Bpmu4Ho6p5MgI/MD3Q4ykk2ZK/G2jwFFdM6sNNPEnLK
xgnWpkdQGueA4f+jBPEgpfM2Vnnprg9R+ko3ToDsJT8+Ns5ycbCuuTpaL0squM1M
LcPgNuCYM8r44YbnOA2o1YUu2QdGp75Bq0S9MdmncGRvQXkgWL/ZPsGo7zw9y2AG
aFPHbs1kbMfg00pIaks61/WHRlo18ygz2l44/MCFJM0fMOxymXa4NZOBiO9PRJ8F
xdlw91eo1Ov8ZQPgZC297MsV2UHHB+NpPXEzaQ6V2xIE8xyzApuQfptqnrqKgMfP
HP+/eDxAB2YKipsQUOaSp1QevB/kgTadz8s2ooMwjOU8YQvq7utJXzrhl35nQ5bF
DqZabMXM0SMQWEQKTBPPVkkg79AHaduwxkd0UCN4/hPMopossXBVmw31/bDPFDWt
ajAbTzyZz/nRnFUuJdsMVVYVeHVcVd62+1n7P9L8N9S5yR1lekeccITxBiowZTLT
loxCGUeQdOzpVuYYVMtdiudeVPTR1J5e7VFIHyx0AKwehe99Ei17r14kUkzVbrZE
s0W9Yv5Z967QBXHJiqjXP4Fa4s1rNzaiGyiRlZexw8ok7NIqv+h6oFF9ovqSpsK5
B7uIQ97syW6AC7mqX3pCh3nMAPN7iD2yRVNe60D2Mn4bgc8RtbhSrfLuDSJPzJuD
dialDTZIXV39vj/1vBNoiAXv/topFZlVr5ez8b3QbZXpbFORFMhfbRkdEvFTos3b
A+Aqfft0ODe4b9z8eaaF1pROx8ZSKFcMvZjQOt2cpcT2RMfjox2/gTg2MxpCNaFG
bJj6/j9MPKQLntf00UkkukZVcGqtu2xPZ1Ll7EJqQdP8gdYXe9mFe6Bdly521zq9
zZo6dBjPVdBEeXmGjp8oRbXm0lmHpfIUgyUmtN4QC6uMoMs0xQW6CAn8DVjPJ7NL
S3JlE1u6QozqP0DNs5LgZ1XDGEpa9YooB8VHsUSPsjArHMvivESFzjWegeI+p466
oyAudzrImjKIN+P53H7+TKR0EBJgCES05QjAwyygtzWnEiyPjsqt/5rPOHSQMl9H
rOK0CChCyKeWoQtEDCxsJheMhaXVQVOCCVTJtqLqvfvWxKIs4ZBRyTpqGFh37Zvp
hvgLKZntl+yCwLx2L+JVhgUqQnRYT9xh3FHw4bjTfVXo7HeeCS1EiEy9onOCHspA
T2tWf0E1sxhbuEzV86hvfU9IwnO14c03FZw8yrMH9Lzx2hKgAjiv4dn9YRDtYZ+M
BDongjiv5yBWeWFyht7qOD2xwIQ6ZKjv6JYv2kNCmyWlwBudvk3gWAVYyI2CgH/m
1fYXb9LTjzjkfX5hbzMyrUnoZM7luZB2YbUjQ+k+A6xkgYczouOvB86Go3DIEgvy
9Ihk8XWdXvb6v5wLMey54LlA6RTPjneqjRveY7wBhCbKPZe9H92uUgaGj4DMGMDo
jveFxDNKpoR9jmkvpLJzG4+t0NClc1lGDWwthnrpySKlxC+zGXE9UaoP5H0rrHMd
FMu9AO+F7dnkhO1ZYSAedfMxxGvRTpT5pnhHvqZHypvbraLz6/D2w3mtOR5DXAob
WnvU56zNg2pXcijLjDbQJa5iT++IGXA1AwM8lsw3+gO1QSi3e3xNpSbwFZVooq37
qlE9Lm8gtQ4pDqBjsLuvHJKCdUyeMW63f4yqHnByZ/HRaA0Fu2OdcEx02yYOu5X0
QQB2KuScd1sKFSJtWQwtpYshqh3dU4vG7Zz13J0Ex+WftRpud6KLW+8xmXj9WgBW
gh3UgUSE6rMKDKu3DoDUWkxtOdNTRwi21ufWnvLbOd+q7cZV2gw7c6gITAK8CZSD
ATBmr6kDc4dGg0TViApQvoDH3rzMGHDIoZgHUzxK5QZHMhDg2FC+9y3e5eoBualW
3sOqEZdlkyih/NPVl8xBMPuzG8KIqoSq4hzOabGa2W7RTY42It0wisRAdBMYBfCH
gnfztBSN1IYDu+atVQG+bJfCveLSJNn1/GZdBQ42LAZbok/mf0T8FzREbKB+q6Cg
TlUwq+KBFhwiwEHWfQSYDEvBL9IDAFzNhrLD4SnVD9wUFv4fegxF3/JiI1pHciE6
8A0C0FheyUa3MnORh3z9fujKL/07Zlj7Y5BfKhnZq//NFNnhAzvLib+WPax94WlV
F3i5wHebmc3XlyicgiB9ewvLfscTcO4UCYxO1SwIv06LQp0b+uuVxWZ8bfeKROGR
ljRJaFG+AbUNeEu/vr/Alqy0gy06MFcTpbR+8iGMwuruaWep5uJJackHDWdBH+nV
ANI8bnaeh02Sj9YPGQ61UYhNGq0NfmxAlH7U3bMN9+TQlj8QT3O/jeFLW25kNCNT
heh6OSAO+ge1jU6NDlYcz32/VCxiogrWjKcwuHwLHaFDIMRY04b9/2BNRGHR2CuH
I5SAyKO+08eFq+kk4BuTijC9MGr5zdVzi0QVslyqg46QJ9SZeikSDeFR7IWwcN/c
kHFlyKpDxLRluG1BIxi+xdZhaibMuSzFR97Ogd4Pw+4uxbqNv+PS56ifVS8nB+yT
1Apzlh5R0l7a1jRTitSpqqW1Dqho+SvTaNBf4l6yABhiRqKGcvCQXyPMzYSdaY75
RCDnvpD7P4/X2XNCjUC1peilrVmTYP/x5LYvCDmMVaRCrTkMPDeUyQ7eUPlyLhB8
CMLA0vv0xMUsKfedSjNfrkW81rQPFFRxz6Z7BI+F8KYqm6GhvryRipyo5d7fY++2
kNYMT8E1yNpbA8PwmmJTJXj6S9icQWSs3RkP0K/mwF16RnRkxBy25wpkbM1M4nXl
DXPNqB14zVI3cf3BhDP5JRZZ0KqqC3ECfiRRQVBdcJJwVMpiQTrXcom4sJgDk9pV
FrEYLB6i/mtpLmHT2CK+ttaV7gTOc7oA+Bed+Gs8yWpw/9df5dUQSS4T6s96Hc1l
uoYzrBkPQ+mVuGQt1n1h8jo1uasla+jreEueHMQfymTt+CJNCiG+bw8jAjOFSzg0
UbmfhbSDNIaJ2kUkAqUlawzUxmyvwXlM8pYaMXVc3mOxNgUdC8BQgKd70OECcr7y
fMfosOuJUPcZpgpC3zUc4UaEwu5+02uEfwLPMBrrWg1FcaIphjYU9ypgpYqwr3GB
9uKnMUphPFiRxUqm2LlRzPUOXyH4/rfjsPYLMPKWHHg+Z4taIsR3jVOnHrRvCEzm
SLN5lFDAHzL5IaI/+CWeIfPLGRaNzc2UBYnFv9iyeP+AJmw0+VHETPl3WDB71wga
GehAT+nFNI0Un9Kpxyw02MbqTfR9tsu/krFtluueZGNDZ6Rb2mEpoIzgvLEscVaT
OQikeB3RgTOQ1dNFV7Bx9qVJWCvHUeySV1KLexXp+Qj8YI4nnoFGph02PG7MqDWr
Z+KUwTX371Pn16qmf9a7PZwuE/xHmjHpO658iJyyNiQH5I46RW7yVBWKqOSFwkmA
Iybs12H3QB+hoOodb+mPRAGBvsqc8OnA/J6rk3CMeZmvsEbCGBeWs/DFZNTDI3pb
bGVesYYiCta7fxhmC7QYlfdD7GLZ6Q65m+kgt19jkPf4pkmvhOVVnT1jr8WMQcSp
ib4SDce7L+n2RFKK3/HSMWEu81GtoY6Lg6ft8h83tJArbzi3XHIyQWkajeusDyjP
FpJUdP9NuP/7H2A3kfsmUBNVi5RE9fvJTP7DrCkY4lbLIzCPplgdbs6zoGaLgNy4
7Gh5Y983Kem5fO038d2pnZ++qjPZLqpQxhOKyBYjZD0hGOXqLzcOTcKDTYILKjU1
aJxyjoBVaGDJQmx7wzCdFsJ3NMILLXlfkm0s/jVhrZ+GV2Sv6fNbsNrhJ+XBWD1n
pDTRf8+ehaW8Q3FYBerQFxUaEdW5i6jy5ZNVvJe3OR+jhVyNt9uSlSR5fgm8V36c
KY6Z03g78uS2j7ADUKUmrKjN3IMBISjg/at4fAvmuh0CJK00i3NHAKllknUaUDxK
luoSaiMbDi4/YsH2IHeTkTOPiyH435Kru0hxeIvWehzojRXMWgMgQvyov0+LQqK5
YHLYc5XsLGzZANPJwLB08dQyB4vBMTCc8XsJRvpmoiCVFyleG/VYIvIHyFGtCK0i
HWJEAgIR9YDqj45IjTY6FbJ4snll8fTsiy2i/dhUjFM8rB32n06BRl6hEfMgq7o3
DMHBhT8wAsWqzT7YnyXGmlCnrOpIuz3sNSZEahz/i2wO9NDhAPBr7h15bjz1Z7+3
GxRJKUscKNmsmaq+R1GRXlKxicEIIoeBRdafdr/vcgtMD3nqJRNGTeLOw59llpEk
Y0r8Ycv7xoMNXLaqeogW++IdhW1rNTKyZyMsHJKlZEg7EizJ6MExeXMomC7VGKp6
BbLNbm3WkAUkpY0k2HJ/ZeC29v809C7hqU4JXRTP2rXjObcnnezTFioEl5T6FSfp
/Qt6/OITC3UpwNbj/HruWxArNklV1AaK99q1Yh4r75sIcCRhNYu+XSm7BdWDhdEc
Uw2AKYlxnTxzc1rmMAbtA3T9/eTk9ULflsiWFjuFZtFmYagD8AbGgT+ZTW54LQ3e
5u0ZX0MjC1xWlvwxWZSl4yx+JGs7hE2e8BjqPYjiDpxSB9jUldD02EvcN0J3Q9Tg
C70ZTTsovt1oBc7kC7WH1Jv7rWFB7lalveD/PV+81IwwBXe9bj9kpg3QRIgaGzZL
6CyV3AXc3gs2qIFp31N1+5tpm6xIi/qFQHnulOns3Qmb1ZGb5XaO9nFsgK/83gg3
LSOESMkurdWlMYysYafMpgeNkGvjYBR+kRLHNO1dUmJcXDMerradvjf1ws2x701g
h2S0uen+YcOpKu5LfpoFffXqIRAqoI1VXXk0wocK5PuZC+kao7Y5eiv6do0n3KkF
rs/+opckYWNp3iouil97e6EYFsvwq3tq3OrDqMO+v6v4cSB4KTOj+97VEUTfmSlu
KMhJSHODHyiThTt4klVQusbnQ5nNMQZh351ItOegE7wdAlwupwoTQbNSTox5Vdck
9oXAeJTUrHCx1RVXOkR+Ps/eBC/k0kM+hg/FEaRmheEsrHSd5hqLTYj0WtOj3b//
FQySebLQLl8O8TauZZ30XJ8RGKZCEdC2+LF9f+XZbXoEFSCMZ30vCfJr++hKVxjl
xfM4PV5lIcCKe/3dssl3pkkiPjGo2l/Yh03C8HIoBbRi1pgXcjuuwWlnPkWyQXVt
kG7mE0LFWL6BbFw0Jk82uFajgVXbIqZkuWnQNnutm8eUoDLb5ZQvEsSEbFgUDMhB
94OtIdTx5mmc2JSVMJfLqeEt1ErecsL7yg85J++yyHD5xtak3J/p71u+OwVjci47
8dSKFZc7p5MfYCfpzdaHcWrRpVzNatkmPMwxDQWFyREY4MKpf8Z6UoqMRjjJkgTl
1vDOgKIuO33kUKPdhrsmE9/KNoSKdG+fw7SXj3c/9vSOKBV9tlV05LP703A8zILw
P6Cq9szJKLdOu4vLhEbJa/TC1FhkN1/2a8gOix6hYaWrvfmB651fAJEfYAGakx4n
ie4aZUE6mrDrAeyoe54RiOJ2pS+fxWbPrBneLmrnOJvLN9TVlqHoboiL5P8ivUkV
HOdGhSwUqITGimsZ6WIsfMK77afH96gUdqGXGNgsXQiknZaM3BQTHf+s5SniaDqW
bBuL7EA34QIRWbBvp1tMVj0RA4FzEZJCd62ObU6nEijLcCtfstpD8rxk4QiFpfYF
64k735HJj4ut8+vaxafvANkU1/zatf2rhzShuJxDplk92T9tY0y4Rj6pcJ0bR77x
Ntb/EAkXQdDTl96DmRZaD9Mmpq25UwcOLgMg+ms+imGgcirWTGbiiD7KKiBebogK
yhtMoHwMHExh/r28XjpIfItORgfgut9oUyAwcPYXyiyq4bvGy50pgzd37xEinFYQ
cK3aXGGit8hMJdIRKPrZcoN5o7vfhyjrGqhT5PZZ18zob2TmTO4UfM0hgVHjfYlc
A2mjHJil1s4A0g0IG870ioKQAcrJP7g+L4RRM1rI/fd9VxvTeOBUfl7tyCWCh/aa
VYRzBg3lVHWTQS9HQSWMhKM4raCyD/OPGbhuvnQO47mQbuzW5FFq3ICG63Oj8GS9
mkpQg4nDRq1mtVFr2+T39I4tOOF/n3CEbZc/27RpnpXQiUNoyQ2n7LOFT8hJJJ26
YaTca6qNgdCHT4GpbLWWkFpwOeVUFYxOjA6Gl5Vds0S+O24aUZb/bp5teHA+3/vy
OdDbww2LIBf2QgCPF1ygqdMfDpzk5SSucHTx1Gdueov+lRhlD/bFo21f4zsX1WHc
/OqWGwjRub9bFRUGEjwKWPXfZ8ItuEVkVIwVKivFqwStHeFkxKg/asuxxiCB67HE
TfJ0BF2/fj5LnqP73TxXL8scA/43ePwGYyophHP7jjHiFTp9iMxcG3/A5hrycGRP
HLG4jS7xBdYWRiAiuJBBITDtg2H5ITQk/wgP1OP9PC/ann6ivIXAEGdlXmrZhXA3
K/DDk0nQyoKq2OwB0RLRpBJfGtVNnUAzyA8Po01xsgAqc7GJlQZTWuCcb+t8KmP7
VdfHnPX4jmGXolw0O1Mt3DUVBr+4RGgbHpG6pRF4I7dClIBVM3Y2fOUPYjyp2fz6
eUpS0DQBNVnLBxbKjCLFNUOGfNQNWV5q3L497mORSf2+x75If9hHCXraCK2ugwLw
ZRiaNMxLDLW0sUMsLyJC7et5TsRfz3zqeNCVVhDLmgm1AjuynoQ6HlL3lfwbRjXo
jsYa0VUdJIRFNTQp3/Q0Hp7OLsl/CjGGBNcwD65cI47G7l1/rf8U6uM7vuruMB4Q
6gJm/jEaPmpgxo91D6USpb/+tuBtuMRuofFrMFfPT/3j31VBF+gkZtfy9n58frTA
yEUW4HpUdX0mC6dy2NHi0SyAtlVogWYpuuFhkVnTMU5LDBgG3i0ft3cZWP3RVyUG
eWg/xW0lRSGMsHW/sx5wNZGMeFIv1vnGkLtNExzWkFpVLDO13qWRt/lkDcR+ZcFd
GHedHdMICWKZxelF3P864DDiFCkE4dr0+aKJKxsWgkF8LP+PEbvAVHjS2N9zekfW
VlRzTj9tE+j+hZFmX5k3LILTpXWkNMkw0aVMU7nGBvqkhjOaJusGTb9LTe5t+W0q
c/km+wFmEXeYjHMyqkSL11Q0YOm8lQI1F06uoZmBNXbPTdxgtWcpa+j3RrT8OuFI
Ug7r6NvVBsjTei8DW+VudmDi2XcWj8cfxRUEDOqQz3UlvqU991tf2ZxTw/Th9wdq
C+SnfMOCIZqgSSRwBFX5R4Mvs7dDFdpwVggDQ1HejERadCyDxN3CATlnMJB8iqtd
RtAtky1PFF/lhoQvv6jsUz+nd0yxTAbTrwhOiQr6L8Fx4XHwvOd+0yPxr3ruiL33
gn+DeT3OVZ/35Mu65hLPwwWF2IU49ufG1lcgAxnCoZGdND4asZlmBvVu3qm9Kg+x
SXewOKZdNW0fLD0QRPduJ/fKJ/oE7x0SL3zKfOQtJ8Q6M1LVvYnH+oAAbIYNFgzL
CYKvAI/ZW2TinrtkkO2oZkyPxhP8NgYDfZeMFrCsIbwswpvat+VHjByMdZdcfBdy
HVnNiBYYYDd57kzBeRo43sBfbmh90GLDpnESrDOscehxROnu1GzE2MHKAs8jpK8E
fENoS1Mdh4OO6LaVq5uMgrQtZHdD45c2Ir5KfBFf8QxMQ6mR2ZOs1oPoe+AxI2yH
HKkYdkav756ZrpK1QJ3zf+FhZwROavZ8vHB2bCfcZUuM9x+ovu7uJ3WjbTcp+adx
1DmvFVr3MUsgfmewL9LYJQvgZPleB++bID1su9whsTHkySw06yUrMCcoor142hno
cN+xyozC8Mmpkl5WIfz2qYsOOjhmUrTX0OY10UXx14s2QGHCqGsVFIamqW4R9go3
nQ6dSiHV8PksL8BOvngaDd4IgRgvv+evtRKpdys3QUXFA2WOo1fT7lv8KbOfB1Q4
1SkI0jyRacqPSrqxWk4/xx1RAl7257UXdRtR2am6KJmL4y6LbxOdKMxLvsC0m9xw
/VWUs9Illqgha8BURR8wgvhaPNW3z5/S0TWxSunqN6Ap/CYm5LmXkfEY0BadYcCM
uKUNZvjuCZmY5svzcTfXBfmwrBbckp8M6ePV6E5euJoVci0q4xlU2BXk1Oh/xRrT
Qo8EpodPXctsnsM3kZ9/PG81fiZMG9pcYJJtPbzGcCw2g97BGZayyz9U98T+f/JY
MMI5pDEwAT1TWjoa7J9hpo+MtWsBFoEXXnf5d19C+sqRkIOdYVacTInfJDCVekqE
eHpbKDjcCUjZ9IyHpLD5b1oBVrRFPy7ozk5Nva27+sRiI9txEFBn9zHjBF2YqpJl
pAyBftLD1iU+N7J3kkgqlRzngIp90wQmCeTBRpMKDYwHRnKp+A7/cmrotTDU2T+0
KL7Zw0D+DB+Vf9th+MfhnVlziMreLMM3Crt3Iq5tGB2vDzr/H1YOw1er78Oiapa0
TB9sPK7ltbTVniPAXMNCxPEzGyQMGgIU8Jsnv+iuBle43+phJfz3jJoip/vQfk+f
vJ9JTJkfG93dohp4FmIrdVbdrJYZQAVc6nre6d3qlxXlXp8jTnxWX7QxoVZVPyAK
kiTN079DNViUeC4pYQmx7rRKrdIVqJgniiZwT4s867BHmKdw/Jw4n7e6ix3G8bSi
OUmV4PPDSFuSo+hYeQeXuwbwyVP2U+5SNajz4wNzh4BA+YoeDPNdYFA8RAHwV1QM
V1WvFx+cotEfUc1pH7mgLV4wfCpTaxvAYkPKFQjlYDbxEpV5r3sSDkMuKuCiKCGe
B+pYCfLhT5EkShPYQAPdpSPsJaQId09MqUTzDCrJ8Z4PLuh8hnmd6KmGYdH7PyBe
HyoIjgItWGE+yQ9o82pp+sfmMxH6ynwKrSCV3SZ669ra1wRaDqjRHIQOS3zc3lb5
dkJF2rdW1fhR8EbWXViNVRIeG7ReSL8XPp/tgqBzXRFihTx2twed2D6+nKoLFT+V
GZNZnld52t1eioswM6nQNMFdJI/CrADb8kytqsM7B15OOHEdunVFMJWnLm2PI3tV
wJR9mpvxHsU+RSQtjS7j8ZfrI2Th1TUxNtOni3W2k3Nts6sYlsO3sbjXeOVHC8u5
mlzUXQmIYPrjAyRO+ehhSS3xpBLbBH1N1Q0Rwr9Dn/9yAf5SDhfeKBLYZA27ZSV0
XQ0yxMxRoxVmHpW1HMu5+dOncFrLGprp1iZazb2raMWtxIz1ggbMiS2fj4GyelwC
eJ6wPcvIqwqogzKXIA9F3GYpivQF4n+uw2GHXskXMu+hFASJVO+rHvuettWwjOEh
OLonpgjoveg4D7PyKvv87/fXzCG3xdEaCbUMb1hGYrK/qVWYnsNynS45j3KMrnlL
R3wuy7xnlQD82CJ820EIDrTMJJgyrZMFEeq3T8WOAmsdG72OodPyESqG6NSTpdIx
8Dvcs5vbxSuavCUv5x0SnQ5dExPS1aUD7cJ0UCMtE8y14XIGP1vat+BltsnIrb6s
2CD2izej4ye4e62ezn29A1kRJuqSwAC47y724zqR1/FVfrmI/hZlAGnuw422V3qq
rH5/7KrDm17N79W6bjz3Xy2UWiPeiyLIIgAHRHutabUOFkT46XBL+W0cKO5y/zCp
uDUc3AhpuE668i+RTYCBI4BJSUsQdoqdwikJ8kfO1hpSKcAN0+TY5gnPAjAPy2oh
5zGwK1Rfj5f30GtRMgoLvnKQw/Xh37Im5+7Po/xs6Zq8cCeAVbOs4W5z2UCYXcdm
lgLGxVYYtq8KMFk4z9S75qxVjsfOLu5aZWzF/Mp79p0nGXeCXV3ZHtTLGIRfGJlc
dPGLkkuS75CNuw9uZz1yrq94aRZkI3h3JlbaPKozCukla6EjgCZOkfY7ocMely+w
WnumpUB09sgmv6IhwlRf3JkaaFB8ci4aEjfTTYxNF96lZax5bu/nsNR4ibTy92IN
b75xz3vD9vX/6xdecRvRpNnr+gXuT0lRi+Fparf7hJS+Ssqagd//VF4sCclxmLlp
oV3mZthWFsLCYug+eauQKOTYhEmJKaxrXk9MSsdEr2r/PNV2O16ehkoECH3IQyFb
5wflnSThWNPFG5PWaZmFP3T3UzVjoqg2t4xWPAXseS+EtIKy1DHSdhYl+QuBb3ml
mQH5I1gcYzT361hy79YZBqn+BMt0kYyGPjWA+8wICwN0eM7DFMhRh6nl+RFUEPvp
ECOUVMXNw9TOT1QopHI8SiLc6ekKGRUL6xfHBFs73I4mfK72zht8vIiEBBIUWOym
KDP9knHWwi3tC65aYDXgFjRiFnZsioj+2Clyk8n+CzU7dQVF4Kfi/mJIiW/QO5Lc
EyI0Xk+D5TjEKKp1/ZwjAQ1AAU1wzPtNb8YXyNete951agGynfLNkEvraE/DN13+
OkD41f7wd562w0IeJ/IFxu4edCzpH9qYiUruG7voiYL/fRaQXVCU4U5l9QPjkRxK
xIMyH+QPxM+3TCTdDmexyu04HA66ETHRJtNjvfC/IV7r8m6R5XtUCHTTh+YZTI0W
GO46lJ+dh0kC6BXvPWbp/AFfKGDYvtvQGALCgnP6YOw6ky8n586wdx12IJC7s9nv
PiyMURoxUa7I/zVeeREbaHpd4ShZOcbDCo5qLthra+um7nQ/yivsHu66QXw1MPAX
JqfNgMo9SFL8mqJQ5VEl2OaXrvRyHjCkxA3AZuOXboFMRR9bmODF5qGH+BAOOlcw
oGssjq26Q8XZNHSbiZcelztLE7VVPUtXLP5SNzvceozVgDKYmnnxHFnO0iF9+apr
EfcWCBgI0T7zSt2LyjctcEa/GTuyxm1hlxYNnUHqxVYqnJl0WyPjAV9djF02aato
nkGAzGnxVMiS2PoNoGu1UON/lgoNY6Ya2+FvhbfS/2OtPfS8GZnLJIKAeoazwK7c
FQTj11qT3EsP1mfwR7WJVYhKn6QJGqk2ctBgWTPTtUqPU8Hf1MFKIq0za7VGb4Co
hOqaxT6mqRq7+avUAJElmzf/flw7Q0jrtFoLSHp2KRdyEhT3GHb4xtA8uCufDxID
i9L3/PKxm+sYraQ7wsR5zNFQJjbp4qLxBYGfVb9bpzJyZKLKdbd+ClmWR0AcgVJl
vRLLqXmhWJ2uuyhYyGY0dw7ePESkiXOzvtgqGsCdcbVP2QDTAnU0xhagidR4iSXm
dMurKH/YREYe4aIWvYmdZhc9sbSKMC6AUPpQUNL1j9m8uGyosuGP4WcrhKedMZ17
zXd2iTe/n6HJYkiPjxYrDNvPT/DIQ+ZlYTxm8vgArmqOr+gx4/ERGsj8nA//B8oS
thg5XDzil439QVv7fuOQoV7PxR2rSk0dbbhSiKyzVywyMtdeJwuZax9p9v0l8sZ6
A87lf8tfXVGKVfkUxqL5YB2Lxzubj7Xx73WAacqT9YLgmrRE5EPhsAbphGFQ9gOw
OXVSeM4hBygLYksX3kcdviT/8woaSRJ0RuQq7tdC8duVTblS0VJ/l1C63yFzkIuO
14Cw/k+IpTJtqOgOc1c9eqqbonL2qn2JrcHj/M1p297e4/lmmHI5NuRAI0BKrVzG
AfrwSG5wRlUrnex18+kgEfwDUpJ+UBpbUjPX6DSCf2t6zBOFAbjDGjWKSRhJTLim
97bta3kCcqDIjDZDZX4yhYTuDnwXEqG1Mhv72r8C4FwAaU//S0hvA34336W6ozia
1ZV88pQQdKY3blee8zr9vlW2Uxih27/KdncTf0h2aSX457wMFH8UmbKuVaQx41DN
oe8aUz5Sd7jXN2PuzhLXMYc2Qh8Scf2XR7SGiJP36sGfXoggGLV4xNk3XmSg1ROx
Nhav8bWajLA3A9PEQF14s8IJiKlP+YIyJ4Ecnn1JpJoIha+yqJ6tQ2oYmbRnhwDZ
7jOu3KjvWQeLTb6jb9AUZZtTkXYqfO7rx0p5jrNpaCC+g3k5x1NKmW6ri0PJSKJQ
9OHoMtc3oUSntaf4TBXs5YUZ52vCZ0f2MD5U1YaT0NJ/OU5jNnJw9O1Ms6boEPl/
5OCadLmee7My+XoQkTEnSB01fsOVc6QFXlBJUkknw86iSzMq4jo17W+IyuX+Pf7P
m9va3TdiBIsnePX1YroOSG0bWyow+dEeTj5uX01bgNKfeIKQ8uQlAdjDHfK+zHWh
d6MUAJNqxpSRgQ8Op+UW2AwbdPJ7o6vJV1ytzDoK/WQjqi1+xGVCnHfleziZ8lt8
xAgOFmm/0o9Z3wPqZ+pClP59Ou82XhzbrGz+SKqLiEhevlclZE24uYzompKREVnB
0mYJR1foQVeJFYgiHhvvGHGoHaZRHoPFqqfsSmqLjjqtuJohVxG11gV+l79xJDgp
irXqmZ2n1A3gd7oTJaoabE+M0Ne+YaslW1+verPhsrXO95o/RYvHhNci0Hz9bTOY
iIISllBfZzb66zlV/W6QgeAbdoFIxDGhPEkA6Zoe8V+Na9+2dMbpx23mqdTQb+dC
sNIj7fNgXKdkXS6tA9BBtVUuggV12cAmIhx0XTyVm/ERmPzZRDGV99CABKvVxolP
5j3AW4glpGgB/IOsfh6GjBwLD9gHlhHAW179OnwxYxUF9gUzepzwXBZcIW1FfZgu
2MN68NMN6B3UpBPWQqPQWYn5sDiA8BNKTUUNKFCz2RTGkHCaXx0XENTQ7NoN2psL
3iLKdzA+9P+vCv6jVJVSVKwQuePJkkwzu5MoU2HEDeqqijzB4BuiRQJIZIkbMZS5
r/l+zDgRVDaqcmm19hciaeZ24DwOnS4b1Jh/wGHJFMyFK/EK045tsbfD85zDSrw6
9xdUCjmYJsTSe4bX1GXLQfZNhit90poYV5XIqqG7hOLkHXg4wO2z+bI6vKdyJD/7
3BvRZ9zqflChC19xBgnO0w54icvq5H7dZu05JGUstnmaZ3IIMfoiSG0yVYcqIGEk
ylczBW9GMPqmzWyM2MyqquhMgkuxuN3u04X1UkwR4nwe49/H3rn5ukkk8un8HiJL
LcUzwJkcyGYktYkt2SIjXf5j9dvrDUWo3TqZYWfaYA5faURJvufMacQbCdKRzpqE
ZVQDbm/gemaxNI6ziDNOXj04ko8LH7si6DKCXH3c+HOpPOvCsHINJ13oUdzBotvA
BH+tHktYdGGYGiP1iMguPf7asP/unLrVVMCWXIt7HbFVnKRm9PdrSu1hukw/c6PU
evM0bvMx4Th7KzNDUnwwRg+Hfg/OevzBejeJG73GE5giuE3Sk0S7pyo0IspOe3NR
8OvvlBW9EoIXLbCm23PX9ZUKXELOWZkZo/2tMs9LVrQwK27/sqg8/CvPjr9JBobt
N1da/Uf3iF3ll/iQn6I5sTUDt4lY/lBDJWwiZFPFE9fg2yklZa7X1bDiJVTiCtuh
EHqoY7KHcWS/TSri2DN7+PR09U3IQE/QaZnwjRswQe6nzOKjPLZH2VnEILWDc7HN
hYNC85w1DAticyIis3So2Gg531EwzAF9U/iX5MxfLDt6ANjivc2UNUWvcbIMP3oc
XQkgY5lCgor5VX+z+KdNiaf6ffVdAf5bnzdcYVJ/5Qm7HThfobCKiq9AYK4qwUMo
fAf/8JWEe5SOMHNh6MZjwhKst4d7TJKePM6kdhYpyBPWG/Bx7Uuaxj2fXFFO2VjV
LjOl82Q/k5SkfKJHWEwLdPAs5rT331A9B4OPttnODO2jb65+2PzOnPrHCGiJeJoF
+dxoEdyi6Oe0zVsqzu5evQG5ALOP/Hnbpp22EOKtPywbrTM2BzNJ7c5z2ir2YMTw
amoHzPboW0F2Nl7jolTfqlE40JjwQQN9D+Dpb9YgfDGlvSiQycb8mMbWUCHy/+v+
UuoUGIHG9kp/0bQ//GVoCclJRm+gu6qv1+EX1oNn8a/JCUxwM5LrFlT5fRXg7d5d
zjPrfzDaj9m6JG3+TBOHiGCljitmCmRl6ObjNjfB2cIx9DorKUL+sZvLlkHAjdKp
85DRkRuIR4RjavSoxaKp5aeURAopR2AIsEr1atFgj1s2VxEBqH6M5xyNQU9d+APH
3HC7gXOvvBw3S1B5u/RzCH7pxPZmYo0VkNi+zTTYFrx820xVO5jR/cVRFL6eqj4Z
6i7I42FoZufJPd0VnddxgNvpbcDwwDwuFAva6GWL4BExJyrm/4P/+4MbVAVcMya0
c/YUAuKhCNBCSLbfZGRBSO4Fpl9qx9kb9VWTcScR3xfL0DkphBhnLrmCIbn55aNk
8KuHSeEjNL6tqVrzlXb/Ci/OLlwyNW52FiMeNXYf5mDBNSLk5JcHF6KQnfTreo/1
uTIrLDgvo1X4gJvjOnjqgoej0pqMrtQ0GkuNZRS5rStY4cFD0gnoUc44G0VDuu31
Xb+IH+ha+ksAoF0A1t1K78fVTe6bEPr7K38kZaYcE10hDL2JAdyV9jt+SyQm1vI1
XMmNJLHxiE7KmmUM1CQ+vCmibRcwFys67GIpB+zVymfRCcyuCY83KpPvPeY8ovBM
+zyT4lXPluidSJhlUBmnZW5UEfUsiZ0GpQEhuWlw66Aqr5L6Xr9m6xGKWCKAlhgi
+PShGhnnylSp911Qs1Cqrb/sAjUVWKHLOg7hdqt2x7ZwwZ8mtrebe8f94fOx8YFu
SrsxTV2avVGvdRR0jxRzA6fMPo7n3lxvWdmu4naTEv822J27ULGtYIPsvaB6eaLo
qJX5/nf+La24uC14Nesq9Ggw3yybywLucVFbO8YSXVYF6a8KPSbwj2THMqK4nGGB
guPdAZ8aXSiStC8W/zU8rx3IkIKcNPyh8L244qI961LYbsCoDBKt5tPwdUrpIxKh
a12nQWyTibKmpN6Wj0vG5gEwCeU1vzY/nPdN+CmczM/jsMwNW/wtMUx/+qdu//3k
HusNZhobef91Pppcb0PfttnJigNOwgU9v9EqnCSif8gfbTWAZgrIbnkdZv4dJDRT
W9EvsnxRMbsEMHH4TfnqENtbYkvm+dx66AMmd9RSG1PeVLIXTajQtgX3tqTyz/1m
qIoZ4SluYTkl6/jtYdC6ERITS0nTp7QmdkXVSeY3WUSWoOzMWnCoaT2Jonits+HS
j6cLw8JUkx8H0HlLyGwu1xfOGL9o6zI3QnAMZOwPXyWvuzUi7qGHPjEjShIj7Ahu
FdGuuWA3BOVTCINXzJdXY8cLA7Rs1RED3FzaB1z2AbEJIggv5/HsbEM9xgOzQmC/
HIVD+DaRMmZR+ZSyWlr2oKuA8cKgW2eBL/1mdrImysSJah8jvUZ25vhNJ7zN5gfr
VDfrV/yg66l2Jv6QYFq9DyIr5jbw45f+d/Vrws3JkHX28BN0cfrXFRyCpV5HEeZB
d0lq9QDYQhZ+w0tyx8zBRJti7+GThTF0nusRDE8pPtuW8nP89bDWxvktqQCq/GjT
jAQhTzlZ/yhb+EJArFqmZMHj/2Vg1DjSPYTwB1ySCyIgafPbRwPIJFhVOI+uQVOe
36hsKdwIhcSmI9bD466LWwWyQwxkt82NSIeaPhErxpZ+b9jf3r2khwqUbuLOlGpe
A6YAO5KHbZ8LZdmljc7MZQ7Zuvd0UY+HDicxXpOn2MENhD+xlU8m/+DGSDP+PHNW
Y+SjjsZp6t7VTr6u0xXZy5QbIJ2Px64Wmm9Z9BBEX/R0/8uWfZFd+xf3YJEGa/lM
VO4F1RU6AYciam14BmsOmidhdn9ssFS5E18PVAoqFB46iRoABUNJ3T/58w6Cxgx0
ah1JHW5Hk+6+i4Q0jmH5pc2JDEaY462mhOl4oOgP38W1qWy4GaKsYxq0L3LXZfjF
H7QzPJLjUtDQAPcn2re5dMeo7NZLCgZWbABxVz5xptC2muK0DbVk2XR14zMhK5GD
/eysidKoG/L42ODKZu6TS++e6tCoXSKtezvtbyYgYTmTFdvvDnEI8w5ufnxic2Dx
VGuc91Atr3LHPd25RAMx62jOWwCTiQCFZPcU0WO+o6YbwnE4ybM+3IGldcWxCwWI
AKpJJYCi9Uctl0b+cvTqvMr0RMBoM6I3zSPzTsIJCBWYT2/t7EgofVsi5EhNaI38
shMcMxK7F/rHq1v/O4wm/lM/xcKWC6R0i1wnMlikKawbTRav0hjLvCBi++TIeiHm
DmC13bZHXKfrhUqSzbw+/UjuWb5lrKvDk8dLqlW5XWateMZFGTJ6cFR2F0DJvJls
qiI6mV4kxO0ibwvpIKyFJvTKWSsB9y7/wiQui5RYxW3GQZ2A6s4R8BE1UEmQ1Fsr
1bR2mWBV2IgJ36F++e6P2j1EhU25oq+rmMZESkiyAFcbPv8fR3gOySZs1VN145wn
X9bgBBcvsymC/Jishxatp2BUiuoC5bT7LBAyuT9uZBn0GHG4Au4iUywoKrVylx6V
SzlsuRYNhFgb/5F879REDp8/JAwbBzJez8Dmq7DRKGJTLIpLQMvTXV6Ta9s7GRBC
pc/DcJSkwWyop3e24WZUk1kHRjElKdLsoi35JmRH66J2FqnmAKvInRqHmBN6NcQN
YoT1RZlYuG1+nhvfwVUxhJgkPmPoCQ694kzKx57aYVVLMAttnn+FpHmoNNKrnjZn
Y1iAf19xkuPoHeIsIUvKSsrbBKY/ljmhiGaYHgsqPyZ+fw+A7Y5o5NSwZdSzM1pl
uef0uBEYGZbRxCy+fIZmo2WFn+P6J/8sqSeDVIBRTZj0ckdidopomitrFi93Hli4
iKNI79LjMtoM/SZJAPKeTbBldvrndmSH6J1UL2emLCq0Z1D4qyxSml86aeLcwv/P
3cBpH3G+B/+thXjUfjtT+prYF2EzAbtkDg3ynOMkE18a0SdlfwRe/bNFCLENuP9v
HqqcOrd/3WxRT9kuxoAVcpPqClOH0lvQSQiSZqUR0wrsTjUNIX3j8gVv350TST1D
slHCCrKeFR/9d9qXjANEEFHhI7FYswZ9lVSVIC1KQBK1IWCRzRdejWU1UlSSAwNM
/oIM8PaEsMfeEtSba+nPQoXD9Yt2aoMaWzZi5Sw8mrhXjyZxXNQ1DF0nwZed3XRg
58GbEvo75Ead3Jfone4d1ZDupf6UcjPtmKqE+tTq+6kyK+PW0m49sZYfPRVoZgWh
/2REu5E6Gg/eE6/JLsr6a0ZUvakD1SBG2nb+RxspJKapS2Eo2sANij+zNRT1Ez26
uU3JYCTfddlDkU6kfrZ+RaScccQctgtzAmyeRHg44xTRRFwDaIpsoVp/w8OGgFbo
rTADuNYLFHPQufVb1HqpIuQ9p2LaUwTiou3TRs2jjfO5XP3eRodnMkL/dOwEnXWy
EavUflriI/57I17b0y1xpdbTs8fqVdVqBEBCV5qB4K9qKAyR+yst9bhxuxZEqN+B
eCt1HFG7vGFegCPzSxMdTm8Qn7UB/ygkEUiNqxP3fXS4RUEMlBkSZZqj/5hjLr0b
9P7gIuKvYi7YIGY1RTfXXMofNMaXumUe4N6Kk+1DdRYshaHAPv+4UqCle+runVWc
7QOuMJKSMeEUNpqdffZXKHqw0pyF/t6+ttjga0psxOCqhhiVkxnF0cJDbb2RjwKb
OCylh8XnICjMWi5k47dQGcf9QpSGZfYgpL0pnjTEm67e1aI1NnYRNzUE8uQhNZfw
ssHgL6Let3rFwgPGxzmeBKgFwO4ltB01T8i/CmbFLB+F4beb1t6FeOm5HQzexXDb
x5gIMGqCn9PvFIN25rkyo5bEsS0bCDKR93k0XFBHtOBucMgBY4y39ERvsxMfXODl
YfxDURoxGB7wkqkh4K9wQoF1X4R7rB0vIkzqHLT2KXpvZdnjacaJcyldKRSJdqg4
xVDTDxVf3GczqVt2Nx+bLI/YSn0VUOdY9WILh6slS7o/s03qppD68jiR1/EyYWLt
u6Byt0v2trg7ExydAZ+K9aazjpsU6vXFo1558yocn9Bgypn+6ojYL8WGL6VbiZL5
goRPL/fRg5pKnk8d4iQhjUsnFyeT8RyuC35P0pkTgIfRWHQxBtc/RseoqxQf2Dod
5nbLje/oAhWgiCIpkDZJ/ys5lpcFnu6GKHQrgABvM3vtbBFDWyBM0bhaOxkJ6M0w
V9TH+az0MWHtUKgA0pkehRw+uh9aljRMbZRW1eWFZZ9SbCWmim3kgjGp+VlQO2VL
6rFXCnpkgy4FpfXOi2VINdzYi9e5u+I7WUwihL9/PHYG8nDGSeTsu0TcWAOvp3jS
rS9J/2h8M0xHTJg1i1BrhD1WtcyKOsPMCWsfALwaxc23EsqE2nVpaTcI4tG35xZr
9kXD3pecMc6LIHkuFpyDw8RuYjN5W9l1JN0fBPefFQYEmuBdWTZGIpAMDoOl+k0y
0NcbF6T8tNzbay05xQOG7+HtWTsbFoEeKCbq32VYVxDW6Cm7kJjv8MI2yujgJQUf
p2kcW2nVpDmnoBIAQmz3M1dDEo3OsYo58c+byBWaM73Sqq3BEHXPdOtHiHBPmwqC
X54W/duWETrf2Jqp4IbqcSBAvzAs2lzaQTNPIYq1q8IUJtecWE3gR86HsFsD+XbR
YsXPCWY40m1y1+kzmpqsKfHbjpz9AUB4ttA8D0oGFT2HthJ+EBC2hc0ZZ87s9nWo
19M7eX14c7hTildHQXwJqZAO/r2PoM9KvO1VCxb3Bo/MYeXOvAGULYKT5XfNbR9l
iRr27JznA1FeXI2698frv8x6PR+Mn/rkakh9RAlgx0nuJWptqFVXyhOoXxcgOA6o
BAmpueUFw9/rW+Wmc/6geQKpmF0UU/0t0wSXHbH2LvJb+bsZTZCjHKNKCi1Pki37
fGFNUA3Pz14sV8kL9veS5ScIKTREib1bT2VOQliko1DerLfU9bk1/7/x3gDKOaAm
GePEdenZtqJlgzM12/BKHHndzF25lNRqcZwgEVSgFFfAdOjh5pP9ocAZiMFKzWj7
wIS4unKjeKVUq2W7sbWd1rBj4YMgQFX4HelNv3WqRGqmJEosHsn0kqhiSYPCYhKo
fTX+ty7C40oq7wZMMGYrp/lhNHwIrO6W6Gp8VeMy1YtPlGWGzcs2de88QU/WOjUQ
SLBEHhbpFuwdrMdSWFKyBnfiMYFMXw1HxPbdMrvTxL1Gmn0rOe2RJ557KGz5+IRM
XcOwLr+//DuN1kihYlbiDRiJhdfNgSEXsuEH8HhFxtQ5EjhiKYFvyorXqvXV0eL7
dYeCT/kuAzl/DDLOv1o92OO5NbQXNQkVqbn1wUKvrjGa7uelEXsIIdaxcL9Vr/eU
pmrbJbhH3Ujkv8FX2ANiLKBhocW/f4O3EqhLWmE3HwO9YGoQEyLhesC1CU1UVBUF
Ep5S4a/e0UXOPwKx2K203xA4AVo7Q2Sl85wmCl4VltEUPLOMC0YBJ0+ewlCfM5H2
jgGEm4vjorgtCobFjwtoGR3WL3L7BGG53yXMOVIphwhHEXhHoNUVqz3YJA6ui5ij
amhSdk+1ygHREpQudYf+8mCPAr9PzW6rDVGrnrWBkT6/OQRP8q+9S2ZZP/sKMHoZ
p41+HsBz886twT6S5Mxyo6k7G4ZxRVk21OCgwt7adykjsh5qIiPApQ7EvTfyRkmO
55zBeyslkYgVOdE76+Xs9D0U7pihXa/XpBXx0ctGh4a7U/HIGTy4nhW1aeed98Bn
wkofZIoKiPRME2UNXIDtqruh3h3Sa4MUkapukjMT/bfuW5Dngx7egM3GQyNImSuz
AXhM33Is/Pt948MzwBl5DPGhiHy34M3cpUmSplLtpKmXA+Cnz0B3a0oZ+Hsz61aQ
V3jPUzNXKQIFdNbpqyG6IjubzXtMgqzlgsFVl2cjBEQkN3SNObkPZiNXlyvQQ5+h
W3x8zRdkPzx2YGyWxVcKkDfAaAcvaOJSwn8diS+yEFEt37yn/X/7gV3I6v3X2zkv
c5BUVfsGN08mCvRTy/bl1GuJtexOpQK05um6gbtof46/QphiM9ABvUREW8UfPAE1
1/dvxl1twZvqI8/U8eoXYzEln+oD00V9GRDPbkP01SP+XIZPlDIRyoJGofxC6SWp
dBwyYiBcTIaXEpFeI7m5RlPSKzBbNR1I+TcV7aDC0442PftcVey/FvXPNqCRcNsQ
caaTevimLwbgLGLcsoBmfv5ysSW9ZWSNQXDlFhureaV3MOgS6LNOlvBtMfVThdjH
MQ56JJKEln/iYHvoaTBoo215OdhIIORidwx3D/sIWm0NfcJRWHmShx/gpKpZilIr
RftItkVD9cSf1Oy9OK3vXv0SL5ozVo4alRHo6MAnm57wiVUP7DHrz1IWTINqRIti
QooJbw2HU15Og8zt06rmMt/gPhpBsW7pxi8LX05wg/XWUG+lrhtFQ1q94yJmn0CK
ZmbelE+WGjInKGAzKs54MkrgRKCZ5dNX5/Ckzeq6j2XW7wxNFnWqI6txLIM8HBkl
HIlT+dbTLbmYE8H1gehfr7ttaYbVg3yEev6ts3dHOxDKL2LPuluw29KcsrcObtUt
tZjnpcg5ZfyTGRVHH3wx0LGm+HooTbFNg7mMs/uZsK7eSpQFkTjqgWDzVTvqNxtd
pXzzM0r/ysspxVrWwb7cM8dHALzFSRSQmGnzAlmJkB77agqsA2dJQq20eU7hOmum
keLmR6WuEm/lQEgxEflp6+v9WeER8/gJE9Evc8olaF6IASEsglK9LRMLuwGeqxlN
tyNLU6VA0LJ3AHc64yC6B+fWR2b7jamiAUyOkVzAhKlo7oMOBWmkQjIHOGfVcN/H
8OXB6n31UMhJFtVZEeSu8KLoM5jLG9E59DJ4wSX505rrQsiwCf1nG13t1/yCa4bv
tTsLodC7iUde7MeIxm/zjmTzy9OnxaGcEtRh6q3XixKOMh7XwOWNTJJNK32Jdiux
JUk1EOf/9QJsyJQ2bAT2XVadj0aw/R3tbbcqYeNSvfvEY3V13LSBQV/SaWLRQoLb
xoe78qB+36nj/11vfgdK+OI1nNykmr6QuC1NnhWTweWCK9TFnO23ILzLkuEAyBpe
X9JhA1KdrbvK+2uInOKIJqptXNJOHU685dfQOnatKatVkXZRpnQ0LwWRgYu8ELJQ
2SFPoi/9hAS9UDCAYJ0C8+srNo9hVTsgw5xzQW8XsXHNB79ag2ueOdlhddRS1dDC
+Rqp70kxmnsEk4xM/K28lnL92eK+8+Jzle3mU0MAwS/xeSzlx4o3s0Ocl93pmv91
RquccmLHdCJKsuzFV8H4b/pP+WOU1b4vcN8DQPcbeDfUwKvAVga3ZCNkKMx3bJer
hez8S5GpTXyCrCu5jQ39QEymhSsUwjfjgsfV1O0d0/E6zPRjsnvYrMkwovcNtMcT
zMvZ2ZFtFR/9pUNiieO1VibKSySdvkvWclbttLv7upFhzjSW7TbmoyIKK13uLMlK
TDgeiUM62H4T3fMOBjfK6MJYvVSS5kPPTRMrcwq9OO6YWZjOTt5R0gXy1AdQA3tm
f9RkRXz1Ctt7LgUkB1aeNRvbpj1rlPcHmk1Cqnfxcpepb1YkL9YuuGjQFuso0U7I
LD7yWdk94NNAl44VEK3Fw6x4hoyNBG4MU42M6yr8aEiBOr3e0UaifFB0BkmstbjD
K+/pDkMYeqUTnty56IeM+Eq/9F5tKZHtpKrhkTusvrY6HdePuDC1EyrpLcuB0JHi
FDBYto8xqPYmRtnLqr0LCpgcyg4S5yJCqxxKp7VZs76+Xm1KkvAtulHkZ0oYPy96
sbHDVsXPMbeNLJFtXrXEi036lF2bRkXbjoNS31GaTU/aEmXKuw9GTbMgo6gER4Cd
rSe36hbkxeh0qVNvm8H3372dzXjhvKDOn8W1/oey4INA4ZVwrfgb0g18hrhZQX5+
FjZN3WcDBNvI4XCNS/ECZF0V5AvXFFVA1jtDCPc+ZX+c6OwK/P2BJTGB/JNCNWbp
mLdgbNd55KwPxcdyTDSWaxvzcgMLY/hsJuVmiU91QeyODTxBmGaV+wxrp6BFPeuf
HFArlyhH8v3sIDka0AIilgMheFEx/vWeFy8DPsWm6+F9cjcgg11zNNyuaE0q6DfZ
9MySknoD5pzHn6cTYcZfP3932hQ88cXvXWYUbPImqWnf2gQ9LBZ2e72+SMR+sciy
HCe187valrzYq2qbZj6jPMn0zfV1097IfWuIRdwz5rguta2+BTz7Kp2g6lzV0nR0
9ZJ5ePA+JiyIe1+hu056IPWyX2CUawOLtmh1yK3WQcarM1USGbHNoENnaPSuZG6S
MSMzaTlWzjeSb3ClA0po89q7YrM8b3EQDU5xF8uW1/vbVm3yO4R/p/R8VRPeULsF
7D6HT6pSWvuH/5eAmxD93T8D7duf1dEqoG2PbWfIwiq/uthEUiBi4fqH1dykSqMX
LlDWKcuOGPA1QyM+JfxMf7X4er8wPwy9aFqIZ1YjRSIZtyQK9YMrjTq8hj4lnqD1
3OCFwzvV5D/4AfbxEn6sI2nmeE7RMxj7AqcUJgGqpErXZehq7MdMR0dWUm0bXBo9
RcZSmpAIBoezfmj6xlDiTy8ujhiDFloP67j8jVtHwyFLZpA3ySKdyX6T3v9+HuNN
pqiWj/Ph8/FT4Sxj6LWZR4GzxhjLws23MR13adGVq/ECwey3yDoGwR7j6YIi3TXV
vFZSTUqbdewLADIH2VvppaPLzDecDov69HIJ61Xptlm3XVL4NcEXGHbJ5iFqyl7G
Xi+8CwZXRThm5bXOTJnqLpt5q2/X2LNOUEZXLBAgNndOm21cMH85RYtsJE7wh6qh
CwdISZoXOMvAgkP+/qLWQF2lyMR2Zn6M/2XjUIKsoWeYWtmULK0+7jadq38DJsXh
yt9r/5TmtiGkPDzeC31FkJRLECf802tDzDuabcupP7WM/vrY7eJXBAVLHtJA//TM
DBhOZNkysTNYRZxszhZwJIoexS5QJdDbssZfHsJ0Og0FwW0It8XPV7YPZyJq4L7v
rvT40wd+R9/Cp9nYEn8hfc82/UPH3n1/oKKvPe2DeaGXJl37D4VuozrVLELVWF9a
N1nTPl+TZR2tnman2M4or8Vq64NimCoR0GJ3pxC5Z9uAtXZVp+6+UIo8dK/a8Rc8
veFKk1fD7WBtXJoUUPQZ7vMCyKZ4xHtWCXl9bRMw52QyAvs/v26wbQuUEpOS65ZM
yE2sDjB1dpc+712c5pnIhw6Jlbq3o8CMIXgsus3ZZ4Sc1cqNRK1SJ0IgGwf+G/vs
6i9HIFWTs++gbMkWhiRfAoZJ6uXKOSCJaHnGdYR9LNPp2av0AiaqpEJs2kV9Gfls
MC9yn3v8DftTePpyH9ym/dkbGMk6WPB0gwQjHGhu5SRh50y0FLu2KW+NBjQsoquV
YO02p5xBctcpnMpM21i9PIxy3NUesLTOnt3O7TI5M7nRx5mVe8ek0ER7prGD+DnD
n6FdBdeRZenW+1RfXaMb0Fr89ciJDmANfqFieZmM72/EHe/1FkVN9V7kX5yIVqBe
OV/xLM2cZIDG1/tTxLuOhErrthkjr6TRcgxvSE5/wfJYiMRuzt7TwTWRFxoJcaRQ
MNOI/tn0cxm7w7koqLmNMyI1Km5/iG0ElLNbgdQvv/6C6JTRyicX35z9EO3BkR0Z
qLA+/IECT9/ZSW+8vkaAbDa8FjwXBh82dMIN1BGFU3YsFzCvmv1oNDV7O57OTp0s
bzTSYtW7EA9wBi0K2AYKPsQ5rR+6MV/CrFqzeY02+M1rgnB5zVUh+DnDpivOucAF
XSwAzN4xN9S1H4OFNDQDq9Jglda+k/MyTp2juGu8jlcDKnU/MH3UdBkuHCcLhBUo
UoJCpNFZxukYYPTSP0MxPtY5Kn8Qx9/O9fwvhEbdst3zcpIz6usN0GUOTugKjN8H
KYFFBrYjYVR37CE1P4a/1zG3rgMF21BsOm92zLP1Us3MayA4T3Q6MMtqKyl2twDE
dVX5wujUEiYVINklY9poKgTvNqUvYdcT8k8qbFjA8amGq122pXdzJe+Ic6oyYlhj
0oCB1wixwJWBnmtaQs/r4aPY8vz72N/pJ1aLCCI+bXHLFv+fMjUnzQAOriV/kEqi
nqOCx+GrxAF7YBSQkESfIaaRBdYbWeVNPXiwPvKLPS4gJPUcEAqawFZel/y2aXEX
gmZM4EnajffgnHdgkU596lP6UPlc31NHJSmWFkOhwoybnPdiaUB0HQ1sWriPktND
nW/TiYwLZ++9NIeECVruXFTEY2H67a9H4N8Ewmk0ZWSgXM3F4FaSznST/R04uohd
wJZX69UrodIF8AHLn9T/xdKpUeE0LR4CyJIAl+zGfiw3T39hgulWmNw3PdlgELtb
2bUV0Xy81RIcil58i3bsCMsl61FnZB+G7m5NkFt8jaB+PMVkIPlxUjqHYpIll571
nnUwRi1HRpmeyTuKqoB+vkDNMbX6z7f3CVLz4rczjuZAeSU34JzzcRbZODHgs0LT
BLgm7azWyNWpnSVC3WwtJin4nSWfjMZ9LIQL2K3hcJRAxcUDR+ujXRaeWuZ/pg/D
2TeZBI+2xksAbne8HnlKwYuMrLfEGBtr2k67ClydMEh2wfXAmB8EysNin6ekhFjc
b9AJaJjJVbIa5yOjWKlqHEKPOWWRPzFrg4y8ztv59f6D9OD4yJNUVd6nsKkjmvZU
i865Pre2lvf773MdKCT88jCWjEGJUzKQ7tFPkaMzk9ytKIhfo1dny33o82iqwKc3
OYr4wq2tutSYDG7lmLvg1cz+EABMipTqBUClb6x1kWv9ofALbqTd0hTSSiG3TfwQ
0jHQAlNCN4jTiRt3I2vs2zWheiHykN5N2shOf7K2cABZ/E6ANuqey7KM+fN31/CC
RhjwzRgL+EFkA+DEBk0RaHbLVsRE80WuamWNxGziMiqzqRmlbeU+mQ/71iF9V1EB
Vex4YrjtRVGGHMqEzepZ6v9Zpc/Ved1TPJnKrMQWnbZykhgzjRHUDppRceJjQ1RJ
17TchrneHpscoHXsVY7PNfpRhEo9n007c1wK34Jjc8OUovYhKyPAek53X+/PvtU5
Lkc9sx3LyZpJeruJkcqdgytsH3Ww7RK3Lbp6Fxij+ICNHJEBERcjC28MNsRp3YkO
AwJpFgXuYiWt/qrQy/4d7/5ymR7GRC5+wVRDfqFSHWSNSJZIa9Ra3MS6k+XRuR3P
4XiH3E7j6Oemb+M1Xeztl7t5SJejvN3bW2ickIiB0XkaJZTrdt1Ex0WHzbhkgCxA
hwOGe1Ylu+fRwJiMrNNbiBukLdSud71Z0/iVTaPVGO8X/8L9K6JQxjgko+jy894Z
Xz58MdCaMRVMCsblD6GPG+wYWat9wQk/IXfdeQgh7bgq7/6uChf2Z5pWdQWw3E9l
TOkHplpOjtAfJscmEECZaw0QwDntDyd6GF5rM3dF/bTIu3jOX2+r81z8iA5VZdn5
NKuOR75HY39VAxHCZL9tSyoWp0oz4YVPeiZSS3vamZ27fhDJJSM1myiEp89qyQw6
//4AmJ0x3Wl0yA/QAuw9QxoA48bQtWp5ACQWd0KyPMFWq+ctD4jb/lYyXi1NXEmC
QpDhV4YtkkWslYLUENPx2PzQGXGIXkc3YbqtJdjJl1zLOWDhGTJa8+4F/Vf61Cee
0pwpP4ln57Tgp+mOGXcKbBbfPYri2JaisjFC+ZrX072yfpLMMg0Hn4CBPN6Vkjv6
EM9L1509MPNFQY5FolqeuhVxBdKnDXbObabVX833kM3I8QrHLLlYxU2JrwwkTG8T
FBrc1hvNinw2g4DZHy8UY97lbckQEXo4Xnkod9D2WK/ZMEEKpzE0sKpV5NIk5TnU
7UqWeR+WSA4UNsZLE4DAG9TDlrKb1An0fKDZTVRIuacWcCJRlJLbDUK7snt65Mdt
odWmfCwH8k8DMREBDAWUJUWgI78FRRJatBSw0hO+igLcmNIopVqB10WZ/2oBvMcz
HANmPvoCYFPNpKjz5UpQq7GeGgI0ko9G58BE2pdXKVzE44HEkME+eHs3wBScIFYR
lOjXl51iqfoqQPN9ZTo0l0zl49hctucqjLhQt/GGMaf2sW42s6mk+ouJG/bZhuk3
wsrxXLbwsDJAjg3hrR2Kw/UO+rDxyCSpO52Z9LKMyQnXaCxcPidWBqZSKVNCmhGR
LEkKo76SfdLxM+Kxm2fEvlrNBzjYOjrVX5up3n7L4/kz6E73MepbFKe5Kh1+MvTp
vLea5dV/HlRhj0lZ/IfWq3PEPsOHK7eTdO5DdLTf7CApJeyR4qNJVepvB4kYL594
2Z0B/N4ViwX4RFi0k3yHihNUbfsF+/3aZyie+ipDqx9mJpmQPCuFFLwx1aFD9cic
AU4vpmJZKeTJYmCLEIpEGBz8O3Mkz6n1nv7IgVbaJBEknlqfWy/xHuVnzMI72tPd
yrsumvETBikCndd4SL4VTPDVuxGXncbE65KekNhZ7Ik+F3iuyiX2e+cctKyWYPAn
ztHzlNvjuy5Oba88m/gl7uv7JBPajGrQh6BV7SuBB5Q+g9G9ljMFlpE9nsQhqM+c
jRzt4in1vqTBCdYC+Z8Q8kwF16FskhSU5S/+YmHB8xjCfn/NKD1PJ07C6b8JqCyt
FC1yp77WT1oWaWaqeUekndn4t2UddMzjeHIaqcJQaN6/MY7v2E9bkIKdBQtpUXw6
ry/FTq7UII1kPaKQlsJ8drsYTVUYCUS4sZjF+GVM9IkSdS/2mzxj/8mLs3sdigNm
V/0uWiD5AzPVh5rl4i1YAnasdi//in2dqXCJMNwl/Wn9DOT4o8W4XG77IZTn2uiU
1r+pe9xA06li8YW6WXK9H9W3nXV0/nCfGasjP00ZGFB5xvc07Xp7rT+d64IWaQ6u
Nnv+WM9C2ufVKO+mfw6Ff9iHEytyhjdaIID0dZz+XMmIwSvEneYLqPPFjfXbVzKn
mQnMem4J19q/Quhzjh+ug0DD7IeataBCRMjOe7U5k3JjPfn3yUu5KGcJwecJDV0F
bVjAZYOHAVhYaleHFvV6+8tKHsfCtn+Z5GCPb2xXjUTSPL7/ERfin6iniMUIi09r
vQvvpoyc/nWyhPHS1xOw8+XwhKcWW3P2NMHAM24aMNiOCx0KAtpYwOzhtWAi/3D/
y5bxT5nj5fbCV4YTRsI6DQM7Dnem9EPxHfkUfcIzfeL/c8RGBUr54hTah+h7O4jT
VcnyhcNbuxhOpn+GV/WJ4z5QwdJtH0Jsd44J/bT9lQy8eMkU/0NUQGYECm5KX/v4
FJG5SOQZdZXZi7xyM8lBYb8iiIJsrALm6kWQyZPTybsPJ8U6QblfuDYBvfdQ62Tg
TMzJeeDzcgvb+j5QcKAK2PtObe+huT0fJnEh/r3PrNM2ANj3ZM+QT7qPvF2n3v/w
wewjhYLGj+TycvjI9ha0Ij7ek2PG0spto6JhKTYDSIN5fRsemhiPvm8O0gliP4G2
Y2KLL2GVb65L4DCAJUCmxC5+movXIRgYAkSBpI0fIEU76KuUSyAl1FeMt7MQp6kN
smMpbfgMl6FqUpKZ1+XVG6eDmzTtlp+uw/k9udjJflOxx6+05XtvoBPPvY50pSCJ
fXa03qCS8UPYXurk324HP9zt1n8yDe/4skdK7A8aX+RC2fLbRmhfK4jEGLlPOb3v
krkkxcad/s5pb8gxo5yWYS+HW4fvBSdDyZa2Njutq27DRTyeuzYOAXcJU9vlmkyZ
bdDP3+kTqhEZSYtJB6Q9rKbGFog5Mu0ff2qqSrX60A6wNRTzRFV2Vj2v7KjC16Rc
8jxcUgxHUvf8Mq+BloOkWMHMcAj+KTXIcGMEUB/XyK5AS3yMigHXf8enJ7f+Riih
hogpT4NJdkDegm+UnHR7vZEtzH7pXalsxmqAgkUrBTAqAkXybzfFXWjEr+iS67Ze
x+RPpqrACiHI5bgOTgBtISms6nVISsNy3+ljNXlZ2ij5mBdNAQTPPAdZ5kE/wqQ3
W8D1mCP7xe0pAEIPlcy+S8xC4FfZ5AYh12IqOgDNn1BMLSvQ1UC8hky1T+8PctDR
gPq+S2P+2JHBglGGg134/B7PsVWuuLEavi2/749CsxIDKnz+YN299wDUBHoVI/eZ
XYCpgd8KJzeKkS+6yWub6ACa0EcZqnVn//nkhthKtzCe33zoMFiuPyU9WW5wkaOO
3psf4tHUvEwAKg4+HLNXBuoUpcpu7lImNdlgEozL2C6Oos1bgFURBkDtOudGOLpT
bEQomNUR9zC4ZsMyDowz2AWv9n44FXHIC97jTe5xOYQmZkf7aW1iJTNLl6RHFOmr
YYrlfZS7DHg6H6Dp8EAG2z9azxot+eTRjqbRk3kdfDLyWa9GX0/olO73UizGSXrt
lian7mOdjpAIWtIjAChTIOHQc6naVWjoQuc4RKlX7nSFBlu94vsegIy4itxy2gqN
Cs4amrJsV+H37+aOqr7UG3DL7CmWItOswVHyN8NsCDgXmsMoiPSrS+McjS4/obo3
QZPC2q/2GEZN8MxHE5npFrBgYKKKBo0P2Ex+oIe1BssU9ujdAFWE19HYeg+CVidn
SxKu8Wj6atcSddcvLHfVhlFJEkvAMySDfAN82okRCVySh0EkECZgY3XLwZceNO+N
tgUa5KjnN+TwS6zM7FfLJtmEQDk7xnBAIol+MVF7HtJFu4ZGlYxR9gNOPfzCwKz5
xPZYMj9wQlDdg9lRLuZz6H4MCOvnWMRYL2OJrIcf34t7wd4AwWjgu2173gByOh2i
kRjTZgN8I5iHrJtq/FrnPVy+6DxAXPQS5wttt+dNKDOLgHFz65LCZhnr0caK5I23
4CoUBr5lVqd542T8arIl6gOqHhfhJKLjjgzVdNQ+3HKSle3aiIP6IzFViEZbyzyO
CZm1bl9TCiNS9Zy6e416MvY+rYrSsrQFF2DyhScmU6Q3L4nISfvBHeGeE5yVTZjY
OPVVF2qpwvH3EeDPJgmTzisRRlS29qG2yN/vb4TDJsIDPpuIPGxvDa3svFX3dIRL
LGTPli7nPk01f39K8i2eCYuphvmhSBeMbe6kV58xVp84SjEEFFa/GZhXvg9vWmCa
PoUl6tcn0eiTFLJe8QZNDWf/OCiokBB0IjJ8Llkf6iiIbFjdqIQ828EWs0rD+ig0
kTd49GRko9/hTahuD/eCg7s97KWG8BVrCoquFiV/WZFyKkFALZOHgJ65mnpM5W/9
im8rnAA0QEJUCQ/gh+5b0aX64tzs44HrlDjrbpLLFGnXxVNf5xS2kuabodXOWHLL
lzGxAXoOZN4vPnZsm63Z6Xgzc2Fvw1wOlUoXpXQNNnG/4msyoxY2jdZvr9rc2+Ic
u4ntDUP99sWihHpzDbYhO8gcV4VB44juSjLVQ/lVgaarVEvXl0z3otMakz91Y3Ux
TtIB8r0RT7wspEXhAFuLuBIzAzGLfCqXEiX+m90iD6WIetxZdCjM6B+vvdvbgVCt
Cr5f+CewPqJGxlycE+B8JH8vSeNmswtxLz8609eBsdI4ErcVj3N+HBQg/m7K7dF7
hmULH104SaWWWpUvy7lRS+ZrmbDM3E4owIDA0wkrelnI5r+LMYFbvwDvLUWN6HHr
m/ohRcAbTBkEjHfcLBbswc9RkWe2+VGZnQOityhkF0nlRd1xYWO5ZrCVmhsXqtPE
ZAfP9WFuAOCaextvZ04D0QlksdYY4DBem5zkgw7COt47TlDCfHnRoxSSLKxgYCNA
yqaGMSl2kpp1dhwU1JwwHAgfFE+YWfuxP9qfCOHnVhOZqFULB9fmQddDWae3psYv
gfL6MatNUF0VAcXfC5nMGfCVAHC9KzVhGq7PCzoJrH7r2pc2N7mnD8BF91M4IsKa
KqDypuufzjKybQhD3O8c9ZPV5GLQMvlnqW2y6m3BNwrkLG15W8ap/UgjmZeswPy0
LR6aMEDUFz0AM3ez653ebfx65F3fTmWQzB3r3i4PKDoZk/chw0AJWh/x7DXIoc6G
pOnuZFBkDJSMgrSCCSmUZI7mzY0M+pAqz9fe+ZRv4BW3b5UPWJmgMTYa0M6iLWUH
6WwPCKA6myBRIB4YA1jSS/wyUEjAGnK1wvdgUpNlpgrjUewBR8xg+GGibhvcF3IH
opFsgwrBSYKeWFM0flKXapq7Oi4Mw/jOebJpqRIovQ4Ml+x65P/UWx4huKtprU3Y
kyn8SqL4CwO5CGQ9lZfXqpfvRpsseYklUMoTPH9sUR+n0eBKYKVRmZDoHXSLOlxU
EA4jFqG/ucXu7sI4N0cEovXfxSmOqyuCmfVUIlzrPdvjA7GNbukul6mouFmnHi1l
fZEXb/2MM5lRpBehs7+TuQsXAMSVx2NDy4PDgY80yQiXjzI36uQHlEbWaDubMSKD
zrhETJlh1HL8E8rLKnX5T925ihtIqdHyoLu1Y5XgfOlEKfdV6GbBN6x14NEn1n+u
T/HOxDi83wIY5c6BXppsbkKvjIJKxyYL4LW/wBBdQyEnDJ+1+zROzQsKB9Qeb/DG
SyaRorvtUO9DiTwb4n7qPwEBREOha8hRsCmyImgg4Zqn5amG6qdHFgdV2PAUsrQJ
tLQvbjs6P6/Vk5rl6YYpqoKq0IDsFZGdJaPeSoGcGR7eE/mhLgk93eyfwnuFTymU
Y5EAM7mn+JH2y6txHBCCn+936pXU96tSt1x8nrTxTkp4Gamw+zz12yB1BxHphAtQ
e3eZUP7ZLABAKXRuTZvWBsrDh6tC6Bmq93QpAFXpDi7XQv/H41G8pG6HxtEkDIrd
bkd+ChZ/NHmGW2Kkhfw7d4ApM8sjiFCqTS8M5kTOjakO236Ohnsp4x2WFQgsgDaz
pbAspT3foTFC4gKMdk5vHlvCg17DIFMnZKRoJ2QixFPuRqUF+P8QXulQp1kXVKm3
lI52+I75fCGDBWDM9/wvW8OT2RzuD9bv+C1hDdxdmgwOFhttlSk85UKi+iDcSOaA
j3fy5IX5dAq9/4H5vBSQdY56OE4oBqE9BLXc1TqZa+v7k9WxeWp4HOC3KMXQN7AP
Z2CNr2y1GDArDVUag4MAfm2400LwrEwwViLJTGy4ad1MMnDG6VdcDeDhFUaFyfsK
TbQg9OQbI5DSUPROOwZrB+SWK5Zk/j2iOQovvOLAIMwbHvyL3R6VTqKPlRuHkK7E
9+uL94MAlgs6u1JzyQLl6GiAmZ7hABJX7jXKSHpZxF8ucB4CI1pCcjprBahX8ovQ
Q52/4hVZx/xlSwZGbo2W0rYFR+MUXpkUbMakjW3JSMpJyG5rH/PM3hIuH/shRbDI
GEtW08muRJueGWX7H26wrdJrZ3JpsQVpDf5+acDed/QYCr7OODC6PWXzODJ4/dcu
xNJ0ftM7O5knkhdXYwCXlITb94AogpxOY0gTl4XSsXt9B4L663gRjYDf2nr2Yn30
SrLfWqIJ4TnJNcD8+dfD2Z2A+HnKsK6RzaoopH0vSbnIpelEKGpkYqCfbdDmwyUd
96Z0A1v3MPeAeY7ulZtxvD+CCUWx7YZintsZl3yr0UeL+SHeBeBqRz+sQDi8QCjy
rsV7pdzBZaIp76/epS79VjQz7ULvwOAVG0Rrt2qC1kFMDKJ1ikyzqN3ALYUahN1E
VIN/PixnFSo9MM9Ohk/Y5qbz196kxWFHy6UlNTDD9iL3/o3R3UF8Uh4dsI/Ivx5V
XqXTH3UdxUTYprouU7BKwz4Rv0diQwJ/mDtfpjCJ1sew0rq7oRYXQqwxjJuacw7z
WSe2ivrUmh4/UyvPPirJEXTSG03AouUmKyFoCtK80Z5X0rL/dqMLmmrFYX4Vb+pI
uZ8CXj8u5jcKzXN6xnwujROMJELUFphUkngoxVGLQQVKnm8CTNB9SyNwLu+9a7l5
ISXKnRwLBH9Xt1Rys71Nv4TIcAayVuBQJI7JY6rFk4CEKpdqY00ZhqOCo3mEozYh
O6Y7qb8O//1frdwBUON7TXOiPiPNZzMak4QBbO+QQO+kdvdXP7BffGixtMQNc/8I
iQGOhIT7ISzzaPB0uxlZWBe9kWn6JxBl/lahh+34wUwc7sEXmrLngTilv6K7r0FX
oXckk5VkiaxDXK2hCpWb+Ekj6ND/+DvJhHmV482m2Y077pTuE9nad7wFeUC5QYxL
uVoQ6Vl+jeJjqifFw2ODIDI0zGOwEWpo+SUnryP2PQkD0JwCJxzsAJllxEB6xYsi
u5g+emGWJ+m3iCfKYGQIZyQIaJI3HSawEhHAbjPY1KgrJA+1x0xwm0x02MqSmZHj
gNuV/r327f5XhsMKHAQnl1j3FpGwb8tdul+kdBfu7p1bNFX+yeZM3g6dzgzgeqWc
G1GfjsONJKxQVL+kNBPwye1lyGQ0imSkBxuPLkjmL38Ur8xg4Kh90xVLHaGmvIG9
yER4L9ZeQYb+aKRVBdIBxRmlnrixzs9XmLMAMmb/p8IWO06PcksZnn7XhT/COrxr
TCDRsOYYGdGqSaspRBWqyi7BZAVLxdxjHHmcm2fhjaXu79autq5L+weeOeYS9Rr8
bNuuayShlRhs2fhO94YSSsThRDTIOJvGt5Vq/XuPJPN6Xzd9zyYCtlRWQxaNtVcE
XTuyAB8bGvT8DdFEdoxw+GtygBdqtL3Jl9+6cWO76EBwopgMyd6ibilZ5qn67arX
L8wIsly8QxJbptjb0YpJgySkSG2WuqOKbHhQ6xNSgFzZ1UTWtB1eFxulU0wDR3Q8
2MtB+HuvNmbQJAYV5CPEa35BsfJxvzigQn/j8UiMEuvMk2NqteyfUr1Iy07O5FpM
QpmC/dY16FWLzDJN8EolmCu6rK0gFZR/31RoeAKthsi0k3lpy14KUv/3QyTDMC4r
ot7R7Rv9K89cku8ejkLGc1QHuxFQa4PLHyJH7S7ZQQISiHvx7nzNQGQc7zF4FJCl
CsG42kFcNkuzKGSHR98/F5JEakLOciOUOlQ1t2tDTqQs1QeYp3VGXmR0GR3YZfar
qhLd9nbt+CAhAuZWEWiaXgHJxcUTbz9HoVlW45DwHjMdcVrvPZ/ugpqZIozAuGnN
8uO3Yh3egbPMfmcES8sZpiMpGbAxaepD11URXE22IXFnq5SjZ8EkI+vzEXMLYgx2
x/zVXzxDQuj+4OVhlHf2pmG40ldEqUdD4XOAa+Ezn7pKk6jC3NaP3NvuwmgKwg1R
inApvHTs14gACFDxCSwWplS3IuJStFTF+yIB0rzrW0DFuwZ5PP3HmR0eCcAfKnw8
5AiZjqNtTYdnckkE1Fep4hsbUJwtIeSMQ1D8tjnA7JcZg5mF3oE13oo2rTXT15YM
Jpgsfhb/UM7MBvFHBqQNqOyRAjVhTHm0OglE2waBfGH+7dEXx5qlD/kLXPTLOV7H
R2Oyth2nMkB07ujtOjtOigWBOxSwQea/a5r1juBwTDA02S9G4R+rkSsRo1ZKybHs
14drcdJx3ZdFvFMAFf9Im3rp5TI+4B2KeImDmv7amfFlTx+MEEoBJj9pk4Cux4Ms
xIs8B8ISGgEpxR/qQOnVl3TScp6WXwMTtbz6sy9P9fKxiFOQRR+ISga4K1R7Egc/
GZVNYCREgPtS7m8bHf/Bd6H4Z2IBtDM4lNFMMnxj7Qjzz8NgMoAnKUZulQ+sFxIe
ecB8JLuD8iwKHQlavjQsf2vcZrUxqLSRGPOU3AK7C61hHlT9/Clps96aYeXxhwzm
+YPyxguCn6Kyd5GQsh8ayseiqpa6LZ1iHZIH/ZrvkKv+KYUD25cyX1cnqRwFAzze
tRmt6e4zAglA9J7WtMkMhehhEuZHrPitG+klazEZU3p95FLAHiZ734VmKHQkO1Ad
NXzdTlPpYrgVCKNLaBAiF8ofC4ICAiOzrgBKlBJjaBq7PEGwwgDfK1Rmi+WATCuT
yBGMHN0rqEI4x6nB1ooJ415EElb++LvdjDB573gewJzLCwO4Bb77JcfZpKGqBU3q
DlPyDfQNfOj/wndQLCSMLm022vL4evB7NFqkD3mPrBOSGl6ONzv90x2LrC3yF0nh
46ftyyIkal8UHSJpoFYmtwtrBBGu6yUy/lD4sDvs0iSjZHKSFsJCYhxUY10B+pkn
pBy/yKNJvER4IpPTESaikdOGFErnbOhx3pEW04SFkgZmzcEyoibvHDN5ykr1L0xu
8RfrtP8qg3A6M3617+VIpaIZphkMEZ1R0MP76VKA1c5c/YOsgcJD30EmhFLtIlKo
BiTG4NCCffsEJn2EWqF+jUmG8JJy7kvQ30bKk/rXEMV3Pk93XG35Nz1C0THok9pW
qP+44KAzA2ubTGySladC5lrNVSb89cUItL51M4ODz4JlGhF8h2sj997JWG1tstjO
QrMhLdHu5YyRrgIsEIgbrs4YxjI71m5EuivS76e+KGbFz0hWIp152rbeOb9q9JQk
yDoohH81zpPzdLQAJeStIx0BUWEOE9D8j+y+LfE8jAlZ3guH2eAyqe4oNbW/GO0d
mfgJHoDMjHZCDK4xA5/jstYPdHqBcqI7bKegdbGzFTdUzfDTEMY9KWNbtCZxez6o
TeB2w39XRHzaEibSrHv6V4sxleCHR4TK8hF86o9VAXjn45QZtCRy+9qztwa6myEd
EZu9TxrLfJChQ7/QfTO2PNLDm74URPI0EngFnT05TWOaHo8Vfxbe4yShMCJKtQm1
jm7O/F2TUVYZ+gNfwdtY9UZ+JUHFZsNQfvukIFrslPf7DnXt+Jhs1R+WgXLhT4BK
FVGrP1u8QpWatbH22+Mf4yEFd0Y1iMYs22R2tELsAwJWABeUzRs8ILZmd8Oalhw/
BkE0eBhG2oNOC7/FdRlSDGp0UCPJ4XfF03jjGR5pxXNIPGQ9OLEuBIzVAKgpAZ6g
YWvC6+OhP9fEVVWyyLi+7yT6McLBeKMBVeylalkCXAs5H1q3YKWDaAS/YUi0LYBS
4a9tWMmzgASiKp4nMftgtCb6J1SJcCEi7kdN9wwK1WfPC8KZjAK1fTY+a8Ut43ZZ
0V0x/9zm2qK8Kiie7riwaRCc62V4V5OKxfAE5/yf5TBGjjEWtl0wORju8VacKdsm
7j/RI0QZcVmykXZ14i4CQLD+s49N5Rj3ydDOEHZYTqHyXV1SbgEqFvDsOOpk2c/5
lOnj9U2/TaihPgcOLoQR8fzfCrWpGa9/SXDmgLh0iLL/AK+V4hSiyYatBt05fN0C
9sy4Xyoq6CZk8aLrqoCpCLTIXiB6WbRtLwNWqa1OH2EMKglZiREMM8Aofr7j72bg
hrXA7wibjWXbz7nXAwJa3t5Y9q3HdEJw5f9D9aSIEiCNPIZi8hAPeS9Fsu41nuS5
h1vcTiXmRaIySOzs99+uU7Z1kBqbtA9m2m26SmrfvTWNrEC/NMRzLmP6idFrs9nQ
aF7H95zeAvnMwIxsFGPlRo+GK+PZjR0ppgbsOoYN8pgLa3M1rNUReZXKKATHmKT3
hoRIz6SNxhM4cF0k21IQGO7vU/FxdbP4dd+MQg7UkSKS29YarIdXzaE53ijDQdPD
bxc6TIpm/nJMaCwh2cL0MbIVFYEZcJlPGPL2cg3X/VVIyQ1UpdoP+I1D6yvjytqf
pDcc3F+2ns/tJCpg9yagdEoqfmuP3ffhbXPInGWimKSJAo/blYrgQTrq2NjIySBn
hO4ctCUYGxnMDR0qsXGY78qKLrT8du0mEAc3BJv2vMcuvRvPIRo2xPm5QYPzFqHv
2T/1NjmmHMzTBRvkuSzTUVFmdmqfpfBkOGPfFReaKJtSAAzhxQ+V6dPL9sy/0IS3
g4tHzfnwjZ8uxofP3ytiSI5PZMO9QRBo1J4ngS4CtQcGGBJH6SGO0mXcymBTOXEV
LdJVPPK0FkOsW51rDQyAEdSMNms8exS8uuQxueEjhmbGkhizH8lGp3lbTFNM6xDc
FeIHCrc2nYzSkc5qamsiT2yjiV0LLhw5U0p/dvwhVM+frWDOStr5y8LHikb8XcwP
BSJa5vPKK7u0kVRxgFTkwmhq7+nI+50Bksl9gV/pYD9GG7cPHCssgHRWXHD4loQi
2zRP1oLDtZwQiVmPWlF3g5QhXRaEyEOGioK/PaTdRo4xGBph5AdE5nFxXMOjUCx4
gXL+W59ITCoyVmjw9E81aENpdxSd0k7et/PEGrLEMDz6noIrlAPMd5GzWARmFD04
FBvZ9pCjEu9jPR/6bLSzBhD6a50ZKNs4kZOEHCYNrUCpiRmQ4h73mPEkqA+FXb4t
IU4aRIxiT5iNMLTKbkN2P6bOf6usVNcU+jA9DZM9XqX6365R8Y86kgIZ/IPTnH6O
n8WBmhEj1nyVKj8mcKclOBot2sj5RhuOxTVlyR5b+NDeDKLiynZ0IHILRkJbiHck
5zsKljwDDAcJ0I+PAXHtlP2+yMAzCibsq4m1+MJbtEBHBAIjBYsGP3rDqemaiZUy
gGTPNA/KmQbqQNgY0he3z8/XjYaN1adJnInMZ1niyFbiBQoV23ezABbs7nmH3sKA
9x537H6j2i0VtVTR63aWvx9c84lNxblciZgyxbpbJJR8sqjqdK1aymEArF6GjrkT
fsHQ3OaQ5hzaOIJvWfnkJjdo5mcYzcAElCKmv00+Itu/dnBOsmuRAMSSBJWDziH2
IXM8nP4QfxddZRTB3sinNeIZId0rKa8Px4Q9NnOPsGyBqYDDv7XvJXFl19embGk+
+1i+Y83BbEw68NaH7kH/HB6jFNoyxcvc2LY/9VG8qWGRwhO1w5qh3AU3jV2UMtKU
o906ODowtoA6B8aPXInV/k3kWHkWCXw1u0vRqwwNwmsc9bCPVV1QNXqNKRymFxeO
03+PjNkUQjfO69/mf2G9WQqa4KgnZqJiVEC5Y7fFf/5FZ+iyD+COK+3Rvqc04D3G
EeFfmmyDr5S9ej3+FiySAVlwL1AZLV0QKoGiiqCtxZX7dL344BTPyKhTxI4D1TF3
Fp/Mb8aHRtbAV1C/ZFssf96Qn2vWLcAz+JwwQuVUtVzHEclQpDvxdyBNMyCrRGDD
c4taw8V6TfHoOCLzzmv37Wp7/iPpnVNGdULJGf4HVgLScTS9VFJh+eE3TxJ2ZBML
KTiaVU7fpmXOxlekj7awIxxDtFTsf2n9WChTzM3fL2bq5fRtgUoQmIr8Lzd1OH9W
ylWY7avImVIBS4MK2yvD6N1ufBnuaXb1iajyPpQxRckQzkBr147L7KEUlJO+rDfb
PDOVbrn905qdZggQjs1vWG6aPodZ6mI/pRfdSkp+Q9y0/2W+AavVkb59Y1+XIuIt
Gy4vhHL67fidWCWjrZidS7mSPTA6EDMh/+/DvT7yXOLVef4IDWDXHMKx37OlDbkx
i4S6EHigrRIujUBtyxqOUhtiiLjCG7JT8jOkYOzvcX4cxOrnBnLSgTwYyMRFcIOG
5Jcfzs1Y/yNwLF2Mt8sxflLheg6II617+P6nRPWwfi5i70ELgc1oe+P0Q+4so4rE
j1RdHV++ExAUmB+GJSMTKh4iCw8sMrj4bfu6vY4tylrkIbu5rgqQUh01pd0Vn23e
VX2xCweOgcYXU1wVrRKbsM/DfpryYbO4uIv+Qv/Il0K3Khn8UQghHRwJF+tQKsm4
ngsd9ydojFuSaLaqpQiFVhIjIxHQoQ0qNiG4oSSjqGbXA+90wkcaRDsLY4LPKwE3
P2Avms+UfRJe8hJLkbgQ8fqL6i56F3/6iuHVdAYo74tsoMlBFEeRYVnldd1jTZ/k
9laa7MasxgT0+YipzVwEBDY/PvEMLdgm+FBtJ+rlGT+gbukAZa7CCzIiCVDD0mGr
rZcOWW98Dm/EANjXclF92wWdXVk6Pt0wNJsuvX2NiyJzDKGk6hUiuey4BYLpTUd2
qmw5bMZP9Uihc+lXRD7vizqxSRfUcQzXfkxnFGJ1JINelI4Ql5jC0v/A1VdRuPdd
88fISn1FFO2HCG7UoMZ/lN5HBK5/9VD6JURCBGOOFeLwulWUVQlik3O8G3qi7jur
NvQmknWRu7zESq+P+ESOEbZ8WtR7EpZIx1oqshHoFSS021rdGqoRK/n2aODuttSI
5rEHO2viGnDb9X0RzY1Jjbs04DvOPOuzKpi4th8PCwZ+MR+g5Js5Jytx/pgl5lZH
QIus5QnjRfJ6x/rxDtBOkN8Pom1qtAWSsLDUwLlHRs0vqtvaLByvdQjqVBAAq1QL
F4Dt/LKIQgwUErU2Pzr23gCh+iRbIF6Xj9EYZSdAyYUkMEER0t7wTkYz0CcRaxGy
YCXBX9sY3R+kvoWDaFZnOo276QTvCZuckaMAWEAg6ageqNuLhGTQpw+t1ZdBf6fU
xKRbnLMAvcUkYUxwb5OS/i2WFQWCh39SZzBwycQWz+yp/AuHe/ojXlMctmIr6QSC
py+AsJNebT/Gk7iXDZWEirvM1JV4sQNfNNXk66O5Ijzehb9kc+sPeyU05qwzgNzz
fOKmzvOh6IfDZmXCIaJOWV+lnsUxkdIWFhCPSzWOjhVVyzSm7sglYO19R8WJ3yv2
sHED7b02Htmuo4g2wEA/Jz8NGV4r14CR3e3/D3C2o9NuSHkO8VUdRHfIkO/YXgBC
I9eVKqtYEAmvHHdS4bw+THBVZ/cBoAd/1bY86iYlpsEtfdEGbPtgRL3qEWW3U9a1
E+uXu43uUTL4TfC8FIOhG5pAPmsH9UDZ/cdP2vAn1dS+ykVQViIGacDidmv44BgI
EL+GhIYnNqA0/P7a03t00ReZMsRG7+k1U+ezU3hfrmeJZT1Dw7P1IyFVrCU5mA1t
fYqXNKyP17vZNoBuOfEYxwkKAQDLyic8OvVT0fyi82U+BHCib9+7aCz7MbyF3Fxc
S/1ZxjjY5ub4cVny0KUQjswnDcZodYGl4tXPPYAbx1+2PfaizIS6H4abUjnAf7l4
1AerQ9/xvKAqye7NVoCTKY3u1wHCwFfde0J2hRuQp9/UeA3WyZZcfOGTqdrWdahZ
P3oIHeivo+kMurqlPJCESKyKHMCqsYV1CrFHw0il/Ovr3Lt1cFz2BoRVMAbTicme
xYXKsm0XKLbemItFzbqc3V5MkTaKl7uMVJLP2m82AqtcF7F3CBr6TQQUS29hkTvR
ou1MVIZrcymAi+2qq/rhS8mCiWU7CLVaNEeWsiVvT9TSucvAsIbmZW/3qsi4aoHx
KYS/uF+3YtKpM0wt6qmj6XkmjymYokB9BIIOGm2seRXcwRbtcNcqXGxI2VLh+CE8
r01eqD+XdHMsI5IuMmGGS7ayzFHstCJJTcUfExQltv09EQhJbSrhV6P30kWcHq7i
bhjWKDtsv8XCD+LYjh6XDUiqaq8WhNZnnm2xwqLxpy4V2IHVLuA33ZWD78eOfBv9
F5adW7Ahz00izrH/nLxiEjPfXHvr/WobK45e7/MkphsU5slvV9EQ+hN6OLMtCp35
1m5Sh8Jt9iOmeR0/XmFrRU7Oeg3TrjBfJCtgNa6bkENYlgSwhxcmfWWZgdPkv3Xv
d2JbsSSWPX4WrKUV4a3gopEcgh+LVRdiWFZJUw5c8XmrGbn72NmdBF4ngjugWCLV
tngVmZkpwcjoZxe1l6opxg7Sf6RfngTTvWlqrxT/ia68WpmtdA4hWc/AyUslMDcJ
aYVBVTx/rIMB9xqdEc2dbb0dOrkOs7MU66AZEtO6HX+rOE8PDmC+obHL5CSTVuEu
QoouHhddGCS8j45/lGP40a/v91WqCJAZI0RCHy1e5BF9B7KS+JvBlsbEQCRRGUSj
1uozqMXoIUTcGFttdRbih4GssEbUEGZbGxUSLzsLJvp7MNaOxebMjEEX5zmKKNEY
hgOQ5yJ1EsD9VmW68J8BvlmHnPiKLyE3by6mN85uhPCifvbWOsAgaedaUE1mtj3X
zA3ox9VU2BZBK34DFRbUXjshv7xpH4Lt2J6ekryA9LRxrz8YjqZXiLKLtnWdfSxV
HNAB5OJ9cIK13g7SijQlF/4P/NCyvJU9+lXobtDRA2FN4X7pvmg5C3CSSjE+7W3Z
NoBvjOaKQiu/Co5xuYJYJbEcwRxNijlh27scCtOeP3l/k8jfG83lBR+pRbrvBwG2
YkjAKKji0G5lcR7/6sMuQYiz+6GFw0Px7q2w38N6JfKbODL0ex+RAsfaf821gDdS
Y5K1xxt5rp9XTTnBsFnlQMsBFM/sdFbwa1FUqICSwNDPhH2Y89MNrgZ8/uaqVLsn
ASFOPa1msrbz2Ea/rOkN51pze5jj1Wr804Ajtp1Y6UrjjP2RiNe+nd+dtp4mRiql
/6OSJFqe/XCPMv7one7T4sq0oYFbEcMK4OHKaHoz4eA93BxCJIqHD3Uf+RjBsbOE
RY1kHZ4PkpmMVGA7TYnQ1g1ufNajy3els04V7kTqHlZs0pQ4Pm15WzXc4wBy+xLy
ElYQcFBJt/Uy33xClui4GZ/cYKeYVUxGah/xz9QKnN+UuxNoP6Bgksok7SJVPbOJ
4uNjb0kk/zcw0W6JbASASEsWSXhsJwjIM5bqNbwiH0AZDY5vpXTnYGb6th78FaTh
R67kQvSfr62mzxUChxcU0JyAJjkRlKwgZPBXlXPlhjmUWM+zp0TCakq293Vqcl/X
sHvPYJnP7URDmb9J9hq7HalzE18oF1IF6sWYHIIqIbiMtiJFoyIzEH9N1u6kOEGx
OPemXx0DpG8QfmyPD0pgUEefMz3ySfz5LQM9Xqs/CCNXMH7lvn6HoLxqpDumHDD+
+GEXwe0gFFMHAk7XmWW8jYDfLUTWyFn53RmtwYDpySWtocXA2kPNITof16cA4C4K
1y8hxdSyoyIGGC+4CbLdXqZ0FA4YGqlxGMCnIik5EZYJKo4RLOtKO5EDYlhG+0xI
ux0wWCxaaGz2iogxmqPa1rGdnYDDAYV+NHLkflNe7X8HLlt65dfzhYRpnRbvbTkg
NpUuy4mjCZ0IaOXPA6Uq3dMk3QEOadQDivwQ3Zm+yb9K0hp8U1c8WoutY4s5r/qD
fuh5LcBvfIQNA9r67QbS0n2MEEeQ3/g2WZfb9XblEEUNUlCg0cS6ItBkosNrwJJq
SQ4I5A+yu5m+7YqShGB0MB8Iq9Nj9P/E1Bu5LVhvnruoyatRmozj2QTNw0U39cGd
n64GdkOBK/VGSpWjPywppmAGNxiGgpyEtJhFq/6jSuhHgh/AXESN12JIiyDmKFu9
GRpKiAN2peCsqKeWJte5tk0XpGBOGYqAvv/SDid7sMVAEAC66jbma3F5elg1+jiK
QA95bCBxoTPy2hZhGXvcgVRrnqNFURgNhraJ2dCiMxnuhk6YuD7/lt/D8wWP4VlZ
3W6oyGC1ZEjTxYktlwOnrnSRVsH71sbPf/FIAGNVdf8s3FOJdwk6rRRKDJRCoiPt
CMqeXfrDvCAmktchhoA+JzkIhI5SmK4X2xpZArjYNmf1T6P31Ma7o2cUJ9bF/GwB
MjnY85k3gt6jStQKAFmkO1Gz29RWX/AcOKBnVLcfMv18Dh5PT4bpjXPuOfg72mHR
lkTHzZFMAGf5hesSvgjryA2FckYXRhPWKVQreygge1ouatyl9Eg6V+BkT6JIyuRJ
6w4elIjcZK8PbGIWrkPPFeovFeC5kCTcxZHfYV3pvmCIe/wI6ILyqlS/jrY+GdU+
20876jx/nDqLJKBiMs40JMf1X9wctqKyGfxp7f0WSm5U7IzC0fLtM6nAtA9Zagi2
vF+jhutbHL+H77SohEh5HG9iJVqQfEuWLeMZ4Spfb29rgU8UbrZALBocMiTqDGpx
GUN/5IIuf5Hxcpc17kvYo1Px/FZPvIU/ajq9k6UfngBCj3viXXgGeqiVXkusbzvT
1adt1Pl+xeG8SGy2n9JqdxH8sehjLm7Hiel02K5OSyzZYXGrLxR7bTORORtsfpPu
CP6Er2KCWyBQFHFNgFvjjPLWwNFAcuIKuRnNbEzKeF54cDV8KAbznMOqGlaIAkxP
hV49k4VkRM7bLyvAReWEujtLJbzXKszO++9In2sKUnrO2k99y1uGygY+Jc6ANtu0
C+masJx2CJkGOzs9dTfjYK/IDiMkscO1QoGBj33YFZW/wVy4Sd5cmqz7O5GPOhwS
0OBSAq63zN0WpKWoC3VQWzN4euEh6PALoxAjqlrrfWsq4alPXn4FTT5WpHZhOGwo
guR2nGNNnw4SzLkcubtqXnp6o3lzqMxyjfgc5I0CUTbxm5VwUl8efSF3q3wgrmZm
Z5tI7ZQFMc9GJ6/mG9htnnBESliaw7lKdmEQHgTRIobuNvB85Kh7d6ghtUtmm+qZ
L/LP7TQETqVpTajAmOLDJdok5OcaJYayqsIE8/9PeZTF9hkAuU6CiuWp5+eZStvX
CezaMCmfJDBtTJAvTzCi7ZIUvkVPhPqbtmlOPMWjEx/QMEnAbP19Hbf1h15jKuyO
flDw2T48dXfdR1fy1mT1kGRm9j60MnmIMP++f6RC3JCJHj/rMNSczo3T9b6b1qQ0
nJaKaVmTfe4mOKMl8aIqBPjzT9F6HpQTj2LafXwzsbLJnypPRTgAjA4h/9VB/lFz
uf9YJD02zFCvOOgLfs7IqvK2p2uXwDiMQPjbYah1jGuWn36sesuCvoKpCwh2+vxe
hQm73Em9KjXHB3kCbfX9MtpSwlzPPx8hshgf9ZExbHdUBffkOYwn6xQZr7fvUmDF
bs0E41/jyV0Bp2I0OVT1WevOkmjvWoQQCgcLKYK8jRNMOzTQevnlk7WTo7t/VC+1
qGYFvvBuP3wRUYdEQNmcBEHCQLkXHBIjTZxpRaQe1ll/qj1KppxJnW6LmlOCuGXf
WUmfAwBGqlZA2y951X/umj6HOwOoRGemC6F0/nY6lkmB6pZG/vS90PcrsX96KENU
SCsCcoN8QDmxT+3OsXxnLGXsXUNh0wIOKXfN8tTZl5EqXojqYA6ff3G/GBldt+G8
7BJaQKpZePPdQCzXFU+xktmy+WNFz+DBnKclArQDU+qe7ZpsmLFfkGlkw8sURnLe
qUIbp9SebMgH1faetu8qNBwSFEBRU6lCNP1flMBqVzgdntjR91C7jgnb76mJKunQ
LECSs5p0DAE0FlkYxlHi4wPnUO7VbNsH4DMJJ0K+KDUue1jqf4EnBzIP2V98uLwb
uwzyspivrP3q6p/2xISEvhK03bkKY7kPSFNCnstjeV+z6loavJwiqJwSzBxJz5eC
zvIlTF/qlXgFt57Vi4TTpCJ0EzDcqHtafHxVhajuiE/WAg2QSAIbVZurMnLUel9I
N2k4VSCaX0sAwl9tt+ywo62dmIkjv26bmaekfmujw9Il/Z7Rh/RWbV+NTF84VGPd
Zq52BLDSaHVCFvao23YkxJFzn/aFEszdIYdsCMm9vs8W3fvunb14Z2wEZjXXdWdh
NarRRQQVsmcH7S8mCMHk16tJgek1o7OOX+CsISI+9aVHPDdtEjS1SAIoKE0raWXw
HCt4a4NrS/qi4IeUROwkIUg3OtuXQwFbew0jemui8pdCHnubyTC1HuSz7v3eQbSn
pIOjKA+/SXjBQcdV4Kqq+mnMpaixtVLoxOEW7J68Yi5+tc5z50l1qzU8uXSQ+1hH
/fHRQIrEmFc7DCzinV8W+ufiU6kBeMnmwxpRFwUd+Nax3Hj4KP5dolLE3NabwSBr
DtZPg1MsyYzeEWTxz1aS8iFnKtJjG30G5yUb+ybSENisxHUGazSAuZyOgb2lv24y
T6pBRGZkLwcSH5S13iC4kcBnfgxOrFL3H927BdZiQlovVqfgTgbeghA90NT2R0Nr
3T46artKcMWMgHbiHoFmQu8HBMFTAUkSA98LzHmQjX8Y9yxrnKNajfKDVQYoyf3L
xGK0SmGQRcSV1VvPwZw6YZaF+W6knszjTs+bjBgXvU6T3UctDDA/gxPcsu8Ugr2m
vJ9He4CFn5uB3RHoBN17kIK3sGDyao3lD0w9FwdFcB7V/xcc51XqyxNzKncxc1uF
VnYUtUdNBi8OCZTy1PfDbTb1Tey67P6gYTFJhPUnsZMM/eaXmmZZoq0PAAGK49EU
ljp/OdcHno40CwazBbBlPwraIP7R4I6bD+AoFkn3ELMmmHPwA8OKUQYBNmG9e3o0
C2IkSklKsENNcgz53mPBjA==
`pragma protect end_protected
