��/  6����p�>ʓ�Nr�]�ƎL�(��#��տ���,Q@�V���!�`&0Z����r�	M*������ �;�ǣ�ga���(�)�$=����������|4D8q�h]KN�v71[��]C�-�P��)ݞ�hz�	0W��9!&����^S�b������Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9�㑩=�<y7�n��;s�ˮ�9�>|r] ��Y/�M�q��%���\! ڪ���qd!�]�㾬r��Vo�F9\zш���-+��p[}���B
��r�����#�T�~V�A�|����*���}z�)�Ԫ{�-�0�/)$�2v}��ˊ��!'�2.�&�I��CI��ŝ�D5�H�c+�L
��M���	S�7p���&�%�=7���>vz�˃���ܗ�W�UH��"�Ri����&gcʶj�cXH!5�Rpmr���[�0Wm�Mwcz�sO���}�`i�LZ_��N��@��]R
�i.w��<�,H�<s���� ��7r�cI6��7���e�&�%����%`�顩�O:P�*7���\�xx��h��M��~]Ҁ�)�r�n���I�ǀ��b�7zU�v�@���_��Ff���Z��f)~� ��pyC����\�aQ�9�;;�[�4���8"������q�Es�c��FDy�֛���?�Q��U�<���Ҏ���x���,ګ�:&qFP����(�qI�_��. ܻG��T���d�W¶1<6��88�Y,�)4����Eb&fd�f0W:ƙp٬���|��%�#/X�s^�����cz�������H3���C�BP������wxW%�s�G���4��mg�����
�Z���V���]rN���d{?�	�9���$�[Jئ5�q�a�8�W
��Cv�\yJu'�H_���C�X�l���3"�ޅ�ߨ�=�R/Zu�,&���Y�Ў��)��Q��׷E�����i�li�|��]{>��W�u����u-Y�f�yg�Lɓ/���X"���e!&˓