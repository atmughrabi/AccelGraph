// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rb4KKZEJ2sDy0dXuNJ+/Myg7wE0dczoRbkv+LQAlAiX+hslPjzRhGYIQWF//iTCO
5uUiApA/u+39AYIqZd+sinxVmNxl3ja3/wwm7PlGOpzpMJs+b+gG6PnFmuAmTohl
ryfftV2Y8CvjIqY3FPnLgk5ba8lfJDYH1a6lmTPZfuo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4992)
Uh+GqUUlBGsMoDxt4UXDAEnJ78D0BjwQKXC4tc5V6+urA4uoeQ70MNU04TpiBR1/
TyiI8aRQWFYullfG0iiZ+x1er++4Sm1GpoxHqQQSk4b2lCHqUuXlxfkdweLf+wnY
X9sFKNl4e8ie1ZDMmCp8t99joz5JF13QMC9wawADNBcS2/GRhzXYBCOf6xrBRQ7G
uzX2lAsEmKgzHsBfpRDxiE6ugGcP+BkqftuM/4NWu7YDsU9nMDBh2z4BWj/nGOMQ
oUCy457HYnNLvJtnGSxfyKYo0gB9ltAGI/IZ1VXzDG6Y3Luya/sbP0mWbwpG7usb
WgCLmiU/qP3ZOvjhBZpFNlTinb4fUnX3JSRJF6yWYHzcil2ZrwIs+0xxD0ttPRNZ
HQjIpiatnK4KgkcEIICPjnnwFTIV5Y1qzIIVCR10nGFpcYsrjXJzJ4UXEU60eIBO
1OT9OOMqVOumuWXtXsVscPMj0wTdqGbqfZcRM5uEraf84HRSNdwRw4IIuS1Bnhvl
lwwspeoXJbbDuDxM2Rq/BTJcNAsBL6CCyaTstLAUkP4NaFyQs5b9jB7eHxnAgl2g
utnxmoXiicJiTobUIPeK/o52C4Hv5Z4ipAjt1LfhZFo5iocyDa2fXKuEzlRWUzPc
fwPxwkDtcu4jAbjioqxTdnffXuKzwIz3bxmTR9WQO3ftZ5hi55rdV6cdSDAdnCIw
RgY7QO+J+/VmTumDRJH9uQzgooMj1pde5JSM/z3aGVHX+G+W2ziK5GbkNtHmin6/
fOETOrST+FQ7F+psN9uqerLgSXmnNguxoeVApIjKpK3z0JARRv3RbtdKeE11HYsB
/Hx/WOrwoJSJIvDyA1mOqEVLctx81ruGSKzR10bTen6QaHt6dzklqwcxpmuVcoVj
64O5Avj5WD66jzJfcXiNdBOjX2hntRFgZLa75w5TslTP+pG7baWrSPfivvWzslYF
AQySNc4pYUsXt/vkSoJLlfssAfgqm9zOj3O/0jOVmRCphfr+2GsMWDYftvDncoN7
Qf8HgJ4DQeQT1R11NWvck04B8fWCDPJexoBlgHRFdLa97xUQE3pIQPODteFyzTfd
WZCVngkCSb4giSwCne0n/4b8rGgnh3QGuknI7TyeJhBCJ3teS4Ee9iFG0nOQ1omO
dztEHmut68PpzpSGoyi8VaCbqLBtkogRDvqUPDJ9tCT8ECS4DUretNIXyFm7ARfq
rUm5cts8lErJ4O2TG2SBtrjKHPn2oHxV4KlhKr2rr/+/3rHurCTilmalYDOiSrZ3
nNrJGulwA2YCIJ6WUVb1oq5xcEb6g/me/Oc5kewq24IwP8AFBgvUk8wm4XX0QCyk
xV1qb6WEAvAY6LRnD+T9pldELCI71IbydQ37QD2P7lMok9ReDeT5hQQLMNqDzYJ2
qzEsdJ+dB+lYW2iKxWCSbsO/mr8yRvjam5mwSaI1xUaarcJAZXBgJchxyMNnNGJc
njbThYEghI34tDKSq79g4BqbJIgzgZog2ZDFH/tlvsgkrlW1FeslVe8+a0nQrXBZ
QbWGxFUuUH89/fhA+HaERH7LfI13nBTIJb8bfkdd70glBdkh2oIxCteepiRay2Uf
q1KK5fbJ1gPF9ILlU8yH0iTOItg/WumyuQM1E1gVWO7MtvTXkfpxTcRj906254LT
Rld40xVgO53f6bQxpolQdX9uVFwJtWz2fB5F/PudjzXPPEyU9x8W6OgNLR6u33aK
fltFZwYhiI3CbH/xGuEkE2sUx37WmJUNtz2czYkOJwVJWVtb3anKWYCwKoe3lJQm
wfjZOBDGnV+1J4q6L+D1kL8N67ZfJCsvpN9Ir+AdxDeZxYrFTMMAU/35aaEqhB3A
XK5am1NVLFOLMDQjEod2NmcI7WcTQave4ak6AJ3hlPpS9nc4i1H92vc/JVITpiX2
JROOGUh6Um9RNOqJUGLzfPJjANafsNPovASXqBdBw8BTmblXmaT62I2LnMXEnPz3
/kAfQWgcqiE28ALXGXCzwHXx4SX3k4bbPvr0AYMDL+yY0RJ3tNOvX6aWF6fBlhwf
2wN+yIN0fnupgxa4RFdpjVdNmOtG0H987OENE4ArwxbnQAFuHglOJyRxovTQPG5Q
JiliA+6wvSO86lXUUgLxx5ERfiuBDInIYwa3NNDmczg4fH9STyhgquUHxAaTWo22
dL45TKytwB67NoRbaICyLkw6wqqhz695M2KaTdKrFu7f/ytuoyYDsRlKbEUoV5Py
aE+CzlXkNnvJuL+yKBtxkF2n8PM2tkzBSUdxZH8UO7OD2GNW2vYbu6s2Aw2QIv/m
85uZJSX6dgsFmMtLLS0Wn9Y4ChLnU3rlxraInZhE1o/ZPo8pXyElcuCyfebzWuGr
Qzrph7vmkt/jaigKOje36UnMAtuQTrDBl+oQO+24n66WstGaNxq8PRkGuuH46M2r
qgPjK/TiS/DZ8TCS5ZS7Pukw6XBY/swzezY5i37NZOa5twIDc9tz9MflXdTlIc2v
qcyAoi/3F2FB1rgwLkZ3z69R5OmxvwD99GPJEP9Nvn1p7a5XO0C7WTENT1DBj3Lu
g1M4jvxdVO2j2AHjAieuY4PwrXxdH2Lf4NrwVZH+x6OmF3O3BvoqmVENgSqcgj4c
yEwE1ENSqXqk/lm+DwdOyXoowItH+C1vn2paL8Umd0HsCBZXN5XJ2AJxTVdw5oFQ
pSd3b6uLyozBO6re2SPdC922xpa83yKXXkBOF6rbeCSB3niCBvdoAoMRbwpTUF2Z
NgUUgg41WfIfYjCo/UwO3UmIelrClx38Ghf5AQpvbbkdAXWOGKwkm/wiVtLVx6uc
ET+xXzday275XHyLdeozkr6aXPSyvbpQEcqIIKY8tYHytbQxVZJcDCEdpkQCF4JH
vVwlYqOE7hgRQbX1ef64oT6R6/8mhdhK13ofkAfLQU4gNtMFlesjvwgGgiHtGsSf
4mFugNH//Cz5lX2cxF3u60ev0F18Kd+12rLKFr0Uum6NA8TQHWZCLysip6hz/BBo
GqXs9Wh60In76hhWmMFxLm9lf657TIKNKFEgmBwxlvSBMKb5RFHWCFf+n54TYlIy
qwiqipO9XRRdMKG8itMaqjPVzNr6ecxvrpVUbSJDXn/mwB/cdlyHGn51VyT+IUqc
c3sB5ZUeYg1Wluu3CWQYh23G4qrTl+wxwLyR41BHahLVFe+sfb4HkcRG1dMP7iAc
e5xaAvi26zB0YLfLSEjowhnrirwc9ETESttBvznPNymUjDrCGlAWW9jc+aOJ5vxB
6aVm5hm1WvlnWpEf0PlbIGHkpnnZ3Qz2uzOTkVV8DXLgxPPACCyX4b6ArNEXDMl1
rKSZPtcTaEA0H0Yv453Fxha7rs5Jg9IJSoWUL/G9Iv8jl3k0tCpjXt8XG+FbQ3Q/
1TYH1y39uMGtbdWucbO390tVV9OdrvH00pV6I83sVW1qGl2lX9edyB6mOF5GoRLD
ls6hWPSGiremx9likEQ1cvuYP/rsapAqkN2NOfQB5eE1rNQRS1cZALa3P30oBlBW
7p4VQo0OgL98oekNuIRaRcr3hSXzimIi527fCJrie8+O3YfO/NlVasea1zogYr6Z
r3JWv9sllMStZBSx4OaNiCMMkGYRCMFysgBy5qUGbqTlNH+CWHsOQRTffb3wLGK3
WjMKYZjC1WAwmHpeqdNi+BIDdThaa1VFoUxxzFVbesBO85jaB2Q951T/8izWwSVp
QWcL08IiXLm1VWz+5vgHzdJEMlMIAc65obKQM/m0sBDbDAcnQrA1HF+uHtxWaByN
baIaQ39LEDeQag5LDqMRjvdc6qe0G6mVgLCNx+QNSqXzVLQvla37CLAuY4r542gg
1AyjnmRIcdrg0LZqtwvxtCLfFJhDjc6Krg3fUMsQzwr171KNvT5cpg0HVEfFkAXa
IuwY2S5LwrFeUlafOqA/BjUceAvMvvL+1J0VSqXrRmFChpIcQ8eleohDcb51i+Wz
YHdTtEvcQe8cG0R3DUFnFbpK+vcKSPD5L7MT7bC/M2cfG3rRL+XrZNBQVx3/m8Zr
BOv5CpM5P+kedstWp/sV3EiJsMntpNmRoOXPtkuqVnDff5TCCfIhCp4PmSaZwwP0
Ex5dN83QXtt+qPaOpFQt2HIjwnYJPFfmhxhzIIMmR09UnmH0NPDAsxqrywpS8Gef
6iMCZ0bIKQEH+JlaBOyO4j8hRpc2A141lzuYIpBpeGo7SpzzvUhPtXdP0eXzo0OR
zk1pJHkpEgm5zYU4A5yqxfACnRF8JdmyeTdgwu5reRifr6bXVeq7TioOmoqItrxQ
FsZyRdqrH5ELlw2edwqYtyLxcGeKM5nPcPM0447g2OYMTT6/6XPgHwqVdUE2H+9p
rk7jvdUaJ7y30Pbgm3bCPTKe02pBeZp9hyOoMlUh2nKoCUygnyv1KNbgPydu8A6i
xwOeQMEwHSdemDbhibcGFks+27o7dascRS/2J0uEfAbGuQy7FJm8ELUBiv/Afwc8
CdjfwG7E71A/e8roqS3djOs4xPpc2eeEXY1O2xCnCp5uQsNNino3YHtpMNIAXf6n
XkGk+0lkELtok3Via3w4i429F5tIdD1Y/0ltvBva+KGjawv3eo0DY6cQHMFK3cHx
arTbmF1pISQdGECjo2Nm4WDW9aPfSkv9zpzAu3Qi1c1rdE4JZUMk6KTEryhrWb7u
K4d1vgEDsY8A7ZQuga0Ajr0QgLfH1LsObIA7amFNIquAr1d3AXWGdCDCZDcnNUVd
5B/AmfaOb6IskDRRUARqAPvqncWhG0JOSrRIlhcSySSkzMe6FjnsiiKbLP5pRY7v
1UgcMbQBMs07GAZmj7EROLYGzkUZpVkzBNMcuXQ1POhlZ/uHfDtd+M064I71mvR4
4UObpTqEC1a379de4DhBIDROaipzpVc1dCWom/cf8S/ujDJOgu/gHf/0HOZ7kk1J
niwYLbwt+bikxraBkuoAnBZq4i2G2DDqAf5yJIf4PjyPFN1XiZ18tLvdRXawM+N0
RNmVYPXV8fQ802v5euWbF+QQDGkcBVHVl8izwxz4EtPrvs9U7MjN1n3c0c7H5BWF
t7VUmkiuhJyLC3OYxf1NWL2BnuO+97sCxZcATN2Mjs/+SJ1yu1CznRqKVzmchwFy
07aGVcxUqul7o/M/jllbbQGhHcHSJUF59yMBGs9qmZY8vqeuqyut7avPtD/TaEWZ
DHR3onNjIYcKITe7xWAy93Dwbv92TOpZtaAwDdxw5TC5SmUD9hnj4lskwvjaIUC9
hx+nry0RxprWtsgio8JHluPMPr5POXotQ7522S+EBKSRy9NVDV5vRbaYoGF+oY3Q
yDQPtU8dsotXXM86aqECJbNeSXhgV4ww+RwmG6sdv/dchyGGnA1/hg665yktIebX
HXN/iBHOHRBa+Lde7J39NpNkTsok20bsAbse0WhhU862vHQKxvS6Fg6GxTKJzNhF
aFlql33Cw7o57RiOdyZlr3eXFsD9HQ5gMlffKDO4t+SjEElbnPBsGv/NJEvN/vW5
WHQF4DRmC3FO3R0TFr61SU8DDZ/kCZ+8o/W2NlhrdQ4GZ7uVu/AEScfwIvqfN1u8
9IKYyoSig50/t0JrIEJc7SKFL+1xrXRr+uvO+aknAC8hHy4uCsO7jALomnfXx5pc
vc4zWdYwPy7w6CmdhIK3Dq4DieiBs7r4dVb29wJ2oLyY6yy7kUmsb3C4rzmO00lZ
rKM6QTdeZ5ZBZ3ehemJJJl1sAgWlj7n/m/k/Lnc0qHq9n4RLjKJKi7jP31Jix7vW
UtLGQ6qyin3eJdbX6JgkudJmJb5M8aAdPkJhtu/PnOSLCrAU86bX+vonztMROo5p
vkrr6HKkNj0X0+ZdcLt+AjKpZOlWm5t4k+oWNXZE49k+2pOsIMJkRO7YjN18Yv/A
xdLgtSabgxcOM/1lmgrnrbnBi+713jJnDUJSJ5zBegiTZdlwZFvlxbaBaZvqcr+n
7RJ4Fh14zzClZaoHms7/MIP3a+mYRTGue/LM7xfcDN/etXFkrVjwjSEDKxHmgrMc
tlXikN+VC2id6orMIos5EOs7W7yWL+OiAmMvd/HgEhPZBJIbdSBmESNjT+1imo8P
scrdtAp3bhLrdwSMfU4RLxlNkQ1OW78V94ajb7ponJJYXSpzYoJZ3XsOPVMsuH32
bpz6KkaYldZ0WK2q3mrV2CT0bp8cFU0K/Yc4CBZYIe+Fj1SBfYX7IGBrCPoYomyk
sy2RaP3SMtKlnZRLbLFqRbnQGVcaYzM5zcHTrMgt3m/929QqfMzYRddDSvg5HLys
ma9gU+mtOr/55vibjJ4G+f4xSngscUg8D5rwDHl39B6CAqmdZJs+3A86JkwMLDET
KF1XkzAEiSfP5HBHSYH5Jv7aqtGotVkEHFjdRnxu1BK05kQEkDZILen9Vyr9m4Sn
sF+7kM5Zwwrg8BXA0wMjxEHO0XJq0dp5+0l8Qo0nNZBRhUNgQamLh+z9I1x9nxCa
OCvVIb1Am0CkQe4gsnRuLOdVoq32XlvJvN08gT9su1Q6sso4Lh0igJ4Pr9g5ub9G
y+0ysVNfCvP10hWXjgflgDvoXHiYvGK+WBjMiS4Gj8IIzmtnwFOe7+DjeVEyEQtQ
TqJcsYy3VGXvFDCIxfKIsZ1Ekrb1dnYQ19wWlPAVbTLVs7slcfAcfA+BTMpC/x6B
`pragma protect end_protected
