// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
R/OqbEuCTVyeGinR4t+fe7fENiddVVx/y4JnCVN9xh+B8xCNdlb9sfJAnuFNRyhNowGSxpQ+YQSO
5eD9iRusD58kFRC4pysW/K3HSISGqSQVCL4fv2S1mEtN8rt0mm63VDUwBhzZ40/6N6A9mo20kLNB
j0VorzsW1LasXrMwdSjH63UzjCR/kYw5736MT2Ds+gWmw5SvYoP3tx4siYj2GVef7AErfEAB7y9b
JnnY8HLphI9wmPUnDFFu8BAPSsVoCcd9juSDiqJFuTgr8o3Q4LT7/LdgJfRWyubzmJ4dkVwbMiXt
yNloJtWzbbqLK1pVvCuBBdB/rQn+G+pyk69Png==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 23024)
Fbyoo0MMUW8+BzAzq5ggs8ICAJiGjjwa89Jd/lrl9g9DNShJhkTuXBxpUL64QIQPDLIz3XEBnewq
+zxMma4rbIri6iNnOzZpmsuKmNdsrV82cTqzP0KPkairrGSCnEQbfideHmIHYBfMYgsyKpMCbZrV
YD039qvKWOWmzh19VcN8g4FdYUlxLHgk2PHb+tY6Qdy9By5Qv3JL7G7Vj6lScbTU4yujzFMDgUXS
QtEi2ELjhgkki5DGg0yKgopnbct9c8BLTDqyqqJbvzjFt1Ji8FZhkTwVmKmL+jmmK39/SEJhAsPk
p0WbHnDtgXBmqzzes8+x2GC3o4p2cEWCvEJsSy08UQp5d8thFc78vKXKWnPx66Fng/b4kRMfLufA
JmOqjQC4ALH40ZN5ghXVY/DzMS2PwRFSxtuZAwXk5IZgV7uI1mgF7mhRZhT05T0ARBsfzKKVNqGZ
d2YbCPtaY4MnbiG8O58cSUG+7fcozYNQzicrXuU8QMLmpRC41W3fArobqr4k3TtXiaI53tx0ZMF3
u6bPoZA3OBGxYkIrjv6d0/Jw8oo0g7cMI46JkOoznfNFeE2NsdrSr597qGt3tFRimgAknGJc0RVr
dT0cFTWE9mHBADCCcqR7oMAqMEafBIPz0cDjrTMq9b+rB3uz+AeZlgxCF5DybwIK4MeRRloLa3pB
5YiI86997R1oTlogBxg8zrpf2eR6+4dvcnsls9KWLTWw00iUibv10hMfjM1hK7mCpSf903kPKHcR
RrrpMX9LQybzyEu3yIpSqxPq3qGsLXxAuj3FNensrMAgOgMwiHLfVmvwwLCKRRB9SDFhZDxryarm
yxlxV/+Q1ocEmwglvriQAi0zdJ3AQUW285zlPw1Q/TS4+zj8i2dLFSnWHXARt6GmRy4BLGlSTRXy
Rcjy/q/0r8gAGDxWNjVutoewoemi+/7Ezs+7WnganrE49bpQfj1iNvfuJtF86+K6ip4MX4WA0L0i
PzC78u6FEnC9r/sR6mSBAuGJt+ByPdWAga8xCn4A3lEhnZlJ6I2VGpI/A90JPDubnwvxDo7uBbtP
n7vEccplzQhN1V/9N0SG53/JDVtK90tk7rWg00RI4Y4Oyj0qj7ZgIN1hNaWcKzvZS0JBosAdBNTH
D0FRbHan9ZQkqNVv7QZeULPJgLmDQv10Vs7YvYaw1snDwjzFKrfzhjgp3roCWGoNxS97U0+3opQA
Tnc12iUDdZDynmd+/UkHk36oRJIWI4/t9UKQi9RflaP5kUiD0BLOtmgmgMkuDGglGm7NLNNSFdrF
bfT1VjUZEZ73gpLE/vyPN/oc/HCCSYRBfS6J/noSvKh70mOib13zi5iigxIdAew21BESAKNqBmPt
sQAi3EfdN9cWVUm45qMG3O6LwlYuTi5NkhPPWVqTiKQjXpEh2UoHQUuB/AYHJa9wtdwZclvwh7mp
8IuG1nd+kF8qnwPVkdU0XpRHZAUOyOMRPfpGMW9vuEwPDdieEDmbZCOdgBLq9QD1mCachNZOiq3/
InWQd53gJf1xPDViTcGiJkCSriRDHLyDFEBcTZmYeUl21xM2gBcyPLlLoOnkUppGlJX0r3lCQEAy
kUOW3Z9ojxi92d7r2GGI880HCQRyC3bqejMhl5mTnHNbLgrISY7eHo+YnfQ22lYcC2lwDryy5x9t
5+w+zYLFtEBE/lBmrgL1r93h8Mp8r8zpZAhIz7Ugq1wJ9rB210u4MbCLZaUq0GDSl3fX6BS0Nkjv
s6EVVfn3DL3dtTlI4dFfcHcoTJ58chW/nBKqNaxnJoqRbJI1gds57peIX22LUFGJ6As0MxocTVSQ
7YbIWeAcJbRxS5LxFkxz03/UUl+OSIKUuunBs1Y1C7rqA1NT/08319HLGH74bHTjhMz3Ul/eXhsa
9hZ8waRRXKfb6otf7AOGky8hm07tc6m6JV7xyOGpQSqkk0xLLy34Su+pBdZ50kEG6n9kAHFGe9Tt
iXQW2Dui2U78dC/KotHYRvJMkJOLZT2WjM+QKJ5kkTBMoGkaiBpa3F3F/F8LCR4TSqilFe66E9Wt
GgbgNi1j5aoLA/KbMd8RnDZPABc5vPKi4V84IQeFyRqoXW1senfO89OcMCsY9tPVzgYI0LpSTqTw
wFRebbjN2H2pYfYMe1DsmDoww2aheMbCPNopXQSsLfOLCwUApPhub3k+mMDEH4w1mcMDdC2npYsx
3Y2tbOGo0g+RTPI1RPTPg9j71d+NbypfIZasN8NkwRoNZLGzAxV5D7ThSu2mK7LwkxFaBwBeX+3O
Y9yrqZoTy3+Ah1gtnhLOvyvzLvLGwwjgUBFrWSQC8jxaau3SkS5oBbWYdS/a9ZHV54B17IjE8LEq
qi1uiAwoqRPEKEm/3ibK2UpMdZttW3jydZSUc8xzc+fuyJPNe39STrMmfx5wBuvmWYTOB/LcyDeT
zM0ac4ylD8d75NhrJ7EK17+8vNbaxrA9YHOButZRKc03e9X1E/Ke8vUIZKgVxOFh2mq/NFeMkeCj
bFYw5dtfZApAgWCGsd3IfE4Ol10Gn2qHCJvOdKkUI3sHGoAdtS/YW7CUI1hE1q6WjnDw1JcSZrZQ
pqIq7S9YtzNaRi4Y7KqsgiLUUnR3z/19oBzkv5qAQvKh2q33wTVtKsx7BU5Mhr5nEmOZ7BbCddf1
5GWk+mJSk+55UkCrZiXwnDHb+CSEyDjqg908v5Ax0C+3YoO7NZkEsZ7U4NJMj8jcWCXwEbqygtTr
Ff7cOI8irYTrxUmmbukEVuo3fC/j3ytI0Ij34bAbyO4gpDkMb1rTWWNinSPABej87chquYBWAgpC
A0uBZISGt/zvFEUyJLPkgmFO945/CKj21qV0RROOneHnNtJ4WG8z05vd64e3aJk49qR6F6assV1b
QLHU1cuAi3hKjvUrImep12ZCip4wB7XqrGQ3WzF8yje1t5oFJnFUUUgOSvpInQ9gTT7pCuF27xMB
MeF9E8X3+GVcXicg26OwOcX/XjbCl8zgpfiELWU7hLeDj4WajR6xFOqnPvOWz+Rpv80VoMyiJ4C5
ozaa3Y1W+S3VIiJAgzekfnXXKrCRpk5vEX6+y7jvgiHoph+YYr/+oAnkmiiwiLttYSaiIPpe7MxJ
ob1rZslDxL7/iLXgGZ2wSrTC86zqz51DPyWt9OTxeOcNashqLzH3FPLiQFMcT+WViDazeE2770aB
s/XFpzyxjvFvlhHm/EB799aX3WmkJTQuuQfkqTpNc4ryFUONTEn3whAazgV9KHkbNSva3Bth6HmC
pKqGHBJFCwyshIboAupZHySXT7A6C03lmt/W61vbCIO8CNZ/l6OqUUFoPt/M2r/KoKhVf3xdG7UM
oR1Ij5dBobiOsu0AnPb9jLgjsBE9zGSHLfmFVaoVD3tAS1oL5xByO4kVjKFTY/e+/kBgo3NBF2Qw
cauIys+WJHB1+Odnne1yWPlLhbrM5ULrPsm0Tp6ZD4zhnMFeKPwZDQnTe7eg48HGGf1rbeDsyN33
qE/L0yMPh+Rce5VWYTkoG6woBca+FdUnE4KhRQrtLDREQUTCVUT5LqPRmKQe1fBpNBu8v0uZWmsZ
wr3rSbv+m/OCW8Pla/y2WwMQ7DP6fugy37lTlWMrGlxeJ2rzWIDJPKF0ciyUMVbVROvBQsY0Dj18
h5vegg/0YdFCaClMgsfJ6ESMPq/BemUVlMyl72QOIQdcuvbVORhgqreVI1J5SVZA53tf/x/gsNxU
gSEjRwadUsYyg9MPPgMMqu66wIlFxK4HH+T/GyLofGy8gHr11cdzNsPGXugcZyLgTJSuXPcS+YxZ
VG9DkD7o45aXoEVndNRwuUFzJfJBrIycyfnxYQ8QKzQ+YuqFYUzGyMsRAWmVB5km5nlIPqx3ajzW
Tqn47DIB2DLcjjLg9BWf9SwuBTRl9e+9IevcHkjTzMq04vYINlQZs/UCWZkVu4pSZkThqTdAdwv1
e0UYdD6aPzTs9x5YYBlElfaCnZA/zFetZizDISYiTnewOr+iCrQ1ElhYDDMsszeUmFYl6Dg/hx0n
zBL55qBwJP2j1hgGujHi17hVR7AcJUKoURShwMQUuR++aPnivGS2crTdIUL5gmNpZ5zqNvCRRefS
/K7xdFJ7CgXCbG7ixZKjCNugcz3l9zkbxXy0T/juHZ4QOUGfPz6CjykaYLiESFXAxESsA5stLDAe
GBTbXK5XheW6ro8lzfwKsNdTZMM7A2OuLdSKoPmP6DDmZYuqttKNXUU7Bx+3RaWBtPLKQzlbsbzO
3XKx3/oYy6ivPoY05bFqTHmxsMjgogCSBSszM1+1RKeEgWSYXRffkhZymNwLpKcVWF0/8qiIfTHE
KKeAPGN8dBU760ZGS1kJQSRMnGDFYlpgkXZcZIQHvGJ4Lfm6aMvFxuanmHhXOvH3yolmI/OcTNYG
sbtZ0IqmUvok/XFKhkywewbG7ir2nmd59qKYRdPTQTuZnpvu4LCHERmbvL+rHzFkTu0HDU1O4rnj
T0ceF7KL5ZxVkSkIdW2Ppis9rMY4n6PbMgMm887rWZX4rJiKHRSGi9Y5yTDJR/tT2pvEEEhCM14G
zExMLgAquLL+jua9l+x2ttkUAGTeSr0X+cEgGB0KeSdtPMoHbG/F+N2KkqiiuFp+YOut2INhTZYi
UYoyew6tVzkAbyY32kSLIAgc1FWCqKIw4TabJHU7d00c97uV4zwyKN5pBeVC0kj0oaAqyAKQKj9O
W/wAEjGyOOvxwWZfQF+ahOxfSJMqNZjgumPCI2nE/X3jocO+1GmMlmZgFVAuPmqauoviKWrHt68i
utUuCeKGMzNXopw+1jF1XXBxvCqKOPKGLJvMFzX51WejkDavIkTnNYReo267uh01zZfQXyMJf384
qHBLXt/ZJ27GSJ+eLW45ZZQyff14LBlapRO4YrwBgC9lul5+hZPxeLWGQrAEmLBkrvdpGIt+wesd
SHUoZX+WdYr5YoZlbxF3UXUioH0Sm+M/sVIte7H5YKnJSTH2kVi8/ZbKQkDWJupIyTUY2wAe05NP
O9rTpp+2fJc/gKa+1TnkFeoQXSaXJBWKEzyPOkVRc6yZW3afolsFdMrLX6P8h9cIsr1lhSC/vcIL
8R6Sh1L8XbBpcrubwL4hDzlC6QRfnIcJzcRMZ4/8lRmroIX+2czM1fawGCWZI37+ggcEoYo09DPt
uN/13/LS2zSxsOTStmBfxK6jiqAuX8jS0u3CTgC7ioH9wGan6YZ4wm6eKThFvdRkgagGtdoUxIOa
wrs9WbajLS7T/MVd8Qv7QudblNiQOGfFSl3hdPJBQNAmRi89XQs556QbIMULNjnq7PNOri1a18HI
/w7kWCm4oBQ6GFEzs9ZFWYRovY4Y2C7Wtqf2TPsUD9LPk20tOhE+1oKPCmwpS+6n/Ie8YEjwKX0/
eowPoL+7UTRCOMx+M+jUoXXjqNuwIVkMX5HMQfAn6Y82dyAZitB60z6ff6AZ5JIs1KAFzrOeqcKd
f2nguzJykobqQb0nWlPCYfsOSp+ktf62FGhvds6bdaU6noHnG9lRfbWHCL4c/E5Fh9zs/kDzfdBV
MbqhGYjAsRVfY1ZiUjguVHmqOIwh9gZI9yJtLIfhGfQpT+H0UAe+r4KTsZoe8XoRqfrxyi6IRGYS
c0Pr76j995tU6at0PfD9FwJNcuRZImAtMJkRTvddtX/hlVO6mfPUYYX8nr/PAtgV8wfgJwB4ZaEd
8rAJSC6d6vPwmkWnc6oIP2CqlWLewH9131D2PUtsY+jjqPguRNQsbIXQ4Z+HHCimeS67V68FzJL3
GhxKogwwJjOhblGciH69EHH/GfoPnunTkw5qN8g0jUnw8UTotzfuMkmjxMV3RDefwwUckshlYiP+
UdC14k78+VB2OxjqAoS9GeDIJdEF0d+Dza/rz2UzOYaXqMp0ZSF//3OU3x3R4alD/sgdkXPk/CF5
Hb2v5SE3Oi9kGtl5P6n3uogf6cCVzuJKccu1mOZOgbH+Hb8g5khrVsVhCvj2AjH5e/c3qXLLVL70
PwTJL20HsFbIIWDZqPQH1dg+WVD/s0NS+q3BzdZVQTRKHLQH70slYc3H2D8ifq4nV0zuPB0GzQRJ
ylVYbifA5g1VKBFx6lfkKDsaQX1TlQHgzHgy2ELv0QrjWnJx/jx/gTiVn0IMqpqySuPuw66K4BNg
KkHy9mFS6PUSFUkKzpIHzBsB7C8u/oqVCN1s2fkNfxn/PKXSs+sS71SwAvCDwDFXLZ4bnuvnTQ5H
TZPdo+l5CCNtVcFiTDOeTyvwrKUkhGQCA6/KF19Scvx3mQA7pNyQtdQmrKJGyL7WBzKZ+Fn07ncH
YEWnHdy1pZjV6UVSSDabPsGSHkmes/tJv4X2bFa8LVlXyS0pDTz08QLFdpiX0oZxl75MDc1BBkjw
zcgEFqSPnNSR2LhY2j73M2+xi0FihzYNk1wqvxtHsbz4ecq7H0wKu2PkrRAHA+RpGzLYFNi4yS3E
qDUphWv9AnW4P1jLX3PrqHZAyxpE2BWrI91m3m3kVotEvS+11iBY3CpBbozmtwu5FuhAeccg0NAP
E7PDh1zZK7zehUl///UvbuOXRn0C7yFBsbQb2QubiQsIqLzWNMKXGp+HN+DFY0/d5LywVRUCoZM8
aD9YQRYKVYN75OsOlFw5fanAp4/q43i+Zr0Of6Opjs3OeagSVt5yS32qlBtymgjtpf2IQQznO8i8
XN/00EDjMk7qMj6NAChvibLPb5nmPMFzJvgU4yW4RyPUWHkGw+//8j7MKwhFGH+45Wjc5qeqsgED
dq06qQ0CPROYL5+1WPFIaSUnp9oXUZ74ToFQI9qBpgPTv1f+RzQukqBRnyVQAWnO1BXf4U6zLp68
TNiI9FkD2CS+dBzO8CLVHrP9J1iqQsxQOoSf47f7c5c1GFNtMctN91OisoKjFb9KsG9q4tx2TARn
YzBTSOb326B4NE86x3P+o/H2wrFDwr68IN0C9sRQMH5nBGkUxUe6e9AQf9MZ4x/Eb1SHnPUeNVw1
lFMoibcsmOtP4iswa1WqX8FsHR5AFnR2OAqzCZJm8USneX9kYUNRI10n76q82H2y9vbEJvnU2A0O
PS9K7tJwK7N6gRlbanqIjgUfKfj8kopeMWVnT41PldX0a1HuSKxYTolBjcFkGL3e82miaRn7yNDW
Rr4n4wl/TBRkt06pmfOSwls6UP3I9mcvn9IWw1Ml1uylp6MseqLdKLq252avUzzx8Ch0NTuHpmn9
AA4kRguRHJI+HRRS3eo2nuDca5yzfjrxFOQl18bvgj1GUNCdtYSzRwX7C1qquCJF9l+8pol2Hqun
5fOoNWCLAwwCQ21Vpqg9gqPCw+8C5xB/o4GBPnDIRkB5cKe2QSoKfVrh6/EyNiKsjxOf2LiEHXx8
DxK4KB9klmGCV6Ir8JigAEncqfULXDWT0qwx8JwmMqVf3T6jaJRg4PKWuELTqmEbgjTNj2JJi4H5
Rmf3W/l5VB01M42StzL839LZ+6r90iLir5akb+h8hbfVFx5HksHEu+k4JB+6XG1F+FXbMz3Rd0mA
iA35Z1Gznbgym8GiXOCil1hopBDhNn309w80NnadRKyDq4tLZBIenfHHMIR6fEZ+iw8H6hSgwpPv
pYFqOOw6OT/FabFhlv6vZQ99t8z18Jov94TFdzvrSnjNw+X0i/9YH6okBO6EBg7oPcYAQtlwKwHF
2+VEyooDrf6NOG8nLQauO6ya6Yrhtm2P23UNKi3+3jwEzbA+YvVf0eegmJQsOScTRPRw0+i/ohKU
sCHsk+snLdch83/S5CFRPvCp8d+3cNE9y4Dtbzd1sLOkLIHiMReVgB54HoPyQUR9ZqQRXbcbyK6Q
su2Z3sAXEVw5VZKMTtO2XPmogYW7BUUA8UV6AjVDivZLA1V9j3ArxxHhttSO/5XqcHpAqa1tLY3N
ACFiefrLcEFYqHZ9nQOmzRLEnm+ynC6uji7hOQgsF8VxjNzwbB8yvDfdP9Uuiu3u8r7XtQdYBd6U
PyjRFEYZS5PUi7lPXPrjHFzIvo6yj6Cs/1IJ4/FMn3giUBw79nFF/km1LceF6NlTbYegDWEA5j4q
cLV314Ev2ExMxJj/b+q3m/XIFW4bXOJbzPYUCU8dF7uYeLJsj90xJ6bPGz/17zS3oKSl94WhOdn9
HJDA/kfmTPn34ksDhUUvAtaqiIk9+Xbhjdh2YZlZfCwEHRi8HmioGZkfo2+Kb4TyuMpo1IC/RVo+
Gvb4pSMyI1l358FyfGZ+SGhhZZcaOQ621ROf9A0sUUUFz4jWl+iv3cbvPGw44TpcNXoDP4roXiFz
mwu/k2FPk0s5mvkawpwlX15OJx+UK58lQ5Ms7Yz+l6aFY4MnuyBiNpgClQJDPdJUALIh4oI4Zzhk
84UWmpfhPbeNiIoQDDbVi9VtBrAEP3GUU/7y8WkZ6QPVN7GCUmTn9+kWpg5JPPINheSgzNRdhhfF
kk3pNF8+FP9H7LwWyemqFnciot/Z0wNLw2KSUdEpTKJ9cXx3MF+xpEt1DJsKq4VpH8+3bfrf2Vfc
HMwoMtVZJCp5nrjo9QeDthR6LVKDYGjVitqnCmufSkY00NgPBysUjxopACKnftVoHahpPKYGJZS0
BOrQsJ0zIE60gIiwgFh9L8AYfpx/ydUtDhwzgNgyMxKp20hzQvfIsium1VHeb0JYEzj1Z7/tbEEn
VdGOOzFiloEM/rza2UYPFNLqvX5VFLN4b0FnAF8limUYfVo+x8q+N8kU0k9XQmvzjMS92pZJjSaO
iK8t9kyUBdEpPPaXRMOrUL+3BE38iyjoLjcJuVPkcSACsCtfvwnAnRRyTVB4mmKvmaIxaorHh5W/
zXd8vnZw3ffX0tLkYQgNHLyAFq6aiH767W2N33p4Yv49djRq1x0Vi2PimfSMftajLN/i6pHt74ar
J3R+kDmrQWjRT47BhKafPTfsANwLWrapkvjwlQ8skb3imqnbApU3w9j5EIKTxw/9FWKVFWU5bdkM
+Jo4hP+/G826MpolwweEt3wydq4wO+Ps5dV2wlKa9w+PbOvlc3x9JqEvbRr2JoR76vR5sbGoqyVG
w1kOVAwdqE/2chb5nxx0GzUZ8QVQU/7Jx51Csm7wJejZWWrPG1gCkyf/Rm0blbTRxFFpoxvO/q6Y
pkYRr18w/Xe2k5Y8sXo0imVbuzYsaTM4za5lQw7JN9OcxgtW/zwv0ylFdbVCg+NC6tkGpRr59NtX
lNf1qFdct646TumLqsgUksjPoeruWn3pXrilHRxGW0Ob8b+IYSxaXG8UByiDQP3NEKEXF4HfzasW
11ps0hzxUJWulWunJt0BkP+FrsfczOmiZOn4WGkXAe1dH/1ejMPEjiUOYj+aNaAirFjvcezPPepa
0I/ImYFkIxEyjL+tUJdzxh1MOghau3GXlzVIIviGCc6Q1ehZlPryu+dXIau0qELt+bWnhwkOJc1s
Nakgl+fVFPvORFznehVH5jJgb+qU05R1XjtcLX/6LnDsdkJb+/2Sd3wyQ9nG0lPZPIUZPAaWxakS
iX6Aaz9q3LDe89Xjj1d0HBg3BvrGX+vS4FBaW9nCr80PRG1/UPmWQtB17rcdzFYnU0U4FLFA/qKQ
9Pmb8OScf50qPTwmdpzPmcBw01Sz2Oq+tUmZwvsb204BcWNDxr5wzoep9nGXnLP/zuXUAYMZc4mC
+a9YoYsB+sjVLHacEsQTXCI9Q1f8w0OeM9Vg74W+V2GgnRFQ5SRnDRU7J0AxmVrMNx2pZLqOdZ7F
4ZLQPe0Xs32j+u9y8h8Ynp+fqbqmZTXWdmBIvNMM9WMrir94HbsSaW4UY5niVrSySWGMdlnCJ1GP
TR3lrGImr69qZputuPQcM+BnsWffSFax8WggBqhXW1B1TfxgEtoi8pXBPplExUUASerX67V7t9yC
Lp4WrFSXpWHRzECd8GdAIvNxL+RlNYPkqybRMYcRmnVh5+eYRDuY7bZJHWCloy8USnsyZdQ/LZ4N
v7cIT+nzDYq0Rp/TBUX9TNMoU00A0MLvmPdKKlCOF4f3kKixU9mVkyRcJxd3mku0cnIepX1T036J
eCXXKkotk1OOESdhFspqwWV4NqFF/Dr9EvOxJC2qLduoaiiNSyzVIgh/T/lAu88NBTIiRBCkGzda
u3bZ476l8KOhoauobZFQAOBsanm7tcBgwYu+UZK/XuzrzezcKvwGIkCEMpEMtQiL2wsxvR5cIvRM
VkLf1SyFhT26WFhrXYCDxTlk7TI/t/FsSOMAvr36OHx6PFJRdxgYQZrbCxplYBrnWotw9bAVPtSO
jSB3BWt6dwcZm1a4tPo9zSpzfJjXqxLMP1Dw9yAfWqZh+DgrvZJJu4SocS84L9SYJ8WQJ9hsqWwc
AiTVL5zP9hPUKGkKc9whknlVJ+LXxgqLjz49o7Q1iWYaap8Fe3s4D566neiWVj6TahR+lzAHE1zH
CdD3ax2H5Gg4k5HCnWM/Xgu1glbI/3mcKYwR1FTS3s2HOAVAX8iK74mp8NeHDo9VAGnLoQorvzEl
DYiwpaO24b9w/u3jjKn2K85QNHY2QKLrvXn9/W87NfRg9Y29/U+dUDGHG+Hy6rCeKHknTmsHIFzs
U4u/gxCBsSQAh7xV7Fuqm9UNd0aQL6740q6NNeFYuU+m19yQMcE79gBITPQz8jyDj3yHjgiS7sG7
sD9s4fE8ffMiV4spqSTKPD97UJriFTZbPwFXaCpWdU1fU3sFzpeiMEPMUe0Ht/l5bp3Ggg1zF/SE
q0MTt96/Vp5n6LJA6kYBeeDuwLRzAKyzUz3gq4QhI467E+FySqNbjgseUXN7a8X430EI62dOVwd1
SXraZs/SvwjuX7HX+VK1RJ59PvPXgOSEUtKXR2Qs96MhruYSVQn90RJiDiT/JaUSRa4vdKdrtlmJ
GkDd1EmGf3piSh5mV01L0HsiedA2/q7DOXrvEGDf6K8uvk6gTL77Sek16Q+tt7B2Waylu48WMPe/
IoYtXw+ckMjCO2GOa4sAF6UByDhTEk+vjR3qNhMRyDPGqsUCkQSkB7ceKMeJqYIn7CPvTaOTg/CK
KCvXEKHr2UcKKo/i4TMJr7aN/a5PzzsGtA0SauE83QZUrXYEeSddgcoM6cvh/Dsu6G3Uy0lufJD7
+LrIh8UoXJ1oTRgy1SHIt4tZMEVY4YtNOvhi/CsCP9Nr3sunCqXTiAN242HE3SkIfl9r1u0Z8s0V
tjYFkxEKBT8gkHMIZ1DeGMnmtk2Bjz+/ZFFVxPl5xNDxF1VYgl9rjIYrxwXA9N8DuJWEkkTGaRz4
btliPO7xx7risXzfdlh47BAgwfbo2lRI0T9VeV0y+6Rin8IMEeQ+dmj/cPPjPubCGJuyIkvMdHz9
o0BeS93Ve9SAgO3YgWL/egiCnoO9biSman8J5WiJso2j7RtfkRFVzZwrUs0EgtOYz56WXtyZN4LH
KjnqfHZr/SwVVmYZiye3q0e2zRxjA/dm7uGKFjrinx+Gm08AbuHY5M5o+aa8n47+fxv5kAb6rl05
DW9PAOeCgHrfyUY4udzHGDMLfxqewzdMIpQLju1V+085TAE172kz31nOb2R0gDmrD6w8g8ygUtEd
72B26ffWvNV+m9F9yeNcnoMcLI+XK0LSjZdh8QpmnbFZzwgnM8ui/vfw3/QlZMBIc9tKEPGKmxXY
ndwNmn9ovR77hcl+PxpMZb7VRYk/Cn7pRaeMdYeIlLqXYqQjLZME9jvnM24LgWBpuvLus+7KNiuK
K33K5jqBy5UjLBJFG0+HVjDfPESE6OcrXo/tBvB1zIEHHAf9jVSEym/p1WZ8aJlt6Xh5KOuvi+Fz
GhCL2qLAd1GHLMdCQooJEWA3YxEv+vY4svXJUboKwEaf3pXk/vCUUHdfc9+brM1lpWZPkOizoDIa
NPGZeBHWmYuRn4w6KsoVm2LLN5Zicr2ptvyj0usDN+Z7GU1i0WvT7pdDGJtyEX9Zz6NHTeOKXsj2
tTVrd9CDc/iHKFL0Gb7/2g96RgTjqZgWso0bCDbuOPsE00C2rtjle75YkAX229Zl7l2YpkUergYG
IE7sIZ1pCbT4kdxsJ/baZMbXfY7plRrqb5mAFFr5rUC3KqREVxxus9/fTil8BDYSaKksINoArniG
LhEDLwLdWLgP58yoUH1hsbuL5dDsLh0QMUC6cxiMkhAw/8ZmYFELRt2DCvrriMbmPkheAYSYLU7P
TeGFdxR9+5SJsxTmQuVqgVUIQ9PiZ39Av2+8+F0nG1bM94FFHgf3GfKAj3ZmHpjtW3xJlWqw9maq
SLgD6oQsVLhgJ3xbzfbX/JMSYwJnGUcfd15lAlxiMaBjfAiXP0fccdmXic7lBManhtg2RS/iLj/X
3L0hgj2/iyw2QLjMUoVxbpRyOGLX2v12hxNL/Rd735vjKZbW2jBJiKlmR5gsL2001LRMjad4mi/x
ROzAR8LnUvvUEVdaHPezOphl81PVzpHPBN2gRWJzQHHCqiTFALMhFDv4CyJTeFbNsDJyqzGdrN5b
lV1dKqkopUv/Z8asOi3NWLU3mgzxRS2mF7yarPaa57GIqyOuoKBpQFnlidj0Xc4Mm4lSKbtEgDr0
AjNO8ohGoPq5cvYKOVlfFLevG0VaWx6OK9Ab12CSO2gHm8hlN1X9fh2nUnG1fDaLxqg53Pra/ex/
A3HK8kpUAvLCs0DMCbPacVD77XmUt+qPyXCj6CnWKMFyv8vZJkmpoxA+jO9cPOGCEsmMniVIi8G4
Br1sqWegRTIJ3O5tKaLfy4s/+G/+zqQKdbMIty5KeRQdTO7M9W5oD6/xxpF9Dx/goxpdyHukZ1qR
ySEeeWCDkk0hJLEswzlszb7EW3rHZXcDlJ1bBYfAijIgHvwEMnoJ9picueODjEhhfp7w4xFBhNwF
c9mJS05h4sFR8WDbFNsySvXHaq4OnwaD0Ijlk4Ue1y/taCwg1RQxPmOd4z8IMo+1qzuX8I3MTkAr
vACkccT/rT6b30iOHzRIdnxPkbTNfioPcXA8uSws4aC8L/MtdBXLAveUEv4c7enV6vx4J8Frh2UL
Y+TZ3ZOEnDu4x1u8v4imgcoSXh0H6ynApcPjfp4ssBl05+QTbhUB6BBjD+xHsqAFhNsQnP948H9q
HBqehGUltQEpwhI8HKT85xrTtLW1f0yU5nJmSYznVZn2rKVPRE0bHya3TcWJTZuV6ehx0bBo3+wI
B05u3rSPPOXK4EH9g/yRLV3gaGbMI8UC8rEb1CMpAuwhl9eMp5tTrpkBLDBuNvUlOEREMbOeV3vz
AvZBYGX9BspvckAGCyEiofVZmV1L70Sidg1xITtFMzF9hM7A0gDXLkvTLkUMqEd35xr0h9m6BUL1
VW9R72TaQXQDVn9Khc412zp2rZu9PhhXpgPgWSoTWtHIZhFadb5TUtzfZg1t66t26t9jvjl5VB6P
CaH4gj8apzUCFaCkXrHPMSc9gU4MlQOB+Vvz3hJyREc6atbF8aqyHf0AzRzVJTdBNoHKDha7xoRu
ynXq80gzXQqSzx/c+3WHkA0f1BppUo0VZE1WPzjoYvlUhjVvNwnovCiHIzD48cjaz96hgcwMVVu8
yy8Nqj/al+O4U7ppk858Jmut5l3jTjMdweoMq8k7i+4k288NsI6wk4RenvUttuNTilDN5E96NLrU
DTJnxEKqnc9jpK7GSpBnTmuY8Fg5WQxerDjA782Zvi1rYhz5JUuoCDttJjwXUaj3r/sX/QlpHP45
BsRMaJ/JlAamMX7iDZya973Vl7LvO+M/UQfcvzUa+CU5nuRD87BGheyxA9/xdoG8tgwNFrgmdLYt
Og9lkIbspXnO2Q642Si3q6JyIsBrkuoTU8G0jaGPfBchmzFHDKFP+dbcXOI4qWOPNGw2R3uD0afx
G6F3ugSRTXWRTFGUe/YXf50xMIdiLWkW4l4uJYq9hbUBoWpLCzWPCNnpQhZG7enseTWNQ6bQ/KPa
cWOlVEGuZb+IuTSYZAF1f1EfeavmS2Lh+RLU16teNLs4b/Bg2mqD+lpwre5PmQWuhBpmTtoehTln
Sf4MsDJT7vHciHmKCSAva7yf6TyLih35KYdy1X5ckEIGQ+xR7GPEggSc2pPSTNEJd7WuUf2TI6WA
2LmlH3YQ389bfI/vA6KZIiH4OYPxeWJIdVT8F58gs6i1MgHujQqMMAQ0c35bDg1oyIW0xfsUdqfQ
O8Q52zYWQ9tfzB9izgTpDpg+fvHSjjuF0ffQUQGLF+EXw95G4/UyCKst4jpuHsEOEHSODSCT0Ym4
P1Bwr0EVu6Fs0ZtY/+KlGE4jlZDG6fBen451TewROTkdeaADupyU51+XV30D9KEz2A4FTs41rXSC
2F59MjRHxW2HytKW8fYx9lhUYxj5bwq/82mfx3gwWmFpFH6+TDGNlpnBmBSTRq2Oq3LzVgtF5FXj
73guRbduoAN80i9IfVWkQHEStDXA8piww8Pn3ujCw73mZadnRRMrrBwojJAgtsOssy8NN+o+meex
tpfaVVIxJ1Uos/1TUvZen/MLNsIRrikbXmit97XzchzXcU6/5DGic1pS6ZX/Pw1nYaL8m/HBpPFt
sN/VODmqtaUWt99cl8I3N1MH/pUf+97N0FVD7oVj/mesPOLzjU4Nty+ZNRV30GncG5YXsaInHtIN
2LYS9Gb1jbPywMbVfD0vw81P33oYlihyx+LjsHpLcDdxoGtxXF1yYKSd3/ZsKlyKYYQkWny4t64n
6viB3E1nHrxcYSodDmfgo/G7JfNI5/zhyFmUnpwsmadzqJwN7z1lBCumS34JyDzbGXPXj7XQHmMW
R6OAe7LBPFaVKJxcF38aqBLK6LBmvMp2cZD/rqf+8R4oXG+62I2S1epgR1AR94hIt8SYvnQRJmz2
/51Uhm3tsCjW+LLl1DYuXNcSxDgnLZOIwt+NyCczXGYZAHDqVgcRx01Qsl5Kg4vCXo9+oqVnTGSU
GE9vkFoXSZWB31dj8u6WLkFfQybSTOToz3geCSyB4ZarZZku4OERCpVBeJ3IR+jNlX/f8o1v/Ozz
hRQ2Cdv3k0dpWyR7ixUNekLNoWq+ukFuxrarZToIPQK1VhodBFw3XXIsTGIZTejWkuO/XUsu4Ejs
qAJDWD/kBT4R8SI/wtkTArsw0TLLEyq12Oz+mr+kp1WtNlP6mLPZ/uVqmyOnP8cgD5nrsyzyMlOu
+yklOSsgd9/e62+wqNzGPVCDTom6IM7I7U00WzUYytLYy2LAOG+0cs/S+iy64s22oXwz9Ixb+Lkf
KcNjk312qaeYLGCAKqiU1lGD2XoJqouZEchxxxyAigXCEAaHm9lffP2Jq37b2hlpRSTAxs7Neybf
K2PRHzCEP49KNY53QGmFjEnaLrnaTpmgJpw/585lWtLQHgI/YnL4EypObOdduWyrad/Y/8StRyme
O3j7ZLYl3I002GAVzSMCz9ESPBjChVhan9XuhiUkG1tWCgtD8WGCHPUqLZbY1U55YS/ns65Kq1rk
JXz9gTGvyVwYIamqtyLbPaVWi04/EO+IZXBS8fn2RGH3bzGvg59x9UNp9sbAONmOdMibkX6/CrmH
1eiP/LzXCFlErkbrqL4f01dy3Hx7sfuNPzEYuyruHkZDEz6i6CFu6cIt3zAc6Bm1tu+q2nb3U3Cx
Vde0vZQJJYaLSBDViMyHNIHh9BpNsLnoLm60J+j0kmOJprWUsk1hHuD1cggZ0VtAmYyHxpGZVliz
G5fV6X0sZ3vOYvYFtHGBlLC+YWgNN7SuXD+FabmHI4KfUzhp+p/4TMaPDzHr3gkSyuTVdbpRNr1u
OQA0PkO7f04Qo8yxSMwpDSpd2J1YxkK0Gg1ASM9n1bUCPKefb9gYNY/lo++WoBcWEhKWLEHssBjz
HAfdDSYWrWjkucxNYxir+1Xk42zF9pUAkpa+LHLcvB0Oi/eolGSybPjj+hST+8kfuQPJQoYBuQph
9MKsA4nLC96mb1BLDeF9El9j5LPBaiT8ES+VL2TMh5VHkL4ioaUdZtSC++OJY+ORyF/RTq/YsASA
+kO6hHwCnIbvkmNYuL0sRxunXbsDzbpMiesDehlKrV8YvTW31BqpDpw5TKtAkW4d6keJ3z287BIW
AR8qUYxpx25NO72vJAV3hkt+4iIActwVu594EWQ07lW5KGLeJsoXXHdiy+Rq1itN02g47CpjHOj8
I86X4eEsyYu8mmTYD4ublWJMMs48pOxCGGveDwkQ1krEV6pXy/tvG6LnOf69gw0adRnkBJVqoQqj
dxY0y3L7VYuJcN80oOFQpm18+ZfEk5pwhXNnXClcyz4H5165GZg3I1KJhpJGhS13rXXr1Fb6+8np
zgjW5qkhssdzM09SfIaPKxIpZUSNuEmHu2qsLFkL/gZe/tB6so90ijM+eMJVOGiu33BcDpCttMT9
haLzjK/s5PYGZXehgXCjVL40PsTa84z25hoH5tF+vhPLQ0/3OaRXcq1uV6rtBglFrynqtUYvevQz
Wnu0KuT1+yJJSLWp3sXO8IO2zSmOsISNepex6ocoDK7+9O5ilYqyqdy+MtjqaHfWCwe9pYADben6
Axsv23ayBN2NXYG67/z3VHEx0qB5faUhEtgrePpFDnu/a4uVW0eUOv0dlrOWy/pj/pMbDXj6ify3
rzQ534/lXSmumZs91GP0e4F7GQetTBe9v/vl4tniRuwI1A2eBg/0gPizTBlA7jcdmo8EsFtSAI6T
vUo/0BZmI+3v4vD5nEgskqc00tyItvEaYlFbX6TFmaM5Hq4ckcYQPhOaVuELZD094gR5AYYWlKmR
zjrbcBg6FMQWTh4T8qCNaUI7ExbT4ILI8RJmGgejRqEhxidUU3dRi4O7XiTKgDtoWtpegnjg1PQg
XCynU0Gs/IsyVYlMvsQsg5s+/DA0Kw4ResnYShohcWqZKZiL1EPz/9bwngPu0mAra1F7WLY3jH2E
3cQcEPQqy6P3NlD058lYzyn67sTKJkn0I1OdzvC2P22LgZM2YoYU5fIC9MCWndGsAXpmf6gUknLs
9LBu9ye8BBh3ynbXij1B6FsTr4jc0IhFi1a+Bf17j/ATSfcbIeRmXRWfJ0IfH23wFpxxI4QhALZo
me2kYszf53kSehisCf1eUaU9YciiCO9Hw06X+EgXDY8EokmPyE8o7oNTjeiCFLNN3oLBpb8BP83O
TA1t+T8CYAHjcHMo8clCtA1KhQu0zrf/NROpkI5tHVenZEBAt5auCJqBwG9dHdNBSMy0AvIJbZ37
wFJI74haAozrePVR2eW0B6U//BFC9QdFUoc+bdL7ZwFYJMmJdCq6YFEmpocXq3f70gs3Jpuvq0/M
8EuKl4xgvwre4rqFG0YC3JwqQu4LNXI4ZhOBJycFVpKjHYLw8+aVKhaO6cNFHv7F7OyrI/SC2t2Q
7F9BkXS6fpvqRpFC4d32Z5UjsQbAy/N2G0z1CsUa2FzW6u/AYWeNynzknGUEDALcgLNRvTflV5j/
ll+njGWjB3KWXmtto3UuHMWycyTXNZAzLEMRIX+4xJ272vBQkRVy/IqDOIPFwn7l7ISeEjRo7xz7
SjuC3bq9Lk3lOKozzkJZ+0a7iM8D6Yn+DPNNGiwyFJa+coSr8KFHHLQYEqiwSGEwpxMf3Dx1AE4E
KeQgS+29jMATzB3ffgWxcuPezUp1S4n3eAH/pS9SnZ0WRhEqM7qKMj5TRxlp/Cgm1a1gEvh9Ik+P
653mTkQP8yTZlLv7r7GxAxa3xMw2+5SQC3cit0pPmbnvtiCWaIr9GCzkGylc/9IfGARJ+zSRkOOz
PsHOBKbYMqNCyOWqlZjefKIzG6nXLfpV8QOqYdXb+F+xaUvkhAwkf5PYmHyACOgv3/9cxPKfqxzQ
3UY2k7qNi0jB/Df0GxN4VHLZQPFbhOtKtt+ZAMrE4ypwdLkJa1QTDXluyW0WZZ7RTMEAocvCNhLi
V5zHBlxvQT6jm9KyUbKqQSY5vHUBEo1QzPlCyNXlQf7gxwK58cEU6xki89aTRMKeWuoJvIfeQ+l7
8oDK3r945loKwLRtMhnrU8DJ9lYPEJLEAXTIIFBE+J/rlhAKAJ1xU6cCho9QZ2nyZd7v38GnJ+AA
fCZBZfMiD9LEbtsmB/7HHnF+WLa6L+bm8PN5ylgQU7SYgjBCZi4BicfIpycBsHbpj3eywJ0jLBdY
1uywSTIylvt5j+kNJJYXCDzOLQAQ5TVVFd/ppmY8HoMk+ObpmnlZO7Fa6gDfBa6fQsE7jqEXYY+W
jb5cvHx5z6tdekIZjPh3dpd/pMJoHsJmWetNh/cE6vf8wYkOXP1mNUVgu/d+ht7FtL+AUYIPuqD/
/CJvK9J5STKEjSwwMYMINN9AsQFK2XXbouUpLTTaSaUWtYn4Kt2N8xFVITTXp7rwqlYOgDVOmVLN
pYUOCWfcsypCJRtmtK05Vhtw0UwJ0USyp5nawPKDWK5ETmUvUJ4FzdeyC5qqezhvx8pmRGhkIYKh
cR3ox4+KLqNY/nwnOvqxAQ1jsJ/yEbX9rYoEp3AYzpbnSoQ+2CAmcp1rS3G2iadM5X33XQgTKGvm
uRtVjO6Oj9iVKcQD8XCT1zZzIxs9ePBkKnBrg6SQ+cJZkJSk+4XXVLsy8YL0Q1PvaqzY661i6s9y
AMkuhIMdeoGVzXo+WN1Iook7xKrKxMEFQ2F3vP8cBnpmjQysXpT8IDAK4ZsD5Y0WCpvdAtLkmsqm
fwiDnr0QpUL5wsTOtRDEB8dj9r32LgC0BIxzjajUZBobk/1yKumy+rl8CPwVocUhG545Zwy/G522
8pWdGToZvXJYI0duU3RDCfzBofVbBYdSFdWAwMGN9JhhFWUewLX3WdG35TkyT3b44GtkqvXXr0P1
XCXWkf9hMhxenbHZB+K9L9vFiJsarGTpseFDh8bL89oJV8tHr2TzmRciaItXlq8hqc/H14GAIQZ8
WZoWDLadBC9VBauX/9f0ZR6hDCv/pL4NmaGerZ8yG44QD+nEGNYaaNSrWJwGm4u6h2V0SLpF4y+P
wKLDnGCS49aA8oG94NczCOnthwjqmIHUCq18MOnWNoVwNc/WxcVrnPcQtsYGW6MUI5aD/g0yXHdn
M0pwBb8YqBxHgUyOJ1fgkC34PrdDEc3YQfobtU4KNGUeFg1hYVdU7LjA1Vrd4Pgp5fHk82+Hpj20
24WrOFf+Y7VHSRWXGMYHFR8Hab13Gpgu1Mur0QzGBM9LtUi9YA/8PdyMsrJDpWYi7njLedm5yYK5
AVjJl73Gf2r751Cc9ZoIsjFY0nTBnXSZegWyCwNTY8nOXa4UMM8qP7fSxQd/+urpjIugtlDoT2IR
YmkFV43wW8GLyH+J3gcYYks0rvFu8spAELXzzxkWAyPsuyzNttatcDGBcoLrMbFEFarG8qc70TPn
wwD5vA4BAcAAQjSw3BFRBku0oV+Llqm0CxwTr573H03nxw+wrdC/QhKbVc6rJpnEd0340Ozft9bi
CieWDPB/skiR7e/j1sRtfpLOSVXw3E9/oeLTAlzCDjpyFPlyumjJl6mnFvflMbN/IaNYkcsWs8ai
dbl/LKo2rCGCpr0NrVAvl6Em7yTFEWrNsK0pFtshuGSWH6ScmA5trdksqe3DVex8xvxcmFjCwcSh
B3t32CBQu8yVzvyqOiY/2t9iflK0h0PGj13szKseW063VbAAoKDwjkCMDZWiezwABqpQjeDkEf3V
USNnYD2fL6jit8qfXobdayg+qtw9w+O+QkJ5b+qyXXw/B04E7F7PQTojii0NakKJE9S872guPnjF
1uzv/ajFyj9xBrHlvX3bwwY+gPpEocMY0hcoh6Xl0K/kQTMPT95o0qg4AD7OpaRtiUtwet9Avtva
bShnP1C9esBn4bxXsqZXxeAsjiPtS2ldIHjUHR3QKfJWuJYb/5Dccsk+H6vE/nHGoFrg3RrMHXRQ
mhKniZTkrOzDeKHevZZZKl+gqkz96ufnEGUo1PgZ4CyKfan8MGeoalilSy+P0HeEWggpzZguXNRU
1iSIpT0vvGYefCmWvSao+FQhdNZitsVbWB9/EHFAkzDpqaIRnfzPpS57bTNltopzDxzz9RWnEp/Y
WEarynKBe8b3FBkJij7/qbodfPM2ce3JJUXA2L5Gc1f9mjR5u2JhkihUH5IsyOqsqYnOglzQ9uQQ
r9I+eI6ZnwQihkXOj+V2ZLoB7pXAoYdz+hTi4tXfq7IBnsKrvLPPAvsypSFQBRtUAl+cmawepu4Z
bTd8xK/kDCcMbCPtw0Rdtpez0gizK670fuOnsdZrnaDBbLC/s1U5ujNtlt067V6acRRy6scs/HdJ
Szva/aLR2yUNv64f3Y6pxdTxRsjev5N2IqGqFq34M3XV4XE+pvbSmW3InD0A7SMsq4SN0m23WtgX
qSDwqYDWJlsFeiuHYQtXxO49yUGZrOw3AFvLpgsWPzXaxtmxDYncpeKHdrmVKwGQw0gxlic3RnLA
H5Sp9a+lCYQreoVR4PQ5tN4j1Q/7nQGzOH40LxQnBQMr2Q4LqVo4THkmDMfff3uD/disRP/pCROe
BxBiihCPqel3FYVQ1zmbfBaOiueXy8wSMZk39gh+oGxk1m2Y0XYi6gxs/x2Pz49j5VX1Im7NMz/8
wtS42iUqyztH7h3x+u5BL5mPQL4qmazBoyWFwQowQvWzN6nbm6eUTxSQpTTxjvyTnW7mnCfB6xXI
J4lyBbxZ2xVHM9WSblxwIqWpyoExA7keG62imiX79385ku37BmQlqiIxN10YQ/bKKj4EBN4I4TMQ
PHKQSRxqStNeqsBVpbTV32vYxq1qe3UHCMZ8bKxydMOvE3m57o1wGUvrf+oM3hcwUt9o5aShdYER
igkgHMOfhX05zFYrVV0058FbxKKFJnz9SCYP2CT9VjqayRUXxGSmrJ4Kn7xq7VY/6HjOULtC0vp9
tEAkMBijmynYECQhz1GVERLkgBgZl+nTXL7bQzKio9V2ynT+hQaAhE5NHT+OLsv7DYT0KXuDcN2i
Zf2ln5qtCpofvM0TIMBSrkXoRDnhjNzaAtnC46+mVE6314cf1vUWsdNt57FoKAwLSR0QY/zV7vIo
QwBM7G4m3oUsnfKHEQJmeI41pwqG9NOp2NqL9cTdRM/Fxmnl54NMDQxS745MMMH4gGezCEUfdohX
ojkvLftsJlyXsfH0swZEC76+BybMcl99H36JG35V3WiZWF8dMspCr1m11A/vZ8uF14NNBcrq63CQ
8H4SjDk2yA3iae9E+/fDML6CeHxFgnXsmjt5LJjHvOVx6aUe4RE8e0FOy4qwMDfnAZEHmKqxFsQm
r/ciSGSP3GQH41MC/h9jeLnax7AvT2Ozslodx6mISRnYFF4Kk+LRxOMOmK/1OGKQLDupFT4y94Z5
19m9jTcFquxZmcbwcZrO+JeJNjwTG1fP7kYvfLga+roPtE+7zFpPELbsX2CGRxxNueAcIaHGxU11
S48aInYV5LdnSY9V+OLZSyzdV47Z3hl7kmjkSVeyc6212km+iMSxLuedbwh66fA1vGS9DYupABNw
XQSvkTDtyuTSvP3OMHhjXt1SJ8VIJ+54A4sRaxmF3++uwYPWhpepIo8YAbbXeTuWHCsIfSKuxy5g
IpbsQ/O1XJ75kAIEXYW55QR4Rf0/laMmYYisltTrfkNAllnlrkAfP8eVXiNSa2XgHt/NMX49ZCaY
23EL28MmIlcZ7srFmKCchXA1WkiIztsNf36N/wd8x7hgvFysdHOnxDx6mk1x5SiUlBTQvYsqgXtN
r2xaQI6QI3tY72WMVKB039RjQIE3StzuXMDK5ikL4ku5ZM6ArLJSLRwaXLB70sehxvgcDvPbJVLa
GuE0Du2mXnZ5f80QSHtB97oTY+GQVeFtnDO3pLbrz5pDwYvbhqHbZbNyv7pDQjLXKj/RKQw9SILx
bZOV5SRfFS6oBCbne9p4bJwn1hUcffQY8/qOWpOElXUlNdGIGLYLnKJ5FL7SyPdadoF+yCqHSvm5
dNUQBTg+iGM5Drh24DO3qr/UfVM5MLkVZg90iwp9Cg7YDl72nMat2dvYwQq0i9LVidcgl/GZ0bCH
SKThbbiZNhjLBgSeyIzUWbch5zT8h0GlMqXaqIAT5kvfppzbk4CCiJzzG/wso8FVLtrYOc3UBK8Q
shK5eEafgRfaWkuZnW3kEML12SyqAXp1U/i1xoz+QVvRCOHmWXRaPo8sMBepk3wauvXLg8VtV+Tj
4/hqw4H8h+USixMFF82t9F9NIkdTAJRBVuOIgVACqG4hnGK6849JgX2UNkktE9lwmtfvn6Co4OSD
HRZe+H1jvuWyYgToM7teSpBUgIKz4Bsf/gguidARbj23Xv1oNqbtYO355yaoyev21Yqxx2AmsHL5
U5sqOuFy7Rr/kfMiBHg0HCyPc5BnVQYpYzP5egzLzYNmw1I460UT5BKMggQvKGQuakqJlwFO5Lo/
MmGtdlVz9XHhLZDYyiLBrZScF2s6iRh209MAk6DSpTAPgf3sU381VfHv18fIHi8vdV/xqyyOHFgU
6G6nA+gEBR/S7FKbYgoRrCS8U20j21H4kxRT9/XhfVYTBbTU/gfpLKd7Py2UzmvG/IdBPTVRByrp
nFJGDMMhY3uWV+bxXoBh7gGe833sjL1uQUwR0VEWXnBKz5X2EsqXRWmV8HqORkxIJkIm+vxJ88s4
xzXSXsDVxg557BJQCBiIn3+XKzQsgeDBezrpeaz6f2XOaA+LPd0TUt+D8NFheDbVeyOcBGQk18ix
xHxztww2sZmXU9X3mshhENW9lUEtvi9rIDg157NTOGyK5lXudV2faCNdKGnWwkkxOSLX74/5+pFe
4XPrpWNRv20MWbo9SjBdLlbER5sJYGFR1IkjqcUiOsZ2l/Axy4ynvzKpUTCsGWChK1Lntc6Rh8Jr
Rx84cDqBETw8Dyxh0hwZwGvEHgarh3xnfV9eVFnCuhq7tm+h7Dyz52MarScFg6Jgu7v5uwhdhW38
k/dk5nIM04w23YaqDqqTDaPDz4bS5B7gIxOw5Uid2SzXHZzUFXr9NxZC1kgknERXnggcb6HcpJcY
+hpvkHLy3r9TT8qQI1Furi+VvuUP6UNy089UNmfY7JT6J6oEo9R+A1d8F2bVo7Qf1J0swMlLCwyG
ErqXCkeDNzmL0GIHBP6hMZOmkYRj4Bb1V/0Ao+EHOMHubVecWe2MWjFITjsZTKLzrlcSZeXw9TVJ
5SczeYbCbQZ1zTRZhAyEOliscukOL/UTmCLD4txAqZ+UawKu0+cq9KvodCswAqZEZtLwOgtusgb/
bQTPJ3OQPveAzLB3IBAFQHIXL4YGrYUJiPgR0cr/wOg3omplL/UIKvc8CQj3mR0FxFSBbt4X7RPf
ijjDBNbNa47D0iwY+1dqKWmpfiX+dy+6ybjrj4pgl3IVXF6Nm413DrZEEcszgeVEondg8ZgStDaL
kIe962G4SNoIx9Iv9BU1cpAnK5PGOpXUyy/Mok9r8dR9PWCyAcj/oKTL7nyE+NwNarQVgWXeQocJ
0fToV2PzImfP3GqhnzcjS0RYiXKqwHqLO2Sfj9K/xWSTZgjkW4RCnC31CS4sUJkm9WBcRcRC5EV3
Vc61n+fVxMZ8P1/Bb+A2eToP3XPcxKI8uYzn7T2inwOR6wDPbreY9N6L0JGKRimhA1B7NGTNfyev
ySpqb9P5wj7JDiVoDYieZoEDQ1KFoiJnxzV/sL2dGJ4Rn7pYmwmdRFVnEqPRB2j2nPwdUMzVUSOu
clC6tgVf+VVnwFICM7oMMcN6u/LC+YiEPoPkAfpDVt2NKiikpYs2wHNJAEdflNCns/25/lvltakP
KrqCkbrUGS3259zQWhggTJ7Xy657xVyxCAVyAzJaunqZYKsiP2WxWnqwZYIu/6yB3ZCifbfC4DZJ
nZFv6RnPr8GrMOsqc/RAFMFOWlxEalIEgFjI/Qmr/wt6P/MUGIP4Qti5u8bJREO18ZOwBId1eUm6
B8O53xHS5b6y4T0UIfH0XodHB5aNvX2ucz2HRS2O4EaWo9BEJCp1jj3tdlUnXokYwPxjoMLlGRf5
c7leAaeZrWjUY8FUTEFXClvwY/fJu4FkHtedNMPGHq1CODEw4Sqv3c00khKtBkU0IcGkv1WtPg1/
z4WAn27+3C/cQEwNrrJzxtY3N9ISC1cUUxu0zeWN4NxqYd6agZVdSq/GUOMQ2nvng9ew7T+s1xz9
Pzs+9hi4SMCFiGFt0vFHPSPp1CMpBzxv0T5BKspO4dxvoDVsli9Mei0psu6Krm+0CLDBvVVn4rpl
tlUdwLbaf4W5fQlmMRR+mTNhmDA41mJtNKBmaPqGHqXPgNkxksNO0lHC0nLirSE7JyaEgnxLNYtT
z4it+J6NuOwCwmmg/15x+sHXI3diyqKo/ilO+6fk/Dz3XoMOqeVFl5n/3k2TjPmZjHH3gAII1lqH
D5aYes7bxbxVvpDmw+cpeTylMbhx6okXzJBCEZmlFbPq8pQ+lylpZGNsPpK8pM7mnhRg+X9NiS4w
HZH2h48w6MYZrTTkLi2DnE/LDYSDjSCrTpTznAB1ip3bncB0F9/J9wl85jlH7WBFi0gv9qiOzro/
8c0LuCFcAfe9t55xptbBboNCCQ3SAj3O2aBbUQhCTOQwI3BBoishwkWSHkBzGk1qsNzN+0nx4Aoe
fng1DoOEJKxnhPHNQstj0+jieMvaTqMvHkDRMjSoDjD1pDK/H8nwqRb7DTVtzrCKD+NyzWKelpQm
9KsqKKNdex10eK4gMSyCP3bAZW1KBKOX0Fmf29uqF0RkEkVPQ2ek0tLoEgIiLmrCucB68iJKdB5v
D/zJYgFEQQs5dNjvOAGtO23jAeJlkQZ56femViuqrt1tHpQff8JdpUvqNvPaI/W9M4QmHtOyUMRj
9FbvG4DEqQpUwN5hMqzYbFPLTKiFIxEJGU1bfEgXh7A1WgOQG4u1fAv51qRKuuq2rV3pMIboPcc+
Pf11hikhU/FAr7JsOTUjscOfseIxJCLismmv6PecXkZlLWH+5RQyC/t6JaDo2S5WA1JRyp2kfB6T
iGWyNO2ROvZ045qey7h92g4LOxaORBdHwTYxTGl652o+Z4Nu70ygXvs6EqQ2U0/ZMtPPWlcj0e7v
+BUnyDeDwnjX4glAA5GqAWZyGzCyXf6Kf90EXNrX0KTEWBvyduKyr6++8PJsINn29QJa3Xokf3S2
a8XCaDQxpKsSVSNK5saRI9trWKIXe6yHhWTKf/mGlk50Jg2LgM6G0XUe/QvYf24tQBmfbjvby0a8
VcjI9EF1+xSyhCXBINYsmc+1YkIhwAtl0oIqpA34j4rbdTX5/uYGXrVq91n0hEokgg50N+sdIQHr
Ske5azaoOyeHeKpBKg4pvPVc1bI7vxI5fiziq+TG24zBxGwT48jiIo5D9W5eSmURHE1EzIG1dMRK
6Jjl3LPXgncGdpk0rIVj+aL01TIiO3moTYGLdmPDsI2JWnpJ8TJjsyFUrczQ2BgAgqQU0aGvwQ+R
lx9VC68Y9xfesHpG9EY7R//uWr4KwOYOc5QBrZe0yB5HaILu65eOm1l94BgarTdoRWz8mTbIixgd
wHhEBTpBLCxdhKPS/OvOQ0kLkEYfvFjJOdfhf8jTK2PLO3o76jWQSFtcI8IG+P8ArXcN4OTevJF2
50lGAuO5t6taixATjfHSQLis+vLWsjpT2C9QYxfzbFEHjgVfwrojbR3Up+ydbm1WZZrxJ7YNC1oQ
0toyyC2cQhMl4cBtqVyyCCz2cZJEVB8H8xMS4tQZNDnMZ7pR/nW2wTRAf2MJNvTa3HzHaNC1YHr3
Y4jl/t0TGArHzyulOT5fGFJw/h6kKoDJCibjtL55RrcKmGRKUkQ7V5u6wwyagoDm2W1IWvrueZfo
gjsVBFrgRA14moTBJA6oLeyQ2j88byWg3/VMWGgb1Y8xmjOF20FYfztpAyFghl/+ZzxTsByI8+Wf
yRgMcwom3IE/PkardOZLrDrY0qd8KyelIB2uXfYVrOSm1Y4lxnonJyChKuBcPao63WibF0/y6gqQ
VM4Dskg121E/PSqvNyOWbBcmvGk7uMcQlj4JAJS9UBHc/5ar8B9QZ3asS8/wDHOkJJ15ICz8fS4y
O5kWgblWfNuuzD4t15xTvf5mxXjZDorIkn/RQACE811AEANkyZsWoc/L+/uuPcxyfmMuPfhR+S7O
fr32DGRaAlkP5pf8x7dNEg6w/2EqTLKxSMyyCXD9Q7hrA4FlHm/9r3lZcHqXA+weuzYt8pxhPN6b
dP7fzgGtQIZqPT1nOotkeHFL1oD+7ihWkTYsXlEDDz3PiTPKVijNkdpo8/g7zx7N9iDGkqfFCnD0
aqetFhYC03injH4EmSrh5v5s6mJzioh8GOborcVV1HF0KTqGt9QBFxFlm6KCWSzP8hhTW4T1alJ2
ExGkMG852iLrmAjTWcJ1sLoxHo+GTRlmghFyZ7vkPl6n2H7C9thCFrcwwp2LVGPACn6STOlR7Al/
A5F/AtUg+VyODhcnpsSdlj2PCwxXjdyyIvfPpdFjBrqstKe9+nsCwF9LymaT9LFbbRSdC1miLf8g
Io+zgOUeQl3vFZJiMIn4sXd3DJUiQg3+ng3pFnRQ5US4an6pLc4fSImVeWaRhxmrKCaBZ+csB8UY
WPHKZ1u2mns94diNsI0CKWE71JB3ZAzgVnbRGKBX2qD/XBum8fFXBItEKtyhBKtdfinWiCtylHwh
4MUnG17+dJTnES6utXQEBP1SDhNT1X2GdQ2bNHh/bWMmh19bDyg6ZXx6bWh9pFwOoRZUFB+7FthJ
xeVVvEkRW8UZRAM83Kyvwh3+kyhT8ibNYnmPgZnvN2RcRLAZc9mgHCaLF2LpGuPasrx2w0KezPM3
GgsSCAkrNADDvaV2FROTCVZ6epEv4cj/nFrBIpA9rLCkifZGbZlA48nkrLPcSD8RXpyFityFIcYG
38hETRhs0NT6J0kKzpXzLWmUGRz7XwEOwyxWZWa5I5EK4j3rDXn2G1PWjZICbC9BzX/d8ezYDwsA
rhklW73P68B+W9JsJVA3h4cuJRii/DEtbq0r3utEoLOTKznNmX65otCPIzdttygiZT3tsuET6RMp
Svr7xyWvxRcGRdE/HSxswIm7WUwgkGAxV7eSSn+SPIQlOPB9uAvk3B+B5RXpcB6kdFraK7PdNwpW
vGiFpeb1W7vqoFvAel9nrmBhYLxehlCS5gJpr3fc5ykVeI7QmYt9/pzX+a83j42TfTQsqAc0HNia
OY+rRq5SzqeWN0QDn3KNKDMcmZwkHnIGxbcPuCtrOT5A8tWBsEJvHBc7S1mRauD3CnFdBPRIA+ED
nhnCKS+XMGwfmKGJsUB5bFEUhiU4ThD1en01i7NPwVsADu+GenbmWZaPMePQFoNuC+ylKD7iIRUZ
hDioNq34LoFw5e7cJY1Tsl5WI+xGw50Fs9AcW6xVwY18pRcRtP96wVP439e3GVfddjxiE5u9QuNz
6wqwOYS+5/uONht46Y5FemgItwSrYpF+Iqish9ZAXSfKcCW+Q923veRsR969BdwoQf8ysAnKcbSY
FyARKrjGSEdCrT+TthuJIDK+DRqT2JrV4VoQt1Rs8q+YFMM4M8vuP6RWjEPfGTPFZZW+srggGRJz
FCx7AhPJFXHMrAiD27scoGcyXdGrhQ3znSW9QOqGnRRSqN/dTW3bZLtIbTQaNDJX12G++rOv7Tcc
li62AbHhJeelPh0KP41Lxf8vGbuVj84YHztQ5NtSUe3g1D5K+Vj6gzSawTErEkwIygsuA4p9unbR
DP2dwVib1eAhw0wUjl6biRvQfQguJ2ZAE3gJIse4T7Gsj/MOjyWZZTqqoBmSgg5HsOIOJqp57gxX
mUF3Vi+AN9jsxLAYO0d1s7r9D1hq6g+C+KK6K6FMJSMB5611FMeSf50eKVxbE4tnJiGo2hIEYBaj
El8OzgJ4MokUPl+AUwE4fK/xSbt08+qWROnWrdShOIhnE/KJf5KvLQip8qOaPUmDdToXT8rkYqud
O+XDerxSmnblZ3kslvsIN7HCczEwi/Sn+x2PhOK6Zdrg5uDXWoMdMihnbABdV4OhBqU6aPm5yeN3
XDCYdL6ezKBvt6o1U0eRCXp71seRdHGY9qM8v/VZR8xOZYeKiUfSUXRHj6D3ohXYoOT4885WYr6C
i/oYo4/E03m4ciumMD1aELpjWVipzFkyf8aKO6EeGrbir1yx+cJtV7B6etEjXao+DHvrwDhFZFrf
UoCrFu6q/Ib/2D9v7h3Ns2UyKb5CIeaTT91GN30RKeVa7Glb//m+Gau+obmoGXhoCuztXm+/PD2M
ZDBrtHdbbztOBolAHTlYMJHErmm5n++63QNRTyxzZarF+Rc7FoZbubKFTdnYzbWSFbMkEWzxPraJ
J6Vru1sp8b/ON76OzQ9KU+EJwOOEzryU+so8OilAQjeleVdVBce4WU+g6eaXD+ic1Di13p4BLs/7
eHT1a9q1u2GfJYatxYRvY8GnOaQjyZRicsbOWCDrAP6hdyyMJ83R39WwQaccOHUx05nH30tf/qBp
bZIBGYgbEk3qwUBtqMLpRhg6YP7Vaqrd/ozXaXd/nS3VKqWXMx5sz9dX2YhomR4OYbUTwLwUrBm6
l8zNLlGFCs+oqO3FO5ewIcz0rFxHiOHW8xrfMokxCGXi6YXyyy0mpUHzArAgl43NcTNGkwPzhZRA
OutsuqSknu4rQzvYARDaIrBTKIOUEeBPKTYJ0YWQX4bopK5DkxRgRyzDzNmLv8XfmQFI18gGQYlp
oy/4JbO5NnxJjz3w/YYVG8diFv01v+BygiSWL5/z1KazYP8+uDxmFHRA6C+HQXlAAXiQdNfHDRnR
ePvnDSVUdVQrWLmGICOXPMPw1yW8XeprJoTuUa5lz04Q6SjfMj7viBkfxllyZN11ogTE0wxGsoWU
WpGBUO6/r7NaKFrsckw+fbg215RHcM1PUBFzvnaVdkVzksy2J8Oi1Ad8LskrYPv7xf7/oJBawsRN
SJIfz+x0CXQOCqGlGD8FQgWJXsL22P8VsjBI3xyaTBI/Bl7AG1tFSX9J7s685Kn9xfXt2a8tl7A1
9zLil6+BuBZHvMWGWO+BoJplzNHB7kx8qjj2q069PgrSlnJ0cAub/tMbf3dV/L0k1K1LIEJ+GUT/
PTmMpDN6s2gLMtiQIuT5XmIVRM+GofAXIAKiJf46kK3KS1Iy/etNvAddbR4uRXlbzJPeKaQ36fMo
kC5ccEV3l77yaJS++mSIr3Io3OdY1yXcqp8LYcAexMGd+L38z3G/mNzskZe2QyDxn/jccl3nb1P+
r+fuIsRfmPHGina5bl3aLRygDsD+/LDCSZpmQ1lrBm5Mm5Rrh7yDLoBxnvuIVn+TDoGEQUaB74FV
sTuEL/A8YanCwlPUEFsY9JOK4Ou4v7D1qxhc4WiTW/0u33Ei5wJSojvkD62FIexQ5THSPxfwwmjQ
TOf+dMV0O7RjeDvMb7g1k8LOO9pmE/mi8sSGVLQnS3jxKj/ZUP4gYr89NNibyJTNxj4z+sHqhd97
gaPm/O4KgyBjV8vPsN8MQsDtWwhpuDE6ryVAtBrNMOPEp13NuaW5NhnZLaEvPRY+vjqwUlgVy/dM
Udma4WQ1Nkq7ZBs/FURKFqpmyK/kU17HB8qY/ubtCc1H4VPzwFtc30EgA3YetjpIllK5fYJPjTb+
WF2Xb1KYQGmusTCr5iyYZd+YFHWKdTJJx198KZPmDSMgKNayUsETTj6pup4waqqG43KQs/B9RD+S
ghtgUWMzvWVOmYf0SBZ0/YAI4lkLipkdwLT2YbkKyLfLxSt6dqwzdbom6OrRNlZQ73T/GxuPt++P
hvN1OgNWcNoeOJ3C5dQU/cYWy/2O3yrX4hPzkpAUZBhE9+bW6IC2uZYpE8p/vNo3sSrayQs5FBFn
fOT2/WGXO2CbxLIRdoTknp1eqSXrjksskYKetkNjH6KXtg9IwL8W3G0eL3Mv8XU2SKzEYKOpwJQn
2VNh0u8EJHLH17OyLrefPxMzh/hcjV465zz8xd95HEEzcebbDFzBYyFsGxISNOuAwSVbLLpDWQIo
wmBJEnDtI5yUvejU5whFCdwd6TEt1+uha0mfPo9UlvkUjoDpESoSC5FP1eXOKf6HTsSNbQpIBt76
RjvGrJVbge/f6ZJLEQ/YATYurjla6QGTOP/58LjMRQHa6UYDKNB6l8FyFdKEx6zq0LOK+r2ska0A
0yPlYSkf0qOK6LSFSfiRSLChyui5B5T9L/itO2CuCnxNsDX4Y0Tv9n7/yCEWmfonfuhn3huIbHnC
IoH9Uzk39+WsNAtKBI8+DDYwb/sNpdfaof1/pXgCAqM/zzaKU3lGa6ANEswu/pHuHpMyRL1Wzd6F
TejcF95pdc1EbJH8WaV0uS/TZSlX601dMGjpLlXTTF9f9cGZ118su5ES9UJaQA8EOWdDlTxM6lBs
Bpp4V674x4yeyZxuGkDTCZj1Z+dPPv7tbOWkS8qsA8W/lqBCd5Pye1Y4X7UU6CiBHdZ9KZkjarcH
UiBFtWo3ZKtNcUkKr5uwkgDxJXeQpbSfCXIXlw9vGdm0Cp6sOhU90UbCEpARawuEqagDFW4dB7SM
uZ5mNdVJe3l9pUgmr9AC0boxpfz6d7D8mFGI8OCpVoFcWYp82M5Qbfh1OEH04VtufaOlTj+Wev75
EcPW1ot0a5R+ekhDg6WM//WSwf1yh1M36iBoVrCPaSCuNMGykikpFGYKY1zzuY/VXQXHw8wIyZZN
S6ZkeE34AJvaguR7coPT6rnLTf728MzJkhG50x5G9cy66BQaOQdGWMP15/Yfw8mD6omLRIU=
`pragma protect end_protected
