// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VOS86Iz8zbJkbWq6Cxs+/b4MJD5o01PGhNANqnMroMA+AZhCOW6EpUm9FXG3YJ30
iWCfFjaWMRWiwfxMjLErp+CZpqaeh6dM7TlIp+Amq+81Aa1y10xdI2CWmYNldxdA
KHF27f2jkkFvoT69yQ2/SFK4U5qpQHOXuhhIXEBXLa0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20032)
0Nh309Be89bRCYhim/iP21Qr1m7/+Y69R5t48Bzi9MxjrI28EHn+f03dQsmARvUW
zKFJOw1f03wTSUWATy31fAx668PvAttVOe3y0Q40aistEFZPgn8EPPgoWwKbiaGf
L7qS83mPvFoCEKxVM3UlyDFHwofrNOMAEKb8qUe8KQW00hSGe2tyJcYhhv50FK2y
1H6BDCwigFY508r5CaUQtrCOPWmc9qX44PaL73BVPhU2r3cqL1K2Ndn8QCgJRllB
NpdZIboadI8n9tpPvtA5ZAbpOdkWemPAi3VyQSNFBBVXWfqL/JK3eG7Dmo2CvsZN
eh6vztNJ7ffpTk4KRUzWDPpa/kLW7+WNy2yd/st4eALsYxswti9dU0ZJXj3eGxn/
nV6hyDB2cR7C3qo/Zx7wQoIceQvrbA+WNqk8Z4OvmfRQSOp8iTc86OxTW1pxTBXz
6Yn18XL85pwg9MeFOAZhGNsWUMLTNanrBxOXpNw8U900j5LUr7uDBhC8UVZPTzTy
renvNHA38tYaTiF0awNIJyXFQS0aoLnBisyKPON3U60S0WxquBMuqsC8W79qESDM
kZRZWnUfgEzvRcKAqmBS4/PssshZL8H7IRVv8KLQDMKJtHHXJlhFqFFT89WdoB8J
7liH+EYVCZXRC6dJHuOR2i76mw+drZLylIEPeVM4OS0RkeGnPeoA6JnJZbMEaZM6
JFbLjWH4tAS4zpsE2+Jp+5Rz7lmQ4RmdpH0y6rI+dCm4QBmd8J4Pw382wiNUl/tx
8+KArjwbrj3iMw4vlnJwc79psuNNkdOcq/srR5pkDqF8O8hd4XqsUa6Unv0XOM9e
cFMwyxlTnyesPuoqnqvFUwxzEl+tzVz2u7ng3y/orw+L20DEs8+cdYH1UWUkWcpS
bAOHxmonsG5AHD6bqoj3fZMf1yH4fovXDywUY/lKsntvFeO0qw+Fa8PM8myYnauJ
8p3cAOUjiAMiFra3Gpkha8G+nY/9dOZjljROL+a3VS2VpwQj1kmh6+v8OihXM1mo
nJK/kT5QTNm+NcbzKFWbglF9i+zomdouyMYLK7xxVtpPlCaTZimW75k2GzUAs9rq
i6WEjRi9w6mth6snn6/SLj86THynKQ68EiDnFCs2c5eJb1+Zdo1MiMc1xRniN0DB
sBrBneYqYGugE10Nrxh3ouueozfT1VnLZRNAErmYBuVXlv7UBMHfqhqrSyhEiyxZ
NZ3OWu0AJSwlDElr8U+V+xEDa7ERqlf6XOKcfk6/Eo/1/DhBD+VZs6PvvElhM/ec
fxOSprrDTWRGWm9nPAIcyQkYaaEa4MRgNzZchcScTpJfBUGcUqEdYBH2gWmIBPnU
p/FYNK2anIEA4O5CCfOvOHHuv1BFuEcEuIRwCuJ/4bboDi6vh/pUTwLp5b4Fpo7i
zIHNifVeqq4+GYjwpnFIS3GAeCWDsMim+hhTIzmm+plNQJR1iUi2SY6MQ9gODLnJ
md+epfbUG4DaEvRHA/TTi5y+dL+EfX1WGrRX0r3qPWhTHV43bSJIpe90FPsBLj3Y
x78ctAPEMSOXVaK3FFmiB1GHvmm+Va2Yd0wGZZ9FPsysPL56iJm7IyRsYEycrw5u
Mdae0qyusnXurc2t6TKlstN0MSSbLScillvkuO79o4P19AMth6bDPIL+cGNkF8L5
ffYrciaHHp2x0PC9xMiaALbl9yNufxcxBD9abTIzBiUUeW/Vo7r1C0R1aWKpyk0B
sZXB+HOQPCjgeS+q+33K+XU5JNFHGXBiGo/UBIxaNgBhBz/vhVS7l255FqKjJGNF
H0OXfF1N0P9yTLDk/peEwwBblhlGg722vqZGv/UEcnMtMm+SP0talS/ag13e8hNa
tQM45rHU/rguCUq4Z+weOxdFXqfKHO1BVp1Uj6+M+K7NOLVclWFyk1WEJJNl4C59
ZIip3xHlnt+AfM90CcDdV7eDp2FnnhFiY4I4pp/KTXDPkwy+gAzKT9TISZo7POMx
p5yspj9lHoM2QxX5h9/gz8cTmAIb/z/AanyRMEb7FRwbWy77jyeCGDMLKxOr6deQ
ZpYdjRlaSdHFpAafavOIA6wYf2OAw07J9XoZ6NmjxTU1R1nBFeU6zSp4NW13i2xt
5CGyaf+XmD1pV0LOPWVbx4ThKJ0yvMp6pTQ67WEmcaL3hRxLOE3x14w7T3r6uOuu
3DUdBiq2iOAEyT5vjkhiM47/j/7QNAzSeNqBvq39Yd70Y7D3igfjwnh7HixcQSqZ
nc4omhqS0AEd1kx7YSy4nCgHOH1tUBByFglNMKdWPxh1Cp9snBXhq5ccFT8GkO1T
q0ooeiLJxUcyujAS14ARli0diXHHlNe/agHu7BFY8+5gC1xAQmXC/D/xUKCYUknv
K0ttBpd8A0njg5dI2DSGyhjRmNAWOUync6YKG0TqvJeQN0F95N706j0Ki+D4tKRH
1ArCI8kDE/Wg18waojl9g0pl34ssp7rMLH5Mm8SO9SzGNpW4xCbRrRowq//LMC0e
V6bjM056aueF/wDMli8QAscOkusWj7COk8QnXZ8O7VmkSA/ak813pSSU6/9FgUYm
QTVCesbockFqFOdEe8w85ZmxuPSGKacF7cT6RqsegzTKfhTe/rq9ijhI4zNyxeQI
J5wZIqwfReW75P+mb+DNJ7xzdd5mFIseJmkKuZePXa7efVu6eAlJbcvF+h01QAgA
vU4KW9MqYTXvpdXRu7SIvmAB4XDAZ1l4lQ6t/Woq+Y6s/tERSVy15fwy6+ypfpCP
fHH3j1vNIG8fiqy8xc5MnU+m3LdYduZWRZQe9IdxUBlcLyeN6tvTS5zM4b+GAzzY
WNNAAGRUixD01Azp9GpsA3PcKa0FOdCJ8zXbYF4DmAKMaHQ+ZHkkj5Wn1+SyL5Vq
4cE1k9yapuNREMzT3RCqSsD+4lS1Yhk22JGIA7ffKBmun7KV021N16qb8YcuCHn5
dJWXnQD/6il631G1EcH3M636SKd+F+TXbsAOWdL8sl2mB8svsnmpVec7mOxdwAQA
eDxVa9lmcxCKTVrQrKBxsKqsIB4R1zCPUO/A4juFJAJYaGjMJknuKIaRPZeY+C3Q
IQYKiKLwxYawOLcPxl3RIAAvi04Ick7OlR87gUdPMQWcj89ciYldUV+y/JxTT4jQ
T/kU+oTu7/aVoY3OjijS3hdWzIfm4GAI7ojY35RieBOf/NpKiQeJAgAPoPKqHQI4
ih9YW8LofgHxq8mK5NRnoERz/plGlzqKpd3Jsf+9YEOXFzPcq6oSQ2Fhq9FkDquH
V+eR0fHmyIivGZJGLSpmry+rfEEIqlGpOHsN/ZRWRLBFmpw1LMljD5TwaLa3kA+w
eKDRZdYr7rk8KWu+tvHpLM6qlPcjvOGf5kRseV3sbEGtzIcpalJkb/WO7IV11vcb
YqCmUK8WI7zj2DSB1+ObKoOb8bozQw6sWXxUFo/xoOAGWVpiKiaJ7fPubu9ADt7V
c08LdzcKIHBQV3toOZ6+M0vIIAD5z6XskfJRLAF8UpwR8l0LoPM/7P3srvMbWCUo
3cYaaJi4pOobQHPtW/1Zqrc7E0OZXDWXz7Mx3VuL1NyRceAt2MLPDOq9pFZygHrP
vSNAuRhu1WmYYDiPrfsrnmrK1SzT7W5earINdp6IXRVNYo0yN48vFyknlP4DZ6rX
5L4u2gkdca31Kr75MlwfTiZZSFviauv5rXuwFATHGphy7MjVk8WNeGY1rt3wI+8Q
l2Q5Xw1PqZg280ikysO6Fu5B8l+7PsujoCyCOOPj/VOTFEid+27MVxqPJbzMSH8+
dFeN3s5UCZJAlpj1iDKO+aKFafZ48kF3hW4pED1j8TJ9f8cInP9mt/aNe2NBw9F1
u3JJ+oZN51y5T2x6OnbPC4VLyEMBSomiQSLTfyxDCi8S+OPtSnv6AzO3qKi1zEn+
Dx0jhfr3/9dlZ6W2C9PfFxkFfVItA/RDteV7DsvQf7XtNSyeePnDurCXLUJSwdnx
LurYe++3r5Z+iqVKwXlaZ8eI2WAvXqjxRqggUJtrVoQmaAiAwomVuaG3ZQ2CS68u
JVEKTLdi+Yj49CSbMGkVCrnZaa+j5fqNtCBeUFuMScCSIxydY8JbgD2QGhmYy09J
L4KT/99Ip6m81/DJc5+KtvPiBYTxnTbm5ABXFSfLn4qu6WJmKGNITolAOLaHiOPY
OLInCWZMW8kKyMKb3UOiTivtWvnXA/+ucsLRXmsY6FPUAUIeSS5klGW7VqalPLb2
ZtqHozIsxxSY2y7DllvXTFGLli6mYo0ZS+kLAiDfnP7ZQUuGYzRjyWiRti3dxFG9
L3loRAT0XwlvQrGonIo8i840Lr48IYxMudNpQl7dtqaVPtc0HTYmnzw40L06czca
YNIgK21SdEFlf6i47PAAJIsafLjW4yRYfIqA0QFs2LFS/hiCNMeQoTxTDFCeFuAP
55uk+1vuhRI/R2uB2UTeBou2f4/3re6xoaNcVLCgcjkVJWqPZ9pDJ5ruZmN7EH2v
Ed6ENXD7Yy2MeB4jd+5izvUS8qcvjEV+NKz/4RdeP5kVCfd2uvPjMHJO12qFyTAj
1+Tf9B5oVNnmYuHGwiguKtdXei/7gXevm1C/xfHBEVTV3qPRAZOruyoJtQsgB88A
yfL+a2b3cxwVIGh2irkzci6ejECdgExxlZ0znFbpnH3eU4ljuuKj8yJyhjMR9U68
1DaL/u1bCcMcxn/++ldnG9MI9wtJs0qbfPrYUSalL1jf9exHOknpOlT85Qe+9IO0
zHNhDS+GH7tS3HPJfj9+CZ8CnEazzcefnYJVqYHYprcO9jfa7emqQAcOhjXs7no4
93jTOTxBbtVQJwg37Ivax/WnHHuvI0qmWo0JHY4KFs+BsVYe3nUTCyIN+F6XkwXL
YCowYHfQmBW20Vvz5m+CGLKckNgVwIIDbH3+oKP2h3+Agh4fc22Lc1znAjG0pNtq
yHEbr566eMs/1RR6WYuQMF6bF8ZpkYGA3RR+or9ev1zMqkJ3ZVe3005lVp8eoFB4
sMfT7diFHBHjAhR7zTYBfCuQLEFIOUo3/RyUMssEugDK9ct2efDpnHPynwnpuQWp
Wm0apoPelM4kx4u61TZsnrjMB54ISeZQzpMQ7GBCFBe/y0a0SmdzPNLIZoqFFcMX
qFvvJpwPkfD+NY64CIkEZrq8UDfAi6sLWZ+cP3ofRtM/nJyyGEUQGaS44HKa8frL
bFuQeAdzl3YExthpbc3jjTBpWh8Q4s/WqMqCyDc1XSdHgVcAupUgXoqEAF40EgA4
aXGyFksew7e7WWn20lJ+xE+8Uv/Nf8mMTkxpvH06ZFXK+15kzGUbs+vunNLTLA/W
I5rE2/xMIK/EGeOrRJEVmmcVlKnYovE+oEStU92gbAzMyvwLQOSCucJkehXPxIwU
RJtWqIuj2TuPU2o7ZjIVKivQEAa15m+C6jgU5RcyW+WGRG6iC+L/ht0ZjArDBnMV
zx57vedPCZb/NfeybQcFsLtouq0b5+yKJFywuKyn2eKAAJ9gSPsInxKxeafNSy0p
+1Pl4K5FVXR0aAR+ZeDDTu7Mi5A2xrqN7XE1xNfILCJXSBDwiyzYcsIi0x/EVkNY
UE89IfN1IMc77IvyA6mA6wVbJzF30Ushltdvt5Cz1EAi2DwLd4BDq3pqhWCppoVk
Tu2Dl119MqAb4WQz/X95qKmiHoDioz7h+C4sVPzebRX1D4lNiukcArFNQSEO/P9I
vKcUxELmD5g9tXRH+TKkcRei6kWZn0xWhHP+KcRkVDgFQNHyWjHlXsAFNUdN4knZ
x6wHNGdo+skgeSV2QCypvk1zqosPCmTBjrKFTyKzjCYvWnuFmbSfM7DG0pr3F8O5
r93PvOZhj9/UkeOrbRNW1Z8RyaY5F5vYOR77tlwC2MgZ8yEvRK9MgmjJsgIjbyPY
+9DFl7Aov6oJtJWL7ug4y80Y/2XBC02eAQEEnfn0Tnzvd55E8RplPdxC9uiJ3wsz
67iyJ9uGMa+apoi+OKxZddfZ49uqOy29eTxKZ/KCFnngNijjlpr4iqmZ14h3g6nF
e42nvZ1EOaABewjmv4gg2zJfjDdkRIbMtjTec9rxIM+GzMr7qqyz3pFoziXFJhIQ
nTERI/0XDdRhOPR2HBcVduOykRSEfGgMy4NVkRKZ7EesnFrsGYnpdAio8LWweKMW
2BoOJJ5JTe4hUjwIbuPSsQoBc4DxOBOvTj/MCieX6oCTdmXEckBwoQ3vf5L0u90H
5H58UDlUlJVKH1L3HUwTYRfCTDfWipdOUx66SvLnKv209mCPJ6ld6eVZK33+yJPN
qhZFYulI7fgawCR7KUjefTu0U0L5+vmW/kUgkdyAg8nE30dHqcdwOUrq6FcusM7V
XZiuir1U1vKlvsoHNmg5MR9KdSlx2y9Fq7kE4ovmwHn2LcsxlIRQlRlO5YvefYps
knpvGBxenpRv7efWNXNgh4J9t/MgahfAQdQLqYl+JKXeyTgwX6u2eYKhH6hz4l31
CX0UBTxiAThinrAu8OXFekFzgAiamYTQ6tlg+dfZKPvfTZzUK4UYId7Fyo3rEK4P
KL+X/WDbl0d4XlHhdi05ALAv7WpeOxHEkq4qVHHAgvw+5Sl5RMPrDu0hX7DCc7Xo
UZcTIp6cZDxMD/Vzrr395U2hVkIQPzu1Rsndh9BNEdmnYiWRiEe4URMG4o2u2G0n
H3DPedqZCaXHM+EYmbODDG/HqaarGpep1Buu6s7fm3358UDYGzLfxjZJ9m0TR3FQ
YgVE701809aOR09++pwLysMvxwbVMGB6qtuGkEtI4nUtM4+znz62qYTqLPOPYEMO
LsTJEXC3UAw5DfRRoPC8nkKDphLWX+FeCD5pqdEmpil1W1zLkyKAVbq4/HHD8v3+
ia72EjAQQXDNt349P1HivGAsljspA3klGJ8lImOZk2qdFUlNuywgmC430IAW+wkX
MGs+EibDch/wmJDkR66hJNAyQSWz/JtaVKsHnP0dGhnY0AP1veZkXx0gBpqoQ/UE
ercNZt/I9rte8HsA/DGdclLZ9/3iCSE13t1xxb4PICIbSCOYt3Hgtwyc4l3wQ3mc
AYqwRLjBgniyVYyB7HjKAGY/7VjEzHrrsT/PTwAJGfmp4lZiRX76vn0lL4cVcvBy
1P42QItrzb9JLOUM7DG39vezccr1J8+txKDcO5IV69fuvUntgMsml/0OJwVxITYE
5Sjvhsl7DwirQ62FT7YhY0q37S1DXjvkAt24DTVsvb+PTeLOYwwifjh97S12ful9
gaB1XoEFUQ1+BuMxBVDznPhzQLVQSs0u+E6a51EFfVX2Cne646IdMmDB2QoVoJZo
plZ5690byU7MB83qR9rv9n4WULHnFr8ajfnlRcpZnxErYYPMsL62ngMoRG2EQOX+
kAJAU2k+f4z+8VrfPpCI008xMDg3JbOlaN2qDs4Ffrl+F8oryMe4wiELO2GBQgnz
kgVpSuiHj0Zdt4DGzMX0c3Pdbr1x3WR9MX/fW3TA4iHCfC6idY2Wkl/0Q7ztjR4s
lI3tnu2hrq2A+c5C0m6vBZ3Tby7BGxuHV0kga1OIbqOv5w00ZNs2RNf8Nf0Q760b
uGdAV8cMqetDH/m1KQ7Z76XuEjrXWTSAApQbUIe9pC9XsI4QhSGtiZMvZgT/yNws
ZYaGQ3BLT6/hIA1C7Fn10vNJwXvTABfitba5I4W6k2yYEV9ohN29XoZ2Ydo9KMDN
q/0iyBdzTX2gdlnD+Nh+F/yi7Pn9erhKdbu6S9xhmMjiWnIR1ZYni8B/XeHjOwdG
PenR8nfx+r9uUwYy2xjYmP4YeN4fXkBlSTXXcYgyMFEjQqcMQopIo4e1KC4f9nBr
U+fyGGcaPjzxjf+iCcikjT1CI9W1wWn1vlorOTEX/UlR1HlJ2Jjb/RbloWvz7Iao
Que4H/gy1EqZR8UP4i3K9ovIAeFrGrvSBNxCC9GQk6xYRnevYITG7aZTRZQGWi/X
N6u65Zg2sAMk1f0FNcBonkg7xKx454xkjmjJJ2xzA1nP5HFXjlf8sRlt99gn6bqn
mVPJ3jvFOBjxvCtktRihYUNRVjwM/k4De2tC0UJgMgr/C/TE+au1f7sJjK17fjtE
ZxhE1LBuGdQ6i4jYV6EKuUIZe8YczBwppC/nxzyEAFHfNsYwXFkDrgWv2o7oazXU
hMwQLPuGLpf91z44CGnY77EJLP+EZgW1osPRE2ZlYR1KZQzdmgIoFcaLehIkWmPR
4n1c5/syJURz6KHTSuSBjzCMskD2leiSnEtG1rdIfH/nlTWsCw8Dtfc3U0367iSD
IATsSnYpxWB7y/Oaj75jVBSR2IjwOEsCWyhcqcrDroNbOv6Nk5WFwSgVz2/VR6CI
WR7f5cLbpuqVAxH6ZPT7zwDv9iCNKHlP8ZYDuwfTLxi9aGke4sDqwFOGW4AC23po
dMe3QXZlXGvI4D/qceylDb1VKqOHl10BjP71jy+G7d4xb7Jdp/j20KWNxSc8i3Ac
/vgHwF+RdAcQxbNpDK+WIGK/rlInEhAOEWcNGGt81++lWDaCnGoft1IlZtk5Sk2F
ThAXd9vnjliKof6vESu/gPynUGfeamGu5Od0DAF0immKKLIS7ZDEPNDxjiZcLj8D
1ujIpiO9jkSwDqe8LWg8K7e8b3ZThtQDKFQl0K9Zxz+SieIc2tWfXc4MnLZONyQF
o1Xo/+y7SV9YIGTrXLwZAH0YQQeBquO9Qelhm1VWLjloWvL+86ASdPt0XPyN8Kp9
UOOyePl2mlq+QYNO0CDIrB00W1dTVDNfwmIqAd28GPN2ibHcyeJwm0iKbQ7NZNjq
ScOowvnambNhAqNmHF7ikhBudmyoVs2u2ZgnUVhcp5qOmEbhULMB4vpDhg0nf7pD
8CVTMcsx8bF4tOHboMgZ4xO9m/nN0k26M/fbSbt0eCem1jqWwJ/IyRmRQbwVCD12
05vh/84emBcm2CdwaJeoplabj2A+4kjcM5JRTiCvGMRX6889Ewj7N0n2kHDnNP9I
wrYeSWQ9zZ2JMK1FJFzvG+we4aAvg14dnDdPFHQX/dCQqZNNwEMmZKH9eMlVQnm/
FRs8KuN89pulb2SgX+06BnOr0XDHZj9ReXZHh5nb7l/RqFRZMpX0GN9mb/ZFFIHi
pANxM0P/5H0A9SKjEHWdvWtY7uRfGGJw6iqOSGi6G/3PzVib4ULNA9SuVzQ/E6a6
/spYwlix0coW+JQAXIpm/+Uu5xfEjypmGCHkwTAXShJ73XmoVsqXKSP9qTdEH9Xu
2nCigOApZM67n6gKJbu7gWrtDP80ir7xMHzIOSR5wz+5/pkWMxCG5+6RcjJglJJs
wcGAHUmmTmQQOJapAKuOEacozv5H7hgcE9qgF3z0LNSUjXr0w9UX0Z3LibO8Rdde
96l4DodYV6pCgO5xP4Q+9O+DiUeJg1+SQ4+kPCQDZqRIiHmTrxlXARJaWZ2McBJU
CN2uDPmD8qag42eqz5v5h9H9Ge6mDc5C+vf5aimPFAzD3eeY/tjSr8uv65JpHgNe
2kD/EFypcBXEYZU0iB2XBmywzLRoXuJ0kMdcxqCgXD+GX4a4U+YsXvM+46FWuOA3
uHXRDoHLkHZ6cU3gkpUjPYNoaavX/s+DMQzYH39zvKQH91wGl6SEwqH+2tXuddOW
IFAjM2yeuybGScUGBgvSXwMHRiqUsAxePQQgrmvDvlx99GI7WlNRl10bvQbqtIvZ
ksVMVQ24CDz4hyC+zKl/zFq0C12wfjxpHnS0QIgc/2cAl1U+NsHBeJEW8b1KEkoA
6SzxdbFqOFGXK8ZBhMwYOG3X2gHSyaCGhDrbMQJo84SAPP6y4MinaAQyzUxRiLFQ
AR+k+QBaGTJIFmjImJOpC4oQl1JRn1w4DrlH5Kx4+AypUufHsBthilBvzfRVOIbP
Plt8Z1P/yFTPa/3R8WCXqDgrz4G9sr/3pWQTPy4qDcGzdV3dglE7rPJRgoKvFwDS
rqkq08m7cePT5Fb1myn/CLDJ9uGYi7T8ouCvCszgGxg19Prhl96+wz839k+ckutv
+XCxVwqpUBAVYZ7ILBHCLE+fMaibqxETl7Da6bbmSbfFEPG2p3tNJm+Q3paCrwZZ
GLZcgdDdw30gPscZ462AxjwvllBh17/F58Q/IrxxxxDIbaeFJGp5gEdyF0oRogi9
clGW4ky13y9dHbDh3HSrITCsnrU5ql4ICJuMCgfK9RWNF4eJeepifG35Y3uYZUXM
erthjgfsImb6hfOtLhHoudIaYyhv/DPBcqKSRq8Gc+svTG9KkERtdPEC3pRHlc+x
gzLSsZtD1phCEK7+bJ+Di4HklpkYHDK+PHixoER7lKcM0UVI5/01kUnVJkaJfhJK
38vx+bT8S1LXyMx4iY7ZqycMpR4Ri5l59LWpR4PHAYpG3Q/1PbvoD4maAbONHSFW
DrsOhj50OdeTFPznpG0+D25hnR8stP501Lzyn2RXQ0DAnfw3wTHKSk4jOBhzsgLG
tCtDYhhPp1eN5VTDLTDL1G7g7OLDBZZ87eFxwtGrTeNhHoBW6++UDC4AQWwKg41b
6ccatVzH7s5r7VPHkM2ADcZU+i/5D1HQkLqAiSrRH08Ql21zNBQvBdMF3bClNPkz
wc2gtdVFkHPGbXuGMy08AqS0LGksfDASrtYJ0xDVM23lkC8nBO7f88L2mzZQqZzF
Z9U14IoTYZpNMt/xjPkU971gOpG28rioSf10siTwgFNdS8GPA6pKIPxSZETy8ZLE
EDZRp02htdCHe4EjInOoFHivodO3Yafj0au5vT1HaBHVjJplDpPjz36U1zVYS5sQ
ugRnNZ0UUlmtmAIsoNUi7mLFzQeuWcYzUk25uK/BJvgYgIZUdzPfhjkyvUjTPopT
OwkAHiEx08sF8ODVQaW+nWB1XBlno1BPL5zS3AgeMbdLAlWz7MzZbRBZPVXS7Xe0
ABXXU9YHYrc6vjSCCn5779kOEWVnOiUTaMegUkIeb1DXipAkf8Pan8M9AhRHTb9w
YU/jfkQw+hdzk3Hquk0yanddJ0uN7wkZ5sMSyI40ml+26dyjNuiYmBBRFVppOaxu
n32DVR6p9lgabJD5KWhudIHyWrcB7KuPoh7PguLzK98gl+lr48iBePiD0nDUvDUB
WKmp9t+3WCrYSUKFVtEke9keK6i1reJ/l8Y+d4hqqL0C3A+mampRH7+sraROWRJy
XJynEDr2PiPqIrpXiy7WhyU3s4XR2lDzw2cIjK6Q5RzRGaxs+InQHZjEYfdsceen
LMK51JRpy3cHpaEiRIG1oj/+/2P5aKdfkD1A5pQcoIhCHMuLw9ycJr3dhkQpncT+
n7e9cdYazWAks1Wad4cxC/v/B8a2dsT6beYhJBGpvg+SyeZp8atOMicgV09f0FP0
JDh5nleKsXMDP01xqaTKOei3Ns8nX309BWonHTfg+ukgrKIv0MphXIAAgENAqi+9
JXPzigmOGuWJR/4cmc4VZ9FtC43hHCQ6OV9D2O3Qnii/ja4jNpg7EfNYGwM/6LGA
w36gwManh72BlJaCSLFXUHPsHZqhHUfbz6FM7DbpFb4MD6jbAlE9JPQZpDtiZQai
lD9h2aa7XSBiiiIxHV7vOKlmMwgmgEGQzeHsfxwoGj7LFhFIdNbSX3rnWGCuIeas
LXmBvffSE0JK69TtCgZ0GqB3B44zyYHBtkWH59A5yBJ8kR2tg4YyaJAht5PljP1D
1V2u50PHRtdh1bKIonXkeTXHsEMUJ6P0E9xMSqAWTDhFwfMJEdynoTqochNEbDm0
jCFX7mYfWcNbz4z4zR8qNA2sUrsu43S+D7yGIAAMDGJmJgSBlTu/NeHbNBnexo/g
xDBi/KzD26lCJ6uDF3xI7E78oSH1XNw4IKE8ovERgaD52U6EuWYPBAS14HtdQtR3
4FyB/y1qii/VrdU6n4/0xDS3oDohIIPSujxKnHXgAM4tmlavIIbGXcV8dGrqlPt7
JFGkqd8aV+Nx2yNogyr96m9MpcT3b6ZpUHV14H/EL63KJXZIbtuRa7CYJj5A/eGn
niEEPKwr6DR97sEDqFnHY5vsD8jV8B80UeXhZfo0D3kHX2N+9TCvrSJBuCVjcH+c
Tlq/3VYRAE/AfDkbSFI2XOSvy2laEJRvi8NsmtU7SwLVx3gMrNQCbGas8jVpcE9H
1yPM4cfpt+ZVmYs4Js5n4hPchzIX5j/FS5ioRj7moNFNvQoZVlQspTCshy3sHxwT
Z3BJjTE0Y1SU7x93NvpdLc6pqr9RcolYBt4blxU4PWuE1l5F9PvypT5YFKXm2IaF
J1Ln3kfzFMzicEVI95RjrSCuLk3RL0t63QBnNkAskubE51TvYIFTolqinA5G+mHz
x+tAoKrp5CjvRGMW3MNV4LDGA5GMMVTyhYzOJsz83YUAMroIbb1QDpYZDF3oVkRn
UhHQsjPQ0jZFjR1jAzR9mpLmRdz3Nea6lZpFPVLZ11ye73W5PUoGK2acsGlQ95iv
su35q9lTFDT1ESBuIJZppvt4FwdeA9QDxxUJM1c0UFd73XsiZ+mHFSWjRGI77uCU
I1K4lNWVnr9HQbngk7GamPo6GttGQU7+fHlxmmSL2puiSdrJ5DtVECXGCAq9Cn2o
/49XJeRr9iuerLykiBCZs02k+AbrfstZPnI8r28EiWOXlN9JcPl5CMNoWdihJvVO
C2naKiev80XRDfCIiYmi++k3vAckXr52/x7tZjo+bd8uAF44hy/CFrzvf6uubjJI
8wQFk++eizlseoaEbipi/OfVMEb19MDuioiRb8Rr8ZZlqWZ5r1Vk3cTIIz4T+E8b
OTfogzWNHisp/QlN+VRnGFIDD4c+GGyh19tZU1p5+kaicrdD4M8tOOzgIeIbTrHG
RjbMCHCXX1HxGlsCi34Px2WGZAmxoPwQ1eUB9MeC/p6KLp53+FuZ4DR88BKG3zmm
3z2Df/rrBlXnAoivqlj3yQbcMOLixnp5mZLX+EmxW9h7I1KfwtHWC+FlCVqRf0p/
TRf2EbDQNJi720GzmFeNgwb8XNNKmrDAi/5vfpRc3b+RxhK/Y5PJ/BHjZf10HDiV
LonNWzTeC3a4ZFrJkK+j/1AgP7tLQ43MF6NypcObmpwHiRI3rgJHF1MVyVYy0J3H
1u1bB7VLR2OQqE60Ilup6V1yur8nDg85KTIxtPOGLKlLYXr7f/Ag2i8Uo2tJbt01
Iy6fYbk6iXzX3LqlqUPBtYN+/INyRz8kNqVIFSY+e/tWc8FxNGzPD6PJJSKV18XH
qNqZ8a8LCo7JfNmtbwEqXagtRiEg7r24B7f6dF/x/8Jdi2LQ+R++vQQYUytq85eN
4BMnMJfDn8+FZvEyXuPXV/B4wVcG3XgoUGr/lveZ/ZN5aRMUTrinhiDZAF+5WBMq
WWfD8fRiatIitXH3vShjfwlQQ2QPYEKm1e7dXvwqf9Qes1UEWd112ZH8zvEbGK4x
MhsSMcp79eTUrMJYuxqJjb/GGaaBgvxtM3HhMe1r23Q36LS1KICwzc5QXTjeLJ8s
w0XAC3bf8vhLvlhass7VW19NoHoVTy5HF9HDi+LRm9ufqwGEoZOXw7c4rkTC1Enc
5QL1PjaHk74K4Q6ve78A5EdTPgtMgeDQpOeXrlEEtSp0sCYrDuCnrd65JJcrqVt1
vvFQ39Ysfy3610eAWNsrg/hPh2UmGhT7woJ5HSJxy5FGEeSqQ4se60K6EGgDv5SA
DAWcYbdR6a97y1T4lUOp22mLt+XtdaZRMlcp6t7G/S07uovksi6bx9/sCAVz1/Oi
kO1IH8zI3JYpYQxq1LLCsJ2g+4QinoxRtWEJL5IA+x0eMqmbVaxD3cGM75n8Obi3
QG0DfkLwLiZru9LLWd+ZW2nNLsrpbOJ0P0n884e5hK8d3ITa0XI3Qhwm866LhZa0
VbSYMVTfqrGQ7dqb3vRCT3g0oeRz0xBdE+8WQtSVciWUYa/8cL70JIKhWgWPKFlq
hft3bOy8K5p8XRfKkZAlV+nzP5grajDZxqgJ4nxlE+mJYfdm4l/r/3ZnjA2YWIUi
f6NelEAeUcPbk98qXEa9BHKZ9ykcY1eCqcagyLp/XtWIKZwml4lfnjXil9cv1OvY
si6HClLT58orw9n8cRE7VOSKstMLNt8+ZMwigKMralP2eW5JGRDrdi6oHhyrPxRo
DlITDgJoyEWGwiPnUZwVR/j9fVmB6XgSa7uHgbf/8chBIyXUt1zMPgzJZe7uf21t
AW+bgDKnylIPo5AtrhxcZwWjhdeLHK/AoxxzA31XZcyrwSsCUU4w4IAG7zKD40rQ
0ECwx+/AIcLZidmJNR6YGWSmmdoq8WCaC1bEEm8X8KZrKwDLT6acDBrNEDpjWzAk
pxxoDeboHRXoZZoss89m1O7Sp1TIEwgknMecM5XdB7iEEv56LDtJ3nhpP2s1AawC
wVOap+g8psBW4+y8y9NuJE24WmM56QEf/W3Gy6yGnZ2IyW8I6Sn9/9pj7CpdsZHZ
+ZA7KypX0aMvv/cJ/cRRwUgXhvGl0M6OyoKVSvHIGH5IftSztncctXS0rcEgZcRN
dYuqk2zaXYbusSLAkMAkKtv5OEFgv9W84aC6cKPschsSLnPk7CIfL11WfOxFiyG0
lhb0M4SE27XR4Of+71NiTWB4xu1cEApvLpMVjLgIx7S8xYgmt1EScLLyNC0wxrk/
jBhf9U6EHdJ/uBw0KxEHPGrvQ3RE9p0TMeO8CHAyQQ8OQvhhbh7yc5jwlixi4+jo
1TSToOTbLZrPzzUGE9MiuGNgldCx9xDS7KozAYD5dnWbMtiAMn1k8C51vq51xxb0
2ZJnKeM8MBS8e3pQ16l2fhBs1mwI3DuGLwa/GvQzs9QMKrGgxN0AksXeJ4EN8YbR
UNw2/toH+UaSLXRFsqVSrOV/n3Pzdiyfx+9Z+7lplpGfKxyGXvVSaWWwXJF4w0w0
RnSFEvxj9KHQuVWtwq4dJhQgFUY71Sg6XqEZuN80kpBb2lSPKm3f43QvyOHT5ARe
qpcz61QkmUuch01SRFmUvcbmDceP4DkulEn5AYIiOlZ5IjSXoycioGXbOx44jfkW
VtcpUwrHR1oVzO4+fmBuWt6UjzxbJzmVMSyYbuWNDEf6T9rlWTfbH33Jnd1MiDGj
kNguRPBGZYgLCB/Df7boU/deEuDEm2PUptIs7UpCXcgnjehiN707Zk/c2zzgdyRC
IdAYsJBBQDBp+hR7LIqdECYDklsM+klvBKjbT9jVvpuE4+wMV+E0PgimH3muD1+i
hMUsyBlYq7N80K/nLPk0uZGCfYkMN2xnZ5RJ6jTytiq6/Oc0kcLABFlohX4NHs0f
ME2RP2fWe70e9smvn2cNv3yYCFz58KWEbFVwhrHRKqmBYf9s+GGixFPlAYWDPLGq
CvVJPApsMlQzL4X2MGciS6LgvqlHMo0kMZNu0YH6utrLGw0NRcD2uS9S7DocqkYt
s3xOInyh1yvCEaHkyBVmUWMZ/6EsliNGokXYeF0qN9ia0mgjywz4Y9A98SBbKqpF
RuKHvriYLrf3FSZuE7dx45Se/aKZmWN/Ut3up2eojbjB4sdyVvyfG+nhYk9qYDGt
DNAmrZtPXxTkAnXTCj2Sm4LTONbK5WlVctoIifRdbikrPoIM2dgrd0xITDv6xxTt
+xiG38RWnrKqsNvrZSZoBIhoFOo1bQLeBodXeucO2px13wNX4T4Tf6/Kf+hI584L
cyFMVUDvAd9pW1qNtXf9jlAaopnjOv2xfEcYBfgkvsu0Z2wjXbJtm4RUDES43Ely
meMm90OxvmnW+Fp7jCpCujqAuGlJEbDlWZgDaQb8wnTxytSWaO17M3TtcyTiMENu
rD+tJFQuSIkMLWyE6F2nuJncJZ/3IaP8VamVx6PmySoomUoUmpxAOYnf1D0Z5PyV
31BCQ0DJmSXhXLxzGFXqoeXciBPiwrWDjVtdqJguujnHs9nnCm73CrIu+uNIxBrb
WQmRkrpTGpt0DQbtYZ5pKptAcuAmsklV4FlFXZ6XHB/9vLI005n9K/Wh1f1NS4iG
X1Fm/d79Zt+SHtYq0/eJh5kk6Op6BIdPrPFAwgKayC3jrSjRLzCMzcZiOSZ8fxKI
CAPb1hcdo1ZYtAkOajKjGPcqsmzfFFa55Fnu14CjdQ6Ky5CcZxvh9EZXeONdF0bv
VU7/M7DKE5hUqdjH2MzJyt3Z1tjUXv4MoB+Lu4SAQC196/+4hhYBvsYlCzDAXWe4
aGbcZ/LN180DmhjcbQGndHvCUvdxrb9xhkooVV6n1fS34/GPI/DU04ikRcII6diG
J3PAvT7OFh7AIyfKTEIoXgYVET/FhWZm2t2ObJn3IbUKuPX6AUy38VTt5xBaJmlF
kEAHkMkAoW9S726VMsWeE+o+thWZHmbRzgmKmSIiQf9X/oV6vB7Jy/lB5qxzo1tz
LMaSP8tMXlvGxWJmwJB0P2tYW7iAMzNn6KLcEpcxIOPYiW4Uw+RGU33Y2EVioh7V
omfto8ne3VzR+GM4tuO8KPVRLdC+xbfulgN9BoG4g39qENS+0E9kwbIOdvdWe8AZ
eQfTZAwGy5UCnpjR/Xq62C3ZhGMHGZjaTHLM5/9esQxtxBpyPXpvAboWMWMTfN+8
/uPRKDF0cc4TWN8BAw4iwXpzFNYp7d+PcyCfAcHPQk5i0zufCz3sMf4GUYUXybNf
IW+6EFSjZQC/Lwsb1ScrkJb3aEFG9PT03qvVBQ/Ee/iH4a1bwH70S9e6BD9iYuZI
duJRrn5ukVHq4QEsbGceW9tOUXeYT94cUCJdtwVWb4fuj6LjurApius7WdO/QBDq
EpCEQa/vq/r+WQM8ZKqxJUrAEjXUONx58VBo9tAqUZKgWUWVQZu4OjXlH2FviaJv
8TR6epFJ88j2uD6ZKe8vc6PTzvbZS+kjpwNbZ7U4pMkKim1a03maMJDi/m/7WwQY
3mghLxEX0evJSImP5fKZmZyePuQwzSeypTbwKBO9pXzByy9iqcrMqMIFoeY6A+t9
KcjPZkkNhmotyF5FgVKSFYTtklUD70GIBnQogwwkiSHGIFeLOz4crQQosSFXb5yM
SnOyeFChLYAwGFh72B+ZcmO7Q37W6rtjZbAtyCFQ7PrOminQYXDvu2r0hxlG4nVX
ky0c/UMx26wTWafx/sGs00flxoPn7AAjVoeSjw3E+qvk/aC1bkDYXpQGwCcFVTqs
rDEd5LOu50uTCrto9jQ0kP/hgQYkw/vD9AZr966EF7qvC0SKce1keKwZvq8F4c4+
EbYU7wVnnebc1JMTLAy744vBQWGT8L7GEmm1ctoZhbVQUgeytxOHzfp9KIm6I0f6
n+UShrOnAPCQKP+2OevlqvDoutP0bFbYyNTFYWviFKVBf2XX6H2LlQn9emNJ28pR
B3DXF5PMsnBrTCD3f8gKmU9od6jpQSveHZG+FmrfgiG0wox3Ter85uVFeErpnEpp
P4577jez3pvEQm2N1aYMit/bemT0KnYzJFp3rmE48vuy6JeofeMqw+FO7GFsOAGL
QvmwO3wdmwqbnaJWSiKMMwrD7FTe94Q08Ka8qjL/O5fUpnYZqJ63I5vibns8Cgav
jlDwqRuiHZT33XOeZ7Spwef01APkR4YUEsi1LOu/Eijeg4uHGb4dnjnyeIaPizDu
74YmU0tqXAta4X1KkwJuAL+yLv9iZu/1MhoEV1BQt7gddYe9x/ri9GyYt5ANJc2R
mSKlXiP5bbpwV/eAQOyiVJp6R2i6rXNUdem9Bx8g+haEfcJjBLmgnATJnagL2pU8
jxFWbJYnhGuTUvpuzHjaKOHff30gYsbauA3aX+bmEfYKojixbjJd0omsGXZctpk2
SIsue/odk1GIOwnI/AGN1OfE05C1WriV+zmsO6vntdUWAL1nP8NY1Aehs2c5Pu0/
iEfM0rsy52TfK97uvTWvGhCknP+TqZuVC7ExKQFs/xRLbRf+9SsiPR2myWI/iG6t
D9SQQfEPI6WefjyrxN/8YAYtJ72eVMwDnjTqomtYT3dcXr3+7oFzfUzXxBrSA9xS
bRekHTdr8S2J+5EzQAUqVPgthuvFSTgoXgu1IoNL4ifBMlZ6leJIUeArmyW8gqtc
edYCetJyjt8MsvODVeaUKXL5P40fvtf0e5EgN5+/QRIXSdeIGPs0io7EblUXZFjL
Oda0CPPWw5knYJM0Uxz5sq0O2s1ZoHUYmEbIYxn+a5f13UrJZDgfvU4BPeq/NuhJ
7IZylOFBMih6NGeYwU7Vq/Bv3E3rYy5EnNbyg6ajz1T8y/dvB98J104kNQyg8L2C
0wibnATLNfMgPfllRX6mi+onXklfF0N33akNpeeHO6ttaveLV7K0yTy3dI0OcJNq
hNcydNun/MuNPiFH67m9kCwAOzHpJYuIxdjCB/GEjp2V5YFyAgpB4n3pLLFARbdH
GUP619mxgr8nu291tbUsyVvz8gXVmPiX3VzNxw8tNTQBeMvg4Jo1mZlecRU/NFwE
ajOPqhF5iIbOF1LDEloo57RCmhwZsj6RsboE4zM7yebDU+TDTJAaeDa/HJ3M3Rqw
R+nCsBWHnbLJPdDq0J4p7dabYzwG0hLwL3IeUA5I2cnTaHV1UfQlN/X50VFAUm7u
4qM4z+d788Fy1ipFOjRKWN3MEQexesCunAkfEYosx4f4R7PapcOAk0NyMN2eXROo
oSFN9655Dec8YMkJkjfNpoZjohDWCnRWAL1SyBQdflxUOzWGqOs4CNzkGsfkkcjU
AYmfUvSwB9HqmFz4ajwc4DhLQDJlJ5So/guIDLC3BVGEy8xH/IG8ffjtcRS24M+L
XvQdAg+NPktPxcT73GDsLfCrsju/6KLyS82qc/BrJ1TGkyQQVVojgMd/9M1X9jPo
qWlXkjl9SmHcrdQ+tUUkgiWXAygrVBfwSM/9MymN6pcAdFYvbBt7B0geiK+RzEXS
K09yX9tPDdgX4/vnh3HLyxaoi3h3PnEUG4CyWT92FYA6dARavwIJ0tH/z5RheFg+
+t9jA1PViOx6eXkz0kMxxqZ2n+j8FWL46VkqxE7NYbhmLm9Yuev+JcYZR1jh0y5v
z3DFHlvRbOXVCSWtRHzTU7dHXcI5zNdtD6Jdo51RjJSxE0t6AFq8RdhN8MF1sWPz
uTVABDfRvHXign6CnowL1Mo6w+NF4An3KNII11Ay/SLCNiAqJaE+yaTbGUZLaUK4
qZLa6J5h9tSjcjybztzw6Y4mo/tYJndbdLC4Cg4rG+M77gPyhob1+IJNdWMBtap+
bWtVsCERKajlJrNvK5DTorL5dz8HLODCLaUKl4pplWH4dpaGp72L+Ae4TIFDpiIc
rZpLpje7d9XodRASubdEfZ8QPiMYMmSAwvwmWzKC/yhjN5jX8jrcitd+L9zP26hT
s+LJt+52KOwpUcXypZ7m0DFqy1JJGD8HS7lhMpDmlOCjgdAdd4I7X+7uE0egDftr
YJjEVurREKw6eRLYpFZWdmk+uBX69CihrGeMMfsg1MqK6j262qZpPpA5cWAG4cHi
UEX8gwHTgoAX8sBzlIqmP+OhqvwDlumFamUd5FVVlZT9CEvWzFYUW44N+BjA0hEM
ZUkn2KPf7tgTXSA24uZPZsRQEEXAem9T3AdEdR1b3mLOfQZmAWpkeaxiWiTJ4zcP
U8w81xwyai4lPY3frjuMs5YOdXzNmHHmMNbRO0kv4J1axCo+S8fvHDojLjq8XmNv
bedRmlDXsmsgX24Vzbx7qAg3CFa8KFjEvu394i9U9tzryfjPlkMoWOv/YnAVBl86
3iOqEFteQXdwCD8lV+6ZQxRhdw4pa93arG4RuG6/4wUqnt17sjvUWEJOJKWvYRO8
aHxk+8TqkjSktx3K+pnAQCb92394owiVdJXJe9eO8PtgA02NaU1tWJZvCOCMPkz7
2DlpnE+X0oi7EjBvtdw2Qua+v37PmMuuHwNEhqqEEpvU8HZu+COLXGVjs7PQ3NTZ
+i8DqRo7WHbCOb8WIOhYWGoH6qiXue8rFCotMjBmyBoGb/2lfaq282s5qCriZ+U2
x4M37e245A6s4ztzCmY5a4b8XCVBVYoOpqBN6J2M7ReTqRmTUYsBs7XdFkPZaZUP
Oac0lYOjAOOEGdNoA/AU4/KmKKZWSOnQwS5iLCpLWR9c8Z9aJ5JlSO7EpztQIbhp
w9yUu4HRwmcnqAXlvvv00XdYTl6IeWVzCxBIkHnjmWIfmU0U9AFXK7tifvj6d8Jr
BP7zK9A8PkKYeTaxaIFI5CeqjpbY7nTefVxPh+ZfWmj5Hlg9Zw/leZf7UqdPWFmD
O+hBKO9NqSy09zMQxOfsF5D5E04cl6RtYQ93zuEe5WT47KtdhSEMywzwALFvKX4Y
2jRX9tNL61LzL92B5dy9UMGjchU4rxHzhKztsrFw+ScL7CKB5AyyoJ5AuJRaPMCE
nFK4sjHhR7IGKiguKtXzhw6n3bPT7Hn4MK4c9lDHsBHCFosW5Ap1+Q0JuJ5fFJTc
9Epwj4EyuyjcdakjMzTvcxNiqbYGYRriMn/YcYoHMNus5E5IBd5DeHf2E3NF0HrD
wbY1qdlj11umubLDOxJmJY2bwi5oci1mt1kuk7ngvQmDLLd+WUXst1DWEYuquacI
rsa9HWWehPmdmHCNzcp6a4AS0v72gvdEEJyN8p1tjQ2jIpZ3qCqfszjTLUlDSM4N
BOQjZc535R3R+Z1hZradNTmFIXw9jame5m3+fmZnQH7iUoYixaBco/Bo5LTdRKQq
Vy6lN8FVjt3wcSVcTV0OBEVt5tuxVtKG0BHli806OHg9I25cRBVoxlyLYc8MWRZf
6P5PdkTc7+MLLqvGUpKOZjAL/4kPRZfaixgJWCV64xUHhW1eKNxQCq42Oh2Vmlyb
RlV0+5xIUlaxEECP/yotANYQWrq8XtnvorbmC1Dgf6CvujW1Cb3sufJjKxG8xFBe
G7kKSiHm+8ertVXHfGi5BtmHMVZQnmHRvKE6JAPZbAuwBx+jRtH/6D1EFPn8x8vA
XCIDxdmR8goNpVIN0mA/GrJLU4WUolqeNPivbfpo1mdLUtOAD7VhL8BEYCCuEAZc
XFpR1n7ZfBPJ0+mENIvPLUso8bP2vdFq0+QRD4pDuEilocoLiSaZT1rVYA229iNI
adfMmVeg9fpIAJLoj3ZCVd397Bn+oeZp9OvnGBexl0+gjK/8o5mYfOodv1u23sX+
fnTo/wE4Oz8blVX3o6vfETpy+YhJIpbvqppsVi41mdwBegNXvjFm2faSsth7bpwU
jUnhBUGuzaYIJ6gve4FcguGMRgtR8asHn/9yph5dhMcPDEPaCjdDp2C9Btw3SqU5
mLfkOEZGbjor+NJ4UxyR0xpH1a1O75j/IkK+Ecvpg8A5XfNSxrOTHTVPz9GN5RPp
ZEaNZPftXQ1vzd33zvczBjHKPHDw6kuetVabRbqi2RipBK04H8PofoFU98sL+SCm
PLEJfnc4cYbAIPPKt1+QAHNAbKA+L6KDSEnMM0mcviYdOjofEpQIV7+Z9/+PSlhu
XRG06XKJTgvcqNj2v8sqAXltR7GBpMM5xwF8HT7elgolXPw9vI3l3p4lIur8fvtU
WQ8uC1H5yE/nse7cIRmoJJ4Is0dbFIWPvS0vEuVxbO4TAbd3s73KpiLnGOt2xmCM
dVJpiUPVkjfUTbPMgnuovlbeVUqYsWjXu+aTsDJMVqZqnbxr9JvKDDjLwgynOPOZ
7gLuuNGOK7v4JWlLwDfmOWahCwF8c7SXuJEnQcBXRi4VM8j4mfUcfYSJ3P+t9rUJ
uCmIP/8tbAJnlc9fQwlpv+p4NEXOQ/y9kFDizyTOwE0y1NtivoJgdC1HRLpZMf+O
ZGYJVZtzdRdXGF1K38nrdM2hUGpEPjajFXvvKHi0OWrimRZSJIDkdNULbLP7zLCr
WPyZs8MmBe0riqKKnJxZRlCYkw5NA1XKntDPxItbciAN9xLdOuxbgumhI36GVy6u
I+GOPINug2svh762Gr6ZHoGVoJCMNosz7E01NpfLOw2e0r2Cx2TQkxq5SAhXui0F
NQ/h5tSg9HnbQ6q48I9s4h/vjFyXQtKCEvr57gA8tl5jcXCn1rclcwCqcYnLCfjA
DsxominZtqCf3ZKPMwnRm8N252/QLiaQ/LPWGwq6Z8A5BCe3DIb+7Cj+vVbjBrZI
yvbwHiD3ZxgM5ozve0xpckRvKjlHpF4m7lEy9KLmILgCF0sKogzZr8EySQveUrrH
mmrrUcUqOKD3MizjP2lfZPSUOi64A8MNMqJ/DsSjOub8siOO0UuVAIT3m7H2fJtU
1LGckSzEm+kv54YQL4Qxoegu9kpoNEGeNvDSleomLMR0xvmcBRgCEybGvghJr71c
xJBJ8ymmU96+trkfGGmhV8JL5V8yePdAGx2/LBkbuX3yBjCFL7I6Fr0sIQVRAC8v
lemM1mMBvN9jfszBITgohPaCOYSP8BqldNoKogsY+qA6L8LNJV+/SfpJmqQVBFOR
4f5pVdFlZsB4/ADa/x121IshdGsQBhyeI9cYLA1p5vCFHHUcZy8c4K0pLeklikxZ
8ZmB0UMx4Fd28O/CnPlaW8/7VY3rt+LQqghtyCMfBJ1Kh6kR9q36ZvYyUFDe5K7Y
Jchmp3yIe4z1kXJySDGvAeYEqfDiWwhKjEF+tYJeXZ9x5qS9OGjmNjUNn/W1Qswr
idIn3cb5XUAVjUk8v7zotRuRJ2viibNlONZz71/E4nH0Pl7M/xgctkOT0ekIEHO1
o19dqp+VgqyLZZ989xeO/8eG/9U7wRRhXNULu7YnyfxnyoCHXBVeKZWO0I/X4V81
pmfmLiyZC7cj+U3BD+rYmtcEBzz6DGRmJMFCzXf9SQU8inM/xh1jRAy0CZm6grOy
duv/tlkZXoWrafuiiJeuXnoWnoRhhz6HPFhUJJejEC4mB8HtpCdS8WGwvbyIlGtd
/zrukBsYnKCS+CCfQh3zCwBeDQRL9chYOlEbMvl4oBqwd14u72vPsvljpVhVTTdL
JgTvZqgNue9lHspZqMgLwQRiTOv8bs/VKzlvi2RPr4JixvJoqZg0CwqQ6WO6RrdS
EmRkAmZ2sSt3tLYg0hGJEvWzVOLh9KA0chpef0TouoGEUxNIntMH+hkNzVYpRL2G
aysmK+YMLF/brch9og6AzVosLc/QBM4V7bn9rt0dKtMheFeLYMHuwzl5uXF8d39r
fKqscwo/LqFluouW9s+hZ54xa5pfkFhG7Llo/Ad9j5sAoi0PRx43DJl7klZ2ZZJS
uWNDqQXbb9aiQQGXqnA0A5L0F9EAeDzZbGAGUMZdTQNCSwtGya0gviTm1cvtmAUv
xbmahg8YwVw8hfXKoFWKZcBjATUeYRLQwlW3gZkHvE2Mm4WAwJ+a6I1VQfC4FobO
PccIXmtEMAOtwL6O/gtWdiuE2d7ZbQn2hfXhRevK/gCSIfi17knPLclMgEfjlkkB
aglmCkVXT4NS2MaagOUEXBbI4uhkbWnYskZsxaoOUvmeOoH2HdVPn7ZpkFVL6RJZ
zhsaRJgufrSBPA5xpNdVUWDz7rLYjMD3y/bw/ugd4zBqFUTwNvAPkxTdlrWoEf2f
WY1NPM7ZoonWxMdH3xSxTh9ffhCyMAoITAe80VlZgwxD2kWvidneMdEHDwo1FsVq
r1K3A4WbGfSnSKiBLavxZ6oOUurQ4QUg/72Dr/10u2AUYHmykxvku2sPWrKwDsqh
95UsGdRFgx1p6gddoYdmJ80tvRtmnPyj8cxJ4MaoYvJV08eI2WK0YcQtvrMPHoEE
FAA/tGoNdimlv4TjzKG0CH2sa2wSdoO685EQhPfp2WlVuneI4woTjY4u6ndAq/b4
HYy8k/KaXfZhiWDhydLczBE7DrTAK657aaJqaI8AoNK1KpsPlM5w95X7p+OYgEax
aCOhojpvVxAo0aNklfVq0WlMGhQMpq1NYwMj79/otxy1LIShoEQaXMkslQSfMfJd
daYanEFS4Zd+496JUv6BPtXWmVIfFlpNVxGcw4007W0Mx0FNe6XJJszyiu+Bkl+b
d6nEYIUe4lZR4wRA85+vZkin+8fAq4AWbd/MsDSkb062zE1YO3KJaV++OLRrv82T
naW9UDJOudDGOkOUnIoD9WsZkYmW3uhfw1ylL6Qvv4mmdBoXREWIaqufv6+YLrjR
0Ax4kgllO8AELdJR9SVb/mWCqtQhoTu/tmPExuLZjcI6QsUvgbByQ7smZhie3YvT
GoR6WqeAVrxUnyNMnromlDhZg4MSTIsc7WDwL9h/GLWkW2Fqvp3+RiBx962mpKsY
oQtywoFpLQNFf0m/d7FlmfurBPZgpPQeNSEgj2cJ1VDudHe5gEqww61QDqGrCphv
XQmNg0n4Sryo68ZjSNQxYjFbk5o0NPCv05YNA+XbgzOZtZTe0sRd3zg7weIscHGJ
t/K5csMDEhC4Ff2FYb9iytLBHyC1PZBl3VARvhp3vulaPObYBdSVomLOh7NmpmXA
PONrPh5ebPXkRBKOHb54l1KbdutnQvIN4RhuPSP/66KwvQ4ewg973P0Eo4eVqaUA
2SEaltaWr6+3WIXYWjIpIFUUzRAw3BYCydzlr7U8hJcel6qccIaqMPgCGKAow1Bq
ZDTf072y1ztv5XImoOfmV4g5Fafd90ZFvECu94wRbQU++aUDQawA4iowd2zLsDeL
VWHlcFmEB/RU5fOCXNYyv8pbVoPb1c3SlqjSRIyg8db1gwEbu5ASUbaB8rHYO9wY
4mYL//dZFVg8S6hZx9uWy/K6/+gIQHYw4Ly70JgeX1s1fHHI0yrFIY3G6VtSBCPU
KqgXS8vY7MWwpy2bGGFkn1r4O6kgrqfYy16gxHJwsowpCpQVpMI964e+v/JLIban
XJnl2b1d/TRzLoklyw4SNpKjZVxSB6zwpySzNBX+FQpkQWmWVswVebSCDJ+66Wii
MxKhI7cGsxuqHc34JH3Y9JmgjN/Q9BlRyA3pIq4fVdLEUOg82OqTQ54x9QhMtRTw
hWelu1oNHjvDa/NfV5e687nLhwzmj5zMJRMfqhHPNHADpwhIlL7z7c+VBuEt6w54
eGjNX9OXrNbHzmjlbnXcHih5GaNaBr28YRXPJz0ljVknh6PbVlLth6jLzLocoPSz
dS8GeFHkqz2Dj+6M/Dw9Ai01eryY1AOUyT+S/brXkHx3BF2C9gyvI8SStFbBuA/i
qFpiwrDheZzaI3G0Sjrg9qtq+g6q7XiKPa4KnoiFZYZgGR2TBShISBul/+lxszoa
xi/0++Dv4yGfVrDGqneP/punbY68BFFo2FAMKdX3Y0r4PXRi54U0Zo1FJIEVZ/i6
qQeyC5g/lD94gJjh4zSB2fyL84o4N7ZG1LtHJaynJI0zCXW6/9OijHYRMTjwCClJ
0SRWV/s5z0O0qSkZUWdQ1nNEJBt6xfi76p32JkzP9grEJ4VxirbMVA0AQL1syq0G
4syg89TsnOMFPsz3Rr6CfP2wiLpM1nlAYXCsWvaWx47+5v3ql5P/3q3+OatLPcrs
owZo+rX0iZokbQl1moPL/yFzXJMXDB6wirCovBj1THmk+vTFxrYRTjMmeufzVW8W
jO2t+vaMFvQO6DiiteGboZUepdqQ5TMMPQ2TTZ77LWm8hTiG0kDKx5KBW521Iu8/
zdoYehY2XMvMS2Rx296r2fGlD/v07QyTpojYNLXFfkD+e1okJbBiK9YXE3K5vZHo
SAFADi0ruv660SF3EVgoC6i1FQbHrCbDoz7e7xjivLjMOhX0aph11gN8UA+XSv0l
4sZ1HFjEFfXKXdLhrMHyYxuCnzfvqCk/hdnrVWr8VpKy+ypSJ84hgen0zge7M/C7
w0qERSJ/LHoDc3HYQG7kAJTC+rq+/4JlfX7EQXIDevena4A5sel3Ct2suzqmetRl
FhtGy0eXV73kdRG04SHv8pe3QCyLzMZYtGDYsxS5rq2uw4uIbeVdRDN2kYM7cE3p
W+G9IzbU9DPVrE/LC8GKQmHENTBWOrMY/RCx23rFCLfATp9uTdIhh9bztpaGF4Be
ry3VfeAG2wZchl9Fxad1ry82R3eJaylWO7rDUWvegDosqjcwfL2pIpw0afNMQvil
4sQXpE0ltmrbO9AeOy0NYQwGzBLOKLnaE8GEHh+ECOJeuj59fOJjKq5by3icDcmT
Ki8H96kMFafvpry0j5dz7ecIxLVQ+KorrPy/K7b04e4iVJV8jrpLjtRftaVz/9/t
H0W8L8bkKNJ6VuFSJVRnSv8sTq6pQA2EiXd/y0duYiwjlHsn+KsjBmpstNlmgA+4
TaP5FiT0EchBXrFUYJItnPIjJRfOsj3wzn/FI5TD7NwIish//iVsCOYE2mQHzFk+
N6HkHjr+aD9vynQPm2WbVognOiN7ipRMJ3gjspaXMMC5GK+Uw6tFLSqp0OAAj34A
S3KvUXzQby0HVHxf8jjxhwNGxh0zvarABNbPz+WEGsblGhiQm+doby5dxVAoO32J
xeW5FEZoGhjaC9OX6Sf9lLdGYOKVQ3a84V+c5gIulUtgnMoNC97UIcQxl6WR2CDN
OML6YINqkljyJs5njR3Drz91GUKvfS56GMO+QcsV2GrP175w7k6rLkhJrd89h6BR
FwIqMjmQuYqfmpFn/nBN2j+S9UeZ0mf3cY/H3hMTw6pOKqvphQy6jNGvyOgzuzEc
A4bdvJQ3Oi7HKC4l+Q3BNCMfB6qF8CHNrB8JdAxkQU2lnrS35pf/wrmlaDC8at4p
ZlaVBfNiRE0lixFF1RSiDrLZJTnc7nArH50GJQ5VKFoUN7AQgF6LV3Yji/4LupYT
P4nvxBzHBzN5gcjKsCl3Hporvf9hiy8g56k3dbwA2bUwFceXUCHtzoW7xTzzH0PD
tZXNxS87Ef5Ek82P95LkCA==
`pragma protect end_protected
