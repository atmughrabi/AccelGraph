// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
a/iPZQNRckoR6PdJDtisHiLJ35tp7D7oJwZICeb2ytM19SYJZQjlkkQhBf3G2QuI
VW0dlYRQFM3kt6hbmLG8KGz2AQ9NlieOyqQHxPey5jAZmU5QXlHIzPwEC2THKCJm
1YnvWJhJEQainh50aEzDELkX55KbAbvwFzXLDPAVfyg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11616)
24Zfwf9Y/DpqG1cpKI1GLinAB28GyL9ndxs04l+9wwe3RbwnHz8F1lq8RuhbPs+6
6RcSb6ykEt6UCordDKvhxC5Dd9NtVmsXnFbd299C2aNul3T0obT7Dv46q2+JRVII
zBcXVpEfiT9YvSvaOVRUgGgza0duP6XbwVeUupZMlwil829PfKSUSvNSFwC1gj6I
5v31WC1TU6ZVsXyPxm0zPjPNFeEvJLFJ/J9AXlulIg0gG7GRheEJV6pTwS0RQDs7
GoISl5jUuUJLaEIG4pdPZI8584OCFr4SbncaDiyQcZDAKx/wsuuASAU20/iTU+Vf
zTy4L2nEZqkv7qB5MUtP0r0fbBhfIphQRI/JkWE5LA3Wl6KIBwy0z92KZDrZ43/z
oMgemH+PEwCYVarNXGoGZQ/fvS+sNn43dcCugjV+Lu9qsH0p05zTPClWoz1o+yiA
mJrH/y5ZYjx14MTLDFuSQ23oMhyquQfRa+JM/IdluQYtfs19b3xIHvlZbj1eAg+l
S4UBNDMR5pYDqGeV5PUiFEsaQVMqZQnCpWATJTifuyGbIXyzTeNTWRQ1QH9NkKzV
HDlw/RSPyNRaOyuCDxtZfeBedhJV263ejMMI726IogF39/4Y2fBGy7VpdsYb5SHG
dKBGlE2bev3W2q2+n+pE3pi2aDmZlyXZDaFUp58cp4GYW+gNCbuevVYpiJbAYLYb
Jtj74zbU4n9gyJZ48fjG0S7pY/9eotHlt43XfDlWALfKlMwPJQD4t3sgZuCppZ5C
L5G4d5NYFbEGbYFsKCAWORiUj+ecuh4giewyCLX8Z36C76ISHQq52kwUmF6tzZj+
IKjTcKZcKVfd9gtl60ifXc0A7fhx0h9Y1NIyJSm31dOG9US1dga+wpexPCE51NMH
B4GqinRIkSyoLpJnrClz+5RnxVBidtiLq2udhcdETZbmbwi4lmnuWvGQZsJEkYXJ
6YBtA3HDZ/wJ9S9EUfPP10iSNKrGJL5ude0w1re8UuEnLcgnFT1NXATf2AD4Bf9L
xW6/AZoYJKOnsJGKtxjA81Z5/tG53DtaJeeYhMOMIoUXWaLcbyHHgA+RbQkk6Spe
uvVLQcYmsC2WJ8r/AGdpYN3q81l//KPLmVRyauTU9mhboq/DMQvQMYSYRAIRg131
Ls40/4eis/XMEVVCAMlz+7rOUEuKi4BYjQ6ainkm6aK8Q35mSnw6cwEYF0gINWN5
rTELqDa6qH1T4a92btR++AKjl4c7JcTEoNckvHHKvbQr3+C0V8BgvXhRhP4s0CAI
8Naqoes2yVfhXv8C5vBZa5IJ8GxsDs1hY1GapgCbMn/YMpjAE8TVQqtEKDnUa+xg
nU/Wz/CpWNJAVFQ/VmcDGvErqtVop322gMhVAs99UUH6NYt0TIsXXzgu7Nt6g8Q1
NqGsA5I2YqXj4U0oJA2/s9lDizHGIfNPa7NIbsuN3klbva76YZ5GSab4NPlCwI4C
Qkblpd4ROJ1cGmbzqRa+JQqpEIx6iMzP0EzPi0KCDSsDCUjUG0aQ4CrkQY0Pm1q5
dT/sdkyPqXIrIDvrPHFpf8vGqE7Gf9gxOgoquspSVM5iqjFF+hkujxEjca/Pyv05
DrokY2D4SLnggCLNe5d+QrVJpGH7NG6Imc0A7kEmlo33xLXuHYy0XjFi7n61YUik
exx9kTevj/VlhPPJRh/fy20uefoWOd4Ae5QlGB1zZ+ylPw81/XN4+Pbbh1lnkSGc
cDZqAWTkucjk861+QoOYohXWN468s9SNAfBdBBiqG1J0PE6LuEZJW/eU31y7FyNF
G+H7kes4wNX2zJpWf8r0DQ95kw/BFkX1S3PmZQfrsOWhLnArKDxkkoD/8EihEr+F
ZOExKWn8QZJnpfhtTOp33Al/9cped4ojyLhgYgETS0IDKHsbQev/5udkjEiv97F7
B3IFpK5EMFBTXS1l/U9T+dvlyM4WgVEuO6BWWipclYvUT039yXhAz+Lgp2OMZPyk
XQ527OOLWDDqKdbWa4IoAX9ppE2HenYDERPONEuHK6r9iFaxdFI3lt1yz/5iAa2z
YdEHuGkHR5ALigd48u08q4OXcWCLq0auQ/GHyMWff42WRKXfV4nUJRHj+pOxqZeX
3jSwqtDzHG/DbZNjFTFlFBc2eEXe26f31fncmZzNjXVlV7S1dVuIh0glRBM7vqDe
3+Ot57tjllUoclxh8CYgxblVOMG31r2xHg7hdR2pSC4e+IvbsRHIDSYX4CRX8FSj
s/mNWeu3B52jLxXD7ODEzmTBFfP2H8C22wb9nhXusj4EaRy2/pz64QpxjbhcJche
S5onJOF/3yMmIQq+cxyhElJOcvrQBHUFaFbLKPn0gMjHVr9x4xVC8NUx1of4GRVC
CoLeoa953JE+0an0A8iyJRm/NoRvoTVgPGPLQLpVicf9xCm2rXXCA73z3RhOgcl9
9AvqCPttIqpi/CShTfKIdw94DQnTvBKIsfLhqfeUisCzNzGj8ne1xDPrUOc5Vl1Z
tVmz0/9AtlqcfBV1sfYSgtNppzzojziASi14mjDBwA+7bljd4fiN1XLTbNVvDzcZ
tUvSR3pCzmvnGhrIoNeC+lJiryKc5gKS7h88JsSC9ngT3gQtqfQWxHsjegPZ3aX3
OhB5I8B1UTEU0RtRJ5N6Wr0HV8FeSvZYeXJuwjFukZkbxLYsYFYUokBmXdDjYRyZ
Lsau9kW6FR3KFQXGEbghyVg2HQtNTtdRIC9D/A6KfomtWGmyxkIAP5VDLb5/nYUU
ADC+z9/E6jn8ATybtnUTuobPcWEINDPnJUpZMHrHvJbfpcJ/C8ZICWAuEjran4ne
RN9Am4wiGNGq1UHjiJHwzaWitPWuswT9C6U0iE93SZToGrc2MaROhIco5PzIvrGL
pYLVwqPue7tKkNWyzqSMMHOiBdOwxX1OWOCDSO9liRc8EM4PhKRoJyZaN13B1+pg
p53mTKA+4u/d7GxbFe9EYLvhv70PZvfp5JirvhZfPmiRFOcxEmmpO+/HiltgTz1U
R10GlqAXAQhkiJdKJnp1TUhd+KpA8WBZ8tQ5ZZu4TLHhgFR7Zr9iWN/HcXWlcVMm
dvE/LhRs5tQ2hbgXmwv7IZWV8TuIclwQn8m70oUi7NP0JZ8LIVskTK++Pu4pjfiH
8XeiBx1m2mWLcV9GlrvDx9cbxypAmvdyzOEihog52e2nKzPz5Yx/LystwJA1h8eT
Bajgexw/4PTKnJuk244nO8/O4kKdZA4wJ8Kl33luqRxe/IAMAB7z/tkIXQsnwwEM
xwk8QqldQYdlrttjw/Na/rtoOl0+ENxvNOLuriL+hSb1f8FeVbm+wj2pjNiyrBIt
A7grqsWU1YDcSBL+XtUYYe8hD2fxZwpE0NzS3h8Zfjma+IEjEcYcSbXyie9i+uKh
2hjxf1aAIHduxx6noR4Oj72eMGA8FtSQQ/XosvaakoudToK7yRrhvrxDFipczqX2
MGW0a8ZFBuO52Y7MBhccWH/BqORo9zuIqMHpMW6uJyWMtUSFMi2Teim+qbTdycqT
wmO26dBI5Th3u05TfESkODvmp9LCJbDxTkYcMaAo1GqYnuHc8R3f4E0imfPunL74
a9EpE+FaPntkfwELWw6e8dYDfEpVGAOSB3ntxKW3DEIbozgWDUzTJQ7lo46CDOa0
JmlYJKdRFZkxSSRKsx75zZC7kJX4fI7dyeLnTaEX3NsFoHz3NvxXl0URt8dZqm9g
FG/HyqKp7G+GhYw7Rcj+c3XbNcEzgmBA8vbL4xz1uEzxl7AWt1Rs3OgqxXdMM2mO
2iesEIbWxrmKt3/Neq8uOuQGfv3ZWVUMb/mJ9HcpOprmvSNHvPa/aDNhJYJI7QLK
qPW45Ys5oz/ccWJmQbtWvsMeYjqlf8//22RQMIQ5e7DKPsVZt+NJ7+jPJ/AXGOe2
cVUdF3sXT/ghOXW2AU33odsunNmd1luRq1+yDscWKFT8xKDGToOqGBA2NA8qG1SL
bAAKneP3g30yKd7aNZ7P7Fa6IqFqZelkapaBN9y6zYYRuPmR3BzDC8BSvKEGeJJY
Sn0KZF6sYxs8+ylzGYSEgZtWT/Dm2RIcI1QSEPlEHT9ZAOEeo77XRy2T+S3vSTIf
VV87wM/k69kDuGk2grxowfp0jxh6/VbeHpwrR0r1vp522fKAmLJIOA2JqJXU95KB
ayIXprVklkB7PfQTCcGFJNQvMCHRTrTPq9704BGcDWTNHZEM1JlM/I9SY6Kl+NEl
IDzRUbpfHErWudkGW+9fjCnGR8kA1VnCDlZ4KXhSE+brekIMQh63H5U/mpBN7DPR
sPH9YH9VH32uS4mItBSPQZOQnYtignFyeEYSv9BNPL1hET9pcKxhDcEHSz5ZfW0a
i7pFm0OlqikYNUkNzbmES7zeF9SNDfxjyW61zd5LHMWpZrOaqwNpSAipq9xuZJgj
spiHaqhrflprPU8Ro+n77zR10Y0ACW8UmCydvzbxT+woyYyvgRSNxNn6FQlnarFy
fjbK8cMfesMIyAiqfYGce2fnogQuBqOZEeKd291/AyRRO+GSFC7bY4V0i3rIwt09
pIjzTqxURGpJMXS8UKsl07g9u3nP8gVXgUOV+zNANKdAqIXiDW8dvFHt1and+9zY
W8VMiMAITZ1GiD75PHMt8N8U43tMGiOLlMfl1BkT6JISXJeMnWkQGH+H1BX2cbdw
NNCED/pCJDJdyNov/eN40qjcTZ4E+9rBDPmVKagmnFqrYHhNBkRIeYg5YtEk5/DJ
pxND8uYZt+4XjHrREh74eoA2ZjBjiOAkxzujFIm+IKOKk59X1wWDAM+ZVSh50S2Y
7u10tGLus5M9Ko0c2/OzcaQYZ/Dp1G3irE6r/XbJzGwI/eZv6Xl8I4VNZ6TbSC6Q
hJUm0JrBAQiqocCB8j/PXdD96UdTKwfxmGBCCoMyWa9Aq6cWsiBH3aqrFV8iEfPs
0hujW2Ta3PgKwxSUeaI/+u/rFw2DgzD7pbeXlwfleZD2o64rQIU6p6Ed42gokCpo
qJ/HN+xUYW+4Hbmu0X/ZjrgesHFWTs2E4nWM7AULDel5QdDZD0nfqZpdciZrO87D
7fW01m5rpB8uAggVpV5bq5pHo+dsVkwkwOM4xH26lwuCXDuF2w7N9Dxq3EbuLpRA
l0boCRMK2bAak1kLf0KqrNySSO5+EuYtTLT227hqvAXLUKIxbQAdwa5dkYWlXLE4
QMCQvRPWVF7FmNWkI3oSlEsOXyiXfmPl9HkHv3to/FBPap4RULXqJaCWzv5pL0/H
FATf5mvZFAhrcwd/6M07xS6+bgpfozduavCSKdkPd7XnkYMPso+j5YjmbfVjgMfL
YeMLbLS07IeFFClzhqlFy5zsLdB+zx+Q6Wx0+oL9FRlqAmLOAS4BPYSDzNovCOiO
LeWReJrzW4n1alb1oBK6b/EwTLINEkx+iiF5MotqfkyHycyMGItEp3Xj7tYJkO6T
A8z1HNN8c/QG8fXzOFLh1nFMzfUd0SzC2oQBsFhdywGqHJJOokOC61srzbA3Ks+G
BniA/icdHL0aA+S81nDq+acJEGsdulcYtGDWIj+aS7Sz3iapVRfk1fPPooldNkZJ
IE0kipGjdc+28YJ7yqqv+f/mvGOGuVUm0dwwSX1taTHdvnjuy2yQ9KbIP+c+cvQo
uvAC3YV56j51edEr8EXv4FK7a0cgjE7qT+/VI9OBrTBQbU8y4dc/NBPguY4EBam0
faC1Vbe/9b7OkmThEnKH432S0hRgYKcqQ7zt0eFuCjrX8yAxYyrgN3saARtqGowe
u2uVNM6aqsvthylm1oxaTPJ100a1f7xDUA0yLDKbhseKpl2LX+rKJR0yftGtZxR+
KxSqxgTi3/KppSOXDmdnW1/HiPYde7wtxY+Z4ro0EkS22My1mKXv4aKtnV3/rG4U
fl0f2mxRz7W5fpOHsUjACXhTdaGhFpenAfIi3V7lE1owhWPODOHOKyDT3nxAA23K
HLy+/BporVevdCwP0e1ua0S2r+btHcHRpYhZs46aIMHiU389Id60JauidQ5FKlUd
3Uguzz5tfsVGnSY1b6AXhO8MdOUrxdI0jaLYAMK5plGxz881uj2sHrqe4S5OxtjG
eRbf2yqbTbTZ24jX+tGn/v48WPLeJ50tasxQHInISMXihjnSM388kPeaJpz3oy7d
OTqxAFRoYAfXt/lSDXUJmcY9MjqH9iLNiCMLW/2ozBfjQM754EXzib/VD4dUOjkm
DWd3m+SmrEJ2TdxBLHkTfQOyyNQFaZorPDk4XaA3sNudINFtCfAC8fPcLBIn8vvC
BERju1ybXBK3pKS5uGh4C+cJ7TDVUA2KEHYgG7KeoR4mk5CJZcx8dBqJD5MEeJHR
R82QTwacu/Hc5TTu6ooONBiNznwrzcm2Yic1m1qNCXctYdqYQ9Ud+vGqr3dF0obb
A3u/Trav8y3S5yUI0UC0Io0yQ6L2PP+x7gr2fMN0xCmlI8lB9mNTEAusi/MGy2FU
oj72YsU5zPZD0/Bd9OadW30x7AAyPJHl1oo6pYuVkz9HT7RNv+YTN+6Mb0EQdXZT
Jv4FIV6iJXyA5YA4Uh97fI7mEo0EjM4igElLZ2DOCpncnOR+jv+ExuDNgVDzGFjS
mA8RLlX5M/kWeg5RaXFXamSRDyi3h9wQFitIgYn3654wRmnmhvuLcKz30H0fG0Un
OdvAPAk7ot9Jvvaawevluz123PGfLE2o/eG7MJXFwfbeaqMgL+xhSl6EBkvSlikH
seaQfvkHNhXBaINN18ptcv1M7vS055ztVdhGM4K7kF9DePWgYH0cqxLGyO8OrqsH
QJcTC1MkMXSvey5Vntr1eFGwTQbseV14MSO2sCeH4ZACFs2vbQKi02dG7hKrR08C
4NcBJVY0iYlkHYNipBu5B8o/wct/YT7cu/kZgJMhc20P7QrOTBmPhBip5jZu2MnG
GKjXA72sz+yXIqa58OyempMu9qM1puOIQUHD78cxLVwRTcKCqIal6I+aXcctX4Is
0XkJ4koYnNq2dn7x3o3kFwHMDZBNpjyvApLOCFNiMX4/ZgTmZ+OIcCl9hJGKghma
dq1E/VixSVcgpRx9gC7bclpm++MfxUSC3XQYGrkbNyMoMI63ukuwYS5/I0she45e
a9ERJ0w35G2O+zvMqZRBcxEqf0RZJc7sAkBtUMK7ow4ybAcw4t7VmJ5qKMUXBNDL
G3lQCRNY8ZHnDVrMgUCZm7h/pCzOHUAntgcNdfHQQzUbi4ZKJieU3ucemWssOmE1
bWs2qi5f9WI3ufxw0vk40aM7+x7k9+DfUmZ1Kc6dYrgDd+uu37brnwhDJkJAMjUo
CsSH6Zv5orWFMk67IX/yeMdwnXfKbQgzKB2wxCEpq6Otq/XRLNcT6tac7odO2avb
sjFBkOv/eHTFCU89U96+c0/4y+snWCw1DlP3fPHogIIoqMyDb8zpZ5L0UNuAMxAt
Lc7mOi17h585/Bf+FFI45DOC8xo/jm5QErxYIVvQKZGooiOJEbCrqJTYgd36zKYK
qOVUadfdJ9kw1kIxy5XtgiWiZFGveF9Qpya5silBmY8FQm3hSiDyqO143Y4PkFQa
XaGN+Qa3zhrd8bRRz6mvTOBaWerZUmuGlOiyvQl1Y/YEy0B3gf4vqonVu9qRj5a9
7BVyI7GYnvikhuiTXH9NWB4Stb9o+jmdzp6TuJs9VTCu4SMsgh/Zt/wUrIza618D
xQxpIT6iZkjMxo70EbYNBLukIV2asNn8/L+BBHbMC6Yj4lGbBpfyJpJfhmhHzD2V
8FepX3ZZPCB2WJmglC9fd8R6GhpjNQp/4R3V42ymJK4ecqdy1ml0kC1iIkbNeTu4
dWc57PwnVNfezYf4zdjRghMokbMBxoakdWotLGKSOne05lJHEsO3d3pc9MGXb4jP
EddyS9nEGyDiad0jykuymrSKzV0xvxJ/+2G+BEJ2fX8UxtroJNHWqFHrFdOal/1r
0TBF7wDJ3oSNRd6CxvkyxHktXNoQYt0bWwtkN0khMUfRiXJPlTDPjjRsRILr5hHt
SgEBWMY8038lGn8uIICp0yFxN1vxjBWXpEFFJITY822KnrsX1w1qBBnRa12kivtc
vj/qF0K0bjtattnStuQpy4Wxm5sT0wq6ToJC0J8nRkUnN7mBfFCc216oxI8AAiJo
6rT1as0MhPnqxQmqChzSpoVAGXWF0aPw0+dIJPrDBdpXqLz1OMd6NTJusY/pwtYG
cSzB35nsB6VGSHtfWBTx3oEFYWpoMKY6O8tjubkpHKvuoK+b55cOvBX5/r69/Qmp
HlPcSPVKTvhItcbLjOTCqK5ftEw7cJ+WaLJ15VI+jDngMuR7KuXGF2IZDNixXBE2
zVErYUstvFjkI9iG7KYJieDX8MhsJZ7yae334dRXi2JaHd5m9S4242+ZXFQCBBlo
6E1xd8J9ZmjbYO4oMs/X+AUdfJzqYbzzsAuUDJRIgo1X0K5K3Cb4tncN2DGiNmHh
eWCuyVGhOtUYYsdmo3yx6OJ5AK33X6UO/8gIMEtCEst9FZtsuv739stp0whSOjfD
Uz1HMW/4gH3mfpSYATR4JRNr8I3h4RluCMiRtCYP84Uz6FL+lXYpvJzzn/ip8Xzz
ogtIkQoRdnkv5JJDc1uBSrLx+vpI4FdTR8ZbRsXBASB6A/8Nrie3fMyeAoYVkzeX
7wpL9Uy6NJYp3YgJB8q6CwWkfTW1Q4+a41Qx9ZJm+vZsAYB+2OM4DxVtzAxP1a3P
Qpe8faCDEi5Rp/9p8USIVbCO339YH42LZkoPJlezBRSyF1TINXTDRNSJlNCcwHFC
zNMfoyUsOmL3ySqiiGKSvpz3W/odJqeaPaML7o2OKbGuxTWq1wPG0jQAIhNqiN1O
MMs5BznvIQrPcFS1l3xrzTZbXnoZUju/3O0goJ33wUiGS5SjZtPNa7pChYquMTqd
FTZPzwc6Ucp3ZKyMS3zy3BPVtLWRu+FN5+LO9s+yNluPiJtW27/cYHX6y7oPytYy
ZW1S/2/0+VgJ4IdMNokeQZfU5HN67KVFT4xwmxRS1jGqmvgrTrI0h+hXCGz9HGgC
Nt8czP3DwJH0AUmzpfL3robE2pTdkc2gsDK68jIqAjajA9mriCSx5sb5gOjFTPzU
uk8xUfM7HWVUbUAC37HG7yYOyRY4eBCaHcqchfwlrbTqmOx7X+jJM2SaJM9Ehd+L
lKAXFpJStdNDDCGQEVH+mR0NGj1oJrLSrD8ceG0DtfsGDVdd2Y+NzHU7MizwwgAM
wDXrmLN395aSRxwL8sgKqYGcyAq9kxxDWU2at2An2zcEOd0RCaaoR+WiMkcOH2Tx
A4nSxKlANN2OnIF0VKTRPYYoTUEkWoXd08ddbsikswcfAI8PZKEc0i3C+E4KsxWv
rT85PJwHOFETpUYvmkqJvuKOWKK6YwBh1xZ+IYQ/04MbKdRcofEx5faTJPu180vK
xk2jlOdHOtDZbxDWnF03x84CLA+a1rCDjkpAuGCWbyiEMSzBZy48UcW1u70ZbWf3
2VfKgiEP5X1zQFrcVmjIp/K1zUffRN2Qz4ijOIHMKUrP3h/Z7nthcr0DGoZwj4Na
+/CyLIGYcPsy/ZNe3Wz0WQji9SzrhwpPjjN5kc3iMXzVRkeEGZoGmmU23OvCEv5Q
ugq3MNvvO53c7eLjKniRWLj1rXwSMbLLkfnCK6UOa3tCI7Syc/YLPgxrU0OlBXr1
kajzjIWPg4tPW/DmRwdGwTeu1A8Knc6ktrPSU46EIXx/fbXZhgbMeauwoxPH/PjN
eSnIXiADT5ie9CmSdry4X5bn2pGMbAgty06ijJeyfYZGG1bF6EMHcqdHp4EIV76v
U1z99vtVQEO+y638zewx7Qr8XP4Ae/by7pGX6tUEr7ilufxAWRI8CIUp7XHKM8hd
guS4JqoPIjdg2fD9XIZZYuPcBbZP1ZW0uwpOGewDJsAvLNs3aBGikXO4hMl/3IRy
BZUDMFQ4FMLuc+90yrfBgx52+ER6QXczxa7VKyvaZyqunNM9uwTcm8SKY8FRvJOf
+TcnANNbk+GlCrxReYEN9uANXZzjg/6sQUfpZSoe5swErCmYaERRn3aI/r3fBjEq
WGgtUZbGh+cgVaihU4jkdFP1tQMvqb3NeETjCfa1PtRevrIeMIK3VrzXd0rxiVaQ
tS8UuNPf+urqrx/xseoFLA+5nzKLNY4PBcFsxz14uvsTO+o0PLtEydVoEKulbV9h
18XYteknn+ucItDBE66ZgMV/GjNphybPIj7tMMcdmGl6PkvHPi3ZeLxG6oIGYXXp
8rn+9PEjCjYAHcLXH5exgAoA2/BXZFqh5gG9Rq7/khPHQd2MtSJiC7xCNdUILR38
tFMSoFtLNXcfNJsrNswMZQPl7CdTB4W2zgzPape3/yq4ktCvXv/zJM0Lrge7+Fs2
7Sg0DsB6H1gNm8bO4herk9BoGzAW7URzAomC5Y/q4GmeS/eTF7NtIDq5/tR/67cK
r10TMrxTQs7tE7KfXeOw2SNGar4aXM1LHnd5sfdwlfD6kgw7pn2x/+hA+eAtSXsd
OKGYEKM2P3vGQgAMlr9o/nvTB5dSAqSJqQ1fKnW/UlOIY1ueoz5gJSbJiXNsXAtZ
cV4PfKuSrUgghAocgOXeyx/Xyi3Bb+JiHXKUXaFbfKOYOdu81/r2IKg7e1m3ryzI
Mv6KZUZ8MW0gqMx6Fp+u+0pLjDaMYkGcw1dQy0sF8xvn6RVpw+NzIX4MDa7J7PgH
g8K+WUMJPxSsdg4IQznXe8wEs1k/cRZF6Fr094gzQM1OnAY/8EXNkrdpL1Y9uH3Q
UVhnCqiSi1uTH6mvRzZJdhwWA7fJHFFzVf9LZwpG7oauOT+vsvd1yYZu1Wwh8cTa
XBN5En8b8vZearlWxeXzVI/cPsjoseyGCAEbKbzlrtdxP9+obfjXyMOrB7T9W6mD
A5FxfyX14zDcCMowxWPUDpafYEv6aL70uHa7K2olukIcgfTkM37gFcaVc8lGsytd
ICLks7bcbXM7N1cstrjErR4DvaRujy4N4QYpqTQwCK5EH/N3sRhai1OmUHGEEz75
EytM8YNgdUEIrRrEuwgptLLjEqEK9Jro6s5Bfue0IgxLQgjb1itRyCBjKmmMBYG1
Weyg6dCBdEFvh59dyjGUM0wx5MvhgiyvCO5cLLwbr54+LuvyFrp20hPMw1EUQzJ4
201ItEOXo2p9cIaBBXeY24N8O/7YBdfQN2ZB1XC4eGSu2X5DlDIrSh7l/biHGanK
JXLNz/CSpPE1bjAgEiotpkVcYFB5SrMd90TGnnIQGIweGmhk+1hB5ZhWn8CKnsNm
z9rAnLpMN0vZWq/fmBpx5RktxUG410WJIv1jGzHN5ZnpVJPOo8smI2lRZKPGAlph
YDBRQk/cEx4AiVo5T/iXsjG6bM4Pu+03IwKdSUbOnkQ+UdmHNsjqZvpWPzbdKyat
ws8vWrbLxCVKuNuJ2kdUALQboGNg4spudtblkDSkYSw89Q1yRQtBgXdb6lfiBrso
H4b0RtOGDdJ9/7gyeFOHyR5eENZ1n5ermXqPOSv3RrsqhvW8pUQMDrtRnyG+UPY3
Wyud+h88VMs4vafUcJsYR1CVOLjdtn6vvVubJsFCDUN7cMX7LCmTVy68HOgmfJrs
dOb5rIRbSxGgUuCSKOwlfGHZg6c+IR2141uZIju4p1I2YoIsuzCSdY7TYZC5NsVv
QKdqYyUv5rajqONk/dMxP3PVUda8eleww0MuuC8nkcbQGPmRYwyVDhtY2eu/hs24
uhCRhHNLiNJfvCLjGEVzNal6DI/qeDpHdT1hpvwl4GqlcoUvqy2jGjfJqG+NPjoF
9y6YOco9IsNO+HNGJJkHOY2txn/DZTvgHkyz0dPqy8aT/Tvves/403JUcbU8Hbdr
Jcos5ApJ8ZTRNuHVh1e1fli7Mot7h4SSni6vX/IyIyosptznVAvJjpnqC1uF67b5
/Z8ZcbEJa6FMyHPOvJuqJ1ROw1dlZ8QuI+zHElzrvAC7sUmFKRfuQ4OVPTYYQ1st
7LeOzQ2mr8I35hTsFXhwdNX671pWaX9UL+pKbYAbwalH9clZKAZ2r15ijGqqkVjh
RsW5J9JJjEwKOrQganEpMmMppFXIPjNZiLg/tMFVLkmGIZ05BNS8k2ro9c6YFuZh
Qfrl5tmscYECVLepRCv6QKsq9osDOwJctKItqc5d+r96Xu9WmRadLQaqr5ehJABK
kk1qH9ayMZ9PIp0hjsnqTIcIE/wBgqle8cTFuaCKPhH3U/bsLQcnszKFiqO6VjBZ
9Faf3RzD7JIK+GYIYT8i9QDH1kZ8GJDNXcnmkkNffmDkyfh1WGdilQISNsUFxNEH
RpR9f+dMguemb02oalpSiN9cVIZia5smU6zPdTY1RMj5x0Cw8hZbuNnY7W8tuMqs
VGk9UJbzKoHbyYuIlK6gHQE0sn5Eux9nYV81rgb4QkgJnW8psQBQTG3pOEsQAcVT
apaxobhYKNJM3AuM8w9I4b6bMRlbrcjIZg8kzvOo8+62p1F+ByEOjaOy5LfDisqE
p+e4Lxh9EwagovJaE6Z6c7hhZwVi0cdek6ZDFrNDqZsGLAfChHiFXFcfz1rHZnSJ
COQicH9PzOQEww27q1/hMCs7MZ4DhX9RRGbUzU07XZsnujbQ+gmpsAWvhMuirxWD
qpY/tdFZOxjCJYOWlR5SUhrod+tBGHb+UD2hcO0RuTfqKDcIvqxuZIWKZ7Yh3kr5
0VJfxO5typHIXfT6E16AsarHNrmEDBTNS2Rno1idibL84TTw65cg0qcJPUEZxuVi
PpfHeVXqTYacUKPm3nRQmEmWMf/i4LbNH0D6kb7rHgdkXPTWl/O1grmvhJWf7KgZ
ZELMShKswWN0cIfVO0tSKI1ZTOyEJa/+O7IqcbxdLgRAlkTmeaz6uuITD823iqld
EyxWW4H6AiaSgK/vSoIOIPnfHbaE7XZcLTww+hSaewf+r7WkAKJmlNcu0uOEAgey
MFBkCvkKQHTBH3H2Hha4KFsjg0NOgROJ11T9W5NNnusMpxCckTMUwl9QZ0PhTnWz
8VOQPZBJIHyRWEKJ9GGo4JJE7nHd7tvX/6X0Vq1QWcuHFfUMjW+dyExnHebZCTmb
ZwWm6vtOTtHPQ5x+nKv2evd4zvlDIjsyVEQkMd080dOZtXvpKs11sXYyPb2A7Ncr
lW9G8eKLZoHhPwVKJee/B/qUXUJD47fbO60Z/WN5s63+BSXKy8ErYol9xh3mlpmd
T44fRiF7LdEzJ5iEDok/1eA+6PRnsAt2bKJw6qIiDfxJ3Ci/7spsG/XnqXthv4Bl
f0eRetN2sJ98Bvv1clyB/cPp2dzWWIZE/daC65NoP5r/YZD/3NNm3zGWRkQJZ2lw
mewFkPsEsbNCQXYN57USaVhS0RQuhzqg3Hu8vKChOpaV4OWQfNlssSHOJPxDtiOB
WBx3X+Ts8I2b7RQViEnorcZXj7HWbXri21BvVZgBL/BwLqthSwEdOKMxFyqo+Hr9
8u3LM7AveXTF+33fo/MTtAmszkGme0xsVcXe9RWQHqKJVVqhNdrd3wOu5oRVWed5
AsYiStjZi7aEvrKheKs3ujwK00g9DuD613Qh3i+2OLZ0hpxurxIYPWJQnRrY+qDV
p5zVBnOWjl818uvcQ5G9gozEcqpgCrkhsHo0Qto3aVQ09SyI86WnD+7rqaNKJNGl
U6+WLdjOwXuniIIvXU0hlKgumOr/bEa+TJvFIw1zmstaKrExwDJwLzroX6uVox0R
3kUR9xrQ+q7E1AHzUF0Pi6WpxGeFA2URurnPA3LK6Z580Kh92SJLbXBRPGH9RlUo
baPrbaWSTTxwF7yybHx6o9rKBFUizrDJp/0C2OjsYVE9zq8dp9+PGFMby5Sx241k
DP+MhvTsGWnIjvO/PornX2FFss4jIxhyBHDgyutZXskOPxHdz4aZNPvpJ+m0Zm6D
kJxWEsmwIMYlfMv1R2SdaOA/0t+UGkcaO6r56enX5hrhSYm5Uz+yOrmw8gUU1o57
u2IK4TC1OYnRJA8LJogk6+lKHBYlNbnClSqrSmPQe3Y49fmJhLzaxiSoNDWth7VX
2GtcBZaXUrSaJSIjTKEerwY9n6LnB6ekA3isgFG2mKSjGcEowq1B/xiN1501MPaf
1ERWvCnFF7ssfGadexNqQeuQUd/+IHTU0FkHImb4ZjR4QmlCL0WgONsw2d25xiyf
Vi2SYYN/gnoWphHr3jBoJURZ0eb1q2gfqWPcJaSbW6aU8+cMB82pp9qpoeJYwzfw
YLOt3o8wui3NFUWFIzstFYLtzISmd+VymPsJ71dgQG3xML+OzP2rqzalIBSrLhiV
lNMi0i00+iWsVHvj6FwcYuLsfDNcoA/SpxUZa13kwrmtg8d99OOi5ecp84OLhZCp
0XkcvHjv3eOVRHPoU5TNY5LI8Cck0OpYqBrvLguKooNVY30Q8ccR3yH22/CibQiD
/Cyo6ySKc11Rwbqz/Dhx7Gr6XZVkr/jdesV3IP/O3EcZWvrQF6OLaN+DbXJBeHX8
l0yg+fenTlyohaF2oV89AiU0Zx7dU1r6J3CzOITBrjrjUvuhY0HtKv3+XIKnBLH0
bkCD78w5LhlUtUaui0XdChf15/XsaLBuYpC4XQuUaSSHstHicdeTQF75IcZdkJ6c
eUSLlzrgeQ24adZdjXM0KMGHE6/dJq0YELjBFmxNgH5uFumGh7Bboj0b7JxizkAX
jSHcgN2Wway3PU35itJlv8+8mUnAkELqQWqgaNC/5wv8a9dMoKNNVx8UEemzLK5n
3pj/gnPPoliYBwU3rroXEoSaRa6XkpBwXZC0PAPRtU2fiWbpG3dqD9AJO5EtfJzw
7qZ3s6lnf7AXSvq2YvVIExACX00vA0gm1sqiJBqL8SGxe+xkvABijw8u87e/sQWX
bF/p5FyXoYSAZJSiFFfcT75T+wioOuM2pRzg70C/Veh712rvnObOXdl6b0oYwZen
iFbER6TOj2/ktqDb8kBwS7Jz3yn0JwjESmRgb2Ii6+dLqxwFLQ6dikv+ckFbQqSH
mX9GbTpcz9WKhquaPjpioqX3t+BoUAiS39CMy8sZ7oxhnofYLwp2dbbMkiPCegWm
aMC7fvUOVtm+c5bvPFFugyoS9GiZ+Db0UyKtEj/pmpMS8ozCbmEbWU2uFVbCobzX
dVcK4QkfQELITHKAHCz0oPwomsUAuGxfr+agA+l1CTD9KLUYaT9Od7AMEiPwCYs9
C2rLP/AFRkddGJwEpWD+dhpi2FMD+2bXAOCAxC0jnOZ0PHQBCk5yv5KpDm/9+Yqu
XcOcXdABJ/ixk+s+rt0DQo/45Jq24xnRsFcfiqDYBcCpTZwCrEKG8MXiarGvNMJR
1Z2cl/E2QZn7Cju2IzQKALlNN3oR6AtyqDi5ty6Xagw9P6OuZRBVuocDs7BKH1le
qQJuGgUMLna35YA2ef9TJlaLIXxQXTOwdukJonzIyt0XXSR1L5msiwJ4iELs1MJy
g5b39Ajt9FHEo6odFePsJoRmFEOz6Z+wgYT/UZ0TEVWUsbG4UKGAKY9tVndn/q6g
`pragma protect end_protected
