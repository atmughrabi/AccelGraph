psl_vgpi_inst : psl_vgpi PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig
	);
