// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OeJtRYV3aIEUBUlYOUO5MrItEa6LfdYb0BuUAUvDHIP+p7ZhGsXP43lskYh82nkI
l5oddPJszaraKEkJmCdGGspepZIJHlwVwzu3Cj4Pu6Fr4h2/J5iNlHujEdvCvFQt
SP15AVW8Ht+BhQU5LXQlOo/xwyHAFRDmB6h9RhmlRB4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25392)
MYRjZwSlJ7Q8NLwZdmU4ZUWgEP34XwTcpngFxVvoTVaHmGf78dx14rCoVmtT0ylA
/Pp3kvjTsa5bwm31JIMybe4X0nWDV3MfEMvUZaqKJvngqRE5ojbQ9KINILuokaOn
t1n7FexzokHvYk4a2/13r69G/KoeUsPU5MojBMxsL5FDl6r6uVQ/ueTkGSTW3Ppq
SkeAM8SGN7WnCQT+FT7aqMrPWgqPt0FjhBU/ATbsMz/gn725009cMsMfVvzmLR9T
tyW0s8p4u7FznMAWIJCHXZSEXl1q1J3en5gV5Ht22p5i1Krqil22yqVvoiR0kxO5
LPPZvV9jUhoD/n/wo6h2/8jy06fB9WLqGOjbQr5c9rQvcZMY7ltZ5+938TQGoRmJ
gjHUHAg9xAG0QqEpACi53ojr4H+k2hnNjLkkTwWn34Qb4ie8LUd9DHiaOwWWSqzn
rMjyyZnBbTsP8xozeHw5HGqqLhizesmn1echkBwNLF2JN4oLwgStEAVNHUgUZR9+
UaTkvKbfn6q8YsCMWF/l/2aWrBHqLCFEs/20IrMlI/9CPHSrGeUNz4I7J1P6Nvuu
b3ArwG1NPFaOzDuVpeW5ub+7cfJpVcLlf6NB95j6oYZESs45bxFTIeoLJHWBa3Bs
Ysz4eW6CNoPYW8KWtamOXZkRfyPxWiJgs/ytv5A59hoJ1gP4YmeXJSwISMZdBz7v
xe1uMWXRYeIkZRz+BqCrpP8jpVj1o3LldTKvV0Kih2yrZFsuv8c4qN3HEwpZI/ez
bA83GXdau4+Zer+XJgODXHtpiBDApjD+sunV7yh7NYyZVMU4wG1WmmjXNX16C2e7
RneGFsDjeyBCxr/O/ZsHmwMqArX3wGPq/r7MIna5PUjm5yJRPzt8gmPiq55hSCMU
66rUAYOVKD9xfgH5Hcw3fJhFH3PFI0z9zI7h/DgN4ycFBkPuqA3mrBUqazIeij4l
yfJIQuNVKe8skRe4G/0JQni20E/kRMdmVKTsMZ7DW1S2I1Tclu8zU4q7qMt7ld83
zJsnNwdq3egBbOrSNaQK1LugTECexnYF06/cfXAkekw81mVxtYxv8EfOfa2g+jal
x3qBrQvKAHr1LBh2cwrQ2ZN2jV2PIv0oAmRZjt0rEImc4lumoxjPGW8z16Qk6TCg
QF1ml92ApPcsng2qMdsDLHf3ebworjZhbivX0/cP0AM8DT0IOCWFBGOAnlwdTZEp
7LZYUx2uaF1DLZPvMJi3P6JTEqQRlFtrta8DjRzQXuGffU3NTUxyJj4J/UswzMir
Yr80BpZHSjtUNrY3xnVJ7z1bYdJAuJOKZKa54xgGpYNPE3x/Z4BAlP2sD0WcjsiI
4WOmPpHU9nG9ycFDeuRSrqrOYAvmek25TuJ75jVMEFDi+bx96qviy8xCka1UIUPA
+oot6JB6AQY8WYtiQJj1232eaE18WidITaslmesJmi317CWPCu9QKrpUYTIdjoMu
XFPWQTsp8PqZWxBEgeOoSNGbs0J0CkhRCdIHyEGOYg2wYP50H+PH/uwfs5/vkJd3
xdKU5pECRVdmYIUo8QqWOPMTTjKklOpuU0jIpCnJtIXemDcK/FKlkkuGeEFWDjDB
P2eCLWu9iPICeUrjQDnumjQ7633WQN1CuIkSkVOHJzmgUWqIHlp6uZ/yrXort7Y3
yAAHniPPQmhg+VVjkhaRBHu/5ammJrx/keXeUjnjQktIciLG5yWjKC9CjBVBj6hB
L78n5Sdt1FhWHku05llBoLweQbLA83QZkkUIEVvQzfxwwS016EVwgoRV7Jj9lwpX
p8OkMmub352ZMYevN72HqnRS8yodU33T+o+aHcVJ1Kb2sIQh6e7Lb4TKj6Tjxuol
1KZcKsk1dYYMWwDbPvOkfAU1Hae003rP2mNdXFKL+qBZltrapE4eKTFqqmN1fXfj
43PQpqym0JCXr/Ww4KIiMZpq7XB6kCXYKHnXuONinKB3ABeE6UXlyqX8GpvGvcKM
nTfDW+bzqSIQE7flhsobmqihEDfGtR/NtA27m+KJv93qzu3WgcuKM9l3SO7LakLN
e+Mwkrm7YULB4sk7C3RAoRBMfoVWeV99gDxQ8yKE96CvaaIsdSWoKUGZjTx1vevd
TyEnwuYUZrRv/rApBVxpkHO5JuWAP7/8T5vxl0d/FY4SOSU2g58IYRgGT0ihkaza
eo5pIha+IPqh/TviOl5kSClDMaECpP0OcbfDqeBTDkx/5K+tbSmLk0gJq7VTo4CH
XdunpRK5veGvyh7CYgyKw3JiO5mPQqBR3VmkQvBW1lJGNanErVPQ2hSM21lwAZqv
/NqD7ga3iYubgPghSsD9pmx+Owf0afkVVxrRA9P/Lzb3DKF7WT5Ez16aVIl4gM8q
sZ7C71htgcAAWLrYXzwUD+X6dj9RjU9B6q3nX1a8r41bN4UBYtQ9Z4yrVGVkMtdS
4G9nxhFZmsvIVm6jBYQazTYQRPUhC8L4aOT947GQzuB77Yq0EH0oVXI4IOkL6JrM
7XrZSEv8QIfbeQbB2lgwYsNs3S3TFNO3gRPft08xGMM1DNp6VGe6ThFl4wKLJzW7
iOcqrIyPNJYP3dljAXH5jc2uqo4IjAN3AY/lZ9+DQsJANyPmeb5nNTOeCG97eue4
qPMhyQi2WXFOi8dSMyAuelg/eCIuOJZmdeuXF7FGsyLZXNywcXCe5ddecugPMw2k
kCJyUaAWhwog22t1CIX6fvM6qzwqMDt9xdGf94gq7/SuntKyiQGAjMgtL0eVyOA3
paN/2clbqtPpHvX5K15vIWP1K2EW5A2nwvjl5jybK8M69rDYC4DDyzIUAEcDgYMG
E2/VPZbhyNLwNul+L6YiirxPGYlGl0VcdDHI4ectmWhkCHq/LEaydBYkRdrkvXQC
erXog5T+WVzn8m7SakL1PROmi2V/IiwR5uq8SQk5OWoDLPoJMT6oacNegryYmblS
NEyOqepMQWBg0bIi+9btcNKb/+1sVQTqXQBdrLFp17/vKyXvw2O4TMyuCwL5tZG5
QZXMAgwBya+82kft6Fkrf3HjrrLjtaEFtzKd0DAwI8S2gdFFueBPrKS2/89PLLRp
N543zUIufXemozZJqlrLEGfKxgoTM3Jz1AGW+lBFb9NSqVcmhsri+Z52Jqslv42w
effqt44HLvSyJBSx4kaE9rNe/Q4SiRebzj+k+1asri8jRo9AOS3ZHgKrnib3k5GJ
MY1du1xEyztx4GU5SPWBCwQaWQkokETjt60hISZP4U4KlTzrleiH58/5FpXoYSxA
SAl+qHzpP0yx/WiGtczRkPeUQXAdkp/+axhQB7s/xMUBLWMjIQhgdNIUG8gDDFOJ
usYo+W3UwyAiBsrWGzOwXM35HbYU1NyU+iG/Mg/YduP8LOrcURT1747pTnAdHWYw
SKxFi2XN86YIiVKP+h95wqkkn0sUO0EnbuJpRR9Fyj1MUZENN56B17VfsX7jvaUz
NHwkpcMmHerTcHt//4McAPdqOs5g/3x5qydEuynDm3NQ666FJqHmPvX/cpENH2Bd
J4pZVvroXPe9ao3LA6zYmyzdla3hw6fBtcSh3LmqfNSNiQ2oI8dqyOaFHIXEeR+7
+xfqKTIBOnVlz2tp8ASJXJyj9vtxl2X3C1/fMnO5mc7WzwqVSU2Vhlj1BaSBAlqG
envmsFR9rOlkqsb0STtIx2LLjc4sF4BYpxtX0NzqKxL94OJOI5WAIbY7v3CBwh8c
P7xItS6/a9vN1tS1EmjtLbLpgyswgaAtxkdh7zyk0hLNShxWSElH0to0UUVnoiw+
eD8RWkwoSYQKEHREeb1wNukMDAUfjfKnT/5eL7MmhkhTz8XrFCsbCCF9YGge2fD4
P3r8qfKtRaE1T7hr0ZFriZNmcNpp47+SbT+opa7LIiJmxpx0MA4+wP6XPgu34rtg
GotIsdVkvn4fi9LfwQoHz5GGGtlqBLvqQA0MFa5Nk5ke4GP6Vg8fYRMIKfo2DTTl
lPXhRanbRf1HJC+6xHyE34sm21xtscCtwc8yfqeBjAbo9ZWGV1/lFhyM/7Ag/IFF
/dtGoFE2tXl986DigbW1qvApf/ewK9uGn4ijy2DKkb98qI0vLNr/3N9uFchRVzWm
2aSrc7AEUlkSgAy22+Juk4uAHFv2gVhdJuE+Fx0jG0w34XTXk3j9tLUTWK7gum31
HK2UAymJ21R3ZA61A7GvC10k2h/h5wSOJRymEKNWTP3oCj66IGkvJrksYN9gK+S9
uXRIbZwmXBnRu7/76IfgsW3duVfcDwtgZ8YpkcHdcqnT/mtWMjIN74BQOhyi1NIa
U4+C5TV3RWrbVM2dlH0AJsfE+kvzb36+1Rb6QXgy+B3zl6gaFJ+r87qVUzHb9EC+
eBeYx5PRPJF10K5DaNJ4kZPLxDHv70sahiJlne9lzZV9TyEaZCRM2ijwy7oTP9CD
uHqQNEJkjlYgNWNfZ2BO0x0Lo/NNOk//bdXvpASSAegEZJnlq8dtIpaUMvG5Hy9n
0eL+1NSDFQ583WY5JheSAkXzZ7As2dq6D830f/W/5eE5zXWZoXB/R3XF/YB5JVbf
N+5gB3/qGY0HZYMJ7ZwztQ7T0A5bEqPxNuqBj1z+ajTtTDL5zK8DI6Y0oQEWZVjX
IcoqhqaVQ+EUCmJ0FDVsHCQUQL/MxbbxEbKaO99fLitMGlT6bf+aL6ciutwrC8hp
G1MhgnHerq+WJQzDvXd0S73c6O3fu+OmnU0cbb/JH3wkWjcmNke8vp7RBJrDG8gA
WjbvwcuYcMQEYPyHPiR5CPRu8QQyhRywINXpyWLOxAy1M08t6c6L/ehXqd6+sZ/3
i4wS5TdbV3qTTQWgAVoqSztzjTZUg7QOYkFiPGiR5P+62tk67c84gwQj3omVptLf
pQM2xwKzRAACU1BX29C8q7eZ42tKtBlezM9QyEruyoYVehhO+ObF8lNwFDsQJhaV
7A/3flBZja0rHiKkJfNRjgqP6uQdlt+Zab/IRgJbJQnYl7Sp/eVo4W/cCrbU5Nka
L9ByokLiQDDUfFj/7cuv54m8cfvnAfF5usnXyf1c60tWdf8sE0T73vqVZMj7EcoO
Ze/OOOBC3pX3UMNGgKSNF33B/knsjXV6Yo/iiMmFprZusw9Zp3vVkLh2ooTKJSiP
plk4+68QF3RydJF8nbxoDNurR0IxuXqE3wANbXM7eFmEYFH/XB4a4a5E0AlFfm0I
NJHAIQyCRENbLQdhaO/ZYKhQWN//9iUdb2/txHRKYyO8r7/Qh3Ez8op7L95IMbmY
DpyK8p/dpt9dF5QHNUMPSEjQP95erXzUSTVqmTP30kYwDZWbWJH95jvpY9AlZ1hT
zC0jjg4ckHXoK1MMUu6LJt2wFBTgVwATzh86b9oaROX5OpmFaq1RqNhdn/D9wnhS
+EB1Lj7dAU/2PEYlb1jWQOU2y49yAWBF3QpUFeen3FW3nKzOC2JZGa5hMSy44Jd0
L2u+8EXGXswPzCef5evEYGKadnH6XSgHid/Y5lcjQF6R63+ziNbpxSTYnCjVhbi/
a7gX7+xtcWdZCEHTsMpc8AGs5bX4wWdfq+yviRJuY/JKkcRsOum6eyGSHEiEizCC
STzRJ3NQ14ye8KQPlsxdl83rdyZD6hlfas4e73l65qGtKT4xMvhQr4gSLJudzl+1
6apYZGztYITy6CCnatCOIHrOMbX21kUnqbEPd02ySIjO4dZAzMD8SaipZxc41LtA
JHI1DsSf7E46eg/hUNlMQAfcV9mFRT2AwENT4EItQzOqJAlLA9+eQB0qoevELMMh
js/Fl4H1V3hcP1KwRv9fKhxQp/gjzxic+zyZoeyn7TFoRbnpWTu47vWUx2xcoocL
ioydx7CSz6ho8C5OoUv+5EsyRDIYmFBpbYp1nhrdeAJKzJe0t34ZGIA9DMf2a9iV
WFi1KwedN2duCDx8Q2IRpMrd8UkgIr2wz8pJm3AuAW5pBjzm2WdlkEJxSkwhEJrc
IhQhQc9z0wQl3iE+hBPuCp9W8vlVFIE8owIIHWa1/xfdHneuhcKgiqGGoEYbGBXJ
sGx16Cd5R96Y/RMdCfjqIoruUFiP+DnHyxTept+YYm2mAlq6S7PgIcPRh7A5gDar
vCrmIZeQzD8gtGmmCDwcaRIS33Zm3xkOWr5voUDAV3Osdw7nt5zB0qogpFAOpl9Z
8QtYr7/cdPJU9Km0rseno0I/dwXMmG6QTL7g7pJeylwJ/33Wj4djo9mxyro/mJBN
hgl56EeNpoIgS7T8aGSRM8sRPhkVzg7SlG5i9HiUenY6y+E8jItXOY6Iwkb/K/wA
YuedWJ4UTEx8FmE8GrAhJYfrMaZxwmRTR+0+3561/QUyTVzA1U/2Vfp0S523/AZt
d20xJMf3mDxpJlXSYxclZRXAqJoPOpjwr5rM2JaC+/9F9jIq431LjdFysa3RXcPw
0Mh5VCCs5WkfRtuT7/PVkBxF9cQ6/LwP/fKUkp7WK9BqYMGMy2aiBcDYU5ivKvr8
G5pwcN3FXlZ+WWOZB6+sCi7y8rNL+QWsmyssiFpV7UGxHR7WMJuRXNHH8eCZ6s2e
Cbe1QVY75crUwdPT7NMrISiQyk3VLZtb800gTU3zt7EM/EwsxD1oE0kF+w6doIg2
L8OVGE3Ivqe8OvueBXQRck4kFnDbne9mY6sHpTAC+XQ48M39hQnpzEIRrO+EmS44
MzHDoCGkjA4ytIXCQLhM84xU86VJneUlRXJL2J4s2Vmrdn9pm7aTGfhx+8VwUaRM
0VOZ6V6dFBhy0jqcsYjEXk24VA0IFEkkvyV/3q3qyWkdYpyHRWNC/12/BemrKc1m
+y4ucqQT3tw49Iu2c0CWXE442EQBvH47gBNZzYQcWBpYcPJigO9fNiiywTXa2P1z
+7VP8x9hvl9wtyQKHbZM0udUnIrI0ub+yt5xrYrflkR5hK2+fXjUE1cX0a6qPUZO
2TZgVvvnH5XTipOYu5einGKN8bawZDjH3Q9QoB2uLW8D0xce2YERQWhEJfh02krr
vaVVNIRoK7/4Mrbb6E4o366vlSSmvchcHFX7bhqq1V1nx/hFmw8j53zfF7Cz2HaR
xQ71u2iYTCP9VIhYzxMw6wPYxXYoSgZpz/sxtP63CKZxcxkpKf1nDhl/NGIs/C6b
ix3RXBVN5/eSx+A/DJl77ulgaVtxJnLkCmHMEYZo5jz4hMqx7VUuqcSShMzbxojb
LoLXhkzdPQ2Cu5ZmwrN2C5iVjGN/i/tJiL4rVTututvZ4WoCxvZwknePltuiv5cu
wUV1gIL0ENzmMVpxg+1VLYTZigJgTd525vCzRlsMQ73qoDV2rDoTUWz2Zej01vID
M3K0R4sl7tckYcPCmU4nfokTz++2r5pO5UKl+iZcGsGux6AErJub3M0w1CuWs77a
2EyjpzlzV0ZvFMXGG065I2HnoCFe6BUobKjjcXVj0OP8x06/iMbn01QlEj/bC0IB
/aEjbqDVHTqkXF96NTomM6HsAdojhGgCQgjaXPgZrApvffSAyKAC4fB/N7nE8tuR
FXBAIwnPXJ6CLNGvhTvm7fW8REXMY9jy49vqWuFU15Po9Rx3jWNQ7TOu3SFPHHmg
OVuwBuSWabldGpOBMKv8fv8vsKeBglJhFYhuf3rdzzzfQAMe3Sg3cKRp0NuTsbz0
T/m1ISBlYIidxmPIU9gjx0dV5hubuIrykCkfteMrtC/dlrDNj0D4MW9OO3KaZ+Y3
K8QGo9uAXIU91MvBvzOGpuawTXD4v6BHOd4zl/2id+Zk9XlQdujWoyEY0GHoMq4z
9ufIpermoW/ZUJ+vsllgvMX1hkmN21mBPPYUD5vdpHVzbouysJasL+MuqZBibods
Vvxx1MCcTqjyz11dioHPzbkSq7PZ+7E5xnrT1tPXXoUGWu3zK2X7cjBQpLtilTU8
kyQRzNAvzWXSkepzU7cA1BCe1E6ehkWVp2R+b5thFl64K+D2s14Vo4Pe1TwJxg+R
6dLBcyIZKY/qLa76Vy54UCqq5ZTCqyD1pCts+TEuWkmZBpSEGaRMQ580jvgr0e0W
eZAUL3phGYxh/z8DzFmb7VONLKtb9z26TSq09RtrPFwOGfKsNnXWCj+ZkpuIoCz6
sONwRc9J+oEMlnkJ93Ij0utjZCu2xaV+qAbnMyePUifVGUwpcmnW9mbbwq5g1aNj
UZPLFeYG9J1PHFsurSSBV8UPlsSBHg1dHu8JvTdZdB210VXQC7MjyDi3dhfG2fhg
aew89h3Yt/cgIlo9kwnFlXDlrxD75iHhu0gdMt5LeAz6vWcwebe5OSNvacx/bLHU
lAp0VyJ6cu54jXoH3kEh4N5ZRfxLizni7V1qifom1qnXthaZBSwq5oOt4oXnU2vY
3zMOlACN6nWEZpIL41xiwtv4bjdhp7qJODP+nHS9mUR5OfQkP686KBeaS7saebdZ
C0Bx8rnqTiXhSd7UR9i/2AMNrfutcC4iMth65xSPWKLkN/PLy6ALtG7YHqhTk5nP
mpcCBF7FEqNgiXrTs5plnfwBVojEtfxcgVCQpEMazLwOT/mUIWxZkSACBSYC0wSG
eSsP5+aV2N0vFbOyPM481CkzrKWcttqUGMWjJb5yNqlFhBPcW9mS7vkRRAAMA/2T
++pMBhWRTJrgVJN1fCYjCzsCVpRhlRUssY0xbw6wNcveVrRr5++6rsDL45GO8ABS
Kf+QMK/EBhHNMkexbsLmab4r18aGtaO2sFfHauxudhsa7/eXzlvojBsNeTIuzHfb
/MT0Mns7joOb0waQkFve58nkk+T0rEN0hXDZwUmehWOXhsS+AscPxUTapr5Y7HK5
234/3W5xo5gG9FzdJDhlk4XPKsSZQJTh3ov3/2s+4px31kbDX442/Ew17yr9Kp/K
qovAz61tMHx8ibUL58njyUDC8x3IFFTQQ7uOlOGRTovONM+YUp82KREpn+6OofXo
bQd2TVaTtHQE1RQEY5k/9GRZHmEmrxWBqXtOB5f7WbU7XJIjNFcaVJ9MTOYA4XAe
SVNpIGjGNSha1YM1IL+PhIf+mvre6MVCAsgiy5Y5InbtdEn+PuLHfFIujupRiEfY
4wf/W1UjnxRxP5oUYiw3AGQK8C8mHTBHN3EuZ4bW7dXU9haJuD8mG5EO6NVCt7c9
W2qMz4fdLsKc8szNAcgERvuNXat6IjwOPyhWgCLB2l8GKghmXIil3rwsMEbG6z3J
flKMSBme9RmHLBIxe+koy59TvuNE5ENETV0HIuL2zhFVSLmISHU5XKn5nughhW3q
22soV5+rOeFjv/ms7ZtaEwJzTBY5rICnkoBCoFSe8yrxRU2uBlYfZNb4nmX7DAxY
CWtn3Vp9cum2mp83W9/xxhYagKEGy2SDG/pSc5EWclZmcL5W9WkQ1RrJEIM2dVFv
jv2puFj4CTtjHiNpsERPQbuz2f25qIS5+peQf/JIt/Y+W4UDSd1lNVoynOk9qa/Z
BMVS2u0JyTLUagjbCHpK5qGtCk2wP3htsIbjWvJtVMJscLNPWiL6Xdat6nQLIgGC
YzMeZ2qOnvtTcN2h+IxGuiNkuhWD7E+MqdEjveHxPGhwWmn90zPcIm6RWwzibOy3
4iWrmnN32EGu5w+/qh+h7nqzVuea0A987BdQuHAbrIzuEy0JMD7ss3q7NZ976S27
Bv1EMUhqQauM2pSj9u3I82AlP3w7d0Wxp3XO/i739RDErAwIUwXo7qL658wxIg2f
bFiCYkUrwQ2dxQyUsl8ZGtdjKh5TMUo0NarXOQifufERMzBqD9pYDUaS0r5B8/br
ED7AgbvzXoBcXFxXEkVhNwEPa51bnzt5vUNCFat/whlUBlkTo84xsH8qr+3iy0Oi
BpSqs+S+s1SmYUb1QtSwjPMBoohVwGLKonQ271qAUfjs9DnyPhNQseXTnS7/GiFX
8ASkU3n6nARBRsNcdR+lUb2pXhohrw7FxOgLwA1w9H0XbdOoak787ZgtkpY0NdAm
mVjiO7e36pI5+OV6EsLeUQk1poHBRxUSJjPPHjxeejQih5Cb+BujOQp9EQ4isQDa
pxfEmZVs27wrUEPbCM6wxqdcZwWfedxvTWv4NZEoa9aFu7XyDO1LGdB1bBkfPFBR
r7rYWkuvqMR1EInf51dtPEHpZJuaxK4oIpO6J7V5BmtZyHjFbIAbcdfMVX5YBzNg
QseTJuJ5PILEJxutgRxpA5rbiq9y6zlekgP/UFK8oGAQK9f0Q3eh1/Jz9oppl5HS
Wzd0PL8ClYMMd+sTsv+7j/3hBhY4/HzO0FFB/fT4q1f0GIyJcbTxPF/yO6/qEg6B
kGF2MmDQDeReWkFec4ZOBr5D05UDLdvPlTuDZqrgnSooDm9GLLurc1wP7r/O/rV9
QzQcMwmryTtiHuNunwY1Z188bidmNmxPRDm7Ru21hYmOIf0RMPdHQiJXGTDboBDp
n41uWgJyu4Yy46g7oZVLQtt66j2AgC+jxLVA5KM9MLIQMwyxzK5jFSpE1oyCNuBz
ffhRzLRsZumjuhhbYEYS8ylhl7v2B7yPv224wQ1N5g/fGpG4o5U9ZMZcOWDzOeFW
TE5CQIXtGc63jhPdsjyEffn5sq4LRyHofqaw42MPyUvehNCQaYcoKo/PV4DxnQrJ
p59OOKfz55GtVt578gPI1jF7M+ylIArnW/WpQkAU3Q1JifAd1IUJ6LBSS64unr3G
Lgk6MLLr8HhLzx8BvO5UMGCGT7z4rlpICcfAsPSA565Rl3ABxCk6YsAN+b/GOJuP
wBxeqUWfKx0qIOInxCXmkYSODrJ7JDrHNFA10/hqBi5zzdxDVq5YVdFpMFNTpFtY
OvMYGVbj8DDnFsJtcBJdlM5Q9Dqt7bNRQt0xZ4vaiTrZtjSeE8dplJyq9St1FjP6
Ze8zT3xrKpSiOOAHDtkKElbwflPoeGYIsFjudMiSfIwWWcbDHwILrU+Zg5MP+FTC
4CtDaR95rNOgYlvYAX7b2Dw017MSsFM3WIj2hX1fzB8G+3DG4636eCD65zILqvVG
wFByJXH+hz+APFScE7vxBi5EtKsxFT+yiLVQp8huexfR2eVYduPVgUFiBAfy5MxF
HJxTTq7inY0KBP1B3Qyg0v1JRRIJ6SPWDgm7R8+DjtUgM1aSLjzZTnjeBLU7KuMH
NdUIf+Fwu0IvSycN++Y9IKy98kjsOrFI4fso4LpstciqTOvJGeXMZWVNogXdGoRH
AJP97Cxen/7kozkafQak2/yDWtjyrXdvXrL6sysatsDuzDfD+HX/oJCgW+fTNDMW
OYexE+DgYoUJuQncD7fp1Q7MhtJEA6t7l+nPPIPLHo0l9VrlpHwfb7QeqCXatFw3
LkgxAjSbR0zyGQ8w2eTHAxs6Mswps1Gg/ifeKyE2eDpOkjbwvCd6t6ZzpntMt33F
BbH91bPcApDIMAlgZLXAVSR9ozETUlOLXk+XMHOV2R8/lv2PHl8zfCcAnMBp/PVV
+kg2YAFQUSx8FfV2I4GlfXAZS4F0unOZCf5mLp3CicXltFenv/pGvip9VU67BFqN
ghs+nEdS9BPwMHgXL5iOT+CLKRveraWYPsn9zSyCjrmXo1j0xBa7zubnyzHjHE5I
daTWo/4Z30QEuIdY9bEor8EJgBBwzPQiuhsrrrRKQW5j1y8MmzeWxwrgwMSXiQqE
Ut0Xc8SS2ptCU5iBKGeEhoVAok9qhX7HS9FMh87mKV+zBHYywqywQ3kMxQZHcPBw
a/Rjkd+f4YnYLjqoa5D1hftQXJy3ae5QqiB1PCbZ8ppBu3WgYaC4UpCkWhRd7+mw
fWUizWW/vcOvw3+6HAMC9pe90+dXyvzl6uc9q89n8Hw8ozA/zc+oQgbv3FKjbEOD
p0Dv4S1nKqEBmZs4/KPTFueLzbV8axTJ4kfd5YBxZNVzn9GI4c6qYK8aSKdtvomQ
r1NLHTu6gS6Gi64y7ykPSa1y1gQAUbs6nk6jBTUHEZ9z+Rn3Yx+Mh/3qxCeu9EYG
ScSNQT5pt2dlGsrKZNGj9rOvTkB18C1cuYKhSYx5tENG+LywkKxqtZDBVc/Fzt5G
/TtjE0YtA7bLgZpSKyJWoHVyu/qfDEtAtPzDbkpptDsaTGr/kf3871IGTr1YXVKE
NNujol2/Um4sbzhlHfIIM2NUdofxaNHT1iGAjmJxql3WH8CHRbE5J2jUiQnswxMN
gXdk++jGo6zixP68Ehxg4R0X+hAtDprPCdEGdDXnS7mGmTXPbrf0SfD5nXQlz2x1
rtKtMBBEq1R4mVD27swb4vkhi7r708WEOKntfSPjypfx0M2FCJI6vTQunrqQvhRv
szHafHFyDETZupQJM0Mes9gnglCbv+bcSNDe9D+hxVuCd3zWOM9PjoihmoMA8uot
kNeKo1z2Q71AMo6FzogeZp+MMIuJm6Ur64ilpxJSrOH5L5uIBlyzv685Q5nhO6Q0
tjEboi4/DBcP/HPk18xwQx6LGyxqc3y3YQPoCYoOJERF+5+HGaMrf/FRuYF3ZvFQ
HBYIaqXtEjicgiCSMwxkuF/ckSPj16CnGO0FdJOOTpKxfL4+2xb4EuzRM8VH+G8I
IMzjM4ehHRZ8nKyGanEY6L8eSfpJXd5uN+nKcQUdr6irojEHEz8s8k6PE3iIiw1+
oJW9xqXxsPqFPQw6MGWod2XZ+qHidlWhqch1+wSExLtCzZ6DDLdP3N1Qklx8fcye
yjknlHDMgZ4u+I5o+OlMGyOClVbgdjcpc0tz6JeYLPidKvPjqUS4X8Y1/QA9vu92
GezM9KnKFGQP4Ra8HVc4M+uJAe6MCepNICOQELQJZmmtA2xFaOo3duITRXbAy2WX
Cjww/TmNgMI3Hhq6Jknb3qSvsCVCF9/uGtN/mXB7BZPDz5X3EUsjxVVrit/4qYby
Xey7jrpD9rdBGRUAig0v1noHXMhhFhMB45PYtLGTOo2KfGI5e64yHFBFRgv82+E7
XviS1OaYML0wifBrAiKJv21za8eveC3bA2QGBYSMg1JnEdWqylPNbF1hGn2Ni7ts
zWGvRsd+oGbrhBaI6WCV9+ADztE3d7LJe8kK37uTSW0eMnpaJYW6LvUgjJh/VwQO
cXHzWNIOpMZfWekZOJgEYmwxAnAElZXn0iEjBU5eRS9B0MNC0MszuyUwsq0wEe3d
C7C/mcpq3OKpwSuI6qiYzj4aE4ty9IawoAufDqHRoTaPDHIY48hUcjJqMRAzVj1w
Krb4yVuI7/QNeDlCKsSiQabbDI/wh7UATm3thmvdb18XuIJyCCpMF9MdIjd9j6zZ
K282/7id6do3ChD/W9XmDK21PM6fxK2+iqaaWOBrZFMSARsTjulm9cbaW/crXAb8
ZFnijKqpJgv1FfrKMf0+c8uxGINqWvE0c4H3DPE7b3WHpZw7tXtNHLn7p1CgDwR6
TdiEzgjrGMRkuE88Pvc4WK7gYY860WzLQZLhJxYbrRNLemHUiGxVe4IOO6YrdEXT
jHXOOks3Bf69NJ4Ni30NSsLeJGZl+huXorJtKd0XBWh6j4HNJkHQLEqWr6Lknvm6
ye90NoIIW4v8QHRCMWH6o6LUJcQArtDXgA4zTH5WplgxJpbowre8fgAjlwYTaezK
HwOJfBpREDqYe8FYgXrXtcZPrF3WYxkAqJbKK0adGTmq92IToDx+E6Mv2jejS44U
7npA8kgJSPWM2NhKphLo6Ud7jgchaW3DqjGP0ai+oX8AH4CL1nMlvLy+MkI7yjD4
imSRQjZkg5CqBF/HyMZUdjI/6865RWwSiUg55v3wS7gph1j0kauRplzJS6Gf9wr/
IRzFdmnIDaPyG5DtVNle13/p9Rbt1FkdhmUp08dvt6G1xNnnbwwOHkwvG1x5Fg2Y
6iuJG81bYo768iL3IXnpY2pXUXostvwdO3i8hYsx7Ia8fePS6xUJtsERHUgfB42Y
OJ/onBIZ9W15ztkjuCYUksRM/B/EOPSgKJcxtRl8GxP0/DOjR+G+NANlKLOvgHEU
GIiKl8qc7+k8ZMJm1JD2e9+8Ai6RvfI/Q+NJ2Pyp/+ylde6Obj0XxqCfS5+7Thg+
ggf+CBokaVSfI9bAn6vBbvvsKR9Mb8WaSQn+10c4LfsJyDtRnYBSEQ/Xz8WY7oRg
0+vWBXTGlkq5Nqw4wkb4enc1148RrVZ1B86Uz7/TA9sd/1PFDs4vF7ogkKT8JSkg
uRG9lAnIjufFVE1gp6LnwyGbobRExN6CiMWxbH+yXBrLjr2GnhfC40RHiq8O9c4+
XmqJVYhzW5k6HgIswfdKtGxW8VqhO7cpKdkghfpMV+kvjUwtGc+OvTrbDflVzqFp
f1dClapU+NWzKfxJr6Ch5SEmMwv6UKbhVjbmmWUEMMmSMdM4TMHeOLo5ho5tAVgY
iPqi0lbIEXjX1xCjET2i4cI+H/Oi1w3Y3Fnt8FEaXOOqXugVoxRKzwMMvH5pWrip
RCXpkd2LvMHrT/6l5p3KH2eYSpu/pMLIiIaPvT9fC4OCYrlRk7CY+fxB6hEWgwVR
k1zUiVIrxCDuCCgTurZqkWAcxlVs5i4OTaW7odPUSjaDy65NIlQbzevu73cyI5OM
1Aw5l45Jj1o6/k/WXSPam5/CDUA+kJUSSXsTkiI/CVE7oWqqS7wjx7gBGjPI57/w
IQPta7GuaJhAFKkuERW37MT1Qc4Ufj09nxaNUtClVKiHLmyn46PoQJKjOF+095S3
jlKnXEDmMWAR5mFBKOkcb9hwZpm1L8M2OLxJRfwAei/hLfQzg+MqZQLhWTYunt64
GX8/Z3Kr2rY0ptOdYfG3Ab0bX5wa49U1cYgU2LdaRLkS0jb4WEqaIWDsoEM3Z4ol
kBMBWaFm4zJxslLKklIBtvK8YlEzrxm0gwz77GyyMfslPAccOvh4FXjs7DSqb62E
cG7oQR4bN3KDpO7gyHDNrnjUNic9WXWWhFiakN3eoS5wulLXHE195OKD3ShYxRb9
X0XLhpEQAFZ7wQ/qGcas/EjOv2ZV4Al6lVbs4VR2U0rsuuqEddbuH8wbmyOvLGTs
3q+dB0ScQ+gKHva5frYpSL1fEmpOtDy3jJDHXqvkmkI1nGGZ1hYvzKAHXQ9wU4mk
ADXQBg2HFyy9ckaHF2okKW25lh77Rtdv8X2GQqvf/6sZxfv+NduIM3vCVkdsTAEa
iBJCvUsY78HiizfFpeaWZOQOn+bSeHomxzGe4p8CHQWE3ahQMrI+3/yhdEttIs2c
m76F7U1o9xLJKiD8iuVeqXMI2r/8M6NZRF/vhYdG515chIR6hZlCcppehK7inxPQ
DPIOwBYn+HjWZ5u3Sj05729lzD78RZz+xZaldCXGGN2TjBq+f7TTi0+gDtCY/J/1
R9t6loruSWCZwl3fiNGgy61Jk9dRQc8R71TL5XE7i2rdPk+bzhxHuFrTmbWXrEuB
Kay+8y1d6peKNojzcnz919swZvvWdplUke03dt0BDMf7ugobfe/UMjIcNhnYBVIz
AWTETvcpWv9wBD7gP86WKmZ6kSsE/IgfKb9Fzrzx0YsUjdAcwvlQlJigdF70kWYf
0JTI4S6FXtWHLh0Q/+jGWOM750V2CxJw7sUrzBF3O1KkscXzk/IEN33vSR+/blmA
rJkWWHEqcdiqTpmRniBcvhUxsWXg7guT87d4K3rEq7Lbr4yjhgfyyWim+DKut6zI
8mBEfFhCHkL4NUcMBEMRXoLEYIshdVdSXK9Pe34F637fqcXgTx/65gFQTMrLiMi7
x45hQNTV//CsMrKHCNeqR7VkGb8VhLcoLGd84J2LqTQ/1WPEJqt1vNswoXXlNAXm
em0eoLrkJbvfEz/lPc76XkR31VozeXbgQhHQxcIWi5WYmKc2aMDeaj5PNV2rN36J
BwPQC9Q490UVoKTd1BPOHe7yKQJxxWPGrfZscMXt/+cu0VAwUPFzfrUOR/omDEk9
QHgYmao+tym+Va3lupUz/1rd2MXPcsiDFY5UdJYnu+iGYxvOcVGlGZkjb/uUj/8A
GXiWQu55uY/XNS8umHhP7+0HG3TQbJ9v5dXOyRCXq4YiMZZjuHc5DsBthb0gmGzy
EEMf+8ssALORsEqJrHKE6oop2bKb/VcsKvOsKzYK4dmy/DBPkjcADGoTJXLAHUKu
QkfXUiljpvRu7l6Xbe1nNMaTmsSADYfEVmb1m9pWkrfl/s5sXIsp8TCf+YfzD7zf
+SoEZkbg1UDgyi53mfa/6djghxirjEfnhlz2Si2qHGYtKFPrMXmhaohtD7vpKf8b
GCsCXajbpudUTZiTNXTWxl5XtGsSbJwDZi/dSCxREATtZrKP/swxG9MGldHOIJIn
Rl3kk4GlZp8LlLpoGeZTjypE0N3DaaCB6W0lg+PyzDMxwu+k6pECriOd99vlxaww
KiNtmgdZnlSp1pjipQyYfE6bS8HXk/rwG+EC2Izt9XYb4AmXWu+bjT3spAcm5a4I
D5vok3iNJzVtdYAtLU7jFsI8JOFERN7VnMuM5N8lk8I/8BJF3A0CCQ/2/NQFq8hw
2Pm9J+9M1zUH8kfMm0nS0FJlRSEsk+0avv4tGARsrjsFcnR5unygtE94qIAJ9qno
nGajmmLf5E9UizjOe3JuDFL3S0o9LLZ2Eqz/JwBOS9iAMKg8jSLqa5/GG+CV126a
Igymx9xp621WELgHbBvpB4ddJZjOgn3cFPCKgAbVGHvorlraKGxbh0tWB173V7Fv
OTu+zxhTSYb9ArAa9rjQowtj6AvnWTlw4jezDzhX28prP+ocNwjPr7LCJF10K0ju
sGFw06HD8oa+hiqM1X0wqh3M/4TKkmwky51p/UJo4vCZPFnqBloTAh2v8raBiEac
tS70veLkBGEjLGU1NkWGXlNFxRghN2x8l5a5bJ/hZKRUT2HFM9hS3unBHopD515w
+O+TqbusW4Po3HtXoEZtlhglFRkck1NdDaTWLSE9zIUIo7QfG2C07coA2hZMsDOE
lKA09wN7sByhLbCu8/OsFZMDQ3nK9AW1nnAysYXmD4akoJ2FHT36brvBnHQnYMa7
2kGmA/pb1geirNHeR4eylV35SeogxNpthLMbbRqPpLAHJwZwQ5n4ZNcA5qD3dJJj
T/+ozP1C055likxf0svPA+GOu0qqgkQ63z7jfbEDGEIGPKrujVQOdoynazaG5dHd
5B1XigNHUiAywXlz9PFd8fIsx3fudz3wvc6KGXXwoAf5sTf/DIErP7l/8w8mTWTv
QwY7rQTY2/lj2ia0nzEk1AI+4YjF5q3zBEXEGSL40KTjXgpTDbwe64c3Xkg2k49V
xXuszbySL5APEhsi5VlRjeRIADnsk7im1SW9iDO92MjD7/A6huffRQUaNBEKf1W+
x+I/UcsXwjELgasFSm8l7ZI2pInOfOfdDXPvwlQlLtSXoc/jVMUhKr0ssMq2s/OH
V5oG8d+MBpDD95SvbOV6kEiP773E9nlajhck7D2GQ0tpRDWYzwhXse7I1IQzYo+9
WZtvL4l4DIWT8DFjaN5NNnBt7KVQdxTDPx3TLUgGE+TsCsAghpNaML7HXODEt8ZZ
3KqKkLXx5eD6MxkI8YeLbAks4YPslafw4zsGuXaMRJbuUJPGK724zbHG38fUL8Hk
CHLp1GjkcsbDTmaXHCgSD28bce8KMpuxMwsrc7Tix1FREOTtiNHMHgCVjH/9oZUC
QNTrprXahGjHPs4YPZPbT4u7P13aWickI21Kojnzl9A3+6BUsNKzxs174Z4ufNZ2
9bQpbhnwgDqzwkFepEvrCr6qL6kTvkKhY3fzTF/56lgTzuqvnTkfCgEhEf8rHF6P
NN2HX7e8XX+gJZgYWoGcIMPqXkb7DpBMMYsCCIL8tYgLK9pZWgo1raPXUzDtdPth
oIDOpCVMmOJK1VnoiWudMZTQVG6VFMh6L2E5qfQ30Ak+7Q98YVscdU9cqIwnD3KO
dTFxO2uXDT+tyV1Lf9heljn2zLd7JbukgLk3wvm9OvdzZzPfJ5HK01AckJLe51e4
r9udM4BNWLawWOkTyNYXJZDZLjcvaQpapYOaKc/CY2nLgEpNcZIco4ZSNGTCuGAh
apA4QU6XXxnnjPvWF6+UkCPkse7lDZbfY6K7Eh7RckEXip4J/YBydWRlQpDfFbth
2+CDTIwMJ4/WYPx+aLqUkNmz+tMaYQ4CqH4EEDoW9V6iOWcefbZbbK6Rq318K0Rd
ZP+cP0fhPJspdlQ12BqXtca2wFTFiPMNV2yV2PYOI4Aj5BD4bt1PbP37++u8FJqm
jyrdQ0s+E4yNIY2pNwZtFelhjaJ0GhJ0noxV+LSGIJFSet/Ulkt8WCgIQd/8Ja4z
pyByXaEd3JffYkbBeOIG22lzccfT+DJb04hN0TOKEcXpuU6cV3k0wC7tSabEW9+8
Tz5UF7I4EKAaUYYib8dnoU1JnzLI+XMWUYnGDlLrw282lyXNn9v66Q8Cz2EMDC35
4LtPYuz66qkASQF4SjjG/JbcZ4337TuSrCJEYqaEW+LIQ8bGJPkO+PrTbFLP4WD2
56umxoilxlokMlZWvmKpcp4Kg4JvYLVgaMxtebsnOt6uC7kj8UMsrw95sx5nFp/Y
g5UDu568NHejIULVKgcwzuTpjfmTuaSU1UI4NvUk0pZnzSo/cxz0C06Ye036TlPK
vIAKwVvi2OpUev5zE0nwx1D8zcPp5tQP9rL2aCe9Dqy69t4uoclyiCWIgrqnkqW7
VFP6rbWHRr1g19ZHQ8XpyqMN7+Oy4U5yxQpTli4r4n9ZmChHHJFcNQu2l09ePJH0
ypsQgU8Z0PGtrkjaJaFQn8K51CDylGM+pMcuMkMeTLY34ppunRCMLXXjLwMO2wpg
OLuhsaouvt+mk/Bga5BeXbTZlpWQyQcw2DMPOw2NiTLLYjDh47hIAr+e0ipXLm9C
VIaOjkbNQ6Tb7Zfd5wNZVXzc7qQrCwsiOo969WvVTHYEqGUxSS6Pss4BZuftMYRx
Gb9ihsnQcLng33h1iACunULFbxeptPtCwME2zoCZYguzEnkw4tY7MWYMdWISgnbS
CQtwXSC5bdFBsbLltGBlz23lnmSCFN9+5ITS3Mt72guUGpnMV0EMMTxxMXZwOh3u
SScvKCxuQdCmDKLPl/appyxurQLBAi4k/a/i5WuLAXHs0yAfUGHhPCJxm4bnf+ha
jHpARQUd7LeSRNcIEeV1SpUyQ5EOnuOk014gkO7kugrHUBCv2pGZ/MWz92h92MOI
itIB6AqobCIvx6DKuatmL+hOOjVwxk2ERoQyCd6sn5R2yQNgJ/fWV0WrfPCCXYur
oVKx15O1b+ThhNwIzatZVwdWB/O0cGBtAKWrCk3eSEYSLb57IV5RL9BqIN+TPpcq
tDskvSF387roerKmujpJPMblGG772zzaDgUrXE0M1q5pz6lZbe+abnVxhVNZUIHh
2mjU8RoxeeaajpJyzEtFpVc2+DO3X0hSsp6/m3VX52b4zgaIsd+6VaS/HqFCXt9S
Sx3cArvQUtOEQpJvq9F1JafSrgnPqgkh1p+uaC0GtXaO6BWmh2OOOPjGGV0j6OBr
7VG+QuGSH32eD/8v+sjzA04+7GQ6JSZwYM2jZvJE/uMN+YKKMbmHxYFdoKCAWcEt
qzTSFbAshWesipxzX8MAPTLklv6tnZpfml7uxF6/QyCIKe2HVlF/93F05VcQEsfX
T35fnNCgrXYDj3NOK6W+W3rDQo+makFISQuIbSzstHHyFe/1xuHn9ciBH8+KJslq
JuRh+cnpcpHq9TUSdS8Z55CKZIUGSsvD67UicsxMcGqa936i8GBFnuI+ZjmL9oSf
e+VYBfAbblRA/JFGK7Ne1VTJVzmNRLVa5QOKpqZGT5iKMMllJyfrpXXXkIJDJJlT
/OzQ2vZLNGkkjhmMldJK98AQf9v5b8sWB+MzQEt49QBuk9zulIfGNuloMq+6NqfZ
OttdEjoMu/G6ptWf3kP3S4lR2d+6gTvLVozVRSrINy73L+HZPpd0av8lJ6jD1/mD
2CeBRd1LLJx/GOlM/StuELUKkADfkQg4bzY7voCpLEqVNyOgf/korj0DJ3+akZ6Q
4MM/rURvahlw1iSB1zIiX8fQAGQCFFPdX9Qer8B3ssnS1smy3788GOlffJDFK/zL
0LAQOLZuk6fOts17U46o8fpGij3kv43oQbqD9jVkv2kKBpMu8+LLWKWVwRTRaG/C
3GeRISIcQxoXaxE8hiDnxXKY/swKe1HTLwK7rx6b2bwr4uYVcewvb0uhY5qSHDAJ
xNWCn7ur6EpqMb00BuvnO+EMQ06oVWaz77RIzEcHc3Ka4kjmTQ1iRNnPrB+Byg9J
nJM+jhWWA2nyV1yJdo5Fj77GSH+88F//K/iEnwFCsRFh2aWvSM7nQVqyJoIlP80s
r+ZBA5b0wgLb89qF8Ug1g7y6FQhIG3oZj0wOILHaakw/iUXHCtVoSqcBqAyCfjWn
XRj2KSGIiHKL4d6bTR0ikk0KufngUEXrBlEfQWq8yDBINanvr1O/FULH/6DiZpHW
YixVEDuTVVzIo5XPTopkXLCLww6G1E/eDEH1h7GDWScnOOziLrFzmY2zFFpCnCdJ
pALA3tJvuONTeiWVM3FgH9JClK3N+jo2eRFT6bAiRLO1kjcWD5ilmW+v5Ap81QI0
FbMyzsUamI6yxkoCbAVLbNDKlgiOsZEuNZg7gzYmF5I3qJ64WDnzbpNxuCX3cVdE
DL/NVkisueS6zir7I2jGvzrCexfIUP3ZSHWoTWJ6QcVSfJMqkc3XkWphHJYePA0e
XpR1AL3vDK15s7NfKsVMKSr4rv71ciJXm2NoAkLM1oH4bpqFg7xF5FI0FKA68WeR
/8gh71JrfUVMHdjF0B50QUhbrKjnCOL0Km6xJW+3Jk3xGquSqnvUVXWIg3eO97OM
Ahu2er4X4KDtrBlQSM3/PNY723Y9zPbXg912O9qhpPZlJlAhDRgGESj8NI3Rh+2H
OW40SIJGk2Xze7f4ZdATRZuhxu58q0GDSTzfviCOsF4xx/Yq7E7j0CiFxROH2u/H
RLNVK1b8dNl9p30auMHw9KbXx/3H24AV/+4/qLENs+JXF0sMrx2btAoxy3D6BikR
pNzQa5hxdIc0D0I8NvuKQgLcjlHkxLVM3TwSNfziuWGkpZn6w4UmprLoFtEXxw/6
N/aMbo2hvXYo2YU0Un5wvn0nLCYXdz6TsikLqF8xqzJGycDsu4GFNchq0x3ILMnv
JiymcPznxS8DqdPZSzvE8YXfQz2y/srfWIZ2+rbrWBofNp0HNunTI7YxxNzVpM6P
uRrVRacrbSjEnSqkKgzEHielX0chNl4pwn9InLJFIf2+vgqgE/1THTvJYLwYTRPp
pGfBpoy6nhJXM81rUIZGstHP7PwyIiNBJrqlyYyqQhSOY//C20H0qx2ZuI8Wf2hi
4P/x/YEJzLA7z3iKzGaloxRsHeGcZ79E1Sm+Ra4WGReclaDdrxvJ1PhgTw4vetmr
gOsbuCQSDt8xrLYmvPCdKHA/ROGgTF5vRYnyP1PKr91aYsfDtTJcRkst6P8wko5M
VVrWZRPiTZnpjgzMjjecKvB5SDM9AtlYQmML6Tk0h4W5fMnrq9CIz4KiPttQwqHE
WyT1R80Z/9Cd7ssMKPUfuie2tNapOpXLiU+aDq0p3xwNYtEmFFbPlAEUT2HZqcWA
qI5BrzSN16rtwHz8QsBGTzoXGYUxZYa9wnmFSAlPb8SmNRSUGPVW/DTg3nbDJqKV
GtcF1dLZt7biw8Y7XIuvsX/xBkbEPcjXQGdO6qTBAewSGcjwf9KvpBKTmWBvsP4t
nN7PcyfKkyYtV7TY2kXSj0FiwVkoZKv1rcWUbnjmYlp2rSe2PPROHK0Mzjqjzjug
47M5b4taqOz1QvwMqLOFazlJiJORc6Mt1IELiKg6J5wIMbcVehxvFGe4yDCiyCSA
90UK50ih1xhPJWR1oOqF6p1ZGBXE0pKki05LKjmxZFJUTG+IT+GO6/R1RdL6LgVO
/vFBdI9OJp7cwGiOo/h+aJtZRMrGG1FqIRpKNGm3poTtpyvw0YVRvAVvPXc9NAmB
E29v2+6z/he9BiNTc7qEuwnhR5Osa0gXquYqCXeF39q/JpzkEcWHYwu0Y4OIiI+r
5/wqsvVzfKTFvdI/jcV9fv71b7Yemvv9fKFNTsiwkSYt0y/qzSi4I0/jEwql+qLU
SxobWPHnDPeA8sTje5k+TTiXll2D1AU0gpvkaweixUG90omFhrhcWSDB05oQrEPq
48ZoxdTQUlSbqmXn4s7RePHUDcqCVHvDQcVZKzp16xC7g5M3jpqQ1xeJOz1w1RhQ
uz4f2+VCL3VK3TF4wxW5NnH064DI0u6riP5a3QJd24HDz0vyjJ+WI06ejgmd5Npu
KQXy1CqisHbbxecEE3rXiq9XjajxWyYB9lU3MkbdcxOm4Hmf/2h5HR+EfYybLX9X
T/g/OmWHesumfIPXJch4EWkvj3DD3mHvfxg7Wy85inhlhK2yhnCGaZnTNmN58fvc
3yM+qncEZmttVZ58aPGJXhlb7Pi2Gdv84AmPxCFasxIqxtQSnlLcLodhJ4gmGATa
ncSRH2eFzD12Thj2deYxdsYW5S0UGRIpOOWLiJTWVeRILs8Aj6tFt9OHLSH48GOi
RLyhjbVL8ygIi5nm50Qtdnla7UqkRnsTslHOP9P1zUPanTDAQK/zMWcrhAWjMm9c
1UUu4N4ahMVCn3MhnZ3CPTiGVx6LoskI2MyhtRV9eHmjIuFGD0ssC62rlzXQL0uZ
ieiQCAjtZPZk9Le/12jcv7/75xGB6nKcHQkYa0ZpxB7SWWSBxpwVq4S6mAqmoZmC
S1vcwHQAQ37ICa1hb4fUYEQI3xBOcUTXz/Vymt1Eh9xWVAUXnGX97iEPRZadELuU
hCzCArzDFV7m3XptAcoAXKQdBqGwYeAlh2U3fiFFUHohAOlH7fIknJHj01ta2Tew
099BP6wrmyBSyPGNEoePd7/Xjhg9RjlXW+lhwclL4x0mQ3o2BcPUqXb3SpPtW3OP
I9TV/gQmkzCiyQn+JlqcrgYL5+G8XW3cONcMtAvFgdbESMOjFg3Rd2WiBoF9vDcB
AFNIzQCyAC3JF9amvkgpZw3PbM1M+a5nlyLbmatXayPgUdIbyknrgQyIy+Mvs1jg
Mz/I6f+/2qMVVWuK3s91ApUoeHo1rUtWzoS481fsBl77s+cW/fdHvU4Hx5PyYDHS
v/mT8VXxT7uc3Jp1K5I6I3Ww8FrsVxMg1op9AgrLvaKwNtW+LDbF3WAFNFSvy9C+
OY84trkoID0MIisrSV6gWcolV7n445t+Y1Srfmb9JwHAZ6osyBlw8xNxcWC5SdQ4
m6xU20WSd8vJ56q8DGIgaE4occX23TUhl5l+bcwNgKNNwJLwCcvjEKOCI/0BZhPK
re9AavXPu8w2n4SLCq6pvQ92x8y8xfTPQ6Jq4VNWbJtn8/CipZ9Et2Vp92xM7NO/
40D3fTvJkqW4S+Ko2UBNmHrqwvjj3nQ+7JvjrSMdVLE+ynz/BMw83C+RNGh5IlZi
geol40kSP/kFRDflF0sH02+WtYwtPCM0HmIuA0fDX5ytCZYAUoCC8A595rC8agBG
fJxKG3FK8msX755cY6CNbUG9ue01NOG0X+W6XPghgTTQMEbEEcQtlBsKCkFQsG5w
6G94H9x3y7DpgvdZB7TKxdvYWRFNJWrl8JlXvvjxEDb7ZAv+23OBJaU8bkaB2zb1
ZoYUiNUI6NdTQKIRsekLVQK9iTcR5mfU3BQa45kagA5ycElnbwzwZs7IqRc5eclB
/R5swWnHDYIRH/VvNKiqaQuuE7WkzeJx03JwqbosGjkuqZWukG8+9Klhq1RwzT54
o4ltBYcePbcES1qKMRihtwYePbcnkkH+kVWgpBeQYGq8v+cWWIzca3Ihz13QijYA
MWU8WaXrNoQAL+rbFsBjD8qLhVtDv2f+lpAknr3GiFLeOgiLPCNwYJknaWg2M70u
dTSLejC6PQx3/PEyVRU6J1DEUz7tzwfnFtyH6dllYzgY9i90Mihf5LBZWnhljWr/
sFmRGAsmbEvwad/TytVyowKHjYjy3Zm1FRybV4oL3O3uCXgV1ve4N0XpJAcHQ4hh
M+Vn9iJIUpw583LnAFlq055UMzn8teJ1fuDouzZaPtvES9QpO4UknDVEO8nhmUGm
peo1EnezOpfZRV4oL8INO20jHbwB7wuOUR5bjowkzv02kiPhjuy52DHQhJCFKKBk
W1zeLubEv8mU51/6UHy8xwE5cprNhIZ4brLV/SGiYB2biBJdQDzRkWJXIvJ+mRtr
LiOO/pmr/7uDP9qLze4FiM2tajZX0Ks9C7+6MrcDWpQI73W/wLQZHM726FgzpX/4
JxQQbGrvPBxo61dt69RnDA+L3Y17IYTLI5cjEr7YzBNtEaoDHu3daw+3s7QSKYun
RBEQRrQ3DT46mmtBJssm/jz8kOzemkrxzxY9G7bXh0HGYFZDGj+DndD+QYSPPAiq
2IRQU41zUyQwegSUKaZlq5JqHvVyYrIz4sjl2nEvv3c1zTX/ijQ75NJfj8h65P2R
Ssf+/yDY6/Tw1xqR1Ogn3v+wHfI1gjrn2q+RnQE9F61DDp9CL7Wkpphlihbh3xeC
2lKvXa1tMXSwIMyXKC927ExjD9gLPYVxB2Jp9t+XAn+naqorwEk4gG1RBooJ2qrA
AziqYzcFeY3sa7rVGff8wHcV9Oi6OQDBQgxZLMtZ9U6SfXjLTEaqm4M3RQOsFgU2
lhLGVXv1zNkqNQDeXDTgMpSmhntG9Hc7rzcIZ/NebDZ3IER+0WojlcjiaFObiLqy
xqKCcVIZiq3vzqgf3ZHPk34FVYx9mXZYFdHXrnL3O6s7ssvGI6iuqBTGLp1i3uiC
QQFC5ODITWlTeq1GYQPwucBktbmm8OBrxOD5PB2dSlHUSUVr4UWH+IDNKFauKRwz
6HcMAHU1DhUox41BUQ2EbtDmdDGpMsOp5NpcAHsFRaDtpCchWMJWyN/1ABGWLu56
+sz+jwBP1f/4EmX14eDYH/Fk8YeKOqq/eg/u0CznY4iK8tRlDvk13TefWO5gKrLO
x712l7X/uCJC9soe4pWR0CNThztiWEX7/CU5SJgbmBjXsUrzF4axRgi4c9o9PisT
Vze87yhZrELopahd9/gGLcF24dh6Kz+egkOqoac0mRUv+xgi57WIjUUwIbgEl7iI
VhewWIJwVGj5OyXseerktHBV405q6b9msdB2oqRDRr9V5SwOvOsqaZ0ZC4VTQrh0
4c74sh+YDK7FyzZ8EQIpkXXZYhUlXfSHfTFJx0NfcZKQqUA7GJkMUPWqI8a0r1qB
y8K+/5Q1U6onhHtQoHVXEQZk1kz/+dVCuRNIzuz8JCYywcKcQj+JL01tHjer3c3Q
cfCRgxNiPxu3KUfLa+JJNMTA6bMOMQcbhf00WX2/PRxfoOj3fU+GaxoCqf47Enuv
XqQkPHABCDKrkSEtaU0aPHw483L+lhOfAIT2j7uyMpTzRHA+gs6slD5dyWhp+KfA
z5/HpIdZChF2ZzbotMLPm2MiKyMT/EFbr667WGZ8k4Qze7EZd6ARelzRXVPb58Sd
YyD0wTqLZx25jBmJkGxrtsMR0y5aEIZebh7b0r0qkDohlyB7fU+xSz0GjmeA+D3D
TlAlz3fViqlihRvhEqUeSvbJUPJgT/0FqQw5xc8DFOXmFku7/fZQFWBOfdlQXSqg
mABQNQKmBDWYHWV/wByA83/LpWpjf9yD50OA3vHd/uIc3G1uN8++/FQ/lpPHX1GV
cMA2zQ9JGoyZWZEoWJHguKwR8+VERfqCXl2j/SWKd5/TVntEt2U6g1AqCHmm5BPi
TKr9TGwBKTLGs+svRGlIzc7Wz0ivXrPFe/R/WrtakRq2h6qsJUw8VYeLl7YJi+6n
Ir/VF/qf9eVJmtB6VWGOga0hz716BwCQbi4zTuCVImDTGZvw2oQuzYBdpeSvKdnH
S6BfBYj1jqVQqW+z8TsKg/Xg2YmB1HTxOTl+piYPHgGcgjNhU9xjfwshKfjfbSk7
73Zj4CE8I2JKPzD3xFexzIw5RE8QD3t/s1VGTSuSzxNAGOvnOsC4aKN5GgJwLTN5
Fs+KVfXQC0aQVp6Gkkf+JXa/Se4bMd2BzktE8aP1kk0fUC278tHvnfaam2LRA6fa
m7CJhkJDT8Mk+sfrZA0xRKHMKAcmsarc0MaqcSgFtpyioMEqLgYolGG0eAUHcSlc
J50fSwQwidLvCCductY+LdJchCUfL+USs+oyMFaqpytbTKoul+8Chqs4Vp2SsAZ8
i+2dOaACGyIEbe9WLbhPYsKlmubOzYaigru/Q4WRh8eWj0pDx7AcEGgutmYuVbrg
/mgBjz6FAjW9enWoBf3Zvt1k+ZpDtm0SrBS40P0M3+/cUpbygB8IIcpWNQmCS3PK
8ktG1yeBhuH4B3OjzjwozQo0o5oQFWJ1vzN/0CP0Sga21eCaseCO/YGnCmavTNmz
7W7vZ1+WdM2E3vSCDsy5WF03Jkd0BY/r0SHgIwaCSJ4SvhLswx/jBCIHQTBFxYHy
/Xgs/r0gbxFNRaR1EU2P5jezcCcynBqF4JfHMeNJwU9Zw6gzLwpMO44DlD3FRYlQ
7z5x8A2tVkfrfhIAkB/9Y9dgCZh2yQ0PQvJl9DiWcfQoAufYqPj9XnPi2ZNn+lqZ
4IS1YDvbyyQQlPyo/hPaljs/dB9bx9Kmlj+OIC6cfG7XEWmN6OBFJBRA8tsnjCmn
d9+LBOP+NbQR2eSqMK0yyb59VOvklSFL6OlnvIdhJ57RpDRPaGW0nSUKz8tj8+OZ
BqTVlMrS5zFIrdNhip0FCLQ5aIN+I7/QugwnsIcGvihYe1rGdWZvMOCVnnM2YCwq
8IK7OrGZXmfOEgIxfR7AqZgnWJiFXjwXDvsr+f7LsI/saymU19kExaKY1W+P0wxS
726fue9Wl6wvs8PYkBiCDCooeOyr3sI+IvSHqnMv7cuyoCBCPB6+UvNxrXl5Wufi
N1xjx/Z1VHuumYgkieo3hkzd+sOAHtvdF1+iaaXzoN6Z6QRnjCDRt973JF5gao5s
6wY1X2GPPysd3Yr6dcVdDLGP1uFkQ71rL0Abm6rABqt123Uy8hbW7PZw3yfiUmLc
++hDlvxqnXqyOvoPV3AooUyo+XQvv2Go23664fOTF/0Y9Xqr8etqM6o753WswE9G
NevwNeKASfMbkvARM+f6oVCa1nwR2vNReolHr0/4FAIAElgGEmqyC8lAUv3BHGd4
EV0b2SNubN1BViHfFhRKxQOs1FSsgbVU9QNHrtX/+EhYCjn5Rka1hYN3yy/UclwL
7f7OfAWReCmQPamQTchFVhHWLeXQsDxa0K2Lxa+Dlvyk8m3PqixpeHSajC88YyXM
dVIfNQvXgZa9Fnl8DrwDr8ccS7IETYL4/W/dHFMuQGLSXeY8YmECfZLJhLjtG26g
XnqUW88XlaWEffKkbb53eUhr71Ui/SnXmnphZ09Duz1zTsQBiSIKcN8MhcCILlF4
ZRkmqyI/PgbdfHYpBfvtxVS1FKGE8WBH7C11hYinb12PuIAGI7QLWMgfIgiS1/T5
6OeUIL6CT7Kr/UsDoq0OcHzxPRDqERlzrGeXu7xK+slwwf5ZLkUoOQ/9idz0AEjz
7JNYxuLX/B7Wehbpk61NCXQ6CuTioownPcE0eaeQXwbD6kyfWY0Y98+djeh/efRu
zx/zkOM1KkMoJ1+NjyRaEmZ8IyMMxjunz2qB+vEHF7EeakI6f5xvIKEx7q3x5y+L
8iUyzttd2t9hV9u/eKUH5q16QkVaSd3BKdrCdG4LGsVbJWYTZt7Gz1iDyKSzIeTk
p5srP5/qRexCG7zs4HY3Hx2hslibWnoebkx9GXnKhIrrNKmuEz0OPVDq14TzZm5H
GeTNP+KiAbheMaFLXLvZhIWStotFm//cfFzh7ldItBn61pgnx144b8YzX2LkNLnh
qBjNuH8Z9bhefo8CJYAXkzXkGI8VWefBKREKcayWj7L5tXaseUhuRyzANXThz3KV
EzQm9ysoyDxMFUdLoMdAhZ4pSJrtpi7sT5HqZhEBAyU0IXIoD4YNaQOpHyuZziFl
2j64BVdrQes2SSnnAssLQVw5Ig3nC8pln8+B7nfZ0y6IXcY9sy6KPT3e+APIK3gX
xD9yGbb8SrQgX4HIHlBjNFOn4cEZgaIjk+cru/Ncthg4TOQ5Ck5Tb1WAmGodSuET
GrqFKfij5iNhcKkpiVzwWQQXQJalQY8QZ/cWNF7BNKQrzo183KnbMgHte4Zp6CPg
XbahS46cVkek/lnxQHOo6dPzeGEl52+YIpUTxnHtXNwbg4/LFK9Bsap7bg9CL/UE
Cik/8DB3AiHQDBF6/eUXMdTyShsUAR4H6mKgeXxlGzZCSBLdfNAD9L8ZRV2Z2RiD
0UGifK8m8JCxlOlrQX0eBBI0+LbbXdtkYk+UQCR/jQ7SmZXmJniPKB+aWgL+kuvg
XpG2KvJ1AyLjrKmHV3qdMtEG7KaxWGEnD11+XcjD3+n3qYbTVlPkcFfatmlc19qH
dUEHUzmM9zAM6a6lx+CKZ/aCSrFNsLu7I5lbFwRaXX1gQTeYalRMYB9ev8jcOZTH
C1tw26CINUEbpxTHQBNldj+PJqA4lhLO9RxVaX9u//WgaaUHvTLPwGK8uoqdOQCw
d4lgCPti9F/rVmvrLUWCIjdcg9xAytelxAO/JW0KrPOSyfaeQeW4kafFIwlHUFW2
tZ+ZgsLYY1XkCvxy2Cys7Za4xUTXTrZv0k5yCYiXjp/CXYB5R89p1dQvonMxkrxC
6cNDgEqkb9X/9J9CtwfWlLYAUZHCw9geadTleawoD7Drzk9U8zzpNqL2e+NLYD4o
PScJuDO8EXftdiIRBROIxvMO7GVlMxAuF3Hm507s3m016R2VUvxQbiGBti8lm51G
GHn+Ga7taL7I7NVHzBrcG8Ae2ZB6gavr8tX3CdFGHmi4VYtMGI0px6t7DLChZDiH
fALuD5mBi5mf5c/Rb7ioHoJhDZUM9AnqX5Ez8dYi46ztXFu9csmEn7Yf8DMcsAWE
Cmwr6Ue+vHkhL5i34ptFEwr5nmEPVHaQeiDgDNFlcLut+z/xat/dvE0u4mQ6Cryv
E4bOmvvJp0KkrgJ6paKu5ngX+UqHNQlVxS36w6QyzO/akMCHzqvTKfAme9VsgvQq
cDm9X8C9yGpWqjfp1GO8Ks7j9g5PFHqzIvWcghEqaCuACHkc4RNQmB4n4N+Z3xHo
/ZfzkCNl77dvD+ynx+GM4l4kqWMkXZH0/hHMCSzq8WRnd6oi+sQNwO25BXvNOAWa
9rxmp93RQ0K12pWuuFfto2fBuZ1yaeULe6nNHchQuTvaB2/IPWha41mUmYtpVH8i
0kF6oUEu5vtbO2G6mTIzQWuRFiW1Sc6VxV6BN5Cn/Wvzg9RIhlGtEJP0PQUtVR7S
5SmBKsmaBNM+3yLBjHU3CTfpbkm7PLnifbPvFSsSHl7oSAbkWIoiLQuCoNX5nWoW
CFDrM4yeLe5Q7+IA30d6UBGC16ahTKnfkdOdPw3tiTSuc5scIv/kldpkFxSb5BWY
LuazztkoZysndUuoCSz/22CUvtonGNf7D9YYC0tAsjNdYiIBk8HHXKevMll6DmCH
Teyviv5gwiwX0270ATkpswIaj05PlNY87NHaYyJr27TcNhIcDM34tTZQXg/yie1H
4madJwfVGqeLLxomZcLl86+/c7vSxQBWk+OhBIQDACVTQ5MsKDBj+cT/uCYUXFQp
4xAAbQFN1A8fUadsVfB1Mzm1epfW3WW87InyGlawODvZN5uwrFz+ka8Pku3ACmpB
4obl2lbxCv0o5wjxAlrJTDfJiHHMqXd/3OkhZoYkcFw0I+dCpupaeHDnvK/j00KW
1r2ID2FxM1tw6RReABt6SNFsSYFMehuYCRWcE5bzzEfLz4Znvt7pHgFTUZ8Rgev0
bk4j+o11lttmEbpIF8/mMT1O6iCvMSnBCVEdE8vdiwcpQohtowB76xXpCPz6IgU1
1bv9LskSJpk5Jj1iLGuCRC9mR6s5wLpjAgvzZt7BFk7IGh/J9tZLUaS9o69zUmmD
+R9xt8l1EHAHmzK0RONzkoCuOuKf3pgr4DMFpvYugS021jlsg2N8lcvikcR+cPQ1
u6lpPTeDYdZw9+HOlfl+nOCrP0+pcptyiIuHESJUYlT5zw2f5EqJ4wURnbd7reuG
31pKAYdm8qdVBCIm2W307xVRr14H3g6ZfEoAfxVf6K5dqqTOnYBVwxDhHokq+Y2d
c1MK8aeIG7ausQlCx2If2Fhh9E+vmDLDoMnzjEuIvGJ7F9vKJw8cNBKRc1atVlrp
szBdZHwdTR9nEP3KtTLSu0I9rj7a7VMvB/ihCdGUqLOl1+jw+U0NqXBGdU2OA0B2
wA9FkTDbfEWkRi4sY5XQC48/Mga3pzrBLtUGe2Mq1P1ZxuY3a8+7uqCuIPOdlcco
YcNdYU71gVEjJ5WCEniOgDQ0BAWF+LIWJaWgQGBjB9KHdbLp0ih8D+4y63dtkKx5
2Ubpq4pqNTkshpn+U80GxuRUVS9vkE81lyIx0LqV8IrMivDtQkRn2WCwS2d7KmlI
+l0U14QNmb1bQgCbVpLU5/YTcpz1Rgtui9wsmbqx+aYpnSARgL1mq3vmHJymmo3R
DFtQ9g+eKqnFyg5LW07HsKi3gNwsH3kVXo3zviTPAKtOKT6e2caIWjtKdSu//cUz
x43PXNmYqwsy25wHPMAccOxeYvNMvRbcQQWaj23Zc63dgit1AyIcmbb0dnx9rS1/
6wIPZ9+QdzpoqeKSkgRb2c9Cg4XntfkM8urR8KqauSwtIDkV0W9Yt6OwSTIOFYrh
gfILLpjRtqImrELiO81w43HtZwG5R9AuIba4FBbz4EvdNU5Rwq1yjRX015DodY7Z
4WiRnA1Zm+s1A8Bf2Ib79bugfKkJEMEU8ifV7fdxNIjtmhrIgvFQ6vH1az8eIQvZ
lWR1KcJC4sGcY/VucixUBeHqScsBLImhYG17Mc4O7dtrNl5U2sXivmqkgob5/SdA
crLq4l5U6VLIQUp4tdoahoHKS4DswJyROQ9q/7XiGarNLmL/sh5v3mxk6EVwmJc9
ZInrqnOhtitT8LccseyOJU1tYDEh9aOTA+F9AyQ1pKMbozzzp/PbIXZd93bdHaAf
DsburhuZq0RD3lcmOloU6l2fi1K3RsmeB4jH9cCYaCCZlt1Ppdb0pklkf+9zFChR
sw5syMcquJfYP9ahV1aX5WGBcVNGcdlIuO36EQlXF9bUuRhZPgbPrtWcgNGxnHfW
v/bKTjmA6g9MMzCLBNqKt5aPOMT9MfSCkTP3bGslTKEriBWaxi0jrAoO4q/IlvZo
VnP9xt5hqt0OKLAiZwEU60xT/V3ACKjqH8zNxDSFSR24laTYkjJEPyXQ0jzvQkta
lH6QiSggxoqIKUq+TsNUIJfaPIRUdSMsCUEwwO6vAMcZsZdPoPg0MvM40u4HzgyK
uvsArect8WwreYtLzXbBdqG9rx8dcFzyDpmMHpz1ckSUtMpISpry/F2+YtRWwoGO
5NPdXGGHLPNEP1hvTNqWk4d/NgoXx2khc0hbvfw73nczyomAdSUWsk9xNIUl6tXV
ojsKFV719TuMVMjzB2Yvv/n/Jnsky3uMQSpK/rLwDSHWI/wL0+wBa7+nKDDlcsa4
vSDkiZ25PXVa/yp2uKq3pJO0uIlIQ1m/ge02WIQeR5T2D+7cdyyavCGYrYkSjMVt
oh7KPQrKMQysRMesTlesLTiXYNuu54pTYGHwODosJGbARv0YaUJzo+SQrrLlMOoV
vfEtaCSxBAut4oR16po3p2guzKATGpQVuSFOOfGtOw8DqR1EUjpgXlrz1MNUP0sV
fPXi7C80+Lf74F0turPmi2zpziK8Q1WuJ8fTsYeN3xMNkjLTdZpfVTwT7WqebfEE
T7Jucac2MMDAW4KsjGwQF0JzCGdKJkNlIR/EmH/uMiu4S8OIn7ojrCKL6x2uNxfX
VIy6UsAVsph11sBnRNIsZi7Hxd8S0pwKer2nMKtJNe1G9Xfxp4xsNLGm0VF6c4lA
D49YrgIi3ALGwlnNQzI4dklEMKOZmMm0j2k3e4Vz+r4qBM4sYPxrlfZKsGK5GH+T
iGjVcdk04WYBo3jc+NuRpbFddULP4j4Y5JSV/UXgHqoz0JteJ0a3VQo5l37LKkPF
j8xaLJJJYGXBHTmR38nzzadqfPoEy0odcaeRzjeiuf27yLx1w/OlDRPV0/PWU/zY
BW9Urzt293dH5TaSO60aVrN/goDZEnCxjPHbFC+t7MIrvops7/TM9Sev501tfXMy
gBQdpsLwbAkjliB7mJRIzHu5PZYSUsKftYSvFOIfLn57UM8x2pO/IJAQN+vyxzLT
lpRMRGUrfAys1Q4wGrzb6q/VyV9AcmGqQHHiPdQcO7YoWjxSY7ffpMjpfJYBTgth
jFYk8N6OJQOmnz+FCtQoG0oQfDgRMnNyBShjRrzj7ku1EJh6bNWeSS+ixBPTm7z3
L+2LWkoohTR33mZ4BLz49LZNfojzR9Ag2snKOCBImKGTGxk6mP4a/eOb6k4zDuGd
yO36M/dmaRdh4iddVXK5MmsC+g2p8QEozQeGFJT9rTi7JXElLNmQLeBWvImCHzTp
vd5eqRlqzxW/j0/e2lI8A9a4E+xve+y1pndi997UfpYwNqArfP7xqikxwP0eonBX
/bEycP2lIxbWKozNDyI5Po1Xsfa778dHtyXe2/dSRGyPaH9UkfF8blPD7fyjIRUr
NbbV/Xtx9RZWRv7TrQqHfH6ADDEWEvMot5ddEx+RGmd5cCikYc7bDbPeksq76HGh
X2t62jbKy4dL0nWMq9anDgtyqSBW8Y7edx0EpAiyPRJfxZfzV4ocorO9Qhecjd7K
Jc/1X3vFc1jkzepyKfIxAiyj6ajwH5f5qJcdYNUYouf5/+/lHw7XbN+tkIv7tVjx
WvMfhk5ZxkuFQdwUvsn7qIdFLtaOZWqE7WPvxjj9B8Ek0tK8hzGbbuMOElyvVAk8
zLuCBE7JOWBfwlhqms8v22XnoYO7Hrj8vReX19dJFSkSKJBnyy6jxuEIhSENRV1Q
b2bQ4z829WBsWT2w5HTJlbTkyHG5iErhnGE99c8I2t/A7/rsqvsjCqtRbNUtKbeX
Ofr4nPujvhvgLyv6EJwSBbBxzCGkyrmBL7BwYFN+Q9IzhDaDBgEArrtTaQnXOpb2
HX8chCPrKRvY594BKGIzLJL1ZyPVrgiD+sX5weNC+XaUygK+3ttT0L7dw9ggku9O
yjPPvStgR1wv25sMTfw71xyT/pRGZWvP634xH0uKBPA0zIAsgJa/0+eSWxOiU7H4
nJ6zwBH+RjiPpEEW24z7H9F9WpWuCKIzIUTfE9C6QcS7lh3h2S6vmfvSQLvomlUx
ZipzG54xJFkW0sI2d7k2ybGlzjOzwxDJXOn8Wn+vM5QD+DzR6B8hzBOWQ7A8ExPO
QvzuLr5SB2fUUTG1poqU1G23FvQ2EPH91yfgAxLx3MunUtSgAX9p+ytNx2w/XgWk
aIixZgKS5N3JuKf5crNVWFUXxwI/HvcUI9FR6V+OBfQ7DkLCfCDwJSP6qeLMfEXc
O3j2v0azmpt00QaIeCVi6f+DyDqp1089ga6/Gjstty2akkLJ7z4+hT+J8Sv4arL2
E3NGuKP2O5jcNoDBCde2NDkUzevg7itqt58GnuohKnTmvc7WZVGehy4pUweQNCf/
x9CRmLJSfovgOi5APkDE0LhAbvNmJREsQ6aKhZyytYaNC9cBiZVZdj/DIPMLZpwA
p0JDK23sMoGe1mEf5+DqC1RYSBJS+KW1mXTtLDXYLp6O0lzCwOxRrDIYRn3fy9eg
S23lP7qrKmzguow58iv5IYJsg2Hk4+iik/pOeHdsI9xIS8ikYy3dQLv1eTQwLypc
u1LDBjAMcdNvIVrvOowXLnzXYzXhkZ+Y5Yi/CJRCeAIKrube0/f4u/4Qh/SFzVCD
lmhEK57Bi32vDuwE9WB7r4qoYKEZPO6vU4aR8JmyaW3LQFAx9EQLtNp02Orq/gVz
`pragma protect end_protected
