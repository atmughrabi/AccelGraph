// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cu46qdG5VPpCk8wT/iDp72+QDavf8Tfos9NPNcoJQ2ce11sO4CxVO7OVydzoA0dn
oQOJCmGAQYndu16UicXUMOGvkhLBN2umjriV00Q4/Yn7g5lUO5lqnnMOgXwH1Ewv
DO31g3ALmXyz+Tu+P4UmkIz+5/hWsdj7JU4oG/IjLRw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19584)
M5iRjc2GWZinqNogYQsDZ/LiQiK3FdCv+s+Mr7sh1VMiqfTtdE5Kvr3ilH44b5ot
C9raiiF5ikcVmxnJyZvBoxUQ9cabf61+G7rBLnadQJvwkcsyr0gQJvE9EHsvPW/5
YwzfJsg1apV6GMOJR2tCHkWq1KddDTR55vvf3koxvA0VWAbLONmDaCjhczD6yOcg
MEgEMLfJd06aHmiHGYhyT9Lm8pRzl4PwATm6bUq7HRk6AKOi1DWwdosyqzNVvsAh
2VzKgtwTL5+009gz2cXRadFfDh7tsfnLElF9dawO+ZLZkC2FJPiA+HRIo4Fmmsc8
497HY+i13gGthvZVCfz1MItTtG6eLd2vZ5rUwRNTAthubWZLgnQflNDpPl+zA4Ul
3G5RmOGJzgQHKHNrXqjjAU0Lvext7uOXYjtW239bxcCWhdMcJcnM5dj/zcY9Jkly
grGAQHcnKLQP8GWBm+DnExxcNc4j4B7Ja1nwwbClZETSZvvDmv7yOPsfs0C5jOOP
0EycdGCdXCvdoi8QuIFbXtqFK6gFsUYaIVtd+WkyPnPTtOS8lOTPr0uCz4nupQve
zrjU+0UVtwI/JG93/gmhqCl9p9LkUfw4VWqCUtyTv0h846WvEcYoIGg5ovF9mVbY
PMuQ4rd3Dmiqk4YSJPLTx5JNvBuLUFWIFkKzqfrCRC+dgnaK90DYsQytnt76ghmS
Yy+W/DLR9tZ8m2lX21EDQif+ClA9I6hVWzNR5yogvosafLatoHknKP+PwglBzyUa
nJ1m73sipN5RW/aQ/0jelRAEcWIKknu8V0kO1iBGyo5jnLbOL6QvfA1YdvtoXWIF
oz94DIDxLPFskRwEXNGlStsr2YEV9N7880jnw5/hvg/QWwuxsTHvH4MPGdC650GQ
sVBJrnBe16xFNicIY37GRU+KunImyif8JJLzE7CL5OTY50DPO7o/6Hl1d9XktIwz
0Nm9f3pwgzUFFWaQsTtyp092LyW6m7xXv0U332z66tosqSEixs91YRnJgkgmTZqQ
CH7i2kQRJus3Ka3e1Kx07F30Q9aK9kIsCJV1twe0plcp7+One66CtIh3JaSBokmp
P3PwxH5wwZSjZ/5JkyTuWfhRhKl6o812LtCBJ6qqstp5tDQovlq/1lhG5QIYoiSJ
zPN9XJs891qC7K3wFaODUS/QAD7d5M4MwAr/ID3MNW5bItoiT0jsJc0jOh+xpQTy
yQ/z/XpzvzflaQjuu2efD5RKlljwKXA+UBEofeTbtxAXMMov+/hWlkWe+4J4q5Hc
39iYzS5eSPCBtPYMCLfSixsWg/8reFiVdUMIChYEsaxZJn16dXFKkrQdpMyeGCiE
DDZCsEV6G1ESW90KQTfAYN5nK3DWxIO75ABPW2vex1MAQUkYE6mI1+vON8xVtgSl
74VsD4ppgGXRmk8ETiGHbtUU1nXsMEik8o8GCz8IaWwSPhcpgRr1awhtFStx/NzQ
OvMYLV1ruc+iaASlJsFqjHm4VtMe4k0552+hSyr1euhqLYK1xTjukPfOGcHlzKpN
gy7NmRIzAbcpifSyxPGM/wSsRx4JkVV7NBvALd0tEK72XZtr5R1zRMPLOx04B+AM
2NHsTnBZ+GguVTqTiKdlj2KEoeHUUJw/+2k9wcJVZMtSPShYpSXQeWzytGYmH8xW
oOuJY8F52DbefZnM3cypINYkjieWKXxuaUoQqjAdomtgMDbQeMgFcFJjmdFXdA0g
h6Wg7+tBko5uE8+LOamIHJuRccYqmg9H95NkJqaBC2kP8PiXMPB8otPxYeP/nuI7
C5bhSKBwIgcadT9h9VkvX9/p5LIZlzrR2VV6PnACzqHWIr3TR3qCFp68yAI43fPV
MBB1aNSZw4UzIx40RIwhdu64d6EQskZFcHjiY+LqVsjsA0rsjZaCb+tE/BGUlrh1
Jg70uqBeFLoGC9tMtQVou4MdKRj+exsIrk9KbLIj56I27dnYbNvXnrsFCUdd7m7T
QbSP05LhwTdyBT350Q5iaoN5iUBOEVM0CTPBUOotKoz2lb7MEWCoPzsaCJ1Xvluv
ujQzIsyEVm0S8KyRSUkYOsu9GCalXmFUUfDyLIWZuzbbmK6w2xGQa+DLrlQSL0Ny
CBY4WmN02l7egJ/3uK4B89VYpWQlVtCTS8HzaZ3Gdutpf4G29uXp8/Xu/nEPTniM
6vi7u0zsReqVMSZSFRon6MBXdR/EfCFdChLkZ8IZNnwAIM/YeIkh558pwxs8CsJW
bEr2PMDkl58QkGYZZ+gogLoNPwWoFchq+g4Uvb32kBc5yhZEnGWPnlXtDvUOaBaa
hn9DGTbdK3lOLuFPFD5DA1r/KCmZTVSu1hI4MakC34YBlO9U9z+/NKv3Xkt9BTrv
niSKQxxS8gfbFa7wO6JfOhoyMRD/0jC1fHo1NTjRj1yzpeGHCTRiUEhzaCnZNWfb
BdDuDe7o6FUQ3vScGkv5xGJrKiEa7c0cL2I5TDOX2HN7njYKwMz8UEqi3hiEPV3+
9OQFDnQVikAG1GQ/HaPXmtLsJGTGgcJOMv6MQZYBeHC8cG++5vMlmDdiyq7zLdv1
IEMNIpiWN0Ub6BZ6///Rt0q9dizBPLeB9gbR+SXzzyLRPKBmPQL+QvFxulBFGmdc
Pt+mvZmKlYmOdI0F5RyfO0Etkf7BqbzDUPl+0FzPxWWz1lgQ+wIMSqEuVlIa6wgd
fC3pVKvtDzxswcRQLREbGeadznC8zfaJUD46Ry/ZljRTwwwO1uJQLkC4KVfNgzbs
x/IiEzbtm5ZC1/dB+VcN/jM3HE6cz+fO/xfkrNibsG6rB2tJkuTAml/P+cnurgRV
KGE+cByIE8B1uEaKR8pzG7UNFhZPUZYZnPB/tKHDKgeyeavD4/3c9DjLQ8k+2tXq
yOZtyeZoFfoZaWvQ6ZdoKIDFhvefanE5WUEPF2UzXK40Qa5+Bbre0YNpUU+KUpzz
OBRViF9/gtiK0vFGJudTbxbeNS5pRRNID6TsojivAtbOXg0O+Oj2/kLYza9tJWJp
zxH7AUHJdy3H7FTnf9qQUAvqtcRkv4MyCNQHAr+0Lk8evve9fQF46OTwk+uVg9wP
0pPAE3ysd04+LLKY4c5SfmRROAkif+CGnTbjqPFNs+uQIODMGMXOCoP95ou3JVVU
/XYwx3SsG39LtXt9JHN9jtYO0PPvXoTw3VzOp14cuX0dFgjH2uhzQQVXH89Jggp2
69XFcMmticYxG9YMWvSbjZB0aYyCSwqmnl0wcQPUZBb7KHAT3UEIDXsrJS04/F7u
OHw6HL8H4IhzofQ/SKUNYQtEkhUnmBa09aQGQNiujqVvYvYXzm9OgfCEUa6o4zfT
kQgRMFZpcCsAlqHQmwN8EvAWc4aYGbO1ljnlJW4Cq+Fj16l31TYuY6FqR9ovpVNm
etf5WDHCOxM3m8aJJQWalYg4KE4sgzH1mq63asMlxmAp+ZPXNkR2IHoA82kVrx8T
tVXIYN5sFoq5VQZORFCUd0W55FfBNbSgOQMAdONxzlM2IsYkQk97c9Pygw7Crx/p
J0wLRr9Q4AAAOQrN7i25m8opK8xKCCqGKoRYR4mG3XmAF8i7tJwgyQ9EFLD6f1va
GvfIRlnUR2xMCOl+AeEXYCTb+8QhhGralKfVzw0Msey8ZMehg1rRWOe7ZBHbXvDA
z1y2LPd1BabYeozELOZ/lDkiuJU5qgXJm+VnzQpsbHqfDOV+/0fDFuFsoeHw2qeG
S5Ra5ZOfYofITlz6oE4HEwT+45qbCgSBFtjVKNMjj3U+2S83psQjOa1xf1kr8WDG
zcSMOwSMn6GfA5LBrSLEc0zWcMog+i8BzjHYHeTViu0I93KR/Gf1uHCLb3LZFB0Q
5mbqoysElbp+zjwzVFgQylbgW5TGSxAIm5D958fkpgtcmsrmmkT5drb53pEj03IW
7q+iPYNE6jvLuuNNB6Xhe9OI3sF6cubTG+8+GWnSwSGnHHxSB2donWoWwq3MkX1P
KS2cXQHb5sAq5BV0TsU+h5DKt/WK/aAyDlQFTfLNRVtmuuXeji0zXJE3dWLQ6n1l
5tIV5bga7iRPYBTWIMcZU2fFBXwS16EJ6Kz62eL/tog/DUUwLMAVKN1RPcm7zM/4
ogSOfnamIErYktS/yuJhRR7fx8SbKxomX4eRrYVKTeEs/60S/YYY67nRBFYgBAoA
hTFvBPZNYmCbVQKwQZzlCGX1it1uoLkU3XjEeAkzG6KY+4VLL9QLAE1grzIVbebv
FDMHwAB9t4w+SiEgPVdWu0cL6dQBLAjxtV1FmBfAdlM5D7rmowwJmw0OvIN1F8pc
t4FsdZWABVKuRASjm5+u3OCSVGJ0VHiNy2jgMPsxole2nNLTtzAafyRqiy+RiIAw
QVIhR0KlBKdv44KoPnqbbkDXncn/xNglDp9WKRRl5Go8mYZUBCQyHlGfSHQCrLeA
dVt7E4ssbtkrULsylI6LdxsHX9GBUdS9Bp/wg9I28oslGVTc5IioE85i4/hebOfu
35f6BVVyNsk1MaWOIds+fy58YFKEs+liK4wewuHgAIjodMCD4A8aSIYhRjTZCHyi
hasiJs6ettHaXUgOKDkobYjYoZ37gnR7rAHuQ2G/c52WP2K6KoPcdMpeTnDrHlJC
6vBijbVtpGWDJt1xYcu2rUmsuE86KjBWDRB02KIhnZ7J046Y+9Cq8dydesRPy1wE
O44/ZxYneXEDHwr76IEAHuK82p4epzrIFzzWNvezM/1abHIJb0+ymLU0y8Krtm5m
YSibVMyWn/ZM/u2KS62JbJINHqcZrs/iymiLPYhiMAgunqw8HH1PL7rKOSyTzroh
AQnLQuRMpLO4MtzGkhoc/efu/ZvlVRi64ufsPP7BjoqKwi0Cndxq4eTkif1AKRyk
FkbfJXhfqEcQgRNlOcuRFgCDQWpjE1hQ5+7rgeytDYsVJyn77rM8hTYRhqbcgpfe
3I+JZwCargVJ7aXMKTRbL/gw8mwwF9KrJtUzAPGyaN00WjCdeANuwq8Ol4F5tFdS
nWxvV8YDoQvI7CiEWw124HWOtZy6EUdRWO2PLA/pUyo1PmP90NClMgj8whRE8RSm
I9BHTAEzu8xvzXMzttMiTdx+OSEWzIXcPl9C89HnEqHSCPik4t4aVLmwMlzz67cx
w5kUi6H3OJq0KLg+JIbis9JEsMD0eIf1tkA6N7lpGwJm1s3ntuFFPJDg+OBOPCif
LQ8egfOwIeM5aYH23IdunDTG3aLFRwcoMgoD92EUvpr/HmE6uKP//4WLVzzug9Fm
VWzRldryHUlkI9Ftc64nry/zOApN+8R2/eivvJOHCBkgHe0Kg3b1huZsovsC62cN
f6Lbq8YiZStlVBmtjf36tUvBfDge6C06QcrL9BIfpbUdh0D580c+ifqcQz2IrFIv
KXcSZFNMNaAtg2eAuvL0do9sL4I362SYz38fcK/BcFcWjG31WHDtsjzF4INxDPB3
YLJnbDqLjhcsfah141GigSd8R50MsmOEsz8JmMYcO9bwGCZiaaXm+dWsCxrs91Pv
KIOZEd5SD1RY39lfFW0WQmlpBTvTLhdzbDCzPYKiy9/kXtJGLXlmoJa984UbXR5C
O4GZ6/Iuj4PoucJv/eZ3FEKstq6dz6Jw6j7eK6qJxICGE6ia3qEJFXgWKcaui5NH
mC1oqyDvOMGpst0UfkSUcCejsfW3wkLm6TGn/4AAow72Hz7sTFw2nMBf0zeA+AAk
Shh9aSk3BFv97AkJFTFv+wtyEeEps4ugxZ8OQNPE9yGFttZawy9WoGGhwHhsh5x1
jLL4ANAZW024rSWEIWTNSwe63MNstmETGM5b/ib9Isq89XoDZ2lfluDFXTaDJcEx
4jlPaXhrREzl934W8KjCAdkKPHuvm+GhkP8yLB00avFWGiY/+3w5RA4AofTHcq0k
wyMeaTwCxvtvd+BDoI3DNMh/061xK580qpK5CSHp/HWyGp99XvrR3BKK52HeNg6m
jXsc4EsyhjqCH7bR91icQhqgfTSftVY3lmA6YENs7YbRy0SebEVw4AMDX5pLPel9
Mjz25w61vYnbvrJK2nNtW+4Iz+axU+FeWyqtapfsG0z+7aNjhvr3cY1xw0nlmLhd
mRZ35mDFT0mGKtKHa7A0qAoMl9ZHeU4XETHv4orNutBzmWqiYH5FTWT9HrNBJDUv
HoGrQcAqoxNgSpyekPkPuv0KAMx2aBMw5XRnKOcCGoh1UOPAihKVSKc8mQY9fbQA
XCWFbQYZdkAcFvc0Sk8TbdyxdTzw8uGafgR+CCu84FdME73z0d/geFgqhYqQds8o
z3U6xd2e8jbVjs9zcvf9L6DgU6ikkwGzCIDukgJvfw5LFcpRtWynnCW3GUk/eBP3
+QySYbf9Dkw9Pbyxw9Vm5tsad6E7+l0MJHsYlewzHgexQOFc0xX5E3+KVSUQJlyb
zJAT6wN062UNWkNtbpHWeiAKVYxWxEJ4zssuWqDr42e3EjFlR6L/+wcFqNB+beIw
kGagD22VcU1xVheIq5V46v4T3ZnRSOfTQB4EP56MGAiwCBIPsMi0VySp66NPYclC
E1tkqSTKTd2A102nFFT9GimkVUcQo1+VtKR/9Dg2COzl/2aP1PBP7BTMWEAh8Dnt
hrwENFyEEQCRLzsTFIx4iAYROP9DfnlnjmprGisr0UxOyPvGyr0xsrB1dHwaw4rI
lEF+AWw42F6tak0vgZ1uaWHLP57XltjmkErhMjREJybSFINl/Y+7iLOgszi5jTzs
jLJtsEBg6rNdLmjDcS9RbxEX1esV334A8MBCqWz/MPHyhN5UPu1atUsKj4zANC/I
opEDnHP8lZvIY4Tj+pA/le7tjUwEYZi0hX5RXXHionhRtl8vCMc7M6VSWcvBRE5r
F14Qyp++KHTsy4NQ3u9ZbirxOsPPr3NLlOAiMmTEPqkcuYy1ADFljgN6EUSHud8+
b5MnNLq5d7MS8ycIfoizV4reRRpGjXDZd6IKVr8BDS/vvlIj83R4cwBxrpDY7WYz
jIW+GFQ8xfmSix0ArNze9gyNJpVI0lwZq9sLPdFjKZGyoFd7WanhNLZxlIOFlziv
smNn4FhvT9npiVUD6ju6DcgGQ7Zre3nGuAjdFIfBl6yu671TS8TI9MrLGEguqK9s
TUrzWVfzY1S4cM7cpZLgkIPRuEPVVuk7oO8d6oDQN250hLPiY3i2NjotSuAqqXCK
N+iLKmgAGXjDpCNPoxwSL1ypUKA2AQCKinoLV1gsAclZSEjExCoyyicq0waiwtsb
m0rXcMKX3DOQJasZSbBd151WTBdnrb1vefYNimWovD/bkKT+E2F63fYlQDvodGJa
LpAil5kThzlPHKIWNQ16CEeNiPoYptkuDTEFIDN6vA1NaCM57dJ8KAtf0X0+CKUm
DBCgQo3SpelWceD6Qrnm2MNKV/cuI2iL0E+8EbHk8h6jm9ATE6g2oKAIOZPmMiad
0L0q9LY4mb2Q1sz4pW1iXlvL4vT7QjwUgO5QXPZeLq9eSZKUd+Tfhzn3vZbRwZUp
mFrKzVnwAjAPTu0AK+uLBK9lrT6BdNVmTF2T3ZIMzyltp/udFv96R3IoFmmgiYTR
1447WW5+XKRDiYQEss0Qt6LnIZSHXF3HpZQjyPeawq7gJ1P/outdW/otLpZxFY2Z
2uExTAjiMEaYHSEfCLlpRFQKU1wPcOqMKdaSYv8PJx0C0X0VCWY1dIAncog0Rss8
pyKufNSs8mF8w45CZFIw673rHPJEeK0GkU9oOGungZCjmeYgn/BX9Fae1S2l+D/P
oHD9ubb+oi7bVL0Wl4KXHZBtKsIQoGLoof/SjbGSUQHN2fIpSwLmz22xCCDxxoxK
dtJfLIR/Lth7Q/kHPLdHrRo/OFE3/a7FMYj6dGWqWSKKjsh2kgEjQ3+I7IQybpI0
viWBDRlB1sQwaJHbuFQeSokBsmLegI9O6XcyFhgtZy0E5BAjsbBqak4qFMAl/nrp
M+6BjrLZaAmKxet2gcQ2+ZoWOQA+jiuv6laGJfmFJoMHzPmaICdzjgdujSKdf2i7
8oZsMSm9XdL/NJc+sWy2aQUZrdBoRyw26y7OqbMaN8T2ayQpojWRDadsfZ0jcj6E
9YrqHMsPjDjl+uaPxuqjttgIRfpNcrc2VtJtpCbyu3V78DkpSersYyjttVwZLFkf
VvuKlm44qSZoROKv6onEFetyfmWolcthgNlgSB/PVVbx1bB3yF1qwk/EUr7pVBM+
+KryCuZMvoF24NFBwcjGztki1f1aV3RJ6zA6gwnK/0u/yYeMHfhbqFfqlfaeF1ea
jSocLLPkQ6IIIbjAlgQrXC1rzLOJa59nT/2LL/Jq6EqthfFMU0z0uEAvFKtOiz1x
wYoH8rQR/e+tVzazeq4v8NRXyRXnmxMIFqgk1KqyLV4rC2axugBAqEqyz65yIaDW
kvIzmQy66g9GyYEfJnFXjmkLWCuZ+yH5JRbuAznzQIMcK/zP20MXbLpTjNKHn+q/
RDXL1OxtxvHqeQY//0Xw1dz2c0l9rdrpwUl83gtiltp55sAR+Hmu8JmxJT+Fsuu2
ulnWcIdshrx4oHqG1IEgUccilMSF5GCOhLB78aaoKUPRcCFl+dG0Fk4mHASq9b+0
+tvrD769Q655E4+KmozUwIAzr4lyk1WzOOSLSDnsEJjzkjhNFquKSvSGghbvm+L9
TEkOhNcqUFaelp8Islmx0k62CR/zU+wt38TIB/4+/f+GforjzoZo5O6ERB69K0I6
i5J9+z4LKavtIp5h6vdtfFGTap7PD1ZCWok1zswQdVjMR7ZoOC+q1TrquRTgqXVa
MktOPCGE9ghQGEo7CsPrb6axI2XeYViZcKO04+sijzU6tpE+n+Q8oIi8rCnzQ+hi
FyqE+7KRWg/cKFPWpeNEmYBhuNsDwpD3umBW71okvyPomb6OJNZGhejK8G4QWlSl
sKQory657dx7ZTsC3/FkXbz6wdpdPa8qcSQLZVdu8tgMZHoZ7CwJKqAOm1lH5f6j
aWymbswAP1Z801kHfMVAinT7wzrSwBvK+jrkwg2iaQhHzMeGLT48yZwDmLkEcZjC
qTAOe/kix+6+kB0GgaCN/o6KNx4Thi2K0rfVyYIYQ9BRdyPrRz1K1NuIm+wPBCac
FEMK88XBANIrJBONIlKG6qzVqsRz0Y7SlqgjvsR2hNtMmdkcsTZ2xpWkyWMCrFF7
2k3JLIBI9PWpYGLlUP0Nzv0NBrZZ3QItY5ppz+JbFxe7g1aLBEK/heh+hJlR47bg
1/HBUuZTuYbrtEvIWOwUw0dpHeNtbIVhHjmCqQkAscKpXC74BxwywnJSAHZkVXoU
F1iUVaM5obUywNVat0tOMynxT/pyIv/UG8PI62BmV0Et+OPW1vrWECpQPqQvDZD9
rSR+TLbkhNnSwlzYmQ+YP+40CLoXuqhdX1FmQ/U2HclkCdj6Le9Vx0Vx/TgY+Ak9
Q/0XEBPK85CwO7SNqu8dExzZKstQxcJuCEqDFKDgjg3AQKe3EOUd8QD9rdCDXYfb
+/BTSNcFRSYdVN/W7xdsG7Da7rbbAn3MJC+tQ66Hjc3SJkMWnNslCWUsPZbRfzKy
AuazpApBMVrfjAm0YCz0h6PHsfa/TC3xbWRQnYXx60o/6Tr8jQVZsgUEV7i5CojN
gPQv/uHe4upfO9CfgP8z80c/b7loJ/xHgyJC4d/4j+MUissx/tk/2nDdY8oHTDKQ
R7eDAYDCMXZgZOfxiVisI+J+5rpduWsSeuuyCqLCX2C+QgN7bx/xzEKEgSafKqpK
fkbHeE32cii1nHgqervtCRfyrmD47jI/GA3uSqkUhDzvOaMTYe2EDF5YJP70M383
UcXJRU0rLu1sXI4GvpxOQnsKa2KTm9Kn8uZNAA6udoJsbFWEgWrw7/zvlLKxR8lT
KCl+bIxdwfe0rBXDzNlAxwUK+NaaRYhFaTYWN/qdQqeNqzUVo2fS5491EWN1FeT8
LluFpviESFutlE8nUn11Dp2q8vlEOa4J34O/5SN7RdV6t8tAv78UForj2j48gHuN
t8l0lXpL8KsvGJLBafHtjkJ0NW3EG3uHnh3FPMhsREO8YpA65lFUQ4K7FdqvQnAQ
Y6joFdYQZO3Orohc+XH97t7X+GR6jHGYJsKbl6HSfdcpcIeH/ybTVQi+9nm2SSTI
HXNOuKoHOOWdqISLpg3J9Hn4GO0GrDK88DH2H3EHZ9Nr13oI5e9n8shbSBlFWY3e
MkRU/fo3yGWfj9JbA/7dz75Y2QJxRD/tVQ3+SesGKiXLnlrWi2s1C8ARa6c1B26l
bWKIgmnJOeOng49UkMvm2wTmSwEsz4GHskiINk5HOpbRgMQgvPuZtKXjJx7PNm+g
cd83XjymkuAbmSLchw0+ATu0oWGe7+JGY+rgO9TKSKenalcvjsIxgzi7sokAEtWb
zQ5nP6c7RfGaxxAC0B0lZZdfToSnwYCsrXnM9rkZ4bRLs2sFKRR0bRI2fYcx2qq/
QcvxiUbLrrmuMiAYUyqokVsmqSDI6XSBiyuaEcTmpE86ZJ8z2h7RGlPsn2dsJDZP
86fx6TrZHKpatJaODMi7gSU5+M4Ye6umFvs/Xxp2d+xy7UTtspbsP7gqNwb4wwtg
VvwGkParTt0cvClewgVGKFni1Z+GUjg3RvHOaXzq1Lxkb6VuqbWCkYWZXuBFZWqa
5CgKt9d4eEyW6+O8v/ypjyNZQXfbgAz395r2K70NgJcL+Zpp86Z8wnPL1W+zk61d
3QWPlTmASgZDSehO2KibhL/InCRB/hQ56Qrf51/8MD9bg4lkZEHp71SUlUKH2/74
WRT1BYVsVCTs9uX/BFPNCU5EZXY7P0p2PxldaV29zFg89jjOjLfhzN+qSN8G6H7r
GAGjaL6+S0fjrxB3na9sILXFkvP5NjUfBjoUUt32gvKyLlUIlOzIvkCpimwuX4HQ
yv5vcZEm3fNcsqstExIbkBx1gBEVaZNi/c0ih0S8dJXQsibq+a3ZjoXIs9AmifV6
Gww0RoMg+zYyinHCElkrdaI4q+3lb/oAe0MANTf3YYTZy8zRt6FWtOTGjmWHXTcr
4kDUeynIXro/RJVwUey9jrP2sQ7MOuqUqOJ/TeM75FvEWYHnQ6NtDbadQWXhq3oq
BBM84ZOpcwhr0TmeBdAZ2x1vZXySICzZ6tKyKxRGCeI+rqFttgQ9JXtPD96gmNAu
tLbiHEmxxjWoQ5xPXq0ZBcOoABIU2xEMMaSpLe41RIFrQnrZLE0rFZ7ZzOklBcfd
O7nZRl9U/8uJPCLQs2BRDIhkReOlCMduyRODroIMHPV10aScSJqftopahrVd30Gs
GqSa0PLpYN4WyQlDaxgJOn9gG/YAjOM9juaFNqsBtgReLqCi3ksFrX4MoNyUGhr1
Ab6/NmbdPbShmmpBkaw3qVa4VuBOaOtPKfSQQ1JwW7mmyVIQrQRFWY94SysMcuKC
a23AXtH3Dm5wE6tEFDW3oiH1LWSSr/EKqL098raEbso0ZEdfLxssCSFflyLdEueg
l+gK1+/Xq7C46qJgNXWwo4ZCMua9AnMez/A74M2nZRVZoF7rh9TM2crsrtHp2l/f
l1fC4BV47FAjln2JEN2aCUj+V70fxDtudUyD+SY1KRR8dl7kiuXAuTSD+CcVBofM
FhpYEpF1jMPXyMXU9q4DO5ExtROscw6LTXFH4ezurajlc9DB1qSwlgmM0wKum8Jh
sBvS8h7/ExY6tmJPTVZHQbCV6PKg/TafLfC95dwdnn5m48BOl62/xS8f7XTCSXFX
DVxl4/uqk7UJjhXnYheFFjNDmSawc8ELtqOd8VV3JEGxgvLwfb/UUMxLt16LHXkq
bbY36CDg72ibXRbtQ2+nISjNjbV+0AGRZLUX9rHIITOPC4GgKubhPHScrI7pubVX
BSZO1NSt0eFRSurWkFtxBzrhpNyR0kPdW4HBoVo1ra3uX78GdLI6T8Pc9nvi2Psv
DB8dHjgn6f7sFlhXdvdJqJhIu3xWqeeJZGn8r400QYUMdH4QhxdPnyeGciUq92ia
n/owKEW2ZrH+mWKpsfu37elFH5XaoNgcN7EYu7kQ/NIPym2JjJYmXQZbZmm0JSSs
89jL5vDrwHERHsyU1w7MqFuH5DiHK13QEBvMpOTxYOf9od14S1TjnpaeTBLXvh93
XyiGblH/NiXIsxd61nJRSf4HcOy7CMLtYfctoFDPC19kCWhmJe7+UptFF9AriaCw
4IJX+jfl603fiSljcVV/rlghqQ+Zu5LqJPnxc1yxspUNSu8aHilaENGvNRXaQrKu
DvtLtFWBJymg5V9uiQ951948bDmV5yVcS149FYjmpRal2lbn9Oz3m/JLTQE5Z9v2
Tetjobyk3FJS9GZz0llyRjBs1MAUv2fFMlb/0j1gqk+mJmmr1QduyQsVUrTXAb7H
tV0EeAa/Ajy0S0qEWIAHUc4u62fz8MKjZ9Kp42pgC0RiWqKQtGswkt4irJlH5v6t
dqKwYNpmfrEbbAeXEoqLmPi6F/858murRQ1zJjuanD1+zQpY9ZG9ao006TS20/wA
REPq50iS0axhY/ehM79KgKenTWvalwtA8DWX0zteyWe3EnqtkVv/jK93wuyK7GDt
CkFssFw+t4z1lo4s8eZzbbxyjFT8rSWiTFrr5p8kdmeDRbIXD0+/efAJfVebIWnE
ytVhJQnKotA2Js4YAnIm8pDCyVxfPxbZHJDyc+++d8XIQVtRMszQPxexxvR7NsdH
nQzWjnNhBfY0nFPL5uv8pF9bYY5N8ByHFZ6ODixQ6iPoWPF1rWbd9LYJ34EvjJZK
e01cUHZlHNX/+TR9wR/Fj3c66cdSnAMHF55baocuirbaQ453C5bPhrMN5Zrv7s4N
OKAaAc35e6g0uXc5NGVNpYqYU9r1aI5M74sKn45kxesj+juKCwjCjfoTWZDEPEC5
1Qitrt10nM7yDrbuNLuOIU04p11m60ZWSgYg5vFlGdJTQFu7kt+7oNNyS/rAK9JX
GsQOKSAhNXorcdZGnLNiPlJmpSx6oitwivAyUE03f/ch1XfCCbmXTwZQU719GGov
RSlBpc91ewLTnBaj1h78ATbPgc21DzdclL3HrSV8GCp3PrkSgAanzHIiYojFMkRw
RUlt5TN36NwQUEcqV2DLm6TbjBimHgI83GuEniwnTyfXp+ZJGVmXckYVemLa2QMm
LBaCbvjsI+DCutdX6HQT5TQ/Ad3MelqdoRet9Ck84rn6etrpcin8mSqfoW92eFW1
at47E1wQ+CY17x/Qneq4i2s99tTAiKkELzgUgHNUFca1kdaBWfia4oGlOPS7bnzA
utZ5tHswOMWeIC1lS75QE65S/A4beE/qFhtsQ0ock9cmJryQLpYV+W7ZMPl/bnSF
okJm/diOp4rqT40oUyJ6tcGcZN3mDZ7W1D6pW+tNjnLB84toGVVYl+327g+SJ0lM
Hb+tzd6GquRTJuS3CA+ANu5/akBWCWNq1WRJ5AiPFsauGNJgjJLE2Agl3P02bNNV
Qga4Ka5fsYORWB0/tagjl4SEczgU+mfLbfrCTExCTA4G2qKLJM3AQci1e/85dKwA
2CImanwEzCISBtWnjNTx8cPB9A1Zs3MssJhkj3ra6hHWoROdPizZelJymKWKMgG2
x5+woyK+vmhHhlo7EUc9H7DK3iAnFfvd14teQLJXAXsBP0ZJk1NKjTlq9H68VGbk
+SlS7yKL0/oqOT20yhcXhjqHU6UEEaOZ7qexyZfhF1fzEnzIog7wtTrTM3naSf/3
i/twgWLI8RT55Bpv80E6E86woZiHAeetldsGdltqH+eGm4ZOLub/47Lpol/nMieh
1ftQfiaaEu+pmwWuf/tja/h9jxzLXDsFJJHioawOrfz1+NM2LFIenkeDw1EApDCD
KACb2NMlKz8PswDVQr9pPdYl8XTD3VcRCg+BrmW/2poGuRvI264bcG8qR0/umDVu
IcBRMWG4d6d0KNAno/nsujbLtjH83znxxYkPCtuZhz8wQSh8nIf9szZAkE2pcThg
oQDflt3ytcZR/Ear3nlvRiK9GpwpovT83KEbe3XiUCMVT0CPZD0orYy+/CYxD3em
M5ZxT3VchymDoVEJbCCmCQH0k2Gi1u7TyskRHKf5jICX5UPxNNq8t1Z1ObE7PeaR
bnbHUZqMzmiLGdvtoUXMOvCQQaFNzH8wvFqFISg5WQkZ6DoDxDPU5BXNDwKJkT7d
Hf4x2fiQfr0vEm811ev/LWl0XskoFQbhcd7XxxGCvVMt6hP3rI85rfX2wu7AMiYq
pLkJY8kiTEKfRBbhZbfby0FDGV/5XeA5NigJgnnQfWsvOww/xa/3onJv/wa0yBwW
2elQeMNc8j6Q1iK9qf7TfhQPPIiyBNJKjV6ZzromOijVRLv/EwWr375YUXUGYkue
rTCvDlS9miG2TYCJKre2Fhw4fGv4k3zwPg7hzrAtVnn12dEtO52fH5+PfgV5zggz
Mhz6iB44cChKfM8rULx0QqA+5dtODCgEZv4oQaum0j/iVbOdLvU/HVWnm2w7DHeA
4jgIdWwGihqXZr6LNU/yG0OPIWoGSDGLa05LRHnjhzQIWKV/hzVxrfrVbB01rj9V
R8qKNSVijDLAhat9Jr3vEWVihcsgqDhj1Tc5jJMnxi99fqXxh9QwJZKlMXO0f318
5VjU7v/rKyjx/3Cv1o9R5Ie518Mo92vnlydDsY5L9rGcEXw4A6Rz0pnLfazGmMzr
iP20TkaHBUbYjb/aHrFxD1/sdgzNe2V6KGe8sCpEPXGAd3cmUv8yAXvSLZNXUpfm
CY7/xyPqnKysxm2Z28nPMRXEkEu5dPzQGxw4xdjc1GE2+pdveXS8GiRKi8FikgDy
z4am1moBkCKxZH5XdbwEk+Hw2SnCOaTPtFb+PBq6gH9soAT+SoNVgOyo0EpE6L02
OBaiYO0YluEfeqe30xL7N7EXE3qRBC9buPY7BMd0nZuPr6P6ansHjXayVUATCHq9
55o+DUnammKQXFrzb2d9bJZTVZ8W3vciQs1mCbhcsPK2/B2Gl0TbfQTkYSeRISHo
ltGqDon+bGBZOYGJTrAH2xJPsM+XiLuXkYqULdLcwOBltbXeLbl12Z+lEw+c0egV
dqtLoRpWdjT3b+tvYNoG1/H3Uj/6EJuP2pKGl5pPozdldAiJoiavH4ouNkjX+v9x
jK72VL13XZfsEnTBbRAwV4B1xG6FiLF2skTbgYkaKcgi8TnaX+TlL9tAvjF888An
pvdhlGbv4tDglVadre7Xd125o5E6kHa7ClpLyImcAUXEPL2XD1fniEiiGt1pzB0E
aGG2Iw6Zh51hIsAajxRYVg1BGNEad5ONyfdWhhc6KFPEbmDmfQl8iDL92EdHGiPf
pe1gFPksuuiouQAs9Mx7CDSK7zVMfSurRDiCJ6OHyCIppxkmgrUs/mNsSiSYON9k
jgyRTIzHHpeIll7dCNxv5KosmV262bZ9U3PE+KlxmikXd0n8Vawc+8oGJ7tRIjOR
AOKvBxFlDOM3j28ofGIK+WtQfZVMmGlre0J8H6RO6Yy0JRaJXfG/dI05AykyLCtM
yUS/hNuZVzFG+xu8ok528wmXoEsSOCeWnW3ga36pphO62wmLVsrhcnYq3Nb36rUn
OAoU7jwzP38KlPo4MH9iWIG+Ah9lyjqhCsX2mh1Tf4fkn1NLkSt/6gq9GoX/IqAM
lGLW1fZ/BfQXVFJP5yicqi6F4J98xautoWUwouk1qGbCywwzqCWIKxrk2sP6UF2c
nishCl4AOUCEPZEbD8ErKS93Ps+k7JOymjvlWLni8XGho003/zrztdFIUGWlWySw
ZO1PB5NXZ9XmfIGSmH1EXPMEQos0XtvtO5FhHY+wGYgB35b9a4Sv5Cl9PEt9yf7e
lYHtaTnN0IaZqHdNDXWsoaw1XxI7mDUNUCc9WH4Lhj3uFYfA+79KMLVFIC1mwp+J
ESwT82/aZeeu8rh9THjwT1WS8IRtcIdjKyEr4/O/oVUX1+SykY3zehO0DSNigKD9
ShcRB0yOz72wLss78EEMF3PbBj19TsuoVqrT3KWrUnc5cejxgpxmnf+jKtf5nAJR
Ga47yt0H1OyEkwcwxHfduQovmkvNwfzQCT3X/NKAG6ODUQ7iMPNdkE50G3IdLhdh
c8JnEkJREDCH+h68H4aaysigM9TDguhRUsI4xTJrmphGFOlElL3dKDn+NTGLSQAz
GLNg8V0i+12idkkJcCzvj1PkCkviYc6BGsb6cGMdHRrhSDR3RMPtf9pTxzrqYxXD
/pgIyqG3V2BRZQTcptqDF7KQfLPAzewNbs1gibGTHjXtIIC9EwppHe9c5zx9jLth
5jAHfeNkS+cYR9KtkKMLQ63l70yT7nAZuRrHpUQVrWO+jmvtt6ME7CMxDBZTd+8o
tTNqEnls4JdPSgim5qL+X5TSGxykO6H9YqrdcdpT5oQ+gzEIfXGLweaj7FtnTxwz
vwFZ7qUMsD/rk25IAqreEEEkLJZkov/WXyLpCX1uinLhq7tApIr+Qi/accN2tfBk
jE6qeDl/IOkKAjakZJllnh4o+JI5wM9pjjfDYWcXalOA0J2s8iG0kjJSDQry41Ny
kgqSj4SK9s05UXyrKPb9ozPcMZ8769L5pbm/NaXRk3p8o9Ms6Y0a/3e84z0nSVz/
RkVtwduFdZD1bzXt1imeu6OIELyf+SZMBwgMsg7d+njoahPYBVK6slJEPcExCCqe
sbAGmIWQ8+ZbTHEyWFzU5ZurHCcRxYJVomsXVdcQiD09IsI0s0H7EWApQZzsnX5K
750bkqJJo168vjoDjM00hiQ8f/J9FN1t37KeBjQUFc1ywZL2BedfiGJjkdhHg/Pu
CCI2rYQEZiDAgOLVGi3CtKp4IWf6b74Ljdn0iuBfEYpfNU/RtFM4exDGuEr1dCpd
yLvOR//x5YgKnjBDTEQm0E6OBxyxvrJk+WtX0Z81h7OXTnN/zkNEpB5elaLiL1Mf
whu/SkMMYaOVF3SinKomvJer87GmYLDo05urziob+pHEIIMXzZPsqDlfrWODxPZC
7xkPhIqt6cwl6L3aPP/5nY/w6fTrmv//8brUuh6StX3BJNzTSq9DiS3jZaIJykCA
wcmXqI1JrnO8TEWi+BXTHmMbYj1KOPybTJXH0dBWQvu1caOHVzh6pTX8GzAHHqs+
LBFVxElVTwX5yOZ6i1HCe14zrU1Q8syAuhcF0WfJrO6VY6hPzzYQxbUHKIOqIoEZ
HlDJqLtbPzkOQBN4PXFSZ66omgfX75AEeL/2LeSU/8nQQxclDhwxcs8uxsirIHq+
GDaV1KEP4PhrSZR0aeyJZtzAO8aYYs1wZExeZfJs/TqoF6F9J04yPHtc8DQQqLXA
wPZxMDbUcX7I7MEsBMmEC7NVDz1HtihVRf54ZQ1stz5znOTX2cbpTkolTlySljsl
Ui4WRoo4F1CZUEa3U1RATs8El+do2xzd3p9iaibnjA+PDTZB4q8+DLU1dG6A50Qe
UUVAK9eWZnkRoDT70t2oTkch1cihoi1lJW2At/mTeMywSUJYPnCAEbNRGvCPcBwt
WQ4tSSCQE/pZNBLH52C/Gb8cvoPdVwyJr6IvKUHYs2rrLHFLebAMQeVT36Nf4nY/
6IxhGizBcHmM6ecrSwxukovhi5Yn+uNo7YR8htZvVDNhVsOZEdB51pqsFnrB6EZh
d8SZHZ65LyYo8Pq7f49M75zaZkc6ADYu+4DyECzPSzfxd4oMsCUmQGyHYSXQOBg0
qe9OBnxQxLmYQTtE3Ade8801NyJLz96Nfn9oqf+u22tGf3SaG4APmyxCDlD05l6t
ZgiBIpjc/6vveXhU5xTCqnfqCX7zXuzbryf2AzLEo4zT76TDXJsCPzIL0So+rhRw
T6hLBkLeJz5TLj8Uh8HMFx1IQs3Fr0kHTFoJtt48AAkkV9PMh0wyNYwWNi1i9CwR
lpvBmW4GAA3Ruil7Z28c2CU4Y8a0ouWl/M6qwTnd9r81c2RuRSIMCkTOj3vT67ED
vC0JnEYm7mEikcQBrH38DUcjnaCwrFAStAqtYCnERLwf3vdXjUKotmXIZF+JXB8A
ltbO9cA5adkzLLRo88Q0IqFRiyRUNHYAdwqVdgaJMVOxc3NDELP1uO/d0RTN/Z+f
a3GAKVsUctxcau7QuWfNPL5VLsYyxYvQxketm6nvGag4ZxKWVhk8cq57dpZ6D/5N
Jf2M208SJsIszXUNC4mqotxbkJsbIq+wD210aP2ycq0wTBUlfAesGHrQig/CWunt
1y1Zw+UpvjFKUJo+YTFXbM323/ToTohtae+myGs9owr94juqaVxL6IdJj0QaeoxG
PrxPZ4g19fEIKK7QPWm7LGcskD+O+K9yBdzHkzoqB43Jz0JI1mEY7RymtPSFuIEq
GrUOo6KyC4+47WhYXZ4tsYuUXbZnzev9zLU3CcsMLCd8kNgIgPIIxCI0HYBe8EnH
rvmKJjusRe6t6U80lSYaJ0GK2gYLOfiW7nuy2N6X/1uREIIcBgDwbcpLvmPA1hy1
5VwFTc8LJhmA+ugKMrcueBfn4NoVqxkpTBDot7o33UHpbcWQEDFTcCnF5BIv0zyQ
wClPsaO46Jy1xz2ViwIorp5hZ3Yw50tEmSgWgo3/mRHn2l6Pr16reh9Ra/YKf6cF
YAO4c/6Zs9uJ/6stDq5phfqHSe0zfuhKcdnxbdR37wpXFXJaEQBdmVIus68a9jMb
FRYsUF9Gr1NwPPo6G63b2YNgVqeFdD+iA5UWV7wHVULeHB6PXjnFmcWsasfrYvuJ
0fS7tQ7fVSMYT/kA0mve82IntBqt2EsAUeK9QLOP5c2sdErdmRF7JLfhTmaldhVb
Jk1WcvBMXRyDzgAktfEFTHHse1S7jxL0fo9IlMBGADbc3nBrbLuzdh7fmjTAWaBz
KScLBmjtVxZeSJumepYLwMlx10X/6P0oHZGFzbAvVE1PvralrrnC2HT1V5kgc/Uq
eTmFQNhbuzheGFj73X6xOHTRtj7lCSNs233Uby6detFUtNezLWp+9qdXKZiInP1k
5B37w8B0cfEj0oCZKMIvCr2Rx4Vo9AfkeFTufv3ycon5OlhcNvhNWDAWaCX3Pa3y
97DcXOnjhNI2x2En/7nt+OThcqsDO9RDLE0QMkBXXO6ENoP7K1m4VP2vgkHFjRh7
gVPR0fQnXlIp6S2iw9aGvc7XbeNwhA7HdM67DoJ/YJbHJdkRVdDbuPxyGHAztGap
VFcvMFa5TZkXZzxlK1jvYOqtLyL7wbYSC64nZGzA3WNfA4b1qCFOkU4+1AJEYQHf
1i27ou3Ykb/ST1r35cqrec9S3o68eTRX8ugyCdnjxIzaNOHlPAgLA8yp76R83yze
8cRfsloHC/lRFBxZtTkZ8Pq2mE/DcJxw4cjEZn0pzHC075WGPWgNiN9Z6szkTVpr
oq/Rs22lwmMBTx+DJRL37nQp9R9N36ZZeUyUZhs1xo/ucdTjBhk8Ch8h+FHirZCH
aZCV4XE23OgFQJZDnjtSP9fFDEWBSaSrokneh9TtsK84YQZF4gRWZDWpZGvvmo0L
ZEwn9vEsKdgeHzGqe9ufDh928WO99gdtefhAliO2gtMz4TEhmMKBqlKYIBjvFe8v
vaq3v1yWQUWLiIszUDE0kEiCBu56ZfdRI/NvtQ1ADeWXWLngV0+ksI5MeWhQ5BkU
UZwD6iM3O6oCMr5uazBLz+AkztncKPd+Dn6/DqAciRKb3RtEg1xWYn3245oEKUrd
guakg7wK9cjDgTWXncdRRhnDLvmW4LmpmAAvhgMIKa7X6UyJhjlePA9gy2+a1Hta
ib8It4wSywOQC0sMGKTp3zHy8BQqgcqF/YWlAWgLb5tnTaJkhxG6raXYz6NlrKe/
pKuU/XDEfvK8lyUd1EkTYznqQE8H4rhs6Hp1+vOShLYY5gOxhD7YGssiI6aXwt2t
wgNvJNb9eSLAPbkF5oO5oLQdzrJERnlaNSJ3ot2Ye592tNG1yr2juy4eCZL5r/v6
aw033SFu1E7fOVLpg5HT8Bi5wbNE29cIj/ofpepRIrjzfQFSVBHZdPOLGvRFaK7Y
bTY6W+RtK/kj27I/fstrhJ7/cTaRg5t+R46cFz54F2+NvNJoHu8+8TjazUyihzcy
pmtKYRkK0WN353r2NB428fHUu7lWBRMQtpjjeUIaV5Ogiw9jpq7owBpmtVAW9fBV
yxtKzGOO8DupnGH5NKBidEW0pg6PoGCbtyHFbL0Uikl4rFn+zIfWpIxbR02eHEPq
JslHB0tR7o3D6+aU/kWjord+LBcGN4EoqAtNsL+0GGh11iEXKzQfPlW1vDSNxe3l
cDn4bnnwegzd5pYbSRoOKh/Bc6taY1LKg4Eisskc0c2+uzmmf8cmg0IC87lBMg0e
+g3Ae5JYAJ2/icVy356/BWqVebzXRD40ZWsiSWzeDIyuKbWzpiBvS0VUFuhF/NEV
i3UHiqaEswb5V0/lO0VhPSAUrZbFMM2GNqSZRRGIXOa7uZhufD+JE50j6UQW7bai
Th8Vl+OXOjCErJkcy6eTzQ5QwxDfxwMCTWBAYz3jhXM/yIdsj60S+WxcDxeHY9ss
beW5pr4M0HHztSKFOc3CiA+d80tgUWfU72toJv6DSeg74ElH6nEDhh9Wrs4nByIV
j+ot6DoGaCYhrL3mFndfQ3Y+GoOqjwL5UjDzg+xCLh8sUulXoS949Zmz4OcpH/Cm
HaUuwOYpZkp4Z+xXHMdhJumFyH0miTHo8Fb7/z6waH+1vD0akDIF7ijLFYtfWkP9
9Bys64Aar9AvWaYWplsrYH0qMXuZnOlW7t1+psoCLQKIu2XB1NJLPSULolrnuas3
Vwlqc4h+kbp2rw6ACcNDbZ08ev9da1/+u0jpxjjB33N9D+gXbG0GCMIopKA/Cwus
j/4MLE5JkZ2v+Hpz6qvd4i5It/IAildq8YUUe8N+zOfV+LT8mqNJJcqOrKsl17ZP
SfhGmBuS9qWzsMigAR1mS0QPrSg6rtpA1fsovXe4D5h6+c2jrcATXGyMIEU1aO4X
2NtTj/e8hd70X6HTCZ5dullnh78cjdV3LPfQNJxawid4xNg85dTN01bZycxIz4aO
9/aKFv4MGLlbK4oubUhLwJWpOgeCLt7EF3nIt42HvKlcPpRgbs/MGLmWHEURe0+2
NCA74uDCurgDaZfn5YWPglgwlZw9usADT8r1FeKZod74KiEwgU0eLWJQgsoQUAEn
50tacsWX9xixehelHiTxM/MNyDbbcpHfOSVDihKSonxrYb49E6+Gn8NeRSaezPSj
m6n4o7Bxq/qdXWDi+0e0KsQOqfedgaRmYnagsBukhUf+Wgl5cbmsuZB175Kyirwe
HhlEwlNLYPZcWXjvbnM+jNPNBZ4p0T/oEZywdKiG8r56Ete71lu4en1tKAV3bhi4
L8+UxbZxQPrE8ZusIoEMILVrHSf3VDlQHHlkZLqyFlcqsyP9knd3xJwoswg6Artu
J0zeWP1E5w0hZG0+yzyReON4fMdHZvcC9GECDPrIZmmZ+AztGCwD7CB6jB+vKCuo
UZIcXXrfOTv13czl0Ojcgwv948ForsttMGO8ATtCysuu+TbDs/G0L08apRgZRSwD
0O940VnB2Tw6o60yF01Y3B+pu0DWeLb+9fisxsA2EpkKG6DMGm6XvPdaU+hr2HQf
4Y9MAJlCPfMGR8BXJpy1OMayLniGYWe+lnagqJcBozZNzkfgUTZU4bMepfZFg9Qd
sYR2RBIgB1ktkdVcev0MYYv+VhV5zb5fbN8r/uzHrZdyr/wkUl/amfakVtuHTE9Z
CApDIllZ21cJKwzO+0YR5p5bHIY78KxmYoSE289EZISwDGOJQZD24LgyMC4BcKLm
X+Qga5SmSrq+5hmn7fQVIxLfnzYyWOEDMzu+P7vWgHKmjQnT5Id5HQ/LNu2scCg7
eW3BOXoe+YrxGST6r5Qcv1iloGIieG7p5/DFo0+81kYf6zCIT7egFUioyHzwrvZ7
pRRumR9R4QuXcLG+aDGL/RCztPlmoi1FG2da+tWOxU2BhPXDLMW//hG4zi5Dox8k
HWQPyAaDFlTVmPClcYYydTa9NPYLKgzq2xT7pTxtz2hQ+S45Z8Ff5PHjbYMvMRur
sBNOkksjl0A6bxtJ3RLbOUqNV7fng9l6cV5TGQAuCpNFiXLDPBKvZga8zpgh1D5N
RxlNDB5tso+Ozza/eQJw48vKSfmP+PLhb5vhJoVP1u4Nc5ffqh/SPZ+pPBmQGopZ
IPDV4EUeR3o5rDOrFmW8cO82sbuITpbqq/oPhrOq/q5jvqUTOOl6uFRzWURyrswE
hguDzmeeBhONWuJmVuu39HZ2Yohru7M1FwTUzczdOgP+G8DFD/WNMb6PEtgZ2gjk
L1sdGg8Du9MRGkahPC3Tns13WvWwUO1M4+PDwCS5gFT1PlQcw7qUvJ4N4DRQif+K
+OvAAU2ynHrhwMIeCLGHxSmn+flnS7oUphJX22NGDB1GszF0Abhu4d0ToXWs7VSb
C4jEVnIk2PToNSBA2x828idfdAHagvOhmQZbK3XuXtGSC/0jByJHayvShPnq95DA
pOROeGLTgJ6I+siSuzjN4HoOfv6Ddv1bhgD7ljdCqsJ+viXNJtL8ei3Uq5n87Iuw
od+atXmiNQhmtnD1WtZYtxDhkfjgGk7882jqMG25uxetrEbw4klVrjkc0X0x5MTc
b3oFj2J7fTK4G/Rab5C9Uwt0RvCicXXZH3IkEWjOE/H/GFkPUZxVAyWSqP2n7oxm
9mLfk57BPaaJ23JZkhtdpH20EnVkCdwUK/SmFvynP4cOAr7i3/Xa/RecXB/LSmCQ
GvLB/hW2bPFNL3d7374Dg5EUqPRJH/6O+HI65me7uU/1kiADqnNurWhtB0OV0Ump
wayF+1KwIS8R/NA/RRNbuuajLGGByTMuWrXMXYt19AMlE3SkclONjf3GP/7tsZXy
0TBdGSMHFtv/qfqF5Ee9pWLvzGz4aRdtWbyHEjWXXXhX5Rw9/J6IugOrBkMbHsT7
vzHQ6KM2ohoZVPNAPRbNA0GCnM9SIivf+D3YVdQDfXAAbdY2lEHQXwjzExrSh7Zf
E7Fm9ReFKPtl3afHJhE2N6OT7hhVqzSo88AjuCx3n44an4uM4sKucSB9pjYGh+wD
XtkGrJZUicl3+O1rGzLkZzHgNMi7NLC0ehCRr4YIC0ITZ9tb8262+lG5Zahx+UH3
pxGfc+UBgtCrDFn5iwuK73jYnSLDoeM8Tz7DChU/kW7aeLgPAT8TJsmhifN3A7n4
GkKE5WpeeQ5mkZ0d+iDfuktZhKlsh385iMowi5hVjiEBCyd1y7dPKznr79rdNeYY
feIcopyKDoJSym78G6PENaGIyExf0e91qbCbjHMbqG80SnUPda27b8hYJ8HCe/ei
oEmsTNXBhRpfg/lSxs3B6S5IohwXsaZ8RKuae1mD8IV9bMSGHhY+X0Z1MVpp76lR
0/6fUXgjUOptspA1mrWg28+bzBCkBsmr6GJMNzw8OFD/Jzrw/qG0eu2SOo8PrDXg
tL0vkomSs1wSltvjPCJ/ciJ5pbcyqd6erlpY/hvVaxkvKixLStZMCzIKkoftfgPU
Tt4/fZfWZcGQZxbYLQwkbzXU6qrSx/hYCltR2yWlrrTeGUG4NMK8j8833qrjB6A8
MEksPXMdBbGeBuNFBgB3Tzb0DSSJ4C2b++syD/b0OlMAnAecusDt6QLsdICi8x7J
t0NezXdC8Th6qBG9qrDFJMhy67KIcrE6IPZ+aMYihUJQ/QFqV91J/US0PRqDO6C1
/+oJY1WW6lwpDi4SZs5ELU+XsTm4YdtzMPyjJ1J41Dm/OE8ihlpcSkWyWnkPxrJm
D+MaWyabSNAixu+D4tc4d4wBV6opWdAfnum2MmQV8wF8mL/r5MfOCXiY/+DscGNc
5OqljYvfGKoabHXsFEOjMk9niFNoUS4Xgqe1G2/f18lvZ9uLiqxX6NnUYXQbJMrN
4CmxcpL8V85pF9FlEcm0+jpgb9FJrYRxVMTjQ9mq0c+aF/dlt4RQWJk7O+z28uzT
rky9GBfN2U7CqtkBS7Sx7SXAUlCl1Q15ySB3zuK9pvYfK4MN8OV5wr96+md4C22C
md45rF0tmbO7h0q3PjibXVIjOPzaer+gZEwHosghVvSKREj98oxtfep1+D7Cvb5D
cuwQ3b/ABhQfPoGbm5XkVD7FuHA2J7l48vxhKW6VGR2hr7HRYpm1rBzUmED+8o05
R2CewgT+AP/B42lJdj21KPcu5KtumCsis0NFEMGfsDEUCwoh538HrFfk8qTiQq5p
mTw/nUYi6doBfB3MJfuvuaNW1BUsimHfqMho1MLZu/UfDrJAQ0MTKAU5K9IxRgBL
bS+fAhIZ+LOLp7Digu/SHEulzdrWZu1Vedq9mp3eC96DC/mT2JdJhkwg3HaGY/Ao
b8/4mS0y7CqzcywrKdzmDAub5lcJI58woM6sHP8GSZJ+mysYE78tJ54P2sfvHfwQ
RxpaHdk9Mp3qH6TZb25/89MAQXzQC4BfTfgd3f2RGad3gvDgPKgNwKJk7cxqwAK7
eigp7nBHL6EcJ5syuccoTyGc9qeoMMYovY///GJITPEYSvedaSpAswJyNYwP2Otk
/nVH6RXpbVxp4E3412AovKh/xKKhypO+ptmscM44naEhMDtroHUKjVHUB0tQNxG7
CxxWK7hHWWYaB0QEDNlmooiwsLBJxlDrSi9bT76VKAvEnVGd5EZoO+4TwnctTW5r
81uemaF6JeSwVcmQdXgHvZdwt20PQfzM1drd3XvQ/fOiAuoBMbNsgT3vJuPpm/P8
0Ue0eHIvfl7gDzqQNX/QIFmtzdaeC6XBph+AER9Qsj+QomRyq1o+/oZDI+XJ2aKB
mzr8EwAfS0aNf/lrzNM0r/y+04NdUOrxxNvez3PY+YbHmhDaSGffEs9FumoPm4JZ
yGhLKBVFebwSeOXqLI2Y1rqn7Fbv/WA+pWhipNuEcjk5RktJCYpqc7U4mKgmvJLn
geK3qK17RGZNbIrg8k+tXanhpN6Q5SFWaMnlK4tlyIrtCU7fTKQJuzNutDc7rd1P
ZTm1lMC0rNf3ZVIM2K5KafCTDjTmioPf93BC1Mw+y5ff6bSpVI+ZCfs9qZCsU1ZU
UD9Z1kMHxSJB0r+qOtuAnD3hNEs3vYDqSFf8bHKi80s/JO7IGV5fsZfstL07QVRP
8+527Igs4+6wWXfIqGN1b55K0IagfHzyvVh3Z8Q5a1x9x7nq97B1VI01xN7yD8vj
n3rT4kMyLnML8uF9wOZriAPfXTWGGsNkRIJrautx1rATG0Iu1QVVHkw9Gh5M+WaJ
Vad5zWv2x9uZdMGKZYE84W5dBzAFZQ4Vg0SG6xAqCMphuETu0eSBUeDkTZBucQPk
nJKfgESvc3JQXwPBOb9kIwOlJZ/EuUvWRYTAohrz8CIDGbXkE2D/zS8+5deE0IUX
eGgwTNhC6Gj9MKrZVa/KWvXzmipZ8bV621ZzuEB7mJAu/8+/oaqfPIt7gcj/cFlZ
z8x2GbcYTd7Yin5fJLQtCUEFdK1z5+1m4XnTQ2sLFBwRu/rla+tcHX9e1yzjSjSp
fQXNhx0yZcJpfJOApehb0kBWDPuzBIniIVxlmUn72sMr4b9iJLDBpmXsnLiu/Lsm
DhFr83OBoatEe9R3sZN17CrkTxwUo9LfyEys7tjnD+xyqvejzOqModzcHa+b3pD6
Gs/UMcwgp+IX7jfKviGszbMJEbmFlUEKWN4q6GR2PozEGrxaD4MXm2xtMrC8S5BI
WriCdD5EgRGzFR5ucWsEdsnV8oWClP5YJzA8DeeW/LV6uchnaqft04BJu2b6eiTL
BsJ5E/yzYeYtMs+2Unep/EWEaWXPFih1JW5vN7rFQ1prtA4WaghabVrigTdnoeHO
Pkd1nEZqwu1I0B/6aMtaneCl6CSKHhPCwLUeqMVyifvMpHkK+6k4d7//kRvHj2ID
yWhJOkjfU2Abe8NUvVvONFrC82dFzhtFtkc0JXHck5YNnz1S8y+rWFyRriUAZ7SX
70erdN3pDmN+3cBGe2EWMgfF6di2BZCkb17WPTnk12zjlqHUl0zDyGdwE3139Drd
A2mj4JCQTdZFsSBlILoz41yTz1Tm8X8mGxWZgbwMpLpW5GP+sx31r4c2qd8kFCDo
9g0PxL170c5C6fe+fl2KYSDctq6yHE+XIbfRk0qFyNrc/+VLW6vnb3XruoVo4z+M
`pragma protect end_protected
