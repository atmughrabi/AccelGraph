// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iHueqkN//tn23Z3itp5bljZAqiDgEr6pf2DxutXegONix1tkv1+IDut8wMinwNqi
1KP4KnXjjWH5Q2GOx5opI/Zbwxg7Zq5a0KWhVzFK0iwzjEAQstWgB4j/BzJMDMeb
6Y+o3oYZROQ/TFuDzODVaBoYWJo9v37wiwNneXgwjtA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31808)
mG72W5WcMkxqP5GzEu5KwOEaJdqIhJ2SAHjbejhXZjokHWgD+C+nKBh3d0vyP6iw
Nd58xxlHmEczDRiCHISSdag9QICLMUcmKURJxJQ7WyDjPaMwB9JQNVfKd1Q9BipE
BJDf2S1d6b0ySBchMQHpEae1XX097StHNTuisGd711crnVpGuOFXuZ+bjTOpOYek
hIgdXtC4zsgdM3F+CuOBXjxSlbPU/OPCuWKiEZ3MRhn/WrQWYGqJIaqyZB7g6Irf
vA0NP++V/ZoAX4eUrNIkci+Ue49EEbLTImSebUCaa20C6Xz2YVnCrYRsjKi65Z4d
Y+Hg4EEND/wa/k/FW9+JndQciL+gWM7En4RsL+2klHUt2MRs+FT8BrrghDRgoN3C
0h86XNJoTps9qqfxLy8cxMn/MYXJilZZCG3HWH65bNcFjZysqDz+EO0M8vjvlewY
JsTvBsy/zwz9ay8YqZt3XQZzo6bG2nE5tCOcvpWsEUpUGQXcpMtEy+fwx0N809Wd
ZqC9a5ogL2esFrDwE3Q+nsYbBLZvpiRn4yiW7CHHeJpCEzPpINpEyFT7N2lMXCXk
UkG+RpXGYvJv9la8aP02HuX2yyRzzeEL/8fepP6D/tsjK0WKzOXyCVeOYTlLijdK
LSja1tTsf2y9tK9+JeTBFkNFI6Nhc8kZ26gSWAR5PMJCYJlLHb5v9f3ss6Tfhf8K
AclNiRDvx8gb8msZHYOZpr8RUVghYQBgiIcxSwxhx9flgUOKVgH238jn0RPY70z9
N6hzn6bbqJRFh88qVr/dS/cMRQx5qAqxdsENyRy/s2iy+d/7U/+1/YaUI5hkMKdL
sOX7e9ebxbGM73Lp7351jhVf+FgX5FoDBzYNszhual60xGOfM0OXDIxm0KPcGScN
ynF2GYDUMA/8iwso7QQJrUB6ZLdeKw+pXF0hkyKFsst341qV5ZoKADMqHb/uQyFq
GsluNfBFjfJjEGwKrZ+0IJEaZQ8/5vSxjhegx8itGRdMlnYYX/DuyHvUo6TaDFV7
8jSTTPMyR3OztFO2Qfv0m2WlVLD2leXZLOkud26vel4/IUnmN523mxqQv0dYVDzP
ec796NGZ920QwPi3crReVXFlWizOa3ThvwXQ08EjicK0bj5DyOmCdquMlq1wP/+F
dxB/nvMUqdzdpuB3qgp9rfAl7T4mRTX1FGcNvQjrzOchGheoQe9NA7MClNk7UB0G
HKF3w0/64oBZajNm1ElbDKNBHngI2bxi9FSLN75Wn5UMaGmqDLtm30Bs7FC/bczO
/DbJaQ/rRnjnOvV8NUGlT0oRC5+EL7kH36W1twoO14pz56VlY9h1Bn8sbBbPciRG
WZTiY9Zxk118OsTXGQXUZ4yVB68ckj4Vto7A8DWlwdzW/aXi0rBEZ1qlEaThaVNh
/imAvgJVAkl2nFzB4SDw4hIUxaT3756W2rgyuTbe0aij2+OR2/GWPDYRxR2lDmw4
KhhDB+KIeZ+8c5rKjQrQKJNKPUvAClisrSMI+B1iy9xwuiK007JcE4zQc1e38gJi
TZBCdGxI6GDbN7InNwLNK70feoL7aPXZV3ORlAr3is4AmxCbQybaarTBwzV8hMo6
4xH6zSWaXyFelk4XiQynXPFLi/u9Q4E2WTAPor2pJJg4YuhtRe+A19F1ihkXSIMB
OqqWhvBw0HplStxHrhTjOtkgNEpPHYIfF2vAZUgMxnXLnROcorFpO7Hq2motSnjf
IvY1Rb/5YslDDTspGEi/xxcGAyB6JGqKWWG3o5taGaFnQjOLPVUgsGscI/lkCzk5
dT5hVRAZ8HAI1lwQf1lUPul7JIkHq2ziHgiCsHrLtZk0O5cRd5KDUlM1hEFy+cS3
pDQdmGnOkn0KEzgwd6NXx0s5EGCAkiBs2wUIi5TdVEEs5LXM/sejeVwxKQMW5iUH
7lsHr852FMbNc7bL88qxIFItnvVZWkpH3g0NR7ms5Sz1g7h6f/Ea4kwagVlFruno
cHFGf5b2uwHuFqXYG4Unckrpii+pk0g/DtUWYXSFKNSzkzOKXHMKF/J907Tg5uIU
L1kWgJo1zhF80G6X0LpAnZ+M7CEV8PSv7N1kELCNnkQj2qGMA5EVgvQjZzchlW7B
EXmiWcYMT4zpZRP7f5Nj/n15rD3gyqyLCiUhIJ2Y9z8oeyia31ojU+pCVwTx9V0T
sVgHmUsawNfL3xrJtH3XHAiHi4iEwtbpaWLxVz1z3Al+bOIdDFFHuK8hiY7DGug+
11Zy5Mtfe3vNykVQKWITXWcRi77EBgOqratJ6nsQ2tdNNIKt/S6gVNE+iWfUUBDl
kKyeWrEFs9kYfjmejxgyC1zcdxBKyvQZpZM9KPmSiIDHk8/ld6sHBBglVUxzKyMi
3Dw5OkQTYdbLTSujcO4mPlworiBqRltEumUNHf3QrOlsvW/N6ywh16XZSy8/OPsc
DDCrEky809VccZw/FAavwLnAnfC4H9T4cuRXSD34B+Sb/lEryqJXgwj6nvgXAxvg
O9ivoWcGmWV/gHoQkh0Yogbn1ojiTd0XgRVr2nzjgsYAqhR1B2rBeLwz7GNdMfNV
bX/nQM5VyDOMLv1iC8o4u1G5lZR/vw7q2bo5+KNbbMsYKmQsWHUrlQ+9BeaPk7wk
Aa9DQ4Uce5PLKN8kHtYhacGtO+Pqj0fDJ71QJtZUuGJqI3iO8pk8QBSwDEklUATK
fJl2C2i4zAIYp/a5nokpBqorVMkk8uQH6S9ij8rcUnNUJpX4ZyvyYIcC6hXz0el3
J8OEcjQSfrmeEWZ5ECT1rcxztvhCFCU5Zvi7hHzwQldjt0eQl7mTFdTw70AXD7ic
QzufNQfwGB41UGMFfACsUwNqL7bkCLjhH6/1IQNk5TxamYASUGwsIFAckNHMBEYx
K3IKSh9QMGvPcfgIqWWFcSbMTt3oteLTAyotM+Utp5LiaOrQhzunFhMtkDIioddw
n2B/vog9Aqh/nwpjxQFsBxZxC0V9bebJGWAPbHZI/CPX/wlfG5i0wawilrcSHmkq
1ple8tze3zxFhXklOZF6G9V5GFPuy30uQHJWoEpRd4JiLsBabzLAoEb7lmPPIYyR
YWXSv57T9c0wtewyy9JgiJGk+9d8y6eef/fc94Tt0rPB1s2tkMFzsknDjM7JOsvN
eh8gd34W8IzzUhw+QkHNX/EZPIZXSNQ7ec3z27fNJI2yIgVoUL5Q8YUPUazHEouI
V5S8pVmMqWbF21dcr7HZ5hUD7ts73mtn5W2ggemtBsug3y+sdGVkqK2hqTqX094r
08+W3VcUea18JR4abqA7GkhYSlDlK4ItFsAZJuGdR4zb65l3xeFFg9sDifVACPrg
z5HeXD1pGUnFmDz5PlG0ZQ4jx2K/WLk0ktAFgE3RJ3csNaAiap+tRDORmmScAp/z
Qj1RqcsfgpvW/Ijq4AQaI+Gfd61lLKLdOR1VqgDU/s7wTI6S9XsjgqKcGxic/l7L
4xuQseT6aMecgmLuptu3oUoEN8fAmOSdYTDVnLjCXtjike4rx7u7wI7yWzkA9uc0
7NTpsX/kz/orE0mMGTYpyF6bAIY12XaeIM1NWN5TsmQxe2p7o/Fv/pGc3cCqGd5J
QBbToWM1yj5EFlvFeK2X1Jw3FX7gGvr7LJpaGHbiMYiyEGOXeTttENNKyT1ydUAa
1qN4nSdJ0E6SPaVbFKeijmmn3iYN9YSp274NgZdtSOwpdWm3cXEr9PdaFo5aReb+
cUruDigGooG5J+EsSVHsa1emySpqVocpzRgF5T8HaKnbWyEF2docZaW1i5DPxAv8
mxqR35JuLHEaxgwCu18VoOmWO0ngn03efivSlyui05snPdm1uK1Yg4y78okQZA5z
3LexnCNxhDGP6qDTedju0GNa3yTVsrSeaa6+qrs+V1zAl9jq0Woz1rvgYJfD4Uhl
L7N3rAXZ/+qAARfquORCD9HTwyf/LTyrrqMMEVH9QzmGBMr0ajIaDKSKFva7Sj/7
rtPOn3uB7FwmA3HEdi4b61EmOmAiPHLVRwmWKM8srV9rjSe8yie1HuDDw71QHl1P
5B3qnC/ATAKqds6zXQJ8WKT+F28GnMcB6mmFqaLbQdk5qmhjAG6Pux3NrpVpHs3P
sq47zEuNWLQYtpk8dC9bnhNc/uFMRxtymcRVlpkLFZFqhPlWa7jTNHtnnzl96SaZ
nMdLoNkS/g0IQGYgtYmKeAJfjlFoMA0MEhV/+ZwQhnmtNnhmBxHVrM2TgggTDcsz
ltBbLS2iMqD63a7hjldKp+ulxXla0AC3/02MCQFi9VO31f419yMJmRrBSMqFRSu3
SGiuSIFTGU8GFzZTpauW3NvLq5GUsxYgmLG6JV9OT60TWz7QJGX10dQ00q80UrFw
XuXr+zAISb0nj4BrLjonbrrwWonPbGBEFZkqB01BxHK2u+ktwjwKC7Esj9kQQB7u
vnf3H/8D3Jsv+DMVfNyqTXQzq3jNLJjsH2DXn8mWKI7mwQzRamypjMR1nrMMh7cK
+718S5lkLy9TL/o9mj7Ta/OF5noFRtOMaCsVFYspU6HNqbJ84Ua86XhJoxa+I0bY
eaxcgeY4QiCNxAgPoRBSp1CwKhyIjvgPvXRhKKQ6qER+pwhgKUYoQI8W3NIkvoBq
yY0bhu2iaGYrjg8PEnggTdIU4NPxDaBuotaTm5ncz/1Zs73zGua7QMFaA6mBVqD1
Nvg8449JD4YZHiA1STIEtRWYGAQ08m83I/1F5ZUYiQI98kqz75sFzQJ7106TWhSi
Y9IPf1lYLlB5A56hWqfRd8Xyi+T2vj7Gsww3/ZSnR2G99BrFxFZm+m4i5zxFEXxk
PKmqq/ROECUC/eGzhJOdy5hMKoWWJ3C8zikQqoU3WblAmWPP7M79+lt+osdyFJV0
3rpfwYpekNC7NuS1KvhyfLG72ALcJGPoMCO/FFpjD/LQVXREyKVa9u2CkprXeeqq
39PqQphTDwZT+WGq1TjHh5YXxlVGt7eTtGbL0yEeLV6eQak1JJC2UyPVgpMZrLCe
MxsA8yHkBcfc5uITE9+Mt3sNglfDbI+6kT/XuGwdhBFpPbs3BJQ/WSm+fq/gDnw6
cqICV1zA6GMl5eXpqrCjx6u3CHxhHEVhi9zooYQ92PiLPQzA6lACnbKEg2dmUOdL
+FI2stzh07Ked4l+3VRzCQJJMUIdx51SAyp60f8lHnY3qKmRaquxz4/LZeYPdYd8
+q5C+exgbknWIIP2RAEdYSVehgyRTmVSdvQVD46grheD0jtbcZuRrGkoOGfBnWCm
h13izfB1/Q8Honr3RA2kQhZ0+kjiUNrmx0QCGdwF0XfmiJN+itl/6XXzEb21naM9
sY7+CdUzS9Aer3BcrXtnPRkAu22CpJ+qWCZNIrdQc5PqgHMdopnMqmN0L2awo4+f
voKU8SYOXe73c0YMsuc6wX3wpeQD6joYhlb/z4wOxRBIfaIg4pN8RhFed0u3tyy9
C4BT7cpqR3q/mHJ1NHMFc7Qjk5R8KtJoxyvrk64UJHuZqCloD7eCkIT5cXljNw26
LNyRgORJ/fzIPH2V9bSyKlP7vpI7YVRl32ubVrAfuyuRfOKF56M8MNZg7hz8yBfk
g/0VaQ+GW3gSOT8477b0yYeg8pxbDGUWe8agsVMsHVZzlDlwj7j4qZ/6a8UfY65i
pvKLR+1q93YQ78Nei+3ma4u8figMb2rqSOoPVFLi2HUuROPIdRW2dB/760gFT+Ev
o7eUmaxRRSNfvTTJRLiQb/s0XtOKa1oRwcqGqV4w5iEEzLb116xA0gncDAioqfE6
eKT1ykye8gP9HeatqGwZ+WpfPPVc+hviNcSRcuwSdxWGqheXzzM/tEj+KU9HnIxr
rkQrziA9jdEna78pxVz9IOKgRBzE5VUCmwjWLQJ6XMs3FhXejRSPAAgybxzsCHwj
/v/l9AzyjgCczK/NTAzDtvkLlyFv72iY9nZibvacvh2+y1q3qftGPvMG6BfujH5T
tfWtHX3VJkh385MN6EiGgyk7hS7VF5zAqdCGLnzap5ubph2iFyBcXxlN9WhXfmjF
EbYxHlNlc8naYmNUmlSTtPxOPp9vpCEC0bKmKMvjpjeGjNTpZva+35WUzru2/lcu
BKBTkTs7CsbGKnDMiACsmMoI7Xd3wwhinka+S4OG0nA83Ifm3MUhnJp4lZ4ELlnF
T8tHQM6Y1OuYONRXl8LSaobGCzvsJ69i49OhEJ2Q1uLNlCEaGOuK+9qxwYbaYthg
xbkFD4HnxUbroxF12xlK2lESP7h+z/MnKlb4Szhgm9BcXjR7Bgf5huTIGyOlP5Qm
qEDG4qhRWmmVEgApp/u74K/7YY1cJaZi0ZIF7feK5AkTpjyJmwKC7Yafb90WLzej
xmLznihpeaPG3Ju/6za51D5HbRd2vQ/CsCQFkwZA1DRhF5s7u9IA7N7Nse9DD1hj
dkf4NIZcBmBy2bMZJK7ow04cx7IVS7ldUxcfvynjOxSD/hdp2lQb5LkgCZsklDtm
ANAigQbosJF+GDGTFKWyLDrkZBZJcFID1/iWaU5biY631soDuytH41KBvWvrtkfo
Ba7mCtmcPqb/RRgLG8p5NAIHkMF5H5YvzqM4TqLn5YzTo4qRNfgFySnXu5BBg+Cm
2djHOaCIukhbL+alfk1Ac6UeUbaxydwpjk3sp1UzYJmAzeqP51epo0MDk2kedQNR
GLbC9/b7Xz5qpt7h0I9ebJNH2mTtXVykLvwXMcQTQm+kEaFKV11EnuDgiaYba14J
vkKZ4PzUWixz76WsZow/0DyudWhWy7Uia7zLgcLNe0dTbDXqdAtbu99ldhmdb1mK
pOR8J7Vl0y8amoLIZKaEfKtm4r292dIFU4I6ap1Yvxvkw2o947iBWunF8jcAX+5b
qNQZXqyCVPzRrDa0ZdYzmRVY2RV1U3ZNxqM+ZAnlv0yxsDUyU5HtYANDsxb/m2qA
EmOLZrH8exNT9e2XWMbT3341pykTkXKLP2f4j3+PM1oKTC8vZ2HNAV6122v98axE
J+y1vLBipQb3N4geg1qP6YVvnEfbV16awCgpkitmvtu6rntbrqTTp1o3M//qRjBp
YPfPudjAGeAunYxYyd/Auvq2N7HIA9QIoVNxPDeUjX1OUJgJrFxZxeQgG1KDypP7
Q7cp3nI3WYXx2UNtN2KwxJnFiko7LJ7ICmVU5bKtNBqDrpM14L9s/mEFie+5YNgf
fikFYGeNmqwMi4sNfD7KDMsomr8IhDD+g3LJyrGUB6e8g6r6atlkven6RvRb7yVz
e8TMzj2atQFze0X7h67jscdwJour3ewBzx/0FfPli4xqThxCWpM5raJyundnGWr3
BKGNkCn8sScNF6zhe3MfoY5bcNAfhKxCUXEmiq4tXrhFpNkeNF6oh/TYARwyzut3
st97sefWfxN3+gaNhD30cy2V0rLHr4sVwClWKaoH38NGqNVpmDKZOhBBnekZmdUU
suhLmO2DJ9GTuoGuL0PtoheqS+Vl2cIA51LxIO0elBgod5rGC+DNb2EkPZt5J1bL
darmbDBeAPae3a4SwYhzphxQ9Ub+CQtNS2xIdkKotWmpYhtVJyqwultYh+gHXhvT
Hv9nPYRIrUMNjW6gG6mtdmbjatBFt8rJZ+VvTSU9HFVuJ+KcBtRalODIhFfurnt7
Q3H+KZn6uVjuX4OwJbl8Qpu7ad5lY347fulpXJ2CMRvHQXwHC007RO/KTvhr13Vb
tvPxGxkJwAEzLeCKP3Vxl3NlIP1z/u8PhCkM8pGzwoKJSGUnxeYjA99EN3lCmudk
mZ6hFBz9P7MNTad3s/OAQzKTqsjJWaJgMppjzXf3QMvfSuSKy/6+Vwp605KoOxUr
pYx0txVkuVmzrRXwbHKEpCCg+VzOP/aMuVpAUmUcBgz8DXxGPB3yDq5zSm4C8aF/
jeKp4gQw7weAHJzWmoZu1M2gRc9tMuxQRjTh6/Ei231U3XQxpO1wvzT8IAIiMIgA
iK7CxYo/vg4tTUYqD5QhLzoQuCrK0GmNyiS2sNDwetCDM1zOXLj3m6Btjg+QQPMj
Az85BdGJuklwKqyZuKXXvgLqw5p3PQbYNMadaRLjvMFCisbBkpjnCGRO4BUAWi0h
RjFAQrhbb3WQPgwK4XNXoHKssFq2N0Gvdg06E28fckwbRb2elD+lfehhhTrhqN12
8KXzVO9r7YuszzMexnebBbpyV90Z4XitkfS8Kim3Vt6HLSpxl/Yf01R8cGBE8oSq
SlWwjOGDnRPoQ3eVRfeeIgAoe1B4i8WgbRtwCzTGuW9UTPWHWr1MsnKNGgH/yp1h
H7tjZ2YGdlLXJnmmhWpC4ehVNBBaZryCLMp+4wpC5oVWuzb6YHpdpzfVTqgMaJ+s
p5Xk4YWrxBldFnJZl41ujQPfHbOZ9ArwWw9896LJWVWxQlQmpDrplXVf35JCUNam
yTi8esenwr+WQiZLFLS2ypsu2Nwe5/VkIbmWfOCE6zR613zo4Q0JPmoE71YcFVyZ
SEuDtCj2YxkI2OXN5hSkxL9InH+Db8CTdJ5qoamCXEY1dXoasvSYQJEy/JstBz2y
+WPqUPwHqNtiiQwUzXQuMy6OGMMKeajvrO9TR97+C7JUPoI6CYscetEOrLSuxbHs
xWF7Wgh9uYAcQS/U7P+YcrE5e/Q/QRiPF6GFSQlELF376nIugFXzRHZcvpcM/Dtc
7IVHLYQnTX7hSG3f0MXvc6DJ7erDdZlErYcOMXvcGC6MPAGAlR6uhR5/lHgT9cZi
dFLl7Ppguajd9fSd7fM89kTgeQlSyDNWR36pzNJvRpxsXaFSZ+qzjDvS1gHFFr11
QIZDAoaFnCQT/mk9IKu52NYqSZfrnSyDT1D48f3kZEH2/ooTb0NZ3uE9xTLDGGSW
sUPf6pmew0rp0+EcO39BIW1abJ3jYF85/7mzXNmlZg6sPEYquadR5sPmsjqgG9/0
FM53x4kSFOQ1jC67r2u4t+F49MsJL4GwIQxKYhyqRRNz5nFR5FKi/E1TzQ895V+X
iGUoBRUrsez49gLuyoNCReeMR8XZUZPE6dbY32m62aAF1/I7AmZTEwNpScJd084F
NdCLD/zOXPUEQBLpm6rhdO/DxbkMAiQQ6GKYuKDxPJkvNGtf93CWLz2N/09DYOy6
MI//PLTbnL0tpKJ/E+jlEybeYnp57uJWwMfaOjQWnpRbjSB6Gb1/KSMTkIqcGd/G
NCYsEGCX2Ejc3Ck66KAUDCTQ5ttP3H0iVfa25wLyFpEsus6NbqhNQoA0mhP6yGh6
6qIpd1wht7DMdJr2FJxg0DyFK9wjDnVuYvTflXIZE2rz4tx1VT+SKoMUo9J9y6ss
xJexNY9Y1mqypEDIALUp99stEkLhbyX4PjkmhVloua2pQiTkl5IvF2RecshfBRrv
nFphOpnzeai0gBB7ikoDJdv5H25UPGRWvwsybGzDNeWOd+Q/XRP+lgN8+SueTHeo
RAD4tnPSVca2uqSlR7KHQbch1O434+86e77Lahh6tX8TJxDCDqMb17uZWwxV+51/
t5EliNrZaFmEjr3lAyPBQzel7Ah+CCB96LOSRCBHAfCaWy8kjLC202RtQxAkTiPH
ByYeKLOnyyE6KwP4da9jFuF3XQHwKQ9nsMHDUt+AmLr4P5MQoOsOQgAkkaOMQZvo
yBz07S1I7we1o2QAywAnKGLeLywYOhLys7beg4piDzWJiH7t4WMLeK6+Y7vqVq3A
S4A7ElxmpEm4Oxof/Y8yVSrN4Pa8nEp4AbHioRdEt5eP5aJKawfmY4phLREvwsWt
JYT66Lma50hqmxFFPGjHLlHAFj+Q07AZlHBkauuATOd+DiK6ODF2WxbjGX8CSLGt
IEJe7ULBJsvAuMoFTg+wY+/9/XGn7HDFr/j6sns1vK4NxMogxY7PrgCLkv0sGXCp
IxoFeTddDfjGgZVSPuv/Qomb1Gbyh77EgRkvaVZVTPkwttcBy1jnvg3VTqAEGJjL
EZnaNxkpS1BYQ273ngWorlHIeAdk6wRdN7OLk/UMLWQ/0L1jcMqcIJ2MBT1sxG7D
XY+GcFoE/862fQWZ0G6GAapfcw5ml9wxRhRyLtEUqJj/VKVxF3ZI4Qm8xO+8wlkb
b+cGCsRcRzd9BOuZJsnKiUsRjGM7+pbOTeU0whFNc+TibWKnmPjT6YmvUXR20OCv
CUja94Nutq4nnJwbmWacRax0L4jbmulfIzUVI9eEaGzZDyVm82OIzLl0WKLgZEl0
OiK4nMM9ik4PnVuAgMf+alUGx+5LUW6BLV8j0YJ9IsJKs5A/8iEgrxUcevrFdRva
Ol4ulBibG3ieuxA6QmOFZs6hgYEJTosB9gTa11Wpez3pEUFCisuLe56L8U8jmSP8
kWDc7MW4l3V+M/cEmOA3MNlf5Lh3mlFoLLxJ94s4cUuGRzSEeIpQpU7bR1Yb3U2j
W2V/rI6q2iW6GSF+m4f/Fs7SNUhjevcOek31MQESbImlRV5sKoweGzTdoSHu13j+
CDYey3PQPaVFgNV9hGVnEvN00p3C2wqSKudHYQlc+pla2ISRlRgoye/h+dMr8ijZ
hiiubg9ZWR8c7ieOGEQZSauvgcbWDoYJhRSzlhEAaqU7bZ5OxDiXyEpV54K2jARL
2wnUgwRwgOh2F6b3NWntQrXX2/SgwjmNWgiTBLPsxOpwzvA2AoyKnqGoJ0EkRbAh
TADqu9ERVsVseQ/+Cy+QG9w5147JhW08SEcG+DNhayeeCe1n7pwQanXKdYSf3CGh
PPsYWq+cbkLyFrt2e1SQ0ir4CYRUGmF18oVuFmOUcJqDDivuUEJHqKxr1njxBqoX
mdbPgV3WOAp/3ZAbVCYA9KamjfC577BXBWxD4ecLnvR1fWCRoWTQL05M38CSJzEa
O7+xC7/0e5M4iiKqw4JuxJwo2aGXfZkhzbBgUo9iVpeZk7NWqrvgNMKPiFazCMPm
49zZ0DF5wGhStDjfhbs0kic99Dzz7E8CnhWgGuyPc4UwTQ4RoIp9AK08gP5F5IZ5
bR+9m5uGsJgjtCv4vSLTAlCQrM863IjXFB7fofAQ4PCb81Q3NTrRDkAnGH4zQFBC
0KjJv5oyPXufY+ocmeN5tJdqcb8HCEcoOVCT+rf1tbhzePHrjTwut9xTOTC5IkJC
/uj903LgduxNhegN5z2aRB4vagUwurtUfsuvCnVrqulR8RaIpakfX8Pg4cJvI/67
I+U/sxfEUzvnL8t7NdsgVuY7UbyGnfoDiEuQeeQZkoLW1dOq6wlv5Ko8101byrKb
gA4WkTPF0ZdaG54lpldz94g0aA9dvVgHlkcjZBGSHzAP+0L5V3Jm+TeMgUidrkq2
xjvEXUM9bU3Iab8TSqakObsumbncCLuX9mBR6dV3A3KcCf2uyhJVMhAH0hjZIwCO
Ar3a7IsdqY8BO/YrS7E2JLMJST/ryP6FJe152u68erB3mOFdsZdMf7stbkhFmJEF
ZZf8+oUhkGwoip+YYtzVp+8h9NN8KrAR+wGSUhx+u0oPMN58GHhdf9s53u6O5/wd
z65LDLzCMhdcFaRFXnbZEJiL+RlOvsCY7C2vCz3wlEkmTE2c5/RfOYiBXJLserQY
reGBj1EW/b4fgpNY4p8GmNN9PTtMqL6ua5PhQmjEGqjtoB6VXmb/AuMnVS4ezv55
HmySNIXdoLOfN1HD+IHOdyImHp8rTPjpuQCSXPwfwmVqfzkW4D2YjAYmZuEDhC/X
KjDsS2haQETLwFUdVr3G5Y9TbFZjS7q9UvdmwsdRX3y3oNlkdaDpaLYkpNVUD5fl
C9VKaYuAjQw1oKPamqVVe4tbUYqKzhWy0nLCKPC5hlzkFTOqxBTLATkSGq99oPUy
RwBcXwlyexlwVWMS3TOzmLoFBnv7fCSuFRdX86EtTnDO/N+eSVboI8vd0pKRThr+
GAsodW1rQgqJjgy/GsWTZedI0HPaxcK/mv51XCOusjeDCMT/PeBV/wauKKSYs2il
RBcBPvpQFtmN0upkr+JMsplcKdhaFwg2sZJt8aGd97BEe6QOaKoRNooZIDbWnZDu
itBtGp6gg3VAKQqbooROJkxJ5mVgPPQ06Fl1lm+vsqv8PCxqZ4q8Yl5WZWIfxJKr
aB/AxLFimI0xyhlbdJv9oivox/fzyBngq1u8FhDR+vwdGqQ7FB/wYXmEDhyXMAaz
uyU56aheVt6wAhLS9VIwgAIhmThuSMxQFHxZ/HVBKu1WMZNHW9kWkH4bpoh0p0o1
1pCplPNH6ZEJLzYBOP1Dq9ArkZ8w2iFuB095H19os835jP4MygwC9o6x/bpht9RC
SLPeUCmuL6CFych1YLW2HnhnHzua6TNItlneRRLtmSrICbot4SLeirRAjW7W9ZdS
sU74ZnISUna/QrvR3TezyA3wo51twt9Ql3oiMfC+nk6TOJXzJAmollSyqkCwAVus
bI0R5/klPuPtl5wBh9fYWAKPQQVWX14DyFQCPgQ5T65IJEhfiIDGQMvUgO48xJyK
WZsoCRHTxvAjE4KQft4YwDMGWQGr7xIrviT0Pot58deN9Xvfezaive8ZEMmiHqQl
SxNUsc6ZQvL/bOWZmky9v+ph041FvM7FWoHLMwEOR/UK2aE5zk6CCknj4yiRlxM+
1C0zV5H/7YbfK3/162FOAp8k3M9p6e/h7BqCa3gqtYIhRI6nH/SZd8KNhHM+36XI
j6RDQlh96JK9NsWjZiRfP/OLovnrtdM1CkiardMjoyH8YbDHsSc0AUm13hJi63KT
W8SAgAcHT4G2KCbpprNlbCSUoxGNhZY9URCtBqb/tEtFdQGumi3Z3DIeokH8J4zQ
aG/OaMxxKt9M3VT1Xbnb8Z9Z9nV9848J2ZM9hAccYXTne6viE9n6eKUjhTFhjE7N
hjr/mqxK4xTle8m7d0aZKntFPAE9/O2e45nC9nUWXGNmVE7qkw3AzFd3pvDBsrZf
hMpkS8HS4ewA+yzAHGhFFvJvTdlGW//27DOFsxFXMcCaNilyXtpHrefAR7SDH263
VOg00ZdjQD2ePW2RtdprC0CbYiTmz4zhcL5t3OkVsX6wRa4fbbiVeLI1SL57o2Ss
SWc5XYK5t1qTSg2vQDvBb89hHcsaA1c+SGZ/EyXUZj1v/+30HYvlptwbTah5YVeU
XcU8iMseQ2zK4mtWjD0tOG78a+YhhyU5xHm+uzonuxOVPfQZOql3I/aCJlAnC8dU
WZyfSFiKrCMPBvVFTsq+bJ0m84Wx/gqVBo1cIh+DghkS9xi6Dr77rorndYPzC6wG
78+Gg1lQfwCRzgJtNOv/wvLjIYf2CApU163ARgsatBe2nMrt10YGm7b1G9NGOlJ6
UaKoLZQROBn/6H2Dsa7IxvGGMpEET75dRbNUwvxTXbEJCCCuCzAsswN5YIMRobro
u1Qu5jyowBlx5nO9g1pZQvoWU0uTBu23cPl6SR2imJR/DG1pXl5gVIaIr30H+tx6
x8ETaYhYEJij6wYULXoTTIIf46fiRND8kInMLPzQIjQRBMUG6DOX73bgzDC2IcMA
4WY+FcJOxl4puWASR0/J1wu6nxMjhaY9eCDtueSsrmVA4Ht/coWcXWEEzIXvTQ3e
Vo50hOkRkpsgeqSlpm0Gw9gjtKI3pkrvr0IWybbT2wL+egI7H4AQXBJEwzgwh8Cq
K2FksDjcByesTWwqhyeH0ryaZYIPuo8P+mpB9437d4+eguN/YYAUc+420nfZUScX
dv875FjVcd/IeHjaqCOKCAUnX+PbEtFRfDRQ0bPJflGhL3KQFcfYsclphCstLZOo
5nY5hiEkAWE8asCwtrBRWEnUElpSH2+EoeSvrwpyIzVAv/KpuCVFSjHWIW72Ta5f
RZc28wo5gwKUDgVGbhlxNGmACmbUiYSm9SWVqb/vvCp3YZ7SI5bmvdOpN/8tItMc
GK5nqfqbRN37IH1QDFBRFJJMjuFctvMllHKeEIL2jfgHBUusKQkY962Vd3LsMC1s
9utpAEOy/K+fr8CM0bt5934Oj+at4OLRzcN+Zjqx7Knqk0NwWnKNynWtX9VvTRFZ
xhqIPOuNoOKp496tuTN5iAArTo3a3L4RV4s5PxMW6ShK8egFVHItZLO8eKI0fW6v
O0/TJIVNYHptVLSLMg0pXkcR2FCoV5d3qEE1Pv0bl0E0l3lpdTJsDefqcEdAo5KS
GvQ/n+8EQh+E70PPNeiqnOhUS6CJhH6ZJn9ig0vgKPvIOo1Q18Ws8S0PyoPzRf+1
pvt2sbUUBl4H0JqPBtroP7wxKbrxJgnMMjbHOrlkNqMy+kMnVO/tDKKgzyMwtXGQ
NrhOlky+YgUTGK2q1YSKWGcRvWtuRUMEaSIITSB4+3GiN9DsPB0SEM0o3HAOtKYl
f6046kY2F1s5asHg+nOfiVsznXe2FHXhAELSiNYOTZbc1NzV5SOleY7ULrlx7zgw
F8ETdULJEOZsPOhNlbQKS6XBZcmQI7JWrdtEERg+1yK7wllT2YXEF7YfZiEl+0MK
IhpAMlbh5YQrOPnYzBYJA4nvVLXuhyjgTYjU/9eS7gMfRdGnAA1FJUnI04tpydmK
FArWhPDdLKw9pyRl3WlBrjxM7johv9ca/5YwnZR7K46i8pbkyJn216wXIvQJD9EB
5MexK98GgFRgKqf5X+nEqakTWxdsIdnlpaLXcPDlb43OKY4qhm9h+NzXFKgkk6EH
g+2nLEEgf/5TBPMWe805y2Jq8y76DzmjJM57744Gw9xhX2yLAUo0BFOyotXz0k7u
H8w5OxjrVvujwZzvDmlD9p6K3sn5/eaJiWQwkeJRqm5XyNvSe/1WL6vJmJ2BZESu
mxx1FODwIwxoqQJPsfacf8WwyhdyC6MmBauwDPL1soVhSavVinUTJb3OhDk0B3FQ
FKSVF3vk0lVpmL8JhMh0t4Bp3ZaAKdwo3Oo2zCR1oHx2nnJXeKAHKUIRELvmGZnL
GSSwqqSC9DtmMFmoTnRFt/sXWnrLgbloho257QXzQHKczQTbFvzY3X4h+YnmI5q5
euCm6x8XmxA4r47N4f4aek8tVFeRJgxgtD5y0TpuFTIxOEqfyuIDsECyVXH7mV7M
SHI3/VNZ15Fu3BvToMUGusX3axib5vnyH2FVXLmDwjebXMsToaDY7GD4Pl8x59uD
WnZ4mf1VJhB1yj8MjmWt15L8Exn0fYIW/mwsB+UYcaSpAnZl4zqupK68aYpCLBJp
i7qCoe9Hm3nOx00q4J2/jhQQUv/zvKyawGVJ5OkC6wWqTAe+iCpyNcHCRfxVuiRP
jWSQl3JJ7JnzR4C9tYT/9jyxUxsZQ/hHNn02Dvsa6+ssAMPaPMvHU5GTehTGCB3L
YbBluq4KlpiKRuaiJiD0QjQF62PDvffsVARCyaX3VkqLg6y42hciocqR158vC5Yp
h3jr3u+M8aPPE5jI5PVQAt4n/U73EgpVHLsqtnaqV4STzr3CjHUh3oYrJaZvKD/C
KHEBSsL+/V2ze08svGR6Wqge9yJnSM5xmMczlMSHc7NTAyOwmAHvIq9WTk7lJx+3
o5ISWkcW0GsIM1qFN6x5fWU4DUeAEpIcNplzXWxk44o5wR0JNlDjC0ke3xHkWjpI
ORNdEDtcceev19lsRMBhoNbwbBNxZ+q378T7Jv9FVxXwpQEr0ImFydtkeb9aPVcM
K/hwYkcsOn2MLQnV6Kx3SGsS9IWr8VhUelbIC9oUaQFEzYvVllnKtycinRU1lMnV
DyCWRt+9PjielW0UhzyEGZhLY5ItGyTazi7Y2yXOy9JDfOHdyQ4/CjRkCcEe1Joh
dd79z50odwz6wbP1KoX4TPEq8aTgYNAeJ0+rQXxIYL7lwkA7M9IQg8FQcq9BFDmU
RnnU2y4fHBcs/jJVx82VeyHgmQnuNijHA69E1iQy4AYYiSj/B0ZEtoLcTmFjrrYm
7wdQjGQvD3FrRN8nSQmMcrjqqoQ0+ZZF3aJ9enrMSlbAZUgzTfmOJPikJ4H1bsna
Bj3NYQqZC59ioxd6xqf0snTisCQ/le9K2Q+Do6a3YD2sS0POpQz6dvmEowhtIj6p
pOfajq4e95K55K7XaqNrQSrl/I9kbiivuRPHxOTfi0IMlytFIW/5ISs+e3b3JMNr
ZFFZJIop5BFzMgmaen3Yyp4OpipO743AGwNWLoH0Du326uQxS7r7eo9pK+bnfjtD
Cwf2zM5mKEOWaeXO1nVqcGAxzjxzTrc5NrbEy97qrAESp2UUhnR5RLGzwdVulsuu
LRtGOwSMKChcWzVkNxJYQjOuIEWZPy1ZAwp/GY/F/hZUykrCjSDO5Tm7KZkMJjN8
OcTNvesXSGKodP/sZWthXVtqk0claWbOiyxeS1iLWTTcUfA265FP3S73gdh1SaD2
kLtiGJ8hkNfQs+QbhQX4hROTdi1d/9e6ePL1TvDaMuWQ9JSrBeTN76yr0FeWTh5t
WX4QEVquYNu7NTF/bHktBcJF65e5nGwImaU7ItGNUCMB94hIxL5OJEvfZ79H9VQQ
ZEQ3XmAF4v93hVXdAHolnO/NHFZtpG1e6lvQ93qd/GLVMsp8fNiGlUOM9NJBbcn4
lkjZ2PK22en3co8es6ktXkY+VkMEAPGKWH/pQDR58o+VFDECrJmrgrLqQ0/hp8Ys
dQvzZhaJHIaqK6pIiePxyJIOfItET7496tfkX+szfjCAjxg0/fDczocX9xtdsM/N
/4LKRy8QLXAQt+D6El6ZQm7XBlu73hX8YY9mcT/wS+2XdnNdb+QEiPvVF5w1fIOn
Lk21Ak2r5HSsx6fxFtIYkHIiWXZwRqmzCeVmcXy/UdW3P6hVVOumaIPNf6WENsDn
8MBFmLHR370KwjA7sIc2T7YeWEG6ApYSNdNx5/9l32O4Z6xF/wAIZc0xjcGoFkQp
H3OypI8RcjcHSek5D1h+PtrdO9ZPN8UpqKcz+IWO4CFSCmYLN+QUU+9DW+4RuLqf
Oy3bZ/O36upVzqr0kJTUX0RCmT5xBkwb0DnW/XYp6l4NIxkTb8O9nvkY+U1ChtIS
MH/VngJhCmxARnsSaqjrM5Mah1ilOGC/Lr6fjLO9sX9qvhV0haafSRoHcAI8rGAy
r1cHDAafvhlSOXBk3mCRjYCy+8gc3t1u2hjeYOyximPg7w2YlJRBcgF7iBz5ikqi
8ZBMn93or8XPrOLscArmuGa6nskn9Ofur/23C0JQQvTVs/zg8g2oQJ/gnmnh0D4T
oy9LCrh3+8bCyoGogPEe9TYjlJAscHyfo/xA1Z7/AkGU1LbI8jw9EueuulhNKVFM
adF614L51mKrm6KWBvs2LewZvZ0ioZVkxyIOOBwlXTbv+kD6RoT1L2/EPeMgJ/wW
n6flfkORY4nz0zJ78Kvy9zW5EJD/QBNtj2tlk+yoeCbVUJGnT9tJRrD6/7wmvziQ
nWYUAtXbf3/KzS0WuwDZGuJvbcGuitdjUSLjHGpDsAin2ISydMAtwXX7jbPDHqBA
SkDn+grpP+2HRuwmyW9k18q+jefWiaxJWaMVfOFCEHEuYTXTIfZA2wzBtx4mhxBc
JJ23d4Bqv9TcNMc/Qr4nrno9bAAliif2XvtRAKU8NxhUI26Y+FfdPRAyF3T5y9/C
nE0EcMeOOWJczinwT7ttIR1PDEBLki9cONf/v+YCxQbf7028QhJnEZzoE4sJTIId
opoQ6aePFzl0b40cFihyDAKiQgnOjq957b0cLOPmelUbSScCvWbjSWMH6I6nQdDP
BOXT8Dn9oOg+c6Qy9MudUo8cAX/eFk9Gcqu89JLaIZblO2/JXDkY98MrSDk2AbCt
nzEd9Q4on+SkkFRQorCN6sAvEzdceq9Smajr+ZNjp2+wBvA+QI8xZtg/1no9F+Vk
zUxBs36zTS7mY1dR+g4/yEbKpLbw7WO1mYeoh73uWLkxp4kYl0PMU24H+CWzGOjh
2CHkXIdkCa4wCkA6dXKpHSNNVQcDRso1KN5IPMbkDWnplN4OnsC9WRVbJ9xCPsAb
LllBVL/+93IrWPFVVuKBdxMbAjDmAyBNTBoA8hxPcXVxkCgovvs61hUyvtqQWgtM
gSNy98No2LAphN/T+u93xk7W/acZIrWAJSsrJN4zJ3UAd4BLJf9oNL0Zzym0/COq
lsKUILorGP1mm/qkXNzjy3bdsTHXiIb8lxipjzen1dmkdWnNHxItLZ9ESQEaapSR
hjhwhTR7rEjFvIpufxw8QF1Ofy7JUJf/eUlRNB9tLTOBYM9zdo4TVyFSGcne9AyG
0GhpEYUb1TwYjZTcNxLTI2g0ZL8TZ9dRFMBMz9ru8aM5hmzmE2nUiYs44ekBbi6T
6W9zGfE4TzNPjRBgjhCaqvxr4MUcAJpocC6jbF7aOUkrlvdGEcfjSGnwhUnqt0vp
+6tZ11OFeixN3Hc0BVj3s95s+OTfrhOY2rTBQHVkIpgss/c07/dXcuhu7p3NznII
NIvcHMxu/rMCE0Vk/SPmZ+bK5BwmYsXhpQ1FMcZSAdlK0j2SGxKw1J87f91Nop7p
karchLscXhmzTsp6dAdz7bwUsKehuyXQZ9+d8Mn2WAhrXEXMclvf4oil5aKSTpOB
bNMZv8i0j+5AqUchcuRq0yTUg/YXG8/0gE+nq/4VXnqydUbUyYD68sA5xdZ/K80g
nJavShFjghDR2upPqD9GplrJPgzDg6ZKa8j2VxDX1dhzVPK5AbCItME6Q2JbFP5D
VVBMcItcEltHCPUQXUXXiLv9PWJtl6YzcPXhhuaUAbvx+JZXdH4sG4Yropa3Q5yZ
ggAajqhzPyQXD65PxcddTyf4LWzyoqexcWo7kNxpZmP7Ea9fNqgh63NdPU/dD8Qg
XqVNlt/MRRGvcVieWb/oKPVUUvE+H4ZwWkRHrHNxfkWJIrO3fYe9cHfOqpCphpPW
FNW9iGwqu/ExmGV8xv0j4j1ts86krFbfsxzxMUL2PBf6oNqUgiFceqxhYPI+2NDK
mG0sglI387Gygy5rlSSSXM0CuNaZ0XDyAb9CyrkRpRWW1vGRyAQMLY0c9uhgIUYz
tRCdcc/nyIvKImQ23pHy8lanq6eOY3N9blZWlKfabK44HBeYSASpeWofrteR/dzM
amyuF2xClSW5rTTAwAsVOAVp36QeqM0OCcvej3eHMgq9g8NIY4KoLMjSNFGJeWkG
NAcBIYk3CKwgFCCUdKsBYNnEHVHOnTxIosgPZnklzGyc+HzD0e1fYnHQz6LdDmMb
TYyPCijUMsHPetpycO2sW87/mwtsW0EOQAN3W0HtobqRy+SLiBVXKd2Yrc6+xz4d
+yPKioSj2nlfRxkHCkgpxKOohsGqLNBS4RUK+YrcWloMtLl6qqYVmB+ItPtxhC9V
xZJYy/vs7j+jHE9Lg2ON5REM+yL1K2MHw445ttrvQuBBlN5yJAM3kasQBVl8DPBU
nBpbruveL6ym0byCa2N+BxIZ/Yph9Y7eD98xgtq7CRF20hka0uUfRKhnPRiE2KnH
AXi/IDSgZhEdcqR8+BkssPQLqym+4mVEcGd/iJd4unL0a4YNbhFcwiQ5FW67fXNA
tQL/1w/JIEAKKN6w3SMjBXmY54V6n5IiipwObhXSqqhSewK69Ypw4fYPnDYlsheZ
t+7pMQ5h3MkuqApaP7o/8pm71zhvmZrxaLpMhub6p8q2cuElxDZKSofkM5T3TemN
cNvVlDu3mwAnqeWTcKV1DXK4nUMVceXvEmXIJ/wVtNml6r6J9S35IEAMwcYCOWSh
e4b2t3Hd79uluxvrTcTqMYfWHyWKJtLLjIhCEtuJUfEu5f52IekXiOedbQkxmCFi
q9eZpKdopgTjoKC3+IOLoDqUdZRuvwcgGLjTDruPKAXM88Qm/HcjjGZ29ZnFTXxA
gxJOMFkk2EJh6nynDbtvzjfssR7AgiY7WpMaBbFOIXnk5/QBP3rTe9uSMzFGi/nS
NB61Z0lBWMBUB42NbWi5TpDiy9OijJ7J6hwBWpXURLXmWMlxzbowE5wAiCQLmWzf
QutBtGQxSmEq0DFaDb69GMtzfYSIEf8h1w+Z5E+IN5F5vZhmXQt9dJoLnA3AYTuy
jZp30LDAvI1hUZ4RJ3F6ESGkJ08bPx24n9oGT9CHdoKDzCKwMnGuQAK634W6K0bG
nVvGp7k8MUgUo8qVpEw5awgE/1wTt7YcY1sHLTPEjAxHFhUaiFHwbDV0ThzfRerG
RmVamZG+AIj6/SNZE0wz3qebEOCQGYZmVkM1ktNUaJT/7kPzhDWhdkWf58LMUnYr
22WyX0Z6i5QxTuuPa5tAnsysGTLyifM6EYsuZWDEkefBNwKRb9q8hUtQcBeiOmsv
GRYA6VXOQxIbcS0eQhPmlqO8QwV0AtA7CrnLYNghXN2PAVfPmta58H0A2674vBjW
ItrgP5wGplsqzXCVgFnzpbLfE34h7KVo7f8O0e0ACAQsl6BuFqugmc+KGTjzHQe3
iwiVTY5I+obKlHpL370ON/3LNhDTd+6WvpeN2kqwqEs4nDHnFixCy3q3TEM6aHHc
uwg8uXGKArYIxM6E5OmUr4xIJXRKntuNzgOCcB0q+QcOpjZJFdiUvaWs61h9dNiu
VTJU0JniyrWvvax42NvMyVnLP+upebySW+t0J2tAIOvgFA8h2Jcy2UW1SI7VDHK7
6nVtpDqbkdj9+FsSdpESFDqH2w93abTgF+rghkAoT7DAcU0f6fcdKVp3/pxfWqZ1
mc2piMzh/naNkELRlA6ldeHmiXJjylV02O/cmYPcLt6UGpHW5CnjeMjfx1GgJirv
7+fybirw6ezKmA2Xw/vN60pbHG+h3XkMV919vrBS3H3qE5EgTG7Qa9SBwRAeSTo6
kADnWpWTzA5tcErfe6UgDLbODv+0l5Lo3TvhuGM1l58H61B7kb4RxYFRCX6YLKAv
U+791J2ymXOnICksO1NJ1Nslir99Kj0inmdrKxKY/jqMj9CgLUHKZo1fTVn97Run
1+1PA7+9n1qCf5II7eI8kVcIap/4kDKye6ayWfR7Ce6hOo+NrKowxiA9EHF62EDQ
OCRVTZEX26RFx1VKcBeiek+1Bm6XSfgjs/i5etsuRdo1Z6sIVT0M2zE8v8SDszUF
uFaApW08587Dp0pO7fpPRn7iQcL8gLuVDKecGDZAh9gD6nYr+KH7CglPkZU6P67I
NO89dBUaSMwp0htx1vCS/LFLXtibThj87jEA1ptilap8yj3sU2/p8RiD2g6zYLW+
drkU3CYYi5ZCyNyKJGyCXjQsyJRLoz82sYrZLO9VeyeUYHVdNuWpbQyssuZIjmaI
S+EAsuDmgwagiqINNrSIf+I8qUXI98rIaICs8FNrf7SSY1dn1G8f9I6bdVHAeUdl
C3KmWKQN+zFrLLnPZF0T2lFAgvjj64tghDUmKiq3tp5uqWfLWyaMb69K3Iwf5jyJ
KZW1VJX0FRiFUJE8ONsCBxZHXQkn067q2u/1gxkTIHX0BPZ0/YMiKkxJV+VPQslc
8DmRpOKfJ1hx9eKxiMydPKLdZIO6zQr0CUXO3Pxw/NRUvfmAEaWGz3pC5y1NwOt6
YsD9XznIu9DZyQ2oBjIeEY68OblY6YGOsgRtJI5gOx8Et5ZXS9VGVkbl+wUK3Df5
T1Boyot22EUj1nxoklMYW7n2rg5p6Zq45t4Nnb5Ad5dm7N/xU6ekFBRwTGoMqrfq
EJXFUBgU+WIlyyLU5t1xctxd5qiQNnDhqh04RTiU13ZGRkFFcFbowoLnSC3qPKYj
Ra6WmMga9CMG5pUYd+fZUssXLqCjXaZvWDoteWqu0pFMy9Nczao/UJD0K4gtm6EP
0e590vFmKxpoZrlqQ9EU0eXeDkx8M5WbEchRYrpDHYNd9ZUywNxdXfEKD0Y1ROEK
2jKyqvb4+OzosZ+2mb19Cs1wkbOb2rLbHjnnYC0NFkmDls1J5lc33isoJ4uyA3T5
+5PcwnNpUUL407+Vo7LiD7nsTmMmRcZ/IGw/SvJi0UyoLx0DmLg1ZWQw1tRCKujT
nkL8FzbC6xpO61X1hRdLDqUIVERkKIBJ10SH6RfXYdOh6UPAU0IwqxzgysG+LWAm
DXS265W1ltz3tao2ORz061/QLRdferZBGreNC7m9jmzufIFh3wUEIL0fwa/tMvmI
cVMZ+bDnuA6A92QOrlxUcJw7iwwDApdIQRkO/LMvQWST8tcPulukZzKbS41O1ZpZ
ov9xuFVKgUePRqIYscu5i37Qf2io1EZnIlTdQlBIJdsQ0oYVzqeN3Hj871jlnvy7
ylhu2QQxDwAAQ56j67m9DncnrsqARA8fs4akeyPcGNOq4ZxqiSe2bsQmyM2GddAp
zsEy0Ccx5sVqJr/ZYURSj9s6Fae+zjYBYonWKq3IkU892s1jb/h4btZlPRmh0Sir
sfr5igYzOmlWMeYxHNMZdtE55hST2Y2CvUdH8/3T5Sv4i5k6BoAdIs7Gj7TqQjBH
YYymFth5DsPFnt5US5PZQTLdgM3jXa8/WJYFuVO1pL14mdsav/XNEt9jQH8/4fH0
2m9HTfhLGLFqxMteyx3yvk0mlS5q82hAEaBx8DIcRQLnz1kjrFjs6vA0hqNiKJEw
Pwzwi/PmnV52xDWGfGuXVA35zIaN/fTn3bGp5nWqLrR3NxLOkAx1hs0vZ4jNf+DL
w/J7wBAgcbtb/f9LKSBmDyYSfrF5EiAOrmvoqr1+kSZMCenA188Rh+Pol/gDFxT9
rrCWRRWSwvNsTTcJV6otB2F9LfGpdaaai5iQ5wGn5rRhvSkO0tj3MCf8H3FmtJhS
cGek0KhboCMfoxpd29MBnmu7UIoEXQvxVuZHDKPCzDsujSpSs+8L/2nKTzZb8dQr
F1uLGbCz+8LQwgj6sCOcxzc+wSGrsumeh9nfGEBgq6T3aA8HKXQjVZEK0IBcARJT
CK9LOc4J+e48hTAmMJPNsnVGKlf8yag9WJpEA6i3NBp5pMbPLmTLGa/ccNXnHRVI
AiVEfhGoz6IjTcbbagjwalE9sW+wYXieu7pscFvJU05BRWk2AkGRaZ7HZfSbrDIg
KnbrVOuYn/HkSHOQvQhwF5PNpR3RHHpj1Fs5QIBQJ+5iYYcb+9ovaPx5t1hT8njh
3JVTXmj07Tq0zyehbpDYLC4bEZ9c2aarGnplAe5fSjhbLxbxYvYinaf8kFKf3iXq
BeIC+IGTlp2xxzTZNkQQDKaLQwlg17Rn3QHApPFWVmMQxzhedqZGf20SgN/IfGbW
hmcOFgP1nwNCarq+cewiNxrrwwSfX1QjFVWYLspCJKOAohiK8xovq1F42HrqjUZj
3XeMpSO9PH80vc/sz33wyN6QIPJbafy1TBzRU/shGZI4UiSvLz0V/1UKeLm2HPvu
xwaym95G7WEZ3istfFcuj9BolAeYsf4VvIlcC65EJSOZSxDalDcIUawr6djxZHQV
tsv/9mAK0zKFv06Zwonw1xvFdqEpPsEgwTmYfIgyMYBcMj6Xo0gzUlw+QdtFsw0u
ROxI3emW5hJ8LD5fSmrU27MIwCHUQE3Qb/zztUii4xQJqeowWuiux8s0ylPESvWY
Grmpf77QxNq6v5NQdsOD+WFLEgPd/+5diIp9NY+EnKgSmZChNueYU3iM21krSEG9
pMGFpApBmvvKO/a3gtl/eGrGxLH9yZUvb2rEQOwc2kfqi/vizwJ4UCYzUvwGxLk8
ZypLbJZ458qS/5qmazLURBI1JIc5qekdTgDc5kIpH13zflvl0D7J5p9uo1hl8bWC
7wcDxB/wYffgM2jHw7Sryckr4eEId2GqiUcu4vdRGf8YLMuU5DzAb4yFTukJ56s2
4w01vDrNqNywb9Wh6qVlong3tBOe0VcUeBSInyPG5a3UACyhKuIZUkDU+sjLR0R0
nQm8PbdmoFnklGVnF5GA3ztGQVEoeQezV54XLH6MvBq7XHoa2amwgAtX3SFWIsL0
y74JoZSLwZUOnDufcHD0l/NImAcDinG4vpFXNVchG740vRohGrT+xj4zpTsgtMls
4oyepoe48g5JMmItX3lMVrAo6Hj+KRPYBmIPWCdRXf46mJiZK75rky5GZTzKjeLS
rSCqbdIIeSOnEYFKvPYIDx6Su7Dy+lWJBKZt2nnXpAwe949tp4xEAiaxk8VLfmxJ
XSyjg8WXB2lIUXfp9+UhS1HpLdt0X8p9tdqlSUhl9tlSChQF9d8g6Niyg+mXpQFw
SdlJLeXY82dUEATC1aJwWL4LMv330J6OA9UHntspobf67SptbS2DFpsXg2UQsian
AokUsaOHXGYGzP0+6XYWYzwFm9jthpBBvevsXcoQAfYy5ee/o50/33Uog0z8Wpxj
U6joDN4g3/UxMPUX5qYHn29octlUpNZ7Q5Qo+UZiKOIML9VDjavsXXbjmCrp6PqC
hk0Py+b9wPPP4JytlvguJiqpQWgrcbwNzZrF2Vs6/KF37VYycMZYqLkQGID9blCi
hqmTKy+y8pUSkZjxW1bCq7TpgI4v59G6F4pxcbHXTE+UJ1IoPRjb6ZZnGYyMpmZX
5jLewI3C2cy6UaGYMb7CWn1H8UAa1tnlL/T8GAnMWMTaCu2OfFYBZgCPEguQv08D
oK64NNK553vWow0tE3cpIq6LhOjM1oRco/Lo44Tid6AwQyng3XKUIN4iXyk4wLeY
64oltX3jorjEVRN8HmtETc0jOIglzCIY8wVc1XOxZgLD+9bR8UTIYo3+bBXqGT+V
B5ekG0qk6a2p10j4ICp+dOXb2XlDe20JzkXsWHHlHbpmpl0Am6iCwHCFlHwrmYTi
9sddjuI6lGk0lKwg9wbQ3ecZgcmeEzN3NuOKp7aDtHkeCh+fg92az37n535GjwN5
TyoOODxe46c6AVwIp4ivcH0wbrREaAtlRdlZcJEc5HRnXFDdie50ZeIID08WrI5S
ocP7Jp/hQ6TOzOl1uI5C923+37QCjCtU6t0CQG0pO6J7vES/dRLVsY7HzLfhiPjj
KY0lFnLPlNUTtNr4LTXBqZtYBkYlS/VG6B/5KXTanXQorixLrrBoVh2LIh5KrsJ6
R+M6OjnJ5H5OlUOH8yS5toP31aOZYuIbi2MQOezP0jC4cO7zG1+IWAc1rZ0ftT0a
gZzrKdzk9imblpULI3qPaqM9xP/mSJjV1j/F9yNpJCc9Vx474kGAsZ10Rgte8Kbc
snPCyeyBusdGZmbm/xYWx2tRukg6tZ+t1Q6Ryp46ELt37YOmsY/9SKG/qdKk47yf
svP7TFy+MBJ/c5mHiID8l8gnDBFl+FwdV1WOyb0u/JVVsIfyk1JgmX2TzII3YUTI
HvCNPZLXA4Gh1nfqAma8ASuplW2ikmf0ybrmWMnBABd7Jqd309eMUM9EdgtsRgWh
hG1zEyeEtyoty/q815aHYIHQKWRlO4Hjl0Zb/3eYc73pnq0h3plWQalEXH4PSTV3
79fz4pr1L4C/BZfXx54y+0sc6lH99DQBNAIMZeDwM+Ehto9DmO1qQ9RrYt4pT5kr
fYW80VqQE4GaXH1EypUH6iP+lhCs52dbjZrA4KwGRnbnX3yxwYyG3uXKPnr4fJdD
GjiD7MpRAQuTVFEg7zzgeTqQB3ut18i8zSdC/HTs/+LEdrAsWOdauhVpDaWaM/1r
41GAYzu6JPcDFNSNDB8WmGhZkLgITYZBR10fwKEo3k01xp0RLxgctu14wEV/VgR/
XqkpKZ55JM7qYZHRN0MSzgXuhMIZIM0UeE+c5dqoTk1jUxTCTOGCZ5PZxz6LbV0d
lAQwwRro+/2quZSEbxg+42x2Zg9Rjv1e4NE89jKnKw8OXYbHxxQTsq0IAqodABZK
cCOj/eINt6x2AMagNR0javFLaJt/uh9N01k6yUzzVICRl3kqj4cItUNsWCZvkNSX
mM2AA76VX2FVNn0F2lSVFScUEieiWzyZdNZD1TlBPqwsO/jYsjnsPUG9lp1Twb32
Vuq2RtGh2DdhxglMgVEvwFRh50BJU2NBNwPhY2vwM3TpBIDXpTt19cgZsiEZB5Yq
M6zemPoGzVqpEfPVFb8kVAGbO6dmLAz4fXWHNmBocdcu8Yi3K9X9yp2i11XN+eIX
DxDoHzkVF7+SK/Sth4rz7ktUy7t/K6kziEcthtXK9zP7MWJZK8Wodxze59+l8Anq
O2MypVDduIN24FxJ2/eSxUYCXSFcbse1TSovkZyGn10a2dqf8juPO4mtupsXjAXk
EPLvXZGc3WdGzy8elOztSS5KpT1oF5eWbID7szg2rWVLte7WbQvi0Wh+bqhDyC1O
/rWGI6e575NPDXpfE+yLGH/XOBYjG0D0YIMdc1Y1v+J/R2LCjMrPPtOa0C+OaFi9
iauIvW8SR7O7KA1QMazaKuYNvGoKw7ojZuI3z6Alc/P/1CI2bgVK5f2nqDh6VzS/
q1UaW8CF/BiI0QXxzqGdYfDqnBzzfhf4r/P4cN6Mj4NajAT6rYdK7NpgubmugnVi
Oc3mvtY0BZ+//99bt/P1Bdlk7Myxxr7vhfQS3Xd2/36qMvcWUowVNHmEHRIchZCj
4c4Gu4FzmuWLJln6l5CgNAPonvEIBL3ueRfJ781WllZxpjrnS8J7uCvLM19TdJzn
9JDfyLk0BeOD4jjM6CzaE/YxjWgUt3dKa5dFBYW+cC2dNMymbSX8VtC18RDq97/G
IMQdi1rPffjGAb1hbbMTk3qAV3+lw83BKitbJgrwA8+htJtW4AjcNl+9paUSkL4E
pU0dsA84lptW+BaUANRKy0we0MSj4Rg+RlmYzu1e97KFQYNcPXWrFuXBXDz1epOB
Zztd/STEf836LkA8ZGckB29e/aKQd0pqad6/82sYU3sVIDAxtyfWyA/b3ELsI7eR
INFAtt1XHW1o+RTUcqmbp1BQ5ij7pJQPA1Kl7sVxpyYEIr/ZYCbCwg4ZwYJFiaM1
coMrx2bv9lDNTnjA6Q4qrqpsqhx6EujIlSGQNo0RNiGZhDwkkVN+0nOLeEwHvBnY
OmB/SHUccVtw0m1Yt5LxFCEkGE1qppDJFdifcXkymjXigkyJQO5MV21aHqkwL1Z9
9IJZ7pTvihNEGeJXifoX6nSCiWXG9Zbs8KxAXMzOmoLEZ76Uuu3dUmLfkrhRauRM
3boAr7NsIfSeZRcKGNGg2ZPitEL6atCZMU1Weh7dMrOSrPwWVWkCykZCOBpWoxSJ
l9bPBbDrZgRR6O38nkJE4yNuhcrINifQVl82wKs1irQtapoLR/KHjRX7tMeasOXx
/9t6yCeUTNvK1j3kWF/FbrWz8D6CUybh+WA1YThwHm/Nu0iDu9AGF5nfLYo22cEr
4FfG0v1xrNWoNZjSSmije8qW+wzqwz2zJxWCXsCAS+mhsLLh0YqwxCfjJMm6d8Xt
YYhQQolH6nrZYG1HtFQeuAk/vGKRuju+wQl24QBcm7pbA/eUofqvddUFxaz9lC9A
mTTNPx+Ya0Vveuull5R/4oFfc8/15lMetnRJfSlSuLoW1/oJAE9kJYc8d5anU9Z0
Eymi7eJYeuKIoihXWG9TbsUVWPQpXVi9742pPVXdQGeSGkg1t4d4gVDclZRVVMwx
p+ixmsv5uMO0VOUaijnXPsFZplTSSp/GD4zUcRRPiDMlV77FUoav1/sVKaYiQWFl
hXJHp5bisKRuXfGO7rAQrQXC34YlluQin5C2Pd9S+rc/W2LcNrPHfviDTyAGO0ne
5mbkEW/+n1dpeN5GmjjZ2sKglLJxvnkNN7vL6fVbx4+clhWqY/Z+tw4EoX4JXp3Z
vIf5YxWOWb9FDL9lfYimy5fTpDIcdfba3Rcnd3u6s1SEut0HwHiyt1yfP+Kfm9Am
Wdt/QMe098o8JUGgH8jHvVXujHAKz6Gtkmzyl8SZBs620PS3Sb9wC0g8vfN4/Bvq
8bxkmBrk2NeDpeEaclgL9sFAcexDAonpQ6pJnXP5zUjK33SC/XjQ0gpoXQrant/f
Trw7KvOs31RFPTe9fqKbcCfkaW2SK3Ep33npBE14gqe/XV6p5X1TPTLL7TKQxxIb
Xl6QVn7wBmlBPHbkcQZ8293j19Kvu3xGnNeNjkEAcuyQIRhR6SmrN5ThJkhkK6ZI
cy/5Dx4NQzG0A1VDe39NkpIksj4WX0KA3KXgvoSmlMBBlS2IV7BbhaywO1yMAhmO
CHi883V7PncgkEYIKmPvZVpWbKwIQbRfU/6baMN3i+W30GUfnn13fc3ZwN5SzU8K
wcfIICFGwZ/J41FLE0S9Mu2jpwQ8IyByl8MX4ony2qHAvJ5cW2CxM3nzxQ8sYQXv
L42ObjIIyiLrom/0M/FN40issoXAUpOiw2kfRLq+0tguyybMK5cZPIMFNqDL42ps
r8GDbUPqKzb3juJKRApNGpZTj9LdJ77onHeHJgZJOfUfWn6uxjPYFAzrQVMGubuF
3Pd8Hd+cP8++dngtgVKL2+PN+FIas9WA4v3DsMBwqlosZP4JIMo/0HJnB0g2ezu4
habcYm72WecJQw1DUZYL1nQBrgOuEmhUvQtColMvFKefoVmes2eO/YWOjm0arfpO
TzM6LE6na9xFUxZk9TH6Z+Fh+MUky1yKnRZQxr2dn1nD7iA4DVaTMKnzH2O/hwrA
yYcNXNqtifRabbI0WYkL/e3rH9QZXY5zH58L84i+A6qcOyZkneONx7YkLf+ntfCk
kz8ZfBxKMUyjv7hFe1X/sNvO41Pp5egQPe58WgDUfwE/70Ts7WUXn2k9KQjurS5r
1HtxYYQtyAl1ndPdIWBnMxaKvgurH9q6UFJGp/fmW+tOOG6vm3RtFD2Tb8Gs/ady
PQoWvi1Plu7uInqqUXQImhUdj5vRBYlO/SrfcBKFItKUnGWRPks3KkZSevFOLziO
LO8ekFW5g3Q82GKzkLftmSwuPHiM9M9Sit50uXsrXt6pA3criuqkiiolBlM3ttoH
oMEfu/tjX7cSqpigXM52R0SLPBHr/N2KTRUujbe0rhn+DHExU0VC5LI8WMwNTCig
DvcymI7fXL/QZYfNBunpEQ4/IPqO+ygY23w4kl3ILX5nDolLHUz8qzOknWuu00qH
8nTr+NREWku8hoK9r/GlkIIaJLnVp9KoxDsCmy2Eupo3ZJzdo5tIEIbpHkY4DoOv
WCJZCbbG2yOv4vcOGYmviBS+7R2A2AKDrKeaYE4l0pCaGGqfer2R471UGEfzOQ6s
a9OR7LHWr7x5w6XtY3p4ESBL/wTsLzA8QfzPxmfMnNxF5TMGaMN4jBD5g75e2u4K
Xl2P3q7oZgLgl4U2xA2WZO4+xpylvaaiZyz9ku/lbbRwprHHXnIsvDdre4vssj7w
ees+/Q72QScaavD8b1uhzaGhqOXxQE0ocxyvg7LauWlLJtyvJKkBU6r3W4HInh9L
8u7vRgVmO6nWnkKZo7rZCl+ZIPwZt6DxtJGtnuhn2sLF8JW/W4HgR7j2PHU2QsqK
BN7Xv/t7AizQy8hzyTjUYco2Guvs7t2Va4XKH48egXdKEmDyLh1H+/u/4RC8O59s
uvcVLcEoJtp5Svbwh+/BY/lY5RlE4k7PcgD+y4d9NLoZYmvAxJbr3rLe+eBSSD0J
YiTd9SR9H0HBHz4htUesVn2isTbGBGyjMWkz1kk/5T6imLZ0+os/AwL0aifbDa/i
tjrNZI0fJuAM0y8T1zi8ypE30euBP0rnbgQwcGqL0TWKpMWxvS84pTrF3NpPRQFy
UWCpFMXWbtl4R01B+VPHXOjXDhIO/73/w+/KYjZbSGyhli9EoXw2vKIG2Nl8D0mV
dpkTR2h0RmmcqcT/0g/2gjNElcR8BPG2DZrKyMRTokeQ35KRVtMtu9X7T8p/AoVI
d+TRgFMSaYlQgBULvrWMyApJSUXVTtCv6THhlLOV4twAAwWIJgqBF3JqP1xH3gMb
gr+NxAuX/lTcV9L1WvKFf45zszoysgEGXUEaKnIpp5Su3NVkBiDqHIXUe4+FlEWC
vpvgGe/HCVMpxZf0MS9pmNadkR4vWuJl4Gkmtt3vWEPDjEPjhtlxwrVn94GX+C1Y
aMvB6RgKCOX0xR8CEM3blmqJ1MIqfrF/1GCOYbdDmO2fm+HY/QS0XcK4yXDFUtV+
Ch9SmTiSMaHTNFHakY+R4xM1h9Vv+AsBC7qdHF1xMzc3xmD6lqGwokuaOYRX7GtW
+E6fp7r7fHoZtOZCqzG1lRjILoKRI85v1zkq6ChgQXwoZHA7wgaQQPTBUUI309mM
C6/8QvNKjQ64d3BLEUjL1Xdzbm28RcsVRSMLFRw0y1R5e4vT4l1+eqZgqXPAm5HD
Z25uIkSX6kVl7P6Nuhgm8avtjtc2GboDLwvg4tQ2IlaqK+yqHbzow2eAcOvfEPdE
aAHtZbZVUbp14n9/Xk9O6aXKHyJzA6PJdwgsZVJUZyvMEU+3VacqF7WWfqmnPyIO
cXXETaidtRF1EEPUgN1MbDG9YY5EnWFEt0SYGy4bq9shSgjv3b0Ee6DKktt7Bb9S
T96ubx44Pr3PNFPaXPLv370i+BlzRMdhhpz/QVn7R3ZFnPlcy7UNqFkw9ZXYR4qC
7I8xTu1rq95w7VAMpPFjP84L6R4lZyVJ5G55hNc59/uKKhvSbEsW3+FYcTa6xLYH
puF2Bv/P7hUJZC65nA+QU/+8lalKgJugcEWzk3esNaQzbo9h9baAVItPQLBQaff/
L3p3fH4SjlChtpvG/FqhqFlC8X8NRF8Ka1DmqOjRscYAYwtubex3bByphUFWccwO
uVGL7PNXCOhXlMBQJ9F8TfKes8IeFgRLNDrjOPX271d8jYRDuk1WvXKe4j+vDgiD
0mtcdmkkpbMCvd3CsN76N86k7+y8t2THX3+wZeCW6uT/drjHbtoepN8FcAl5may+
vMdlSh4M+ZcpGA8LHtUFtDzlj8ENNLdPk/gqSKumtXGNmuRRbzK4tH0cbgVQKtcG
yJSZFGlRdEElv+XOeAiNKkCGlyHCpGepZ+OXg03hCBlYr70iwebsfEUGzk00gKfb
EfNyYF7VwAAI+t9VeUcv59W1q1GUW26Gvdt2RlGjnaJEORjH66EgPAumj6IrqcGf
Af4aHDnOvVh4ayqZXHr/Hn9wNNMKwKht57g1i3UTSwgQvCX2u+xcVJ82b8DUD6z/
LTX3Ngnq+rEKqlWaC6uyMsE4y275rtDVfEM6FKNSfBLQR0PfHHhAoxJk+hsSJiC6
IfswKlmmk0F/k208CjvgsCOA711DcGX0zdcJCS36IPTOEdc+qht9E58HZzLKZH9H
GZAyy4pQstuRk1Wfstm1LF9t4sbGv3O1m7wAXSrFIu7U7S/0c9clBgC3h3pxOwS+
qBgTTa2KRBUdNaxxePJy231qoyYiFrGLwoebpGIivJsHDrjez3bjLiaOgwB58FE1
BBq/6Ffgh5y6NwMToEFal0GkqKrwXGDNmaqlsZaQe7e5Nguy9VDz+b4K7F2gmjJP
TsCWkJXwO+2U06dkJ0Xg8gOEz2B/pLJ7DEZoaSmPKLUuhNSe+l/Std1luHytJr22
8Wb9vYYa9Y/oaKwFC8wPccj9uBWkgUZ0i0PlLZLLv/j0FzkYKvD0/PqnbrStGkUS
3YRBwN2TEkRi2tb9YZ4KTGspY0dGnDGvQs1GQO+Ps/y2k20ToNzpaUm8nUo90y6u
ddrXIH2ZlBshMzlO9g3Qw7scG7i9f65OtkFvq5Fd+fX4y7N9bdNgSWdSdWn8kotm
GSIlARjcI6uCGa88pCHmkTkA7xt2Z/t5h6JmJptOaZz1L6c2vn2xrDcGDCXcjqhQ
GZOTHTC/56XA/D+yX7g2Xb2BlVzkzhnmdBFsLIdppnFxjI8dkGvlmP15bm4P+zQO
ualfDB4SqYPT/Z1hwZjrNeIk8zzQefJi93LWjz/MO8bayGp2dAdillaS+bl509Py
ya8cKuWAoXS3Btpxe075XKC/n5mdjYB+yaRQGDSmSAFLO9sHUM553kbGd3i4PKJJ
NoNaoNWS7FizOHAGDivwpuLJnVz/rL7N4xEy4uGOxM/SZNOv7MFXlWHj6GaLdxXW
N9mOH01qYl/Ib6URnqvUxwmcbhTUDnPRbhmqcCgBVCXoRUupUGCEXqwVqNLgMJ1z
dg/XSBku62sIlgFWOCpPXCPFvtFjDjGxMtpuXgdwr4OSYdhX27GT0NylegPSOWKO
QrwVIF06TwifxWmLHCg+xfRdrDGau4oAFYe9LY/VW3t/Vx0Xm2sPyR0cVzNQnB/Q
ygSrbW+o55WXE/EDvCVJtoa/1t/USeFrC1ZdLHRqcdcEXBaLeLzjX+VX/mPdup+h
8zNJJSapWZuH1hYFzn1KADqs6OuaNV152FoDRA9GOA5dBKNkXj2pUDq4VwZlAdOZ
wHSkbtYax7qU5yMY8lVUAvIKJp3kq8h6g1RssmucWeYCgDXVf+7qZONOJAgVCdO3
Kp0QDXA4jYqi1MCwVdpeNjyatT2N9rUyy6FEI/IuquKfzGM42l3NAKdLIiEm0VZ9
JddWWKjcaruHaIxbEqFU0NrAI8T7AY+ahwY+u2jhDvl5E5Mn0jcNnKhiF6OlCOaF
pZkKjKvMJiDfsod8fsoqjkxq/K2+OwGLl9EKxVxg1QjrF6mFyajvLbEyV6M8aTxy
BE9cSdVi06n6wYuweTuVnEFVAR8mMVAp2mSAHEpzd0WyX9FmqA7R0BRAWoplNDel
hbXTENiEldYRT79rrFm4EAYa5l36S/iw0s7dr54fuIbXuAPkQyFqYSxEq4lbZyRU
eM8BtKcjrBcuZ0pglNjISsGqJeWfDAq+3Ep3oPqQySM3FjVnwc5rTm5REBJ8zeyS
rSa3ul5RFWyxFc1y+BLPBCyYN6jVI8czwFZUEbuTVkE496UF+2RoTx8JwqjYzUNJ
c3iQ84Ym7BybzISH0ChPNMcgyB7CHhiNEzvHYhdxbslSjmbYzsGphay4wAm3wGA0
PcVBlpNxkqwlbuPoygZIAa8uwNN0WqiqmqbXWrapjXoxuZIjDd52LiXBX2sjzRWD
cCf8dNbVq3UO6Y8p4aHTaDzJk8ysjPJpJllhW8eo2XM1Q665LcGhyvSdtsyZwzi9
QOw7Z5yZdgQxvSy0MUB66CHiNjrlcJJEwTdiECXQcAC4ro39XFNSJxCeXSl+6iv2
9wm0SEvwzBSd12zJ0iNsM5bGVvsPzYqf8Z55naqNO/jFUMDrdbzLN0inpgNi4Rj+
846JbaZxZ/rVgRYW4VrD/g/8xyj/nEoIoWQ5kxLVjMQPWE8VOiln3fcmapv8Ll7S
mj9jwEGG7ZgXVweeJy8KQNJQhSYM/KAffuyrMq4CvA2Ab0RBvCgn/reXNaQw/ac4
n19uyJEdNDxptwIrbGgA7DgusB5vURUinNUyRt1uZhgtggkTvyZ7nQrfWmp22JxV
1yxMYxY9VvQtJbxQT7YH9ZvUutctWymBcJTiV+ysOYeefs6ozdWMT3zouytzylBq
VO43IUFDLztY+M7jWyc+9SFc4x/BXD2TppPj0j228GQW0HyuhGqW62oFP4NbL8nz
WwOZaRJxEFTvKkj++pF67TBv7VYiRSQXdtkCO+/vH0NpBHRTeAergh0S0IYTvLKG
SJfnHPA7EO3MXCyX7VW6oO6D/VSrHFDOHQbdtzXqT7ENc21ZfclwsaP1Aphj2rqe
nyGtFj2SUvF+wDC2FmIC75RhNk0+Bqb3t5OQt7jIJfXmVXIoPF2JB3Hw9/S+xXr1
1FQWgh/QHheQttO/pn03Z/GyU/qGZxIIl9yinovRL5ItdaeffT+/qdeqCnyRWdWh
UBjVPxBidZKXF5AuctT2I/rXd2hYEOh2p5M6JsAPkma2Gda6YEuLUA5hCUa5OTrg
H++KUG/Jf/mWwcL5sLLGh0q9dt5qR6Wv/GORfyhdQYFjGcXNdU+QqxpYj28oh2W+
n+102Q1peIxVeqOMoQ1tfcxTVR1ZBygJaYZr3rYQsq2+Bbfvkpcj0Uy8WDGzppq7
VA4nXSzEqV/JMZ+FtXyPG5ow7/059bFCjif2OY1zA36rEl7QeXz6QEtEK9R2MuBz
wK3TFnM4i3eN9OO1qnS3AvGKRYocq3mB6ZnPmvXdrtOne4GFMIOa3E5YKZhMsJv/
Sm1IBdHbkFWnvTx/C3AZrvNGcqh4RFXSq1NptrCHqfUR4UAGT6tYx3hXmi8hefDi
iXL1qsXzYtVSygdgh0xBZBzO/Gnxx/SoMPSaKxQtoeJXPeLy+2q1XQ3yDrDhM3dp
2id8d6OboodGr4KgDFPJ3azNd+VRww5fJayzTfvk6mfmjOwxL+R0xFXzJKrFsBGS
eng0QI4lSeBD4G1DMPkgY1oYXtTKkAV9Qm/HyHm/P/pYj/1DtJSBv/zR3cKL+rH9
9wxlhxq1PGx4paa6rDo6O0fQUrRE37WihmRrgc8vlKmJojEXfvvYTPEnH3tqq/7I
SBgdYY8Ia4Nha/LF6oBSfIkyX8jxz0NaDh/tt3IQjgzj+OpzINRcaMkf8xnzsDSG
FywGNo5fwHOFiQ2Ei7HdOlPBhLJtTnBFH+2sCQfA8jFzJ2phziwYZaTXqKUz5pEw
7R7WE10PjGnQy5hHoFiCoWPAA0J3HYJy+6xqEg0Jp6P/HQoMUxe2NQkpjfTtMVtk
kfTA51T5e92CWTm/b5E5XYPry8894rHLMNX840Svznb6i3td1gnHAJ+PGFgNNF5O
XU1+ULWZugPew+7D16Hj8XV5CgOoB1oHQEt69HSmN8H3te4zShubvzgoYbpgevb0
eUAkHgkP+RAmjY4YJSt9Nwu8Ke65IoLrNqa8yBRovvCoZKCeMC0TmHdZQP8uXZXA
qJjqlmXYQX07MQXYD7BsrOBUP9O0PbyawGDOrVa4tiHai+UOUyztF/iameFauKXQ
eiGI+160tacU9acajOnlXcJ7cRGO7IhURtw/9sKv8tn9tNlS1Relg6UqRoz2XZn4
X+1/ygKOs6cptakR+BNGeKqX+5LI1DVfSyA4CTGaiel1GctEpTxCtC952w9DcevW
xGcKJ8pCrzIjqFxtuwK0bfu4YT1yXZ1IRF4ussdquN6NATUUREcPEWAnvzvaN+gz
b2v+PcIaKcC89gxu5cOmjcnkzRGzoG5jl+zOpr2KyPwIvqTXf6vUnuPoHOeIAzkN
pqXz0ua/Y9z4AKMGgRn7JPwDSSNgaaE81/dWOQsJNBV2TSkHZ+TWLBx2/WmTb4P7
nqxpG9v31k8bj+Zw/C8vTvuUi+F5eDr4KGpJhYvkOgMfm22RJlVEXJ8mOmwMcv8K
bnZokRQZgHbNLmLk0XQEpdNbWefXnTnTSyfJcy62+0tDCRKWXpTG7+31B+a3guMF
6G83gYFrJdRFmzuyk4913QAecyZc5hSIHSBAyK1CA4fD6KI6fBNzmOfxAeXlfG7i
p6Wtcp0mdQECo4I9R7ERvuH+I8oB0ykyKh+YtxSBgweE1W6G8n4qGytbilmN3lBX
npcSOP7//X3ZMDRRT3C/Obj6AKp1lolUbiMPXclPgczd2Z/ug6+K0kvb72STn8/w
lJVAm1vZcguNS7K/2SxGGobkEd5lg3BXALTRih2KPyNmpGmdE+pEIGjYiSJW8ByF
vhMXd7UwVtrH+4pZYQgp9g4ozgcnoIbmOIV51ypBSWkFz1sBiG38TWuz3C8S5oTm
HHQUin3VaFqSkZ2fFxsCvVskkCYIEEQLt/hqbQhUKMV1L9eA3WYlv10U7fpnnvWD
EcXh2PMBDAHKanrRf/yg/sU6TvulMKzNpaDlCVj+tCaMY7q2EUyPd6/NVDuTdNrV
6Nb6+mk0jKYZbw9b5vh/eyQdNsC1JoBGp6KPuSMLtA9yrh79HQ3AsBsUPUHZCCA3
YLqoP+Ee2Gnk0yU1vzL20fMZKTuIeVpOCKbojdNx6tdwsfFCehACBg1golGPxsTB
6qO0lSGzDZ7nVzoQe+uRvJBCxBxjZHvfvdzlwutK9D5y0WoqCyIsl+PoDrw/HHT5
oM3w22+JcUbwudC8gSa58cDGpVXuhX+TlkuY8fN8KED7GCwjV3yYSb8FwJyhQFeQ
wm5tRrKXmgcutLdvq51xmfZU2lTkj+xuM09TLF+pWxreQhO0TMhhSYLyCtyP3aE2
OOunpniHjlqe+CoJ/gmb8+gfw6W7n93CUmWJOp+l+hwTOdlpRmd4VI7/+zek8MU0
tJjgtQD4BS9auB96/UQRlZPwhCK2Sfwo95Wc8HYjcjOY1Hd//7tbAalp521bzhDS
QTqW+GvPvAmJLcyndBvZWDN9oiMkXxCr1yC5Ny8qF7WX9Y0jaOo7pcOA+ZCRqgLJ
k5knrk/6gH3BvSAfQ8LsMa83wg55PtIWfFO/nW5SOmF+eFNepdpeA516gZLX02YN
zkPK3xV2SVRx4ACwO43Y6ZOkF+kqu/ZYgdmfHSnZHDze3jDEKRImJSn5rzHBMG9G
po9zkbyNqNbxFzL/rAvYu4/j/oZAquRyO/9KFioSPyM6RR8KCZL2OlJ8B7uQsewo
k5vD0V0J+jzm/EoHVYTq08OT5dQ1OKSqDQFMqhRsnJWPftAirylNfvU6PZ9k9M8y
N7CmW7PV7qxH4aBDzxLNO6x33rX/eASBYtM+SAtYrtotYbRRMQusMDuI7kNXX+OT
GEgIpQq0FSeIh63yMlFP0dB0gy77un31kTLSzlyKoEt++WFgYkvuvBx+jUukWL4d
5pNKy/rPt9VWPmBEHJU9ElFDXSlI4fTeWCuLKrbGUtuihRCg2mVNYkMnD/DFw2XZ
lHsvXY17FJx0n/8rY4QQIw0xDw9iuew3OKEvEyWhLdmucPbw20rGfpT+L/GcptuV
tvtjRiRSNe5hYdl0ICs9x/b4/XVtoj2difY8m66fN87i6rARLVxuRB1JmfZijK2H
ZIjnh/D3LZCdQ9PauAA3SXPMfdz0LM8h4mrM9oddZ/vYLU/GhDCsof0PR44HXtpj
XsegzY3Szq9PdY76DQlXyKbQdRqPX8rgDoVwX1f5dkSKo+EX8EM+6Vp11Dp5VAoI
aCwYb89/SGjJpMSPD8LsEYCfenvl2SK5OecT0tXzPOIzkYGzKnpmju4n4fQxZN9F
t54VVtnSpSjY+AIw77IKYRa15cPCo4eKv5hzTj39TuFkQdQti2c9fGPLDa1/8+at
QO+eon0DqQ8I9dAh+cC9ap2cAjE+pegpQFrtpXLVWquPxnD6kzqr6GBQfr15YAy6
fzNq2ysJzFJkdJGQH3oeEXagegrHOZY0jTyozrHt1esw2ofasMpYsZJpFRRuTl7l
XKTj2O2Oz7X+YM72zX8MOqqCeFEpqewlJfr2shC3YjWVLgvNU0jHXUD7eggejJeX
49TKwgKbr79rstKxCvNrHXOCyd5GficzX1KFJrjeEPhQJJ/PPgF8Sqtadfi/n1HV
x+BvCm3Wv+s5Kq4K6I/LaaoamXveW8TNNqXsR25bC7Wpk1Xz3aMBMgVWG0U+LgAZ
GWZhzwU72HcRylJOJ5zaH6lgAwEZp2gLzL7YFgovVoF+yyLqd20xsvP97VnVf9t1
VeAQ1n8fe1zjwxrLVItDxQ0KUGSWQq76L0agWeXqCEOHqhAr7yPSkgcFv+prHUG8
VTAbQj3oGP8ThK8vmLmYCebVNYEAfBN4ZU3nsRVXaRhyaiCowWgwFNcHNN1n78un
uWMQmQglQoKdJ4k6ziOeAELQEarFixrjLuCSqna9hPlTvv75TkQ1N9uhJWQOP07D
Gwm6nt/0r3TzehyDvkzeELu7g3IjmDshCFsappbA1YvSo/9Cu+2SVv5JLUNP9bjO
Gqy67u3BO13cD95kjMN5b3u9lcXaPWdoc8I27X2A2xCCuxdUWiPbGY8T1XgascEc
ISHacz1n8Khf2cuj7aPVFloNXVRYfThvuI3Yp8gnPvvDEP7B8MuUiH5WU/gIQ+8e
Za0tvAfS60ia3SJqRA/3U60ozqsieF2NigCjnQg61bZKpF0X54ZsFTPpjFxVeNBV
AGQHt09w6zf/MXfhFOo3d+BmcUIFlHoaNoTZmkCmosxdOrcyT95DP4T2Df/jg8TB
/j8S7mWnHnZsgQZzPJ5Lhk/QnqsE9+nFHIuyDWAy2HedxAjNdfwkbp4o1yTWZwKG
mApJdMfvaDIgqdD2i2l8/CWZDmNU959TTDIYt6RfFgdB7rbwy+ttlZnqciOp0HA6
8epAf0zPoXrMTCeNBuWcZaJpHJ7na7S4GhSiwuvbVry+tnklDoeWJKwt55AkXdvT
1R4TzN4nObUfPqgOykQM0J8GdZIYbMPcnILG+XEIHZEQV7GLDjKzoiVlTJn4LWrJ
j30k5toIL1HXrI8FTDmgcDJgikYv7Ks/96SoiL1YNwVHU+LYSC1cvD27qcCg+WUN
d22toJe3pQGl+oG3elZ7ik+B0g9JsMcr36OwMXaE94Y549CVXpvfIspFFSDhh3mJ
D0DD1hpc9V6xAB/q/+p8pQTxUfrxlZRzbUiXt+AlQyclp6qoDiU3Wjj3UTfnHw9A
obffSu5Y+tILNX+YUXM60xNQx4zwk+NW4WEDPEEIgBfuOC37l9iEq16J7pUBxBy4
ch5P0Cg3OiwtlPjhVKsWb16tRgq2m5P+tp+b286O9V9w2qJ7RL3RqfKNGDG2f9k5
iuAa98qKQddVdrSn83nPmXX6n60KxVNd04dq1efrWAy1L7Xj636D50hmmlbBsLsJ
hBbI+fX0AztvkFvOT5j7ggEXm6QciVbksC1mANCu2Vw7S0xzOdwet7FwY+dNcqoO
A7AxCIBLPWmra7KoK1eUtDVnl0se+Rn2U0ntO7CFp+Bk3v7D+lnYsmhVEH4DwrR0
lLFFDvA3b/9rgZx/0lVY5W6iGFffd4XaiuZ/2SNAdwvTrRLUE4wwdxZfFTNvwrZ/
q2rqiRM3zkfMny4YZ7s+KkQUpGatwdxugKthMkn6L0DegKhVajegH1ahbCaGmyw2
BiGN1VmjOP6q7DjfeuFHsfUUp1bgDeBolkSNnEQ6aQr6jLUQNC6sPydsdXVLXLS8
KLczgMjPqKQsT6pqXKMj+n+D774sxpWfnp1SNhZmOPXP/dxdxL/qwnbyjnUwUQPf
g7MQ6YxuBkm43LaydmYV5tRQn6wXsBki1XfmCQTqr6NxgXgErLD3QyYmUqEWUGm6
Ak76cqw2VxtSYyCCjj7cuKtcYWdh0bKPy9QLdrdNTYtDEam3M2k3HWDPvtFWqT9M
/FkRLRY6Y6iDLEnlHo2MUthN5FdEwKUYj6k5qTOrIrMW+OgnW8QEfXt+vY6SEYTO
EKbP4mf0KTzB7SXPa3RK5nmH6BiwtGFHgFqxius32DB/LBeocl1WOdPr2mvaRtWb
/Vv7lIbosCmjsB6a8LqcHyW4hKa57RFHlww5SxCRtR+wDRrmuiksvq/gTPQBg9ek
mh87m6ahjSKthUr7TJmNkQbkFnG/dONZ3dO/wfC7M5echMGu87/FC9N+t42MEmPf
9X5xhFr5PIEzOFoTFjN/cN3y/dfJ/Z701J6i5rzSK3FzueyfaCRwkZG892rMsN1v
/02w+/+Ggtr0v3ygluBjse/mWFpdma/JAjRAWg3r4a4Z3n/yLkhf1oLveo1/IyoN
Z93hQ4DJdAHHTitVOREdI8p/k0OKiirGhVkSSitbMdINspv4yT9ux44BkieO1fYR
HmtYuqngxgda/ZUkLWn6oj44NOZHju8RBny9WHhADjcAP28Qqnh17pAqxaS2zl1o
LYeHanGAqNl2ukMlX5w9mp2CRvMvlZ2H2S4eac3TWUQYzdBc0saxC2GVlVX9x7rP
BIrCzXJeYjFCPXeSJLnFWPXKtu7Yk7K5s6fPdS9vcLfzwn5IOmRsiYiaaG2nnhLc
fJ5+RFxjBv1MrGG4LXrLeVAcN4F4JsSh0FSG+pSEAXfwh+kfFQnb8Id1FHhgnkL7
gW2JgUXRITp2kb4Orzu6f3au5XcpU/RcB2AZM1ptt6pfG9vjfRWReD79uF42rG5S
QlUpYZu4xGR8ujZN2uKxN6pdMDkbxn1S4wI16B8440xR9jLIDeSAO7tkXJg+Oa0D
/MhyqK62L5YBI0KoYCkqhJ0D/zjo9JUIxGeXXcYCNVnxoiNPtMF/5Sdbvdr24nBC
ZxLWXi0FSdZiVJQi0rNlVHROuul4BqmxQxEFseWhFhyCQ//bR3YPfLbQuhCieBV8
5diMsoHfaoyB5dK199UWKgSw0yiWLeIP5DCD7C8X7t1nqJ9dtMMfWi6vpbLrqxcj
ul0LCfhYRBoisyJWxwjO2ZRWi5KJSHKw72Ml8nA56Q2gE/pJtOPMDSf37z2VHven
22uNk4r1kiyc8Ta09vN/Ea7zjC/+z0CnIM6tTRtHBUPxbg2Xt3LnVB8mLUnpfLLT
kDeXJSLvIvBZH7Q91bvtqjHtKX3rgnI3sACBQpjJx0gkc7Ej43Y3RdD8TDX6xTit
6hPf/IWqzGaZhOvt6Dhy0tJJKMW51ykCPj5fVOFUy8VDhruOxMucfKyi7YA7tScn
DJDQHBauFNtM6ITe8KlAP7yU+X5nSMUgyd5yyVVnd1jc09MYii678wzLMQ3YrfD+
J6bgydQyubsYBrwsXz+Sae2JjebxKYPXh/A2AUwVgH1c5bGH4fVKYXco9WXtEx+M
8WBZv9kIY6isXctC8Ea9ZlOtcrYgy8cWrHjWlfF4CzKXT5Ermi5J2bPTrlh/lfcw
5mf09cidr9GqiGaq6yqDQu6kZKcR0dDEJKA6Ep4EyUk8tnf41+17SNMfZE8Jm2Kb
nhOO3NX4G9e9FAVxfHPlTjMBHaDAHg1BwBTtD7N8FRU6nJIJU9p/zqCIaNz9KI62
5MBtWqpvGgwTtxx1tag6GjfjOp9vr5ItVrT7dpPLhl3oJMyCbbusaMJsAmOP+mQv
jKh7m79+j8wY7n1SW+XUUitEyyQIxqBfwkUuaSgxpPqSgKQmLylWUfusp6uXr2Ip
SmK9kTO2v3Db0952XGn1TNxdCFjnNv8p68wagfQt6GkG/w9NSDnma753knLq5wmr
dtmPnGVLB/gJ/+I6mty6k4r622G7PBT4p5gDLenSW0Kau9daYwDCmq+PFuvnOIzx
Wv0TRWci4o82xcoLld5gq3ZmiRrfGOp7YirLr+z5hVlnc1tQrswV2ZQ1ObUmYCS5
C6popFVYUfGDKgPLiSCJjGqlN5xc2LFwK8DB3EFQFek+u4JuTvH89tFp2X8r1uoX
/qF3X4slZSqIlHtsUlIQeKddpT0bTFYMo8qZs49evmmzA4JPZrYP0hEbwJVx55AK
0Rtz7H2/U/E+H7TO0doInkCRavgn3TQq3FjE8CJcDU6NeIRzvu6Zq8oRWnDdYIuH
PLCm6LtPiJvRVF9qIgmJY6svz9nAtmy+ltuwfyhWIZgGk0rG8e45DeX0gpiskzYk
avbIo76Joq3OaCzpVNxJNzytXvmY8bRtbHTReSrDXGM0RTAiufIoesrifjySOS0X
jCTt0E3Nt/LghUBwRh0QUGYmNimmwbtuwmlMSMp0hHqsENSIGalsJbyv6ZRk6Opw
NZKy+guIU6WHLrbA0X7dFB8dD3fzb12wz/rMea1EiN6Tl+Sy+i++i5OBqcM/0koI
2gx+xIFdJAibO10ge/YvDGb1RuPmdUC2BCAbsUcLvxOyVYQ77RftrKMI7Pr6ESGY
Vrc069HvEBXiH/J+wHik4tFHGVsAe7dEIMVBDYeoyKsp5pbCtlgZJUIq/lYW1pdl
Y/9Qfz1p5w3D2JQcyKi/lHEAIjnGRfYla2qCuzTGhD0jO2PEMtEpTq7Voj9hp1Rv
usc+qGTg+rCNobScvrwbocOk2wOzz1D27zjU0lPctNfUesk/z6zoj9g/+xog7urt
99ZpMpzpkdpshGGHAsa2hbutXCNatjel42Uy+QFtgCNcLLpBYU/MRN8eF68bipiF
pPOPtPAaPPpHHTgwPrWfmL4ZudbwFmoLmgxKvFZTCWJ5Jmg/jZlIZR9X4uxkk8F/
XxOb1F3D5eaw7qAAvLGiCVFKjmBas52t6uLLf3sAn0PTWsnxpBGksAlOYw51Yq9G
JSbK5MvCjHgNMAIFNu2P+hOSgPZfUnsBgaJcUBIHB301qmItnNX8EnJrvEJ5mDEe
LhTiFqd2vAhW5DqeIMP2IHTaoaDUuG+nG/gXTuSAzGyHUNjlwffqc2KJenNU1Xrv
RtOe3hqjpQZF4qPa8RkNEmxCjMxidDQ7gkptTOzxTQKJw6Cnf8HISk7Tb53N5In9
R+PZWxqoGupxPZxU32WBgnkjQveKChT6K8JTDHkWm6nHmw/O42xrQqGL1l8SZWgF
X2g7HECxBD79kWWdHXR6o+eRC9INQIN2XGLGQYg7tSxiNA3Amz2j3HdWmGGBDjq8
zRNBgC/ly+7GOGl4rnVyEKswSdjfVBnQI3nH/tHJLdN+b8r6RAuWF0s/7dusJOCS
cxLbaDC+tlZZ28c9qNLx7CTL0uI1WPruqeHktk0cIluYvOOFLBEm05k6tXrzd/AI
7UIqb6chjxnWnf3WD3Jrrwfn3vlSulZKGCu/CsOdRLH847suSDJPWWOISqQnZTRY
6ljBqTLO9PrIu+KPUvJVN9ypXELyaIOqdQwU3sm9DCetbWH0V7NkEQWoZu6mOjDg
d9O15L+/88hYNa5Nm12yOHonyEm0Z24yRxAF5K0tpBns9EuC97wrL22NPVc3WWTR
fbgK3ofzyXar0NwwBwUdd9VBfomps7cRoNKs1s6UYfms2ITmoQ5e5l0Q2ZhgisJE
4b2gmnreDziG2LRNfmjhBBUmKbPbZoXNc+5HQYUrz6g=
`pragma protect end_protected
