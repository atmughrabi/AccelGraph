// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Dt7S9JZF9YaZDOrO2tdoZoBVbp5Be4Mi8asClmz9zNUorehDvUPsfZHLw5f/6U93
uxG+gGSFa1OHXs40feSuFg6uK6IBM23wU3QC+qDuDBahySpqZBq/ANUQM7MUdMxr
cNSpM1sdKDVQwsm9Pn2HZB7+mzYxGEvWPRDDGujTUIk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23248)
olUzqWi0vDxsEFYJeVgiFog7K13szqSmogWtkXU5p7U2X9ZToQF0Nyep87AUZHzO
ZI+vZ3iBOs9FkB7zVyO1zHvSMoOLuVELa6L0kiCeuyzwFIDIEWI0KWbRHPR4zLSR
2n9h5DO6CD3ViMUP5xrn1TnJ0/ePWi3jIXBSaI8IjMWXbnjIMsg11k5OWLyxJnVk
QWb78U47r9FkbFu1r5EaJmAPoq7j7G9jyomySJcwcEEPNswOqshhkq7q/4jChDsf
Qc1bUUYLqSncgeuLij7muVKrL0sGIgykq7VnAbtF85obZYLw2fjpbQ+xLtxP4sPx
u1j4NQas4nBwj/EQU+kl6gfJwJoA5nkan6OOcYZwIWgKo3VmbJoU6Pd3R2hmEkNR
RmiN2SLOH70rG2DazCRZx/sWBeEZ6J3RmGfOgV2XyQ2Yr8EEaxg1jEgHbvYwqlah
unWuhXDYIBFz0SsF0r628pUGnw9qev6OXQk4X7KKTnMe8w5XA3Wk8t3+WznIlY5R
SxQEEAF1UV7RzM40UoC9HP/otIK4aii4RGynTRmzI42fJhGL6MEwVBNWjjae5/ev
xO9yZLTSgmwR2ziZicMVUNxdL2LeIO1Q8vNGML9BtOB2s+8pWcy6vbHK6quZ88El
rDeGdjUhOYuPX45MqtX90SdSJB0kH12RAwzTEa68s4M1i6TwgSKnJh7zawcmo7L6
RhdiN3s2ZsHQQkCHep/m7+w1j4gtmQqOlDtfadIUARmRUS9q/8fcFVeipCiggjBS
NLvCBWe1l9vaNShZ564JUg2WywrfmRVfNyiwIA8N/dI4F0gYjR///jDgvfNxN2hF
TJL9V/Sma6PugjqeiUp6Gg/VrlttNA+WF0APAEZrqEqiqfbypejb3SuVLOewV3iC
UPdzKXxCoLFa03mt5IK70Bayaa9SHNi7QVkuBnZ4nmNDtpX6+nrLJ1+7j6kkMedQ
5IoitR4HacA0Lihk9uU/NOgPToy87Kw3Y0wL2LhNZAu2PEKNgiI5bUtmuS1NG+0b
LzPJxyD+PdmgKyT2q+USd9CYIJ3AVXpGs5V2qR+uGx27o/mHp2D8tuVD8MgMu5Iv
hM1jDAsFRSRRc7o13oro6kjZ1kOrHw3tyOTj17M3FPhgXiRj6TgmCyhNmSGG5V4B
5xwHZBrv0dC/k0uPkjz1JNL6vvl3vkABC5zhzlNRU1Nfg5oHJ6B5s9Se2KjEf5tZ
KfqqNaHWeyLbjkwPLCj6bs3MR3IFrh6iVZvImoc3Sp1E00gcSL+idsIPTf52yMFm
FQpLcoUX6MSIBn3hxguaHqNpDyDmTRQNb+4XyJmh7JhDYMd22D2FYGiS69Cp80n2
8ietAmQDdCJcnuJ2DS+3aCqDxIGi66uvjt0+Peu8LOA1zY5UHLnVBVSEqYXzPivv
AHan02TWR/hzRN1WqlsTfpBmCZ/WitKTQ3rXakmzClua3GkJnUtQRvDqPHgut257
Wb3pIYp33ZQoWmcjkgKc0stz2c3hVZiS/4bUVtCKnJw2nk8Tcb9wU7x+YMNjvpER
PZ70kzC/Mqc0+gZbeRunqyY6sNJ94QIC/dtqibZ9GD1kDtGDNU+Q3RfdWFyTFUjD
Rl+Ik5XNOaR80KbyqPlABdqXhqjix1zhhtUMdnXWX8ZtX0ffxAy5M2aRQxfWYgTb
xB/q6+GY0EF6MpFTDAu92vspW8EIpqukB/BDxMcuYJ6EyihDfjCT4n9zylxBPFoS
WEuAjr/uf1ieu8sFd1vSUjQb+R6rWzLmpYy1/Su6hMVzaYCaJA6LnPndKVowLKIh
J9yvCNoK1k1xcVgEh1o7HFWKKERTlLpUjsOIKHXrhH5UZfq3vBbh/13bgPj/Q9DP
zbO+Yd4PnNQQMemniUK60s7NGbIzFfRG4ud3eQsV5t0mMX1O4VnOZkJLJRbOx9LB
Pj1Ls9SRBryzTyqoI8ppe69Fi6wLEqdVUHnDpNYbjfn5i0bPF3EGSVXEaGyYsWKS
ZO0++VH3F+5XLx6VOPVngw0E635T4HLVtqMPkBwX12cEoh3iDszUAt49jTGjdbbZ
0Cv0TxLxjmUqwyph40Jt5LJOns1y2dEExqUjFIBALbITO6RyQOlbiesjHKo25KKh
4vPIiPyHv/X46BS+J8UvMRyP1SPkjHIbWfstlUaNIW4Xy61XH2qdrzSxveLrobWX
dwXjtQgehvZUeDGSPzgfVd5RCQ+6nTIMJ40aG7HHpJPs6RorRxsPuqc4lDz9hqYx
O20RSL29gwhOGS9AuDhfcZWpf9YKMIl8N+m9rFxBtIUhQiGXuWx962L1SDN1fH7F
b0GtsebX+CA0OMPolZIiD5B2JibCsxLRWkAlkO5x8EAc3GGc7AdpLkOzz7ZwWDDJ
sQvBavAsKqkdYX3d5rLS7GpkR3tuzphBwxmZc6sNVmaKcxh/aqtBMKuiH+tL23ND
iFpheGe3Y/J3CpkyVyofrVTo6/GGzUzSjUCs8vcQleQZtheXex9Uj5IzD5m/Ewq2
1ob8jns9dIY/XYa1wVB0YuR0t9a+3wiaWH3Ldsnkjx61LUZ3MpqCWysi0BWgYeb/
VKU1ngngaoJlPHSOpNvZpQx2EAHl+Us08d4Q3pESvO42FdsY18pgYIhMLBmZcf4V
e4xetgi5NgvM1JISiKAvDQRSmmq9etp7OWGx0H5Bki7g20Ml064OWVMUgAY/XsK3
taDVIElixM2kYrlJD8KZ+90dyYdG9jT6K9iu0+cI/B979Edc+dEkP0xwqvHN4/FZ
CmnZkmFXCX74KlssSJ99wUjdQYsSIA44iT2RpN5h32d5utlrkF2dBPvp9QXTN0vO
wmMNP+2NHbro4Hcpx5lLViywbGkdD23dEPyFzbP1NUysJrYhTfasZ3+lx9jnRefa
RfI/NrSF+lhZdvUug3LdjgWU00jToZ/HGEVBv1x4uHNlFyvRAqAwKZQlq3u9yca7
/L0wR93m3cXWLxvEKo7KqZAZkcxG+iqWaNFLkrGayma2XmVPU3L4Mv7h15CcDZtw
f+HedJLSE2IxNcEwzsxOEOlZJD/Nv89PNicmB9+0D7HsGuz1gpZBa9dy8CWw0K4J
NVu8X/6BEejWl8FP6fKcUoIwQ14VmfbtN1qdK/jUqgS6av/PNoTsxfZIsHHMgBWD
47ozjGFD9+buwYJe2aRvQNTkOr7r2uwpGpLIzXLHOhukAW0f7xiNWb8AY1Q80F1X
KLBPj5S00XgCEQcUHWz3abxLWome2FvNuK1kkxcXRn6eNwxXPMfomjeyHApECc6S
JQrjN5RsZqbvJ8JcK8FYdR9NtK8m79i2Gk2tld45bv0fGj+JPNFQzi4Vw7vDmxes
7sm8BcwZQ058gHd2HsVHYr740Mm6J0Zsu6eOVPXrTeLyW6m6b1ajcxdy1wok8T4q
9jhkX1T9irmhxdQ4op5wjBIwmhJCeqHFSCjAjwL/VAiHP90RkuaR0Urn83QzFc2e
Q5dcab9zQcEmrPDMvSjyysl9N4pdsJdJ43GvOV7GNwYkak2fFhmqn17Y4JTXTSB2
nqPRFPvKLMBwJ6iGoHMLhE6Wtvl8gU01rh5VwX9wg29DUt+pHS19Hgj6qWezHiIi
xLKhoExU7vNyBQ8B6svV0wUWIwWQeEbH4EUi2V7+J0g0qwwBlls9684l9Ibz1CQJ
I2Vo3rrA1MeQweW5/PpF96Nf9l0N4aDm5RhTIOwfEKyCpGhjQRb2+QGw9TZl/sJZ
tNMCuiViEJLQpPseTRVqxnyJLLCriHTLndagOkNlc8bnX+k9Y4/3OCFZJjtlGMbS
axQwA0hQkFRiXnFPu4jA7dA3KWocrrHh1Xhwy6UfrMWHA0IL56Ar3p0XK/MD3mbO
LISvs3RsLlT0aFFpZrAV8ZIAoetRqMfA5BErErtostMjvk3Rg3QUleP5i54fa7xs
EdvfbILH1y9NamdP6h3lwetiK1OrAENXO/Q7vwFphEl8nRrpBUyjQMHpBMRhfEz3
0lSSpl7FamuB3ozMez7aX0kXkc5Fte6U2lRPuti7RLKtbi++Y0eYYoenAZSvyyD1
tSxu36C6f7AiJ05KmutFaNwBKFYUEjtRqcGQa4pOJDRF0aK974ZJosYuym0mY7PK
UOdLBji/hEZCuPiPvypFdCcvgYwpoBaI1bjZNWAx9nrSIwcJvyBtT9GAKPj9JMz8
70qabMie5qsa9RF0u35owpUawcNIik0QjEj8FHmP23RyTQ4s8RaN1kkd0gs+zAul
5N18DDsxvwc/cXtYyiGjIIpVuOcdulgCWalyFo3ufMHjbl6qT+BQJqOQ1JJcQduw
Mmbt7H85z1ppyk9hqyTvc/L8hfFeP5/gD2r2TGeaxVnetRt2FkzyDuSdiXatXwek
FBqDry1Ey8hXYeDaAXeagUGuwKA5fn8PAv/wt59W42hM7BVkKROw5vCc8MVLUpkH
x51Sy+McFoUNr3RKYoXZf6ibk/yPprXWwVSwPN/kyCcbBz5rhL1SuvCi2knCN8f0
sPK2tuPeXLMNcHFy0RXXto9QQXHIIGy+OJIDNPTEYmEtZyReloybQxnrh/aflhEW
b9CM9S7jVU+JnIBmBrpy9VlbBXB24hdFcvfmIQXEJ0C3CWu3bX/G3r30K9h6Srcn
jnnHiqTffYInSbSRs9ctc9ytTdIGhMUdSjWmcCkmnwLay/cR4aynFv9/DIvd7Snz
3994oKwPf6YWP5uT0rAN0jgafW41PWXadDogY5OWwjq9/5o9WzYJhKxc4u4Q3D4E
E+ux99UrqgS5qPDUEwvS3HsepFc9/7Cfwu9/fzi3CU8K+HRpKwbRqFu4pGHJ0sPF
s/go//ZDvxLPpalOLQJ1DDd0q45iwNq/7MGfkucb0UIPlJLQ9t4lxxCNvRFELTvN
RP6ixM1BsXaaNh7q5+23/WNgeWqBeJX8EWYR2zCH9z8Ixa0/eBWXemRY3u7bjCeI
DmfwwH57L6cj96Rn1S0lFYAaP1o+GqntGUV0xeMqQH1rO7OtMZAILlKzrcoyZX4T
wScNBeg+5/x5Va31oX4HM3sEZH573ovknMv+UNsgLRr5LUV4Uu7TYupjiaX1wrkA
BOwy3vOu/k4ayqMvCKXKjqEwZAKsZQztIDr5/mbfH8LfvRxS0QiRoUR4tQIT0qBV
5s15pdzQeRsuMXd1hIiLA+h+BrLp3x6nACHNK3STl/+jSQ851FxTiy6eXMGJXiZA
mWJeMSMBdFLCH6Pqb9E4uQf81N6rwagvraF8C7ONc7/ijbNKweQ7VudAQOldAsuA
GEs6cekjwXSdJiD9N4x28e6jy3VseeM1Iht9qrNgWLwXsvWEdwrwumNWob3xQnVl
Wtc2qeioEUm9BSDtfaMVLmqaWDtqUTf024h9JZ9Bg2l1AaMnCLzt5I8hPJpqPioI
PA7CgO1AHYxwddKav9vezDZf7q40RhxX5q0FV0Vu+QPaYV0Z4rdAvdpJ/qdiJYUo
NJg61JA4dK+EVMgOigaz4MwNa97sOLfSaousGVjrYE0M6FlFwQNnkSuLyRrpMDGt
iTpTNzlOdXfiezGRMGQcE/Hmljl/gN+zeoG9j/1oxMAvViJcaHygzyz4OJS8QcX1
wImd9+qFQ3R4MhKpfGsWXN2KNU33yfmqtxpqdWn6Yp7IR8yxrRCk+kscNzEcwovj
ZFOxP6cxdLXwPGKfLniZxzcFDSzmXS0hXh/U9CATDNTx5My3UHDzMOaIYzxGTXHa
aNs33/oB/c6l7GZh/wBGD/mhXhDw68IUE94nRjvBXsRmkIAHyQlR76AD8VFdqYW0
p3f4p6TEk5TG2Xo9gH2OfYR9JnG3riXm4Q3jdeguUZ7uOyQaBjq6ZoP8BRVPcqsN
F32DZsONTvReZIOmJIUW11DCQttXHFMlFCDAKhlUKSzsRm737s2GITUzcuHcNSnH
zXk2VWl2nqODNpZ2iNc+/aLGAfdR+V0Nd0QZxYDQH0+69vLFqS3yrRcgzXxY4jEy
RQst4160fYWuX7EgAqduFaI4yvUM6Mm2HVXR3TerVRfT8K8LuIe/xzNKhxa+rqNp
GClVtyYdMX4TevFllsP1ZPxZZOYTba2hO/9anOf0lXh47iC/ZR+vtoqT0+ZCSCcG
FqXwQ8iWhO9pVL2TTCAkxwVY0+7uZ1hbgJLV2sfoOCnPtSLf0GrtnT2jZwb3alX/
cF7yQwoqalO5dBgqtu2ncwGnDrfQNDB5ZWotFX0p/Ovtx2MfZlQMyZhKaxPHkKJ7
Hpd4e1KksyaUj7u0oBHkD2m/IyVcwU/qGW0FsA1E0IHcPD1HbJtja5TyZ/H+40lu
bTVvVM3Qrq4EUudYKpdYZ72rDVtKc2EZEylcM8TqyJyofWY6/brTBednaJ+uzwpw
haz1JWrgmi+eVw1J5vtbbPRsq6T4gqxteZStlorQxNAXiINvPLgqDsc6dmiJvFkD
thAHRiIH+eNNtY97Px9RB2THmt9hpdvGvCr4nph0JF0ewf7TtdYtWgpG8nSI3InX
RKQ1Ztnm2qVpxCS/7sTTjk38s2J05G/ElhWwAq/rwjM5UdSshuKcS6PtO7/Ddsa/
bunL4JLzp82UHg2JeSThYCWY1tmglM2evlHzbSGkbb9n5NbsnI7rRHwhj2PTPYvK
jzoseZjZmvqEGntLs53B40mxjhvPMFJkcK6MTcz7SwqwrMyKZ4jppAtR+w0hhAC4
UmBYIMUMBw2oz3ebZ0e584aJ/MSvPUXjoe/hTPbvXkCgsQHC6Qy3Muf4TOfA0nBE
LzIDiJamqOuuzrtDRP3yDzyy7ZxsJAXUUAWxYAxjz68aWYyogY5DXwrZMfZ0r/ER
EH83p1tRsPxzCBdq8097CZR11b4X4HTEa2cqTn+AeQzqq+/Uifp82e0HL8DTiJs3
EtlUZvAhjdSa9yvDSI2sRc6OHIKOv5fc5jC3Kl+MnxYBSbpi2QZDeCMXsUQy4ua3
cZBuYHLYKIft3uAqiPTVR6sPx3YmEZHRJMPKwQBT2PUuSmrfDWPMeOjsxnmH1nr0
fUmHDv0qEjidQV3m6a4x27Gn7mlods09yIpI9c8ICW/6PMmU4p53i4/kroY2mDtr
CvmvWyge1xxtJtoAFi+qZMHTVkc2BB0OlBcB9F8PqcZ8AtTfwoiF5Vzr7sNZsO4u
ys4QFp0/kbHE4u0AS1gemSZLuAozNGIpAWGSzidFj/an9c+PWtXd+tAUsFDbyhzn
qc5WQ/Ysz6v7ebN9ylT1Hr7M6koDpfGJc/2GSGzLDDjJV3WQintFbv24MtQqJBqa
ys+27+HoldD4vaYjshwoa+aRbX910YmjPUwOytDOAvj+Mw6IN7sh46rU16wzlmWD
2JeGE1xaIpG5je25VsTPCr7IQ093w1t+m4Egv4Us21WJQruiMSRGaMxu9MeWD2Lt
6T+Twr/bpTjXqK5YUsn6EqDERVzJX+ptNwtcCu+a+Ty+tW4CwhPAFLMPkrjKiB2n
l19WRfJIuTtlcjKeSYqoiZzRw4L+PP3Dnr5EEzfQI8L3KBYqUkREYPWDklje9R3y
b/BBVJ4nhVqa6TaSfGBgH5i7GCCYvNlTLZANW/xKeEq9iRVmwguKCXaJ8mJXMRl3
s6fDgLxTkGQ6wXk2ISEgMGp9d6mY5VrS2F2TxmUdoNl0XEC0v7Y0cHsBlgxjMTsh
VXjeGy7/U01HrP1AEAj/0YK9vaQQtusfen+svDuG0pYTiwjZm+RTTSvPdSVHe5Pa
IJP8XvPaijPy0g8L6wK7s+M36WSAXcLXJwM2xEwamm5Oz0SWpNb2wXPoz/xIA0eI
SsiYRvdeRhOXrNUrPxUs6JOR/ZG+Dam6k2y43AkK4gUHxG9UwTXeV+EWPgJSlsrS
u51yh73FoZ5c493HAPvQmrwWGIyOAyJozQ70f34WNbc9aDc3ajqbfdapOFhWbZI/
e9led3hDxIEKpYfwXMXkCRSSKj7acic/R1xWbpzvUhVMoEZayu8zuSoLoJi2+G7B
pu/lB7LjPw/vALSpNEwRJLVv2mpqAaV7ZzaPtFUWtLBLBww0inek1e3o1/e2DGEu
wsLLRoVonWhYloH4U3xOUphI0nimZXaCF+2j4LbttKJkW85U9C2hM2ZF6GQwBw5M
Feb6GrksUUcCRPP29SP5OAsRFIK+VHiSUaTb2LVTaYQs/prpurTvlW5KzgoMsKQD
CxO4MEyoUbIpSUmFVSHn66/rYp52BI+zV6/T3lL5ZeQLDpWvR5+Oomy+pDrS6VgC
JedtxdJaNb7W6y0kC4/S7FmdcunlbqBdkJeswDixWDNAUK/9HneUPeK+LtRDUhTk
0vWFQgEXPkPhc5PphZqiFqRZ7swJuaZGOVbwE7GxBaQ2lq0MgcElfcT1FQtF/RCM
kJ7ZRGm5XQ9vsaYpnpDjFXOJSuEn+u9cIjo1nx9D5aDyK57NbbmwdeLF54ClLr8U
7gqAaeynykypOHK3WJxoIJk2HjGVwjoOPmyFsi6Fuxp9lzBd5ukF5p7ERnQh/b14
+SRBhkLIELlbtOz/Oz1rEVGb9V60sX5JApd+Dtj8Rb0OnCefucbsq6XWGwO8fBjB
0gUUM8p8usbZgPz8+5CPgTqTGbVnR0Ty7DQMvfeufEwLVuQsMcRLwgKLY5VVpb3z
dXJHid+lvxLjx0MI6t/X5F1d0GfIesV3eYp+uzsl3s+i0iCT5u/pXmiFNEmiNP72
/UHYOvLSduM1yJ0vH/FTZViG2kjRMQlpxADWVOKiUdrTepMbXDlDH9RQ/Pi8pj9Z
HiKNan0kXnF9+E4AwAT//nbR6nq1wqR/cP2sCgjrDOnEPBEbaXt5Rr+JkWFxxtjc
Iq13SVHxJR3NEBMdcJOX40me03hJIBAbv2us33WTeULP9lskbyxbFcs6bx/XBFWV
gytQn5R1q9X0ooAA08kvhzZZoEbAd2YTtxFb77sTwLOdmgRcoiAWuTFupngOov3y
VZJRx4K0dAFq6XlN8NHQ1tkcwMjpsX6v4VLtNtxs0eQiIS4grN3n0HRyZtPinsMa
ve3mEZmeku4Edua6b2+mfReYZwld/OJIPSO1piMx8ucrQTCYOgCSSz0W7Rnbkwj+
cS/ah8Zxh1gw6QwQyEJzCifpCbRkZgWPpb0uMDdOISKeYvdN4Vhr3gWJxnWtLZs6
D8DfP56LXPp+vG7V++4jrV6bcIEJT+Id0h7GxKWaxSffuYVG+wJ7qOePtoe+IxVb
GcLVOC0yNHrjx8/C2viQs6Om3MXsTcDBX56eBrGJIKzQt0jP0HuigDmIQdr+rd9s
u3W0YswfkrO42sjtkGZ+OvtRb1Zi2RpX7115lWwXF4zOS6jdmnZgJqseNvySBGlu
O0tiriwteWm8eVQr6yDegsnmhuOW6T5w7i4FT+W1nhPGVeEcokYIglqcsHR+9ggk
sj+UAz6sG0tULbyioXqunTHCeuXvsHWE0gA6EwiM+s6gne2mSIdiYNCUBYt0UoZE
2UNsLa0x8nrXKRGO4zJEwjEMARTSYjr+HQqSWO8ceZYg1Oz2/QzR7dH3T+o/aL21
b2sVWGbXiHWpjsw89Gibbi/FDGCS5rZtektfNtiWdrnqnd4MK1H4ThnG0YM1BMIJ
y3+WlL4ibU0yYOLBVMqGrVoFW7sPdfFUmKcbm1bS0M39pqumiCBi2AjfODBrat5w
xunZoiT1zNgXYFV9Y9t2aK/5pUMdW1vu46fsn8pihsYrnypecg+R/fkH/YFKMvtJ
G6CXGvsJBTvtTXPMBlen34iD49oJeQXapKnnPufIafdKDWpVUosrlQpbvC56iR1f
H83S5HVjaGZOwLrKPSFxiPiia71EC6mkzw69Yn1YGld0BRXdKjKzgjfV9GObuhrx
IlliDdR8fah3z5bq2Ejbqvixb1659+xktm6SNnh9C5IVTrAY+JdrF/o28kb+jsX1
wCDxo+vCU3wlTHH/lKTNTpOs2k+P39e73iYMDrSgLcUYo7xjr9JDCdzQh2OkPdcY
c4lrBtJWUicc0k0jXpytl/pMJRCbooB6Ogu9XHKiTF8r+flEkMejSWlUY9S4lQCR
ETsDXlZ3G8bmCHBZb+xRDg+BTQAbosDq4w+R6JsOvC+nUOlP45U9AmpuS6t4Ozhi
XJb/tz7Onx87t9oTKBs2e+UMdAt7DX+3DU3QSB9gzQryS9sfqK/Dm8XY8rZx11ED
smwwUjrh7o/oZU6GgkXta1cDNGrR5GgCJ37yjTcwzU7fz+zsl3Iu6US2a+EkhNG9
Y7KegPTRlhA5f+7zPWdRKXx2VzBbnS+bfWo/luM3RAFWQEXR7TEy0i3Ky9iaQW5K
hYK+lPguJodHPELVLb+V0vGgKv596mdniywYt7nIO4RlVTJ2GzSSY8ZBIPCzWitN
JGyXNc4w2qKwRU4uiMMbiHkqIElkFpB7jp1Myixb7UW6pcTZo8SpU+qxuDY6D0FT
V4lTKPQ5K1eHzXYFwTnJO3vChAko/fzy3eNxKLxAt55jgAw3wZ/ocbhzP83Co/RM
55aEOQ7nUZMw6GxOTtqqM3yGIm7Awf+klwEyYkwtXiJfQSYzm6u+EGBIDJhmRY3G
Jl9JXQc9sAUqdbGabJnWtbNAwH4aD9gsYacfmhFCd9qedqlQ62XYP+NiF2JjdbY4
lHbXQJZ1PTeAx3SVugVwRrZ9PQgY1uVclPMCW/HY0LWg0r1z5sLuKAAcx9RAWO9v
cTN1rFp8PljmA9+8IeWcZws56To8moLE3qJErFNWD7ipY54PZGEVTJvArT+cI44w
rcXZhoXu/FRmHUkLLdW0Ce/nKuH0pxq2ywd+bP/k0JLnz7TWjWvYPUPDV40058ZK
zTIlRKk+7GFIfAQ/KqB3kctgM2pJPe3tarVyy15OtkDvftL3Q99x9yOb0PeqrMrY
LSD4Sn7d/NmNzMsqubpQqNMKChifwHFTB7IkdiVSEIern819yeb8KhODYVERX7Yn
003Q47N5S63IXnVfDjZqmhF0UTZpA2teKioIAgSHEVlFAjVg4LIautUGAQAk1rkp
qByqRus67hbhgWLPoQ3YriE+dhz3TnZOtTDeDJRHch4l4kXFtLRWjYlYYcn1wKp8
F7yjRhSG0zN8VvLc6EqyCYERqKUnTevDv6kc0Ek/qQXa9IgpXj0tCsOCNHcwM73j
e8lhrfxD/ArNnD62fINujmFX+hF0u6SO333I4JbiOJKpoqGzf99pDHVOgCx9yBGQ
SQmMd3a6wXBot+WeOmzCwG6i6Uo9i6lMw/n3mYbuaCi2UUc49jV7+N/mkynQeobS
AJrAyTGs21yWFbhnBGTwJWvquVMnKM3FKYDgMivN/h36yW6Xp0uRT+nYype21Vkt
H6XD4ArRSrQmgYLDdutufyohD4ELM74B6J+dSKaUTQhKEiFGdPWGC8ppIrm4zCB/
cziLWLwFiTlt34Bn7GVhVLOBwFHgnJbSf6TH3vMfgcNcSthcWCquufcO4TW7OaE1
JPqVrzEEPBmNxIv+XuTcdthaKhx3dBCz6DbwyVqSjDFz+UZ/UKIFf9Z/iqn/MrH1
OXW/apTHkNog4+W3YCGsaMhKz//FKDvaJayF7Wft83Iw+1b+WpAY59Zz+KDA/Ec2
sPbzqrqIeXdwVrPRCXQAeUmN1IGT68Rm1CXwfr3ExdsdIq5K23IfBjIPmJoroSOt
Njn0izp+c3p7QsWXHO0ELpPVAjACXtjwBYvh7VuoCTlsLHG9QkyEjE5/cYDZY0Tt
9dQPqJ2IUV4EGIeUMAElrqxdUgIq28D2s53O1K7K/+pm/UJtF8ezNk27iZRKjhCg
n3MpdJD5zPcWnWeog2cDFa+jxnSptGXy4udRd/LKt4UPlUvcv9v+5L1p3bClTo/A
AiLFJ5skC32JOUBZOKpCQXGqf2pWR0NXfDLvqExJMm5+MhLEt0GGdRxe+kxknMG5
Jmb0Y9qdezXJ0OXPMkTCguSMEkte5r6i+ZfR9OWBOIllGTQYug8iXec+U+HvX9ZJ
p2MY+mSbL87eorIeEsc0Ih/ORdeFIt2YYm7SYTwLnyP6KXx9kNBN2ufYjATrqTjh
ROsEMoIhywSnH9raCcdjCV2W8baGcJt6McV8Le9Td0FGH6L70/fo2QeKmpU4de+c
B3v/Mg4RWoHhviVj/INkn4fXz+e4UTYU5bqmvJVVXkyrcSWsqk5729nkYNq/Mszt
VZcQ/o/CF746SszqtGbLmpH1tt7yCiH8HKN+5vju5yC3gsQZ1hXeixB8kW6DmHJZ
4wC58k3M5QnKJkuvv5WBpsGmPU/C41c1gKgzPRLzUYlL2OIWW1rVHDgIy9aV40Dq
caHLr0cw7mi568C18Z+rJttrcEIpRiLKaCqyiHQRkdDanD9IRgbUaIL/LkBEddgO
C7MasCEs+EXNzr6QC4SdTlkGzVoUog39RXZcXNhSATZIk9MyRwjFL/P+L7vsxMjm
ADE8YV/KtKzYuUQpRbI6IatQR5W85cKC/nsm64gIfwn7TUyS4tTEQV/7I63PKmXd
Uah2qQml9/xeHXXxnN/f2qvgcoYruFvuCItiV8bQvL0np+aJupQuQNyzvm66kmDD
b8MNdhvo9ROphy0+sw7iv6kQxUGQK5nkadTo2kbKoeknmvABvRrRev7589MSPyY+
Y5VRGHfOepbHoJGlaiCjdM3vMknJAhkwI65abu9yq+wPjEzndaqtAcrtY5p8H5Ur
dofgRFlY02pJh5BUkIajSt3aFUJs8+dUgc7kRw0cRtQ969PB7aYvIABi/mQupISD
XZbis3//sx9B5XJhXLau4N/EeIwt5ToWJAxoFKQ9CRvFtP+Ten/tEz67XbXydMOk
4uerD6gxNcAWSXeYWC9ex1Pcgc90jmTnXclEmhGqFwXaokHHhPQkw7i5YmoPwCdS
P8mAbkeWngvzyRRZ4bqsAnY0rcdItrJiRX+AUmBsiBZ3u90xe7nf/zV8uslFsXKw
sU9kMXMaPaNE1NJDShbyPi5eD9txsQdj0VF+TUTpswVbxcwbBd/Z0E6gw2+3cYmz
ZKPUMmwYez1gxDtiAnJVnqWDddgEogfdTCNGvHuv0QRRt0KXTLsdTkmSWxlJzuVo
MtG3J7Lg9YIuuu7Jr1p0g4FiC0TVHAeYuW6+aL4GQzFxuRDyVMnYON07M0WoG54v
OKri3ZbdD2at7FsDwUXXTXisP0+Tj+7Qb9TP+O0yUtttWdxXMpBvHNCeoX2uU9Ir
fzHUWi6WhRx17krPB+ULMXDKNqlp3EigoWiqYyaqwaMBrt9NwXkEQUI/32WiAg1o
BoYm70ruMLinYLfTJoXjYQKdRcgdYhl5BTjiv0JBd/DbGd7EpL2lFCD1E0q1cxoN
eCxOMjbXzS+vLZLiQw3V5+lB61FFXx2pU0XUjVpl/D4ey6YYxkI8zjIQVehn7ZUi
oGavIRfWVApZMLOYeID13+qYBMMZHsLaae3w7GplLkBGKNQBD8rEE55D+HeczNHG
NznQhpEKxU69QvvX2NYUCU+JrYkvU3KTNwqrGt8QWEXRytXEY1t4laqyCisMI5zX
A1S1amUuVOrDWWfl5dzRtM2jysaDnfcYLZ8lX6R7cfmYQrhBbSXzFiZWiI4iI58Y
zNrDzxutDPvDWc5Zt5jzlTf/1h0fnemgQNwuKOMIFVAwPbn2sPQJpQnK5Si8ZhJx
+wQuW9Mm6cvsk2IPvYP3AJU1I7vHqc8+yBJ0oMrGVNaMK0OxyaJPbxvYOQNBz3km
4TM9WVjZux2L4ozNi4yzptWOj2KDkSLwR64tP0asj8sk6hVD/fRuarzBoXHIODiL
TojPdrr4QdQlaAlptHHSGHV2LWLelh6xTokR9zkAoPQPSoYjDJZg2pWoVz300qR/
s9H0I+RhsbIebn+QrlxzjNFWoBVgU35atTYEYwKTLQTKuUtwuLHylY35Lq218xTi
FUzh7zob1zPOEOjqtS+2q72iGcpVFqcBBXHFQQ8KI5+HbFcTvRPim8sV66qoSJtp
67WQl4b4WJLw/2ZRcG3z3Fw6x5UbsTRbiZR5yx59p6LfwhoFkdDBLRfhX4is708M
qBfp5eXRPzkrNFIpX22Tb2t0FuuFzIZMpp60YnTEpi9ZceQeu+QHCcv3IMpv/ERR
8q2C1tQEIBrLGD9qj0N/kkHHOg4SJziSqL3HhNHe1yjcNSBaYlfXF1gxjWQiaj/e
cyk1OoZMp8le5sTQguNWnKElfoirPwbp1MBnlvV0YsfP0oxRIA2yJ8KdTbxmKOOl
3Yy+zV6bMSEUHYnIAdD1Hy/dY7XS/kviW9prSMngXSTz9yrgFosZDJ6afWtiUTKP
6KupVhOySIVEcL4hnhYB0GRM62fr6LzGFuKYVpM2f3OpVqX6BjjbnHjrlLb1HoRq
Qam90dRyWT46I8NR3svMZ29pZgx912pF0UElOkYqUcUSPcWzCyaoBEARcrT+kWjS
3Z7Zc9LX0LYgoq3mDaqQN7HGoRBY6wARj2XUDxoETWzyrMdCLCFG1AitIJiGrPi0
H6/N9TTKQFxa5SRBxCk2I139ULjIhm3R+10nwz8GSN0LTLXBeYm/KZUNJL/iqE+v
Q6cdxOQWt1DdZ+HTm6tCBU1QNpKU/L1M+soI4rcYUPHFUo+/cjPXi7d2DLaiNwfG
vueN99NGOIXW+D2ukSQIEWrLImdgxuxxrStUDl4Oe5DalyThf2jDjzXjokaxQL0v
JikYVoZVXeGzDd4ZSyEbySzsN5poaNzhS2JP3dQ+s6soQfanlm2M0AAPFFMGzhab
vzR/zhdAz8hRyHjy4vOqAucoLul6vnLHxU4vqXTcBsGRLN0mALRdUiIVKf+nd0ju
Ug+IlPeZHi6r/vEUlvaSRX63BwzEknURuL+U0JBWfKN1k7OYYT6gLfdZrdxns5EM
ERZ0eEio7i68gyT75ig2FPfMKGIb4yLZRf1gIuRrtvvkJ6o06dywsp5ygRf+C2It
rYYWo1s+jCKSOBZ08QovQvoGlcVfe/zqSv50Ym2buUCC4ybtD+uP5hpAjUuO0jcy
6J+SUM2OiJ0mGA6l9IPzwSbvAbDNe6drBNiOk5Vns0XpAZKeqwYBYpK140Qp1FNP
6rRht2fx7C+Z3R20XhTufjj9fVcLGUsCDjA69NkGS3f3RQOtQjyL+lNyOQ+ltPjK
f8fjLHChepHhcg8f6vTpH/A2cJE3qf/nk3znZFY7BvlypjQgmbyMUc/RvF6QXUPq
fYsqtAPGgYZf1BWe0zwk43uy4hGnxcL9XTe2SsmsUEQppN8WAbC/Ul9Farylb41s
aBrVpjxe/0HGLs7Wz7wi5VYm6rHldK2Fgyy71z02Iilg6xxjxW0RXrDkE0BGrij1
B9g8PWDGLvZYa7xT3v/ygZ7/S/ELD+nl+saTs3Avsaz03xp+200DBljcL9rfyUYQ
NkhN+nY4BB7X3gMsxarwvBaEUI+R5C7j5CXm21PJyut+kaLt9iA54bfF8i/sOzgy
rDOfHm/qbvM0C73GcappeX4eAIZl0eG0DNEUn/gQxirFF2pTyvWOwlg2n52V/4Lm
g63aH98Z1iRmG2pbOMATiL75JBDGzT8+0imzrOKKQQGSDaVHbWjLxalpsWBAazX9
6TZYAtdI3f0ZYts97/vS0x8KafrMBv9jW8YI3mRKsLVjijUUOSvBfKhtYMXQJOdG
82+XYw7R9lV6x50FIw7rrFJM3g2wffFjnjCACJ4M/nbyANM5gv2XOpWit/qRKKvk
7o/SHzLX97Y6bpwYo+fzxXVSIrF5MrjZf+maCagqutN99ALJR1CaK05CwnfHu9r9
nYykjxsG+GK3ExguB8QC87aWywmu2OYVUZecahIqIa/o0Avrkofe5nZ6CSjH0LcB
djTsROhU2j6Av2Q5hAjL3mYOLAlzY/iiikH92FkG85yMPZ74rEqMhmByV0mm5tnj
ImTiNwp1bJ9r+jR0IIIYC+WO9p8Oyw5sHR04uvrb8nUCRI+RJQyZPP5e/DBjjVeS
AArCjYoSDOZh8ZsAA+HvU95sE6V0xbH3X5DWUYISwF/QG+vqiVqJon03Z/k3G6mt
yT+8D1kjbNmqhC+47E5nj5huSUneCcXScn0PO7X3B8qhkkHzsoUFtaU27sDy6hQ7
SsKutsvonoJ9EBdb6M4gRaq1MRM3gQNtB9qqHrVsIB20oMjdVuqa3LFM8fed4NUt
3A1jjKYszlsGYtEDsKPQ9CwJmW/MnyWXRqtVvzvT67Lr4tC4VYMNnx9sMd6y/DxD
7dokK/ZuprKBMd2O1x1YgD4IRgkKrqsj4z90eg0yBJA4L2zUCwGF8scVor4akARB
iXMJqMDeTsJhRNCqAM410pJaRTmrfQcB5DkNMud8F6bnHXykMZ6lmip9t5reWrDJ
1Ass1dRV56egFIa7/f/l9PiVQKvVIYWm2WItNyIf/qYfx32QpojFrKHudO74dK9Q
2zxL2H1STcwi3RxtDWdVaTUwAx1urbfFPHlGpZw+9SKz32x5gT9hDhlNvuSCXozy
vifPKsg2YakuKvmnTdMwtvfaUxc7nXNE96Ik9bQyhe/sNuNbBFCUQeM5g3Fo13vf
l+n6CDKi1E6dbr2aQNEUiU8FajhWz9sdbQm6quje+EeHPBlOU7IB95lnII1cJZEM
EmP1O6dRaTWW7iymPdqWHvFK3An3cZrY9zfFkhZfkQx2Fh/SojM87bASwmf9u0lB
ElajSwmhShRIRR7mX55/S95u5NCP6Tyyv1nG6gdzRye/dWKnyigSn9q3v4oK2k4m
MtbXqv34TnGDAmdbcYy3L6yHPLHOGLwIEsL1yUXhd0YbS8iLOTdRN1RhDCdjPb/T
Mqbe20/L3ZpyAkmn0OFYJ0hUE6f0H2nUOMWR+CGy8FlLw26PGck9bIOcaZyUJmt9
FPdT4gR31zAvILeCzwYT4ZTBflB9MgDiIvfGHrCVC/TpPkwXlUxsZfJmaTQS6t7u
S1KVpCl/daIGls3DLSW2M/C2ZYkkJfHgfxC3rEsPg6f/sd6NabCCPeTlB21jI5gR
i6mbYr2jywTS2elPU/Gju7Q4Wx/XYCuihjEbnmKHUTBTs4IGHrZyJdQgE8N/Mqzv
n5shgJA5pShBhLTKljNm7tZYB6kCVo2cNJKMfKwQyuCuoKwb1Seutv3EwuwooRh4
Ie+sxUv4wwIEpVp7kzwvF6zM4VZcUn1eTSg8IpkmCkJ1YjDXQ70cqZJHka9OzA1b
BLNLGoS3d8O7mRLbC6Afeoy/c5TecUxZd0YCBFomC3qPmqu3fwSDquM3oIvYlw23
FnQY1lttp1NHkA3seOjcDKoRz4eYVCny3+hWVPAzzL3tyBcw8HFY6pwkYo28kt7+
IpsFCsUeT++cbEaVQwnQNTFYdU8UqTJcn8vJC5pKMHVzKiAP9wTEBfuLS8shsIZ/
S6BkVdtch7YQ/fIYOhRf4WZ6rXGEguKUx+TILLWvrIeXFKKS8uh/3Pj5ye68fwMF
sOa5amjgKPRDRMbrYEb0nACsfWRhva5OdU9EXeZWpRmH18P21oDsHfW0N26ugoK1
ZpdY5qSwnxKa8Jla5GGM30bCIQjT2C8aWa4shi21eA96YZ/Sc9VwGSrLRkof9062
5aXp/II/O99rU8+xAtLNQJ9Jt+RsDYkLyuU2oGP9I750f2q/Zj9MuguIqEHg8HwO
DksdGqRbotMGixYJoCkkmqNlDSAfNBC2oEeu442rHUVrJxGIcd44emM9dyJXF9/D
QBfkiIHd+IKf2ku4nwu1Be0+1whkp6Ffb1BVECfw4xtgFbOg40VR3mbgHsbtUNIN
bTXAPoMtxZdJ/2eE6qduveRpneB8qinVN+KpRJ6zYHtj9V5GSMURFJXEtiIOLyAu
U62CN1381l+4rPS/1gdYd2Hf1tHaYEz05zrD7wPkjeORRNC0qHYDySc/JmhJvI8Z
AzhFHLZiG6tlZx+F9f2gTLdYX4d9FBw+Hg9oSjutu9eVyBHmeFeP5kc2jqh0ch3B
8m8/pYKwlUT4cielJru7IXAJZESvADqsLx9Ii0hexzxgUE0trXzH5jPR+aHAZHF1
FrEkv+SWPaetHItompY+KjoPFltRnvdbEu5JXwZFmzb46f0djeuGJFUsFS0DIpuI
RsOBmP3KOQThaDf0ooosViGXWyp3AsK8bJYL0NKOTyQJ7tVcBEDd7HYtOH7/O/lk
ll7/x6uBoiHR+x0la/wYSbN3clx/cpILyQ8mH240nzFwKgCALpHWxWPn79WXtcqj
0od/L1fryBxK571e5mjYFDnt3kJXjBCk5KhU0AHJ6iqu0LCiUeoj5GGJj9H2teQF
JCaYrbMr2EyHrBL8DCeGAonYWmzQzRaBxfbF2jJHkkCN6Jn8wVIBUKl7dFDMB4HU
CC1x4CNBh4ZsyUaw38tmTZbyVjnAvdxZfmE15++JemmH0LUHZdOUdBIAZYnxh+D9
RKrAMX78FbkgOwQeFAgKkP3m4f3itsHq8IJzRvjM6q5C9h4bWAEFR6wOSPnuozDy
75sWsGBn2lC8uwd4Zvr7YyKLyzZLOWRwPy9FkeAhpNKVX32/ysTD0A+xm+jLI99f
Mvs+Ss4TqJOJy9Ohg3LSU1Ea2VDOxST8phhoYfukVcuUQ3+dLAhWHS7I/vQJXM5c
SiPuBv3AVXxWGaDBqqjmC5y1nFUVaCTh3xIwVqRLnS21pnvrQg6QKXTOjTLPxgSN
yYYBx2S5jxw7OodqITj3sx+Yv7W4w41x2ShcBtIj99eS29PNSA6AFOmNksDauaod
75+t4R1ytOLcF59jUlvM5hZx7YKhKxt92jXDOuLYUv1Ryr8lE1mGamI9qhyL2tYc
6dCs4NZ0K1gkbSkzxDq5FteJyNTgx1d+7mwiGuywVxdmTB8XXgixSeFCg8cRnkHF
twm1EJMgbB4wNX3V6XKv7+kWwLl0O4NPjoxSAQiLSq3znd1F93t8NVrNfZVmD6KE
kEmZmVPdMyLXXhJjVKoDj7N8aDT6QjOylayg6vSTxggBU0MyD8AQKV4u/Ya7Nu04
dYAq7bEcwtq9w/ArQqmurW2AdnfqwhiX3bIf4kbjQkNmX1IRULCqhSHprFn59p/l
0AY1ZvnfUDkwTrntb8GOwkOIEavmztppSfxsoLokL3q8/2aljYl2WnvXbQaozWUr
zLoJIogpqK7oGcfIq2ZMItzUMAn+aQz6d10c6okbqIZkJgMH4q3uGIbeeXC7MIum
NgGmK56GRbdFA0dk42mulM5LCDlABdeC7tjrbXgQxaamV1VEGrIAfSv9ROH1ZJPr
LvFqPpTzspT9bnKXXJcnlbxqB/uMwK7jRPvoVwkEd3AEXc05m/VSfC3F8gomdpqm
jlKlWgS+0lX8ADI0euNYrcIVvTUK1NoDUlEzxPtN3I76GrOrQBveA2863MoCzinB
Z+rzXZGje6DvbLRhUKJfBdg/uS+PYPZOnY5jjBk/20LM6tNjZ1KfMdTIvFF5zt8f
y8Dm+paDMpX7Vtx0dtSKBz/23k+e7po//YRK1oYkD3PuDwV0vLGPQK0IBaV/0euf
bStit6J0plG5QKbBwwS3/Cax5prGe85siFUqrFm9KXzf1IwQSMcYGNnY3AU4K27n
miVSu11vxOUV9hN1aQ29YGtCMFT7rfcuH9tuxurDc5LFGEFQ4QrTVLniFMqdG9SG
oW1/vbIPMwg4DCtt1FAVjGMqTzLTEdY/B3fyKQMxZXgzzGNHN5y/pGv49oMbPuTW
L9o0n6tQyxj0kX4bDqmr3eAwasVnv6h5lOb/X/CrlFFRhgBqhC87J37l6WiAUdQQ
RQ60mW1XWcVJEuYyyEGL1JGRL5lqrQ2rzXghsHPHCITFfg7NmhXTr4yMgHx8Z5Qg
Y23nPnsV73Mt/4WCLa+FV9ji3M04HCMwQBdJcqylLe9SBTzEx0/OhJD9fNNkdeO4
570g3VFpWv1h5CICHI6TevtB7Ed+87fBJVW6GdjGL8RKMvu5+5A0KbI9Fl1PP5A9
aZ1qR0S2jwU5qXzPt51cZAwhStJJCNZ785soUo6OwUd4LSScZ6XHgUHPopfT6rei
W33v18EdUm0FKfbs54zAlpIi4dtYSDjLPhqlRrRSyPeqsRaqpZvV++dA2K3I+Xdm
hNMTeMAys517vd8L7MIkMNrh5keGR/7ufSr6mJAXzfW/zQjRnFg03cT/C862D9y9
R/bouJ08/ZM66PBPlR4ZUsVLQqiih+XQjqPVh9Tp5Gmq3ZGsOIxQobcP4zUjtfFm
TkfbN/ZVmF4bDSX/NaQx48RhTg6g7IOMzCrX8KrotBDOTlyY23OhkmNo22Mh1qXb
rbV2lc7qIuBU4OipZn3zKg0cLuWjDcdVNLkw5glDtRUQyvy7HPdCkxtgyNMXXlal
YbuA96xhl03MvOqv6rZSZRijF53Lj5ShdxQsMjnKEnTCOKATUdBFmRq+CmHzlaOt
ujmloVAl9MPyWFja8BqgM5FzSrS/XYh83rTCWXJ6cDRddEXWiEcpbJJEyi6c60+S
IAT4amzG+/BKgqopYF2yLEVzLxxdHZjZXIgSgRbKPUBEAswxkN2NAlIYBXACUqyL
iRQRQC9d9/E3NfD2bxxKJBKrakAekAXSDu8WdPwgjaej84wp8RnJCZ6Ak23+yBjX
6enhrjYebk4bhBO2ELZHUzbXb85NVpXPHZT+LiyXJDVlsPnsaIiT+xWVjZ5vRy0g
qgYPXKx5/V0SHAlw7VnFWshFMcwIJ5pWhadlEsfrjWP4tU2q6DiWJ6o8PswMBh/g
OpLnlYghPty+9bJF1Gl0l3wk9xu2IrRWIjLCsuFdYbniNq7a0NHCpJwefrlqQbh8
jiFdAxOhLqY9zVChT8YOwCQ5oBztA4p+C/AOUJXH0rxrg2sqURaUmP3UgJfGX5QR
tTN+T4EbNz5vFzbIS7vKZzBbiWvBwUwU5IoBOwmh3MMvWQvgBkZT6axN8RR+wTug
umnWS0/vIiS2iQ95xhzdZ80RIoxY0sM5KlYVSyLdXutUd63ocsZttNlePVRgmkoy
YYAoBUPhUUaH14SnXvXcuGa4074c8CsXS+7Yg7uf/nRn4iPzuzBOUNl7GrmrOqmQ
dplqxvLWAbajy8G2KfEFw+wpialLiVVzgNGNK/7Lse3hPFn0fWGV6fTkaDdQBk4O
sBukW61yuDZ6zerLocQLxFCp8u8acppCLdym3oObSNM7XMoYAm1NExQFpb7yfVrX
X7IHmCmOtHMapx9nSrD3Ci8vzkwKqkHBkfRsibF2JLpTzqild6arxqb41dLBaTB5
Ev0UXxCGBHCwbBncl39UKgNx5XPfJ7q/avCaYNINv2uHoWY8O0tMFUChuO9bsNq0
MLqDHHe+80/HIufqqsj6fF6HbnmNl0SnZYsmJWEo3ss63B668LcGAX+V0iBYYOvU
fX0ji/h6/XMTp+R8iR3P0HXCGP1ibYryRyM8M4bP51kd0CdynSQ5snmW/AJYLKvd
6PL5CHodlz6Rdx/ByCq92icwkg6hkALhzge45BwhXYlKuEZ4W7tt0oCFiA6uUQT5
HSo5UK8bTtXX4//sclP6gfu+kMgCqD29YgggJ7wD7WNrMF54PHgD6Q79wbFtr91u
IIlPjNk7COVIKjzTTCSrzziPv6i0AJtI5lbvqEF0ZEXBeGyMaNftkERVDo4LooWl
Sho8q6zTKTP0Bt2IuawHscqc+d9Ni6k9x8TcvgIlKb2Q4B7HaZsBCvQUIKBzohyu
v4lrqj1XpyfE8x1bOE/3OC/hcTzzRzm5sNk1h5u2chhKDiShZhHzY6Q0EhBDe2En
k6gOlAU/279+NwQqNFhiTuZQDJB4+ttXj9VEbczvhG2Py1ibII5U1jcaZOZWSfEL
mjiDE3Xuvyon1Yii81qP1+vWnOIQycQgkf82O7ls+UrgszAwQ1MxeZWabUoCd9Kb
fsbEb8p0peZezEFE2xKAt3oaHj5paGYAFP8PEjrROoHz9ncRaZhWgIVp5Oy77tpf
msMG8brEdM7M3tNqWLbqVaNrmM/kRsFFOqAfMnPiy3m1O155bDF8rqo2joBoQ6iG
KWAFFxdWLNLXLoTvLsSFPZxixkercYk6qYPAMDtUQ6qcFP0t9y912zyOIycdZWrE
KlcfdtpVQb0YdD7xfo2JlPyEIizGJ3ezHRMrp06F/2cLu8bpbYqBDzoWX8FxoSij
J7FzqplrsrxOe0/0KbGQYNDKCtY1xE/fGw0cDIZUkMI8UCW8AkbHylhK2oJu/I+b
mcPYx9ZS/oYPOOzhSvs72qKzwicV+RoB0iI542X/ndoQ6A3ZlV3rTEC5QY8lZCQw
9xd0MhlXqoKcCoMEOoqSQ4FjnfQJPAb7b5rUN4wUG5QfVkvS/X7WzNblCPVqBNTo
nij3M8sqz4mb+rjN5YN7uVSGjitSDH4C/C9TEtVq2kCmbrX1lkFFn0InX/4dfOXS
o9s4eWyy9jV9d0GHyXs+VsvQ6+zmnLbjnI+YtqYBAMcMks2tnhRA/xxhQwywepZ1
o8N8zJ+NdQhIBFIr+nIr2GebFe6mksF0kceDawW9jsHnIQkszFFYZ8iEu10ykjJl
Ji8bSdwTgOwNuKC3XZ7Q9yVRZsS5LMcgrzi4Iea6B7ceRHrFOXm8O0jC9lvS9+zY
KNq3xidvweAkAuf8ZhiC54zIIa1ERn5aWvFWtVuYyH0vw9izb0+yUXAmjircP/eO
dJQCM/UcREN4JV8842lrxZy0fHUDOQotlI0oYei7711mJTfzndNGz0BA5Ug4Mkok
jK/ErLaziXQQqtgRhIiOss7k+rjduoerWrBFSi/9ponAj2fipV3cc6hNsFDejebc
0/sTH8sQo0l/JQTfOPIoup9MbV37ncTlJ1ZBst8k29xCTad9eCK86AxBu4BdamHP
ltzKhPboHLcsmj5gbc1PXfbLiyicBKYYMP7wYb5t6xgrb/yVt/NLo3wTN4bPbXcs
sdXLKNoAng7ooUFeT63d8wnWqHBnohRqmg083vkCeEb4NRsQlenh3pbbX5lgVXaV
yyKYRjk1JN5X7aKrwYNSKnUfm1NICWry+OIzWdoKJb1EM9L/UCSjF3cN/GZMvWhl
tDj9q0ltNUoJoCPXLjswfovVKPcVBKU5UKY8GawHOY+tOw+CavzXZmIkzo/LQadE
cn4TwWT4WbmGk6bhqJZWbzUoxA0u7g3UddPx0Of9XQ/1leqNz6mcfUNrOJrUgmLf
xobdfaafFw32eN96ivr15DqCOBqKw0Wjd38VwVS6+E6OZMOp9/W87N19W7VmUnXw
/C5F3ne87YdPFu+N97MTm+dd2EcmiUM1+56hHyRT8rinwkWjHvzWhpOeskliKkh7
FknZH+OT+GvSlEX3L/ZEe0vcOFswdODExrkvx5OmOBy3njNIjW6Qk9+UNagzduAc
ZY0xnOmLzmVrx2maXqg30P5BRvPS5T4Eyad+fh+eFgNGceLDH9bO/JSP+zJdceH7
u7UsuklidKRfrqZ8EsAEIXpuuzv2bse+LlL8JA3brGNbjrbgFLrv3JmR2t4VxSvI
Y7E5FXDdMZa4hGVlLWrcUjY2aePXvcAU3OEnaqx65y20gi/TzTwYBm+XY1TeQAOd
EOICgnhRR9u/kV+mhHdiWO+WMBU89NtufKYWwhildmZE5oeMih3bAfVu5BObwHcn
IQKE4ah5YIrOrEzyiLWK0y4IYVkESC8Cl7WruyGaKLN4vywdtZk2tIaJUoghzIVr
ppGyEZqcBCd7F9RTF4QzrP/2b/+7+5OtUIoP2GK839eArZKZBRLEtymiZtqtCAB3
PkNR9j80pa/jCWekwZh1o2hOVzduyZQXx8XLhJyUVxuGxvqFtJQDayYVYD1Ll9LD
5qZ3Lhvq4TOxghBwaYOLFeqSZcs1qFlefZ0k/8vEBafso/hRDkifSpatjV8kBl0y
doQVxz9grzENaiQCO9Df42Eo+23/hJCNHkGQ8vaNQpwcBgnGPNC8Adfn9NNqH+97
J+E8G1YsKbfGYP+Gs3wH7yhRp3JcDCZClQrzY65FH4IeYGf71HYlyaEEZfndiMHV
Do7tCwvQdhULn+hzcilZ2LEqYy7/qQeEXi2wLrGiGl2QCYAIxwkb96OqHN3vwr2p
Tjayg/bs6/oNqQ8YZSSBb6VgqhjF+8vN5XDXNqMttXU5sh78hWkrizQVdsd1Uybk
HR7FJmQZNIcTYu7IcHt8YMR/Nco9beSSJUd8j/Zm0JLUkzG6bk7Xuc8dWEery8Ln
xQjC9z5cBr7Pqs4xoMISb9kdWPWHPQQBpusbGVZ1Trm4hxAc3TR/ivo7pSl1s/Ud
XjTqi36aQwU04QhQFQbaA3l55YBufLX85NlZULLbPkBzmGnktIDuYJffN17XmN7V
QzxrGSv94sBPzXbS48aBY01vf6FOXLy9soFMShy73tGhgdy13es47W5iYI5NB/qx
PTu/hXkb8S4HDykdn3kg9EZEGKGEOVboiPVhkqu3pQb7NP9fJ8jARw1uwMlMbII/
yC79qrEOts+GXpmuXGw29e6qxLoVDLXBS6aDSou2zFbeVtiFM5nJSVtJRBSft2q6
ti1W/45r5udS58oklVAAco1iTBhdh1irMJCzpq7c+F6ITfcCQfo4vVcgo/I7bRUs
E4d4im2OreolfTXvc2utJqcedPMD74B2HnMx7/jKPTci7cgwLRAbPZiEIriCtf5C
4ue/3+Z69L8TtR+2KZaCsLeGb2stZnBiVLqhhSRLtcE/4BWf1D/tUI6sbgJLogmr
7C99+/87FdszPbKGdZee1c9FAgGaduS+QsqjAzVzpfv4QBy1a6nq73l33jZ5uFQk
O9I90NxW3YH9w6Da8rsYNf+Ev6s/K/n4WPs4U/MwkeQwho+wO5BABX/S6Kqii3cI
Z5+dgQnHSkaUkl9m68ss8LVpnqquYPxFiYrcHfkNwNh4XnToviTqEkJnpcDlmCte
j6xdJKzg1taofWmV4abK28g5EOVVdkVpqeVJP6kRfRNBTBARqWSOT6ZvWmoHfeKW
+N8Htj3HyLNUUPOW3Xg6++zcIG0o+ol7h1gSQB9UVrNE7SHVVKtNDmeVbSY7KDQy
FLKQF7FvxrcuTp4RTWQz/jt899kZNza91rG4K5N4n1FhghjSuLSJt5/5Ptkn0AoD
IlHp7IRIz5YH3gl4D69Jlqt5hGsvyruGM5HmzXrepPsF0YqKo/jkgzTWFui2rQF5
iiNoGPXq/SZQ+q6cEDISwUvP0Er/72qHEA30k7GyDqutMq7qHsvhd2bUm+sMjKqs
7XaooVr1rZrzqg2SfHYs3dKs37GGuB0DIK3B1BWCYxoUKMj0aqN9BHc4t7obPLrZ
lbk44dwGh58DyujWqcGWwQf7jK2AppK83IQa6cFKaawgEsBVTEe/3FCVvsLskNDC
WiIBhP7PGETB20yFDzQsqoA2Dj2KjDLPJKrgJn9BR0Jrh4xTFcN6mTIUfXCweCqw
/8OBpBWbj0xTCK61pYrwNwiPq5+5f4FQdV5jiavHS5xHUbuobycWynk7AQxXOHUP
zADInIGxQn7x0eCrL6DpzjBG+FOdchBVTM+uov8frce72PV0EqKY7ktllvAnawsS
PgHYEJVtBZpmRMPQljw3JI/H65v0kgD8FyFleVu5dEaSfb1SUBzCimCsSrTTm97V
EdEym/DM8XJ/8s6TUSvzLAH9c0blUISJm7dUI1dmot6wzXA77B5lQj/Y4qQc85p+
qxRhaE0RlW3izRsBGVHrepMbhnQDUYoNS3Fv0c26jSyYdBpEzEUmZ2iZSVK0vziz
6g9xutPfHlpMXXnKmnE2U2uUmueRdspjeMJvetZuDF2aV28bWI3oas1GJ4yigYwD
ck0ZCPyIY2KQFcGBal0KOQB+4e1oSD933Et45q+OR+VcyWX1vb7ErTFPDyqfoNB+
+Re3hUcIVI6tBaqtzY4Fqciz71uoloOy6ROz52bcuY73RkB3nyxNJ947Wg3nFh7C
cXjvMlk+6cGDEddT4X65lW1nTUZ/Vbk+G9ANkOz8KVMOPaHy0iFoySa+Bt/k55Nj
nmaXOQZPr+LzO76Da8EUs8IJWUUldKS2WG2c13yzdsNs6pPAfRiuVSmtS8cUZW8N
92iOgo8XggHxl+SEyteNhT85FRUxyTwvbQ9nLe4TEQWoMnp1mxvfPmCHQQn0C0tF
lekqhZsn+gqFTt/4BYbhg38g7e/kSUc6rsFEs18Cmfk8cvgKGfpYnnUlLfjleFyJ
mt7nVif/s1mSMw+FxlAiKtc4JyWjRVFWUlO0OR2guwk/J4Opvdt68ahIGmtz3t6l
Xh6DEkcNvzP1xYD8lvxOtYuxrLafYCH+VFEu8lcA6FWPuoiWwUBi8da9tGod/OLI
5+RsLY3z/AJ/4y6IRC7woEcJUIoROdZpu2BmoIP2BK7f8l8I/mPGLDW4DPd1zerH
wHh/6CtPtaSHphICWaNxNahphqr8UA7QuKfQbA47gz96CVky0rxRBAghKICP0xXe
WWobzABhXFltRNROkhMWmAjowiigNmE0fsEmiyXFEuyQU2Ma+85L4hDTZPrV81jI
MwXYETtnI0AVYqwq5iZje/w95t9n3Yl5PyXLuumODc/oes4JpFE9G+trBkLLMZvR
Hh/AOw59vLCb9b2QxDDM0Y70jctU5GkPQ5Qwes+foGstiR9j+88v2MaqUhdKryUA
tlvoz8a2hVbd6RYHYug3gp6efTcymWKInRu0xmq51Sa89XxhSAXXaE8oi8UQGrcz
5wI1Ip5I01gJPcbxeirtbjp6VCSZDVaqSESFfdSaxQjQM0XIAq0Wy0rpPjg58CHQ
50KO6Kc84QtPh1/CbA7I1MBQohvDmFuozQyhthHCWMCX7NJ52Awj/p0x/1shudID
7/6Evazjzy2CQh5fjGnMbQyDCFLit0O4Fj4npS/cvYzdl+f4PL9RyB3R1M6arBef
je4ZJoUurCs1LRY0WdOH6NsthzTveupcLGKhZ+m048aY7FzCEbe3SZdyLlwp1avB
b6ogdZI6YoKOgEkkUNnCc7dU6v1Qjp52BSfBVxj05c6O6N2ndkyLCQsTCo25lqXG
8rKUCCcG3aa9e4HjfZfL8ZIJFVA7MhIYZhBdzbqyz4PPcFOTVCNw5BjMMUETxZJy
zt/ubP3B7XF8bLp0Q4+7S3IlLQyJ6acNY584oh4KSZHT78/VVVuxi7RaybWpNUfY
65hQ1c58ntz6IaMQot/8voauHx7E9KMo4OhO+lAcUoZLdQSHPFr383Fcszlid/Db
26pKJr8+fjdykoOZJJYWD1cVD7gEBso5/1cCbo7ldSFrstHiYVKmFEvrKtybMC/c
99MQEdpBQjWbHGmgAQt95U+O/G8CwKJal2i0sip0SprqPV1M5O2qFyMHjYS9onxM
AHDcQiD6j0B9qa4dzr2q3bx4yESNQ+n8jvLZUPZkTK7R2rsysxsdxdqRBv/RE0hD
NqL/PNPPCHTZyWUoJvCuq49t8rht94l49LnnD5eAewn04Dl5FYby9891uCptb75r
iwSlJ5a5jsj6vvCcbRA+OgKm/aca95Hey4VyGv3LwN1BZPNvqzDFxKmNJ6j5dL51
Wd56WfOQ67M9a3MY+1ftrWPsOIIgvxvOZS7Z8+tKd1KO+9GfXaJo86aYIdZoSDc+
yKuewzSx7AnRoJCDBqP7tZI0vs+UFKHF0jqXujCRLQThSfFEU2Ul/c6+vkiUmrgR
jm6/Da67Pl13Znacl/eUItBtgSt+X+EsndAzQOVb5SoYHHjkRHKkKs8QsJKc6pXX
CgmvSJUqmQMBk87QbxgiKhgLuYhgPE1K6zCKAXh3JnOMLhJNIqpQZLQW6RhSep8n
vhSI+uNiXC/CplQCV5A7Blg1AAzNpKv9O0+x2zn3A3czeest/qs9A9Qfs5PS0oe4
+EwNNfcbyl7fWKa95bQE31lyeQc6zxdahrgnfeKNcs+Q2om4HUWJPje2DZFlrNcv
b0TE/UtFs4abSlQj8PZpZp8tisRtW5HbNslThZczKQsUM8JoZ/IQ91SOaHd1oJBS
XlJhnOLcTV8uGdqlTxS6VKJQMt6wlX3k+qr/Y/VYzHXvjV5+N+Qlu/BY4iPFjg6+
Mw5ITM/IEiY64tLVLQW/7L+441aOhuQqqMzcWO9gCfJ8Q5vi3kb94f24TP0Ucf5e
ycOkngeJFyn42gK/gPd6L49Em9V8NrI5Ym5nPeuRBzLHhpC3woKvoEWo5PflmDEV
ssjxrW8gIylKWNBbuUHOGGaflRA4jEUgMOqDxFZIpvyPoS33wjCfJdl6a80CqPbZ
3/5FsTuzdFM9tGcq8Hv69si1uMRJwibNb8xY6ShNfF+26fwHOKlJH9bT3UHpBP7K
4afzwCPQnsGM0NA6qC20VG2fSTcTm5J0lLzEHqirwXWFz+j6uoXGeI99NyTe4z5T
6BAt8Nm7qgD9TWgsN73XeenfudChAYuSfWfVFF1CIrJW9bmp7jpZEOGl+Fs8iuoD
jquFzcJFSNXkapMPxaBWbgz93w6aPfiCVC8d694eDhivR7W1vdFEoo7XJEMyIZeA
KcoCC0lJ/G9e6DRvW0DuZeeBrbxRt6DCRiXaZGYc9pwNDrAxg0aAuxZPWMmCKqqz
gheIGQCKtRQ4v0Cxtljg2WcYrlpWzUGN7AzxelTIrG6k4REmgNoowMNNVnbgjYYa
Hkqj2l+v9RkuLxtpMH/CfSPgi9J4+YpviBy6z4ucdpT3uo7YjBN7hvsUVdbcqkxP
JkpejS7TeQ78kkNeeg4gihxm4/sZ+qDRcTc0INMReX4VIJuYmFV5xtwPV4Wfc4Po
S0EuoRasPQt2wrZRQZ8wPfFDyyuDft0aBd5tY42Xg+1F9Ckk/zFmIlcBRmgSaWSX
NKAfDLcMaggdeWUpvepBrYJsPaavjvY8vEhkm7BabtZJPyn/SxcZIh6FAGlPqqfx
0s1gdTLwTJ8VMER8cqIAs26foH1nY7+OkDJlwcTPsjqWTRT9eqYdZnVO6CO+7Eub
wyKq+xzRJ8Pkq+ECxP3wWq6n0NcKaYtilF7puSIOaoa8oUut9NayIvntGf/9oGw+
y1Qf2G3NxkLlHaoqjepzwheFT9pib9Ltle3t3V33O4E40CMP//97IzomE2ZclBtD
6DUOqu/1Pde+WB0Du7cLIBeez7trxOtehT0WqNAxBlfp7D4ePtGfnBWVwN61xE+u
u+DeM+75i/pa+Jfb0Lj2/HTqn4mnR1d5tk/qMxYGjlo3NCt+Djfs4lwU4UZyg1yo
nlMuBrqoAJp+QNuk+zWsSsHR8Tak+ViXvqC6yuq0Fi99MOLKEISSN5TL+ZPrz9b6
z43xiVOEa7YHdYrUYl/QcMNamxN4+6HKkLcwvA6Ojczav4hp7zkkofVbUkr1BTMC
7cZPjuuRZ8tzIeWdrTudlN0cyM4+fCYlC/wHL1d7wwbkputHW0H8NrgEEK0kWE3A
aFIepv+HEilqeViLh1VSGPv7MFSiTHV+1sjHnRVr8chBpbfWmjR+byeZxQTyiwp3
30t4QE5o9AipcuzBY8dfOmlOYFtsUIoo2TWXVv+omcDTPbZIc3aB2+6i3KL4nN8Y
mO47zJaSuFiWsHE5R4WlMT4Rr8A2pHxpE2CnjXHZp0JhbtTeXLQF9FZ0FgivlhiK
sfedIF2aPTsCrsjrUkC69aBN33XLa6chDpo29w/A9av/t1lynu1Sk9sej2lYmxGy
kU/I27RyB8wCE9SQAdTlG8Ha8pszTMHTFxNYqrkctgD5vP6zhHdjf+d8K+Sj9U63
XGFTVSryiZTDbYtH/lXc2aeW0scS+G5cCx0BJKDYGJ65GLKUlZjN1n7jVCaRCYe/
3XwfB2b1vS/F48EzLShi5ySqatgOmQANT011H1btwdj5kkPTMlA4LEQClt7O4dBD
jpUnv/h13rKg6oBaWdrqQLx1tP8AWS1Fa5zb6VofIw5UNOXPhOGY3a0QW+saS+W/
BFY+36TDwZPMLmc1H4IBVEFVHoX47NJoFHyEbC8XxJ5ZKCbYnO9u3yEzeRBR4izT
WKjRG1MpkEjdyZ1rPwHjLG8CwWJvkdfX5RsEetFLRexIHaLVPNmrgbMBT79HxsOG
UTBiSO+12wJrz28YGNkl8Q/e609sjvuUjq9MhCjC3YRdsRxbdURbjHNppaSWMIbg
UqdHYw1t68lLxxJzw5Tl1T6R0QZTfaj9IKDi084gCGHdBjPWNJc1TSrJsDkEuWpd
4c0rmRrcani/e8Px/wfl/Isoys//SJz0n5KizsktOWzieQD3gf7GHPbGalz3VW02
f+Vcd6c4ScGdzySvaxOWulwHJEWWnHQJPD3dvwKCxq3ZMWTVhDIO7HlvZI3Ji5rJ
Rt1PzxOXo4vyCXf/nBkqAJYWvn8CZBQXWnmrUfkiDDd+0lE/s9xAseNTKuKpUiOe
Lx0d+jP5JkcNsb1nYGYoQH9LvJrKrBACAdtU/jcd96+50qosTft1vTzG/1zNtTty
Vd7nO71pe944llvUnZadx+qTHzPmoVR6bphdQ1IHLkJK76NXBJlRXLvxuWVZZS/Q
NqkiMZ1v2v0gH7zvHiMgbxUj4emQNajtGacU998j6FJkwGZykB7ZjVovg84vtmlb
RePcRu4x1LTGbSVruZ9qYE2pw8XJ6feTD7YWMqPuGTFUVAVQm+qr+IWnHi1GN8qa
366UoM7Eiwyp6rVRpmZlCEShSUISrL53YHLnMiWw2ujj9u72DNlgMgHAuxsXlN2t
tbT1VNzBYFAtij+F+BU9/5F/nUVBFCY3Gpb2VTHE2SKzusC42moF7WGgUloJmDAS
5QHLMEwvv96CiYLCc78Rr4nWmJAt/7IUJCAc+oako0y/0ltNHH4yXExLu6c6dCj6
6KkicTqnIKcoS/Hvva/JrQf1gvTdsbif5spBPK6BeVDVrd35G+9TWgVFo4cLjDgA
KBfBG6U63HkuhOoc+EXa6FaBx6tKrl1NhyNIDpBRgG12EKFslyrFVJw/gNamAAgC
qISMH7d0E9+AHG/80gQpKvpTRIqrQO/2qwDeMjUuYynPlehUtdQU0uCfJKZhggnp
5Cp4tviCFa/nNVCsym4gmGK5WQzYP3tnpMvLGebo4v2OsQn26WnkzgfxX3A4QRgP
2klc/vshpn9YSNBXVQ+0nZAqJ1M1hPN0COWPGu8vsyih2GybsXzCYanLuOy0oUMv
/ClWSffu8/vp+eC3PU5fIw==
`pragma protect end_protected
