// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NzOwuvNCibby3FEpO6UbTcrXlfSmizhSJVdBzNwEl/ezY9BhjtHy9rqZV9BmCeuC
QiV8aBRcThd9Pk74NKh/BqfHuH9NW4imdj36CttMlhBkTqKDjBh5DIyL9QQrRm7G
Xae/F8yRC1SBv+cI/z6ZLh7UWvqDP9OFL92azfcd/1w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5648)
7G1CISnefEmRTJkvcEr7M0BTV7g9xTQyYwXjv7/ilcQmS/wEWuQhuPzYOtuizO9o
CcxKEv6EOhleucBCkAwMyIMU1CqdLXFBut4DTSnrlBLfcpLOvSMBcbq/AS+TDYMo
HaTMBqwwheRU8TzH1CD7DRt4ocU0KvkqPkWWortuuXecIaj1foa+52opSg0TPkus
3NPVF/1HCzvQiOEUbpjzP2eP2Kaxt1ryNEHf5EGTmRJxMP1ZXuGiv6JLUZ0V2/g0
2xTcy2GIhdtfnui5+oQPqSCd2UlBSTEdVldaNi95ZRi/KzwoeM/XnOyvdbWn2GcB
CRmviZv2Ec9+KjiNvSzCsUCNsjRoxlly0cJ2WBn254cc6NPIhv2DjfRnPj9HgtqK
N3/N5T8kuY9o6uuIlXphdOgSf5BcomHviy2DCLmS1VeIArOlcZDSwzNh5a8QjOKm
QfYudzv6kCViI2XGALcoYMHwDWI/rodTkxzG23ykU3TWE50BZlQ9ehXr2hXQGANS
OF/sP5DWmBO+EtPkgSCzpCfivkZaPmETyClJTy9nALCp7IP0qczSAZehLk2IuEmX
8QKKrtc/DxefzKNPq5ris7HV+rUsvYe7/mGGfy7vuKoxN8RcafzMn7aHQHCMx5qj
d4M8DWQdmhj13+uXNt8pkU8mGaXN7bv/TmmycK0hNrgFZ8DuZDYSR6QzmvSj1gfJ
UkyLdUrDsyYjLLj8NV6Boo+B0YR/kglB/OSjHA4iscESuWUSBvybxen6RHnl4m2M
E/3ilE6/XqKs/fBLleGffBZ8tb0nm3FBUwB0QUS/1h3sXPX6GC/3kXFdwX9ZydU/
yKOi9gfV4yLDhw9qQrN7HJQMT+1HEfOjiQOFVAlt5+XuNMG8cmfwutl3aKt1V3sD
SScpysKFAQQ1bGdx7sJqTTghRpYa7zZ6LH4K2Jp1hiQ4UvHLMODnnsu+vQ5QoUpN
SFN7lslibPedEXIzVW9WklPZ4rFtXC/H/gFpRPBtrxCHcjjiFoZpfCIlELoUiX27
T2dJjc+cKb3s3Ofkv1UxiyUq2gHNB/F+EdHiJogK5RPTau9BrFTBot0vJCP/iVsX
D4LPusvyeMYEMk5CXl7NAAB8zYF59Z6nga8PhZVK5afgXcqjMGvvkXaqtHNftZEY
GU47n2k7Kf+35W5POIkGxa0SRuMD/CV32XjYoCmAacQfFldKXGv37CSBKMcoSgQM
b+n1D5KXN7Kie3Y+rvJvUI7HynvfquT+P++/DLCvYUfOIdBgrp7LckKZMm7ctAO0
/2aOAEvXhfQERvnrj4is02IrbGeA0kx3aE8uW34+qwyvCya+t682Mdtph34WEHeC
6u2SDJFKLb6QjLa+kCdWwEOfKNuAkNzb8k6PGtrMHiHrzdK5CEbNZeqxBd/OXWS6
VhFbwDga8KcXfUd0BbT0uQHyIia8IrdKn3/lfupJZ71G5UVJ6BZs2vuPCB4JZt4M
p0PDRQmEbL2h1OLbkpgcWbG5+qRmkNuF8risids/V+fnwVIRiQniHxa+Bw8UzLHt
NGFQZxZOOrU1/jsqRbPQa5JIzQghPs28PDgIpdbacrCkcDVJDL8tdliAoc4MIS6r
j0eK+2j7KIpPPTmZ+G6ykzVYBankEIznRPIzaSv8P9kcpbsIDcnLpUeoTuVsr55/
pgP2l4Q5g5mHa/QexTjQmESHT8YJ9z+gk8wNOXgIkYP1u9wwn9HkvOBfBelcXufz
aOo71XsNRnCgUTonbXdU6e/bpD7/mb44poXcTJhNPfl9VWM/hsUYlzWnluAPxXB3
vDEPLviAmkfdT/dbEMpqPsHr+79RmgQ116td4ItzJ6c/W4+QBVDWCg947mk8paB5
ChFlj9EnVW2fvOKPMkcanwAq9uhsYq5krkuZCscMSSllkf596b7g1Dj7bbNrB5vr
nLCMKQBAKFlPJqaVnyQrW9OlPKd7V30qrrjBnPf86RXfqdfHnnHwn4ZZNbs+rkKl
cItNXzTCRgfApBGzHACfOlIcadccVRHuV5jwKv6qBYp6VR1wqAj2Hp0k7dY5SLSC
tfxbZEyCiL9kBvMB9gej/KHVoPqg9guUXWVOoFZXXeB9ww5BG6Zr4/kiUp3Dco1S
9sMneMXEyCipEMDvzc/0jUZW9cw5AnvzeoIO3TMIMVSdBAe/0DH2atsAmToq/tYN
xH1r8xihmydd1hJZCX+5/1eDdEsfmzQWsXRgRodteQ9Q5kEhxCyQI2Li8SO6rhHj
wm4kEKywD/mLk4xNipzpWzgd/kQHPYoVgrj4XgHlWusmpilB4MMgmHgETNbSCEtX
6PEZ/EONB+och4T2rSG+BfwU/l17Kq290BbCCLO2lfXNH6UivPiaeZvD2uK4Ba6Q
LXDdF5X73DQIQMtQ860K9LznzF1y+jGF66ee1DL3vM5MbwC8rvpN2CYFo/VSMr5H
6+4JyKQqEyqizGauajRDiHo13wL8Ecj1oX+7QAXaDk4iKOyQUJ8iILt8R0gevMZf
BVgi1M2uXig6WVFx5+mpQnGZ8P9WJ0mpVHvZXwEA6EXJ358l50cRovXk56PmK3Qi
aopXhIgGqOrROW8kM9wlfLDizoSViCPUZr+F1w/mgmLCNG72XkuEGF0+RmHmE3Ci
Y3Od6Mxq8A5+m45ujaVguOyfL0+ODDBipn52dgDrIYrjRs0ymNXPxFSkWEUm/+5m
AwzwNQfin09rMuFAFt6bRWpZnrSweU8Qferyw83BbsV9JsI/JyHuKJMQMGo6A4U5
b1t7eJIwkHKsSqgIiOXWB/rJVi7FbrjYAlAOpFKnlXMn+0fFZKySR46/yDoBg/fA
Kcx3MoR+xDSX/NAwWyCB0lki1pJpfe+snq6UYY+5BsJfNELUO/XAH0zso/pSOznw
14vHV84VCg+QnkBI0M3xLIGet3/VI5FybkJuMgWSt4pfFqm2rLJU3EBIVDK9UqpW
inmG6R4cZ8muX6tSPyakvBxgZ4cJ6I2x2QGmapCVPzOrcwp9ckyDU7T7YNtIe7Ym
XKHG++OoeJMWzhJBUDZpHk7W62l5nuC+wZW7MAUTm+eDm2ESVH80vUOuFQ3c3Y9s
k+WjmkibNguFzlZyXaWjgvOoo+g1Gzzf43t4RrtffEiyRH/ZZCpmZPUXfhKjGMkO
RF5GJ5AA/0bWrsUKwB576z/QvqQRIKPFjoQgpMlZThsZczQFvL4iazNHwQHY/g3+
TPGigLQdnD/GqOvJzfpCHETLfDH2+0o1nmQ8QpUWYbZE+r6vyAhN373j3OHfRGlL
1YdG/NBrlD+4sLTy4RJRUF7zm6J8aX1Sgi68SvsrpSwdpwiL/WHmCSU0/qbnL3Ap
cPwAANUhAOBK9fwDUKWjjzJEWSJRfZtlKWtcA17scbFTsRo/EQkT/JPKo1n0uwBP
y5DhVHyTiQIhFdlSwB/e7fqb7pwGZ/g2VZ5H3o+Uic9wyTYfAoAT8BO45fMphbPe
KawMfD9H0wHoXZw5PEcBnCqZKqeZupupNqj6etlg5cAJF+W7Gv+3htYQ1PreCImS
G5k6jH3z3H0a2FaVPmb3+FMFIaQmuugWPwk1Cd1Xf5gDaT8qN5mDg2GMwk0UDuvH
SM3caN2QX1Wnr/GT8S94iydUuGdDIJe59KXwRyfJCOxml2QPZj7t0dT0iGwjmxGW
qbML9j+yq9lFWfAsDKgFANv/lYA4DvapmDemd1teSRC2Hc8pUo0Cz1MMHFCUCKr9
pAsPhPCc9pXJVoQzAXKEg3+N6EL5zchcWM4iqts3GsDWOFgaDyD5S9Ll5VR9jmbt
VbsUseOcteVNGG7h8dC2KJaRrB+PJyagUXpY0yTTg4+7k9NvZASVTCklxoFZRMUG
c5zjGM+W90XO+GXX5mEVrFfd3dlV7INGYl7JlaThVojPOXW4XzuKXrtKD+u3/X9e
0qaZ2bm28VTqOk4Bsb2VRjxnh1k9euDZx/YawlEBQVCblMYxZ2eovQfuvASu1Tbw
2i/Ynm91hzNNNRaNBesHUqdx5r7HdjvPwsBb6y3h7ZGovyDKANrGPjwywCT1V8XV
Ev1YXUNs5NQtiSD49SqTMZvRtM8bxJLAO4+nXzfkqBW0fzVdHQ1yTy/Km/lK7XIK
HMJfXGY6AX00ph9IYhirU2F6qwEj8XnDgfunTkXYpWHOosrJw/ygo9lLbwlZcwWp
kda7n2iNciZLPbxWj/IRO6oNm3OLfbdOhVcRi4xTILPDaUmbX280rfdtH3ajcPWF
hs+HLT+yPm8BjSC+wI1C8pPRZpljXHElS6CHMA+aLj4UY/Uz4T8VB+x5dTbwMqS4
0F1GR4p2FrkUaxISRN8cXxnPw22V8D3gW9rZliMQ5YPmQUmAgy4cpEZpGy+L3M1J
4x4LTwme0mJQhtOFQ10hAIZrUgX7xGjYtASqVe5sm5Goq7OPFLaC3j3BzyZHT4k5
ivproO5WpOhxkcmwqzGizWH+ru5QTk6UXfjhopvuXzi+EkCFwqDzHnZEZtnucrv0
Ho+1SexrvMbmYsYdvhMfY8i4mLJVJ1fvZB8QvUIeqPn33TPw8IhIeXxhSyokEQQG
H1a80Poq2LLb/OzhR8H6JTG32ssFaavVBIRlyHBTmbP/45HCLM2IPLHBuPLi2wfK
vcYkIzDn73kvy29mMIvGxkVP3Ut3ixgwydmbA8BDH5j0W5y2IyAopuQI71mg914m
jeUafOdl0dlpXe89l4uWUSiWIBuftI5T3PXMI2Z2PeRGF++XqXe6HXcYwdHJLTtm
0ld6xGCgnJ4ZUyhLcqeL69HJ/UhR3HLOyxJkrLl9No1onW1sL8DihmS0nZIsOHEq
Y5xMstfMvvNFT38hL3KXqQg4TEyxRq1Wm6adQ4wPKpigwJlbcKhpAJ4GJYLbhFwt
5TPaooxcN+7Ub7ZN8ECmOWJEnAkfHTUtjla74beeuQMZUIgVCZdPqQn09tXji3R4
rZnC19b1yJg3Ot3VAY+McWhj6LnvcgrHb1/liOgZqna4tUofEEUTJWrDXYaYtDfS
ihH7xkDv7iIoLPKR/uZjJEJmbEfYPdx0ywrlA2793mXSCrBeF4Nx3i1dNFIZeEgO
0j5yr3cZ3FNqezy+3n8iTIq9dy+glKyAYsRZFLlPrpeF5wr+oGJiiiwM18FilHiX
40xPo2Q0SHaoa9DkrfvZe0NLy5ZJe0S7EgmQzDXNYm8Dyh75yesxBLrWedIQG+9s
KFCwgLEu8RPSAwN4eOMhEGvb35Nd59d1YlCleHQ8Brwc4AHSsTK/b3GmgY9nSVWd
5pzQz0Saq5RA24E8UxmCB7e20qpCxuMuRX9AdiwIt73fTF1ybqG2aUs+8dReMhLX
S7vj3n0BJ5eDpUJytjDQi+9mO1dOEiCptvKBxv9zShopEpJaYMqlf8UWN/3pcAxB
eIN5WpcUW0b4+clY4espVu4GCY4S9zwl8drU5xoAMhmCrxqvOF0cAT7Mvyubd8mj
MrqRK7J9ZadqX3ENEUJBFNFJNgGXIXbkcLPafltC3unRNujkvhUJRcEMOUN8MpQH
mPK9X6cNpd0AaM43Ez/kIG/sEhby24EIodO7SxUg2ygDNo3UlIf/w+EqRwBu60pY
MoGsE1MsUA3dcOg/Tn9YfZfb8g0wfoCViNgGzuF5N/bbJdnGgiet+7IGpfZccqLq
xi2uD6CVGjSavwkcv8TcAZJI3OTU69EUtq8VCq0BliSXmfpXptX+V+rRd2cMvvSL
MYbkwVC+0bmCKyq768vFmdyZvg2o0Iewixz9kyX3BreDXckKT+cH12IM6+vx2kgG
XgtchhExUPxtOcPyrXG72NZkCo8CcodLHrPhqSsLSdapimTLLLS5V0aH5LuXLUy9
larnzxX4rAK8+LxqZuTsSYcLgDow0ypXLiBMZ2C4GmcxgdPdoc9sviCzKgyB2UXc
/4DY0I0jvF74bVWlEhy62qhiHwnSxazLMX5KH6jv39hKiOKdbYJMSa/Gv2E3T6c5
5SzrMwGBWZyp+L50BpHPuFF+fqwTC+c+UI56CIJxB4aa/l2dZeERGEcH9BHYCBas
YS430Gd4/hoJTFgu3/skgnWqc0Z+uHqKefr3LU4CMqnlnNR+XqPmAG1MB4frxdnL
GmQEcI4con3eTssa9+0Xq2zo1ZHN2sNK54T+O2gJyzzQczcMgHncBH7sW8Kmk1gc
d4IPqmZ4XN3pj9YiPzWNx9SXWeBF/woeD16/tHCnsZ72O5XJsa64mOYxp55CDLJp
6eJOFWV/K68OtTj3okTvXb1uhjZHHkY/d7W5DHhjd9opeQxvCZs8OHLSBbZvA5xV
Js7fzGmWihTityaQsZRXQAXRjMe+FOpz4hwRn7/OhHUkreAkor2wcYGD99UElJqF
WyfKqiztpg0WeK8TIZyGBQ572ucoQmV7Vb9q0g7mXy3OSuvqpjsGVsgD8/mNcjDX
amm/5cLomLk7MLxflnd7suLSA1hbQyvEQD1gOUFWgm213JqopDGlXg6RVhjCsD5M
wtzoA/V1j6EjaTnB9Bd7HEmVj9HC2iLiwPDcztzaBj0Q9zdaOrzR1GQfCVbE/P9O
qr59ZPeDVGdOXIi6u/T9NRHF7PJjrYcVZxP6mmjblX7J45jE5l+eYKR5uZxc0vQe
s2RCGPazNjW4as0MFpuBHkrHBPvOT+fSDJZX/ARS5H0S0pvEYKPFhivRj7AkMQW5
HEKF9B6gbUNx8WHHcoWnskrgO9WRfyH2q9JrrI3PFQpeVnQ/RNTXBBHdGuempTIL
P4xSicG+ix3UAR3SjF8nnAbv04hUc+73eHHM6Vp9hAlDO2kumRYgQNkqBAwGps/x
lnDyQpS3p9hpzlKQYJDkijX6IOYuNAQzacjKEzFldkj4RpDEMNLTWCyWK15D8N7k
n70cyX4a8rX4OomUU3Dd9OGaYb6ewKGvyHNYYyqoIqqnao4o4rKd5sAYarQMzIH/
+JupQOydHJe8fjBaacfXzbKhDtrN/zPSGaXydX1AZ/fBMBjgvqDLStuNRVqTnR4v
7PMZO/7/79t7+T9icOEYzLlfIG1zxDrxKGwP60kJzf+E0p/ZDfVJyniwNTD0g3cd
9D+N8YGzghe0991sPW4oGsTEukYGHnfqjryCELhcRHP+vhMg4N0I7bdCEjnY4yrN
4vCM5lZE3nNyKvhylD3IZBmYsAQcBy3YFFKnBn44I4gJM7iF/H3PrxCuFfd2TeDZ
pmJIBU90EyUBFaPxYmt6vI+NsFWMtwT/8lNT37IiQSghI4eVyYuuqi4mzbNILlXf
kNqJw+KslpS7NK0z42JNtTPA2kVPZwj/RvbW2rnfrnTMlccRpWA+8zPMf5PZnLNy
cJkqEXdIjUDRcoqlraWxO1t3MymoVqG4A1AKt60GT0j9aUZF5WmufDvSRA0J+jII
7NDuTzP4XvbKh9Y23w1hztJnHnZ4j3pIBjzwagitUVC+DaR1tB5Md1YVNrnSxSCs
SbfHsyepYBpCCQSoiFhfyNtrp3mhwNuxGdnyCFEV1bzmVOdMsZjDNFUW+OJ4/rqA
1AL+mE04EgMVSkn8Xvnxwfk8a0oWjvEew5gUOYr13JE=
`pragma protect end_protected
