// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pu2pjQ6rNS7L3uYdtW79ogIjvcoIC5rL4HgfGMpGw+P5+xYMjn1q1+YScZ4fo7bb
jm1yiDrhl50GXFVCZVukeSrnNEWU2YUVqRULFaUj72Nj7+7NOlt+Ie8bAWssL6Cz
P/Wrq0Dyzg+klspScPWXIXbz0ynB57o9FZ2+tK7Kf6w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5504)
c9AK0AGd/n9uiEZQxOyS9MzIsiQEsXHv02Jzb8EY0cBGhfu3vcGUJYqPmYTRLO+/
GagKMeMjEJldONdflJtalByhW/Ka0CCi0odcfB2VSptTl4f54+dKsmg9zSitvmP0
jU6xfu13MMh+VHlGODcXulvI8gBOcKBJzqorNNfJUtqoQEm3qh1s8Bz4Mw8tNWfN
T3KSlMNCwzjSXoOjBk0hrgM/6IYOzY32S3Bm3UHP3ehhswQiHyJhQQhIkT2u7PXs
rnb7L9biOwNFM0opgA+aOJY5gXAa+7ght/dOVY1N4zCo7+8zrS15aGpbL8Gy+Ck5
Vqir4h7mWhZHLojLO+WMpjCuCen+Cw4ls5c5hAYX88GrD7Ubfl2LnO4WoDGNo5jz
WE6I58zctQ42hKMxVejLK3hfjuE6yfukWvLTm3z8c2vjlxYy6SDQEvlCTrSvetQj
Fq6uY6RkUDpvcN26WSLLZh2+hVqWVq/ZSrRHYcA/t7nJjica8ZG3Vw6Lz2SaKlB+
AXrTeS3XOKHOk9UkJ/lIjdPk94Xm4s3jJ2sMlBHM+8I6roLomq5xWTpTtv6THW00
m8dptfuACjKzkTdUFOxkjwzhULhSTsIcleST7wpa4DghQYiwwsGzxYaXZ8s+kDeW
PAuBBmrrv3Vx9KU8OLi0u7aTH8P8o695HFlmAR60MWJ/XbbOdKZKTXruUo4g23qn
rP9SdVtdY4AldxKbxxBrxKJ2NQEyxMMLMEDSTbQXzhvgy9GPPwkP4YAuIrsvIBvw
sNmQD18nkZnKFHcgpmry6KPHxgfwkcwEPUb2qMdH+qfEGEACNsggWCWQFiTGKJ39
vQT+LzxdK8OPZVGkY1R7gOLscyiqhZUUKdWh5uIz47A1J4V2H9PEJlx6vZdwqL5Z
io7tdyOsr3Ha8NiaAt7Aly2JtkrAbbqCH9vSciPE/iMyBlpLEiitv25FxJG53vAm
W3+qVFUywdGy9rkw6T57NUEjvU+Gr2yq+DKk0xVndaTunJgCLB28QooxNM8XXRne
vc75XzpbOuBB0Qvz3ejdi+J/u8xAOyz0JBZolQdvcZTC1tNSG0W61WnLNde5bF5m
ITpCLeCkwOXwjg59btdar/f6chY3P0pkMu+YrDLjnJZC42kA0r4nZQb2Z4j8VvMY
4oA269c8bhSgiSnuLsLIK021c1virxlkjKw1bAai4g8yqXREMDTDx54UF72diPh+
dBrS3boK7h78jVKKcYkUYWTxpKz1p0IkRJk6KmjDqZeZYzKvPjGw1KLWhovlbFK0
4rhZg3CreUf76+4HQkIM8EBCHit5lKv8BJMSVKHRfVkEhTRnQlWCAN2qJkDQX8KV
7LLdbbj6X+/zGvAmrK1ZijL8nm0gn7vUYAgYLQ3vWfMu9BsI748X0Nl+N44L5XyU
AEl4or6CoOFz6sy1Cr9JYcHleKGCKPDlNXVfAsg8S2dBMu7xCoB+FVt3O4x5P3Za
KpKX9kjJ8EQDr4xjGnncunAvNnLUlxjAn+cv+6EIxHVcf4krJ4Z51mn7xPDn2Kw6
ukkxsNgEC7suwUZ8oekK+GN8i/8nP5rpQMPWMbLSkqi8CyqTSSq6UfWfNTPlCDbi
MgKELuEi6e+Mz32K3kLU/7T/tSy1OTAp7quakMZ3JWfgD7k9nioS5OZX0SeIcnWd
SULymSbqcE8pgjTbhXLmKBrXKMa3GvfhoAD9BH4cETW/4CAMkoggrKe/2TDTckhM
RGsKQaKzWL1tcLMj8OVI7ee8QRzeHAlh9DFPzopjd0y7Wgm0iWCdCNeFRQp5RTPT
BO/qju0qxP+n796gYQUtaILkeblsZnKBH/prD2kw6FnAqztFPL1/fwTeerJ5DtDB
GpQ8w7TbmkwJXXD2hZLEfEjpsTiD6rr0icVATHVn56Sgumgq/NBoh/YpcMklJVWo
vvvFYxTdGjZtx/W+VY8kpI8q3hFs2xiP3Egy2FBBDAudcwXEPeS6Df7u2HAjU6l1
wxnrLW5MozsoqnuUHx+JIbWM64c1soeWUfj5xpUxcqxrivIOB2UdRk7NVBzHUseH
YNSNi7TkB1fNDIY43NgrP1oi19JyYIqx3bpEGbOyvZpjCofx9pV8V1Cc8bvDB2Ih
KUpS3MFpoT2roaJMkh+VNI0VyRUulLpLLxRJFDMJkudyO1Tw43akpfkqeuh5Sf5z
RzZEfZrduoZ31TI7uCP9hddv4psYGI8SfiSf2TTT3q6IrDkdwlMEs/kIQl0cfvvf
IaDyIc+kgic39utJOapNeIeb6KGPrj5lZ4/TonznqymMv6Ty7ABnygEIamAWR3bg
ckuCv/Ji86uUaY4rKQBL93MYafZK7xnfnfEXis3Hcm48hulE8MhhZfaYT2207Biq
cW0eCLbGO139JHCCf/wiUGN/ZA+eCxa9jRLj5r8LCgrHgjr43EvuXwDPlSITbB5c
tG0z07O6+pdE3lzHxsZR1W5Ess0vlYD0SPxO+xqXJX7CURpssEapxxHS7Rv5hi9g
BfPY2NO4edSaK0VYnmpFTDJzQIzMUm0ysY4Q1xShKST6mk9SaQ94hLRMXcivydDs
UATtqQMJFMXKvysRNhMr1Olv/gSxds9BTXgQPejSj+3X2aEkl5cGftedJ7wWFwz7
Uolr+RrQObH+09MJdzVaIIc5C6gPUDv0qO6AgUB58m2GDZ0Jl6GaAJrC+NXiDiN1
2aTLEyVjcVZnH3i3ZksIuFz+guVPEPSp4r32LsZor0XQEewIhXouyy1ejQUQ9N+H
h1M/S+5JxRNzY9BBeg/gnmwyZd4ja6RuuI9GmXfHXl3uCA2kYoFpXHY0q94ULd+m
lFT45/kiBUdG4nsPGXbNBxhatbaWnU9X3bleAwP+9G3V8gBT+mzRmkptmfFsIuw2
MxTXvncpQTtHso+kawcEAUDz/O2yoG5NkC6/7CQ7zM4ENEB9+W71sKPbRJ3JUF7V
qkoO/C+qLSHdsk12z/AcMzTkeOX+e4nG2kPb2QZ6e94CBhJszOXuPm9SwKEWBet6
KO2oKcFym73WQK3os7NTuQtRNq1Xd6JUbiucr+T48no1Sf2IvzcaEqBbKuka5p6W
UzW5HsoHG0apaFrNNeDMkY0O5AzslMckv5wyTvA9XUNoSgzm0SnNJD3T7v6Mqnq5
qEkLbvMwsY0odPUOyZTjSggNN1+eFertLHqNNNN36E3iVP6PVpJ05RKyRzJBAFqI
zrxGcjaNguE3vWau13Cp11YbYGJKxr3cBHGAcbokKHeMhll0gsNboyMpZeeZL42d
5edjzxS2oKUVFj8T5Hyo96vjbnSdYyop6WV0pWPgQJhEoWO7ou99cEzdrgnxHEyZ
q9YU/dL3fadWWu6AN3eDX/23HbTQF8Ge+YH3zxqATgXFe+WlO1agZ8ktb8A9uppz
vMVkJnpo+6vZjM7HFvUB92gtdZ1GfAvYr4OlX4XLVYqdG/gHynZDlE0mwxNFONUd
h9m8UmATUm9ohzROw+P848bC1alj1itjvIIl1RqjrFFAj98g/FJBR+94hBloUM7U
bEHtKifSEsVpQ+COwF1Jr82EmjAfHzK9IDzAt7leRFUbQGZCpne5gCdsSYvUTGo7
uvauSUYNigJIHSjMe06cKtfgzc9iboeAegOuAA7K0KziC+cuPENgso2xU0/GZqUm
ClQ0OtOLJBAf17sSGOGWaefMwcuuFofz55ryFFGCk5GzVL/Imd8TSIWBYCKHmpdg
Tmom0Nbes/0zHoaCoxFons1xHpQ7bhBrYRPJpJYT7wnds3dRi97ijS++14lXYWUx
u9R2AKkr0feMDXpNKW6uBKufB2cmwCuyzyrQCXXmTBCJ2Gi/yU7WtPYtkfnHW+og
hIkVQ+EsSM9lmZ76D8394tT2hiZzk5VhuH/AtB21asycZ+zPzj6Az2N3HTnDGvb0
4Wr8u3YOt+c/Z8bOh+0LDin+anXpwGbBJOF7TZWbWKWaVhcfHOOSkgyUi4BiVAQO
+3+4gphmUfqOAH1PWyjIFMgVgnekCF/mTCCq4elOzkdJEVP2274StzoynUvgW4Ir
z649sA8yu5PfoAcMQM1/RctHIUXonLUmA2p+Vb0aciNvfKALL/QbLhLsNzIlmfWF
FRtrrhrWhV+QlBhgFFnI07LGwlEzqJMfIzB6SwI4GTbodGTiu4nuhivrvPJMoz+6
7zy8dpnJDgygbtoaxVaqE+1Cps2YCezZ1GWMU+ZOU2NPjxD4Juw1TFocIKEqbDHx
Fft2CFB+LFqHZi1+OE+HZpmnliCbTKnQa+otUTeXT0jS1f9AHtV3I8pxPgRqG+kT
WRw09SkFFm2BI7XCibOioqrzGPyw4x7302xs1BVDNOSwE+zTHJkZtaWmjuX+WopD
CYJgMif9bbuVnVN8TLBz0T7pHzJPQIDjnRd+jA3hfhWy7YWPmuQjT41ymbOsJgpg
LJUdg6k15OgiROP3gN4o9+qakgMOJ6gg1VNjkkleOEnlFB3STGULc5+togzkCkL4
iaL4/9Tdd5d3WkxEdYCJpjYPk4j+We13y4f/lfswD/tL2+mW7+2C3WQfgztZL2Ec
C+GikoMcASfVdBQdHz9Zk+Ydpq0GEtDUamWUXBfkYqZ+4OvA1ymCWxu/JiW7XvZ2
v9J6HIXCVweVScSV4vcN+0QX4Af4dVhHqoSiZ7iX4LURQHl5YaxtkgeGlKlUyL8V
zJ5AxM7qdbyIAyBUHW0YXTKVgvpIzXnjnCwaHkk+DJKj21uca1zJmy4CVDUXkm1r
g0/JihwJxMPQu2DHeEAWXUL25sIJtH7Cne9KCETlVfyQYLexaMfubbX5LkEiSEO5
GsMxU3EAKhkWq2nt6lG0/kxq1Sr32HJhlkIHTh+qCkj2n77DrMZ9raqZLF22zbWt
YwqZ6LEUztbmRjKKIyLbfG/9CKpC4QPsWI2sxxJYjgXF6oIbOrLGk1c9g1VGUMSM
RqzntbsRuct16ZQr579LLg6bPbREEKHuxa4EYIDE8Gn9vAE1nLpLJMW4+ZxMz6I8
omZ5a3majuucDhymoS4yVu+0TjAHZocZtbUzwPmqA9TlATs8z/mWaXP8uZMD3NVg
I2UMDesSNWOQ6Lw1vVSo5/xSMcJuzl6Ndf9UO50PmvUFGGzfZkT2XMVnveeBB2LY
aHcjcD/EKiW/LLroydTZ5toM81Kopo/zXMP9h5NbVNMmEv3nsj2Y0aw683xVaR84
VctElysMkrqA6lVRwDeaLJ2MFfL7+wRsmTBdyEUxj5LAUIB6yEe6IqPCExomEfr7
YQQ0cmQ9pGXS1+XdePZQyhfMDEyQWEs213TMYM48h0fIwC5jjaUzIP1AV2dO2WnH
Ez6ghASMZBdCOgIHbzey6Ytp9c1T961l/ewts1CXIBzxN6vE3AAKG+KY+g50x7nr
QaGY5VGbj1mRt1NMhKt3sj3JqxkEtu1Kxacfn9WV5V7+IAlcdczRqMET4eaaFqaq
Hl/C+okr5i6jFAaJxbMJJ0ZpijQzy0rcKjJE3+Lrux/lL/P7fLGN0YvgjxTDN6CI
4E9IqatkbKE7JXQiWG8rgrVdGxSLkq0+xJfLy/Z+B/zT4oHmJqLzJPhVZCnREh37
ot8o85Ek8AKdDcRX1ewshfxojrzIjd2jJ+ctx9tc7z4TLT+zgJEXQNivRr6JLAyE
nK4y+U2OFLFUoGcMD1jNKcRTzvetTVDoies4rS5cKxeC3WADpWVde/0ok1E17GVZ
31SQuNbV5KaailjM/PPPrEh9kANzJjTpGAMRd87Im6DHQ0FSsBnOdydTphcSyjbx
fhJDzCGCAROFbho29mBKSv8F2nE/xnOPok192NM5xh0kj9zpQcACYG+tYsLl/8LN
VhNpFuvo6WNR+YVNRk/vW9JIgHKQvaJ3mPuGFia8Tcc3OlUiO4/rrH8oYhe5EUD3
OWUjPMbemGHPTs0uG8VCzEYgUIosTM8HkI7uftA7wreYvf+78ZU0OxwCXPG92r+A
RAAx0GChbfdQwEowtQ8ZaqZg1Mtrb7tWZXVsTayfaMA8QdrCNZxOD1qe4PUP0C7y
oF1oOMdS3+FqOa/oBS0lVXgbkQgQ11mTkfGFXy2j04QZq4bwgJSpW2Ap6f78U1J/
PeudEe0lypyfRv5gbu46Jry7BhcqYGxiJ6yNrX2hCXBgQ3O4r6Z6xlpicGQnV5Ie
2+htdbEIVCfWlU+j9ianzpQjwl3RYPMYK5mbYj93pVQtFqaPC7zLEL7Ptqbh3Hiz
frA3a6DCnRed0ioi46+IrF4+zOickmprTREiM3Pac8bJIniewpVxUIh0+G03UHq0
C747vi462f20pYOs035fx5aojrBD/3DbiUxSN96Mh4hwo+sIs3mvRuDZw/YYlbFL
abLKHudDE90L4qNg82MbGlhlqFmtA+hAEbRYbHcxkLkJqaUO1D1Jt7I8vUPuGkFn
TvhBuAtuWiPtdd7J+vNxVTTPF/ghNslTjumozlyjQlzd52qYfI9W8oKC4x1/YxFJ
qdEvfnnSyK6W7QmeNo+kkstdfHQlpfJXH327pH70pgSbfKdNYWUN3ef8qMQJy1jO
WwiumaiAT4XYWvZIK8XoiKMwbY+SGXw/XFGJ63yJDCT6PJm/c9nGjp4b1AIw7xoO
74zHQnxYk6wDlJfMiKTKeBUdxxr2jwM0ApLWGyQo059Mx27DMddu5XM5DMvlVVUj
AexlTH4YzXCBDeF0NRjCiBRaDTidYElLNmMNDrhgipQKcvY4JscCjhr0EgCk8Rjd
Q/AY3VAWg2vLtDnQfmVl+r4HvD542qjqshdFgxVGzi2Ir902DRAVpUNBNfh33hb0
jgTsWt6HG/iNnjGAcExs0hMynpvREoQQCWvlzQWRC6hd6KBo0BY/iTINAhSxaThH
4eG7HNGELfL47MHMVWVq7G0NMcSonDQY7/8X91RDM80dgkLRNKyAg88rOZX+uAJz
461UZ/5dN/aArA33PiFJqJwd5RaisGw1QGc8CQqQ+3+ODi9WNMO5e29+uFNLEcMy
5dugdRzEGsIWVb4DMitNIMPj30csf2PguXuRuwIQZfLeHiV6PaSGdkFxVUHWAvoM
lbMG+M495ODxgF6OyEzF2lBNmg53mWyONzEqoJhvtDVVzVR4bzaMeujB52wwATdv
Kp0z1aOmxS03bduuVqHE0HipWeDXSzkSZdcu3dqZMBfphKf4kfozpN76qJSbqGyw
CdNISdXG6Ye0qIZrY2pbWmDGIONu+/yjCsjBKXkAM9K4lI19q1YCzRiauj2RnAPM
7HlER7RpGELGhj1zpxCobNmGQViikyv47QIXIMt5CY5jAL0mkjCq4erFLYNuMm7r
QbUbFGl+jduwD3F4CUBwVC2+mkS+qZN2Jovi873JFgM=
`pragma protect end_protected
