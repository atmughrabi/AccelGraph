// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
KakQHPJxpxMA0CETfWsMCgUS7kOpj3AXD6N+X7vpQGtN/CQumCOYcUD0a3jWD1u2MWfL412pKBMt
GhyfGSGUMuitycyy0LVkLeSCcCOdllwR2ggu89lyYgBiq7eBRjtxUt+EgYhiHfO9hE4vvzx3N6EV
yXirKwOqsPc5tOj8Q6ASGLfwhH+011kTxBiN7+U0yQthRSUC3L4F3pRItaUkaZP9bG/yNFbOCbMV
hn6meG75wMN9QzVJhGaSaJIXjkqsU85WPYR5VKpRfcjPqNHDQ/gIcL7Vbdya8vnx85syYSbU/AsC
94FdwaPT7v5mYCf2PEDuUQ5wVobSXa7OqA9WHQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 46080)
cylpGfU+SgNPV8bBFondd7hvz+mnJ9EMCq0snE+leb64ga6inRKAXwxtju2qNTU1uq4xQGCTuk1B
YVgs90K4jQvSZ+Bt/G5rsuteK4qkr5wXO1R8Yu2HhSYgVkYDCzQNMvcPgFuxah4Bd4XdS7OBDFw6
96E5FSU47fngpiGJvgm3gDDJkgjq5lTbWiJLCb9Wjthy08lXqVBnNmcs0kjt6Fb5B49gLAJq+eu3
hNBhkWcKQNFEy3Px7oIAEWraUQN48H1vjnLkQrYOOsIVi4a0T9HWiw0ewmpRDiUGvPoQdkQODFUQ
oRy5lIby9BUJxZOk2i7jioRPEbrzzw96t9VzAFvtdNwNjGqzGq0z6Xko7g6ZQxV7Uhg/d6UIijsv
O8E/p4NOUDja30FYLH/SZsH3mGjLVUKpdgatYgWtNzF7iuzilK+3msu6S11Bm2YXo675a/LJm1vA
SONwCTR4FW4aVEY9SUTYohP4nSnMuPfIrAkUEDx8x04IR7N+7he5CtCpwNluaA1Ce6Xe4EyrJwmK
QgcWTPsP63ZTTXQW95HLGGnogfcRYuzLbfUVZ/E5I8Y4YY3+KZmTWHrZdlJXm9N5Hhm3l1QjOdcV
cBHHuVeYuc7f1/jxJkNZSMXG39qMlOM2ASiHk2K4x4vF1Q7KUwvGhKYmXw+IqDnZidpd7qFhjD4W
8anCh5tmH63T376zu2QRZKgHGKIYhc9uO9Vn8bm6RuQncpmTZHkklNefcyLwvDcgrZdg9/nuTJLw
Io/1rlaQFbEIDnUETgAT5vIKsktNmAfmiI1gUTeroHDlApO+s7kqlvj7ViXrBAeW9j8qZCFFBUH4
55dVajmgjXmRh0CioxezSccQqI/j6ikE9VckdqT04Yg8yi5oYd5dNwAJaapIuncGASrU5HMrRE7U
0Tuou5LSgtfeF2WA41UyElyKuaDXzEZeFkWgr+KL4qLNQxBSFlqgVwg1s3crQ85xZt12KWfBQgOv
zWsqm/9UCeifVrAG8jETgb5yNe9L1aAbr98dWp8sUnJyH6SElGLzrrNbA2CIgktn0wQq9vNKHpy0
/ZqjZF84ybJ+B3a3MDaSz1vFZ/WrcMYzHDeQn9N6y0tgnAHyXBT4n8BPGnVO0fW8b8lutuIxY6Wa
wDH5Em4DFgIsZOKb++qPCwoQhah9JZkcHUWTJSRrksuWllBvVOiwCej5HFv+IFuxiVG8XxZAlMqc
NjAsAkfzo0sczkMHof/k5COYiavexf6BxnUG/JweF/TqoY86aRPv9PCWhwq2ZLx3mI5lYSQt0k2+
EWzQSuEAudo6APCNl09n79TDti3C2pYWWQTgjwSfZAbe1mG+fNz9wbxDy5Qqb9AoCNQVKjOHYUom
/jUG51ehwvnwfB9tdUYxq2aVQRJPfXmq6ceCKem+PPKVovX3HhShkg7KIwsOHKZYqpdJnvNwW25K
jWoZKB2VmvEMhfHAdPuLXMO5+/1a6JHXwDcCKwumhvBefRTzhGr8/HscD35a0fJunjn76MKdkj1Q
BbVLRmDB2FDLrrxqcgqU2hcOTw09oDQGYuZtqJlodxrFK6nQ28KqRHdFaBtyuFg76/RNDo8euGP9
/m+1vzMMKPAU6ZJebHEy+cnM+K7n0d+TSztcvvLRWze9OOUn8/ciy1KDJ0IJYBTyb0dgM6i6km/N
QRLgrcQHjmJNc64QDnKhDLyFrfQb1+3aIlOiyfFlH/gW39NKR37SzG37d5rPd6gL3f2BbYG+ttKH
xMlmD+KVg8xj/BF0AmbmRiuj2yOYti77DiTEVHUOV0AfWbyiWRUraxSrerjRYqPica/w5q0Y3Hc9
HsFu5kZ0OTf7M6S0O7o68e524G08enwo9fl4bqzGvmM+azY3KSI/VvhpXbE+L76XaWL/9tq+6+Nm
jAMiBOCysecB4kgG5H5XVXmtfvgcDinqyEBgWuFGmOel2PDGxTiQ8KexsHVBYyl4VdcOa0z+nb5E
qHbvQfW0ov1jx1bTsjd99P9MxyUOr9zYP8gjq0QTEqDyuiRnpPmJRgQYzHqjA3tQlmGBcnOzI2jf
WUI2tYTs3Sgy6W91J3XOfpl4HL7ge3CvoR9o21A+cS6w+XoizRZdOMrpRL0SHsTr1chTw6CExebr
Kd6/A0BPZU5kF2MkUnhC4RFbpcdfujKfIn4hScKLSTJjyGamBYrJzA2+AAX85Gw5BzwsJWonygP8
2Tz7uWPpeQtXaslB9tCF5uLVgIbAarqKsNYHLB/OdJS6AWnr5ysuUL4+c9L1vObx0Kt/o+ng30Sl
FNEtvxquXaRZ7qQ1wyrAHCA1G9g5n64ws510bROsTx7bBsGuPjsc+BKKi/yFFOWqbVQATYl/yug4
DWEtPIVc/Tb46XmykXSJUaLVAjnr6Q/+FRCu0yN+3Wy5QXZ7NXWFw85pMWBYChL5+Ej5rAoMBQLh
OjtWNnOS2turAxAXupENI5sXTN84vUKTvnCdUAGL6VQuXDGjj6mgL7UZjgjgIZiXUY5H8RwlvSwK
JFR4Ru9oLV+XBoa4ln/BB7pPD3sHHeR7KsYLPP9FdNZqvMG/Qw3jwrdu+BwT6QWasSNWe+p/Wpmq
jvldG0vYCDo3ZKLpoGUtHUto50lmpEDmcwx782iIOSTOFtW/OhfFRYYyYmMM/kzZfbu91ONGEn2O
avhLLoIneSqAIXPWLlmqhpesKAgv04LLRPB5nch0l4u5QZhTs3wVLUu699HZXCjlpI69t01afeWe
4vroZvR5geul30sUq22oDbTpGt8u8DzytFQ774rVi4WEobUIqw9asnZjbR11i5Z11n03kgz0ly6Z
vBov78SssKASnw9DBV1ktHeH1DKdI7h4hRKZxjfW4pDgUYkuEShLlUHml7H+0SGzqIouTUEjL/d9
T6JeJizxiJmTPgHG+LmV/LIIwwCiY54x0Ehf/m6kJpejXiyJVkAIKr8506//NEDrtpbSFQGvPg2N
2FpPUx0H5+fp9jNpwOje2IDyXAm6L7H8axaWEXB15dPqEVwD88v4HRXY0vdiOfJMe7spPa7iwkUi
TVvd8cKmBWqpuB58AM7VZhIrrE1YwEqSCqOEphoLyqDAD7e0pen6ddVwDNQ4rE4NVfhbZMkKBfWr
QqMfpcOp2mCTECNmipJlHxBxpsSOVXvidcUhEuO7ZbG0FABdJoZTXWVt1y+Xu7DTlz7Anwm/K5SM
7UUNt5iXxkLG1z0LTQOZsUPJcGLxLJXO5OiPUIof5t6eXXh8HfG96lit5fxV30tefnzMIpw10i/c
RbJoNKJc4kY8Ioct7qByJLA5rRzcP/pPrO303vbNhKEr96cI4S3QTUKfZwj0spyavv6mGxXl2sAZ
epMALIGhnk8VMC5+cT5Hejl/NsGGMXxnC9VUMwI6iiQMb3vLqoeyoLhemyStAJ1uFJTgoP6M0WJq
SuouFzmiqPfqi75i+uKf+JUhXtZR3D/vVHca22BulaqR5x24hfpcvRNyVoOsfM/jAv44araJetRb
cL9j5WDf9RI6huNaLWlZo3bFBmvZNMaYQQQ+VK4i3DiwRs9eOBfiwA+fq5uBtQddQ3vOHPH5sz7r
XSFd4TRnFZlYV+Qxucglhq0+amnZwaCFBP2LTizxMjqFe7yICaayT3ey3hjRCbGGnjKwC3CfRTgi
aN/tu5yI8b/rvIupaCPtQB9e8zIJv+mzNK8YgqRH/gy/+TBT9135uvtsaOrOHNXtBEFk1h2Choxn
YiZO4LWSP15V/ZGkXSZNF5bSBawnjgcyfJAAx91Xfdt+oHi/4rpAeScY9tEiXUr2O5EJot6fA4My
fZRJdpXoyELLTKi2jIrCcnpnUiDqebHvvjGjaZF7sx4QMSkVMjwKDyJlESM8eqt39aWBzBwzeefA
A/GZ/j0AvUdC8ecQ7T0Ehrvgwdox6NKtDsoTbi4but+/7chXG2RNZIyKqOpZFrW5SdF/++Y3zXGa
xsK4KQPik7ojyP4Ws6MbXSAIZYCbwOmDnxr0d3IRLBRyqx5/sPVO6Z5zjh50AM2Ikx3Hg7d2zPSw
pM8VPDwZUBBH2xh0MILDm3/mOmdjuNwx0p2Ao+XxIu3g9wpoH3F2flxFVoKxL5FEBhpBm+Hi4L0U
fxnKyVNt2TjAeKb0RZXy8DpLgtvgabFf2fqNWFyx39L60W0q5wsYW7Lx7sbeQwWRDrsId+aFUb5b
pTliGnHyyIgS5OmcaCISE4KwpFcLx7+eR4+YGZ+jbHsx7goGSSr/44Fk+2q9n1qjBwJPwhDsZc9e
cYI8FzCBkc/1sS7OBpP39iIc/bBE5u3TYBQJ2ly4Yr9VdzP0wTlg0k/EuM/9fyqcf1SQYuY3hFa8
IMNjZeuYyKbMhkaE7lc4dyqvpOUYuQIwD73OBUDmZChC4VItk0ToKZa4R8jwmeGGzvSp0GERoUgC
mgNvyum8JhDMjm6vrugj7aMSesHCkTD9UbKFkm3sMi9Rah1j+4lcHI40muCGwgPl3XmuuZNNQZlF
qoBK1aGh9V51WUAiCrdsN1VBFugDzZDEjqSYZZPoPIcfaSJWpykJVAFBLoCH3VZQAKF6ksIaB+F8
Aa7R8BaQPMUGoMxWFj9DyeWKqkDd0rn8uRsJPoSI9w2KSBlpJmm57GSmHtSKurZY7qUZIdKD8mu9
AbQRW4u6B20pbkNp49As8Goj8sJLEkSYIhI6xutX132ejAtAzPWnPiH07gd9eFyZBPEemm9Keo0l
t+tK4Fj00n5Ja4u0vPNcdqNORw+spLSQAd8LjgqQYZpNhMXBGzKLM5x965tcLnJ+45zcKytJFpPj
TJ5zWwaff9Wm/EaYU88T5aJHr2b1jIeclloah3bvh2hCPBhaBBVzx4CtBmnLPBH+UkF12U+H0M0d
NXs/8SYolINNChta3XT4T25gfpMF44cAOyLThYDlgBa2vTI+R0TrMAWyGFTvTy2iPqEQ5PUmXZCU
z8Vjutqwi0bVN+eFvJ5gwGi8EAYeXxmNJsx7xiqbKv1r1wch/RNh2RqPwGCyImM6BOWy0hpcn1/h
hym027+0kFNN3K+b/AWs+oI5ldr2Ih21cL36PlOuzf5F+gOSDScvl/ZBqORKcmsSnspVnHOGEI9k
R9JM1FjC3vNApXlQVStV9eofvauRgPDWFhZFVM+AyK5j6xwgYNUlsCjk6OuGmqNADo0Yigk3eyKC
wRMCeT0pWtsm3eNDpjPEUjx5Wqt3Y1Ab7+utJbP6aByaol1KehHpI2IM4c+UteIdhPSWQGDWhSvL
P1Pmg8VCLNm8EgprUqfGbKMsX45ilr6mBHOM/IlYoBX/MBv2gPC6SAnFu6W93UFBHvVPH42J1TZx
wU2pjB22CFI7VvArJKExMRkQgR0XYzbw4ZByyxHiy/8UH3Op40xM1Fx8SAwYuaLJQVCvLvhAp7NF
3FrC9EJ5UG/1iWeo8tYRWwuJlwEsd+isEAC+RFdJVBMGt9QeQsvyd5kv9UFckp3EOJ53xidphKsI
HsciMgVy5iDa7K38R1PvZpMV5eZEaq/GXAakHr6dgG+keLs2N05sgrQIyI1f8OyN2VtGAFHxy9oy
4lVowE2guum77lREMNCgw6fTw/dl0v+i9tpQis30+lyP6McOfnYS5f5Ik5rN1+x+/PtiRRnBZYht
xKMV5tMqOGYRzbLUKFTJMQ7NmjqPVHUNo7A/Ikmaco9RiBAvShkEMWrjEenDcvAR2TX+3oluLCyW
Gz/YB2gY/NYpdVewET7a2qt19SPjt/h2VrXZYM/bA3sVC48uOewAKsUcufr9MJh+2if20Y+o4yat
9R6o/2Evc45qRNq5GtUsZfxBRGKc/Y0M8C1arN+7QNJcxwuNR36vu51aIWqkjO6PRzGwYecFnpsJ
IK+BkF5EIyM+0AvD2uTHtgWmOgMP0zi+zW74VoyLY+Oa/L08/NRbfmI0eWeJ8zpG9B5fF0FmHgsr
JZmJuJjFkjhPC0SpnS/DLhdKtK6LLRXBRI39sJkr1t4bqrUyO/HC5UoYvnnHcBHkIoe1tBXzGgvT
mo6zK8u9/kKgzwcaMvnXttQ3ZWbwQyNo7eCS3RcPRLBjPSEsYog1SsS68oK1oXg8oHomMwB3DkFn
CX51CmQGEjjVU5T7kfyZrSvXfPtgXVajZHtPEDT60M2onGEXy0Xunqwk7bFbEg5f/XsAFJzVdzfC
qwBgMBJiwP3bJ99Mkv1dSsLJJpU8wGX/QI7R2E/l6XWHXiHW1l6jndSmLTSqj1Tb+Pqa3wJbhdZw
XWGiOXeaKt0Kn1uIvulZWiXC0SEKkKybfz/HvtBltkNt2jN+KiJ5f5WwVANH6fN7xuZxxTkgADwX
xFxRmuohF8l+h/dhms61C9tL21kIhwz8yS6okSjWFLgS29z0LO0wUFzCkyvgLppTlj0GK9NPaJix
BidZZSeED2wm1w0yzlC0ZCIDtait3cglBhoIXBoH+cIZw7UapyvifY0RQ47PNmtSCbWyJ2NPGVmk
F2IUTCUZPJF8nIC67r6RTrgJ9ewRXT1UfAgfVRT9vgnJL7Akp5MXw4SmP5+FzrKy1KhTaOSM+ucl
fBLq/iCE8bLGKzaG0auSOAds41i7HZB/93cDqA82y3T/f9NJ8JfDv0ZpQiZ2ZtxvdATxJRAl/xWC
xsPNjmAojlVyW4TR5PsIFz9neDM1bjNhRWFiJ3cmyZjKVhgSHKl0FWdTiNM1ySMW8g9L3oqU0Zde
fBTlGy5lZsof9v7QUuPKtpCRlx3Fx+bJeRpXZd0Ln5wC/PsaUj5Qc3841vSGOV45Y3O2AriW6cLm
oo2tddd3zuLog2GoVQlygfnysFDKbY9EU6Yt122iyqLSRBpEhXzXuaRh9A71nCuo4aJ7TtGaamOw
Lkdq1I3G2ERr1v6Js7Q9a/PT/yAJatYhmweOvynQLYbMXJfQ+1Nk2ZOgz6mPvkoAyEYT36+DnnEs
Rxthi4Ry7ZymryG+72QM9LYH68y2IRgoYnwibxnoV6Htr6G2EyFZ++CIV3DH4A95gpk3fqcfHORK
pyIhYFe1iwbYd3Ah88Buy/u/yEc0qs+qBQBrEbCH/WVb3glkqjHpWpjH3ZTfgYujSSw5Aw4ZGBbg
STSF3MxAG8nRX62yzovcCFtnvMnkNWE2puHU9IDxBtQ7b8xdxt3xXTeDRQ601SDaVmyuOoWMWSoF
GRpC5JBy9JCUjaaGzSc7BwCwcH01T43O7hq1NrjL+o4GlBm4AOjhnHqqjv2UDerestq6AnxTQ8m1
UzG9bmHW9uHG4jDyfOrQjUrpL81FIMcrEXi3daV6Wcn/m3K0qO9GXmsrD6xOh4sfzbBPlXAvJtRK
75W4n/VGvi3YcBTsMWfjhehgxEiYZKlhjWVyOPfBLBhxAEtbgy1ciOIxsjs/HKWGe0cVgXxGsh1+
Htn9YPUhAKuaNzKAat2DH4TkjV7t3YXeSmrJ/8J7/EXhd9VdszD2xlPOdDxDwlDgzyBM3oSP+tv3
IwB/VDmyv952vMzromfopOeSet51pQs6VM+OgASivGiVESRZ2D9abC8XYmizIKNAURCL1NHiYThg
I9C8KZiD6Wfb7fQXUcFDcKRmDWA2LFeJF1aP3fgFw0XtNXnLoeHrCDT344PwdQKzhemP8Ik0DNe4
D0HNPTutT8LfJ9ILGEjaHh84iRkmOtfv+NicQ2ul2fJyH4OZbGa1aksIGIM1J5wUS6qS1x/IfaxJ
p7lGrDENvP0nKZzsJhdfc0q2In5GO9zQ5HNlkrhePclOSDuHK9eKCaKvf7z7tPqe7mqFi2WFA7hh
zTef/uh/NBvgzGDEHYEi5APM8r7AtWPj8W+YTvUGiptVVX4fF58l7+huG0nzi5QnbaQP11ahcViq
BW0FX2GkNgAVA7sGcYVRI3yEFRkW8yLYXoy0cxdTJegL6stEN0FNrrBmm34lv95BvYufHVcfoOjs
VF/ANeJ9eM5E3HbGtPWgj85k7cWoCVzazvJ+mhVJgw3Oy+gnjbBk8g/xMftu2GdqOlY0TNqRF2vZ
XjFep1vaYRE8BBxxmL9o/bCIwX9eqhReqbjxSjYGrNEihknQu1ngi9brRIoCzFb5rAuh2XOjWIC7
Cx59icE+QEL4A0vA+68kw633Lg9l5UhTxsTYrKiEv/N2xeyHrJt5zkDuCScxzM+3dVFNVkQKcHu1
Ys0LPy/EP7EqdDUBDLz+vA7U+5/iQ1PPojQJIqDdxFd9PhNj+NhHXBjwvyV+Ui83AEsUWlc+cav0
d/VvBw2ATEtKd0uM3fhm6nBv1kfNcEQiI9xy6MAVxUHQRVJbflxPz3uHDbNIyqaWc9nrOG3TZ3jx
fopy0jEKrjZN321oo++2oJ7dbmWxn/B3fd7bxZRf+K0almQE/Lgf7PR2Uces9AvmljbnsKLc1xMa
lEQ+73aXjpYyy8V3kDWIBfdNM+Cl9GOp8pSfQxI98p1d//7SrxSQKI254kXphK+rRZ6iG+OOx/Z4
VyH1VeBGpF1+N4rJZKcYOozTGQ3fOgc1/o0+moTBK9xVgqZr0/5gh7hyoTxwOTjXaajd2H/Dw/Sa
zegOHoUvH3ElDHSe2l9aRqd6w+lVPRUCu3xyug/tZdX6X9EqijRAez7ale5lLPcsMD3PSOIoTfnG
J+z4i3/YPvq4vjQ3CwJaZy8fZKW70zLvwhzxm8NJbxypzHh91cLcV0z0Uoe53zJOe06t5y78BRPb
cIf/EgHBhIITNXVrLEEy9OX5ILBEOaJLGyLGPmqFR5Q8k+YiQONeEVvs0fvu73UedJ1eRqu4eFBO
jFnMi78Jgu1HxklKWNiWBwsrIfHXvihiltEc4b60Q3rftmDoo8pUMNVhUMMXPa2IC5hF0s/rZ0ux
NRMXKGSx05C/wD0WwLZ+SCTfuOEgdio/wqDhn4Dtz3DavI7SKYVV8tYFaNzwG+cWWmUre4fxFBi7
l9WP0pPKtd5597S2Tpv/FNrHtiOHcbyQgZdVfwCrz9Fd8HX60W2edXqYizWkyuNVC5kTBHkjszaC
8yRZ3p2h3C8F3G7uZ9/UMhQ1XRxkwYCUFgnmWf5IYolRnlc89NXi2IePTv6vILvgdgqsC6RomzYi
weAy9bLQLJVnSdMf7zfNhEetb91+5Y1okmSt4dwOHWKdrhVzJnh19FXqmsAEQFz0i/h9JOSbcGWy
TrzwiPgwgfTYc7Oq2Pz1aAMTqS/D78fwu+UclH4c2B4YMBu8gM9KHKhhoJI55mZ2zTmmks7ZoIUp
ZFrEdiACRB3nl/TwFVcFkNupv6coevlUGLCiiiwRsMt1KcVh0csSZ5tywAM509CM4rjGezCvn/QY
Qxhrs4v7Gz6hTBJjHKofLVY0NWH/1HmGYXcdE/yemmhjc+rGwVzNVNg9BbS5xKNW9lMjgpeOEjYU
k1rVNsR65+FAbJ/hbopmNH7PNHmvMByXD7cfmDMff1S5d2OxKKG15FnvITq+opqNNmIs1JZLcm3M
Ah1KxPTRArG14LyaZfXnrvjfIeYDztcRcv0AlE2OaGYm1E0ZeKMxwIjQoWfVL+T98eVl9L5BVA15
TSkSSsghuBc7RqHG3st3SgKUvHt4/77ujhwuR/oAj46+LS6HXB2frSG+UupBbpoEamltfUct0qwP
XXrOejB6aHe7d2/BWpbBS4eQnY5pc02HLKK84UvCXiPHMqXjZFdy+Ebu8CBIhlnEISKVigp2ANTy
uT2Bs2Qr73PuCOafBUW4kslJc3uTtmDtEbk7bJM3wU9Zxz26nWkiutUESvrCA+QVPLCxO/ugqiDO
wB+BBi07KjvLf8zefEcJeS6tiC0mEWiRGadxcaCPdxkVMvO1d3FnBpnqn1dZ1e5oLh0zmSJrQaUf
O2lI09m1qW5XBjJq8b/SbMjbHfrAR9va5XBg2xEc7oHJTXkcAcp6iwLXH3PPt8+TNfRuU8rWVUKN
fLHJGFEbEDx3APBNxpE4V+z0FBydutLQbZDxYrF2Uivt975VC6Bp/pVfhMdUQFrKFrLGr5cArmmm
j5wk1Wob4M6ldO9CySl8NDKSN19WdTAjWlv03gmI8kJ6K6Vv2bvjENLvkH5TCECE47fMbljXIpYF
fRjJl93OVqra3IRlrABfxEAh8mTbjSNOyk3bSLQGRZ1LC98NWCu+npygw5vpVCEU0jDrFFmYjCnT
mGAP6KNdZXnGvR+Q5Oa8PgVb9Sw6ZMfNOVmCNkPqiYAd2SXR+iorVs/l57iEQuQeOULdgr+ZNaZs
fNnPdNrSsq2+WlwxkKQeNN0fE8dRrnMrQYWiARCAIg9uc/mW7ZnLmpCyqqwwCfBAaI5bP6z38e6h
9vGVpcUbTtaZAKI67drm5Jn2jLKJwkcJ+LqjCkQr+C5ku6lMHKjwX5aGehajDJt0cqkY9J8ApmL8
xftwE3hHcnL2WxnG3r66a4fnCvnQSh1I/VUK5cOKZcvAIjSPGlBL3mVQfl3Ptn3eTRjdiw2RHiFk
8tSAoL0RkyA5xecOhBi+/tjPt5qX1baGNHW5KkIFOKLJAJ7xenzYsyRrRzU23VdcTm0Q2UEz6HF/
GbI1eNOSdBlGJzcLnOvX6mwlxh5rQ6thZlNjttlp4SPhha2x6BlqSVmCbbnDS+hjnh7FeQnRmHnj
ognQf5KNVzNaUoXWk8bIzpA3xbfsY/hETSvPFMPEExMFJ/8xqjwaz/fng7LLkFl9k09KYEcDLYid
ZDwmUSoaWzPhItrgp7KOu/yTjhUXVQr/mptIQOmGp7DEvbLCUAR4bHXoMJPVpfbogN1obGQwLeE1
vISZpMgwmP5LlTC/MQiEp2D/5ppPKeH9+xrpY4hzPEBGu/8LxvkR4rpWkmQZCm9pCxsd7SGSrWVM
x4VtdhbHTGp1moQ105+GwgeTNHWrQ/ERJPOvFOo3qf8GKnQ3oendQaW0A1+IBPGv/jaZa7wAatTq
dMMYw6vpLuyq838mzXUNQFTYZud5Z4PjaGq3ZxKC6DXY9Wcx1GgnS8gpUK4yeNt5I8UeGINUUqjm
1MML8q2NUrUMVp8hmd4tfbkUldb4ZoSTFejpDnOc/mI4BPHeaskRmW7s4T5+ogkxMh3tCWqMXT4d
mZ6j9OE84oAmKueB+dOOupqkCePxHeRRih4HFNtooaBoZuvQMRyMSX604AxDECEu48dsF6blM2eq
tjEU6GDKwPJG32N8Dn3ic0O8vpNLmVXEbXueTZ4uJY9ZbTjQA/4e3TG8/6YVVm1wtiBIXvzpsA76
fSTjEW5dMNNJ3M+pEcdaeHSpuDfyACrEJHPHq0kPL1ep9GxeG8AOREOq8CAGDpJHg1z74SyBogjp
AY4Bytk28kCKhYFoeuNfYo1hU/H9Sqje3aSwbIeRgk3d+5lK3/3XlxO+/8qnjB5dpR3z8XBv8u04
tsbwOKS0Mw3jT/fQKKZHdibcp472tWnS0P87UTsa/3KrV5rlEXGiXwvsuUacCiavozERal3Cl487
Wg3JNPv1gb2uShJvsPxiizfLVTRgfMDGDUNzibDMykhChI07wp5fry0W6NWC8cFnEk/R7Q/RCInk
BFp57B42H/NZTqTZ0FCVoABZ5wEJIavH+jtTeTi9a8aTv2MVcoTRWNYVv7LKI1xGaestjVB0huZF
jMoX2hZu+3xDmedKTEjHmW5uT6xnzbh+kfS2cTcSwjzj7EUGRFKLdh1rWaSMecMksIwC4fTZXZsm
wkbx42nchziXDzh3VJkUF9PI4UjhijiZo3dBEghCjmuq9dgHR5kiYeaLuY+uIhOa3+fcZMmU4PTW
BQQEVsKleAf2IqL+b1pxlTI8Tw1AiLQpA8aVNgI2Qb+wZG3jQvqwcRUC7jl3IEA7l7eMtqFn8cHS
32KVZLcfG5KGSg1rs80EG3ScItb25Yye2hRX7FVGFVx9heQzc49a3kYIx9ZhALFHdvk3s7i71Ff9
XBT2FF3QwRLa7cTSSGKz/kH8Of5rFGeu2pbG56termrMuVX6fmMCHI4yXqTewQMsPkVHQUuB/JoS
i3ypeTSMhQMBaa0VH2mOYh4sgqD4ts22sAZtpSVnj6KmvMy5OX356i4G+P2MY0TUg2oR+hvbKHez
qAq3YUE12pIShcSAq0HbSC1apOx3xD0Q7KS6IDGrVA/88XVqpn2f6y020yprVQ0wSJLWMbY0nxgu
gzU4qGnjIGR0OQp7ZJSarjsY9dS4CiCmdwTLAScfw+ZAJ50fKgT8AYYYOq55KHYD/qBfBEdZQSGn
8nGh7t47V7kdB5xjbxfrMGwH+JD8MVLS8DBdYJk9PEODzT+DALWEPnbsLwYgJs8znSqVp7oGY72v
qs4Hi++vwcF/nq1ZI6Kiil3MEbXt8qAUzKP/cKUDknberALWXAN4eGin11o56foqEjZbo/ME/z93
Qu6qwaXHfW2hWQySFazVAjEjm86RFo/O2h//rrUh0f3x8JwMnk9sh9GEqbig0daV/q8mV3vk2A1R
Ikg9pzccmD+o2ZoAvLW8gLT3JEVyRytmrSx2y+lkvZtWnYqK8OXQ0aaPzUerWp9HI8sKb6z/PXc+
hdHgEGS8uT3pAuW3tpAPonGWaVTs9J6tvda7pjR9e/zV5ZVdC+EjLPQFO8VydYwxvh5PCqB3HD+B
/YmzBQGOLtw+GltGrZh8XGLXjepvf4Oqypl7SHPXla5EgrRa/tUU4nH6+H0ZaWe0e1ywU3BFgVf/
TKaLDfZ5vy+VT3VPzP9tIxOs1lMVLTaIA+MMQfxrnQM+eKYUT53RXCQGNdhPnrIRXEI7GckdJLLi
k+VxJJwZT2FEnVn23DxHds14bJLIsB6yjlCqRKjzQHYAOyu7Al7HHo7cUBqrRXAlviNkXFIU7Hy2
k5k1t5yqjpakV09JlvAobS4ppRJXilvNRPwWt2suF/2Fm34QYUkSUKisyQZOtHpmNVJY9XqYsYhG
pCYAK9tFI8Lv9eMw/Fq27kgrMqYyGyhvXe2VwbUBXmh/jxgcqQGu+ggmsvfVcV/qpkmO1g7kLvgQ
kRSxhRGBZ9EDX8JJ8oCuJrB/31t55PF1US7q8yHBYYQpO6aJNY9XcuO1nDXALXeTuXAGEddWAeyh
93l4P2CX0WLtP9jTGxL1GEw3P/lya1NGu5fE1zHtvn78CotHU++a4L2n7pqElpwwYxXBv2WCwAnM
KshxAGZLA+wodFnHVoUf+8EAhIjM1LBclDyyglI7JOrml7MwGCjmL2bwx7iFd6h1ll2gm5+tNi/z
4siUfrrDM3Th265VGOwKHG6hRRw18aDYIxM0ow1g8/+IiI8MuPeo+Kd+ZM4aYY9JR3DCwNr0O7tS
CWH0zm3wLu1biKejoVPWBPZXKixzB79GoiwMaXIXjhlZFDSzZ8nQPUGtMbRLubyeaVRJ+G293tvp
lHeAShCN5/dbbHdkNcupKudD0gLE/zrJ9Z8KNIRD4gP6Ro08Fjk00ACqh5i4E6DKsqRNnXPnJj9f
EaHfD2BhnTo+A89DwER0fX1gM4bFeoa0wHtsg80JiT5w10GBJ3RDULdz0mwxPCvis8IULW0J9ZiL
suKodaTcE9+jcEjzWbiXzqdDfWzD7WMwLKQc/lxs5uhh0ZOnG/xAUivugdsEYWtfgLYVFf8z1d7W
Q8nX00jt7Bq15qSGd8dV8uGhUC3XcP7I9meRw4Lpd7nnNXNj4wEC4S8iO3azPojEz2JCDCwHH1Hg
OfHE9EjbE/II3Xnr43IvLaSR/EiHrqhW7X0cmESi1jzTE8OYasupYrS8Nu1n+6ngvAUC5f0qjSp9
cXgZCB5Rw9YztmrYDFFsn5Vxju5Ljxiy/uXSgavg97sOOOir5ocXZP9IKto7i+sKDf23SXakwzxo
xvbwjymvt5BiP0ik61AFlz6FZKwa9r2Cm6bRhts/RBFbb44066K/EPGwNHjvkh52TTTwVpe5sCni
xLSXQRcBNrU6X5rNH0o2TophMhWmB/VeCbKcv7EIMRn38dx8NyKV5ooRA5xmySIH1KKWy0wpS9zj
lv6meVpV0hiaiGuIq3eXwlU5U9F/ZT164gnnuf1B5JVuYNbe8MVV/OOMOJv8USk8J+Dy8MTUs8xh
/JMAWjF5CdBy7kDz9yrdGgj0Bm1Rgx6iCgxjUje8E/UW/FWhNAQ6DTUhu5ILusYYBJu7HyKtBUu5
mAJgWY6v9ZaWU6eKaGbpk37HoDavZf3t6qmOigGxi9mKneda4kbaLP1HXNRaQu+CCd6VyVo4toGq
mw1lxhiFS9pYt8Er7zqL/ORLGzQ/DVhXZifXp4+o25uoNoyCVIkTMSBGxdWcogqLdhEiBOhJ6XEk
ADWEXA+SmC2qScRdQSzxWWcR7J2XBDf6BaxWlJT2OAttai30CkjqbUoU7O23+fOU2FGH9RIXe34M
RfqgQSTY9zXEsJcKRaLfJjvgUtoUgEVvFoya+T+aIQRbAfhkkl+6kXfTXmcdxjHo0yECWWbMwUTx
GjRfNeiJ/nj5T4IEI7bpPPzzd6QYIo/SsLCmiIp4VWAdp8HZDu/rUWqJU4r6xCct4OLjTueJu0jF
v86FiZwjijHuOVbjzMW9wkOtSy138nvrL7BB4QmmvdnN1/o2bM2VSgF7j6Xaa2YeambmV5U1tfHI
zNP5C6oE4SeQD0veg1RKWOyJR2ie31RVULXIBMnM683cJjO/FB5/NWbCY6h6xRVozZMK5Ksq3Jr8
SJU91Dlp1edXVYqen+TSzgAMDHKzIW2ipcBDtP3dswGqQVUNAduF0XbBPJaP9r0yAK9SMJ5YS/lw
gJ9Z0vUX62mNSfhkq0sqrR+2b41+8pdhaJahzZ+dUCpNQZvajU2VSefdLIZe26BlX7a1lja616ZH
//FWATRMkwwBKFCcXOa0DhOmh/KCYbQ4BqUFwf+hqocqoIQ05zvSoubj9+4UBHB4+5kx2sGmQL5h
hQQBoqBTY2DJgsul/mhWR9HbIFdbV2Qzqe0JkstrYDiGNNV9tE5cpvmZbTuwsXc/cpmcS7Z8+5WF
2rzbA6OlKULF398fE/aWAyZFHcL4bB0fbR41mTslfeyDNFDWximrwf4LHTqgo7k6iewfFwWcbijS
r9FFb5yL9gxEoMWcKDuxBeidl5KYXL3WvxaL1SvTljv+3BPtN7LnT9s4jBb1gKn2yPJy7er7/TiE
bmxtYH+27MAUCwam+9iTFoFGS6qLzO0AWGrPnmhoDkGwiVKIRF6xKy4ly/ftJMltxYuecfIsU1jQ
oB0o50P5WE36dlGi6Ir8GCiK3KbMK7wS+OxaNSIJvWnu9RLdZZRF76uZ+gSWRlvN/Ek+2nR85Qfg
Dt/gYeAfpZGgYXMKiSDy9ySj7SSahOOUG/kyG5gxbC+a/kDldL4WpRfAIgMxtWYZL40tF4y8Zy42
w00CvIQIYCvIdWKKlqsWeSr620be0rmdZJxUYCLizZhUP1IwEaMLOv+yjKnjqLr/NnvKKwybNdwm
5jvZ8415VGxS29jaRH/mGxEgUvFzHFiF5P/5UFvhZtr9aUC2/g50oJpqY7t5LNmwM7PQrSP1/kFq
VAjhg9WoyEI+26F4SsGcz3h5/CHAV1QyYbniqSvc/GJCLM67PEiJv0k3Cd/i9UQjJQBmnxUEFK07
FizH5ekGkstQ+snIAfPA8xqk08u2OvKLljHlV8Xok9ocbJx1h9OAppZgJdIMUO1tpjfCGuee3LZ+
9MvnzsPj1UyJ7ZP52BS9oYROgye+/piIxRQaKHgu/5gzl9cW5x5T7PI1WNnSL78JMEOFxRBOYHAY
i+LXVfbzPHG2qA9K1sxR2nTPW9CKMNCmT71yfPmkdhDh63Aev7vV5cDXoPVcQEt54NjIMB06Av8f
d8gHzqCO2/Q9XGkcjkpMcst85aQhld3W9DdAiLPGYqoa8DwLuR6/gApZmEFkknuKF5Zv/4OvEPzT
8QI9rWtNYb15/hEnRQFGRAItWAxu+SgFMbC+d4ncNkiWNOzeflokK3uJDJEhFe2rsY6OfrIbZVT/
+81yTSuJwN7j+PruFSfu4HaAt9Lq+rewZ47l0byytJ+fwVY834ssCdky/WIo2nJmnSAxPVqSBPXR
/ceseEjT2rzhqs2IZeHZuUwZYwOhWfnDfhOYoeai1f4D9tGywsYnD3Rsym/Z1QGT7U8gRZkr2yq4
7dc55KZ3GxjvfnbSTp/bMedkoqkqVy6Iy2sZVhBp6mnthx5mVfs8UOfxzQJNf5oGR+R8VTpCKbJs
U9fB5g9nNWynPxrUksjuMowoH2t05dDiLwV/iRgWddXPWhcecZIIi8lMYd6WMQIMjSHr5cuWrNeh
W7aqaBW5t2HAm3h1W2ArNUNRls7AYkzVA28yVUyT2oEDpvU4wNHOGcWymDDKYFEidTita31R5CSp
lqY9xGV3kNhlKwzC3UUsuxE2WMc3OlfsDJsxFFZY4KC1bndyJEsi3tlLbFgMbhJNxXisGoX8LMNp
Y/zVRlxa8woJ7wXJjV9PNeNe8GXlyJFrNqajZz2Va4HlRPWLzzKzGFCwICATg5nXDxkvOD7c/nYT
AyPwr7M+EfvedvOlauCLdiQQiYINJtKVodRCuTLa3P0R9b4gMtduw0sjZmd6OSKPUhBX5TxYaiXx
FNgRiafDC2w41ukbEix9Rui4EBLp0Xn+biR2a5s1PcTbKy0OslhFcDkQbTzJymQPveq702+0NDOM
M9I9nFjc9kjTVeCvigoxlcEg9tOXDmp9r/EGAjx9nYPmAoC7KBUyu7G1qW8m/kxAnWwPQjPc2i9c
gFRHRsM+oKerEY4yFjMAZPeHDmmykbizkbdMv0ZLiDxGUMi3Prmu7ejqKCR2PoTTrLlcDSdZ0ufd
UwsSKf5snJbHTizYOhzFc8icq4u4tpFQx2HJ+EQdv+Spt4Q5s4JTaANi2kcu/7b/kF7cZoq2RS65
UZnhi4gCwIn/EDa9s3fJK+UhI7fQaRJ9gvCk81tIEUMVnuqo2dZP3zAQmRCe5gsOLMrAqFqgRgrl
Ui5DQB9QukAQ2GnEuItSdiARTLR+CPVJtDdR+k+83MriZ7WG08x82RLm6DDhSjPcVFNX2rMr+CrE
VMA41+rnp944M2QWd61otgWXJA58mtwmdf/nEjCUIxheM8Zw8IJQY1eLeOVZOBEJEu0U7tVEgtoX
JpHxvC/H6x+crke1ZopAO11yLP+AGh0SHKwU0pWhcLLDC4exocpj7Nh/Jw1xfq/WtJqgx+reDuj2
jlANvb7E9P1HTJ9ZmdjhF8+uHk0pTl1xYRMfTUeeIWLe2YWyPm6ifJR2puleteSdgK3GW/iwwpsR
+6mlSR32+YhvgQNJ8q15oxrfIRbWDuJtdxQpNkfVqfJOxxfMZsHZUox17B93CknXBpCLizGoR8hH
7Xs6D/1B6EoTGgPBdi7g+XjP1iR4A369CWa2c8AU/lCFhk4Lxs/njmNucUfXdA81Hs5eaLC1vDXl
TOVT4fPrjjVkhuc6BtUgmIpDupeKbIbtM+jyNfMPwFNcujwgtnIpZH+UMg7h2al5BOMVA8UP4fUD
BCI+ZoAIlnAtl83u9RhTpxFb9y6oIEMrO1Q2WshLmyqhI4ZiGdEjl+7NkTbFD/wJi7E+lq8eK4RR
2yxr3opvS3I2pb/SKzDOj++srNdp0hITLmbyyXg/dmSXGG92ahQfrKbf1/bl4Yj69/BAWm/UFA6g
UYDberuGenuQeLTF90XfxUhwgKYr6arM9aDEHnFY3pWKDkgnQlJMWSFyGkMMwVVinBVyGKgwPTtu
XUT/paLhCKYwsKsZ3cv4ztTKcCPdRrKjm7Wkg0ejXdHQyE+FTOKHaMMXpHl1U6e2CTHcQ+RbbfZz
QAywYwqgkVfsOgMfP/KOr8Tedbi5gblauVk0oGVgxdQv2Ivg/c8LJqUWcpGyloeYXXygRtJEgnZe
3V45Vr76Gab2GSDouWJMFseMbtyvkaILampkSJNr6UOKrc7gZAWlRjF44rOizDGOGXLwt6tbSFwx
YPMbD/hH6IqpNaYS/B7V/5NGoIHwGddUAWyQE04L7KuKA7L0VMT/Wo1KHp8Yjb4+UPvk3k9vMayo
fP5XwI0iD4obtPxgqL1VvYMG93j11/a/5f1olzS239W1kMZeTtclXZHIzlL51Vk9kc/y1OuADTgW
McHfd7zUH8yl8OPf9WwajiUjQg0JnMnkj/3qHj4GnfaEtam24REtObONiiLfnDkwdY8pHUkSHDO8
VhgXmbvXAyJdQtNC1g5V2cAhSY8qXOhqHsU8wBYW73iKAg56rGnAy39zg69q6mSy7bCEnMM22wzA
3oUy35p+lOQwCr/hMTR49mboVPApBoW8afOoM11Kpxzx2eUU9pjAcLP+bgGECJr1selCuJjk2Vy8
s1ppvQVxgPS8+5UHEd+TIHJFrHzE5dMKUW8YW2iOoJG5Kje79PZlqV0lWoI8Rzuie0/5HH7WBwoe
OEN+T60mn+D5nfHRRoES8qBcRGoWFECSFNuFNq/kMqQ8qkVKvF4QPqjn843iz9OgcEU1Cos0Ba8o
/8GvYEaAXCY+YnL28EM8O13kahv1owNzcxo1uvSAX5Wz8AyybJXmgWiyv0eHFV/8s9t9a1Emmllc
fSTIFCCtJks/fnbF9xpyT9Y64H9uunN0dOQqvQN8Chfcw8ZXLio6eouVBISWdokK7a3MeGTiyDlu
sEtgKtx7qB0kKDaO2CRlwQrZ95vto64eOruht4WVGYHJ8A4BmZP9NnYT/FPYv/3jqPmcXP/i564P
xPmsDigvpIo/OIKrCEi48bdezs+wdDE4hMJpDeXHZr7vm5mOMB7BR5v2eoP3FlJ+HNjVAO3Kq88x
UcGymhKg7d0pPBvmuZhGMnUxEbGiVkKBBT7dXBh0VhNAZdr9sLKWHWtFMlGlQyC3E0Hqxi9AJJkM
Yw9Jcj+mEurbuuu2MIiIZOFBxUW8XyMicZz6V6d+yMpXewsza3nengsCMpBYG9JSPC9gOi0nFPy2
kCcee+baemS29Qp7912JWC7zL2F2kh6uEG9DflH3b7QNl+lgLUQ/PelClXPDJeSokduoQuqcIAbe
AX7dRI/AH/S6SvRUhWDhvYL2lLkm+nWZ1npl3rVfPRFlJsr8aIo0fiS0Rt3UFasXw2uceAoDQl7n
cpAD0uiGgVwOqYW6fE0N4WLnIq3sxPxbu3Q39XZWYszzHRkpw4b22mbdprGBk2awQwNCnHGROVhW
T1tX7vMBPF1muUp8r4xEV4U7CesE326j9FJGcK/aUEhymbKmhETygUmnYUVMOwawl/nGomCQZQqV
D0z+JFmta4JW5ub/YBpUDM90hGmrevlt2mFv/Z8QLN6ND3CCuUmdxSEwjKRya+m+e7DK5SE585hc
DYGP3NWJOvw3Xg725nEjcs93/GH3ksM/RoC+QSW/zpRogfShQU88HVmGGPh0YLdwUci7KEvfQE4G
8qWeCzYLyMwkyaoxd8pelwwE55xXqHG6DXdUbNPzmKzcnbCyChhtATOR355iqcNtEsc7wBkXQ17p
09AXhGePsfAIbso8yq17iEr2EDXLEnvCVCEAFWTS8ThGeOCIc7cqRoL+YF95zwm42cBETeRxnL1N
5emKPew2gEgceMa79+F/IQ+nTvX5R4CBBqu+MnibJqNSbMfz96xG+m2UtywJkeUAPsdAAxxs0Aa4
kIX4Wge1zEgJvhR4BK9OVKScoUHd1Wk29KWJi0gJNIKieVZfeui3o9hjl6eZwFlC165E+GK1/svY
fkpLk7vNZ15T+IpVvRxj1AzkPFc3zuYa0aqbGY77VNDg1txCeI1pCxXv9sbLD5kAt/NU3JY3sj2o
rt+D1WUebFN4wnyJcsAEchqqM4gtIDTKKXmPFg8TRFTUv55NxuqAmLa+TnosuW1JW9Nz69w5C1Q7
WXyb0aEnfrfofKZIxmKCgJdLxgbWg6hCNZeFa6iIabgScf73JpDmt1YfSICPqg3eGhljoNgqZAR2
5hBsAB0josCp8coKd2GE5GBXD2bdmz2mK940NSMhGPZ48dI0aA1p9NfObzfDXuT10r68B7v1xuci
pweinvnAerMhdH7bxBDg85TyYk2Jm05S8W1r+5Bwed9vgIjMOgqsr5vx7b6ZAteMu+4TL3H0T9y7
sRFvInmRZusZd9yySYI3Vi1Ygq6RDyMwabIKcwZyMPmm1y/CYhna1JIttfZdvMgMpYvqOkXQ0no+
sSLW/U2YMh6XMFymL/AekKwnlUbLhFOkz13tOYWckB6JsaliYxJz6f9gfxB5cuJSvWzhBiqo6cSm
lLAWfqcQbCx8iGrSEU5bR3yShw0zaBRs332YE4WQkQw3KilwpGdvwTH0dgw2WZBEAdBtAuMZ3pno
NJ23lN2ghBzC42oRAAjHr+Xcvnl473pFyH6WNHmufuG6jS34AHeaxIhXzHaFc7JE6STr0R4EDu2Y
89vJmg1gww92Hy8Zht1YvgP2+d/DYD+AogoIhgqXCfAFApRQ+UWMiae+s68WulWkrIFGHz0Mf9rC
Gl4ob50SHUx9RtVC40923ajdbqkfnMw5KbGC800/8qDG2meu4PM49LP2KT5CxMEsodTGV0humth1
NbggVZE6P2vsSP5BHM3zJ/vzuyc7W36Y05Y2wmHZev3OxHXh7eGGQmuvDF966kby+U8tehm73Ukv
sethWdC4h1RizmhlWjfa9BN5nLqjoTehNNdW+NrTB9kYf2c+GnuTEEVZtqXE17Cg2LgTi8alvama
hHBB18m0peAc2P3E+c2Ear6pa+tfy6c/IjyGBdAok8suFbG2MyXuPAtVKbyBR76LA3B5tJb8nGIU
F0tt5rcU4Q0aeu1/uEL4ezKDI7jeoT5Qa+BrFwPBO1zhVDB0uXsU+8X6mS9BL7YW2LXzOJqCtuk/
T1Tixzvglzu6HoOQFPg8RS6BJkpRsw43VObtXEDZNXM0dOmp92my+UvXLur4gamXvW1dLWYp12d1
W/2pmebmDDCmztge2oe7zoNt9vmJ4Hl8Sk3k3DVWxiivLjltLKCVK9XNq7NABCsHNtOdgkYNYwae
cuLkXpWs7h8nJbP3EvyeDhRnpAg45GG+K0i4gFuDWIsp3Z45xQ1UYYAlk57429PQJYz/QozkV6P3
HrpDWdjttP+DMkxcnQMFFtAd9ofT36a5fMCPElkPV+Cmnodoq0hnW0Zj0eETzlGnONOCBa5XNGNT
L91HKlfA6c7Ron/JAhKb39mw7a+Z6jG7DO0URkyCmKPifVCse9ZkFmd2S93layymF1EqT5VndC1d
QUKMR4N2NWN5w3V9y7sY9t4gqXX3U/YtHv9SmGMAR23FsU9GkTUuiLg2gGk5nmNEeoqbMGPtofHE
5/f0DjHwUlYYxvtOlQZQgPWVmkEx5wuZtyNFxBGo9kPmJOJHxMbJej7wRHPWtHWUKPiQbp0izJux
r7UIis6sr+NTZSaw5Ue1kZCCAjfwKlCO09xY6oWsKobJMD21e4uiE39BMfz+0TsMRQR5WBQpXo0G
PYmcmm3MxppfeCpUEffltGUm2Gk0SsG4IZmuifVAZHfjzG9Zt3q4BEp4uijO9pCe+0bdI0XJw1gk
gEjre6LhCEMKTqRm0jizTHV5u6THJVuYoGPp1bw+SOV9k0hkV2B76l/ybLGucnkfZi+pQKYeJR/r
C/UpF5iYEpC1FgnWA45f2ZZbiC7jP3t0T4rTtJFBXSqaat68wM0SsiPoSXnggu3rgxl1lxEVWPES
UhkhzSrX9Kgt/KjFz3t8Nsqn3E5cN9l3nG6RPTYH+2tsTAi+Xo40LWKH+D+Eh+5cHogE6bgGSIDR
JZ6WAX0w2tAq7ZsCwiWt0an69Eetl1chUUF06/3E9/F+lIq3gf9/CaSsqDUYX1aSnhb6j5LDPzhN
ngxccGCRdHYHhs73mefbiZsnOInTvySn4S52hQCZjONbxK8vSx6nW3LMmfd9C/8jWFNC2Zr/tRGL
Z9GhnRidwQ5z9xG9fbXvv4b3YcB3FPBbjZokSnWwnU24/hk0xVB+qLyvIK7NnVHbnHgbJbu+IJqd
o6ECkhqcqT98pvgK/XWS0eme/seKqdN7IvrCCfbHdOzdoqKv1GueFLNlbwLyFXN0QpyHvIJZ1mrt
eoLYLJYnyG0dlyKrIuaTujY+uG5Pm+SpCuBHF20nMhujCLL6dt1493UpAxJ6ze+pugb3zJpPq7Ph
p5dZRctO+UMxYC6Sz962WjMc108TDPe5uiuRdMQl/GOvUV5cuQOmKiNdvlh31l30t+a7bbaN63N+
HScoxzLKAbOSFRS6ENackYQd/IPnOb73tfc7Gfcai4R+bpEo0gUn53KZwwQRRtW3NqJrz3YAdPHc
75vHraBXz2xKgdGZvLgeeeA1E7UOnTnsJV5NX11Kt7EoQlVsHiiBSKlB/+aChkuGGum9AUEGyV6n
r8rZFSANUBT4Bu3TLDcY77PWCr5smy4i02cqTucdabnV/sJQaqGJDCSdRIQYNifZ5LcQS+y1KHLg
KS4EIb51iujLLt6I3Kswbfd735hcrbXPSxwTf/sD0B/Xxx8s4o7n/t2Um35rhoI9mBPQfPt3UBW7
qQ2CtzvohaNdHsSZKk4JjQGJc7L+HxG//1d5lC05sfKGNxA+54O61TmV5cbrgI18+7Hp5y3PE7cl
Ld62f4Djg3KkH4SogF9bEkZTQY9/1SHEl3I1MptFB/PAz+1IdOgOH5Dhm7YenC5lK6bkrppEiHMP
dxKImZiKc2UU/nO84GrrGd85/6+jNz/Qh6o33a9NDUIovD7UWJX82GjlTxHyehTsXH81Eq468zHv
mlKNJ0GhkLITzgPoDy+nB5xM1lJ85eGrlfHiAc6lUnAaGJ0uzAEiU72borEklWFwH92v1C8mz4nh
oZP1R4yiJdfoWPxL+FIWINtCK2zmLMn/+KNKgljEw2lcM/5u64Y6Zko7c5XamnRsjAp4FpBL2QX8
xJgo1gre2Vns1qeo+bELdhLXpejXbPsJowcdcy1Z9b3NrvZGBTSzM+9m+sWxrkmHpwGfYMW13SpW
JLKTwSh+dbMdkfyqMY+ENaYuK1hdvsuXwaEFRE1rkyJBWUKPmyw7DJj8EpY7sWOHDiAOufFVSWRq
ToGdeNNU6HI12uD33htidLsqzcenFwGFNhxpAkDlaVm2rNiJM7x1uCOlan+7hQ2Sh0g3SO3AiqyD
XunejfS5CS+FHtUHlkskDlCQc4Y3q8HTEhJlT/MixCLs7/9oNRwMQnTSkzkBhK1XrHXhjWcOblYd
qTZwhTsk9dUJhYIua+L65WgIneTGmLkTqHegEsRx9UCEK2POWwVu9i5RmiHq3ljj1TwOwToyE89X
DZJpNJuTTzdujIlLSowEvZblVIDeLUqWO/7DZTQrny8ZnR9mB3Fuj0DHVInpByywC+QHyPB3n9DG
k6dmTZI449GxwIoPtVoXLWIONX1550iE2EGqCQlRnc0m3OaH+r2uuxfVipSYNvXaGqoL37QRSA2K
0sBrAYCSPmShmTbo3GomYoTF/ba+ODeLP+mx9PdSDgJk/vkZCC99Fa5maqoIWTq81DryMStxDQTB
R+5d/EESc27VRGvH1a3U0kiHRW/0eTihY9SnksF0ZkYjeEf2wEWjatOTA7EEZtiOe8kj76F/EoGa
TOQaefzhWuIajn+cDjwLPp0JC5Fv35OcKtAtL8VDgnrp14NGrvhSVTRsGXTNUY4dcm+fiIstAzZA
RUV6ye7O7++n40u/KQxAuUhvGm/m/F1z6n4uNo9CpFH+eERdxapQnco9YyRK0OYusgZfR91Si8pZ
RWROP/OjA+afXb1ZMYmk7wi1ckbZk13w7I1Epr9HyiXNGe9L+56U7BvyntO3+Nu0M91ieeTiV4NR
gVRGgpR828kfpG1c5B7UjuAGCb9Wk3+Bm1U80w02qGWEOhpYItMV6vu75QNsKZkKGdnXu69leMRl
2ya5PGoMIu3TYNc4hLBgO+q7nhzHHaoNe3EK8KyAKpUoAN/5m8/mJjFP1u9/erLCi/LKAF9q8DYp
6k/coJHeWpTMZm9VIcE41sXMmiTwj6CkFIc7ZmfCdbQ+CtXr3IAqegejrD+0bhn/Obznoh2Mb/B6
KffBeZdKOd/blJoK+PvTu6JIlr5rPNoxqRVu1IYxbv3Z0qZG7II/L8c51uX/JNhVn/CF+mOex5hn
rtid800Xv5i1vcb5mJ+FCEbYWDJirh+aOALiP5J/qY49zhMpYCV+9l/pAtpusXNYFGRD4c9c5AOO
k5G4BUceb/0+oS0WzgwH9VGbg5KRCdR0rrVrJJrQ6Tgdl2hgfft1WdUI7UJVmIHHkeNiIp3+4Q/L
IcWYErPiJFtXXLNVpaIABmRV03PUntJGed6wu642bbfaNYqlUVPdrHiAs7+j4wkb8PyIPpIXeF7C
wAXBCpEzZlGtTDrSl7xhQjR+6DgnFrhGNtv97XQ4gUT/ktUhcYid26tIBqLC/ULEMVr1YT0QG/Ep
qO3Ko8sAIwmmedPLSi25617ZdexlaNd8IUUCCmFvPxOBlEb2/XsDmU9hqpcXsKpreXAxmJ+4Jtw4
woNuqGpgN6aA8pUjB9bzF49Tj3/oywoRc3K9ygoupdMAVgbIRm0z23qKBy0AMcWMkhLS0owVEfFS
qLpSY0/QKSigCpbHlIkZxOhJZNpKJwF3jSDx5VhhfFpqn7+M+G3VabLfpoNd0EH0+85Q5HQ1FgtG
pVv6khP3I3ISABQjAn9td8hqMR8kFo2C7iRcmTtCYIYhz72Vd3vN9xktK+nJter5LxgHqtlb/c7j
NW/J4VSbje11ZxCBuP2QdP5mkoiUJFp7yg/fQ+o+lbAkCzTPwwV+Vg+2sTdyNali0tB3l5Fg27r/
bbJTwQ4REL3U6jQMABkGIztf9OL7pXzph+Ic24kHrTW7IV6wn0t4gLyjeEmvil3hQLWNoJdyBm6l
mn7kUPCDi3E/cNc0U6Ous6502sqalxKwbbmrLDtIgex2JkQ69KIC+XKhueP43CM13tkg15ZbKvWI
W5vbCX1oFliagLqT8wn1+PoAPKsgFco6ieubixW58puh1H4C5O9x7vhAY5lsJHlhd0AGHB1r6Q64
oavR8n89TXEZdUL6ow7jitBlII3L+OTrYXv/jvfEVzD2xiFB9kToEMFQwOGO8XcSZUL+paUiKmnR
TWCAHDcIB+lcnykYo5EfeTafVqtskvJ6c+OLBAimt9i5Y5V3mPrkrM5dYG5Nk27XnaLvJ2ExpOEx
HdBtozAnQkWUeFQuANOhg5PtBoXbHRf01wcuK0XSoHO+B5cNmj6UCez4XfYUrJ0Hpz7v5XKUIwsZ
KRO1puemjShTaAkBrOi7ONanWpJj9/BoyipQAY+mBUhNfhnF2fM2OlKiKkNo6eMzD4x7qTumRADT
1S/Bc8YF7krj53qSA0dZ98e96+WjTRjdm2pvtBbIzvLIxRvMdyjOAQBHqNd/I7O+/KF11UyfUX4S
QAmeH0/7qUCV8V2TNi3b+3vLnj9Ue+0BpUv37Pn6P1Wo6dcbY9OG/iatws5seFEuj+qYirsfD28h
lKmwVQESxTNN4y4ONyNPWSuvDSseFsxPxYZY7N9leuvsGCfn4jp5E8uRXXyiXKL6eRsuwmGsdrC8
wvvByuKnlt2BYEmbSArwosVIhvbIBYNl25+gzJAvLgiIH+hvMoxWzYBulw3weftHFpeCmXHOgu7u
U/FIxzzUdrBDwiHFpsZvrLg9bkwELJsglzwnXkqvB/cN9dNFzGIk/WJTPXu69P7Kg6VkM64NG/Vp
cdolzls+3UEYhb0ZL4N+K9Mu3xHqFlewcU/3Kr8ZGqJ8qrrRvzAZk7s6rmdJlvBzb9VeJmzK034n
N9yL10wLMvm7og7XsTV7dFaPcc+iN/lo4xJqLes9WW9VxcVqLWK5Y9+3UAQilvNxXRFOUKwiELAl
KGSj8Q2r6m/8aARemWrPe6CfE7DrWS+EFcbm/G4usVuyc0p/c07E3AsPgDpMwWEqE/46eA1NMKQO
Oy8EzU3mdluOugQ98svLomaO9kVtWS05jWLzGBcr4toITTkKLN/FM3lhGx/IpEqKxvJHAUiaZZKz
Rts+hdoVUz8qZFs0+4GHRXAIM/hylFJ/34yRGP85hWg7H07tWldB7XoTaLjCgCUiYPn4iLtU5I76
QEFdUQy304UNR8ZCCQaz6IUNAaAAQIVNKj8lTjuBtooCKdh6NB6rrjGrKiYOZpZfXlJ06KVBkQrl
c7c/oP/dpp2Wsr7yG+ZTanLiAR8hDcWQjShY9FZvtmU7iHfQmlvCA9kXWog4ozx4GF0+E4cwyIZ9
1Yy/+v+fNHpz2yzGKvTR8N5Rq7YbqdMeXrWvHUBnLsF0TiuEY/eX42T7KXGo8gUNOy9maane8h39
DegGnx5v6xpQQa/aaFrfGLrdclOixYIPbRjajESTibL9/MCDu20FmgRvYWxcuottVOXPSAkkP8HG
bEixCHqbHJgwz9ok3BY6ZQj7Z6Is+Gzre05xjrKens/gvF4FKzAheBzaDSNPyA9CEmia7i2i0s5W
KF16xieR/boG92QWuogByz6zep5e+KNviL3yrAw2lWWIaD4apQZRc2FhItzrbbg6Xlnj0AO28TMh
DIYKvJhg7vtIv90OTHRmqsi2h8fQ18S2EhfXg1cYPZqWuIjuAfqBirD2TTRb3tc8mHh1sOGnNoBU
J0RHHJ86jfvzQoKTxD+FLxnJdKhTVAtDbO+cYfVUL0btmNwuq/76FFQ7bS+bBXRyGQRdWIG9PHhT
2qXatFOt7pG2Jg4C8iq5awIBPn5AFaMX5QXP34XXkLUHqZLoIc0q293mSyNUZ9ezMi0l7b+mgiGV
StGry/dHDpH9SZy6AJjafSLP9ol/AVjcF5E1Xa1rB9dEYlrqwHHEKw8V/kMRlI4oJZQISahuU9L2
rNqB6JoAVjVXtrtaD98xAL/uXJXPckHJd6ba0kkxOYftKv587UYDe5Nyd4+s88YK5YCc8HE1Br0d
6uAOvuc0RDhiatrsLNJWbCyeXXfX9A0O6uhk/YGbBzDplfP1hTi+rMJD41ZhrdwPr7lCqGw22Jxy
OPTx3gyiD+i9ODvG6xRsWawGd4wV1nGFg0YncDDhiyJwtIcIt40p7+5y5kUCfES2XmOWfCgnfUBB
ZUeClpKbQD171/VUFcGKJS7a1pIfyWj+EFyhh9LbEW0OM91qUq0FymSHoI5g1JLt8eJuq27E9iu4
sBx029cn7+NspfNLC00rDSRR3a+PRE3EX2ZkihwrCJWlUXonlQKeC5nc39rjdQg3nSf8KSWL1Tfy
aUWLXmokDw7+jLICiANNNeQbPaLqpkMWfoV4/Iqe9+nyD3J+UsGtAo7EXxC4CLIf1XJdumeST8xE
zMjbAeHtGw/Vx9L45Pfzf9sgnX9FVz8yZr0c6pJVjuOkKrdZP4IO/F9gwv5yzEI5pPdIhU2xBIsA
ewyGSHU1dBdXw46ZVuOAR/6XKPXFeIF2/maxqAhV9pCCMO/gsoT36EbXsDOFiZYGA4AJA7EMcWUt
4y1rRmwi2utfzcOvDGELP93aKe2JKZMaaNQXm/Obrwc+dO8VAOMOGE4e6z/595evAo5hKE9lcLZG
2Ov5pSUXgTsKYdu549nlohL6kwZF9HyIZSBVN71d9nwU3quukgRvQjRzpJlOAwwTGCDGWdOLH7Z1
YGdFBvfMY2US2azxNLO9PqnZdXZY2cL9uaI6m62BcU5Rv3NK2Fxe7SVNvH/sxRkwTigGNWZoZVBQ
95PsH5ms+I5l3VyO7fHG9u86X3nJ+DOfPk0jZmB9KyV/dxFUKCjZLd4tcJxdmYCtgyKjhUexO2gC
UDZtX0yKbAXbaMj9ZriZmAZuL1Oa7Y+3Q81aoNxokwWWymtxLdNf0IFmW/eM+5susg/U9wf/0esD
JNVGDDgQEbDQdYRo5XeYmdVfx1/sQfIVV9QPwOX/NTEj1OIl+6Vq64LG+s3VaTh063JNoLj65gBz
XoLgfoq+xoqi4uaZsl4vpCsWHZX2YfVR6iuV/57gtvGCsCxAVUDYWfjlNNPNIGEcG9HgLlAmMPWL
3hXLvQYQ95kshqyrPDpl+7tJIE1jVMYij2jOvRgDifJ/UbEcLU5DvEWJAFSAfNDorhUXMpUhqpUp
h7Uy7oF3FPs840z0JcitGRT6Elxczx2mSo8q7OZm1dGuSR4SCu4ktWuI4EnFoU9ASBVK7FvIKYEl
6TLdPkNh3mTctqIugYx0aaduD72B1WB4G/i0CCXu8I40Nyf8gUvQ5hPCeJ9eI31r5nEAkSkxER/r
lz2c6F6wrBuaGnFB1wP059/ugtIlheFx+lp8OAZU+Tj7qpicgUdm6m4LKwTVxqD+lv9iNq7pO1jf
3PSRjugx2TwqOoep+0jsKhQ5hbIoaIbqKbx8aZRH55b9y2b1i5hzraG178d4whMyA08uOQ/zCjk4
qq792Qc5G+ihDykrWWX3ECC+NzK1WJjfdovqZ51hBqNZSVFt9ZiQPvQCRjsmeQgvdcSOc8Zv4QP1
eXk9iI7Mn3S+LeOA5gAF95mnp2ypdxd7Y8YEajg1WTrQW5bLfUUnQtQDlebIeYrqPKCAUbt5B1Q+
Op3fvl0QG1tzxuQ0Xjq4YQiRu14w5apMeCrnYDhy3K8yU4r1+NnKiwsLYtmVV7DWMhAk6BBECg6N
5o8LEKmtiYBvYUL7I0SxR7b8RSQTjAisy/XdL8LtJeQIgTFaf94cqbRxH0wbsA5eRUkpuVFH9pxu
uY2xgv12v/XTS+iXpDY6Q7AluG0a47eGcFVZ/Pu5CSbdNMj3D+E2LvnZO8Y9mSJ14FpHXaFEAI5x
guX3Ko9K6N37XZZIFV8S1E60zehc7eZctH84p8QoO4vLxP7podeJpuJ0b8L2uyKjU3MP+wiWmgNI
29eb4LtvkB4ylGPaRjqwt9+yTWSjikMFjLMqHkYXp20DeIFK5yc3jImw30exrW2YZ6Tl9J6j+KKT
0HnpQpK410JxG485gjro0KeoMarmRm++JwmK6AptD+EYcQBnLOIAJXwnGZGoLRssW8ZMXXB3zIAK
AUY0YcHnZBiKSI/K74hA5BtA1DL1S5rZTBW9sNkwZESvqegPbdEW4QZJRvKcXKpn9cIXDCBx0eXI
rujX+zdI8SXLKwuGTkXPVKJXrg03pHi85HYkaHEK/RRbcTtU5qi41HRk7Dl6eegR47OrzcT2Hkbw
tPZLVlvoqqjZB/8oU+4RJaig7WKsqSqj2DvyBNO6OG7IFM2Dzg5RBtQjzoR7FhWZO9T/ACxeG0dB
Bvore02dyw1ymDPMSXSwirTtlhGlFnPW9ek1H5TJL1oFmp4WNn2vPxlqOGDTAFTMf7mGEeDoVotj
eDiTnFnk0Npk30VIa+AuNOyHU3xYHEYIpjziLS/oEVG//u9PKust5ldJyIIKg6CyxhHLhZHgqxJw
az/o6tl1PT85t8cyvFZ6QHdIXH0GJkchDS5pEDdP6EWZ/+z34rtIc18J38McT+/h9+L8BrzKRhbW
8e0LI5IzWpVqA0/qCAlYKXDhIfnCzYdeU35id8/jMxHMW3vKWdAzwgoTQ4XYkJO/KM85U6UbN+bP
qIDrniEhYv7qdwBWIiJibP2hab2Hp73WKmqCiKbCEjgA1bW0EIg84LVFXSoVasaXzA45Sse7Uw4J
bFajaWSm78bYgTNf7gfdNr/Iya1V4mr0ZhjPltiWFDwPGBgroEeijyOCkLOOd8gRVbP0TdYoejw4
1G9fdMx5VSoM1fWenB7nB+qyRkc3lGLnR5XaplusBDT5PFRAMU9vxxjA2cfeKgVhL636Pg834S7r
e37eZbLz9OMqX3AZOEG5CCOuUULNnr+MHR0jP9Z3O8ghqPVJA7lUQBmF+nJGKwd2sx+44pP0IjrF
z8WCo5+gTOG69ymDYVtOntHHUIakG/uUhI86WDg8byPDLz8ZGIjF4B9FuIU71huDZkWfmly9jb3G
qhS1QXnbpu/48glzEXS8zGcoX833g0sA5d2PJp05zUDgO+XmonTnFTHTcWoeEv03DwO5sN7O55aR
SBbBke/UR6TeDE+iJ4ElZnxsHLahyQcG0BT2NAnIIOR8nfqfkyrsoefGE9nqtPLmEP6vnhdoggY/
YkZx42oGMdZ+OhoNyE36P9aTXuCBdwj0M3516XsWpK4V3IaQQE4yfWMV2aJ20ti4eKwCXERXblTQ
3KM77PgqPII2TcYl+5UlRMZgGYqXW8kMGjKyQ1JV/Z1Sy4tjnj0ZCg33jcKPj7mDrsy9QyfZVC0h
cY64obGgEWdHHDapqG/KCunf87G6LpxfimGdrZaY0S2tUXZKnUBVMp7a5KAE7InlFULpmGivi1DB
UQbJ95gN5qvAWlv8EKKXZvnWg0D52Gxufg4wvLT7HVI+5pcmCQ+wQ10SBIX+3i3ezDXFGWbxaOz5
gRurN8jn3vvD0Ax41CXFfyTQf3fFaIL+MHpw1TRfFAtqyyWfM3GiRdeltr2MjbDQSt4Mfg129RPW
9NqI04L/gZkLJmvpNjA2bvtp03V29RHw+ixyHL5c1hCPjRbauSxDoOqO8y0aNEUj0yQkeTMw1+Ck
L3S2bpXYuhq8DkxhBBu6V3hcRxsSOvhdEtU1DZUXg6y08jhlsW23CCKDBz1xqREKJn4cxAAFldS1
A1d73kCo2DjdkhoXusfzR9CJT/RfmrPCGWHHCaBojjKtHMJmAFhSVDPYFlPB6LroZtQcXRI1Ua/z
0XNxfZxUA7659xyAu9W1EHzWyWC+NUDFgPV0b+rlmMxP3EqkMG65XwvRJF2Top9p1ISJ2h5KgMuX
azm2taZ7N5D6NRwH7Lgv1Fz66eu6R1OVTOZ0yu3jQz2Sj87zcVjCwpnxo3K+SPl6U/0zaF88Vx/E
fy261Lit9ygNxQ2qOLs3FRJMOUJ30u7ovo/kKKtlxQg70R7z3NZC1JXswXHwXcxH5w19sQjqDewO
oz2/tmy7hxSE9SOvlw10Xf000K5UoAzmr768XGDD00JgKu3cUsxDbtslloSUcBjz9t5WM0zyForI
3AtI5cdn7wNLbQR8YuzBPSAj+v64M38unnSnm1K79L6mpwplefPnRh4CqJP46Zv2GlNQLnqgdE6U
qBmVEBe0BY/J2Ke88BLtfR/gkRiZfB5NjaQlZhSytlGbpyD95O7mgVs/hNueXPTxnTaXu9Rxowlx
KOJDCp6s6rjucmoIzabho2M96vSMqq+AiFEwcOJjOJux/jGU8tz9nbGseDxR7ucIjojbADFTFETG
zBs0jTpO5xnQ2IT72vj1hXCajM2Ti07cG1B0mah9JUqj2l1Vt1eLe+PHk/R+tutm9ZohQcynXo5j
+AdOC/9h7MpS2rv6snrdfeN0HUESHYrq8oRVNsysz9R47IRzJ+awgjcSOUOaSYFfEqjFtSxTqi4G
r7rR6QYzYb7Bz8fNSi9dij/KH2BYJZX1ZI+QLJ44aa5pRatIPnTOGGs8jH/mhhb0DapooKNapwlQ
09DJGlCc8uP1nrQeto8h3ZUOReioosRX9RsMMfTncgWwPkhwz7AfC43JDpoyQBzVK3auQBLO4pFt
+qR7vDFMTSMts8ViVXHgW8jhge5+j2Je403DGeRbTzsiR3Il21Y5WrVNMeLuCbHydzmFVhk8aXgZ
Q2U1uOLF0OH4PnY/Qo4s/P6jd/GOoSZ5hsokRblZkJybWrVQ7JGUBDLmRpK3flKESVm7G0qxZtE0
ZEcRFKBwInuFRejsp33CReiPlGkloPX5aX9lXNv+ocYRCPMe3loMKFDcD4qaNTqERXfiyzebtWsf
sTgUEUwiy9NV20SY4R+bljYvI/s9OSrW83wdnR63/XehA04+YrftzZHpajoY/qF8AOoyZPjK3OeC
eBG23djuJvsQh5cUk1rb3Kf5DdySR8WkimAiycAyiuO0flW/MAOlsT84AYTB0PB5DgTLl1PUTFb3
94QuEJS6UOyoYlWCqVzLvPOJEe4YK+qwCkdfZw0w9u4Nub87E2/1gk67YOsVp3TJydCv/a40hPbX
IPpMJLGHk89N1TLyMT8OBcomhmsF7cWX1NnKVA1446uBnWD2g2BUpgKCQj3tLXqEEzUoNmOWqCVx
vIzBdAWmlVGgPgPr1EsSqOlfZOgCGZJ2ovB8dbEB8UeB1GiLI5CxLJ/DfiCpMwasds7oyL560Q6N
vtkK6HMfwjDHolSp9oOoR518CJZ4cNu0EJZMpD2xpivAEdK/q6RO7sLn7Kyjb8vhXKfA9NlhLRwZ
WG7Ta6P+3UASw+WLl3jn+flFg+ucHUJVxSK8UVAgnad8CT+XCVaV++wS8h8p0mCS8SHeJTUzd78S
43IR5/wCJwEll9yC+VD06SlpGaAVSvEC4bZmGg00xSKY2H6WiRTe/x+HA/LfDv5dFfajMFlpgLPy
FOWdlwxmYlSwIO5KB0w7N00faPQo3eGIyWgg6tYAOs0IffB/KuYL3HtfaqmGhgmbgcqWLJ1Ao2g6
8mbJDXYm24u4ljVhgUGZDemoObUtNKQWVB5kXjPSo2rUAMgR4PZiv4wMe+hoKI2/mtCwHBxWxEzx
jtPvS5/ykzxsvrT0lLCG94Js/DEXChL5jQwF+ThFDtQADfoOuk6t3I/S4YnZQooIf46R+5tzjpiw
bS8Emp5OUL/ky3MvdFFc27Ogb1v+0hsjdSSaCE0b/UIxIfh8P7lNimJyjOsoPWDzi5MFo4V8maVu
NXEVgObUKmFDCeSjqdSyvQw1bEmFpqypW/zgKi0zwMIZ5AZZpdALtn3dW0lWxVZWSIS6rXiSkwgz
T1XbeJ54feL1K/nL6wmJP5NTzp8ByU1ornlKDKfy82ZnjNNTNK9RxuZvczJVPTBkTSrmfzFJGja7
JTXMfOvGFhx5ZbABCVDWbg1IW2pxotM0nypGBLwEFLy81EsNYOie05S8DcURMIRroOYbsxa4oV+r
3rT/iR+EEPxRIdfZOojyCFckmBWCxgiz20J1MrwGbdQu00AwpbkAa2V8d7hfpdqUHRoTatU9z8hH
HPyHVrJ+2EISLgZC9mxz2+pYQCWiCfLb0425IiUChrd4kZyRPxN/gBw/49tQfrd7A/mgQkCegKF0
H4IkaKf1JR6g3IbJ/tLjGT3tBrt3cJEBlgdYE1Yrs8zfPZ15bb05pm0RJF7yZXbJbDo1aRqwrpum
RjFHdV1PjR1gjVd8Nkmja4GY2gOqqxk9VYJxTX6fKjFRdhuKh3rfZ19xe0/r7fZNQw5yavdhiivZ
t03YTsd3hlFy6aOGjLegePu+Edost7syGvAicuNJj8tJmkcbcdHOnJiVyRxMc3QbkHWFlvW7RBnj
MMirIDs1Dl7Nze6rWulUG8SQCwKsBsYhI45io3JsynblAIVuVDlFEqJqmy1xE9qsiQjtBlAe64p8
/aZCeZ+N5yqLlgx4s8AiTY0Yeijs0fqyr8J3ztjivuE5XdVVwpAfbvy6slEgTqRX++VEBlcWOVqa
SKOVgbkldOq821OkckkjLDMm4LQffwzVwwjUUGmXZsYvpCLjY25dZZ/2vU/HZtqPRzZ3KiFzG3zh
VbG7/qD6rYKUOXCG8FBCwEWGjkPS8MQtA4kxP/2Y2lV6kCsFQJt0F7i1i8d5c3/D9n2H8T42hXA6
tdNm1ibAVAT3Nh+cJVHMHOl+xdbzfh1F/Lqa+o2BoHXejANo1JDVYtgo6K9ouM+DAKNWkFFVAMOw
M+WO+67G+NMDmko7GTWM8rU3fqeAoyH42jGeHRCsK3GaxCM0U6rCTha+kEwI7KrgctkdFQHVrjvf
dCGVYEqhUKhou1vK9GGQHYR6ftE/peMvRh5KJJLgEk5MGVWRniVi1ejEJm0JBujMT2lik7B7hq3O
oCUIZwDIVhyPMRFXvhICd67MOcWcLUO8sgB8E+BOr6yKbpkBoIA4digpE3mvxx8Gzyzni57459Zs
isTf2zx2oDYD4LiXO4ZqmzeYi+lXj71T/M/SgPC2vHrjCQO+0CsHoQW/b/yvSVeIGkHIBdOMfuWN
zsKObc2G8w4z3KTqsOVxTKnC6szqs+v1euJyc2YOO5oqb/a5e9H5WPT2StTShii5/m+HZ2zZ8bl1
/I5KxNt6g+X8WhNyCijDx7m1glnd+VDC1npk+CJUVU2mt2LjG1aco0YgXf6ikdvq77X9SFQSqcWK
4QLz4FgKvxuSJdGCgvacJMrZge01NcGXYRozOECWSDYnc2vZU2rzpsD8aSc8lBnF/zRKhNxxXEWF
YsQijA7AKEdAgJImCLqUy4I2lAui8Li13d7/rsGOHCZs7W1GeAnO6iWCArBbl4RORmte0vfcqnai
vUJSQ6e2faQhKpQLESI7x0FJPgI2yCIKbEfgQDA105/ANOcxXiTL7c11w43MOAanEJPbvi4RzS4G
iF/K94GuWCx3zCE/fn15e8C+U2iBrVqaB91OEnizGAgRxp5eu3/IKhPOVsuspGL6SrjC+8aL//pp
r37oL8m0dqa8LqRlNolKZLmN9L+oEnIomzVAcYRqta0eHlkY7Gaf2M92MXrIWd/lixHhczwdnk8/
Xkx1eC6DECV8GGqVHzipEj8R/mT52ASzmkkHI2Stp/kznp75e7gpI5rB0UKzzl23NxvwbtblXMLd
jiAZsRrJIweHooSuM5GmVIwlJA8Kb1s6S8yHT4Wag/j1nT82M8y7CxLQ7H85FMLe06oeUODiCb51
QeFY9mo/jzdGbCgGAJ0G8uA2yTY40DW/lEgoqjrjlL3O+B4r/oEBdQ/jdD7crIDHH+0EPQjlpVb6
369N4cSxZ/RpFwxtpqydSIzevj7tKJyLkPLqWvz32iuAiJf5orXOwrvWK2vVikUQ8k9yTh0OcsdT
xK2pQEak2SN3V7Q2Y7fxIcM2JS3ZPZIuI3nssbAurwDP5/yZGWhupmLaN+46QA2A2mjG0kcbMyyc
zq1Epeo4mDe3eexZrD5cI5PI5FslczO7FS0xawgZ5KVLOWL43yLH8jhbtSH7gNX2KG8imAqLzwuu
wjm9MZcszsBtt7v39QLNNkYsX3yITJuSXPnQnPPNmT9rqujNrUE6BrnMPTDO4qZXhBOIRZnKKHpW
fuS3AlVpGMx3jDIgt4WcCRJXP8PCYszSKhqSPrcFMUgRFRCL6bn0eylMN38k5MXucQmhs0Av5ezP
a7rHEnPmhFiAXh70dMSX8I3F7ZhqE6xFAgA2f2Sz50SvMs27u7D0eKNi2LLbZ2IHoLEj7JoLmGHM
dX9fbfGIgD14NVgRALjkcuW9XByHfdAjplyxvsiK93wdyFM3qJ5VnpM1Itm5zn5yqXYa0dEIrVHu
O2CxtEI4s4NR1Z+14d/BPnjmUMTtoH+NlR6s/D7No3UgZXK1zf/DjdYI0PojztN5v8RLXeHvD/0Z
ot0fN7g9/27LPk1DZiJel+wFpt+hB/PG4QHpu+Wo3ZifEz4B1NlFD7ADL5QBrWiCuMTVeZ1uElc5
JHOAOIpRtVJGwCi+oS4xR7IQCwbaMJ2rrbkTTfRudk5LsmGk3VjU4cBFXxHi4kETENASxCHZcalL
EIoBMLYGVF1BkxG0wB+Zy5I88A4tNBiMBR1oZRYSrdUYcdm7PbAu+OXeXW7W/J+YW7NGr0NoeTWv
93mSpduENkg4Bkxqny8ajP2NKOR7Mv2i3D6ZWZAbrn4t661fu4nkWcQzFBjhEidmeElXQTAu8IDH
ErIFfoZgh4YeqB4Jwk/fSH+8jc8q6y2DQNlGr+Pfx4Jf4Dyhjrs4QsMXiZd99vM0Ily7OPb/8O+v
oF63uAXsjK/NJOll5sHJkMymf+5FCTdPc6V+6yNSEWJm8J0Zibn13xgG10ew2v6YnHvCc3whQYYM
DnCSVxzQKSY8MhWgi92UlHbcfBKmoKFZB6e6YvZVn3zmn5uTZlAnOUMEiNIk0Fve6kGg870FPc/F
2Ve7eGnjxJcVtg4Av0SC8h3EeTi3Usq8epaJrxksua7geNN10SvYASxFfVa2e3XCwe65LLK2vLmb
C06JwHmMQ7TNNzHdXFEqWkOK71VP83MFlirDVc89X1sbw5Lm4HzOdXN+EQrgz345JjWHESB4cBRc
vcvx4wKz9iky3ShoHWMLDAqlmKItByXT6GgZlqzOBaOOhoP1yFQIOMDptlgOQ//OFPA6UXiENsUR
rOWO4w/s8/bz4cbZwHtHoGY2BRjMEwzX9pruTsbu4rU7OvCDfKTFmIMAMjmnMH9Qsf07qpAnm7IA
6aY15O7PhWtRZPV4QF1WKfUs92+QaBzvK6Yy/k8nlnySHqBO2gc7Z9d50y25kCOVq49g1ALClYXf
N/LaMgZ1wYxi7F9Xbc2sUCp91b14StvBRqocPB+dadsTMoGxpPfzOYw8j/dpkgXI0x8v+gGTIwTO
DPlvAglssE26c85696sQXaCrzXOGqbnjA248MOvpSVcsZElXKB5aiXA0mAj7JFAJFKDmFuqhoia0
6VmBKqH65x1GjJ7GBmNhc0qlS4R9ZgBHNkAzSy8pGOIKLj5cFSfbaIwKSJMQMuT5hhCrDKOFblvR
aeEb39MERoMLNmAALA3trci+3+gpjn5eDLb/9ceYkJfHQkeXdWJTjfg+pssdogwNffUqLUqsFAgX
vwWvfqBMQ8G/oVirMPQtECegTKY63zXklt9X6MkNvS3h14b+NOvZxXNYuKLoJlLqtbYaVWXJht9S
+rULVU7qNrI/3TVJzqml1WKoSCgSO+vW/hb1gTjk3GmOtYUXSNhINMyxuIcmCFtXT2rUi5QUUxP6
wQmMKCMIxszVfkz9kRZQE+N44oZVyfS1AClIKBNf0lK5KDtK1uMi4XgswY0eowN8LNgTR1IUUPJg
gDAGrh3z2JYYbPL9Smz9laHQ0uUtxJB7F203GyrIdwE2krjRCR4J1JhUUwOg4W63QPKbLSfbdwQI
4qEfNA1p8fHmZIu5sT5ZcHpWiIdYUKK+HA/4xevPWOOrDdrWjq6QxK6F62SYyX2oe9T45HQ7GryB
/ErvlivcomVdL9RAb7KYHkiOV6PExT/sxV1yJDtI+c4ImnfdAR+orLB3PZAce+3eNsBDvGsPBOj+
cbY5A3taBkLgJT8LebkLKj7tYhiNQ4WdxIqa5+cnKWfw31ze3so0jyjwTFSyAigEfo/wTv8k6zik
dx4OLX5W8C3Yt8z1O2Nr249bh6k+FD/xamnbkTkCiPl2eyz7OEQ940iFcYzF0FhETK1Nj/di32HN
Oy0ajJOYHZKevnS+jzQfTZAE95eNGLvw1oO5lo5xf0sGSxW9GJWo6pR3vkueTvN9PJlQz7r3Uq5n
yQwHKmOpk00ZqKqQbp47mtcqPaRXIecrfykdW89fdkOQhkzk3Nv24FoLGUQ7GFx+mtDsFu9EK58y
Mr0jjIG5J7fJztBpxb4W1apoHVK/HarnYSsppiPOT8mLGlcRDRyo5kDVlJA13KCsJRtkhGTucev3
47STmU3LK6N455Wk0s95eZpcEE9p+4sR7abHUKs8IKjPx1lGKZXulGJuEfGCMPnb4/VuAfjecspG
KgISIUoGsjCLnapB5QxlFIsifD5DQa26J/wyj6AEFGcqbLArIdJoB82+JNmOR8znOoy0sgJuN1g6
ZnyFcryk44ToU8bDAB2JS5+vRVf0elU2xUOWrvF6kLmppybbzF+dVANQOVdFUZoZ33LvJ05SCCVp
IoTDhoQh9CXhdL6/OBbtI2oTXLJF6Zlv66viQN1EHmU7lmLLGftnqP8bA3bnxrS1xpF6LXlGcubk
W9Tt8OBYqiTTgxhSsU2RsrE57qCgtZ+SW07vJjsc1XyPJXAnNuMpRzkC0rrA02pkxvwtWvttj7/P
oo00DTfg3zb+Invlgs9/Gr/3uI1dPdEw+Pzj7M/51P5DaNGKDbYcPonvCDPs+cILdbkjyB4TNdBR
xlel96L5oFHOJA4BRkcrVwYc8ETrzrrFYEFrUjsiFVxly9j2SGqdiXxXVSBFKBcsdtdgqFXr+h7h
iYJa6nRmUQT5H77wXehykzm0CZLJwmdUU/+R3SahIK5LUJMeLiez30xDdqPd2XVD1HPrU3qyC7FN
BTGj+e+epqItwcmm3ZAnQnVni2pqR1ysHjeG77GHxYa4oEXYzhJ9a8GEjWovo2Y13RSho0vJBjy5
bBrwG+VO53q64OSYe85AIJqFeiOsLAbyfGbhJbgW+aUyPaNTi0bY20g1DpejcNxSym6TUEx0aSI8
E0NVr6a5TIvOZAUmcFlJ3UBLHw0ZR8+GiaAWh/IjcTDXQT+alDTMp12tg/CMlXCqpllmhEXt0HaI
17C1Clje5pyaEnCgzCX9rHOBxrLyf137/+9pJmrFExDHj0qONc2HRCNS5r2MnjSXsen+pxUOXJlR
G3QpMkYJSixkLPzfI8FptJYRJwRFCmnL4MZCVmZoEKsc/IAkyuBLlUK1n3BfjIquK8HtnQkxz2Ru
C/uY4+ntl+ogfCw1sAcJgzW9es9eCDJtzw7BEQ9xdO2zCAsAg6HLOLxD9LXhpXrRO6TMf99978oY
9qPk6DC3wwrtY97gw2y90zYcx54I2Yc1l6g/R+r5qxaMFjI+b1UxktHtuTJGeZzZm9bQQQruzQx8
8ui/8tW9Ud27nHWoRlx79dh6FR7mS+sqmi/HEzXFnzEPGF0L2N4zCo8a87Cm4MKmh78KRUAg2dUS
gtmKFVCcoaodcapskYcyvR8/pnfC+CWLGBKNit45DKxcfXCkUca/7z2vJXJtKtxfLIV1Xh/2wUsN
ZrUXW+uVtqvMJGMLHp8jbY/Inv6ZDAF7l/d4YqGUA1KHTrWPbPZefjSd3oxarJrxH3fvAu2ZERUa
Y/Sssnoby2iRAvseCKI3xj0j6sDlm8EQl/a1rFFiLzjUKrbyv8bekz/0WAJY9Y0gZa9hphmv8Uzo
GZBvzMRjXLtdI47dXQlpakaWbSLBC6qe+9U6tYXKzyL5leiaNNeYNl5lPoYVEce8g43lMzjVTNyx
6ANCjz3vPxwWKmcsoqPnYtml/6fqIWPTabc4dtXrrog9sZ+pq4MH2rSVpYohTTmIcjYYgbLiabPC
MlhYtP5DZuQGOePkB6xnS0IT+KLkekQU6/LVXRGeg9pcUh9lo+NTjb8ezn9SgWYwTRT7wuRMuhiy
W9JZEQzGJVQkQ7jurT45Q/wxrjqqzio3brJrTW5bhjPj4A1WSrawZYQFTEip7l6GiasTN8gkNTTT
6WdHArOa8DUbAULNjcOKmM6jSTMOZZTm1a4K7n4gBkDu0OgGOC7/dhbymrdZWg5oRMnpFDazYmzs
uXSxUKcYNjQ80UJsj5+e7OeJnfq5Py1veP/N/fjhg4G1tbkO3/DRvLunNoQ+7M/Gb7kuakL1g4sD
UHBwhCWm4MgVCe3dNwwslcIJhnAGaoSEW8hbqYVdza+1wpAu3F/39B3tW5Y96LJl0K6ZW3HhjJZ4
b6jCItOTjBLYU1fn/0ZEpCEj8RcxDKSD4F3FkWdKKAKPjhirKZ7PuXsKbrQKZrpRgyD3HcnpIrqf
2qiPFoYe3Bt38hKvI752WkJA53neQAUz7nraEmwxExgDRRdYxacG8azpLDBCYK3Cea8yNGNKPqWk
d2JuojrEs1zdlUyZlEBKKbzR2RDGEcEhcXh9JvXkJM7J6yA4IlbjaOpkiwc/S2XemaTmjHKgO9yl
1QiX2Ivy3sWWVeOjHEk+H3B/FnAx5SV/N2catfxmYLVu0GMBuWy+xzn5rqXYreznktQSiuk0+PHE
zTMhXeVZlk2Ba2wnd88Z5TYgiWflROcqWx+CGXLOYyjzJtysOzVcF5cgjCaNAL54FLeTZzoU1i/o
FlapSaYXQ9PiWLgy5ZcHkCq0Vq77WlA/779/FuGMg0vivo6ml2mM/SAoQStNceI5i2Z3B095sTV/
dpkmBgc7Cm3BN6KfNHBH6hAyPf+We6xiPbf6nFNzlUghpF84ytSJ7Fq1o6tS9kYycyX26soj093M
mmMJHB2Qitk5W67LXW2rBLnH74sb371ubi47PNys76yEcwuiR2HCK5UVATahg8kXAQfDpq/0k2tT
y4JUbJYkRHVMM9v6oSzPKcKvz4p8js5US/tWoZ2nibZwYvRWKoCSFk8ui+sSP1bfh/cDRaITnGn0
kk3oIC/+yyb8PPicnlR0p26O4dhYLquSAqMqcnjSvk6H/5ZPXiY6FZiIAb3jimlftKLT7PKPVhe0
sCtjQJspcGZEe83mZ0y1sZUBJOB/CH4p8vukQqly19kxMxG32rxWXH+QuDVXplokO8cKWi44xD5Y
0IYvl9ss1ns0JG4QbJhCF1uiZkbMsSrNojDX4wHGEH5GkoIVlyQKDvqyvXwoIXOdeyKo/VaJFwtL
ew74p21NuqV5lrMXPIBSAEszcODgO2LZI5kv9EpE+XoUl1VDvmqBF1S4ZD+Fleoo4oowiAQaH8UY
hU4ZtMw4sKyxmWNrIxKe0TZ5gm7DIo4kd7YClL7x3bTajE3kiRr4ZN2C4WGKSTCtvY2x/aqZh6Ii
lRBbBgGOLpmQqng32dkMed/far+UzSF98QBhgebsFRuSAh0ujE8poeunjUqNsomhUD+twmOBiKQI
1L9nG96bVMGMMHYQ7GO2fiPCJ8q5xM0YgTwFhfdyg/czFREolDrjUAsb9wXmpheGD6xXvCfPJ4qj
gGRBuztPMp8+HysL+Yf8zPGSoBsSbBvC0dMfXut6QyFWK75JgQ96XnsCaJ1AK5SEJ/KjgjWwjLxA
aC1km02F1sToVAv1ws9kFpO+Fy7+Vl56t7cETFmKFvtXEDiPw68M3AuiX736gcv/jOWf4HRvDRwj
QVG9jbeO+e4sXKYlvogzaCBnFuMxGqwnJNnppwUNhddfB97fad5legZIcq/VDAj8Bbjm3YC24NeE
F5G5fHfAcrtuhc8SNbto46C0ixb0BYWYCLzUIo/mV8J7tS2MfacXYUfag06gvaXaNRfpW6rQspjd
AjqkgWba2fGzvosACMRNxrdsKtIfO8rUVXF2XJmTUO6KDvuvEpkcbYQ0nQIJ1kH6vQGCF7WWJHbl
5sT/zuh6vjmiqD4UYfiZEwxtFXwkP6xFc4FKRJn0k/iEJQLUwpqnnQjQtmca0A8CWpbZFmTKR48R
EisqxyhvUUHulzLOkdkp2G5UkajAJnpSqc6kLitZKUCNLcfiZQk+wvpx3Cjj6pMKYeGxksdKVyq5
YhBTiWVDEFTWbEHY2VH58ek4L5/MYWLVmMNer5AEdda18Yj8cL6Kjlfu7lg73KOisb++Q5fDaAco
lBPL+o3MQOwivlaldT/1BIeXahvrlXQJnYhUEoZC/gDdw57e5FOD2hOkF8MVQV4jxQvbv3qx+Quf
SG/tyyCB9JL65898ExTMo4s/Oi/4fhLnf5SjvbuIZIEbu7qElABz3syejKnicqi+85IkVn6tKW1K
muagG0qu6NRYjWajm7WGXT6IY7qmJoIBNevZX2w5eIUxIiOW3sPboIoY4BMciZit0gL8ejGbYTes
uYXwpLFP1FiHvqNiKyElc0BG1ZfDO5ZYA/9K9BoaEcYpI2QqIL+fa7EFCgma7BQWfLAHs55YMXoQ
2/5oAHriZPgmUptS8kcFP4vqpjW3qX2JKwU5ykZ1rADEG6TeqCbycKpkM3sX9kSgO8fF0O5tsPVv
4ujSqELzrwwGTyoT5hMOqQlj89MB5U2DThiwbM3rYnbCOgU0ix6T6HIXSH0QuOCRtrDujxS0eiiU
ble3Ka0quKjK7/UuLxF1bhyWQ7EAC9Yp3u/TcmoEXFaL7rGXnw3LsI9gBPC3A6aiAEbTNiq6sfUg
A/zpzvgNQrV9ucEHLxljbH0adohgK59jmKGzeOnKLbdOv9vMqC1dF6Cbr2lv+3UK0+Jr3/NqS1ei
jALkuqyvqT4wpMMlyMveoXjuWFOFo8ZarbJ3xX0covrgA01325BIAj8ynDSWiEvAqlY6C6ysLBd/
fUReTgwb58qEnLeN0Tc2SWu9oQxmLqIiUU4A1dY3RaTUPdYSGSj+zxOSghoB/Y74jGOoC0NhA9L8
pQKOAW4S8D4nOS84lTpw2+ZM0Qo3HelaenQltaxg+AwggcF6Jg9VZDlB7Jc3rx/aoNkVpExTo39+
ckTHewExNEQuHEgBaVAk8LX81F0OS0obKVTQN4++SzSzboZ5CrH7Aqomcx3x7W+GqP27iObr2CTR
U3W3E+i9jba7uEEroYqxGHNJdrUG2ZZwz78BEB+pMyTXOPrY96C9VC3qIWmSiyAillITejaSKVpL
14gqemEZPn60nGTfyWoRPby10thfIyTyQhwhr1tsYu71AsD4C+E5MCe0ncG/HGT37TJre7qDy1uc
9D+dLIJcsdsQBI37lJS+Dlsz1gGOK8VTpkjEXeLpY2Mx7bkNQrDhx1Otw4jhtKM4L3I+8eWZzxnK
/Z/SeLoz/LRYW9th6Kpe2j8/ibUtORSiyjNb2VXgZ/7VgCQrbMfaYCg0WsSJyuB68SNEggC0EJyE
1RD0AnBRbLTgi46T3AzmAqatJI4+WbPrYr2D9pVuQo2rneGkeCboxO6zRaXtbk+lZYqhLNSLP3lE
7+sd0eWx4/XqdAQCrM1mBb8Sr2TmPW95cgp8UUP2Xgx+fGlb5ZNuNPKVYCD8SvSUG9lhNt/XqhQK
z6QqmwIG6PuRxI94jQG5hIvnU40pBknnuDTbUPbwmmiqaSqzxglkWTWAD0+r4IAoJTjbJC4DQ/oX
3KOUEp4t4q0ZOIr+imBFzifiv6U20VvDB9ld4g0O3mqnaO8AIliCnEmC7rTuieLyeMrcxwNS51Ft
PmqcoysAOS8A7RJN6WBtqkZx3roYbChBg4Lxw7hPkUu8dEqrAl3IvE/+YubqGx2DrcCtUWZUUSnB
OvKZZdbczQongd1gHfY9TCLWwwWDTkbFvE433P4gltnFi2lARLYTDvbZz+MEfIOWhLXzcyJ6C0HM
xg47YdyExl7FhumOk4zkxkTuVNmSc5uGmNvEzZk9urFNjOwb3InJFkBS2L+1mHlxplSqeM7LKDg0
Dia6qhbtfKsr5PHkKik1F/mtnHSBfpm+MF/QkkM+86a2xU53+ArDQ/ZTnvaSNLcE9wRQo/lM67Kw
n9Si61DPv0swVk4+ycQ7r8+4DrBt6b0TYaQvSKdHhyGW9VXcFnehdcQaVZCSBMXH82vLz7qejqmD
EiVyF9XxBYis8iBrq97BGiZaEq5stLDrx67HGzjuIvN8bgY6sk8AShbgvIdQch+3J+J0h31ryekB
hZQ1sVov8dPE7YJkLBQzSfM395o2q7cFCm+zD/i07bfpkeLVaTRqRGoi4nLhT7AEtI65Htyc1BkC
CN27Hac7O2a4fVOkT0+SxOwQxbnGG1G86UpRHODZbAywngn/ZgZ49f7Pdxi6TdwOtXXTlZ12YvXw
fGi7/zj3NJEpLMhDon9hi+ROgQkJ1lc684fev/vyOU4Ig7Yj6X+rgjwZUX+/iaE0J37rG0xAnG1b
JrsklGXF9ctWpvOzblQu7TpWa1azqCDEGvGgoWZj5XdDE1v1i494L+AEHhUTvWjnoXqLuSU9dxu8
djphuCy+7/dJoKYLuBIuwzPFBuPKEz87fc2fkcsTZfZQKo/hK/+etZIgirEMpPeV8FCYmqoNVPbg
mB+HgxIgXrccqAK3GzeJyNr0YUlvbYlcF7BDyYgQ+r8WnjNDc4TqfSWHUigiCy054xgIPGEzuXy8
POiKEFdZ2ifqwDhlyvFR7HHaQT2KEj/GChQ8YOBvkgqEtOBRsgVuIKDxEXqXfBk++YfOtIPupW22
pxtOLMEWSWgvTfMjirSzAZSq3C7+bmOHRfxhW2JtAQ+M7IVX0rFhQZ9VsBZFiaC8lEkhQeAUbnOt
oVsTcSWVG+a0kFwVDQbmMfFK5wQtN/7i2oVe38wZmJJjw160r9LIo8KAsLP8xnNkJPt6iA2Fx8ig
8FzAbyLYIaiRS2fvThVFTEf1f81ypE9HmE0KE9CaPjrYIEozYpm/je6pSw84YoLTqpGKxxvXxp9w
+KH+34zRMebUL74/cXBSYBQZaVzLXufo2LyMYeMT91zYRP7OWGch0lSRN2evrfr/EtOy1vXPt7K5
gLl2LkBRybloIWV1safq8s9efoeMlAkVAeFCJ8jKKydoLY9cnYieVRCs5LF1LvjUVU8lOJj1GQpj
g6rEtS+Y/VR62Wc/ZPsAB6xaBK9iuKZut77dNQdN8pclyCzfoGMsE9YO7cgcE5nepHl8YVGeJhSz
1E1SExS8/JOqlWhEXrp7pFVLa48GmpIH9tUuCN/q2sLKK8PzoTpoyj1fcEf4Dzhvn79fSW9AXR3t
/9dGZh5DQppU/zBdVIbziForJaETQicxkKZzWAeRCgXQjnrHb2qPZo/Ood/CMOqNAvZahjbwgZJ3
fgUydWMk0ztv9vWt26zFqO2DbKms5xGVBrI1JhzBzexHBSe/YVCfIyauBl80f7690ZQ7FFF45eK8
S+hZ41UOVsHRqLs4MGmF9vnGptDg/Q8UHDj78QbCUwAii/2okXwhk9gs1zglAR2cR0zcKu67t2fC
jUB5lFK9NQL2oML3J1CwOJ2iaZKhLTXGst26CAKOoKVCa2P5ne/brWHxf33zsrUIdvtbEub3xaXW
oKFjeyOV1X6gJlApNoTGJyzaQM7PlqJTyHZY6SD0xxQk9Bj4f4VyJTKutaJ+0y7ETnk1yu/BwPvb
W0mkBLKLFoIuRYTkEvOLoYRey/mC6e1chGjymYLsq37SpbY/fhsd/lr+rNYvPC7mcDlm7VOlUQRc
oFzTOZYrAZ9ij+kSX6nXnvp4OPo394McwqyBjQxd8ABKfE+WXTFZzrL5TecuX4tCY4PqqGH8KABv
a2H6RFSvZUT3XXWK/frfN1vzpr6L6PxDxIekI9deT6aKXQ2BSEpKTHhmCKEhSwohH4FsFxcf/zEe
U+g2THuBOfnRM43UPXyPQwgrPX1NfuHx5YoqceePrWXnEQ+Z/ztSvzl3cJBSIA8Px3FsABWoB1xH
p/lUGwWrUHnlCRh+puDByqmtWcCbya46VFkh7y1Vvu8EUHSk5qjPTCziWNEDADiOaUKqQ7xyLo+m
Dnba6wftPtheqKYFpWIXHHez4fAdt6ptvvednqsIaLw2+WtSFQhCAsRWTPNo9htEzR191vSx/bVm
E1R7rWK4Z+Y/MyELetyELa7bgY9lk4U5mFBDoYIsQI65xqJ5lrozJ/9LaKUwrkfqK7jCaTQ3PGRh
h5MHuugffkKJ32U20dHsz+MTCpRd8mL/mDnUJ3LtRXQTD+jZzK1MklajadTbhUrckozbVIuW7FD1
s9urpakMSsIzg/PJwMNhkPze2ilIzV6349ZRvd/dwERdJ/rRjxNEvuKfd7nKTHtDlDVYszA4UdaM
lqIQoOuJ4PIa8UEEkPSiIBPow5NJHbdaEhosIQ+bnZ9jKXkVnKI7IeyV9uYqDLRiuIWZBaLcTZ+O
CnY3mSV8vVKG49FXUTChIdB4DSFleB6tZUf/84wdY0dMgxn65lALLIOvc50sTUISgmAdCM94cMxa
p7/oRAxLii2VSoZ+Ky19bC5gV2Oc4LqkX4IEbbod1ieMnWCqk6yqM/xQXGxT/+b9D8gwO3YsoODJ
TXTkWyUbtbpZsvDMuidk+IPUYOjal8ofwuBTWsfVD+eQXDB4ZGT0x/3tPVgCXkInkijPhrfCibB7
niLu0b0BowQpOhQuho0V5x9K4yu1IAWK4pCfdFAFLcc8Qb3DxNerCmis4aj16+ncB3GYYtlBVVJt
ldwupHwtzcK+JB+zbYijzWuDJGP77rxu/FaDFsa8QzCqFvZkC+3XHHadcPBPU0FJrhZ6/MQA2Bbc
MiNooYOOyDJykGqwWgzyrKj5iH10RE7jIoyFAkDuD4XP7NAriHbaNk4zyTY8d3X4GK/5FaeMmuCK
m/NDSGZrLwcFYo+2AgPW9IVVS7eoqsBSvoQQxk9A6yVG00QzXjoncbn17fD6EE+qrU77HoKMnvJG
tAHRclIAzWvQHBxSIvdH+SDhRLxge1DahMXMriS1cwoiwuRnRAErr+VUGqdbv+scxHt94ND70vZa
sgMJRXFcDeMHvp5HYGRQ9HQWXlUMM1+xysGTpmXPs+9b4Um421VzxfkpIFFRZsbSkK7OAkLHJEya
xDUkpcnHvdG+G1E0FpKzm4pfojC6yt+nnJzrbayDEuAx67s5mndp1l+tfW13SmTWHwbzWh2Ggm3U
iL0whj/OQh8ZNHLTEApPXrfsbRew/t566tC/RyU4NVLfI7SUdWNHZOjfveH1tDZSjUuDB2cVLGay
cRQvxHqMiGOxIkN0MER+pQiEtKHO2NAiLVX5yIwnIF4zF9EGKNhmfno1k5iZkrdmR1DdINQH3b4H
rxyb8kTTGjkijZdrdJqDcL2iXFrr/a3Fr8qdez4tiWykZsnjg8v4Ggkz0hBSTzQSHmSISEKGrTtT
8dAjutP6P9qfMmmWwY+Muf1dDfbH6l7xTbNYjpZCYONoPw3t7VIAxHgbAfMpBYznW44Pkl4HH2sl
BYHP8seGivqVOLGaCM7UBMypXvwvSFNodNXXNZioYQYymFViKw7whARgrQ5MKP48ppIqM7lYANgE
mhZnq4CyBQ0oRL37k1AUpONOJxk1HRrcq8PGLKkmTDssD+eYJyKhvykkbwEMWWNyWZSeW8IE6jc3
tH6Qlcqu9gZXHs04MITr9M9A2EwgUxOqWBEZ1xpCTKdgJEVSZa/3JJfAXqRnW4Bri9cQwlRKwuYB
ZSXMItXwoiLxSnk0+c5/k8ui9Z1GixaDQzriTCZX9KK2zJ4qcQtnaNaZSzVwrlkvTT8fmbS6Dem/
QTwiV093YduAKzzcDU1EP4F+esRDvG+MOmk/v2oyAjAj/9deVUBH2q4Oq7XGmtmXFpcbazaBct5R
ubXfWsyuaayY/SEEClksMs4EdY+EXECgQCzd/hOblHTK9nzRWJ2kMehxhMGIwqXzE6cEcPmSKWgs
m95sEWGhR/HEcsy/BOvUnUGo9+Onc14UK/+LHF+6PR64pVtpfSYWyGHnS/PjtzI7/4A9cAQ24H2G
kFTNeXwvTpQ4u/ODxGDJcKBBtER9rKG8K0ILjqS0TgXF2DEvOy3QQW3Xe0c+TtIIlzoq6GwMyc7S
cozvuhV/ff6haX3gWb/BgYYjcBiefi/d/fe3gBmqRFZgm+NAxmmueD6PS26wfNHuwHiE9b3K7Fji
D59ekRoToUiwIO7rs69KN9IpFDAQPhBWhGzQ9faU9oSLQfGko43sPMd8u+idTF6cl1lfGH4VTWf4
1BBfCtmiRifyDDaXU3UPa9T2pqbsuC6e74X1zFyoZh1qkGe9lecaYFx3N6JLD5iz+v0V1bSXnCLd
o2NHO8t2YNEb03NrRWcsZXyNPaZ93pietIAt138Yu/zzqb/CFc517NGH1zZzAcapR1n4IXupMu1v
S5Be89kCOumCErGynV4i73dAAAT6ihrO1SqDobueaPas5PZuge8Mr53imKNSgu6BKc5RgwH14rEM
iG4N5MYdVbUb0biCs+HOJXh+Y59C+oicvn4JSzboCeT1RNfwqrNhi/qt2Fp1yIvxpwkkyEFoxDV4
ryIN8Z8fpsCBv/C2OlrruiPaWG/ko0nyWKKnH07mCMYI5rkOdUkUNVuEBnsQMBefD0KujV9ppY/i
TW5/Ye/DeytBPi09HTfShVVO1mvRjCMgd574Es584iZrcF0H6oqYal8YeogT1rYuDpxHXrZL6wWA
o6O2qCQzbVkT4hGMRkIWlSCGskovIfOyndfscSa61uvcZcjFCfBPWr5Lo4JpSGMwUz+0IbihHuwg
ZqdYED1QaUpvR1bFDSbzZhQYqv3kvrMQmiP7nxcpOYZsx515gSemQfW9RT6gidBBJ3jS4p/gZJZS
rDamcVjhT6nWz0dFyU4jOG0KptL0ME6CXk2zNRhGXreZxnAD3aUiNFHBU9P5+1jKzWTwp1iWlCvx
JSeaolSYmY1rlCmcG2Z61eDgMP0n++fZ+IOI9o0maAPpgPKvijnVtH2urysWZM4hcZjEY8XXmds1
zgzqRbbBrc2ggtGvnvdC1HHWcQvtlpLFUviCILwGqICjeiIHbfpS0VmLTiLXCn0UTGYnS4Ao1/H2
6TbnqmLkNQtcUQ1sLSgdrA7mwpa+xLSKlB+mBZDTePTaUExE7I1Ae+Fe+Srihl3Iv8PQkxjuhNj5
0lxIb5hZDJEPg+Kvvo4yo86EeDrj+f7R9pE7VFTu4cfa2nRuZrRiEVwpuK6hnt2XTOoKeoJ/VelQ
P10e2XyvoymtN14o6GOWRBEDQ2ZeSWhygn23Hdo4BfPt/ENpm4CQUlyPr06frgbm7RB75ZIQ8r1/
GtABFAke2ICyVSdF9SfObcir7hZRVaRIVof7PKKe/V4UVTfRNZhzbRZs4FLd+5R2RnPT+1U5lRcl
d5CohyXUSnH+/O6F1CO1fZwwAxZPiOp3kFEN2YF4SRkUXx4CeI5L73s8kU08ZTLfVQyq64S4LUP9
kqj2vU9XndJdXjqA6lLWBHWnBsLKIERp6F4kQzfFk9gnCu5r0hZq4N01EoncOf6snirkiRMbcST8
gv16VQ+6Bf6idilMP6GCqCoVnjAQ7bhHWKNQKzP2lmkXS3a7ZdUhbKT0stZbe3yc1x0JI8PPVPXm
aBMyfGhIICJ1eoI1wVddSEmZTOYzSTGYjJ02dnsJmfMrWi7pBNVsPvJSMaGLKGGT5dbdC44tZ6rp
mh7WwzrnwwBgfii8+BomBoWInWHvfkB/a5qCr1EdnIvOGDvOVeBSAImn44dii2jPec2fBYqc0vcf
ZRmfyciNesy+5yncoWTACK2TNiPT45AABkUL6gCzhx9S0ZwHkXo3Kcz4uYyjz1GHAMTp4LZgzzoM
mfHRRWYRk79NTi8Eh7MDtUvx7XRADhK60J5vOpV25jBOsYKXTBF+LX1kF8T4VVw3zlrBoivE3GB7
FEH5+2VBnJ5JHeWA0v+zNZOt4M+SmIvEwUowYSa2Mth7aTxSFM7/oyMqWK6SqbDhp5OE64FcmInv
2/dNnBfHG85lfXDCegfC9pwsIPtNs0Np0ZpZIkxeu5MvQXjOcDDwGvsyiNiFcfdBTtjASZ9OrSHy
E7ma/rF30Ee3St68zlp+ZdswT4OMnfNQSHSRpFPVRML28JJLJ9S0aO3d7GUM72k6/kmMDGM1hLK+
8ZE8dbvpWS2wZ+GAo6xDLl2MKAmwBf8EPytX9wnShr4zNEUXDsh0Erw/acIwZ0ZGQGQ/YBTZji6L
hBG+tfAG6fhbWGCqcV8+tewL+b18VgyIx24ac5lHPs6bQEnKjwwe9EcCyAd/mQ2zYqz8+eKsOTkF
xceLvzM8KywsrpcfeTJHBY2SZ3TusPlEgWyOq4yTpSbz7WN2ChoQoHPNRRj7ejY10UAA/Bd5OkTY
FBA6pvSF0zYg5zEDPnosmOem3w3by4QIEnqbcP3FTNFgBCT6DwK6CF6e3edit0rkM9W987Qyx0aB
e6i3BMy80tB+3Y1PiYSTvOOd7RXHMaCoiYBInkZSiVU4bftiFHoGLyBHeqZ0wWxi5y6Llr3fwuWd
w794UsGIiLlpbc1GxknETkKDYioRsbKKwa906E/3XMFEkWA5J4Filz9y2CjKJBypI7Byk+QnmWwQ
t21nsONfb1O9yndVEysju7X+/MiZk9lntv+ug+/NhZNLZclkv0RYIBfa3CCUC/aHGgJ0ILixO7AH
/8KC39mW8UdyRpy1gtkf4HnoDFMneimwFe1U0TXpezgVFyn39k8rOPcaoBcD1EdbbyvOPW6Td/s0
maff5uhq1s9bDZkJLV7YASogNLAI9i4Ky4QqnZVb93tMezGU2ePunD2oud3Dhz/gLDvK6eIfwmJp
H0sxHXBPxidc6vV4y7rMqQMkflEHIdm0ql+x35XaHfu288nvAf3+So4Bm/LtQvJkTkuo/+tEa++2
t/F/iu656Mxj8oxo9Ms7aZ1SGZotDdl1/sButuXnv8+xg7xxBlBQjMxgSXAROpvco3cgROqaW81o
etG6ZFs3s+oqiGC/h2N/J2MWQSIfUm/VVyQri7JvqJlq1/8d8MnoJ1N+cjiMk8FaELLrac8ZJj1T
RTM0QinQ1qmMNDQdxFBDsmvpi3o2rIHyS12U9mhQXlxLcncTdo8YmuzZENF068OEwS8xiDFNxK+U
MbKZDYlC/c4BItdVXqURPZ9uaa30/VPeaAY2IrnCnxrwnpSfoRLms8pcyELZX3D0GiE1H2vw6A+l
sdxoCbtXKOAiDdlBFo3226P7Rk1T2eVtaG07v/JfL6Qcn3/SUw/aS+cBQkG8BFgpO+2+aOot4AGB
mqLoGx6pOfYIf8xQSpiAdLyU3do+QY3L8vvC9yCZWQ+aA7onqQBg+ldna5PAZL9ZO+ZZuGruu94l
zOC8rNSUUnkk3JjaZ4c1U4FefZDzNLP839nplULEMdv+ElZbN9E4BI2wwUJPjiu/AjgGgEsJ9+Pc
iy/0jTaRV9PUBqPdUmoaWGttdB66rIx3BANXmvK2E+hH/6ogfbKfbn0o46X9ZYqi+LY7f/X/+VE4
Kxwq+cFO2wVrxuU6Dj+gAZyw/Ivl/EtUseMmpjX5H5kXQV741/SpbX7+S+0Kd/lPcGqS0Nq5EsQJ
tZskEDW0WOd615iSn29xxjXyGYumAZFLWsA4EbU2gOSn7r5SXC4EH0wKIddwf/TuNxvmRY+DpZ2t
ZNGtzpmwW8qnaJo+7GNjkgZ0pep15qBWKcZyQN3jNnk3Fq6Ziy2c8qskAK7tDr77oQeauket32B8
+0tYeVmpBX3quJFsnsCiNDNnWqMWH6SkBJHPh8ldNAeJVilE8OH3ds2wWLtmo15lIWCwByJKLtUg
rz8lvJypGGYwW0gKx4a3e8oPvV4GjyS9mTaO6BEtuCndoN7smPAdy3mWRqS9zTn4EEZ/eMvp58/3
qP2Oq1Iys708YNCw1gAc00ijeqFq6SYtXEMRCB2BvXl/K3oTIDFrqkW7APwTjq8JcCqLT1N52OhR
77Dl1hPmI20yR39DDlRXhQV5vy1VeqIO4rXQwWoR2RRzfD2E6sbqnmchmCkkEvOn2eNuPBd9kDbo
tSISrHeNsds1cx7AE843RHp0p3JmFLdcslE0FxXJBTsSF9OCeBkZ2dkci1vM/cUNqS5HGv9KUkLo
6F2QMRkAYt09TzOwe4HhkL3SpLFvRowIfRquXhL9WinaIad0xFdmVGfRlg8Q4EXjQgt93U+OXpke
/jr8uN1DcBe4//I3MNZVUV96Q2tcRQRo1c01zKQumDXMLxixqZAaJVTDsPFpKjS8iJwX8AblPPAL
PYBDorkC95ZivyQjbLbhZzGVziadJJfpVwclKAsySPXAdu6ebogjds/+EMPtlbXo29rANEoGINvB
gADIzI8Gx0ps9Fo/ulzIENFG0T9yEJofIXG4ckm+GIRMjy+cS+YTnj2zazmTNwYSO9tsIOZUuMfA
YgzkjcmPOtvI/YV4A0ilwmXt+R1/ib/uIWQnnFo7A+fmuRgfDfW9t6pdNQ+5xe+3cyXjsaZy1+v+
udrOLpdlMUC08vF+tO9GqxHk85fesQbvhZ3d6SKpq9ok/1Gy3AVKO3zVRgz/inGoPNOuxFXqdJGC
GE/cTh6fr1j8VKeS+evyGPb0FaL7fqG1Lbyyf+uazxOLWyRgWLf7IXGXHgvKOV8hhgC/PRQP7Vn/
dPS6SbjvWesI0k8QqUlyan9QZPXajJvPMNQYNyusWvnySvLM+u79U2o3poS+0U1p71FFd+Zm+Bub
A/f0tOSPXlle2/Gdz9lwYy2uNtmIsJteMMSUe6C4BbSg62atv1FI/LziV+OIE+MeWGwrtW/l85KV
WSDJSJtUoPRElOj3PihUnsibDXSjOacSGLPq1OcHY2prRd1z1IeNO78CNn68srAmYYZk5NLQn0dy
H/MqqdJ1V/PlYY14NhCe2iIblrtjb4ybddvmn9i7Qh80VgTKa25xVCQPvKVgJRNnyyMjPzgWI94w
n/Wy1m5xQnEaLGo7cNnPmwEt7YlASdrAr1SyehIi4aMq8r2d1/AoV02DEMGg+D8eUYpGcVqJX4iM
5ZT9IzW7tgszmg2+ap3mB8Zw+Aja4TRnIuxq8LUibvYMyXdqMwruydKDFr0C+69C8cu+yYYAlSYF
z6U8m1DdaxAX9rwS4g5XbmLS/rywfRS8oeganmAgwFQo4kD7NU+s9lThclz4ZrrR5uI7j05hLRgs
p6g/ByeLLF1NdjDyzrsPZZvFYCebdaUGG/OBR/8VT2vz35HlNWumqm0wfJxPhCjwCJIutimt7Mhg
K7u+p+hbt+RF4x0b33scx4UDKs3q4rDXkK+buNynKINVKq9lBclnYKO/gFkj73lQsToDRLY2T3Qc
WxeP8QF36saYOyoUnx2k0YtNwyzqpH+I7raWbUpoLZXN6nQ3CyUi64aCrOOv9O18FyZM1PtBqh/j
w7g+yxYBXFyhUaAZ2r2exWlfWjAb/ePmYOOd3RAqIvzzLQp2byD2uKkWavhsv7Z5vdLQ6BHEJbpk
xgVJPudGQx3MqDTa1pnneePGsLd50fXkfCrU0Q79Bgw1AptPlcsHLzAykw3DlZIXuyYtV7TawW0k
mXE1AgJdaghZBidZsj+3Sim+n1sjpgty7YE5fCXCNdPrT/+LaTm3L2aufjJwZLBiWs8NMAKl6duk
bcg5CFPdC4seurvcV6rkQOt6odmXqco0GRrLRjOGL13gwJaPYC+Ymf5U1fmh7B/fNjT9AyBYk/de
F6+6+AjS26JhhCNCIuq/jpMt5oK+WaAY6+ZEjRsXxjZ+ENBTUuJp9MklHA5BZ9+V0Y2mJ0wpGkz9
ER3s5MQ2o8NSJoku5vLtmN/7IRAZILv1MVWhNrLJVWjnLp8NV772vI4zMtkb/X0no5D5RmX12Iol
JErS4VA+Dz80pDKZV0HN9c0BmCATvbLmzrUEsBiQQf+Y8coWMbNOyKCWQ9+hbHc0e76vLrmQbki2
6Uk5U6eLADNuZMkaYdUdCNZTfevLEpM3gMr8OpfQUFhYozWi7Px6sONO4bfZbHMXont6Im1PoUDX
+zYmfW91e76sQtI3x//pb5zvmBAnmvrCyef1VDJEvsnkB/caQ7vsk2273PRh99diHnhJqL4DDW67
liWf7pctODovoSBz/dP5mocpt4Czk+7XYWnK02F1GJav20sgaS/5EBNkJ6Cf7Y0+BUKbd9SHbrs3
RncRbZRNYiEkueaVSrjtrTqycAskBJWiU8tfALAaCtFNVnY5fewqxfbrZs7Zb8pk6XBYXk5jtA+I
BkU1AMUjq/5LO+prynyERDCEdtQd7t21lVTCt5FPWT+AHYkpcOGWhFyHLfjkehtzuuMrVClsH5ne
ugNZCAI53/cPIyEeNQqTGyXEDJuo5KUFXsjtzKTGS125NfyiQr8m4SXx4Ia9c3n0+mSxXj6wzc9D
nj+wKfzdeguasJDqK9nmQgeE3KZT3c5WOjhrEJzUCCfYOqbrYjRRBl+eXFrGn+4DibNDn5s0y5D8
SAP8M4bUAKjc4tbFo692nfP8hfWKyhraAIrCcpz4xp9fqC5r8m1eVxekS/ucwWuxpPMdlFlKvJ2r
jjAoLgyYkrxDb7tBWbzIT2vvq14E1zgS9BTa6xeQ0GN2wA1Y8d9RjJbgLCcSoXRbyVm5Ek1LoGuV
lPAfnkGbXWx0EgIjA5k9CEjGbSOFxXOrquASB1PwRMwEznjkWaNqL2WfuXEZ9TFQ1CQnMKjOn1Bv
U9AAf4OaJVR8izaM6josnkqdu99yHpYudhZ67EOlMJcTVXFi1IUgJx2CL/Q66sK34XO6K+9y3pzG
DnhpGpJGleP3YZskS4aQwrtQKnvpuuwo1a2d3Cq4cjjBWeLAJ0ej6P87rAkhAVNRI7vXVoH3uiWJ
qlg/3fTwKuhOIlyVx8XdV9rqv71t5FxTeZpKW5SdsuhPE3+sYMaDuEHw3xm1od8BRBOVAlFAa4Y/
DpOFMyWLPa+grC8oGn3yu78D4qscPK9grKsKVc40FUXTOrm2EkhiXtHwsIonwtABnjq3c7zPwlxZ
WR9LKMwl5nL30DBEAYvLQAgH+0YvwIFVC3IkmRxBVeGWnMoHwDE7M0b2EW/+jmrB9Be8v1o/0fo6
TPZI+hZzLOMhq+VzvSkPA9vieJmWDsG8rIDdoO3iDBcZeYGaZ2TWJrrD13XwL+mSQRBZnwvjS1w8
Wu6EZXD9d6tR2HgpwmbEVOuXL9DYf3wIcSMAr7ujs7dbX1T4hbRMRSrAIbx57wDQjeMz2SGBSZRp
jgxtBDSP1uTEMb8dDCTbRwrTylf84vGoI8zu913u4nQdtG6TN5s9+g3zTxJgt1um0cmNsHtDotl9
kf4WOEySQ1TLmWP92oqL0zF6xKwaCgHM9GC1Xo68ua2Db44zX7nZtltpBspCwZ+jeMxtxsEKwHDK
SX+mn5hEhJnXgLuIiOjL7LdseF/QRrsgTh0Ox6gFR29lPBaWZxyVHd1x4cZbwck+SI+j9r4xhpdg
oPAXyTCYHY6FjVgyl4bYg8YWK7kGPPyjRXWSzC9tzbKeFuCJH8ZSRarU/X1JQ1FBm7BOGZhn/aYI
uyZeEcG7/B+kh6SdOl3JWJKt4WsrQ0iT8wtV6Mz1OQ+9/tOsYOyoKpeyzP2DsbMRCaVqUg8eh7kT
tewPMsQ/jo16bTZVH4gfbU8I0m1h4SlSn3uzyDk/72oVY4pm0RLMg8fGbYjhKEvdB7fQlTRB/xQH
oYdnge5Lj8obPHECe686H4Xrvi3vgrPUTiaz8k+3tvg7SNUp94ZIJQZ9Ne4NVzYlHSh3/cqgjjrG
ECvS63yZjXMKuK8w49DFj8qQjokGQefSiX5DqaKSvvSeQqNkE0Duyq0lkvie8QxBhED0Axk77UvY
jfLMkCye1P4MzinKyu2I2qztKSL2bEG8IZmpNBPwGexjz0lqEWJng/nTirnHIPB1ga3qVhDbZluK
FDeWyy+80db7Tg41w1JRCYYTZJ+cUJ+wkgP0XpZfUgPhhBWSTdl8uyy9gEqk8mNMSo34aSzTL44J
PUcq5gMUY/2jGgpDZP9ZIIDtQhi5yUpNCUsmu7aabudmRRT3uyr/Af6nxeaa6rd89fdGOOeiLgD2
NYYQimMhJcAuuLcH9n+pKqgP/I7yEfvEGMXej1dLwtu8nKTvTAZRkTTK7fJx/bEolphWkOTivqv2
TO9c9AquZYrwF01A5owakFVGjDYNp7jpTTZ3gZgpPmv9CCSCf3GdsrtT76KmhFirHC7NRoRTY2fw
OH5fzmJnlVKJrpv/Nr6r4ySihA92I4Ur1dtuLOG386vjB/e+QSVAAfY95pGyjWKvoEYk/o0JGW07
5rFRnlGdwC5tPnfwc4jXHpyu4q+Izok4toGlyJy7SuBIh+I5V5SnkLVEP1LdnarapO5U4KjmzY8E
ZYoxE7W/NzqkPSeFWS1T3vGhnDj5KIYhZg5oCMK8J5jMDAOVO/1qMrjwazrpQyDVZXoqFoZdkf+e
6rSMs53sKYDFWB8A366B/hwCyzjbfn/o7s0LcwXeFw57eIVMUgCi+RTu96WNLgv4kxAR400mbvf9
IrsaALdChkepiL1JNi+sDeewqAWdMtqD7UhbQ7FQLsY6eavhBGbVxmwO80VTB+bHNAuMuy+oMi/b
Kcze05ck6AitqyQP5E8C4sBMrn+GsOYati+NcREWEkCfTbUPCMwNYSy24WyF8BV1wgpBtoZXX8Le
1hOlWpod6WRTs0wiYpXbhSTTx+8oGvy6+wwFVgLNcbIcqXEZsa5c+cbDTlh5sV5wIexE0vyhpmLA
SkNFjaRYpAwDSnqeVYnxECw25HW9S8XhnOWT5tEi9Ac57QMi3KQ/bW2g5ygt2fHGCnjxsGJwGB43
inkVDifuZv3MVeMRfEIS857UfcxU0VYdccYQDHIJYrFfYjGRjlWZn+XgmiZGMl+iEH2yXPXzAseI
xC+b6y4IvlSBkvVKEp06AgS/JZtOKgUZUIUEf7zhkpzvWAEyEfn1XMw3fjnt4GUm1J4vctr9bi6n
0kVva/iU9xd2aEYv+8USxjxx4V7gTElXFKxTZqeCdeREWfs5rEAOs8tUNihEWXLADVWgYYaBdKTA
7zPWlLPs/AYMFnEjNr2yLKFdtsXjoMQ0d/l5cVZRIp9n0ZUmk8tTaN59UbUvDNl/35jVCWmboVAO
mdX3m+YO72lagaIRpKTDQSfHm+MFHpJNbXM0DVU/zg/Af55l8j2AkVQeATei4FIE16MSmyQbPEAW
6HHh2BMYDslurVoNyYlQumI1cBw/VjZSmKkgV8pxM6XkSvjdSKs9CvJEU30As8ZO4Cn8oi7DZwgV
mchPiUJAFyzwN96WSN5JnRSUyU+F+NAi3HguX0/g1TZaSbwIRg3QBIdHeFNVvuZC9JKoTnkzeSZV
ksKMvCEiiUiznEo3dsv+5YSCprwKlxVv9cFXmbRmBCuspjiHnRHQp7qw6ZXx4Ma4msMDUpqvtH8w
rxluYgBiQk3FZ5BIpcDPc/M7WRl0r3szKhSIzNM6Hr6qfbquISAPBvgV9SDb93IgeUMbalru6fWi
Z0vU1eEusx68r4rrvAno6q2dXATPkOFdSP1gAkPEfyEeVfHIk47FE1LNFIurZFZq4x7leC3bBbRS
FRv5T30gZ3AiLoWKPy/M9psxvPy5FtaApMmtOvrOaw6HepicZCZG/qu40AksI7ADl1ln4TWI6Tx1
1F2/OAhVyDkDcAPHFnspdJdMjXGqes0X3vmIhR6yhjVk+wnmNDPKkvymg7Kqa8XwfWXrzSJwaEnl
5XxmZjYZGwo4aEUXhpVxgL0gcbu1AdkAF5Z/goI7i4R5jNRt+LsV57uBzrCcK9Le8gXm0Brj2jRw
gE//o+Hsb2TVDzeqOxYcD+rb3laKWRVk82sD3Zo/p0FCnTK8u6Gc3gwxL0aG2zm/igqBUL+vg9xP
OE/mhVDnjOikbs9o7+SUc7HMrgfVbf41U7WpDZh7KLNpWPocgjCkcJFeaGZKm5SIphC5H40nYDU4
9yoYNuNQ0AztLOMGFC8vRh46PGWzaKbGupeMSf8SI6yaA19oj3wVkaO81xlFizibLoCraAj+ajDy
77LMOVg/nsLm8KKD4w5r9k1W4a0Blohf1U9s+M0+9//MGjLbx6jOQJAgK1ARjxjD+9zkxxaBnQsc
/mLH7qwB836Hjms3e8vKx6UIMQ98YKcqYhDzfoi8ipiBz3XirCfl8TTlSyjaxNNt4FSL8F7tBIde
A3wKp8gD8Jx7+xkoo3mMmQTsxYaywh2M664uoOYeIuCe2Mf3XdHocMUVx49rzupP/xRtqndDXJr/
WbCZH5vWUEeIpwmvu4XfOYnz1LQpFtX1ThbOTjtzM7Re5qupvgcxksl2c6/ZOpln9EDHYnQWEWyN
F8Q2b+p0d5mVsMN74qTccc/UKdSTC0kwv3Sq5qAi9wodh/B9Lgy73M/0rkfbprSHAO/r8OtmJ+Fi
1oS+rrmSWtxzo6aShbJV7vp1Mmf2VZW/nVJ5ZOQK+HVEOHkbW5bF+vFOLRjPaGlODip2fP98e5QL
k7HCo8fvc06jyCWe9c7d51lr37CsYhkm2AopLWju/J59kzZtkTItCyn2sZchWqL2KBeWTZuNFfqw
QnUImqHiuVyeG7XpLLv4DZt7OFC0YH6nTS6NVEGtU8OJkPXPtovVcEgXlLxbq1janzNypk3If0QP
ntuoQyVpuNN4iABGJRY2u5AuaNczQQlC5zhWcKO/wadLDwXADk7oABkWmYIUl6lXyCfAETn+sXIW
PBYd4I9iok9DJYgTnF64CPeuYpfUHSDECg9ygNZHT5z9Y/A0wVTUaEqzemS11IuOdIDm16BX9P49
mjmEZ2JOwdO0i2GMmJ328vU82U/NRFJazqJAdtYK0UJr35bFppAxlMkoQdJHMeJDLSHVAdl1fbDT
miytLD0XdHyYkWLTx/IE0oN7XHXVjBTX6c4emsxuYRR9kmwbaVEfPHpuFfg3QNcGCCvS6vGCrsyR
JV+LX/gNcApsPTzVv5Vl4eTJVRvYyHucOCfdL980sGiwT4h5lGFhVPmZfs/jlbQFpH11P+Mqk59c
yA1Yc4ByKBHBhTpwEKo+0M4be+ujzIQeEhIEMFm9WRFAeOQ6/3djiDpDdyrj4/WT7KPw/OlEKPnL
tkpCIvUS6xPFOwwvqk7fiMlTtLC8LCxnnMefzkawCQcKt+jfqPMpe41/WSWM/qKGFG1B0X+PauW7
68dFZ4E6K34Wq2HQWnm0zDEf9PX3CKfDsL6Cyg9c6DQxvFgjuSg19UOgKHco4P/NPt/zXOpenk/b
bHCFc81gEPlZov5hy0GMZpeE6oBae51ucFM4x4V1fq+/GpR0oyiOh9nSDhxrUluMXcvv/5dZg8Nw
Ntsq/f2iG2Z6LCzy/slVVvU116nunsF/dHtWQ2sx+CtRZyr7wg25QBXqQzG6CteazUmS8gjAPbC4
0Yw1VLBNH5SCi1T99dm9WHtFh9+LiEIrYJinkYX/6cuLgiAaYrMOhqAm2M4V+I7SrO+uf4vxZge0
UQKdu+wo+WyUDDmPgQjGURkrFJgaJcKq1bUxUSqys/9uy/nfoLpB4jKk/aPYwcc5FmkpjFu5y7n5
MTK5JCs2NLGaUA6slD9zz/e/fqM78+yOIpKwse99f6Qy5aBFnspJs5jyrfRH04F+BxuOSwPAUFQo
G1sfAWJZDbKiST2ZK+WsOdt/TdWb3R4ihDjN77wcHEPC1dykdzZ7+pbMTqSRndqwRYZykgJvFT8+
g6UTIzj0mUsnQo36rfhUG7jSB1im8HsdLExW4PJ5PeIygikQBNXR5JQVo8Q7DXd+wA3ID3OQQEWA
q+nl0cY6X6AYcY51gXX9XH4l5J6smu3E3I3MTu+gaW/nMqWAtBYKs3HbBi+Y2NuPQI9Ow1t3pIkk
Z+iYdtf9KJpoVxnx2iaqZwzChyd4554d7Rg+OvsjUHnzgXZxDmK9uFNmjw1u+W3oOhxTfK0lhS96
p4MMM4Iorop1Dzjl5fOXujM8xfwhJyh6Tyz83Xt67+I9zxxJL/e60UbCwBYIeK8b9oiG8j6IULS7
APSZbxL1Mr1KTl09YT+YnYlmL533woiQhA0HLkQvMAj3nEqAn5NJ900yLvSJJvjU8FpAOKc8rhyY
c3Pv1xpJc6OnUn0oReiA7puwDvR07WMYBbrjn5+10rKQX8b4Sy/qodjJn75C3MVV5keLv17IoqKr
MLoqB7Q8t2Gz23KsOMlRAtkgXCeWKgYDpXRL5SxOgmud9GC6Wz8q6Fa/mMZd5KCJjKNZtCOxURXz
3w2ABK3sxBSYD+XhpUdzpDCpR/OhwbvemzwBaQL1lgLDDXL1rluulzw+fcoZxp5Chbgeqi18v85n
Uk2Gli5AkHfWpaEgd1pWKf6eY7GpcvI2HFztxLvTMhqWW46KWbMi61gSRgPsRauXWH4PUa3d8pYQ
HI9fW6jOozB1Tl0eCip4Oq02nA7+8q16aPdTc3tQhIFVRyOsRBHJrh2o9TnmlU+ZOA/5EfNysexQ
SsXH9QO4j8nCMWRwY1kkBNLMyQjLjYnVTrfLSy+C6CopXRv9oF+SJJb8DclPWAUs/zdYwHQXbM4C
G+SeabwcC+IPbK0cqk+B2S1zH4MPsjAUeoyeHSBI1iGa/A2pqUGM4Dxb/2VliHR0wbxJklcQ9gsc
Niv54EExvWo0/m4au5cnTxJWWle9iQP6teogprbBoqbDbIPgEkWpshuFH3HGXxpS1o/JAjmCifev
RXnR6lh6r0U5CX+lJ95wovtiMVNJy7w68KbSoMLWhJcLd5401cEHMy095sZFba4BGDWONKeANMr7
HOiwAwA96spmPL9sAF+pPhnKjTJ1kWGitMOJaGiExfwNP+KBuZPXUCTqgMxh5hPVniRKIb1+ooMN
VjcNu/kdC9SGhzaioMAt4q4a4/VJNvzmkZYe4ku1i2tECXBH8FAqPzMI0sLgl5Ql7Ah3d1XRG22h
PKdFmnk7Ga+VLxQfx9pDJFC26I6frOMWt1EdaZFEfsMUzRcKnhiEB0lhWxUKXqbVIg09BvC00XB1
MgTHNNzJbD7Uo0IMsNq8wm/npXzPWaWgcsViEHqTv2vXfkhG9LKAif6wGOIQqAysyeT5axviur+i
IZgfgYeXoXX4d/JDDMtRUE1G8APeKvjKiO05vh06iTo8/xxEDSFpU1SW50OEkEyt/t89w3QhEr6g
pPVig0Vc6AUdnzSZDmeDACrP0f/BLEVTvGAQhFAMgPhrLo63NW4juMI5jSdWPepKm1D1MpnTOWfa
FBLYdGJfl7tpi8X8UhzE3y9XmQPNGU0UFLqJBvXWjCkQ24gEWEJkb80CKUFBt5R2yAXe/JxsOhip
ewIGXAq+coQNL2idj/j38lR1JtXxknRYZf3jxlYn2ykXexj1MRdplufB5qbpnru1DVzymM+u9SWu
tTCy4rxIEOagaAs2Nt2BdqIUSu/BNAmaxPC7BeQ1DJqt+j65SW0BiPwyZ5rq8wMV+cL42vOVZ0d1
JmYxZcpnjmkzimRxS8HIl9VHC4NOSFCGKHq+9MbB6FNWmkWLvUuac+zgFsHSuEzHK56L/D29D09Z
lpuO8Y3IqA4OEcKM2p8W0BLjvdg2PxKJOPrFEZKh8ziCg3Nau+xJFO5++Tc70RFXhyB/GFjNfK8M
3i6L5s2oai6aXl6c+161lGxhI2wciHJpmU5AB/98X3OyBNCEi8tQCQ2p4RZByJFYdf8IXsFOKQ/J
2v/HlCbjyKWJjsameg1fTbXcnOt1cV46aGInXW+BYcO9JtbQBwJO5y8Hzl9bOCSktj1LJnh8k2G4
3zt1LWSGjzaOxFh3MSzkxxRVrlfJOSZPaA/VFQT6dmV5Q8wqrQj/MdnK+4ovxtwZZHKqADZE2oi5
4erQE/d0x/b4oG7XyxgvmTk9VX/4Y5rP3kXhR94fSb+f/tTXd3scsAt/fXZnPjnZ3gdVd+rnj4Sh
4QeHmFW5saZT4IRjs3cDfNodnhXaXLCPWR5XGjYyePRk3M3hdD3obF+XSCKzsI8MG2et9gYqO0Qv
T6sM0AnzIvjcj3aBIRi0xprfM+qqopZLFHmDDzbFX45IU5jt04IsELG9Yb7qP7DuieFUolbZGExJ
9Doh3FpgqJ009eIUw+0rrFJCSHsfyfbfGv3ahDZDUGWCfFPyKhTbv5+42TVGhjDY5cA1/rRlXt+9
MiRYUvq/gFxhRFGrZqNjlJCv6D6q0uzQFnlwCuBsDsFuutxodSkcn0zCZjLV+TuLQ7N/yOistrrD
BqFk8gNqO4AmeaflvIZDe+9zAjrVvGYLcHiPW9a2j4IH6W6sGwC1XM5rMVkv86z5gFCHocXc6Jra
JqVdE5YpEGfTestb3JWYgycZguYI2gFwOmdiIc2qIYhXbFNYXgyogxCj8BK2yjzM2itmUjukfgkq
d7OZUJ2/3oH8JgrOOilt4LqJzHwrnJBhknQIwzCcSMzGjb00WOS6MN5DMiOxFZSenauli+Tax2hd
nZhOvBhe6GkCKyRJTKmcklAb0SYcBqHLfa2OVvud9/mK/52KwHikKzbrHK6novEdTfwozOuMwfoN
dowqzjor7tD0UH8zZHjpjMLBDvvPG2TzNptN9Z+FvR/v1DoVqelkzdEMNmA+tB+IObaUOLlGOu5n
MdTIl/SdNDBUL6N9AF4zPR3pj8TkOR1N
`pragma protect end_protected
