// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YgL46umJxDiYUrCIrymQzsgmMI7f04JTaF/fqC11I54wIrgaPYhOOyFTIHorZ/+5
Iu8vY5iy0HgfKMEBHwCq/Y4yftnvwfRgnDqYFoUU9tNgWt6dcb2ZjD7ttZD13a87
gkIKQ4ZB2uTde+GJcGsJTJkmdqhiMnLjMFYkYqYNTTY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 49984)
4AeBwOXCNwzpjDaZh1A4yoUjHLnF5X9ie7lQqaBJR5EvlXV52QiwyjrRt+0FPkfY
hCln7ENV725xDcvJlT6rxZokPMF6ZBfwzHc4FzM4gcKV20ZS/q0aTFIGTaZ8vQSC
C6JJ1riWMI5+9nPuaM5n4lxTIPlVRvjDcSl7kQ+jhbBGh8m7PbE3vCIU5g0w4kUx
sO4UI7AUa9Bv4fEgYUiXxRDGdwRsJl4p6hfNcqh3rf9ziogWq2JbaJcteFq5QgXh
blZ5+4Z7w4qaonir4Z2P/LZcL/IE/2mdRN/a6ZJNF/pbLdDowGMQkbSxOoL+YsVg
0gAKZUeZuyipxrMp5alUS+GUYIE+aDXiKRN+SQSsHis0a6+IHMA60WH62Gej4bse
eRoxpqDWs/8ebPMJ/MHkPuWxQt+z3gcv7GI8mAfrPMp+j5/PQN7saqXsNs/9EmZZ
sjPesTWrNqHpR9OqN8ZiwXrV3SRnRVGf5npmu2eSZ9TgyBpxYOVkv0qiwb6eo4Wq
lX8P0tHfnA6O3MoMle2XOG801z0bgfwdDqU2hobrhWrHeeirAbZ74jZpC/YN+6I4
gJm7qjrYAzqJBMIytOKARxQNSdGcsMnMR53zlvt8Bnb13iybnGFtgARfIw+xWuQA
UqJCC1+afFo22Wn86XflfaCjRHB72YNk1keAHwWm0wEPBsoh8tif8Ss1gEYaf6U4
0Rpcx2C3ogxhFoADpMVq/vHI/Q7lDUUkN7VJ/QDJRx9GlBsABgu7TWZkEP5HOXiO
+o7UANwZA5vz6QGoqrFEowekvRLrqVvD6PyBSyxq91488KURdyOJ7X96+xgxI/+i
ZgEXBqdpTUlqFYEaPl+JQebsR/1K8LE/c6FpFKsL0q9OL3coAFyfQPbvLJ+dvCHw
7bcJiz64+M7jTMD36wP1maWhlGbIqb3DajkpTvFibe7OuCtKBubvDPfi8NZn46vY
dAWI8DWOlDwt9WFLq7E1gLCDolVTIA+YR18u7iRYw68YfZ6g95D9YS5Gx/IYtjuZ
dPJ69olz2cjFu/35rn5PKfErW8J41/P74KVz56Hvwzdt5oayJZkVW8+4P0TJfS8s
uaOIv009t6d3kkm76SdftyN0EY3BFDmFClW39g2EWProHxghBvRhUsRa2JjqYkyL
X4kCERSZYpkh+E7YzcYXIaOVoun/O5ezc7g30q74KpCS1pnE0sVrihuFR7gesfm0
o6Zpip2R2Y/hzADj012NMOYm2f8xljdhwK3aKNQ3IUXfImKBq/ODnZYD2/lcDwcz
pjiqNcPckn5Vr1QiRoeQyULGe47ZbbeXDNaUNfdkHnvz3UxI+UteHlSf/h+BBaXS
BGhapdboAnIn7VLSUfNb+HebkbRf8sKWMEwfNRJQBStFeK7PsyvItXZ3sleL45CN
AYy1m4eG1oYnMRemOW0ml/VsA4ijy9fFIcYh82hm5rxuR+OJhI8/B+22/JAV/cJA
uUMAuYpy6zO1h6K12KBNh2PRJOFuXESzbLmebLlWur+qyHsErxBHMtKd/h8E6TLB
rR/b6X/64loRG3qd1iQ9z40Inr5h35jAbw3NdhFpFhG0OJ4ZT9pbdTI0xSAs3/AA
d9B+IoBYpb44lpFdpfICpx6p8BtzMmYj4k2ugyvwO+0048+XOFR4ZV0lkbNo2Tkb
M6Hu8hpOT4cFo85F4BEsY+jTKCEqf3Fzoyy0DJZFb8SjpXgGKLqPFpmHhaKZWY7O
BtMbRGo433KrrxFpdgK6LYcLcdDVkvS/+T9OchgBo/P9qNKUhn3v8ZHbBs67wLS3
beMWktDRpkHcpQvC3o/9XbxKbM8CjecFSaCxFgg9d9F5mxC+7FUhoicH2f1iN3aN
d6qi2xXKhA9VoTSNcypbl1tcLSEEGII6HcTkpsdW0SomcDeOPNBkWnpwdIPLuuSj
cQeYVLgnxRH8hGJcIByuyzCKLn0IcHj0g4wkxjD/kc1IPpCQMa0ukKulUpBCn6Db
CQLKU9rODo2xbGXoDQQ1KFlJPXpC3E4RP9WlFWEqdvkg6nrPy2OQ3F6NmU6kM7bR
aM2N4U+aSAVO9B0sb6Y9LZdbr/z6EQhOPR5Tx5pEyvGivOk6D6DwYWgM5GU83cft
iAkebWPnwyjdInT8VMf3mNHWC0TODrUe3SSntuSYxiY/QykyDyGKuVt4vCoTDCzW
S2d3k2LWPR2O0+CShHufkzXs9hsR8RBhPcTymyaUNMAt8+4Iqid9JmzP6KY9FjN2
+iLcINovSLb1SWtKPN4bsAdk4XC49pVd+fRUu0Dg4HloNQC6yCadt6rmWYULZgGL
IkvxUupwKp5+z27eDPRZksQUdJreNih/6B/NncbY3/zS+4txR8vBzOZDQMZEqcfG
RUE4/3n4S0QVftTT60C5Cg5Pm3g51sB5pgvowLKdmsnd5H9/Jw18cR46YwZQBHWY
Z9f2vZYocHfvL6tXi9+qSrueBoW700KcSFhF1tBUezYebD7Sgk4pJYzUAwXqTj+W
l5NWtAhWgMV1UxWR0RX7+GumVzCSI7wjtlQZyDlX7Hx5UzJdXtOBc0XEp5e1aWL6
6BpTzkQK/KJ5GW/1gzba3K3l+ubLJen6WlMevkGhng3O+8auUIF/dVhSuLFRkYxL
Zo2bGu8a28n4RjkkdZnuvC7u6MfbgPZHXByTh+6GgWHCLHPylCUUKGpMopkkczqX
jV/pXz6863rD7DPZOjLYsf9ftCm7Nh38Zidw7kZkE313rFzM5l+dRWaTeTDsuHVk
L5058HZ1hikgekw4ErlAYkjhhakJ5seiPZb9aIIdWLhETNz2FpZjE7K8yR06FJWi
OK3rjFgaQec6VqRsO6YCtbMyy1sikTCYupyhkGM9IDa9n7J681xRWyv6tb1FbrtF
uqDDTlQBhpK0Qwta281kpoUdeZ5yHnN5zmXdY5e/EBcqQ1SD4/F+UDQGCjKbCxi/
cXvLnc8ljqsfPc2R1NLzLQJ1HYeGww62WR02IZfr+uOdCEvpE6H+6UJfszT0Dglj
Qn89tO3ihvVQ4vrFjjoDWE8r8Sr/zC/x6paULRk0wKu6E9VUh6xp+27HHc8FlKPt
sba835ZMsFc3WBFOBERXoFYyXtO6za/oMUzsOe844k+YkbU5tWRuOcBMqCIWVVrq
5J/taM9jl65PFGu/S1neUrIPY4gfqv4H/e7wZej/IyTFEafzV+VPh44AA5oNvwzv
GwMNJ7SNXgwq5lG2b5CPQvbvpZUxDg6KBWxlOf54eIgP4Lt3r/iiXv+q/w831ksf
x6xFchwyhFaaHw6v0ti08LCIicBF2gkOJeFTW3+nQBYcU9ukLInTytP5OKw9J1On
ngEZVwYat+G//C5z+b+HdX+mxlOOfP+SIN838/UZZu2Sn5BEQI8Uu0Ony5oh7OL4
VHpYuggfomgke8moov4PQscXOuNBrhVQ/ehXoCIlzaYW+6uPAuRw3InIesq0Fufx
C6UOSzetffslAV8/4BoUAgECfy58/3RCx/qaahAuuT50myU6DVpH+7TWIRxYyAhs
tXI2ZdjanILI17YE7UJdYZ/690YwJ5Edo9xZa2el+3qkrx6Nq9FZzfqBwgWF4oLp
8Cm0LMcCrTPYF6lWN9bPvDsTEuAosdzVAKMefc7dp0FTCbKDe7orCcW/p1X9nHNj
ilP0K/4ppqM74w4gGe1klWmyw8RLq3ywngzpYsLis1p99nwFDVfDsO3mcnSNDRah
OhJ+5V9xytjPXwDvdtfEMNUzgdikgIH+XkmGf5AoaEhxYfk6r1XwFmRk+S+ZWz3s
/o6hmPauAM6n4o1XYTa3YWu0BsFQAkxOjiEYO9CiuZDLt+XrMu//amKgQ9Ljqq9i
0C70bo1MMA3zlOlYSBU+O2qEApg74M5cTKdnCvoqA7gGpXnhpmaCCuLa9gX3/L8G
U6Y5W0oiNeRIvupQBc+9BNyIDVM2He/67c2ceQMfjv7TT4PygO7W6rz4CVf6MtIm
xahBvCPnOBalHgryDQgzAPk1hjmk0EctXAQUauvIk9H9IqQNAHOmaB4fCiiqhFtx
KDozjPaQeCouielBjnJSEXsBf5nxJwVI4xqJ+nFSUZUnoydnfscEIsemKwzYmxvG
BVcFzT7VQ4fZzyp0lQWT1UwTdML4q6Se+sbadH5ZgdSAShKzrWMBB+rOqxeJx+6A
ix2IZPDrC+krgyjnCT8aV/IA0K338goBf0xdSbGOoiO5kNhVH8PblItdaNfNHt1j
m55MX+VUHvDQPjRzt2YItoJEe6qv/Ddg2/0axWYf2K6wkrzDDB+czogMhHNs0vRE
LHDWUUr778qMw/AbdrKLS6DAUQQS94/rIeL7De+8w2MiHAjOaac2nSrEclfhZUa1
VEj3onFxU/KxE9BuVRrLP/gTekt9PQnYYRlcjxdk1uRlHFXk7xwNneWO3/37xWrA
j9HBnd2uwG4BYsiDqPoi/rTl1sYAePKPHlR4iT9oEll2/YfAWnw1FK4XjsExLJuY
4AfANmELny5ufVWGFl5sO9+2C/Fzl8biAsKLcvGttxtRypljwmssYqwvNyWD0b+m
eat+8u3Brtxd6/IhEM9qlPMln1jI/sDDPH5EyTIuT0Ff4BS3XVn1LGHso4B9VkXV
jKSejpRjC3iNZg6zpQz8qk2M1qQ+VNDXVeiKCuVgiHLpc17Nff6Ix1ms0nuyRTry
Qid7qiSsHaMbGP8Uwl9Q2rxCMccDer6VHDrkjUv5qJNmgQDlQnF6aSj4Gzt+qIa3
4TlPZUEcpO2SDzx+JgUulSuiicWe27WTJlYSztvL04pzbAWGwQzlBNZaTqGd7acR
1+SND3SkY15DvrLGjZN5yFD4IPDwPBHiDPZI1inunXoIGCdVJIteg/FvYjTqIQrN
EFgglilV5rc0boh3jZasokjBRME8LWpvR/3Ueu1nwOijZXRI38OBhY7vACGfWw2k
iMSfxgq3eyaYnR0Inwwc7eL14MWUrUFXM5vX4wy8D7RcdhQZPnXXbEDydzw8eRGA
fNZ/WoQOZ2ORqgWg9haoFZfmDMByffWOmqxJKlPg1ZAERdl3KWu9AJh221qRo3dO
ZqmlW3VjCaIV0d5ZPgG4VHHMYS8iiBxPdgu/og6eGVa7CGEfvJ5Rd/030qNt88tv
sfyAieTcvgtEymG0cltbWQCeQywRhCyVaVFE7pVip6g756Mgp4k6E6+K3ZcS8ve4
VO7Q27adPA3E1LVcbsXCJBnZ/3B4qEDh5dOTDCzSTgdueimpT9bP8HXBhD4kDOMS
VTs6y+Qq/OJChn9XBjYQItjChQFORYh9vIFXvQFBv7xbKLMKz1l3ra0Sk+f+UdzT
IGtq/qEr/0WEVRz3fSQAwEAjG2pypAjqC2EpLBb7K+1wU+PpBnkandpb5AkTYLLg
mRl41gEiBpZPST3BJxPXoDsZQ8l1RAGF75+ppmbkvmnoR7TYB8+yU4RqEBHEQ9RJ
yhZxJkMcmBXIlxPJXtE5e4HNeq27KU+uTIUk20BNsCJYMwrKz/apaSoe6vtW6O5b
XTiVgY0yiyxvuSGdY8ADxOSPXGuRpHDSAjeNnWRiMUNhlKmVa90uTg+NPJ+VZJKb
za/EJQSwRaw67rjvmuORqBAIfAQP9Y37Bjs00EgUgTxkucMxzZzbv2i/xJDGR8iJ
AjFpetp/e9ujbTh4BLusoJkqSyvNkdY83z7n2WuyaYPTca6gvzT+opHqx4wQSPKh
VcFnL1OcilZWNunOlKeiZq35sBXaOYrRbm2NAM91glQ1ReSyrQe6jKR2qpB6iE8k
3yR262GqB7YvxJvGYDUAWj1xq5WAidD+Vjggujv/cAloLsE500oCS1G89+BAH/xF
EXa6IZg0i2zgAmeQ3Qn/Ylg9lfl801EcN6N0JcfhY/+9FiKID3Dv9/di7e8eVMkk
yITeGx1ziKcT+NXabG3uemN9HM2CL+53nqf2yJ/zISzO9tcBM+tctA8IwOQNw8Af
HFaiMzTK/9xbtFc0NuFlJCUVGleojVSn326KrUaMtDGiKERxuu24WySrfrSGW0BH
yzMICgbZf+z5g4pJwezru4/VsDUi6WQ3iwPkF78888BOljWETuLz3vvfDrZjJriM
Tjqbpzb/Gg6lqyVS27rGgP7Jo/BrqxGk6IBZM+ai43tIKyxsi0tCgb/L9ya9Zm0/
EbxEcf1bzibP249j6/j5utVmkCUgRq/TZlEEf8atdKXf0qyR+MuS/DgDi3QsYQ/2
z2nuSF5kLyL8pJxqZfGE9nC7zd63AbShCxzRvsTtbQaT4wuXf9ktA8oc7rzwoHYJ
ViGci/Pb+ZhV3DDbrfQDo4N3bV5msaHR+fRaRBXZoWl9sZpKOnLdZLTgaBb9xP4N
djFEd7KhYPHdht0QVOdQdzUJHClQK4gnLMb1WDfcehqT8kJb2DpyoasTMAP0icJH
ZsoLvY+4ActR3s9EFZ7FTRk3Xvt52TIU70jFaOLcbvi2A+X/tqJfhVmMp3J19Vve
h9dECFwAGlRqzXXxwVuPub4q9ihMkpV4ZSXrLxHThLmZpnbdGOEwYoi6nsPrGCop
hunJHjgBuiNlAC+tdJDKU/jzSUtWrzqfNliWmUG2X0QvzoAGse1GOpRx29quH7ks
IqJAczgQrK5Ap3+B2fthJfiFR14Il5/wcFd7JXNc6EIwKegs9heHCd4vCufbWXyj
Yp4hRnseOQLxitBt3RT/g6d4UANj8tU5oLMFkbz8DX4qT6jI1Pp+LwPdRxSbsWns
6d7u1783fx1NU+6GGUukWTar8ClXqYcgq/oPzawNchBFY7t/3n3PbA+MwY0+yq9K
rvvEtJH7pG8G+ZUNFPq3/rYNnIYepJ7VpBBZg9nqwx9nSZCg+GDEfy6adBUS3YR7
5BGDG31oYWkKdOsynxjkUGY56u8owULYpQiucx8ZmwJey4Lzfo0iAaAT4T/Wv752
x8W7JRYHhuEAI/tPNMHwKVt9G1Sy0IK84Yy9lHtLxdZguSBnGi9U5dV4BPMHkUb/
Kl+PZXmyWOgM0Zpv1tNcGrwPmbQLEQQ1PuOniE/WRfJd6VHf9ezZ38adpD/4lFc1
fhbJJ5rj7ADqhOj0OgXaJtyUHlW+hlfLZ2Td2GveR6vCGObfXnufLuEx31Tp5fL2
gMQOrxczmk+yiNacxsDTyMIvg3JQjgKuct0vQamYzIwIU3bJ613sNbcVZM7G5UdR
UVud8IiyqIqtUrde4TC7kqOdQQPGcfvPTgcOWvfQn9e4dwH7Ne/KsGXxWjnuuK76
0dDiknm4tSMN6AkMeluPXhXYDwDCS30fO7CvRfYQb5NFoBsvxe3RoiBnPyCiwcvr
BWWjPwXVKCajHusYHQVT31NpwkPqzeVK7tPEaSvPfpQFCRTwtTvOCAgBmttXjjPO
3DofTwt12CxV9Ht0Hv4dZP4u+SQ4h0ZFvbNK5l4ZOkw4Pd+ANNr9ZnxdS3A0eUph
Y3q2xJORZN/RAL3XDU0CMs+ybXGzAGqfN6DeqTFtGadxtX6VPt23LHeupRnY7QYA
ofFDVPjIlF5uktPMsNu2vOW8gyRIfMgTXqfVpntontj51v40fCoz3vJhlz116f84
VY0fXG78Kw5t0bD/Vy1BkSv2PCZw9bsrfLJZ3rggyj6vDdXJ+HKhoaa2W7Tkahj2
Ze50m97JzzJzxEJ9tqpMC0Z+TtG43tgjgRqJ1Mm8Ii7KH93KmxBBQQpXmwkTxpRB
JLDUSQ/tynbW3BjpvgWGNhd9SWGOrIJr892qJ3kaeAjp/+cZZLQpMtm9QuX+P7nc
MEHAPTPPhOa6McN8etKwOMt6TBMNb9ydEOzonEgUigxhhXIXneeTpI1JcGIQJ9Gi
Jh/GqWH5Uqa4JgYWAGjlwdAL+xeMt+jJc9IqYPNJuwhuc+xQaKBR5WtmkImfMT36
kEule6ep4Vvo8bGiB7tkrt3QY+5tpRxpmh20A8iPlGA7YM5LWe0f6XeYXwsQukeF
UCw7a7WgLRHVcahtN/wInFpgxq+ygPpyQuq048OFi7UeHL3mOk/3IonUbU4wP6uO
VIVSJdfs/quRUXtOQIiSj6ZDI6vfCB9h1HvrBJj5cKSBixilcRDCe5nSmcOiFeQ0
4ouTsSTZk4CGwg/asERMTzJq6UIz3EOSjRnrhTYqylF6MLBL472J53qMAhgX2HT5
+s7NNoVOUvrTqcIW2phv5/i3V1wtSSsZiqWO8rMsPYi7qPeR8Fuuzz7Z0GoaXnwy
YrpGdFVzZgxBqcQC8EFafs77nw4ShKXoeQslaZMfNz6TYms+NlAf64tRhIPW+vsR
fF7SkUpR11C9767vVY6wOC//wXYKDY9c1q4+v0SUoAZn5US3uZU+d4x5kbpaxwNx
hcIjk4YuzzgUfK2I+LBdzUoz33BVXYgt8srPgUXun8EINqQU6tXgdEV1NztA/jX2
Wf/84vmMcxVs4gouUBX4WSs4buMKO9QSpZ13sKMJ80gQa0Tk/8OXhC808hquQNAs
MPncN1SeVpvxCdl43zOguiVTQBIrl1z0HDyKIYBvEiVj2XbostigHCgmjaiDLa2N
94n+AfgXuJnacobV9zw33wEkFavXePQQlh4Y6ZehRQVBh1A1d+3r/PeDc2QqViNN
0MADQgwByDV+RLDNFvGL2oEj/IIZiFKXzhBDJjz1hn5tLoexOHpSNBrNjLav9PhX
VPhUVJ7wLzXfl0eMrMMUTYUbhXL76y9Y1w1s0VFe2r4ft1Ho+LmRgo8oR0qPiPK6
Q4qzVcGcIVLLF/QVHvMyju3zzLlHNfe57tLp+ouhNWS33Vy6kpuKhxQyoOgcfKcN
agKSUuz3Poujr40R/IQMoAEK2EA4LqCI9Jt2SMN5YJF30/6MOe8orK/adQd2Adz/
jA1+q4aPxTlMMlTddqKqMyBvRqcNguqsD8V5e9EB9a1HjDTGtvDxGgcFUU+U6Lp2
aDmQJRILKLm83dDMp6fKr1TtqUZn6Lz1Z7PUgg2vs4nMBtCe8Z6RxJNr2Pe6HHOG
d5oz/rdqv5SlYSfv1M/IRSjnMBOa1A9dd8bwrEX2Fz/acTAlIl2pPuJxbymwku7K
QMHVCpAUdQ/cMWuvK5a7Boe44hhaAjJZukJESTdMYOqKfze8rb0dFZFhYj24Iv0/
PlHfRtD26oN/qmmZfdyAIBCeQBR/ABSL41DE1qe67nOp9fOtbTJjTNcKczWrJZoA
XC7BeG7vnQE7WzQQEMfd6HXTs7ozB2geSRbw5V96GXpcP5bFQ3U5eyNH5C+DOHIk
llwb0bC1gnUFK9RxFJZQyT8BKGDsO8mp3gDG0yiivUHMyNfle5QyiZk2RKhGNI5a
o2pUmgB1Ua6stE/fnBu/KUNiSGBY7tJhCcmd6V/cG9YotpTYwSYtXet49GJYe++c
DigWSkWDNZUQY6JmUbLsWN1TFVeQvqm/6CouJePFnk2zFrBhb8ACEOjIItHdB2UC
QbHuiR4mseenY+TZwe6yHW5y6qYuKg7+84AsSohUgN+O8F3tu/QwyXzgBCi7lByw
XUWptjgipQSuWIl1jyh2Z/7bUSE2dZY+3jP+kb+z+hJpo8zOWuxkVU5PIRNuOR0X
EXaauvJkIQhGcf7QuBmVa9M/9571II4PdhB8VvGs+Jqji1hsON568KooiFPmFFNA
JeGdS1Ft8xXFk0laV+TZGlaWDTrAKqOS4SoKYPdxcj+86xRt8iQOBUnwKTSyD+8M
iSWkVvkWDtl0mGqVsyubL3ViAuguvBMjYI8y8pYEWU39Us3F3tOS6+nplvRztl3C
Jx47LPn8wieimxHvI3FYW+A+XmAQVLX+pXBt/Rjve6C/F4YNlatmhwCu4lTGpqt2
kiKboisWZThtm+GNcAx1gLLmTOzUT0+q0Gt92rF5yn2buda35F2ot1nVoC6HQfZL
rESIwP5uAmBTNqU9/ARFIVr0MANqjnITma4kJGA0DwdZ8qQj/OAgGFUbGoAkNRBP
X+f5RRIHJHqJ4JDLvTTJa/448/tAWDqpmEJqTia7Y/rL2oGeZRPaS4OEgyP7sWWu
665xPZ6tiUkv8+/twQXMHH4HEO2MLFqXaxs2dcBQuIbRWxKWGe5HctPrxMlRNG/d
RtPl4zH2HWrOc+zb6oA67t7WNJJojHQNWwJm0YI5JLZ2/ndyZW0GjK8FqMMx/dUc
HFF+BnIr1oC/QSj7htuq3HaDybUlmmRHyfZgDWuJW8J1TeonoSM4o9OnSHWMwQlA
cbXWUD2xPCplqGqqKHBolGjPO7RPh9sbeFXpvEQvVIcnkuVXr91X/A45RjM9osmY
MkGcM15wZnwtyG7qjqXQxCK2qZFrZyY2qFPbChkMTvOqxy/yH6YsET+T2rx1qTl2
iu0xDKyEdM7jrn8IXE4ivEyC8kceFnZNSX6+03ITgJotFhtilXWLnpwobdfz356w
8o7WJPMougguhPJyVc31zAuMZhegjl9YaiHUJndruTQe1HvEndtF3ST4SnzBACWI
QXjPD+TU6E7uZzOrxnr+PBVC1FTNDkSaw9FwMc8JfvND11C79/aO4q4ztcci3c6p
zC+4cFxfDXySoAjUoc3TKV7nlvr3rCZUMyBiFM8SELM4sBl0enrzNqccgrh6UZeE
tOjEj/vRlEThyfgNoUwdWyBtyOZ7JTilqDPTO94GiNnGjnUtYKW76+8Br/LlqARI
r77/YochWFAfGXnLQ/moYl5KXHCE7yU7MXn0X2OjUTS9vkdocfrb/n7pzDAyisIB
eM+r/puBMaVSYYuTUAQn0fbzxlwp4Px1vCg+1OJbgTxZ8NDgqqGDL5MbhtghzdtB
tFLM30kd7rYnOrqnaDBgWbn+HTp+82/DBMGOV3kCuXmmJ7BcWCGOSBuz1hxPL64n
O33EggQ0kcUSOGIQ14CRWVTz7JriT9YygvdezcQyQ2F8FkI2MMQYxk1+vv6Ja2oR
CEE/X3n+rnpzkJq1Fz2He5pGd63bvhhpEMj51BVpaK5Plif8ZIurVeiiRknAeHpX
bfsUlpdj3EljlYf/dwh0ZbYNF4uAuVRw+PTaYChbfMX3NRMMl8FMTArf9J90qYaf
6onDwLdDX28S34VccgRKLwZ3c3iZgGl5NIFlfmuC1VupNbU+zC9BLIwI3Ta9Qpt0
KTs/xAaoNDP+PExLW2r7XYctwu0XBFIVIa89cKm/6xFrzmwCDSFsUBhwwvSa52CK
Tg6wnIPBAVI17DS1Z7QpefJORtVEYx5b/on8Gjh8fFcV7mhT1GC+JyuGCCUrvloE
jerDbOKuvgGgf1fvWginpvnu5ElfekLBhbBOzz43fOUaxDWVgPeU6p2dNlQDvb3E
HVnHxuOxvt1rujdd29tpGH1u/4XqybvC7g8YVp9x9au1CqK//wGzfLy2+hxGQOYY
3ctO7oMzgUq3S3LZDkcDRv0xcUYgZ/dEj1FC6k4er3ToZ+Hf5PBT+6lZnm6M9RdB
WTfuoLn2rLZJSy5zdhk3p9SlDJkMydW3E08EkEtf2sJZR8784B59nrS0dKCL1Gk7
RcZyOXDSRgOq8NgXNryhWJYGuuE1InR6MsPm5+Beusy1d59qoAIXgC+YHtWEMN0n
VkRw6eVe3F98qjC1CplvWCGefcxKxO/gezm8xLaxd5a69c2sTTLeGs8genWRUkD1
WjD8f2837eDbyuDzIJxNssocIoVmcQV15R7EfARkcV+VA+8fDmvCa+1S7RTGCIOp
LVYVWNn/PCCj6Ed9Kg7kbsK1QECg3jWJPAY/wQcQnU/ce0gm/5WyOrkbtYwUDWCb
snZxxbM9CXeLWyMQLmvf19YNhRgRbv2iwsD2yhSu/QYaftxVnzmL0Bx6CUbx5Zma
BVRhNxjqtMJntzowLYx9pEEJeQ5akxv38TEdvYDg0ygJNxWvIgOYD8kc8H8hSVtE
IRCrVviQ15soGRT/FX/EcJxlBAPDVW/+YYIEoHl69VxC3JluLlpVUP6UI+d7LVSS
Cd/ddm9TFDkcoRxkxRT0bMvumkFS4MrfnRt9F4HS/+r4PODg4Lj74EbqoiNDuilM
UaiaWqI2rKvV1SFSE0B9Wfa1qrSJQTrHjYhWxSWlxlSUCIm/MAM0nA9SDgZGGDWn
zJ5IG7I7u1XlspBNPrmtLrWVwRqXdJLzHTfBOyzltw3Gjv5Ac8RdJNqPqlLN9Una
HWII+IuwhBdJ3U/Rumll65KxU7+TKH2PayP0wN5QsKQlhidGYY62J4LRu4dffy6Q
0Y+fGgJWWrPWsovjM7QlSw9bGUziHHBssoYPYRDWYhiQVZGehg+/jrb+6KE9a8LX
DlJdghVo/EctLo+gRawV3QxCZkNfzCnC8BP/Ff8tAjesLYueNFNqanLBmR4kB2Kb
OfF7u/kZxhAQnBTcpRtPxz9thIz2b0hxLmLL9sjwnjkd50eBgm9RxsRgbNCn2L5C
dCKF9Q/5nQJ50WVKeSHrO+prsn1UQ4GKhJhr+yNu/SAGJKrjYjbFcO1JXUj4H4f7
ibHY+/aKDE2xViVOXmQYRGgZuVkjwTFcVbnU7wKTCT6Nd0NCy9/te3pw3KiG+4jQ
qIPVeKUMw8XN/BoqaspDh+LA99hkPxIPEPUM4QuooRfgxqwmD8lYggZ9v0KRQNaA
puPuRX1EJOszIngO/cujq9q4acK4+Aq9AIeiPYxjzMDy+pSaln84kGHR7+NZlciT
u/+VG8LPp1SvGs5KZ8p8rMf7PuhusWY/tL47a1MrT47iqICCQeiyKcCfsgJkImN6
GYfoyu2WiIZeoSXRUhhfQ7RDCUlTR9QCo+CFvHbLvhZy4cq0+22zqiSH2XufeYfs
8cN/4VW6rwspDSIyoe+eSOMPr8QmwRDx77NUzn/xkOLv5f2RmkJTN/MbA4SBMMgg
lcCXXxCsMrmrKhy3Tk8MaCsr+5kMpzWvTSe9s8XQVSV+7lE05kSUUHOAd6zM0+kX
0ObVKgV1Y69np1bRp/jZdF9cD8RB1eFaVdz9cASTmq07dFC9q2XPR1q39/pmcQk3
xpzlZV0m0psUjFsF+vVF9QLU2YQ2G9sFa1WUUgzsQMq2Qhs0sZ5D5pUpfKgaACV/
Btx+ZFZeFnayAz8qk5yG7C2fk45U7bEUaO+2MezisDRYa4dkVM8O5NFunnb14bDv
VK7cQow8ZxdUSosu21z+0nCeBb8Bbwx5jdglx2RM3jCozukrwFKprBJWpo8o7BGq
zsZovaLjEa8aioILV1q9ALN4Zs+f4fw+WE6jbGRiO5YxdEq0rae3THqbblJ94PBd
CS0Bp/rvRd7d4spzIvouRgRwYX+1lBiBFAGz7HJvd7jzKnlktdCQeJifvochn4h0
3BvoqlHpub7iqq47ogUFGvI0ddN60xn/4Zv9wjjW24soPqdoFaIg5QR8L1oN7lBQ
GiyWf2rIB+NzNHZZWO5iodILKQ4Za3pOsw+aUgi3KvDegPnHCNrzw8LoAz3trADx
WrPX7M76BI9UwdXQWR/ilcjVcrhARP7cwuNecB8oxlFNd4FYT6NsJcoBvi2/+KJ9
LIV0+7Wn70M6QVMcKYXoBEzHTZxqsi5zeBNzFN2Wc8AKhchKWKzKwpVTGI6Wc6hg
Z7rltCnGAwHhIK5lvaCUD7JsHpel6FlolGvmLJKBYyAclDFRTAji/UonJiCvEYCG
nFaNQQipboM/OaX3U375lRAXz2xD3IzepXo3bo2+cKFtlG4HTFvdio/Abyzgcx+u
ZMjWXC1mtM+laJocd1pusDRwe8eJNCfFlK08MpuW33bXeGzdHGOm/YuPal+sqpHT
g6qKBqRLB4Ja6H0T/skWzJgLF3aiZT0BCObLCcjlhRtvvILQjxSr+A904JBJGhPW
a3Aeod/Dg++YoBGSjapmLdjMlJN7GlXuNsb2VkW+iONgI+/TF6eg5fAY/A3exgdD
f1YUwdRsXhWz5lZ2Ekjf2iu1M4KQONqhwphumePehEPoAvDDA2UNKBkNPohrmxjI
sGs9TEAPQlAuOVymAVRT1kJ2aoJ4JmOVdl2J03KPJMouFWpXqcvJHxjkzHsn2/Ec
IVv2CjsAsPO5KtThc8YXPKVo2LYh0KVm/0kMk+ioazaePcBQEzJOrW1mJDB5Jg/o
trHFZTQkkKnkscue6cnF3O6lgrKr0K5GT4N35hPlV72lwxq61S/c11ZYa4QPMOSG
UmuT9aZqOIk6Y54WgxN/FwkhIDEAS2sNY7+EuAEQJ7HOLseb6GUQEboITAq/6y72
FYmxuBVkmTcBi6HrCTw1CXIZVxKWhGdYHGpG4vuTOb7NmqiFjXjnkoSgqDeOfsp4
YWnkRUKn0j4iDFAO7A2TKiE3THDdRNRDbaab6WJzX15gYpcTbVbz4SxhjZpNVg+I
oXGAqHkdhTRFh6eqFcv8TRzNlysEu+w5hmUxoGFyZ21eMDbnBQSNzVf8MIRvo8o1
obegK/NP4NwKyCpQ8kX1AGd1Rfxv6hy7nPy4QFyV5GcXK/aEoGiTgsqgyRdVY/zs
R1Jpe+17MOpqHayFmZNWP3dOzEb6D4vsdoNW4Vtew1x0yYTs1cbe/q2l4+LFyoKT
t3rB4Nk1bdAusA19KyU0qNLSx6MmRod9VZlYemFHhHRxHZOo4Z1QeLivV0lrQCjb
zCQDCGZa1xtQdrckVMh7qySXtahHfAetCdrh7pxALA76NPGzv9lBHE96q6frPYnT
Lrgp203PGQ2T6sGbfNSW0p4e6IhBCSnnZbI3KzHcxKhF2Rsc6+w5ENGaXVmG32R2
A93nijOaEeZcDg/tHvNTN4DyrkgjV/b/GIMsnRfkc/VgAJy+0JHRyt32J1DIL2tW
SdaS7CxLzASHoMcMqfQEIWV1L17dn0MsY3enigNLFSFmDGfzHruZKw4symunbIWP
CQwjpH2ggyKne6qBYxo79MnyN9QfW2iVfeUsmxFtTz0gdVyL5M5tK78l2qgfUbxE
wdjUcfa6i075eUeFGAX7L0yM4cHk3EKp6t65XeneBYYVwgZhOWWt/LYtpJmcD6Ai
jJXmOcWb/eP+PUZhTu/onz7nRYCwDp/AWMPzVXh/ErlG6NBvUEb+7qyd0en5m/gl
HFb7fTHPTyojEFbskWE6HmxpVMgEH9g8foyT+O1P1IWNp2BbOlWne/QwAUqjXO/j
2hou8nZqpuFCC0/ftuQNdoc08OIPhKm3j6EH2get01pv4rec0BnyAB5LRq9bjyl6
n+sQX+Ef9jm2WdvGHpNrTfbeKG1/o1pybvQH+gjYP2UirAjKsjshTxI6QmXqVicL
riOLwFNwaxdnKosAk2QT0VDx4CamvPRsTZ4cmcKdlWJc/wDqlKK7zr0/oD1KkJtc
xoUmeJ3ROcu5Ipkz1qUJfiMRYH8vFj4Qri3NrZQQRN15/FlRoJsNIsUJVpWaD/X6
Cup3ypT/xKfQT5p9k4fqTZeO6XPWK8y0WG4AYA6jlBQRa2476ANBaeK0oFa+u/SS
s5yo19/794DfFHFU3vCWgaS66rLx7DO+7REqyuHlQX+DUYKRJ00f+cAjj1gvxpMr
PM94ZDqI3FrKsPqGMNN6AcHcQgOw6yYLzZrPk0UaxRLld9dFNbqGw7Pgt0vGX8FY
0BUw8UKwnn04rBHHXDzbIMoY3GtyXKD3FnmgaUrIU8UipunVZjX/DPECu5w/fiv5
W+4ENy6I+bn1YZ1oayoS+Uaq2rEwgc0+gJrIzpRMv+3Qrm4yotZPL145J4eRRq2Y
m9wfa7A7cMW/sNoFJNfWJhQPvZ60aCZKlyiIehUYyYd0VGYzMwHmaIX/7wY+hyvV
z4jrFyfyupb+mQP7vbLznm6XUW5BTC+xVYmMJ4vU/hxel8Wa/mC4aLoTXMyReMSE
gw4QWkRGRzzs9NoTtGw8VN2vuAd0s5WbeuTjP9iIOYnzSk3xfJuQN0a6CVgvPPhg
IpS3OykkkkQq2cTrE+XL8fbAujWNOIJFLWt5YtBOicvvcKMETWxLGv99fNrxwm5J
5IKxfkaq2NLpJ1YwDAzecL5ftnT5N8rpFNFpgLF1mgGVUg/fHo/tMRZsE/nEQWyL
0lL8WpVkLsAr2/ecsvWQIu37qo0lqjNCbXQmjr4rTgcohEmCQ3ZiASxNt70mAapi
UdHqIUUxCFNBjZjIJcACdhCWTkCTD/rcv4Od3/KmGUpHXb778MCnI7NqCX7kP9/K
QvPDjQwRi+OrJ1Cmy8nBtV7bxqMQDDTnrjUmrV8uddkuocpNdWuVyRMxGPusPali
sCKre2Nd+16Msp6XOgqDcU6zLZ9fdRLLu8cLbUx9nz3fCtAZjP6Dzx1A3Nv9jzRW
3jpLvkj1DwpyOqOStojbvM8EB0CMN55/xzOLCRPKWFZcwtGZj/iZoyNC30Rlkt4s
82GSi58/jzsV3TfWXFfNIsPDe1d4KrpOSO4IB7Z5YsdTxti7tMLlUoFA8krrVUv0
5z6lIErh9mLMIvZz2F09F8VSpKMK5BLsoYKoS63oTJeKE4us+SvdZ4tcNKijeLDd
cVjcnk0wtwpED6BYqeZL57REDcYMvhDPi1VRcAqB544kcD5vkYYuIQqJPGQT/px2
pe7iwV4t6t+5p+htK0oTKGFdrhvSAbW+7p1ZxYpPC/8zjUiEKxP9RVOUeVqeDOWk
NJP0fiasz/jxrSPjwS6IAiEG+pEO+398XOM8VpcO1Lou0+uN+P88tVTAGErf3RxN
MrwDu6dJ8UJWuW5gAA6oNj9o0pqpkrcGWIOQfy5vvpg58VYj/9b03uZ9FTivlqn9
haoLdqnlN55Df8XZPWSCmkj9UIZsQu+lk8hA0as7QvrqL+V8fJ2WXA5Kh/Qm8EkX
Rb1Kh8UN9BUWGhsQOdaiL0gLeennLd+EXWvlAAZ1Am9jGcGhuhOi4UGofMXmZX8V
Z/wBzFhLOxSwp/8mT79VKeL6bypR4DiE81+gknc7+yq3ny3hlyBOj/S8Z4FYdu/3
8UncCcO5bGrHg68HBE4BgEjOmqt4/KspXZbEp6AY3SjTwzmWwuv+JaUARty0e4Md
3UD3msmNAyAizIaUoJi0C3Qna2Y6+A9HhE3LpNDWJThmz4CHI5zlXL6sYljD2A5F
5owfxPk3u/DMc4ku8jNgCLii9ohBOJzWH0wrCWWRxBeu2nfHdL2CQ7E6kitMOg+a
i4ziC2XtlM/JSUghM3YdrWOcDHfT15FxcCns1qtyfLD2fPfR6n8VQWWqOGIgRw7n
EFx/SXXIo1JUKkmN5Cl4gNWIZxKQ+m9e5D9sESEVUiYrc+oWXcHLo3ScmhQe0yL7
rm/SecVQxdWO7Mln9pwK7Om9zWMSxXdW4FeGcKtjqt1NLC7YzwVEtSj115bVjmOQ
QHqAmi7ljam68JAJvd5YOrJoEacqg7YQjlhe6RfK7z0Riy2WCXEtgxV1/bcELvSm
arnUDa12QoqNCycata9seeZVa813P13knKApbzFQDM4iBsPuTOYdQXOsPJtyz3zc
qSet4K75O4X5L+ic3BYtfdBrrIeJ7TUwEaXW0p8ID8xDqZe/1EEV3I7LlH/0n3j/
XzHuEQMk/9uAzuhEuiK4Z3LhJGdvqmaXfffqYnl2VyxkSRkwPIC8FqBIHdY/YvLU
pxVA1KHmKsveI396nCCgRGfBGcoToDH7KXZyq9R6QxRrOMYCRx2mnYkX2FBRYeYe
IPM1LI+yZORxEcd0MAx9wNYGJ9mk2aoiAaBe7e0D+DnH4RkP7TxAj/LczwWyKbBj
51wiPiurToj4htQuRdnjUva+rihhRj8pk9dCQeHLkrhB18wiau7LCynYL0sxjE0r
8a4RPH3qyiDi9syrEjnCAZCBr/Xn6uKJRXiwwcBpiUq8IC8nsc0R5Go/dv1iO8fh
JHrazuh+ahxoef+BjUr0JEeGchvRLPg2YGTGgggDdPqEPpmC9GvAgrGRmPzIfqoX
0R5phCZXLJ7TCrrbmwcH2DQqfzvM7bSvaRNHmBCTAa85umFiPm7ONFtO3NO+Z2f6
FxYA2SYsSVyHkpKbhAZjutp3yQdNQZqTOLcc5AfZnN4cSWi3erMWz5BcPUmwCa8M
A1iTzc97sPg5EO1ldeTgFxHpJ5u9QT3EEpFntj02APXXHp0ifkD+0cQk30BAnD56
SRtvcxaj9HBiEb4WBP42V1xmTJduoqsAgWb38EHQViiRmNU9/lT1P9oSj4xRG/4X
XGG2WT8/w7hBiSdrTO10yYVPWfNZ0rAF2ptSx5ZdY27UPDAW1MEUPvI4Ta+bPq9+
hW2V+3Q86wAmPhPD3BHvYBt+SdCOHJQEgJShG4wFnD2Fn0w1/WVOo6pVTawA+67d
E3eosDBN8xYfTXpmYCVuH1zVsWVc0j4G8z2ULKR5KQZTFF6VCI9XECQdbB/aYfFP
srhB0t9XKQetHr36WGpv37acYg4bjjCc/fxjlrQYG+9hImLopB7+fxiGdup3A5rR
96hkMIwfky1mo31n5T83CjyfKIHqRtt3pGS8MdUME5SeAxA7ShyVHe1ijBLEQSw2
q/mxrwEM9aTnj+EvYGrMxiwe5C+TA2zOB5vlaPZoYRn6f3R8mg9nnWnhx3rWqRGq
aJBOlb/qpioQzwgP9v2gYX63cfQLTzVgGOhxp9xK5/a4OKgfq2HAIv6nkB/dDVnR
7fM2I41ISnkG6mMMSOuV/GRYrrkKp1+6UbIZYCJ/oWS2Kt7A3cWy3Y3T/FnaDP9p
3gBF0w/KE7tqLGdH3nNjCTAIhAGORRWIajCsfmvM1awcINoQADAT7c2LgM8GxrQS
rqvYcKtWfWd6dnG+ZpDp+hsMLUUlj0oUd8A0wQLYwlf//Xql2Uzd2s5mtueaWW2V
PUERBwX1KRthgtmw10aaKdf3AwQkyOJ6MmYtH+A/TVb0fxk+fPaZnrDkLfyYPuV2
mG9e6ePmCmfv1BzkOq0u7ijQvGVnqiRkJixybzhhp3tO6ZOzsO5Xa8y5ogwsrwkb
rpMwpmVhosTtNvdyVHH6uYK5RsqrIdVo/J9hIlD4ySpJ1FDV2pCVup/s0VtvBxZO
vxugELHkdQL/repZFuq4fVvc+i12w/JMn+iJ5zh+OYjIJLVGcNvYHBrjB08qhJgA
BLQWAM1Zy8M/k0XIHHafwjiONEE+T4jvmRBzP0r6ny9lEyHNKCtVp31oMsJKNO6f
LnJnhwHQQdNWnfcmT+dnGkswuoYcYf2YK4Xhrzg9j8X1uqEoctADJIBtgb48MwYc
GgsZSMbUxv33k/Ze2PhcKsQPoWcMB5SEedYPHEyArWJVaXNblqol22qgI+el4f3b
mqN7aCrwauCPhc6wZBAc+RU2WHlF4pRWfuUrwJmNHwbODoSOpKrz/cXuQNZYDS9h
DunmpvDKykymjth/t/pHVokRd5u7Y4bmQH65tdjMef93ZjA3EWg/caUqLqkLV5TU
A6Mz002GeWt6atIdvc/+O0tJFoeilSaKRyLAHtBxLs47Ub6wK8I3uSgaT2MEX3e2
n5xfP2RE0NwmVa3fGvWTWz3a8qAsSkSObnH5zFOGK2+4AhEmLs40SWryuC92M5ot
DpxACkqlUIiJaT6S4eA7eVy580kjuW69gvnBE02+y3AVUrUz0wV040y26OtvufEp
mw+5PZVAdpDz58oeJNNoNgOCdGbWjE0gOKTv1xQFbusrShbxi0VwO95QoT71FW+u
nvJyh3TRJuv9dW8M8yiHX7cK7Ns5T3JTYAB328/iAhGJL5krx12mVOZisO16zI2/
UyCpfOj9+MWL22ZXqrVsIu+AaN/VTfu67z68KUcMaKCgsymdDWS4/uof1sZlYg0A
cz25bb8DOUKfPi/Q+eOoqMnClxRAzU0SgF19kmhI/6xtHN1Dn8MbjR3N29Na6jQk
nAfa/LNeinAr40lrWF6JQjgrWah1Kk6ZG3cteqyP0/Hvpht5p9TfOKCzh2iDRWOq
IEkyiVrO+yB9JjNZDv7x1Lh+d1c5s24PcYJLoqlzs8x3/dUOGXsJ/FAcjSf2dEW3
AN9/z5A1QVvR93pxHF65TGTFwULIYQcvtqDh5Dnd1vN+o9YSrRvbU/1w+BHOj9hR
5NBesMaw6gu7itExfCHOVBLVmnUmI1CxbEqHRFsOu8K6zUJNv5ddvDz2CukV7jcZ
GiskzcQBkEpl+jbo8Zge+SmwakRSf4kUycgO+35LLhprUy0H/5YigVTVLUH3lZgE
+/7szCTR+7vDvxxo+ruTlkt4A9Rx04F52LIYOlwBGfLfS9TBXPFQQ5giv5DxnAeu
P0H9NVb2aYffEV4IZsDxWL5zZhe0BLSeKZlNyEkQIGPLcCK7z9YT/IpwstGsnra+
h9uXmdQZP83FPGtlNNobfSdf0iUw+6XT5BMKBDoD+1XzSGrH62khqiSh3oiTyQjy
NORoeCroQWIbROTU/tLmQ88cpvpiL3aWKqLw112Qu92qiRUbO1ky8Fq7qt0l39GY
8q0JtB+Kvma1dXOHLx/J6R0zzxk2FM3BblLZb5UF9igBZgWPgmTZP3wv5fFJPWUP
ACvza2GrfwQTkb13vsY0MgUP08yVG142At1Yu7R1NqlTfYglhn3dD0mOwM8wWFX5
rNBwOyYYNwmILuQhFmgLkgL13tyrxKi2lAD6h4EQA1UfpHQWFePp8y1SEyKb50uE
kwl4whUXl5YpY7vttI8lMY/+HQLLZNoEtoQAFz0gypycAuZ+vfnNk1hfkfxu22kZ
inQNKOOy0dFYPOFERqx4qWEW1peuvfU/Uogx+Vwr3eFIxngmSV8ZKjaQrFaKPYUp
RpSLS/mwQTZDsTd0YoIoc7h1MBJB8yaNvewm7KDkHhk7NeCaWhrNV5TiIALGsPan
h4YU89QnvlnozDnlbNx0XiOMbfiWkBQNtPCLNIGz/oK8r98k2WqsEZiVxKKkowM1
lo4tsdOlBhDcwII7eo408XNGjgachyErGOniM5vOZ1U/Djp8nLjKpmJ5xZsoVfa4
pqtTWOxSV/QgRNTT4opGtKO+tT+i3GSb4gifMa/kZhu6bHO6bqW+U3xXu8kvd2cZ
b3eHKTU/LAVxLabxKnNHIs8t5lYXjHxCZmpX3DtCQd8rCWxwboTuKKqwY+qcxe4m
DwEj7UYvD9uXT6qb3RUdMBWRq70CHycGUCI8byzfS9lmWZP2NAao7O2BlzlH+eam
57iBcAqrKARtlvnSp7QjsDAbCaacTrtXImxjc1pTjkB0roIzzDzo3NrD5tUTWfQH
9tqSvvzGPjQb/V9FzAC7MfuHUGz7/P1GFvRv2iTGpGFkofiPpt2Ah+2kNwEieVVu
alOjFsW1CU7jXL/f9VYrnKmqWJtS/hhsddGYsvMPPSO3XFmSV4k5eaoLNlV6wQk3
SGKie8vcCk+frTiVycdIw2XDjwGOeWO/78//VF3WFeKzjmMmWWwCVxOHxZN/BbTw
ZaTemigrzpx38To2/o/B5+GUcircLyrCL0lZrXzIOKYDeKkCoQnyU8pi04DWUb14
YOR8or4sRBWxVQ8fQFJKdGo+CN56OSWPspfdZ67oCIU5mXbmej9GlW5yf6QmZMhZ
q/7wJCHx3cpGJBQ9QUs+f82NTGta49+HCILZqSUjnCHTVURjuApRkHYLk0/B1+43
VVJ881BiXDSdrIiEDFixQzyThhTqVkPhoE5zYeb9jqMh5zhJiIMO/c9sD6GNI5PO
CnrmhSDroU+OprzwJrWHcd5fJE4dOiacgeUjbx1o8rihIA0+g2TE6AzwHrbvN1xe
Ck6tydopN0aAAhDvWDVHCwWQmccyQ+G8Com40nH+/0ZNsmeF3n8s1pmIICnjPtpH
nMgCQLVHR5i9IERGSG7s393jnxjfp80pZvW5h9dvDfuSm6RxjpFsdnodTlOkbaI8
teTr7OIqcZeOwEqoxdGleA88g2fr5pAoTgR4EqoMhbn9YGMCKvA1+BZTff1gFFDn
SVpIXoa70VVXrwTdwLGLaDIGqbvHo4AY3qm6WGAkNS+2ZcHuN1cCyQLvgHwgaZep
oqTzs8K0NKgF/OcDoAoaboV4TpTXnl79tlRtKfB6qcVETyIcmhAlOGaHZ0wLX3HG
N9gPAIW5d2IEve1Jdx3VJks0k1n4WbbMuDwhkQHPiTZVNCK5uufxJ0nZ97p3wuVQ
NzkmiqohQOHUYuDcAbitnsbN+Cmkd/L1bcCuu/jLGdWg0TQvRIfM/bbmZ6wtdwDY
UrG7uRP9aAWD7MI3AxwoHNf5z5WzsHRoHm+k152IUlFJWK+WJ/7HDoJGIJjWaNbt
0VfTSNT6NL376PtuNg7sR3iesVZuiNRJT6rc6J7Jb09PMkhPszkCRvE43Muvt1jc
jwjKuHQMgGu57nz8bGOGAl3n13aRQfdrj0bA8AxOpgmI3VL1i8xsNBzm2QzpSXGH
oy79usl99gOI00a1RggYgoe1sFUOOtCHftV7bMgC3b1HUoTl4PepPsMAzHXYARwJ
piMz4zePFlujfoeji8uUD92oI2wld7Kl8LSPqrJpE2mpcIb4fHZcDwU0axy+wvtS
i/SuO1dZiJGIncElIDz248iBFsqrbta1oR3MiH4cOxDXxGBZTPccJLw/1CaQ7pTx
svO0xs9O83x1x4qqpo+cFQDyiwPPYbT6HHF6cYjlzIxhZ2xLaSbBVEFmIKKdWs/z
Dn6y1ESi79JnVDXkxLKp898rkTAw4j4RXCfgNLRvXBCGxsdov3wMU7k8pHb8aPoG
uKotQyBW4codkw2lgjEOMh3sd9AdzOePrR971uBlehytEvWgwMFvYb+QWR+CDhO/
JE2iTQ9PiW9BfzRxSFZfcXdfSyShN678jwb43J6Tzqn5joS/nBhs9zG1iuzV6dAK
DQ+2vI+q9bzngdfGj32qe23fYDGsgwdANlPuFQcMqVL0qxT2hMogzqtQcKa3IgEZ
t36nPgTlob8Rx9znPkMiAdc73J4byXghiUAMUftvNlMQ/pBT2v+wn7/xPdbdLJGp
u9GrrBWVRz9tBq7EoKffkeDukKNDscYVsnE7JHedQQOuJg9YVZVHfsrlfoVX6JpL
SlQcbH3AZcvRCaAf6ekIEuzil1bWuPj5t6+64dewe4ZTgYJlAPObgAg5RD76vKy6
CGIzakG1/A8mO7+Q3TYVao0OAza3U6a3hGWgiaJNqxrBfP4XQutnv/izK91WXMCy
PBHvhv8WiouAa7Hbejaxn/gM20eggBlpOW/dd9zdYhKXDN8QnIqBlTzJ1NIjhQKD
Dl7QLeSFQ4opCWyDj3rFICR0lHmwXU3PjwkhCRDmiU7LGG8+QVo6Kh9Wsec0NLkR
8OEJrxOKQKvqPKAjcnoqN9jJq8Xmy3B5SScAbwO4zDh5tv6QtbaB+SeRA1TVtYSv
xt3lhzimKTxbYRkksOfjMjfbuNeCAmCjBHWMofyZFqF3cdQ+2xyjcZPgzqzVLidN
27Uxy31DZ2efFfQtSCy9TW3UhIrdGLT8a6pj4FJtWOayDDe3viRf08Sr2NR8WgkQ
u2NF31pdzWdOvgrfcXzRT8y4ybtq5iLe8/IlaKB+SoMPCFY/FyYVL9d2NT1nFUQC
aVvwbD0WtmP5xFqj2IeKLc2Vf+jsIxnbAjrCnSLA+YETSkLNGJTm+Yb9KXzEqNVR
Z6sUDzO1JLNdSgus/WKG3dxpcWqo1x8ztpYA65+P2uEffMpKH+S0ilfiO7WZ5lKG
iTB56RCvxJjLcrZy2QdIMBmkvyZm1yLl7KgJVh/YYZdHTBINnPF2oAXyL2stvPoU
KMC1NbTNN+rcNJ6a5nmUUGnZyyWF2tEEUypuzoyeQqHZb0OHO+TOgfiyjWnuVNur
Y9ymAnZ3wIXpfRs2z/WGD9CjGGVvYkfefwODoywO7co/greZ5GfTnzEi3w6rszbA
w6uBwuOByc+6D61eUTASYBs5kiHyH2g4r7hEsiWEfwpVG+871OO8rlRgSkyyOPfE
CyQp01Z1kn78hRTrTm0KBEsMM94s8AGXlGCwMEf5QWC+GNcJGFUR++qTbjCbIaBa
lv04t1iieAnukEHeHJ2AF2yJEP2ois432QH9K8F4PSOiYCzCawj0mdSx0nCexCi/
FNIX5X553hftVHSwUX2b4Q5dAC69vL7HA1ivsoj3ZaOvyKcDfL/vXNTpQ8B1aj4E
pSBrwM3bRmFDoUNycMJqAEOFbzqOrb2h4megtEIBku0DELJ1L2LusXw7p6Gz/Lpy
GqQYotnPwwmSrV/2saIj83TlKKOsIPE/qfSSKG+fidk097FC7gZuhcPLDO9tZ9Sm
T/CemxbqHRdB/E3Vx4zYzB+QBw6j7CZljnmVt+pOUWkar3rlUTUJNRbtInDh4P3F
Pgl5XcMUnB8rC2tDiR56OKfeePavuVqpMUgFZL7H57pvaxYr/yXGTeJ+EoR6xP5S
cG2oXSzExgb48vSAdmaP2a+q4Chbm5rjE1t7R49RLX5nXmJ+ZiiL3g/c47R0/erU
5dpe07rNTWEYbD7gQ3N5Hg2OtTfmbGvJZqSPqHIPL/Xfn/cIAXCQGgnzaqBH1G7R
ZkQfQBBIUs3rEAR9dpig78JlWcz9OBoHKVl0UGVsLtSzthbO9WnF1PmSH7696hhl
2hqTQaLgYZ7+KVjv6ZWPwwl6954BOt+kYkcQfU9afuyEurZEXQlFSztVvP7OujnD
B9gFm5JrA4jwa285+GvExPo+QKeYn+He+V6d9GSXs72NknPOHHP8gsfALWH8rTWM
wZHgB+RjF9rT/W+OWo0+MPT7jhpHqxDB2BL50fQ110L3sW871X4vqHTti3oFh0yr
s6oiG5bqBgbhTWEUvwQjHh+Pz9uybI4MXv+vHqb+gZ7sJvg+aHsKcDRUtDgQtAsN
wl5kaTxOqccMhuOGJHd1MPAbbvLzJh6ZYuKQ7fbBSNjfqTInZoQqC1dCwTIDLNSJ
mi48UaKVkhnkj0pahQ0vpiSrFJ56doN5SAoEi3pu8Ac6mTtkpu6YnHOnBm036192
Fg0E6AvOHyh6DbrLn+sSWEakU6lKw3rPouj36LhrKav4nf09DOZ+9dJBvxcMUtt4
D3ICm6Ia54FObzD3gAGv7BEatqOXIqqywMTrFUT1vfoSJpcdLoBDp4lWbDD+Up6q
TzDyrMIWLLqsPUymkneyzOZeC92yF2ZsZ5ZNMn3Xwg4aX+LbTpLfXMAj/BS+bEse
GLuuyEq5VjsmSLMMVVKgA+l+jLL0yU6SHZCVAyLlEzKE2wpn4xuNlAMoFi5s2lhb
vCdJOuGBAFeQi6bLf43PZ+2i5uCvrQZO4ju7Qzf/hS+CacTsgzDDh1/HJYS6U0vx
/4SPbtOf45IgKzBA6oH9FnxaE2EOOg4y8190bQAqaxVGB5JWidwCauqbY+cLCvqH
ekTxUp4L2q+8roix25VDhtFbvdoN1h6XjJZFfpalG4AaLN9a3fH9c+jWBfKgZWSu
9+uygaxSyO7prfKq9CSFhUmtCGiVBLZgy/ok4w6kJyWCeimIl0A8QTcVRzTnQM2C
TLna2BXJQKDGZUP/nrcp/LsVsnCgI46A5M1fKnNGNe8KLG2Ypak4+kc8W+6q6qut
TeYC0SDqQOpNeX4EAj2zmcnoPUgMygcnoWVuVkFa5a/trViSwlQt22E/Sj2akZ4J
MAt2FV6Yvu3uCtEMdCd4hFfXwU9PbanTsh6qZO4eqGXZWHTL9ooFQzn17ij8VFB/
Xch3nj9QeXswn90vAHIUpillMsrfRhaIOChWnORsKL5NCztvnaYpQXl99Mm09T45
1H6cjY0x43vEQUmHjLmhz4kMvqogSAn7UdDnlS6mJe7O/zG42kFnhUrwBokNuBZQ
dEynskdtaGNJmFS+yaKPdpOaPlEzeY6dly95dpxaY7LNq/iACHSaNUi+8IvopCQf
+h/i3YHJ56RJEGnU9+vbyxAexgZyFRQfmmHbHGomiwtV9fFhvjX65eM2oiyJVgrK
7nVadTJmOzUEsGhiavghsKQGBKMFHFBxCaj2My1XtfoHo08G0J5b0D3rgPQqbfWX
otJazI7RRdW0A9P5ztinVOeNVYBvLbxDmMxMoRgmktAolK7Jprh9tWsONUjR9H5I
3OqY/epCxtdE6DEHpTKPbW67AOEGOqlymTjh/h1Uh3WwiGeUPXw2kJQGbxtwVfAu
6jD9tGQfGTUKnslZv7D88XAHM64Y99eMZfk+gtQOw7HpdFQ39r/oQleQkwRUsbcO
LPM9ZNz3QJzsCzTlIrHkRjAVcwA2HLVScEWqT0qQYqP77A/WCTI+QaEEO0Rm80Oo
jpVpF4nbXR7X7krTGbU68UXinWDuULjF8Qzp2wBYdefkOZ4F/n4eHnMIYoNtOeUm
MV3f0HYTlSwbMuRT4rRNzGkpg1wDdaXmGhxTx1WH6gMAPIby04uCobvE5Hdm1S41
f13hty4E7S+hxbBzwWScdYJ4XQY/N7JCQQ5ktelZYdplrOgPeVtNTFe1R421L53h
E35hq3+4rHwIQ62EnYgEP2O8wedzpj/o+xGM2jvtNbJXATcOubMC2kmIfur/Y21y
GNv+V8EcYjbq9AJgATSP4G8khaWqDW5l2967wQKR/+XYiq/0VrAvrO9+CzjIv0b9
5Lb/dsqDFLZNDFpMxYbtcSQw8sAchjCkShkCQmEHhoLLKpTWIcSi2Q+rBENWiDsS
oDCEZ7+gDlZl3I5yvZJ9KyxvXoYcuhttZP/5GjgOsdJYs4JZSLS+Arg4UEPxS6A2
tGxRrWU2QFpx+6X0NGyVRj0WH5Yb8nqQX+wKba0R3E4RFq9sDr+eRITdOEPTKFm+
TSDAahvrHgKwEwhs0HRw/lM4cIMSSk2/sQ/A3qJfQyxYLEWdCJxeRUQ9znb1hyip
BzC3PEioc97WqNi2OVdWgHVducnxkVQ7vfDv3xfg8QOWIsEf8tIAMM6eUQ8FVoIV
oxAGf91ufGXS9wIRGHM4F2ENp7SF77bJQmBppRx/FYtFZUvFl+4TmgotCd37dDyO
CV1hvzX8tKYpWbr3giDUGbeI5iMwf8gz0637PRMduJk3JdWGUj3B3bMipZvwQyN2
xIWrpJH3ZAP9EMc4z0aCdA6ZzCLIbCParDKgXOLCxpIa7Hb3rVRArDfMQsV0EkS3
lDHg1+x/5TAvquZq1BTuhzo9Z0sQuRYo4qBbsNnK8+G2Q9eGocOqGdWnW6R4KfPL
/fLVFBxP0hTGRRyWpVAHSDOPu/bYQYJqzt18DIp25tzitQfYUslCWujl7uwKAAXp
eAfuxeCteRrkaT0UWlJ0xPEq0JL66abDFjEMYl6+cMFJgl1HqLT1jQAZ3ND4dw19
B8BH+2+pimYIUl2L0DAmZtabS13Dnlac/FsV1NYoSBkN7pkyQcwVN3Wbzh6MVW4U
LlEB8q2kUOdwl6n+lXedUmV7kQB3X3XNbL56+mSGkeHk7UYkRcRs+Pb/HIOW8vav
v82+mccnB5D/ZJIzkBuPy8TxNhDJAqvXMGhkEdc/Qm0IZhibyu2qKm3WJLucVsg8
USO0TuZBgYVt7SqBLuLqVWgVBajRRJpernG4kInP3fAfB31rULr1etWGER7HnCVv
kqNXfjaLT3TNfMWRstmi7zt8JeK2TRWyf1QGMScsCoZ/qDclnM1L6Wl2pthwyXcR
WktCUUSts0YvUdcZKmUUJhOgFNSsDsBxq679aS2qLhXfNB+cXDPzgcPr2NJwcXca
yRLinLz4QtEwtxAJwiUD3JeNvUo1vg90bbC+eJWWyOS2/1udUbq45Gbrnbm0gknB
zBAiumbBFViVzY7GKIVzNqqpJMBTKa9FMe3mFgzh3PMxukU5EF4W9vzGIAllVm+e
NNnqG/aB8feBdC0zeCbgxItPc3qWWUSV+ftnZFTMjrXz1CYgVUzhbL5IUXOnQMM5
x2L4d0UWi/MBjHqaWc2Ut1/io11B8Jee1bJmqP6EwjBiUwfL0vPQ7DXcBJE5vkHH
NF8xtoxwtZctWhS3VF7XT3tLRc3aU+/CZTItHWVIObLy4uLTZ2/dTJ2RlLK6WJ7k
4XARESMS5rvt4pPJcZdymWi9AhpsbFc307apfVOPwOVQKi0MncTVB3dalKRH6M3m
iBc0gKpj3uNKT7TTJr43Kc/0SGGGJEpxPv7edR5qeu2B4jE3FdccdSh8TN2Inhmu
FSCYrSRxjKh182xROus2mG+EyPHp3C2N5onbhcaN75mV063OIilCgwEgA0ZqmukS
Me+y4fgp06EmPJZq6sVUAgaUlMgWqxLzBIHlqWDKkdphl2P8nRvQpaoeZ6OQRMnZ
UMy37nsNtnYhVdsBkeKa4abzFZriL5F7GwUjdFTK8QX9Pon+nQlWYcfu8nJ0oHAl
qGbsyaJ4td0BiMEOBgTx/COgHIsKZ4rzyvYUFqoiXjMupV+ovapWGIZ2MwMb8ZsW
SFifeevtH4m94bKne1QKqHiKjcXC2GW+Oh2wMZI6YFSN1lUrocGhiy3djAoWyLmg
fvlBoE1K1vEsI1YngpB155qoDi/89/SYK4v1rNP9n87USYnf0LMnmIVHQOl3nY9y
rt+9JLie7uf5pKnEJyR3co9fMFHG5TQAfibaw/C/ZJLb/Sc/Xq6TMMmkoJ3OhFao
TUTkPaIJLIvsG8d0uapN5tNDVuxaYLSDDdLun0FSp4TdUTSNBfy+yM0OSHVvD68R
6DoYSKfzRZ61mhDLqkK6ksdMf1WxlEr25cjgCYZtHQ9SFXtJmJRH5B5hvrf3fwV/
InQ8Cq8uzStTM0/oCmcDznw7nQvkELPuiFKvd1Fo+4M/Z8Yu3gvH31YmEsx/1CRB
dpczMukED7F59AopLD6xdOmlQTRHwt/YUz8FS2A8yia4zFc1jyYCAT5qqxGiCRzg
Citj3Pi+CRHMlhCJoZ7+ytiCJbt6T1ICe8u6YLnu2i6tysIGoZqhyPJ2eiFzP1bl
h8F6mBf5nbzu8ZXZTB1WDrjSTt9F/8dPLx7WucaJd7m6c9Kvd3u5kLXuF9qJGPaj
cx2v6upF/IpaHnXE6n7iHfvh2M4V1YgDDKV9kQ1JGJI6zHF9hGbg5njTaaCPhXWe
Obcocp/NwHqfxQKZD3Yocqy0axmyqaxUvQ/GH0Hxq+jKu1BRKo9gZB9wiPtJ/TiM
YMsF9C3NdkGeVoYd1nOGYKsWzwkIr8Y8IxbTvQ91K/xy9EpQkfBixnd8toL5Lnog
5uWD97cSkLY60Q1ywsVsM18HtxasByOXAx7iXyBPGJsCO/bxldcwV+Yy0f5wgAnL
sZsiSb6tB1zlCRrSTfblJk8KnANXInDQrCsdyrddlVIkd/RHwHRCWC5cfXxjXOGX
ruva07SrE0p12uas81+l6+EsjLWyje7BlO94S1C2W5yQbk6uo1W/MPo5vm5GejSt
z4kQ5e9dcECrnx7EFd7pqIY2la+KcaeZLTwkZiv7dDLUllP7pmsDiizCpu651zAT
C1iA8L2POzynaXjt/kevHo16xZMZUFVOEyE/HZb7vm5x9LvHMRea0QDOuwyMFoiy
ihLuAxbyF7zyikyabk8BYHfPef1NjEnYD6hKEtQKa4nhL3hdJ9kUILfwcR+WmxOn
dYKZr8ygdJrnYyKTk4C1lzJGMlG8cqnFTlJP9C575Ej6IsS1ePaJsMalhJV1UuWE
x/f0cEB2dKaJs6n312t5ZgB2zVJxl5+NdQzK6e24pfNEERo/d/eErWnPsOwWbnI4
Jv3tuymxN1vUP9LjmbED3aw93LKmkMZDCO/QAJIdJovFhNJBqyCpPuKFeN6kKdKX
AYzReXTg/HstxS0oB86yxu0G5Pjc1SFQEkiYtCZNB1c6NW4/etrKlZq2EoreKqra
Ha2QWlXKcfdZ4VRcP3ClPFrNLnSMwlqbbSUkRprt/Pi9sVueez4Qa8yJzTxnYGrf
2sjEMEVIUCVE2rJGmU/PmS1y6/qXSeeRJ6UIGKsMp7vSk4iegbjjbMHQ5sHE0lVI
v/5rG1U168Fb0RRXi/Uvua3P4sQELiji5uO8JoT1t/ZwlbQH7Wzau7jA0GYoDOQY
3W6AqUCtkXfTDVfDGGcsP9x8UtecxVkGFxg1UehQJJBFQOpX2gfn24nA5JzfDyfM
IG3b3vV/HwU0fJ7ZNpo6qF+I9sDY5u+y6tApJ4jXdjfCn2ZLiojNdea0gWhrt9bA
cTAoeRCTZ600aTviz8kj2+3WokoPQZMU6GEQTsqkvjiw07QdRnMfQa++Lw2c5NPn
JXt+Ztc6YrQhTUC/F3RocfwZrl1JNkUfISm+iVnXU0OODZWv3UrR26CC7Y5xWo0E
wUb7sR6XAygQK2pvSGd0oEb/3znBpbLdrE+7LAXmwRverUjLakV7jLRCnVl1Z+6q
6pRhAWefltzH8icJDJ/6Y4CKXKznab8qr/84hDnTNLVY8InJSjWO/P/pcTHjrMQ3
eHk+BibQIfuL7wccqORb9llhK6bB5GbS8IBjKlS7xE33JLqtLSSmsKlMzjgq6j5o
8GT5qMPWLzfDBfBkbUK/++E5K/7hG+UEMkIbx9ZKzTZaE75RVXG2t4s0kIixthr9
f0v9EXrulZgeZKYY3jWRxuI/i5FdT/3kHcvF+jcPyWkYu4h1KYyxJg/fCHpt7Q24
tm7fPTpPJ7UVHnrAypIV7hk1c6fwJBubXTOO1nN2DOr0PWtXyfPV/b4rXCGKyZs1
ZYP9SA/8Iq9qnrcx8xIcXdobyLIDEEhv6UOfALV7A0JAVDoeps24co6w4t8GYn5v
jEuYF4LMfWteelqHRaJ9zy/R1Jze+zKy0iRP1+kHDENJsHFcBFkWQ2qakxZceRbE
VkZztfkwabNJozJUc45k0lWkf+238b0ZdYHcWN56ybKBvtvK2LTjgu9HDvB9Qs9g
ECZzoGgYVmNIjyuzBIvim/R2Fh8N1ahE1osqI5eN/8kWATy5gpr3Gk8uzeikTpkg
GE3KboNqow5BiYsyAro4+ACgnOQYdv0Fi5yqW6gDlgQ5QIUi0SjvtHLJY6jazxzX
XcMfqbwx3RX12O3cgvgBfAIDjJvJk4pb6ThfiIsxfSvWEyjBn90KOFsjEMAAT3uS
GuPBprOcwKHUgBpKiLk4qWJrZo6YaZyu+Tvb8oWkqEEeyt9vngYVjdaLEjoGWm/k
iXTMXa2sc/hfu105kMZJDLJ0TABibMPOvkiSlHvjZMqH7X8oe00/PRjJC/5Vicj+
5WLkGP0GN1paRQGXuEf9yhy5V0ChN7Nj6B/nIPG0oSUS60HKM4dOzlqx1PXEwiWT
oNuFp6ZYHMl02v6mKCRJ5a5G9WSpIMcC1ub24ELXjz8VmPu1M7BB5w1jA0XWjt/b
2pqv/Nao79ZJsdhvfXb7/DH/LDzrYW0FTtYBfpnOncwiSK6wb3qbkpMy/VtOI0Yt
sJPvZojvUa9ug2UsSxYrgIJY3CgB9Zbif+IOfU85x38q83R0EBTadM1NMFmD0YwL
8pI+oEjiMvNMogF3N/GxeLzdFLvOg7g4ijLdmTbbxEOwL63Pc6PwcfdurSZziuC2
N/kVOosUOnKxyg3g9HzRPQRk6zaj2AmoQPD1IOcU46/QX3r5lhSVGy2fWBZTN/7W
nytmefPZ4fNK17kHWnAqogm1Ix3g+lGvc+CbhCh/eBE70wwjrbeYP5mae6rmlzzk
B42KrSkJeVsVyPaiKo9XnDfHcQC3IyiCOXqHI6BIUwtsNyqD5aYtub8zHAZS3hN/
wqQ+Tu7yAIBhsgJ4511W1++9ypebY2ef1O5Qlw7xJwNwp6gYo5DWPXHI4AGd1PI4
KkDWg8KcKwzHl3CTuemCBT5eLX3KearWDYrfPROSLbGcCUUN5P4M1O+bU2M+MCBg
Vl/xCbA+DbOP4OfxrqpztuxCqwSBsuxW9JL6rdKhtg8k6CHsdZfwNUyi0oHxn9el
eeI3CBxpD/IHsG8RBhFG6NXdv5RGrxXHfmWo7PgjAQYKX0HSDtJ8pva2mrX2FkHl
8mYRNPbTJA2w5zZhN8a87CdRelHA66EaZTXQt2vMKft5iIUdfZuT+nlCR3AJ9KYM
I7ii4SI6n3xzvTE2mF31apUxaCDuC7pjkLNH/XTzO4NZ2KQ/+3tvwWHub4+47DOX
2RWay8ELoiVerYrVKtNlXdj768eJGcWWM5YvF8XWOe26gOq71NtGjIm+WSmzy3A3
gXtCCdoxytQO7BRl5bVfvYzSK1jAcOuQdnuYUjAyHgZqWyjiu6O369KLVbJQlbdo
2cRH9LhnSS3jbRT2voz3cOLNFKvjYiMdIY+YgzbjUZ6vCu2G+5Mcpe9fvYq8ohsB
NGtSxlFvp5MkNJ5lAYKBkicKdkuP4rstAwfowYxG0WSKMKGGIEoBIc2TJJgVhZPp
+YtMSuwIb/vIQBNxAbHhxA8qUdPjPupyBMy3klvl9FTnGBUwWe1TnyvIeDp8U1ib
ELtu+e1oZDUTniMIW/fzttK0Ca2ITFggdERs+OCnRIWn7Z2bdpxVzzyGrSetdIGM
fWXy55HEV3GoUS4tnVnClI1OVeZRweowmBKFN8NlGmSSruW06zAgT8ComL/50n45
ZrabmIKg+JioEcO0dJAgZZuWTtn+tFmy9PIcoK6Zuycd1eRi78xg/i8CmA+uRZHv
Z1q77gPT8VGIbBCFqpPVRUXBLClWBLXHQGUR8WmnxtD0gruynPBKSkBNLG6madr5
t5Sc0zPRVe57+VxGnXnaspMO+vqGGcKz1Wv/TXO2FsS/u/i3C+Mbs/XrGG6qSROf
dlA9CcbEMzdJ/VexF2TTo50bQgkjAMe4C3rXDwUmfWEu2j5WJCEuk7uxrwvGOl1Q
Fape2VaZ6D6udcNzym+yiR7J0EmZrXQLFUyVKFNQwq1AtrEVRPiey84VjY8qi5sO
roeTtHlTeLKUW6dk0PWuHvdYNdnEQDZA0VfuuNcE4AkGKjOeJmuRyPmyxPvn5ekn
4HxuRM8/h2C8irCDIHA3Gw2ae03+c2rS6YpjFQ3kIyVUZhFixsOkNvRZIabtoz74
1qqWnU+tr8lafYu1+UtveSVghLzGLAaBnrCXveigB93TfDN9XekDkVkSIavJItK0
4wtjF24+W0bE+2Smii3NdX8gpYYws7E2eGyK3M8JWhhFz9UindqBQ3pDI8LAEXf3
HCuhesOZhPG9HVdbLXsdxIGV5ZCWZVJq/OFfbsCzmbDay+vXsyNZRR6rZb792X1+
TblxVTwHbreq3VBeYTpN96xRCGSB1qvvKXBMRQ51VtJKkHjiRFyyuw0EmDIpplII
+DdPDRt4loYGuweBBEGL1ohUYTCorcZhjxlumbFf3GKvR2eAIsYvdfzVAMES65my
tlV8z652KHbqBu+QyQlr7zWaqeywI2C7mWd4QYHTSjHxs7D5Ckz9GN7y+cnb7r1u
I3eFTCGMxph2SUPtVcOZffCuXenS1dHJrI1TUg09JQCi7F4HaseuPcJMLC/75YUC
/eyEhuwlhEdwC/XEwrkPJiDpBvoJs3+ly2Wa+BfZPm09urh6Lx81siFvr+VsSsK+
wWEmYkLttcBofNqL6GvqQl3TrTwRB33p68xNk3jMuUXw4UVEOygK2ugb7AaMqRE7
IxQEga6em5XtM3AitwuGSr4KGkyzQPMiX4LviAuQMCHcHnmV3Rbu4GSK7zFq8Q7z
MCAzf0Ve+JegvgESQEZaJDOiN9Y/GTsrjJaPoOmOX+hvRI6u03J2h2Kr7Y/XNwY0
lrL9byHBcRdD+aHKXeQCll07omdkCWX9D5hPw4kZnSDl7/PYTvPV7uMK1iMOqPwZ
8GqtRQYFRBdIooedQzoaVQmWLmpb0d0xk97WdSYliSkr0KBuYI8kW9SY+n/sc5OB
MWbJlEH5cMGnSs4HGvBe64QuIbAf2Dm6fVxUiEe+X9VoCdsLpgd/3h5zTgJTBu3d
x1YQ79oGnND28oMv5v7p43xcMMWf5HjAFOlJkx5gmHXNe8APnnSW4F4mrsNiI9uO
LND8tcy5GVD3LXTIBh02jkkttjdAFR4WsXEzpRcjcgpILIZKWZxT1AC9HX9SI3KO
y1jQtzGDtbS3wBVzGQkC2ctB1qQifyYIOGjGcW535xHPxWM1mxXcvHy0gr5xGxW1
/RFj62wfnF/X80I59O5OEkcRIbTzOv249BFj6AyLgPsRYgu8u8PI7VE88oLFfEtw
D/gAUQEcvTCvYkXvuF/zTniFlkWnKPlN2SJgFhyuYQZdN7c4D2ZMgDKQqovUplu+
HEg3VwN7ZUrUQCjz9rw1gRqX2DxThZS5hmweOLP0R+/VClFUJWaDaxH02Vx6AWFd
bNmZ0zvBIkiHnuZog/H6KLvsGE1yaDCb8G6knNa+J5e4+KzPAuQUD68U+aCJsSzB
LgVW7i6cOB34jIV5uAHDKRoAbFL4r/Q4i4kmZ+0RjX/af52bXGU5ZJQE8AWYqTgU
a6DWpx7jt0oNxhopwqvRjm7yYIAZuWR2skiTMZpxixtxlBW31pXjyfyZUxn0T+Z7
7pSJaspO40v65FMu5evJ10AvMO/ev0yVdMR4OTqCTDxlbpxdtUGUTzmHJ+NH+TNA
5U0ZkSjaAAp/rXEz7jE2kTYmL3CF/i6z3g7kBzMMqId1jCqjCifM8abfffKUSt51
QEfPnSufZt+c58KNC9AEDbOA1HVj2tm7X2SyjimoRd8wris9EQcF3KcJd6UAhrFM
ErIQb/scoALUEFYuYEo94n7+vMZsUHnOfCKeimsPZ8/KQF+nbAHdHk+hLcqQ3VOl
XV9cVTF7vP/tbIcVyOt7zthOJm66KDsaM5ey8NDxLHpiQISbF9obBudh5OGrthhH
lAYOfTAe6cO594e74nQhENA0iempWGrOmpKqr6QBhgFlzdfoNJ1+Xvv5Us2oeUDQ
ozS22h3UkjPrwRmfuNbmGYB6GWq5eaK5iGE+HMO2yidK8XFDYWS93oqS0pMal0FO
80SfuW5G2Sg1bDq21oz7jVszzdPmDBhmAmyvzLWUNTIlCcdVyq0xlSJjHLLO+zTB
pzQPU7lGn/AN3ApzwqtUKjlh6/2FHFNDJdQTo7KAknvPSfr5d8l9HLCNPSLA3azk
l7PWk7OI+Ze1uVSu+Z+qqkXUfZBPvzJZodwrtK+81B2gbU2UjolNUwg0LHCJ+zho
d1gKhDkd30KF86fGcpTnQYy4yf0beZB8i84rrjC/sVB4twSddBdMb2h3wyZgpRDY
sa02sAl+imxVoDo8JPNaJ7PJzDTooRopHx3qa/9KyBYc0027WzmRwiTfAupLgV+P
jJAyB3afr5SnXiQ9czsfyxAS1FrwSy/Zi8itfsE1hSMGQV3HNHZL+QbBpn1kpEel
SUn77/+Xk5UuFhLauc9kYf8MqrOYS3qTjeEq8GzPiEoMud1iIM6uGrTohjcUhfq3
yqUO9OD03a9ymF14rCFgphZ4zsBLjYC7R/E8Jj3B8+oWCKmsn83CEzikYw9iVfXH
NngleNva/NKP9bmV771LI7tksvvMJjL9M/YOsdl8WYOIFg0Vo9jEGawWdXOGkEYG
2/tt1yTGVOhfPhQj15OWoIC+gesBBaPunzEuPisBTSu4XRoTmxXWlz/kX9wAiWG6
G+2mWcfWecqo+OLqp818YFAArHhEyy+2mQpxRXJ6kEavSA6jeNLR6FXn/uNmI9jY
i9EmS5sTAkoAGOVW7TNReLxuqHzST2Y9c6PwZU1M9yfc+EC6OBgP5IeYu3QyxFRk
J08F579R5YKBorx1g8/jsSeNogH0QOjHrf+hFkVm5mkZezucRoiZ4ikJ3VurSWsz
Voay+34/lZxSYhG8CSjucTuVMZ8vJzAEszN1GZrRBj9zOkab3QJl9rD7wiJiTHrm
Tj9AqrQ/hXzrVcmTg/2q1WP8k/BNPByLOqK9RP8VsczkB/OymoyDg/4n/ZomTC8S
e9Z9Fddurt2Jlj2WJghEOyAlt37TMmtdhCfcZ78ugJBprWSw9QabA/gKvEz7mUnF
u+Cv//0/1ESrPJKRLbB6gFy6lOpTAVMVZyjuQi3zJJLHc5zjzfx+VDxC+gduYPn/
sr+GugI+QDjL9YNnoYATghn5zkthh84XQ6dPFA2jI3StAtbRWHGHtFoxqPQa6Ju9
JLe9TzuCik5MhaCLX4FdDFq8Xw8CpM6MM69mN0PjNd9BtWDluinuMSc5t2oonAbO
qzRojHzZ0fbhXxVk9xXT9Llth9dXch2rPyNXz2cYkdWhp5eGarZkariuQy4Q/k9l
IhBniv0EnNZNu1VaNNzXUnefTli/Q6g6H/edJLB3TdvDphbDhDkG+E5sZ4ugA6YD
qyJpWapEYbjrfIXTYNiQTZojAgRT//NYKlsJssTEvZ2+6+wPiaHIqzuK2g/M4JE9
uGnNZBF7SxZk6/+OWWU1HcPeioEPLVaSrDpCLHPNY5+CbPcsg/Jz11cJYwvSTQ8V
utkdBJS86aFgkyMv0lRud07xzwza7EIRY+D/dM7A9tDQDqYqjKxtAm7SeSyXBl5I
ox7eO5w5t3cxOcP7CUZwpYwcLVD7iZ3+VFOBDHFG5rjXzoUDE/de4HnIlxuRkfxu
peioqUB3GKvi6rkX2aE2O6q11RQvpA8cwywQFytlqKtJgAHfcNYA0oSV7qBGP/Hk
L/wYBa1xUE5lE5OABzdogBjJxtPnVgXAb3d86QXfZqEbyoQkewESwzDtDc189vfm
xK2HE7dlOrc4nlBD624UUUvQ9idvcwkEkdTSC6AIRFMleWXJOMaEIM/5Kv8ubDld
QeRd4KVK+yjikMSbr7MkSz52wq2kqRafAS2X2qWZG6Ch4jjolSoHPj6P6Y6uNbI1
DwFUy7TvJpm6SfIy0/q28tFsAnQ9nn57n37YERziirxiaQoJYr0owa9SoP+B90xI
KUX3143KtdnJeCtRaZDMMJUoj4g91wyZTrZS/9u8nftPfcnuWuj07uz4gx/vrvDn
k/Q3YxkDB4GZ1P1QfJ98KFUXc202ucAupYjLryjSXLHY1fdzzghY1CqDysBCBEmx
pSJqmF4j05L4n84U0dzMVtLFjQbvb8IPMNE+L3JVXfG7XXKAoZHmzHdwokS5rfzS
oeNTetEmQh5txUahXazS0EthKSc663gAcF2j2xM6Se1ekIiZfgxAV30Cbq8xGqLy
QW/x/84DDhjXceal5BfKD5s1m/7vl7d/jfJTrEOswFfiDYN31a3qDp0oqo+icZrS
JsnCRfJYQXsdLhSgU8iFE5bD+m/3RBfQNnpsBOrn3Dbi33NThH2cyg36S5yfnY32
UbF/wD0ZBV8iyH6W3snDjQEK2H2ZYGg9q6vbHQ4v3L037JUWsCF0BIn5PReK9x9B
eTzkqUxfg5LyVTCF0XPDr/nO7fREMvbEO51sGOrNC9bEkYqH2tK9fCRFxswpQBsV
fbQDB7Cl/LcbgZytTkm8caAugxRX6J14tz6x5Xsg7ZZ002CCXTm9zZ4XtVeDK31G
7brhXxagxRAr+wChgt2jlq8tbbM6ldKH++LdXxWwCPUVEs7CPdLEVqzCH9ZgBKkK
hk6zniy5rIZJKAd1JrEa1au+ob2n9LNlNxHDCALN8GCPUZNj2Na36vWol56xhIsP
0hIt4jVZY+/Bk0JIqkzQtas5F+sWyX2J7lSmKzKZWm4dWv+hffe/jKUagoIxXB7a
yjAzmd6z6A2HRpG1AxES3nZ6NJPz5D8WRKx/AHZe/4r4mioYwgDTRGMeI0K69WV1
QIsvTEjewxAy6NLKOZ8CmSUOIMNm/v0gKpmwgMSgi+3WxrHLUuGYtAp/86Ygsz6E
Yclc4InvHtpmizApMVjIukKR3FznEPzqmHQ6unxW1aUdm78IHYZLbaayZ2ofmCOk
TbHRH2y0jhZUBLC3zFP5NMRhSYqmX//6Hxee96Ficl2cAo7e+OeZEA6BJWu5nT5R
qWqbthE/hLHRz7wPcgw1u/wP5bpXdErCaukZ2lSJisJTU5QYBjZAUczhU7y8Mfl3
FaZ4+4pvLUN1j/0MVyMkjaijqUJ+asI9e5jViO2+vww2Vo2Hxct4ajLhF3k38h+n
FfTQ2RTIkTLd1Eaut9Kj3DnOHDfEGHZ44vx9lOadO+h4K9RgNIUSemr8M8K+6Eqj
MI7XYFV2+WqUuKVO6yNX/vxMfEIUuT46JU/8+w8lfLzlQR5FlPaKkMv5jqQn5h2t
CF+4WAxT5xvSo4732cjW+kEcjL4yTPKAiXYylNEOgjYhTkH23n2Vl/Sr8tGBv3XO
SawmnM8+rJBBJtyT3bbRxeDo9INb0tDAsaePcBvkwItMBcNrKyxHux3f/AoXXKVD
jpb7ce2qQfEJj1eITZt4jRDEaSGNzWn1vyPZFKouuZsCtExW4g0L9iwQXon0SKLa
0Y+hd/4/xMnkI5sNjTniy6gIGWpzqmkYoVNXeGr6qmuPI55sLEUFT8idiLDH8agh
V9W1ZaKOJaxyLqvJRzzg/zhkP7FN61bbGzog73E5htEZIaMhR8bq4FL9h3Ws9/2b
VpZXKQKNtokWMU/AT0E9Si4aK0cfBLDb5xBPMbErKoRrbYNG9zX5Wc6q/HER18Qd
YUtwTB7VH0eqM2f5/o5nBGiqvFfZj9QsRHZxl8VAdPNwnkJvIBnjXrMF3LqZVQxm
SimmkzU+T11njuNFigi+7vlxczD9OBzsbB8i8m3XgWb2+oFHOmT+p5zjB5I9ioy1
GqJtREWn5xBgDM6uuPwkISbJFdLvVPIfOpBkEQmw+Ozo4Cu8SEoBG/yAPq2KIPA0
qrKGrV7qQi2Vj1+5IpB08VhrkrJAIzBMtCOtBgy3jekWkiNuXzH91kmgqrWRPHBX
gf1Xo8MbgH6hOr4Xa42/x+jldMoUoADKJSUJVFXWQeBlrDx5NwU90qFqkBA7OV5I
M02ZuRCfsOGs5Gnv66+Nfi+kdsQqR140tjPBK8IQPusiduYFJnOtp8Jj0x3HlDjl
r+lwMvGGk0cEI1TBoDSmpsBeZXyJIPBk5o9BNfarJaMUcsfogzF6xZUuUcR3oVTz
knzTJToXjdf5G1cuYf9c1cUuJxvO8q1COfAYWYEDFrcO3nSlmDPD0gdiYaL1uIQU
kqLI5B0pFd2Ndm4ynSk4HLoExag0D8FReVtqXd4qQJeFtiNs3xwg/0jOj25oX/aO
jMkoMhRCytAtgM4xLbQ88Wz5G3xbqaNI7MQibVo9Cm28gTtHCF/pHBlnEX0R2z/d
wJNPjjicJkVyJEoQ+RJ8CQvOXbouMBLCShBpOlPECPqn1KaP2lnaapPLURttCUI2
iryYKdTfRYx6Q9WW7pRaWBDTuX5VE44XYoqbJi0HH/CZHEEEpRyKJ53jBJ2cYqyA
OLHtl+aq9O1/EBrkdEBwpx2fewa4Os0exvEYVdR9caSz2DseLvq0/9B1hAu19MMJ
iQYIHdZAL0K1Cu7oaXmIvegqkQhq8s5TFq3gYpupBWOQG1WSnztbSYjI91dkI25I
75aYwrjbxZ3fNpy1ySfArclGrL6mgEiaRSzQWTilc08omlJEEeI1YAH6g6HRuqTu
fKhUewJK2LgUAXRrkx/iGuDEwTPTLHl9EB0fy6R4MSCe4jDnVkPQ4E/zl774KFlo
wq6WLSoZ9W9CISN/oRlSXILIdq1+/drcXcRzo/4ttGL75p5LxWUNqQ1dwyu++iqA
/wEoKgzPpU9Ss4EUQBkKBP4C056ZS29mxT/TCSlQS5GAvEuun5JQruLKvEvIw8M2
vJhAwf3qPnKLUQvD87cQdUrJRlYV9Tv+xEDzscF2HYLIYWkuWGwjHhqg7TuDcUrE
TNjuREDq7Bcq+DlwlBfEa6dc2On/fX9Tbp4AQzZwYGEBV2q42wQDCeUWGqaBOPTq
PaeYlun7jXoAvwuVX2PxHw9aeC4uTJ+gW2rybgbEyttv99xY6BbG0Wwkb/Qw5jrn
2GERqLX+5U+8kn0s1Lh6CHygPHyIpYfKLyoG9aaTfeZjsf8Ys+1Fk7mpV692o1w0
v4olSrl3Fw+FBhlJcyasq0LPHw33nHxetYDPUuybqkIG0DApuqz4capHhTJQDC8A
77RpuZWxgtO0UubbcWRqRH5TijUl2S63i9yZo+c+f/wkrK8hxeAWfH8C32HPOZbh
VHbfgM9RSfu2gzkFWf6Is4IYaeLBpz1j23avKXIbQ/AWCbj4hkc4KClB0yWAGLOM
9ZpQgf/vp3W8Tl4389gV8Mxip7dfhWlLzA3lfVfkBFksTxiZdtmDqnJvGDB2xm6F
pRe61hVZVCzsyBgl+1zBQ8EcaVEP9briQOOG7cFz4K7Ua2xyvVHFGqyoPSEbETmx
PgwRsQtbcrAG2x+HyTnmtDFMB2m62XH1nz6jkWy5CdJb5dqP+UUbuD9S5qJN7OOq
sTnKvEiK5QptfuMTJQHYgc+4mgi3uuR33SwBqihaHKF8gw9KP3LcsnZxN/y5KRou
Y5bzG3UWKhV0ccrIgBzoxWSE6Qhp5WTjU1Q1q6wYUSC5jrs6TW/HY3pZshHtDfDd
QI9w8qXdggwh1xX0uXTkI+MhRGWFVqtFWgdrbPrtsv2/Zk77WnPNRx3ZZJ9gcES2
ToqVH37GlRJPrICS8T7el1ngtpT2qqOqGcygOKXGHG5gsyYn4VmbFbeQKkSO7Bof
08FSREqRBj0Im7/XXgsezBpzdOXhrf4evhTtx0NJpe5hCoJ7dynWxlSv+942WaVK
YtiJCv6LAn2S9xkx43TI+oCeeCbuj1msshCWmH6Ydp8YWYuMhUf57nMzr0qWT29V
ewL/tZAMgVni/8YXXQZRKVDc+TKYJl0gJCN/R3qxCTy0V4XYDV2s/oSVppuHT4wo
aVYejXdtAgp37CZCNmItHKib8W1XLjib0QARQf7UE9GcoFJeAma/3S3Zgd4F2nl8
SLslySIk+XjA6nErVPZg0JHo637XkckfljvWM1le4nDYieISKs8iw8j+Jic2UJ5Z
Hy5waTLsqftWCbFW+LEtMHgk5+akPEB9N3RnH99xjTjHbRp9R9YtsmzrwJyQmjl4
M+ePO2/pNxe9i+/az60dMuRwdbTU76AFWuLmzEqnOrpogIElXDIo7uwVsAMfESni
fX7++rWAPLKcIlBjZXVyYV2O9KppPWkcADsX0FJhf7Vqatrz/Jesqwk3rUV5a+Wa
bgZfpykxX/kbMw8iIGXRx8TXznbJD86cO2lkwjAYUgmOJ1OalJOYtBmfyrNAD8h4
gRmk5ZQbqW7FYZAd+MTzYI/rNO13DRyqjzOg9orycZ9LKGkG8bX8hraypSxufgxv
EcG42qtt06cmrDdsvp3rrx9/kUH7vOxNXLovEgtGhWsmx1peDQVTMttyUAaeBUQj
ZBwxNgC/k9b+pEZgr4N0jdAaU7EBn4NYtDGxhdRFet3Rnw6WRZXwOHb0V4Sm0fRj
9ZP+tPFcZ1ATfeMxRXcq5aEx0ljbgnR6o+xqI9lqgMxIc2Z/cKwUaPZzfOh4GeDF
CeS6x3iGc35eMahn0WqmdOb6DQC/4CZrKByQUVeQUSRKUeJg6QK5pwcvWxmikfjA
q4OiSiCe8RGCdugyIxw5FTYt9KXmmCse61hIpev5LWiPq8BzOISTlcHEuvAcYaoS
cZdL1UwuS7L00YDUCDIZRFPniNZ5MBduFY8Sos22RZRF8qMiMyoiTM/LSYGgSRTY
4ZdDO5bMOaD2dEzvebDM6cZUIhdjPzYdk/V+2MFSHComfFTnEu+hXt8iPXGmFiAM
eze9scmXnUVif86EInBFDuF54u4pjD+CJsCwf6fCaH+38OLsxtJpRc8oXdA3SOWP
ObUNMVMjQX0ngJjpkYwaEy+D5FVQ7VNr8LTZ3XnRnWzfMB/t3bm9VZfqAS1YfuEV
1+kpaxQnY9GeNCdI36xaVnLsNJ1fMM/gQjmHFg8YgS3ToB/9Ka7pQPZB+CjUP4T4
5OWuvGaLDgPJiO+TBkFeLamyge7tu8TWdBh/NuB+K4dXyhjRdwjA2a24sLoO7Ky7
ZMFHjPD1a6q4+OeTalmSigE98StXM33lSKb1OV/akUHjfDFkEz1cfmfV/t+q2BwY
U4g0IZDZ/qmJkoua4fcVj8kWDrU+5X+umk8mMOo6yuthJlQnY9DqeS8C4vCKPhHo
8VgN71uYhMZJtIXJTRyKpD5lfCV+eOCZ7vEVDzVXr9jj3Us0V4a75jOLIQFgxjqa
nOdtwGPVCmKy1lMaSzdlPRIyUovpxcsDL8PVbg6A456USQFuZMvqLGq8tfuHy/EY
wsba8hRr/LCHnVLj1zEjUlTCT6iUoDmJNe7qFS/6jos47TprTeKsIzVyXOdKYUZe
/6HBCPi72U0/R632TDS3IR4sx66hnk6IZgfMiqiLlReij9fMMSjVUFqw+KL5wrGi
YL7vo+4Cjyi5joZIqjodhZIG38Pmb5GYeiCi4ENdkE4mMu0ZelFTRHIdV3ykGo2R
Ct1iAkFo+Ak7IAIiCESIn5JliYZHaFHGsVRj6Nh6oQvhAbsouBqQUgej9Zr+Cu1l
A1EWQ5XSlFEf6jwZfv/AyT/FJqER1gjJ8QbIJvVmDXOzD/nztEbOkr6Ki+gcIWqR
MNmFsrw5MevJ7asn1GcFlqLjMFDkQT+llpXNYYLmVGHuhG1mPJlaAgoEyVAFG7em
q8k8BWBGr0PQujzwqPWC66Y3pxpUqhqBrybbqIEb+mfodribUdGZ4Cr/pFu0Fjez
LjU9WkCUE8/5XgqerP79HTBJ5lWE5cwgBPVqMXGTInT+rVSyel5Y5s09UVOEye0Z
STc6y/AnybcBJWpYudQ3Zn5of7N7OCWvFQcB9AnVCTdqTNdB+jpjKJ/s0gJB2TWK
1vAf7WxkI0+J7MzVKn2XqfSojo9Z+2tgPRDxyrDXXgWwJm9HDo6soaOCViwZjWrg
flaG+JSqXN+X9CmTadckiWmC3sK/tkvG8L2EXyDtd9skbga8zg4X675pBRHw7T+u
f2Mh+EwJL3iFjKymbousPx15nyQqohJ6gVIbUiFUNSPjlfw9/m4MxucpFhpxIpTD
t/om8+hXLIjoq/SceG87DSQSJhu5+9Zervk/ZwzYXzUikxPRTOUkPyk9341e7+ip
d0WNrwWc4kLgrhiffdMTBMuFwrlxf2zIvuNoprcyWFy3pCVcxkYQKXlunIXtNzpp
bjjEH6q0qc2gG5IsIAScc0V4NUTVzARF8WyjT8aNFK5xsIp7VgG47p+p1RA/h/Rc
gkpPRGEHWvWGHPKeW8cBWufB+2Js9YBnGe+EwleffXPdm5ZDJ8VGVRk+oNXKtMXw
LhTDUxHAlasfLyj4xjUetSG8cIDXGHMAF0Hh3JW2lJYyDtDtsQ7AI+ZoIrwb3vNL
eGm3BkQOvzx9VyUTyTiLY8p5BmVCRlbk3FFhsItS3slgdKWDtZWgODI0rhNPNQ8x
dyr+Gn2K7ijk08g0PtcfO/XmEzxMJpm1E5aucvpi8eEHMdxYJEZH5L5YJPrtO8+Q
6rEWOUq9JkFL5C12YMTPot3sqGkt+n3oNZWc/Y/ynSirsjRsIKqLIHFp4GsPc8/J
hYsj8rJyYAip7WMHSY2uoRSbSAnlWyPC79haB1uWfD/Sb89AwB1BtanELiWqMfI5
/LekQNUBT0ZO715pFGcWIxI4Z2cqAqB1ALIsM4KYGoZJZcf24bzUrbIubsQzvZRg
LvpZVKzgPrPzTo0vaUHw+qThKQsuwwSWkkwVAgcCE/Dv2QkKl/yIcP+q7eqyVyPS
6GB6jWWTvsoYeRpU3WvE0eh8OFalsS3wrUIwK33tRAEt1GRy7AOJFss/Z9qN73+C
9QxEZzk8Hi3VGL+Kyle7XYtUWuzcdWU8Y4Fw0kt7jaYMykR7ptTJndEGGDkcDSI2
lbz2iuakvJCIn/HEGV/6ALT6hvz6xGz6QFnputiqHJbTEON6WqbeusYxVvpVLrje
N3VU2/fZP+XyODIwAgUXWtkYHDvKXq53lzSrN1Wp3aHGZtE0N8j83gQvry/xyTIU
BHyVMtsPnVKDtEsFN61r8bx0/mVXnADSe6AB6RFkmAV+LZMiHPq5ygekpVZTmAmH
ys9mUK/zY0hu3xp5vAFZVq04YeL6jxEQtp8wz3OWjCUoBYqOnEglb0a61CPsmhcm
Nj/XSZJ0hVLNhDQm5BrVH9Uk7c1n6ny1o/rJNu/lw4t9hcRz0fjNQ6G3JDfEk5R1
Iu0n8qyETJs2gYj59+CosUjRSXZl25jW8KwpEOVM7pgIu7FKThdrCveL5Bsrsmo/
9GVjqVdDc7Bz3HAY/qpX/1VDxrsEuPiabK41JcSGIQmHT90cRq3sXYuJO5XyNe0b
HpbdDx38VCtZdeJY3SX03mm8DFnT4nqA14vj/uHz7sJQyZBVcF8onI6xzDghrjQa
TAojbCvha036uXowvIjgWaZvJrKTcTp5btYwnbqB0W4OnWM7hpYI7EOt33+eCajw
ryo2H4q2I/BuqYE6SMTr1vOvKP/kfnFvZR/GtDqgqLH6jcer/yO/ZNyuBUEfmh23
ewJ+h+NgARAkCey9uQF7qkajlj7ZzdbvkxuJHvp31iwo+ou2QrS7rr2eyVl0zZFn
2ocXUeQajs3geOum3L/YCfBc+FCX1f3ZBXcU+QBniJzJXU4KxGF0CGjiUUZAQDM1
4Tm9TDR+G0wvKC3eiVJOGjtidk4lgp4nwjI8esDVIDbeBwZUfZt/7ejlduycFWjz
nUKt0ejoP5GvKU3G/NWc6rgeFCSJuFeF7ixODBrNtTxBe0XZEBppYQ2bjrO/+FfJ
lmQ90yqpjk6ojnVEVROiNkTzTWmss6hUpWo6CnKCd3L9hFPlAspTN/HRBEyOWxKM
KvbvhuINJyL/ohTH77NOah61y3EvbpLw7gOfrGjOYJVw1MvxLl1mBOhI/L0wmk1i
dNZq4U1vxMllXJaj8EayYBt31c3fXvaI/5hljzaOZpFwUnYAgiBcW/oSG5y94yIQ
uzJztLeCGIzxEwa1mFiL8YviT2F0L8OEBE61RRk+cLIMpMzKRHyOxuuA6xWBsAJY
coK+x2FsHtGDSxXNhXga6jqyD7cjA3OXLQuyePbIKN+oNdEwwRsImoKH3y0eYIbk
PDtqt1P4ZY2xQBuZardL58OuKTFrW3rfOwip3Kr+Ajgvtp87yXPo5yd2yFdLrVl4
mIT8/UoN84sfDECndUWVzxBS/F5/8XT/YGtbaqf9xbSGKxIUpScSWuEkRvfjUWyD
OoWGCDbE19lM4aTGuuwFAlsvMcJAeIXQ/Fxev39HxKvJ0dnyKbH2Qe0f4oknyVU8
yPWsQazkGZUec/V/HLLjV1h7VZGPY13xYUwqWzrovVpnNBqSAFvLrzd04PClNu+6
THS8r936Beg+2MlGWR5ssBroj9CNrwdGvJkNeBx6NZ0QlA7ZAphehJqos6vP7o2A
ehoWoIhVrgAVAtIBSpCwqUTBwElYCmrtKXYqlyVfRY/quZqbKoY1buWvIOMc3hH8
WD3KV8jC2WqrTVeAGyISwLlW+sEml3UcDPHJmi0S/gZuZxrDRpWMYX0WszW3QvGg
8sNU9KTFjgBfDXd5iutIrC9ImN4eCy22oW6NPG10Sie/Ur2ntEnjdlZ2vFxJz4X1
thdtZ21H1ggeDhlB5fh0lfwH3M4NHunDtvjSDy4Mne1JS8Rzu99ehYHpscVBV+Rs
i+Cf9cFSF+647vABlEiXDLeV2GAQ3Yvo5lshjuLJLuY/mqWbsw1QUiLThlyVn9vV
L3j2e5VRNXGmQIMXReZsqhBBE77JSUy/RtXvnOhIbfr9V/C9xcaEHjKi2mEYRRh4
aMCYLQYNvu4GTegNj3AH8mekznEPHSTA8hp+B/278D1jblW2mcNmrIJP3vhPKMaP
PQYOshJp6HWr+zaheSC68dRrrEKE4ahFDn1xktj3jmcdi9EY9BvFDZXausraXEPq
7VMDKRHDHr/8M2kzyV0hBc9l+vXP1hXeKXsEOV1gAhl3PJ63zXy/PWqtxFj52wiR
sm76LlCZL6ME9Kn7zstRVUFe+aMtYsBhk1Da+nZ5iRJ1fUMT532J18lRpU6WSl6d
yTgMfBHczGJjlylZ1KolDqYiA5iDG6UlD5neY/27T0siD1FMSd8FV7NouFjy5s9+
EI2z3rFmAVRg+xYK0pgEdCAcaA/YJAMzaNyUy5OHqy6ZVSP+cdlGLOW25uACB2g4
Hb4PD8i4+B7v+JMmJD600mNx3VDhiFxUIzMFdqCgrJyamIQX77frk4wcjawHBsph
fjrcQof8lbLAN1xQZLloX8aoB3xleijru0Z06RwZsGoPfanMdExXpKAxeXXF8qOw
mlfd5CIiA8BJzMJcApk0e9i+iLh0R65ymJ3VtxCdPicx7f/CEiSLv6AYKfdsYADW
JtH4Y1Fd9lbC1WyJ+E8M+zn2bqBDrezMiGTKAoHf1r2ABnEtTWE/1dnO4g+yadz/
Ht05VKIqH3AGGokFS0tfBYJK0cPor2oT2vyrg1kTur5zGCes/KB7bQz1G1cwIXzF
kUz++U2HTc526FIpKtFkOoa/9qxRipjnvmUvyDy5l445HdsPEC4QgBrUiPNumoVM
u4cxQ9xG45sgI/ooJdaRA7tBiH0Sgi42Wmrd88HtzTp1IpJNpzfMd9KZ4aY9SaRi
yjlNnE+IJAlU2d5Gj/GG0I3CNqC4Danhjf0dxUHRp28hTpcaaIWvq0aezkg44Oaw
aXwIznyxrUR7GpRk06lYQlPV1NafbcWo+blsgdFtBrXRpJRxu8LsHrAA2Zbgi51R
3/cGsyi+ZqMa1BKXjdxvNuA3zeZ6WHTQV2YObGmKFG+4EVEV6qLmCxLxJ6jPxqkw
vteRvpKgMPlc+ea1+ACEp3L645xJ7rz7Db68cBmcwrtZCd60xxcC28tBGhW4pLP6
2VAhKA2EYGqi/d/Fo8HG9jzVul0lBS/hb6V5OWbkfuZB3i+WoBPSUfdzO/xz2E4d
AlF9CYL+vVx7ApAmVAwobVMZp59VmuxQ1vIbIwN4Vj2BZJAWCrX6DPX26Vsm56lx
d/NEymXceVjtF9nhDyo0y4EAmYOuLNET7MwlyQmLwFhMSjlyJgdMN5ldoWMYoDMJ
Fnj0fjn2/d2lZaVlc0doVQ2Vf1AAeE/ZkaQoAIVIshVvRvDTs11rvrqMKrG3f91N
BV6OPZ2D6Mwv9P89s2tX/6JbOU9mZs5TxfhKkC45oXgy7HOXFpD1feHWjIDVl+gv
pysEclf+RSbzUPb76JQMXoQdlJPP3wYYtJNm5JYwAP3zdXFmub2IQJkeLcg0g1Ld
iXO937JcbZyk//9pOuBbHnZXRNOFgGAvu5J8kMVhcz1gne3vGJbw2INugrvgYgDb
jGjFSe21Tgw1JJhpOOipTZQLRTX+dcNuhJ+LPtNFZm7D7ONTZsUwtZG1BEjM1FBx
RnTF+mipAm8BbPB2C0HbdQz083J1ACh6H96HTsf9NiWvfzntO82sY+d5Asf05F3f
fWkVtzG4ySrVp6nML69m0VeYsaEg0qbxiH5qAMNFkkXqO8PmKQRrZnTzoTDtfR2d
wIQjgydzF7QZxUL7C1C6bf09akW1RM2buq4QM+Qzvf5l2psoAWzrN7r222gbgqge
txxMzP1WlYfkpIDh4S7LahVoYuXAAoB0PtpVZbb9HrlfFNM2oyGWaTi6FZmJhzSf
Tnp3/OJk0RpXV4MkIl7c1vqY2aa4qBbyENp8cvFZuM2//h/kjqqaqbms7NPNffMo
eMGj55gB3zMnwKmgjj/HFfj6PCEx2jvnuu7S182NObw8DXZwM3w5FdUL8ahm04wV
m/gxP6HtGe1LvQtUyFuxVfDjGemoxhf1CusW6AGeu8c6fVhQMqKgvOlUhsC5BM1c
3dSm4Pc0LtM4pg3uG0eSOo+xdptJPCG5d8RVFyBK0LXHYWrBK/MheYLH9y9LN8D0
evnLyveGw/bcuEIPTkAKtPivJe7F1wq4nHEFHOmj+qZKHjIEZXPFvVSA3lKyN5Dt
5jcdZ+68Sl1+sd1GIzTVVNV2YHqA7Ie/b+K+CKDXNBYnE2RKDwJJvXfigr4/9c+R
tdBjUWI5SavxZ3wB2MdJBREqMbhh/8/9RplDTe3uhjRRuHNj3yl61eng4/S+kgFt
jjIws2UUftgjBWc0P2ATgCcILqs+WYy7sOXcvphM6OsHQvHf8jGwW+BsJCCO4Gfs
I87Sywrd7MIEcsU6mPfBrsd/2YXgvYXXDUiYqeaLtZD6GPKx2jzGo8X7AQu6/rFn
zlsZOpVkb7RtKfnjSVso7ejFj4vgMMYmw8Ime5foKQs/ddoWT0LwUanGzWFFl37Q
31Hh66RIKR1a6oLvxNSCC36ld6Crr9Rv4yGNQVXB+DHTovpuJCQJ8VkaIEQ3Gs8O
Lp7kZkhhSZgfC83me6zGOZUgazwDyyo29S3CVxjoP9qbA+U0OdNq8g+mkKu6FDAX
fZdetejFIxd8+tlsiOwZeFvUUa3gl3/5SXsyj8OqiuVYeoSrG0WcJ470Th2n8gc1
d+JtC/e//qvCm/zHHdlQ/qlPwIEVxud/vu/jRR/Il0AdH+zrJ/Vcp+hsHLfqYamK
Yb97UckDgSu+pNIxqwNyii6FbpyrFgbu/N6S1MjXR13z1+QCrNM9LnTLTGuUpkNa
22H9kBNHPnMH/hCYjdn9ZdcG7w6ut+sSHslmV2h4Cbv45hUsgWvtrnp7U9szu2li
0WMBnCIzzXYtFVeCffPJMF/K8nw9zR94RZJi1Gow8qtEN8hZqxAmaIx847Yf6SCo
sHQYHgE91pBXl001EaovGgIQDJj8uctk7XCtv5kU1UAhZSy3b67cL1tHk/xoUgUH
9vGXU7PZWxcg/YordmNAvj7xbC46R9VUquzZrxHNuTiAIJdqZ5zDKcUh4gXv/kE1
WO62SSKvg5sP4WUv7HJZVpZICHLaLXJq+c8m9mrYyMYqjNSPt+ktJDDuLnEwXogP
F08NCoVqCubPRDFZxZc3FOYy+dagaWdRZvaOcGTJPjuy0QxWzADi2s4YbZXhxu69
WhBcGmOUjDJtb8PmupDXjQzDR//mdjSxcfyJd1Puxrl2v/uNnqa/D64yJYJnvul+
xa6s/tTQf97OndjUoeK+LZWq6sEybSZktwGnjPMtREBQjaQUJeO2JQW9WLOHxcJR
ANiwXop6R/IjzGnlX1Cq0QDxaupDTCZs3xkHzxQ3eQrI7ecNlLgPKttNeTbwNlQj
FyNbVfbUIrY2jYJ+nFFrGKDM8O+774x2PZI6vVltYqF9dQ/Hvn5i3t0vtmyXXax6
a3Na2JJj8LHtRbkS6iWtT8ua5zlD8v//JrXtAlT9hV6pRDf55ci+bmUgYqSWrsa+
g0xB5/RGBxsf8CZCYrrMfViMp4FJbtOhL0AmiQ6lQIvM4p+nGRqm8Y/eo1ox7PZE
YGA0zMh6XwpYh/UnsmXgRc2rBg3SCNss+ZMahPH3yrLl6d1LCRTXaOEeRRksWixL
hCcSgkFnoscgGMTGFJ3z+QmPcW3q0EfGMVjmzNLwlKccLp2haAV1EjG/NnXt1nhM
HFrd0iL8RhGH6/4CqxnQQl5XQaOdb6wJQpHWbEkUUen2/mrTc9PBjUf7PcMMdpIr
Tb0nHDCZD7kSJu764MzNdhgNl4IzcBhYW0sNjxyczXghrgE+AP1KN/KLS/71adbR
NcqQqcJJUamX02Gsd3wz1RYUJEG+jV27lPhH1EXvV9NDk848tXn8/TchrFX3nwKp
M7dooox0pT3s8gNccHXJd6+WJ12cQ3DPz+OTy7ou5WPm9+QrUNVmDn/kwIRuDE5N
p6wO3VqI5naunkf/9HJX0Xcvf4NSPm4wbl0mzf+JIRx5F8z5sEj1xSgAg2TXmLBG
H4UBIUyx1KnbXoigRD9Y7na/8q2cI+RUTCpCYWAGWLbwCqT62E/iR1ulOlx6UcXK
CcV6OBUpOnZ1iIB44VpQA674UztC+P80PgxHnKuidwfSyyp0O57Xr4xsNJjpr4Wp
0lOMGW6E5sBdwmUVphO5WGszhSGOZGzJEQauZGz7QdpUKvecUyHawzQ6t0NqH8K7
Xzty99mEmICRFWJxVhAhttJx8cwn8dVtMks5zxC9gWF+EZcqcaO0ISTCzVRG3kqa
IrqzcKSEG7JFrbyhHpTYKHxTFyZTK31vZNxDpdH+Larc5Gvgm44S0TcMU+d8m7nm
slz3MrboL4AFJl3nK9ND/X4ulFyrYVRHeJEkVJZxyKa8cZGo2vXna3nFeVOxluAI
Q1lRxk5wYW/HZVIEyHsy+cPMPXPDqft9XkQS5yuEhiPNPmXsB+MJp/ec6HL9NOkI
F4GkPmojVQCtXYg0ehIW4n1iytSk5LTAui6DwKr6BCOL73kJKyyJp34QdqzKKoi6
fQzq5y/fuhahpjXrrITTjT2ok3MZNyZd//IY7Ac+xGvYs55wSr7kq+Dv7OgotM2X
Gvxu61532LiMJtYgiQTMgiTzIwkuNzvKoXDlQ7rV4r9kYaTAmW3L1Al2ITS5MHi9
lB+XhC1tNLHa4aVznTdMydzkP50m/cH6LQCm7RVZX7I4kEOzSoddteNd7UzGsYYb
6P2twqHmsqPmxNR8RDm6RFJhBzGlPE7/v2gOdi7yEKBaZif9iLIc0LwHByuzD5z0
A/pBldSUv9JxyjZOOTYToSpGDg/c/eaRwT0AKID7ZN2U31jg7cv8klg9NezT3+wf
egTFphY62Fkggd5XBtRWBWg21UPEt9ZcHw+gESB+7SIlEMskEKAcyFVeI9lu07uF
AGGNe36cda0flw/HpuWz0NYlzULvTNEeWc/ntZ7bWppo8U5fzkklFd18tyEen+8A
4QzGQirzdkFvVxs1vaYBU0dwZNoWoaXNBOEyvqcXoWi3OvAKRe2q6Ii46jI77DPu
nxRvf9kogC9otMOXCkIGqc3odXnKhHOZrZXA6VX9n6LupsuRZvrWgkKuJuBr5Hru
VDmnnMaRucMiJS5ImrNaMelB327cycdUFEHxdKbPgW285otRCUO+Zsjc6YT93r3d
wb1rUXzO5V8WM3A0jS0FvP9h+MSxtdNFiZU9BEBIYAiR8xFh/kVyuaK7FMrZNQn7
3wgDEGA74zJv+xHrtqAtua5mfOxuUevkpmYAz1nNGHbLO0EgzdKBosswgohtLBOa
ZHlVwMOhKNOGIv70ltmoP0bKJ9ZAWVUlLcoLzjK89i+MjIvOhuJe8AeMwXClHcMN
Rt0iCM+WDPj99OGRkM15LNhnxtt9fhC4Qg4PO56C3/L/5mRExF8KgtI1RnUAAAGM
KumRgX3Z7SjqlTrkhz4s+ZT5pyzJZfHvyDZBklToBxFcnHTH3IPEkZC8pob6oEQt
2REcS/wgdGqi9MmOesL3elRSetqqqURMZjn3hjnJAme4n8PiIMHhVCHuokwyumh9
37B2FA53XnjS2p7AZW5qnCZWBfHAOxUAzAdGRJPIdaTUd7Fy0mH6/1EiZt8o9Jn/
07LyZKXczXEepWqNbLhs9UZvrQeScKN/1NkaBUL4KtdIzlfaYiY56AgEqrcLqfHp
I2s4eYW46nQcJAcjQTA2SVpBeKSH0y1Fx951/eFFG29OuviEQzpKBvppom5OtbB2
XcoIBFSVU+UgHoqFKT6v8I3zttMPxVKIobEha6QUqYxG4BSsdrEM0WBeMUcv8FKF
e9L02LfheyVYlWdGFUvbFyBZ6dKTk9QTz+axWpUe5xhN9HXVhEkOtXQB8ik9+oJX
7y+iOjuF3Fk1UqcH93U4tLY6NSZwJIQV1KrC7iDAJM+cG0jPm+fV8Hjm2qXhtB1Z
p+idgdNA1lgbTh0QGhOKesYZPm+BHlgWAW0iICa/GCtTf+7PTlfW2ayEkahSEFXZ
KRGqJUg/Is+IVSutzqduNaCcoW5lz/WxXe5AVE/xDMO9/NyqvhtOZjfxj85jgvc9
Mtel4NnbZ+kvXY3r0fm1xeTVyMlINnL/job7ZbxtWZo5ZUNz2mBL2h2VMCt9B4yp
DNnUyc9T6F0HeuqZZvPpXeCrNjfUpXfDG1uL1PHkxY2JGV9Zew99hEumlttHURKG
/9jHHYLAOZ64MaKWD4l1wwdwBCMy8yl6RLobw5+PWj/YeOsf/EqGhTrId/47v/yj
fR4aFhuGHoWLAEDO+1BpBmwKn0RkfAOtjTNzL5wawNjChuoGCiLbGXMKp8tgkAyc
sh7GCpK5ab9k+q8izByhh3ZPnzbQb+xqahG5M41Yy+IdOIaSgT4x/WKhNqBbITRT
xZoVexQ2xSTKEVzukI56i4qZVyJikKhAPzWODm2s3RNeovmS/SdKgdVeCOFs4mWV
pS8vBOzp4kXojAEBOwu+iOLvkGJSciO+7/4CXkOLi0CsIa6VdtpKn7c37fBChJPb
l3/GdVgkEgONPprSDH12xJpQmBemO26tZgp5xT3joq2+I/CSTEKwS7ISX8R+d+9m
8NjQNAivdPJspuG8X22Bk2pHmpdbvtrcaEphmU2uNOk7mdbyjtQ98S7hoG/VqUIs
1tDHSM13U7ofbKCtdZNwF07XR6ZsHmxfhgV16MAh7RF19tHSkYWYuWJQeKi80Tik
QzrO/HCrwYk61/wbI4Pl/nIhzB69BBMy0eiehkD0vb5YwPmVe3kNhCSX/dF3WnIl
EWa4y6q3KKOKO8Y1jTQ0YyNoj++Ur4MNybrTWb2S7aOEILvyD8H/8xtpXUaGbiPt
uaH+v/q7WNrr+NpnOM7ikvXHvetBP0hPh1n3swaPwkqEw7bmxHQ19TGpuSDO4nQX
+N8MzyzbnkdO5CVkemTJJ2ds8jv2gmJd+JBap+3zyIQGmLOUFGpYkItG4H/pjY6G
yitFhVTWFIkezIx2hBqLPczLswoga/ZNup3eDSgGHLPwm+Axz4VWdIBHSM5cAmc2
WI/fTKDwBkjHQ+vdNUzDD3TUh3rVROHWEaMRsj7f8qtP0ny1nipHwQGzl+OlFUnF
tuCq7iki5sb0oSlIYEiGJ8/Id5vgd+UdNZ23Tzamz3oKFWdEz07C1BFsW3ZX0Y1C
LpfGogm74DvzpEoACr4CyBlXKhJnMdJB9OHqb0d5mtCqtmUjkc//xn8uG8rbQ8Fg
CWJDazfdelm9KgSQkUH+f6QfNaI1SJfMni8dqMvL61G/tBQPURmiDjoeM17/9gg+
tHrVs4bIJvfdP77lsElMhMD2dRH19Wm6evG9J3Rj1YjgvRRkcPGRRyzahVejhtvC
ZjLmsbzpjagW2rvQPRNG0cEzAZuf1oAKRkc7P+RcCzh8Ogp06/zGuw+00Y6wX00D
Vv8HNp4bdvQ2iUgaWw7ZBBNOk5vpikh/9in6QmUDpiCIgz9AYFB1zFFHi7TpyRO3
52rME+go+le+V93nEUb259KZ/yknn4NyhXurVhPYl/l6l4UTY/I6Wv0UA8GAq9jH
PnEaUsFBNPexzz1E9A17dAG+y7iIRwPv6s5QUEvYMmdOdLiPv8z/vbXUlsBrZSZf
zHw4/aXjPskG/b4y9H1ghBQS6vw1HT8THlUBIqXP5yjAcuBtZ6QvOLnNN2eogJes
tAoZyaIXPlRJMcPvQuAgvpl6ugC/JmAQD/+V/itLDZIiI89g8B5qNZBxOkW2Qir8
uA1GdQeJRnLg+h8YkaS2LY8PvE/a0BG5AH5wKsnR8358KdNtjtvFSlbyLDf7zCA2
ZofWB8gnN2w80FEuK/2vo3PdZXtAsvQ7Xndr4fkJeenMObwNs0ZEHi/7fJsSNFJv
O9OC7h2IJPHW6SiNFtiZ+Yl8cTPCe5DnezGL/hB8J9iGc1ildLb944ZIlLUsVyBf
tJP7mSDoGvjAnT9Z5gfE2EeVhhnvOlTGgr3c7hfy6AclNoWJXeqBxeOpHXoPeW7p
wvaycx7FZ2NfB+Qfuwyjkob0itOFXIo5kBK6ihiUXeWtT6lLTrKXAk/tkRqqcpRV
Y1WSPxYk0fibJlBEFSDmYvueCMNxLMWO+WJFvFPktBxqM3nuPhIm04ipLqfHblq/
ZcxvjRr61/IXxD2H76+ORIeBSVlqvsjH4V0+jmeXoNYDVF1BU4zlKRYvGaf3YGbR
rsqg5aDKMuUBIIvvOp1BzM6FjpINCyE8YTdnqnP80uuzvN38Bwq6wGTYhZGyQg5s
f5n5WNmcIMLGi8duL855lbiH0yLDv6ubzTpmU37SXM5R1Luxxs1KyI19x2G7CRfv
6ohBguVBvJg9z8K53RaVcbxH5g34RiYJJhcSXLvp18Z4Kt7F2Z3THk7bE2S7q7Jy
1yWYSNm9mNiGgBsgqiro03u2PJT2NGV2cGUJoeGaUPNWL1fQ2QsUfp9BQ+4EuUq0
OdzInuKvOuh2j9dSGEk272/6jhVzEppD6fUv33oMy6V8Q2t8oO/IMRJ4BEo8pqT5
2vtV90MEiQIrZYG/f+Cu4JO51TEeZc98YrzNF3sPgXc47vjTZXk28GMwxV2UZW3z
KDIxCtjdcafLgtrxvt6isOgbH2l7+oc9JTjgLDuj+zNw9ERKdX/G4YHFl0VxMJ7a
ZCIRddhMQjLaOjhUQX6kn/ggTPpg9Kv1y4r4YzT8GRrXx6CRtMSAOGNtPCnUcFfu
d8Pp5BONnSLv4dXixOqSTfv4flDSrd34Mul4kd96iFnzRffnHRhTnCmFfsLbt/9M
FPlpdssFwIK3jYfghj5qBf+pZC70CORLwPhjFfnMY+iNQKsBAyw0O8pw2zmHF1rC
KxvBzSGXC1SPVkKp3Em+iOBUAUCxmSxdVUXmUgC/o8AeU7X0W67CJmqI/QfILkS6
7+taT4j0GKmrp17JO6T9Q45s0ySDPT0XmZYjhdZ3WFc99U8saqEFQEq8P8gzMg6P
ByBwnlYHW5kgPd7LqxFGjZI9D30mrrtUxo/ybAe52HvVYFweaESShJ72122pG5wr
0d/VnKFYjWDT3GibcsDaEEajV2HhMEat632E0TxPWu2HF/E1WIcChw2TsBrHzk8B
/pmra99Y4LgCceBAtK0dR5GnAlvdvDgPStIE/I4Cmq3aiCRo4A/1k0D1MvP0OFKt
aUUXcXNcoX4VksEd0Ia5pqxVC5q9RpxJ9eB2fnOVj3inuIAAOF4ujJc6KkiMnwYX
LvInh2A4sPme1qsJP2Q++wB2GsWzyoVbK63SzUQqhOhE8Eb4ncDRHJGqTTXCou3r
SSUhZyBmLIzflZ1/8/icAImmLOUMRh/gh0Aa58Hgz1QhTEoHxuK5Mm4UhnTOoQ+C
DjSMVwohAwNJiqHsEjECYrj+nueODXjhVbP6cJ5wM2Gprf+kHWDh93QRXvYP91a1
K9J2L5yXfz6Z6kL94jfRpp8E4dMZQPppe1nzTx1LZdZ1JJaTBIi6It5yD5YXodL5
pT6Nvho5BAcFojFcBhwa6qJDKfwFqEGPXknpojNpOd3wqf/oIu0+DpSjzJVEU5XK
N6VcztviGj33h5wue6jF4NWAbg9gBtEg9AeYHEFpCt8lLniEDO8f4wI0ROwqu6Ni
aPzFw/DZL53v8XMaavgdyhQyxOj05nGVmtNNgoxIMh1H6Nvenf5JwI3wFF3i6GHu
Z5OnR697VZe9XK22hBpoQGovlkJvaWx4E5hRcTI1o/Dk/2xETAsLRsp1mLgNO7YT
ywU2hHgDbLvUFwh4LwvZP1TL1zz3oxCvev+J+GmYSWCK7/MXwwiLom0ofZLAWfY1
mJpM+GiImI8CqsA+jAPG1pfhmY7A+tx2GIsX5X1b0YGxagvl+5FMLL4KvYwDNdp5
t6QeDrJRLZtf9dcIS7B2vI4SXTzZylmIVd1WqA/FS5f2ra6eAuIDqpaLED4hCdmW
pLkj4BKNEVVQ87h1tJ5qWFxdLTv4JujP0Se0W7vkPPZweIMbFhqyfUuNt8cTyQMZ
GA0AofGusNkYmrV8A5cd4JPIIcxwSFLY1eK+/3Tt/tH5P+vnsVu/67TwfEAIcEby
2UbPvCK3PoatNjMtlje8uaOMEgnAPoDi/VvCNo3YM4GRJqH1cWqGZReEu1pci2vF
gIZWgcitOJbcYh12j/0w+f2ooMciukq7vqpdxOQzbXxr66X+ouNCdB3h290ZAZBM
DoJk8qo+N3c6Gv6eaS7vAusV6A6BA+A7TVjqzC7MQrpJRxUD43fGq+tmRDNFxoWZ
K7oZmhPBaRW1StJHylls+Ub7TjaxE9anCjQz21lc0UBKKqC5F0celeVNqw7SM2G6
Ckon6NG43NUu4j3zLqu4oNGJ/8IaFNrEVEpVgWSOZIgUt0r/vDP1DQquZknAdcA+
jxZ5XkvntFgqEKqpVXm5QafKxnWb2cf0K4ZZ//Z0WLtaaXxL2ZQXeixOEDgYjbg+
AbS9HpZv4XQMVAj9ChWaWayZRx7t1XVZQVYAJ7PEYA4npCAA2XmdvzU+mVhcFe/I
CNpoeoTBFNfz8ESj6OOlGsjs7VPePgpZTiazPPLJFXs9RmDLsjejMfa3UqgSxY71
6pO33fgN2dvnFS4CrkTsFnaMU6/ZqLdTWx42t+EkKqVY1eoAC4GtiRzeTRYGNCxf
So2jruusE13WinmH/0cEEbEFsoIp07JBcR0UqEmFzMvyJ5Mkgq0BrmgR6GOAlSwy
To+g8L1S4Dy4pPSVmHXCkpIcViTbyWJ3VWQVaYW2XgmXqglw8iBBxm50wi26cJPq
LqYOV/n5xx5xu8oqN9dLIiWd8egyHFJtmic7cIHNnnYKyLvXpzO8FVE+fqM1TC5g
Cul89KbnTtSxkuCbbvhZvT1NRzlnJ9cOLzppOzUr64NnJgJzGIogD031bmKpNkKw
+AayHEP4kvZP3O5nj/Uvl9Jvd2PctS3rNVlKzekXZK1Rvh5hMq0thPuUT6FXK+k4
Cnntmx02nYLuo5G2pkAXu7ozdC9bsFaowUdWvWuZBP4npH9YrWYJE4QeTz08eA8r
MHlR367t1z+ZesdDFKXnTp/4EvE66rJQRo/bGln8zyKo0UOku6LcYmLpS7qTzF1i
keHwhUdD/rOMDNBis1tBQwKWTZ/HcC9aWJgEN6AjFVOetg+5HoM76bMqX5llEqk1
7B7j1FGig4cQI1xaRewHMIEXCLWRMdmeM46DQmsp4k9ZKCWqw/fQ/2GW5bbHhFqg
BFXK58m9O/29ECnaKf0udoFvUCW699Nu/fr/GxMY3N48ZTn6rIdujrFxyJa6Qqou
e5gS2rtzmXxyaAmkuFJjla7ETM/+OLCn05vLTGNi1cCZFqwzJbzm++bVceZfYYLa
QSLm18S7dGMZxnPaLKtYHH9KsEe7odX+BO70z4T8e2N4kGIcQCjfKcT1OyUTrF8m
ZOtJAeNiDMf5f77+GkJAAVz26rV9iO/KVyQ4pPqq7Ex3lGOPktT615idWkpVbdFl
eN45ZneL2eqWzWRDEa0a3fxHNdcb6fJL4UtQ9+oNb4k2TySjjhD4kxjD9ZOiNp0c
lYpH3RCBLXov0Xq0tA+et31G5Gzi+xrNHcDrZWIk80swJzW/d2JVtZRvHoV/Gw6F
xiLyNnV6AOCdPtG9wff8iuM99hVHyIYKy58lVRMsX8Xhrx0BikwuHgHi1UD4n1Zv
S/dub8BbQfBQQeXoota3yIlpc0M98E62FyFq8ahPrSLoz8tlLMM/8436BzqSKaXD
pZYEmExXXeDXDzpdl7ri+9yP3yTGhYsLOy2bGscXFARJ2jbJ2XROOs9hhsO0tWbu
ErGnxt6wXjrONgOyVuvDwgw4PZUcaUm2DL9iT93d4nmMRuLP6+KGDdZfQZ+phgLr
8OrWLE2v+9fCZYLL1aancqFMa4tQgeOY2J+kK5MkZh+3TW5z/TSYOJPN5MZqr+i6
pjpy21cHJ8HjWRQDoNXOd5zpgCbW4YroXtKt7rtzGAFPWBpGoQGGoyy8hqrN/R1C
MBRsYFQGZVnrs2A6fEjNTsSYr8qiciMbHDaToZox8Z6eHvQI/RtSK7UTyzelIonF
pk9JnOSz7LlimKlImgMzRgY0+DhSqUwuw6se5z7rK6uKRCeG9nl1Gw00fPGwI1Cc
y3xi4bq4D4Fm7B3XYKo4g7B6e3q246sKks3iw/v4h3jzTFtTgb3Pgc1Y7TQtWxAT
/UqryQiGdmCuOmUyXIVhxAtUFLqWKDQcCjS/bXunjNmLeoR3n8d41dWDQWRm95ip
+eOhbPTs/B+Ee/CkXSV4G77UgD9kRZnO8BeoaABr9gY2Ido5SmgpHZTIl/rbNtHh
+YXf2H07doePub0zXfeE4uqX0bktZbwHCnvKQCk8ZXTO+WkQ93NOgYH5MvpCcDQY
eLaNrvPBv54W1f+47rPsXYPr1fy1IlUpy8j55udAgkn86GBsFEycp+fifoyOj/hq
Pf8lJHqgpUaebAv+jxr1d/UDqEfFXVuPrRaJ6Cdbl+scGKqF6He4x1sZWRhjpEGg
mv5IzKet3z/5uz15f5dFVbLfu0fzJbwahIa+rv3fIcF1vRjXprbrZHC7tq5W/87t
VYEr5L/yCAyjU58mBtccDbnPV+PoH8JdP3OCi1nC8a4LKlRBG8qeG+BkDI81srwE
1nPuPwE4k3QiKJlOOKNOezGDJnLrb+C1I1Uwas/jZnOILjcQPgdqUGMp37ziwpZP
xDIUvNCm2JXPeViBPDj0CxIDYRZ2J0QSTxOrDrLqrLj/XmmvEtg0DPVKR89vExpq
2tp93Gb5d6x0f09u72mi/9oAyC9kHoHsx3QjTENUlIZ3Z/vdYRHXfMmU3R8C7U0t
CQgKzeVPmKd5U1dMAd+Qkjuus42fP7RjKI0SX/AA7Ownngnuqa5brdC22AEc0VOE
0rFH/uD6ZMLm7u0X5BtEyRRfhp/2U5OVMcLGXDaFodbm8sLarrqGscTTZXlQo+XC
LWmHd0ZGCmdvO4iyv/4UsgXAqtl2SeslSmG0wehhgSkhxToXhZEYqkMKfAWELnF9
7gg9FZA4X3FQ+M5oBGLBLnD8XCFfpkpCZt/LOfJq+nOyOpw5/1eNvIfCBT3/4dfL
sTEfy10h7b/R4uRdzId7En1g2c3LfjtoLHHYlT75reKC9a1Z6ThtylHnD3nQQORr
o+hmLKkPQ+oAiNbDNBfSDzhfcSgLTb11tFxcjBLcTjF0nKYTuBDMWkI5J2jfO1rn
TTUDGKNVc5QQYBcBOO2cEzbTo/OVA6yVWwwpgc5NfHUuFb+48lKstLKGXX/0f8AU
zrK/AS9JPmOlOpcPS62WGDhZlXWy+u/IbQp14+nu7E2oJbQkt+RdPJuajYwvF84d
LARN/haCSRRXXtqJKj9skLamjqa5F0/zDX/3rKTubxKwUPchDBecGcRLjj4jTC0j
Q/Ygyp2zS7dIjC/fYwmIDgtSfaeK7Vwm/lfD/Tz7N+UaX6U0Qd+K5R7PGFWta5ve
YdGRAnmeRt15zruDIrq/PSRTZJsRwDlsPiMrjL9zjhl5IoxzFkSY8MmCWUdZPLKA
m8t9imBlOYxZpSYvg7qMllELW6hvrqQmKzf4RWvBdynbLwMHxMQvIamS1f6n9VyI
9smEwlAj68MsQ0uAeCc6qLQImBYAhS8R5L0nEocbVocEdNnI3uHtfh4bF7TqBThy
wuuLNp1HqxlbI9aKc2jpV/hLFDohxu8HM/soOIrsPBS+zQb38Ra2I8hFwnBn6xul
yhmTDqrMTX7N+FcT2b8RW6EuQweGVhsHu5KGu0Y2tu50yBWHWNg0rZImsmB3A/MV
cWE3a6OemCVE6bzrQD4GcCH8hkiC0Pe2QSFzo0z82LAQCax+i8M+EDLIK7b3RMve
qjktdVKApNMsN1Lf/9Zi5nYUABOWZCIfLbxukcOQHiCKqGE0li7BhhJT2IVireos
4SFWykCG8Ly4y/jqZEyuFrm/8fZRjD/GeAfDBerbDpl9ldu0qPksXoJB/9FgZDin
1SjRQknyHJbK+gnVjWQUvdJhn+XiyL/oqDnFI0/tjN7wuGnWjt/47jBB2tLDErsC
i35Y2YEPHT04nel+clJswqzrcTPyf6p+hFuxwunAV0ziZZ7JHExnLu/GM3mf0drc
adRn9Y3Y6ERPiZlmCrBRO6dZysC2MI0UnDhR2r8IaoxPBdd6HQcNAKmuK3WMSHGH
qWgO798fh0tk4CYU8UmJKFOO/j769ZkSv5ArJeOxzPtIjJfjwIKxoNjcVP528XAZ
4D2BRQjN6TH1GHJm7RwoCl3D8nu7HmnmU/Ppql0hWHxnPxbgWesMsqVJ0Homo77k
vQrHVGTCOp/LPQlQ+20PHu+0yNifK9mF5L322dPbpola+z/mURZw3IdfpIr5PTYa
Jb3bZUBjA/P5UPd3jgddWULwJ1QUBxatuFt3pR+/btBxMZ9pXYCOiOqkBFtwAJM/
6gfj448nrfxK66MoO+xSpLOfUxCel2wXhhz1PZyoy1hr+dd8ZgW34ljCzca3jucm
gM30hb0xiFqkh/bJi5Op5y/YPEroWxzsOwK/3Ej/xPm7tHLTN1aB+fmqS5CFcr7C
yLKbolYDs24fl4zYIKFt/W5riLyU88POAaUja4SnV19EpKNDgiyhpG2TcbEfk8TP
tvhoNVr0dJNBnpA0NOqw6IsNp2g2fPeD+C+ehSIBspeKFeApLUHfGEnPVAzcCjK0
+FUem77OybCConR10GIwy+6Lwpkht8OLnxl/J3ItvxoGSh7l90PHtLlnufpiwCxl
hmNYN0J8DIgqpWeoSLdkRNbQijJQokbNLg73QmzCWaxmBDgc1NZNK9cG3JIVf3y6
EKiPy/eVOaH3LeMqMmq6bnGDLJstHexxX/qAJCzcB/BXo9tNOZjc0pofEOR7QjfV
xNtZqm7eIxE3aj7QHiCHi5J5/EvUHOPdLrZm9WczXuEJKPE8SQBbG5CFvYOJ7sD/
jCdyBkR5lBy5BAvzJHImbz5rBNhtux/XxltZGR6fGf8SrEK2vPIoq1YzwTKB0lxZ
5asYnFbBZt0WVVPvIsRlXxTo5YGEm588Rp8xkbNMXknXzRlGXLdQ3/Wkz52rhCDP
//sZZsnYx7NTF1iTTj/2MLrygaV8vkTFX1VHCHhBgOLI22fJmYwPuSp2VGYaTz3x
UCPdfEJPWhzc/4naDR5iEeewRe0NJd108Gnyr97Ds30wAK/8YJOUODHl6KmkOaIf
4UcKTQwe21jmjcCqLgZM7ra78HB4yhjWm0CxVHesbaOm2onoaqBArtx7k4os05Pk
JpkKTNI7TmiXFm1HoVt4uwLdopcl3d2Di05hREUaYDx8JgVUwndh8WA31WTx80Vs
LoOsRVeX0fmtFAQKcylVxFyrbDsJuO70htwCPEiCzdi1rfPbqpcolsSt+bH0BWOA
WtOYOU/HA3l+L0ChhSRTH2njhWHQ0lE71WKE+B+nHBHanR9MA2wr2C830Ajbt2na
Up/sz5sDv42yCxG/ab5NPjryGfLaW3oDcNtGn2W4aZ0bFEifTOR6egy9a+B+SjHT
cDlif5+F0oFyWTEnWswFTn9izSjAMz/Wo4JVSO6/fvRt9hWxIRTopZSmi232GG23
lcs2vHTAXbt4hTpEO3+vbj/3D66lPbc3IUObv+MI0zC3gzOdajT0ixoeMBcz0LBA
dAWMNIldw3LIn/BiiImjzP2Fqx3zfxcNjVWirWuDay7ouHHcs9XToXeKc4ujpsAQ
P9zwNv79uCqC8+cFJ1il3IAB35ukzihY+/VLehCXJ0/IwGonTZhHRTh2EkwRsKZ+
khR6aZpYrK+Tt1Sn6ql/vQHLDIHVLzBfGEkJ4kSL7w7wd4ivBShnpULZPq/wUFy0
ueikTvbSye/Xla+75jzSid0ZS2L71j/jC4t5usNP4tZDsz4IQDu1TInexUlQ3p85
wUp7UCaf9CAWg75RzeDt9iZNtdDGlaKhKF3poOytuTtLXdgYrLfRwT3Nd+ZyURu1
EGVcQy5P6K0q4tM25EluQOwwt1rcnpYYduh/WD7IlJchJL28rSSQejRrCoG5/yIi
0PHBzDFVRGuTBmxgdCp6lovDCTw9IZgwqjPQe2JT1Le6J9PeHaeWEozV+p/MniPC
mojwIi1sA036wgT2FA0iC5QA1eyhEol9n3pI+eZ4SNjicleZURMFRAwVHbIIGi+u
bQE0WkkCsNdh1Fd5C61ganbwJGbUCVzWv4S5fJMJIE/U1L7RHCEI3ndpmkDzgsvD
BmLfJWY1s5z1632ocLF9FS/YAHWS/T2wubVTnbN8wCuZpRe6vwAf6zlpZ2MuvE7u
eYDx7SpWOLp5jEa0Ljgw3/S+I3s/M/4GkZUnU/Yx97AKOhXDEtfBHD1HFMZrOt93
ZznRLOJ0G+5JuIA/Nwr3X4VMHov5l9DVsAWsv++7fT5j7Hgx2DgvRnCSQddABiH3
2B3nvGL90ssrcYhbqbndBYGwCByhNkf+yskTSrU5PYfVkZKCS3GjyR0JTXsmLNat
xSdZ7L7M5RyQl+7gvFakob+cSf2QkoYccIfoyXu8JlhQ8oS2sTZbI4R64yCUTEM4
ngAbZtDzDIrbPYN1iWohAWKcB7RsfmmAlMCkwlG359yGl5HFbAqIOoHJlosBsA0Q
v9CQmG9kZ7KZnSEPT55DW1IgGvyBJvD0WzdfFpqOoDt9BKCFO/RljEeXsaAB3eZ8
+irdDW9mNf1mhXKFRh8LuqP/pa4+Dmd8LGMMmMqyMrizfINGkTFJfBaRLDkJIqLY
5Tldv+Fnl+u72HofA6zyzPh8hK9+dNRhm3n92FMnNwuyunXLrCrrFU88SoQgpFDj
C31O6fZNhZMTUj37Sy+xlUSLUeir3+S5UGBZatex4tiPhpGz+gs7kMPlBbjZeWiJ
YcxVk/Ejt64oXxh2kuI9bhFZBYHUbV8enwqiVpNL3jJzqPseR7GbqIgNsNcB7Xgm
a2/sMujrazsv0j5D90DESFrfhzaWrxhDaAWGmqy4A0EJfJnix0cgWvWH+Ag0zDld
s3Pz6FPe8PZFb0aDdQUHQ2fJ5Lwl5tF3J7dGZBcQVhujo9n7ZoSNkdhlDxfveTc9
7clnkYAkSokCNvWEBStrAMKaFIZiVoGqEF3xnVh0UiXEBH3XAHVTV4lpMqpHoT5K
HDyoBwyDfUrPrZmlqqh/JcLlmJb4U1wvR1vU4lUwK7dQlXqHGULqkZcXUN3iC9k9
tqdgQRVSmY20vvhn4LKUG0qNYgA4yNCvFg6Ym+QRIH0KduS5geqSKN5uYXi+G4LW
dEDuZXk++Qo1DDP5TFyJ4A6NypTl25s9j2XnwB/Uy9wT6LUFXOEwXZjOYQlL/0A4
DjTnmsai452MUQjiijJYv+Ro1FUq4/HPBP7LudWj45fygAInZHJnQfQbE79KWhQO
fMvITo+IclExjahB7XIuP3g8byv7ecLa1Go8A/DDCkZatfVLFU8QQ3kNslck5GiR
sKMonKZXlvbNzjia2TqiEnqpxl/EdwaA9KY0ZThTavyvNFJIlqTLUNPkHEfjNLjy
Fq0uK6uwPSHouXTrBhj4f+JvByx7cLykijbh+aW3UIPDZwuYZT5xwoxXNns2hnEZ
Hq1T8GWlEtGGb4PBEeSOSOvxMiyAbhj7u1KWxcZyqdY0hcbVfSW+tA3rO5qUA/tw
lVvPFE5jxwmQ5Spppy7EiVU+C/A8pET9wo0qf8drhWMIiAcdoqoINx6GZZywJ1Qy
rM6I/btv3oEB5s3JCT+r4zGABCnkCmM3MmL+JF4FVsnRBvVw3sS+4nr2D+3Vg6ht
XE7Xgvft8i+cSMy2Zxe0vkwM6dE784VLeDj4Z1c5ncNSSZ1WfH7Q3+MTEISCpfkH
tXkj89VmoFi91ehoEoN5cBSMlh3ZP8uK1/uihoN3a5TC9f/jCGIrj1+5EUElU8qv
d3cpN3Q/DEqYFfY7k+z/galXJpmESm3EeB0jG+1PODE6z0Dy63eBH0mz9yVlHp9p
4+9HMaa/99Fer6uRy9c7rf9dVzUIIWtrnmIt1w10rjhE7g5u7aehYwb3Vl0bqGpo
DVnBO/UJbWsfgqM2VqJmC1jT4b9h+KKny28HJ/fqprB2xSgMYAxTvnQuvh7oDZc4
/IjyhzqXefnjYeGhs5KYlFHsfhUmy1QAM3mgQLDjnCrt5CmJ1uvd0Raug5peEk23
FI+iEwSSbPCAmhV4OfL5OSUt1MXueWlQuw7uKRKUPSdOxR2UVyrvDnSFDHuAAI2h
A++i7GRfbiytvmMkyQQK9eM4+wD+GKBwuScBGEnj2CszGwlNJ6IARG7gqWMsrff6
OCz0ld1DtdR6t3EwBaOc8Y/zpwzBF2x100hLIP6DumdcQomueQv0mO+eAGHdLzar
W4cwAz1EudVEJXa7KJsNhHFUuJnQ7K3TXRb3pMnTeyTYAXAW+TodMeQSJl0So4W7
usJ4JnipPBbz13D1aFQONudRQnlnCsBcPA/+wF0BXsR4j18mBof9Lv0PYjcxY3uO
4LQ9Q6C6AimYCyczNXrKIyOJdJ3YQGJR9FAgbjVUATSd9x/Js6Bqvl5krw9jeAxa
OpX5/wyLOZEkTBQqli0Pp4P85gjLgbZEx+IiN0W99+8jBYQMMhqu7TDhVNPqke8i
ao7Buu1Bfo0ju8wFq0aqWYMTR5apsi7tEhbHGVwPNF6y4gFu2Gq7fAnS/vi6jH1g
Z8s4setMR6zbR5g1BzJ0jf03ltlJsx8tT5yM1vEN2IslfXeHhTqvzCsZk448WN6d
DHRb/1wz2XzhnQICEIFtGInrbe/BHkh0uU6jiNJAC87QI0qpl5WR65rW+cewJBZL
IznqBHPV+Q1nnXGOPeZ6EjMAj3Tc/b2yZjosrqF1M9zW9JPh8I14XKK+stzWjiZe
rHr0L7oBYTlC4zoqdMZNeYQXY0JLkgnHwCZW/S+YMYXIbo3CVlaLCGTaE0tBzRjw
slOejbcXbud4xeZy/9pVIT1TADeXG7HcCOW7ibXsIcztzGzb+hjM2JPNuoMrMZRP
T0TQkEnXz5kW3QAuu6dgaKzTy4s1zR8szQMmc/n+jXi+mR/GPRBeZMqaqBV1gzfV
FQfmCjLL3+RtExey0vA0pNee3IBBmuS6uNtB6MJZGaow+0QobaiKEFP/3u+hSuER
xp0YPCSGEShO47MEuHJNdadTC5jY3l7e/Yz3qF3FFHwuVAgCdt2nktkvzevBatOa
TRmDHjx4LSzJZ0J0xFU97mPERikafHJHQ4dhdCxQj4gNqM9NEaQM0ikWJZOYu/Fv
phJuY+a6NcKRM3VQM2N3Qohco7LlXzKTfBihOmJBvi2dZNOb08011q7mLstuFkFM
APnkR8abjUJoJ8FxUd5P9LaGk9LQiGBf8XxubK/RvEsdRNp1a6/+fZko77N+7kq6
4Vg8InawM9vXLOqEVLwed7QH30bOcI36DWwaH+T0QN0SMttaoBfjKy4QOkFAr5MT
P9vetJooC9HQ9wRxdpelerCZ4kMQaDZQ6FMiOvxdiXOmREVL8eHUte2ohuGNB0yS
XToYsrnv8STzprsFZ2z12kMm4vGAZbPI+Z4/ctWXUS9hQfH+C8LvaY0GWoZSihur
DxGvM/yVetZwdnKM8KVInNIz1FK0e8M7OuxZ0WEMCfM6tSNubX4cITKIJi0cJGPe
Qv/smE7/pC6StiKbZE8R3vbGHtW7x+OpCG6tr+ixO8zDeJ+8466ZnNlO4HuOgGxV
bZZiDz9h1dLUx8zGUrvcKeBztV9xYnTZc1XKCCchyiGIacELmLn8zUzherILMWT+
hmRxilobXcTUrelQuJTtmoLZswTlzdRnXSox6NgkTERGdw840tO7eouf658Gt5Ey
DF3azFWsBw2sT9fu4oG5L+ILHovRZbJme6W0abstvshXEri7D/ca8GYiKnAoZPol
bAVjW05QpRxCVDvsHOh3jMDSXm1ft+++A7IyBsY+J4l1Bq+ap38hE0Bctmn43okM
kXk2XswhWdKJLdTfaAIoxullVgdBPddPciH3sfmHLl2d6Bb85VYNgKolKtTvYJnD
v0CcPryvHWf2iPXfkdW68cZq01eVIIq8tIN3CJOI3OP23x3RLaD9QeAW9yF2bK1y
odca5VJN2MqmX7XQeFggEy++S1uuNG0y1Ay5l0Ova635ndtlkGrFPNpvIWy9CZWp
ndw6OrhrdvQZCVgbMg5bA1PAc0WKZjem/TrMysJmYNnBFTy+kWB8EVvYy9Cb/+QH
JACQ/kTNfEoOerh78GHp6H4WeIEZZwzhOYv2nQ3QuUEJKOpLafC15G+BLew86Pt8
ulyhvtsBn9xZGMeJog3X0nMuzMPFQx/b6eWxBD8CpYd6x1pGyMN53EzLaau5P1yK
gmhXX2JQZAfUiwWcTa65CUfZaShUr7jY17jKDASRw8mamXt4AY9JgEo+iWnX7Uap
CZpQr3Zm3h1plYkGZX8ap++D3E5xuiqBwEuTFrpGIY0OtKRgeWz+AUbGH2viAwM3
OYCB1awewifzZU0Cf+d2AcPO1OQdPA/3nKO9CcX8mrWcJDLbEs0kVdd4D0jI42T2
EWn4iMPRfSkYvLdsFqPukCGchp3OimdP5teUDaeiiQLCJefUkx73qWB+kqNFD+Nx
IIvaUo5026HT5wckd66OhabaZXDUDRaarP0wdQRZTiAQihAgWSMx/frtVYRIXUw+
MsbYVwjFg6w49WNAWgKw//115ErQ0koq+Gp/UQ21+7N5Fw7YbKGJbtr1TToZ1mFn
NqfaQiscx08vhaOl6x2tgl+pNTt7EyLhRXYu0HmQq/9lvnITzia3Cxqfdy6djO0l
vdiXogE7JttxtxvLe8z9sC/3XpcYeYXndfwlocsHwuMfQyUr5bo+GStkt5JOAVkf
RJIC66tS3PkiDpt/WYSTr5vbbyNuPAjplJ1zLo0e04h/lBp/2uFuHOIMlTrK6Zwe
v8SGnvXXDVlAqTULteg6nMCvszexs5DoJiag1RN2Sjp/7U53PqDKj8Bk2phmEXBW
+17YCNG9yDv7amaOddWggV03kiRbMOsX0QjkxZ8FfcmjT8gJckv1SHCbS5Ab35s4
4KWKsbdTfajXb+R2vDfk/AEgPaePJUHm/mheuh1GMz10m3G6wv/sLmQKfWo5LyZr
xLlmxYP4nXhBAbfK/rR0hcWCAwWbHaNYwpQ4fRre2D1l4AjIhyjvggnpY/WO64+h
RkpCu572G1UPE7h+y5WLSrzu3IMKKRuZbQdFmDWST3oT6utzIEcpgB3MD+z+pSDr
INSu9znzT1efDzPIuXglrmcStcnuz1IGfvx7qfaK664eMgJu8pj6TSL2gdQ8E2ac
xJhJQ5dXEvYYuiJp0NuwnA==
`pragma protect end_protected
