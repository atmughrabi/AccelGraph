// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
h+Dv1EUPFcJKKA6V+DP6Z0a5III2ROBLtEBwGitV7gX+xOW4mQ2WaG0n4J0aY1j3
Vs5K46zytF9YYE2NIEbpouybcmafNAMU/I4YCDVQiCP0FYLVFCYSPwb6N35JNRjX
ikOM+BgO133c16jC53TS3ddRRC4bf3kHICf6I0TU8t8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 58032)
TItYe4ZhDGrE0nGWN8RKvTQK7MoLJFG36fZZBE23ttar+mvsCINj4a9cUIv+bSOq
r4r1aeDRqOUxtuwboGkRMA3+dMeomtwKRzxgpY7QAHLdXuu/J1byIjeaTasTAOw1
apsOhAnaWjlGH6dBphACTlJtf7oG1zpKwOdsVR3gsEHNknaWrfpwMNPieduktT+r
yUImgtK2a+Z14N3lOADIxQqObizJUkQ+/Le/yrWOFeq4/Buqc8WWY1GKcLjB0+Qz
TDlr5pTyhB7TnxVfIfzqqAXCR0il6mgZhWd+A2AcMH3ezlh0h/q63oAeuT6xWPzg
8XYVLvcpB5seynTvhmZCSDd7zTrmIr0as6FODEUmonHvSaGSZjupmUrPOk05b5wG
WkNxh8MVQo0T3A20WCkQrnznheWNdOCLxyiLbp6FDhHf+k0GMIy1uvhhoRyryTdo
Q4Tpn9Iy9fI8q24Jp1/VLLUk++J6zjrMkn83pM/XYHQcrso3S4crHDkwcvZzaHLH
dDKVlhEG9ksl78v3ZXlvhgDxTHPl25yRWrnC8q2NSfnM+fdagznng7Y/g3vys8Ad
cDyr0RbV8ljZTThj0bOQ8rOm42NpicEUcZFn90o1vSeT2RQbPOFSWPVVcqQAufmO
mOrTU34AwTRBy3c+ZgktaOn6TSJaU0ce1fhoZHRLY90IfdrRP6a0w/F4MEmPrk3W
nr8I2EPfNXN9FOQAk4MU+bBvukbdWW+IaEO0n1EVnCC3VOiXmtUgkU5BMCrn45PZ
O1+yKrryK3JmvWCLvcDkjwybHFlD1szWc7q+w+kSpGqkrFfvHQvrjFsoIR6G31/o
dtR3LyBErOAzXqfCm2LI6VH0OV6C4t36oEA2iIoLEc67C/G0GL9XpYiwct/z/7Z4
N+htoKA1grYBZbwKMA2nMs7INhE0KqvmeEUK3S69MYRwePSVWzHm83nM14gj2g1M
vj3EwP6rmhhAX+4Bqi/+utV+wP9wC5aLn/2Ko6HwFWSe0ZHkJ9KunZMSfmd0pIFa
vT/QoeN8P68y4Eu9WdnyOAaCZ+8/WWBpjgOxUUWyZ0NISMkBJSbxk2xXc//5EzeI
PFwqzJE7HY74YmfoLm68BLcTTWwwXjvgilXWexTQKxpvdwjiSy78BBbPGSflJ+Oo
gWjzeqlEuwSQSm3GmQzTtkx0tqkzaXpuxP71z8rmikpUDucLlWWmUkPTz9jDz78P
oMOOTOOOd4nPh0So0B2mN5Swt6evB97ye6ZKZ6aHpHBEl17pLEkt9vJNxI5LesCI
tg48G0tToCxv33FpJeqbKGUpQRpbhDxIxRrf2MwAesF+Ngg3zw/WYLUtcIcPjDZm
qugufQt2SXfs1vFh7y8B3LTVoTTFdKdVhP21mOQXDyB8l14otsxYBds++VTlS6T6
havxpOwVsH3d7ppSdD5us+hsdhVZuKJ8zWdpqXHvjpA1mdgWiORkJnWCghr6vt09
XLO8CwcM9oK1pbVrEe0XYGlVpMEqO3/hjqfVpyHdgrcUOH9qJzIsZw/RBcXa9tGt
1x5shOhYeMxG6IFqSU7nlNYnWO72oAvmHGLYo9+aMp2Vdi6Znreww1yWPm1/Gh49
jQ5VzTz+Ri54zbrsZs4jZy7PAE4OJmXAZkr5fotY/CNzQ0PlaDrdfhLgiZx1UYC4
6YwzrXfC82AmyM6nwJLjg8Sfh2KinugX/tKQl5dd8hvJq7Lj7KEWSE3MsfA5WgS7
gIuB+BJhnCYDQ0R0mArg80EW6z1OzsYcC1Hdiqie5tYrlP4XiSySHFvTXw77YTpH
BHycYaec3OAwof+7PWr0uCpjGum9NP5I7xb8VvEesV1N32QwQLRRPNHYbysB55IX
6dvMh5FF+XOJDXibJd3B1Dwzl+LUFnM93aVVqVzHOFEvynBwRGwIEL9tLyv8GbIe
qe0fTN0K6c+Jw0x6mZk/ZcmwxpA5VpL5fqcjIgU4v37twaSOeqQqoryisYBYJyeQ
5tSo1DCbugM82FlqYYl1KTqYKhGNFbevx5gV/xdOBWz2kom5wi7HIuI6ho17pYj8
gTWfFeiaEUuOQgUKOp/HGACX8rdHiC7QqRDSminHbANQAf6mU/X5C7zgNtzZ4jhI
/NaW0zUZ4DYMO3UKj6vVhByzUIYYhv1D803EcIewXml8odvXB5bJQBeF9Mc6x5hf
z5BCmc0xfVK94RIlOsr19+8k006E+lTiHBhx1hO1P9ThOo16c8VeO3RJY+HXMfDu
1yeoDFlpYLAW375p78rnTNqeo/f7LgwxjBZ0TYQqxRnt4oMAKcPSRzm4QZPcsKGy
ie+76jZJsqtrDgpLNheaUqUOWkHCYl/JrXzlMwpE45pGnNNNABDhnryax8AkPoLz
5UWliidLgdnZTMDf0irWcegjXBU/j1ryizSHCpVLlTjYz43IJTCzyTkSPC1SkWld
yQFkGSbjgGTHLCwyVPK3TPbUegkHIEAgrakDvujAWZh0ERoGydWS/03RmJA7vCFh
nEGVHlvHOx9j10XrV0WHUgCIwhG4EwBNrHCOxdoGx8Be9zJ3fq7H28s0nBc9qz0W
E/uS+dxG3NUrfQc9L4rLWZT4xaYaeIYv0467mZNR0yyDF6el5spQ2NdK76K/ymyw
NigTp8QIW6OyPxJLK9M4ZJH0yysAxbDQeArM+3t86zToIolR3idWOAn7by11Ol5/
96p+oC+yN5tPA1yWN60dXAZrK0K4IHeKFjxJziFCr36XxMrACisC7zNfDlK8y5K5
CVrNxpaK/qt+AvVKqDQhscA/czX6eSkgOq4K/Y+rK5h/ygCzw4EJTrJqxnyUwSNQ
KIqZ0OXsXMzSqjR1SImBtShn0/GNesAL1T5+mODV1fJovEde6KHoEPCp63vXfvL3
GFLzlqfqy3sSxbqRmRX9IrsM1S1dyXkbjPSDZN3DtU9g2Z+ijzPi9qs1sOHyqSCR
RKqYhKGAeddx7ZUbQkNgaIPhpRW3rJgg7av0UOU6lncj8R+S56egaTs3sfK57jXZ
XaSrmDwBae+GxIYLeFjIS2UZYYQiUOj/Fv97NeDMriQXoxFdSVK58E6X+cI0pc8p
QEAjPNH6jiiOHMnW/ggwiXVg9ji9VckYw91fhmm0uTfi71IsSEN/HSnn1rimQsM5
Xi5isLJd5i4c74wpuY4Gr3ZNsV1Ya5qnvkeErjgulby/AvwZ2qT4HEx+hvryYZl2
wkTC8CzpWtufx/EO+RwHli7aj7WGOSyfOMAgLzvYDcTP+HPqu5BVA8hOdVzAg5b+
CviPl27ID2olPNlkB+F7BdqsXttZu0PkFkZtnij2NLxlXwTkGOh4+fzudT1yJ8nh
mNvl5LtP43IE6b0TobdfFgnh/TPPYutk2uzq7yRPq3PlnsurcHdan5hQ+yrsX8Mu
cbXaJjQ58HG45F87Z5ENxhpNU+ywSCTD77q+awInVhg5SgTzfybDFdb2yWlLn7QA
5HH09uwStZZYCH6XIp6KbioB/fHrTB76mGt/b0M2B3lSmc+/N+DUy9sbTJmAtkbh
pN3hIhCLpWv0aiqjfhGvW246/UVKB1Yadx96qffbaBInqMg8S2/nuXDpQHcIo81B
lkb3zQq6KOHDqCYy75E/Qk9IBWPyTaX6hPn3CwB9YDGPUNtL9V42N2IktcLRPUtu
Sp396qNL0LxKeP/43i2qNjoUt7ggMOvk2P+7Xzs2aDlLB4hyjtqQI+s+TmkEvEeG
bXzN2s5JfhyBypAyysybQBsj40F3yg0pcodhgkUAaqR8FBoe4NaS/4wcX4bhFlya
2tencJXkhlJ6N+gEWyc+Dzi1AXnqKm8MLtBV1Xl4l1Wya00nOnjqsbC8Y0REzavG
ySmnepk/zm398TfmtMDk43WpwnIo1Wf3hPQnrQTFDVwOxV4GzQ2aLLJmR8MTYIZg
f/6orbMvN5xXYNQDjYlUqbqPwqfNFMf4k+T5DZKkHbB2wuTmwvqdgXLQCGOyx1Ry
VsM6WBotSdUsY/CJsCMpKJ2MkLXcRuHB3n4/v8ko51cas6b2P1BDi4todLc26PCu
s9Y4UWViMC4fCyGYHRakm5fA2KwyR0LsuCuPu2m2XMAgdj23WKZdyM7rHMpI4Zwf
zETOa8dm2Jv/U9kbRL4eplIkcZDSc0UEZF9Sv8/+3KdNNu6+mNO5PtCWTnXHjzIb
DTYqyw3UZkmPV9a5AjiwLWrYXsuzMdq35lkjSNeB5KYk6yQHJIuD2LURDOupFxvv
SBpR1lDEczeU5f3qXgwRpPcsmfXffhxqJrm6HXtzXMhMCtnFGgskb1ETHCHVujzB
niAxquVShs2D82mG2Xy3p9rxK0IiHsS7oYzhcSbBrFu+dPd1DB+f94BinAVXqcx7
49HQ/W6HpHGKt7vSWcPKBFhHjbqscW+h78HEuOISQEP0kSoe+sAnxT96TlSHwcct
6CFXHxdo0BItklDKpwTDbq4J2zzjlc2uz1BiRtCFgFfpVkWZHe2/D+DzkANFEX6I
W/NqzcHAxD8NSw1rJHFHYim63SiPSv5S4kHrugGzJA4mOnGDw8pmDohgwXvyDgwL
01oK4KznIcZarI07pOmi6tN30MhJL5MBefzUio24pH5m67Stu7jQvaakK0rScxOc
yb7hRtyvg6UIznTi6iuTpA3fLqcTRNzQjgLPO3eeJ0S7W/jWeT+3E5uy2AHCjSwq
te8vlL7kW8P0sLB4I0KlSAD+9doxgapsQb0BMFYEDaoVd9VltabJ8sg6pUacwveQ
Z2mKVgfoVfE8r9AEr7XdY5TSOf7WoRQi0y8zNvi96JXrYjXovX0v53n0AyQIxUox
dns58boIfcbZUzEuO1N53gaH/GEk1StlnHhJLFxpcg7GjQ515hhlgYThXSOPIJLw
oPvf38ur63gW+HmfhzKdMv0GkPVpUxDzO0FkjmZf9Pc0UF4UI+S1AQah8GOiGgua
XNOBjmoG1+VSDxcBh4AyzMmu/aLKmhLhABZLhDr2wjxvQsg8JPVPnTo/NoqdOwyL
LpBxvavN9bmKVwoinXYiHyXdPk4Zdfte+s7TX4VoFasz7AHzm0HhNEOejpZG4ljQ
MhoYcGuFd3A+KVqyijUTFnOo+u2sM8DWMF71Xie4Q96A05ehgR/eMRCwwigUXUlG
qha2fuOJZHhOCwOSn2iofYa4jURyuy0dXLYFauf7kkPpmhCLfPSuKeIYK8+yzJsd
Cxp5w1g2FG1xpc8yOaSF3O2MaWnM/HTO2+ex0AOOb6Ig9CvpJzvtCT5cg7/g9pEe
6z4uL+CcJ/d9mu7/nYSzPJaUt6kPKg+EHiwGCbafIev5KtDGR0BSEHeIDdKwUUCp
YEC4gNZ3bwRTh7QYUmQuX9g2VbiTwRFfiFuZe6Lka/JtxCAMa6My+bdrdLYtRc/Z
fwke9jRGBvFeM4UdnfP8dI8qs/f5QXNWZ9TGWP9ucr047ljd8Lv9YaVUFi/Yz1S6
LDRMEPeCeKgphjRiq87yWTWlp8WtCD3IWbmjJW8Fk4Qi9gd2czdkxAc+o94D6R2r
il03atrxZ++ltevXo+kvb+Sm3Z9cNBaniuCT4xFJT/Mj8mROiYyCoomwKO9j0VIB
VxoyLB1tudRvW1nZ0eSOc4cblS1BK4ktP1C3qYyJE3Dyz8pyCih43mZbWH9sdKuI
gCeYUWHepFijYrxXx4LSKSkqWHWkDXgGjbpBvHBHBIEH6U8tf+YzaR1AIDJgzlOt
tojPn4j3k6bKXR+q5bMPGh4OmUFluwKh2oU6ejw9B//OzQTD55pHSjb2nPNrphYr
P2+iDy8iZNrFJ0YBzy4WRm9dcgdAAZm8CGZF7PmveNRcb115GPD0WbqZmlOH/Ogg
ncdgUN7BXI83puK3pTAYQ4oxy2df3yvQqu8YoQhrzp3QzFsOugK15VM805rohkwe
RtnVvL62sAirb3k0Q1uA+x2ICdLtLnV0lZFhmr+pJcIiaMTmFbQ7Mswm8FrDduPr
UObJSl2i+wSoCRCJ6QOEuVIgfJxAURo2aNrvi6Izki7xPcS9uES5bW/GECJ7Txvt
3LQIUt2vzlwCW6MR1rA0Ft9eTzaS8IrzJVdd8ZaOvhHeM/0DW5MaQKoArtZpVqhE
2MC8bRjCUZ/w8rFZy2dP1KkRD4yKdrZg0K7Sv5C8uKCt+8D5ZKm8me2X+jcUWbFl
070GH5oDBuKkaZs2qU9oQ4dI6+KBWFVe8Vzo3TmkGOXR+Z1TbdwyinkT9WKFDoK/
F2f0uCNiAU9Fmhum26hK6dWhqKuYenG0TqoPXVCZzGfcPB3tWtxfLAtqZ+soLdim
5G6UKP9GycPUxdaqq6ZHIesPgXi4vc0K96z881xfpoYvY7ZmFkWrqUt2m4ydZQM2
Px/LLuUGm57bbuZnbt7mWnqS+aLLNQCOwQyz26y/7oxTGocCbaj2AMsoX3tP+L5Q
ygfZNbRnBqU5fuJQBIowpwwfaIonIwUVZF0Lvj6ZBEGtD/ig7PyD+X/Ldu4ZKOkE
p8VJYHJ+x4odCi2Lqm7JRJJQo7e7zAPkinBK3Fg5o7obzKy+HKBsyLK+4q4BdY2q
Oweg5vtUrg032NVAqD7OoZeNPhWoqv+86AIFiXK8n50+YCZ6ZV8x0BWOeNyK+SL/
YxS7wwC5IF0NNyju/wTwx0CFAZHQ23xozWzozaCxeuNOMqDeg+sCeHv1cQVpDRKv
UVXgB2cgDX7RsGx9rsyvTGbMTmODa85pjALaKLyMEv9KQEhivswo8yUpGbdrdd8X
T3+EP4FtyKNoAUKHvtyO2SlHsuaHP8wlV3wtMHvf+AjF+Zk4+NT8ufIfDX4mY4Vf
FuiXbIST1pVwMJDrm6xWaeCLM1stLkUVYN+BehfSHYJYqEkKHhY2AVj++mNEl+FT
tK0BMEUDqbI8EPrR8cDUxqTJccrkGiRlAQ+Z8AthTBqSCHmfStr+vR7Pndtd2lXq
lpBTQ2Eu99jQNEGFKZZ0CCjrNVmLBveFGnMa7JumHv3amFJWIMJuKVYv+Taj0F+r
3l9afRtaWJ9+rOiR/U+iRDo4YozXkUrT/M2CbNVFWAlNrHFmxO1N4Gx50toub1gX
WvXEQhiVgoMZCzBJ0lAz5D1jY7rL/faoKNG1+pcmSQumHsYfDIg4mIT3xnG/tUFS
dytDm5qX7C4tNaMSdddoooS1WCCFDKjFyiYSKey5r3esz7MrgkqOe+aJmOlO3jzs
h3PuIkwZ2rdBfoxGf+mdwK3VznuKZSnOGydPTkTMeTsebAOV9S3jONt6sHubFIlB
/L8S+NX5giIZY4bUmsFudQ+dzv1aRywVlGfM1SmCEKzXkF5HDpK+X2e9ihJUta9s
E64e3OPHYm1QraPR8YTxweyXiVeIS8ccHZU5PoMpZp43+ptges2kv04qfDyd9cPN
J3kSg4mlyXhJxjqMNEsnDiUsw3tbnQARfOwTCvhGXTyseTWwatisgGBj45Vf9fsE
hrOeg5Thv6QtnhJtp74zD4RWqZuVuh7ai+xu4cB0KfcGqoedQM2cH0RfESP00i5H
AgHlWYg/5MQrVaZZHiNW42Q01ytuQWxs12L3IHzKANe/AXIZZVRXxppDYWojn4cH
vD0wI1U+lu7QeLVtP/ao397p5LPe46PQKggQjZ6gfLNy2lGEY3o0nYSeYRP6N6qB
0SD6JLw+miAUtYUb7K/WE8fyWB+KMCMXgjS9b+ck9iSf/r54EQVJCDbUnjM7CULg
JCHZbaSii2grhM8ggcA0ESlPrXbd4wh2+A+3xGzW5xF8QsZTf2+QWCevnws4q47W
9n2lILRZpmRkTDIKL8cRkIwx2weqjZTq+KDYYGsNNG2I9/oyyQdCdQLbBOSlnWZv
9FnhKHqGaNQHVafSW/s4jJJeSffUqinnKpF6/LS6aJwDCZB3zYykhYDoDasj2s75
8Ed1fYejmgzl0eJPRoVnTs3e8sNe4BECoSRNIqEEs0WHK0iqzAdVypR9TGJj+3OY
TPIjeFaMNRWp2D+tVn7gAROvxFJaoAbEHuaxuMbkrLdNI4Nk95BdOztXgDzNrMJB
1Vk5X/gY6B0LK9zae/px0NvV/iBH2kJmJCzCdyfSmHbCypezvY4MoDEyczV/FL0a
vql6YI/zy+X6k+wbNjCqbc65czy6T9Hls6M+SHZQJa35cqip1eOJu/mwrW4UXMEr
9mKyL0/WQByvZkQcAU4oLnQMfZ6aO65/Z1Lu/bmt4ISwdZORSVOfFrgVfahbIT8b
gfdF9/tFUH2JoczLrk9RKFkoXC3q7Ujb59jwoc7ETY3QE6P1kDV+YitBs+bQiJhw
tBp89IMmz0hiYWbMUzjYkMkbLL5oVQ9L4VCjhPNNfkHtzlXYDUy+jY30R6c23aK2
BSmRnDR6xk9CdBtO4y8p0UVxMeyZ1fYGvegmm6qjBeeJVgvOyWRuRBmNpCXhMvBC
tranRkACykJ15Bul1n83PcMZ/ENEBte6PclHau+WLTGF9GsXt2iKW0j+2VMNB1kV
YQZAZPUwkR9Wf08uy/GpVeVQiFACX211Fiv3Alq/CLEksyOcSRORn6aNTT6EvBHa
CDx8h227EC5fLki0Q7cDgnEvVZW2c/zhpGbATS4zpfXsJM0ergtuOzuYYUiZWf3Q
EuphLCAwgQLhSXofb6kYa86teztVczrkiPzlHwoJ0aa5NdWbvL9fwD8YHNrmVUki
p8cRenm+rquOhtm8HhqSLWMiSklYF/mngS5mhsqH4kwjyi44Y7LbHjuUMi7CCkPg
anyfB5rSuwKV+G+jmTQDOlnZOWbtj0eVR9hJw9LImDd/p3p05ink8or+XdTTsWZ/
gY/bqp++8ds0IksL4jHEFDSDbhaRIUTIUyv/CbBSckru1qh8pukB2Y7BLbVbYzkm
r6i1PXR9LNvHpEvNfiXORAbefpaFTVitrCeYul/K7bLRf8bMWBUv3EddUd2IZCLE
QbjqbMexb8L6WjDLhnvMK3GRMFhngWvfXBiqvWxY2GSImgtQn4o0SPa9p96uQLbz
UfnPvU7riK4D8LOx3en9dwhHItu1VBpZ6uuNKJHPMXZ8dT5+0xT+MyyZST0UEOM5
uvICW1LUJb24pwITJn26y587i2IWhmLcfGo1fRL+KHxI4Kkoi/G3TyrQXlK2cN8O
NXYbvNqOBByyLTxPWaXvCV+BmbStwrGZ3lo7HzrVfLGVg3ToQ4x9MO4SR6+BSVBs
9jjRebCxaCZsjE1hD/8Tr47zEvRRKkfvZ9qhGawt+lk6wb1RL12lgwb/nRhqubMg
AevNI+YQ5zWKhrkR8CS3WjFXS3a/er7aDWY1qSvGDftUlcpUy7/wYUqaTITJDBfj
PS3H6G32lAWlkmtXnSHCOUTRYnMQB0M7ggvGgA2waKYRZxu8KPWJpTzaB9Ij8Zjp
XF7zl2NHAesQzWH90FLMGPUJ9PiMmL/2ke9d6XJRY9Hpfaw/KYMMSaa1gjllcBzm
HFL7Cv/JZips0rYyu1ZycDkBREkBQ7b8zoKcQi6bbyqBPCXf/wlANatg35Xjb87R
GlqLiWMtB5tbxDQH6kjWSGNhoRsBaQzC+MRH+MI2KtEk616d5C/gdVaekICb+5Vg
j5rrjr/pvfFofa4ZhsuskuadJAXiHJkSxmjEjy28o9++VTFpWqzF9ru3Sg8bRFAH
J6p4NZheA05hu8R5kdvr7bnvLH9+a9RZXUw55FqGhGCD2KisyejhYIcDRDswnxhM
Z4txHgS2jSZmE5uFk0d09/YiUZOdjSs/y6W+OEnPYe7/pzljPxp8MIMQcagxyWT4
sNcbAk1suiuUTbsMzJ1BAS0zJe8UeXn17xutrAk8Ft3tx2EZKX5g5MKeSHFF/LVJ
lxYQDOFCEhKu/A2pJbEOxU+Id2voEhRgAsQAcSmf1lHwriLbdo8XbiAMawxZVvU4
EdY6eS6J5ejkNwEJW+7uswGabjdh1/uvsHUCI7EoR82sr8WK6y7uzkS8bx7XOzn+
6vSyEA0U6ZPcHFkgEzRxmeIM4y9BUTKRg3AGn3qD6x/m+0o/iIa6e6sbYo1uvurC
BTh3rPB2q3f9qkhscbbshQLggII3bAj5gYWYFxsNRj1MewYVuE19SydIacqSRGKQ
SVqK26CEotanfPQKeSMlPCeZ0BvEltlWf3g//5MK7HZjwQPI5kAsyn3WCOfGwkIt
FtDWNIghYs8wb3LvIB27a74Lhb/tyZBvN51pMRkWXw4wrsmSX4KRlu+05FPiu4E/
mAqdqUEEY93WT2QYqBTAJPBa2rW6+vXWoW7c/YdILsTspsdXhQWK4/tAagbsR+lH
8AKexNKht8xKPJ6Gg4fGzGr7e4kQi+K2cqP/Cf5JG2YB5UbqtrjDLzX78EzljWLy
dhLWcZM0n7b/1E+OhnahZ9aizKPRwFWIvvoNcESsxnfJQ8t/1xX75tjduzqR2eMs
z4cOa2RX+pszt/aNAmJ0ziR+PEZqafSMoaHowJgAl8vVs2Rj3X75qhe7f4MQpBFv
1EdE9iLcs/msflPFy2KIrFJ7U0uDJsnq95chZGnPofoldL6tmO5rDLpbW6yUaQcK
CZvAlJbg5OBTlspeYuCvozTC2E2v3ehgdTXXZSSWH/MYTlmLXYrNeJn1IOkypXa0
WVDqQD5X5fUVvezpiUHziAQsTTjSqtj3bBgVacDqpV1/2mfgqxzpOql8yRrsvYWg
SP+4qKlpJSKHQZrQ7XWoETKCVLFLvh3nVqzWYyC8w+YgnIxS0fm85GhEBHpgf6fF
7uLXjpjskqebQEIl4z60x5/aYiOzmQVgMqni1DGR5HUsjfkCKqzEvmR7lOLuHLuB
oF15pjBECsEfT1U2hTZj/+P2aWUaBBMR1d9+jV0ee+atDoJ/woEe9MF4LEXepv1m
uAcE5hsxY17u5+9kxvYssq9EzER5IWhI0/QWJ2ZmoMx1xHg59GYfiWKxxGeC/T+m
bsn23JPx7x5PS8HspSPOoS4FHlPXzoW81eJCqlo+SsQBeEmvYpbrZg8b8ASutPjb
8fhss1rGdOJk123p2BL3I5tKIE8H8anPoB2XoGTUjO0eN5NamGBWGkHdphU3rICN
zc5a5wnC4HSI/sdQbgKi0fesea5g8X07LP/LbN4mkR7wotQKytHrhOPICWcOOOJx
4aCh4bdNgtKp1sgsnIYj+apNj8JZ6zHt773qgFnQo+uVN84JUh5Uzdz1YwWS04YL
/oracdBL4Uz5hdPrfLXbHG0vYnmouJNaSpyJJPEzCA5lx1SCH+gmxkat1uJdHR67
6/F8KCcUlav71yTuOw7w+QgeNjo8QIbZrgESwNosmwf6A5+gnB5shvL01lbOuII5
raufDXZcUmI9UDXxSvD/0Ask7uFYW7dYPoazt9PBvyVaDrYVAQZaZyTcIwtig3ke
I2PFQYQAuUa2V7FuNHLLKt2Nls7globmItH2XKevRW3EuFAfXxiV88G+8AlcjL7C
E3ChgDywOGXg27zZCxtiUKPlVE1HwHnVl6sR2LHtXK5wzqDMJEsXvFmlEJBHF+O1
SyWT1yXrvo/oOogWsp0o75k2v7bFBAAy3dVWr9rKFVOH0S7NKJPYsW0r+vAHSSkM
WcuwdC+tUxYRXYRgyHRnYPLY0+DWDML+DGYOnkTvn7n4A5ryzH6rR0i6DmPmBoMY
n8nMZhifSVOOMKpW3/IcTmP8QEG4Ea5uKd12f+rEvSFHWb0T4PSrrRl4P4gG18dy
RG8bx7oyl5exUMarYrEEtHdzU85/eHmI8ogLccJlzu88sYzGoGssSImqgO3DJ99M
moBYiof+XsrHT9NxWr1LGyLu/22KiKbB/qYb2scW3wMFgmSdut47N3dshq7bCuR0
HZp/Kridrk3k+86jARBZaHZU1DeXMc5tFO1WqJdQvLK4svGBZ11I9GFlzzepb1zN
PSYhEmxuQAVBm5V17c/dHTVDYu8BlZat1zG0qjc0QqiWDBV+szL3Gp2hL1lOxKHz
UCLa77s3PekkGhk851hukOTycCxdHQ5lt7/BZJmQ2UVuYQWxkHZDOAOFwJFT3pL3
YGC1BWcfN6n2vAwQcFW58qv6Xa9DIUCmsL9agIb4D6/Tw9Ifs/NYaiebHywR2sSH
6yboMKchU8c1ZXb2a3qV+8/LEIQgRBIqszQtW+cPGWqyac7ccZUI1hTiikgFbxh3
vBfhYeu73DEqujM3jMxsSppGKv3aOZcekFz/07vJm1B3nhR7XTHVELQbuHsC+7dx
k3Jc6gOdUMKvuxYURpBWYOm46rCoO4Hc5UK9aEj3PUL6vXsYTyOzCTGAJtGSJ4f8
HxBB7gyA+dO4GlU+Is8Wj/h/Zz3K/aLdgIgD4hkdx3l7EAIHv/CmCAuuqbpKwzDQ
qIIyUxPJIoUMnxp8cfjH/GP2VYhldlLbwNvz9rCZdem5broOjK5NHgsXU/K5KwDf
6SzXAcO0zhcj98cj6ZfMRU8RjIYImXTxKiK24TyoCx9CaFFAyBvmwL76u1Hqieo7
URVLKKCMvN+lHyxDxBvlEXjGNEZA9Cp5ioQDuzlvg/LSwBeUXTeWc+l1dLO/8bOq
IF2P4HOZoCa78twdCaJy8q+7Gwf65wFwa1Eh3UkWKbr4GLaD5lKYYSztBmljdG5Y
IXAQCamSQcM71KQ1DOYWP+Iy3zZq3sK0L4X6UBGGmdzJX5zG9ht/fzULTX/cynxF
giTFKstYEdfk77xZKXvjokq+eaFDnly6ta8JDYJns12Zt+SMhR6W+a2Rq6ZWgY/B
Mcf/CJJvm4TDzEPz7mRvrRLJYB9rZL+Aoofy3Bt2nyvPXx4uDLe1Otq0hOViKexO
wmkZ5mbugZ1t2rVscjOxWsU+SerVEJdSbp85gsw+n2Qm091mNMSDC0uZJW78jZfC
Ihv8jT/MK4uqgToepcw5bh9eVn+flVLi59kf7e0ts3TZjpZgnm42u8SvYfllxzIG
1SPDwjxvJgsnWWd+TkwAdFJGS3hx5MV5M7Sc3mfdKjyAwZWXW2M1OnMyF/cChMDH
hpxyM4mepqVimSRCn7m3IBhjMW1IJE8eD2tItle0RKPTSM9NRWHfFgqjvTuxiff8
Y5l47j1JUdKoGyn4X/dm+Y+bsosk6biTjtcoyHumLF/WDsLtYuxuWWU2NzjLL/Li
GTa5XpLvg4Xly6MyTFD3+16jGGAOTS5QFIo3w4tI/NEiitPuhy7m9PaKam/h8QQn
4lFKn/E3g/QvVEe8I/3044ypYt23oMkIdSEgZJjJSZOGHT33ev/J6nZAaxoKEC72
eTKXVBuH7elhnHPCcVY+LU/F+O47U3oJ7TsH+TkdH7zMhI/yzdW8IbnRlr+t9iN/
4dnovuiR/dln5yUmWUVKN2D3Myqfg8E9oQULIvPKfFJXrysc6lsSSNwLY2Y6R2dr
EOQKVa1dKi1cddgYkGdorjpYGKPhwDN4MNeDsyGjZL/EZbtbCjwrXSDcMq3LOEQr
qGk53FRFBRIgA4qWn+rwZzMQ95FKQU5tP6f6sFn+31fXc93881E4oE1NPERdrbU7
YcLl3TFVwuEWel1dp298aBWVUn65NCuYCrKnDEul5VQE/nsNDcnavHy/yq8gF4J9
ePIfd9QmOF4+n4R9lNnXwu82i5oUdKv0MS5bJbhKriaK7sQUl/tLYazPPvYmQv1L
W8Wk/1fC4ft1DkbWBkZbneL+5xNUrMy6p+oJguQKXDJ9AQXqXQA/m7ul/rXFQVy4
ymOrQEr0j3V++mKQ4jb/OzxYn7azHZ9yeSOZf+de2KkaWu2yYU763anRb2FDNPhV
HmD6Eaoh0s1u7AaBPIni4otGtaALfnx5ylZSpTa5KcrBPjH6rKbmwP4XiHOD95D0
KpGAJv2WJCgXwZW9aQ41ZyGoAUXu81/Rm+TXyhWySisnkr09BOkc+5vT5OCw3dNY
T1ucR/fzzQ0M8XJW37I7bFsHuy0KDZCYbjcKz9/ZiHvFTwx8nNYCIrgT7p0I875a
XXHxdVwey3ZYYsBGBxrHWkpamQEe2r6g1M7Sem59nH5/qaSAX97Oy3+m1JoCR21a
cY+HN1Dym8i3XSwQMAwVyr4IMooSio3klh/owkSodLDbxqdfosVNutE6AGfUwXxB
W6Hxv0RSZPg2ttHHUYtE+9jzBcS5/qPnkXIeObgc6J3u479C5xhcqiFUi8md60Vu
0hYQfTupovoJra4CSENcf4NyGlcyYxdNIub6K+ljfG8ktXp/0rzPl08n92ca5/5t
KLSvuFSLmKeRuSRY9sjT7ZaQYXUkFdvjzxLlo1UdjRTLds89n/V8W2YfmmkLeCnH
OQm0h51is9DU0a7RHnwmjBx/AIkteX1UUSBSmlotClGyXJ1WqrkRHH3xkh7iSia9
woU82KD3poDi4FpXA7RknJV+3P8vVZSRwAN5hpckO8QjW4fas4lIXHbXpQDIt0wi
ETmb68o8WGyyf4OVfSkUPyYJDWyxaiT5lyDEUK8YDP0a0LRQIhthMKYv1iJem7O+
86dlnLr5nzZylQqBTzNORzexYWifprFekTWOSP1O6/rd95SB/KGzkYtks5IaRJjv
xqWI3HYsQDA+XrfetQHCJyEbE37jxaA9w48zN0X/XO/hjGBZ1J2a+NwoOnNs/8Ec
kMug3MYxzMWeBptjoTO8Myo7CAG6Sa6n9MoynogVUD0tCkh/ANvq9uNNI3bFqUMU
WO8jAI5HIbm5xS81GEfppCaIx+PstGU1nQ06L4uiRr9u8rwIZl0mL0eQ6LU2F8XD
NstbFz+Dfi2lo2y/7cngBGw/q7jdv+Ow9pq09BRr3+MIh6w9UuJOq7yH3PBCk0Lm
Kj0Z8dWUYee+Eanw7otOtPvF92+b/yR390zzh11g40WSLCE6eIs8hsoU3QnnxUog
XRmgLIMSGUTv3/99j2WczldhRXBAqu8viMoMc/Gc7TdkSHmQIes4MlIc9TVdf/15
81J5CrB8soSmiIN4YqhNoAyvvvU+ZRftTl8rgjMSQurj1IXAO8viuFF1PrGGh12I
/zkZ/SqIgs7pGT1YzcOLqLTchq5hiRUl+uT4SNsr69K0p5ICcOkMxst3UnC7qhZl
dr5z46Ekur2wHsz01qVBEl16je0ywsRHxC2ZwDCKPLxee3aaa2gMPsRllRLgRnG9
65CQvQcksVHSmmSsXFkT/n5uC/QiJoXC2/kh8gk4XKYvtVNy88IsZ+XEHsAcGEv0
Ud85jDHMTQFjl0Ons5pXyjCpYYm9M6+fUhl4QfgcmDhcKDIzCdYyRDPB7W2dH9nA
lLlIltVrgDY1KSdlDs2P5+2aEq7KWhtVnbXihHrgCj2awjOSqS1WFmQ+uZ4vTiYF
YOccQcgr1AZzxBG+ZTd6GMkBd/tV9wcGIEaP6D5EcCe2k7cUofBT13D5uIPdLOLS
LuAggskuKOY+FiAfTjWeeVfrepK1DFuCcJI8IrQMl099TVOZUe2eJtYMd6JCdCyE
znkSGvEqYG9mgoUuV+lLnHOkwFwPCWOD2pkBR9dzYCy5r8D1laBFl0YFrAzrni2V
N3xoV0/NhqVOQ7OPIz+nytVrhIGUSuhHtcWgYOS0+g2cP0fcyx6qvp6Clhs6k8jc
mqBBUnIFUWK/I7B3+jIe6Y1Mt4Jk7dKf5IZCHhNQTEch7p6lffljqyCzBeECiTDC
iw6jw6PaytTfKQ51fNbCuqgDzD9NSQ2ZWYFwkzBf+eKdScPJ4IjXH1SejGG0IFxG
Y7WXFk9ygVwTSfXs3gkJKULt3E70vhJ7dwTLmfiRqiXzd5Y6IOZaDzLxHYqgsaH7
NSLMVDEtW6udf2nNcbmXocG2vbmiRIznpdcXB7hmXq2VTTIu/J/vReFPTdhoF3T1
+XK8J1miSk70y/XhrybxvurTIvIaFeyN4G5Ido9qS/XyBXwsrR+5F0YbBu4Fi3XC
xF3C3cviMq79OdXnr4yLeyVbkiDkWLI1NvbPNZj07y87y0EtfZ/mCsevyuCobCv7
6OnvZXH9UFRa0vYjvHkX0KBO0J1b/fecdrdeVKvHI0FqWph5IRAHY7mRJgAFzIBe
ydoCRTxqTwd9AE9MnQ1UdDv4YRK66TJ4EJXmExfmgFmRWQxeDTeLepRBk+PE08N/
kFIT8gfwhg+P8weQMuNlrtWfk446bJ+0cFyBFjiGc/Q+cIusCSVfTjn7yPDDi43H
k0uiyyyh4vRSdr2Lq02l4zXPACG7HI2IaaOltoYxoSvjSjRLVGPU4jU5llRsISrz
hZhf9D39eUjpBvrRevOiwXNjAzlMIHvRlKG8PJd7JtTU/wwizGfsA79/56e3nUgD
VeJayppk/JubJYKBjQuL47Stqr5eC2v0i1gGjEfuE+5TV30gvhpYMlZrZgMJ60eG
UbxcnCJYpveAjWegG14th0DbcYWGbNJjDPsmM93ZoQylwliwRhnYPfhOjKanUnn2
PrJXF7Orz/OBKweGmXu+agULv99Ne/FzHKCc6PZZcWZrFUmxcQjvUmagvMN7ZVo3
1WvfXLN7M1RA9ZjKFoGVCv2T5ayBU/k9c1ucBwOA7PrQXlmx/uPURkzHaJX7lSLt
rndxRyW0LeiFElciV/ov4i8UNb19cWA22Tot/ZNhXd9xblfDz+Rr9C36hkAeTKmA
6wKmCT7KeguyDgko4WqtlFrPikyTcRtoBnEb66ZPOMksXOHIwa2n5NkuP3C8F7OD
S8GtPpvHdMbdrE17o9VLD5qBe35XnzHDuFuVB9D+3X+H53wII+lXh91e+NS8goWm
OBFUolnsSQHYUnvX/GaDU/Ri6TdhIaUh2TEZPs0urMUy06K+EWiL/+jex4nnBRHv
s31GGaZxdI/F/rllrTqQ26M3lAwDjQzzNEfmml5X6NpD+F6ncYOGJzOip/XV2qf2
fG2gWHDy4FWmXye5J/XsFRyg8ZcWZyuWUzJgQM4vjz5efFArJ38+YwaPaaZ/273E
8pg6z//eFboxegpKIOsLnwi/aBVt7x+peWjcbydEXdo9dOWoGl7SxaG9Xh9c0PJ6
M7VuCT8pP5OkEH5HP+zyOuGAO1ETeSThDCLkB+ZX1Tp0uKT+j2j6OMTL4lo9sVPO
dGpQ3pUYvzJk+bU+5H3KwEf0yWNQGe7snKDiXlbQJGRBjoY15KtFQvgwDBXhsEPp
qH9A9eAcF76QEvti3iNwuWUy8h0gFrWs+n+9OcnauOm+xX6sRy2/989IMbm3zCqK
uKw9nHAn7kS2AYsnhm9pQvGt9Cp/QE1PSezkic1Wfw0D5oM362VIu6r66+75Q8k/
27FlnWCi8r8iZStaZnfGhGbvM/J6K7L8ByY50B716IQVFRsosVJOiA+m5RYyfoRM
uIBe3anIqlHXdQ4X0/fgbJSkF5Z6jwAiGn4uxRd7gkTZT02YygifCpAPIWki22zO
PG4ypbnAAh7VDyCWQJ3/g5wkr3x4hZgzQjBJ9TE4nJRQAKgLE7YEXdl118AvrKNN
BKtCAh5g+AS/Q3H3SHI5vclMzeCsMR7MjEb9Kt+UhhbhkAcQyPOvojP3DHvTfyyX
BJQ1lvOpXs7PGEph6K8rs47C06G5fAI7o3h8qvGqJIuYy6iHzjuoCs/sLyToMmMY
zwjxZ1ScynZ57QPKTIKUMO+T3HxYPjWMMAQjYDQYhvpFEgG60JcQoNtNLMKXINcX
9zMtADu84iff+lQ5PfrCrO0giKsEcB2YoXi7HDSvRD6+vrmX0eUisAlOApmKfbQN
jKIr+k/YOsj44njaQEAE0oypXUGMc/sLhG7vyoj7L2P69PwCY0g85P5fuZcKmOly
kYmyCJ8CFp3c5MCd3+oxSWnGqDcJRucaEuoazy4uMpJxXkQRIwwNaYCW97zlfbqt
e+h9eu8nbKRMEbJI4MfMiusrG6jw0a0d11EtcPNY6aS/GrnbYUY9lPIhaGATQX4m
NxMys38ix545+XHHrD+bFTEcvhOuy65tXdkLF8m4qNIHTALRaLNSyKmJ/w60yDBd
yoB89ZbK/zRdXvrriZhaeXp3xzHDRDbU8seY0nOkP7/8H763/B0k1WHQ4G2L2Vqb
3zTUeCTKjh1oaKXpZRYD3PHuLrDu8XcS6I7V7Z9kVb8zhtg7x1KaX9/q22vNK0yT
tnklOWV1LOAM1D9XJzT+O3fER2sdKv7S0dqOssISDvlH7uA/JuhrIRbiMWrk3TFx
3oZoe1OHPuXFME1WaIiJeIgPaIfbXxNGQUoaSbj/6D3m/HOBe8nSyMlZjkiL5PYm
f+bCMcSFoGO2Lp0fjsWRKrkLLGssuuLrQvL1doGKxMAHHvJzk9ai6bK+7Y7fenjX
Ro42iYa7L8jZaTK5AOR8AjOgZOvG5LzEnM9Luhc0qj8MtFekwmVbOgPataApyg1c
5IV5kZwgPyxwi9rmcVRv0p+WwJ9CqwUH7lC+VPS7n09GbWw5vHRK9ox778cK1g/b
e8UlWH7MLy3eDAWEdo3gY13uRxbcWYnpmrJxx7irmXKCjIRQpc0+Z/YSzyovtLQr
20EZCb6r84ZUf64pNb6TYkpc6cheYLNRIE5OnAsrlaJFE/BazyDTHE0QpS32JBYF
nV7TzWLEIX0C9DtH2TkIXbrBClNS3MOUXvFLCUbF/itqlv8DAObjRzA8H6VvZUsf
4/kV4B+GxoaVzMZl+UeI9/ijKOmQBovZQ1NN4yEQViIvErpe1SFQKVqJzyN+4gb/
R+X53bzTFG/Y7MUSabbtWR6UUZS/rWhYiOFLmnPAJ5S/2Htx+f4FnCDHD3mHLkLO
jc/MhXZ2wdpq/zU9hMPm6slc3qRmjqfd+ro59T5ZPvMkNdiX7w4HchLzRVjjPVwB
l9z5GAfeVXO3DJAeXzBMBt4I2AkYbxzdeokdY5IjeuIFlPheVe13wYszOnppuXmI
1A6nx7hxcGn+8T5VSKDAaMN7PLk7H9W7IVDRu3covu0dr3cZlzof9kZblNd/nfls
MWBf2OccaaXX/X8pmUJ9vX6jkKb75ZazyepsJUnHCTvVFeogGNUeZyTlGhRU+UvQ
a/bcaln0Zb8KeWn4vzENzBBLjEVprQgApg/M02I3QmeWF57XkCoqE7/+VjTbWIkG
rNaDaWL4GR3sAQz6/6+8U9ym+7kCSJxaFczEPKT10kydlLWLwFjXeIORC8cF74jK
SYFrK1/c/iHf7k1GRF5P427iQIhuJn/LMhLmMSQGkVlyJHQ0g63bEFBmcK97n1nJ
KSqygdMlNF+oiEl+Eei4GzywAqEPkN8AMIDmaaTyphulcB6DdpRTaVBOODadP22Q
hn/Z+nBYLAuMqujDOrRxLyhQGLRbzqlafL9twnY0WtNGdOH31mCzUZKkI1Vm7/I+
A7eykDe7TXzMN8+I0XxC1eWSb2HwHiQW9H4P7em9+A90ZBo2CtOofvileCT7hi98
udrPc5LytviUk1dJLKUK3JsmKso7+/mPMCzITiA8Gk1YmFeqiBxC20AGXGjhkvFg
J+Ky4wwEeSt5HNrGjaGVBLBnaoARQWktjQ/rAb/F/IwsQ0eNVR3fp9621hlQVnUz
DTkfMyOO4IDHZz291m2fcRbLlZLQg9rLYffb2UL41TKDNFJfX5SgZzwN9fVmcrYZ
+bmaiQjt1q6VYII2qivTisa/igyrxY/lJu+vpqRbZ7n2daH5s0ySocmCrnY9gvn2
Nbrlfhwd/FroXSpry5rgu62Fyv4fkLAt9fKvnPDmqGNZIZ7mcpp2nglh83HszUYP
3YCbC2PC7QV5S7a8mOhQqyqzWZm0S4v0PknBDijAPvGPJFgw/vqXKB3sCypSRPZj
6o5UFxKzD+44mmSnTUl8wZrOUV6ST5+cPI94ubaIyHOgYclgFfs99YVmkw/vRL+g
av6jQ/BYCkzz/eUqiBFoTFnxtWbxpl0X44WbWl0xL+y+kHYH9cpFp9oIwmpkkood
DzZirwAscAJ9OD4DNjnacmNSx6IZuIoqfo+xSqcsTdBSBgTJh+sMHk0gqyAnq+CQ
ZpI+QOf+Ims5vAHsSs55PKkt9yKBjx9dx2KKmx2xAgxdpkePdRqVUMdsMqQA8Mjl
vKONC5x8j8n55+IGwf9mAKsgQZqNnA7NeFckx8KWmC/dkHq9TWq/scSlWfDFWNuY
PH3t3RQ0ivRJmJphbuNCcEJUpRUJbC2AtfTOqrDv0E+C/AdVxq50ShTGjLfux7VV
KlBDHnJBGmRw4ev2IwOeS0rWtT2xfivWQYukoiQWdCP/UCbuhkoLwUmDASbqgxhC
i2qX0IKAJBAgvsSW7HuEytGZXiAYLD0l1dBg0jyGJKKnaCueD3euo34+aI8avwUM
bo1buMaFVxAt41CHsTU91TDXbDIoUKdzbFJ81oczIGtbJZsFWsORwBIVCECy2z1b
m2lQHLkMp0AoTzQacpQJlzJu1OwNo2TGC1pPvEv/ZnNuzvBJ1L7/SeILqZOSxLnE
ErUBKh0lHARyRYYffuLBrfKhlGUPNbi4jomxLkX2ebQkr0uc5cVfcJAijNLLk1Ci
ORUsiRNwgqerikw7ptKQl0joNUMq7U5k9i2pxTJHIti3CvDsUzpo2pUgsBpMgow7
sXE3Zvj8EqAZHigQ6FOO778n2VmI+ocHN0BKqPVCDsfy1beoG4gmO2pirYIw4lS2
vTwuV/rbfbe0aB1rkYNW4I28gQab9CcPsEpN7uu2Elgk3pqBPM3FWDTgytYP0jC6
Wem3VC1PeKficARAhhaPwBoXeREIPb9hVQNm8YtPBI5FiQMKc1NtqZAOVU+ySTMh
sD/N2/IU9lklEDlBU3IrY3fk6O197RUKXAR/MZ5EitEgLP4sre3qYSPZsNVHZXTU
JJIQs7T9Yms98nAcsyiY5X6FaYyEEHyGbfv/rMemtM89kv7uG3Saq7D2TR2v5amb
uputg4fxVCLBq1vdMWHLZoZec1yyd/JKE/NC/XOMA7q1NWjpBdXRe1TZbEEnTQ3s
B2wJ6iN0R7mppFVuGmiqKwMvSr2B5ZnVxvzOtVFX6na3xJvwsQBHA6Mnr8yEiqIO
TbP7GHaLM8p+6dK5hvHGQj5bTmeDzDGiduHG7fi9PEKsqBdYMWe3lcTuifre+wen
Qdc5f8KSTziO3ImotTlKdtMs0k11v8uyV9pampgiAU1pZe060jjgelCHQLdc/fFW
TYFrG4L/ZeTPTaLkifJNZfz4K9FNfnvU16D/ujYjKNmqCyq0rVIJ52q3eMAqaMYs
Z8qEe+GijWW41SKr/R/6OTt6wOGj+S8VbyTE/o+SOI3DnydDUH+zpj/4tm4uJmGb
1fRdQjfMAfpjjioyAUo95BoIQRJdvjB7jbr5wNK6rRZSYcDf6gtFAhfZYqyC1JJ9
nhJDaAOgw+1gjnqf8GKelizU438vJrxqVZPcpV/K/pqWqJMlTa3wBSJbc5EDlMz+
ezRHuwLnJfy2J5sMbQika94wfIrUnxSjb14P0eXN0CKn6SVV/2Cd6qFmjGPiGahj
HhTuny3UmM5R6ZP6emmk/mlEAJl/Z32Fm+RvmxXrWytxBfHB+kJcGfIhFbXRj8oK
I8cWxVT0XGYz7UjdXa/Ej2KplUefYcgYPlQB69zBo8akl2o01eiGkJzx2OfbhMFM
vf3m6rt4V744LDy7SNrU5gkaVnIROUaS9dnMAph5ds/+LvRYA0sgy2fyARtsABCE
WMIu9iCbzmxJKVAUcrVWgjoDmT6D5EknB2Lbir+MMiNy1h0KcWNmYoKixZTJTgZl
VOxpWEbm0Rp3jJ/ayzW2tkxJYtRZAavXXn3pnbaZo/AdoAC4OTl3WyxmzxoovIla
5VLm/HisSaPfBkUxnFAGSUvVQLiL2drmL4tPzwZGFzwPA/4XLqDFtQF7eMewjwq+
2ew2F/S0o3Lc9JX0qz8Fn30qxXblF9YzJoMJv9z/0tnGyp69c3S/ddXYcMoe84bB
CucD4ye2WIjyDCNr+0H07JJUmu+NSiwkP7OlVa4uX41zKgIlyxZrrz8uND7oAdUl
g53iXNFQZs1aH9dlE2SXXlKDPQYSJDHFb+ilB1D82BRiAp6h+VP0Gu96vs724HdK
0UwLAz762yYXlCe1VhWewq5mhEoZKChWJhQpW72MGHex4G43cYdYix1egfJ0DXm6
lejYu9lFNqPsz1yVT5vcz0qBv9MPrJHHYZpBpA9G7ynQ0HxwSc7Bf0HBQ+CoOpVq
EGBIcaDfpPf7APifUNfAnRznl1yMYUh3YAve8BIdTg9SYYrhjNDMILKUWU6/C2Dw
j6oGVrmGfC2b1dDh8w28xKbjhvwCj2Y9rbPaMCI7xDUQ3lIdOWi8nBKV+Z6AkPjK
meo+qAaSW1uHXZEbeXcIb8VPplhrhuRCodLISEbtLhYr5KHpCZ27NqZhN13u/Sj/
wTR0sybTGLVq4DQUSPsw5lmyLbpzfbpTEebjURlZjt1uqj+EhkF97rBuV5rvXvpR
o0nBhfM+JFaBp1ZMk2CnalWZxBJ/aJvKXg65KnuWmvtBDGTSRY5KT54/mbrM/6Pz
edccmrVABeX0cZHgEaXgM5HNiBQYFinHr4QVMs4VSYYJzamY1fBAuhzMMH/yEP7N
2gY/4oSy9Y3LbYJdx301hR43Rq9BfCMDoNX8CVau6dCU5l1W4B1/pyNrpFNNvJr8
ybnh/NZQKIKKg5jRRAmFiWj+disYQpCx4lb9E6GvKl527YVH0BzP9RQ5J9CMtBhW
h0K92PX9+EJdc/d8WOm4P2jq17X06uMkynPYtUjJVE3LRlL5+GHbsGC2yyjjZpGL
WC2wKE1FRj5XtiTfhAjaxnztvjZ6+K3yc2BTbS/XEw3/h2Mz6bLmA457f6YTA4DH
vVqdkezZJ7TEJyL3Q+lbiWIyJ6YBWn6K1CUXlpfn17sZ/PFaHiNrVBOD7oaCIlBY
dJOdZt+ioszcq8CQURyc63AZ9RGNGspCQi3srqucVqAVj+6VIlCAZEmbuCUIF/vr
SwVsHaKO+uCslWEVedq6p3aUwdZvR4jUtJ4UoGyDp5Q5uTX+mNRA3pQ2qxyeiy3z
mwcj8zSwk3ONa1/2ayizwHslTZ1tL+1XzVcPWvuqbmAp7SvBLirVmwCNv60xWAz9
7ghFwhEBC1XRm5G83fgnJUWP16wlDK/5smnIOj8+noSjWQRQHqCETL4NV9mvjQLZ
/p9v9uM9CqcwNRs437AjaYOOUJUoH0tinrIyYTWvaIPQdQMuGXAzJWrKKsDh2It9
xp2QaL9Djz/fra3q2+jGOGSc3GoVjJT71KhqzZJ7B2rhyWsgMT83SzIn396gn+Ih
2RahoW23Z16I5VTHOc8GtT0q4IAKpBkSc+XcFDKzveyKz792Xwv4cOV/ZkzDlA7E
sMT+FANvRiSmHwsKvFWOUGLXVJlZCXW4msZ7Analwb4DH7thQvCVwn0EXodm01BI
ZNvfj2ho/XIeM/QdvTy7jdHKbQTCNDkfJhe/89WQLzm4Dz6W4F8a7csQbb9quwGb
4AQfkSEEWLHNoGaofxdZrMnSuzqugKKycLflbxXlKEc/ZFmBtEAop+PpgFfbM2Xm
53ELknzZd7InLvC3SPBArMfhpnlNSgAPBUReqa3FdQu4QyYeo6DcV7TBEkBc2LkU
ULiInaCOT3ihBfIpNSGMfdCxZk/vixCSENj4N5LnRvDk1Uxy2KzotqMjuWb0OozB
F4WzqzAlRcKwRQNtEfdAefZWOVo7OjQwWI9VKt50Ou8Y1BzLYXbFmUT8nSJd9CUT
PgRcpm/tLtRElCVhy2oEU4c2X+NU7BX99yKirlNVFzgreY6jSdepImfRQYirh3AY
zdQqVfEkmdoJ97ji1FrGjyf0VzPD0kYGlYABnjCa50xO9Xj2MAGguJXhOrdtTf9Y
u4MAKHtLuwiMErrqhYR1CngIOfQKLZfsuDKvhUjw1hD9PXHo4hflrPURe6ewEFk6
7ZI3jGLSFWHVckKlntAXDzO+8kuF8qxbJjzlmv87CdDiQpC9I929fJY30K5rZ04l
RFuyjaLzM76cEF6KEd7SF7/FXDdZfnYIETI8taaUx+xUyUcA+OIm8DvGSNx53oH/
OjsFFxBocJ2Xc/d3qAcc2pCLO82RqkajqOaadLvD0pRSsnzEzVedoVL2orBrAEpe
VSMkV/IA3P0zOUzalxEcq+/bANWtJ0CrsDLoPHzGQy+UrouBSzCj5yQmEvml9tKT
kry8DdUcEmQ/aFS5pWJ+UQRdiCsdN/OgsMQENTli/hmwn/xegYZkPN66V+FOQeL3
LoyqYIdzK0I6OwBYOsa0nDsdfsO1PH6WH19PcUtq8SiQhmN7G7gwQvnaPhbKl2AQ
7+izsPvaQLoqk6aFOYcg38A/Noyf/fk+nNCqtjs537rDOWFD0RN9zzscy12DZMhj
uhJLHSQCq2mtXhoStXIk/rS2libQJHeebIdVrCvrNC836Hyxh8t8mx19ScXRbcf2
mFK9sSYvsWku9gZaxTExTZpFWjt5JLmZxS9BOHIyp+YrzijNh2Xl/WZphx64AQH4
QKBX5w5PWt/CBlzyNMBFoTDckKw16G3/o+KG2+m1NdibZsO7FRjPxdlzOBed3rQY
p5I6WQx6kesM2tLFu/9KZuefHokhi4jJtt29y8WetCeivmEqSNzrpH9KxDF/8mGE
EsC9VOZG6hbvuGCNbPE0k/h+eVjJQCfnH5q+TZs0Mwpbry1M2ezPEr3cq0bLMucG
+6X2OrSQWBVI2OpbQfjy7WAiXBhlqsp5w8WoWSfkUscYVykqNH5KBVLsNCZlv2eE
+lAQ1hVSE8+G++UD+L4FiNmoPecdqAoDLa6jqJymcD2dXcFTtDpAa9wqDE5KvQgr
uRQasTFyhI/aRMD16BQJ4rygjQr602gN+UXH+yqqUKtlbnRliKj5FEb9z1Wo+S4E
pqvyzAavilVxgM55/gTNd2eF09SfvaRBeFzqgBbcnjYTMXB7zxuCRZhduzQ3yD+4
JLiOr0O9HB48RChrYUx3YhlRZW5q2/3VuihbRIb0Mej9GNZdROeUcTj8A1RwP1uT
kTHbSyOmu45gWt7ndMBzanvcg58Zw/+Mg1NU4OfNlrLjgkuROGu02/02EGbNj37P
9ISwcI7KZLgS2qoThXQOQJhuUrZ+ienYSchriSio2ndgTarmZEodbRkJNKgTtKee
1qoLAK6THvb7OWy2PoRNbDnIPHwY2RV4AQiL6NwmqOG5nQ5lMLbwDT2jZkb1ol0K
uqKMuTuKzh3dng/dlmhLb2I/U0GGnFwLNTpvJjXA3F2CX6nFGCWSs9V9bSGJH9sj
IanoEDi9FfFzMKcXoOzVsT+hNaM1ZTyQA0nXyK4nr6Y22iBcNT946bBcycQaY+gz
gRXNq2IMf7PEN3gIdfrLcg9lWp/FeGscUH7BTDgMtEly6jtA62GbI57oIkA+skIk
IClN/sNZovH1bu12P71TFYzj757uSfvyfRXSlvqrBKKNNDcUHZPG5EO/kIp6nnqR
PusR+R1AZdwSdzsx4mWv0V9a99zYc88EwbH70zcTG0EP8ZHmG0MA9mQW0qcCiamD
NROhf1bsyqJAkSV6yLXcmzoledV7uGNeyxj1dUz8eHj3ES1XSc7lI6ofVreNdc3B
/Xf5XJO2k29QvUXk9+DtO+6kDQoFOwobTTq8Hp5ldtGvvpVrGAf4IIYfD7Ba1n+U
I3F5o0i/RPMPKQnjcfHhNegLDbAoDSro2AOjGpGBeVa5kvi6yxsZ7FjbA95N/SBA
i5bhBtavDWykmILER1Uxvfek6UTUKpG30DiG4U36CvWdq5gmbSABxo75IzJ/MiJK
/D2DZTboMY/U7U2MFVBb/wHk123PPaiIp06W54YCLJ3vZB17t2aVPFwwwplpjbmO
MFyH4Ii5bfr5Pp6j2hCqs9P8tgRu7nydnWBZCMsuLVwm8EXrmHmFxcvRLSgQhJED
H3UTvGAcQEUf89wsfx9TCHlkb63GhAuoK/MX/K8syrrJHqTiPnbzF+/2vmMm/sK5
QtGIGzp3W4K31OTB2jbV5Y2UsjGy+3+f45bGqc9x3QbZGhHYiRlz7R0k/19SV/wV
6G1YHjnGe2CTbFBXyBLneyx6NS7KiUJI77Vg9CzEpVfwGgXd9LjqB8iEyOqcCjiu
CdohxCgYxuehZ2qFNTEjANOw/YMvqGTQ+zS3zpMhQDu+zBGMGzgUy6BajbW0CHFH
04MJiaTZ9Goo8IGwlqZtz86hIV0pZstvRBXWUwQ3Qyw8tGW2MVN6ms7jfjwZBxLw
VOURMliMgGURlYSl17Lv2+LzW4Ihlshupkq/EYtBqubPxWzBcFSAlEcwQDhzwqVK
28xlHCPtGComZ1uJ9nGSInWAe1pRHm3GXyBxsrviHoeAQLaudUgwR9wRTyMcRLL+
ez+M+G9sTe8njr3Q9QutDEc2KwB2JVfztFOtJ+fFmmy1u09NzApdRUETEKlP3rEh
JWGTARr7JZlAxWNXYGNExn/QXOmQCOhTTaN0qAia8ySatrHYdf1lXJoK0ZCEgP7M
aXeGax9kbRRXT4+VDuHvGE5WPZzn6XdZmNasD3EdpPptQV9VaroGlmRNJcJfbZyl
D/cxEJNbT/HLqwn6O3hll9a5WpvMphPdVhZoPQHKA6q3L+SMpR/v3UyfjwMrebTu
t9N8OM3MY7uieBtm7wyIxeuHE7Yor1ZKsoqHyEgvvFhL1sOymtT1fsbvK+ApL92j
Kb1+ArPad1bq5HE5oK3vO+VafqaiZc5BSfF/moauk66lXfSGeHF5b8ry5SOboWPV
7crw9GbIvTbB/5kmZwUwNluEYZQkPk7hiYUJ10gXPaPxraGDbL81kccS0A2k7M7J
YMe6+WtQJ4uhRR6vrWV1EZWrd5NfdN+kQvmRhgt3uqiI2yrJTcdxqg5b4RWl3B2y
imJLJtno2aWqOdR8DR0t//y74TTUFl+OiJ7OVvVALQ56yMvwHzyrMH+qhpFoKygH
CnHxPCn4Bm4scaHyI9MJb3YL5qIjhvxo1+E+k7dUVsfvCZuu0PDSAQ6mHeWNlWNu
F0voJ1LLwPqlCZP2k0vMwRX5/FAukzidlbPNuE1a9ZVODGwgf7/r41gG7MYFPEVE
0qgS02gBBNrzTNbHPfbesB/NoIA/J2gZMi/ypqGB0aZVM5yOkB97tk/djrHhTPgi
beiNwsFRtEXZPdqfxkz+VKjgp8LZBdtT8/2+Bakrjl7z1mNGFAWxSXkLhgkltDGT
dan5Da/D5ekrk1WG5qdDNZKd1Rvq6Lej+7X0ZBbx157lIDHH16u16m8gtk4/vzm/
OanX2DnmX/zQkJj8Ydf/yXrCpsVJgciqjvX/jsN/aOO6A7XRCsC+1OQRTI8XprF9
vc5arJOPh2npL5DUM0h8ptjSAHsE+d7eB66IRyDeBplfV1tE8b5GGgmXTk8x5PFo
LW438Z8lkqF/yPTDvFF6api6VDNCFVblGbdvHfDS2UeLiHrMKTPywMSVRteMvDf7
F2mu65S7Y/UkovhvbBP4v7daAkYyhnBUixSmfJfk8ONwebdAFtWBt0w+OYn71ksQ
BgMv9lv13aZ/ouYh18FouRjTQODMzrQ9sPJAx2bl8npRtDZeszL1TEAjjCYGS6aj
Hm2QQmD3NrtUn9VzMjzp4DV2XXbhnJJvWUBYWx/VJWv2sqgyXp5442HNp7/5AtyL
0GkBPUqZaXtZwLWyYLGhLkqNB16QBsm9iRq/SzUvcbKfkLcO6M4DjF1NpkdcNDXF
3XvmyMcZmZxh/zl2YfUXhLnyLfhXMllJHIB/T5yu+N9bZZdp7eMuEzoEIgs+dKCx
TglTntBJCWFMg+bIWyhsnLRQzumxOLMBUxbA3s+ECP0iIC9wTJ9rMcEYS+TRSYR9
kSuE+DvsE+HWNlLkqvU+aUn8MQ1w+Mqws5TvxBIYAay/oxDZLt5kGJyQgT51m/+0
6m9CouQHVf3RatFnCP3WtJgiDyDiEDvnKFx4STXQ7MZGqt7SEfMMFbuF3pl2Q7Ss
qJfvUJV9XqOgg4ufpQutqKUqPvpryIMu2Q+G/THwwRAJnh56QxbMwp/KmqNWf99P
RswBPEx+MeqYj/lwNddsLQdoGScuwciEDfEDlGaRzlQrHJd/PQSgzxS6tJ7WGMN+
MhCXv3VeBG08iyTq79cMKPQSl9Gy+Bf9RLVM7Q4u5TeHIRbpDrLbZKgQxcs5X8lM
qNOHWDVpQdGbtey2NFinh0o68TgM9P1pi3bwX/lAo2uLJ+yhmKrFNpZR25Um5DR8
pNUPUHG3sXV0K3iKCkPF+rVT6Y9z93MGekD5mL3zUybc1K3ihcCcYCDF2r56X2Aa
kOE/LgSYLptxYaF3SUfdVXym+szaqQaUkA/uXbTQYfNOPIjpnOYE6V98mYdFO9f8
uJQSFKYPYW4nLCEXAYZPoe8ajsmvzqdOQKORC4vu4x68ldrcZdfPGaHqfdT0Tw7Q
YxvDfijzhe7dHlnwAFe5RBovBi+fwI6KX7eWRFxpiHcBdzgYySp/Ml7FRRCosAbN
iK9T0ad9adWx4krlvU6UK1uytz8Nq77chbPcndz29YI2NYMsKYxFUD9rjNhLNV5X
zmCA3Ps+6lqDbu7rwJ2t+qGbYOVVdvRjf9pFkh+HWp+SjrU2/j7PgkkjFTUp168o
GyDAX5/wGeVgkH8wfPx3I8hawcjsO1ZOGApvLjnuR7ppKpBXXwrUxROZqPBDDU3f
CcrdSU+r/u0wskUyT43uUPhtX++gimSdBuMq9R8AoNBREyaLPNGPMYfPZpSVuxAu
UowPbSEC13E7Iy9J1bG6nYf+Cmkr1UQiGAZ7J1lZjKoqQS84bbVuP1KKyyyA/yPd
ogPCzoXSHA7nh0M/8QcLobbnxqRo6GPbrYCdpithIWzdUcpfN8qonx2cZtSH6aE2
p6JUBNOycsK8W153TPuRIk91pFDKVBbwjfv7e7UD+v0QhQdhQGoObrzzgmtvaRQZ
YiHkmre34p6F/yEdkbQnhPeV9e53c5QTnqXHRgN5eWiCLSsSLouuq1BrwZ5/m4Z9
mbshb8gI1TYlc0P3r6nWGbHX1x71cW7YhYE6wA/oMxkxXABYQQoXZ6M+gW4NQl/A
F7uqRQ/DG81rqxDA4TKTc2NeK2pGP0Focp8VFrMPrtMaXxbikhuO4FEOKOWwS573
go42fHmFKIgt1lAyGbWgucjgYnsXuaLVRdyqvzy3uCOUWh0jJ5lxsh9k8MSCoud2
IKp1H0I3IUB3Z8e2oyp4siKQ4Ml3CpdMHAHRVcBWT+mIoLH+c8xC0XskIshE7gLG
QZHqJfkFN35X+MgPjpvZkzFbqzlRV7s1pRNjmuXVS+Fbmwbb2nrsXKP2EZP+EsB1
nlebL23YOMMrnsehlv6IWwMdvcHDlx75MICMCkIieGaGHo1zAo/zjuBfWScYYJUi
+WkLymqgqv4sEsK3wFMzDxqEVAnge5k/PG6sjfv1sVjyWz2pNybLQiS+rCw+CU6S
OspdqUVMAOmODxsTZV1CfeJKn+NUha3OiEbK4DDmn+jhvoSbH2MtrgyAd4Aipjty
Rz2QMNgz2AgJBl2T+eK/JHXP09gcoVsL0wpNKHT7zHWhCNOupMcsnUoFXnY+nMp4
5wWunOjG3slXIjjNgwRqW2rhO4cEyhmEPRgG7elKXr/eSHh/j6KeUVpWG5rwFBW7
wXFrWIf2Wb3YJaQNhwy7pS+m9x/T4W42yXKFIx0W4wCd5stwuyVdWSKrf22AJIoN
UQkj/rb0vPphk4rfcf0x1YdiUMDVfIEOx5568+WJJfF3NJIakYbMgpycu0J2zoq4
8fUsh9S5DUG9bQYZAD6wgVCXFqIeXRGRUN0o2FAqahJdD7anBAZ3WbUAnfkKyeS/
kQiyJP4/3YBR4SGyLx5YOEcMyQoYgDA/6mhciXVLFJ8KQFYoJmQF6pfgPfvM19LN
sKwI/4ik+ncMyjeHZm/3tlHSCameSQT9Xh+SwFPpUiwZZG1TssMFEIAZlRsXdlHN
E8LCUf2x4v/F8NiJZ+pI/IICAQXE8iocH72kIHnuPKewuRER+k1A73CcU7VIMmCa
eN8I6cn8qv40IC2/WCTt05E9V4VyrSt6AC61yemUyzDajT22GiT0vXBvM7Ht++/u
XIXLjNgkeJzRL1SMATBDG1BJeIxXw3YvXAxCCkLKGZYPNcTJfyL5JAN0RnDrYVQz
7tFrKw87yBPSpT7NwDSh4o7bQ9SjuNQOy2j8+kX6zV1yxuX1fxgkihYTKZPMVKHz
k8aq0yWyaINAycTNVr5J9Zus6ONot0x87zyd5W8wb/23xzsT1YZV8CQ4hnkb84h8
D+hOFSyhM8RwrgqovsZSTrlLWZdK6OQPsLR8E02jSCKVI7fCbvGv32R18gklP18s
sS2wqi9wyDohFtwOxtzoznOFbK4rbsw+y/VTdpaI+dUizdDN27h4YrWWUtluXoYf
udpke3l1jBDNe/H/m+u8oFOtyLGYK/bNlhCjw/DU5zIVwaXWmv/K6bO9bnAb+ZHt
9CdTZxypvv4Ihu0udm/Ox/TvrBechrmLitkAPC146IDRzpUz0p95oyQJt4euNa8I
jI7UA2zpsGI2NW0qeXPzK7O+57+LsbVyUcGn87qOFWyGjL6CNOXoMV4KZUOz1/ea
2in9dQPR4Iip74URngr2u83HAMBFSZGxjI5Ya9NhIe7pht41SVy/bf/EUFqWoEQZ
TCrVQjr0mKSN+q8OVCtEVv35bCf3r05j1ff1mbrcmZG3gXuVZZGtKGGYMPuS9B8W
apuF6m64BnDx7FpBOQ3ot3IfI4C5VZS+nV6kmi7/XhAhroOil/lWJD7ccv4MG8Iz
P5QK+5tc6vH7REGU91/cocvWJH4+qKslUCI+jst5TopVx8nntvLbWowPavBU1pj5
05tIVUZwrzUVupKWa592zUghGNzoMP06VMlHU59gXv0mXMXnJIoH/ekfeWMFVl8W
SY73ql/S/nYYtyu+QmhCqBbhw/gygJP89JYTFch4zyh3xOmlwjodaXORPchSyuZa
8ps9wygzAli0oh9sJwcYBwWrZ9YyKAufZKs/kcUaB4UqP3SXATyEqI9xy/5xe/cQ
WIpxXo+XncBVuuVwszPZR7IFKV0VVVimFfO1vrqnb34ysL8/4rq6NnhZ/7JjW8Y6
Y13kxsYnf30zD/Nvv2FMvNvDSlpA7Da7hCd7HFJxQW42Se6K6bHs7ix+w7M/jmnl
Xo+tu0gC4xvcN+RX4SpZvCn4DZP21XR6glX5dNyOjdwfNVNzdrg3v0Xp+Tu6rq91
PMB3bV5Y8JXFiYK5gZophtjSx/xTp9T2X1kjzUdrCJHgB2FsaCYcEkXI8a7nVVLL
vqYwva2epra3Afcc74MO4JG1A9KcnETmEwegA8i21ghgA+12FcbeGQ1RN/Q7tLVo
9r+dOOl1HWYXbh1EVyMkz+rQ2vyI/pC4uLzDXWzrlwbSUoerxG847XeGfhZYobSR
1jMZcZcG8dnpziRP8evt11YuNxyy0l5B1ChWIz/+2EUHrD1QXHWAsRgsFVNy+ein
eyxLfO2WwqMsXvW6Qq2auxZURb/GLUQAYeQi/0RfYV5g2TmBwN3KSYq4e56JurfW
fo621Lnaa4em05oIpWVqrGvjIJVne28jUNGakR6cuVdOPOYKtigXDoaN2ZBi51qU
rQxe6X+sdM9YVcDlLZBJN+2i75639825zZ5gdwirEHMxeL2LyVciUbsn26YJx5XN
yLkaSLlT6ElrN0Yan/sSbJYCMEO7dpm1XzWwQMKEQ1CJLU1I9F45bT5lxPsB2PQR
ArMGBJiIx/+YHa/DIe2Z+xilmbv8eoqGEzgsfKdNQgI3b8qPlfETI4NSq40DWsqY
aV2lJ228ClptAOH1w3DqSc0Dhh8A5oRWaoq8DQdHiQ2rha5svR+AoPfgRNZbCvZe
pqzO3VGS4/MP3EdMCXRZQwu7HcqvsH00TVBKWTKmpIl48+h61RYaaq94u/yYjKKV
Rp2u7e6pXlz7qdqKnQ4uhC8XzloyGdaLPhpD6fRhYT6a+rfe8jjbM5h2Ixobsgxo
sn4sAGvhlfUx12r/mIRS2KQ3+GsYfzb5NeY7o2dgljqWaWoiaJmYzU/CMioTE2OI
Y6VmV888/7QNOKRLzhMGdG1mAh48u0AtawVfWBZFhpKI9J3jcpZCzv3/wXWqCsGM
41/3B7RG1BugLIJtN8ZjaQ9MdvhUEvC/BLjyMP0uEMja3ezNNfcVqmbixKXddwMT
GbYQ+jC47dgD7JMQ5Vd66cZdW4tdyO8Eajarp/QrcrklR+e4cd9jBkvkqcTFYLhA
ljYa9zSoExvjsY6caMKMSZ3HbS0tvf4TnXhMXPXBpdlIF+ggkQUI2mcDRLzgZ0jF
yz0ZGTP+Ww5Dd0WAhTNoWfSUMDmhmhUui6z49rbsJZtQ2z8FIcEZcJTfqaLeU5tT
n6Wq0Om5SvB568sfCrUGxx5hfbpTpDP6XTxgFxejN96hggceupTDwPwGI0UoR4h5
/BVcyN8FFL3qCw+D9UfbCC/VlPatYWx/UYWI74pIvaHoWOy1NeZgd7ok4et0NNSY
i/ig0u9xmsbFu96qzk/I7cUkXyL6jjelp1vLFD/xrX5YTxoW2ypInwgxkGRbafsu
P8gQvuvlCc9H3+dJ+9SRXGGfi6NTqK8mm+BaLM+QXtmh81fOfp8DCaUA7IYSPscZ
Dg1t7NLaV+LEFzZi93GJmQvqkvisOTA/X2lbyZbUQjfp6x6tmBW0vOMYNEY7IEmM
hqDK/gSb8PPtYfcLjIJA2Ssloa3B9+wUrkRSvDVNguh1vVL/7QyC+02zePJzLCq1
mtxzJDt9L+MJqgZPdKJ+Q5PNbXx+4BQnuNtO4ZgDrditQQjXGSrqv6iqE/ZTS4Gf
cZJd2nVeFL9j4D9oyaf+Au8DRspZ6yGd/xzjhNjN5mWOmKof0Aysoyins/IXN6P8
6iCaQxJAl5Sa8JmbaZJj4SCttSXihXiWcff+ANg+6E0F4/Yr2ooxBaif49PZBJLw
MKuVNG/NG/gU3q2VuuiRJ9oeuty2PySL8ZTJiAooKIQFeSZvDjBuSVTNUx09d+PB
GuDACtvCdhRhEr0RH13FzHoN/g6bx2RNlTRm8qxjIC5hRYVudFDn6s+UTfgrJ2DR
1jGi/Hdub+QVMYeh9scRHqeqygzQE30J5A4LckGutGT5CqPqQn7Tuv5ZVUuiuu+m
3v/imuLKJNgRJQEADiSaUuKmUEMvd8v+XNHqWnFhvxnK2C85ipAu+Mqrwq9s66LP
twnoJ8DGKoo6InNytyK7HiMnBYg8ayUzm+CJoDaZteEhg/S8a6zH8AqCyDoj/CeK
/RTMbKhkPQT6oR4s3AAgmmsqf/nos/gTQ/8yPvfLgZOWJ6JKtTQryL9vV+D9QOHI
Lf+4M4bmYtu4HkvQ6kuhO4lqmbVVY+Elr6S4HTwms8oNVXrEP7AppaVt3mbRDfy0
71dYrGCY4B4abLitS94zSmcN+fbfFBxmAvcgbYcWdV8NWiPb/wOi2d0LtrII8A6Q
SPh/PYKtjWPPs4pS8g+Bc/ucvcJC/7K9bMLdtsuMNkYlgQSL4Ml2TCJoPpUZg+4b
Z9BQNt8sK3NaX/30S41VITW8NKTKQTEeAFh+C8Wx1zrfPOx4i3Ace/Wv5G8B7Np2
cXgzST4166PXLE0APyuVXHQaW9o9p5skYbCSF4IB0n056uoXSB6TqcJojFL+UV2S
Uy9KCWkG3zIx3MZjMoXaX7OW07Tl03G8wosQbBqauBCfviJMQ6XXtoZnH1m9dM1r
NYReax9g0WeSlAvZDqXcTzpCo7FZnOHv6B7n0RGbC9Mwv1RPTv550QkJUtXfkVQ9
9jgCucSZAFJGDc2GfsU48c5WJP3RHsF16RZQYnMy4bhENoNf9lhKhOrYuKJtXmrH
PvmY6lx8VgyJlckRgAhB6yfzN9KXCECoyFW9T40imdFGwzccq2B2R+zsnnW9ZZKI
0y1mMbS6bZ9zJ8kjssT2xUI9b6qgzYyFuL6oLzGHvuVqVCjXhbhbHq6eykU4sg/3
jbwODJ0Wi+THWQNFr0ynM6h+Pl1BUQR/UDPx5w6TtP0jK+2xhAQbjIx9ZD1iBWeR
nga0Twc24xCF+zxN3njenmDDgul8Tk/Ua0VNs+kNPJSLO71+tB16pHoEbk2DIG6c
5PWSIrf1oDYvxRIOSU20RVgaxKRPNR1or9plxrFCyyObjL3pcZwzPbvJq5cJnY0Y
TIGGaJZ7iTGXW1mgFdOGRdnAOQpGWaRCy6dIVDUmrqO69RYrNa1x+k1ZU+e6gNta
776+JUM2vBxNiCM+sCN6sON5iik23Wz9MXoFTtkLV82YSoL5YaJNdQxF6HsqczVi
pqrKK7l99+tgGCuPA3kRLg5IKOBmHZfOfHkhUbfHlskFK0NKtd6QX5+gq8DWIe+G
ODpcyEnKZpD8EqzIk6dZZJTMsGhIiZ5GdSafrkGTRGWqp+aNM2S0zEplE7WI49L5
OtNki8Vwupq/7kNJNsxtzNWha/o+hPwr87Rp/qK1/HE/NC0LWP0p7jHeJDFEynLW
SpYditd5OfbdzDI3H1HeG0sGIwvic6EaiUDXkpZz3xcawkLKo+bQtOAyANy/VISh
KJ+6rIwzW6xLXVVSFeG6Wu2+ny/7HbqziYXZSU71N4te4iNsqs/E/8VUIOMDNC/t
bTJQc0ALAVoqNXkmkiePMpIs9BzUAhWFg0ZcxrzLaCs37c1CL9wco3t89mL0l5DK
k+VaGSRW1tNKZgb/0sC7Xaf7OvYG1agHISgXHftTrl9EgzGQIkZGD2L0Ac1K2Nca
4bu8nS4KU9Sfr1V2Ziw/0X7RZtL9fDLlr6uz0YUE7jQ3PIvabTpLWsgoGf+1ey2c
f0IS2s1nfVmjdAcsjCbACz9BRy4DeixCwr7otLkbIyeYAkXT0IsL62Ln3nSq5gr6
3wnl8XgqLfDihCqt+nubuhULEWg0OghK8rpdlu7lcPekti8e4L5q1X9bbYo2qSx0
lepM38hG6VY+6rz3DkU2E3JfK5Hb39XTeqkMzhbhtZjPhirb0ddF394CygzH8G9S
nvSmc5rHiUfL27L6usjcUi0Jo9VI6mpInoVKUgpQ6zdkmgX9x6P2E4vwxjrCixLa
QYfNZ+CGHXgYkddaeoDoDySBjj36ZpXt1fyK86bzGOVYyOqwTzTUV6c8nLyz9Ljp
mc8101TwQHH23CSTn3245MYYgStyM5NRBpNZ1abraK/+WAeLXoylXo0C93DMb6SX
V7uwsMubOQ5Co7usmmja7lA0KBm0NFnxtfsqhGUNBy5cUSHpJ7dKYFk5pE0E9+iT
mxcAgjUzkJchuFr+XxDmc68MKDkKpx28aRaW5QtlTg3S4H8CgKUAL7Edc21M2kdE
z0qxxCC5arVp9GxFvCMopXNrzY5hTI4N/S3l7JC7caw5ktVsOus/wBNi2tIHNkmW
Vm9svc+40y305LPReHbMIQOZt2ncm4HaktAwgAQoSI9HAk+9NGfheAKCOXCkfw/H
jAKNJXeoIKEL3bqG2x88NpSH6mlc3iB+KlyhKzkyuiLRZC5PSin4z6IDBxHU/jN8
eGtiIsh3RF+xN8qD+cQ2QnV2LmG7WHbwv/sq3wGr8NdMlRi+tu/4c6cWyg9pL2Eb
M5x0Wm01p3ee+vq5gM8Zq2jOHXVVxUIrgB8DX/y9cvJGlnqSBifeu49Cr+h0i0ti
Pag/yOHW1rq3P5D11OJ+v36dHwrmQczQGWsI9Vv5SUaNKRjUtGROtBvprN+Pu3jU
k07/ZU9WZunlHfZbOoYeoGfHCsAPmF6pB64u0q9X3DRTzhTgF2KJw11u8Z/ly+Jv
Pqa2aUaVas1EJ5y1nIZ9Jd6m7nHopdXh9IdcATJ2qeWmimkT8oeO4ABHOPRZ7GEc
jWfFlwhJjmpOzCKqN7p376R/uxaKoI2H1ktg6O2ikY4FywnwjqGiBJmIF8ASixRu
r5GDjMpKWso/v90BMIcT0Tgj/41IiqZJ6Wh6Q01pOW+i8zlIIlmF/pKh0M+6z9mT
LJOquzQy/JZ5NzXEVDSF6PgVPZ9+KJRz0NeefPw6bqBmhe0ZTWjg3hfu9tQazw5e
KK/tHEKEnTmG1FC/XLuxRogH6H9LJprPsXKyHk5NIvbYEiMmkB1v8UqMhKn3/JIl
HJ4EwRMfw5GHO67Eg0bZD1I8EzjEfXeqmZfKUkZRg230IF5CIJNm25C0VLv9Xbkr
55cE2tnDCWZ/or0UPENC2IY7P97WoifPNU2ZF6gI3bVEf/NIO9Yqi2+qMkrwmyc2
Y4KtkLNiHAdLLyNgB9JvdXfCGMq0uZZXnZ15mpHcfF6dlmo/v0yWZVmY1NlogoYp
9igZswA+gYQpOTbg/AjpW7K/ro27h9QQV5Zq8gPELSMjthwfOFkGSU62iEK/zkVz
ZZXoFcmnMMW7vJNVuGEp6+eqQFNQiwI70e48UdSET9VRpAEoAO63FeRcIqGlYPIf
Sy207R2tcIgL4dB4P5BbZRBC/75ZepuU/sPUlUR1TuY4aZHpEYU1zZOozHTVPG2B
oO0mrm8CdFiFI8dNNpbYdNHj61kkGlHatDpP06Fks9ruGqxMn8lxOY472v2Pup4x
qNfqF1yY+cmnQvGOMb0BJDoY9qduUzc5C3nzIyGBx9dIWs+0NmUEoGdYY2V/gaMC
Kb1KFJNODT4BWKCqPYaeXUirAuw+qogYHs/ZTQq6LlkLKCi6GKnOrbWgVs8ZjnPG
ZoIBqqUkDUB9bLGaNvZQBhNEWJvw9HfDLipS432vRRDdCjmxk16XnEWrayG0ZekM
a2e+hm20shUc3ymqBjDtNUUgQ00qG/JVRqcgmjFejZ9tbiduMNUG+nC6s6BEnlxu
xp2ivB66jAsN+f29yeUhDX5TCnqvsNcN9vqGv+oGm+00Sq23yZBNTBjOLIHmd5F2
Xp4EEH+I3Cr/MmGMIOHduDhy7/LtTg37ANjJHYkdLc/cPSUA3L35h2+3EXv6pUxq
HG2DzQkX46OdDg8jV2cYjVDEvFgoXf7ai5c9FvfoLAQ6ttDLMB4T5196GZAUgXjQ
5SaYoTqCMuEBL0woKtCpi40u79hRAyDnQ7updUJcgeSu4T1wTEjoPOrDdoolLbIf
KJaza769MFzvYP+DM1lNmFjiR9x+YOV4vqF9DJ054d5rloSjtln5PQ88Wv/9Geio
zvCdO6Ii9JFmCnnq8BwXVb4pIsXkjcdmkQ9Iq87lQkQnSZP2gLwynsHFtw+eFd6x
5++dYR4fiQ2iJ+UlfAKV6KvZf/htBvc1pECD0de9GtQy3lLoKGPLwB2Hf/5XtyN2
BOIdrK4/2l9Atd9T6Kl7w37ZHo4Z4zmPnzMV7X7y4peshQXk0bmTCZHdnEro6N5l
31Aon59AxIZPbvnGi90NkJLtueNZVr01GtxLWda0h11mBq3hN53lCiq+usSkj5co
deV5LGFU7jbJlAt6aIC++Fw0JMHdyETXizN2mfywXls7/ogWnDjtLBxRWDeK9Rhk
456WxXjO1xU9BjadvUiSxVpBpZdxLmP3vrwY++JQoad9/HKPoLMNxBB21aOjKevr
Sx0zpEWhH84XpkvTzYauAUoJe0LNNb5NSMVMpGs+IEr6aIhIe1w6+NTmlYDvClOU
/9GWigW04+T24e/rF2yB1IZifQFvOTRnNMjJXBaDRnQcCFSmcx6jP7pKyJyb/DWJ
P/LKMbV51oFjRLkYkGSuE4sxzr8oSyaOSmA5FEiMFszsecOBbY8eChczebS/MhOB
ujNzZFjESv7eMeZR4eyftLokC9zr8OpFBbwLMygwqpVJpq0d6d9+9RB3WOITVYeZ
FvE933oDZvGLMZk8pVcDp0dWQmfnF39fTQW0hltWVVJig/j4ZmcHRFbBdSNYBvR+
U4JbEs314eLNtmW+ILZWUPzRpxQ5h46GT+rZiBIhTcQHJ+oAte1UNvmVrqUl5iUp
Fd7A9YWnT3ACi+hhCIvkUTn2cwo2rDlDETkcc2EY3Iplb0ViieVkizJaSjNhRjS+
5CWZ+rqZFZJE3fiVv16sq7/rFnDN9QRVqvdoJVIp31M6/C6tMoPhlBztaGzl5LQV
u+HyXhfF7ZQGQpNXIC9EIFnztcp3I9H9ijKHgwhzeEwXDQP9Yri03GLv+8IUUrJ1
6npxxXINBoz/vdCtES2RlZK374/kQVJlfQRl8oPmxlvM2zEJsqbTeIGHhMqr0hkI
EWEcRPUvYWDhnOr/TzhCvd5tVeB2wFOAE9/GQr384P2gxLihwb3/Gl4CJTOprDg2
4aV6nWEboib98f/NGjCM0+w1bF4CjxgPHP8zhfUQkcvmCBmTgPsfewFm3irXjrAF
niTr2gARwb2UBGNGvlhoN0PHlZyy0tt0UKOLT/eIGFamd7U8h8rzegKnh8t+0CGo
86vftXjPP/kv6/+PcHcn6NmphiRnqHYk5hw+dJ7d3qQkDk8Oc8si6LqpIdiZHu/D
oPv/87Y/b9jsMi4loG1Y0wXDhSXl+yA7Rk88xBnM2yeE0KXnM0Lekaq+Q9z3912J
FwV5k/53zz22V2UaoOArZIfipb0yc6NKSv8dKQJSNChwYz2PnVtcQhpjr+qm2Dvj
NYmRRS+S9anqCY3SD6sFe3VN2hnNAuartGukUnwgMih5mWyWRG2+RP7lkmTsNmmh
k+0+dFceHzjL9UDBkiyst0EUCzn8auFbOjCMAuBZI5Vw/7yCFo6Ojid+3evO+su9
lClgcZBfX89H8JejxgPT4WMNws9l9X5DLhla9n13MnJq4eb4ZSAKvCQ7M3wRfToI
kZENF8lVkxgeg54siaki6DRW7PSlzAFAvQofpiuTzXGu5W8mRWR087MBpTzmgZl9
1FlwwVST2U4kVGC6uGMScK77Nh7/D7uTxjW9h5sYUv6RrFt3qZy6DJiKxUQssJF4
sxnD3raNQzzS0JPBfQXrzdC+t+aGexiBsm6NDE0Is6EPGXKW08ATS0WGqoMr+zGp
DSEub7Pb+hu/1MAQ0d5yTfnqs+jTYeJJ6OHiUr33U0aU/em0DYICUtRfwkdxkMKJ
/wF/QD6sNoLDfTA6PfzLf62uHn1s+Q4z1hEA/w2bj3oWlDX5Zsd+tr6AN1LKsH2j
jHEWaAU57ohwblTDVmCjenS4M+3OcuI/XOkz9Hh8jmq/8aQr1/8l6zAn/fDPFkUe
DavTbg5DfU21yaS79KE0Uz8pJk65yEiONKFVRJxvRhjk0L6DVWPrBzuLsdrKlcBw
IW+fR5g+hpRGtHMbmnuHJk5u+hCnbXlaTQp1N/d8EoCiHlo7KHkFH8UXdujfKAaT
vFr7GM3uwOIE8mMSlKKqP6PXta+Kpc36tMUBWzqiNNcLVyf0RQcBPeyxsXLaPueH
ffBPU7HYqswcTBMjPA8d8BknCxCyul30u08luJqIHzXsSgxlpSOwhoCnTK9D9pNM
TS8vSpLpbf7bMkEIVvDoZefzdnH23rhB+vZ/1vla6IChgtxlxQLqiZljsorh6Mex
qR2ez8jaeVWaLPDkO40hitgG0kUG50N3cIi1hBq/N1Kp+Gk7oXcB/UNGNljNxJh1
RqFpc1ljC8A6wyCOV0fu19oNOG4IoM/9pjKnIua5phsrhrMjleoPAbAnntM8W4My
jDXX+LuHrXeE3SCQjvhMFlykAWSqlLRxOh7fLRgHswkCtctBQhDh0yanLwuRQvCM
I/awjL9wR6GEiI2mtrBLLM9CtrtJlTlrE+1wfo1XfLpQiD71na7N6qtGNbZVt1Pw
0nlBC5U2VLqlr3oAaf9c/JNVhJ9n+ivOkoOX7Ok1mUvwH6/T2192TR5hRBrW+fuo
zzLpw9bGpMS3EjXL7WGiKb0t+FCNrAZ3vEwGtxlFyQR9ryWsoLshRef2PHyM/1zI
Aq0ABmOhSHZ6+7IQanrOd1e0N3YQSQuW4/Gq6zrimR9ndfBUGVYK7T9heUFWJHWc
L/QR82AKkTRXHvt2kobjwiAQgKHgsSHdSniP54xkKIpo7dBpOidYA7yT61MRV6G/
umoF56IBWla4SgaPLLmzytuwKWbOSUvtfJGRgw2DEqbDm57PELx4EEqQsINGUxNH
e8UTySy4B0jTm8IVRGvtPkY2QJ4Igt3EBEoz2NFpdHFoTt/l+B/4y0JMUiaMeD9R
6UNQ3dE/Gb2V+MOS/dQIOXCx4KEhioPVVsoKMvw/3JNeAqK6dHyQ4FOWOWpFWhc7
608PBLJZ4G52uMYkqN3Mfl5WFBlvIA+ffga4M8XkANfoyAwW87hWKahku0qhaMi6
2hUTvNyjhXEMrL34asW56LUVWbOy0Ldvc5XtFII+TNHyRCNlgf7cOXaqlUeoBCTY
TpW5w4SF+gxIPHtoi7ijMNFWBpAJZ5yHYZUzABjJDHY5p7iMR6Lum0+vOelqQ0WQ
yTs16yj0oo8AW0kOmPiGWtjV0QK+eIImiClc6d4YRKPPQD84GUq1GsvTPbl1W2V+
GnNlu4Uq1xgRb6bmaQ/RbdKPI+AoSEdHe1UEjnvRv2SCsl5Sbjn7KSdxa8uvccNv
DBFlV7fsY2XgcwZLfR07p2xEzUtp0pYKqerfihGK9RLoQI0PLqA+HdVrkC600Tvm
3j95cfk5HgX/CizPovhX9PEx6ARTqufOXAQUS8Y3jTxKNjZKi0TCkrDNzRPami6F
gNTo71FBnGPHqg4hSnb8hAna7AZs/dX6TN2Su9jsKIVpFIzw8/LHAD8WwFSn3KLn
CzHC63jUAUDKN2u6tvBqe5uv//r7egIeC753Ji15A1yM8B6HMF1LsYFnzcdSgLV9
I14PSX47DLOHE6Z8jujv3Ltlp6MESMpyRR+1UgF/qyzePn10UAOT+y7Lo5HISicW
2ThreOS0CJk/1ZCCeti+CCSFaWmhJfR3r9OHa/8PW12Hnm9+6yOhdBYff2oTLg9+
rUcssbw6VABAHmp6JvJTSDJ6xLMIC9v/7HNMugBzwqGxIV3JM82GMj+bXTskXnjT
fjnI3Ulhd3RbnKh3XC3ItPawGxtFo4JqH9VX/B5XOjWrZE4Z83VJdrpI5oWS867/
hh0d2xSviUo8IZk+zRtZCrtOagBmT7+qGHfT5pbNDOCHPz+lHjOSa1s9Y7WokWON
xNuW5URcHv2DznhTlGqTa4tBIj4HlzfNMS6ZYDwICRnuKqK29kkVWV9rESaAaAln
DoducqYhwCTAG15TYa/YlhJWEr9Anug5qUOPOLj2pFA4xBtbWqaLz1qbEAKS0sdZ
eNRM07pfzCJ6/jzQsmGCNOi//n0402EgtQ3CieTvTjIFi1aT2FQhEw2t5dnpQLI0
Y1gTOhXYLYodfJXrJpFY9KnJZAB6w+5vr4VxkQ+t2NHYkHuuOMnh3yKiTyfPe0mM
M3vBP9ksguw9Y92UTbEc55D6XX0qk/DcXjEvfMvA4Z5+DppPTNoQNkjAYE9UuwQ8
B7SrdFTf6zVPJ09e32EAVjfc47JADW2r98FY5sOdgHMisfXWmHwLyD4byEP79O0z
PHDia5Sj0CnHRKqlkbLXumSfg+daCssovoiZJMpqt5UAcP/udFeXqF2lG0NbxPZ6
E/vQXkc6z4vASC39Lrk0du7TSS1YnhK24jobgRBiTsMt2FphyYYSWZBMG0lUXz99
etlq21klg9oDZdy5U8+82tdoHjwrazPeZg+n2Z7jxx7JHZGxDBKCXcVy2yY9BFTM
sux2WsVJcJzjrximsScocBkIY5R8Yb/uSAw+S+lndcUhK7qTP8cmKcpcwvjhLAks
ZdU4rrgGM2mVFvks4ObpXQPqL5wzI53x54SQWQzSoSPqZVVlcvSdXjzp25VmuJ0c
len98rY5TC17c31l4rS7qmeA1oQ2Ud/1NK7zV1BsTX1Tiq3s//x37YRTWxFoJNpy
jUjBIfoDe7kNO9TDRvkP6EHwNdM6IHWfRgw4tQakcSXvpz9ygsoC0UM0Otvjqk6J
j0D0AwWYNIapajtwYv0wCcP0qDOZ1OpggpELVAFNN/eo35Too7H3ArbAbBIef3Y/
VSZYx4/mlfXL2ckhds0ioio5gI/i1qf6O3o+nbg4YhbMO6OjwktE1aUQJwnDakXC
wdVmFa/6CQk57P9io0zkhxvl/AB3fcGT/tmmbl4wZzfblbh1diM51xpSdTFbTs25
zsjOdmOk8yMUD27yqOdw+cgdLtlv541q0PzgpWpOvKM30W+otbCZYB++jm1G2S+f
B4gwac5WktQBeflJcjxBTOuhXISfHPzjRDYJbNodwadjzZ8L91EnPXa1Ymj+71N0
UQvvUWINzFSkL/ppWNk66lQmXCW6nPtFogbboJEiIM+N5DHc7bQgnkVim/I5FiSP
yiI337EgQs9kliaKk+lfq3Lf97zOC6R3s+3GMkmoiFjtlUJleAwwUhWF7hFd1xcB
QDGgTLwhJZFdn9NMvhpFR3kqUjn/c9b5cyjoYeMVEEiUSTVrOrJ74jnd25iKsyKN
893RlDeZyZo7xE6IU9qHt+37Ly8ze3QkoJd+BkvK2MFU0FQUFKsQpbGaH3JDAgDC
x/Q22Y5t9Bz+FQVdkQYh2QwSb+6jvf+ZhyfzV4X/neHxQGzJgyqePR0ojR4PF4jd
ufjKEa1zp9zIRcRhTALGMKvFhvxiRamfwljIa6RX4+FqAs2CbjROMCN3F2l/GSFL
aE1Td0wiG/mNkdGOp71zaMu04xovggr2ptY9AVi50hUUK6Jn1XtPzzx7AVlKR+or
BOUHCaA1NjcSMOPoA/I/r+5Hj9I46BrajdJ44kbdmKhGTtyzAgFOPYpvPgWAhIfT
/f1h7nU4dF5IF1iXmblNRmJ+nILcWnTdzuJ2UkJKQNqhD0llz7rpQsfH0vVvtqDR
Cvj/Hb531wYdRlf8ReooCK/pmVDdU1fE8TaR2tgvqLAOiy1RWl0l4kdrYKcEI3Wo
LeRAEmqlwwTAz/CS2muGq7nGgxma+p2p9S5r8GF7wfFwUnn82hz3nB550DQAShDx
QSCbqSZIsbIwwKNCCfn77Kvv9dcbMAWQWIgKW8dN7F5959OhmJYuGMbia8a4JwAd
BV5zcHcrHRSvtVePBBcjGkmltUzRTiE2Z/aIvM+DBvz/0xaDYQW4dnZLMCie9GC6
WQtye7hy0BqPGlUw0RScK3CRGdYFoAJjENdFD62pZ6OeYa+M7r16cCPqVTdohtMM
5cr2dM9eCFje+WtfR9QgRP6JZoI7LBbrogsOfX7pZwOvieiTncRzMBoRdaxe4A5A
0kx5wEC3W0NRAVNxqE1R37qgcX6N4H/YIsbIpmkUZVuhj1t5tGrS5kdHj2ZqQaN/
RYJUDLX87CV3u/nQkeA0FKsoHTIf93pHi0xS8RI7NhzlQBA0TSO795hRtm14rN1h
kfb64TnN146fq/QglJR2rkKFTYh92xOSQJ/+3joUhyitqzhYlcdhWCZWAHYhY8Ux
5aPjJWEqNnQu+dZ8xjP9L59UeHpkyzwzRpu4DQ/wCR7DzwxSBvP0TLa20C1bAsC0
r++lgXkkycFhBnC6aX4eGO0H5M7EqMXmGIrGpiQWlesdstZdoC8CpMxHYWJQzj7f
0tcbtuGuXvKaCw14VCJXUHWa2Umk5qfzrZAZD+0gQsj2TiAKMf4zJdfisrzfBbs3
SWNbfAhmSA79YzaJgGjMyTULPYew0BrkPbVmmPFF0+K6qHoXb1yWD9+8+rDimb/3
S4j0hvTTU1srjtI/VuRrakneD/bpJ6kSz0l1jQ2tSmvAuK4IOHDWSnm1mU8hbAFv
OMXKUxOiALoyva25TVj+ja4doxR+DsYaCgoHNNSGjFId8pKBdi6Ozu9V8xvNBN6X
e95fUrKF95Q672BJ2+pjwCPUrcb88/0EQTNZJa0N5v8hWzSnAi6Ew50/Mwrkm+5S
UwKScOy99yqv8jLl6XJcvtd5eSu9OTMKZgP9BBYdY0ae19tTDGeuFAQNtoBgFPdN
kuPalC8mPtyWqLeEHPOS9u94alYd+lvpcf2yIn+ODsDdyJvTTjk28FrbC2+bXRSd
b05uG8ayPaxrRCkhIOeGs+2EdNTqsW/lMu1YUpbOhapzILkWDT7VJLOLwcL9zOpr
rhe3Y7wgGrxT4wo06fC61j9aLe0AVXj+KQWmVQzcv42ZHYMYcgtAodaQ/bmvdhMz
slcXN2kw6ExAdHUE5gazKgKTXXV6v4Z13ilKZL60oh3XBHhq0XlW9VnuFUKIObK4
3PeczFFXyzjBNl2G2Jgz18l3PZk1U90yI6T4I5VHQhv8QDPb4rxv4FUeykLzJslH
KWFvlFhThQ8knN69XVw/49aourTkTpInKuVJQPxrxzQKiiDOBCJtxeA0dAuKLbNw
SFe3gEytcg/HBchQXn7Ik6ZcZ/kuwp9SiZOnVozvHoWJX99IoDfrQUQdaMwWBlnu
yzo24so+gPXVRscMQ9XYcdhixkeeHCD1N7RAOpwqKoIDSfQcAu9tdPi+cWERS23Q
w1JeTnyzJA5V7k85I/RfWtrJo4ZIocsyPcu8P2yWz+lxhz0LeyDnEqbs/hWKssZX
RuMtljpH5EQgxPfO4gRiFxCeLv/vi8Fnx2tvLEmAIszWGlGNv/qWBQ/lw5tfS/hE
LJWPTzewOGgXnKYvydgtrBMQ8pK0aQBP84mVyJkkkF3ddpJ+YC4P90hfxVZ0Iy+5
vgFsyKCxWnOpUU5xc4CtdVXSB8oV+WAn5hNfVTEMYWOeMqD5gKc/+7gsc9wryGwq
l4u+iJ2HmiAOLS8ZHJ/O8BVnNLCU43DoTI/Kmzywk4Z/FONHq49IzY2tIm9d1B6f
cxShYWQ4RtNCW6Cg6sE0mA/r/DFpC6U50VpboGSxAs+4xnlF4p0nni/fqWeE1uF3
odpOYrjwINKDXbQAkJ9p6s0HKwi3HO4S4hhSTV/fqkgM+u0tlrR7FYcJeQWeEtv3
Qj8qtbdIqFm2Ikas5VdKd0EUyqmLqVwpFKhk4KMWk2NAqAIiwLwliNX9Z3vVnA+5
8tqx9obkBvCYBFaMNCpQdAEpywwaddnAN8f2BYPNSSxisEXuP50hgMKyQeve4qmt
kemhnTUKECNZEH6Tm8jsesGCT/wVQlSwuCAC0Cwu5kAUTm77EfRyoLilm2xKusLO
nkSBCH2oowwIm89JEk9C1vr/q9NtOglkbhe3owqGPSN0iekJxKgEOpT/8thzaKQt
cxEd6TWwxeRMkhI7LO9Dn0KgOltSGlqx4iUPH+cNpL2kT2SYb5bfK59I8n4oYcs6
1nZ1tknZwVEJY/93PpN/chVyDoLCSee3WgCj8XDZf4nCyf8MrvNXTvQmh28ZcenA
SES+24Bpgs6z+U/iCBFnlZpGkEqShVvgKgaFi/fjOzvqWYCjvwNWn+Dp0KkH1uqs
rICRmrDgEjr9VRK6gVvQBPfyxrxIOWBujhgMymlbQwfrk/GEhornr+0Td8XC/SBn
z1fUgQjSm4HOQIjcJugja0NPitfzgw7s8xf6wuhKo4PZwEhP6cATCOCDy6DU11Xd
/0T7sQceBhCwYHOHuR45LS7H9Ddr1SQNRveptuM7O8g5KU3reN5n/SLzN9QkswTU
Ew3R4aPMDCZWBlAX/I4qjDe+DvKewCSU3fGvpSHjtEpJosISQraNxdApr9DVoGi+
UzB0KKztLUg1e1gCA6ea1KyB8WrqCautFwJwMev2dmEyQtBl6X8H9tWLociyDyIj
WHGjTCJDlAgRzOcaro4KPW3OR/7J06qCc/zZCur86jDQImDZIpEUj61RVzNWZJgL
l0za+YHj5223LWv6NfWl8i4M1duyh5lEbu9CKyZ8hqt9Bih+J3d1xnYndURjgBEK
6Fd5ZFSPbJvZ3m7MVEOQNCWVuQvNd7huEyU9A8d+WOT95/fCiT4jsBfSNszhQBQC
KGoF4YE39SCRE4jpE4FO4/h/ipQn/9zQOZiufLIrRsilhLUIheC8/IlkqADkgvLy
s3OHLlnFC6E233uBZ7Ada2p18TH+W90rvs1dIdIvFc02jnViMHZITaYNyTYMGB5i
D5Y1rwjrClkikF0qTvuSJSSJbe9Z9jMpTnFqthQhUSIekb/OgElqyORWE9+e27pn
UCApNquSUSNaSFrOwlfGLV9xhwujo+xnWJJqVK4cdiHADvKwsjtBS7P5ARvnxvea
Ht2RP3pl/Bkkg3CM5ijlJRBPl9ZSNYIg4sKI8+tsAb2TiKL2LOYAkormFTmfuuwj
r83S0yqXa6017ZA3s3W1K4sMm6Ksy72TNSabgSbtaam4P4TWhLn1id0fjoeSmFS+
X7hZgRWPoIgeR6VR8cu6+POMfZ1xL6lS/aWIwHhTOVh3dvNDNu++q0zB7xuLwwie
VtCrKRd4TRS6G00P6EggEKgYSa6wZx3WlUX3Vm1vMU5E4ZFDwll+jJXMxnXb3Mgf
RZiZZRZP7Rw4qX3/EFf2jF1+qHYmrqBb6Q36lViPr/1iA1iLNJMDnrcfGcFVSPf0
iShsbtXOSAY+Kv4T+cqYlFzicOdZufp1uVh60sEe0LjmTWQj7gIVbAr7lC0J8FXo
a10cQgFwYwA6zFY8agvp9Ag8FfnhKeSVK+ipwX2ZHwWE4RtygLi8xShripXdJw2h
HlZ6dL7DKQd4YspJNlcIopgFkS1NkEZb2H4vNtLQMepYTa6zsnQZjgwlvs/6qDVL
MPM9mcbVf6UQaxh/SPLEVygWFf/SfT9KRt3EmM+/YAJQ6R/ynMGDGeFe/KTgT9Nj
tn6bqNsWdFB4wgjqDY2AhQK+3VFTRNr7DYqM5pvvM4K21oI+f2uedQ7JoQ80nYI6
CJfxi8Zz71UPKTfP10SNByhwcwW/s2M+AhOI2Z4ulNMe2Yi/f07f+b/fUlTTc7fQ
wZwyNGk5vQgCRTSnNeHkP2bwm3NWZ5ueBAXGTHek+sFoqLuZiVJ4c1vP/7xmGkDg
WCczlAOm2t4gFyrXBWTGXaf/k+QxnktQyfQiKFElB+Zha0oOIt8SqIhQpSn1NtJB
RwXe6nvQcdV+NsGbuSKb3eA7la/23uAhgnEqp32kdM9unOU/RL6R8cSPXOgTJBR1
pMWUBzLsdZnBLijrEN9twQg3aFH3hCB8jNe/JAE46rSq9paqa56XnbPGmG9aZzbu
0hD/br08EiFfbwh1NdH7tDkuZFYVGAgqtJGXaBg9oL8YAS7/UgiNk6LXWKHurEf6
9v9oVkbiWt60P5CsaMn3Fj1SbqJ973iV9kkqOX2i2/HU5ojc1AT+cLHNk7h37L7C
wYiYfMuZRQECcJU/6doGyDHrqaI4KADkfvYaU7xkmPjhKpssOE1r9cmT5aiLpqCx
+qGi2FUJyHDERwBOGCUMWbws1yPfRquwE1tRewmtlS7WGSn5UOYPUrOCKmBvwjt2
Fzp6g0gKDCpOErPVP0ii3Hrc573IbcDTDE4ODwxS1NNN1jkQ7TvP7QQ4K6aW+Y5W
+C2x1fnY/QFfTnUjlxBXMzhtf3IJyDHCDCTQMIstKCDhhYaYrNYo9HIhIxzB5+95
7kS4aq/GVHZcRsi/sdT51Mnc7/9jjHsQ7jbO6ICDzSeWzsyjyY5b6PBAi+cSglhS
/0+aGOKCMWDYZiYj0skwV1Ap3WMslUY8ZVYG++G8H7KPxgM4lBXqWZ7GMiIK7WHs
krr/oKcSgr9OHMbJdAJFztvT0bSnhwUNlLk4OiTnBPUVNXirvY6gUNgj0IbayhYu
mxqASqhUfbZX9ERMYeal0tex+bqGq6z5EeaGskcSvnix05DrUn7zljKB+No+Br9d
nBuOOQ/3sFa6j0MKzbl72GnxbGnJZJM3TC+Yzbie16M/MAmrsYImsjJPkL6Ljjb0
cFONe4LXFcxKHNjKcaK3os9HiRkwNFvP3nOwNNzNoqAIVTRyjmrkjHtchQMVofeC
SnR9Q3ipfBiyjYyfqlHpH3OH9JdkQb20NoItH0+xWV+Y8ROELwOjtvEDQqHST8ON
FplUrX0xEfsl9754xAVPHez/qdL6ol/zQ5uCKEeWzx9v8HjUAogoWmlI3Go2/6uF
8/f6Eh0nRapKM8flY5delYUSAcBq9kLtoi+TeFguFM1rtrvgdt6nENjAPT0bJ1lg
879hA4hePFE/mWINg0KveSsBP9IAgCSn8LMuo7RJdbMP5CapX+4nmSN5REiR0X3O
sFXQeP3a0Tu8gPe8sP5eKoXXgRbePLpGPPKfMCdUtdgntu076HDLLh/ho+T0v5Cr
lc+H3iNpH9MqxwD+XFsINBQcwkAMNmVdgGXXH8dAE0oUUNwJBqlp0ri11l523nCB
UM08WG8IaxShSq6lcyLf0dvrBj3NKts36MUp/VlgGLhVNMMc31mSb+Vp8vlMnFZJ
rey/YORkTqto/ER2SpMozeoBLePWSC8cO/hBUj9vsNG0qI1rd1wNrKC/3mVVa6gp
RERZPf6fep7zu8pdYqf6vpE5iN7i94lN3VgZhlRnF/+szQL+qaE3tYnfJnOzvcbC
8aQtvpEdRUs2Bh5pJtOJJZIv/ySpwL9PeGpXl1qU4as237K52gSRvoJSlIl6RXLp
djHQGy8w5Of5DVghKnqAbh2wqUzp+470rgFsxsfzbPdtU4cxsxYlJ8PgaOfxLymc
9VRSc4QS9pCboKja7seWT+MFNuaLVY0ZzGEt8sAl3aOMwBjHjPulVjYf8S5/sKxQ
t4j7T9/YUWuE0FtDhGq3WNuBFY/gyvizKJINopbGgU80s/Glyr86jeYmqOGxtS3J
A4iQbZTkRycw4MKHz71arfDzyIC1lTgx5okAlSqQwyJ/KvbBKFIIAJBLt4tCfWR3
kecr1INhMHpId20j5CMZNetSrF44IIfzaKVPIlpFkfCbHqVXy6dnv3L1KeTYN1Ye
oDknptpjyoHmb7ZbwOQu8IUcrRTV1+IRW+Nsv4e5ampXcXk8BP35Zn4ZTpxPlavj
rbvw5qe4TuSXP7eCHEgPKjRJaIPxgyr71UIlzgDVYsZoQfXItyVTjtOM5d7iYYiM
oRg5I40UsJNpLW2l1+q4LfX1mCYU3cN+rPbu7ByMOYg7nsOPHpcZc3x9MtjeaoF+
CSJR6MCe+9/rFOop5DvjVvZaSb3hTx1BinQP2IO9p5Ag4MstS+1M2tCHiz8qabon
m8XCVS7GloKFqPQRYLmPQUkmDBhPbHcrMUgqcp006K6x/Fy49xo33foZKP0CtFD5
4KBZVSZXqAplF43+de8DZDB9HsxZ+7R9m+gG1x8q5HtLDqAp3fWOHcB7nItq1Lvt
zpqvg0xdOkgphIGEEWMjalofC/BEFp3b45qPiGAKsJd/NgUCMJf7xfMYaqLG9+TG
aXpsMTONQt9ERn87bksdOO3m6fPOIP1h80Id8zL9TdQZ8lZQ+ntOsiZZ+kOnVLIL
0jPvq7F1f2F/Na3tX+iujiQnOXC+cDEaxmSQrfMOjpZh/ssgCdYCDcGwXoX4nQ+i
5QsrebFnyVKpiq1H5aEkJ75tU8lHRrPRm4zDaFh+KkuAwVxfxJwemLoTykQQJt9X
9sThRpbn5W4HmcIidg8WL9EtAvjJd+TEdv8DVDgcO5opDmuT0GrirB7PK02HYHYx
KQgJTrTLPF9SH19UWLzLnj0Fh5GXeP0D48S8VV3t8iZZhwC5VYFsInhkFx7C04JL
qo3kOXpVuBci8Lfk0g6vS6LUM8MGWvHbv6Ybpa5DIDZOLKKk8tSzkQYAnbt8nfwc
eciTg1h159tdRlTMT/1iNepKP4hk4tvYXfu5DdyvVJqNYDme71MbRliZaKuhajH3
Eop3l9v88S3ejEn3NbHEN6ItPBwUS6Iz/vIbE1Ok02ivi+Lj6R5uJfpCl0qDR8wI
BTvQqdE1HDdo/17upgurCE/SB3TjMdMlp/y3YQj/wC0G+gKIfqS+pr7aUobUJohE
ktZr1HZwdvyqlv8Gl4PFrvbP9EmEq3FOJ16OUWuqtbPs3rMHEyEkuts9PoimrBM5
r2GkPYi7QYIprWbQJqoi6qkr4CJUsOPy6Ar9/8HWUHQ6WYwTvDYbkFcefhA6tcwk
b590fRB9yOtnexosAncD9ah/76ykWof6f+L0Ude/oBXDD+hG4mca/vpIR+rAc3VA
Cw2Zdti7p0rWMMRxYP1xYuJnXb/MwpXO2D1BLp982m6ORrAw+fSXo1sypn97M2SP
hhxw9ETEHaT022qjFdiTE7MAdDKnVlaqSeLpD74bHD5lpaHuioz4L8MsP3qbz2SE
ZCiLc/EBpjjKWVtX1FlXoxTjSOUKoeWf62uVct/hskuziKx73cxcCF2yg9OMxfMh
Wjw25NBR0TZJFwvZ/7K2jnk95MdEgT0l5pv7l/nakv03yl0Ri8nGYnoYE3n9IYvD
Ktq8Vpnraif8QhFluGNS4f76Fe+ust/B39TrWiZHj4aPbD+b64/ws+EuKc0VYfM2
+w86l+bDdUjliLpZfMqyqZNOvVP1o2bFUO/TYm5JzrSnk4IYGo73LNK3fga3MBEc
fRI1uh+BoKSKExIRWd+/1DqAxiW1CSNLEEmZ1h1tFV71o6LDOfRBOPwhUe1KE8Eb
OuT+O46xDCYyZB16vkFnj689koy2BGoqBa0e3IH2gRxTkv0AlRDlpaXEa4GULabw
/AbFHNYAsdxg3ISBXds1FTv2cSKRIdY2JRedeYcy3PQSTfGT1qgxpeyPQ81ayPnE
Zc9dAg9361K0lpQ4MSoKlkwAh49zBzM9j7bvgayGqYd/zpoJqJBrs4Z7+jynO+Yb
HHq0t7RcqZdlmD+RNg64Q+wKpc80YhlBFkuhursZ6DYp8oOWiSchzLGjfScjmPHI
G+z2Ck1eEqPPHr7WMm+xTAl17ntG48uqiwgtdDo5Kr6/enZltztirET41eaY99Xy
dku4Ct83I7I+tBWpuYHKD863g1XEn8Y/6sP12RydHfybW3F0TWTguJ5qXDBXpL7K
XdejFHUa/TJb9TLkC35s8lhGKXtPkGtq6PRKH4czrIAVHBsRuJbgTqG8Zr4sNm+1
3Fs4xjht5PfpqRBwHVs356BnQWova235KNQxFvulG4t7z1kZuug+i7hGwvehvIGZ
iyZ+Pg9B+zKhDrzv7WQTfJ8XiP4Esoy0lVInGxhe8g5Iq0p03o/x0f8aKgqpxAP/
RHh/QOgu1IjMF7iVJ92rRKWVtav/BgCJItxMm39eUEIq4DlaAOUAmL2L0TEHUaCj
pNZYDXHnw1zR585Nb2wLFngORGXVginlA1wKBlMQ6J+fq3O/MqYIByG6hrjpiAah
o1oJFvs8lvgGSRnAVhxUsq12fP/uuIknNhMSekeF7jGXGPyyn08rCLccaXz6Mgx2
gZexhqzeFbPfdbIhsePyyn2FloHwK4kuMJbVrB3LPmfINy3ZqwCJwrGLWkQq2zeT
1JjMuDL5KdyKGmdWMelE+3XLHvOX8gSMmbwo50zN0AalHvRa6bj44+2PsbrFihcq
lLjSr/JGerA4fRcPhLnuo2ENIbtxXYJrK4CmWEPGsweewePmJpPaYQcQGznaX8MO
clvDVtRi153V1/W0FzvtAv/xKLLC464XXMVHH4TDL3xbzx/1kfg+v9nwOt6D15Z8
WesD10m+2avCs5WXZchnYEroJz3JpL8+5dl3IU5eSGJUt/UnlVoZW5ymaxoIrDaY
bq+nEyeDbbPN8Qa27Ad5+ZOdbhyOHWEQYL4K2Prs4EylCXnnhX6F1r5H/wRD5Upu
0YidqtkO1O/bd6e3I50jxg82sLaeA+jh7Ap/fMRZD4CpUJCsYZMPL2sq4Tqr4/fV
GujaO3McjwZ1kMTSi+2w7JmR9V+Qe7x6AD7bfytZ9FeGdxaOhQcIGrfFMM5DhM36
KSBguIHmqIZLeO0bQsDUKhK2WtA41VgK+8unQ6euRFIP0dK+Q/LYm7869J/XrLTx
vatta7pPBe66IBVog8tslmI22GBZkxGKdnh7Xs6Tidu4+PO3IwKHh75jH3z4SvTN
yq4fkDbkTS7lC/d6kbFqsYsAnKBByGkaw0Ky0A9yB/twYrjKlHsLy7K9DP1RHwGm
6tfB8WQAnXuvEXpSXhdGj68kbUDxlsGLE4K8I9qwaoTVdfEVV3tzBmpcy3C3sKNk
kEmdUGEeDwFP9vnPW9dHEB4nexPSSOChjt1FNyHrryfkeGs0+qiQyXcc7yuD0qqZ
q3Ws1BnqVa3OEi6qcHdukRrQBVDmRfyRZQUZtBt6ih6Umxhs6XGqUHuG7JdRphiB
gojnoFRrAWiYvEPdkbh5AxicQza5gRnNAU6aZEne6tSJmCf5pD6OtqmUc8gVz4xW
rDoElDZ3jZM571IlHxAw8VcJd/+DDIVFQtuALFgegT8F7KX89cKM6nhemc3rIDLH
RsABsdcOQuw8P3/jkb7R07NCKYtOtSL3oHYjyVjTc3TG1OxuSfGq/V8T8u5KuSkg
99yaPWF3Zfp/77XV/8mGL3GVNkDDPCYP09wRgutfA7LcQqZH9J20Uptuq80+eHt4
Aiykgv8/AGW+8oR/wXY9+gOSgpDi0YnBBrAiYFgJvapHD5iK4EaKKR+EVxPbGf/Y
K555fJmVFiI4P7zBjwjICh5hp8pemd7JB4+eiTWCfiCKRPvXiMXDikcAU/79KQHu
u7/4JGMy/H/VJgqeFX63JttrV4yYznFRd93ujdG+h3GLTiOnunYGRin4ObyBdxcL
iOga0fbOA9iqOrC9xvgzM66BEz9w93CQPBFmPeLdl4ClCWB+IAgWRvSDjW5uZ6ws
4qVUe+yka8jBa4hXirNA7azHrwOJ9VqPS7WJBD0ZTlF5MWoaTJjcITx2pe2qgQ1F
YgaH5pbz9aV7+gMl3eU6Jldb8AUg8zryMJog8S9KNEJqHgeAMHUim/cLms1ZFOnc
4DUShdHG2cLS0LZNkZDiXLrOnA+GOZ4l3l5KW6hMuJagUGyeJYK3uDkGal2pR0VY
eseNWSu3/COS7QaJAYYmO32WwpPFn6WLpEca8XWyfW+eLjjOYtKCGIdtag7fioyN
xIvTY/CtrhTiLyJZPsPJXFycHZPB064jetg0en8csvJqfrVOpVAqYz7JiZ4KjzsI
ZI9HHHO5Pl4vC5c1mSgRWMiB/7DYHgA1osGsIEJ2vcM5KLYjwTEoGgGEQqyzO3XR
hdFaSVyV1hdBt7ZL9Md9AmhpOV0hblTfEillQTxp8Zd6QtfOK+e1qdPGBFwYSCFE
Sv8/cp5hdoGXQS2zIvHMkWFWORiVSiNzbYdpJQz5LnUmt9wl+LtlyDb6IMYZwPOA
2muly5PhuX6Rtoc1rDqpVOlmvEOYFzrHF8q+Dh5BeghYY1wG/BowgpzCt+bcCGMB
RsiS0PrxFFe/3mjam7qt3c5CdIkvTGLv/CWtGwThUOn0rx09PuR91o7LdV08Y8hI
9v6pOtF9I97uA8vEb4ukuSx8jqhkEwroXBbrej/PwAcyqxkatjZK0TTKPQ8bOMnv
yjZ0z6X8UGfBwsJddHGZ/ZX9t87kcFc7RnySnYX515g2PGmHWkrQoN+8UjdS+YUW
KlB4wQ5Te4m8z773D2NmTi3ZHHP8PbLkHTrI//yNhGuma0dGX7Ej3GalUpcwPqls
Km5pzT2ztoVuoSWMYr/agFRbW8MZrUkFvzQhNp595B9wBihQpbP9ewCC0GFFF9H6
zw4LeiV84fTafEYZm9EABvxBKJvmnV0u8AsOCtdjdO6pqo1dhU58OAq++Ybhn/6W
kdjk8ExcPBf46oe1y4IzSOQsnbWd80A1toiylnDuzPidXyMxh8SUok63aDYCyy14
c/TfOUOPT8YCrD14tUeuWa0MpytBPZ7+lxdpMCtyvc/pCiCnbcFdkPluWcOSGShb
4VZIU218GZYv+dVk+5cd6vk2pVdYrfB0EVsr4hUoLSYBitl2J4zMkvfMKBl4j1d7
R6W3NYo5KyLk3TvwqlhwfErykCVJqyQu76iVw8p5DMgXHeZ/j7lpdbEg6Y9FSmGb
flE79s5wBqfg//4utGCunR89CjgufO4CWOBUV9iVtWxBtBEO6iSxuAz5omVqZZLG
W7akWb1iiI4HeWZztkIXkkrIsmnpcOL11ylY+TViwUdtTt0qysAQM6Iq03/y9BmE
JLlPLjXYLcdLNg1oOxDsjZ7plzWj0RQRNF5xJQk27EiHR4tBbOe/SRrzhpjnR/U0
bD7TSmzCrubs4SvMbIJdJyu1KwNt03nlsfSrnSKI6tv5IYhcrsoN2y9GG+XRrlSW
ZpsI+PfSVwzagdcFDz1bc0sh6puZCnbM4cfPtdWCJHEaP0vm/lK0m5gl8mvZ4qnD
5qSaTdHZS0FRBwGwJQd7vYRJnjwWNqHkZnMspg8RIjX17QbZu0a8PX4I2yIaWQGc
pHo3Lb8db4ekXPYbBXDS1N6w5zOUwLJhNy1RnFhOOASoTjRggN01uKw/GluEjkKV
SCavACVnXAUZbu3JYul8MXwFBLDKqPxTbNkrk0ytKY3jgelJIPkzDVRnSMQ2d0uK
m9OoU3XxonRHfW/CfVUB+3mvQznYwFL6IqMSi8H0Ub5Ga0Y/BnEr7a/7lfHD5wFb
AJNAsExhUqBCKML0xEtULT+zNu8/N6avoZNtTW8XnKkes0GeW7TWmVfFvc0q4Jse
Uzi+z3aTTm3P4jyxG42M1wgrfqHmqZCgZGlk9Eb8ENGnuCfaMA7cMiTi83I1ZqWM
yKRLwjWNzlUfbaB0TNLve9NEVvKRoohAndTwazp8zT+P3HEKHsLtBotojc+Q9uoJ
8OVtGMi98GJaxMm2rkbcl5jluLCBQ9ou/7+BHyOOgNbg/hJoWPK/6Kok1zzi1kuY
rcZ7iPsszkYyqwr5H8nsuRMswjk4hl+qtuUNK3nInk2tNGc57f8xjYwPYhIN8wJ4
8NlJOKU2e8lbPz3O3yzKYYsf0rMme8JVVWNHTGmzpSMZC33FKcNIh1dMrHV6Cl/8
mu/vUmXOLuxnxm3x9wAmzrhAO7o88EqFRt940wQc4l8QQAJeHPE33KGUzCCCqSva
2sqZ42FNa+82JzIQXXkMPLgkuYKnIZsewkzTnmx0WGG6nU18bea+rqn5Ky0Q2fq0
zR5/blF7Jrsdu5ZXt3zh71SVZwqKkXwRiXHyVxFCU1NWnLf/6Ift8wpt2kOgeGV2
ypHsAsxjppCB+0B9zhAzLPhXggKZYUEYFuT90T9UVHeTaVolzUdXGn8xG9frXb5U
ET3chNqZy5Wr8txge65F2clYkPy/fwwyvWzwVgq3UyB/Gqu7GnKBj+ZKLbx6jLpk
7SuAwIzbmOWs4HxKLnshnsWXlCc+LTKxuwAZ8QWfDmrKFZq2wDEZXI9FeyAMVGoK
p9flubk80IDtuxrQ3i5dhkg9q2mq0VFjspZ3PVQyuLkc38LsP77px2E5o387WW6x
SgJ16+dZD/pIBn7Oax5K4uazxoc72vjdEA1ELWpoWnFLE+64eiFQWrHu2OhMeHdz
vxpMMpDheUuM5vMa/LES7EZZRQorHWvwXeYIgE6VG1dZpYMmnOK4I6CHP0tiRXe/
dnZfKAvS+2Mhcp+PWH8dTDOlxRLO/Dzi78LvYBC+arprXL5R+t2Yju7MdYjkmyq8
r/MV9ZuqWvMp7VJ6sCWqPOjWbE7dVmRcEySH63J7vqPJVEhje46eQZwWvoveZ+lD
ftWKnxg6AgAY7v4lUI5yVYntey4vS7LQ/JLU3Xtmetc9OMco7Pj8GjC1lrmW/Vvw
lDez7H5oTdVVCVCoxKx1jeNJXasHCX7ARQBiDUywLzhr0DdmB/epBzTTn7v/ql4H
4wCQdxkTYYWS9mo4U3HuQs8mRAO6J9gDY0lP07AmY5xww4DQYeEc0f66YO/lUXoO
ZeQ4hOUdC303sxOSUm75liKAJIwsEeVHI+jNKSEyEwkqrLjhlafz7LW8+ZKllb8i
Yhln1AchUVnQPBsybGeEJS4OMWnwE8HgQrvmpm61IEaPMFwSDrRIIQzf2qCulWdf
rDywMCF1Uiz9FFmDtrELzqdOWvkwk0RAotduyd938wJEEX3imkWFiebHt8NwIF+J
zy/KDPQLOg8JaPgfcS4yiVO0C12kmer5DvGEZtIV9obIpCxG0nkONyd67OaI/fZq
Zg5t7xb6zBL9DypaXozJBlmOPdCnk6kGMXunTMY0WB4+VS9DP8I8buzjnzXnq9cL
Q1toEZAnqPDFREgCwvCc53WaJPvv1RMH17VIhmMuAGnolqsocGsuGqodRl3wYlCj
/TxC/lOe/1wujwB3w2FfPUUP3bc54vT5evexMbRQ3Y1QE+Ag9qSoR4yJ+TGKbDEX
7AYCAxqYNAsDmjG1aZ+KpRf6tZVZmykl01ZShDIOZLD4bWdFSM6twVq+7FI0f9Pr
PocwYxS1jj0p3N7iVMkZovlHf6i+WtAIkzFD7EfTA5LCk7CKCJfCS0xZY9GewsPT
6mC6D1rUZdsf0W610eBhzWyu1xOcBmJ3e3kbMjBSJpVnuf6CCGW5etfrTAUeofji
sEPXUJd+WeuGH2DSwWpo9iw2qOLdIFc04T5GN+v/7M8cc6n6KMGJReUOryz8sO3C
bfqpLNfE4xLAPSI8T3A+jd1S5nAXZ4HFucOr7lt3iU/dtBXOD5UUDH9nKnprXoGr
Zh9kxICDm/5zuoYby+pdV6pzs3p/yU0g81yqNWIEbEmxAXwtnDcX9oc3AgTsLlR3
eGG/KKGR+rYpiLyaS2BnJNDKhGzme2kbgQ7EICzI1JRYN/eBCbd6RVTuMeVN6Gu5
mm1gjR5rKib2r0TGFMwV7K+t7Bx+DDZrgS28kD0WHEmucCfz+j8C8B12K8kULDTZ
GgoOBOn/rZFxlzLLKM6c1xTxWo58nPZGD+90BmG1Fbiv1mPn4uy0zTkUcfbJU0yV
+Dr+/+LzOkKqGcSNr7iJfPmkVmqRZ6c1TGNVtPauwcsKnmxrxTXjuq7pXzcnXOO8
f2ONEOapzqRnxk7w/l1vlQ2TOnvNtMQLPHiEW0xDAdo/C+HNjIkWMKTOG/5bTZpJ
D0kbcZYgDKQQqFiF8sQovM1CluVof2cqu996ltvOBit+U2UM3sV7rtEZ8907xsbn
Aw+sq6ZYD9Y0Vvnp8ECPY6PDE4DaOspcWvfzsI6ISNy5678G4ocxse9WbRnqcV24
r+Kk3mGHz0F4/6/iL4y85tsYqEcDtizwl66xKqwgbwqJACtSnksSy/TqsNZDobAE
OO7Om8X8KRMgYpbMdkZOR1HBvdG3XP4uErGVzzfedYCCoEE1qPagygDs/fIiOecC
8wfapRIJxVt5nxQVMfj/LE5sHRhnJcTYxXYKP++Lc7+GELFYu+zvWlq/FNE5i6r8
+ekW5iHJamC+v0xxZn2hSvPz36436EwTDye7L8NraDT+eAR4RzSRQCKNqIDhHVOP
z/Yd+mzq7dlVFI5YDrxyztKSVscJbu36IE1Xm3Ms/kBwqJVvkoXz90L+TPX+zx84
gQ6Lk2FrUFUYsiJ7RID3l/NBNGah7QZCtHJm3uEKdXnH9IfHVDes2MPY1vD6Q6km
mqtZnkXlYuKoKAIuXtlkV+WQGC9XZ5AMJlJiukn0Xdf79N21DxmRK/fpLNNu4/8Y
6NzZ/qYaUSFteCb9rjs3f5Ofr1ZdKWLt4G3nijgVehCkPw/CVS35pUjKHZr7tLfS
rZuqZGLWKZ8ZhYD/cu4o9wnvB3qj4/k74A6FgaW9hxjYqqx0KziG4SJ027hOn46W
PnZruq2iE87fxt+BzPt+AoO2WvaBmZKfmfmjFqQYchJPm6iZEn4xt3tnS8F9ZJLR
Oaj6OUYnZ/orp7RBy9z9RnUDGKqSFos22GPb5wOWh/TKqn5N9AqPYoysrvkSVlOX
RmuWLUiINMQMIp9DHgpQ/X75nQkGAt5ceDK9NbMiyoVAlnGNsp2iKplfNuIe8iDp
f3x+QL5QNuTRX7lLKv+ri2hemuZzSOXwk7cbE6MP9cWYPXygx0N7KqhwsyjmyCEC
xrx2cY86nNe5vyShgYpGK6OrvSUwRLXTudMgnjXl+IgniEhNTLEnJA3UfDa4pF7/
54h7preuP3WwcjzltH4qd13yXGnNlDCpAjySvoJ/Xx/GTYeDWL0TaqZwQG+G8Bf3
aSzYPtCO5FbcqNeoNKr0Z5pn8MT5ya7iAYWrbonZyxfiegaFF1kY4NDIkLwMKLMf
IrSYY98Xs+keK6YT/JfU47s8Ace5jp0UUV25dMH4yd7aQb2bIIqNgmsTLzaYfZSb
uz8PKZ81dhk9kdkluuFV3cyPgmOMz3F7PgH/MP3kCSLQut0RrXLh0ZDldHjCrWhy
HE8SbRjFAQfcLUtO1IWQgCDn0m/GLZ1y//5ssX0zNpZM4pQDlnYcpFWT7qYNFV5M
hJSnVZSZX8UcC1uwjgOBUMFl18Qu+oZSSof4G86TxMlLFyQtDeNXa5Y/TGnZrXUX
pVvNtnXTG9rm3rRlaiuIOtENZjrm708icsSOa/GUWIKp9vTTPj0CNtgWloI5Y14S
Dk72HoPmgtUq1llFj5E9N6nXRWOBMv+uZvHwF1gMjJBNpVyevzRVzekf9K4vXZYZ
beT+ZBaPm6kLE4cx3qXFPvgGlGGTNRceG4iujHmRJ/N23oB5CqhGtMlr3qZoDXUA
/ZXDfxCvxIgQKzMozB8UqvpVSrxESxUNl2LElOzOBG1WZfb9lqz1hJ0TQksoS41Y
Qn6+xZw9VIli2F2S2GNYAgjd7xoVrB//Ke16NlqCMrVvuhR4fhON2XXZVY8RJJ5R
HS35RayDoonJf8L17njQHfUErdkZiv8HcT5pm8CexNmkhtUQ+DToJ1CoXIeoUGg+
Tetpn0V8Fkca883aieukx67UnO1hZv7h+ZPcfT+X1U3jeVe252uhecMd3ZQYF8Ko
Dl8HeMTfPxm1zkDcj6b4U3SkGhOSwuikFCqaDvGB3YdOrTzM+UKeglEzgR/mmDYc
GfLRTSsw9lxMYoWzwY71GS6J3XWi3Ahtg5ZaNaUrJ5q9L+x/TKjqJIZ4+lBEubHe
LaLIV3g5vnk04e6wqFn7GSKBeEGpJ+Cy9RNcUt+9IKxwsep5/q0CId0lnh6YRzgA
z2kbB/ZJmw5y/wy0kNB0C1FumfWwnVUEbhYIvh6uyYDfoQT2VHH9Ln8vT7FZj5Mg
8+BheN0A1ZlkOphJiWSUYHnh9dEA7TIuH9UqvWtq8AbdWzEfjzz+E0RVZ+XXS8k1
j0Qk4celDC33aNcB5h/03IET2MCZhCw1r9HQsYILnJk2s2QRyw5T1J7gEH0RZD2P
v60ixVO9ukI23YguMEU8WWnJtUMMugD9u+aM6xdnNuaxr5Agqm4tpdwee0hjHPWG
qWRyJ2T68cDoDkm0fizxLMX0G9nANiwQ6jFUfJ7fo2iAe21145bA0LwMxoBc+taG
caDIn0ZXoQADhO6wOfspQZfCNw/lBzMitGsMjr18QondbQFkFaPKPq1TFPHxfiU/
hxN1VjLNvkiJ180aPkpDoeeNASsVOzqB/GI19eqfHtOEtzmyUjzI0XTKL4QJHbug
9sUunB6daT+Py34MAIdPsummgXBoakHXNKrq4i7tSK7KtvBQx5qvF65389swiVYe
+jQ5oERsw5VGkrCVoFM9qJ6cV+voQuHJ361rX1FFSqIzlbUl+mL8ZrAYTpLG1wiq
1ghoKL0HRH3v+KSln2UBmtTnoeDVkHOriFdpcmfKqhOu+HleRQ//jpwcVoP20Vtm
ZFV6oOG4YI9uAZftfPrA2kiLihbwPpM70WJ+d9PGUoUHFiH9gJLN4YDVGZ3LwfIS
DIWKzpkSsqjNOL47cuYYU00C7Em6UVxo/hThftVN0ciKlAN/6VB1oaPae41o0pxH
Wbc+Uqup6FeBY8H3jryHQ+xUIEk7cRAZa2yGVikyKlpvcVWQamtPxo3khGXS/BFT
5eYZgEN04q851datOoOjElT0p8GVjMBDJSSlmZZV4GwawH8MO9IuUr6iVfC0L11R
V5moOicE15Dk5Q01twf533bWP1RePmsYfR/vBChc1MtQo4nGQcBTCJkI82Jjoepd
7GCh3QXgUZACTO3ve6JYv8ZO1w2XUS5Z9+aVBXjT8VdpcaTriIiUAqNlAPPSMygW
0Umdf/mpU6ftbTcU1CQHu+f5Bn3dVzdJOggOWpPSC2H3RLNX91rcrSkF7a96YJXV
a8MyFMxLZvLNQr88DQnr3oStZGDSxJ08NB9AeGjxUKN8tY1chzwla2O2DFGd5WhA
ekpiml7PUZ9ydIT0K4sHQuwsBxxtdI/rFQ3hxLWNYfc36h9HtDVvPuE0Al9E7g42
O9FVPElWAwkMgQpDZK0G/ToRnGsgTQ/GMmn7QHlnCVb0xKRmxb+I43qzBJ23Vfsc
Si1lrP3DwS8mg181ypNUbHBcN4bf+7nHt6Tp4thqVvUMwNyEsIOGK2WcJK5OmJhc
Wfa9BowELIPFYUPsBBuxLGMPDDafw5x4teKM93zsNgkUnMn1zLmg672bw1CeNqEj
WRdQQGsZG6MatLc7ut1bezvlxT7ik/jGhwApcXnsqNM2IbQBiAsqqkRMtC3mNL9j
Y5qbIURfB+elNuBuF0fj5u52O+Fx5ggu4NNOjbSwOY7H+mjWrdl3M89kofTMapnn
cbLr4gGKVJXtIBOLtGQ3/IH36+Q5LzwWwW/cOBSkjTD1FtB/Z/TYXAJqzmR1Y3UR
3wre6M0/YuiVxi+qyo4pX3+VSa5JQ5UoKPujqjHXG4qFuWh79Y1k5mG0D5bTOFGu
cUBWRQyEdmVb6weU792aDKYSeASv7qYMwUcG/EEV0OyOjPzraYHO3bTbK8845Pxl
ZzlFkeWxVLJBDQO+kNV63hEBfHn01W6v/lgIoC8GZLPIsHWZTDfWuQSKBR1EzBkA
+CVKCoOdA+S5KIkFYBfJ+/Dhf19bSsZ0mJAoFAqd8m6BTYSmN4zUciOzTJ1JIy5s
KdJUPayCS5wSixiOXS/magDVPdF226lKXtbSEw92pH+w1nMNeneLKLFvnA0qzxxU
Rr5JkaXC1RfEd9vNQ5fVrp/YMphWXnvTuKu6EIBBb8Hywp+i1JbX/njFP5USJ/5z
s5h9OXovFDbB4q5+ODm5iqZCjGhR7ep0OXyokA/Z8Bv0LuWUlkXUyP79Nz0Dy+Kq
a6Azeyos4VPqcfWzlofshMOcTIeV+coBVwoR+yQFpfxJsaqDp9FYXY1iDwfYrnfh
E22lrfUtCGOu52UKu1WOPjhlFlLI0mPO2F5RbJ7AV7PVLBbhoZBPtMlQisKN/vnY
j72H5L4P3agIyC3nKcLzazeJRMWunj9p+vSUZKknpp0DlnyEZbU7cHb7pSuK5S7n
cJZDx4G45zNoud3y7E5Rk0txVsTsLSHhJBN4+spfBFPDt0K+zSsbqq2ZHRanIusm
2kw5m9gyd1E3a1mYoHNT14vxmOlaSbrp10f3SoN3jsAyId1KHhvDFYfSctQyNvTO
IOBn6AXhy7lONXDWArnIWpxX5T4s2kk4QY2IPtqbb8O/I9HsZ+XbnS+zFMEDa/5L
+Oe8CX3cuEDzbp8wshbkPRdT8d5Xj6Hoc2Bml1/3T7f0C30H9Q8xR6DBi5W+pSGS
sDTe0G+28HwdCYlbsQpsgjBO1ipqVJFfwNvobIcBIHCqBMP2FqXHv81tCUAo312t
mrayDaXteOfI455e8tmY76n5SRpkcEryksN4G8aJD2oi4MAyaGZEPTizcZPFlMHQ
Kagrzxey+NnsO0IDdFKdCuiRXxtilDyDIqSstlmRr1UucaBmzzTUtXvhLMhpHjcm
/WHBX6LHUnBNDBDlt6/+8c0s+dPq04B5Z0AG2pRNnvcEIUDPtoSl65F9M/Fam3ue
mBEwaV94XeJIRFhPYwjQ52ky1dTqJ7LcZgAveaeQ1lyryLkupYAYnIXv4H80qki1
3RScf9FHWZ9OerCC/qGbQf4DotYoMYf8ErOCAnVmfoPh1mPBk4J0AEaA2k/IjNeF
rxri29eVZ2U6G1UyI/M1PkOkYsoBXrl3pdWVf8Q3qRiuHSTGtZINtrvHgT4tgnaB
G75oPhqaHgi81zlonq1xfMygUzdesHjT8YpJ2jI86f1XvY+Kyhpg+UDXdor8PSHK
oTkK79+DGGvKwjG59h9xbr0naXR0VoJ3VJfkBXs/fA1Ve2S6TeT3BlV0hZNT5Oeu
Uh4wHs51W5ZIQ/7pd9rrw7D0aBBc01asZLPgFRlToKewDIYLQear1UaX3ZHkZNVg
0mC3RDBHOeA6inN6c7pjRhezkQE/Z7PTnzXcLOD5v0kJwKdB96d3q4eT5sM6NVHn
SaJFtIz3h/nJq7P+YsM9JpnC/rsjWDTrEcoLu0tSMuSARrlRZU1MoQS5Q7OK6k14
HiYUhjbmwWx0TpGz7b3in7q5oXdNwtU+lQx37Z0L75/Gxt6sq1UU5qen/3dUT3F9
p6bxgvZk4EwHY8OUJi9DvhtMn6fS92qt1gzSVF7uFQVibdROT07j0DjCXu+2Xfck
bDP/cOhvUCKnxv1K4kN7XWS7yoJWcGFkheaJBwYgUBmYRX+81oPAZLlFHKhc7KvE
qkKEx/lmx2Tpi3pzp7i/jJj29YBEcrHb7bg2/LV0Bfeu//UCP4zz9+mMgFyQTrmM
i5zgMS2GMZ7iV64hXY4k0RT23CcaTdNMpVClkm87iS/TEM6PzkOLJB15/oYv2BPJ
LV8mKl56tlHPVteE35emREt0xU7maJgM5FyI1DdddR12LTsu4pvaFiq05Q3yYiyJ
3G4Nl61sDNjKhTitIz41qgV8eU62qZFa7gtq3UjN1WRJWh39JYLl+IzblD6Op1Nn
FMEHWQ1w8/seUY8CN0aL4CsZloAgrkkWgDuCZV4BCxhuq0cYXOgFHpu10yioC+qp
MhRoU+Rl7rC6SpYlg5fybgNQxLO0yxO/R9ioNDlrQEYvl9F75MK0uK+qOS3rCrzz
JknGfTgd6c/BKi1P+88FkTZGD2Efs9uEAzEBjj/Y20n0Wt5vVvy8w2hvaL6PYwI2
FDyrdSdCheBMruYrAYd4kOAKcywlfylGdnfOXDAHGkKgEe5mJsH94XXYy0Kk702f
XZMCEMJPzYsXRjxa1JeH+hbTJBHAGL3j1dH7dKgXr7dy0tGXUd7Rj9eSz0BmvJ2w
nQSvX+YBzRbeSXlI1RTj14uMIuwbvaWqKRj5Tlvg6htkkEOXb9OljJwUv/T7nCE2
K4mepu8RDpFA87wOz9MrUb5QrJ74wPXznRon/YYP3ciKtwwzPHnK4rekuLi3KkYz
yHD3/KZQYtUNs3RGAuqDZSpG4TPJkwEJspnlNB27aQsLHcmt0P90/yCRCjF43Q50
QHFfxeZ88646dT/C+SzUYxVVt95lzSkp/i80f3HPf1T1BDbtuu5wFBfXreHsUgfr
17Ro01mqVqGF02NAq/Vge6AcXu+wy+/HDKCtoKed0DDuG7NTBbwxWDbBxaw6usoW
gzRX57lpnMBP2BkYmKyWISY6y7jA5mXcXnmNYMZcxbeFlEYrJN/JUTIcwY3+/nLh
WxG0kbN+PWpx/F0WDI5VvG/WUAZzPcRAkc1swRFEfh6ap0NPGxUfv2HZrjTLcgAn
lH8gO0gRaOx256AHH/LSGkdOyWlB7oQh+Mb1m+SdcU9LflmKHzY9B1KqyZOtLNE6
2C15BvYCXsmRh79JSiTXN6e9UT26nryw6x5aST4P1i321TZtHT6SLtE8nKfJ9haZ
3PkdUotWWK145ZjVnxMF4U9H059hUPxg65JdQnflSWQvVCDXE62ITXIQiUcu4m03
tPc5nILBaeLZwbEKSzl6ojs70ZLD7+UFvB6Yap2gBaDL1Ty9P24yHnPuzuuhDE+d
O/LONTpLjwq8s9yuaB1+xUr6c4bK+xkF9jBBM+9KHyQzQZCKyffhUkqrBBhB2bt4
tALBYb06WIDQ9ZmGRg7d8hoxZE87IGtErEVpvEbN07MTEAg/SUUZcUiC8erDoYTz
9PPc/rRUwJ/4/pwlhe+E1rMP9GWLS6XYG0RWxhaZU+lEvGV2GRDn34SwTh7Lxn8Y
TFRl6apDoR1MZJIiMtsjn+iJf+W9nHyzxfm9ydq+oouHvVwovGRxT9Md9Fcw+ehR
Z8oCKdK24QVvS0OLEJlENMqTKpcKV4kVJfKgIVz4BllJGhaAzzNkLRl7sELq7MpH
pBhg9R7demeNwirF6rLe5aWS8OL27AT6Tt/m0re1krFWEzGGParP4X5e4TUuGeff
nyhmd6gjxxnCyh6h1Rn6oKf/rK8jpUVrzBXJ3CamPdgKUDrRNGbBkwfbGEzp8fqZ
Luo0e8WQ4BJ1/Z9aMavD2V2BwcP0ZfywmnznMRVvMX25frCZQ5R2zkIzasvBxrqF
zVvCU9eGMQEDnzvIBTDYmnfIvfEWBZlfHnNDwF1k2pkFC6zSvVN8h0Y4YUciFGba
EgIhfr8+KScIMEmZx5fyWH277a0/xhMr3Cofb9ImrFjSzC/mcYjj8y/oNLnuAPVf
JaQco89yHKnvqIB7vtxfoYawohXDsuxVTex1tUNyRx/dhJJT62OD/PDWJYU1bLBU
nHx64tpOaaNidhW619Ol/r+E1Lwx7NIwcNx3ifYnCHW6135VtEbJszGSlT4ho3HK
22PsLWll22zAUhpP4D4VpQxczyzrLWtOT5h46DJUeETcJEk8vzG1FvtovxS8oNQC
A5QwYBKtb+531EMKjEbZAkg5du6CmIZUoztDXdjPX0gdSq5V5V0Uay9kvisaYBqo
GCt503BoBcyiu6Sum4Oax6+mkXIPBMpjmZTmhNwtfs5IhR6VxbWyH14HNOiBrY+c
LVdBhj9swi1gorO1GVdj2TqCCIL/HCFL52Sn+by+L4B7s3Ew0qhldV+NKfXAkv+s
cXpMKbC6jzgygPzdEYHBqn23Z0FxOzUX4WiydouA1Dkl6Zg9LaClFJe9RoyPjcme
cR3u7EN5+NGfHZPh5BsG/o9FMMG1obJqvr7iYbwY41kewGV/NqazjZnWw1FtnVoX
M2CuPpjCzxbXi5wGEw/irSCO5lqw6kx8/A+n7vzKqHNS64uNjOj/3RzJuTmTTmRg
VhJB6Y9W0iKQ2uhnFeZK+i38691Ae1aijhVNVo0Xo/LsO74ndovGbFkVFRcxBII9
5z6h5MTEeokW4fMLiSJElNy2y795zDkBWWlAEgBLVcwGGln3weNwNCgBpLcylHXj
Xs1gfNji3FvTvDeKgG8L29KmYGXcqmltfsghHNyeB4oPw7OQbzVeFlrJBCNyL/18
sqHzpLRFq1HL16DYUaEhynNNGL1+4QSsY/sUfZkKvXdXSaPwg39D2JUV8tKqJ8Jb
ahCCxaxcMbIvYgrQz3Okn0LEy6Fndf+1ks4kTbZDq+ttZZl+FuE3JrmSp4F+P8i6
DnfpqCqBYotnWeu7UmZSJ4EtOnbi+Pj+t+AdaqXD7Okkyg6xgCrv2AFc5P3CX5AV
3fmikJyjOlFGPz36bWEbYsLmWI8/ML/bDeTm+i6vYskfbfZP9+ua300igkS8EFl4
wJpo6gNvmVExczjZTGx0au6E73MRhsZ2atmO25m6WU//t8XcQ6TpuLxWRdTBdJLt
VX1B9JH8ldsf3bnQL0Khn4ssVn09Jp3boqiGau8nXnsS4Sb2oTbucKmSbzaiAwEZ
JErrOKWVi9FQjjjD7zyGUNiZuFcnId7ZxRTxhbndVZO4hDeJFBbbNvz9CskLNoTU
nOOIqv7MLLn9tMddf+9HN/juFqCR/VfkTQM6b1pqBglWBtg3qqE+SZz/9/HRd/e9
UbmOWaySjdCbD4pQM3DBkAlC13TN2OWw1IL6sxhMHj6VfrulagsQEyTsx31yDIFE
uEHfIl5ij3V3BYFuuDD+iDp4NKLdTK0SNUJHYLz0514bU+qoErb+LvXZ8lyxTQhV
1tSkDaVFbgo/9XvXVUkUGXfwnHQ+F31Cgx/eHlOeTd5zAICbOsEcEtLderQO1vgp
CoCkZU8WSeG7ib3SW223KxR085O7QADC3S1HOXIVQrLhWRvHrgNdqt4gRH6W5A00
C2A+Mo6+DYaqIJQMv2cQSlY/oRDMQm/1eBiCuX2gIrrbGEjbAAQdACRPRBoSghxR
G/2twk5dPsYKwdq8TRJG9PU5HFIfSI0tmujm49Zxt8Xnyhm7KU7rFXOoWtwDlQeU
kvvv4OQNnUuRe4iosKsYao5fPds5WElJ/LeBzj+yCYYoQ/rXjFbYjWHzjdHWKzPT
YvPM8M8OG2M/nvW0YqX7SPr9dmKgagjAe22YCz1OsT14WqU7FP3dGyZhR8t+s2Tj
04dOAeUXftnccTurmVsx3SzDOlLPUkCZSFcb63dWioeD9JtiaKynta8nfSeHkrQO
HHwU/eY2ChoX8l+EcTXwL+IuPBDeszcEtEYtrloDaAbeZq8ukduQslsHQDxAfgPB
w0pVlnXKGJRHw/Itcv41qSVP/aUseAuRRib4TBB+nopMEi5MMcLVA529mZX56jeI
bwOp0YhIbYI42gEVOx6a6Rj4ukd4s0xD+p50/24YahyAu3pKN5s97CTbzx2VyvZk
Fnf4k3qH2dApTVSUoKccVNFvvcyKR65c6qjfPMxjJEcpozGpIkcMphfZlEAL/ZUe
Nc7MvbvxqmDoqat2sN8CKmv+1mukii2j30vJH7kJCuUyga30jKdn3IkDM5OGUwkt
HiCsq2NvOKotAHz+nYXEyzZeEC+F9IU+Y067Duy1qZoyO8I4O9rssCcxa4wfUx/X
pPCXoLFC1S+4d02qkYo8F6MSNWCDEDRY6JT80U+udrKUF8tsn8nWfvoBZ5CrCu6o
jEsAclhHaP4/AH6VxYJ9D8giQI+Vfk8dvl4qhaUSu2nDoniyB0wOs93aDRJPdPsH
3Qvyu/t5SsxD5K7KeBtK7MJ1TqfJW2sj4FEm8l7dILhrfloSt8xbZsmieg35Pm2s
q78mwvrMWyJcdd9wE5UWeIRgyzebRnNaBqs1iCRlhqRXQiULgEMzV4f2d3meDkvQ
Qm7e6SkU002v5tWc9iaBeAANd/2cuk9FSoh5FxWEvBJ4DDxskD+7fqmgAaE9xwUd
d6F35AxvWq+8vSi1uJoztN1/DJlezxev0mItB8O9o0h7xHacy9c7O+CjAR/HMzjU
IR6aGrv1TXkKOU+0TOyT2Lin0fHgIa3/OKX/BsXmbnj6JruPIOKNVEAkSctJNLKk
+ZFylSdSc6xtd2rPsC+xYxaa0REkcfqHkG5MmW6YV7bFx4E6YFGuNw6W7n+M+6fJ
xhzYQLHhGjpq+a6xlJNEQjcM/1GlWgJiMVO/qMjn5aXJGooDi6cHf0nnnMD2r02M
DPIu39Vou4QYrgAYJyRXLykyYNoKvruyJBXY52VcG8YVd5W3mgsiu+pmgU44SpSA
f5uYqp6BLtHZ1spG9DeSLQnaulk5fN91zamfTLetmHjQJt3lkdLhRVNW5UTCwCB4
RlQ4xEKtEMIztFpnI+r0eKG/MeGPppCwj2AHukZ7m1bioEmD4TIzSYgEDa8d1wkn
Th0wLBgPvvPERI1HEb8sZ6wuLva1Vogevi/VPw7tPg973IJAFO3oB7SR7WP+kUDE
JbTZ3CNrfgVUKd9vkuTM89aLckYnkUUX4eBnADLUNAfnDDG5shhOf3fDW6wqDPW8
/eoRQfpcKGSz5lvoY+Mr/+mteRW3vHiY/aHhDXacGMDtXttlGNi1dfC2xg78yB62
pIVYtGhVhuRx9OG/RWIp7wzaljvB36LodBZKiFh2lH4k53hTzhamu3kWfiNNPmK0
HlSklmZXlP3+auJvWUukx71p5aRxbXLeBFulkcp9l4SC5tIWGOuS/uM7ZczbGXR/
BLrZVMIZYeBAyZyryGAaM+Ws6xNTTfpfrCBFjPIjNqNUeO/nhssTKdcQ9auM67K9
7vgDkiXVR1ttXnGSZyEaOErBMiEGQiCb6tTJE/T/quqxtx7Z3/xoZj7ato+MSfC5
YZVI9BeHJTLBzWiMEsfKBM1P2I5l2NZKjWYzk2R1TLv4CkGsK8B0f/d9Tkib4vw9
ljYNfr1LOaX73qoYJHkN1a2NnaZ0/dCO2cwTvvGvpvnAAPyVUR/bC7Cfmx/oO1VI
xu60E3uN7d296VoJJgU6Jlrzud+41frNl3CRwK5Layo2F9xdc2R350Q3hVg26RbE
ZplNgLN/ViVkmhY2wNl9cLqUDsQSypUPzZ6cM5sMvhV3P4kg7NHoUs9rYE7Xcr9o
MrFiLrIWkOnUiTYLY2b5K0mtKeCz9fOaOE1qf4C/nQA93CKCEWxTPrxWTVJ6Y+NH
nznKQd05apTulStT77B6DbS75OwwWCN5itLy1vLXmPBdLSpazA3SHYzwh/lR4uZB
jyOStOVcAr3y2z/drijj2VbuoGSzAm6+Rf15i6zyhZCRoFljWClyoyD01xc6lRmb
Xf50YdAZCfpAaUKcf4FefzsLhu/5CZVO20FW82UbJPVYolX+Psv7jTmS40vZraoQ
UW3XoPeqWhZuYYvFcKOsB7lptaG+5m4ExiY5ifyXVPBj1eCoyMCkUDhMKwsY2RPp
eQEejixFJAJjZMlSXJ8zIy3zlxPdcKN4B8GnGzxByEvKQfE/AjreAo3XLuqOWMZv
hfvdzyPTwRLIGVQnqiuRlpso8QU6nAonWd+xHUMxlugTfb6m4Ufa/4ILfMLWrGjn
7RXIJB3wF+2SwgYWb92F+YcG2t+8vHN+AW5x7pUVBWqa54I+i9a0xQT5nwMysL2m
dKdOkdaT+8jRnr7qN6V8vtdm1kAw6+aDruuD4hX0auqfEzik6TbID7tIf7Kr+/2w
o/EmVGMM8YnTHGF63/FGK4n7X5KAFc9RpAWy76DDEpSiu5+MkSM0FS+LxXioRoSI
L19SBTCqaw8I4Yp3lesFSx169zC4P8zZlEV6Chjkjb377P5OJ+6KzFK43CSah/2E
GIvUrxy6OQ/EJUA392HSxvpVJv/WnkeV2+wvh+iAL82tBbVzCxTZFl6HOKCNll3D
g3q0wFsVxtGBO/hte4woMpivEpRZlPTOj9wXu+RRyyCIU5cv+d/Hzg6q58KYglDI
e6SEPS13+DYgVd4+gNi0pkxTAX5sU9t0DZbC8gWVhTOwgGKUo2bMn27P9OP6Mz5l
A8/w2zo8SH/pgvyDNtAqAdOqmnPAcWkvukwsuBzYAc0MMzKQPRhd4Pzjf0SmG0fk
Epc5rwkXIDuQRoiFOdJnTl4EgVX9EKbxDRMvMZgFsBTpaVhVbP51G38MsskDHIhm
6d+KXm99vrtwJ56g9yFQnr5yCQUToE9K6oV5SzD3OixkS4ZBaZWxCCFdRBkTGw4+
uJc/+voihBHk6NaUIDbZ7iiaa7NpzqCmQVD4DEasaFowxs0SIxxxCvgDcrZ7+jSI
ZRVZX4AYDWTH8GtXXCkl6lwbup7KU5J4ls/K44Fq0efeSXoqEnvmUWKOT5VWe48c
SHzlrigwWQ1ZjLBYhoGYlgHYjHYKOi7kWNEl7sy6u31ErsJAMskTCNV8d9o4ipB8
5yKG7TJmz+v/4wKlR1cxei8UtnsMEy4D7pPBeXc3hZFuQDAOdE1V66tttTEvFHhD
kLCn8B8YrgCU/GIy0F7ibXlp2ko+qylkZqsBqkHCtXC/Tkoc7ogLbfWk+vU50yfq
Qs+/DFstfvrqy0cnzDzAsqDR9szYc0uXXXJKa07hcewODLV1vYJxOm7sNUVb9fHm
4pHOJN042j/KO7D+07er3nMxgVho4n3D5VP7qv84A2rcCwA1o5vLN3ATwmQwX2Nu
rpb4SWlCUafMyn6h0MJHjwAM3j83qglh3UO+o6+DeyWeO8ZrYWK3yiX02xspAZU2
B6R0fhClEBsweDoEvmO6UuY41WrNZHoVSLhsH4Oya3bgQfxSr0J02rHMgAkIWKPR
V3qkeug4R+Y53b6m6LkgeVuGMjXlU+oSmgfwEY/v5d7XMD0BBw944Lfx6ru5KGb1
digWsFu4be7cizK39g4olIkn2+yttQ2sAhmnjz29DEi6pPh35Utw1BtPKkANKXsU
2BLal9rypgqRJwBajzvUuXhIa8cnB/xbr4J7zBG03f1M93/2GUZPKFQAKH6TWnYy
jUqbxas7BBg3x2yt9lxqt9z7SLs5+7EXpx4jEHWIrrHb5z0zgc882eVfigkzvScj
/ZYOhHBLLyfqpJnJaYRETC2RRx7wpxSrvXCPQM+V+wRKNewkjwKx/7wS6mimgxF9
9R5ytbBZhhQJ0amiQgFglFtO+bD9FSgiEFv4Rfesls7AfBdE+ny3Z9lRMvSui13H
Md1itHRxgBHkNUWstej0FZJz6DMzGpQP4fdUDOADTB6QoPpCMsRvfSgtB6wWxU/7
tnr7GFfE5plyN6mCQTOO6g0M3hRD4yvIH2D10oce+UABl5BFwFKJWr0vFDnUdFA/
Cjwa0tP1kcGGD0oz8H2PkdH/WyS/pvKMW00OIGNZLPexFos/R2H5xR0FuM3R7aXc
xHfm1z16NewKr0ULHMG0t0dYr7/bZ2eFkYP6BK9KNcKBG2KYKVUyyompeJNt8Bc3
Iy/KnuwQKV7mhk0TuHSfd4pa2otdEoMh6vIayeD5u7CiygDjRoaNLh87iSh+ICqO
4T19UrV1mNZm4PtQT56A40TOgGz35HSzjT3xLbueDFajoNVMvWfutOnRZumEFpCY
7VbaFv+XDJ3VK9Dpb2c8tnuo9LXFcUTe3ForjDzfzmP6Nfs7NiSj0SlN9IG7i96G
iz/8o0tbjWG5+jijuH2QHW+LNjWFxvH2dKjFmo4jJD5qiLyKLfXxSidlgL4Nv344
9hZI0Qov52zhtOsJaT/lCwlFJE697BPO0IEoYTmuQfbmiTLw43f9El9ZM+cYcFqT
1kTox4ORyYgY13ewF0MLS8T8SWazaoHJiGrbJyMwSz42zpb1116xiy2U5dOrvLXN
Ok/HcbxbneN1/YtjUITjvuYhpl06T9hQU3oS50Dkp9UCJplR2mYtc/i8fFBF4P8A
GSqm3GRuokrB+zqSwy1nYRFNOSl79l/8oVRDH3LRnb5nyqvzVPWHqqycx8PqvRwv
ygSgOFlbbkjc+4rVMG/L/gNNLJZIGP9b0DoBs8CHDSSmvn3D3+jkQ9F1fnMga1RG
oPP2I6clT2jWQcq5OK8BJEWf5/AtOXq7S9nfjONQTnF6dmrvma6MZTH8iNv/XyLh
IA62OxtbydpwGhQ7fJizRDKQidYJCWcZ68dkmDKVZMP958DXQHH/VTNkYvndHVZn
N0QS+xgMNJ8YkPWER0aFoN0tkCj0LZvutqcV2YfZuqyisqUd8bJ7ONbhW2upqqvn
MAFwB9QPs83JkZqUoOAacJDa2k9IkTLtn6UIwOJT4DUxEeIw7GLyNSldSgf+Agwy
KAt3LZcKv7+CPHzJ6rUPhK8y+qlHZsTNf6ifs1cC6cvk08eC+Bx94NLeCoXGunNa
m/cAenpuUGU2ng/IFelHbUbjepvWRk2BXnGjkmsV7lBji37+0YQ4PfIORuUN37RJ
pKUODsVNXHsu89OVEfktFmx8H69UFdbkwiUWxvjupfA4RyWSNES2guzTbWEdE+2k
ULPPXDWx7djDbvwHn+GxnWz0YFwU93DL/awFOTnTXaDSGQqbiXUyPh/2FyL6vvKP
G/yymxGM9mn8xhv0tnZ7BMcXQZGQR0CXWebHGqFrAohYYTHbwlr1eYpT+VpEhvzu
QZhkU9E0BO9KqZ/AnT3NglGGjA3cnKintTfeoNFqR9ZyvOTNNMlGUULaisNlpcq8
MlqosXYXFn+YBpFniPSJQRRPund/5HK30CQhpKG69oSk/4lKBFHkRDkkTTntGsFL
8Nqu21INlo3iS/tb/d42/0rp3hQNNH7dYtv+v4sOZeFelkU20Tg/iR9FOKYZcMyt
ungE46EjAbSPEAw9vMn0rs+ZKsLNGMRdx2bJPUtcJ0pyj5alUfiUb1XbaXg2OKAc
1SY8QztSt6HtvCKVCnxbgg/ncYAel8KUbE7YOE43+Q/QPzMgW9jwLc1ktzSKUA4f
MFAqdE3kf/lgurNQ+XwBcy3P7BhH4pnxKwqqKqXyhTJxG3WNRRIcuRS6CBH2ElL4
9MdQjbcS+X0Sf0Ruxk6IPgxnbRG1PQbuX56+drjZvUBFzX15ok1QjtP245u78lUJ
dlWJp+d9EfC9X/vpYUrLghZaQLLfJzf3EucJZK1uKjUfs+EZ/0/HO65EHFgX4hnR
OgzNvT8bOOMvnbQVVpzq1zlNMTWvp+c+UjawlQchk0KLaytnTfh7LKdj0v3yLYw1
szqzSC2Ioy67q1lTMxIBJpVpnYRqggoH/wkPX7LJixeViwKb+OARm4JrXC1nzMOy
LtkkcMMj9vN7lUfFmyALU+hh+YBaq01N3ef6ltE7FY8plsLATkY0qRm2m8M4daE3
uYZz/u2nB0effTflB3XxNdNyzet8ej4EUmZQ6yztmG5593GFLQRKx5hHk501oVEA
OeeVMZ5KwOFD+devxsBYumuFBgYV51hqxijAjpRXrbK29FTd/PFO3uyzQSaFJk6y
AN/gNO7VJ7XPVVC5BNYNbnd40Psj7TTYJa46JNAZREFn7scfYe38oNXtbMuhPDNu
kvRWVqvNJ5o/LMKf+yd94veO/j6NSHI0q1b2BioXF0dqTp2yacQDkQ5Ldi+crcTa
6PRj7pVHcgDM1BO7wxOGwpgInZXtBIsRqp6xOVkGj2YvDa7Xfxg3uiAVdxAY+ZrG
1Px75gbr9eEwO4VxFIAbicOX1iFLKqteoF2K804j75Ua9JAFbch000gDfO5NQ0Q7
c7NHEF9tVHfv79Bhrzfe2rCovv5X4YKI84NCggaT+9S0+qc2JDl75+kIyk9VYzQf
/nsfOvyswef15ikOFQcwsGXKnA+kN7q63ZVIOylUvkY4y+5cBokVKnNFoLnEj0eE
H4aV8ae8Q1XtpNj4r4g8bj9WNFajoLTpItAbWFoq0+cdpizs33qhupiwHx6SMtdu
IG+3jqcwwP/TFYRoEyOCjYFBoUvtCcKy1dsUcg5VTVETVyBNGOp04ca6IBn3O4oV
/8rgvsl+tNYRAZ1eN1snRr0tuf/p1ZcB3PKWcgZo/vR++vQdaPZ86Az0ijjQPRcT
w/z5oE8xVmr9F5+LmhP74bdq/FU3G0dlnFLRiVUI4AT25C3sCYMhTJo4nuDLY4eQ
MkBUOp9NvvRP8/scUHiGhFqRtLrRugHDhPCh2aniWCGTfZGTs3wM0P2BjgWIpN4w
oYi+uXNjBtDpurWOQ7mw1+1aJsQnXayVZ/TyWRaNKLZfTnXc6obNDlk+2T4/hqOs
od5Rtf068rGKD4+h1qOOouzwZdIK9JdWi/dFqh19VJSxTElcOoxx/NTJjuMucJ6i
QZ6w6E0i2zqAk40J355h068HPRuV5TfWILOVZDZ3QuoItd6L4OgbUTZq1ctN5gS+
TlDCTZyAPd/A39EOL880kydlJKMhUIRKPNmbsusuT1Ucx0s0EJX8GymxEj5br4Qq
/G4W3VJgiEJ3lO8J/5ZqSvNKINMq9QqYRAIs/rMl5OjxM0p4iMQlTXl78vh56VWW
G8ryfSqb53g8tl9l/PKFfXXvpDD+GqUOSRuFJFVHigMsyPkVM/ad2/u8Q+yWIvIz
2YJnMmAxp3l1W6NKpP+GdoyWjDtecF+HYQfwMS12DyM5Bp8Opi8YQa25OsS4sU2b
BLiaeIw6G3sbW55qQ0HrmkSAXNs2p5q/V8eyAhYm/9J8Nshqa5XKfegUK2JA1T6C
mURMSjBa2yOOHAo484qlve3kXrsMwZ744KUaTWmHyfX4nenSDJ3Kt5vcOWlWvaZL
ZVuGXhIQiMh2kJj+OwTGQUc9iTmPVq3Oo+0FANNLK5fIh1fOZ+mYt0lIrAf6XZZ8
Wz3/AwowetStE88rH6JHx9DZ7fYEERzFBNIDwfJ9PGDWUf+G+oGDgCKf4hb0AJz1
nUlnmNDcOTBLa46ffV4+u/BGZ/WxbuEQibaQeAspUXaW8+zWfAD/qThyb8NSQL53
hrsoDSP2svNOROPjFiH8tQXZaZSq+7fCnnZx3oROOzaSNG94XQ+AeCU9gPABrtUY
BPkLn9zceAjDJSNmWZ7hdGIAf+mYG4t/18Ixmh3SjAzmGNkYesqBpKdH6YD6sJNq
hma0l0xyc7giKDA5XziJ+cDSVZQR/4fIx/8dU+2aZ0OANfFCyG3FAnYBKm0t1SwM
x8Ses4R77GKKEu6isYGmy7hvhtdmHGEt4emoEs5p8WQOBxDmliYJ8lo6ASKmXJ7U
sfW3iCLxPZtUcKTZy8PpQKJFkHYEBsBMB8FrWmfR2o8EdozE7Z74jkDjllqt6I9z
GdywFZu1uBm0ltBrl4Z5ROLnjo9BrrG7DsJOOCfXEO+bdxZB5KBRkKzqiJE2fzZQ
opOWS2csLDnvtlqevsCz7s0+3DOarIJlBCETUVl5bkDeTkxNA7wbRf6QxY0sC/Yd
Ewvl2/FCBh/Pa4iBVWqF3DkZEW0NOKzEdY4SN/FuHYaC+DwQKSOiLpmCuNmowGBN
oXzF+rkWKFnvzGJvSxVRdvbXyGVS/Gesf9s0e/QrUaySE6qzcfGAKMKMpfdQ8WR6
mqIgNPv3JXSHfiTDkJEvITfIiVgqQbsKjAKW0RmnWSDZbs3il2DI2U8FLufkvZMj
IfM/NJQX2buSXxjOiWtAtbPBLlf9qEvc/W2M7Y1sd5cHwiX3iHrXiWswf1OIEJ+8
mENmM8jgXY26UsSmyUVjZ4eNjRoNHYEXvLRLzrEtapkpe/I+UGdSlO0OST3myrS6
mbpePLIjJ84psJKeG5MIAu/7p8wxWtLCGgadbsUoqmlW86cuiFw4Yoef1/V+u+qH
lqhj+KSa9F2BlqtKfgYGwptpDuLNE9218hXrVyJTKdbCG2+c32BbNThVwv7cdxxy
d3sIFAlhMCj/n/Ydv/BhPHk/Sllgxm+sL1uUtWFjtNCN0MFV1wJbsul8sXMgTDoM
0vsySI2Q6BHGq8MHDTDY9FlcLuXscsfjleqs3lT+a5nywO1zY+b+dyFp87J2tSIO
svWcpliJn95cfInbhAadE9uOHisZguluvR8fqTkIB0KE183m7NAPyo32mda+k6L8
SnZuyrW2v9/UIhyG0zczwUp6qoKmty3u9SLwr6NLgtJdHU5hfnjLrTJcfuybYRvx
ic18MWeMQJnCBR39wNMAQd83cZEySVhjbtTd2fJRzncdhTdRozSiQ2EXJXKkAXyc
3YgS2BvSqfVXEhk1G2kJI0W5UzzwEUpWNk11sDu2rDTiALJzQUVdDoMl5STj98d5
jJ47lZsxldkh2BhetN9zPrfurCUJNQrPV1RCkWITPPCO1LqvmtAhnYasx1qlhHea
KQX15kRZdw2tXAkQiCZpsNfUmfP1GTOUPlDM8xDRow+1z5nHLFdUEt8fndEWNVRl
e9pz2ArzTEeCkIW35Yi3f5aAgd1CajFad7gfmPmaPGBe/Tv7s8fwpnjXnCzgdpGr
HBgkBR3qj5rv3vefwM46HiVnjv0mmLpeVs4B79JNlLU8VQQ1nq2HYEwSakrsGJB9
Kg63Vp5lrj/+KzB0Q79PHJFTwAbTEX0WK6yzg/CISs1wxLWaJJfsBIWpZrugFi61
oBoS7iDwjhP/27zfcU3X77Fif+R7FnOhwU87DAYizrBuc8AshAsVEDdq6OS+pffG
4Lc6MLvkMzZDj3oy2Byj79FXjWxHhzWED3HPpTZbrimnHaXZ4w/FwH0UNZWvfL4H
6y4WFXA6y/AJ34zrnxtvps5mqXVP8vhXCZV69pnlf6lZsZ+ZQ/iPLrJdPMOEEsTr
MD/ojEcF6QT/ASyleUFvHVFhfWZhF95Xw05SHB4PMOde3NTUhiFTy7O8I4FL+dXW
YZf7EHwJAr5rgcjMeB0ALL5zwunwAjvt+IsDUw8vO9t2vcNlb9ToPxd3zeth9TqN
ZkJTkQG1T6RVY4ShqFIsXhs8hyX5vqL4DT8lrUa7P+ION9aPH8IYndM5CfVW80NS
4bldhy+33RXtQwGFWfR5UiIeXVvFOL14Ppa/D7BSvQHGHatmPTs5iAOEDEVAiRBb
yY8E2IyrQXeZs2M1WfoLA6z2Lk8Qi945TaMOcJDrLaEnC62CdIy+/3kwHTFDi9Db
0nbLIW0OGwofV6TeeREvBMq0P26bqFFRoOGqijukSsOXR3crgNLrV/yNf4kjEZO8
F22gNvXza/v1e2m4AA53S39oGpDch0BVHrcH5slWzn9bP5/f7PQXEZSmJD/LKCrm
0qmJ30nDIxB38i1wcuCZf6hGC1SKq9YsdJjN6/QKyfXQ8IkZBipk3AwqVtipdIjY
Sqost3UTsStN6iTep3/zoMMpYNpn0fKk4TumuqD0h7ECtD9+9UXGM+f+8bVQmL83
knZ0DRjqboUHIGdJJdYW49NLAan3Zb1/BnNtcFOsVf9AzRiNFNtLUPySnu5iMNo3
Cg1fMagjkj6jcH764TLLVkXkP/LBk1g3Y9DXDMts1S27y/Xoumw/0tf3l7zhSWzc
zEK17SCDF+W3deH/IbGXno0W27UIPbjaB2WKRYkEd+B+bxgYwSqHxzDSzcjcB0uZ
2C6ujs1t2efJu6mT6uodrYfCgOIQJPCOR6tb7pHpUm5QkmXByHDNckOO4x8M1/ix
GHwvxDb1l7cmZ0j5htZdbdbQggfn/T9cDBkIbJgTv/0obU1cmkWt/ehDtEvxLsHU
sSft+sSmq6zywE+1Bgw8s6k4kqwLUWJofou8vL/srazgENY9ddjHqYbgRSjK5eme
7WPwolDzbYlXe1qSmRV+TZ/GXijoGqCOoh4W1pl4rfc9EwnK66H8iv25mrpZL72D
VagmA2kVj/s5x/ars6cIfe+47r0er5io7VjOKst55BujihQBwoUJq+XU3HAdlM08
0dLrUdSg9dkkLsRrsyjDDwJgZowginZGqNfBo4Eoo3c9yNraLEylJVTIfozB65hj
VuNpuqTCmyhG/hjKPvwvMtoLorKXRXIG76dmcfj1z3YtNRqz5vG8Gdoucfby9ElS
SQhfgM7uyyNYTYDdpyuZzuzQvzNai83Hb9hqOdszeO70KRKQwTxt4M5mE3re2YF1
eoWJ/c+SfhhbBUiWcYW41J7KjaT7/kHVwHL4pV2R8W7sd2LN+6ULh1u/IlZBMMrh
VEGxfUTiml03WZDr/G9Ca2I5DML/GhY9ngALBL79STmWtEznAeWZgsdTC+347l1c
cDYOuoC5G3sZE8qJ7fK6m25OkFT6CEtRyzc6yyGWa701Mv+Z6UzRimAbJ+jK2Btc
DMVjgj7+QOwoHSQfp0Hdtg2DnRzH/tKaO9qgGT8hkoWIBH8uWzo7Fn+vEv7kbj3S
ATWdNmEbb4z/t8GKseDKlXuTEzk37E7Md8/2gT3WOaKQjLQ/PHzdELbz5e9qL0e8
vpfYhYtLIRG3HdCkzBRz0kGWzdVUxLmtEd/IfoXAUgcuQoutMt0m88iuyXqdNyXZ
06n9DBj0JmNN5Qj/3koygtTFalsdGzenpIEWdrChSLsPb0lWSDbJUno0lOWciHmu
9qnStrQXoAxYXEMStVx63Nrdb6GxtkE1z51j4HjX3/U2UD8eowf/81cspN/q6zCr
qZkHInPlk5D+fnpMU+5ZRB3bnuJXw4QyeoBQVVwb2QaIu9Z+nF/RJX7KRP2wLlU8
/nARsbP9M4acEDBZpKsMmlj2OIHz2V6Fq9PfNvdy74jJN4Gr01mt0IOgYM8tu6Az
KJZhH/qDjKyb7Pi6vQtgo+4JbhDQy/werSo0yRPlgbeydr+pg1uWzMxFmxsotepy
zfJddcs2EGqEVAXfzaEoyIKgbAFjWCHb/A+mnVL0kfbKztE6++sLWxiZyan/jA1E
WBc/cveWFPYs0OT6kaBPSS9BESSrJhSpJKRMta+mhWOYumM1qZ+ouHM3oB7bE04h
`pragma protect end_protected
