��/  @9�n�4��XCֱ= Þo3���M}��ӭ�W�8쉂�K7�`�'�:d�%ga
&���͆��h�ݛ���4S��R˖r�	ru�LA�s��oh-�����-�FrI�2��vh�mM7;�H���<Is]I'�#l�2�E���_d�%X�_/��n�)����Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9�㑴�7e������G�L�k�Y
\�������0��q���Pª��Ю`��V����=kK�lM���~�ۣ�8���M�y��f��L�_ʈg�0QA���JR�U[~�+�O�ky�Ccyx'�F&�f��L���Qe��<y�o?|e:�^��������g�L�fӢ!X��&�d�.���`�A$���Y�Hbk��ltN�N}ξ́#�ߤ����"���ȧ�=F\��ƕ|zy�ǌ�2�ͣ�s�#�ȓe���GS'a�������/LI��-PQ=�)�e�C��'z�Q&���r�=��H������e��d��v#4�'��y����XP!u"�g�7��!ì��O�P0E�j�@�I5��m��RZ=;��d�n	ª<,<6q��Y&lC��u��'B��1���L���7p�=>���8���1��'P��
����ܥζz}{����?a]z���am6Ɗo�Q>��w�ElU�<p�A{�oSF'FL_ӓ�7[\�!r���I9�4�jшv�+���6ʌm�E��=�5�Ԫ��;(�)z|����L��0��&����M�Π��OvN�-�]�ɋ�.+	�#	�Mo�Y��	ŧ��矒{ru��p�(�,8a��������B���̅ ����0SJ���4ja�|��]a6�Kr ���@,<Ԋ�\P3���RVĦ ?��z��p�a���肇����'W��Z_��(ձ���y�qmY�h�;bh��c��<O�)���D�,��^�'�#��CJ��w��G��:�V�!��C]���h�S���f�i7b/xZF�q�3���W?}��qH� �fbi~$�U`���o�b�`��!K�x�f8J�k������q J=BT�^㑏B���ŷV�Q�y�lȡ/J�P�ܛ�����5�5�5���A��"��z�$������[[�@-ii��l�Ѹ������fY�ì�m�=��\L��g