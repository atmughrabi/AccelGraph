// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CEpqGZFejkfqNdPLT2E4Wo/cIdXiXmidXfybvkx4/x1WHnH6fTNywzGOHqqmmLz6
8GK8B0ZuI6Ibr+siWHZzT2xS7Mt+F8X8wOxKjjm58zpJZCYI/PQHkxMjWeQdeQed
dMYPCLvZiEqIy5qU3RA5as6/x7tc7EX1rjaTKhNQiLA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2144)
P7Ri8MAK3bN0za8ztScxLUN+gqtl/prAZH4SQ3glVF8vW5wH45H09kG0rG4/2k1A
FG791MS+WM9d88L+5QrFFVqvbPA873CKNMpoRXq+ES305PPZAAPFimfaZc1sXa75
Y3sIzE7UCVIDyCYhIO68v1ErJufXCJwRAG0p/Zhzv4/a5NOGGRzCwQ3NwUJpNFGf
uEZZP1cnatSWmM4cWWKUaTzaNla+9i5xhMUmWN05ce5Mg7FCDmATHYVZ5vlFCVQW
DAr6t2gg2YmhgCwv83Q/D5NQyleDX+Lf2RxopUdZ8EkCvnwQsPELeNNdNK9kMk3U
ZpSbiThR/O2PcJilrSw4hAY3wIvdFfre7cfsCHEfZPGmiqoN6Ny7iev+BmV+Q7wN
4R3rr04TXOxx0Aku9juMzKAabQkVpsnubeMuty8Ue8K0+2NN0OnNWiQ0kIZk+psP
P9BUHISijT6eWRlNLQNgpK2FhS1kSanCk356vV42xRORGWSZR9jT6uwfWeHigeXT
o98x7YS4XT51TnBGed+drVF7FkDw5WyrZM4P9ikKm5InWOYcUIyegKyOZGYSSo/a
PgsAXAkwho/DsBC88RAPQbqOEve5Pm5HEmHuPXxBXkGmgi2wUt6ipFSBbROKjufV
edwMTtgAG79tgLTpc4EaFLJUp5Rgzi9RoUA1YjWYBEdxBuTb1sYr9jFcCWm7qtpp
4I/sJe3td8I5UPArnnWHbSDgM4rlMmaCpBpyvnOTl0DR5j6BUHAZqbgZohkYKdHf
aQJ6RXxAHceNS+XS/FIhPopkZB1LAsoTZMwBrlPm0RUVjGq7W7bYSOKsi06+Rb3A
OLZzDGXAu2jiUkCtE6eYnEKNULvK2nPIKc6UQk1PT4y2JqI74R9EoK+kLGL7iaO+
aWGIbA6+oS356ByktMdEiNCM8YWZkQN568T4uMAplDK3oHqw0aqhtuTbfOF0FotZ
tnEzcshOiHJwfr8/5sIKoP6v62RHIU/YJr80RqZ3+OkSwCarVdvOsLXK6154nrwF
T+AjfuLa+mGm5kLA50cbH2KpBGEBand5JqAmENz8nAEHlijkc0Cn4FqcfRFoBQiF
9/KRAZiyilL//qKkD9eLRwcM+S3JZEASgKOn0PK6fIUfRdAoKN5Nik5gF2rpK8VC
PP35D+b8h0ZlKfjA1tL4pC7HUHTaQGKkTlThMvV4iyuDQmGeS3EOfKwUn5oJIp0+
B/IfWLaKYlEeTyBw7cuzijGln/l8SAiDmUN5jOjZnZagv2w1Vz7FzfGvSVnOGOYJ
kCAJ5et5B69MQlT0dFzHXJKltMkmI5tbEr1hOUCshljKmRJR8ERQywi5mfXxIGdq
MBg6m1VnaK/43gxDCaGQQzN+YQGe7POWMrb0gbjWH2R/Ug/Et50qKU6M4CQc3GHS
uMWQPx4H/8XdQDCLRIoUjXAyHFNG4bF5Wp/nVUzUoKqygeEAgxIlS+FJKUaUJWAz
ev9jOij51WmKX8o3tuvBb+DnWg4qXgGo5jP9sCho1bxGOkTahqAg2tH9sJYaIKNx
xtgVqB1IlBhKjE6M61/txb/3BzZVNdM5UDyo8fRNgBZzAI98hNshhmZMw8rOZnvf
EPEhxOJO2r3BVuxq8B7RQklgZjTdXXop4GH96autjyz3MFTtU0JoWJ8mKxH5jEyT
Fr8/lkWZpqU0VIbCditx8XgJzzigidr30BzZMOcg917OODJSCU363nrdwXfjBz7r
nLWvyOR/TKCRErFj4P/twaz/uvCeSXXSiIqMq6c/Qojc351Dy0VhtVxQirScaisC
WA+FiP8Gedm/Jjo+ICejRuPquoos7bSOv4IBKg3jLTlhal7Ibdt8YGJsC3xnGHCt
N6idyLl1Op8kXhirrvjg+wzti5IjAg0dz3NCMhj+OxAkvjcJdLbpE85m3Sjz/aXr
WJC0QYUSnnTKff5yBkdgoRB7/tVOOPoD9MNl3Ch8zKFxqI5axp33slVnxcoFTYXs
mOG8LEK6DH3MS3eBVZ8RZI35fISkNe55mUD+AMLopoyNRjIgnpM+gQf6hN7MWDP5
OvkGQONo38+Db7VzVqFD+S7xGDmfvHoARoVZrE/MmLagkoHRJXnW9NEBhLhQxXDe
lbs7DGqYgxmFsDyD+b0E8Z6gdTVuEIA/5Tz91FAoIhqMitOvi9CVC1D/v/UBAnhO
LRr83oV2RdQ6Zfk2a5Y6MMXOwqOrHJJcIzVay50CCmAu2Qhxd8/U4KIjaeg7o2Vt
eAy7XCiEUE3DUblX2sJbpGBDnAAn511AEf09UI+wvupvNPXY54qZZU+dzvJCi8lF
RvonwHNuuisONzd8C1YHlNfRwINSV2NDe3jWUI06lqschxM3noT8frd/QgX+zFbz
4k+8+TweGsB7jaHkIWS2MMHQrEBqc8gu2C/UILIvSq3MK/lSYXREC1m+mYeMVaOn
uq8IahV/6krGFXBpoguMWBBtPZ8KnfNxN5xu1xPzcHOkzlM0/8UIfS57NhCWnzBF
TkDI+mFXdwuFsMBAYtfmqzEoYznVF6wnRdaZXQrU8l+RqSIf8GqhnAjgZ7le2LIv
yKxOJ9lKzlb0XnLmr+wxcymy26F4X7kxKHpiw8QCy1if9c65qhf/JDAE/YQnIT0O
C98E51qOss1lZweUs8/trjBZCYPDD1sE1kw5Q2zrizeUfVZ7zxyXdCywnk5QRQ8U
0JFfR4fk6HExlazmKmjmJ4xJclr7SMgOSu6vqY84K+xYzxqnJSch0knmrVp1lqBJ
n7z1yfxKai9j6TvsPdMhU4IA2BWvcsp+WXVF5Pwyq41CreOlWV/CrKYDmWRjYtwX
OxJfpxvkqfer3OM0O0FUE2ETpN1UsZVmaLw0yPwA5O4=
`pragma protect end_protected
