��/  �:7D��W����);������zdZ-��$�d�D ����bG�,�j��F�@����)�o�~1��1G┸�_
ìT��@D��n9���-�}-��o\mR$��s��s�n@w��d>mS��޶��a1q=t@���?��G:9Eng��L��)��]D��Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9���d�85��ͳ��Pn�k#���ȀD\�$�0�����!_L��� ��%����Ny�S$�)v��v�ն>���sZ`�}��x͈7h�t̺��z�É�#��m�^|���M��c�	��u�kC\5�7bYi��J�6u�F��������4�o.�Eu|��fNі̞&�!�uO0�nF~lo�~Gf���ru�4PčG��C����qE��>��h�&&$p���7�"~�_�\C�Q'ӱ݊��Z��T��9Z@�Z�$+O&W�]�-0_��� M������V(�T��\���p�k~%(&����|z��#�f���O@,À,�8�W��<I��ᒑ�;P'��#�7��	{E>���,<��LډHwEѯ��S_[���v�pp�[�9C�H���p�d�ֽǕ5��uΘх� �$'&-i�� 
�؅�Í$���	k��q�_�"R��+��5$��2B*���]J�_�l���pMO��)�-��T��́YF]��6Ѵ�ˁ|t��Ke� 
C}a��?�u����zWȮ���I�p!5ԢU~�9�|���;䯓�$	�7�L���ѩ��H�K�^-QE��5��m
��D1�ڽ��]e1�]��l9U��S�?b:<?P]m�1���o�K�/Q?6!��������:J݆Tg�@c�"S�o��s��톰��ޛ����F�zZ�0@����OA�{����X��R������ק2T�\>@���>M��4n@�a�\�{Y�?������GG$b��#w�uc��I�����.7R@'�u�K�D��3`F��൜�w�x�Ö~�+���-M�*��L��Z
A;�l�R1�?�a�H���A�����n?�����ê]��U`0�U�4�V��9�'?���}ǝ8���K'r�^ݝ��EP�}��0�\v�T�T�,L}s��Zo���վ�׋�e5!T�$k�r��X 0����F��6�NTv�f*A