// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AN5PUuJvO4n0yu72H3lQWMSmGwdrOceh4bETK3f+E54j6YUYYY2Vy7B9WWmsFdxZ
QysBevMIgE1aPkh9q33pgEY+BfjcYAirUfzSqF+aCmFp7VhuhBZ+EipQLH7xZcNH
cmJ8/GEtk/cqCnnUUX68+Q9HrqbFidkOGUczXkBVmcA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6240)
KGRytMAsjcUAzCE9NREPfRuNBFzedYetmmUq+pds7/a65bGVWV5sbZ/Q31p6X15s
8RXajrZl550olixav0inCUuFjMo7pM8ZWkdTxZ/uMMWswWnvfkC/XlLDHsqlkDDa
J8+vFXcATXLgG+dHxXr/NY+F/+nw62Lo+TUM9ETO+MbWYjk+f7sUbBBtzPNNvDrD
TvXAxtpCSEAnWkYpk2jR+m0UZjNzhN+Ii/EfHIYXK7QYzQSc2lhHRZZOHHPh59tr
tuGCIvJw61FD71U4KVAap1P62WUm+0HgkLLQ6rx2yLryya00NhxYvrT0LRdkJSwl
hHk3opNcQf3JyaD3nDBq+P7ZNPvfYp2xT/Gg1Jju4d+kAwx9w8C+7KvxblUg2SYU
+d6Ge8vyChICrzEYux41XROT8NUJGB1BxyXzhR6PsulK/XAhMI3MnjYjC7BpK6kV
jLNFU12mCnA8pmNDgd9WvMKKenAL47uwzugy0GdhFLBYOrrz++NnvOK9R+oJHYlO
GYPhff+susPqWypJkIhXvLQBrsd411TawwtYY9GZTDtjGCpXFAmBVwk/IQIsKZ/1
UbsY+ptvDbceY6UrAOx7sSmxnZo5f7XpHKshpPg/0JWFgTLk8yGhJ5Z1w6mMmgqD
vgc6EYhRNtW40YHUISvK6xOzN+txSOjCsdjnFxYKXChQ7Di/X+bbis3gipyGz7Wg
yKtBE8or716Gmbapo0EfprmFfZXi9iOCepFdM52JvVK0E5Q0umzm83eF02WCt74/
o81j0lUnWzUhWY/QiBEuwyZeKOp10RqjciuJ3BHLkTYjRJyw3j90MTdGsQKkj0Y9
ziOo9TVljNlC86SG2U7f1vHUMWW2Vvw8lolNBrfwyl3X17vcKdqDLFDiEn4ErPLw
bg8wWpNUGOkBqU1p3/QaAQnT/uJ54JdlcKcPnYaSa9bJRbd8asinlG17hWpQZbhs
Fse2QnLyl/V/rdWsbhV9tEgVVVuDG5QM5TTxdekadMqLrAf9XfRrG9CkzF5slRZV
swXJ0BYb79oiokG9VJtrSNFC3gvrq3FDEtrWPcpkkSb4Md3J0rHxDgVBQE1ApcbA
wgpTbyQkYSDFEG+3bnQJjoH6/NkQwpozDVB4XrSM1S9WXEwSBFuQOmRift2fLcQ5
AeJ+jqNe9U/y99e7FrEX31k11gJYSzGXifmEUYRxf6GcNHTgp7PySosxO07Aejlw
QpgaC6LkbJucfoEDdf8L04RFx69gCBH5byspmpFTouLIMk/q2MgisRLXXsz/Tcfp
c3gmfut45DVzAPxaggqSwPpnqM9DLaDFrkVrQ4lKDyiS7rEJxhf0mY4xBHKDbheV
tziHGoqPuoIcf8YCujx55+izDlCkJepk9GTDrBKdYziJtv2NU2I86ipgHyGZbe1j
SYcC8/fC8FGi6TXyZk16q1E0VDRZYXI8UyVa/e+9+rpcP0/wKpObb0T9uN8lhN2A
KURWLYL7rHfEdydnsnUiDg1+eT5+Zmo52DvrUkZj0VS8hEeCtNtnE55GiLOY4jOf
26zDJk0wQsIa8seuSNn3UD/h4BsMqAfykFccrcnq8ICD5Rkxdn4+y6yweO95fN0E
0c4bYHEgEZTDqQ3ChdMzpNvBnvb6dGGrGzQlbVl1QJYKZ375YlMtWgtduEE1D3Uw
mcOjAWrMPpi1oEIgI+jYLRdSPPh1T6IeJnYM8i8OuvnONW4T5B54CZ5EPDZk+CGA
LHfe1/+Wbs/Lst0Biucm9oFRdzLSGGevHDPTPq/Zb6DaDfIJYqbbnflEGKVBQ7tt
wTGsz6sqPf0MolkLA2wZqU2wO797cu1/zElb7wkU5jeRdG6Y4bZE9gyTdkCZjXKA
/h9a9ujvrbmvKEnPI6e2yfhdjebAC3uDkxXM7JXJEVOvGmJyxEe80tVv/m2XEGs5
Cbx92Z5m1TS59nfQcABLt3nyjlvgIyxIru/sobPx642JVbVLiIPESDbyaxQdTqFq
PtTJ5nU819rxqJqRvalW52BSTMPmHuQFtkxprOmV4CEwH2OROOcLTS3ls2NpsV5+
YqkD00R8SwavpViFVebYBh+jaQYl+HLkt6nEsj34tJUSY4w80/+WxuCpZzRtz/gP
mN9oXpRQzogsD5YCPeSJYVNifPaTM60ZtvgqH5tBKfAqdjrA4KtAPhD4cE1O/MmB
JAM+JXkC9dOnHMP27A5/q+doBGaK5uRQvYXXcYnYSJ5hTfDnJdyzhEG2t/5JuTPg
QzQZWVIqWHOo5zo354TiVOu4j9ofyq9skNgArFXriuaIYnlGhg9Uz5L1EqSpyQd2
Xpw5Lmi0+hvQdVZURqdn2nh8amFTCQGHAUcs3AmEuDfLOjZCVFogObm2dkEs8Hpe
dcW3QOutLFpIfHLnYtdP3lxnhaC8ihXS+nQzdre3t95I//XPpcl5tok2MmagaDJv
uEE+cRTUr0qDFNjV9r5mQnsHpQemlnQm7V5bMtynYsJra9vN8Zb5+AyCViMaGX8o
AcncPy0s6wjSIEBd/cAtIlyvP/oJQuA9BVvQVXMvOYPt2NsseHIo3lmIbQatyP0b
9i4/GbYUahSN4GxtuWUc7MPmN6kRK3SZq9ILLQFBwsgfLSSHyc4l5hG18LmqpXWZ
mOSwDulD3+pRgFUlwW+Uqsnbj8xj7X1nrp0201W518kuOi9BnwIS29omZUhKaWSQ
uJ6CCpWVyAHg7YGsRqSgFJH3EJFqP+HYl1+/uFPhl3eYyoLPbWpYkUS3I1a0CkJm
0uL95D49QfmuoXQEz3JYpqqY+bA+MgOvnjuSY1SZreCwT5s/nY5qn9WZIt0P9UIG
P3xx8tYvF7c5iZ7pEZ9z2Yw9BVP2ylueF1EDWnHSQVR3VrawPfd3aSG2EmYyIJml
juErkk1scj1UmWWBXGjcJ28RY2DtUQtgO3/s8r7rWEm0HULPp5Jx/ZU9iBPK1w5L
JOgePgcMVCTj6Afs13sk3ZT4T73sTUyJvkjl+d0i/XiNaTxgTNzqIdOg7nNdhzyC
7pKk5ZSM/cUSQ/kXFktTIyMZRfeFQzwlu9hTZWQjqRqsMy/dSDjYXK3TxLKSYrj0
RpEFP0KuPO5ik89b7+1nBYDFAM24HR6JeVfN4dd1I5zFgWjIIUpTR56RnAHkQ1DH
QpbDBY2/I14Ubr2L0XcWJC+uRLwvQgQb7PIBn6BcIeWngyA1Z7dHebGTsmCl2HhY
DDRaKY3vEiaadxAnhsxlAA0aI5+MR8mZGRdtyS4yWxaRmCy63OX89ruYGrcLpm+H
QsWs+PR8kcupjKqR3lSkb9IDaVf/lZDTEhPuo92juAHEoeL+20bymepkWbdGB9eI
IEUXoWQXRXSmaavHREPhWWqgUfHFaoQAm9oI0FL8C2Qgcn6hiMOBxrXwiOKfyZUK
X6WsCp8AS7D2YmHGuUIpmMC8zfwZ6e8mebxuPMwIEUvi4+gQqWHM8gHPe9fbHNnR
99aNQ7MyK6HH9kMiGkLvCw6OOFPcjU0SX1pqoBtZBNeStSWxMftkLsTa/oT5QI8g
eBcOTo/tGcCxn29/66kryNtpZqFAOsOHOP9sK+iSsY5fEUyTHzMXEMYcOL9v189i
1IEGNQTTgGa/tT3cf1Xjb0cynK7oxvRyFWbwzTJ1priHWQBmNlnxpHERq4nMC0JA
hBk3TOkC41dIfKqE4hiMfZ0KLImrJKIWhRWTZcLgHPQOCvtB7H5wY52qd6C0MugL
3y2f1bz61UYnaI2L4AFkSssKEt4r8dmaEkOObY2sMLWU7Pw5uE763W29CApKpP3Q
QJxppIxgymyBDR76UUH+PQRkz2rLMek1mtr4rn6FCn74PP3CYJmV7IfoF9remHsD
8RN4IfVoYoKI/WcRKuOKLZWTNj8eNLXm6Qmd+LLda/ErjrSv4ws0aGRh49i1wNyq
LB/Y1hASgZhQ44cA8+po8gn3NC+r+W3efNB1aDPZqeTRROeOfVRCbH0dN3YaBQzD
Xk79wv6VIMlNLFazIATgQHLpn4BfjpirK3tIeVI8I+qqz/AKK9Sqk/PMxDnwbLNq
2k4thhGBuhuUqqaDiwa9Vl0CGhie+gP0abxuQQ3mgfHm7nlpzu3Kb8dBN6bb+XfR
VSMigET2vDu1ROdM/jdLybw8O2UB31FKHxWe+XTeXUapOmJLnOZBMtgKmkw+KfJb
3NAxi1R5AGUEt6ljA4eVPsaWew9o5SBD+jvmnecGKtiBfEjdKh7ziAaQSB7+1ewv
qUhy8VSX3acEzicCTqbEHw6nA11jhjwJjI8aI8gWIzWUVaTLNQWXT3b+11orHWma
OqdVSYuN7rK5uUE9egn/Ja/YwnhN+ABj6owe9UVyGmRb3W+K3okoZpEDTbcSdVUO
QAtC9aN6U+d1Pss4ydMGqICeQqoz3mtNuwGCqQ31UPbVmSTjMJ6nq6fX0X4aG8wW
Xl2PdToq5IGcwMMV5k2SNVHqUs47dDKTf5zqiLE9+TeQZCNqnrQXvGJGhjlMibwe
LemBMnNTxcCE5LuHWaNx7aFFSNxiAwCJN91elmRa66at9GiSwNGcMYi7rqbeDeh+
SHRJ9odLYgvCjuzMgoiaUxwi7IzCURK9Rf6jpDofcQnaSQ2BPO/mAhuDhn6cfIhs
JCgT2j67ltnzH1MNT6TeX9MG7uoNcGQaMC1IZwONbYwAuClWh+GaoaMXegbV65CD
k7AH2QWJ22B1KIun5Lg0zv+arZDQeRkYdw/d+arer65THU4RUixUk34Xdsq5m/Rc
Xw60Kg8SNP8eVJGm0GFCM5502rQZ3kTwaGs8otvaSHIv80TvC6YNe5AGDxI+aOy+
GkuOoJkkLzyyLv42zWhPAYGPHU7uVphWT9HQexnGGzM/vY5zUIAWrz+bkmUECTe3
znEwjhIVpPmP/5/PaM/k312TNRnIPvj3VNEkIRV14usbfxQiQO4danc+J4j6QLnL
naFvw80AlGZ4DKEfg7Zn+AiNewGsnvJPIrwML5L6gLkhF/4Uj5irY6AkI8jtehrB
GOcG8coptKqI/0ZZFxOggj4CqAj0p5aKdTdR3i3SHmGsd6cxzRgkavQkRW9Ix8qo
BYGhSNBeX4oeuHeL9RWE+7hk8cQbA71MQb/v+I7yITaaWCJzoDO8Z4RIuP54/w3s
B1Tj9HRgcwq+c7t+6YDI7ak1b1YfiiUxYsm9CXQpmYqyHSld3goVh9ISQs/dnNEo
EQ1cJzFyP/u6UeJfBnLy5u9VKDR1EBK3V+EWGZa1yXKMJBhLacWgrLor+mNKNUhF
tKa5c0s5UeQXV6FZpEkCpNjuz4VY2GnVuCYtjnaUO0Rid3bXh/XrBiuHI/kkM5SY
D28E5/fadZ403icoz697fGwxTvtmymSA5CsI0JFAoyT5Tb9zimyXc2p8O77I6Rmc
VaR7vqWh/ozuHVB0as5ox+WY9bnthMbbDcRYVwVeWdW2lw9XOw9melTYMEBcweaP
JaQavYIkQQTSDDXtaOsRw+kWvTAmUCXLuifXnqLODvtKKRgoAt4h6BuZFCVtoIRz
5oUolZQ6izdoOjVuJJMAy/R6NIM0o4Y8FVsyw3ust+u6uASc2QyUA1dxDyStUixy
ecMMRUN0iD6iyRYR8r3wAx3rmWO2Cx2OKkpm4nw9riRe5dT+hQKoQkDp5yaQa3vu
AuRrxCEaHrtJD2Gdlru1yg+da8trgQ2IK0HomfabRdr1geCX1U/s5HlXAi1SBVSV
pv4DSaJqoPj7SQ0mq9NXIkM5AVeMzRXhYVvqJDYZFpuKsxVh2s5NvykNrYikPeaC
Oh/ZC57uWIjXgb+KVSTg93wjsZWvjeVrssmOLeqOQbKQCTnD0SYt9BVLJP0zlQL/
2fRxkUd6AIknSPPE63RgXWLFwHBRSgMWh20Ka9IvZP/8Td+0Za+CpfjzlQcgKKj4
6Y7fsEmZS439cmU5uYViawk94FkCqfE7tlR1c8m9CGvyaLxAXx7hGa8ovcu9yJwv
O7YOzTRozbA43iQMKTfTPinyT1DEzNpHLkYBljbw0PbpcYC5FvzGHQIdigV1mMyM
18Uoef2thDRaWgFN6d8AxDS8pSFcyRGAFAjcml8M43kzHs054ZOJKwDSN4uNBxh8
m5nfxVZ1scvmTTeuCl/WTMaxlJUwrfFvCgAvXOmcNzl2m59I++uGY8TnJUIzvzqK
FhxDKWVtwm9HGzMjdXSUbb5f1vfT+BcRpvRmGkOybmnfr+AtZebAvhgOSDS61Hhr
W/fFssJI5XSy9dgogAmZ+b2hKeYaPAk37H51Uup9tAn5yIbfxNVcyaMD746B2sET
pMMEFBMSExVHrod89EhI6aF/RfILjZWDxoTPh07rYCY3ZgprQhK/zrjyWgy5xJVX
FHKNSLFH0bz9pBHSUfNbdtCrAUrtWp1c1Sb53YtYUEgNEFhZxaYuuEKQAEoZofi9
Xm/F/jzD7GIAOmGK8YBvKjMcCfyOMGHJLCGLutQDwYmSdTUNIOcIoQCmDWrpFU67
iaURExOzgC97NEg1iW+VKB3fk72omntV6ZgdtEWzE15wnkLE4g3Uzg5RjmOC53sy
RLt+/FTjnRPivUnF92UrxJu5EGs2CvG5+gT0kMMlOGXceVdKt4/flKFXjlb1XuGk
NSjWV+8T5pbU0QjfCNJzJiZ0SFDQ/+6412/9VKR57C7v/fCYO8/anqaeHo9UgwyN
tNYnzeiItVuQB7VMTpvtRVYjtAC1qcShExpTpWC9Cj/g/VJCdh52FtnaIQPuW4Gy
vHxb5JivY6t/U3yXO4zNx0t1huEi0xZDMnfxAvid0w0B0YTMKsHzYqqIVEB+AYg4
vSLp1MxcVDi+m9M9QNwSIqO3INFvOAhkV6hh4jc6RPTM5Pffzx1w5q4i4580/IVn
ery0qUCw79t1UER0fjiZrTSAWSTb9PjppOSD4KTmbcr/BWMPO126FgtB2PuW1Qch
t8k5d/8URF55GWeEdqtza6mwzfCc1jnm+yeBuBhGlJzdiHh/bfNF5ic4oo94XghK
R7EFwqCMIlwBF4769BM6eeawHeyOPjROuqPJH5WQ9/EEIByTKmG4oZCC/kmfDDXJ
nriwUInse83wHGVS6UX+tyjJVSlXdgZN1Elpen2caIWd693TDaOVH99UBRYLkM2D
DBEkWry5Td12LpWSFGHcynPFc2IYK3m4n0JrZYu3bGrM/pdJC+js10Zk4nkHbn0+
HGWpsBSfQ/RL0NRdF+HuDTX3cNboxEh4eSOJYkMIiKWIYUzzN6w5LqzRqSLd0bl+
uuy/ASXG2Dioel3YjEjrkhOHZVVAzib6BiSrNvWsvHyVBRZlSHu/AAyWYltJz1Om
dUG1yfHZnf1HfmUhYqZZGG90xpjsblmWwugIwLDJ5gE0KDKjUB9w7T47KF7oCTIr
QU5r9OQC0WaLsfX7n5u8/0YDpsmEi4AsgiF3m3YuBu+ianure8TMUae2dJA9yiWv
r0FAN55qL2yKF6+ulbn1W7zlWnf/tRfIdRehC0xROz5/nVpWk2qis5L8OavgLFNt
vYels1yVpF9fnMpA+1MayogSqsoyjWOfVz3X8uCldfMZpvuYHri4CBRAkgqup9va
+mLcJCx77uTfHTIGKpReF0wlcD25DRU8ktJH+ehY+WZcriHtYycbxo8Ke5YUvJfE
ZxsuowUHXi9Zj9OEOKJimGM715RvWhi3zmB0wb9UBMVWFJHr0SiEG4hSi1DvDUNu
rvaaUWyVZA5Ilghr180FUKcjseN9V1h0FLK+oVfZKqNjr09813j6TnEXWWObeg/u
2kp7BNrAnwPThaw0t1PKU9RgGo4y/CHo0oUt2lefxYyj9dCcBPnhkpx+cSKkPCE6
5/2nA8WW74msp4/z73271tnS8l3mfSFmbudKQGGbgoMlgcJb9ZRDdL5HoQhxQjeS
lOWTGGsHe16ZzfqUTgKeOQgIrpZNy4hVdCMox4b2NAZ2nR3AHihu6aMNdlO8IkTO
FFWAlKr9zaYSs+6zjgnTUkDXSAqUUi6szWC8WsY6Uv6Wt7fbhpq4eoNL2//BqsUF
iDzFWgUlJiRlbRXGL2BelFu3QdiGofDTZ6eERLC6y3n/h2ZTeqlZOcETlXEFGmvJ
PXqV+WpXM9ogwriRs5kNbYeSG8DREfnW8qe7E8yCNbM2igAUoQszYr5G4pvSNV2t
wTdKdPnYY2GCWlKZE89GhvYgVTADApXklIr64Xu8Ha3a2VtLvLRya7bjZgJW4IWS
1osfRsjsejqBVq1EJRYWKLjP6lh05XOZ9FvPy+dDXFSqgKbj8FxIcu4nFZdJNkxI
mzxNJa2/hV6y4+sMRKBzzoVLcI8U+EhFV8fzoVCClqdNW7LXALztKgPUy3RBfeyZ
`pragma protect end_protected
