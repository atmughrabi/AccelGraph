// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mD1WR9EriyqDkbK9+uVS7z3ZOohte7sCEIN/BFM7PxsVGFMVFQPkO6hYIa4MWmBv
ARJNCY6LhwBPmdJSTm5sy79Wl+Z97x1SGbsNcm9g5KLTIkUxnAL7bRSpUesYZnpW
lYxMDklhQFXgv/FYV7WownMhX/YnEKKxHJVUDAp+CBo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 193744)
y3aM8QjG3B+6MkGm8hGxdzcKgwX16Caic2snAyAar87AXWTd05p3V6UQyEShLG2G
V/l9n5DRzv5HWbwMXcUg3s1HEEwwFW2vuWg1MLnFpheX8Q3c3JaCCzg+U5fBNhN9
dz6ARb7ReWXBfilaU19pkTZXzEaXPwhOPJOmCviE3fZMdNfVLlXZG60QT5bSb045
4TEi7qMgZ4VN6ugiSV8IFMPWGcw128SCZdPA2q3wzqSoUjrXqEKgI2mxiEAwOx6A
fNzvhdgYNw9d0TQlItyvm8XARafuENH+yHmL6G2YFxb6zm/S03rv76FUfavy4wsi
3p/NYBYplTvtZJcTs81ccnKsOJYa1fIE2BzRHMdwbrpeDdzTl7U+HtlFEY549H3m
3awhGVZ2iUAfeZNnjjHrDPuQxs0QBNKzVu1SzlajFPaCSrr8zrbh3n2zCMo0myCO
3oXhYqCCWB8fd0NYt14TBknip7qw3aKk/rRsh6jyutHG577zLsS3BUlhlS5QKNx6
2g4zMverRGwrDBMzRjC27QUrkDXg/ed8/QllhATmt6fIVP1inGRfsOSe2zxxrB9c
LFUYRLXtVc/cCLWg2szB1Ft+eqpJKmedKE+zKzzQOZcaRmmm4m7NWO33+PiomV11
ja7A1PPqwTcJfWHgL+NeRZkMHikZ1HocIWMl4nPE7SAZcFlAsf6NeNVZvHU17p9G
TWJnS8uo/Y0z8wQlbMx3GdZEMSQXbpCMw26teYst603rRF2fzNmRHg0g5unf7NHw
Ldx7QKVZqBTLlBCrMZWm7by/VTVYHicPih8zgzAM7iqEOKKuXpwazl1m/BpjauG+
eVD9czP6m8XqxsIKJeP0u/Kf76n0/Yg8Az6RaHok2FiYr+qZiTRix0nS2PTh0NU8
GhfLjodGUpv6HGa6UMhoKrCiK0Kuk0JaAjKwuynToRMGIOp8WlizUb1vsGn8VA8f
FqaIbUIE/LF2iaOMt5582SDl15yRqO6Tr5CMHrhB+LLhL4lzpmqL+i0C9K2rwmjP
bBL6c1H248JHsLZiDhYiOjh0amgLSy7eBr1nfjPBXKXaoOSrffWvQn0+hHDei0Qm
6pKw+MPDh+8HBzpixT+p5ZqaXUTbaEpW78dGZjNz9yA3db0g40FXefoFrI2xo0Bf
s/v5HRUmCEL9bXXu6a2wtktkZRbgZdW2SSu3vKh+QXdn+vKIuX6xs08FCtqeCYKX
yYvcVvq6qa/DP+GUf4nrL/XLwwH4sTGKcU1tSTdwaDHO3XzKugpvEpHr3msF6Zqf
7dJeWxTVKE0xmg2oTs5D6gUJ2thjA6U/K0PcHocdYODGOGlswtLObwIuJyQAXgaB
GpVcsi2SW9R3kjhppbLGxPGo/BoCFFhJ/sX4jOqmS2oFGSvoXnt9WKloAmvl8yhs
q3ZXdWzt7U6KJvn0UGMJt/+X9Pp7WPcdHu2kHQZg6ew1ISrcB+j1mAUGIpZuWWU9
NObFE68lbPRacSv+USITZBBoSYZ8Eo+Ovzg6ZsoiIWXZf8l3+UjulGQkKsyUiawa
tvWVupDLOLL34C3uUWD/PUyHQz7QqB58FbYCV+PXHfyA0lsuh9jK5RkghzNOvKhv
qVf+4F11ZAa8Ri+zwzV0CeB9GKEwwRzwYZ7TPMtFDMG60T8Cb0wLxikZ/7IdcmOX
UQqPc7k/sOmUZM1tcblwpcVRyPUAbTgjdnPpJurCiFdxG7mwt9ZbKppGs0LJPriN
ghkgT6U0+AKSS+T3usMjh31y+JziJG59+WQESi+YuqE64oSAtAoduRpl7jUGFvws
j5HAva158jKTxJ5SW/8CeRdkvtbpc8xdyL+zPMGpJXvQbRHyboNFeiPWKQV0jPbB
25ir71TengrJsyws9lfbt4bPPn9X+ZgL2HQpbgY5WXEOy0Hz05kRBvEH/pZcDmjF
0rs8CyM6kokG/3POtnPjK1Y0wdeEBwnVx2FA0k2VxwllewA2mgCme6SkdwMibGPt
7b37bzfTJjWhmEQTG8o+Tzw+3QumYnxzkFsXdBbgQETVGicwRyLOfTll8vxYgAlk
Z5VhRHLJfHY0LjxLrdAQx9G6dm5KIKjEB4zRCEoZexETh3VG6Duz1AGZFl5skpI5
3fu87hTkLklclh9cmQFZbktdXa3ZLSQGdz01nW0lE137ucsCDYiXY2qCpgWb9ME5
V9WnVaj8UqjwSc0n0Jjl92TWcfzGL4h1r5pAu7UVEl80Xj/2DvHSxyb2DtpMBiY8
kxBzNWQq7qKR2yKfBq5QXv3w+rMOInA6azVQNpFnB8U3+MjupA1riBRFYdkJ+3bg
7VyoBE67EWwe09h0c8NNWurObtOJJtaotI+/MfvecY99K3P2Dn0A0N5xyEJ15UV9
GKQhyx60VFz9wqHIS+CxxX7ifx10uOIhHANldGahA//khhKWLBjex/W9aok4JgGZ
W7YMzsFpDPxMm4mnUMMo2P9jp7LLDJoB5h0zJ90gpM0uzuX8KCMiPE8iWPdlZNY2
l9BtdwGDtSynw0taXgtRLfR6YUgxmy1zf+O9EMgEvZ9Y6KKfLYuo7o1zr/Xm2FdX
xUKEV3BmeWMaVeBFLGm30uH7KmbJC9Iain2pj8UWKgKfKYwCqMfiuF9E7CIwnPAm
RvUH5JqSCM/g0O7eX3iPG43n6Nn9pQa7o7lGKAln0oVET0iONZsyhChAMJSHfZT1
C6QFejnCLWXix7pKfjtMuRA4/o63f0JvTDkLAf6AvfbeMtp11+LbhhFVyFmVAatJ
fKG367rzqTmRD0lVbH/twZKIQFogtnj+nCgNiu8ZFsRkqqUww/EdFGhNOP2LN06Z
VwqhDdreUPFaGm8iq9jfJpIIlSr/H2KMKPGAm69YOLcI0t5qow57LBm8wHpQAGYp
wcqxOc1BeNl/wbdCZTXJNbWjBGO5zReU8tBw3Sznb8fWW7mPAV8dB0e3Zvj8lpgb
YWGSQR3+WCwILQBiaiCckIrSKCdUE5vGzQiZso0t/FbpdK/yeg7RQiKkn8f+Zxdv
FsITZdMRR4gSx+LSwJQItskUDuyLVDWQQ1wHBvQsmnK9ZYDnakCGXJqsVlBITb/c
fOvQP1e9EQbYyrD3u9+x33rxHsaHFBZi2u8SWV+Hq1AQC/p4nZPS8WjP9BBA6XFH
mW2AyNKAaSZp2ZxTzjNKY/1a1Dy1ww7VejBaZEUFJXmtGnjb4bXUV7e2zUSsYXnz
okcuCEKnh30RXslUZMtMHuRqkZGerFXupZFoD45wEFr9SQvIKacTlqW0miOaG8/0
OL/gmfYjwNze+rKxN23wIWioULJwCen1MugcCtV9RKsBkaDODbxJS8ElWo2qZHXo
kN3oF8qj/F3vl0nXHKQOc28Jh+Tn6qGAd9EfN9jKzjWNUn1F5VP93PImxt/TcdpG
2EQ3p7HZeXBBqPYXcXJPsfxJLa+QI48OwA9coliuP6aYCV7zfeZ/EKJG3l9cc3ap
MAaE0VChmfsVeI8g1mDiIvjakHynQFnE+5vlhRy3pB9fSl0Gm8af/bbP4QevunEu
MeW6YerKg6m8W8H36AsDSU4S+F34WneNZEClb4ihRWmM4Q9OpNgAgI8cNmlcflv8
oFT3CjAX2J190sZ8f4EPFI9gKPAuuYFExB6Dw994+LZ7j/NSFZjydiVZfHJpNzYB
q7XBcfyb00GLjoVfmtGB1RbOh7DdP2d4ilrtAqGwv+h+lWhaHkZv2Kt8MPSn+AuZ
dxX7KJxUVwaIh3wRrmvCSqGbZNgWOCY17VKaEyFX6INo0sDdoiQudSlt3MXnMtc+
hRmpnw/5zfc2KTT+VAo2DdHOmpH394Sc+dU8SeGQFTVmoQgw07WTKwCubIqTQwZV
DqHHagKW984rNO//Ku3jkXCmn4YoglZRx+IVrAEQ9mbahIrMSMgY5BJ6rJHTiPoI
MxVMMkXW4ZPV1Zk9Tz0tX5luakwfAdB/B8EtbNEZKW+d+8KqG3BAFiJmD5YrN8Nj
vjB6TqGf3dcstVXulrXGRhjhVggYi8Gero0o7inEyfJIqIm+e50JxjbnXjBSWHnr
Zg5DjRE6Of8XaeuHkxMm5ypyZZsD6C6HmO9tfWGhcL/AuX9iikkQakG2uCrzhBzS
hp4xkP9Iv5euryZuTQHuPQoW94OCJrbVzI3IIaW5Nyu+P0lf6FBxA8u/EPYidemy
GPA2Dd6SDwzW2Zpq1XM5zkFy/nXjv1VUbPT3zXbfYGDXpUgmyZjdjqdGbZGmiZ+D
MsNmWhGg7MUGh0xfbtwDy+nVS21txgKdUQpC09LShAF2z/mTrcQNXasCpr+nSeWU
Fg6p8nTdz4/P7qmV/VEa9V59rS2nanMj5ZcMXdf1f/q+cb84dIGLf+vfdxdb1LJz
mYJn4wc469+1u1am3vLSKY1K7trzfld/6CjC0b6K0waz7F1ClGMaV7MPd8GjgrfT
AToivrE5Wa2K14evdItSMcHBpnHoYh4LHcWYHcIHk/R7Bj+p7MpHUh31FyXbCntH
gZ65PYCmlmr+wzmLr7u4FnVJ8HHcDbkwigefqVIkc7LousJHuMVfPTJml4OWS6Mv
yv8W/1IGoJPpCaIWx4jWAeXudeAjC5pguNoIa+dLZRdFILPE2oxA6ujaEkSIzCCj
sT0Leo3LKDZTClABLYWrywGBEIdcBzAxCnh9H5pNzOpjLwbjLnJ440F4GGOKzRyJ
BjfoKSIx4JkYs03gFUgsiNJQ/LHwJn6ZyIfMgPdLViMyxxJ6DJvqsqJ541q/vnS1
lEnsNYupEWgWLIFdVCqPh/5v8RiZIayX0nfYMiL6Cc631lYgg2nZPDgtMKTP2A1h
LWEDXMYhwdWLOJ1Uga/VCXQgFQyxY9ZbtGj8lOkkzJMDlnsvqQmFgezE8PaS81ma
0jJt7+rQEEPtbzkbqE5a3fYILSu585scsmyUF2Z/QvjDLYw4QXDrhAyIlHUZAyAQ
F3W491oDlH9WxtiX3XE+gzKnXxDDS0s7sfZ96yFWb50/DutaZXE5k5Eqs2ilcmSR
eGHIpweNXa/cEoAjCi0H0gGpWOqej6oZF6YJeWQDc9DcfwEAjAV9o0SQ8qGu4wWS
sa/qwWH4pMWx6wbHpEMKyhmcJizrZJZROMhHcxGE4TMS8u0duuv8wZrZ1wMRhQ/E
/jtI6utpHEw50vpPlRK1ONKYk190nCqNPLHSvACo//NVqLmtvzySacEKdZ8mtqJ2
0v1RXbjHO9HixIdpCE9+SBK3N3YUGYmpJoYt0dqrh9HPxSESb5da7TVXZbpvpTAB
pRMv8Sn8qxF0H/IkN5VNmHpzwZSIofY29XmOzCEuE3YW2IhqfSvgYXpkADgpaAnf
huFbUEIhpjv3530orWkUK8vus8atLyPKwL43u+XQm73+ZopFRKHNB45SOOGjlgcf
Z6oYvpSnH78MUwU68Ptl+1LkaVdqKfVixOdVn9gq/ZF98YLHsbRKEVPuNSGjwlEq
r1W4I3ZgxXyH6pWzbwhrRMyDnI+0s1mDt/k93I92uBAzW0oJ7xwFg9xB7PZ6j8yr
XDHy3GM8XMNMYL6mqiCK71G3B0Ygv3hO7UKJEI/WzqVXh+SnofHHSZFjvZCF9lK7
zo86DyinauJx1wyAhQp7RnQyGf7UjjyodPKteHjtAppxZr3njmrV8T6ZlrPdeQQU
qiAP+VwoTGqNhi9AIdw6aj2WIDpEzZzujYd7d3t1RWMl9whKBUwhTUcpeDNxSr5Q
BGFa2KM0hVQ5hNhqDpE+uAwtpM5bW0yMWZ62AYrdpkBnyb8Q/MLR5qG1xWO9wk0B
mQoVcVMbt8x7y/xK8d6v0BnezPCbXpW0ACC0J9JEbDubLx3spZT1TiB6yAL1Ttkn
c8brhqWVqp/xQ1pcq8JkCeogpgKDzff5/UGy0y/Fuh6r+TK+QfYM1l+YGYXSuKhM
WPLBIO/X/rAOxRkFm+Uvig5gdgFce+qxO3oj25+2Q2/wa9U8K3/Ec6tsC6cOHUkL
aFMy+ZzbrDGB0+KzoRCd0xrpf0d/LPs+rntGq/TB6wlSu3kmB0EVumuQBn1DmwRh
E+5285eWRNzloJw8si4rOcctPgI0AuupRcN7Q89FAo2rS74lXSeP0WijRuDnZxx/
npwCSkWqFoZebgkEAfM0Wz3OEstvLV8GjEQdwLLWavJeZV1gBJf1nAsC1FVuzb4X
Y8DuViURYvSf6x8DQnkbsAE6KRC2IgG3go0GIcdS8Ux9uab5n2u52iKHcMS+YKhq
7PU9IFZoxwx5PrQ5nL/gpgHnzYu+KPUcwWoHvEoNeSKRt2NzSmz2JSxF6aqnVs0+
6soAd4JuTy6MIHbzqpKe53g6PROr6ILUXrxofUvLOrf32MnoM0Ui2Ll7MxD44VpV
OEvu+ZmgiLJQcqltXgSARZFvso2Mz7gdW+vbJQf3LioaFN+ya+3B5SEtyGtjKeWf
eTaUD59twY2mqTWx7ZQfK0WTVJxlrZAJyNTOojc0kevwxJJYok6QVTp1MkhEYA4w
PXq9Gzbg8etFtcC0zy7DVSuD9Mqs2a2ISqju+EI4xuApshr6pyfQSH+bVPmzfYDC
dypne/I02LzZnuqIPIPmAE9b4T0wPyw1wtoQu49zTfdFo9QAeeQu1TUU6L3tdNr4
tFTVnvtrKeLbJJT/KYcozR7sQyP/EcCMmwPG1yHIWXjm/hvcII0f+ne90YnNsp9d
ueZ7fPuLxsupu75nW9P6yexgRe6aRowcqtMJkhJ65pWQxV4K72H/wUM88/CX7SlV
ic7U35Aql4UkZm4ZpS6nzyvHX7rieXTXldBJq99yxSgoQoggzWYIJOOtJbyEsHfV
fbc2F/rx/ns7TOgX1iJ57zfgAla73TXOj6choCtYzrkOo+DVbOfPNDBeJUjQdg11
CJ4KZen0d7kRLACtwEw0Bte5HbT3nR8r86AJe13f1nmJiR1ZG4S36BeJm39yulfs
cM8Coz2VB7Gyr4jrZXff7nHRR3nFMKF5Jj4zpUkPZoBDP31vmqMEUHeHERAUd4DK
T7yiDygwl8WK1KMoro8y7C8am3yBy+xuy9/mD8o1FkkZZHgZ4XPtvZJ+gHsU4+gR
9VXlrCBGqYlBjQ0P0IwDcKyBAkhbsg9zlMNx5drKCUmQaOASQvPM2FVJC213VvUH
QItyFpthuYXO+anojv766RMkWi2K43BaDiTd3wghd+koEd66qVgAV0jIYetM3PUl
hoODX1aVV4lBudYvcUq70t2PEDqsaxviVBLf41DLNzT8sRToQpQHWB6sOrbwTPeP
EBcJ9Sw4h2RpeAvcWcJTBaeBhp9QfDOLRXtMHkvDN6uiy4+sDRaigXsdVUd5EdPg
qK/NgNw57OlxbCD6qp9t+wuHbqZuR3+u8W/GPFjdPiJ2N1ujVrnonnrvXzP3HsOn
bwA3a3refemncoz7gj7HiCNsSzAkGZfrv4r9kVw040lCncoi7+FlEB0FkNGvV/83
6w40rI16FMv9SFvqwDaU6/iRH2mNE5RTRSVQ9Itns0gPRm+PrqKoHo+uvZ0R7Um8
zUZjeF5djNC4xRqODH3n9ZID6Ld03UhwbCqXDLa7rao4Suk9S4CauQJcXO87tG4V
U/LmbqHNBNNFmduml/jpUxTsYzP8Rwb6AiC2HTmMsmhqtp8cWHNl8GPW0QAmkajd
JLysI3R5M3vvM9GXTun9nIgBFiCaYuWV6K5UqjDKpVPldCOEZWJCEJSyYym8M5Cf
hynwg7FKggfVabndLmZ9W+ZRKnGCMRLw/RPMi1gVmgSooUwy4pmOfB5bbJRiuhI7
sk6v29oQ0XCyG7Uifr25eCPEqNtR1CilkVODwDtwzoGiopSjiBKj9RHJl0XnbeCv
bzPbn/wt53CWEVmG2c4ZYdrdIB2eHUjrKOeorxKWpC9ZPmssunuwOyoBJk/97Bd6
MJ2wB49e7b/xoEqDyDDboU5QFiJATHM/MB9CwCgqUpTyVf0POz/xa8jMjoTzb/Ge
emjVzE+Ar48chOlvS+japR+X56EILrAwwsIjOaTSxMAjUdNrqggUGUjjdek41pva
tPGVyAJfur/H99d9ofKYlAqJl+rtAJi0taUqnr1TKNNyQZU/OpjAJnBpQHPehQGj
04NhjD2QZsBDc7lGvS/FtQIOobw8QzNRBNqqXQr8qBTWoTevTWMCagqhsIKJBpr5
tgAxtTEQiSDFJt9jGE7wWB5Cywy+AOi1nLKIPxWYzUCs60My1Ul7XpEUGbAFwwOJ
Zq8hINm6LHLiK/f1vauQ59dEYBP/2Ill78qyz4LLv3GG4bsaOqk2AWb3uFz3AxNh
GnjdvTl5xN/i/WRecZrmfw9hVG7K6X1SUXVf+B9RvA6CM7zjd1sewE26XwmY/RJS
U29jlQqZq7bzMWgyus1j/V8JcB2GXXDQMX7g8n+SCBH+wDggEY8zqBrNwUx3kBB2
/dKd1gYF1HkKaLD2ESmk9lFaZvwYugE6Uls1NDazv72+gY0kpeBmEFy7TjOMTCBD
dtwNxlqzlVEzzqlpqa41BTG8fc6Slk25CMxqscBg3iMPr/ucyYpFGDMpOUegl3el
GMx3KPsSQI7XgO0zqVdY4waujqhhC2DJFM5SKPxhgeZ8x0DF5YZ9qwUf0akM8Xrp
qMgz/JL0IaMM+Y79m4zzoiPbV6TNj9kx1FA1o5Oh+hF8hn8Y8VbntEaWMFiLlmYy
tHSEZ97Fv8R83GX5pUviW6uGyUmJreDl4do11n/910Y3hGZ6Nu4RzlL7AvE95oBD
tCGnW8Ir8xAXMpy72jqDNLX0TPSib4wCDk4EdMvxGMj8xmHxnUPou/x9d4/77aze
tzH8gtXFgS314HF3UDYImazpu6et5UHjansVTX97MGHfEUJItS/pJierqbWMBZwj
f1LrIBmpwxkgF55saWuvZjh1h810RqoazW6Y4aBMVB1ptCQTzNBJrPpZrBgOVqA5
07YGzpBbnd23h7gbfrqBZUj4Z+bNE26g4I3nOsGYpLKV8CTY11o9KcPmsmYg3V52
2i5ETjhLymWPejzXzYFom1DR8mfiPgXOLcUJdKbUn0abJOnRo3fvYUKzRVazvcOl
MDIkNflGzToNLasVoqQ8AGdYjNnUCHz8RdlHJ5q/Bunzgf7JOZXvCba46nv+P11W
DD8f9yO3DW1XVZCdaoOAaOXJQqPGS4nEBLsmZ9Hc6nAwK3A4PC58SGP0rpFRNIo4
05YQTU2uvBZVDGCGEHM30/Kc12nFRipK5ElPTY9bzbOaty1KeoNox4olad5sc09C
EWqGHospdMW7ykBEk/105REibTKzgn5Rl+sTeRSQuz8Bb78pjJdGWDpRhmhLyAyS
Z0A4bK+3OLrIWKOhjN5BRTgzdApG7DicQZ7nfSPP/fAw8P1QQXGNWzhmcqmMwUB/
iroStCpmUluK6bmXPO68kQxlv0nMwrAo1izUDD/cFZnalP7JryalyQ3CAhV9kQBj
hzcNBnjbiABFEHNKZzGQHTYzEl72OFwYmjkjvzxVoQQUXU5Xtx1yq5jjNbL+VdID
gg5UEEq6lFaClupGdAFMh85MLBucqAR/KdfiHnNyfpomcUPqZ2Sn/3j2Fcv7TY9C
TWeJ9qou4HS5wW9nOnT+BHvRWmf8MtZfLh4W60AVlvoP5WYOXyoycZXTABXmhCIv
+fBtRo0v/6FfUDmpdE5IY1kZsrnBl8UV9xIPC9gyuS65Hm2reOCpMDleEoX5soO2
xbzXoyDloC1h9QBeYwLaZi4SivQrdDYQtiBYdzgwK8joM4yR45Tty3ntFOlzuTjE
J/J5R1DHojCp8tuv3cLojWtZH3CFH4K3ec2lzqR8RkmlFtvJMFHtfyW3KdltzlRQ
V65861LRY4Z3z8aMSIaLxv+pSNSZ12eBBJ5OuNzkSwXJOTq8Fy3wZOAAzx+EMq3j
NXEJ71Qk9mQFOq2C/S5NKxhUe1U85ndUNwl+ppvJmdRsCnfO/TaxI2cPVD/2raS0
Da46T4sHFZHR4wXSmmQ/5nyu/K4qQE8T3jyiEndow74yw4iPKsfEwez+brQ6Be4u
VpVV+2mEyyh/k7u1HH0+gVRSocuUfHpBzm0BKGz+friSaL4M7NwhOmVssH+Ok4DX
RRg1o3g+Faoa0zawsVxNoKcuPw8BgauVvCP0QM4atVmD+K7ohkP9u3e/I8jT4jYU
PQ2yBgqhZWJVVZBbPHuasAhpuYbUAhEKew45e8gItCn5fWYHDO0JKc11x/Cyt4k/
QuvBUUs6c+ixpXhC5OGRk+tM/W8ok72shi0jgraKA5/PN7A1Oi8mo1qfgeDIswyb
fSvvS95R98maCtsl0BHpLYhkcQrkYpIeesLj7IB8Y/Ay2Ji4HCdHrLadbFHlk7zp
CS3TvSaoXoM0EdAqykDglztiPPYiJAqEItrkM4Mz5u8M1x16FbYCsvm/gTZWIZuZ
tiXMFIRR+wh3f62ALI8vyqnYku5BaqvTCKlz4umqjMLS9J7z9jmWPwOC7uTQEBMo
1m8QCDgm/01i+xxCcpS/ifTA/J5M1rWDzP395gvC3QZeMkAJycgMcOadn2sWkJjX
6Zd0by5x1H0U6cwcDSi9Pr0Lna9oQkRFrTD+DB86mMxkssD93l0cOqPAjmcTsyGJ
LdnFnFubDIR/s28NYS4+LVrVNIh/VcT+7ZAjxFP4J3zWsBffhOt+8fxYRY274yIh
3hjESETOzEAyAOrcnmHDg0l2evDHRZ/zrxLTh7NZo6+to8YGO4g5ZtZG22S6VVr9
kVG7cnZfo1/gjCnDI0KTNXyiTyQzwWZz3JzfQT4wxHqj/w4eTRuB1uuTD/u2UkMy
kV9q5Y/+e/DT/JZwt7+98fe4A5F9Iu5EnKBtLpXZsWxdSrzce3wu/jdkk4kaiN6f
cF7aIr4CXbHKf6tDulmn8qczLXXPl4cOev28vnW584701BPq8a4rwT26cdBqhYR5
nxgTlDzRoDlqFzakpVBsKV2ogPVtviZjSl17p/Wf2XXxBc0qvH8nhmHZgF1q03WE
1xGJAlDKFR2ugd99dhU8i7uJKgZIgzld4NXaAA2s1uc/Q7hYwi72TGEc4ekn5tUh
4Z9xhsn2MgBfZNUJuDYR1TMJZzo4cB68ZHThvf+wi2DyeyyEtKCPINYyVlNWXXL4
JBMQD+Um1MfbvP/WPSI+m/XzJjt8nUYk8VNJWgAlaJaDjg5D4f0+v0dSBN/3Jl4e
tYUUgnmHhqMHIfs27dkfha6/NrKgoYQlnpWI7pY+sw9eQLEPPeTEiH2BbQQ04qjh
NbgzpnRhLAvvaxBuL6hM8EKFkGrliyM8XH13LgOsYE+7mmiREGOjPAI29RmzwIas
YBV4kS1rIt8pfyC6tFaIUjZRCa2MBXxadFuv9JykfHKqpddDXZGJOGfSdi/9tf3S
5JKumNNz6/4BQlQYkU1cGhWNEP8vSS5gF0lepF5gvz5NMPe7GUdiHs+XInVxEo7/
VW+Q/ae3LvAoq/WCKbQu1iP4261TZO6I19o1KToVf/pRn/xRt7ELdNlWukxjvbqt
+G6Vi87dxKZ8Gi6aq7ojzTIr8zV/KOxD9zSEUCrGJfVL8OO64w4oLoZqfTJuVcy6
ep8JnF1VpO87xXsfNOr+elnAOQCnKE24nEaizLpwmclDF/IXjkwjzxM5ELmuFrJn
kpSpO9BQbqi8SfBC99ijdlTn/JWaVVgkP1Y0yn5zYKUo0fYMYeFeEr/al6FByO3U
LMFToVulybfu61ON3JImSntuALZIu7E8pos4i5Aa5IriGinizx9WiJ4Ia0FO0oxn
IA8+uCFD+EyirsPtd8tM4D4DD1nzMTIrxE9dKwb3m6tKK7cu8Y0Z1GVSzR9OSzSI
EkbqfVzEfyUyvP2gh0gInk0MkyHwe2JghlWZ11Gl0qEjonEyMeZdtPX4ICfk6OGY
JL308rwdymxs6q6vf7jLZ2/RGKxhYdqlq1iJr+uKtB0K9sGOMmWtVdZZCLlZ/FEg
T/Dwdvxqxg5T+DuoJ8aLIxLzNtBB8bK/hjTMGS94/YCcYqnAnHog/17k2Dyn+1aI
VFQVXhHsf+YCEKI8FPDFsUw5B9jTmHmQ43h3fF+ELhZmdRCbrzNflo9SmIU8pZbn
s585ANVFAehpoKK/Rzl7A7oi4gQf5BSf7BUwBX/me7mbL08TvbT5wjNlKP3FZ3No
O0t3tYwMX46vO/w1YnpOrk4FlHnVCwauhDRmPK64QFNYw+fzUvlQ4CCMKQ07xYE9
bIe54CGNIhwZR41XgP7c1LnNwNpOub8DM4Oi2N/Omj8A6GWfxZbhB/o9hOPd8x6j
OmoRi9LieD9aYNBOPbzV61dOWSPsZ3Se1niGQzt//6fAreTO8BPCe8dTqgB/8x3R
TjQsfyGbpEuWbPRZFCMm2Sf6g98vxLRRXU8vE0d84W+fMApXMBZkv15SlfG8yxEf
+/CWCbZrILUbY4ZPhjBH8COEWy11G1th7urCQRaaY7tM7HOQTzTQF/C8XsZUy5wD
m3BzawZQsaDn2KDu9tJ0PT771IWzdSIEzv1o1Pyx2QLaAvWzhDbQxEK1y6xf5qCl
eJy4/posX8W+017ZVgQMmYz1zs/c3uUzqFiSCJqca7lvfaAigJx7R4Fx/C/oMSzL
gNJyp0wXoiqkusqK0ABJEG0BoRT8F6H2N6+d+2+LdhGc9782pA3LXri2g3Bzh1oX
7GB8Ikt2WjOfvcavmMQuM6EuTwsC1r7eTmLOEex0q+4CY8a91AcfP9Rm8i4VU4Bm
2eV/MKtQ4U34j7gf1q0FisMegPqCWIFcAeWQofGruyqABUICpvvwLfkmSHQ028W3
inOrnsQQJuw5vilZ+OVx7AOaNxKbbdmLb8PRGQ1fXvbfx6p0bV7II8DSHSz9gJdZ
vDGzuAaWPUoBZx4vneh6kATdXHxFen0PJxFAFFHHIUx/0VbtUCEjfLKWj9HpvMod
IkNhiCqQJ/ATPFJM2fkGXlFaz3wUHfQGCl+6olIHz9z/hGVfMU3XFX4ugvZAoptA
0rSYhjsl2Dm/pdarXI0vd7lTSwbUcsyBqdA9CF0YT/EEHGsdDTRGBR07F6ILTo6/
9Oqwknndc4Y7M7Zw/BhSliHOFph+t7Nv+1y9qu5sBaZQuOfIfqQGRExe48tTDlRs
nNsSLJyZaur6b3/K7FZLWKrBJpdSOCSzgoU+LRBw3ASwe3+SSiVr6w8JGL4Mxysm
imcdyjQxP5LjevKZXaAXLaD1EEhf19Oaw2kFxajc03FZIVoIiVYNFNuKy2rUIJ+9
rvDxqZXQvm17zC9NY5rehM1TH6PyHwWG871UgYioC5Pj3t58u02SupaxET57+6VY
/PnZvhTOA7ajJq80LT2ZH57naQ0paNxk8CIDq4l6/fIl1iE7gHJOuZ4HXQA3/yMS
VLbWW4XEzu39WbGvT5ew0wjBsqWBMT+z7/tzGt6ubwOLUtB9I8cPB6kCaTbE6Zom
q+06QrprFP+FyvY2vIGNgW1gfzgtrxBmYwQpLWWC2SGaOtAJYQtuULvISsAgeK4l
U/5LzCmpSpisx4xml0J7Z+YepN+1ql/0cv8fYGRPdvlnGr0jnK78Belu0/MzprVJ
P4Ejm2onVrlQYnR3DIydtWlDP5izDSkncTLpSD8IRST3/BPxeUwTmedWnhtGABep
f1hMxQ7ghBJJdZWua8krwV3FVkYlPKc8I3lAi0C49Gh+PZ9V5KfmC8VXag8yoUA/
NDYQsJbx51Z5PvUUYSLAKlmhFGG1+g2WHGbu7qJnpnRiowrLSiXsfAPgvkAny1R2
CUDzkQNl+zKTUg70JDCP7xCEdQ85meyAAFtwMNLeYYwfIdxrysCIv5aq8LKgBt5J
QVLinT0PyHqZuzFZAyURcHuZq/TleYvZ1ETX57f47sYd9iUeNq4jq7mZSNlUsLiV
/Ru8dyN3IfQtK1xaeG+xk2VHLOX45Av3XSpxn81O+n5daYQotYdnH4iokQRc/JXd
VoNxMlR3gE87eNjWZYzgYZ0Wz+DclsM79YwIcbHvERUsiDXpRr1eQdhPMkps6sTk
cBsVl/ZapVqLAQEX/6AlyXU3aC6RfPzGpJdY2oY1VYaOU2o8nGxzJL1bQel25xHh
nNiu6QKBrMp8PTeALNVmnqRleN0oKQ36IynvWTtSGZmAOqJ8nRF59yuRSP0G+RKq
j+Rh+vU26Y5eBLBZwLAsS3wKeFRAuLa7JI7UpSQqVOdPaS9FJ5ZurwA5yapEfOo9
p4/DHO0QjvIHtbxu4rlr8c2QTdq9JKegR1/2KW+h8UyABj3EZkhnvJyeFymdMqJL
OZEr+2g2Ng5qmWCPf1UEvPw92tiY2hoBzCjcycumfrzpPdA7i/3AO5N1EhzrZdWT
TJmiLw1RtoEv3Trpp5+X1AsoystVxs160WRGN5VHZacfNt+LTDe2yVesxBlU+4vh
blNItNVoO2zPv2WyRS/p+JZ62QievzQBw3v8BoKVBGNF4NhJvFAp7h8whU4lT3nH
LsYTeeY5PobT8ElW29n1LxKhUwlv5H3jUaUytHqr6NJYi0R53aOpAgPvZH9/9CWq
NC+dJeq1fx9hvIX64rZmkCr/Z6mnSYHGBoXG5F9tsYOYkdpVLg9xBXg+B3yxVEek
K9Zrwz9OB2hdLuFkhREPy6FnYnQDrdAHbaa8Gg91w22I+4tH3/9PfdxancOq7iTJ
iMZEI4mJHNLglEMiHKLbz/iW7DhZ3gdljg8QkcV7yaiHLWRpWTtel8vecVp5uVLI
JGQY4DYkWrFu/ZLo/mZxL2GoevBBlygoNFORff+AdjSMcJOH2y0mpnLCivi30aJy
iFpoh0Uv8BC8KG6wzL3VqqaHQ7ewXtsKcUXBDKdu5nsKE1fiTi469qY0BF/vkBXQ
vrmibVrGqrEUgpqbLhZDz8CTYfbKmiTlzj4ofZUq2K1s1Rg1HYKOZbh4qOBTzCZ0
Fug2kW6H9wHT6FM1GNpiTSqq7Vz5hJ299+FdrgNKLCn+lL3t9QB8+P604Yi1JU1h
6plkmOw/boeTFHdM42nmUct4oRmDZB5XVn0cI8UdeQWGhLr21ZGqQvlhz2sAgFzP
eP24GWx86mGLYZGzRdV2l9kriSvOEtNJpZo1g/Yn33POh5bljFMvmtaNRni3UurJ
sB56gBkFEksvq4G9FagpVilCDT0S/7J6QZTm3PL7lIP+hoNWCOWLD2Xd9oa7zrVw
sLUnqQmQ94g3uJb2peT1eiVjPljbbkR5WgDhlKxXS50Lbih+TiQZleiTcKzbDAQq
+FPvOwgpjhdtZO+SUSpZHz0GmBRFWev5Brldr/MGrIxv/5J9+ENF8/dkoe88ODcw
WzT/9rxkq9JZiz/LE4Z147PuXNgixg6O6uUYFi0FCx84UauA8LgdYeQs7oTBscnn
bzNHnrXM4CFE9Pgcf+n/lOTHUH9cBZS/iWH3EMZWbxpWITh6yC27b6cUp8uWIBdm
XSKdDwCHGOz2viYNdXveYkUdJIidAkLiHsPeY7OoTW1Y+tfl6yFdZJAJNSQl4U/b
xaRSabOab+mn94R6gctk7EmomiwrXlervO9gFz7fcMjB08ea+toN2ACH+NHJRt/f
iLPv8O7NLr8e6FqY2gSd7V5/0bNbQtyZ4/urupjtvvm+3MZd4Q1AlpcZ8OPakGGd
1oNPCYA+5lGfvccao5Ua4MoKwOPii12Eu+/Ctg9hfWTklPF696+XEXkpMcqzWDU2
Jq0k+L5vJ494v5eEh0aleglY8Kn8BT2PZHQ6VovCj9pQeN+eMx7B/iPe4n1MLyVG
0a65wnAjk7fHOf8eNUvQktXMfxWkQnVrhex6xIpC6nzkIjCxCy+XvzgTWN3JfZ3K
lxqBT+M+xjGGcG1JpazBvRuLZDdiA/iobPQ/hlWlDPJZrUOvJTx6yZn6+89ogbrx
7hEpOtvBo0rpDi4t+igX+AwGVhtcTYtb16DBr5rthKCgap9xMHRKOfv7zYLyUb6S
JSXjdAkOm63Hl9ut+enx9l98ZwbkhQB8yXBUStjQWSm2+V8Dz62Kq9rHBG8DIFvz
5hClxyrTXpUY8irkAqzhPVa0kBGqa1fENcwHk1JAaNCTekqDp9l4U8MOVoo+zXtf
XLHtcKbnq1QUmbmYz+/cMK2fINEA+0AStAz7Nu2wmhMYb1yYDYZ+QmWIxifobRuk
ODb87lJH1U5rnAkMs+mFPrzgqYxBts//7cDQmB3DuWTAzEoJwygKTWphPrVPvsCi
xI/poq1xzWQWVPJW8xeqmfWMlorsTVdyOpL3GiZZAAtkUm7g8vbqttcMychPMukR
PqeWXghPrP242vbYD5Wu6KyCIxVGpseDdF4ey0KofrgGRMQ734pU0pULwIFr6KbN
Tw4scZxcxx8qEjb4yn3G9Ch+eIbO7E6+CfmC3JWc2cRdwHCwdlJ+GPRV+kuEFNnB
rN1m2ZuOmaWONvBQoenWuLuebVi144oCCczy+Sv33PWUJ2fdJk9TTgS/XXI+wL3P
vLW3ZoXsGnbPYWqEWTzemg7Xzni2fRQSYb9Vo1WI7ZP3g1bcZycwTWX1MCkGI84A
zlm6RjMOSnoPsAoZgWZ8FUcgFIsR2SlnY2E8vByEse+YfD9pnbGd6Qxq4+3Tn2dx
IS723BuPW0iTg+Xer0uRt515dneLK2rGw7m9nibrvdrzBhcADETzufezZJgOKxjM
chcFVuBZIts8D37rIWkryRG6L0hlxd28ud0igDTJihS9Xi2AfLoxkjscn9XSY0+o
PvZ1ibrds91lSTZ2OumAXoULCYW+NT3Z0IniXWL6GNZNlEQoef8/5nSHgsHopNT0
ac+cpDVinSYjU1QLV9j2RQsX0lla/44TkwvkJOWimyQ2epcYs8mnSRZVpZkAEcMx
GGSS7/8Fp32OFDeREodcHw/8DUJgR40ghdfDYjKJbxszR9dExRHp4yqmFUu0P+Yv
lpB4IXCA/n8+fMAZFj/um8pLDBBxdXY3tX9ZsUGrQ0VdeoEOJdpcRZKrAokrtdwn
OfxEML6p9SIz26ngXzwAX74IdTIeosDr8skZR2CVgKGKwTrD64MIwPgFkGkmvkiW
JJWHe8rdtA99mtH4xy6iMrvoLgCvYFR/Amjnb/7SM7IaQMloDB1B8v/tbCkVrMKJ
26RbQ9QYVdwPtk3uy50PVyCw30XZXKO+b7+7xpPY5pxCG105Sa+Pud4PwPhuwP15
8C0mfcZbzDct390WNa/wNBc2YAYDV8jSmT5vTVX1Hdib5dD2qpB1a+997hlVpF5s
Zp0V74nLrPL8UwMFTSHEm1JpMjmXmgTL0r6uCpSIZO5bhdqzvIo6I8Gvb7ve0RPl
PwCxXlX7l/QAZWwqFCYeqIILULzLeZ2784ZRpF/Q/J4WOJ82ojbDRD5B9oWL3WZ9
I88W1Q9Srfqlu4pW4Dc87tMB4DQ5Laz0CxTozMsSFAZOsQn2FUidcblYS3sLthIU
smiRALiO2/irfif87dmDHghORe0r0HHBWIW6DN6/VXNDLPFcfCNgGtoxXScydb86
VomgI2GPUQGXl94DWLmpnNogyCowNZCa0izb8VBbvDICilvVdAMaMwTRX5BQUXDt
ZVFfPCpHH15nDuHPKstQuL1EV3DIAftHGRjOfmlCUlGYs5z6+8JznvaI+bDNoWPU
6rbMLG+hsrtnVVQzm5cs2+1/JCc5aQhBzViA/ICBrK96etY9yn2A2+kL9jEu0+48
xJtfe28UoWMvnPt4GaCTJN/2ZGQvGlF/fy95Wa3BsZUcnLRAp2Owwd/3LvsWSY4l
LfV6V2wBpSBZyhOiCwtw5s3VndN5KTCDWzSiXo+vsnmmlcix4WmPSE6djBlT4lDj
pBBfV573iU2iReAJXHtUjPoTCdlBCdcveBRyCaOCTjTNcwUVAvbrIufe3x4tDY77
zhn3r0qWJI4DemudsylzlU5sqV/gl9bQxuT3M/ci+kr6BigjWmXITjHd06kux/xv
8R/10Gzmox+50Vd+2Qg399P+qu84+5TB6Fy1DVTQ8E+JxHLAIrdgzWelN6QZ5jFO
iGb8VWVTom6gMufw0oVi3FYyxgMXlciEkJxKyX6Fk/u0vE/Dtgu4CdXOdkx/SX9I
T3qeHc57M53+HrtKk8tWvBFujQyvSbQFgQDgOFp2aCHdYetrLwT04j0d6e6qwdYm
Iyg1eiMnMK2+DtIZRSULugVmel938L1z58yfrATcotG0wOpttoPBuBbfgjNaHWxu
80jZxsPpXcExFlOXp/+lnG9FMviaKzFzQayGz2yLAQKXenFX2IWPth//Y1zl9Zn8
PCdCVKE+To6djAxAMtqTAUFrkvgx9qV75CgcnclzblsTEteoFVGTENjhbf1wfHOw
3hG1OG9o3glXe+0y53ot+6hImTIhYd8DdXmKnSLGqaVfa4pyhxQMkPy7O+D4DIc+
JW3J9kit79aoJxAekqnoKUcPZ2iXpJNMx3h5pfk6Wv50X7TyGOWdef/OsHWQILkr
aOs/hw0bmoteJy1Bt84uNrzLJ6109pBU+k3AiIK7/nON7GcgoGwldYsNVqvi52sD
P1Xp358RZRc1dPfkeQYoYAfi18bK9IAXhNNnOiYMuE4fZEcwqxYCrwKwDq7c4CDo
IMAIsQDZSCr/8Ei8Gbrxewhp4gclAk9OQ3D3pjmxviu38M5b2EHxFXQcXeTgJ7wA
Qwc/W7EVoKfhNLEyeaijdosHdGq2j6FbyNfj5FIMEnhLjjS7Kta6sfRq+J2duLOB
Quu+oEIf0a1c7YW7J/wadcY2nVeSN1jk1zK6pq51rG/oIHxld4fTN/IvfKtB2J0x
vnkik3Q9G6CxkEElugK2F51zPKcDQBQ8e0RpDNkRnLZcE2GCBIgUH0pFkBgK1h+Q
CmDUpWY2ubPVVGXPi5iQsllB1gD1b36NuzjtMpF+LuaI9gyBXko/IrcL+mYSga2B
h5LKhnARn1OWB6bKKVi/Bf1FpAp/2itMESrtZ8pGzFOOkZK3ANKacN2fpJYjNvAW
evAP40bcEHDRGpeK8cggkOpP6Ao5aVe1vdjwYDC7youRoCwxTN1wM37BYEQFvhF6
NCA/2i79QnLdhYk4guuEj+478VJdY29q9Cmnw+rrOrU6vwOek9IGcVcbM0KsYuJ7
G5pWU1m+V+l5E2WetyLZHyFHOUvjmXNKrotCMjAPs8Pvl5os5km+V0vPfZDBuynC
j5OU+rp6hgkMDzRzZ+SqkB+unBeBWIC0lWa0TGR9BiQ4EHuU+AUT7Ug0+UxVjz75
WMm65wjw/PnR5lTGgBtH3UuQxuHmnDylMRZWNpdDrPX9/4FG2gsLEja7fnWfLFz0
M0XCaYYSljrTXEB2E7GDyriyDO9Kj2QTjlHf03Q8gI/PRvfvKa0NvrWeRiFNU2qm
4FCEJsUGtbtcU3Qhl7zIsKW2HalFLh9V1vB09dKuzX1AQm5Mv8NETED8He7ffu7d
gENH2tKxDZLb5tuaQ7iHuWqaqb3cCONlRWcKgKcV6YPIRqYBGz98Jw9mX8/Qciq+
OSPFMmJXtvyCHBoG+gQKdL18iaXzyjT/5xmwrArPUV/Y64Ed0ibghJ94w8wqa9JM
cr9V7o4WMvWZIMi7ZWEU9x/ZethPZJiQM4VZAlqwNdW5NUd2xivPhl8j2Xei2HO/
9M6ne9WhiIC3WAjrLt5EZ3MOo90PB2cYr9QsRWlvf91I2Q8+RwJ4F3Q6ed++ar8K
LFQk28jHZKFcZIv3oojyLPfVc+V6Qb2Bb3i4EKjmV6cV863O2cGSqeyD2ovjn27n
EwJl77wwp3VHPh7yz7zQQP4o4sVejRN/nbWWQh2bfrsBj6dqo2U7gzVvB7Apip6B
wHOXQwf025BGZEy+5sN6NosalYgPqt7DBPqFPa3hhSm5sCGfEuD0nHyNVAi5jiE7
xvjCiJ0qO2zARk3BWabWrKxtUNoiAtO22FxFxMP68b2VkQ4TSQAEyMXUVUS5JkyA
ywjDThRO/d/ve6SQF4wmdvDwavUtDRWIIM8OGvSrilY7Qk554cf2pptMXYnlSHML
xTXntXC6ieBOqt7Z07ZRiEQ3fQtVjTyx1eyHH/z3DjhAJouuujbTzqLIDhTXHdLM
gk5ERpOBLYKByS5gDmtDSGDsG0PHZyGkUIrj1joBqwkPa7YEYdI7hyqoAQnkTR+L
XTkd2UNsEUoCNXya6TczXjlxlsPmWw9VtEnHWv9SUiDjvpPclfz7V891nT5DxUIY
JIbXLqZ7zETg1lvVIdI/kiLjHweU2VtWPZpLN1sAmiDn2gAfS2ZqqOrCEEGujSbQ
sbP5kqNqS9OheYapm7Py5GmdLhRSguAcwqWg0JuwwPUcDLACAGuvMzLtWV68AGRa
C3mLIaUm+NVs8oFPlVXvMqeUAf+QTHAwlPyDwXuzxO4xqIBNPmIlCOc7yoZDSMAH
oouefL+z6AHT/68lkmXMKEXu3wab0toTau9ew/+Ovq04CO6CuS5tsWI03D7+yk1C
wPTAh0JxtMFKjW0LGF5n6iFsoscD2FSouoS1cI+f96xLnNrvIiFN96FqFVF7Qc/c
JFlIeX9dpCGi9+UMDSivCmbb9fcLg4erc2gsjU4TUBOT73KtGgyndDkJFCg3RFE+
quO2TsYAPaQlj0Bz5701yHgbwfTN7yPd2zmtGMsxqb3YgrQ5psKKRZzErVi1bdpZ
Ay/gdn4yzpyT0k12CY2w7fWpVZ4QBIfV/XP1Qx4qkUk4icfmOyrvlgfDLGFIeWou
lW890+KiwjXWGeydBRcSDG4wSWE/HzJTXSjTouK/fBJdKuR025LoEmfWElIZ8V3i
OM4dTYHgk3H9MPUyShlopWeC6S9vxYpR1spEsK1w858OMYxrV+T3UUR64DPuK7ph
BMuPKBHT2fonR60Pf30Vyd6sTQkUPdpvPk/rHj7WWBn7WPiegFrsgk3Zn/B9/nKF
WSyASOEj/OkM2mdMVR2UN6yBRs+LQ2CMu8SAVNxe9YsIb6/GbOVTrCXKM4ONpY39
nZL+dN5WNIJXPF6030XP1b5UOT5tuTT1IjHQOx5dOZlDRQ8F+oLLF2REfPghSYb3
5gowPp20EU689qTbFIetWwAdH5CuucHbxwvtt6BIlo3y5BeN7MPXXLsM0AhNpfJe
3/RhotXYJwMfVx8dhTblCqWYKWQVv1edmN9N4YJwRF6R5yT0PwtZ6FpxYIuaTnD5
AGzV3E8Ysg/1FtEq0+0gryZyzJN6JI76KpkD2usJi2UlISve/EZ2YS8/mekORD1y
eAc5e47/qPlEW+5uSwRz3BxhKRsi+IKZ3PX9H1MK7FhjT5urHSMVk0iBa2Pdg6JC
XxMBAtKXkJFOohmEAUIifnezmxMu01ABJV5Iq9DFLEbI/kGsE35E8adDV5H6Msim
NjCgAbWmaFYkDiUqQ00EqNtGHOyI0btkx+gh/CJ6N9d4ehm+/6v+5mSpn1fxPNaQ
UgitR68W3egDY9JrRPzTprxtDQjZ7BhzTuOhxlLgEAc45hXE/P8Jc18XlQqwtwRv
YYDS7EGMldNAHxbQ91o5ONGX4lxkMukvUyEkNsFXAhOG/Lbp2qJ4rsXitWiHxUAn
kuYTTNCIXKe0LTW11Y3+/xpPx/J9WQglng/MC+r8d0YLAZalaQ/rcs3eaOkU5BTA
/SdPuTPYOJk+lnKY473qmLhf8AXj5KujlEuKVwqjpBkfHSzCv/+VXAXc5oYmyJUe
Rm45cTlLw4uZoLOSwZl38qaA5ThXNazDBAgNUrYRwYpP94vAJmnIAqZeIodPeQr8
EItYFBzhLhuAsQx1W1Z54SCrHX4p9aHmZydywAes4WxOwSvXuu7ORWZZTVncLdT6
8TM0AndWFvDMmJDF5QN0VNt2s5WlYK2YkBc+YqSwhTCZ3iiwPI/p0+2hIZZSPKgX
wjVK1LTzvji4E9ySH6pHitFxbXBOZhH9I5g94hg6c5sY1iF4RarZlup8VnfTnkcj
0tz0YmybWA6kxapQLoEvhvk6/Qwotvkxgdz49foFarivGhy6BcOkAEe/AAuWisFF
xR0zKkrzIHTHCXOn4u9riITXRKXAYdYM2ewyx7ZHpIKTLRL/C1n8U0BLq4htIhy8
61g43owfNVeLCUQD1Wlzvgh8L1F8bxCqcSIW998H7CEoBrKNgYEjdE8nO+wJr5Xm
XgZRzZ1Yhxt2aYDpCUphK0ULFvyxDD+itnV/1gqNpCo8sS5BHweoTNhOkeLJmwj4
5+c/xYd3ICSk1UNkTeOxabVh2UeLSF5ssBo+SxHzVbGnGbnbo/xHmbsB68aDNBuN
6ll2dzAojIvLImQ+Xoqj0g27VGameHRYBPoVt3B9gg3AHf6b7g4+tf5lV+R7lMEP
2EuiW3uN/IxiNUYVVtauGwqobXQV/AW5seu4U1kB1wVld741Gekpq/MkuRBnmgqf
tqJANyywCfLl6noXI+9x1hl65eMiSicJ8udoknXbphj7Oom1ZvLVHb/GbqosnQIE
ZZ7ABay4R1FW5Y0tVhxZ3ASsSCaZ5BAA8FUuUyNc0gU2O1nRpbf8uvJRwrgz08gx
O1tlM/3XLYRKUjT0SizqPmBTZ9Zj9BfYlsLRUa+rllpyeDWqruHoRmXCQDYJCHMD
ZEMrZFYULtYjKbor6i3O9MMPJ+2NCDG8V59l9TICOHgt0+c0t5KIafSDrmIFqtHW
ZcxMT0hoYy81QnFxs6idGh6gbb36kzsKNskVSccYAf6GzVgnO88htK4uUEhC2mc6
WG9SDxNUOh0UvWb41wjA3/kVxb+U+OtMCxS2GeQu/eNEQCpT2AW/W7HmPEaZSv7e
MngBeD2tMSpBFeDlYMN7oduHohnai6DGFDv7AycqmLq27wyntl2qAw9qkfpL0CML
lKCxxVEgoPUe/WHuPnUXQ1RCVp/kEH89+aWNRUWyIwygqF6Qmb4gZ+2WgDO6YLre
fRcWGJH1MVvqKjZFYS4FkHlRv1h9t8tjOz6QGgx6qOe+Q64u9aGtwPF+oQqicqsR
Rp1UzTcA5rtgbFtJW6rqKsUMGImfqBxroard+nJiVIU+s1Erk0FBFT27FW12ANa6
L43VUSBP6nKSxX93TWQkFerLcKBZ7rQI/3p0h8NUK+bpgDIiupSSd30WKsGVd273
Y/dxMUd7T4X/otJswf0RztK7chE6SVka5fFnw6y7YtqxZo+5sIJNGK/1PuVDb6Tp
5cUDIDVCcmbmdDix0tkG9orP2GtAXLrxWdAjXDEF7uS9EIIZ2+E/EGI7PeOZnqok
8GBBl9zxHzucZ9MpO2bzP0ybuoZBpmoIOkmgV9s3i8WOf1pQ9STPmR51xM6rwvr5
2LgtVI5acGBLbpN/J9fHjzBeY52DVSdtekWi2p+33k5AMtzQNIAKG+GoJ9JKY5ea
Vgn11VQBmlYTlNJvuDQ4XRk42Gfmqy+9kEEvT25Va9VJqA+27xhCG1hGOuHr/mud
kMpFCCtqzCYCJfUqZ4mGVNs0/hD3doCQL/1CmWFa3OlqN6A/MJrAB7ERS3HsG0ED
l70BYl+ciNNNwRMRYODT3o7zff7EytGdt21XTIJ0LCQTquy5Uvt06ZREN36Wjgql
rZsYEFGfTaHL80an45tWx39lNhEhQbufiYfq4Y/EcnoLlEcZ4ffHqvUI/uCqvBHq
zfoW1Ro8WMgYSMap06B6B7/v0o4wg1XpHwGj7mMYIiBRa/WKwbu7iW1cBSJ0XUWN
M2E3nXnmVhSt/wMWyKj9ZnYwWkaflF/OOoD7hTDFfoaxiQMHoi9Wgk+QnLofi3t7
gQhOGB5Dl/JSs4F8HijJXBghL2fQ2wFf2cXKyYj0CX569g926rqrfyVo3MylYLpc
BPCjBT1UXPZndrR45/Udq3qlAnwTstiaNSt0h58pslXWjyV1yPW+Fh6YlmGVmlgP
BkZf+g46+TWIqXD3GGB9+xAFxu8MZXWoklj9us01GYLqZ4R9HQ4KxIKieLOGEZwU
pxyVe+YAA+3RjzWfao7ea/jYw2rZhf3J/pCDIhrwTF5Wpx0TlcMCqAabg/TlM045
8oAM7PT6fvXPyv/h4iaM//4JagUNVnfMq5lxYPbLu6M5ZjhOYR0oPlTGBRBSNY0A
gzHSjOyh1tbdDhsZ4l62/JGUyEV+coDve0EGNci7iZD856ftRVaxWwigGIvEkUz7
Y8wd5fdd3Fw8RetDrv+Gd42RHnaFyIS1Zs3yAThCgn3o0N6kQgYMQ5nQGdWOZ0I/
vpI9httThSwkTaRjoOQ4Js3bmIXUUYuo6SHbWL0JxprNNdlZdFpSBNqp8fO8p6jY
R5knkwK7WkW0SCDxSHXtKMM5OTjgduMDRK0L1/VSQKLsYWs7bBSRtRtHuyKn8+1R
HoBbO+It77xTmHIBoh80ZGDZ55qkWeIewYdXkW8p6Mmxt1y5ry1J88RsOx//XeUN
AT/phPW8q/+nt9dZAp2C2Dq/ddQF1J1tfy0I018As34Ddc6zCrGA2wP54LbBLqUG
zf30jPmm/cXnjGjNplZPHOTBDjUBZxvI3sRzH/ZiAEHZDu2fet9la0qI/fMhxlat
5qZzjv3PziLznlR0Gzu3cJi+1sdQQyNtNXmtK+E9wfWDXIFkUkjTWZTK7bxoDo+s
1riGa/1VYwLQACBqMzbnZ2ZvVR29Q3aFM763wlFqfSqoJ5RPRsrhyTTkBowsfV6H
dVrXzWmpeVX2vRqQscOff2ZPef3ghJLR5YgHFZ9WmkQobvEUumssOWr6X9B7IYqQ
a8fZRvLtpVRZqteqi6mI1qGjrMXJSwC8EI5ZLEDhnACcmIvwaUBpDctU63wJUoDR
3107re/IE9Tkff880DzwOBLRR5pWRb5VI0PqGG1pQqLvcE0P7SoiLviSl9UDdzcE
L+yvovFF/2d4os5Q+W4aAhXCC/eLyymIVZkQx1zhtPNUiQ1iw2+Oq2gFkYAoWM8z
WjaEoV5DIHH8Dn6dNSiL2grwg2PNYqFtXYlqkOHFlytCCYmEcGGHgiYefgfsODB1
1owsdv1ob/c05asBgz8PPFHDlyn19V4Aet/GiIaCoFBS5foTnxwTeQ89bFzTdXzQ
EoloxXK1G6UtvLS8n02UV72fmq2/Q12wfSRTHuqgA26nvtyl3nPuY903wrGpUVno
aRjL5O1FH5sBPlazStO3Ev5mDmW1JK7LV53tkbRqkrd7dHYygTOpNjveo8W6yMeC
YAROG7pw7B7gW97J7uo7elcyDumqrQR63wgyjPmTo//iwImV54RKI4qW7k7WTatE
fqQV7wRQD+y6o1ySZ1BR/vNFFrWPOjDGEG3XvlTfgYzgXmXKnCSkgtRMNIQHIZvR
7bGOj33wDT2mncNlv0LLLs5oSUlMGkxIhZiWFKfKjBUrf/OSyyfiojxad5m484W6
Pog3Ko1o0QthtSxsBvZ+XkYSww69AYAjkHpEK0mRRXkL2vd7PcQf0A1ziXmbHjCV
pFa+ul8lsRz1GF+v6UbNCAq3kBajqjIkNa4RqU8Yrdg4a+ZwTIasxMdKp7NNDKOI
TZdPf1oIGZLmiEsBUGQR3/4lWgohv1NigQM/rz7Svb4B8EATiors85udKGuXXPX1
uwcK7c5BQWjcrfqt8jzpJA9C4mCeGuFkM26GTUg0WboM68PmBbaOieF7DcgNTxn0
RKZce74NjuNkticNcxVBxWh5RTwJAN4m7dfUYJsWNwO5dLhW4Lox3nOzLuS2Es6w
2a/g/hsXZ1WgTSl5PsgAwcb03MUWgt88uPay+CGyscRcmaCoWfD6cVxufowkLUtx
17VcPOTtlq/4v1dFuxn+S49a4MceQBuzpgQVduVu0hoGyAqNq5Bv+rpT6E9AZbvB
ln27rdtH61aJBeAD9yJsI/CDP8trxJU7y/4msLW6tDoosaPXxxidTXksHU2aSMow
keFbG2JZLmEiKknANGlwcdkUZvNrzks0jD5xTygzG1HaVMGhMh/LoJNEYNjakLui
d1JiQJ0NLgLn1gfxhiwTCRpUo2g9RaBq9jC+n2+a+pTRNQM/Iaae0ZS84nNS8Idy
3XY4POUpQbKy9E4T7XI3tyCAfLqju3YjbCEIB13VThRK8ozr7DZlZE00KSbCXKAj
+V5JA9FnssGLsbXs5Vd0x/dtamIkKOM20RUi0C0O959B3SSDRwrIFK415CfToCvK
Kn1G1gXqr57ER21wK0nfRvyyamszBkM0qbnGdq9Ul46w8uDEjFa/42w0/VHq7kUz
VWsXNloO1QHlnCmSCfZO6BRQi+UaHV26Okq/AUb5Pb+Ta0X5NU1NFQVObLxiDrFB
EVMVavTf8Gt89MNbS+GI4hOfq5IjRC4DptzgixFyL97HlgHJbH/kbblnOoRf5CBB
OGF45UvZ0SyHMYWz3MYWe6a7jBZh+7BIWFvpztiTLTPoWNKX08nWMRVLu4T9znCE
RSXcNxitsPltJTwiW4FrV4OWJUCw+7533GYbaM1y6J+O2rr8NlHV6Yp1axgnlXPD
/4f4Vbc0SznbUM8Bk7kCRnEIy7+R4gxv7GBEm8SGwCDoJk+zlAbmDeXFyBUb02u3
GDFenJxezjJnXvl7CzwV48ho9OulSia3YqHoker3G6QcIiHy3/cAgnbaL3LNskys
2ezVokBnnghgS5gvvC8C8kkcuQfEdmxy9pdJ9RNgoN/LV014I7Nq/JRj4sDbzO/I
BKWbbzL4+WPdjbxZxODviyTKsKMrDuaDQ1rza2F/JEhIitcSAgaqfAQZ/HK3M1GR
Kso+e66y06f9yd+kInc6JZ1M99PRnhBD0uIrLY0nY4HYSuovFfLcV/3BlIY7l11O
vkChd/Ca13ljcsYl6RWI5ymfWTQrNIjAo6sdn8jaAyXkGj3/EXAKxxNG3oaT8WW7
vOnB/misLmSFmrF5r1r1FnM3MFH+HO5SeI8xI8DJoj7QXXv2gO//liNF5hmtM0Pt
1boQdsG961XeFriPG7a1zOFKNmfpxaMIR3iS95dUwafJVmNKYzeNve5japAPTS5x
cFKJUyMvIy382k/+WELPoIqJLPPWkvrwTmJChji1HAip0a0afHn6AOP/Rv2Szq8f
2v1tDaZzhRugecH3IdHl3dp3VJI/H7mRssh608jm3Sc1jx9PtdyJk3kWerr+OoHS
7Tcb3XHrryfwu18jb3wXXwLeU/5SWciUbp5ak1YwAM3u+1IgsXwNVmfzYVtSAu55
hIB7b4W+rs0Ju30NVTHjdhYQMpCJAAVJ4NVkotIvHxPLJ7aGkI3IfztDVGa6SuZT
xQ9qfKkldYAEhY5COk+2PQiXBf+aeP92OtVzizMghrFG7kxECsQ+4i1UK3K8XRtm
48VJJEPUgBYpQNUDF74F/zbL9E5tTqX3CgiPH36a/2G0aD4i5L44rGFxzX1Z9q2B
jhF/La8OuiBQ+Z7eDEqqVHLyXyV3GcdB7mOEvBlS29oi9EVkTDRpsGiqFSJvVBCN
VN/NuM4KAzDLBgDawsVk6btKvmWYMuip1ehoqpTJ8ZZb1Elic5CSZTCeIbS8Urqe
G74WZ+3oK0dd27QL2fSRJqv3RaU8swaJO8iERT2RzkFQoFpaStwdPEG6RYRyhZw2
mizQ2K3OkJvMeSOj23z0224hk11hUOWxVn/T4OCaL6qIbGoMBu00kbqL0CXHpDbt
/Us8SNmXnNI28fOw42rsDLWl2aG6Ss4+zoMlVaqkLqGZ1PIRsmPH2QsaOY1vLIBx
jcLwipTYYMjoIinECTrVjDdPbD6gpJCAzR4j8VzedRwAHZgZKySLmkrAg+guysUl
I2P3+3cHZ6WO+tRYjqE8eS5BiuHoVbAzFYcMih3HQ8TAinIRGSQK34jnoit2u8mi
tNZzq0s8eodAYFQc+LCsI7mO6KgiT/8jIT/z+hNsMYDUAD8QiF/Dj21vG7+jJ79s
NS/PnfTl4JuM9Ho5DqLTsnYU7r6NPrxQlGKihEe3zavXOc0BtiypGZuhKhbdxo0I
IUttYPOeufgdZvRjjnc7S5Nuij9HUytq8Rs2i8D+hwRgHxv9XXWo0GNctbU7cqdt
M3Diy+dfurRyMGEsf2eVoe5C2KXPrWQnXULRt68IZviNOqSL8UOTHOD0NxR/V5F4
QlPOERkW7zvJquGLEXxYApvoKURcr7V/H7uDxHVQn1swYo2ffxDDM0brfhzOYCOL
PdPwLPaJpZ3bHsi9sVdZfclDb9KZGCzVJGyR46NrnUwRx3plhsYdMSw6XW4XDrhh
BuE6pwJFLQp6zc24h+GJzuEdoeXVBra7Kd99wKmk4+fwJhSeqsR2C1Ld1EeJp+n0
ok/IZOs+mTw4U57fVNlg6ZfSpo9KVeuQS/PuOYvGpKFeJG+rmq6n1Ux8Xrf4fPYK
2Iri2fnKtt2wnQaKk/B31NBkZJa2JzvrBQNYNw6mYfZzlrPsbezqd592mPhle3+H
tXqmR+IoGfkN4S6GTsdYjzcyly/rN09t8A4dxkehkkM/LyH80c3BELXYUPYdRltm
0BNtzDlkl6LrGsrl0Cwzy0gBNhZLbfBzwXZqr1ZVejfTQrte8TETqSfhsz/EyII0
RYugJ0qq39XrDM03aIYU9m4DebYkeYvk+wIyETCbFw1+0h1QIXhgJn8DE4P2doVf
C0O0uOsAY/GkOattYIxBsUfwWslzb1SuRihJHA49LIjXJzAa0XGEX6V5PE/8SQLI
ssAMgUv1aNaMg2CSIBu4Bvdn96NZa2bXOHzIDATVSqyImIWuT7Um9aoY+IRWN+uu
dF1Hr8BURoFtIxuHkICIoyl0Dh7TvQgFO9HxmL2NIl21QazX2KC/Pqqmvu+lOmjl
7AgFTjMUuKCsM04lRq5qL0fYmOpohSGaneFnCE0iDnDclTU5t/eRxPkUTsKl/CQT
huO1bGdSR3HbptNaep9VmIBnpQTMZqU1u/lqTbs8N8/+n6sY1DKGLU2CHDu3bPyd
weA3W/9Wqct00bc4noZrna/rm7mhP6N6QE4/dCKb8Hbr6Ar4RWldafagcitCtuT/
YXRIJKbyZfj4MY8COME9bWhG1jVZN4It2kPq1KtLK0bjo8sC+QDZpc3wYTOtVZJx
Egvvj1f5P8PPLf0SQ5xAheFzEry4h+LOTz44skC/Huhp9y0VXJLQM62nv0453pW0
mvsO22e5rxR0awQhAm5y0AjI4XAntP6bh4PhDODfXKp33ZsXuJZILXZIgwCrRT+f
ldQs1TSZY4BTiBjet6kNyn2pXqRzKtnDFIVyqcgxTj0y80X7iB5MtCddlNjfzd9E
Jt/fk59ZwUFDyp+20BqPn8Os9rkIPob0ahE08zDOb689Q2uHhWDu7zPJF3u2w6Xv
AqZHUucWTLqJz28muwVukn+ZN5PgadU51zRxZAxBB3O5FX6nAHH+JOP8naO4yd3w
dx00jswVNLKwh1zvDHIZLA3d+n4dEp6vy+Q5BrTv2cyJDJymxWBeepshOcEmiIOW
rHINdHH6Pa4tQ7CJOGIqOhYQb23e6iAtBidq83fywywPfUOOxhPtbhMz8UcsJzmF
KnjOTbQqbDj+aDWGL7wZLB+yDJaZY0ersKkcrSMfBEgetAqFheL8oQbhoWdnbYQn
UWI3bftbKbHCN+v4UBFtCShpTIckSGJ0Bwejj/gKD05NnxnDUBJ6LFokhcPtEm10
hJH6z47masH9OWOZsxvqIxEIWzv3e4r2ER9R8ddDKJIYcFrKKISL5TUK9TTpnVBF
kdegG/v0GYb7HnAIHKb3qtS9Rac+ny38cgvYQqMqTdMvy977Qo66+d3uFhaog3tL
PcGSN48yd3yf0yd9WpBvCMjVkYNr8m6B0ohMddn4SjhS3OqkTKMbgLf+abs80+J/
7Ztz9jFtFIep+NH9XmYZHYMpbopDU8f0+0UHJ/yAeGuY4HD3qqj6naU8nWGsQrQb
wk/43cLQXcQENvGuelJrvYh0Eo7H4ZUODwrFvBZCoZ5X3bOvXsCcSlnDJnsy/Kpu
vNTnenp9KKBa8p7s/nvQSNduqPny9Lkaon8+tV+Jp2a9DoHAmqvQJL6U8CYagg2U
095GHmLCLJi3HIrFmzAJJ9Wj6DAa54202CMQ/0BvAJXCb9VRfp+Vk1DUu55K+nhM
NuLCbvb5XJ52Dg5/9n7VC030rK/G9f3q/J7FoJ6C8l18BmCklpmuH3bmAG700Wm8
QRZDiOJkg/nCVXSxzA+kFR0Vfpr9aGT+kiy4/MWxsJDhw9WqpwoJ0vLvn86FZsAk
AwYThYvt0zyZAiWuTK+vZKj9zNPd2fL1/O43u3aK+5a6Pwwq069pXnlyWwHYr2OP
9V6OOzq5Aez1t54zhMNSGBrT0vugAn9F2m3zgIOo5iuu07IuadWQjFTuN1wskUpq
TKjXSm+Ysj4WDx6uaox6bGY5Tj+rhy7r51cRPzoHGVrp5vMhgRjmJ6wYsqlKXJGj
SZegeJvKGibWf7u+P58kb6RngUWnMptiNRTDkynWwYfHk/3yB1XCoDcNcZ1UXJ41
aKGQBJ4sf1Mx+KIEjp7AY3pk0x127gxCM6a/7npwfY2Icyvi35lQt8QmhZfcK/Wt
UeDZlRGhKjNw0jZRtdVWYD0T7kbVN/kHCH6GqQESigJgntcQ9T6TSMuYqQnEek7/
6laWbc6rrdFXR7N3MgKUmNCSlFI5NDyAFvsjIVPQAYSyoowVKsy5K91zkVuWhpzW
TyKHs43mVHZGeqOobd6mC2M7oBpTSYX9JkkGp4qVdC+nm40xtNVIHZQ2E+wl6vFh
SBYgf1pvfAM1LVctsVbMSFpjuMpbztLs6xfPAcCtO/BrNapymuvBtwzfyxph4NaO
S6JDYLhBXflpdvBVTRI0hze8Orz+EAVR3biGx03+JvdXEFvlihkw1cBl6kkWrzsO
tHMyD0c44s/jvrZM84M/cFZAVjyMUW6DhRlq43Vd+c5bcWDbJjewnhpds1eB6I34
uyD8RBwidRQ1b9DKagRd9vSb6seydPE2pCCR2Eh0NuEECUF89VpWgV6VJwQqtdwl
68+mv8MBZhf7iRgQ1Tuly6DZQYwqjrdlc11f8n9peVZSYztwx0wMXL7hssokiFR7
Y3IduZWmFiSAF1s/1PELD5uc4B4tUyhjoo87fhWXVxiJznxFys+EKGfdkblLaRXR
xg6B6bAPWXbJ3X43b9LuHy6x1qymkz3oiXLearNlemC0bKw+FD2OsXe/IJriwfZj
FSscsZKnTc96KYKw2WWBv15ptsM54t6Blu9jHyTG4kT1YiDdODx8961AXV0uYsAO
qUC60bI5burOthhImzzEo0voo67J9mzhWxUbsjU3ssK10BQYXoPbeCFOFrNIXT7w
3eaPg2paSZ7tcv2JspOnOXhbMDJmGmth2P66PJcqJdcAs6SrUWFvBpIQktWAvnJg
U8cgGwsvrJMSVieISFuh5BEe/08FVhuROg0u+EFS9sPJ1ZSaNO+QwAhYiJxhffvJ
Qlutqz7I3xxvVpggSeTFijimw2MT+5UW0RzowxESd7QLVfPuUX12F6DsYLIhVsZa
az/4CiQtDpmfjSDqwA5iULhwSQyEaQ+9kKQELwKcHi8D0QdKEVo6zM5Hd8kV9y2m
aLmjIEKSmiNX1esUzXg0cuj2Mvoy+ErnU1CNxroKxPSHJG/NTmAEv87E7sQNSacC
G49N/KEdhtteBY8H6/mkR1QJgP721EYCE0LvKbXVzs0VnOZAPbMRFxCrYAw4zuQx
UZ8VO0Ieb3ing1Z6rmshd3FI4sUqXULQD2qYDjkHnGRNQKARLYtaXH8Kj5tb4ZdO
8kWWsygnyHd4ieXnY8bslKFVxcu28/E0NgG7M4lyjVT52bq4edvP970Wyd78ppOv
/ZtaH7QSHNXUmIe4Z+6wLbB4yoAo6jgnJS1W6mGnLRITltfnH+r9juZ4D4QIfyrZ
V1y3IWOsYfbqUBwwGD8IlMCZldtIn2aiz4EdRxZlGSmfoOZwkjzrVbVc7IwEGz/b
KzIHlpSPD/2V1nIVzoC71Tz62HzVTSt5qN73Cgvo/t15Kv+zxyB2pdFCyv1P2Uek
ggufyy3rJdV+/6NG50vhrg8rqOpWWV6oUen2vFOzTJwsgxQVqwuDkfAMYOD/mPEf
xrnaqJBRaXrFi+kg6yJk9PryWh4/Brxg5BsrftKPenQCpNjuImaHnwORo/cAQYCW
hWrgIxUZjJ0D3f/iD9ArpuIplLNV9RUjQROl7Wt2FA+S3VjKE30ZA4wdHar0NBht
fjlsHHOQKgrgPnpNdG59dYKdED3BN4X7RiWoFk+AWAXunWA7WQNGwKts09Q5ccAN
zG6VeT2dmi+TXlC9UadkFh7F3DKzB9bFuOeJcgFkLWuUw8UAchrOZtUJL2ZKtOGm
vOgv6ppaaP7JRulTj/l2piLiJ9xARf986dmP5N3UHOf6RZyLlsFjG6vcDh0ymyGg
sGvEn7VrxlOQKa8h/LDEs9OxGJBKhX9Ib17pkv/9/uO22br8Ug3vXiLhfHpPom1P
0+cPtDuaUPlL7d6ciaGppXrVxY27AMphzdjigPzE7gEn5XpsPxeNue40X7fviMTM
9MSmTsmUTRhAW2VHNbz1UevN1PXIufQeVwxbZsUDxRKD+iFLlQ4P+chBZLGVM+yz
c0qgRNOZbH1sQF6jfoWU/oe43khltSktvS1brkH/rL+Rt1g7EAZ0/3LH5fS7IMw2
b5wN+Achzjngi7hXfCbPsAi4wzM8MmXt0YSyVm1j0FtQgBN0JY8UIrUkrQwQTeIv
esQt5XPFJ9T2F7q3J7oDmU9Q48uShsrlymoX8oyCfFdvvrAvJFaeMuiX15WwCZ3N
puX1J78buoXxxPQmbJe1ajDfSh2u3q9WcTAK05BstXG8RSHRnn5XF6Wq+LdLWDuS
r5tV45TGwEhKh27KU5NnY3xYxWiAVa9MTcle5J5n3WgUrNipzZlg894RamvCKqUM
J+gks+dXg+qWCgk29SpyNKK/9KjO5gC6mmx7MiTnFqCUdRBshcsnPnQPtzuV+PVQ
NEeKsajGQFaWEwSDWJfPxqa+MkXpdqUtMSTVDvotjPQatTfZKYvw3wYHXVvSkam9
k/LM85dc220x/Edq0ACY0mjyeI6Avr8/C12wU8E0i4UY6TI5FcD2/pPul+59Dt+n
lq2rTUKSLvWvVhaXl9w7eUD8JJuTnsWUQJaYYycC9rp/6z3b9PJOifFtGJQ9ivVt
GrjfVsYryjsfzAP/d4b+toKuxx0Ea9KHVObbzsVTWjxZ8U2VcfZk8WnX82ANeju6
PVP4565xuLO+SYxIhwSP+hDJEsCjxBNQsdaHL37ve9sji3xqZTzO4M6DHzDtsd6E
FAltm0PT6f0FhXCZoayD1ya7N+3iC0DbF7Y+w8mvx4D5ATKfaftSJFWolJAyIL+J
YyefDPX+Qx2kTKG86TrFv1KIPfX7HX10oE5EUassEOjKbgfd6GHKaYQL1Dx6tSsN
l9V/LwIWjIoktJFcRMroobMH68Vb092LMmGA2L3bBxpF8UK8N/DLzKzPDwKbtXAm
bcUrw7/CSP7HJyVP4owrwAzSMqR23TN9T3GtzTOfk07IMl+Qsn6LjL0qszeLkO2G
bE/lZhQqM51GgUrbNSPbPi1Jy/o+HZ2t0vvUjyyxIfb7L2kRafxA4fdnDxXUVsEi
tjUa8XzNLoHqLO3dEkmi4k4x258EfErI0FRLgw+GPkTl9PAzDAptAuCCQobfJ65h
ckQphelWi3b4kGxXMaHNw9PWC40572/089oYnskz5jfgV20oQis/N8efMGC49STJ
g2x4RE8kOYMp6KIZ2m7IKmfpR2ptuUOSvbiPGJe+oGVpFTmjvY6x0+giEtg8ZP/j
+P6SGLUxC3q/UH+CnOxL2qel5xFdTw6pXfEkQzfk1k3fne9zTEkrOr07fAxGeiHR
qeUfOAcBjWc2gn6MWRE4cRHg7scWBXNm+vmkFmGPGS2CDvPq4oQNk2Hnf26VSo4+
7eXJshwBJSt4qO7/r59CbqW6xVyaWM9YjSyHzpo5MOzGHgG0bJ4WJQUOmKDGuwbR
zT20mEcTA4J8hhPnDbtGEYycM+YsfXRG+m4N+R2ne5P4QPUY3drwpLZCRUtGWVMF
Td6VpKsd//XFA556b9GNhl+tFAKQuo5YbwxdQUL5e4xGjTjdQK8NPH4z4EXRL1PL
S6Z+YswZM9Nl92eI+6CqL1Gh8KTTQinDam4d7+kI6L2jzqOB0whcFRrvWC+LyfRU
uNu0CP9qjZAgNn7LpEItsL8nCgT4pacdal98Y5vsTYgLcrdyandLChoKOc/YVceC
s1WhH/193EI6sDIin+LHdMHfqzw1lDZ/fI35WqouIl+yCBnfN9A+21Og3ZT402M4
WZcIj1hmSIF36ra23//WbVZSRQ5lWvMTU+FFlRzUVE75TACpR+gP2yfWORDF7L+p
yUPMOyp/Do4wHt1SxLpBHT3kSLpaK0PpCItNdH5mqo0uAhpxwQx5dLaM6r6EqYfN
AWcQZwE/JS1WW8tdUNzMmbsWUzUTc+AFCrDq+gG4xWFfd3WrOo5jwIggjeTHzz0p
0TGpteZs6NIfr/HFH9hoI7MbMYf6OoNxRFvNtZotfsUso/ApF8oGIOqlJp7qM43M
BDJgsMQU8MqrnhgOOpHZNHCOhGQJdLwTmjaoOQ/44DVhDU1ONoZRLH86rV6t7BGR
re/lYc0RdVwEjto9Sc9lsY0ZglHQz65AbQQqSCBj2+peKSRj1gunnicS7o1XEQId
fn8CfHz3EADUpeLuMwWHrh59QVOlef0HS6AhIvghHvZzr6TWiV4Dqpc8Q+DGP3rA
CGO4nEQgyx0vrtJ/vY/y9yKkXRf/26NezHqRywokUHciJcIFP5X3z5WxbMbS8nPR
vw0IzupUMqra6lCCEEGgyChI84u08uQHShA1mGceaV8wEpCJpBgpsEqsRWZkHzh4
Yt3nfzo/qSgACr/WplZtWDl74VQOmLys7boAVR2OmLaEPFUx2g1/PQf97QpZ6826
37DCJbNCMIv6QXXevI4+lRETLCyA8wzWM2ri0C2sNSB3nnqKHuDmfkQOc8LPgl1Z
OftCecoe35UuBdN0QbqjG/iSykcLpFninKjvcvIAk2CdPYj6xFrkt++scivHLDps
CIHYqOhaz3+NtdbtAuMgIqUW33UvG1RxaMQ3xYWRQ0JqAc+s5zfkW6eCJOOJ6nFW
SOEBY1VvjZUr1Jam3CbiPeaWGD7a8U091mczPv67mDETiyYjwMLpzCOMvJYbR46j
1g4/UcUmVgzO+32y39k2sQHsB0johlXrVJaX5uQNOCMsHA7uYatYX9OLXLtgp9AY
6Ij47VK1l/o+OQY/zTMkxAaj4zJMLAL+DDSYFTfWwwPV9cYGqZVEUIorEY813q5z
h30CZ5fjAWBw8GFbtSfIXWmapoTacwIH16RjDn2z9UDH5ofsbYXK37m+kaZoLcZ4
xX5d3nd3z+uzZ4RUeTXPU7b2YlA3tma4pYx6Wn5imYTNnYnwc5x6uKJ6pdv9fFpY
ZnyVJWan1Wg64hHu9MoBEf4TaUWFLpz8hG7B+MG7Ym6MvsFjC7O1cqcObCacOe3i
9lEtYFk7tuRAVK9zWkCBg3y5M334lewfmlwt4AjN/eek+8mzRMcv9vTBbQ7k4DcB
mRuT2KRTXbs49rihY0Gbwe5TD46UUbKWXjIjGBzC/zCukEJZgCmlEkbZpiHSjHTa
tNznTnSveyIk6NhM4dCbO9YJwC/0tQaGY6VdGruOAfti7lbcrqoeU24HQvOAz6/9
0gr+YTdrQ8fojDsJAZhXpJQJZlDO0o5g3r8fPi4skOEwMPbvowNSmiQUWuDUZKEH
vUvyyP+wPYW13lCT3qG1iWWHuzwgPjii7Hw4hKRfZn6yKTThbA7R0zHo84/bl0EU
J+JWW0l0UijPok/Btt0VdJM4YzkQhTZ5X9pPn2ZHXfQfLZ3LZVTdtuQ0nfO30FJu
c81YPNC5C+MD/eHdR41qocXslliJbY0BNFlPJPCskRQanZtJhIUcstC9fLSvn9q3
ikRqsH13XrcGVbhiFIpzj5+Pry+xVce2ydw+5Ix95C2Pf/lgvIgcxRqLhcupC1/W
sKjO2mmSGqczn/VpB89bWC9/tHUS2vC2VcEkRgt51eyd9CBLFdXlZjKhdDrjbTDV
drvQnJMsYG/ubFc8oaAJZvVi9Szst8Ouhed05iGdQg+Lt5vhrUNX1nFSWzBVVTXx
DpbUN1v6WHABZDdP7s0w3iNPGPhk5tItgKGsOvlyQZCoubF4THKGvS7ByNkIver4
dekvdyo0pRR/fQh9qdcpWYELz2az+pmRBGg4bAv+7iTBsV33HyTGmJT5fg1lbATh
rZeqBu/8VuTYsLYtr1324P8RcpZUbWWLgwYGflHPRZ9rnBG8vuAshpWODZg3tC/m
HBIR8B310G2AKVCueopO1af/J91knWbJxRiCPk/Jcg3yoR8EE4dO6sLQZCA5hRA7
nUX3HNbtTkIlmcCNeFcan71QAqqJ2zuzSuqxtyLlevUBu1gmSUi+IBLsA13LmbNn
LY0vZ2EXJ9xeUl9a8SJXkNBQxc/amyeNEIypT8aCkjfga+UIktemKdvBOMX2r6nl
/AFE8PZ6HDt/vEPCEXtV0DAnjbMKJULT/dSxFD1eRuA6lbXRavqLvyKuulibmmYx
78Mq8RAFdPZ5+B/vmpSOjlIIvZDM/djermetGUbaxCEzFeSp9Aao2YuItOK9tTNZ
K3Gw+aMnQQNLWyGfbIL1OX3I1ig13Iwouy5VRZshlrn+EM7TrS0ru44DFqpe8WO1
UyjOJ/vWiVV/HiDqFC/3k0LghG8FWJr0xu7cTJmGpW1JEylDqEUf95rvi4n4oa5k
10vXcahV8fh3lUm9v/qNqCobEG8lLrKf16cbodSo3pnpAOfRaU1ToLXz/C6v4wvg
HzVkBGueWjtR1G8iyfxva5MXsdJ4fmOa62DW1OVCa2l/tyIGNWjLdciLLoK36r8A
D7mcYfy0+KzHqCwf7//RbhvB4RVszM7mHUNcO5Wxk1FFrRUu77+1Pb9FDN9A7LD8
Dg6e4aAjFb6BzXcDpepoNmXDtbSu8Rq522xPs67isr56ouz3tnNuhy1Z/n4V80kE
r23yqMGUpCdTyW4+Lene7Ohzacfamy0F951uYy06nZYxpoMnh1LUfh2i2n2HDM3M
LhTYBGza3ez97Sm/nbH4890yApXO4tPixgBXwi63yeWWadUA/TXplVkqDnAtfW1o
06RjBWC94lds5NqJjYQvGnTH7O0DdrgVD+H2Ds+AkFxhrF+NjsUf2B97iYGHZ7NZ
2aDWiIwa5IY4MvcHsWbLveoS/PHH+GrEqFd4K08pdobih6QAw6OpP+VM/TFAVrXJ
ll/dqqHnloYbk9pD2TtzqQbVleAXcOUEFCtjy+y+8ddZSlQ5JRaRastC7n3rsyyP
4x3tZJvfhOWofThv41YfmX/cqQDbxxNMFD/M3fmb19AkxexZyVngXdpUzDu8tBzW
mjWC+IbFvZUeZYRSeSpemV0TxWltMqLqI7UPlBKQ+L2dIgbBmQ1Q/SM1PlfzZXMg
fmYSenDWFCp37m9fLg53avYimXCL78O8LF2oiR1c/NeLQV1YcGkDb2nJN8ozRz6O
CVlzdl3UqHU/Q+emgIT82SQG7Cf/KETUQodfoIcJqaurnyMrRLuHTfcF795WphHy
od7OGvqbP12O0qLbYaUh1JhOvelrH6ydYm8Dq+SbgutU1nInTNLaZzwZx2A5Ft/3
Bz/MzvAFpCL4rDNss24ozbiFy0ddlPliXYzT87O7edgp3gQ/IrLtaiOjDw6SlzKW
8LpeRTIFwR80wFFtazFYsqdaXosCN8MrSS75iBpcS0nSUACH5DryIPcPrlkhWYsl
ORTiqeW8IDRreQeYFydrBbqvtXe6YDlghvyrO55M6seaLYfWhljIqBiU/1TUvj1D
nOanjLmzNfAKpxsBtgkUnKhPG8n1y3nuM7PjtrZMDGJfcvUdCb3mswkrCwp3WHEi
JpGsw+p6XuBjtp5NckI9QZobmHtsKOM+kCZ2pmvBNtZFF9FnNNvrd6kR2OxuGbYt
xa1+pVTmOjEqNdJTbaSRANJZdzeatbb1h21vH9vjavw8fodCMywqSSXc8M6k6Xal
GO64+BYbs5YBnug/GTyOPyLeUr6uONplw63Vx+giAANRLRkQdXA/Jug0p0aLBo85
qVj5+qtIZS1CTiT5skCCRPb3cLI4uvk9knyXxThJrR+o4vCZVU7/WQ76rb0WYjQ2
0GiTgmEe/RVUkG7KnXev9Er3wuajjoV5jPk6XxjDlgHUAgBh9rCdBL+wZrYcIPtn
6Mnn8mzKMXditZSrf/WVLrtUp2lpIGy8U8EDBUJqrzM6lik75AOH80ExjVj/G2+Y
W/qdKQOEjJTWzMlP2kaN6TsWbVQg5tapS+OMCK1w9UfEFcSVma225r3E0DJt4Lx4
Z/G+MzRp1Ux8dMpRlz4K7FvICRmmsL/086hu+GvHi7d/GRkJC9IGMVWFQMB3driF
TUPWHKSEt+4ZYIH19BU0Di8EmOXxxp8me6pzxdMvLDPqWRkmnqedESXifZx/8J0n
/pP8hsvHmixm5JV7jJZ+D/t/eWKZYvugBMAVauHBtUIWPEJCAQT1N+Ls0uvej3gU
BeF374teYKlDRqZ+7ZuZoy6QNJ8URQB2pZhULcYVjZDVJ3/B7eq2c+5GHrqbRuOu
ikClPjYcHBjV0NU6uaJk37l2R4MQSJBJH5ZfXOX/9C6evpN8k4JapOd2+jZm22jW
yqIp3zISg7U1jQXkmd2b6IjzwB7YtIjR4lW2J0inTveyqO/rd08m+mJhByu+pN0U
I4lHkBtgAD9Hol4iQ91QnwEAm+vGU8nxShciKQEoI8TvMWlrnLQ/+lFWJHvH51F4
n5P2GiXfAQ0Gobr3+ojJ0V+C39V1nJCy2sYMKIjGLJhEdRssFqzgN3XPdv7sv4kP
TF/y8Z/AiYKf7/rgh5dML2hxx8D9MUE8yPjMasv/+vuzLkYc7xI39/s9fovM1lf6
L/eltY2kJTnIzGFlhmh3gH5SdvDes6xSLjoT8iC9ZrXg+YLPy1fViWyusfSUycFT
OnDB6oA3HNrH8rpZGBCcFbLrLTgobbMse+j6CwyvpQvVBMuHUcqRJc1HFityqbvB
VMZ79t4Zc9OZohZl10DJzOul7u4a8t8CivbStYdxQxfje0Jt6bjqd1sitkLSId0M
OTbTvvIIM6AxqwRle1aZ328xf+spMjf2LOITzWTmZytOuRAqyeGdjiWsSKW1xjhM
zXPQY09plVEQLfhDJ/NzZGjJyKuSsxrMCTQd0rxTp0PXhNB0S2+NjSQYxH4K94iy
iaMX3za4vwKUxTZTCcHDeZerce+V1n80406jbD+Mo5kCVatRAZxbfDhc7tsELybn
Txmz74MvFTDdZ7swLG/6bDhN17Se9nCt8qaVsXzeL4DMJ98OFgybBeA5RcXN9J4n
BTER7da8lFg9Tv2K0Cfs0QDa3RbuG0bCjbDWs/jCSTyQbLK+JMsLrKJG/qEYvLbG
YHUBdcPX5sI82S8AIEYsWHDQKfpRuOg4D9zSyHeVa+a3YshUyzBw6VcdtDzPjh/5
atrvFUNXd9V0XIu7J+HKsuskq0IVaJhioV1gnCU+a2jA/4z+KIwQ4DGYF5Zw51RQ
YhzURD6MY6KrgGMrtPuU5zKoGMCXO9X4nAxYpI7tXcVTXMoDEmWyDYdz5DmRSJdK
hLPW8a5tqTaPSeIbaRhhmuLua/KCvaXCt3G3Kct7Qbnz4NBU2dq+lcuMMTLQPwGy
56bux0Efv35XPeHtMe+efYGR0t67iAY5Cn19/iIXaKZ2Np/62cokOvvmBwB/t9l1
wVBY5MawxCW6lWhyAUFK8Vq+xC2Hrt164hKtrXGCCi4rWSzoA/g25Y1BOwHi4NVz
rILkyi6um44gVE/Tv6FWypX1ZQUpKL/k0BaSA0fdgm/fhBDT4N+hXskJ3EIdxOc/
9LB8jxGAP6Cn6L5qE9hEfWgm0+5ECRhC2uRFoUfxhFYD/fFfZDuMCBWDBS+CgfU/
PCdAHRDBGCsjq3wny7I/Tw+Ginyw10m6Kug8qExaLNpaaINjtKD9WjHAGrT4vuvR
J8bO07qTlwhud8dgBJpIzah3y5Nng5PI66pvo801+WlqyyW0svfsoVPRvgu6X+no
9tbqM1OWlsu3LquqwrIto79uv4gq32mMexBM+oH16Mw+kN0QjYHVz5jQ5YDqHaPZ
QHfZ7H0O300sVzQI9bc3mwDySJPtT191Ycoho1YHAR9k+ZLGdKY/UVQFlhRoIRkI
xeR2awklZ06zYr5fobTL17VLRI8x7Gf1JJLB8PngMnMQbI6620L3Ihh1+rR+YXzd
3aQDETSH7xGLaU8F1jRmplm41c9a5LoRaiuCvaQtGbLX41IstGCngytXcxY9itXk
kY7VqdbRhLsNoztG7XV6U14veua708lO9WllknvGkotk95GhSnOIIJlLa3Cd4QAF
gmkQpMw/EgbmFgMqzhx8jwpUFi/KKtWRDYvnfNpH4vYUFK6CyO8ED2N1CjLQd0D3
XeWXXhfyQ6Rz/DUvWnBKqGSKu5DLneAWwoLAGEduy/9l4wX4S+Jxf6Tr2QZwp7CC
7EcnOpzvUzYIigFZLKJT9mgbNKy9g3OVUa8wIaRA6S7/hubtM4TSRdrlyikAIi4x
Z6RtsKkKxuenHdg5Xj6axuiSbVAu0+Vv9BbTVlweCRFn46EghT43Ar+xw+XK0kkX
lU9Ak4kVIlAf/8fapu4ajEREFIZtYf5h6K+tw3DC9UKyosFZ5Jt4sq92BjCKPFx0
uHKkUd/CBRUyBTOE4k8mFhr6KbAwrp8ovYxOLXEeWHL9HUA5jCema/xmcldIiEYW
qlS4yGDtr8Kyr/kIneSt86e1d2VdwIr3gkJ6RnTgWIRFuRYvtyTLWrcX+Gdvmrfu
VcL3zUDngcJDM7hL5ZSxdC6CwrtGlc/fu40n6d50Ru4VMNFT51OXNimeoxM1tDG6
5aUcbJpILvUoO3BL79Ngg/JKGZHaoxOwkoWWES7ylWNU5p4T3mRYZvECjJKGcoaK
i/KtwlHBjrbZ9tXQXyyOWt6MZeoopjcYa0lQbIEZuKhAmntWFhsMD+2rVhhEbGPv
2I7sK2PwqsCd7msbwEbXm2lLsnDSePq1LLknj30PX0ucdIymJ/n2ZebRgmBvyl/r
pHu7jGsljRCAIHTJDEMQTjNmeJdFlcxRL2LSAmNXmwN2fsOJwj0LCZFAI5DS6Mz/
leXthi0aRRDFi9Mat6dQk8MCAnmy7hQVCR+kFgfwMwf4lWAyTrVBhi2y8r+AoLOC
vh5uVdCP57ByuudcqXAyQBdDl46QY0ugfhgWOR2LSCEZjiM5Xg0eF9xlldQcbHz8
U2Bi1P2oQO9e8W6d+nQTA2CgxuvhzDZmHaLEu1irFeC0SM5kGTWaPcAsJFbegITo
i34Cv1QvQfUmjJKdQOv8dgx7zbBx1QRnaNr2VgCmBccsfTlgtf6ub7MFh63/e56I
19Off2cL1PkHEG2l/SgCDSp+sdhkuBkdCb3dJB0wzwT0NlHfAEaweLSVgkZMvC9T
sAxJICJtmGyXhIxr4E0kkkSzMKTbAtQmCyYkS01PBcvN2w96iAyvtFbDZ6ExCRA3
tTf00HaQV8UFHFgznTdl59NNPnfPx2cPZAR112Fy4k146V4rgo7KBcgMq4tDkWsC
zBZrtlrSEIsTFIgPN2c9AMcdH9cs6iTqQ37BL/4dehwInqt5V4A1tK0NMz/x3Slg
JvqhnzFNYgO2HfNdnzOY/C/kzwNQVWmIz7zLNms5pAO3Psw3QC+3B+1c1CNZwm71
CQuKhTMyCdpTNgbH5PLpSvWSEcw+XiIQ1xUraE9nN1zDV+kf6bbmShUxHMAqUH6r
CihgENyi4Kz3u30WbGF/f5AzD+cmluF5ChedAoImVxu9Zjeta60HtJOViGQAlxju
t9p3E7SIjNIEi2/GQmcuW+zDamQggvHxRV0nmgWHWulXrBL0jqC5CAvL0Sm/QIJ2
TbYTLL9r05ecDFNu9mp05mxFUpiT2PueXL/j3xrkcgBvPXjEjpAqnp9CBSd2TuhH
KrI0cropHghkQeQFbZ/NfOBmv+hAbKrcswt4gzqxYq/GarO2NZQ0hEy3yRERWsvR
wqhwwh+1aOc4X29vutw1KM7ojuPZmJpXuAz1Tl98ot4Qgf3aFGXE65hpOpc7P/Mu
qBdFx6FYI++08AYYh7ra9TmRBKWYsRo5LSvFiGGprU80c0Xx1Sb7SI8/gKUdlbKs
Aatvc2CtwXuDWhiPWkRydZKZ2x3on4b6Ut1uuXz72Kc6BCG7ZDwPGF2X/8s3Z+sk
G7rXms+qnvBw3BVJcsTuBGcesnN/dkQ3E17aAnOP3gHX8vC+jWuNQNJfwp4oF8LF
lgwteGsUfAF8+3jzA7HgNR+DfYMQuoiYCBO/ubfE1pgeXw8/zzbKD7kds0KnZBXJ
S+kvgHrt6H7s8lvvIG5dZPt70Vot+Eq8YC9bNYmgVelYqoIsySLIEpnpv/xtRjvQ
njx75FP+yQ6BtpuxfQoQ9JsX+/15v6E7DSAiE9Y9/+Uw6vBqz2lCikiYFm7M6UT8
7ywVDembTE7PbEOwoKI13gNna3m7cDUw4OIIHlv65HSs4ZbksMMuVb3gctaMmFPV
rw8cBNUFi4yAT8aZC2+2ZUlGZ5y5i7wSOvgSBzPusgla4gdCVTL9DhgJxsgx3RCW
KD/Et20AphxX77y5eYqWkyjpx0lSZHgf3o+o8lI7VJcFbWo43V0mqDAS8/a3Lwmx
ZI9M4g+ak3zhZCiKKykqaMu4kZCMyu6caSHqgfnn8lJOh9WbVdaFfTNLyv9oNyl/
jdnlX8xuOe1T0t4n7PRCq/nQJWXfHX2sz+1pJkyz/THvzoJag/nudxRscTanWL6L
I4ptLJUq6aa+0Nef/JVhGSekdwSoMq8Vr1XmOt6IEzEspeZXfe6ART+YWCF/8PmX
aIK5AUWu7jFjJNd7OLy83MbvkzuV0hI53HNiVS/bcxBUsa/JER1PbPTzYVettEfq
bC12oh8pYMElfMWJkSpVGIhJB6MGReTNv4SJ9sRyQCf6A5ho9ys6Flt9h9KWETHm
UfylNR2j61vhCVCwRXGAFbnV7+dhXfjJSeveutSz4LWYVV2JWosmVaTDX6+OVa51
N6vhnKFOE84JYh/KJPFGzmWFK1e1xC+9Ij7rriaDWUxvoTJMrctanCtHhRT2n7+f
W5XBlsWy2lkvBCSx6l1nhiswV3R7k5ViCqjdjwJMK+IhRXQ6yYUiMCmeaW9b/0JT
yNi8oo51tm2hEGVe0OxRUYQEivhCrFxUlXP0uubwOmRjRUZDzTLjqniU5ONgHeFm
E/j4yr6vJAGwgdNsxv/g0uhXdbgFdEt3vJRvpDuAtdDQTKCRyG+bAEZSrcd0MKUC
rrUMpBQ3/EhW7VT3g1o1/DZibRM19/3wuz+t84SebBGk9hnAhKYSs8GkMbDZr7I9
In4uIXiFGVZIhwmLOhBlDTFCVQEGtyC+74HTM80Epci1k9GVI8XK1xwQw3z248e/
XERzTdfO8PgCzy+Xc8GuZbYup331TAnXOHdaMTD71ky19XtqDHmfqTj/Vi9dUsqs
WqWBOCsAEI4B3SFqVd6Atgj3K4hjOjNkB/wr7ahU65dGOqWQhkd4OkNtYne+u4qG
UW/EOZNgDBXYS3UFvCJUJ5N4PBExxXB5F3ACG5JGxD5zIevgI/IGPcbCYCiiv7Fg
NOysc1ZLdKzsSBw1oCRRf0oYKvG1WSU5UkffkYan4GZs/ImgC1ssHF7vx0/uC6W1
cv1RV/K9vfIpzFLVqwYpHtlQcCE9GAW7u8KOwwFPiHeaHGFwRaFYlbqEyOJgBXe9
IWARD+c9Zuk/FSNlLZ202dLcaYZW7nmS1h5tHXcQET42fazBhecmTKqXzhjBJmWD
BplSbZ/Ne6EsjWII+tSbK7vyWy5kM7t1Corfgpb2c5y9sbU4++QShk3T4g0v6q+p
XPW8ZlMPSDrr5XSsj0rIlh1J6LkDlGzms3Oey+hpI7HRz78SKsv4nji2147qspPZ
OSkY4kGhrPyQZCdNMjP5MAW+Gjvx6yFtow06mwWR+05WgoRSysjCLwYnU8d80cUR
wt4segUKG/YThkJfHJJzqo7so0X8HDYd4BsVUMyPVYRX0L6odLZ+PF3PvOBGaf5j
8vKESO+yYevb9++efgOnDZyrTqmMDSMygq8ef9LCjWat4wsfe8WIHrxO1JPFzif+
Jib3mk7CG/Le5wWZpVU0kO4eajj3B3tbcoiWRU3jwPwnLb3hpAjyBhosNYPF4GHf
v709Vxq52eU1jTxLfNMaTV4NglZXhKMuNoyj9fM39h5LuUtsB5KU+DGF26njlfvU
L/J1KHM/hvV51at3No00cST/wTWg28d7ffMq608lfxYkBdX70AQCpf6wnxML5pBi
naPc4zqlQcUg6sYpkiQqpBZytG4W8a8UsQS3bEJHN3l/E51Fxq6AFUkBYnRYFM0m
/G//xWNR0RIM62tIT4UZfe6xSbWUNxcNm9YYjmojZFnVUiRsm5N0KMOCQ4prjuPP
0Ya1sw7taurpgUoR9bloNEE1vMn/tou/wAk6mL+VcMeVAroUiewTEXneOaeCgRqG
xkBRkqEdXL4+VsAvTKLvN4cJUcakHpXuC+7+FWUK0O0ofb148c7o/2KHuWcSKxHN
8ZdFzToK+CFcsePSGObBjdXN1ty3GbQMkvcKb9Fxg6Oej6Zi/bf3iNB98e04RmOG
sz0uImPtXoanbXNega7E7nEEY2YpbaZWP9kX9fEhImbHB/ava0e+IxFAkW+cSduf
DcfARGkLe1GMh48N23vml0T+nTBlW7HTpXbV+OJ3Tz/0IM9vaSEI/oiz/jGlNLyb
FsABWIkzqjnRqXtGSmoJrTTntt8ntzUMOrnScexzzNyDJQxYSunp31mPvQEjW4YI
A8AnnnWRB0/t8sSHE6dyjNTjOKxUTmiZbcghkIbJ5Iy/b6oQhYet05bEFlKc35QW
fPkP/FWxiTA/y7tmLPq9uF07PQKhe98Rt8TYUyMUQuY2HT4cUVg+mRvv2p1EERDd
nSCJQ3NK+fkWpH+ZSesOaXTTlLhDq7PtgY9sOa55XxEy+cx4TW+owNpCsapG06rR
cuOOy49NZ1RmngW++YDqF/jU6XUICq49yvBlODfFFL2uE4YZlmG8hspjPmrbHq67
2dKE0RoqHQRvjkLD+b/sUVHF48O2twtJ8/e9COlAJHTiYOI5i7zrgwl3RtoOA9ut
Z2Mop9H7Bvzrx6Li4BBAv9a8ILMFBk4ANj6sX+6smJvm7PPe1Gp3L9PtoJPOsX7o
taYt9NjoIxJpRC3Rew8Gs0jQtOPk5sIT6+z9O2VAG82Dd7QPZsqtgzmpiyZF5aOr
LWjf3R1Ab/Mmrd6ObwqKDnLxn3S/GBO8gWLqei5/fQzEbYQArJS7iHocIukTHiuP
ptzOonYIxi4kzgIup+4n0YYvtJYQel7WnooE3H8cK13BFfH0MnAF2DrhxJjsCebw
z8EoOyHvg8IcX3Jxb18nDbYDH0ozzd1wtVm3Ku9prp0iTXIFIISx71uDzy2dJFls
wsoyuWOX891TuCRqU66RhB/dE/217MlO/21jtrJhw6FBiyhdOWoxOAUzqHCWvZmY
kqyYinKwH4aMJJFNn3PXjEy8rHMSz7Wtzdg/Y9cubI+kfWyLEeq7eILzIiqKq5BZ
ird+7dwyaD5FiJIlFFHSKxSizPRj88KG3Spdo4Qm4e73N4MqjBMkc8GYW/6tD4H4
MlyAUhq7Y9hWAhq2qAtnvENn5ZUvB3aKCfCaOmUacsp72sP+w1TG7s7SvTazDZss
6vACQkUQU0/uQUM4F2a4g76WduKu2RAB+SbrA2ZG3eIZuTWPVdTiv1Txi7zbZye+
eRjNCamE19zWo70wQjVPUHG0jO38TlQbCGn3T+N2upEuxFsZBjG8+KFNhb5PVcn/
RyxBW1dZzljUJr+sCIqPRtGU9PP5fl0SK7IoBQxa/lRlGed9Kt06tOj8IyUZgrlZ
K4dn80RaII52SvNbOD9cdlnDHQdODh+PbVBlNWcfvfHIWILQDgYSabUqJykve613
6U/zUISz5RNTxpHwwPAjeggqKZzy5sQ0gHLbLnUFM2P4t/k9n4xoAHPjwYy2zcci
MpH2fBTnsRTYBDM6QeXjTqnJImjW8n+9uQZbA8yFYe3nN3q0OyfotalClgnkBSNE
ICgqjxhg4M3SHK5+dm3fXVH86KF2/nyfooJ64fqnZwDx+mNxI5YtkVDe4MvAgrqN
1Y4l09UA3O5RPRnWwZQFi7OoPLpkwzPRIHwxQc5eZJiAl+wd+aKi0eCN2mqOQ9tA
N5z5nQRh8OkNaq10Gpnsz/PDS9CnfSLiAtqsDhxfV7s+Yc3AtLcpOC9FclL+Va6U
L5b4wrE46+Xi3V090s7tx4gB4dQYgU6n30CQ3fxwJaT/E+7lAmkEmKmTy6ESqG1o
RapY8xoKBiL30OYjMpWZtlYrtQumvlPzq8lRz378X3zXS8ZkmZRWLEqXEl7mfOoG
ScTWQkCBrICe4GpNSaoV4Tj7rgdoxjkuhHxzrwQBZjnRieLPSZhB2vi2GDMXOQ0V
ur6OBJs9httpPViha2Jb6cDNXAeMPzGdMhuoTN68v4r8h2M99HoxXNgg8Ti7nwNH
3ujHFfHbE4ps5F08VJg9EWwRUuw8FWRNyQ3YWPukZe4tWihehS/t0OKHJ6ktLe/O
ujVrZlI8AvKMbeNjv24hvl2JwMIrd6KRqbs5znKzq4tOCtTJEZIosaPXtA0O/uzW
75BwdXNDVwhDeOfJ0TnWT19WsCBV8oK+EFpCEWJvjOy0zG2DlqT0ddK5Qhol5u4R
sXnUGpe0Fv9bb5TGOYhUHdKxYvJnodh5ACnNYyPWn7PmlW1rWDbsOuOI3t5UxG1i
+1h+eKpFa0gd+6gzwPTyiKQ7lCxZvrmtYhI+QEN09UYSgW6K9hEIY6SdEF35PFod
CeN6tgYDTeDHXgXlYnuqYMkT28uroL2IYUB1Fe/dJJ2Rr1CIbr9UmVL74PAe6muo
xxX97O4cK2ECFyGj6Z36n3eiDQ4hv8B9bktRo9XrbmSApyJ4N3+jtYY5lldWE5Va
wJT8yvRHP+lBrU1jdTwXXZWuGKa7EAZVMc3UvR0VmJZaXSV+MivmLO3nX9Uhmy6S
HqZ9bOFHvAY60Gs2uOFeUgB1cOsRT9MlPLQ+AsD6vhlAyVMSHl9eDsgSR337Kei8
zZp3QG0V9iohpsLRkTW6K5So1lsFCLzSPeozl26bj/C10ajvFBlXX7Bg6+uVmIjC
GTP6bFJO8hiBbgPULDX5hRMwrr2ZY8lSTcawBnSWQyGIITmL2fQxPmMUBDvv3v5/
uX+dAyvLgpgwWFJSqrnZ+E3iaZJOF8/8zJPBiCsgyUDtuPF3K9RB2nmQPgvT/Pnj
ZCB8SL77q52o1RGueIxIE4EY1U6uPYtpORO+r/r9PIz5nfVfNlGPYAYKGJDxzGJF
e/P0ZqusW1K+o9vzy27C4fSthh1/QWyq3LgGnvMx6mSKwrTKFvtuYX/Bpo0q5cEj
cpcK1agnJBp8qpWeti63ZiPFZqayVygZClo2csNU87kVobI8AY6nV49JRsYiDnZD
3QgdE33jnSbrvGO8OXDeYH4k8sWbhlxSAhYoG4wLXE+YAavfI2P3UA3mhrgeeNi8
dLK3ee95leiptKvrFrm7lHXwTYxII1x9fhmLt8RN0cumBjYk+1xLX+HmLaEGT1M4
KektNoTQ8tUIIrXvX/Ey5Y2i1/q452H7MJ8oMF5CU/b6aJMbI88uLGDmCkjkjFgd
xR/7SZB/A1veYyKeylX2CTP0MfjFYocAVJJ9UbKd5zpZAtOPd44C5aJ8qRfGzhSe
IIynQipNnZwlEnvYSZsC/3imZ1rB/Qg0tLgkHnHR/+YW3PMm00y6qhrKO1W9juLI
6b3Z5kvQ/Jrz7qQA88YDjwGHQR+LqVAtrdfFUNTaN4qO5H78Yu+zTVJ3iUDSvg4o
S/dr3OhWc6De8z1KNUltV4ZChUqWcKzY9lZoNpS2YsCeASwIKO67AfhtTc6Wvi7Y
MlLKP7HNcFaP1LdcaSZC8CTOYKSXeW4ske97Zp8v19E/dAjXuy2gHCoDpaxJUrl9
RzsoqvL9wMKQhxPFLH+m+DY9rFuiEUVVKNrXwBHXrHWTcHUWE1JqPCfKaXybEfRd
GXllfstTLqVnswb0fXydWWIVtwYQySBplf0GLB9gjaVe07IaMsnGlHIdemP3g7D5
ZaJ3h1KdoWgZvJaSuiXbi9IXef1kOeZSjWmE2AkVE8UI6HvYP1B+af2IuowjZdlu
YOMymJzbtU6xL7S29lerD69weOXl7+Vm0AX33ln2RxdkYd6Pr/TLqMgTB/HSrNps
0eh6LI4Liy2TTPP3RH/v82KhgR19MNC/3zYXdJlXtTku0njCFOCcvci9x6fj3Uzy
kxSw/f6XqGZXs1zIJubeow4fMbNdd6CPSEDXlIeXUA58ceuLFF+kS9V98OVVLle5
ysCqauKoNkjuYnykJVCD6Y4mlHHd64Z1/tl9u8eNLVPHUSk4ISZ0nfsRS8rRVkV3
Rpj7qn5ytM8v460CF3STft+p4RvuUQkZleZqSw02s8zYRkmYPVwEmF1koGSe1V3A
v2xVJtW//gArEF+2Pq8E4xPAv477rNBa8rdKmSUCAysSIY0hzzDDAUKfJmSACAvD
lOeDAfp1ilwUI+xfF/lYitFsvDuecqdecm3ym1bk2moLowIkdriRn6iDJ7bjDljp
AXoEBk/jbnfrmP9xlaiCsCtlcYshBCspkvwlW++hsC7LaNl57T8VYrx6D2Ja7xQs
zelu4Bs69NZsmLDtZjQxbKdA8EAPWlNfWBb/NqmLKWtzs6LSnJeeolYzntcOxJK0
ggHoN7lbQW3etQ1i6qzLrK9L671QuALcwUKb2gT6cc3Y6rAqsOEfkagyD9JNsNea
NPUf0wRHF6tzAGaBq3juixS6pA1Ucwwr46x2q9jyUbZxDNVnK8W5Oq+QhKCJsIja
y5AAHpFKuYgkjYlAWG2rpnJuiM3R9KFTQnmRXLw6niPtipVT66dwxEngJFDfD5kP
TO7l0iDs8UYGX65APsFioFRNuqFx79EVMvprojI8gUIsW6BNCYF9wblW6+4CIx46
TPIQCmzKmIFPoFG3LucA0+vMIAClBUD1daUbPNi9Wo4g9cmOBBd2yUSzS1jdGbaJ
8yJMCBccWI4tIcW8wpJU/4QuJgiWViIFvWrGLoCqnBL7yMMU0ohG9yPM6EaRbr0j
scQ7+92SBs5cI1cNuO+t3dApTUduWyCGCJXrvuoQRt7e7hwZVTn9wsu389A/z8AL
sI9jTvrT6PYAAR5jyhBfjG1saKqYQkW0jKgBKmN1GWrojZ5BxZ+5DPAE+tAf4V9R
qZgx0gBEuBElVVSaaN5PamCwp1SSu4q5oPDzXHzw5H1CiCiIQs8KdRbEfJEb/qpq
FeNUL62zLeB/kz/ocuNLajwTlPdvXiP46UKda+MZ60OaF+rQjYIjB7LQjJkjqceY
Vpuxn4RvPWqS/W1VDc4H0YflIU+KoXoE7LWUq4KISopJyhDTGmLlzO04Nq5i9veO
saop8wfG9gxv8aM3aIWXykvq7w2QYWSWjcKkICGaZTeJtNj5bGynSmvRg1OFMYpe
lvNv85Pbk0dKTufMCVZlgy8ksSo1wKfpsblaDBI/qXDSOiil/SJTxcKsFEJoQKyV
BMGP98eTmBPU4E7pB6gQ8p8MIgo2GE6kKf9L8jSjRINE6wv80q2T6dw6IALIGm+3
fWMJ/w+mKtVxG/LiUQ6zm9vHU+XHMr13XuzElfQZSa+M5DAgUuNrONhVjzLLT7v1
pRMOB2UdaaV4m9h/LuWWlVECmiFQUX6frVhrENJ9NE2Lec4W/ZLpjwpQqhO1woZO
+HPKXrm82VZo4B9jdYzWbXxrC6spM/6/Gyf5r8pXUnwVbTjM5oQOO9E5fY031lT2
dTeMzfbhS0U+3N1nBHPL8zHr6GjQNu7E6yCgXfyk0oCAEynUPtUkH7Ci/s7//Ziu
6cjK1b1e36mloKdh1qhFwNzKMbKhMzxVT9hIeWSLwXlu78TCeNw6PMmGc708T2PW
0mz1WePhGcJmoubhcm/oie9fljZHcAAwu3O/YTkpdKzF596zH5WmeQgZeU+XIrbW
jMDaQGfWsXVclNFi3NZZeaH0kxa5vp0lUBJud68coaElqTBPtdUY3QokchTynR1R
SpCJBZs3KYg/4RUg/6E/+eWrfij3PnzXQT2sjQQnp6CLqgXwvm/qi2WlhNHUfCYG
n5Gu/U9UupVvjNQxdo875haJ8YgVQhNTGU6j8L33Gx1Ztl5OKgveodqxEFKIqMTa
VBkR65Bz11lD1zQ+D4jayevUFqDI8TJEy16yScD4oRmUnxhUqWtEkUpjm/dY+EfJ
KYSfrJ/288rFuV4eM/Ua5vRAH83swrpJcuA83HntolB0cVQVOsrXZYfpC4ohTFYc
IEZQ5livvutoEY8MoypqEZE4v8LrobcGqO+LyLL5//2dJUGDCnxVKME8i0nHQnYs
KMtjOBTXysdKmLy/qglk9WqwUU6DmVHtF7yg0T/0cZuUkwTLCwPVS68l1kFtccX2
7X2izGzYAjWciY+2hS0oS+yuU69yiaiFmOzsb6PXuJ59Gp0P7oMqw6bWPro/bKXF
rFey6tvFQ8ysG1QQvlJQqj12dy5FrZCYWr8DFz96KkvZJ0n/TH5ZvBwP9UjZBcEQ
3TXKb+r9K3POPwiD4/yWYEgNfJaEFDnwlyJqnasGrxeUczH6fCRMjxH7p1gsb0Bt
4tdp+j/LjV34b5h7SYIywcBaiqi3Dts2E1HFYJGXRj0EXq32awGkvGuTkxBDcIFx
KEhRKlhz7UAl2/V89Wk1DvJCb65QCQ1MipvAjb6D+kM3pRmKmcw9km7EVl6yZOBn
Ozx5zAM3+62/Gl+1CXmmUQov74NKVRMjGPuWoDpdWdDARUltXw04u5S6zyQL4HlG
5KA0JeNowKeLvh0IQU7Fg4lD2R1RnuVxrGatkvYwE4VNPc8BKT5fGmuZ2Ytn/bBY
it9NgmrPHrQfSkB1IXjd2b2EOtV/eE6CO4Iy6dUC25vquq3O04FLKgVy9Qsmrt1a
R05GDk03lMgGaEJMcjMaWuZvdKug/qZM5bS2CRnJ83U0J+tuZecHcHq4ebqtDNLP
+JYt0r4c1/CIJunF5F212KEocn4Vmg0VoGLq+DGvne2Iz56oXanOWBbC2qF4I9NN
VHsyiffu+HA7Gkn2US6F388a/lomgzTEzODko/C1f8f+wh9paYIKixtOq9T7K1th
OWjvKMnxtTlTlLplfGvZXGjbnE/rIzfzpyiVYHonAAAhIb1A2yF3k+754oCLTUT9
L9heANBYoNYYUvYec4S+gDo7wXgk1XqYka5slmAFGTLdOZe0ASUcaEkg8OGJGK2C
nch3KXapOsLXVezwq6ERmfk+SmBvXPQywhu+LqLMvSYJEOvP4jmOGRkQ8eqi9k7b
nAnK6V54JhDrvbwDmdj3nASx92ZJHul4+hNTQ1lKzG6rH7Cu/cYyC7DxzbsY8C4N
vw/p4OeOlzH1MUpEInP3k5OHFNPhOWk9/cKw/r9eTr4Cq6AN4aDHwxLptUPtu09w
hqwcd4/SQ6Xx/M9kwSldKQfD9utTL1TzdaXCg5wdvxyNDSSSUUsg3FV6dQDRAlDx
ddgjYWBfBLbDklyhxfKHoTOiLOY7A+NUMOr+Fzfn9rTSZlUvM5X3Es/gdncNJPx0
ijsPJIq3mvhBfuqVJDjQ6WQXolzGA5SK1Hu+x8LBjUO2NJLW7bkq8Lhasn2bqgyG
qIl/SY/icqjBcU0h4wI1UEbGBRuVXQhomZ/3/2ph6OL02pRD6VE7vttHrgSSkd+i
Chqec4vQ0KNK5hO2G8z6Hpt6c5Yvj+Zq0H6S4GXJDq6pDsOjszM2RrMigaggMnWR
6/pZ3z6kePLC7R+qALcZMUICM+skACWUixcYWGGVzscFnMn1B1ZDyu5+k9lHYs63
FRUzWLKWx04+5PkDtVv16WdjXBcZB9TrpIpUamj0+D7bnXX3ON5s6CL4HyIb40Kd
9zGNnA6Lb1rhz4nEc7j1njplXzWW1acCX6YUko6E1xKubOt4Pq/FiuBpv5x9/L+g
pjCTcj25JKty9jmXdsCbFkKwR4GVJ826gUu269WDi4jQ5Er2GzuHRA5+C3Mtvi59
PT9/kipNnwZRFmkDMqVGclxUzqTO2rw+Q9HzAaWYatA+VI4YnDI/qjVzQ2re785I
5x2lrnfDOSXEZ5sT/bYKPJvK49kmckeP6ZkmR1tVCZAKOA5h4glEK2Ly3aiNCt3L
Ky3EqCZCIlo+6uVl00mUm099Oa7QXLu/G+6z7XnBLgwm+JDoCh5CKOnKCj346mNg
W+mstLoQEDSrysRMV4mnxPPzDxe+iuhwtNl9du8sd9A1ukpPcnEIc0wd+7ox0tl4
/LTRybaAIvDos41Sw6r8FTno7jolMKQUxySHltv2A7yWoIns75BEY70yLLOFJI/A
vHskTW5INVzvtcA8gNiDSlLXfaF4X1/ZT1qTB7zICpzuHNhoAjEX1hss/XrI8oLd
nAQviAruswViDWxbGGzZR/xwrrK4HvIAQwCeq+u5osKW4igolkD+UTN94jyp0L9r
mU4VQfjBsBvpTEHW9qShO+ela8PaRsRj0gJXAVCGwlproTLp+dYfelsSWL1pmYoe
AzO+hTp775t2ZRM7TifQ77j+uID8AmIciYNjwq/7FyUO8n77jwFg4/YkzOXfU2fJ
KdiDBupJCOWtW36Y1MFOJY3GAknQK43gwtZXL9wZLhmxEcGt69S1/SSydmtOG9ZR
9ClaHPYfp6tgrHTddxU8pBx/ewQTiqt1nZmZTgyMbNNym8S+v0rb4xgvhDJBpCfX
XGde5IP0Y6HEi25d4vaAsfgByneeLSx9F41RLT9VJhADOLIL2b+XCqk6QjPVqyib
gZTqdnP/ZunzFDighql95iVudxa6Njh4tZ1AbEWgEs1+a7XoA3ipt/qN45mc1v7F
gBRqv+wzLnbg40l64Y0RFtT4yobtu/OyPqzPoTbFF74vyXt2zD77uoqyrxkp91vX
QhsOQ+2C+Okc979sELGU/v7KKfqkDNsE+zeRbFVHKxL+KtwP9Uxf68CXgghckeg6
TspzTITNsHSzuKzrSlBgGymgTMmFzsaNFDPGXDlNUuauKbinnKc5zxHOER1VWos3
3uDYWd0w0cnD8wBnKao1ZICKeOCrxE1clMCsjJZEWydI9b8NdoYFoUycRE54tnpK
qTbep9ehiNiyY6Ju6q9hx8fjTiGrxqEJKtjuMZSjIkSBOhTdtY1GlXkFT1v9INo6
zcEP1M/WZVYnDQJiki/ZpFzVB7rLk76+lIy8syS84jIQQFO2bJ+BjHqH3YP9/dY5
Z+uUb0aJM88Lj5LoVMfaYTaWdAX20J4vuou2HRlkvkDnBfNqOhyzTkqTD8JSMaip
8PHE3YK81GT8/gKsYAygk6z/qebf8fk4l2/yPmzPXtd2QYp4V91ieP60q0XMSECb
+JTe0qemGviT8QEOIVrR3DoAERJG4ZJab+f8kktRPHCffldLJKKg3IFS/8BiwY2I
a+DzbRgS51KNNE4eUKkS5/nwohp0J40/LpIvKMGMinaFp3UXYbQ82ihYW4UXDka6
zLs8pvuZmEnYm0Y2k6oU4j5q9TrFsTb+HQK+fWSvCjFcsXY8ragrhAj+m4zS2uIZ
HBoCzkwgzoI73MUW8QIEjOht3T0tHuw0mZjex9+MmuvdlDJspr9VosoHJF5Xx+NR
aYd/vlprdv/7nCZKo55zxjKPNa8wLAh3JGlzlHOI/ezXPZzIgH8JDnI+1+2njaeT
lTZt/659xzn5q36WjC0up9NYGlU8zBlI/QDpgQdz8Efvrh3+QbwBV0/vBdN8kggC
K7FPXN/S5oCnuZDKY4b83S0HLYwiwAsEcjcikhCa5WFV+Cp9YdYtj6NhwcID0sbz
nLBqpWIwyDR/tz5+PhX84n2FDmWYloOdMgtxfHZ4Laq+gn/kfqRHY4rIkYB67POu
9d1PJJP+4xjCc/p32nlPAkKFfRQPH5Iuy+ibRBKO3HLsFXFn57EcZYdJgp1lB+4h
oSoeNuLUFZ9NQV+71Z4wegsRMQuVc5ro+46QN2XjgJRbivzSNnmBfyNRssvpxWvp
qyXzTbaUglPukqem80j/1idjjyKWW3gn405Yii75ZufZybjoiM2Cz6kQqKDH9v6r
YHuZDqNwnhz+caXTmllXerBnciTYBGgdfX1PYQ91ZiMVi8LGfJtSHME8B8t+ErFB
CtlIHoFa4IZ1bWYJNRz5qH3w8xj0RnMUdqcqfMbo/rENaExiNdTwsMbgaUV3zlah
mza9OF9lis7RxiNSZfYq9nbFujHrI8vF2o1VTkL9i4MZpuOx+qDx9hxDbakPvuXX
Le9cqGLXrSXesL1jl5l9r2pHau4fMW4UvojII6quui1GoKYJ8K41zsUEZrlLpzvs
kitZvvwoH6pk30NFn8npp/1IMmBq2/UOP1N3u+WPads4w0/BLPQFrm4//RwFrWpt
cCRH9GdZvTeP251kTC5YFA/HC6oGqo+CM5kBE8jIDPCIAroOG/MGAjsvhWR2sBDr
SFBxhR6dAMBFonKu3TGchV66Ym4mK3wMD4MuCsx4AGzQ9CAbERV9Pmz8kFqZQhef
4JGvWgyKtJedIeRhvYozUBZGi1jGadKm1SNo52jw+pJMuCETbF5aKvX7y1CSBb5c
+CuaaC22RT7c5hmjOtk3VwsFWEKUzUYBlIHPh7CIK20PKHhLEpwmPPtJ4RA7vJYf
k+i1l8Su4O6o2reSwyk9IweTLVZlguClZe0qbthnfxESVygY7E6SPRLE52waqWbE
SkHXk+WSpgYxAsk26/bkQc6zB/ORUijhCdwYMj4sceeCTRJsOQlJz5u5lporO+Qi
IAX472Xi75Wlcjomt68lX0G0Xw1jkhTt2kk+GTD8X42hZazklmEjSli4mld0wfkr
NBb7C9IVF9/oNzooZK+5Pm+HGnAlDgWu4Z5WF24fMW+R6SwBmw8ESru8193uAa2h
r2JjPvFm9Youmrnz5ltyoKSPo27B3i1snw4Bo1esdNiI4gvKmLPukANQtLbaXXqp
hsZ55TiD9UNyBrVuPzP8Qxp5RA9sELeI8r0xT0GRL9iOOI++Cll35r+HQ+2sY4Vq
10xpvOkfs6MY3nOROF0046v3ThjdDAhmoHl3AdkwNcY6L1A4lx3sLb/0m8kUFR/W
/rbGBBR1Itpb04SIZODkVXCpPoZG9Le9mv+rMj+msJqF3kjMsllvAsXXcZckq3Pg
+o90hLdInBdpVHLiMwtlMyaTIeoquWs8IoIh/Za/QqWNdr3aHaBRaDHIgtfPOqsJ
r+up9+YRwocx0X/RaM8uQ/yCxc1TBC2WZ+6cjusiNgHM0shW/VgiuixnK9UsV4WG
nbVxHWsY4mjz6eyynUariOQX550zUPGkOm63fN//eh4jFeCvvRpUVzwPJKCMA6wA
WejTQN4s6jXmURxY+SJauZIElFmTpiBldR4e4lXD78Ef8TzIfGc6n4k+21WmxpWW
PB25oiHCpXaST222W2Rc18f7vN9QovH9UMWuc0NiK3Kskxzdvzy3cHLqyGCPGgsD
n9AhCTz3XsRu//if4KwpYfVkK34xmjVEzR5HsH1vJDnbSg6TfwYvPKK8fvojaXKq
nA5uQHqZgbHGAEaoMk9Nys2IlCA88w4VSPGrg7eSPS7LG0D9IgCsrTwN2pCZpDhx
ywyuDdOeYsmFwllnS/ijTx9quptxhdAziXLWr//OCdB5MDxo65TFPLhC/DP1bTdM
4io+RF0USCpV4HeM/umGR7guzRm9bBTBdY2rNJTTmhcjQ9BLkYFd82NhgaJcU3dW
27na5IznyfgQmiEnQcFhmqKlYd01LATItu7khuBW8N6xYc1rJHFnvnneI9LexT5y
2ipU2kKJ8vCHB5pL5V/9jvTUevJpq9rqFLyWr0SH+0duLQY2oEmw5E0VCRD1Un0u
Lc1JdZZNy522sndQGY3kfhXQ796fgEibPGbdUsf9aOxVSF9V8PrdtM4UX8qEaU7Y
cnRp+slOEhjfmRaxfUCKkosXCTTl6r+ebITHo8v2YCgxOFbrEN8gplLuGOB2eg1c
f1fBdSdeVZtmc055jsPF0oaZWBhrZ4EpgxAX0iMkh1InkKWdx0k3WTDXozAu/8pO
PsIb98cK8gw2kUoVghuWJA5dKrbYyVyvYFg2YCBDMCgpFLqxVeUeMH8Gzex9BgPS
NJZZf1lm4oGoZUNYadU60mZWgIjvI4NKbFWtcTqL/SjLygVvsJRRlp7jjSdmjGrU
RbZxfiOJdLmpbd9zHjKaK+C0G2zb8GEh0USS+/JXZG6qU+n/EJOhO69b7TWG1x1A
S5w+8nQ37x7+5hzV94cK41xZfpI5YjBp/FwD7fwc+73FiCXzi7/dKPvXn6CqCI5d
puxmAtbA3Lu7kXsVBGsLWkQdTczMoekvJCK3T5nYyQLjQHEA0Wudqk433xWL4dNO
FD0zW7Uuc0nrnqICy+pcTUiv0olAVDlXazvQLpTY4kJH8Pbx1zz9AbvOTIeQj5MZ
QBpitdKMA7h+tfomFi+A9oOHjAjLjog2PCq7dVfqJii7KbY1ds0HRNztw+ftFnqG
Gy8V/PsfdlqLeQF0PdonwL4nNYmQRTghFotiU8HthGfECBldP5DXySDQFVNUWVT4
PL1HVVfklCtQnF3Vez+uFhHuxrRSS2DDpELG7+8CO6iqvCxJm1Gn5MTM0Swmlef+
HWTsDwN0pjRhIuyyjKjlg67Rn09Tc47pWt2cAUntf3g+Q0vHjwr8FOUKdELItRXM
MuaVdzcVhQU0UdYrKgIIjJj9vfc6x+OMnd7faK6sPLYmo9QoLL157CNvKqf57t4A
wClqNJ4FQQFk0oUfjFIxwhWWKUPrKMYByAc+h2nfYfFq+1KUupF7ye+Yu/uux5NF
tLg8XlU/lkSwbWRfUJuqE6SasqlNtdTNcUOYtBshaQyid/P1z2zbLX8DLx46u6Gt
8i+zKOavWCdkMeFg+MgatAtLTuiVKo5E8UMb3nYFSN31JcMLnRs/WxZNkgEqj7jH
Qr/Nlww0sVnvKs8THEUqx2ulYNSxfAHJ1fLytz0HxfsPDdcnuND5Y0kFgwaW0w89
8ZoybnJVp0dUlqcVIOwzw6PQCm9NFxHxYMBO4geF6qu0Lh2wjEbXhQ1nJUyHfsRV
3QnjgNzwhiCELCAniPJJgMJ8UGxWuqKftkPd1/PmRQFumIPWtraJFaHes8uNB6ZV
PH7kNC8hMPWv/QuAJjBttrI+A4gg7e/FhRD5+TtULPtNUTEhdkhgPwN7eUdAUgbn
mNoGItvgwI+uCtCqsKP0qpQ1ihKrItPR7BrKqWOh3rwf4ak7GzyCMIbj0mjgvklk
q1+G364XICCIXQQIQoVf+dCLXWiEiAm0LidbUJWkqKJkblwRSGavaiWICW/rqaTl
2OccYu3EsyLwkxL9hVkQx3cIeLyux8tz8zvCq8Y8EmmTQA0zl2p/fKtBq0tT8is/
pQ2VMZgcB4zf87ppE5cGkccWcNCyIn4Fdy/OvBdW+QqpJ517aRmoL1lJnZim1eQU
V/eVxruRqDi5PCL5qKQToxHONjd1mMDseSyOYPGYQ6hIPhjYwtU5gh6X2Uso9V8h
Qqw7/izyAHZgl9k5F2+dZFzc37bqyque6eRY4QFrOVBm6ega49xauX/ZzPYK/enl
wWEQ/rifDRg8NO0gdv8uz6IztJuR+nSPpQs+kphdiieGouNuYrg52vngx+dTVArl
CBN9Y/IeYKp5RzjHzLncRx0Y5SxLev1Y9uWgPC4ncpojd7kjdrg7S/pK0T76UqLs
NwhRz4d+LCQS9cw/9JjoqtEy9T+Q/kNtlXwT9w/ezRA6WINuc87+VkChKlTZDN9O
1zmC/CDusjOCu42vULp5xQUOfw5dDy0CWhxbH2t4kgE31D7JeLzW3jsc2ARkEfjd
AwAqPyTv6VLkZW6J0O/C3++O+oEhsnLzgfo3e88inF82lv5iA8jPaIHiqQplUqkn
x3XS0tDQ32Fb4MLz3VFNhEiWS4pxiPv9ZxYrQJJhteN++JWik0k6m14EgoaHsFBT
CO45I4r88cqDQ0ToFkgUDRoBrXxz2JTb76VHA1mGmahFnfkggKPobM1PZiBjYHFl
QmqW82+u5bi2v7asb+bAlSvE0CfXhiAHOuK+wma1mmFaQREaoWcpASWIYShPOgLP
FVzLdtkS2yNEZ1mrXuV3Rq5fr6n0dkxVGUnrGiyuIeybJsfiv5bSu4JjacmDcFdZ
YD3UGMIyxhUuEz1vZdNFJrM/SaqCtddwPTOVyKzxq/nnoLd8U4mU8AiSABufzV0q
RVkOgJJgqfPUNQFXbgmPg3tpmkRS5OUdeMOShOviCen4pMkuGqNYnnpZwDl8ejyC
HoyVzECPF0cf66uaaObeGo8PRhUA6h5rA98z2Od86dHva4Y2H0yaFMFodTOvxPwb
rSmNTYEWSx73aO6vk7KDaQpBJ2zn0WQrIzrKlwEpEbLLLGgizPGzUj37hcWpnEks
pBkYyMI/SOmBXSdiYOnA1oY6zFfyDGideo7gGEnuckRHKaFf6hjW9K2VYQ5tO/6F
ym1oSjeLW4Q7ShWCWmL1wgl18dJJ8rTkrvgGBFhZWlJgI6ueFVwPlpNPfbISidW+
qj2w6xnUTuNjXgqbf9mKWud88a8T4/xGIsrpUfBb0lgboW9vIHoN5sgjHt2brVE5
PQTjDNm6rKIuXS0xorev4hBJFEowGDoOSeeZ3ltMvr3AgiaRpVNuoWAcbD8HeZCk
FqBmDZk5clDdwl22D6vtvwAVHRlnrx7JMC8W+DvbwSYDmGry4nEab1lYO3FgVb1x
1RQ99uo+dQd/jDbJnRx5shgxp8NkblVHLqy/bBb8zmg8fmVccs5TbOXpUL9E1637
H6bEb9T+w+9TFJTeHe6sQ8icI0LfWUPUTNKQnVIu1GIcDxp717iHbVmGyUy2gJmv
FZ1k2lmrVu7s39fY8FE7TQWUOG09fwt6gAwt//MIHYrXTfJosIWiF9o1VuuXB3Wp
0m8u94eOs/mnxV2wswLbF17deC6TBtIJunl8jO0wrMaGDqtGPoRdAKcaExdTnmet
0MAN/3SJ6f+lcQs+sTTQUDkCGCthl+WEmE2mGtIR4ivGNjuXA9mgFVRP02wAKU5J
JGGEbAgv+RgKO8S9dLj85w/81tU60JhMNWtsAB1UIbLHdSpCe7UKB3cydMQE1OQL
bWEbGUwVsBOP9EWKM0v6vlx72zh3jJesfnkKFlsBjd9YEcIBIGqMXRxqk3JPf/FI
oKtyCmyUQl/eKfADMXQr8DGKJcKMdo8KXtm/FiwsqRucWM9EgrfvDohG7X+4LrWY
ANarPOi52hLU9lq9UCeecREoU2AeYOD76NZXa5/lGYnlQWNTg1YLaK18KcBqp+pE
KpfrsBxCulNV68deXJp3a0j6XyDJ1Jzu9SetsUECZKghC8d0cdSqGdWAKVC4+gNh
cd4FsNWf/0juRiVfTlhQsTgCA18mwPCURjbhAwtUtxBAgcqBHVtdKmQapO+Ftpmo
hrlZqUAniYLeUMOiHHhQ9w6PJpFncQ3/nSLINGVttP/czhRHt7Ml8/HhFUuz06f8
eDKa3WfEf+NhwwQtH1nrC8FvBdTxK6+TxYiCDprUw+xvQO0d2mFolU7vtA9vHdcR
Y+xMKGOk+umGbeVzJbT4uQ/OprFIrmY3YmG8mLmgtAKy3mQUQ/DV7PYy1x9uiav8
6KwMZUCFHtEEIaKxtudaCeJPHO47E6xVeiDZmVYeEB4qZm6EBjc3tueQ16gBOP4j
MCuLuIxr2Mw07CDDsjZOuJ38T7alKgT/14ye25RoWaFg+kBwSly9OfC6hvBMSdXu
2T0gS9lWgeTNmfNaQFLkc5kk/qgVe8mPPhrusDt+rWwSIwneN+5iOttb8TUqf+D5
6QwxIaYc/9mvQLS065UjBXNkmPXMGasLTnwfJluwNM+5XZ+FfoccaPAwatkFhd74
t/mp+MupVjKXFfCEJHongDkkgpj9nkY3btrGVa1USOxmhcDzhbJFEC74VEldvA6k
6mfdhfNwuCXxm1dbnY5YODXt9uVwzE5QkA9YYFkXho+eG+WdxOwFdtDU4qLdavS5
QBPZBNOZcUAT+Qr9kKHuWhWsqae7wVuZimDlj2ifoEcbnbJWrN0ROWafegNOCRTd
bLXAH9sGWhSPEtaWRp6eDhnA9vO2MpwOvO8++x3dJM72brzC3vYVEh51unzhPZAU
GhW9RVPGqVujf3jn9+kenGrLnPcyUF1yB/YDXPwbTxsIyu6NC2T0wGCfneWSz8wR
sv51fG9C/gxn+90V8ll+dxUMNv7hJASI3WFjvF2vMkbbQm89VMHsQIBssGvZyuL2
gwW7g99m7Y07qO8Nb3SCQEYmIwX7dA45AzEr+ZkksA9LvBThmt/xPQqUeB5XPf5C
BGpzn3KpOgweK0PFyx9ndi3+nW5+sRi+WjhmfWS9JjiGOYOl4JjH0Bok9wAu6EBb
PNb5yW4V4Ja7TRV6zN2hZOImMfw3yNyfrke0U85QCf+3Q8LIQ7QgKjuXgsnIv1mA
zo75z9CN2jb8BO/B0MtgCRk+uNGPd2tMJJ1zJZnyyJhG4kO9OH4MxZLjjgilBojC
46+LUujpnpbqV7owcKTPiOevVQY9uxfSjcuPxIWJn2j5MXMxWcsdII7Q9ixdn8RQ
9ZHDDnzqMZVDXd1Nufy5CaF/J26Df//tLF695sZHemG8PcpciFOojgtgdf2FWNhq
OcAY/jCsWab7cG6/30V5jYqy/bn7mGhqbuBBx6KDUPcBEjdcOy75jKEW5CLEcF6G
3BK4gDOTwzmDhrOx3XVDfR93oUFdtCLlt9TblvrqmOsHrtMNFVh2NBGhlTqd66Zh
sIZEldlVxsWHJZlbxzEvU6Eqg27PmJl3dbQ0s6UK7FkdGf2qILFny3VP+7kbaE3j
fud3IcVyPTSl2oWv2mFGrt3RWfLwrGIgUzlopFXEYsFiK3C6Cf6ydyvT9gWDkTv9
gVEA7k3CWEJeK89L69VkVqdrBkJ8kPKhHfKM1nl9Co77vhnvIcn7gDZZ1xIsTfK1
bCRfn/8C2NyXhs5RtNPxeMtIwAywEjawwBCvCDPBZep+nQD9/OJX5CABx9nBVMfS
XkYY6/ObHidjWhS2DwXnh1QS6PXj9xvHe+9zaoAGi+B0OMuxln0thff/t8gh3YbZ
CbSf7h36O7co0+QXpXZsYDRY9BduqECOWL7dHcbu6LPeMdPYY0iBBWfpiV4fzhLC
/gEE1sCULrng5XgjMd8JTR3aE3pXDjxMzKMLjIoMgX9+YyFFQLkiven1eO/jC5Hb
YXN+4Dm420JBYtiX0wqoEiLO5iRCXy72DLSFZpNV63f6pqzQxWri/kaUW7g2fudl
RBgM/5J1E4Jkc0QptUKfaGMWi5Vxs5jsD41v0Va6vgM5dgo6NgsUkl9LDRQufac8
IoCRz20pwx4/F0eQMTbfQ3yf3kJp/Rl1/ilLYaIu4ppeZ0zLhybu8gwoewQLtWgY
NAOd8+fgMuJvdyz+EIFNJURbZOPoT+15LHwyV6x3CZ8ar0YBaCgFusvURE8jmlkF
OchkKbhvE77zImxNb3EVOJdGaCZX0Fy//wO54+1NVKgsszx3tA8RDLKExZy+K9+M
KYS+JJJnenrLkMJQza1eSs9w5065AROF1AS90K2/bG97jyM73GQFDSN4TRxC/yAt
mZY1a0EQajA8PH8tWYiSdBZDIZl4kwLvgUmohGy1lBOYeq73bknJyXhXg5G9gFl5
jnnM/veNezZMH1uGkcN63iToYjOJCmpjWUIl4AT+hijKOk8NmeXuXvc5oohx7EPK
dF/UUZwlwJuvlN6vNky/vW0ixSe49xE9fH9QuCLEOonXOrnoeEHaZgEfXfrJTFez
4VKEZ4I0eiqTTTqWY/W4rvg8bMIshflfXDQXp/GhhCNa6j9ZXmVhM1LXQ4j17KHW
3NEZjQJaRJ8UOVCV/LkvlzfIYQrbnVUfU04P1kmAlAr/9YwrgFjj6/iP7AJykz/c
cCZeMXbggrTcc0Crrh2dUCvGBl+TmLDvHz3krueaDQ7LJm1bNPsmET8+YR0DaA+F
ImTcrHe28+AnS/3UAlWncLIKg9qVBNQGDQc+pY1Yt9R6tttimv9uIe+8fUw7Y0+d
x0sunm2fYssUnP1E7JTHZgB67YWCTwEpF0QzCyhMPd3TPL0LAhLMEzsc8Ap2vSs+
ROty/rLFwy2tYOdXsH/KPyp3DlbVKVgr5USOwHiOnjagIY8aPbSbUw8b6cLsSuMC
uzvW/mbBYSCVyLHZJRIAKJTRIjLq0x7/pW0BfpyJj//fCt1d3y2OfHNEDh0BBUwB
LGQeN4hvh0G3gTNqIsx8Wu+nL6NOK0QUXYRHtJCmOSRmzkQS7Ds0spsrblQL9TwX
keY0i3hwwStJXBo+IjHAID28kTrqP291IlJO8JaUhtm1pZRNZxBzMNrzBFkBCWuI
dC+F2s6YxUVwtgc8FnO41loHsfZoDJLP982XlmAQpwZq3HHBuvyNfcPQukAlxjHx
QhSjsElgb+ADZuid+lMrma2+VIuKhprmZgSRHlE2pR7+n5iPgufy31F4suWkO5gy
caPAJS/oYrMK2n8rlmnoxSFmNscxRFCwQco1nBx7RvXz+P73lFM8JjnP1LaBS8sy
IA8E5Mvr40LeUyKrbBeqiJ25zdY6W0wRF0mR5YVCs66mGZ6x+5RQPkde5FhQUUIw
YcQDK+lUk2HQJl2jCn3mrwFjm86PsNW6XerRUxLK8EprUpNkyWk/zLJeBUeE6P46
5NkR/AcDwSCUoXiz5sfQO6ZKEyaKI0XjJVRgHpZQvJzR8Pjm6ibD1J2Yjn4LdAvt
nw9rjwSGZFnwML8Vtm4xUTxO3aKpFtRPJh8oSzBkv1Gr65rGyqHakRu9MQLuG7DC
fk+EiNSSF7TVwAH7+eyx84lkWDx2c6SL3qdi5oAlWbUyywMcJPIJYnOUwtk3IMjG
eybvbB4vjVgW+SWjExVSgj/HYqz7jvMVFpqr7J7OfqZu4UK5fPdQaUALldhXYDGZ
PLqpScug18rigyZxJM8NZPEP3rSkI5wqEII8I9++c9+D+9cO7bFyaVQSOPXZMUry
24sTQj7KFPTCaGZJ0MqFd9YmFIYgf+IymyHt90QujMNz0O84NJ3CecA47QB/DOCs
5HWu1RqGszGmF+Ryj8/YwwIXovRZ+evDBt+/CFiEleMmYZ2nXoYe3nMBlyKkuk/H
YVE2jqpMfM+JiYrjz4nbFLL+QI0hdJ1F5NERfZELurEl0L9miyNLVK7qR0h2B7Sm
vXq42bhbusRDH81qLzfwSnfDfs3NTOsnJfxLEtKweP/eW+QnYZBab15IhSvWEskT
gzkGs6lj+kOLALpKepck0z4OZl7kLgTC/1aPc9/wHQG89MXUgnbw6n4kGdVNlAYb
QoA5YliSUm6qI5bV7F5pZ+3iAnoWt3jbz81+ZbvF0yZy5TU94Ao8L+ubbqQ75z12
icjB2HQvH0w8gkVd2aIKkFxN1Ioh30okZ4QQ2RyXY4toeDip24ZpoZBjoMjAP/5y
opcs8TR4AAskBRPBmrNHhDh5z6s5Sv4uJttOtMpKzerMOLOIeSlakTknH6wffWyN
kXFJucUlmXDcE6frjRduaUKX1V3r/YR0wN5E2wqXQat5o26uBZ3oKVZDhUBngGfM
lN7fmGL3k5fxoZ1M0kI77hFuQky8fbLcS8hwsBTBvxGLIvaUlwK3KUyMvqeYeJBC
3dhk34bE9ryy5HI7quZlOxJSiNJEEiOtXAtpwUaskyvbvfHw31UlGvVZ/HUWeqXs
6ZfmpLT/3Sg8RpImi0bbedELAWljBwn8QAxkNKAMycd460xYlKOJRSwobP7YsvtK
xv7RIlzpkVKLVG6Qn7cj5gN0mmNMnCXXHixBfA6jnx+BWAK6TgqFQHpEqMHRk/pZ
lyC6u+7cIPsA4oe6PDkzIX8AZjPv10mZUjpL0Dg6r5xQaSYqy3K113mI6fMrPssb
y0KvTjWzlUIv30UD2zZfqVaiDLXkZSYY8mbbun4BUSFVi/R1XBP9VtQcpahTkfNx
FDxfrW496vHzW/rJmLfNrqErHpsRtUAJSBnMkDhkz/9+E8YCbUgx3jBaVg8xFpi3
MihOFg83L2X1qhkUqGG+LVB6t3PyE4wGcVYwnAoDeDmflFLorBctxgc3tmzYXfIe
gKzzn3OhvNaoQ3hdbVMAdIcaNSUthZXDFnrOT9lBvgwC6rZEMCvE+H99h44rOKkT
bC+ZZ7NejGdE1t4PA9Q7hoetyuvLIbDgHxjdIPyk3G01lLive2ALvNUdx25tNlXz
mB1emhvoqIvEmDwK35PQRAjuWChJsID7pgvuLq1oOA3yWBjG36w3ZbuiCajnS6ke
DXw9Sb31ySny9lnCOe0twc328gsMph3nOUJBmJMuD3eZTlfLHj2tIkD9rTpT2D06
j8v+OBw+0ouFohP8tH3H/q7H9dhUCSeJpt1UD1djHVgWlj9WZU/GuPougjsqR2M/
FsHajfo1d7C68uxICmbyjDfbarDiprhRg//v3A61oFL5vW5Ko09YDHuIR6L4nd7L
VeibG/4GbQMFZv8la6I6oL6CF/xhSUNJPUFGeLpHt2u8wIBpzimpvliXS2mqlj6K
9jjpTyjtcOTcBzFxh6h9N8i4fOGlLAyAAilqPjTJyV0w6OebVZR2OCNdsMY70Ovs
RucXazyb8oqvzyQSL/1oYQ+qSrGTk45y3kPut9k8AQUtp30zadnJ9woMeU3bnEre
iomcCVYV5PryQvuxJsizyG23+BJmSDaAZwRgq6h6Z29+KGCzqr/fWAvLoHrAO18I
xXw82qr0UMcnQkURNUeAqAFWsP6ZRAq7kP2GTjl3Dal8JP3XnYFZwGo42MyqM4aW
FePUzkOHSxJj/jIWZL+K0bwkWuNH9RCxRFutYLnlcFkN3UAAP5FBUTi4x8F79H5H
Dbf4CmWQSDRXC5ANar91SZaOEL3vwTvTSetn9RR+AVgJqrs3tz8KBjqK+gqAjtm0
7gUWogVj6sr5W43tGA/7T5lUADstMvfyBMdh+acttQ1EynlXTWjB4WoGvWE3b4PU
f2GeQhNFLQoJ2pvcTlYBsM/kZL8Ev54GKP89inXVPLYD6onyEFIdWRDiiOgUUfa9
OKFeFd3aDjzLdLjuHa6sCRv9GJEqUw96TacXH1dMtYABN7/uUsStrUMWbEbzJUIK
UlBME52XywEbgaWGM2anm6tM6k/VxSZ0c8Kct1LU2998bOv3JRG2WUt3IJ8KVjUY
qVpVip0cfgJCwF3mSXSbva5iSigR/51WDXyP9sIpMOUwMns6sVGBdfOTaFqLrdlz
64K8Dc995Y7Is5FYsPZYBXuUbFCcZ+jNIDCQIYBaioPURS8iJUOhv/lpdLS7x4aw
/HjGJ2BvaxleRDwty6CRHakou5GJWEBSlpGuLPDenDEK+pN09Q7h+UYAR4QFILm+
CDf2nqDWdFmOIHxusb2UrQz03JxAHoxw9hUDJE2J18cr6tN5dLG4i4l846MyxNL+
BvX5NLt/dHa9xSlej5KZoIl7KfJ6nl7A7xFv/IFdk0YvLE336CAyXkEbBjVw1TqF
KxGBqDsrk9/SpbWlB9RZq3xrE0BUl1jec/dAVVBWvVgBR+S3VJiEd8bKclPZJs8Q
iAJMlubNu1/izib8bDpPxP8yjzG8ncZRi8jUQ2s2oz2XAs+o0HdTUxY1DOzjo1P1
x3CMX9sHRcUrxFNnY3OV4v61bPnooC2uwHB31EqL6hr6ac2f6RcXx3Rfc3PJarR0
T9rVL13sJ8p27A1XZLa3vfmmGRIIqTtpIwN9WqwFYwKS8uNyqlb/C8ci2Afa4yic
WmacZOk4ySSDqmOR8TQw+mWvH2iRcViUNwjW4oz0xOAgwCpKj55EnbTLqQCaKVGx
EoYsUQXO+ID0gIrOogq9vbt5/sAALpkn8+1sffMdNG3odKFQiujvPhKWLjTukFSL
14aa3Pa9vYB2u0zAmY2D+RnNyZ0nZaDGCz4kWmec12XNAB9MOCQtNDlUE0x0C36q
3BpnwPjFwH4UA/7xQlFrLHwROQbWie7ErEgvSZH0aWBOwtHuKqQ91tfGVEEsoLjd
73AC32Ru9lxE6XNwiPNn2huM9vFrd8Ub2V9t0cLeLNf1IcODNnojadOmdcNaFvKL
Ec4vaWfL/NHSwKYuFzkO2RSwievON7I5aOcUUDS+S1aUnHCfngpyENYLWSVaz7sl
BOOlWLbFpTG8MnNbh7aiuRvg2XioQLTI9yCAab3h5il2N8Uif6SJJkEcxvk6HbGg
IFaD3szxyZA4yPa3lq0y4rNNhJnzqZs1y4JKSxIKDThK+HfxeJ0BV4UMQyzCHD12
7plKHtK8E+Yg+4HXVG3pUpYHsoQTCTOFiavNgUGk036WVg76l5iWig1L27KvofSm
NzZ92WEQak/gHif9I6ECr+Qafg04z19LVAuqDGqdZNAacztQl7jwWfoJaIuRXPxl
c6E98+LZQaSJJdVjIWhEOYOK/bvY2bn/lDzJGu/kO5XhHqVxUkky+jQInQpuQcOW
Kbrr8yfVw/wRIGGljrXM4y/TkamrRaOSrkZL3djQZP6r7ZJcMBOesFgGzUtvKp99
1tXCE3o7mIYe+XVwi7118I8t4nUHUL21+775x/v0pOWaEdWqkHTwWZCvqSNl6JZe
KLnChG0HEqZ9G/bOTiKPYbW8UOKnqAEmF4q5dnPJCEU7np6jVMkyR6IuXxFuZybX
djdDHNf2mLim0JGJD5UmjZTth9GPKOYq+dfF/jdBcatYS0qIJfQknqMnOsMZLx/R
OdgFt8Oto0NIcewu8fpn3s+o0uvheb9ToZTBSYY1Wv4jOVkNQJLtBviwE+WZYGem
YKsHJYqcZVZ2qo4H77EO8MPshHsiIv1wwZk61VInoVdy4tcGq4LJj38ulxKGkdnX
jHzktxzyjhbieNFhRSYY8nw9H3vSAgN2Yu2nHSkWrpA1Jyb4hJSsLYSkWJpJnS72
eFnKHQc/gELioteFkUc6SzMVEXURxP0+oQWuEFiTpbwuKW4qc7c0PUzfE2EOTy/r
QTjFxSBCr3Ov7TJjhk9X0Jl3E08l+kkc5ARzxDycDlqTQvicSV2qXhGwxAXXZsj/
HbFCm3WXJxPFVAzw06EKhzvQy0XDmG5r1KksHr6d5GQH+gUlSLzfYCFLF+9DQQda
0NgFnJTCzBDmfFyUDTPD1dsVkyNJd1aXbJmIAv+7aWvyYzpsPDvC48IC9IKoRU+8
8Vk7jlQ7BPaTRxeeIzanVucIhGxrrgAiusH3xZJft5JCZKTVzQoq/8+ApwfziyOF
8YdRikQLZ+Wc2has07CQV4k5tUrig21cM6PvdwVYO9vmE26DESgAAhQgMoLPvzsC
0+DHqXnJnP9Ncyu3NCiijiFF6hJrXeMHyHOps4zV/lYGFOS19t3yPhN/3HYCoVGz
bfPkaHR1MH8Mt1z2PcmbRL1SZwREpZz+pTFsAukb5JwWpuFZV0imyFqhomyOVOZN
1mHEcbTB8WQ6BR6aIW9qp6XmX9rY++t3TOhukgeVg9puGT5yYqwvco6Vgf3XN/i9
CL2TjDAd2VwnjZC6QwszANr1fZtFOh6zs052oUrxGQFgjf9dASGAioT760OrUHe5
+BiCY4V3KQ0RdLmbUkopasfB+pu4hrT3dHkK9kBNUYJ8inpoyxxqCVPO4e4nsHTh
JYds+RONdBmDUVJuU/t8FXV2Y9hYbl3jmEvy2b4QdvwH9H0PUp8n0kOEaZ3Ch5E3
fV5Hn0ysTsAmUogVIOgth4L+DEmBZf/r9Xeifc9iyXfCybYgOE/nmiH4Mkm0hM3C
/BanoKTFHyT/DJNtdrFrJ6Jv1OFJI1R2qbj7NtA43fhnndAQuzB1wrpk3efTXjZf
Hl7mpcLygq5BLamMbNdsANc7uPVmua6k9er29buYXFKQGu9kvYm8lP/2AhoEuJl6
sHdEr85dastcsAh7T/LJUtJzUnaiZr9O5HtSwu91khg8Dccmf6KBgP9QhvZVpK9S
y3QjmJB0dOzm2BdBaAwbb23n4EsOF7eAvQr8Usm20gCbNEn7O2pTBjCHRuUj4hbJ
vGoOYRGKeZSxunNJWE/s0FZlvBQKmKhuFjiuwgRtOeiUv9HY9CObXymRBaw0uqgd
LIZUzz/FqmaTFPvmqzny2bUkkhbBbnhoWH/+bFJjZ4VR+KMrrarTc7xsNfRew9jO
CMEp54HtotFI0tvq5kUQSBi2D7aJihDMS2Lh8BHPr+VLgB37gflDyLBYDCYhVNyG
sgcYNUc4QtI8omYmOjh/s2URlaz0JOqbO2FIifpcaqZ3+D6SFLJbx96myhSkNcJt
3APiuOfGkgeFTbdldS1+7I/TXiiO45NbmoeZkULZ9ossnh1ZYPY7ZyKMnOXLEEmW
8A1WQ5aDxFSMYs8emdEjWnWfHpg0E3cEueYbTtsSiiE2LNEdsAIYZI/VLaoIwHOK
WApj9mujNBPLXPMPIbi51FmXTtHzxtDyg4N73Qhv2vKFMp+JviR0QdwRu09Fi809
hyTpDbjT2VoAjB4vr8FvF/atWo91K6hjoO7eIIUJXMdV/6MyXZmAQSUqSzlNduaz
valIMKCqCGvhrVJiC/G2vcdjCBd+ZSaFSl7YdWlqa5ZUDbfKQ2XW0hg/vwOZm4x3
oImRtYROQT6DoedJ1Hvnw12/XmE3KkfSebCubBS2S12me3m3I7qOb23Rh1XUcrVT
ksQ6SjYJPpnaFhEQb+BXhqAVDEC1RS1C3+kMWgXBY8u3FiB64YtDEgVzPpCf2dHQ
zD6MTp3bHhGNVhNu/YTgErjxrwGq95BMNMj2QYuT+PekX8PLk2rGgpF3TfZ/pjf+
rTjKioyCTIvM7m7EtERzIcini+m9l7Jf6Flccr0A8fgaxOjO6H2OGuUrBmOLPwdY
PF9xPzpdWv9FxRhZxZz2KqxEroEMwj8IY3etgLapEsptgksUF/qmSax+eWsG/hWP
76KyVaNi3FDYl/dBvHfhXeSydePebSI6H7S8ZLKwLa3eynq1XKQcQsQP7oHTER5e
s0TveYt4CdJNtT53BpG0SQ49PTGbYzz0bupNNnd2LNvjr5klBL7zMs5PQWMT5y4I
IaxrHppMiLxjN40pMs94PIn8u+JXVlnEq3cnjCgjd6HjuLvXQACTTBfSQ50BJWAI
7v+ZX6DZXnpS4RbdlmcRf91fao/1ty0cmcUj/0VVmFQcHoEiL7jikvCqWSZwzD6a
H6oH/KndnEbCXN+ruuIooo7T+BNlMG6cxgqyUfWKn9hjNovwLpllH5rMLqKkpZR0
SujUjrcbSMP4mzfBld2UOQTe0VitzxaK3W/0m8lq46IPHWHmOEcykv1Q3bP77HmI
pOdSEnfeSs/cO+YdF8AjmBZO5J0wwvhrrG4DwN8pE5wIbExRJLaop54N6mSsxNAM
jB/Ajihx73opibJa6BXZKvxklM40Zm4iY9svWa+8CPHYRQOO2cNvwK6stvyXfDHE
P+JmrS2uiMl2acEXcRYl+oOSD4MFOBx/29M5ao6OK/PEPlci3i0kcS1INYZr2lNN
6xX6DuFeSH/2VLxU8xTRZfoIWf2bE/X1JodjHqB7yNYAlod1W3D7vdQd2d0DkKWC
IDAk7/jkLM8nb+Ym+6nQZFl1N8BJN2ujnE1q1bat16hBK+FePuYnaJSAd7JRxLZj
Z500iuwP5kqUVzQLc0MVUayLS+l1RAQf1k1OHYs8AicmKBWm5kgJauIClnxN6jaj
KKbjz3+aGRB0WcZs0AbJIo6iXfJ0YPHdXCjjXLuM9AUDpr75nBxoyDjMjNpkG+FU
fJZ2ZVFWkQ9BRazrU4sJeAf68EDO2WuKANc/sgo25iPtrphWYLFLS3LJDRFGSYVv
wIxyzBNT7Ikm6Wl8z6bAp1b8LIanJmotGttrmPJk/ifQoLzXUg55OQPeP1oKNHo3
6jO3ME3EboIBVWPRPZ4XB79jBQWeAw8JcO7nYI2zvxl5AWk4RTjIzTJf+qQ1B9+L
+n44xApbKAo82OVRhsk7H3ukAchfdG29XQu7Iefnjm1M+z//PsFqgGhx7eo8VWFi
aOp1l78qP03rQrxwfkel6+eIIVL4deRdxOLZv28JH11G+i4/fqfvrzLfOIwV/isA
Yhp87XRWnnSto11wfEFPBKBnMEU8lSDkr1qGeIDiu+nvrXZIC/4JEv7y7WTXacqy
Mzv72mJsDZDdMTTmp3DXQv301g5QZ8lTtOWAg3oEqi8JJKyzjRutcxliAMFQoO8H
MVg3IUNfCUd6qZHGcu9PFfGFn8EMIA3YAhIOvVhVwsMMc0y3kiIG/0HxcTHm4fq+
m6nmqKJCzKKn1cTXb17T/Ue8X9awulBIDKKzIFcaaxPM+LXzV4zDTkQjixyvdV+G
0KIvhVmuVuclT5l47JageY9kZxKycVj4vnCRaxKZ13wyXuj33R1MaRep/78CcFfW
pK9AGqTCbNZF18WrEAtp6O9F5gljSZ/iqtOQ3IVCCN8+Y/w+ukNLd3eIcXr5xQK4
vmp/Z5suHzu0/vmBcOONaeVSOm2wqozqidbbZyHPvTy1f1RmgfmJKqlpkXKBVi4x
HWV3FrZUTZrhZo23i4WVlsVolVmzkfbxRPeWWVfI9Fugyh87rhaUfE8SJT09PoF+
/vi0W9YEL2Z0VJ6QpCQQ5axnA4VB0maGxp2OptYH58jHSTvsem24afqbK1yDdn2h
puGhuhqF9DveSZcljvyFz8yS6sp415pU3Z8IC6xkD8qwqgNtCHsph343TMJLh99+
bkkRTh/VGnZB+9cNSzCXStpRkpsyDJUvJvOcj+T9yqquCifaDSTUSIP2hzRPTTvU
CN3/jBHI4oIiRdDdYzm1Egk3dyznKqlm/fsvtKY8w7qsyFm8inUvgnpK3PmLJjyR
NIDkA/piKs9dZvjgmX4Jo9ptB80SVxEZ0+CTbhtzPgO0qjwchsAgir5YbEaRm7hg
lpvdGMfa/BCBI/LOEZMQ3bQqPcijBnRmNrfeD3rPtk7O3Yr2s/Jc8DDg3fnhVlbz
8PAU6L8t4W4IIgvgRiyRs8+VZYByuTGNa83wKKzSeFkoIoFRooDKUflRr0/Y6ObS
2Q/6rHmmtvEf/Y3S3lEvZr45bICHC/bTWUsa6tLnG6LsO4xFHw6Q4RuMnKS6S8Oc
By+dErnwfqoi7qw3pPFJAiqfi5qZXDyO0SPTnosw655mVyJPltbAQqQOS8MZs0hy
UNDz3EQWh+ey6n3U+iytb/ZPe9vlo7PGjlpSJqjiXTOea9VyBf4wBJdllB170J6Y
sTklnhyu6JMRiDgdikVKQxbsepoAMLJXnf0qGRq7+hdpyaUntB58mDp0a/im2u1X
mey/6Y4St5v26kvlrMCvJIiNn+NGmfZAhGST/3QH/0nC4sWHwjqDkoWFvcguT0qI
RSiVPdIO2o61mVFCyXTi24AS2gwK4J/HmZFqfXxVoJleRCIYmJFxEwhx2wHuNxVO
h9HSqr4dGYwvRqbtadqqHE2MlvoI58hO0ZclUr80w0DQVnTr/1NLol95tf+1/ixV
RZCp0ZlIxIS8nXHC28Q7vU979e/mfC8HufeJjlfIMxXD5B1XGdKD045JlL6nm+hr
zdbk0H+XpyuKFQEvW+AjcKudXXC2E+o/jbk+dIAN/hW3UC36oPHjgqUZ62aS+WKJ
78pRumLRaNQpeDN+SLL+foz5q18iH+tOcW4WRLly2g+wtVLiSDAusfO0cdwO95jp
ccuJCz5jhpTiXFzOROLhEdkedu2hUsPre65ybf8FATTI70S7LaXK2ILCiLct+5CF
Tq0s0QIHu0Dd3HxSHxvI11wCDxFOJAo0OG4kxDofweIocDoQMBpgAtpb7UsTbZa/
rt/B1CExUOiBj38SW9r8bGKaaxRdZkpKtajXCERnxx3T5I4c01r3++xZ/KbsKrdo
GuQmAQgm4S82+OAOiLos8yQ0riTe5CyrTFzFe34wWx8ZTA8sJdczk89TaFr0LD+0
WJWB43rdMbsKA6kv+P6/R+XeJ8LYQ5F4O95+qXflUk+mroNDJuN8qHzPh+fYSruI
aFbzuzZOZ3vnR1PhRhJLpiXF/UaEU0ZayIFNg5CRlRjKlc9QHUxnRQQRG8XY0CSm
OrxJ4VZWxiepmPYZbsJBH0r5QVI8vhIxLdLXX4Gjhs8sNWmaeBY1CW1qicgBBWMp
4rFmr1w2vC5rfpqhc9qMCYkRhUCIARv/shu7LcN8X9WkNcPWdcjsgpJkh43x3Mq0
qoWlPBWS2smrAgS+OIpaRj+Jxal7lgQkPxAURxM26sD4m3PfAfjrK3e+xc/n2NzL
CMFeUTUMF4xNDSKEJnU7posAfewzaRdclHEWha/detAgWy7ZhHcVbCf059dTuTkm
EG0136ULsVZE8J3ApbDGK0rzcMutLH7s4xbesSBKGeCCEHYg9X4OEqnwMvDivmju
YnFHeXmr3mcIyaIYhOdB9Bm09STfwdFGtdwh3RuBLzO5pRKsMYpd40dzwY/Qqkq9
u7m3XkQVJrlI5TjBJzBbhIAC2mSva3+NwmuLIz/tFxATuG3eNlesl42kJcPcTrml
FSbaFCShmbDYBD2Wu5iOoGPQ83Qxzm58mKJhrg+beNkadKg8dk2bp4gZlwONDaYf
a1wTL0WT9lXkcvTi2l1U7zpOqNpnDkhH5rmao4eTCdVG56jRKtQdSy54RE8x8t0I
iJuqAuWMS64bNhLY5EjdMH7FzeXVjk1JCUjA13lcRFgpGwSHVpxx9DnurDbidZAx
XlZ5JUMh2KdHpmzwZEngb0b9JR2qWEj+TWnML4I99bUnYel8xCWA7L9kfOUeS17W
MKYIC68sSePqK5aDqgDXWsTh3V/JoICaGYYTsjhcbh/9OtKrlQMnxg5oAfi+cKOv
t3ha9bmqKvGgDsWd0qlg4kIRA2s4FHQtacb5rG21zvu3eyehI/zcmkLd/PmVYJPd
ic3WtaKZkPdgGbQXMSDpSI1ErCpaMRcUUrIkrmDYc8PYaNRr0Uf0bQh3jyDiRxGW
kMMl/d0yCT6GjuNNNc5Vohfvrc8+L29RX1nyLW/GaoSsu33tRd4MIDe6W9eNqQtr
265sHd1J7iFMV+J3KwRzbbMjpkRd+JMQcxheQPBS6IuUXwoaJLBL/JM68UTFQ7Cd
hRVbegT81IbTGbQWDgmIYmF6gfzlG6A7CxAFECpo7ZDzW1M2wYIahZiYhyNA4qBH
5cn9PzJTU9v/cahnQjUMDgjika6aAhcLcHeno4r9QI9DvXJXomyFlXvlt2JwdYE7
k1ZFoLnAfWUNE+6/7ZfEeTNhUjRthY4K9E15sWLamcrnYHvgBMzL3fD17AlKTtlm
8X3WAET+mkbfdWWITGYjkrtG/4qZIEMFegwwj21EZ7eokxXdEkFKCQLeHRKkOhgV
3gwOo64VPUK6UOnnA51DeM1ZPVz6y2Ge/31ZcEIEH/rn2iazoXdm9VHeToqy729G
lSFL4oSpbco/UnkumSq4z4ntLTLjQ10/Trzkt3eJkdqkSnBeGUJ6rjHPooh0ENcF
GzHOwFaCi6P/fQXkjtvBL1quSVnHXZWTVYODvc9AO0sdg4rn/bC4pefFR7eEaq/8
WiYxLTwhnBqz1uKm6ZyGtOjkgd79xs12GXeC85hQh7rRdsKjIoRgiqRzGPk/82MR
Cu0Z6C1Fludcc5J160DhaCTpNYV4y2ra61wD7vbhAa/6qTx/ZkKbCJadFNZ5LcFr
La0XL7/f1goesbreDBzHJ2YcHQNJnziuFjb/y57mFIPt2SpoNodVGxS9qpod35EN
Y3IKe/+SLWPolRkfaK0Z8kBY7etSRpP9W8tQg3xX5C0YLlAOChAOP7QIJhmIN2CD
45qYKU39WvGAE9i1+G0AFp+rRgGN47kXAm+99q4JIofP0jPPLfOv72v1T5lujHYe
nY/R0/UkM34mtjnDn46PnIR4LhBDC7lJGNgyvoWwffUY37o7hbacHbR1mkWsjjDz
6pk2ePpKeAYhO074oZSIfIFyafH1RtBS8WARnnvpw7FqJ0PUjKZngqZ3/3gN3nDw
5DWFT0FuPzyKbdkLc16ZnePeQKsPEPsr/UD4GSuU5PD9AVhdXdApis5Le/y1lWze
PdcV5O29B9rN+fBt6PCKUiZJfoSGgZn30Sa2ayFAE78PKQ7j5pDf0lSxAe/BC2lN
A0cW6OXXDoEMyD6AfH4y20/7HEbJcZ5mGEXktwrpZlt/I6RCOTiut/ZB57Djn9Qu
iZYAwhYwJ8pGDt6g8lFMMDANAtp7GKIvgxqNH8UOUAhjl13X+9D/iIVU2mYmKsp5
KAlc7BF+e1ORQBlP9QCk0G0Lgu1rH1dg+IvNJzw5q2eHatFVij35W6KxRsJnF6Q1
4hBqok3QNkMMZE+Gs9a+Iem6US6ZYImP8UkPd0PsirvVL0KPYocawaYSLnTnEFwY
79rLH7DRVd+KzxzMZlkLqJrMmkXpbl2SCjV8YPvmmFzUIyfYl1sDYIOMzQfeW4hH
hKGgwJM70LpV3FGg/AY3826eKaiVFF6K+TTGMoZNE5mv25H2p2l4FkNLX/GTMwap
/gPexZfRd5KPP6IxfM+KpEXW1FlIPyJyWXqcdctsyFdIj9fgAfsXSCA8GMRosgMB
Kgy8serUYmEtysagZtvZfVdbNVdlm81bS7e8/yKsmM/QcwmmhbkZHOzAH9Od93ld
GtKhd/MUz5FKwN84f9nlBfTUxjYn8Vuogy0prAitdTYCeWmgEWqSvu2O2pmgmJDQ
EI7u0I0LotutHqGgYIsBI4pvdUTQ0YCDkKO0x9t2QZv7PAdN7AlEj1qY8g3BHF1q
a2y21j8fdGZBR41oQeywJKgQDbUVrXoA9OB6x6Eu/v6euU8TAcxMKqncA7FKYSiI
2Kjmka5s4TY78GcbdhG4ATBuRczHxbs5DKUX2+qz3MLJFUc5f1SYaLi3hEKaCDCz
+pe0hhjM6YuC9IwZyVFpE8NZeImBF5lB1JEMxbblQsOUyU29JwuLWqgttrDeJYuB
ZJNlwCHf0bliENSMBfo+cjnjhcoGN/cAyKCPUAUANaQJ/8jt4tEEnLlHzchUBNJC
bOlBLfaMCnfyJea6E42DmguCWuBF6e86RcXY9oxjKvOHyL8ih8w8udKh5i90/Bgz
Ff6Q4Wykeq3pGl+RzoFTuaAzWTX0wi4wmcSkzLWMFSbv30htPFnCayxOSi8LV4gf
4LA1DX296AF5OnpMR5fGcln4ab1HdK8Gas/uXnLuwUr1eGPWAbPtahGLo/Yxjv0m
H1d2/JAWIWQZFm/C8UHfYC1ycK32EPgU6fIFEpzuz42b0ltYljdq+TuyOjcqwmVa
22tRuvlMSzfr8vOw9YMrNfB4J1DVGXknBFxwKU3ZVCGh/QAsos/8eeJ0JyIaDj7z
YqZP94CwZvXwSrqMAqG2KuHK7cokkBn6F6R91JIoF9h1remC9m7aaglQS9nPu9Q4
sbJiNcXlDoi32vTNlTJjY/0MOymk4pcIeuwI5zjIp366GhQSNWnejdpylz/n/LtF
OwYxPYZQ72BmAbO2koNbqorE8tmHTTy/OOqFW5L+dLHJFzisbkOctd3BwkltFc1i
uopDoV8aMnFeC9ql/+/lIdAx7KiUCWBxVddv3ViqAWF2olYpqHSezZJml83uIlBs
/MJ7dvmpsro9q3buNZjU17FYkCyLqR4GHrQdmQ5sRiTNl+91pIAFha/epOGi84Er
3PbUsRWZ0MONnjGdSZfcKjVNMJlBA21oAyDdwr8lvU+Jp16Q9yAn2i8LH2eAHQAU
5FY8ICE5foWs3YEXMwdn8ZxXw5bFaykUC8n1tTKu0xt2aMaSbRRIK/+FM7y2EKR6
OstIbpkKeyNpFR1d1TFO9Ep39LQyIMS60LkjRV7jc17zN/0sDjWbqViXsrP0NigV
GahzxT+KWwymzjHXHjsyY/NzgPf0feu1JKyy2/mg9nJxVVypwj0XxP7GfSeo68vP
QC7qNg8YsQGpjK92qrFz033bYR6SDXMzEemdknIXzYQFBBNtH/DkxzcR6Pm7sWmg
b71t2iE3lghwCJJ36nwLDEpJYSnLWDsfNc2ufqWB2YuIfkvhCxRKIX1a6JkU8GFY
PvpqUPJKLKj/rV5KsJjCTF+E92xadeR3PjwzZTeYsZRNFn35sN9I7hwTCxWjGBUG
sBmKoKiDrvr8sVB5GQLbHohBanb8YbvJTyQbiQaUDbzxzc2DN3fvQmAq5dzEib5M
YJ6il0rk7WsGCr+ErxbWmcUe4XNPwC6JtgxuY6OcM4/4nTlbOrb7j5TzlOUdGmyK
2k5H05bw5zVbHT+AxoI67cnJKWxS2SuLA8EcFAyp7blzrq7guGYJfQFtch53sINA
Epei2pUD0En1SDASSx8qecnbUgpiVi0ibIhZAsYDSn+Pfu2MPkiJK6ttu6Gv3u5M
TEE0XJTdlz1SEJSpH/34kpM6xPAEnGVKWsQIXeCoLm7T3kzcf1QQR0zcSsNYbeEu
+zb9bNvNeF1/WtUpYL2kzFZG/+P3BKM9SFcJn+ecQ7Xnk+XmPXZZl6lRa+dWTNbW
J/bXQiejE2jixyH3KmKnY9qxvQYqTqUhgvGRnYtqsYkdU312nUoJYckiRJbH3YiE
KKQBeiL75RzD//a1Hxyr+WVahPUEkR1HTVBhrQ9toMhRx/mHhjApGXDMrD742/xq
uwEf0OY1Wvyzekfw8Zdznr0xJCHicT5JDm6H3nIOkesXUZIk2Zs9WQqZhf4wpYqR
8nk3auLEJ9DV2grvTljzw8GYtMCpyOnGRm3l2NYmRjKQH0GQ2O5q8nROWi4x6+0L
/mw3FxHmoIzJBkkANLKgI2fmFeYk7TJXgC/F7oyE9/mQskP//S602tn3wONnBiyC
MlpRVdyhlkpdScTbYaEH+VyXEdjZ96tZSiDekmtztKlNPiBE+2hvF3NQpX10KlF1
mDpsr1bofr7OTdY2d6FEexrQZIxg/zMrlnGlKlNmuTXCdPSaycU1uK4p7tSxDm5W
7hPqfVOiT2xo3Lfqrof02p22udoCVEae5IDYoG0myp1lmh2TAJjNR1j32lO3Q8A5
J0c0xd/8JPpt8aSAZ3bUOQ0517io1dhMli7IPHki8E+hOa2QPpgscCwlXBllLC/J
VUfa2B7h3naNtAOJPHzpDwVxfEhWskqhYnOT+PzrX2RABm3anRUAfnUl/bp8g37u
FQnN82ikiBE9sd/oosU8RSLHxUX1ByBW4StVMCKQlAVAU6bBiKoxmDzim2ZQbNQF
7v2Ezr4K2fkkyYWCfWBV05eHVb0gK10sr8M7B/rv9WlGrY12qpWDoIbOzmIvdqPE
Q2IU8OtxJ+ZHYAmg28pKHHOvsIBYzEla6vrtNd79AUjUtYIXR2zxQfiXBlctoih2
jdm6gf6Qqz3nxtoGJaJRF+grR34+QB6K5i83NmBUAlnXPKPPDkuUoWjkIvcCjPXK
AVVsGqwNlUDAxvOBEjZEREFQa21DdQG99QlyIWhD2cUAtolnTO+eHM/sOrN8Xudc
aOmKVFBppnOwzlQ86O6uEJwA8GP9SR1PVPmqYt8LpA7E8D/nqWaHEyCumRcAiGdX
xS7eOirgdVGuWu1PelBJsewWBE9TWIHWuBFnFFrfIOUC5lhyG/sEYPkfT5guARGu
bGp0OMZYorxCJdQotrBTbgW0LiTGatOqyVt3yhQ85mjQjzmyW2A+D41MHhVS9oO4
KpxZBXpILP8hxfVDtAQK9kiA/THmi2n+LJtsUQj/9x4ZxuNJpkigUIbhFaKPUXLj
HQwkKfdMCCXhKT+yH2VzZzeQqjdy1qhjURVNqOqZwgRy1gJnYlsCOy2a1GQDFBkp
yiyiE5ZvVg8Yh+NQdCUrSDKfRbcf+mjL0Ff6mc2edkdFzc9zGixf7L0mfPBXuy9l
UVc4Ie3Jt93CPCk/Ab7jvqDCI7qITrTRzngNAA4RYKqc94GlZLfRLAvJ3D6zDT7g
1TAst1wch0MAyRsY+uPfgplMjl1iPa6TG+oXrvlNCjb9YIGq2Q+5DTRVNU+KX9rR
eDoFSGSZo2TjImVSvluMZpf7b15rhEVPK7b6N3z/oZNqQCig5WGgie8DuN6Wz4Ma
410/pJnt2ZNwjTLMzNsJcWvoqtEVypyOBauf7297t8yuqBpHbWIlYBcBYf95lsa7
2o46VZy7QMBqfTI+7mcWq5izbGY9tdfBpIIg9IqXKhxraEN2Ts+3+2jiBBjC4FYC
Ss+HbT7wrL2yOsImgX/7SPIfsF4ofxL9v/w4/5u6tF9AY8YM1b9McbQtWJigljMM
fu+a8nt+PbZ6WChOAlX1Oq/iYOSLQwvM9r5Fky26EDuB3RXYfMjl4Xv7RU1I1VKi
c11jsCZuIC7x8IHT8fMKgliFErfxe7zx9c4A/L+xWBwFIkT3Mov32vnIz/PG+6IF
7fnJaSDVgYzGLoxfjZfQBR/u87pQvO3nUHrJuAILZwkEzWkS2H4e0CTVWECA9tq/
wEgf2wnV7SIDuxq7XBNPpol8Kw52/FDg6OZ6zebXB9bU6l9bazeycoOF0v0j0mU+
DW79lmMtxYPa+CJ6GPl1f+zeTpGztlMKG/78zlovrPJXREWMYz/qpc9MZKo1Zq/d
l4a+t56S6bXeI9Ds52oaxAmPPY+Gji72/BshG6gx/FPiw2TDcXfLid11milgD6PK
Z+NY9ktslPlXZyE5PWgSnwrU3EeLKneltIvGObBSUQlz6G1yGH7F0O89w7d6sEsl
yHBF2KEzfRjaDLSKARH6whzvDV37jATWaD+kUsTI3IthI3dThQVeen4a7AWAW509
Kwfh0WPDW3yfEBJpdH1i+C2yc3e1ZimeLUP/OU80QayuI5F5J7MpHHJ+rr2ph4QG
DGJeeXTdRTcFJi+Iraz4EYAI1YZMVMA+MFG1JiUgPJ1dyLJfj3zLV4/LbPacealk
TybRiOOrC9RGA501AVgD8Lrzq/ojvuejK1V/Lp3FjkbcnNb14msRqwH9I5T7UWT/
tPsXojDLq4jqexhmQXMVNiQxfpTpgAGzKvqYFtQbAPcKtqMN7/7p7tHwvAAL/wkN
ks5iEyVHul71zAtpHSw4zugCAjSoiDSo7JR8N0jS2y5SK9/9IpLceqgQUujKqfCa
GEjV8Us6Ba7/NqSnlT26YFMYKwJ5gdkMEVBEJmJs34TE2h7DafuSuUVEyD2kzuH4
i200BWPoFMEoBs08Mo2VsnM8OLjK9uEN83sezS2NZBlMUjIICUv7ExziQeZtxC5g
IctLgxsTnZmQrt6Ff4xqmzO97Q+7H7f9bVz1QnQPW8wRxn1Y8j9C5JX1q7+bbREP
+yr3zCuUkfRf1hag3uGD2RWzS508T6UPGWAwLIFRd/lMUu7K9m1LCvPy5/9l7aEm
NttfpPjh4TURnJfgp1I6NkMsgL6ERmQwU4g4DWvNoluPSZZoZy1zEmLBMIdcGua3
Fl/Z+Wwe1cnmhx7MjWd759C0JkWzrBRZvpbQORsW9Kcr2FCUBg6FSvpp0YKLSCBi
nvc56IKR3x38WgLPiALOVfWzeyG5iAZwkgh6ePWmWUAeyfNFpC/WxcRdW2ecfVcF
gq33cju2uKFSjXOP2frd/wv693N1N40m2heBhJxIROJdRdeh09AETHZwCvuOMZYU
5PhxyEoIJwnKbUMvD4sKZTGXqnJ/MpJXW4oSoH3/C+Ym8qc6oULUHbq02PJmu14D
CKvMeYnIg1eiqErRavfY0vsLhMVfcz+UI9Q2Gl9sftVF0KEXCRqfRKmZY560+kK5
I1DbWf+KdxB9XbkkERacx4PntDSeti71B4mGb5S+O3tfthWtGne5p9qcKsUMJZfl
lvSvt4lKkqccLBEs6HE4bnrIsF7Ows4yrL456Z9VvYQCYHfDiyr2RwfCOWY3E3BB
qRsXcbMgam1wKrQA04B0j9DCWGLferq945jKVVdhIZa98kGC6v+cXDyYpar3vvqo
uBYzpgTC4d4DiUNotCerHQUkU9Oaa7ldgPmPMhjcmQsthu+5FqUKHnWtloLiIdWh
C1kSvQ/1HIOjBqDaNr0HV1htSYo2ouJIDve2QqfSt5dUBP49Feea3vg2Kd7jiPTr
IH5X8FpR4qw6+uTOuSGYYn7LA0yb5EKQEpX6B5BI+QV0Kc/La5IiBmJ1WJjlWR6z
L6JcfySxsOdqVTDKFZdpGD3Oc3tqggmYg/a0Tz+u0CKvBui5bCVMfXZlDJbLgejR
RmDPv8rrdr2dnUssD6FNrr99m1ZfL8yQ5C7VkLEeuXXnbtMsS6Sesg46qxyZMSkU
bcVT1WXxngtiBkIti5iDrj7JKcIhkgnH+MyQ+dshHasBnLwdJeHgjepY1TFKh72Q
EPiD/7l3pQvHeNN7CsFyqWw5zSs2Jo8E71XXFBoR9564Sr6GA6cgnJnMWXu6jy4W
owekGA4R7e6KnJe4/mGpvanqVfKG/63ZDHRrRggAuC71p6Hvfb3N9/v2BVn18866
w4HOOGUoYMo+pbUrVkvYY66A62EGolwjNdYZWmAaim0CC7YjjRO5UjdHaIfA0yb1
NW5tBnAEdgdX8pXxOt6HkI0ofmEIhct3UlFkc2qkWoYTJb6taj9rsTZoolxGMrAU
kSDJDerYXs7PPX5sYRvUd52ALL6Pm0XwvwQhL1HOG6AyvlHpcqX068/WyXhP9McB
RdTzQAIGFRVWWO3hPjDLXvawraPNgU3K3jCLKDyQb2FjVasRiQRkpfV5YXBhPCwo
/o/78eL2f06DvcP0fGbXNUNGAxe3PdqRghMQdgSgOHr+qRAAky3C2IReyNUoq2Z8
VLV1xO7yPUl7/QrrcAW3/LaNBXpJJfddgqhy6muqYY4Xve2jTnEPPcFNFciEE9uE
WhNdTE/t1iVOPWNJ6Sthz64wRcdByGUw/6ggWKEWAA/HCPoaw1DAoRutsCTBuuz4
OjmVzyBPKy9GFlbjWW8ADbbX/TqQ9N7KTyNy1xMYj6tstk5otxSqDVQYzOuYjE88
/YXtuHl2m73VBFCrbGR3OQTWMzkb6XnARISfs35bs7Mj1y5iRl01JO1NnHujZe5Y
Ju1byVXBtNXdHusw9mphE4nWXjvjeYeI4JqsFP4ZodxR4S4giOklJ5rgO8ucIfWf
Rx3g5Sh5pVDGRy+roPQdq0t+KlwLQuUeLcEcjj85sMfNnrPklXkt0Blw0IRsFRmy
mJQfrvFnEyVXrYmmepyyIyKDFuApwatICMoEEfcaQVy8bGInNUZbqNfgaW8yvN46
TvTUh230oowQYzDXbs5n11jud4OGDvbikKkft7nEiFB53T3i851/VdRq+Q5shaXL
2O5ieC0bLDe5MTnwCAlNKsUAiaX1Nwd0QVqoXdS6B+i7M4aJo5y1GU8LjtFFsL1k
tx6Lll7VUm8Q0IwswcK+ZGH+OUkBbaEIm/q3EKWmZF3hse1UKqTgQq3AEBtvmkJ0
fAEECY5ih6qfrpM22WvcT/hg1hApHsuR8ZHEYv3KERoYzId/rDIRN3OJufXc7jor
Il8VCJvVPZHtjvFG1gH5jI7mz0unDDSFZpCa1QamKvAsjLB0Czlvpu/lDG6+WdfO
bquVgM+idK5ejr/kDcUVbRvhbNTXrGa80QnkQUH5Qo4jPYP6WGStdtGpxszepe7W
Eaj2leTPaaQUwt77Vk0GzeucQCVQPIezMbPig/fzAsnXiTewbXNrFo+H/n8ZGeEm
Y/V6VUEstgcVz+8jr1tJfYYG6ZGwZoTZYCmzVIiyM4RqCIuqydjCyL/Paezb5lxP
MxAhHiGt2bJGFFWv4JUstevViwY6DOmPd2NEqZSiNDNmGWmQweQkH033A/1ICjLa
2WSftyGYdtOSm9E8N5PuvlxF0zUovIIxNPVeK2p/6cWACDR4kYWSJB+02M0FenzN
Vbn9sHwifavuUDhcf5PxffoOV7DwGc9Cf/myHjqjxpBNdd2ceUISrgnYzEnrliIK
DYntiiTCmerX5cU0hAcGTNAONHRaKh/aWl5A82ddGBoRTNZYZL7LJj+7Jz12wBkf
Q4L4uHkhHbrdq7eqnISTDWwrfBQrfU/sSMOHVfcaP2XsagABaB3vE7sIbPCoOR+Y
HsPP8f+TcmGvVBUn7f2ZTWb9An30Q/dA+/yjJ93cq+NQmf5Z1hh56LLY9k/gxyqv
8o87clng+W/DZZptIdKnyztloEFzDhf827xAYBIyUEaae3HbueB2lv6vaW7dpKxW
C9sRMWOEwfqv62OoMGxPe0dvj5QsZq4fWGXyVn7UtytgRyxm1Dqyyl+AO0DJJIax
17MHjajdDuDOmyS3tPS1LVeF5zOvC4v9aMj2wn9FBOoIDGVRPJiImzbL0NdEl5If
IIawXo6YFob5C81oJ4j8KgJ47mCmNESvaGEIQvU9QKI/ZTK4aCE1rSRojx7yA6Q4
fH8w5wlhlBVILLSSZN1B6sGtnbQf4wfX7jG7FSiMMjfUSfoM7HxwS3JdJZyV/Uk1
o/L1wD6cRibo2HQGJCsuZB/HwzPdgHSGubhL2TKo/5aafsbsqKKVpNyIBazQIvvw
DOVpnGJ1gcMHIUye/JQB+KR2jg99dQcvkGiBpOzlDp4ZUtwy/j2IEL8TQtvYGV/8
9mCbLtEc9ojRC/pWgWcaWetopqgRIJySWO6I2LBCIMRjEb7PjRQAYN+NoOggdRag
I27pDx7sQpr2GHMrIzcPyY8Vzj6AqVZYNQf2CxcebDr/BfVcKaGy8HxldnbBBLFj
KJWYgYz/DC69JnSMaNBneKzmRS/laHRbWt/EQugX++Vxwo9iXyggYiOGnRmz8Zeg
0iS0pWGBBfkOkFG1x9mGG2ijLk0d8s4RrqwtMd9c6Jsov7wSxWJLIPdlVBcVSf5k
dpASROidXbMhsWriAnTmAneMxNPNIFnS+O3A7mr9/EL3oHwFBZuPx0eZYVy75asj
7ddhrOEUNikJt3vv68TIxIA3cshlsRsfrsptxZ6xwCzIieejUhplmFSgxRKdyIdq
/Ey+9p56CDtuOviG2D9/OFhDfb7B/Ly4q2JZ8i5zjbF4CKl1SDkH8b07XYqobAoK
Dyh+eJIcvU9uodpSusQV9g0Il9l+x6rLj0WFxCIB7ew7IYqwswMo5RyH6LHGg5EG
1u8P++LkoxThLA0Iqk6dJPgl1TiWw+x58ltqnOlz7qPWdpM5Wp9XmPX/qUV+5b8P
3n2sFUuWYES9wHKHEoi/jTvIjNyp1bNejCI2EWhOfQQn8qv/k+Sulk5dtlmzD3dy
QeUnEFsIAGHmlI0Sdgp7B+KkuBIhyCvoQTigbksg4pI1lHRF+iKs8N3sA9iPBgt6
gpAKNwketYsBQTIq8MnWY3gf8AQaIqe3TKrEP/ooC1LWGjWuqBjrOpjI7aC2O7M/
uR6D996XuNDSYrtgG0C8h6Wt8Golt6/HUrvMC6ahJap4zCFqPAkiH/bPTTZI91GA
1oHKJxuziazt3sNp8lL51nA0f3kpI1xWvKqkFtuLb0VDirGoEwhC5oICWb3aq4x0
2gCxKWsr1MTdLh4tba4XKbybpqG+CcuSbsfhWoaQQA3tAWVyMXxfDIePdyWeTLg6
hzgasKL0AyEIwedVYIM6J7Xnl040alrU9skpOVpub59PPDDarKOqsiTNOPjEPNzT
tlVMX0o7I20axgmlgRnREIA73f9ddchCe4n06RYH8/11zUk7uRcit852RETuIOFb
xzfw22OTxHoA6T5l19ACblFu3fBNm0qSKksUblkAyIuzj1fWr7X1psBjRt6NQndU
2ABGrzDx6iFWvooG3IqdwUwoOpM4AONtdruPuM9yyOZk/N/ECpIywkLZ5OHI2kgd
13FQpAi1akBKLztXHCcEPfm5OQ2OmsSuA+8b5jezIbDgrP2bX0KIexlUd+oGUKtE
gXJnFtXlvTyJ7REW3MzV9CSOcswSAGEOVCj8OdqXPXP0EkTxPVKlB128/1EdgMWL
af8U3MeQkRLxSScO/iysLOqm90G1uNL5PwuBH5FMSJ5W9BM/EbDGw6ChOs2gkCv5
Md2R4DSlNawxuoSyCQXrhXZTEGY+kaZ2X+J7kpfJDZ8gPW1MkIRVSQRmU9Bx95qp
rvO+OxMhFJJ/fZDGQohdKxbDAyO362naIwx8ONWRYLhICPgQPBr1XEKyqxDRNLoP
qhpIXVaINhlCjocBtsGuWywbRDpnIkv9BRiEa/LIXkXxoEq9fLpPI2yUNXdnKE76
QRAeY/gmbKgPdGu2TOFrJD4tKG/gQlQ2RFOnSMn68n5LKPyF4PXHaK5zku2HIlQa
C7aFM7AfbrBZtD88Z5RagrIST5h4I0QKNdrPWJsi09FLilkT8HNmrAjLZcR1eLmo
kz9IwkudO72Cs7e+onANCMWEp+e5gvSbRnZ4/dEEazvekKB4+zu2yhER44fSzNy2
B4+gBitHF7iZZS12Rki3J+2ial3uISMypy61n/r0urB8k8+1YJWIi1TLGgODOZNv
60coJjyztX2ZYSlE2UFTsnrJg3miLHmPGTcZt26QhLkDzJXVNiBjOBMsqEBLwBzg
dQpBvE7Z+O3QW/n3vrsQmfIMmyI+iRmYF7vG5bO4jaUco15lFkKGrdgMa9T8o5QS
9gc2vrND56QommUJyVNCv7OKI8hD9pHVh1IO2hWneuJsPGG3EKe0f1GvVvpx1ocY
ZwQv/xTDwqXDWf7v/sy8WRK1wGHPVPsfzsH6xVJWJKS+4xL272t7FYkaRjirmxrm
gJq1Rr/LhxfXU3pYWIqiS71WgXfVwqfmCVP7wzJZsUzPUQqOY2PfWhNFJRJCdVfQ
WtFdVAFnjVngiV6FPidu/AT9vN5O/c7Gn36h/VVfcs9wNLiXJysLfE8Xaj4Z9s73
6qAltL1i6tF5RXy7arzITlwgNreQs3kGHY4xpP7RO+Eo/ytn9aAXlEpjs7PDf5HU
Vfi5yc+BX79s8INLZPisyvzeCqHrIeKpAl3TmlNkbhg5kI8yhL3kh2Pt+aKzBUta
Uri97bisgxaNKE7HdKWtvtDeEweqaH0kI1rmlkF95pYIKarvN0TVq9iOPOJWAYdn
MybckGd6TcvUikC05XBLHXYiw/PN9a4ZGQm3Cif2lVAMBeOsrizvRddjObbiCeDq
iPQ7tt6bwLkwy2CdR9HesOpcpKFwJpzB+mOw934jLZDnCl09+Fwdb5T3ei8omqbc
R1obqhMX3ejHYpDkA/EUp+EO7OOuf3RQexWYopc/wEExBNVQO232NMKqBuctBnt6
MXHXO+IR9INfueRmVydv0WrivUq+rXrey0SeXF0OdUsCRbxhSGuy2kxU771nJ4Rw
BF4TxR2aSX7YUVaQOUrC/m9Oocg3QTGFx9QyeN/xFAmAlScMZyTy5M655sh4q53Z
gzI/qFGJTnO7tLqK0jLFEvGDZmM43c3YEGU/n8ufGOGLMRuSvAOins65N/79Zi3f
YrgCgKbbHnPxA29tSVTR5u65e3DnkfNsQiLv/GkpPANiEN6WXjnNnAvXxN9gTcCL
fhGQIOKvEFt1/3J4qm0p/XONQh51/TOgsj46VSrCGZQcbp3yL+zhx60x+3WRYADE
+WCA3Bo1yVHsWp2Upx79o04It+BEt7TPBXGwxuv0mi7pcrn5VAFMSdRB6vuiuEmx
UOxnCwFWXH8LacH6gsSGwgS521bD1O6ss6I+mWK3x6oclNtEiaFv7no179DzL8Id
OPXEUTvXRuCfN+YwsCLQRS38SuFv+6LBMGz7OoHkY1Zt8Da3qtIAfvRKuBp7GdUp
9i/8sldrfc37+JesR7vN5QwMMq/lcfgQooBfG+28WJF8A7lG0UofFOZ4VAurctOz
5JN0gsNZhNgyqN2oOJEHkSwRmyeFcGhV+C4u3cyZOhulE17cGJmbzgY9XCKAgMpS
Gk1R5ncFclzgqCAQGOYyUJ3cY3wUh0BpX06N9vZGsz6U7EvE+hoyHIJMILOHNyvD
wqzzIR+9FPFamShsV5Z+muk5dCIxNzV20+55APx+I4VYTvkXvX6bnBDALLQ67b+p
U53vFFEcOE1cldjRLmJ4EaE/8zL+YDN/46rdnjzpt/PT07LIUcjVWyO5d0IFSkZN
oYdeLKuekn0I/ZPuHNjyAMmtVX6H21CHKEQIR+OcOEAOl7jzzDTw7VqBoimpA1dF
G7VYFjEgKU6eHuzflDr5qwY+m6SbZCGKZcRRhaDghQ9VKDh8dyYdYWc+JQduWXJg
k96QulJ8x1g1WBy8FMd4pAp8n9keBkGN82673wEziyCZjt2b7mz6M35wA8z8jXvD
J4qiUJNR6TZvn7Nomar0qAeWFfXSTifnDaR/L4mJOAm4q2I02iecuUWWLzScbFn2
8OB1uEqE2c7iccElfMEaqgttDlw2C/carJdh4KopnkNEsOzRifKWxt1hUUSy9xBj
3ySreTlmzHD2azHxWYec9/H1qwgiDzs5Pujd7HQSoY8MhmZaVxEIXfcno/0kDXcn
HY+8w05cfvLpVZDhisVWZ5cRZji36ZvmpMcLEH4JM8PWe0Bs9R8eOwwqessgBmSj
pJv3k68ev29vCb5o8vzbayG+W/mLgMOwkG4eylQu3nPS+Avr2fe6+lxcPw8XZEkV
L3SW5PLB8iJtsvO5GkKuIBKQa/l4/fiI57/E91Z1jtqyGwQdkGIDS/ubmjZ47K4k
qHR4dL7Qb6jw7CCU9+Sk4M0xn6Zf+zJritad6bGiRce4zHZxp7hwpar4Cc3MI4LS
5fydOH7hDnGjuFrKkUgESoXh3iqyw+plk2lpVihDabaR0rKccPF6T2dHDNGagllv
C3kM7k4DpzfT3jQbQj8Dy9sK5fXZMlo3sYoWrA6Jxh10CXNz1scZ2NtEOh9jir2g
OWa+yHP/lrggqNgdPsCU5nkGTPCAgT/VnHAyByLpsX7OE62wfbj2S8k3+M1aK+rK
p4z9fd/Fiew7QH0ms1x9OWDVjmDtoO+WrmrLzpiDcW3ErS/V7lVWiC685WjVWNSi
LWKs/ALsxDLUTQPPjUfEX4u4TlaV9k1sRD20N/4cCoAsT7mXnLYLFRhQ7ogCnt9V
LK4eDkoOOKUJHf0FC+QeqNTC9xYGJZgaW4+bzcrP1wuEytBQmCCAtxUqWQkH0UCk
uqgG66geBkiQeKLrh/Y0FhewlXy1oSeXdK+iu9Z5Yw5FVv52ks/MD2rTItyC15Rw
pNHhILYeu9o6R5EVAXousJZ7b1dsSSxaFwFQ1jCJM0DRylXYSWquJ3ptxrPJsAHG
7XyuYL+2yYWaNXRZ6q0Io+TDGPhRKysT6gOcSlN2Il8VkM4PBRXjyLxMnBKRM0Ln
Bw99Sd270cKNIquuFBM+7mavJBrzWZa+Q517D2Q9UvC+T4rFUns+L4yQ03wbV1EM
CadONIPTyU+CVQTy7jLNfKgaGRVrhUETFo0FLmnscTnUiMVq2npVcV/wfWckXhIB
Mx96ixfFgoCh7qQ032pWusyVuM5JXSe8UzBaWvS0cRP/H7XtbEgochDas9vQt4YR
jbVIQqinuRR1Rh4R96UKnu3c7DyaJzUzIi4L1QHKdbJVuiPSvU4d2ZWZOLIk7ysh
cjSSyiMDABkGALGYTzW0NezRuO0Qkjq2FpdgWT9nPBQ+i//NnRY2tFQxaxqNpzQ6
BYd9jcMLvkXJB3GF1axmwfnwBbRYSC0e2DB0bkcytJpwhgBz+Pq1Ib+PL7aKFzZj
nYsuLYYIylZIylrKnv/Z3NDnTohztzzXeaKwSPEOu9AK6MM5sp5uRMGafsgs1+14
vHaTMdmudVSKq5FZTrbllbd+Xj8DC4GcVSupix7mTogJq5oAyKauBh620JTz8GSo
ZvMn2+Qn4TrqlLHwJqk52H3XztSpyE5HMfTrMGKWtNMs7kmRitPeeNZZ49O6kiza
DNmDrKnVsG1MmotYjqa+dWAy++272aAuz+ZFvkOvjvP/voRDJGpmup0OQTwG9K0A
3DkBhcCXhDlmYUa9ZFe9oGNRwM17f4Jl5TWOMLr1Rm/OoDnRncO+Vhb/psi7JAmx
15d0AVjFXc5TG5garqVDbNcQTHj8yPAVo8UkbiOJppSu9wUQVzSkdP3704AoQeoT
ZSO47o9A1MX3qs7J/BQjHZ+Eh+ROtH/4PlojihiaH84obZbrieIPoP/8h9FWQUxO
q4aea0RNVkhaeXtA7A0M2FCsCHHOkm4C0RnQRGIag6j8VX3Tw8tWVl+A51nfPIg8
6O6hfZlRxY8/Skc3cedt7oOXsoWFgkIawn1Lrgw66Z3M+QaLWtF1IuOjtVIeCFRD
c5LWtVxgX3XWTMKLUCUW04w7JHyVgZkPP+X7UHbeub2hQmcvD6FbL9QIVg85T8gK
hB0I/tJ/ELBynJI6PdsBcxaNUsfyK2Bc6t/5PbWPpYQ/hEig5Ql+SDD19iwVq5WW
QFq8YW3ONuLjkPMU05uJrZJjEWSJmg1lDi7x2Uc09dqb1P4cBRJQWFnMwL39dMPI
Do9Z5GhxVM8S2HwQHH5DFkkjKGQ3HRj21GZInMPoLc1BncLzOW7U2/FlHtREnOXr
R4uxGNj9opgtPBJULneaf9ACludrG4POlTTvEPCrgY2Gzz1jnLKjb5WqnIoND1a5
0b546XF0mTDFQzZBks6Af1PiTZbOjIxvBksiK8S3kIdMYMgyYtuHWhVu8bmEPooQ
csRwKVzCetjnfwI+7AxmCq4ykCNj8QXkKCUUT9sizgZoKBXoawr7OioG+85HQNMz
dy1vLSPOQ5gzobPVzSE0R/YQOdy8/heJTyOLfnlGfOSsYJoxQ+OC0P4KcR65XPsF
VYPj5iwcaqtEPT9p9cBwzPZ66LR8DLbHgIOzjOwJAUVgpACkXTdZJJWlkzFjl5tg
o8M3MVjcBynz51C/G+TWjvSj3HaU0d8BunjkE/czTw2Ww4W+nzmuKStpRNUosuaB
fzlZTZCCbC1iXByaggOcAxz+Syx/olVQ/0a2Ta/szO037QI2po7BDyDsJMrIcjX/
DX+TR0WF7Gj/JTWLJJIXH8Pdl/gVRbEf2HEnmrkLm5xdcRQF8J7exNN+cl+uIJvO
Q+q50rFpwPV2NiS1IiBqJdWkuUCXStOoGbMOXENa7dPEhiktWiOT6YXrU+/mKlEX
olofe18ijAZOj/ei48HonktkMPJNgN9I8f3FOCHhJinLmYBL8RoJlGmL4dcWvcZY
U6IAANgmKDx917CpeM1esXQgku9Su+XYzsS6DJWc/BEI5ojLQnCmRZ58Pcvy9iME
QIxt2NWdRhTN9RvBGAwyO8CFGPV2d+U8SXDb+KWUjOVMG2S84U6HFDsspHVLVdKW
EXPmcTelZcXbpi3zR+kf6c1rNnvaWl/O7H5rLGUPKiQWeuz1OAvqwzqpe+QbM4bN
otA9m8XLclnx5T2Wahfy8eQFDnEaP+FYpJ9L16aJ6brpMLH+JkaL3yhAzSsgJtrh
291IJdU3YqL/hKVVNaUmssQXnjlpd4tiGZfxk4oWBTJP7BJ9l4BuEsmapkQ4gnvY
6zdVX57UPT+3QkAZhma5+GWH8L5Ca99cm5YP6mNN6CvgbzLugc5Xd2G0+AntE4JA
IHKklNR/+6EHQrG3x0GzWp7MrnkxHym9o9lcn138LS39HBs5TwKD6EC+PHvtiiHY
e4Le2kWIosq1kOnEiQfAmXBJEbJB1M2FvoDTDRuZ7bWwlYViOuupJHJnMGa+RaKD
jvXrMeqQHKTPCULoyeC9GuR7iHUQNSNvml3+WeGBEVplUObMRAf6ihRgEWqUvFwy
c31PNR1xLovF4bJ9MgQv/MSfu4l+Y/VZv+fbuh40ZUmhHw9un9ARW8Q+7sxYblnD
vhAqAC7LedvN9/9Lcbhwttf4R44fk1PrZSUtRqPIZvqWOk/PGumoT1a7j5MrvhT6
/UeWGg5CchRBXXrH6NnM4SqLSJARlbAfKoc7kTppT+DrBOdNz8A39BidJZ8Ke4qD
entIOFNVRaj/TiGQokACI7zl50k3QHUm8lQRT4roCkI83HZR3gjcxakLYCPH/Ohh
EvQl6hGYP9/FPV/WYQ3QBGhf/AcGhJ2I8UKMYAfEXSNwB1mnOYL5K3YtyyK8YBND
F3sJ5HZcR69Zgs05cpK/4NEazbC+fjy6FuvNXmqegRJ47b7e9bl+wn4F28Tq+c9c
1Rp2FVXZzZEt/vykbBWn4hC82dv9SzG82aqY4BXdYfTgqf87t1wcGunQLIqMrsCL
oWRfbR3ow8zMLaN5QPLrZpjR33ghQAc/yA5QDZB/4qfjh8aO+iUAjifWiknla3XJ
dRwtlEjl96Aj2chDEL0fq8lkcD5rb2j11VPfbHbPrY9dv5/nkYkGcyvLihD6em4s
qL57X8NbJpAu7Nr1ToM7jITdzPp8rW3emIvi4aZpkb6yqzc0scheAJCeMg7jGWLG
emZfGv7Z4s3wvMmLz9HAlC1EP82tBSZsVvVenof/Urgh+g4k2mPk7k0K+W8l4Pv5
cclCWNPq8GEZTIyPML9r69gjuUsMG19v2FCD6nsrz7S90pkxABxP0bvQGE84ZB3s
4TNGkN4xGagD7s3Tt2awefuCzhEV84yAlllzqON5qPnepI4D1UNFo8JO57qYVu70
LWeqtUYiG1f93AGWvbwMS0M/iwdmRQ9PVpn2ykid7rR/Gt0/z4447o/pt95cKXmt
4MYGuzzQknsI8j06LFLqpDZpilEya7Dp69okM+rq4M/AGLr4bLfAkvqzpzOo94hq
6Ospqgv7sgoFJQJFntlu1G16FfWYuFEWFJ9Gg6iLRcMmSDDSH8Oqktazt5Q7g7z3
9pIVDnGnaw5zmj4CtHthGFgRIQmSq+uwvsSAA481/J0BgjaTlCuQCI547ZFts60s
XAqAsR4mh27oZSt/XHc7eLbl0cLuhRb7RGCRZgJEbZQL3YdDdjHcQjh1K/hN56gG
t7S/OXihFHcHn7UYJUgtrDGBQ2hFoDJPYiE4MKPR8+pj+X6m1JWuMWrJW+iIwOs4
jj71T6Qjcq5blHLtvlDJmioTXT2zctX6Vk/izW6z9NPcXYUIjdJaunO5f0YX7Vfv
r4oaPOG9M0CMGY0hP9vIfFtGHy2YoFiCKJAMb8sIlYQMLxBLfY/0h0iZOcEsdkDF
yFfcLQFZEjdLXjfMEQ1pB+vUug1KoSjWdGzVFXEGKw53XJu0golcD9qymBx7WhQ/
VF1jOyAHZ1JDPo8h4tKYLoJSnDNDdkX509QsQdyns+gs2wtAET/TAVp67xypjrvS
qEJKoigt9kyQlJbpJDN88zktpb6wO4K7KmYwhYyFmHKsy58zVMa89QzE/0HC8HgP
haOLpKaQ8ykRD/XKAXCVj79g9riuBzFAGV092tmyhQh7DLcOm9JzrKolo0mjWk5j
xRDzJYDjzXQe+i4jarnvwb1CZWe2gObUj3vO4Qew8LJr7jh8FqtfEq66Bi2lgFpU
Mnmx9dE/+JK2eEh4ErW/hegq3MHqzzOkezh2sAMuTTcqpqpHa8DjPNXPl38PSKjp
Ljq5DsI+zbg2yf6pqJD0TMm/AvjsuSef5Jdp2cmwyy8sIjujYkgENR3p3cpQqMTq
nTvViR7SQgpruLS768QQLXa3iKvRD0qalY3vGnqtdzBoa22/ogwol8fEUdN+TwSB
4EWwWpsQqcHsDAWxeiE3YKds7XardGdFIduJfY8LkIHZ2pUdLBG4gsq/d9s6MTKN
ugdUWLkPhq7yyiFUUpWKI52BE5xlIuchHd7k8vj9iHulGkKRP3/6IZwc7cuV6nKZ
BJZvY3uI2aDNFq6PuO7/gZflK7FGSXCCpuzLlBzB4vn1q9QPUK9lWOxh5X53dcwv
06RO7RDavkLBx2O7Q+XOmH17whoFczTK1da9HPLuvFsC9HJtAruloHJzFvhhashO
qwqM5HjMmEyMNAftJ8endE9nGPfDVIhFd8uHzDZGVrRlQom9RooEjBi3y4dyd0vm
RbgNJ7EwaHxkVy2JvSFv9TcljoWb/wZHH6JPM0A2e0UkClxtscNxSN7S+fXwxU+Z
00WXcjOGj/pkdMrIAltsWnCOs60m5D5VWj5a9vDEEH0jK7tpwHzR6OfaMgOj6kCk
M846wtXg8Wa2K4Y69PqBmi4uz2E92Aimn5L5HjlmbVguyUeN3ipaxU5hnOwoNvUi
Y5T2BErM5Cr029AjctExF//oCOZdJWszpzcdikYgK7kMCZz0lwPA5VGXTt8H3TnC
GYB899tZii1hkw3ZAI0tHy94rOUmInilJ1rjVmy/2/D63LSNKHAuEl9CWfpIbbav
DK1uHJM4yvhI+hunbe5ElXstDXJTcGDMGwW7gxnQTSTfDIgRRXXwUKRBSvU+wGB0
EBrI9G8n/YnnqjiBE1HvXxF0tn37wowryg2gb3dOZxYyd7yx5PxKF0HyB/wKqhos
+S3VKhNLlX467DR435PsEXMTyN6r8FMiGXTCVHdDDhuZCVN0ZaC70VG2od4rFejD
Ne8yRb6TZHWkoLqfOhNYejpZDs46tRE+gSglrcWL+Txvb2rJVSzsfVPMh3I/mikl
RUVD/59vO4MaoSny2w0Pv6JtXiw9Fx4n0OXPG23WzLzL+PAdm19Vx+d6TRdLg6uP
rzuQENyewUEStb4M0F2GmvAasfISwYTcMmW6Lpk2ffG/isv+5iWevitdZ2v5B/Wo
fNGatLieo+kqGiPGwe0ea5v+0GfPBfEJ55WPfFjCY6VoRer86pRJum6w04z/Ext4
AyIzeCr8aDnx8j5sn8gqltPNO4YbnBopCwcevZdBbmB2ggHV4NNOb1LRdjXroy5f
upsieOjQIuZmlIOk+Rwnm96fKuVBrO3QT55wRX7f0ctlokz20tERj74sc7HdZ2iF
wIYX8/eKIedvPLQ+jeWEb5pjxxAdiITz+2OL7HBLwD/7svUqrB20GH6fm2Dd4ibE
5OMz+l07CPl4HS0/+r4CQDy5ZefYT4tF6rWpoEeoJEjw3WUWqckdeEcD1zlrbUYI
0og470d6NkFs1x0MtLiJs1wtHqqfbPTJuHa2eCuoIEhFXp/zg3B2tlliwrSNcg2S
vGV5g5xqVQKVDJy8RGsRfV8QxyhZlQffAahSOTUSWF1CwYsuQIVpvYwzUw/ZYwc8
WwYjnmbcfveEBRdiTksjVCxH+JFndzUttixoPGndjXpjSSc8HvEZqAOC3gQmCrqZ
SGNVXv0eqmZo4p1OnV99ASkXRnqXvvCRVyEwvntSFTvFjjqbNCcl1IXmNdLHy7kr
Zmh22qHg0SPv26yaUuh5ArjFCKuNhP32SVa78mUWGiDSE3lhT4s5f8pFjYHm+pcl
6se+fFGiIBsSqxSCrGTlbm9cFrUgvijzGZzHRnMRClhfMZryogK7BevXq1X+G37H
MF7tgujA/5mlNKkZ3TllugB2O2Yy7wgwjPsqRTBkrE4vwjJraK9I9R6smBDC+xmd
RrH3S9LmRDCWDO6Cvdddw9FKcAqeIRSNpch5mJpIjsvU6iqz8TRH9jhM8wOhwXRp
Bm9o+ifpEJwEFSUBIjhyqY+2lzXbW8vAJ1bBCAC9bifUj6T9MKZbJLQs6Mi1NGKi
GmMISdsl7s/wODk7uXUFVl9BHdIh4+z6n+7reMIFbnSW7SNmvEB7pMoHKE3FpYYF
2/YzkWPlIhKsmMT84eECguD8vUUvxKsf/SeS4+e8xsEGkxJ5Fq22EK2gotdYChap
hEkWp3INyLTCTORvh0W+SsXzBIduxkQG4EzK5cfvDmYg7GbLMO9g1O/FrDueAOBB
PmLPhnE1cWYTF3StCIBvKXOVUuqMcP2xnOk9uYYhjhPkUvhi43yAh6CodLyaQHRA
456l1p696UUf8UUs6CPcOwzoB5EiLfcd/WkyqFhy+6GBSMTO5a6BdNzl8VCOgIpj
M1dNEoxcKIRADmtPM5hoAN1fCEXVMW7S7206TsPotqsJDdr4yfmayPcPwq1uwIlp
Wizmz1LF4vsl4DAgEDLp7lGY+nSNyi0yEX26C4K0h1obw0pA2xT5bhTP2e7lmMyW
kzRzBkjCRuiKHTM5z4L0jr7Cn2bC/USrCe4LyDcv8rBMY+7Iqk7IO9Ljy2y3B9dp
QskQkym+dcwIjcTglwal5/+OR38ZfT0/KMO7fA8X3BlpPe6/UPsEn0EurRRnWMt3
RogBGe6OcUMn74V6fHFtC2xiV3eRcZLRduSCAFaoC167gkwmH17DeEBpSw/sqaHt
D5DZkym8xK8h7QgLia7PEUggdUpesMsdkDHAmlFnrhnRvND27iuc6wOLbOZs1w+b
yjTEtZGXpLoMc3RhWXApAPX0A6w54mTU9Tz1/9lOfqrc5bKZFU/Npw6sKM2rf1rf
oGkY4wBlWDJ8WdhYMKvU6FPR6TKnDvM4KNe4RQJLIU4Jt9TXUGILjdFsYU5gGMQ3
UlbdtBSZBgPt9otYONx46f4P856oVjBthfrYlO39P4kVw1dG3sbW0ZYvQqPdvOo+
twkIL6/oIF1obu4MrIYuuqme5/5D8/Ej3EY99i1BaeUE0seaZ0uCfP6zdthkuw8Q
wotklwe7WfvJMRgPIR8qRiGM9MWKC79Ud8y7O8cDQhb9XrxTmE2OsMo6/nXubUX+
+rCeq2CzE4kEZ7kSCQj/ZPQ6OWSV6wZ9hmeUNRN+l6oMm1FiXVM6GmZ3849cWMeC
I3h8p0DGkPU8dRg2QK5U1dBetT3oTheHSlQj+GkvQtArCj+6oMAZhFxRwRBcXVoA
/9tXbxbYxTFmzEd6nJnVjKw5K81vPorjrSw6dvzXw4/aWMhERyKzj9+3qXSgJp/W
vyn1dawDKOv7xDT6XwhDQXk8D+j68MmnT/W7KnZCDzL2ThyaBJkutzWvvjISNXgB
9GXfSvKAIEVnMaXyKQ3Gd1Gp/SLIWH+6oL8E04bLkHEpvxJgsqb2/oO+kAuF+eet
0dpTHmKcdg+V8Kxo4hqMHJkEIBfxrC9q5JQUQEmyH6jAhZAWBLfZboQM/CRu0fvR
tjlE51b1289teZh/0aJXDym1LKCpK1cs0M4SOK4D784y8djiecclL40l7tawez6t
dPaarDfsjAA60wf1E1obhNG866CSK+ZvEeYvRH0A6qnCHMUua1tCtBz+67vojupI
1GgT9mI7NK3XedDFIKRHUnrDaAQCKk6t5a5pJ/E4CcNLU2fZYoI4kOiio27VyXmS
O++PD9lGmmXelJyCelCwpGkM4kFJqZa1OH/t4UcwvQ4jE7w6k+d/IwsOJ8lJg2rK
RbVqbOXm6rNzms7ID2YnJJApEoWoZ0GenzVCUf52MU3y/K4zU44VzWIbKNzr7MzU
lqZnDgxIjOiW2ozX1VLHbbDzPEPDyka/c86xFNnvXTStz4Kfs3cwaK6wIc6ihQxc
1L5S6mq6YATxCjoBuDFf6pHMvOWPcrJ+W5SKXioCr5mmr/aLQuX2Vlm+0YXE+1MU
fnTeEAymjKeTILubRwvAqJmnBxuGgTHmdPQ6t6gBCkCoMTjDziD8gJm5xO6dx/BR
3WXSVCkAYAOfzWmP4YWFNz5WX2gdg8MPOcXEwpnF1IaZDkKtJhTEK3shPTfOXcnl
aQXHu045ITCNpzF/2U+wMdmXHG9AH8NqY6SBXz9RKVa02tsuLhY3MdzzaNkQawYA
o3TCtGh/Jj7WwyM27HnZRmXz5Ak97hDFpMzG5YVERRDralas9aTv5S564yZstAjG
x2EzwUnfPMfwpaofrQRZRe/fqyo3BVqMD228UYb7IxDW2J9RsTcIsBZFoHEWPDIP
u21wyANXEP+VPobbzFkk8Nywa5gvISaJWefdBjY7tVxj2JjGRLx6l+14HU0HUk2T
qVyqAtaTLlKIGNa3EO6UqvS+u0HLSWkfIDpJ97dm2mXp0CVNlY5NFCSMWxY7AZrz
nVlXUa+Mbj6DU0O8SHXFasPPVLj5uvyakak61jV7pWSIAizueRIyc2Qj7FXE9S73
ZG27FaonX+BHxK3N3NwaI1+g0LzTc0j5b0WIGLLzyte7dRdDRXNVJvBQtuCLFf2W
EaewT9nd37IJgFyg6F97fiK7XXZC1s1NaYUGyVILdd47AcBSiONHsrdP3Y7B35kO
tiTLlZ/6IDDowJ18WLog5v8QLLzyqhZ2Bh6VQt336/bPyosUnLAuVY28AFbvcYiC
QEgtRsSydeKpT8Up+9+z7lSg4CHef/f1Zvf45gDg/AxUh0BXVJAPEklA4OIoOlla
Ba8c1mpNYdHioRYDHtsYrjvH8YnTVlhrmuxng5XfYljadO4I8LV8B/pIW/Amne7p
pj98o86umq4SWNkSMCk/dtfANdvvvAPaNC+t/mDYaBhagL3CB+d18yzUTH3xC6zR
7gE4T3AQaVVRj4aP3kkRRWbIeGalBTarc6ei93gwyE0QsCmhSewZGySgnuBp4NX0
5ZYv7BsKyYa90KYX8pUPtWhgJJCSv91khLyjm7g0VTa7uHTghZu3RVwMlzjmy4U5
ZFULNGcxL8lrobzkI+cMtvsNizE2m6R+VdkZQDS5fN56XAZHXZKQ9BKsUF6FMAKV
sUDI9qghyvJOac9fc1brB5JAi/srxDXN/vuRVh0fY6Q2+u02wSx9NwZQB4DMCxzc
6uzSs9KgsSauPnhde7aRivANbrFNCwTUg4hkG8yIud4Ld7VZpX332nNANXDRfFVj
x1xHs7mYbt7p7ifCzpk85wY4UYjodE7iS0E5Fiv3w/Ha6fsoQgeoTg4vedytK8aY
l1HICwahiXZu0j22tIQJkkwQpGKiami9bxytQBWseQzNlB13bSMRmiXFKGoms4Fh
S42WUgsbaHefQYNiBDrSP/pWFqvV+BqY88nGKEjZ7JMbdosBDdQDH5xYhwDn+70d
L7F4AX2N8I9aVyc95197DFVm7MT5hBnRX5PPJhtYGNmRRTVd3E/2VV8m+FrOjmbU
xbWD+N742ylBReqV0ES/w4sxwGK2TLoPKCtmSUTBcjm7P8b88SRePXov8HSKNYwu
OfT06JtvnBd+nFCUMOck3Oc02/qiFhqeCgn5xlSo8qoZACYfNGnkBxfC5KPFWawG
WDvu7LMbLpdRl4Q3PyKDXyQ76c1kQzxw66+I/Odvk//Q8ULDDkiDSyOx+IcdPMh4
m3PmrAgXu1F1mAnCwnVL8obZlhkBYjH87P/Tsc5dqv0aUaV8VUUPdpf/t0BqcMzC
jqw25/dddsBPsebC1zaasPNvIRstHIcW54VKuRjVWcC6m6yMhNrDfnteongSJ4E8
4RtvTHpaNDr2xUcYJIcPjt0FMECiVoqcsWG0yruTWnycxYmiE3raMrp6x1LbtKlR
TNYGNTpswE3hfhj6fAAakWlOL1p5sSD42I1i0g5LhySLD/nLZlxifEkEQevLjsFD
/j6rOJy2WuHTw6qq4dIeqoMgUBFTQE5ZTKbNpQ/WQrL+w4aH9FUDs0PgZ4cqoM5M
eRc36xBhgtaLFufiM2kjBENhitDtiLVtCQVGrfS+NbEgW+eeYybleE2ao89mREZG
t+zY4e/WXoMtMCpMdLhXTZPJVEz6b7seV0rHXpBFwl4oa8uTDU3LlhiFyBplSZZs
l+k1lXcmrQjyhMFxrHYLohBfUjkDUGBjtNPMviCLWZSD02b+nd3rvI3sDmp7TLlb
Z7hMQ9KbEz+kpjQ8GgSYQ0nt1bC7MKg+P1VjIUZUqQa6cstjFhy9/cWHhdqrmi1K
7V2nfWkZi2Mi9hkQDcHqlHKIhstnKl+gBL1bCi5rj6pxVsis20ikGPi4h1tg00i6
NUHzQ50qStzzrcrr1WftDjg+R/bt4PzEeKYpozZKH3JhPkDbWC+w3z+wrdsSXV74
okbgtcx+Da7lLpKhC1LQH2f4G12MTTfO9DOB38rmq5ilr5tWMcpywrr8PrqwL4oU
4jZBtkiPWO8QfKU72yaLNmtjfg3gHBkXwZuj2ZbRzypZnyzMybaK4/kfwqxYWS/n
znI2D4WjqIrbO+r8ULkTFkMimLYW+OG+HIPvnOK62EQxxRaF7/rgWxuckjmnbOIa
zV/U79O0D+EmpuSHKz3J66DRKrfr6K0Mtlv8EuRTFLdGQoMO7RNL98d8pxA4Fe5l
y9EX6TqmuYfs0auCGTJICIEtdqQUmrXjFxTmZygi7odbCPy6awkzUxSqqJrHT9wG
Myzki1loWBHvzVAJTUG9pfi9injdHvHV2ZoyS3bJdARO4L/xzMMmighkA5dZwRN7
EOLlfiHf05TLpV98P2itk49dcEV8ZKj6pY/Zh0WbDb/nXcueHo1Jgg28ehCPJwHZ
+7E0RwovoIHtqfaL649zNtkCuMbIB9HQSYv465avSnCmVn1oC985a3no08HSjtWi
/vZRvyzjcroOv7ZEnRwwVz+RppwKR5Hq2mtRDcOFUcMhtu5f0E7g9fbX+iJeCDWg
3YS7n8wt+CR74lOEgQSmrNphtkHHVSKIf5jKZ138zuE3JXz+x2hcn5c2L7XOyf2P
VU34W2VLiv6/E6HmA3I9l6ROhVMqN0p4t1sO6/8r31C5w9DW/lg+2HM7ZgH0c5jW
JSb9Yo7R0+nTI+85h6zoFmbS1s4C3z4S7ME8ZrsTS2SDlSQlKVXgwdabY1W70k5F
WSLjrPSynNLue7lJ6qFBf3QUnhPqmIgH6lBfnBmyewPbou79Wcm0eNOQELfjaZTI
N6+EkgeBj43SEqvNOUlJZoV8UkddFGEQaLzMvjMB04uN3TpjUUPb3wv8OugM8ogM
huN9xd+aJyUNeJ3+DROiUa+g4e4C9D83kYyYJoTS25M4vKdLMveVve6HfvQWHren
N/Mk1oShzAZXjYh0smbWiwNrpwcKym/8KSsVMEB1uMBWyXD3aGdrLybcNRrrd5+9
6NkoxSPZSWQ0B1tqIC52mB0ujavBv5zNlQngqmsl7UaUQLCLJDvp+lzSXa/WrFAN
UIm/IU9rutaUQYKeYk9dmHGsJUcQMtLiXpXjHMhplTEXB3jYLcL8hpIy7f75z/ic
0RUpSe0hUhtRvRiXrJJKAkCRFrCHb+MtdyrtnwmRdV1A0G45+QCOI4qeBnG0GRqZ
Ribxt7omEZFD0JfTHRIaEaUwIJa4El+aYDqop0PGxVeBIfaH2ExjbC02iZFDbaen
wclMjMBwW9xsLviZA3KEQXNSKOv7mIvvfcUHYNyV3IKLDm4xRCvYZ/Jp9HvA7z2E
+42Es/ZAmfOetQGonRK4wo0CwuegxfoDJY4v+xVgrI3xdqDSbnNmEQTNf9hhdh3X
p3wS3MPgPwPTR7eoQ8+ECQTEjShGOJ7I06Dy8Ir7ZLS/jfD5Hy09WeHd8+vHcFTx
IbnPIrg0BCUMMprGU7LFCOV9QONIra/HbSwD3cUJXkzUXjdGXionqmLKxe7Zqj3O
SG2q32Qn1jweEJVZiHATP2mlGSIZZszFW34j5YAaKzZWtchb853F4FGodXQJX8HA
V5BAcgcPB9wO3Aw8A9iISlF/YNCPkFipy9tECluhxDMT8oKH3Rmy2iQqqnbCOz5l
Tet0QVM7UEuDKGNlaQEbKeEYiulCbC4WZKGe+qBWpW4PPMqvuR8Ss/N/gTiLQY1Y
5272kwBf9QP/L1EiqhYzxWI1BpzIHhUK/7+/qnBG3QS0Od52/Amo4yVqqWK8eKfg
gcejISsI0TlIiC6Lyg7RpY8NMAVJsKfFAdT88pKh9pGBJa2+SH5Ry3aNLRAo2UzT
KKGlVTMzmO0A9WX2nCE87Q67W+jUL2zwbYKLVqPJav05Fv7VkRnxHv5Cr/3HBQxx
CIFhqtCNGstKnMigwl0pYzIJG4lUkQ8x5nFJ66g5EL5K0eHYY/XfkEzX1dlSxfBp
d9CNrYnIa5ygsNUySZnnw4hTitAWsAT+GbYLQpPbTnNj/atqKeIXAq0s1tUIZ19y
AEYh1x4xVDSxTE2q/HfKxR90vKtt20i+eLCeqT76uELBqTRxkT/Jx5KvtroimEuC
CE34XLTzDj4G5dwp/FE8m6+40z0e0DsSorov+RbxoLayF6LBsive/Gd97VdFfKGI
T4wFVyexHkueibU6PkE6UpUY7u+wuEolpMjeBOD8frlgM0eS5zECym5UTr1N9Enc
vINVjSIKFqnfy4GBDBzdIlZ4vEgwqJIbc9VzYX3Ptazt9QDHSZBoparmcCuIkGdF
0l+7EY/1EGVekdvwSLMOnnwsVV20+FdToXdHKBPuBsAKTSdPRXVNV77SN8mt+M6U
9AKGlaMCpFZ1AYIUj8Du4wJ/NDF9ug1Ku018/hDaLrXoPwdQkNBezyt+ckyy/MZF
afjR2i8UctiBNgzL7dCHxINpx5CMmscxBI0++Y0aEE/2ecBUQyXAsGMj4kVcF1DX
FYrkZ1aBOixgQ1bUQn4QSD/Un2pb7MVMUxKqQwRT0e1wWvNsha5huUA3fNoY/rVt
KMZyyOozzU1acAiCT3oi+tuVKvoz43dOOnQsibg7j4U2Y5lJWdWOP65HTQZBXfyn
MLaS/+gbfJB4FLNYimfAZWcBcLt/QCsIU0UiIL2h41mLB2HdU0o4iuMHvXvM4z9l
/JZlZiomVn4VRnyp2rOToCLGfNRTWl8KWWvKQTc+lLWms2GmQRNVmEw7iY6M26DM
KBrxwlZP+FuTaLxIACnrdcyscpg1SG6jFxxsUXw/shnTtz4l08URjniydiUNPehb
jWBkB6KueHY7/HHp5rDjsGP2eFoXh/rpL4SRzzOV/OSS/jXJcI8r9Pl6fey+Zf2L
tq9Q/4TxxF6VLXH9MneUPZapjgFbkPxOH/IEJq5FqwIc38Swd65PI9lSAZmqj4+Y
y/QN13eciWftSB9hXckDegorAR/CY68hcXOXDd7MYakwTc3UVPD8j2HbhPSIAaW0
mE/Eq4K/tcW+cXrqjPGt6bi8tg6WAfSlgF4+wq5zYcbNVOhbN49cpKD700TZaMZT
idWf1rdw8D2sXbD2I8MWBHnUkHKL6SOfGrL8nRJouAmgTFDc5PiDP03saTKamnMe
4vmkRBT+/eLo5W4/T8mzcZ39ZqqzpLNvGi27ubKPZQ8Ica8mF6YAPnkZvVSsz8a+
6LyVn7yj+hFJ4DOBp/9ysA1bi2myLQalf7MNCu6EBUbhdF8dssJv1ui64+T/1c3o
9AIViePPbZeUTbtERpIqgghwpuAnYQmBa1XglHLt1udQ7MsV/JsQyeK9HivbemVF
R+NUZHkSm/YODps9d+qWfT+UAVtWqN8ZPlhFYKpH5+6gDzw5QEJz7QWACMpSx7tZ
grUdzgdEw0R4Eb8Tn6AHFUuEliEgYmyP+g9A6MCcaHtJPLCKuVEpgaHKLLnbI16l
87nUwKDLbmUiX5sv0N2hTeqv8+MC05DvMRhdIue2cLmt54bUXVmpqCIJsXmnGmvN
gpf3/RwfLzpkkm1meAMafq68f9G030kz21Asi4jMmg/Kt6LeM0uJh0eh+URtmRCk
y1einnL8/0HejgKyqmAZ8IpVlV+zTPVK38BZzYaGd5EZnD6wPveCcd1R/Ld3+kqI
XOWm9MptRs88lYu1ce6nWvCWlGglSfySiNqwN6C5Kt9brLkmkH6er+qmZ5uS3TFa
y28sOnD40KTQbYJRsBlXjkpkYjEPXooGam9dRTHW8Mgfcrhs3zk5nMnTSEJO20Ld
Rt+5PORsTRxSlIwCqK8PObqA6rsSUxivntBrOV/o40zWXqIwoGADrTgRFI69lcKb
B+AZef4w0kpNxHnRC6524xHIOejsFDKziLBTgheG8KuAqig/HI2F61BFzyCnPimb
0Lz8ntZJ3hG8FDnsEbx6Ay2b966gG5pjp3F8z+ajIJPwfSXlwzL4PUmFiC27106Q
+j9vgc3l+JRaD+d1ZCCIfElQyPMn7Q02N0PTeyPeMHqwaH1X5ni7pg8vy88zALPO
q295tvsBHvA1rGmIQ5Wgh6S93Zt/qCwfQXW/EizmpMXNKphzOWATUpdEhLhoKRfL
zd6LdtWU8eYoZaKF+i2+FKYUNWdVDyvvwrB/WOPMXfSL5SM2akCz06RptEWBe2Bi
kIleWaTF7TnMbVtY5jWPLZ1nH6fDJAyIITm6zh6KbJHsKrsmFVN9d0Xc2l816m0z
uW7HR6z35V26GvoXxoEF3ZZxZzYZCqzuwRiSCYK/Aw0EqVIp1VlrdIw75VuP9yf2
J6X634itWDX5pTWmAy7fYKWEwtrnZi/O02k16bBLHglH3MF5sqc5yX4f7xpnvGjd
ydBkmnHoVmNPJMzX6TalUyHHemFFBnVqIJxeyLhiEboO9Nrb7qy8WgNBF00n2RWN
/AFSSzh9021qSwY/j/hnCZKMtqEnkQcc2DTBFmCb+hFBcSP+/AKq33dCULAIglh6
E/w0sLsbITI/P1/KWxS10yIevUYyuWllLYTxNhfLLFkdUjjFZAR+liHb018IOk/+
Q7eRX2i8gVTz0oAuBVlYaI6etIbKc0m78ojfK4prpIVGJ1pBLAEYIQknljEjPQRd
WsjNu7dL2COIA5xgVsWRfwLdQyLDpQVQt4E0JDIuvi9mc6oPd+t/JY/fOa/WJ7Z9
UqmSjcD0iDWM4yCGo26At+pjyEa3EjA7GojpsBRWjyDk65EJwpR3yplK10jpxcSz
oY+XSC7Rl0GumpSWtxm0yJ6R2MnqLS+zP0tLiz7KlolTUmb//+sytvghzpfQtLhJ
7BH1pMc11WmYg7I9Vu0HSRuaDEM9WZ44dLW4gweUF/O+RMlofqRsJ9UeJmQQwrvx
76TnA+2Q1dpruvptmROSCs6HsnBWO0znobkb34qlmD88AYVmMwxGCQ63A0uswA0K
x2JLR/nuT4S9Iy8/gMBdeKzPNvJrnXpkbqWFMx4G73Wx5eqCJM6nKs2kkU2rYUcL
dY8T6g+54JjLdvG152S3Rxes8j/ijubgM+7o2NAsWHeLI/Xc/DAqbmCsa9t7nMe1
lXVicuMNU2UjzoC5ayoaFW8fWgaAHEaM48Y7nE57uWaaUgDocYn9P7FawUMXtLwE
U+7OqsEphhyCx6HdAle2oN2aYC+3fOnfv/GiZq9p6iTfiqkUmr9DmZ6jh5x25SZQ
C+eGntj6JZDlKySSUY/ubluDTkPqwy6wkj+NSYfmtgomR/YZXA4HZzOto8bJZeFL
GBzJ3kqGzZSsmhTNHm9XYedkOeEHPF6mrJYmaHNEvvFjNdwq8frS4q/V+gdK2crZ
Bt3u3FJ12tMeL3L0qeqFSo5CpOowvTRAaJ6xtCW6GNR4aIaUHcZ7nZZdinsgXpC2
uyKzAkbXLm3IDQyAm+v+RsERFuyCs9Qa7dzNnNHNTlnXLVkfsRWrNeljl1UEWjfs
wn3/2mT0ujnAYosCirOqG8QSAbb2V5rjHh5t1yGqXwExwYifKoKpfhiEEfC74gSk
cZeBDiIBqi5D8/3VR1QfenBxFjYplmGlV/+U/RkDyluY3PcSIjDJg0Q2MbIp9a9s
or32tuKa+6OAtPi9uLFWeQpNsVdK8Ym0nuvukC8j1FJAbnK+5O4ZCck4tTUSHIUb
ssRr75yCO6ADCTbz5GMoD125DmQEoRVZeGNQUWAEONnFzxGiG62pGCkDwILhfkvl
wedkCb72BjujMo+S0y+Ho5ST9NjYeIXljOlqcs/hfTo28ko+u2r4m0yAaWCmjt2b
uXiVLxM8/iFNHPVQySc/wyv8g+gu6ouhQ3WwvlDlppbcCYihJbeNTnZW6OjyaTZw
cJdb+kTugsd3oQVF8GlI4msv7D7L9sKroOR62Z9NOwEY29PCGkHeWwp8G7WsUPm2
H54ZkQJkzGGJ9iNWXr0an/NAAHy4MucWp8lN41vEXFZ2VBw7gETyJD04U8B2F84Z
pEck2qA11NMiBK+EFM3/JlXg/AR6amhCJFfAz7TNswNMHuqAlY58Sj7YFfcoSI27
RHBFe5OcC4M4T2U3okevCCqNsLErrnGAjFgRJ2PGdVwdtFxzcwhCcADSz4R977xB
1HfIrTCt8cTpkCR9H3qV02kG3FGbMME/2q4NGscs9VX1MUKYWSghpYZSr+o9R6f4
kFajvBrq2nY3kEncyyVAcQyjuvhTedTbLZtc4MSI32u6iXsp6L/AatSjIGNHgNAc
tcGIeiqotfMncmXHRznZu6xZCz+RSoYaKNYbzwxlrlTOHV7mP9fENs/uqpX6y1f8
d7/5IJ29KaLGu9iI77lNaqAFK7LrdZ2K3IhiabaO0BxEs//dRE1D27e8JjecNxQH
V04hMVBKz8rkuW4DeNTVwspNyZmSIeerfWecdNrm9TDeDqky0383Rz716i8IjKXD
Yvi8L15h5XwyT016NjrjkoWigYpsjwl4mQBRY2IV+3KHQ3S/zz7hMQdfLWKP6tuS
w3aV+3dcSqsWLK7Gq+1oJpj0O6xGnLHo2pnpgFhUl8EQ1eDvVweNEgi9YkLFY5Vz
ci57YgSNSGG3XhSmeTsCRcva/4S9NDUE6XXQhPL6f7AOjYG0NZCPXgnxp8P0tqT4
DDYRsapQNLI2w8B09kaZSBVNEQei3BTEN6rkUq+l091scgUapZor+ZMbhIghOEql
r8x6wyAkoP1E9UPn+bibCSyrQOSppfWKuDHC7p8658igmDAlGG4nskc6hUcVCtZ9
Jnlg1UBqnBLB2U3atIaH2UCHGqCxEydf1uTueivwDS0uPQcPQRQmSYzdP7y5oKgZ
pXaGQ3FtNlcawO5vETL4MzGLlEwweNp5mvfRq0IWoMglU8tr2MjQz9Jf3jF3SaPb
+nN8NXKY4JfCnlscz6ONoT51q8Z53uYL3XvnmJEVfq0hy4UM6oiEyAD09driVxCC
Jl2SMSom4GlfLeUa2Z8j7VwR/D3V2ORGbRn8Tqqv/geAWYDojJLSzDrZl8YkKZkn
X7Ns9GXZEeUVcYarO1lfsvuxnN0X9wo61fA1yrqf3CVlJ1fCnDDrREDDagVlxoM4
EESH9HYU9NQCM7TuTA5R2MOCxikaFlQCJNNJEtedolVod/TijsGrA8G6LmhNphjB
9WwrqU8kCibfQJ/Mnr/uV6yh9ojTUW+odwRr7YwCPDWRO2cixmaYR0FagnrfVnST
tDkTeNzcE+/PYhRXMAwADjnV0seymzaICxuhloF0Qo68DcARMptqGGHrGPqpAz+1
1mzEsLi3pSvata4iBBBZW9TGQKLM+zGDWxdLIu3+R0F0fnM95qRE2c7gWWAUxF8n
mBwiT+y1cxUbf9GfcS97vz3eULiMMwkOwip01n/ztEpbu+OSiyHYbPs/63pNO0LG
UWZpyAlb3tH0UaP9d37JSNgMbMZKE8tBvUp3say6wWKvbrr8bD1vGr34IrmhKsdr
Rd9ZH/nFrV2CAWpPLsqoqPlVNdYVrZN/iSjbrF6XGlUqLTkcVbkFygCghyzkq5EW
GKR6PgLJWOdXfVN3gM6WuJ0ey7P/kmFhDSXCRX3uiHUpdA7KYU6YxABLq62q39MP
t0XyYROudvpRUZqO336LXv9laez+D+7kYqU6M7hIo12eiyWxp9HmCBeDV78UvH7l
Hm4Igo9Y9gfIOAwfGEZjOoPcS4CHqoDdN6F7ZwPT9TBteBFVibQHtiWCI9YZBGf5
kyURAdzuj08Tyc2BGVfxR2Z5Mgtpw2mz2eyfdhIImKbLLhzlGdrZbsLsPG9/1fTv
G4gWZMTUmc4ASd9Sy0ZQoHBVcQNx1PXLVE9dCYZ2tgWsMsPJJVcmtXFzjnXpuP3l
hvbDTDAoWz5bZW6P5p4A2Fqj45EOo0bwNdrndcWiVxuED9b9b2bx6LiKRa5xmwdz
Yz6rLzZ9AYKWYm2VFWcSkESj7j0Tn/InK4Q3/gHlfJdAQel+8Ur20JUOxDc2WdOX
T4vu6/KeptfrFluGlhJfsqtei+7GimaWoN9eA3dtQzvNM644IysQKXc1OPckJ5ys
fAgoi7CK1weSNO4YEW4JuHfzJR37oiTgpzs9FI7r2c3/3k8i7zujiHPC7+/veBLq
kpdDIE5U57YAOLWbhdJ2iVPbM+nkouqYVJEESm+/XTOcpiZBhIDBlsqPVphVRxPi
H/5QctIxMolU5ipVZzKqNVq37C4gxyVhpilJ8ePraB3GHdtBY+abLLU5MgzioKMt
D5BMoBWjeTA0G8/731aH+Mg2GWqo8n41cUC4rhDp7Waf98eg5DBKi6Ge7pbEvX5Z
2aBWpO7IS0iL592hdRnY5fi9rVa5Z+z5liATQwTTUzSgfHRQIgaCeHEfNr8sx+sw
3YneM647Vv7sB+FBkNPyFvPEmjT2VFbgDQ3uJ86fb8J7HdEIfhwYKOS5AX1ZKrEk
CzEFgNKGvQ83lPknTBd4vcAc3vsdbi9tR8AjoalBWA5PNx6i/DbgMtH4V1b0ny4r
3i8CYplEkeYazyO6pGam45d64Tb76MpT9ZyuIHLjK6VERNWjNS1zVSBCRcleIFZB
pNIaZ0YnCFnSzUC8Qs4U0BW8lkyL84wO2L+9bUGRxeeyJrGyvvHyNCJAO7cEiY57
Gxu+eBqICgfgTBZWjhGyic6YEEefgSN58XZc1/0NfjaM4+1Vf61yfRQe0L2nUYr2
shrzhcJfRXsQ0bFWUjZ7sPdv11Vw1uUQ5Iab4GoYfejB2owUrBYux6Yyia6NEuUu
etzieSNOG/J+Lhy0ypcUhgWvjfY6zxFONRth5I5YCwAfegjk0uYpueHoHM2ypYFS
eU7ap5u5QYhQ7p2zilXJ1HAcqO6qnRKw5sBeW75UhPTjelMUtz2vI4A1VIugTu8s
i+/X7Ede6+u7pbVdM28lbkAjwa27qmyLMDpv2aePoo10wYSKAYI7YwCQspIu7bq3
KAgxMpYkWj4VVju2D5wBA1tiFSogUfeUGIkpLOaNa/6k89cKUErwuT9QbxKm8YpQ
E6O+zwxLDaCg5JR6idK5HJizd/iSGN1m47pIHyDYC/u97NFtFO/Qf/d3TfBkVXZL
KksW1GU9k+PWCCBqRpff1eJxnc9GbvmLnDMmS9KDb+yJnL90q6GXmT9bpl+FML/1
c5wAv/jpmXe6saYOxqkdlC/BDh8PZ5tGm27/8G7I/2aVkMg6ITPKde3lY/ypqmpu
IyNroStkoE5NiZCBClgKPohriHWDis1gVxEfq9ur2IF8gS1fvBxtwXfkDmn1RzUy
lasTZl2tPYioZ86T0mouZ/d4/2AocLRVadXEn7gaxuq8Hb7qIpd9mX/kpUl7lET4
Vjk8PIwcawq9D68fw+zA1UKqhuVkb2dytl1flKv82k8/2gHeIS81Df5c7A/E3UWd
L2Q9MdRF4A/qGp7X4UYFkaM3VV2sXSAEBK8XQ9OnfA7PtLt6l7thvOkCbm60ARkJ
Xpwpaykcx6T5XykkFhLtooos4J9AJa/Wjmr8HnCX59jDedrX566caUby+9064I98
IJpFYqrVgfwivvC2lG66IwILKtX1DFqtmYH9SDPKg31X0WpGSmWnBgHXgoOAgBWm
LMTdM6xpA3UwaFIe771xupLieKbONXjUmWz76dDb7rKb6hACM6OiGj2ZGrN98xBw
i5n9nD1fmyg3ZLe6STr+0BMPT6YX2mYy0HSfHHb21pFD6ytUBsxXxpPt1rgUYOLf
zU5fzZ/m4kkbJM16mjcQc4PpZotDeeNfPy5BKl0lCLvjcWvoOPTPa1FsWPyWNeXC
wWme/2oPAtG9y+6csLe9e/JsJ9GSct/Kpk23eoqcm7qQdYBAekuUt3+HUWs4H1Xd
vJkwdasCF8gT342hK13jXDP1cw8T4K2X5jr5cswA9yePd1x+HUolG2+5JRV79REK
s3l7pIa3QtW+x/qB5BuiYo5heLSgaNvE4bJLTpjQ+OM0FGFT1ML8IP64w4mHODk3
iaqZ5fXFj1x7FMD4jbKw4JbxN2xEy5izSvcoE4DyfaW1oAuRvLLQxCrajOhPAt0S
sURax0miZzg5x6hFB+/Pu3ENDawMo7yjOebQact0N3aYF9G+fjFfzy2WCquZ9AFK
oUo8D8gwviGqOrM1C1ffKL72UdVCNE2DZ2p6bBYn00F5hb6SdD2XVUjtmc1haw7U
SFeOJKTSB0Sq+DMV3+BoU/0UDkI9+XHEzzRgF02Qa7W7V/WQ/YYSW8ZYVmyv8uNJ
oU39LYD4TtcPudRj94S9kv62nwIfYhZCX8K6g36Fz62yjodNAnnuzKC9dDrYHLNi
zlij/cT3KFdIRBClnWj1Yo4fSiuGLUf8yxNMbPqtvONbHCyH4VcoFLogY4bWyTvH
15eILVoD2Vis+0RQPJ1upBjAnISeneoPJ3RL2d7V5ghKXIILO494kWKbsiG/azD7
6bpx4CJnJiYkppBQpgDopR5YHCppdkK/cU5+u2xJF5hIKzPrJJRaVjCvzkbSSLW4
zXoYb/drYAkVDuf8KGFuZSELZcGqamkytVbhs8pzFzO6v8nwjCyPij8aQMLvOQD5
nGqBW09oTOVo8Etl/xfpUi4PYwe7VXrTj70fngiKLs1Zr5YZSFXtnGIp9pK0kfjx
ttSfdb5DqalqBkwDpx/EDeL45BSb1oV6hXE4nYRjFjLDa+6ZVmA+DoMj6KPqt4zz
y5/z7SyjUwcbUixQwcy9G1I/91XkwepZbjpfbuUFYBfSOahJ2vItrvtL/7FcRY6/
mt6ef3vuWivSO/VJc7kUwnXy1tRVBoex143TT6Zfw5bjY32N+hmwmHYzFDsSE3e/
5lHH6LIt2xu98ehdrrX23W+hByrGaa9lZsAH/LVK/9ZPSepCVviHwIUzzf+wvM4Y
bwSzHlw649hyHwuiyVUliEU0tQ0kl46OmF4gNVb7DGuu9Jt0MMW4hK9tMOJSgTWE
WltXMfd+z9c7UZgE4MdTaE3x6W7WnaECfNy77rJZv0LmbXmwU/URbrXI1Z1va6/W
kQVrYt1xjCJlwzXmMzrVLMGaxPZTuIP0b3DPmcRgySmz14bAlAYBpymeYa66pf+p
LoxNbEr+oNq/U+dlKUsuNVE2wH1+o59z5SxWpmT3ez4gwH6SEgzZKPR+WiptDpWy
6Pka5amFVVNAB+jC7TEK26HSgnygXIPOh4XUmOqAu5XDKmbahq+wJk7rPjC0YXfz
sPjB+wR0b5r9HSmg1w3adPtpLFc1T3tG6nFlWPLxsgDXwqucFU33rxk574oZIhzr
F4ya2AffYwMB0XA7V5jUgUmjmf1wXm7XxZn8i+DxwnahVf1woRyS3v2SR0EIsY+7
+V/NY4NO63Cp1fKn+hUFSOuG4I1k+NQw2g/gCmOFmPFgANh2lQH+cOVZNJrfYend
Zbu0IbwvfXVOs7aYJCFmgLL735vhghFkAOcX5PSO856Twkjfuh+F/al8IgdzFDQm
liulSxhDHgxx9mnEFwds47Bw/PHsrptniKT7wS8bJzTFnOvM4Q4z4kUff0naHtj8
w4Rdiv7awrG8A2fDWIanq/lrjH+etu0ZG9yH+GRu9wKvkCgdQY5+8QMStNEIfgdm
nUkRh+0/R2aiHDjCndG8WoY+fCFH/PsONQUAMkn2zVVfzgz+ZEHiyLulTQpb3v20
0mlvXXlLAAvoDPBG+I9dxvY0lU7WZ6X9OEqGtvbBE3mAZxivj/U7Ln7523JcV0+X
c037grVLZjf7J+8cS15sD3bE2bEoUqImgUhQGFipuetIZ2ChSo7XM9P+7MmmT1I4
zirUzqxIOiOhl/jj5JPQjHytZecRgvdzCXBj3F1asGXCkG24nwyx1LJJoi/SOJIw
+B4LCPHSv8TVyC7LmA0c/tMLqCdgCEVqEz2nEEP6a/jAKdGi2B6SDo7qrX11irGe
bTxCxpYEvhQox3gCFzs7s1IoNVQNuzMI53/834jICfPpkikAtuynz6pulav/RNQP
tiqAa2lHzKBTgTb0TaawXIeIxr5HgOYhwLdZo1fTzIljcmAwIBdtM6Jthu4kb/9i
+1S5N2WbHfaDAYvqmokN1H9dPF6L2oIBPt5+re6n4IKr4RoN/V9qDCFdl7fF1ej8
zVXkPv3VhkH/PUgKKqQpoPSbmunJja9bMv6IIR3ehh3oFalKgBoJ7QQYplRsl6jY
3ANFTttMuHvewWqLdhl9iDz8x9OTBT71d3ZqEec5EB6qsnvHzBHRllQdMkrI+xeD
BL0dhZBckoKBb4lrx4CnCVg1kxjUED3vbCGOo7I05w6W0+b6ARZil4bm3QPrTlvr
YNUjLTKDPlb1UIPh8s2Emt1te9SJDm4+d0mvqyG2g6MpIQBMVgdBG7YIPiX75MZv
E7j+bfpVJLwhoHCe84Nr8bnHfFuIx9piyvAH2Zn29My+hdRYPmtrRAQ1DbGhpP7b
Cz/kf2BfwXEF+1NeX5jML48NaBukvLRduKd4OfDk9nK7FEnxT5X0cEpgoXveWDx4
clu2t9NNdABkLOH5Uy93CBXJYH4OId+2dAi6U8bIxK15cwX1xJWPh5tchZkgz7VN
gBnTK4ujBMpc04xEwqpLkskOej5/IXFPDCmCTKL85oHS4RiZC0TPpLFnXk//PgeP
mcRPFV7wOLR3e7ndaud6I52BksdwFH7fE+DJGTLyKzq6pUgraMgICOFvxuITU6CA
6bdfrElbKZwiOziXbx5kj1Wh3QThcq+hts9zmvCLzfRUg1kocAQTjICKDVqaf/jz
dbuESV9B1dGvIARHdNSAGVcJg5PUDBtfzaRE8Wb8eXlCRaceGtzqhSltoNSYXfgi
pKbX0ap+v0WL3hL7A/apIZSasTvfRYrpVlybN70VL1jf5r84+xt2PsNh/eGNZeuy
Bv/dIpJ0au/8Z7ToVrn8yVrelXR49jGQTklyFp4k+vK2UCC5+O5VZv+QPRJ+9evo
COEE5X7dSSS9jbsFg9f13aw0Q72kgIxgicEBiG2b5EdA25E4POoQhroyaLviovHU
iSscOXryYBj1yq3JYfhtOZn8r914CDgNixdZf5pm2KF3NRN328DEvMoe0N5nQCfo
VZaDrgj9y4b2LpqUlhz5x7kRpHvcEgs7UQneh+60yPRGyDWOgv/3fBXtNz4h3cta
uTMoLMok41VtTlllo73rcYtjXwg9bOp0HG9AM27FUgsiN4L4XkIMiV6knrapyQm7
0mVcRB9vYpygJVfoNrCgOdH6H7i8Q4jDXmmcOxmbj027r+82IocCy0RZ2LYwlQgK
XfqOjJCFE84y46udP3FAaPZ4NDIpSxB64n3sVxHIuG8FHmS4Fbx0/G8oucFebbMH
4sYRR3gja6L0+vxT6U5xmk75MsbgCCDUuBfwsyD20wBLcP+nvCxq72XHqtrW/5W+
+4iuA6vJiaXsIp6vz+caB0HB+gpsIlEpwSYB/POkeJsOh2s3uUbAleX1RMnjCfwT
R3Y0Ml3DpkDSxgzsgUMCX8ZH0Un6ehDScPyQE0y/ko4iI5Temk+ebrw5PqoaGECT
pjo2PUlQt+jjIl3kzL3FNfKq8/j7pdrqqVVErSrEDQSwlaACFU+lYWtyvdUrNASB
A7u1e7kngffXqJiBr1vlDS6HxTVChNO1v1pyZxPbYVgd7YWaf1dNts/wLPVsPWwH
5DDqtpK1b4e5LMXxPWuHgt/92HekcuL2t1GJ9K9+CxlXSJ/MrSjZCwHE1DMcnBfb
4oIcuEfeUP9nepjvEqBdR0jVgxUj/nCLziFidMbzVRRZZIcrWYbezuX4tdyw3KHD
TibHYpGVmb+AK1kszy+H2GYrqSrH9Tgxm/ajh5tJhaG0Ndi8DqNOJYbDjvJmRQYZ
FeoUQQjvrkKd4xVAp1AI5FYGZC9r+4K2Qc0M42QsI0TJ2LS6WKiwmuN1e76sBEtX
yI5prOEtYxyTgBtNvLA91ahOio4uAktlcEU3mG7N3hCkP/r74/MgY2KcowcXcMel
GoTaW5AkemIE0bXRqycvXuPf1x08Gxrw2wtsfnS68cJ6g6gH4UeRnSLb5CJ1zT+E
+zlJ0wh6kI2eu9/GcqARfOukdquytZ5bABi/g34R1ub0E87KmV1ld5qgqozZSgwY
wU18Gwi0PT1taWo2Sk2FlK9wA1pFe3SBhJNhq2PnfNnv1nihSsgo8Jutjbh073H3
1jIL88yKethSlQu90dcn3PfW+MhbpUKu7lq/WZG+Mxj6EaSqq7SenMQDgF8P+Ifo
zYbk76GZ7Gwjm9Z9ArLgeJxpEYSEcu6IiLKe1bYfsdEl3c6z/SjYc1f+XbdHPXa8
lMyJA8Xz9aSkvZV3aZzIQEBavUuP+9A2lcxeHMO7/N3x5giVxpNpMWNEQpR7VY86
yyECo330i5AbqSaLnLo1OWb73q5epsGT4XKnbA0E40Krxusul5yRKok7xJWUUJPd
Pw5r6afB/R7idhZqqCn5zvxtwt1Ghosmb1YfNh9phEvZehtO9hwadwNVLiF7DhDW
vMCj7294kqul5AZ84lCVmij5Y/A9KHIGxcRixenoXVNNmRN+mo2YG1AWR09mNnxB
Av7qXX9AGGRyJDMBzwcVt5ZxdHWIwnQQVX7+zZBipLNWiQ0P6x4/VR0v5gdIi+x9
X27dx8KrmhF6kOwJSklJzDdRHBtj/O1ZeLoP5JBD17fzE+StCTw1xY+Qsti/2jgH
zq2+Dir4TdFnKzrs57Yx+YNdgTVtYNv7WeW1VJ3oaYue0tK0eM0hkzVPOMI2XnS1
yghA0kXIKOjSAB/YfLL/0n5wNJTRoIcwzoKHVznkRg9jUyOHD1G32Xzhu6GDmZZe
ZSbvzwzBS3w5HZDAAPM/9qhIOAd5BwBPFiKGrG1NqnIvD39/Z0EXffMcSPJn9E3+
+ZWtw3n62Wr+Aukdaj3oXK/55jypsZl+ue9yS/hW9NwVFBXhTUygRhVhaN7TOey6
XqXHyrWZotluopklzzYRaTPUOI/5e7y3jmpkhfWdu0fd6pIv8/jy9DXJ5V5v8emA
XEzQfXbRxK5S9EJ9JYRpWv4Pv4AHV1LoJQfs7e7dH8bJ5v7sZd7k+UVf+SDNwGbU
sWWyYFX9AJc9Vfa0P2m0KwijZn5+y0puas3rbIsUyFOLIvzU39MT6Q1JQKm83AnG
mnDO3aEz4hr+3cv0CmDYpVn12EIKcPYEIud4OJABmrgXCTiXDQcQBuP9OauAplnw
PIWLCm8HcOmyYFHvS6hJdkdjW4DMQlDCksgVKKrsx8Z8D0v3umktRjL3ZiOL4i5T
EXpQQIBPhPxFuYYl+mpdxqvUjAHUpo2C/b7jChonCqN9aKLzYkOuSh8HiliyWMc3
eFeZji33ZflxAGBMUIK1thY/G9nzGkwqS0mW6iYf7jbN5n2NXYWa2iPJ6uMnEJ2F
gn63Z/Vou4pjvZEPnNVxRJtCdIht6qcwW7zK2sMRDE9Hv82ae/MBEVWXF5OAaDRv
mWk/re6SHPsV6vc3dUAekG86MSgfVFVda15mYB0zueNJdTWc6a3OWpn9KBXrUKXm
1LFlKv+k3aCovalo2OjuCgAD4L1Vxy7ztcWHbxF0x5vR3I5tUWGyaxA7DiuLbY6/
fP5RC2q0kxfuVgFmMMYzrDuYaZlDJZNO0fe18sa0+O7U/Xu1J4XRyi7vnYn8Ej3/
Lxz9CcQtKxO25h653sekxzkOql5YeO4o8L97f3oey8zY1oJUqxhUhj9Mw9dYDmCS
i+/45poTcp5kuQ49sIOZeLBHwI/BQUmsUolfw9Qbc5sfylqAtZQi/owDbBsOoKje
yNBgDMIBschpcWkx5qKtgVtFRvtFMGOsj5GgqAOqJpo2u74ZSyGEQ0Js/qhgW8Pb
frTrwt6ZUjlAceeGnnsGeq4t6nrq/swZQWd14WFxkgDfvTUOTfcGcIaMSPKmuqCj
HIVbkaF69ZHjqpJVT2s64ihi1+gB0vtZLvtPz5uBDs4LMHy0JMG3NU7tv+XE27Zh
p/l5hu5aReFKQTabminWhwvBDzQj0DA8N6yvPNhJA0e3Qel0XuVaiFZPDvgWMYdS
wyBudlqAYrp/DcQemPP9rhfpyTSeZsUDsGW7q7UR3Wpw6Tv6dQaV+svvx8ZLzXjF
FB/yL0o8V+KRQ9yKMgfSw7r2iDsKgDbvagxw8ycBnTUM6HxIv5gGmNjx9DcD8Muu
WP3DCovkli9u1nXKl3tDsSkbIN3Q9ktEF1OluR6I6BexPWPr0P2SGSloTfVvFMfD
UwNVRV/xHnGQQxxQb1EZ2924M5kEQg51xil5StgCR6K16zGL7iDsXODXWfEHjKoL
86hRoiZojy6k0H0DU9tT4kXzcG7tG9RYfkzCse8a/Y3tPzrfo4HryekWfcda3B4E
n9Eg5YogqNI6vG5uDd0VBtLWyjF1dxATb6QAPjg/dEX+BOrAK8PlY195qI1EiMNt
JDZ5NrM+VSwXRVWff1/Ocrvgfahg3yQ/fHogp8vF4ZzUbHVhXuc0lIrbKCl6CVQn
HFBuIUKRdbsAFMO8oqu6uhdEUaJWuDgngHZElG0SQGht5Uc6QRmuhedZXPGx5MVT
9acCxNC7rhp+c50NPz/izOAoyQfXjqd/SZiDZqZiUzrgM4HCnxJTAWIHk0tiFCjS
j7JYzyfAbDdqL1/fwbKnRjQStu9iQKZdOe39GiJLz+U9DBGwB+2DMQPxd6ZtR4cR
mVgikjQ1jRrxInZ1kULvj0kHYeGNAe+vs1L9m5nnEF7Gx9nLWtK9LaiZvJilo+R+
sAF+fDZ6KamDcPPm2vDu4DQlyPqXZYnFLd/iYr0oSfvAUgnLG3/TGUtCgxuJF5DE
4xPNtGzsIwGhQDFBwprgNC0ftVTOGGNa7LsLmcaGch4lJD59utHjv58CcgoLPoW+
sPFZSn2AORUSJ54bIuzVHOMnYGrDKvrK6Odm627GXwN0tl2131+RC2LSJoD4OoI1
NM0wpaQ8AHEg8ZJKpv6mgnY5ABgr3uTupkjtkOd1U5OyzgKmumdFeVjwTv14i550
Ia03svMJ63wFksiLdjSRUXFkXyGW/R6kghtJ4vH4f7hrX7mb2tZlPhkF3VK6MD2r
1hce53HD2lTs9UxFwJZUgOR4bJehFDsId7ySMKekRiAm6B7vFLnyGhNmgp1bspg+
ukaIDo+24lg9ct+3ohV6sIl48OviBlvgSGtbcuTc2pwnGo3i8S7GX1ohDWHiByuY
MK/4mGqpRoH1q3tj3qRy+wlYsQkE5uT2SZwGMgutqI1vxifOedXCwrKqR12Tz+Fn
9CWeHz5+lUmXCDhiHhSF/fKLCD8VzyaB7o5t1gDFNsK06y7OlVg63tre9YWAHPir
oaWR1k+SR0geUoiqIVw1mPzvcor4V+S4eDAWRRisa931Oy1BlCVPa8YdSCBVsCzO
6MfpN71i+QriJXqD7/BLvtK5YceJBMjsS2C5lJJjf5J8bDiOYZX1N+2cEJWiztGs
tesOZS/51zfQOI/V9OpzEmowzOmOq8IdRt+gqtj07+bBS1XpjwpnD9jOewAoc/5G
QyN7NHp7ooSi2PNA16eXEb80Uxq89X8y+8VO2NVnko3G2C2nuLraPe9TxFRkug22
ZOx4fS9jso2HQV4Plp4uS2XXzw4hWJ3jcXB1YVDUEZU3YlBb8Eb7QQ6stJW458K4
QAe+eqpvQ2pddIDzoCa7i6j8Ijz2PRofhxfMSzbCArdtK4JJT/UyHTdHcwW9S4Yn
rbatVWL/JpvLQ2CjiuIrpv/L7O3495aCmvlc7afcSq/7wPW1Eulk63G2YFHs5ET5
EPocmIj3OxeXjJf11ipjS0EIk6S6Y8cqBOkmBfI+a2GPOK7mT8JyLYOXFGmHilY0
iGJvpv3RvoR3fF0/BgKm6Ub3N2RN0CVh6w75ZNEz6BA/lrBm9mSwux4i04IHYg5v
1ipQaa5OrAxTzZllhx41gGUjPE+hMr5VymHJ8/nshkYGSPe4hvk8XvnnT9UP19kB
NOK7F/RAn3h8XdBnZ2dA78kyBbwV73RPa1zfptnRCLjApTv3Dz6e8/l06vfSSy6I
ceFo9k8csKaA6no5wX7JbD9dRVmLUad8aoh2Nhnx6QHX9X9VuMEC5AN8lWNMoJ+W
xZHo9lc1a/HL61JUnl19ftV+WmFXjYy4bgsLOT8w5gMDy50gr5Ucnmc/ygrjVRnu
1X01BHRWjj/5b4yiAEfvLxOUwLPtX+JVzJPxJ5nGq7Oq8eO2cARuRtZF14qV7FKu
1e7LVUnk9MhKO45MIo4ELwlVzUsV2SE/kFFjRTu6UAc3zPfpxLJZY5WD8MJmE9fQ
X8K7Izv1g67ifPWM/PlBepyPw6KcIQi04qZSQegCnZXPv58tm3scaslZVCBhK0VP
gjxpJAmDplKF6Os1cyDTDgeCkcnEBJxGIog5R3kR+Mat+e+lYkOe8HojLPV3qmu6
sSwNWsbdpaoALkrFS0dv+6Lf4haRSXs0xvLTTQEU4dEdpEjJTvlEj1Xyx/QNBAgu
RLKOVZcVYp8Qmua0NVrGnnRDY+vuRB+m0DC8Hw/Yv3tOQ61f49m1IcwkbaVbCrVE
ifiG4l12bkrhfO9zn6WcPs5t+oqmErcVlRkmPXa2T78ik89dmEGUf45twoJoVJQy
48jwMlCBOjifk1VBSlnWit7a+HUITDFJbcNAaP+5V3ZZEoAnh/F9UDPIOsD41y6a
OeG6V6p7cBjYTKi37kKDal+NajkXoTAvoEczXA650Q3O9WJ0MQW/L1/8PuBrgrvn
pI/9/7mu5vnivN78+/Z68bipamSIfXHsCcZ7gleJi9ac+uPBuzEq13KvRrqigKKX
KR/WTOyVWCz4JZNUmW17o8BZK9YIMss71QtshRkjDeMm3F6aZZLMw3guV1SFfpwU
i/xapMIERAvsgTIgM2/UB1QCvkVF+LlZAoArP2FGyX93PTdAiCo58C//GlqtyAm2
DW8hAE4lNlFisTPxOwOHaZYuVTdLS12+xuemCcMa27tK+a92Cc0ZZZAudTc3huE/
daQrPG5TQXgkQQ7NOEFX+6auS4vfwg6m2bhHowOuHD92ZEqryHCfkZp0Ub1ikccR
GzjMmqRFSjZ40fgYrUguIzvrneBVwZ1WhOczpMfFDLcLeovsROLnOBQoDHp38wYQ
o+WIWHA7OOK3NOb2LQJQEQ+xyR2Qjwp1DIE/Rlg++Wvbx9r/BRlvmIYW0R8Od1qF
4D2lmcTW+e0A1v+hMJEaB3e0azQo8thgqdln95Qly3JBZEDC1MQ+UGdYyePwLXm+
j/LhPjEvRdlk4iJKKMF+t429SZWihnmPj9dDZJVeIYIKrDd1ehe+h04K60rStpq3
gk5O6fHOx+/hGEva4RdRaTK8ahGv6+43a9v81Xo3rJ/denS6QfKFrcmgTNmTyzFa
LjlkdYC0xab5v+V31A5T/2JMcaBSJCj/It44UXx8xwT2anCnyZOkpv5U3dbhZb8Y
0n0Kag6dX+k+Lq08A+IsVD/JYtTyrdEMpEzkZlR1jCSS33bdZe+4zMSXkV9qiD4O
ZmYTCv9bJL91GHnthv5ZHS0eGjUZAa4uR1j9JrkZ1foZffcz6Mh0LZg55YZGTNpj
MvY9F/PpPVu8KL3D95/Lc5N6E1wOfv0EFPQhVocSGtVDzbPnXhmnyQBsLGiINIB9
/cu4DVYYY/dXnnazKd8KYZmhiQWXVoO2/g15Wi9+t7rUQYpwdGlT4bmdBTJGPy3+
sJMwKAzI8c9/ITo5Lbc5KHImlKbPwj22EIu/DC4jWR+G2n8c7r34jwujn4bHW4Iy
A/kKF0DuVDNnhJD42y16NkCyPkb9+7UY4cEF1pD1czEUT442ci8D7rxpyByxz1ug
ap+ZFJV9zl/bghkfiyKyXi+ZiahZ2jf9obLOugXbUqTiWLuj47+DRE2gSo34yXZX
N4cWrXn2RslzJHl+8v19nIrWxoQqSUBmJ/wm/gFx8hcrLD4cboKx9Oe6yoP44Syj
y2Av58rBkmj4CoUAmEMtRZbvkT6OE/jKgbj5SoFraGZipeXVYgGoT+ZhwURp4/F2
KSCxHG+R5/MlHsZh/WSZzsTXHQdY+l5VvZ6Qtdco7RGsYfbCdPZRpu7sLyyKIZYv
K2QODIYwFmySI55zzmaJoa2+Q+LOsvCrAXErB1IknE3IwuP9wrzdF0PISJ6M9hBq
mDrKdjU8oHEQ92kK7mEU6rJys3A+dyPZvxTEIMsxl1hNmm9yfFBv1s+TQWNTWiXz
BhzFOIMmwcQi4RHzn5uUPuY/XxS2rVhvg/dS59ayglAL5nCX047Uc9a1IiM5SSIh
ejxz4Si5lY5LGurpt+4u2dldtaCOQJzmnyHzyQdYqDvBbu+ZOy1Ub8cMCGQgqrf6
/m3FNvJdZPdojDom5DQDjgIAnj0eXJevwTuc7FsGUHgHXdfTxzmMkZDTECFmTdWk
Loaqx8F66OM48dEXKCBZkZK6QvxhPtMaTz1ZEJbAwF4cGvoza3Grfm2ki+8JHN3s
/hJmpj67s5xW6wFJgNeD4qtxYRmNl0HXSon+bmF7OcFPYaOinuQOj17svACzH3Bq
vDLmQ+cpnnb855zKrRHt7qKaxqhu5kau+uTYM2eJ7+t4T2THSIvKzsqyKClQbJdD
J4oqUlAI9YUp7axSPSi2Cl83Tl8YctHiA25Qb4mmavaMUASjExbDRVybdjoWiM0I
KKQUIiC1KuJnPgpZI5cEvWK8b1IH2mOnaqw5l6AJULIgVWivccVsGHYcfRiSMsLa
UFcZn4+vKnkyXqr4JYQqXLWIVtXGpg2bpuX+w6rsSo0JBntxQSDIviNg80QmDVoc
drC62oPfK8u1Rj0DBM9O/i6gnqkur8ss2sN6jVbC4mJyWdK9mb7o21Uu7OBg9AbF
08ROJ7N2HWHFY44eXnv374HeaVLX1pzQSv/MeENoBeXMHbDb8fheZEnbzsz7jVLf
JdPTfpg7kHfLSAfFeQ1vqJ6sD/ZW6G+REdvpk/blJjax1EMRmR0Kovc6UiOayW4T
xEiapRbjId/yl3PGZRrNDPltvoQqt25B83rsfD1pjEHX5az7XJhmefwFc1HVh8q2
lr2j2k3qr5QdYlH3teu4AOFajC9p5p0E0D7d078eqIbVOOpAjivr4n0d4xmgrvot
zWzO/1Byi0S0U0XWxjFXJdoR3sPMfJfFRntBzYvqZFu4PvoxBZlTv3Ja6nmcPSRv
/EeWJFVgmfBFYd1y2gwzVy0HSnAmZIkyLN8h5gmE8bng54dzQpLzHnlXGD8uS0NB
X9ZWhjayQlJQOdGxNDJyEmAb+6zfyXI8Q6hhfAwkKAqL/Ne0hzJrqz4JzHk84ACV
OsRcMqh9e+ERxWPPKscvMY6EMk7UtbsxRi2g8V3KOhK3Vgki2Vb6qS0EtfRIsAV5
wwDwQfraNTMDP2W0sL/eRizvtWEMAhcOFPI0XB8pLLDg73KijuUq+j7R/jbZ2VWH
SgW6fLC9SYIRv87q2dPQt3dLKpKPBEtErSu54MTBC+uXhWQX+6BjkJ269uL6I/ly
luQdqeT1x+lNl2+efPvmepj3ctM66h6XH7FKG5KvDTaufcAtlSLAT+tGATGtJz3c
v46OLPJO2zWZjXILF6Kbty+cpJpzQLNJON5lbnOGhigeFz1cBy7X4h0eggNC7mJK
fpiFU+K8/U/pRabPUzV1LRKmPYBvy+T9Q/1e6Aqrzn/ToU1HpvjfUWgCuJx1u1RZ
XyOT7N/2y6lyIG/oVn9bBmnNq3cdQZoW9LQGXoCrGGF/Ok8iDorgYE5r2p4JuVWs
mvRf6smsJDhY1vnPQupNv0ZbI7eH2FGmsMZbTrXI9AY5GFML0icZY9Qwdnqv9b/Y
WYBqjHFogT+p01ZrxybfqEasCyBuKih0HJA7UMEVOpFkmkHi90hA3WK0FPU2ODLB
yyyP+AOHdkb/3L6wPA2ELLlQoomPajYJR6lRK3dFT9Jh9p/NqkIX/TzMLqWFb1sV
tyNSI+AEhiaOxP1ie3Wo1oIRpXxJSqlU1xiOwAPPlRuhqGyeA5G502yar7myJVwg
sUOaJgRLBF8fTJfc+3o0XtNOGWxUvkvXUKvaaXatF+uasFNc56UtpVbSnZn0SlfX
QbEAU/XpLf6HPKGTQc3se6Mi6kRZuYaVIZYILa95JSf10TixDZlp3vl/hW1OtUOj
XMcD2AAmaNOGHBz/6Hxivbd69qEeWpFRJ0JHasbLqU0IKo56y+fe+qq9fs4/QhW+
6XEzJu1jjjuwoBoK5f7Z9wvSKqbY08v+wMY2VfQthRqolFj18gVa3pOIERkI5aH9
SIc4Dp5gbPAi2z/0l+LVazwdNbb5N567VFoHAzGZzQbWPeFsTxy5dOPxx0BwMJP7
Nda4W1QuxJegSX2ur365cKcPsiutaXRCwUMeVmjQq8G2osybNKbq7Ldk0to9F4cF
YtAQsZgSofyb6qVCV5Ji6GyOaVPuJPOKOCzTeLXMm2PWAFQQJA+fTWVjCBNzZRSA
mSa9w5TmiHg1qZrTkZiAM6UH4tlz8aUwTQcOc3MfdHWvXF6foY6Rf6c/qiibdoil
aWAwXvWkqFHEb1m1rbyz6dvGrnFBtYtMEG2/TRr2YHlfhHotxp3+ytm56FjjibYr
NU4WWuIzDkHL2NcuRza8Nm1Gj46jtUGpUiUBzYMsWxizp6yg/395BW7tMcSonfuT
Kd/R85+DfIaqSMbWjJ5ao+vwxf48AwSAwGO4TpglCzaUCQmqOIu6b4/lg2cir+4u
VAD2mTpFW69oaXj/yrieVtYwexw2M2A5zjPkAfxv89KKabo/Z8IftuEFgRcEdirL
ykjLv/mHxQFRyf1S9cQB2WxjbOZKIe/JH/wjjDhYPVrLcY8/mgGAR3WcUbBinl5O
xybh3zaxipDUi+jzWMzbznpD9SMi3kfPIphIww8yqw8sK8SmfWsWJ7T4P3rnaobI
HJa0RZ99TK7qNnmYNVQM7iLYwGh26axdBjhk/6Nn8gMTYi7U5ipc79MmldPZcw8M
VeFVNLZA7ZYJPFy3OEKfBjpKpUdhnWQ+gKs1E0b980YujjpnkuHHw0JT9NhTqfDM
gLB7no31Iq7EkFW7nngSQnS2bdiohWd3+dXP7CtcrtV0ClI0SphPz0FAqfKJRO3a
kgvClYwM+LTHlR67ipf4SfYshhrrwy6mk8MVxs4rM//DnAFsayRKqwlggtJGL8r2
oyKNdL12gM+nUNsZCb5BgnBGynRyU03AzU8sjQc8VxTxTO5Ryn308biVkFVnmTyK
ncDZmKXueh9ekK5X0eaFA8arFVYQB3beSQh9fXrTf8EaSblGDcB6k9JUR8Mfwa2A
VmkprRTr4fDQPs/RyxlDm6mqBmAS2u5BIvZZrfU7SfOWIaZk6ChK6FDejr+I2kvt
JbGzVT38eh7kBgTD4iA2wZUnbQ7yjr5LtLThDi1bwlQ4ssIaTgWTWD6SSBI8LNXI
Y1UcWSZMYYRH786juanZcHrUEOJ2Pcx9LGAk8r/8t4bnc05l+pVnRWTiaMlyt4yV
OdiHvhoQ98q+WEwMb4XMnxsM9/3yIM1xRrZzyDOj4vt5j0AxAI6aETlrAaQaAaBg
m2ERnQ+HP2U01/1N7siqSv7qzCvsSpE6rZgut74vpTRhdPjCEtZ+wGpo6Mh6hxi4
U9WO6W6VGwk8k3UCZC96nxz3DVLh1Hz0bUckjl3KvlSkVnc/CgdnK1XJ8KwtihuY
ZedwgooqBCrbA/E6zP55ssxtTexPQ+ApvLThqf/4jq+z5iTi1/dN9WuJFZtL+SgJ
JnP/fqB+yPZiTQUtbljcDSTgSDh5xZTmkhgu6HevlLIftCbvdo0rFNR7mlotVj+X
zu10xH7gyHmbJDgC3uAIwZgOTP8qHUqdAROf83yCu/k45+BHXCue0ub3qqDZHg/f
wSgfCzuBw/ouXhFV8ZwzdR9DXJEbrJhqtnd028nZk4PRJm/QlwE1CmA5G7Snlo9p
t0p4uLVKKL1ByoejTXuTLeA7EclR2ch+GlDyMukazx53OU8QSOhLOTY3Mc5mX/+e
JAd/0n9zn00DGpn5wDJGPFcFpenSrHM6oq8Pblc8ALhKc7K2KVIk0cooDK8czbZS
yncPSv1FMQr8pKHPf1+nsPZTf8v9VTlLnqN4Dm/OafyZMP5RD6kdXTvu8lB6cO9s
TuZTL895+NPsT8p4tV5zdDydSgU/8g9gEoDpEHzCtnP5MjTy4647jasrvj2Askjx
YwV3pux31gV85wZUeZgzc30EptJLhwiinQgZZEcYT9ZdSUHFJDMvQp2AjcGSBq9Q
E6R455h55bPm3t1PlDveoyrP0SeHtS5L6MAOYQPI6lD16m2abf3Iw7Dn4wMlOUqi
HGTOGHW3cHhgQBr7IguxgvcAdWmBbJYgnQL8H8WV75VoQ5UOMA0sfQSaZpz56qmR
i0yb72+cUqPSrW5H05rYpD5AOKQTU2blqNG2X0tS6+lB2Re+LeO9z3XhtoEuQVVZ
GabjMlaI0amCKzSvhl9XgUAJqsqmJUdKGIqiylD7dDNSEFea9nkDFTkhAUKPMzS7
hiSFoJOYjkeCdyFZKeQHlGwD+++Hgdau1dasMS3MTjV+5/3rmDP0d6PGWubuLIMS
wlIRSuzREM0zS4+XpwJRtHMUvw9eddGdXlii4UuTXupWJy0nF7L3V5BHyy8qqLhF
BpqF6RC6bJfX8nWYyWjp0ueo65TgxlDdSoAgVRigqa6Gsm/JeDcJDbjRJ6KwpW0g
PvSFCuXeJfx2v4n6M9XXiYjAibf8eFiILIXBRFnbhF3rWfrkpa+hdvBG54HspkDZ
HO8hWh6h8+7FP2ngsw++dfpgN+Utn/Daq91iJldd6ooPTpiADX+JIB4RsFmbx6+l
9845UTLZECT0uLo2C55xYKe/QQgfaIAOnX4UPjOlohgGgQr0TKUxyQCJsQ+zvl2u
f0bgez9alP28o0JB+RwR8EEslkRbH/Mz0/DPLDV7VBwa58QUHSa0FM81loQw/4wP
3IpsyGRKkw2zl6cy02j6zYBEOSaPBJWPqp9gMjHTz/qBztwMw6NBcY06q39cPXD4
xu6wTLmrz/W6yH/KeXjBwWFfVJbeoZNudxmUnY1i6N1JQGoDUTaynX5h8RUYqYls
jPloE4cGuqdAOmahypC/WrELD2/CliaBuJjLP6EO0I+TQlqW2a4NuKfm1kZ3ZT+v
PsArsiQbP7XL/21trq1RnCzqlFOnEDoyQQtoJSvci4t4LsXfyyb1U3FGcwJb7CZs
C1R5vPWwABjkCPFOk050bJvDX5GP09p+glxFOEcdwe4mtoxmlqw02DrmqscMg20s
gtNrVkkVw+PKnhX6K+MTUXmoQE0UNzFi4qn5Q1KuP+wCdhg0CexPy5Eyp9og3+Uy
jf5/ayTBYAwq3RLgXp5EVigwqeevd0PJAhRJfX7cRoVkxRwh9puQpLpfkTgu+CFD
6OAs+4vHqkNcKUsUZlgPyoGk9eBHGkUGWo90ZlLsUmIxjQY/Zn90oSoJTAHHD2ti
4AhhyEGIEPhVsCNf7mXsMyzMnknFxMKhMECYCrayQp22c3UOjdEqZHXgvJcXzYUk
mTKpfUCNqMSe+m6AJYZZCB4rf9o3MnXz3Z+AJXD23ef+8ZHX/DfFOtWv5RwcV6GT
cpyCpwaZzGKNx9jv6H+iRWiHG341bMuJSi7OlYFQL9OTHpxCvPsoPukf8QIL2Alj
NUJ448Fsp4JAWAsnOXQqstcnihociYgmBihEJkmZR86QXWuC1CcY0OYT48ujN4TF
bUtUmKVe/KFJ62uNq28w/Nmx3hU6aD4tIuCkQAy1gY0kFfxrinL3S5wx4VFAEL16
n00Jjczi0x2cJqCSEzzm8VlGQHi3Etsmv3Hvn9WVCitu2kXch8sQfxvjYYjXN/4Z
EKfV6ECjw6UVp4Jc4XUfdQSE3iuGI00dS4byDuQYBSrkg9P34aiY3UvEX0krDm6X
8VzOp8siAFkhNEx0iHY3O6EjTrxtgsIyIucaoCfGhv08ubv57rg5fkVBBlgexVnX
yQ1A4ei2dEWUEVEsP1byaR83F6YglkXz1KDRlxGUoCZTA91X7U9BvK3pNRyZ6Uk8
QOzCOVLjhS0hEcKWB1skz9763P2ZqH/Ycv8AqrxVT5aatGExVbj1qsL5AcE+NLvI
OnmFEYd7uvNJDDWCmMTpWBhAvU5d268chWSfVc3HI8+Kkidqo9PinXDUcqZIy3ag
u6hNFMQ9aTTzhSvHoMvsxMB+B95xfN+o8c2bmCTujSnCaplcHWNYHt+s7IY/SkIP
znSWS/ERZK8dFX9qfR7lVsVMTcGJIxGv1OQ0j8gr2PVqX2aRRyAJQ0RBezAVayEe
Q4KxecDNy4pROQfLLGGR022Wwcuje8+HkcBGPhZ0NjyqwIKrzw/BsndkLVXKdbk3
+zrM9zzIit2Rrpu6C3IZTK+XgikCOHTWjI/EdTgsFpbdfTkrtatzAofvhTzOMHbL
OonXNfX54T0+Ax+mqVn5HGIN+sXtRaBnEsQmtuHA3m5rgHvAW4/npvTdJD7CUVNi
79GLBmoKWRV+ROh3Xh3M+43Icx2Lwk9OhDqRG/CW0gOMFLoR8r7B7u/xTM6ICEm/
qGZ8V0oYoKUKCZY/UsLLMSSY2D2uyn6IxLl6bUpYmM4xwiEacLq8l/9Xi8+aGBev
LokLTt7cnglc/nf8myoDgz6gRiBuQbuELOzgFlWJM2NIYMcsQFHPok3rOFitNwSW
tHHjNkxZNHzVNBti9BDwr9VkQ1GwZLMsyhe08lz2Jbki9R7YnjQUx2FGQqy6aO2k
nRj/X6NGLHjBNdt494Ri7AFitd8/+nN0CrAf/ylHL1STgSV6/3o9BMhrUFfCQI1G
sf9qTN+MaGNwD9YBUPsUN2WlbzeUJb7/mGttk8/OriQIlDtTNL5WvKtLTBrttbAJ
Q3jUi+XrAfBJJXExVUiF7olBYONF8UYZ9mVU08Shx6VCEKKG6c4jMQOgdI58mDW7
y/LyEReJrJ1Yldj2Tbd8VqUogVL+aLB1w5cu/Ytkce83mu8pKjSCKRSIH5He1L51
lz/qN7bzwG3JM3MMONmsH5IXdBY6qL+S5hS2uaQD/o/Nn7hBiAApKES+EoH+Bt3n
Ar/1kyuS70Hd9Mv41CvRSsIwnh4W54u/35Oj+zMfVrEEnXRuixyaNhVA1a5bj9ky
00WsOPCrUkZoIiB9/SvfsLxX3b5JVTQBwKoAkDZSxUQnLlQKn4PALV5t/twI8P4V
r+F1mdPJ+p002037jObAQIV6RVEcyz/Hr86veWEwnimJmydnogBphi/99wopP0+Y
s2zKOlIbE79seCofPc+JjnlDH6TRz44u3dR7x0uLZ9yC99Ty1M9wE4ZB2PGGYm/3
Pgt0ppnXaXulnvRtk+sPFP3p8QPe8/uSVuGjWY1qmLyPhrXHc4Rux32z7EDJqisN
U3qLgYR0Pa/RkH9EvUrENtboG/FVJqX9wqFQvAXeGHGCk98Ha4NhIegTTzt89qHF
DT9+0XgT4hiX0KptbmSQ2jdwmkMiiSL3Ur037sY93S3fwxdv75qpCdCqsTwfGb7f
Pe44pDiQr1sXCxeU3Ix6K+iCQRUDBQv0bMi9OqsHPiE7frkgDRrtGajkaNmpK2Xb
n1ubVfSP5fK/oOSYthDl6c2pHz5veAw/M4+jwxUrFMLRar9p9RdTYs+lRl0jiF7T
0x3xFq4svtHMPgjyxmOiJkq0dCEz15AHzNvfa06sZUdLpq1NDCU+98vS85vOTxUt
szy1CI/X3xBhPASm2VqILUjcO87xYA+9RTG4E7TQ3iGedNtWbrOx/tW7LV+koOL6
1X1HL12BUz7wGftVEyGzoYzeg2tcdR8pHy4VyH9FWgfKSBGSguEAgQKXwZRv6AJE
ZYS++neiss1xf2iwdU4WMBCVnsytXuNeF8G+Ww9Ao2500xEqVU0CYpChBnB54g49
79pDzO9MgXgYnKqqZ+40KpvAMWa9pI8aVYM5Gq4V0960Lk7sfv8v8lwOU80B2GK0
uu40Oy1BcYXB6ApBLV7coSXRXu1SR4uxwaSZ/c8bqdQUn+Vj1TK+hAvhorwIaExv
FoYgfG4R6WyCX3TyBxz0WfFGPwwfVgLTQYx62nVJo+hTfO9Hc9ZAI/J6Xqux8df1
86hm1xl/r72KTXf+roRLrIgZryazcpgmp6gLcrxBkfflKg378mLraxP4lGHFjaJQ
z8dLlSSKqJ/ks3PBmZ08jXzTcH36ydXU3qmySMlxW9G/IdhLsHxTLtoSEDPxw+Iy
WwFVhKK6z7uRtl+g3YIUlvfBn5Be3XSMra/e2+aSzFMHPgJ0p1SD2YU/R7xaX8uz
1O6j4yhOGu6kCYji3vOfH8zaPPi7pFicqnqssSQCtOtupXXr7CWgduk/1eMY2ZA4
33q5VhBfBmLRrQ6ux+RXaQgQOBx3+f8ErYeYkP2Ap5lqNVz+Y8n13v90uY98C/fR
Jl2Sc39cxsGBMewBsXRR/my4JCVqosnaYMCKWAiUfLWtDDE3b6vSP9lHyQYycKVD
umEd2EThmztPYr3dygOLWGA6T7YDO2RDLJC1tiyaVpoTVEkaHlZab5ykKPAZque7
yS07ikS0UmVJ22tCDcpHJYrPj953rhrfhrL718gXltQPrgFNNItpT4HUMFUrodsp
/jSCRpzj6rxlY78FA/fQvKVn2c3CijHe3MsoyCHOSubgye6Dj0ibx8LRoGkrowIN
nwp/quoxM7sXGyTCid6PlntBgoTANaOcDSQzu8OzOA1fijNVxoFYIUCaKMuE/X/4
/74CWzk3peN9tNMtaV5mWugaeMRkZ8euXVW+ScVtLLKyw8kw3H2vQwDvIqD/wxOz
MFUn7HKzyHALnuzmMFbHFeV+ds5EMkfoBSh8wxfHcxU7RfMTltKPfRM3p1VOLmKL
VDaneRpyJSfJmgg69mscSDhR0ABpkL9nufJdGpC02B+44PNHOsb5y88iHPWVpuBU
QJckN9oK0MY2cNLnpB1fVBDb8/IHaI+ndI5NuAmdynpzHwjR5UUuiwdA2Bh+AV7/
fCqg20lOzGGhO2UR8CmGit+AqerI18vl1bvWRVApaWHjUY3bEtyNlaxqeUwkjGAd
gvKnBGJgDIDiJGyoqyTXAsW8ClBGRe3AmLaPl4TieBSVPE9sfjE2jpgqtl2gN4Ix
Za0TZiGQpJEWSGWnHRsHmaF/toF0rfpfq9HqBAKNeBZj0xtyUmbCXHn/+UDhFQnb
ShDNAMJFpKUmNt5xtqzbwbxXSEVh4bstGs0BxGAiq64RvaIH/8mtDG8DnMGMDJ2E
vXLXmNnL6ngRO3kEifZ4fPboaAAjO7qiupHpqp2XENflZgWSeMAF5Vvol2qzBUbk
H2fBP3+f8bHZT/mK4Cp57opggroFOvfrdY5BZ1w1iLepTaySn4KGIR6sQcDlYFo9
ga657MHFp5JRRd0SwqH/8tf8+f4CDuQaMAIgKQk2V3WaN4i2hUWL/LzLuQPrilJI
0xoRH2w/GXflnJHAwKv8G8mJc/GJ45+3+EIh1WJaNnCWsATQqSFeeLryhzeiu0wW
8ipWEOkn/Fx6rhzY5s5/8bc2NlDyez9eet4Rlp2hkTC4bJpmHfrLeG1PxnU1vHvl
r2iRlZBES88tdKbCivt/BdoaePa/aotq2XM+4b6oB+A77ZKmHop9d4u8h0cAxaN4
gTUk4XTzm3BOfOTbYYF+AMD9wtEXQ7dntUmGH89HT4oz4r/bxkk/R/hQpExd08Ti
UvLEr9k08UxlbDgXRVBwRD+OKnGx8qHqio9+2MS2i09q2A0slxcvh+2swY/UoeRS
QpdV7CO5Ew5MluCTIbNJPLR4RAK8GRZizLn0bdhDwQymeHcX7oOULG4YiqgpgfcA
Be4sDR8af5K3ebNXd21eYoBhElc7LKcym7oPd4Qk+Zcz02mTWutLHQ/S+RcW7KhF
2j9geZCSXxhVuZ0NFSZOWXcEHItj1+n8dXnGFnZMBbQz3iLSgeeofbdKh3wwmhmY
0aQXUdvvNjgBBT4vWj80tlBE4m4QU0FOCKcXWWeGfPUTEwCTll9gC9xiGxi379L0
JSsOe3sVbBxl7iXLe7bfbBwKYCvvBGzkYjQo2tww1K6UDwIRMixQoItYDlRQIBs9
nO25kqyQNYbUQjSWy5uBgbkAGhSEIAz94/6K1B4Fy3uuwiKnOiWFik/yIwA+p/xN
mJcySPs/fqi8m6DaDT685jxoHff/jSapvPDmAeU7Vw/mx+bnK/6Bgc1OB6aDgb4A
Ou5TX87c+cW/0KarzHvaxvpkgbEo5422NCAZ+IwZ0zatEf7rlH1AjdfngD3qiwO8
EaDEDxft7ridIQoneaoB8fa7pmkvXrjw2ryoqypEfoZZ+TQECGdzvJfX0XSv6NH1
rx1lS21S+ubmME406bwF6/o95apbXK3Z7fnkO+Q5A80ZxQfltOkyD3CGCAtVSoSt
oMbbUSq7wIUDJ5pemmUGW8/ZIjzxk9DtxTVLVtTR0sJpK3mmypmSsNoea4kgRD0C
qt4Mav3DwMOvVIabl39x+wCny9NNN17bBGFLemKSxuhtqwdNAF+7J2QEmJmrE3zA
6zI/QDOHGA4SXpMQBs+4V8DNGgsTdCwpkbK+tLx/Ahh4U2+UXZzOWKGH+JExy6nB
FBvq5AXOKTJ8ZbHwLATym/P70QzcSUXRLqQUAVxWJfnDQPUn3dWK9tXoqrYdYOtW
nlB0IILkoJ4W1pobRqniRfLJKK0OsyBPswOGf26aWIfXYc+QUyE+UAePQGf4ewdE
HIna23Bl3GcKFiIouEXuDzeOgfmCCZqgnx5582p1hHS97Yh3bX7bLWam2eloGzTx
nbrz+eLHfHrQL6t95x9nR31qZGT1y17F0MtwS5kXXkA58cRy1lq3pApTJ3/Z6PZk
v6XS3ssm3ewYTm666H5yl+zHf1tg8JaVNMDcFGP+ZpD3/pVFJMq0+uJjLVP9WxM8
wJGvy7zmElVmRLCuYIb9j2r/RixWsDZBPKOOWnhw4o2JnM8qdfsPE/xosYKhnDOO
U06pLYce6jgWVUJoZ/Kt1yUVoTf437+1ypyiA/b2/qgive0wQrKaeA+aRiXI3CBW
IzOSqVDYlu5GX9Sh0nvEndBcBvn9oUE2jSF/YckS6cLTiDHiAY/LBoo32M4gTvLM
1eu1/YRnm1Qvt44yOqS0/iQCKU/0d6e9q6wFbgYIluDijVjFZVmB6G618V7hGJbT
OJf+OCTndOj/lLg+R2mUrxEO3hrPTQ/HpmnelmfHqC9/+lGdI6Hc87zkQgxfLBkB
C3D3LUR5EEyAbp/VE8oNo2oLbQ+qkOyveJ6UaKeeqZwcCWcxiCA9pIYorUpf9cOt
ZsxnPLWl8/t4dxIYCzF2HXPWqvuaI7ufRsXyjNff8YHiB8RoyeOel4x0Ihs6XHff
assTvpKAJUm14uZx/C4P/bozV+AO4KM926gYuBaJu7Oy3/rX/eD1DGIsTja2fU0J
k4J+zs2ZgmW0Lw0v8Rr2JuTs2/seFGDMkjL0BkgBlbWqddhY7/Us6ROphYWSZJli
N/J2NucLEWVkAe0yWqZ2OMwnTUqthTUKeCVvWvEjhM0zcLtyqK0/rvWQkk1SDRLa
IpzUNewcwPbq35ykYbg93CCNAIxiBri5yeJJKxBBiZtMjlHVs/+aW0oq6G3mHZgR
rwjF7Ln2GTZfDUwnIXcE868NfhvclPB3CYhRKT5Bt1rEUEXQ3eoQmsnnueQABAnG
KnO53CbAS0DWziNn+u/q8cB0ayLsUCyIbOAtC+HmsR/vxtoDeoWHv6AT0zaQ7ZuO
XIHjqpi0kRMH+ii+hYZmWJqvoMrbRxGpnwdOOophLiCgFv8Gft3vd0qln+VRYz/i
mYQS4uawMMcZ5mcoFLnmB17Hvm9sJxRj634pl3db57fKb+fqisv9UTbBv5I+/+9+
tlrCIuV+xouI0PiFs8XuL4A9/HIgWI/mIm/J1Lp6mJHX6x2iYGB4LDWpXBdk/AvM
ocg7qUSRAxwTpaiP4BYV5q+Bw+BxLWdqLqwGe0m9F3kg6SX4cYWskHQEj8jsTKGw
Bnveg6He9hmwyQXG540j2vSC34rq+iGUMLm1N9I8da0ZfGXATnLjt9AatSn9vR9i
dw+AmrxCI9PFBULqNbuPeNi4cBvVJUUZWPMETmn9Rx2Tpm91oM/X4e3SLMfddr1r
/knHYp5tN0fmUGXZaL8xVUR8TEqAuMU2ANQT18v1qq2gwQNmJ09SSuNRsC5E258+
JcyIFGAVkol2BD2c7cOW3z3pbxaXZKIA4dgizeBy2b+GWNGRWygbfgIKCE1upMyM
gXmQoWynugJyEF1Ojs1GF9eJzsnApGCGBe/R0wu0LUPmsgBV9H2vKO6y1HfT3Ssp
oC3p4trwG15kVC6e2QQTbminWNdjIIJ93jR+SYQ6vPBBib7FL7ruHh68aVxlbgx+
Rwb01Q2SMQZ7IAyPVOK2U/0FXpeFG3IaqLLpoYg1FDLttr+b/PiNGHAp0pfzvDta
wqdshPau4L5ZdB89qLufo3Fq3nHMKGrZrRHyFSEEiPwYnSl+2kQ3PWXDYsMJbcLF
p9HSXTKBR6nrLylA8hu9/6zQhaZVthxiEnZi8QYb45dVZT5DmuvMWDnSPlKJYY3Y
Sx6By7N/c6zpO+1SfGsh68u7Y78HgvS38F9lncvKidoeTDuAPA3wlJnJjtH1XI5z
L/Z3z+C8tmDV37wT1B0vbJHB6NickngMf7a7OrPlK5SZLYgaAtyXsw8MED4dI7O1
JMBCCGf1aF2nxQrJnGP00eXgz/9HuNoSE5zS548llA2heJYY8zgwEj2BvsjA4P0I
EFvNmOQCLiaRlhbKPN5LLA7b683Fd+HPEknDsWxzALyghS6t48onSQWBaLUSXo9w
c+tCC3dk6DmTWnxKfuOqrmIbPlth2O3/cQndaWsroFlflaeEcv1ZZ3mAMvvGPx63
DBqsK6mkFhWuB7BX/8VMD49ni48XO99VgKDtUZIqxLNoCWt2i0CsrieQBd9aB4if
8BR/XcaQZmVOqvGtQbAmkWuOMZqdN966HxTNg6mqWHjWU9xFHDCqc30t+y36MWWF
XnUIgYBqp8YA5KiYCcurpPkVtpBiyZz3KaaFNu8q0UFzx4w1LFfQYlxPobrbqauA
O89+ZsAi/WeOc4JQd8owfXfrhlcJ8fLdB2hbFTl/I96LP1zp3a4PN4iNNYseD6lV
rth2LuydT+rqGDIVSN/OAlc8peKRfeAh9/pfCSJQ9V1okS7BDnr/9xmgtQ1YRKtz
xVlqlfvIrdshnKjSonJLpJJbbup9+NuWyGK7XEQlFPFfk/vsRtCaIvpfWV7TkEiA
0Cag+RafMyA74Qd4pktXGtSAvCri+9LDswpy5yhnmRQlieDNoLSqKj+ac5rX9Z0V
VBPBbOjnq0XsJ6dQlt3sUi4NPfzTlChGDR47pGQeA3fPM9YmbmhJdfUPzehyV0HO
nb0yUtk2UJ9HkgKEk33t0ywa7XiUHVFx1mi2xPENeOurHeZpHlCvylTInuwgTbOK
8debxgi2Enm1zz2tNySbvyQyRZwfZPZt+rQ2f92IdJkgOcI47zhamMJScXJJgflJ
YbSCLtNuhdUlDl8LLHVxrCuW6/kbg9lEJ3SpWvzsVZJ7p+6g/p1TiO8tSUlyOpX0
b5VixK8Cu3Bg4OudzAufc8kiMmQTVEz9VCqW/jlG6MvTXSi8NnNI6ei4JixpOjgc
Qh/daNf38Of+IXfPnbxv2X1kWbXi5etNthqpL1Zfwc6FgFB9nfqOCYQSE2te6LW+
5qlEUdBPiIHAOBHN0n+n4FKacLc7N8KTRhybWeCs1ClSx3quy3AGBeA3IGxozwN2
/ZbTEmKIJ2lYzJ5+Hw2BVCane1ZkVyoGVZAdhi75kJGnSnjBNi52eqh9Y+Cdc8pI
p3sPuDsUDHzLtD0os5zGZ4eXAGPFNQb1gI4dP6vqtldukdQoM8t/uwNxq1TvsXvs
I5+kzR/o2wAQB7oHj+6o9pno0B6SC6f1y+My++eKCgIUpXU6I4KQCuTBnQzcV8+N
BA9rJgVvibLyrctINc1q1/1Hpkwx5dH1AK1UBC9ttrUbemMqJkwEqAoq4k286BWZ
aDZTLs7Kmk3tgWDCSldFtpp58/ZC2Ls1Z/orlK00Qp/OZ4DpyKSWBNIyuyyX0hio
HmkZNRvfvfpPQTo6h8Egnt9IeB6bfbQGShQ2LZ7XAn/Y82C6fOrFdBcXWgBXB0p5
6wu/1MN4ruMRTHAv7Q6sFyPHInE8UV2HDSk7/XLSWDdFWkI80JB4GD/xvdSkp6T6
YxK4pW3nvcYsSwNcp9T7KghAP03og6g7QZZPw+IzInieTRb4T7mIn2uRV49EOM2a
39BFMb9xRnH3ZKXQ/L5PGv6o/QLURR06H2QniuU+xDiO8wE37kKxkfII4eUe3RP5
vZ8ScnWCl2WDJV3fQXbMHkRdaT44B2lPErWlrM23qMVOpLCjytTqT1ysHAw1nTUv
rI3lh2snyDnOGMBSoiaaCTc6VTSioEVuTxSpC5bLr9Ww0K3hLmbP9VSuoSZeD+n/
XizQ3MqiZbIIxHt6o3YXFqhip6kW1NsRpPDS5eYIxIXzL/4UnVMxzFugn69VHB7S
0JlDZNRzfOGEkATRwQURAZZ7LALyYnIVw75OocftFmc3OzjM3k4BLron8faZUBmm
FcTOYcdASeaqjItiEKo7b3/YDs1Kzp921QFCnOlAQ7ZH7OcczIOakTV4pAq3R5qk
qN7qiNRGkDS0ur/mEkj6dwtTdTlhJA+reso7FFh8QXjUaoVQFPKGJEQ6+glUzN36
NIhY1K54moOhQVp1799R3St3jNq+wdUPqZIu9gor9GzQkIdTTgFGWIlrZPN4FFzx
noXzK/7WIU8e4M3sQDezukEQ+dkaC0DKktZ3vZLrLSCOSBQtB+055iVbT4WL/9LY
YMgVjSJLXHOER7Ic3Z+9M602XFugljQElIhl6i0rSpLDueoK9vjJM9dzZ3eBZPC2
bADAddMK4rTCyYzCDGKHd+8bQsvGfdLqtnATOwVTmSv1XlHLlDSIn7BMPiZf76un
I8iV+eimWVkB8ri+/HrVpyw0SmKFRK52BUVJzXcXnOk715aDm6upilrmn76qumYq
g8b0lreZxMM3QIexAif0XZUZmVhkjVw7Q6p3SsXUTMGhmkPuXT6NS0LChRa1EX/o
CMRq2iZumxDNkZnSkoIZwmQnfVqvRv4u2cxg1RUB3Ygeqv/pOm9ciKqM+Izwkc7F
r/WvssWVA1jdE7sTYpXmMPKQz6QtAWmdQb6FY2sZstkqCa52KB7+Rwl9PquGRmFU
kAZhQlhey2YwbWKoFdyKttFMdjVcAm04JiA1eMXQZKWkd9H6ZaWvwyeaZ1Wjyu7U
heGpa9EPVYTLC0vnEYrHeVgxC1/NFX6QPZCi5EFCw+EOmMuzq3mYITNyNyM4GbbW
za+4MYWRj7f3u3CDESvHFuIoKk8ghiQlo4TOfHif9F/KD+DHTkB0YYAkA+UthrCR
Lal0DPLD8rHzpj7K9cEDUj+Do7tAQB6CJ+M9l4zBV3jXSgacb4qhnN8Q30FEbfoI
6AQvBXL/cwJLTfeXvhf1riuHSgq6E92UbrA2KHB4BSP2NC098JYhfbEKFagY7JCz
SLYK30J2tEpVZInpKZwIpoHuWiB/Y/TXTRjNcw4nPtsNM5TntN4X7PfpZbOBYMdM
9ZSFPxaAoyNPMc4k5IwQyF7cW4PdxeIR1mq1i0OQ2BkhSrbrYA4a/l98ZadPSt23
7lf0zx7ANUZP89AcFHR5jBQ9dpZKdKU2y+C2ZjF95/kQYwgo35ZUegHG+XjykAb5
7pcKfMszT6BxSNXZuMsw6kQaX83tF/JPf5cpFpHtdm4tPeW+ugxuakZzJX6Nv5Ls
FVLMgNi4jS0/lAsAxVto//azE0SpwhBJeEQSBjObEGORhj79LqKZZgfbO8tCuKhJ
jWFAfMA6No5ogUxFBj7rpiT2iVH7BJXEUeXWsYWX501CRsuKczX7b5PeUzvbVMHR
LPNyMFeIZxuOsifY8Wf3YLrNh9GRlwK6wsjqcwY0A1BQPOGgYXGIItKc8J4B1HV0
0D5wN/eajHcezcLxxGWKrpG7NxlbGEIhnvPHCs3BJCfCpWluAHHVKvv3j//pfNZg
aH5RUnKisABPZb4SttixpUwgBCHMxNpIP2KvkVI45MOKBKr9FOJDaZVIFJ8hgjId
ZimmAc7EMRcuE6LVoxTftAJrWMzRyB1m4BccDAvBn77lrKjuOUISlEgeUiIuOIKF
9gBZVhtykxwOLqJXUxrOR1rfdHT3bdyJLG1WE2lFjMu7FCuUdx29wHtKW0d1tVv3
/T7W7wS8Nfrm3KQ06Ws/iq7WHm2f0A1vfv2f/d/4m3SKUmxdgOtY4m7HMsL/XXAF
WCtmwLqLpb1vvXoBn3NWud7BY3l1TJ3NzkiJ7liq5DfUMbqMdSs+k6j4KiKOz3PO
8q52isf5JeLmdxqjxP/e5udarPQ43Md0+iDWtxzKoqGcLajIwcb6ASVA+knCYXkd
57OBuI1F3siXpfEM3r1o+RgZMTLf9jh+y5Te62pTwUqHwyasNIAGjHUOJEsY98Xc
zeXwuDqHO/ZF7jLWhaELqNDvV2IjieICxOyIBB5WOM7i9dyeSd/c8vsX2dFLk54l
DhKQNlm8tgcHUkEswMljyyUwzDZViEy+A31EThA6u1QtA4rw5UqtlOXW2GUEPSoT
Wtw0F0v/VqdjVt7vP2FEEGj9pTBS/Fa/B8WA9eug2gMvQj4TkzGEntV9HZaD0oID
HHTbe8wVSF8xpukjHV1JXf7KAt0pItdnKPragSi2opQzGp3Cm8BOH18qet1UakRz
S6jbNxwB9yJV6v6mtOZ7fVttR6SjTgsgQDPwdw/oWnLqOCBLr19z0ZS8olQuc/yj
+/YeOs3ISlxNP4Fbkp+t4tcVV8/M2dt+8p79hInIBFfPZHcAMxTCIS00arFxtWBg
gFCzm445Ob+Cm2BSxBZsyJIMqfCNbtv1YcTXggjrhp6ks7RUD8560ZSy8hGChYVW
MWfQ9AwdVOPS0aToRNdMdPMi7KIQfb7cUBVrHln7YRlsea61bG5lC+sTxcPd2C2+
HGSaqXeNLQggDNyr2etOlNgbfOOAaSyFWrvnyXHchTPFRlHQhrfkeuLsNQ6ZBgSI
qDbc7FUKPlV9dwpkl6WPSv3tA2YW26XE6HCzHQ2lLtfTiyYoe+Tlure4e9A5M4su
Tpf3/NAmM4oA4BfvEi5Hsi1dL5jR/FS1nSZczxX7Uko7ikgkheFuYBOQRdZpfcXn
ii94w77GzhLK/CM9q8VhNJ35CrAubLag2AgbwTkep9fST2c66mqB2wkyUb59iR26
bjAnb7KpXE/radX6yWHGMUuu86FQ7dJEGwv/Eh9F767SmLfPYLFoHrNSNYlEZvuC
jnCYlM6Z2hhkBW9vZWzeBgaNM/qZws31foI/1xnI7MEOZo7ovUcypH1fhJY3REoX
SIP4w6Ipr8FwqrH3k58/mAB4wMvRc7JI3jayZu8/9D9oT2KoFUITw3a8yc/aXrwv
Xs+2Q/1DeEDa3UmNjZSoaejvAvP8s/Ox4h8RTpXGBS/8PBJRKw4xlYEnivTAWMmc
qZ0UACXmyvX8ABne0+fLIVxrUzla82DPueI3xReda37an3nFwvuZ0SGh4zhAXjsU
RYKUiIiX/Mo1iN5ydi5ptDJiJW5uURnlha2Pmlg5f0/BMQe2Yi+JvYxDeA/jjRX0
5oQsN4FZLfFRx9blydzTSim8cDvbE7QtGZtNY1vHzcKU7tKyq6apAESKxLiU2kZG
qVWEP1xoBE+8GWRos4VieQ3rdwMjZ0pmHifRhyVJPRQKJ3OB+gid9FEgTSoMwPQc
IBetAONPgtIf4qgWMqiAvbMc8Br6eB9rD+jwUOZRuqWsoj6kD1aKolsTzfe+wyup
vDtE+MtZ5scDoR+EjkbxaoVylUhh3j6bp9bw0q7SIlpO9BZ7MiV1dqbA0NuGuzMP
7mQp/C77ZtNxauZJG2nJhWfHijvrSlaJBDVjyzqHMBRMA7puVUcjhegc6FpJX0eU
qJq/f3jXGlhz/bka+rcVkR6H3wGib+3PMlLX5fhHoVftp2FSW+kA8flPmZc111qp
rERxy+qpdOpq20HqT9AddV2otjzah1xmUMi1G5w1hagJ1wGt/qPE4KEMty4PFW0c
0ggFchmDERhfOzYTaWuEkDo10CDDV9i5bXXqhM5Xq7HwbnwnH1QMYf6KiDftDo53
g1THNw/J+WEgZIFPxSulXJl8gtr9DcGpZDBPpq/XonM6YGCNeWqjkbJEGwZPFirn
hHZXPU0SNPM5bMj8p4Q6j9GjIgxTqyCuSAuwleOqnA9NM9th2DxjkTnz+1EdK0jO
W1jpsdRxObXXCCzpx8snGXeza3ZJ+C2btzZObW+Ki7XxWzrjhFQW9+XdPaIExcPZ
WITIyDvu9O71fnt/nMQ+x96ME42eDkKXLu2REuVRvaHFDiQip+MLtcgvCLCSIP3X
GTAT6RIqucrwhbAN0gh+NR5EJK3+ds2ReBbU5xVvbg7wwx7CQc5QKaa0bljJXmOn
xwv9H+9OH0XdPdlbt3zooo0tcc1SShjlSqKPn0x/xA52/WKkmPrBbWYosuZvCRDw
q0T97OdcziIYwfmU7CyyXv/T0+s3Hs0V3IXXb9t66nI9f6zaU3Z59hdhuFG05qlo
5ym1StFMDG2qVmxRNVTx4gjhfta4yuYGutC4Db20Pv7Ah9uXvex6RMpFy4UJR07O
m6sgDz5o0iNCuxvjJL4JZ/Lrx5B8nFFotvXMMCYvqh6hYZYvma+avrkhJaakgrqp
zLs3WmTCIa6NmC2gk7XgopmK1xp0AEdvG0MrIlfLZKxRBr1jN8w1XdxVIC0n8DeR
AB1hwe/B9HCv3u7LDM92kJWytOSiAB+pTXQF+XopI51TXx93vJzTcOomtHlmWBc/
6seR0F4mIV30mS0dhSQ08dR7qRNLhqkhGG2Bp/vFA/EkfowzCvf5MGWf0F+A6TM/
uqehBH1XoO+nmMeQFvJAyJd5XamiiQg3fdE8jo37LklNNbSk+8pOhiCZ5XNd3pe/
hThF/aG+n8JuoXtCZByyH0BBm37qh86JfcKkzMXdNlxGOmYXC6zutFdXGJAHMej3
uC8nvgnHo3s/7pfG5U0Yv+YCFKJ8txYVcyfEd93dK4xcXxw3WOjPBCs2Os3hSkng
puq6NPRJPWh5IUB5WcbfOHUrBLLbSecQacKg8deOvn3DD4RM7qmueyxfvBWjoTu5
/mcgWyux5OreWhNY7qnuKvxvOVaOBDKSIyqQTkYyyKRO9pAwZu/pNA6vq16jzFp4
5acxV1mNUJYv6Sbx7zR4uhbIeByEubcWpMGwS+/qwCTayb8xS8JdcUlMLJx5onPl
D0OtoJcJyfVM4GaV3AavWnZ9mcFZdGOJfCtqOE+WzR7UN3M9NqGO3YLgs6lYf7We
yZak7pPass9f4kLIt4bbU+jH36BXFLA62bi5EFuZIUznpzD1Yg2xdkM/zt0Zx9zo
O7KO7ab88iL9TOb3JDPJOdnAh9dZSNA4CRKz4pfGTp6zDEMBzgFNdYADdllO0cXd
uwMisAqAkbYTYEjhN21PUqp7L9iBJL7HU3/kjDNjOLzubNhY0tOwDVe3ouFz3nEC
r26RAj9IjYwE5wY60asZoLgtukiQI7DP0jLa1FV/9ohhQMmaVSmzv0vdLLpA0TJk
+O+uhPEHWKPcIXgQLGrVQ5haVknHWCZwbj2vK983s57glBVcl9XadYmGpYuvlcLp
TJykq2k6Xsy7uB5q48B0JlDU9IdE7sJQhR7tvmuRvCjlUqnYrLu1dPkstQO6JVm7
m/ygXj3NMLvIUK+VeysZGf+28KD+V+ouYpV4IWWDyK3kNQg5swhIogVrM1u6zKjL
o9t5CDCkZrOgwDR5DAHFHaOMxI+C5e3tbtXIn00NJ44f01ohnIYtEz8nQQpM3TFk
H8Bu2aMGO8LNyJlICY9Xa/oyaWQOPOYfrjXwILtSTMiS7uS/7VFJjtfVWMQt9rlz
MGWWM95kOyFP9gHree17t2/Zyf096CSrfyJgNEmwMDPLYkcT1o8/kbqLXcqadVQV
rTrcLSgj71hX/2qK2Q0NjEmWWORoP52QRR1MjunOJIytW7snIShrk32MMReLcyuL
HVzp2H+TYLe5P5IoXAfhvGtsm7oRoxNgpGtiMO8ryCS9pV/82pfUgjbKOQLGsDd7
jjRwvWp5Eh1+WEmJsqKsN8xfcO7PaKiylFtx1KUtXSSWXFxwuaEAeY60URA8CTUM
EEI/y/098xIEkADzuesm8s9Ua56Ojmq+LB58NSGDGh8XuMf7KearN5WfQxsbBFob
foco3xsnIiFEj5uKyz/kNma+U4BAToosP1D2QFgCKyVbLnozcA+1sA/fwZIW/+pj
9lWj93T5RlnU44qqafxUrIBjcOlDIidAsUY9CVvo3ODgU1izbPVijPnRb0zM6vO2
1af3BQWSLxM5P/5oF59lkkhLcMb5mYu8RwhILFLNH5wvbReNpLV18iIvMqV4Skgq
zpo3RnU6fv6oAOB18RB8wcNZL61JFwqpsa2/OBH3nbNiSrAQYJZ/xxIAdI3G8lvG
Tb+Gt0PRxZmieCYLcxs2ZYP8jCSzMLZg2CnblxX3uPahL0RGkMXJxnzBxPfVLkA0
YezA0Wa0udoOxqeZHrMj6CjdmK8ILPv4U2F5iVowWEr3TTkhwgGGLGrlAMTfAKLG
AStogivXpogKljoblWcHryONYENBrxjvqy1CRauJ18KbcZNzG9i2J9CGREjyWxsJ
f3fXO5k2/K0nuQQsKEGsKBi5n/1XX/fBZQeGlsjVgtQ1d9JogpYxVAiYOIb1PFlK
vYp6TDJ5fpbMMAtItb7JA9e09kGKEEwE+fptBByDEULQOgYD3+lKYmwSgy9erAur
jNgZVmjy4hRZo2EHStF2/8x/5qM7EICngdrvhcBqu0NIKqEIzwQpTdyWPSLCbiWW
42MW1bwiEzxdjed62VkzSrqqoFAjwEsVdk0yNhs5gXGc2NogSukL5bPH/nZ4F8qQ
RG7290pbzHYn2eXBZe9F7NpXrF2YJeCH4lcb9xg/JlDGMDGbhOm4xVYjs7ThfS5e
D8h5vZ3wqmz1QNSlZnLVo0v8UCafjWk/3GZoVyzhpJIsDi1GOoj+OhoaLt4uuukk
BK9P0HrRhIGTL3cTAZotOy57cecQhjsOGpnWqFJJQBk0nTOTkPOy7X3FJvs7OxQX
mSqn+uMNFkDyba5/zD8OEDVj7yCTM96BkhSBTtnBWQifANXLxlB1Af2kLo5qfsD8
kmKNi4KDiXYF7JcCJNZjH1xiksImaWB92JS0YGi5xc+tRyl2LlzTYNyb58nBVA/0
GIa+shQCktLV4RvBSXERpQRRqZhxNonfqhcYY+spb3TGh2wN9kTGCqSI3ZmP+st4
Rjc6PtEPJo96fqEYGMJWZhIF9sEvz1XWJENegAYRZdGRjSX0WBj9rvQ71ObtxQOr
jYPcrvJih8s6WijecYNycRY+4IZA3aco6ro5yen0YMY6Uk5oGdeeGwNz2UF2ee0P
fWtO22LXlWlr/EbpJkD1kSYmN8kbN6BdTYhDOAr2K6FyxwGnvTJVi+TvJDgHrE1D
twfQyaYIqCBeSchVIVhaYS/zSPGx95ydFZ3EyorxQOPvsV90gVSYuyE4UayJCcz9
528P3QHJnhjjuf+pCEIfav88TZvM3HLXLn/YKocsfnIBnY0e4MkalIIPlhJNjtST
Py/NTpsfNu5zbG09HSgKEcx5iXgbyhPbuDgN1jh+C6F+fJX6P+P1e92Ww58+iJte
LqqOtIryYW3DeEZiUqIy0kMhMjEzDWqOH9I7gx8FjErEuJBF3TNcHESfir7Tq7D2
8tvvF0mC1pYaNNEsgwuJWU/9aKK4oRSXpdnYupGDUqnYFg9xtaKh7GDxHmKh6iQe
8n+0jOWmPXZeg+CSXqGhpgnZVxPIzKrPyY/X4DmG3NNRhMudZ/lkwNzRyiQAs1JD
SHol9Sg1uJYqUU0srNH0frab/hQhvqH8wuNRaI30NDUOjEKSjZoQ1NSgwWUFYPZr
YCJ5+DHHUfHtcemV3bEC0uSHULYr8oGPBNx9kWtd5egspMW9xOSJjSr5coWg7ifW
3PkzJBem8ojEvOiqi+b0y1M1L/kKgqQAksYsvQISBNi9RwHS58hCaU30Vqv9RbIK
C2NSgJE5tcp9t+2ynFlcphujSFv326gG+/kE1N3Pbt+GWyk7bGIbzTclrWGHNpOH
ZnL6hLPaZRYxCIkq9sgERoxxTsXirV+qEF21aErlswrftDuWEmv4h0v6Vea7Y2F5
z+0ONcc4cMXfMpZeUvQNAQKEQaCe1rx9vMZaZ/D/uRUirlz6IPRiF3IZZhzMV5ir
+XYkYiHttkiEQrl9p5fSImmq5BptbGQkxVN0BBTIq8Y0pnsCSKCud0QCQBmjZ7Y2
tkej0CswRmS8yuAEzFQAhr2EE1Y6n32yqwvnEegVNKmXwYWJ9UDg4IIIIJMz2tC9
0tk3Q/jZ3ntmB7QPaDZ4wwRvI3166FoEY9obGVKuBN4NkN+m1tmWibMi0x7ob6jr
EhH2uvme+5Xh9lMmHZmFXA6QTjgVTsHIvb+IUKjofkZszMoLqQiCIyLGuAWJLRB/
jhRUgjK87o98YAWtZ5w8pmKCcDql+TH8oVKPJ6fPKeWkofnZ6UHsbhb6aNGSPTCD
a2JEI8CixkDY/yAPECxYLYRQUaEOtsLnGqxZmTDf+xuZ5LbT6VN8zUDnxHMfs0eB
hPASQcvw0/Rnu9jEt8stU0CPRRMrG1820B51zjiCTiTahLO6gamOWvhHnYcBzrag
Q3RI1k6RF4fGyQ8Y/uSJMCycCy6qbUuqzwc30lj/8hCk+Z07aedIR0pTRZ3XAyVy
JKRgAkUAyvLlRA/pAlNgcuvqYqsjAWwKFzOKvjgX0n9DKBziNGe3gI2I1S3kGgsI
VvwaABLcLd0mfiPJfatIMj2I30crTxT25qLvDdFCRvicSL9aete7469dqyw0CMyh
r2K94TL3U8qphzMz8qir3aVvlO/umeeMQC1Pf9pcv2khWMxtCIA1WdfjTKamoG8x
TeH5MI5N0MNlBkPYU2xWmRPLwY7GdH/rjIEeJmzdBTnEQmaAsZWmoZKTfUZgbm03
QEjV/PHQZTIwo/5lw6QMLiJ7BvdLLdrPQHkYnUOmjXHODLV/dFL8fPz+aM1wXBZ/
LaGzkEpEIwo0JvQKAgccRFP8GTLAV5lhfB2Xk3f0hNRxk0PK6XQT2I+4xH5/+e0/
9H+I9hT1RG+IzMuxLhvddGwCX+hwSdKMFzQSjcVquRk4upFPo6OqmMdIx/fYI5JD
W3hEyK29Yrndyr2PVPcHgh+QjPrE4i+oF3DWRJMwImNAEyHK2YEPfSosoL7cpOwv
uPFgLjyekIMuGMhTa4FrLL2nVV797rlLBdeT4Tzs2EHjP8BCnp3vKFjfvfVncFNx
et8TZqhWg0GxOkxi0cAAA6fn+UmiiN43RlueCXUNf6kymwtN8B20SQfkJijEobwF
TuaiF7NXu6WYJCkeVrIyJBnl4TYA2Iwd7IqWgWk6gpLaZNEWd4+QWCU6rLdTIcHK
JU4JpmdZmYbgSCQ2gCRVJBsMkvtlCxP7R0NbhF2O0hdw9yMg/UI9GB+xJjLexq05
cBns08LV6OqomLo/OAjvwp4U2d5JVljQndlxTPYcotBxGK9NgiewJSXeNVJ1QXy9
nS4kdoO5yHLjygOygeYXVQbiempx9pjPhFitCdk1E9FFArrjm6s6JZTf/YYV1c5f
+HBx1oUujJk6midCeWJE0u51bToC9y8OhLvtmarr61qhnIDS/oIMNhpDJP7ZjMbh
psrWV/xBuXy+Mfi7euoSf6uCDEBdtyJYDdS5WBob9Fuq+9AvdlbQ6rS28KEpa+SU
HeNrgdFgf2BKJeixIJQxeohU7dbXvPoeox9ks8gtiSMBYdP/eW2joooNWrIIS1SV
JY9TXodTum3ELQ/0XX+14DJTKHe2Fab7tZ6M78YaArLwJpTwfj10nMrY2V9JADgG
8YZB4W/D/kIfwZiGa3OYIDv3hPvGXBMkJoQx8rWsCFxwGM5X7i9P0r1ju0FkrZcc
lElaJI8n6swVeipNsQfmFRvJTtAsgNXLmGJDfwYyvQbPzC5EDQJB12Im/nphg4fI
9D3tAM4TvXIPrX5t9h/2RsP16JpMwlwITJHI3inh3y5C02iK9oMQiEfCQTXjYyYz
FMWUI7GpfA9YI0FqxPTvKEYKUdytW3GjO7KfnrDk+nhjIb4sb7dNOQi1q7ur8onX
nRlScsgo4WcpmfvV5THadu9597Zq07vq9PUxnGv+JSKfXyEogUtWIwi7KaKcQdrK
iIu0I2fNmRaOOWqt9qEfuc2otGRKTxQtpJ9CIT8j+JyuvTpuoW/KknGUWTprcvKA
HWVwkNGNrW1cSEibte0BCPYIkiNl7xkiD9gBDD8uoZ71XCY99Ch2JiTPVRB8kfUE
23UM5+I+UVtH311dTnCJBrTjNkzmeocD7NsnKfcsrTqP7fn+JNw7HY1GavA+STgt
6JhNcfas7IskPd84hlLFF5fZp13Rx0+eB8F9KCc+MjDYcGb+zyZ9OBZKqiFQY7pS
mDvIx2jehC66cGm/kBjjrtf1xK/+zbN+ZNlhqmeSsBduHZjfXZun/YtmD03l9eIF
qxjBwnIqowI4mjjZIMIkr/Q7JoKd9IUop19sZZC2CUacfUJ5u5Y9ccRpRxRycMbK
rphq4y2B/ImpMCz0vQt00TJPKNupf8aJLWgjxmHNjbfiyPOJoAyamrZ7saAyNpuv
HhK9IYtLXj+zIsNpGFsXpS63flIdiYmMRrJA0tm5nnS/yNvWjq3eLzkVrIT2lMrt
1ZkSJMR8yK1ywkWyNX2oGzcUvVkqPnVX8Xq1feMHBwA2reqwxkYFlTM20fYb3lSl
RjLpdoizC1dXEe1WlQyOxlHEcn+WSphkRdd7c05xQSt9LWYWQWw90im5izSOVUNW
i2ZDaWsvuMhfzKPIbg9RWyABAVPXy6DO60T/3kSZqPtbx1zhnfMpyd/z+V+z4qSY
GVFCw2F2pR1SsxxEDB0GNbSvZTXXfaOJzpSabuD8Rd4GVvQvo6POmIOFuwEpMzwN
pocbpbIA1afDZ4ZsIf2dasPPP/FZKsKSPD/QIrn4wxHwZdCU1lVgDFcEo8FbmHKy
9tv2ejAWEtLQc6MGx7SYVO1cjpZlAODrbm4hUwMPk+3lvicXTM8lpZX4j1FcHtCE
AvkQmF7JEAtVAs06MOf/H2xt22WC/CkptTeAT2nOLBpOlGHP7MPQl6w2FwuvbdKb
uXeJwx9dCcHShIHszcx+iQ00Xz3R4Y1JrCAXKdgyPodD+Iz94OGfZjoDMmAnZHvg
UJN11iplASEo9x6lM525NpsoJhAhqHy2AuTXNKbe+54HvRB9lGZRsKaCKQAvTVQy
mF6pviYed8NyQXBQ360sDEmp1TjNKsh0aD7BD46/QdHN5OY4FSPthY/Lh6Vz0y4v
hM0pNMS3cEqnQLdWXWmO9xEUBRtVYTIoik5HPJSJguWMk3rLe9O/KXhsqbOOZnPH
+kiGhT2PcgC/EH34LpR/qhxG3PNiJTGlQjf39TAZNfzrqeiEDaCYQgZ1qbIt0ueQ
y3J2R7kcMCFp5s683DjIT8uyc8hXfe+jws0moAfKXNo8pDcgMfmc6rXTszOXR6lg
1ty110BCWC5nnh3+h7W+5q0Q29zQdV/coQlbNLYH4kpRws5X09vNLYbtG9oODxES
E7Ow819gsFUXuWNtX9QYCFdR2LGwdDyQN0OizK5p/+qUPbESYVcj+cFImkmJ8Vev
+Q6IUoStQeSsCc7gXx6v4S7Y/IJk7zqwnEh7yJ6Nq3M8iqYG5n9RD3yxJx82hO2Z
ghTHBuToBOAJOJgg7tJs8nXerMes+aQ7f+eboZPtjD1uzaGanGmEDST8Qa450CgI
q9ByW+gK1tBNCTkYM6BijaPyAXHEFrMJ3g5BSO2MYoIL7y6/VIgQ7xSnAWg7B10E
zEkoD7s1rUmzM1bKu76iWmMP03pOb2XxAuTjOjk+EVQylSMlmKoio5vohDMoK2C+
kG3VRq3DZsnZA6wTUNJ0oWrxnuiwoy+Jt01WgveqXmYUgoMAktuPAsFa+KjgeACY
qyqaOiBZiKLDS+0ZKQZ3YzNVGdZM+tFSVPnBTfkvwyuRjUilz2eEhob+K+MopcoF
1qiL+XKhAI702/b86oNJvpVi9BxKFqnQjn+CvmQtdKbcPEb1x5UhmYFeGyBkRW1H
OJ2Vtp6gB3KhqkxOd0PiC20+JxfsLxXB1SL4B0nW7rXPSglM8uka+AZ6rca/a22d
1sai7NkXw3MDpaLUwTc5+WSXhu8oInvmyS/dAECuYS/IpVkMMc2u+VbaxKV1zcNK
yPEbwhabnHz8/3BzUkl/xgBcqmH+b8wMxMU64eAcmipcnYThgi9oU/LqEm1DIs72
JpG0l+7WN0Jdw2YPlI40dF7bTMWutHk0b2FYHhGxuPBoHI8EgMz89ZHOEixS2/u7
VKPo4mW6H7K68+h2aNWDQ4tU6TWG9VGzcGF0vfc27PXZxn2N1jAGKeAXYBuYAB0g
KbGS+fdDfqhqsBP0kv39rARJAwzODJbTrdE7+9AYt/FYEhwf2FO2Aek3BrsY5nlm
fCezeHCHpOk7szhuG5OLNRB+6whK15fbHtvHMrHfaFWYsW23Tk2AuRU68H6QcfaQ
6/lAKcYOyja6W6ZQlOtx9Q7+PsxO1Arii5P+t27Rl+1rO22n0+eoc1ljGpD27c8e
E0mp9+wJYL46tOVIAJsLj7AQJidyGFZ6bi9G2tYWWxvrrAE2dp6VrXXqAJUY82AJ
2xRNZhfi8AwV5XCcyHg8wV8+TZ+hAIwdu40V+KzmtqcjXXLulAAYqDlOzyoZS8RK
2OrBQftmM2D0r0aYkGRQZa1CvGiJBXi/n9EOiFoNT8zNBnZ9kVQPr4ZPSy28Tczn
rtEgt893+rrGjGB1iZWoLRkcHWymNhVnD/rFQWO4PEh2TxFak4w8M/+Mh24h+wo3
CKfU2O4mkbSJG9wgq1vE5LxQeaD6Zb8V9vqPDfaqlexwz3Sx5XQjlTRS29yvMQeb
EcKOZTxqpTLLMmm27wolS9u0yA1DbKChQhDCfZS/0lk919Bpbd20hSZhvDO8DiIz
XcV1ePCWdOuJ7Or4DW0rBXvw2Qbd+7YaiHvi7FH1A8do+HO/jIj1YbFTev1Aqdn7
rbB81btnfrPsCqZqC58IliIv5du36DJBy9UeUa3KTVmP5m1O9blBHx/Jz0KuYOoV
iAboNS1z4RC92nprhM64KWO+erBcdFJ2sFgjCWltiyP29RacOCY6Da6MruLC2E1N
rE++MZkiz5xIvO43U6OFM5Uwownd6UtFzm3Su17JDKfQt6UpEI6u1rfg2fnn3znf
F/41G/3qpnBN7SSJsyg1OcmNT2i6ta5kmhZGLfYdopwjqNH/MKEQFJxCRXXtJGj0
cYBd7waRAF+btca3GJrMlsFWhtqEoUq+O4IHaTWRdwfgzLjLzY5FROL7V4071uRM
qbPxnowVl6ra9/huBWYTDZrKMOGYNHcLh+5aCBWjQTrbeRbEaXOAl71A9coUBKiy
n/4ElzVpDzftUFhsbTj6Usv5zKbnssPimQWfktzjrlZGNPHRljTWLw0WDLm/b7Bt
JVwZ+D+1ZFTR4WUrPJdfS+am513WlnR7amNH66NhE2pncyIlDHGqz4sa9M4Pff66
FfLmnbnlHsFniOzI98lOZQT9X3qBJc+Wob+ao+qXMHzuBO3+DVTMi2yklfI3MyuZ
/WsEApWBOynHl2Rzexjk9XHrQ1PvqDHGFaHtUp7oDCxskvBCqLDRBVz07XKdwxDe
/jDKkquT9NtFL/vtT7BIabvKb4n8vLQ8nwWj4oYcNDC+6YkP2Mo4JTKXaEjzWgTP
uEB7usVIGTyo7431cLffqGl7Gp0r/tOVue/++Qx22yKGfYOIms1hkXpt0G6wrI7W
nbZydXHHY9jQs2e9CTxykpepBYwIY3taflvHg6MFiM0O9r1GB6/ZCBY5ldZVIltm
FbsNtHqrnStaLMw8BDtzWrR7l84/2UxLXmzAShSOJQlujmcYF7SdWHnF4ZEvJn0B
o87fVb/N3MBUWc965WxUb8aQ1eplCb82dEZ1f5zCMqbE5vFt2OCs5NTvKxqiMYY6
zH/7LRBt9G0lnQfxGmT22FouAGbU1+CjOvg/ELQG8jUxIN9fyZ8lvRl7oGkWZJIq
lkZyPDE6pC/kcNZ3MKEeMG+9V5V9ulWof545047XntuSx1GIOgGFo6CgTPA8+9gn
bJysGFOTsWdt7jBymYcOBDTuB5nhVXp0cgwjAY73B9w9m0ZOKJzK9mumIbFv51F3
s1xibIDCN1DB+Yb3csBwnN1vyOU5iEuERwHj6S6v1Yxz6qwl3OIAOxHmFIEBNmQI
grkTMpTPH0wvLeCYiR25GUJVDuUPT4biaUfNLuDay44y/NG3E3Dj3u1jc9py9zQc
rpT4eX/OY4OyJqMqfpEoLxHpu6b623yGl16601IvCpQCdBayrTaJA4MBR/ne6nUb
0s3XXV6FMujmIrB3mClIbhNCBaNm5stcyTpREdvssjQSFlTjaWnAjbD9b58+FmQS
frBUiWbvlH7YGFntkpO2F3INRPi2rm/E93PXGDCyD01PPhHLA4kgQXCAQALNH9MA
ABFji8W+oD2NDwmxVE2JaBBen/m+8r13VUF0hUt5Cpl42BiTJIZB5B4qdKPLfyik
t/hJ0j6+vsyF7xioa+NFEVGoUmxjdR8d6LsazssrfqmSU+HjFuuaMRqYeXKOSolX
4f9U6h18Emwzqpaj9iWhGWoulPkQcM0AY2wS+Vpm7qUMlnEoYlo6JF2iSZAv2udn
PQi3wtdeehXC/7HPnXMulUTqyGg8MPeH1cvy+H+5qBJBQkNWCne84ofoIJtusc2W
jOXQKCSpmI0iHPJHmiV8gcQegLiYDwUveV37M4irHGYB2urov8rNxAQZqoNktHAV
kE38CRFaPO4XOow/QmNZcKjABduA3V/3xPq101Ucp9/B7glOGJNIqx93t9cl3rzD
BHRq+IWflbJBEgz9+UCCPA3EB4bhPRgpHRNPe1gDxSIT+kujNGx4MVpliqGcr9LD
L53UrL2c816rwOpM8jaRXDQnf0z2m1fuPSQaQx9Ou9yShnB2CjBEP0LS6cvUYS64
NttlzGJ1zuy24tTSGbaAHdkujSd9ebIPtr8nrWvh2SlzrWSK+eHlRyfPvY+/1O/1
Lor75AP1VRTU9bKTgaXlfQxN0gJaN30PYnLvFuXBPN3QYrJLE//MkP5Ydz5hUVcA
eFK9SmfWnLntXtnflw5XSB34PIoUJ3/xIyo34bzDtl17rXkaoJm06Hxa90CwqYvn
PXHf8EKy/jByqti2N7VlR282kHcf5rIdlYlRCfx2WLr+8hdcdV2oI489q8odvtQO
ydlAW/AZPkNYLsXDL1HBK78W7Msm2XSkDekiAKoLliLdcQf9cXBDOKCjVH6VyNEw
QCq+0MoERJowXd4Q2aGeE0IP3IDFJWCTFCf9V4pC29MqTy1O6hF78atWpXq288V4
YuR4hm7BDJ4YphvBYZXgXGrJOuga56gkheSpd/dQiQ31kwYls91Rgb9lOARlP7p2
kRao2eJCjfo0VsWDtuSC6ntz8Gp7tSngAF4ZgriyL1KSPVuA7AxonEh9GIbg+P60
XKazGo/Bwxxm0GuZe57NjcVUGwnSRjcZDM300obyjFt+pYjosZH1UK9L1KQPu48j
8sUISHUuHr/mg4FX8Cjlc/PqYFLd8I/cAr3Pol3Xl4QJ8Y5kgCONlJibeKKnsCAM
SuiTztQFdQNAhncDpWQ0yckYQ41OkaCCe96vs8VKbbpOOU7D0VaNlZRNnZmlzZnN
QuVPZBdT5Kl7oFw7tRJoJrH8/ZadJzbKvswpNjpxlpc0cAwWA3B3JgVqpBVo8C5U
4Q1iu/jioGoPaTLwoZ7frrTnI37WVFHnIHH4kVd6Q5pEeVRpepBVeuBgCDESQo2j
+/gNrtPg40+RGR3tRWVO/KVswEO4WrFievH4oY2Hk8GTJDq9wKrQQBWNApcz/7tr
oNwX3DT+eXoFP2LqBhWYdKLKZWn7DfdtbDBK4yMzoWdZgGc93T6Y6rTQlW7Pnldq
55zlsi2wGymLN6cWm8VWLKK17UNd+NSx9gMtw8J9ipBVCe7qXpXuGIpUbM+pV3+U
45jsFTh1Hsjg3b+9XfE8u/OWaH9XO3wzCGTyYm/8wbFR+Lid0vU5OLwiOsJoCMtN
+qaFNwRL0pR2DKM76HXlhTYo2OlZIiDjza5pkjuipQv7FxhcCTmkO4Pr52uPyisN
N+Rrqz4hzDjE0uF/x3r1becPw7QLGK1aSYWrHgSq4VloYZauPyGVIDs92B9lg90s
3cqLqDaibZ4W4xBefq5rSTfaSi0XFgVAeqwtz6xdgeWY5eG63Cru8KXhXBCHaDDW
qvFrdPGjzZOZ0IESTDlIrTm5R1CaOtVPRYg6M+nXG1gKtzVISx0/qex0ks553coX
u56yaXhhzxeyzZsUbsBo8U6Eb9/5dMEQPMt4HprGHr3bAkxzJXkClvtqr82RRdOX
Izo57idvHchMdvG6HdVBbH6t1QDcImC1UA/9TP6vBE6rbljMZCNMBV3fhMWzBuis
NwRznyVdEw6PKlJ2I5tkIOTQMBbsi1ozXwCZffFE3P9u9hxgR5sW/PU4UJOa/yOQ
LDOjIXo+OUoMf6aJGv9kADBlslDjVgUr2VwMRDchCApcqQ5xRm+THVhBke2SAFI2
cjN9aOcl9Dbek8oBY33/EF6ozCzcm+dSyDVAM4GtqTRBq1oUki+6oX2QuPIZRFeQ
2TZ/E+IMrj9HtiG4ecTEcZOl1cc5I/WMKyCG+JCclLAOS1Q/QILAnyP9pAoM3WlP
RTqGkm42r96Uqh5lQkZUyCOgRi5O9xy8xVbStp610Dj13Rr4ZaFPhK7AQEQt8PXc
aTUrQ1qkeIEoqHB6w2SviORz7/aYd1xOpKM56lNTByJccZNTbYdklOMKitYgMUeX
HXuqHb5R99XwYUeuMFLXVAFBgEjPfJQtHJP5ZvONKhp3mIJjjAXUrlxXLMmb12pa
YiHAz700RSsSjh2a+7JcVe2B1dAO0fF+uHJuqtC/ttlaQEYN9VpO1FI1Nh/podiU
NNC3V6VLYSQfAMWNzQ8DizUQs10SlVIXG/MN75oA/JhDCDtiz2HmdJEuy9TvgRGE
5d/2t847GsSIciaf/eM0J7ur6aKXKRg0RVZ9f1Az2y0/bFHjwuQvlD+wYx/jCVFj
wjYkXpGifTzm6IDr1vWMPmAdxfEbP0q3HsRUywOxS1v1gpI5UfOOKitjIKv7hjWQ
fb+VCeApn9LfsxdyMdhghQsYvsFCnG3Qaex9a2veJmdBdGQGjpV1nmaM/6CRY7dv
GcR9khTYan8UghaQ9n9YoBWuXZB5Kq8OYtsvUSURfulpiYdefacSOvpTzsKOtqg7
5hLAILFAQdNcWpbFRI70U0h5jB3vdpjVnr8MG0b2qCsL80n4xLsp0VQ1WMPcauv4
GxoLddAvSeXr5DmJWlbXpwUyVxRZMS6cX6WxBxUTHDpJLBqRYO9ADhqIWU9GhJl4
hEzE4f5LwkiuFL6TKUcp2AAir/frCnu1Zgth/rxjLbIzf/P2uAzUN93KmBxTwYlR
Mlg9sxA4A7xZvgXe5gCupDaKA4xY+NT9EX/6/vIkSo/txaKytAUr9qKaiTOp3WUs
JvADacXragmOkaRlEaZKB2p6hsbz9+hjMRSpeqImJDTb6ZhlJg5TjIGvjcHozmeN
rWaA5BrcM+MKnq6j2Des9RtU9ZqwQJHtjoZGL6dn9LiGSg0iVynPrk0uiqc9D3Lu
OxCRZ0FqSaUChkL8qBkl6NWwEcghYWHZyMo1Qq7h0H7haVQVRHnN6fMATyfbVE/e
COvwJdGy60jlABeneJw8A59+1Nb2FgzO64BcidiMRuqHxSJ9m2Rm9xeqZPET5TLR
owNAgHlRP8mO99abw3Ok7PzlM1ifTvhA1UrUbN890RhBsgqXUJaPFehBmSRwXIkS
xWF9eb1QQ+R/tDcch5YB8RM7zu5dWhtGqnvzKbSB9Y4Q77VjT5/fkbLlhZomonI3
rANB2BRpLC0AP91mKJss9hSjic+QGQOsnAu2jCk+0L6BrHcZW+HDNm2oCbs0N82P
LldASu5iGqRvu8R2DHNZ/FDYhCwFWNZH+NYLX8w5aejOjNFNvIXQYKR4ZcsXNAH4
IBrTxJsirD+GOt+aeATj8f8tXCfikug4mGN4/2NBVjYoQL2mEZ5WjTpjT8HJOb55
TfP+8ELHPRw2IRhy+1PowHsUQ7PjsiA1YOZEJQ+uo9apGSUARfLGq95x+shXAIcy
76Jjh3iSZN/yuLE957vQ+0dVFx5sDGAfqiI7kOAxX4KWtKtjBmEw7pm/zcezygR5
vY/tW+csDaFQXiNWIEGxMj1bHlam+Zh0KxU93To+8+EK1R8LRpd2k+2m/zTJIeUI
Os6rzBxHyBD9Q6ISfED9qpbB2e2QQsXhrpBd59Ywy6bxcPjMMcn4T7fro9vN2TMo
P2YtZJ3nagyRILRVKUfzj6CVtpAXZcxlU2THrazNda16nynrFOvkTi2jDA1cqh/y
nqisVxNCqDuxinG316xylbFICf26xkZ2iUKawbXrBqOm8Z7ZkLoRGQjBYKKXCefo
q6lASPS+Vl88pNlD+2Z1hKhxnKubcgcWAQV9RBCSlWdY0ovlraUmKx9n9jc9+BFi
pCvELFiA2fs3+f/2mji0/wgMo1jvbpVwwv7SkCC/VZTbWNCelaYv9NN2YUF1I/Wv
UI8+3tDLOXCnEfYDWKQPAkEOcoinWHWrSWM1SuVvedSNY33e4iWjc+hkKCiDLjN3
28h+VwXWv+P42rYofPpb8agURgVdFDw+n7biz+dZsM2SzDCBZfeRekyuXJaqi7p6
/xNjuGPecHPrq1Exs0q3VopwRF2v8tcRjfN35BN6xvbgkXds3L7++Oi34Lt2HF0Y
l1gOHevNdgrbetUCdL8jDIab5q+d84ODztAX+q4fGj/b1HFxKY+f6AMAHeKtmH5u
HBNeaYw1V2/oL41PZfjcE/8S4alktXOufGIPi2VBpg9J/Yst4vvwZiDNWZvsPOir
YHmvP/1Sa2alnXB2nIYeVRKq76YW6IsWVy6D3yKGr1TJMe1zlkX7MqeyH/KLH3i6
8yYQ8aLSCnxhK9nmVSfJOBi5cL/MKJUxiGT5FLyQEORcR+asDiDQXYKjLZJMjc77
VpdckOeiHdq1Uwm6noAh7LHpPWqeYWDCa4Hb5cJ3JMgLdWbOZ7qxDgjHXtquTdfk
lcxGjuQbrZAoWs2MYi+83Wk50j2busP0UCGO+ox7XjaYxA2aRr6t2FdXFKMDR/TH
JUWgA8CmgPD0MHipVfdTS1xdEtuAY4oTtLF4Lin2MFAwNFPxIkHzNlxXGX1UDrnj
MASH7Lgxis3SPZ740HMiOQniGPi9uH0TEOPf9En1lK/5xGK6YHuifhSEPHZDIYAd
LROMRJduE5u514L8s8L8GTbHR9fI+R96d55TIzb0QfdM1aVGwZhniK+AGIE232wj
fpGrraHa1NtVPP75MhLiBrVwnGmki+WaJzcMx9qDO3tqyl/J9RI94s5rTm25ZudM
6iVoFTEA/tBo7HNPnPvbqpFJ7vYxxox1GSHnpUNvmW6TD/piTmyakx5Np7+rJSK3
KabaegfU4qrNqxOJ+PxQpzP2V4bHw/xCU1kbAf61jr99L6pBO0MBl+s7RGteICes
h5ZbuSauLzpE0ZmR2GNJoMbIS1qxSid3lmu2c72WR1+sxp2NlFacN53j2p5/f6Mx
JP3xFUd8pUjyPfRjJSCxaKSFqEiIi2IwwvtRoI4ha8yJyjqpm6EPaPciV1SJzm9x
EtMvVWiu7Yx23t46NtQnCOdicPuY+jvRf7GpnsFsuofCcMElzBzXLuwUENH+C5qC
+TbtFTH9VJHTSyxTqYALjbOioxi+IYJr1guw2iwje7510PlbsInM8UaHQ39g4PwG
8TRvs07Ly24gOBdYvd8XNPTAaRjAkP5f8jdX7y5PTNRfpxzH9DRYqADILBoc6Ibb
VNx8u0MOV9G/0FKcsvYgJMkKeqSZYM+r5WWApb0ohaKf+73XPrv52imxAbHB632N
I4mUquWBtw87dL2mz/GuAwXza5QcSIfCI+hIYjuY2oBfMs/nr7FdVldqDqGPret1
RE+oZrERftP0efGkUmoz5PwhFBuSKW3ZcSILGHMQNNuH/3xjofMaHsKr9/IerQiz
Ji+RC3LOJMa+YKtxNzQL6XGX+8U8XgI4lVB6xnLEE4f0MaL6t8qXiumXrVMtHVUl
DCMeTAe2eYV3DpuNpIt0RjmDvAWGIF1BF/stN4hsHTwGHKb6R8OmFrB9wziS3Guj
mMmoq20Pd73/SSZSbL4NyQGHm92Enddhxble3K/Ke0JV6HTK+z8oBiU8u4WY6AHu
pqUFS8YMIPto5Sm643hJjxulYrEvJ3cCSd+PmH3/lvPsc3UZwT46BhgzndEAuUm7
ol/UTQPwCk92XFXgQbd6I3IpZ6CpDsJ7aR2dv5irBHTDPRvISkR97xmXh3M0M87R
PKljtF809B28pqxXy37YMYJuGWQQ8PCSZWP23o8O+ubxTFo+Azgk6YsqcXRqKaHR
DIiSVMZYjU5fkzejSRnKnYBe2XRvMZmmyRVj/WSEk8ZyhmvRsIt40JfgsS698+7a
2C31+tPOvXrAIx2yO7h0RMjuU+FCtwZxW2INOM4dgO4/mDbN3OQOtlHHs0bSutFK
7kBvslfr1ZOWD1kbi6iqY+N8miZ4DkEgbWAEvX1YIemH8vq8F2oArghNfASBAV+5
ZgYWP06ycbjFtzzu1psNQYqrjI9pMDw0TjKnbtaw/jqqPwU0VETQpBxYd6YorHvk
5Y5vgVfYkJlv2nPeMEk9747dSX52Vc/87X/uNdXPOg9ViFgA+rEFMzfEN4MMjNON
qtteoZDaMELbimFDjwfSfvZS6aBvxU/Be0RiW+O9xwA2iJqIagkIAg54kKJJ9Ymw
nn7GJVJtloEWyKG0EhHegFjfjZpihWRPi775wcipYsNOD5inyEje/BOGUK+QfJ8x
PxbVSArqREA/9f7j4vXCkYfhtwa/rWumf6BxDsIgQZVGSLAVBE3hWL9vq3lCazYw
a4oXqpsDTPPrgW5rawuqL/I82Og+NK4Z39phgOCx2F1nbURDJvuk7v2KRzfoKYJ7
6P+wr/nQKi3Qewuh2NQYzGxhEkJzM9N5aiGcUIe7o4NGTNmH0MS9dzYr/1HNTHTZ
G3aolmjMO6OEn34IM18+d38SR1xxq4ycjAYV0XFCoH20cwlfwlf1ojzt8wvTOzPK
+lan0uPUc+e4wFdc/hohuRQmAs8mzvtdSppCIW/+JsXMHPqo7GNJZI3unATXckBI
iUWgqNs8lXnDT5xDeI3PgZx5HaEiNVvTns2WPqZ1/hW4F1A0R2aqOmmt9EeZ7BWO
ZImTL5z3taxdzfbw5TSzJzg9FWaOCdS2qM7VubU6DNYOpTA3XVeI78sObXuw2xCD
IAmPckjfaWl89s2WonsZ6kCDyBqzKVU6c9wJKtxqda4eTqEycXOtqzhxN6TzQaC2
MaAjSMthvu2Bm3B7JXg3zxRICn77H619x5hRZdgm7XagEgZdp8z1+EDy7VYembaL
mTmWW+Aa2+H4O7hZuTEOYxzVp5/u5sued0svja5Pvq+uadE+3WAe9d4gmIACtliT
dfEsGVS6RyJDlSe+3gHbWrM0bR0KrBnX/E4STzpVTiOlTQMbymwHJ/kSzQzrFoa3
t7FhQ9B9oTS0/qJR7ES+JOoALH3smIscTCXcRS//zkIgzPmHXnJYLdiDbNyzQAG4
g703LOtlh6INI9tUk6+IELRPW7wYCeO+x0aaZcjFyh+TubUP0mGH/hyf2loi1K/B
VELYhyQZ1S4gpgT/xvO7O2diQyrLOIkT5sFfi2zyUDzLP/70f5ZE+rd5gr63rkYR
tuWe+QfEOQCkKTuEEDR/+e07AN7ZlWwewgX3vKxoX7czYtIBohnU12nfQMj4CVTG
tJPcOAXnLrXMwzpiO0NwWurCayYmkm1WrzSLy6xQvA5GGlg8iov4gjrxpCtZCFpj
qSxK06A5UFtDrKd+uI5PpSHcsnX2F+CgwS1M3k+KiMpTZN9EZYyyRqRLd9eHM7qp
akdvMcoS3zei6dUXs+/Do1QMea6Cv+MEzIthA2nrR8qT/nEEn1icskcx49EL2FtL
lk1H2iQIaHNK60TW0VsgyNy6n8gD4gJOf1HI9sbgw4gOD3SYew3qtIMhU8P7vIzc
9xZlL8ovMpclz4QapoNdTNG3Xrfk9VdWa6puEgx+OvCD0sHU9WI1NZJ9YuWrD4wz
8BGE76zRPyyR8GGAhr6gSEMQvYt8T8ERNtLZmPrzTtO080z4PsISvZpTIdW6E1dp
I5pNgxXUC1l4gC8gjOtELAyh6ls1l+aD5Qtz5qGFMxy2UXyK/eS35tr/DhJzUiS7
R7S0ZH2tK3lKS709k3y2wyjOERhUrXqObfmU68be22ALyDfqjj0Yze62NNzArkSY
+6aRqltGd3fyDUCbyArO61hvRg0DhuaFtfe2AuKiWWDhgFOT0BEaO6ei2I0fxgjL
IqEcEvWx2i6NkCdLvU9S0+9Z13GU0WqzJG8K27XxV1muRvAUPgpQAmOaV8l21WAy
iMsm6PrwFdi5QLfHx3EVWDprbY/iBQP3vRBP12+yaxfLBk7qt9NBW/QlS4ikBBqz
Bp05v/L28nUzG8qc7hfj257DkcoFhbDiW8XmBCC14YzminudzN7avYURMl8KZmqB
wSEVgpxmdEXJzqxY+CEfCutwDL+WAFveI0/zIqNy9Tn0C0Iep2pwdSHUc5zFx89D
mzxjm90Jfs7LB+9GsKRbYHFB0tQxwiURXt1zeqQGgtMoKGVf/8m86utbnKKfg+Dy
CVEVhjJhTAng2Y1n2lTZZ6PVlpwEa0A0ZUiNtJVxqk0Dc3iVhaYSRveHCdFOFRGV
yVPr5yRLyeHkxXaClzLyls9ZXSuHLOjCUee/Dq8IcfhX5x4d+h91u7GkX4G+/KhA
twSNaB9WRKyGOb+telNUuSyRi/h/ZRIpcmHifAmCLGii1Yr4hlf+E04SKZcyvDst
lIfFqZ5QZHPT9VbC06uGLvdeX+9xP/AGf729iYj/4m+ZQnKwkFx5OT+jgN/fvAk2
2RqJzWNa7P0EDQ/S2Hvkuzv1D3U+06YqXweX9SE4VZExV0Zg5J8VwJC3jd6laAwu
Yd5THMNcPUDIGaeDMVhCa7PW+MTJLXQvc4l6iGAxcJf5MBUbcCAcBrqyeqNf2A/3
ZEA3mGam3nT0BXSJTwgtxpo7v7Eb2riNmToQWKpBXbPYb56uVcqMqBFLtSMeVg2J
MeiiXoOWcKN1EZxxf4ThtxTlAcAtCIhyIFIFm+dITYJI8Tm5zqgjXTK/ZR7/9Wub
uEDu556L0Dw+lY/RTXBd1BsQqkI+VuJFF2N1nW2lfra+RJ9gtYaFEG9XwgMdj+Kw
JD5UoT8MNyVtATBuYOuQF00Iwk8P94WYx4kDStdjGo/yB+48VxFrsy5qK0c6QYh0
kLQSSsm2LuVYdb7wn1e3ggS4QMzb7pbSXmlSB5NqE8UMXP8WGyqRnGN4vjgK7a4G
Iufo/+EE5Ba2X+xaRx+7e/O/VdsK969CuCBwUkkFWbtI825r3KJanhpHNgXTpBB4
IuIP9PHjWVgw+f3yKwV0qsB6ukyoQS6gcaksmneNFIOEmjSNMXLp/yTcAEbPK5NG
kaosXIoeSFbstWGrLQV8V6+ZJIx2dlWKYjMHJ9Kp+LTdS5QLZbbx6nuyEJjnaYZO
RP9FzOYzsD58lIV0lDfuOkVzsMSdLLumLE8oUC3QT6WL7TFYz/f3OLsq9GapLcai
df8obQKXHBeJU7rWfHGV639W8cdcF9h40jZpCZm1nrz/O67cTqiKbcDXv8lJGFKH
1zH6W1xfGcSxdVs5QWY8MxCJnXjViwL7/7Z/Cyda3o5Y1PnkcnThmlQTaeTiGEbr
L2nH/jEzIrsopt9PMb4gmZ1KHMBK40ytwatSXPt1C4ugvS4vhUwh7SkNsayC+GmC
KLGIx2KxaTS94XTAs0rXZwiuZiDXuLBwun/aIqU0B6L5Ws7UO7unVwRzI8bXAMSO
33xXwu6oZ9bJ4PcilRZp73YkwW0GcFj+v010oAr9UcleRINUefn2DazajXtvQ88u
tA/ecUHqPSm84iELbbK4Zq2wid90rpOO9Kal2dFUfhaUwDa0DsQ/BjGsqB7OJ+cg
2jV4dDXLWRSS5rRNFwc4OchpAogBTor9C+w09lYsBCt1GRvpQ/kS+APBmxhvQaSO
Ddqa5H92rStUT1g+QAZcaAVAirZzoAwH1eFFOtLCePz4M+4Tq9J5FdHyMcHa5Ofc
bA5ewAhpqGyB5smAz6ijotXfJv7WkpA1UkDVUObb9uCO5c+BdyF/OkqIo/VWeRHM
2yug8oZEkIwWbnNJs/vaH92I8xSg29BPHXfIWNZmFQtFFaqH29sMCbvAn1eNPmzV
MDyDHXxxeALHUEnqGtT8vwCRb+uKgtAnTMCBuS6gMBErdarLOJKJZ+688TeTpJoU
Q0rbp0+7XvGgDEBmfaKzloWN5WLSJU9DIdyWCwlb707Irie7UzGWU1AlPv+HZMGi
0JWmfGbYclzQmCPMzOGyvugIO1BcYj6jqXq9hR4hfSjvcnaryFvSZpz42JH4+bDP
GDoLMKOQ4vrLlTZ6MnGHEJD7wwrr9dhDPoRnTYlGXSqbGfgXAn2iIXxzbPnrMQnC
VpmY7QuAlsWq4um253yohAmOLYg8KRcHtRlWcgjqNHzte2eUNAT55my7z4wFcRyQ
jyPVq7EMBbrxgWx4hKHZZhV+jiv8MB9FobBSKl+X2QgxyY5nfQC1gSiw9nNHsbla
8bmGYA+8c2BAPwnjUvji7InlRVu3GfYDBNpvTS1994T20GE2LG9dPq39cBDB9XVV
EXZGCzr/uRQ1il/GTpDaHgKg+dOOB1XtosEqXdt2KzM03OU82SDgJftWREX+KSKq
urf/Kl8uSN7YqoO2YVNH8B30+qfmajoflYeeeLOfVhiKc8VB3yI+s6K6omm0x5wz
5OQ3cmOUVA601/QfrdBuvJMNUEdMWjWsuQ0JQwD69+XYP41Y+/IrLA8IaQyL16DH
MtnPOHYLWYM8YtKUMBy5nzLEYDFXZ827N5Iv2utbVFmTJ5/8IpgyopAs3gsti/26
A7VRkeJPQJfBP6k+SMUNiG8fs4X8h9uITuIgjjksPu7LsSYdSvkXtG02EWvXYiCj
wzIdvebxukmpKhtUOjIrm3ALY9/eDLUG4XEfARD3wxASS3eypvsHqOnQ7XtmtVhD
8VR5XD8LBnec7iqR7dj2MrM6O9wGWNXQDqhGrzK0kw8ZYPbpP7OZ7SAIItd2P/LJ
j6LCNuyAs6cJmHwGR1tEtBdQW+L8xUzxKthmFo8RDLtNcna9dfZgrI9mmojV8zkm
Ywolra+vWRaeKBy+TyxUi+SSc1LaVrVEXBPrOLExNM6x9uEs+ucGZbkA48uz0gn2
8lmPZjn1qk65aP7q1w01ZFC4E0kAE2Dk/Z4frYp4oB59PaPcCjXsNZu+nkM/ioAz
elmorb0AI4bqRvQftEpS00kZ/mo144Ml/XWgSTJnR9YCemdXRgfm+tu0tFHOL61M
0aLJr2gyVqcgzPI9mTrMeZls4ZPFMwR5gA/gCgZse8abSKkX4oqvH+cojBA6rOTo
heFh4yamlpjtA8a2OGEc7NA6iplOIZAD+U7YRSwmsL6D44b24KTcnhVRhuidH2jC
T+3I7YL/Ed8B3tfB19m6cRMQAQnH74pYUfYp6H6zJVN41qCkOlp8uuwNNHfeMKdX
pIb3QnuXwTdtgpsYHJmwokO5eBvYDlNixeiFXCpm6yU1uPFlrhg7xASrxB9Qano0
6YuA1fr5Q7Aw24AoIfTHBjKs68ZHxcCMgfWlSGJ4w9t+6NAY8CWdnIEfznC4ZiP6
bkZLc02zR5kNGUrNXmFA6ijcQyx7JL+9TPwCbDIHVtwVzsYFeHQG8IdZeidMIakS
yd6bqLnxgJxHLTeKjVQSeyblXcOJd4mFtH8MInxzhkdA4iu5lfXvR62PSS0WrwCq
3LLlzXC01+CBlsvqk1Kj8/2wOdPh9oY0tly3LuwxErxa1HYAiVbY0HQu3nGGnhke
tCJ/qvs8ELRQA97zb7qyI+OTtWrq1XucH1N7sZVIQB8Jgj/w4SyMQku3ksqMxcaW
Ok0nt5QhOChbS8DlP/3/tRnMQuLksKCLzXJpgeiReYsNCJgSE7J6AJy5CT/iUFoe
A00WbAXnPTV1btr1sB1v38RaoMM8rfo+VQX03t7C7Ad/2Brj5zbkW/g6Zt9eusxe
UTxjwXLMnOFnNrfRGXtD5yaiHlEm0Sx1R5/T1gH3klSstyrMimvgLiYIZTrz9iUH
xFSjdzJ1D0XZQBHBrpwYZb/bGe1k4WDWPYVpcvGuks8B8xMBi508y7YU5tFWhJHG
n+Fid6yzEklEjOltcN2DHx4EL/wm+ZHdwROUX4MVL0Hd75fEEfSrJrzcwwEs/rxS
JgYbubk2VFW2OSyg674pn7vI8i4TOMOt4uC/3V5zFrQwGXoIGYYPRllvCUZwtKpc
YqOydoZ1PMFYZxf6c+t4jVWOKnYMRWYN2uz6IvmYoSC72tWVDHeYikcYL8v/JkJS
x0/wD3j26q9dj8mWg62NkdYnuOqb0WgJDrEg3jpEarGvpNGILUrbaqRwjFDzxeoT
IdRL5uN7mOFfhkOmO8/TZySQ0tNWunbzb0vMK6fqZscrHIVTE4Z720h7xVRaMXG3
CRo/N3mhEOFNDKRsG7c9l85+ncbq//4Asl2hhUFhzB5yKhu1YxrT8lSALxzUTsj5
pMaw76PJq+sPbCHST+HlbUtqiSxad75WnuofhwfL7OTGtaEChQ/x1vGnlCI6t4Tt
MPfbi64qorUYTTUStE0vlVYtNuAExUJ0jVbISY/In0AQv+97MaCa6QLTBGONqVmM
OaCYzIyy2ZSRU1afn9egIeJcvOv4BlNrqK+DWMLkg4MSebOgqlvuIrKelw+XWmW1
dWH5TjoKkJDP8AmonP01Lni+wOq4kA1k6iKWGi/+dPahewpj1gho890P2f5/CttI
oSX+w+DgJS/yb4uuQE4mIydXz3YejxneDCSUljuuHNkS6e1Tlyp2NVPTZ3LwpezG
lduP3tc35fvSMFNKDFzBUT2N0viHgt2PCdlle/c9lQkoqgV16btddZW2+BHmWZdP
Eo2oLUBspQmQR1xwVGpiAEoOe4JYmeIbHfGK+FwVN1SOndv6BH/if60k+6y/NzNI
OHhuKHcDxlu+uDZF+M5LRmy6A1vIIr36271pF3DParEa489n31oUlsCwwTY86w9y
YxOP+qwTblD+C3SM9Tc+xUAJkThanOV+hPdiEolmqXJ3fZ7s12clej6129YhijWn
AEdqStNrciz6xU+CivPUvXKx5b6+wTMYy1mLVk2a1RJqMKkqRLI0SO+wU+8aKIny
Pkz5EcF1PoXbYa/K58WrYSs7UgEb3iwBJcREJQAI2njkC2zWutZKPSbPtQ+REyar
MERmffjz1VkEXZIxjHs7rvtgHklUOm5lz0eBWJvIsapAL16iGtNKdJcWG/OitEQO
gwXSljQkWKvTr1zso4yMaGkSA9lAbqYVwonvp1zKX5IzGz+X4aIBfecXHzrRUryj
ADX8N+LFHUCE17lwQ1aem0wuHHjrq/vD2b18gK/dNcvIc9aVSVJKw+WQEgHGOfGI
eh77WzRzngIzu3+icooe5ZWmH6Af86l9DsKJo599bC8xKDpk3RC7R513Hlatqav/
xZk5Wlm6WJgTvEL93MSvX1EB7BpjHtukkqPZNrf6g8GRdscwRc9qEfoOGrSy545s
Luj+RCVEPa9DejsFtzzPEsVlPBprIS9SwZcE69VyJimnDqWrw8CPtt0Tccr+uQ6Z
ddjgC3bmPxdOZabc5NXnn1NythnUIWmafd3e28DlK2WmanGQ4Sy8KjmSmbHNytEM
B7dMOLrG0KP+Qmwp9TSsqxyfOX97CnzbeSTVzuwyMcqwvrGUQvibKQ1FEHwujFs7
6tbbGtvLPhnvjxO1Tz4MCdkjXXJRDOSupwc+vHA+EtH440rubxkXm0ZNy1jjeiRE
HDxxW8MNAjAX4+jLCI0mmTIMv8YAR1Ff+qxALfXE3VoIh7QnTUyYhgqyfcFRrYmm
l+KP19hx1KkLTVmVb+abqS6B5DHy1ZLNkbqSfFNlc3AFm9gNc8mMe+We0ZNm1KWN
5hyUjumFKnqAEGIPNCAeKxn0Li1Azel1JClj1S37iNE9L6o5bBGBOECAGzQlhBLZ
1DqGIWJlJa+PQGTlABs92o1U5kDehqkKGu0kizumoALCND6HkFCfovVjBf9bhx7p
42nS/ldXKrOlw2chNmQfjzbWYdGZJ0iURjk/RW9rkgODwYNrGy3RstGUDK6ayBA/
X/rEfZzorlwvHVozP+ydrgWQ749TtiH0GmY7AJYpJGjbzdDh9TqXdX2oMW1EtvDk
YHQVnlVyP2VaMYfLbx7jz5kMefmnfaZ2qLSxuUtDXXDEeQumbyVtSseb8PycL3cP
qFnhlFinxQIdQpsy3TrQedU6Xy84pY+PPA2UjKd7uvGJ/oVTENpCqDHl6blo7pT+
s7bwSXSHdR7Wwk//tQwl+yGS/THBWjJeHPfpFvPYq1Mx3L7BUsuV0hSi8ZNmiSJh
ErUsV/zRBobmRRr1rS4jB4k5UKUBS6pchNnvKSPv8IadH9tAw+xwNYtJUtA/Dq0x
nClbQH2VItW40gzWSuue1oLBMiQvMegEhdtBrM1I5XsNUV2Y6DYkr17O4Dp36B8C
tOG1pk1mFpr15UGrZy6GSxs8vEMHTfosydLQH6krSDizhXgsn0dSJHPrhQxxtQu/
mU3l6q5V2Qi0bzHVgGOgD8UfyjfvX9vL9w+bb2XEIgSsWy+ryV1jKxkmzp0hnjzQ
mKM8UHgDGFIn7k9lrna2fIT9hW/sNkS2MnlUbuMBTT54gdPRnJsI68PXzvghYvGD
QaR8rxV+SK1vsGP/3m0vC22tuHCgKmFhgtJPflNiD4DY8neBl122t3gElSul0qnw
xlKlHMy6NARNz3U9NXEjDMW9Ns8JZYJXuVhQ8E9GWmxj9C7tsqFHFMviKkCfnVBy
kgvzNEcuQ6r3E5TO5XDI24l+xaLpASwbQ4b5kAXlhyEExqGb4SP7yafiUi5Rgon4
+09WeQTpwvH0cUzmnU9EMp9N69HmcFPzP7b6pEB0j3bTBLdQxMTGqLG5/JXaQwFR
9dlWty+6HMSwFfkg9CspJj0aG1GuHqNdTjCyMLA/pbeQDrP+Z2sqDs200lrS38Fd
nrJAPOwGcbe5JFGYlCXOMjahhUyhpdQ+2/yiDzValNLCWK8YlJf7W37H3XT3anlw
VGcIBZyoYKEYUsQ9Ry9gGz/Vahr9dGUgSKy8XtOwpISwtYn3jFDTJ87MNhIcGTmn
N6vrPqpOG/wGJ4nwMjvHEpfBn8MJyRJaX30b20H9tdqSGHcTTWyfEodHaRkpG3tC
extYumSTRnS2OIA2uT3mfe/IwLs59u06RzQ/mKXzRwGNIKWDd1H8G9QI0vWugo9j
lwHdX/xcDbPkyOwxaHCiid8Cu3OdQCMpP74rZ890XbNkNz8GI6NvrjRiPpVZfIlG
YD+UynwbUywTKNoVkAxhU6SyiVSk/s1cr0kYu6GFjCIkYW0bh24rECLqYl8255+3
qwtdbsR7vB4CcGP9Y8nvLevQCBBqu2c8++pJGziyskYh2x3uziftTI5B+BcD0KLd
NdBWe4Jt1gMjCPEcGlKgEQws7dSy8+YLjeeXqWKtVOyOCGGJTvV8O0+ykOolgzGp
zgiGhfnKm5Z4NKoDxQ4p3bZ/eH5Shcrc5IC2lV5N7aleOaHSfice7w3fEDGqVbew
Q6M5FFOdFHLnrLDd0Hlyk1SuGFh5Rt1mAyAUkl2OoF9VZ9v9soqK/wM/EnEZ+AXO
7AOP1NzWUq1ePuvSr4fiRkHvdhgjMOJgwOFsFYx9BzdrkM1NmTcyzAWkkCSp1KEB
6oG0GVdhNsJAhhNZJ5jdKiXLZOVXx0SHw7viumufD7LtjVe236nr27SozzTTbMex
bA8h0cc/iUOvevlAkqTmMAl7n8MjKdHmlOQmJDbNYX3Qw/UMXIy3n+bVUODJUWkf
NJGISrKHGJmIB1W6pxeiYOdcgPczQq3FI0kSxNtWoeCpaKVObWYFGnTDDoMXEYHw
wXIx8H+Sq/Wibu+T9p0VWvN2QPiKxSg6xLW4Bs9EOFstWp2+LfG5dMikUmx/qkwx
RW567Jb2Gok9NFgc0n3KU7AzH7Onl+WYnBw7BEPacjgKErjSI1EiEpOIOZzZnw24
R/zOYyN3pMmjhrl2Ff+os2agdfgCKNGg53csdz68e7hGpo2XyBiDDdl0d0DusPfa
N+tlTPx7GWT4km3yi0j+Rz9Hkx0XUB40AWENUvR88NaZh+PvaXQv8JKlLfyMdWzj
mi1eGaQ6K8GR1Oy4Ct1nWEw7cnLEpPXsz89lsqzKHrYbGEqC7ATCDXJOoAvBxG7m
zC9zzsnX7pwjpfPRK1QEC1eCdXkLHb9KTzm9/Z6uJD4fyAkOttPjeb2hS3UVhwAM
awp5fFDqKkHSmNlVofZR15ZXbWXvCoqlyhtdLA2lrqJv6QqQYmRA3FUyqteeG2U/
lUgfa+jpKmHe/WEDILDu9WXjY47DOd3K/WZlHRKOLoeIE8UcZpvX63+BwAlJ+6Kp
4Y80AOagpXLZNGG/bGJf60qQANI8KaYsqZDSGHWREoirXMp99IrDyHHB6cX7rbMR
RtyNy90dUEmsZx+9qFjP0QKB3s9BllE/gzGiHXWng9XsVLsi7rGLg9p5HLoGB5w3
1afp3qmQhvlxXsbsHH6LdV1n2kBwAJ+HKrzXXMH5gzGcWrbaJH7A2Uu5hacuzG57
3djKfCs/EyH0JFwGgRh0z3OG9J9NwsVqlr+IO1CFP8U4gW6z7Hdr5ftQLXzgzqr6
9LStCIMMaJGXRYvQiKBbQUjha40SJnfswcAA7M45GDqedYXJuEjOAPB4+tFwtFjb
oziKnVd4YCpY9MohPvkQwb6HCLo0lv8rhmO1Ehivj1tuzmp2DYRADFtIVL3d3rEV
gCRPzGCHqVhACoTcXUkK6Alr4l4iHRBKSCXy9iZfkXwrl2VRTYXbBdMtXlpgWIoH
bBEblndSufyURaaTogyUGDr8Qt5Euk1d6siz56H8ZiwM1Wjzf4gI8vXblSgun8/s
qLbyvz0QTfbhE3tEpcDfuvpka/DYGK6Fe35Y1mP2w4KSTwHG3MdJCtbjGgeqKb+x
jxy0IFIzdnjt76D6uKpZgSKtBiKuyH9CoqCgAzaWUHGGu95esamoRzNki45xmIrb
Jsl+T84qiRmPknOEq5em6CK1KIO5k2jCBtu+nkm92r2zL7X1DIBUBOu8jf9S8JBI
1PpywfnjbmbJqCAKimyhNXUE/Oifqcjszig0L2LH8uU9o9gE33IUS8VwLma8E6XQ
0OBn1xisHj9BP6PhkQJ5IFM685apQtgoKSXEAsICZkpTYjlrcrakD2lm74cVoGla
VCFCJ1rd5UTFL1p4+3jQUNWmAqrLWkTBgI6+511fPyTQSt109/TibMXt14nTAvYm
P2P9CsMQ9f9C5s82h1ozzP7eKIEmUytBQ+pAk9SWzB8CBwlOk1eTaXZGsqg6C3FY
xlcWJ3OPhN0eiluc9chKpT1PXuZ8Yc+9PKJMOPRc3c3BJsxsWtOFYzWMGLLdEomY
qRaDSUILeHLxxdVjzl1B1DB5yjRL01kFjo2btpsSEgn0LDJ1eYRgS++zvqQmVU8W
b32Vh0hFvtZZxeqqg6Mn+egc7fK2lYWLAyR7mAoeV6pr2E08i+TDL2GVfiKI2iy8
RuUWJSKyU4ZIbnhjvTDdBtfv4ztzGgsf0jve18o+//hJiex5SYal4j8ktI1ASnCf
pAf7WEaTpa5RdUSf6TFq6o/U5iRSf4YLqlD3ts6+tMhhGiOe+4QhacTftM8qWIL+
MQO1NGtkjEvXllO14raNDkdwuW+vBF14CehKmWE0o8NF9IX858LGU0UB44cWhf+F
EJZuO5DfmAhs+hS0jHLpj4m+MflwiIfCUccKRqUeeTwlnJ3UCEM1UhnLR4oSV1/P
wHPVYCRsXKEZGoQGzXMv9URsIYJwmObpMdd+voQI9a3eVnQ+0Lkh6wBDGVJf0qo8
7TDh3dZyo+n7dL9616jQHGMFB49TMMZVgzB85rYxmisAvfUReOpx0Nl+VZPbHwtw
WQ6pf0yMj+FXRPjrp7aLZPGQP7nKhZVd7XCGs+HWefGQ8M9MRbs1FvuR+LqZ3hrO
vdRpa+6DExDn+kwzckGWiRBNHIXmGQvQNhqXcWQFsSTgynyBKTchl1wOveR/xnkU
YuvtRRFfij5kYaGAD3vjsF3d3MqiK3hDmufKHXYQ0oG4b4MgpZtghfCQlft7SM5C
9cgQV+TPGNfaiON8Wy3GieGhnaNhhiYb/EwJ0snrwQ4ia617PsH/TUUirZAKgWFc
zyNmx9FZ07YuhoQMINCVi8qlrmGLfdkRxb/rsibQywnRabR27rpkdU1JXRkV3anK
WaHkE4tFKt9KgcNWWnZ92ocEicSROGRKvgjJJ0ITm4KbOF1Quc38yuO1TDKCLsoQ
75BGcIBs3lb/lV8Xv61AtmwMTmEtG4n64yyJGjYksRezWvXnVPiAiD5pxUSxGaLJ
vbajgQDv32h84JhTM3c4MT8eQQsAs2/fjpxzUHindGZrcpTN7sIQzoLb5V/F+tyX
7HhoLx/qaHI9Z++JHMyg5JyDPJLUt2Jdc3C3xVOFeXQG5T2c6XwuT2R7GA7bFSZ6
5Nysz/q5KOnc03vXOv9qmIFXXZBndX8nBEnUmA1xDmOq6mKiCLe5j3x2GPWbrp4W
vRhksRBW5SGVLXTXGnkHYKwH0vMOwLLIwVyaWt2x2yAasAY1W53aUOHoeoM5Wygw
0pifhpl3Tw7K6G/wOr1e1stj6MWFljxJxvDYEQaukWVG5RamqhmQYaPYtlPm1Dj9
/hFsthbGjMQTkJ9bTrJpx+XxAfGhiJTcnbIhJuPHb6iqB/M7O6+ZxNTnH/IKcjM+
4y/hBdUgRag1Ebyu/+C1vo3aP9DQmm1BcG4mbNa3x3ZtSYjT7NqCgUFskTyKqg5Y
sKOm7uvU0bv1a1xXrs8Zz5+YU0n3XODax1AfTxrl2+xlSbvMSZfl8lr1IEQEuoUU
ylwVY8RcaYAQy5RjBJxLNgW/oUWIgreiX11G5Kul4gkjptaGdk5cC4yDckda96a7
tRr/0dEXVZLX5vovX7qS3B33k+JbeFMruIxDkQIkM0sHFJxLKworLwABmV50zE1q
nylZg+aa85Vr7lWTPtl3iv8fBIYA1aP1hCdIiP2SosHbEeicT1mAj8C5ClPlEg5Z
d7QCFO7AtiXCpvOkeWKX8LCSJXiPA7MhOWJ3qUGhKRZuJfA8PN/Ly9ByfsVM5P6O
sYD6ZSZ0iwYo5G8zVO4QQ8TcI+k+jPeodXNhYHktllOhnf8urqT60EdLlNgL6LTi
ML7NZIRv5x82TyFD3LWlZwJOSayMiUmXVW8/CMaVWFdezLUa6A0t6D3mD8xeO57d
69QJzv+eKvcM9QylXAyNAiuNgevMmBWDVr1bM/vDNqE3yph47aigX2mx2Vxj68Yn
N8/74CsXPOSSFubv5e4EuUgueRkqu/viLaT1Nu/wNkx1kUj3ryrdZXxQ1UYOR+Nh
L3TKbNGHPHSc5omhZE5iup9zOShTsWdyqmurSbTy/TjQRtOXtc5cfwDfYpAEiwh+
GiOja8N+k4TiIlmRn3zAAFjaKYHihUfiZg0D9+NutaP43JwsjKqZ0/RcZiTMgDL1
gSyW3tXMMbSI+AQ9SL8o4BGmEdagXEY53e/AwgUlvEyzmcX5/E+8rCfzB9jVViua
DuHlNGzSVFpuHswnvsvKbkG7xNHy4+MJq6VizWorCiNUToBAK88dNIVyaJdz/IOa
QDhu0zUPrwcWggtYB8bGc4EvUMLxTfikFPaG6Vssi30Jpnp/uNGkANujgQ3bjZZe
xbdEf4EuRKts/L3O+DDLrW7b5NFhGkPJSqt/Nnmm5BtaOi0YgLSfDSV9NSiQRX/a
CDTmHtID/DclDh3aEF18liT/JPzyiwY+8X6fwHdlonvPrPemSrzy4VAW+ki1qcC2
kJa1UoqnDlt7dzfx6XSvsGO4fe5D9+B1q2VyWxL7sy2DfOiTJighlHP1BPaFtPhR
AQSyPq0ufZfOCW3MgwsHAQYXYu5nqxW4luDAWjxOjA1IhGAdGN+jdiy2snN9E1pQ
C7pWzIAfKIpUIFh0sIX/K2kbJBuSy5KHSlYW3LgSYt2dapKVzR+Sdthhfdze4+N6
rbXuAn+WdxioIPqGNs2a7LpyqWgKTB2klJnxQ5Q/myvB3MA+rNUFpLqv6WSKgRCJ
FcybEeBO1oaZaP1L8fyyYul2inqjd9y1lQc/7QsImWi9YwgYRTpJhgUbf/XqZQHq
CYAG8/zKUJOa2nQk8XWUMDXjnbdMNBryHgxKtMHbRyc0qlfrOhYLa+qr2e1Vtdjc
+VOdnDqHe28GkDIi80fNdGMcj0zMGNVS6+gdKm45N8WkOHZCAJqFC3mIDzDUsB4M
048Z9roLHngSF5Si1qvDmSCm0PbzR/dZf0W/XldGvS8XfgARzE9vk6z4mh3HBZ7y
WhdN9k0btmlEBD4zNmR3z5HxyJ/a3w1HYTox0BFXOoeupu+MvGdVV21s2N5xGiCX
qgb0tjcxh4m2QNLgJK+GMCsqyQTTxknnA3MBvQE86ZONsdHcQCgiJqJLTe6KAkvM
OZKLGrwy6hHC/kUixqeSyLOvFqXecxXprvHTxYcA+G8jwMeVItlrLNO3o9ucdFsn
7bVa1AzfkVSzMZ/BTahvMY2amKTI/yoi3Vkzt32T6PKI3X4jRwxBb39RtaWSdB2J
StB1YlBU3MIIWIGzRmGU1/X2fzUyzHeQ9h+rTGhmejC5N9XLY8Vd/k7C+0B0yaff
KfAuO0ljdHaJHgqnkx6DOEnTqN2fIAbSLZuWyQiNqiG3eHwDNY69RFwfCZRx6ekA
bVPUz9iWYGHSkHKtxBYO/tS0P3MX1fwCw5ueC5K6sHiZ5C9dLsZ1kEq6cVz55y30
ISi95zAD4pZlssIosSgkygKMvbUK30QUqi4JSMGXDJHFnVKHH1Nn9/Ze/R2G7hdp
ttYftVLl3o5R8DmauO19hE5iI9jqTFKDaM0gVnGNSkPZOAg9tcA3vw0cy7puzm+K
jI3JyWkPw3IyTZLaqZkzJ3ba4pLbc65leWPgXdtwV8riBy6gqTUtlC3m4rWOcsLL
krIFbB5uG6lRl3afl6s4P+fF9FEkgY6YDqwnKX3nTnAmUIy8ZTF573qU+wvpH2xi
p7eV+PAx0U7QGq0QF4mlgXuLveE3OFfUHftDiNPqskajnP7L+InqfGPdfQ1AlUsf
WsB4jTayIfM7BhqR07FJWOfUf7rgrxbXcaQidceAKQMNWg0dhmsW8yKowwdznrnX
Y0JOAxuay0PupXjIteYQs/L7L/p4seNWmfn1uE5Z3pim2TzQGjJymDZuIUDHKzTr
tdQW6Yjo/+9y3Zam5plX7fBZ6GbjGeWMnNac4dpT6LW/XohRi3wqEAZaV5PtKELq
io4jmFkSDLCp2ljpIQFB/wVvFnp64EFl08TsZRJMtiHUHQEykUbg2Rd75H1JYlAO
1Q7jXypgn4eYWktp6DM//LO9O5TwZCGsurlSYhCcbpukHzG1Gf4AeAe+y4futEVs
AftS1O/JMYN3Yl+iEIBNb3MguSVvEBDbuq8kkGC0UjZVYt54WPmur7l3yF5BtC3B
9On9G8h0Z/l7vL6kSQEcddocoHZMuz66MgtSnxiR+FvvcPSy2lKuXtOGtwPA51zj
GQz6P++bmNjfRO1DWArXu5fxwXLYEcEpfAuO1QmCY8RnWhwtuxXgQeOLO1jjZhGE
YFzz22BCH1PXX8t3bMGDU1TO7skLkm9pB7arjgYTV4PtAylPlRySseSwrjF9juZl
7KJiv6xuxOQ/IdUVnMeDwNVw3ktZRQUMZB1xBfhk2hN+J5zzz5CtcmCH4R+kW9+x
ZCmoIzPxIC0M0uxa1WhedXti1EffpU8x0byy7OcVwPgmG721J1jg5hb7fV9EX8nZ
28ujO31cXTQ9+zmeF/mNVyLhi0XRwzsOxAsx4iZcqiq8l1adt1LnMjFGRLBvmlCl
fYhb1KdJZCPaE+u2llns6ov9xZfSEkbVmAp+8XA9WNgQj2EOlCQpubBqfxueJEtQ
xKOFZXVlRJ60TSNU9NQkpnQmzz6tLJvVGZEpLAS66Do/JA1pCx/GzonzGJDfj9w6
9THRbePQvb8SUAkdkA0b9D8+UZeT90tsIHHAcdgixHXlOLhI8q/HeLQ4GXypOCyl
dcB4JKiTyaTFYop1lYrT22FhlHrLeTPUx5OW5jWDGMc1L0lSAfv1W7Z3sMCBl9/b
3RvZXZN3XNQmjo2eud1WudOm8BMR+vlcX68KYCN/DvKgdbxEGQXSrTyVEDa98DhA
cmFRHElI1nWc0BfGsvq9ABOEr5PGwgBqYzUPODeCiqEPDQTtVNWYfkJixY3HBQVE
4JHh1HNzoE+7DGqGnuWKAVmA7fkpqtOr9AU+jaSFwqNNnA4k13e+HNV6Z39toUG2
gZjp8MzLj82Bo6hsJoR9IM1lSuF+Hw1I1qbfN4cwcXDRjCusyxKplpwqWTZf+GNi
jpWopwto44rvZ/mWKQoea9Hek0V5FbE5q0uk763jLPFdRFkzxrjqtKG7VwcUmtA3
rDf7ZwLEL1V9pULdOT4VwOxC6if9fw6k8bTCm+wkfKE7Xeo58NchrZ4lD7nESBt6
dHCK/z3dQQLwjYxqZk02zIP1rM9+0CKcFehAXCBEOZ8hTtC2M0oAz3YKKaQ2+U3I
hq+37R53+RxnW8avrutDiygqTEfMg7IkuAkltcClfvXCF70Dxxkg23wo1Yn8MUKD
WtAtPSUAd5q2TLS13TE7UrjzjGumyfnmOwKoRFRMbi4ecD+5p0hQaOCjn9YgKYB1
Dr7LG0tY4kGcRlItyrUItDcvvPcRcz6Gc3ZjaqM1WTPGjgUj0bCcpvBxPH0qgSN2
bzepn26gxqJsD+IKTZT5extOw1mhrAix8lorKIuUdO13x1oQ6ZWRJ7OS+DOPPeSC
tFpD5qXb+CjMj7I2QXY+6fWJvGH13j2z1o7tlQm0JouevvvtTqrDkLbhB7GFJ66y
nSVTEvgr0AfYW7fbxZCQXdqExRuqFHUdZUzrvQprOIkv08kE/IY57EospphLYJHW
zJIYgem+klCRb6KtNCv9fQWArnISG5EgzYMMnF7/TVrZINvJ2INZZqOa5xb9ePA7
+40ObO2ABBD23+5wIUiIIGzJKVeEoOcQN5QMgee+so4grk8Qk8VMPJQf1rTNwUyQ
Q/FMELCDjO5DXbbQcF6o09Pu+yz9t+XeJhxgGnJGlTU49OM0urph9QKYBbs5c644
XwrmLkYTGdo5qUnik0LcyVITLQOlhXs26rSD91MCIIWqTctvbHGRi/H+6XS4l+d5
1ckGULYpVTinA5wJ5ww1dH9C/EFKPTlp3uYf27+2v3G3bZiAvU+xgn1uzuZHfe05
p0/EY1oMF5ck0aZreWHuipzNCo/YVLXc6ryk9mWgd1wE5fjONwKlYSZalxjq5NuS
8tsZIA69ERq6oEyBuV5hHyWOtoNGeUbdkdvT3UE1g6sJswttQh9NFy8iQ2PkGPKR
rwMlbs2j2O5qunhjoIrfZ8ye44LkgZ5uGHLOhNMiDTV538++00BHIDqRonyCwC6j
OREQh88GCog2QNWicD73WdtcvF8vdhe1IIoJ5oWBT5wA+tK4yyd2fBIdXrZL9mN7
i3qWLnKyTBuU71PJ5QucKt4YNgKU6yJvRkUIb3P4JbnEQJz6cQON8G561UOk9pbQ
Ln2aeuyKRfQc6X/LGCO/j/eKsYwvgnoJPAoMwx5rWM1sNZbbcLi2pg8KRVCAMGIj
L80basviZYG0cWnutW+n/0LdXe2RFUEmUIOteRWdioBj6n30jO46GkfKJo2e4a/l
jxSH1jNX148yFCh5jOprjtWv3ujCACwupQZ7thSu7L/F66cQ2PGI1ruCF4zo2fYG
IWfyiKkyUAi6uknkMMjtaEAf1sMnCVJS+CXxVNcHPvv5qcYUdgNeqooTXBr/xbik
gyr84DRIJxN42euF483vv1vXcbb/gSueeUQyR27rQ9WFtpJm4Q7u0zCRg4ghue8K
D8pKMCYmUwL2dHT22UwC9TEeUuxJ75w01jNVXl+OWw6q4MksrHAV+5ww5p65FGtY
FkB8fs8NdJyqrysafBExSiCTiHf372ZCBTq+t1oePdRn6chMYV8s553jSV6pnwb1
bmppXBjpYyV+F8gsIvd6WZjcplfigalf1rdcblDtAhpaqFzi19keQNKxSDjNnK+U
ukRH75lIyrxKixR/D2hrnsuMp3JjQMrGvd+LN1XcVh7OcZqAjJmPPOUeowW8wiES
OWKy1QPCertIxcHhvVJHmidcCqfGjV1SGiH0zQKMMfZB1rs2fV4jWQLR0bDwSPrk
2iytpLUNr4pYu1xA1w+dHQ4ahOwH0Ty936KWhS60DkUW9t7UqzMogaH1QlXI+7zo
6eeyULhaFBb4R8n4H6/BJtqoXEUnCk3q3c1xMUP1qkH0lW1hD91LgpNZsLQXMQoF
JiI+FFEdmNJtm6YXA8t8kyYbNqJMzn5qytXaPS1v/R9MzLjo1YsUzhVGH10T7DkA
5o+IxgrzkiItOw30sz0ioT7sJa77aBKWCY9K7UQbwDPOoYnjInqiNFAJsMNlF5cm
YJrJJblkEDOt6TkzteLhJUVk1xqqD+dQo5BRKyEDPu/Nb/5Su2npxKEAHJfnivGI
qwM979BRmyeQHBNwJSBE4kPgUuM3vzQ+1+R8+t2oqOh1cARj6QnpoQpW8vo5FTsZ
iV9CgOdPdSGvoIhQ/rmPYNOa4oVzMV2/J58JEWSqNMuxgA9NCVUmev7Ugv83k4zz
ewbo00sQdsRPHPXSZaKe921VSccgaGxgPdSj4Q20ZnLUEk3yuKOKw7Kes9HC8pVt
BSCvptbi8xBMKoahXj8m083x9rIQ6NrX4B3Bw+cf/v5l7w3shmtd3mpZ3CYOpP1x
KJgPyTwxbwTT6LImIT4rI5iiqy6IZwGC0Qm7kT4AdDf32h/XO01z+h99obtEhmjx
Yui88xb2rWdH9pI/5CZfL7waa/hEC4732S+ZtkmrXRDXFD+b19KAj6PKgNnQNQFF
OxrDB5PwE7sAViRJ1HyGJ/P6tByEUBDICVHvzSrWNeykMCkvGw8vPaFA2CLb90j6
ieZSGiRADu41y2mVPPoijET1D9W1AUWpcE9m4ELMAfj75faEvQzH0E81tPCMu1cb
mIsuykPHsED8MgSNV5iGCOmY+HUmk2PDl8FzP8dNnWq7IkmdQBcMbEVLgdIRRlTZ
J0yY9FGK5DZ/Kgn7nvtnr/Dvl3xGbJLQIP0sPfnKTFgVbhBg2UNiMYXIlJdMKvFa
/UNxVfgU+kR62oplGCY3iO6Uag1wgU8c75DVTE4eXMnJaRtcNjLc9Wcyi6ucrgGz
iOwcU1nGuFJAGyx9H/itfckxrqJdO5FElSzjquRYtzNeuqMeQKcuiFunft5u5W7y
GZB80boCHkpAYoesaeYFBx1j7iCXLPf+FVij4qQ3Hg5e4LRdDiocXwIBSIsPiaZn
4RD5kwJQbvHbWEmtlKmgxqlkwErqpjHzv4hgEo/13RweVR9EQ2CED+sJSvqplHQT
skmYC2nWIYFDuHOUx4gtei5FVDrpfitO7eo4qyzhSGjjciE6X/LDZ8bB0LzY9xTv
w3JKYkMh8UOA4Nd0/EhXUYVqyuZVUPdd7joPmcIHBpuEU36Cw3iiRl5x59wjiEl0
4MNolqpltMyTsBrDIBgnVhoRr74gl4D+5zuaKABLjoRpv0ajS9VrrIqgxvW+bHIe
JtIyJ4LbUKDDrlf0rN/LsT/df55C2rsoK1PRfjPI5uGBA9I6UOYCph9PurhDcawJ
j8Qh2uw0ykJzTCZa1fCrGfkf7azhMWCTHGjCQ/pcmeNqi8NIMXHyGHwga6MwKgMR
P5eknNiQrRfcw3Vn93MFPIvLKvluUD78/QzMzNo1/cCAd2bp6wrkPoHeYL+gdZEG
LpsiDiUYBwgJEFShVRr6C0+VTS632x+0HVxdiEHqbXlkg8nHTOLpKCUY8QyyP8Jp
t+faF50ePIT5IQBltdUMcpFEDuIoIUj3UO4SgS54k/mIv/uVJP1D8n5uWmYINl6a
eDnd3lrT9hxBuNF0RbVzzjxPQGQA0kql/riFdcne0zaG7qPGuKZoypEp9uEyWGob
vwXP1ciP45pTE88tkbuUnGz6zxLFyrEhX+zj6mwxULYqXsSGZfDntCCg4xfiq1uk
s1QCqSKOdmjDLUSGsGnT49ahXvecpYOpbSWsUiBfxYB711MY/XoXSAfXGJySyXpK
O3uxOucTN30t8m4sAoYtt+QAzConKY3eWH7k9Lzk7kyAwc0EU3sqr3ktLvzn3mH1
NPFwrC1GvOiu2PNlZcs87qKDL0avpQPWjY/fBf6YptAeZu2uMiLQjfEccB3NKZxC
wa7Qvi8GHycfRTLCCckMKscxv1TO3xKlCHpSKkQtjG/vSiU/Lpmwsns2r8UNIOno
R6k1jNMYITQSL1qa8WMiHw4lYuKsQVJveqpYAn7GuEs/9nPiwYJQsz0W2OOKTeAh
7U06m0WgHTIYI4W3pjON2DYWssHIkXNmjgIsuIng0CcBaSS8stVEF4HIyAyIsnvl
nUeeklSwHweCocV4eISovP5SPAZpHZA2pUkLdjbnBhGNdU4b6Hc2fxCI57iSauW4
OpXcQsRJukNzXDrQWNK8XxFzd1nTrnn1efd5VqWRONcAEiJW8r5nFNHvRzVNEaXp
xbHRBxMLJYZbc5wgh5yXnVbS4EnkYFhvB1MLqg2/F+x29WzioWNYLo9SSh2MNPC5
xI44oY/Tkko8JGUchbz7rbqTHwIyqa2hffG/qAYGN3RI5/pPDrkQYTNmIu0qKRnv
w6cYb5BSMlPDhV+13hLjncbynV/yNQ8zl75z8Ax905gruQalv92EQc+O2kRcHZ/r
yOiwq4TJs6WYM6BWscQKT54xc4I4tUBMZeHSeu2WknxXur7lPCcUy0wcQ0Efze26
EuLsm95QjI23IXjS8UXHcyKK4bB7lXwLhP6sgFmyB76qqPUI6NHMSEiDKzlm5MYr
AF+zx9NLzNnM+9BNc29joWtPV3vK1VuEN+FS2HLUf66JJ77RFVlU1KOgeOHDsuwE
R6y0qAlHTz7YAHZkweOcLRIEEl58+clujE97DpJ8qbOGo4kInL0ayKJjSRNYVem6
hyV8byq4ThPl/uLjLmMA6ETUO7V8H/jyzkNUbIjGFYgWbbkmY56N31S9wO7Pfdv1
jtV30SDGVSuNpAFevEjxKb/cyL70Bp2Rer8EJOZW/8AQ+fbXKHcbk8ZN8qMh5mpM
Lbi2ploi8YukJ2nFQBizKjPJwt38+r7znFoHUcL5C4oXJA2egcgEJhhEh6EHHSOi
W/Vxk1orIkWEwzzWNSdot7Yz/lCTzmkKyRhmdi58guGrgrRn3KZI2wwi+38Y4Qbv
JUhgfcEqCCeA2wPXzj16FBQ3A+GkocWJyvB1bi9dmIUwBwljEyUenOi2Im2+vNit
sVqYdYwojRiEouUJH/C5SKowT8G1Nz8FFFgAIx3BR+X4Isdho2lnur0vOPnZO7w/
pWFNZ7Sp5yi0dTwHGxVgtvuNLM1bXv3eex4huWCN6mjr9DvF/v8xejvMGv7EPWrX
8xb17JU5mUyCX6Mt6+53NZNwRrZIRA+rZrpko8l6gqak6uo1tqI+btycYI1LQ2GS
BRDz/NnlElEnn/wUMfN5X96PDE94iM3g1sbAkFDzIPLczqh1KJ/nydEfaWWqKyEK
62yyALWtLzlvnWc6xoiTZ/baNSnrwvNMyT2DJenmaKKzFm8MuPFuDNcdxWSSNI8B
GNDG484EGwqMP0dsVDMIWCPGLXKq9A5TMuTw9R942dRdDK/swAm9RzO9AwNJ+GvE
rePWupzROLzKJiPnbt97No9d/tiRT1tP3G73yvVkQCWyZWCE0mZU18fcrcbcQHEX
c14pItYN2Lcd5eVQ2rYmQs6LY9wbI1J0px11Q32Mr1Ijri56jMq4oxhbAdVqvCN4
PlwlKiSqDY1fJ9GQw8sWf5e3c+xwyZtJuakxuZroolOAnNQG1lNEzhI5uRGCPXtg
H8UcvEJXRrdNlansTIr+ZLZMg/FiHHDuEzy6etdGVkOQnIUqevsJr0QOZm1z2SsI
ujJQyUxa8HZ9eZ65MTdcp+X5HXTtJ0cE1dsRxEA3FJ28llDqvSK251HI9XKES+E8
ru6luKclCOeV4kIuQRE2ziJEfHMgSLQNCkvZRSSOA4sL01Fz1lSja8jxeVP32Zx3
V5h9jRJzD8AYXZP55HmPYcskip7fjYm0aY98O7FahwOV3800Zut8iYEMQWGfd9Pw
e/aZnmAbKB0HBAPEBQO1OwX6AywlVb/DoPTBGfIlj68ol5lHp44RW7+JvtmmFK9K
ao6fTudM8qQ6PZQhCvGYUHnGb/7jkPw9v5U6siqf9h8EnyMqSXWUxlStfzcIOKVd
dSyMqM2GeNGU/JHTGuCaPOV+1HFxBuP+nvhD2gnp6vUaiAa5tqRpXGeH4wtu+QP1
e1UBSWB5mDv6o9vbJxnl8zBGnMjfCkoryvCz8ZNh5BzNXr/6bB2Hu2FoiE601gql
1TDi07i3PoP7JY+nOygj1f55VmTYMrjLVd2ibIekPBBFAaxzORN/IW0I67OwewJL
jUS81CV7DC2JtjLhgFrHVHj5KoxckAbN7yYFuyyj773u+Ey+S21UXznA04/0U0N7
GQaMwd8JRrz7nmeeXqM7c8cejz3EjUjRv13VVdml/pRFg7YPyl+Gbl6KVwRFtR+9
tWxrdtyaw0xJ66hxe5wMplRr0LR7pJdFtsk2E33YpNN1dSEQ+ymyROel0I6ymCNM
r43w2nzvZoFjdAMG4lh1TgvOmhwpKOBz0A84ufWxfOwX9FzIPOkgd5weTxWZjlhm
7fQ0YcbSbMcCBfSKTsli+3pspKaGoqb5HYdkBcUfjP+wnB4ThH3g1E8EBrobglxo
dXhRwpzII6VHqrkgVQ1MCjI6kOPWUyiSwL4JRLPT9fKEXbLFF4U4nzEMPaU9Np4L
SHrR2QSbBlAOWQU2m9WN6kfMVikrx0sqfvg3EUvG+/34Kj8zHlNqX3Sfa26eFhoo
8CiCp0a0dzgrQuZdT5WxuHjuQi3OwarDFn1S62PKZz0uNUf6BfdSPqpaQFhLIGw4
OJQoNOv19jXY5ukImsagE2/Jtxc5iETH7exQyQEhMeuxcHvWez9HmkEukeROKIvv
aL2Fz9IGXPV4IpmAbrrqddWXknp9XHtceOxFWTkQkfWlUqtOh8pUrTPVjgXx1uHG
J31OaheA+rd6MvkeUyrD8O0wqLiKN5vuxW9WlqAlkxZt0HkTFa3v3xOo43fIvPnL
4AIkEBXA7xfJXBFxkAJiKv6DvYP1S58E8xr11mOp2Js4V7iIoYBeYqCjYJPIgYrT
zp21HYEyFMDZy2yIqABOJlwwOMDj2lM/jPCMVKCisw5osTAbTn0SiTL0kkKv2/YD
RqjT/iIY+z96tZggRGBy5/dMupxZ6vwZJjRrMnBtWJ9Wzq0FaI1z4eLcnJcnpFo0
vCiQe3+ou0wJtJDUnO1Ox1SWs3UObn+psSmHQEAbR7M7ExQxVaxxmKQjQFthoS5G
3PbnFzNw976Rux0gKtJIMLUUuIDLURLK4h9Ah9yimMQD9FbsjGAssM3Zy5fVSbna
7FiKfjIWIaJrCYCWwqVk8ySi/Q5PQ37xbbUTQPa6vyb3sp5DCZVUGM0xTc+It3dW
cs355ti1+51WJDDs7MI4ykEAUYMJWU4pSwagNJ8ekOlz2kfatDjDqqneJViW4TpK
XhCHKQTiAaNyIgx6ptDA/7j8L1QY2VtBMcCstSG8xNRuk73M5KQmM/Xrfj5XtYDR
F+xnAML3tVt0/uPXaw5ORi4zwd2c+OxKKvdYMLEirJHWAERU7c8aJvAjMqV39ihv
MSXuc53gB0Hlq9ghVAgme/tpU8BOKkZtu8E6hLfPoXTaCw7j6n+w8OpZOZhINp0S
ecNbPkiJV5qo1OOgzSKpq3l40+0sLF/mcw1GtOJZWxy41vDXgrwKbQZA0wKFyYcZ
vQISOVeIp0Dt9PVf4tAs2lFuqA8yoMe8q55tJxcNeLa9wI1QJSSSAENRWFilvc6o
GJVUKCXeTZ6pUlJSBpnrGvb7sTor1Cbm+KpH3AOGqZXQk1L7tOrVD/fqXfuaoiqf
+Ssq4rNfybFe/aE6hfsFXuAiRxNtx357QMnae/q1Gm2HbGRBV4A8GscaqqeS+hbe
gHGCeREuw9C0rQ3OmTOQasBUyoJCQT9MEDlydQWW7O4451z/TZ/jKHOip+KJEEop
JWjFZGqK/hxYka7+DbRrXf1Z2fEb7z42Nq950WJ6ADycChUjAD2WARI1tVYzl+fS
5qT9VMzTaV2pV1ANbqd0+as2ZWlICN7uu51CxrDctkTdb98UD2+3fRrscxX6+xCT
ErTzBgti7yBoKwTHvBGYxhqrQHJ87RFoEQ20qotyXmbA8mG+PG6B5ENaur85csnq
VClLWrnx9K+Xg5duFYHIC7ZNCxwIg+ro1UymfpavOGpokjVxzer86qd/qbrp5Ku5
BaJi8bPC70DGoOVXcydl0n1pit0nyb/IGnen2pULdfCvcakNQkwS1Z2ooDpUq2Tu
gGd762jjjE+0wIwsBlviY34CcUYF/TAhK4gT5ma46GpsmZq+5/uToBSEJic6EBcC
Rz60lKiee9bZ8W4Q1Zwo7/In5rQKPRcan2ZSBNly5lbogqSv6p0fhBmzy6yy4y25
hJet1UkaJQNncJT6Iio5OBGUEDZgcAvZl96WTtaN8PfWqOOwtRYR46ZA/eWtPVGK
VT1bT1QoHE9rFvW7St+pQ35vzT5pe1GeoVD3iKsBSdyYm27tvgdaJ1N7Q3Vql664
is/mpjG38Vu3pcSOJjwC3SiAR9eAMP/ViyBl4gYtVaNTW6cmmTSNa2TYCn3kf8Y3
KheeQXhNbFpg7RPFqfo6V41OKvJ1833m6JY6Vxnf7k1CWySPQR3fwVnglUGGf2GW
g8Z+poIoIS8dEEambjd3mvrx/j6YSr0QyO9CQqdxcMqqt/Aa4C7oBTxryoiozwrn
c4rrCcXr0zwFy8ZNks0T32A6OWyiHrvgEVCOwe/SoCoVfrk+3h4NQmPLqqQIKJcM
3I2svts1ebtA6jRdJ7PQqrrSsb8EXsSONHg8MwJ+elguMXnBdk42FmOpEuP6qYXZ
rWUxZ7hBgV1m5KNb28HDfkZa+ybJVvu/wZq9oFQnKPM4PeTeFw+aTfiF3+1S4191
xuIw1utjtoUtgotJEnS7FBvSosQHsGQOvOz6pFlHtecWW+rd/DYwFgAndeQUhPEC
HLBVVTc6IpI1rh0ssFohUbSyIB2wFOFCKCH30Loz4nGAwMmQYRvBTE59DL3U8mgF
vm43eoP/e1PO22vWjbOt2oO7yRqy5rRkqlOh4bsx0SUK88Q6/r2ccScYB/TMHU4T
v0LUijfZns2SDrJSCYTwZ5X7FTelYNNHWpixSekAk6DiiAPRJPxYleaoYjpRCH/Q
pCW4HVRZKl7E6ji75Jkt1waESTKlHqMoPpcDN9npy5eWfv8N/XipaUXOHiaizKla
LOUV4D914r03dhpSqPGH5VYj16LkbMDsOHQl1g4O+4Zo+ib3HYIwXQ2Fu5BxJ96c
qqYf/fmeKa7hn3ujPl2Vx8OjdJSnSApCjfr39Dyv7MZ/pXxDmgczzoirFD9oPUUj
02XdeB33c3n7cdWkZtWpKXC3Uu7n9sN1lPm6Cl3ixD9rwypeQjtlgmVVr9FVPy4u
OSsf1X1FAiy59W5Kb+pv9dJhlkCTsMahTXxskQHmNDOEzmm1x40f07piRsPYZ5Uu
dXnKunEueGU7W3sKc6yqc2r1I7XYyZZxxEmqxUer+Vh8DeJqubAGZLLgBoHiiVov
PWiG/UDLVFlYUqFBkT9CpI2H1cxmc0FV8iNEm3ISfDU6wZl+E8rXBrwHWqS4XN6i
/HcOlYqZAL8fN7YzcchxbDHJNSEhtRgS3qE7Iek2CxysfFOEpkRuuRyCs1uwfAA7
3sFc0m8yDnxElyv8YfbmnqpNedIxZNFF+rC2nK3anGIfjbc8hGkuog34/LWhp55n
cy9gOg/lZro6Kmo3wARStnzfgtkEz0pYFQV3Y6WWjXgcI7QXzGEssd0WIMRFkYBm
pMKQo5g71AFrPg7mKICo6Us2BHQJmhX9dbKVxkKcgZG2AQE8cJCrDR2+eQjil+fE
/G52h5xrugdnDeKO7ov9dplBm2+wRV0GhDyh08e1AjzXxYjlI/grZO3nov2Q2bSw
LuIbVOSBqa9wzaw2aqbYjV58tyc6b4Oeq+G/W1kq4/Zo3GpGh6dkibPuLgoPy4Sc
Ca9Zx4Nr4FlIofBAFGjqDgjHiCL0jWxncAK93j5feS9zdyubfK8Mj1SjuomSshuL
/4ma0zIgWaQi87YVRzCDMkqRHLJdOjEGurHJqGOZ5drNfXzG72aquOmCHsdeDdaE
9La/rEGZxZr7DN1GtG/TZTJTtyvYJg2I5lj7MZXIs2QpBkUEk7/TUD9n+OilRWsk
JY1P/DbR+lrOZWlbo2an2BJnpfS6tIZXFTUKxrNFXNiM/LZR6Ee/j1+ec0VuvxBm
VuxXbg+a/MODQnYyRH0bJysHNezb7HBah0CHtmM21ImzaNQs6snLffELHXX8S1yP
Slj6tswMTEz1vmp4RtyU9bFjHSN0jaxV98uK0lcswLHVRfDUjsWC2jHoDU12NYmQ
8oWaC5PKm+vTfPCtvAufSHbjWQ9ayqgihiqOv7PRYXfDcdPYnrBX8FCJ1GAH9kkJ
EQgBQwuSpAd2zmOBV3Mtwh47V5GZJC0lIZmWLPmOR6QDny73zTp3YsZO8C2njdAS
KhJEIWwN/6TiXjt1ePNvcrgbHvx4N/JV4NldNQpWnzGxGLgODY+h2DuGZuOmZIit
jcxZFDONGm6rX5GmvuQYm55T1zSf0UX4IXAG2ZE26GW5X69lRhtbalmhqvUGLQoC
ZumcW6tRH92AwVLNbzIM8FEsmwUDZLcEZBllWUg0z5enEZpqDkL3vtQFdJDH+tPP
WcjYN2GzL1iIw7ZqYKoUKUzUv/qO0yR0kEFymTP1kz1q0ILzztn7CY3Tih4sdqKk
Okf46aZ9W516r+F608Y7OFpjJNnwPRXqXPJYMf6tMLtbHgeiTBu0bejRYyKUkqed
a6vc7PbL6yeKhHRusEQHtvc+H2eMEisWmm10hPZWwqHS/MMIo9GJeYmBWSzfcqn/
wBtSG4hI05Sdo9Nded+mCxbqOItD34YRtW7EqucMRHDQjvgaJ81si/tLNZt9PVVR
app/BLregFibzHikeZCanCTasx9cGiUy3jEKwcGQcEYw/3UGqcpRSLDZlXDZBlKI
KwljuZZqW4j208ZcNGFp3gY+Z6r0GuCxfjxHiAMRjff3HVv6kvglLk+hud6jYsXD
nqCxAZseK8VKfqCT7yE5+7TKOFLXWeO+Ilp6+daL4CS1e9lLWbegdIRobF6mgaDD
mc+d7fsGwuwY6aJ04N1Q50zREMRLXnrOT5r9SdZaOYI12rYyOaEW6WdKXe8rxcn/
yc9HOp3F7L1uXzbqgW1zTP/WAkFuXoHYoDxeP+wdNJrdwQq1aVLV1pHJYxnDhJSO
kHHvzwPxPN9Nmi3kFAD1pQuqUeGCVRJJfosaI3j9Vi6bH+WqmsrAs4vExJlV5oXJ
We3K8jTU3dUsKcgEtHW9lZs71oR6U+5XI/7YE06Zf1rOzmnN70nWeLFjPlh7CSqO
fLFvG335AVd9LDK0NZDwZ5A7eftKxU/9J2sYD0E4Ybr0L2dLCuaG3JSFIKUUkj+A
bGQ1kFSMeq/vNtxq8KJ4x92GQxORbSwJyUDuzbes0JJFgGFTvDakzqOxj9HL5T6b
UNhdjbV5jpmK6eFpYAMYNorGy4imdNODYBND59/EKnR1IeVYw+nOwufYRxFCXDxa
UpY5xBZC8yliVEMqpS6fPKyDLOPS0cxJktXCTyLJDPXmH2uOfGmEtqom7YPFfnm/
s+AZB7g3Gm2qdY/ejgGcMqZ0zbwPc8JelTQSOTX6xSDFURh6W412BZaKlWBuHvv/
eEypduzVqWrapoL2IRQNp3DwoSdu6aGl+0fhYsHOM4vZtP9zfmNZEnFzPDL9j1x/
l6NeVGMWFZtvcCDUTAFl2a3LUUSsO3WwHYt99vBCtuCdMSy00OlLbwkmRniiErM5
YQvp79j2uiJs/LNlNAhE0W9VVqHQYP2L979yLw9i9MxI/hbTECjpFNyxwpz0NRFn
OUjDHz8zZW3mxOSfY0aiGunoIdAVUH3uoVj5nho9CsGgcv3+V957sy1hgOjIrfDE
s76keMTz8PwXsrHndWAmKVCAKUIj5sa33LsTHkcV3Q9+RSE/ejsewAYh+sxztNRn
wQlxCo57hveqsQdyau+uSZJr0RbORhBCziwgfHuy37qtGIJM2NZHrFu9VRzco2gu
FF1ug3cxBzt3BwbQwgrZm62oJNhgu16JUmk66iy4sRNYNxtXD2WF5b5ljloKnktY
S7QHqgDhgCLuh7DEoeLKXychIOpy1yjqDM32gRbXcuO9VjDyWPRYqTpURQ9waUJI
er18n++LKHBja4QnCBIoWuO9cojLD/cJY8ctl3kL9qGf5obW3uq7kuvDufEZjn9s
wMB2HDuKQFUqEZqCU5FRl+RnPmuvN1byoHwMfVx5mhxy+W9bizegZPbGUsTRl/BK
sdDKE7kHCTNB9aD3wcWqRi49f75I5jyZwFxHm4DDDeTFs4erbsw+ZkwhiRj2WsqS
FK8UY5k98rt7WK0M1u+dS6NxhhoBlo2sPrT6YJtyXzKbjx6wtdXstZkJUpNYCVpT
re641A8W1x0dxcj4nBjVtO3PIli106uVMDAbTdb5FYojfLFL/+0I5itJ3ZxtSwlO
CNpzUWZXHVwhLsKU4TMLhkNvMLQUn9eOZXuPpDBsErxDjsDBBx8LbPLJlvz6XDPY
EsWLr6Olc+JXgx0qD1ico1P5NWptfF1q2Xm7pg3JGmTiRjObiBk/uXqHKRXvHzt7
OaZUb3AkSUeF3xlmyAnZ9Q5Vluge0kMGw9kcpD3amHD4NJu05Ixg2n1RM4yG8mKn
RItjE3DsJMjmEmsMVTHykUn8Smm3SQ3F5tul3GLSym1K/ZgehI57TFdc+aqV/VMU
MxgLASJ9/ENhUREYPuVOohYiimA9wnvNlENiPYLB/g1GtCaU2a+c3MUs7IGZi7j/
mZF8AQi1tYE19YtOd9XNBpFfxb6Gzn+EhdMnEqZXhfUyd+ov4Wh6Vy07A4Z90bND
mi7pQbHXVI7qdgcwcL+PCnD9ymSxGVsv8wEtfiS8M0ovlC2PQ3Q2zXB7te/zbAVE
TlGdPqmiZbpujbJ7EDiGfjCAK4LZgeD+mSbKAbRKxhEreOwvpwnTnCYfIdzYclWw
dMlp39YP9NijXrlEnSrIuxp4CGkYaJffx56s/UziR/a+JE4tVXxqYKGjhKWzUrPQ
Q/laHevVPEepOgbrC8Rlh/k87TGE5OLSylZrfI67Yd+BCrm+IhBJYg9TchgV7lbk
8KIfksuWZjHlPk5qtMQJaLWLbefYcULs9QKddDJk4KK36TpFb+uDOKtBdKU9/jPi
c1OLGTfBjv6PxFsq/0FAoRnMjolTWpOCx4bcllfpS1e9eZFwgZUKQJVhhaToPPZN
pYwlbIbrq1rSytlyWisxKe+b3eu8E+sT+47BufXDeETjqAHaCQw+MC+RvKBJB7GI
VBZGktBhIsoWi3Tzv9LucxtpSYSjR+dkXpLPvzCntvS7RehRPi/BZo16rj42CkC+
37jCvcX72cieGapMQ/A2CvvgF+W5vjm5as24jLRLAuPv+Z9dwURNum8QHrk3erI6
WBjd47HTwaBtDsDdJPmA3/Ky3b6RXsxoaP9SgTM+qW1VAS5u1TIizyvwehH2ReM4
cxwiAjwEnFvmQQ0ncUE2tXb3U0di4Si42IOzTtWI3yOAOs3jeKgyF4/TVZ5PcvR5
YPt9yD/M+zOpdBqtMCCP33HEqZ/0y3AymEN4RcfPejaskQSLSiGEyN6G9VRNfsB/
qckxEqxTWpCc9eCg2LcXGXPS+M3DNrXpYnLBhq9d/kc0WekId03twzSs7DXdgvsF
vQztV79EmjWlXuSC9UZJMIquEEpFsWn+n2tEE9r+K4tZRiOmG4MnRBIw2Tg3JPnf
09DMqb21jdh0IpYI5iHHlbd3cwgtkXR3DvlexxT4Yic/celm1RXBcz1SYyrrfuUZ
VwGqAsx2ZEeSzcGWeSAcjI8Yv27i/0gdzKIGrBNvFwOXODHEHFhIe+ION6MKoBoK
0cyl9AbeUfdHlWSGfMjnakeNDVi0owasKJDoJ6ULpEMDgz1pch0CDpiqAi1h1Fhc
FehKCvWdfGDGyp62nT8uB7MQFE1u9X08QtFVGJ03XRcZREvCvruSf5tCM0EkUlwD
L/i+Znf2HLJItdHZ2u3R5R4CowVIQRio2COJkfIXFHL/fd7aydHI/Ybf7T0rdRvi
71KJ9n64Te96HNd7Had5kZOaUjQlHZMSZ2IalK2WssckDxEQedzo537vPvUa4Jw5
ZwYPjKd8ndTgETI9ttMI+5FNylfGit/+DfFSqJj8qlOllP4sBOyRnfppxH2DLoEg
kGveDYXloT2RBmgDl+QH/wRoX0mvi4LjfyOTlnNfVqdMR5/TXq2myfD96MjlJjNP
PgJKCTwtVCO6ZpastMeRlWy+svq1Mvsxrd6XuqyNhwG5xKMBOaCgKqNpmDzglrlc
2QI7wKx8nxOhUjShI+qHK8FsFl483+ItGutG1/rVr6Grxy+wQjPdw6bMtzNbi7uO
XgM2ez9xblD0/mtVCZ6W55QoNBDI2rmSuWlvA2uBOfa0PYSF/XqfYqOBorVQjMKO
y3RACcmnFzSepYhbax0PQ8cmBbTltVNGE3WYpaQIJtRixxAb0QfT3Gp0SC5BMzIE
Bsn45YyYKnqS2kZoJi1CuDzTLJcWg7z8/pIzP2AmG8Jc971eN7uOfAn1JKIXvVgu
Xwd7aT2Tnuanog7ws9fMm1NJ/DPthkrqjjkkZlCq+mCuD/v1IwPPcz4vB5LzHX/u
Pw2MXd7auldsqtYZY9dBOkO2iB0sKxsk3cphGcX5p7jz2OVOVvz+P1j6pqh6e1jL
bgSIza/8Ucj2+OgObJCxJhMCkGWL+hBKNzRCm9wDRTo85FqTKsPjFle1BbYwQR5W
Mij0DIURZ2hRQFnOhUySN7ZercgiAbs+4OXEY+yXS6l78yESfPEbWFkIT6hEE9s1
Yp6k38m4lcyr2+FIVoqemVwlLYzajkKVdDOmpgbx2VeJZS65j47lnMTXmiY+s1s6
9k3+QDF/4kgvwiX7znd9QAzmI4WL+JxuMWcaaNiIE+HUKLF1UKT00ctQfDypGLPu
CXPF0SkugcNlMDHWPkaMpzFwM8FPW8G6LgqJy/6F3ihWjXX00TEwoOoVEywAVoTj
+ZD0fKm9tWO4I3fcLEQ6Mp9kB3VDPorSEveEPR8FVM3O6pp9Fqb1Wkfy+aU2ZolV
+q78Ddb4iqSE8QvVQvNPCMo0uhFEXiq/7VHF5+j3mUfvocuODiKMIT7BR3l0lf3A
MKAbeY9jjLB8DhOXgIJmIbXU1Klh/ENtW2kt55HbafQskyJ90AxxrU1UMNNm0AJl
CJT/PexixlDUHTNWRaY1zaANfCEDOlHPND7aECqHK5Vz7EaZ0JvTIGrbjamr3X+n
FPrghFpHbHRHKAQwiTRNXwDMoaUMQSUVE98ihQw9uPf/Az+WLeZkT/CFGhzcUhbc
+/K6gaXBDe7Y/ts8KLbbHE3xdSsLALLMqAjwjRkOfns4tZvOoR+l2dCktCdZy7TK
7CepHauh51STHlUIFYDgwHwGWb7PANjgBcrJY0lMDqpIDu7NwwWneqJ1lrfrlX9e
q4yudD2qPXmFTf10paqrGruupkUhADxvIs0SPNuKnHYt6oSGOj7y1B0ks2M6fLWg
G2pXnnpuSmtyPhGVvTV7enGsT8ELt3TWU6jzsvH5Eot6ueOBg6IrACxxikXfe7xz
OjGdP8gtyU9MwWVGI0JXCm8MYpUorHXdONS1OvsZF5LpXcUFnqTDx3w/EdnTgBtr
UQ6lvK7FruvgHBE4SX399M8V1nDilh2MW7V72UEIKjKywANy3fQhs1o4x8uFwNib
SRE2yYAuWLNAkBf6mNF0ak42xyYozqM2mayjtipZpE3T4vPFAAqw81VERohlZQYO
mXt80NPKVTIGNJdr5itti11WBaEmUSvFd9fAlxNfu/66ZNUHWvXDBo87UzlPe8e8
2cQ14pVKH/IF7u/WAW7SFUISUKh+Je70KjHeQsWOsDlgdBbuixrLkCYUiSyc2ztR
8UUr8MUzuXPsB5vKuJ0o9/1dEwlxbESdZjS8o+5HgfxwYXZlgSw0xDi+P7fgF2jS
iQCp68NCRajii1++ZGu1eWBbkO1znGVDnsPa6oFwdQzJUw6DgnMyIyIfovOMBvjN
H6Sfh0I/TTYvCj255lJdcBh66nRvMZUZSRGwEjwe2jHDFVIgdn4FNJkImPZkGh+/
sowkFmRlFK2l5XIFCBdBMDxm8hwEQB9VejRDy8UlcXWhRB3rkdx24MRg8YRYLaLs
SrIQpuBrM3rG0dXxggppjz5eTgAreTzvj5gtpWbHpD6iQmx+NWjadBrK6B6OaE1k
sCiuUBQSdMRe8CpYZyQEYic9sT9FewHdeQWhl6SZemINWCePXHIWY4OQMKEJy50g
8z4z7SYagV6jjgd+35Fog8LpfwO4H6c0zr2xqc9dE2xJ/Rs4Ahx04E4YQejlKM/3
NyxYMwzFk1le3GGlKapUiHzwkbbOigwSM08srxTNGwDN7skkfi2vCergwXtILie2
6i1uTjfHvhk6bh59bkvL28b6eojDYYZJeNy2XfmSkVIHoAWohFqfBA10DF6n9G/m
GT6g1F71fQxf0YAATk2KyJV5RWP8xeqcpZE2Rx8xZ1j3L1xs1ib3CUNEb7YMWaR4
h6KgSDx2hzoP5qMscHDdQQI9KWrsm2d+e/c1VVengEa1gLvwVQoGg+c5rVZnPeRX
KSt1m/RymaLmV1QDmLS/6sF4JoXV377sh6qfbcysppvBnWEPS4HYfqxBMkJy86wc
/Y1qEp1BqW+5bJyVFA43zhouKmdNSiOpjF5Y7XdA5L53uSMH1OzeBA79Ig2j9U60
mQkxBA8c0t0b1BCzGf59CFNuaocpyjG4JbNC1BrO4M/aa9O8JdcWWLJoRV8PNHTY
TVlzGeBq9UG+gwt+x19RQ55KAW0ajaZeZUDHkndCVtgB5MdHR3iwqT6WivQbCxyR
95BfrAjlPI/4tHD2M4pIFNI6H0OPnkv/lhu6zuMnqn4e1fNU2Ka5ed2y1vQtweU/
2GsyzJG8s0nU621lpURZ6p5wd3Rx4PChycxpglthVLWvtyTV4/2kX8b+FKEGLa+l
S+lX1CiPdHMdyGSqCInp5X+SFQkAVqY6XCjTjygrdq0doT8tkukqPdyaNWCoNsft
9lUkYganThRrms/A40XxVOjJQQFsSRRjgim2hnKliuPlurD1F8G2dKHCcvUZBNzs
GDtKZrmFfOuE62KxiLXdgzd+D2DWxpR2FeChv0MfzCk5kg8a8qr08+BwkDLCcNFQ
k5OaIoQ/oozdlC2QteOLRY1N8RcCOfq4yLlNP1gKhVvmQXzNAdug9jpSt4Es3umO
A1ledBtlir9YkHNeqDa0oD4khEcV4g9jEhZmat1H+1kQtkO8Z6UZ2pIWpR4HbKpm
OT/8/PLtpL66Ebz14RqvWXU9qjP9312gINPAGotW2rTiuCdEPGMdgNdIAqiKathG
XlZbzZR3zHfFzCSG5dNVAfzmGwk6pRGvatEVxo4VSxcN7Y4u2rUjUYV9EbqSvR2j
MOX/uOTBtLgZlyGHGOnufKGT6yiAlE7JkMPLYxUQjqrejWfTWT3nqMQ8gr7gGh6n
zpabG5w0HN1RucF3Ec48Co6oQaUIfUADDad4Y7w1ndjCLqpDX7ZX+ChIvw1J/mj5
uOrKyNU6NJQp387BO/Hx2Q/RfLJP4afv2aa0tDwAG9xOuPNCEnEYnILT9jyMvuGC
Zyxb/DhK7SZ63/Yd52bNeqEfFNtN4VyVLC3Jt9axFEw7/5wxuBvqV88Hohnnbtmf
uLBVJeEK/Djetkn4gPs/EkMAhuqnp4Ftey1m5wWRCFJDogro4cAv/iIwpYNVgnl/
t0S8xYznTi08mGftIsbAH2bpDM3WxXfuAftadM0Zj4J97tN6ph6Cy3VATaNEIEp2
kO1iLeGGK/UrMDRqNm7SLkwOT+A529FfGHG3fprsbFiFNNN+Rsfn3mYOBMlMQxRx
vVOPfhpfdoOYy0B4jFSlwEJMhqwoQ4jhrKmPZh8eT0kRBd/GsEg35cGfDPGo8AN0
EUkj3SIlpA+KQqLcieAGlVWFaDkco18rZ41G4Y2giqUIpH987udD6g3aR4gz+4Yq
7A+XjaBccySzytn8QwafngAlIkCIhfKfGTX2kE+pH1OmhLZM6YPtiI74X2YrYla5
8xjhGqR80UHudlF3ubCFRnwx+eehOcuFlWIz1++cNZEXeFpZ+panREtRsl8o4Rtn
dOS/lQPioaqhOq7iQZglJUv99tbpUl8ZNyaBugIyaruL/HZZfs6p4uD7dvYuOp6P
TOvUlo+SOpXaf8MuD7Ec4eHju0/tggyI+klWXd63XC+nNDInCd/dSi9+gWoqtRqM
qEXPTeRs7w3zd3fw4z1G/E69riStA4cK/V2KAw2GhBz1xDiuC4fapZ/j351hmBNB
CmwQdjcMdngUIOleIEaMySkcV9kCqbKu5jwS8JVg7gxFNjbQkW6eP3Tst1c3jFj5
NixT5oflLDGKv3LEoO/k0P3ru8csM77JMBUvYjLk06q8/0iKR58DanXkjEbcxwtS
tiWDKwpYdBdj8rq0qaAL0bDmzhN8gAniZzvFSxhKYWFPKItIpPJnG2QmK7B5huAT
vAw7zto+fVUh37Z5IWYnk5KsayyW3JTMLB+nGg+X4HsBZBf1E1P7XGTq8mAOSF3x
WheqVIOcMAWiiHVmgry5Q4rMqhfu64wsdvA8UJvq0JQph/jWEiV185JCbxtzLNZ+
TrqtJcVUEeQTvcxsbyqxW8WNbP2oPuanVsPoIGzF9I9W2TOSE2viiVtocEq9Af52
RO8n8usntNDkjkVYLTAE+uhBd8eoM7zHMkrmBjMnClz2VkaHpZG5RsQZjFC4N0/S
RhOqBOxEUluUVe4B0K47SEi+k5YrV0K3aMRycCOJRJ/Sfq2jmWsMkJgYDIqgrEsS
fY7ZmOkK6MCMR3xs5TOlPmi+1EIbQQWqXBRSPoeJTChDZ6B+vZKgtxyl6xVdaNZY
OSszMM2sv7fInBR9nXeavFr4HjUUhb/Jj61s/m9l++Wi1K38qxDjxYzNIkv8aY1v
Pxj9DM1BLJxdlNAhEHLmSpq55Q0/w8v+7SDRXjU1GTUSXI0IwAV+JmZAHB+Xa8zP
eZvqqy7LlnrkzsyLHjTU7AdrF2ylBdqvOoxVMp8pLCE9q0bU0ucgTMDKIt/8UVrt
TeJpYVDkhbVECLdb3aVTmMT4G0t++ZgYtc1Pd+k4egsU+NoTsMI/XWpr3WAHSc94
iUn1RBbklLo68zDWeuBC+tXsjM7ch1b7ubjoddVzRGSnJL8RqHX9TzQAG3tncQ/1
7ehBkXotoIrK8XjRbmJboDvVtk3VRr7BKIhIAmuKzkEokmfgKxMkq9SnYrxdIIAC
3JIg2ZtgvmgUj1M2MLpRB/V/psgjscDRkIFKEqIOMzcvKJHMTqzTUgdbWHAxdFNJ
F6w20WA20UkaDPm6GUjpqDIdwmr1i3aismzWXKrolEyE8Sa+7ZtziauWnoPJupM3
6/sgGp2cnWzUyM5il4+fjPYoBe66b+g1I/JfOSNeoBV16DZwZVlf75rtLpaVsetl
a0G7pnDjnFfFk0S+cWdGTcNARF0RP9EC08TzESMOPZKyewktge2XUz0FcFFS+vMM
Go4jBXmdheoomrkHpzCBpWDMrboB8avPNutjjEfmLqnXM/UvGnIOV4z2eI95R11S
zAh3v4nCa7clljBkcrjL4nxrJmrJ150z0pnwB6rqq7pXVPLCYSEwA2KBbWSf44b6
oTsdqIuFPnmixecD5QJBGluqMfDj+7T5pf6q3UeExXTy82pF7y5zfa93CfcM+yF4
SF2ScCCouQ8Ahuw3rVeljomE0LmnM298+dYxL1CPw9+NkEglOQ8Gkg1WwD3RHwPE
dwXxPXp3bkwRnVnqoGhG3Vg96iBYsTsPq6lsVvu9crH8z1xGOqUXmqZAbGE0p1Gi
PK0ROJyKF/d3chu35dy2S0H6eXLB+c9t7MoLLjt1ngNWF0bCn7NvfJD1O/c9abX0
vcukbj3DrBl8H848QpQTLP07BK3LQoBVSCTRY/xogM2gcAHwejh//ypXCINsQO7n
JGRq/Qfw6kKfJbZpNUmouOKIZlifi0OL2nSgLpvTBQDGP9daNruIEaqYoXUdUfKZ
/EcuBubBZnfZ4znDkzWRPPugHahSuDnKogP//r/IstR4DtesNjaUYfTefD/dd8mk
XbP6uIpkEZO4z6auvLgCUIWmlaxdekL4VnSaibjcotggKdOSznKIHz1nzw+aLQpG
6+oYQCNLMAQ4kAlpBKll8aywczhueGqyJCe7gbsnQU4Ci3otjLDrYd3ljU/wwQwr
Qu5OV43EQIx/3Ecf0s9hr5vPT9W4h8lxFJAgVp59mWgCscub7SWnH922KtshtbMn
ssxz5kPe9WmPXuebTNR2k5Jc4q4PANw/vGKIN6XSKdhRVHWyR5BBRTaKJQ7uatNB
mv75IhECXpIvCwx3OmrEQViRrmVG+fm/oSwy7oQdDBcOkHkvdyxa9oh6S7D9aD6R
+YX2jQKkc0WF8qVDXnXTRvZcQH4o49b5I29XlAt8TNzZXEXeJ+VOQwvYGqGcL063
ICYYDUb2cbbKLsN6oRjj3CPw17oqrDeFwGBwIUNR2MxVn1NKp+L5i7ka5/CXA0d0
NkLFNoxFhavJmhhv+r6oLLWuL4bYvjsMkSxkQOgtnyFTd4hdn3w8Kn+amq20etQO
+irdSzf0ROp5joMe9pNhzezIulW4CnZeCwtmNc596n8Zc3KOkvIxGaTdIksxS/V3
8t+5MIcVwX7oE8IhC5ne/wKjkqkasVjQeETtlAmiXehgy1+EYm9VLLMYvrY0Kwxr
DINkpUINjpRvIdJSYWir39GbAeaw2MpVpBiRXSygPn2DSFJwkJBkD8YEMY3QUcDX
w1I84kx+ohFBSpcXWkgV5iRIdkSXcJfbHlBkrw0/5xfX8+rxb49x2fQdw0VzzMOR
skEClDhxdZIiFW4CSrjHdIs7wvtlgONvzfHaEF9IHbRH34b4tAdgJqDW1b5Qt+/r
e6dBBJqpNKprruwUhHfglU+l3DzkQiV9ffrCi+KUoQnQiL4YB9ihGxtY/vd+0CVo
a8nM+lB3lIqqssTzC0NCs7FdeaWLTXOoX/vnV8KxnjChg8yJHjMzQ3WsSP0Azy2w
WhSeh3VMDRu0umzYnBxdDXimorXuTHNCiSgRz2+dwVDtiJyy38BuE4F4qVtB5GYw
9Eb+QG62MEiokJPKfgWC1e3aiQNYaQdi+s0+gWtTt6vvYepldu4dVubn0T8Rv6ll
ScBPP7C8wAd6m6fV46mqMth0ZKb9I7cKE659z2Xvn6B2YpyDe3Fan/tI9SasDhwD
IUROPuBQTT9YwIleNQMtzmwArmZY1GqVVgstkSWRnHYWXzUdBWfszBYbW/mD5TH+
zGds+KRin+msmNbKUQYhV+ZfCvEVegRV8xengOnpDPh3/buo2nrTuowc+JA4pZ9y
X5ZFvqHE+EPfm5uMpcYVMK4VHSzWer1lAPFvKDWgTEcec/wrkLRZAsPGb+b8wMGp
TcyivWATUHRHsaMNI4XTiw4y2cF235Bs5XySY+ECLiOk2TroArSo1IYZ392Yq4yn
6Wpobf4WXZ5KrCXSIXvACaz1oif5z7c4Oi5+Pd1ygmXzICkpcch9dSM/vFvz58Dz
tRwR0dnNik4YAjXnzfnbZfm3uicolS+Lj4V7xPZSgOpp+FqTeTVIyseADvSOGq6t
WRA6RnqzHpVhutBx710/86FdS8smg3FhPNUKSTlYGWf4/r0hfgn7zgLx+UefqYRS
93AAqHPtJtVifFHbaApeQttOuneFZOfKJrWkFhb9uJR2M5ZzEhqUHqYQJS3bbrOy
vtw6JyxWdXCoKNIN4B1aoMSKprohedEsgCPirdLKScj83QX9/u9F9/3jzuy8zJOe
b/Hun9U3m1tMF4M/Atzqb1owlDS0MQ1nmB/54D/tqFYw3aJEU+1LmUt2677UCK/S
p6aznnn65qRjrKMOIHEIYDdVYon0Qc7cUqMb9hDQ01Xo+C4E/5MaBa3dDP/w4PRL
nCsq5MYEamfHAocI0e71PjgrIOir2D+MZy2ldnoXdtlp/LW7e7puYg4qwNji2D8t
S1CNfTwy5Zrax83WxTwpOcXF777jkL3qmAG9oA8njc0GQ/CPORXnfc0pjOwkfpJh
GitkvwxDNsF9XKjhhsgRxxA8YgTmGkIwW6q3vxI4OIQz65VKOUGMVvdgx24Zzq7H
LYsWucm3dkrKIhX9ts+5k6/n5NWx4kJ0/PAsR1TBH7p9AMD488ZzfFQPnbTz3E6k
vpfnRoj/p0pEYtlPWpMaykGK2swm+MmJ5mmt5sFf2qV97uqlQ4WjMS9KsE4ac2Pt
WDaIBl6+gP4bRbt6qA7lYfwnlyDVsm7VDfZf3UrU1wyN8VHRYtwbBwxpOuIgMOcl
foFbpY3Xj4gWoZ15qaX04rBR7/MOIt0j1TTv0x90/gWjPd1GaGLPfb76vScWqUnz
NIYTWjUDNx9e2MB37ygdfyeClINK4uyh6rI2W5AOBymoqRD95fRyA+7kUkLplxlP
YQOCMDenCMWyT3bzs5/ATSL9ammLDg8TclrCCH3CwwE11sbe/dXSkgWbnfvbAjra
wtMyrYSa3p1xurfopzvfeUirz4ZlvVeV8iD/lgzL/vYfzEUQ2b6EdMkHfhc+M+OU
p2ceX8uDg/jEY1BWouQbX76KlA6oJdCc5/3myLNXzsBof4B8eetoU0Z+Za0hFhw6
GqRJCTJizXgCaqZoXkoo/Zq9V5WUk7cz+5dsguNUBqUhAKkU0V3Ir2hjjSxiVYT3
CJLtL0rjjqvnPz5798itIOm8nJwcFWtSo7vsmkO5w9ZZFDTpC1Ew4bUyxFvhsIY0
NOz1dwGICiM0CyDtcUapvYV/G3kYszKgdC/2rnY37fbHQSehnvG2rnxg0DLv95cJ
n0PQjjxQADZU9Xgc6S8oNG7XNJbn8AcJTvEFSgPUF59A19pJWwAvtkIas7OoQ8uN
7kqUKMWrgBmjxipfcOeMxKjm1cJGgBWcFvXnJQq/vbNJ1b/kvBM1pRpcOtPng7Ud
TyguD5L5zg3esLF+Xa7p80E8Ia22tF25yZFdNW4VJn2xhxnfWg/B66PaWABzpKSD
p330V0JbI/T3HYst+YxgNaInpX0l5qQqi0e+G9IB3C3CCjRoLIynzF+5irrQa++E
tsPXSRDW5Ejw1tgq1ujvLteH1/NlapLSy0pddne+hk5TKZu2r6PrtW+0FCbwuN+w
rNKl7uuAXaYo4rRLi8feAgjZgoh21t6sZ4anz89EvoJV4fYX3DdQNH80ho+IZh1g
cAz8kMbKBSfixwlIpuHCy90WLAovMuhQjkSPY8zyhL8XRk212gWpmTdIgsCUcDQv
yKsO1/EAP9xHq0hhldiovjryUvsgCJqGZ1blUYZ6BbHhRDo8dfj4mP2yB/zTUgXR
c0BnrMiWn3FO7MvFEh9UDLwgx/pubQfFwq1zHJnPfevn2pNeFwY1KT/p8MJLNkL7
7j2NNEGvHXRJiCbVH2O367TahBO305gtCSFZuaMTvFEpOE+N46IA5lnB29zcCN4f
SR9+L3euv/LaqFS7Yr4qaDsqgEcSHRMvj24vayPXChjVdZAIzITXyGwIWhLr/ufo
1TvDZtAjBWHwo/v5gXZ4Z88g9Bf3IVnbkND6807PvP2EfV9S3lENTfqXSon+0mNt
jgwfA4dAnGKJ+pKR2O43TtU3ShiBBCRA7p33SPQNAw169KIF+yq1LBs55gwHDYBu
caay4YFUVvoIL6qFAHUVgjjWXSc+kj6lP0xcTPGdRkNyRbj3XWCHsX7alNcSVmg7
a6Xxz8KvJ7pkKC/xNFs/fVSg3Cu0+hjRhwMv0U+3P/UVoURCRgGi8YkV2ZDjBAmV
lXz6Mw+Xe2vaZiHfP7rjEiFKpJNNNGemEOYY5fwFqDcLGpMkrdtXSZ6injP/NWfh
QhqJX4p+kqE/XZDxej9Z8u+qG/A3Nno1wJrKAFTwPYduj1HopKv4C3sqTAw8n3vH
GJSS4r71uxZ0jnFnWqC6Q+6+mh8cQ9S6/Xd31iMsxGI/Rrpa9/HAckM9WVx97ckP
LI1+vmiwiA1NJ1fQXUby0pZgmW/XEINirGqjTtarEPnMFLOT+onNTp+yE/VlBndk
ne58BIihA4n+d9IfZsDS0sfKzvR55FEeRV+jJHQRTEk3Ctlgqmyd/K6lOM5UjvZ/
ah4RvnHaNscVtdDCfN8KNULwFPpxxZxQrOq0WWD9IyftG4dnAfwvaBpSb2P0hFGq
IqahhbTFQQtXFtNIZIsWe6wL1C0EkxNIA3+kXFk1HxGOHr9TYHyiA+WfqvYVeFEX
rOj+77XQ8uUgoKvpjjPB26eBmKYH9cAKshfGbeP4vOBkM5qfvb4oZ2NcxnRhle+n
H1PolqFSw17YkP/N4MmS+axcb0wava4RnJPI/pshEVI1GZ1JZ7J0PL7FlLFa66RO
LMp5hycJwV3HUjh0MoWfBRjAuh70UKv7Mc7G+tQzO80cmnqSrABXXkd0buAvpEMY
psu7cngX2vbUsUZ58avrOL4e2QbXNiIQCBY9kHWj6Z+4QI5h9NwXgSoyW+ngp9Gj
QJ1DCGW6pqfVZsj7o2/6FPuri/xwq+KOYSiB9Ed/ip+qP3TnMLviWHxhN2wtScDC
mrXYhDWouWkspn/6+xEr678Iue1+6GpFphq8agcMZydedysN/OHFz45Fp6QNfeGL
NXQ3GNbJAp0UVi48CIheti/Q4Szo5w1+dlnrn+DouZA7xS7XDKYaPa/Y4vkmRTGT
Nyrw4OEG5/zyMRiel2fQl/bNu1mZNoT5Uys2p7KkrFIyQYwacztedL0U5tAb0wYq
DSZofzCrTJcZ+PekbW8CJU+BJGSPhn52/Pke85XW/0rRVRx4PuS/eqYdhHR2ba54
eQnShep1Uc6Db5VAVQt0rsJwHSKrOUmFRkX5M2oB5U54cMUKfVQAznPEvaMZCpaS
fbugKKJIJ5+mD0WJtYKRPtEFFvuG/swufaiTDh7D4MRmnlQd2HLQzF9xNQs9R3Og
qsKYXU7RV6AlxkT6R+hP4+BKOSBoRZY8ZM2klqh1xrqrCLAi/TPFnHUOw5kjO0qs
PNirC0srCBHCP9uiFGV0ZgyrvQsNA6SEddyh47Xn2UdXcGsMLwQ5/dgSwC2XGJxy
gF4uEMzvJdducSip8Jf6Xq8dAKy/vdOgNWesb2LYlcBRjYG3XNlABi6ey9UHvvGj
tOA5YdpGmoZyOOxFlQJNTWzWDFeRhtF12+M2/pMZv7rLdI9p6PVT/SRr3399zlhz
0EWP0OOeWdG+CyV8Fw6P4VBYu1ujhKjAGuaZhwzaIdWg1l9dczW9myXJk1MF9/pn
vn2WXCmFETLkEA0gCfPBLOaWC+QYKb3LFsLPEHkPDwlh1LHHKutPEA2jFSKUWPxt
fqA0ezNmejPr4zk/98YaMOwxHS0KeX7tgjzWhzbR/g5y993/tAQW/726XKwTUZKi
+e29xmzNFZ6sZIuIGW7PTI/8dKbELQ+DHwUCB3Udb43yCPWXNw8hRJe6VgVA62TS
rQt+I9JPEdZIuScyywxAIy0kkHuBUHZhYufvlMZnw1NdBypLLjyq0fJsaps5Zo48
n3Z9l9f6aZw0Gi8crycIU2zbpazPeC8YFsjaXclYAA0fPfanuWeIGSXkSCU/jbHQ
bRNItWMA9HwwQWqAeb6A6bUoZ3PVvSQwfWZb0Y1QRPjBjswTc/egMFDQb58N5V83
hnDo5V02rpD8vUR9PwOBks0emp1jef6MJDo0nho8xB7HtlGcCnB+wYRQlc12BZkn
QN7JtjG2G62vak2GMWlc95CRIQzuXrHYOYBIN6EUqU86WOqgxtpmRlzoxzEPccYJ
ZgyQThXdgeXFNns+dqXOx9ZLIZMhWgnenldFWh6jrWmBJoRZW2yP0UnowPHYnXsF
GrqyDmcln4I0v5avLAR05Hz+sdt1xvpdBmBe6B1MDGI91+tCDk1+kcXvj++kb9rr
Z5KaD2xmNsLf0xCADzbkOyGjhgeskabYDK0kG3wZ1ZdTTRYTetmA0WfSfHljme0k
/DHJGShM+y6dwuu8h9vxrz9DDIYFbQHAJII+UbfDzuZ5SGWU/VhR2oeIcV1mfInS
QRp6GI2OH5WdMFhzS1v4gr+2nR2qaGN+fll+9A7BAUVdtB7WMHeEj4qEwV6er94J
F/2hv1xT0nzQpnYTvf0X8kTggB1LAH+EprRNWsHxkTxUJOtLjNk745Q2ZLNK2/Pm
xKoyJ9QwwPto6UBYovl8VMjAUpOCOInUte3RXdA+mEtRUnw+4yvyFISB0Vx8xXpr
CBpMKcEuoUAwEwqkPcy5L0aG6CoKLWuV2pSiH2wZeK6YGRnPSoMSfHPZKf87gOZp
AGWzqIMrZXnDXYkN8rnsLZrdhDvAsnYAlCQotQPOI22AhNuDj5XbIaJ725hFbPdP
UjyA9h27+Y2Z94Wj7AJrqK6p5a75ZnPIHrdUBzPokTxX8kT/McWv6sYOyS1l6RTC
doDqPPAacGZy7GJQohDcP/k1wYp1DmVo2ixj669ge3s+xDK3chA0MpM+T0Tip69i
NH5djS69UMgK+th+hvTVb2sZQ+VhPVSrRCMNHpZ6+FjWFLRESI3yGJ61h9wK2f6g
PDqGe9BQUyL3N680M/Xpj22T7mV7XZyx3GItmZJF6quX76SlJMOk4dyPfRQHNzKJ
REvW3MVHi+kFPcUQuHoQlUKFax7CbDQiItN4kAdlSDCd61aLRvoSmglIWZNngntF
nes3KAwR+pCbANMtOadMjphyFXP0eHG8nhRMubOYwJUGkWZINgfjZfBptzoD1XDM
IjBkWPiTzCG1IhSbp5n7t2HPISF3fJXz5GMpU3L1TgY+gZF5fYoMv6YqDTSinszD
AyKeVLWoXuIlCx24O0L0IoFBdbDbnxBqREmjmUUqvYf3Ono3/hepYx7UMuGgn3V0
ev3xEOdkD06R/BwMRy4HaXMwRdi88F45qDT2/3l8XWxbRSLVpNGqqN5USIYIv226
Ek37VCpavcxUnSIh9o9IKD8Q2/quneKumEdJEnLT7l4fZWwFX0o5DnHecvWetUyv
nqtUn6WInkZSM23l617QX6EjCL1823MDz3yX9sUS3VN//oXioMWj2TeszKE9PZxl
vpXT0yJyLOXmHl4uMlSqZwINMXsx7c9amLOyuZSGdMzzv1OBwVeedKwPwPxGcNFH
FrGbzMQ9WmJIkp5E3lXlyIv0wggMcPcieWHUP3ph2YoTzRgqX+A+SydhHCpmtRNX
ru2zmr8NhR4Ub0L6c0orLz+i6CSXMjI0XB/UJcyp9XcairVgELI/KyR94Qpc4Toz
R5vJZBiKe1DFyG0cMf+vNlBBAaKjzH8cKns29PnrdJgRUoGHwAObM0nLHJ2Sl4i5
v464qsftjhixNmjYw6ZuPLFgbGw6iAd1RXnnvz7/2RhSJ54lCQP8PSwkrBauVPtK
m4rRLSmDO7PwSIGpkewXPOAiKqvn+OChnwdWXd/M5i/QrOzFpQDNHm4pqOb0W7r9
MGvY7wAgONqbpvpTxNzfcMc/6Wt1KYDex6X9Y28raZDBChGCovYEP5DfUD1wOS3x
oKXG1Vvk7f5+u4BMj6W5X+Z30s8yFKgr+0lfTDL0R9yzz+FmxcFw0XB+CG7nYWKT
df651Dwx1LZ6nhrAPYTiPJ+Z8jOf8OaxqVFb+1tvQD6pLD6mxx2NLqkAqY9emJNi
Cw/Oui6UorjZHJvN3XUcuGBHh6KxMfDNlAnIg7iLlHjSku2U8bZctji7+x2Nc254
2sOoI71MvaSIQlVe5V0Fqefw4xlHkwcXLc5oqs7lXtI5Fa8mWYcu5r5sCOSUpuxf
/FLUnBUsls0JSH+qsXLhA/t2vZNK2RMSyVMjQ7IXCqtb/8LLCWbhkB0LEkRnKOLG
Yk/AhgLImVX59gVNyvnWbDBjQ51vWraCxKcrWEmUDdIEz+/EXwo1OXb7qOg9eQRV
ke0wRL7DrihF9+icLa8RparqhEMi0jrp1aAEjQEUxJNbGYBDurFnRefo1ymIbDyh
1XuobXj67zFiFDEYxSVYdXjZJHaXiaUzCIzKM/HvhXIhR8ASIVApey2ge58TcUfO
L2y7Dp6QVJrJA9SeKnL9jliFBtzyj0YAcAu2ScHRxPrQfmFA/qfajRhGtKq0T0mH
glBXNfrQx/Xrxsc5RS+pULRuzp5S387Z/RHm2ZVlT1hgAd9D/c+Rjm1qBBYwRzQl
BeBgtYSMqu252bgZnl9QgdnOXMBObLCtKPs0hEoutUwVyn7GDptBf8vZ0H9PVCoC
+AcKN1NJbXwivpjwI8gc8VS5RpnjrEY5nJ7qc4pGyxe78uV1is6aKLPcmPrhXBbr
6e+QTtX/Ol9na63ZTzi298+lhOlt8rKt2UFoR4x9MDz+TNNe97vEBpxqNFFrEr3n
sPmKdMilmuQoOqDILSa6fwu/ipZQantoV3SvhKlUPl81x/DBmOjq0ndmrIJPczPF
X1ZVSeSxXd3YAIPIiKZ+YGzkM4HOnWI4Nj8qdIr1miRUTYs2x2L/l7kI8YHBtw8W
AnSDbBdpF2X/DbIUj4AHxPsDqnbDleuQvqqQFQjFn8my9EPCWIAW0cdaCS21ynw1
Ol8K5HfhHLQpBiBpurWc99YlpC98tFwK9uG+bTpzqpGXPuVD9zQEIV0M23kwH6du
mSuyTCv2mcBdwYZFt/gqQhn+f6bmLyfu8e6IW4bLYlrnCGkz6KynuAEkLVwyFdxa
Lp4ldrLoB8NgSJ72J8Rr0lHp9nDC/eB1XwXgoS5azWF42dZGHdHM0u7+2/9J1SMx
tr7XFRVsuXwsjhJy7KDHP7NLP/w00mjZx6XrIieVFR3Bpf7RxoyvyCDUJYZWI92w
6qIhfQt4UPQZTKRVlrI+YKrn7aKCrQk0XsYVwZGzUfzPnmkq5zHxOsBSZNLsxQPs
emutttj5q7YniWWN59cwDf9XG8Z3y0nZbGtZueSUpGKb7JsDKbyvJV1/vlFoLjT6
2xnl52mJij4ISkqCGG86pX5rCl2Tf1sZW7yh/gAcXgHsN3khF6wPmE5gEUsubwUG
kTr3chowAXMBF6LNOxL2fX1ZGnVhZCAIeW3GxpPzQQLYTN/EuPrGK6FIfiJ0DRXv
jRZDU1tSkJa7/Gcv9l2FOHqw6DUBNnDnElpGM6MzCCX9dttpZYrMgRwJF/EVWoHB
SKb/SpONuj6h/bz3Ic+olz5rmlIW6PQNmugwRuLcQSZ6mdAaDuZSQfrlt5yams9F
Pk9DM6vtFH+Z6pXNtuYUN1n7RcYYnpC1TjeZhsXOWMF1KoYA971xfCp6ldcD4Qd4
DOioGQEssTCAHdG3LWaWB7UrbDZbFdO4c8DPTauuBjVvmF8J+okoO2ppTBxoCUr/
RZtf11ZqHl1MmM/Yj+AuYeP4tkueaVJbV2qUs47uo1lbcNDMZLd2uBEU2V7WGcFn
EOAsBhHP+z7qSnkUHI0S6sOT87WZ1Y5BPq2aGCBIddeeufe4UR1f7qlAntz93RTq
RSjQ+1wCsTk5R41PvT5XRiOa+YvZae11GtVTzefh7g8JOxBHePCWoGsS715LxaW2
5kEUFybdIkRDy5FrFEvGe9GjMTZypu46JF0U7nWJwecUdepzMBDebngLE3jv+OMT
tMq6gc0UomsphIHCw31UePgRatvz+zEqdxsoepxCd9m+UVBAfGA6yry9oaPgIyuh
OGCXNBlSPMAZflIoEF8XWHtEA5uBGpWv5qmD+PglJrGGX5uRWQCJ9+0oREL1hp54
GrfQBlaVjutfHGU8ohY4kGYTO7plGliLExHCOWiKVq1OcCpyjDb1wGRFQMXNXWIm
AqcJg1PpuuBIlQAs8bID5c8cfbhMpwgQ4Hym9PEQv5lE4w0+/XCClXjGPUN71FJt
XSovy6EcrmnuZoM+hxukcrONAb/vRwtaUc+CMToFa/bhKwHC6aWcH/SUhOF3TSEK
OqYOL5vn/+a98AI25vYhxJSKT9KnR8bOzjgxUJx046XsH+RRx/DuDOY3mUIf96Ac
HrP7TLC3QH4ZdlcfqIU1jrGa9pRzG2iWGqyzia87ORZXoL8qlEW8mtESoKdYRKkO
bxwuXgGUYaWdRwj26bdb0QH2ZyViVozHEpJR//SPvzIRucwJiHJc/qfe+1uTPdnB
vhopPJyxLtKP1KsiYZuaMMTWiJ2Aum9mWuBt+JJ4vlV+iy8kjq6XcaB5qhuAuwPB
DJYFhZmL/2PVEXpuHzf8vi6h/r6YT1j3rQW8HXRur6kP8eti4lvH6ICGO29HtdsS
L5+NxQbXFDHXph7vKP9qVMUQIaxW4quMdHvYOFUWR0lPD+15dqlcOc2PCMQwYCzH
Gl4Nc3mMxnmkxzl8g4riPpvtUAZbp+W2C2iVoJGR3Hf1orOWkdJp0DI2zkor2YGp
6jtu+Phy17+gWP6lwZRgr7kkKkK/VZIP4BwvVOmeo8dXzH8mErUnwT/YDw//H3Dp
6Zt7Xzs5U2uGrh6KaUPzR7ShoSA6KarhBpMHiWSlOl8Rd8NtO96SQikxuRAdRxDY
SNVSqXtiHuWDF+vpVHiPk126mrBIJ9aoZEMEgNyslF+Bs2fXf6r1iwGNOqJ+tIoQ
o20UMmUqzZd4RVxOF6ZXC1ivBA58EHenviH+ZaPzKnoNK3oO0q4uFcjD11fDabaC
bt51NLSonYFuag08KaXKwqruOFmYCIAXkesP3Iz72/z4vRBru7JFVFdso10gxu0I
DsuQ24Lp2TQ4pHAvfNwKRyMFWwp1PMwNoAw9YcUjaicf1F78xnT6g4PC+HY/hUBB
jZIExkgJj6lMOSKZczRtNvz5uFkcEdmvaThOysvW/QTokzfjwJDzI163tsyXziFH
SdTB6BoS/EBUi4OH8+eIHwczJz5fTRJxP8XttHBNqKi3FpEe021DBmpIKqQCo4HA
8VSep6dTMQEDaUHiVNtPFhRlK/6gMQZmbS38u+JT6A/3YdhA4vcy35StbP9sJAhJ
zMVB5mdVVqdBz6hoLw28aRr+SWIAf0bFunDi4DP0YCgk6gRs69fn/zZoSx7eiuYr
0FS1pvEMbXLZ4xqyYxULKZ+h5uRYh721aSrGCgzFgz3W92LhCm5kjhW9iSjd8mY4
IQL5R0weLKUgOBpW8//l3V4GPtNdIPOzENaUnmA7xqM/7XfFoGgBbsqFRIvc2Bgm
QFhStGT+gHHGyGnQVwjbDKe6H6ulvnLMNf+fY9Gf5HryIlCPwBZI5a4YwGfLj2yn
igJMd6KD1Qi3W4Wrvv1kavK9P/ne0LncwloXJysLnM5ml5z/wld1DiOBZ2xGk+c1
69NjjBCNmSPvN2YJlm+m8VDmWJgPmx4o0hjbgNZvCnUuiwasCiPe5pqg4a2HuarS
fks07+t9ncZ6ThOsFHCZZSN2RkbnwmCHYXbXCObMKY8osY2WTw/5Ruqufa+9+q4C
ihQ1/+LsY9hPko4LCZ/KPEkYpL9QX2zph/6S90TrNOXKTfYFo/lPrPhvtX1uz/a2
SR0k4IXNdQoaFaLGmzNLJYAnzkbGJ0zB7ervimih6wjtJ9S6yYdKNCdyUbh7SErO
jbMp1KXW9PQQEZOTss6xMZRiSaLOMnPYZTY/YJcxf8uDDm79/hT3oF8g8oHrin7r
7Ett43AnsLE4I0dnoBFnFeuJUQTJzJdIDbZUwSRx961yxEMr8XDpXpyL2C1zTZ8W
t0sNWjePWTLmfHT46CquW+aw6+FkUxowKz3AolgIyjD9+aPfhkUmdQZQQSZNNIB3
kIl0XHSGm3GeDKWCrvwoDR5Uc0W5uCXk5XR5NDkxf94kA2/t4T7KQeClilzbU1ix
GABgc+pX8lJp/Yslw8uvJMFE78H/jaCveDcip6pLfddhL+/jwrn1AMK2SyalJanW
X8+DwM7epiTRaH0tMkffJIo5tuF6CyWqB0iZEud+52DLBGcshEy+ffv5Iy4+tsqx
mivoU+pZ1oUT7GYQLj/Q+chNaiopBq+oHBR1cwkmPbl2X+hwKqsylqa9So78yGjT
2xO+ExP8ORo2s49qsPgAkrFz8QUoNOuwXVmJXjnqpDjFm4VultN+p1WUumQkTNnu
kI24yXdpcRdTYkzTgLv/xSwXMzm8IQ5P3toEybCLZAcrKWeXgXtRDERXK6R9A5Go
fUrxjNSz/k7HukFZiDaszomcZoBFKulSmLqDviP8HVnR0VK2OF3qL8tp9GKiEiBp
c9Hb2SzvjgGUMo/IbFpkDIQ7Yae3V0zI+RDJ5INQcsw+jq+co3kfxYIaP2COJ23s
6nSC4Mg2WULRtPLAcI3a+Zxxsm0eNVneW+5rjvQ6pKPDvboBFFhKzCdrLUUh7jGO
VmZxL/nuTH+KcqxYa6FFIYm+NJMdL4dvQmoWQ9kOePMEe34GBLwZ0vCKkvcK2o3u
2ovPmIwwe9RRNLGjNGjiisOmUenxKShtkzX3QKsaxK75FQ3nOMkCrxEFilt29S32
fXSMyqrQU89iAtdlSDT+DVuS24WCMUfN3MOetwOe69TeUlZfdbTTmEdtJzMhjAac
FmPUZLCRefszRmVnPEyZxUDB04oqzPiOqqMa6IimMZ4baSd2kpGD8ZXRpLdZ8IkK
+BJDiPGlyOsB0cVvOg5NI7oFxFhI7sYwh/2f5DdIHMDMqVxLC2mBNhIMU0Nd3u4+
tvUCRc485juSxDzttShcitiHsilWWRO+w5Lm7tU3H1t1fxE154U2FGo9XgKkp7nj
iEqPWlTToDMlsnByHwROzoUVFatPBnQ0+1QhRg9tr+2G/8CM93ZZSt8+zl1CIhMV
nP6l/ibZ7saCAVBq/iychEUqlq/D1Jl4dFxWAsCgaMOCb3IbkO5AB4wmH7R9AYEc
OCP0y36Y36Gy/xmRLMyvblmdEDyCbJ0TGGpeefVfUwJKc4BohH9fb7YB7KUvEbz/
mDNYyrs3TmO4ZOcHkKT0bKFcGNh1naqXE/pmZ+W0KAycBWbkRPu3ROXCUCsxTjMD
tQbXZB3B4mnzpFibOgziDcoRywtCydJeYksVdkLIpy+hrhxHWIQWydKfKeJ+aN1M
Bf0OXNr5s1VhlX7BAdcjeTBHWtV70Vbl3Bf/0axrRrC5ZjtuLiDRICFhZOitlAJK
zuW/Sj/dinSJ6NvyDW1Naet50qyKhZd7V+IRkZfG6OTe0HnR5eMPgh+5p049xfHC
sVBS/xcOl48uVzzshXurwbRJVKkPBm/Ac9+7JrRsEoQGUnQPLsdLuDBe4UENdYud
gNRbghDHuyenZJB17TNObIO/3FYrUSvflNWm0+avAP+fZ324HeMlOVS1PVobRjJp
Xbw/vtMuKwnNXJxwaJpBLpMx91w+/O72Epjd5/aqE72Pldp/7enD7v8PAlRTW0Sn
jAlAqgVTxmM4W2CPcST6IgDsJthWX301qDsp1TZRc8cYyJRq8tv7AsJZeACpldyE
A0GLB/3E8PnsbZNnztvK/I6fJCg3oFD3eqW5Jun0FH8kk1wyq+6nSRG9vIphMhCX
4V80ayJji8yeZduzCwQOfV9Ll1AbOVA0OH87uqvVueE8fvW1yaCvuqFKKjkyeAwY
94RwEj0/xdfG47cSX/+J9/BH67kunFzyE7PQYUzWvYQGd6G19xi/Gd8ztELICR7r
EWo5OGfeJ93khYGNaIAP+HZLSKe95xB/FuDJJpIraHWf5laGilzS7x8ySakmsvoF
+9gEKM19cGiWbna4CpH8Ub/HsTFF9SLxd0gMEnKGmW6tmyFVbTR2aMJzOFgiDctS
J7weFDnS1dp+lyahSoDrakXxDYbIYq7LWIsRlPVIHvhVQ8j5XGZ2h9iUAWCcWAUb
EQVd9lX96z0OAhxCSG/RoOkFUjmPAQjHNt53h5i2+ejrTrcINcsuTTe7LQ76kpzk
m3OMzccsoVI4oleg2zD3WGGrbwuaD3D+6maMMmFr86rpFJKpR/P/vZa/swgYJgSC
BlMQ/H1P4a0ZNsCugdvRRMVEru6o+Sw7ckt8HXo62JtlVWEERtuvS3mDd8xGPCdk
aAiwSF6mhBQ7AazYHVvtw379+xu19/PH93c9ryturWztti6fACNCDvdkv2Civ1l6
yEOHPq46NAx27pwce/NreHEyjWxMH2vjxohHrZoQPXj0/MUD9oSELO+OxczuIhaX
feDwcnCHsx7irBHICyEJBxKI/CY5Wp0xcBp5gROFc5eIRGEKy0PBMx73zGbQw49t
J6d1IVrDaWfUjdGQLjG+pcWNs8RbbgRBVGOfr5KGhVmnHaoiUUphOx0NZa0ISr3i
swuUtlYb2Jyv7DlVp0SqZRGvpi0UzCenercU6+FIiyaOFEZWisxVxFrBazcQvXm0
fliQoRkmR78SkWM4OCNV8JKwvCVtiDKJBDOR3s1BsTLJg9O7BL/oQW+Kyvn503Nm
urIFNfUr5AyWzypaJyiUv+D7mG6wB4IIenxcYMaNG+8FQ0GlckKvFvA5CMHphhKR
CVD9OkVLh7VcfyLcFpZu/aX1u5G4UfvySBSriDh8MpAIkO1+j4x1mnCnpg3+cLyU
I+IfeY3+7+3oKXyqg9gt0JBW2HGvV7JyHyDtK326hP1Uv/SoDRVd/u55TxZB3Na8
Gx5CMsvWXleOMR/852r+W2UI951Himol6aAXWtXrZdL6IAd9waY9yduFlFIVtzOM
mRfYkVpQmZVKFf4P91IOjlKwKkQUUleCEs1+i7c6lsy0TBOHFe40cPCQMORpmatp
1Iso+wKKJO/p91JN+kAGoEeWuc/wcygfLOpL319CwU9E0bYXOgUd2SoxFJ40XXJ7
X5VQmaVBHt/PWm4i4AiKEFqPAUQfBNsVYxtNhIPMZs3rYldNwRzPEI8GOIjJPT6G
faqGF94Y0jWHU2sn38J6dYPjbbrn+SPHl4ntpVExC3xbx1yAW0ELQhnP3WUx+1xg
CJIE/92X8lFjOsOxMM+RJ1e/b2rhy3xnAcKVzT3+XjwI7zjKsVzvUBhqMRNLDVaW
s+zHn0UBIBLBfEEyMw3PvfVTa+C5ASb9ZPVZ697+iuzlCCeaLQOfQ8ZHmy4FlwTe
ETBh2ddEht0UqoOiNcoK2+2zYzl0alSUbbYDvSGNohJc/3GHYUzBxwfBjICSCRmB
Tt7qcy8JBa7XkuvJmGQ49PehpU/d39c0Expp3AvjVO0bdFlMiPfwFR4SR6y82hos
FIwuxkgSiDBErmm4QJd3ogFLETU+WcqgYZYWDm5Xong4IwemaJ3cwlLoXAXi7Nob
tz/ftXn6ilCjJsyjttXfkERXGg42MXPQ9T87rA4B0p1irYxdav7zfz+gmPpSVGyQ
rREolebrREKVSglebOPPMrp9vjCxr7jhS2/hu2n5mXl6gGQe4QTP7sgx+F3GCR35
vd1joYtxOs5TPA7j21Kb0sER0M5YONXqCZLj3rBNjX2A088G1wd1rPi0zZ5bIP8B
mvsFQWVWImXPGpdXNflRRqnGCBmP0wNq5XVU7+aAwGVa2dE2MEJwdEfuHYTKIRjJ
jkznHElXmyZ2o4IX7NE6HUgov+ZwKYWFu866DZAknDy6GIhAJflQryB/Jc+TZ92e
VI2ijKRcOeXfqgL0avuqxAu5d+MFG7vVXq3M3bgjyOIQU4ULhSj+L21zSMGlnbc/
u8KzD95GOriezyPyj1+iGnO0Dm89BGcYEDRjSz8InPLG5ho741DI2vgFUdt4p8UE
Q9iYfRZ9NWndIJrhBg4akWupWQSGZKoXp8+elsj7Pt5acnh1GcT2HchQzlazQjs3
bCf1oufVSQeKuX/9oAXIDVHfX1gj8sQ0jqe6JyloLYgruXPNiBPc7co28gcFGZuH
+XDzQX5Bv5GFF053Smcnb2IycypIWIQFnZoGkNM2lBymY9DP34uTpUYZrMqogvKR
38GuqEUtn7inW38HMchV0oFuHuNEnWz0syjeG1uP6Gtdgsc5AsXmsqi1X3xObBJb
0U7BtTXKZO0qG7IIBRfZrcVQ4m4aoa84k2Pr+pvBez1RiVWfzCsiLM2FwiJJpEkx
XbrBzvPgB2h17XAkqTh6FbMPyMfFa7llaKVwWiA4g+omWK6nJSqTMARqqyTtDjVc
pMCkdiQmdZnpfZ6Wr0uVRtyWDarXw5NAK6TPHPVn9fNZ2d/pNrUwDMUepIITd88D
rJl0uBXyyrlo3u0FZuZ9DXWU5laVxkvG43Qa0U/kC3aQHhoJBjeT6b+l7sJHlbJj
w5Zqvvb62iO0ENYXLGcRaKXVVJMEUuCkpbVRuIzHEDuZFO2pfVvTvb8yr+R77dfM
NjsHQh0/5V7cLmjKGIr/vvIv87TY1ejooGMsmFQV6yvUWdSk4y6E9YumBfguYrZj
pbm3MKp8dO/x2Ct3EIoccPjGHl/FCY+2uuw8GszzNnZx9vnH1TxbRO5+70kr35ZD
nI9UjOMhQvhj/ia6lm9hgCpVQOg6Dwcihm1qRCw+PhZ/7DxKtDT/sKnNbgci2g5X
/EwNNC9hq6mJvmURY7n2/FbXMt7BcKR4Henfo0rssBpiE5ytwMnFFzbPL0yR7TXg
SF0/YuTAHZ/26sJhOJXenJs9t76UVIurGv+ZORwa0+RIwdVCOvdT2aCdt+C8Eq+y
z+W+5NTTnVnDfLA6yM9t4jAP+8qAovlfkO8RMGawcdmPa6BlFIXAYs8Sz0wI+kJo
ms2G90mfLbwRuDIFXh2uHOJm9gPjYGap4wI42OAyJuipKN8kscG4JtCzuLxD4oUQ
Rlh2vdXYYnI4pwj4PkVX4P7tIpPrj8DYu7lgl0JZXYa1zyvcCiU1enqAak//Purd
tnJa9aW8Fc/5LJon8WZ2Y275pYeCRlXCA+MAFhiP7fpZaZ4pds+C5YMG7xFPfoTi
Tjry82lHcl96faQvpUTEvFf3ZiW/b0+z0YyS+lzY/IdnG/U/XXl4avqgNjuwpXdm
7jl2gPBKaXUbINrxW3C+ZikosVOwsbygL1++mTguhEvn4hTz61aaUSiv9tGQzwza
HljbjUmbEOFFb+pFb+Dq/iy09qLFk/dLa1YhkVcLOzzOTlxFM1quyoYxk9D3+8mp
Fp5nOYCDEi8hZ4s7ymd5DCbyaZ/u377HXqjebg1gb70AhndDt8Xp702EMUwALW40
SalqwloO89VfUeUxVQCVutUdqjytT7YUQtUHLy7MelMR1/JNxpWpo1DZWOv1yoCO
DMPySgCWW6PTn2PRhyFi93xFCPJDlspJpfMMzThayfU+8yrkFI/qT2TuxcBU9jPT
CSjocRuOkHs+OivEpFSlQ+kVow2rdvxr5tIVHj4WGPQo9ZQny2v7NjRdHzCtbnko
BTnHAfiW+2/Np+k0Jyc5PvXYg90IVq/IhOksOCW/u1neBw5MCAGSswz1pzO8ZurI
0NrwVoFvAE+bltQST4J29JXLPd8v8VtrPX0q6IXNtc0Yv1/wnFXaCu6QTWtfgq4E
CnLuSnXqQ0R5a4apY2Dy2mmGtHogadh8RinVA5gZsT2LZNBHC8rdEJ/+h7k8gn3D
SRvAGXsubjYcdVcj5kwrOSVd1QuhqwC224cqrH+eSy8ME4Klc8FvgdeqCd/IxepY
gzqpo3w/2vT/q48YymucNLn2ZOB8yDpTfIJvfyyyeFsX3Qm5VTWXnVUc8qb26T32
+eS22dyRCqtVL2TxWWTHNfTdVGPLMAYZb63KifPBMUdlkTe6L2K3hsUhP4qSGVFt
Qa3xc8I5l5N0V1vJfsUso5LiCetmy690yRtvcnyHtCD2rtbAJvpgI4KgABbXiTQJ
ngl+LVa8dbSwl39ZK9GTd66rmKZJMIhkwANcHvRbvgq94M/5fKRNaii7LN0oAqum
0HNMAUaFg9bBLgymBfX1NDDfKJtaAGuiIBzJZRZO27x/5ZQcTLDGDpzRqYn7h3Ng
+FHAirYe9HjNtQljCQivXrigk+HkTSjgReKU2c0CZj4RSiBJMlcCNJlPVdcZo8zr
7DPuukOxF2Whl3eVM8a6Yp5IMGoc2R/mNxe9erE9YPCGOCEio1QtDakw4PDqxyrq
ZAlOUyEop/n7uxLKtto4dRPZ01WFwEXwPZGMEpym13sVERb78lUGWV3LSSrl8CoY
DARq+HJQfn29EzQEG9YLskpNio8KkUM+MBBaX7tDtG1GSav/ZEVKkDaKGGwkqoSn
84IBIfV4ms5FXuwjcsk5m2W0cHvVrlXYwYs8QHKE0LFpDDUh17/BXfWdDjI2hNKl
zzFchB0o12cIWd1Q5bTCKjJv/lM0R4V7eD0tLhYwAyhIS8TUU8gRjw6Npdnl5NsC
V/xkM7j/lA+f05vnMCvBEojRAzkrDyCSGD5nq+wVBpYPx/YXsACXw1pJHmYSX0iY
MRR3rfCilaLy9BpRulXMJZ/T0tpxKqszO33iDxkSNmiKlpa3FlDhVMohKfW2uEwI
SscqmwrycgcRqRSIiQYg7L1R9Ubqtjb3CoFxZKEexiJmwAWAdyvFtgcipsXfOYVi
uYOHRiA8kxxvQeuO9hL83KVT4d3DlP/34hKUYYpWqZ0PKfyj7rvU9i4khtr+Na+j
X6az42JTlJ4JubbWUjzK6/B2L7Sjy2ggE8t1UAzETpyoJSV1IcT08Q+C9ZTlr96a
kyDeFf78KB5LpI6mdIqMC7mxA514QtIKLxL8ID6Yeqnb8g6JxxVkeEdndtaomzeA
cmVbb1C5roAiy18WwDBu1vNEd2DWdtLD4Kr13/0qVM3aqPQpjAVHC/qiBXHCTXhc
zRbTRMPf8PiouhznublIs7i+4QM9D+/ODyhCTaTfwyheVLua07g7rvGHNkVDFWpO
IJ0nwSWH3K/Ck3RXdIQNaBvAY8pkBu7Yt7eqGP6az8//S27BMx9IGyeana4+sPcc
RBx4fN9Yn5Q3GBEU32mnAlqfR8r4ryyr0JzJ4grB9NChupT6OYj2eDaaQKqr24Z2
eJuplTtqzfxJEqCMFuZRbvY+gl8tK5XuMqnlONtfaF6uSS4Iu2BTxbW/Br8qz4hs
603WWRbfzmlS4DF7uLJxe9owMfroiRnDqudtBOS1FUXNANACWirEc3esU+5+ZiTK
6ldvs/al++98cyXeyr1ZZ2mTyFupzBaQ2IRqwP30OWgG8Kljx1lTWYhqqB8/xaiJ
UXAMsHWuD3RFM0GZbA95heaDThEF3fAhj1PhznmvCrU1FFNOfYki+e3LxTCCExu1
VeSricytC7p5x93lxzaZscAqBEE8UcCsmqXHnaAbB49964QNYAiAsMsY6gf34Zu5
/cfOIA8RfqURB7mp9nn+pQv5Rj92NMLB6nWyqjzEGKD55n9q6qnieo9aE1J6R8OL
UpKzCD+LopGzXgS4iR0F2WEj499A1vfYkCpMm3AigTWEaB1G5YjRTH1H9bDV4Q9v
9unxirWy0QRR2PAeinYJ4MPUoot3hoOgFzoOgL6oZ6bpNJLdWdNQAW/yQaYv/TjB
U4NDN/hDNOIBkAiBG4TOr9nmPyRM51DqLrBSsUjTWfIcjhsm2j20oq4+zhXeInm4
IgTfpegJbiWsObpo9viTIl+MsqLmHKw3/QCNf4Qg+7ZF1CKSAfS94sHGs9JULN+d
C/BtyJkVTFz9ua5EPDX+vlJ4e1+W85PusFt+f0jS+lJlq5bReV7Yn5GWFZ8ZfW8U
zsQxZfCniBwHqNQ3JxrkvwmBcka1RWACk1hFtt1GuJWyspqutvKTVaKiH90s0Erg
rdP1DqT0U9SurqIxrPlWyk2CXRuBFRMq53vMPJf3AQjYJD63wx/To6kpRa02stMS
77W51c32ECLUiJpbq9LxQ6KpsymEu1MP+jvHM01QfghPXftQ117+fhNKDSsY8GlW
KXVCGZgiAs799BjEBSZqYVS6PVLfr8j0GIhblCHsm1aw9k0em/b1s7113y3qBHjp
UtHn1AcqArx7dedvQRfFSLZ3z73cD7aB1Z9fOeOb8U99QgDHe5wJFo0EcmCeIQwj
TXUFdTsM4/5TYABnjWO03lzr6tPdyWAXFJhusMzRhDxMtRxpRQ+76zP+eEwkatC5
qX6aNJhlpzJDHPR70qkW+1AIpvShoNCiqpC/7yJIhBIUEfc8ia/vJhAUXvRZqrI6
i9U30nBFLbdUPoIot5C21pFxiLSl2h/s0xeIEU4JwAHIOa/XWREYOtbg/unEKP2z
+fy4lsEhTCa7jkL7frxCHipw+KPQEqK6eiwAWR+9i5MdLP1nlpcrRZdSUEuXoPyc
lxCbbr/WODxPYow6sE98Su6KQ9PRWP6jaouAjXsRmF1DSlOBJxf/dHZDrZIMJ5YG
uRKnX7/N/7z/tFcdLmDOBSZPmv2TznOafAIkhyYmD0KJZnGXEo8ClvQgC2ClTOXJ
FzKIA+ZIKZR0GZ0pZtG6obtSPZsdla6xSB4TYGyXmiYqRoxWieEzhO6TooxXk2U6
Q7mqX70Pp0AtwWVSuS95LWVsvaFY0yC9WCJXEPeNceMYxj++ptzYCk2y5g4j1yZj
qSav1AxvqhFRqiwdsZNhMv+6ZcWauXTu4anY0ut/CHjhjQmJ0yygL8uHV53JO3Jl
Zl1JKabf/f4vmuFZAG/XhPqB+AQChoWYviQZNEwNznNJafoVgl6jeeoptdstyzXM
Aq3Oqwg/S/Xz4jZPpxl+X3eazBoFe7DAYNHwS3tE4yi7AEnlu6TICoEonxDvfBB7
KTKBM/BwLwwBlox/zg1t/mK55kzv4Spefgz7DKsWKK7WGOtgChQ33aRiCcDyEJr7
74MYJjwTV1VoOqmI8j6qQjBaLsN4MO6/qCP721QEL4Y3Uj3/JimqN+rKOzhabGih
eB9JLMQk/V9GgxB5QiVQr8ku7Duh3Tkhq7jhyHcPZSWfeuLfNASuWDQfTIBVIL0j
K8uU6gtDCBRxI1gwlT9F97G9ypD1jL47X2gUGEcFSARCDYstK0+DG65esO+hzX8i
k9UxNOPvwXHJIFE8w9qHhqNUSkQ9fnjuJCfZj+8MRItg8Qiq3Cjgq2LewQPotisg
lLwl2GFl5+b5uQXZCUDCLfoBkse9aRt6e91EqWnn2WP/jA03P1x8TY8axj4VL69B
FDCAJnQZloHvkLPYAEuDIWTv7vRuMQCfKcATHGiAYjHEy3t1+s1QO/Jt63AjbQgS
7XdBs3EgedRL4mR4rZByGOILkPdqSp8V/QupaV5DXufEL963cVFRsvtRzlYw4laD
XcIQHnwuXp8PTRmreGaHGDVd1LRu8973E5SiltVu6xu/glFeuMB6jw9gHept1k09
zVTJGHF/HjcdcSPreh7Ynrxj+Mu0SSSK4SwyqFHkF9nckKyBc6Z/S8ais0RQeSGv
aKW9K25SHlfsa07lHVdWT/lh15tgCxssWXrmO6hPSvaAkNJQt5SHmRe0YHJ+q2ay
MCUbWgT/R/6O06hPQi48gm+Z20ccYXTlNZaTARGilMYVS1NtU+LLt/+4pSdSbwDI
Z5zZ+QexjNsPZo9d+XMOjSxqXeb/cMWynnxXuiG6W9Lod1Sc0z5+9Ew+S97MaHuq
CjJejNfA0pvvHZZj8D6n8TuZCU3d3lb/Nh3JoU3U8eABdt9oI6cG3OQuYFj5fn2a
dAPNTiloa70708Jv3L55RJ65/pch2lfKbDJg9dVeggoDboi65J68sCEOtGYmjYe8
8fN4ufEHgpkajq6w9JdCzIIZ6Y+KmKrj3jUmLvn+iBuhDxU3Gxvt/OMUkMUyixkf
7QJqqBF4jsTlSanPVgfdRgUJuF0IfDDRnAa8sHAIICbJelGSitLS4IguD/2yo3RG
Oi3Z5hMjaBvMQjVVxhPZQ738tSW3ue9b1RPe20ErJpxN6rHCdV3DjYUWl3dbCpsP
/AE3ZA+Uj7i1QgE4OdbzF9xJkBnox/cAbMd6vh/qRl+uLQM00LR9qZEyKESjyVck
OyKOs4oQ/XoPPcRjytoVt4+U01XoFDczysbAMoYrlhNxhCeB1wd3JxfHHv34jXUp
bL78O72Cg+9t3zMUQG+WKIov64ITTgRBo/gY+E9yuErkHJ30QJ4ch7SvcXsHepJQ
jkoE62St40hIjkJtL007BUGS66yeHFUtj6l0lgqXvYFRuv/G7XgMfImXlWmBNUh3
EN8TuMktdfjczm/i8bo7O8n7lmAu/FtcnbkJvt6UMolBvyQNYNSh9fx9LxboucrB
9Q57B8BtgwSljxVUVq/G7SXzYcKgNo3tkxmU2pL/l5VgrbHPUYPcvBdsXzi6x9rD
GxZgyVRaDQDz8Nd3ToJ1Npwa+5MKoe8e60lee4LoHp28OdNZvSR3FTZEQC8rxMq/
DkESIMFKJ9Pt46apGzaf4H/AC6bLBcl4vak4yj1+03+bjtlefO08Va9pCKnN3yCZ
N3PHPrfo/uC7suqaSyC+U3ujifuzxyxsPBYVbVujPfjFr+PCLNRzuUVfCLEQBlBJ
y5+4ZIjBVO+PYvjPi/9oPneIO0Mjt7QR5whonvYIFDBq72ppLL9GzaD59XJ595ST
kixzQui2VUdTnj6aIiT06fk7uXlpixoyV7H1gJLLEszCnjEjWZ5AwytIx8GA06X/
oYNOXYChDIGxs36H2TwzZi+Dp1+2RQP39WWkbqcVr7YbVlVVdVk/hFEsZGuPl0TM
bEz2r6X2V9ZbOHmV8ZTOC+QpNKtcu99abnipY1gfoQ5LYB7m5NQgxlvps4BJqJJd
TQYYafzHYRr824w8aYZyOF6LxNcRT5l2CQVZQyb5ovVWvLqIgTTcDEdG2ert0OlQ
lfHpBFRoDEgYarp4BD/BwM6RB0tyyxi89xxKeKmlK4cP12SaKTWfNnqn/YbZWcam
Ucj/faXwtqBCCtHIYNIa3WndkIB1/s2ZNvG8vNVUq/4BUoFxxvjE1bdU2Imt7Jm3
2Z52V30NEOmu25dyPfU8rX1xEnGq7KDBlv2XL1OFM+LukxDBFQbONhVTxLtML3C4
f7/ml/B4rSmEu1xzxs/4Wpmt+DPZvj9DGjwe4D5ppo7qO06jgtcNQe2W9C7PW8Fz
wRb+mabblrgIu0DjHThLoLHqsdUW84QPtGZj8ejpc/83S7IZRBuRbEzGNQOa0iPK
wp4+qWBkbImiGOrR/TUQUMD2Z9ZmVheZ7qiJ3Wm6dI5UMo74HjewWia8MIFKO1p9
Oiuet9h2tCQ9VvsfRIUEGf1QE+KMOhxbLSykuooV3JFzl6hhGXqUqeu8l63pXYMF
5stcgRHlxzz+XzmwyqebRLj4JnUc/pX/9Fj+fLq+0j16dfkfnvQPQGWXvpXW5BTj
rSSLBd9bK0E+i/wTQEKg1U0nGwB2ZMhGDat9AKKO6vtQJCR0lGlN+EwGeDRcmfTr
K9GyrTpBsyD6lls2cTt7zDE+40WaXU/xxVxHneJignZHKC4VMI/H3HQiFDY0lmkR
bKSovoZmYtTRow4d9RkKVyFjei0bA6KhbYciQnLByfe8K3cdcs/IKReWqIHYCfZJ
fJq7Qs0ELWmAU4gT1xBkPcwWYdbdqTV2MhmA+bY59vYqC+/c1kNl9W7nWOgha/NY
QmtuFKXf7z33txX1TAsHUfsqNHHKAqI53qKy4FjiuVZ4kfehL/j36CQnZhk/Wq+A
g1YekGucGW8kWo9bYm9faMDC/nSo2jptyau9xzXmnBycQLOYrs9kujQphTCoTBSJ
P/2WWRLgzVnSGNvbxTAyhix0MJH89qeErK7oMJtFY/t7DSMomiFs8RK1m1OQIlDX
BN3DJ/TpngfJ4KCpN6LM5+Vpv1aYL0K8ghskr4Q2hKKlHH5Jo+8pn4w8sLKnn1CH
pm+cfOQiQL3snhT236ZkKbgekIU6eNiISgKObBN5cEDa6kfpKx81lPSCP3jI/9g+
rLtFKq1pieskYSOFoPM9gQJ8zB+RIFQnOKVI7QOPs7rsf5B9P4/xCF9wzuBl0s45
BhDB+CQR4xQVX605y+UOX2zx/e1jMG/mKvIjQdKHOC454HfA/H4RuKVgxR7PMY8G
PRrPvP2LoRAw1kzDmEZPtSb7xbhSNcppGWIblHpHGZmcfwOyCA3HYSsBuyqbZ2J1
tfR7cKo859wqAHfyk3f9QZ9+dL5kGfEadNvyhODNX/mJEluB0o6TPUZicNUEQYgO
ahaj6a5a3l4V7dbTOHVXkllJDZxe8rLqneWXUlh0rYFYKFxoe1WU8OmxGGpcwO+8
5YIyJnUEAojsi9j2NgkAPcdbU/qlxyC+hy/rYuyBqTvlgrZ8FYl6npyXR8VlRYn4
uVpCNTTzGz906yNV2Fgqb4Z+voUa/US8LVMwWr7+HsY9AbLh7w1c0eNw9Zts/vYY
Vw6Z1T4LifwMYI6wa3hpgYN9KJeb+dNyUFERDTg5Oh3UPxGpnikX+iq238FkZREH
/2HxvDrG1VGUpuCHkpTwoXaejEw2MBwp3VSJm3SOIL96esPPgq5VESLT5V1sZL2G
bjv8ZpESsi0am1l0oE4+DTYXQZVkHjwPn96IsVS+HjkJLOxnc1IKMBRop+CtanqV
u/mwcMB/S9Bz6vboa+GKU2uAGX7HJPA6SFixD3Z2lQO2aiS8oT4u0Vi3Ss8qRALe
7Blhtz6+xnmP8HQIfG91sd0Vx5i0mYQfWfUWhMbedC0EHV1Rf564ZImEuDcC3Acp
t01QyW4vuHoBFwkEWWIIs8JMPFKtepeWDZFYll7/tjEY+LKDAJHMmoIaZ2ApzYYN
GKiMMzmnDpdJeviUtoyxq4x5cOaTw7dK7xPd6PS6jfzBWzZcEdtxrivCrXOlJ7XD
knWANJ6VzA3kRA6ef75dCB/vaOj48UMMa4Bjo4zsrrDTE9WKhtByq20UyL7MjDPF
IhUT8A7jz1FC0H3/YCwD1CVMLlSTvGZpjBnw4V1NMh780/oLHma9NjrzTi439DzF
/0cGTTqdZusTej1t+8Ook4e6kyRmnSP1N/q2tb5ukaiK/EaWXOsEQbRi8YmvqlSo
E66aE8jVcTWRosCok1/kdmWQQyhBXO7/6+pjEXY8sBxt7acXdUc2yHVvDEObT9Nj
AZPptwqo9jVnXE06ETx7LqG6XwijxZX+Wwx7eW1Ppy+tTyEycUTo4qawmLpdhhrk
ckf5P3Ns+DSPsRNOwGGbp8EBYIRL5KHfBSp0LUfbQEEof12DdRy1joDOVS0y9VPn
2yJWUNc70Wx1YxkZ5BellMGSFd08OoPZB0cHtTl53NUX1Uj3Ak2zVVb/pxwpb8ZX
Ha5dA7pgLLPpS5grsqF4ebJlIwRUGi2+O2Y1+vLc5BFh6jmw81wprVEMQcF70l/j
wh2Bie3v+KUqLVVsDHW4RM4H/t429NUXHv1EXSmJP1bJ71v+5+IPNABvNQ8wrKmv
FOywra1Ct/nwoW9dtAmKIhkKYNdApJYlhP9fAmfBVf4qcfsSlywvQXaMErwSGWcA
BzzUTClsZHjgmIUakYYozlfCY7PnvNzqOwIHyUSoyESw+2t67wUbJUO5ltX3ceLD
OYIqftqvd4cD0lAtejRe8kxr1JRwwrJWHCpCxULGJQNLA05F4WTaREnX1/jUFcFJ
bwrkoutCBYpvGpGEbYwoAKLTY5OZyUCeWBsN/28+FeA0arfJ174ywtlF4DENDhlR
Zcr6Rh8EeTf4VIonNecO847wgkogWDP8HCsXP+Ji7dBRj7QcTHmKiLcJD4DdIfxu
iD+X31dwn2bIrFkvCEYKw3dOOGduOEcMBcMu/VT6TVnIzWx9jfXv/C/GT+gVTWT7
tnoaEWf3P9OwhfES3Is9qHoUMi+ZPB5Ku2C7NkB3ImEMgvvCR32azIeTSQVznfzC
2U6bc9ZrJ75aDkDzekXxyGJoL1/bVpIMiSQAOrgcjslSzPyuQ1Z7TDIkRUYMwTbJ
qRa5XdnHbdx50j5Z1PgB+5yOfJWzunbxrk+K1t0P3+E/8CNsSR5Up0QRbcD14m85
6Wn9UHfpivXQtUt1yZtQ91KpexxB/Lw6W7uq7yHQGZewCBmQB2LDiPRYqzCg9Jjk
AYrhjOwD0EmMpT4BxWbejxNfVIlS5aCWdG94jKLuVy2Cucyg1CaYkLP92vxWJ8cO
RoKQkcb/RHppKni2hEBRxE7IWWGdiSWRcPXkoJxEtEBKD7yPilcQtSnNcU6zLBNX
cJZIk4ha4+hnrwZhWc17fUBp9PD7eEVlH9S3r+HMyExs8z/3ihWgZYe1UonDUOhP
ipbZejBIBVUtPmZdwD4YogJy1Yzg/4qJD8mj6J9SKBtpIRCTlsEkOY9hip4rZFfF
1eSTft/+nTujCG/mFH+mS6GRCn0OR3GPOwdHIGoZdxVeWVss7SruKiI0xwZOfAQM
f2OIopE+2cFQEKtpdkc6a4Cmw5A80mq7L3hV5bKqS3/UIoaVCATuMwiVQY8EFupS
Fvwdx86uZ2Nd46QD2zh9zkiEWfHnvpcJ4iWWw5n8BGPqshXhmXds0VzDcga0FuP3
zO6fiJIisWJI52qI29wX8KHa8ZJVri2bAbt36fzLDc3tn92Yh1VFcgQhO1+hxef7
2VLBIWrcDA/r8LugfnPD9uyQd4ag4dS9ryvJjKWyse3tQBaX449Fn4rVdNL/RnJA
FZqRKWfJXZbOMmoFtaZ79jn97FQjH9q3Gr8OWsv3qkjVpsAJBbzzMclxFMohIPHS
4tKiEtgxEUq0MGoR/YlKELg0HW7WRV2RarCh6+2cbMnd3GeRko6766wUfxn+y8Jh
UWhLwi2YZ3LkpRWfCzs0/MdVdXFvRd6whtCC5Vyy4yjSyvE5uwebFXM4+nk81/ha
LwzP3GtAduEn/2EUYOF55wHsN0+GKNEGlo4Haa4T/fjq4AQGpxVpm+iSbHf1n2A+
YXiiOVKc3QSe7drW/bzAUfyLFMGkaVegZ3amHrb2T3vbsXD/7h5KA9ezb6a5pk9n
ZAOOuHR0sITgW0IQX5TJeMaM5ZwzQCPo1pkt3XnsHqGfF5fYa1oO3q49Hnd8PhEo
YJ0dpU+jWGcJ2hxNjeyE92iIGwkrjd2Z6T19CjB42kboTrp/IOvmD+frejymW9bW
0qOQpVZBYR3RjypXTRlgzfjuNto8dchFGpAJVRX7Wa+U9YytITUNvCTmK7ykZTcf
+ry41WmcahyIj+Q9Q4xV91NuotVepz0jttCGLJTUfmehEaaM1I8hJfngNCvs2zd0
mWnGTjAUsdr2RC3eSWIer5C/KrU2M5XuFoCwVc6C/fr9lDi6vkNJBnTI+nC5GrZX
ofIdQeo95YCG4jAtN3zcQu+UvBDTweExctSxE72NKhWb7CIfTitrR7HwhWZu/FjH
35YdwsUxOw4pLxgI8mbAeQLs8Np+3mdBtYK+w2xwu29OrBAvZGRz7z7jEUel5Kof
++qcqAuDqW2ZJvJKOGKadulY5Ju6i/QRc/nERouPPj2xcQyQOyGZgxgs5vYQabRM
El2hte7p/FmtlLY+6U87Has4m+Q9YhE6W+DOZiBpmHlPJemaWUeSAcJWi3/sikZ5
Hu/YGbxxUbqT8/RVAj4Z6oJrYsvD1MGDgQT5IFXGc6bJyPcvCO3graNImJxAjiqC
dByAUMS+/FCAqym6Egt4VQqybTdY1iJD5PNvlGI/IvZ8iaLteQkhuPWbsDclEHAP
ZESA3fZwDs0z2njiRPjP48Q+dLDo0LN1GiI7+W76kq8XPMCub1qAOYL0iWzorhtN
0OR+Ye7pziRL/8ge6CeLBMkMen4e0lOC5lRrp7/R40AcOjPYfUgAsy+l2E0qGGI/
ASQuE/LEwW9yS9S+Qo14WTUcNejZnIsVU/ixHiiQA/Cx0+/DulA6StvJbUIEDUnL
D2JG0LNe+KsD6p+f1vGmBgxbzQvcC4LOKxFIOAeYuJW8kZcJdpluFOdl/L/QCBfK
ctDJnu0EsF22E5qkS82xSeLPpqEMEbvvVfZ/SPHAIvLXdftDX/B9u2ZtOmfLHvNj
c0ZI80y6bJHvowsvZK+sGE1LShtWXynlY310ir3defuBRt9ktjUB01JroCAFQ5X5
41ayA2TBZfuwW2swB5Q8uXGevXJHoYqLS/pg1WMhrUqp9p2hV7+gDGf2tN0HNheC
tLix+4mZSBf0YmLAa0m1dW0342TwJ04jsDWyrCsjO3iD1u2FK+fOcT+qXVqAVBUh
5UB9bQZF5rwEiipFySOj4Zy9pH3137guOozZ835ON4BfRiHcWAT+MlNUtduTgHkj
mrKCTTjIJtkk6vY56xmDlAmQg6e7iBnwGcztnj2QgPcNVlPWUH6SY2EkFiHPAfV/
25wrEf1w7baxi2okQSXkjWUyZ1tPmbG+SjyHbnmij2bU8DVJHBuItxBFqFBD+nFa
ISXUYK20tpQfEca5r8wyr97vF29SdlOx3tNb/ABvWo8ca1v2WN+GIdLexHzUCN1l
vCvOjL/SnUhFd4/15wEcS7o5xsULx0Mpt4/bpfzSGgUOlLSVcjoP6aRRclC6otP/
MNnmFUhvjGK6d6/iYvMgF38pdat/F31+w9By7w3HmleU1ng3PXlcCzsONMrnvXy7
aVt6k+hqnOPEgmtoUrpG91qUaz1FPbEkt2F1s5iWRP/YHyxS+dlyQT/bEqRIXkfq
ylTmZolN/3MwfHpU3qGwfB9lfelC+fiDug4+MV5VWeAa0p/PXilxHfkCbGECr9P/
hnAx2QpQ1z+fofBJEhZp/nbJjbkz29DsQzFKIDZil80DllXZ8zPgY5FHeP+I1sO2
kjd8a/gUNPbDAIPkgMUtUsLpoQBLQPnkr8V3WdDWHBU+BlR6+0LqAOLGikxz2cOZ
Sm60mj36rXSCmX2OdqTlSfyHG9yWhefrWW58mh/Kc3tYPvuprkjXeqSzUTs3n8In
+0Pv1ZMjIeuSQZJViMI0tg31gSdI3/KCCR0harnsyO48fitE62J/fzn35CPbqydZ
XBBTzjJ/AzUVsxXO0Lwg1Xp4ta1CcKYuYscThU+v/oQMzIaj1zqJ8fzdMjsScXWm
BgwUXLB+UXg6ZI7Cty+pOYgQYVD39byGOMb18IoWdAPJwGiaVzaLxMtZVGs0ynbn
4ZHmDJo67u9h80SqlelVNjCpVVbOzYjm3yb4oAqPxdWRVvoN75Jm9eF9ZOvnZ0NQ
2Gv9nvqop0SL2VaTfpNT77FVbBxUPHmtgPzfDO8YMWvywrXWM9AhYQzrNszDS8Oq
W7mXYgSm0kCLJdnDBOwMT3csGIMtMu3JKqrvHIOfoDBBM73Eu+/A0fUIy69+W5q/
vef8d2T+mKGPQAWDCjVe64EiWoU85IdnG3q2NW8DRsNPLg0w5LtnrkVbhbb7EPeO
hYZnrATlC3T1J9um/oqQTmzHckPh3Sc18eLw0v1GdCtBNxQV1L+I5c7Xz9oT/nYG
72SgP4zP9+a3zExbVdglwYI3NEelRaEnatw61sylOAisdvG+dJ6Xs23JBkK1HHo5
/uzttxSmMmuX57iuCakeLiPPFSNcMW8BFbPXXds23gZs5zTg4MP5fQSm5a0zB1xU
BfXwyL1CM0SKvY+fcC6kC5Bds3PrhiVSrCpPZE3eUTDLGGSGiCwt05/EDox5ZeO7
C7xVOvaPcrMVUiiRFZsg+cnlLh+uors5GL9zoWxTjP84nb2AIlvIyYfouJupad8j
73CjGQN5sQ4MZVANo3xdM4dE0gkiKZiSAt8X7X3QCqkDn+IIOExrE13egzTpfjDG
GKpQLbbdhM6V+DOgqci7J9aR9xHQ3Egvdb2kf6nB6Bd9jcNax6M0jt0LaXuExMTv
JldK6VmVeREeEuaNRZ7ydyKXmeuxzj1gDWjlx3DJPfXzZ+UDiHOFZ4fMTQ+XRFc/
fJffGoQgi2jQpoLUqTtqUBIQOq2sKA43b6mUTnp19dYXPzL1YbjJmLuIzEuKZG7x
xiVCQh2zyMaVKuACi4tLvldqm/3Qe382eDtenK0D9IMp4TaSnmWUeUvjHaRSkVd7
JBb4Ut0qi1VG8DpvnnXMDuGHUR9fBw08J2GAdpRHuqmGeZg38m8rY4PwlbjxDghd
aj5+Xy7t9IFoBiVowYq4EIAd7bnJFQjuLGqTmE6dJBkhrnAtSdhDJGs+wa7V1dKN
eA9/srBiwa9N/CDDpu6+vLShPtgS/GjrPdS4Wfz/DHugtv6YxEmMLt+JqaXlbion
1FYk97XrSV0F41py3rN6xEwVqF84Z+rLAm7wpxZiQLYMVfm3HLO+NRp7HjPzTfKt
cLSQqBdxz1ODNiJNVaLUm9wKAJX/omvzHiyN2yY63F6X7mY+wtLLzlSkhA8f++OU
DNBVEmXe617WSlcxOs3ab2z8rdykZHKI7qigCOjeSRc5Aj76NmGaanJKDUDdN2O/
HEhyL4sSrZsc6643yQg1Cxa4QoPJoRizVUzcPEamS5wEyvDDWWWduihJ/LaSXIGD
Kdb4faNrVHWE8VdrF9yeg2bER2qRxFj2XQnpelaENYyLTK3NUps1iy3YtCK1gw3g
dEdigA62zmJJ/9bQEHw3SzjMOEsF+8aoB9eNq5cOJmuWb1kGuIleEhQNylAPd0+M
Yq/SNr+VDAd8QLFkKqYi0W/4+25yRIM4PxdgtNhO8jAvysy3lOqMp8J11f2I72Kp
tOauOYzLUQWEMAeRP8JFkPILEabr3+0Z4CpzKtBC7RPfPHDlEN9chRUtJEj+4vQO
NjyQlGE8yy1z3Voi+ZzI9QugikBFy6LTCYrDbd+pLpx1GWNmU3jD4NDYhKJs0dUH
9kf69615Xtbeg6z+ApdW7+WIFICWx6rmGSMks65bZwepEQ8Omv4KWnkaiRuV6NXJ
pcrLcdR4w61EFIhWc4ObrBnvXsVSWbVf/2UjR4WU5MwbYu/fvkR5Dnp1k9Ojo8wO
46ehMvzzD4nAqMc8b3YOS0jipxkvl90CMxtB6t/N7A2eowZcueB10FRzNAD4IAwz
n2Vz1JGPkXQHhEoZy5S7DD9H0jnQksy2gYZjHNZdFK2Oka9rbCPOHhzwDwhSFWfr
ygUvecAdpXEMeg1ZxvTdHg19EovQQU7LH/Yuink2CMxkVF0YmSJjDAEjfnZ9IYNj
6PU2REduSUyLaqADi6GjnSRLSVVPjHIwIPg9zXQBAs6p18JKuIlg4dcMbboDnhL8
HRE1Iiwu3804aXjd2ieOUKqmkvkaJwrHqxqJbwvXs1yNa+LZepqWAIKVTtzTfHbW
YvzPrPuHNI6avodlbcvzIZH98x92EntIQAloCYZx9raJlfnSVB96IkiQg0UbfmTH
rt4ojSn7QVYXtfEiSNx4SeHUzuAEDIoF5jd4PSFnXWgI0MEfeKtEuS6sPFTA8cuO
tVKHXy0Fn0pzFcTX5an7zOfX0qyY/0V3ca/dstHSt8Tyth1gY/FE+8hqqGE5oHCb
KSwEorznWDUYTpl22+YTWdqk6jYewSmB7Yg7ysHniR9gvDPClMWj91Ouj5IFazzd
OQI1NxvuSxeAHeaqNuXCzsWEXJ5+rHGAndxtfL2fcsgjlTu+kxNlbVyMGR6SifR5
68qzzpyqRnGo004cD3HTTB3jvnH7NEjj5j5ipuw+G5Qb6Kn9hW8a6vj1uN0TR4px
aezMSp7L6EUFPZLSdLpZlnugOnq4El8IL3HwWnE3WjZFATkyX3bzLHO8bgmhbSjS
kZZiuGV2SL6/kE5ft+fDu+SejcmD3q2qf7aZC7KCKaG7A7YAC5eZBvGvRSKSgrEx
+lqPcjRaO9xGl0UV9YEP/2TfIffIgEHiYkckHoYCtD+4fadRkxEPD04bwhbNes5G
HDO2TubKB3I5aTti2VFwNKjov7YkxLH2+aOqnwanzYe2AAdlAGKQgLrLRxowC/3/
3dXAkTUMSpOg8XFjBDb1UYHMuHYJ3ZSn/Pzx8NqLfQpMDU6naedlw1AwIFFyoxO9
qNbhwI8UFogGcIZoipJshCrKfJv3/4/sjDPj2o54uRNklGwk3i/xN3estIDz7EHk
zKwBbvo1VTLMZjeWAke6iZG/JZuTU2fUEDoAPYOOGz5GWEW/3AhguBuPRMu/kT+o
brBjBd8x7AbMQ77ALBeqvAOM9GfddhsCdmrwX3fPafW851rYRARDPYGMZ0KuYbqm
Y3igvpYFG8iMBed4P4NNxHUsWy03S2fdHtCPo6WeSM9PUr+19yjUlWsJ08/sBkxp
Qvw1JqwN0HSf0PaXnetfXnHDcn48UcCSQaGXnBt8vkh3LJqiiik1PvZBVTVXWeDT
bdFBaFgAW0EZ/bsP3PARc3rdr1E22dGQFBCYs/jXiN83gk40RcbMBeAlAubbcPCa
GCrG9R/M4HUO3Mc1zSBEPiftjKUcaW38Js6dFujUliuWoKGIE2/gNFsmTGpCzSPg
VcvLSXQ4chDe2wybprWvnu3fSP3ubhYbHO7BjPAkFcGH4OnPjF8ETKriJIR3LE7s
a/LyUO3cCFZlb8CWpwGT3NI033kIOM2uwxAhyVFJv33hhIPHjTmZbjS0T8086Ys8
Tvl0ZTxZxc9Q6DxclucrORb/ZGVmnwV83Nn1CWYynSM3K5DMCqmGwd8q7umIBajn
J9K5Ub/bcCgqCiqoJRdf6DHeayarmDSu3PAunx53lFtRp18lSep3sodYxZgymBV0
bHziWx4EW/5P2czzjZHfHYyDkKJ20iMa60NRIiVkv4KrqzbQBnbOVzkY8JlFJYtX
9p3BbV0UKMxC3BJtcZvKTpz9syTicG61X9ST9Yy3Q5M35e+Xdi+vRHb9fzyind5a
eE2GQlAatwwNKsY3V9fIuTqAFDqoSJhRE73mMiMd9cf5BHCFsFZ8aSN129mf1bwD
wGfkNSy6T6EK/PJl1Ip8Gb0B+TEu+oTHsWGqDVvuBRMFA5V5ClauJkriwpN6gb6J
8/pEVsR9TqztK5TbCVVp68ji9yu7vXYItlUl0KllyohXNmdRhG/4voqG38CtDAmN
q8045lBnW1sS8jvZ3gTMw+Sferv/142Zo8M2CIUG7EehZkrnL3AmRCD9ihB1RnCY
6Rp4C4aPmNMoY1lvay8NL5BlSiTxC84udgUYag6RQlwe9UZI5nuJcDZrAHExg4Rn
o2Qd5ZuBvwS41sGi6D3u5uDZqCNs+NkhhZH1mc/9rBtwgR/aDnew2/7KL0VML3tI
fi7yuK5Vt0+CyYcM3anZdPmA4FJaf8GjLeug5h3f9H/7PNjT5GQdTPHdKMYD8fH8
4hYSO+zyAfKp5mJwarnMZAH6lkkfWDzoe1RAnZ+iNNmvumauCFO4a8QlHEBSVwvF
XvQjexQ9Wuyy9381XdZcMR0SUVfuQIIEbjzYv/CGe/5OngctUjsdk07prZJraOQN
8GA+Hs6ECYfdoK/CuTnzRisSZbv5KKJYCJz3NkNgrn3pYf7fYmzntYK4ExdAwln4
w58Vx9Nk9z8eSa1D5SaIp+a9JYMf/FF3vkVq/ljq59lWAEdELCleBDBxrIp6EQl3
2XFQYJqLUGndOOWYkT7GLs02cja/59aEUm81KYlp9KCPb60NCHp3gVJQCu7/eyjI
zmBkf4xAlDTew326vxNvDInkvJ9GMjzSOmX5Jk8A3Oopgw0TK/5xNSlsORxHOO+7
LkXJ4WXR0B8Mp+L2dHkahXrwdOgJ4HBNts/0t8aYNk3S32nA7M947wscVRGI6G5w
zSyWRT/CLwZpElwPfm7k0rPd9Lm2KYi15cOQnmCzF9f2yE9Uz/FcyprzBZXom0B4
6cX1HSZGgp9GZ6iyaI58iwoSNgfHLf39N/WUCGLJ71z3GHxWQDXOGec1g/bja+aO
79zJY0kVUHvQg2xHKxAbLvFzOSEiO3/O5bTGn9bc8CzLLAhwg5Rod691T2ZslZf8
bfBz617KQhC+59KlWxEtT4DpJnJL2XPAg480YdVI2WuAxao5BvRyCcmv0oQWg/ti
agpofvOfX72FFBkT6F+V8LJeeRoPhnIP83UpEB7CV0IFb3H5cgcay/ZyZ1/zLO0K
4KHZYkSSrLz6OwKqlG7JsKzAX5GcXq9fGumD/kM/EnnsMBUYHs3ThF+RwVaCkY0C
DnYbOb/XbuR6XpwiQNww+HEZHeqDl1kKZ4GpL6HGTwzda3+q0lk8rOewazBoiBDs
F6bXjfIaT0nDbNhp1r7Asw1KbkSBxR3k8/puDeKcpECDOcyBJJqrU6S7wfdS1WVj
9+YpOi2+8qWTeSpR2YZH6mv5CUXLSiCsBoCxJWSTvlV+Bd+DasH6vhL8UioY3goY
Df0OV/lXWNKtXS6Nx8b8qwJbgWC3AuAAZ75Fkm63xm43lSYoeI8YRgc6ytMe3iC2
9W5v4Djc6/W6DpajxNuarQNHpkqnfambta7j+o4hr0pGyc9WhrfcNz3+mseeDSr3
grrZx4+gb1mX0vPzhNJKcqqV0AfhPM7P6jsjgJFsfAvOXiojo7nKwIglZa/Rn4F4
Y88lNN5s0ndiB1LX6y0bCsvdgQiOtMfbwRyKhhiz6ZHXL8p+xMABodH30n2WXszh
4LUzOJjp3WkjLV4ncxGhEHNzEwk2OZZ6YB+x61PSVMbo8yAvHKyBQzZWkXVVZJsK
dzZClxdKBdYlwxZoFux6so/DYUrcpGTGJy82LDtkOoDj3uNq3TeP3i05kSVeImt7
DXr75RKuuOC4gtu+3zZ72V9rkO9pzLABz5vrAvNgbaTZjuq/ThXiHi7ZahVcVu8g
T8Di8Wsa+X/MwKSdEJlkXyr5ELKmND3yDrIflcLQA3A+R1Ka3CksR2FxB2FuU3/h
VHqCEQFZsb6YVqBt2JMooOyWWEuS/djt1r0dtAIioAIRg/IYNyEdJm5QRypNOaoN
La4Y6mfy0Ht3WX+/6LcyGkL+HQcMuZYeRmgiIfDq/NRW5KSsv3Qb31Uvhzat9W8L
sIYZRDFqyBZzzVWPn2G6kZWicpKN4Jm79MSiYDmE+TVtXbEWTxvrM69J2nPqkGkj
Uao883QCUCAbboE6kwK9XtogbgyKuS+ux3eWI0MM8vuSy7M2xl8jVyKQLcb82Igo
4pNN6SkT3DZb0nkQe7RxSMi2u2CiADxQg7IcDbZ+ktpyN9nbqccw0nAgrKI0SSAu
nHxb6bK6WpFnUtz1+NJgHIQ0+hj+mZ9SkMzPPmJZlmplgwBHXORA7w+T956wnglV
fAAvT3JrR0VS3agOhFBi7bbVhIhId7WhAWj/cFCwmECSQoM6zKwRqGfprtUciQOT
MP9lCSkFSCL8d6mYa/egK3+OURQOUX6fqSI13hkBAI3j27BVGNuFjdRccngllXE9
23nSKayZXz3jqPoROrtvZt9NiPuTVx25vhT5Ct+yCJjVTY5SgiTJrBX8Ulj/2LS/
VHiJTnkD7iVmwRy/b+U/aa1uRTDnNKDdEDPH0scncLPhRTjbIY4dEj+uSHTSLt/7
URC+PreeDL/Aqw6IK9sSWgIdfRhCm2FCOMjmeLtAM7Z13WcjIwraOezwwWH40tY2
5kLnRrmExbmoO6AwWvwtIMHHJOI+I8xvTSk3ogtfVkSg9dkootiOmycrzL83+hvd
tmju/DvgvyET2lW2yLrjullogmOn4XJ6j3gEchywXCp978ryI9BztXUg4F5mcybq
VwzLKlrnF4XMwm8WxRM8bTy9VPlO0pOhQpp4tQQK1BjoeuW0Umim2vcD6OthAcH0
tNlj4mDT4mujKt0r6a89PmsTcoZXnaThrwcg8WYW8ppvtg6C/ygzoMe0HfCdIpEo
U+RnY2LjUSSqq3aEYoPvCu0hDjLVjLhZ358lzNBEluECjWgp7N/QvtIO0olcaO5V
63DSFYeDN3ZSD3eVbMz6EIHD8og8sThk8yW2eHSNFffEtUKvG+qQhOfB7Jhp8YA+
hYkd/Gg8kQZjs3GQq56M1L9AR0GBSbXlneZL081XBB4MEeTaeyDA5WCduqswjvDs
7oYfELIsH8FLFVF43TSauc0qUcdSqkefdzrHqOEmX397kqOTIURT6sFy7UJ4zVho
WcBqshjuHQb7U3FvjUqC+bZuM2e3JE0IkSkTn5yTPJqy6swMn0sFMUSGmRuk7eyO
9WKMLwslv2+GQg9rRR+wxtzCotcGzVRpKE6uor0BmZLmbY/6DZqjN2xOgik9CfT+
CK7JclUotiCDMxyGTl0+n19sv9LzLtpQ/IZkGoVCszVx64haKl7i4ikHMCAeZ/gv
7bOSPgtmUj+Es44jL+mLLFBy0/oUK/4Bcl0MP1YLC3vPxITQZ1vjO+HF9HycFlK9
zd4FzB6hcwncRGxTSPGvODSsKYENKrYYZj23k7avX7MA+DwLlkhSjiPgRhIoJr7g
BXAqBixS0WIdrfm/piGOieoD/TksLqdoZ0NwVWkLlJEvdSAm+kaF1QxWx6cIOgNo
ixTVFTEmiA647pQTOd0ry0sjBKe5U3qXLVkHKoqI89T598k7/AJw7J/mgcnhF4Lz
sGrzwbvU+j2xFrLvd1vwRVbGKNviXJVd+bEQqoptaziQkBKuaIGJo9+lV7KQnSSl
lEJS0sqIPh7wO4w0QUd6YXDGsKtPhOcUeNWEu9TbonCMiXpoz1EzCkh6sAIxRhE7
z1BXMSVBZ8Qt80v7EY0V38q/yOVCyp0F5A8ysWWuizfs4QUX++QW5ejUjHZLuyqF
4rxHdEHtyeqkmMf/ytZTxc96pSm7XAjeDgRmXJtd+h4TE0RjEk5x4D7FhvKLATDh
rXl0YUB6DKRCdlzZGumA+lJG4fi7lhIXdbEaJxrQ43jMLNaAZrWog4flBc0xjeMd
5tE6ecWw+Z6bKA2kj4yCdhRkiw9rHzuRHuBEVgVPTqd8d36Zd3EQoMBcE/CBQ5AS
ixFRjnOFTWWoWeumj3flQdh0+iFKXST7avgTuy7Bp/y3FHx6jZyqjMgQ/psa4uA4
GcEvhS0Zs56Uyx6Cq7wl5uDsXnX7nEOQz/tpIQGUZAuLBB5xdHVMAS0ixcIrtskn
TPpXabu75tprcW/Bm7O21b4s/fyz6YeO8LPxuZPfdi4RvxtiIZ427O7x8Dl438xm
WUp8Hwv/zdlyHlInVjDwOfBocfKXFiOVR40tuDZlabDrQuI2pNoWijJiDrkAl2QT
LDa+JX+XdgEoClObpap42YdWvD5TAoTXJu0VWKZP+ik54gss2Ak2CXwd6MP6Lj3o
SfLBTT3b7bQB4W538NmRcDlFK2wawiBj57U4ARHvIzI57fLwXgTuKfFkzs6RINfd
UusSRRVT6fIKGgDhj8Cv6NBqMqgwjcKSLIwn25QYCVCO1BwBo6pIGVMLDHqONt7I
5pMYKANQd1eyr5K70XpDWCzP3dQa9JzdKWs/M4apTxksHRv40KZhDBGIZjzvGGm/
PfqPY/OOHJpPI5YtKq817tiR9Ra1k5aboqtpN979uablfNNXLaaO+xjdnsNIwh8a
3+9WwgIhgDI0fdIsjWUZmXANnlCcp6zvJLiVMleoTvVl9fxOjtX/km4MTHaULI1u
J4SkxCx/mk22eOaZi0M0EPINxGSsqhK4vj8EJVtXxKa4SmTH6SGSOg0xpEmuXDuq
H1hX1hzoFvcBWjIQErJ7ucoB2IGk025olBKn0Y/3/Hc5lnYYv7lfT1kZKi4wpms6
6jTRrnZuHfhXW7HeAysKFUC+yI4DO0rMBE5l9XxXmVuVhmz3Y89G3sWCm4ccqeKN
5wlLeyZjO6rbIJcINacJmnuXAwdIUfT8fK1ntLs8Rs6NNZUBJD8+vO3/PwZKcFwH
Xhwhzn9vfjNrO0ojFker+uxVcq8w7zrhvi3GCxEIA45C6aWyhoc+SC3i2kgd2M/U
FsSH7weUhe6JE4Er1pyk5c40ft/cMRryxs+JmuxGEvFC6uH8IyP6vQeQ4vLywZ6W
cBCKHFU9hGdbebITEeecMmjIgzibpUFPN+NysZhaJknveyGHOSVde4IUVKYWwInV
719gbEbsfjHOHcfIgQzt4PCFSo+cT7zToghszT6701QpztvaMp4EmyDNdQNKGNtP
NyDK70kLQ2Ym2iC4z4NeGlFFdy6AKxh1pRwy2/bt34al1vgb/tbxFCOyA2ddhuJ/
0hnBd81m2+7ZLPkBvE7h4fAVzoj2OzYmIOozTlZoXc22SSS/4OLzAfxJEUeBD0lV
cXuKxJweU7STtJvOQHnuiHxLzyi5GmNZrIEwAb/EAey2eY2b6g2c1fF2RAfUcn14
oaPIm2jIQzFF36WDe5vqAwK7ZLWNq6BBLx1XOCF4Q4k+dJ2DC3cjb50UAJEXuFxX
R6WAUG8O6P7uoah77J/x8JZ1yBdc7VGLYqCHbvcBea9EXtAbWpx89GxDPAMyZc7j
s3IoCgDz4FF0XnXgY4RTx1iU1UHLBiy2whUj79N8BiO+mb/7VYNM8notoramETuL
Y7AaSCNT9JL/nv0SWK5r9eYWnLFpAJYIJW3GxnV8jyrzveGkChvvo4IvZRc8DQXl
DZ0dNrqhwSaYpd3S5ozShsPSgMW9EawEY0rKw3SdT59Y+DDPavOA3RMUCfaIB/8x
PcZE9Z8t9iapgaIEMQ+JBWvV5Nfe1lAxBjACOr9p7cuNCLEj6VzKHcErcn0GU1zE
cQLNfq7g4amzaOYg8JWmZUWwfYUqOjUj9H3nWyF1QvYL7QfUA5AQUE8QDRicCkcs
JM5Q2rhIfxkrzQTAg+0DF5j+Vl7plehAvCS+dKtw7hcc9eloZUGTU69Auuw7r/Gp
f1bRdQG3GYnjl2+zIwUd7oRjUV83gBSojr4YVgTBuoq3SrHBeNn6xZXzlasp2lVF
hoU4+1dPKxeSsZ/wcq60kptWtA0x4OpUpXhZo9QDdoQJ1+k1mhvocx5AiR/wa0lC
xCjUzaH7jggU5FeGgjmnA9bnVDdroLhxFkDNXqa7+s9DvgmtOTjA+iby0J7dh+UE
S8IIJolkEo1+lKsTqopRJ6P2rkwbl1lSIBfwL8OFQzo9MRpVVCcapOSngbdfp+Wk
zQXTni+xYimvy8rA9G/3ZKg5lnWhXjvN7xaRoPjQvF37VSZsRlahcHJShxHWEjri
+7TGVjfOjZPXFkCvNdpCLH/c4nknZevHw0CbmYYzg0ZOaptbjuuim4DScnuBx55F
iSWAUkZzfQjtFih18D6UcPjIh7muSU6wLF4LuLCWqpQlJeHaGdCqy7zEOLealnoI
v4HLwbxfv+vh6/KPLSjbPt99mhA0DCfeFmIHHHKSXN0HLX5cfVXvnThcr2cch/Dt
FboI4+/yqe4hHMtDdm9AIEgAiW2AkWuhaBjntQNrVqT7f5al+hk7v2lXJyZ8fdmo
aTGqH1RPbDZeaAg5AqUcorxiuySlSHV4yFNbAjJMieK4kmssM1XUVJuf1ZSEPer3
9+QJl0zz2uAZM1GTRWDFKqiKN/yrxAI0hQO3o2QMBdT/RBcWEP0GL/HhL6xuGdM3
OiKIg5NJX1JW1LBB6YIqxMXU/1WKxv1QizNLNNwOczp/HZZ1Hb0W/S4wOJrrgeDB
LZdpYRXwR3u4UxfJufMxk3Nx5CKUkwDCId/WrW1Zpe7nYJAVCdNK7g03u3bG+mTe
MYBogBAPV12VcBmMWAzO5zDkmO+max76NjB6hg6XnbVY+rpA54Q3rXzKB7JRTede
guPSlHgTYt3tEGhid10JfGrX85xeZn46JVDV7l9+Cl9itFKAAhop918JksM7+NPf
bBGBDpX+Xw+PWkiAZjuHjdXz15xqa+h/3iIJkwcdVh0sGcczkIL2b+HuA6cTaGdl
FVimtdm5dZeXVAJauTTmZkJECIXXMd0XWxiEoSJGC9g7V/5GygC52N8KR6u9EPhy
5nF835osmQvkajk+nlfLvqe3pdtmNVNctIwpaqHjxLI3DTRgBF59oF4hRTG5n6io
8SAGHT1X7WecI55Mb+0YXJmEFe/hEFxZUfAjTY5QiLqWgVAA2GxOcW0698xWkGQc
0PBuD1B4WCXorfGvLu5xZFTAUbWamdfGUPA6o6wrN7UGpgjumlN0bUUV27Hn8bJL
gwKLbIl4u7sWd+nEcFUwvj6yM4ITdOYol+DoY/1eRlAh3VOp5YumUMH55aeWFjjv
WcCIjCHsBiOn7162lquPJbTxkGPGa0uahzy/+3gIhckix64vk1kpRTUQXKIa2Alk
pIt6GGZVB0W5W/Ioa111p8SanfBi3/U1nbWzujEaTxq4pIa7w9Yj8jMTXbiRJOBc
2rMvxY1OWY5cqdTBnqceIl0MU5bRN50J3vw1ESZCCUOQNJetDtjEXT6Fx6cJVB9W
h4FNCzzy86CXAroAq69Tg90A9mvCFn5pVINYyYYLjffdVYZjLSiKlQVvP+nsuUs+
wlCDAdwmGsjPzU0gYwr7nMZmOXxFXYHvJKrvWSVKdrPuqotsuqvpZhxiOPZkFG2E
okQ6CKTFyVU5K6OvLoaqwIQitFvGvJ/L95if1fxFuN8L6xxDi7Tj+oFQ0WqRERad
741oH7n/taHIuh4fEZRnpMkvOrIKqV44T3fP9eMapSdBUdRQImNhHWYef7V58v9G
3Q34/BIEBfrRV3SWKpLFaOIsbQ2Cozxa9VXhj/yFJcdTUW+N0wYKfZ3Yue2VW0k8
m3k7LAUOR9aXNDxyu0ln3/XiKxkv+7B+++8kQmdVkeyOZQ21TuEtZcgqaP9VZmHP
31OlwTDC7lw2pbqu2nc1QCI1e/xyPfR2ou5vM41fjPtMkSK6WW3BwVCT6HMOLwog
aLzbg8L4mfybrmtTh4b6oNClh2QkKXN1PpSNZdjx4q/3/LBB7S24qjQKbWHlqe/6
ItnBLNqaX/KSRV2LoIMrbZxc2GW+URA1L0F3Z3kDcf2PAcIja2aBj+Fn2Kt+0QGW
44vyGGuYpToSo+Ekk9KejRqoQRWI+hTNk+n7uWkKtmL9QETfOcXJ1pCSoyiKlhDn
JkBGWULGMsQYwSHrBUi7cugVxoQ009TCbu9Csr4Q4fdZ3MGbk93uY1dCLtRm4IkN
7bHyRFDWkFOCX1ZeEji/mXUNwd1N5Lx7l1Ej1c8+9lFTE5hHP7TZTasRDw1m26CX
gxHy1uFAo6k0IuTzh+kugrQ5BfX/F/sZJ5MZ1OoTs4kp04HfAyb3jkjN7SP14R0A
RSuOrcPFYYblMyEP06vBtdn4l2GM3n23YsTRWo+rCzVRNqFPytepa2il3d4K4CMd
uGqLGKNZ3D3fHGreduhRvDyQJPu9EjSZjyUzBoAU5lSex0x7wn5vs1itaaFrMhQE
qvaQmqQzn5bqRZGgbv6RV8eaDSB/1PcBe4RcrtSsJLQFlVtplgZoJG2yHPvFMK37
LE+GJWkk/0xYM8Bi2BR9Ph6qwMKKllCHp+C8ZDUs9/f4vGTbyXtTnDvxNVvHiYYr
CDFn3tfa8v6OGokJc5ZJQzCZB/IWUjBaJQ81f86a1XoNhfLMrxYOpAqicwGhNzWM
AiDQPJMxcIgF7m8TuuYcRqAvmNioitCQG7qpzjFmanNoRhivq3QdnBbsEjxtFLbs
ciaWKDpbtE/wqCuFdSTy9pR9D7BPtrpoux0VMkKQk4l2aZEFctxZz4xF1K2gJCD+
aa662eAODTolRyk+GSlzsQEcFfI9F+6Tb4o1hv+uWPmz4yYFCCVHmQ28iGYP2rH7
POpsoaoxEWV25wc52DT0qWUiDLJqZeo4CjdbfRMOS1Y0G73kf7d2DMHq6cHhOVLA
xK8Gq7hEOTjMHKv+7eMnb0/eGK6NjbY9deLX0g61g4MCnEqzO+gVfs6TUCBlXWyK
l5xaipg77v99iMUcMHGWY1v72Y/XNYlV3JclVQepnqIy3SUgLujQQLqFM7r5raA+
Gpyy+hu7H3By83+QfFhx/lDb5XRNcuZYYhnT4cZXllL8YwCrHs5qeS19IaB0xuJC
FNCmWhLgsAeeXdAZi7izSbICm45Ub16XoF6CDX+9KIh1MNOObrYUlIpmNWFT7huq
1Bc6GQ7jNLr1fxkrXRyY4Bi3u+z2nxC80Y6dUziAp60cm6wFBPZzUSyXG58DLJ8G
iivh5dYLrU1hTlwEPo8EibQo60xkXUlICefx8tZmUA49fvw3J9rKagnatAa3YHPI
KIufXiShsng5REZglqtMjgH4+SL2raZGlFQXCNw+RLP/OgGW3+kpcwD33pNBt1ll
SBFMOA41wHfIFsJibjkM5AneU8bQY5Z9se25vldpFJyt3XWgtDyYQ4mq4wNZad2X
cNJjmz7K2pT8MjtGUKdIJi0Z485V98rrO24qaPnT+v47OrvEOwEzgI7JkVmBU/l2
ueKZjvN7+Ii59sqJbOgOVtusUOAq9jtQqu33sO8/GVUjzh93DALQJXCXALmVAg9P
oPzw0VoTGoReyA3ALPHlgBrEeAhRiHwRXAYzUNxGF8pgumj3+f61OvLcMMfUkq1q
iwra0uSiE9zaSiTCI8lTTfs/awH1NeucNy1KR1tY3NWwZXS7wrPwsndDj1D1jHXp
i86hP/E+6BkIieaGvjRULMnqH9HR2e1JDRe1X1AdCVfWPn0mPcpyL18iHUtWidPh
bjDgdKtxlNCqR6S6WVkw7Fktl7/BaV8bF/KcKxP3NnnXTSD+K/9JhJeasGuihTIZ
X2rex/XichmmmucWhntyuFG/tGQ4dJRWCAtZdWb2Kyo8sbxIC0hZSDDhfXhUkkxd
vrfbLLXhBEaOv/Q9smsfP0JnVTMOdxgcNNsxhzzDKQlAdi0AtrUAEsh8sRSO5FHV
/Ieb60UoMJZNP29IeVsutquglMSI3gUqCu7XNCePc1EEnsQt5wdthsuT/6UWMWN3
MQYK6oQojNpelrfHozc2OXds9JxQ0aixHwf8xxQqRp+N2I4ZGxKvgszTY7mGIthS
UWydcYf5oDofcjOvgccf7r7NSPVlPafAFr4hU5DfyVhVhF9ut36DL7MvW5LVBh7T
c9an2v7stzRYMac5p7+iokvU2bM6HowFPZicDTisubLazaQb51Rljk7rXCzVF7ey
OdWodicEgc8RINJoClr/uUdC/UBf2Bco/S1yFLCGsVTgt7UOym57KpDGUsgndepz
lbz6Tbq0rrQS5MapEZVRvcvY5EPPCBz2blRyAIjz8iNfz/dF9Wt4ge5nrfvOEFuE
tvbtgkzHHjXCbhMliLZxo7Mpbim6Ke2ivwqhy+xijNoWtoirjznJhgbuF4wmkj3X
l77cT2kwsfW6KpPzJ/4/PXDYlDbNyDYzukZm2PWvSdCdVMKK/+5Y0un/aiU+C3Df
xPzq420C7qp3eh+JBFeL5NNOsRCs8kbItMGT3JHzs2skk/rdHaHdCCxINwlWw5Yv
3r7/oD50WJFoeNuiTn9DAi2p4DC4Qdvyqs/aJquS65MNp6QA+LSOTPIuV5601cmo
bZLhGIRxterN7qXWzZCVnHk+ahu57Mr9cX/ZdUOcLvNf1PI8dQ1I3JAHOG4IEya4
zAP5HsYPZkHUL6AxU4lratiPC9IfRBx0KWg57a5HncWhH1XEJb43H5DMxypdsy/R
pRnNzxFh//5yOjF1qKxn4JXvMCXZCoGSEEA0oDZ/0pHcPbwPYAaTwexSvB8JWjVx
yivWCHiGoAfrA+t9L3MNDDMj5hpRqJCdBM+4VFstGMS38b3NNSkwtjRxQQK1yudi
XyLkc1sKK4/g2C0nU2KzvtpiYStelzE4BGQSHo9oAXmPtq4r+3aQSHlH7JzwT9pc
EIyV/3OcNSejMuICds1+SyeOB7Q87UOL4yrzNY6rI0fAYbX+DeWD0FzTvNeDGeux
RJjgngu7jLEOakuLQkbJJwSaszBWfda1Y2S/QjWwP6Fbpaxk1ipn97uUqcWpFWmG
HPGbZ03o+YS0/lVY8Rk5JUXDZYznF1TTQb6ATujzXEt4voqUXLL/uRamtta0Ezth
deE94YNFmI0RvohWKy/wbdW/d3ethlIzwUqBopz7Y5PDZ4vDMexWBS+a7vK24e34
oJzC8eyu4XYM5yx6DQaRgBsXh7R16rEYc84e9U18VAuNZ4cpyeiljBgxVA4zrKZD
oHzDGM0Rr3O1+AHgBOY/Pf24qrBW7O7cRRGLyzm01SdrI0bwEa6KHsBtXQe+ch0P
BXFKs/M8thGLaOeu28reMbCpWri9gx0iNWi2ULtOhzQO7YWEYxIdypG4BqnMlyDw
rr3IADyZiY/64eK/fFZEhhcn+r3ZUbbppOq8BTeJtDVpow9yUtYWPNcZQk0DXIuh
Ntd8FdCbv/jmMiLXaPjiVe5xTkHQ1o2L5MRyH6Z0m+sZxuMpGtcp4/DceND/bQaS
uaw02gPRRGBf1MC6Tbzw/qP2D7uhQ3HtODTRnCExUcGOUXBKATmTS+kg4gHCW37n
7JH6JZ0yyx/WtYPPZEaEiydjZXM4bzPJtfSeWV4E7Kb1vprHBiORV69BY8/kRLgT
RYFZ5thEzS2n2BiMMwLSq8iSBLvB7UbF34WCQswyZwqQNQx5w78EjzjOVMzYNtTA
jD5EgYJqOr+2c7akigYjm16NWW0p5EWcb1WARs15c9F48i518UStux/vgyKtAWW4
w0sIuCUpDh9hvzthLUDE/llIbVwngdR+Ge1YpAZMBTPTThnyypeFnYnGeDMiBNo3
sHRR56g9riS+cvnGYMUMOfFcipy1RUvMPHXQFBOV/2wsGJ3weXe3ZU7ytvwdJG/D
6DuHnu+Gtf0XZvzUmqpoOdHypIZiZGxkA8RPLOuDQB7PRiMUc9+b4NRaFn777CRF
iBGHM6kXqmJKIUS1jBSYwX0ZTkM2We3DSU/16TSoiquK6W2mOjHp+oxplShDHw/V
PkZb0X8ECA1Pqc4VaBnd0IBxG2v81Tqpv43fg5wqx6lP9g77TPj4T2F14qnZR0MX
Or5M9tFwd2ROhspR27E9RRJDsNw8VFJcJuDXkyq1ej1SPtrByccQMLTODp/x+aER
we3w7LpbHQJJH2PCZDWmHWpDwkYp+l8FnjVN+lWkrO02W/tMztQ9EQYF6GKFeJdp
pcU7ghoOpTwIhGqfYVcXvsbQg5gT9hzuRpobD1IbvnLTbeLqrsZTTEseode3vgyg
Y6P8NnU58iWpwr8GXkV2INHe5DztlVfrtmsXqaLlcqQovQQZlRebaFbzjOcD7VfP
MoOpgOIQrfVtuGYevaClr4ELpLcI1yK3qFVP9b1SCEGgC0i3QmFbw9RPJ32GJHD+
dBmGqUXzycijlyn99oEQvUZv9U5SVjKIKqNchwxsDQKdy70fI0DJc6T40FHkzXkK
MKzmB9VE/iuOw7JFfQoAuL/LfKpW/pPYr6KpqS9IbYM6xRzPs+qxK/zeCd8S4UF9
F7hggFwTa8qhSkwF9EJNJn2WmwPRrEzitOTbYdVZUrHKNEeYjPQUnb9Y2plA55Fm
75bc0HZf3yVONBwBDFsMBHZWI+yxsPGPgRLAcrVsIWjI1eA6NpJp2ykKUlowy+mS
1SyU67SZA5eIbU0q8QM3d0BdCpYhB7Ju+nH7+r8MI+/psv/jjphnBnosRPW9qWiR
Gi36tNB/nj16TIo1VOVEPHUCl2DkCUI3n7SrhTYWJHR5li9aP2mc9WA/THaEh44N
7STYrQQrz7OjJGLV+Xu1nqkA3y/bIjhL4qfYUOUzq0fMWmGry/zKluNO+jGhFeJp
81N8KHCSX1xsp0S9Y9DYILfMVgxjlhO0ByNxwVpERjCcBv/if9KuPa3r+z6Z8kgj
lP0gLqO9a6rLxfrEjxpN7f/1bw3LCsS6OOAlRMAxqLwSDo30fcb1sC7HM2e5qcAM
lauCb/n30LODcosh6szBWyazvm0e/L3TDEF0NX2b7n3mXu7WmfVx9WBdoJLxxc11
tn2BpgIr815TeWmRY44Zcm7IkdmMUjrdSqN7PpPH621IrmyIMhCvZn+FEv2tn917
mFdH3lMwAmwzvV1dAJyVHwSjpRQZJAkFCCbBZHgK5mtQYp69qPY2jjzqhIxZRPjP
supCfFBXDA2wN5cxJwbyCuLjsUBomtrVLjzV1IYWLUWira8yFrBrvOSdzQ4VMxuR
l3g1wGPOAAfYN8AWhjc/nExqSPJrl1Y9AM6jNzjvcpFyxUlsxpxPwjSqeZtoIfxW
E24noL8GrSpW1MHcIAqOQY8HL2embm+Fhaca1NfGRuZQzJIcEYLfDjz0CSjrPsyf
eMkd5AZ7qN9UnqC9KFDStMOoAeHUrq8X1a49CLTFMwQPE1Ndxt0F1IOdGzGAj2nK
b8B+54h8g+5/pT9sd6S4w/N7Q67LvVeGO/7nAELiEG+VUGrWmSkWRXBH5Z+jQ/sU
PZX3F41XUV0G+Lw9PSjvIPw4Efb7wvcIy7NFjHbavKnQoaMhZkehbhFmf0r3IdPk
J94v2df8NUGWzO+4dLmVpb8V1QRXHhQ2L//iDk3p9j+iaXOTRJKnDkMuErxrCnec
F5bqvTizLugbGXVJVXHNK6Pmsi7/eMGeurWN6GBaSRGsvjobvxCKETPEbojXSkWz
d+h0mFQpS8l8T/ChkuxKT76KWoES/Bg+gPB/Z7F2yJzlx1agOIApIG0sMOGFWmbu
bMvckKgUp7B+x2DoHZpfBvhWdPlRsZnkXEd3V8sIKEOXJu+jm4uT0F2nssfSKfFY
ex+xQ1DvwH6O+UtsVQLKKgfOD9seBNRBS4FvWnIeqYOI0zRQIkK2Uftdwok9Puzc
vU4/fqeSi7TmNbJpMckoEwWefEZ7FYzJk7KCc9whb2RtkRz7O+F0L3susDPLRS4C
ac697dQzOFKHlYHa+a3T9tqywRjUfRPdow91LlYY/1Ow66W+QJfLmiDHoSuJWtRL
LZZ8UWzgwEud/9CSCFRlwkngoqTbK6hILS1sVahzoLxEaFzUj/YgAfDVCILA0w87
1W0TONn1NbdRHdiHTOTZWzoz3v7T7PAj+WNvJlenMTXz36JvUrsFrxVIrDvLHdXI
xtHPy0jXYFcnzOYsbilHJ9B9GA0JUnwZDGSEFRplu0/+qktKKfKaURFdHXCt9zA5
lfrz974h75OBS7kNLvVzrulpmdm7H155exF+Ep1k+zmpYHn1vdUbBGegKLzv5XMt
XtLgieR4YK/xO7oQArYTLbCsVWzkTaHnUIdPvPWFXMT4JdihTjZM/yzIm00Dbsto
/9Nrg/h2YNNe3NVrl9/0mUcAEgnk9fl1mdQRJ6zf1bbQtQNxR65RK8UDYiXnlI08
V4dJULpXIj6xzRYDF+2LRNaEYdKWqYns8NzS2by6i3DWOhiQkGsr5Kc35HIzhiFM
FQrSYfPTym/l5v+eLOJZjn/ooRVTnZUvDkN5PJOqC3RehlRCfIC0ITjqNVXv/rcG
jHSsO5ClYQwQ2w1e7R6bee+4CuXHQc4YncGYPYEg0Hh4qU+6vCZeaexSQnBddG4P
2DwCnWUsYIzMpthPhczkU9IUfl3yT/gislWWWmWlfsMwYOiwrdphhaSXP0T/goht
cV8SmBpWWu1CB0GhnGRjNud70AXYEHnXLbtQXYRpqecus+PkGJ47Fy2G+sUom16w
yYcdqZ/oyKW+vpDtspIX8d58kZKwmkYN0HOAmWw8mUI90hpH2ILuXUjv7/OpYQvi
Dq6+9xSIXt8oXlexD7DDu5K9ljYfqJA8gBcEmKGnKE4qJvaNLsxq4ylq9p+iazNk
jDYlryADj9j4+AcJeJl6jlAWIpL4d1unPp1I+qi6rZWBGIgkFO3Y3hUcy1ChhY82
s85Au2ngdZw8rsvRZQcfP1VcxU7kpMZFePiQ5xWxED3Qun9+ErevMa66kWEIR8In
iTicUeMVisYetZJlz04cfYm0tRigzN10Ub/Zu62CXqTLb3wHu1Dj3LZO2nU3793M
gw2CppcLyFzUxH6qGGo3/2pgXlTo5n/n+RE5XjEmo+zoXCeFTvl2VO8tDK37leYF
TqZLoUFfvlzO/0hPwBI/hL6iktFZIdGKVGHqughpHqNdnPpLvC02zZZx20lDzinB
LeWdsGC4ov7gxoFd8FCL3XSnlq+IPjTBwgXTRIMafn19cC/5fZvfWtfAVWMpabsl
a699Vm8/lX5omARKvLw5ghqJt0dvdqE+9PsH5vXAX1kqp3/Jos/QZtUBJNnP0O7j
C+k3ORhCXQz8a0PJ1NyMvPm9kB0eLacig5IGIMGjyTwbQ/xGi6mMY+LRNLUbblci
55M5wg8vkkBWLa4RglI5x5gE+glP5INNkXf3KSflg8TGyKXfYTrStcfNFYzu2HUE
MXvC2WD+Dd2BJQIEz3twAbv2pfKRz6iy4+Jbp+UMnWyYy26BJVPm8VxzUkKV6+54
vzS1K+O2SX1Xk/Dc/mHyMfN+PmvlCs/6azdBw4YnDdD7mj5SP25bFDRDmMK7p/Ki
gt4r0vxuwnHLWWgI2zphlrZ3D35rDS56FjtTrKovamuzWbTPLtb82mMjwrS9R8IX
ZQiw5uM0hu/KxxSPr8OfWwfjZ471rrZ6vCKjufnAXBkRq+UHWldKk9HPdUbKnksC
fz1r8owthh+TGvwpVnvzDb7QwO1gKJE28TUHFvrqYE9LnwK8oVMfKkub80R3gtnp
WviWE1EmN8Pt34VdVwk2MfwpMCl4EKAO3D+6nHG5eBvQZlyaBYVf0OXYcHdCCU16
0j6JqfxVJEJumCZVl5FRUfsCHeLG171A3Vc+3d+vGNvQr6eNx+4EVEFezwahaBc0
GMPu0WNPz8W96/H9jrUWzOSwxMVrGHt6f9vTZTBP/L88NvQewsO/bbdJlMBMVON2
oLcoGilh720q8nRjDugns5Jjv5fRXqyKAULMRir7r31KbNZPlz6/BZuL+mFL/Wrd
4Pa5szSZMZVPS/CN/fkirylK8KjDPzEgYFlnnLLcGQ4ol1zmnL5X+8U0TDdUeRzM
6QgqNuRgY8XxyTgK3hAG+J1gCw3oLUCVad0GmX8ZM3c8adKURZWwOk0NRcD2Ktv7
TXBsAoaZJH5EpeTRXN0Xy+DrMAygm68QaZpu9innekhsnUbRrQZeAE/hUDIyR/Ve
W2b9vgEfu4+mReOsm+7FjCnS7W56pQ0y5gw6AqVGGSufor1YH3a9yLy5xGrV84xz
++qaqLwcv0rDJclSvVSgod9LySFAq9jgLKCVTJ3fcTxZAFs2xgdvv80x+a+H86mW
EbDDonzod4WFeT4mxPiNZzTNYiYEORPKzDFwpCouMIEDyyijt4/J5YtmlZvrFmBG
yM4WMJ3Cm6GC27qayBtQ42m/F1WqIsXPF6anBxuJPUebojWNdPZ/Mlqmx4Fv/jOk
qeo2DVVdxsZWGGpWM3mHEnJmXc2i/ox3l9TByuWBXZnqNLcMTLBlJR5OXw2Kd/Ee
3UvJPyijjNl+nz+dGVCD0DDactxlcQuP44R+MyyvIQMEGYOI61gWw8Av94pgypP0
UXLxmCD/khCjqUkT7vnYF8Kjy+cGUiUt62jBevpIA59dH+zb0BWpNRx47hSbFycH
sRXA3Ve/V3T5MxZrWqqEWwTN9Ka+YIVenj4ol1UHt/JTU+QgodHf3W8L8enVyWWe
PnVXT6jCYtjulfw2vjHI2f96rvJ6EFhgAE8kWwBXINUJDfztvywoawWykbfLDdKU
u6RtaFz4PwOLoN24Peib5bIma8EVDOSdWZ3Xho5qX4KagZlRfdIiC99PBUTn46Ka
pwZ/Beiff+uPFa3RKwaJvaysoqN7qiKfDqoSgPaCInW8cALLobnWcnp52S2ZgzVs
rdqedL+rkEAbFChvhSAPFd/rHPGQwOZ6iM0j6UpPVIL5+0M1gBnJmfffZJ9Rvc+V
SAvrSDHqym7XFCs4Qip1J8lJoNMmegLSWALpz6ZcyvP0Gj0XJJ10x10K5GD7sIx4
PNMiIuUwPFgecV3t6A0ai4K4adDgv4hl0uc2r0EkaCbOXx52Ffr/PbjZSuwk5a1x
lWXQlQOraB4O9zatbRWnxk33oapOW1YKbwOfGdPyQ9E5ie0HO9JVobiCFl6EdjA/
wL160xS++e/qEg6hhE/UqCqA+Wnnzf7hHZV/WkcCA/INJ5h1g1r9XSyGTEXG1dVk
R3v+X3e+kkGA6XkHTT+mo3AfP5iadjzUXtZa98K0JtQYXi3ulqTadjvicFuFhnds
s28wSlBPMWrvkiavzWzsBcc88LpklCl5AolZoejDPYami/qCh5rpyOOF4JaStOUZ
kKEv2IajRiTfIyNrwgfELpGbiWqtBUVoy2itxVCOVrkjoi3/0+Ml55Ys1dIML7JI
Wc6+dJsXX3PvLPjpJTAKoRMOYMpdMGvLersf7cRSMPXfwmBvgDdTouydkYQ2qvQc
L4V6bCBYSCj+4CrNMmLB3Cq8qmAvT4WoflWr99BWIoBJ0bx++mgNpLYWbBp+otow
isBYQDxExFjJTWcIZEVDBSJh79AX1+VMe0J9QilRM2QY4983ns+IRDVSwdX1DO6Q
89LEExTlddQN/j7nWdF05sIA1plni2v4tVmoojuCT3IQS2tyFzFVGg/ZF+QUXhoj
wTFDOSSlErldMuyADH+9O89oph15FY4XzNmKu5tx9V/Ol9//LYLCszrik1vwxc2W
xVkKLKN3FN+gEAO4C3H3euOZv3Igm3gTuj4VS9iSYe7rT6kkLbZR/+lyTSuQfx6A
pQT2HDmHb2Ua0WIR354qZpvnHlHU7rjMQ+haSp8tf6usKc6yQ2aaKvD6MZfaxIl/
s9GYJjE/k8KSFcf/Hz9lbXGteQEsQ8uQS6w5t59mbnGaFtTHF7MKogGgNmM1hTJr
GkPqFoX2S2Sgc4IzloiGpmxn+qcH63d/DX9R2yK6cn3SR0jdd+QfRAmtih/ycTGS
WZl0CBQFmShraPQRwWcX6SmVAS/dn7EihzbqTWsljug1VVklj5f+oQ+Aq3I5ZEjd
ysAL0nJNyprpWMm2P5maHhzLDLQmCFkPCBrB0YgJ9P25KlooQRLgjE/2lB32bMyi
cab6aUtp875BgY8IxVQYmdCYwtfiCE1xC3HzJbex6bQcMQM6PL3FJ+SurrY/g9Wa
9ckLai6Srg+3VBE3yw0XNQH0lHQ6lP4jj1WfvfTcoqO4/jU4OEZjzrmld8srMuAM
Opzt3MWoQGQxxK+WX3m5FBA+8v08Nlj+JOFxhrhUo/JpRASal8/2pMDtBz49rsFB
z9VNoM9xk19IWjnWPfnB5rCFNp0mM5q+SxyVXoPraCuMPNNislMMATqzHZDk+0fR
LRtInmIwF46AuBpndE5TFZnN2fP1UC2o9k1sH9NCF+uV3JuO4urPiD0OzjDr0s1s
1ASmsWGWDNTl76RbGuHbDfzsTKeLF1cT8YWV399G66VU2ZRBgupSVazubGD91gy8
dMHT6/6A8em0VxnXw/6EZHT3WSm/c/1PqBVrlNZ9LcGPsT3/zKZSfgm6rZobgJUo
1FxVh1gVGJJhpM5uz50ntzK8z3LfpwTLu0dXGaz+QTBKt7uMh58w/PNsmcWqsBu2
HAZvIrl/2cIMmRwjc94tQi9mUyLeshmkvUnzNSRGeYznnIxf/8VN2z3me5+PwGtC
mMPtBdkcBtXebuo9ZiIKjTw94vSQoniTCYDHPuz5aEbbdf+OeGD4zoa60lrM/Teq
GbJhkQdVU1U42Uw6FHpMR89fZB85ormOXut/NX3z1NrDRbW5dpEsox6SHVaqkTYZ
rY3p0ZCyv5gwgTssVEv78J85vlDwWInZCo5/9wyYbg/MrEwd5IsI3EUpSyCZoAWa
wh+NEbsTFW4aU8DO/GzCM+GXAChHPD+seo2Ur5hjyMpHeB9m8DxPO14RIyy7SGlS
uZAl73uzWlL1sDdg9ec5R2fstmyhz9yiTKcxbFMxya8vwW8l4mXcoIxQd++H3omb
YyE1JJ50/BaIYChlj68bvM1eYPhNbvsGQAi36SPnL7FhhuDzaY7KzMepB7eV6XlI
fBQEov2CDtfKAHwGDoX5LxMD3Uq4YZGFHZqKrBmEjJPgcMy/I6R63C0BBy3WZSc3
L60Y78fsPRewNgylopI2n6NKxeUqtSUMgNYU8pYorPwIHKwA5qfLQ3/2WZtQ3LnS
6mLdGzAbP81E7VCUz/HyiUv1hhiNd3wBnnV2TcOwo01QWcI12bKSkDCv/D0mkTmD
hwh+4uA0JohqzNt9rtKTie9bPuS2zMY+n1hfaFbAMdecKHDALloNOFFAWV9xqVVX
JVWjyXevK67CM5GnNT9IoL635tmmEv+sBcFSMBhhc1cDrZB+yZUuCe+oOaz81Zog
ee1X85RbYt7XdMc/FIJywi5JOyWBQTWhHEs85EmMyouiP90DDUOBepmIHNrnIeon
quiEXaFWGVwPb5HIZlWbVrdqDQB3eVW5YpaACPs1I21dGKDTsu7Pt9EZc3PvyrJB
jA+KwZB7Gs4+i/7TLM+opKy+L8C2LtFPDCqDci2LpYqGV7DgdJhPKADZD13ELk9A
dNvBQkjVLAnD/um61Qstb5WVipQ3KPqxbHeYz5htbjEFss5JzVc5g6n4wOI6h29G
yoZoelSe13LLkWFcbE6oLrwYy3Lb+gnTXZTvppqNilwPcixP90j79GXliaF0RsMG
guBqy7OhDuNoSMNarfyOr/gfcLy0WsHh8C+r3Te7Bet/9g30J/VGqhyttuYlO2SP
Ua5qVMSqJa9sHtaEaaXrmLzCcSMCQ7znHAPo/H6JDWjF8y9AN9Mas/bV6yOK/0le
A+/Qzsw723wUp21DkqT1lTmOk7TwVCMrZGqo+Zf5GLIUSUqg+wUvycc45yMQV/jK
V7OyBJBZTh/cTjnK+DTez/L68L7wnilUclR2/1E+3NiiINA9Zk94SwhaGRUWbhdp
DPZdhVza2tMLA6Ko+wGSi+1f/05m4Ity/yfL+/4yVTfKwEymS8y4oza0zhanyuke
ZEdcg1qucM2Q/zCZvSZ4FBTAIuUF7HTPqAeelwg76DDECOmFNn8kXehD6hygNBhC
bbizBPKll01isc2mDRl45mzZPC8D3A3LpjlG62wJJnY1LNjWfwKKE2psx2gLH71a
FoyZz1sBn+4vFR3nIRIKkCdJrOVamjzvU3VcW2NC+XMa4x1SdCB45V4YIk0KXTSR
QAjEwDM7+/UMUxgavDWgpVbjOD6cxLLIBDMU4p+thzLBkf0Gr71pmCh8pKi2E7AR
FHc9izTo/55pApHqX+/oBjesTXzDS0czkNJzLSEEmld5O5nuYkbwVwRaFgXSqScQ
MB57iRIHVjUR47zkWPIRfyxtaAK5WV4BfKjaaQeTt3ergpOiTnuyQxsxyWC8yNgA
20evHUxE+T79nDo936tbaY5FbfKxqjmTGWI9H1rNhCfioke0vZWWs8mLZ2eE0mwM
F42lQA3TduWLIYMAKgpIbFV1443GeIqN7nT3vvDCToyAeejs1O4PIsmFAzMLGdRf
/+NMHbydfHDNEwyXdn9kbSY8M54S+hH6sVTkD72La18WG0GyXXu4l7tBUQBjN23C
lJ2C+ciq+kBlt4pynfeA0Y+D7a4p5K/5z8vAm+pIk0iWmdbN2zC/Q5VyaBX7yWgi
B/lf9HhbUax1aoCInzGwoRs4QUZeJFXbG0ir/zageGCYm468mt9+lbZPu/AIJolp
1wn/xLoTh1Qota8XhqsYjWwoLQ/HB1SUTlDz90eR7XTMKea9Rx4CSn9pDiI68gsL
XWwtnU78R8Ypkvw2E+DO6S7N1X3QIGWMLAxJFdrkyWJyFwRjXuBQP0/Le7b/7ser
757GDPSZzifFYF4ctEGAO47H7KKRswWb8106+U13KN7dziADvh9cjc7RlUlTX/PF
yi5f8oj0AmpAE7FuB8q58N3tOO6XiijZoiP4cGuOtr60jIcpXNpp/bbtUb2xcy+X
ctj1ykGZKEeye1D4WFAhquc6sxHu95wx4nux8+Yj1AWskovx2zmhxjuVR+KM1H1P
EYIqsoxIXZWCBdlPQojt+7n3cvnY+Op/YXB5Ws0W8VQvyC0Tte6R7iQeMxzY1U57
gKWNq/mf8Oy5x2/ZIPFb2S8SboMNJ38pofGPPBNGnFDquOmvvU03cXpJHXuek8Vm
+LfGavKkfEDAcV/e0rRT2hoqe4l2IqSgr/G6g6IxAQKrjLYXgPmx1q1kM/gDPqt1
3LzlJrZZlNSRcjyoCRDhCnF+g7r26dFADM50GQerfmHaVXbbMc9IiyLhvIXYSVlY
lAljc04MBRbEq/rKQCU1Fpjjpv0ZosFEmDuttbPmnMIAeEjKZS4kf5EYjGJ5SOpT
7HekbhNBLt6KvCBj8lzKxMi5t7x3SvZlTK1h0KBuaq7DFXl5u9Qh7qzjXOJgJ3PV
/jJ6d2ngyNJq2fIy1UcoMqB48F+p2ll078Gz2WlriLe9cwRi1M2LfBpaBoevAVnP
uF3+iovAQ2+Xj2kFnG/NB/nwYRsfbRhCLWxxfNNiIRq3uguXJhmyIM/Xb3Zsz0OM
r7ZyY5F7rf8qy0bA5J7VOKqlBRuzRa4wZLEl+TMbvmJ84gSZkHgTap3UrESdNNY0
cpVFo37Dp9CzRZ37eYRB70SArT/zMCkmKuob0aKyx338QU85MborgC/ZZOgLceC9
Zif1+lzSWHoWtyzRBQqmmNGdXfnwNldVbd1NXq8a8bNu0My4u+yd9AMB3fF/RB51
awBsRH929oRlJsBaAdLLEf6dXnSB89d5mqRIb76A2AMvH6H0znLSmfnFNtQt+Eow
TlEc2OpBrSptVFAiWxeQT82bs2odNgtyYdqDXT/7TdwgTFqOwInCwtgsMSvzBS5I
JNXTQesqFnl7uQfUJrOXnYzyz+N1INiYbtL6XXiHQa6k2K/x7FaTEUrDAskLyRtg
+KKE1SjsyDfo0MixAHk84w/2RXrrcfjM/1gP8ozg2epVDD0bUCy+U/TeEG/tOG/U
ODDWwrcYdl1n4FIN9nFeT1ajCtufVKSefZe7AQ+UD2TPygXx/FuC0KDkuOriu6oT
SRaX1a161ak/WVMB3UPD+CR6yTIJ0dgJFzZmwbZaE9xjrrwKn7bU69ZKwZ6JwljA
yf2xRGJgnPNln/vBJDI6gx95W57RHhEDmG1lKGa2UNSuH/meoa5kAk3aj5mpBryz
k96OK2XHNwuB4Srra1EiQcUqKSF2bIJ1xnv6SIxuhCaKUD5/UWp+o0ZNKGRPhzuj
b2uyE5uJ7XsrlZ+dbnEg4M9mYKg09ZQuUQgcgfEVlFhn05vp2tJTqYHJTjWclst+
H++KNFgtwGeVl5D0kudUGXMhqjsbsq9OkVTCksHsq514edF0RhKappdN79J4PqS2
SNKUI/Dy0v4TMmlje5FSMfp+uhVffCki4dgrgqZvr32G+t0hc08KPhpYzG1f5+tN
6jgVIaoKCM5uEJEEyylixWCd2zx9Tf3VeH+IA9PvT1hDsD9D+EdwoUFGt/EHR83N
1v58kC1AmjYW2xqCH6zF04yAm0uSa7eZ87mpL+x1Tx8O2a+rM4t6EDHo0a6dAkSo
qEzefQoPxB4KPiokVa9wxPinhlIoC7tEu8FccNawImr/ehCNQX2vHcThXiefcuzL
+FusUrIPvkDQxZLSlZgQCDdFTBOeoW8LPJvPGC4mxxQo1JLSSdH58qkVlAETLXZd
lUZAoqloF0VpLMUYvFLG53BVc0zFwcTp+04MjMAZN1SOs1zsHHxfEQCg50/zP7in
2jg0mIXdR3K8xZ2t+qMjYuY6RjFR1rdcsnpgsgw9FHTfak2bu4AvIZmShXRSfSeE
zFac6Plo7FaKNcp4wVg7apueloTInVorx9p5ewW0KZ3JvS5+7kFTSlkcTJhC9dMb
EoGMqyJeB2X61xjM57NJs6Vi5THVnFBhB/nyTP0KLoJFceUQnJ9UKX8Q3UJR4aCO
H/MrrSAOthUNV/LnaEirQJSbv8g850XkK8EZn5elA3SUji3qu9V34cHn8gI3RXGE
izN9xnaJlwICMXHjf5LLpGhS2oFXSdOrzty7B6uAqM6OhJhGN61U90kEH8GLOTdD
/8VHrepyN5Ewcx1tXwIYSyPPLtbOqX6JxzWd/OuUKyQlJcEkaqliUJOXqra7YA12
nxxtLsCvOMqsu212Maf9qZzCkfgNcAakpmYizVAC3LEAm2jWLf/IEDaKDe6orisK
OzLrgdDvr05cHwpjg/w1PJ9xOAPTg32jIhnIWGFHOS6pG20vAb7s7h7BmCITZ41v
W63LgEknJvXsYVxiLvDlmLbEBFixaGuccwZK54f40KQ38G3bpbRc+5ouQPZj7jXO
pKDtwIQGv8AuuccFJlRIScE7QQVLlRrDzla6mdYSYe8S0uV7vcYQpI+mTCVWNeYB
liP4w3vmMpx51LV6J1kEkgnqW99umG6M2nC5p1QvX7SeRcxIpasx+1ORWkUsna8E
VXlMqhbIcG7kgtt3b0Tk+RBiuAunyn3SEQzLouLw64qToEIhq//XptFbZxCt6ISC
zFrZQZdcS5/slu0I/w0NpDoRVzniVOWxcUdfNoeZqkCx36CPqA48D/YuT1W7Lo1d
4/6nfUN/7l2A1LZBOavgZKLm/0EZ6Acx+kkCAzeXQYisfEz4LObENunYefakSY4O
KJfHuuDkRnDpRypne4mU9WsAcTNjYG4U1bxM/yXCICyTcgwfCEGkewwrwhiiWe25
jAnXnpsE+LVOhhzQhrTpEh2zAQ80/RUfwHBDSsCE89ImiTAErUECzFAF2vKE5UMX
rnRGegd7+BwQB2tn1i3Piighkki99Gp9TX/XFxZlUhUq5tbgRA5zhExf/geB5yIp
wlTUxd88Q3yr6JcR5mnQbiQLwpr0FmgF6pH0ns7aL/IYFIAETg2rW6joVGmfFwyU
3+Yp5JMq8v3PrRdnPM7/4S2ofyfrdIUnLZ4qumqSofCFc0H8SW1s1jiUcCfFETYY
NfUZz/yOPNbETI5lB0h2JwVn2w+VQZkE93KjHWIKWrqo2yUmFHHRNKlyB84OI/m+
Ezl/76vVBN3HgdtNteQskjWXmB+vJF5iVRsc+UrntvzTJo/wZ/FZrgg+muFw7rdw
ztAvIQwioA0sv10P7AMmydZZB8HFQpp4n12mymo6sWxo1rwl65MZnqV69KXpt6xK
lKSkDa563Feb9nNzaqLYLjyPAWgK9sMBexhWgHTahPfVmgDLSLus/NRljCT2MQEu
TGtveLFGTpjT2rbV+vNHTWIlbeMJeBydcnkOCX+yoQmuW6iDV7nk8BzEUaZifm8w
a4Y4R/8v/JaAEplpVFLdg8VAqL0VPkL9UFnUmSDOcD/Cl5Do7H19PZ6yqSAvVZnu
xRy11Fl5gtziLfa4JfzBkc0WJLuYtE0Uerr7sIJOrMKNRB0LfAsXrkwKprjG/gRd
4/UPTAcq2Es3X0jG1HWL5GVP6u0uW312nBZ1zY54RtyU4zZyKIWz8oMCe28K6NTo
JezyR0+7YTOj4NtMYt4ZAIwxGo1eJnZSl5RUR9blDp2dy7GxHmgIUULK4Bs2sBxX
IemtKw7ujbluy833leiSwd4OvVAHB3zn+2kDNYCJYVNx9cPNeJ4G+oZQTBVYtYBY
teUgqQUT+HVSv4Kyn9eJcEvEfAs50ciQNPW+atJPBEcL0tQaqzSBAZAVcUNp8zv5
JzBUYl6leNDXLGh7B+EtIVrKH3zRH3SJJ4Ji68yqshuqrJszMdhC8Tbi/7kezsDm
55R3k9kVO9g0r79ZPZHVkU3YrRWInaGscfZxAkh2eG6EWZYLjx9v7wJboTcY/St5
aWZy8edWAltIL8yTFxuO+HwgpMe/rmvRVOI8eYBU1sQcEyjSMMtnKTzVFpmj+kJ8
rDKyc996jzidPkpq/sIFWZunRrEtqtxNCCGe7XmK6lmcdD4sohMi7GXa0prlwtYu
jYkSPnZUsbGVT0tJGyI466FNcqc3/Gl1e63GI0VkgkBrfw4UnPrQbbxxwiTNxb40
m8bvWzYEwSqU9QrzIZlTNXDVgr4DVTdpQ38oRPmDxu36Kk1L//uA8BUSo+C/ULzG
dejaSRMKvjd/VpN+qguX8dfTd9Cwr9Q6VQCdNnF4ZHmucrQsDyk4gtazTHlJOWHG
ozM1y+uwt/KCz+xBhEUtg1okJ4kyUzwzP08tGROq3KRhGHW9GfvV5NSVoqa1qdPT
oCkVjM1JFYhiRnIfg4NIK2OUX6hIVCqXOpY8M3WJO9JhAplhRsSkv8w+Tv7p/NyO
J6N024n1JFvf2rdDPztkBx3//WSSO5djaVn4UPjb6tmfO9f59ByiBrLqprHVs06R
SNel09r9N857JETpmrjlKWFOGBcL3kprR8dLmZNqB9332rwFnIRftHHMQaJE15WK
20bl5zB3LyF0ICrOsrFurPPbovCY2lUo2HHjMnqz2CTa8rabqhhlh0+5afXZGRLg
6kS4BNV9z+SYgjrGXd+PdwjMrK+DR5+5EEzHGuyM7h3YDf0W4aVfI/Hs92ROwfdA
eR7iPDKGB92nlo3ki6ZgeZSqS5xVUu7+8hKdKj6ob3br11Y2OovNBVG74Tfnpw1m
WXDfvQmPiJrxOdhA0U1DMLMd7FW1SoxGPqELD1YJjll/WmUThUogPdJTOm6fwMal
eXP2IxpfXKGqV4SzbMzP0ivFGBOjDNyia53dhEJdJ6CU6fFsfjFZe2zr+aWX2tzk
g7LX7kmwJ0W8fR32PY4PVuNerB4349OHIo7FH/Hvm5sKEs9eVXLFCbArC4hO18hQ
qeIBG+CkRsDVdy8+vqX4/8I3K5BKoOzdEzOYCfdg6h8X09JU2sDY7bTSIXL+zXav
WXGWggGCJxoVIPaELGClausJfSDURtGDgEh1OfNmS8O9xSHqEwz5RoTbcYpFeW0c
qX3jSmr47Abd1Le8b9iv0lp3LN8QcbJmt6Mg1M1oci4Q6tBUh43GmLVR0Y34t7Sr
y+pkRe8szp640vicaDmyb09U+ZoRxb9tMxhxu2mHb38BI9EDedCR0Ufgg+yDd9nr
NwRdMLwwQOCTsbszAPllaC3RLUDNImZ0ieKvzq5A3gQEZRIq0ZMtX3tiK6lR5op+
lvJKkQ6wMnOpNnXXSye3GHobHlDj18NxRbvO3giHGf9vqebTRSu3pfjkwWvPpjVO
q8FOsbonpPipRxQfI0GHaYHXzbumMxybkEBRWhVMao1SkXHMhy1i6ph99QrB9AxI
hywoWO4+npT9EYjRNzPThJXNNeA1Lmd83FMTpy7a5ytbFVQWYP6zeMcijyNGlXIV
NJf5BnQCnul7W7GFw2OjDyO4SCih+HmX/kW90+mNK85P0sGtUKSZVxNXvtyQQ5iK
swE8F3mlGRmYwb5DgayCgTCv7PRdyvub2Aa0o4zBNkTmAmksHq9Vo6tKZNMplBej
+rzVkxhTbqCQRLa9adHm940g5tUMCRlM0e/SzoXAEeTqWLLKHXPz3gCAZtnJTac6
e1U5kGhddUo87rsRmkE1wt9TwtchXKg7in8DaRrLtHi80lc7l08AxZ8zdSKZtc5/
9Q2hvfcRLJwB2/cFhBypFTOE907Yxvne3iEntSTYZGfFAdSuA6TE7Ylu2ZFprcur
ZHAmq5hN2Z171hJmalHmxwCAuIKjRR3ex21W/vJM3d0QYspVoZP7hymnUtyjKwx6
HkO052V2S3U2mG7VX02lvKVuBA1fXaVJ0A/WAcGeYayOJ8zQzrv8spzBWxRT4Agy
jOFWqXLefaIJ/IgtrsIit7XhCzy0K8Tz2HlCphqwhQMGnzISEo0982aLXGjNueQv
OcM2jvviRu24jw3NT3PNom9QTPCcagcgoXBw6DY5HE0JRvNDG63iYu1AlvTg+6ct
WEsnCvzmePu4MVduGRSKRoGtOSKesutL2gARBwrwmjwusPHQluIWUMsxVwkGSRoR
7YUEzMHhCHsPhgApm1HyMQkbosSxCvnbuLEj96+G4eU3Mr0L0tKsTQHSfSGtzA/p
RwLnmdyY9vEHDn4NjxOUZlCX1RYlqfZrdqLm0hP2MOjtMxJy0/pFubjvBHthr6pF
t5Sil+zyAbM74VdPaNKa+KzDpN8kkX6yIVhzzmBMfFw7OOiO3ylAno9sCqIcwzlZ
wbchI4kOoFCeT5fJUust6qJS5k3HE3vOQxRgaxg5lyne53sdicVXaMWOYMpNj/YL
Q5FF9uoiHmhsmpE9FXP769pZvZ+MdSHqIko414zt8GzBSbyYLRwmKD3oB+6F6VDn
MlZM1kFGS3VI/ZsqKOB5o3+ltA4J9YaCaBYihhg80rL2unvGuMO7sA6Foht5Qt3d
bUhbOByHkT/ufCVebXGDN8jglGJ/tfhrkTVqiVTqu/VVYsVGE0SrBrUkEA3Z7y4n
T2kPj2/TJSjshkOyXKp84HSuIgBrNkWS7E5WRBz9oqDWpx2Lmd5DgJOem//lqeHU
50K5eovC9UMzPY0Y6YLtRcGYkpa5z7zBrPh5uqYW5t/OzlPZfY6UxfvZUx/UrayT
HTYcmWImkuaJ1mhS4w81tNx+CuPG3UEEmkvdOUA7ACzOfwqBtTlvKZhAYSTUsHZ0
QHr+4t8Zq0UvEfYLQaQfYz+TBdfOC7kJ7xugISGEIzByiO3Z+apv0BdtxKYDG+Ix
Mq/Ou9cu8aMNV88vMn6LmWeR76hinbnT19rrRm0f97xIzZRBV50baZP6cJbx0D4Y
mb5PxoJKFOIaysXd4bpsYSSDld+YsBlqrnWbbbovVzNeteOHBud4vZvhjO2SERDs
8ssoVVnxnJOGgP4Xeoi0nqOWHLkCiXxHt6hKo4fReiFQ9lNeD3G0JCAhWAOWHK0C
o85Kk0evyz0hcLtPoUaGQdgg4hcqCmkM1WG6u/yq8WT1q3KBvlNs8VxrXi4ReFUb
gElsPrBy8vzpBUX7SmwiU2X5QYM8ZPL4Wi5L1fCfCkNQAT6MwiOgXfTojQNF15N/
fU3NpZyz7LmnnUCnR46poaFTlWm4amEc39f7NG+GzQjtBP5p8FpabnLxYMH6qva9
wcYZXzXj7nw/5j4YPBOutSNOu9nREIjm2/3FADDLXFYsYJfvf7P5RzB5WQoozsLF
dILAB5aY1dkl19IjL+1bckc9wkRNZQcVJ2vR6PXfV0bPkzSdPvpjL98O2piP7y04
Bq3XqVXwtaUPDgUH2FAbqmRrHWwQeWtLY1oRe1auT6eOULat3fFOQ7P7MD/TmX3T
zGoLtB5cZJLd3uXhMwGeA+ZsW9pLzxAe3b1IXhx17EqAdtqj9si8vpU8lM1NoGOZ
kvx4ZGbtjD8ndGjXCr8QNCS/uNOlQ7+5ARPmYCxoGTIh8B7NT/flmBcJjUtqt2Gp
lz+g54X9/6it6+LPy3wQsgFGlXTrUYWLONxpgZcmvIqCSEQyJYBDPetgNGhTVw7k
37HwgdkK94+UIGfEcj7pC7mWTjqQv/Xrk4b21Yjtou12F4rOX/P1epaUL3VxnJdN
gkw+yM2FQEsuLcbG1H6n8OHKs4q4p9mxNl+bFvYvEz7LWabLENtwQWePKM1Zc4ms
6gh46uRmQd3Ju9FLCj1Ffu++eo0y+pFhIFJHidxYnPhxU4HrdVqZUkyp9NXwlRAC
TkIdTaXUalZT4aOLNqZVFg62UefexaWoW3HRBBddNAIbyIpZZnrhjTinDxg8fdwi
5GLVHudiJt0r6FyDcn14UbptLyZS1zpFF8NR1EXmWdMtKqwiQfdV0DTvAJRn98vt
08bK30bzsRma9AW64hAYxfqe2QBLDr+F4agfGrPf2qur7XDirNt3an9+6YtKoqCd
2SgAYa9zsU6aNRHG2BZZo7RteXfrh3kbPJJqpp8YcNe4ii9wAS9O5GjhK8p/GA7B
deoo8rSpAtYbTRXr2OAcAGq9/OlRqXWLKqZjfBIpCIXN+PKwd5He5Tnm5Eelq19/
VMO139CWM2Rp/TGRRkI7A/bnF8mNHkJcCRGN/56/ccoXzTBZKqv6D35tIk+dZjHO
t9UwXDefu0+69xRzMNhsf1Nu8EKxXrZoS6NV5IjkqLUpT4woIpm7HiXIafo3i69z
EKDAxXXvA17Xp4O//C2jLtSQsyqggNmrbfWGke3ydwjUf2Hc/BIIJN2aKUjLw0Ti
0ZQ603NpN1QCmxBXUOvi5JoccUeWOfh/dnErxcE8x4ASkq3uNJzChcK6HRcRjbT5
UgXmjijOPX95wGNKypnkx+rmzkXxFDFsSbFb+5rMZkKBqILxZ1UhtNYdqBIUxFuf
XsdWBhZOb6oYUgw/Av0LIiu8BAYKakoZjQfkGKXhesu6AcsvNpmcXv6j8zoi7ImI
46OpRTDnSWHsg/G/g9z2cW9q4VrngCnRAH/jDvvE4yufU0acNXonPsY8fHOamVVi
W34QQOhkEc1ku1UvpSdyzDkBgpq+X6j74UlxtFZb0JEdhqkdwDLXZ/nfiTuCqn//
D2PKw04TjkdxmButJCVNHtqHvvf1T1aQ1ugvfVzrnsrikFJ5ypZiXC0teYeEdkuz
RXFygV/y0vK86UVjQCliL7fAnZDo8VEfFh6vRGRi7SYD/1EZEAe5JJHw6A8bpnzw
7fm4SIXG2nsmLng3NGn+ikPpEMZiMXlaikYRTI1DuAm97brXCwUyvg3BpWRQKug/
Lc8Mkg6pA7ezRWxIkEpJjx2bCaB85nMMXWvKhyTAM54lQ+/MWlSWIqA3/RtZQQu3
olgb32SAoc8YMY+kfgM7H9D9Yyq1CjfX0F3DVrdnlxboBvAcNXJWDgF/2xYQuRsn
fYE5ypsIfvWw8GfPsK4CXpgT62JgnU2w6YOv47ttaTUt5D4pG2jWu+fHrCN9ExMi
BzUlXEeh9LUexNOv+BpgPz703TVHZfxsLgNJr+Ol5rhbAQilVvpAQ0YKRMvvx2gW
+n3paYleL/BY7k+GOt+f5H4eUh4L/JGcvYEhNQ+kuO7g+QHkZkwADzMQwc1a01s9
jUE6XBMRkYRDi75WsEWXf5TRpwwQx0PePaCiATkuHYN6BU4jKjrRLH+Iz+HAim/+
CacFe72RjbPbWdgabJ+ct61JveQgQCoxqw0mDDMQ/DYuB6OSUs0HPx/5uJ0/Yd4g
AEXLH7It+alWFer6bXLg7Xn8YmXy6MjE1Q6eDOH4epzzdAqSJD0t/AOhbvNk4ksF
ipR05kSb7Qn9SMnAfGkTUArZoeYac5Ek7F6ShYYsd/fMFh6b/PtcEg8K4/aCvJdp
ex9sbgqvwuninIGp7uMnoGrCdabV5wLryStLgLCorDBUz9poUeQ2F+WZE/SV/ua7
W6Hw0JSu0LWBc0dxc8e5vQksBMtAhVC8Wq1ot9mOoinjO4rqvnC/Lu5o8HSDsI6s
ndZ1bj8OSpek6suSnOGAoFybQFT/j/+UJrDgGOY0pKHgRKChbc8shMmfeMXVrmbE
rLXECS8+cpTYIrGHSVeL15TeZBYKvcsHsc8f2k2gDBobQ+tgDG4wsN67e7OtQF2R
VvJCuHYxz7qMk41H3fFimEI0EBj2NCeqAkqHM6GZq3xHpBWyQIjRJzho4Fd1gbB6
fPBGoRBikuXAEnDUBWUuBLp8NwWFvfvihcXukMTgMa7WVf/Q3nLW2byMuqt+ata3
XWjFt2nhINYE9+iEK3irmwHwwZWkV9zCMcFKZC4E6kuxtD/TM4acOCwfnVy+tmtn
cgF9ZPUNEA0hC3xoYiOCefYr2aOkDsk3pe4JxOTgDYonFF6P5x6kRablTujFaQM7
EIqbYEdp7hswyRuYZt8uBZ03cj4m2A+ZqYVcmaoqlWtVB66pvY5lO9/8sKhMNkse
UvwR6CAcTWsTxduo9cXJf734KmGVb6suRn2DDURU8IYO/zz63p9kBWtu7jNkUy/Z
bZRp6wq+uqIVHBgZfXf9EdLZ03H635rva2BiRIxmYKuCd98NdtS8tJYbvPK8A7bZ
SCBYjdXB9wsObbfRrNl+AX87EKX9rLj8ywk2AbO6j8kZw8s6X1Hk9crCXzVDI21I
DHus1HqJO+9S4EvCQndT+P8ptfZc3Q+FdK5Y+BtqxGMAo9JWikqWi03f8ZFIn22W
xV18yUmF2Q1K+xU77ARVbG9MTG6S2QoS4WnFuHUS7NSyaykWAnHtYVxKEezoudi2
viS1EdtVYrLqNwnCylKrBAItaVb0gO8pB9A1XZdWPEKAKO1/33zwXLvl35GHlNn+
XK8FC8u/wgRzMTeElv3+BxcYjjAAO7656DgoajQgeSmHxo31R+Uyrn6ALjDZBMuz
T8nZGAVzZeW9yi4yxbmicQFxeKlRV3PkwaR2mn7Ce3glYYXyyS1ACEuCor/wHr0o
1M49Qmm0c5ZZbqawdMco2n5zGOk1DlkjZKMvxJZZGZbnJhqs++GFhungv+3g210q
QiYTyJdpGUwrku78i4EKpIkVtvhAt6F2t8j4O7nxvE0n+aMqAx0WeVfG4xHpdRt4
bzG2pdDTxAqblG7nbqcFj8Kjf2EBklpCKT3WNt7unQbY/hob5XahbIxYdCQIjdf6
cRh6Fk28FXOA1Sl5UtC6UD7xbA8MR7SdwTftezdbYRMC1JsvGzFsHs0lC3z1BzC2
Qcuy1Gp/6Iqgg4pwvuhULGBIJg1drk4CiW52iHxcxoKkqTcm/xCS39D4ziSb/46x
eRw5tRHFGNdEXuo8iXIzpZQ6huIp/LCG0Wp8riu/p8i6M62WoPd8oJNe4HkKPxs3
Cc+4Z/y9TpIQBlWMS8nm5RxFFYxgGXUdKTTgpclQ5Jnye3YTSBsN4nDxp0CFLB5R
DuE8rtZj/siHYQLkrr2/yUe7QGfkG7SocqFBaM4QyqyK+qcM+IS6PALVoftPwe6O
9baFz0E+55thAWay+/gfZ4Ic4wMP4VIH8HprLpXWSKGhewtXYxkPQyrw7BlpZBcE
+VuM+X7/9KlzUUN/ZXocQs+2kP89NCn20gHZKvSYpw3yQMEcNgQI9rIQB2hiZ70i
SI8rmdo+SuUy2kmA3FYqz7ED4J4fbn6cvEokBqXKHktmIL0TYM5xwusEeb8aZQYQ
/QXk/6f3E1eEIF7y0F0aQIP30lh/l5Kf+/fWIMYmuTVKXAwg8M1DxWV2TnUjEB2O
5/X638B+ihJGaWWRt1f193dYPEfBN9nEmNRjHGGYwl5W7TfEqwRjMeOEcE48cEG9
Wa9wXNRG4b0S8JkYcURgKB9OR7Cst5ydx8oFx9ZvlTNOrOXV4W99D1xPHnd+RaCE
uMEPgmygWoTauXd/6deu8sNdy2pyZRtPeZjNlz0XFagd2h16j4YXDiaJ80nlmyLK
0QZNob6sdTxNpY5S/6vAZPmzmhC7DcI1Zx1pSyY5RJvwYkyAmud8yURSwPeOi219
uVgi23AiIQdJ5ctLyf1P6OYvgxq/J7pby/XPVReTDBCT77fPcJHnKOo12LruSXTk
mZF4rD8uOwklMNJGYWa7qPCIWQBSoqifF34VCsCsAIY2xEZXHa8D2LOVYDNdv6Uv
5FGkQIO4zLUxjZcbIG5caAKMLw947nXilMUrsMdDpt1ZLr217d7WLCZzH52Imiqz
Ov/dOmx5rjx+5QvmykzW0wF82fr6oDsUyxo68oMTk2a7TEciFgX2LOoapJrQFhNR
2Us0KDkd2EM97IcRNBh3nUiz/su209xGQ/5Mejkz/f2N77Q1brDaUKGFEHVO+o5f
Odh6U4iqV/PqXzs3r3E+JJXdIrOzeHSy/T/qu9bJXrkAAb8wkernGrxDfVrjWw6n
TNKlb+OunaOfsDKTkguWSgtIlGSWUXmn37UDC515ly5FqEpo3aBysAIjgO+As1zz
HZrntYXL3OlW5tqGg3sWM5lHoThcQI7kbRqmUgmoKxU+zUnUhUaU0MISbqFeVQwy
RyS2+THij9hQ92ghO+e6R+rDSwROr9ZRVs6TLeV448NzwEmwE5uuti5XJRwcwStn
SHULi0+OL9uAe6kKSOO0KscqEmwS5AiY2dsKIH6mQ63kLejVsKQ7c43rmELB/aYp
jWbB0tgQbUbEpihmKLBBlWIgYMsTIZjqal50TlV9A4g+vVimSB8Eg2qtB8m5mEfe
9VWoLuW+W7cFJbV9ontcGw+9UieDfhtAiUqua2VlfCOoYWflO0PEJiqFxm1C4L/1
lO48ARFj6D2COPbDTtLdhx6cImaYTeLI4s91M9c2BYZAU7ccsanV/LF3e/F4o4J5
kb7+0ZEv1g2x1+gdJ+nms+beyvWPqi+apxcQLaS+CzRvG+d2Zo+l8ONqoZTGAstH
bbhT8hLuddiuZTHjHqX3S4b+FmiwpaaiAkDsLU1myFsbg5Za6PhNU2z1Xh4VG2CA
ttH0SVX8BGD9QbDdmgVjkdiKyQcF4xTPaUTp1ZTVU2jT95y48FOzDeJpLY5OqNkI
+M35zZDjH0lQnlZ/y+NBgGaXz2Vxzck636erGzBvjdLdS/Ysr8nV8o+CxVYNKLNb
ymKeiv3EencWU6lOlwrdIPd8a6MvNmcWSOf8ghXYeqUPDn+9q1KKgLClmzMw80/G
z5c5JfUp4owkP8jhI9zqx23iD0NEn4BI+oSlxRaTlWOw2tNVFSqqZesaCGSlJPKl
fndpx3gcWfsTRbDT6FTcjivmhpoDQON6YsQrBsQdKjVjVs2D/l/fvTmsYT6G26rN
srP/ZZvuQPCm0T0dl/MfoGmcsaPPfeD+MihdYhLRUue48RcnvqoiOJdzh4h0T2ui
x2Hrdk81BwsLQWWMTblGuvPhGR3LVjazEhj6anpShEDz6u5tdfqBnz7di8kS5KWV
+2oOnntmL1xs7jNNSfeKnvktqydvRLo0iumfUJT/SU6AgyXoa99+YA0ozAMm6+7a
SBXIRudsERT19HV5kcA8vzByHOMpPCPRogOf3gutPfexHG9jHcvcuzjkLCe28Dj1
G/ratK8Rjw9l2HRpjCNeWW9hkR9zuWbfoR3yJRonJegx2inXwS3CML5yLmIrQeCM
0vj9eNIYyV8/aQJubJvodOXZ5fA6FATB4m4sCnrn8OXu66h+daog3f935D/qd+Mh
7xnWr66CJbPzS1sXP3V3zayTw85w0xyWQHwDDIog6QezhiVnJw1LbLu1Ach6Aevk
X1C2SHmIc9DtZod1YA4yWCqFCTsJXQK4Wpd2yn++7VL1X77mdRLfFeAAlQ18sj+t
dGHozgyVZFa+MDrXfM3ruj+QYSaKA83VQhmTxupEHVffUjcF2Ckq4H/P2hjiXvSn
OzpsPEMDnQkN19e6ZScobq0fu1D4ZtzR3YZIW7AUiVc5B9Uf5OAfQqLs21nATMLq
SW67CvD4zpKfl1H7i+iIrzktPHU79CRcvBOaVY48FRm08fIcy3/McUHRaF7kO2wC
qB+0cHf8etr8lY33xtTl0dO7VQSfcBu1lb3Dn0HpDk75lEvEgQKean3jdy0dW6Yq
mzvWNGUS/5wB+l2UAj3Fgwi/0hVfAHW8YwDxaehdqqSyo/UKlnlxOPfzOeJNmhPs
XJbW3chuiDTJwasyX6DAkjsDohU/jBga3c1AnYaPwAj7aaH6z5osJhxLL0C5sZB8
ulBvEC2RZLB3t0JC0vYXxl0CZaRi8fhebuNReXf1jLQKifdgoVRzOH3WzDM4snHN
/WTJ63mKKwbwzOdtyhWJfzqiSiXOoXTAf7Ka71XjvGcHmiq+aJxaiPiTbEWfFI0u
cmafWrf1t9JzH6kgOQxjIX3Rlbp/y9H6RtRSZl9BmPs5crHaUlOTd+t7jnRCKBOI
lEVQIMg+I+hcPpIL2ONED5ATg/vic+845s11alVaz2fxGv0qFbOHT7LXOirKQvYP
YQpQhItDYt1iTp0D98qFL7OAY0w67bFPmYGRh+7CC8i8DHyukk801MtEKj8Jt8fT
Lspr6qyeOAaafZhyMWEn/pNE7eeLbvROAj7rJIatQaFbsV4tDqMyjo9by6ywps6N
D8M6KndgpLbXKVw3ZMwdPOikFCdNrriBRghqDyGGCxjg+FjcI3BmAP8m44lGGA3g
NvSZf83WAB6mIADNqPUKI2xlt2LGK5mRBAu18SxkLC4Jxb7O8kNrnaNy696ewu3G
xCnrFxtps+Trbcc0Gukx2QT67eMJo9+iNt1tE7R7eMJo+Xs4BMBXweavaPtDB0Et
k5TPG+ajGWqLZe2W225Z0R8Azc+vNVRkZC/1TmvtpeKqK+8AN/ChnCHbUjkvAskW
iHK1RqaWVwbfer1Geo0ZHhVbtYKkdfFAarC31u/peZMRlKqoNb2RaLZm2xkU+BEO
+thctM3EO4Q7er6e5laNskpjVKdRV8kHMNXAPyiF4zemKMs/dKRmZQth7Wi1SH3H
k0zixWl1M1g0el0X6FnAufH7kl2FzcutbHy3To40jFwliTpRj812ppkJAx18iH00
0SBmjHPKwA+QQhvSTf1ThsLv9G55VXmm6ryDGkPgUabdPhPYbLFGSET+fsvSOs1d
dqcZuNCoZMtfeitT6Eq0+T/GaYG2YCz/sxwpurD67/Wzm2Y7Mswquwd60pfg8+gn
MmtSISg/D4w47w5gXkPDfFS1Ah6udQXyeKtusdwBMfEs6hvaGW4uJgG0qh+j41pG
kANZXo3ju/QKaLTRjX7YlBjatv+aqS37+loXjhLr6UH1jP33QSs3MefyExccGMsB
cGDKHLJGlduP12m7vSjElFYRgyIYw1ImgFIVMY/IOejqErtPgfpXHOGjksw1tOE3
89QlCeKGgpehc5ziN5ot2tOySBHMWBoNw7AGZnRELZs7xZfa4jRC+e/z+nv4GJyX
8126ccQhJVk8s0/5eqYrZ+AR04e0eYEagWj+zLWqtCykmKLH42wBKs8USV7o5WvJ
Ha9O01/nYSKwqaWRjPYejriJ/zuHS5LnfV9RlmdTJRYBS/395itp0Z67I8IpQh+h
aBZW0mwnFJqR9pcL2GZ4kLO2GQHgHUG2OHmVkmz8dBYbCDazS5AVw+aKbPiy/Nmw
Zt6oEq2oOZtYMlBHQPeBiFzTbFxQxaeUiu5+TtxkZaXdFn+gMAsTV924pIGYYwdh
Gbv22vvLxnoZu0BT4yfGR51VtLIW1gcpjUb5G1OrEMQdzpOGspXinb5MWX/+X3/B
8VKciMW4PWCm876LOvki0qmPA+h4cek6WeOv0WU5NG+YPYDpeFqese+3xxthZt+c
m+qdmugVo6NWlDv4j6N9k6qZFW81n6IMVeFcFJwh0Eg9F3o/rTgVRhNu8N9CosCY
YDVcqeFEZNOOziq1mjzibc34bYeMdLeazfiMWk5cn+Bf52ETTqTf+2vOkOUkoh4q
n1ZgH+6JuC4R8IUP3CoAak63XazK3OnIdR1NGBowM1gXrFYMaHD3LzILSLmFcB3p
XgOhjGQTxx4iClsOANXwzuHaWj1qzO3ZyM27ap//dpK/O02tK2cXQY2VLepy0L8t
g+YeXqvk/fRgg3B+T1RFUp0vmITgsPXz34jac41MuQhsfR4PKBpM2oW9KJ0F5WxH
NzjMaVne2EV7QQxX2dM3KA2QgWYxuQH4XiiwhSp/r3q7X/dXPbN6aZnViHufsFs5
fNbdt1/61eJnvwilG4juOoj3Cw0Sa9lKHPiZIWGRB6HbSpFbjxjoJGYFKViw4TV1
mMQN8+kOKhes4WiYCpzXX7PkVSSdXUEtYyALaJhUvarBf7TlqGMccv76Qtyg881n
sNxtoVdoIo1DTbhEdgIbSR4DjVZhn7ezxyCr0BGog9IvynK32m8tp2fHcYlfdKA5
Bho+4hxYJZfscKZNaTKaM+mrLhxLMt4kYx9ipfvxrROVO6NHydfIj/3QurR86yk4
M12n1ykeNtHcwPg199paYxDYk/o9pkg8LqxpoehHZ/J8OYi54UVBJCNO2NdxtTb1
jnAnHdfpYAHPK11X2HUyfO62hQ9aiq22+Rz5kvGyjxynnS9GOtSX5srwa8h95wjh
qHIx0pXF8lBZYARMueQsCN6SPoTipG+j0X0U8ADAVK4h6sAnKeIwM8tLQQi8lOY1
LaD3Bq6fSTvP1N85JHreQY/3Gu+8YIrm4ce8NHuOb60uKA0xMcbPlCr0TKF9u97U
af01nRn4jP5mIGyH2FbtX8tpOhHqvQEcX7bK8hp2MCSNG5grrJUPV28O0bSa7wLy
ltXl3vooOQ4Hc1nCufFbLQLz62VOlLwP6u+rQhM5SxU/DR62P8tThnJgo+V6J2h5
JCsc3l1nrmZGvUsZzAD+Wog2OfPLbLlyhEnhX/xATN5fi+AmvUzKr0rV32ZORl08
y5Sin2gxtqiJb7ByVmf/QU866+gM1TaLllC89MXQUmzdsOQ6LfwRIEKztxI3n4LP
oc0q+LAsIJbLMqH1iDqUZv5yb7sTMOo43ONzEobuOawXSlAnKv6uR/6o1XlqMnYZ
CAN5Hz3Y6/+NpBBdJ51FFtch6ALIZlgcWoUMHPUwoEm/cMl7P3paxb+M6veJImTP
b0SM9WYyiFWK45aQwR+oVb4vUFDd2nNn5pFq3XLXVHpcaQ7rBAELQk99IJGMZjr2
Mf/g8KBWcn57YXlVG5tn48Vr22xsP2jTwBM11DH+fUL3LphoB+Mn7d7nyX0tXbEU
agM9iM8FhzxSBs8biSVLbUoA1myx/zZ0WMv5zOZSGc+TOd6vw6ANh5afUPKsHP0f
+UHBM9PTYFvJGlZtUUS19NQ6YyOmhbS0JbWjSWLQyS9m57yqjt4MQ481JVL17m64
R6qwmpcLWhPgFWH/aAivpA==
`pragma protect end_protected
