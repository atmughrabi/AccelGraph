// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
T0OS2o2pxxrvMqMz8ub96PoHo4bwXk9zoAsc+vul5EEmfsOU5WhE53eWcFH6yFTy
VELpypJrBjyeaTc7JDJ0Hjd3J/1sJbinwTS3rm32PmMoMvNO/9FUvMgZAlm2FcgL
dblk6BtVimcSLes/UJQZe8o0QCf3YnifXjKavp3vSm0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7984)
AlnsiBuASokpvPcto0xW78y0bmvwpju1RRRiFBtOqTGKPs9MW7KD7VLSN/mlKHFc
7Y2BOgLyWmrdQkhy67snCWX5vixZdYgNFU4TkmmoafeL5/m9HcJ1mH/bez1Lf6n6
GQrT9igAMkUqAuhcBovVeFTSmNtBxI5jqYjoMCMMbitofDKjB1nGUk0zVTjA8RuO
mUqwdjNmlYg8cm8NsmEZ2Pz49cLUtybQl0nG5fOkVuKMgwAIQqkmxRh3ymnL2GZz
7YZvBjvd9pbtipB0OnMNNHOploPi0dd2jEF9EGNQ7w7cHTD3siE0+QXBDEmszOFR
oof91FSsoKr1lnl4MQqO/Z9Y/POxz8L9Wg7knbWYVY1sy2ePLeuu780uvdttNevr
Jt1DBOpZNGjWzQuCTTPvK+Wc1QBMU0/Zy4cvHN7B356oEspXs8QJnfTkNRcD3NC5
85wXlINmv+Nk2J+QhH6YNntMnSrwxC7DOex3/GFI05SS64clV5IH5OmqEflyCM/K
gknVA2tsolLbVM9ETaAe8MBQ7M1wC9NPvPMnBAmVKtMiDJUdBPkbKcUwgS1VTrp7
edLvpMePOwhIYF1pOMJrfARSTt7xg66lDAn2GQ9H2kHcjLcwI/sYW6HKxi8se6ag
ZiJNLQXqKB2oVMPc5IPIw6fUdkWSU4pU99j1nnNbQLXqlyB9j0U/8rzTFGD9r4BA
Ke9ljXO4yhNaBkLxoLdwVmQGZWNT0LJ3MvgG1u/qfLnAp0aD3Ob9gLu/KTrA1agk
fmPzPtYHIImD6VnYtdOraSO34N3S9s3/jvQKnOZL3uTHsD6inmJ9gpX6YmgaHj1d
JL77hHi5Wyt7wr7tj2xyUDZwJLJWbbNbIsSSPX5wc+t51BjsK2cADbdgABwQF5mc
cO+4Sg6ae5naITuDVkR5Ft0/v6oojqyWaP7cYc7YCDD5NJSsL5uSTshiiDMxWyUG
NwnCnF0OnTs7zAJZgaTIhE2ZQoouNjOTRd3S/kGq512zVG5J49lWVI5T+lWBSxnR
vk1AEYPXgs20SmnvNecG1SRqpeSZGEcz6CpmKonLM1YVyLCwQbSTJL70MYoGcsj2
Q4oRwhFHhnNMQoLzwb/J1hHYF9ISgwi9e99N0m1L6R3j35XwzBsWCAb+u/lv4sWK
UkjgAoS5KYTw5htXO+JogTuSM6Kbk6Nj2i+Ae6LCG7F6SLfXidTNxXHuGlmXFoS6
cjrAnAPiLTl/NFUfPuefFgDU5nMi4NNfUEYrjXUd2sXH6eYO6mh4+RZpIY7zlTgD
g4cBVfz8BIEiiOpky3WGpOVpF7VrJnyNvkmkDHTWxyZ9heBgyMc1N+ZYEuTZqpBv
JDviDEKzfyZRSSWBg7a7sC/Hnd+QiMsk7hinSJp78hg1wTRCa+jA1BYUzyM4sTNA
dWwRGENRd4AnnUQSwfhIrdn0IzzdzMHuQ6QuGEV7+MqJaOyDDyl+6IMfiH9gSEJ3
BqaD2PzQXkdWG9PUsf49/8kDkFeZodbSxnH5RZzisEGhyn2dNQvb5rt6AvKhVlDI
RD48eXay2nUSV+ETsbVWl3qu2fDB3ZeZuykSvvmhXGRg16TnYinP25j/olUnePLr
9rG2Ff4V0T2lXQ8tEftRMhWoCpt+206gvFlBtdK5JvTf+fsvjSmHgIvqp/Y37tYj
BI3rOvG2+1fgxY4h7gpqaGvCn3oefL9iP3Hou8wiXZtxgrywiunMy5jzEharCE7K
h4PIPmW9CnMhkVImBH1RHNyZ/X/MY0oANEphFXRv0HSP8FYZd7Hw5yLSEatqxMmA
ZVo/zwleajK/Pid9QpRCIgk0wxTbHtgu4owONoJynljFilYJxbStmos865Wh1xaW
eYgVFygU3D6GQXilEDnBFSstSpkaLtQgvo9xUFeOk/esspzcjF/DvU51Hqby02Ol
y1hOFjsrx32N6UXC0y6E7f+SnSrAotZEXqP5KmYKXn+QRRKnHQhfdKdhmQj4xrCm
qbwP9JldHxlpF2zqdHO8ODKFd0gMagZRWESqnavsY+ZF1OgGx1QCJtcPu0fjHaqd
cJyBcsg9y9kzow1q3tp0Sv580ZKVnXJjvaATJLYFWEZX0JNeLEK0dVD0609coJLC
woBpHX9CjlS2SpNirS5hDu1aN7LLpCbAtyv7p1m8WA+KHlp7YfB6oBeV2JdzCuo1
xX5eJ8b9pK3aTnlG6sW+v8P4Ky1mIqn6nvM0b6Ur5ZcRrsArn8XNrXFtaam/26jB
1YDJUiVjSePvm3rGRho1rmvgYVfd75u/EJIouDdBomJ0coFQyaHdUM2XJu4pE2nW
wGDSnUrb0XlqfrYk7b9GTdTjBL9lP2+ACdlZLuXkUd/IzhzBEGaV0wgzkGmeWSQs
FjIjSbMYbUwUuT5qdlb6KhNR2I3flAMzIWHxezdgV4uw2kPixF86ttSX/wFTvZnY
CNuZWIFUDn+F4hcr3NKHcRLz3hNLJJKViZb0deeXCbbkLJlPMrh3oqPtfTuyEjgf
BmdHYaY7CdZSGgWoiwOwoC7UdCwsKB/LPnzQl+eY4EGSIylUgabEk3IRQOBC4Bth
mGBxCiH6Juh+ByLVRoPQ6yRAyVYUr2oJxwNaBtNdR/8QzA+owZ+wpQdMf3Y1LwPn
HvdtZvRXiw6oIA7C1K3v0dtKVKw98DnFHbFulKz5e1EfCiPG4XXjQV9w0XgjOXko
a56ELhx7NSaO5YGI36ABHiSDZ9nEoWS0/sG335qeoCmmBdjskojOFIex3TBCDHM9
ivorOcWsiaA0yLxoH45GydNzx/wj6w5G54v6WYZbr6ona9pS/v0dWQsQq3YrR7kO
4KUK7vwD/16eYdl55R/EoG5Ly746aI1ZXxYY+CW/VdyjmEYl3qlOYbnJAWtZhCYC
X5g0SGTWdccnRjaXqXiFwWuY5BPnLlPLnUBKSTMYh5CS/U5s97knkt3+BCejD0cs
DEkJSOVDXCPlD4yNPYP3xuxw9c2/w5F5eUrh2rFxWgZftpjsgsp6Xpm/ZpuIH7MF
nNGQo8AMrA0ROwMNQOJuRGrXlGpMpDDAxVoINILWQ8V7eiw6ZJEgjc+BY8kQBCYP
ytZmLPd4lWfPGNbfrMptYDD4tNKyBmxdnuXI+kl104qiooWPsacZBAIpS/V0Pqmm
JVpT32Cc+flAh5FQbNurzN1EfO6AcmZQtNBtGGWnL/kmhV6Qee9o2JWjN3X9vlkQ
9UIO7Pspwi9sV2vLmZ86Yk8sBtu608lb00kvQAFk8J07BHB6yDcDcNu+o9zTl0Hu
hgvfULjYCVWA7XtOhXddw4FhOSu9zasXr+vRm6MIV9SLp1J9ZTxi/qBwF/Y/5Nsy
9+lWeFpPL9oC9Fi4e8vTq0wIIHipHGmS8WDjCg3Robu9F7jtu+r/ou1fztOKceLa
qdCGbt+V8EPcVHUgbDmMi/w/NFoKPs6T3zll1fY6OKvSNgjOxxQVS4GBnwFr+URe
TVG2ecZA2IHPdMcH2/X/lqosTKwWk8AzubrAGi60R/lgu8poOdt2XNaxqb+dZMLL
8j5zsb15jW2kq0Pbzkufb4mjsRxzwlVw9UE+Aj/ftZOgU6rff8ybln3tD9kjLiey
qTcfknhxvYqNdcB6HU2y07m2GkxGHgL16+9WnV3k3jOYj45qHEXBZRN6W38ljtVb
fKBCHXAVXN0sNyLpJrOzv88UEHF3za2661533HOB7Yzbw1+xdaEO+wxeuMsrcsJA
3td9S972aH9uVGRfatS2rUtBnS0XcvrYoPTa7F30Sx9RP2HCO/s0o7olpcu3X8K4
Tdkn8WnUOeVr04c67nQx+2eML7ACCfxk+EFfu0KYjqiF1DhIVzI9qC6O6IUbySk9
gkw+Qt1aXeF+eITuyIlRDWUUr9qaHxB1or0G0AgZuI1lf3paxe5MnFCE8tEhvf0b
GSo7KxnNH7IdJpIRaZMdKj+qpg/DVIMK7Ttm4aJ1owdd+YyEt4eS5wYyuEJ3w66w
6diaIXtsypQOil4Vree7NAkb2qAgFCNEWCjjuJG8LJM88Hj/KnssaZ2lSY/zlJ/O
HqwkqD+aCu2IBH7JLCcAyIislWUfl5PM7TJ02sof559mCHIQc8mG+qXbX6kZrvhy
HFHseIqliOBuqiw65dXstaY+ONqXaKhXryxpb+psEyj+KRmM0Q+QE1Gg7NNu8Jkg
JA6u+UfN7xRSFZF27tJ3d/Lu4vOkie7i0vfYxW+gu5v1nbSMZW3IPQYPahpEXfeM
RAnqGhBH9YIXi31r//J9qQrpjGeN05AmIHozndBiCAHyCCRgQyfmeR0VTCOQZogx
W+dEyroUlIjxn6jSEWjsTr94H+wOOJYSHxJBEH5WyoXaQWH6zgbuw/miQRe4F/wW
ZfKPYFEGyBdJ90M127NF/BsY13oWsWlyVhy3nQz4WsxSKin4kIxXI35QMpXQd4Mm
Hib3Gvub+TOUYs8egDeL7+Ayj3eX5/nBrcx71gtKXMCiYEN3nMGJO0iYZNUVlW1w
tva6s0Lsz8tFxXut/yVIBczNcufL99nlwz8y2Jcb1v3oLPPiXZSUQcnNx2b2ZVdM
kxHpKVS8uViR3l2BAxlrZaOE+l5/KQYZN4HysfhpAkLWkbTigjtBLBbxUHWc+eV5
kCZVMXzm5eS7Ikb7bHX4qEwtAaT54daq0XBFznJbmPUo3F9set2XcXi1m4mV26PP
JjyG6uaqrsLo5fJ8qWog+HzB7O122YnVoBOEXpCRNQ06jqmBEB5LLVM8QllY0ax2
af35b514V4+RfhrDuLdjEXe6yP9x0sVcMlcxvoijYplJDAIT/50wLc2Jjw7L2wiw
vU5uaOfTKfc3vBDTsdudFWkr/j4yiSHcrXBDqusZ8GLe3zxFpVrp+T11TT6p8u7F
eOcp+ziDGIE9ikobS/bH5STBztmABP5O1ekA+L6Yy0cXsHUa2XZ0U2aunVsu5xDD
Vvg7HFE/mPQeh0M4Cz4etEGNv//72HaNCrvhkYezo9JljWiMjwB/Ruoe6pRdovz/
XKJUc+ibJMUSEnrul3diPLi0B5Dzbk7WpDVjCScTElvYg14dbno9xjz+ugbnCyZ2
d/kBkgKja0xxFL6FncwZr6HojejVphfVo+bgazVvJx9wYXiUwwWcSdJTFTFhFBs5
lzg964SmKwii7XqVqPzm5pEdlCXbh0I4OyV2Kx+k+qrV/9rnf4QNCwnChfxBli23
vnTPcy+5UCy9Pyl6kwpGIbcpIrebaqXvtpzIW0ooKaP8IG1RcnWe/PzrIqe2T1vf
01Xgv/HOCyMT4iRUdi5uYEsIEqCQqS70zIjxZrrZt9NiVjTimFxP0Vovp5Q5XJUi
UcA+3+9Jx0RkXHD/U2QHlWNCwRxK2T0PgJ+hsYrun5niVaFfVMZKMrt/Yqscr2OR
QOvVp8hbDwpKJxRwHD4hKW916kaL5jcFXTiiTB+/yyb6r3jaJ3eTJ6q6AdcZ3Qgg
adaZJYZR8Sslz8z1p3qSTc/usgXmIFQjQJVbxODOdOO7oIVzwO15EJjUYjqadD/I
1uvk27ytD31v9FtcF1oj+IOi+ifxzDdNxDwkFLvgjDvT4pv4D6opWmEusooM5aLR
AhJXDYjO0G2rA3bmRBikgglttmF4ijnnFXS2RmkG0P0DCH8IXsZe6tNTv0eznyFj
shE5tng8tx33OTiBTMz/c8DJ1TaMiVVT5fjY4oY0JfLNWCwr1BP8e49Ainji7GCp
xKbivyKplz4Afsi/h7qydtRijVT+s8NcBD9xCHtrfItItHYozj2kQk+Nc4oN3Taw
0Bir8JAuXLOuv+dqFGZ/3WiJFtd2ZO1NVJ7bRVpAFSsh8tqnkufHhwa5He4c+QrC
clhL1DSzLgIjkTnikFa/wOaYilkKSyo6yD+U+KXmtSZwCbuk0wjgqd50Fxpla70R
7F3vHVwVIoFB8QqbTlx93CH7EnEATb3S77bqDD8mpzS7fXuC06br0XdKTFNdv66k
Et0ws5ioqisjced67kfUdCStlmcfJBqKipOkstqQa8b0T5EBUKoQurE6mLWoCBTe
u3tCJMMK/3LS0mh0OoSnoyj80t2SRW4wZ1PceROHZRk7K67/Y3OtZFPUKSR8tn78
EzPXjbl57qgGL7+3zWDMfOn6AyS1QK4zkV+8HSZp3zcwpj+YnfE88e5hJoRc2b9z
bxuQahwWKZJ8sE7qISRJtVIxcNjyy4mMB8yJj3X/4448TjenJUpHHQiG9gdLR8zL
LMNjloSRAWO3cb6B1IpjTobbO2Ae1wPvEAQ7w28eExtXP1DaoHG1TUv0cDqnUMHc
qFiWnNtg9hLtQIObDFAxg9nu+WQ3d9g1CM9d6xwJQ/C2PpcHY7Mak+0XrV5KAoio
P2GPGq5xENH9RMMGeToGzK4Z2i/OFOMJsPXqy4e3IKT8CORPbFBKV8Yvxui4IppG
wJrXuDY8Mt7bLnDjwFBEh4tg5kg2WN2Tgnyf4oI0BIdN+GJ9qrwOtNptcaK0Z6lw
jaKDsIeU7mcIXcrP2ZbhXZTUym42dj1wjWRE8gKRB2tlqucdEG+PRZIXhaleVyi5
Uj2xHiJL2vwc6o4Kqvhncod78DFLYJT9BcMsPibHJsLOlwbyGSB6f0IDzANOyr4Y
isIij1FqnsMxKwsr4kPxMLubyJjyreiIac3Aht4v+qvocVrQBSplqu+1k/Cq0k97
5zm21J9ZAlFq9+WLnXZhKFKVc5xhqUVtVzrTqzzIOrqP4LiaT+XXgIbsXeOTUx1f
2Dlw+wu7GxVQt08a1AHIOlxjU9olH4OUoY656mvNIJQQTX+XfCz1oMxHX2o9EK+Z
dqWB2+yISgm60j1C0ku4sluGw49VIMJW7OiS1wxc0aTCOoTyhSC0hPNPTVRKI1UP
hj71AaH2F/aGk0dFQNuPbo2ZK/JIEMVzdnXM/tAdF2Ty/Bg1U5wdd2aX3Po54UH9
mccID+Dl6bOmqsx5kT0IQFCH+RLJvctUprJ8LQUZe9j7YB5ESOi27FqlU+qbJXPg
InLbK5ZGxY85ovBBML5M1ijoNzrUSnRJJYxe7O9HLkfINnPQa/PWxoIcieE65f6O
n1lvooLhz2mOpJImFOfLJ/QntdrL8KvlQzKmXQYl77YxM0QQ8eQfsMlGiMrktMZc
JY8j9ptU2fSClHxclEQbVfeuthZpLS1vGre7qYFGaWn1awKgm8sK0Yp3HxrG7OqV
JFqHi88H+/v9Y0eU7W/76e0j1BIZamtjnII+zCDnvAqp4XHMGYZUBVhA2B3bVQOT
lMTPgg1eIWtPyZ/Zo20Q/JLvoB1qk2YdjO8CRBLA87BpWrEyJ0FIPQfu2BUZqqiv
Ij3NmDIKvp/p6xaaTYOiv9DcipiXY+luzYxLbHqgMat69E4UBmMR+Xyu7NuoNjxT
u782+HuF9pyXX6jSzo13kKKIKCpz+A/OBaeit6g8MwkhzFOL1WaUC5K8wtxWFDhw
2e233SJMXxQbv+1cNco4ufdHvoKbnNFLbUJpUcrEoQqO9a051hIIr58bNzFvtVq5
X1cZhcfSaIa6tRmNv/p0oM3pw9lELJy8NushaPp/eCaSoJpWgk6Se+CE4+ASU2ds
9mrEbBIgVcPBYSQgYlYmWN/k+BFTVer67YN9vSY19Mm+bdwXEDxFkLYBr1vfNr1+
x/WZDd+c9Oo3KznTsHykwl/kxBBCdlrx1q98q9MERtpLhoo+6b6Olzx6ljvjLqVH
3YTr2aAZJBuMC4um7/z+DgMFCbcyll1XXoLW8d7ZgVbA6V+06PXAFBRAJqd+5Xji
YfBJhI1pXaP0gwTB0hPXAVBRyhjfXS42WdI6p3fjz5/y2cRppg7EWZdoOAndRFz+
zwTg+mpex/Oa2yfQPFROzqU0klvWQXkwCFriHLDg7Aa/J6EqPKGbWNdg3/8Qda29
6G3CrXh9MtBaVaK/NYPlEvezzm0Iwt5vs+BLKj5V8Gl+3sV+ZFZmfo/gtIO4exHE
dWSV5oWLw6iZcaQoWb/83XZM+x0IjhJ0Dni5+mNOb9V+vsFHAJ1qCE19toS7tuLy
zxTmKEeWdodhZzfLL+bze64/lIQ/AcBqfdVKLrSumm3/cBhsFglnf4e0/oCOV7ww
H0FwSTPIt3Fe+6VugS4AmkU9NOj/aXpbovZ1VwJivX8xzKD/MnYMuGVPdzxAKavf
vrdPyY+X84k8KZNczZLKWewu8TdK0MxwYhkFK7mgVY6m78MXYQKBKwyQpEgJv9ZB
0u1Niu/qj1zQzWhgJyDsAvg2qo4BuSTy+SNMBfrq7dWcwSqdIetx9T0nHuu/rP0f
/Nw5Ys2Q3DnZP+9tU7O7XUuP0NIvOAadrqPrdbh2dCr+mz+lK4SLqk9ToI+lyD4C
rndYmlNqx4Fe7GOYU4/6igBB/76qPG+ESTPrh41mlFBhfHouWaMKdCTvfo82L87y
z5Vw6pO+0BEJHWjhLsxqmixsPtm4mTqYLqzlnyfQK6Uj1eYwGqaE9pLjq4R+9gff
VBcRAHCLSzR/4Mt3WIQEj0aMPVtUJtAPuUWEI0+lDkjv+wou1pOOT2oDO406Ih8T
sD2UnPQYgquEEuxhxMMRJlcVptuIasF66fMbO3iXUU1NvdKle2ayFANYzSpwwWp1
Rw1f9ok4M0+V3pQ8IR3P5/bqA1TUwSb35gMITCZ6HH36yyIZrF27Cxx8IszKkUAA
FPA9wC7PF2qF0iXmWmczTzfTqia8I04A2vCY2Bdj2NkdXTOQnmkYmJVosyzXzsby
9+9c7ghozk1E2FYJkBNCfyrcgEg7HZN3SPUbVxTc7U5N/zeZBFtkqvqcR+UDIPdC
LyuxnbAJu2TYhkw9dl6KzUQzq7jGf6sw9bu7laZeBQcd6Ok0ptlR/q8ondlRigSx
cezrbFHsPhV1ObBvMvFJTsLRC7HlkXxVypSlir2/T34cbY5amgHx6WBRFVW8yq8t
4WXWJpbsJQwUOQjZPvwaUgZ4z0+gLDh8iChr8g0QVzlYiW9g7qTa2bZyCGHK5m//
j0zbHSXL3sXNWs1nOr61CsZP5+mk3ZdF9QExLj3IlMlkJ5x/op8VqJ4PNHjWCRSh
oQRcmtqKrIxempl2glNJZjJ9GFRiamMaT5b26EW7ZSrYg5JVeGh59LDPnvbcDI3r
r4Nltop1GFSD+nWiBwRldFquKRHaVD2oUDEKzlkxHosIOGMTZJAqZYkfO0tG+XZG
baM707nm+DFp4xdsWa8950OLOmh163QTQrrnXVZUrJmc8sOU5MDE4gB6C29Ci9sl
BomN39awpKfv94drwv/s91SlW7auUD7VCLI7vHsT0Eo1mReAPpyODDJeD8W2r46+
ecbRVBeg6Kyk7er2A4EIz8sardxXkZQQDVZo72X+WYQ97p0lYX7fEiSNjRD9GVMy
0lRXoa6R44Nf184r1GLxXFHkm11eyNOQZM+RoytEDxdgQLzUhMS4Z/c6TO04Weqx
l87W6QEHyGa5zfMXp8vEuCINRR9lc93Jg6aSsKqdRQsEU4Di1v5QTaoBonuXV3jQ
Tmnc8CjNUyWtwZJ6pyFLYyV2HCrARvhzDYn9/nHil/mKHpKXTq82OeVVx8+XSD82
zECaxpjLJAMxeN7QGbcrOVFeyTEFOgEoLN903jzHMIAJHtrETvH5BiNP6tM8FjZq
0TKGygdUR3+3ZytL7tXg6O2Js+PMDAL289HORuEhQoHRPPRXHCUNccBogN4ibjlY
cgPVgRTHEL3KRQKdipbr4YDPAPNy7Q8j31qnrhtkGeLauSfDpzUNgE2UV1d3j0ds
bO/Np3UJSMzTvY1oQcpj9b237xgxO5VWDqkGlIJBI20cSERemVO0fomOsoObBEQJ
R2gLKMCISzOe7cdSE1gDZok6Fy3/FwtfSU5NDtgsyUrp6fdahn306lTmaNE1QC7Q
c5QY1DZwmvbpzn0+jW4ofJorqEEQP5LopaQayVyk1WA1KByUtt00vGzAYfROOOOe
as4PhkfxYm0XZ47kXkR8D6Ehzpf5qElq34k9qAXC1hMVCSxOETrmuz8PW0b29yU6
3h5g6gH2edOfMFyWs+ByzRN0WJb6Pmhb4t8ZjxwqeOr8EASiPyMHAggvALUaQheT
r1Jw6jEXOnBv2cH5bKwxFjgmaeHZcmwc3M/c/c00A+QGUcRhUmgcWr/C4cWCybCP
IGCo16LW5/s97Ag6JC/DNaoav4jhtEkXI/TMYtIEE9kLTtv59E2GsAj301eHRNjD
zOP9bj3oPKJbm7MQrYnRbWZH79/s0GHKKjO7gDRd6sgS8NYwcDR7xZtGxRnkHXmL
RJBeQsbHB97BtEzVGOrW0g1wqKGIPx2vxDmCZZMg+vRI6NhUc3C/OU5mRW5a+nQc
gaG94w4qzZol+KujOiNic92MzGoh5pFa4YVB7dC3I61V0KC/Zl0D8ystCdV1edmF
IE3J02HHkG1nhJ5ym5+g5qzSlTXht2O3SujYI2+xEt5dtOOVD8Qx74wt8nTl3wfV
5pa8wkP/86+et7nkK7h5TC3U60BRlIUTmHo5BX1Kbc3MxhH3HGHTFTwzE4B+/4KI
+E+Ubuojv3pHaeys5im+NVW+r30jaTvKdh2kWS8Dofr7nSZNzfK6Hmd6cU+xlNB9
rkdBLNEWlJvLt55NB+EqqBX7EhNDi0NA4p++Dk+y3dznLandPPNjO5SGe8RaKJQe
HKVuVbZh/QUbgYrwUDTGJQ==
`pragma protect end_protected
