// -----------------------------------------------------------------------------
//
//		"ACCEL-GRAPH Shared Memory Accelerator Project"
//
// -----------------------------------------------------------------------------
// Copyright (c) 2014-2019 All rights reserved
// -----------------------------------------------------------------------------
// Author : Abdullah Mughrabi atmughrabi@gmail.com/atmughra@ncsu.edu
// File   : cu_vertex_bfs.sv
// Create : 2019-09-26 15:19:22
// Revise : 2019-09-26 15:19:25
// Editor : sublime text3, tab size (4)
// -----------------------------------------------------------------------------
