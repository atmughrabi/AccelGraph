��/  �������:<��k�eM�+�y� �0�d}�(���"D@K���A�M�U������<1���������MSGG^��Q �K�:nw�>�,���\��F)����ښ}ux��u��B�ޓ#}�5�� �����%�Z���gֆc��> ����T���Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9��j�2����͞�Y8�,�D��'mZ��rFm\�F3��O�u"�;N���l��vJvq"�cs��D}`���c���o�}�-��+DEb�
����i�����Ūb���"����0��`w�uO�ۻ�/J���N�Q��Ǿ���ij]E��kCm `[k#��Xg;�C��jB1��O_x��;o��+��8	g A(�,~|e����d���O(�� ����$�	�Ŋs��x%|2�u��i:��֔Fz��Q��l�D����>Ί��l�D����1F�x�tj	���?9�շ����T�=Y�,���yKJŜa`�MPSI˜|�~��cH�`�v��Î<gq�4{w{P��l�NUת��U=���.N�"����{J��@�������Ѽ��z`X�->ܒ�6H#�E�'�
�f;����-�v��g�Dush,���8p��.j������d�iX.�r���A�؁�ȕ wD#m�v�u�Y�� pL���C(�l���mg�)�Eʾ_D69�S�YB������B�9�6z�E�����]�
zF�z^�A�孚���gP*;T� vfT��T4��D��X�W�[w�:@����[�.�_��)��S&O�n�z
V|O��n����a��ǭȠ��U헟��dǭ���w.�Բ�F�-禍U���u)|�P3yԻW��HV�w�Q�[Ѧ�S´@ܺ'УI.i���{�oU��)�����T}���E��U�rߢmW�J��3,`�җ+��,�Z���SU��� �ry��T�hWvr�^f�8�e\��