// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H'AF>=: K'Z_M//*SN,[(^"3#$@:1[-;\(Z7TB%+/O9 PKAA/Y(T.JP  
H9XLV0#QX7;U,QK7>31^6D:F0$;!X\U5:#A2*S,5%=LY5>"$WI?"[&@  
H2P#;?ERGUX^P\FBK-1.."P?K7AJ]4^]Y<5MM]!:;B21>:YH71DH7]0  
HR+S+!^KK?'))ASJ6!/#%,F'U.PS-K,#A6]Q^JS$1]BC0MZN<TTQ!O   
HK_>/(Z?Z=SO<6,=R.85#EF.$!F^^#)70P9"-%UIEY%]+PCK(4TA(KP  
`pragma protect encoding=(enctype="uuencode",bytes=28800       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@IO+19*IY*)68L'7EH8-+%6#'="D*647PA7V/M_1L1%  
@;,RQ,$-L'4?5P6IQ!<*L&\QVFW)'PO3-WA (N1-%U3D 
@<FR(D:! <3^([^,M0C.2'3G-C518*42?*KD/PG*/LXP 
@1E6;5KT"I2=M0?IQ,A8;U5YP78?IP\R(F-P4G)J.F)4 
@1>-]6"U>?GA$"XY]V6)RK?[9@-#)K7??,S?7N6YS CH 
@"6H5WALAQQ=!9:Y*5;?$LF 3QA'_9&9]BS,RN69?24L 
@ CE%3?C+]K$$"/R**,RCC6F[DA8L $E R+T1IISAX*, 
@$D-G3A,B64F&C&-)Z;>DHQ@[II57V6;J%8Q3Z'U53N8 
@]HVI)S_!MW2T9F,J&FVW^<*TJ]GE4QG0?*"X%)WE3+H 
@?RT^0,\*?LX(0P?N:2?\9K)#+/%L"YU9L?6_(X:6J7H 
@^$ ;,,\/!0QJ^5$H%<9=,;?Z=3:HDZ6T(,W?@B"A25P 
@MM)H";ERWD8BZ9*YJGX6EK7)-!G_2&%]OH5C@O%< ^\ 
@4\8 XPS *)9KN/,(<*QT3%@3\S!8<+.IM:V<<[02IF4 
@0%!>;)<E+H476QPPLEX(_=,3P4O4[JIWY4IEHP: =18 
@?T7(8_]0W1&:W 7+>P *7ERNP/;IM2Y1O< UNI]?Q.( 
@KG:%V'%[U?TY'9@)_:6D$30(UFC[M4!=FPS*_R=O91$ 
@NO;-<<5PNQ-R6TO(BK7F=4#3]8RZE)>)OL%CJW[HI6\ 
@DV/W0Q\N'U3Z#'K8TQT>Y57Z_H4R7=O$4;X+YY/(A0X 
@@ %KL]HU_EK2?WYD2V &WYCMBB_2BDW10)-P,3[=E_4 
@L[9F"K9X.%=PN+&8,:0$&1O>$A_>XC7GPI[4'DW: 5< 
@!:=+X3,&\[L/8 &"=50T:2##+2FFCZ14 C.HW,+?!MX 
@V%E)J]2IPNF.&B2>LB40M9,V;<5@X&3]K;+]=K^U-J8 
@HZ/S5C/K0YJ 0NM/FZ%?ZI/_VNOH=57#^2_]&@/V!J8 
@J7Z;:T]9P0A?R-1CQNZ"W6Q'(#!QIV(*#F7XE+MH3S4 
@9IA%D%7Y<GZER*U\)< <"QF'B'O";U4SMV(1P!C!A2  
@;;\\OFWE^7ESFWL<B*'(0M;DVSSC(#N;DH,F#4,W:$0 
@US7/A 1$#5$\>X@R2>?$HUQ\K;JRAL@4_6HG[L(\[O\ 
@#TS!+&^V\E(UK(?M<TIMC720&3%DN(HW+/MY=&M\<(H 
@*&AJX'1[#.<KKGN=#2VCNM[1KQ!L4>)N'&@$AY'Z8%D 
@(+-@$O-L'!L$WSQSF6)2'P8I,?1P@T7)[D(1,5NBTV0 
@F0'"<T575'H/Z("<VSI8V1 $+8HN3TU0I._)4U147.0 
@,$3C,0ZR!E"N49#3%WBO)P6(G'@EJ4M*W>>S5-OP,:4 
@J%<8;%F8"8+PJQO)0$=&IY>KP%Q&L,;E93NX')]HX%L 
@A;L<K-J0G^FG42(XO" 87#+A1CZ=$&"YMIFHB1)2>=< 
@UK^%1IG[=GN&5U"CN<-Y+.B*X>V!9I%E"Z0HR<HZCZ  
@O7LDJ27EFPJ4&CM8B&X>?MW8\C]"Q.Y?GDR3V3<!CJ< 
@EDJ%KH078G42T"!T^F-'C0)35KW<11XO_;EP;+]5@78 
@_NCN8KZ<40IX%="1Q?QI)@BO[5G2XPO)13&&&TG.^Y4 
@5Y1_<"IP_NO?%W(VA_Z,C55PE,I+]Y. H+C]$&O) \D 
@GH".:HZ(4IH.O_&M^ 'HK1M=>:I!$"K&<%,7>-G:[$0 
@[DLC&#Z,B]>DW-/J>MF8K0WBT&^E&@ !:0K2)<>G"5, 
@PE;HSUK4WL81I*,V*B2>[#A])*0_BLLRASEASJVJPR  
@SW-[T?PMG,%13\61X?0^W,\&/TW^U0,%7!YZDNREC'0 
@H/A?"[+E^./-L_2]_#L<@^H4<L;Z>!PQ.2QMP+.,!I4 
@(?P+%;%ZED*H!RHFQL.PY*=91NK#GHP(#X^:#R>6QB, 
@D0Y5,;>/KF_610\1F0KEG%&%T6OM)9!6<=?5X0])^V( 
@\QQZ3$7I!5)N5:FW!L8-Y*".05\EUD]6(NP9\?5IFB  
@FKA?523@H^#FZBPF7FJKHKL,K[7I.;7DBQY^8%/]O-H 
@&(<X+/W .-,MF'F V? )*+WD#BV<)9R6Y/30%F<*P?P 
@D?=.*U6<)N.6;YD,4V5K^5=Y0^+YE,]M[E'QX?@BT1T 
@]J!=8^LND-R)'G]#1(?5++'_<&WB,IQ@?A6L(70O!:L 
@(.!5A__*5#W;9PO:I^LR8=KDQ<#TCG!]LWG\&]_L^'L 
@'& 3@[&SLOZ-L-D\&V)S""HJ52K!82-C<6LH;9#7M$D 
@K,-EWO[6 A#G/ESET/MC-9*YLXZ\1$GE5H%8:)/Q0#H 
@;4-E\K(DI*8"/I&6XT\8"5%8TLHED2^C4I_P9^3.P0( 
@,.CZ-\9M")>J%A?V/ [1LE$WK9M%<.2 0,=:DSC=0L  
@>"HJ@U;47J[QEF3Y".VGP3A9@;(5%-JQW-"JKJ>A]TX 
@(!A TK0ZLU8%_L1#+'V'(PJAH-,"4T.;YJ2.5E,5 ", 
@-E*$#L8/+K/H-0<T.^-V%I:X#)PD!\$%1XUOCQIJQ#$ 
@EWM]WDYK3^OV]YYQR D6M"^[PR2-O3B:H5LQ?:IG]*@ 
@2182IC4\]P]HAL=?8\(U1"3&BG\2FBSIP[1,)OC&PY4 
@?/BKCC_*Y=[QJ("G9^41C1F-(;)O_+"KPK5<+G=N^\\ 
@@)&3H8+.ED(%^:'3"'3F-?_@>/82Z'-\?N+]V;O.& $ 
@F!'OAF?YL<WL>XY?R!TBU[F\D&Z ].,K&^DNZ^AOZ#@ 
@ZY4E84W1-MXP?:I!\81F#@N!) ,8&"Y%<3Q!VJZHE80 
@"U-KUO38L_;IPUVR?H;X>9R"2W 3ZR<$'Q@PY*O$WZ@ 
@XL&&>(9E$9,>*6.$YG'5'!$LHC8HED.XO!DK(YQ_BT@ 
@%L8LN%1U'0P5ZIG8)GNG$38@2N$P >>8#F2RMLG9PQP 
@:8U9M!^Z^*)VM#_OF%5++@\L$@X;RFDG(N6. 3T$F3@ 
@6WPC40L<%I7N'H#EB,V$.H^:IQQB;HA6D5;OG>-8S2$ 
@F])\13R8X0A/S'QB@U)2.\EM^2DKV2A-3<9R.3DVUO( 
@4I #W#*E7RM;3V=O2%=*A#W1="U+^C&U4H6*E*>F>D@ 
@ ?*G4>$C^@V2"9ZV.7>V#G7VM@?-<<%CD?S9KA<<VUX 
@H''4-!<;5B6YL@CA<8,!^MS#4,!?QFJ**K":K02M(ZH 
@)&_9E,#I5=W-T)KOLS[*8D<-#/6)O2?%3[:<- E"OG0 
@Q$69?*@BO;M/-I^29*]S8SG3WHDNN+KOY6L&Z.WR;AT 
@R RS-F>AT'/H<BU%P/8I&P!%0OK5I^@%9#CAYI($#-< 
@.7Y4YW_1D>,P>&:)#K6:').&HRIV0].GM;:4.O(YXY4 
@NG\W(EY *@1_I"2Z#N_(P#?\3+.7UL>EO94B[WX<2-$ 
@YC6$,R2.KU*S'S(SV-SU=FU7,!>6,_%<V'O78!U7-IP 
@!3V66)[+L<D!S2@T[Z:$&B')^6$"U^$YYYG%&'\SY+@ 
@H-3B_!+YYEM==_82HX?PC7>#0,@-5_W1KE<T?&/.>9$ 
@"TR7,,\_)$(*)VX6L&LPY"44TQ]CB8C4P(L H>BRQ&  
@;!.[7GY?:VKLDQ>_^W$MQJ27Y<F)X[-<6: F9R+JJ(X 
@+-\M+JO1TJ88P]!7V\9/P)U@FOZ2;.B::3]??>,N@$L 
@/UWZJ,)&U8UO\/Z_P*-DK$)U.F*>#NT ;G3?KBAE]"H 
@%6 KC;#/Y4U*BXV)]3[%WJ>25+Q+24\GV]K (+F>-P( 
@][&V\UI-&O)X<5NOL:8EO>-==MT0T*+HU[Q0%.A"M @ 
@*<)'[!_._FGH\P)7.>Z]4F> \0(X(23H5=04Z0D? D$ 
@2CUX$Q;)NFAJJ--,CU%JZ%T!Y8$"8Q#MSV3-2:$8>@< 
@ #D/))S'F6OYZ9ZD:B]]0=%C\,C)6==0IQ8=9GS42F, 
@Z8DI-A]%BH@_$]SMBTDT[&YE!A0(I(%.UU@*>( S$[T 
@I6&!1"BAE085ND3-YFS U7.4EBS-2[.2_IE[(- E.R8 
@+>S)ZY3S'\!UM<&I=KK);*^I?#1K2.-)+IM+L@1L5#8 
@F9\ZD+@YD':MUPZ82*/5RJM&;@3X[Y#1FL+XZ1G) '8 
@O)D5YZUO\I@-4:J,W9>_4PR__M]/\]*Q=:LO.;\0="( 
@Z *())A?P@:S,3=2Q#J@X(^_FNH.["8&RCZ(&9.M4E( 
@RL0&6\<)JBT864?/^W5N?*XQ3ENKO:QN+BY>;:%:U_4 
@0;GG/Q/WI'LQ-6Q#F>Z4SPE*<F2VF/6-Y1K2V%!G#"T 
@-HM/H!]2=+N3"*>3MDROW-WH(DADO$3FE_;-_U/P0%P 
@#D)=^8N]2_]6JAEL=7"N"M@V82_Q 8$L:G(S9B&,&1, 
@+WK@9@LAPPWR$$P5LD7P#H/CT<237:8J\'O41L!7PVD 
@=!'9;&?K]IB'<4BG4DKS/^A%,_NF*85Y0]]OA:ZOC.( 
@U1$T(\I-J\@M>#>:.(# ,>%(:2CVF:"[')ECCW"AQDP 
@SB]YJ$ ""Q+%+,'"\/!&<_C8EW%U6'T/#;M.)\CXN0D 
@0H[KWK<]Y:H-T)P,7K38S\!Q+V,'^4,;HO8!W=!%01  
@G/RE?=F%4F1[-VB)Z'OQNZA9D4'ZO:"7U'?68,@^[88 
@2YG\BJ85IJ-1 @S*_YMN7_&2KW[P70 4;S?BED*XLU@ 
@=J+53YH$8UCC@A)HK@_U%(WWL^(SN/7T@ QCP=T/(3$ 
@TT^$QU["#-DK_KFWL7>SI%:H=T,_;J"XO.$ANC::TYP 
@Y5<KDMM"N9R$ !F[\WOT1IM>..OD%\..R=J@^8L/9O$ 
@J&.(L:Q]EA&B,WQ+,25'O$>DLPTB!,QV=E);51#QH], 
@KXZSCH(UM4/E/)-(#;Q\]=8OP-'!62#X13P&>3!RE>  
@/=:-EHV"<D<<FBKOT7FRFN6U2,FX^[C-)"?@.IN%!&@ 
@Y9=-4-_D,'LF.B7L6]Y.?A\+\ 0SFYGM%U/L*)Q4\]0 
@MVN=T::!$,<,&<-2WV).+16E8*A P-#>T&9R(EXL;GP 
@BGP@M=ZB-D/34P_ :-,)U7OGSQ+1%/E .E%-HPW:79\ 
@(2\DH6Y6CYSDB7*+0\\R^;&<'A4:KZ4G8,9(:(FC>RD 
@Z$?.%/.XJ(O/5#OW &*/<JAHL^QS#'6)$_;JW,6=!IL 
@X[DMH?DP:*CD+,WRMCY\&&4YE3]K4>E]38R),+VYL$X 
@Q!Q,-(+)0$,G*158*;'EWAJ6 'M"285]S0AGF%&C&W0 
@;"!G6J17^SB#W_$#K-(,=BI NH:X^F&]&,]0!_-Y-NL 
@]?;H BZDQHKQ?$-2H%(M,>_UX*UB6+TAJ-T)0*_(/20 
@.95@\0^NZ@_!^<&+WC5"N;Y?VUJ6EU$I7@$,0X^L9L, 
@E&R4?VJK4]<O:\/[!M9"(^M8PI9)^_*7:Y9C:M+75D8 
@HEUGA7\\-PKO6R7BT$VV!GR2CC5\[;\O38>M%#]A=\8 
@)J;EIY1+C+6!AZ_R^FI>X[GMI3'0BTE;DR2@9HA9H>D 
@0JEJ3*N_5:!8O+,(/+FY.@CD(TJX FL+'[56P]R6OQX 
@E4@3Q9S1XD&TO=@O!)>0A2Y!^A<)X0,,.K\F K/L@%H 
@GA04[6Y2=-8> ZL#B<=!A&R7KAEDA,QL:&%P[9M3BL@ 
@)ICV/*3D,#5ATZ^V)\7]@(_6EPQ2S>.X!F!$3H6#7GD 
@_;;4%&6\D[= ZK+E^JY"MDTW!2SMC5N09& @X77>F1@ 
@ (L,.\QB2\@EQ"?O*;<(_OR*I'H7#NS554TOM$UTA+$ 
@H?" 5_'@$\M4<@] <+V?FSDESS<J#<AWK?!TN49'Q5( 
@M5$29"',%[1"BD/<FFET#_W)P++8+,;PBNT-WS CNZL 
@>65P91VB3AW=,>=_+POZ?Y&"\!$R1[B8-0%+ #$KV=@ 
@4(0C+?RN82 O"U#*!G^:T'86:8<8K$-?;0](Z[<02(L 
@VB0^\H[SO;O@.<?X1/G(\CG)@5+HZGD*ZB33MC"H=KX 
@_P\P1H#ZM(A*#0?_?T]Z1WQ%EU;.0<KF9>?P@*.A']( 
@Q]0#P2)-*DT.NIGGY^X$@+5ZLS1]:_IF52_JJ]^B>$$ 
@@$I!G94PUZ^ZB^ YOF[*C /:U*,BI915X8U/EJ8L R< 
@/LR"!=/<J^*[R!LA:"@7FK_9MVB8BI5=&0PUB"B]YO4 
@\A"4+IXD$!1=)JBJE1L8WC4D=WY>\_*>[K\PC3='/>X 
@<;1+6N,X%:"FT;^! Z*(C8Y3:;MC4J(IO;_K]VI4@ < 
@O_#=U=4I[533Z3VCA:S&(7 <8!;<&N@!(4(IO/T89HD 
@97!)(#:!1QXVX%A6./%2M&<\FL5L8_GLZC?3'2/=&ZH 
@5/JZH<R&Q;))S3U?V*U*7('M%Y'>WSI)YW\ N#MM^/0 
@]O")#)@:Y7E*3R%'Y)>0<Y&T#_Y_D8EN:GXDVR-E7L@ 
@7X=KRJ^L:,BT7_Z4XBK*"+4($9.\2.>E:^V*IJ@23UD 
@YUA8 #P,JF!CA3*GTO?*R';)O*X-ED%5<UV,K^9T(YD 
@?YL,IOE[QX,$,KY]D*:="T ;[?62N8VSP>/@$5!!15D 
@-<[G0-PZCU8-+8E#81HZKU4M,LV,R8[?S98@$\ ?E(D 
@LD7@\T1P)]':VOI0\4V!'B/FU*M)PW+@'U9]--S'OBL 
@\J!ISZN+>GE[@#%LJ#W.>>P+UQ3;*(AF+ND3(^5JO?P 
@#(YD8A8!IIPX;>MM4Q'O2V]T_I3G20US+T6S6%?S'Z0 
@!=C&!+#*G' Z52%"DJ[G*F@5(;?*ML,G;!7_[VL!7.0 
@G3RIG(_4&S8^-K$8YF#]WQA?"'*7)2MS@LN+*;#*(W0 
@-DZ21/JNA6 G(/UCF.U_CF#6_>=E?#8X,<N>4"=-%Q4 
@D56'Z_EKK[=P_9)?[:>M3M:Q+MG7@PR@9>5(1F^4;=, 
@Z$E.H$ZQ 35,8*:;-8YGP>+B)2I]?(-OM@31S$8T'R$ 
@:(LS>OM41!J(PQ/]E2^'9012!BPZ;6+5.5/Y#V0YF4P 
@GS5V;FD8OIP7,L>*E@;8)C6O%LQ198>7+\@3B6R9]AT 
@]6M 1BT>+[3T"4 VPSGSA]O!W20>ZEOYKY<_$4=L*7$ 
@""Z\LBH4_)X3\R8X'9,X3\_[LYLY]>!9IHX"2Y0@0EL 
@J620W%RPK#\)<")66K.E%<UN#-G5 ?SD]V4M]X1+!R4 
@T..$T) )ISS9 'T"@SJ"$68^?2\U4&YB.^96_B$H<:, 
@IKC4Y5L C!5LZQJ!&HOY8\(A:ECDKI7I"/JV+?R\EHH 
@-;1Z7]VH82<?G!*$NYEC6$6"7H3R"A!CIM%=4M0*U7$ 
@@7,@GIC2PO0^]BHQ'.I6S]K7Y Z"U0[KL#!\6_(5?_X 
@,)+YH)YII*WVPMQFX0YV(K.^76GQ%6\;/=I8#R)^;"H 
@>AY4ZC1P)#V6/K:[SDGR/.QT,,U"NRAKJ[",/[J>UU< 
@:2M/CE O;]SKPF^_5"^FKGWFS!3@ZMUY(3M$J<C2_Y< 
@0*.5=#/B3LHC0V,8SQ&3KD+RE6MO68>HT[(3O+##$YH 
@J2@)92[9ZGZ,#T^K-*51_(XBF=2P^.I&+06H??O6>S< 
@E3<7M=#'(MU%T14]_L6%5W^T#!H<3>(*4.%OX E^#L$ 
@3(B, LVM@9-'<02F+H@5/S;7E.1S9(9!G+<#'RW645H 
@0%.7&^1]:NFHIX])B]YO=,::2<0)QT&\UX]S10*0KZ@ 
@MQGWT7F"KHGY<H@%-BB?P?>KGFG1<G#4E?FCB73PX64 
@CS, JED-[#UMF"#%'7JA<SE_ZRW/X#:,P"70#&XB&1$ 
@<))9*I%"EOD4#X1J^8X*J+1./!=FA* -PV&1CG-M/O  
@$7ZIHDQ39.^P^#IU4%5Q"A\UJ*;Q@\F64]T=D'J1A_X 
@2!(G'&!G_D\]^.7DBM?.O#TCLE;V9MQKL!FD2(C"X7P 
@L7+R-NABW,_C,-\&=K>.3EDIT2CW%R&(B@\INRKD&]$ 
@6VL$!]QN,//F8Q=]M"P0/ZI-.08,BFK7\BE>"/%M_K  
@&RPZF4CW^53@CXQX(X>TJ??/*=QZ^+"A,_!.DCL7:04 
@S?=W6E'5CCYO2S] OR!>[2_] F2<.]B+"XB ^AB&4@D 
@<R1*B$E5+ ,'1GD-?)D\?/<D%X,\+L9-:V:*@N_3X)P 
@P7]>-FQ?D(H<;SY: AD/+)%+,JX=BOHC]51P?Z53V)H 
@ '!37:?1."",N34?&7:L;Q"[P6+,V_IXDON9]?-W9AT 
@9?I#AN\ =939K7J 11CZP?\2!,Y<2;TX.):D?I$V(=L 
@#K_Y(D_NX8F#I IH#9O7^#C.8^ >\K8^+KN*N#.\WJ< 
@M^W^8ZKL-YH=&I X5,WAW A%1#FP; +[JUSF:J7S6.< 
@]B=S8_JU U.=E5GM_WL]=0>@;G^(750>,LS%[BNLT'8 
@^OX312* 0N=O=+DL:OK"/&YM5#7>SZ]'!D_QH(D\]&$ 
@OM@T]9^PN;>@\IJ)!.FXO']0?:@JV!NOG+#*_,#<7!8 
@5MED;OY:4[S_W%C1:D_\O#B>J&YV'GZ8E8VQZ6;S,U\ 
@J2_"U,<9"I ==\9JTON_N3B6LY2"7\YV$;^LA)RTF!0 
@7H5;J_L]Z$U-AS&H:6?[WY=O32O;HDW)SD5*-&CJI.X 
@K!6*U<LI,XFWI34R*11WX*?EL1-?L\%>4 &K@E5*P+  
@*:T.+&!+0<XX1$QOFM/T *?("IA/B4XBWT5\0DQ,(NL 
@;[FWLE/,1?MS1 .$<YG=>(;W27ONBWXMGNFE';Q@NP  
@ \*/VC#93,NRD>5N8DHG*K@ 2S-A DE>6WS\:5(Y^U\ 
@H"J.=82V:JJN><@Y.[B&V<D2"8<Y<E SV,69L"XY QL 
@M_%1J*HCM5.F7;]7U6FD%AJDCAD*F E\T N/QW5@^)( 
@!VKR+$8%*)H>;/2LD#__TH]C59AI)O!6A1\_44C$Y:, 
@*#J;82?^(XIRIJ=*2]5?6G&R+N:AT&6I1/MGJ(P3)*L 
@BE@CU-1O+.9A.V?$Q5*AK+ 62TU5\EHKC) !6Q#C93H 
@7N>65\<EO\;<D0L4^9Z]JK27A2N/BG#R@><*CPBA)7@ 
@T#Y?=E(Z&@>+C8*T(43EXCRE06HSG)@-:Q>+=A&ZWN( 
@0Y%4/(Q9;LH*.*Y\J*J?)CHR\COWQ;P+_2"=HBX\3;X 
@ 5V8/\,Q!Q5(A\.X%<:N6I?!K2YB8"@IN;;^":&!;F, 
@:\3^6SYKG$BWC]HLCE KI_FO!\%]O8=)6ZIUP_K#WJ  
@8]AJB9MYI[]"G[VZK@%M(>-C?>_W<,:P93EP2.Z4:,L 
@S/?1X>571>VPYM\*W\,RG3E^ZH8V@6O[0L+B>A?C0I< 
@?1=N9MS5>&2V<B1HRJL\*Y\)U=MC*)0YR/$XM_>?7[P 
@'=S\)1&.R:76?VNI]%!Q>?+=Z0WVH2CPCCFM9CC?;B< 
@=Q89A35446)\BY?W);FM0N>':!',P')MU)VK8_%;-P4 
@6B-G8CLJD<68!S&P]QA>?"G)UD-7IE#6"L\_YD;<8T  
@W1J[XDR;: Y0\LV<(/;9P;@O7H=/! HM#0D05LK;()L 
@G@_+2I/,V'RENO!HQ@2:XK?C+'$!RP-"^"P*8\EM;2D 
@<M\'!#2JY?3;LM^!@ZBJ>*>SGKF^C!HS7N'7#+M'&K, 
@*Y%G>3\)R$;(CT3J\U4R.(KAW4JH9ZI:*&?6^V$?0)0 
@$H!+CV!.+XK[^K2SD;DTJ!JB%WH7G3BTLD%.HZ!T#$D 
@"\R!N)T]$M'RM)^O!&>EGT9QV'731_$9D\WGF_PB&;< 
@JTV&S4F9J6HXCQ0D#4,+J0<G@@(INN6%]U.VGCGE*2X 
@@32INJLS6>*R7JF*Y.O# $.1CLU+8T\F$4TU%\P@=DX 
@D&,]\5;5#Q=EJ7)V4MMXCH;?JO;_W%@BMHDSFR]"6G, 
@NTV7,=%0VP/(UN%A[-H!XU5%V#Y.7HX$:$Q\Z\UB5P8 
@$0<W-!B21\PJ9]BO^$!,4)G<7QYM'_>;.$1CU/7GLZ8 
@GKW49F5,/WZ*M0V%U::J%Y6VL^C74;MTHC-,R6(TQ:< 
@#I_'^\[<SI(S?)9 OOGO9CUQZS/7Z;(=:/G9D[J90 $ 
@7?9_9M33'K81.-H,/:+L79M3^G#8\[K)%EFS$!=CUQ8 
@("PJ<MH5"%81MN11W^#&+\"..Q.M)F(>%;N"4>SFGGT 
@DB;<.6W+=8<=8Y23^&AQI"$[@/*5XM6F1>';Y80@_2H 
@761(Q/'AD@DH3J/VT9J'K YFBX*32G9!F#!38*HC)]L 
@F"WD)9[%0'>7$1:G&K<O"5/@VAH$+R4*Q<[5=K6/"'L 
@ %GB?1>05GY$%'@D-'CUM)KGEK;_>,\:;0D,(OQW,@\ 
@"%)QE#E9/6.0KBB8HNFQLQ8%I&[@LSNTZX?-X)N_X:0 
@-CT&#(ATU$;[ 3#H?Y4@#2V27#(G22$V(U9U=OF$U*P 
@ER'"W]Z\$RN9<*@ADO@\VF!_DJ<H6O!N)V[_*N6'V6, 
@"LH3%9;VO5G"6"OBO)8YT,*1,KD,U!0_!SRQ;J*O -@ 
@< %H X$#XK?>W-S8C9PDUGHCO2Y#R+^3<(PQW09BL>, 
@81Q898A)50_ V "?-,B+__/DQ?=0.W%%=Q'?+M"\@S4 
@YI)0,57$XS3<.C\/FO&)R5A Z:A!UY,=XZD!@)>DU0  
@<LNZ0)RK,]4O;7N>A=MUO86UAW@)N403?J34VNBBY3T 
@[LA29BO_.M4.^![(DW']2(GH)K5B*CC;)\S>U2.:>K( 
@?@2G=&_XQ*<'@](KN+B\2\HJ,?OL)N#_^XRDSSE.:A$ 
@@!\4T9]^^\'C/;S:!?GN)WEQ+#JVV[TU3@9%CT/AZ5  
@STY238BHTF9%14(D AO(>!=[V;F@:**,]AW(?/%#D5T 
@20P"L5(9H&R\NM-'71>Y'1X+#WW>LY,TP=-CZET7Y2< 
@:!8YU)%V>EEP\P'M>+#M*=\\$D[H,S"0**4/&ZD*3!\ 
@ C ?K*P;*9<>#Q>:P90%EZH9PWJJ0!/DR.(VTDT-E?D 
@,L<6*M5BFT/^UDZ&V6\/ KL#\O]&?A0S1V[?2K\^^WD 
@]49CD%<Z2+K>;L>A@^@F%^5'$KV;3+6&^QST9&6"BV8 
@?+'$6J* "6$L=$,F%JZ1&@F]P]%D$8!>_7;SL(N-2*0 
@G>=2[+6</9:)UT3F\T718M6<37LM%D)=+ASF37R#N<H 
@ZN(-9AIL68?6BL:'_R#0R 757P6;>HWTVJU.IW/MDT  
@=H2P=!GR\#MK#S<>?*1'O:I6RKLI9];'S>_C*D8,]U0 
@8O[QQ288)YW8@5<4;L3*8I#,Y/-P'YK1(F@_VW/AAN( 
@%(^";V$0+0.@ZBS3C;DK\.#EAXJ3)Z*E&[K*Z7BO5I@ 
@\.<H)%*:?,$*%W:XMQKA]?$_1![8<+@T?W'EJ9JM(0$ 
@Q?CZ]Z@\>B-$SOB2\0C:P^14?E2O=[BWTM.PHD ZA:8 
@)$9 K!QLR*Q95EE LCS2M>-1J)7'DU90XI"=;@SCEKD 
@^M'S F$#X:W\9L&I/9A%>;EU,ZNQ;0$KY4C<K,L?AVP 
@4Z-N!CS^06.U=6 @O*[7E&4PIQR=3V\.%N^R2Z6JN@8 
@X@P)NU4SVGBKR'UMR[WH2ZMPIHK;;DW+V.K+3C14U_0 
@=N6#V*&S "GO)HVGG<C/A:5X=^ZRY\.%G'&;NDIYREL 
@19?B\4@;^W1O_D,>6J#R*J+N9/TM$ >WT:",EXV[*$8 
@BE2Y<%EWPRHC%\[5HIZ@3H:PE",C4;!RHVFHVG;=G?T 
@V>N-! O[V06/)M-NZ'2PM6Y2J2CY%:<_6[XJS.2UOZ4 
@2DT?R-]< J2NDZN/Z$#IZ)] 1Q(^N2] .T63M49,Q(< 
@'^Z4A^8['PN"T'V5BBV6ZT3*LJA&^KP/(=O+5#V&4,T 
@GP#+4_XI'XK%#JJP_"08@U\BLQS1ZDR,@D_)IT*0F]T 
@IOP@M3OH2[W:$"]&!K<"0S6'=-8TK)@@?(KC .?S6H4 
@+'6D[()<LEP*&$.5T H&T5'-M3DY7)IDL/8U2[(/:+< 
@HO8;I?(\DI[)MZ+&%L$7S/3,/Q+QDT(V#SR2 N04TIH 
@"I.&$NJ^HU\66<Y*]82MKNZGC"<2MEJ&BNS]$ C^<+4 
@F"R!*<PM'\C%+KBV4"-ULGE^! *@;%9<NFM+9ZH8H0H 
@?^5?V[I:E5R<JD<UX;LSA4>N@*!;HHOPQ!D[YP,OFX0 
@M4/-1V6&4X3].3]H%GYWKX*/X_Q>;A,:M+*O]H4O$M, 
@BK;O/#BW3"EAY_\VDW/S[9I>V"GK_6FCM=Z^F,"JZJ4 
@L=BIVHG5Z3#"VP]H'B5J\M?%LP1_4\7"QHKS[RM#X8$ 
@CW]+28@I'SIFC"Z(Y>--D*N;W.@0!N$Q@F-I<-,!.W0 
@RJBX/C@J6T9-:<@MG1A^A+<YJZ5J)RC9MT=FO>6I5PT 
@2W[N7*4\9/2KCTZ$O]MD9(!^$RH1.593%TV%I%SY!0X 
@<.[*5QCU#OS0\KLZ07:C?$AC:=WQ&T8725%9KFG#RMD 
@+TXTUDI](?-7:(U:;YCQU),FN#FKM ;3RPW.)8#33]L 
@DF,]: =2$I0!MH12"Y4M16V=+*##CFZW3)"@?SA9G=T 
@4M)#^!*=:43LT+J8$"X^*60E[55I7](H<![I75;V]_( 
@Q,.S]W=7N\LH$#CK5I$;O.6QE7&_^H6<#<K:K8,U5@L 
@U@GN#+R-C&1>?&!+NSHGEPKQRCHCA($N^^)]J.@F2AP 
@L3U?@Z**J UA>4!JG[;8!L",+)RBW.T%Q18PPQIW</4 
@)*-4MGT+H$0 ]?@G@N6N#:&(>1 ,H"?+^Z3S]+,OHFP 
@U._B8"U5Y#PU%<N02IOCF"8*3R,ZV9:9S,655^7X$IX 
@M9Y!"];_-#SWR2&:&V>;%"_LY5-7<>=/NQPB18LX(.4 
@1/S\882P#T#?YPL2U1/,E:_B%41X VB['!&N3(<&F1H 
@6<)2]5#4."WKQGBU27IP7'_ =<,%FY#< S^IY;V@E]@ 
@HUYZ0(.[/EHTR%_$7<.\:5FLD];>9M6*]W4<]P'U;P8 
@9Y,BCU-5AM*QN9LS!_8.==:HGI#0)5^)2X1]U9U4[@P 
@M';=<[0JM3?YXNRVA/#%]I1E:+;7L[R*N9*'4\J0).\ 
@AO &9XY'0UZOM340V6Q1%W\94XFZ* )!V G\\K@'9'P 
@AA0^ZK0G9]8SGB,<]V>-+=.KXI^ROH(RDB2&COERF+4 
@<&I735A@&GNOJ-OS;GT+X/&.+!E"3O=44A'FB ?%</T 
@6U(#^IOE=YCGOR;#,81?>@9E4ZSW"S>.ZG?;K4?V8WX 
@K)Y>6.8E-R;?F W2FDF_?(.![7HG0>CX;7*<ZWIM''4 
@1Z/(C69A  < C0_N@_==P+[D!@@9@05;*;-.?"WC^N$ 
@:O$K=6G,XZR1F;+LM)M&=@S\?XP#XR9+ /<.!7X_5^P 
@E+IGF.MD>JCE4;M ><S!EE^39U@S)/=*G"F C(#]B=< 
@FT5SHOX-=$.&/UGN=\,H_-\G2W<Y$793XDE)!5\O1TT 
@:DV?>=U0*7#'T3 XS:7+ D0+5"7K7+=.=Y>GQR99-AL 
@M_&8DD+<2]-A&9V>#OQ1JWZ1$43O3W4B.U%NI9TLES\ 
@,W]KY**%/02S XP#T:)! $.A +D77> WF:&RA2A,$.< 
@+[EE_&4S>')N4L3K/B)K0T4:N%S*<;773-\AUT=\RZ( 
@O$QCL^5^[KZ)+;!8L/;R'4SL<=O57FDI2C81CCX_<T0 
@@AV#_2QB]8+0GR.U@=8DC>?[6('#YPM7%,VB-W$W*KX 
@Q [*Y@R[)!<5?DJ7GO;2NF<[;*E]QEHJN5#7$73PO=4 
@^/F%(2)-U'![$VJRT91%\(93Q(</8;=> GZ<&)QQCRH 
@,IN733-?H<Z)<!UU0I/3BO5VU<R 4P!B-=L8>!J2,)< 
@[0 O2MQ[L5@)-_#O<](G_O9I!M&"\ E%[CW?WUPXN(8 
@!@SN#$;G10R"T2:1ZD;N;AOS^=569;QCV*,= V9\$%\ 
@;"SZ<252\Q[@-0%$<+$K@ <\WQJ=)[3DT(R4^@FH)"H 
@:\EN@_AM-%&-\A4/;(DGPH(XZ-[_:,-5.MWKXKVO9/  
@NB#Z[0*^UY!-3*96;T4)E3&+7DW*XX^G-@,U9<:@WZ8 
@T+L\"FW/H'BP3^^PA(R9X>@?;( 0Y0@2].T2YGH57#P 
@7=$G62%<W1!+$E EH"U[>44GGVK>A5#J!"$LY 3C\WT 
@7:CH[8E#XWJX902)E#3D3+-R,RG1OVO0CMWD(&Y^4!< 
@Z7#,HZ4W-,&*YC]^]WM,3D<+$YR+S2LYE#>%^=#L[QL 
@?E0I,$:S1_:=ESAI+IY@U>'NJ4MY_)"6$AC-PR>"8%< 
@N+!?E*YEZ&UW3JT&JY:?UTF'^;69,@HXB9B+7RGRM/, 
@"H@(]@[.F40S+3:3B(+(VQ9JC=7ZSNJXV?Y4<"0S\,0 
@ZOX4[,E(<HB,L>M0Z+Z;^T)!C*F</4\Z5SM$=V?-RTP 
@5:Y\!6TLU3?Y;D$]%?G6) CO ;]V]TOR9/RQ4^9@I[T 
@ZE(^B/\=<_1,; Q"&#OB]\7.7!!#5UR[&4ETK>V,Q^P 
@ON>9R=-6H&OX__LQ;)J6C+>K'6Y:'I!R(]CC"^A__<< 
@I0"DB6V**\]9Y:V<3HPUW#L%1C,M2N#6?1()63HV-R< 
@"T'2[6SE;A9K P/2AM_(H^97S]@OU;[ZV-/)H91@6,< 
@N\;8!GA!H^<@<>(13W;93(RM(%BMY\<]S",;H:46"6< 
@@FQV2$S3Y,(-Q5X+OM6(MZ8BV54DOA)Y <J>GF8L0V4 
@2EJO;\O(OFKJ*F=, <#&]_B>-WSLA02))D*V+N?12MD 
@#GXZGB>B,:Q$6 >>0XB86CZQ#4?J:>:;DS0^.?AE15H 
@AV"X^D==/=X6O[LZ=0R8G=P"WG?Q+2Q;+HS/''9#A?0 
@1]8*",&E^_JL >$)BTWA-8Y72DO;&EBO>C4\RB^*5NT 
@M,42PD*"#UB^>RCR([QX(K^A6P@!".&L-+0Y9XO,3%8 
@U!"?G=H PRK ?&,&R90,6AL@;WQ&J. 2.=WYF&D"X;@ 
@CVHL[ZZF+ L,*N/?:](! X4<8-$^X^!B$V0\<SRRNMD 
@COV7%ZEXS)F B/<J6B64J<$?;?=X3<Y#,=+G-8RP^E8 
@2XPKLJA&\I<Q\-5N'K"RH,^# -*!(T&*LEJ]["*.CM@ 
@:0? $)&LC?QWN^ABSX.;$*7/,Q).[_@*#]V5%*S*6#< 
@195"!][IRZ4C:%FTW#5_/?<?=J;_5O)JS2B'9SPE!&$ 
@.E5A4@LW'@_?%/+0$0 ^9O);H(CIR.F[GN(,=K+03$< 
@G!;II(9Y17;&>KX[PZH+G6'T>#(#%)$47:F#&T4,B40 
@N"#3M"%X0YN^CH-=#IP$34Z6B%W3ZV:)$"GI0D  /(8 
@NR<<TK(!S9_5$N+1QXN@XQAC>[W"'494EZ 8O%4[4+P 
@5,[$6U_ZC.D#T*=]9A#!<!/NO$E3EGB?[#/:-'AN@48 
@1*539VI/,"KP,W XP"<:L[Z=I0_3E&T7ZI(H2C?.(4, 
@3WVT1@7,3D.>>7UXH%>[%9EP&47SJ+L")WZ/6];LC=T 
@WM%7_VWX5@Q%J0^!%! <$.I8TE>0HGQ"&\T5\K]28_D 
@$%=V!DT$KXT%WN%C=OE<I2*!S_3EM7:GJ2W%U30;A*P 
@>@AI7G?!G^L-I3<G_) S<Q$\2 FW"^?,X1:G>_4V&ZL 
@MSS7(R-N>5CIYC=U?/L-=-^NQNS/D!?8I#&&X [T,(P 
@:P<% ;\LV*L1R_7LV_ND5(70BD"ZAVO>8)([&DKWNJL 
@#FS.4--\#>>\C<0L293*&RR-:?+:[3&9X;+EFF_&N>L 
@IXV.DL4!=3RH=^WH :<>UR)!RK*FO9;/SYBIQ,7%OQX 
@CV/R@#*U@ORB\OL>^29TA96(+DJ^&IAQ[1?O!3V 'V4 
@CI$0.\5##N37,5):5S_X=SB21]FCCA0A)E):AD%SY&, 
@-S0Z?T'NBV&=&F8*QGOR  *10Y'[7MFE2&H,KS<R]70 
@H*5O[BTU%E-C=^;Z\NY,O($N?N<=1<O[*ZVW^Y<3,R$ 
@V/Q]Z\%EG1@BN%&]&H(EP8;#,..)DL'$+5UC8NB@7>D 
@CNF$V$J!*2)JWMO W>3=F=U7W46ZB.H(DN50$>LK8]X 
@Q/R_PGCG?T1IC9=BA06S"HE EXK&%7E]UJ0@&@;:WJ4 
@7-GM0W3=Q'^8=15&I@%8,&U9=^':-H#?,$LL_%#7T-( 
@2%F[ [$VS+4PVX>R8*<JZ_R,?$3;&1'^D\D;X(9M9U4 
@,=,/;'7M<*FW:85^;%A3KF? OJP5T*VZLV1VC1#P-A\ 
@9_+I;2WQ@TFV7:5M;D=FAV:>W4R,F)^'(%[[FLSW-9T 
@BY2),JZ;"X"&(Z!&B_'U&QK6%H(5+>?Z-WA(N?>3L;X 
@"F#C/PO&(E3 )%,)QA9*(!&7*"K9Z$LUD#Y*N?=H_EP 
@1JBC;3"F='^;84&'H""JC"G62"]L9$J([%2UIP#[SN$ 
@*PM%DBP'JCO0U$'\P8S<-8T[Z#;]8.B#ZYN-0QC;6*T 
@%B@>J,&(5OTP19A[4YMD3+"D/E[WQT?"MAZQ8^)5@>0 
@/>0Z.N=HD;,'TD\,P\U7@E=/L"+]+7@.U;N_!YWA59X 
@1_+\CO+_S[&EP<#MS2_I>6O0G[;ZZP$B5SY+=%R4E6T 
@3:7BU\TG_RO1$0G"2"7PD3YF+&KS6_;L4K/%DO1]#[L 
@X.-W8ZPRXUQ8:4;;FD7%;@!38NKCF](L%N$$+Z#V/(  
@A7U/OBGUB?>7&YQ8V6.H1Y@&!?Z9)3.)!<6+X27^OX, 
@L(L'W_]ZU(KJJ:RR^)P0;-"H$:(GW<=XZYBIYB0A"X  
@]*RQ-8"H<F!LNK7LR>LP:/&%7(Y#3V;@6J$W1=Z'<VT 
@&2'_DT5[P/DNB,7Y+ ^U1!!U#GMEK((#Z*D(/%J_>"8 
@RL@*"7NZ_2>F'7F7:+-)'BFIPC#=H_B0PD]2)%5H*#  
@3=6(@LK^BBY3HZHC?1 5SVFE@AR:CG&,"R^Q;+! LRT 
@CSK\?*"*T-:?U'/_@HT_I"$2(\ECQ'1K5>1"4,MC./8 
@EN/-),D_U[R'0%ZD*]A7X)Z52MOI=J<53]T884@7 4\ 
@E^#II\90R=L$[P,?7ELFGXQ?QBPJKC"0*_$&I,5"3@4 
@BXDFB0FU2>!-D2>,CMEU.<&F$):95/#=I^1,::,-**8 
@DO1[KRL4C>H_P#LG_WE'G*%Z7<7.Z_-,T !(9IG^-:0 
@3?;WGP6L4.R<PR4Z:##\IAHW:&#,N%V8=(8,5[,BQ>8 
@4:$3*DMGY]/)Q\FAZ1[L^'5B10E %;DY:NWO24E[F6T 
@THFT-. )<RJGXWYIEREW<!# S0+NI+;@WZ1]08*H@*4 
@ $2W6//!KN="9OX>$=I< 8TF[% 3:U *156C1+>P)2\ 
@YMLA:/,*_%83PE$-JE* 9\F;?M?]M\II/HCM%: 1"0, 
@NC<JFMFBZSD%F0%]?2A42U:-"(;[%)0MP\VX/'B?JP( 
@/)=M,;ELI ;X_GP&]Z0.8=LV?_3SP<C<;,6[!LK.+_@ 
@P@9YMH=JX]ND!$:TM+R=3P*)FD!F-$C5A>-<EQ8?)1@ 
@R6TSSXU1[K  MM.F;D0KF6$S1=4()'>BFKHT_A'KKOP 
@598.-YO<T*EU<G2'K&4-ZR*/+9!W:;N8$[PF7O NP"4 
@9SDZT<41X>X@%R?Z*GJS,AON#=0^.>YR25Z5T6(XT(( 
@-:N%/.F][])T0X>W0&C&)%2ZDH)QMQ4;%EP+^OMHT^< 
@??P[1% ; YP5I7XA6<B[W )H6:6SOE977;9"QGWZN=< 
@1'96X>\J5^E[8-!Q *<W'B3:]X-Y'>,-&AX5KW6'?&L 
@D+"_=)JC(;6I#*J"FR>!^.T3%V$'P1:4</HE*\@87.P 
@F-%YH5YKJ+=<QQ?_.&[V#.2 ^5W:,H P)S+QN\^A!/T 
@848?L9RL0)%&X"?(3"=,?]/A%KUT[&?_%UI7<MEQ4%0 
@V8M1!C?Y!>TN!^FI=SU5Z09^: \_GE2>:E:..M>]ZZX 
@CVG?A_J-A\"CSL-@>\"3PY6BT\=6#RR!V72;3L4)[L\ 
@N30IZA$H%N> .IX_<LHW%_B?-0JB8;-B7<Y1L/!?M8, 
@G34V $&<O9UNAEFXBR:@6)HKXLFX#NOS5Z;&G123!\4 
@*_+UBO[BN0-G]7WQL^:P:DKCRW!?VR'/\\AF:;O0_TP 
@>P 4G.=. ]'8&M*PW(HA=?J+5.+H7P\E3P&[K^W!!2@ 
@WDO"UB>+AGC(B;RJU-XC0S,JJ&RZ[MPRR7M^>CK#(-( 
@8%1C4XGG3)O+%I^OZS_<\J@GX7F^#([S+<K/0GG\TWX 
@8IT=S22-9_9/U)2)7CRY-8<\D?0&T/"V%T:W-_7$B.< 
@RKW#^O2"3%=CHG;;/'\C1GOV=0>H."7)960/P"9 9=@ 
@_@SA>91WY@N*FIIA5N.C#:F:;:'L_N]&5GLIGS60EM< 
@UX"C:?Z:M.:>&T-'+2SL?L\[&A_G]N@WVWAD<-$,,^4 
@;K>Z_1/ )0CP#XF(EV0UPI3V_/./K483+BS/WH[^<A, 
@"O.#5:E''_VCFAK*EJQ-MA>-'2@]I2NFTPD:QN FM^( 
@+1\98X+S=PV6D<60X36UNBNGANA'+#7Y^:G\>:T2O34 
@C^ BT;03P;:WTPFC(<(:M&\6C@?QG5A<DJ>  (<]U78 
@,GWM5GBV=&)ME?ZJ^FH4&V.%H,?2PH^"78K<&-S<F>T 
@KU!+:>MT'I:(# ]R6"T;$UX$ -PM=W,,BC<V")I&;H  
@(+UL7@R6/09H1375F=%9;\)\,-$!GWSPW\2UI4^DGV( 
@"O]@,*I-NGR?)/M9("+%"]76QV;_MD KP$*%O>IOO', 
@+ZMR,84.,6GVD&&M7NT;,313#U@774,3&2QH849W)#  
@H0,%8 S>S57&(L4PN$U+KV!;>X:.+<V>KF5#3M$U@:H 
@U<T$NOXAQ\2%;VKN0;KOVGH>)H]JY61;1$R,F4,#+EP 
@4^^^L+3\6.I>SD._-A,UR*M#6K0^(Y+0S\?G978..D0 
@'F&J,!FDZVM[2\()50-+)M3-KNBD,S^;A_ [IA*K*(D 
@^N'3OXPKCM/%?BJN**G2*R3^J/0V_O]LZU157CD-&P, 
@I4F=E0"0\; '2\%][@U_-J)PE! .E,DTK,*N)FX0&', 
@XOA/?&%-.:R#L^XMEG&=OL)3Q@_2;#L#WO%6=9*EWMH 
@O>HXPLCC)G8P#,V&"@>RF. GBA+02"O(7,=":R&\H#D 
@;3P]5I*=;A;_[TN63@?2(D(?I>HO+4B,')I5C[CG$3D 
@"6[#0>Q-R\$5=."[0__CZA,<+RB5.KC];.20O%\,(BP 
@BFE0WAL(RZH\.ADUHB;A!K#^+..&5@FFP+ZZQJ3V[(( 
@(".$OR;Y5A(?H6"H=SLX_QR]Y\+"01SP\H42,>UQS'( 
@HM%U4#1^H5W[M16I@VVN]<;MUBTVDL_%,\BB3BR[E"T 
@^T2J RQ5WMU^17\\)@.MEB\7+H?Z-,>W:_TY=03H $\ 
@6-H<JC!%M=RQ;C[=RP5LPN62LI.-_+A1AP#R0*CTMDL 
@H7#/(!4/%"YC4^^*MXJNJ#):IMNM+H60#UX&H=]3M;, 
@*RZ]/6UYFN"9!?>E:? O8?J5^*J0#MPYM73^5E9=,>T 
@IBD>2@6=C)T0?SV;CW*"I;2;!I>>0B[M+TMIT_$4UZP 
@,8K2/Q_FK(L ]<@_IG@ORK%#::XA&[?W.G>&$C%DAB8 
@$&WOIZQ4SI>JZPBT-9R1HV,<!#E$F)*;E^T1/S1(NBX 
@ .^;PAEVB'F6Y:XTA(""YN;L;7W?8S-4T,MZF,F>F$$ 
@KSN>^%Q+A999/SF'G$--NY,U^9/,E_G_!M0T_-+.$N( 
@=P)VA6K\'Q1=-F7[E"PP4;)F(G,/(.+5W6)#UTQJLGD 
@88XCQ7*J"=(%?&)B2(_O77&5B3'!C'+C&SR)+4$K&JD 
@WS8U:QD/14G>N;-U,&5(#W"&;0V%%GM9S\W0P_4PO_4 
@B!*:#GKY>VXU0M5(0CHSX--@=!FL/A*/9B?YF;?XG,$ 
@L2]'N9C1X?>K$V[N1!@4J36;:?:5DDH\QWA/K&ZB][T 
@N_<8>I)PNV@43N'ARM"[H=@(ZN0>THS$0.94:N>*QX, 
@C'T=:IZH.J?\AQ:V$3[PKZ1 0D&H#>AY5<D0(<!_D?L 
@_ &:<P!(T,N#T<0TJ2A+GT=J:_';3S!"=MLQ(:Z9W;( 
@RFJE*NB2Z:= )<.E6I1]SPY*$T9S.N*[CI(9GP =L1T 
@CD!"B$]1-8S%J]1+S+*T3JY_:K%Z*[KMM:OI,C#MCZ@ 
@\N#45<<H#)Y?=5YZ%>1"Q._G7G@C\33WLQ_L7<&'^+P 
@E(PC_=-# ;. Q(E$#E;O]L[T</'464T&ST$$7%^^E"( 
@V7H^(4,XDAV!PV_ !FLGMY#.](TQS@S.9R.)*I^L7[@ 
@A$;-1</G4IA[0JFS/LVG71_8%/\Z&\4;>"&]FY5E5>L 
@/4.O&50T-=9^;N8DW'<#W7)0),-5+M)S[92RA*%[VAT 
@N! "]P^G<>,1;LC+;@]F9;H=#]T7[&[+S(ABWN(0^SP 
@I=O8BA7OT/M?!=J]C="&/=L@5T#2O40K+*5!$#K"WSH 
@1S4:7K0_M)&0-\[$K$W+SFGD ;9EVBWS=4C4=EJ0K"( 
@]M.A6JJ#@50Y"FS?O= 6H]AP7R+)6"IDC(RFY:@'XX@ 
@KS.FB7=]0S[V-(&<X7O^RF_RF:MRRB*RKB)]]8$O%N0 
@>5@)+LD?XHK!%3KMF2 IX/#P<6;R"OD&0"^-+=3GVBD 
@H>?MK&K#V>,B4P(564\K!^LJ^N H2Y'-!TZ/Q:Z>F]8 
@:-0B.@!P7"0<D$=PV#8$\W0DJU$DZ5%M69VIX?XC.IP 
@=9976JS4B^'(G!#;,E%993G!5[VZP$XW;U_\10Z/.Y8 
@]H=OF*J-9,;U:0M7%6J=P[CZKR%3XY$G+913"6=EDP< 
@PO+EU JY#5*OMN1E';IY?-::.%!1L5X/K1468/WLR&\ 
@T%Z0,C4=:_,RDQ:391>"1XXG7(QP%/&E\_^=WM$"(DP 
@)I&QW-$OH4H2LN5V"4"!+_)2K1CZOJ,L[*EQ'Z3%GI0 
@K8+F$M"A&(]8Y3;[.]%G91H;Z%;0 G(/KS"R7;HI,^P 
@>=LN4<":<L<Q?!@BN!P;51#I7++H8M1X?G,C'P)2.WH 
@"A_D>PVSITRN*'!<9RILC74H6%0*=B,8&E;,MF6BLNL 
@M!@+L%=<XYV$C35A&G4/\;[S^'9[I,\4F4C$*$U15O< 
@Y.<DI&:'6[;#TK]LOI:_N\J73\#.;%OK>&+2K)NNB L 
@H#*C\9$HK#+/=WC2)A4/-'BJU^^[UKI3D))S&YUBE,P 
@8>/IV8.8)(V+*1.G<CA8NHP T4F"<+\'_81?]$N^TI  
@ JR3_U1Q*'3=>]A71N1JMV]"W]?,4]L*P"^6-,J1+40 
@H2L%IK+5UCDOO1VZ,L""MWLM=H:^H,Z"?Y_*?<+WG_T 
@AX\$S*%GP 5ETZ;._)@Z-5Q";6 3J*V@(H6:\VN5J[, 
@!<2K8+R\MZ*;)%931_X^I9_[#M'9P'(RQ()")I=2\(\ 
@/;=$I-64DXJ86[.%,(CW3P,I=/K1%XL1#[@4QQ-0R-\ 
@.K^SAPE2%61#$T'1K6Q 3[)8.=+N^(O'6?*V/.3<)C, 
@:S*GZ;\3>74.9F!#$Q@+*IBO^6[?<0_&\K]F<M,QLQP 
@ G/A8*+>3"GUTSOBQ2>MVTJ;R0]UR*/"[F#DPV5%&O\ 
@PV'.&T3^CQ YR]MMH36*M*6T7CZ^FR/;:'J^#X'S2X( 
@G$)(8QM,6 #] 'NZ%SL]A6KKDM &*@B+7'8F81] KP  
@FTKV@$B08PGQV<QZ7\[';<E[W:4$@=;YYC7=Q=A9+=@ 
@@8&](BUNPLM9KNG_<"'#G%1+Z8I=9KI%UL$V:5>U](L 
@?ACA4?_! $TX:?PG^)13B"VD+8^3QEAE@5/1TZ"_4;4 
@P1/R;CWZ'Y/0O_VZLQF1+!G(>>_5@K%U08/62@@L)SD 
@PL,>+RG&\Y22M)!DL%PDP*/H\K\_M^(G@$30@C7"&40 
@!3 #=UCJXMBY[!T8,"%%M'U7YY$V4W.JG&E^@#+E[.8 
@I2&D=?D7(3VNMC(7:AT Q3;X]\ZX@V0R?+G7*UGX#-P 
@H*N6:9YY&A]H3:N"_#N)2""V-WAT=7^!I&!&P1CY*00 
@X-9"EP19N_TCUZF.7+I1GH>K*MH]2,49]<9G^)XDA[X 
@IX]<"!3V"Q0PXA-'_,A3M>!+PPLYV1>/ Q=K#]?I<P$ 
@-ETW(H/*[.EA189KDDG.>( OS4KVB-% V4^YL60$4"L 
@]Q.X7'J,._)$!G6;#E/TG1R?8]_=-X84)"P!\7>^Z24 
@9Z;AVT?U;XAZ)V$\*IN+[-^M&7(W7\&$V- [ANPMJ!$ 
@?/#_6%O3$VWMGE/LJOGSF 8"5%O;*[4*DADQ#Q53\.$ 
@YV45Q]'ITZFY\@."B<[ W%#K-:,)H\*V:$2]\CP4'/, 
@9*<$4<J4][&T3K2HH#GQ>(P'F$I _BJEG4(OKM[8$/8 
@,^@]Z0,$\DI><.Y5\ &(CI25A!(,H'R!;9]MDX3GVT4 
@_K';M-C\;WG9:%CYT0&4'4LC9F>4;ZL@04-**#,;%*X 
@A]"JQ.ISO5\IS( (+#<TTL^9#:J=9;$#6PD3H]+;+?X 
@CXN4_<IP)5#P[&[+ E7L?@O@<T4>*;2M4B6E*19V&5( 
@HG0+@68.9@"AY<&51K&WU<JN%63QWKVX@[[Z3A@, I$ 
@G7U (VZKG2LY7K_$ AP'U9*K7G?.4.RHV=%,6@6AW D 
@'%J>']H5Z.$1)*:FO579:CF*E"0,ABAM.AB8<#<+*F< 
@5H>B4^K=W#N8^74WGZ54/[ 0]()Z@H"G)[#>N)[O)UD 
@1=A;=ROKWJ&,_PM7>VS*>!P?BT,#B1'HI4XH>""[AZT 
@O;N<A['!J97@Q[A_H L7VBS+ PY[:A<W//@"4QH(C)D 
@@GI0A(^>NE(E9#N%MQ; * I2@(*6HL/6#XIWK^W-$/@ 
@09R8E('ZN8;JDS@'"HW205.%0.!A[: L&0#8K?!R<=$ 
@Y?BIBDX4%PP3.&"-,(T'[QKT65JE"]7\ I$B:TYT%>4 
@T*HS*#3'?:>OWPGWB.YR=,64KMI'HQV'//@F'^:U=(H 
@&:;JU!WG;,5TDMBNUPQAFLAD.+?MR<PW;*8']0AR"@  
@L[Z*OQR*3%,YM#]26@-OX@6G*!D)J\.5%8EIK#$5WF( 
@1,:ZWN##L-8S4["&8&K(MK_(+&K^/S[+*[$O3I@F-XL 
@V,8UNWLJSM-&Q2=5HD*K&OI5_,U#.$L!_J<UK&&>FG8 
@A:K='Q^7MK%VZS%5*^-Y=1KK5 +UFX>Y&R]Z^KSGU,X 
@3>B=FR1U =7)Y1$'JLO?UO)>P&&$.P13M/R*<C5UHOH 
@QHC_8PJ'ALWW K)0A<.8H(4A^\V&6%*VVYCT9PE&_VH 
@SSF>RW3"IIA.WG<E1YH\$F!2:*&2^_V@M@+G%!(WGZ< 
@P7HC1_QA#)_SY5:D!F^']G6KF)+@@%A1JK-=";W>]+P 
@.T$=.]_1+8@32=\6(W#0EB8?N'SU8^1!)^>J!?2AAN\ 
@(-W&OT)/SJ?%Z"!YDS57#3N[$ASRB [8I17ZSDE%X/< 
@ /)\L!CNTQ -[B/A3ZJ<PB!H>%FE#SAP3J2">/=&B98 
@Z0YLH3WR;_"2[0CX@>G/EFHG[O7[IRCK_<HK6L#Q/%@ 
@:BZB^D/N-VS)5CF2E0"8\/)J'(N96(.DJ&96N5\&'HT 
@$71%%$DU1>XQQ4W9%9VE.V<O7>G,7$)0U'3O9J\E(T4 
@[X#ZN<X^<6WAQ*':.T(+?501%ASICLIYR?,!Z%:=)AL 
@_366*%HA2M0#W!(G?T89P3OS<X(H*4XS#I[*UK+[^YP 
@*RB08D1ZR;C*9+:=.5=[^^ J?AG!A\XI"DABF=3YH^X 
@';@H0F@08H$D(SB,XS&>"OEER7M=:[_X4A\IYN8A*0$ 
@O^&2:CWN-\0:&3,R^>MK8@,EM<*OZ[8GY8Z('1L$\A\ 
@YL*1]?=TG =E!NPF A2@0$]4EMJ)U>FJ4%>S*G$+4G4 
@\12GQ-#M\_$6!XI$P+"R)WBKP9I/$###CF"IJ>8_G\T 
@%]+#BK\3UDGRC7XYW:FC?F*G>9<!'P!%QLRYLY\%G&, 
@?-3O5WE1B(3Y!H( 4MF/HY"VYO*7TEP_O-(0=F\E3/T 
@B/T/E6?NJ@MJ+'^&K.I5)P;CH(5V]:URW"9@L:'0>0( 
@^V"K8)*M[*G-L\<!+__  $V6RX<-MZ]/LOQ4CH8G^O8 
@8M<['FC=0SJ?$V\:D13R0'GN^8K?=8=9;38DC.QU R0 
@D"G+K>-CYT+U!@&J@'MI$PZ)Y#]$;8@;6WAR$/5Z2W( 
@<ZYBX)*&L5-EW*]E,7+$U@M*9\C@5E_*AA$ZPW+$[U@ 
@[I+.V!"/*%3'6%T6VMUY8Z57J>[)_9571F_NM4MHA]0 
@VDP)?O(:D#^$-_*7L0%[X;G O[G3:;<:N=9T)R1CXMT 
@-<]CNY7[:<0?S:!KDU(HS:1=<3E!/?_$@\>Y[A1,H78 
@+.6,$Z JN-1Q\IEEH.Q]D&WQT(BV?2*:=;*K?[3,2LL 
@T"S'<S"Q\3L0N84,XO%45P8M3+RXR>QF<'V:J#(6MS( 
@3%!TV$Z70!Q $LLGK0*PNZT\FW>79-30P?W?*&+K2^P 
@#E7$,<UK#K&7QI?._0^"@.5L6I L/J43_-=Y/E_RNY@ 
@<2C!9I%Y^!P*#X2=G_!8AP#"01P[Y[#6@;B#U(XNUU( 
@2 "6*&07&IT_PEA8NMGOPQJKF8:&#$6'F<%OCCT.->8 
@]:(+7,BZ%7:]);"$@:W'$M6_>+;73(T\URHI8([G;N$ 
@(TRJMV&2O%7HLZB\YJ$O=S-Q:F#2:/$:'M?CD-/FB\8 
@02G #13?X51(484QK"-:$:UEFO5&_!"XY[<W_YQ'&,P 
@I6PE?.K2L(M2I*_X6]8U'<&J!7FQJ"3#'1R4#]>*_"8 
@K\SWS(F?\;[MP4DA2'E7:NEW,K5JR-0()=YKTM&Z%/  
@DA(A+ATN)E:^GZK3F'K]I5L:",8)U=K=E'*D_FES<), 
@6*8*I0[;*R"E5!"IY!"PB-BA/\[*1 3.1VG!Y8$Q"+4 
@;OCJ>VZ?V4F;-K/,>4']RJT%#T7"(K;A?_88S&0JKX0 
@P)$1A54W)(F]A_-+4$:6(2NIA[BP2L78N[2=&N%$*^L 
@\\S<V:0??*1GMGC\%^[E)>Y\<QB'?L8XJ'GYV@!1F+@ 
@L/K1YM$_?,36 T8KF+ X)!-9 TY=S]@\[^T^DNWVO9\ 
@.J3#MJ@=!P8)VA*ZC+TV^6G@!"W\!/(84U>&3<NF 6< 
@;:5<QH^P-.D'Y-6"<,]KOY4X[KM3"P3FH?57JMS7SJ0 
@Q.#M\$LN.K)9JAN_UH3M^C2'!&S/5JC.S4NJVGR<6@< 
@B<SO0JIT?+GW]F><T6ES WM=6ML2"53* U[,]!(!):, 
@"KCHPR1T1BP\-H[7NWOV,L@HV[%B79N%#[=$@(*5A(0 
@A+!^VKD6)RDXHLK/86=%7([?(2*=HJI0V\8]5;]3#B8 
@GE-+1'7&,_##N9$Q:Q=4?47M^!D(2=U&;0.BQ2E.]-D 
@/Z0EA?)SQ%4N-6 @D;;EMBKBGS[].QV!IVL#%@PNM?L 
@W!3,!I=\WNX+M()^B%=2%UMR@+ D+/2ER$EN9:+[(6  
@64I,KY%>0V%(T_V9LLC72/WN96RJ"?5HK#Z)XIG'<4P 
@("4E4>/Q]E,-ECRTG"C7& 4X?AU^G4]M!L*GU^3\. 8 
@].Y](EL#1KLU/(A5E6"@#@O@01ZHBWAS*YA,3GSVX&P 
@A![9C!.^B'.!YP;M]1:^#%FY.3A\GLWZ"D^%>93NJDP 
@L&G-XZJ!2#/7EGVVM$F'D7[3GDZMS%)^)=EO&IA,T/\ 
@93X9X["N.WFD1X O_ XSB6S32N73Q\$VB75  9D>.=( 
@*.&15M+5L H_T(O"P<&8TF*@H5*4FH+XD0K"WL,3^,H 
@1"/$-$.M:XQU8TF_K("TRT!8W)J!V>K7]P+I[E,\@CH 
@1$-XS@ZJ_]0O#&AD'C3[L[>]C5B=IN0Y8NYC0@H6@DX 
@-I@%\ >,149==3WLOR3,"^"A"P7H ,7/;B2A^I<N _T 
@I'M@*\..#LLJZ,S-5/,"J[.<BC"0;RZ$1@F;?VY*Y)( 
@KG?=$2K 7<1=1"PB3&H';@Y4X<# N7$<D03(ND> L/T 
@I%#N@8DXETZ+QROPUV5-TX&8PH:Q@< >6MG\T:E,WMX 
@:VC[\!XB*1.#U'@6C7ZPV<W>>J,T8- &7LY+&-Q.!Q@ 
@\P$%T$AEE.X.:;Q73 Y=_KQ%*FJO!,PP%W$SUK#&,U\ 
@,ZW9W;00Y\LA=U9]VXBIX&&V@5#<(K#4YWG3Q)*/=B@ 
@PWPI+*V#!I^P+,-;2<^5#/8LVMV[@>(Y06:"]AC=8UL 
@A/$TNJ?IYD'V\Z*1I,<^DX6: M$[D,&E'<I46FHY[]( 
@^G]Z^% B)W91".)9!PNKTL=OJDO@IC.,@0Z? 4U3G0, 
@: GW#H0PUTU"3BLP!37J#\J-AU<>_IQ=P %NQ$/@CQ  
@R,W:OGQU6;QJNY$SOC.[^M1])*LYY%0NQVHQM?^UP)( 
@DN_$"E$Z?,-!3OVDH)PH6)I?-(9\8EM%#*1>?@*$(E4 
@]%P!RI3(/4?,Q93R0_[3D!-CG(59/F;^+9>B(=V$Q>H 
@*:7T8PR#)__^[$C<9"^L@'2,W)SN?11:J& V#XN(FS, 
@\2EOM R<!E(9;9O;4E'%/4(TWAS11PF1B-@G@P=V6?D 
@&@P.=S:Y'ZO!L$<NQW$U.V#>PLX^'W/^+G^ATG)SK^4 
@R@J4M(: &',57D-64]W/ ;N>DX8[G?K Z9 :ZM><Y(4 
@%S? ZP&KPFZS<@%35QA8B)%KN;"/N.XB&",LA>!!OHH 
@&JBWR*5X-**C!)V'-/J52TGS!R*QQ;%"Y8*XLS^1U+8 
@9U2#==C,5'( LZB]+[#!VZ4'6QT2<L5&4IML*L:K8S$ 
@=: WJO0]\=U261S.-S<9@+ GAC(+.&=8OI_(NE(3Q0\ 
@NV\+R]M85 2!!<[*MBQ-6_OI&@XG3G<?!P_X7/O7 0$ 
@D2)*#]$1%AWGC\"C2LL"X;:U/P%#)LA#!R;-[S?")W  
@:R&0K+]"E\E.;9L4"T'E\ BW-?HS/&.:(/LS=-Q30M, 
@<4PE!&[B:F^@BG\018E+*\9N>JQY.4MH$&>1Z=@<WO4 
@PP-FT+9ND6/^[]=M_V2J,#*VD)4>29ZN(U% =C:E RT 
@0V%6&\.;HL^]&<01C@ -=2W ,BK&JF<UCJ(CY@]%9+P 
@V*6]#KB[GI81X'!*W5UA\>J\:!E3URI)>[+']?B 4\D 
@F'I9Z=\7O+#N"Q&Q@C#15W=S<M\#%4 )%D;F%6+;7-D 
@,H/L74L;FGCU[8AQY7!$WZ'G"#7@?V=FR;%_YD1^;=X 
@0T9NPA"("6^6$?9=]AM6".M-WA=6AV3>QENR&FL8_X\ 
@K.VI<(A^)W%(._[NHHQ)Q7T7HY24WC@)VHJ%TP5MALH 
@>V [=1@++"6/[.PS+E&2V3MYI*4.1<^.:\(.M$M/P6H 
@PFOI7I_$=&=:]1Y:SJW3B8^0/Z*@<=1.VUJ<1U6&)2@ 
@4)[(5X!ZUSN. <&4WJ_]:K"*:<KXGBI6("]>JO*ZFJD 
@M._VD;&LNR)%GZS6\16C9GB9+4&Q%QZ?W:T%=S36L:P 
@3W%M7Z7[NTP%Y[B+S6PZ4JR66Z;WAZVKIC.$0@PU5-$ 
@\?C[75Y4\([MZ H*ZR+2<[#/P=E)/2OMXQ2@NI$/QR< 
@>X:UC@5W:^ R(9 7)HM"SS8+SBFS'LBG%CCDW 4DV-0 
@OZ+25(B\).2Y-0 WV!5RR??YJ,)MZ4G_)3F373)Y"CL 
@LRET.+L] ?8;'[9C[?$8MR;G+]YS_X:VA+\H;6RTHX0 
@!1"SO; F9' /2X PT3[,15GY,K!].UC8.(Z6D?JR#[4 
@!A!3SJDZBC$&&%D'5J3+]#>!%S7<FJWQ\11C_K7;"T4 
@@NI]>)>XR19DEP(0(_)=1*4$S46.#0@'+J;RP0M]1G$ 
@LG*Y_0$6$%(" )&3T5C4Q+PU1:WWW >I?G7#YR.LA2< 
@NCKZ5S*W6BIKZ?MIQ(R5]'%EKLX$NU8[P#H@'BZ219X 
@H.;0WJF1ER-HIPR%P4NRI2^^C8ZF7OY?@;+@I![F''X 
@/ *88:G4B:IM"]Z#7MC/=&\+H:#88_^4GNG:]5.4ULT 
@\;I[I]OF$+VS8@H(Z]%1#?0LA;"S)(P_ PD?C10\9$8 
@)*@(%+V,OPT[^J/6KI.Q<.K%#Q=FANG#U),E<UL5E*, 
@G7C(K3;/>FDG-S'/5X*;TF>N$-D[8DR6@W"R;Z)?6,@ 
@QU^A[<%8N7K%1*Y>.+81M,QRM%^7;4S@=/]2_W/Z_0< 
@AC'>AZ.-ICD1AA&.WOBK_M&>E</%,Y1C.A$!!6M8D:( 
@8"X0N]-Q<[\+'S]Z)?\@G3"^!>,%/=\W^:;ZLF7Z-,, 
@ 01)\'JW00P>$,JT8*)4'IH.+_SPVY]S>"_7E&=@I&\ 
@=]S1)Z4%_V8L::8XZT8;0+ 9P/<.QR.]F,IT.), OU, 
@#*RK,K_W++:,;)OFC<<<4B6#R[MB)]!$O'!Q:.Q,6+X 
@D0!V[F'N5;W@GBANAN> _IX=9B;55,O@:F'.O*14)=  
@O,2TWU\&3WR9+O>J@_LH=?#? A9"\//3%^CK@4]><2( 
@Z@0'&R/,MR;EL)/K?5U:;!'FZPUWQ:#IO*XB=V3(GB0 
@3C)_E!6BU&$E,;4'@5%#(1HI V1U9PY38[]?:4H1/]8 
@Y%HL5C?&(VU-QPL*.!M_6S$B-H1+;(VW?RUX6Y?-P$\ 
@5#KN%0 B/0^Q7>6E]^Z4BT2=?0H$^LRJL"NMRZ\C,CL 
@TT!, K13&M*<)=/A TQMND'UI&5Y!+#QT!>W4Q1GUX  
@&@RYU=:N+O4Y*?R<<EK@WH[K6O]]&:-O)1WUIKS;M#P 
@B ?/,+>F6#W#7_" +H4,!H!_R]*:$DD;-$*G_16IG@$ 
@820*3S@TD_&N/$RN"__[9VA2F+5],;@'2I%S/\ 2I_X 
@ZZ_JCLX;72 'K5V]V-N>5"2;S WFQ8,#__H22]=9/KL 
@%OU:/=1>D+@KIV(TFH(93!0UW9/%)3Z7>:'<?LJ,M>4 
@ZJ7P/ST[14;KY$N2#E:K.]3PYU$ MVVXJ*9(EU_MN(0 
@!:C/4#"25CQC AIV6Z(A R!9DX5P#8_;*32SU5?4!,8 
@&<55G!H1-75SU)*$H) C Y1A6TK+.611Z+E"!Q3OA.  
@4;MOH$!\.WBT=34)ZOQO=YL?'<E1P1<@Y_5$I0=(].  
@*X=40#O"D;&E?D Q#]5N.C(Z:,L^%]@XOV$T@DGP"E( 
@\M@EN!'>XDO45@/$(:Q4E5ZF,U(VRC!VVAW (VSM-$< 
@#*=%TL60N;@!+,,J?B5D2!*..W/G5,DR;OD>3 CJGB@ 
@?)>F'I8,:MZ:!KC+_G%F14GFS!J2D;$M"9@T@7=E\M< 
@$UGW;0X/=X0+8@BFWTF?H/%GGNG/MPBN"=(,,<@029D 
@-OR6H0[)CPH@_O8C'B_!DX7NT//0^'/-\35&Z'':YL4 
@2[3;9E.N;?:DD:,CW_1[  XHZ]3NR683>BU6A3<!QTP 
@SFU!*ONX+C&GZ9F\"*/F6P]_Z-,F*9:]H3H'ZL*1QLH 
@(.1BU%^$4W]]>HT@8?++2%G[+QHMN-9FM8,T)7-%F#4 
@O>%&4#L"VH6UPWKFTW^PX'6Q1AW%AC'@.I$\).)=Y%P 
@\_]V/3!V$^=3.3&Q#\H%NG0TNBXX)T7W17^0HCF,\@, 
@/ZFF2QR&%)06#VY)+0YQ].W>OCQ)+8 H/EK+<<4:W)< 
@3%W:HU<IL3=TRRJ"'-]Y5K/H!^_55J<$<B,6WB3QQ7( 
@"5?J$[!'_BW'0L=5UPN;CL>(.O)='MIIOL+-<V??J]P 
@&$ [5>+D";)7>AWFF/"=#G:VS.24?I%$T3^'Z-D-[6D 
@(:H:1FXP1>[6>UN,4Q_4;G78>H]#@=#QTD(4.F$F&94 
@4&_X4]\7_8TM$DX,.+>RI-0]&#.A,9BI(S=5EUM#MT, 
@7<JN1"H1M\XO'2;7'=C]X3=,3^C@GSZ<RM*CU0]Q6HT 
@C4?[XE(.L;N;_1S("[_AA),Z[Y]%&=B/+VT_-:/R2XT 
@#"&$?SKVBF$A*&^\U9!Q%TH+#> R%K3B^UIEFSO7].H 
@?7'%A=Q)"R$K66Y9D34J*>2A]/J"5>,%V9M?@9RL4]@ 
@M'#D)P>386)N%-4SZ3ULH7Q5IB *M'9M+AB0!J5..'0 
@H-/5 "\]'$&O16I<S#0(W-YJA!^)W7""*$/18F:Y@TD 
@R?S,_0[9"X%9;IWB)PTTJQO"G0H\XYV37Z@A;\#\4+  
@N;E\,[%1,W!8WC7CV'",9^PF<.DT26%FR?05KT5@0&D 
@_^=D1 9?U*?Y%:;=RMJHE(_?@2P.DZ/"0-,U-Q[T,J\ 
@^<^GH@*1HG-V/<H!PGB5\QGE=DK;CEXH/..7P/B@H D 
@&D4+%I=BL20NO#UT)2A,3%4AQ_ VB3_XK<:@'JD?03$ 
@>9FI@90-Q&OJ_U,DE6:T'94@PB;DXS!>7WS^@4$@F.8 
@"P.9^W;ZW7UWJYBY_533N,'*I'!3)+TI!)?B88 (.8, 
@S3!IV4$/P@[TS(%=8O1(Q_@^BDK?REF7%:!)=+E,@8X 
@214NS%-? &,"T,#4+?.RK!69$+RLZ:,[&2V/8< >%7, 
@P*$VIM/+$O=WR\=LQ)R8@ 'DK&:'6G_==75F!F^*ZTL 
@7Q->!2*LD2DV0JWEOTHUM0BZ8=S/6 ?1^5>!H44)4\P 
@' LFE9",=5!]O9V,1#???GS0Q4I9[U?!$T' HKC*/N$ 
@=Y8L<"A?%$3$XCI1W+E$8:0CJ0*R-ZK3M#M-!&#F1"\ 
@_!&\[7:CI2>[C@--IYM!G92TTH9'-STE1;WM'PK#IB, 
@/L_+2;9XP6ZP:VK1;& EX+J6< B *XM^!F/<0Q=I3[T 
@,]5@*=1@7GJL\[(KB/\M2FTL1&+-A_*:OD%X<'5Z63X 
@GV3A\61%<B>FEQ&,/U"--4^[*B02RH4G%6YD0C& **T 
@ F*0H]7B=>I?^S^PQ&XI*7YJ1<ZQB:U,&5IP6LWI>*0 
@V*]FSH!>Q&WGNJ6 9$8Y9H?AWS6/(L"Q12/TM@57N4, 
@NB4PJ+,WX0@QK?$=F"51J^&?ER%E6+ADUKZ%LDO[SUD 
@FL-=52 ?Q-\=Q=]?<9EFA746]$*(D9!X6FRYP<0\KX$ 
@+?6VQ;P!& <O]?J__!'93<2+O:Y[:!FQHUMNC2B$074 
@'"^%+.>X$U&57"C,  X\6ENXKM05R*"R_KMG.7GS#]H 
@IU.<F.SD17>&N>\MLO:(^OOS"PC*E:;%+5#C2'6R)8< 
@_BXT"<Z;;B"ZBIA#!$D8OG73"K'! D=+ 62X9[[TSZP 
@Q!91HT0-0Z!>$U#M@G>*8[7G,V&8D4DSDNKGV./9EG( 
@4_:,C8$5S5)YEMP%O(X?2_;,+[%;KUNW?>2$J+$!KND 
@-&2U=QBWSU^6F!)QUBU6A99DTMH 7*YRK#[0N7)D*0\ 
@_[<@<.0H:<\)^#$1WI#,V*O'$$+"\XP^O2XL#&CA#YP 
@$C31>'4LQ?1+<Y4^P ,D&,_-.S!G)V5V*Y J8[\1SR( 
@2%!GK,:3$7H[.]:AF?+>OZ<0!<9\N;OT"^WN62/#Q3  
@NX_;NC;J(16-V1Y7^73OAQ!OR2.VIHUYA0;<:KZ5SU( 
@J.[&-2'%$O5,7U"H3-OY3]IP!6N%#NPRL01R]U92&#D 
@_T<P'A,3UO%F*_T1_+WT]MY:BYI427_05A9%8[:6:]8 
@&2Z>(K=E<(4V!SA@@TJWQ?"+3,D:Y=W5)X&_\I(H69L 
@S$SZI>VZBDY>;&Z_22J0D-^R5A-> MLF:C71K\;:I.T 
@0E<C%LCOYDQ<1-0P*$P5+&%%8:IJ]%C5],+/6O!L>1< 
@I[<$XS5_(DF$<7=Q": JE3I,D@U&5X5WB=E7!571#T< 
@*<+^>[XS]J&I2Q>E$#=]@TE2]:D8^^Y'2_;#WO,BN9X 
@Z/.:.(/XZ7<<BF"$I>U0]JL2OX8STL]0RPVC/C_,4M\ 
@E$V\Z%J2'S53/W\@T+VSFQL#W?@/I<X?&#H8(\J#8%H 
@0]&T 6FMTUP#Z\1)<)M"T261'(V[>;T@Y??:UM:2^94 
@FD,NEMA*C&S;U)SGQ?"_W:!TFR7$_!R\)<=1QR\K%^T 
@)LLSQ4I=HP?&$/B1S/X?_76W<TF-89AJZI<:MVFW<=\ 
@%_&A.TKE$[(],<XG;J6":WPO"CNXA=0_V8DLUY/=YL< 
@7!U 9$JPK$^ V$;X?0M#D\9 $G<<U\NZVZGM8XR&""X 
@P2BW3T%<C05"E8-#*/O[KO'6"+:0DN16DPC]&1JES'4 
@:!J1#C:Q]\ZB*HED<3!EHC]]^&/X"'Q!4F?5T@F6B4( 
@H@))#* \.%@6@.)%7O+*_,VM PE@D  D#Q3S''E=%^T 
@-?%)7, WRV+[=6S_!=S-TE$2)RSZVY?,=,-+,@DDM., 
@[#FE]"V=,'@:T,^U3B;79!\OM<[2)(/K*^S>--<%A+, 
@@KF^R"#\YV;40QB#-DUMW^HJA"6](BGI]6A++EBE8B@ 
@0'<D#9)[8O[GC+$_L'"@;ZS:KU;]J\&%?EV6U%D?ZMT 
@$+GC$&V>4_H35'Q7/Y\.R[=[NKW;P!@SV5>VLTZ+0UX 
@N$W!;SQ%H"YG7Y=60^TD:"$[SN@J3/^ U6?O,%:>*N8 
@Q;LMB[2,A%6.X>9.<N+;3])0-'$,[U;"HVT*92M;@Y4 
@KV(_&)&7+::Z5=<5?J%0G:==VRBQ6#\MK@98L".=NOT 
@.Y<6I(8M39ZK+Z!AEY--K!^IXT-.WLN,73UW'CF[Z9( 
@S[ EI0N$3/$A/5"&W"6BV/.%N-:.'W\"CW,^5[,S3]H 
@O?$OV:!,9O2>!&QE"5NY9]X,W&^H(6T*?S@K'LH<XR0 
@D4S//""RS-K@I"=+1RIQ84!G'29I)Z8M)RH!G'KY[>( 
@&P,VQHF!=1P1AT,=QCH;Z28S'68!EKQ-,FQ>SIOUZX, 
@R9LGKK%7&[3Q#Y, ^*=MV+Q?3S_78R9'/,/"A4]8*JD 
@GBU5MD__:[[)XI-Y1;*!"!K,=%BX=EUHB'KCGOPQA40 
@BFK%NJQ^GUA?;;/OJ9AH/B#X9&L'PN[*:=&&P"1$'ZT 
@#0KDR;<+7&*>SMF=/ 0SA#ITB//Y9J9_@M435*9R$AP 
@%1W,Y%[33<36GUMFLLYNM@ZDNB+67798H[T< WYT8LT 
@,V#&FF(R"MJ@QI/HG><!AEG5*>N1FEPMS"*C-X-]QUX 
@N@8U+SI.&Z@NKB?SE4,B78_*"DA<E1<M90^- _2=?!P 
@]#32ZST[_C&(M)^CH04$<[!D=YP3!CHFW_/8+A@)U4H 
@KH)) >2T&0:!F6*@&X^[GM>")926F%^1#J )-RY2%@  
@ISRPW)6#@]8H*/"2&B/(2)MVE-B:U2@+,[((">BN7_$ 
@8$.]PUJJ=;SRSXB&+'UC.6R-RH[9#?Z7H7;"W'%,V,< 
@Y%0D_<Y3I&-HR[=_D<=WX^:60+&VU"/N4JF24>>M7Y( 
@VY'_CM*1!P#S[:QAU0=#*IW8]L&&R\7_1$]P4JA?@%  
@%A@V9R('"&R;:4S3T*]][D55P_1L\TG%!Q)U)./\6$P 
@X3/K6_PUPB?XAP\YJ%J]E@4]:H&\D>Y*W9]Z%K_>#3< 
@'702*T,!)1- XYK[3$R47&U&4?A#NFDT;#'PZ]_^W.$ 
@(W.9H03"[/&TED\ ?LW&/@WJGI5;?G76%,'ID?Y@[QT 
@0'Z-*+H"V\GXL?##$_SAB\DY]IW^KP0@4'7$__*?<$L 
@."9P5K$%^SVYKU1-R?<?>D!8U8H0L%'<@'XZLW&C^6H 
@TDFQ% XH8'C/=(LKYS2,C^>E^GV@5GLG%8R&!;D*M2T 
@*7L\?L<35/6EM#/=]]L>]Q2QYY/'J]D!5^]98*R4;>( 
@=&.UA'5^5Q[&:%-CA17C_BPK6**)QZ>RKYA11#5F=:, 
@B_U\>@&(<=GMD,":0J*=/U&:JL"\&-[4$81/!H"#J3  
@%0'2W4_*VG)SE_O<#-]CO&1@OF>A/E_??YROS#V&*YD 
@V7V$R+/%+1G>V(L'&Q,IPB(4^GKF+GD-<7VF[ ]@+"X 
@+(7KC_1:2'!GG_+BQ.VUZNK) _V\9J9A<,V3%D=T1/X 
@9K]<D)F";Z?;+M:K%@@].!54?.J +ZJ$M\(1V=#7,Y$ 
@I9*.'HC[@HN)S9A5:=8T3I\*3^J2J9P;9/**419&V<, 
@YIB1$1N:>=&] 94M!@$T""<))]#,KFW<^X&H.?([W*X 
@\?'<@X;#4Y+*\(&/^)^C'D'4%8O88(;-U=VG^O"77PP 
@^I]5ESOZL.J$=[D=CA.(BN;WXT[]]A]=K2-I[A#^-Y  
@@U^<7434NY45\D>>P?'$>1%I<88D7T>S*FP1)KO)72H 
@F3J="=%HR?(:;I8(W _,<,PQ&[VI>T+U<EECGC>)0;0 
@PN9L9?P%T<LA988F>R]^)=_MNRL-H"C&>D>.%,\V2(X 
@MXG/[_NO6P@,M&/36I6:W8T>EPGPCP&GR$GTA(!G+<X 
@2OSW<MDNE@);TS:9<N\Q>6E\'8?="2.^J]E#)_Y W,, 
@/IYW/WN*;8Z;%<EBH\1CA&3!7\#,EW$E1""SL7AYFYX 
@+TDU% 0PS;Y(WT<=!4IZJB]%A-KR*1)7A(G*'TL@E L 
@OV%O,UJ4M^7RLMVP4"!.JKB5$QH(A?UEN'FL4L]RL@D 
@@5>/-FX7[5_0,Y8U!-L-+:M*$O^T]9L@J$N,#TK2D34 
@\]U1OHWBC:TSP'JKN4&-W$82[U!SNP*%'KPJ(T3+\TH 
@6H+#$:QR2-@KS*E_:3?/951''E^:)F21$KC&6[ASXC< 
@,.[^:@#4MT::_B"63@XATPF%:%H$X8<S(8Y<#1$IV(, 
@1 JLG8>E(97$\X!']]$?M$@M\VK][?;H8,F0!1C*C$8 
@#OF<SX1Q1[FA/XKF*Z=<3RCF!G@.+L*/RK<P/ '7Y:@ 
@.1T5"))*V3,SK-+8F^1B^CJR?1E2Q&#ST@$EO!4_^W( 
@9O#_8XJ+^Q4077'".-X.I[X$I@/+5-)/C'L\!%\C*#@ 
@VUQF+Z4,L/6+5"^PN> B7O&:DAL<P)&4 /V@N N0$%  
@N='91/?JC&%-%%XLHF,/R_X)(_AQWPMW8UY)D.^B;.D 
@\YD6=[J(M'8<V=R/#Y3& 3O$<&M84FO!1'_Y  27E;, 
@^$ILP4\^LTLDU'F-UGW2PJ+%-$?;6TKSS+>WD*TQBI\ 
@@1#C6G;T$G4H#2?+F*C;5T?,\;(+&^%)U@ND!*]M0JX 
@'PU\D,AB-3$9]H$9L4/& &9J_Y&OKKI9H0#D!K%!0@8 
@7Y&XT24]>82M%"(#ZC?47P9_GC)A<RB2C$W,J\^"L"< 
@1P;UQPE*K+*6\ 4:I740<&(4XTZ8JF<\V&)7C3C??C4 
@38>=4W5_YKY$:QHO20W*&B ULN^]\S3F&+:+I]M@%&D 
@DAC"D#'IZ;[,0#5O(.V6JTB\!,$X&DMW.,T"%_:0YV< 
@ZK086,36N&TOG->"S#&&!) +:64$1)=TV.8-T$T15J( 
@&>V(=5+;2GT #\KJYSJX[1O_4NT+DO2>61<-B. 0M44 
@CON<^_IQ)YDFXOB(,)S-WL=B&,(^O!VO_<D^9GW=*1  
@.O&QK8/KM.RNXBM?CUBZ!:J?!!Z,_.">BC=XWPM^;@0 
@C=L++U] QL]S.E_32[[USF I;R-A &9<D/1]":J$O5D 
@XVY;J3FITO'42($\?WNO%6'<<M"-GEL7%3K ]8W3<4P 
@J;1!7:2%CY=9867V=UZU"*YO-RVR:B4!&!F]F;''*^@ 
@I^]Y[!LO4ZB;*$;=T<S"B;0-E@47H,R]#6(I&!"=ZUX 
@Z+7#5K6PP@4^);W6>12RQRQ!.I.(;>)Z&=RKG*<)A"L 
@/>5(\&Z5)^CZ-@.5)=]3D@GCY@$AO>49Q[!+!ZN*\8\ 
@EFVC3:N?O^ ?'13:2^XBW E2U/#RN"3VP0L3R+U"-X< 
@ I] :#9-STDUZ^(5!<(JAB%_3Z@2->3";3,%URTII3  
@XMK2E"QF.]$<]1#'(_=&V;;[-'DFKN>BH;E,7"P\8>0 
@VWQ!/*[=0\O_EB!2VDWN;(\?23P(KGQD##(FJR>^-.$ 
@H;GJ/O_!.LW% B*EY/")>QW6X$:BN5J'&7DJ*YAC$^4 
@-2\CK.NQ[,%5P/3B9CB_'<X1RS 7C#K M$K"73;O'/X 
@BBU=L\7@]X7YN3!0'7OW6_M%,@7E]30+' "EFB4*HAX 
@",AE^"SB4D/D7WB<^_WM%:1"9(JXP>6A/ID-O?_0Y'< 
@WOD&32-"/5B.1\Q5]=W#WIG!;2!)Z0(85L64[> D,EL 
@J',&NW(B:M'V5[#.B$7F$"I6AMU;Q/"CZ<+*\RZF2)  
@@4:<>1(X;_ $H[ (10J]5_M/]RD6E22$EC@!_E*)+&, 
@,+0!M!KW3Y,] SMBM2= P7M]$E]#2.+LSX!2] 5,N2L 
@9-SA8K-.]5NNE_G_3_I#W(_.%M"[$NUSM<\S0T7MZ:< 
@&ZV)6#HFT(K*=:_G)$XZVU;>'/#O(+4,)SGTNCMFQ7X 
@159FI1D6$7WH1YE;HCA<O$Q1Q1#=\N\YEHP4>/E<Q@  
@9*>:LQ$OQ+^Q"MBD;,#1^WV^G(4"_7@')NR-I#%7EPD 
@_I"A1&]YQ?)N?N^-SBB^X(95<_@9N?HSKCW3"@165$  
@-E&D1(6#7\QW81BM+;K"<PZ]QSI#7S^W.8S_::\025T 
@DDZ*NAC8-NEDNE2-"6ZE](=54OS"+0$ CBJC8.9H1'4 
@B?S/ PVJ\R0M%"X2P&E[Y7[+,ENV]$Y0>[2Q+A\1!)D 
@=6'[/K923 >F$_O^D?GW^/]IB\MQ<N9Z8WBZ#6,OO$$ 
@#T]I>0I:[-#!9]S5U>S?NI)6S=ZZR=,+1ZH &K,U9E8 
@A3S>0Z;GV95Z^KZ&LF1C6H^IZIG-'!J=J)7=Y2+B#;D 
@0*C*1/\"XJ^:!\T&_&5N3V3LPN4;NJ.4CN9E\Z*O?V( 
@0U$01OF(]AGS/GLSCTKEWI6U)IECIGP53L64YM@OVV8 
@?J24<BGUZ[#6 / :,Y"%RS%0]P.^RW _)#5-,S&--=8 
@(9!:+)^3'&<VJZ+03/^2B2JX>C*2K;1S7KP?3,:QF_H 
@G9!#8>F&'HXH;- DB8-:Y1I/ZI&/PX,:F'N'.6##3R( 
@.$TN%OIJ\:K[.SY7!S +D[WW-&$YXA[T"Q#%?_+3K=, 
@5I<%!UHH][TK2>,NO#2(R/ #D0C1NX7[N3>\?]V"O$@ 
@=7SJO\)G::K)$Q$I_E'TJ,8OW(QZL;F0\WGMA^>+%W( 
@B=3_>&D7ZN(SNJ'KCZ8&"?8$/B,3IQK_LK3H%,*67P0 
@FBV@W-!50#X]G3U#6Z0X M9O382O3?.O5&7)PQ,U><@ 
@Q80AEQI.:X%7<JH#B*\#VN&)SVY%-VWR>H@C]'_$!40 
@O=2&#I5J^)=%>Y=_)?*ZD>'5NRU_7\U_8N8;G+V=P6$ 
@8@8Z^"H@[5%:Z[7)>Q1>;&K@"4@DRM^;:>NSY]?L%7H 
@X%PAG_PS)^<*=7*U1;@'A5UY-T]LH3&''NXTQP^6C@$ 
@1D*<ZHV:(,N7P!%>@:-*UWY?%0C6$D]@=?J52#0?!'0 
@!P0<Y/-73VMF6XM!/8I[XZ47&U5!X!X<PB-X.[JC/5T 
@I=;"(4X&ES9993]A=TM![#UKGTOO<?F+3/+:!VXN;$\ 
@EA(3@1S98VB5E7O[3]#*M8G\*<#8?=4!X%>(FG*598\ 
@==;^KR;T[H=-,V_0TKH;=TK-F5^%"Y6K^TA8KCR&BLL 
@A@-B.RO+[Y4R]\W*4+(V!F,<$O[VOZT;A*PKS."ZD/4 
@*W\Q9?]_+\?(U%,6C<6R"7PW9JUR9),4 \W4F0I>7;\ 
@K';LA>0O#"?QWI!/R#0S'I7%":F[%U2W'W8+9RJZQBT 
@C4*W(\I_CQ9?,XK992H4NS;!\5/!BPB1Y*I?M-4=7#T 
@AGEJJ>^Q?X_2K,+WL6")N2Y7*<).4SN79!YMTE8&@/\ 
@[#04OOKBP\ LDXVQ&1\H>K(EA[WX#X(E4<*76"BK Q8 
@VX#$>W+9X48"6\NJ")C"%A4&LJ%8"0E)\<#!^-#=-!4 
@*J$.UGW@A6&D\XSP7GYA8?EAM5"A),:TKRW>WZMM<KT 
@!Q$@DP#JRT]+.FF]K#??9GMP_("OM2DX*X+JG?2Y\>H 
@>K_/%U[<I*QHHESV@%D'%7G@W(YB412[=5T]:8^@@]H 
@<P^I+8"B<IX%<>5A4P;+/F"=\ 7/(>G!6=">0"7T/,( 
@N<?FV)%89VN^*^.$*.?!'67=T6!Y'-4 _U1=T.]S/(0 
@EH%<#E;?-#Z5]GNGW;MQF-<=((4+].!4&E:Q%H&=M9L 
@+B!QE&&.8__PMQ7<HG6=.%7D(PO?<?J=PO$KN("D,AT 
@-.:[21PH#K$_9J?XA NT"PWZCS-\I.>I'4G#O#[.F2, 
@%  UX]D%ZK'6&&X:H5&4TU>:UWI M%]-;.31:^<\'18 
@Y.5NV,1PKX6>E;!09WUB6+JN;'87F.GQRF&'"B^SM 4 
@_<$P35!]F@,QX:8S1+&'W,:OWF]?//4.W*J> 9WM<E( 
@J./<&LLRDY7Z+X'/$D!^-\.><3C@CC\E[8<UT^U&,DL 
@_ 0!G[&[.J9&98/T 1+NE:P$!CLU<3A,>8I#B^>2 M$ 
@>-4;7_>/ZE%G UO2TKHK)L#L7KH]^+#-GBX=IY=3<6< 
@HY3U641+2#I[4%5.AFK#5><V^2:;OLQ<[!.UYMQ.;#L 
@T$4T<RNY\QR@7&>^?IJ;.3LE-(=CH+VP[81''47T! < 
@R=@TRPKRWY/!LE[ -G*V)A/KLD1Z@QA#1W9JZZP/,B0 
@6UTA;<Y9<A?<4WV+%N3.U'"/Y.W%4.<XZDFG^4EV>@D 
@:&QX%/?0=/(-5$I62BCY+%U ON.Z#WZL]M::06Z,3(, 
@/B=JKME.': 4#: 3E*+4XQLLO:;CFQ? VVF00RQ&5FL 
@,DI]PDI5,]QLX$A9P!LDO[ Y#VQ\DN.!M\8RE-3?14L 
@U.C!L?*I0G[9H?1='W(=I@JW<XP4G,M3UZ?RU4V>'#$ 
@'G]"-EL:C%<#_U-./ZC1BD.^:"AY98^>MZ..OSTB;M4 
@F00U"7S5ZO=*F)DH;]>-D)&I,I?%N"S52,?<2"3%(P4 
@E ?PWHPW[S*UD=CQ?\#(2[ Q.-:)7L(F,[+!03EX1DL 
@ 1I$09!_$H&C>BHRD0E51D"X'B8J0WB,+?SX]&Q#^ \ 
@8?W!=HZ(SWDLVU?&>(D(5(OOHB*8[ 2M1->>6MB;<BL 
@8RQNN8@>0JB3PT&D 1F5N:SS$4B/]4PJA=[&/Q7[*0< 
0=!:/ HJK3"X%G:U>U!5F5@  
0J@5@KE 3G8TAW?29'DX;?@  
`pragma protect end_protected
