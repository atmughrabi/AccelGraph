// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H&(T&P0E-P!>YM"[_H7;!QD542!M]8NA5!&'WR'4+OQ'"HI.PJ-GD60  
HE6]#2^!(XVJWP6N./3L6.$K29U(AY0QI_7&^E0IO>M1;KE#W;HI(:@  
H[2XR(D2]YV(U1=#B8HM\\4+^U=T^$3XT;59JIAM^)ABHBEWF*Z_=8   
HXV4%CA %#_M+1+"'$7=G1]-ZD?X:WA?^/@1K4_*"'GF V0[*UNJ!+0  
H49&'/HD;'<9/8[%VXR>1$&#^<]6QT0=]AC+ST0J!!OA,/WQYE;P29   
`pragma protect encoding=(enctype="uuencode",bytes=18032       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@HX9^C2*H9:\[-55HMY@&^5Q>$\*+@"%S,UGYL1J8G'8 
@*SE[%>RWLF='8:8T/Z5+)WG(2QV7BSK0>B#1S$3^^.< 
@5#<.P.]+4(^3 (7U!?UQ 4(+G^DMI_6R2:'TUT$*J9@ 
@C*[5Q69'1D^RP<>SF'=O;&LX1SLJ#5N$).8$X(9S#=@ 
@%^F=J157^EX3035A"5\+.CGZJHED+T^M@:<MZ6A#25X 
@/ 78@9H*?Q%;TQ@&?QJOKF;VH#98U^HI720L!X[D%6\ 
@/([*)M(#_&=VH(1GNSOKR7:B O'>^+?*%5OD][CY8A  
@,KHN[2H)_G&3A6AH]HOTALY5=S#$!._*ZMK.J5R$BGD 
@73*]2C(JP.3UWXS%<Y&JE'YS,VS]^N.<Z=U5OS!_?6D 
@1*EG8,;P$U?AU9ZAT<5.*'G@P4W057ZC^E'!.,<^?A8 
@CPU\].T2+99)D.^E$8I"GY9,V:.S]!38 "FA^G2O*E  
@6-VO=7E:0Q "/8<5 COSGE,9MX5/K*O-A!/L1RK,H88 
@GAU'KDZF(]/.8/"&NPG!#,G<R;ZGX)\9O5RHX4U0PEP 
@^I5BR[-$,5XEM;PCB@1856&"&>853(#^_#]G"8:.N 8 
@3K<<LTC'"L[N-SB*!YP;Z4W/W[1PPK:YXFI]ZJE@.T\ 
@*24KC6E6M"RN1%;^CY>$1_$ZCW)<E%TF7!E\_/'%4S( 
@.OUIMCL\D<(^(DUS4S_J) 'Y4FZU)R4+2(J$K:J+Y6L 
@)J8Y'U;2;TEJW*$<?+O"N],W40ZQ?>UTKX09DS$^)C, 
@:5^N6 36#;3S%E^8]"3K.(1AW),-2_L.M398_&XR5C@ 
@\8:5/#D@0K?P=JEOZUSTMA!4&DJ%1DAV:\4VGX+%B!$ 
@&32>D T?21QD=*9C*'Q"VV\EQ'L#KE:Y>XE*'0,=Y\T 
@@]'CH4QZ7-3O%D7C-@H?:TV>[U,F?N2U#RDC\BH9 BH 
@5^NHHNE*DS:ZUE:.Y&R,0FHFV'2<#V1J^4.!ZL=-[(L 
@QQ_^'=G4<0$Y[ 2GY780 &L+[$'5A65VN0/1J*EZY@8 
@=LMU@NHS,+VEG\?3A_Y'=:XT(PMVV'M:<M;3-E9_?@, 
@"UCE_5BPA#DO#!&,T73]3J6UVZIF(C)H>!NT*$C'D]L 
@RI5 <<9E^RJ9MUB+.#D.5T**R^H[A%..U%U[V#!TBSX 
@ L[4C8_:F&_ N:US//2[0)MG&\:%H,I "9(-JZOY0M8 
@ZFCK(Z6+GEC^O 3$X$;"Q(>1+OXQ4CF.ZFO\'SS??G  
@T8W:.,SDI+.4E\%@5C,$,A_E\BJ%])2==92?_ZZ+@FP 
@H3K.VZ!HHQ5;J7I!N%3241,%TWAXWIT!_9J>4P%F3:H 
@[7H)]3Z]Z=+[VZE(B$7K:7XFC6T0.6OH6O1DS3Z(W=( 
@" \T7XQ4? Y"9^ 5\$!E7Q?!"@_9@+71940O>SGDG<( 
@ U^-Z1 47LVB@4I9KHGOHW&JY!<@*UNE4G^V?/I /Z< 
@I?<):R)?%HVBI3(J=G>NV-?@#'_0^'"-8J,73L/^CS8 
@/S7A R1_H^VVA0BM>GYJV#%^#JYIFX<BZ))PL$=D2Q$ 
@A)L2X*#M>;U!@&@3S^E!I^, *MV6>?^@XOY5I3N)X(< 
@VKL2O1D19-4,9<?B]&X]'*#+,(3!2CSG=1EX_851X08 
@&<S%G]$0M<(A>AT$7%/,S1(I2WX0-D2$ 47[%7(!!>$ 
@%1&XQ*W\US6LG)U0G,4B(2X 5M]Y!'IN]VR'L$_=)VH 
@0CV\4_IG-?+' EFV.M8;Q_D]O*81X$?-FW:OPPMY9=@ 
@) +T%UK109Q>=%8-8!G3"0QAQ4A#--<6V<U,].L[HZP 
@YP8Y$*6CH%)!=8[U4F=P\J[59#C5_9""E#BAE'LNU=T 
@T<A>IB#&1K]#FMOMOK!H!*SE*0N8GA\7A;>)\ZUG*A$ 
@'E@Q>396OAG.M4#XS]2+1-L+U&<34:S+Q7OPUBQN3RP 
@A8U]C=+I3;41(ZS#)VKO3?1^/5!49R&CCM#%R(02C!@ 
@PVALEZH_1]8-ZTI[@#QR,.R@\)I6,*2:>$QQ3;@(7D4 
@(5N4B@+.X6C(ZB1WK'?\7]D<ZD9,H;D!,$+#(8CT'7< 
@C;\YRQ^'1?+QYDOMD.:2-+%^JNV?WQXG,->1>;6FI/< 
@,YQ9"?7<!O7!^GFX0/QF#]ND7TK>LC9^FW+,:GR9@ZX 
@$=(KIAAO:MZ!Z>&5" C.1MU@4F+? \L'X:$G\A4T%1X 
@FYI7YU57H6'^XG[.T%)B(S"#9#9FHS<5AF1OBFP'K$< 
@,PW]A%G3Q\<\>E_W_(,@H_[?(ZOW )4D ##I)WSY7YD 
@YVTZU/IU'7 B?H*</3UQ3V+Z>+AM:I.F>1KL [(.PX( 
@7YN)??AZ)Y/=C+P]E_'ZC#]C<79%_ U+UKN52X)U1?@ 
@4J,B,V^W%$AH8BPFSI$$(U[,K4=XY\7\D*;<_687U4\ 
@;EI<'E9;_\&U(AVH7T">P* L$GT?MWAY<:U0)-OQ7H0 
@IYK)L,^PR)/P=ND(-MS[WKWI/^0['%^S=>;1I]Z-Z%0 
@\;*5#TU4"6!11[\]PT'XQ,W%Z@M4+MVR<(!!QF^7D^@ 
@;[.GS+KX&1 WE(&!F-0ZBA3QA0I_)95&AGRQ=A\/K!  
@@TP2NN@LCM*ZE"N-_/O(;0H;77!)</REMO;Q2:'Y(18 
@R2HI:2K4Y[1<[]7VL?RZDF43VKS"8ZZ9#QI!BUE3ZK< 
@K24%-MU5M'R,;7B@+):HK8"\;<05IZ5\+^ 0,Z!B _@ 
@;$<\LSZA5KABGQ2C;"$6A \DU\<0V%7@;2;>LH@:!54 
@K[$Q233::1MWI 18V9&6K;),/F,;9,?IXPI,83^JUHT 
@ALU_XT>]"_K=-;/GK/UG@'-YSFC$!"!Q+J*58]C,V+X 
@N6UJ:]*X%0_#"G0O*OD<'6"".^XC+<$7\>XJR$Y!S5L 
@5YHT@'_.=$?\UQD99-[1D[UNM0^PA2_@I?: 0S-Q/]L 
@[K=SEHN/)-LAEC"NFM@$).KG(J^5&B_#TODT1^%SS4X 
@#V=),_38Z_!#BE" +;Y]CMYYQ,K#A(0R;48/$7Y0W D 
@4S;_EF-"H+[S S473!NC ,.$X^>%/;LEW:PVM%IF([  
@7RK'+FM\?K(_ELV?D)^W"CFEU.Q3KS6X32(]6*7GIZD 
@+-8S6[4P25O@[DO.??3_7(-WCL50.?.%NSANRT6&S=@ 
@6"<S(EJJ6&=B2PD35&+-+P-U'0F[U@)'4:N\]ZZ\ST, 
@01QG:N1,TJ'&E3GRF4D2=OG,H":[Y_!P=<;A["Z].+0 
@/IK"XV_0L]Z5#W$LND8J^!XPKB9>&4'*Z+%])V =!^@ 
@VS$FV%.&5"W-  :UM\+(4*S[(8)N:<8!M4LL[@CB^,H 
@*])$>L$Z/-YSEB'1&KU?$!KMYF<@W(A%34;/EP.W-@< 
@Q84@H8,K,[[$R79N=I6.HH$ @7J9[%8PX1+B**3OW=@ 
@-&801DSTZ74#4U%7TW4], ^:F<CHC$U(<J'Z,%?!_.4 
@#ZYLD$-R;Z/?& SM7LJ6?U88NPNQ!(?)94?/20>=W 8 
@!D3 .NVO&L[MFRRGNL"FE=3YB.X*4%D9-N-BWN!.))  
@A*?E 06>\_ *A^XRQFC(\]*^CW6SKT]6\-J]T', ??D 
@9V].[\ <#RMN/LMHP7?Z\OQ6)'#9-GJW/!.W??,?PS@ 
@3M23OSM$Z *%K;[Y-8<G8G8MYRK</0Q_R@,;7H^/1G8 
@6_Z88<B^T/2"[0$<0P#@KAA#]=29H J#&--KQU*,GJ\ 
@R4LHF[^-R^Q^+2!"732AF&*C+T,'HWC>=6?Q&64%<8P 
@6]E[HJBE@J=6@K$J0)9EN>1W691*@7TQUG$5IR2"E>P 
@I6H9+G8[LD3+O3(@_,"=1&VS K5C](S'27;=R*)2TM@ 
@MIM@7EN8?NR#RXL$-=($.:SZ)X4+^<N@JU+HBS4-Q>T 
@^OI^?L!H$S=3%RG9IS_Z'_,ENXDMD#IG*B,49L'5+%( 
@/3T2[6^?F(5US(6:EV@PM@(.E*GPP!SYG>JE:-O@ B0 
@0A-RVO]YW.<WN^V([YQTNY*A;"%<J)?:#>K+HSWE.AX 
@!ZP'.7DW3?9$@L5T!"VZ/L8/Y!JZW69OI[V3^IQ%?I0 
@=^)5V1/'5QWH@V;DQ&CALQ0+WBL;Y_8>;9#@%2/P#7@ 
@G_;\3R05$T7S@GG,&(5,5C.U*9ICZ5'\:+4SDC,7L1\ 
@%O:URIS<PX5&ZHBHA 0MZ;DS7T((B[&@4,;B+4S])2H 
@2&.KG U/T8^')(VN]2>T%?;5 OF<65I%LM8_.G<,U"0 
@$AVJ#;B;53*.>R17T% 1R!X!%$:W8[2C%XY.OZNT)'X 
@&M7RB!4 9]1!V+?\FH5KBH*#"VFX*+]>Q S!<URJ.'( 
@Q]>)=S-1N>ECV3HYYQ$B6'2#@M:*P[$? Z,D=Q;T%(@ 
@C+B=,!I9":=5V'$FM&%= 0T^?\-W1GHA-,%_@85'CPD 
@_,R'0XI*ZC]\4@%1QG%7YDCIJAR!5&G/J,):%6,,S<\ 
@[02<XTH4K]:]9[W2DQ@<5Y^X_(E-8*&-XP2*:&I!_%( 
@+E(3LWJ=8H'5!;Z@[OTG!8=-)[X/^5;<7T'UT\0 Q=4 
@@V[W$$]?<8OAK9.).D##+D] IRIQ_3<8$0=QRBK)MZ0 
@T I)Z%5QRS^DI6!:,5V+-6DX%28XD! 'Q<EOPE)DFI, 
@6<B\&/R@$'XD/T2O6+W5%5"W@+ 9M^]X[PXPR#C5IDD 
@.?;B0^B2MJM<36V"G_E(&0&RM/C??%$#H=]]Y2L0KY@ 
@J;CPV=9@?Z,#Y"E^A,:OTOT&_S&4F')!L2!<XV5*FL4 
@E8E0T GQ,ZF?58S"0/_*>3"'U<"T[M=B?=<AF.E5P@T 
@R.:[U&8N1,Z8Z75]X6I!@H4K:P>=DT--MB,%#$,S!$L 
@;K5&4V*XXJE'!TY^L)>.[21OX5UL+XFFS%X;'7KVTL4 
@Q8J[&=*I$0@1)!M@#6!Z=ZA'77;NL!F)TN(9X4UHE0@ 
@WNI:V9<EQ;@D0^UA%[O>%+N[<&910Z)73-CN23LSHZ< 
@DKX2I76J*'?%?(Y,"H)#>Z@'1MM[Q!=S-[%R#_(/5[P 
@=JR#[MX=3JB60*\JD"UM8;Q?7V9NM['6\W4]CN?,VXX 
@S5L6U%.A@/5V6H+&AVU@^@=OIA";I."(U_Q7Z?#P%!T 
@7GY18EKRI;\$=NL:F0ZPM?8:5^_975?45W#ACN3:H(\ 
@$.6E,!&'86GD/$YZ:S/+&%.[UGPQE5@N3V#F=?9 <_H 
@E_M27@7[*C0"44C#];RQO=F*-#S6TWKTP)&X959,=?T 
@>4&U\'*.URZ %O@5G+;($1N9#$M,I%'*8+W2CM0$9Q8 
@&UI;?V=2$? .-;HN(0YM2_-&WJXD!0HSU][?YC^?"$P 
@!AY&+Z73,90[5#U"V@Z ]$S:U6(">\*H^6)BG8;R*E@ 
@Z[!=MT#9P809?W8$="6AR*.H9:TN3,C$QFB4@YM=.1, 
@VY9&M\])/*SVY=8"7!KU251=:SEM:00'@[38"8M,U"T 
@;&^CJE)92=?Q\1PM2]R*^3Q9 Q/:!I;YWNPJRC_<$!X 
@X(04T;[EHGI21:(P5X:%S.1[EUI5Y&[?N&>2) B #S8 
@%CELZ#^78L PBE8058GMH>PQ1BV-<C1H0+!=H&&DX$$ 
@Y&4L+^Z*B$"8I4QRK>^?7C0S?QY>U71^/+TCL33/*.0 
@AG%*?XY%.W#B!6;"2=WEW\\'GBG=^2^T4XY[\O(POWH 
@?"&P?>#./OQ$C6X1507YM'#&M.Y*HUV6SDCD/ZW*2XX 
@FVRH/K/[HT#*-UF"&4-T,OC_G9"D'=X4"0E<M,C57$P 
@1 5")5XZ7:!FS7?0()+O%VGS3!<?O;YEY?UR30!X:RT 
@V@3"T%R1\N1.U%[]1:+))\0*W6C:(G-%L:BHPN&\C_P 
@.5]E'&^ !@U:LQTA4+WD<P5[J.G /TD0HY>GLH\0%GT 
@N$8@^TG^T/OMMFX>RR\I:+2;33\?4P7LJA_>DSG3C[H 
@@$6L6F0S*%C#B6^W5+M!V+,B?,?&9O,XQ0-4.$N73#P 
@8"M?/YGSBY@67;/'HD#<C=G9\A]= K\,.X^'B=%LY#0 
@'JC%[2Z]@DZ1\L7T%<?![(\<6T5I+)XMB8)L_6G\!0( 
@I]> M-?FSEX>4>^:4T,<8 [F AWZ7W,R_362IOITG[< 
@ZNH8\,8:S+'.0]0#=I8NJ[\A 73H,P^E[O3*\!Y4!+, 
@-+*ZKG>Z@#G@>7!MZIN9/:,W*OOOJ[E(D*"#MXEL83  
@;$3&-E8=W83%T,%Y:84),>-+L #KC7R]['\C<5SH']H 
@L5<A@/W><Z3R'A(1LWQ?2WZG.2\,3KQ,FN[@Q5_JVGD 
@E$=/O3F-"YXS>$4R'[RO@XG'5+&LD ;@)<,,JK(9;OH 
@UP SL'>QCM]$ZZF]$4-?@V]C:!%&H=LVY^MDO\Z\':, 
@:2SYV:-TJN9/MOI-"<UCG/P  V&5B=.],:95Y=V?U;, 
@ 5@LPW8$A+/<N?&4MV\&" 'T(KP<ESODN9NA*JA\;X\ 
@5B,Z(\V&?41SD)ML9,JD 03"9]JPPD33;V("@&N"!*\ 
@UT^]82_M=A[:<[$T&4.Z?+>V:6FB\O!2/SMBN!M]8;\ 
@]W2\@CB$9;F+IH$K!TEK.P5J!O6#-@CE)[Q[!B#N:I$ 
@"BOG,W)80]^S\N<0Q+G[*$P-:]2:3.^L>!IW^GI0)_X 
@Y7B<SI_G]LML.<YUT]L3XK-O7Y!)5RR19!NS=II='6, 
@!VS$KYBVI!9_(Y_@._6@H5]2 '3UE,R,E*ZU[[?K&KD 
@U:\,[OJ#-HQW5?F:T'FB7S%NX3HHQ,&J&/3L6,S1/'< 
@!"V?B/.>Z[4O+$Z;Z5K^W&I\(<^$ZJ$,906AWB;&^L( 
@&*NE*A[.GJ'8IM'@7?E U<E6@4O\/T-YWYL,SU),28X 
@1IG3!*N<#6:#2-6^9[!X*3?4-.!#'DUJ!33IBN%F6@$ 
@<##L-?O 2W;EUB29B\49UW9FVJDA-"JA)BY45S=!Y*0 
@!#BY;$3WI"C8?#Y/_;\!]SG.6'8>#GUU7U4B?:B'-48 
@V6!13E<BTM9:R<"N/VF<\+4P?3A$IY$2YV/_$#'-'_H 
@+K'K!YLUN7\,4R312TDI8'N'-FJS-#(F)$VZV6M.K'< 
@"&UK4S1Q%@/I]32>=-%Q=")V+MDMNQOQ@]PNX LS"6T 
@X0DOHE766!MQHQG*C/_JK5$_#5CIZB!QVP!\Y\4TR0X 
@_&#^'Q\IT<LH+?'B]:N?FA;'>(/A[X>"\Y0/U\;R&>< 
@^2I+,+4W_?#W^Q&U*7.=2V!TW/,>CS*)@<N!V4:?L+, 
@^A"]0.0<)((V6(KQ01*3=4S0XXB6'"_9Q/-=\5A+AU< 
@!B7!#!BQL#;6%WE3G,I;(%RSOD.\F@W/SAJB8R_2RF4 
@M38&J[@%P#%[:'!DKO8_5P@%XS)\&'S0RNUX6WBPA@8 
@Y8.*Z*5&J\*>(S B=,U=-I#(9Q"D?0\UB]H;9R?T\,X 
@%%R(B2>%9P=0U6S*;_#;W>V#04ALXLJY[N!$&>I"2JH 
@)90$+2=05*(RDFX!G$>[&O%%KHHF\:VT^_;OR C9SNL 
@UR/>W5J@\"N2/2/\7FS C:M;$!M\ (\%=MH)27 #4"X 
@-%WLX*'9B#?-1J\IKWPS"C(*X;X1?!KEUNBW5S7"SAP 
@H:FK*)[(-'Z)%)%F[,,SQ>KC@"1!VW4C#MB\/]":G*$ 
@HGX(A%1S<21Z1[ZF<6X9&$7,HEHD;_EDR&TNS-8>U,@ 
@P2A8 !_R*&3)*\V_'$KB>JNGY5P*\I8M%&VP6F:6F;H 
@NRZ[:6/7;JF-1S7F/&4[=8W]353<M3R7=:$X31F6(6< 
@_I::_31RI'H8 @3"ND97X3H<*7TT8/2=;H/:V@Q;1AL 
@*P#<@X#I7H. ;AC70AK6Y9#U4@]$KQ/G#ENITZ_F>U< 
@)\=A"2M#6W1=9O :*J-6N-3C+]!T0;&FF+KYOJ,Q;K$ 
@$-WUE2J'\_Q>A[PLP)RY4LBV?7/W*@;E5][6(^.7&/X 
@/,>T./E *,M' @ H D:2QZ>!]%ENFM@ZAK/O%D'4J.0 
@X&(B9N\(P2!VU]..R*WOX&]=N\*M0GG)&2H@,3=,ZO  
@:M3UW0 \G-TQ"5X76]8IQI)*AXUK#G1&T7KNL.#E.D, 
@6&-Y1,1W?_6%<:]ZK+3*MZMP2A1T[NG#,[@B<!;/_3T 
@E28;0V2%1CRPS+U5_\9$VU9$-=!G0&NR]40T@*=X]?P 
@6<?#P40FD'2#":D3- X._H@N2B04%!MM%E*&TOG7SV\ 
@C$NF*F=YL&#J37S!NZ0^0R_20@)IP'?!0/>^F1%^5OX 
@JXS$O?U+2NVU];YD-?[8,*:NZY! X[1ZB)OC%]0YW(T 
@M,K1H$440^N%9GE;$V+Y! ]FF>2P;)T.T@A%^./N2GP 
@LHYEMN?6,FEH20YD.IR.4;(5YJ\5 ,"X>WJ@WFW?8^X 
@B?F\#\$5TPTS!MV<Y4/DB7!0#@#%N8J #(BQRTUBQFP 
@C)5AD>V *K1=:PF2W X5?)AK2G F*D(\-4B,KC&K'%, 
@!="1^MH,I^P6R(B)QUVZ6_DR1&O<B-XL=@Y,7_/@F4< 
@#]Q_Q),<;5#T0/&;6QW<1Q"./.T]GD58R0G1TV:?0&0 
@#I%>,-!51 *L9J@*]6#OI B=F=$(\H#8CGJ'/2-^2/T 
@DU39#(\KG<LM;NOU,-BGG]2GB_Z<%FE/ </H@3<'DRL 
@K8\3KP>5,(-D" U9M[>[F21+)4OM!>_#$3)NN$>(?.X 
@>J%F1:TNKBA.8Q\)YM9CO=;RR9T7B@C.NL?I#0@2:7X 
@B46]#:\+-US@\H=T>62W8L#777,!J5+O%G>ECM%=LK, 
@1S,<SS&,6_COX?D&MM$@2D(&,U"QP3Z _\.BT&UN:)  
@3IB7GF@ZD6_I]1J@O("S(YCW:H0*CO94M^:X6UE4EV8 
@L-RO;)G->X6A,?(>SUZ6U]*9>)M?1W#S!QWC WJH24$ 
@.M9/[TG65PE"<X[V"]SQE,]2+>*W6Y."JR51)YC\G@H 
@07PYP4_"7=N6X:5.C;!+?FB\Z!P&B(T(HW$!XX>>J(  
@UU>=6IXU-/-<J:]W]\(VQQDST%MN>GMI]X=WN:E.DO8 
@8H/2\[?AEP*I/&[#QC-C%=K9^(VW,46T/UMF31U#S:\ 
@F?EJ*6LW@3<.W,Y9,:<X>(='V((Q4IZX1*OU3ZY'IMD 
@U_=!P]_9,?[1SR#0\<>11=QSV0ZQQ;J:N"+3OM3K7[8 
@]<@7B7656@=>19X,J,F@/-M/0=HYC278T0R ;Y_=I)8 
@,ACO%H5;'+]GO-B*DS+;M3:1[8X\8&M'))'?5[KX?-@ 
@\K\E;T84^I+SSTW]J?>IX!%579=8<(JQ*+G7YH%113$ 
@0Q]J0P&4>@5DR2N:8'YK#7V2:..ZEEZS7OB:4'P:0$\ 
@3?NR0E=\NMV@L?$SZJU$8DW#)ALRIXE-#T6B?DF_S#( 
@D6$/\+17T&SLJR-?YDT*,^<9;XH@F88<H1O",9<"8IT 
@Z67X*8:@H'FQ3R<0*1ITIAT($=7(X+,W8$PHB1#&WO8 
@6:WINANY\R>W"O6H8H&["+OI<N2A0"RN"F :Z^),OG@ 
@NFH#0-;8K^02]8\TXI0YDIY5?F[<GL<"B77MR?=,/H4 
@9Q*;>\V-?+"95;[#?A_+:ZG41]1Z;ZEK47D%\2'M@I, 
@BZ*PER7B%368>B?_1S1F\)_)/,T2%MDV#C><RQ_5@ZD 
@I$U:A*XH$QVS]NTX/CKH!Y&AI)T+X2<6>LKQ_'OS?10 
@G6A*:%NLYCDM[37@Q>TH=Z%(']TB4(UX2STQ>&^/X", 
@R]ZXI[FQX"E[J%&R2,L_UX1A4C@>;<\OWU!<@:':6%( 
@\H[SZ]?+DMQ7=(]$,:M(N<%H]VT !)E>GNVXZ#>F<4D 
@AJO$_XQ93:33:,*1O27UBP5_\FN3?C%F"&8.Z&L_0N@ 
@V^94LA2,<*+5"4"TU6,%Y\&N8H0S-08+BZ:XNNXK@%H 
@"+1A[:.(1F::+LD!&-7%[UI8L]]LS&.F$GH6"WQ$_'< 
@G=S4E?.!%%S(N2ZM9\TD=S^*&Y>&2E]*].G:^/*5%[X 
@H#RWO:BN%<_I[)Q:N.MZ1162A]SY77V8<[WJ7+RWCZT 
@YE]^GJ0?A2;.,M;4,D).I ;?D"$ED9&=B]Q$/+[XW40 
@X=(O6YB,*]G)?_MAUL:O_?N1FRHX:%F?  %N%YLVGO\ 
@G,5$ R#C:NO:V6SN%ON,PF5E^M9A"NHQ'_XQZ:\M4M$ 
@NH-':&W2S&_LK9R+0#926;+BD<W[.D'J0_=CCDKO )8 
@ZDC(Y*?H_92FM!4[2DI=*7]>E8.PDY0ZR-SA,SYQT^4 
@?G'I)GU[J1.6;-A1*WQ'3,1]A%G;:+S%[A'["Y_R?A0 
@&&;+.Z/1OI;[S*SE4$8":40).^K/>V.%"4 8A\#M6G@ 
@G,E9=YXL@$2D.PMYU[RUF_BR1TT>C.DIY.*3Z%QY<0P 
@J\XCL8^;:8ZAR[%QPEH#"?B(<>NJQ "HW/4&9\;Y>>D 
@,;WN3\4UD).ZL&G>*:KT%L&@]E[AKL<#6"\3,MOLJ54 
@-YO3!>SE-=GA'S,'A!0]Q#A:[?E*ZN_![^);OHR(AET 
@=QHVB"#:% =YL(<5D>JA,<4'0V!< R+;*^2.8P?<WK4 
@>_JB89:[7HB\_?.IG&L'IF;NDGWX8':@L-C#J3 1D5  
@ZZA)8@C,=OD'ICMGCZM3E#Z6AUA=:$<3J8)E _ J[HP 
@[;9L#76?]*K_]WUHOG"B41B63:3ULO--J9J"'-J]=8< 
@ZX;B)K<#C*KK,_[-='X4/\TI"KE.*\XM>.X4\!D3>T$ 
@1\2QBP=,U!#3&PX\][H@4&>P@M$3);Z3#*9JTFR9D2X 
@3>*HJ >,+^52]IG\:G2J$B^B ?:&@1RH?X'UC4@XNL$ 
@9[/*2/P5 O(1[5"N1=:S9ZCG<K]B 1+)(B@4]#!B6F, 
@BY#SN%:CGLMC]?(L3U>_0GKBO\>@BJ"+@@6%+4Z,$5, 
@]R3S(%NU7-0'Y*@<D7']!7P_,-QRB=9E->/1?3P_&?, 
@>5%]-) 6[@E;XTD/D74+*0UA_N<TJ6_/[[$-!/QQ"68 
@(MQK3FW J3PK_":G)% /Z8WBHW>>.))1'M [H(FZHA\ 
@;U6?]\/N'37GL:>9@@9@33,-T-9@*YEJXSUS(*F#^FX 
@ )VNZN737@6N17YJ,&#AD2<4(0$N%HTC-U8]>8'3NXL 
@FT;#(O*TGB!"#L+T2;7$6;;;LLGUN>9OQI<\%N-%XX@ 
@3Q0OE2F;9'M!J:#^(N<#(T<57R+_,0M.FBV0QMK:)XP 
@+7<#"\6ZB,<\+2SOI0&!M9EQ.6[S*1!]5K;,*:<&M9@ 
@Y>4-Z?;36R6Y)A=Z5IDK])==5S\_M?FSR0(5H+<M;(T 
@X@IH1)_1_XQ>_$QC"ZW_)PL"K*@ 1$]'A BN 9+.JU$ 
@%^*$(XJ([6HQ>-.KX:(1K.$J@-IN(_[<Y_<'.](0/Z\ 
@:6]V)6.'!%*^MXO$FP(&5"#-O*Q1_!KYPB#!F,:-)9$ 
@'T,(QKY^5R34_.40/^X"W["M\TP'Y$8$[ A530!<K.< 
@/BV*1+RU7>!(B]2_YL0,6:&W7WC+ NC4(#H=L0EFD,8 
@#P?Z("WLO+HM4BH?9IU5W<;B$G?:WT2,YN$SN,;=++< 
@>)0-)L82!8WCRVYHPG50)G$$Q+**+WZTV\V>K=>H;K8 
@5Y% HE30^M1KA(JT[]787C<B=F)GM[)GQN8E+<^'?S  
@[9W'KWDB,T9 T8R-0B9JWB^DZ7%#GO@8U""M[V8?U!8 
@+M'7<FQ[>C-"+1B$\/CNCQ#V6YO&)+E:]0;)+9-']B8 
@'>6!EU8)3\^??/8S/>P=[2._[Y8D,20(-DZ?HY#RX8@ 
@TOM/./'A#-B:\-1:Z-AF^_]*W$851)Z(8$01C9%;2N\ 
@<=^2G@1^WYQY0DB)[C_U0X<K_S.I.(Y>5_=9#\I+A\@ 
@M'[ 5X%:-^5R^KO>#R(QOT2S.'BJC<4)SXS/\C-5C6@ 
@)0U]/@???R?_E_QK*(6M0UXS-'/3>AFP<8_P6U&6<!\ 
@\QN.PY']6)SJ[-^=/Q#YV*=HKJ&>?;('<B8%_N9;/X, 
@C,$43+_&(Q4.3SRV\Y"BPUHD1Q "FO*-* Z>LL^8;8( 
@^"[]R9D[#OIN/1P]+P_>B+FW)UB7/$,Y(\M'B\1D^^X 
@SYU\)E9\Y@[.YL185$<%RX.["U>=# =+HC EU)D?(&@ 
@(T%AOLU*T@ A\6:O.]6(SXWH2CW_CIZ$SNAL]J51M8X 
@2ZN,)/JX%)BO[>#:'/!GNB74*12$7*4/"=$#^JNF2S, 
@$/T+$J'_9P=QFI-E(RL2]0CLYY(KU9.-6KGU'H@7\]  
@)S 7.L$0H0&U0!Q![.]B[^AW#:"I5(?P+J*/;&O.?N@ 
@BYK7F!KK8V721<8*%".-MJYM>I9R;/9B D+(W7Z@RC0 
@J ]XQG\0E?R&^6N%ODOXGPM[XLV0HTET_:UHTWRD03D 
@OLOR)KW']26FZ1DB6_Z[,F6N+T.R2-8V]K<7X"?<.WX 
@V95 *O=RT6'3YP>!D+ S<1.Z<+N<A7UBOJV/3M>,2B@ 
@ATHW.TPA9]?^*?@[K/K0J-'EQ+Y^A)F0%%(,-="EHV@ 
@']WR'*FMRIBQDK-""; 6*@#4/T(O2^RD=*=>VO.SQ#H 
@7/KA<*9?[7M%6YG+FR+]P@#79LU,/:E$C!3<N<<=7H< 
@YS]$)ARP9T,#XY3Q3*6DW^_ J7!B<D2PI"QTC@FHS0  
@NY_O+(B_O>"<'9,3/HWU>%??(&ER(!_(B=YV8$QM:T\ 
@X$8FPM>N_$BA:C8C]%54G"'8<'=*S<S3M1M& BL*R5< 
@?"DTMTJ)MBWNAZO+2)AQ%0UG\)H'>''U2<R>#((Q:]8 
@FJTX&VO2AXT0SU34I[3FU5XL^2.+^*_C@O("*P&<\!( 
@(ZAC&6WA: Y.'0\OI(@V/!)G1$H:O/K)HW>>=7ZH3J( 
@$^(JOW]G:\8=S.;0%FN18*3H.H*U +$$L35L4(JH+X8 
@Y&"91U^"QZ6N.I:;8]I#9NP9O'R"5+?'.XA%:I1/52@ 
@>:ICRO^-V#W:E1.+8_E,\?3N,,##TK"?L80XH4ZH)T, 
@KNT/=#(Z^5)MA!*[_O%XQ#H0B7+1]$A'U%H$8]E&LMP 
@ <Y$W@^5@X))I(!ER1I]D_?+0P=1]'D*VOY,*$G8^7L 
@,>CDTJ"'GG\=/*O@3\(S[8"X.BK<J1[#Q9_%>9'U=Z, 
@I0Q)!,J O!US$,RXNY3\3M'U(O2,[VP%QB?]SM$<V!, 
@@0)?8II27J9/B0J#$Q::8>PMYSNC*3W*4GLCNN](.&< 
@ ^,H-6ZB#%S8LZUWM,&-WX1?:?2J#:D QS-?%1_N"/< 
@G_*T[%%I?%-8@VTR.%T333S]N+N<EJ]4D[?LQ:2U24@ 
@$A5<Q85@55TG)+ ]"L)0/?W59)8]'V<T1O[04IOU==$ 
@X;8T.3-I0"5X*Y&DT8?-X)[/T/'N.EJJ!6G8!-H6Y&D 
@RB') "422+ENPUC*K9-5L(B\4FIH$2S@W-B'!1C"[S@ 
@-0G,DZ2D25GBPX];^F16'5D7#.LVXO'<26'$Y4ZN4EX 
@X+H+3J8F)S9J&,S-Q!VR ^+3T5Q=4$4)@0J$]<9@.*P 
@$( \9C.=14D%KC+A!C%(ES_JWI1CMI<R^?\<\RJ N;H 
@E-B7PUUVQ*]1C9F96%D54O'A[#Y@,!'DZ6W>_#[;3L  
@A%@3?;:A\H%=AD"6H]F0LU68^^E48RY@V;VWT#$3@IH 
@JVT"+C=0"Q7<&Q*RJJM9E08*XF^-X(I0BJ(\10'85)8 
@W3I<L:[&,KS1\!(=FXK$8!RUQ^*%8\O$*+@IS199??T 
@KL\04@:G>F8Q9@K;M+XRG[]I"IO8^W*_C>L*K'GKA5$ 
@8& ]2W;YR>&FJ'7 !P],![J:\\BT)$P9&IP'C6?)F1< 
@W^\B'L;VS::YZ2"X-(@54+NCWU'50I6FM'[PC,=[%7@ 
@<WV&>V0B8*6ND^*Z: A6,_"99JQ..$%6V]451M-ZXF0 
@RL$^"I'QXJK/J0*5%TU6_9._#TA2Q)^K"^CVC4H6)-H 
@SYL3!(VOOZ+T^W$U1+%:V.H^]JP!?P]96;YN=VSECC  
@>^^ZY4(TX5'@565K X!]P/:R=BVO+"39HG)10@O^ @P 
@S<K>N8."8R"G%JJN_WW_O'IDO9L)+0WG?3[ATB' %8P 
@@_;3!1Y@.PM)5FA5S7**EXC$S.\^?@EYP^IIE_$+$JL 
@IZH#NUP\1BB]QK7KGQ(K;[]]WV%FP1>W/H**'3+<D:$ 
@G/:2;];4O$4<FP5[N$7Z>!.-\ /;V(GV/+ @GPFI_@< 
@?YULZ<ED^[.FX3Y3L@+3Z<:T'K+B^HF42B5/98F%IDP 
@'8VD@KFN$/*+Z[D3K>.7:1$]@3OK3(LM *RN!BM85B@ 
@=N/"XL\<[7KF$>T@CP/$4#<DFX1>07X.Q*=,Q[_G^7( 
@=2CUP[4F\.1%Y-L-OX=T\YR>J2K,9*IO4+.X,&RZ^LX 
@F:"1KYJE?+SV;1=2V-H=9NWZ'1LUP__*PJC5&#'1$#0 
@6N8)V!;CB/ <:6 U+(3%F)URCS*M;1&;=50^2'O09PD 
@; K T*@=V&R!R&T^8QU3VC49@*] W<IC0Q821.Y5)+P 
@VS>WULXD7/<$)T_C ?(7=XR;4TF .N]XT8SAJPK&(FX 
@6@Y+&O#.6XW[,@U=+2Y#%)QJ#^,#RL'XKV6U/U(C?FT 
@%6W%[Q,$A,3&UK8:*G%*:?''[D=*^#J]_Y&65DC.']( 
@"*K:)L-+K7Y-B\@)C4G579FMDE4KJD]K.OSB[TT-#7  
@O6X*TF\G1F96>VY'DEOE=?=MKZ77;Y#<;>^3WG0JE8D 
@)\'9%W3\B 3\@%9(#B4@C*%<I'H*5-NL[\/,C9%50<T 
@M_@4>9=&>H)5++\Z?TQ:<Q/J$JR 1[4E!>TAS,9]Z6X 
@HAKL9#X];_CZLXW#J[1*,DP*.\*H5M#U+Z>=+ISJ7I( 
@H3I(26A7(!71C\>97"$I F$4BXB "AXI"&++U$F&I[, 
@3B2A*#,1^/WT8MR!C:@T^89$,A!&0$*TZ?_"B'0!BVL 
@?<;]. I^-KEXOE]ZE^E"J81HBUID'?,=H^0POZ$!]S< 
@/A?Y*VB7IS\HG4IJ[\D2T)$-@LKA8KY*R\*8&R\M"@H 
@_9@Q;O]O3+7S,<1EK27U+]0K'1H)G VHT-9G-&)4P*H 
@0D1_HR>#LW)CY@-?S4;!_P=D/KHW57GB$5_E5S[F)$0 
@=*_CXT8((_6 ]' 3* V(O$<H$ '8E?4]V<X8SH%_S\T 
@R5T9W%V--V)F0F=&QD]_"KO;/7;&B?0%FEM.ITR6Z5X 
@H!<4I-QSB6;(B'*<3BI7^OP*@L!Z0W5,*O 9[A%9S3( 
@ZQ%Z3I?E\-%A-PR0=JAK^IBVH!IJ) X?[J5;/]/%,[T 
@[;*UOL(^/+V%_F)8W3UGT[^^'IMV 0WJL6,?+E7[6)4 
@/4S3XO-B 7*8364ELA?/>W<:"G@OM"Z&LP7/8$C58E8 
@<9B5V-=6,)J#/\[^6(28%4#/=PVMP3D=)?,@V6^Z290 
@$7'0A>PL[T@E]BD>E+HN[YZT]PKVHQ4%@*%GOZQE*'< 
@KFR#1L[>!CF.=3C,RL.K1'?=7S1L#GRG(BF' [RZLTX 
@_.B4^ /9V?7^'-NC=V)/C04/.ZNMY]G-Y:O>O\E.5V< 
@A="+%^)@9\R7*<R+M?5G)/:V44R#]U;#40TE)RG]8XD 
@)?5\RPJ12Y4M<XNMJG#A=R=MC:!;K4[CP.TZQTY&JV4 
@^.CG!+?/\/I5E[?X,T.HI2Z;%;<C=LO)!Z16ZD46X!D 
@#[Z/]>H:/GI:-/\:I<+7)BN ]*[_E(Q,RTM+/ZJQ4<P 
@I#+>:(8F;.K0?82&;0 PLE0U5S,-0>J%EPE!%O$NJF, 
@(66$7K*C(KK\U1.?R+RZ1&TIVV/0+K&DU,$VM_+P&-H 
@4-@VJL*C'88WFRVJ&JZZ-HF<!TLE99-Q_A6>TPH!T04 
@K\666<RL#PFS7% -#_O!Q"VE.EE <!-21*"/^=A=-5$ 
@YBO0RG1 4.&I6!FG;SQ6?P724@]>#\U=4Q2-[<S&I+\ 
@X#A:\*SO@RO7#."_)0>8P$?'U!ARWYIDR@>73D$"VQP 
@6;_)\V]7JV[UJ.K @7D82>[=P $+25-EZO'%^+* SG4 
@ZCVE,[B706FYX3*-(=H.B$ ^M?JJ+UM3$YU/U4TB;&  
@'<9P7UCL"%MIA@AON=9N'(Z'7M"=S0I4Y=YD9F*MGC\ 
@/\&4I -]WY, -H#J1*<8["OR-0-&["7?=HN>P&%O/SH 
@7S-&4&.MHCDI"04^9#IL=;P)$Y(5&]UWD^(UR@.5*D< 
@$&<+S=Q.U),C5R6H7<P4J%9N'I_%,LQ!HDGCA$\Y3#X 
@7[%^4RLAZ-\O6*BZO-<9BI2O7HA 'M?1'I'@XH 7# X 
@.\ET?G[WG9"M0"VO%3&;/UHSZY+L#WB\9ZD-1QAVB)4 
@+UIU-O.1\X9/Y\=[LO.Z#O+RR\6<9X7MDVH/B;!((=8 
@-CILDV:WR)C=/PVGX;AO'Y(&",^I^LM!)=PH_*P$SKL 
@P]7/W%'RN;&CZ.XC3MCGUS1+'^??X>TV,>OL.E0($0L 
@\3.K\H=U]]?1X]:U-F9C5SZ)ES*W"0-!^,O)C50_^Q  
@ZA)($[V]2ZRE3)Y_(>>PF6]_LI:1IO"[C(!=:%7(_:H 
@N%,+?]/ ?]HJK8^&'\8Q3::MUE<EW Z94FUAG.UU^4$ 
@3,J@\:#6S%*+7E0L5<H.Y5ZG5ADIJ!Q^KAO5CF*>'K$ 
@:N#$IU)M,-D??>[JO[M4/&1L,>VQPXK6**7JJ0=MY0$ 
@C3*\O9=^I>1TQ>\TSEVHO)S$89*6>1&IO%UJM@_+_:@ 
@_274)Q/4+ GL&J2D#T<M^84&N-?52BXYKEP.70!=DMP 
@STFKX.*@ (W^)]MK]NHUN:S @SG0%_$N'=Y1D<O20&< 
@ 9FF(62XJ&A".3<;9_U4M;AW2>'_!23&8O74[@?\9UT 
@+,8]L8E_D]W,8_/#M ALR,$-)>5UE$].>Q6&7M]&6>  
@>^!Z\KC:OJ\5E:0:*"D:SJT_"Q:SC%P$.=-(AQX.EC8 
@V)5>??(34TF2!8^=(]NB=!.2EZ9@[840OL>7@_.'^>0 
@L)\B*<EQ9)G94M'6>PJ(DC(PL9Z/_FI]BLXO:06>PP, 
@39JD21<_>Y9%U4LS\A\]<ZWP:MY2$W#.[!X&@?"$8QP 
@%@YW!)F0Y< \"Y5,Z'N0_I'NN,DG V?M,W6Y!%36T"( 
@>:-7ZA]'QS<F'H4/#A?7 H9'P*/=-]8Z'6[-8]_4DF< 
@)ZFH$@^EH6Q<UF*2?Y$0?AK?;7T)B&A,1R=C^<J+!)$ 
@L+EO*1G;>.Q\T(S-GM\;NM3NU<E/9[H- R,^#%?[5$< 
@C@ %X$B6?2R2><+?J]56.9G-Q]"%7W([PC'Y""0H3Z< 
@PT)ZG!+7]6VB.FF7U)(ZN5- \>+:BV:E<']ER5M_3W\ 
@XF\B#&/(DY"@C^_J@=&<^V)"-]=0ET+IY0TMTV0KX:4 
@N'BS'!H:<F.H^K-9E>0+*%#">4#$ECSUNCE,I?$T!3L 
@WHX=6?T)[CD2>Z76%.3=+>*?'1P BJ2*!;?9;)Q_[OL 
@78\Z'@@^38LBDE:P"6*PIF>/$Q?U"IJY<9'.S_$_&\L 
@^/'LLZ\NN1/*X#-+'%&"C!L]=J)WGV"!<WN_EK0> 0, 
@GT.7@-F&1H'LHTL^]KQTO.RK(.I32(V7P=8T#=OY.)4 
@E-I0+ *!EOPYD%11_+88ER3"%I,]I+SV#6,WC7C9#B\ 
@A]AM.X] N+\-HIV)G<_\*1_WO>D&RFN\6 >394CM9A$ 
@ 893\TDJ:&*BL8O_(I)G#\19ARV@)PV 39T5&%%"WAH 
@$5-8=V)22$^.5N;FOR0)8/#J/HK ,)N0YM)*R!=+#HD 
@@9S6I(G8;HHA=J6TY[D=)3] O(B)9<WM4-<<D1E:.,  
@OP 6[ 8\W7^$8AZ1 19-BY1^B$5(:,:GO?I&4YL3YV0 
@#IN(HN3AC2P\P?$R02$+Y_9<Y/!I^MW@/\?R36H.)J8 
@-_JR2_I.6IS(/=6\\M1K6'>FOPQ5VK^<S#Z0C]G,,WL 
@ .>SKY]K8'*DQ5>OVV*W+#\XG\F4J98V'.>K!,QI'<X 
@=T^7>QUY?#1P.U?@PS2>)BG-*$/*T'B^HC.&"P8*IQP 
@JS<-R;?FDPI]3>WRP;93D@&N5)&9;,>++N% R_.V%VX 
@7V,KAYJ(#']WZJ8'@LU@7=1;19J%0O7Z9CFLS1)@]V, 
@DGPXWQVJY[IUT)6<VA&C#UGH%ADJITV3< .G]>UEL\T 
@5NS4=UP);DOA7/MHPS%XT-D5.=A8:1?Q> I4@(B"\@, 
@\+#,>@P>J3@$IF- %_NSHDC!B3G)(-%G [:/2?C3(,T 
@RT9"+@IHP[;>H$P(3)VGA^FO2O4\"G5M9W ].<TK@[  
@UPC_,+*QC-7;<0(0_%SCZ%,V-P\0TBW^K):)]'*$5?4 
@[(4/8J%Q#7#"7#KA_T=\ 6JHJC'VCK:;I5/D"Q-/*>T 
@^U*;2OQ!O&[8U0??*8,$.#'&2>&"IYY+WS>5->>5^*, 
@9Y_[96!A+*"*"@@L(U* RT*!+,2XB^(K%VY6@O?%K$$ 
@^'Z,GHVSN)WG@D[_(':T)"U90N]=#[!L-I_9 D<-NEH 
@\DP4CW]%*]H"JYQ?$T0TT&7>DO3[=<+(!"IZ(@!XM%H 
@@&T;P6I*W;DU=ZF*&&=:^"KVY@>SWDP7?BG9XO,AB2, 
@'EG>#-8X,C)3ZMD;BQP8">OP4Z7<)\6C_;D W\3[F6( 
@!S;M52@KXGH69B+.TL],*\-S^=O=WL)B?@<UC?M&%>, 
@FQ(*L5J GE/J]::Q6[$Z$G"Q.ZH368X>?T@+>3 >H,0 
@?H*,4/=:,H M-K0R_A"4X G;QM/+V9OE!0 THKSDNW< 
@W=:#Z%*6F??++"FQFW4:Q=IO?<OZW)TB;3W9U)3 \\@ 
@4SRM!"0!:RY:#$F]UQS$@*G8RW:-MD0FY1^<P-;>[)X 
@[NM6I$NU?]42(-'JN=-H<S04\<$3X]II#D[?P23C<G$ 
@*XY33F8Y!IC/CP-A)$L)%F:B5;K!KFB$J;J6J=P(Z), 
@6+/#6FNCQ\L+*6%.RML$_;,$:]]1"N<[.2B8NBZ1H(P 
@*,]_-NX(-ZJS'J>S0<P#$8\!)6[&_2U#./0%#\ K%ZP 
@D)%$YD V38N2\W/;'%.M@S*50TZ+]$8$080:UN<(<7$ 
@"I!U>!X_)GE9J 4=08H*/E['/R"$YZ:D"T!=B7=I1E4 
@/X9MQG3^.[CN4MQ//=RS0WI,@OY\/BMCPZBWX&O9V]@ 
@%:]7Q99[[)*3>H6LO<2S?P519?!ZT"(W9Y#U!BCSQ$8 
@GZH>&<$&K(J$^'FN\"SY8PAV)"NF^\)EC(;_.3?X8_( 
@5*BR0T2)F"]:H0_XN5E)['6MH)_Q!!')P <VPELBI(D 
@>@;CYY NQ^BBQ%DI._0C>%^ (^P"UVTU&F@FYP^Q25@ 
@O1DS_Z9L4$/@84!(IB5J#PXJ#XCUQ!DZ$%-2'*CFU<P 
@>([=#9M?Y:GB[-RKI%31\<5'1>]ZIL1W9*?/ ME29BH 
@!3X59DR)]>8;*.$19XW(2IUWJOU33%1B)?DS:7C0T3T 
@""OS$U:'+J;V,_'>/JX8-!TD3W-FM@<7B6"V.#/7.FT 
@(5"ZCO9@2<:#<&TJRGC'; [,[=IE3($_CJFE2/\(&>( 
@%1+C\D/'!L_'D=V/&&N]D'W'<10VC%J8^7?$BT=8=:, 
@D_D$#(>.>%8.J'0-F9.OAK360I'DCQ]HM=2O]CPU3C, 
@:@;4@@)FH*)6C*K%&O VL'!;3& 7=^FOETV"8&H7-TP 
@6).$6S;XVM0-_L;O\)O8,3K9?K^E"E36W[0K:H11G_@ 
@#1$)9R8AA2HG8X,4J!^M0OEZ8%_,.L?EJU[:T*+J#]P 
@UHD4K*IEI62 8H]S'J$>HTC9 :;K^D=#K/TJD34*]Y8 
@'K08MW1-.5-)+^CX.%BJRB3_%[ HFOP8M&2=VS4:[_4 
@#WQJ^B6:,(@SMKIN)O(#T>CIDHC<RC1S\F[T6S=_.-, 
@PMEAQ@S$E@44*ULN&>W,!FD5]D'GL\@OMGF:]#Q?)Z$ 
@9@)'  <<($+H"1TND9^QU[[!<@;<TW8U]'?"PEX.9%  
@;"UQ8H+EJH)I?UP#YTR8.9:O83"6FH!9)'LH=Q).;JD 
@UPCV_,%R1&O0S$&*W$'&)G*Q%V/""4-4T]OR>BL.4.\ 
@XF%6OFJC"=<7052UUY\\1$*'+.2 :5%^PKB#E9.5J.P 
@M0M;=PRM5+C=1Q>?G60X89]3ID8V+:XIOFSB)U;0/$, 
@,>E/U6\P=A'LD@=MIZG"=_B*B^3>0V0H/-A)W_M/LG@ 
@P(5[7"M0R">KM<WIO1:<.4?L@_44*R^2>-V"=&Q*?0H 
@G$MC,'#/)C58\Q.:.9V\$L>WD0 F<I\$W!;@4?]^2V\ 
@;TVO,^/:<^8"NL7?N/$SKB&.#HKVB/'VM6F/OR%RE5D 
@[ELP]\J&O+1SB G2,T90RH63I%441%RL"*_2 [MB0JX 
@ SR3?A6_X%LSM=QQL>ZXF80T:'^?SH(G-/"*&WD/(7X 
@>/;7\D#@0Y8&%;1TS?BA<9]XRMXS'7G<R>>!9O."NZP 
@'[UXY3A^"KGLX8VYF;X$[-D4:X#SP:9Q.W68G5]=";( 
@<I$\P9 ^CC#:3/#CS>TG$!JFRNYGYU$J!8<WGCQY/7< 
@;US#8"% 3^!2W-83_(8+TXXA#C%K6?E5 >:_%KYYAKH 
@%25!YR0UAJ=3O)R0:,S]^W DWJ(!?R0I4>3R#1Z \RL 
@$'0U#*8YIM,@4A3B$AP&?X'W\WC%'^,(;Y'A<M5H-U$ 
@F;1#4!>;4ALTD"*F:>FC)<D7UN"]I8M]Q0U*'VYIZ<< 
@C+PT#4A^@SH@R1F_%W(VN+@,TGQY)^7XN\6,1RLDB[8 
@!AXKDPZ7):7J'*)BOV03645(%GW>H?H&>>@2>S%9F\\ 
@+ZS!"_D1>EM1,"&/F:QED%K*K.?H6^]X7A-\_CTZ1QP 
@SNZ3!C<DEZ#.]%8X^MY*HYS  /-'COG\Z5R)/P%(XQ, 
@_2RE@R-D8WW&-MH[)>"/#2W_J R5C_%EN!IX8YW!7]8 
@8EMTH#EO%@QYYKE_BY7OPJ46;*8 C([KPJ Z:D-6D:T 
@6,W-3-SLRLI!7!0](QNL3T&:0%92$R^_@?@5T2$J<-, 
@NG<6!N7BE0%I&QL[<;.9@BN5$E&#]@D7 8%K[0_L?-( 
@B0DMAX+/789L(:Q\5(N!IX&=!21QXCB$OX-P]V0[6_( 
@XO8E!.D2,DI )Z .4 8@YZ@JW-S;'JJQ99C%)(M4,ZH 
@S:+': R<\6;)V3V&CZU#W""<N5& 7]+Z0K .0MR_87X 
@)A0^F"1_^=>C9B[7@?SC'MO G?IZ&D0J58!5"@O! 5L 
@N?)-A1:/*?18'.J=P7A.@IOI$9%T2RJE>UB9I746SBD 
@6"=2>%;"K7F#DMLT-(.N?D41Y?7YGVO62QY*N(RI;J4 
@ W+;UBZPFKW&$;"K"LE;0JDBGB/N_B89N]/S&KY_1?< 
@IY-M4""Y]L<CW8U>+5237Y@0=K,7,)G<!#<3+]B=GX8 
@<_0X&'-T98C]]>+;]4T3ERF\GJ^Y6905I&2BMT("M'P 
@O-XKK0K<!TH#LKUYY6[C3?C?(\LNZ5$-KQL?RUF^@\0 
@FTMFG:"OE71?EX,2GL_E,/L^38ONF6EK,D]OC"(6>PP 
@9D0?K,4NXO/_7H]'OJE;#98-RWTLO+A3VU<@>J@.1)T 
@13HSTY/&=6HG [1AXFD(;*(&+NEOH?R!BQKJTYJ61"L 
@YUU\--7YCVP/<(%8<S^!)C8T!R:(AAI+J%+9!/28J<4 
@[+=H"V0W:4X_#;4;TSPLD?/C:<"@!S%=<_!B*G_V0[D 
@=S2IP0[[:[0DA>!.SE WRF&IJ)0*LM"40 J).2"8?2X 
@\:XLIK)U-KQV;4F2:\_F*;(%.#7#(^U+PCG?N@CI72T 
@E[(QUP(J4N^V)H[TT'JA!CXJ:6 O1[T0(I&$/LIR$ \ 
@C1[E5N.4YAOP7K#78XZ;Z"DK5X!0<5N;\SG>JJG!,W$ 
@C2S101;18I5)]>[$=1>NE6[\'?89;*\U_?LE85$;'1L 
@GJS^GE[A1@:)Z?AM_T\DA8,AQ$ +,L]C-M.H.WI6:R$ 
@SVP.@><6%Y:6.9VK&O1VF?2,EF1/[XBR2UCDL%VAYO  
@\U-AP'64UA:?9X'U IA(GN_ #OVX?]@+.<RXY=T^P]P 
@SW-CD5+$'TZGB53OJ9>+-XRM117#4Q23NX%9@_+VR:X 
@[_Q^97:BI3RVULD(RY#$#XEX*F)_P,I!OL6=.L;6(Z( 
@"!"A2/.K]:?Y5$#[;TC>>9,19K2R@A><,OWTXB%+:M\ 
@26"_!@(MX2_ZVT0:)SVD^Z/^R&U.</%6<VK.V_T5CWP 
@2WHLGK0FC585P8955R,48E+O-817&D9Y)\.3%-LSHT< 
@::2/?3;J6&ZIT9:+SI5 RY;L\JO\E:%^G8N-C ,D[O, 
@?XH 'WHNSDGY;P,GNYQH8'!&U>HRL!^1'<BJGTAW9T4 
@GX3/$I7Q<F*Q01NH,Z>;V>/F:3CK+07/KF+4GI?0+G0 
@XB>S*%<+0NO_]$#JLH&\)X6F#U7_85%\$>[S""CTPJH 
@\8TPLY'"19>/9TUC$Z3+S>24D"/6OZ<8GZYN7+9K'.< 
@4<'P\F^+CB:DPJKMO,9QSM>%2ZWJ%J[@[$$P2A">T=P 
@U1BI%Z,;X3U8T_A7UM36J-7T:;39\ %[@7%X^HLHU]( 
@%0$M5QSV%L/H*:V6UP?(/2#5X"Y.'1;E\[\$"8E87X  
@4AW_&![!B\O2=TU3T/!'&\+)/])*->#9UW84 >I7Q7, 
@RZFC/#.!7AE$2_SBZ3J#Q7$6DS;\-WFTXE_;_OLA!6\ 
@G3<EES=OYY*F897 :ZZ'0IGH(,AUPQB*@.R'%34XW)H 
@7IH0"\76@7++ Q.*TTBE&>4VDES/&4* '?"C!,;R3_\ 
@*[R801;J+%Y#AUNFT3RLXV:<>IWE@=?S,S>K7P.CZ<4 
@B<JY%+*%F>]J4TY %>*>\ X:=WE']>7+_UJV3)_+)0  
@.<V:UE'@AI$U4ZPWTGN"N0[I0W]0@,[+.AIX^ *78 @ 
@2Z-5'[72<5F4RG<E H*EI8(!DH@J._$-C6NUH?7,ZT0 
@"ZPD"3?L]&T35F0K=G89OOVALA?T?P% >79#$'Q*)8L 
@^7OO\;J_&P)"DI6-9@8'@F2$?9H5237HVNO3FP_7Q$@ 
@HL 5-RU^<6VSC[8K$@I"@8+0M"GO=K)HNXXR_X'0T20 
@]W!0;R_8 TM\V)/G:0+V [G K^DE?3%WSK3*YW#GV/, 
@2_@X 'L#8C\@,K[^D1M6\+0 _!1$51(4+&>7*I(%8;$ 
@G/N%F<M=UWJI21EC<,*&VGCQQ..WBJWX0L58J^"#%;\ 
@\*C4KV/OP84&1)61:$,N>Z^9&"ZWN8UO(A=K_2#558L 
@IA'QK+(>:D7\UI/)4H$F;.*CXI<VL9)]/DZ487D#3=, 
@FI@\4#QU#>CEJS4=G/:!Z='2_"/Z0Z*(DJ[O\A#XRGD 
@]V:T[1.A?G],P/N>.#+5FY7]W#B[P$5I0L1'844GEH$ 
@U#!>0>L6'5]6L'-0=M69=+^V<YJ?]2]#<>W41Z;A2<P 
@OL840PX#B.N;%V# BL$-$4_D"JEVFQ$HNU4T#9>!P^L 
@]I>O%R0D5-%M^&15;LBD'Z&A9QE=L_" $I\YE7M)2/< 
@?0_<8^]A!=*N%1'KR?F\0,"I#1I%R1*G)<QIWA+)E0P 
@+&TY\+K^CYV<==,SF#]:'^VJV-,#=&JDW'?>&DDWHLL 
@'DE8-?FXPK$F2FNJ<;[M4>Y!@U ''R]3^-+Z*]9[X_  
@X_;<0R*2N]0DM<9)$Y>[#>YZ,(8*&I;%'DI?O$T/,&  
@JM$P,3/T3S(+!B?V/#KX@-$%$6GS*"XX/_G!SXC]X($ 
@',C)O+YT150>8HV076R'G/F[MQZ?7RAB<TF.7+7I;0H 
@L]9>P-I?/EN<.*=&N8-NAT"RM0UOJ1&&VG&@<]"K%!8 
@ZL?4LZB+*EM]J@:3X;!=!F]BP/HJUM>"%CG# KJ77 8 
@A#'E@U6X,>%-M%FVN@H5/Z\,T^:^>R,VP)PHA5S04*L 
@BH=(W.\^[A7?'2"=TCX 6)CL!QKZ=G9*J=>'H[7$2T< 
@802*'(M/"9,G9XD;$<#/%9)IYY22JRL9HN&S?3LQRH4 
@*((U@Z##"X'::&K#P>T_-_E^K]LCVJ8+IU=#1I]2+MP 
@/0# "$':A 2'A55LV,YXK2::@.6QNB9\>8\5;N0^5!, 
@:\RY(CTXR/J+2C7J3W G9H:Q$SM,CXF,QUMR<\D 16X 
@"SXL  8#C I+=7A-NS5],DL-;SU\F=$2$O&_/++4HP\ 
@*" #^=A7)47CCA>G68.^"D\C5@]U/(T Y?PZ-M,PD?( 
@M=U@#A++/J9+^(:EFC-*#FC5Z/+O9:9;0%)_-CU&&Q0 
@RER=HC4U7>RFRL,%UZ [8,LQF=@:51M]-$#YCPR'+_< 
@;[DJF>ZJ3A@Q&#:6WY.30T.:W%@OG_N3&O=8MQAFDC< 
@I]=>;0:EI36P2)-#[C@S= EX[U7[VOY+A3RZTO<>'=< 
@NK#@8A_@.BFGR#=$H].ZP.N1GDWJL;K P/SO+_O*5XH 
0?$98D)L=R.;1NY%@7ZA5*@  
`pragma protect end_protected
