// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DdKLAAZOlaN6zsihWgdSsNPcziL2d00tWStTk5TBMraOIHFd0KUP/nMxmSkJq/M/
oXLrd+i5kGBj+/qPITlv1WKhqvjWyU1GBvK0x0japMOY89Kzl59uUfF/dBUmEIsI
cWHZZ2uEt1vVskUfXLTOmtEpIXkJEZwDJJFJ+2rhpeI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10192)
sroUbAxZF0aK+UMFUiLxMyyH7gIW9Z+EwqzBGCSi5sBiI9HcXeYd/dbVyX86eTB2
++SE7t21Q/9sDnRIZpuKrDmiR8X+XxkEvbfrOgaK9pWWgIsqChmEPuLKPpWq7KI/
Y5cjR/1Hpwrbxs3Haciq7SYJeTI6q93K+zxuXh/CZ1d4dJAZE4jZYICbn7Vmx0je
lJmovuFBLPErvTlt2okT2b6DcJcKY4qZg1j1MK7vQcJ4l4cMgACQYvoysU3UI2+B
S/oc9bGpLLB7d06Xu187WbAj8R6Bq80X2OqFmJMCj1ymaCBMFYyNfiseo6aoRg1z
CLkxKI2saAueMGsZIjA6GjM1Yxe0gm7xTW1L25ZIInHNMnoDYgPNz64TDLRMN6XC
P0GkMARjN8PqbrqHrMKsNpig8klsNlM0diWEEY5NmfhinDJV0O8hVjf+b0rpFY3G
8hhwVtIB5BchBXtnlBWCsORsZ2mUKSDudKrNlUZmUdck3Z8bvYY/QAGikwrPlNS9
wAA7VnJzs4Bi0KR+UCEnLGEjPssIKkOkft61sc2Rwsa+0olFDk//wwrVwYc+NZhY
y6wdOyvqlV54N4DvsgBtX/VnJyG8idXlnZvlemWkWvyYato1ApAcwUPvVJS2y83J
Y4Coo9P4XguPvwlHt705eBMoxRZJUv505Lrv9DqIphVPzvR5W8jGhTi5B62OgkwP
6Vx4hYnmGLWiZ8qUj4M39QiBjujqREIzxTKXxSvnqhyWL/XAkPHzqmfLk7Eu0cDp
HfB7EDd4reXqP6DbUo5/WNJCaN8QBJ1UeB+F4G0E4jhjB8yaw4UMTkF3Oi/pYtNl
MR5jb6Bp6Ta/BNW7p9fVkS793SP2uLsR1fk2b3SS8ZoGjF3RAE+56QAsm4pXTlQT
4nKmC6P8fxNXQXRs2auaP5E08P44dvOC89FnZmHuq7sw/gUKmE6tpmvOkzHN8lu4
lBUHfE623J4Ousn5k1qW+ku55KuZWYvgI+Tk/+dSOCunphtGM4gR2M1JwkLVlOD2
ZBVUQC3U7KUG72qASI2h/oAm0s8u7yW4Nl7lhBZeSBXbTdQSxvD8b9GCtEIZ8nDS
bD9h0VGfkaH49dVMAIaA6GIIIvHiRZt7ifDKwXgmwkFdzH3mBZ+lypH4+blyFXcN
4p4BF5y8KZonp6ZOfQBDiaZR1hJ+UWCgbiO2J+xywwlwpe5lTcp7s33D5wukh0b+
jsOJBV4s/aN0Uu4ynS4Gmxb3jixHn1lwtfLtFZP2Hq3Cj/1co7JSW+9oux05lUg+
JzD7P4wDrMSK1xAyM7J5+YCOJZuQhm/SoFcFHRxUKGIQ0JfuMWqOzxJP50MLlmwI
LeYdA1tEkcQV50DpxTkLWpmDKnW6TQtQsVAdGj/ZniccTbEfiBLHYAJHhRHJYHKU
nXmO3eCyPb4emEtBEQbfRKmqpFg9fK1civAQXh6tT77CYeGFaWp2CdLliqfySAey
PitjnsR93XBoUI8vFHrrRqyvoUruIr9VVu9or4SNnMwxgnyq3km5MnN96aqQKhT7
2yuID/o4jPlr1YmaAmfnf0UppthI7viDjTKk+YapusiQf8AG517myQrxcpMFxz1N
Wg/FmScD1hqGwK29V56vkrOwNF1FpJJnBNs/XjDqvdo7y/QxUvjlNHU5NfM5qiOI
H4MP/XbQNjpL1F0zwb2ViXJc5VGDRy4l5MMZJxcBOQt4xWCzi2w1g8WdyEv//g96
tlL42Hqc3Sp+mqVr4/pNs90Onhni6gO4WF0AtXVqZnLjqP8Tu6ACSIQxeBySPQ9E
9lFh2+g/bvI3/fiXmJw0ujBs7r5bIa1BrND1B5NmFnRsjjECL+xtUUJyS2vz1+xF
q0UnNufbj4+jqOW9ElcOcx1z/iKN91/gPBeYLGennhdBpQylsFEXekdMLmLA9EgW
Hj5vkTG8zXxj2aZuekHDhoMdtAKfB7HIS2eupXJMpolDU0Cvfx8fL3dY+N7wfQR6
4mQdrH++iQNMi3ymy4IdH804jwuR38qUjEk145rUT2GcMv72ehY0jZ1P4r3lpITb
EjFIpw6OfgXz67hUnIPatxKUywkzRD5Fc2kkx/tHjVPeQUT75fbsEP1kGGj+wQtK
np1pqqsnb2Bqn03YS7ROyGwWRz9ffg5QMeLWJNOUx/zj1sWjkIMKv8UJSm7ctVXe
FLZQlewOXbwzhxJ1sLauyTt3LTrbXEEXGG1acSdPw1g8UiILnG1Fb8n5dC4VrsLF
62BMgzZGYQeyfll2LBCEg6QaP93LcHuAR9LPB8bp9M1eOuaMxa7kUmbtrHab2BN9
is/XPeMPX43MYlORZfNJFXunWoxh3GpveuzY+ZMjP4CVdWK1MTXB7RKvDG3hfD2F
aW3jofTK9an+XSFiMqMEl35GM3JMLQGMQ6/oI4SCkd2OJqa8w1EQRFmz0cR3lkUt
EED5zDhS0AY6Z6rh2k50Fhb/uxAW/uh6I08BMDG4eKb+fMdd+283a2RORUGpgVG5
2GA0BUQ1Uyz9Xsspa/tLFh0ySFG8mz+rqG6QT2OBJ8lPVdbyMXb4khmR2ZxuiVXN
IXmlqZiUaDYAwZmzyqH80OX6jRVfTJBurDj6VCZsjMz808wuFX7mCLuVCcHqSGqI
OyRookYHslWrT0lSEOJ64+UrCzHQuhHULCkTugv0YJzTRnNsxmPSAsC3CB0qlwoB
+9x5+sE219S86Yg6bk8O87A4tqkwtil4aUhwi511IWZ0xvGWhlZiSKIc6LML2Bkd
Yp+mSwVj0sBRAxaNbDtK1pMo9jmYYbBaWRU+PcUPfMH+73MTzj5gVqBk5oAEcLxh
m002oRheWn+OJ+ne5+APkUrAMl+TaWPL+l7LjnfN7J3I5faYyjJa2BmSU5j2KThh
fUByiaC9CyDKoBa4v5P/CopZJjM89ejmndQkEl2i71OTfoDD4VxqbvhuBdJ+gxAx
gv2gZDgUPY6JwziIcUjaHGp7cm4GyLb6ld4zsUkTV3Pt7jIxXHwu4cSfcjQeJL3f
ySypQjL2RW8yM8/t6qVEBMnuOfjMia4RE+VLXgQthyQhkZz7XG6wDjpH7nvITpdK
s17MgeQsfTq0TyjQAyOfqpyPTCiZ+XwiE8IfBz3z1O1H67rqRA6iyMuSEGXiMsbn
5k9HvlILngrw7mvuvhPZIuS+ClvzRTgxeT8ne47Sabw6ezEAr+R1U8wQoQUzH3RN
NuMQg7GxOYQUmwLvfrwBH3bxxl4dZXlPc4udOM9Reo4QCj6HueYKvANx8LepFAzp
LM4GjxMpmr6GWEBMDZB+ECe2Otp5On2HeapCBFSdvkVnuDRFszoRsEza5c7/Kx3F
o/jNXxpQN6u6RB7rAyvHD2g1SQAAZ1JQcnPk9rc7Nk5waRiBRIw1i5U1T+zL+Hsl
gzxgxjXGOhuS8feJbhd9uBVI3kUyZgXkvHXJb1lh9kEKL0Fm+OQ2a+EZIILZdjh5
vNgSJ6P7NAsFPKyRcFW1humFixier1gYe5BKa9g1b1kUm6CjUiz5nNx0BtAypJX1
P5Er32psU4GzZFvuh3moTv/2Z+gXF54iINcIXXd5KXlZpRkqZuqs9dyFZ72byQVI
a9GlPw6jLmZzhOIoCrdmYf3w1/r++C6QZthz+eTL4Fd3TOpiUOif4hOefKaKDn9v
Ndsu/U4mCBxFLBacT5W0jXVfJIFncytsK+Sv8ehpWi0kLjFRShN2lo6hIc/9X+K3
LG/7nGAd/duemjdSD5e+YoVpEpjCOkHcqVrC+yOw7wBb+LeqDPrSeXEyWhWcenP8
qiBuxRtd9nvzMVyIHknR4wiBPxbOVIFzSFSvfPII/laWOe6IcRg4ZA/8YwoiU+nP
0jLxhZEBkJHoWgsktt9Loc57mJ0TMk7fNWdhkWq5Wq4ey+yUwEqgT7BmsZ5j105P
2m8nTauyQ4zAyr2OsPirrUWQlAbVCkvCK0itQzQbdZVabDaAFa3TByuiDbIhIk3J
jZYCCrsJvvEI20RjAvrA5+gUufJAScTP6Aa0/hu2VLUmN4vTsnAXSLKgfHOxFh0h
WmFOhSRk3Xhkj0nBTyEVes2UUHfXdKgO1KdV/9p/P8ioQ7BWxqe2sbjSgZg4EtCb
AVbWPhmOv2RnTQ/tjPm6Ox5ykrBUAk8Cs/VRMk9k7tXadg1TiEWsOpwYbg0T9bi1
CwaOfWKq17HT/PpnOP2d2eijHSTTmVHHvsYn9w8P8VWdYqXbsvZdX1NMVkrlcaZg
WGzOVpBrG4lXm9BiR7My4Umw5DaIk4A21qC8AKkiEJj+WiejJ0v9gxY3lR7FYgOd
pv2q+4PpXglGf1niGJb7qzmXKFyHS+vHIGaRS6KEthTLm+VW8a+mE/d7+QKxN1Z4
tt2pI7X/nwUBWEejBLoSVkC2EN+p1ziXSJrlHrM+u/wcsDASBIDfzwUGnWxCwMbQ
AmEZXUIUtPlmsoGTlJIDIHO7JYE7UVN5qUcjCVaXm+4nNKqqWMB4pO3uWm928lCi
XvEFq2IycDbK0S7nTxqD10xtLAII7OQvaH6dUfXO775c8cNxkUpmv1CazkpMYD0O
k23/H3V+kMIS56xnhBKe6HuEeSu92Uwma+wHwH2Yec/As3hSOIiT7ap3wJLw2aFM
OiKPPY6Zyx28NSMP4jYwUHy5ZRhES9VMnY5p89Kn1/6QIVyC/g4Uh02gzuQev7Pc
oaYHsbV6kM7kjWiypz3k7/tm4jES3ks4ygOImoHhf94GghAUKy195d5pwIYfHzvQ
qNexgQO+2XKubHLsdedvsI1V9luecT3mJQa4w40ZEM55XoagYiXjTDeAMBS/2S1l
ZVCbtFXTC/qakOAR/h6g+YFXeCAXXSlZ1fgYTgHcVpM00Gr9VQt27yCEeiVtQv2W
lEQKVgbsUwzAgUxydTqjCDquHWR9oavRRNUQgB0TmqoGpFmBLK136dFXMUXrPdsK
wTfUnssrpMFdKH1kFo4vJQPCv9xL6juIUw+Gyg4YGUrQnB0uQ/Tgbxs+zUSRp/dy
Mkucwz3fcja4oUkNveZprQG46HEiJT7mz8sS91g/0/thp71bc+ATtsIXgGdIn/C3
LU8GNxpYuXg8dVo114mDzWvXJi0JNQj7cGTFjgPARnMutBYDG6Qv33vYKiVLO6K+
FAwIxfxCoLxdlgqYmktAHglyHv/+eQ8UDuE25pE5nndGkDJDkaqXTIrRM07q4KMQ
k3W5971VuxWaLxGE9er3dXUMO84FTePeD2Como5zD6ldtV084hNp8bIGLFAZF50q
Eilf2UNTg5EuSVNBuxnBQijrEttjLHbIrRdD5CRCaCT6LMk+vHkeqw/At6BXSHPl
RZuETq/H3uuMCt2xV8SsF5CrxJ/DI88JnjasIjSKGZwwHK6tiFDE+VhwHPaPjeFp
6UAyVf7ia5psYxy9GHoXcRFf733Zn29b+RRSEwCbajh2rIu4wcAM1ROfWmKCXj0b
9emZlJfzcEDXhAeAp5quGJnkjYthHN0WMt+bJs1ftR/OAH7WZ38wbG7UNiqNBGCu
wf4kOT/OL163N/mXECjNYXsqmMu+WjcfhMimlmpX5gxI33ZO9M0rHLc7r9puH2yc
fkbTqbbXsio2tUbu0dL87iWdIB5BJ7jp/lhWU7ZjbOl7RcZpHG/OKegCsUbYJcxi
9SinbL0Q+xgL3XTY4e9GevpWHEBoTrbOmv8n5438vs4AJIZYDJEimJ5sYWRZfddw
v8w0+0dTp5xb4YZJW5oV8Z21+SUzZs5P4hcd0spRc1i+5a6D1zNbqhYtGYwiAfzE
B29CMrpmVQrABed6CAJeK3MoqCha/vDASKcHYjCLp2gGuFT//SPWv/Gog+FXihTo
LU3iUaVzQ1OGxy5i3R7R98paEWB6W7Ny04LXOb9fhSaxlQXo8REziOmdYTAoFNuJ
owf4I1TDJqz8f5fWCebxOqxHygXDGixzUD8k709dN48dYCnQ/Y/UrNpRnwcUcr+3
1eIoieFit58xjeeecoWr/4wawE3XzwpccIaardiXs0oP6FVVTZifqPsMyfqOWs12
WcOU4N8ckEY7jIAIP/kRWZJzMEty3DxAimyPiM9CtvXxUkBMHnfD6DTBT9RO42UU
2je6ylUfLwchh1RkJatpMz+KcYLP0qOfD/CxPl2K0jfqqvFFLaS8QhSnXIxGz2T2
RiWolrQsZHEUXcfBk8itezKyLtUffFIDghteYVAn3z934Ay4OF8HslQfdl3A/yzw
AoUfCsl10OdNXikpi9OaMQ9jjIAfwc76ttnInD1K97gXCdjGDYwhu41gXgLJAbAL
BYQ1kKCcvbMCACUHtSy2Z+JNgxco2lrsWmWRHTWvwCQuJ2GfN7u+3QNSvhKHGtqZ
ke/ZLSoQ7nFOIA9XZrdd7/AXZKafBFPU9PyrBpKMkY9o3Li9hSCAaMGeJi/c5aJf
uxqDMyM1MPlRF5yd6VwKrN7KUHQQJFAl1f3Dz7x3RK7hw4Cdg890aqcfCGYe4BYg
URgcnnIXTQ/ep8+WUbHJCfl6sfCPf9CcTNYJMIiid4DM3bmAM1uAxNw9iC4e2eHc
Z0lFn6V4BqT5W0QsANdwKMEkgSv9KW9BBRlV5jM6a3cIauXAjEjrrmqkkMjBJjwb
mMnRxjIKW5sAleP1Xi0ZhTGHz35QG3HVfn9ebXHKxw6/fn3zH4RaZVpIP70KAMac
rciYgorCeY28CICuV0ahIaqnMzLhJ3svmnYr0jkDVApX9+DiLKUPuR5H3fg0nZOT
/RZiTM8XpyuJt+M1kf7VnmQr8+FoPvPOOs9GbBlnJX8Tmwsj2dIPuHJ0nZ0nRlM+
ZVtSrg0Vlhp7TYZLXlQapvjGRi4EwRPZR28gotFHoqgI9bI4HNNbZmBKgwjGXc3s
2z76aB3NhUsYN24CZGXiU2cK9RMmYQfp8bQ0t8M3G0ZbBupoQuPefBuDS5Bzc6bN
CewNlBy1nFmS54UOv65zFfESa4B0EE75UkAoOIqq33JNySEZoxNOlikT9Rp2UtDi
/I3oJxbdyQ1NRw1DZChXBSUtpshvwnoeKvXTvzl4jSdEOkhE0PljUuAg1qf9k1ou
uepjB/hI2J/eAOOTDWDWcrIsMVNkUrEd4YzDKdPaBgWI7G/yZMoW87Oe0N9+tOmH
sJFqZlaRWw2iWI1ynMDyJkcImLhjamNCO6+OwPj9NgTp1j2bNom4hnGuoFICXihe
48rXrHROV48aloABE6tqo8CFdRLPql+SWbiiBFuGKVphNJH0R6T7JFuWxCs65ZH6
7t1oWqkry9vlo1WGxsIBSM7t+hMTyRf9Ji0vi9NssxjSg0FMRH6jRY/CkW0xGL7j
J4MRHkFoBwS/jmf+AnuxHCB/3Ia6gM84yzLgoiP0Xvyb53SO61URUxxKH9m2kSIo
iRyJPagb9LPa+R5wLYSf6zspl04e3Y26ty7tEQiO8YbpsPqa80k7nrwn5ERRmE4D
ed9X61WyY+MiNbUV0uJt1eNGJRVK9GpJ2Cp6x6CpLIFrm+sW9Hrv+e6PoM8vINom
Nkx1Cq9A59o97ILIDuJaGpk3/4NL/XzOIK1wn7/zX/vci2pKC1Z0fjQRY+UTsJg/
tH4jEfqlozOhj0IaO1bLcJDrs3IXeYslH0qxH7UnWXNDfWs7u6I/W3rh6Z031fQO
b7mEm4X/p2vxHCINWadR2x/9NL5W1YvS9psZok0wZ01vYh6gG6iAc8CjxtPqEDie
852M+Aydim2b4KU5UjjXQX6YOrklU1ONqWL6XuK9ibDME3HjqdRbRAPbO6P7dtfY
qiyAPzOrR/e7N1LO9Z2VSKS5JWWvTnt7PgErHvTyVraXmQ/mBFg7qBkvPwyuhgEm
vcA4wCVYkZU4Gzt+nafekFKF1BJg0VFxrGpvLtdRnTNyqkwtpQKtujO3z747SvkW
6IRURB/wSKkA3vixudkyMf1wYFYEkll/0laPzowo+OHJvrG2kKE7tfiMrNm77w1x
LCb2rMln1qDn3wANUQB97WBeA4Xeh6Qtw3tX1fhGB61Us62MA6AsuxtAsiVBzFtv
CF7js4anTJYvBC4kj5xXDE+7ZvBKcN7RoWCJIwx/gh8HC0u4Ds1c6ImTwINZlTkq
pwWPpTMht3w56T6Xu+ArwbrH1zDDKMV2eskGJ6/6yZ8Bc6R6dPvaEQPUcUkm/VCc
19cHKqo94cT20JVhBxFT0j62o4rbLRqKjQkKS/VNWy4ZcqH24s+p9HS5pXcGOwxK
5P/8KhabBOfp+95/bm7OOrA/+TfSHKskSIliWmcwUcW1zC+c2yT1W8nGEYswLF+C
cDSSPMBa8TK5YaGBQL9MAfTHOrfACC7NTqR4JNbI6Psx3lwZ3MClbfSWyQtwTkeE
yWUUy3YwOw/Hcb9AD8hJOa1BpMRNtYKfp2id2Tw4N4xFO5Jng3pG54MUWXoBf22r
Q6WTcUzpjjz8PqUKL+u4INXI2JG0DPr3C7mlTVYHfzuSObLBls2SaDKzMekJHPLc
17c+t+so5j1biWRKQVjm+O5DEgGNfWgdxGbJYdAHTvMbAmSQz0DwFdk3J21jd8U7
JCJymhzWiHdPztGdtBr7lIorapMyBM54xNNfxzMmlRNpjm9qNY+YzQcqChttSfz/
d4B0uhYoyJxaV3eHNKKfhVsAhTMA0BzSgN6R/Kwruyud2FBYcpzz63WLoY5fmIdX
Ckz3e0dPgQLLjR72/41y994n7GoUwm5/EkYSKsawtZXFEKBo9VW0dZA0sZNlH2SV
XYjivRooD4+cpKmYQm0fy/VI50T8c3WZvw64OlPS5VQQZRb5tf6tsFXKmCLqE1HO
deo0R3R9WfCnZPwVrwvP9NHXudDNPfVZmlI/0V+YBrdyYfnDYo8v4U/2awdcNBuN
5TtNwW6Ny7ZbbDYx0DnMRKyKI0BvrgRdVkVxugs/yms1EDJ2yC3TgTQTtB36F9a0
4VMOfsVEgJtKgmwOpkN/DI7ZROKawVkZLqL5jtRln7oXWGfMzmO4OkOAma0GDmK0
Jcs5O/BUY4pzE6Jyjqei64XrqpyqNjb5hkPbY8jQbjCB+G6GfyYLKRkVsFnrTkF/
ZPRE3uNAGINoNlWElqKWz88oEuAbdknpGx9vlAOIxm4TTyQnhfSbgQdoB6MBvlqU
KwiSd9/2lafwmW/AxbfXwjIPhg43xDNA8Hn/F835cTzjyx+esznA0y1eclmFkpn/
z1N4MgTkqCt2H9OhG89jct5PXe2F5PN99edplKz8fzYP9A318Ya7ZB8l8hV1gHjY
EO1Nq9BYr84kA4+kiLMrl2G28cYfxuB+nIzTKETdNZJi484yQ24EvnMYoEWznFja
rqOCJE6T6HnIk2sVuH2ZYiX/Ex9Vb/4Wv3AYthotw1PAaXX7VUgaEk+5t5HFtbiD
RvQY3Vs39AAIcaQDqgRGT+Uq/km/H9DoPZhiqMoFCX68d019CZnGHWaU0MTjQ/G2
pQ9+T33qRcTp0ZfC5lo1OE3A8HsH0STwMVbSall0nA0yjPv+GQutEKQXS1zNI1Ay
Zyq/nYRj7GHTlaFZE/isv6WEMQhAeTdLcIGqX1YigmXLm3CZ7YCjvi43KVZ0Sdok
x0+YU44IGwAwlfMj6dAZ5Sz5H2FYz2pr93uO4Xac81xE0p9OyW54LRGpHBvFAhGm
gBKg8J4K3dZf4GbCMxKoGmAZzNlisJy8nV4mVFpZQGLt0fgjirpBwtB1xD4Jy6WW
PH0I0BY0uv3d4njmOEPV9YtMERpXLuZleYKJtDPT0pI4CskmyJEfaLZSwhk7dxxE
THjGN1zs9NdP85DQrFacQkcrAFiDT8fqyJBcSHBvZCggLdctFLZqCeE5FdO6hNIC
Gk6/EMkwpJVp3Qwh/NnkrjzC4/Ysc1ZcyZMezDDKsriGivXm7WJUEdp6FyaF3k4T
bRId9gxcLxiDhnb9J5XR80Y+my361sUcnR8Bg73eUa57kQzNwZe7ImOBJLvBhvul
bYVc3ctbJKt+OnqTIEMe759WzsgY6IHKPLQDwsAKC2reEjazRJLUZJotJgGIcVIz
ezPZ9kHxN+GzgFOrCKLc2V0KYARUoiYW/utPH07QfJqv23Njr9kDXWPMC0WMw5V+
q9WujAGj0kl9Kv+yvnwrzxkhG3nzrFbTcf3Hrq2g2ga5ospGx+tptEviUF4Ehhxu
s484WaOqhCCTerZb1W4vz/ZruDvy3ua70Tyif+etkotn+YQ80N24eGHZmdSgI4WW
lrrIZ2YTH6Z7cKvxOm5pMmS1BTUGKUX78NSKQDcy6KwFpfCEF2Q+yc4d9hPHEd6M
vq6Cri1rmC2DiEK1MgRK53Zf60poDVOiUwfr7Db60HBj1t4fTExTdy6lwmpRH+4z
WCY9AZp8WT67G7zHqzQpNs4rmQIT5LDnVJe27snkxvUhC0Js/TjvDkQ4XBS5aUjg
YGRcz2DUfK4n2sDCaH0DkCXa5xDD2KHjhDrmqsOzhP0LBDgZDaDYWWGGlurYbLvL
t90q3KAglTc0uEa0l6ohFpThR+TJKAX6b49KPcvYBHGtAxzJsf508kbxSLRdgirY
JUUo9HA2lokP7NxG3ZETVbKsKY3zn4NJABkudc8kvBtbXp0RMZHkRdepIOwYgy5v
ZN+R657x9TyyWvbb1ZMh0L8k+h2l60cFsg8pRY8QDE5fuqR9qX+NJvSdbjFuMPKK
nsO8dsl4eV3Axgd/9kDc2R+s/xd65okln8qMIZbfk7iqFYYC63VOFTwTuYk+IzBa
C7TBlofo3yqReVhCISpgIN6JLLFcrcIRXFStqqpR0EDbYfjPq0Nd1+kmZiq6ieeS
n+y8NiPNw6sRtyFdE5ShNl4VlzmKP6jfcz4AqzYHlJ5fzEgewIbanRZ61YxCU0P5
0hsCXPTNpAYIbyIZYICNgSNj0kdSY0AAdnK/dzqeaumrXJb6QinGEQei6Nr0SOaC
oyFWdrWFie2XOZsWs/+OC/ZnF+8DhxmT4wL5UbxTFbAdwuoPpmYzL7jMsj3BxBl9
NApaGFWLKaBU7pjkNLNGfqQFmeWFSoW8DqotY2aZLEgMrelBBqONX0N9KrHN1hjA
Vg3V1fstoC0Esl+nngOoDQSaUQKU+r0hjzKxgS+vdvuHb61UVmwggvfMy96P81BC
uG09JkhtLbt7/GIIOwKcD/obQdUs0HnLwHNQDo6Vaq9YhmA9K6xHtTzzXfuGyPCT
pOjb/cvXBoxDFrW0jsZN9nA3Q7cK373qGq4F77Ko/GIPMDc9X9G2RJVR/t4wIRrU
wlCDmVkltp/diiHdH1HmRJL3/r1u+/IVuEDENlL2uJ90WRlQFQcD+9XGgjb8BB/g
SkEN9GxJCaNOVPvs67Ba5tffWNuhEgKOQLSQOeCgoYtFbOnW7C6yGMPm6vwsDH97
uDxH9uTHvBm2EOICb6kWP3cjUdDIuHNaBhGVWSk6cm5oYhC++XeWkY4KJadrZPeP
jAa1hhT60fzOkTlHs1Ivu9VIsoBvjFhKhJFiTe39Fq/CcQa4+vcTHhjN+Vja+0SR
+0LaxP9gX79sEfdrIVJizIYHuTcYlDqHMLjj+Ga/jXvXq23QLLFk6kC3kb+E/Gii
b6S7gkLdXfyd9fNSgwQ4SxYVBR8EEXvehvHj7Ne5f6TuEG0jVTNE8RsGPb8mHfIw
vuREZmhRJHNacTgbHPTMb+eko8bCU5anBin/ZvJ3E+8hVkszxQLZnpiy2eaXJu31
ZPbkfOWkwoIECAZD1QNA6Bp/fahaXH/fjS2meyBEOmYT+Kg2DhueJVwpBmE9tqu2
ZUScz3b+OXhdILKnZK516Cw1Ba/yg0y02OF+qD9osjCRQwBbBpVKpoWpPxaO21/B
AqJ1xTJk4RT+w+Ik5rYVLOur7a/+w8f+iyeg9rks9NZ8aYPnbWwJIzTXqSdwOdr1
CBMW1IzicL0XD8x2sasGdoerVNAJSoT8E4Hn1XC204Pl+2mVSYgIu7bDp3aqYG9w
NUkSEgwexEHmwuQPcRLxmqPO+UOUG2//DVGu534an4d3MWdqYFrXionvS0JFJcjB
MG2g7rzY3z03jidE3fr1dK7xUxGwpypFMsHlNLnzziskAjFl2FTIoBRZKpqh7scE
A65t9MUCboB3OlMsq3ptRrWBnQBJMJx8XG8NVXIh9Rd+oUG2RjhKatsjfTlhBBSc
5m+sR1YRg+SQVkVwQdhQYvv+pYF2adTU1YXKNvuTmVbgneQD4w8DDwNvO1Txvz/K
9hITUx3+LQMCBVWnEoqN6C/iXdvvRtagfo9ODbc6i0DY3PTsxIcX90XEpI08jQ7l
4DBfex41rZrchZ/jhX2QpcQR/4dnWtdwEDU8gTmYnFb4eC2HgwVW+lwCRGjDnjb5
Mqtu/6C4UPcZCPowAVBjMa2BmC/WhATC4Ryf/aBFRupCMTEQYC56M3oJE8zEtzLg
B/GsJUSoER6I7AlE9Pp6XV+xdlgw/I2/vvd8TwRP+g8LaOk4sB5RiFPy0MV3hx7E
odZT+0HcL/PtlNX0416zXcCs1p2ehItT6J+h9+1qp2P7q8TScLSYNhjuLCsIt3oC
sJdVkXjXKPGMoww1ZPpe7HyYFKcWbZW7Jj868xo0Mk0CTTyaUvnt5F7zw/I7Yyxr
kl6W0aPbzrK0mlUSfNH1dQ4xV2KU06FfobVfRvS7I7b5t+H7han6lRdsgHNTgwr8
zFJ0Iye/h23SXtvb4s2a/9Oh7E8eKNSDUwL8/aISKKs7zo60fs4uT6fRb/4VbD7o
wyCvkR1tjbMq1FtTKDOnG5GldQ3aOdLiEC/dPG75p1ORRU1etqzI9uuKdwMxZBnq
7dCSVgS9jdLjivaPoshQVr5jdQRXHihobyVK1jv4XPyu2QzTR0yff2JRtvdrAMPY
SkS5+9sodS+00GY0F4dyLV2T7KrbhTFJdP3M1o04kyGCWrRYjYx6YhQJ33czkxeB
GiU0Z/q4oPDgrBSHFoxhpbqFtwyz9bOxj//51bgyf8FBXcynb0wy6213pBal2FLM
Lx0F5QdPvxdtvruuEYmk7dB7HwvOo/JVIkF5N7b46LFJQ6SRq/HMqtTCggneaYYr
FcmbDFkBwyetIbMLDc/02mfB1mwKL3H173b2W7ZRyqQFWRNF+MPBkBryOhtIu0O8
KYk9bmwb2zaz0DoVStFD6uIeKKF9YrK/Zv0w8FPfD2UgwNBBLWOZ3J7ZjnByQagL
g5CyueR3ydi4vkYYA5ya3aVpO3dlpt0YySQHTUaj6fQ2Z5mfknx1Fa/f9jx0pmSd
4trlrUtKjZyMOc8m0q+0G0RJtxojnvWwZqrZ89mPtemWV/W0OJwhdKJM8Fa+j9nT
1AH/1Ika/znVw5NH+wKd8vaqJh2gcKjVH8IMLUVRla6PLUmGPPuMXNxtip9LKceM
FT3EFHFWBfqBmuK7lUyBqNCNpMW1QFiajoLN0PcYsLpHucAArnjbPkhDb4rqeW6q
ob8QnBDeE0GQps0+HdRr6bX92TyPCYwiYjhNjwTEmUEs8yMMB26ex8Pyh5MVE/sZ
tHFNwYjuj1cm3VKFX6qNC0iOfM0VXjGasNgNpKStxFHiXHNIN8A0RaD/CoA4WR6C
+tIjHjECqyIeHaB5Wn7+NrqnWilIbyS1BrA7LBURPHzLsnHmLYiW+GlaaCdfYQB0
cPLU5btWYjvt7sVcfQa31Q==
`pragma protect end_protected
