��/  ��^u� i'���^~TJ��t6��O��U�]��V8�S��/!�(Rݘ�1@�gnѼF�g7M��N(H�YA�[��֮"4����'����.6��{S���f�F�q�ߠ?Gc���R���q����k $��l�t�ض˺��&	z�Y���M\�9߀���Ơ�/�hLy��8��֥����b�q��h���H��� !HO�Zc~�c�$� ^"Ƽ�����B١A��Q��r��M���C<N�����Z�c�wg�}F�	^7��WOf]]�pg�O�����,�S�E�Ҫ�Y�K��b`�k��E����O����a	_6�CF�ZIqx��R��$cuNjmˀU���(�C�v?%,D�L�AD����ǒ�˃���<���+�X��W���z���Y�e���q���7Ph?�W��OE�IQ�.�q�����<G)=���?Us�� ��faNX_tt0\t��N�H��Q1O�r��9<���ã��As
.=w�0O�tg2��#e����q�J�tGCFex�>��m�b e;:1�>U�����&b�IꇤS�g:0\.����lI��OwK���`a�@$pC�t��}���0��5D-�.�Av�n�$������m�b��↺�,��E4�B� �n����R	�cpE�Y5(��c�P#��|�}���ޏ�D���j���V>��6!�n���q��PcO�e�Uh4z�l%�l���Ĥ'@'	@L�%D�x��-��N�U"��Y!=�a���gB�,�N��f�j�K��'$	��|A8�B�?�9sʳ*�_2ډ3��m�Z�Θ]_�iZ�=��jň�M�1Fb�{�E�W���[�[�g���` h��T����}���B���Z���,Q)���^xı��p�K�f^��"��:\y��	���I��14�PURB��k�A�)׭���I���<��`�?��+���L��l�,˨y��w��F%��۬�&4��e��p�
��F p0�*��Uv9C��%��gt�1�9��/��\�7/�F#ƞ��d�}�S��_,-;�� ��h����5c��ꕲh�f��8� P�x�9~dS�.�$�έ���E̝Չ��d�ϗ���놾��FU{/8D��q��8�v��8���o�C�e|�9�7�ɿ��@��?g�I�|��7���.�[o#+�oܽ���y�uVTE�?�E$cxQ�>�m�޻e.�YOXC���퍵���x���êv#���i��(��G��i{4I<es"60�Y�]�zj�7��!;ܒOԘd,* ,P������yM���d��o�Mѐ.��o3n�e��̤��L:~<��[)��g;ߝ&��<�&n,�M<�ո-��7���S*�Y	��NN�Y#!-��:�T�n\���͢F����A膦�apRP�ٕ ��2Lɘ3��W��e�q���K<�0G���|��,E�P���ƒӖ�FpG���Y?��H�쮩	�sS0gM���Z���GO�x��Y��4�2ay��u�H7����}ɘ|�?P��OkI�Ϡ�L)�s�[�RZ��5����q�x`@��u�I?k��� v�5zb ����0�꘲Ef������̼�12�K�d�'�@�d�A��A�zFs*�z�)��)���AĿ���b�D���4�T����˝@�)�q�oqa4V����m���Mk�&���ꨓδ�s�;N�_�R�l"��Wn|��Št����8<���a�b�>m�dB!G�9!��#:��yy5��/��.G^`�_,Gm���	W�^�k�7~���RIg^e<�4]El�_!x�|�Խ>���RtaϤ.b�����g��	_�9�
[(�7��{;�5An��
�|��@� ��r����
�M#Q~\��q��zK��.ۤ��7��d9�`d�_ɀ,7�x�+�!�M���"yH�W}�h#�0�~�����K��j�I����W�DÂ��nC���Ӕ����H��)2b!�t
��>X�%��gf#�lw�OG�+}Zp���jFhO�3/��G�b��C"0�3�s�������P����#�4ă�CNW �����[1�z����R��cY�Yd&(�}��[m�}�/��E&��nm��_I���b~/���l��	~���+nk���xk�ħ�3P�ێ��-�� 0�N�{�f�X��4ێ�`��톣o�|��k>VuA�f/B��H&ۢ�m�?wnƠB�i��G�������P:��J�l���(��n����&qq�-�hd��z���Ͱ��s�\i=)Evh4������N���l�����D��:�?��VD���7MH����C�$��1��2f�S�W$G
��LJ�:�요�'Ř�uhkȫƾ��Z"$�|�IhX�iP#���a�X5C�l�+���f����
�&E��?ig�ÀI�e�1�k3�DC�l�������MJ9W�g�U�\ik*q4U���ɓ0B#�Ћ�9u'�zg������Y���}&V4�̀�>�)�y2��3)��;��Ƹg�2���ϸ 3�c����Sn�y��]nPl�f�^G��@�V�KL������x-Dn�ZC���7�w�'����S�r���*�\��rX��/s�?"�c�n�3���Azҷ����!T7b�����~]����3i�QiP��m�-� �`gv>U/��`͡�_�?A%O��`�v�(��'�$�c�x�@'��]�Y΀�'/ih^IM�-�7��� d�=2�>Z�'��~�=[��g�
�*�y�>�ou�I��6�]��l1B&jPj�B��Ç�ط�݌�x���'\,'��.�ꃿfX�G�g�H�鏄�PUYe��@X�	ԙ�����oP���+٪�}�;���ង+��Q��t2?�6�@x�`��
�_>"�!<	��B)���}�؂�w0Ӌ����#%A8FrvEM�F��o�s��`�T��7u�m�m���֯P%>��	n��a�3X��̐�!ְ��@ԮK�,��8�.����d0z�f���h���gW�}���( ����e�#�9F��QML��G����Ó��3^���E �t�Wj���Oh���9Bf� ����(�ܭ�l�L�M�
(1������#�� �.3���������U�73K$�`M�C��A̤���e9�]D��T
$֒��z
)��ћBV�\v�ʴC�<\@��7%h�,P؜�)s�*�mHn�D#���a�Uv��t��l0��U��o<��*���od��EV�v�>��t���nֺ�~��O�j�#��|�O��*Uhů/��5��zcf���ӈ����Л����Ǹ��c�d����i�ǵ�9 	r _���>��L��t\�_� ~�l?�(�a�[��Z�{X��m��<?��%�P�Ø�� �ii;G�7����%����{r�:.����C��y<�7]��B8���Q�+��Q4�`�Om�b�ɧ{�G.K��i|9�rt�P�6c��]b+��\����H ?�~�Q��w�#/����k��2�Գ	>�5��q*�ǰH}v�@���'^�t�#J�Oo���f���ۣ����Et�'��.�·��m\ �+��`��sKl~�H�g���	#���ҭI[ 8��
:�c_Y����f  (�WxSV[�Ida�J�(�J j��7Ȳ;G��5��u57?%��(|��OY3[5FU<�����8��ߘ�p6�<��g�r��%�7Nf0��i4��>x�z��ck�3׳�=�E�fykе�����|�" ��-�����L��؝�Ȏ��:@M��)a�*��X�6�+@�<��OQ�k%�ûA�m|jJx%��Vt[���r
N��g���+E�n:���À���
�ڿ�c��*�0N��)'!��8��.}Z?w�W)���4���@�B�o�s6$�F�����!y��F��4@�Gz���b��p\01מrolձ3�2`fUw�]����|����1��I�bg0�+{���E��Fai|Dq��I¿��:
A����$�q,�l��ף((Y��Qڰ���C?c���Q"����/l�N�s����{TM�S�m���� R�����F,.&��a��%R��rJ�Ӂ���j�ٺ;�ʦ��+ͿUx�-$m+��#�S˾�P�m�����E�洊�q,LO[�@�nP�V-l���X���9b�ߦ6����d��M�6��N�A��K5.?Z��c�$�������Y"=?s�e�X��l7����Q�چ�9:Q6�M2�Up�M�����h\-/th�Qj>��=��x9�����7tO�Q�����]2�U� �ܴB�Z4T@�?��\��y��4�TN���v�[&&��Y����	��L8���V��׬�9���\\p�ބ��)U_#���o�C�VE����)�j�v�ȣ���uy�ۣ&x��Ph����
X�|(�$�_!���in��Ɣ-�fF?�B���\١k��>�\��~�޷Wԣ�ʓŠd�+�Cd�A��oF�u����}4��U�P��۽nrJ���c��D_PE�a��b/6_�p[1��Wυ�<�eMd ��.��$W+!��gI���#�Z@ϤM�&����M���Bv���4e�����e���_B+�=㺆w��7�Abדo�+5+
%�]���ٞ��D�Y�\��萅�i�,�9Xd�x͍��[+#�(�+0�B/h�j�'���u�~� �o������\�A�Hz�-q����jm�����"�Q�A�W�ү��&�Ȣ}�]��s�^A�b�J{ �[.Ú3w1^�%Ѧ���IW���F5�����	�mx\.���2f�FR>��7����4������ٝrR��vX�co,����	&�ִ�ል��;��'Zv�%��/�/�������b��Tum����l�f��iTk��Al� \��4[�b�EHWzY�����6�$~�XӉ�Ƴ�r-���ݵl�R��c�y`��c�\�P���.#�& m�/�0���	��>7�*�Tx���@'����󵎆�{����������9�F���G�l����'?Y��V
WI�#���*z���r ��|��`�t�U%U!�b��%w�ߑ�j�����	���X�/f���(��t����;�r����}�r�˃��@�m��`��:O�θq1�&
8�0Ғk�}�yħR���Ӳ��P� O�/�F�N{%�Te6F�h�2��C$��J��]�u��''yIc��b4'�
�J�G���q<w(�k)/L������H��=q���p�b�v���ٸ�����W�o&$��x�����m����P�f�1f&��sLi��+!�J��*�jԢ���,:7��bsW�q��4E0��Xg!�CA���.0[�ń$�к/q�g#�T�,OՅ��0�y��$V/i��n�����"x�c�ܾͳ�iP
�ș���w�*�(�,��ܦ�� F{$�'l��ιbx��S��RE)c���mW��
ƕju����زa��L�V�%�Qp�=W��)S��������PEx�g��=N� �U�"@�kS�"�N4���zR�Gb7z�]��ͣ���H����ՁP�Ȟ��lQNM�_�j����o��s
����2KX6��
�
�te
2���L�����ûUU��,S8|�A�?ʗ�``B��Jf�����,?�./M=9:2>�J��7�J�D��&\��!8��,�`� �-ʦ$�>N�B�j?b���ų�W���xES-=�l���9a<��l��,���}��J���m��T�c<�֓�԰�6(mUYoa� ĳ�7��n9�ƈ�6��=��x7�n�n }�>�?�)�׏p����PF�Z{��c3��vq#�嵾���.̇q-*�@�(pE�[��af���VoE�h5�.����'\7U��n����S���Kl�����F9�QRiʿ��xU�[J�B5�Ѽ����ㄴf�h���Ŏ�(�f٫-*��:go����lV����Ǌ�!�����Hlcƴ[��(�A�E��<��<�%��,���#HNh��~ؒ� �/���ͺl��zG�͡9+"T���b�x��*d}^���?�H	C �����0�����,&)���������ϛW� �ބ8r��������L峏\|ryF@��)I��aݵ I��eO�V@�0�%"�44������s w�ͳ��T��皘��-��Nk�z�X���*w@Τ>4��F�G��;�UmÅwN���������,ۑ~�����Ժ�[�,PvM9�0������o/�-^����$��y7�9���rI��K�C�n�z�rl7y^�~�5y��&G���1.��<���&��X�iGӂC!���������h�����[&��+�Pfr�o�3�ͮ����_�pͭ�x��%�r�\5��rh���煚��ӈ%�C���"&o^�>*b�k���Ҏ����((dG��� �����
�i�*��K���}K�IS����o����@�]J��V��t�����,Q$j�W��}@���O���Ē<�z$�P�����ꍄ�۪{�ώz���D{���Œ΄�ux^U�
�E/(fA`j��L�|l����M�^Y��x�������Z��z��uW�)m]��+S��ѭ���3&$ U���/��������ϳ���bxzu�8t1���/	�A�:�o��0pE��7��ß�/(q�[��c�������q9�M�%���ۆQ^.���!2��#��xbeY>>�zWH�ӣ!MV�X ^o��?5�/�O>�!�z�=j-Y��ū�f�o�Os,y�U���_d<��f�C~�n��_�88cq|��5������[��a�:�; V6����qF0�陑�(��N�Ӕlg<�O�1� �"�Yg�;��j\���kU[Ƭ�y.'f���b��Y�Mz�Ocm���r 0����g�����/-��n�x�{�,�����E�@զ�_|Pʟ�6��/f���V6ivW=gͱM^l!�I[�ϕH(��MJ�;���-��P˙������E0�'/7���sN��i��:���4�:ѝ��2��xe���`���.�Fr�={Q����x��+	����<�k�W�s�0���I&��y�"@�� 9t��j{��L}sM���Y��vƉɼVP_���Y�(@����L�0�bbw����p��kV�#�����:�޽i]�oP��~8�P�0=���Ki5�y<Y�.=3�Y>������a%�bE�վ�P7T���z�,rJ-��  ��5�OdE��gX��e��"t /%.Nb�Ă��QaÊ���y�^�)3��=q�E���a��7�#R�Xn3]���6_,�C9	W,4U񍢜9���`cͅ0	&N���ߩ_�u�|�8v1��r O�}��$S?^[�bs��5����X�KM���(�yz�����fS�?��S�g��܅�}!"FW=@{r�U̣E;-ko)����(ӗ�Q�9d�e�+�_����%�5���R!co�� �wT����VO�@r�k��N��Ť�"�4�ް��kL�=z]�a�\�O����ɽ�ת����j�-��M���z$IVpt�o��G�3�4�Ī����o���z���<�i�r�:�>��N�`'�y�uH7|PcL��?Hs�uLx�}��R��~�"��O4�ʸ����G~?=�){��$�hDd�a��h�Aq�����4�V2|4�����֟a�b�,�l�ˢ@�$�ˊK��b����?n�Z�����}tx.JX�E��n�u 6��tF�Þ�6����.@�k�r#�##�o��
j�3mS��J΢P�ɚE"F<oǡ����#'~\��v�W��!�5S����<k� 9���l�NEщcyRx@�L�!Eu$�B=��̳\�t�$�s��4ϩ��(?�ִ�L�:͒B��Y��H1�ÄTB�C��Ʊ�&w�`W�U�e_�i4T�^f�T��d���f>C{�
뻃��9�@��p���ME����j-%���������=�zq	 	�	��-Z��>n8-�=b���5o��ɜ5i�4�|H��ŏ�{W3����ðQ�/���]>^�Ļs���_�ۙ>����W�a�ێXw�}��E���2��	��纃U$��/��dF*V)=|��Y��G��>?z��9��X�$�(^8�Tk�3�ݔ�x(b���٥`��.�x���EeWik�W'�\_��邒���>I{�MT�H�k*��,�~F�*=�a`���5%>��5��������ݿvL�2�����ZႠ�^�[�H��\�$Bݞ#g�ˤ���kUq�J;����J����(����fТ0΍�f�{�B�"T��y!a���@�=��nv^֚;r��k�l9%%`"{g���s^�����3��s�Rf*`���j��T]���`��ag������@r�s�c�|�+[������ |+���I���
��=����f�9ʪX���V͂$�pR��l0��<�d�)��blOR����~}ͼR�?� 9���fA�DwY�(�g�i<'��x����Ku�9oa���Xp?}0��n1
��(B��3*�.�}b�`�<�/Љ��C;��+(�Q���E�LA�9#S� wx����u=Nd]�E*�r����nO�ZQ2TkÕZ��?Iǉ��=�N�ӳNW��R{,�e_�$8��g.�'O��T��M?#=j�ۖ��O���X�0=~C���*�}���X}�<bX���1��KP.1@Q��P�$֭�����:�wi�M��zk�,�,ro���v�����b��q�q`X취7F+(|x|�M"��]<u�XH��e���ւz����;��˿��\(Cp�d)kV��V��&|��U|֭����6�|=�@;a��<���a=�'���mꉰ۾%I9�0A����r�+6�Y7x`j@h¥z�M�����ːZ�\F��W~ ��X���J�����jٯ��X�z]�F���` �ܣ����r��%P��s�4W��S���i�ɓ �S�j�&he4�ڵ�	����(|����S&��^�R�ɯ��������Y�K��μ
�S=e��o	�h�>�[@ �{�By�M�n�	�PO"����Z�Ѓ�ax�`�l&�!T9,H{NE�p4�]X���N�T�]\��s��d%0��+«�\�5x<�����qN�.]>�ʝC`���ilz���EM�6�	u�$
3��Gv��t;��r��`_�R�l���tl׳_���i1�0��8��n�˔W�_8Y���h�o Q�@L�ы��х�ɷ����O�R<�UQ;~u�u^rNغ���V��U��\�
�,���V�}F<��v�%o��Í���M����V���U��z��Gg��eԝ#ky�7xEI+�/��~��+��+�����0����f�'�,TM�Bwbz��Io�8彨TJd�
�E���ڎ�_�O��M���u��R����gm2�QI�i����/��"88���U�:=#v,Be?���K,�ݛR')����3ZIF�BxI�'�l����AJ���>�T��}�3ܡgeJ	JX��>�̺����Ub�җ��:��q�:��v�R�:f!6��+��]���w@�Jꢪ4��C��3��{� �챆9V���.�;v�w�[�W�jd�	�����ژ�*^��[�G��N�ߢ�8����ZU�R����+܋���.�{|Ձ�a�]�	��'��¸7T�v���I֚�ζɲI�$�xX	�\,��_o��)�js־_��R���<�[�W��*_p��&�dÚ�;C���Yn�Cl9$0��YRf��߷_�L��H��5�L���p�w�q�/�8���%��3�t^�{\�w<�u�����9�aǒvd�Ȱ����p��(�!��d�^ħM�\w}�1�q�:�u��qOsn��Ɩex&ɭ�t�,�6��������sq[@ņ�V�rgY��Sʿ�"�{��|��&6���g�c�~o ���?9F��ƬV�ԁ-������>��q�x4�v�+$�MS����u�{=�g�.	w��Sx��eD��P:�\nP���Aa(� Y<�� n��ӕ/��`s`�ى��5)*),��~��H��垌B��+�qGq�R�T/|d8��:.�i��I�6��z��ܵ�����@�t�ٚ�nݫ�b�;�W훞�Oy��1w������f���k��\�֭<yߺF�:iHY��VFd��#V�^���P�.����ĕA�.b�y7��M���ϋ�^{RU��]H����?k��,^��*%�%s���s����;�^��Y�7�?�F��ʜ��(AqO�<r�l����Mf�F��16ث?I�d�>?� V��0����<�u������Ne[Ʌy4����%�^�p��T벶�_�Rm�Xv��<I�M�q�Y-d���5|�w̒cޝ2�Z���u~IG ��)އ���V۴\if�PC�<N��BQD�[�hN�I����S�{�	�RO��M棓�C�x��`�X2�ۺ#���2Qm���3�a~�R��������A��)���̏T96m�����$D�P0��X����I��kM�qNR�dw�%���ז��ĕ�|�D�_�r��>+�+�%��AG�[m�u{VT9w�mݚ��
���?��D��2�=H������ �]H)�ٝB��a��Ħ%�NKD�Z���3'J�a�F��˹t�џ�m?h��^I����H������C��r�kg�L����[u�j�pS��Î����]�F��&#���nG%O�>��ؔ)��b�N�j���r��9n�o9UjE�bM*�R�f���P�k�)�1%TT�٘j�է�d�q�U�a"�Ϣ��+|�z�F�!�!+H(�]���{"���x6��%fŤ�d[3�)V����y9 ��4q �c�P[����9}�S9*�{�%|�N^|�ꠇgv� 7y����]��l Ӱ)��+z}qG<�l���N{U��ɴ8G�q�[��҈�ܽ����;�|e��C�ȡ5��k	�Y��g .sV ^2i�J��v�x��tV3�oEr�B�����,�QC�^&����W�'�e8���(���N�DM���|A&Ӆ�M��O��X�cj�E��uO�Iר�\�ES���8VH���͚R��Zuc�$�ս�ڲ	^���O�>W:@����@��[� +�G�wމY���g3L� ��Dw��ˈ�NRfΝ9��X�]:�f��<,1�6�P&J�W?���Kp~���_���Z���1��K���4�|����KFč�Ǝv���|Gu�O,
3��]K�0m5�36�u^v:=
	vtO�
#Nڬ1��Cr�M��IxW���_JS��M'N�!O�@��T�o�2��b��;����ݼ��ۉk{m��҅��b �ś�_��veX��>R<q�w�;{�2�s}�q�I�����r[��j�3r	�ꆐf�Q�HT�hX��f��@2�K�r�|��~���1
�n!�r����;{�Y=SO�[T��Yv�O��O��>-�p 'U��� ���I���A�xJ�p���a`�+���Ycr��Mmf���/M��nL9�W�/�	��z8BpȊ�V4��K8fRddU�<���]Pp��V{�w"�9Ys}%U��J�B�����^}��;�{�1/XZ�W]�g�V0��"��s��]��T<��M�nP(�{�JK�; �aɺ�з5Α�Ȃ»oT
{���m��~V�!�oÜ����m&B�
%���M!�Z�Q���`��.���L�ҏ�uh���)�GE.���B?�pLuK��)���Ij3Y#��шǳ
,L~��f�5�d���2-4�^	P5k� r'}H��mTwJ��n��4�,ɍFNUv�Gc*0���
�]C/�y���)���aɡ��_I�!�q��ʪ����Lw	]�o�0b�;>�OO��qtTZ���^B��K'���g�]l��3L>��^��I�3��7�˙@�*"|a
�ojƫ���Aa�b�xkU����*$��e���X;YŎ���|'�����ڬ��[��8�>��F��ݟ6.�A�5����)�/EǇ"��E���ޡ�S�g�����O�ݭW*��x��G�UQ4^m�4��wfN&�im�t���ّ9HȌ���U��t�Ƭؗ�W�d,�Ƅ���(�������޵y��]H���9���}`��ÔDw� �\����ޓ����b�cr��S�:���e� h�y���A�D���7 �(o��e'5��\`k\#�|��5�,�/Lwt�Z�Yk"�\�J�NW	�%FJn��0���l�H,� ��`&ru+�����<r>��W�.�(s~8KW�43�~ ��>��:�l kyS�uH�b��,�>L�;��=�b�^���b���Ջ���'�d�|P��1���Ak�yl���^�H=+��_Ox�6��'�gίE�府��9GN��a�D��*r�@�\Bs����`2Ą����A���9%Mg�qŮU[6����;k�rs���5~��I '��ٽ	U*W��1t� ��y��oXjM퀋�G��c���f�0#!�����ueY%�~���a��q��Q ��wмS���(<�Ľ��S`�UQ���6�_�D�(�������K�,��0���l�5��qe!=��.������p�ߖ~�k~i	C\#^��"X�C���Ԋי5LLnFNߜ$�S��R����O���9�R�~ �5�4$��4�@g!��N�4E{�ӌ�5ҥ��fK�ƻO���E�\t�������J������E @�'��r�=֏,wATn��%��t;�Ø��ۿ��x��H��_�.�Lqc����=D�H�j�Via���������0;nQ᫔45�h[��ԩ_ 2K���l�v�kR
;�]6������
t����4����;kR�y���C� ��7�A�.�����m$�J�RG�w����Akj��c�5�0�~�:�?��V�՗��=���>��'�=�D��m�h#O��G�厨��ZM�b�KR��u��l���ݝ�u��:,�eٚ����v�f���uߜk9/|��]�X�����b���R^�������@(㏤S�tXG�N*(�YU=qRc.?�K-�\��]�֢Ph�����@8:�Q�Z3����R����4z��`^�7^p�f���� ��?Q9O��َ@���!ܡ��R�Әn/����iv�#d|�E�ۣm^'	;�Uz��L"�u8
�
�����M��� ���,��>���.L��ŵw�>��x��K���;�I�N�K��Rr��k�����ty0����,q�)�;{�U�?I�z�Ww�u_{ԟ(����.<f�ipo*|?�q��B6��؏g���Ӡ/�/���9)��������J�P�2A`�r}�ߴb[X�#��2h�Z��$�4�T賣4��5
�e+�	]�ovISwC��ꥹ;=
6��s��xv��6w�s&��FA�������)Š����e��M[�P@y�j˒���%�ʂ��2��f��	���cܭ� �$�ȹ��wO�%��K�@����AT����)W2kux�[;��\�_�ͬ�(�?W��|6�6q��͖�����$��NG�M�mF�20`a�ˆ�5�*5b8�~�E��Yd>��f��e���9*�'5�$�{�;��ên准&�X�XR9�6Y2$�q� t��ߟ���YI���(܂��bF�aQ!����0s�H8�����L2yI�7�y8`L��Q�gN5��>SwNh˚�wb|k��Cb�A��<"}� S�� ���>g����[B��A����6�?��Q���,���t�!���>��5�S�{����m��6kD����*���F%����m$	q�:��A�$6.��u})����	$�����2��
Eڒ���ߜ��4�T��ȋv��1�,<���NҠm�Es Ye�X �br�O�G, � uw��a��'#P<��y3��i%��N��3�9*�Ѽ'r��d�ý(<�T䣟�(�QS�j�~�<r�H.��+�)=!Q� �
�ۢṳ�4�������zh�����ӝaZg�B!� `X>+�4���Yti��ʁ
�'�{�IG��Z�sZ�~D֏��3jS�_`ZC�JwΔc��vn�_i�/�>�|f�tv���X��!z@��"�k�]�c�I�p��)�r�P�D�R���o+��Q�S����F�j��p��\}�!�"����� ��K�O��=bf�Ҁ9F�ni%i����ڇk��}�^�n�|��7 �Oax����щ�M(���u��IU1��>������`l)�*Mk����(>&H�)�ME�_d���#��@`7���|��DjA�0I�H=x�.��B�x'���Y�8ܛ>�7���X�[�.�zgf��"S"�Z�B��v�߄$�3;������!h����k$����G�qlW~�^6�2��f��u��8,���D�s�pJ��_�:p�}J������T��/;�Օ�QQ�"���m�k���p�U���*�.տ��;��ȰO}*L�s��*n@F_�r��ԡ�t@|̅���3/��?		`L� ���w�X�'���T���h�i�*z�����p��Q�N_���63��m���N�A�_�3Y���vr��\���q��z;,E�$L�n�La�H��/ji�j���ݥ���T&
�J`j��=�g�(����t8������L�A�(1
ơVw5"�TY@�x�~k�ܩ-�]�'��c�H�"'U�6�Ԕ-e�F�*�'o��MS�X݆���4��%��v'�e��2�l�p��V���� Na�*todQ��I=g�\�sY�M�n����k-%ʃV%m\��zC�򼆾]���\6CYM��1!�������z��ݾ���S�80]�3�3]E���e�o����Mnп�J�e��Ne�c2+�*��^\fJ�%��������J�����
E-�x�W�FͿ~ժ[�bߪ��-��O�|�2~����_�ɘny�����S>g�I6�BW<�̂���y��	!��խq�<Xޚ͌H ΅�N'�<U����_��`ܒ[3��;�p�9%�ͱ���(r[c�ШdA+}Ҍ�I'pʛ�_9��n�����w
*G�j�i%�mv�rK|z���j�H��O@67�	"�,܎ƈ��&ȶl[��Q^��}��8$d��)J�BBX�~(�ן��u	�����<-�����	�i,u�۫�ݲecb��M���{�N�9�6����N�9a �	92�	�r ��KZ��i���0�	 �z)H{�
�F�J���C�k��6e_�6�
v6־l�}��U�_�#AdP���� Nv֪�,�*,�eC<A��#J��ZL��%�m��#��/��(rk�opi����� �^~�̄o" Z(��S�A7�|O�s3o�*�qm%[qwm�V�h�U�2���T�d�5�a�M/�M�c	�+1o@U@ %����yر�#����PIQ>�4ĉ�D-�
/�*<*��~��n�3]v��L�m�}È��:�
K�[L�]X�ycXFQ}WVubd����5��ܬ�~-���ȥT4�#�c��"oBQ*X�����
���	ȎM2!�g��l>y��+c����]qrs��F{���ʾ?,��"i��D
��	m=�O�`+�!b��M�+%"3�Z���Qu-�=��M8���l��=���2t�@M����
��^���%�l��3�-UHsP��v�x놔Rl�s[9p��@�>�F��K{'c��t�#��ϺRB���>�z�D��T��d8ɹb%�k|�}� ���[�^N��* �sC���)�M�$~�I�mZl��_`k��e�����ꌰ҉<�ټU�Db�x�C*0O�c(D4�"3�5ԖҮ"f�S��S�y�p ?#�GitXo�q���3�p�		bV;Ƈwg^��7Y����ͅP�4ƥ����k^���rh(���K������ю�ݗ8P��z$�	�?+P�l��rXm2�Ek�6@d�S��R�H����%߇�AQ}�oM��x�aB�̈́�Y �\����o�4��{#g����v�I�m�G"�ϱ�~(#uy�����z��$�Pe>�[��Q�Y�e���u��է��<��42ႃ��5�AJ�n�p���mG<@�M�a�ƹ<��&vW�NVЮ��H��kGv&���c6��:�s��G�i���yI�Q�(3F\(>h|�J�,>�ks�}�cw@�4ߑ`o���:�^��T6��N7��>4Ttf�/g�
��aȿ�$ݤ��0��Q
ye���P�aQ*�E��\`�!6uF��loz��U����4;��X�t-C�yi��D���<���Ƥ��դ������1�ÔP��2 ����;��{�k>O|j�"�KU�Uw��0 �(r[�ؓ,������6��H��)��� ���C������{��=�୑�����U��S��	`fFK�9S�<�t�t�.�9������ZV$��`�0����'��k��{S������~�t���D����m���>�Hb0��r}��]�ǲ��/��O���iF��J�������ܣ��/|5u�� �<Ui��%z�l�ڝv�b���=["�~�$��m�pfy����9>_h`K��� -!��}Ey	8F]��=�Z`��妿b���I����BM^�*���@1%o@�u����{�ئ���!�^�ɋ7L=W�1� 0qS�P9�)����Mh��Xy��^�n�-9<m����^���c�@f�Ի��䣨���a�\H�����{(/#��<��ɝ&�(��]r�$����u��ȋ���we-t��նC]�n����7B�*Q~���o����^�P��>)��w�\��;P
�FYC����E�B����7)x��^נ�h5������Z��i��XY�" .�9� �N�K�e��Ù����Ǌt���?�3�Ѩ{<
+=��],�Vx���l�ڦ��us��3�'G��۵̿ Û8��2�����������l��p[��R�Xv�	z�p������Wr�/���_)C:'9��H�P�K��{X�/����y.�OHM�M&�C:���.ژma+�雎�;A��aE�5�7�iQ;�U�g5uq
�ŧѲ2As	f{�&�B��JR|-~��5C=�$�n�m^A�d��*�c�����7����z>��Po�)�Qe.kSn��b�DB�-���/��^�p��.-+�
�e��٤/�h�P�����FΙ�~�+/�~Xlm�E��ΣD���(��/����g�yP�
���_5��C�_����`uE�XI����v�I_F��͊��oʳl�6J�4��Syo�τ�N�c��Kt*�'�Ks-�F;
It)�- �2J .�e:���7�~8ȃoc׋��*��̑�7Ֆ��oI��Gߥ!Y��	4��ԓ'�~�XN��jܚ��/E���'�Dx�����_��k�<�v��)� @%y�!�t�)}���Nu⦦8'�d�wo.�y����y����E��L+�bp!�e��6��VpsC^t�U�ERd*����qd,Ӓ�-s�ꖼ���0(�;�LӘ�h���)��H#&���t<?�C�����*�&;���}���\�	.�sQ=���.��J���sEh�Bf�V�oΙ����b����^X�I3π�*ݔ
hn���N	]���-%��Q��,��Oߒ�"�R�4������Vqw�y�ZFTE��7+:��<�gݞ����<x6Y��U0R�h|��P�T��\��� �CG�<�X�D�ZXcE���L���U�v�4�6�����mlp��2i�K�,�R�-��n�LyIƬj摯�3)��wb��/e�X�W\�{�PA�� ΉG�sb93ka#��	�N���@�a)G�m��+XT��u��TS�DjF�䀅��g��~��,%���$�	,/��QV|���P^t+~���U!�#l��=�#�#�
ҳn�1��Z���D@3��Ԗ���g���P�*��~�U�x�E���C�ø�����u��C+��V �v �.��N`X��/��R7��?����ǰ��,������o�:=[����t�$�y�u�|�xP���� ��J"n�����K�[��������ߪk��J~FLA�^�k5���0��G�}�KDp�N�j`�gY��O�ۃ�/E�*_0@ۧ���N#�'�%{1���+�؟B�j�Tտ�w1�a�9 (G���bԙ�!��0҃un�\�j�j��M���{�Qp[����X�\ 8P�� /�n5 Cw���h�����#ѥJ���\���G��	�,
M�	�sR��!�Xn�I�ߏ��nDfo�J�IKp��0��,���y��B%K���gk
�;EeE;����v�/<�'*�k� sZ��Я_��%!i9㸽]gt�ː�_�:�5#�˄�a�oj_>!Y�W�$ɞ)�����8W�t��<�����N@[O���t�ҡ��W�SذԦ�3����*}@'�ZU��[òx�zj+�.M�::����*|�9�.@1C.�ٓ���S�@�SN {�c�˽@�NA�}QM����j0n��i�g�̴��������:�+�7��!*���ƣQg���&C�8�c`%!Tm�&�n6@Tl C���^��_d�,����~%�q~���{���po#�Ҁ��:�կ �5��+��B�ʶ�2�9OsYh��ث֨8�f�pQ�D= -{�W����#ƸT9�l5/��[�3HfAaM%ı�q����+I��4���j��Юʧ�i�u�sGG�޲ZdQ�%;XAd���T�tn�K����L.��A��9���

e�|k�U2s0@Ӊ=�� �@�j+�ڶB���@1@���~��jω�L�*�Eh���&f�a��XJ���ٮ�k �2[@Ψa*�w�L�[���'��Q 4�W�P��2�OV��}��r�%��	���]3$�T�x+V�0�c��Y&N �.$�^��i�.1aKw��:
x�L��(� 5K�B�ԟ�B�(XwD"�U	_*7�Ɉ�䝲��x�F1�f����ƀ���N׍���wψs.E�Z���@)F\d?��m�VYx"4��P�A�/o��i�wЉ�i�}������>�l����a1o��ȧ�X,�&��/e]2�2G���G���I%]����F��&[轰�0t/����|������#����]]!��6�eei?\X�q�㒹���W阓1x��Z1͎Nd�"�A</��M�Sܥ*�O�=��C&��4��A�C���ź0_&
��o6%�$�tN�������ɔ}��l>2w�N�-��dE�K&kM�0��{6F�uW��W{_k��AB�����(g���?I�:5z����E��'�+��aw�y���4ݐ�;���3J�%4�d�w5����'�`��ӧ��}���gؖ�e�Z[ޅ�K��<��
��k���[�e�r�����sa����O����S:�\�c~���7�_:��vt�8���u�E�E�����;W�#�\F�xu��|�@-�����f�]ƛy�{;�E>���է�2