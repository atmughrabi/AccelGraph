// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:45 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aS4psQF9GlQcNzViuRBuNkthI51ExrQKvhUAjEFI6px0XXOYWOKblSnD7+gSTNq2
Z7nW4wuf8UW/hg3rQxcKMqw1BTPbz4Nstlg1NZlOoD4rnDbzsUVb+HMuxmT3fuB8
yyUzZolGIBZ8jf83Kutd0PgiIm7IRGHhI4tNLlieXF0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46800)
hoyNFf5VwM88FfTRzfojUVCf7DQGYD1vvtkugQA3bItbQO8Tw9nL8CYoEKadFMNk
WT/pKK0uAJAHs+RPU6+OMV0ABIiZtcXDVI17xy8qITHAAwR6RHg4p5agem4xKVxY
uFIzkbJiNetaFGACmcZXrszSxtSTK9aWpEnyhpWpqahQPqs0Kgqm7fKJot2uDxhp
a8L6ZDLKLs2GVa4p7zKqvBnh6CHvErc7wJPpqv8xJ7jmlhOiL2PuKmzcuOlNRwJD
p4f5TYVFa1dwUilcGIgUTg2Ot2zI50UXejL3uBEtANcRd1BTGXkndNHJnXf0NBuf
lLsPOBQXzC49Dqf7a2zynP/e22KZPP35l80cLB0DXY8XxoXjneLUkKYhuj75ndnv
f2Mlr7Xi3EC44nZZcnYrhQg/PIX3gHd5GRBf5cfEjjiiZaKrwaNPS4S9puoGsYC6
WgRbzXEjfJWerWYhLvkRV8ZuPJI3twbDZq6xxKsRqp3SsP9Krl9X74JTgLrxtxMS
6yf/hmLPVducIyXcwESgHOboJxmtYIqE7RwGDjo2Qussh5/2RnbrfhkHxhxQRefo
8kNU+vCdf64EyhcywxF4+c0B9mPigiE0bbYoRmnaw005mXwd7y0U6glwWjceBgsX
g+X/wl1TOazH3VujZt9C1yIsmjQ+bvmSjaflONCZkkG0yXOPeXzdY8whr5Ngfo7Y
4SbrDsTkIpYZFS4aDP64UbgjMVNdDUejUHe8u+SWtrm5FXJdiGMNeuIzd96Iz495
KBjKj1vyLWYh7Sf3lqxrRwciM5xM5FZ21RuCkkTG4uDinbQTyIRZuHw66hhud5CJ
fCBEMAef94pDa0gMW8bPaBfEgKjv1//2gRyhu3FD7TeeK4QVhw6jekdg4sQPIVGy
vP3wQjB5VTtSBgy9NC4DBlbqJF5e/Fzqib8ITVHNxQJDw+1bqZq28geMx30BgvsP
TEzIv7YyMJEDw08v0JhCYkAtci1vg51bLBxQoDNd+OqyVrMq+uqV61ZfK4l/Z9jn
7fJ08MDxA5R0AklIguF3l0nXSbAiBDzmVhe1SAGaqfbBLFylM2tvEjVW7YdM9k7c
x480sUqcM1K/Zi25DEwWgqO+MlSVwfhydUaXto4/uFN/X4lpuUtzxiIUan4Ibvgt
1c+PG3HbrDLm9ZHKJzz0hDB75wEW603nkQScmg82Z2n+D32m2IblY0DS7PEf086q
XO92mYs3xAiQ7O2gDZXF0pnNVrCp4bQyWDtdKANOjJY5Sen9+Ec0ccGkZo6V1Tyk
Ch60cRVJAeXP6IxxNb5hezsb8C5Cy4fkEOtO0MTzYlvt37ZaHsMFC2PIC57qrp/9
mJi2DXss3BszJXg5lu7KLk0e6zI320WB7OB0HxpJLGCRYjlydC9wZIlRvLEpNuFt
bkNLlbWLjlQ41YcxiWctIwyVLDog05XlXk6a9kbK3EhWdgTrHg4Phm20umbw7mw9
dFVP1r62HujK8PVMy5sxFJ5GdaZO9Fmg6xQn879v5nUjX3Ky/oIL3o0B1xtHsDZ7
IOKz5WbIGmoqEsD/HDPj1PVyDbgXjjMd3LvuVw/XYTcsSGxzwx1q5mLa5eSW3NLU
KUqxd/y4gvaWjp70L0vaM85y2IdeQb0ysl0kIPfPsCCbU6uiWPWt1QdaeNRC9DIe
0HA4kU3dqswPDv90hHEd4OyeQ9lTvgWFEaLWuOuTGQCdKNPYBaT/E+DpHrcQ+61D
Nzy8j2AoEb+S677NnXX8fXEQ6pOqWy5AUKGMr4FUTRm/uPumxWmY0re1r3gifDQh
N/+Mywjys+7ScVSAITbscvv9vKNdVTU5ugk8w6SRv7T7knoQt4Mmol72kZr1ygN3
c7YrGqoNivDYxuLChUV98j3pUrIfMfyMN7DaxzIrHoZpe+kTMNU8T1hi6GOgldCx
v1Ke4P4w442GxcUEDtjJVua21/MREuoYHGTQhnFFMmlja+FHovxn9Na39Z3kFaTl
FI2y62BkQeQnA+9wHyR5rwd1CekQbQ2bFE+H+nraDX4yUZjo30hwtzTdDjCfG9Vj
43WaCERSY6mLqkT8N/ngsc62oWROx40mm2GYn3GMD8sbO2/N1ExweJy6ucjIRsDT
4qnA/Vi7lkQDwNf5DHSrMabFBWrgJFAX2iGE0YLbpOeeyftgXE3FnIvCBqMjpyKO
1de6dUL3gK+6RMdzH0V3QLrH3SaX8q1BWAq2mbzzq7KRmar1mbd0W658ClxsmyjX
OAoPDDDYB90N64F6b03jNxmp+MwbUg3AU0EYDtf0h0Zt7xi+dssL56N99T6bOtET
xxVzYQ+XUaZHogKPx/1n75X62RhAGtidvZfUmdUwp1KTxFFQVH/kaoaCo1HbmWGF
O5hR+yS/zOPc8iKmSq9v+FsLcpu9K8cg1NndlQeqrTjLT/2w2NnUin0As5zXIP/J
CC4ESYqH2t/0gxlGt4O23k6wb1eyo1kCQMLOatpFeO9P3UTijmWDXwY+30dl2i9D
alHSo0f30zZErz63bWOsX/L8CXF2vCG1OJEX4fCmzgSmuFFp51iE3bgzQ/w70Eqg
OkWJ8fOj9gjgS6jandoF5ivTzgTxlWF/Majtga1rED7rweiu8ckS/EA8DG1tQzR6
K3pbDX+tvVzk1QNjPzs4oOaSAAd2sn6iUSU5JloOIHBDfGmVaHMX2vVZ2qDr6YsK
RMbitnWj11yLRumWQnaysw8EjvRoD5cDTX4rymlws3ls48fFZATpgXy2c2JcAnxC
SC/KnNRg5JZs0q1hxOxZN3agBIPam58ic9WrRBEiLl0g80KRBht5Q/XXTFTubLmX
8g51I3+7vAVB8gFvNDmQMC1xs7xFxp0YTGbBmWYDbbaPj/vMbfy+bSEAJd+VPbu/
cHcPNAZMnTry7IG6YoAuBPLF9bXcOKtcSMjSGKMeJlz+yAYl7rv/s+qOWAwNlNrD
2+3q3AlJU0nV91fKniYy6Br7D4JS3xy/Mezkalj5XRJ55MycWhMavzoBcSs7W+j3
HjmQic9VCbCzttjhIZfKJUuCZCAH7PiHAsEYsXbOZ7P+axXmvxPHbvBEOQraRJkH
WNSimEtSZg6MmCDa8cRXHG/8KdvYtYC/usf6jyimUh6tPMPo+4I2+aA0yJJ1mZr8
AeneuLMMWn1ohwI8W2+NWkzdUBgDZjmymYtKmdvI+uYp1JcCv0qvmdmy4ab3fN0n
IZoQ/isUW0LjpZDfg1yuZmvH4nD4MpgYo0y3gRhtvOshW85mn7NRsgz6lqH/MX8l
ONv+IF/x9lFr+r9TcJsAqqvm9zqVqBEh6T/ofNkNKw0FbSz+WMM5DclwzedDikdd
fAV+7NR6aAmubD1EKzwFc9oiXNVBUUyzrsg9bWJni6Z1HA3cW34y9ptOwlE7aKIg
7SVtLz4Czdbdkh5XzBzeiLfehNXa0QGxLiaT0pNcWsh77Th0KyJNrxWPBGNonLam
f3nKrm8KxyBG90Cy0KJc2Juyf2UBEV47dZXXQw/k9VJMIz9TBlQGT9pCkhwWf/L+
6i4F8m4ALr30GPocsR/jt6/dqkxLaUZIyPeKp50ylFqumUolpMdPvWykI94COCNW
RAhlMgAlDqe+9sQHaheccjp5MD86m6G5bgyFGfzOfSvi8/McDr0+zGemhLDy+lb5
mrT9oiho45LQkLWGtO5aeroc1K02Ukp1dL+v7q5zp2ByeGqQW1I2m6y9OV3wF8iY
PT8pQMiOemQHYSt8wLT5qeIgf9jGomd1MQhaDtYTrXXT6pNTqNIcqLycrF5xLFK8
nnujuy0r6WrpzkNAVSYRYR77tA2kvIAnX0p46nTq/DH1/hzdJgIKt3NzyzCy1MeI
VC348Xn7LVqW+l8nP0fQ8+mqksB0tTXL0UNro2f3XZIF0K//NVP6fetym1aXXh10
U8cwu0UvIW2z7pW22oqzP0NFRy6N12gQ55r41V4Itce62dOdqfImcStMvPYgp0/Q
PjtJdLRg8FPhpLdc49L+cb/BQlnXS4yhm64ROojdkOHSXs9B/MxaveYGzBpkCSux
OuDoVRjvQyxYhKYsj2ATHabDL0apLC+KgiR+n/0KW43+vgCxku3a4M36z12j38GK
Luc3Nq+udZo0drUtmD9xjIn1AQxLlm+LUEio9MykkkQdy7w48sw6gw01eR575Skt
Bf1/KrUVFqk18p8gPZf9jRO+JgbqgE4DC+s3FYC5a3t8NBBVlkDhY47hJ95WSLST
uxWS9zqw6zCGa5Q0GN20oGaxPAzQ3VZuDWngSdyuPdn7ALGRWHfgmSik45kT0VJL
qpWSr1Qgy3jrtLFogpejTpVRXdlmLSacugyJ25mpQlLVuqZF+9gxTzZT4n5f9qFF
CpvUZ2ENgKrizVx5ssGiAL1VufGAXYlOmDFVr9P/0gkMDnBAZe6BtDgMx756pV/8
mWc0QwMlYbLygJUchejET8V9tiesfJzzCQL3FL3jtFIL7h5udWIHA4RdPeabEVLE
EtcdBGLiUvjixWxN5v+DrtkG+AlOUltla+AfBA/OMJGwFFjAN8anKWk+Rcy8rAX0
C3Ne8t20ImYn0KX4iPmObR4t2GtMR6kVzMejgSaeUfo3sk7gKPszOVe1QpyuJAX3
f6hYqkT+ROL5aVOu9qP8+Y4pyw0peRwthkeoPb8bU9MAFehP5dLjJBFlXarVB5+8
K253TNyYs33ZICHu8TOnIVCuNBR2kGEEevsXvEdbSOp8fOQxrs3c5IVy7rPbaBrL
0P7t+C4awb37pHoDarn34YYAMzOfT+CySU0RusuNCYktD48xwgjEL1lDVH27WUIe
sGylKafedYp15ieM3WUnd3/GpeDGMAx3Yw61xX6nKOMTsadtaDkLdahxXzqvVHCE
yZmuBIyNJu7v1bSXMHh0555xI22K4TskTRSnhxitCZL4jPEMBE0CHOCXW458F3uJ
4Be/+r5vdsxhYP0pQSP/FPqnanoDnbcmTeo9qxyFoQ/kfp8kPK0Qeqwp3ITcPGe9
qmAE6YXsE/+DcF1czEc8xVobAMH0QWZANwoZ0nzfpW2mXXjBHBik6wa2DG5LDf93
2nle5ppIWuYyyhqsE1Q9CtXBwzhqQIFH3EMUB6bDvZFBoz2XKohzJwXlx8iGKEhc
DR0ll9XCgJe5br9S4WfhZnVCYZbfgqUSiLEwEyIvmnqjj60h4NZHmhOyryaD95N0
abTLi++dHOBQvAYbKhh03Tds75JXD7GdZy+6u42tsMaEd/TZ1qITrSSkjAFjgaDp
/VSgnxYmX/qYLazgoeQRC1ZzJOUEcA+Xf/6ZUzeWjDMHffuHUTd7OqL9gEiugufm
oQ5ozDDBpixfLyZ+LgfPAZk7FsyxqNKOy0qOkfb9foRKxJhMOB5yVk5lRhx8mx7M
eXqI++b9BdAAuAXxla3B8SsAywkfll9NxtTpMvukza9yyd7hGZZUdllEH3pez4Kj
bojPEm77ZITfJf3xUWHiA4lV9oehQGy1ZSTEPQsl5ye2TbskDBeIo837nwNWAh8k
7poy/TckXtPwv7LOB7Ovj4vxhgssbh1vALNbez66CTEHYX3u4EQtDep00qRQkm3e
Cos5qUKvK0vDXpdBuhzrF/+fhGwKfQWt7SoLlYbuYIS3LkeUydwEE+NiOuzBf921
zrs8MwSczjF6Hv/uJnPVHyDH2JGxDtBPlL1uUalHvOx30TQ0fM/m8OuF+/aokvGn
4ieO9YDJ49leeUFDmWVh0cnZasFWrzKoO/NEq1+lmcQjJqCQOyd6yeesS1QKDS0r
/RybFaGUbUkEJVaFeWECr0BDykrN8ALczIhXEFowO5ub3t9wyDv1BjBt7BmpV9r1
JiYj9ZA3u7g3PkoJepI3HCNHg6zysxdm0PIIl15W177IvJiYCnLz5LzTQnSOLPKZ
zab8Hhy1ACIeqSohXjjAEj3rhs6FegDMRdRGpsn8kD8N3gUPzYl5rXgKn+IEoPMB
3sGTb7WlBOavyabT5y4kZA0m/offPJFj3k8q+UpJOrPyRjbVWnHZPQWLyprCBPql
ry0P5dX87yQToatuo1pUF5zjpXB7KPuQCrN2ZJGbJk/xjGwz9Nz24n1qxs/Ma0nb
5WtqKz+aRBS94acmlDWV5Loa68klSRmXvWZSZuq4yPSkr5RyxusOZ07z2axjT5Tv
FM5JE0ZZKiu015Q+9ADZa+rMjdH72n15qEh0Ra95r62/TAycr6Z2/ipPfG3GIFXQ
ctCVwqYbftS595ZVvCdov3Kc+diPvcKc19/B9ZB5CFGRQkhKHfAv7pVDg0h0N7Nc
/h6qJHk5BTdyNxGMEP5EJsPyqMHIVaU486URHxnJA8bA2PYgl4wLeNQZYa4wy4ub
MvxORdd+ngT2NVNCRzsqEhhtAw3aLbjSFhrqlKHvcipptyQzu2WkkJbpuev2c26e
CY4ZeMgbR9uU3NPiP7Y8kRhNrhC0OJdXv34ZGVBoeFBYs2Lxu8o0FjMsR9tXBmaT
6yeJdeYeRvHA2cX9N0ykIppcXhe2NH96shg8fIYJsNes/TlxrhBJG3zBDKhbd1FI
tGyXzfO+bSBsuBLNXDJ1cN9uEh6/UCe6rsp8rv1gnHvPpX4IcWf2XTxacmjmrKWQ
+9KlVILu+zmmqlO8IDa2hj/XTgHAqWWVudPOzlS1kgb5azVkpnCQNoEfp3EcU6Aw
Z5MLXpGAAK3C5A1tqyTGxu+XJ+hwAX44q4xBbbQx07njetPqxnH+wmSRqigGvTdg
G2/hv9kVnjfgtk+tkjw/aBZLD+uv1meAs5DB9wNbcX07M/CGXozRIUmoz0TylIir
UQ8OwchQv8j4K+lPE9LIfVNDiOLlOPtRlhmEcehxFPSRriYzqh4VkPBUZFkaqvmd
B0uTi3byutWrmRv7/OeGFPToHprfx+wIxEVs9MvAcwOfBTL5Bnfoi8GFYTrGW3tP
RSRqHCUnOT4XjDTcCDUBXFKVpbmzwc8C1ljQr8vYtiTNj0YNLLd1YxEM03m6v2+i
KIiMwsN0ed+EHXMTH52ZFzSikeTTC1qCi20LhwMObzdCl66JvGRcJNT5yNdQ2byd
P7zdHSLgPLbLkwMrj3EGjmcFWxQo5vYK3j6Q12RmxRL7xbTIFSM3A/c8xC62Uv3y
TKYAxx6GzsRdQrFswO+RliuDTYNaaOrsmW4BpkKOTjrqte1skHLcAQzoVyAU8UbZ
7hezmp03weDlN/vPKjxci7CEfTFGZ7pOy+6/M3Gy3c+PUEopQomf0vTtSRMrFfOo
J4ELuSmr0yfaLZM3gdIk/WofOpR9WtAzXNXPh+jUqWzcaqRjpt2jjLrBWDCoJE+x
ObxTBIhwgoJKlXv3+S8gz+rP6vh5PF+z15i/HH+utwZgAd/m6c90fbkZmJphizkN
zox37+UacfWrmTdR9OGSfEAw/eHp5YjFWY2LiOLzBJ87VyLADo84RXvzS2GvHzRd
E8zR/hw40y9nFLzOlVeJ/zs1gyeFXkkO6c8oB6QvgIL87aSqfavaHigq7kJYY281
tXDDaSewiSKv9nTn9rmviLm4zt/PIgpNbxxdXH3MTpU26U3VhJ/mry1U20WJKin2
xbujawRQYfMjyzDXhgd2vBmb9Em7NuJi6LYL0XxZGrRt3oFLdEvI0mcirVYP2Tlx
cdyVzCBw5oaJVQS8tC5L4UM7o5Po8d00VJ5+IxLRpUUQfv4FR61DFdlaxjE+eZAy
QBxFWzTOZaJjvQ31m1SqJp69iLzpUDYlH6UYwdeEi8hsF8Yl6UVFosAryhDWI3eZ
YVM6teVNdVxLfoBbrJaSWJaowu7rQswjzjZnGnYjctEjiqTkIoxzdELt9RLC4Oym
myxqkdCWSI7A0IyIESuiWBB75l0kIpoC1ogYk8kdNoENHj9SYB4gKHPXaUi/gNGR
P5tQl974C5ymn+FcJV8mdEyL+wOQfcSYF6SbnSUEgFol/TqjdzM2m6vOF5gVE0k/
+kQgteb2mwTxeg74R93qlhShy06mOSi8BbeB+JpznXXq7k/RYsZBT7sSkyWI1RhT
f6KlV0QX2RRLg8zm7Nl95ZiMYGBP8KVWNfvkRnG8etrQtPtpiAFKIGlidyr6trBu
S86FG5BGbHCmzEN/EE5g5wWTh9Yym3Tuy9EISywAlJOMjhUIHB0l/BELVPY2L7GN
sC9saRVywE3X06/5naJzx2OxuNzfxF5jeUd3HFpeGYH2lSNQCqGtKhQbAdR/KDUU
zA8O8Ph42gfn/gGmCEux2s/Ob7vqWdOCtax1M1IVVIu5mqToyoJjpKMcQUxbU9Cx
lkKlFrPAa1lGatHT0MqKkrdjL8QrqYHZNz9mhb221zehueSZYQutuEfubYZusKg7
vJcE2Skc9E4qAJ7rHgl55M95RDgQYq5WOXmoi9T3uxGdfEsgW4fy8YWHDIyMdxhh
sOUYRk4gMX7NqcltGiYo6plPypsl7jxH3BfNJ4IADJHjCuXsSWYkvKMRC6K30dFM
CVNq5jYeZhSdurJRf3kCiB2Cohh0zzKjPMvJJHClST817kuJVfYnTiBOfb4RScX0
+7M9oV1kuqTsxJiiQBqteVZKycKIVJ0TE2m45RVqLI+0G4ET8ofqsfocu5PGGZNA
dm6TZQqS7lhwvFJ73u6ZxEvk97rZMRYC+x6oR0GTMKLIEWDLGkKBK08kVUAuRklE
igKcv4BXu/MaBDPk99KPUGADct8fMORsBff8yBOk2JLUj4Wl2S5X9aUc7QecBJpL
p0MqFluFdxOuUIp4vK+8HG2Vgf9b3q5b1dLiSJeacvJwW4m1sxxoIHARav1SCPEG
19JVRT0J15S9IFHvLp6WCbavfR+VKDHH8Z7hC9aNeQsxK9X+Q9yFTcyi4mHXwu9t
pNEMygzKA2aytg0tRch9WUhRo/tMbaboyN6gV5kJaJYTrCXR6a6WNk22uPEqyMh9
SdLI6Ftj4F3ZzZPpI1ObOHtiFIVa4UQQ00tpM0lDhFCbcAeGBSnoiKT89itqvTaI
K3C/MTGp+OY8ZKp11r3tZFV+4e837xqXqdHJPTa2Ax1BuKgcijn2tkmcir/gu0WX
tis347+r8NF7nLMjn9eBpbMCRnkqeG2u6uyTx/AvspnRwgzJ3VhjmaH9ILc+GxK4
xGBe2iswULNB8bnk0Z9Tzr4SgbeercQ1QVmz3IjXe+IYuHzvtkmrKnhq3ctIr9+S
6VeqCiJN36uR+PQ2WI9GFQIU5N7EofrXQHweoc+laSYPlBV7XezbtBgqxTxwOSQO
aMjasv8Ls0FqWg6GUd98RQXttFEi9V36S+PnvltsiyuuZfN0Mdef32c8CG9ceaea
9qj72AWxQC3oFPKRXLUeOo+HczP2BZ5x1xppLl6+0kAbUa61Jp5xPOhy/e0dfy+E
/ygRGt1KgOTaWs+xK8ZzkmFoFT3rUHlRYi0SED1Gkd7TNp5+LLp6Hw4B+/y4wmcC
833zdA9DMd+Wc2ixXo5rhwaU4A1BEjfrSzPRjKOKJXcOx6Y/DWs4eHZcxElE0N2E
38MKYSSH0vEHgHDvnjFL3mlp4BSKhLFj87K4+UBBj7CnPT7JtQc1TBwAagHohvhN
BhdB1o+ZUZ7kTLt8jaym8hPTw8FnYx8abQN+/sr9wlVI1Hv0ZeZNc6MS0W4W6FRG
LPY/3Ufsmc1E6TDQFWk60bcEjimi4F8IUQ+WGdo+B+3HkienFSJQt6vSl1og4xik
xDhIbJQv0/8uSkem1n/2xI6gih60I2o73lfv53lFSacrHsZX1A2aiJGcnwUYEYFs
y2GyEinC04hIV/kUo8FXrHfYezDqyisyFwR5T9/2Z7gvfFwGZoSdqDmNShmDOHvc
wYhX0Byd6XOCapgBwxw4EvDa3kI1xFy4aWYzwbR01YT0VC9UaWBICAtqcVQ8LkdS
BP1pyxP8JltnPUqMLLf1sO8Ne/duU9K0AQdUqS08quaHbwhLML7uiA677r9F/XGK
iKd5vOmgjxFXTQf27Q+y2bxnKyugoH0x33I1nJ9YgA21DNFrxlUf+9rxAaX6SMYP
6QCbN27V4rwc7cMkct/qFV1H5Dnl4M3BTLfUvestavWmzy48sVtFWzFg1IpbNuGV
QVqLA5mG61IuA2DLG6wqww8DhbKtir52XudP1VeEjIW/erGn/ACHCpURgqCdOk+g
xGEdl2X0HV1ld1Lg0ZfBak63Uwetr7C68MbGDRp5PsujJT7N7A3Y4ytwSEEn5+Z+
qHMbYtQuPTRDMJBfii2ARJ7Bw0pMKqXDMN7zMgIRnXITtsDF0HHfu/Timm7qJPHs
+6XkP1On2pEuKIVGCcyZBocXdLDSta1+hJgiC5PnfRqBtyyBQMrBXIX5Mtc8YsHs
3k4SLQJcXSsIR9waCgfXiqHzLT9T3PTyiE/z7nDKwTrS3v6jbe0occ+wMtO92VFY
uzAAYeHVLWCAtQD6xqzyu5yGiY2jABSBoZmu4hmPCqaKhQIg7sfzUgw49qKPZDXO
B0AmuKBM4V5AVsrPNSscwOl04OuKBgTDNRw4YZAu1ejxB4CJu4chUeh0PaHY5AV8
mIV1DsOHaBV1r1V7G+DHDEcE/cAGxhnYtU78CqkqP5FTOYYjG2Sb4C4ntOhEDcyP
E/tDizrJ94JgsMQ5M0nYdiDRyVfxf3kxQOtnHFOsIjdix5aNMh+LczV4VGsmDLfw
vJ7/bXdhsyY12vJhq9fJ801Dgai0jWF0MSKIwWw4O/jhlljKzH1ziXcsy+rYdw/T
xDadq5EAYvxaLaqZnUR/GxPnWt9U6Q8MwCqDJJHrLvP6CW5Y9gM4YbK+SXvJTR6s
d7BPKufjmSh41OebUP8KTdClaNFHR7m9ILY3nQ4NUCX6TFiFjjnSAa+XNsV4d/XW
pwAZu1Us4ZsZX7qLIwAu169VXVtZTsPH/dfGChg9DM77I3RVdo9NrtyPuJdwOA0V
JuW7Nz5d4We6bPWz6J4xblvP3xCHVjVvf/umlMS3qTQzqVSlX4KJ29MFhRzb70D1
Z7B25pvg5CTr4YRR7D8Of0fv382HK+PAHxwzkXP2F5SrTvrwRjVJ56vhRSAi0s/P
df8OKW8mJcPpMx55hLDJbUSoB8WBv/gVI3D2zs6ogyDpc+47C2YTyrOFvdg7o2OF
5D+5/VXxuftLQbIDaxsYgw7DkFrSzpEy9wl5WYYT/VHVEtVhAZ0QIrA1OxhzhPTc
eiGrmKM/CBzXgqFGmu+uc9SKDrCagKHPGXId9lErLxcPYTV+WAHpzYFhVY+D6AF/
fNpuoLPz9KbQRfD/++8W3UQ26/ambitew50FpaChrxNQ736fYJTyM0AnGwzy8B/1
ZG/lSUTtL6lZ8676GD9GQLEefOXZhL+zlRtyrcGMqq5T4EcECut7qXJK1un786K7
WXPHFLEGnN/fVtI376B8FL406Q4mxklzMqSfqT2s4opj5OrL1GB+OdijPBCawzsC
xDT7b1nXpr+QEfl/Ji5Ehu3UhBP7e3EItmNJZ1Tq0DBy2p8GUJDpNkOs4m4SbCXK
1EsLiXR/9OKt3oyOUI24se+cyJMHhmUOcA1Gr+ksYtbM8DpPDeM4SIktF7YzFZgQ
eAWgLXX8DtuZ0vUF8J5yJvjgNbVCGFI4NIk3kpItBa55cdx8W2ZZFtn0gmxxd5Xk
vHeu5UXv+PDGNpi3Poag8F4TJaLzvlsW9ob0LxXIT8vFDURLZya0qYqFIeHA283S
n6OVxN/ybwBOOr4TkQqPWz1o28Wqbq237bP+7VVVwrkZck80UP32JKd7zT5xOyRh
REeeyic5iUKdEwwFXSW/v5rQ+a0gwR12WLh2QmI4ANKDluAdvcL4p3yJxtA0GPry
c429nt7ngCQcEMscGwM2k0FQsJmSKqGGWMcvIl9HiwfKTkStuYOfgIa4r+hLyXJK
WZfrHZA1+7c9koARl+oZeJ1/hCTMjzwLeHlIIA0rll0KW/9QjJTr5NklAS8P19k6
7a4tStbKCs8cbFwydJviezPBaUyZ3dFapnM/0ThkoLiSe5e4+fUV1egK88Yp2+vM
GUEMRzMa4lgcNEopvL25vAH7Pe4E2lRRGTC+ERUTA0uGcsG3dsrOCW0UbZxE7NEY
SIqFwjXyIuKFdNV9CSPGzKbKrwfLu32B88/fNX8QC+qxusqjPr24RnaT+Xmq2ht5
bSVskkJusC/G3HqPOa2KVxgMTB0We6X7pzKnNM5SWMKvCkeAloFsGjad9G795A29
dGvuxLA3pv6x25ADWMM4ZCnrLE7EW9EIsME4ezGSDWsWAOxpLEQDlpU2ehgHlp6r
WhuLek9VpvfHDOY9+7kT4ayH/cdS9k0cFc7jvAXyTEePR4zcFXo9Gf94h8yawChb
UzKBwr5AV3hX62uSz+TtxTdv2/PTP2nHBw4pELf9cM0vrThCyD8prLwHYHKrXt5b
q7XN5EcwiVsy4bVk1+LrWm9QtXKnVXfXcOBNFB6d+9t3Lxlul4zvTGZ2xK4bS729
d/C6cvkVqAztN+5NXH+3uVIIx5YY1dpErNMm2dhfoGOLcKDIj7o8lmJ9Pv0LZdwH
ZPIcotYI/Oi0S/K/p5M6DHgdgv6KWDZcceJBGVpCX+LMgOy8YenGWjb0AKgTk7vl
ZmZNkBvm4VLTSRMARQKsdwdxcjMoHiQDsge8jT7YsM3Z+BndToBSAJb15RMmbwUC
BOhAq6T6L7cxOvd6rTn6gFc7XIyNFm4yzbDBfVEEfd3Wikf6rkc16mZRdYRGTHNK
MNwKM4xlF7CRdjvd4J3s52VDU1G26wWC7uAmvw7gpTnDg6zymptIK9bvzILSRU+T
IzT1wKaBaZKAwnpA+uZl3uHrFva7eQIpIU5QJ27oSVDv/c2RsKjCi7NpEVT84Z0F
XPmvaO2Og+ipNxQ96tle/ZQD1hXB3iLHHtdrPrI3ZDwEd3ldNKiX2o7Sacm+EP8v
edUuteUKrDZcRAIFg0BmRD0C32YU5wNWuNJIrSMdDynu2tCu6CjB4/p4S4sLkuLy
nnFu0+RO1F41Q9A82PeHu0kBfKjxBMruDsv+2C3kCAi2WgdQutz+Zks4vgxKu/Qk
fqymQlDVYAJccTEdvyVF6RpSuIPbboj1mETOzzxGU8tiXVjPANT/GtWf8pYqlBsO
s6/+KXMMQVg+FQRf4o/Y5by0FkyZd5apsA1lFMy7fK9zEqAPDIUe264FQAyveBfb
SgbfEUJFHmsoMTq7P4W6kyJIQ3/tCr3YQ7CjSNUn1QzDo+OD9eb6U5XbmT+grFo/
bwf8Z1hl4JOITVkLAqnDbGncOzg4Hl5bOwJpKuVDQs8DOD3Zrd3OIdOe9rpXb1RV
Pe4SshDgUBlV9tukUFA97Zye8sSNWuFg5DSPYqhZwwHq6d125dqlRE0uv9NmEOuj
83Aqi5PRJxewK5Ms0BIK/4Dwz0CUnKGr997/HGpClMibhPpRX3osSfnVzMYAa7On
UpHlSuhwXBInVOP39LFW11XQ+ej0QykBBdnAXeTYPMYz1yp2o57eqnL11529d3tO
mbKqG7cNx6gEeevtXV8wnIzioc8P/hDv6LsPLpIec7NpFrUVKvWCAEvYoZN6s0CC
sl1+ZuVjv9SwPqxjmxJu0t4P/6ckXNJzUCRc10egdAVxdf1Q8vAXtmpX0uqgcZM6
AKof+XRdcj+wC797VmLrA4GpvzA3ld+uxg+S0rj+xI2sQTEKnec7Bxp9b1jvGdpG
KOIhWnG45CPNEHHcQTg+J7g113rxW2gr6u67dPvL/UkJHAP49183TzKVc4IQrTtR
R+yINFNaSCmitSTNw/rUtSIwUKl12tr5urD+lWjmElOVwbiPkcfrjyY3S82jHwzC
i1Ozl0SbPFjkKNbHMgccNQu3yAaY6zsOwg/6XXBFv6dV54c1VnQVUT6P5xqr5WDg
zyUt/E8URuN8oXbHw0a6OxIMLDjFDFxAwpY+iDmV6qKf7xmMRRo7hXE4CqNEYsXW
uUWdHfK94EQEjZmA1Yyhx2O0Ss6AqcDlggwgoZzTSwZjV57ilveTOd6wezlLT8XW
T7jjN/xZ8XCLqdW+U2f0lYXAuQZ1rRswZn9rAnuhDrfIMai8XlWD7R5Ri/l7QZfa
ueP6rCsZDVG7hPUtiT6Keaf3/Kaj6NINbRiWpewNhZNbglC2joCgP5wsbO9/oGPF
HLxDmCSzSG9g+AK3/vyObiERkYRplDIy7/Qfa38+41wwoMGsZzpKXFvA66ojl0eo
LH3gVbfmwW6tYXtx3yXQ0IUas2HoOLbD+r/U8vZHdn1R36nJbNK4mjw4b82b7gyT
p5oiS5IZ+QFSLo7yhSTU+ZXInn1FHKIk/Y5jz1OiyNYbpir29UrQSpCmyrkIFnfv
E4jNNv0fexlua/GjInGN/K9cQPXdvVLVDJt4jWr8MTzcXoYqVE+KJ+YXteFGs8dE
/XDexJfT/mGJTMd/W1RtdYqswzLixy42incOtebq+K+0R/6pab9Fv+fpV3PYHKJB
b4JdNghJA7c7J77BSWx4MFEKUcz0lUSQkNa1xgJMBc42XhGGn5nzJNcZmXkytBeB
CsJJLvnKKvSpyyAcme0y7mSreJ4pZEczAzUrrbjAjm6fLwTj68sjXfkimH21tWKN
GY9Aut+iPcsemV9QYpYna+6BkR9Kvcl649qjSPQJKaLj8eUiE7poUbSbT7qW4tEe
PL6cpX2/Q/sdISJCcuVb8KAaG5WcHYzPfteTVUnL9tSogkogOXdHkMBbXoX8FxTR
guP2AColi0pWDxhGxYOHf61XAFX+4nPRIzsSWl+kOu3r3CEK96NfdJz36mrWadTq
J9xwMJUIAIi40+FTCA2tp8WgI1tmJNb2QruR/pcYNleJkjFpJNHMFOnsoTTv90K+
VUsBUuOFE1+aClkfoV4Sgdxe/ygvQ/iuHtmOsq0eezazVUXuRDBkQXJ8jNlo9lLQ
7ospWv/O71gNHxhlupr2vO/h8/EdzTuMYLQTDHQVLeAbnooBex+Z+DUcFMsmkceE
j7pHvljt/ydbIZcgFBGSICYPCeVh82xdbetVUh0k3xriVrP+XNIK/F4vufCgFu3r
jCe1B7VzTUbHkXwkYzNEvkbet91Qqcp5N6H/9pME4d+QeQr9VXfVtLIegWjnf925
SglGt6ev75/4Dp2IZddSknVXYwIsYddyj1pNTmt4CViozzEhQawNBKQSgQeDyoGH
NVExB/LLH42QKlaPs/7bUKelj2d8MTy/RRHF2Jlgi/ABBr2ApDn+Ybt9kKN9kQ1e
uA2UDIv937I+Ce6uaEN85+7DIsSpnMjun8BgA+AbPeiaRiqLLsPWrOjE1mhzlzZu
cyEzRpE3E6HGPxiymnJGuvws7ua4/YSHKtNwmbt1dr7aPQ7b5GU4m+09IDvZVKwN
tzGx1fxaa0YIfS1+6n4YQA6s1i6TTK0mRGw2E/V+mhW1V6KmE2AoGQPgU60+40/g
liavotXC75GrIFlXeF3cxkKMVhR3gcfhC8R1SIVdpE5ntMXSp5c8zkZ5Kf5RZWUH
RB318QMpkQz6XR1sg8CpZ34yQ7jQZaqSKZi8LGMoEtIk3U1hY0KWYtFxkKqJifsc
zwTdFNLFKmU6wlxz3w9AOk9AuvFdwiz2ZfI0Cr10sPkxWtL2pWD10r35dkFMK4o7
7RBrJTB9gIug6dXNMDZLEsXf1eoPGuOaH63jGN64OzQLco/miKbJafJNDA/dMwQr
FHyGZi9xHioelFC1PHKpqHWNOROFcOLQwcvT/4o2MBlEfM93oT72ifztphEHpwpQ
9s7Zm+pbc9XdmRD3GBJ9WgHJ81iJ711zWLhQUARrVP3PfESrU4KclNlNaCVYOONZ
h0pYUEY9Jv4ej9z+foqzf1KsP76Fnnc7CC4VfHbwCZnCJyG4+vZJDeWNvNLNOypO
2GLzbveYke76YGDN0GlwTaCV3CyS3cigSCTedxCXo/kyI/mhUxg+5KnA4ghXAyaq
R1p0j0JI6dcFuy/FdXSTWR7VbMHi8CfWpESl3zevW4rr4KppzvlHiIX7hl2uIRb3
7dZHzBYv0wYeSMDEWdiQOlZhmaoLAGsX8b8VsIhjFxpMPIUxy2PVPnTePw3BryB8
sewPCXN2vi2ivZp3PBVA6beNARn8CMQOwQea8K6urg6bw2nCDZhmS/R8Rb3yT2Cd
yF60YDWnQt4pv+eYhRx424uu37nAM6TN6HqIhl15ztwdkA6AKJhhm46iXRKQWhBp
s3AAoH37aRBaZeuVGJ2/l5hNU9mfFLvgA/hxRRX4XfsFYeXW6RYKrfYj5akWZN6+
z0IxcHRStvevOcmhop03WNxoudLY35OQoWDKsaLxt3HSCye10fep9WjRto5eJQ11
GqtAdyy9yeLBEL/ayFMv0zTuwuLcqzxP2dDtl7XAXi94lSssdYFMlDhgxhp93dp6
sQH1RfUHY68ZhSWL1u5/hlSm5S9OO8CPD4ffubC/bQ2s1YYX2OhT1ZL0jtgQBoTH
BV00KEpElnWUuJQx2PF8kntUWI7pH8ro0sZo39N4sSaKm+kKr+SmE+OByPYfXTIY
K0LaLvIRqVOqODXnjqYFdEM0LmXFLVnaaPiokPP5H/hyodJtIDQgtDAfZLKRZtOk
xXGdPRjWuN0UtV/0EqXAwWQt2DflftJizdjlWD5QaawinPcY7MkyowyLKDoSbQgD
+qrPnkToHLXV/vXIB24X9FzOB2noqqFvpQtdV32pp9DoWhSQgTH0CmcAsEY3PhVN
UPS6gP/sYIgH8NdMryHZ0U/STzQYIPypIXkXebt1udT+qeXvFaVrsLhHMYvl84dC
VE5XJX8Aw8JfIddiOz3qA5Kv0jBD/OSxw/q83uT/2s3bghixSIoNXry50z9JZJ+9
gVoPENELdDXLQ7+LZhFfHlXfKk4VkN3kqKnf3KQan0MZK/3oSqOpG0ZwjAYZZaQv
gh+H6Ndo+sx6YReiTFDQSQhGMw+Y/gcJHa0wHdwjyePqNsxrpQVZihqzlKGt5v8F
rl/xv3KL9QHHAEOxm1l2lruOEJh7YNPhZuL++bHAR4igwoFHsEAgWhL4EYZFw9Wz
jp4NI+b5kX45UZU8sxl0xCkOfPGgNBpSFPZu+y4TwfF9c4UhquHipJvAyQYtbkdP
1QPd5wESOHWRQsFVZi3rynH07roVcMuxRXQgN0T61IYndrm8jxlJddnXRgxcWUib
nkWRBtT4FgDB7UA4rt88CXEL+8T1hBZXXTQP1pLt9NWs9zSDycMYvCcMvqQaXzpK
BlpZ1bPEAkWy47S0VE92vRvsc/RGLbLZF5NDYT2MJiVaT8ThiqN9S2kvPZPJVgTn
ftdRmtpNjfi6S/pwuOOuMHvuAAl2kdYyAbWorU7wAGPWiGXLjUCWY8RoCcsj/WpP
SA1hi/6MitZmZEw90LMpRzNC582mWTx/OZ/JleZ5KkdMsGM5bGokURDGFIdlKXkI
JNsquuyEoVf+4PTaEOf+2J241cGyUa67kxwYvpQo92ViKoQb3VTxQQDWZNukQFuL
dFzzgpmX3qGEZlKSexL+QksWxoV0Nrciw8zhXLu7j29kgNj1PJOn1dfOH+6u0Xq/
zAjTK6yXMKYwWmvfWDLqU7LfXJdZFdLXI5DroZu8ucCJ3KpjsmnXMeteFaB871VW
jlgoeHOHndHOSw1LeOfhBhq6fbk+cnB9hQ/JN/gzONIzb4VF630DLNzJJWhfLcnv
SxJqv2shW34aE1mwa8XBGP+3MHepgQNA0jmTSPv7wNY0vyBtL9oOriltgnfDZ208
lx9mnRZYrwd1Wif/ZBEct5DUkGWSVUrUuJIbxrHmz9Zyhb7Fxm6JRbi1x0U+oD/8
EBhpCxg6ZAxVE2JG5A3JzM78nbrwk/QQhlbQEtgIoU54/FDabfAWQRXnTD/rJoQg
3Z34gSN8r5+Q0OsyJpXqfi7VvDeXmuuocgPZylw2+to0MItUlotLcr/J56yFosLF
P1DOFhaIOfAC0SJ8RlOEUBj/l7PcoU0JQ1VVDY1dcFTD73A1wek2wuO6SEg0jAfo
bYZmjAWPyK8Cj1v2AzHolJSM4IOwRYNt8h856FIHYJm8i1ZMQ8rWK2APY4iyqWke
f7uTUOLh3zErcd9q9FJ5rfZStbkNsWSgh96x2HzPi+BV/zzJ8ei3cLzzt9XmaL2o
N37uatnKk7i0/g5St3NSmSdlBnMoUkI0l7TSUy4VJBhGKsBFtpEUTXox25+N9xw8
PTb1i0wlhWCk7zO6Q1Y6sEfGg9yUAz/y1RF1cMRtxZyJDsp307Kch4RzQjqpajEb
nvm2f7Mjdf1kttQwxq4zuDZ8Abnppx43JoBkMZUWa0CE87Zb1Q5/zIgspB45l4sS
Od9eGCBuCIdfmUJklqb0bBrzhMF0w8I2LQ3TI7b5xpQKYulNvVMpC3V25IcKnHmi
FafJAZ9rEAes0PwsUjkK5sOvvmZ9E9cAZ1PWyIfb/KBLUUmgZg43BMy7b28hnyxz
bvI+ijBXmd3sOw8rJxef9nByULOBMqwFbb8Rmy2ThMNuV9qzP2MbT67HsSX3kvZ6
gbqX3bup6TQiOSBq9vZtAOzPA21U1F/xG4//eV6OBKgnftSaCXoZcBCFHAKFdO72
nHq/SAhwkRACWfe5IXAj35nCvCI+IG537a2BTwiKU8pj/zgS9K8dcawGMeBnXPXf
30u1r0DdthoGh8DDgya7GhZf9Vg8rP+gk2+CKIqTwU895A61eTDsoyLKuAEKvipr
T1Ff3bvl98Ds/D69UbAntFXrktXoof1pYmvBMxpGmcmfEtUEUE0BnAe/AIicsFFt
cn2JgHiGk6DVXAUVr9/yxJlhj94flY4W3QhqK1dM/oxqrE7Hv0GOfJP9ZpgsjKeV
SrlgzPdIqPKStxP1SLhEanzBEVS5FVNFoVzQj0xtAh7EmXOE2xJ3tTyatB1vLMME
JdKGY3QSKAwtJB+i8WxMivBpYT6D5ghp5XWdeT5LnnHs4ZSofspB9pWlDJDFNggO
dgaqq7azI8cSQeGkkkvFr749eB7UklXsafwl1OmyZLiK203LodCWcaBBy1Z0fseb
aGathZHMDzqv8s2QaXI0eblXnwP5RwSGiOOFSrCvXKwP0VPHA4q1e0i1PlCtqDSK
b0vX2dgyQ2GYSwWAxuUAEFnLCc40fRz7lL7hEWSHJnCXtwU/WnPauIX8XSqAqnvz
XLy3CpoXFPOCpViVIxqKArFaY8eYG30pQBlKOHXTzJ5IC//MX5WER2XMOnl0+vy4
7gZ/deUOu/5fWlSQcBjvhI59DLyt+DzfrQAe6BAodqk1hd2r6WXy3YyQdDUIHLOG
kYDCtlSxZYn7SaKUR39JCmj9zLUzyD0niOWvIECYuBwuEBAYNPqcTSKrpWqRNxfh
RqWmdtB5oDDTDUU9ej0W/8ToA36x7l0DFBFer13vrE29g2F1suWbIlOStjYSqjtv
/SgT58E+EvEqKsH7plv12dErm5sPRofdXcIHwsQ049r0kLM42UecMIRk8SIfAPjk
9WbKCw1wrL0Rm/1EP5r+3KoBEA60vfcPwaPYqkB06je80PdA69HVKIPAoWWWMXbg
xFJTEimtPje1HXKVCfG6DEY3vN5DYBS/SywZqnbAPe/6gxq+n0WX2foV4ktcuQJl
uZt72whFCO/a5D8ZB+NQRIpW3TxjSrTp4/Pbdi9/spwO8o0Dv6tbFsCy2QXbKApZ
m2RZa/AjmYEUGJAJQS0WMWRnB3UfZGAO1M2Th6tPqN8UnPx1KL/VsO8lPx5YNiA2
AdVfZ2O9C5W+iQNI8iEFwLsznxyvWvCH8kXLOtPMz35iO6wmUhFuIUzyiIoDZnK5
ytbFtMZLSKyGJuMYPuVqNdRzYIO2BlpUSmD7c+VRzxOM43AA7xd8r1T7Eh+Y/Bq+
FTNiD+AiInSzx0Kw5zuGpIZc30alDyDaaPc/hRj29Vb7SkxfZFZaXzcehoD+8rQi
4dyEnxqEBwvq4+jGDkKgrFe3RwjeE6mSeFUqwmSeApVlntI1sCJBzguL8peUSxt7
LS+fdXKRaddOe1JBSgZtDQz8wgJ1ZrGMsgVebKFaYmPFRe+6+Mk9qwTSRaDW6KWr
6sxvDMS1U819sB/Pt6ZpI9ZIdfNADmhu9Lv0A6gin7Qlin8DGcURgpLhHkCDCgeg
dOR8D/jBJ4uFdwuL+1hzmlf9qsOOZEbM8+Dqk1upN6SvsJktO3CT4tpxPbCfvC63
wB1QovEVnT4NAtAK7B6NfHmU5YBvwGzvai2VWu/zti60KmyY/wfk/jbcHkQ1gY2+
VlkJxG/Ga3FexH7Ev8ga80PfPU86EeR+HDdg5tU6SuTyyR5doq6Scl/n0TGqjmwk
4Xu0Ng2Q+9S6dl4m1fIOtVMrNo0TKNjy2mlZXxDGsz1LTlrAzpqmcqeIy93uH3+k
3mMJNCwtUDJDXhnUfrPwEKeRDG8upIhlpMxlMmaoMeHcRlqPCDSIx9yMTDP25VJC
wPq/iJvHIt397QNc1fy6Ws8N95OL0zdeN93UrzKeLiQv4JBfKXqOOQcdJTCgQkxj
qFUF8gzKclWW4zfp3kFfoJVrBFz1YKh0S6W+byDb4WkaYOgmH1ZCwUem2xWlDA6F
TyKuJVM/ZhJOUO/6P2u2bFDCSXevOPhnEuJpCgbuC5/jkTipW1834uBdsAEsKlko
VIt6XLMMrdt34GirwR/67+dTMu1ANfo/o2S6P/I0HnQ0JiNsKIEt5964VhBCca6I
CaOg7oP6j67T/YzS7fsz213aN6hRXliLQhyhcL6quvLHKKgHD5WnDhZ07JSPiE7a
2y1xf3cp+VmgwSY7KNKt/wqMPC1BCXTQRJRs4eiW8b2vdB8tX+ioBBUgL7ZuSd3X
LIphCzfHWbP92VsaUMatQ4OXF147k1oTyeFW+Yh13S0CkTceR3S9m0fYfZ36m3Gk
fVh9O6N4f+HzXc2viQrIu0TJnzjb94Et3cyMEst26QdWzvcKjslC5WXa2gJmGdI4
CY6faROF2025nDnhz2QKBGPWmVsHGD5mCeDvzoEPNK8Ixbxjb3NGOKp1fuartay6
kdXPTtS0XujUOviPV/v7EG0Lvqcl0nNVn9q7TKY7/UvxT7SXrcYDShBE4ib6rUYx
87Gg7RvsL7ezpYcTFRS/Ffal+129t2UsZYckMctiSDcONQyBDquixfQi/bpGlluT
UmAwyI3Rc5HYjlpWcx6Ih4DNE4dLtc1XgGTvUxDZTVkRMnz+W6QD+zuVq9/UHWsm
FwEoV2p2zaSnYu8VK7zVMJwtjWahZeO3X02NEKT1dQT21cjeJjPJowfsRxwzEcc1
bt8mq3bL9luMpIieWy6tx9FTThMcnQIj4FDC+q3MKJUUGVV0qQRkDxRpCWPS6ZxS
gxCSS6MbbebtzfUTU/7WUzdiWeRNryU6LKEb3xlfRf71er1sP9k+wBlMD9aX8Xps
jEjdA4wlw08/48kfwBk3TbhuwTOzvMAbHbpDIl01cacXqwG/TNUCG6zNq41M9yVb
3hcgf9sM57raHU0UhLK63EDFCs3274D46Ns7iHx95A0lgQWahFALdNyG29wJ8p5M
J+5sYBvzucTNFsUWEYOOUdh16XcHejfwWdLN38At2D6Uh+75meKZllNR8aGwlvvm
uxPLs5D1PpL8vk+/6Uf1W5bGp0ji2Flne49s3wXbxciH24NwZF6DOlpjwrZTC9OZ
MsxedYQj7K8+tUIp6YTybZLor34o0Rryo0OL1Isyg0qL5/WsfJJQbr17cnzKZKd6
yrsHFkiWsa2uuZUyx4gvH5ePH6X5fyh70W1KMZa0RtrsHSnP+s0JgiJ6I4dvIdS0
tTPgK7+8cEE1HK+dhs+8iwHWgjWmJGtqpOps4UPAWQInvFSfzLULusECQkdZ2yiG
qUjzs0jVr/fm9G2Nuj3+ZofYeSC4KeI8fBr+DHtTYpQxOS0YzE1VCWIX4W60+mH+
QuSQd1plIvbcng6sUYtesLRe8y5UPxa9xx2p8WmazqrPso2rmJGDkyMb/IbkzzZO
2d4nk19nuCJkJju8lDQEBpbMnxLEiDK5VqdXe4y8yQe1YC9yhLrPD5rL/rah4fvz
110WAXTvITmBBl5hvsS1l6jz+6aT/5nBpkkrbXlNWuwbbuvNkQRIB2QgGkV5bFBb
2/835gA4dJS8AkfiOzif8xwMgLRg3JHLAEtPgp6bss0HAxdCFSgCne/UzeCTvJvA
KnUdcvsx9lXz3c53fToiGYxlb0TsDLnLC1EJFINYl0ONDBzy157BlZ0W3DaanAiB
0vECod+jORzUJEugeMg9uEZoFEeeXI+qf4dQq8mydllVsz0oauZk37kWAPN+K4+u
ROVGAdOW6I+pVWKZfoyfxw6dR7xu0kQ2s5FQx0ygPpo7YOjFqDBleImvjHDXngCB
3AUJei5yMyoZTF1RbBfeagvQ5cQxFJofg4V8XSdAdQ9jlW8dSUCBDEyflUzp01BN
zuggBnI53hVQrZQce8fslNeQ6BU5yDRi/F7vY5tq2h3RAqY7qy0qCfimbFJfC1cJ
SeACAC/+Uad2co3ztdNOOqV2VH11kfPSujhAkRF/0dEFDjip2otRAuPFQAWF0tV2
vCTNWE6QB5mrAu0EURbi96uDCZz89ibljpWcF4VyT4ynLlMNra8iHW0qR9bFmHap
/5g0KvUHanmRX+xdbDRGI28rcXzR2DjYkbC/McpMwm0SkxMSnO893hQythXMNAHA
ZyvtyaYuRFjidjh7Juv3XZ3onz6ddEA1ZclMJmbxQmB/ntR1/SpPo8ZoL76m3S+U
YLBcdx5tyh9gT5Ag4Ugh9i/12tctvOH1Ocx8DbxIJ1CAUGYL37EJDfadYSTU+BLM
5YcEAKuIdR40F+o9TXKuHvFHI95C6hy2zbwJER6yVQicOis46V3mPIyOsRuHgbS0
k1I0OXM7lk6mH00iE0YG35COhwfTnw7B7w1zbVV0spnEMlPFCGhFfZW9Q7r/Gh6n
1X/xOCBDHuQacHh90kx48OLZcC48rtf2tiXQjUyQoXAcjenq21taHMguq561LS/w
NIhD7xXeltOnjkZ9T3Vl6MRFvOQsKKRXxcPWzFITJR1tLPf4ZuvGg1AaWKtWLDHx
QQ1whkrolcFBGxZgJ+Ny8AuG9RPhzQusTs1YlfqTgdHAM31qUsV9XCfi1DzrlZ/y
+kTayh9dtanwqrkYwc8NgKLbzk8BOMI/hZyCNJioZ4p8W5i1iMUqZaqi38d2NC+4
k8/czUwJDrbHuYJZa8iM2daXKAvLsMcYFjoEJiBiKED/l9tvX0gbFqu9JZc7jLPV
FIScS9qmOlJ59VVo+C/x1jXozKo+oUgUc4/PALMwRUVpYR4ocQDmQorlDAlKSpmk
OyuYZXJaLVD1uyu5VnK3PWqV4v2pVp7cFOH2TfnXXn2St/eAurZjZ7B3sBmowB4a
vX0IK2QyjTDQuqAw6npRwu3Y/VynWuiB/lterKebUXGxjSo7h1DB7ZMiO2wHyJMt
DL3uf7/OrgMP7yEx0f6Zv58Tbl6wcdBi1SDQKI4c0r6hFzcNp8IHglvMg3CxN15F
FNdGu2uUpLkQD/zM6OJTsgVJyJY5yj+0/rEMdAYIybsJGN4nNehov+anz3GeSq3M
ZrDxPpC9ERKOKQa2gtOxkSnsRmczrHJdrgLGkAffokdq1E7HWqeygrtYjchIp1iq
0IMIiOy8lPpx4Uce9uJ1FSt9yxPBVLKQDfLV+SwBY7t61r+nUUwTLftfZPxuaR6a
p7Jsdpzadi2q/8leoYw2TEyCo+Sfd2I434xzzv4JsYJl7S8oeQxY2OYPfjPQVXyu
Mo/nV3BpXZwgcZV33g+cExT4z9AYaFf9ubQLekwvk5W2WByk+mUkVmLF/7sVgZep
sS9MkkGwf6bd7qgpbVNn2w6Tfiph3PEk+cRgl5b1UFPUjDCGHTVx7LVuW77uG0xa
MwwtN7QZvOj9atnXu1fVaAQYPdxp+qwfdADyLB2hGOjKo7NKMehd/xBAsjFpiyza
Za/rQ+ZE1/G/+gKUsSyRomz13UeDO94yGA/TZ64iTDmr1L2BHkKf/DDLqAFB0d+x
Nglfo/s/ye5KmbC1TEA6zsmb4/pyEXBS7X04/aXVYkIbepLFTLxiASjXvxuX3SY9
2exbc9y/GtO5ThjRcyKMakMBTe0qmYcgkiGF/sZP7dhyeswGJs0ZcHU9MQjC1IXW
tInKw/P9+42XueNZlITGtuXUKc9o/bLV/O6JN+m7KPhNdXeEmauA2TXUidUyAK40
Rbmr8eQQgc4qAYK6SKi5kLR+vfQt37gII9TbHnca/nwqvprD66qCPM+ONFFl8Hz2
WXEs6rB/691VeDKnWtLFIW0eE6nCK5vmG0kF59scRTdq5HoYSBbqH4RiYITJVLp3
/m+Zg/ZTdGPEgHviugSVN4qYPFS4lpJ0jq6XgAXrQGYW2tMQp07kIh7Z6VHluv5X
v4z5SNr6xR7WkhTGRb8Q5iifMAJ2kgd116D3KBq3XZHIyMxOzLEmCKLgjN3IoPUQ
Bavr4kkaMZBryQkqpKmqVbzYd4c01aP1GD08qkNknZEeMSqUrs3n82BGwZ2+u1Ag
raMCSF7NQcB1+zsFt/mqnrtUKvxaLkFCFrQhmYY/M15xv7aA+G/+Z7gB7UilDAYW
gJucLq/xnnwINcFiSd3APUbyGbQMmTaY2NIe1HATMo1dQQ9MGTOxKIE/5TQqdlmb
LLcf24cLm8X9Xgf95rLt5RX3lAueT8L4gH9xx1G4bDx1HCvdoqOG2v5VwYIe9MD7
4mcAit5qT52t2krHW+ARlzJmCwjZhkWDrY0FHfx2MUqqkG77pxAU+s6WA7R5QfHC
hkmcJRERjGRfCydTOXjOa0nuz2bPbdiVO7GCAE7X0J1EezKYK6wDyVqN8rA9mbjv
pa0ux1QpLVSjntzjjJAl5gM1cUHkj8Z2ApruC7rshiepDG1xOoTGQv4Q2gb37PHi
cyihmbX/b/YlpVog9pUQoWZteFEe6o2tohK7vQH4DIXT7Bw4Z6kSfs2rKEdCEEhT
1LK5oWcWSFcMtuYnK31r0kcVUORtjXyAAxZ5gC0ou5qXUg2jjfGaolLwi/MJgvsU
q7YZ9rv/zhyy0wopOGTmdiyj+RwJaOpIbgX1Kv8t6Uh7pUhotvkFBPOwzlZx8Qg3
pVqB61bIg6BzcKiKZaQRV62R7QzjLA+seAijmxy71fWGTRqpvsDvEMx5Dqw/9D0g
Z45kUmBqX7nRRubfwpHGE+avTl10lD+ShBSdcUsirB+6hw+gusGWK7uAb5pXQAUA
k+XihrttP9ZcT7rlarS85zUwGET7nHI84Of5Q2FiV7VY51KpN6dOygLei2xJnWTb
ycbR52vft8VC9fw4HHGcrQ45Gunzyb8fqHq9uudkS+ZHYq7kWHMzRuIRcozI5Psq
iMAR6+YLcy3QSXkBLb84mQNSob53Dchvu7E77nr80yt1obVXDK27+P5UZgyDSPLu
yRpimWnhuoC2X9pMSAURL/KmM3r32raG48qiZudpFsXqoSPxkArPtFDBOqA2u/sa
A84Bw5hHFI6YOii+Vr5peEKW/TPsxw8OJzU/Zu5P5NNgGt3ekKRCpGpDqP3yVDkb
2P5a0wO9TLo9clNLEI/TiatR/r4IfV9/TIkq160MFO3fbrHbnHKotkWZfQ9VPb3y
Y6hOjKc3qaql2OyEAKH9M592J5vaweJeOuUJBQOO26G/Q+BrBtNiCjKDzAgCD4mo
sykeMD5jK1fR+6fgvVKBrqHRbpQRPwxV8HhrpWSAp+dq3BPhpJlhWpxOqkiiNfAT
P3OFJwRbhqlOj1JeOlCYFEHquO1Prfq9riy6kubddOHYPlAcO3ZlIWVhaXw6ikfn
/5YdLh205HXo8BZ9F2JR8BuBe+kWTG6i4lYd2ifebwsSApdqBvNZCazZFlGXUMnT
z3QZTzU/dK4oX6rWUzwXRR96LCLOgvG44RwqEJpvz8lQY4QlgVwRk3eMh5w3BdFJ
YiJf4rIu/TYrHSW+INoTZrfh2d4LyCBnPbJLLm/eXymqHdRYNctxkXSbbFwfjkwG
/xLrNuW424p0MDAatQkDkZSN7pdBtS9mM/hPf+MK0+AcSFWpxFXNa+vsBKOe2RxY
avz18PWOhGUw9zrsiBK6/5me99EZsU1D6OnyFOpF6PDmf/j+qAtslh8wyp/Aqze5
fVW9KzfEQFWnh9YUbtfx3kT4tTqZV9rJ0sCGAyvSvrFiygka7B/ICUwPCN3CkV9t
ec0pAmayPQ+1uvF7WHHSFOTnEzfx9OMtQ7xrgAs3ZTYRto6RfsmtIcYjCwFWZPYK
g9A/YNqW7hRE5vrHbLrHNB7o9fhsWufdBt4W+QSLDlFdiDq5PFzxQwxYStFgoVjs
8ffDNwwnXmR/SOLLtAXJ0jjM8pEAptn46zeZZNU8gn36BeUWBv+ZckQP0SYEwK+B
i03YU+tnGWFMAI9n5wqqX5D3Q56nUivU9SqAlus7qyMcViMGB+WPZErGjs7BOXU+
jK99+xm+s508MAcrpevCQHDUuwpQmEIiaQW/rLWVZzg7Q5zEACS4NSXFRjlgifNO
GIHHuOQnF1qExD1lukVqYTYpu6PeRqAVhB0YsRICBJLINOszm41bdR/EK4McJM3R
EzEXULUfY+m1bo5dTB3VOSSY1uLrfQPL+1eBmOm2dQJB1+VpacDuHR9KaBtDhUsJ
9MGmccA/+oHQo0sXk82IUyeFlLS9LLd+OWr9VG7msrU7PYPw41EcMdKCyRfjtVKT
kmbjRSYlVBRBO74mWelYsOFDpVpkHltFspactVFRtgIU01GdMEe6p65xmSCWXpZE
NgqFyBME1xj/9arqNBefKNenlUhMZ6exX/92nb2eCjSwdnY47d9w4GJkiN5oDims
QjnHMFWHVdtFeX3mZVQkwoiuSdW4vwA/kJrmbBMOJ0kA1oZzbEmQ/n9A4CJnYzhK
Ht+zLngquGPTe3rFpEaA9F4YX82toVMfSp1yIkEqQSI4/hzztZlxJGrwnQMnq0aw
Evv2M1W4ReY5HIrN+UH2Nbnhin5COMXvMQA43n1+P4eIkXrjp/67Q3g4HAZpB0cU
VfztgzXJCZG788GDOuB/JXtwFY60u6N071g/xokKW4KaHEgq4qiB3eS6Br8rhDfZ
6me36odFy0+wx8xIhUYBwr7VYm51R+zQ3kgzm30eAFXFnBgRzuU1G2FNIX/WI0A+
OpcUFCdmW4Kh2fuVT0zOoa58UUmW4k4T/e4mTJjlp7gfwQ4MZFCZCNG1c8lzFvSD
n+YBkYK3FJMwuRJn3DJ449DAK6ZbbSf0xdQnz1Ze6ZFZDHwo0tmtbyJIsDyTmpuq
lTfMRJ0TyxYnsN7g/k4FZrDhKqxIczm2JHCV84IfXcRuMZMYv1DWGoP2evnjEdoa
1xJDL+wwBMYY7tEyolpgjFSW5IdfCi+NF43CwBbb7txeEHJ1A3MCJFuFigrByrq0
7/2NUMiyyG8dP3dCUIlKnZ1sz1vn9VnTcRo0FV7SCfUUCC70t7ydnCAFlWLmo2hy
CYSOP5x5NVIur8hqCRolPk/R0Y8BAjF48sL5Fv0J5sr6sXSbnPhUrvYSuxWbjXMS
edfO4/tKxOQkMSmdvSbweATI8f2BhLdcZC7bEkusaqTZebXeUsZYELNhWaEbRVll
2Ip1JWcYLyxJpZlle94s2fMpEFTLYrvO6aO/JdzUyuob3eStULZ6I5/+eOU2v2bc
i12gs5T+T4tWRCgECgLUndqmvtuGEj2gSbx219wcrj7HWQH9CVTbShfEBjIXWHGW
OxQWQPzpxeDXoS8j6X24qmBW3la826wrPXfWL5jtW6Hco+kYGeTBRIXk9c8/eWpQ
QluP4WEB8LXh8aT5zupY0ZHY9C9TcXYVsJ118I6ZeypeZ5xZvO1pKIp8XFaACYO5
qA9EWVOFvjIgNVA6i5OUbpvcGJ20htf1oYoP7zMLRAxfV8uU2N4rQ//iEQETGCYb
SNWgsJ4IXvWAgCZYFviIn6rhtfEbVrs5c5PaDuGcwF2IbpS95Xn5tTpuMuPn865I
J7I9rcVIUTYMIi1DlvNcfh+FmqHvMaBX/uL00Sh0SLEN9DyVsBSELdZ47GmwTYS5
WswFQvkwLauLjhJEqWh6yXiPeEvurG4tB11e/ZesKmgWSRqmnMtcBlb46vGAEyPl
YxmHikOUEV+CtKqc5Dv8Flma34O3qjtbJLYFu9ZjaR3mNfy241F4FwpCWksm70SU
45GtyBdbVkE+WSD/fQcuR+IVxKZiHCmZa2ceq1mu3mWlsAU5DSS/KnPwmOqkm0j7
A7781SYri3VvIn0t4KC5ifykT0fsmlNNHj5QcgD2oeujODry0HxUt/EZ734t/YWa
NjCuezkckiUEycRgbt7susgtgCBVC9aCLJ9z5veW2lyjzCyKPcYWn66E9uExpfAr
N4IZ6OUZM2rjo4qXc6x2Lfarcr3MjhQc4id8N7grY81LJ9rQWXnikRKv9H2ELtio
GFbZ6/Lsn0anxHBIpDe6m/9QIP2Vbi1cgBsZUHgZ0ZWIjEAFmDl/hdp4ppBr0eHR
UVX9y97tALdAssj3YrglzJCT6W/MRGZK0/CQNzPeIS5cXFzkP2Jdbd+KKUlqVtYZ
fXTdFf9Qg3UYQmlYak5Wnh8mpSSjUKkDA5YW7l1zwXkqn0aNgPmTYXsvgWwEnZqO
aa7Tf0/TaSCeqaH0wH1lddGzTrlHJt6LHebTNxULMCVtCfczRPC9qs51+vOxtVR+
izWjal2k0+teXEZcAqDsQlcocg5XxTRVviXLzJuNYnnaCCAb7deVoh8fBniNPxkl
h8/KZZaKhCC29tUHgtFzXeG9oAKD1BWialB6HzpnSnlzrEjJo301QnHdNeI57rEh
+YGl+R+nR374ZFenmyDsqivaoeeXwJKgbeTK4+Pu8pfHY4RQdi66UdgHACLv7/mm
BIZ5+KeTfcHxThPaMMaOqbBzFn7jVvYrRe2T11Lwdzj000iCIQu1Smtr7LsLT2/l
SVPD/OaLzERNU022zfHtgX66K6jSVsi2LDu3a0kLj0wlhSQIcHfBGGnZlxai9nuo
KNVCKWkhYYcCKaFmCXK1xAv4p8QjJFAiKRtTUTCMDUHeaaQMgAfp1mHsxWivH9pF
S5U0MimdxVOKXuY648thmDdwMKV2GP+AGawPdx1rG1YnhxA5ldHGJjx7k6XvdDrN
zr0W4UEVcf+oA3pug4qv6AwHbdAZhNKq74GC25ShxMEIcFkzEvNeZZl/gzNsUa+q
GLewEr9C06eR5bd93Qbb3KTxsvlxPt0caY1fSxTLhYDeJK29V15sRuCFlpLaPx9P
IAXmHz36xvBIDnexHYHR/Umh24UaXSRYS7ahhz4w1naOoTH2JZh2uxi7uB5eifqf
+k1bwrA4DZARQGi7X3w8z4GXTTM0735q66zrTcWMfrfZWJAQiO+Wg0E7jizJMhV2
P4fLoBWOZKgBZYW/8N/Th9dJDB4V7xbgSsCFwZsb+dwEfjb0qxlyC8YXm++4+OhI
QPre0+ObGJV7e8oM+CABE/7mSpXAGAss1huiB6pNGpeU19n3hpWq/YigYOefvWV+
IWdKabzA4zfBndAT7mr1W9+e+qH3XjcAyLvHjg+8NDvgdDqICExC6LkTPf5wBbLO
NDM9KlO6l1G4m5tcNd42ptxlcLQ+Qj3fOndtp5dKuGgXc+X0COBX+oFZqQDUygR9
JJd9lkqp941FXglLEgHzaLcZYQ79JuG/ITFoJTChXsKJ6ETn/AbcEI4HEcJjc3dC
+ibvyqB67Vb8jELofBXFx25G1K6DttbU5+3qP0vJ3THRSr3S5wbjPo72NAt4hq3Y
uk6IzfdVKOXaFJfiRSc0+1H5OIcAO/hl5YNeW7YHRr9XYR52nU4J6EAt/PFx0D4N
iVvB8UiLxqb5GfyPVTE0jagRjmvw7w6eeppyCulhZYK30Ms9qgxpgeYi8qbqwrHF
SZpVy7RLB4IWX5+n44NNU316UtEUgzk6lYxT3mVmWqVDgou6FohoI6zMr1s9Vpgs
+59cMrrXGEYXOBONhwtKn0lpnrhrUvl57LqTN6JcZ50CXnovwBkXBqEXOBWF/jvw
dkB7lWE5UXNno1LtFgnxRJjcLHIGpcEfa2q688iq/udZ/GkZytk+l5/f7yWSH99z
MG3dpDfXjOAZocG66sgS1/qW7aXemL8yoZ9LBrQIngMHkZ8TeE2T/amBiXRn37or
Z4s1yJwIGX/+AupZsRLu/7mAG27s07gia632IAt04UhdiVXwlRKsWkknbbWRxjWu
eWrsHnN7nyNnO3sHedydV37JbeyLkr7Tyq/Y0rHMt7XX+7DBpCZ6ZfpM4Ap4g09K
1pddGYJSDsOM12SDzaI7TclXUvsxBtM1ApNB6Tubqm/m/PKy8yIfBBkFp1gG40kp
ZdMUKFCzOKSJo7+LZISew/BwPm3QCZ87ZgVdzpeRHBuzQ0IOozrcFdBQ6BfkdeLI
Cu/JM+zs0Cb2yxSyWNZTlY/mkCJWdMWma07f6ZXglg4rTiFYtxkLs26Mg0E0xNiD
TxdTO/hmF4oxGAf7y1wg/uPsppA1ShM7gzuTL26FlqwGSked5pVe9snpaUPfsZ6Q
YHLnOaY69j4+P3keM9ElaCQ25r3WlAsyfYWxk3TsxlxCUvwQ/wdZfkVjKUwMjDWU
UgD+h0UQHjmSvbeoY3CiSI+I1ELpNzqEdK6HrTaAjFyk5s4MdbDw+gwrqTjuUUIU
F/sDvYBHom4EmWwadNqOLyW2dWdMbaHTC6bjeOnimF+Vwt5+Ezr7s6KmmHJe/kTy
H5tL090haHL90POIgq+MUaJblGgjAJ8PNJ7Kx0IECI6nCFCOq1N7ffyvQ+/dpbkO
0FMSrM/xX2YR2gksDZ13hUVO+NDX1qjvn8g64zO3Ldx/Sx57cqcP5n7SfAPuLaL3
mCOK3vr44mJrwqLZYUGsOIwG4xO+5k5R3W/1JjRnSJg2CsS7Xyi/G2MnMTZSYhYI
cCVSN5AJWHOZrLuelmZ43GoG5A+dFjrQgKDxxxeqYlO50AwAKRhj+7oxNhqbNKJp
hNQ4FWTpGO576JnW13AtEgEauu+wI5hf+4S07EQlRlEoTX7JIVdl54BWSG3OzeXR
mL+Rdx/3QUwICGtVyF12wJrS1dp0oY1vZLXCdGT/8DgcXmsC/5KjKWja7oxdAbl7
1c80gmwfrssZsLzub5yr2+Pm7yhWgM4FVFK/zDWjJMM8xZDTkJ5Xhc4djoNIHDdA
HtCpi1RRhCpqRwvtfsT747KGj+a98EZGtGpRPKk7AzX3h52/spRrKxkOyZR+XR3H
17aPsUcFqoWaeKShS0wQujIMVtDPWzP5ZyPEKIk8J3Iwa6UxwcFiCgzacDmLBG1y
Z49MBGT2McsF0+kXW38NC1QWZV4+il26soeQyoEa7fG4Jb0Mskz0LvbWTiBB7hLA
3sJi5HoIpI8GltgjNwcuSmBsCZ6kqkSpc2sRjQSE6JVlcUb6xgt8NI0UsiPTQTBE
qs5BcM4nCxL8KbNr00ep29atTCBq3eei84Dynch39I1js+ToDHX3vK63C0g/kNNE
anP9ssTIKFPzdRqMJZfACDImz6jauD5Vu58cRRIhareaolhXJW4W3yOFS1k/sEe5
Ol54jegqOO1mSZFnwhxf4ErtdERaOKoxuTwj5+iPqWzR6RtR/3hUegh3v+or4xg7
qVDJTXUQAnLWygQPoIk/10lw3WR/VM0GrSHeBXEnKw6g/9hHGd2jXyFTWZkHcYmz
/GH0aXwnPdifiU54jrsh8c/C5rhI48r+HvtAAQSE5JzNcCoKbwTdEJLTfKDn8W0O
q09meWHOi8KNIYEPqrFxjA7hAYhDA9ejgkNjllMElPCA5Y0mWYR4Ttnw3pf0hfpV
d3OUZ1wuTcYWzW8dmCnXy0B5s0gbgCi0BjYYFEEN9h/RzEI4nYZ40ZSaJgMt21gB
UpM6y/q5q5s1lQqzYreie3NtmxHE3cKzuaRLSWet6TfxsFDny8Bvr2XH1YQIluwm
1CdtYZJ0QO4GaXfv67Eh8DRs2Y/l1PnYcSdUOaoQQlRAFZYLA7uuiOmot1ld8HH+
ZlME9J2aDD1cmxF8gEZxbpKTv9m/DelNZKmjijYaCeJ636X/CjjlDjiruJ/3s6+w
QavbHAmpUig6ojKDAp2Qw8/hNy2dxOwAZ4vnBXHQl2Q5rcNghpXiPuPNI3d9i48q
k3POe7GzELq6TUOxyJcFUW8HDLxmsVhd32QfnOTdaGv9465xqLNb0TOo4lnrjeEf
7xwrBLAoZT12EM8YYleHfwuRx4u3zhOW2txQMchOn35Fh58seGBOuhrQPeATqFNn
5hJ9tb1DdjvJIicEFl7sZe+s+hnlqZ3HlDCI+PigoJFmDpxj9fnuOc1fMVnfen8p
HdMMWCqblZX+LBqUYqHawaSiPgZ+EIQcGrbBtt0cRxmnsaXCsS06VqJyWVhia/lj
x2/epgIgpDx8zZ4hnzKLtL6qIifKOEf7KQkaUyMAne/apjfrbgzd/AEzNEmS2WtS
AJhPtkZc+77wNAcde2k1HmVyVd6Q4dd575gn53OXl51BZi/oVGB6gltvOSTv7Lmv
wys6XvZNB5f6PP0JUYP03v1amP7bFx/C/ucJ2btVU9pYTEkG9JJE0x6erbUPC+aZ
R19aPqkB3NEIrKroLLGOMpb+e6lVMzdiTRNSMZXEqg8rjGI5dp2NAAokVJ3yRoFx
l7zYkYhLqmIkv1EWxvMjreNZnK6bBvjwZ61TNVdm09T62/fy2hHxSAzIq47nQzaD
lXQQf9te9nGS7XN2+zcI3OBV4WZMESznspl8iZUrh8cJ91xvhyJ1hW110kdX3iFg
kGNauHIXLpLdKdq4EvFDM5XyXxe/QLU464L9UT6MXVdKR1rOqMMnwcL97LjBXvrC
vnuE33RqM97NXOl0DsAmE5+RWlTlWUn9KiNKsm9yA1kge6TKWWuJLi6bpM8P4zOx
u+AvoTW27Ah2R241Ib42iwLOx+HSjcL3Mklx1tHex7e8lw7RzrISy0wHJbbCSMap
n2rAmGOxiyIplLYxlEhs4gljG1g/hoLZNHfzM+sW9n2WKQ0DFIrIYiYPy8D06+7n
mI/+Jx+qhOKsKXjQgeJY3SmhY1tg+HZpTQJjPlg0mcggptSpS4AGJeuQrnntXc8C
mhBIIFZEB7m3eMqT/Kat9d9DTfeoQvAJBe+UvslVoaRQqKf/OlQrcEltaIKNvxJR
7mSCM4UO9nGDUi5TrcQbau4tD7Mcm+FOQf8Rc1686sPnwOsqvq0HMMFQEB/gcJ+W
+haWsMQdTjoxsPsZ5BgXm1QQ0s2omerz06KVBwJBHJtirMMicQtc79sFhAip5YKq
Wzq5Fz4sH1IAImMMUJeolk4MbAOFTjkuqHQCEMAP+DVrs7+Ynib3oPIRMIiaDX6a
m8J/ZW2+39uizdkIzfyHP4O7CltRfC8ITQy7Tq35Y33+LxfylcgwEmaelLC7ETDl
m1N5UnXFeklYB5H3KdjiyK1vTNcerB9CBiyjPgDjbxFAFyIQGP2EeCqTm5Vwzntt
z/tOMhU6srAdRfNUoonw4MVdduVoIAvRbURJZm9XZRKUDJGLTFc10elLtDrdAaFG
8f149hzkMNLLy5jp6FGUl7e16b3amHefrRGu9RRLIQSsEIfbYPoROVEatvkFCmJZ
mkfbPDUEyc06beAO9YqZDVO1RHy/5twvZ1qmed2AOst0wHw7OmrKliPpWp7eZLEb
NG/rJ5hlxTl/OlEGm3jh7Jg47W9tVl0b3/V7qKMu6PH5DX/dw2nwYH2cf6O3w+Ol
1+/Dnhr2HBE+YzwvJxlrtST+WO56Uwr9lu0A2zlzVBd+NYYppr6EMSDFXoFyocF/
lWfW1J/JW1IXCddYMae5CMHfpEeApWYfTV8SX8ZcTFXQJ+KQKE3hTIVKVbCFeaal
V/ZSr1JpijC24YI6CxR/nc3ExEMud11XqrUK5gSxhBISR19W19EVMmkgYexrq0Oo
GveWrcu7VFWD7UGZMQwXLe/ZO/URTrOFjZqMQSdhfXJePMLDIglJjPtzM/8Ovm5v
Rn78++RdckDmRgx4chCQumHhW293kxovgsmw+qnP5iLccYqxvuIjeio86tiLa8xX
JR4bcSp+R/AQyLdRsLJp1ywnnwZgj/8UzGbYmmfFoK36LzZ9JluaR4Nxv7sZK7XG
GwB1LBtyEbYNfFdi645awtce7XCEvHNOWZCBnLx4Gp9VyQDtITYXNQlQB6Tjf7D/
8jmlZy/8brWPshHn8fNzykjEkccz8XWl5mL0mlTahAi5LgkILGXlOK2ELMgygqu+
vsYERk4FkREf0yeccjnwRMR3jYzKqPh0sr/FeBM1baNrtyahUYwOLuv/5chbkuHr
9Wanw6uiuKiqMJGEGdfqTq8x17yJYTwM+GKeSIosXWRrJzcPlDERRg/jqB18/Fme
dWvi3Bn9l7+mAd9iwEb4PAiPYMFrVVD8Sc+nJfZm76S2i6PLAi2HYTLI+kg9K8hm
T7I5sEujaEXhRSInUUnss05wTZj6BwC6DeJFmQ7edbYwq2rBgsyLI19ZNbD/XIPT
ia+e3YTVpDUTn1HWb0qxsUIdJMmoUiA2QYLoNfIetWxfhallDlREiDC+YCk6saGz
/omn32+XsPR/H6y144vMzjEMGRMdQRMrJZ+EdqPAqOB+Bj7HSxb7rmNCWRkGl/Ul
tL/V4Ad6+astH0P+8B063HN9+9s0jsY5WjIlvt1tdOST58AmX+JjzukX1Uw0yMrb
Fj+d2dxktByQbjqmtlo4nAwuKOJh/XazhsdrHjZFgqFch25rwViYDXPTc+lOGqN/
Fj/eBzEvGd3tuIKyh9uUSRqDixorMoQcWsEluz1dDc/oERjR+AeTsADw+9tcgqNo
QakDt0OQ3UckffLPycvu2O6VHcPVS7rFl3uqJz/bI0f03sQDl0b0g6wmYfqm/X+2
eL28smr34vM0O35MvzPt7iiQMdl/+e9dEdvDOYzIzshbPMrjP6JAMa9LVLOFRXCn
C+8YKsFP/A7OeA1m5sN50CiItwgFEBAP6stl5NNe8Bg3CsTsvToVQj4hjaptMT3h
zk805DDEqYAI0Dzh0X3VidliFsHi/AWYF80j80gd8Q2w2niVgWv9B71d5LaOyvAn
y/Z4ffo3SoGg2dQydMcUzgeK4yqimDYWVWI0qkx3bVGtT8b5LbXKOrMq3Y/eYfx9
uAshwPEqGHhL25gpZPX1OE2ayNVcKVyHA2TgRZZomJ6i5DTCyA7eUdZ4m0bbeshN
4CpvKpKqNYI45anrehuGfU69DcsDYdRMzSs+1CswFAotdnRYOS/gxI06SCUsBOsu
ozQTlLKTEe0moYMjzV41cyUmdncfUYQWAdldVLwMptoVqmzDtGPzBJCYB3+sqq3+
lqHRD0C2VGOoJpC4NYwmnwAIKsPOLQeoKJNt+1MRLTiQgPFL4M5hCXU2tECUZo9E
9ODezIS5lcFWX8/qvaQfvV8MsuqeV7cbMh6W6BTPXdx2T1WQWunxauf34uIeez93
ZI31EtmUshRG4aXjyMqK9kWzJcx/SirMn4hmhQdPDbtrZANycJtZO7GDk04/zand
kiVvsYSK5NEpsVZkytobSANniHeUHG6lZY2Tg4tzXhK72QuZF0mGzhQMtLaWRuiI
7OPLJ5xb/NRFyeaU/1lnHEBZP9KefvEHROlNKsZUKPFinN6mA/XUeJFqe/mfj7DB
x8BeWj9lSnCxynvY5fg/69i0lIAIbPuvf5qHK2oGh0mPkdkIVvfLHnbLRTdip77L
yeP3JegqhrI9SKmIlayXewLfq/r/W/h0I2kZfy7iktSEixVFg73uB3Db0+pdZMPS
eYKec4RXUnKsQ842rb1zKvWtQtJYxmjmZiLt6l8pmRpYQIWyMPh5N8klSVVb55eT
Wg0SN0McWe4VqyNwnlOZE+9sPfE1oxoBK8ZLTZR4dnlURcAqdyCVVuySe5ioVgqz
w279Vav6oVGWKeW4Mm8f10NSwIF6ord0KJmupFrkDHJFYOeBFGXt83IB+WfTapHb
+HarzKqgy+5qykOKVqSwy8TYBe3UVnIQcQ3XrBGokKyNQJUMO2FTJiAe8KgF4s8i
hr4zZwxSBuhPar9OVN9e1G3pZA/PePz0lZ1tJKHWwHq8TTASNSEzf0cYYBnz/Z1S
v/K6gtwDrss5G7FiBI2jTHusPtW0gzSMvMSTXJKb9wQaMxKQ/VAJrA8vT6UISNt7
nIwct2M7UTWlUQa0QH8yIITT/P8XC8tEyKKBSz2g5j2vMyf/bIDhSpcAXXec3SOX
3YdZO59bfAHXbyr6/TZIHkP02tV0BwELWxHaLrfKZfjKl/BEZ9tEpQ+ez7li6pd8
qJRnF4tmhMAvRXUmayatytgOSQDCEs+TAnR9jdQO5kx2Kwihh5H3OuuFVvjRwh7i
jkCss99oEQBhBfaE29g7mAryAM9BcfUB86j4/Rr2JY/o8hcj2Nm4eac1XmqGe5iw
g9Fp/UuMeZnH76MEAQVJXmlIoPIbtnpOkN1VCenfUb08uEkIMe4pkHTrAxMIODKE
22GaCk+RiPlL62/t/fK/n3+mLn7bheElaIRHejIfWXgMedqk5o/uTfVJbagSsrcM
ACWWATN+oc2aLl1aM0XeytBrOZNKm0sMWlr67185T6iHcI0kDwmficCJhE1sl5SQ
v4L41TYddjf6Pb3TPvWTw+GKd9mMiAHKA6tXDI8+tpJ+UUeVUrjH5dkIkW5wABX0
e2Rec7O3i20DZzkjn3KXWBKcntJ04WkS0w8eQW8+jR7yCQIUams5FCigaytf+9Au
5S5ixSfmAdNGQUGJ3xXoRpxIExciSCsCezg63nc5qE1/MVxuN+jJc94G5jdFTIZ0
uw2K3jAEE3C8mvyGEq9TJskMzgEppdfIIjyUAJvBRMSCHnYF4I4MTICU6FT6ZqJY
3AdBmsRS/wsc7RDtcDoOqmATxrQ0D1+Z1t+nTSF8XlQ71rmuh9jMTmcd958kmfDJ
98ILZKKfcNzxkTQQYUspuiCV+6IIGs1KuUHu/j2vksECCKsRtX4S58xfC8WAHeCy
d/RTz2Z1lv35KNW2W1TDyA4J/sZIZU536u6Z54yhkKTgUCBsO4Un1D2sK9fczWnx
BI4Y6uIL7ZUyWS9NyADMTkm3fKKzCwR4LZo/IvVYoBMhQAa7KbowGOZ1H6i4sERv
sU77+lOIlqr4nN7U39BLKms8Y/SapbGgwvED04mKYMrjZYi6etjoccfxUCg+8nNI
asz9IqgeXALKA0fqg6cd0zVadSK4MyOT5hKkke9pgdjF6M7yqlVOKa2MGTJph1Dm
vAsmp1lk/5qWw9ByIvIJiexNwwPThmfZH6T4ODgQ/Qdr3kn4IEGc640X09blfSvr
XdJXCqkFqx4nXef9gIoXp3Q8cEncDFX0oTQ0N8scZPI3nXvi87fO3R02S9WCtC3y
pSicq/vfFwFESL+M+QF9SjRr8kc+EZaK/3ENkKyX4ORJMFobS7qM52iOg3ZrBIw6
mbB/9U6GRcLQnVQNIcikNYjh/AP/o/3o9gL8twyMvISfkemB55dRQQlWkFQZqQlN
ucbg+623Zu1HmLdrKSN9/SLtun6Hq5G2xlTVDNT9FR/xbyAyFrZ0lZxSucbO91wk
uGPCJjR6k0NB3oLNxxzivkuh8OnZsmoxu/sxjrtQWnMsdralXH66N4EbF2Xs5eTH
IDtnXLGe1uiS64NsE3jWS/J0inORM6UU1WK07aS/egBeIIyOdapIOAw3G1X1xpCK
JSfsQiv7zrCN5aaUpeXdKNmQM7KiHVp7j8CHXplNRSmCrhwEBO6XKZQ7Ce6ze6XQ
IuOdS2rL8SChPut2L/c0wRlYtbdCCX4TZg7G6J2Wr8SfTMR1C4etLS5bYD1JNm6J
Nxl6IKPX97BNh+wOnDgge5cFvFj0I1Hm2dP6Cqh9BprFSpicBUBTUYJSbgmnEF0j
dBQDpcgzbL1Pz4nJPuj+4Mph+zeqU3qLJXsLNW9tNGpsrW75RXtkjHK8RC9uwPdn
O6YhhwE8O5J8E8n00aadqeZap8bOBDPu/0QKypg8WVSDOkpHmU7BJD1LsxFngyLC
smhT8nHDzAEf71Yzp9ApRazDpXKgUi1yOMkSMrvI1oGQ99rCYM5G2chy6IRXIL4t
IgNA+iHov9CzetGyODEVy3pzS7HL03nObeZBTpnaCUesRydWuZLS1OmlKCBXZNKM
2E5HGcIWKaaSYCmCr2ojRV/ah13E3Kd7xu58AyUv4hCSQDMXuZPERdb3CAALkynX
OOl5D5o6VLDFQ34HpgEcQLx9OOSTXJGxbzthDVCRvTGgVFaY9YbEKnQc4cuEEByA
agxbSIagbdfV7dMshF3klUfx5CKsYLRvL0YDX7jCJ5ucN5xR1Q7ewfXN1eAsesLm
aOEXQTFgTznUky5fm9vblpaYfKi0H3PIJccJ40kK9i4F90cJxkerThcQOz7WT+uR
T8oog98V6gVoeFc4I529LY8NhHCSNxIS1Mp+2EphF/07cwB9SRY9Bkd3/RpIyztx
7ZIxzjm8hNubblwBojCqu/Q7l1vbEBqLrnEel3VwMwbiBKVqtNC58vpEno6stgwc
fiLmWE8M46O5isQinSmsW6RcgiY+nl72egyfdsGvgU7EBiSlQd0dbL3h0P7do/Pm
WUvWgkP1uMjUbqkPjxOXLbHkG7EdckGBxjnU81OhsTpLrxA3glo8/uoFQSxOFblX
W3MTADR/5TgeRHSwpdWwemvcAkkTG1IOrld2Y0boIkUkTRHohE5xWWluJWdvWhzx
vdKqokLaSP0ycp1Boc4IIi+5uh4umAv+TatnKoErQ8hKZhd4umQAF4l8/mmnWfNN
GRQcGkhTuO6JGjyRMp/GeXu3zftX5eNYtseIfyZvq4oZ4FaPWRe8fDl2hUfZ6N+z
UrgPBUXvihubg6Ocntz5WtZz0jXIJCdTor/Hug8V5BmxFv9yk5IziPUcV7Wk/+Wl
itWZ3mhZ84d4E1oTe94zYbuaPtAbrISwJ7gjFpWeCv+f1f/jp6Bylu6eYZYeFw8R
+8bF9h6BrOJ2u8+DZbMiNNq+rFzvMdIgprOHjrZQ5cXbXYTgko+MtRxVGC/EpK/J
L+CnOnsrbxO9kKBL+rXCb2205nfQ8i/Ahc1PRVIjmpyW9fiJNeIdrc1Mg6mhMJzC
PjL7CJghgq9iIVdzM2YJ0b+M8+kGhRDQVrzjEsZ4ztY6Ymx2KgKkfqbRUailQ3zC
quLsHBsP6Z7EYES8xA8p0P4gNcAOWSMn5Hif4xztU79wZWJLdixov39cmCIatmkc
Jm8PhLYe8CcjKyuoO93FBetjfhE7htC5vHF1J+g9trfn8j2svD+MCpp+HC3pHCn+
vYnhxRRyhsCgZiRkUYzqczQlI6krV2WQzYQ/Jx54Pez3pCcYJsIeOzbPS5wDIEpB
oS5fEuTd7Q4bsSjwmoyyYXF5p6gmEKqbouJDNL65xgpGcZxod9BquwvggJbTaWLn
G/2CL/K6Kw0L6GlUS0Z+n0lxv8UIP8DMi+ClJkMKT6iF5ZNGyuE7gcrgARi1EbjA
4uXOYTerFQa+V6roa7nPik9AWFOJWGq8iQX2O2rtFqUS34QE+vUhCZJ/Q8AlXOTD
cTUCAOP2uNxoRtHQ8Wm/PWRLvgG2Y01d02o4u63Esg9Dm/erRUA/Hf1wkCXe+HV5
yM/FBfUknEv89tTyMGXiAbENOSLtXjnBvl9rTe/ftxvNl908cbk2jcBqVPslu8J5
rlC4n4Cr8X+b6PfOFdTvNmM9wMqCppaIFx198JMzkFy6L6W1M7AjJMof8Ktop+Ai
jwPm4N+Tnbk45qA+qAC8e3IG95/+WkROsyU6G592N9xa0ZVrZVraSR33yNzvo6Aq
vf7FJVlzWBWnOcqE/uDdjX2xKQ0oNp9slQLmPVycB1j6pjmpa8R5P9easIr/1ip6
bl3UOitZBjEsnnTWNYHv7GiTfNVwBfD/04VP09l4e6L3fY8IBNahmiOWvrj+x6Is
dFAJlpDxIHg4iRbQRLKDXI/LIlv1orOoanIvET8Lw10nnRZ0L3bXlLf6jzKZ9eZ3
PIZomW+jBCrjXeYRnIg7oRCFN3Cbi7+Z/730dW0gPkNkKa3PduEWl82iUdU5TySL
1jsfUcDA/eA4jbEMhRblaJov1lPTP5owDoBv0iaqnAVKk5Ljh0UhpdO/UmIDh72m
6AQIp+O2fp/pMeh5sv7Tuv2hXdgcpQqILbU2e9nzOJAlWaZd1L7M9VUKi900x7iF
Owol9Y8uvmiVd1+83tX32cxoFudaXRtNGfLjdxGBoeQhy4zwWowvWrAuP/i4h70A
Ss2OMCZizL3rnNdwd1r54FTkT8ApAs94coqOF91ILqkMxXnfud+Y4sJUco1CLr98
aaxyIJsxrRbaAFWI6Jj5WY3eg7kFyLUXmgVWV1Ki1W0fnzPY0WIvfGtlV7jj9Qry
nrkl4abLQ9PvphuMM+A2jpxK5EZ5eEPvWBGXakD01ka7vVGWnoKSjDEMgfFFNSCR
0I9ROeSjmlA513IQZjvA2uW9nkkg2FdAFqM4jw33IbB9lICi6cex04SNue6n3dfN
o7++c5KpaPtC1N5d2ZyPJMSwZV8h9u0KP6UH8ytWOlKjcKhEKgIfHjkGF2H9p6cx
wEa3ivOxZc6oeXNNmCrglh/srV8DI0kIfNCrTgVYEMDHwQXmtn9JtQ7reN7D7UEJ
7pGDkJAqhrE/hK6oySt7zrt1ammwDnS3Ld7kRumN1dK6dk2LluSCWtCiMpECynv9
Om9icTxeSgyaDoPyp3UVUqeeljFdltBT02CN5xfrR8hTC73q6V4uVoshOSQos5OC
rHMHMEnmhwduTUKxbOpnGLmrTZJXABKLiu0bAZtTtXcwAO/lQMg9jeXPy5aL+KRq
DSvxitsRM7gy0Qf/aJjoq7jSkNnbi2/+yXt1FghKO94cH4IDlUgropxDmL+gPgZZ
p7qFYZLEzd/ZSbnq63JFVayEHe/NtRlLD20gZ8yPzBSPke+cEAxTCYCt0aqK+vWQ
BAUXC1anQxToy/0k4baLk8uaYTRSzAfZbYbpXoxno75lAQv2f7KHelr0BgwWHQ9F
3Avy/DHuqXI3vF/0eZTjCWZIDoL2qMT2gjzXZpe9W6rxJlAunPoAoYwGKUAYAiQR
mfMUweOrcG/HGzB0rD8rrl9ImaRedE0ACl9XF6V+O2zv3icT7ahm0QfsxL3nKG6W
vQ0grDPGzS06EVMXvWnr4O/Jq8IiZPw8b0RxOARILQEoNOqiA56A3JULrPTHJz0L
C8ywWwQKF5Xn/z/9tT6Ce/X6WvwwQGDbpoZd5O16JvmNyU2iBZLbjOd0LhWxeDA9
wolC6LcVvw0m+dKxWsdyX3YW/FoPinneP4izUe0hHgvJn23HKJdVR/Tlv0793hMk
CeqRtsANhEH9yNvkjWilJmzXJlgEkZ7u3fjQ0SmWxiLYALEi/QRnRE9TSbkAYFyr
yN4ExpUgZCUAeGDLfwyBnlqy6NmBME3e6oJUIc8ni6Uv4yrjQkmHYO/1RvBs6w7M
qrLWkU2lZqxziwVx3Vrkmeg+bpPuWEupyOJ1cYzpS6amFpq6xwZSL3k+nKgFvFCf
cx5XofyU2KXgGTK61dIcof4Wba+A/Ix47vwNNoNgj+Vesoq4J3dPvgBIekp4kTQi
G42ieuz7XbaUVGw6eivEBtXtbdZJJ2zIj7TEzsoN3ySnHcaPFF4+c+iwkt0AxGXP
jZj2K5fdr4anSKCQ4z/5yyrJwM+/WeyzbfqyI4mzpRFHDAx+fX20y/T9KGT2Nb6r
/2AXQkmYSTiQ8Mqh8lauJiM0B3YzciLMPGZqGpbT5LIVdhZLqiVmH1pkhMM3V01p
pFlFK+g7n3Q0Y7LRqXLvg8ylk/oeWc40LQKbC5gMr4QuM9yi05XQogNDGrBPif4U
M712GxJF/c3QcdRRYUCYaSJsPfB6HnY+EuV5MCap4CanCp9dBYDuNws07YwYXaUu
ZjqDP9beS8JmPvcfeAQfMTQ1Bq9sdCcq6GDi0gb4n+i4VAsweNscRi8bNMpudUfP
cg52T6aokZPuKQvDcl2QvaRTa1jq941NQus2ueZclDgjWa1e3W2G8bE0JphC3p/h
9mS22AlFYoEfDJaDjPkV1tb61qD1xHNpAqTnxPAkW86xvlKVqt2Y3jnIz1UVPHhr
KdhoXyCadPMeF3rgWETEmTtib5Xuho8Bsw2MTGitco4I4RnybdBl1xH+fukF410P
nYfSZ37tvYedI9SfTuPUxse9Y0aCwncb8bBY3t9cw7xrqFRKJMOU8sg7Zvofb7Nq
d2ZUhWO9wGqU3nv+ksUJrGMYLtVZTGtO9BGaI2Ra43hx81pFEq+8oNzBN3UtRipN
WKrXYr1iEXoEqXnRoQ38fPL8M9MICDq3o05/VSZhrnQgk5i9BOOUnQ7V6xxCGpfR
Xt5/mt/SUGrOY9cCO6C2bZQyE8qgEbhniB1XqK2D/rvbIMdK8lLraMOShbJDfW84
I0KTl21IsYt+13+Vv0RfJFmmLZZ/etCF0ARtllCfk1w5rNvABn8lLxdV+Xf6Kf8b
Mh5NDKFFe66GGSKJFwHhnrnszgO0rzrI06MKkJMIbN0QU18Y2nrWMCfVQl3KOou3
Xc/7eG1nexZ0FcVc/2GXckXbdlCRI5STzCZApyl/JwKpZWWsbHUBnSjBvBeXUEsu
0JCA3Kw5skNM3Ztknkb5zwl14azrpnH2tvQQmJEWxfcMTxlvG+SiJn9EszOjPZtB
fNg9J6CsyNmxzZcthjwoEZUdDdTndlTY7ZBxs5PERdiNu9NgQaOv5PC9Yt+X5hwo
IJ8bYfCY89KaROwmWj6hGc1h5wj/AKMs/q2OJNJeHdQLsYvOnKxnvasffqdFHrky
tipLqf7UaycprdeXfUpJl6FMrO7gDkUEYkaYLOPc5QfsKYB+VX0WdtRiCMS+vW1R
RkzGmymD74Ngdgac/g0b+wlUIpTNiCZW2X7dqijL3SP0Sj0pQquOT9oCZle2Etgf
o3mjNz2rUDRUVRRCxTYty+yKHigFy2SLtBHI8cqmH+jQg/frgq+7q7QJOWC1Np12
+ySSAnQvqzfwTqFyGQWzg6TtA6s9AKVv1VCO1CZ/CJavMrz3jI20WOb6b+xcov6H
6UF6agCMR1cVamFx0NQ/ORBcxaPrm/2zJWQ4+QD8MzFDj4MW0jA+ygY+9vlTKvKo
FHualhq55Y7F+OaO5XAXREDsW+OdK5uP7X4qEhhZ7pQPhubRu9MNAJyUcVG6WvwW
/b7miF6GZ39pjhAjgfJCWdUGKj1i/Df+PV0Yz3iOTeyBJ5MQf7phNBCEPzo/OhSq
vAqbSQgC5ndYCAQCdIIGLXiLyWnlgEtP888cIIMqikrfSTzDUpgi5xaTRzdapn04
gVqgktNbozxl3vDy7TPG1uRtgEGwZJqQ3lCJui+3Nj4W5lCBKq+Mbjw7nDBE5opd
AbCI23QqN6bnwHuCLUkPknRBUJOtbGkiNV1NkBP9fKvOYIZNGimtdVjPSu7RVejK
ZhBfM3DXNY5Rvi4W0XRJNMsQI0/dyMLXaLQAobUVSP+h/OXWJYA/twVTo5L+5ZOo
Q8FhgAMDCMjcAQAJuo5qcv0OMYZVtTjh7CzB4IpPTbmsMA9NFa3k+antcdRZOT68
RAsOAd9w0fypOXXwVIgX55MMMNaFbz1kWeKVafH9xTGNtAq7oVXEz15VEY3AwC/D
AbqdGmyOxfa8PIUVkZx0ULnZT3nYEwwZejiIGWIffxoIcHqxkGjVXzRDIA0EMVpC
xmWgviPLRDNnXbZDF/CBzZ0oxZYNlCwSlJsn6v2X8rSAd9jooJ89xtVhH42XGbv+
3w25/LBdGxYcFbPUTpBPvG0bUH5gs8iGVAbGEjlTeZpbHostwN6rmoVexbG8gevl
BmkMuYjg346eZ3AJCFs+7JKXXBdWSkETV9CUR/7id/4PwdDn1E5VRI4/N+CSh+qS
WUYqBjYO/jf45T7HEtFHgWLXMYbMjsjPNvPOD85Kic1rQDx4WUX8RMZTxomHKl3V
milzkOFbhtJHsfSwGlCUN3dX0Ji+vqTwZVSCveszAMLbTJIfwTln/yqD/4rRFfyy
KrCFB10dqxFQkScyw/5KBgQfXRmC9Jb0xKYBehModYq3SS1WKDnTLEk1ufp58Ifq
onjlyDSfL50CTDbvg1eqbRHTBVrG6nQCh8y8AGUqXn51tsgnSy3Odu5yTDtQqReY
94ZknlGDotUVa/ukDC+vfaoD+lxsQumGDazMJKIXhLKRiXQxL3YEKjHWB8oMofdL
iSIO12FwFkEZBAdoBdnbiyk8omcXchAq0NFSR473Rgdz324Rv9+UufUUFMO8u3zs
/k25Rk5wX3kSTjRwgEekPEyIo68rjUoCSngrI4dNr+BOB0avusqE0rqpgnAokBjF
RwGXtC5VYCMYgYAR6T9SjjKTc1neW+7DuxkGKIj5e8F2Xu6e+wkNJM7CTkIvqtgH
ykSA9qIT576vU77lnDdkvixbc784pGMLirE3ED3wWvQEFiop0WCUThDW0JYlXvSq
yAUfBKF3b0iyG1U/h/SqSQ03qCzohgXehtC7M4f6YEb0XIzPbE3mJ+gDsE+EggTK
BMAqika4ZYdjtXhOhrvSDj9cmw3/uxWHJaZ7gUQMSnqwFMTl0X1YqRU3aaQanZGe
JZdJnBP066y1Onvut3lv9HqE/QbkSiwgpy9bTWhVr+aEk/IrXh2iSovSPJ8S+S2A
TQd5PEqtdy+ujmrsML0V2FEymRMucx2zPj1KiDN4IGDnF7gfvrbf3wP9Bx7mxcaV
UrVZjiLQTYCs+zmYTalgqO5gOsGWtEYTUzXg6wrIHyB+X/g9SAj1kZsm7n90db5e
7858MCn3sTZHO1Xi23YEHjl3kBU1EiPvGTxjubYlNEXUZhwZu9vNxN6ZSNcb139L
2sixNJcv0Qkc8bw7weqhDKjRt+IhwRM0ohsOoZEItUwrOi4uZHyAI/hRGpt+U0kt
0f1Negj4iqNAYcyjvFW0GSSVUybUwPVOfPN7DmuPstlipIz3UkkBRNWL9ykVmYZ9
tZ/qMZJgJnyCeYvzh3X5cobHU5PfbsMTEQ2W76IlAayyT0dl1zIZ7QyRcAVURnb8
6//ipJIFK7BpzjGA9jXsbbQNTEbU85Z+s7iKabNdnjYdI4n1Z/817gQrpjGIh1iO
8TPYAD0FdK968UfcEYGiHPkJ7rbHvXw5eSRZ+WlErYMPU1/gaapsMXFkUcJHdoK9
u71GKUGVQad+pogicA5dxgzeDoUu19E6/CwUae83CZ/f3vrsTFQywwoZNwykpYu2
2CKL2bWbbs6Hh3FafgdFfJWYFwqFsOXM8R3rEmq7dlXyZoHIGS+MrCWNfS+CdP+S
V07Dz3Jcb2NSfBXrmsNscpvjdW8f8aQdrDbe2gheSLyOiAIZCgb9wpfOKk34RnJW
4wqihLQNmzOZ7nOZuDiK61NlSWDyNOeTlK96kYrAWJN47qbzO43G/etjtRh+VEP3
wwdcYcQvKTIQ+tYnmrDjTzK6t/PgM4YuwmwrWEBdWt5eD7Y3svTg/MX4C5JPAlcN
93ucSIC5AhGsMIBw2qhHFCI7dNw/aYkBo9p30/oihjaRYN1aI/3pdmnjXd3daIYC
MkDawrPm8sg3gRNHqgVIjsH34UquEt/DuA+dCW3IcGlxHCFeemQvIq1I9EdhUyRZ
fngwi6t4YjXF9tN97DII21hmnHxGHEw21QFelQ8ooYLJ2YTMzVjnzo2f+SoQLdaH
zw9nra8aLlWf3HRfrTMEff0EiJi7DKzRo9mzh2EvPi0fNbNA3VpOoz1eokImbvrX
Bf0cs9CIW/grhJVmTh6dCwtm4woRLvSkRE/lvis/C3YCxMYeFuaJdFdBbtyQRvZn
nxaW71pk6SlIMWsAPfap7AKoVwxvB1Q6H65N29eiNDzIDELPC3reiFIrI4ZkIlRw
7vxWOYWJHQOorY9YgJBsTps+j30mkC2esxwVf1rryCZQeF9TX/G6UgJqZxzoeq8B
AxDAVvxAzwN8GytMRyMWLvcryFO85qCEjJw/w+5+/1Lyse1qxqGrF+JxKPDxHsm9
45FFz4ySvau2xVfQmwBfkL9YHlHwTmFGydKUgG1WcEUuX3kFpQCNrQpPldw3ma3v
smgfqUoKqKco3fgNSDH5sAl9MMxVMMg8jbV3uWIegqvJsDcbszXDhxMlKTgFZ1Ap
tyyHUzxjrI6ltMfIG4apnrAun3c3IWILuls1NttplezMf6RJAygOUtiLDlwuFQ5d
msyQa2de2cshf8BVcMXPL87m8I9UOUB1zqwMvEOg2PZ56TN9NW5syT6u4TFXGnBq
BQTDsgzZeCOL+3aQegxmUVW9Eo5ZYsraq6KQOV0WIc/hZauPpM0bZZdZUQlqVGkp
/S41QoIx5hsPdOOz6zgH7WBIsOvDFW5MhfQRrqhsZ5Zgq4hEIoRolDsBiNeIFf5K
V7hFwsoNUf9wFxYTRkIJBwnwo1+TPWVNNr/PzkQrBDkSijGXR44NVrZ62fpnje3w
G5h9Xq8oOg34G+2e7ATI99lVegggVOjyl0eMEOTi2RZs5n0hyaP6FPhi2o4jv+gg
lUgVD/HpE2WFeuYm+9gI+oy60oO5apMg7gHSObjyajOtJW/LrLECXZGlncFIQSeH
AqiAJUaLQvdwXcPlN/buC4dNbjfEQLRhGbRo9Q2/Om26BFiuhJzeTgt9JeH9Bbgj
+3aW+ucDjTy4PBBQarmZ+CfxpMiF5J4sMlPPeVb6o0AJZr9f/xZrv7WFCi9Z1bbo
hgUyBS3Tonn7GoSFnk1DLgmZijAuwoPruVsiPBBfSgxFnvXk2oqbevsm1b99z7dp
I2MhOgU/EzmDV3RMCIk4IAeoGd/mnIjoeHGi1PxOSZ221NAJK06b19YByAiM8Mbo
cSbSYH6/cfND+/ZLZnMzX+fb/LF6XYFJVC6KdBiD3ddDk0vXZZ0PQk80Dqeqpzz/
aNXAKL2oJY3FQ46frjmho8QI/zjoXPsfuDqpZYVlzC1JJc24AUTGZ42SvAOshdU2
WNHzazES/Mfh+K9aBBhZIgSJoVFzFmX9Y5BT7rg7zPljBlsPQkjscYcxdduRKarR
cUoAD9PmAE1lhcWdN1l2T5B64Uitdtt+tWBBzUbnoxA+Vl0KY/MhVl3wwL2e29Qu
8JKxVzNtrgd6Ilq7XC5G5FSbw2eC8Nz6Y6yHUr37JAsCf4l0FfSvjYwgQJZCjrWK
/8gn/CCCGW6Q8Z92ApH45gIOkWaTKzJ2fy23p1RdkiTPiZe2ogmv6k2j70VvqZrz
ey2IPe+/tyBiFA7f2mSU4OYRNZyIIELk35OyubKsbg31i70iHHMcEhrRag44otlm
eT//RebbDMcrrKScymvshlE2ZIv1v9RnvsCDhFWUnGLq75Z4/BUxdZf99rFj+8Ag
oTkWS4HYQYPt4l8gAjgnG2PL895KvW3n68slOGd7UNv1w1Ia3OCKOgX1/R/CYubS
YOh0gU//rtDyDba2nh6rGmnUfdmMRfrHyA690H8hg8z110S1lI0wfiwdTmg4oJFz
olBkD7NDc+nWGbUBW90EHdSdJD/U6xkeYhv0cuVU2d7eAe7TmEReinE3cx1WlN0o
xCvFHC9B6/tLPNN4OrigCBhY+VHQ1knl9S+KtTZe2X+nkYGGsW/oGCvUrpK3vABU
1xfoBaCr8fnvwPvm2O3QTj4rlARzLUpdf2NSuVj7S18+0B5shJLbMnsxE6Oj9pHl
7ol5uTpwD/rKbqYiJ127miK5ufFXf0vRSidfqIRENcQ/xDJ/hiljujBPohRXlfL2
QPsXpmeSHGHUIORjFI4//2JbMXgbY49t5LpmRW/1uBWVH0YreyVunJgyvum+Pzzb
Wh43UOgoa3DWZ3Hz9QODykZPudH3++RgEgkR7d4B6rdKFzQ0ncbnp8oiR5MxacjB
0V2KxPOvKWEcVwyC78TKtqJKoUurFLaf6t+PV+xVoDX527gZIwXtbnHlheubrF32
g9qo4cp0soHX+FbQGBcICXV35Ppkzl3eUzaw7QHIthxRH3NYdZds4KWnSVMWGTrP
gjB2QzKTERsNdBhkaRhVefyrYgAW+MWTHHSGhIkek5IlwVF2shx1jcsXdznVNz2E
Wwrv+9IhRRewb0c4luFif09YBMAZGim1/NFty0WB2WNhoEuAQukw0NoephPNWyZv
MY9IE1dWd7ZWL43VIGtQTVbSI6tRJcfcDqJJYYTJAFe+iYqK4y0iYAunNXiFG8pW
u5A43F+Sls2uIOP8glbCLvaL8EYqTrC4KD6KRtrfVjzgobGrgDtvWmrjltSnyNtG
QTZC53uzyQjvh+ikNRHP2VwUouvyUC17VcfwR/TcacgN37ABl4Y1+6UdNTazr1e8
2TntXevTBiUuKnmFBByuSjlwEBfRDtXR0pSmelQZIL4mciZVf064H/ed3Q+KMrje
3jyy5TtuzfhqYTO63Rnp+W6Prcj3DkJHmB2Lx9esTIaSZhN438uVx46UzcZbPo1K
O2zoYfJWj/jcTetuUetDVECjMGX6Wvni1JN+GDWiic9jjK2HdI//YWf34kRbLzxl
Ov05kByMjI0iAk9SsL+sqiuAZZite2dIOu3RfNawVBL1ZiuTCOFETxFBZIS9FTgO
AEWhiHfTySEPSdnTMeJToRaD9YVEmnGhqOLXMMSxkVaOEFxzaRK2YQonwPs3jmOQ
Zy8ZmBrxjKyTP2zbzK4t+oi3VFM674RDbFbkAhdB/9wYyNjMDMzwhpMfpO1R9cfS
4Ga3qPmB5aFuwH8/VsiRy83XvciuiNhGlxBpw4O3gd8r5T0ZnI9F7HsGO5/fbl75
yYy9OwPftIYQG/Tf/PKRKROntC3zfIGlGNH0kXyy6bev5mrnAxAy/Vnohq1JkiO2
KwTBbNGIGt1fj+rR8zP13ABTTmnnL2WC/U70XDQ08VZR4/yy3qyXAUBbEJ84/iIm
JuTR9kLiSewLwp02Ty/2vj5lduqkxwYgUqV+ElzPEIXmFFZMlcecujCs2Y3+h6Yj
X/R38rkhjXeqTmON3S/bDCjYLfzl8PwwLbjME14c4crZPCq83wxfxiGO4Oa7dhmd
8tVuO3bpW/z1/YeepmavIAm9uaILhb43OVqP8dc2y2aFvctFY+NXlaficEHYr31B
TpAfR9VcKRT6MeySlx0ac2yy8ATk1OoE6g2cjvoSRSVGqI/ueM4JmarnK3C6L0E2
AQwzyVezGkuBVkp5dGPCY1It0DkVXnPCflUR/TI5kTthkYRgkwB/t+ThkJYIe84m
l3PJi4+hOxlstedYCcHKeSMnTggzyHAGq6CVl9nQsmC80FZR2Mt07wZAJiOZ6hIU
hmjzMR5AbsKobtOIRlOq++0yVyXpkc9JuDRGFR4z58KQ0VDSp9ozf1MfgBlFOdZ4
PTsvgf21riDVQ01BkZDsd6SwqmeDZ2M8S/FCfhzmvxGSoUfUHfIDAtJheJvZ/GFJ
a52DU/rCY+qFPTp33KFRERmIaJJ+pu6DvoOmN+U/0i0KQ9lwWkqd3buu9TIER+64
kq7MUCAQ1/9Vp2X25qqGiJnb+o7HSo4OueFyfSCz6NjTIpyh5NWHVLA9BgA03u0U
f/eCHLJpLSBt6z2IfyB8e8C2SAfzxrWo/8E3TmLcrOk572ZD++onmemC0+b1o/Ww
vl2OibmDfqxlOLVulEVWn8V9xITMp1W6mcq8OnPS7asiakDrVJujQt3vyHEAuCYE
xuXNDHzOwhLRuZMIGWbqWHmPGAQmNJGkDFyBKc2X3B3r/qVpenA060UB2gntNq+d
6v6Syd5m0wBWIJcIzmayigziScaq4igDISm/MmV16FSpRTBNzYpgEW45/wt9X3zb
Hw25AzxbmoCEer694tqAnDgpbN+9T+opDwCYFFMwzB5fSCmW5Bhz3iekIWJGpYdP
jjwBp5mqcKfu4LYoheG/1wFVfmgs8PBuZedmx1BW0DFwnatjreuDgp7Sz/i2sBl9
C+HfCEXh2i1/fig7onbdhYgFczB7B4Ad3r8AqnkWaFwhIf9/XxI6Pnm08i3Yn9V+
0qgCuKSTNHzN4BbqFf8DRwFNLZRkwWxg4KUVrerW5Ma9CLsSIEsv5v6c8NBA28GY
DWkSPEVSGf7VHY+TAd4R+ze9sUke84tkExw39bCW7Lq3o1uZudKmSS21Vc4OXoGJ
5BAscD4YHP3CVv+ifSgv8KVaUWgYZGfDn+I2E1iqGtgplhgcQVlBJOl0q/KQMsBX
42IwiWb6uYrIFxxhgl0IoPGkzkcia9tGfDuCVQId8/BfYyPzG+txNRzXvHYnVyuZ
MGaFgHdjHjxGrYLQh/Q2Nbgqw3yDjhAa8Tn1dPiWTUcgX1VRicQwdvh5Qk42kxqL
H2YlPqv2DE8kBPKvPdO0Op4Ln3z6ZwOAtD48EKhDqP4VcLYIRZDvlGgoOpm6N29D
FRXHhDBOylvFZN28rjoDEFb8TuGtG/6+yxeNwuR6uiER6IQLX3hV8mBkuyyjf3hr
2YZ5KDY3hfkQJF7TkrXxGPYgS32q5DNp5PH9M9ndeUSYBgNRwY3ivvcnTTP0Uw3p
FoEHMKEFOpvjtmYAPSU6CQKJzTkVvu7a1qegTZgsGVdkeqAU00+Y7T2fKDg7wEvz
KqWhDSiBjerbLytyk8mpy4gw0pllcyVYxYb8gnnm/HvHkTPKsGcxHAKe16/w5N04
Wf8X0F+/aA2pCEhGfNkmZAqomiikSiouF0r4bk/zJxy2S+suq1Yg2W9YeCmjXBdP
T68ZwiPXHF/UFXuscnEl052CDQb5skFKJyrOYesL6GDHDZLAtOl98tI0wwNOyigU
GsxUgg92QF3KP6yukk6u6aRlvdOKrVLQ78AhBVyU2qSBcDQYWgr+jT1pseqnlJSZ
lAxQYdETJHswtqKSXt6mXGa1djpjBb2EvEpZ18RK8gPE6dcKzIZBvHMVeiojDGmA
/9eAi6eGbqvGU44JCRNrijhQfoyystBCc0MxdNX+AV/jghdWpjLNqpvVkLorkYED
uyh7kTSnV2wltnK8JtibDapyZWKiOSLc46WDXXWeFwEzR+NON/13Ta6/I/OY0Ilo
AnenxWugxm0E4sQlnHaP01uVQefDlOcVQUkRWRae9m5UMbnsvR2sIxLks/rrH7FI
bYyMh9/1XAhdA9dblmQ2O7H38HnUeZB8gO8Yp2GRZNTfKfqUs/CJd14IqvJxi6Vp
ul59SmmEmA0KWwezBmbZ2BU/b5BeIuxZH6tgiwdfsvEkd+bx+iA9JsIgnBxkB20c
eSf14Ta+JqnAcQYSZ9iE9Riy1YIgPafou+4pq7szxduBOjEl5LCEezRHFzA8SdTp
tUa0sMQbL/2f+pqxnGHrdTjWHSjHKYTXbzUv5LZuytPuq4kq5BfCqpt+I81Y4FwP
SKDLkQgOLzp9N+Bb1JkR0iwAIZcQpa/BbtRAmGvgMz8ZAF27MGLUApiLCCrqpsXr
GlGO3ci1bXOXkOskRjBApEkrsyACkH/1chmZw4RYfZToXDlATg2LbEhHTtAehj/H
jMXPEJQmBlhOVKaOlUp2gukGhJF9KxDx5VAadMSnoI69NpUdTseeHBYRrN1rBUgc
r+9gfFr/32mQANF0NnlMQZzU9wnLqd9yB+hEfCYPLCM/JBPP8Ky+IyarkDYqQG3N
S4U5ze9+JenWCC/Sqf8p7xTdEfdUqYKPmA3kFxQobZ7olPxxfSDXFmTFndW0fmCL
M81kbnemF6rmhaci17I1kfOUK+ZA5v3YpaDwmbRtSY+cvydX7YFopKOTUHNO/pCC
D3YqBl/EN2tobjADs/lvx5nIZFwrQEy3Uoz5MD2McyXCpb9wJyRvozHXwHr3DRR9
RxdKGc0s8pJcu1RN6vRLJjX5oNKT4kPR8BMhK5lcKI+h2AsMTmWWkWGlbA5G39oI
gBcJoAnG1UgrNZXCJJ/bADC4+R7jy4oRlgM4dGCbEJYbwLGs9RbJLvSjpurH1CT9
TqGDUV5lijA/xlzZkZ3SW8bzXQCydeGbLluBHQzhYnAyxBoIlz4CSub7EgP7ZRx1
DmPj0ok3fDrxGXU6qRKOdiKEwEWAaVwjbLxWaZJH3MD72KVf6NXvUoD85he2gJei
MjESFNcpQkgW0tee2lUZh5GbVfPgW/lMboecOH9azWlDgg+Znz4Q2AHT6YqVs6Vw
p4Iw5HVsCsvrqcgP7Sj8uHvK9snCHkO1kCbAlvdFK3hB/Eq3PT5sQLPSX7wGKPPl
G3eJlPKrFI6FZNNscMmAN2FqUEjRaa3C0UpCuf0xpB74eyLH3WFbUlP/eTt4wp7V
LkLD1EQPmhoBwjI3j2NjxA9Fk02jfgOM/byHRtLE6x4eQB2lpqwaGs7JxhAN41BA
7JhGQoVnErPm4slmJ7hO874abqPLipFwz8E+cYoYkAo/LkIUE2c+7ZxFLQo94oAk
z09eiZXLlQWAlFbeIp9aYnZuYv8KvC9u9SVJHIWcaePWD0QgvVTRMt7lX8KyabXi
1xuD7mnO+YIVCNuJe+WvVMXcazDxuKOBb2WywHou1nB7z5A1mF9+5lZ8fp42G72M
+BzLSx8yv4i09hqJGa2zZWoX7VX19HuZ5PE13pPQ9wS+s9Ixvhh6D8iUz3NTb9CV
UyroUgllyEfzD1BjQZeu7/Y1Y3Gt46lP39NUZFFTxaagpRqHf2GbcBBMeTMxCLgq
FBBJnZApdOlYaFLq248q4aPVi7rdtR3JzJ+2fTm7uCU+GD2A7oVjgDeEHdC/h4xt
3qZn77O/iRNNYEHElM8JvDWMbY8iDEYa58YHqRRozYCv/ucy5nhkKZTKFwIRJudp
r86lPGY8U+5YdeH5puXHby8wrEz5stSbAoM8DdDP/SzVZHAyaSbE5vwi7az9ChZv
wJ1BNhuZZfgVuBHMBQ6gPqaSbrURnX1jykGhk91Zpdly6kgWlTyeeqhl120s7dol
T5P3rZeCPpfXefepNCuP2DPcJ0tnzGyCsOvLD5BFFzMqmrDVN4Q8K03slbc0FQ6j
k/1p1bh8ubt1bwx/6Nc8xjAUkfXrlFnYqf/YcJEEWWoiEmFzWqEm3XedrrEqqqUk
dlZM2N3v36yS503tsI2ezl3BJEZ1y7LeZUzWAF6H+e9EGrIZpZ83yMXda0pQEvR3
vV9SsxprcXjEYyT2K0gDiBMju+lCsx4uBZ9xylIamPwlTzVWTh24zLzW9sPuiZCL
vj0h77P5z3bF4jGO6Sw6ilSjBwTqGN2ZUChuw1z5fGw1erc0sqn2hidhgZ/THTcI
jphu1PmMXIiRKKoQ3poMdMYAtBChZ7FdDGlInc/krLBSbBogfCBPw2RNHE9eP4GM
EEMcaBhJgO36IRm7GYZ8E58f504cjZCS9xpPvKxfqt03yGSsPJzHKAPQ2pp0edd3
XtC362dDe6d3cwoZHokTKqjkb3J8OxCLF0GGI1Kx9rV4XknOa7wL+55pBXlE9lE/
rXjX2IaVslNaPmCu6iiLYlN5C17Nc6Ax3NXNj+ouYjbFdJOEaMJPXj9+cADX9pTJ
GK/C/7zvtoH+Mm3qLdmmxWB4K6nbQHmOtJUgAJ4FfZQQ565vuxdvdDVTYf/aB08q
SKl94oxAxBdiaJtCdLtd/NJRQR7uuEcRP6j4KsnQ+IBfOxZAwQTPtsZYq3WN/U33
pnQzqbT2tkvSHydR+XZafvFgx8ZtjyTzTHf3wMgxtNeOCLbwUTrVZW6/XChPodjX
K40GviTDYyAObV1Zgnm+CXKrTRyzjzO/Txm6sNgyJeYEMOhJdIFmheQl9lV6Iu2K
MKup+l9ZTCVv8hsaK1PK8TBkBDepFjNtOjUiKbLhmPIYfI2kS2Ttx+M04ZMPe224
vWYx6UzrKR2+vPyTW2DwuW7oj4eS6/x3Cp3pCfhjj1eWo3gF8L7ZrNUUldzsXgkM
4AVuLW3rkhpfgroL0w2G/TjL1NjxChHPArdIfk1z6ZlRB5o3Atl8mvsKHntLvabX
Xyv89ds3UJxGQmqOvaBfhJh3+JU+un4uSQuwUQVu3UglsknfXlrOq1miYAHpHpS2
ybrYXPk2cvDuVXGu8NeHa+JM/7lsBKl25C1GLXWIdya9n5/KaPYOaXSDRMIHZWZ6
pQ5me1dHim/Pzco7tg8vn6szsI8FNrP7eH6HOVo8nns+5lSR8odCh37UP2rLypv9
5KYYgYf1Xk9gesIKRMXPQ9NEoHQBr55Mth6rzIwVNNBB3rVn87P7YZGfgjYDAp7h
cEKoog+pW7WkUBkHvrPh0PHk17i+z1j6ddKajzGsJOjqUovzcaenNxT/Qt80zQr7
hoWTTpqZ84hFKiyWBC1CNC1Vscasyz2zwAahsl4zgtjH2iWah1vZL5VNJyBECGUQ
/eysO+lRuwcbN52/4ScLn76VS00NWO0OF0Y4BwFtNAe/J1wUWA87Nyz+ZzswmnYD
Z8GnwlttuWdB3ADQO0CF750oCrEjPq7NTLz4E8hph2r+9sL876COZLPrTpA/LH5r
mkaLJfsqnA21ubvIRf6dtHCtwS6fcaLPLOOmm3RxfXsTwltMeU6/Ap5MpJ0daSg7
zyY9juJdIHr+m3Mx5cW3Wp3RIorczSOuw/BkWcZIJgjT5r5+OzyL2zrbDH7+m8uc
O3E4z8Gzr7fD7jqLLHEQ/woLvIurlwhWqcV7LU1fNLNW6PBAkCbulg2XdJjU5vzN
5W4wQyYIX/e+o1IQ476YxwqcDwukRo7L5Qxk3rxSF+6FNPqGAUz7d0K1CIUAjgUh
GPznWzJlb7o29dqhde0/65cibDxUxHSHFxQKSqW5WLqtr8MsCkWlrhPZrPqaMixg
WO5K6rSQa/lfB6y9De3pokm0zaM9vww+gz4q/ZlBHaTCw7b+2s+FvE6mmfFATz3n
04bttvKtP6fp+1zBP8QvY9ToFnY7G6r1CGe1JU8tpFN54Ijrh/cu1rGFbb2lVp1Q
8YPdsVNQ7KqFAzPVS6igetBzCn+VOJWsLuoGh92+XIUGGLkLYz2Borg3vVSc9XuN
nzkal+RjLINihvcF2H+h2H6UtRw7nLaetJzxsf4FlT+FBJRXZdWQIjxeLtcVJnsl
Qmxr21vxnZBaeYqyh0EHfZYRgOpwKrsGWV38srgUD+zPoDheWAVB7aRw7sUZqvd7
hZ7Q7ifkvxpYGEQgERK0C44KzGPx780RDDu9+QV6NmBR4vguU/wlGrvdNRqA64HU
CV3CfXm90ri1gww8mHRZNsbQAKtFnCc5HVRUD0tJkBsM5H3/AzStAaNxiPnAtdu1
XJFAlpRJxXhjvgrrMeSc2cHqPjOAejSaEDpL6hsBSa/N2jVG2d/CQjScsY2u5Dp2
1ZcMmWUWLnQYXbswEpBUzqlhAlOQEfVY0ipCsZclBwzWp4CpWVDj/28ctGz4hrge
tpKTl1jxMt99K5p6yKEad1ZOKGqxUwM/D+/vPaMY4EMkhLrL9g8PEYattDu6USAo
gLBSHeJ+dVphX2TME0mnKR8PExwdhNdPNWvOynpYWTiIAz9WpC9ScEyujcyccP40
9g24YM9eZSEqVikW0Ucquwu49jkW9EoiSaKmmMq8DEk3Cv8M2dPVtjycEaKwBnYD
U14zoilsgKQNzQBAKo2ufJlVnHicrCSUkTsmso/VOn/YEzXD/hCsZejAKq5dBUrM
k8esMWI/ny3CiZcYBMLcYA7DdH7ixL7+T3c3BZbNkA0LFzNboS+Xcb8x36tg6wSi
NVYfQ+yqJGtqL5t+DDwycYasYyYEepjAD4VIGPLayZXpAcGExBsvo7Ix685kAmKU
j9ZE5eG9iS5PctoMRynPB/kQ6fhtr6cnk27JyGXNUB7yDZqHBJ+dm/PGP9jdWt7R
Xckt42babuIF4wP0X16skcbOwL7/UQ7pmqDgkIxNfhFS9tAGVYDZRn7T7zOvxEIc
AekM4jyPyB8B0I616F3FNU3vFlQvwn/Qd6erKJBcNIQAEMnS1jkTXbgW57MrsOJ3
Bj/mXmKLn/2Gc2e3XDDXH0SRd0WB5YRItO5s18nfz0dlKABD5hjFCEq1vNvkDPG6
gLqIXS3tkbajRLbd+YMYMACAqBEWeiArjO3P7WgnUMtcSPf17a66TMggC+x5BXDn
ctDoneQQe4wdzVD+tMCWBKe/S/MNIJ+BAVc7z6lPC2JEgEnPDLOcXvmRbKB8nJDv
1BthJ0uaT9r+TSfbsUEzqfpSI8EEcKlbd9WLgxAH4OJ78/0F/zMfV2JNpiQLbzX/
yco1527V4EC0MGjPoBH3RTPxjawjUKqJj/lga2UJ8Ljkkh4/Kus5DdzZMvFao8IS
kc0sQJ91MN9TUSZkCdwH+2/R3KLNaJiwfvNXtcaYLcCkebtTMzByA5syQMUzkhir
sjz3KhDT+K+sphUuTIUizgKv6jdrO1vDwKCdPCKE2sfx/3ZW8nYHi2mQ+1N0OEVT
xFpD/4XKw5xsL6jjNThXvNZ2O4HvswMfShOeoYWwt61MyEziJaCkmr5sSUWzqNd9
h7MLosDqASDJ7D8hoTFd5Z9+z5JrI1sXxK+JkSOTBAeo9A9o40GZPibKSrVS5ysr
iLmZJZewUCN1U8FHl7KYQsHM13HtpMkZwXnCAButpNrYOl8FRfM8BzDTlYmBuXj0
c2bpjnFvwiWqftLF82KHEMSnXp1z/5IcKnmKJhtrXIBi1KcuZV90trXmBtJ5OTWS
o/qwUeSFVGom0ZOmTHHf7n13HeyqWAT/Dtl5kCTv6eTbYHfqFTs4Nyyya0rBLtP2
sC6vrja/i6PY98JDaBgUH3MkiO/kWRWWMSw0J476LJkdBVtwf99bzBLv7mNl+VaP
6jPew1pYszCuS9M3MsAgyu8TZ4ukC6feuw2KtPkv1nE+yTJhaDDaiRvgSuy4qCuF
9rGTFrxpB/U6uEjhPqT7eTq7U5MNHA8mafc3KJBlwSoSDsP1FBl3Oc85annfYpJn
FnBdLSGx2reD93J7BMGy2qPuz8B8/NyYGjZzsR4iGzSg8FQehNKqLnOTPft7vRwv
arUMM6GmYq6X3Z/2Pr3wTCJgGfkbIPaVYObdM8kWFXt8FtyN82+bLkav1JLRjWFM
1ZGkt7YmUzq1+axEt/ZnGO/cYvP41kiGmXsVxzEXpclWD7IBIfc6cOa1SDVLKQGb
+PVdvBq8mwaVdVFGOgcdQT/0E9qh2AvsDdb/GEzedDy5lncEO0KByaJ4UXg0eQlT
koMRCo8h6/kM0OYsJgxMsgvQsXguwwHDFBrzQduTvhKQFCtClsQFVbgLne9WIZE3
KZEtZ6QR2PbNcKtJeXeI3M9tO9x6V2uyVrBytZhyybr6leYuho5olSPLhiprPQw/
k15TdB9Z1poD1pDgCYI+T0AUlmIEo9SO5vx6hBxQmRh6mB1KA0xlCoQzu8p9q1g1
BD22nR1A40uT2iDs5iq5sdxuBs5Z5naoU2jVsyQsIwkmox9E8MpOPaL5P/TIE9G4
gYe2wXmIOST1MKyil1PyW5I8n3giW0P6nQHpWGXkI2YVFZLZu3Zsb2SuLY2kiRTn
UOwS6+fVxX+kYiRhbhd4WOUDqxeo9QkWj5Bmk1V95RVHJmV6jjzIGcrv6BnMIk0b
MGfyAqq/DEbLn58AT2iy1nwGt1yc0zHLSVniR4c9H5mPLlcMMu4S/vaSGbLDbbZW
8PnTD7oDOh75J7D9nGpHcFKAOfaUFM9hjIXpMyKgQJ3irCm9drGL7ylW30SyQYLO
6Nlz1cBZ1CFdz670WzCOlFqAr5VAIEYruHFz7oy7zYFEgGx9etGpfAOkoMoPGOFg
WKWXf7YmEsFDHboRwTubVClZZ54ufFDAeh9I2GTlSxftF2daXGGtKIuErum79ouK
P0rOZ7LDAMD3V+uDgQTn7wCNHFPyqI57TFA/9TZ4+V4m3WPkukJ/BLK6pe7OOoVA
q7FyT8RnKHTM3Q3MSs/NgnZCmGAc/NBAwq4o7vnIwfeUXDpBn4Wre58dzKPQxLoM
yS9qaeTqHvmHh19XAlWD6fbmQOFSZ+1c+bjFPQF7raNTZYZiI0EDWusjxGj7vdxl
us7GMvxR3kISEMN1/jHpSPzIcJ/r6B4sP8Qwy+nkjogkksxhai5T/pKV6VKoY+UB
jiMURdVUGD8lr7sJLi1FG52z5O3mFTfMAwtgVNXWj2fGgpPUf6Sr9X2wq30RXVuj
8WItWByZLbEpinHT7nkIHn2t16/b0oegv5GfFEETfzihc0Yyy4JQnMkU3I4AmJ1O
33BZQ+I4IfWmW8Ttv+tyc1omDWUJNx052cH8y0yzSx1tXA7vAIrV+0n45tmNi7z4
SpX/IxqTVT2lUkOmg0ISepe0OLrrW/MtHwlq9qQhjdBcylQwpYieIsNkqGcXYSEW
iGybGo+4XAzDMDNJkcAt0pvi5NRYZH0MfDTN8yL2lmSKwhI5HPp4/24AESxiTZzV
pPI1PRdNyb0IO4h26vwN8EF1tkcLUZDn/xL0NdniCZWnFwkE91Q2ZkvWN8VhpjB1
3F7HMfx2ewsN2Z3/befVPtE1NQlcgs7wcksvu6cC/jl0g0XVUkDK6MgQM5JcqrMW
db0hgR6/6VdnB0LphpjyGuyBCh+mSq26n1r8Ca0iZ8iUWjzD+z8mmiGK0aW24yGw
Pcx+Ecb8+KzEjhCsp1+YAQH7nu8Ccf9ZbQ9lo6+WATNw07YjzbBeEMeLHi8pheGP
EjEetbSIgDBJwmvQU5uduNzNEBj6Kn0YVBm2yhK3uX69+Uo1pTuFUDyeUcgkdFf/
fTcVxQlQ88yBoGFubKxbmb/o6C3p4gEBpD1Tklku1xx/Oyytz1mTxtCR1pkWYCri
VU40bCc/5yJyca7/OD9uCSUVefH0Ww+8Vi17pqkZ5HfhoN+8NJedrhTYP1AsiUva
ytuCeIIBi8Ox+O0tdCaRwIGjipXZ/05fH7JhywHGIb+EAhvI2rHukMJ1vkpAzMAz
ZlkOF8jRvazNrZZhCVb0nn6gksqG9pKVQUJyKisdClhTa5B+DKcvN87hD/kgqIfp
/2QD9GFxtiMI+J3l5xhGJtRlwgH//8kmZ7SXSa4jkKkNh7OpXqvxIyij+1OKlpno
yRioiAnUOyDfGxhXtJTNsQLkf9zazdR2DvA4j2y1xoTjmtfbXggbYgmGLPk1VIR6
13WGJC67cXojbs3nmtLBqgqW7Y+uGFhKc4T1ys0w2vx/0xp7LRwCXH/19NAZDLlC
27CQ31TNGGN6BCfhi2uF/H1pR2sfYqJ0/J1tHkILodLNjmqA0vgzsQiWZ1bneA5p
JwVquY5gNrvw2c2tOsuFTXoMIbBmCNpT10MSxaD5dwKeDv8ZkFd0bwofiW1ocSAO
r0vKxtANhjaGCsz92N9yD34r3GnoKu5hMWsBs/umyshwv/G2fnT/A2heutiAXFUK
LC/QPRwZSMXC0P4Y2b5bKLGo5P7zjY+u5EXl59upiI6pOEEk+Q0QRbRnTnq5sSNv
ibslDe9OtQOzR9QfT0HFDlc24RlWQzKvY0o1o9+/aqDdSZl3O4RO0EOvuMzdlDiG
y2TLznuHAXuo6EJUzktBJD/P9KblW+L1IYnoog0YR+j4Ep7OoubH28BmxM2wEYNp
np6O14dOPpblUAoi3Br39/D/elTZmoeaR0/fyYuWmRCawwhHZ4okddQcIIqqwGfR
4lZ375IfvN+9Hn/M4B2VOdCJ/m/S/kf1ffyJ/2/yK0S6VGac9PX2HjJpyxX0jq5c
p8uRVIdXlEKsfhDLaEOnhnxZV0dBhCA7/11eHBZBEi55+Gsiss+829+W5gZPUKuv
/feJii7rD0McJKvMO+tBAjQ89sGN9IDaX9H1bmdqDI1ezWK+K4cwMEHNRKmz6Ndc
XQbfAyQgDQrD9lrEG/4lvmaLKImuhE1ujOB+fn+w3xScV37z9//xBg2wFnIuEIyo
lxGrpjFn0iDyOU79nvQshgmMTlJ3lxy6mHaj0Krtw+SfQrDHRKIoo2bj0423idOc
tzJmH4akTJPawo7I9c8O5WH7ASNpE8tTAH4tOB4UMrNa+Ih50qVFpbMT5P1wZgoM
Td6FiUROprdJnnqG9iqnOET35RKucQXyUk4vhe1BCUvXKQXJViHnTtsMre7z+/fi
NOTKpZkw75MvQg3UxHGJjzX0Vje/qXbFcW+n6wDj/x3eC1wpiLsVmXm/a6Bud75Y
7JPk4aoLdMME6iNHrbk/D/cLVcThTFaeTPuh0vC73Zmk1/hee6xFa81dLKK2hVut
8baquHXtv35OKbCfsL1YJt3IoBblxN5p9WJox5gxRPk6BqtBHy8eOjME+Ts0p3HO
zAVaBGQMIHF3PCv6IuckxYO/TK309B4j7Hco5gLCc+J6TAvjwmS91b3v83nUw1LN
zw9AuWsxEb7qUC80t/AIj67DCK6x5+123fhaGYn0f/3PYP5PaFjJOGzKvqiCiJ/W
o7EL832DyLOEkadm6iM2relEAMinQE6f5PUP7ksC9nfbr65q5eMf4kgozLAY1yAS
Hg5AHNn3ABzJu6W3tRmPRMziFiXVBYx4YSap49yfV4UzkVxZr543TmJ9nNmrJdNd
xYxCfoCBs1FwIffx9qpKpr3cFdZjszSQOHnszbxjxmjAfOkYyydku9LSDfU8nevA
eQYe/0uYazpT8XEA/ITTNgAlMuqwwVuDJl1EuDalWwVpmbtRBlSEIm1uuO3BQiUx
HdsoIgC6HjeiWR0yx5GQcNAKYazroJKqs1N68d9pAxZJGxmCryp9TK5iB0byw6Bw
W0BZUfvwUGaGGp5rPHw7n0+55wlZ89GkJ2sMjQ/8UT69bx3nEyjAiPpWfjH+PmvV
A74pqB5VwSwxnP2czrwpbJwjnon1TKlhAWwHGATeF3UKZFhBYV4ZJS8gBMXPh5Ir
lQ3hpLmA+FsWmRbD8IHpTxkwwigWmXJNTKqyNkmzUpPsIGOWJtRD3CsX97ffVwYA
6mM4scMiMdO/j1XeIA+mz4biZ7+Epml0TcQsHrRlFyTF2RVxnmJkOhja9OWcXAPa
jN+0DgONpPqwd85pymyXnfy12+05Wm4hW59M/JTU1SwBbsCO76xlmud3os1OR+7m
7Ucs3vM4O0by5MaK/wz8DE//LJiH5IGefb/dSIHIIV3wIs9sVJeNqz90MnWFSyOa
w9YbD/TIEytUHbR33XtXup+4UcUKU+aoY5aZ7QolahfttZTaWaGDvxRpupjbcBOL
JXEB1ORNs5zCqj+CanRf7C+IdDFYNjtZnor1D71m2udf5iP9TDMLzNI17WppUspF
IgEIH7gV5qCD0j1xYQFcNvYHt1U5GzoEhZ8DoXJTn/ei8M9hIW+/SUpFPXj+fUR/
SSomvy3hM9y0os0MswiH1WoBmcv4z2E7aVaNaYIwGesZE5VRPdHky79DnipDoTFp
IKdqINFHPRX9DHiq3NowrfdayvKCWbIjx6dW9S6NTNwB7Z6lfkdKvzyT2E9GA/4A
WsW1u7VTrqGbrXxyeJMcsQcsKYaNp9Yk82WZVvHlY1uOvCBY8ey+prE5Q9KGJ7Ng
N3XOqfuPx/D6kmQ9tZEkt15NYdViry03UlhgRSGLAkkbsPsQrmG/vo+bsWsLP0hX
OczmqkQ25SJKpzscOe6FFAYv9uLftpYmvTlfuV26SgP/XgWOzuICEHnWZgjSG+M7
AGojbQNRcSLtafNjuoKQCh3yOgol8PB+IO8kZCHvl66lDFXcxON7JmNg94zmk9D7
pN4WxIlqcQ3c+PQVbYgHhXIaUHadeYdYQwgbFoWKpdex5q4pkLJzQco+YsWVVWxB
akGCc/m2mWEseh/mlOIWMKGi1T42NjySmK5fwdqnHu4YB7cbFPNDTnaGPMB6303Y
jZXkeJF+IrTrBRNTOlVr+OSfj9XO13xYzrqa5lvH/9ZYV+Ohiyz8hNYxbJBpxGvk
OL3zOpktcoGx/ZDKdbx6Vn7q+1VrMjHQGh1b86cm9LqHX1+6Mpszuxqn7aOfy9gb
o5fATIhl7/CC+E/PSbdGHQtWTN5pnq6NvFCCMMEsAK0pFLUWUKYBA/XtbBFvE8qz
4pw78mS2DH9Z2Ia/WTJ8nWqISpzE5P2cAuOsQ5BG2ZRPxtoWpl4qKTKDfMAeuY6j
16G0kcc92BGkvivm7lCqCLgBbKhxvwVtVXbMiTjlBW2puKVSE2C7mXsued9lJCkd
jfiwfRN6SfSc1tgZ+sF5VpBCGJEeHHCySCF17Ob6K0QlZBHvkuwlkZLQDrQY2QbL
OfQ9r2a0YD1gxNChNxoDaBONeSr3RPa3J8wNUW0doUoAVqAGH3lMs35nujawjozN
KHOXs0LjcH3pM0lIHo8t9MMpPOhqI6RgkcpYLSnXvbO405JDjBgNbz9r/BnE165T
aS3ZEPKsyTFIBWhQUhzFR/iPR16hR+BzPJq/r9bFQ38IJuXdSbj2axiGJnegFSWZ
5byRRM2x8l7nnM3Zf87l+je44gC38cU/GNoyXsIRtQEnaI58VZIAKKJSzvoXBF0O
jhtMYoxHoPTyBI73R4utInc0DWuFxABhV/H2cTK5yP78QNTqTyBADu3W9m1GHpwl
VTgSxo0ROeWjpJqnCWRx0k4U/XhxyTmKUK5v5oKV1JkVS13dyH6um5ciTLPLZL4y
`pragma protect end_protected
