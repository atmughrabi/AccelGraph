// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LbjYgd3KQ48lO4ccyKbDW/9ErF4g7NyfIVWME0zfDGN5HOHtAFdpf32UOlzGRn03
r8CPxaWRhiTM4x/3KD1toI4OKj52FUalT3dx9kzVDEkXHw30erUJywIOlUaNOxvC
DZ1ND28lbGR2M3liXqDriuRxn+cOLfFIA6AYK4oKO34=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5408)
YuhaUZ1lJXIkMvWcIp0Pwdn7NTd8NqlvyDN9XkNbhsB3/gl27Arxsuvk9HO5TAR2
DPJfrBbeHbIggs8jDAFRNlfNdG8qFpgwXxTbvskEnm1x5Lf0TOz1MlWdgjP9Mifd
NxEEBLQvMANm19Ze84GPN97erCg3IvXiYG1rNWatlZ6AQU6lRnlODV6+n1hL2p6S
fwqIQGVofOp1qR4smaoHsnRyuP4vNNxvsFMfqRAKWvyym+6XNEAMQkQy1cOokrQJ
agFW9XLiaWuGCngsx3r4HHjWnpkkhZr0AK2n8wTj8pN3BP1RsXlQh9J0LKJRObPu
afAzzl2sprsZNvcVU1gi+JzscMIJoGFvr5elmOp1AgELnLIg2BIOu16/O053AlOY
cld1mmx1j7tM7sdTVGNpoxEHS2DQJZ4KPtWCqAYMRW3JHZD6IuI2kGH8BzxsIDa6
Jc164ExlaG2Ew+uXw1ciOKliPyOlesr6odyocX5F/wxD6krpQOgt9Mfvz1AbBoF0
uE+ap7Aj62aeHSTEC4Ho8UTjxwMvmGA5eCe6H8xIPue2zGOxoamsP7tA0mWeDYJe
Hf+4hFyhGjYZ0T9AJXWpS8z0TsIeeKVd8s4vTVlnfcd2sTvEjb29RqPENrXgFhqN
CUI5jlb6o1s3QT3aiXDvGFc00gQ7LMKhNs43o9pAUAbhS4kGTDBHfcv6f+1WmIB7
DkGs8kf2c2Z2nCa5t0esp2VWYNbyYEkh6LQScrT9ZA+QWSJAx0oQYafezp00pbXM
8fTq66hloRyHNo24gdrKtdma0xE5wc5SCRxMUNmZRUDv/3no5CvzMcU19FABY4Sd
kAEb9dCCjGQbmPf9OkK9pcKqBodowTwpxfX4cw94M5iuLHKsECgeEunFYFLBvl9W
JP0m/9R0Cd/muOVxFE7eLnogabsOnyKAhEFcFe3VImmOeiiHWqMl+1hiwGpfA9rY
38iD4zzIbtDdWXNWTQjFgvrS+lm7CGHipksplcWynKOMp3nYuMMLnnlOCzveoSAO
fLddWXT6BOntUZhCbJFi6IqDciL/0AvkKBcxbPTyL0PCMI1utWPOtjs98h2IDQTd
YUliyBzTPuxh0VjhSDdZ01GyDP3hHcwCdNcDfmkRC+jcUDrJjHtguLQrsvQtoILy
OiFQhFXXomman818C7R/Uxvw7w3SNr3SuMM/gw9sUt8T89GEbWLSpnjLNF3GginI
M4potOqTO/cSYEfHbWox9RhlUQrp0qRNdBPwHUhXOqNiNRFimAQYUEgCjDIzHYkv
tDejFrZqMByFKF2ytVCTTV0FwXgHbuoDPuzxrLzADkenrQt+Y8YsnmbxZ5w7cjuE
H8LQie7SK04TyfDEosrPyUEpIvbwIvN6Of9er9rAAxrxClkfJDa6FR4HzET85YaX
/yvvnlHkKNo0a1GVx9TrvOuL/38dgQo2KlMdBQyVzxEuc/MmMLv/CjiQLvyOslJc
mx1FJ/c/s5ADvGwlYGJHd4ZbDJkrXYYEsrw2I6XoQHXKzw3VCthIR/JvyI4+RKG9
8Kbn4hbCfhfWzaBYC8FrFtj2pzJMwmzSLQntaaKFE3J4bhyLfBeKigG2aht2REUS
y5fltaoHhlVDNehU76fOCge7ISgK1ZysOoAjm65V9cLJYpa+Mb6vKs+Ex8bI0Zu7
UaEboysYfNCit8+fExM6TT74M8trY40Wr9ORPh64AUOVCCqZiwD66x2VMwzyDW+A
H7+euqw+cF7wkKPBytVST9JAnbfPe+K80mgUhUFYvO7+7ispc0vSoM9ziE4G6ANO
QlBaKQe0fHmaCAfmaWEiCpIJ9JBqGG0ukaK6hsqfW2IvNF3h8yeNl3nP5//msplP
7gH9DNYFYNZe1DkDFXy9iB9/qjvpcwM+1goJyIvfppIWYT8QpdTZ2hnReRGai1XQ
KKQ8cjXCcodlr3GP+eH/EvtpiNqRrzY5kiVUAD3zNrTsUnKQrcieFaaSCHr0uyMp
dduif9clOp48JgriYX++an6argHtWKVw0lk+YolGNy6EhpqlCMh5uOpWSs2NSAM6
ey0mP0t2Rfdg6cgU67rxhoWDS9Va1UnAJ9ClSVmKLrNg7kUe/wlJOvZLIsuLZNxr
gKaBTXfsotpWxrdtcqpOVWHtGAGSVFl9oS2qMuJ6TrnPsHQN6sZd0I3qDb1xA9ib
h/RfOaBpXBD5xEwQ6txdy6o1xHfBemneCtlSDa+9CWmak1kPaW+vEEYtjCUrOx7Z
sAYAZ1SJ4NvUs+bY1KE3KEPoEyIWZwxIzhDrTvK1U3TxSwjC2/PO3v4vC74EHedM
r34A/Q4JxOj9BQv1mtBk6PobMFTzEs8Rv2s0fhN2J6ojuK1oMvJISHiMTmI7KJNj
+DBNXcr5PHv9fVaDLhnMPxjgmWuCnTRJiOybyZyco4LD6uHwYk2uzLBXwcxsZv3z
1C8icRJe9SK2gzFrIoktujRsfwBB4QaAgRnYxrV3RopKz3qPZ/BFFt4329s76CN/
w73hwPvOeCDHT0zGkDPHARktXE9EyLS8GClrQ8JmfiEJsir8p25HwPqzUkt/213o
ojYPFH/2l+1Fpr/XrPnn6uQ+u5HUG+3Z09qzzxyqvsTl5WYEWIQlNIRseqzkzgvd
ezfhzZrQq11KbnFvHEyszQ3aZtsrSIyAw0ErNPLUjZgc79VodpPTDLCKRmmmUUg7
LODg7U8bzhDjDLCRrh7xEJLV8phF0dlFL9AgomIyOX2qSXQULmTp8j0xwQAyuXms
9bezMyawDnnMgfdCwZQNt1g+0REOYbM7eoFKA2nrigyAnIT7V0AlkvcCl1kBNjrL
du4ooGF5VHWDIqlwPySqH9E7KED2+GtRPCtftqgKoJ/HDlrPmuCmde08FoHy+2fc
UWGp8kpwDZN70vO3tc7m2GJUdiZhDqzYcTLpG5JvnVgAl+gXJBd1m0Rgc+m/4Czq
JLsbpzf/9z9AqQRJWMelI7vDmebWuFgpRiG4W9TvcnzIpxa6OfeI2DPyfjdP5Oba
cmca8TAvWNl3rk85pVXYz9ipIuMRA0PiR95dfLLgU4TQ3uaDoAqobM5FeS2fJaxc
a5IkztQjOZqX0LMGS/CkrRhsy+yiMNN13/+jCvDlmoHhsW3QCVS+jto+cq0dW6mZ
fw9xW81pN3R6J2yoq7cph3SWTur9RZV404ZdpUHNJ6N/47K/7HNH4ChicAo3X7Bt
Xwk6RDdy3nrTza9ES+ciYH7Eu0z1pbsvPg7DLJyk1f/XNvxmPKYCu10tlSvoslHO
H1lg3QrcdDgEZ1WRlQNtdoilKf1bEESuoldr4ZFtD6rOZo7g8e5u9F8/iABCTzld
tL8T/FlG+GNdi/vFGvH5hfXWtZhM6v6IkZQ+ga2OyysNtYcf44uWTspf7xWK+esL
/mCQa5X62IiB2PD31PXUNgr/kq5KvQZ1s4XIFoes2brDCwOs0JRPLOKy110hc3sm
qqF2IqyLiXGaazr8aiClC7xrfmG1nkNjJSjajtR9y2slx1bJu7gD1DoQzelGck07
CCl6slRH/rK0v/BfxDofHXaJHucqXIbj6Mv11JBDXHkh9RQ/NpRof3pegzq8keCL
IR/ueaUf9iVVRkmbCsVYLdtXG53ADI+wmbXaSUx55wgCL74CAySM1GiyIlSDG5Bs
QFx3K6vKi83dB2DRrp1qG86BWmxqobG/3zy+hTJpbnGc7TSN6FnOFwJPM/0cU1n9
8gIk5ZRrL47fQxGTAEFlR5Eicm6O1A0kifI3cNM65GaAcNb/kHcxbep6jxp378HB
CJ0+nZuVCrhc5rIn98CWzS21FsNIaLP0nHocLv0fp5otKkfu7d2ldLZwOZAw5J9M
1B6Op+QoWeZIKoG2wb0CNYKAQ7+cxXHwm4yuebwINe+5rdSyO93kgaPLRR0ybiCx
OikRHtHmrcCFxzjWtdYvIPZEdG+tJC132d8k8JAf4hKLSEHkH0viAI3x61Sor8mi
Wnb7KbNYnvfTlrSs5f2h/x79pu9iNTEVnnVbn1QiRUFMV0TTA3VI6dl5XpJdhzqI
bk2oguwIZ2BV2sB8HxoNqGdMqz1h7M2JRlNqgK737mxETAx+raBuuNdZe4ct1zX9
uXgyR4f/DBMcmM3KU7JmYWYd5MJWOMS9WDZqDHP2SYf2+pYhtXZdKUcjDMqItpYu
VVVHIlXu660DgQjdSk3NTkLi9phZhvEhzlEjOMs/nvmAg4WeCfsIOa7OboyQWlcv
TSiZEJxPTSsOJ+WPvQevtaudEUstT7pE8oQO/zRB782XxiREjzjdbQ7z+I2eMT3h
dDgr6j0KEq2daPWTAGB0OUxLIkcNiXPYejK4Imzb7zGDcZXeBnpp7VU9SYk9qifK
tOw+CrSM8zWlxDFRThoyCScHeGQE3hMYCWzpz8gx4I/3tYx4fYcy0DIn1bcMGM7I
/1loHhC9+G1bwUhni+vj8aGQmyiRXuluU1dnungqKS13TcGjIx4M98LmKnSd9qAz
dex2QPi17Tu5fAZs4k+EX1yKfA4bOBUGqkLNvKl5GLMjuKMlFqVegw3Lv78vV6k4
Kl1rsQPKDnj06UasYkE2XSygJIR63m1RbhAbVX5CQdB3nOtucsKk4B6sTGkHU8BU
21YGXJu0L5v9sf9NjN6EP3g7BGxyfz+0y2jhVVAnQLsPqAVI6tElrl9AUzb47Agt
9edOyhMwKoWTLm8R1Lhb/IyIcf2gXAZAr5Ctfih8Cg7n/u/on7F53nRUJ1vB5Wcr
ve8s96vNlGGsY4RFKxz85vBD0/0pZud5CWJ1x6YdgaR3tF2DHi+4N9GlR/ugLQhF
wolpN76LYRbvYBqZYx9tZwINWTafz3iNu+SRLBDGM6QE2oi/N4N05aKCP4Pw4BrE
Ix810TSXaHGhb3iF5lkHKjKidaXsHWTKck5QBVle9asqaAX8SY3lXUqsG0GQcCai
IPZnKozIBcIX9CHrELioKik8Wn2gwmyXej/safiU4lYDkB3WAOxuHVin+EosO1J1
TeaN3cSM7nVRo4ZRXcF3tPuce1GtSgWbzLnlnVQyPbtY5GbF2L7ja6+XfYM258WE
qRGI0tYs/uj4N6co4pn7NDTWRGO0iU9AzkFTXB5HTvz+jTofkMR8Xem1qMK/o9OP
vekcq06okPr3dwLeiOdvJC63Fdc+bB5359YvLhrBC0uP/gndhitVBgMPP0txvOam
WJXFJU1p6wwQvP2S2Fr6u/1E4uFwjqF+B/v7ZqkdDHG+bJ+1aK0jh7wifNyRowZw
ElJ78ka0qojUYqlg/eOkb9NAEDbHmztrg4YUxvZ9fyn++ATY2Jw+vSKt1rP4S9x1
wCQaad0r/O5AqPX3BgVeFTl1kOK9goaeKzN0vdflbdVOjtMD9X7qsLosz2oW9RE+
HAgBvZ73rAsA4iLT5g2pQ0Lbt0PC6cXWMxE9vqAF/k/idp//Yv3oFabOav+Y9Lqx
ghVEbT7E/U3YHFE+mtwBIFZPOFY3ZvEXkUW43fEmt6HEvZncvR4XgOiDpF6g7KRt
d4ID3A0vKztp0NWTv1mRRL8AALueZ9rtfoDrCTVRWFPFyQ+U/6KWD/ViSE7TXC66
poLpWoItMdsuEggMRBE6BliJGWJvJfJhBV8aGtOQaik6aerCCbmYPEV/cbk51SGk
KDE5k3PVQ+AX2QELLJ7BjuOH/+YtDIQYw3JlI9bsGn0PrjV0nvwooKuTuuDkF9J/
rSsyKVC7sv5Bx+WfC5xyqa3iPnxZVtDZX6qgJCRAMkBnithbGmiXCNXpRdPNQyvl
ozPARa/9+XBeEhu9t6VsGKZikI3zgysRQIedjoE2OO4Cnoq7OCvEjDgAKkyIvLBQ
SbMKv4y7eI2UsAwAk5ZNIu8JpjxRxx1DchC0KKpSJcjlpDdl1cc/CmC/E1Wq6Kjk
4dah0djB8YAjYtkbiuFQlITmsHa7gPUolAVmZKoO8+LjI7dbLq7mVHuS/HXCcojY
KkHA58IM32uwYwvBiOi8DW2R2rE1xLTvlF8vu1hnS58PpJqZSbplbtFbhlkFXRWa
TDX4Kkf2SY7l/xSKA7M2oggYAZckDjTPZ9Bd1uBdL0flS+a165bjnplZsmhR5kMh
ppha1BgHcORQzOcLaOAaDiU+O76Xo+9gdrXINvmXfOJON9vyfZ4l+AdzpLtWNhmY
57zrHg7QDQg2ZJpq9ZqDCbgOucRnMdOcvmXrJ4aU3A6pTm1BSHEqn1EwUTetUYGC
o/sT8Ae0Rrhp4nbrAw8KnO6XKVrlkiafTvMTc5X7qwvLIjhtVWNYsJq0bnF1PpRi
pIYu11IZAqm1pd2tCwC8wNH0XuBQD9NFWIe02p3Uz84f0TZ4D5mbjP+XCivcoPSc
sAP5vgoaAUL58EVoliXn5FBv87jqwDYo7JNwXI1tWCKT5so4M1LV9g7gtkhmXxsX
2+usOQ2fx373e67Fi9qivCpSMwLAUsMY2rUBGWRBO4+HPXA7MikzfWLU73vQV3tY
ViBn4g3e5klnXxCCqMdBzEIOqUlHxNfQMc9TxmdoeNFi6cW218bzKGA1UIpFpGlA
hq0+3S63Sy3ag2fch9wHXo/n3NVCPQofVV+nWeU7Hyrso0k8Mt0Mn/FvJ2ZS04sy
6DJ3JcDWtg+06pyIdw1aG9mtZcBNvM+wliLv411YFi2renqgTD1ZZiLHeipSWZY+
U81h03pJF8lc+SajWM60eU4I4a+kHxXbYJAbr9v0sq2aiybUIM481qDwxgmuEKYl
2o7ghxFp0X3OdDlEprDkWpneb6c6H0NG3aTFh/QiqRb0gUp/q1QE7LfCzIypWd4c
SV5/xS34NA2rTZWE0ltq9/bgsxxY1nIrhRFGLh1KiIsp58dYE8ENDDB6Z4DNYQv+
K3Z6WHivup4gaGKvtmwbBUbI+1uva5yytLR9bdi709TmM0qjJKIFQ9zjvDAKM/gj
sE+I0OnAcaBcNwimgBihlXP3cgE/dhqiGyxFaW3YulyymiZN+3W7KNLzfJbQZtTj
pWraqo5/XipMPkD20fqhBAAySjZ7GHnGdx9bE0FhzqYJcERnkIhPRZUYtEpOubPR
me0D11Cu9r5GhgG75WX7KQkDfjMKIyIl8ZL5jsdshIOuKm2Aeh7qG7HOi4+qp6sk
7ZfDvuH/38x0JJTnjndhB9iHn/jeCYby9RXWwW9Bs3ohZ3XfPoq3Cp3gkbL7MzED
+up+ubedmhodlpA2ySM7MWWgWLOXfVqK4dw0+6gM/pQ=
`pragma protect end_protected
