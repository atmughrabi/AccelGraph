��/  ����qy;�0��.,l�ٲ�U�@9bS��
N|B�f�	��#��0q��������!����#�K�f�,S�6G�а���'�~�!˰�Qy�XK�C��d}�, 7�sÐ�����d%2wԮ�����w�3��)$o�[����擜��Ԋ����H����#{@��)	�<�:3eE��He���#��� `�IY�ݖk�;;Y��Y��;Պ_��	�r�vmW7z�ö�%~�}=�S�3U"
]�/�
��
\@�;��`�(��f�y��.�V�ᝰ��dП4�]٫����WvTV���ׅ�8����m)|���j�%��^/��LH�|1P�e*��x�4i+�J�ȇ�! �r�.�ϲ���K��LN���{�l���r�.sM�%]po@�q`�h���+���B� 9���hu���v��B�)}\��+��ZB��q]![+�3�:r��^�>��Mh"�U��/]��~++J@F�������U�8PZO63���'d��T[� :+��0.��Vy���{9���~��Sc
�خ�~� iЭm;�Ri�l��.3�+��|BW�C:k�%���-SSF��Xn���9�����N��plG�g��l�;�$jL�#�s>�{� q|�
�����zI�MN��OJW���l��=?�G�5N�8�z��;�(��n��ܼ?ϝ�CrH�
����@ӱ�B�
:�����Of�f���T�)}�^[>���/>{��K�wr�`�=��I��m�親�|ȥ�4�p��P�M�|�����O����x�Q�y����1oaF�y�0ݒ:tn�'���2e���/H�k�H����Cń���&���F���6F'3�)���+6?�+Q�zl=GJ�ڭ����c�c	���"���ղ&I|�ǈ�	�,2�`�bƟ�d~���)���@\N"�Mr樯&�K5&.rW��f�S��<�~Q�Ӧ��1��+�t%�� �1�3�Ѕ��1�݆�	Ra����n +�+����۟A?�vR�9����v��~�eħ ĵx�53VG�e�5��ƏT�즓c�J��,#1F�{o���a����Xm~ ^^��,AA��Ŕv�§TǑ�R��֍�sȑ���Z��L)3)@P�,,њ�ٖ������B7�|�˂�~�Ԑ�iĩ8x�!������O-�A��6�g l) �	6��Zo��jF�p��C���p[D�^[�+���b�:����&�j��<=xa�I��O���j]��U���G7� ��#a��O�Gb9 ��b�p/7���]i��}�0Y �� =�S:��
>3����~}6!˕x�K@:襔@�yFg�Bwز��@&�`uX��s���=0Q���Ե�N�T"�2J~v,4=�2`�}gݩ��p����Aՠ�b�M����S��8E�2o�۴%q�F9��$z��
��'OBbC��Y���L�-��~_����oC�L�A+rbH@�`�q�aAӐ�¯�\��eumձx
�<�O��(6\b�}7���-�m	�l�{)=���Rs7H�'Rh9�V#d�)ʈf�� �n(��#�?v�S�zU��\����I���2�,��T�)��8�6���.�A������tz�Ɠ!Q7���:@9|�R���0�f9���a�����XE_�Ȅ�wyXn�5Zd;�؆�������^G-/�xJ[��N�vLIU��՗*��H��$r�N3����L��ed(ux�B����ۏ�64�K��'��_�(OU�(��e��_�2���>�kk����6<D<Qq\��#2� �E��AZNG��'��5V�L(\��V ��K�k;(~%�Vωd]83�3��Qv��W%h���L�@E����H*W{�X���N�vQ�m+pA�9�R|)�"�0��U�f#5�}j��g��淪�?Ci�`�k��}Vn�!��'T��Ne��;i��=@�/~�Ѧ=��]��)jiG^���-��7GI�X����L@�Y���2*°R�,R�/��⃦�L�YI�ݛƖo|Ô�E0��t�p'c�㹣�p�,�b/�8���>��-y���*����ʻ?��U�7E!�N��RY�� �y�%5�_��j"��DHW;]}�q�m��@%>�¡��g.x��mTG�C�
�\Z(�\O�kQ��G�(^�#3��C��!�+��L�L������;�v���,a �y���#XU<߸"u��ŉ�ѣc�0X���a���ߵEO�,��o� [)��$�+Y�f�J�*�<w�*������&���9���x��������P���Їm�mPH��M��JJ����B��c�g�!���e�����̬�L��q�}���Z�w�O�j��O�HV��M��u&.��
H�vx-k�ڸU�XU���z�V�?G:����D�2����z��MQ�W�!\��I����@_�>�e���fόj�X��K��x���ّ���5�8�ͬǑ(c=��i<r�i˖�����m	5QN�:�� ��c־d�m�۵��-'U��V��;��
y.����_K���M���ћ��@��fe( �����Pv��S�w�leͥ�f��d�ҁ�[�R��Z���܊�<���
X��|{_%	7B�)j��T�����L�Nd鎤H�R�+ aJӾ�\x��rL��)B��[$�P
��XRe�;-�ȰZ{��W���#�1z[�K�m"wH��MR*zmkU�S6�ұ21�v�`�ks�`��M���n?u�KS�= ������
�5n>*��F*]������#x��������>����+�R�v �0���V�ȓtX~���ۡ�OC3�1|;	.�wMBT{P�DW�!&0�?�ހ��GsR8i��phI���s�v����i П:	����4$�5wv"$�+�Æ8�9V�[8օ�?u�U'���Rh�d��d�i"ճ\x�����冹4Bj���m�:��L���{�7����Cۡ�LG&�H<�1�iSM��UqN�����4lW���e�R���9]Jj�kp9�}�W��	�w�dy��H|�ugS��.�F�V���w�<�r[�_�]녬���_?��Tw��t�{%� ��ؓ�6�vLQP]4���6�&!�F��5�M]"^�$�8��+�|x�SEO! �h��=�>Ε/fo��X�N�t@�#Z���0]��q���<�����%p�&Jp�F�Z�s�g��asg�n���6o�U�"|oCv��'F�ܙf'�)J�!.��CY�	�6����H<�=QO�4VU߬M�	�^��f��suD��
����	s�!�E,�H@Du�'O0ֱL�į;]�Ig������s�j�nH�����`6���酻�j��m�'ɢm}����F����h��{3�Z��l��>|v*�j<���kW�����KQXq�oR���rVq�k���\dT	#sq'�GDQ]?��m��%X*�+�!�5.:B�֪�,t[l�C�M���&�5Nߊ�	�$�T_}�Zkr�,~�mR����#����rDA�Y��:�����zW��itū^N����
�htw��; "�=Gz�v��fXξM]�O��l��᳿��4����8�MH�L&C�=��1��`�T�4�1�N
*��2]�n�h�T��eΔ7;F�-HD �<�Gv�)�s^���E~\WP��KA�`�{��ц��^�?��%�7V,A�n��[Q�?��Ps������n9���=|X����A��{7^
�&� X<����+	�8������d\��u��S�q��_�wY�\�습�p`��4�ڋ;������)"�"��*#����ĲNJ���C��Hu�"3ck��m������а�h�i�1�������Ȕ�O3�=�?���(gQd��90��)(<�5�.��Y�_���z���x�sPڢ�ӛK��b2�����@�%�}z��fB\uJ&L;� �-"OjE�8�|���+��p�)kdf�c�EQ���Ȼ�+t"��hCx�M���k����1{N��1��8��`�O̽I��}�~�|�Fa�\'9R�J����a����o/^7ۆ�ej�:GX�}y�T]�(�J�zj]{ϥ�g��<)
��y�� y�˘H�=v��FCp`6�D:��β��V�9� ���"{~`rg9�����g�uZ��X�P��?:��Y�!Dm��b�2�eU���)��|eK�i�^ ��U�<��D3Fj��T���	�xb5����H�!>#�Ǵ#�3�x%o�r1V��eG�� �2���K��ܒ5�oGQ���]s�f���q�J���z��ŗK戼�r��
������X\Qo������ߏ��_!�n��+I5��`�o4&�|�ћ��};�����]�w��"XwܔG��ut�����~��z�0l�)��V�Li���t�zxqyj-yo���% L�8���*���K v�J2�c�)�����������"����&�u�Fupl��p?9����#�d��;e~��wLS�x���{v����(�f>� i �}��G'��;�4��K�:�VQ@�A�u�[ҞT��и*�?��$,���c���[���mB�@��`*$�.��w��s{�I;g%�D)B�.�V�iF��dm��4�́�*adt�����Re ���������I�M�N��ݕ̡vLVczY]Z��B��X�2�[�y���skx�c	&��� h�k��1�E1�M��nI��C��-R��X������w���[vu�qA��LUR~�c�Q6T��7��`a#y(�_�K~L�ņ��@9O����������,�ȟ`-����փdЉ�uAn\q/��4�5���"5ݰ��P8�_�W��ҟu4�R���Nf��+�)p{��L�MH��Z��i�Ti�����8a�#��繳CI�m@X6z4TC���E��F�V)0C؎�F��Du[�zk�Iܭ�(���B)�7�Qd������5L����q6�#��Fy<-dGw���,5� o��^U>(�,529Q�rjVt}Pk̬gn�Y��j�潙���
|��SހIP�����g�'�t�ͭz�����KG6�=�§#���o�8��}`:�h6i:��[�����'Ge�-{���4W߃�~*�y:��"�b��~��i�v=��`�j0&�f��`z��&�	;�FΖȃԾq؋���h�����`��zx�tA
u�2㿊Kv�~�.I�m�.&��~h�q�=G&0@�5��ք'�S�I���;��oa͗�D�1�4�T�Ceej�o��ԋ���c\,]lY?�i���o���>`My�)0����ʎ�C��X�H��'v�_q��=��ϣ'��[n��O��Ӈ�����!�	�JU�5#��uLܶ�.�n����Pr�4�?7(uNa��扇�c$���-Q�JOWB��	k��.��C�3�zA��6Q�ǽ��Ln���a�p�k/�`6g	�pQ��-[N�X�6���x���t<&�X��^gMs�����ވ�;�?��y����^�p&|L##Ԁi�u��&� �&? 8a;#'=X���4�HL?V��WG �Im��J/ �K:���0��?GL$4!ԀgWUY��?� �����?��,^��Ǚf��;c2LA��B�n�D������-�R�l!A}����h���p� ]8�[\U�w͗1�̵8���Q{Q���� y &�oiG5bGU�<���%V���S!�&PK�/$���`֞������o�X�ځ�kO��Ts-����ް� _�C�@[�!����n*���A��IM=#�XX�>�xY�{��ڲ���@��4EJF, �:W#���!�e�(�A�<ٖ׶��O�}�>`'�a�QZᢛi �[¾vC%*>%��+�>���^��ٳ�U�~vm��c<k�Ѭ� -i,j�1�e7�Dƨ�{��|ͳok[̞��#B#����%ŝ�H��|X�@��Ĕ�(��/�rO�D���{��FO�|�.�e@m���u��L]bz�d�V�h�H��df�`���z������Ǧ���x��ǌ݇4B����'��'D�m��áZ�� �˨"�ߖ�Ǥ���ꌢD�61����X���	^P�)<Ö e���n���P&��T� ӛ�Z���;�nZ�N�d:��fV��P�+�ʰ����K��_�F*����sF^�ҝ%��k���`�a���C��n� 6�fW�l������R/Z8����dqH�A��m[f2�~�ToS�B����ͯ�>��OQY"-G�zZ��֭r�Ҽ���g�:���.�Z:1��������;"n��>�E@����Cû�ǳ�9+����f��SA��<����V���g�>�H����n��l83�-@z�^��Zy)��Zv�<Ψ:���Ƀ]	%[Ǫ��>%�I��=�D�ɀh'�2��᥉Î0P�-p��IZ�4v�H�	 FN���E?�P4��I���E�m��5e��x'��[�Hs���_�ﱘ�7%r[����N~ �����Gť�����J`���=S�O��ps�%��,^��@��Hv����0�0wr�@���f�ɛ�Hw?�����U=��ҬG�ϔ�:.� �:��K3�+,��8�3�~��t{/�+�i�S�S�����=��2I��G����r|jl2e!��5S��s�\fj��)y����K^^�kF!���	��
��#�G��"%_ac,���7Q�ɰ�+ſZ�9�x��IN�"�q)�L�����7.�oj܊n��m%��s���p=P�����1u]�
&?��$�}��1'�$�T�)��q���⭐�xe1w<%t����+.��2s�گ�����$�����v����|�^a��6�>���{J��n��2����G���܄i�aY�-��/)	l��8���{Y�K�'r,�/9��9x�:/b �.[U̔gM卓ϲ�� ��8J���� �t7��w�=�[i���a� D?��c����ۉ�-��]0oi�N{t����K�h'���~�$3l�\����*�;�����}��Z�4���4�#C��,w/n�.��E�/�: 6˽x��؎��`�X��}~��UH%�P/2	9z]Ϭ�0�{B����g'�Q�m�/� �>��>�"��ߐL�-����+8;��s%�T"�͑iM���	cZ��T?���̟�d*#�$���)2!2#�M$8�iop�ԇ�f��mM���#�n���,�a|%��"#E-�l�fP�g7M��<QfD��>BG���ġ;�iC�&"�A�-S��͌1��u@�wB^�GքW�j�p�"#�IJO����x3:�,8fUs���S����
]����@^��N�)Q4��-�����@���P-,,#fJ÷����X#$F{��}�Q�0s@�]8e���j\�����^g�D�H��P_
�4�G͗�������@����2Y@JC(#M�u_����+�=�����i&P��%^_��%�Ƿ��O�������F�`����2ŜV2�8�Ŗ����穁�"�����X#Uv���b���0�p��/�5�Ł�z#\C�;<�v��*�O:W:�����Y��߂�~_b�S+ye��u��3��p�O�i��+�g�S��y�d&��Һ�gH���h�P�t�못��IZ|=�mNo{W��x����5������#*/����ކI�.٢�Ԅ�ilm`�f�bI���&�������������q�p��׎��A����h�g��n���+��|�Ŝ-e3�؎!?�Y�M��af�o΀V�E�$��۩9��k�w�u��ת�9��j��x�K��:	��M�������k���]=��O�8���t���B�N�<�G+T�+�#�:~s�99���{>��N�#w����I�a���P(�*9(���ޫ���l��Bd#U���lT��J#�����,�昨�b���+�s7Y��\Z�F���S��n?5��K
}=:�����}M�~��W�W�Z����%�=,��0j3�;��@��4�Α���7�$����M�ݼ�՗���q{�-'�kS2|N m��&K���;��FU_��Bs]Q�K���� '"�A���x�y$ ����P�&8�-'�Lq��Hvc~G���K���٣y�o�V(�}��*��q{������*�I�+@'xIA�S]a�p�8�I�R_I��8�I����6~%!WK��[c���BW�J�VV32��gl�9�bG�Z�(��)�x1tP���E5�����.��h��R�.r�RF��k�P�b	)��,�&y%і��H@�޴K�"�.4���in/�n�O�`����\�!���ry�q�5�����ꎿ�A�*��Q��c�G.W㔰,S#����%Y�5Ӂ�c��'�ߎ������v�Q*@�H�=�^:ߝ���u�Q�\v�Kc�r��X��_��#��R@B[��$֜VQ)c���uJZz��7A;)LŎ)�N<�v����3�\�������P6�޶�"����F3����ԧ>`���5۱��>�"���N���Œ��/��<���\�I�6�������}�6�.������uvߧ��+nF��V���8���z����0`V��-��6�n5�i!����C/�0�ݤ�u2z
ͺ\���Ư���-��8�2bS�M"�|@B��qN��,�3"z%դU�����������mUy.)��uc���X��]������e�]� ����s���f̉��k���(6���-��ށ�yl�C��3�7>�e��!��8ZvF��R��n��oM� ���tk�1���ZO�L?���G:+6�o�l]o�I��ΪyЍ|!��R����·Z��H	U��^�mJ
���ZK|X>}2�(Zr'wA�*�[r��!�!�h�����v�20�>lX��!���! z���;�-��V����)zD�+�t�w�\��Jl��m㕌o�y/��`]#!4�D��_Ɯ~g��N{_�%�1h �z�V�U���m�9���+�!\V�J�{���������w�)�j�eD4@�A��Ͼ6��<��U'�ޟqE�3ː�fFW���Ԟ�IZ�xt��G`�V`��3�u��@Q��xsP�=A��>�#��'N��LX��5��{]>&B,�ܯ�|�ـ��0���NI�-�2�Q��q{ɞxlI:KUk^��`TϏ���-6Sve��o��ПTI�b�w:/�_��I����vH���QC�Ӝ��f���NU �q��g7��[�D��������Lj��/i"��U�Җ}aĎk�`I��ϛ�u�_NǺ��7��M7;�l� Q�{�t��oe�wz������������]�r��k���D��]6��A�f>~��9��1i�.sb��!�rXB7�Y|A����i�|��~���Ey̢,�Ԫp�gyo`G�8A���eVq!�w)��
��Q�.4���	y�M�D�x��#�(�z���
�3`S�c'<_VX�������� f�>$��J�wu"J�Q�VYG�T�TR�V<��HK�|m-�c3	�#ٕ���d!����H;�pNG�"�!�7��/P|v���u>�;]��A�f��co%�;#�-X30BR�@%Rʬ�>�1a���L�9L��y�	��s\����f��N�l¤�3�[:��K����s�y��m���q��餿 ��v�<6%��KE�N��!.��Z��X���d?��fLR9/H��hY2Q4Qm�tb0����y�9$�<��?�N�i�m�քgw`�FY-!���㽯�.�B�>l3c���X+l&]d*A!Sk��?�B9�F�0jm�Tp��u�ۡ-��#�C̒�g��!�ѩ`���������໲�*��ʧs��R���D��O1p�r��tLt���[��#����Zב.���z�z=4��
�����s
���/f�����y��Z;�Q��֞�lս�"�XǧɳW��o%),�}�h	�Mʗdy.���yi)qQR!��O��mZ��0?͹|{��Lu(=�S|�"w����"T�r����'�'���{!�1�}9�U¶���­~ӟ�Q*HB.MHɭbb=���Y��/
r	T�Q�u��:����q)6�lvY�e��!ο<���V�9hAd�L	]���Kk�����Ȇ���z��
���|C�)�Y��M͋L�/�����cS�`n�,6���O�Z/U��gn���h��n����/��J�w���Pa�V���Hu���*&,�w��B�J�
�)������W'��į�tϺ�|9�I�p���7RU���S/_#Œǿ^z�g�g]��Ž�R��kJ]��B��u���~r�hXŭ���-��c��e{C[�1���6l8qOf��"oF�E5d�2��m2 ��h�N�����
��v� ^�D��	r�;��hs"&;�U�8��_�U�t���S�zS�{p
����T���EV@%-���г>p���q.�qƧu�P��{,���+�)�S ﲳ��:lj�砗I|���f���|E�(�PO����:�Gg}A�O	�����'�FRM̌�w�B	-������x��r�T���%&ǧ<B*��ޖ��_�U�Ěy��蓁�ч��a�9����+���C��-J�x��p����g�,E������W5�j̣�q�o�f��NT�:,�$@��$w%���-fO2�����xR��vn��(hD������ߋ�Ѫ�4?�����-ɼzV׹�6^�Oɒ���Vii���{x���&�`4D�	�3�.�5䬪`���^F9�_���D�>V�j7̃/��8���}���g�>�Hl$���hC�؜��f�"s�a/Ӑ�2ry&/3q�`ގ+��/L.�7��CU&!^�Ks9��nT��I%��R>�q�I|��G����{8�����﵏IM������т��R�FΜI Ag��d#Q���:�����k<NA�K�%O�S�KL��) �Uo�G�V��v���,������{�7v�N�k�Fz���o��4�æc��Iv%�A��82q�7rW�y'�yn�2C��08v�>G���%]�Z��������M�������c@J�W�B��'���� 0�a�)4�*��p��?2v?�/�a�{�(�\�8�h�7�:c� a���*RAWM��X�K�!�����0���yټc�4mD�)~y�*8���=?m��n���(��˘��}�gk᜖��(v1!S�B�A�ܗe��T_#�Vg��%�\!�6'�B�`�Q�;�i?^"�ZP+9r�ܛd	����K�s/�Is�u	k��C�n� ��@f�A��A��������),��@ځyS7ӓ.e��'=�1p��W]����H ���F��~!.4�=��!d��+ H�UK�S^��I���N3���.��,�>�֯���A�zY�q����>d>K1g?��)S�U��1�z�<E��{-���J�Pu�AT{�`���£ؿD}�$ո��D��/F6].\��wO���Lq��Op�F����)��9�t��w��H�Y��e;�7m�����p:t7��FbL*hW�=�$�\��U�DBH
,:nh�5�ǽ�P�*�s:{�GQμ4��k;�Nnwr����n��;�ï8K�駡�"sJO��'����U��K\U�Y?i.����"��!;����2s��0x�����=1{F�(=����9�"�=$�0��H�ڏ��#ˠ΃����x���<��4�3�9,Lco�5��c���퀳��Y�I�T��՗�S�"�}`��! U�k��~�̼#�)A��Zv�Ce�����@����)A�4܋{%}�zU��s�bD�M�0؅�h($����`'83=��F����i7 x�^�;'�/x��`^؝H�9��z�����=t&����[��
N��n�K�*`$a�f���ҍ�HÚ8���)�����*�~]�S&��t.������������"ƈ�'�Χ[[j�I��s���	��J�R���X��"��K<���:��F���ߊ���;��B1&�"�-	��$/�+�l�KRuMV,~P�a�oH!?�s�U�V�-^7L����l�����l����H��l�j��	�1fj��c�υ�g9�t�Ӯ�s�~����ƕ�-��<�������T��l
������A�Z�d%4�A�C������5.U��	�ّ����� C���C��VF��h�l�궦�а3?�ݷMݞ�Ѫ�S�@� ����@�2[�b�\6������j�ؖ�M"�q*��G�i	�<�[��!�^�*6��!�m~z$&�Fq�	-� ���	J�m��DG�眩	å�5�	�JC�&���)r�i�K�=�kdO�$+�}M���=��N��`�
t��P�iǜ3���k�/~JCÛ���/��<^k�g�V�: �X9��I��s���1�I��=|qj�~hb߀�z�G� ���42ؾ~���R���;��/�-l�"�)!����廇�~�6�̲b|G87E��o��D��0�kI����ҁ��;�m��A����`w?�/A,Q?H�#yx��p��������t����7�0�[��:n�������.���S��Q���^f�0��q�j␵��?�0���q<���[�
������vS9 SO�wH�bK�ǴiC�o�:]*G!�v.������o˻ov	�M�H<J�=5����xߪ��@'u��E�
f)V���i���� u����вSR9��U�y����&#����nER<�	��ru�x7>l�S4�7��ی(��S��؏�3�I��ԗrW佺{����\gzFr�0b�Y�8s�$����Uu����og��.b����b������,t��m�K��Q����{��sϿ�`������p�t=�s�{is�"X��n'�p-�9,�,;�䜭L�T�a{���	W��I�����«t3�f������UY��x��$"��s1�Y�J����j3����2's���oo�,��WÅJ�J���m�4cM�}Hg����'�Dw�C�t9�@K��#�� !��P��������g���ܷ�`� mW�)Gzp(]����xq�)Ht�KY������W���:;{h���+9�k�+l����&����ZW*ȭl��^��ɯ�>(�b\������﨣�����!��z�f��7B�3��YaALK��Tq��|�qq�B�|���`z��"U���t�ɜ���GX�44NHIV%:r��H�Uk5^�Gy����*����(�����2۳��*����x�DM��"�?�9�0�)� `��9����\Ӟ��ms�_¼�(�jZqک<}vc�
���=�7.�YH��3���"�I��D�	���<$� ���RbS
C�_��!�|I���雄�@6l��5�JzuGu�q����L#�G�����j8�y�t�"�g����V<�8�\�Ӈs<��#�˖,+�q�0��G����jk�0�7Z$����&�.F��s?Ы����D��'=����MZuT�7�h��V>��3��@�Pr}���*�n�[�̯}���okϊ�ިʝ%7��r�V"��x	=6��Z��7�L��Tԇ ?�O�Ϯ��s�
j_ob+��T�qGsˆ:�x�e~��I�K'�Yx���7�����ܛ�nݽ4F�|����#��t.��A�㚏FD5X�~�O��*�^m�u��On,���O�+�ύ����s�-~��}�nO��j	u�,����v�Q�7;�= v��� ~�f��-HbH⪠�2Пl�c~M��rVЦ\���6?�_{T���?L�g14���)�����v�K1<9�0O
���ݿ��Ɵ�@X��@oV0UHh�m�D����=�%@������i���>��E ~��KEO����Bx��$������}&.���q��å�u�z�HQ�_%�	2f�,[w*#Wq���������mӲ@�%P����|r·N���h�y��f�(y�����:�N��U�.5��l����yUb�"�؛�ݍ�	YmJ"usf�W���o��_)�,؏{j�%��:u�󱗅g`�0+�]�k���w:�Q���l� m��Y�%�R�Sϊ��m�����R}����8P��zC�(��(;��.bͪePw�%"P�劲���-հ	�u����}e��=#a�����8�7�@�納�8�9w/�Mi��H[ ��a���`��N���C��iUY�C9z�C�i�$4�}˛BÁ����\`���ۨ� I��$[�@��c�9�������r�Jj��^�Gd�0���0�ߝ;�;����Y��R���m��3��9)��g��\h�%=�h�F��G�
R�WK�JER�JJ�K�zoޯ��/2���J�H�58<p��^T=���?�q��E��R}#�Roҷ�2O�r���d����)8	{&�^t�F�B?6*��I�5d�5n���r�[y+�I&e��� ���V"�mFv�ɲb�ԁ�����W�3�1R�Q�M���g$zЦ�9�7?v�6Ԛ��k������x�2ag.�hA׆��{2_��U� ���b��~m�3��S�p�*`�o�q�[	6n�`�v��x�l&��Z*}�������䃸����S��"	��W���;�	Z�QF#���]�Z2(�M!��/�p�~5�G[ؘ��� U,2l���m	�K��Y^�r�$���np Jg��%G�u�6��>�� aڍ��G�=��V�&�\�6�1Oz�TI�KnK�ѯo;W��R���$P��K�/��զ�P'E��k�|a呻���-B����ӽ?ղ����O��'h6xh
F輬cCvP�ush��#t#�e�g�WKA���rci�wE,|�6�3�v�4�פg!-��K��%&nI��J�XӦO���ߑ��������}ҍ������2�1�O�e������ ߒS+�m�t��̩��,���P���C/B��9�$:{��d��^�������]�Z�,Y�+��9Ql�9H�T���	���<s��'�8뺨Q~Ӱ����^��7�i	X��	7�D�jj0�6�rK�?�c�ꧻ��|����W�n ¥�b��S��%��?粲�(x�7<�fpu#8Z{�c��ρ��vV�^j�I���+.&'�X�PJ�0�l����O��b��"ߍ�u���z�ti��/B�~T�~}�	�.ks���◌ia�I{e��*��Q�^�� V��:r0��z�r�:M�=	(I�d����@�� k�9`������O���.ݕv��B��� �VXd� 9��8(�5�+1j|V�"���c�x1���8`�+�M��!���h�>U+� %�N�3�9��G�$�Z�v���_��L�6�s�Xi�D�Z���8�`��6cZN���=[��Vo��JJ�OP�f��՝��a\��.�2r�S\��A��J��\�s�r�0�j��P�oQ��ٔ�5��l]��Ʌ,掋�/�����������Q�N�9T�h�W�iupP_��]�ZV��S�Y�@�U�<E\������k�Ŗ'���(�X��f��c�1�+�X]���C[>��;���G�jV��� ���j[�`C���șKU�w=?�&�~��J^Ei����L*����Br����"�-��mll韟�F�(��ZŖXs����᥵����e)�j��@ZU��>rI���nP�s[�h�k�4���%���f��
��kr�c��+9��ⶍ�z���Jj�%�?	6�9�H�q���@II�^�f([t�p�q�s��҈��$��L�@ʞ�yZ�k�'\�)Z6�j	��NYS�۴�� tS�D�ԇ��W���M�y^�o�T��O'�ˡ�ʦ|v4�yo`�RR�`+f�ճ|&�苣[t֌�e�S���UPK��=�!�G�����[�f|M �i�6*}�p-�����{��9�W��Ǐŧ�b���� ଩����l�������Ƴ�c:K1˜k	იC?��OK��m���e���V��Po� X��DzŕBs(�>M�@>�&<�����$�J@��'������^H �M����z��2�#�Z;��o�Gku��D�8����l���.����6�7&�
s�"W>7�c����Wps�r`my��fo����D�f��-M����ʜG��6b>��Q8�OK�:ە����]Z��󒶠�K��T�ffT5�L��֯�l�"��f�[2txi����)ԁW�f�����!��p��eH	��\�����q�X�!h�Єe�����8�~'f^W?n���w��<&����I��*���w�����큤{�H�("��$�2<��W�@\�讅��_QS���� y:���Wd��iw8�G+KV��2�K!��y���L���6/rƈS�v�W�����-j���B�O5��l��:pbj�)�8�>q#���-�����0���쌻D!d��V��0��>	��Ry�<���+�W�1a)��93���]Y��,��f�:�	5SAa�-7a.�N��$�]9G���K�2xDB>q���Ж���zL�������=���<>:��(����s�mRviZ#s�a�9wяĉ'2u�;]̄ۓjF��v�$|޼�o
sM����I�v�0�1)�o :�t�]�7L.f�2�3�B�O��Ku̞)
h��n�N2�,x��&��Ԅ�@z�~7�9΀,��AZ�_��M��*�P~� ނRk�z5^�%�X�T��MM~�Er���9֭E�s�K_���C�i�|�+t���@	��6�_��]�b�K!��&[�N�)���~�o@(o6�过1z�r���.�Ns�w'>K��&H�ĭ_h�z�l8�@PI���}�)bv�N|�{�Z��L@M���e���?,h���{�e3�\P�p�Nr='�C�B�����m���;�rpz��{QeSB���*/�~��T���QA|�����Mrx�RT�B4�GC���]?ҍ�0����f����!|�9�,�'	�Ӊ�H'�������	_N�op�����g�����7�9*:��E�=fu1,���aN�#�Z��@ᮈ�)�Cd�.요b���~�u�sɓ\SH)Hb8���%2طY_���F%��=��FpG��u5!�+�3�큧����̓�'�����L�ђaC�u���#�BE���g��C�j�z>�l��&�p�㠺զ�,e_���CY�*p���[
F�vߊigYrџ����>��n����渣o���~�U򪉯��I��j�ݧf�y�]0���q�پ��O�{TL�	r���M뚱�lԧ�E��)lܥ�T�{����5����fp��U�g�C�a�ӂ'D ��0�����&��d_�O�ļ��n��������h�$:����/�0�Cq�4md�]`M+w����D��N��eO|����+�1{�g�����	��Nʰ�����e�C?������X>:3�������f6/v�k)���{�|�E�42~hqz��F�M��-5�\Q��x8�7n�}�����\�rwY&_#|n�(���K8�{��;�Ʌ�?���p�_��֒;�AK�ϴ�Qۥ
�߼��0��'��v���<9�?1$�1��<��F;S�u킯�O@�P�@��Ce[*"+���p�7�X��%F�4o1@X&�k�9���Ǻ��ulS'�q��Yo	��i��Nob���M�k)5j{��	��BK�@�,]N'��$�6�!����5zȬ� G1
��ˮ[�I�fKK�98���F4i7peE)4UZ����j1�I���G^���ȶ�y���*&yz�;,� ���<���w�.Z�{~#�i�~ݰɢ�5h^��(��>ЋS4c3w�"*��8;��+�M����],�G0Q*w���\˗=A<	�(bd�I9g4�R��+�h���µ'�H��������F�|v�x(s0�`���8�!���L�h���ٲ�(�E(.�i~�b^#Y��T`�����$���[��5����C�u|Բ˲F���d���U.r�C1���]����?W
)��c�
w\�\t`�T�ODQ*�,U|MF����jU�%NÑ�������OE�{:�� �.�]�9����ʱ?�@�xS����˻�����rB�pˆ(Ia>s�]>���^X� !���Y��8H��}�=2m�s���W4�m�O�_�8Ea:�މ =�[Ӵ��?	�H�x2���&{k�O� ���x�t'L���V�ؑ�Y��#MD��ob�"��*lQ?J����/�?�[L�MO�C[��)�� ��� ����Ͷ���t��v���P�Z��>��Ok~�{�� ��^s��d9SYl���̊ĻKhD(kl���F���^�=���O�����V9,;���~6�
-K�Z�>�Ł��)�Z\��e�b D��xw���הE�S��ʁ�V�	9�1���9 �(-��������������W1�)
o�����U(�[-���� �7�k0C+߈�"����s���?�g�������� )�>Rb��F<��m��^M��'6*�C>$�G����K���ub�Ux
� �*g���Cl�mEm5�X����{_�{z�ɨ=�މl�J�����ex�s���ԡ�~���H�T�e�C��*v�mD��RU�,E�-{�T�*
A��/�AA�t������A<ge�'�֎t&�0���8t��pqP��;1,�z�G&L״w��}g���B1)�5 r��4��ː��OߓXv�pA9P�vV���$9�����)��S�O"*=��}�B�m�k�E<�q1cJx��Y�H�>��U�_4�9Bj	��r��:4�Pw+0��m�(�b+�wq���%.o>��z��5�@<)��"���[-PNc\���w�<��O�_��$�3��J<�;๴($�8���z�� zG�D�F��;$�W:��̲|g������D
g�}W�)�5�Jk]q'��������t��^�'1\��i�f����x��p���]nn¹��#�ǁS
8����S?�ZTS��!�}���^��?��N��Q��5iOL��'mEB��"K@�v5�>4�D����$OHgl  E
θ>��; h'�*֗7ަ��BO	�@���'�,����F�)NI;!���K��\�t[�Cg<��sF-C�-n���Ȉcp���(�wW�����Z��I(�@�)?|a���ӄ�n���)ya$%��6-������\�<vzm��v/��W"l�t����q7�[����LN���*����08N�G������ �V�g�q\}up����߻|��GE�	6�T���=�"�.�b�~�Ǫ�E_��ջLf�@�fY�A
>��K��:|C�>_���S�@eE��54�CcpYq����]*`~��'��Q��f�B�������@,}�?T�H��)�_1JN�����|�����]Y]f�㲋���
�>��`_'��b��2HV3�
���obx)>�˹��EϬ���� ��
N��K59��o���a#����8x�~�P��R�`���2��ڥ�k���D�����G��d'j�ϛ�d�ƧO��� �ap8������@gR������e�S�M����g4ĵޝ9fno\�nR��8�_;:�����)���,>nju��0���1�v�[�Ы�#�EaO��W*�Rc�~��dd��Ӷ�Mt.����\�^�n^&/��S��}��[b�)�;�Ik>�$���ܝy�����wV��#�N=�e�y$Ӣ�
:����EN���T�%k�+��T�Qsl�b��	�B�|�83�шJ�7?���-/=�T1�5[M`~�����e��[�F=l?1��mq����̽�Qd?t���3���``w*)Zl�|�I[�1z[��wGh/��6W�g�\i�9!C&"�A��_�}#��������ɺ�mB�P��I��-�v���?,X�o��>��Rz=	<�3���b����"iLUL�����VX�K��Q��/���Y��f��˖) ���]��"<K��~'��2�\sddH7\V�"�fM #��'�vx^I*��ѻ(45?
�ߗU��v�@�����h�+$�+��XUH�o���A�R�gÍ�K؎^�F����!�ȕge���hp��v��Fs1��`�.2*
v���u������N���g�s�!q`�.�;:�e���4c��v��uR�uL�DJ*�|+�����m�߰�jҋy�%���T��~��}��E)ȝ�i��|�Bt�F"_��BlJWU4f�6��w��{KM�"X��������Z�=�����|�7<�g��>j4��}���Ov�C�~3�-��������Nx��.F���%Z���z滻j1�ު�ፏ
0�����m�h�A���?C$ψ��R/@z�����A�^��V����j�&0�����ˆ���gj�8���ڷ�ݧ�pȏ��8�"����Z�Wǐ��>�]Y	�|}N�{��*����[j���!�����y�g^�x@݃24.�b�0pTqDN���Un�<����mZ�-;�h;{��S`��K��-8/�Q����m�-�9$SqH>�CB���A�6?�:�$���WSX�	�90� ����ٖ�X�߾y ���3����g�eП�%�ߜ��`�¢�gtZ�>s��.\� X_rօ����c&���t%���6z�@�.A�Q�ң�*l�U65b����
?���ѩ�c��z~]L�j:ͬV�u�VT�fc�O%�( &z!]?x���m5Q)0//ԡ����զ�W���$7�P�_�[x��_��~��S�sġ<������>�̈́