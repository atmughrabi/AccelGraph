// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DaG0Wda4hE6Hb4gyvpYHVHI3xLPl6FGtTEZ87MzZc7ScLMfFuBo0TaxtvhvtaNxh
N58GA8oS5Famfx63ylDGIf23EltYbBYKidJFtkXoXTWWyybSoLVKlyEHuni5ckmq
zbodecUp+ILVsdf07xZN0xZIG6n8BnhE6jaa4kzZVnY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25440)
s2FO7PQ/5w3y8p0R6eYHaF0MAJ/hLTHbup/vHWOctGiObnjMUwi+dWulXGPsLMPy
HO69yOyx/Ln+wwDKRygsXzwTCuHeS3J79QEYVp7/ihvKJUbW2YWJgySDVXFcEFHQ
ksuptlGN4aoF/4om+tFEKkYdy3+rw0q7xK0sbF5XHFhNVEKZAVEEd3+8mzfklPaE
fSm/+MHDlvz7kjabypII6aWPUHNSIHdp2jBALKKEzlP/XoyRzbGvEP6fmUe+ss1u
dmisUVlahVk/AY/LWdNtG78Bdudy+eDWLFO1TjoaHP1ZE8xtMBRLtwVEIQsrm/Wy
e1jUyjkehoIVzMDIebaZ475qp4yYAFknKNtJkQH5jaTspBrL+yX2+TU1c8l9q5yr
xpaLY/OKbIlWAKD1dCrgOiOXPzgbTbT7XWkNidtvWk6oV8nxU/0qHKzihpPP46XI
UzQci9udy87wOCg1soyJ9LPbYQBkseyadCo/wKGRA/2EShOTlAQXJoEu5yULDCO4
wN7+DZQK9+9cIQd4m4keW2Q2iX7R06niX+1K2avhiCSZeE9I357isRRn2dWhqHYp
I5g389BqGHP1Jq2zbFH/xhDAUxfLS+YaNCLJjLfdyE6yDhk3CXrSjh67DyQGA07x
yGl7uDIfQEWPV/Mp4+4ok31CxkuYZx/Tes6IYaqjlNQYsgM1asIYRx3HM2iQZ1fw
hBVE8gDAy7iQDYZI6PRCrklWj9oJj51POdwy5ZO/EKqNSGxjZoUv7dyIc9cj9BDE
/eG/ytp0PZWuwCEWxoYn5eSM1qEwLsYo/PUCOiMP3CBVTRmTyl9VK2dQML+67a34
UMizxq/mXKqBGN9/xgdLJwgcJOfmwEw5UJJXCTulNu86ogrklJW2H00yfaifujXf
5d9GlD0xmUOR/edAqofo29xqPCUc+9Ea/A9XwAYevZA9xPHsttdXmp5BQTrrIONI
u1ML0Yd1xgf0XWqnOjgN5GHGDgkIvXDeN9HEK5qjeSTVrEkz1na8fL/L64Q3uzo5
Dp6TnNvdz2UFeFozv5Rfucl1plse6fON8I/gf7wJU73plHSNBssD0maWyuQ31MGQ
yOAC3tNOBQhiFgNz8Yu3vT47gxROecB4plLn8LIv7wG2ZbssvvBeSC9zvvmJ1fcw
j+uCZgc/Xhknz9Fbl88m3cOOB9EFGKEqQQ6rBiYiIHYB/TVYTT0S99DTtJYR3RGA
T5e4+Ap0lsLHW7nIZBfIFsFhNQr3HHsGzza3WUcAH3iAqoVx/IzbJUUk8V5bgfB/
VpX4jLZY77FLpLwz9h5YIfLiAjjydmo4QladrhhBYIpWC5qg/jiwH1UmoN8liuuH
8swNYWuy3+o1P7sO9IyyULqBv04+cDWa5W1tkXy1zO0IhARZ7O/poFnAA2a71AFs
4fehS9oFmY3AOfxVHVs7LqlJdUV96NS6TKKrwyJDhFpRsMd3f5k30TaJa9NeIhX1
U5yKysYHGuYs4IfrETsys1YdbDEbFtPfm3SzB/0l5X24jEIxUT3AaeciAygyCB74
9p+6bRBevyW201lFH70sFcle34xzqn4uelc4G4v6Dfh5hzLRNkdqG7t5/0eQlej+
QQX/W1tUH+MBAqkxhS6BnZV0mhICaodbrnbPR//iMSFbA+T3BhJ5p/Nedw+UMpll
bctMMqcrrWa3JU47oPk+PI+2RJx29YilTA/wuqkbTm4GkBAB9YeOEd0csMmM5u1C
aLa8wxbQgkJt/YQK0YJPvianS8qo1RyqfytiTHYs9Iq5rDOE7RH7ZTD+1l0iQPnC
Si8ssB0cuO//Y40VHczrd908QrRoNY5DRrbpm0ETjLnF0bNAOCp3xwFt8KVJ1lGs
OBX+UE5h/4bUCvZScrR9eIm8ARgAWHWsgthcnwtdcJAm3O+l5J/Q1p1GPnYy5iZb
mhLEpbGu5oLc/2NzhCmYoKcenTkpVig9xltyQOo9BssOvxBzKf5lrPB5w7oMnsVQ
TrtHQHUd8bk54iwt+lLiGvGmPh+bsDYGPYWd01TDpm9oEWIy6kuxEr5sRwmQkkCj
EBJ+qOlzO6FoQHsMskVODO06maWq88cXPTf4LBaIaxr8Z4CqGkGAbgxrQfCEPPXx
DAirPiEMxJX1VggrvoFdRUnbkKhqZXzYmpf/L1XSkuGNqi+l0XQRs5e+GEcBU/Yb
HyrYGMz0hwrjYIs/zKO/BmZnSnHr9yHspPOHRQE2mmxbCK3Do829OeXU453AEJ6p
pgzgLu0l63uc2QaecRszUIAA9Fo/u3GaS6kWQsV5PXtfxi3tixAO4TxcoeS4ob0+
s/2yuKzE37HGjLDGH8+gZPexZoHvS/72oUH/S4raCbQmUYHQDbAzjVBHaxtotsNa
g5EiG9ZWsanenmvyB1Ht7B2QEIau1/CZDJH8mI0sfNzqWishucpZtUogH3YJ2GTY
hotODE4p8B2fnEcXuVQGFS3ob4fJ2earwyJ8Y9pOEoHqi+mAzQuSOnSv14SdL0VH
EPKNP1jHOVI/ee6muDcr4wNeolgsd5+LuY3QsVWowh9GdC+WsJIPEtPkd0D0tS6l
Qx/WKCbDfUpC5AGhYtoyB0JhJ0TZoZ4NZbpd6LILyOdP0cyMc7ecRBqVYCSt2mOD
/mCQk1OxEua29aGzVKZeCX3jWJ8GVQm8vRzpKLYQRZKoNDffl8z5tSWjASQtJZx9
UIfw9wtaotkiqV59cLSTK/HZt3C8FMRVOegT4vaw6/ot2Db+ji4n22+wm+8zfxQW
fADYkVcxjcDfdlQJCMwaMWc0pQQaMpRk6go9ijc0ZT060eBtDNyJgx2pY0ef4/Yq
x8062Dl/AW7CauuAxJwFkTGYyn2XxyNkFo7Ln0v/js/1Lj2l5nuQ7QA+bkHAlLu+
sE35k0Jb40RV6quA/ATrjbGsugJvSzDUsqPOyNl+kxGGs0PLnz3nMriPkyo5go0g
qpdD9yb4al/uVW9Gxa3bUNwoLfJpXxSha0vi8dkBh3i3A6izetNtuDKvvKueXPm7
WqDU4HPvudHNU29BVsrXd91qGuVS0QxNCSYkSqFi7Tvo4SBJc6cGjDdHGR9uiKSJ
gwE1klqxZeuf1yKeclIct1j3YQBkIQcPY/2xy4rhFX3HYgtU00q36IeZOtuw672W
6Vi8Vspzjnz6akozHr60zVbHXRcI2Une7pSQww08XwrIzHeIin3/VdgRiMZAzjtn
iKre7FzPTdrTtmD/Too2ObfUe4kaZ0Huo5wplq94EKXWF5VfbaoLOrLoSrFRUvjZ
bkd9OaJyQu1AHH7ezvJ3K7OXNS3z8htN1YDQ/hfbRAdhq+aBLsK32FPoxtlyPMTi
nKAG4uq8M2EpEBLioRBIl/RfAF1c+yk5csWerBd0jB+LbK1owsImU/O0wL2wGhdy
GkuQ0hUBKKb3UDuM8ORgyRJ6i3ATdE4A3r9fdCYo9ZQ0enRbHCOJdjpFkOFH8PCo
/UIjLWXZwjbhj581FeGWM7a/4vLw0sIPkOnY3EfPSiu96ZFWGvJXamshsq+uUH/l
f/NCtO+L8WpWYcxc1DIaKxmpXJAmBzh25nkAMD0PtjhKjKc4ebEehzQ4/BfbH+Mn
CBTYziTntiVaXfewtlituF6CzTFg2YHD5mYcrY4heGYe3zkl9gmxcBITg5qfUx0O
vjkiAQM4R3WC2ya12qZOBQvGiFdlxnPB/jJnwSyMdGkjB4zJB/YHuA6v5J8Wu6y2
JDMY8Uu6VQHMi99RZdT9eUXDMvghEbMWqczgWXtzrk9gxFqOiexLSWJyfSUHNcgd
M1burZX24K1wmXcJ8ZQuKfI5Flh9LBaH2RiFXXcxo/nW4IPOFUmanZeDVSnP/9+U
8Ty644p1AjcG2EaLKjcm78FOID/7JcE4yRiKxD4KsBeTjF9F9BxxaTrvhLdu5Ikb
yba5hB1igpKmp9Brh6vY1jG1AyeCcBWEwCDB2i6aXduCXz/txq7ERQdMNNgICB9x
nIUF+LhL0Yc18O4Kz7sPB/3LbEM1rzUAOIjayIaOuGOeZvQAdc6rIe4Ve/hoNPRz
y1frUGXUZMJNfgpcR8H/CYg85wtp21UCqpigVWzIV0yGOi7Qx3lvmku61GjEEPPU
63L//f+oqNQ8gkSKrzR7ySp8HeFkeV1SKVrgQt/Y9Y+4lbrYreimwTNbdZQLu5df
z+QSwASC7PlA9J704DnAsbnorT4bWzPbHhmPuHfFTxUelyEwdw1hVNAqJ9Qp/m1d
tO8snPhBvZPZ6Qe5/7KSAUjmH0on0Nrgn95IhWXMUu851moLq0DoC9ne5w5Gdbrp
mm4SbTeWzGWKVbfHsrLk2l4O9iLOO7iQzINa8BVPRhUlD3w5UhoorZy33fGWoYW4
VqaoLVYCByheHoaL20d8U4fvusFHeTdtOBbfzbcOPk0oS9vVuY7vnpQfOm0HvD9r
q6lbmkmQn36VdPbNOdw+tosb5fBzCLNOC3EGarI6j4bX++3pYeh44/WheMzgQ9bh
o5EnbKcjKfbynpQdG3k7cI1zVg1SBCMyAOzzNESGOxKkjK8Ao0fQDlHck1JvVY9M
znsxz2YQpdaj5yVxX8hTe0kTaPzQWDLuJOObGl3u+OSJqe7MeiJjpWSACzmd2zEd
9eh5B53rd4RxgBx6uwdhXFx+xlebPZu5qPLKtRAj/k60wqk+J0SZvXpvc65S3Lqf
uqrcvi8/6Ovd7n+Fq1BUe+WH28IS3FF4hWxwlRTpDJvEcGGdGgftfGtO4NaPefbP
6Uf1lVz25QX8WbQ5vrqriFJpkT3c1dviRrOk7OYfTolmzJLM6PmvSqiLQe5ayRWz
cUH8+HtcH0ZYCfnK8aH0yc/VUoqH6AMRuDe/Q0AlfMc2gAtBFZzURmo+MgUQ9mfe
MizL5evi1Lntg0REhnbmUO57Itqtt6iggUMa+02ewtu8Jx8zfLZau1lxApWcc5mL
AfedsidKjdsk57ULt7eMed83EKf8av1bZwrMm41JBB8xo/vUImeLBVAN4SasHCnw
lt51rsAlL/di6O5btIhtdn9hw+gYCW8ObTm/Yi/24JQVnrrnDDWjTwAVJEpTcIgx
W72pM7a2XU1myMWplUr9AqrwRhNMx81/DHRg+BzUM+PWsW7C2yqEDPLGlUXHvzDG
9f0R/1siFlM25p+Tci+AMDgVUXUytkfxxeEa6CEEhw0VkKvXCI6WgZVRA5kYFK2y
qrGFPupCdQ1kOCOc8KlluH1xUVE1oKNFwD7qeknqbDspoCFRRVOkKHbobbZKL9d/
9cyVASqAQWEuHu3eorddcb0TlEot8jk57eCWwOTosDx3JGUBkNToZEU0pH5yzVdP
biKQw/pZMY5bM2Nnw+npS78EM62KrODDMDNmbzGtPosV9AAzq7srlXnqdwQyQ0iO
EC3kY0NDOWL29lsUj3GLq1eZGNaAMeTtRmyShB3RkzE9Z7LsS6o+aG97QDSoUMcS
9KMJe7+RGTpzsT9S7yo5adRxU7Wa+cEM8mVPuc8o0QHK0oSWLcqLnZ4+jsaFpIGy
lPUmnU/Q1RDXaAurgMHS2Dj20LOr2z/pq0kxQR1DRzHw1CU1DrHVGbpN3Q/h4Hix
boyzgDgTUuO7rDakdL/SH82GITQCW3Jy9rqAIjP9Or2JrrDE4bdjiuMTysvID8OY
zJheYO6AYvZ9YQdKMzKKqqWBDdb6RZFz/dMXDarC591XYeXmodOf/afDY1GL96Ke
OpxjCewAqBdt+S0sjRscHzHW2kNQb99tCeUzHQ7PNXGSBeasrdlXyq2NANzauAYa
kzT5yUQoH7IwWKNgPe+RbV1wPH/QvgrGV9Q1uxCz/z6kvw2rCWvnewjadqdn8RIV
3JsH4AmFdm9zZAvL/mZQyJxLSurrP/J9RM8aDN0S9NQCLMhJYLmLXwYM3RiVdQ88
8ksyk3ne+WP1B19vLysgIk5s9uYkYmCiNlluszU1Pq1x5lgO0HVNkR4ySnEP0wE6
pA+WQxpV6oSRBHDBJ7QVlU5xcCZ8sQQCflILAtUCi/DkbmccCODXngb6Ic3VF4IT
w35zavilqCm1cmrKuBYTjKMUpiCTY6F7ybD4+14uOokt9FUC+eYMIONzguCXSYQE
jiIb9826uu4C1FyrCTIxhOJjhEmMvjX6M/Geru2k9g7IOtIDk/BOvJfkcsJ7pWPR
nmVwTFzQuLhXYTPcgI1HTIfgrDDadTfpZEaMlblvn8A0ta+SIpVYKMv28YDLQd6d
X7Z6rQEOCHOSu3Ockn3Um0/GvDLv4xwYca9Y69bBbfqSpJrb9N6EG7rNlD2MrB8r
GYPja8cW/1l8g3sepR3usFRwLr5+Sex6LveeHoLYQTGPZdn8CVc+sv72/iFE1DcY
lcf6fADAB3owANi/U/r8fw6hmxg1uxKxfL9muJonU5vHs0Uaf47tLEZ4mLZ1xlMw
WA/hDjB9CjVE/H+OYzVj8a2n4SvlsMqrB+5LRl4k4tSLDxRIYLFoyl2YFPTCv4sH
mWejVIVfkUff4Y7xX1eoJ3H7BsTcH4Sn0SrwU1kMxq25pMCKifWR8Ai+xunvMlgt
mbiSRqchyjRLCl1wdfCF8BQzEulqyCzAn1CmNB0TbtnjFzoesI1uyTiMdSwjCfoC
sAD816vb6Lh/YE9Ujk+uj+gNUZ9k7T3RH9/bU3HMYQM3nDEfj0ws7C5v3fpffIeU
IaD/fFt22fR9C7O6Xs7eZgjN0Uw1RiFKR/RTbB2sllYShA56em2xZrT2hrrOsd7d
OcHoqtZSf2SQBXXaryuBGzbFYoxi99d57Cu2YK6Q7xJTYm7mhaEDaSYvf+LgxNPI
Tu5VPrs2iwPK8NBpgq5EOrtjlOU/wZyTxbro3iPGrE0yAhk0aLfmrcG/hClRqoeA
jjuk/IMB2il/nyzXvvQNBmI2Jjzl5zf7scN4Q9ETlyTaF4ARJ4BDikl3KGRBNGZS
BOozKv/UClacRZfUd87/Z0s1mhSXuCvo1L2E7XQPAwOsGgGwTP7JgupBC1p0flxE
6Ba+/t+a9ol0yD0tJMluSryVHCBqHzrwFBxkSnZy/rKKq3vyClbtHkUeZOPmJ9AP
t+qTxhFzcC3mMWmQH1DQpfBOc57cfXsjhTTdMCEnQychmyJJc7+JUYgqOmTq4BS2
so/9WlI4GkkxeHhVPKCaNWXkUftoClP2LIuojoKIWymhyFKiwPTwvmNyd2cOulDR
qrqKzRifq0QLdDMF1dNAHW1VzKlE3HZiz1MwQltIIRigiJRqK27dk1lqvG38aH8Y
e/6AGM5H35CWYZjFxO3o2+enqGePcDzntku6S4fERhJ3KU1Pn7XOEwwC/dX6jT7e
5IRoJoQnnVPz5dj9Qs7EtgPIjCPpOONN6mSfLFf4gQZlxITwr/s2Y0+qnNfHNLaw
8908jaCqnMseVyxTgwTHRGfpGuGbOyuj5HGuiK7MRkhcDvEp/pLS4N6DiOLl75Op
vIK/yAsmGv/SzcuBxAlqrdKwBBfkOTpGwhaa4lwtEwxXVrjlkc2WDpD+PNMRZDXJ
oSHnU36rckL8vI5rfYiMWh1zmRHXO7q7YmZuSufmLmAMK8elmoj8IuzNKk0es7OQ
ymqCCIQ0eTT+7JomyFgrBqi7jzNQ0HMnZLlTPqqNaRaKaJQjPbKjYHHFX07oYPAX
YgYcK6SndT7HyGb5pCzHwN2FtNgN7Of3OLMLW7fUCUWU4FY/IrRd6N7DLsMii6LA
AzyAlAHQzsh6+eMe3JZ4nJwtX/CoRgCQ494gxowXCb0tWGxSAswj7wd/6ybRvgRs
Y6t8DJvl5kD9QoSx6ye3jl8Zy+GEXOORes2G8eWn0mwaoHpu8ybOspDxlCr6o9h8
i23RvR+3/9h+Ks1o1VreUKvMqdQDBgnhy8MenCRY77ozUKAfMt5JoxSCC3OrMc8v
Lh5fU8jzLY1/MBoCVOn9oYfYbKrFnEtcadsZX2lKR0aU2JrnmbWu04WnY/8D1WIE
ofgH90Hyyoukp6TorPfuWx4lnU5WwUVQYXSS79TDEfMQO0DqpZ4zeb7LU1AQD4ep
NcLLkRHJKwkkw8OYIETpwfrX42tc22BdrdDG1tmpblmK096WdLNoACBFG0QMxTmH
oVczXOB6dgMNekgiOFvhuGEwOsDckBjxCVxhZITl6CgZPrYzHO6S+Vd/vZ35fB5I
ahh+N/7Oqbi8BviQ8NDx+VbY52fp3UMNTFQHZnqFVBWF+tBrq2rpsqjoIC7GS/YX
NlQpYAaYEHJg49n58idZhb2ZNyH5ygGnRbMOPHm3pQrb0foKKS1sBLnri11E8Bip
hGx6NKy3nzCo9a8Hhu7nuRwNaIdHVqckuABRY7v5L7sLjimy7Qv8H7GguGb5zl+O
GbPAVsZVXDZiDcr23Bc8N9IL48H3LEU7qjVEAZPQzqOk8+F3R5UwlAW7naYu8SvC
1SQFyrrzcp91lNYjjrStCHNFUtujpTPcGomnlJDB4VtZE1E7epbr/ajGFDG+SXf5
srOM653dtYvaAmIrjeYWfvtglYSBI4SW2knHqFhMpp34w2+nL0exeR4x4U+CRNzf
BFLrEFjooeUYtAIg08Rpv45Scp+cRrs/b7oKUUUzEjvdD8uoLqGOI9Rt4Sd+8qyH
Qqo6z+2BBMYdWeHFdgq7R21BOlMNgYWx2c3ziPnnhG2Ab1aoS+8MgOXHNN/2LBfw
N0qW/cqc0I7YZIAM9rJ5omj8Lm2qEaq/9OHeeJNIaRpHYYIqfx2v/G+DX/lEwvBp
oqksvLbY91kKQRde16XrOt1Py6UQ4hAfIm9Dm/1p4Yl4K6rA/MwXVF9wxS6sEiNH
bv6vBcMjY9+OMS4ki3FDOLMKopl3XGDih7XyQYMXXFKLofUXD5G63L9aNlDHJ6be
TxIHlWwnm5EIqschaap0ifPLw4vqa4lqlJfKfPEUMnWiSI2UFzICwDds4qw5oy+R
lQeGxLSL7RavO9eKAVIGdlMvY9Xan0RE6JFa2KLuV63/ZCWGyhMG74XGRTk/IhCA
YBggN8zk+v7SmiSAx8CQa3d2rXaWjYT4HGc3juLGpi04k6G/rjZ5ZlfOvtEj32HJ
JwVk0YQV1H98Vyvirmt54f3gZQqqEohuXqjK9NX0rHseD/jnAoGxKfUBALwRx2rM
XBOKV6SfslsOca+hvazvmPfoBWQd3le6MQD2LsHJq1EBNjXAQyY/Ax1Apy+VJRDK
gC1mi2m91oUXRTDe9Pbz04kXSHUGy4gIvRiqWhRatPOwpJTYvOQF+fnLLnT/ENgr
kF755V7ZT3v6BCv0wMUtsgo7MU0oDZE8x1uhzENCtloqM04g4WMG8fXJj2ZhW5Tb
RZ5RmhIuZJb2Qg911hphEBEVrk+O9k7b1jBPLnyq2UeKF2U81iO+hCDFyv6o+pgP
vOoVbv+PSvvPsmL42O+9Yb89HJcOPp2vFnERmmwSDtAFIbf5Z1nr2Jjgshe5Q2PW
dOVF2iGMKGcsf7im/gAbm+tvVVrf5/QO56P21ElKIqXiHps6t9vpx/pCi4IrwctH
1KXexur5axnDkxBCI0d/oqqBRJft0bHJGuwq06BiubIEZBwSR/jgrW5gG3sG0sQ1
iRrYpWwHq2XmOALl+t+zoKcAxhvdKKKtt5ykJ4zLtnw+p8Bv90iLL219SMeo1cgt
I/0iY9XykHOE9z1pinpzfoe1159S68PbtSGSL9JySJX8EAKDIbn5F0EDoHphf2dF
98XBc/TTaEIhPggrlMXz5x1Ds9TRdtWErETDjXl8wY+ICLcbqEUwzZPg1PCx8Euc
4mrrUH++OIy6VsDlf7pMQY6ODvHy0y4VvnQGJaz2+AnjfOcQ6NuFC+tYZKiu/Eap
TD8TiF7qx2dg8PDZy/+Lip2rkROus9f1ssQ8lauK38e8sZHHI/Sc21f7BJ2H0eKm
OxUE5JiW5bwe1cFRun1jpRo+vT3oXSlfZHPJdWD3rv3fZXnam4CU3FBuM3okKqnU
VlsRKDUAXAPmcS4pYPivklDKbq47t2qjBRirE5dUGLIYicxsGrVwHygsy2siR3tS
Nx1N8l1zcab9Adas1q9YA8BVFjZEyA8VrL0NAmoDaOIwxeE/RnFbq8Du+8UiYnb5
1HvkcgaXsy8RMMsWEYeKSexR/QWQZkQ54GglgZSmnxifBKV77rTeepnG3Kdfb00F
v/yUbYrtmHXBt+2iXhhBkTsbcYfEBsL52+cjndeB3ED8QWRXSXzAfq3Xli5KftC/
dSbWKcs4A7t8T68ksHLEn11n7g5SFOZOXhSLOgAQJzCIM2+Wsbe06jYlgzQPM3Rn
meDeTegRY8ZbSbwaRMIk4lekddzt+28SZn5XuOr0L1VajBGUnKPFmhJJt3h7GrL6
Un5Nz+lVRtqxHhlFwkZUO6FsGyeWKDVHSsYTgMgxfTL9AkWr0napZnkUHzlWFbZC
XkTn3iaDokt+2PdJxzRLLVLTDKqmQWaIuT72A15Z6MJWZuskWzo1zrgqDpRDmY7D
o1fyET+bRWD2y+twsm0vIVwIr8BWnknQG3U/HXnKZL9UFGqIKERkgjZ+uyELxsWj
VjJLm8XSMpXfxRo2w75aIUoi+VLACrNccJpQSUIrWqBBV04ACjcZiPYAg3TaFzGr
TzBO3JHEWnom8BRMiaMMHNEYbErRaHukKezly4ZQOhQhb4GzJAy8qzpsMYhUqmpi
3pluubYqTF3VVNCcIHaIJrLz34+co7mCJW2MRNANQbBusMTiBc7cX2JVnOaGdZIo
nfnk5nhzTFBn5JWxHx9cIOKzxe8IuEWvEdJVMRHydPlmhcBjkWPJot7DwRQQnYpy
5us1fqcJlT8jm3Xm4J/Nm4A8VYA4DQyZZoKqYspAjKVXBBKaFX8icCvrRZ0IOxhU
oLnH21jfxfu1L8c5NejnOqdprCODZIpLkXwqw9MXqvRITI8Gr1DNUZK5z3Foyt9S
qGB4FRX5VdOarq2wleTwxvrz5g2BxQpTZ6eC45ZLS0Ke7ts4exIbw7s1lzimW3rr
pxutdn+jVU0Gue0ik4yyALn5SeaqCQzwJX+xdp4ifjTUud+hhechUQXFmAuV6dP4
+2FkVgFk7UpuXp+cmISVBePanuSewMWcFXvaBHGhMi1K36yaBzwPeRkpp6MchbRn
zvynLu2KKgdvygNYypArnXguCYHJV7rDcABvD76AIXAUaVrh+LZeIvmSuv+Ffa4B
hJvHBHlXZocCrqHPn2colWopbaUSaiZeMCUzKgV/2JamuFyIxqy0EqaIzNTA7r44
fUC2A2cdW0uEyPvlqYx7tid8YC61mjcxo13ERX3nd6j7qx/fqQGZeHjZcCQLG664
jCZsrrNFNp6eRFa2pJY0TXUUTpgxoQrQFTD+PvgFZVsjZCvs1yqI+gIfN+71wyDv
40k31T0cw40BTGhAU4AKOPm+xwmqgez+2ByTCYF89pYoVfnIRxiKrhPqm5ms2ArJ
isKsZYUa37rmuVJOAmXYoPlUzz10xmBhRbr2ieKwphrbqe2J4IVqwo3LHsoEIJ4y
DtZzDmn8KUvA9CPKiGWcBuNGmVRakuqM7UzD6jZRO21QC60paWj0OwA2IwtZSQkl
PpgtrwkUPXdUedo8bszyMxpwhaIk0lEUxfpK9h1/VbDyXDqHSApueABC3yDS0Kn8
xKed7m9Jcd82REk3jv5ZJWP58b5N4zDBs98c50HRGnxVHOH3PpsbjXN65/MD7prJ
JMDB9D3w9/TCt09gxcSwOy7G1QdlIksdg1u15RAGHfRziI3oiq5lxZOTQGc+VinC
rlVkqHXhNdvkArGwnXmz7bEof/yl8lfbBdUVxCWmDQqfKn+BxlwKiQoO3wwH4h2G
8ANmqh01DqzY9VtY44TBaXYqJOD7leiy5cXGwyjbxEguc0ktVC+qOdHwuk1P8ScA
EV0rWHzHXKlX9Qf/54A8RAJZvWRUfcCVL9EnJaPwJhdWelsbmCvxgYxa8KdQXqLt
tzARkV2MLoap+buPHodqQWG0R8Nxc8o1oPO1dVDJgiBiFaLNMgPhElIDPEBzGsRs
Iyri6ytc0GDf1UNjn18RW7NA2wpgw98qWNZ5Sm0j7GhGsgr0rWtIgtRSNH7eVcVn
1bczqzyW4JcMbXAACRB+S1zUYQRnkeiHZyIRPPLkeqh2x6Y7iMUyJsGYJU0jTrNT
kZUqjUA9G/fvyPEF371t072oz7l8SqJYPJ64bnLJqrRLYTSaOLHGVCPmiN2GWhy6
9nraJdR+smDen2r4jaRRUtiaOe4TJcbTFCk8NPc2E4oVtUNE0Oj6/czuC+CyeIa5
VldGUerd7s7j/DFtKyvnAtg1eGUT+cZZW4dHNt0DDSbjzdZCiFNH6TQSyK6F5fQB
uj9ziN12yIX18UmzJbYZjC7D051rw8Htu4taV0rPsY6N1k4w2duvuEuwrZedicmC
HA9Vw7un+2lReAQjr70vwS4iY4Cy4awFBrp1Pt2EwzBOv+A5sDMptvFs8+P3BsWc
x/U0aN79x0EXC50+fyxb9/QT3fVquui8M12xdpyr79FTFQjDs0VvYP/QidG9UbJJ
CaecyAWa5XXIbjRICNXhWESHTODf8mxC4jlClStcQ+qiOlvn1vXfH3EA4H0o6YuB
NaTMoequAyMLc9UVvkEhdZxqqfSAeRFShQdl6aD2hphXBGi3obZdCUei4AmMMlUg
JBiGlEX/bM9CAge9aiIOIC3gJpMsXxOuAhAiSBRBh8yINOPZNBIymscinnWOMKWA
u5BBoAFnGqlbfCF2+ceNig4sFPG/ympTsY5pqP/ELzGMXid7cTael4C5p1ihqTn7
J4hXdGqfmaJllXUXGJzXyIc7Jm43wrYJcTOyuwP4v264/gfMB6t29NchewXIf5s9
lb3XgVKXR80ghaZ7Cvs7cx9HXtg2fy6z6CQ26x8jbnIzp9CMZgwIcF1EElHogJUg
yyrwFGO1qCPaPbmDIvrESxzjQlgthJYzbmJt3YeB5MFUDBgUtMBw8ZGfU6pZFopZ
IwiuHoG+HbXAO7W6IjnAc1EDvMPObt0X6XkZA1K60Hix4z0YoTdje5+HNV6QtctQ
2hOxVLQgB9eGjupGTZPwt/0UznlEDdTarZODSqTgSIyQsnIdKEpK/nKQrdsGFO09
nxpWxS4avpzO4hEGiN9GWSnl8VKf/XE+XgHWNuVE7T3Lv4wQC/lC9J+AJ/Tx54NO
L42pRX3EWg/dzeRul0D8hAvoIPbdnVZyHBYGJcKKx8OPAM2LorIaFxnAwjuD/KaG
LARVKVSIbp8xVtt7hlzWOyi03pAXxlvL3BoQUn/Q013kUl9H9lqHr84QA/jgJYKZ
wDd9n1Q8G33krG5poOz+mMZRWUT5VOCoCWdHdlS4yVfmBzHlyv1S5xEd3EZ8EsXo
8tjOQ+GAcgzRaQkCcD89GUKQIA8g6pMNeLx3RiG2VA55JaaPndd1E8zcwaRfpELX
iwaiJBESECy0BwgtVYVpqn1BMPJmFw/Wi+A9EMcpczMtJ1y141OREWgWRveGwAl+
ElO5HOnk2soC8qmeDaChEE0MwYikzSr+QEBBJTa3df1du1jHwZ6/cjcys+WdhaLs
9VuN/AQxnRn1du+7hIZog8OOZAW2Uzvslh9ouZob+3dQ/ZgOkSyOwTxEQn3r7mSE
ujf8OAtOfneTLBWAagdS6w7kG7kl1sGsCvDTmL8KCqFux2QNeX5kJ/EqX3EoELOQ
INaGEIImOj5qmpDNhfIxL/j100gPZYEin/HbRMUgmb2Wr/lz4urYxouFeodp+EcH
mDvS4u1ATp3GNap3vRx40F6LK3WFKpNT9FiwqM7ccwe7Kpb3z8dMXlXCx3nR61CI
GIzjz5qXyd/g3v2/pfOtv8/LPNT6TpdwiRkl0FJboWgtb8Gkt+J7dPMeZmbYieWM
i3HCEdeSmanMpKjCgnhVppSagFUAf1xcJO44Sn4M2T7V/n9RqiPJe8YUwphsJFtg
IctDswWKUKqlBhaZH8aYRgdyQdmwwdMn5EpBxZQG0d5ULLzzyt5ZLs1MQMAAoqnA
QQGy1VvkH6YBKR4NMSE97ROj7Wj0mqObHJ5g6yvYPbC6btHCSX9kp4sWa3Fjwy5d
ScUr0JlG07SRNHcwFoTIvlZyZ48N2aDA5kqW0Fe6/frvm65qYKfVwAfQzyabWRZA
kO1vnOurCwIWgf78k2hK+LwH6B+dFNd4Btn3DFpz0JFaS2h3aRjkHQvwaKo2gGUi
OV92pHp18WKIb+WZLW+q578AOih3u6UGVWSsq8wamiirDZRwir5zPXQkeu3zXfJh
qoZ8A64JkICeunU5EH2ISV9StRMRnX74dQaV32xSC41Kw/U+4v6uf4jx0oI1+elt
8XOB+1tVc9p+6wm5oF/13jNs8NZKd4Q6vz1CSbd7DG0a9R7+LMe9A3jzY8IwYKV/
3l4KiobSQW8S1vYnbjiAK22rrBBjrOEXCwi29OFXIKWqIIXHgrWi3c0tdtB0lLtn
qPobafoEE39szgGdtEnkHf46ZJfGDoKtjBN3SmgKAHfZof2vlAhmapr7sVjmI1Lq
7nzduteZ+lHOZ0YWQY7aeFpJqS80bP8Sp+3ky8SG/GmbJZo/3e5FZiVaA/P03VfJ
qUj6y4o3eQ7D5+N9/J0NJh3353IE4WTbpo66M7jSxWhVNntTFOdKX82D6oWv49UZ
FzJS0sJryLGrroP21egL1xlNhq6Vk1NizTYe/qcL+jht2HTGJTez/V2LcjNGidSc
SoaWt+OLng5OdctlsAV3FTp0CpkFagsFTMzD7tblNja3L3Ue2hGGs3xSgar15Uax
1reyBPrm3Zt25neGgG74l/GeGGW1Imc2aJQnoDos7z/VODECXtIraL5KOKbYtJ3u
3eNkHsFL/W+8VKIJWSJQlF3AW91NrBKTIH4nLvlJ1zVlJO7F5nKeKy5AjoT4lOww
MMkPYdPbI6rMO0k0kBlXjxyvwt8U6CVH/dtlHmeWGzNFCandnf51j1t0V1dPMloz
LZeNCPIMpR7XRSRTmPAaRBxkBUq7NAAkhTOpDJfES1kEcG+mgCCWtXDVN9F/IpjA
XvCW8WuHkxXDTgB0R8hr5zo2zm7GsO3LllsRbNAItZzBq27QjhkhhELLOY9biNFZ
LJ6VNBaKXq6HtBbYib86469gPrVnI49JU6J5jPtM+OdCWhBcV/9TnhlMuDlq8F/B
NSqZetcvY3ah7rr8pP+pwuHfPAN6ozSnvgYsfGBs/mwBREcAoV6dy9Ff4VBvA2Wv
/Ay+07mv+TAVr1cXd/5lKDJSu8YG+nNs5cJ4fehUqIW3Kh23LpKk+RIGAzxpwF+Q
EXbpbR9NyNHxU8GX6YbjOiyvdcFgUrAsFCZW679WHyLFbldHHMhmF+xOUOHyt2sG
WLA41WRr+WhoUH1xBkJjVi6rXVPtX3+uSFrn3yPEmBCueGiRphMlmtpNATqfePf5
2+yjgORUnIT3j5V8eai8o+lBIQIxv/X9gd4jiOMlMNsathsNu3Ixltpew3sU8XKF
ihCL5sucyC9WzQXg/dHxIDPhzzdBx1vh2AX5iRXYdlfpH18VxE435gtEWbJo1XaJ
mR9zu+NXGqa2MVOsGtTTLfS2xy4VU35GRpw5gIc9u6wqiQg/rjjqFD7U47mLIChF
eXANBS2R8cn4xCaSNCJAGitw4PSjv0ptYJ7Aei/XKx5e55lbc7Dqugv+GAH4CjVp
p5yo+dd3lMvdLmkA/PRjxVNx5dvRNa/DOTJngnyO0aKHa+2fpP5rxkMGNHJ84/Rl
KeG9UTP7uiS4wLbV/pp3Nvxsqd7EG6/Rh4tOchANOmf11FzIQk9hAimmeK0205e8
EePpBTg+ACe9yVHHS5ZVM8P7vgrhvRsmEyyo8++J3YelXAvEdZfsmMLIfOOO8thr
AWO5SLy0wCpV3ZTKG8QuIhxQMQ40I//zkGMU/J5QHangZnGKniVAgeYM8KrzXgXX
wUevuj8h9rrOMUEnhYx1TKSEYh9TT4FNwcfA9DWmQTF7zWw7c3jdDe3zlMEfGTDd
24q5HIkbOxwIij+YCfSfuk4oTO2/MdqzRtw7tZvctd8+w18r9Dl8VM6hXyjTmLch
MWrKLdTkWfsCzlgiqo02BoTTnWOObmRY1zCClos6aj7hM+eNF++Xsx6lhyAb15le
R8tgcXsCLc8Id/HRuxNo8Dq3vDNyqnKNvlHWEDWsaEVuDh24m4rmgFfEarVrdYi7
dWt2iMrdp95YNGoON8d9MynNqxUySZ190enq8bLYdapmkz8tK2rXELeDOoSYN00H
KOTW1BTj9OhDacHPi7tmMxbl3wnn3A9QGP8JbJ9aiwhZm+vI+9x9G4rXmt0ceY/u
+6mVah0SU0lZzyOE3AtNB28gkpB3Jqc7HNc7ht34pwfHo/A/LLTaxINeckEvVwsp
RweRbeT9duoA2RmSUzwXn179fWTl0hJs7yaUpobFwH+69cr/Y7Bh/JEbHmvIzsAt
5zKtTjkkXkHoZszbgA7IXZndC0gLxFB4TtjxRNhqNEdXO3r064P0dnZYugW1y6ZA
9YfwHIKTo5SBjTJAi+HUtu+Rjroffe3TgRkrMDW7nI9GqU38vpzcNhKQ5pTwje6k
8SckMnwp9iYZER7Mez8UO7lEjEvKA5tzDbuU3EVO8vnBZDnxeoFgNpNJh3Lwkma6
ZDdnzVj3SQDI+VCjHFBIA5n6rQk8XplPZXeUwR1I1Zp03+3YN6XR9h3Qyq0PKiYf
QQ6zraob/WtWwK7cAjAPFd/ixaAIWhE9bUUg1Ug1yD4RYr+Hts8G4KzVP0PhWjJ9
mDwHoMRP8oRAJolZSaNG1aS/ubCTwKWrEhSyxj+nxt+lpdRgyq8TqddMGlYJTdpG
UJ3Ivr2cHAKh+PvKES93Ba+gdHOEnVoJg0VHxiIIFVq0hWsweodDwi9MYYWhwuge
Q+hG/nVq3XIEitBU2ULT0USwRhbYNMZHregb+XjeVM3TLKQtXLndLcjdU/x1SJyK
mSBZN3xrQ8GLhZfDzsW5LpjLdtWYrMlw88AVlAL1Q6H7qmP0/Zv0PaOmvQB+nqNp
Ob1ZUu90vTF2p2aF51o510Vf9TitWluosnOtA4YTITvoPZVP1mmaKoNuNtBs4bFe
9RjGpuZW25+uhMioZwT2Nnw4E+dCZUtYEwzupv14F+WJIUKC716EMN8c/B8yxU3x
Xsj/zrMcuyMSgyorG4yIcoEp0SQ8Jj7jMedEPsjGBDzVJiQOkr64UDOJ03x89Sy/
Bx52MZvAMRbeWSF8qDljHgbRvEbHI3GhZnkIbKscORq+Mgbwj46fUbYqLOSaAEzm
dKxoD/X1iEsQvnbUPf4b8aORBzDbnXssEKjSeTpyihzaauflz8MLkIE4/aF+0/+z
HIkk2PybZnE51F6hY60nca58XIH5+QhCBrvEg4x439eKOpx+i1ZNQIyc4r5FzI2o
7mannB2/XsQQe4ShAOGayTReGcwjJ4I6CowGV9r3fFnlpLyDcP+OJkoatCgJh2Qb
ltsvjrTIoSYk0MLco1097cmE4ApOFP3mzmxb66UxbznI4M1T3D4Lh/K5sf6bv738
nLXey9TcsqKiL8xqDZqey4kr79HZTaBWBe01c43zpwUtcPBgqWf5acoWCbptpxMw
iEJ6j7kWKy/B16PWow6VPiAoXjKEfBnrMH0DIwll2TrPybxX9G+lge18M+4SYYB1
7IwI4yjsTAtoYQB+y158obpCcPS1QdPBl9sDES7wRlJMOqk8FflWx5M8Ev/zLdS1
bGADlWa/b95iZUlZ/7jvXJ488L5Pg7aTNd62psWVVGiEx1SAxv2d1Ww1x8kv+nax
kXoSV8Pwuuaa8Pu61W9lb8njGP6qKyEQTWjU4M50IJ870tY9VEA4FljWFBaZU+Q0
ytI05XMbhovFFq1x59z/JapVEvdbT90LmwHCsBq5fukHMh8/edwN1qDcQKYADDnu
Cxq8oowQP10uNc6SccByosTV/qF79DhBdlXkGw97I4JepjPgxXSgVTIFG3WqVgIj
MYRoTkCDFxofbZay9aXEMcoT3WIVYKX1aQ7pL7dwHydvrz9eIQIU9aCZ+Qpwjy/3
uKb9LYl5QH9/YV1c5EOOlny794QCLpLOJGgLxrPlBJhKYgfqPG+su4GswF/W2rP6
/Sv6ddw2tM0Ou+GdT0ghEVD23lvoR1tPoH3Uwp2MubzXoJ67m7w0KkwcOTB2tF9I
2m1ggs+tPzYwSjYjFtGjRRha53F1jmyW7PAhDTyWluvtREdpAHIfgBRjEsKrhzkr
igpURNy7C4/NbyBkGhxvb95WUk76fnyuHvVszBa6e7Bja3RN3w+sb0S9nWE4YFRp
s+JNqKGW6QetrVbjZvt2h6+yaqV1AbjDBPi8wfJZmBkbiwALk6nDmRE01mtP9GDl
2nyFrrGtB2Nt5Dfpc68cZoQkfV/ba8LkK/s26K5Uype5vchKwyGu03UrOZTJ+sLv
SuQOvAkCWzIHxORgDJUYpJI58IhtipaJW6422heLSSSevhcJPLOe7+kIFE1+eeAq
KSfyMJOZw9Wc56WkV+yT0cE6q9LkZD0P3GNT6TgZKPcqoaKAfe++aIwy83r0DIT0
Dn9HpDrR5XxipQa7V68VQVpZXpa9SA+RR/JK54Ql2KkcaXIvY463Ef2hP9XHyZvi
s5XL6wMOxgLe5uKuOJqr199Hm3L8hlgNUQR3evsc22A4Ef+/5ZVsdTGV/fR/DJSZ
p2xso4tH/3xPpSr98P24SqGMalAbPucpBQNLtGpEIHvYifjNXuPF/P7i/HXtRMWl
W6R9SUu+GMBtyuHf/Vq99i+xg5JH0k9oBmPxeDx1NXpqOBJoz7Wx1bn9u92YxX1T
vvGiSr/Mg8n6MqCmBD3J7s3urYQAzlhh7R0AJbwn8qjE4F/H1HopHLn8Pu2AFYx1
1K5Q4NFlmT6HSqtLnGiTIUjme6BLgBnBd2mhIKzfvSPmbimmirVWTa7zY4pRwZaG
0aK3dW4eUb5gPRuLLUN1nCI8RFkQXAAhnf6aNGE2BuR9fw3vnh94Eijx3YqPbASY
DZVoyDEUqf+I7iqOGegmSLbkOuB0b66aWvfHnJpqe7nnvOYeuabYExamCnQUoIfP
VDGawax1CA1FkcIUNItWCFWLemnveOUu5mefZhOCf28rImXzIpSpcA5NGJ3pCLiq
WCsJghsKcq5RFfuAro1gtke1Ug6qv+Mrw/phYs6Ra4ItGSO0fujRJUJtjVHq1pPQ
qx3hi1OoEri34BSIkbtOLMRjUffLtX7KkZMqRPqAENBZkH452e9juFtYKnVChfbd
2TakaMerjoy8fq8cAScFKndEF3nj5lWxzRNEwtmBnsAnoH3K6uo51C9LP4XYCnvG
buXDxwDedUY1znc1cRfK3nCRTJTmg5emDzbOxxgne1xawPoc7DdTjydahmOKhzXf
YzgeJr9rBLeaFbbUCSNNrT4fQhE+Pnysgf8n+am7dDlcixm7vgnes0X/ZOIZopHG
bFHl7C2sIW3KfiLcKaLCX1xRFI8T6N539eTsO6SA/hPx1Pxlt6nB+dMhJK466uz4
JnS13ICBnj6MfrYfQB5Exj3hvpXX0uquWdUFiVJvjvggbKPKxGo2bs/2s3cGeqRi
B+45MVRi+m8ipAwQ3SdS00rDdXgee6VbXXDo3cME9cXfMGpBi2jcQ2RKMpNgZ/b5
GSDvgCZrSNS9k+NLCi7dgg3sN6RDMbcmHSsavhERf2+eJ0zazEP5tyMJxEpXssVK
vSc+0xwb0WHkp0zcEyZdp+X2igF38ch9Cn+19fqoG289a1iSC4m990ifiVb3ZZgE
iCb5pHTEd9FxoK2C9VLguDZqCa4xrUdgQZ7Z4zKOSIlF2kWEFTz0zz6EvIS9IT/z
QNysiExNUlklY5hGaKSVqo5u7rAAawTG50q6mGVizJ94kDSDOgq9rkX8W3Gfzzqs
ftTL6Oi5gRq4K/y1ckTdkcWKveKGiOLU63Fa2CWL0mWT6w1Z5Wyk5iZlrfRCMVhm
WmW6LwDcuY18DpUJZ6B/g31wvRzlabsLePQzFGkQ4SHuYxc28I6f3It2BWQF8J47
ieHhnVTKO2DRxahdbjFaWojvqyOS9L9MWR4BKMhKQH9j5s3CMB8JPb/Fbie+CTZ7
OeZ+mRutihSaDnG2IpBJ5eYQNZGaEddObDpFU7rBtHzN6ob/vuCyiVOV3nlOF5N8
IUOcho030xw6akmXC9Cu/43AYtsZp5DaTq6VC5H5lardJ/nWSy2ibHPGLC9RKdUC
OpKvS7pTtCc349QcbET+7BvRLoBDzPt7xpd/JDQxEimMKFCE5U33lsh00SqjS2CB
Aov6sZ+HBD4Pcd8EhunocAw6RA+O69nflhjvXgujDfGpKr8ylnjljpDkISXH4b10
teH4WIrAPlJqKxsFddxJ9NTtjFFoDg7IZSv2iIAZa8uUjtEz+YFtLFpVGslZnuKN
aBnTLvjXzlhLMfRoCUYGIb5AP44FsmnQcRwzaNS+x4rxLRoA9P4uLBZUEEsmWtKb
jL7LlRFO9w9HiEzy+l/5ntdioQyAf0dDoxgL0QCnGcL2HWDvTYPrdifuWD7BXOK4
MKIwewi03F/pncAYZoG8n1GeqmdWDwoUB+7F4nj/ZEtn+TnRABTnwlXaLZR7vyKU
3fzvgUbLIxdK5efQZ39dH+z02KvQJ/sRi3q9Aw6aQYOvVzYhQ8yV9MvIucBBI0uF
vn7bTlFo6Qbr7Wijro4kXd30/Zx1U3t7meaf2YF7ppQJ6aupYQI7vHNy0sQSHUkT
sEyYtjq6h8jL4HeaZtXKVlJNsvmJzY7824HJiep9nuQnOIM7yR9iCJnPFAxZf2aT
Ik3zxLyLJAHJp0T2Pzsa6DtOSR4/6WIUd9aBEj0/6VENZZMBYfll8z8Twik+DH6x
4vv6DsSMAF83OsFtdCQ7t7RNof4q7ORetgoadJHbviEOg5aGaep9bFUZ6uFC94iW
CU/h0ud84hC5tqV7LszB7hsCtEaPI+YSlUCKxu4kMDlGFmFSiyGr32ykl09QitYe
YqgfnUqDvXzubHzCapLwVuIkloJ4CJjm97KnS9pESOM3IjooHvrXcHb9jV5WbkyK
8iYuH2BlclWp+De1BztgrU4uGReB5R4PPGBJbR19usleK5s5+jwStm0oR4F8nAA3
7XgX9GMQhwndh4mFoj156wsnRR79Xbem/raApRxG6197PUXQjRrZbzDTifl1O52+
biXF0Lw6V3IF8JiU6W643Grq9UYB43kXnwpyPds37Ko8vC5NZR6IKAziCHBnvEnm
HaZlt51cvo7RSuwtOKh5imNio3/al2hAObkJU0UHCvcFTlotZ7JL6Ha9eCtO3uLY
T9FLk1oxv3RJG6f1k2QQaLTQ8KE/C4ydliC0sKOb3JIrJoaYegzqVCIHccDsfkhn
oJORy/MufzN2cIgw8qjX7BNIYYMc3LjoKRAeQO+WKsFL8LFb9msSFuGoQSP6aU4Z
XqDblldRzYUaKqAhWeJJNiTa2Ovr/z/IxDMAcJQk3ridRffP9U4h0dyrDDq4XsJY
nKf4jVf/RPY7zP4DiVfNVejm26TZu1H2DoTBhyDcFwc8FGxmiMvo5JtPAcpEtH0E
gXbIRXzUGtHeNZ7GD3V8/CmKMN6ObQO8lxYquMdOi1DPMlxg6IqX+9hI0ybP3KuM
o45NWFh8yaLXcM4K1jveLSWd1XANfJ1H/FXWKGGrfkCcwBENy35OrR/bl0A7kISL
5zo2WWgYYLEW221n5Pg/PPr42hapqdZXuNat8Tuy/rwhvSyStJuDudoE+9QFdyp8
HGhXeSgoUMqo+Q6eHOPPn74sVT/+IJ7RNzCQPyXMeSC8hGFUd18CcvEDUf9xy8Rz
1z0Q08Pe3t0aCTwnlooRYVvQPnsPo3lh2NSN613xOwD/+D95GjutDxMEhxX8T1bN
kvFuiJVb/V1x2MUEiUhwoouweV3IYW6RPBihuQXCz8RAswwgOlteQkclOc3X4wac
x1fAdSsnkBMyoNFQ7BYJ9JQO0ha98JeH1INUPDZ9qZuyINYVoApC1iDndcj4t/rl
lmRsP1EHb4gUiPaaANgw1ODaGvg2IGckNMe5XeKTfMQQP0gSw7N/QJbWSDQbo6qs
d1FNsyRwKhd9ywjmqe/jh5i70Y1UiwLX5g/Q7vtY0quygO5DDzGVFwh4QhNtJJ6/
IU7fcgR7PiNATL/CAco6VbGpkVVQ8vyyGwH91MZrbAFBI1kxD2yjexir5wCDUJ/B
GivwNppF+OnL7NixGcPBgdgO68BcjR9StLsmo1hR+Er2kVNdEnzJL+Zs7djty3mo
JlncmxZ/kByJbcHv0bbs5y/TNZ4mH0gZGL/cpGdQOjQCUjRq5Zkrs7mlZ2FIhNXu
j2oPwV4qJ4in0pObWgG9OfXnC4ElHxX7J66Ls0Sy9sZU5r4nZTEGOvZ7oIKKhBS5
Vl2AroGOgYqMv25Q0HS+rW5pxvp/Nnw8M/ds/5dI+yS67miudJeqMUt03nAAQDaJ
/1ylvZc4jipWmgnPcy91Zmsi1fSKNOzdP6I9JKyjBTX0TB4Y/+JEAYeIMyuVaG1g
VD4xeeVOyCg1PlMpqidEBWsl54zkLH3XTey1i+NOXiTeepjGxx6C7AKV9rJzT3Ul
175eHAvxsEVncV+cQRCBZpavFhxUKUiQ38PlG9UZyB6BHiMnzIX7Z7Y3vG5fZEef
eon8Rf7HwluVoWcDLGRcANQCWjSArBPkahEikDYXYPkmeTtq4vsD1Cn9xk1NMGvh
naY1jXYH+ciScjVpFiV+txtU5EIfnYhPa8XG5orF01a5iJRK21yrMhni8x0vPdzx
9VUE+TwQbtB7sO/cVK9Z0G5rUVufoH+RdSa1lzsrNM3lptHEbm+BUVMHJDorvgjh
oaYLtpVLfc+xrKzcE6ZA7u9Iim+icx2njSe37m61pvs/qP9JvBX5XgXBcm9qPYd5
zd/CgBiiKr/Yj8deFYdvGVpAcK8BOq9aGCGsm/sEGiMzN9Tk928nOI3YDR3H8CbC
ZWDyZy3Rw7SCdweqgiO1Hb8TLY6SAC3quGnYVV+K/vhM8bSl8VjuByGUmzdWJZoM
3Gpt0sG6Rk5J910Eg+CAAik6oaLSUzVd6NlMZ9d7ETgF3Y3AJ2VrcIow9NgyEDSR
ga/gKxwNwA1xgE/+dI17EYbHINsjsDy8Gz0c1+p5r9WOEEJlB5SfkOA8CpCDKRqI
vFSkmJ0+cXiA92fJKjXFXtFgp6X2c39Ct3FsT1eXBbJvN3O0gQbf5MBHPwm7AAuc
HftANs2E4/lv73lvYiq/x9rTU1/b8UJSbDIjAGXD+qxtgUFhOUUpdLatI1jIwGQC
6WxesA3Ma5B/GScatlcMFsEtaOBTvMI8ejcE7bEaX7TQ8Z/jFgvee2AIJO9ywCmB
aO0sFpaUhKb60jpoQoUC/4ULdjRX30HXm+uAXCs8btsO61Wv7JfUd4OvKvFndgei
2dUiE+AixcAsdKfvpcbogn+aqwihYBtg1iO/GemMyex+/wzoQw7+Ku0LKRNIacSV
gE/DYW0LVARjttyEfVsPUDzuILDO2L2BcmHA+wox8D1vZY66b/qpxMJzCyE9sHiI
2LvRzpcwxfR3L/a7RG+npUYnwP8kyj4PYxCsYBk+cKLgnNb9boaSMZ7yZQm/triP
6DvOH37Sz+hDpDMPnCxWZ+6La4zQaXnRzPWpmB5y7EOmK1Zy/Ut98/xTrO6toBlF
GINTM2F5vnTeYxosYhBJhg+0SQmSxyU29aT0+rgxeIzdgswq5iVMuIY0gw4XKdG0
yLXVEN6JYhfDYei/VgT6Qt1UZQkkpktCtv0gGVbKDzCLRdxnWu1aYlyXpiH9loPP
P5jMSQ1SOnFwMIwb24xEsQoBhz+NCxW9CYhqLDCyTz77wYEIocW/eXxinMaNd9Ev
dJ/KcgLl8aegTEuPqE3sTX59tiQaJ1jsAc2I2IUms2qtxLQzDRjng8VgEcq7H6LU
9rfnI2rmGXdSgsvIbRqyddYYI63PyI6qeq4CkujJbM0CnuQPwf6is2gnvJ8LpP1X
ap6UquyY/QG9LGmOMNc5BrvVwLKGYtBI58gu+7ugiEv8lma2zVJyWNHO7T0/qGXI
tZQgoEcDBgEu/ibRpydPUd34jxg4XwORdI3p7NOfoN8XYUxTsVlilrhtQCLK/rBX
hZyqMbjfpvn/r5SXu/RGoMcI54dnxZpGcJ2+V4TZl80v/N/UV+nLUN2x54FhJj9K
25mVPvE2fBd17WjiI/q/aCbmTabRRnYiZHYzzyy1UCzfTNThpz5oZ4Dp9SZK6Ka0
XPz3GCWjGIdCAgr4SLMWameB8rTqn06Q3AGNTlu86rzg3t2HNjjTdY1hNmJZkM0W
pL2X4ee1UtK3ticRLe8/DflGPYRd1k5nOcfjz0FG1xL3yrsJflKAP7rh+B9DPcQY
vBseL9aMfjuTaq33qFVHY85S9I2aT/CX3Jll/GA5d0nN+ips7kVphbXxakVPpKYe
F7SsFS+QkRT4Ty775GU3WJHQFpnwl+ZBnRQF71goyCsF0GpbVM2Qbu7EOEQVFw23
fhUCpAqujOem6PSjiQeOkxKQy5GXKYwtTXNRtnh7lhZPWnu30dsWunNhagflTICz
vkUXI0PSR3t1AebppHYtBhvGDSFD0/BkmPZMDwcmyrrFVfUutU35LUQjA+pR2Ly1
0/RNE+yjTDgvUVzaS15WmrCxSkXx3LKBsrEDmkMjTBKhZEjJQRM0RoBxbcQHQ5pM
HbTL4IntzVcLXrbYEF/Zsnu/6GdQufM16Uyw74FWuVOEzeLSaozK77e8HFqfQxBB
JaT4WI3kCuzBewPKCn2oltd1he7kXoQQJTooEZNhu6rUthLqOgUogKMiBSa2BLgz
xZ9ldWM96bNn4Hp+JQAn0uZa/qA7YzTx7TrdsJeg9m6MUHYPi4IqV0oOFRQgM4J3
eUO8k2aGdNFZHFhip8vkpeftwC0VRJRWNRiuzxQR7qtlrlM+nE/jh9qxgFDOiFAF
J7CG578XIJQJzCQXwpvlMphOfxk8WtUwxE1tFFtTNDv4YBzri/6fY18n5p0xiBFk
mTNBBj7n+Gw3lFaCge4F03lXukiHkRiMwvM+lM9iCAziOY6unW1Yt/vkjKV8CjYv
XlzblzEcc+89ScaLUlx2mXd0vcxTjbw4g48eUrPgJ6S4cCw2VgFPOcWZ2Hjhr6w+
w8Xh0482usrlB/dzpfazDsXvyP49wUXJkl9u+ZH8S1MRyqas57b2pNCtUFYCDZQ8
1IcuVNL4JhoGYuF8rh02UB4BItq3TUJtbdR6CzJpU38aARzBuUq8qgukYBZqsGus
WqCK0YKhaskjxTbt26PqYx6BlcjiXcgvIOWQ+KijiG1Zp/QIO7TyxJQ7cHzQL2q6
8PEYSUYhXZrCK/uztwMnMFjX6iAm+493KFBxWUhjMJ4B3Ftiw3S1UNeIbKkgvEZc
4ZlBTLv4Q2+mXKbplKNUHxYwOl0StH/ocKHjrpSMJWMskLNvFEHuk0oaU184KuQP
s4srsaWBgTuJR727RGQ2/r9NPBZaqrg1DMXJqU/HK6LNmwK73eC/uRrWRUZqVouK
YarebVTdvG01NkJDZwWwlg8rgRng0blkDO+XJnvMHXrmBKxMP9NW5VRUuG+pdQbJ
PlH8cLzLokqmYu3DxhCYKf355na0fMq9bF9zH6rHz2txISo1TNtss6LZaif1p0qP
INZ1pZ+JwShwdcGpD0+77TBK9JVi6ar/8GoaetroOcCE0W2UROym7sbF+CKW5Dl8
Xwbr60Ne9sOwgNYMzV0OcVP190F9U9MEf9bdbtEbRGmXfta3Kf+W28AP9w3Ycqlz
YMq5/JcghvXna4s8Uujhv+UT8ViwMsFKS17r0zvpr3a1hWDjNMMcVAw4XYQFQBkP
8LkmJxiPhdmYa2aU0rlF7JwtHW992TveugUZrs+yDU0Igzq9SUJY+iwq+wDvnbIs
BTyh70KHIeO6Svsgl5Kl4aKxxgATPy+wj7IGA1If+uoreC+s7GpndLNd8ARS2t0n
LSu06k0Osy9Dmc7ixICfz0CjkedZXjL3UMXVItZD7ssg/uZ1/2JwMrwH2G4yDMPC
AxQ/5OVVIbH5JVSbVB9wcZrC4Lr5NKecGYsgQctgt9wylWYkwQU6o1MCDGjsDUGo
2EOt0VYIsQK5nDPloLcatEjZn4gBJUmLxFO3xqGYlLK/gDzDzpD5t8t4/Jbr5lTG
D4T+FjmImVK+KFJyoZnuN6yy21Hm+wnavYlE9nGO+dKYh/QNhUbCQyQ/NiYOcAPk
YWXtbuIuJrJ8WWIt77jlv+ZvsRE3CuSwSHUYTlwAsjE2z6LI38f4O2Qw+0vhYNUw
q78wkekj/zrnn5DAJM6rYugVT96QCuhWNp5+X+gNmK2Yhi8kJEuIhb/d2sn/Mm2e
VqsufUJ8R/H7zIhQCpe5bVd7HcYgLfZsVhXGL7sbKrgHjpU6jwfq3kWyEChFnZus
YB3Ij9GXHUuwvH9thWewS43NUH/oeEDU6P2O/duH+puVyBhIXFS3vi6fWn5uSsLX
/ZJYz7VSweB8HmFXZ088OeMrh8J2lf3Ko67e4RVVqrKJ9M/l1HIQ92mY9MK6Ysr7
pS2QWgENc9QO+tIcKqUt8VNR43OGKWLXdgrKOhi0/Whu94yoHs+k1fwIoUy/Z6/E
k5kodICdSnmEMp4LtcAfMUJc+q+SaAiOMOOXa493Fwy+NcUWSR0abRgRWKM5GHfW
teyymaFPwtu9b+7thkpxh9fh8pW3sW54zwmA2tfUAQiQWayAFz9NiGygUKIMa3tf
T4etevNbPntQc8xktn5e03pFtwP8fTaMecEbW53TypQGSf4Dp7XX1YAwYSW5FI5Z
bYgv/4ued9MGUtqKEMmfxzc1iuJ2O6d6EqeUVljTrHo+kTAuRVLncByzJrk9Jz/N
V7K/E5SJZ/FoTo30cgzA15P/WAfBgS3TwfVxIaEJ8qhS7tx6qOsYl3SJalJGKGLc
ZWj4KN/FAjyapNGtkUyh65GuGYYTZ6KxaMEIB44loYlYzHRUETdQUpyUbZB2R4NC
zgClkROxBSvCkZvPUbI7wdAynUh18MEqB7IK5X62Ul3djSzgADtwF75cO3igMiUD
xURbqSofcM/obiSN6kUmg+KBllMbatszv/q+fgeOSwVpNK1ao346GzApFazPCoOD
TFyxgzT3ex2rs5ggVM3XzJIRZ/fUKqlfkpDzYv2VruAVxRgPYosbcjLpWM/F6M6T
AUFIBek4Sdu7ZxAqJoFrtiQDx7B1Uchgsy/ee/3zEMgehm+1gdUpRnRqGRA2+q2g
jAYMt4fpsnKYCF+vaAwRy3WDhc07+Zfqp7eFCJGL8ER9pAg5kBoqhK1meG45xtZY
CMUuNYIEwfptU4Y1Vx9mg3pwe9lEJtff9dkzR82lmZJ686C7xoQgGOLHuaVPeC4t
SgMYKBMToWDF9bu7ZUQriYqppzEXA+L9bh00XaziW08RRRk/bF6aQCMK0McCc67u
xpqgxvXkaIl7rQxvL53qeYzMF+cLJGZ19lKfWcKdkOoXLHjPfa6EHxbLCSiEhRBL
dzgdwhkEoVZ8W4fAU6TrpIxlcDEfu1DMd8L76fDxSuus0ZqD867AktDPdY4+deh6
m1Zs4jNqDvLmq8mEsxRFyPtMLG8Q8omaadmEUNQEl2ijjwk5zj3Rx4MN0my1iI+Z
KbcC5ZTxyc4bekJZ1qcJNK9VU/6ebs61eLEfSwhN6oFCp8gvq2v55PnePkfgHur3
eVlPTh21gAOxfmnPh7JsfPkDVx/vm4G6PlXiSUWbu/eftNVlyxQLJ+S5wRgm0S69
vRO9SOuvRzBPaVuONEOZRUhkLA/2LPA4vpFzLQ5r6Sj3wULfox0F5WYoGyCBwQqv
MQQZ0STzreMQwu5W88tm+nyqGtOlzc+tPr8NymUJwJAIWINgpj81N6/R7UZooNlX
zrGKS5cBgR+ShhrD+9tDU4phFoTCQ1NpBxFwWpd1tXzi65nTKiY0Ri6ABnypLztv
ogmmQxHPBCvqOMII4JG8MJ6Wy7IoM5RtEJJYAJ8olne8hXptc1CmvLPXoRoRJiwV
DNI3pwCE7LHbhw1mjqcBl0xeACfJ6TXoZoNrZmAY3jhsicMoL03agp1JBKbTy8JK
QnmAw/mNyUubXeRS1+aQ+2pXBCBQs80VuozusCbd5NCd3aumHvKx0BwfQRSGSqkK
bap21FHwJeEGJgtkOxffLofWt0qzAMwvd059MEE6w3OC9Ht7kjFMPoDXEXQrVjql
B3xugl/jLB/S5aENdB6fGNVcoc61brzUIm8ohjE/rwxQXveGppCoWnOVAXj46UPm
Ckg5T0eJuE7zUGbHsX21uARqpogf3uaLIX0e90vYZGmhU5LBROT/zKLkdncE0Fki
ZP5Ie6984B3KP0tpU6rxdwhXDrusfw83fmj6WFtxOiXH/nt3GgCEk7Y1b/QG8uHL
KrBS1eMUw6Hcj+p4Q0PlEjpWDxODXfe7jTu+ysrxk4kINX9tg0T4W4APPc1oIvC/
FbeBPp81GTtR4p1AZjAOm9fPM56qamYKEEIHgU4xUBOm+7ztlozA2tEa6Ywg20oS
5J0iD/mDmuOM3NYUflsLnIMoZVpfAOPhzFlvMvQLzMERsex9SsavGRFTDxccoHw8
csEDjvEMBl6IqitvSrSHznG97u/tvo2YMO+aFFGNiHVE9i39ae50lHpBh5cRccmn
sx0M5XcKRbLrKqZ5Aysk7xiAg/pCw8OqTHNLY9NCpmNZbiMqXWumySGW76Pcgas1
fx7shc1zDVz72UpSm5K5bh8A5sCqTXeXzHYxdkn7go9Uqpwhd+SVb6BogZlsH1w3
h3Y2lXZob78g/Jle3REU4kyWgnUDps41LWpkNHuaqxFykfKIkneSZAbevj79UjwA
nUwk8XPzTm10sljfKWRRe+26Mjt1VHStKDnG+YQf9jZ6CWxjtvCoUw2kPPU/ZDof
3lZkqNLU+C+zttuhs44awTsXBzT+ojY6JO5SvzCybkk2RmWAp25p0eiO0qcDJxHv
p9Dufu+LZUBWR6Gug0jqCy4cqlACqMEXFFL5g/Ib7ABRjB3lA0LFOsDhPXMbPRs1
qeWzChMxqE1NpFCL4NV0/IsM49hdQixXo1xKbUm8mbQ8m+zrLbMTtRtpojtLMv1G
CerFZpTVDlZyqVFJtvTIHzpQB+YtVbLsjo/d1e09qPZVjU94YJCs+OyIVWooXHt0
OnyT6hFH0qLThPrLDqOxTIZt2mq1cxOVfrhgVvey4+3w8xp5PHNboVfdyj7/k+ds
XnwQqAlA/c/i7kBN1uaK5wRIgAB+ALSefBxjzzyxVY/mwdKpMxW8LpPbXCPWfcGb
t8KiTVCSIY6qLwvKRX6rxywIsSnPSfrdsNjJXVc1en5T42D/GIibBWsZMk+r0tVR
WilCNDDLZw+OQAzFZDnsMsGZpbm9zmUACiQ6gUKkj6SpJ1AxrYUz3CA4hf6YgLj2
cGDHpmsJ7mr0qybIC/2JEUk036yDtgjmfDiJmiHa3pllyBMOo2/ppiKIkM9Ue7eL
9iXeScpzdPA1T6VD+kcVb6aaYWXq/+wWB4g8HzP6VE1YdYLGCsnaDa+SaLFO+N8v
klWK0auASAdlw0Fwpxe6N/CjyMdeMphBNh3cgsvKiG0aR7iBwQB5nBBJyd8WG62p
fB+LVoswUt4sEBTZqUkWCw7WHiNCWYg7BUMjR6jGQ2yoJz/Ho99jg5ZVBjsAqHmm
Z2+gMnramc2D7/+P+yRuPr2jmMENmVHXeEazbH02a6sVa3bipojS/gyg4TqLmdAj
khddHGP/yQq1zZMzaserDuf6mMf2It36uI7kNdFkRcHNRJQCS3rtFVBAGE2+HLHR
pt7//2GcUx7qHUE3q8FTZ1haOT9lRr2PXU9Zt6RLxHQIpM4cC38XmzWcbUMyURxH
d/KVs1AAIWR3RXTROB6SzC4meeQjEv/sZ+PYcQ0mjtJZ96O/xHab8W1WLN4MJv9I
Alu5evpi3xh1oKrmKhN3zfau09+4tRDcMp/BbcB98JxGp1YNS7bQj/Xz9MXF7Olg
29TQscEUcUZ/IwuBXrp/HT1Uv1t2tSIPDn1iqYc3UBKYYj+2j7+f0vPjelrEbArw
m5M8qo6HZc2KoulCBkU2t9EdAxuLwqMfW1XlgQNzmDA25C54KndTM8M5MBM7EM4J
kbL7ExZ+AH5uS1ueUxVFqOknu+rTl9nxnEpfkK2HkL8cmxBz1f0xpg6jdYwYT9Gw
Mdfyo4WH6XBEkurz0GID4OYQxC2JWY9/pggJ7SP0Wly6QD6cZoi+jZDEOo4uVPa7
WHHUMzL6C6r/GLNSgpsOtsy4pxXfpBcOFTqL1uBpZ5vRKSrrKjisyQXYiqBwwPht
ranM29JrcnbTowczRD/BtfTzKI0kOHYfGENovIKtIDBg3f8cbjQUKCMTesa7RXu9
XJc/Fobv6uQxZfgAAL74d78plDr1Nheop6uVr8oLkYdrCemvgZuZT4BweRsWyw4a
Jo8VTDAjmcmx1Qx9XzokWDp5D4pNvKC0LiXFKY2X1Z15re2eTKfoRpfYBy7zVU0h
sCnzgXUov/ChFicxwoEnYMloX3D0fYTQUKfl7AMu2OQVw1gut1RoxFBNrwYOtvH1
ZZ2dwVcMEdb2LK+wlbRqFWi6Cwyn1fA6VtlafuC6bKy4SThGYx3MDgddwh6ZU86r
psjVGP3LxYzYu4CF9rIp/GPJOVQjMX/+WzYA15tLBVhut1u8uvKE/Ar/OGU+d1m0
9Q5oQ5HBRLns9YTZWfVwNoarr9AtHF7k0QCeLoelh26zrWfCIs++ISPiKABiXzs0
cA3oMksHJf4/xj8Z/u0FcT7NRsJKVcSTbIgRmC52MSNHW8QaYKtN953mVEV7e/1n
saRQn698zhG2+3hUt4SSVjj9+T60saxhvhO/GeTPjsRdxB0sm71PTQ62aFTMTyZP
ONDnw2Wt8r/9auxpGES1yOx9WMZ644ExokcpdxOCxgI3y4PRQKAZRt3sNPpqY3lS
9utG7d4g1YNLiBh5fhWURY4tBC/eAxVO/Fc46+KcUIaVYJh7+mwr5tJVFz2/U+mZ
FayTq//IhNWJ0WJGcDbr3guQGMjTixc29A8DZhAu4OHn6iN7H7Ps7KPOAQfHu0xV
Kk6bVwAsR9AEgpdGwMT4C06nwc+FT8FWmgxVpMKHnthXF7A+rmdhwHTyngYjap6C
uEbIK/k45+w9vzyx07/fJ17fUPxQf/Dm41C79H2vHYu/AOdKd2H4s1v/UQTtLZf6
MTcEIhUvN7MWnxkIdxl+t02XmVHWQGBhSsPvdaptK2q+8PBWoIOKe/nbZim8i/Ho
OQ3uZBJTdbWEUgbFYveswd1on74TX0fzeTnUhDPGJFVpUKCw20eAbDVny1ND8dTD
VblwvN/h0nRQlP01JTxydv9JN5mdDLlAA1eXqS/0ueHyOkFZmi+nEYWOeNolEO9m
7yvC0Sqrlk9K1MOd6mL3CRvHrqdBBSXg7Dzi/bv1+NrUHROG/OtG7SLYf09kn97V
kQM+nWO04SVgPeJatVQ6huVNVU0HP5pgTYt93ZS82c7mG36q2+zI4n48vYHhgCFV
5DI1L/u2Vzkg4Bvrgn5uPc9vCRIK76w7p3rT/L2ol20psHnrHspDDzSeD4d2kc/o
9lc/tiDheFkbJGIc0trfnXC39ZR8TGlMxVg0rJ+xpyeSB0v7wBxgjMpZOSiHN+DZ
XmvRcdRfiqpqGvM1y7Er6/EcmYp6dfu5rcN6YYTNnDMf9hVCK+2G5axrrH6jy3V5
xKXF1DZMFoZy5Y4Q7lR65SOJbE3P3/S4pKy8MuaL8BtgHBcsC1m/HXR1ssrTweX4
RtW08xIT4/XLpyr7facIlVFDnkjZ5qDRtiZ6pFrHG2qVOZlQZ1vsS3Tmrm/a9FtF
tb4IZv5CBqixM82hS5J0HZ0CLyeSXfyVFi7YPsoHpP2/eGJI0ynGE8fQMkUGIjVa
BglW83NI6yXAtwD5xKtiC4Q2w/yEjYKGCdjLskEmirxOCG1BhOU8g0MTUpAfbt2s
apepWcXMCGamWWRCeLwbgUO4i1e8Gr2F+ElmzUKlh9PMIWgNBc4ON1v2040ZWnKi
23VOptFXmPTQEcjDtAiAidTmWfhUwXvomixNRkRSdgXAvHgNeRNn/+fc/tiKF7cJ
mGgDG/jfsRu1LYEbQMj6ZaU9LboE+9wJJzjnapzwz6dXf+whRmYr9GDOadcMoMd/
b0BhjuBWpOEocmnwtxJGXzkh/o+fGl5p7uNYqo495IqFqi9GtEPWKQS6psfACabP
uxn2NwJxrUbkZhAyMZLoEN0mxdQMKwbvz8m8mGS562SY/Le2WXipgEvvXLco0n93
vaQ2MJUHUj/uVORRkj8m7zkul0JHVSXz7gVecPxJR5Ki0q41KcFL/VzUymx13twi
FMQRTLeNCreF14UWwB9xg2A39KNAdf06Z2MQy+apoG7EUEIhJAl26Q+mI/w19znX
yeOWhyTVWe3xe+T4rqAMosfMoT1J2kBPWNxatWU4SohB3zQLpu6eepbgm0QjJWZ9
duwZ+SrMkzDOrVjBFIx2ToSs7kjTcLUrV+F3/WmAIkHUAYXT2CxRkvoa1IUAxaS5
cqANsxAT+roYL5syfDicsRt8T0WWy3qmqmOgoGJci8enPRhoszxPAskioDMGYQ/K
36ED7ydB9bve8X09ycpQP1CH2YwVgwk+IhFGPHfdIDZvNdWGpL2qzjJanTVfzBU3
kfqkU3ur4BHvFzBzygIpBu8uuPcQbVTs7/cN8J+FdqQI4L+AdiC8/I0ay4yybrZh
e3olWrQttdKYX/qvKu9UYwRYpGwQyGXL47TpLTqv1hRsnf38abXTv9SdlLIBML+j
ZIjIJK5LZSkpH9PEwwxoIR0GY9S7KueuI2JboUGfNwFuYibxdgo/3fkl8UcXa9fl
sizCCp5TnH9QuESQGRXwwvPdXnxZf33j5zAHyTeiuDmBxJwDEkM5GqIvVEIAzA0c
WcvqgjRS+gDCyBCXl1Y/BWvLvERBtHuXoMU22dkLK4W4Z731QYNyDTdZhcnr+a/b
um8qclcVfDLuZolDfN445tRl4FjPHDJvz3wP71kp5i3vqPlJxgF2NqSlr5T7jbnU
fMNzHi1G5cpt5C1v1hLESED5/3kq3ZgooLam4mjAHStB6vlxzreZ1GRsWr/N6ALr
CnHoqykJBfdJFDS9xQ80qAw5OdiwXTiLyQ3KjnwoMz/ZnxRGdk5nuD6WL1oWk33o
6gE8XjfcNLZgfHcrNG4ZW2FDaM1tRrKl6bxbp3BD5kGrMbijsNpaSgqRHTs0oik4
kGTzRn7onp0M7xKT9fwLM18rnugVQBozAaNk4MMLuOfQf5eZuCxROVw7jrK/6K21
1rjTIITYhvsbUoQeaB3pJ/0NR/TBn+7GmB5QYMbyD2icDUiNHfRyOBRI8Zj0i+fD
+xnODAP+64E4DVbaNzOF/k2y2COkoVk0DJVrKKZLpYDiXzkikEtDucYqOUBYfhc7
mbYo8dcIZiKa6h/n3Wc1MRt2nZLRx2GZTzrilx959d9gMcrSTjB8M4cblh9DYP3p
20FkvXJdGOG2i3eb1PHAtP3aEuykOCp2vEn07lsA1Z1BPqBF/prSzmqwOHOXbaxT
nhsYa3AxqXreEzsamPiCe/spnkxwLKz6js0qS/SgCM/eHkYZ6tR0xzeyyw2OOO4Z
nnh0IwELZCpK3Sa7LuTnst3xpE3BYaRi2OdesHS/gCCbiw78Kb1MXuhcTsvZRwO5
DAKtTR+SJO+t+nwQ0/qFYDQfrpRNKkFo7+ANV4fZzCIWY4/rEJKwIIc4uow1mgwy
Uk2IhoI+8E6cnNRwFpiL3YlQfTA6j5slqKrrdBc2SvBHntmU3NVrhNr8OZUTqGeV
fFvKkMR9+y7C5Q6U6e7nWwCtzTVJAj3D8yKXteRBbriZXEGTba8gN/x7jy0X1Q4H
TMiqCCZSaHgEOVD17iWD/K4S565GmGH+B8w5LwN+miYTFAhOqmjschRLfXt37jYU
`pragma protect end_protected
